`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i34oGvJMIw6GlfVSxwLNY8c372uKeSWECD71UIK812A9Z8w4anSI8GkzK7nFrM2O
kw0q/2kCyJCfoD+4hLewT27PKkBCEdbxGXPqrwDOiQylUGdlaZz7dSoa1pWJLJ4f
0JnKsT44DL4WVvMk7hrQn/5fsFpec4wbkU0CvFH9oFjzOUD6FfJWg0JdENiTSnNO
Skhj+KZmvDBI2io2CgcSPmIjbBr7qplLbHpCgAm/qE2nkHhiGXtKwkNQ7oC8ngAw
QG2RY4dlDQM7saXdMaik4mcQccUMoIfHeIbXwLSoWE6GyLCq8oEBsS9SR9KQshsD
6NNxZp7QLq1CHovdmfqjgaJKzaO3ZWfAZweNAfmk7iFv/SLmTVlT4WozHqtiZnuL
Rk1rPwxh/XiXXyd/iIQ2X99OUkl3qFNRl8GLmdIhe8GS815waf68+dBL7rvxTHI3
/6SyhBBLbcM0CvX3oZoXxo4y0OO4vMQEV/zQR+mplQ7sk1IezUyLGXN9b5j0cGGG
lBoL/IiHS4fF42XpoJdYyDTYFq1f1KqaejY4DA7j/11xdL0fvZhw+nlTL0lYEnOP
MT4xPnQhw34TcoSJZCXKTWvBqos5YkIpMdPULU0B04OxkvqVBLm25DVaCvdipS5z
8a1YhZW4CHoSpwm/mW1BnhdVn5Thznwp/jNYgvWdJsqBaqx2SRQzLIWtc5Sgs+pJ
HIVmp0y8+g//RgX+QSL5r36jlawcGp9NNl4asTp5dJB8NnsjEczyijbPbOVkW519
3Bz6xL5oA0hK7xF/gsiF/UvPww3ROs92sHxzADPiLMXVB8ReqM87wLpkMOsPSMkK
CPv/ATm04Y9dcbDkuSlmMSwnwPRLy+OeTGCbbKLpE5P8GDvld9doO0daCCEkULzE
RUHiC4vgUa7aho4FmrFDwzFQLJJOBWxJbdcHV5uxP0uJK/nqhXN74Jvm1g71qygW
eA1P41MOkw34/vFIoZm5To2kc4zSFdnnVaUlWtCoKmkJT8kgSIV2PPw3S4n/nh48
Nxf6ZJU3udOSTK9e9o6r4B8FkGXQG7mDtQAl8ojuNCq6ZXwzJEuoKne7A3e9ayZB
wUyyADOgrwRGaGgC1/8vL3Z/X4RZi1gizNZ14wpL0ve7rgcjCJpzKrwb936G+edk
eMwMgTVBXwsZ1UV/vA/cYQSmmQgUqNs+5hbrfoE+TRe8N49IvkzS/3/yfCAKSaCP
xuiyWE0xq7u0gw/8O3n+n2B7aK9vayp4Wx5oCd1E0VGTHDwFeTW9oNJLiKBfchHS
4gek6grUxPQDCsCj28hqBGAqxrLVNfJVGU1Vi+nA40K51U1hz2/B/qSvOnUOUYfQ
NOL9hR7dxUoeyuPxptUfYyvZe+pnvFwi31X3WC+VKE0F23b78n5l4YQSxaPjpoup
ZCVMNDy4VSTpvSB/IRlw6Ftle5INrgULS+erFBDgCc1mqBAz3nXmIiOzq82knB7c
zhw1Vgfhi7G4NkJlE5/ExidmgIwnHZ7hsjBV068SMIf9Q39/aSU968St5akklnfb
DiTICvGqTYZfgRtxaliaDalQt5KLZHVSzmJ6wzFj1ii0uV9W1nxkJmUD3FNolagY
MfhBBphwB6hJtE74s5DhcFBTnCFTh3UnVCRjOBjnc4o2fFeZRzUaPolmxTjlqJ8G
oVGath8pHVKPplzas4iunfQZJtI+sAMSYd6H2LonPRh5xHWziDQS67DibzBQXu8y
ojerXzZwKEhpKefYdtIru8PLEuWTN+q13NiqafNEFPK4M6pHYkyZ3qqZ5LVkduWP
nmBN4gUgM3GJXyR0DiB51YJmnz6mt+ZR3hisP9F8y0YyKOY+brRbAohACtTv2frW
7W2ISczgZAVR76nBvr8yyK/shVECT/O58QC6lhffIusd70MnHfuilUovCLg5wTlB
GT+xRhK1rt5819IzhiinwNB5hzJY3/enMMveLcjj4emue8etHY9XaEXlT6GKH+bp
8SWeyWiPd0IjxpeaUXqNLBdj9DL3kSGc0CQJBxZ+3ZiqM687AM4uTJCQyoNbrMSe
vZeirOtwE4jw4/e/qSq+JsKnNWDg+k15fJ2vDyBGMFhZfdZlbLTttfUZHvTMeRPE
VpF2+tb2LQncXOLRqX1AV2zvrlPnk5s56EVcmpUZ2HgTn49O+kBnk7A5csGW5rwm
cRHkoCaWwRX8XpRcldNSBze+5wRrKIb6YO/nHDoOqAoxovzs+To5as+WdViQVrpM
VtbCbgmP99pjyR4W04eIsjla4WYr2JiApuaHalcqWTHavHZOORwS/JULN/71nG85
idMjQFgSMtwN8ZcaYve/2SQZO1i6HiyJG5F2gzl83Q3vNY+MsKnvVY0WE3UWskvH
WyY6AO6vuOzfxW6iNFxoX/KyawZpRPbMp8exfCbbYnjsCzOGJRpXgtpPmuJhAYuM
yQFpXE5gz76zsd9GT+bJ1JgYEdMFOR486Wo41dS3HZg5Pg8vZ9x2wwmYPv+w9QmY
3sM43J+MkCbbq7Sw7ZEAwxoYJqVEYwPW8LT5bd2kCqmUgeZfJaFPDP6BOvzChvVW
izMqoQk7pOLQyY2UrcGh0TV7ljqm2SLw5/Vxjy4aZmOmO7L4mhfYAANi4No1HDbC
nuJyxBmDZ7HnuUOUtvzbcCAxxAzTy48S2APTaWGmd55PBFLB2xDW+W2p+m2kLMex
vVkZgEbNMFPsEzp6V8ayDgJWSAU74xJI2kF5w9E4VTEgkaO3Z7dZJX4yGTw8gVj9
3v6fm8K8Khhfsgj0s69MeT8gAkAiLqPd5yFO+xY4ChmH6V5jATydKH8lG7SVEBLl
qxnTotjQZ6y9PeyovpJQX1im6Ijx5TVohLh2SeYEejNbp+mfsebW0Mc1zBfn8drg
Uhq06JwKvlUC3yh/f0Ve6DDitnZs5uE8SLZiad76z/XF8Ox5H5aVe15u0yhhM/eV
DhsU27suJX0Df2l34dGbb/sY9cWXN+NQK28hoHfcqhjV3HLlJlTFAFkiyOlWEkWb
TpzgRrXvGfZVtd+s6sxfwk5JQbVl+gZ7lQqnt24w8KcxBOYP/+7i3apmnCQeE0GG
F1U9yvJ8dSJHyf5Icefg9QuNjzKzy8uo+Uc++sEELfzyvu3n4ZP996DdlwyLZ7JL
HnLWh7iOjLU90BKsQLCNK4CyinVY6Gwc6gpx7QJjOkshhEMnn8bFNfmX9nchHATR
z4N/zsG5d56aw6Dzagu1Ccy0ACHpuHPWQ5WJF9/vuk57QfL+1KSf5LKifUJFwqHa
zWwpO4U5Osy0jz2DUCxYJOSrloIhca/5kLq9LRoHD1MA69ldghe5s7whZLSvJRqI
/Wc1nwzr+Z0Ic5Aw8uMD+IT3Kqb96mS+MJKfxg5/cFZBc/dJdWCbRbjW6jHxIypf
ni6pKo5a1CRbTi1ZtFrY/ftwYOE3pBifBhQozSLXeK/OXJkpyfPBoPsgxNUyJO/q
/UNpOLOl23WutbvkFGBokhYTFMqe/LslEpsTgjKrAdEFe7tUHwPsMOMvvJGgT7bH
EEBYTGXz2dgg+qpUIl132gk8lNtGkgiqYaathdz56l7AtSwlZckFcuEpIw6AbgRk
gXuv9Up2o6IFGibofkU/69irwPTwSiAyLO9qwC/PbLkRBzEioofeKG9oBwZEh+zy
vFj5AqOinwPvsh35jvy/vrE9qSWTuH4yyf+G6TNR1hNEczaaG3nljQ9vXC/Oa1jo
r0mvTqN0ghI24Tpz/We++e2AQ90Xi0RibcPPykaHxpxUOLfkh3uXUal6mcKh5KHI
13gAXM1kh6ZivOOix0qu5lEtMipMFaLZkI0mISZCqGSRS4LIQ56bvLzNO2vBMXaa
Z7Z3GjMt1f9L4pJ5fsS3+P4Tk5XtmI9nyi1C/YCE9A6ppWOOcee3BUV68SJINogv
hiyhnCRIoJTOGza0Ms2+TAapwTaO5DAuDPSEvRHqXrf1uiB+qtrPKVUIBi6b+AtJ
NL54UuwU4iE32hPWDrVKBLpKzPFshS+wllkMATlE//GfvIbTHsF0AQ7PUGEEuxeA
N6JmLPnCGO1A4V7a/Ep/sOsRnZLyilq+nmZCrYyFeLeLnAbDsrrcLkkKhCod9x+u
Em2NFWsqOiHoHpgNsRH7Y20xovIJlfVXtG8/Bg79fGxrwMATMXMQyyqO6PE8BSxh
0Px1oVpxQDvMLZsE8kv8B5TPXWzK7Roit/29iBdoFSDwQays6UkGJGeF5whDU/3g
/G9pOfj9iHqLsMejEVFKCtLZse8lT0UyJIwf6dTaZcbzCo4BWDZPi9wDVCwgfZDB
IUIqCrn4ImAiakUyr9TpdjuQJVpvTY2Vndqh/lx1hjxsZVc2IWOWBIIC+qeRgcX6
Kgss/fe7MPltshwHLUx+Co5J/ZMrf+XfSj4G7SOZlYC754HI6EJcJlSOddXPGA8R
QJVCgoeNzDEeeSnpFZgwCjJYwzHXRJi/LIU/M/GBIWhK4hbLAFAO7qE2fneBat/c
Sm5omDf/80lO24tH+x7mvmeBKu2sgrEyR8pyFUCgVkYwuPufUfo0o+BFZb7gm8fz
2Szd8KNHecm1O9R7/OXK/GaKQK+kt2ZrCtLq7zSHtLPmgr9AfmpWjCEC+Lmv2XAr
qn6AFGV+NaNbgE8e/p0IPL8r+k9wx+/93dIyV7KzZNW/JjdF0QcWTIcUYy9qoNCD
2YSD+A1GG48gv0JuGx/NVnkoLqEgGCJ0qsUwDqGcha9oOuCiWcTEKKyIESwXnSFi
mS+j4Ho9uHaMH/NOrwFR+pawdeXQ6vlCsI74wJHidsmod/CmWkXMosuH59RNe5WG
laBF/6hENe1WwR4ukr97cOnx8v9fWrI+GgmU3ow2iQOtd/Ypm5lAPzL2yQ/VlMGp
OFOl/QjPbBgIWix+M8RVCeOPMEOeTDhpfl6TJAtdCqtqfdfM34bbpjBzxVo2nWat
uNeHZ0l80rPgqfI97ae6f4nyD6f6f2g5IqDvh8ufAlBFkOxpg7Er5Ekdeek2DdQV
Ut+JAQhkhjtTfvPJRmgaxp6zc5Qw99kwViDiUOMPjWVIw6dbUVI/dHaMO2UPBWt+
4l2jY1AUhER2BMK/K10fxP4dtFim/qP8BkXkOGA73SMHmIilxZewK2RYyfiCb1us
XPtQRNq11U1JKEd4Ey7gGRLBnQ1c5HvrSvWSXSr/0/4vnAKlHpq3pGE7HApbzzpY
nX71xJgz45iZmbgw9m4HE9IlguNZqV12sBX/6BKa/4FOlcSMT7b6mFFMoA5MJiPY
A++LwxH86yWANypNcpilaVh5VyazqKLaEbG7Ab7QsIWPuNRtM/DfhGwrZSl2L+W4
KEPOQCObu1WpaoXfTBEpG8nt9HtPF3cR0yXM+jkOUI9xs22U/BBGfHSMNXnLkIw1
UO9b8G18q4exoAUmgLPWF0yr0m4od1vt9FxJxXcYloub1Q5OKcJ7DURppxY9V3GD
//snGGpRcxKFZWuODaoGfuSl5BZi3N+kfscpIPnWXpEzj7BENNM0pJEUGymhpUJR
pIiiRCltK34nIvXZEOmhEYO0Yik4P796T2le8sgPKuK/+iQ7ANyK/V4ZjfxF8Iz3
2ctg5qUwNewppoth9Kx0MRRg3Hzm5KlPwou/BYj9yu1vVL8ybcVBLcRxwqGol8yx
KLIK5tZrEWbnLN/v4IRxcj21aGaqlibchbX7RzmkQLM3qwi5boUT5XjAv0/FMWWv
OxF2DxyoxLAKqrZMFF9qh9+gffaGy4VJbjPR0VE5Jpyowaiyh+ZftqqeMYWym4F4
S39pR7COzF5jfwLgc9lxMGfd31PgHWLoF1V5/WMdDYNS2jA/+kJjX2TVG9eJKfJd
li+hjhISeABarWpR4P2g+PfDqZVxcdWDgFHqUHXkfrUgO6/+zEpAvfZ7+9eyFCWj
v6N1wCNwHSd0vjaFQETGE+g4lgKWV+4gn+Z2s7qz4fk6OotYy44ok76oo7FPmi7r
BLjVjfP9tfOGfCDw5UOt3iutmi/Mqe6sAqJ7/KbZjWvziZitY6yQ7S1ZHVhciZN9
UG/LLi8wqDRq4uyGeyRoMMXy+vX7dKQnmcCb05Gotp+2JT0v6CssXrpjcnbtHNXc
EWhzLrhkBRWRcjnxvYUNDx7TCoOT9AmbRZDp0dk/4CmR+3Yr9E18TLRiIN1Nvwf/
5bSHSBfhauK750gUiq9rxr/MUu6zpxAPGNqZyqj2Neu5PUnfcy4IaMSKNmEXvb7o
ZBcqvvVdNw3PTjQd9gLp5RKa8C0M2d9YlRXnJlkqRV03ugqV6spmF1GQNVLCBfhl
bE2PpjVLoRK1I2bQ9J4TykW5NzWawBL9H/vBKM2vKGanVi1UDejXAqB1M+zp0KqV
dYdjQkyqH5ii67KoqMVNC1v/hewYlchbfvjAetAIJwOJXKuFbXAozw+gk2jsktaC
XgJfrZhuLm0kNcgdfEdr4I6kYkHMKTxL7ca5L8plDRodcCJqPzormAjMrtknzYeS
X1kOBoyE9PJ89J8aM4MaUZAanbsuUp3VztbcbjpSNMh1hSWMV4/pls1ZNXZAAd9n
+WZZjCCfUrzZPetUpsVuNqrdlcrOHUP0dTYh2tEGxUvfBvS7wL+YoKhif7zh9TyB
5ie7yB2Ff8kWmqqpseNZxdyvOEzPwy51swpve4+0KScfUvKhwYj4z0PP6mJnX0i/
mtNfI/oMMv7Yxmlj4XBWSQY8T3CVkKDEBnZ6RSXwAJtLukSxy7KailZ66NaAtflC
8+u5YyfTyO3oRtRSweH/l7MYzOuexCvfZAI44Tc5suOWBHsW5l61IgHbqjdhWk+w
a5+3Fmha7qNpbbeJFx6VqoqtWMvalsC1GqTYsFeQO9UQTRNvJhwh3m+vfrmRbo2i
7OahGRORkhaCw7W867wpmkoa2k3aPoqlSraRvMoIvNch+CroWeXEdkU+f36jLVWW
ZMYG6CesQoTtA9pS6DzWZWvj5zjjQH7ulJVGpkHU7DmJ5cki/UGs3L4SD3DXtxWt
0/0ZdALyFuEJ80FcY4wMwm+FXAaWAO0AAFuR2y9QPgp2blV+pYiiMC92aJFeM20z
LWf/j/91mW9ngISVlEvsIUDofoG0RpeVAUsHtu0jXgk4HSQyswnux+jo0PAp6Dpz
GPTOL/xB597MTqLpoWWUjIhFZ6bxF0TJCcop5DfWBPMfXe8RJwFylYmAGPkOqWH8
oWcG21ncF2dtKtOVDbELqykTMVo6FzA+kR03A20aHmhVlCYAoWtVat93sxjxmb2+
c2XK3wk75Efz8WXFiOXBqnJGAAJuvqvuqd8Qa7gRns8DTLyR5hWyQykYClFGDeYp
9BtOtpuatsRsRMUeXAsHmERzol7JBP/pd4IPbALEhfevMrI67ZSLIo+Y9aRKVMjq
umMttqRaHyr3bPGHTGVNOyHG7IH4Aw1VdN0vOHqoEGzKySHTZxEz54s+d9mxP1Ii
b/AhLG2isqeLtzkKkdR1owa6WnxOQOIs2psiwxaYCdDpM5IXsfjsaHC7eUiw0Zgz
uH00u+aHjNunA41cnHFGn6tFIMWI0epBfNrmzClBR/Qc1z4fivkq2+mbR2NYD8/V
I7wgiuilc5FK0QpKrNKSh6ONh3f+K5QS8eMrNDRioGt2rQMDIvTV9TpWrVXqs4ql
IVT7CWiqUojM9jQ5iMlVl6Hs1qC7A9KUeyafDBk36Hx0Uyt0LRMzPFU7a3SMbxze
yXTjYYTlVrlPtlBxQVgdqpYlVtzkHT+9Ngw5qqtilIg3iVWJjt5yfpBiIWx05z1V
myLBXT0ug58a2qHciBOntGAnUBA2ARqcAILtwn/F380ozzys19Vp2bpAisgXkuJy
ru/vm6NulwY072gEZhfFXfF3PRPrhwKZxXfEbWl+FafT8LRRGZm4v6SP2KdS4CqB
zBiG2AYMbPZgHjMhhS1byRrQea5TkJv6MBQ/QpGSF8DmvSDadn0owA9R71TwL/Ng
vYTGQx+Uta61a+9vIfv1WtaQdzd6J1tGik9anpTyX/e9ub1K5OWXkJK+Lq929NWf
u7xjicysJ90M8U/jAMBQhqrE3tacpoAuPM65JVxI4I+YIbKiHUdybWkQXgLC/ogy
pvxL6NfbCWIugftseBqTKTmT5yLLKnjIjHPIRcRI8eDYsurINrlPfZV5f8nI+TW/
CVIk2tuzU3NJeR+ioYbkDTevRZ5F7EisoUkuft3Kid1UdhSRG/n5TZERoK3ETLSt
2a7U6SnHqvn36z1H+62r323XYUibY3TTHcaXt8akAkt+aBQf4J8bELK+vQ61Q1rr
`protect END_PROTECTED
