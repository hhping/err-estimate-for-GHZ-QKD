`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nbJGEJ+HgPied6wYcbEMgBcCH9gjz+gquPIa7nUUGBMWWH1pUepiCXgsikT4OuZ4
knLWFUcTcR3r7/wGOlkMp2tr57NVKqch5+VRf/qkUdeH0ACXZh9u3ZnOx4JV2bIL
AfW4vqPofHhSVV7JE8IXmt5psW6X99kBcb4OKpGZrKbJDFsWtn6gBlXIf9SsrLbl
FVxo3f8VcoO5+HKB7x3n3pOpQvVNqUw1EPGvYG8FifiOR9tC90x1I9p1l0nRsHHW
EvIJI6qxFwAAtxl7IMxLWBpf+ZHzwdCI0TUFw0l4Xg5+OwrABC35LIl5MMqrpcK7
ZOLp/RNdwAUsLwOi9q+VwO2h0xm5tP6TLLjxbAJRu8gbW6LgoyoIhmNiuN3w7zvZ
RcCQYKYRybfq3pjE8K0Njv8x4rh1Ze22vovO9IKQYp7MsFXDH6NuE6C4n229s+ms
eLdV8uZ+mOV8MMEFxcyRakBSBPzwbNgg2+WIS6GJQitNtihhVmSXdcRc2mQAiy1T
+3nFiDwDKwIiL9TjNBtUdfMHDwoSEZoIRZQyipYTUUg6J+x29j1AYTibNDT29S3b
VtR8Xnr94jQ7vrHh6ItOnYsy5Iz6tJfeX/0A5UVj4oAAgm6ywbXzK+zNFQEp5+zI
0w+Y1qA69Qre8ghwAKDcAsuiah5DpGyUkA2RXfLHJSALcsKFDaOtkQ7hBKfOWx0q
TPyotJa1AVo2de8BpucxoV+qu9/wlp5UkktAYHcRhQG9nNzhpXHyBjns5pK5Vx3J
N3F6FlChofMVKjixi25jcNQPpnnTvoyB+8pdKY3obuk+gykXCE/YrIxMJesHLzxi
U0jegcEjxuczYcYgdGlq1VP6nkvpoMGHm7DdCPNFtN6Onic2GW8mJHFr8tYv/0qZ
0t14G6IE8v+w1h1itTdBGrdoh9hh4zb6TEIneHGwrK3EOEjxeYaRo7CTFErmnCW7
qJe3p1rvpbPHYubhHVpQfX38fLRXtVXNvCOp6zLH26CUKvpiqSUcpMzbPorNRtPm
zJlYkzS/YqmoGat9WGa33zdlwe8AXyNjBCcLl9GOc25FpIEue+8pa5QXZFn8uhbx
wAulsGdr1Qg9MJP5pRqpDsV3pseOH/jVuuNPjRM8PzZvDRLPZtEPBNXgGkcG4S0B
5QS7Zo3e0j7/zAttovuuDRX4VuuB2uNID78eV86XlSDFDCGcQ1REiH8Lbo6wo9ad
tFM44I0nz7zc8LOESBiScZoKchs8HF5w1QqTefaYAXuVzBCDxhF49/AcIDLseLeY
C+N8bFMR/08BnD4AI2ltjr616TK3cBJ6po8b37dB6HmKUNzOUfib1PNhxmCKYh/M
6xYWufpjizwGKH5P4MeNsl+YRhYh7LcALY0VUKe9AQnj+buLOw0aGxgFuWTuKqlg
`protect END_PROTECTED
