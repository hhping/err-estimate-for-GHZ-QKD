`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fML4qw2DvU7dyX76AXsKJYMz64Upfd6LJex4UH4GWjJEXYWu0PB19a8YjYuT6PAU
BsJcaDDVeMOpvbAxD5rC1psrXT+u0VJnJaeZcIWLAwKKCzWe5MvliyidNcJz4Psw
yRFFjhHnICiuryRaReLb7Wk67mFuIPSY+PQGqNmbfzapExhd9ewI+5BdUJ5KjTol
SwL4sfJALiK4MpfzKLJPHbHtxrgtx0YexdAo+frN0yb52+kUHbfVRcTgQTio90S0
uvkw3A4Xl5XJmPkvjD8Vj0GRDszdSsDbP8EAjAN9oQm8xvPdbx7GaUbwL+uPnZba
F1DJz9xCEUigb/Ivja4K1ayXVTL1Ku6vajNPVdxi4FUM6GzR4H75RNdPJ49T+r9l
jPKLAUnhIEK1krewDxj2KMRQdd7FuAQDmPdQGBrGwD5QQaELhVbIVCv6we2vLGzV
DK1J0kOgIWj28p84L90t8skNpsMoLoq+OYNulFVwrbFQo+WjR4kKH3zTpDo9SZBM
5QJpGX6SSshjY6I99Wop2noITTI7Nu2aEW8y4Abk+cB6L7ER/mM+U9nxIP5Q9RNg
2KA0jWT+G0qoa07zsQ9bDdFKB6HH8z61WjJH6QlfqCPQiKZwy9MUuX7RMW9XjFMl
C25Dbr4AM4dguWyGpbSp0m5tRWNJ1Cv81VTRlEClcO1HpluMQJMhO/LkTKwQ/OYv
KFBmC5ZmO+gcrwCc3pU8H5pKyOrtSAiZ7pPHZIeI+paV53jjl/643H+KiPT93vw0
f95wobvCvIReZnwKL1yQbi0QglTrYgWy5v43fpEKEAqNZsWnAF3p+7vNIj/7eaiI
3S1BKqwv9MiNw8Df0Nw1HFuUqCNRBemFJnEEXc9p7BC2Nqsq7TI/pnJPp+JNK47d
S5CDnW+Mfy2TX8pY6yNP3dw+hvy2xRMETD4GrRf/n7+xLMoE24auuvVVz6VVGjyG
x6iAYLfbBmeqUBrSnUIhMZrVhiubQoYe2A1YcGrQRYM+gihXk5OXuJbG0Y3J51Ae
UnJChMug0UU77WkHPR7fkP5KHS6gYAodIqw+oLDS/lNwX/SuEfARfLBiHNTH6Inn
Xey2bF7fpd+t3xEly6LrrDZ5lEBaJiB5/oMbWwtvRO0ZPZOesbLpR+sWKOetpHTO
1pyP6Khlw8ITZEQbchXTtl+l5OAGQW+nWAUnRzhLLOe1u63NzJ01iAR0BXyK7ChX
O3LVU48tqmlDhq2R8oF1cxg8+KHRPNIkg5mpP5glvlilMTdoOFW5ymEaHZLwRc0H
KcBurIzLtrvbgvv1OnwZQcT9AoDZ9eL5o7fzCS87qxzALh6N6wBysOjKcvcifkjg
CM1EEPpNjKBTc4nZiLsMTm3WQ3jAnhkn3aJA1kll1zQufSHByIvq+j4IKyB4TEMB
wDko8iLput9duRRvFKbQ+ONSBPskfdCYKfjbpHZvcQGePL7SfZln9jej6qHsDnLA
z1+A+jHSmBij+ArXv7XtUkkjNHPp7vt4tuKhKGvcOqXTZ5Xtf5n1kWcrg/kqBOK/
Bn2tk5xg2ka9ahcNdf0lYl/n4jhX32zT+y+KjZmQtVvSfksRkne1eNh8048d/cpQ
PpRmfk1NsPJD4ffmw2ihN2RDcEO564Re1kuYlJXDIFriCjoI4lIbOWCaOCfsytNO
hCUhKJa2t9dRRMF3tM1YSFsNGcMoateYGAA4HofE5j1n2mUfgSrfo3nDTLjJyr0a
6lnAZhMT0pFgznM9Ngf593G8iWAsQna0HnzMzjHr7KP/zxsWMkyzfe8yaXjXy1Yr
+7BjMQYbtYST34ApAuSpe1ZT3x5BIsx/FWJ7akhON5P4r9l30eWlQ+QjTbF2AdLp
L98OBcfdhfI97g7CRhoNmcAt70tTZtIvBgeTry/CgeK3gV8eBdV6P8UoU/7RBm8W
fxMoKsCiWl9X/CyXz7A/tmuYGE3mgSvb/umxbtDyW/i4FuBT3iRtNHyTkYIKOLee
k/tXlJF+y9Q3npa4FRshUCe7N75MgZZW15fBHrdXqTaOyp8iAa94U75RPa3tilfE
vZ2avZHJwYC+hxeq6ryeaoLW/W0u8me65PSZyoWgv6eX/si4otMzlZ/UyVz3XMBA
1clMAG4fFTUrYbp0QT2O7rs3VicDHywSSmgMCeyQwPZp/Rlw3KlKfspIw9Ff7A8e
NcNdHp1fYn+W53QyHdCUpogt/wm+jYJvGCprI/PnrVQMUaVstar+vau1XdpkKJ+F
U8JZ87kSgs7g6BUeX8xoRsdubo5CebAhIZW5bBfIAUPDiKoH5e8CoRtx1kW4NbcF
/Xkjg7jTWwCDUNkUTegr3L1GKngoms/bTkt6o9426aiEN8XRrFuWEgPrcnuaoZaS
eozUw7DGGx9bkdNsNwq/hRx5NIBLkOVkn8I8l1HY6XtGTstywdtbWHt9Vpqqn0Ye
/GdO0UemJuLYG25tEgipk6Jce7k4wNM11lq+eWn4n3UCq5HZ2OwQvCjlFw07XGXV
7bYl9MGSP141xFF8Rns/aM3jAjoTqdeIHUu0lwL8nvndTn1o175xg6iqSjCuGYBP
bax3l7iBmNS+5fzXiPrn6tN7KLtyPilnv4qZyr7q8VvFT7DboRfXnF7zsgcYQpE5
vuMdv6OyJzSd5Zdy7UTznfyJddMZzlpNxl6/je7UUp5Pt/U9OnKrqxzUFVPFN0U4
gn325pGo8NkAVvYveW8B6IEm+LIGjZ2Gry3S2HI/JW35SW5zkraHeJpN4FwfRn2U
pcjFukEEQlTCjWfewKFBMDbWGV/5twW7F8fwXrygOtoWhU7vgiKHtHg6UphRogGk
JKA15KdnQ0DJ+/XSFclfRvyR3eFZEEKpHlLg6IlXhKgFe595dFkCgHlK0dogCTio
OJ865i9UOp/yE7fzgYJrIojOQR6xeEOqDNl4bahQo8Ls6kXX7jAHX5U1c4iN790i
ybxYbnF4RBljNZO0MP+F6yslLnJurghznGrf5CQsWT+b4QAEKW7G2DcNkIwB41Z1
4yXVAmfUzSSCtZc0jCd/jAC8XAV4TSPBEbGKQOTrq6jDE8mS1zH1UfBYZCG1hpz4
7tlUP6DsbUha6n2E9bGmqxMfpaYpKP3a3NisL58/tbLbXy2cW+YunAXcqz0CvNPi
Bd6Zun7eCvG8cLaFEIXzAXe7+kGsY6I4NXeNdvDil76EetT1CuD7s90xoi7zksrD
O/1FrRWFXePqLtP1uJchFT01nvlVdRkRdouCNmrJZ8xHEckBcP2rmVYucbOndQ9C
Ub6flquWnXtF/dspq9MQt1HVzZ9bZAl5jibbzCi+fTandisHruech+m7l9lnKzcG
ShOtCi2UsmwdO3fQWZ8+4fbpkxQsSwP8yjHq2iUOkQ8bUgHq7PRISBtRVUbGWxCO
FbmGA6zS2SZnOXR3ShoOf5oBBkm2cbzymArbM28StLUVhrF/THmsc4L4Ef+ijFUp
ttxUWGDNnVJW38ALNYwYqYsm/s9L0hSKqnYAFLXBij7F7vKJ84OvzxnOvcOHMqs8
H5YofhFlxvi98Dqrk37GF9ZtK9BBWhmDpybj0ZVhPn88rJ2JzZpXpznPcmc3Rrwy
obP85p0YQxARe80xppyEytUmFvNV9xsLJVVurP5NgeuJZ9ibqz8OHTX4xNjW8DSk
ZUdgl4EFBHdfHpbbpd5X+V/d6XoYXS+VLWsZJSbPmWFSr6WTKJuJBniwD4W/pal5
sVl0mCxeNySKbYmNsMytJ5IP7xzX90z0yf4F3InA0luaIUUsU+I2+6hQPXBgW8va
AGKVrdTQi53cFVQV6yW2NEalyZeG26S2f99k3rO8zLEw9sDh5RMoOPWKNyGtgvWf
HBZmrxBmfaPtE0GTTPJiTAD9//pZBTsbp1Kpjq6DPUK4DYAgLURvAk9Ihv5/cBsD
kir1FbcRswefSPqgWmN1pXypHgVyiAODDiX6Tn49vDaBcThn9FWNCaU7lFbPjxmI
zFCdQyK6HK4+ukYcYza2BGTW6JmouVlIPHuzcmrot4eOKwgRO7QFRYnVB/+usPUq
ANsXmcuv2zKyQB89D/iq7n223fIB3wBo7158WbpEc/Mj103Wz5k7b2J6qBKBHFdH
fX54iCMs2m98e4tz1dVck4jWNmGNMAoyw7m86sOMsYz2rtWMoF3swVGdn4WErY6t
d9M7dOgpOOYS/cAsDUVp+fdRgjqDZoHxuPwwh4yZLVyS+xmjtmDB4EIzkL3RTH9i
FVnl6brMSc7QmQQpJCgQbQ0N6hP8TUjeUD0vUVn9DHxPZk44w5MUww7E+AkB8oqJ
lCQABm11gwBY8bh1Wv+XYPFjkjN/w6YWe/GbxfsRclK91d/hgHK554+ydPSiT5YV
aA9g4Piezu9GK3g4aPWNkfiF0NKoBzZR9EvjKVqeN6oflDQ734qJY0trBpW+zdY9
51YO3abjwI2KKCeFvmErCslosQZ7BwAQMbIJGU8O/eiTmolHQFAzILWBk8rshkkt
87iif2HtgVrZuQPyynI5dV7yFlvV4h/ue5BhXsDSiZZqIsJCNTC/il9gbRnBmIuG
5js/bKlWMuPn+Ulg5iRovJdwAtjvzbdk2WLCI8E6XrTtKzLZMFLwV/1uM9N1J94c
LamjoFhYp+btpR8M7cNwInMcBSiyU0mqP934hBrrXUxFQOl9/UWRkjLfofVLtDL0
`protect END_PROTECTED
