`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YUXiL3LTGYja4m9DlnhT4ilpqlo4s4fkps4wuiDGHBXm3nAb0jYCX/5w6FvMrznd
IrY39GuMAUNjv6T4Ar5e8bNM1hbADF/encSOn0EKFEQLtDzM7i3UJXG+x3QZgel8
M64fETaUM1SF3o37SVO7lRsNqWM5+Q5wBYzDmfNuxMTuKSHfBGQXMq18ySyJrsNz
4TLSUjamYRG8oOY37iW88TGvSnJwXSP5fb8vlUCz3ovKNekXqStkqSowQVswyKVT
7ngQACAnzESfcgKP9XggiDs0o1rxvACxAPlFjqCt3FiN1JWgk1oLLPs8TfWiiu+B
Ugkn8uI3DqwFagE+FdkxLjBvvyWIxQNyh2BNLZlX5xBJo3WCkJ17Eovh6pNwb2rh
SVi99wsOcsIFFEfJ/DBgMdX8eKCkX2gvFy5c1UJyHNr7RxAarJHonKw1HrjHqbLP
Z7qA1l3/XssaMESkO0GYWTfgtGtEcHTDfNCFUI3kCD2te0bjQ1zYQlxZRJZetyN/
/nH6N6DVb6Pe+jv5UpaXKyYcDNyCsrUKTgm0pDmtSmxxqIsfBkOhn21x02oXpzhR
HNepYAge/6TpZP70SfFAl29BOd9MJc/LJ3lsxnIPMw6BEOnegFDGqGbEXJYODtCs
+Mn6TD+C6HyTd6qGsgpjxLZz1u3RJhnM6zLsUpSWYG4Z2xBFyrmzBeKoL2dOJICs
XDh0E2v1jIRxpuuqYTwak2EI+Et9JGoRq+BvhHG+30D0v3cSlxXvJIAb2Xw8duZ2
/Ijfw/GflQ3wo4fDc6i0obHcvEqeKaQRZzvVkOSRK7CiCRQINFW4EPrMRcBwnsnF
0eYDb+d/YxVadl/kFJAOL2IQFmt4nQx0a5pk4Ad0+BY39z5389Lrd6bhoe/jX57e
Jyuc+Ba8wqDB5sKD21hFURlreuZKE98smRjKtM6i7AWuJPPENZmfLiWQxUTMhxQx
ObWfDJOPVya13Fstq/8q+naBTxMw3GsBCfiyNM5S1H+udtowBaTwEitnMX15BfI0
fhQRY/uNRU89ybxbpSfHEZEPRJumrXWQTE3UIAAUECjfwbh9SnKW/hkjM42KPhQT
fAtwY7FxBdWcTX61MF9hn1GsaYmPJM8xyIa1BSuOjcncr2ifVI0K1cSBLJAX92WJ
xVX+hnsVs6xhlrIUQhqAdTTIJOI8zlsd2jNhr3QVBZydihjokvrYzZ8U81AArj/A
swB+Vstq4G7DDnrgQwb0SNuimHUAcquvLe9qWKwXEIcKw5bvQoIUl/l92S33l7mE
izmBEjy91S+SyuYf4jq1hifR5MRBrYtEWZmoDQwbRHjK29tAlis29P948iQ3686r
8Bf6rw01TzAyUCScvD1hFKB0G6g7nZQ5OzK7a6vBk41DsiCyDpsk/mvA16kMrSwI
+o+aN/44l64xxRHZuN6e6aevGB8/VmC+lh+I9yWS+kpvmeT+zLF7rs1nupZpLu5b
8uQhJFfFeNhpwLQkbIhgFpQc4WCKwbxzHFGGGRgW2NLKqBzMA8dpEG1VKkNGp0l6
x6HsMpIEdnvLUOml5XQ+lhEN3h9HcEq8wUYsZzbplabzMcSZOwS74sOE1csyF+S1
XmHlH6MCPpJseA+GnbeFQs7aSHb1Zlmuo3hqrpCcqpjB2q1O4Le9/oabXin2DHO5
8AwRxHbgELHfT1GLkaTc0z4WRBa9LwAW8VBIrTtaJJhig3SYuIEM+NTMX2SkS0/D
5We/QZK+ofaAdcM64ucnTg==
`protect END_PROTECTED
