`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5OdaJ1WtLDW+VWPKY3XbbB8BaLOlPO/OgwSGFBk6M6E3ZNkZdeXoUHMUrno35xRs
ppFLf5hRuJpgwh/SksU70SCdiCDGj9EqQBGDqMdwY9MQ5S73dxU0adm7QG4onx0s
b8KntNvNqJ2LRZwei/tVUqs0fmyRUJ/Q7Zw6BS54OB5Xc1qNLpZ9DOT6gh50nB+R
+e7Cx1eFLhG3HcMQjETgip38uzwyKQWqR+/Zc5FFx0ChUJTxdRlbnC+fkJOhAmJ5
V5ZBXjjTYmwQLEgpb/xETK51pGxP4mjTy0L83/vs7cBBtKgppESqzO+1rdGDCoM3
Z7HvA4FYsCVUSvkV8cLHUOshU7gLWs6x6oyart288HwBIzW1ZVWqOGvkhb0cMTd9
hJIfQ76eOLvr1PJcREEXo8IQsxCzbDZ4waoE2OgHe3rs8Mz2euqiv6gZ1fz3iVnB
zvhtap5TTAu1Nj2xHlEe30X6Bqrc89JKyCozUlvZVJ+llCZEKVQsJRv2oGh0RgHh
q7NegG+z5eu1WEcsGI0cywDduQIbNNJRJ21jvB1gD2gihlTVgJlDg8zfv+EmTwoJ
hFh5zRw+3Va0PGZmEZ9yS7M6bFsT9qZiUf5+YvXj49/sUaHNNeh5JSYPdhCXsFvM
nQIBVXxl5p0FZerKqO2n7Mz3TCmvhDioRPVNTZuL3Q3PFveWSIYSglBQdsFypKBr
2mVwrchu+BahDkNA2U/dmF8yDBIZI30eK8KClNhaWqX9K5eZvdIdGay49dBcgcvF
VdnBK5K0J5MbW1pcg++jcYR6xtW7bIaFvQnLIXmn+KZq+cYUALd2v2xgGm+q2jn7
AeLxgs7B82Yu+mvoXth0eur1fEdk0Xm+yoEgVhpPoWOOYOOU4AZf8SW0S2VFmmZl
hc5mgepJqDm6Eas+xOE87w+xlfCan1o8xUcD6rGbTl5WxOyP47Xm9yy/MZndnStT
fAOOqvPyBoqO4IBWConfovbmSOyh/jr0TNv8GW+zNnnfTHPKMR5PLBJjiSt07rxx
1bxuadEurCPRkaH30z7f69pqcYEdzVxwqeJQk5WaWopG3AwC4AludecWAMmLuCdW
+9lEdOMgVOvUwM6qT7zN62lI1Avhqti6OmG1/V6bHwknC2uVb7tY0lD6LALlZ+3a
+Jmyj6Ayiw2n0YW3WxrBBkXrdfabjL0jRmeizq7NWEkB19YmDamkA0hwVCwQ1Moi
GEK2ozTW/JxmBqb29NUvLUxDFJH+OFVZdZSByJE/wwk5JuQP/Pkhpmff3ncAJehq
sWxA3yhClj0PH2KrVIuAfqdsJXtxrRQZuA6Lh2rJuK2mxsMB+FSIKNkONTAo+T/t
mGR54HFWW81xCqvnE5bvkz5LowCr3RZVDmcFU+yS65qPKNxbMUX4mwCmbufAWi/0
PS4QolXJfCjP+BzWb2iGI1lEzuFiIGCQGD0gHzRfeNUS0Nxhy4WUor4ZjUlFTBra
U2sDZUPrDpG/OdKMd6sSbrAYYE7rPe4vb8T8sr9OXp86G/Xzay9qbBcZ3BPoOuPO
8W20vAcMpW1JBEkcYjLGBP0+phhi0POfuqVPc6OGqpeXOJXYsXMJCYna+hLpBpjI
rgPZtgzqsLE7SPNO44YQdgN9Cmlb/YBoxP9oJVS6+SgNGDP1MvZ2oiz+JuL4CtSc
vynEFSwSBZv9NvQiYdxjQUXer406vepb3P2hMjeR6vfXWqwhp9z2NvGMlH2m1kf2
3MKhnvk5Cxn7z2hzZJZOFnzDABDvi3G8Y0bokTFaxbCfa3yFMX/pf3pEkOkBmyo9
mIKoHH+28PMWA4H7IERNkaJs8QzLvR10CLxTT6tJdREastHK3biWA3dL+TjEAoA/
UipAuulfMQGZyyPCl22qbOko8neoGRWTdSkI9KLHaJ5/kI1O7dwQOLqBp+mRDpsc
vqJse/7SbuBJ9hReyXsUPzyY1IpDt/Fb+GihdpovKInp6dupdpZU+/saWU2ItTKM
VCTqN5l4BnJEyFt3bRSBtbDlJUYEAluOMehQC5/tFl+5oK3eIdd6Xc/jJfvwHEI7
EBe90iLMrnFhc3pL+9yMexj77jyKMJVguxmXEZycuN/ECe66AeiyKVtXII6zKeo4
V06bPlAj9JTZwdvq/B+fPAoF8VfhvPsvPUbG6HbIRJRCaqHPD/TtYw5eUwiV3IzF
4D2AKZ/0QKdKx4ETzMPssjtHqzpjDVYoPTMObRXh1DCWxXo9q/tZRYsWV/2SM6Jm
AlglLoFByWuGMqiRaenjXN7lmZvN5O+PkOGMmfAmFOY0Q4+2Yd/EQZyIuyLn3By6
6qyZtx43lqsHouqN2nSGKebBXzsCGLz0kuhYEQWGOBizmH92La99h0C+2VdVyI9I
PJprfjb/EJk9nBQZkY/zlbuhxqMTVpF9hzVmSA/REO5KO8xJ4N8XlLb8TTyEsGYX
XxdFcd482tJBWJjBELRRes91qgp7YKukVSLWhndi2m786lWNi43Q8prnysgwoySV
Ywp9rVhOzArWuimA3TK675E1+YPmm4RIBh8JrivHiyhZugXLAlHlejBDZGSsVlbl
UQoNnugCFXmd76pdl/WW4VqwYEljVXH3w3h3tKiUlHfOgvjC1VsubhooBc1VROL+
8jko+DT3CLffxmDLMG6cERcQzFaZh63xag7ShbD0iKr9COQzGKNk22yUP6HXyVB5
2Tz89q6u8hmRT+bIxtY6XBRMovzNpPifGKwRIHrz/W2Jwtglu/Ep18UwG5k9f46G
BhW4WsJrC4KbBwjla4IVHCBDIFp6Ww8nl6yE5qZN3niH2k92RTlrsOMLK0FgK/xd
E8AoJ92V1p23JvsNRUsyogl1D1NXPWmvfKdj0RqA/8Dh+fO+I1CgimftemEch42V
xK5Q1rJS0J6lIWYJwiMjmwq3K86LR12Vjf54jr7Sx2RTvTKYNF31WamsvU7p38GU
GlgmSz4oOcor4TGpyF4Js4qeG/2m0JW44ThrjiyLZBux/7rKODqzlpmeJMv7mBs7
Algwm6IHn31bKkMoEcWbxYMD0Nt373kK8Fw/NI08ktFoPjWoQX949rgz7sglPrC9
6rxHJUB3e7n07242l61tQwctEWI6U7OIZcF9Ma9Zpqtcx7MQYJU7tywysI8vmBG8
tbiSVjtFujIMkhxsMdK/HxXDI6e+KQ0GMsYTMj863BdDWBQqwzYx6lCjc4TVzbsB
8pCSMGmJwZjB1PJkfiUeA1k/hAfuAIE2S/ypPZHhx5jwTiiZ0zVhzAk3qBkPO2j3
wCGJvZt4CopC3Qm2gJynOjjfEIvJQ2F/2HWe1wI97VTuKxe6xJpqjaUz1P9VyTFW
JDW/IOO2Q7RmuOmdLBCRMG3SfEE2CEbJlCnMIvarZ4sPTo2lWTXWzOu+OZ6F/WfT
W1wZWW3YOxmxmIG/OF3QL4fIU389V/lz0iP1wgCL+3el1wfUM+ew4lhWGKucClbM
VxiYGEifwhIxQFRv9xGC7PWMenz70RIB51axUAKj0vCNJXs+O7/TUnCojIpHIbL4
mIPHQYefo0ykW5OXtTEdR3UNBR0QDVKALTLY3x3++rL4002yWylf5nEsKsyRV3Bw
pVZqXuAEi1kGbiMXYd0IA+bzsfqMtHGow/O5SAD3+ipsGaUcEUQWKLvbxZaMm6Yo
XPTXWFIK69GbW3A/9kuwSo+P3bfrheXQazC/Vq+cRkDRoMRpf6rC231/oOjxhs7J
gOcD0BQt/34+NE5NjRSy1zqE3xffr41lWpL5kTvS7tJ7iBKOevYEd3WIrjNtxgNi
kXzEF0VGa/Jlcsdfm0yirs6s2vvi00ikRdymdxl2Ak54csj0VxadzFpWVvE/z0TC
M3vynTRsOocTnzEMHS4UodDXpHUZK2PDreZ+qwdin8rKW+lZ1n1kXJs+rlDHO8NV
EqVfFKJryyY7TVU1wDOrHH7FthpAFyW/VY8TC/fiq8yqAunD3jvLEXb9Xi7qCQpj
0PUMN9uQsBmN2jJW4w7Vz4O7aErlAcbHO1yCzhpclfrrK/DzEU1EtXrrayhQ7KlG
ncUgAp4K6d0L9qldSBbvUQBEEgtJwAFHD++9jK9S0XvFKLhxQJ2A7JRFco4FW+R8
KfBKBPWy0IcJ3HBBkpy9YNXzO3SS9JlMDgdzy9768ApYxCPO8X12PweB0udk5Jv+
X7He2voRZSbfVr25USf+xoBLomlvknRFq1ksjFdrXzhr0HLthJkTyo5v8lIdyXZ1
jh4kqXmQ2yCF5tX6VmbSS6QO0K9shB2P31V5csTELXfzHNrcPA02Na4eedjDyMlW
npt2VMja7OviUxWfM9kx1ZClq6ySErmXZgw68RfAEkA=
`protect END_PROTECTED
