`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HTjDcsm4IFEtcalSVu5tfATflTDjDw/YMBMew6rQ/LEElNSkgLGjL0nmy8T4PnMf
FlQtMjA6dgHqfLQqMr+7ZxDXm2AeuXN9jyoYd8EkVLZispCfwYT1xzTM8Wg0Nl+B
pR2S62g06tjOePRU2c2CD5HZZ3PSyDbbyAyZkH+xIxX4Kxg0bjJnsZMbcmxo5VEY
mL0CNkCZ1K7AfcRkGU2X/GIjRJVhbXajIza1bzkADcfyv9w5bBYf5vjCSXWYnNxY
EuzhC//12IKdUFnHJvv/riSk9jFoVCXuItbA+Q/LXSZlvoMwVbBImp1pRk4U1bJk
iuoIcxVLd9Cz2wIHRlwksAS5R8GEVrpP+wcUaRmDZYm//DKxZqz6THomlh+COAiq
fuVv6abWzF+gmvkX/1tJdpFMqx7u8G2i1dwnEXhnagWofAuSUktuWoas9jKdrJTo
4yfTbI1gbPGyZ4dL/U9WUEgQiJbn0TTHQ0xsEIvLWGX3fZG86cp7E0VlbUzRJn8l
ot1+CLED+3eTqJLSHbwruL+6FLZVtShWGInmDMxgVz5biMOu1BUy6OeM+i5Z3sUZ
3cSe/3m3cHU96++u/zHfaQYvD6ZStgP2Y4Gfcw2PCj4vvzyr+njDEz5fZcu8UZV3
NQGlRvtSY9hvofBIZq6aE5fI8xZEizKMwrmBm3aUjWD4xE08m5PO+Ce4QvWEpR2z
7l6xPbfpvO1wahWLKV2WfoRsc/pTB/7U9Iq91pExJsIS8RivFrJbu5tBHM/ldrTB
Dil+bBF79e3lUqJdUefYOUSgQJFmfcq2D8+Oq4L9rR1UeqeDOZ3ZHrSQEaaJ9Sjv
7rYWuTGJ/Ml7HK4C+miAYn2AdOg3gg4CQ3+tb9fvqGXe9fNfUCUL9y3NS9huU2Lh
wcPXps120fCk6oJm0tOZe+wD9XFzXtCxqVnjYLBTLPDFK1uiofmsTjnyPFVPL5xD
9+zTTrHxDBbvBgMmRIjtbMoI19nWV9HFNOHOeVXZtsJonXFgaZ/SQAQ6h0RWvt4d
kxbR2CBLWDJEAzwD1gKwOCcG0tehy8KwavSRgay+v8tzaTFahohqrJJQBDuq+dNW
aqTu+ca0uxdClcmzzWw7W4CAqZMbDmGDpTzhnCPcV8rJGEHHn6DogXWfcvWPL0wU
HzBSQRGHmJzou08/MZOFmSW9Kh+az0DEztECDtXwT+0C/WXtQ3YHJjY63yRkAVQF
ZBfiU2iniWDVeMWFELZwh5S+PNySzAVgN3dsZzuDwXDhI/Y4uYF57pHkZAcuonJY
1vQW0ae3qNwvtWofmDFO8BNJxV7lfjac2WbKbJH2qnAtLjgc4sIzYbT4s8GuukDr
`protect END_PROTECTED
