`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUxJcexD2tE7yH0g59O74HwB86SLLpoPZvTcwqeUs5lPktqwn35/E0By56B2FalU
VDoWTOcNPr6SF/QTe6MiaEOseVmh0gMHFPkoP9KnLkR4P+A7E5eXVsn9w+Du1KVq
k1MT2BZAAUV2CQhkxyslU2oJ/mIlnZJh8iZ91njux/nlNjZEKt7R7qYmX1cRgttE
TLQGsCmMWbg8aiRKGau2zmro2zYYCcF+Jlc6t+fcMv2RmW9/goiVc2WVXUvyh1KL
BbgQA+rHPQTYpMJ+wySP+FfLPIEY4BAij67rJGk46KQbSbmqsQ2rxlSRmnHxsTnH
EyfYoWPAU3bsrFlj5f8uVqL7pDw9VRuUDq6WUbONT9G2NDNCMlIgpwqnngHWSW7d
ifaIKQtMu10YYqzj7er3Y+c42Qe4cTPf1T/4AsUXo1fRDF+oGzZs2v3OOt/Yg5Y0
JIBceDi/Nubjmu1OPHDu0bxsSSL+tPi1l7whulSmBBEAwwKY85cO9pZr+rsAJwJ3
uqbJah7/VJLG526C9xVaGSUZgjrjLjMLxeVF3OwnKveFSQT3RAlT2sWApHAnPW+P
`protect END_PROTECTED
