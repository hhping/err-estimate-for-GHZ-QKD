`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OwRFqF6rPNT8EVYfwxdTMEBOyvqD4ToXlXbCg/6FYZVySbGHUqF4su+8TJ/8zxA0
1bBnxwcxXcl3EuNmVZvwEOZsXHbL/1/zGkxoQHW1F5W66XCWjgEkMZ7ViLOgEi2W
QsHQV/bFrcqLPb9TB7R5Fpv9LIkCoRkM5rIIrsh4OCS1MSooALCX28QbYepV4cy0
`protect END_PROTECTED
