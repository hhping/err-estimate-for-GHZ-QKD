library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_8g_tx_pcs is
    generic(
        enable_debug_info: string  := "true";
        auto_speed_nego_gen2: string  := "dis_asn_g2";
        bit_reversal    : string  := "dis_bit_reversal";
        bonding_dft_en  : string  := "dft_dis";
        bonding_dft_val : string  := "dft_0";
        bypass_pipeline_reg: string  := "dis_bypass_pipeline";
        byte_serializer : string  := "dis_bs";
        clock_gate_bs_enc: string  := "dis_bs_enc_clk_gating";
        clock_gate_dw_fifowr: string  := "dis_dw_fifowr_clk_gating";
        clock_gate_fiford: string  := "dis_fiford_clk_gating";
        clock_gate_sw_fifowr: string  := "dis_sw_fifowr_clk_gating";
        clock_observation_in_pld_core: string  := "internal_refclk_b";
        ctrl_plane_bonding_compensation: string  := "dis_compensation";
        ctrl_plane_bonding_consumption: string  := "individual";
        ctrl_plane_bonding_distribution: string  := "not_master_chnl_distr";
        data_selection_8b10b_encoder_input: string  := "normal_data_path";
        dynamic_clk_switch: string  := "dis_dyn_clk_switch";
        eightb_tenb_disp_ctrl: string  := "dis_disp_ctrl";
        eightb_tenb_encoder: string  := "dis_8b10b";
        force_echar     : string  := "dis_force_echar";
        force_kchar     : string  := "dis_force_kchar";
        gen3_tx_clk_sel : string  := "tx_pma_clk";
        gen3_tx_pipe_clk_sel: string  := "func_clk";
        hip_mode        : string  := "dis_hip";
        pcs_bypass      : string  := "dis_pcs_bypass";
        phase_comp_rdptr: string  := "enable_rdptr";
        phase_compensation_fifo: string  := "low_latency";
        phfifo_write_clk_sel: string  := "pld_tx_clk";
        pma_dw          : string  := "eight_bit";
        prot_mode       : string  := "basic";
        reconfig_settings: string  := "{}";
        refclk_b_clk_sel: string  := "tx_pma_clock";
        revloop_back_rm : string  := "dis_rev_loopback_rx_rm";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        symbol_swap     : string  := "dis_symbol_swap";
        tx_bitslip      : string  := "dis_tx_bitslip";
        tx_compliance_controlled_disparity: string  := "dis_txcompliance";
        tx_fast_pld_reg : string  := "dis_tx_fast_pld_reg";
        txclk_freerun   : string  := "dis_freerun_tx";
        txpcs_urst      : string  := "en_txpcs_urst"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        clk_sel_gen3    : in     vl_logic;
        dis_pc_byte     : in     vl_logic;
        eidleinfersel   : in     vl_logic_vector(2 downto 0);
        fifo_select_in_chnl_down: in     vl_logic_vector(1 downto 0);
        fifo_select_in_chnl_up: in     vl_logic_vector(1 downto 0);
        rate_switch     : in     vl_logic;
        hrdrst          : in     vl_logic;
        pcs_rst         : in     vl_logic;
        pipe_tx_deemph  : in     vl_logic;
        pipe_tx_margin  : in     vl_logic_vector(2 downto 0);
        coreclk         : in     vl_logic;
        powerdn         : in     vl_logic_vector(1 downto 0);
        rd_data_tx_phfifo: in     vl_logic_vector(63 downto 0);
        rd_enable_in_chnl_down: in     vl_logic;
        rd_enable_in_chnl_up: in     vl_logic;
        ph_fifo_rd_disable: in     vl_logic;
        refclk_dig      : in     vl_logic;
        reset_pc_ptrs   : in     vl_logic;
        reset_pc_ptrs_in_chnl_down: in     vl_logic;
        reset_pc_ptrs_in_chnl_up: in     vl_logic;
        rev_parallel_lpbk_data: in     vl_logic_vector(19 downto 0);
        en_rev_parallel_lpbk: in     vl_logic;
        pipe_en_rev_parallel_lpbk_in: in     vl_logic;
        rxpolarity      : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        tx_blk_start    : in     vl_logic_vector(3 downto 0);
        bitslip_boundary_select: in     vl_logic_vector(4 downto 0);
        tx_data_valid   : in     vl_logic_vector(3 downto 0);
        tx_div_sync_in_chnl_down: in     vl_logic_vector(1 downto 0);
        tx_div_sync_in_chnl_up: in     vl_logic_vector(1 downto 0);
        tx_sync_hdr     : in     vl_logic_vector(1 downto 0);
        datain          : in     vl_logic_vector(43 downto 0);
        txd_fast_reg    : in     vl_logic_vector(43 downto 0);
        detectrxloopin  : in     vl_logic;
        txpma_local_clk : in     vl_logic;
        txswing         : in     vl_logic;
        tx_pcs_reset    : in     vl_logic;
        wr_enable_in_chnl_down: in     vl_logic;
        wr_enable_in_chnl_up: in     vl_logic;
        wrenable_tx     : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        byte_serializer_pcs_clk_div_by_2_reg: out    vl_logic;
        byte_serializer_pcs_clk_div_by_2_wire: out    vl_logic;
        byte_serializer_pcs_clk_div_by_4_reg: out    vl_logic;
        byte_serializer_pld_clk_div_by_2_reg: out    vl_logic;
        byte_serializer_pld_clk_div_by_4_reg: out    vl_logic;
        pld_8g_empty_tx_fifo: out    vl_logic;
        pld_8g_empty_tx_reg: out    vl_logic;
        pld_8g_full_tx_fifo: out    vl_logic;
        pld_8g_full_tx_reg: out    vl_logic;
        pld_8g_g3_tx_pld_rst_n_reg: out    vl_logic;
        pld_8g_rddisable_tx_reg: out    vl_logic;
        pld_8g_tx_boundary_sel_reg: out    vl_logic;
        pld_pcs_tx_clk_out_8g_div_by_2_wire: out    vl_logic;
        pld_pcs_tx_clk_out_8g_wire: out    vl_logic;
        pld_tx_data_8g_fifo: out    vl_logic;
        pld_tx_data_lo_8g_reg: out    vl_logic;
        sta_tx_clk2_by2_1: out    vl_logic;
        sta_tx_clk2_by2_1_out: out    vl_logic;
        sta_tx_clk2_by4_1: out    vl_logic;
        sta_tx_clk2_by4_1_out: out    vl_logic;
        dyn_clk_switch_n: out    vl_logic;
        ph_fifo_underflow: out    vl_logic;
        fifo_select_out_chnl_down: out    vl_logic_vector(1 downto 0);
        fifo_select_out_chnl_up: out    vl_logic_vector(1 downto 0);
        ph_fifo_overflow: out    vl_logic;
        g3_pipe_tx_pma_rstn: out    vl_logic;
        g3_tx_pma_rstn  : out    vl_logic;
        non_gray_eidleinfersel: out    vl_logic_vector(2 downto 0);
        phfifo_txdeemph : out    vl_logic;
        phfifo_txmargin : out    vl_logic_vector(2 downto 0);
        phfifo_txswing  : out    vl_logic;
        pipe_tx_clk_out_gen3: out    vl_logic;
        pmaif_asn_rstn  : out    vl_logic;
        pipe_power_down_out: out    vl_logic_vector(1 downto 0);
        dataout         : out    vl_logic_vector(19 downto 0);
        rd_enable_out_chnl_down: out    vl_logic;
        rd_enable_out_chnl_up: out    vl_logic;
        rd_ptr_tx_phfifo: out    vl_logic_vector(7 downto 0);
        refclk_b        : out    vl_logic;
        refclk_b_reset  : out    vl_logic;
        pipe_en_rev_parallel_lpbk_out: out    vl_logic;
        rxpolarity_int  : out    vl_logic;
        soft_reset_wclk1_n: out    vl_logic;
        sw_fifo_wr_clk  : out    vl_logic;
        tx_blk_start_out: out    vl_logic_vector(3 downto 0);
        clk_out         : out    vl_logic;
        tx_clk_out_8g_pmaif: out    vl_logic;
        clk_out_gen3    : out    vl_logic;
        tx_clk_out_pld_if: out    vl_logic;
        tx_clk_out_pmaif: out    vl_logic;
        tx_clk_to_observation_ff_in_pld_if: out    vl_logic;
        tx_ctrlplane_testbus: out    vl_logic_vector(19 downto 0);
        tx_data_out     : out    vl_logic_vector(31 downto 0);
        tx_data_valid_out: out    vl_logic_vector(3 downto 0);
        tx_datak_out    : out    vl_logic_vector(3 downto 0);
        tx_div_sync     : out    vl_logic_vector(1 downto 0);
        tx_div_sync_out_chnl_down: out    vl_logic_vector(1 downto 0);
        tx_div_sync_out_chnl_up: out    vl_logic_vector(1 downto 0);
        tx_pipe_clk     : out    vl_logic;
        tx_pipe_electidle: out    vl_logic;
        tx_pipe_soft_reset: out    vl_logic;
        tx_sync_hdr_out : out    vl_logic_vector(1 downto 0);
        tx_testbus      : out    vl_logic_vector(19 downto 0);
        txcompliance_out: out    vl_logic;
        tx_detect_rxloopback_int: out    vl_logic;
        txelecidle_out  : out    vl_logic;
        wr_clk_tx_phfifo_dw_clk: out    vl_logic;
        wr_clk_tx_phfifo_sw_clk: out    vl_logic;
        wr_data_tx_phfifo: out    vl_logic_vector(63 downto 0);
        wr_en_tx_phfifo : out    vl_logic;
        wr_enable_out_chnl_down: out    vl_logic;
        wr_enable_out_chnl_up: out    vl_logic;
        wr_ptr_tx_phfifo: out    vl_logic_vector(7 downto 0);
        wr_rst_n_tx_phfifo: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of auto_speed_nego_gen2 : constant is 1;
    attribute mti_svvh_generic_type of bit_reversal : constant is 1;
    attribute mti_svvh_generic_type of bonding_dft_en : constant is 1;
    attribute mti_svvh_generic_type of bonding_dft_val : constant is 1;
    attribute mti_svvh_generic_type of bypass_pipeline_reg : constant is 1;
    attribute mti_svvh_generic_type of byte_serializer : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_bs_enc : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_dw_fifowr : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_fiford : constant is 1;
    attribute mti_svvh_generic_type of clock_gate_sw_fifowr : constant is 1;
    attribute mti_svvh_generic_type of clock_observation_in_pld_core : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding_compensation : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding_consumption : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding_distribution : constant is 1;
    attribute mti_svvh_generic_type of data_selection_8b10b_encoder_input : constant is 1;
    attribute mti_svvh_generic_type of dynamic_clk_switch : constant is 1;
    attribute mti_svvh_generic_type of eightb_tenb_disp_ctrl : constant is 1;
    attribute mti_svvh_generic_type of eightb_tenb_encoder : constant is 1;
    attribute mti_svvh_generic_type of force_echar : constant is 1;
    attribute mti_svvh_generic_type of force_kchar : constant is 1;
    attribute mti_svvh_generic_type of gen3_tx_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_tx_pipe_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of hip_mode : constant is 1;
    attribute mti_svvh_generic_type of pcs_bypass : constant is 1;
    attribute mti_svvh_generic_type of phase_comp_rdptr : constant is 1;
    attribute mti_svvh_generic_type of phase_compensation_fifo : constant is 1;
    attribute mti_svvh_generic_type of phfifo_write_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pma_dw : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of refclk_b_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of revloop_back_rm : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of symbol_swap : constant is 1;
    attribute mti_svvh_generic_type of tx_bitslip : constant is 1;
    attribute mti_svvh_generic_type of tx_compliance_controlled_disparity : constant is 1;
    attribute mti_svvh_generic_type of tx_fast_pld_reg : constant is 1;
    attribute mti_svvh_generic_type of txclk_freerun : constant is 1;
    attribute mti_svvh_generic_type of txpcs_urst : constant is 1;
end twentynm_hssi_8g_tx_pcs;
