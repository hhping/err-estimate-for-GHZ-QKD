`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kTDEC+LxFIT1uplcipVvpohbK5qvodvK7FOCvmtFwXEh4zzd9xXQM88j87HOgd3F
Fv0tvPWfQvvtvazL/YyNTGmM5IZX80GLJhN492GZIgS4G5Pzy/scAiWncTM9WwNT
aIftOPSir1XtRDpUoyIoFg3VCeLLxFZepvSQG2GpzEW4aoXA5OAWjWgu3vWSBANb
ADuqmkg7KoLjkA8sUevdeJPy9U2CBKjX0zA93NkpPjzoDQhwxrTVctp4xuRehjrp
pF0rSKKOnK4MCJHP/HyAUm7EbYJZEF1go9JN/LDktm3ipUte8BflAcMxmBZXQ46D
Fw/U77BLjyRQz4k2/RGjB4236+YZcEZCqfpX0EvmJ+NMWlF2snaCApRRdc2M9wF5
GJB3GpOwb1kHwN75i2+6hdNunsGeHlj3Tr5b+eDQihN6b2jNgCfadw1Z7kAeFGki
eMtPA80cQaRkBQ5Ae6UE6pwVunN1WXDdkE4UroqIPa9NAgkOcPtwHjBu4qMcs+84
9I9fs+/jpqnU5rUsl3vVE5FWqgm+9rMbfAkz/YtIOwHAHVpYQCI5lksCjrhvfMWc
5vNTOB1r6Nb8l0mEwt/2cny/TSRhZCtmYaELHN4EocY4gBjT4GfgPkqvTmufQvvi
TZiwAob8tDoXxK7qA0cNQqKY8CTEpZP03CjhLIPdwl21e2yS2EE2MIsOEVWs4iBO
Ax1QYQpjdmesdXiXW495JOYygR1bN6+MpglGY27GKOvTRX5TOWo7/f5lOoaSLrHq
l92yxUvqyIREwRE62GxifVij/9ZWJBoHfmsEUkBgXhGuztqVGeXdbW9ZfrYPQX1K
MKZS/kyrsAbvvv9U5gJ1z8yURRNquMXHWSr9r1rAhIgpxYuWO5Cp1D0y/o8B83us
aMUsYvcPC1wNtQnlJIKvD54yurj+jWDkogqPPJP52EGrHmJ6MXOHXLe346EMJTQe
Tvq2ukHVTuDQVAtz3eERzPBhQNpo6ibjxIxnlihi2bdCkVpVKMOrHDzgICbWVmXl
ZDam8RmMx+8JlMdty1NWud9AinhfMKddZRu5UKABC0Cvn98REVYEnlEmaJLNtL2k
pih50gYkPGTzKEAqOEbkApHI6Dv/umhTRHz3/Ae4MSGmRNIj+ktjtPlwxJU7THb/
j/ssK2LLa0SEWWECJteQpOy7akKNBpA1kl8vL5Kr+cbmEkbLIPyFh1x683Op0wEG
RZ0dsrNP+TfrwavURjYvxotQh3EnTG/ytNBSksiBRIBKlQkd4fByLBZjSxjMDUZn
d8iZxdpEtWenbQEcWUiu0PBnp/OJ3MPK0IZ7ZVN+mt0IMJVTTEg19nofavjjBlT0
diGsul180896t1sUZTydK+y4fc9N5HZeuVHL0b2cHpkhYJbSc+4qIZvPOb9XQcgf
fvwQUgjO7N6uif3N0PTS9nKHNlOYpCVNGDEVx0Sx2eQsznSv+gFvcLGG62Cir9/F
t4sush6nocMqIZq/9Dr9gNlCTGXz5zgOAvEl6O6JnXsQR0MtHTai+iX7gP/CWg/M
AgMn8cVbMlei2P4g73g1s1wBpubRe0GbFkpa71NPxDP/xsOzWzvID4Fo0TTy/oKN
cfVXSMOAqBZtwWdIug2f2Sf3Dy+LCjwzy3br4LflCbKem98EFdQ7NRKYckkiTwrg
5UFStegsWSunWYAOO8afRdyQS73GT+jCkjv2i2JWCAOrSBP/BjCAEFid1V5X53tI
4ZPj1Hk46XSKMAXw3UTfn4RCzqCYDbkMJKD2YWJKgOkUaYuLf0lZfrmrfdcobLIm
e9KTV69qkGWA/6zJbzqfODOLihf+fDMDdcCx8KeoSJhvU0GRgLrA7iWI2PbGlolK
cbmzwr3YHr+9Y9jQ2CGgBjlWQD8qoUxtcgqEmRZDrnP+8zKCE4sBBuiApU46rp4g
8/5MWtO6O4E8MkPaDzs2ztFJXYjDpowRIY6z+Cu4pnXiL9pKf8tCLP8By+TqQM2K
hm2gRPuttXYcEi4SnuFWzyH8j5Rwqu7oRs/UDuaAKQSAjHWVDyDw3bmXQwLTLd6p
hafFIES7I4CC/DIFIooW+hOqWZTddzdP99s+vpy6syeXqNzD0QzzhvQuk6YxFiXL
FTjT6UHz8Z69BDjwa01AXcBSJGQlz/2gKD+ij/RSAk9a5gjIbDFyjTQpSGYopLtf
`protect END_PROTECTED
