`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORCLFpe3/vDdbTVRar6dFLcu+7LfF3BN4Qzqggoi7QsyUCq1S/EFd38AMYDl9TU9
KBNkwjue3kstuPkFMaZ1JD8F/DweL9/VFYBfwTBfWi3CQ8OBf/W4foYapr366HDz
gm9eO9TAG6pKrPN53H9PvcR5Tg9YGf2q8EzWeW6i8Pk3McLQ3sieBEI5/b5+SWtc
q+8QXokLYKlf1qJ9q4iseIWATtiQMeMqzjWy9BqDNFkLix9RmCPxa0iCEk1fH93K
SNVw6wLxJyVtPXfnuQbGijxYWPS++MP71voIA1oIFAtoNMvymTbKmdGRp+4h6kMW
msepBon+IUqq7rNFpNOgL1pqQqvGiwd7iP/WLYKuXLgh2qCfbAq8eSeIplgrhV3s
OehdUyflWPihF6hk7xdRhmNaw5Xzq4s0v3pKg2Ac27pwEw5pLHLkjsW3i5e41Q1j
pdCQL70RivbJXZfAgnyFtvHyBTY6wcnITM4Ucgrtht7ybacvzbM4f3VcRo4/m1Aa
hpHQNa4TefO53Y6tzHKUTz+gp4TYXIKee44yYD2aruMCeNPTHAHX/HHcYrHtni0R
zj6bsDAm9t/lmm0l4FfCjWey8E4/S9c0cHEhiu61bOJeD7mPiVcfx/brxXu9od4L
SvExg9rsUTTrwwuwr8NPMIghQRqejG3K+SVbL8ktuMBkXuFBTqAe2OhU/hc2jJnA
JgMShM6dtwxjklF8gi7aCQs9M4LScXpGRKPyDkCMbZ079H7sceVttiOXWt13UGvR
dY21EniKusFJc6wbOfY3BUbiO8j0WM8trZdQ3TYP7QTOYs4C7ZPbGsOJ2rS7gF4y
0oQS4JiG/3Te3lcm8fqdy96nQ2V0g17EBbw8HApdt/QoQy+w93S+UWzMfpDBOrxn
sZxNneC8rToOeuWFQhJ+iZfvf4DAw0Qk6qq61z4n0getBSl8JUUtT86+4XsAXmAd
PdBscL7nxI2d/rI0PcycnvPIEP9nAXUvHZ0gL0ARlWK4zRFOiGGRLrCDRXqhSwMr
6ceENh67ewLTpeP9t1ezEnqcQ2m6mWFl5yQ04xgXroFh0Awx4J/Tag2PbseCi975
F2tmW+KJBbhyVp0JjkuJm6r+6GHBUYi6j2PHwkSRzVScEtZPDW9i1JsKkWxf3tID
D9SLqLORADZkNYmCawJFAj0ZIPd43zcf6tH4x5vV4n38pNTmF715+LGID15BDDCj
U+O23mGQhTo2AGczmvDY9Fg5qWx/Q60V7PRs0HF6s51Vf4EWxLiuxPlydHQfJ6XS
YSs63+IcWkY5+N9eRtf7bw==
`protect END_PROTECTED
