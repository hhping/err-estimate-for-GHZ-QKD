`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Ppyl9XxKXc8my7O5yvRV8BRjx9ZCtONGmBB2ZnIlDEXmTAydmNjwzoWVK1TzdjW
RycnS3yh9BwRS4GRx+DP2fQZJE/9oUwNomuJVC4X1t/S+is74sLRxGl1PmeO9+Po
9MM2M3uti/anHAmJQxr0G71adeXSit0mVSpd224RJ5khxtTBpQYAwyUUg3mKqK3Y
Q/QTxaYlYNfaUgtHuyZ7k0ANjID5krYXW0BmoCCiRqvGBemN8xUyPHaoNP/QS3MY
9oM3h9j9ffrdq9dSQ3NmwETRt/xqCsyVbGMTb8mbQ2tAmV8bO8xKEb3nuAUdbtK3
2HruKpIt1QpblugJ2/+aeKQsKzvo0olJkhpHIfVk76Du9+IKH6gTnEDfErIDZzcZ
eAtVt6joTZbyId2e7db4W8DMMyft6u/XEweC/Ngko06Vu5cdie/DLiP+eOZKnDBG
IUfgJa68fZdeZ15RMJp6vA4q8c/PfnEN9n7W/Ms6OaQjdnBRZjkgNaE0Gg6J7231
mID4JRbH00q6iwlXfKMPbRoKbA4rb6PKzYEqydX+CC4vkYcPIPPLoV0A8mHGsXHc
t37wDcNB721cqTbqUmY4kTMOBPXm68JS+MyRvc2RkcFUM7Xc2eQihKOLI/haJwdy
kuCNmD0Vi1UKNslo2W7J8+i336FuTGzhNe21mxRf1zII/4fVHSAYLpFz5dhifthG
1xgW1+ypjuT/zAj05XWZcvFiN8umKIVjk0QFoTNMLPG0qo3guCUL0Zz1McOCEwO+
vgYLOMiraWo8kmcQWRSINkLeuj92wSWo4q4h/eR3n5pu9F/KFbvEJ5hOLLUcIWIu
uv4a90TuxDV8NqIOiuyQFrUB0noSsNF2pHj52rFnOlEvqgsYTBXsCZuzaBDCbpci
RG7MhvOnpiwNYFnddiiUo1hyXLpWUm/a7CtGVNC4oBdyGLmDv028zGs+IJ/SEw/X
XFRY5xbEDhKh/xGdh6FS+O6AIP9TZANr0DbAV+tuAdipgQ+07Q9trOUoT9K3FxC1
Jw83ArPYRYLbn/T79Ib4z0xZcfovG5zzeK+Sxan66kYYPUbzub808O9we1dfjGFH
/iWOd6gIkLYODxFyUDshz22LBbJwhTmLvNiJ057R4ZP+QaBCNRqIYMAkGxQ3u1F0
6yG7EqAJXMKaxCj6AaG8goC9JRkmUPblHtOITlKLmn5+X2uzPbF2IcSbOZy6CjZs
2ho3GRE768O3GPe+lHW35mf6OBumW+Ys2QeUB3Npfxu866UIL8L1pAwdUpX7fTbB
LzNyIEY7sRO/MVuC55U4jRhn3be6qUuvmm3wNbBqCKfPItW/SjzAvsJ1FsPAUKAU
YhHnFrbE94K4ABw4BqjEgQr1qD/tDI1FkKktg7lnBn4F4mgQ0uIAtatKHe9uJxsq
PBFT5kHu0U0cXSEsnjv4tVkd3iB7vNCwwVqTwTDqmF8pAVDTJqlQHO6je8mhVfef
vaIbIUy0bNXRS+AEBrSK2YBnJ0MWvCXl85EWrKgFtuE=
`protect END_PROTECTED
