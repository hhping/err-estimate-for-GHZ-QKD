`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsI2iEGrV/yHnkVllSKxUa0WQxEZLWijSur2SIIXaf/QsAQ/sCFvekeuVz0pThcM
6KTcWD2eE8+OUxC/+MaJPtcJne67XHM+H6hcjyLDGytikGpQXyQ6ly5KrEK/b+eo
XQXFof5ME9Qfg62MGvob/tsryIYcYaIZcdftVoLiuTCLOdhjys8J7cHI+NIsqNJS
/XR43xXb2BsH7BY2yN2Mhkcz6wnOQAHDFsxgPIMHPp4arpJX0B5XkxFiLJmo3QNX
OdY8gZUAbfuZGh9fnjGkujwTjiYAU+zJra1Fs+nc1NbeqZ0LdRgcmtNYRqtAddrF
dPfrEXRtkFx3PcBOs30ABum3Df6+H66b8ypoVkjxoE1Hkgbd7ix0rcCGj8JgSw43
dNSbEE24IbqDIysyFAeqmeJZKdSXNRLiyE5hTgnx1r9nhfKTWd9G+TnrkAZQkGiL
7QIha8WAWEH0EV7jIjRaWBmIrKuiFftE0wQcqS5Of4Av+HUuoJUAoghOwvRhfsrV
Aij/ETlH6cM10f15GdroyShWQ8lNcK7KbgiyjnNKRzu9PqD626JCx3y5LuFkRjPy
77M8uCXn9WbySmxWPy1LWqt/hYjMiQvv76CtDtgv4Q9+m8sLKSsCvOcaYj6+szDA
QcigCEnXAqQIDIzB1b2+ptpY5qVqKbGRVcRByAurT+gct2HWBAciKMcuzLchQlW7
B+47x5ZpQnQ2QHFxlDuTAdmbDffeQPEsEHlCMumLTni6r+xAMqQBA7DzPbYKkhp8
yNkzGcWmReVWywfRJOQ9mHsA8PrE0w28MjNzcOXgeSYpD8SIbszL/ZeDXHER8H17
OrTMrdA/6TZ669yZL2i9kfyNUpXby+qNrRpmAghC0peji8JN+oX4L3ovch5bWQO+
NQi5NpErfB4m9G+RCQA/84gfPR/ZpFW8zYyXRK3CNTgK1C67HHh/sTLb/rZkyXL9
WJ5xvWOP6niHDJXcYZo+MibbdQ7lsIuI0T6lh3gZ575wQgCiq8PpAT4gBj86V/GM
sefQ38m6uxJqBtcgnWlN4h/Ga5tkIVO2nfZynMgSyZsx2MJv/WYgIJpY3kTZQwhi
50B1bR5p2ydaAQG04Qc2ixuctBlRjFylaUBjEaJqG7wRoQxQFHvFT3qd1FUbYGZs
IjJ+1dJf33V5tusUq5cZrNTL3NDeYtYyF5Qpe3ZaBNkXLXSOxxJuP+fCdRho+4zV
SOi2fZNET7ZQ7PmN97yFRLXcILeD70UcSU487vl0n8dsKEfr/jFBDyhmSStRFeSL
1dhQYPiiW3lxnIsTPK0ucHJxa7VHgAS6Xg/62ttB+V5Mm2kqgdN3yHnZ9lics32p
GhsZdONU5zZgffh4p3hhPKr6uy/RefNyCFX/7P8ZyAO3DBdtPrHB9nzNwHvveSKn
7aHiX6tqO0RRqI2Kvw/WbAnukvgDY9LOKb/UqAlsFcjoD3kNiCQE5Gbb0vYE0YUI
vTnn0tCVD7zB1wUa8PFXrqp4Qb91glRntspwj0Tf6CSeZLgSnS/iOXtxzcI6CEAb
1lm/re+YSBHOJ2xme5gTNt1JPLMuyhty/7KNWcddJyuWSkraig/VkVB0FlT2gOtU
3qvTMt9WixSyCwu6k0lRBu07l7TRDasdLSvalOw9czy82eHP28LJMSODdIOoPZ2K
QcxLzZRZvpcZWsKvFTfTvTvkHUjKaFmqAvPfFx0NxzCA73eMxIh9+uIiigQjmLNg
DkmE2768CbPgjGItQFxbF3ewaA34ZdgbVBnOEONpYwAjiLodurZ0t5kF6t2rEFGw
n98L8Bshb64c5gp/t7sCghibYN1xTjYWY6vfAOXCoinanxRjNapvaEJ8jil8Iwyv
hLzn37urg4FtSmMFwL2Ho4sC2NidLXbdHx4VdJTF4gfDwQ8VW1T6FMft0Q6vi80w
JKYXDOoqFVRvgIMhgTXp22Akmdx/fvdiyYaG1ziqfhDxPN+r7Vj804wPi3B5eqbD
qcxT8ABB5170FLUQzDJsqvyLStWXEgxTfOeGARxRKMIptll5nc75p1KJOmWWrc3m
3uqQS01LJE/deMyvgEpMGenfGdxxWRimhLoylZlZQPRi4I54bBPkxC4noHNuoMOn
2lQV8tHeZqo7AddFBIuGeTT/zcTP/ijMrZ03knFLtsFHL+25OG6XWMy7Fb4/qVJS
J58D0Udea9G95i7BVUyUQ0p1F9GkoDxgqqu9icnT6LT5tlr2+kLw1eiwbn7qJuIr
C+jWc4OXu3m2eUpf65VQMMqVn3ZLNcgbAsx4pZ2fPoUgVvFvP2VrzWFNsuspHDal
MYwFi16kMFfT+BuL1RMcEfAr4UZOM+zDCFkBBgGTIx0cK8GUQcK1676YoyyrKCDS
McWL1fMTpwPvjkE5PvmRS7N8PSzO2G/FS2iwEL+lrz46BVyWiwr01Re8WsyBowOA
mXHbW1zx3JmstEDsLMvtZMDTo+6om+10hSRsGjpKN30Ez1rOI1ObNpx05tyxBWeh
thDBRsaukQAJ5xE0L44l0aAzdTyqzKrhAXA2ajybUMEPZnx7vEg12zAvrs4thtd2
K6RcuLn0fVKBf2jPvXZxxAr8dm0RbCFlwmO2YM+xsC0lmXXdLCXi9A9LeBuSKV+b
0URAiq1m8zLo9x6xlE8GML8QcO4PugS92/nMrCJaJCxAq0BL4eF0OMo0Kpneidg2
i+wm/PUBx0sbUc5kkkoQGKo1e72ZctvWH16uQ0Ae3oJmbrSwIBYsgiG+LOiuW9NQ
UD1QEhyVJbyhyZXLyuKZW10U1fPy1IgLJ8Hqc1tLQXIi4OdSCmLSs5xYG2VpSgcR
Vx6OslEuXvc5QfvZT5Q0dRsgswnhGBm+aub2Wny9z1aS917oY3O4ltnDWkjnsHKB
9CW+PzKN8tuOvYe/ZFiAf+4geVQmO6bsfi2jK6PiHJyRL4m4QmfolGchS6kZOYUW
tJCr2vVo5n35cOoCuDEXqDHAmr4Rdp2BkRMyYXN9R8SJYU6f9F3UJR22WKtnDUyq
wY4j8aKSt7UM+Gy8h5dRETR0bc1a+pKtvWPR4yZQKA+qrfVT8Aj+str2Xj6gLQ8j
PTYO/yBQ/OgcY2DMARdHzsar31ojApdSgx1APpxGUblqRtTUVzKBTA0rykhpA8Ge
RQhfWkSOf5Qd5ZfQv72LX0IPxKwLPmLvv1EKGjOSWzGEKHHVPQUK/R168OMy8yAD
1+HmOmUYtOxqgrkHLIZXqQ1QANBATtHVYoXyHqZwtvlyn3xKZD+vby6yCpdg+zso
jmK5YvxKeEFtOloB//FXYYFt8nrMLAo/HJvl+9n2yWIqajBHy5S9oYXLJGKW++pt
Kyd7GYvf/8OqB8nNTvqynZIh5woIb26eLYIostnWio4DD+Akl87/XmS71DkoDp5B
01caT9h/nLYaRZ1QALgj8bfuATajeMa62KTgRKBI0KidXn6VJDSuecqDMR2ixaQi
`protect END_PROTECTED
