`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRGRo5xEi5LtvjgnYGGbw+1fve/1rRxSDERm0cf+Bd9UHXtDhKxsHG8QweWcJ4J6
f5LAi1QCU7CC6vlDViNBkp+NgppTv0Sqk5etHvkrKEANBtJH8BN302XhBqAzUn/W
5Rlx/hrA68ZXuJBdd8NZiLr56NyueIMSxY3GPKOJVdhvCjYCw7bSq8RHGv4b7Zz7
Hdb1mM5KyL411Y6me96NIzpdEwd2aTyIfMrgREf2VcE/o6Dq2M6xobxNah2d5f5F
jmOozwHCvgjn/z2niZEXxVJ7m6NIgQqizZK/xXUFEmtruZh3Zayx9FnKSKCp3frb
Z8KIWJIHnigjPfD47kL3QDWNwy/dbhassg0S/5PXNWmAMOlD4f87iDgygDhoEJee
oeJI/y8AFyWurG75unxHpc1pmb89BAIHvYfvRltwX+SNeTz1atrbZdUB0/Tc4OjW
pEZ2WpLttteuLO3NNX3W2gtt4uPmVN6fklco+5WHaC04ZabaeLubvP8Tx6JMsCqq
R0pwCqBtWLahVGA9TilqvJr4Czf7Fdvrj6JWtpmvmT508a4R6ricsO9kD9RAISL5
xN2PxYWdB/UIz5ZYqAhYDqXQYB8zboZyK5lYs0DzxeMOaRfGnqCrUYHysQZFwwxh
`protect END_PROTECTED
