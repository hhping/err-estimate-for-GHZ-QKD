`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KejOOqkhgkxMisjJjNVl72DMoUcbcZLUgaeD3TATVfRYS9bwUhbw/xtE0q8rVIOz
9hDbc60/spzdgR++T63aKzyfM6/HKKH5O6lbRjrZx6ROzFW6RzmFenH3im4LkibH
cZwjLua30apq8jJzATQaehRfBo+eGnHZdkQR8N1xgno/4VZPXF1VE8WaxPBpXwqk
ojwV00egt1Ne9YWRrunz0tkFUFYdI+ln/gemiaxt21OX0aryu10atcOHZs1kBkv3
d7q5zMH2oaaZ8Eik4nGy68mYtN5d9nr/orLh5Jl5eUKaS5NbOvJipfbY9LiRTOUv
VnoVSQYZl3qR6kTVJprvkg4/P6m5s84DReDwLKzX0VUYdvAHTYXstWGPRMNKTyB2
ktPnO09fT1l9/egME9meIkYQa7OljRWeD5gpn2NDD+5kQ2ci5Csrya/hSK9yGuq6
zoGXjRVHoXXZzlnohHMX8Ezbpph7cxC11B2PVvSAVE5f/781uiMiYkpmTWZHzO8v
un5y8r/EWqmzMX7GsIUEmRUKrBHVoksp7/FYwOYsmScLqqFBQHlZvNCCSNrNFsZk
TeQ5go5Ht6T22gnOxrFI/SM+0DzUPnrD0cfscy+uDJqbQqq0teZhKbs1s3F0sd+8
RO9HKzpx5QB2/vLHRIMGsoT1/FZfqaWormK86U5hZyE23hznen6rKVcbJMKQMNBD
WFzFcEvmUeKJEKthzyiHA5a6yNbMeamYWnsTUm687b+zw4okmyOYrCkvcAZTeYVe
JW2KY8mgKFzBLMH1Os9ONi46swASE/dQwsvjWGyr5/w=
`protect END_PROTECTED
