`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsr6qMnT4bpu2ASGWgz9J0jxIbBfaQHVzj658Ykc7KJ6R8gN73CEfFu6sP2sz7Z6
b6bm1G9rcSi7sSUGbYozKyQrM6feGTdX8e4bujzgZxRmVzufUkCSJwgYXIYx9HNt
C3TCsrBC5drkIbXDMIDj0fD39Kb+eBiMUtDtj3GeK8ifwJ6MyoEdFBKXYNyF5xSs
AgNuVYJRaT191ZVcimD1TjNRy3ci9b3aLCDrZbIqjMxVGO6BDxO0IYx5DNTsepYB
ezELM25ic7Ju5Jzu516UP1hLVdcPFM62jkVvuzPzu3FUvy8B5fQ7x2oR6O70Zu0Z
h1aBd/EjwfkiJCqopMcmVqbkeOwIDcXr3flP27qDkuO2JZ3exGSym98PZ8irbq7J
gaOb//Ot2uqXo1a4SYpc3s/6yRfU0/9lsW/5Oughaod6c/p2518x8qhSp12kIB17
lkXioG5hofNsmjJesyUk+gxD5xip+6l77hr8VBtxCp0uaHBYYTPSrP6QwrrD4i/H
5wOHhKqGHpCQxqqI7Olby07L8mUnA9+U+1e0qxJZX7wkAgvhMzBVttY0Pietpxh8
Ri0W5juUtbkPITpsSTE5cNOavyGHy4RBDMTFl6cgCi21ycK5oEMOOOXPlLixNWK+
DITTFHbqivlX0aEcnyL5ZfkSC+0T8BvDJRAKcSjh/e7D75oc3S9LeBDKo/69vEuI
e/mLhTmpe5gbgGNXglZVV7/RMuadMisJK+GIhuEnmdp5o7jiI+E4+mHrJyLcqM0H
mLzhPi6iiWF2GELEFzlEMmlgEXaeppqBFGAYxv17eqDQVxDZLcaB0cA5Y7UlHQ5x
hl0uC05eFVMqnsqgUxIj3vbi9jZgx4cRCjbShtKkcvvKdyewFkY5oUKgB8lNTRji
87GqbOvliebyBfeNJAmfZxTpG7ai6hsqFQ9jBGo6HKFUyJmEg5hrrBIEqRyDrE2s
H3yCzLAAU299nWiQ87PW5KKfaWb4NzUODNdIjynHtK0KEshDRLdMxNwq9EuxGmpc
vkUFBeDQEMiGYP0lqIOBYJcY16r6HPa5OvkunQ3dbV4ua8qN0tkJ2hahWJ8xgglR
D9OgEXFE56hK32M5Erel9Z/Bf/nHl2dOZ2jZz2JQXVgwRNsRkT8PjIrpsEzzobpr
ToHfMi0GuKHkaoZX7OLcZuSg0h4Li1EM8rMw0EJcJ/SSgFm2rKETx4jO6GVaAxkG
2etaUG26bakurIVxz8mew/VgHS+Aj6sB8c1AhVs5FehM4dF8XfuWlN85Scx7nGzs
ltQ2OGQW0MQOtaf4DSNkpu8BUBWIj/W7PeubJolLf7BMPl33vpI1yzgQgTc7WHl3
K9teb1wILlI58xWvSzxMsH80oOgXvyx/3SO+McKd+edTDdfubIPJpZnF43zR7B57
VOxoBZ0AwSKgRAW4gQ9XERp6ml3NhEoIgSDuy0tb4rjn0ZSgjR8iFUjAo7lL95tI
9BdRIiLotlGzt8LGw10iiH5tTyvR61ZUkhkSCLiKz4+V2IV9sjGf4nvrfmn1Im/6
6YF7P/yc6+2TJ2xgc+b0Ofus+ush+S4mMuoOmP7Mvtp9tk55Emi4sv+oVtCAen8x
NG/hhQJsNUeP+qym06FqVV+zgaLovt6YSZ8cl3N10HXX5tTb4xb6Rk34/w+T3WWQ
9wtUtQd251moVP5/YWrMd/bKpwtkQQO3lbqYOP8PsvVcD5XaDuJpczAUoQX8DsSw
bcqgaKP9zGgBbXljX/iglozokNRDhCKdbLCFYTpFlHN79WtKfuJL8i22uXewMCv/
wP2knQHrlTQLd/PxSHCtShRNXygu6RvAcrLcwe5s4i8kidh74pxXNNohfkrUJAJu
QjGrqDzigHl8npaZtVfIWGg5SMqVjFnGN6MVsUr1dj+q1Svio7Es/qViaB9O97vp
0FrB0PTODROCD70IdG5yFk4JkNg8wgAfaRtK83vERpuhYDyecjnlzNez9cSMONpq
c5iatnBT+1ktK6IOeglmPuxGztIZlmPblfipaeDtRihhkK5tBsPLcJv0SR5YXRcV
syzTyu7W2HKBnDuxeO1RQgbupHHAgEJKK3J/AW/uPwBl42fyfUDjCa0KSR3kTePK
KNGL7QmktvmynwOw8qBY439V1ISbO+/FgP8k83+sZwFeGWcuwE11h66ZDW/8SF6D
bdMAVcyGzSZprWsmunVZCehbX6S9IvIFOt0K2iirGajYCEOgj6SSWAiq0u+R9+qD
ZhUyGrlM8sFUthB4rJSQ8g==
`protect END_PROTECTED
