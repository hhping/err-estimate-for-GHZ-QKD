`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXMwIJenfokx88+9YF40PzMc/NbKgIuh9BCxmAWDCTVg1XPJVHuZ4rwNUuYSWemM
1XnQThqgfV5c9ilYY3tVDpGE/API0R8s7xrgpbRmsNnn3ZOIc++uDsZ2T13HKO92
Nok+LHXWKDK8ji6LPLAsktNhpqhkV3IRWPI02bAlRjzJ5uTxIALHKnzxklpzQSBE
vYQfLvkiq8evpPLwwBT9S2GjGkAyFSMD9gJlB3tLgYDVH92Le4b3ilv+gh38ppB0
TW0+fSunG7Dau8E86Lhd+Bz+qm1h+h4HGBNgyqeUtj6CRN3v94EhTooQ0XtTPUxG
1D3n3SNQTNCKShYCXQ+nFeI9BqjjgtwZRoqzmcuVWXbcLGrwrXFgCY8fGOGakuaJ
Icz9jizh5CmwInLrDpwBhDetbV+vRjVSr5c5iysWR1GdtWO/NG25jImFXLqxh+Iw
TdyP06b9rEBCEjK/4hDrKdxQUStuPV+jSZ0XnYbpVL/m2JSvoWxjSCepXANm3SBA
/mIZ4BT3SvivnKJQ4E4BVqc/cXFrkTaTW/zdfySOYuxSNDgxUgOhMJesGE0ei0mZ
f53uNp4z/cYnqWve7IrDhVhbfvzVokJ/WJ9IkK8MnOLITQOgFLCEWFCNBXyiPL+0
T0GZRpAbzy4RHq4jjetYu7afPGJq657zX+PjIwCyNO7NaKesyAcl5KVgvNUo9fQ1
jVlQlclZS/Z66HDaL5MKirkEABFkHbDZrKdxdYINh6Ugedbx/zJcuA32o36FsLM2
JjhPVH8soE3A+iaNQUjLavhqfa7LYxbAeNJMBnqzygTVOT/wJ0RY4DNhraSGq3HZ
YhFtI3ZVpHbNw0V4VIAiA4QZlErODE4J/teY2JiUk5OhnjBIExtLJByxKuW2c6jF
49enleQcIcI3KI+ZAOKqoNXE39EzdpgAPfVvPn/54e5rnZzWGsoWpGhOdJvXvPCx
CiKccAnYgas2HoXDmadQFZ4hdoCibjlNCSzjgEmv5jWcDGq1Gr7rsijOMojLvjcZ
dNRkntop90Oz+m+xesb9ysNaHfO5AnOydx2O6cJpDIbW25+ezl7/X9k+mtCFr6eC
ZO5R4+5Wq2zo2HNjtowjZkID8bRDhvuyLmPWkEGehEM=
`protect END_PROTECTED
