`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGs9bdTtBYT5iNrLT1WWnYGhPvLys2MyjcrySSi537ELgtzP1a3y5YiEHmhaPflb
1uZboDx10JDT9bDTflKP9bxdoOTIlxjAkwHiVM7edBk8VxX7IPtkYv0DJ1TYQT9I
hhrYRoAz8t0t9gV7zaolDnaBtVRZ93kgqpIHjJOi0DmFbGrfoHnIgNX5n5EfCLkv
dfFPs73PdV6yhLNbO8uhwCKvsCFeiZK/bjKQHNcqEFPbL9k8gKb7TM1sb5UmCt/u
mPdw1g1ctGTh7n+oPu7jb1gsLNzUOInrk9yUecJwYuJvX8572hpX21QqUQP4Y8AW
o8tvE/pPIhOllTj3FyT3HVXTxU2p79Av5H0m27ouFDsHMVL8oKBMvQo+CeaS2VQK
uQu+8NT5oQqqnwb04XLqNR3VTul1gvVQ03NQ094Lu5lhGJFOLypSHyHgKEsvI6BF
Vzbw2FDT6xeg11nlaiSDpeltd1xUdasG38uuhFMUd+ur+ik2KS1mwiB3jO7BZC1p
Nrs9mm2ix/vdKTPwN/5/ZK35IGSpP4VkoexTeTSdMiF27NFiqvKuPOzYF97xdoY4
uWwoTKJC7PX/mZvTK3hPgjHx5MMO9CODbe3/p6sfmbLx2LUVkKzqb+A63Grf8X7A
tPdt7m7gSsuQmuJikbz40C1lFbopumwDLk213wT3yBfTLEwhjtGI+qts9+7pn6Pd
QUi6iJNemaZ5aZ+MD+DUbsKAZxGtP5HLHD5WRjgMosDnhEq9bXm+kr9tSHoA2e+m
VnwBLkjEXWT1wlVQmvAZBKdBsxo2bPTewYAObQTpWQJn43pe0qtFVg4E3gW3mMc7
517rVmVoQNhM0m9MTyuyLBdQ63hI4jYg2L7mySqFhgaC4u//jBkUFeKF31Ezxtnd
BJkgnOVnqQGievMQwWmMqLcF0NSn1C4TUc3Gz56Cyc58khvzx5mbxUaz5scEypgG
zguetW4RaumzAprbhTO+pdTQpLwb3FuvhiBbfwpNizWJHYCo45msSxUMtIEvrGaY
ygOp+pznpGj02wqxTReSPj2gV5vh27DFSscuaNuqSZNQ1mGLeKI5iSY1nor3R5AC
BvuMSd7BBBrmYiu21JbmHCj9TtS2yHbV8zP9ZwkPteYkAkBYRzl58eN02O4gRgAn
BtcK60XMQvdIPdaZtauvuIhcBKRNYcPb389P48wGXf29RBCy9qRVNh12mE0yVt2O
BhMix0pbzZfcCUCypgbYeATz1CmfNxLflbi21ZIfmeK9N6cCvCRhD1EZktG0sGZm
VbSIekciGANS0OW73kIR/wVvtlsSZnoDKW4vEJujYAakqAw4hWzNOcKbWELBSHEj
cV/5I06sYVl7KWfhFPLnR+zmlEv147m6Ow9POwXGEOYnf7cf0DMb3F7ryhufXvTv
GNbsbZwK6BXoU/5L85QcDjPhYunkLwTMioBeKAsw9wtJoxWRjGUHW9gT9diO47YP
ekem6o8uwTAUS/0uUG1qR5znL3arS4PN1iQkp8er1AmdZ3g7abA+bE83iAl4TZCw
49wyPHxrVXITSMY1QuS8g8fbhG000J7JIDi335ytQB88+NIrhKv78hLE9xE+xHg1
dMa7z4QXkcVs1eAc0duS2W9eshYP8aIcUPScmj23d2Rtegex85hTw37BQscfhMSu
Yt3SAooNPmwK5B0RYJYSTF8SVo3moqaA8698vdiLktbG52SqAQxXJaPO0t9hEX5n
8nTYBnY3GaLyVb54II/P9IOC3xYs7pdh5UZvGL/6FtRpRvw/tf/8HhnK2Rysv04W
rBoP5Jbag38Jvbdy5rlRtMtsB4dCekfzxDipEpnqpjO2GvL5a2QYCwzG+s5fFC1x
RErH/jnLwr370jHbq4NO3vYdN86HDHCv8FntXQWZE4ZAHQeWyvWtJZ/LYvO/11oR
RHKWw0pTnIFCHL+dcU6IQiNt8/0wTtxrzCzihYSHIYcaA9k7IFn0+8gI16I1bNhu
xwfhDcdJNcdwOBSAGkHZAx8lExvYh/a/SxW42wY775ZrpzgWaBOlzTlJmW13xTfh
KQEr0itx12CbHZUCfYCLtp4TgZ892mAxZbtCxx0cT9qBHWEUaW+9+oHeI7S/ZPAv
SM1RrKQ3T0dCudP08/KrgHQGgqQVBsHmGp8IqaYd/19ulhdEdyppomis41PAEkYu
`protect END_PROTECTED
