`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RRg+bznJmnoBJ/B0BMTjL1EXiRez13LZgzg74EVi9kfVPYSBGEsNwLmdVnBrd9FX
FK0EiMCncHZZjK6dtQP5vZIizdVQyyxbytdvk25HyHQaUy9BU1SLIplV/5ylJw/E
CU9HQP/qvhNDJNpVI0Wt+/QPSRKObUObAJPRuJbWLUFFqa0RZ2nD/NtZA/Y0Ai1i
Pb756IBSVaKk6iyKvt6/Ajdfoo77s3OwNuxtF//TSC5XQDz6//mi7Qe0xoLpLrau
4Xw9zfhhLSzfq9U39Or44rbtFn6s1ogArUhn7U5RrXxqaBK3g3NSWlK9V8zyevQI
XAlOyelOGtyu9E/l50FXN9fWP4gtuv05XEj4bHLB4QBduRVzcXBRldyeK6X1czJU
DT7l2P5qf6c7yi9fytUgndVl+XjB+L/9KYUyixzUnXnag8MTdwKXiRQqXgbxYb1S
Q4P20zAuq6PczLWjgrLpqHSPFvkKL7CeKdLhMz7tbeQh09a+mN17N7Za4D7b9VH9
9vUc2kzFnAqzLykJOyFfr2SvqB/3uAA+rRqIgJT7mNSS6EJ76+zutS0oNUdEJ04I
tIdq1m2q95Ps3rrHN4x6492B9ehGd3QfdsCUrBjItcJnexwl+2m5xUBDryeuynyu
W3KYyNyb8mHmiOwQUEOQCUD9H4TJ+QogodH5tq9uDGM=
`protect END_PROTECTED
