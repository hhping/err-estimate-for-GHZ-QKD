`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWeMVA54GTEMSR4dhEfDXUyCI5tqS4En/Z1YN6gCOERpOCvczDofl7YDOzPI8rth
bVRBsSUbumUeUJpTXE0024KaXSohxGNTQo0RgS5zq+wW4M5U1Lm9N8aTsa/fGH3K
Cak0gX04KenKbEMphDK65ad2kdiS2hrNKjuHpgUrrLnCSyyObxj4iVjENjrbMy6F
VrR4Yp8HEHDad6ADoJYkY3c0JkaIvMrusLu0RtEgmGRplDB3XHVgi+xBDm3cAzOZ
SPLHTjNGnkE6/XXTF4t328kwbYeJe+jMIUIemOVxXL+4E90vyE602KWI9pRycT+Y
oBBaR7TOtjEOdVJT/Tqej9xct87NBr6LJMjPoRNmrhVRW89JckEEClsoHaDD2TP6
FAc4Y2G7NTusEwV+DauEkT+Sw5LHmtcPjAapgQxatLyfSbWxdkuNRNZTLfXSQUsn
T3TDynpi+rif0zT/d81AJnF+FF5MMSunrm5MdjTNTd7eYtq4o2KBgm3Ki+/PgJXp
WMdTWDti0w8HK71/py7WxydITXuVIGpL6YXidBme1IXiAzpDcKbgQWl5+r3Oj7g1
NeeTDHzBAAGhgKgq5IIkWSSdfz1nVCBbfXxx8WRsBOtR9KAnqqX5FgB3p9FuL33w
`protect END_PROTECTED
