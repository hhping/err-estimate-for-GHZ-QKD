`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i8QysuQ4Iii8lEC5OsmyJ9HPH+ZWYN2H+HgprzLC4U7iELb2uSPznCgV0Xzhl5Jb
AMaDFoj5hVOiKz2xpdzvdtKng9RWPb/vIazxIH1lV25+UxiXBsFXa1xvdXl3Am+k
AjCLB7HHuTfJlq73d0MfUrqHerhIfD2Ih981pcZMovXCtE1nORx7yw0gnN5iAgR9
GXxO3k0vxb1QACeKPUAtqfTQQZRduMUhDcbTsxCB8rlbPApg+21/0mze/RPrCUmJ
A06MFbh1aJOfxxLuKt+Dsk7e+jCSS3BzJNuojJXqMIfJuB6431kUI81SVqhXYGUk
KMQpfNR0EQysJnHelFZunrau2uIxOOe5gnmvRnEfvxDlwU+jSQqQaHBoxQh71BSk
8e6QQWQO5m2OcS4mKJSO07s5rwGQWg5HN5p+7kMS7IVATzoygrgr1jwOgmSN9mU3
V030SuXYB/aXenAZOPzLFc0y/lIdHuQTP94LTaoXZr2khp8luJSh0AJSwswdSctQ
gR6AJeOFX1rTxrRmuhzARqO8BHPDaMsO8QtuDBMnK2fxGwkk7zpvRV+W0R582dW4
wDZ9W6XkCiygjbXTjUwRYcpz5Mtuqn7uMB+VjeSVdEbtsMgM+fceKknTofEG+QVl
iu7tyXMWG6kUP1gkJg+YKUkwwBzATrnJNgdFuV4LTkfqOtOnNS+twe4GwLuLz6/S
L7vWIplRu4SqtXs/9ivlMlQXLBuIo+bmGykAxNsenvESBDIzznFLwwJRSEFDzDag
UI0VifZn/gkBuJko6WIcXQW1iV9lqhkTGKs0JABKZ6v4jEGihkOprR0ibJA+TYUd
n2l3sIQUz5sLRmdRrm2e1dmhyb9FE7g+In5qSbrvMfjhFrRW7geShqJrsuNdul+a
S9plNqH6XiL1uGg7rSyuoJV0EcZYS81Yo9W2B4FcKeP5uYz6csi8TIoQVYZ13BOC
ZE6p2z1NdisLagocov92oilTkaiZPtR87H8+MoKJqXREfYA8v0lPaSVVRobb9FtA
JOGulRwK4C6wPTnkVtrYoWoLLivfiFfV0mE7ddCpUSyqLnZtLJoFcZA2/pO9ilRl
bcqD/TRNcoBpOBzkJiAZcAk5Gza15KeVzKKAWiciAnJjQaXYVwBxk0SfYs8DZFRW
agM+vZmvx5pQ74dWpPn5rOZSb5Up6F0ZVQ1JdXj60y0oV/f82oG4eMOgvE+1APwl
PnS6074KxJCL7qynIgGFTXPQ6AGoUkU4iYnY73CW5nxpi1eCZ4P02ZaIkKQNIpoj
iEk7ZOUQ7GHAPPuIEuzRUHkYo7cjBXfkjPhvanPk90QuK1C37zK990WpMiFosn/x
DQ/9c9GCfwzBoT9mqp7rbkknfrAxCywfI28IXVlYQKGQDkbqQkQX4BQnhGqJfXlX
4FNX9qnlOt7tMbVT5Ga9eAVi2xIOwVIvG8mUmMU2HTjoUiQ15bQ1CFr0cLJeOG38
31AdjuRMVGJwyyTdrYD6o4ss8X/rutMruZoz9cLSRp8v09cvdn+bwU7nsiU35MsJ
57JMSU7EzaHC4FKRoybM4Gj2OQS2JV7fGIz+mEqdgdNaNPUl08jUZgefMRKAsfOg
OhwhkbF1ehZI6LsZTJAECv/qFwCTcT5AhUb4g+7N3v7qDEtR9ub+LSs9XrezmDGD
IwHyeDvjIPEUq0Qi7/vw6Ivo2dDkMdSHKiKjW4d26i+VBTMrM5GhhGkSGwECPOR8
yxHfd1DYYzJruSkMQw4wcI/UVnZWi7ZPP11yme7+XHxfI43hFiuvMV/Lh2BQrDPZ
bM9MO8qT6lQW0k0UXPJ/rY/P9B1wy9H558AOZjLVYp3EtWnOB0XDcsCd+457zMhh
9TnqYQQn3jyQfFKtm6inGZ/KENct0ldpQxXLq7XwGiE/9KCPbKABnt6ae1s4eZKu
YFOb9FCjMIfv7sXJpRbYNg9XgUlLPog33yVZhGfXA4jFF5HH4yU2kogWnZmmIy6K
9c188g38HIDGHDNeU4Ocg7L0vdTp9d/7G8AgLEU01wRjqOzlB/QLH8EWpgGrDJhF
fDQrRHeqamDyQwWN0WVKR6WANcr5GCnYS2EP0d8DYH6LGVGv0h5UV7tB0vQ5FHrb
miAfKCxP4qONyzR5ucI2AFza4zSlFCk9JV99tcxKC3qInVoKyfrrUQtOG8+3MaJg
6bT+XgIt5R7LbxoFNxEKxTKTQuBFbIjTC3s+zJdJeeRJyliooM1Y07MubFwmGJHq
uJmTfHwWlQNH/UAxgrSWwNzN89rsyB9X4OFaEMBTsnEcTgocrs2ucuobeOpNVNcR
l9BOu85jj/DakI1wGkA1CLxty0qCmFu24u+5hPR8pXw7VXXbQb/iur5Zf7itepqK
`protect END_PROTECTED
