`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CrCoCvmbK/6fBIRzW1b7fWb+Lim9igIqbu5hw9FNwNYysHyztMAIY/0ETXmjQ+Rt
x/3lUsBurv6XnT7zSIRw8dU8VZbdaKq/jbk0IXlwqt9LJ4yFcXYeRniCjc7Pcsvp
Vgw5v6IpyynQCaE81DpJJnsBL9b7ivGXQjzN4e2uB0s2O0PrKPgrEE4XwQB/bg8g
9fZ3bJfwiBaxZjqQ6iS+38lh4Yb5+yiBExnSXm19myTc7LxmpteYZyCsIEQc9qkY
e+2mYEW8LuOq55mQ/41n1cOHP7q2uO+yVoIau89t544zyswtalnN3R76yLjR/lZQ
nXRvI4TC5xWJrHNSMuqskGxNqzbIZDFE588s1YhnPMtPM5czvE0aACERHJLFl8oW
`protect END_PROTECTED
