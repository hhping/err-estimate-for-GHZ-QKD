`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iOoJrUe/9FqE9QGz8BDJhWpJRol0BAOIB1RYaaNCQWg/F/ncdSsosf2BGNr59vnn
W5W7Cj1wDCUH4zA1c0nD+pNWsu8rIRH2+NVw2aMyAknCljOxSb6B//XcOHoTbtC+
LMRXA7swC6TM1Z9LR2L+45hptsAJx5ihiO1NKr/dTuAnNTUVXz1/sgV1BQoGgM/S
7KKTlYBF2X13qCaZvXyDQ+RvbtSGVoLZHKVHio1lhQotcynYDWSJGKeGX2NpAM7e
3lgPskDXZUfYd85xMxw8VIWfE0jdLyCbN7SoaLBy47gF7bw8IgBylHBwsDM/LTcU
0ScYhRpY/+dapV6NN63VTv9cGtS44gCfAItSqKuPn4zV+Bc2ZjTsbw1VK0J4wve/
nFnUZ9K6Yx1q7D64kWKqoWsrADvCkY+KHKXcPp2qnMQzPvE6RZJYhJI2R5VF6Idl
bVMoUTrHTEIA+p2Y2PDL5551Z/lyvzb9mKfxLQOMICiLAN5y94vvU6xy1TYd9YhU
f8H1zHguaT4o2e/RPUUwv+EcyULYJvVUXSzsedp/SkCTjyojAdYTSDfe+cF8N2KD
mmw6f9CeQIhL66m8LWKo9RjyX7Coke886VJZzoJE1jRcJbVCZVe3p/pkfH5w1Fji
OvptxOABum7NnSkIme8C4DyguAVymau8EZtrNVhF/gjdc/lk4gGg69HaNBRFwOXt
49B6O7O+bKD+2bGLj6DzB02B758MI0VvDJpm2ZYFom/bRLI6OBCGDkX7dvTuxMCd
/dlFzQjeY9+VEfnFygGAstt22bqT6hKKZce8Du1HMDLB2VxthYDXgbsu+Jk/jFoS
S3P3adM29zjHToUPR74KoDbfCgMivsK9Kha9xLv5mH8fRjeA0IwvVo46ZnYPME8j
rXUah0ungGJae4AItGl84DZbhd+qDqgeuHB8aEtrk6NK/vu25kML9CziV7blPTiw
YDTLstOOylLM+XiPQthejUKhMaD3c4EFsJGfgWBMuS8h42EaoUHteQhFCbbfDxkk
5UNMs6VgzGeBX7t0S5AIcV4Q+0JUbikr4hs7sKnFGWd/b/dO1m2eSRlHjIQo6KC1
y39fcI0IPTyaUc3AZh0rNhSjBVfSg5LSiFSh3L+p4KifxC4ER7INFRlFbqa/mgSC
JJWYWX4TE07bXOf6tkx2kO0H/41MV62FTKD9WCN96XENF1o1WUlLdcJyovLc6pCc
nHtx/Q9m0UkdDAp9phvFZ9QeRGdIeMnmZJ4GYXEs8kB1sZW1cOEHIP730SBS66B7
sxfkc/DncwDO3ufC2QJydEFLNeJ/+r4wRrSdQ6uHtFN5GUZyiX9Fd143e/6MPiQH
A4Q7z7ij6Fje330L1ITp6Q==
`protect END_PROTECTED
