`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDOZ2DTGvI3VVDd+9Qyj00vFioOLP/7TCA4brQM55aKW89QNyNLDqZIZ7CaPvEVt
xDJN22/YAccLxDQyCK5g709MPxMaK8oKLuXJyhqvTw2YO11u/pUXuReAaovylYSF
yKC6algqy+LeTusqhXX/Eu05q7cbijufV9EcpZhfQCVWl1IEp5Ryiw/wxL9uMUJA
nDoqtnrAO1X/S+WnMOmmN6rFCVgnDB/o8zuRttkcUgsNaAZmRCegWB2k06kUrhuf
6H6BK5z1SpslQpCI51zjL6kmBVpXjB9d7s+M10XSe2gQGnoUUH4aTmLandD8bYR7
13xXJ1YLY4PfFE0eV3b8rMSQhW6Y/ERtgnAa6/6C2p8/ASQhe4XEqArsKWsWfcan
+8PaGSMNOeawscmD+q8u33o09z4FDJFCwANcp5OtCWkea+UVvsf6YPgwmQ+eUmpU
+VZdXXjX4rS1hrOdDnRKuOU/wHweT6i+XCM2x0A03SSXTE241Mg8WgzFxatbmgdN
1jVDbSivJlc3R5Qmcz4HOWv0zLWE5i8QyVmr1+QE5E/g9ipbRU6zp00Co8X5hLDs
NspkFiA7turxxG7TKYKLwpu+ItkbpM/T64tCyMKFiZe9XFyN4qK4rrRMss9czNKY
vtW/tjutisZUHAmIZ4Pz60szsbbcD6RXqxc0PIfvpBFnR+PD6gud2AR7z4TFr2Vm
3eJuXTobKqps6Z+/ROJX9a83xE0Wk2h81oKNuCikLg1GeGuQRm/yQnOp+GnsBnAm
EvaHzeqHcn4gG4IMoroV3cSu4qygqmd4aEX0HlPbUheb2PKkhLjJvY36Zd7dni4k
OCclB2+e98rrlWf/VS1gXlGMwxouaEWFfKFcH1aJXshG/MU3mIw+GoqSwko7eMky
CzH832YLrfOqocUNZNrCVd7SZdFG6Of6i+KA6kVtMpaJdqC3OAaPaBem2+EtxR/j
jGJF/lbmfRlddnHUjl2NpZ9dD66HDajvCap1s22VapFQtW/NU8WwIU30bggmy0/b
ASj31XflmGmuzQ12WzjV9BqkZBmygDvRy6wpKTKJkpBZ8goN5ahfqjczjO4Wunt1
ZwIl7v3HwEyWF5tWsbz+RImzAJCPBKUJdmdlSmOj9Z3t8LvMdiDd+9E9bloaBIAz
y+Z7OFH9y1U9RA7SjXDE3g7bqXhftRoZMwPBmG1Lyv8yM4Ob+PG0rg8FObwS9Q1h
2o5WwnHg8nWW8qnu924tSerhJm1RDyK6tYSgQ1GoXTRU8P0S7kU/Y6rj8iNqErz8
rj/jZOWfYa3nvk0AH/rX9jBxqmWDQJWjEqxnAlJg1Y/u2BYY2O+9Lb2uyy9HDScs
bi1/e7pfStbYnN3BlEdwQq9vdsLI9sZpCAy94d66WHShfb04f+xJfSpL1m7i9dk8
C005vYPiwUBk3CNx2pg0TxVBQjN8MTgz8WTq69Tdw8WkOhVo5vCEaT7uMJPcpCFH
W+fvvWfNSeJYSBwc3L3zHfqsD1n2SYFV0wV9zGzt6AJ+FqUH1ptpvqQZo7wNEyl/
eXoX6Z3QPrl0/YKOxfFZ39mvxk/Y3+oAAOnbRdV9ge9j+xY8yCWHdh2ic6XRw31k
UDlnGaOdCtGdF5lFFCZghLmp6AbSrEPtMDQiHmcceISj5l3YDqGXhRQDde0rb8Og
YJSaZV/xEyUhtHyw5wobrajISeH+Fd6GDbX88sYP+uZYGMMSfgd393je2jTD0zVe
bUlhG5RwI9/q3Gph5BunRbg15iDUgkjc8ryuLSW2RpFott9epkb+utee34nVKsFx
wLOPQRWQYFanMn/hLvClc2OQp1LOyNIZfJqVsAoAySpvUqGgeotJMYZ3KcMFo+rH
piw3Gv5f/+EqORyYj6bnYX6xjVGrDHbhHRJMdid/qT0a+Jce+bmcirTdG/hqeJ04
BV5GlFhvTNqj2470rQUDbbW2/wx9dJhheVs7WEoCUmc=
`protect END_PROTECTED
