`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaf0+EpaubKWaK3Fmm/2QTmDmzOxYMVi/58LUFqPIVwb327B1phCquleAMKEbT02
fSIuCyBaC/GrfbxxjqeU4s6OAZ0ulUnS7fwvWpWqV9hTRIU+GS/xtugqqWCLHlXn
78s+AJnl6q23rp75kIf+6guOfl+KEuRS3UyOohBqXQzktDwk6S04/w/fnPMbrj+2
+0gjvFtW1sbkPHQVJbiN4ikEFYid+bdy4/OmUMKuRshM+y9B/kLyOoXTaZJ0CCVj
lJdtYuW24V2RrRTgUI0BHJAo9xsDuCpZBvhB2DJbREm5yC6To6XS9i2AhsZMSaL3
KRc/mzkSgfYWyR3BmiZOPzJtURZHvJIK1t6QJtPhXZ4PR19tP/EvKtfXpSvZYh4D
pbuN9LesuV0eeP7yRvIccyeSiyP4smhHbRXPbsEiUQSCNvFDk/PHp+ZV7OQ51v+C
4xmnocgxK4GDyCu1EMraYJKonH7SCK6xwb8X6dRn+NpCY0PD1KRIt8ax0nGQnMWQ
5Dc0StmURGuWyzP4m4nPQgSBd8UeODpRNyY7iBW3czB+CiVBS+yANBnzakRW2JqE
VhhES4mivlKxrXlEufQaAtRJAZWc7Kufyw14KyQKhwfrKIk1nWZnruHBV4dgytby
`protect END_PROTECTED
