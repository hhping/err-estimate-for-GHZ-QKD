`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qtRvb3RaEaAnvuxm5N4IXaxVl9WCgt2gl1O5txThJ3uq7kp9WnwV16sYJu2k9wT
A7pwoNEM8ktWnvxJln2QaU3RNU/zkqH3PZElmGQ7MNoFypPTJh2IFe8iE4Qj6T41
OwzynqnASC6Tc6Xu3MiR2/YMSAFdRSDI7w81HE8iS9BmBffsOPHHwVFpDujNM3go
fcaIXJesgrk8aNsZuZUgq7t/iWN4DkqAtbpaBfzEuylizqPOD35dy2aeC5cMdIcl
ult8u0fwZFfS8BPQK/wtfLeoM1zr33pdS0NqMvP/lf1dVCG+X9H1rmO12CJQxvtr
K31TzC0yJe6p4VsTkcMRH0ybVLsR7AAQ8xW/a/ZatEszankqJy0NHy3j47uiliSr
Ao7v4Akz+5hs0X8D6evDMPmpH6nX4hoCHRBNWKdxti56l3v5cY2paLZoBqBWs/gI
eRLOQlW5qf0KV5oHPKrVIz/gQKTgtTyudzBLMiniif6iloWuFd0WWLpmxRrnrEvd
Viqt4U7FiQvAWKGwWHHiB9tZumTRR6HnSyJXeLRRc2GJG81k2Qme0QSacMIi2BlP
DAGixfJVBpQ9LfZannvkoW53rfQAexcLV6BI+YLkH5wYiw2DrjMHrStrXUOVCQ5K
QLRXCu2U+HSedjNR0q5u/WVPIN8tTpLXdgMP6/McR0V6Cc1r8RV7+Sqa7I7TVTVQ
6ZhmiflR3J0X/zp6qO/irI7FgwvN5iZgRYfpk4KZqektoqLQgA1Rb7VNCYoDEVrt
p9v+2FvB2eBCh1gfMJ2JmX/ALmjYul4LQWF1JRiFXblE4XOscB8ME/K7EeauKB2z
5G1NcEafPHzA+ZCJuR1GM1ojOHfuVFgQh4SROax0AIX9EKs0TNWgpNCEcrbAB2ri
nsq5cU2IXvcfo6y9GddOYw==
`protect END_PROTECTED
