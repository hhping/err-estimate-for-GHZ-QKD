`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ouqjJjko8kcW4m5nFJTDIZtIwrsW7+JHYqPQvZx2mMCTOYsge1SnuTOY2e0a/7b3
M5heoKQQwSPBsn+OWvfVN6WzeHLOL4ALkrhpq0akWwKpaPnKmvpJRN0Fbma1Rov8
wAWJYxoucm6q0PbPEiyN3+Ro9dyqpgJ0dLJ0JR+hxP/rYLyks6jOZLVy6QaXTYZ2
kfMLh6JYuMOJgjb0C/D5zGWybzi31c7h4wRRn7U8KYs=
`protect END_PROTECTED
