`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+qnykO4nJENaZ53URPGmQLrx9Jb1IkDgNt7KgdLrLz06AUbSZh4nxJe6Nbrhhng
ulPqH0cUcTh/oqPnTH9S3Jcmh2gpjSKwisJS7uNkyVknHRtVjCqdbTLvMHLdNtDd
OMcmm13PVDV3rFsoZ0avLqRIqkXEQjObv1ydLOzvmdqBTgKuLvcxwhRmjYEMyPCD
ls6m5EOn/uLku91V5spx91RgZwPfT5YZkPAz/CXQn73cWpUyjuhliOyAHt86aaVe
gkg3tpI+QwQ6LAm/nXyu8FNr5zKBWYkz9tTAuiazimLIBVAgSdUUyuHHLwQ1FHA5
IM38R6crAYPVWsBGC8rftHtIV52oT/JbUywwQc9UlJ0OMqhoukdWmFYltMjaUEfb
ZyXIhwEZK31jm9ALIXdsstNG6Ovc7Q69iKUxQw4PfaMO5OTmFfJWL2OrMw7pIqtP
rN2TVKuHAabWl5C6IZ0SnTCZAc1xO/9EgrbLCrzsnokGsfmbOFbZGt4O9/reYS/X
H+TBiie+V+FOtZOzE03F+L5f2bG4Sep8r7BTEdIJWOyAb6J9RYy4qGSPDP22w+5+
EuWIB0wp/2GFZFuLrfIP7pUB3QvtgTOGk1pS5ON8X5oMHaXY0fO7jIIOxVuC1nhc
FD3qJ8Yh12qG0SsAmzh98/qSAuO4MsPfDygBWKgX9IQwPh2cnjs0bVQYsSuyaNHE
+t6XLDxJ03XMMtuBPV9d3mvgFstZ9P+btaYwo6Kbec+oOwPSiTisAUVW1OcETMVq
3g598O7XyMxo+HvURRPrjmqPUb75SJwFLh+YMIjnd5PicdmsTVyayqo8wrHPIkHu
pB7d3l3X/OZCKgl+yCmzP3d2ZnS/D90ipSvQL39NEDI=
`protect END_PROTECTED
