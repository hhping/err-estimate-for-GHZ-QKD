`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sKTw0c9sc7GXPVa/VUOH0WeuemLf2g59n7tF6K7zN7T2f8wPSX0z7r0ZWpPQfnJy
lvKmZKyH/jSgG6kd3VpEyX8uJJ7noyDXhKKeCeS9Yi+WMZuiMqZNvupeoOIs6oxM
/j00uryp+UYzDKaxfoG1LtrIkQZafLpfXJYOT9MZ+NY7ppTDJ4pv+4+AV3Nw0zu6
sA9BkDbmJWAfiRKzEENoElz5Cz12MM+4lrQJXlsdIuiB9TBNUv3zS0cgLiCO2tia
BUCLxUa01F2kfhV9dV+UF7NZgsFzykZSOIFZ7C6P7hsvB7T7FnEuA9QJPxGVpTrY
n0qop71dCF4cjfzHTG3lGD4bwDtsNu4INl1JNGRxUfk1UuD+pbEHQ+zzoOP66SiL
l+MUBPl6RGhfSz3IosNKUovt8M4acYiSEfJV3TrwkQl5WaZ3tUuq7urJXkXF8ZOD
6nJQ+DtjfFE087ilDU5ecxbyGMktaadZa++bHqbcs30P6mOBBgvCqNrvkboWZQeB
JiAB7Fw0pKhVpj+5fMQX20jmn/vsmVAxjhk0qjgxUbtP/XQfkB59vGGqkrytgpig
S/m4Jw3JjbxzHs4DJoWutnAYUo1zob7xD2zopQ0vYGJzleUScIp1sA6MMO5citf+
zmPNw/7/bnairZCzlZ2ubCX4BM3EtYdXV+wanDnmNm9DxFQ/C7JnWeiD8paGQEXu
oGkTB4BwSNQyQOrKUV3Rt1RwwgRwCbv/q6Xz7i2+GaKB8x+1RzRk0G4qmNMozBV9
0YZKSfdSJ7HsNq25t2D1HnKs9fiIGGUROOVd23yctwUwmvDQgcE4AyqgvreJsv4k
xPqtO7/uLCHVtnB+E7KGFOcBv41gEurX6wFW6v0LqlEegy032SoZwYgs+L5YHh5l
EHwbbNaqJ+Kh8Yg6i4OzjbW+Z96wjvvku6Jk/SMgqCvaIyCbrUoIq2w4n3GQkOOv
mhetTTa3BBG6aEu6TINkHjw5DRcjlRIl43Cb+kR5HyLFWdWNERkPGtR/DiFkhLx7
wn+k2tVcfBkMxJHzlquVvnU33r+pZlL/xOYa72BIy7+d1h3wPY3ouLAAIRSvj8Fg
S6M9Tmk4GISA5wfjE5EcQcCmK+ml4wu8wbyCnNbzwLOpjfeDkxGrLm0IFbAqMnsx
fhWag3jyZnFQ6p1mmSM3lM6GlwzZkmtHwI5k9H9su8/ImGAb91y21+qbtxStDvtL
RIaIRJ9X7gVxeNZTI2TXVuuU094EIuR0PpOt3+QYnzNoIvsnbqKVwlKwEDyjZziK
r2kNi2fgPfqKgK6SaTVrr1UFcAZOMQkyBOSrCenz8t1AItFWyiIH1lbj6euwrKlT
V8N+xNO2SCs6IaZwp+gF4olFdmK2qgmngKdba40kgtSpppjtcbeCnglLR6vH4J1F
/YKtL+BU+yZ8zdkoC5qaLSsMmd1EoO4yvyPb3cfThZhXWZaBuxKri03kqyTF8gz9
tf52/Rq+RtUAgXj6dnOfi+BzvcReTDlqsekROPd0v3nWQPu1CDpEfHUguGpCQy0S
9VXnp4a4Den4wTwquTfyhYI/StaSjZ5DhIzDBrmfXG7JPlX3dpMN0WQ23Qz5u8hy
xhD6SgSCMXFXquwGsnk1L39e8OEiifpTf2cSqTqtdhTnYniEDPD2SZmmcURGjsec
yOBrSfjVajsrPDXPLuJjGpUjoQvA8YYdRWUICKrDZ2n5HiaPrQu5pNsaoO2CTDYr
BksEkqra6Pq0+Gr6fT+qWbKuV5GtlSjxeebERrRu2dAUl9tm5NABMOSpotsvHC6e
a21hwPqc88Wx9W5HGeXQ25WN841TOhj0HM/QIkVFA3X5Vxz5wqvAv8ZN1o5MZMqi
KZArdHbGgqtfOThjWZzJhPB5FIdjR2BHoo/e0ytqXxtupmzJVEvIluT76z+V3Be/
nCwvtWIQT7txN/SDzCCFH4MQXX4vxWQ6ZZ0f5j3YtA6A2kPH7jrf3oLu8F7YNxig
UQuDMf5im60GqAqG6pcEp7YWHxv2ihbhgHvH8Ku/FAFuhm7xw40dkwIqKfFVw1dK
nze1/PAs5NI1S/TRzr25IfuQX5wn3Ph22OGWJJLrFkpTVj3L6JtAh8ZTgr4E2k6k
S9E4bvVAXmpzPaC+c0aYf7yeIGnkPNTJyzYXfUDUQ2yKMuAHaBDauHIECDSoiWN5
SWWgeQ/SQi3K90TWSzVQFi2TnPzM9NO1W/RlEimigdg4OGRk2VkpNtvFfViv/tYO
8NbllAsJovynbUTutX373+Nrb2tr++AnB9wHVGndpJkctzAY6AzeNzewpEQiws5m
zI7+LfHJ5bw8cYcGxrr3MNpFRTIHR+YVRHxO59+R00hq7ZilNcXuZAuzzGcC9o/w
a1z7BaZYohmtQgREKTvWoFwgBEu4Q6q7sazo9UCRz1Ov3B7cvcE4KxG6zRaebqBi
HiI+GgIoRsY6vAcs4pELsiuEp4O3niD3bme3ppha/nif+X4Gc1ik4YlYzjJX6sKi
lZjeJyem5CIWiTIJloZxXoMlbl82A/4Qk436YZv0ybzK9vODKivu/l4jpCYWNRUT
Ow5aqFUFgAc2MhNsG+U8sq1ZV6d73iRsSpBNaQ2WhkoCotqt7MfWPK0gADaO5f4q
argAFfMqYxWkYjcsutq1luve4gW8yq8QBf0ME1ep/OXbKONfJFek3sT+V4Z68gJ1
uxONrlmQe0uoxrdYtKF7y0kKw3y2Gemu5OjBoQ/72xHdWgZQ+zoFNDt3tjWBDA+u
ulndFjyZPD4CRFhSJeOla0vzhuu8j0bBKGlZPp1Y8yrF+sfIab4IelhGrZwjIsyj
rH0jwBy40ASXR3wxX6fBfm6PSPPuYv5yTet2+06aeF/qI8v91L2vUFWyQY1dVyQA
O1jj7fjY2T5sUQBTAhq6eutSYkGEHDv4IX730ogk2rIiY6NkL/CkeCaRLvaAZlqP
fDEleRLnfXUKNjuq+iC0sEidUafBLbLV1WGv8UbKeBMmdP5ccoV0kEKg5XpW1x0u
aFn3HMVlSgpvEuILuzT5phVRR2HnkLKga+HKEi87TuDutQOxOezJak6fa8VWgsO/
gqS6R/auLjricLcB1oodB/ktdVbdfQ3uDmqyGLubKXIfYi4OxSDIIvWDYstosXHL
oIhvfeW2uySdfDUDhl0pbKk1Qi3z6v4Hx3sNUolbQG+6CY9yzpm2wqp1Mwyo2BUG
va3cdeJ3PW11ROY1UXY7S+czMFdya7ruUeYWixHqr5yRTlgvuw+lzXoPVxGuSh0P
Ht4j5CTJT+T3z87QimxFSJv7dLw7hOgQsWD1BtIAnzmOuVoiod31L5jiF4lCRiG3
I+F6E59WyjHrsx4RbAaEL4A4IIiSXG1jXkMb7WzN7w4g3v6hShtzHESL8gjIICs2
bTiNnfyljneQo4LiZAShJicUCHpX6uAnWka3XhGnuAsKD8wBAP5TR5oYKgUP6YIF
hvlWjfnK8h+X0JLJMdHqteVgajVAVcGQjiGTcvQWm0iH4LmmJueGqf5SENZoUKqS
MG0KtTaKcpSFCubFimW5oEQxwKKymYnm6V9pXw7oFW1DF4T4oWfE9rn4kpgByPsE
jA75Vt+H0uePEbW5DIL8bLG3Wto+WfDGXhZT+ru4qaOb4xkUsxI0sSAyBPx06vzQ
vIytSgP1gB2x97VGY8uHpjjPtMijQeL7GzJo3u35t8wUdwJS8EN+uwAUaRKICmMi
LjxFak2PIL9xq+oo206G7hlN7MCyRR51gVl2LRN2CSK/Pw+0539rh5A4dQGGPrn/
Es9XKWwHZS9f6U+YhUM21TQj8O77VsDqxv6vSPiiJVxRF9HSj0tUx2cgjPYtaS5/
APOIDiWcgAHqmwWaIa93Ye0A36fn4KnTCG3DDK2E0drZhVeAG2iFCdFfdL+DK4HB
G24gU+fnXORO+O1XTl4attEugcOKwNElsLT77DElpiPyDGKRVdwZvRbSppP7dNl2
b927EKqPGJ3Q5FIfCgsrHDFqISEO5y1pyFCbR1Is8WcjQrRP4qUGk8Zk7Q5u9e5b
/W8/XItjbr4fFsBbteB8bd7l9W6ZXMNMR+Ll6FhRr5mUIlfpHn4BzrgBwVysICOk
qaw3WuTfsoI/Lq3q5MWVh98e/roc2qGrTM9tpTAG6VA1Z+NRLQE+3CZhwD3KTVBF
BtCfbmQXA9OQUJ+1V+wttMQUkDcqMeBPGiej1DEaCIXRfVUzXTYuuz/5vYfT3DcJ
NTlQ5RMRsCUWsACvfHA/IILESDPlaUYUWDk8W4wOeUK/RXxfmCkZ4s16NL1CFnuE
WwmS3QdpUmv+bfTFJ+h/c98aTY1flJDgL7UGv2Is0C0JyZ31Enh6rMWeXri1Uz92
vnm5Rdyx5WQLfU9bbm4/uNBGXJ7N2j9GI6VQ7TyEp6rHwH8XM71DArgLYqxJ0Vf5
5LM8IMWEgat6W6PO8tFWNfxDu1iphw2SYNKcOYsb5qipysHuv+W6EkrcP1vOvIdU
lbOS98tWYORL7uI5NVTtb+CYXxrOLuLWlGebxsi+slzIp2z6O3aM8YLtaBtDygrn
wUPj26IgPVtkiNl3ywDV15oaozGIXnrfynahZx5RnH6NdB6bzP18xl16EdXLlVGQ
WUxlAAZvNWcA/9GRuLMjxFx4RSw6+BVVmd28O5036fY/fnzrMyZPx+i9jNQynP1g
bLu5O52GzLfK0x5tkHDT+r3C9cggtckWIMrbQI0yc8REBqsRh29ToZeEa/TEqwBc
c3zwCqW7P5Sqpf8elAL9pAHtH184YMgQ6jCca75wCJZr6aBQY2bYROLtyY8xAaTH
uG51+yU32/qC/FWSET/2oH/gpwHVNpFl1lE0lnCB7RFVzRQUArjXhR5SjUs2kkNM
mr56KU8jFy4xtgF22c3Mracli+f4MNj3a2j1Pkv4eXIO0NHoBo2Lny2yJsBQmL9F
TMAhySIS9aOg+tHENxCDwvtWg2U+HdkAu7eOmdQYneB882f8hCk3AKdwxTl+e78x
EretNM8RwrjOEDSSz0nwkAJHnmDuSRc8V50Es3323YNOUYZknSdBnuYb0VUKod7x
AymqefDCjAdDme3EuRP111TJQcWxiCTThHjW567NXlS+5pEKrAgK5IZu5NhTdP79
ITqFzPBk66WIRNvBxVwLFV0RZmYyitFrBaF+ABkVIooqIEtmZHIyp/Q7ZpOIuB85
4gIbTjO+6LiW2k97QhpYa/QUH8EVZg7ogGmG8mnAmfsxsgRPmU91WQepr6NDoo4s
j7szKEpSqo3QwaWvpud/EeMQsXuA6zVxthy8QDLJXPDkGn6M88n+W4ncsrzKJ10p
qhM5je+ZSjiqlZRdJ+UoMyyrb6HMf1T++ozYRK5Ef+YClB4W6tcEhe2trQUDkHjJ
uyU2+dYtLQxfrk8aG7a6/+zhKv+bKDHlxZMrUhJwYRJcd5gptO6KodWjvddH4v00
UGTCuIuv+WAQCdF5W1mYiV1d3ZQKA1tSrmuoNVsuhCBN1Tq5CtWqpsaHaz6ErOPl
4UndRDWFWUzJczGREvFg2gBSd8/VwuoP2vx8rXlP3/yiO+hsmjWowkiOYEa1tLuK
s8IboLzrwI5ahW/py+5lGAW6vPti+cTAIIjQF9KQtaXToWc2rTbSSDUh+i8W5rvN
inTLDDvk9a77iq89fCgIDHBcxxosQZF6LPLhzT49H2vEy6GkrT47jvn9lEodiDvG
VjuGCpFqdtYjvdxjdoXGHxj8LN2HrT8S5GWrDrGZnQjQnIfDvqAqz9jlcD1F9EWv
2nfplcvReabLsaFg5JJ0v7n5OmB6JEAQLn7UbKE/wYEofg0CXHmuhv8eFAFA4TCg
rJYgnHJEPYSKStfzfn04g/eYl3aptA0m4boYqLp8iIq9d8nhw27WTUUmXQRrsp8c
vGDG0EJLFT8+TeOLIRpq6jBlehGD8cLZg3kp4cRVE4l0sQOuC1l1Wl20i3cbqeoM
UkgxCGNHBY/gMLcFQOqcdGB7CeP3ewNUEP7SAK43Hc6FT+K4K7HHM88V9b2v0KGY
HSzmY1cDcRm8lw5NZJ6TIeeuwLjCbetC68c4kL3uULDU+ASNY0MLsbYplYr9HTW3
kyNfhaHqRHFYLSmdJcLZwHT1R/Sevq68d0KiXsbFyaFTWdhvwz2yQ6k4KIH2V8FA
/KsYlgRkFQj2rQwsWWUgzTPqsLzKnpCBk/jBFoKwxhiWvAZkMLpYlL6zlpwA9cSg
PsuNQggTnVMmPSp3mceyrMuSm4kq2mp+hNlj4tQoXuOzZ3g3frcwmNoeX214p2XR
r3MO1tq+ZgQU1DIEk+/+9GYgK8ZKTc81HKUnAltkg1Y/utyoFEYiEI3LhNnvQx4z
B2f6ipZo+JOwEpB352N8W/TKhBbNWURSmYvxCouRNY9Iafx0MWHQLh9t9tsSV5p6
DDMhUXE6xu9jn8TsJH1hYnut0ozH3bdBSJ1pbLfKgRc3XkNlnZEjWByvBxbPIffh
rP5vlh63K7jMUwLawB0JUOTgrB0EUJ5/7pqZYS2rBHsJr/BTlc1NRnR5k6GzOGd5
IQxAJpvmcEuxS4Zp13ijTk1Y+ufcjt2yvPrcJD66nS0695J9zKXdO4KpfVvpq5HW
wD6mFept9IeQGJq9FXfmykxp0m4KHsfUBKyD6saMwPs67xMB3OsxZhbcSB1tt2tv
lOLe9/AmC/ZM3OtBGb/kw3IeqbiOHl7cCzlVZoHzEY/7eoINvySN2c7TRPT6OXa2
D+vX9kqL5RC1tfHZz8FmsMtQoLY4Eor++XP5tby2hMnxNzlQEnekAA6+40k77u1n
oI8XKGENSxQMUTV2ytcED0x1I/sQxgzHIwgD+8ygVEF5wBcaC/c7Ymaiu32b3VyU
iuGh51rDb2HvftE/RIXVnxkzYBAmery0YTSOLKrr7/CETNTR/9ndEkbhCUbXnTIF
FbzKKMclu4XUy1yDPv+oMblVxbwHCTRjwWCgklaBLAjAUh1d6opN1b6M+HNNdlqj
GwSyE2vZwNPCMUevtQCETPwX6GbSzNwwWPS37NkIAHUaW4JNc3rsh4+b8PBKdqwb
TEtlzO3WOhtbAZa4aDmUvS8hi1HhH2LJayvivuzCpDRUA0oB0zGzWddO7oMeqRow
`protect END_PROTECTED
