`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X5aq4TwPMcLRdR6LISxe3FwptD75HySfEc9AIFSh8k+uxPs6VwQk4KK9ItRTlDST
ngnfzoydQR5EQDlZaBCBIiyWwseNEaCRg+6Oaz6fGemi00f1O1trw6JiDKLehBi4
qmWbo0rsefi1mqecwAVRdLjT2cuXdXt5Q3queCjwKlbYlnZPwH9jqI3O6mW5n6JC
CYC51GeMGkeyMvrJfSnfL2G0og3RZE99VFlwSbxroZQMgiBaZXopNlDiGVFiPwCh
oP6tfh5EhfM2fls+7kR+IzTRPz2LHcpu5wavv0Cu6Lr4CGAkNYIkShTuAOq3nhBu
hR+CdAVosiHiNmRSDY0WN9tkHXFpxFUs36vteL98XfAiQK89+dFKbLEdSJLWD6oh
IePQH7HbG/t+lWkipCxeBbNwoPynlo43poG00Khw2DlTFIZALjbhXmkD282vWGFA
Hs5ykFu4PJr3t1oDVad+ob/q9iKsKQ3t7rSGevFbV52w/QvEsxr+KaHcEyGel3rp
7laaR0e7zRI8yVKrStsSqQeBRly18dVvk/41MQEHJBvOlTlk8Oayxjs0ZSkx3mIA
Qwr/41YzrYe+hsRrc3nCo7h4q80cj5FPxYf4951POnMEUCYpmXErHzaPqMZIMNyd
IrgoVyvlLI3fq+XNDP84IybQ5HbjmzGSaKmaX/cZMWy4KBnzll8qjoBbdXefL/8A
gJ6nHSDezvK1hhBdh97EdkPdvesmwyPT1MeNonl04IXT2iPGdJOfW67FgMfYqA5Z
+SdT+L6enLFOKC6msNzR3lk31rIIP91JQQYA9wh6Nfo=
`protect END_PROTECTED
