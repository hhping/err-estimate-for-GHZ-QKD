`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0nR+yuoKJ8OfU1nkVfPCHKz+ebFlyg7Rlt3MEjIcdtC5iygzSwNde2YLOob6PddK
cuzmjf7KapmpwaIC1vLqxUQ9r2KvosfytnsZrOuksUq66+zzyuwGvD3qf0mqRCR/
vUbO/6HdadbMWL32sHlaCZyWnHdNMlF+FFFEZ7zeBHHZ1J7+sqtVmSM686XBZvvz
hnZBoK8jXiYx7YAMj5hBrHimXCEVHcm893qU713pI6lxfIhybSRfDaAPPwKOR4ND
x/pYuYg1MYka4W4g7GRZiqs1CWYBMsKj8T0A3cDNpsNr/XSNvrkoxE3B2IMEDag3
2Dl+CBXq0OXpL7MuzTzk/DyRksR21lGZUT0Rkvqvgt8TwQZUniXCuwSMQ4Vn/Uoj
vnjynhHXrWuuUvtY/3rCD/Esr1Kk4c4qWnhDFM4gSX7CsRUHe55vSig7fNq6bE9j
u+a8cTPeE84rA5cwObKeI5Gx1vdzPm02qKE/SufmVnqXJETKhwBuWtWaylcomUBp
lYlfLdNa8+orQkm/ly7mMsQuwVIWSNmZdiv4uWpNJ6/EREone2Hzt1EVN+VIMYLA
OmA0IgDzIXBfGd2Eq0bUD1CP6NprvtbF7izvO0t6za7bmcaH2P+Zw1btietFdaQo
TuaOBgdsn+NArSp88AKuWF3pv9lGLawp642RKWflDtB4JKVapC/zdgIvorEjq38D
bfpX+hjHI5caT+vgRVNt1l7N4cvFXm6pjHZ7LwvBB2jp7GGrSrK5sXAalF38OIlz
xmkteFZRGKAiVv5KM1O7x2IWi5aiKyoaGS9bvM2Yn071k//hVBOEGVmguWRpV6bM
5nD9DG0j3Dbgre7kXh7C1aq5Tu3ZWpzPvzYUSROqSIt+F4IYfmKdZYE1s5fRAWFl
D9LqSJOPfDq9OaFG74caBNiX+tgzyzxYaJbvP6JjvMtp7Q2JrTdVld5bUWcAlOzT
7prBLzoTD0PK8NUlAwx1JYWOm4UifuF85DvHKMthUmux66KUSgIjJCn7Hnl2Kdqq
U6/48ka0OvdrFMWTP4DF37BkLOJjgjKmrE4iXgT7wJYdkLaOIX/0PwkDeJHP/i/Z
S6HD4WjXCiPkk+AQhzqlAAWx/oQBikOSE8+z30nKE8bTrmQgJflqSbaTorbM/3Xp
KNkAdcOufQbnQHIzYDpNcF7qk+z3Cfan1Ts+8Fbw2Qe4ZLvn6WGwcOnsdqXOK9ci
QAzDmmpADisAniGb71BP/Wmnwj7cYXnChkHEQ7juJHInt/+J4HiXW9EwwLUHW6WH
okWdXTGQ129B7HhMSWGjb/v89GVeRbtaBv3qGSUjJK90B5ABE1/yHIhG2KRZkC+d
Arp2M9L+qFg4wNl8JHIm7rUdS/HivzDbqDatuArse3RlObQ+filDT/5hiWNltZdB
jTh7+JQbRLj2lsSeXDo4S4FuHk7BLcA5B6Kq6Rm8heknCpp5BCwXnm9c5swwM+1k
KBPjvDDAX3PK2owOuFzPAPYUqUP2vwn1Vggacyhr+R1CyLEtxhB9hLU3dfMsIgda
qzJQTsEl/RTKWdUOZseqwJiOXonvB/l0XQ56YvtpMLfPJkjJ488p13OU6gpz0VHy
eompcpP1T6xbQuGhEqtPzymEOs5kQUgu1THo6aOKAyL/voD8U/fGOISc6R/ROuBv
l5JR7ZeUk/KEMV5/nRLyWVodvySgfThW6vsh/pdtbDsynrfL5tDuJKxkzX5dEzP3
rvB4yx3qJSVlH3tCYYWUM5dLk4RD8QQ+UUDcX84009t+QqN3Ff4vdEdibW5J+s2s
ajuZZnQ4cWrg9hOUArblhk2vmV3+3o9Rmg6IjoyigFjMwGaqDkW0y81qZl77uqvV
nL80R4crzYVsJrxeuAJgLhVERtW6PxxwA9FOUvtbCE8widdDj1goMsa8XrqlAwAX
tf7rC7ll1oIu2eXYhw1b3mYPvPO1s51ctwgI7CV3BTLEk8b0i2ev1h7XiX4w+ALR
aVdwkNt5khJiZr/R9Bg2x6oRE0iuEunbT2gxiebF92VVxD5Anjo0n3j1a3CLtXY5
xPhGfQ6mO+WlJaHxBFROb2l6K6Pa9OXvLOoC5zEDa/84CMELoaeNCEcMCtfruTW7
GDJbWaB0O+Yf4fzKbf/kjxscNTz/u72SX5//RnRjPuOpOrFvM/CpvJEPzvls8G6o
zjGItD52QNScxFSxB45ssP12t5/qeE4dkZDYQDS5h/qZFQO4On0I/PbUyrvxrEjd
xz2n98UuHNm5DivBN0xxP32iRL7QvhtZw+xjU5VxY5D3umdvQq3LIJVZYSF9lxLj
SA2NKUcZKx83Nm9koQx0kZbH1QU5vTvvAjc63jQF1kexh241q/2duHyugcviQF2O
rXB4HcehfkiVgQSNxfZto70TmgvA1N7AxynklPCzCwIaro3QVhcAkfU+RJIw8Gc4
yiZ5l2T0UM81s92sSsY1oKN0Syebbuo4iJopMROIl1xFMGb4hIPrmohTk5s+S+gO
UverikhNnzqrMJB/rAooULaluKzmM0TbOZkSDNSpegzlma9msNh/pB4EU+ycyPh4
xMKIitThALnbzYdtd+vpI3u46pSY5yoLxr5VvNG9MUpdkUmWnTtgPAB6Viy8p9CN
QZFIV9dUIhSJMu+zsv21+gS31x/PjP97isxjDLAbTvgpJ0gQZhySMUgPvUfUc3cX
sK7cX1AeD3aB7V/p/acYJQwGBIK9qA5/7MkGpKAhi7s1jqkSApkSRWFhQnJ81oFf
X3DpSZjdKWAYk2NtKzEWpU+eKtwHF4z/bhYlrGKLzRxSGy4f4Ea3e7ihyudnGMQS
5XOMaF0PxTaUkzz5wEoKeBh1ZzH4IfuwQ+RlcLVddulYOs0JWw0ledrjbnUIykBz
j3GX3nIeKH9hG1qzFaEEwNHI9VWuOn+29bSuVaOcS/lszzoZGzwJ/HpmpbIqbBK6
Qv7KE7BcEqvFGPvRIQxrtqOL3wPYptBShw7SoLI/xYh8FknQvWLkdu2C/XToKz3H
NU40p0iOlCGVFmeZDZbdCUmg5b63PtjNXnS8lrcQWVHfQSAFQYSa8JW9jQrfNdsM
R54Rqivi2xxCSGLoiqFvDkFH6bZzGjGB2evlcXLDvp+/I0VaAgdI46AnQzy5yxLr
dOgFJ9PDYU9URA/Fw1kFR4Zc7SST1sQ8zrcbX4ADXcs8UTzrW/A15MbHYAWJIAC3
hhe+ly2qrlzD7TsP4R3qXPHUXjqpCcxm+ahScERXTf7HG9j4Rl5I9gxi1dv4NxtJ
3gi9fXiWIZjuG8pzEvvfKJfybir7gD1yKT62GdfHQ8y2azU2iMfwPPwd36F8MsSw
f/Tj8AEv5oqCeikYZ6J6OE9lmIrvSlLf5A+xVJPvUldWlyBOV5uW/D7XlaDH7pmh
hj9ZhLcXea4vVd0ReLaYweRaU3dbxOH1lYZEPwJoxXpEnI0fmLUZMTbK4ndutJFJ
9VgRW1LKAT04ukVqC1FUVKtuEYJdqykrQDaJthPDRdWAvNLhIzLzc69y9cLdcMaq
Ve547sb1GrVaWRnNVZ3q8a4BmlmyZKb6Gofi7BdqypHaGh9mt/VxQa5R70w04QaL
LJh2hKFxQA/DztX7CVd+VEMYJt+pdCHw9pLcnStOWPKR0NSppGGzJNCKJ6gJmqrO
RVfWVKMCp2sC8+GSZQKBchttptxKb7Xi5n0byTJ7475GvoDyHoAGS2QHT5fbiheC
GT6CY/eHe1il2FcpqMxPW0yZXTHBbd1JSZ1kuyl28BwRisO3g1Y1m6z6BeFJQeRO
9CnWg+K8noc0uOMmgxaB22L8ShmdpXEAIx/E6sR6iKdTOmcf+wO6LXBGAmiB9nAV
kWMIbvoj9gDusQhMTGTuUfyKExfM63BRtK/TBeout/ND9KoMhNubKHpiwvZVcR/d
f/3ww85fTCaSpeG3UjMfnF/TkTHlCBgA2fOwx69xq0AiZAHgK0s8eMupYERlkFOT
npHwzDZMuUKAdAOwk9vcy7clL3QUfxX2DY5FSLXVB+QWXhnxv4v8Ft4TRcOr6hdC
10y9WTiiRld3+qf6Z5fuJuQqKPl+D6czXzooxWZ13qsy7bEju+fZKH8ch8tQzQfA
iRM9oBltfHbutuLN5OAGDtYjMnNGF2+MbIWbUedgmGoWFifuJpoE+iWLmMX4M4hd
g9/URbISIMf93I/NKR6p/1Jwml1LoqJZ2mZclp/SsnTjjCeAfZ+3uRc/qcLG74PO
GKXCs1NoFxMRd0HxXiKJyKsjMyXGlAoT7p/IMxpddOJhQRPQBpA0yIPop+sg2dwK
5sms0xG8RGKzxtsWtcXbOqtYOhmRm+bQZbybWEk4aS3N6jMIJBAtT8EyFFmwhrIP
Fmm1xjMwSkU9QlDGc1NJYG70fXMcl2yJbt82hMHWqhxS72c4GG1+8cEZNpuUN7Ay
do1/oF8QM5u5F/3vdT8yoI3mfekDfhNA2exRfqexAEGqQ+jcMR6ZdsT0PB1e8Qdu
KhhxtajnyiCedncSrJtFwlQw1rq/G8ZvqmX85zVCkCBNSFKO3Bcw8sQLE+VHWiNj
q44wke2vS8yM0IpWNXJ/YDZO5tDwGc40VOFgHQIZctwoqtb1djZ4qLW9YaWGsUj4
c37g3oydm7De5h/P/G0GCQhxgS7sbtqIH1x+NiaS1ERDCs3oWDqs3EQgaGY+IlfC
OCcnuGKRJJcU5hW8bT4g0qnWTRYkD8xLcz8NcdouKaR2K+R1T3kfmtUHvgobAjkV
pUvrcCScq3/Vfem0+kGFLC/wZZ7ANnOHifinHiymqYMaB4YJvaatZpDeASOU3F5z
+a0PPlyXeNYb2vJU0PHiSxozabHvITnnoAMBl0yFdWcT5TwHAogbeBPUk5UU1mgD
sVwrPqtIgO23Z1LbDs3jvAHzJapBNQj1bJyCRsr9qrdETQzd170OD938LbZ5Uelz
CUhuZaGGGYC/ao8V9vExZ3TzAuk4lSmDrT6FZ6VX6W3bWYXK8euOIFQa3tnxLS3m
rXR916UuxuBQxCZOwFqXEIkWUroe+J5RWIUUdR2BtHwXyVe4CoQXVtBUQhNY/jtp
cJYfdrNhKPTvsWDt46MQdaguUF20Fqon1FUsSuMydDmKthalQAlrWIqfbN3gAgo9
D8Qk5zH/mVqfx8ELkeTvJwRZ1wBrQsIqZrwPdgldNgzC2BSYE15EOkZL4OCTQei7
mUwteacyyi8fndo99ETVtPgTGATtmlu+djSRFbUG8CBzZenKmSTeWm8oFKW82ZjN
ooPCZL0PLM2EWKWj7rEbUGXrnFdekTokhMS0+mKubRIvPYSDjRUnwo5RLfhmCgXs
zpD47Z1JRuf4sHsrhHf33dXv8kuVAi9daqUq0HShQFLJTHLvfQKZIpE/1PKx938R
GLXlOPffMKNfQk4dL4J37S+nsvKyvrfWhVFsy3vIhbfpj1WVdxfa48S6Xd7V4zgP
/04Zq/34rbDGhSkihMnRyEtwpGhnd/OC6cD2DECDkFC9Ig2WpXTbTFQmZMEzzhqA
oKit40ACWEAPCl/wn9uxgdxMNNoS3MsVXSH8QVjHz+FC3IFdtVPwAWn1JOous8A1
scQMXVHsgnMaaLH2u2PKw2xukBL874PoMQlKRSmkBw7ewsikvRg1/b4GwqUfiX2Y
gSPMXXm4WvNsCFnlAs1DN6CMjARios7EEyHHJiRyY0rkAkz5H+tjU3zxRuhm4UdI
Tun08kFJGz/Vjel0jLUlkJYP5q3C9RJgAb+INPjqT3DSW+88iXk9KC5ZdwCSI1Uc
Hcs4wfZASkMdD1YYFBpiyLWlzHMck5NOjuDdLa0PumEJm1rsCsJjmUbClrry7WgZ
B3tA2swxIv658/mJxzfqUErBgCKUxkTun75/xBXMCLn3KqkQJokvYHcw7ksAPFAB
ajEumIY9M+HhmQBC7+rmss9DBFXKK0Uthhd86teVwGpFuc/t/9dVoPOzCaZhQkR/
Oo8PrGfsc8evhzV8Gz3OHjXt3zpmIBIjGWtohf0oJs+H4xyu1VQGEAVAWH9OaEjS
9Zof+svvjZZc10IKKDdXOOXsQdnT1zcCahOzfeYcgWhY94u/K+ucaPYfAn8Q1I3n
lR54I6JivPIiTRtOdmD6Zw==
`protect END_PROTECTED
