`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVTGrVgtdl0NlMO6HKgK2daOmSQLEh8NCkhJJ5lpdoKeMT/f7RZvkEV6zQzkvHDy
Yz52yATVhlmMLKJZz2LJCE4/1eeBSKr4FTOjU/n2VbDC6ii1rnDuNBpl0IL07+gj
v4daNBlHJWKKmFXhuqK6ofA+yzhCdj55pvH6tANpuvikvUS7rw+/45RUiLF1F6ah
EdFrE76tOP7SlBe9nmylySlj2lnYFd+jQIMiLBa3+dMrFx4RAYG/fhflD4wvVp46
JgvZwR4BDAOLd/J9PO/Dg3YlnwohLAsf7znyJBO1SRWwT0wwl17GPDirpCcNYrbV
+RQQ7rW+aUQJndXwnY6ENg==
`protect END_PROTECTED
