`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZy9x15IpVNxTaayTsKkXHw20fvw0m05FmLeXZna4gtp71whWSFJLC4Qu1JHkjTh
jnz1OL3Bfl+FOODqTKGjdVnO347Jt30bNGaT34CSZ5sDpzSRzdiKjymbC5lxsDXv
Y4N7O2xKxGznZakguIXfCEMTStpshjeEXLzs9nG8DpV+jxLF583yyfH32GNAVdqk
t0OjSTZwcgCsUALVIFIZXiKp19ltDYnj1Sly1fOEqmxM4NeUn02G9l8myVdFx2N7
LMrdhRA01VTtlUxzDb9m26Xq7NvP0iYQlZ6RXYpWAP4krQT/pOIHblPMZDADspae
80ThTXfoBurVaRiDgm++QTMOQpW5jzIXODJQ6L5vQDRV/I0ZDns89xfzeKs2t8TL
Po8V7ETtL4jiL1ECi9lpCALTw1PMT7JGayQPbZyTYx31YAzun8XPGP9fgNqpjSV0
LR4eQIlAGhPCuzlZ089CvEALzzt3sHTXEt4YnxMuAFDU7HEt+8SEVMVBnKdc7LHZ
dSBGdQw4MvdT1sdd3cT2sYMZJeXSavfmmIgXEEh+vWwvBJJMiosaBToNPD49oRZE
E8gQXJulq9VoMxR5FMWDwLhQQwY/FlsIA3TsZN0j14FN6ssOa2ZQiCYA7GZ5nWG2
wjI6kIrk45ffIjOPqgXPVYJo2hJ+kmbSrnSBfGyvJlZ9a3bO5a7C0d+ADfzclVXc
BDgvHXFXzDm1aO65iDr7b1bc3BKONM8oSeV8k5GuyQk/m6PLXaXTUTFpZI2aqEEl
fq0ZZ9kTiisrGqfH4bcQLp+T6J4aJ18Jwii/z8OO3ljOr/c1p2gZUMOmuNuvCpUb
xRKRtiH8VHfiJJhql3i4qLFp5pKpUjiOEbgT4pYwAIU5fF1Ujn0/kF64aN2TM3qp
m+ToQ6jo1Zpywspz5RAAoc2FevgHpmNuZmnkVDLwlgK/WmRjL2WuqenNhXrN/h6V
B556RZX/kE9XqdXr6JxLFl+AjpJAs3f1oSQvweGyyp42L1Bj36bN7kyp8SLAG/Wk
Cb7m1ZSZtKygazGgs1zJAePLEnODO9j9CIX9dm90G7ssj63Qu3Wno8jB306TgsMq
pYtOUip2zccdUF3cD8h5sIURHAaS+T8dpizmMdOyNt4STgm3iyi5jqD1OOxSRcfr
GHgUTOxOiov9GFTus95UDHHwCGzAD3YXoQKsnel0YCVerecuBLtOUhfgiWxUc0vU
ZIxKL0UjEGLF6JwdHuMCAUoTGnjTqkLblAHBcT1KBUyAQUOgt5uXRsv6GTtAt/P6
fT+3yFgNeRFuYoeTH39WAO6vssuf12RAG42+vQrdVR8OrkR6sNGEovPLb02N1+dP
EWG7j5KTi3/QPs8yPnv/o9ut5twZ3tRVhfbfIa8c2UNR9tPG3Ih/2h6TyCu8/VB6
zwb4LgW/Jmz2eNapquTL81BAGawOppqhM3p+HUHn3qI3W/nGmbJ98+L8BqofnFx3
21GUW/BV9eyzU8rvnALgA0bZ/PAMsuZrOE9uv5ZsvLCrP2QZp3Pm/x1mC1nbgYpj
Ny56keS+cW93dnY6xtXmt1nlZmuomU6ugkYLauNRJ3EV3tCEOM452178ffWq6hQF
MrbKr4Rcwk8ql2lSbc8/zjjuJ90eI7thliHiE2pvreVuhRRyLY0zybxa3zTs6HUG
arSaD4WtZLEKNYmbxRH7+0zyrcWTRz8HIYj02NxeEPbdnLf4U8HG1ML7FwaKDtig
/0tA/UaGPfpRUX0U6PA1MIk2QdbDRj5GGW5WW/4b0wh7tgXG7gNBUR69BmJPBbET
wHS4tSsWnVTX8gcPG+83EYZDq07oVeleQuFNWi7bB5oVXtzPmS2OmB5y0F6Jam2h
E92c5HVNA41Os1rPJRMXgsecsP5xvX0wHeUx8qbiW8JCpwVACbwvvnr2JuzjWCzw
Gi1MHOkS6iIYdRT9ZOb1yTmrIG7o4i/R7LYemvKBPgZsQVE7PsIVABErrnD3n6AX
VLHR0bXwrNuwq3VsfLtm9LUogWcXxn5HWiIPNeX9VNR0hTm4RGxzOLFtxDObnwQK
4qoy1EFZAmOau4vZlKkE6o9OnqjcLbpxgnYTARirI7hWyiHh0CIsgWy5PodZ1J+K
svKyxK/XVKFUOnTJSs+wz+CQBrAI8HEg1ek3WK9Fmiznc8FGCsv2wnwWnZRvorvZ
FoOl5ysQVbM3f/63Y1Pt8v4yFdo94ZynIJzkrooX6hDUhLM4rz3hc/fBMmSsLdQS
N1wVazjF+KxM45u0luMtTAK5oo9AptV3Z/YzspQhUsG5Oawquygs+OpFEAI9KsPr
ZBNxo+SXAupJJUSPbPtsafb7GakMB8kgPknysUp+i4pWYfz7VbFthGGg56lfSTEE
yrpjSei+g4sz3Ruo7C+EJEf86uXCQd6wZlPUg/mFK7fs9ihWxKqg4jCksXs2Je44
Y6YyHD83a1DiAg9RlsCfz6M3hbzxro/fs9OA6PkkYI+hgCdAoiToRQkOdnIlfVvc
cwe3Cmb9Mv+gvxVZYC6XFzdnOsgPiAZE7Nf6qLwyLAb9IvTkGB5V69ARFFg5a7EO
8ZXJhHB9nco06B5Hyb57zbdi27EWon3m1iDuhR/rtbfx8BKj022+qQBJsrO1mVtI
0Z+pbNbSHruS/Zp95FrWeAG9oRfRUXqwYKupxUKNwuvcsvNRxDT4k3t8IFbFl9xz
ZaJ52YAwCgva0yK6m7Sp2gjxm6FfcROId1tLOXm22soxrpdME37CsA6YyTKXO+Zc
NDcinRKtbEcn+mtLHuDdmJVgkj/AQPcMbA37m+37nsgSzShXIZcpb6dvPretqIny
jGnazFvJO3TApTivNNqXZgZ9xDx/QXxcH4Al9jmyToYclWcD30ZIhR7A0lX7ZIY0
PippI8Tw2K1QcccFvs27xm8xGcFAnShfwGRkBPCBv2baFfRBvaTTQvJHNAKudEYt
XrjZ/nVHSZienXnmI+UTQR9P+YcU0XIkiQ/WMAQxJgXneTN6V0l/P0crQPoS1UKH
9OoQXfQ2tnr+1Lq0Hio4XI532Py7WGfzskjwFPF0HVuvN0bFqeC3fqkOLXVzE1Fj
7nZ6jELogeZpAtPwnfmIfzc5DhFn8SWjP3WaePMuCzmBtiWRVzIvcxq1uk4rBowJ
leiEkk8l7SRhjzhRHFO4IZh4dqXdkZ/quLFmoHl0ORTK1+O/bJA02/nZ04iLmeNH
ssrv2+lhhdGzpwG2rNf0oV/HduaOdoFDb9QRl/Ly/vMmRQxSUcHKHrlRAyN1nZ38
Gedm8RfEPHQgPIuxDnA4UOsCw/vm3NfLMxLvJcIlNID5m6EXfchmtC9sZLBXyCNO
2Xsg8eT5n5cu2ZGMCMLXAGhdvhDQtECGrZNvOf93siMN3LooqG+cv3aEzEi2dsiF
uUsUVlTqcCCmX3aozdbdQvBp/hUiCLnMnAIH110bWdq131cy1QjudxYpkgwgd1cz
gGQ8R7ysvLu+HWyPMX3e+E5z5Onx2PgbAYhV/b3NaemP0ITIIccTuE4bi8cP68U1
tKqnODrI5oOeYMMUzdqMkX56hrXy6IY+x9scAv1huXVzhY+2p/6IsflcKUcNUPDd
DOOospQ7z3KFHalsa435BzzTPaYOtfhJGwY9eDOeS6yltRzbGmB2pUIQxcNl8j/t
TXEkq+v4GAVEteFCR66MTpoE8OtNF+oG/9nI1C8FHex+mmUgoqLfHi+1pVSb22rv
FBtD+ImxiNS4pwf4C1Dq+KOUhczDjLCAnLd7eZKVLxNlvVXzYe2xOvPRveAGocwA
S5MP3whcnR7tP+voPkPD5rR+9MTgDLj4S+DxDVSKJ+rzZGuBKr3Higk7zGhBvkzu
k4Z98pg7xKKbQpzcuBHmX0ck3Pdg7v9v+bOTrJvUb1nzNppVMXLYUmyZ932LPeot
mvGXNRE7IroXc7MRD3LKz5LQzhE9OC19rhcxLjE4kw0R1iknPSfeqpAsQLqrQCfZ
8gUaDRpQPoCfcVu27md3XQRnhAtnGauTMQqZUOrHtT5t4kmns3n0yiKpCU+THoby
MV+EVWmhtDOouX5HWhgg8XMplgZjqLr4KGk4rHDiXAL0thETYIq63cDu44kGicIh
vUYJVDxMn3vD5R3GjT16IITtVo4zApxt5SJnkF73jUNh2aHUsSGppHu9fx8X3uP/
NhWLvDX0o4IRi+DRViJJBE/ypBftSuDJYD3ky3Td1sGcdz52ItESSB3rLpWkh/TO
eXumz8g6pS/z9hEuaU8iFtXiLejTkmrr0VwbSl3FoBZrj+yGxi76vKwSFnoCZ606
c5rtz7W+Ryu8jlZN0m7Uk4j0KCZhAb2YME9yMo53G8OZQYIAKCleJhzq7OclqDuP
oRCzCMVdLdDtL/ri5hnngsUIEkcQiIh9K5cmSBaaN1R5VxAtiEC7nNp+KD8k/xhv
1r6xSmufC3jsuC4f9zumD0lzvw3kpL9QfYtFOc9RtoivpGXhI2eTnack7at2xJK2
ynQva/4pSiyskXQGvwoyDYZ7nFhtltFj5hUQPJ8B2hZJnS7Rn3F8Sm12kGa3shS9
XZGMBjVlL52OoNpSgtLLoWXt04SxH1Zc/22pNVKiKCU83DR1Gnh6qTrzYS958vjs
QZ3Hfy27DHgfg7Q0j6nkDXTUAbuxP7zYrEFqETsbs/63B9bBJMylYhSE9XI0LBPV
xFYS9VuGINwcp3phELczHjUHDH0iwvBzDRyZiPieQZSVmS4i70HhFjv2tErI4vNd
vHP6t7p1h9fKF9roT/Zl8YhsJGWMhGLKizS24m7CFkxq4nIgUzUZwZhGxI+RRNVP
4Rme+ZvRRrUfslyOc1BotUlglTiOHj8YnpJRz4owpOuZVoCwEKzVCnfy4PdrzSc0
E5dEzuW1SsZ/p0zKqr0pql8Pbs3JXsAkKJdXDUzmW8tArGQKb5ElE+YtXn1Agwhx
9mlw51S5lmmggIxAW6pwrSm+SKH/fboMGuKH/vnT5Q/8UBJECCcMAIglIbkd1rQs
RlS/JmGqZ/S8fdoWgRqmMycCaAUGYH/fydFHUv0s5CnFmDAck2oXmRujJF09SEGm
zIwYuBoOTKw3NGEBXCfkUnO4l71vGLH2qMI8/73Z5ko9zk1uPXjcDFzStHcWyWHZ
TDSd8jbXua/7tPz4RhfTuR+tjt/BFbzkeSlqbD+PWSzCDLz+pLGSNQAnBEzRQY+6
IfyLKmDIuNiAXD7HYI0QiwPs6Au3UN5dTUbmAmdDP1WwV1Io/7rey2ud1N0Ue9+5
sPZhcuqcoUsjLr3yx1oTIPAlFzh8GrYb5HNggtn6hPycGDfjyOYzBN6YZh/wr+mO
XaglL3PDzH/4DTdFxHgO1EdS0mVacXP5gTBYI2Muydp8gDGXkZ9QtP7nE9Yiolfy
bglENlAl9SxFM3rBsuhLLikHqVDPFDgI3Tal5PlqxYDp5RQUo+9TSvVEJPruAG79
bDqHeF0F6n4iW7C7t02iobc3JPOniFYTTGXwSqhbboNlI7rF3F0kp09ISncpIfPn
qDaViNy4h0ohLpvpKStancI7Gm+WGqYTBE37H+SL6RL3yrhD6j+lHiEiju6IqFne
QhxAyRFwF+Hv2HHwjW4SLIE0Anu/OzUZJ7NxSHzMV5IdiIzDW6Q/Mf/cht8YYHDT
roHVYfnY5wghW2klyNbAeoH5SCSlqyKhGDFNixSfKlhNzKWGWwVZZwkoPgNsY4L7
EMBTYKTKm97MDoxjHeTJrKAY2oskKK/FwpAeqJjB6jls/oLY7YGp+lvLYjxwaEfs
Iep/WhGMGlqrXUHbYaiMSFYBKh0P1GZGNFeW4TUZREp8ylu+MXEbv1nWcVS8USa4
CtXJFeGgVa4EmPyMcKKpz2o9Dxqgj90ZIA9doJ/Wx9zqvi++HuQUO0G0Y6IgTt5Q
qj8O79V3Nz/RkXtEeNUz7NMo51SxAAJX8iY7QgxeZf8a2e3HFWA7SUSde7KQAc/3
+TBIY8j6IesyRSEHmoDBnThhjNLOU4BGCysYN9fzLRSd49UrdEYs5ScsOcZVsnTu
+mvqcxz4d2vb7Aq9vVWV1ZDyiNaHPVAMELLPLFSS+En9Trou7655u53nqBdEnnV+
YFOStsYfoxLrHcoi74HukRb0McxWkUDRhHpbCwMSkfhCkF0l/mMdcROeF9ZVQsKk
eJAjCfF0DczMje+WX2AdyXaTURGB91bNsawswBucSF/tPNpv9LLMlhVbc38NyfwG
67vLg5kMz6BgBgOsAfUOEGkC0U0Sxw3aTe/35XlIT/qaFaTBw087eBxP7AG493er
/X3vimMm5AScXJcBIRctnvQvfE/KxA44C590Pg7nXYcRFep5lwIjRyUNUblrbwT/
BK2n+6dBI5Cmg4uLfSwSI5BRbdkcTK2ndb9GZuT7XrhV2+UFY8B8LDNdVyUj5V9S
0v2Fvxg+SImxD+OVimE26PWmtjeMorfwN/wRuP6Re1ubP+uO+LE0cWYnQSrT3uOw
xVJ0Cx556HjpYMpft0YqFPoibdND36g5HbjATHw1OnmRgP+5ZEMXRvr+fKH77iyx
tszsc3qPhFNeMAe6i7qInWIOwfBkgUb0oOVhKu7MCcdxSjHxjqO1AoEPRQnOTXG0
W5NbKWOuA5PsUKmbaFr+Ctr2ckFGcYXauyk43RMnZ6EnHTcZ1bns9dQ8Uq3dYx5F
iTI4imXnSc1KW1VnbPo99gwM/HVxqa2nvExhbUjLf7ATJE30ET5ao+V1UPxIxMGa
n3WlD03JPTynylVmJ32zcIJol4GwL1ZgmOr4OFGlDK+bSkLaqBYu83K2k2zJXE+8
B+EVgJPvooTueqhNAQRSQnq1aJYli9+kpqI5uqdHHmALBWmZSLz3Y4VNw9nXrnoI
+YOdkYzDbjz60a7fR5uVTXhDpSD/17ROqYEG3k5QXYOZJTCYg1Qo8S/+o4vMr3j5
Usr8HyDWtpN4C0Z42HzbwbHbbZ/aNGMLADK1/gwk60JIVIppBpCdgp2NEtpRGLwr
ZS5KrHYPrkG4IfK6JznDN9fP61i4ukWR8QHyPXyyvbpsx1V+qQlXvncJU+RMQEAQ
dgefHzBxdXT1Wc0cGpRxx/TOC5VaZjc2fFJR0yQE94ZSube1pr5KtebgZ8KfYmLO
+NbPxdSiW9aH4I8Rw6QZsaTdc+uqhhNkk7EsFYTZl/Jw3u2aAT0wEZFUquoISt8z
va5k+l79noofabSXnovtZpB5f3m2yTKACLUjB3Qw64tGHqhMjKB6vcsw+naHbTqt
NbiAN1DvjOaqxBSBmwVUWhj3g78kDinOsh5loq9P1R/ipisOIxWebxfRVyVgAhuV
Td2QppbCjkuUKqO9BNgiGTRnVcPj4MGJjXB/I9cD3LrL6+uI+G7pefcO+UExY8Qc
HwAX6auIz49wbgLCNmLP/nl9ahECy2uw6E4ZZc8X/bQMRa7RHyQJoCjNnSa4w9mz
Ke32LGsHS9vDPLu5LWxdjGUOEYCzi28AMgPyHu9mEZs6m0LPXamw3b8bqJqk91nT
yiNrzppq2VxLYj0tq9V3c6ky8B3bKgDAP2q1pUOwqWv4M50hlw/U+MV8mcC6hUKn
F8ZIdiIOMaqyXaz2QovVsCEnUhWAk6skhb51W/YZpM2LSBfs30KJRCI75Q6moDRW
eGZIkSK8e0XSFfXgHFHBEf1/GAX6ls7WupNISJz3z9bFWMiHZzuSF0CG9yEGFFFA
xa6c2LHZTPmq2K7u/UyULfpmee66ceHSOdwhXZSrLqt4GB/WFztnt/tu2wv6nz22
Y10ic/cqhgPxxTp0ANsKoD+7XRXVCMaet49CYIkFN5p8xBusGfx6kLaIZaRd+ITC
9ZmqbtTd0MVE1qPQiPySQBz0P/lGIKU4xicnU0nr9oFh2xcRTUrdl+Xq0/ffEhXC
XZvlAUswtx4z4EYvSi3mN8tAKClcdEaMVHCs/ItTasrmipj5X99jnYrGnskFk1CV
wHzdIsedSujt4nAcZGfWFK6RE4qQpNm9P8bK9PNHC0elDdxqFQ8eKJjYRslmRKYY
twzOK8QoUZa3vZGbhiHs8XK5XWYuqtqAO82A5qFBbW2DAoPdESULsAtONq1PVCqw
7W3frFK3KdG17VOYFv76JBI1lhLwF21mHD56jG9ebrSNUuVM8vWuwXlZ236VN8GW
d9JUs7U4Y1Kjgj1yQDlrQxQ6cNn3ziZOCYxopigijdIZO7KuASl1T/+JXE7s8eT1
Wox36B6PKS6SD5Jrf7NKkOuLom2F6yYBHs5w/6aw8TGBUfRGa7bgzlABuqDQvWIj
TMPK6Lw9AgxGsembqMlqTMQh7F9EKqzQC96tR/IItWasV/weVpOdUX9yZQ+6bl+2
iJqgaxUtwR4L0Wfnmwo3fZclm7lsV2m/FCcMCO8jYYKpavGGNoiC+ihjpj/MOvkC
aDBb4TZPunZcKZyt+ur/b7srvojZZSl9cw6rSdk06sHfuPc6O1gk85+g43queTYZ
tvWLWIK0p1zN+a6UtGBr5LfX1zrRiDRgdmbC7zMQ9giwpzcuD6tGV1gNrrM3TUIK
OpSyePmeKa+HJxEUN98SDRnFQQ3Ks+p8+p6IKI7mtrslFmA4QJ6S9SbgdijzxAmM
GdxbP8Ib/W0DqZXEennhgoVIvfEawhac2YPiYNnRIcW7QEZRbQR79qktM9go/R7H
nWyj3wobh3F4eWpVZbykjkzAAcWFzfTSFGHFrLcNz7CE8dIhyh2n275KgIcCLVhp
FyWoTpe2bMddbzSQaT+HZbEfpjmTHPY0WGkAxZ6ccdj0xQ9jJCuHVskZ0ALA+1vq
bXtOYtzHDCUjZYfByyquP0KnR6Ej/wMDW/HeJYbn5sjfWHsbxaEkkyUe2PsDRjlQ
L1ydAf1v8YrFotrn7//qiTHv8kmClP8RGrhxbqWcbxNs2pSsKhRb3987yzfCS+AK
8/WV2SxY6EjSK9C0W6EHUjc+PUJPwRDL2kGHbCAmt4N1Ye6+P7Si+Ru0Zd6eWNcN
aqvrk1rAr2CgcxNKti19DuMWEFZHVtuFlSzOgQtoihjHgt3MEXnz/GXuPO2K2/Oz
EXsYJ3pnCP+lzQ+aoANurSl3WRDhj/HqvzF7oWoebj4NkitDiz4eM+0eCLODVdzR
669yWubQCoCAZq/Mgxy4aeqCD67+7f4S3CSZYovlQAK0f+bU91ipYmzgkjmIoAkW
ApyktW2MRHmOf4CgfbunfvPaxKYqKTiX7WWd7Txumq8jtJZeyQ0tTKQrv2OrI+81
nADdqv5TnWKmIEl7odJf4bo8gnkiHFqkiQV0Fq/3mc4tNNcibSIJjt8g99a7diwy
xAsIaWScxQsnuXNiQRnfaDyP0IHnZ/X3KeWJtdrVGt8LThWudr7CqYtX8djd96Rh
LW/uXtYkQkKFAuPxksm1Y3qeyvj7sRFVqhVn4iypo7ufcIMUDIsxONQ3cmu1Wxar
k405rZgTXbX51aA5+i5hxdBpjDl3N8x9CjQ/JsHbDTgHLFmdxj6Q9WakHk0PlWsi
KSEdgTsjEL/eGq2f70duRzLj7IrF7/f0//kpICxnuBsYKrXBT6jcJqqVkhDGOJqk
dDJdVqvB75l0mTqoi2Nt8zUECPY6orYLsTlgkL0cCgmPX+W8NL8jJkXzzL7FiTY4
W597a2mXc2wrHuRRe1dyRG9gA7u2elYzSDFqpYhWDJWki8+4HdvGyyZKynn3eJtp
c9hqmSp/yx8Z6r6S69K7rvffgYt0GsYyocBu/ZO5gY3zB71HWsMemrLgEcRAu/bS
cfMW0sx9Rtuygg1SSJZv1fDKy5Jy7i7832//5vX0pdOYwfOFFlz8nAbsWwSbQqQO
cci1aSh2dIM9ridYvNH1NoH0pNZRj6oGx5qbs9J8cl+mdZDT6HK5C5JpCFq2teA5
4aLnrn+8lQFHuuSugQxQk3x6R7kq3bW2wTHDTpybqWyCN4OLf2D7kk3fIobwQzwM
WLC28cx9wwculsU1IZ9Lr8dzzl+qMQ2PJtjk7A/JdvdKjfI/UF0rc2LPtg9omEri
mNObDdafhTDCaz7HFegmKq6+PYtha4RYKM0oc7U1ZJQzK0m7qqu8gSYmZm7h//9v
ewixaARB9jFO94hnNtzVgv0h1z1RC44ZyarXAQhVEiDtgQJMVOrCwl+pDb9554ZV
QMwjCFeLqZ2GtD/p7G/58A==
`protect END_PROTECTED
