library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_gen3_rx_pcs is
    generic(
        enable_debug_info: string  := "true";
        block_sync      : string  := "enable_block_sync";
        block_sync_sm   : string  := "enable_blk_sync_sm";
        cdr_ctrl_force_unalgn: string  := "enable";
        lpbk_force      : string  := "lpbk_frce_dis";
        mode            : string  := "gen3_func";
        rate_match_fifo : string  := "enable_rm_fifo_600ppm";
        rate_match_fifo_latency: string  := "regular_latency";
        reconfig_settings: string  := "{}";
        reverse_lpbk    : string  := "rev_lpbk_en";
        rx_b4gb_par_lpbk: string  := "b4gb_par_lpbk_dis";
        rx_force_balign : string  := "en_force_balign";
        rx_ins_del_one_skip: string  := "ins_del_one_skip_en";
        rx_num_fixed_pat: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        rx_test_out_sel : string  := "rx_test_out0";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        data_in         : in     vl_logic_vector(31 downto 0);
        gen3_clk_sel    : in     vl_logic;
        inferred_rxvalid: in     vl_logic;
        lpbk_en         : in     vl_logic;
        mem_rx_fifo_rd_data: in     vl_logic_vector(39 downto 0);
        par_lpbk_b4gb_in: in     vl_logic_vector(35 downto 0);
        par_lpbk_in     : in     vl_logic_vector(31 downto 0);
        pcs_rst         : in     vl_logic;
        rcvd_clk        : in     vl_logic;
        rx_pma_clk      : in     vl_logic;
        rx_pma_rstn     : in     vl_logic;
        rx_rcvd_rstn    : in     vl_logic;
        rxpolarity      : in     vl_logic;
        shutdown_clk    : in     vl_logic;
        sync_sm_en      : in     vl_logic;
        txdatak_in      : in     vl_logic_vector(3 downto 0);
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        blk_algnd_int   : out    vl_logic;
        blk_lockd_int   : out    vl_logic;
        blk_start       : out    vl_logic;
        clkcomp_delete_int: out    vl_logic;
        clkcomp_insert_int: out    vl_logic;
        clkcomp_overfl_int: out    vl_logic;
        clkcomp_undfl_int: out    vl_logic;
        data_out        : out    vl_logic_vector(31 downto 0);
        data_valid      : out    vl_logic;
        ei_det_int      : out    vl_logic;
        ei_partial_det_int: out    vl_logic;
        err_decode_int  : out    vl_logic;
        i_det_int       : out    vl_logic;
        lpbk_blk_start  : out    vl_logic;
        lpbk_data       : out    vl_logic_vector(33 downto 0);
        lpbk_data_valid : out    vl_logic;
        mem_rx_fifo_rd_ptr: out    vl_logic_vector(15 downto 0);
        mem_rx_fifo_wr_clk: out    vl_logic;
        mem_rx_fifo_wr_data: out    vl_logic_vector(39 downto 0);
        mem_rx_fifo_wr_en: out    vl_logic;
        mem_rx_fifo_wr_ptr: out    vl_logic_vector(15 downto 0);
        mem_rx_fifo_wr_rst_n: out    vl_logic;
        rcv_lfsr_chk_int: out    vl_logic;
        rx_test_out     : out    vl_logic_vector(19 downto 0);
        skp_det_int     : out    vl_logic;
        sync_hdr        : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of block_sync : constant is 1;
    attribute mti_svvh_generic_type of block_sync_sm : constant is 1;
    attribute mti_svvh_generic_type of cdr_ctrl_force_unalgn : constant is 1;
    attribute mti_svvh_generic_type of lpbk_force : constant is 1;
    attribute mti_svvh_generic_type of mode : constant is 1;
    attribute mti_svvh_generic_type of rate_match_fifo : constant is 1;
    attribute mti_svvh_generic_type of rate_match_fifo_latency : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of reverse_lpbk : constant is 1;
    attribute mti_svvh_generic_type of rx_b4gb_par_lpbk : constant is 1;
    attribute mti_svvh_generic_type of rx_force_balign : constant is 1;
    attribute mti_svvh_generic_type of rx_ins_del_one_skip : constant is 1;
    attribute mti_svvh_generic_type of rx_num_fixed_pat : constant is 1;
    attribute mti_svvh_generic_type of rx_test_out_sel : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
end twentynm_hssi_gen3_rx_pcs;
