`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UaWd+EP8wMACTO+vGK6H3Htxd6IsVso9MRCfkZflsA1SdlO8CK3eqeIsK/AVXbaW
uXmFiStK2jcgw0veWPWKIu/9Z+JUmE+QJFF+W/XHPTg0Gk+YgY8nHQ1ho4F3EC9v
eWAwL06JtInu4rlKsLEtda6v9HGJM8+NHtgTMd9WznTzJCfDZNla9iW2iyYBSN5I
MykEdlGP7Tke1SQ1D3llnI3nGJRuzPFDgp0GNdQAvCARahTfzeLe4CiLcgXAoFkp
8FnMSsqfV8sHHOD1dQg/8bBxJdyy9na1+KYy/rUCectJe4wuJgzvkN8z28nU/VXl
dKcWl3fHWKYtXb3E4eU+dg7KumfMfqs+Hj99JI5L62dlwDtb5JVLWjfRMaUzby8b
bqCVyJyPHPY989QhvXoTGaAD0q7yGfx4cYDrdsSLjOuQF91+oh7WaLt0kC0DkUI0
0mLx6eeBVED2UX4UiXhxidYxEJ2kMHNX6xKoDxfHshERdD/ml5R9ayTQ5s0r9dR9
fIaOH8mrw2aLy4RGxGoBXSk4dNmUzAWtUMjbvbRggrgU21dl5SoTDRQuq8EobSuC
Y/XFye5Krr/EJgAySMLfiXAn6uiZJrgfE753Uv16eysCus6BZhDKAfD8oZMIWeb/
e6TYfAJevGiOTwmALBRs5qps2wL4Xqm2Pozg1S3+X8HBZQJJ7aVMDNhuG2k9ifon
FSYrz+37Ga8DGWGg5e/8FToSS+CKlt31C3xwooNkpgx2WnJz0/sVb3Fgf/P7dnkW
Pw79gpbx6Wg1+4lXI5Qa7CZH32TNgwzi2dcSZu8yw8dwvp43RSaMZxxFLOJLwUEy
YGznXbxikmwXUpcAC+6FjJIJgJiTDNrJ3LiSBNh+AwGMx7+2xtTpbU6jYX0H/AsZ
YoYWJx7VtWlCjxyyddcRVU4QZxC1YEf3aNKelYcQSIXQ5WUmVBSONBmkVyMDT3eE
FefZCLjAY9LkQBKAMIv/V9WP3aqUEz8n36eQEO1ET0g=
`protect END_PROTECTED
