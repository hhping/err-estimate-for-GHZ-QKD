`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDJZLFRfuGbiJby6vU50nTbiqHPQwMfEycJ3pKH21O1736YED8wonI3B4Hzl8JVZ
zkDv7hdtYiN4LmyNL//RVDkA32/rs6hP+JZexSJ17xqdjHpxcHQubu+JeiZ8IpOT
1RaVNHHlGdNwTvP3tCA/ZGN0fIQdxyUQwJUpDR6/kI2iZH7i+KvEiZtYdMgxqAAP
jhwtMK0qyRiPQyfanF5WDinCpZjfeZ0BjLu+jfMsMJVzotXUUik0qLhKNK/ioFsI
sNy5jb4qnZooOkJAjfrL5tSBWH6oFY7XGXm6lT6VXu4JHFSvjgsOlIGpIOYS3W2g
IAjkDUnDqCD3ZOZb8e1pywb9HDNVQWuhX9vtCkaFj3cCoMj/O36q+qfVdGHdd+rX
BWJZngixmeW8oI6wNu2GBUNk9bCqIEAtWaQSstwt2iKaqRn1a8SAWycugL7ObR2t
WkU83ylLLHJKDR8k58KUGbPHxjQ/zPIon47bbG1aicqYyg2ZYFROh1H4lLL1zqUK
xjFSAI68VtHots5Ed5gTOGRs1v3uSItzYOg0ZJX0CilgPUH41zdDL721h5fedyPy
imU44L14xvFU+h41xsOgR3x2WdVW3sKIcz4lFAeDbLKuiyRG0MMgR9gEHCX5B3NQ
5fG38qsQ6krc8RMPbBxuRtpFq0QkKukSrAZ24Kv/tHyJAKA8qursLY2jtlD9RyWw
b8Gj3KjBussdYCwA3SE9E+VD9z5cvNwxL12rKNNKgImXoACw4X0YaVQamMIIT+2Q
VEGJv1eMK3epq/atQbE/bMkSQ7dOwJSjSjOPtnaagAQX+JOHwX+vOIV0YaxmdNNO
KYQCw04GzKFkcwgnvtfQeI7vdMBGOv09gDAteGZxu9jBPR4yXuw71Hh6vz6DG2Il
ojTAvI68N727XL9/uAxboNSqMgd4kWf43/VWnlqwEAzv1OodCVDSYJKprFmkLdEQ
nJeYEkg43SQ4QXivwuO+/ngEQp6Xo/m6MQruX3Kbz3rkH8mFTtFPX0fqVoNM8b7y
zgFFeDnRDQ8g8qU/fHPb9+HhHyz7J1wo1TCpE602a13uanG5GtT75C76SEvyAZ50
4LZnnjAUQPdh0cGpOnhNIQ6/7YpQ+3wsfdssLCoReBKx5PNw6PTqo1bck8UItvQs
FNOw8Uiv5dydeIbcsBJ3AHWxcpMhCGTRbcHWYF/HPt2e9s9bfkP4PLABjw/vPyaW
aVaW6lX6aeuHdaJeLj6r1Grb3xiBaNvGhA4vMQLI6gN368q0w+rM/xirMMPzyOi1
uL7SmSdKA54oOURH2DRG0ODasLEdiU15RVlptHK+cEnwBCPYNYeUWqYtM92eHDFi
GD+MxF0xp/LCzwKtkuXqgEYgcFxtMG0Hs0G1PaZ9cY3BlHb47GI6t9VynlOGrZRl
gctyol/yZSatwn9Rg8zeIJJ0ncT3ZYsl0MLePKp0Bzx+ewLS2yh086vYaFR7rLkP
89lRN0GoQ6IrbUCotbSVqOElfZZiuT6l197wA8tW3f4ceBDYYqXwZH+7HxWFVxz9
fPz5i2jaNrI3N9eALg8aThQ6vx58eEkaNiGl9sopgbJ/XOI1GEJ22OPCqREyH9T3
0oD2M4u6W55UcEFbG0NC/ba5wsAM4pESVPSUv7WUKd/OIVZOMw+bhPJUzZ+Yx4nu
6DSgbW6mUrdTfoMu+MKuazdHNBRkDg556Tc7LZrQZXzP1hdC5RbHaVc8fZA7MztG
B3QsFCn/94rebP22b1KFD6qgIzP53NAb+r9Cj9LCgirQomcJr7WsQF/VyFEaZ7c8
vLj3fmCuPqy9+inrBdz8lhDsx/Ej+5Zsy891tGemzKq6Ei2eBbGaEYKGRV3AulY7
EktHbtwOvNOvSc7T3rErFUSl1A4XrwI1qGD/C4GMMO6lmBiLCFDgrT0ugrv4Edvp
5VoE+qku2go8Re5k8A93XsenCJ0a4lDVJTWRc9jYnakrWRxTB8I3S3bxaQ/khDF6
bmdB2ZasUevhX0hhWNJKutsYQTqfR7RRPdt18CoaiX72ca9iQbT7Dlhr4RyCrDvY
G2UlzSlTwhpCRNIlTTZANwaK18hDRqT87XGweZdJKguG6RcGZaPOGx35HTmFbkJ5
NH2PYdYHLA3t8T+zUm9ZiUD861vNQcOK7Qw6f6emdTUKH+FiJH5M8a+9WztcBD2l
3wSU89IgkB0m62LjqG+gmbE1RUc49KPNXQ+mbIFfrVN8uipu3XazU0YSBgswpeMB
7m+ms0kFOB+ZLQ5Ky7K9FsmhKilvxSguGjM7LWdCPWg8UXH1O4a64mY9Y6hmiucJ
JtB8Is3O+7/l+sWY+O+GLm0qvyfP7Qd+j6U16A/dABmieo40X5mSB8G1Adb0jcTq
r0V/gG1eGdh4aqBveEb2qPS5M8cGfFXKvxLlfTM8q+/PWa3tE8MIFx5EED/AU0iJ
cDjBKl0DqeIT3QW8vG+g0lUET/PkcjG9zjpTcyVFTdsonVWeOqwMRBt3JefcgYvo
Y50SfNBhenL5Q0t8cf+sNcXEIpyoUvkLkg+CNioW4kr0u1KDamdVYwbNxWKk1C+v
NTW5aTKy4BW9+FT3sSrgo058Gb/ap9NFOz94HBqgpTh1b0QVbHr7H+31pW3VcChg
WCJxWjOLMxYOsrPraDZOPmV3OKuwY3qtD24kzgfRpN0VSeH/xyCHF5T0cQcAu4Ll
xScYMprN0fNORm4pRyXBKwo345kjkM5+hXZ37sNhpWTiTYchDNfIDyAlKMQgNTRM
Qa1xWZ5/gFPZ8zqxeYuQCwMPOJIZXqyznFuTZ3XfiY7BJc09fx8othgSFdJmFQGw
ZjLXRwlcSh0wMCLq8PdI1nwUHeuC/ZVyC5EgIXqXDSmY/T2W3pMpO8zm4JVtdP8n
s9LmFJLDn/GNxYchEod7r3BPkFg0FnU70RS+4f+Y5etQaf6L25ykBB78H+QKMF2v
nz8sRHDXNMJYPrRxrK5ZtQSWwZcG4STQtgIC6Vr6CgpBHDZ9lPVJ+rqypyPNn5IW
0Tz+LQORnOamsmprzTTqATpM04R0YrlwjFaXbWc/ijr88/WWmN2+zzj+G9jd4bo2
T6v+4qsmSKLrfgyw5uSDJYWV+onbUdEa2aULvLEkCRc3nYcdck8AvjArIFhEjCtp
DjkKiYM8RS17v9pvajjeOL24LWvWnwFvPNaDxQrbT8U6iSKHWlCJp/SWCpzqvfZt
xdsvOJ29/iQ4midKF90J8w==
`protect END_PROTECTED
