`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifkSDKTG5cjd9Akp7p88iHrS8T4g3EX7c8+aIqSyJpd7akC9fkY2zw7R3LKgfuza
e4+ZcyExNh0bofIzEE4G6u7CR4chpurv+zpqo85axFXn6MZEtmTUkaonEV84DD5W
3io3uP0pGaZJbS+Yfy8whp2a41w5p8m1i4PhZqJ92SOLrISLrxjFPDKUDgXVO0/R
fqwLDcWOwmNaXzSPqndWPXm4dxesvgm6BPCdAQyP9vZ7LmBO9iFPN2iUj7lQqxFj
VGBQzjqGn+UZO1NEK6tj7xZSyvfrRQL0fURhl9Gw6chV9ZUdonVmX/ztQAjTKAf5
xSO49RbL0nW6S0qsuhFFMMmwlMBPcWFROM23PevIdJZLTBBQ6Bwiu0Wn5D57r+GJ
NKYJg1D5+pOLo2XOETjwxnPLniaOeSppV+SHhP1UXSIXp6Q5ThTUqhwkXA/y3lWg
3wKwKYciUicZI0tSdx53a0yyDpSrpJO5zzYkD7EoC+2+/vdDsDGjqCI4KoQ6VY5K
5AbIi/kOpcKWyDKMQeke5rnTzx/+4XYDfoluoqe6cpiyyElLbBoOfHtQY0OgIY/q
N2FRL2blnfL+lcuNJ2Xg9mctD5ZFXTZTGVIlXk3XSKZgfLOEyBuMX/jh5QVCE4A3
C69qFWuGeq3X7bJfbf6tiek3CGeEnHIS0zSNrBQ2dY/M/lswuyUvo6CLoVe6LT9f
6+Nzd5qvOsW/bHGoZsx3nX7V9FxpB3IT1RQyerX2BCIKkJ0+7vJwdp0ynyWTlAJt
Sz0oDSJZS3Sh5v151Y3Vo7PbZGwFQnU8fLhKgeWKiPlJgWJCprv95gbbyIVFE2K/
4DB4ZDK6xQEgiVJvzMaEMgvicaOd3/zjs92kMeCOAQMmcVkZu7cDV8DvV84L/szC
i55HwcsZu35WTYKL+1C9TIv2ECwMfJqHlK7owwF4/9o6LGskrqrQ5znDM9Br5Y01
7OzkiDXm0UU4FSxdZ8IzoeIBguBwdOeB/7YYuzfliDjOxfam/vcaTpAQrqTsRwgZ
813q8U0WWvyvfjLeuXFzf2QJLxXt76myi+Ycbx4j6gmayZhPnonnyM2z4ExU0SeS
jiYGQGhgQXi610xPvtzYJnDr8q5XoLLRPit+g/AM8V2aw/pD15uE2QlIuM2lcrfY
1+7ILyjNiOGeOGFkvudWbEnDnz83YLo+3ZjRn2gF/UtU0iM4upOkVmyV8A9ukx9r
h1zQNKddDuCqFqpm5AzRO9XCOmOurVoPETAgUczaK8siPgseZXd6VYZ1sJrB8ctl
+2MUeSgRhAAhf8JkxIJebHGvqmZCqx44WajkkbO/ufXCqTeBCbrg9Ar/yfmQ3Egn
rx+QvhP7uwoBpMEP8wXkud7vxItJB4D3giMFxJaAqS4LU6v2gnJXdgUv+SJjKpnH
eElwwIrjgHTvnFplxd/utWKl1qdF1TFy0T5Zu+FzG3qdNhTWYFeggMCfwuLtM8k3
tO0RnChVoScC9BYONkgntUTkFFloNFrvl492fp5Z5UwQReX2yPS+HsiF/UcOwRqB
HTwDRSy0uLbNPU26TrnTq/eeN6ym96Uawn2+DIjuGtLGbY/PCIerfE4bUXF1NAdf
xVTl2hDVpXrNGALR5R14KJwBnyRHYGVLBOYh/yYByLRbtDudOoyMygPJRk0Xm66o
Q0QmdYEr9wiUyS3r6+u93ACpjSdXNankqp1NhtgnuFnw9aVccOUtqFa+k01wmy5e
V3zK/hcMiGvPFN+qyEr4gmIXdnuJQAGwB0gG/Q/JzuRqLtKLGImGuk440qER3ey0
TVNg6W8JrHn/NoSoyHGmejGrWaGbD5FWGgHjMR2UwMF1zNyRKKyopI9bFDZ9o9Bg
8wacMvpsitt7I8i2fcdBTKIGOwwaLV7rQ08uaVibi78DLpx2GO+E+kX6SFfVJrxY
brZEq3l3aPZP4B4l037RNsDOwqILgSFPJW0i653mx9l9zNevgsWo6/i3Pvx+/ldA
`protect END_PROTECTED
