`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZVmNRT1o97mtCYxnjrolkdIveNirFzAfFubrg9WXgTtriC3gLq9d5AgmQqvhDOt
Ovk4diC9ozEvLKSGGPjhTt4l8+21YW3mU6aCIt7IfVz1J2AsM3ygMSPb82xY0w21
cd2tcwJqHkRvYhnheV8+Be1r5AFi8DaQ+2PsvBbOrkNysBQhNuiegFhVIrfyKIyh
skxjMc+DaJRPEq7Qlpxu5kbtyTEwSKxsV9rgrPwdIfONd6lqGjyqx9OqfKFrJJpU
oFaivZauJw9BoOa6vW6MliS0RgxbQ3gUsEXqGIa8IM6WkKn2cY8Yk37ayHKjP4vK
Yn/EicsHjWHkrapah/3bPSEVsmeU6sRnW7isuchdOnkZOnRK6VGmcB7gFF75HAF2
A77Bv6CLRscSOZvZGGXsVrROuaeZRmuWTHiaeQh1yCLP59vRlYjhScVxU3wlkxT3
SJK39YDvLzLO/N1IS3hs1EWMpk4NOAnFL5ZfzA2atzfmVpIU6MjrS+1tQ7EWMF82
U+h1+hPpG8FzJBJuFji7qNdRFxaIpNOpptm6g3z4PAr8dtppbo7E6mg3q0uXqc93
wSfaLYmnltUuQnocqNY/bhNs1MRQMjZwxv71mwsgdHd3sRhvSKBwGHmC7NvGYJsB
ZCNHepeDGFs7gU6ep2tdHrZWzFOBZhpHXBB8xlD8WuOhOM5ONAwjYmSzHhttfjFT
PO0JamWqDCz3r325MGrTUyho9yM3lQ2CRFzAvkxJq19MMrzyyroPvKetMzAvjtcI
`protect END_PROTECTED
