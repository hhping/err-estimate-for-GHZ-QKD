`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXAs0svLXTjLc/KAD73eNBJSgTWWhioA4VQhLA6PQbbbyUH3E+PX6cIf0uvvhTef
A8SRmqnaPrw3lM7nY8Jr+fckji5Wd3pRGWiktlmqIHnqdBO5sCETrtpZfd4spX9I
sHaLNi0Y84AbztdeY+kSxRztNsM+ax5/HyKtVoX3plabZXGH14U5xPKNoG2Wbdhr
8/3bIovYbv0Sys9V3vWXpA8qStY0k+oXS9Eojn2nmsjIgFHmeLFdSFf25wWJu50k
dB5rb06x9kBv/XsosPq+ShIO4Q0eURSLsz/VBfsLzAqGWuEnurRCkx8F1UEgRnKQ
Yi1pSLzO+gShN2DQwicovk9JA0DgNgcUuM6rpdzNP5FaZRYYh3nQAksXwHibuTgA
epsr89crqAAd/950bqWX2GJ3fByFWjMzFdg00QEyj1yAYqc1OfAx34KfFWgfOIdh
p5btbSqWuTDG+/n6d7ELhbLaTu9eKfOzsfs+oOrtHcf1KfuTXQJ1LMDaRvJEtjt2
7zkjTF955tmX9KqOY0ogJ+kiIgtO+OGb82kXZ8Kocq2mN+CYThXNEdjhydrMpkG8
0Yq7xjZ9z/6B8J6r0vUNJ8IuIqGtkjuvDUCInGO0mL2wNr8cx6Z4hNOvDOOwYdBz
ApbM/zQb8xvJ9QdW6O/4CoKSVYWtrO4szpu1ZSA4wH4BnP5ePDOU96o0tyD+uXEh
LuwePz8qDVZ5tWfv3q1BLcpCkgLxFWFrwDnfxaQu96Zfu8Rpe+z5s9FzSjX7l1sX
`protect END_PROTECTED
