`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aG3Ub/JUll/+wRK0yLqT89l0bUZF46+QvwteeA2/YQdA4WRuPWUZZma/h1sJeT1M
q0+OzG9mwu2gwsPT9hs74lIlU2BIKl1S90vYpAD0f766ER7yO4S8MyTkui/iVTEj
XxygyFxzG5ljPPDITG9xUQ/mXsygMvGz2S57oA3370iy8oQmw6eYuW4DhsmPFHTy
7eRRnsg4nKOzgFY31j63pgFFsoik6eHIhctmE+eAyWHFXghzNbD+TitSKRSuWJZi
Zzce7P2dYHKEzN6/sXq9mSTXZAYMLC/7i3I/Qmp/Pqszj+Y3bCgtvYgTs+VAv/9u
W7ju7nu3oY9+lBuWqcnTAnHiKThEa6zVB5tki3eH/+8aW5LYAsU89rKPDtCdi4Fk
tn7MY7izNg391KtZ2wgQzcYNlye0hX9zxkfTs76gR8HdCpmoRKcwvD9P5dwA9G0Q
egK9ccpwIUgCALWRpocmAN/LhMnYTPtqLNTW0i22sWCZQOzj6oascgjGg+mA0tVn
/lbe9CWrN9vZlD1y+pyONDpVgmPvyN3VGLpIQ0Vojdgrub2vClWLeCu0b8aS9a+g
XeFkw2gsQHbFAj1k08tKG46o8ctdgNMHblj1arGkF6wd98R1FVZMZgkJo2i0TtVj
1XXP0goh4AJv/yt8HdraVdETvTpPSUA22tJPBdoboQozQ1xpLrv5id2WOozpyMBt
EaD7Ky+RFHNa7pUOXRFlCsItODpbM8yqGHdimQDSCYOMk7XI86zZgU5RL1PeTEWh
DpbFJaEHSNX6WmYosaqG28Px9trQhUf4uDi8FOryDVCj+8QAj6c4TmrjGc8tdVdj
8IhuFCqx3mrRi5E2mHEP7AAYHOR/pIp/alzeQUN2jS2E/sCHKswk2wvcDCFKc572
bM1zQcfaXz4T0vC19bKnZ3G/gjKsjJSOW9Y85GFkSTU6loXhKPYApJDPKQ9AzYDp
zg2L54gND6IINueGbejtLPAzP498FkeCSVoK5b57UJbwFtJMvP/fTAR/6YgtZ05O
fm6Yx9PVg2TqPkfu/ZhFkoSZySI9twoh0AkyEU78mhEmcW+w5Uc5n5NuMgadUPbt
8+x1o8J4YmWO++LSprVuA9zWPne67NCuxdO0MZVqxHCiPPHaj20yp61SThWR2BZR
EfGwwILeyOVAjMQbRUpPmiIOkAGRhX3Jthqxl+lkfYTD4YFipL0pjVppWVwYRVaG
U1llmRanBXs8U7wJ1SaIdRlx26j+fP9PM4iMK5E76qezMyw//giw1cKCSfyeRxPE
R/QbDtnGIigokQiXnwIguB0mHiFcsN4E8RyX48MugW4m+UVOaAc7TlcMT8mVCu/v
iJYLByKMeVZRegOlWjFEYIBB7p1hO4hQs6sprhqna0mYzaFb0oOwBRUPBni9MjoO
0oLXqr77s8/mrRd+lNVmsmGd313BLEW00wzmI45tFqabSTyEDePUxGMQBxFrx4M+
R4PO24x4UxkFqCex2hWHBGfNC+FuLwFq+RBj9e31R0U5toMbRyBih6qCWdVWU7cZ
/iKtt8jzQyicSVB2nX8hZklCTRk/szsw0HHrgCsDUs0C06rHwduc+BAG+QXbpAFi
GPLPuy/Zp72kHLs//dTtVABzL5s1SU+Ji6mK7ZS0JghFPfeMhJdEUtXtPnDYN2sx
hyVrRCgFknaZTsvx03HLVVegwSWppYRwWknXJKaMly6xD3HBD/22L1Ivvhl8c7FB
24WLPVR/b+4LNJp3j+S0RSKCb07Je705cN4BVVknVnzr9dwJPmQvN4XAvB9C2Pzj
0VToZ/WYDiXIg5hh9Ge0gS4jGX35jSkQUlOkMYND7La1x9bOzbVVmknfG3gaTTuk
rLXjTmRzqR0yoTgUcYBUN8e28t5e5kszF7xeH3xk7RZ7ZSgvcCzFdENZJcgAobpY
9aJLuWHK6Nc81UZHYbj7rZ3ZMw1KxXnMEM+Dw+u12bhc9or4SLVRl42gpl9tZOSV
KTOQOMvckvRR6WH+S6C2ezAP4KESsNei9EPCLqhaCui9yKi/yPVocW+1kgwu6rNO
lCwFI+NShO2FQoM/L0tMxJXJF88TYDmyjnh6FA1ai+QZPAaogPX2fRGJe9cehsqR
w+L3i14dvFNrH/43C/c2BYtpzycMr+iysAjJRzzmZcm0oMCoLv1KXx0//GjEX9SH
jEp4uZHXNksq2xUkqIbY72ekgUnnWwOOjZFwgDCW7rUa+Nl6u62JEaIiP0Zy0f1w
Io8SVRrytrPWRwvCBqKbmBDqetU9wzK6FVRACgoNXAXwLRJwc2INZ04g23ZE12Re
zu4rFXFwjIdMiFvc5gHXuEX/xphg5sJXerGsAzqUpW6BnQTRydJg04xfS4ftmDPh
YIXWfq2NMZA3J1MRKf1/za1yzewM/Sf7LJo3T8ZVLHyQI4lkhEv1kRkNh43XGZcv
A1rRVi9gSYIXtwKzlyy33Q==
`protect END_PROTECTED
