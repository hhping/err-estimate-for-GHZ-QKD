`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UFD+X3pp48Dav5hdcGKMrqAum8g3ptOpdAiWDjHUYQ0bV2OGZ7Vxjo12cUBRoX0r
0Tlq80vlJxOXeCLsFV5nfIydto6IeoFbaeu96WrtjE7D8jUI8o945odNkS7FQRig
Jo8TQkoAia2tn+7orgs2M9vPvJC9Ve+JhjMOksmHEDtyVoFoGKZHp/VJWn0mxN5U
KnVhyvlfa0Y9FK4+yu3iGGzaYvZnouJlF7UJYIaHjZ0oIO3Q86A31FzwKk883EL/
nO/IPdm+waqS8/NhbJ/6LcJEjNqisxkv+du5sLU7HmJEAVkL4I4PTNviAyD/9KR7
Wz2bWJPGQsU48fg1guxZEy6hcWTfg/2Rsfv4GN1PyMbnOPCm/btRhOqqopGJt/Yu
DHDXvIDS81mSLTwQd8ravcO47+J8mYNEqqaOekGbbawnUnlAQqn1VC6jQeDASgBF
4b7jLe7HfI1LVFjMpVrZJkIb7pTugAowi6ADa8KQuE94xTd7jXCLlCfO3QrfloIb
uvdpcLqbSBdNuTMalMBp3VSJ9paitgfn05x7SceIK9+D1wGb9Y2NiC1YrvjU9FsK
CsKOIjPKnvatMRbcFbyTcFO2C5IZjBJ0qBuddRKWZUnAbmCAqG2PW99Y7T+UWi3e
P9BQPVNqF3etMkZTq3/OEg==
`protect END_PROTECTED
