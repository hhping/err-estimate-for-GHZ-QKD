`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
siiHPxJqdMypwIZW5A0LyAuxHTf9Ckao4wtZviiRU3F4VCmhwJYfANXShI7hdVic
yxgbKjReQ6yYYfhMbwgQWVgNXpC0GMuDnskWPlAnXkWdyKZsSOqHYovhBf/JnkpT
rfqYzogvGHRw2mf70jUjlv272FmKZ5wcCsXFFcVEVulA6JImgeV9Nh1lmBX9cFxS
FMGfa1kRBS10wpFl1rptBjb+3Z1z3dUrc8wLD71kcpAJbr6ncpv7Qrs9Es9P77HI
74G/z/HzxsPg84kh5Ks/EG/vlmBOloayOTGCJ778wn6BRvu/84clxnQ/iAJGX+gJ
D6Hqu1hFJgXwt4UERzfLQCozzd8kR/aIhjBUBLr/x9Z4ZVqXjutNeKe86Cr3NLCo
7u1Zy1JO4Z+NHj8lh0mIv5elnD3RK+OhNEjJURsC6kUBnbEpXD0zKajvJOi60dSd
MiOgO3C2rrP1WhP0Zr6ZYjgAaUklRs24J5f5cVsMNPblCzBmi2FEzg6868AvecfW
jazBzk7pBL9xDdPSZyS8zFs9fKeN1iiGxjcfTWiqckPeo/ihnY9N6SNLXpWQAhfb
7D8qbcx0D/0+hDGxJ7qvTPkXFxJIhaISg/HkhAhyyY9xS07kZSlIzIlb7bnUAitn
mzWScnnBi7bb80m1+2MF/wefXzu7WYGrXtJl1IYomlZC89BVaXMm2yqyUWr4pDDh
LglsoCxp4arZ+eRBSFdXSAi6HDf+dER/uHSId2aadqduQ5qEtvXMrbjHI5SWXe09
yelWp3T8DaZTzUZ0wVXtpz4jsPcLtmA9pvmCgQI542xfbrN5jTKAIHzvhfWfLczn
M7Wjx8IrhjWF+PEAMuCrR7sv8xVzJ8JkD8PZ4WZ0H9dO1KzkphxKDYbRmEcMNsgV
a8TG1iU1uLTrkIyBpagyNuYCQYwR2ETPHAsy5VJIXNZSz/3t8bq0aqO2Ro0eo6oa
shaql2Vs7mfiRbLrF04AcjtWDl8/marAelzG1/mjO2a96Bezdy7Zi6oIpYPDv5Qf
IOSFuIJq91FbW/0a4X9AwqjDXnLvAarHI0iifYxoTul8mw/gLx6f1iQ6SnIh7cJP
2SeQAaHcS93+jadnklDX/XtL6RGlUyqOo6oyXTsHKb61Fcur3TlkjpFhgow3gg5O
RvacqxkvNy1VBLyT1rT6PtkYh1++F7FYd2JRwVhicEoHgI0EJbH5vttuG/njRx3S
IAjntSr7iM5axUKSD832alhRjv78mUY3aTPZ8aKMhu68CBrJz7fb7/1nszmk/dXl
tpcl24JzwjobsdTbvyOMqBEZKwl1VKMECsv+3wbXKFW/fxbK2PS8QZl8unwI1mGx
53rSt0gfJvRIon+j3+8z0IAIWgJRW9FcRIXQxO0gOmx50UXeOlu8l+TFkq2G9Jpv
kUUVTTDhsUuxfsmuV9fA9W02byIFjUaJbyPZaPpv94mMcYv0YzExUonW4RK6wkEl
bQmGBwPI7o66EMXJJtAPynuj2vRCvM9AuB8YLc7yIaFjPA/tOPIoJjMD9QwpN6NE
rrXlsShK78kXcNRrhMoDDa/6DaJF50ZvWhqUgpANZ2cXUmBBS31gRgi2PHMU2Q5H
z7n1Xuy3z7Hmk+U9TLr4d1c9MZ1GtuhzGtDv1pRuxQsMm3NDWpoBlhkpoU1FlWU7
0p0pLcOzHuQoHuYue1Lh4A==
`protect END_PROTECTED
