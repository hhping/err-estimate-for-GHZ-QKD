`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eIYEcwnZ525PqzyZiW8Ft/FzErG3O1kb5geEj2FS6GrmHrsmp9/EEdBZyMbIci1M
eFw2hWqH4P3sgg/rvOnxVVYpALvqkdNeopRSb3zTc/gayTzslnRupRCAeocir4Q+
pKCtYA+ecS3CK8zuehlhOU1vOY5fGo8T18CwcSOAJwLcqO2UWqkslMxwNUVPecBT
sVck+Q0XCBH1BfOr6FRc45mxSiU6D0EJTFWNVlKdOml2iPEOr85Lp1OATkUxO8a2
4p1eGM8Xl9uoivpLE5s+/F2ybpvCjHKn7DVU5gXfjnBfZ9kmxn8B83XaIYxhUBjb
JPlFWTPfxZBAXHxKI7gi4+37N6v3S566ryBe4MBLFW+JaCpdP4LF8LSb6sj/XIFR
/hyaE0hv1iFSPegpgSNBWraYo7DdN7TSBemgaH56ByFOBEGgZe7VbyGWX8H8FYHV
ftNV9Pm6ztSBY4YiYHAEBvxHUBwcJbrunentWZhQbbQtmtqLAbO8rTyEr4pRh05X
nlzOswM/FY3rXrJXUA329lRwG2YDEs/NvBYFbGSgV5X8hNZZ7lhJat0CacmNB2YI
CZlPJoChhzJDY74Glk3YYgYrqqc7k/WTmADtXn281UdVvbmltUZgQbyWhocAaByv
G5tXgMcqqFmPLmAKEgVFpf+bo8JSnTYVCtjRMJnDL3YQoXN9Fl9LSLJUrEkkSMJD
8A0Il4jUc883Eme2zy1s7lcJunDl8GmuUO8oLjhc31Sn1LX2yrP+E4ki1Ki+4ZIE
1LiapmgqnxHh14m7U5maN8bOqZhci7KMFKRTkbv55z4+nlsiWESdlHa7S1e2GqTi
AbH6dXlIL83u2b3yqpBc3e1p5dHy4DsJTc+PJ51it0/+Aampt+ig736gd86wOcrM
o5ySk9FkVTPhwcciIPP1h3wIpbz6glXwSthHrYHbpjmLq247q2R5Ci+qg/V51ri4
7OvPsHQG10wq48DjhjVz2nQKzr2OXMN8V4b892r23WlhsjY1rKeBucD6+1Tw1Rkr
/qjxm1/uUuhysvwsxk/aiDY9jHS9viJvJlHhWHqQ8eqWSGofqix49vBtXWVUjVbV
QeegulC1Trr3v2Hr7jdGAyUYMG2naZ/mS4r01yFeUojxeLBrbNTktoU38jHHtrNW
iSjDjYVyTvaJXZXjRAQP72w9oqEcW5VbsUaLw33vk6v80sUfNhZ7jMQJtmtrA3Av
K1/9NZd4dEWRvzthHBLnhH6ndTE7AoZI4aLXoljGVXDml77kea9IyGyM5BJREhdo
`protect END_PROTECTED
