`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v54O1HOrwkj/IYl8xQEWaqvpgpveuTnGtLeoH/K19Gku3wVMLAF2p50Rc6R1sEad
IrZ9rbIISBheau0nNNdfRgdB5LvwjjP9rF25sZt6M9hu6PRkfhJACwATFxcrw+vO
gBTqoetIk3ZqLH613Y0QGHSV6rKACZ/0/Fz2+0k1OgWpxJ0PvkQtIRNhw0w1btBr
HLB/rO55FhFpOse/Tz4FVAMyBRbzruCPPTuvdOaTplo/SnshW6uwBJzAhXC82gEv
Qx4xakhryx2FDmPHOKHka1OJtVl3iDrp/E7QPWSIVNu3yFLWwWDmo/JVteFO2AUr
kFtIDN8egYdXhoPPLO3KCtRtZuIvgH8+x+mO6CB0Jmv4Dy9h1qMM4xZP3aAJYLzd
wnt/tc2XoETL4Eu1eawBAM/t2oVITbqDvjhHZGUfMV5gAQKiD+d4EKyuOLBsVzUh
x8DWAY7vCrVpuGSt97HEqL0ECAR/M9p5JVbdXcK15M4CdGUvMoh8lUBuLX8h0rbZ
AZ4TAMGC1tiG9zeDzoUgl+HlTWEbxG+cRlA22ktBXNLumC2OUTcF48d+ptLzLt2g
St2A9UorWnvVviou2tsdVHY8YxJCGPbkpDoYUiQunKSvY429cSm0D1FsIV5a6qqq
CmJmv+dM9/5iarQoni5aPk85AJGd/dytmjBVoYs37Fa6+ec6nZ7ZZ0j/DwY3pQM0
rpduPOaXJU0dIBR+Ma7nFdkbtv48FE0fY7MCAaqXHmxU2Y39S8vKi64U/cfYWigy
SwCAnL3gmnTOcb/ebNhzaXMmBjJWeTIVMhg/IscA8ctC/iKH9627nOcpD3gdMe1k
Cq0DKjOyqVwL8jKJ2uBGUhuXnc1enCGuh5ybV2uDM2C4rHnFNL48zIuUpv/WTVnI
kF3ANQSBK/Nc+q5zh75SoUC4G0sALpKnDdIjR7/tuLtg4fq1mOJNtOVyYh/4mF4+
tzSqv39WZSk5Ve7tncvH8G9sW14s4HvdxamdSFPqb6hQA9bVeXo0Ta9V3Ts8Mpip
1pFLPIWsgcA8INR3u3MwcxujfUds54kEbpKfFy7SWNvikHYaMDZSWxe8K4M5tHHo
lUyZ/5CtwWAqhFaSMcGxn/A5Y+9MztyozI/xPiP13An89xlgGiTqVEObFRdQ7mT1
BU1dntIN2oR6/ZphyrbcbNCwyWeOwoXj0LUi1XZZShafKJB/Ho/GfnI8lp+2oXV9
5/Q8In06zgfJhG0RpPEAm4JjNqv/rmZ2k5dpmghTFgX+aYdMBHsHa4a/JaLUutUh
yvgFdk5QOysoYcb5pg3fjFNYDF+Z3WIG3rVTyPtGFKaAkEpopgxy3uWe3UI5rcW9
oTbVQV78iZA2bs8cXg5zRovkuUXgggMod2RpYl6zAyl1wZ0yd2VsMygVw9GjJ8qo
mQzAKrJ54MmbAPLdbua9rQbJ8q6NFFfNc1Bqs2ZcZ0k4pZYZUq/o4fINvt5bGDpz
Tb39ufby5fYxAJin80IlmaQ3TERdaXS2bUlOkiUsmgOTKX5zRsreI03m+zj5J5ju
caxXJYouoUrGq226/RlLpAEyU0s+hG0n09o7fwQI4cCXXBhXTHXFiXpohSkvAGmr
60hv5UW+6GRYkdQq4/jPYC9uKkg5/Zl19XT/UDhQlC65rJD+oUzvqRXwl34DIDKI
rIOJ027duhRzT38HSG8mqzcU69nfrFTMXywJDeu1wVcvLyf1YTem2iXNNmPRIer9
TBTaSPbwdajnhH2/O+atxTRzqpIoBAm/Ue/cIC1IsM0+BfPhoAeoGrhJfyJzWKN6
Z64VSY/YbGIphYK1eTd2b7exLD18eYkYojqZHx0s5VJUGaUj188RYTWuU9sWh7uY
/VuQuOJdyHPRCKmbEfWfWFPKv6YLNs/AjxJ2npJFCW1Wm15vrgwwufrv5JGEiDRN
mb38PZGYCvk6moX807dXeDf5chI7xbWluUY6v8Kaz8s1l1Zrdf5PZf2c2dbFQII9
jdsfTqapfI7apR8KCvUXWb/N0sVCasAsBxNr3Juk3Y/1NDUPvXxmrHBT0AV3uSEa
`protect END_PROTECTED
