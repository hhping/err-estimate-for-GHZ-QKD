`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xi2U2/pZAyRUKeSaCKohdBofKnrCzAAn3YKQwYDarcmm3POdnYBrcPIoEwC8MZ/g
0VjcZGBkJoO8Jo2UV6kyVr6GsZZTUpxakXDCAb4NR4uSPTwqrXfWFf9r0gLG6adW
sc2Y06TXkZHDXfdr3tyelYFE+FrmPUEGZZi/C2QfsIDAbz4ni82//PlPulnazul5
w97NoSj+TSe4YOIdc8G6ZnZYYe61SY+MgrI/MeVQxkYPGI6G0ivRWzkNmp/0rA5L
w9miSD/uIwHD6cgrkd3k542e6GVYN90JMP0HoHB+FdmCqP93M5njaJwAqvs00hgw
36xEor/L0xdU1VBwhtEjLEhMboFcSuQAwH7Q53ZH8cQirwiE5unBX/nEvAuo5pm2
MOt8oFeYQskqJL6sFjeTjFcobIz0/FsvgaUMt6TfMj5MTYgtS+vuCyqvRafO/bcZ
+xrIhBPMyTsFtPYEHh7BaqnZEPAMkdAelO6/K7i+8BfHMS9tE3ragta0m3SOG3oi
/11XRzpcIXJuNIEaCKxeBbpV5HvFmfo/8WjcHoLOmVTa/HbZYYobi3AjH8UPXTa/
hI5eV37xcSfO5tl0dQ/18O3ufaa7gPWC8ZXd4izjD9KjlOUwi094C2NCvZvnsmFB
N5+O7xunTieeWQQL6QWo+/TOoy3R58Myuzui6x3Jo+vgRdbNZXe0jp7yRgPxI9rB
x7L1+h47pxmOvZQdsu06xt4NkaUSwBVfJLXGw2T3xn7ES+0+MF01FEwErDKYVv2M
hiG688x6ZrDOoxx1mqch7jUDsIociw3R3TXbLCYMiZo6R48fxxST2CzAKR6xkJa2
jOpW5TpS1lwNtds3pWR8/nXg3UrF2E8iiDwaxQqWI8JEYrw139nOlE8YnfJ/XKSs
RBOTSZe510s8W+aYgzNr+pO1GbIVCFZcpRHWd6xmVaojyC7lebZCpRSKFnWPpZJx
DfvnbNMAcxYNHr5TOIvju5uqepAP5/Jvh1If7CYo2UVqNZQAiS2LF8cmlIL1A3Yy
2JuvzVr/BvqLMQdnNbNv0VcmF42YEILmqxEh5n5890mpm2fSKqdgYUhAhqDaMqdl
yXPYc9SViMBgkAWDUPbQmDXWjBf/VYoCfw2+LCmfnvwdREFDJzD/Qy7Nj8otp5Y8
pm/+g0f3g316r5/sWiuRN1MGHKzyVrNpeDieN+1YXYfB3TVH8C5eLggfxfPEFkvY
gebyoYrERxKb9qfSWXbE3udKRIePN0zdUBmwGXfNLc+JRBz4PvKb1HPuOFcnmdv7
EBoL1rGeAY225KfVY/l2UAvnuVd3uacjFEVegCjFkELgq+qBxa6PXFwNJmdzB2F/
mFdbzNSL6lPeSZAmK7H4WHwB7YEYuP/1/b8ikA1nQV0HtTQ1gtMhiypjcLSnJJcN
mnig50CroVKMkKeG+AtkHtRGj8oDaze4JCbvEJLJPJV1pIAk1Xob70AmJhuTZSwB
yyNaSI05AnMh0L7/civvOKmG+ygWmmCxxrbLnf+DBNq/qgfM/vVbBpYzcBGB2aHB
okDWO6pIgUtHNMnxvWiywFraSSZFurLJSrFGoo4UMc3RkuXq3m1re3fvkzWn/v7v
W0qYsMFDOgGbtdbWObvlFyDVf1TSorwXTK4xUYfjSdXtlw/Bti/0anOz3CQWysHs
wPoxbll2qLk9tfmwcrIw0bhUgaGx1ICVxoRo0fp88PMnRCeZJVjtXZUBRYlbYIKG
psfYYlSH+xcSTGcUn0DPxZAJfFYbBXDQnPYajz3Bzl7M2sDFbYDzGNshy8p6dqEW
9C1PD6sa/+9GonWMh6NavAK3V9JWuqShiMncz5VNjy++GvmC6+2f59SjMkehoIu7
lC1HadTeJ3ROCjyt0ZkVVcHGCqRyIF/4VdY36NuVu/enMQpaHgSf6UX3yntk6Xfw
UK2r7MXY5c0bymf6s4s8NH0+jsQo6AypheA4U8y/V9Bwg352sd1GeZThGtcduOgX
eiMfdWJrckoc+1ZIr70g6yUXKgahByglVJaq/p02Rh8Ucexfmj7izP3THWvm1iPm
u/5OTjDHchCfPqMKqI2IRb788zs5R9CODP0cJVRoOHSP1EbN4MI8w1MsTPS0cMuv
O35dHunGNjjdthRKFEYeMt1uK4ymusRthulkPJ66z/How6uofmP77CqLUCUEPL12
25jbmB1U8+t6G3xPVZIayi9sa7Ba94wt26FP5BeCzxJ1aKA9kZZ0v61rplKR7V2r
piSyatHrdMq9wfEN7P/WHR7PzzL6jAbJxPkRobYR5gE+hhjGLaQTkmInTVJUOQ1A
YEpfNeDwATPedzEw8bn+BbZwlq0P4jiRa8UAaZRzjzo5NhGOWXtzXgvIeA8mMKs+
YBM47JIEQEwL6zd5rJXDTE1DTzMfMHPBB6g7MYGrsk/ZSsZH4a+ZfWRI8wxPmqAg
R6etLzwCZIANLCV0jvZ9YOhNrSYUPNf4WMYsanwgaes=
`protect END_PROTECTED
