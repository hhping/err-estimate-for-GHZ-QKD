`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8BjsMrKJNLVqxZeb1FKfqOX8zWJ0x9FK0UT0QFM7nVNN+I0YvpHxlLkbACsF6iee
q5BZpSMS14d2iPxcvVC0yrAjHXT6Neht/S3dv5cKDxhEG9Z3voBoSs2lvUqMPc+0
aNYiC1mr5KgDU5lf7tuAGXA2eb2vVhruEpjG/2FO7d7QCwsL791yvZf47FcJi8FZ
fNnB4f5nprqHC/KICk7W1/a7vHiq8h0f5exjW4e3QwhXlWFf6ucfdmfF0p3Dz/rX
W9nga9HiiqCT1XPtrbWR/rP7U+xHgx+V2duNSFEwY9bQM9R64aboQgZkApZlu076
hrVnb4WZ4yFu7XoA/GtyqaEB8YqtDJALxbDJ2WvS7uzIsNruzWzbrijAQIneUuov
s46qqjv48Xv0PQFdO0xHWYwr94u2YyY/e8tMvII0E9PZ/pwHQtSsbXYs22pbdzSF
s5CEjsI5vDzKmRf82D9xnZtzCKyJUo/mPscx82gJ6zqBODzd+C9x0NhT9ErYdUPh
gZFznm42PgdP/8aNMeKSEuBfLUiz7ybQ8W5ZOt77DpbdhGZGuysa6ZF86BLdcJlw
wD2QzFyKW5N6RuviiF5IkrQoaYwpRy0GfkReExu8lCvpmEP22PrfHcjwqfY3xBYx
vdAJUuIwLxLzbB/ZuwiaWStYM5AdXyaEevsuy+b9e0uzPN1udpnyXM57kO9WXxrK
OXt+3YZ43OOu1liyXP7pi2jfTvmcPC7WcQpvfU5ihZY=
`protect END_PROTECTED
