`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j06szFyaqGWAy37MtCrdvZN7VozjfKg6MhSzcBL4Vo4OGGNPvn0W3aT0Sih3DgRc
v3XPs9731fVNIWddk/pBb9Ju1ZLDORFq3O+AHPy7djcKdgGwSNqQ+GWiy9lJPMb5
fYFCvSRGxuOkRu0AanzWDRb4RRtJa558mg9tLuhb/f8Q64Cr/8tI/4Xr4gk44/jC
bFSEnDr7qBDU1WeWAKuSuikKpklrQiDx0K67l1m+VE4809jwhG6kBE4+ZNYIvnnU
eJdhaaRt7IdSDNvG7nUiBWF/QfOBq8p1Oh2RRL3fj+kGuS6tbwKzscl6L/gWmqTd
iGRLpc/b4G9ezZYTb16zXGDArGQ3BVOJjEqlLz/9+2gnv+r0qkgHJxL2TbDVUQYU
uZYKswYjaxghNAHIE7aZcbmOCImCt7w7eaK+bYX2j3YqK5B34c70pvQKIb08+ww3
kzxxYyRsvD3/Gpyz8gbyfoH/bpi5qC1zLiGfYIFhxQAVJ/hYRRiNixZyMSM6j0OQ
TjVMjFk3Nap1PlzcOj87lpsvShSJI/qiVi3oZOaYZvwTFbtPXyeK+mLG8rCZino6
x5sQn6pTSnu9pH/BPLHcr8n+WLt48+Gc+2V8SRU9Hz2aAnjDESkUmCxoQsoQUf3X
H9Q9LPWdA7KIW0/eHxk0jbmrTQfI6NmoudJwuWpRd1Ej5dBTWwsKX+Izmf6Z4eBO
rsuT3LL/kKAgSdS8ku47sHrxwEIfywm3aURm0xIfIXo9byNoWtXkRktxBQlo3bdC
8ajTXvMzRGx/qSmd1wbcY3M59MQeZdB1A7wBBNf6AUWuCRQIbeBj8IVL7rR9awDs
nFVljJ6Iox2RvEMnH2gR6OI3lSjtvbCSkDfR5dZeFw1MVnr1nx3q4pFB/8Ab6cvK
cdw90NPb5HUK8dNrmon1XjYsM/XpBAml6kDryepb46G+F8f0zvueZrOifuXI80G+
DWewi3nwVJqTwVNQe+2yDD2fQbXKcy1wzmsyn+CsmpGD3R5bFhwNN3QHqFNid72V
aaDnndS9eISkbTg2YNipFA3tt88I4uL+SB5NG+BhHFA9fCWV3aQMbBInpPCSX4h3
vW+760umapchTXPYYflLJitugJ8FjtUHZdtFde+Uh+2Wcf2dOB7WXlNuRUqxz5iW
IpJm6hnjE/zorKDWcHptdNvgqaVMHCcnU8Z0Jt+IxnfWAXjq5FWTkrSrOsbXTGpR
6JcBysMR4Mj2lCur3x/luEIeWdX+2HR/YNAdA7owu8URT3gPpBUe2Ok/CnoBKNUm
PEiIF4W130/XbXRWFCwgrGvzJmLb2m0+H/nNuLmeNSePJXuSj+avgAc1yD1TuE10
f6TISlqk6yxMpUaI2y16xKDmHSkFx2qnoFIwetSXRlio5HN/Sw6BIYvv92Gp2w8S
2cbNaCb0bzfbyBJi23TVsYa3TPb/ef+x9nwTPTA2J0H4dLd7JugVDQOwNztwFdks
FnMjxpx25WojFopJW1aqTaOosP2sywlqr8hZfjJWJqLtlax/sHleiTb4eZgqKuZg
crOW8B1ouo80R1x8UGWYg1daGPZORtkWOITskNgDXnbHa7fGQu7JHMKVLW+KVg+I
HRgbKPLGQHvFWX2R+hSPRv0ezFvl0JdXkLmkKtDWEYU1CORhHCtZ1/zwwXeLxNUc
`protect END_PROTECTED
