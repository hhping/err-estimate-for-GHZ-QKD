`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dr0bcWLoSFEnQr0bVTqgHhW/q5dfNTFM996NoLxUuHBnhAJ2QyYWYV/o9bO0UJaI
NiWIIiFrFgdK3tsnr/IsodNs/5JQ4eNedSArNXHUZsx7HsAIFZRitIJsBdr11w9b
JLz9+Nx0Orjbt/uodRQl+E/kjIC3Knqr0wG3o7qEe49+1wIDrYTko7lzE8vdo2Rm
58Er0cGn/ZVvwrgC9F6WIfoafgbRcYPRMsjOsYItXSg3Bf61s3awFqJvuVlKzUF6
X3oa6H1/H4dgLN8W2EtT57jaIgSMwzazQ2koUnzf/DRgOaMYT1LuBgJojHKuwcsp
XfoKRNxx46EZ6XZDFpmnWVrrpbg6rp5s18lmUIFGSn5yDhDK0JlLVdc5prLhtRxX
4HPcHjJpeM4ZIB7lIBdovvC5sQm83ZRCNUVD45ity9hAWCGEahXWvWQgyAO7X96v
lA9sD/wlCzNvHqQ4jPa0yVngTIwmiyN7Iw6fOSKm3QU9xvzZv+7+B9QMrSNLnb/L
slf6PExP5qnYlKn5ExnmE2b+n77KsryfJO5Yh7RO56g2q4+ZfejpFUkh4shp+bpM
xW+3lKrXo9niC0RogH02J9JcO8+YX8TFlM/KueMZEw1yz1K1bQbEYXhh1b6Joqdp
96wBxZgDvnCFAUXmnJuNkPPIHLlirNaF4oNWp5IFUlkrnFrf9CX3kz0oMyIsvp2C
ayq+dij7C0tlIeULxRkU+2N2kFzgE2WQPwcKGVMsbX0C1DeLI9heilA3sMPKVZUR
ajgBlNDXxkEIup/dtf+48R3vFqiGPSMTGgWEQoBxtEBZulgV7CWjKbdeJOEKg4RT
tmfBRs/O3wsf3QYq8vpRQLz6VRUGb3423kv63E00boZIahMQLx6q2GnGVm0WXkqU
cyChc3RP2D+LEq2vRFLWSpgIB8jiyZrup2kC54ZQMdu49CssTnNaFogsEbRVuKkt
P7ptB/z74icVWm+wmpOQ+a5zEdcYu0+DqefgOY6wd22eCtjVJozzs6lV+lulMMKW
Q0O2lxEzG4WUOsMWLX4xSPQdUvhs68PNvk8uSYphaxjoprGRgyIDKrl7Eer54T1N
VD+DRjJEb0aqqSQLVPpaSGpITvpTZTiVSKkR60XiWDxMBGVxla7i20a7b/zUUBut
5fMjl8QPTAl+QPaLIOHWaxrNDS2H5HIa8ZOakoSk3LjuFdr6Ze8ZXkoMhSQKbpOj
2QOxg2TtN06RO8IHF1OJ4/7UCzLKYn3RkvpFeVwXtc5OjCCwZys63jfsMSG6LyYQ
ZpJByhkkCr18kGBXHk17b3GQ4bIdTaO39rKSasHOdiRfzrYcqQ4JqAMORX2fbTXN
S6wi+/o7GmGzdbQbs0Ng2MfSSnVLQKARgI/5T1P+uSjL5m/wt8YU/Ky0kYKU2tQ0
0j5TV5tUGPqVl8/s5M4kOaLsqNDdScefgGiMpmXnFuOiXWziy6ZY8RMkxwZQPT+K
c/h4LL9UMh90tPCXsjVXzqYD2QxQTxjsTHVsdKq0GluakB1Civ3JK27pZe+5nxxi
ffDvdIlIrcVSyjbLPZVqhSBcoDN6fuc4q/Yq44lHb9UCCw73/GDGv+Mjcx/KopZo
x3eoibfgFBBhDKhY4owqqOF6BluGs7of6LsOCqG1iV52Zzmih4cUHzpK0A6W12zU
yqRvAiQAwORCZkymKrJB6Tl69prO33RG5zGeh077IYiz+CSXC4dm9ON/sHzoEDF3
flepzQqgGkgKHLw81fyXbionyP73E2gA5mDTJu5ql4PvLn1rkJPXvo0uHf35C9dB
xJkzWz8sND/b6XkXvSqDLRYKsheVgQk8cI/G3+mWVMslsmv/VuoXwjwdVjt7o6z8
M+PTcldF+7GTZFhH6nUkTIuPREVBgbdX1sEr4d+v24MAZMI6vI8Xx8ZC6JeBeSEa
46XGyvjlIKjl/cAkuQ2oXs1f/1TIicwI4bGzIDcxwMBtyexZa7rtDbDiqbIYft8M
wJjMVzYXx7o8Cxix/iG8rzIPQqj6D9ZO18/PpYFGHFA74mqJhJFrpjSkhshlDLWy
z60H+NB47iINuWpu3EZCH2fdpEkXoghrTghrYz2QlofdnI78Y3ulBvQRL0+FOyuf
812JY+NIWS72xJLZRpTJOifXn13sqdTxEE3M1oIYPlkLkimlq73hM4sUBOyQHTRv
IwsgoW6j7nMyxtcLMRcMoG2LfRcg7WJqnxaMXBVYhONgy9Fjr6PkOVetvIBPng2a
pRVNdigMLZ7UjElO14L/dA==
`protect END_PROTECTED
