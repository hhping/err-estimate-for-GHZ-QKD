`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2LhBJs9p4h5n5Y+LLXpuoB+0/iiMZqI+6HfZSPKMPm97n8ZFRSq+8ai6TMfFuNh8
o+p09p91mOsc97jL3ztM8lXxmuPtPZ/WlGpq1MMx2K9nLrT0tzdW9oa2oX3OaoIL
Vyh4fZmJ0DLSnlVxkUc/lH1jucSkj88PoHm1szgufHOKD2H4XMZRIQfUIw/islb4
utGExlXCVrl5NaEArHebM+YD9GSiDFVspvv94sqby7drgyXyeJa1BEE5hFzX8hNE
IVvBvc+ud7NHMHZ3+4XzXQDNO1Z9ohlLdpOotexSzZQpdvTB0+wx79myDTb1+B65
0PIR9vSih6xUWIIB9sthmpw2yU6+lwG5pPzw7ToWyuNr6PfcqFlxDSVMfP6RWArm
5uc09gNXIDusFnXli3dZVErlY6XGv8LevoIiwWkfk+irR1/tgzcLHFQD9WlNBzi9
ObUoiDny75GcSEbydbt3R30Sm+jy8qW0QMiujGhKkHPqPREm/xrfwnSfPCxWuk1c
F6aWR50WyxlgiFeST4VeEnrnttnpZsRgThSj7wmsmFyb/V2zxf0gBGNZnpuKhclV
`protect END_PROTECTED
