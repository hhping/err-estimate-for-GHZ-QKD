`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+f3/TJ2MR9NF8prO3LHGY/rVk+2qSMUuLhXi7Zwvefex6AqYu+7jXjy/WZeDOx2H
JbIrmewZ8SAIqI2jx/VbZEpABDC/R5ZlLZD4u+nhUYONo5/BqMxhY1N3+w4gFhlq
MrAtxkw8ASpJLyoOBem1v1HexexMf3WDDfsV7Fqjs+HXPVGJBrpuDpvGaNrObM+H
i1YMKzqeP7OY396jOa9yAeI3gP3MoIEtyCJKrwKZ7bv4YoE3kdaRljru8wRVHqWu
rDBN54M1J0jZU2cuuXtEuO+aWVdG6CHuHjfJ4E7vTIXuvHUGjvF/h1qjCmhVCbKF
YFjYwRXa5kMxFMF0fGh/nNNlB2a4ZqvivJNvLs7eJ97+y5XEaCAydRqqQH3m9bqE
G84suUkmP+xWzHJbeUCReg0KJ6Gjqtvdh293SleHslnB4wkee265BojL5fL/jelL
MaT1ldmuIpBEifDgnialArDFUL6A65QIJwkWFqHN9TQhdc1ZN2G2EixY6LKFuO0h
xMu/83hxmLKLJvEcgV8SgzP54R8CF5RtGhBWE8HqHR9AQoibft6B0d/1BQc32HhZ
d3r5bR11Fha+MTysrSKq8qeZJEJ3lGmnjQU607Mb6UnpxQKtAtUhh5NIkejlHrEn
DarBzZbofow7ZIllgogmnmoZHABYN4W5Jb1uMRIpKVzQB0jdmF3coE0U/SSB4MA5
rv2FUkC8yYjupPPAZPHqecw/arPUsr6GmYnruE4QKKi7GU1tG02FpwKHvQAdw0L3
PbqJvm1UtNeKJVudlWCJwDAkHCLRwUwnCPTfeJ4kTxDf/HqkjaQWsWuD/FAkv93F
CsNxvVkiT605VYv9JnOKLGL3L6v79+BbXbqsJ2xwpdYMCqLgIR/yTShHkZ7IAdYT
g+3WvFJTrC/lcwq+K1EtfORXTNTv9nFD0Syz3QBb4PkRqOaVlk1NStckx3QNx13P
dhN0usCEnbX0IsblFok+Xdo4yg28jeoEp4baDiw/JYt/Mx7s5kCNeITiTt/WSpEU
seS9M7t6cj3XFY8oBblGgAZ9b13Bxl+pZxij4MS4IaWAzbn1KZpfXod0Y0VP210C
RUmtmOYdOStpysInTalLCqzcNobdxNEEwfkwhgKoLvMs/BUvJyY5fot/pExYSmYQ
YgQAhLM+7C8yLeedin6SCwvkplFBGznseWOLW30Gi5ecZFet4vodSlAik26+6Duh
mDkU1r0p56IvKRA/FMtS5ruwAifZXpLJopWkwdaW2T5wCXEmhu/HUw9m420+ZO+m
zc616msyDQTskV/Oo1Ua3X39RWVxbPyxuoCcUpiLUCJ/5tuzgEGaHxQby6c1Q1Ju
Ei5OGTHeTkB8yFVjozDaJ9A0uVNRWvAxnN8y2TolQeWYTXsXu7fFuNfL+Xfd6wKr
6FSHMIsm7yq17F5vkJsDkXgj1ePo7rNP3sxSXz5K1jYDLsO7LY+j3YWQxJOlFoPm
ng+ShxWanni/C/W7ntFB9p4meXl/EmcELnQSDPNAca5IKB8nEblCNjvHB+suHvxM
mXiwK0XvVx6g92o9amNu8viBoIebK7Hiz0J7an1VzRy06B9Okjyya8d8Vb18kHs9
3rlA9qcLb6HeSV67pmj7G3csYBhWLh0lYXSZQGSQrQsrmLy2NKHSVurQtL6Vkqe6
UDZgEV0HyakBJIosFYRedW4imX/jaik5ByVx88aAhoZHoU4th0XX97UByqHFnqVN
AkIkpcgW/ZVsmmRxlQFMm982dXuCz32kihW4wdJV+mZ8fL7zl75O5WqTpMNw9Yce
vmjaWgwZSt4pwBvtZTESiCPDU9MvGgcpmKSml7aK83UTdGvB41d/WPqW9IHlYNma
vlZqDwfXxdT9ansZXZsGU5cY0kjazc4zO8Rs8xv6bZ0gvOSpk/Y1TiYvSoOrTEbc
aYjfMuKmSpdPlGYze9O5xpdpeCmmtMW2Hd/Akl/zs8PokAtEU1d344ITTPB9N+Yw
v8jZN1gTTI0B300G2zw8tj582byLB1Xpn+kI3BPU4HY5sZpkMMHMvWVjihEap48g
6pLZvzZlt39Nbn36pp9wW3rWpR21bi2bzFXqpEZkBDleOR488fI/XtKMlgkhBfj9
CJ+R/aP+cLp8rf9gUDeXAJ8Gg7mETHxWdv8e0I673q0+S3aO6ZFZsBvQkhk0jxuf
FT/9b97bxbs0h26lhVMn6QqV4j/MbM+rBiYuFyC05TJG1odkq//gey1zRBLX3c4Z
QR0kuTjO59iK+66lmW3IZdueKEFESBn/KDHSoJdVdxq+8wcYqjkNOCH4aJEYn1xd
J8wpO0jp4voP57FZMuv35TYapWV8xk+zklAH214KV5h9wf8hA0NJoFupUASIBrJT
sJe4qEkb7S/88a+27an2q/XF+JENufCCwJByZhO2dbU/vYf0dqSoSrYAX93X6VdM
D2O7T+wIFkOlTzOpRz4ONZ6817QtWPK3GP6xWgy5U+ro3GF8kOQkplDVRoiDG1+s
cOQONX8ivMpa4OzVJPXcgV18APgZHiI6Jaf1hepxiqumIxhxqHPN6bpPMRaSpKlS
E8YmLdzL+53GU2soA6BPmlOdgnufXgJkHqppgT0P7KKBeiPTRaAz/zRk0wREMWRt
SxvJmYVM/+4m5RcCuJ+hgIeHp2lGyuUlL98zvPYo3HP7VUzYVsJ6judsjnHGssF+
XQWzu7lw+FcmiKLfNIGWAFDjZ8+N7FcX977kM+t26g/IFwTDONicu06kU+oP6QV1
yEhv6iC5+FtYrNPSDJdrCrErb121oPnYtuncrPe0Gatxt8n/E2ifOJa4N78vkd30
B11VKxGhP4l2gRN92+LNcOjrM2Kenvphb2G46G5PPpdxD5pt9pfTKgdWpNHgVoEW
N6IDhEAkI6SOT1zDnM/cfLuzYbzJVFNeduqIhadi8lUEgmloDnYro05Zl3Ucszbq
HiI+UyCccpSsEJkdTMjjNc+gWzQNL8dJ9TiT9dLy7hy5pOlJnBKqnlGO8pZBJsy5
cCDdz71uVvZuUhpx/x6zX7zw1xkvZTCY02WMsyivb+BgVRI7+tvfAyqUqi3Yq5iZ
Fsqb8PAvu4IJTQRj5GhFZD0Jf2sAGc4gVH3C8KbGXJaYommZq5JdjrMWTuDhj77j
rRMWl3rEv4PhU7Mdt14NQBD7Y2jZHSSPXYWzfGQRTEPdgJyXQIsHCa7tzG4WdZUU
Cdfl4vYQHLdJIAkcKg8eFM64w9IxuSbqOlkpQIbg1gg4jj2dEbqKsrN0BsU2ZqaN
8do6a44sRsE8CbMMabhQ3ZynS6xEqJf5l15rEzpLAwNiw6oU18eYw5bKSYBYFckE
2vXRgXmUIJr9Y+0kXo3TaNNGOP1VfQOQXozIbCkHxkL5j/1zryK/LNXx/mHfQQzA
ZnTst3il+EwwhFcuYnOs/QXM+9FpucJwwGXRjVDoWvtfbN3TBv+1yVjYqDNqoutu
JMamcBvNFtC4ke3Ke6rYY+sDE87arF/ulTOpffD4pPOeSbrNFa6YZP0GelUozZXA
HV7Z8nruB27b3vBXQ6ebHFoEjQ++h3yUPzWUvWIrt769Ogvgnoi2d6Yg/bPIkPru
P8iMCpaw08mpwx5s6M0OEhiQQO6nIb3rCuzyTBp6NYh7LreDWwhSvGusf2ZMUd/g
wzkfR9CjRm88UjvV6R8euK34yQiYmElQAWI1uw40s9Vms8Ffs4o+Kwptua2GaGzs
vviXmI8+hbXQa7wWcY0vF1KWgXdPR8dIsExX7LoeL8wdjIjc7xJF9TUIB4+te0z8
clePuYOXQcmISUJ4EHRLr8NLU/7dw+aYKE6SC7oXGCTbmjzFWytMQIJ6Po7zNUzQ
wEKfqcgeAUVhP2a4ACxTuKvqsIH6cGW0Wklak/XaPYZQlIebFTA3rLFcUctWKAEL
3TTNfbIcvbnNakLCU8oRkAHCTx0J8G0g/+YxHw+I1iuWG/vqa06aKIGvsvSrJfHw
95RxzokWExWk736QLLNXndU3pL68S6hn4c/+HV95ftCMRZ2KebyZqBUYJSImAOtU
Qy0ds/duI4OpqqeMNR/GYk9WRURZNtQZDNuqM9Msq14hQ/IwcEOb/vXgCNCxqfhU
l2fuuApeasHenna9wZ/yihLokdcfXep1n/+doyb/0dDzBvrOclC/ZsAw5cKxgfeS
LHJ9WIhAlJSxkT4KywAnC/URNTnZxmeaM2fYwwHnVqzErmHTNa78zy65zHceyzii
uHpLi58Hl3DCWHWrZRq8jiYguNHjfKjjxa9ezWcjhv86RYdGinnR2or1CKmlfhjq
/Nga3F9i6+EBWw0JNtZhSIX3mpgGtxjYmgGrQuP7S3qeRLw6qaFcS7xbmEI850n3
KLJ9hcInJpLdEfwBKPfsSdWS1/Qz8IBUPBJdy1xRVn2GLMkEplpJ8J+8o8WDIcJA
pwJZ65fl7QCq8n3UNZm3mci2XLObL7Pnk9zGtI7mJ8HTy4cjv3ChG+pox+0x3lSH
5OSPUH0Yar2VOru1c7cjK6hfxRx2URiWSA76A4ywzSrrU5sp9WNFMvK/Joai2FXa
ZeUYgWP899JZ95NTEuCjfTtA3nMJh6i9+S7u93lGk0XCdBITkk3DLqg/WuJCz0Qb
3zFbUJi7R8n0ij+SBhjpq5iq/NOWY096UeO7pMBMa7mvNvl3oeLweYw5gn09qa4z
w3l3wPQwy2szuJvVvaEFFkdUsqeDPdumXOQg5qeo8lspb9oIOrS48Yv2NoFG6lbQ
FABRXR3XkgxDAXT/L35xMjRk4InSP+KMB8b9GirfaaRiq2wbO6H2yaFGr3UssUr5
+c3oyOYRT6Lmz/4tpfO6Lwpab2qsvMc1dBin8Xh3KFp14b+mxkwKvMZtXfz8Dt11
vVPKiW/qDpEeiJGGXeau0FK3Lgg2O5MIxzDGzSJcb29mIAzcdQy/cnRIn1iRmHFq
YQweUee73pky7ZAegZP5HcuJWC3I2uNu6VnlZLZx/OH+1rt0u7Qq3NCYk17/uudp
wUC5oa/fO8kwmdQMwpDBu2TJSdldgSxJU+Bv4HaaoBknsUCI/PH7R+rFKgosBwl/
hu7VtycBxfgqzvkgjx/rw2SPBFxHjoSbSoHSa4KucxqqVY/SbZf606ser5VsvKgc
M0zKsobLlrZfE6KCy8ErBDzEbMxjTMbo8aacEx/YQazkPREgx/5GixAzVPZsfJX5
VltxrOr+hBZuoFlc+DWkYIad9IlSWhQanmEpgtKRFmpdTH2HPLKx+RbuEHs+7dfr
YOb7L5xkXiFDK8zy7CgcSQr2KPoRsMvbg1YyNmY/FAJciDgQxZQ7wQIQeS2V9gIW
YVWN2H4iMc+SLD0djKpe9k34YnaFKFTnEUmKazSLUD8fwZ2wYXd1tWKY81N53tZY
6oEfsZKHhZt+cTlweOWL1w9xEwcWhcRpVqfvVblDdG9xdLwlwJYSnXlUCHPPMWD4
wLDbpatS3XnEh9s/0o+bDSg2lrChqmPrK4OoKdUllVDpcmAzPEn3TGzEiGGcRB+6
seGXdV7dVVTmMBwItPCnily9pxTw8uw/ncfWlb970ta+SgVemrmp0iXQQGG5Wuxl
8V5ZuK3VlPoPq52E0YLYw9gjVqCTJALcpWqmAVZRnBq9ZGCa4qrKDeOjgX4cLDfT
oITALYz+8QvhE3f5/tzxiTGCAcmVWzgK1n99rPQK5wqdSoOMkUxPIeWyFSrb5Jo/
K0ybh87RJIqbX2SKL2KIx2pyxNE5Nt+2aqJ5CjcvyNSVB7JQ8jdGgaAa0XwXZ1u9
bhHdKq+iZ+50IFvElEUOcvMR5u5vnawZbTzqN7nmGO71YZP9tTU9J7YChHhlQ/FR
bepvuHgR+qvbhV3jhwDqoksWLJyReYs3M43azp6G+quY6yw8MonCVIni+T2mS3vC
sAz0G96y54SvtT7F+0x8JWC0L496x1ztCu7MJ2GIMVpdGpLgZfdT7f0CaZbs3/Yk
TW6VcZrJ6la1L2a5iujXCwQOFcgoNpb8gTn54IFVlxZUYjlAuGckc4ohoWaWp4ZW
f7KjOlCIoDlnD2zXqKLv7mJw6TOI1I1BYs/iB3BylODQCGrhY7HK1B1221Qzrp9M
21ZuuZgRt/DGQVKOKHyZtZsXMAq1p7vb7SN32yGw0Ux+Bxe61lfU9SFXtl600vN/
VXYMgCK9jBBWcJaFXiZ6iR9k1QbdDliKF3989WdAJqEryAIpppavXclcm4lZiLJd
RYptw2RgYUKdlB1+m2c8jH9TDG7DvZnC1N5mEc4+q78TgdjnerFhRuVBbBo3ucB/
2Z5xZZgw+lIenpvBAubyOE1LcTp1i+q4+gfsOhMnLb5ZwUoQ1tCn6zKbPA/pcUU2
bHUD0vUPV5JqwuluwduaVUnLIoImdgESOWGlETq1vL/lc2khdTekscVZBfi+TODs
WsVE4cNmScja1nOCNVvI6BWhrBs1I4WVGKXAuQ5meS6Oy1YYQEo862BxcbBeaaMb
IXY7zIKin33GxoXec8hK8ue2ylk1pZ3rq6zaAlwVdBojRTLnOKGQVggbK1wDhesq
HOfokQBOHsL94wD+6uFGH7mo9VNILGZUqX3WK4QIktjKGcGoWvLYQxNNXADhqnII
CG0wyOWQxHydWZKXjO5BemkF1/GlFtBnk21GCo1AchmUUh4nK/jPdjHkP1s0EU0s
yI5GzIhg5UNfuFqnDuQhOr3WRSSOm/M81+3LRaPc4j6kIYn3KLAxWoH07qCEGT3R
f9cXswJjDipKQ3MJJXp69S7Ut/fL33p4qje41flFJOicYtYO2BYS9YPMXTP68fdc
7IY7zWRYtL0fH99RpEdt+mmQb1RFpk93od7i7UNRxyqlyj7A0AWs9g4rkUZmyFfU
uPdxHtXUeR5duWZQS0AlBZYxe1M9aDQkYCBY4lx1Wn5av535XUTE0jDl9/Cc9K4y
fAexH/QiM4rmV97HHJ1fWv107Cp7Kgz/lHVvpcjgfM/4+ANF88GPKGqRoH8IVl4C
rrpkZYR8Ljus+VvtarSZaBOtupNs2V0ITtQragri2dgQeodYC+IxLnCf1DBeBKSV
/2u+WdDS8HXO+Og9oVaYXlmPE2js8ZrhNzJlQGLveG+PteKB3tB0SEheRM0B/nih
BBIif5aok+2dhecWGz3KVrUQzF+VuuwO7nHcgi5VI2lsulO1WprBCt3USrCd01Ny
gby/YO8fRkyroLPHNvajD0TQuDGV9wOqYH18/mH5R83LklHms0k0qvDIoqN2alIk
2Gy/41HoxCNrEtevf98nLFfyTArq4mgr/0rYwRBI34ej6As6oI7kT1b+KKGKEhde
8/sVpXlhHe4XwFYrhDuuSKottS+YdhsOzjlMtowJ+mBNg/61rkcq3nhEP/+tq4mu
UmYGYB5mR8S0jucTw1nw5/jkgS8aBkCfPvtXv4tcG0To/QXekOdkGECF45R7bv5A
TvX1fTUVuA6zqy+uLRV1ncPlMbwBWGxhkC1SiPXhglTroT/6wCZlLKwKEoDYuGi8
wkM9QgrLqvBkXogscl9mEqSGYA0bw52csFIF+YmDAB6XUxcbeyG4+Y42mD30FH1W
MApG/1HFb2r4ub7dudwSRzxX0BMVVMRgMKbmn12LeH2OiXxazYgCOL+ohM3O4dOf
KQMJGSbB+ovfXtZPyJN0EMMhjG51oerBi0KOiRYLcsPVksSI1SilMIjNcH9pYqkE
W/IttTg3rImayrCEM45tX2hdeks3cA4lGWzHUmwXPHaV7yl+EV4zxW8ojB32x2EF
vUyivPJLuO94DYCPZfZWnYPDpCd1HsunPsJ7azu8kcZmzuY2V2Cv/DxdovHG1Kvg
Vq5aTVxg0JdAEz3gGtOMLKvepKjPsp8/kNoQtd9LjXAUcp4kc/Jx1ifpkP1qfRqV
eY80bsb2MYnHAfZmAwcpDbSLxu89UyKQVeyxEzzvqXw95i5onamPaCoxrAAuCYLB
qKdFpqB17KTWEfjGpAJY7X2kOg4+uxzXyCVDUtDkrVfkWnPyWBk26SjLg4JKGAAQ
YFdhNP+gpVC2BiNybTV2LW9C2IK9SAg0FK/b+KyhmLkAxD0HWynCpxYl4BZKDGYy
fLLEnnSETFkEZeVF82R31EDaXdqIJE7xyXvAi5HQS6j+2d5FE3iLBayiLGg7jyky
F9PAUdWzy29s8/dsAPR7B4DETFD7mnVphlipHAeAEJYZlYKt8H3LEernVB96qgAq
p1shOXrjX0M6G0Erpid73NwzsKCT6DbHmhWeCx6hrwC8OilHunM/U/DiEIIsC0Pv
c1jvUrjYvkdxjIxg8nxq37QClXnauhYy4iwfa+q0iMtWim+B5NUN+r66paOLsHWK
vW/Tlz5zgP99vXCFVXOZpBx2dfbCaOQDRqFRNylzAitZGpygaviQomGTLyfdrrMW
ikwPmhj5nt6IQPiBe+diyBV3rjWaVcg29NwQx4v8a6fzRrRROqOwKgtni7GN0g9G
H9C/dsXroNU4qi/VgjvSpHkRFSXT7pIEgbbBwUjs6mANUUTmT+RoTVkqJgn8tCmQ
HGVETaQVYNlui3Pnf0kPLE0GCQrvMTz9PMh3+sbVp/m4T/2MM+pKNk0CtK5XItoO
uamKg9M0dOQc54oloqZZhNdUjNeERuEc4RyRVkdIbEylfVpnfi8xjroownEvA4Fd
C1KSLg9b/WdoSPJifjQjMJEa9i0urzR8gbMNVYV3R+BdrNwLd1tjc2KS0q3AHpR5
suNRglRjERA5xZCO/cLUT6A+eDfexFdgocIXhKXTc7NZMm7BuBci0SXvEadgRoYD
/iBHfcg3f+fXGWkO1J1lmOzPQNjD1GX534oH5FMZ33xHyjAE3V+dnRiZfPgESSfE
0c9SB6UckkEEMIISVXq8u+kdxFGRNtg2+txBOH8z4bz0bHBtbdLHi8n8hHyKkzWl
3OGuv9AQ6HjUTzUe3z95k3LCZyEgGKlz45n63rZet1QdTc2B0Q2vuVCnniL5L1T5
K/rHHdJRSzfRZJZINQsqu7qpHsG9wJXif/y1xM2UK72CIFdDlnij4epGqnH6jrzE
4g6AnELP4bziQ2EfJNLrTUWqoeNszAmY8xxQmi6HM4xlbFtaqE0yr1ANBbTIvPsp
usoYC7nRaQB2dW32tcoER6lYDNv7Cr1uTFE0OpkMN+k65/EFNv55kYzdbKBaiDXk
p44i9b/W1jqsduMr2JE+9g+aY/3AZ1UDQbEV8LhVhfLpXLcSEnNzWzDlv1eiwkEt
9MGOxI2TxA85RCtLSB5h2YXpo0qS0P60JvwGopPJ1gIfkoTHDKThZK6/tFgVGlLE
I0oOmtq7I2ibIVxy6to3+4UkPTDOGHZVzYebIPE62RNs9DsRSo5Jt8QoJF12bD3Z
v91n64xW8Y0CIqtgmLKUzAcsmVXu9n3hHK9md7Ib/KB9BPHCsimodKw4V+YQ8pOC
lhR2aPc+JXOHNqc8JL/+mhoqr1bK/FBB5tUF5vgGel2odRlZFIHHDh0rhSAf3f2f
Y9ZjgNhjRrvbmFWXpxn/AL8f5nag77Bdiyj8bEFslrMJPO1lfahP4LeaUgJeVocp
Ezvj+JLJxXJ1Mz1zY/ckAO5AjwYWFvJ8F4Dr7x9KyciTrcOEO9Tfy/1sHebd568c
/O/9/g8Wayi2RIMGVU9d9uWor6iwuulWu94seFaYY/IzwjAMb505LauSJ0uyIfbW
GwxCipdSR3iuufxMQmBCUL5yOJXahfrACv1Efz9XapLjY770vPRzSEV5UipK0zVa
wyHGRSjI10SGTWCybiWKpjyRyCnH9OfIE4VDv3XKuJk2JTGJzHm8p3tJSx5Ko9Da
RinK45TGs6uKgBtBzuFWz0lPtc99n8sf1HMvUtu2odh/zi8WHcd3dJU+i+P82oTs
UJ+8lG0p5snQGvlQbxlpLAH/ZzMhU+K/0kdAJMPjbbJb6gwgQd6c6d6ablbEi+JD
JQLeEH2slSFhgeNxsI7ZtX7ui6wQrRii8CHJCwgD2D69nA1juKOJwHZ/xmm95x8i
vNY06PlbDZW5qoTi8CLrRHJgZFRNzjKHf+QbwxA5rV7dwTvkKXkbeZaVEeM9HSze
aPWa8WOimJLJcl7RumI2LdYXHXEzksIDgrrAUx4Zycnt3h4VA+MLJ7T11onLAnbT
4D8118cNHOzDRVqW1ptkKaPYoAgsn7bQgAN9E9ubKJP5LCQd9GEyhp3zNSW3mCvW
R/Ipd/rdompOUVJi9/UkwC4tBHV+v1TYhyqF5eFlq7rpF/eIg5MO2J7nJgYU+7T/
8SDmkzWuZ5K82vWUKQsNSV5FjIbIzNMDiJdu/e3PfIlZBxvUhwta+Lr6euSJR101
0huyjUkIlG5+wRAjLxzhlrGz7K0qdgldKkSdNlIXOGeh6g7iI5iDNcfZVlaZYrN7
v9CwMlDbUsHg4dHsL/Z6sjn/MUqBwpG3vRpWPAd6Fbn7kzxJDXg7Wy70obJnKlYl
zkkS71ysCPldaKrLcaHHKo0Zy1+EDU00eZwHYhgGOo2i0eleibt08SrFqR6eVw25
PiSsG/9xO9mo1rxrO4Fh7f80gAid4sPcO+ffLFSJpFygvK66Jq8nyFA4tKb05Cki
6EGtbEEMcaujRngUMZBLUmFrdt2/wiLag5fcbvmqIMZfR2L28ZdbsHis91SzY+3p
WNCZtPKgpQqwrpRtgRPuok8O5Ly6Zx5r90m4lwStt5gbxxogrq2pGFzXN/7ZfViX
pwgWXKdwX6xzw+NnRJ1iJGE+pzZ8PW2Mgk+peWInczEJQ9mMXErhEmurGDxgLsu7
nj6llexQhFD3NqnXFpYl0St48DXIRC7crvBL5voCFDxTxAenM6JBRX6lUN1kn+Xu
CCdFqTsA3WvXuMkgIjDaibrXHnARs2mx/jDZ9IW7z65rD3zOUkefcMHViZmvU2KN
ukr7UuvJRVkOtAhkCTcj/uz48UFwOena6l9jPlOu5LAoPdtPEAyZ0vPRDLehwIMG
dvBXZXb8PYhwXAT/jteExiLXjY6UB6d/HtebNIydhBJn6+3jGlwlZM5X2fLx7IzO
j9ER0hCw1y8UevJ5qSJSL9QH8BBBxWwm66unAziQ5mSJpYD1fXqJkjLfy/pcPx6M
oVTWk+Vd6lGB0DKZCXBuYIYr9PbAsUrggJryGmnV0r7TOgwPlc99mtXiNjSQn0Nf
6TtGEuOxc4WVAuMJdb4Jf4zGZjGAlBiZMqTsAbhTGj5SkJcIQpnGTEsBTkFX/+EA
JHrhw5egk1AHtUbvDmHJpypChn5NbHaxAc4HMw9wPB8dbDoCg13XNoii7EgVxlVv
6/xEoHN1ZQaeJUe7evCygGpczFiwRbJox1Bt+xC47knEc5oKo+J5IHiyZrJFJxMz
5OnyxXUQbY/m/38dOtQHTrN/XC/MohQ7YFZcNgb04ytNFkt1TMkD8ETwWp/7PtUU
KLpPefPOb9RkZGUytJcNMdSqLJuprdDMcb7/u8d/Dmn/eQbZH/Pke3LvEIQ4PCJg
1GisClZh9aBz/BsM0FYXKg6oO3Msut1B56ezqUE/dPhusFCcGJ9gsoKAWd5dzfOc
h/D5zyur/XQgos4vsz06wxffE2pkPNchLull/Fy0jXIcO9gqqg/0pawNihS3jcLl
6QMLOo0K59cn19KYv6FcOYF6uULuT75jKC40HhZzL83dwtH6g37dO9E8KIekwrUT
Tg/9yL6rBnb5CH54lBiJGLJXwusnKaLKohcSaj5NBRF99BHKqZhlV4jOxZYqrhEE
g5nx4hwb0XbEZ3X4mFKs34Av6ZHgdkoexgkcRYpg7XDDqAWWsOyCQIdRsL2SREEw
3mng6V2X7RGsQLp20mLS0yy7knNITF529pEbotpWik9oqGwryU1LsRM/Y89DUiJv
W+I641GhpvIKtzH/ax0hwGNPqtHedrvdxsyh2bpLHfXT9Pfgl4rNIOapc34AqS/T
qQa+Z0IhaIF1Wt2TFWqYR0b36u2d4AxRO5QhurpYLMetqcDfENG6E0QRfV8Fnrji
6PYiSroQWr+kD2chLzwFysudXBWo7sDATXoWBIIylJH2dL3BYGia67kzYyXpKHul
unHFYysQ0tkIJLL9HJqK2TH/auISmVabUEeV1Ca4mCaUtpPOUvEFJ6Uf5mTaUaLC
7Ckhlsz8+zdKqOlF0mPdKIxfFAMjsDO0EhmfUpU4AklvyYySNDyNCiPXDClRgBev
wdX2sY2lDn12vW3wfcMgyBZX1xFEF1feJe+ZBTNw0XFq3MlpnEF0W8758XnQAgO4
NCl+EqLx0w9EdR+g5q0pPnfrfnWBgfKHpSMYGBNFo/86720dLTRgu8JWUldDu2Jr
5dhIaJJKv5PQ+XY4bTZAfQUHQsf1KOPDhrBn7aX1avmXP/Pjg3xU5zFuLp5EfL8w
YORxrxdjiFCjGjgWymsReQAU7SLcogaeNFor8pK8iECtxSF8+HEZ+rRTzq8UswCV
5WwXjX/rrRly8c2TmjcQhAKjp+YuQGZ36s1JIo9N9HZXMfVz6stzel/OfI/foO8I
d42r197PHuMs8T3l2UA1x1219iBEi4ZNO8Y8KXCJNHOOzJZ8WraM/Vu1FFNsqR9R
ZmwvpbpkkOc4jJAM2mQCGDg+GgTYYHUufMRqBTPOSZURKlA8l4Jf5ye3uEt3z6fE
N5L7JTqj4JjivHeXKp3bkYvVjolCi65hEGxfDyg6sB+x6qEAGtTxDKBeSbFO+k2w
hX4Bzu4lxIZynID2PbH1xOs80ZfNIg1b11U0K+XEzgF4kuo4utgnNvtWGiAE97rZ
M14CK8V1oQJe/YLUmp0IbpGRlYFzWoXuDP1+AIGSvWY4jUkTpT5fmOJlfgBrQMpt
Xo0ZRpGVf6JUfEOI7XfARIEZDjmHxFKh9YivJz6Uvdqjej4Snl6Z4eBLdbJXR9Rh
WoBbrEamfNNOVmjTLK7kLnvBqF8G/4OBfszYgeGkwN0408IMAQ9ZbyHo4qkEJtJe
HDyXYbiuO68Eq8SZRrHmAmP2iEPMk9J3onMZxAHhE7EgwSgq6gYgPY7AfZbANJ28
d0OcmPeLLNDdLdM54/J5tjzIv4CaLsrMIlYpqX/GVMEGigDVfjI2AvOXJVmrrFOk
Es8OtjxmcwMPcOdUcb7LVrEhRLXA6sEOQfYrQbgwzIkA3dqCqYXpqb1e3jBGaNkq
leipPdYVjViqMsOJIPxYBWKdgkB6b9t/TAVqNfl3XLMCdYYeNAPhWr9zsLChzBIk
Gz/ivkeGzA8BsDlUkkldQ/tlGPNC8fB2vPA6Lm7Si1Wx/832C8FkBs/ba2rE1ski
VI0d13Zc9pfCeiZp1g1dErVBUZ2AKbIwb6ci1MATN5SwiDOJkslH8GS6aX6xAMSp
hLNwMEM/68wtXKgnwUr1ujSC2nE+q7D4cWkxarjXM1J3D4OJNbSckuASA2Ucnq8/
N5pAH5S4WmNk0VfCL5stfFLvczaZJ8dwZHjBGZYYUDGsA5K9NqLBXIfDEp0u4nIy
LquqRIYQ9xO+qlCNp5OIfosySenFw2zVpA4c0OVKYEaFPT6+MkS5+W3IPZ83KehV
RiIFIGOEVzOrP6yLbNAqkSBkyjTI5A0CCmzaklfy5tPSnSWw2zTF5sM0GH8PA3tF
hBv2G9RUsvelO4xOGk/16P1ULs4WYCExXFqLxzVrPfgNaBQOpx2Q+JZIRLvsiM97
mGICDe6wbPdREIrBMEM+A/FRPDzJj0iuFhO9HWIIO/NiGJ+xsVJEzSG5/52XgBxQ
wMRbVNYlAuZc2tA4T0R9Ga/avnTWRUkpEcwB7tqyzgbef9JqCjmYwSzW0k3J4s1K
lxxl0e8GcoG8Gv4ib6ONBNXpNfC2wfnkneS0ZPcWJ5kvxkNBotBl4dCzEF2hwgo6
kgQTKXZC9FJJ8SWS2mhb7HwN5fwOSNCIvcQUMF9k4O0pR53e03rCKL6GkznA5Fjj
c94yqvAWkvs0bTmrpVDpKx7dlSp9oSSciocOzAIfsnFjD3AtDbCoxixL2I8hIcUe
7DeyN/igjzpPK8S9lPSkNKyy3dBcdgBEH5GIFhtknY+xlSUQsEu4yNtF7/7G/bjP
gpb7hIGG6Qw+fZWQdeD9hWFtr/GCyIh2Yp40SHojf6zt40gG4FnDDIq7tcwJOkt2
LTBn4rHIT9CI/ORvgdOG+bqUeHwkS/UmABEfAU/AlWp/apV6LZcijOQeit8Tq18l
8u/QjjSc0iBYmqeqs4AwX+9MvRyW5ICzRyYbDrCQbDxxIt81Na80XHk7NGX7ZB9e
2JU8W8D7vXTi7yEs3VuRx2DipHTw49FvNYfxIB+blu/o/EPF+MMVWBQ5Cz6fZCue
MRbO1/LlOLiiFF6KcxrM2NVKuMDbKo2u9AeLdPg5fncEHTLL7AwYftLwLX0exaFY
VWgffFNCYrqfPnMQvrb0YnJZhTqCh2/nd11wwAvUnlY1L02iRR4j99opH1r0wPfP
QkpnZe6joydcRQjH3yXYM3UXNFDVSdQCpKPcGrJG6ZzqZA3+4lnwpvkCrJLwW9zy
3v+6O41zmACUpuEmzex6UtWFjWU5nWcRwt/ehc/3oZLBs9q9oME9HPit37gZEfUK
tQV4yADjlv/y/qqgBDhaUecWXupW9GNsPVikazufaVt4lDycXW6eEjVAPOeceyiE
qwwznlONtZAg7b3ieR2JeIpsxKa6NN+8tBFxzB7O90VAqnJFQEps6ryMfeLdTK/e
acQpEOgrr2mDoBeTa7HjG0jqvUOv163d+dvKqI9w9e4g0y02eBu9Y6NXIMLNGiRd
Gi+WLIPdwYvJhegba++sVZzrB/GwqBD4UVeM0h7mEYRskCXTzrM83vPQTPHpTwkW
47qu+K70F46RP5m3+qQ7VnOt/IXS7oiO5ylvKR2RUnLZHUsarCjFHnymoUPeaQHL
RT64OdD39/nzhL8jrV4aWA9Uw06O4AHHcDW4cIdJ9yPDBoxFtg0BSqC08S9mPwfq
IYH8VWmOO8uFNtlTxqQo2NlTLih8dBTcKxtvQoAtgXCd8PjwB23dqQeG78gGEfds
r2xylOEhh16f0iLrNC+hOqbf+Vs9jiPYD+lXOIKliDUdGluRmct+M4WEvCZV/HwN
zPUI73sl0cZDDS/KiBjiz5Ehsmaf6HZ8HIAG5XHBc8z3tEHvwmRLm+nCM9ReCeiU
voLTuO28GJzhFIKo02QPUNrtQ6NTW7OvDCyqcqnaPbIimFCqnXoskCxh8dj4PS/v
dVc1RuR1zTK2igGEefJncHtmrZbD8f1JVi2ytJrVxsYrlXiPh5jiA8aIqp9psW6X
mtwXTDkiUpnjgKdW8rHI85iFYTCHqm8mcQwYpxGuRtQTA2WKPSKfu3mNjk12YAEv
F2jXGiO1CKBdnLKGm2q4gGghKG2P8qPF+uv60znatPR3pgiHUWpy2nZkbQqChO/o
1Ct61qHTN45UZMbdyOgVYUd1Vko7NtqXjc/G8SzaD5rFmfWRY1fTkjohjuxtWEeg
HJjT1nkPdHv5EFjS/XOtSUWwwJVKyYVfFDKm3i4kHxd+ubRSjm78Itx/v3k5fzE7
5tg7NZ473PNZ0hpYS89/ccwiu51ZCNIvEAK66zIzRhMvayLEnqCMnVAhRJcyXMdZ
tqCzv9FiiPDz3X3oboHhSYuA8YoqYhIvjwnNW5iTpfnrX/Il5UOOY2LK+3H4aXja
3u2o4hWxtQNTk666KTreMbG8uQduDr6QrM7DnihL+YejLbUw6cFXHNDOjeyAnozc
rLzKUeMzgvgOqWop9GMDEUF7H+qH+r3dh6Z/k3CmiigiV8f8ASk225oBeAQfyQGZ
51b3AZ88dOKWeRLU/P1b7gSxfyS+CrN2W/JZK+yKuij+Eo5i6jEz/8J34bGpjJij
uZy2q6qR1MLnvusCBR5iOotWlRz0W9foipjjWJAyJti2G6cuk1vJ7SO4+N33ngD0
2XARA47pDosl2X5ebJ+lIA==
`protect END_PROTECTED
