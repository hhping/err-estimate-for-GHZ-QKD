`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmuTQmw3ohCeWfJDnXgYM9CH6zZFFk9dd6hRU4zwXBBtLkSv57U1yihXNWXHI0p4
q6cTpYlU6ErxkQ4Ydpqd+hLRWhFVhEpnVoF7wkRMBWkTsyH+rohm100ncTZM0fIj
QoiSG9I0memVcyAVfjQYeN5kOlnIprv1adWEpN+bKB0m0RiYRzprzr4ESGvWHBUV
UIY176t/wPjJAPXKBBZSkoWhYMBQM3aNPBNQ8pzNZKN52evkDx6bqgKiSt7AjvU1
MsIqjDwxKbIfn8TGvYATzJNUkxdeJyzhwf6EdEpjNuQlNpWxlvkNFGxwZdH+6d0b
YPDYfTpQqw6m8PH6uJ8tKGB10VzKoJObP66wL09AKWOLMjO6iaukhl+A4F90sg9q
qIJ48x4i3DcBD1jTHnGKQj7QhdTfyTj7Nu+FClf6GrwHeqrku8OA8Ts3py+URwTX
e+hnmlSRkYugAQSwCivpjp+YaNBy5szZELEpsvYYAsYNHC2HA18dBTheIBuPQNS9
0iveBTXOqEOE0Lb6jKjYhWcfxeQIpBWL3kx3jRNrOE4tx1uJzrOm+v3+DhGPMjbV
XpBkX9FukkZciHNN0Fh2yezrWcMYAvGgn6Q9onZMIpI9npzfafxgr/PL6fKxvGW6
KczPOOHqsrF3PKYCsk8faVFr6SewSEp9hWYrmhm4HwLdPbTxwuMIDV9+/tMpKLEZ
XytfBbSclYxY98Av4i9DBU6Gz+4jhFj+SXdIDC7JXUMSPfUXtqfy/K8zbgWk59eO
nGtkRk6rdOBYAf2rX308x0lsqiFZWcfer54QK5p3lxvW6Rj759YwnRrq2u2Jm9oS
ZDU/aJQeHfQMmbhPKdn2SpbTZMA84FN08t4edM74LVubczUvd3Sx6o8CCPE4Fpdx
uFttAVScKFpG07Lxl2k5qX4W/w7YlQLwI3858HIK4Pa4Ze+TZhGSQdPBW5IBvJ+m
00mLJF0AiFEFDdnHc2i/FX3GAtDv1LeK5XN5xvcCZQvE+ZPdtpBBWWdw4tZseKPq
FfUaAoHotnLEUk2Hz9NiRihZLzFubQaP6a1Ok3bpBmw56AXzFiLftLD4zKV4tUIQ
JOLQ93liE3n96Yei9PxIsB+al35ZtAPmFE/vSJ/VP6EY3BzZp8c8JnZL/rlc/SNy
BJVDvdciit9tBKC3r9GHlC2iljp7EeFHhfvSxl8Vu6qAvSLpz8LhDezDh+MnSrHK
uC+zzZsO2r8CZ5uKvjZlOZCBIn0zzE9sw7EBFkEurzo+BjHMexYzJZTqze6KHSyZ
A9QoWfWh4+d6cN53cmgjNdpWu+1bNLhwWkoQZU/Yno9mZlB71JB4Z1j/UdqjI21G
7Mkr/39Tn1vfNikEI+LnvparS+DAhyNTkrLG/4cm5BOAfws2JhdCY+OuXL2hF9uA
tCFuHp9aJZQPVABpFUlMxbBphS8VIuiwFDm0jCL+KalS0MhgZolBSmnL25pv1Usw
GVAxJY7OZGy6Fd5KEvv3+9dzNPRxFJx9O6FsVp4r6+pxpecJTevZvmHKLwr44vCf
ofRyvM0e2HEHRBXGfU2jbrMpvUnf8LclWboh6LfIBjTkdFmmTcOmywtfwuQF2bMj
8AMBqKBXoa7eEDyk+o8ebLJgCb20ZLP4o5yQeMN/A8Tiqrri2+yoPFpmgY2sN+98
cJF39z2fqUUTyWdklsOpWn38DpAmzU5EQ0xhFroOHClwX0nAw/0Y7C7+aYxQllpE
qlo+TyGvBoKcW5XzDNH3dNhM8OVKMwD9bK2pVzd110MpXQpwaf1LBNs6jKoDVE9J
RlPJ7Hc/NJlBlLAbrjyAJNjij6y0t7VbqKlFQE1AwmVm9GQxOAyXBznQ4blzyFBi
sz2TsRiEQahmUfoV245TwKIjSqFl6LcOxDwiE44H2P+WabaY4+/gt16RhLs9bhhs
pH5RcxSRkYGB2LJMjcUiBoTSAmKrq1wPIoqLGroMfpXpC4gqT29DmGZmuOKpKwIe
tyAS2nV+jsqGVYxTA+6EvKgMVZbFMrh/cj11NGpLSIEzCXDVCDQ2N5B/a128u7jm
AfG8lypdNwCBQ0aqVTg3sb+iD9mpSYzeY+mWrS9YXbFiNv+oyLaC8PYLa6/oA95m
FLK8hwjUuEb6eES3CzcJh8bzzlvc1DoBHmb8kU+5LW70/k/vnzzlinghkvbvOqbt
fVmtv7jCM/mxjw5iHmONFEYrMzhHD2EQQ6mbh/6N3MSlpUzjfmbf3+B1EfsGarFC
3OqnSCUE+asEHzgXdzEh3s03FOm8RkL2jXDEUWlueauRHTG7e8khQACMUghjY9O5
F65L2zwkKIvD5ds1R39tlQ3wiFWi3jav+zf3CsixCg0=
`protect END_PROTECTED
