`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEX5MJK/cLY7nYPFCF6lf+ZeN3ViL1zPV0LV9vNNI/+Z/pATth9peMqexkdbqh3i
3ZpbOja1meiMltkKnQYkOpjr4uBm+4OgSfrs7diYMV5DxgHLtUipUTwxK5rTXOC9
mTLqmoj3HiI4FuAmYQO5+e7B9/GLPLG3IbNMfTGu3GuKXimNY1k2oC56hClnRk8P
qqhA4meKx0fGQoJ4yS44+r/7sO6g1G6+rCzGFlxblvlWWg/nMVWD3ElIHVJCuBd6
62hybdRXkwskEziKB+Ey6lJkyJbbaTAX1v395vEQSKbz78w0OPi29Wt9f0U9N25n
6d9tbaScO1s4kEBVtYNkSSmS4M+ew1Bu+Tn2zpKEUIRBdFkOsQNQWEi0UmGgipke
xSfL5DZHGvjd/OhwiVG5n/y/YJ2vbeuzX51mIBhx7vdCs6U0FN/roZImzrx/DMr9
23MF8GL3vaxGIMf9y9P1wdU96E6xb3zgNGfpO7R+GYsUZdRyQcXmgjBU6wRp2ohu
R6wxXAsd4mPwW9oh1L66yneI53E/i3GlUZzF4qvG40mGixsolCw9xsILYj+YIac2
gmN3gZtNgRUPBC4jfH8jdUNxVfAyT2ew1kNmQU2B156HYzuKei5+RaLbf+gEiFm+
U0bxF508A5Y7QkYDZ2nj5iPToKouPqJ9OrT/Vrjyl/b7cRrFi7wtWsw0Z2o5NF0e
FI0Bbbcu3erT01c21iwqK1tY0zbQNwe3H9mQE0ozz+PVnn90U2Fvl5wv4bkL1AWR
lea0ZLw+MH7goj9vNMQBrEdpSbve+IHH8pQq7CvFlAf64JZTD6HilWCVv0/PkUQI
FcJGhZPhic1CRUI+dWd3DfGCTTasIN0WRpgi4nLXR96kqBJl82jybrrujY0ZqzpD
4cK09E+3JwBx3vGqh9YVjxCyHjvABmxsENDD29aj/kCgvGRCdH0wNOpF4N9gw/yO
7JGFRJXlaxhS5KjhOUrJ3lLw3BBzMa9o0TiQBfTEELmxXmRst5avaOBWjpsiI3Wq
WV9oFTXCllqmE/WSwLZm1S1TBjieh2VgggGW+3HoHGow+5cQLyXsRRyFtR22iqQE
ZV++vZ0k+FJ/3QOCtn2TurkZDFSckMInc3+sqBHovBhi2RZvZM536we+FzUAfKri
Urs44RZRhPIWInBNAFmZN8qZ7XQwhL/dDMRGgEpQi5/S+buncjSIj5WpDz4F9IEw
Hr3940X5SarGx5eHoqSmuzmxNaPm1ER9JD0JjReIHsBrPlRVg93cX7KPZUEqlHkm
TneuP4sEM0e56pqMyDZigfhAiMZiFkXCn91DM5caClQ0MOkmVygjPEbTlEdNq+KJ
`protect END_PROTECTED
