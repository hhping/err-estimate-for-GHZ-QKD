`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/raCJx4DcpmHtoqMZ0fB8MbYCJsR4PQc2GqfCg7VzA40xZIwkDoETn2vKfbBkt2S
RII+xCmfCRLx76Q5HxEiD4lyLoW0FsHTZL4y/K9rZYcPWdU07Qu1EMxt6Esn346D
28YfBGiOGszxrhyhi1yUCJEr6q8SBO1ZJTF7QnDTsqtVik/Mxk2P6QD30XgmXWVv
z7CUOxzEGSXUJAsc50Vt4CvZIptBqI6qbp++9bkoBGfQEHRtWVs/ZysoUZt8hwXq
D1miqNxAtvknfDxOpZOc4+QzmiR16YXsJPejxjrxz94WcIiLuj4L+/H8J0SjQCqJ
qDtCmGfSU9x19JWmnw2S+6R8KMDXMO8VGQNte0Io+RpxLWg1sqOZzSVHQJvJT6nG
1pbNvATugZNDGHMMY8iQwNdyLkwdxLciyfBGg/pkQMENxp76W+v6JDl3O+CTo/Ox
fR92hBmOsPSk6lvsxRGNGB5Bx14vln+RL5uT7JjOY10vE4aqb7OJOo3TGDe89xP7
/bFn+HgBohKL5ALCoyKKZj9ZCitAU+M65PAiHxEOpyB6t6q8sOq/wDQx5ZE9l24e
Nur/bbDLVSQj6hN8maEUlycQ5jGDp2GRrI35G/5NrcQIoNLezuhi0dvMvhSVsr3X
jvEmJLF9G02MjAmLcHGPpgUJKGuNzIaUgqeubye7rXpd/ULvQFRJd1o8m0f39N7d
urm4Plx4Eg0v5hY9/zwlwwDK8RCIy3l4Cu/GxIIQI7j+oZh/7QsFgkp5OgGK+4yh
y2uf8R6/P7fx6UwACYryugmkj5VEB72aUxFERIpqZ0UGDjmCiXgvEO5e/00DT9tY
NUoItWs3BpTatvqsS6q4zozuGNbdeW1PawdHCz6c9bwbok42hM9YJmTAkpeL64sd
hKS5q+oyeLeupff2PvunpTaGkha0XBTkENcp1jJq7Vy9wP27IguhY8kmgqIvPzu5
/p3A/O+WCExYCnwhsAYv0Eq8kpuHLtiBF+Kb905UzEIfIyPTPuudMM29E3YuCajF
pdHooT5C6bT4YvGPejWK5jd0lvXhHekPx1ap//oXoxOY6EkHFa2zq8ANlTQemfom
ldEP65fG6kNu8t8EI3gkL2GZe81sZ3EzPC/9TlSs6eNR0kjqXSQLn4mhJm8JH/ve
av+qZ19CCkafTLz75FkPM5EJuBImP2oF2HkBPoKuHGnXNpw+Wn0oyD3yO2PPLbv6
X4PWj5NFMQr9OvZdXWo7frMuf/Bg4CtcUwjjMVeP7iu6L+fnrEKT7qfY+MQJa7gl
/cu45YoDUrBwya1Nd1U28HfzxOXnFo1itclCpfRE5OvDEHWLkRucmrBa+mxlcirY
ZhgL0tA7GUoY3TvtQ8SkWafb917kET/Ni5N+QKOdH/GVmNp45iuazJKpXlTPk2eQ
fj53xuVYlXSA34deK6+1UErhqxG7ETnpr0kcUiuMsuyYF0sao+N1o6SQaGryS8To
zBn9WvR3kWNulh+VEBQ2cR6Km5ZPpmi0U53+/WDjgGMusKNU46bv8k4YNOv0xtng
zKRI7olLM7MFMXnH+mjaDvGX+hztsN/2P9IN1yLx7AYU74SbxvAD0pYnExkHnII6
SjcTFCavhdNAMQDHZ0y9oZmZ5vxijas9WIfj8a0SjXWd0xRKJ0jk14ki6m5FzfOk
v3PtscGwCS0PyVDGzsO4Pj/4vKv3SYnsZIEU5HIw5A32bnq4e6O8ntwh/u5xMqQX
Qj6uxItli2pEwwrMM36X2RZxabaS8HClXphl/NB38VpUK5J20U4LHqReVWzHr8fG
fEpTLxpAUJI+nFajAKeNK88LpWxWEnQAyI86dhWbUfuoPwyw+xdHRjjP397x9iYd
bvXTQ/2SAr1b7XF51amAlBoj7loIriM7KT+zrgrerhFHCDXRaxcn0UWvEZuevtII
tTTC4MntwN+mF3exkoPpRLyDmOOY3hqq2RCldwScuVaA5L2Pi3rir4CBZD6nJKWk
`protect END_PROTECTED
