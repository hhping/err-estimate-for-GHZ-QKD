`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2NIzah3e3MP+DaurxYwmCM3mt8fz6wLYd0Bukd9qeaqNJUVOLvxtIvndE5A4V8NW
vWXo3+w2nh+dHLTC5Vot3LeugOHbaNSQBS0d3FkvTftDfCQmw63XT62pimQuXTB3
UnKM+9p2v5V6/VmjMwBpUkpSP56fw9M8NcwAp0Uh795i1NS3sGisGfzDmgCWs7AQ
GLGjklGmv12texZ+0UXW3BJ+4QpXs8cIMM3FFoNIb9yW1cod4HdPEQXA5DF6mNba
djWDlAuGuBKDevGtkTuJEWSlxg4Ioz9baSldpkc7boBRRi+kDKV09lenB7zsdzdK
H6uatJ0P1fXu5hMuazZ5NdPpCPygt1msRqe02FEqcwDC8o726svFSdbJq90ULl4M
KYQKGkXWm+0bDAik8+EPMm1goawiO0TBr/h0mQQSkjAaBO0NA7GoMREM3N7LBXd/
r+GqAK5EhEog4yEQWkCsuJ2+6Gi7+HLRZFwN9NGsC3hYtV7tdUD9MqgRxiQTbCP1
1Qf+ik+O0/67X58iEQPbEcpbAxawAlKwQ5nbjL1C8vICcyMnp2glFVwutVUBW1eM
v7chkGo5H65v2J6eWYIfsxYOwWpd1JNHglIBRP+b6WhNmaZi/tYuNK465UrjL709
A6xfy93foGEKAeXO2hqRZ9lbdh8Xz7BLcvSdCHzwOpbN2y5aZJU7UJnQ7NZcdyCu
zmulimuFRCnI5PC9nTeEtBlakY/N0iDWaNQ8UgiEf0uGJ88SiSzV1yl4rEJJ8hXF
wmZlYjxUjRYoM2Gc5Ka40x7QbSjaruV/Hj75B52XbOEbJ8WVr8I/deEOPnfAxfoe
GSJD28jjdZMy5FDacZmRgQ==
`protect END_PROTECTED
