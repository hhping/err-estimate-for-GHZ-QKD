`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cjGACmCyH80V7I1rDiEwpvLoUEd03IKa3LOMF5jNAd4mIkSiNNZ3bToETgTkCya0
J09ZRSG+jMT1catiQZS+hDbsd+ahemfuWUlOkOLFWrio/DIPmO4UokLA76Ko03mw
tQKNGOCdFx2DDyTG+IHH8uyJQzJDKbgfyufyd+EgKr1FxA3NaAzqE/6KpebdCC5+
GsstXL69FynEnJCh9+IMhdKh+mvY4BTAMZ+YpNyPOkIG+oQVs0v+OzuIh2XhBJiE
/uD+91geYCwuhVzqGkEy9vu1TyRNz4hbDBj3hk+1iRfgEyCkH4E8EDoyHKUNFgP0
4ZNnPpNxKMZCKDAOPHwret8okf9lrzW+WIj0LgMOnkKspo97CXgNfIW1ehkCA1Tl
WL9H9xenR1fNxKBmX1dkJJg3bwRMhjJvgdEFXvZjDwR1HhwRBmQmqwAyeZnoh1+V
XzPKg/wDV5EH/Lc+WMfqeePjMj8Odk+9nlQJ6GI3acTW5Aj/5uX2DO77fyAhHXbv
tRcpG2SicafSWyyuRCUJEYy2sRW7E7Hdxqws26xD432Dj4UoCZNlI+Xv2cX14rM7
n9j0fkR3GTkl95XVVk1gCH7eThoWC9cxR4Hl5IvFr2RRld8jE3+8EWHHW5leYzko
OBj+BYC5vXAQhbHbQLruFm/wykdJJ9XfLiLW49+Md1ugGzLxjQHVwNB4QJ07i1yi
a9JTTJmjOsukxc3bd73J+0vsnu1b2NuE7NZF6g1iD/LcV3eI/DTeSbKEXPrbHoA4
z3y4FBNEP2yKhNeFCk2rspvt2gJmNoUrN01Oh06pK8F1e5aSqg9s0jlp41FDPSHB
w6Hq+vmohi/mJllhLCdzUGbDsrdeAJxWuSyOHWOhh7gUC2+4jQM+A5ko946iQVLG
nYwN4oJEPDQM9Ri++W5qd7apH/oW/ccIzuM8UUlVjWfkPVPGPyXShZu9nfixziM4
ny3TQAnv8JNAQLVKlGUjToA/CTOay1ravdTAJzp8lpPvf+FyuJqDuk9DDO9BzTK/
2d39HZozYtvVbuMw1O+vsmA/PRe2HvEcAQYAkiohppGlo7MoV/DcYlt3CsBH8bvB
C8fqiw9m/c3i3XE8VWLQGtquvpKI0QSHbbxvkCF/ZEopSI2PNgoHaaKRZG4lSJw3
23uPL4reR+SDU/QPUITcCFJXJexqT3DroD9vb2zpfB7gdcEsXHJUfhpLryvlMQZ9
48K/Bpoxi6XsuiZ8xG7gWFjIlZ4+irzmN0Q255781CEYUcco+s1+dYmHnbta0XJq
aBtlc54eXahqvyxxTVUcG0GN2YnUWlCEMFuJ1cAOL5uKgUF1i3e93tdwu1xQRSP3
ViU7Qsb9SQrT20Dnar4GSMa9XI7Qn2BtMZ2SQC7QsFGQ92q6MM5yVUO1ow5Klglu
I+cTKRXioMyBg3fmuGlEEYG3eBL5BF1HarPQmuS4nggSkbryrD0DXN98as7/5dx5
LJwDfFf0m3InZiSxACt8NtOqiGTSBMnuBwMU3w5mYyjKz7ntMsQxz5nCaxvaKIW8
Bufsfpn53Itre8FhggZpTUfYRLNSmdIyBQ6ZnHRlRod0zZ2CkKqAAXgvhMyO5EIo
+ww4vIwsEGc3xiQ3z5Xfc7EtYrzFrg+vRc1nsH+MXMBH6XXEkK7Eugyx+JgPw3NV
eisEaJXgSIQUrza1jCcScS000u7CwnxJYtrOHnafQIp4IX52y45keH25GzhwSu0q
RYEsuXyewFP2/PDdeAgSCS7GVrnVXl6vj/dv9C169Lr534/9CRjWriJl0OqEuuHb
UVewU4/8AmnV9SfplszcOlEaHJX3asm6oEGHADzubcI=
`protect END_PROTECTED
