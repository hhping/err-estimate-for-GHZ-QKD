`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6WsVNWXM+dMBdZ0lN1qpcBqj/e5UCbNjQsaDWYuUqDlaS5f6r0TKnaLSaHMfGfv
cFMfBkTTnlHaVxwKc0tXmkN7+2qP+vldbnND12Y1a/XqNnYboyPIm9vBcJh1Yi13
sOyfO8dkhmde5HxrklUfk3ZKoZdyvcpXn3bDqoocJYctOCQERTNt6Q2qEkuSGEK3
LCJ+mdo803nUOfAneisfODIRfvm4CFW1ghQO3J+IoiiQ6czk7rxvCkExiLCyhp6z
E5H2DKiXZdKFMd5AmABRStoR0Aoxv7VDJXa5dY9ZN7PhZseyNFvT5otIgTJwEt5U
vzBKGniHRajRooxfzR1YgYdUu+M+pHF5gdJaSdIrLCtOhtxUp2Lhw+SLiaadcENF
Iso0OJ2DQdoV4rR7Cwr0LpBJPpobZuRBUX6lE57ZZNeF4zci3ND8jr3X9Aru3E94
jQSwQw6uzYZocoGLKvxFlKqADUMPaRBtbxrQzmD7Nnr/pgzNiLRuOK1R1RB+F8fu
k1i5pEh2qRQAEyxrNCp42kmzipXZ8I36XS0+WwDl9+MWC23Cp2vPb1V+c6ce6iDu
MOsFnWH9gsSLq5YZuAxvTzDMy89TFUnkNKMyW3/fueeQ7/ifoQ0U026oZAgmvO97
ZeGyoQb9T/5Pv/4QR4NEzknI1Is5ocZfvlzqkqRh97XbNsDNBZa6YwC155zjp8tP
M+K9a4KGgoShUyT382PjbBwwZXzm3LbW+cv5/Gb8ArYU7z9Hnd8QeYf+shTKkGsk
DY/MI2CSrSWgF/eHWOWCM94UeMOSkeh/X/JoRkp+TKO+53T2pMDYT1Lf84oSU8UJ
WW+HIjk1ZKzd/JQTVSbekyUgVgVzvejDHYdILfmRdw8CTt/QJtxQKXzBPTZjDJe7
ZXUiNMWvErI/yyN2+w920oJ4/wN5nQPHWZBLaWh69UV0Cq2bRy5YZPm2hleES33s
pUlU/kHMDtCjYY7FIaOfy15AAC5hn+sQJKRXRmmyqX0290s0U8W81wirIR8QMnWP
3vpsXy7uoHHsD4Q4E+C8dgcfVvdlcjiXvF4bgFbooCs=
`protect END_PROTECTED
