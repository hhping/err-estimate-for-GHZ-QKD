`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQttYrB81+gneXnqVW+yWLVmDxQzDH9wr8FojfdIBFpVGM8cC+xk3rO+s5R1GbkQ
/rPQazUFTeGsbGP+RIIu9rlMOxiK1tnYS/c7rfGFbg4u01GRRSzG/5sj7lSve5Ks
J3oX3ha+6B03aJ9nhVFtpgfo8i2bHyWs8K2M+IKS58c=
`protect END_PROTECTED
