`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xv2ICawsizFkmQSBaiRitAkRnAwLAM23OAVl9HCRFVrzNidUWDorZGnL6JSHAmrW
FxvYkaW6hpDS90+5hBEWegHhkmktE8Nu/86tlD+dN5QczecNT812ePx3ONFPoDt/
HNDGfqa7svT9QWaCjiTMOGjqdsLuBAyx12muu3OcIsVo46U4e9Cp8WI0CEXRpCkH
7d5GjrUaboVamINQkkJQcrFU9ZhxH3+sq3q6xQ6hexJV8c+a1PBKmwsDpGyxx0tI
xkpsLKPk6DTnsjcL3XrBS0V4T1mlDjmDEpEAWa8DuMXp8niQ9dRb5jbYxgjPNLXl
YbJ0XgRH0o5fqNo0noavBWYiMEoZsUbJvs8Hheqr4PE0KQghww0Om166PglSv3r5
PBe7LNh4urbhHayY0/NBSKxPcPMjuiiN9Wo6uR0Spbx8UP2zebxcjNCUx5kGhQ98
CK+sYtBaRfcWfzYA4cgvrybpgqhAnwy+FrId9fLiatOz4hl989UtIAcGc/QJBeq9
LXfedcgwKm764XEboNYEUYvY+DL7uJImg6BFwwVSUE+FdHGZCXRVfSUSHcixdVhE
3vNxxkhjjW+Jgas1cq75N3MMmZk2ZlzPSbgSrPXUTN7TnzthEdy5/st8GDNpnGBG
NNXOVWSjgKkrxYTcGxmN0y/L/rPuPbCuOBJOC15iTgqAWeIKowWAvZuvJ9xTFUG/
dzav76cIEuZzxduCJVQoJBA2r1YfKk37hMWi2b/V/PAu5dFwsjxZIWs7rdjLDgBx
ZVZrZMmYt8+1OZQx5cL2/gU07wdc6nnPnCzTk33kZfdfFZd31i02pdNQCSMn3EDM
cif4ujnMLdsoLXZP/MLDdPVFy1QIb39cCQRn8oPXo96SkmLgpnduQp9Ga6mo8lTd
+H+EhgIyr4m7eaEANm20Z552j2rd/gz+hZ+wxhb8w461Qgs3FyDnOmiqzbIvNBGD
FOVh3BRy8MEIXPvJ5Z8y9JTUgheke/g2/MLId0wj5ToYlmBuNWYWJdzjh47hZs23
nArmEtY3DIiU1mr7uZmKkUdy+9obiWNmHdZKmMGkWkugdzR9BJJRo8/LT1tQKL+W
xCKi3Q2T7VMkQQkqZFptPajVANGi07NrKw/RqJsul1E17lKsu7R/Gz21KrIP9gEd
2gyR+cdjrTj3oM/MsOtlCOkLnw0kuZnjmcmQNRbp5bbZc1wgvJyRyvtqkbZ18JAD
GVmTn5URi9xkc+7guAMGxdtNVjWZNO2F5ItKKws688tkaZv1j6EH4Xny5HtYexUz
A9dD5j1Gr7XbTAE4+CdMs69ezqejAfDxID7iHjggvJt71IoYqbmBqDxWhX6SXrL0
ieo00AQDtJeaRaIsFpSPNHUYTENEb1T08NrELX7BaMc5b6hLgJ0N8Dku0vx+YmNT
UhnksbZtxgTFbLUamK85pz2jAKdCpx1ThnlTxbFwSPTKBTBXAgNQDOmWTFlK1Q4o
hTLQAhyCnUEBbv4notIomFI5H6VZfwRt6vIv7y5UinB2+jUCEhS3esM87Mn7KYzT
tequaTDnotque479MR5YBgztd0MMwR/jfOR4kTVvaW7XUHa4d+jenGHWz/Z2sMh0
O/TsFeDJRLhtVoM81zrfTdUOn487eJNdIgRQc15Vdb/MqOIX/6gisgTXVsCiJIWi
wembu8x/6XYFrvUWwVBO8QZIePyCPHszl7Eigvd/+y18nMLvJTI3nX4dXqE3rPP7
aw88zmirJm2lRHO7MdzGnBnButrcagkUgqywe3T9BGeX7yyc7f2giRm4S78kpiGL
LAvvZNEw1Ich/lxF8yrfrGwYquuULhZ5CjRID8kSC/KF39LrEsC/95HOLW/LbGeU
OAJrbfSJZlww4cUrpsN6RKAE5Qhcl/NrqseTy4qKDA0RPWO6eKfeawYcJv6KB62z
EaNO9bin43s00uuT5QDkdcHaPHbjl2D22GvnTZmLVGiiTF+T/9D2XHfuRH1imA/I
Bb/7eE8Dx7tOgNu1leTPFh/kQbf2roZz+75NPfzW58gZmgYjpyZ5XteDqRB2aePL
S+/s/Tl55M+WO5kxBIqx6P7KqzNjISR92htNvwAajbPEBhp1XBAo1fIZ4infBFw/
Z6uvrbWKtQUlUVyAVnwQK+NeyxNqqaPowxJCs2+AXqZkgGBp/uGmdrbMP60TbGhs
5vp/NJx/n2ZiifudwtlZ1HYzQoCEKQULbXiomTOtrnq8jRA2+4B1+aOby9A0fcJi
3j7f++9NBl4svw/DPvXF0gT2zRC8/ZJyKad3nEOGIAj2SlZa2mXG6Yo+yHSperH8
nlGYcYYi3xDnr6m01ksNm50oFQAhGpae9vVvhWUz3FhoBwI6LNyHAdSwA+xEqpro
lgm3HBB9ZnYkmQfmlBoG3c5j4+oCJVY8OPdFO0e4eTega6U5vIW01HHAwQ+X75G3
Wla5P4AX8vDA6F1GLO8C6o6fAubgvNEbbc2bfJ5p9yvB5Ajr9Q2CqMuSSVor0Aiv
4tG4yb/CE/mzrmdM7sq2XhBgutbpZn2/+MaFGJOOtlCaUphSWmoKq5nca9fm1a43
izZE8eJpvvoneYXV0cy3B9BFXw+FUlSX/RZrQEdr7shrrAI75zFaKL/nU1fGiuKJ
4zrhr2/ZaaWWZp2O2TbGZF56RbJMfhATsBSL7Gt245//1Ub+y4W3weZL5Sr72roS
waPoT5ic4TuH9G+TjCR5fcU4xXA/eUe5evidlie8plOuEu7l8ldDBrw+p0HSYLQj
Ywh01cEW1D4T1lEHm3199LwZ55UbcDmoIkXP09qO2VbEEXr7zmOm/g5BmhJf8RvK
8ZtZELUWhc8adJl5zT5+C1zFMy0lKkU34loSaxhAOlQmYjyGpix7eKAOyhIv783E
2DNSRDYT3DtaWB2jNAxFpk9uDqhyU3rnotFgsbou6B2uEK/Ho2sRxQ+7TfNYJSvF
e3ehi9nb3SVkk2rNJhlaaNO5J0HC0OLuRkD7tW2K18sKDSBRcPaDDw+1IEa8gWTO
E7sYdDpvQ8Thi6BzLA7tpLfVSjS1lDyLRaBQcW7qCab9vHeKlRXeVoxJ29ZS8Gq6
nFGCNwuKOPPAs7V//zIBIYLGBFHSzyfNfxZty2JAWQ1lcBjpPhjDDLg8d7yDrLsN
LshSska/xVbh4p8BBW4Ua6B7JmDuYEOwTczG/OtElyQEyQvWH0Wjy53bCZ0mQ/B6
Sjv+UUrb0eWdyoQGD/fXGIdQQwTnTqWsA0+2/pmjqzW2fSIhx8zNx3TcfjyeYlLT
0nXz2e9sUQJVu7EqwS9fBYiZ+FzVAM34NJ79jNXJY8lux4kdAFzj9vBK6urnUffz
IuBHRAK1ownamMkJBIrzXY6C99aezsDxsorbjSUVODurcrXKzswhLyifn+GG3b8s
9sDpqu4NGFOlh5gtLbkLqxYl8Cnic7kFZSJiDQlFVtO7aNhI7GKlaY0pzAt9jd0Q
JCB0K2Z9D3bYq4795apXTrmE/lqINejpG7OBKFlgHYFSIZ/GAcsvHAYXb82edTsI
WBNZ8GgAfPGeqoVFtyVuJsBJoNP8XD94FUzi5z5HQCwLNZw38dDCJOHvDXjuKmEv
Rzb81cnR3MOJDlZXz+nvG/zxMbQ6PpTwDWgqzuFKEhdqDZXkS0sX9vETncP5CDrg
VtDJ4qxJEyP76BhVRVevNUGFXfoNKE8mnmf8SarbI5FhNRZndiG84e9l271OhpM5
aJvqSiB1Ys+j842sU8aIhUyJh/ZVBOfACxMiFREaF9iz5ip6U6mzsTMff17VSsPP
1LdsNKrAHcD3asR2/oBin1WPn/3Ve+Z5PJwPyGbYKKwtc5Pa7XtndO7YSvFeWlem
5fkCk862emnVBGxM48SbYxlUwZ6cZecI1KEIJTrAqF+0pTGksSvYocPaSahdbtXW
LhnkHnL6JXS1CgFbM+IYZOUghA/p5lO/cl2229n5JEvAwkERhhC6rOravPwlKiOU
NvQQ2pzt+7b4vrGGFeMfIMgfX0jT2MuMoQL+Y3b2JFMjr3+f6Dhbj8tuzNiG5HNn
fgByYjUgl1QOFKBa9XEeqvVuADWObndeYeL2XUmIzbGn0UxHYLUQIBsrjANBoAl3
cjdYRh+Nr+jqcHtiWfIfAdsNS1WglKIJrmCvgBJes+Q18emZAYH5nLUYzQ77AKdV
WMo0vnV6E04x/oLTtozRu6WkA9I9H44Q0OTJvS10URkcFtJsdAITUaX+Kn4vMFY8
SmvU9dmerEVgUVgkIQzA9H3QqXUI/9A9dqyr6aCrV4IzgoVsXYgrbzvuuYSJSf+3
tFOtCD0ZNxZQyyOgJVJUTsPPXSzQqeaaiJ8N+BxQ1bpDm9822nH00rcK6fXPOtvC
ne+OgIE5RHtcx6jEen/wMJyTMr+M84hb0vkHf+9pTrYWPQP3s46wWm7mWIkUoqCy
tF9jGe14mCz/5QFzXRHnhKoJBzOCbrVsHYBGoZX5YOQMufzN99MIs+Pz2y6j5mw0
Aj2JtayWkGr9rd3BT/YJV8VOlfdl6p539WGgJ98maiY+3DoN0CldBqxHWIOXR5gg
9kI2haXxbD2iFKvBby8AU73QcQiKQ4tzld0eaShE7rFQ2U/O87LhNyKATvGXWYnh
GTMvtCiq8c32MHqRdMhHt1VSezDXC5cl9i8E5AMQVELSGMIwy125TXeBvQpZVPpp
sgT5sLQMC6U6oxxxCJB2eR+QvunPS+Q83eYLkr1fl2WOU4UAr/Xl9gMcpAJ0C4Lt
C2gDpWsTUEmxwQIumltntRwPGa948RvV8OeydxH1A6XG4EMQ0cYfAJ0XAiscXqsH
GO42JhnVEsM9iebhFLU2+RFPA4/wGJUCz64SCWXuf+OQsm+R8gIlY7d0fjicWOE+
mbQTsHYSbYVB6xQMYCwYkxi0OzcVCTuO/KgKOw2TKC+gxXh0O5IygDGk3cj1BmPo
CbQy0pQSy7Q3yDP8LMj0dyyKWfcw9OyLCDEFH09YUf7XDNmoBHYft6vdMPpNjgd0
RKdxl+VttMiBYHO7sMD/unHclc6aGTbZH8mT+6XqkzqU12sHmtAvkAzFVxTKXXRF
RVpTw5Vom3ryy6usru09H5hysE3M08DK69m03Fj3aSq450MGGiIsxw+RMr2kW7PO
OANqcwIwBpGYChS0Cn1HIJXaeFXoaZrQwwT4FOLS6CdRdztvvfuZ66B8SNgg2HCW
w4BM+kMiCFD4yeG2C7tl6rLdMUZ2+6K+v9xHxCWkv2QGw+TitWhgs0rdnYtF76ES
JgND/6i+yMFSOlnR6j8WI4ysZk4+ICOSmHBiFp33co23cjNjJQu9A7frnjlZEP1t
pCYPxiJDTvvIf8wCckHMnHYwnrbyC+70nmtQmv5GhD1081kAKj3bt4PUoW0OUAo8
MTdaXl+yLwRmoKBDrEh8ogyGzxsiVtODy3EC7+pPQENAH9HmnrQeANSxlXFtLuxq
lxA04LOv9NfR1IJ8X/rFRPwY0ZgpjpvCmPAO6qVDR0OD5ilCdmq+3VsGNMf+TCeD
/qOc5WMH+gXMEIL4eRrWWtNl/16U10Vkr/vuvVLooGF9isOfJBNPjlJhI8XvLe5k
jxbh1QM5QGZ/oxwHoEI197K9zrdrf6vhU4yonP/YW6Q9aWSBs8vPU5xfnQQJypN4
NyahzaWhCnl53iHuZOI3z/lZ2LwufJFwKAOKADdxKOYV+gP/ZTruDyW5C/JAFCvS
Ett5x+OCuZ2anaqa7rMTXb5k/jusmaKbuC7KQzZwCjBoYRsl8UGkYunAhZdc+WDg
CJr15I8sDWE6R/MTbqHRTh4xqLFMTxTTsUCsjfD7Nznsl2OVtDp24QOaASKKiaZq
vFoIsdhUZgDKp8l1aYA5qzMnIoZNByb3Fm9eZh92UsvgAjPVO0goV20TNx2UzWVr
HP73IcWZBcqJgEnTw9ULtZjIJUzWSN+QI2I73rJHLFvv7WVGkNwfAaVuBbxrQsD0
lDMMY1Zm1iw5i3/uYVGKBoKqAETWXRfa8NJu7aZlRloc7XbXnXAVwCTV75N0rDi5
fa44m+Sy0YOFbd5Enj9n+Y3AAyknsLwsPgoCW7zD3Q0nyrVWqRGR8KEwN6pTb5/0
E2r65PM8T0ImeZ1BVpHNMb04raCDr9b3PzkHxWEu/kb2y1Rvi51+4Ah4ZtFXruu7
1QT/M63pZrN9vL5+FuXwMJf/b8s0AggokYvIqv9TgpV5SvkJYMNUIqhRXfTU7y2y
mkP2GHj8GpDNCXxxgz2N4J7dmzOPGM2sDf/BB6tMY9B1Ly8vhDVvRoKWQ6zr/UQy
ReZR6i+Il+IbwsmEaPanNFLMjYQL04si89V2KN0cyB0PcGP5oPBxIgxoIlGypCsH
r/LnfLDNZhySFlFPkZYL7XrPdRNIV8Ynw0dmI689koFuPCmhdxBh5RapKB0u8ibT
rFuFwo2TWztTwXdMYP8bQf1E4cTlIvFP5vMGuePbWI3Gcu9LqYHmvNHuWIIB4q89
f5pG75u0WGPvvbaq1duerjPQMDLcLjx3d29tW1rQbmcKWx3BYsXDYpBcnK0jrlYK
aSJ9ULoqpL25o5vPupZrOjHj9pIqmZolj/XBR1ATQlRW4EzwtpmNkhmAy884hUe9
mcNdDMGyompyQBIxgAhllbBZC6yrHH7FsMRkNs4Z7RZa6dfMFkP5nMeounEUBFeZ
ItKVipb+DK8OeJp87K+R2XaRFuNQ/Aw7Hls6M42vvxAJ+DdtlwJgQI4/xdCtAsfZ
BObpOJdDFjQ15OvscNdM1PtoU+UUgSjOIWIEqPujdvvjREZ3R8ONcKXUzMRf3RFM
kWxK9fVXIOil/ElFCj35vr96ueVH8pDQb0UXzKuT9foArwO62GRtxQvwF6oyDr0V
Zxi0s/nXvhrKtMymd+bk1PwLKeHBUSvinVeO0cCzkNlS2lJtQYFl72umBMoPvL5M
MiPmRqeAvIUJqQ8R6MWWG3MAqcTl95Q92uNQXrtZ3RC9/jsbBqe0pn5/bG2suyNj
64rhhUQoCP/PMrGJJZv2DyUwxqPjLPmvb/q52TrYKfukDMRnSIANGMpI4xyngyhj
zoPZvI1RotFIz/ofIn9Gz7eHIRgoNYWUg/04EN6on2QLNWZ+9dZ70AWVBkHPDk/S
k/vw+6A4pAdjZ3yRPK8qXQidximkVU+uWV/W6v/Vgp84Q95Q5idNsodf3n+Qnrle
dqk6xZ1NyridO5nLwiuJtx82qsYSyLnSwvEk3Fbk9w3Sg5EQ7+GjGlI4bvddfXA1
K6GDRPG4dnglt/rZVv6THD2SRafrDHScyEiZ8DFFCVOidhXkAL+D+1pbYEyrv1oi
+RvKiXd4i6H/MUE0NoveRAr9/LMTBG2EQeaSFUTLl9HC8dfTHJw7C6NxR81CfmFO
vkmTFdiFhkmSJSmti2rmIl0mPn+90t86drCHyw58AGhRvA+S71wXDMX8vZakqdT7
z9e5QkKHYDSkCGW8Di36VqtRmKFQCpo28Z7P0WWRvEyf0vtEZE4WoxrcbtGkoP3X
moJn2WItPw/mnvVcI6/oGjL40EGkOCvDD2NAJUd8Hv5u3yCjRjuOsnZbCSfnWRIv
8pyP09gE4YPy69gyh7B+LMlWAM7XrM8UznD8YsuyydtBZll+J2u4/t6Z9N0wm8Ln
h+Yh+w9k/FdZj1e3Q4Ue10KoALKs1FGNeON4SD0n1GKs9ymjSXwgKkllB/d6DoNt
Y4Q7TLOSwtM657UY45d0OlhvHMzk6N3n6gLwTnu7LWvpvbk+n2nAbhB+jrO82zg6
IwuMZfZC1s3Pk0BWt7tMvKMrcFQxBnu2/uqAi/FnmvtgEJoyX+upQI/dOmu0G6Eu
22eO0bgx2VmCse3zNcC66VjDDNZ4X+lOpmzkXzrx8TUms3RKE4Mf54gK/c5mDdW0
yVwj/nOJkoYSB/pZeqN/y+YB2bqV8mYdXY8QcDIFJbLyHdLnxjZRH+RnQTBkJBNw
qlAwFGqWYcfRaslIiwHRI8zWKErJlmFBBxj16ejsfldFy9y4e91ZxMrwGxZ/buUd
ZVtSTEMPuY3CRm54IygQ7Gf/OsDERKZaXizeIXLFo4tC4HFm1tAozonpLYLPGmbd
9xQAnMsGOfPYQIOpgSmsxr+wQjAwfI8eWC/WLy1gMcOB+fKVuHb93z5rZ03XksoK
mWyPbHA8dli5JK7XUyY7plPHfpu/HM2y3QD0Z+/sp5Bfk38Kc8e+ABqErfWvGxFZ
940evjlEk8KyZZXb2ZB5/E3yhU3TxzciQ3Fco3UTwIHRC0CYjEtUCXhQNaLJL9ZP
QQoAGvL4PLC2fj9b+jCnpF2RibMQnlV4dFtnFsvaqe08ppoY6JhUWPsY/g9ucIIr
mDx0nCQ3+MYErDwcg4xYSbp4S+YKUofLKBn81xTjx1iJz3SO9vqfQ+GWlmwHBs/6
0RWMk2sE5r0fKLE7m/zmwj5C1Vgzgzlx5EMlRddWGEOePkpLI5o9BgnbfL4sh3KT
JKINyPZs9qzE7XY61rgBGQE8uueg3ZZTCbCK2vPW/a29QcWV2gBH3nvN2L4bnLnr
554KX9pPyznW04RZTGCgRp5at2c6ghPtF/FcObMJKa8fN3ao2XDJ0fKxAazmzgWF
+bCDeovKWTd04ccswPjeP0Cq9zxxLUmq3IauS4CZX2NRPX7SXhrTCKDuB4N0v6Qn
KtmhiddqRkeC0AozccF6riKdj5+7lHqXwWy9QBJdIXXboNsrkyCKU73K56XN/d9X
x1AaObIBlE05af83t3YuLKxjW3cUQnIHERAhw8Cv2SfEPX9OsP/fEOplsDYkay3X
+1w4csJ9TI0zrRMVjPXW2Vd0Ur+ZacA7qoVK/3+Tqz23YPfHPWhFx6/wBC4u3FG6
0h+kxaIBzHNYEQaRwVoHO4v+Wcj1n5bN+OkAbc65nxwDxDIdHOPVxgJOvMp8veFB
0MB0A0BY5Q4Uxf5nzYZORylUZ16exJXXTFhV7Rz3YrHeRuCt7Y4aWJ0Eq45ziTeh
Mc66B5jn73+VtOdr9PHH946NQSpVXaJROO7ihkXjnqh6+qXaCdDMeaGKFY9kJnDg
T+WBa5fznt+e1/GKyKlJaue5uxNVzZbYy85Kz2FFDNnRotU9KaQF1Z9nQg4tiogE
PnAceQW/NCH+dSuPJRAQOeEQIkSN8tHm1JP1SwiI5rUiYXfmx2FR7xZM/RLtW7H6
6QNXgN5oxnNcLoegyfReYxQj0Dh8muO4E6BMQSLbSqEbl157EQzrbXY4CIMRIot6
7iTO+fHRHHTM7BGKd1fK66AoxmemkOVqRdUF7ugZaun4cbSnqKAFD2QKcuctg26B
37W8CFnYzu24gKvsmx8G+BLx/VfbZy12RGJtYCv3LJcjubZDsBjgvS0LRK4rmBV+
tRoJ9ov9k9Uo6PNagjoG62yHn2JW8cY3jjjaxg14i073tQjXi0LAA7wZ/Y19AGDO
hY48RVnZngydcOFUvZPIswDszYXCt7n82aLbc0Sy61hnzCDzmCYAJG/OfdAtyo8R
91M5uZvruesoct5jsz25HtTiHAy0cHyZKqFvUH46mqqulXT5DwljMXNWBX10c85A
irKm4Cc4t5PGUJQRqB/P+Jvq8MiDIwchAHaCvUVoOEJY0CxYigUwfa0bsCkh7Xp9
LZkooVYr0cdGf6bTNuF5N8Ha6aXPHy5wnwfG3a2Hx8sB+4nQWX0f2aZyzlInwgan
zqVh9WfLkuYPrUsbtSKHuHFekD51/22z+n1LEwUQCNf1szpqZfQxtra3M0b+T/nO
R01ByxxUFEmJ2/WRUsmzwXUoaXNLkx9zk7qwO5mEOek2qLiUEi8dGF384f2p3S1a
8iJrLbGaTivZC6ETLOxViOuTo3ATv7zd4QtbfAtMrynbVqaL5Ay5cPbqUSGl+ELp
fxQYdtcqDbCunBioUcqNMsYGxPEqNX8tyVtyN2oc42/oHnBAOjmWYqSC9dDMzMjs
mb1h0I/FqB1RT8XovLWyUPVOgfeX3eoGwgb/2EobPz3GrSgkpz73sxM5PMTgtWel
7q66YTTsf2b4UDW+4Hm65O14Bo7SxRiArsj/ZrAdbPnVhbbhYj3Q4LqdGthGb+J7
ahsWVkPcqhDnZaCJTvxoU+vntoadnSoIpqXt1eAw3dDsCkjY3laDXRwZ8dBPcZGX
PSIUeUebo1/m5gDkrHC3BBvgB0cFfqnWK4xBoW6SKKeHwCPhY5EhHV+B3M6qke8L
V8UD5cWWoxpjNpAf5JE23VRe/uUmsSrUcVnQmTl+6HlDpSLWD2nyaGgABLKnmIjK
oRd4SM3mCQobM/6w6IbnV5ltbo1GU+Bho8fe/gPOkbMKZIwsqTIsB2uj0YttLN21
Yp6DOnln+rJ8ctCMQSKyzFve2lSHhIbqRkOk3dxtz1HsnASR1f6KkwpcWcQ1J6J6
lu6Ep5gISFPYpG2QLN3j1UvmAUMyPncxfY2dKXqg+Ow9lgZAExj+/UxucRHPt/0+
KkP6KqIoktFANKRljrPs19TQeRIoPCfDvpLvL4pVdiOlDUvcfhVuKZSrc9XGgHkt
joI9uDVC/N6G+KwKiYvI2P13QdwGOshtZAwn2Su2YGAvAVi85255hdfrkZnkJtd1
fcsbx1eoE9Jmdr4txA13BmuuDy2xqwesTZjcemp0vMGLYiP7SX5whY4MPnBqskHA
8dzx/38W9fSQa8ejWyYFKxADpRkIsXdac+ujfDwiK8+lffjf9HRg6yuTvq4Mz7yN
VABjC/NoXDmphkRcZq/5lDpdRjQ4XTQMCVvRCEDbB6+rfcjQ8wFLdFdk8n4gLiGs
BikYQDGg5tSPpCbgBA9BUAGK17kaN/X3Ul1JbVSX9XenW/Figelm9g1ZHawTimLd
KyIKNQD9MIP4sSuOf21ZluJnovv+9Y4PPyL+D3ciuN7kWvJ9nUwdziimCFVRoaLw
rAvGjRw7hH8A410mHPrILrpyPZYo/Wi2qqnkXXDnPt8rhm88tMow9X9/vAI1q0uB
secuxUGMmESR6QTbp5gTTSBqPAHbLEQINp2otyvHPBT2JAqML7Mb4mQibr3y3M5c
wM7/eKNnPiT9uGkK59RJuiFtQCTcfnzvJgcDf3kspwZQDH380occWFIMDv6xD808
W/hEIecPnNwBRfhjWYPwqh3vrLJpX2PqchdHc4uwZ0aO2E9eXJgVMMJOsytbAbOZ
1x3ZIspI0ol9u1a05WGd+vYGIcDrFANld6sehMvpxkKOASWah5IAgF5yjPuE1GUA
JPQPhWk66vzC7GxAWaRU4PIb78nrTQkcjngVuA9GcSEqmckd+c1BG8UUpx4z2QZE
T5sU7Ije60/sjaIURIBgZlj6JzGkJcukYa05kuXYkd6w/IOon93bbuSncTN0TPj8
S4aehIemOthbGGXRfN0wy1yks9dVJP9AsU2MuuzsfIrggADuiHdnsVS7oCiRL3FE
NuhInT7/PLeDRkob8moL1cgSRLAsNO1qQJhBU0D1FZDl4wNCT/sAS85xpx/s7cNa
wTMFSkJ/WjW0gvU5HrhA3V8Y5lh8dbNa400J1+AvkzMN1fR9TrOAdGoZ4sk61uwN
gMVqN5V1ctpcx+E0E5K8W1+iOYa3gWYwDjr5xeQiAsaATdE/WDH6rmC57AOx6M26
XJnlrUADf5ssoEaHEgR/3r4rqxxODCb0XpFkbRUZdKtqhrQ4OwnfvrcDu1OYk4KI
1CNK/NhaBC0Eypr7LbP5lbMV9CzzJyWoSfM3WBYKuVcbNVlOQD+XP6dHjQ1CKfnQ
l0bsQSTch07W2W+5WHHAoxiVCwLej6RWJwkwxz/SfkXWHONVJIRIePkvf1VlMHI+
n6z+N+n3DB3I2uMZKIgePv19Bfc9HofuhNsLScGKKSVZ2QgCZ3aK3twrXIAhUnTp
/CXYfpCptjCQFIOUSed8JzahfUrX+77clEd+R4WzhkggFf2zyD1NJVx/ihkhVmXp
sz0SndtbaNEXphY66s5z22TE40vPulHfvfr7NB2z9LKHvpVhAsYJP61xPD+1eTYj
VOXPlTZoSQRyCfbvheWavy1OnkiHZKv7v/JvsgcZb+GU2dLsdpC8Z+MAaTJazb8w
EnuIKvII9XaQBZAR1uU4peBu8tzZckTswjmDzJCqMOM6BrA6g1LFIqooWtNfO2eu
uwvRiWYIcB8qNud3p5kpGoMLLfdcU66+Ec9QMbeUFO/MPwt5dfaruNObRN+DoeaX
DLmxFrmxoeevuKK8RuwU7B4I9nI/jwvhb8vugoviwlxiwG9uybm+AYw3VTeFf979
B4ks4fJFuxcyu/vcqpyXlse6h6HfsSiMYZooIHK2wKzb9G4e5CRu6S83EgK8rrqR
zoFPiUUVPv0CkzBSS9svTEBfTJ7Q6GCtpoSbD82Rq+78/lK0+/RbE1uhv0WvMIn0
K6N7XF2g7MNIcwmB1HIKbrG1KZmLSVI8UcaRiTk98+DUCWe8od1mh4wYUuhkFBcL
9FfPUsCUiSsJ6g7kJ+OX9/x9LsK6NLUvCrBtJ7y3KkNoSsKj9caUHhZOSqDAAO7s
3zjV5PmDDSi/l3h+C8YJP5LrmiON/fG+/g+9w5aY7hKXv5mJ3Fi2rWgPujHoOYiw
ZW+WCnDBfQDX2aHpSh83j+vva+uW57UeYvVEHmilqU1QDB3tYAdr7foW35pSzVHh
vEp1/EPnRmUI8oR4YCOx0UPP0IdfPP4n8afMURyCoKvAo3xOIlLpVuIWMWlEEk6+
Nm3QrtHRSqWGjO9qE27s/Nmsu+FOFqOFINncTCHxzRhi92RBhxsDR+MPt3XWn4y6
HTbQqcVhcu9w8EOJE/q1ypqJ+koJAMEN5nE4ToC9cHoz3C+/QdG0dRg5/DpFyUui
m2lyzzC1LGm/qup6XRwhJMM4sk0Qncqz0xaD7zjUHvdkKjwZikfwA7dNh+H9rpaI
PGUQZOLhPlFX8bODCOyB4fDS40M+j2KrtWAEKF9FaSsoVsVPO78ROLjeRIWrAgEU
I3MAy1WCv48YeU7yu56q6ZCAlHcPOgjSTlGhzhzDOGONfAe0LYzTReGDM//Zkw1h
xZa6XG9mCfjtpRoinTe9WzJBvFlVV+z40HrhZCt7eHGg94YtkEEw26qv45TCRi/t
W++RXIWd+aynrB7uac1TWMP0LtclMH90HFUqJgnXDTJqz6ljwB2L1ewuVp5TYeuu
zMbqYl1/XYfNDg3jM/EWj9i3GOYbpx7CS5tCcrqUPYNntDG8SlgMMPPql4AM9sGM
eOMAca+LiBf5kwzQwYu15Z3mcTc0m5iSsJyFDHpOefOFJW9gW68MWUs2c5fgXymB
KcXiqLRdFGPUg45JKWJ4J/Sg3JLxymWSNQp5mPfJzsnb0kI7DQtY4VSCUca36LnM
TsLTfjxovxmdoxDB6SE/6Qqo7+oVdD81opP+sIuLUyQen+olffW80/jBCkcZgxj+
xj2RDPelWNZvB8PdhOoZvL2bTpjNQ3exNBBVW3BtsbVzz/ruTGzWl5U7pQOAh0VP
de1uyEi4Lvgoloylfdumz8JyC6tgUE2FIopOthu5HQ0dmOSpPByAk23SKo7fpj/G
SZn6DcRyt7ECXhoF3uus4ggOvbjFG5/5ywLAVfNZ9mtsww+KCfBcNwZHLOvWnidc
PibqGsK3XmW5EM3eCKYgHFZqhCFNDZvSOrR0VBIS36c9SEIa37Ch3Gj7pdBqC3As
nb4+rgvROFsgilwMkggcRmyBGeWvZ12+/ev24VixHo6fvuZMnVUp2dH2plX3GgKP
0CbzmDS7xaBlYCtIopQSoC5ESyNELyrV2KTgtD6RWI1BhpC9zKZXV1cFYG2Dnt3h
1oVX6tFjJcEbA2uekdvKr+ROQucX0ZrSMvKco753NY2C3+3gfJwBUGheLk90riFx
cPpTbpZHF1lkqABn7ZS6dvnY7Nk5WIPPwTVffMNOdkbd47sAOTpSZOPPbHAR7whs
QnsGm6YJa1g0inR2CjWYbeejna4r49TvV6O7X0u8yoHgwWl+Ap4gk9Eneet/eF0J
20tOXdCzP6T5JwxTwOM0NcHsrG/aVyJ7HW3DsUGkWR04HhGM+ruMys70YtSOqELN
8g0010SuWI6gGpuic7BSM00CuJn0klAyX8lh5NRIn3uE1kJgTuf7IFpAgUcMxNA4
AtMsX1x8Kz0BAhYVMJoh6X1UDccYL3X3mUcEOsVqhiSUaw/aBu1hM72RuS7d4cn+
3ZanYZ+ajqTZUuQGirTGzPotaxXuKGolxLJOByZi//U4HxzQ+DAMF2BH++jtKIQe
uRLsf21EZtIdy/0z1H7n6eyGH7C5I+vCDFavtaA7rTuA5+JyvXDGRGtIPwh3JtEX
EMx2XWZv2/E9iHWQfoMWumeZwb6Hr+dQaI52p0asgnUcEJasdSMD7Bt95pe77H4s
rlpBr9vAJ6k7ikQCvTGfcAWGQqcJ1TVcy2t8UNomksSq0IehBaeOFykVPGm8W1os
EWsMFGsv8nHFcUpYqVtcrEimNcn6hVK7T32j9H3jfAvy4wgpt/mSfqq451f7fCfp
t2QokdWc3R3Pl2hDrJaVKItMmYJXmrR8AUPbyBO1okQPnwt/LR0P2v+ZJWt7YlLl
7kIsUpoFNnclCsTh6fDIAMUgW/JxiGZk6gpTlBPFQnu9Ye4IGAVyLBW1U5QXM4T7
m5mZQb+MJZ+ykBriZSgFOk3pMUYKeRkZbsBaJcBAFB+UzzF1wIEibBSGrBGBq6BV
sXxXRSfvRSHsr7azVT+yMnDh2+E60fKKXrV8xSTv3iswANDFtLSOC+Dpa5lBzdri
da/ADIbWOrLU5if+ckXgSoUN7kHlBPMacGUmeGKr0tHFwrwJd46qg+9paJK+EEYo
MR+mOZay0VCZJonnQUBSgeXvyzSi4neYoGIzY3MAkMVPOn1Ops0AAhhfkAKeHWpd
m0Qiq+oS/jCkeuz826AI5QfHXOUPonUpxlyqB2cpIx6YoJtz6UskCqQwFlaK2GaR
mq6S8Eb6pY/g0/wwgQUCjcpY5RRVfmEnpBXjG1hJEW6LCoLy6PKa5HRyIIOLNen9
dQd4Q03FzhCZR+AgfdaqqGIZOD4yTYeESkf2ugmBP6+dNXkYTyhC4G2R5y0SD5Qo
XRr46RPRYlnjsy43GhuuGkKfMS+WW+jO/In4PZ6HGoyIV2sSHiuho47PxEBIM0c9
qpw4m77/gpOWZIc0iRQ0lVvGqcOqZIz8j2cFp3YSrgE7NiVZMk+LDOdizhgNO632
VJ7mwVELHoYVD7yUcSZhVzjM17N3xGX822ph+OHNor29TbqEULRAFXEVNdxdRC9/
9Phaes7+EaWIuz4PwJ68m5SQvS8guDLf/8V7Jm1a54CDOKvftBLo8e7ctFUNKFes
pVtJXTYaTn2tUlSHLhZ77UMXTXLI/qpCv2w6yWpHycSQTdsjirzmAZ+BQtddOycf
e5IErvE549CkmILryZGxsJTKCMpQbEN//6uqkwMxhh5EiuPvOzHudhebEHq/GWq9
FbJnL0ZRQ7jMYwHkVXovAlKQQFph53RoPKH5+jAQbBwgS3xFj47um2VnopOl/hYA
lbcXFE+MIZnD2Yd2NB95xNgr0lFF4+jX9GdHaj7lxDEhi36P5w/4sO68r1/L4BKS
OSXHppc8iasJiGLU94UE647ATkQSQfYARRRNq15DiSDv5NhG+hmZ0HqY5VNWDQZE
s8gp5EAk7Mi3z6pTABGGTRrh8WmqaZXjhopuNceCxwLAxRENP1Jq/CIVmWg227Q3
3AHJt9P87FBT4uQa+sHfdkvpiT8jx+EmdOwmllDaYjqFL/Q76SRckP4ByGHdbUlo
xkSj880hCIjZSL+Kq9WAwYhIQrJVCEF+evRqU2YwQaMZH/bIiti1vT2GXK1LnqsH
X0jU5kqs/wGjKu4OQo938qjp7DlTnBSnH3ZIWMzIfABb05Nn142QLS6sAVl5CC1S
NIzC/1/wPzufM0B09YjFxJt/ZCJbmUJmUpQTNeoUEcwV7PL8aIZCLgOo6dcIy9K0
G2EBXIPz68xxzWnkx+iyMMvk4tD7KmeouDaNh/m0FrPhBu72t3R5LuOTMQW2Dta3
AksOygfhOLS8OK9An1s2rhFflbrxp7zIi0srdR/1lZl4p0JD2cpbCg/64wR5UMCx
j0VBBnH7PsQqDkjZ234OSKqzb+WY9xFkOT1+XHiPCz0JUtZtsDtzBgQ2lBVP5AMk
AgqtcboAzPjzv8mS33V9KyJwymmhrTJwshRpBGLE3NCd6GjNzYL2CbmjUf78jHxw
myD03jhFihtSGkRyNjapR+X1UtzqQ7sWPohodScLhDW9OrLc13TYreOVbKIXoIKw
kxqrOI2YKRHJOiMbxywkk+sdirXXZ0lsaVs2GiNE3qg70XTimKByN1fKXTj7u7HU
Og3BqnDF88E23RKu6I375UM18c2Ctzt49qZXdBUWN4N/xToeQwH+VNOrFvCufvYm
zOnmH2krHnbQMcWwrN7e3y8REYmiP0UnrCWUoNDQc7dRIYTzoHke4BJBnSt8d415
/O/M6+AQB6TchUDa+QtaQ8dAyza+MF7cLoTmeg3kiTvBWzgZzSrOnTS631IatW/S
PVTj0kGucWPI4+85sPi9MPNE0BkBqcoDHeYS4eHl0FiL28/S/FhIeyJ70OZw7Ynp
z4foGJEgz9kIZqMpF2Y/DAbcOFmxd2rpSnClaj7Cyzl36mfmwm6UesRAYGtI5THa
WIGHrVQOQRACB8UORI4nQi9q2f81N3s1y/AeqMZJLMAwrIRl/nhqUnlHZxH0psWX
EKPr6UaH0KvW886xwLGyjxPQgZeBBCxkkdUisjob5sjOkaLhfp61NIgMr5/UuvmQ
SzjG3oIb9g7P3ZEQHgUCZNef3TrzHdNl33vFkf6B+68Xs1Zy2LwS7Dx7zRzRZJ/q
cMeuHjQgpbpm+Y9/rQI9g64WQyn4Zr9AQXvNE+SiO8S2wU1xdRvbvCqUlvOMtZOD
oyoJTvlTcCNFoBKHbtcnmsHtVFcDqDREeGDn9v5oB7aKlkrZgn9rKpGYPZOJCN9h
N5kNFZ0xV8g7FKaZfjYxjSofnTZiuRrL3WTpPsAO5jeN8Cww7g8bFbA1WPWcm8E3
xAgZfNkLIlEvAg873O4bUp+tMnB2h6FdUHd+wyL9XuPOmI4JMDkh3/FsMJPyKY6m
ymD2TNczKa2aNuuWqyObl4r566ZrT2KHnd9dkcB/327eT1Hl/vKn/XX61Mn3E3j8
sC6VwMJ1z2y5UCncHQcW38UD1IceEeijGYFqeYaCtr0TATwdxqftdZOCbdUOpz4g
QHgNmJ8iLWmz0cnkz4lV43NBsgyzGRy9I6jWidVBQf2/iUYp/uPOmsWwr/80Iygn
YMIw+sH/wy7yJhFvpXf1HEzjlqOE5i7q1wydnxo/RgWb7WjAJBMjd14dEmdEdWw4
arUVUspn9seM9Tn93H/xyFKQ5HolHWJds51MGTVHoV/eHMxeSmCY13AsSly7oFDY
jbWG9T1kzd62ISb0EGr6dTpbTmrCxs9D4Dc5USPAgFHzoRM44iIfwzkbawCBER1r
h+9qcdBrqX9T1aeDWsez4BKyWCBFY2u3WFNJNg1szppljGHKoXx2AYwMiHhsrQQd
D3Bf8D8B14zi/BTV2jtex95GUmR0UZHDM4cb/ictHm0buCIl5XfVybfJNX4Udp/o
5Vuq0exdfiTs+dIT6jzDdW8uLjsy4eYXLP1ajO1C7GccTCql8NkJ264+PUwwEtoA
WJb9772G25NBMtzQWMJE9Mbjln4l7K1TRy4F6AYpLYlC/3GF97aNhVrZbjMWl5I3
VoYDnTFNMjvyzzZgtWMJGXGQ+F/yFihQ3Omr2FpKtBsORtOAkcdaW/6292H/AY+m
+XGQ/KjyL8OpvBCGVHOjFqS8AHsA3cZbo63CdA2zUveF4i9THoMPK9Rx2t0AZ7Wg
NL0gcdVhjAXDKM03oazqSOYnesD3zdEum/jOZg1uJNM2j263gQSLM8D3P/mOqabA
O98zWhxqHT+UzR8EQ4fMOYZUnBikczBS3evQvzkYZ5G8RSUXCx9I1g+T+peS54nc
fKFYFH8mXk9I9S3FIzBISGRjMUzn92Dn5vUhK7zi52zJ3AgH5rLQiRtpJK5Vs1iL
eXlimkVMFQWYZZZt971nCkmD7fZ01QLdBN5XbBiEURhoNQATJxGJvUM2rizhaliY
/dj/qWLnIgvfIzIWEj91tsIBYiol2WchG8rYdm7f7rFBthtBZfgUCEPHPf46EG1A
AisWDRA+LskbAjUzZ3IUsJBblSm3IucnQt2yqipGM8xlV6DdXRNW7daIG1rNxz2d
Lyfvp0C19MLRFbnELdGebv1v5+wnVSWWpfsRFlYsilYuSirvkMEqCQCbXdE6/wni
3hu57isVjNZO7RY8me1lyC2/2062Fg8WV7xmJOyfeoCZmQe78opvPqJ5DsmbsYAE
1zc1Z85fT1QbcMmZXjAcn7c66+arR+cbY68MRx2sStVNYYSjGleV4XV2bO9NCiFg
+prdu5TXYYszXsBBzY+1zSu2dd/401SZYl1Fg2BceRgH+wL/FsWbmVkNr+GxaDcN
TdKfNYOVhuXOLRhWryiW2vFlDO0Vh538pYzZC6S8aGu+hv2aTcunyuyKbbzfAcny
E4M1INAEPvaCbhabjvXC2UTxqdq4HpSwcjJ30KRU5JRoWmYGZRwU+A6Z96TETKBa
x1zB2CAJALnfQBAtvYyVITk35DWkitiC3u6f63AdvTtLy8ptPsrOFis7i9fjDrL/
gQt0PHxJQj3gIeKECatcxfcxC1sLMGuFfKvnbPblvAcHh4N3MTIDlsrYn1P+Gw7A
FfubxmglsYvm8xncOs8Z4LYqbxfbrsFd+iVESGSsDcJVZT+aFKqgsgnvOVmTDNpF
mgvb27nKUWloUvqa/W+F5wkn03KhIu8Fog67UlTlN/+Q6AFei2nuAmDy7emmd2fi
BPJCHUEf3QnKPwrR5UkaEUwiweCVrW2X/2M8ersyfgekNVb8kLlEwvgRv9Tnfwig
7bEVT3/U15OMZo31CUMFVHiqKj6d2QEtlYM/dFUtIDxQINBLddL3vLexb4cO15cz
p8eB8JExXQLETqtS1ZG+IVamu955p8q39UhUY5RczqzQ9hcLHRD7gTa+62E32M7b
c+3+CrnXg3y0LZ6RacFUVyH5pgQYnJwX0oFfisJlxz5qjaYKjvf3eI6PEvRMxGkL
Pe6H5/r4oqi/w2z+JqUeskF96dIdFvJEePRgt4abgWd7lHXdntHeryRpnxjiGLxY
CAGhyXYgIDkjpCMGl+1HGq5YnEVQQeU9Skzbl0/vTLkYiyrWl7NXm+CEpTiVn2Gg
5ggYXGIldr1wH8ivYPUqSpvoxOWpltPyTO7ITnVjuqk9lew4y7Z6y2oLQMep3Y6P
qsrxBxuC+oaxVDqysPut9o0+Bcms+9E5NOJbbjDYWAexdmWXHzmBdBDG08GXqcSY
1lueoRZFOXWHiJPkA+YuoK+5KvMNUcJapmz2eh6gFv7FtW9pUWrODy20f8iouK4g
xMrno0FIU1KAqVg6cmQWph/Ns/siPQtgu5wDbqsgjLDJEJtxh74grn3rBgsf4d7R
po1YK7iNtGh2ppG7m11Otb6/XapKMegt9aTU+BNZcDbY/M+YMOELu4a+KO3grAzQ
EYg8Xu3CVF9GJNmy/cU7p0rcrCYoqdDSdgyse50ffJFckg0Zk0jypyX85bHjUsSF
K4MvRS1EWuHrIIEzUGjHxoeGR6XUI/bdnHB9FcaiApJP5DfEfkwBvjqv0txvb2JM
D+Gy2/fP66zX8FCQ77h80bjYP6nNUdgrEXZns8NReTa3M8mDdvDftypRy5wL+iDZ
/KHyQ5CXhBoU7cQ60jtMGL0XaZssd/qV0/gdQ7WoaD/Vl0+jb8XLIvj+QX3dls1E
96j1JMb/TjGfG1RO3lRlTTzziYwuUbhD23WFg5P1+gR/Az3MGuVDCJ3FLHJpC6uV
XfGBze7aDLZSx4kFuYl+Y/dJJsL0XKC4A8bZKIxR0AeV0D4nGVCJrsQ0SSrpAQC4
/RErpr/1ZlthBjh1qFsHXDFtWu8A3GATBv7nHPKJKV0RlAWJFXo05JI4Pnp0pOwD
e2Mf1GygB8l+KgL1mZJXjer09aIimtHm310ruHBI8ePB6uwwvR5n3j0yeocVwAKg
+brCZJPu3fvj1Eioch2Erez9Ua1BKBj9/MneTDR+jaRsWorqZqWgE6FNNZI0D0B+
52oDwQaNHb+aHUUAiznjsyMClp4iVdVyKlfkY78e6cvaa676lcYqyCF7ml/dFiFM
AVHMv3kzDCMqYFJ2wTdxm2mw6NhxwPiFKEfeUtho2RMZ0sq0rK56b9+mcVwBajA4
zfY82v6w1xd/P4NgLWlK2VLkApG0VpTGbh0S5kXUawe0ikjItUaqmk15Gb37x7J9
TsfLKHX9o2RrWRLb6v6I02/iaNFOymYF1uTMX5UMxHZWXhCztAZUbipSgn9Ysmpk
2YA+EYAv1W5XrxJYBTnVyMGRsY2mkoFcVqk80R5bll7L7DP/CRNd9PKI++uwvZ4C
ny0lMMKkOle+H1Z+XCACghgCyzagwpYegBOU8Ph38gF/c3ha9NcZ4RtSY3OXyrus
7wVtWBE3uagcHqsY882jbvdvh3hw/2O+hmd/x7bs6VKZdbaHyeQ2CXCii8L0D0Op
LQviUICEKvJ8ereiVCWWPfnY1uo62NyX65OAa9pms7//6+JzG9GXvCKRhDJ8QEZ2
VS3CyT4TQGuxiDhDPQE6zicmSsrW4VKxZHirCQ580L2Cws1CC9z/UzZc4+sEaTCi
xQHteOX9UY9tX0fqejeqidO7ahiGEBKp4zY0R5WGUvTNeuRmv7OLj/6EW/NlQP3R
MhNQoXr20nmlG2CiEdRw+muqsh+o3TpOaYtlktUyQOljMwNhwwkm9xTIIz8DJZwQ
Irf+DmyzlIucM8lz4RVxGEHvZhJYrT/ygOg6LthFK0SUwDKHadjlSkzzZ2rWTyFY
cglGKZevJRHYMq71glFu60Xk66F2OmKanmKVn7N+Va6ijWpYA9AKSmPMD+rko9Z2
MFrWtf3juwJ9bvkkjRz35u0DyzqX9XTJhg1pBsqaiwMwHqtLmn225ov2AeftKZ9E
3Rn5nN4yPBTl3t+Lv3qPsQylXalPSWl+tAUzv2WWqwb/9+C0gn4zuVp8XNEB5bHv
0JHkqoEi5UZw4FP4CgGLxM5wGs0Gu2g3vybDhTweQGv9B9n3dSyUZ7f34QmV1joU
/dynSm1d61FefXR3HI1jwFZQZKWm3ysgqo+Rcb0/CiwbiPKoWiLklmm1NhxmxgZF
qLUY1d9rZ4brBuzW9uVu1wAXJooVPJMfXnCM0b3+wSVKi88gTBvpxwpoPoiyhFJk
ecPNOMM5lUOEsCPKidVs+JLgjzSRUdE4CIvb4MgGCtFT94jD7oGO5OfOAJj0yTUT
QSggBWtE8RXvM8ZW4FFUj0vcFyBReqAtA6BdNWoMM5Xc2cw0sQZU4MtP69yYw+7J
hPcP4lr8ACnwZm7bZVQPFXw/3a6a16MMhpRkHSEdIFpDpdOAAz3vC2eu5Oucfe3w
CJeAOsdEjSSynq/aXWhpOl5kqBOHtuRtbbFzEMEcnechrecmk9WLVii7dewTpFeN
WOxboo3c5fHiE5+OVvwVYkGd55C/HMSUoW0+smypmxFr7foxJBx6fkY2frwkQfIP
R76P3YI/0AYALOK4HoMHrgA18f6is8dd43ze2SJ7bykkh+UwUYNgFCfB30qqOLfb
hXtvUXjx8365qwt038m2M8IyASiIQiSPIs75NIGZUfub3/MiMTi7V4wh6GVZ4m77
EpXMykcEYfIWRJ3pACfxWuQeZNot1vsnI13EU1RbAhWqhF36ljq5rcGpQPP3sgwb
DhIk+M9qpSteAA66u/OpivIh1dp2mQTpVLDOAlmjDui8n4GtKtz+simhIik0GCy0
0ApasRN1CuJdlahHdC5VCbrzyneujMTbr+2hAzuybB6VKGNWag0ALvZPvue9ksgd
ndHVwFcXz4Oumd4aXyBEJWmY+IyludXgu+0nVBcBoC60SjE/8/dypYbAlXt8gGvy
CiZxS9g46OkJhi9A2IPXMHYUSVDcnOcpAOTH+IxAr/Ke9Pp3jlTsE73hZm6aUAqm
N6S93SoMEoTdjenYD/VBlWk4DcgDO0HwU/vCtQkqlJQJgLDRjltEI6N8v78n0no1
8vdWwO5bwEg7klMgsfQ4y2CnabP5kpgB8dXT82scvRgvUobx0avShfKVYSIQax97
YszpVq/DMD/AAV1Lh4E2Zkp2j6z7w/QeflsPSvyFhxdkN08B8Y2JTaQndQ2elg5+
BjawcEUzuqzA119hPF30zkZ7xB7EpMUWlO2g7ipdh5X6ngRoW6k8SPHH/tNJ32fk
rHYLgMkVpeCQ4F5A4EyybzcMq6quJNju57MqZUOVp5R6hGZpnz4VXMbUYTPxZBnk
7FHYJO559JJT0n7nr2JIfdv0Fsx7kzou7ErWe5BX4ENU/QRMf5nZoKdBDeCroMNU
Gbyopo6OhDDtMRuOitwQn50YqmGdoQEdLbgS6Czd7GbEKXli23eYd42h1S4blSsH
zzlA3w0gNzlgg0XC8exzKU0aJWZlbWBEvozLJ51gqM7JNZXFxZlGdTQ7eCZOHEuY
FQLw0Bd857JkD+UxKaGh1r5LyXJ+4iD3WgziJ5Uw6sjuPT0E8MqPJwCVOGOMa+20
jXTD1z7sTLA7VSt4nvShzCvTHvVWHISSGS31lYrGUn+E30OoCnJW0aZiiNFeSrCt
9xVQa9EU+3iQ6KHZI6AAW2FHh3gK2sObhln4Tm9SRxqv4WmN1ktSrwZWQ9Sy5JHk
5K1dCjjP31Ymook+d2U6+YSNgP4QfYdAiWgWnhyyxMpiP/OZunhBG3ig6h2++wzO
g6EpMx5UlhQy620xV6idqwMtO/BkZwlVG66/GCsZoYrvA1xkcNCTQDCbwiO2zy4S
1YzhZv5qb3uTpWYfiUs598eLuZOOnvx3MWvFTdEvi99blofynYV0uHKK8t69bHCy
+gs+oOj9gnqdCVL+6RfhwZRQ002xWMVp0fQPiDL0w2c4CHAN+H454W5IK7pG0tK9
lN9noCZZE7buS4jz+HVS6dwl6vfR/yHl3/Tit35xBNcFN+4fHVRfMiqOGCf0Yh+i
SVMgI6NKwrn7TKe6OU0Ys/gqv2xyksBCBk6CykZ5Am0V3yX6v3THT7aKaPo6cJdR
3rCsf0n2PjCH+uADLC32O+HSEnpIghAA1wffAlT57C6R7+UwydwBog79uX5E9aTQ
rcm3d508S/OsY46Kf0yfi5OGID9uWxV4duOMOD3P0qtuGy+M6lvW1cHsf95HwGNq
+OgBKwdTa85cfNHRnl9e9lRmZ84FxTS97a+aEY0pPpoD9pqG7cEGZl98UsuDD79h
7NRzodDwB0RWVZnoBoVEKLY5I7S08ydW3lgqjp49qO18JYI5GQ2IzH0ua59OQ96U
K0loyApFpdoN1RtzSDAN5yKjzu39l3WTaDclWWp5nBKMUk+Lgfmptgw8wn9IOvwj
FeEOKZFo/jhNbdzFBZksT18dY7DV3xyGq79Fx9pYT0Lg7FYoXhYWpnMat9WFrD9z
XIyJiHd7louWFjVEmTVUoA9mULehHHVvWnWDeWniuZ9ZdKT3HdYnQzeB7cDLB6ma
cknTQgwO1lHtr4cytPb52OPLfCwv5Ncsy8PvPZlmFDqMbaqVOHTKvVr1z1gMpK0i
v+D0igLiRCsZvj7QNq5lKF3wOATPKEffYQHCJzohcfRtjt3/6ixsYn2jxlMOjOhu
/PVxDTPQ7d3nUHLv5m1WklFH7NZyDmT0ykhl9dBePosUbmF0XqAoWQe1y+VgMmKN
cjh1tHFXE0zzWmR4xHpK9h83rV1avpRQvr6mkjlV1OC4owQi1OA/fKX0aSkx3WP6
KEMIydFKqWhP9OwjaLs8A9lLbiZYxpYcj2VTnj4KPoyKepp4pkCWkhAWjpF95cVf
ivRDvAQxi5TWeglc8IQalGAPMLPA6n22pJfvc2hMCrfDfzOYiPuiu9zs46p8gQHd
pdMDzYWEs4DoFxO1UhhFXwIBessyRadClCvUgw8bnc3heOOmEsLL74t3p03LHTNW
nnqK4Des3Xccwc737LrnU6Rv5YHSFGJZSEWdQHmGvOP/PdQd9BOU+HZqvlkkSQg/
jTOzTKTSFWoHfaW9UVNiiDZLe2rL2hq5C6rdbeIBpvk8D/7a38E2QX6/wJjuuKL9
8vx9nOSrbTGvBulgPLkyK3kB1esRjS8nmT94jm7LRxCTnV75R+63xAbrv6PK63oa
ix1pdxzYAsy3bxEdS8jL1XOXwJWAI1OEH8Y0PZYes1hV6UKl5vLBJ/0KosXecwfw
J0DzB7lHSy4+81HsGtXoI+ltTm8kpAz+KbqOrSCZVXCRCzm/dCqpCtTLST1R5brW
tuSg+fTmENwFN/kGMcSWDY56MLJF2D4bGPoJ0u5ztF+0sAdakcEH/UuZJ0ZMW4Dc
m3OpnDl/q7fL8ewuNDqTapbIJfzWqXndrOLaEVOExCo2MUxjevw0McjahoUSaETa
gA7KF/vkWKFJpMsHPQaAW7uXylSMGfoeyeKGfZiRdpRns7yqiWllZU/GGzfZFpL+
8LVlBqdKRLEvzskQpIHKRtzIh/UYrgUG8HEN8yNmXcbecdvqu5mfNrXQr9U9+YVy
K24kJ+Zpwgq27LN3pIIhEG3ZZekoPtGj95yy/iFIx9AOICa3BALO7XYyMxOSId/2
p014bODMc5T74BO/vv0DrR4NglGeuQpZYwpVOLeUxV3gX7XUl71w9jzRT/WCks5a
z6FCW3KI6V8qUEsuNBB5cDfQSYl7vjPFL+4NdS8RnzsTdXxbUbgc7Qvk/hpd8Udm
Gbs/Dejlv2G/zuhF5tNYztfqLiuFGlruYYc8i6LA04MHtCmTFMus0c+gilMyuDbF
O/zFK5xB8wY+F8XMDf9uKzspzQltc4ZVjJng6rQBOY6ZoLSam2qwyeCB0UP2PvuB
3tbCLAzIOKIX8LFPKOji+1TfudCUCbP3f66pE1VjhlgZWMfxyZeM7c+VbwImsUc1
IcyoFL/9VC7mZB9IUZ5QZQGQuT8KFOFqZqbgI0DXH+QaTfmJXtg5kL6u8xSpiNYs
7jyAcBE7Py89E6CtmbRTrw+HheFMzS/EOZWvIRIs1wdMvbe5GRfcWTxXqQQUaKJD
VCU2kSkscvFEt3/fVDg0W26aUU0HPYDDMtctMgn26xQhwI+IDs/u5ch3fnYmUR0S
dfAebuzAMmI0oL2aAJm+/IKbksTtliMNLVvXP2sJ8xBv5CYiGkPUd/qOHWBSBocL
EcpjNRPhHpofOoXF2Hxuww6MdXreqyUhkiQq4d/KjsL4ir8V1XQk54XGRWFW76WU
VdyEf+71CJxy/2QcwT2iUPmcJInuOjFi7clsY2M9tuEia87yVvme+txQJ0rsMYLN
AO14HbsRAstwzdhjCUdsIcBeEuZODh1WjFcGxKf+qY+bRTtrajqU4J4Fy9XHXGOM
5qEhVNfqZMmZ/SedFB+LcIFEYJcKtDSCU8C2QeDwaTlpHN2wyQOA933JPrySI0wn
VExSkMTvERB2TAwoZMlxoT+0017I1367IEmByfBs72Rv71i23v1bTFCELHmAmggI
J2SSn6F2lFm57WY/ZdlNHbUHuFM1e0iI/99p7tOBbkyoT+uCMTfoTks5ysZYldyW
e3cKQdxf7fpcUm32ACQQ5JbCHWvsJos0HckQ8CoItl/AQ7r5bG+IjxiqKEI54elv
6Ho1n8yLI1CWfgTO1wNBvBRzT9gW3hYhCczy+xZWxw0rx+mCAMu2jCoiLB7DNeTq
DhawljSaH2i0p+7DYovrozzaFe68l4Vcu7EXC/EQ1eKy2Ls/tQQ/NQ6l6yM+HDXS
WfvRwM+/fIrdNRx2jBmNxqQOfnCyyQer+JPfyolGb7qzNBYDvZyjmflNUMSOuGr2
yt3nf2UChChZu9ov/3iPR9518qdL+w8SDeNIbkUe81HYHvwfyvoT3MhYmhHnSyWt
ApYkorpsD/FsDfPpfu048kjrUHezs4nncpwnDeY6TDM0Vdp/WfsvJyaujzB+5YuF
t7F54N6uomcCZ11INDQxb+4PmN8/uKLchZPGBOHuqb6tEmLuuYDNbYZ3lNI6hckb
Ir4Vlm+qVESh5Fxe0o0D80txTthEBIwb9R3hXvwXsm+ACL+jlWv7Mw1Hwl2j3anp
9y3+8FLGlMapcZzl7BynEPsOyBxPSXkX0d02VjbxmZarcborNiUDcMjximriYZwS
gjZ3makOk6X3oQh8DQJSEAJYdq8FmA+5vyYOBmOAk1Hd57m4QPnEPezscH24M/Qs
cW5V7MgbHTjiHV6Xa2pPhASzw6eBv3PMKASpa+hhtOm0/NODli9PYlVb6+s1Ivkm
8Bu6Ri01w3Yu11wbvzgU28bWW8Eh86QTT7wPLMZsmzXRl4KmoYnpwuiLnho01BS1
8kILhRTvPKT3MqOu1j9VPLMKpSkd/ZKC5fiPT576UZ/PD8kPJLFG/3cjxZIb6W/e
CD+b59iG1a4xKcEk2E1fTX1XJcTP+peln/SIfHdp0hIw8cEW2KliLE60UqXwIwMg
KVckvVtmfEOZhsBtbzOw57Thl0Fdu2qASRnkSBEkLnFJLv6VR9T7roXR65AJkcix
Cbe+cx7/OF/gCZSmJjpmm5fLyKKZODMAc0TzHuQQG32rQ9uClY1eKeJOdxJRDzvN
Uq+n5HalE7kbnIy+xiDAgLyXnjvK+n9QYM93pETTMAzAHKy+erHP6bDTU7WlBvXP
9XBO/gezHG3+NK7pG5zu6WPMmVBl7GviRC4pRJT9gTuLUzvwtOyB5epwVa0l+wJt
MgxG4HNorCn8FfVFFQWqOXxHmeWBLPOKkTsJOcdFyFgOuInvHyArPf6IznXjWK0A
pIVhBD1of9Gg4ixvlREy9LiibVDpq4Xtvw5dSoP6qXdU8DQFRnKz2bFNRtSoxDrt
xxOP5p5rrG3/97cjsC7ITG0kUEOMb1rZqt0TqkMAa1ZC8mwtvsrwf5eox+t/ist/
Cv2NtWUWMHrzo8goMnAkpqvLuqL9DxLRMK3FHzXe/VB2iym2XoRAwOTM+flG1gnZ
p6AdUcFnRfYSGGL2NzI0xSr2hQOke6Qsy9KBzvi7y6STtW8iN0JtnKmwSZttI5p0
IDVMg+mi7rjRDxDdCidH8M5yx/4/iHMyQDgdnJeZ6G9trKI1Iqmtq1fbL0PzXIcJ
yEd5xlQuMaqhQ81dHUNMlRHwc97ysH4TP0gEZ+2wjePOHIfbKeB/cQ07HP5Ko51h
Al+DwpHiU5QpYQAMoTos9CjImFp7Hys5c83Y/7l8mSxCLbaYyWK/WgViOt/mDusG
per41PzcTQ1RWRGerJaMSVltyQ4zVJ4QQYQvtez/Jt8J2eEMFSiw2gsFdHqPokXP
AAxy0LDzxvN9RwcExJLFar/wUOXKSELkgfgF/rKt2g5imYJX9XwHIkZEs1HnUjD0
rB3vm/6YydyIekFcoOIxuFqt3R2S1fbcC0nm2A3R1948fJrYdorGPirLDB89PAqi
tWrOOM2z4tDq0eitDXfMUIXsCuQ+q/VA5k3M57OScRoID9+qkpIaai62gyMABn9Z
UkGpm2A68cFd02KYeTYGSr+MAveWkDJgOenRuZWApdhg6xMPKoLiHCOy0+B/KQpX
MuTlhcKhGUt21diDrxmm6O2+ZIaF28lVmsNFOhwmHfsBkTLpVm9heOLmPxb4hYtA
0pPe1Dvh/8/Jm2QEgmVG/LWnwoHWVEFThJ6e3lU2cIOcZNHN2EtjeUaRe5oCEL+S
6Ss575RAXInkM5AZf5woD21pd6MYh3fTI944waFfEzMriiFJJraFnhrccMWbghiP
Sw7LGSF6Tt3zEjOBFAwRpbmPO0NZUtovYVQ/id7GcPfFxxkoEaRWIwPlu/OWZnYM
y0ObpWUhDUlAVv2sV2B2fxr40bSQ3pxXayWkt6nqAi8abHyyAkwiXGc2Aw6krEV8
3YWyI/ZQfw1sG5TJQ+wv06h1PFQJm2bx+xYFcjwZPOmTUlpw+1a5xLaFpqlgpZp7
SR+6B+na4wK3g6/ruiV/mExLNNPvLkNN6jiBGHEOQfZrEnBBLyhgdpxMmg/8GXtw
4bOO1EvTxodMWfYKWf57sXWDBEY/npb1gH06+HHE25Lh+H0FgcGYNoUFSqGxBJyO
C7E3D2aBunuuT0QrVHJ5AyqnHagNgkqY7WWduKcahBMw1Gu+9I1Ui/t7L5gNatkj
CQtmlh1v1Ui2Fy0GDc8dqtdAZtGjqr1iLRKi0b2ZaLGl549IK88ojr9oCKXmAlP5
Ov9P55I17hE9npvvRaMpYWJxEwzRJbYh24XcdFzik6GVhXDBY3c3tcZ/PAZz03zY
6fEyT6N77U4rwXZbfFXd6KI8V/AKe5vuFy2+G3uFPI7XZJKSXVnqWFr6rmMboF7o
k/MJhzNXUhjO/M/dsp4Rx5Cn6BTHnEOF2S26DUr1QAHLfwlrSBcf/h3hdP/VVJ/j
X/N+f3ghZxsqx6eNBEPNkMDHc2cK0gAvUl0N+J2ic9ZplFROqw99jcUTBRbbetOb
WsfxW1VRR0wBEU1NrSSCROX7BV/XrCrnIQCwJkoXXGi4rxk5Y+C7GYad1nfn8ca8
bh50fwl4nKp0qrrWrVze8UGuos7DbtHt7vmtTe4SQ34JRGnHWljbTaAT7uRhR1Ej
7Bf61M8IW+wgXbJcGWATXtaM8x0zjkRCSY3P+utgPwMLKrPTOg+zzpZIp1uym616
mwOnMEDlBUz+nNbFtGhH/oIrRLJYXZA9kvGxPoueNjlkBonfVg+iE0CtMfX1wdVR
Hniae+FVATOTYqmJ033QVtqQa1KXCe2eagM3aR2pzRbvHkaXc4J1+N6fV+3f68UE
a3fAbY+AQIBeFfOR4FB+rPvFhF1OhroXRlla+vhWJrz5JW9ieEVykkxwtzLkEqc+
AFwhHsaBBNncHcfvlA2GohwkHIEa27evfWlsd3f4Lqfy4eyVzMzzU++NaFomKKYf
wWPbG7fBrToLgPeubOpJR4ucM9ZV5acoYCTrd9MTMf77SWIO7fKWep3Wgb222o8I
fTtZG8KKekTlx3g5KcHSUG539g6Cry3f8dNimKYrgPBxORrkzR95ZVi8ZLW1SHq7
7r3DO7dnGqRghTI1oCTVQLxNQ9CsowWgdIr1g0V49JPArxWbOAoTrs3B8dqZWrYR
fT/zpTlehsR4olx6z36Zw8bL4ti6+TfnKlB4xPxEDfBSQHOAbs9gnN/AqZs3dTO0
4O1msuGt9b9zk3xC6UEy/QnCmvP7fAoErjrzDqpmYWmW2TkzAoIFzJP2kGMIPExX
K7BiQOv1gjfp2I6Mn+MbMfVSwKc9LvCpebBXSTOwFtXiMLuJ0ca0loFtxqwNVsgt
lRSEy2Bs2SSYZHjvpUQvTBXaOWGyNeuQmQxf0oCKk4IiExtQDTEoMFrM6K/owGYH
4+PDKaFcm1FT6haHPCYiikO6TA9nXJrCPOOLwD3d/u2JEEfz3URaofig9Tc3hHmH
BuT0EnJZc9ZvcXjNYL1R/WtbX04LKJOuObLnaNq24jl6vl7LwwqdXMRS4d8TIHAe
jNMMP03PlRvfnCP1kb+ROURMiCRtjFvZPccA6Q32qjDPbsABSGyMM7quRRqlvY6P
Acn22RBi2UXPzqDO7OLX6tfTAP+ZH5opSQQ/hQJBVH6aCuWd3oNZw+khWk3G9FqO
lc9g4y5FneRVFeQfxSh7btWQxPUua4PqmBVZpJeQZ1fKY/2wUQ+CiFKEnbcULo0N
2wquwuEAglVTi296kt786WtO2KyCnOHHEEk3gWa+L6h01ja/4l6l58AG5zjOLxBu
0/9zJlNoyy3oWDyZ50IanAV6p8EtpUiJI+tU9vpFCciGCV24oNFzkV2fLBIBBIHs
cUCaP7DaYdEeePM8tLER10GziShUwyK7s3IqfDp4HhHzFBtqr/4EEc2Tx7wj6fcF
ZDJocMQix+2mllw7HaepF1eZzZV6mqwtVgxUCYMiZ9uepKuKS/Kxo346Qjlvuuic
+fNUodqcUC09DTF55cSEWBmCVKbd4bi8V+eOgC3omvL6KjalJmQ+LFBfhzMsqTXX
6a6KreSHEKyiv8bpqvJzZXAbnpHtlm1LB0rsioC/N7Ww+T5pRM8n6vgf0jE//HTs
C6GBcAfzIi6h1ZTJcMU6IKMzo0OE0j874NeuctIkRn7+/RlnvSdkZoJX/XaQx4IB
BJJTkBoGUk6cmKDimSj1QdKoY0u5htZ/LKfwfd6IbARhnNVrZi+cfsK+d8tyOZuU
Ea1TeU3LDJ12QvkYgouM59ZSUJq6NL8/lqGbMzXITgnabUOyGMJ2n46SWblJY+xx
Yp8k/Bhkd3N2EPlIpDfh+AB4AKUvEmBFr4QKWaKz5zeKR6vdEsEgTzAfhugTWcj8
S2S7P/B3i+K1zqsp0bbXmMaZh064WSxHawQIlfmMACbPeG9ISpgQ4cYREvY+zpDk
6dT63iJDcaocA1QWULVpA4NG7e7IaI19uX0aMTlCOuWt8XuuvixFo5Bc9zPABort
8z9Um3ve2TGEVXkBcSiYhBYhh7ypKm0oypYUjFkldWwiQDSppFg9Y8Zhr10ILIz0
uUoBFYXvedlzmcP9Tv/J7tPDhsMCgGDZvsBIYfCjsCufkl9UBy2gdyjb0YX6W5qo
ZAV08J7aVMJG7cc4GJaQe5v+rK/8msSukVggJqHIXFmXMu6fVinSij6kMPPu9K0r
nY3WfOFS4u58igLKdY1W9+WmT2mI4nN8uOyEdgeN80Of8NfzmDVP0U+oMUS0gr3W
IfXtiXudg9DpFyI5F3uTMckbgczJUTVN1hsnRO3ReER3QIriluZbHBZko5q4D8mr
ZfpnzINdDFfVQJU5IEcDF3rLpYhpRrY/p8ZQCxZIXE+BFT8KrXUhHTbskjOkTFfQ
ZFsbGEmjJ4dzXn5H+TpQoIqB9NcTpBaqeBe+kdbPOYW9mk8KlnusVXceCqBYkHd1
dQ5fGieuxKFwSPyT46H46nUaiLWxq+I1H94aLw7pG2rKm6A9zJrlfVccYhTv5UES
uL8YMSNBGQO2MOP0qRSicpE8jwWB3K0Sxd8a2mN3B/WFzIUJVB8KbG/80sj40Rg/
w15rEzWnlFUlGu/Q+Yz+FrsqHthZC8AVp1aGwUzk/x8v2+ULNQlnqaQezOcsMHsG
O6M374cxTa0X9LtFeREDBkcKCx5xXWQMfbMxquMWccKgX4ybTJu6csb1m0XAUfEX
pIDs5zvPR4Z6xDq+auh3sHHNCTHqLwZESdofr6WrHs1etxllU7ICT6TTm/6wUcu7
fwxGVcpcOhWLpwQF3Vqal5wrJPEd3ZUdGZ2YCRK7ZgqSXsD3IgDlQSGiT38X71Ra
qJI5CrGr3tftYyxzJJ+3TaoElF6YZU6+0Bqn3KfLHneqSOWr1CvvNMDFr3CeD01o
udp2x5E+eNBNFVkLKBHH0X8cdzC4pwyp7cMy450Zzg43l+rQwtGChSfQ3cMCzVDb
F/8iG0sdjAqb4rFh5hLr0QJw4Q+x2mZd4AkHiCOE1jWnPftnsGI/kaF4jn+FlUJT
ihjkJ2542k5EWJEdY0WEoFXUxd3LxT/TOjC0D56MyJrNif46evnLJuZ8zLamEyhv
sH9kU8nLSCc9dG6ycE3GrkFRhzYpqAfqYs0im0U9G4Y+vCnnxyKViDWzR9kpvI0h
Qoxfwf/ctj4/ZNkY2W2O11MNzUG+3CwlB9qn+3BOc/ZDXS22fObnsF+9Lqpr9fRv
JI48XW1nv32tEriVeFr1r+D16eB/yiyPfXhnC1L16rw3yAVxvArFddsGwTlzatGR
hP3Yb6AOG0JBrg29EHgOWzeEBX9j1X34ps/bayvuJ/rtPN2+n0mUBNtSX3TKiBvy
6Li3Zlh24nzG8ovtZmIXKKqk0K1gYvaqu6+QqNVKcwIeLdFBz0A0bZeqg44Y2rbc
NxfNVlkriFSM1KiCbO7tPcMrAKoyDnb/Vb0rV5olRpNJb/AFP+6T51udLUbneXMQ
7Oj4XFUhl0PPOsMFNSL96EqnZ6THhNLCiJCCvdQvTvcoUTo82SJ5fE9g1jiFXKdS
Mp2DZifTdC1dIwGenTmz4pQr7K4KTQHb6LlWWt6ngqHrT6pg6dW8agD0tFqoVHbk
jncU+zF+p+BOVHtSmSG1d4ytqBjej9JGR7pHduBgVk7d8P8BQCB8Xa3sh322jM50
W47nQEKd3cduLoTj/4F0CSSH40vX4vZDTfe6FU1NraOgDYpVHFzUYBIo9LYElEBy
YMCtr/TJMIvS8N1+wEAD1qbqru76RIsdVm+Gfq5zmwMbatOsAdLnRHgZJ0k4w0b4
BoyGMeFx752RDi8kLkSLBjM/UHFjxfggvNvrFFw7xXkeKipqtpa72FtJGbyTLu5l
tZ546nPNOTy+hX/RWSPa08vcRsm4csf0ERPlZrxyhSFQPdvVuyDG9xDAwm/HEZqV
gvQhR70o+PTUK/nLaLljEVTIy1iCwXYhX2A/gUl5qBTpeepzjodneJBGKv/wOl2c
cNSUIsE3Flb7jJgxt6DYugHEjR47roUVb4w+SvRs598QSsqhdNCkI4m7jH/mcUJw
P1p4RZw65q2KYfVleS4NaPCkJ7TZ2F4G4HUcfmd3VEJVY3eDEYKMEKkXUydzc0d8
XL8cXZmP/O213tpczIEaeM+RJflUV8ZO2wrZ6ONX8v2o6Mz7DyJsvLkZtp7yTWP3
wgSoVqE39HLJsG0qmDpHdQgSkfUVnN3tjRs8+OignF9FaLItM/vCdcocTdc/gvaa
JrcWaX4FnijAYhKO+oKSaEvO3tCmcPJlXoUq8rhJIhaq/N2syeL2Xjz3a+K5K2+S
kDx09+KOsT3CjJ1P8BWoKxHReX4SBWN9MiF47yNc+8kSs+ItQlYG3X9aITDRWSDE
nanRPhAUXRPYdrGPvpyxo+eOdwLSgx2qsTvyoGS2MHMsk8pSgjbtxKtoQY2S75oY
Vm6010cVcbueO6vv4qRS2bObOWsZBqH6g6nNRa+oaBdjNox7T21NcLb6xgVeEKiX
a8M6b5CBdAzLYQxeOhqrCc9PeEYIBXVIVCay4GDdrn6DWxpmXX+MgenscRYAvxVM
+pOCL1PzVtbPpYlrtuDO7oXFhUDeNismYUCZo7iS3xxv7B8u4KGb+/SYqlBNJbO5
WC+jsHoYA7aNj8HAsPkj71fobpy32yBAF+VUUUK7aathJXvayipdTPb2O3xtut80
XqCdgO8R2mB8vUv/mTTKjydOpYbf1j7XzmX632d2mYp2T/Ub7ExtGsV4dPYubxTe
6uzXdmCGrWAO3R/mz1Uf2jn43g5DTWl1t3m77XbvJ2FAEbJ5xX/wr075wfRKlVgf
CCpUnaosf6hLbDSZp+B+PDmqSzZ3uHHdExL+87Zdn5vK110UTIt2nJdd3JNprsl4
i9DRMDcKHRgELqzeg27uCnVaCNPc/KbJcQh5yCQKCbErGBwQQq30Y7A6USqDzoN1
SwF29Tpy0kMMqBKqaSGYRqzxApkePHxgsCX+DqcldRHtsU4//QIJraVjhmOdAYPW
bE7/kxU2LiBbHcuVAJLUKpxiltnxH8K/WmUKACnmKXLoilbekvbodYNYSZN59R2u
OAIgHa7LsP2oYg5Wbj+t00Lqh4DR4XFc8IdpfS3JBTuIbN1rJV1zDzOXyTKNNIpd
dErtbZTyZ/DHE7Z9aHhovwxiXlxW7jXOetcGaGxejycYTnh/bTG5ppVFk/FHAz5c
6VIargWW+bpg7807W/G+hxVhcS8kKrbjxvL8xZr6tqPLiYCVgSFfTE0v6HLcIbKm
sE5tzU29kabJqFCxM9ESm+xQBM6XhE09jDurTnAbPlz0dbV/XqQxLegv4OdEaQ6O
FpDK/DuEZ4+12b9dLrtCB06GEtRjl0hUE48lF+OEjd5o/vq9czfbSxpOnwHbffY1
JUTj1fuG+4R3cnE2uklhnhrsmHA2EuXpn4UofnGh+zZJ30EQWSIwq7QuESeZkdgP
FsTYW5NZqbJ/70TPU8CJ1d3H6NLYaERZSwTPtHggUjRNDyMrtMdGhTLL3B8Rr20k
KLi3zoywSoK+WU/24tQ2fq1qcYDlx8ISExzjzSnsVTQRw/IdTq6RGCHEZhbxQi0J
OO+Mbd+NR/RcDQbmmFxOHHUfVWNH69Bd/v9vON/anxEaYeIiRr7wzBQiwI0uggfR
ueLpVRb/7csfO7lZUnD1sxH140tM1nVcdSiavUe9vJfU/HTV7lkKnRvOeOBUANR3
kgLAVHUBKe5UVNEHli6SdGzww/aCBpy8nArFud9cN6wOPj2ee0d6RkN8STQQET+4
7jD5M8gJboTOYX2z+/JDUisw4bSHLcvDstzm5Fn4pYZuztjlsz9s+1x+I1bYLVYG
nIg984hDok3eLyMla4FmGKGRBDIc/DLWZOSLpm0Ww3SV2qHom87gRDsNc5JfhijG
+E5Cl2RDFZKMyZbY/rvvfrsGQH5w0WrCMMgM+MvvoctHRW4bgqcQAxMr2MENCVCR
zatqAX1APtF38INyLWpHQ6xH7TEZqnzusdAtadmhVoZNV97vxpDa+/R+AAo9Qxpa
ISCgU3VfT/+rfxNe2xp8HT+pWK95Z5+et63ofWBufgfttr31q3oqk7fzzi0B8953
8SikRNxgKwdO7LhGMZjIAp52kO9uFSbJ2zZh6c5sXk4Dv8Ymr9477SUh/+cvCGCK
6AmOQe+0UVm/OpgiacqTvgw6lON3ts/A2pFvXnEEt5rqJSC1tt0UVV3lm/3ybgLU
1Q6zuuoUPvs8879S3L1/Ak5ZyUHFoW6GZIP1ebX3m4sdeCgfhndP17JaDX9xxkEZ
I74TRgaWfdzxoHxn2Fyj6sVMVEGDJ3QRK7waAttHGuKqo4i8NkS08Bvn7qUXjjij
0jsDpqa8O4qKCOUfGJdbfH1Jc06Jxy7AyL/ptNBSsWepEGgCKTG0Z/YCDm/gj1S2
mA3ESb+W0Yy9i6ex2sCXGLm1MTUAt80yr3dW6FAWUnQqGLVkhCtadWIE0VdjpWPa
ZidUXkaFG8PNadEa19eEhKu8WnWuhe/uVbFroVRGiNmOgYou7sHLVUP0j8aw/JBZ
3vFttilBvC8KFdZbpbPBk+Sd1QSivsMXzyyOPDd/d6NS9sSqDugbmFe3De35NOGi
WGSmHLXkQKXrfS3I9fpk2dfbEdfmKSUzmCbO3L1McNEiRMvTykaRStDoTTpfHX9k
bNlyJi3Qs5Gr5tpNPycW9FL+g632Sju2GWBv7wAwPB7UdmNm7pTOL8OfCuJjTuI8
MQzyuBaKCjOnqraKaGbdpPfGXUL7fy9z74B4uzex+cG5IHVYo39qVCMaPK+rR3O0
88mDlMGQRCL6D4jiUWsCWrsobtNJNfmyKuHdKl7b97DYHhpDDh2GSjmly79VK2wg
BuZ4B8y7KLViI21z4wbqq9D05nubdS6cripQ95k1aXKMpsTikZlB5PF99ht43yiF
zVVqGlwqwbJgO0TXTnTudlRHVhkdSwb5WYmq2TT395+Ir5VfP/+C5azkAGXbVlxp
iIPTHXpWLtvuS27yNA+JBBgiV7c7ukEiF+YpeyzibvmvRD+VbT6EvLyFJWppAlLJ
E67X6TbK/wZa4x3sdFf8UQZXqITyzfpdyMIjjNHuYVdaJRlW9NnZwBeIwSrb4n12
PPks/B4ZFIVSFdBsaJogecHuYvs3qjCVP6NnJAEQth2Tj1y0mSuX/B8bXnxuCKc0
kscUuWzLRyd4m2GjQ2DSr+v/V2ngZo4HWHEJWRmuQa+CN3SNZT9o7U13e81axAdW
ZE5LewO3rsTT08jsQjs+svxvIcTCKHWcP7MxWKb7ob0/ueb5RTeFTPrBV5r6DAyU
BR/37DWRSYAyiSZc85yhMMvlEO+/7+e/wQqJOC4ca29aKcm/HwtNl483DL8jhDkK
R16Ej1b1wUg5muALRskZBfr2xZdTJjI3L1w7Pw+QJA4NPemXAwN0FxNeLSU73exO
xUwwdYwmUL7FGnqr8e2IQ6JWHMblp4ea3V/NAhzeZho4xBoV1pPJqT4RC9wVWfxy
m5kg7LdBASOhrCMNgOxdm09CGbhKM5dFMmzW0vxNmHRLwGNpE1wg3P+7+FW8KdI8
RBPQB2LZZpCdgUJr19y27p5Mfyc/cguyOvDcJ1ZJxxiufolcBCErnR/n7o6a1/XW
bvnEdaR0KLoazv0lCfTbtIA3oyuRmi7p92v3X4Cvnu88yLgMR9wtDznFLbTebOb4
ZEsxSqDtGNkvHbsE4yPlpy4i9U6MajlKi2luYRGTkPwMzbtocOxDMDDVBIo5W2KV
vnKhKkZG9z0V0MdBQcHYBQsMhI2YPPVqa5icefi+eNKoQ7jC2MBW8kC8sDwB729P
pM7qv5+jB7ePoiPvs+3ZbIjywdvIMcz5gr/Kn/3yJRmQVkWY1B4tyFny8PhUwcT3
Y5lM2r6iBDcXLSDHHv8MwWkTyWu2bjBtNmIrmYPXJuAjirSjVRkqSURhxWsJEWpY
CEkzEynr7t15OnYKT+cYkwhN/Y2Pl6aCrRuqh3bCpy57nsBFpUrSzAnCKXwbRRpD
AM61vjRVnDfWKi0pr2OQ9qyglklLmKl+nQgoW7rX3Ol3A/tHeVYcfw6tprrhczKa
Vw5FISNThInow+V/FTuNfAoG8lX84gUq4AYVXKeUUFjAaZb9WIhX4rrB5ImenhBa
cyCoM4eMMiPcnO9LZqHmJNyPT93kVc4K21gCmseNHLV07mb33w8ihJy5C6WxSmPU
14I0CkcYLaTSet9dKfglb40FicQt8Gle/BlAX5HEP/a8QJkGYZKeIhYhLwaIevKp
VvXxbI7tK9KP/9Jd5oeoCFoiSOSmAw36znN3F+MHrULA5k1Yb7aUzOlIQ4Hk8UBX
duHFvIs/JMHlpr7J6TD+S4EBPHLJVW+PndTkX5f7XTMtQZ26AUeDQ9y1d0PhMB8k
Gxs9ONGHsR1VU+c0LslkBVpFxow+tWCgaxbCFdwDdzSOFP0UeHjV6CJNfO6nI9xi
Er7p99+igpKA2N/8p2qa7fZ+zQmkRPEGv/gsZ/BU//Gj5lZ9Xxt43LqraZeE2BFe
pqQMH3sL6JAxseVuar35EZFVsRyQ0aaCpya03RuolT+DWbEkF8wuV7Hca49sMz0S
xOKgOK9taVhRT+d2upp/Dm68l4jJJr4iyHdkCOEwzhSRQJQEjOaJxEWxbJWdgYxx
SN+7TvctamkKiQXgeFapGBIYkvCWh0h9zTEtDJvgZw5DYbrGjHnbTthDMTbbO7wW
a/zoDvE50sAeM3JZ6BBfb8525XeQTeIcvm8VVpFNzuWmqR4H5MfDECxHuM+PJlzY
QOheG4v5nKefHSn1Qp6INQNSVaOBNSa3CP5/EvBarVOpfHyBMmqXzDmcwv+aHTfE
+xTVC+FA7qqeGDhHEoG4wvekpW7kK8qSWzVRLKONGYRw6kh/bU96NDSxAmqBL6m1
nia+pmmHVwQSLi6ZpFupUOUUu4PKBrpbJUsKH3Ha03zhiu2FDheF9tzaQnu2f7A4
FKTFLaD7SRP8Enio08+3rNV8aKuEjv7kRoqHIlZkht9kcTcXuTcQ5U7UlgV92QAJ
nKkJ4Aa9oxRCUvfshytyShSXoYoEHAZiaAdgm5LipsdDg0/3LRy6GRLYDggXHEbx
y8x+aTY55/1v4Ap25wyU7Ti9LiMTcacDIpXF3W7WoiuAClYX+1Tjjo3HG/3zuNR4
5j1MhuClv3aVIBQRg+HGUpYlGFwOsEJ40KogJM2c1TCR80nj47sTPCbDwYFPJeB4
btO+eUWS0ZCkfrWpakE/on5eAyKUYEsro4AGB2uRJdCAtSwcImkjSbOXcLK2EQeD
eSSssuLGECXO+q67LUVKF5hp1JoFfoSNebEOsQszRCECly7QIDQzGoMwVvxWS8Aa
JzowaoJBBkY3Z3pF2oLZnWfexKY8OCN+4Zfs01LNEmT80TMS0meUMM9hrezzEJMc
olgSy2eky6QTcPsugRGOzT/FQgo2cr93ZOGJoXgxgcoNETDNSuQ5UTY6p2xtDWG5
GZj14IrhrGa54EpkVWIvUZy5ILkfdrqeGOPOcg7lKejoQFfJiJfY4Mecg+0b2B4/
ZskPcZD5ZNtWwEekZZw9QO1b3AzLqM6dS2ynuRM2dB9QPF2yTjtq8q74Pqf4FbCo
doa9kNFTRgxg2ZPFSKNOgvaQM7pbRniew3BMO23dPVdwpSoVFu7LTbtSuYvTPcOV
vJj7CR6vmp+PMXDhuv6wm/T1bTreVJ38y7xONTa5XphjSOJ7YTpYaz9RpWtADo+B
sjK6UURneK7QdiZENFeJU77fucl9+YO9M5V0DYqKaarFkNLM2TwmVChr8LVtKQbm
IpRFKQh8dokZxyfyRUene6AXoBG/3zvDbykUlmfSaz8ObCq9AIrnjZeVcu8q/jvI
iQXx0w/kAJnmGYwQfaWV6tArHKAaJH/3UuwfEt4wjnYxl3NROzL6Fy8tYeM042yU
vO+8a43L9ROMLqPsiGHtfxuC4+nAFdWFEAoS8h3KwOi/xCPYSGXuMk1/QvHraq12
yD6woTk3WuemXwIbGHR9Lti+SIAFbzK0EGoaQcgAsoGAk+y4cueJil5lgYRjZrbj
NKNH2ip6triIsX+6VnlfsGU5t89pA+ipCtwAGiYkqX29Nphw7lcd5oTan3EoVoeu
3/Ea1TrApUqbj1JI8su5uRxfaNXPeCZr1ANHiiu+65YkzEPJ/rwOtHxLhYck/IcM
yIyc2qcRbUAimyF8yW77YTmWQJjnTgnQXsWZsr9tSBaD6JaOkBVkcfxU0kXDUNwL
+BPd+YW6DVRqfjI60mp6ilfzoiez6Z0Empm5N8pZXR8aT4tV7AnIA0zbc/Dbw9Im
+cwJirB25Os+BnfjbBPwfsyAr7y0WYmhsxBW1bMijl3W21hysgACdW638nJNErOO
BSQp8d8+Cpu086ahL/28gUsZQK+67C3va2K6ng7bA9WO0Lp81rG/avVzPCukNFDW
tudY0WDmJj9sMrVMRKKrYrTl3wi2fXVOq6TTyMuFmLQUH6r11JkPcNpxU9/jc3LN
DS/OdktC0/I2xaMjghFkIlYmywUySwBT5w8dGWuZGYqLHkG8ZjnCrz7uON/WuHWt
ILz7DhaHsw3gczobQWZwlhwTf2h++qmtkhgyV126rS6N130SfnrnaRUBcUJGnAga
iuQ0glhtAFwDVSy24Ir1Il7ceLehf+IgkJDraUVqsrEO0wRs0KMevPrB/5Arjwgn
P8fJonvWTWHG9vaVZ3i54Ie3oigsGmM75tgtrQCMKLRpdlxQyHs1oAIUY80g3gSe
97ug3qiyEZG5QxtUrHezuHVN6OebnJZwxR8FsVr75VCb80/eqNIBHv0XybAa1AGi
wXm2/6L8NK2/eJ0W8WqCub4QSMnNRar8YalSPGeNFy5LYUoYfY06p5mCdmu23wmf
mxYZGfWcIC3RvulEqYnfPHjg69DbpYvlSbdJwhVAszJxYXeB0U5GDBrOszQRnpFb
8OhHSSA0UTrrYmedWKoPWpwQNN9N7mbjXO1PqOEH8CK8FvEGtXnceTM67fGUzmFA
LAfNRQZwEtuvpOFn2ZK4TpI6ezwBlE/bdIfcYYsLM6S+MQcA9qKWK/xxxONfi8Nd
APZlnvtynnfcCxuNzRdDZDqZqf32fuP2WfKyhr0/oCm5O6ASKH+PZt1gemaYrmhp
znvA3xbxMG3JlVSeFMShPfvCtbwKjBQK0iIBdoU1w1N3mDulay0ZqJ6AInGe7v2h
xScv8YDXsVjH+30SorBc3oT622lyKUwOzCLe7mGxUJlM5Aes9rrFEaVGkCTYw94+
/+iRSgdJcCHNEeAQpMg6c5Tz0r1jU6slgAUShp5onSFXE0qcYyG77n5rtIKmPVpl
AhGQip8QrJTXuwSMcIyY74CGLIvgcmCXAAAcOzDpXg+a3YOwv4pS81Lye7H53ANV
RUoKZb3fDu2Or+qEDeji4aPXo3OCjFU7Kkv2HtRYqXj8YUV8LK+KHRyPf9G0Dsdh
91ZC+HYzIV4yQ7ywmM8HCsyltk4OnCD7LdSg3ojrvycM+mUnksaRcZHCzjKyCs1V
6Lsm2MlAsEpZxwmwQxYGfrkB/ooQUtZ8hrz33X02Wk5i6mWxOF8UiaQ8s9B/CAxo
au7EjwmWBfDkurUhXkRE7tOUL1d1gNS7AnK1KBViS3qBfbLRTSAY7it0xl84XZyv
Unk3t1BpXTlQSn+ZTEzcj0yKasiJCXnF/kJ9kvxF3KAk8xoQEXl3EUztrCLuDakj
m9aEw3QrAc2Bydi6rWuVLsCIMnjYpl1AXBT8OxOpwWgGjqS1+YuGBFn/oTU1GEw8
d/Rpn/nv9Sv+nuuUkD0HooML0tCKhVojAGvMTDjYrxRJ+epk68VvUjIm7dAc0B6h
/wWdB21DKJREBMuegp+kOdCIUAyUGIsn1hbFh3lKsWJmVNqiIjx4Chj8RXZl40v+
ePMnufrFrFQXyibDjSoAaaXi5mb4zpLe+G6oj25YavL+gH5Z3uoStW35/eMc37ZD
HjEM9r2FdZofrQ/nUG7UuAH8Pt7aPtL3UqrtAixC6IbBvpFL2DGucitlw9M29PCV
G7u2SS+hOVbMbb3L61kJ581puw+bMpNz8zCVwdlOmcxo7XMJJlZ/4inZBI8/oqEp
y55Nnck8e61HioTNC6ME9i8Z26HfS595qKHsM6heaEzqu67RuoCTUCX4HMDrsgU9
oNulWn9B20lGoD8nU1Q2v2dCGtQyaf1ZHwEo840GvlqQEb/p6e6kgQ1bz2NPs04n
H58ZiQL6ugTtSq1VoRc1vhQUDURaPE6y84tJfFUAWY3GkiNoVc9wrU4CyIRYe4nd
zpR1HofJ9NJWaUpQLmm8jJjcoI/lUMJ9/Wd09CkGAL754jxMkUrQIrDpyElQO2Vi
WkmeSz+WCYoKNUB1RFWqnRQstMolCr/cszUUlEksBqAFaVMfJCK8JHXKENdFgq1q
VcnXHh6ABlxXpma8SMdY65OwByuac7LCM/uVxBP9yWfXJibMIxToc6kDHYscT8/+
U/DCi5DZJKtzkzAWyjM/Xe6oB7pvs2uK7413I4DHHJgNgmL+S7+xcS5NO9v9dc3V
8I5m8dZJ8ccZpU/UUH5fNgW1gBULqHq0T2gn3TD5GvN/B+SlIcTP9acz0okeLuHx
WaIyQiHP8lnZ8qCt/PGXsOEUCZ0lu2VwS5uJk6eHm/owFtlLIBdu4w5K40VqzUGy
Wl2yfAI16QkEahRq5btQDknB3YBFd5B/7Ti2oyN7HRIW+OS1RxQZwCO9swTDi6Fp
sV7ovvih4P6KWcmGb/S38uTPOSBga4OPlfb5/EsTqtivcsexSJvA/wXuiEaErnZo
8NZp2MZTLjMDuAzvPnvR09kRE3s7tA5tlrO2iSNDkqA0o/xUP0R+jPDfRiEM5kvB
CfFGJwc2VTEEX2tbCdO42gB6zpOJO5WQnoSQ575lyxntcp4lFLulfm2UXae9HuPr
L6tKwPl9Wbm6lm1ws/6n7qWmPzd2DUxxpxDBMZErlj8412f0OJsGMg3UlRjgyihx
AXQz4K0JkQWC3oK1L0MyctHEeggm8R11uy6hcjOMaBE59FzV0CeAqQSBJySuWAhl
5pwo2MlsaAeV7ttJ+teQ381MyBpoBCzRbT91blHOWXjcCWrUHbJwbDu7GQ2YuA3p
dHGeLGuV498Mz9prxTOTKiqG57g2yeMcZOMloEOzvN8rhGZZuOm01SiNSSrbsjgI
CwD00vi8xqjeXw87kLoraPv50t2V2A0Dtd57lLuNdIzsDjCzIdUiDm2iUVKa4gL1
fjvSJxipoGu2xAgunY+iXGZL2z5XPVFYfatlR1Vx9abqgwYiFsoQ4hTtng/zAv8B
u3Uh5CRl2xpYO7B4oJmeYGr9WabWV2r1tUSaSbis/WKGfNIlwyH9clJppufA7Ish
6Of1takHjzBRAy/crFpIMG+enPLfsV+K98szXxY/+tG/0ZgMFdGnfrGV5bRBsBHa
hmlO99GMZyYuVs4kIE2FsulF2M80gf49HMSC9NgUOGmoGmGk3CzcLcomLsfhu4zj
g+P44D00m83an1WOPFclWcjjphFZXjEuY+L83T+7hQvas0pdH8b8N1mzq9P026ur
gHdo/nqkhs/t2V3CCNxkeJO4cuFjMCEE6fV7tLyY07odmKKCj9NOh/Gu57yohUVH
BinpM+xAF/XSUmDFLLGdeWGk/6061LSm9+3lVe7h6+rlyLENM/ha4DXv6beGH2R9
ufGgMHXmXS0buAsAGS1kKGYyWBHn9mkKc4Y7Z5Zkmj4m+2ksTfK67yZfUmKoxjCu
phSY5OHavosakNmCcaRfeHmYf0a+xDDO8ILYPtQDWpZUGHwmnzDjV3sl617QCuF3
mHwCv+2uT2you+tCykTrfSO0GqIcC9T9T+fqVjBbHLucqseMFHbz5njycPlGeV1p
0N0D3gQnY4YPd79w2uyLqIS3a1ziWmJbj8E0Leqr6NHJzsf/kpfaKJFEm0Of4EIk
HBJLp8vcCB6a+aY0yIAAuiHMle9+OnGX1fH+O1x02Av0AYtyn0KmKEO2uSVMphQH
abEcCHGc3R4AlqfjFNa6SgdigFVGqkvQz1M3OgfYl5X2Xs3uzptavr30LKptlEbq
mx7xAldNHQv8hYIPh18gcB6VK8l6MfGPSVWfErTI6zWYQr95hF4+d+lKh5rWmnA6
IU6ZqOHY5eeEkzonul7LejcK+sZB8a7CEYSSCnDirhRpe5smqYxXF23cSlaVvBtP
qJ1hz7/xzmaipLLvnjA5dw5ZQowvLqzOotm6vpbisS5BFoD47o6F5HOWgPUSEt3l
UjD2OKfmQqL4mKSomUhb7UPhXxPA2rNJu8hevsLMMyw2UUL2hDxrb7DvAZySybO7
WUDhacNpPgOwGBxoZ/3nJYn8i+XLvk8anG4q1q9G9kP33bpqHUkRwZWeub9OIE10
x9gYBEj/F79tRjDpFhyvbpKLhC0EKZKtklrHr2cbDB/OrJjQTf+w3Mrz3YncOyvc
3IWioIOVwnY7j+98ByT6EciPmgpsTcCKcUT1ag7GC1EVP9mfpRWs9kuWnoTqGrwS
qUWZt61T6jZwjtEGumn3jlGKsgqi6V0E0svRFXUFH3ZHKYCWmclgbRtL9ISkwE9g
dnGx4mexIukba422ZxhcWvNQs7fC92Eu+UjukoDivK+Ubi+c4aIRWnzmj+X/PFrU
sMtZIndOf2NSJ0yK+MWdvkSBXC3BmUf6JdZrDxNoZ21WTRX6EB7K9W35JKac1Q95
eUUcIMRS1GmUY0y6mioEhgT2kGJawdfPA/KIt0RfLzxmlMg4uFSTjjUu/ZpR5OqG
qKQNcKhqYZEZUHEz8ZNkshmaE61LCxIsGjkQli5vRfg3NpqNhTPgyOQ+EtUsfE9c
TOkp8AcSlZZslwE0tVy+HjCZKXqsMfHx4RtGRokYoMXK+DG3Kdp+843TkchfG/Iy
Wyn4IC4mB4ZeWxPJNxtzQbd4g+iIioNsOsY/MULO1i9gPhCNp3OxFBJY2qi5qz0N
7O6EekwOQwd0iL8Sk7qDyzD205yV2Auf/YIAdmjZlkm4ArpxVXGmVdY8/6AbKweA
Yh4pTSVGB3/XVjyNFz/4STmmGY11yBCpKcJdGa2p9vzktnRgpIEFN6LA+zgDNYV0
m5sPWeAOqhotnqiK4n45QkJwdAVNjVDsIgLyTpQiHO261vVuh3yyYKofXFyEFSwR
YEK3vzzrGcaYDDJP8eVrV9z0oAsuD8hIHur+VYXbk+x5E4taOi5VHlkQd8dUMuV8
zUijCHVwNpbMisyFUHUPWUnj+sWBrhMaB9sSssDuk47w14Ka+pg8YzzQtiNIG60R
UmQ6vEDQDsVhG6LFgLt6mucC8Ipk+DfMVKp5wWqgwtUITGKKMXXF1/K8u9FBpTQr
ioKoWCSKV3y4zDFdM5XN+UaGM3L1imFU6FAdhbbZyxclk19vNYU9B3Lx8sDxZ5zF
udOg/akvcSYrPYkjPMmGpIYLYkhJE+ScneE3STjApXSC36nRtA4E8HaZG3LcSmAx
5erlXYFZH+hxTds0KvAE5DNVH8ztBwGGM7vRlLWd85+9yrmWCAxiaV8zs02ZKpPI
a6F7Dik5nv0kFn0cFJNsHpBKpNInjb0WkeN3mVDh2HdCi+EQuUc4YOtq9CcRfUbW
7OAYimpc3xDDiCzm4oE7jGyU031N3AeBOwVmorRkrG5SkBRcRpr1eRqHdX2cAHup
YquJklVbIUOIogzseRIzwughLU7D/BNq1WkiquociPssZTeksoUpVAwStN5gdkFU
Tetk1URyGX9MvGi6G45/JXzS2nen7jhEl6+DnAlTgwBBZ4MVrfVmGu6OSe8pH2OO
1Arnf7Dw9lNCk+ZqHTe7j1YJBS1BQxKkq8rfTAWJrm/0Acg0hSqV00DKsIrE7e6t
ghQbzi1NNSDkvdvbcVYyTjsznSUUT5hLR/9m6GNzpBKt/CZb6UA+ma5g3bHUAvDx
Lxy/dwnInyulq8SB3sXk5SGezkbabofZyZ868KTNkIfwKIpc+ESBErBVBCNV1Xl6
af90AdgZ/Bv8+He09ZKUFXzi4kDtO7Aiq1kfyWWwbEphxtqO9RI1bDj03jtkie13
xDH5IdVsM+O0qwFhvkF9aoTUwI4HlSLP32pfN1T27QTfgm37GZ+0tP4PhCnmDHCq
r9pZqkX5NYKrUb84TiIs/AveoXO1Lj+7lLkx4e8Q5MZO+eWTYyNBpwlOfNFiu/Y/
uyLWVWtGn1efHT8oU+a4mOEHDRUwOGoRWP1Zw86dmZyCmCBn4ziahWyCGW1v6K3W
CMd3gDxvBL9v1LZ8J7Mzsr6J78B8hqRPrmceDj4KB19pbT/BHzy1nBeDJw2ybcSl
MtxDEFnTR9gyi7ek84DXBVsReNey/duaFhoVIPtDSB/5CnXmVMdctKj3Tc/3eI11
iXqGZaX+C5n+7Dunpo2KkKkE6f5YNo442o9B6q8/Se77JqcFSGhxE+ocVJROW1gt
vi63Lyyvm2h7iL4lOZs/JGf0KzrC+19LKa8PSVi349kMln2GPQMSDJ19KoTsoZvd
hcbXujk+l7Edq3/Bbg7BcB+NnW0xtzwJ0IA0NV8JZYk+Iz0jlaO4+3T/WzP7/Gr0
qosAAEYuD7hd6QHFL5cJGOxmfkPTrIFTMhZwPnB8x7yQvsOWAM1Wdo2LiQfwVN1v
wOY8kXToeUzAsmS+QQ03uGZFua9ra+XOtKHOKNt2xD3mRZI4x6JXG9vyWihXZj8f
TxdYtqxRl1oEhjzeJVh3ANztjEuE0QYbrTEtbZcWdOByGJQGhvsM1kDy7dN0gxJL
9Z6iYSyHrzZc0oIhmUKUPur9keYmvKUNIr3S/HSqp4HTRUjZ/ATh3bkrWMaR4vy5
FahAir9zbTF3vbTmYNHrjXmWEhep8MBmbqmXd4muQnBOGu05kcj80TEsXdTnXN0T
sfzzCqCf1ZSH6XRwPF5Ux88GoYPrjKqVZc7nS85Jw0FdofwTYmtw0FPjP/oc5uKH
YQmrARv1cqqnk8vaO/9C2Dq5LDB2vM8YvAQnittexLuwCztE5tOiUFkcW7JZnfz8
c3QHWseB7AoUNlt8IGE8DifwqGTTsjencY5GYStLNnmwLqi21+1zY5VouzeyLQ9I
lYmSHV9dju/PuV7SU+rde6BOSxDtT6jmfV+8n16mkaM0Wbbdggbp423nTaEsVgAG
dOaiJ3gNg9FYrXxNipSLpmctsSpEATCZT2pwHlMkmhUXLodVCYXDIVEhJrgxZtVO
dwAjHyQxpPyNgjqSwrP2vvz2v1mE78tfNBiIDtPypuAn5TCd55X5BinRpGsdFEBF
R4HdKM+EOSwA1en98f2AnEkkys/pp7chTfJx/yszFKBefVc14+ksBweHRr0VXdLm
5i4EwkiFc6QKy91uTX9bu10oG1Qb73We14nvTH/45DUdG3cQVr3aohqXL6FjBezN
vdISnJqX98qXDGVo/ux3fN3RU7nziQ3KPtZfBUvfPOtm//ynDSOXBrlr/ah7Kmjk
vwZQu8pmWdDZ3e/w2B6eYVgnq5hgsFgVp3ZzPSE7nQKWUKnSLo7MBNE4w4eBxhSW
YBGOMCEs/lxjon8jih1CsCHNvzLMgDVegBqlvLJKpmC68tb/Yie6ThtsxG4j+tES
5DkElLabLM8KkjgF9G/v1erJsUmSd44X23J4VnzsUZaQ7zqtbeJiYS2OdH2envEU
/OfsxP2yDLorU+et1H7ao5tzc6tjhFJtXxm9uPM8UeuPwZwW5YRa79vv0QKkmMEe
ELSmB6g5AcUby+3ZgncHQB2h4+HQa2hZmbdZhE+Iy9OjUOh5X5XMkw9eB4PCUy5i
haRL/id2nuw5+MTfdBHko1RH4L/kqh0q4IBNXn2j2ZNZaylkv3nb4+I7SQ8amirk
KzCgOoEUmyGqQskhevIpOYTmS8q1wntjpVmP764GW/lEkxUxeGbdKozpj6r0nMHp
yw87DHPAXWKVIRUW5PqIbldpnOZ1Cfg0bqz7jUXZ9dUtxw6N+c0V9JIGQfUkGkaa
9uQ455CUjO3bXLQaeNSre6q+PBXPeYjf7x1WC4SkyVrjGtzkB620VLkeS5Zy08UR
YGlGZHMPpfocaAW03ylDhp11C/22enSTsMfXUJTURLx0p1Qc0NJq6xF9EyGg/+JP
hokBhLc817isgGSjzbeYqZv69HCd0vwxAc+SplZhGq0sRBfx8bRO8rhqpN7Ir9SC
uJsuDiaoM/ej3TquDfVNJFe7JhQi8SDvDHNvIuhWtF4RMPZL0jvYZZ9wk5ptA5Qq
XEGEIg5uws4Tg/0r3O5yUoQhw77QorVD8uay0pVxvUIG0cj98eqHMqRU8fFreVe5
Q0ciZ7Ixb0UbuN/I+N0TnjbmcJcEpmhQMnRCekMP9G9wjPeSXGFpe4//xfG9i579
hysns5DIpaVcGK35XJULXthNZ3yds3tF/TSDf4LtUXA8DIuq3uL1lr34sIFi60af
Sk75hqRf4Cr1johpNmqwDHs/aNXPhluwVs4JbDUp6Ycy+MiJtPHiLiRqShD8ulPd
Iy3i/9FYhGHYZEduMTRqLDZmBayhmw4M4epPL1oDV1/O267yl2L0qPNsprUpBV6k
PQNMEYWj0IPdnSurX8HHVotk0fuMa2mm15Em7oLvK4Dox35lsihDr8N7S8hx4dE/
gkjfMKo3eufbHuaMN9Ngasje4G4UqOXFPhRNgv2kFYDeU0s+Fim9mxKwHmRA2OlC
J67G+9a/LVoz068junUBeyK+tt+U9qWiAvCiyYJynL3A2bN6oIDwcZ6Lf2czWYHI
QdZXZ9MCH/OE5xUwe/A217yYkrUcuUzjF6DQnN4Iy+EYlpY8goOcJ+nqwkoiU3mh
MYrYy+4cMNMPJmzs1i91jlJbH/+mG0TzqN9VnmKRYLy+J3LxOG93X0uo5Q7I2oT9
Yp4RXl+VuDH+NNwVt1EINPfl/H7ST0suoxPy0l84pM9BzDHauCK6OpeCEul79hYI
oOTfdRhNPVeWzmd9TGthxPVZm1Kh/3qgAHyHstSrl+36xkluPfCPCPhVjnf5Np0H
i4WYrfOcDVWhS2BICgV1c0lvYOqyym+tA90Cl2wCkk9hzM6A4Nyh/Z5akOHsNirJ
wQnxavDyl9m22Qk4tEju/7UmdV3BHiX6a+H8+Mg8MV/EwUicjyBERRRs0iJzm8j9
DiROwmuN91DRwiZniHPqhH39kai6QuYSxefkOffJDc3CGCs2CuNGsqMJ33QtXzEy
kQRs0e+MNN0cM8x49l7PWLpTqoBqYEw1hulKSRo4x5nr9hk2bUAbFNKjFWjOx0AV
xUBdTQsJEVZsgRFmiXPpgd2OkoB5Dai8UW4dudYlDXp2Slavpum7G/GWn4I6fx5C
E8pilNG8OrTI2CiWQjXKluKExjQ18BAAe4NIgy01c/jwUaHhaN1D9FQPh9oJ645R
CBF9pSokfj6VFtOV/H3RE81JgQ9Pjphhdm4WqasbPaQ6DD89FoouMuYyC13022nL
Ce7ePVMFYCVaQbqu1n7Dc6ByWeVL8n2wEKPPhn6N+Hvymy5d9egG/s+eW5Qfv6zs
+ZBi/ltqmVnuUlHx65ELMSlBEXO47R5DKTA/mNwWm3miE9gl8rEDDiZz43n8JDOS
MgBdZ8rAbKEXJNP2ZAZecwcceSvGwSr2Sh1ZQVyt5NylW1Ab8VdDQdgdzoq809ou
9xvnAf/zQuLrQmLAghcCdwX/QZWD6QZBPMBarm2FFlqvJ4wicXCSkJ478J4vdaon
WbburB0AVinvwryuHYFmKrHFJvf+VGGkm2xwOVq4N7IqzGsACxsWjLT92juX2w9W
r6+zdbZWqfuXQjlinyQ+ABltexGXiuBbKFBvtTcqfo/46nKfwP4uUMjxAat36HCc
lkHdEFlmS2utYC8wQo3AXlm+XsMnQ1a3aQ5aKWqbtmwkF3VIXqkNteJZ19IOya/M
S4fFnVgS+97xrHahkDHCqhVZouwLk4xipeBOKEgWFT8mdWq/SanffPOhJTqZyvuY
15bfHBnh6AuivcXlu5tAybwk2h+Yz57dN1jKh8XxVsmn0biChU22nvXIbaIpVVfJ
DqM/xtS352Jyo8jgyAbRdKhdiQKQsg753b7AXIvLQ5eFJRiKZrJzc9ujwlTsw5Cp
/UTODfHUQnvVBB4NmCkqF3fxbB0X7U82/5GezG4ZqSrsaTLohtDreXk+uRt1tV7z
rWRGL+AXM2SKvD7tF31EK0VABp0RDo5BwkFwgWXtgHNcSpCNC3Y/FMeQszPaIfSy
jmINrFRuxhrYKTkZ5GW/6Z8mzkgGNUQaUZmUcPyelSSqs03saN2QDzN7l/YyRbEi
zi/wVKSFp1RQddmPPC1uOF/D33FK9qKnPI+AFyX0HjbBYnWAKT1tJCCzp0+jodEI
KBaqRILth5UUMeti1NUaqsplZILe8/W092ZtW8ovo6nYwVjID0XEW4Y0rwmet1k+
mnFTMJF0Xm9bFTWEduDvn5NcPyLI4XozXUA5LZ30gc1ajSmapu4hYbKs+LQqcHAf
cOVzHUZgf+KT4exWk4T2UWBkT9kaCjWFDDJo5mbpIjxlbggIroUjfPIY1eOKhRoZ
XUA4+3nVQvJ6R6hunNBksCo2k/LO8+jBgQvOyw7YpXiCVqq7LEpHhWrBP4J+F8vK
C9Da2FjQdftVCuIXNgfisqr0msljXtuf+xdGityZIENSXIySjJ8VOb8vwMJay7+X
JDF6WF0quVkdsi8qzJY4CQUm8dLlz4Vc6B6H/5e7XDmnsQk54QXQa96tDXPxPoSn
7kOIy2J4Br1FCioys6850jS1MUNpaTR/wa0yMfhO8KA0icAN4nPuYabZ1AGeC8bM
ki7SHdrhw8CLt4vxmWixoe/hotRjpFfBcH5JKR0S4jwh3IG+fR4MGeRMf3NAgK9w
yWFOtMltgMdvjZKgKFTxp94Bz6AaAwMxKMIAtXxd9+bYYSP6zllEq3qmckV0piGI
rRL6RKEPlK9RjwGATnqPL9xM+fmc+ll8HO+fM64yTH82BOIhl13eWnfWwB0YUneb
5dHw65DL7Lt7KwwY1uPFyFJOeoWppJ9GYXZ2unTrZmkgKIVSqlsV1XRrE6jp3c9q
Bxb3QDyL3nrB6T564frGG5GjvPLKRTF7E/bnzQPehoF8tRW12M9oFaK+PSwiWOvi
dgXIutc6x4saYM9t2tJFCohJ5aHKNiurs+iUPikT9FjiL/wZ30YlmjumdYlyTwk2
Ihn6KzCqQbS0Z8ATtG25LSthy6mdHfgQrOmWQgt5qAMBtjmip+3UzdpXLT4IpldS
ChCHS+rQPuS3aYPL/EVk6nOpxZjETb5Z7jyhlVQ8NtbfACFXd8a7hetyQrP54jTG
DOhgAqwuooCiCNra/VRU0leYYHsDffbB5zHJNXwUQQVDkT7JyVpAh0iRTm8XgNKg
zQgOmfTaRIi+j5IyuEw8qWjDDc2U92EZTx1nt2UEGTNfs9yNh3YjImFOWCPC43C0
Plq9wNEVMdkj2GoG9hACU6AcAd9SZ50Fe3eJlAU7f9A6q8L/tQmN0nxZfhcdtqpV
1tWkDJ5b/TYHg0WtwMc355zLAK6UyRY5odlsuYb65vnnE1DVjWVE844RsVsyYtJK
DFsxTIWtlgEWzFYbgxK/mfkzaPXDQ2ZXRLUPnXP/gkt52SPv/aGwGXG04k884Rhr
TceegjGVB49ZOYT+rTG7TKFjRID1QT5CUTieqC/qw1GEq2Un/a0C5oXNsoa9O94L
R2ehAuwJO75V8u89k6u6TrKhwwbYgMPN1T+MWo0ySSXcDgubq7o0C71HvufO/OMZ
O2Hi1CiUzknXLQ0rrFWdYMrAdgoIHhCJV0lmYsyNk9eoQZrFbGhYfcBFMyWF8W+8
4GZv9FdNQP6NYP9KU/2lWTeynEzjcqVpiyqQIC9p5xYtJ07mvQfEm9+NebT0qXQw
5HE9XvKu1WSn85xljVxdQjxnvTtrKU1gDVn93wAkaoHWxchgrhUiQDnaYJmq9xNm
gCT7j82cb4DFTOYtMQKma0HAuMIQmYh5uKgQxs1VmNdJDQyW5paQqJIip3KYmio1
12VqP6hBJzCjNlcJoJyzTZX0OltlS++/QkVzXAoHEIn14Jgqvpgf/FMk5iQY+gBs
vVoP4QTLURFQqFn/tiP/0sjCbZoTwjqQvVrqz+Uc/BREH43pb0/qGTiFpvxsatUe
mZl6UvJZkU9hrZL9utEym5ivUhYPVf2MKbqJDj+c/qFuWeduveOV77snIOLlLhJK
lUiae0kuctZBtqZ3r9TYVHIxop0ajtlEtmdnpifA6x6hEkUEKcQ1cXrfuRK+eBOa
3NTqF6JdLk/2xZrb3/6J7lRLL7Kt8h6dixbUkZF8rVPOjrpbbVj1pROHUY37Xvef
VWR6yUep1FOn9LSV9I2+wj7e6NG/O5XWUjFTo9fjCIwsx4tTrha3LYMNhLd0ut6d
3wVkPIkONFAIuCuPxCTzf+GW4bRW582ayU5mBssNYXWddMnEzhetc0LFBOQpUzLY
nFZkb6bXpOQP6Doz0ZMRzqmU2SRfxkt1NyOYnyHMsuRlHs4kPGdxa9B/RGhktDW8
+WaXVddB2I1J9p9YlgHq6xpX8/BELyPZXeFbLNFocZrM4XB6nrrT+xG7+lWQe4t0
Dv3/QcWq/9R60R+5/w+nYdHrYhZZqyo4/rK7zWUj88KA2heLC1D83FBo8DsstIub
L7xpdRpMokeC3KRuX+3OMs5xjaCrg5ctWAPdr8LMU/aafjMHL9fKBZ9uNPaQB9j0
dQEeOhvEhwH2kBVNT0mUYUTJj5N8jdA5tuHbjI2LlqASLlpx7ULv4gze4DeOMKHm
N5U2izraMwx14ilP5ha9oOzQMeB/pes6hqofn86AzueeOzCIzBmcAor4gxZKBNLH
KkeIo5FAP8O1vil9PnFXkCyIIZWAFAUs1dzp9CrsQYpOCM61FK+kMpYjgCPFNACz
Hk6l5BbqumJiJ/ErQOHKxltF/LM0wG0qc7SZhgMF553lHN6FCpGgVgzJ9UQq3h0o
A3nWYUHcHoRhYh8WiezDJiXdmSyFI1HKVrLnvaza3+JHmOk0lnAsv1Mp+FT3SBJ7
+z64l1X+n8vdDR6MuQKv50nxsH/M/pMc5kQeRopOz75vGUJPxtD1G7oR7z47kbMb
i9EpU/Lhacs4iealT/Kgnpf3mV3BDAMuc4rSFVYQTUh0GbhCpckU3YSesBkC5fXq
hzw8mEpvtK9Suw5SotbncG5uyNLiodG9ZiebIin6/yOoTXbScTJp+fXHhmYbv2Qc
4q1CSgMV4bCz1tFlSmdLNB18oHowNoDCjMEdoAOdzZ2BxSwC00Bv9u3HKnI2P4l7
xSanUAlPsgKGxKyPAa8spci1hg80g7jamTE5USI/AFEcNJkdQg+L4KImaXmJ99ZO
hjJj3U7Rm6fPNd1EMbe/2xA8fhc1zdZMDXIqTRrlA8eYhgf1OzPe8eFcY5y9VxDR
eVouMRbUenvjsthzZDs/+kWuLaAO4WDxIzyz1MmNR2zg67k0xsNHeYQqsGzjhxlK
lHnldqgUNrYWeZA+Dc5AMNQBVu7wlh1tIPa05sQDXAJt8u+PKhQzSJxFFb8lYftu
0FLRHldrYDzgRfGzJRIwaZG1OtMubcATJmzwdegEnVOtiolV5OjQPcUlUeFmVlro
vX8YDZCrCXRkXCkQ8Fn5U7vA/ExVONr/QTkAqbljpOCQ3VGNDeKPiPWjw9dToWrn
o6yTNI0QagO/2oZoVoSge0eZEUFdqUVsWv39FIKPwNRDlPV2Er1QxkONzEbG7RAe
qVl4qqUBxoGbmhNPzQhS8QrEGqpi8svQ7bVCuAlNPZ9gtmNwaaAorncltQEjx2CJ
Vjx7HzHfkyOMqkrG4JvA7buOBhfMXKbQAo2uhpvQshNEtU1FLkZ+8Ah3NK8B1bpv
e598r6kv24FTMn6aAHWtF6rFbH3fxbUCLOSxGENffsgE2GHGZtvg/0y6bEof6GNl
TsItlZDU84ZpwLgCKqqi2pNFty4eoLz/t0vUC8INgHTyLVETkzRJNVmIPJmCdOXK
06ouR6DFzTJyuXNH8zP8kfgfeFsOqdJMb9MEAYIvxZ1w9IsnQWAgz5iUW+EE04is
W+fDZPouGxlnXKVRAD120NtrrNKLRTIeRyfWjg3tDYfcjkKAfDeB2paqUQUaO/53
K+lQ4bVSUcVTI9MKDCTC4xUVw1223H9cbp65LDh7BdbGEyrO+OfcJIrI/YfyzDHo
F6eXIt28d79iKgq6DixuDm6UsjwIs/YG6LlJiyppWr8fJdkmI5qhhI38UTfuw8JY
hKxWK7owFQ393VRgy1EAcohDBmufUgj3gasXKIEwpkPLnS+C08avyZ0Zz6cdYMKD
ot74HIjuNh9FfEIWQU4WRpeg8OaR3dtkrAJg4EBXhm42Ndns7mdZ9p6uf2bV0AXe
dviFC2QYeVUIKUnIJkiy5pYW4UIXhvpwwwh/8vFnbrT716DMGQD2IVlTZ9yJYB4r
rbWiI2kVWP5eC6c9x8xxGt54G6kP2RRJdHS5y7y1xnxpi+RV7xO+iZq5qpFHfDOh
MaoFGlqSQdzR2+SrmBJRS07dgirZxfaAn1IjdE18lkIRAAC94hXU8mMsdnshBu+b
AucOU6gfycz50pJjqnMm5iZk74kX+rONo+dA9tW+hdkz79oXsDzhKWk/mla+Yw6q
fbJ3v3Ev8wGNtsM/rxwL/0+niSrGzCzXc2UJUkiYuCImJURJ7PbVhqM6BFAuCwh1
nR4zOyA9qub3wd6xeuD/S1nuaoB8Y4CbUkxSkbFSYlJrQirbdlT1bIf3RlZia3Qn
DU7ZIn0GAY/17uoWjFOs9enz3dBw7kcrBiRY7lSWCc9OitZgNhrls1jkl9sfd7lQ
nyNc8yI1X0cai9LS1kNLcPDO1oB2UxdsKEi8diQoH1bAbPEXGYJGiLjHPsbhH2mw
m0vmc4xrV/jjmk/wEwc5M5ohs0L+6AM6+ba0vyZIpHoO3+eABXoqMn42HJYvGfW6
/YQJOpUkYQ8zaH1QayqvYVs2l/cdUeCuhQlGfvEgsYn7IKOE2qUO+t2jGfvWdGke
jG+sWjpxp3mVypChvDrvmWhu3HaMDSnfV+P8ZPr4H31fNa9r1QNPkUeFsDcdJgNT
uHeMfIJrlmP/kH1/hVhHk3h829iO9YhlGZjveZ8YAmZsi6kBQhTUAvtBIJF6t9mW
LzsuxtBA1FKxanuRUsHhzuD3mbE2xgqQfDj73G1n71KaWDuCQwKDwZjiSz9XkdlL
lHK4426MGHwHulWEpn0pF07IjxTi6qqwsB5D7Dlcug8VGoclciAcoudXcwP3sudq
iKEg2QrJS+2ZT4rimzumfolQYSknFWFlrLPQXB0Tlw4ZFc6+vUV1ZWLzlES39A8I
KpbTEimm9I0LFLih83efz1Hf0gXCs7+M7tKDVcDq//TBqwX7cCr3xukBfP3thqxr
2dGB09PFcljLaQRMm45iah+DJjQQjOhLLTjc778O+DweNv5ltypF0PwncMNqChN8
wFnK6YhyBat7KteqL6MtoHKzo5nnIHNQd+JaFt3WDegsrEKm8E9shklIKhvc32EY
fj5eDkLtCLnu0t9vnKUU2lijF12h5pWkzDYbJvRE/0UXENy8s29kM25Jbalssay7
VL0x5u0Fdh+5sYYLlxT/AhxCGww5K2EYBhqqZnnLKQlM4nLvf2V0Ap5Dn5J27CcK
40Ozeys/IIr6MrmqSPOaV2jung4MdVclf5ZRaesumj82auy8HrWxxzpg+/qSEzIF
hcQy8CdeMV60/w8LnyHbKKY05TsDzEQbYU0K/D6mR4OotOi2ssb3H3zD1QtNNme1
LGJedxm+BeCQWxHrUSdfpoJaBu717ygoBSOxH0d3TVe8IgXUlfeaDjTMXBLsAJe8
uhB2i7/l5oQMZtln56rYxgc2jDxGq7xq4Y7/y1FFltVvPPLadNLNi5eTegBMnvT7
nkkLxDCCflkFgZmGEEIvIw7BpKTKcGzgQunZ2ZPqzrjsRcF2kj7VSgIYjLlgNGhV
dp29AZ5cH/97vRvSgQfJ4SGfNbNVFYoZjGjQeOqr6X3NWdgBqKsb39cK6E7WuL7t
fo3rrK0tamlOR4vGke2yxoWkxEB0Hyz56xm8xK6Bc4K7LuCLaxy+nIsEHK+MdWWf
jkcOfxLroSAgT0Hzh8HthT5/HrgyfFRysJiLhqEBZVczDLuZTQFus6kR+kszyIU1
76fGIbAWcKSwoE+lcCe0Hleai9D6JCeaNIymiwlkhTrnvGx3/Veun8uVh6IW7Huu
DLOdJjfGXU7kBjXLMDfyI+L/JR1C4Ii8wKtkr+0/ytKJkMLz7xJ2zE7ndE/zvzDR
amdVw9ZEN5K8Td4/9ZOHXga8OiDqCvpi2AQuS4PBLGpNIw9mce6cqQDks6gZufhG
s49UWW6L9PdOfnNehPHEqNa2/X1WyZqZISBwahjSy9oaTeN5NioMBZeId++oVen+
R4HY4DZnWb2/bgIrKCkuawsJx/bzvgzwqWhjU6aIHA9R0OQFgwtVJeE8MhDw0M4t
XnKXuzLzMzJnatP2wvNacr2POW3lHxgaBbO55XjQ0ohOS39aXU63cCNU6XBH5YsC
OpZvt9gXbvyWyngFlY+T/6HLSsF5YETnAglntye83fUBN0Y3MmoU0eI5qSfsm20Z
aUlOgDi70ybu4u6Em2ziJvjQFVauISxKWxIH/aa6Aj0T5ZuJmQmN7Ga1Cb8oz7wE
09NgbdRIoK1PjFyTJ2Kf7JWn3aVEQLi65d7gZOTlIKTr2ctGUeUR7G+QCZW6ZR6G
Kh1NBK+wPpqQ/qV1+gZO+hjwAMLnEAAa2FmcQGmcUdRRMxqvpBFFhMZ1EWQqh868
UONysVy97t4KZqnStp8mTw+eJhlIy1M41ruM0do5YYDP9ut73eSKdp490x4MSSP1
/zSxtsZFMIwb8JWbQbZKHWSwVpNdOWrvg+haapI3ipoggvbpc3ZUoK3wnIuC+v7p
LMKRTilMG1RSZ6NqxKo+nd0e9gNpx2MDPmA53caGQSNZrzw/pMePoWWWcCml/c6j
gSj5dpafyC3CnaKhCsSO9TMc1veTtd0NswDrBg018I8bqh4G0LnyySDxNfQ7PNf3
CnhEPcwsf13UKnuxaL2xzCVRQfS0q8oroopuPHrZyPi0A/9GuY8x/VbfY54Lx4KF
T/Nb09/8ZGVUiSONTilV9xfwLW4EzY4M5cHxMtTOTPcEfawo/l5OdUGgOdX7g+R/
RSGJ4mYfPuIEC7YcPtTXFaUBnmJCevsmmgKpqZWnHK4XoaExYLv30QjBFSkfZo0y
8UOKfCYZqcEP1AvqGOAlyZ2UgzcToRFpTe17hGegY7RD4SVVOxv9fefrUweQ4g97
G6hVSQ0UR4vMCZ6wRfbeLhBGFydOH4wMxTTToiNfhFocWpFdiy7UIXo7SDnbMTBa
ApXoQ3lFhWK3BWQw4kgQR8Q6d/WT/d8P4YeqUIq7ELbD11p00rWg7aPLNZB1XIvC
5Y5S7BjxNkJclt1e6ZGO4vpxG6nFfZYAS+25svwgfV5T+/BKWhUbXfV75AgGcgh6
sgwT7o0ufVoBOw/N8kDYm0FyWwDFwo6SnvFiiQBZAoJLAu/wjHEXHiqVyjByoXn3
1swuj/Asi6dCr12aCFQeQk4tP+LAzB1l0nAvbjxpJD17aJL7sYiivlmdWW54qTSk
RNNdoqYWQ2R/e73t0E1aF9w+160CzTEKobDjgKC5C8GYv4qkxmy45+GsnB1Q7/DM
BfhFtkgVJ9u+6OnJKMEf1s8ZwjPSLAcUZnucbOm8/X3B59j74FshHsIPXepDjFH1
8giPEC0dRNp2CWyutsn4lwN6dqiUaFHsle/4yJVwaKgyOrznowsgXo32k7ihLNds
uqWv5mgM5g7KJeY0pBde+JIpd4NI2bIPrzRXvjZZb5VisNtjwoMb/7tYXaREyLsC
XWCCD5r/yfXInjxNdhM+chi6iyqueZRuDv2fKPmSsYPrJm4Fq2WYS1GqTe80Ok0b
PWd/tKhMfa3AsSvMpBdL5MlMg1CGNeLjkfTF0YOV+55f0mSYTZqMjFRJHNfAbK6E
JCkoW0Dp7Ol7jvbXfM3V33BNBz/le7GMCjRrL0U5Z55CDrVfJscWUq0TDFovJTbr
GJ8qCMoSxLZAeulGWWKPGLVqfzDTNjDGd7H2eP5CDgX9nwpsNU9Lb/GgfLUKgdXy
5iWM882T4XPuWJ1R/fvYjs9SV1qB5SCrYLljgDB/oH7okW+z9wa/emU5/K9zuXEZ
P3dfSVdvT7xa4QyeRa2zRuwSvrKwgoln9jOqwRYyLoxX76D4VfszYHZrxwXTE8WV
i+l6jekO3PNaeR9RNfo+72/7SWwWJDSlkzZrqFNIq+Wf8nkiRS+q4GtpyR29frDP
95yaNpnw72w44eSQwMc9ZnoINfT9Q5FaWWK5sHQZU6E+IX3GA4rzOrfGZ6ifT3gf
Xi7yi8N+Aeq8Yqhd4nA4gD4bXtyVvOUOu0CG606g1CIQUNpAQB45+j9agBgMyPTx
ZF8rpcpWdVGvg9qck2QsZ6+QPNdZszirI5yJoHxxfaVVwtk2zyaXuTUOOc8ASYBT
71huT2TQ5EU0OAmLeTHCeu4khm90OT7vHmIxfTLdkTU3cAlceJYLlbq0Dpbc+KG9
hD6BmDEdZCQgiNmCGC9CJ4MgM2PzOwltyffXvum1FggLqydtGUA1AQbklaZGaQdy
hDrUmKJUte2SHqP9/PQsG4SdimpRKTzFs+ZP1WHmYt4EGfPVZtq1owyFTB1qmhm6
anGTvlzWAhfmtUnAKYNQrHoo2fOzqvyQ3ijX/2mT30wMDGOmx7wZ0pB0/xJig/Ez
xbdvMYTy7ZUSk+pq41ShhQEJNF6S9JZ+eN9tk51LUCp4hiaeynzDzNwUKVrKRFVL
fxD4P7PE/zwNW9S0slG5UE5sIgmPsl46oH6o2VeTmPSSaf7xlO2XDRKJRnz9B8ll
JxxhBzEzNdIznF6sh1gia5a08Js2K/2DdbyRYngbRbeUP+yBxy2GtYqg1KoIcrVg
FtsM2JNlNZT+OOtmB+gkVErM9KfiHjBb7y2jdlJOwltwbG0v63gzTeJFfNZXXIsf
QpX72QCT8l1+MLl9Bmal5kX/nPa5xqTAtvifKEu72X2x6Cc4CpApO8DMiUxVS3jQ
EDYgfziZ5JYu0RZ9qee3kUU4iQZ3tfGbEzu0B6ub4li6E17dkTBbZpqP2bGxzugf
sr7j4cHeRsOpBWuVh+kNpYkNqFCNdKr3301IAvxOhFP4EjxoGg2FLRyglGbX1I5Z
WlOsxu00Ue6Yu2sv96pK3lm28XaK7jBYeTrNIYbvXwwAvio6WyhirmfoetXg8K8a
9ZUfE+HB5O3Y+lnof2GgOW+4sCVTFT+hJlt79T9BkK4qO9INcmaH9Sr7RdPSrx/8
OzRIMhEoO8++ntI+U+JdRrfyREfdg2Qt7GupEtLVMWs/VHGdBK7qH0hG7r6/TcpE
GExK/jORoi4Sejea50dBX3ZY7xsgnpoZwM1ihrL5KWMu7S7SKbF1QHTX9Od/+ONe
fS0AI7wpBy/C2useAvhuNcBwiXk0KXQ8eCPYilpAl/abGpBJYIKmwkuXb0wU1aAe
BAId0v+lh4goH9fDG9k6wRTjZI2ZF7U0/jk5l7oJt9/9WPikTrwXSlTZ99gHCbEb
k25bJBiiKhEodAo2BCdTwmv305o9FeRzGZzQ3/hd7FysPqpMOgPowP8skLZEoP49
IDnot0UD6JPLiMnMjn7MVwmhaLFaf0KprvfC+bDVeLGm+txPoX4gb63Ivut4Di5k
/jypvJAAtC6mMYEXr9KBqZVPrueyebebVjQfpHPTXyM38GWFWw0MLYmKI9MRwOho
D/eoBeSnSDD477wHAOPnw/Cq66I9N9GZPxDhzJoZzEEErpxbBpIcdyfDfr5PAHRN
vctBKLIrnvivx1aOUiLGuHqj2IU1Tcjsac9fntf5qHLJ7cejCHg3hBNQlD7QSAK9
nt2lu255hKfZYVt+F+epRiPrdzGv7GhS19EWhK6dItYc83UbTU0s8Mvmc5QAvo/L
hsX34RASZ3Q84vJdwLLIZEk6FT+EaoauCU+zr4UZEMwZRCbTyiH7961GSwjmih7y
d2pj8yeEmOsbHJeLe4t04UQzd0qM12+U14BolYE4v5p61PdM5MdyrbqKnBq57kjC
JfolMYMVWyFxqaBn7N4FJkgaAXZE3PeMUEPvgiPhYo7bIc2+CGSkUDCPX8dHglqg
oqR3A7ogjQ+IR6MPAbHQop0F0QandmscxaEwNmnfuf/VXSpu4NgUolXaRgMekZtV
MmjD3yFo0UbDFZxD11wVSMEKS8+k2FVCuptXKyeluRStyPtgqZXpdEJyY5K2rNZN
A/uMFfrevbuU+16xCv/8bqa1EQhVCXcQ9zz4ygiVpnEptcF0YbsDBMUTubp/ANds
YaUL7mQZgNEXF/dt2R873z9+y1LYuqhCDJlk8NWcxCElQvNjGCwRX6G24S7xC5a9
AzRZp/1vKbRdGFSWC14Rg26U6V2w2jY7YOWCT18iKAn/1OrhpkjZPJL1f8OCRcGT
wR8S3vOatz3zDErVHF13X1JrkXcNFcV4abnWiCqzvbShoMUgrFYQje4gx32cnOa+
yJ90KeIgzEnUZbhvueNZ3I1buQloive81gt4ssk4P3IlcYGMtN/U6dju+aNYPlni
lYu7n0+or+NDbDRmwYpQp1e3H/w0C8W0DW4QXjsRJ+hO9HOxDWX0aglbW0CpZfOf
ywowmh9tJkhksMiVI+a815i/Zq8ZTr6Tx2m8M/vXzVagp817Ldw3DVwOS2Nz4fZL
7H2sBkxfPz//NjjhSGs3Val6ctiz8iQymQvmKwegsGzLfhmr9wPoBlLxjalUqW2M
VA5OZj5ZuRXfYuJmbQfH+I2g0opUwgX/N8tw64HOoNj/EaF+JX4ZukkesoN4CixG
/GTkuRPK4bt2AfK115+FAGIlzu7bPjn4pshK6va+FsposBuB3HgBT1psbUrKV0sT
VRnHRM0VPSHJ1bNLSgTXQUsPIbFz7yXFPfJclh1bMzTh91l8DfTPcmTG2W2a2jum
yPp9Q2a0+Y8Sb1nONRNJOcoqdOYYE68+wQlN/xAOXQzie4/a66WmB2y++P0qQBlQ
GsLIExdOgE58zlRiT8HrPvD+JK4wFzyK7llqKI5rJt+LA0eFM6CZOETKPN6gQHQ3
UoA8I7QJzjeHOooKUvfiqwYPcN5540KtKb/z1/25ycocAYdf1207ZFQBDQ21gCg0
79PKquNJ8bS5UVaB94vUhlMD34JuKu+W5eORDYWJvO4UZd2AIhmrBi+d5qQ/v5bm
B2c2zCtoOu0qIqujqMepnWt/e6Mh4z8TfReF0SV0LbctL11X7SvoLDZYA9YgBRxS
SZFgGULjOksWxUa0+VGNCzp6QD029fJWHABWes5AaH5Ve6E9u3y5ChEN4FZCfWKk
adbijY0QzaINd4SWFPKx1E+rxgQ4K0OFgh77SCaTdDecbmoXtEjDQg010UVkCUz4
ZFe9eLw7/9uqKvs9lbs2EwV8u8seXrDpghlZFu3WyQv7bAzUEGbN97O/pBDKifj9
Ucl7l11i0uI+MMD5PFxIUA18gmXhnTYu4+Nom3iXzNSDKKk8MoORp4y0JT/JHMk2
OCMshPr2MPmvOqnp/wuMm5qLS74PMsQj5/MPqVr7t9a/6DLSKHOR0RnTcTrz3pch
4wf0bUYzHfCuyeG/eq5zJ227vwIhAAnJ266YRYFvhTIOpxtIevBXzHNg87FmkCoM
ErMMZ5/M1NwHGJD70Jvl8wmGcp0xulwGBI2Bf5IqD8NPHmhReDz9VX3lS2b0LX9A
6Vd9zX1sWIdeZ+uVU4HvzSrPgEXKghqqn7mPu9YeXOUUtZUbY8mGIejqg0tQew7j
x/Hq3fzwUGRg2WXKJcQ/TQI01ZMu0gLmh+pyKESCYw0SJdHUzzoi0OqyvGl397cf
nggzOJd9t8GD2G0IS2KSperAgWWSzMJHb6fciop4yB7yQz2157O1019gVThQQr1s
GK5SMO0sZzmMU6BF5KcpMABKCAJx3cqu/zB8kzjuUc3Et6bd1PPcviDDZUtFXMoh
9rA1yXtpKEYROul5+G7E0vwtzAYypRF2kBDwvG2yIIcFlus+/WY7ZfAaByIUbDap
dca1QSwbWLqB+lyQwv+tKJTor8NwGIQVosfbD7h+FrRulJaSOiX+Jf/9j/GmmhLK
jfqMD69bjmBmdKTWYzABIRVNxt1b1LA9mt6o3+zXndnNh5fjbXjbWTKW3fOVSpf9
/GXo/08F3arzNcHvmsg3ic+u7ljjZ6CekTvrHQevA1ChMhX0sg+BFp321zkZiday
C9yOO8LyE3wjv2+h2voaE5NkJqu4Q0iCmtjsU0/JP6zXQgzdSsSsX/wGtVmZioZ0
CrmIWgBcmJfTRqz1UCXyVtXbe/iXxBYnn8LGdGazpnYWA53B4x4uc7saxPYfvzE/
f4p0QB+NSd+yz8wgpWWk2nEdzJEFwjZjoUnpvNyHKhnLsO1V8vALj6wp5MzNYe5Y
FOHy+r/zm31iry8QoI9B4h9rDBnVm1++tkJgyxSvNbuLuCfbMjq+Yiet1Dz1NAYm
tWAMOg08HdOxvjYv32xt9mq5rF3Gw5M8ex2QarxPWQHaaCFauPliFALDMagvsJ4x
KAqpyBfOMrgJK8AM/5BcyQG29s6w8hbQk02djAk0Bll8s1mL7WY5C+G7BuGKFjLW
s7wKqYbdjWH/Ho8p9o/o61JBXNJRnAWmYOC5zKznpxb1rlswiJoGBPC8V7RRWgbz
0RS98HwDLMRk4Vp4w+w9kR/bfVqVtWlko5MhM7ysWwKXNNGniV55WCFPddx0FB45
7S8wWM+9BBirsC8X1qnnJv2HnjI68Vx/GPM4NXhS7j3K7/OKoPQdcRiNCjsTzYhf
K7zx+OdL7Ae+riiieNHVUW70Dqhy2yI1sZGjFa0uihFRIc2UuZrPCqst7WXhLmXk
pD2X9Xo+WLCec0NluOBZLNDL501y4WIeL8foeJJplwSWVRy74OPntyzOkjemGRS/
lGCPyCqtoTHHjiRozo7d3ExOSPKlkr3jM8T7jqNWGtyxdGMmkTurTf70ASQkR99U
cgFey/t77YMmKCq07Jz4/voAs/Lsp2pkVrvvf7Y+fawnSsx34c4m2GsBlv74hy1u
x0CZmtn0GgL6RG0cjw5/panqOAnYzBLn6cRn4QO4I2rMvIDJI/vtTXKAvHDJxrXN
0Ptz7Sx70ujj87MVg2NV/Z8oNqwBFaXbESjIb52a9Xqu9VbMizxRfewkrZ7kMQNb
WvMTBWC6OsnNrLiXkS2e8eUNuK7JfyrWYWeMGhsj8hOs2NvjXV6imUJohZApJyF2
TBBUAqEq5q8F2ShVCZC7oenp4GdyF34d4jMi7vZJ1Ww4ivT22thMqJ9G8lAEUPGC
phFOLp08lwmLQCH3ARxF0Rj4kKJMwikhAg1qMZ6lEHMdzR6sBl8ZZS9fAw3thg3Q
2Cq5EZEISlX9/Y3t/i+5gVa27iPQDFFi1lJeOdyWjUaKZnoJZnrAiouQnfZ6Z/ax
j7+ExAxmldBbEJMn6zxO5NoAXcwe3pqtW7c0sgqiKD/Y0UnB9WkMaC/onMUUdMc8
WZU1GeLtIVlKNv/z+tY6MpwUxCvprPXKnVsS1d5dZ1FOS6ThiMtivlh/8b7UvxEr
W7T6NcPIb0DLU3eF8U2mwqg3WCLAqOzzpwvtGTgCxBUzOYD1TpdsUKZj/jUsjtvR
WpCR8O+4YpUMoQmoW2YZU31IQyH9MDjg3GQIBCNrLOI2cpLiS660H6oQHYm+EEof
sYqbkEuXjlcHyOX3DZn0VuyKBCZYj+kK1pqYM8aZ4x4Ug4oYF3ozgWoyubzC2UGD
us7I4ERMcbYia3HkAe/lghcoAK1gS7z2g9AmdZI82yrZpc2empcn9Ptu7KptfplV
QryXRF1IvS4tzVsLJ4GJaUpFdz0+kbO4iu3qmijjyYAaKc81t5luOth0lNHTnRO5
lDXuuwyeluAqk1jzeKZMwhiKm2Q1Q0cP9LXBDC3tbIOA/kVqdsGvdsomN9jrsAdS
MhdzxdBuGp1VvMSfWbT4qqdKI7Un47IljGfVP/UUot9i+a+JxesKQf9vmvCUU9fi
6IlAiw3WIcTXGul9pz/D5AibGdWLtDTmIcKnXKCxjx+PbeT/P6ysPybMxGakU9Ty
t6eOUuibhiB0WQVnO4c4J8xxPpkpDAk4c+9uf/kZJ5RRT2FchSZfhaUc/rVNkKCp
uaH4HTiI3SNDISu8cOhfp4P2cQqiO21P8cb+uaY/jONxLTPBXt2Z57ZdbOZa89Bj
Zte5WgsaEgbeOCfdBixtepJbyf+sDwmS3JWdol/okyCsnLo/Dx7kFikbaj32ghOz
iyNs4iXA4YZ5hKjAcKRLkwrDNE4JcNSyVX6cQNFAQHaiFmzQLCgKQx7kX0R0xZlC
xpjHGGUctsxOiqgtLNAD964IDZBmCvDuSd9h0YWnqdBR2utaKhjiYhpbOdZQNnwu
k6mZQ32y0/BGbO7fRDhDBqjSNbWfiNlhjv8caKtvXsTCZbOjp9qJWFilcI5hQJ6x
X5tL1MAbK36BWQ3plrUdlmI0dxANqruFvYhEJVGuuSYhu/R+v565iv2n1wsz8otl
1EfrY7PFy71Ba9TBQh3be+M0d7V7uwV5K9hNbgfYqmn/2SHsvYAgcFv7hnmRBFTm
g6hEEnEFrqAE84+WNJx0Urw2jOvu53+bdNv4BWCSMiiOSde+xJp4jvhcdCev5HLn
vRCKioj0hmZ+11frltxVIHHAGzc49iostA4noHyW5OV5tSIwrjPR+npOvTJXR4eq
wvCWrh7MfyCa+5RpVAtAX2T6dRAGM9tcSlQ5a7GAfOtOMe9y7Yh7aF6jrRIStVt7
CNuzUztwKnkYn/758mCGWvvkNWOxUkLpVhdI6F//Uxi3M3X45D0ivWuVG4eMI8Rj
7wv6qrXwAnpxzYwl5NCgA7j7kdO11Qm530RvbjjY3yqz9lXo3j+mJhYDLIREvSBk
44iiIetPNgHOkVnAypn/XQCnOSoeq4MHFa/CiptUyfPi63KnZ2IblRtndjX1RygH
+d/+vmx706R57vrQL+zd8IJrMpPPuFbyy4a2Qge7lYn3FFujMEp1XTixYU8vA/wQ
flappVLEzK6ueZrLd0s9MI/0B6INzYF/NNlNy2ufEE2YxW36rgLtchv0HoX8+2zG
mI4xSY4Yze0k1WbJf7b1LsQ85KJmDowYlWBcZwEXGTtwElSkAzg8gJ5FElyQ8NxM
En0AJJwlBUE6Q2BPshoHdWE4T8ttMF5MUrHO78j5UesfVpKRsYsmosz3NxlFbUdv
2doc3o0mcAUI3ChPRnfiqPDVmVG7fXxbzLZj3Hl1lt6jTDZpTRqRhB2VJwWf+IOe
AZnT0ILrHk3BcurPGyc/WL3OO8u+kjMqaxXY9WCjO1dwX2v7+2B4UNbr4ScZ1QID
p2bw65ECSBfakuv4RknHQBqaiv02Nhu4/1ZBONyNFprD7kbEDAh2TTiG+Fz6Rt6q
AwNcdb+qRVWWBekaCum9PhOYd/99V4H0iOnP4peYuK2PpCkuhtVzUFNPkhwYPlxw
YsHJSIQUT5MjYyqRxsMrZGcyRRw2rbBNseL7p9ZbtP0yMD3CYdvXLskxQyraD3eg
sypPAOVf5V8Sp2H3Yv/B2RsCy7YgETYicxCw0HM6ryg5KUZg0FikHo1Fjgk17YDB
yvUBjyaKXqs3CWz2rABvWUw4U94AvOEc8054DSGWNta35bcSW7Zxu2OkjylhPEo9
PnTLNU7x4AADJXfg60ndG2mAzo4Dl4a5CPNX8lrUwNefdS4Tty4G6LafQXYSy/Vr
8R1DcjVeaLrigVDwkHY4v9CbSDy0J5O718WjNEyH9825kSEBfoVHFfKiP4WsY6DY
f/k3qjVf6scBtghVdMdMYVAYzUEKA+P4DJVeSicWrVenMY4AYYRif3vAp+1GzefG
oxl9PZCNHAg40Y8CQPUn7SbVBmlIGMHA+oWTuLc1BkNM1YWVq0RAuNfnb+4dv6tI
von6RYWMmLBfbmIorbnOS2vUhhSNNxjSmRjoEYto0CSDihYaO1YzGmY2G09teBol
gxE7DmN9YXf4S9fgpcvHoIQrhm+tkl5qss40o6tmQCA/IWLFgdnyKHXaAtQfZIaF
+5wwFoqTyK4A7gKFbIOobPrpkR9zIAHOlI9XIi3jp3yjIPEBIiTARFi4U64vwoGe
EjBLJHipMBgta4meUupGcq+5zP5hD+9wZee7vSSHC+IOXq1l7MfEztABPc1H53Nm
BuHScT/SbQGVbjAyknS6bcqFkwdchh16c3pC/I3zn3o+oQHTNRLr5T0DqNZrSXot
v+qgNc9d3S4zqyo9tN9U6sQXzLEROGTFwZRhBarnI+q0PDaSexzTl9uiPBmH/ILK
SB5aiGOJqVq534T0o5dSUWseYf8bXe8j1TdX3RwVPGS9JEKwVBLl44TKOVW/HAyZ
vyi101KBC5y6l2Rqw5ubftkyeUpz1uUaJYMzGbWVRUdZETNgg1JlmRvuQ5NquVqF
I6lfzJL4q7GNt7LSn/Y01gfX3s51bNI1UjK4NkLhEvNO4qFcOsR+TCDfhqUzSqrZ
rpeen4CCw8mR2u+Zzl+lqq47ubTFKxcmA0oflmXdHqDBWs8Cd7zSkO17/Ivlvjwl
wp838VAGXxyfO6k1a4ZA18zijqgq61JZB2Ph2J1NHbGcp4r1JdUv9xwQd3gHG6Hb
Y90xPT0pnLRU6g/POzROARu9dXA9orF5glkdWbuEUQBSQn7AylGIbuzW9B8u6Jfk
C0QCAxshhI+HqHkOr4KFMSnwUfOxXGoHzHudi/jds/SexboEOG7MRFMJCcoI/a+h
BODs4V3Iq3T64bh8obRCD0L7SnZ6FIJWpXGGGTEsJBwblfE8E6BVYc/F/FYRwGs0
3/VlFeJbK/EVU1o6YF4tbGGgPVS1k1W46CJnY2vd6ike5ROX5zJyDObyTSndS/pt
4XNUTj4q+A5bGS6PUOjoCQQFRyHeeZdwOT1J8ve+fFM1U8WGwKYV7UZ60JcG2xQa
vEsP2pF3V978p2LVWaoEbf2WW1STvzq7yq9SY8pCiFdN2p1EU/i1a5bYFRCeKY28
Z+LDqFFo0V/HLi62OCskZQMut1LeTA3CcAC9H0Wehc4o5ApPVAJPMBaf6968gi/c
Jdg0Kp3SEuUnEmYBmudI1OQ9Mi6dJPOmJP1HL5IBZVWORvh2BuWaRKMXRUPPkPyO
zRyjwUzImbjLqmPyV2wwLde/mKFypj6U1sFOajWUMlmtl65Z45wzMohYPHgTRl1o
dKeJjPJW0IOjPqzfFAlCpGO6aJQfvQUxgOEluB6w+Mje7lxqtTL7yJEHoLR9qEc0
o1Lp4vaZM2+MRWoBrq/QdJRv88KlMegiFQvqFAxga1Tbe7goTVkYTXFI8aUsSSop
Yj1NrjeGrS/0uEosOyI/HX7EPglZ2fs9dnzSQAAopsbPo1VudrmDpOIQHg6Bz0B2
4p0XeZTngq0JucG7IJQ8Rp+J6zPGr0n0pw/dU3Wl+UWkB12m9/XWmsckjia4EoI6
FQNKA3150o1ClWLDa8SBiu7kB4IBtw0PIa7H64ozIWDyrdfP0xIjbmJvsPgH6UE8
b/aNoLe9S/UztmUr9pR02T6vW5TBl14ttZvnEsyusVFaVg9ETaKE5XCtUooHM1Kg
KHHgHLY/FrbuG8WZG6VIEWQGClzSxDbbn9GNN0YPrRWh4xlP9UeWVjH7Voz/ETHS
LAcePGNfPvcQ8m0DiEZDCFYfEQEO6GqLv+nB2hG94XNFbeDC0GPjps8hXFYDCZEa
nb74We3G5fbwJuTtmjLJNNcH8viCTIyOJhTzIh2IrfGmi1JKx04yyEESqS+JkNw9
Foj3UtdwuDZLq+fENf+R2fE2+z95tQBUPyoGv24GG4JmWNJwuJ4gXQir73t75tSq
aJVHV16rYDWODLOT9iCgBOe+EzFBJpbqnLmq35pHZeqz1/nNagi3fc8HdDo6NZSJ
PeH9hMMRYAGd1N/ltc7mxLvipR0zb6l/8aQe585mYWNGiIsh40his2eO0HWhagiV
PLOtV0adLRx7AUwb1/zbTduU+Ip7P1WnKAyGcveLAq5MlzN3dalipPITpSrHN1JV
tnfKMx/wFQk0SDTgHFFmhfFdmjQxFWTdL+RYuGTT1I9OE970MpeEDFwSFsEJwUaX
2fcMv0jXzSzF3oqCKv+qvxzGG3sDh35C8WqPHZmgBYFoxGfL376E0s1IkcPTDA8h
4sQAJk+nxox5KOAi0aLNUvyMBcOugdN+elHzKPp1R8hNxjme/emaphfghmm5Ge4d
ZSezoUbkeWWL1TjaxXXk1acEaJPd/dsgMFwJspHJTj7h4m+GB+TiFqjp+G3sfXBW
sATKENWIt9a9FM7gji5qyWleY6K61jkagRIut29IexVkCHbfedZ++kAQhzCRxMdn
xn+aXuzxEIf9K36eem5yg22Z31IL4o5sSh2DRFfQwvxs8Mngdm7ZbrpW2FDVyXSH
PkBf+veOTUuOaCUwsX7j9xpSzFdfsTqueefypp98hQqy5eluRSruzFD1nIvLTDIb
NLtxZa3fQ2HLBxKv/2e3MBqaekpBR1zU8C0QAvzTd+WLoKZdBQ0lYEuD1DrosLjn
yHxI2rFRAZTjEqVC38A2r3rrAWUGl9rX2hnlabwF2VRPU26dmM0e6TMvCip50LU5
Wg7Y1YJl4IcmMO8wP4A7nhApB0OdufnJe7C0wAZiy92LIeIIfTcICJpw4iAN8YNo
Mh5keok5E/vroDR4ged0xLedE3Ak4yJkPiEYR5PrGF4NAKKfcS8EzDF9OU5kWExg
C+X3XHAdKrgBn7M4LoqeOOI9heRjqgBSc++E75OA7i1BZ7DBtunDRXDN8GmJIbZa
+XyhhQcJ3L/TMdWNI7LUqqAu/R6lzCuJcywzGmd/VXo71s5W+IaYU3/3iUmcy4sF
3infhzxZ9gJgCKMfkXXyvJkYkswr3je+d0LCW3RqcHkUC6IN0R+KIlpmilQFd+Pw
nDZe4fkZv0FmgWYrEJ+sn6By/7eiBLDsG2xTU31flGUnKXOBbkYVBmRAEMb2QXHb
Nb9sJdOhiB8ZoUNE7GA4FhOmew2Wizhjd6IDIvBSz7fZ1gnoPvd7rJ73gQiiLMJI
6RdjCIDkVmRdwwQsloSkS525F7HTiAGjJAp7fsWKeC5KED1M4JiujoAE5WsIwaOa
YyeM77WNGb6D43oYwZXnzyxmxLfVE+eXpJDG8zXi81yvMaGHawqRvC1Pfv96Gzkx
w6lGEIhK4UoXmra2vWv0RZwil33u9rYVNMX+rhqjdTzMrHX5EU8r9tYYXH9uQ17p
+hKo6i0B36MmLILJXzi3uBb1wnN18tk7GSIrcwCvhr8pR9ya1re1iJhcBXQwpR6W
5STp8mfa+3/uLJedqqeAyAULSmeNt9rg1oQF/gsSaawmeCzy+SEqqQQzf8xpst7b
ZnsZ4ywiKigkJtrRxMm7ai+FcxMHbJSQmgcuEMVCe6rRqXpEyVOx/L6E3VnKcQSA
Xx/6rk6DTzC6OQgoWUK/NmMycRwhpO2UGMPK0sHtzfTyzulzCy20zv5trAf7SOHa
xWtfx2D2P6au5dZ1sDlZBToZMttcDNu8LjD/FVOE4HMxS0QlUrkloQcodfOwUrUQ
uh5chyGrCi/tPP+BxmMQ/E3l+2n/hgMvWwyv9g3McxHAmPdu/0sSpOgtNVytCSn0
9gCG/CbV0dvxEwbjTp6X9KoOoXnk6uAlVCQM6LumXS3pJWAwH7tWao2zYARyGCpF
3A34s8gKWfIyg2ci5Uzr3u6KaYOFxnQDdtrN26ViRRDWG5RVwKVd2Hpd+89T380q
gmGjNr7KiqEbJ3f1nG+KNbUppI1OxKmbhG9jp3GCJKvJZ558fWuH2bcZmNdXnCwz
+0WiUmLHJF7XrOez47vU9EEIKu8Emr7/FB1YotD8Wn9Pno8U6utI+Ctr+Nu4MEwa
U4hE6g0M9xVdAWJkT4UM3kkmN7WqragIea3b1RX7AU2CkzaEpP3ATDKiz7qyjN+L
JXg9WTfcJvxE2LOS9WsnDjrb4GxjqyEAxZV+Zd7eBWfC1x8/2+ib5kR/vmyD1k3v
W0Sal6lJNXlLhtN5aYVpBHmC+vPmHtkADXsYYFebJm35ZDuQVbXTrqECa0QalQaO
SVzREoXj4GniK6QR4TuiXGFrr8E79x13BJtj9kiOKXVHN9VEGVrFPffNPZQzMJRy
VoVcRnvztRwjCEzAphDuEcMngeXrk3Gcf0X3VoMRr82lXw7ZD2/MLAgTqCp7z1LP
y7RLthVBLujyl+ln3X41x8cN7a18zog/qDDs28XeL2tRA3Z8IeorDpjNcx7mmS+k
Y5gThOHwpec+lspVcEzbMtzfN+edgz5TZe93AS8HZmbg5lwvFeYnXq4SXFV/eFeM
jHFUxM2C2J5f0TALYWXL2VMHZ4WF8Xf8140c7BNYjdvwGGANQxcpkdJ0dsJ9Nb6e
0txj1CPK6FAY3w7DHNjVeOhwJUPugsdWP40iYRrL8RM9VWnWRzosHVwaIfjHsQ2/
eqIbb9Go9wQ9xq8LQKOPtKL6rLxd5h1PJFbxiM/uzz7HZ3kOYiSEsVBAEkK54VzB
pIqQ4Ur4nxJjWKsBTL78jQvuTpkJUrZM2dDCEiGuTGYmwQMuI4rZjv35b+bjJn3h
tSCTTBcIoKYUeUgbw09IyvQUH+162XiS0P5QzC06bXzdZ0RyJEuO8QAUoo+t7Zfj
Kqn4SUJ8jNzwDZWoKkf2UiJE9+Se3cIfcLEBkruAvGhn1uf6CpombZr69NSu4BWi
yF2MxycYwX+2SJJf4DtJn/B6Xbe5WRzdNOi9G2BG2ZKONNMhLeYcQAtiKX1DPN+J
7aR+o79g44T3ZVaH8lTGmlxxjQ2r8qlhSBh6qAkuKMuvFXIofCnTIZ9KbckyY3Ak
dMME4SmmswJVUYssjIlb3P5IhUi+OBZjP7Hk4uu423rKtSx6B3gazyd5fQQCPvck
Jb5XHlWnvz5aISL/N/dyn5n3lzGuBIuIpbQf4AK5PJw8XHeULZY4FDdY57L3ivAW
CWpSH4+MbKheHYJemWj68769mDEbv5ICFclg28ccF2ExugKfza/2g1D+4JuvnZZY
nKY7VPudG///KJHjx2mRu7yX0T/2fysjclf5yNOA6PH6KSqdN8OCmX2zelGIqI4F
TKVkjeyuO/m1s3WTa6vT/hBDF+rqSGRypsXkrpVfoZx+lA/4oIz+1798wPQS/o8w
DDkAriNx/eHejatWZdkYBTjvrHXSolhM2wzG5CpKwDur8/qispJw6nwFsKdVC1UT
sq53Xf3Icqju5RbK03OCucMwlh9H3vAF7nFlLqFNffOm5iApkYOQg8pp+TxeTXQB
yNjE5HjHClN+doqEcU21khdeoOR4ZqHYZr86ND5RjAP54Ix+gBWJ6JAFcy2bukC8
yjXzqrtM8dCXWWGDeE1o7FJKSoGO6+EcGb9pIPLagDtyaGaukNe/qrJP0dAj5EeD
61lJHMWeNOU+GgDIPVDrtO7y/SN28gxDRXuu0fawXbZ6Gq9JP58gpMy1WHiqpaGX
cafj5PynYhLb5VhS2Fbp0eoKzSSlaDrG91gQ+caIc/8qqPh8faYPZ9K1zOuQUjNB
4qgcAZqSLrnKJC8CUF8sM1JS/UwOT6w+Fl6sNWboMUz9oJqUCweosQw2GopQ5tUM
EWOY+MXwR32P5M4k6Jg3h7Hf8/jiiIg2UvoV4FvCpqQnkOtAf4grzWnbNe52LYPJ
E5GOACgOwty0q0colu3TklJs9lCOyqZgAuAgMKHqJK4YSIuxI76fJ17RRFYR78B7
VTR8d3xVSrw3Sx9PZ/3faSZ6lNN2h6ZntY8ssd8vUgQKtEA0ufk0L2g4BAM1ExvG
CCcW7lp4QvXlMbPB/NJsOFvRFKrzFOaooR6gB6WYMguGVxPKr2+m2KbcufKJZ0Db
bJVCOkQEqUJwvHAxfQCF8TiYGxiYdgQ7cnrh1rZnJGmNh/ntNuLCg4XW3xk/8yN3
yMJ/8onbGRueEzQJ5uhpF67eVPCUcefV5fTRSC608NXdoPYC6I6jOVOfKGuryDlv
54p0PyVOcgEJ5MmuDgdnZPM7ETU0OHWeyg8naSceq5frgjnLWOIDVXV5+BO27ner
szD5eE6gv9ElDCFdRrB8mZXrBNZRnTClZRO7Bo4aY3wAjT3qSTxr+xZBjyz0M2XK
IvmCETiVzIg/UMwftkqu2CvEmt4N1+WnoAMdVn7nkFQKOYYk2OaeDD2XebdLM0S+
IPrqCrXagvCnk0YryZSHcnYehRz32hfPRaD12lwHwvn6WBv1CdzZXpoUoTFeb9WK
5Lc6QIQOZaLNNhjWL+bEBmvb+lpguVourOI65ZnSHcv+OcvkwaeVT4A8+XSkCR5V
tu6zluNYjCKs7vowor89r/L036ZrjdKZedr8qCBvONu0ESp4NEYz8dm6XuGDnG0y
EJSv3O7g/2d6CTLAJgRI1jK78v+W3FHFF++w3zbkJe8yjrxt73O3WfknwhG7iUqd
uECO/RDBzY5rnxSNkVfjZD6B1mHeBWHk9VgDLsFUq2YNn+6ZSmdI5Q3Sr2Q6JER+
dQz6YNwDQ3/rBjrSLxzHM1vBbF5b48/aF3YP+ZNJnegxfZaQT1CeFBj0p8wi1WNj
PtLIoTRtWAiQihAATJ1mJKhphdgWvAmFqrVDuFvOdtHSjpvquS0/IlXeGvLU2OIh
Ne3Y0cthOQ4XyCvtD2RakS6YSB8D3EaqcZW+UsrEGN7xFxsPQDNYlRLEIdAkfThc
6AarC7g2aq4k3fsQ2nDIQtXhSqFOpNla8YuxaDjjEbrT9m3aiPtkbvJCplY6+f1k
HIxaOsfcxzWDtEqFSJuzyL69vSgbOANA4hlV/KzwtrZC82VQjzTrhF1hUPGg+Z6d
IDtgHwnihiUng9WmUN01s2BzC2E0q69YUCq5KqJH+pomiLMzsmqreh06DoTN548f
xO5PLtQ11mJp5Bhrf3C+mY2ApEKzsJwb7EwMdhRnVOXX+K4sXrD0pjfyL21hsHye
W7JpHX4GkHNXtBHcwCA+OzmG+wJKPS9gyYHMUSTmwVnKOOwPoWfULarmJ2czHUWi
+3LRAK2rD4HAz+4HwBCMc+m0vEjdI+W8RUHOCDDULsl7JVRlcrCdl8cbMCacnfUo
DKnvXpLUkoDUGPGAfyZ7JuG5HMr+SdrI4IKlSBeNNA5XQ636AUD4gwVVd6a6M+Cd
5h4HezwepWptQ+iRLmjEbRDh6sbDpf0Ez/eauX2qVUNx/zuZWGmBF/eBC8HvslQ0
A/14uvb+weuAZjgeNsUpfkzh48FUVy7++GFLfbHAJ1RODARAjB8dSGrmTOwmrIwg
kGpaeJFTotFck/RIzBGkdT3YCQhtK+iHMZbcUeWbuCv3waNjXCQ/IdCGC8GibREh
hG3s77twI/XllNBi3yLe2Dp+c1DP6REBOWSd+V3AV3A6l2b0sXfpI3XFPHw+caMy
20kbMDs7XN3GEwwOxmipJdxeLCCM2f24uZFYTBqQiu0sfXTIdtMyGXb3ibmklTwY
ZWK+nlY9pnzoZXepfBgCj+kCj1pBAor5SHEJCP1LM2xTwhkGHs6U1Zk/HeByvgki
AQOy/EvV6SCgbFU2Pjl/+tgr8STdubpLv83IK4i6bV1emtQ8n4nWCBYxHf6ATtDU
DMUUslpvCyB7lcCz+TbUG6dRefjtTDnKnhS+surPptkl+qH3df/N+RL4a3pk+t/G
KzmHlEsqgI0cr3BthhqtW9Ph1sauLJIha2xvQxEPFf46nmiN6t6VNwS48doD2gW1
Iag2gGMNzehddQfoEjiVHfx4sMh33mYb5ufpzdqpuNGirstLB4Oze/0cKom4vtGR
AcHptqgV8pHa4DneIWLAd6WAAzZHbNMFYEUDTzn6bt37a4VJjwVfOxl+NkmFzSJZ
fD5n2Xnl7Bhc9X3qo3sLi8FXXm/N6G7wWLce3M/xeH5qxF7NM+n0gD5Pm9BztcrP
63adbvlbc756h6Y1xdFmd6TWHSONzGnCXk42eSGRjxfRl7pBS7BHjAxpTMDzlXEq
w+jBmlVXDokFAHl01kL/kxw3Pz4RZ6xEAfY9ScQluxPcXdO+MFeiR947Ar7yk0TW
bNKh6ViPRa6FHRukY9AvkDZlY5hSZz+GmaxEB3BkJtGtCh96YbUbbDIA8qYVz1Zq
E1aS0p8OtQjB+MrcbGkE7yzY1VN5k9hq25ZekNiTsilps3aNBWrmiK7IVwCuNO+Q
M8XUIXlNloQ3y/QhAxiUmjHHfq3+aJ+fv3OQ4QEWpolTf88iP5fZGERWgau5Qgcw
PAC1H5a8wq90X5bpJfhVOFbi/htM/1YOuluY9Jj7sis4KBMzw0/yfN8awOf+w5Hu
nAw3ZqTQniBkIJpwMLSGwdRW3hTrgKAMlfWO2fk8WrPyMzq1gsY1maUa7Lzfhj8G
f9WaFyOevrj8Fp9RMG5kGt2++zZkHf5/VrlecfJ7W71O81l+IIW+tuU3H81ZJznd
Qg5taOyxltf972wY11Cj7nZmdXWCX7gZSi7UqHNeBmnZG65bk3ZY7UVupd1ZMQ/q
4K52QC3ZT3e68xJtRgaGM/NMDmrytKBf0IQSkYPZvPZutSH6hMBuDfTx0ok4/7vA
2tHQDyVQk4I0rJL5SF7Lhn6I6F+CBVPIvDoF7Tnp76o1v0D/FnLeHcZZXzUGGIsb
uHx/Y+YCx9I9dHeraQVqkewTiY916HsfdewL7Xpfginr9fVRJFXg3UEAOP4M0xt6
wvc3pot766WjBv+n8G1WN7eCNwU7gw/FFKC0GziGuuJf37kaQ53tDLwcJWXVKRpH
Cm/WpxtMO8IL+zUr5uSblSebhRb2i+zlKlBkNddr+V5vwAoUVDXJy7W8HySLWC/q
ED3AvHg9oDMBkGoAYKBr0ANriwRlj4v3pFRFsZGoAoJMOnbhCQRbuEP9AsPIMQG2
GN9aTKN9p6JZrw5oPB8tu5c636GXiIXg3gv9QBgyyBbclttUitCYLnaaSy1Uhqnz
820nJV3R8Z8EatglyqrgPIKC1Y+s9VdLTxxM2Fu3tdCaWwD6qvXnYR64xYcqK3rX
tAf+2O78Dnoio/jfTrEu4/HoHNZ9cgu4mqKZV0NlKamtLnhiqMDuY5zZhrBmNROo
FFMluv3yQwNP+qS9O8WHveEPBOnPqEJeu4FPXlqcbvDaPtLSei7NwpFgpOShi0Ny
u2j3ZGVvCY/lx0+7dfofUohInOdgxAr6Mi29SL9ImwPpmu+gd/KcKPwVH2A6Wd/j
5ZZzAYg5bjgbGsfi+cm4W96Qasu3Qd5yQoi6crX11XMw29nvp4xqjPD2Rt+b4IrF
dfLAM8LkLn0Pf+CPRamAlJ8X8MlJVa5qy4OSNM+7NHpiHLPJrw4OTNs7gEqhSux6
Y/Fylp/yZQjVGSfGdJk/d7kZRMk3TVUh0MauN5DoQtRFjODW6It1sUxObLnO+Jm9
dBlq2Q/Nj5JoW+XLfNs7S/+1V2AGzRJklU77GjZefJBqzrEMF47BdPCjfbb+t4pN
wU0i762oKD6xQ0V9b659HiCLLjw3+NYW150b9gKr6ZpLmCGAsIrSQIS+yOgoCfUH
7W2aT/Wlx0+WAT4KddDFT+lx+TY53IZGVNhCoIbdK3hvMR1opJwbPo4y+sedLKLP
ply6i0bdUL8UrA+7FB9vWZjuIAbVNnPu5kz/mWNvze79tJIqPKjyWP95NYANlyB3
L0j3J5g+/lmAG5OY+57GG0h6cFv5vjuW9vSj2clMt2JcoE8qcUZshy1zMXioBfqY
wejdAR/k46g7JuFtaMKwmHfpkingEk6wXhldABc3GhgzYqUUgUez6yF7PhxyEw8n
Wwmm+XQli+65odsHCHtG58L1IIZMqhhOXvD8Wy2y8WqWNzTUMPI/fdcnxFoCGErb
wgrTAekfTynBQHVDR4S/PFQOlKk8I9VxSKUQQZsY2IM23YUM2W/w4BVZbHU8847M
56UoNO9r7dNxIVd0n/8iguqS3wWwTiUb+guJxXRlvEDsJ/O3bo8oO+PyWnEFrb7r
hyoDmn5dq2chlZu9QkVZeYXJaf4LNIdOTabTn9gMRoOsVVGFgpEn7/sXzqOw9LHb
3W/9rJD7K4qGRGZdohNtiPVHAQ+b0ocI8QigPXG7NSGPg8ue9z+NBY9ALN98q5Tm
YCs+bu+010474hOl2I0tvGKdmID9L/IcVnK37WA0K3EWFwH+cbolXGHZn4FqMy3H
ye1p8EpYWWykD7REdLLdY3MXvFqARjGNwkguLjmNkfVA/Gdi+GO7pA3ucIvbIPyM
HJLpwDsgU5DTaaq5URY/F6951tTSVcsYsLM3LKsAq2sGPm2mqyHaN/uNgv+bVyPo
rkMhY9L3K9kSI0OFo02kcxlcEq7QniwWM03MG6VQqtvKwio9KTYNtA1IXKkA2vf4
XQHGKAVC9xrfz12xIDHZDxMGA8ftBBawAp0CrOV+zqAQulM2rQs8qQXkk+r9tfrK
x0TrO5+5wrwnh7NEmbkvgbzGyOVbjsMlJFTicCpzHLUIMK5b2bPraripLHa8eaAo
UHAEqD4K9sP8D08afH1dUbVKOQwl9s4WDBOykclzdCSxCmKoxRfw4H+Y+v3wwt/A
BWrW5wd2z1GQaRTlIZjGD2+hcvCV5YS22sYzlowKeKo=
`protect END_PROTECTED
