`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFZo/c5R01DrwmS59mnEn+VufALPRxTIw3B588KMmWgXBxsBFrO/PVvUhGcNM6OC
G40iLCcWcfBfwcNTA/fqQtd+vc9PVrT3pDQsTeSfQslnbMO6+q16CIet1WZV57Cf
vvHsTfOK1np+YDpMhuI4NEexDW6+pvaL7xMnDXD5T4eGv7xVQMFyryxIPOCiyAad
un4He6n2+X1NgYRKaLCrWn02oullH5irEj3OTuwvHH5CHvCTFInx2g5AVFe0UPoW
d27zDXP+WxSo/o8X3XuViwrJ9DttZ8Vq9FewPH/q9S2oREOQAWl3UDmn/ChUd7pu
waG0ZAaRIQJAhblkHX9uAQzRIFe5HqzkaqAcwj0gyHjWYGaCvO75cOb66ZSF+wj6
Xe2oaiVjzh0gKSrxpeTVlczLKemWHRIBcpV/dY/t1clEwARd3vxXPivyImcqOuFN
zedJQN570xhY/XLd0NSvIf9zW7npLcCy2Hz7ZD61XluKO0lPLB5e1laPj2xUJxod
yDF69soqA976+XTKXQilH4lwOIflxrpFa4SQFu5b6QBIxrCj+S1CxKYC2UnPxjyH
DSZQf3ub26F9uY4dPqO145+XO2JQgmPMWGfP9yXO3oZrTEE2EQ/KFW7Erlrx1UdG
tVHpztXSnNncCLxa+jk0W/7ZTxsjNqFsY41vuXg/O6vcmppHxlCc6Q3lJl5EOxBC
E6rNbT74rHhyln11F3Ojb//LB5AR6cql1LidlV2wQJrSgzwF2B8kZpXInD1pG0yO
m574bs36TzxwcrcspP5FNX5hHEYciS+peaCzlw/0LMtmvpzKMdpgZKMtcpFo4Lmv
tZGfSYuBiXA/S6S4bEwXGJjPP1qRrHXYPgoUzdPTAS70Du/YyGwNVmxkiU68F9CW
WXISxnm6WCss791vuQpj05yM072Pr/Rvsi1CBy7f7P16ooXEk0iYHxnU1/4Wh39w
vBZm9c194vkJefwoLBhlg572ZlnQKZq9/XXGvunHASK9EIsnnqbWH3ruFI3D6bNe
xZpnoDBIO0oMFzThWIxaPNdQ1hV3TOPovLrpiydrDcC6h7axMTIqmdghiBOTreSm
a/66ALn1w+G7S0rp9Q0C0U3Ay8QIzTmBevPtSt458M68BHKuERzUWju6J3TxomsC
SChrZSw8zr5nE7zM7oAu36kNXNhKPCcEPsizDNCi+RqUaGWFzqDOHXxu45cVPSda
oEQPfHdAPFTjkb0FaNnPUb1aTEnUbOMHtx2HRe3lDfzr8j0jUoIdhjBEtOqE/LdS
9DDMzSuIU2cMTfzNgmOgTbF426YG6gg7LuokAnb1iWPncSyjylZMj6A/vzGtwG5C
mVt/S+NbK74ypjmQTgBMbNpaBiay/nl1VTiC8Axq1/v62rgggpvl3G9BLDQmysLH
wn7sNPF3IRPUNKiPOS39hCbZVexlSOvB3je3p9His39jgJ87s3VQGyvlnIO3fbku
PChzM3u40WrFTu9bX6cHWUUHD0Um9RBwBDq8FrgWA/fLtqC2iIZ7wehY7/Gf8eoq
0E8VSs0Cgl85TCuupUPGNjYDKDNFGBFurZHu1SCPKBgdyeFW30tty186XQmtI0gy
D8GB6a3HAVbXizxk7ETq7T1PTTsVKsB4N+JDIGqvet5DLA7eYxfPng25wz9RtTy+
WgP+5RY1wWvI3suMQetO9WuBkL9cDg27Tz3Nri1pfvtDUJSOCEQ//IOT2ehbwlsI
LPD7LrdIwVDFEY1CfipaY7Om1MzNmky9h9I1zh6r/4oSXxM/CRmJZQG3GcWB694Z
Bse5609ephYreZmGUTztbV9Z/WyQfywCZPcuSwyPBdTGEtfsUjmXiYUKd7X3G9yP
UHsG5n0IJskepNmC4UTq6gdACuBXdxDb1d5gHcitCposN0B07Yf07nYNiG750LBj
hxq6l+6blAcwaQmen/EKuzn11JQH1FMAksfgX3BM/vRUg1zkEXux1L+7l/yZYJ2W
i/i0Y49so30w9/8ABEWULfUkOdMKJznFC4KJOubR0wJlGbgYV9aIEBOQwrzmlqju
9mPtwOH9nHNJHOEkqJCwrwv4v+CdGfEvLHBMHqajESOoR7IQIBDB2YEbUpvgrOg+
GW9BuJ0JO+L1Gtnf1OXPYdBlkJdjbDrc+E1DufzTsnTTwoVA26RdjoOqEcJZf+4N
8euRFya0J2eU3dnTU3P3NOfVV5UmH3+AvSXUqX3bm0xcqLvLOypwDK9ivpUiAmK8
2cCrQiOEoGZHOACUeYTbSA==
`protect END_PROTECTED
