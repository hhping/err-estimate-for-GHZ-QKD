`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wh6UK7pVkXsWsGkowtcvZdOFeGh1FdiY43w1fS3Kv7icUQoEk+w902izZN87PvZt
YM0RPoXsmBX5UvsQfx1pl5rBu7+/6X24a0PhcpqBlktUdcaP2bcsb9SDWSIbx9Ru
1DmKEd0QSJPUmf+f2UH/Ayzg07oud1oE5bAFUJPdzng4IxjbMZx/gm+S9Z3F6Q6B
4wbclWxdO9TS3NhUGyqbIkzg8r4fPVwwKqCY57M7IZsEz+Vv/jaNnSPD23TROHbE
k2v7k5hlYJr7eUpu02C5AdSnKRA2ugiB1r48JO9ksGY1X6rbSiCJCoFQDt3AhJCL
txKu1YQc705hiZczLZjCbvVos2DpOebSPeLZq8ZYiWwxgRNSktpS62k6WjT4o7Vn
cN6sde3VBtA2dUfL79N3a64nnLVBiUg04bc8Yhcr/qsy3d+r60qkCFIuYSfaq0/y
eMUkIHiEn9nUzSVlsoSX6jZKNssSL5QIIQ+1Xs9PSbL9a5Yq45kjaCef1KnrQdE7
StllnQzNlmdWJJERoEz/hiCJYtnP1mJ2LY2ttzt/f3WNb2JfCY7zz7gFB3jO3euA
iMxSozwFFLS+5fsUVwx1Xb2tusLSYaUloJBUeO7Su6dTBhQ5QNO9aSe3vBCvFz+6
eD8lN+u2zPO541Xz0oJvuHGWLx1ImpjTdUrL0TAJlPR9XO44Iv5jEOz4lbjeJThf
waZ/RpCACtvpn4LXWTV4fWorxO5fFdN9AA0n6DyjScfiHkgntXxrtjT4WFJYT+ht
PLNbVExJMRsucQs9LeaoDe25EsU2ykCNgYHLSZg3J95AjmRiJ5ddjHCv52EzrjOs
Nw+WoH17REgSR4jQP3hA+oLtUr6vOfUD2AweYCnnruhsczyiWIvI1PbsQws3ClRD
3/ThvyTBiLwfe/8vLtx06mqPpAq9fv45VocL7e4pLy7JLOTFDiQKkl3LAYPQCx1P
Z8MHWeg+zc5Kz3gONOwgvC/6MfuFaZ7W2BWNfUNlv/f/Xb//U4B4lcgn9XL63bYl
gJI+qEGffMz4s2Bm6TLF0Q==
`protect END_PROTECTED
