`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8huSElbDhWuvsuQGmRFt88ZOBIfNjDkYmZX/t4wDLJ0OoC1FEtP1yNaq/CvdfEzA
KZRgkqIWekS6V4YklvsgUl7gDe8PXJNOnRegDViwht4xyVEv1UAztkOibWR4za2Q
is1G+1/kIBA10xMbk/8Smz4Z4obGg+MVLpRJ9eLqpY8nGjIeUA5L4Z3ql0wyzMoj
/96Bw3qBvjQ+u+UNQvcwJi4k0R+vTj3Oscox7RjwG88wOPOfSML9l+82rB0RNddR
KH8Yw0NVkz9I3IV8hIfUE3JA9hrQ34EwP0Nei5/7tAEGoGZ2xpGCylluCeffEbrF
m+xCauBOC9bVi1UPwlxzBUF3WwWMLxjlQM9HMAgvHKmSd0Mpaa0jZTKKtAL0rggj
PKsPgsnmq5GSOvEjJ/RmofzjrG5sHfxxWR3PluVMTe6A5scK07xM23+cCgquOT7q
f12d68PjLBBTaWvKufzbd5YElEeIvhaYt5Q9lhTOGB7JVp8PlNaLoQ3KyZAzERLC
UpE2V87HoNbwODXuyZOMnUqRnoSneiZcfAhqQKKWr69NnemZ6cnMo/9Kosf7M56n
gqKXRg857NnfsDkWrxDbj+SrvrIvKFv8LhCJWBhXEog0AcNKC3KSlYpMniwqM2DQ
yioqwzwzD+txtP7bz7ETiOdgSgbcu3b88iqdpEr5M2fm/yknJukRuJQ3CbRBRn0k
UtL80OckzDdFS1Z4VwbrAUXx08+itMZm2iePp5RsBVDntKs61d4/drq01jBW50uA
u8OoLPNHkEJGsm0Oc8WClzlQ3rzoZIiv7LEdmXEh+Gm3HEbicmwIM+jMwAlYrXeP
tmT7nYK6RTRptx5hxnk/5jPXpYwoN6LiccKxoBTF+GXkhlfwYj5KjoR3YpYsDbeQ
Kn5GUsNVUYx6o4oNdXMETzPfDFAJm6miY0WRGLiXNTu12L7bhf4BzDS5KrJqu5MR
`protect END_PROTECTED
