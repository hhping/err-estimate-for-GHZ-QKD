`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTCB2jP3Qi8VKX9rRK1RH73SNVU6eM+SjH6jsi28EkcGVgKfYpbjCwWHfSYmg/wX
OfA8hs0ci7duky03Y6B/MAdKbcRAuYzkOGyYKYzbwG93VL93aWYqk/WRROMivnfz
uvBUobfolyRd3fHDh71VH2Jz5j1NW0Wf4gdRQRP93lqs4TtyG99OUi7TkHQ0zWPo
35swI9G3toPGc+He//sO0II2jPfPCv8IXAa3PpwLJN8TQ7oV6mJY2cv9efenv+zp
w4m8kJ3kge9Pfz0TLZogr/a9R25LdgMesyvxQ8oaPn92eMLP2TmPmXri0OWkneE7
ahMjXN3wlLSWMlmS46O1T3o/7mRiupKxwyCI3kAurshOlBqaIetHsUiO1T2FOP5k
rpGcylSueFcPE9x24t1aZUmhymHHaeVKohfoyt8NR0w0DEAoDFvUcQJR4UB72qvb
9x67TzOv3SowtIZ5KPkaHrxG1nZQzoG9887ELq4CFXzw88fdU0Tzh3LiuG+LV7Uh
2FSyGTf4+/4xwtZcVbAIARmmLNyZcifiKe4rXiRVc2rtvyZUhdNuqTbbFxk0MmER
xSrGJ/L6A6WOg9mAtGNG339Z8zckvNKyd16ZHn7ZN6zotjBntup5q4gWWrMa1DVz
6t9c789fBSM4B0le3udbtY15cnkOphrCbR/lVlXPHzghS091Iuf43qzSCWwlf21a
Nlua8bCsCp4g4JuW+MXbAd+tGVACMW/U2vTFeHtoQNa/OxLqVK7nRzIb9LM0v5SM
GmqgEbmwAnP2hIw4hu/Q5g==
`protect END_PROTECTED
