`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2LR5z57b+/xxDNGKfUyUP1663abpokjtc7aDYaiN/GL4FRhPeP6ljrdiVb9B0fN
xmzHWaOZVmrKFnl0D2/6EtfB0jQS2wjzQQ2HphqGsVxGbyI+7aPEn2BaSnAwxqgj
Yrv+O1nA4lw8vlwCmfN7jjzsXzNlNYJ0tn259x9OJRxisXXNjcQadyNtRBvAWA3p
0a9BJw5gVTRXKPnRHMMVqFq8R0ruZxXBpcX+rCqttFEjpLRXWDlGDydc7bls/33v
2nQTn6WFGwzzXFJ49cv04mdqKBQ9DorJK/nvvsGM9yF/2OHhJeli+mD+zMp0XsD8
gEOjEu8jLcRh83mYgZu7UgfJtHmdRDwwOc3JlIhLoiqM8Uc67BKxk49nIyp6uNwO
ScYdofaZKdNDUq+GNXjlMICmC2tBKLK+8MBYY6JUxsKi+X4SyQC0e22qXi124Ewo
0eYb/6/b3eDl324X7DczuOuCEL/vkIYMWraw0Tb3M/ErqkNl0iyUUrzGNG4P7Q4Y
g5Gn0qDBAjhrzwx8NA4BaMpIbAFMfg0U2zhMTsQBFPrGdaZwwX8Wg+L7VkuG4SIb
bH8kYp6i50S5eUbkhdFhVllJ36uBG0KeV7aW/etQQZlqmI2Y0wVuYMLpJvD3/5QQ
H+0/5H3nSFzt1x3tworobwDEHcK+hFo5s+WtrR5PapwHMoz34gzTXLc6cRxoDuQ8
oIFeI7DGA465mxqj5HBoWrGreX9JzL3qR56qdnbnUMZqmzvzeBdY4KQF4khtz7wm
+usDO3ANSQciD5+D8TXbwzDgbYp6FHF+3INvdiGof/oQQXpGgZOYJ9fkIA65BCYj
GAKY0gptXnJ5ztTvWaXbCRUkKN2TDkhoOhfnAZ8KT862kHGWHNYbP4UjBqtNz/G1
6nzUd5uJDYPvBY2PTim7Ak/WdAXSKcsKYM6V3MgXGweroBkltIjSaA8A4vy4wEMg
U6Zp1v5l94PXUfs5FDUi4xL45tH2nDfjlwAev7s9/oXK47TASB0xCl0UwthBHuEw
YEvDLX6KMoGOfcc5ncWI/nEbS7xL28iMaVZZ9oCcxZ7U9WcOQjw6M8wWBReKan8F
V1Wj21+KbYp1/yGohJAW0qRjVwktX4hk9cH+LPJsUpaFheQWqSwge7CR4xupqjoV
DSJ0PVfSVtw+3/OUM4U3sg+ipTz34MILI9yEYfzYVFl0p6Sysp3WnWHHghJDQJ+x
uTzFzlYoVn/VYhKsaEWIk/j1XGmwzHQ+v/vRnSzH45hpbXgzO8g5zVvthHaDXJ4F
wMQR1EFZcH5SjpJII6c+y3Ok7pZgtcfwoHALcXkUP/CmM2KNhKJxIafhG+4EZyB0
ZddWjAPfzSqbCCPK/7yEmQ==
`protect END_PROTECTED
