`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SORTEBa8Yni8axC5UqIo1fZf5MGAF0SYe89cYaZwgNIGgYaECfXQYGKsyxV0Wd8u
lW6YJqM2hjiu0vw+9hBMcBaJnCCp4Biktj61yahvlaJLNTNdR7F3sjkGjvFlze/a
FVANvUg5WWDSbn5PdoNeYn99jMBWD5c9SEC9eTrti1i+UECN3Z/9bGY+7PG86hoO
JlrgmE92jbIHcDWJB08t1nNNWwGrVOvJYahVeeBtSV8wc34ZSVtH4+/aJ2N0znnc
2r4bGaTAqPFh0HJzMXJUUEwcyCzWR+TwfsC2NAqMtZfacz94KerTAXtcX7nUAROM
zCiGADfeVu9ZM3K30t9Y5B+JYnd6vsZ4iAR5skqObe6FbTWcASYPOGNopAQQIIfx
fp8bFzT9jAOukM66BPBO8Nm0TK+DcLHn/8zLV4XetuHndl0c/yYwg93Tx7PrlzZQ
6REwBfjuptRbJVvCpbM01td6HVMAT/CcLxv26pz33n9IoE4L5U4fuQTyNcnJMqol
FHvLNCfilWEpcpcy21ZPC8xs9AYNC5gVK8wylCV1tIw2imZk9qwbL4OYPWUv3Qho
cX+Oz6rjMnC8vNcQeZJsebGnN8ppwiIzAR6zfEFaCVm1WTxhRygUMAuOlRasDrKL
vC3BG+pCRPlrlS39Hbr5Ig==
`protect END_PROTECTED
