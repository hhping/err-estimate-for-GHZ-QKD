`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5M3UNlwfMSKz7hZVjYiy9y8Rzx28Ooa2vlZYhO/HceVhUwqjZLXiCYqOQMzSmVE
2D9S03FIjPi5u6KkaYNmvIZJ3vq1yegnvb2jof8lpFJ8s04chzFdBLGUWCaA1w3j
jdo5YjBBN0TtQba73y3FKSlHMTBjm9FVUmcIhpfEL6iVHv9KpEEgnJ4ObyFnk/gu
3mHPqfRB+EgsWtfMCbRtz1ZNH9qDt7pwB3NPA1VAHruLjlhAhALOaDIvHbbOpklQ
6PRW1X8opB2DxSrsU11l8xaknfwzfdcm0uG0JQaqDiFwGeEzwLOYTL2QgA4Yv5+K
jLqLT49M+5L789AtYCYP+w5ryisy9E5IEfkQKgJq2HVPWICpl9tFXIFZniGLyYRI
oLjqSzW/S7o7BBOhykNqBSO1mH4kV4Yb+ze1qBB4jvaXACA+FpcgeJ/qMW6FQ9Ts
xQ5HxisXGyFy+w6gLcrDgfQUZsT4LE2OayJkYHhgpYnBH5azwB4XMH7qeFnPwzHT
yzmCdGBGP+uKirGdhjYAMdRCJo9t5j3+nogA7J7+1nbXzW/xj0Swx7xh93ltz067
H5DnJY1XP5CbDV5g/t/gy1/RRXy3te8Txdq7YcJhMADe94ZprKNuEocGP1A9/S6E
xIt00dYBf5o0c7y6tzvOQf6P8M06p49egwK2hY3mtTBrqJX+CUXDcYbKn3+lJ5d9
wbhRwNNNmC0vyh62rBaXrDCDVvUlgoLvLY4Mkg+XSzmORop830AzNBj3ADFY9qUc
dTeNd56YTigiqyHzWLk0MBn4WqjOeIjcPRhdNhhWpRIP++CmbZxKmXbiLpCwISpW
n2weGC8WdZCYHF64P5PzQTktzMuWKD99Lq37aIDioM7GxQ7/AumycEhq5IDBkMvw
wrJXCzv6PuCjr0jC5MGWahwAmVVp2j23EdVXhKAy4C/21kdbwvh6AjSQNuCrVbMO
E9btb3TUyvW352vgfgV41TkZ6eqs7MzrXhtRRJqJH6qvrKKE6tlu3ZlSLXkv97Pe
9BsVzTdhRFt4lOTeJUAnIIAZaYQ33TNsOOYxEwiwnjpZyl7Nxmx164OhcjyKFa7h
IRMQWHMg5juiRlifiSyNTfi2YkwPWK4PRSit0+EF2cfOSms6A3eBof9i+zV3QYYR
kVEjXRjXMBK/vpTOhq+7WqOF8meckHPGjeM/9DpVKVY9sz/L/O915FK89IAsgsQJ
zhDIAvEzKffknG/rmyH49y+T5SWIg6ZWEm67ELU8plU=
`protect END_PROTECTED
