`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9JUUmXrX6VPOAWxom09R7JsyFZgSsw83gpPezRLEd6VIhOUYc5JQMJeXnUfxruP
wThGF3/Y41tPUHZXP9fgb3YByd/IGwqbsBlXIdKN4lzQ59PRtidl5SbNABcRZI6f
0oyXwBAZsqgf4aQJUrtOKP+oq99oW5RcHQ6JvGRxVIIzvnoBx36lBW8L8hzLKWha
Xjxvn/i4FOKWx3CIQT2dwM+V3RfcngJJzQTXzHm+ze6AOVxx2nJsbyZfaYD6gW5/
OIoXS2W8f9RrB/nGUKvi0V6D/r4e1+YRisu40ZHejzBwzFz3JpAyPVy3vLV+JPi8
fVl3c3Rcy85ea17DbdKFPteDdCLyKXA87OKfOgVMih8=
`protect END_PROTECTED
