`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
okks6qj/q94oDiHuLNQmN+YV35RebgPkxcAwtQs3qPlivv8/IdLdR5ZmgOMqlP5w
Jbk+IDwwXUf6ybyMrwtNhqPUV35wpCLrxFs86c5cR7Lougy+No+t0eTfrqvZtmcz
fYT3yRfxyQXvRxv9BEEfrYp/3QK0yQqTFDRKGH5SxU8YBM+CAClnu1rF3zEs203A
CKPRfHJpDos95g3wS5VDq1VzOCKNUDJu4N7m8g+AXxx16tB/fcTsNXlqUUWVP5tV
MmJxT7BYL7Gd5tkobcmp7d5kIrZyI8xHRgtKihxg90yBF1iMWXuO+D+f5KuONyN7
+03is+O3vWKuv7QNT6LpKm78nZHRAh/Zz1p+659tWywMxHWyOOy/wvkQ/OG21bKX
0e6PFjpBH87wW7GHI3J3wYNyi67A6gbCsQHkf3eisJR1G4cPCB4NMPSZCsHvBc+9
xDNDW89G3hhchjAGeouAFMinBAF+FY0RK8fTFsMca4O6baP+zuvSY+byF1e7HqGN
AjeMkRYWPq2UM43mTKvdAxrBrTmyDbw0X1Au5Sx1YYz6GSSn72TKTEA5HSJynPWf
96ioUpyKHAzdpX0KIMSTx/KfImmWonoiq11PJpLv49FROd8GopJ0AqmSMQr21AYm
8QqjTwFmxoiA8t+sVYQEyHoEPKYng35gx6sM1wka7kW06VSnjxX97VM9+N2AI+A9
tfJW3XbgrdbP5myM1mOLoXwJhxl54OVptKjuG+/XNwXMKcRMZZaV/ux/OOVINrHQ
6XzDreHR9mBoLmnsr6vP8fLEdKF4o0rjO12pleLPlNPuh4bu1/fbtCH3sSrNv2VO
I2UpdwAKGAGYpY07gsUtX21gAEOLHI5IxgsFOCFVOAp0ohf3kl+OUL79hmOM60EL
jqMz9Tva5IpdHOWeB74PfLULfa3W4ulCsekQGvpT/iRhXnS/teS3pCP7xsg09kDM
8LT4BXVQKJcpYzkWBOzBb+TjEKSGEG9YTQRi6riymg9LqlUDHHqjjQ3isIgdnJco
uNa55oLgBePLUojDACpqjM52ipO7Veob6HuRxm6SDEZCroEMIRX0bPPplExTx4bl
5pMU1xMiP60Nub2qBy9Vtuc2kvlQpFHzwBvuj3S5W/H2QUtqiBZ6UL167BqRZ/9/
fzEIhHMJuWrONvLkp4Apdfx05dkNBVXb4CIkVMzq+2I=
`protect END_PROTECTED
