`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4t5Vsm1aiiOyZrb2YlHOuhVI9p6V35n6caPrXL/QTtkyMolaplW34oFKTd6188d
i1MlJ+PjYbVC508fKWyjAKPdQ8KBkHqXCbL6ykBrONHZI0PFQMGDnbJujmTI79Qk
zMcXgK0hxl9RX+DiIhxuyn3k2930Vdz6mtBFSPM5UF0GkxiTZDhxhnhhXDfO23rJ
eOnKj6zXgIVhA/oxVdlQ8UbcCBTL4HoHM+X5/oYV8XnMCEWMr1bui9MBthdjG/YU
KAuG4ZtCAqmcu4HgkVSFIJX8epRFQmk9T2GSJQZ3E3GMta/0c4+zU1kaR76CVSk5
al+5VqHeDaz80OmuKA+GSJh/yWMSh2hxgdfJU3agroI6FRBUEGW6UWl9AkpfDTLK
OVmkP8h4t/HLrl7LgcUPnargQERqJXhPQXsSqgqnfF4IGK+fSpyuzKkI1EXtRnA8
xFAwKVzoBFyqzlP+RTKlKhiF33/Q8Vjq9MZLNaQFEDzTK97IXo/YDvioKCihVdRz
8CUPsWFky5L17Y2dVURm4S+ALWGO3I2JUwMmhnvPUavXddTp6gm/rGH8rAJi9zei
3tS9be0syfubNuGp9i4JeQwx3HNujKcmGlp36HbBkiD2/cnjO4q0SVRJaMPkuaBe
CZuatx/S/GLlzuHP6I+Ll/3kwzjp1/5dkGgkYRfI1AJBSE+CIdAtZ2zwqgdXZRJU
dJY0Zd+o+nH9dID2o7SYK3WL9p++Jx4oaP7CktE9D1kf7W3OG1QjjMAeQBGFZshb
2DQZVwvieIIm5QFxGU0DGYkRn3FnpiJFdJufLJ6101g=
`protect END_PROTECTED
