`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYiQpLsc3pULlx4cqQMAG9b/ugnPUh/N0WiAc3PStCXHWV80MhSwz4wrd8bcYPQm
BhQpWv3bE+1E6jenTxrCRjhQcvXBgHR6xUntFzsknQTRt4cAKBAa6vH/ha7kcbh9
eOxWsgvlmltUTKmFkOuQppA2aAnia+JxITrBkoYONAiAW6f2OwvylyFaIZVLiS8D
y96S3aJAInCZFz6g84QXMHN6s/bfSeBDNFUmc70PxjQyDOq/lyKCWG9GMPhqQAYw
CZWUCHYNMBrhRFFQ9qJvD+9b8U5cASMF7KHMV/NiNzTUBwzw3oYeXMmLEp7w5V8r
/Med08DeD8BlfF1Jvd17pGPc2RjuDYW26NzwWGtlH6IXyAWJMxOJM8q1sWEh4pP0
2sPNJBFmXCgd252I+zh6WeeuR3F9IGSY+7JxSItbhyY=
`protect END_PROTECTED
