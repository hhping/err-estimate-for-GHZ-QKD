`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ohqVigdhHwylAGu0kyQCfLzODdVLXxzBUbzU+OGdHvK0UCGtjbcNfJ2uzC5gfZA
S41Ir5ZCij41tX/261ek9ERGa+CADUW6+qC+S+Y0XG0X26g2mGllNEardjGrpr+h
2tmI3AghtIxOMPRBPx/SvRyeToEbxPdkgYFvjI6i5NlzWfNNPmRgdDC2hcLLvlVf
MTewu0x6qhahvqVo1jj3QzrbnOQJiFvBIN9L1fgLbFPUeVA9ecWYVhMsl3vdV2Fr
kjxrunfstwHouRBRGUGvZHOuG1sFuUpku7ecaw1iNsid4iU7tZsBbrmDEIWLxrj+
oMRXZQsS+gLqtkk5vj3ChHEX9kF+/kMKviHK2qIq+YqU7uGbuqMUEXx69ULtKNiQ
d0e/cK6N5IeilBUT2BxFLY0p8n66qkM3Zi/WgIgrJm7a8y3mLAGFSLyYVp6+8Baj
/4hOGJ/AMtgzkY3AMABuJkx0xcxk42W78rMnAIqaVRE=
`protect END_PROTECTED
