`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2N4a+wHInAM7bku1Q912BpYFtpfRgGMHSHF7e2D7BzDTICpZ6g6ic/+IzzVGvgf/
nZjv04TS6Hd92C3zjUWpp1Ce3E9jTiafJvKaDwNI36RsR4zLriabgmOY5ycmt0m9
A+3NWkhEUulmLWLoG93Rxm35q92ChQGDVMysVs5SJzo/6uKfQE3sx6auTMC/+TII
saj9on1UjtvcG0efycJKg4BBiaacjKzdE5JEYtAXr1p95YU+HkSI7w5uDxicpzfd
t+jd27TrUlMH1YtJI6zCQ1ZygGmyukQcImNwRYtE/gKc0hGt3mwe2QaeRc67QGQ/
PuGJmwUZBQvdMtvgq4yGpHVrAUDClhZGfKT61V9tbRYt4i5BwcIv4+06okamRDOV
A0Ws9S8OPtiiLnJsV80fhash/JvkSA4UgL3/nSKstysHs9cFGhMX+mcBBzQzA3O5
JRIJBVbOvhPBrcSjpx9CiMf8KUFvGV8um8Kg35P02yaNbB9LK1fpn2xpjtAkIEKC
BR4qpiRRfG6RHAHhPvqnjz3/nzdyG16P9Km2nDbyaC8UiUVBeboHRJjoNmQlEF1j
QTHXrghmE1NCC8o8cPz3Rw==
`protect END_PROTECTED
