`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUGS3fotEVfDYCeH24fFUUh1hTtqRgf+Q7YKdY33IqICeuuhfoqMeucLUCH3nSL9
BZGhPPjpYp4oxAMqhFG/WP34VIKK9PLGd4yMVDScoAINe2/XZn5RZoEQ61vRkFK+
4kr7FyT8RNf16RGUUKXRs0mr7VMchAtmGFWjhhXAclNaAi97VfV50I/nZ/KrGzHJ
QmTEyl8Mqidt+jjAKSBUrkfblVx4+l48qdowrSxGSlfi/vvbZv05IlWoOCr6G4kk
ZGmGkSGPnJJKG0vrPPvO44aW1tr7oif+nZ0p97LuLlWSFCPr7k+C5dW8zlQjav2M
5CRggKoWZOhi965vA4QQsT3vvGglwaNMM9GXgxiZb2CoeK7nxHykN0q95lqhLR/m
mLFbhTOU5eSZbSQ9TMoEBtKaINuO9ELSq33ih/wp9J9eENr6+CiCQ79FUyovfuQX
hUaeGxhmWz3j9u00hghg22mqqib2ldogU6ou2TyGhbf7170nB/ptgk8yDAmPaAlD
R9Pk23034qtb+CvxUxtJpSWU3kgnbBJRaEp2a4NXTTW26kBgTJhqXa+mQCDeYSDD
eznLUx1rXbaz0j2oQ9Gk2h+QXZcs/HXuEsRvrC1q9Gpk96uCrS0P6j5NDrrAWtu+
u5+b88jV7i+o0u/ldV3Lf9cDiAYYt9yh5N7u+l6JnNKr+TbVcv0bMseGa4zksfVu
HgDyIkLNWO/keK2ZFje4rX9L/i0OFTmTmyOUVZogqkVLGRq1/u99qMUpNf6NGNbU
749NAOchEMzKgvQaU4pjwaThMXwS/mlC9Dgd3qQwCFYb0YvTihHxyaFDivOF2sc/
KXDs6yObyIX+9NJwfHlFAgTnGCx8qHbtnL3xxSxdhydPcdxgl613eNAFgWrF5hNO
DjnmT3R3A3bpLyjcJ+3B9Eh0C9qzb51WalBais5KcfjCmRdgGEZ/ODcrXIaM9ur1
Lid1YtpIt3SJztmKQXl7ors5IqBrO/fdwjvbF07YsZDLNfZ/PNwlRkZ87L4O4Rbb
XeIqIBcH17k2RFPiozLfL7ADADQpK0ctRLuYoB/5lKbkJwo+J/0LyskrcrCwTmKN
NnSAPN0oClBpf2nFFJRcQQY0bg4ncj2WFbGpVirzz9hyjwmlIQXshchrI9XIxa6y
/LQsiZZMJM3Z2i/QSdZeewcN3DQg59G4NSqJlDsgtPuUgKwVPNs9M3ePaiIYJCMG
OU0eAZwTkF3T3H/980OKEw==
`protect END_PROTECTED
