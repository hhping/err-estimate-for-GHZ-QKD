`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5JRVNUmhFpLlNPbLXpPcnz/d/Q/fPwAbgqlc+llMJNhOiAsU8Uzm9qmHBpMRmNY
lArs0AJElllo9G6THPaqjQ4SSyDhJcq0fIZP4CyX5YIOH2431qP1MBkUxwBxLVtK
E5zgXnKLkl1E1wy6dlCs7XMqPvlhcBN0XfeiSHNRet8w4nCIB2IqS9qNRt645nZI
wyNyCNc57QIKvCxa37v51q7tCZWNolOOnNyzUKsoe8SLiHKfa/42sqed7tg+vb78
7x5HzgDU/ai/e09Q718i3MUboARyg2QVbxfmrlyHOXUZqpVQSTzOmIlKassbcKxW
4R5hyw9lOZsmx5j5ymERafy3Ou3pSuyW4XYyO3eHGCJVIfPHWqNrYeH1s/3B45tq
9H9zqdx86/9nClyYgVlk6Lhfp2i9PzIUWzhfN8UYXFv28qY9RTtZWZb+PmUvYA6R
35z55YcgdU+8QTS8jxic2qM/9glHK+s40PSzpWbin9x6lD8mLPcRGR9HGbK+l5hS
0lqkX1/U5VZRZBkW11GZjh5qw7MqDaVH9iXTY0G0nDYGlg2JYBpNrYE0hWbFAkcM
LOs+dqaxiSu7j7HBP8H7kR06vDZ30X3QRGNWjE3nFWw=
`protect END_PROTECTED
