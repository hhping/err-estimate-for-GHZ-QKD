`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/lkZrYnpK5No8bkJsnqOslqQ/yU5ccgXBHBAdtNu7KBkyLY2fcsPj2LpYG/0JWTT
C9ZYzeeTkxSo6hArp6vJP5o0ankYyRVNUFEbm1wcjj7yfU6NFNa4MNlJSScvZ4B7
LY4wLjRw4qMJvV7Ht9rje2lhKRnnDqMLxmPV+G6NtDHq4zd0wB+Duiz4m1RLC49o
12NDPgoq4wi3cwBKJmp6vxoerp3Khsl7kw7YMKTssatdjvAiDDoy/XyovQADCtqF
xWNu09MdfZfSgt2KbMTRKQHigmfmrfS++QEJtc3ezU/URq13VYmkb8vn54BDTRel
NGnWzojivqk1g8neaZaq1X3Us0IrIMdh5LAUvgyXYR7PW15132hy2E4H974gk04R
SVbGP4+CMT7qVr01N+556s2mcih/drCbEsTeL2LoSYFPYV8XAf2F5gVL6QXuqxEh
D3Cn3HQG/KI9E0xjZS1uAbooJvB0BvGUkgWhSIln6/GLjyOwWTTlWQc7e1c839BL
MPrw+kWRLYP/gUkS1nbKVtwhGhjuP50E7Yp9DJ4r7nRKw0AuFhr6N1MSs+eMdHeJ
+fpdnwq7I/Fb2a24nCdh8vZ5aGy+cOXyT3CvqURUwfKedYf+e7jCggom+AnunFoJ
YYQiwTENVtU3F1xYDR5kG9qDXHjexESqu7G35l+SQ/DjzzyGFABoOqPablD2wleH
icOo/WtSWi8WIDWqXt3++kwGQW3UyshPfFhicYTBX9t1fNr0E0bOuHC0x0WCHqh9
ADGL/K5SV1kZ9XHOjv3Y6OWMqa6uE38lWWlZCu8oLjW0aGoy/W46nRZpNa8TM0QM
Wy1d2rruF2FLuyZ3Ic1uZz03f4PPHFZMEG+1rPDyoAOfuDZrWZXQ70QGaEMuNlBF
22hsRrcbkGbuA4ck77RHgS5gavq9kGbJtiAH1eHRxVeZJXYRo5MrtizrVUY7kYb9
uTIR3uRjvnTKVBXkFloBOAcEqYn8uO7uLVSQ+4QhoVl0LkNgRh3JJjk/DmtOJ+pz
dEHtJQyMRS3AgjshpmbLP6b4bXJWELhdo4o+IlNaEWjoLBBMaSoxe6UeE/AeWk2o
Ne9Sw0+7/lttVjmxhWqMhIsitrvCH456HzV4//RwecxnJBFpRs4rcS6UAHiUEgHZ
7Vle7CbXjfEzM5QcNIpMa6yxwPIH+oLocHoHHe/vOI2pX1jz+m+YrIGj9/RY+DGc
/aLnXcyCCOAnXvR5wZhOXLHviVazhaZ8OaAGBUDIseWcegODF1NCj7SUk7rEBwyk
dBLYqiDv1yar8aWJEdm3d5VKEn6QGs9qjnveWKrX0/erD04fVz0B5RuCs/wLUBVW
l0FIsVZUxsG3EAqc2NY584U4mi/QUSQFsHWJHFwJ8xkFtgdK8wCwu0KMiN4QBoAP
T9srbtISnTw/AY73Q7ChU3G1D4RT/kctnYGFopExulRW8HbaBOkt9jG6rfGmMwBH
uT5MXgT3oj2hdUXN7IDJQLR+N9JTYm1NZVMgL4oK/xt6tHf9nKXmLjr6KgFMZJcN
G71S0TguB2Vz5QJBvsctYG0xadRC39hZEVBjVzIfHEevKexBrsPylyrxDyePPgpX
4coYyHBjjCfm4r7wnGKs55E+na+JEf5zIcxadFrzpdpmHkPgCzD4tCSeAAzbaYyO
gwVW+2S1keQidAOhsioGPJtQEM82T6zHgC0eBUtAx58MmDeNCM94+mjr7V9yyNMd
Rp7TTFfFAgBmLQy6hMD222QZEkinrcQmjCs2XgkD7tb04mWPiXzEIiX1OLrnOB8M
o8Ly8F0pUrUmYE93MApV7rmGpzbTcJcKI5WtMG5RYtFrKaD9KtGHLnzproOG2eig
YdeVrWBh2LTF7KLlelpxfT8WDiF/aXCP2NqLh4tmnju5NuC5WtNjjWLVQJGBXd79
E/PqmulPKqB8fHsIjBAOFdwSDRPktyRHEtD3O+H1Y4bYD/4FDc+hDQG5VwSYZjB8
G/XBaWTFyFEmjjYPd1GbI915aD1EJb3DAFwoau/R+d3B24YUnHjw2/9Fb2/q6pU+
EkhmXFaRsJMXK/ZUm5LsTepU/WTNB6cSoTThcZenpq8trmU4tRzUPNT6PcxnhGe/
qn2qoDk3sa329cS4nClb7qLepVf7EKAxPuymvytpKepAZsRP3/djKzhV+gQZEknC
uHtpHE4tBxM6PE2HuyAM0ZeB9E/aKXed1I1CJqPL5d3Xf6ve8rOw76FPAgYgkX2x
Kk8UeOxgkZyl4h87IX5Cg7fcz9iFqmyMBd/ZK43Ek67e5B6REpP/sjYXEhqz2Ap2
/qc6DljLEFyYllrCs0Og+gsNd4Ak7+9ROfXDzdHFiSuOgq+aJYu+QktIEiwlfrzy
v2sFvhIH40F/1fJRWP0zDlhfpYwZPs1vFwBvwsdYnToxR1sMBNsdqPVIWz0OC1mY
oZ6gQX+oXeadg1q0BojHdPm9aBgh0LZgI6tjMNHheDcEXwbgelh7LCUrYqmzdtiZ
VyAKYlfrdzu7S18j0714r7LzwLoNJmeekelJAHRdJ5Yl9mRW5kkerSrnM0RFZf5x
CxTUblXrK+Kl6yHfvaFOHHRAl3IjQiVux+17wc3H4fJUVPzgqdElg15YDog7RZ1i
rSJ5rH19YVfXEyDrtAzkNfjh/0D7x2a9FdnS1dyXohqlkomcUU/rdVUwU8DiKYKw
fA1oD7BWz6/BJNTFlBsNzf7oncH8vPi4Puh9A4vwV9asmRpOlqZ3Sl9autBh3sA4
5kzf7AM3hm2AAGcWX9fRF2FNnTiBLSRwoT7CLTLtvNx4g6xpD0b2hx+MFPtqFAdA
u7DLPDr7jfEz26bvn37csZwVq9zDE191W3Y26lP3vlintiG7wHF7CB28znFpno1v
/lTBf/PTdnGC9UMoTDG99W9z+2FeLgAsKTwbaoSpDjGlmwYVdYVzVe64ffLjEU1B
f/8/iPFCssgVhp5EnQLXdOtPCmdQKJQNuWFvMxLRJEevomcM9cg84+enwOzcsYOC
`protect END_PROTECTED
