`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eiv/CdsXqclqNyR1gbL2bSttPtNQcRD/gRSu4xcfBYQ3p/jZX+s/BR8n1qwt5dN
Us2jgZeeLixJZejk39q6BlnfEUQCJkN8ax6fpj+c96wpa06b/HcFB9vHOvNb21i3
Plv6ROiNNuGuwF8Gkzb1Ds+nUuF4FMl7aLCruT6esP/MzTm7Od1/X9khsm7N+UCi
8QcEZFvB3lFfU6cndYsYYpIc5Z8L7pLvBW+/7IzZpHbHQVAzhIEtdxpDKng49gUC
14Q6/Xe9k4uB7hxf7z92eNzynTaG54IolURw+yUBNkSQ3KpnZJ9icQkJlKiOniHZ
O499HvBMgwm84KMspyok51Oy18v8LLHrqWVoKXXkCKVYjWrkRRzrgWRUsUoaMKh6
YT8Z5hj5/Sbqx8LyToXC+E0KThxOdt4lp1kH1KSV2rh0PbYp1tfA0xCFiIoy6IgH
nwDc8FxVIBZ8sblmNOo4qMhG3TYp7v6ydk55XH9l4IDqVIzzybOQa92AzFsBJrUZ
chzqn3y32AQfcSLi/m3etHzRMakCX31HiF9n9Yj+k1JVtdRm0i/KA4P7WQvyfeLt
des1K7LgKvy/3RLk67iMPgzMGFzYIqt/BXl+ACfAniBWwOxyffZ9PmJ0qJzntytP
9ndsRLUBP6FgioSxlwqe3GNf9Sr7xfOEzMjOyEi84Ki3s+iQQlUQxzCkXCaoFhuc
PqmFZkHZ6Mb3U0OG9GY3EqvaxId8nUFfPQGclBpuqxQltAL18hJlUQcDeZOGseA9
UgWi6GnU2IxmRWam9M8EaKQ1Eu7CPRvouYgJVcect7VAFpuRKutoKxYhtxxjkpN4
4tFDydR7RltSjm8crY5UwXfPRhj4g5AMz1fSnnSZM63NO+3BPLGJivhPQ/h8d4HO
C1Q6GTTerIhlLmZcF2ycsOgvVyOcxLvmA8bi8LTJHxyEKKPYL88UxXpYi2z4WluF
2A2d4jW7qqxHspw+cHB6+T+o7JMvEwx7Pvd2zgf0EQGXzwKn+dhaeP/i0rQV2W4p
s0xTp85lIRml1cYaQz+ZTflYELA/+y17mU5MX0QNJxoEhopGpkGEZAyZ1UzvwKBV
w5ppbwKUCo/quoFGWhVMQTb9RLZ/QGs44jHHnDP74SieUdaGiUbwwDkqZerBlyj5
nVlNfKGLL7PMVlkOlR8GmiPCLg64Q2DFUYfpaqHDU9N8vvp13QKLDqMf1w0HBKsI
Cwok2daeGwErSVFaxKBdADmeCGa2fwHZcODQQ6ncqrUq7Wm1ELOFrHAqmoklYw6G
R6JrrxlAS8gJU7y3VGOC6sNs3ZYS1k+976uB3GcMlJ+Q0oMGHSz0m9jkV6u30pAB
NA0V3FiOlHUGlq/7ORqjCiWimSNMAyLhR6y1X5B448yDI1t+hIPzbFRF59IRiN1r
IBPqVkVrwzyvLE0fDOpsZ3xRDgq61ySLLVAV698fFZIa5rJdW7ybOPnaf+G5ATJZ
WqukVCQSqKgLJ/y8QJ2dG1L7GJim8Xl8EbRoqMbTD4PoiDhwYMb6jlsl2fLchvG8
iDmb49m37J/DEwijvWcIregIfXy6415flEvVMJL5s7ky5TnmOcYS9T1dyLUeyl0n
mPwp093IpVQQe5t3T/A+vzUHbZ38SZChWvRd0ZjxJTAMSyUTgP9/LCQGFI88bLQM
crnWHSwQmWamZRerrG1fUhVJ5DPLltMsa4QFYwr44hDYU0RDXQz+H9dtudMSGx7Y
hiRHHFtNK5zMCDdnFSxZpR5qV6mV7upFXGUr//AhMbo/p6Cdg0EDQd3GiI8LW8FS
efh6J+tTGS7G6K/fzEV4sZmbmzI3854a91nk+yJNYdO5+bSaI+muWt64SNQVBKhX
p+FG+nOsytNgmqf+B9XZsfUma+x4hSjdOnVYdhQC6o/Yj4lF1Jt46O2AFyQvoAN7
8BrGU57ypERyt9ZGaq5S/33rqoQAM+oK4nYaqD8hx4M=
`protect END_PROTECTED
