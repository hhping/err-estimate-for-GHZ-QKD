`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+wsPmhFolOZ1vIyhCVhAnwF/AuGu+uwJlQGNsKQ+DVM9i+m8hXGJ4bKbudr93s76
RajRb1mBkEyafCSPRmShJ9+lamm5asecG4os7mmBNG5ToEKCLOnhnFj1o1Pozdc1
psVxGm8VZi6ps30jCqbronwWe4gdkfH9tslZyp5B8C24UfblpPOSfESveIuWjXfz
aksqrr1k5IS0gxzjtI5K8MiAeRMVtkjYHI5TuXqXawN/puRXFdU7aZiOXy+gFywP
e5Xo0dh0iCci+wGM/lvksG4bHbEbNlW4a3yJ5YATEBTOXURmpnvFnzt1kHw8dxoU
3LvzmsnNMuJNHgRmcztPpuS0w75Km8f4k6lhxzpdtiFWDk/0Vq1fSKQJfLwCMzu0
kWiyQnnTAnNXyC0Qm7WdJVqYxVQU3oj4nhMdNMF5+gEQjL5ReodEIxhpFGNcEJ+U
28xJbPUeO7CaF7VflfI+GvVg28aoBPNeHGuFSDMkBBqgT2JLn5yYbtqcRtA5hfH/
NvhCbEn03w8Qujpz0AfUkD68eMe7UREGe34UswhaEo8pemg3hl0yXt5JZn+dsEWc
CMWs1Quunv6idfccB7pstQhz6zBbK73gZYZ43/ezouHiIdhtzjwNvTec6IcWBLcE
Veiepr2XkljqvyQtvAtM9I1PO38n5jtFBHHhEHmKreod4T6TJQKSYjvZF875enXw
4UY0q0KvudMW8cjqB6xLc6pgNYidCvU8cssY4qF4mVrPjPMZVaTn2qMaDRrQbSQU
phq/qDZsJErhtOJzCAotRenGdw1eK6RGWFejtSTYcVuFiVKKxqhumJT4EyPJrA7b
N8r6ltO2lQpGQ1Sen+x1ZeBtOV3Bj6UHkN59DWLZtps7ER5iQTNedWMW5+DatVSH
4qIKge0I3hJXkxlrV9vgyZ4EMGB3ZxzbPTtj0xojlFFAsh6kbCd1963QxPVPUoG3
ty6iry+hwr5nQpc22iNIb3oW9K9sR3MtGm4XHaxGt9VePloiE3mkLeLSbCXpnQb6
aJQV7zrJRAz3O/gKai2Y06tHrTrkWgBotbfk9hiagwjcDWeO8zDuv/UWhWfRqCaf
wR8kA42OCiXWcMCRXi9mmOTDgoSnOpT1JrQ4Hyv5cBqzygGOkaXxnXwv0nwRKAqs
XIiPRwQFNGo+EOZZyTK8IoKrF/J1af1PFlPnZEy0MYSyxOM38HjK1LCw/Jxbqlxn
kWvfSuEl94fFSePW7z5EpY7wsJAqguhKcEQeBjUKJ1mMHgmiM6YA6IItckXAl0yO
UDfb8Sp7sabRG+sWEv8QS9GfkcvuJFuyRI493DJVzeHrrxDNb5yDIzzLQmOZCSEe
K2LGB0xLiivYfR4rtHXIvvo8fq+bShJIcLuAwzBPAXBZYCTvI2Du2TdnRCWyRLmk
G4eZX4mt/v9VxKo50yIh+v9VlEsebK+vSYNWgppHvCid6oIvDkidvQZAc31PUXD2
OXnZkQOOBeaX2WTIZlAwNfwqpq9/B4KE2g/64pr7nbDFl3tOodC0mtla7r02cyqm
EOB5Ac0kTS6cIXC+450cRKaXIeNGnu7Ngg5gT5Ba+ZyYSUjYto3LpApYhDya3TLy
MI5VLr63+j9rnTcih4UGuoAq/VGHd0Q0TSk2n2zGmRalHlbYElu0KHQv6DIonBR7
VpcKu6tjJwv5r1LWp9bYF0cD8YKiHVEr2Hq341vioIh7aNKN+VKxuRQqo9FYWYjE
DPTdLgNsfkBOYPofd5t271AN67eKiBNpzQiTOVdVP52LZdAkId/FWMcUM/TofMq7
zgQxLvPBiYDQkGqUGZBEqmwVMest2N2xQ5/2AI3zSNSLJhK0wsdg7jYMvPwXbZua
DItGCjRfpiaAEInETm70ADidSZ7g80MyCmCmG+OWjVk6vHElnlt/kRnf3GPV1HuB
jCAiFCKckBpMbjr5zaHl3isnrALH7hzDUFN6DddFPhse9uKBxSmxXkraDEwtJEEG
8SrkNlKRY2yb6yk27rtrK9jSF+0n6WJ12PhzuEJEzslu460+PPuO0Zo8unGv19Pa
tNm4UEWzb+S3uF9UR9FUSBwKcPiqg45E858wbpNLlQMiER/ovh160kFbaz6kvT4I
MuQi7GcXolG7RTmTwtkIl8nS841jEazqc85vvoukQEw8X+hKmK+cyd1OdHtxyCWB
OwLBEfd1/oqNd8kFrIKkzfbSG9mCzo7gXm1OUT7XjR3fkns+66tzkZxRAwNYPQlf
R1iOYbT9JHjvYUmIsCcFWFuwVleRa5+8vqSfv7GBIrSMzJFESRjq8YD25eyOhTqm
kMU/S1nGlxpO5giym/1OYsfqT9m6hjRVMsq86ILhUDnwUk0ObvTRhy7l2wYqN7mp
LHcHI+uF+HhtcnFNj7eSn6giORokV0iutP6on2BHmrKreexTakpiR4PHGA6/tLpZ
dLm+1ZUMrJFYdVzDXcCycAbotXkEN9bfFp/ZS2b6tfg4bAnVQx0YkpU4BvvVvhtQ
meZoyCmuWAgCK1AVlV2OQIvQSz1kjYZxFB+m8M2zCI//LaWO9mSfTPW6Tzw8tbOG
2ri/DaMlAvWvtOGCBS7ILppebw7WmAfhsD4uoAeDxKfL/RW3nT5cHktSEEWCrZlU
k8u0EmNgvtZZ27l0XTStCFWbZLEaFvO65LpH3+mfsieSYBKzNCvnQavSzUnprWr/
UUoU/VwLkVtyc/GCyS8jDKa03QNLOKWmll2FHCAE0y2GNnXV1oDJQshBcBmFhVlI
oKh0Ao6a4GjRiBXHFrMEMfZ+eLQ7IvyB9j72BoDqqErXG+0ltdTsHKXlokpbaXIu
y6E+8Rmqf/lddnqEp5PgwOq40/cpB29rK6NNI8TusZ7RQ8/4TjMAz0OlEnplWVmv
RiOiIDzTwa//YFQeGqjSrJJ+0ngvLb1MlhZz/rpWlmneUOLicwUxmRaJg5nPbI+q
fvsYzhahLIl2CJdJ8JIG8X1CWaFQ25AcGutdR4F94x6+sIx5YTqOcPUjCbWfVTjT
i8FLG++MDwufuGw6nAWNymjOF39Byo+bnOzEkpANfzg0uMmkyXgpnmN4nhqYXpyt
Cb472KHpzwtaxN3cMe6jEgF3VNS+tI2QiQfWuxG8QPLsZOo96kEZXdrrN2D/HTzt
f7y4xhk+20tHyo6S6k7xvWgVl07vbfguQzyJPTgAMXJS5aXIZ4kKwwn2EEDnodts
5bzksyelS6eyqk1IJW2vcgiSUwd+reyUhsAVDfeFdxAtaFt8/kEodSxQeimPQyI6
KpGtJ6uLl3tIWMt+Tsyyg1yiLtn6npT5JFfJoma23FXdfhcIt09VgZeQc2jKjJRI
GEtC0th4cmlk914G1bV3zBPJ5t+dmL0N7FyByz0TssxiIYIsa1X/+t1nz1Ki/tW+
gRBH077FGeW/ENmEC/jXyZMZ08gmqg3KPMly3/Mz6rIZ0FkKNCe9MEGanmKEMuLR
jznM0+R58vBiokunlaFy7fKe/PbVp5fZqGfBBzB+rlqaHs5ny347/hMimmJXZaaa
kgZ72tTTkQOWCicFDAYU2U7lvZBVA81GfSFHaN6eCsSp/YJP7fEqTbnvxcC2x694
aosLm1PlJCOfyYBneVHwVmP1qNDdAJDZ6QiWguIK7SlSWZT+sQGmf9w9FEhRQAEk
yOjsFOooJ/BrUzAa3c3uqfMQwQlPh8Yxx68tv8K5fEIQ42HFJuHAgijmzNoZmVin
fHGe5RZ5JdpveB+YN6z/3u8MgWp0X7EzhG0zDWa2DHQFqsqc6/OjsRgkF2m9Eca3
VGieQyOFbAVE0cOpazrICEcgryZQ6lDrnqv96TxMEynVs/vjNfuiQmh3QZWg61Ff
JoecnITobxAOc0vspoTguEi22dO7q+uSIAQkiD8PRbO+XmyDCH3DmBxQ1YzGRKth
JsNTpnVPE7tNhgcTmOVYjCHhcKOFI+K3Y4/4cD3zq2n5T81MOD5vlS7jPBsy3l8n
z6kecoEjYGOdE3X8QwdRrCfcgt527TawizpdcMf1ugUiW6KfSr7fi9yRO8knECaJ
4ws8bfsXL201sDCB9hJGQzKGXGvnvL6MayeVO/pET7UeU/Dam6Bo42bsa8mgnnjm
Gx0/2d9xZUIpHPcfd1MBcFpNHV+6UIIXNU8zDBKxBMSvoSl0BYGYYznRD+DkZMED
y3iS8w28hREdQ7dOiuuO2sKcRlPl5KeDuo8OxEFG6N2as4JqOuysXyGJnULcQDyM
XKfNTz4YyHlV3Eo7fAsSG1dGIJNX4APlK9aEPODSxuPq0REfJXTYRJ+vd9IRDR/S
K0CbDxNQetIw0SX76gAFPVSZasLbHkhvxN+bg4+nhg1CiMw9lpOuwRrWP0B044S5
jL6jdlnFLLiVeZoqkX2ajY5bKy8YTRlXX6DRpXBuA0rivONcODx3o2YAvhBFMew4
JQCX92i+IQkjsdIcnDPnZB4UV3jjTRd7VhHVibZh6KW3wDZztR568AK25q6/Ww6q
5jL+LpV5s68C1GaWvfCNWP4poJNq9gTWIR1qWtqf+uTiMMf07ncRJq3rZYxdCOrs
XPGneg4D+mXKxPRZzMFJtSzFiJvuiSmdmmnWbqpfV22wjvE66wovndbWW8xJVTSn
Gz+leGufw1FrAoo0XhHlobNoPqbaHoFtrc/fCwr+kRC0jGP1SVd5DlHCgbBp3lyl
128sOy6+r8EVfXSDsvUDwtLMkBi+RiA0IpUZDRhVwk6IP+ut0VVvtHX6ZCw0rdBp
1NGXNfh7u+ID95G//miEpMjn9GR2zlf777RsQQWllAKKF0/JaQYrZz/z3tw4v2Qu
2OcnWazteI9N/f/uEEASo+ENFSX4cCrP9TD7k9rSa9EBOVD4t+UNbAyAQJ2M8DU7
UNYS0R5NVMRIOmP2MbXLZGGprHfgwgK8smKAYALqVz0TlZGXfnvKf7NmE0sGEy9Z
8zoBL6QVKgvH9G1rNvz8rZtFtTMINyDHZARXx1MOOZFbPYfGOvSQxABcjIXIYbr2
qNhPSFOuRVKiHN95o3uNrg/UHhtcLKYTyq4QcUfEOWclBVxNdIBA8Lp8MjD2jn9H
18dwshGg+34PtUhj+Nx6GU+j+IlDslL4HZe9LOC67xU//uIhDpGTf29uOdVxeiI+
gVjDQkC5LrO/fHX1ZKDOpwEKWSdwAGNh10601e5fEW6MsL+2ht1ZymmqRcirn6FI
Bsf1ns9ZIbJfjkKpvDxVIAJVA0SFD09nbb1MGSqaCTx/8BgZpe2+bm6mhlAumaGd
HW1dKKO8WT3lvoz5qpvtmXn0A+g192tId2ADqZVeL4sD5DBsMgoJvd5deSjgSOnh
PsvqvpsjbEcmi98+i5j46248xywdcv4P1aHHYJz5fBBm6PPbzOUpCkspwoyh5X3B
7qsVZOQM3j+LfxCUy0optz62YtsbMGzj6x8/HPsbS/RAkd6PWUwfiGqKoTlrvl1D
CToFTvEdigx2jjfm54LLzjNzmlSklnCyUG2OWQorvYzE0C8CjSVD2f3N2YmAKqkn
4E/RgXFZEdI8MimiqwoTtaCRWuX/9VpV5Jv07pYXuLw3T+1MFybkdwIkhZXNS0PI
OpOlPc7xlUCK21lx/DDJtRlTJCLfofQCpwz11lFzjn9TgpKxvwQwuh9967auR6kf
VChkDQyTjX0OQ4Nm9VGAr/1FWYcW3dPbeqiMgnfTpdgnRTjPInEnkYcNVYhIRCHH
el7+v4sd8CHYd8kr86cavwL2t+Ddau8QJa8Lt/Ycha2jLzYsxIZKcW4tug+O5WUD
hixy1J3YF0RHhkI70KD+7D7ZLizzhV/eGBbb0cySHc0XQ28vfPDI9e5iGSwYHTt1
lIiwWnHPy0fCj4SGs6NVetFGoWZYpkXJAC4wcI/RvhL/IphEuvYr4lS/V1ImIZHo
kq+x9AOIh57gdWphaK/XYVsNNY8Vyz9Su+zXaJg+GsNBxe7kbjZxz97PEDzRYx8C
dyX6ENV2y0L/1BUOUyPsYupDZ2TxNfP7kXdIt1R5k+r3ycMbw5qnJOp8wLDgN1oQ
XUctZqPSvY0Mz9mBejSn4bGOHnDRSS3s0URHdU8CiR/HZ60ZOF6jjwt8q9KbR2dT
6HkhSxz+19sgbjDuxu9ch9IqGtHwp/F1QDophdYjkLzjZnAzkWWwYCe0BtuP8Tyi
VD5vbSfADZSOSP1v62kdRdqe3qCWnu67Uq5fjrIzFKydkCErAd/sPdIyDizLOfaJ
PHTClp0b2GP0578GsUq0wo4GjNHd4lr3uSD1yh5y7HfmU4YRwdyWhJZ7XUPSK1Oe
6ktagKRq4+c2RICDA8epWHK4JOQWSpD0QNoS/eYCsE0b1enh/XAcBlMGUy4btY8s
jcKVtXnY+eIFA8ft5PnSdT4nkhvp6LHHW4R/5Al3UjCvVRKuBZuWyfvvuDnKmKkw
8wQ/j6pUf38ajYVHRaeVxJPMGi718yMwAfckbKPLI03DxEGD9ZeC09kGNc4R2KTR
cf32f3ZQq7tKkUxtiBKCakkECi/TtORWCqyNGgfgh40fA5dekUOgENY92BOVZgQw
juYOVeHPR7lcFFj0pyh/QEeWrPgBydg2YZCkAC2k2umMzrGZTTlTFKZAuKdlrnPw
Q9VDaGXcy5lcqa7ASdf2Uadm+AYt7vq6eVoSb3UTONF6aTFkSlBoSHs5U7tsMsbk
JEU6Cd0r1j/Txm88qa1aMgzEHkosNsQZZad3QnWFc3t8LwrYGiThKQG9B0yk/RP0
0N7CLYJZUcTh4rcLeQs0yPJjXmN3f5KeMOYgHRQNoNRNQmMXFJEklCxCQUnA/wIS
AWIBgjb0RMgDa3PX945C3IYYlOm98NGNH3yDZosrFAb2CPOc3v6+joHVZuK/ACZT
HYIqh+6igYU8TyUIJXwqGl2YnUMtbXz17vB7PvA6xUWce8hhplzsEAdA3XzZ+GJ1
3bXU6hnqrIXMVylL2YnBzxyzPuQwKd6SlqTsKf4g58TGdXmNaWuPLD5VMao0h5xf
ftfn8EUFShdF7+hUK1nEIt5NtMhNB3cUJF4xXdVawIGQmStvxGgyTqrbr4apX25k
1YQEbQcZkFEDGPngRBVQMPh6ezrNHtZZFuBHEIbYX4crdfUji8uFVfMNm6IsIk5A
tH321ErfmwdbNhcoNZjEB+Nc/hJJEk0WYoiky6XYIZVNSAtd5dVMPsYOU57AJ+Jz
t665QV3onyfuuWOhGTA4XOYmAzZ+O+yAHqII/mTMYmCtG3IxKwVe5tXnGeTc0Cze
PPd+Hu8yUAath7oKRL8NsyOPLxXiP92xjmVMRqGhVtX5Fvn2l5AfqCZjb8XBkzim
lEZwmtuqPz0qeoiDnBF294sOck1/aEE4pqqClS6bcYdCH2mduY5/kxuo8SgzllaA
ZDurgMbFyIwvZCMuperrbLQsPLQ+726uIQaO+jhUAUhTM2HPmojH+yVP7FaWZg0A
SVQM2ur1JGNhpoHxld6vHndcv/032Y080XSOCVQOXKULSld0vo17nHVKdLrn/d8h
RNoL5rm4Cm5uhOWuGoUc7Y8ia+pZjf81VWmYid2ERux8GBhKhPpM1kHmfjwPXlmR
2TZcH9NNyYaUcb2fA9Wr5FhAD5jlQoMsvskQXaojkJzx0FcppAmgS9BgIUxIUFyw
/ybriWRQhIQSz2ugfKXiyD6CNFh5PPCF4/55N9hxssGWqxEBwb0f9NLCmiPhKxcB
3NboaQArUbmK1mAzEqB62RRWTB1mleaKYJNhpfJtja2VuKEB2CvF2DjKojMN751N
n0LPYcdzYPIxYp0a65cstXKdBT7nf+SHAq2+MyO1hMQfszw6Z19LGdJQkW6HAFe0
SSyZeodnXRzo7W7gE/ACGJZACjGi23ChBYk1nzdDz3h9dPrYgHw8I7pHKJs/7r2G
+osXLv9mZ293HnffNX1GNgLJfnOZWrUxaQQJPgeufQEiQFc8/NYqhZtG3HQp0Emd
JxKul/jE8K3RbjpSSRRwfpbDHayVXsbc3kWXTycbQKbKnSYNzPeZZPp59vPD27UD
1PktVAvw7Z43pmq3whH+DwAYkf2f07I1dqIRXyLw6jitA7i751Iu9bVR2oH1dg4o
1wg8Yo1M6jmKmKyZ3DlTSiRVceK8j3/Y7DTyyDqoiuV0/6jXkgnug66Y+mJxj/6g
Dry81UIcmhQ9NEbTnfncBo9xspBShfvnyhfjZNosqJzbUs0BhZ4Y5jtPLAoO19wl
3Co0775AygVwraRZvG3Kp8AxRSgwaYNu6SrO7KH6OK/je5XryWkzc6HcP6Gg4eUS
wrRnNz9cqjX1JBIMPsn8CLCYKhnj787j2r9aXDbmHNCg1HqUtfd3XxmoKf/jWTmm
am7ie6ppvHoMsHQggfIsZfeRtP8BCeIaCRMN2c73JC86Lhe/4mTfjXAC99DOBJnA
+kDYjO09Y/4FqKAtbaaTevV154p6mYuPG7L32uig6rtkNS5S3BrCDDwOzzH5KoU0
eCIv+AIWFdu6jU3gUdcQnjrhHxXgy+J2TLRSFTh3sqrJr4c8GRf1D27x2JFW6Fuj
lcCO+9Dbg4F81Y6agV1z1hgrU12ERA1XnyLaJ8B6Zz5DnG78fqH2HaGe03clymJj
ng4JkBOniynZzFxOi/cWteGf7uQrA7K+MhXoGnLl2cuf3TixRiESm+4DqXbuo3c+
F0BeSsJK9U9wVQj6jHxi0qZJ0LwSuSQGaktLYVRLRw/YYfx1IJpdn17CNQT1FLJX
U2MPhNkrNE7DqXK0OnH99CSia9a9ZQUjFBTRg920MNwWi1FY+zYrfIYT41KK9MyP
aRCQBlqOqROFoWe6YViH6JOzsXuXzB9keAI2RcR8c6Z9HTFq2kCyBL//Cqbb2C0d
WSZrnugl9G+xsQXqFyyHr89FYG/mpXGfdcFQcFqgaJcDAgaU4LqUgthMdR2rWMvP
DWbxitYtksXK0CcSUYAYx34MYZQXg/kvt/+227s+w/y7U8eax1zeQpxA/pcdem/U
jwSAw1+lHLAtFr1Rd21N31deMEVKVlbUj7RbBlhNkS/DR1wOz1XIgD/JgOrdm6zP
jPJQiotTTySsSnW3/hk8LA+DmTI74cGB5gzBWlZoRzBGSpqaUUl4mFZDJrU6ZDlG
O+Gk6DzFziSy+sMt4XcXVZlxfXMhb857Btdo5YFg6FG+j0Yf3shZbKtizg4rTv+/
XjyRs0DEJFrLXS99jVii+XtByQQfak8WhO87xfSXrlKBE+Gu6mg7JKbuc2VnOA/o
URgIiHj1fVH34M6ldBqdiLO0PddqHM6KSnmjZ1wCs3PsBr5POHZtZaSdyzY7FG8J
oT+6IjWHD/FV4HXs3tNvdpaRz2wxgtvG1bIFJP60bCB5t874t9rJw1YYVs2RWY6V
WjpqLEZ/duCEaNdwDPlS3CrxCEgmc3MZ2dYXhbsPZHsk+JVKND+IbSfO187EteCZ
yFqv6k6r9PZqGwF2OfLh+SMdFoqgmxGGVquv5AtGsac8FBeUE64ghdhEaUtJ1Sek
6Hy2POxc9u9//82Hhft6pmt/Xok7wTRlbZW/++YY2T6+4mmnKWOWAcVu6Xgcjq1M
aoicoETqgSTpHEz3jF0xXfGAx5RSSjb0oOPwJXIaDlRvS/Xp8gsvF2k0mj2P7Rz4
nL/xednPjCFM+9IRswhl/+mdRkRMs6bOqLIyYA+ye1ntlUcAMqHLYIBRTeIQUUf+
0WjN9ZLVWJD7s2nM1cN26dzyjxgMe+UK7bNrti3VErMvaRtm3gowrEPf49lut83e
qrgY3M34ZUaVGV/vM9TQ45hSAJByHu0HCE5zuRs2rTvrI1wqNZYGYpXdBfl7Tdq2
Xsy1p63yD5V2LN/HAbTFADfQjX62vvqPk6ZykQfycVvy12P30jFd1Hl+Q82amZhv
amVe7EU/uOn9xKZcOwZ6/AYI4f6V8KTVlXDRHjxlBQjPR+rr3MxJChstwDxtiYOk
WijVYck3pV8j4Re8gLKMyBdUmp1U4wgNqyQBhIdHut5qPX6h2wgrzeFue0pjdSj6
ZFb7yFrPlLdyuyEHNLtOHfuDgaOG7FmwewVyq0sKV+Jetx+c5EjubJd8cbdOMzOf
i0e4pDIaZlF+0fOHs/ISiWh74EazP5ETVRv+G5I+3eIMTe2eZfnJCqJF89Ez86SQ
P8wV14LcW3xTWmCUay+1Yd1jB3VBloIi2B701/r39yNxhOhzEDMlJY7g12s+gpsq
M/828XyfzA/5/CPSvTcYeeH3YnQrKArjZiR405vpNShqaYt7GwQUxAy5gumZSyIw
DU7c2KVhXTgPohmp3nGmuPt/vM/TSL9px4Rf+0D6Z0DCQQliYRVS5wCbM4rBXPpU
wgpMPJ2EKkNq4IDiv7XJpaViRuJJifb3Yypgx6wfV95Ub+dx1XhuYrCdPYgvMBpA
fU/rm0g4eBt608INbk1gRC4QcVo6roG4alc+/n74xmEqjh0BYGxbcW/m5e9X1Jcn
gkC9iqA6cgSINM0YONnL35bNav/B7hqpUwupIHdnQ9ry/SpNP0IPqtMY88zbEp8Z
blaBaosdCpVbIcVxczafTnHt66NwBWBU5xQBGR7gMrzT+ruA0PRDkEYVIhh1o3/+
S9sI9MUQaJlsaDE3AzHW55sIGKbeCSBhRmNC489Kj9wrGWiPYof+0MZqwfp7fG0O
6XXGageD2FzmxBhSPhPsnmHsuhyltQjcAn7+uAmg2SbOUH6gAnubzOyrvmgyVBH9
0hTKs3QjmxRmxdHBh3PRtHR0kv2GAqc0ka4gD0cP0zIb+Q1C0vsFApodTvCaafnV
UJx8dG0Pcp4ci/eWmFGmPKs8/EUeEWWHc7D5Ujgg2EbRqcNP5C1uRwkv3HVXIRIF
xOWCNOnltmAe2jI9js+r83YbZ4APSGmCAxGxcBp5BgPg+81hIo6KWCdxry2vFRn+
VKngmUDMaRPPGiAReN7BwAifmyAKNx1mDTcOYwc6R8/4YQZNfTUA46c+XkXeEE6Q
75koGtbPBSQOMGELUOtMhQSp+I0oJijS+MRZ+5aS53qNGX5J1wScAO3J3T3c5eIq
L/5aeldDRqjxV+/0q/L7ZZwvemVthNo4fLiELbEX950uIB6g1Ku6M83KnX7+HYMN
tRx3SzKeBI9P9a7b1HlPYGqi7lNAMJeWL5nyyD7kELs7Jep0ZjOorcUpYAShB1TU
4XjcSctIBzGiEbl7976tTR5q3/sLFR6CaC4hxvXNJw3BUIlPLrdy8VdXbz7KmXpU
VZg/RiSbcTjMFAeva+hE7978oaX5e62vMDKS+eI4zT3JWuO4PKFeVrrsWO50UE/n
jmAE5GT72qyv/sGE5OqzxyWu5aO/Jb4SXt7KxHrmqoScmv2wn1AVvIQOGyLwmh3n
bWEcJD6hqvSxAN8QKbkrL/Oxox0aCJMVL72lb2eWA8JYBgjMPLLYbrcWy2aKkbjk
+PcwB6Z9gxtGhMVEtXq1yiwSRO+1j8LbnQupWYIQDGoRv7/J/zR1226r7CUo2IVo
ZVbaANTMTvCc8Jz2qvtA4oW4Z/WaIgk9eaDMCxNW5hTYCXdQTJ3jT0GWnUSEabOQ
VZIkySH2wX7DCt4oF8lRR6yfnecOI6RH3GrZc7SuzgD2YvN+mj1WK8J3vUYb6H0p
yi0l4xVT8741O0oKn2wJlXAkVfoXZA94t1O7Kb5tTRLZkBlUfFF8YVbnGDrx3xPe
uZtWxfhBGKP+nz755ZF7DfnaV6bbnlSEDgoJvqBZGfYsl85+RvVBR27ie9vj4hUQ
YpofiwVxqwdxl8zA+IllP/FfRrh7Lo0+B7lDuRuMQafuj5cp0ebX2qYu8vK44vEi
idZ1O4TVxWHx1NaZb5el7+tcKi60+k2edthMfKvTtnasDuoGNGJe3HLVYolNScys
ZuxqcYlC5CZ1Pp6n/bjjh5uuoXgNQ+RGR32Bh0tKoIkiN1krygL/HpxaUuah6z0o
diVXM+WyYHbn5rZXWOe42H/lCzcS987rQ3nh30JnUyycXrIIi6S0W+QSxXQOD9Bd
xdjyBfJd1Jp70wrUTA3aALSfpzXtkMsdZMxSbfAMXUTzAA4y6Qgy1vdlN9cWdVxq
hxHP0uQt+ysO/cx+I0sPiqFDZEIHFjkWC8qJjv4lWHi0tPZec9gJDnbwfWwScnZ3
B490jRjIeDmUrbZPO/49rP6HcZzC7QFXP7kfJ6xaq/F9oQRqst/orc/sfacZRgqa
hTqUMBMkmxCu90BemtMZoAuK7fKC33SV4pYORPBlwvCAKyTT3Mpvw0ix0wbE8bMN
C67veEjulhok8k+hVRLQ0h2/2EQFPuZn+8JCZIfax27OFnzP7qXZEI1SLkBOewGw
Yu59reXwXEtxlaCoPaywyxfDdmCWft9bw4GhbYd3m1Yvedp55SwJnnefvVbKdygB
p8wc8IDRvdJKKWIwQgouzM240VH60kOvS3YSb7PaJTpvpn69a2QFSTFfiVdQc0QX
RdkN8XiyPIA00HUZqc6KVwGtxfnbuWgrEOFlSByKi7rZBTauDKlSlEWOmOQKK6NC
hpiNPN3F3PSp4fros6IRWQkI5HCRlfeJTVO5GBOA0BCADBV7GMVMnnzH4a2aa1fO
bOmIuZNaC0dAT/j8WtkBoOZkw272cqI/xZkGP/vtgbsJeMOtwaxAuPE7Qt03RL5S
cnU4rrk+9nCmvZfOydxAx09uvjNydXGC6/QZGEvwCJibWYu7gnZN7nKVQEMCq3oZ
Zp8v9CJH1OWjJNHuGyhJxqZEd+qDqVB/VilJz0gRs9iignVQJyenlXhT0CxFbpoH
Q1Lkvkjkw2fQXkhjKN/XVOca8vzqLqlD+ShkYl8uKN2RRnEBwC8A8avcyfe2k9+U
wO91VrZqpPUkaZdGAwZXOYynAwcfi2UEC0h5xVfYtR29imMzeWsW6StCYLXIZadP
H/IUOPaGD4SHbkWMGZCP/A8uQKb3StdKPAeE6aypLItyq4TgnOQeUTcrEvPou21L
SFnT3I4aF/TO67Ce+HeqNG7xSZzSEZ6mdEHGV/dzdrRhHtXhYQlIryzCdNAcy6ZV
WFhlszxWGKc0eV3vAk5pNoq40q2LgTewmiMRhI08fnthJ0fzYddeHi5qyHlLMclJ
mNcGu4Dx7VmM/apvyJKqGsQZsoIyKSh1r/DzG/HgOCRRHSoWQI3fPJvbkte6u9xG
vfU7LxyVkxi7w5KGbyIwqcNFx1CvUDptDRJzMtWOCYiFntJmz0YgODZfwhkBjatW
NB7TCOcrGxMREIpfZbBAMoAyEtTJXl8XJoDukU34R6gsZDNJpZTzw/geOYwYxm/m
de5dxnXPhO1+eRRilaoPbacH/ZuwbTxToS5Vf7IbgYtUNXRoR8nrjQOY/RhjwZkm
MG7RVJKXn9lSc6xsIopeq2SpdLCHhUD/o58Xhtg72txmqFxowyCwh6lESrXIHyGo
ob27WEfyjuJU32SNidRqxgLuirJQXJgFBFdS9/zIurqN68X+uBUJ/DSS/gA2FXeC
bsgsibBCSd0TcNnYtYrpXhZSLrQo7nKvom8kPaclts6mGnYSRq0C/cteLXUJ5uRo
BQGts6hYvP7zQwvXMBAFKuVrhwKaTUQYWzBn3MOsuCJ++VAWgoRQdHzH1Kkay1N8
ZBtfFkMxLWdASh0pAZIpBElU+E4LAbIpYA/e7c3/85nCNs+e1BcBLrsJOXu3Ux4I
OUJ5C87/ugRB51Z/rk5IRnj4eboKN2U7nfAfkuAdMGPQCBLrXcXkLarLB3+FOU4W
mUhPU4+0EH15ujx/s6/Fl8v7HYBmKO9qI67YCaluvOed/NBc2cMSTGCoQomEyZEc
olexTSuL/NkbeUpN129rbpQkoNI3MGOoKjsprsRbChPGAbwywQEOdFxHwAB3fTvF
uxIf18HrbK46Wa3C9GXlAJsyPDj+GC0uo3HK/cXyO1ubaxVX6DGX5p62WNXJG7rl
7Uh9ZOvdKqtm8+kZXdxa1BdGCXs5qNwCdYQQSS3e3fEwUPQttABP4IWhhdf3lZ5J
VZ66lfYOdoED1Mm2mCWQkFMyKIcdNVf6EPLc8fIZ8ojUFDvFoheRZbxjOukIrsQU
SDVq8P8umqnX8piPifiwcksWUU5AFJt58EW5ok2irM1a4KrAs+nHSMWOIfQm0klb
jWYv9w2rrfFgBS/t0XYB1cA5UZeHhJvzu+31RMMahyc8cnAZH6kUbQDobRf2m3iQ
KVUR5Rm3oNHGLiFBYm//+ToLldMMLrLOKZKRdApYAdGGqEP0+BmSLDuqc7tuELm3
LLz7+L0eDUlIUh+RcdTjDMQbQjzjERkuaaAtxvXgMyg3sHQHsVlSJgp2bsdds6xA
17N/XUeZjIhCZ2eYAy8J7+SFo0qBx4Rm9+otYbH11vF8/MfkkwIS6Wojei+NMUIp
tTG33ie8TqBeLV9yOnoMZ8Fv/uWR1bcBl4GR0H9P/zk9UgfdhaEPpwvxAQ0exeVd
xLAxd1apsRPmJ4ES3JM7KpZzFCa6J9PLQ4vX1qj4uwQg6SM2AvUu+/iybEEt50dN
m7VYYwOVJyzx4D9HXheKCu3iJ9BpgsPcw+zAmE3SWFuVi9+FKDeNUs14y4xbMBF5
+ncH6DuVOV8aCR4pNQthge6w41J5wqESqSM8EWfGUVHCjJ8RJrbtJgXPBTkHfvon
a2wBRzbFH1BNLvG+jkaLA460VKJlJS9CXLm3j8LCsadmVHojNOZIGmwyjCm54nTT
1wYIskaAjbQWtI0x3BcRKYnpkB5QFNqgpLL1ZYiCMJqCiSGYH7+1BZTqxSO63/Ce
ofZ1UpE6+mli+Qf2fIh3rYiwWs19HBnkbZ7nLJaRMk/xu5MUdckK6t/Q5MtuwOnQ
WwHCDwmzq605yoBeFZzKHK+jqlwHH2de6M8Oiw4dPKFijoDe04lyUiIlTyM0upS1
s5yr3Gbe7MUCDoHuQGiCoyPNXiBmg5vYJ1svaMxVsCStgwrzuh75wDkOPef3JPrU
/3zGvHyQAEgvwqSB92hCjyaVsvAwBmgATWvn1cnSJ5jawUuMQ03on9ApXq9hNPu8
MQcuEWSMacx+fmkp7jQEqs1ADZ0yJGy7BzBKk/mZWLG6w8N7phoqIVyrVk4QDSfh
9TRK1yoSGmB6dPRt3ZuhSJLo6tTyHmrMNawuTc9zmMaZaoyFtRquAPjNWhNQ4EKp
U3nwUozCJ57Qz5rQuq+VCmsx6FrDIFnEkuTC8ubBCiWwqylcAzIDIeoHBfuSN0bL
PpjTjW68lb8ed+chwaso1mfa1XdXYclunvLwK40+P1effVij9RfnsCQcgiDDbMJs
b6zvflfNDkaZRnAM48vJbA3gYV9O143gyLrAWjzAu3jbszxZQwZRZcaA0mwClAGI
MZNSYOnud1y2lldym8BkIWg57fuXZgp0oaVzkne0d4ODuWlWr5nIUvQG3cswiTKT
u0dIB5X9WFyf3ujzXEkB0SAf+xWgAcQndMPm8oJ5OildbX7UtIXYI7zGecIRhpsk
6x7daUIwdaRzG9Fdg0UMnSMpa6OPjxucYHadteqJhLKf75HyPvAARQRNWNxw1JYg
bt7vs8wSOYXFnG/pxB/12yMjPtT7R5G3rtYt7arhSsvJF1TYGJqc/Bihruw0hOPA
per87jJSHuy5Ol/eOozhTJXN/ZOBlWL8S8lj0CASdzZI8mITcj8f4PUJJNczrbF5
F+PMT5emHKbje+EGXvUxrNEFi8Sv+z1u6GF5K9jDEPElD78F7qyxP7QKpAVhDSPP
R4dSH9GvWbav3VCmKELCEhrX9qVb8OmUonX/kGM5NI/chUaOjED3s8Rbf08mmSiN
30iti3dcgnyvonZeaqcTubBhi0X45V1kUUnCCM0HamGLmA1vp5uNkl9z/vHFRxob
scAaIWaZhPJE0QYA7zXI0FPm41iyI4IGWqPEF8559PFqyZwNrsh0JDAUXAlzQyRr
hZoMLnK69fSDzUtHZT3LBAR7jwhMPi502HF1lzZBg/m7EnUpA1KDB29zI5v9BaN8
k7HMoZlK5kGJgEx9AghrWCDRXQ2T0ZzEYSUZ0mwoC14r8TI+S4XxLM6zPUhiQ+8y
2vtFOFbsqh/rJ/8/O4lYvt+lqdn4uh5yJtlP9a/pM+fc1k5Xj0ixwRmHI03Gd5PZ
GHi4rRZDnxs4fqIISxBpNKlwJ6c8XDWsSk8jSJrHB0McN1pk+AFZPBNPMckjSJHP
PSTDg7bMaZCGo7J9Twbb6L35h1EehRi3ZaKbL9fg57ZzYSxM86ZvuOQRsl4b7hxC
yGU2iG0kxBPdh/Im0hWwcKzvTVnfmpeQSrOTvatQZOhK+gA4tpJlGnCc3e8TljeS
ngW3UzH0eF/Ss+JRKX2QUziFCp357wQl+z3mU7txb7U9O0PAaibttvSnJ1bMybxK
4zDe4pXYVfQ9/B7JwI3LLSm6vxdwdbAx0+Ps+wZfa04ao8UhaGgjfJTQRdRPI+1e
wWTXMGu2ipbXILNLjTIUJYQ/FP1qLxk1zFEd+UT6gQzdQs9UnfxTfHUzpGke950Q
UysrmlWi3gKgEa6uYfDB5XtquHjWPU6ZEEkfuasstQU9VeIvpUjqd6o1/4g8HKYl
hSlDp9oRrqrvnPoblMTQmkS/C+LQaP47D5lcgUJhUFixMcVht7T4FFh2nwIlz4yD
29OXHuXLDQoGHO6rAP3SR/vAZoWciaHzu1NhAWT2hvnhjen4X8ToxxNsPcpc+6oU
zSYHGObCBR7lgg0dJ87fIH+Xd3U9J7z5nwRlXLRxZDw1wKxuDPA5Ne9/5kmQeeWa
iHBEtHVIKmTb9OqiTtvSKKEXk97y7XBwE8w+VqYRX1t2yg1Y9M2IIenXolm0uK+T
SylsYZ0CTF93ajAcBl/Efd5CxQa3Rk+W3btCWMjdPygPC10Eft94h/lBSiZgMKZe
g0XiexkYwlrc7iNngO9crXM24CoDnUP87CX3liYLjoA8mlBl0neE6k6hIYFsiPEi
3CcIKupXFOwa90vbgcY/jmxJ4BtriluE+/ZoKcMQpX1qH7t2lcsSxSANCHP1jf7C
OV4XGluKUqyurNY2NjhWrRFJYOFEFfpG1e87Keqx1OHEsjpgBN0itsG4IVNLYaLb
HV3sF8xhwgcIzIHAGJowRucinE65xV10rEEfXPjTycIEdkKSaIevU//Q2HFExdy+
GbVhWqwUrU/taOUAth0wYlVhjuD2iRX1e3/GGK2Ps4ORWXKk87LvBaDsGBly+OZU
UxU1BBc7e7FYVf59RbwO4TwxobMx8fYtGIXMt7DcIQHkq/d2SyZOgdgOXwFjp3ur
fLqQAV+M7VxaZ2scJ8T56a80Ti9osS3VzuvK9Tvk12yQ0Y0WfdTkx4iFXn/g5gte
cp8psCb/i2X7dbgCLrj6MuFsBmuCFKI6yWaunvkKhgNbXJeAsBfg76SRhYiEosXM
M/VUBdLCoY2OqHSl8oXwhhERcwkCOr0e48ERDB7zXMmlE0CycRudbbVU5/WPeDSX
QK0mxLHrQZrSWMssvld90Vf0rDXwq+Nxb8ix6+KIYQQb8ffaM3w+U/7SPXjgAZ/M
ZyWh7Mr4j6pjOWm966YElkMTcjRlq9xsHHNgmwj5+1hVxfQ1xkC6uxASMIMbtsut
XRhbfXHHL8ZFgRPZk1qabOEn1h65iWWCgUL9mhhMvLWIz/Y2ZUXXYFdHqyWlO65T
uad88Q/0zR9s9u6xUVLHlTBWFoA4cYRGFGUiRE5gNOrf2QHW7FmKgM5a2ZT4IrAE
gD5/5rgyIQb9oM4ysGlw0go7/VGabWtLaUa4RSBBGJxmOmZmS672Yy5AvnrqWCuh
aOy4Utr3L/v8sM/A5rO0bvBpShl+gIF18y7z85Xwun9F5120g4WpFDeD87HmCeuQ
OhwHzB++4CE7OY1XQwR+asTMoZTMPk+kqNVkSt2FLQY3+N6/u5OBKCQcUtqAlZpY
6nCp3G0+m03zEI1yfwX4+flYD1W7/+1uxkdT/aNX/bpt9AQlMGY7ruWU00lvQeIG
RMbvpQpRlGWD3BgIK5ZoYWnp6retEvDuZwtrSpK0S5akQW0H4yrGb9KBFltv9c/E
Iy15h8HeLGy4zlK+ASjnveumlsGZNIrH5yKvggOFAVnjIX8hQ+kRxSIbI/S2mD9v
Kf5NOUfubLok75hU3pIpFzFHLBskn9fTOE06v+4Q6XqburZRZkyWrsRSydMjt1Tr
L9bT3TOGCSdUJmfk1WEPxxP1C7+aHPAN81ViLqCe4cPghtPPYf93jBfzCVfhy2D8
jRlQEP70KTPuHWypgVjHMWFewjcjN9VJqJiwy9qFDMDnJHTQTeOhFdpbjGaN+BT5
xRQJ57K1BV0z6TUQUJEjOwiYSPYdZeC3QIkGpSkIfaXQKdrfXFP5H/LLe8CQD+jx
RYRyUk+ZKezhpn/CZGMUklh6YpeRQkUEJpCHPW1Zaz5lagXlqxhlfR0oaiascNcF
pvPGX0+YsXLnI5/nd2WWd0HYSyUFg9TkdZSsz2rC2pDiBUii96K5PLq23zkYGj73
g3ejoWvJpe3VGxhJvhsgQD3SLCEuKI8mM4MFqAfm/+pMGk2l3oC7CRDgPreEemkG
upZt4a1323jW7KX1m1w2YOeWn4c1pSLgZyy/vj9PJQNKKyzIjRsutpkZndgRKvx/
ZPAnGhXjhOl6C8QxXk+9MAZWSOF26eamPpvcDmbgVv7/6ZAwbnpBk8LUlZR7OWNO
UQBrs1bheBopaqK4IAKKy8CCx8FEQIoQkL0Ov59PTs69tHRyPiFVtSt065z/Oaa2
a9bTcnQCp0+7kh02VRPrNomINMwQMy3PwmjXTvfJp3fx6RY+51G2n1I/RmdZnXoW
97BBDZ9y+G1j/H7V2AzCnZtxb8rfPLk6K0fwXV1eMVTpxe22fd6dBKRvIhb5FfLY
Btm5329nHr5pKXpwarBJrfx+gD6SGgO3efpLgcfW93hCQ3/0KQCI6ljvKwIVj7bg
ox78ABt1QFaFW155fz+Hck0cquXLwNfVZadwzyEATobPyBxaiUhUQ+VAZDxBaglX
G+kUWT1XCAqAkocfg3q+Zl+smZyeZbwvJHrEXn9FPBZdRDWboaKYFr7ucBf7F5wW
jfJYCCZqKxosqSX/fHuqQlOS6Z61gM9VTfPMeiaq21GvC/OWKzeNjMXHEcBJr44+
jn0VYdqndCv0iJ0R4HgRpIwU37khjnhNPl+ymUt9jJ6eavxEANkKmX+0iEqESHtk
m9v9qn0CL32gLgzAcCzzlT8TTQUcyfFMNPZMaNrT5BjKldnl1klR6la9Kiihe7yG
FRZmUgPA2Uj+r3mGlQPr/clIYfvzBQLg6uXA2uNKP0BmsZ8Qke4NZHMYl3zjuoUK
Jzzq/w8keA3sLayGrGVI3TyRldsbUNdN8VRnLVkOzocXL1VgrMzj94dCfkuQ6lgl
WdV45AQcQVMGIN5T8rhxTx8aBJTWsMMZALTc7KYrdJV9VadCNQX2JyjueO0vnfE4
IYk94akYpJJ0q96iBlAW73gh0xWNgB7w6t+yV4G66g4gG3SKrVvJOoOYAPqrUQ6G
/1wnY6N1puDPCxfMBJNacrf+MzF0WFNo6qXVFbAGnsWHLGmglLvDl3rffFJjLox6
XK6w7gfLTmzZYjJAcXJq7JqrcqRIxe32D2NJDA3CcAyNZGQJqqMRSoGGWj5KOSb5
8dkFf6zhZnSA0bbqOYkB2EI0a0WC3yotNAjHjDHwufoBB+L73JlCg3ALgQXJFN6V
2etfzkRWuB6ZcEKV+QvTXrWt/Tm3uSzciPIQbZt5kfi1iaYrtghx79k3C2g4KdEw
AYxXZLDjel4fOnNd55sJ+gWHqy5Y9uGYCSNPSWNjlDe9PndN9w6jX2KRtJPsyTp4
0TdqKrnpnoaom3SKNcBKb0VPBvGumo42xHaxKPGXmnr4IKecSUozbEOyjdbwvPlP
3qa8q2RgMKaNZ2His8B1f+i0VP9Q12wCRDhdk0MzXJpFRoSroihf6weMg3iijVIX
2SfBqZ1+RKAOtO1Zp/C9j8+Mzd/XH3Wl0s/T/7Nv4CASEPihAYkTW8yt/UwVWPbr
8Pp9wbxEhFw7VaOz9CET81Z977sryZvX6exnDHruDymjeMkpQbeEVCBUu+q2EOHs
ZiC0iZSWz1cQMuTgyuJGXEXxReM02zuZFoGIvfVuln0Wkm6pM4ym19e/AoT5PtqS
FvHR8Qaf9Q0kGrsa+CaShz5mH0I1uaKqThPl6A3btfx+6l+5zwFcriLgVAzfVf/N
tVvqpKNBOtGMX2tqkAVhqJVjoJ4zOnKtFmaaJP6F4LG9VvgsItKAmCabijIPlEV7
tY3Umzq/PZMUIHdoWVpqi9OqQfYbRLYh/43ajaL9GSehbFooZCoAUaE5SPyVMJAf
rDP/H2KXvuxZuSfoK5KfHCf36/4YOU5Wz35Tf8AZm8Z/YTQ+X1Tcm4hQTSnZISm4
G5BPiTbVEiyv1O2bMy1jtpcTM3dhJxMtSfYxwOWGnKn5exN3oKix+lK61u+lXV0B
zZ4Y4mZjGLW0/IeNsc48U23fcyopPV/w1MnFK/XMf6QIOQGu3dIGZ5pYdwB9SSYw
ctq2DUxNG/s53Q5YtL9eeRJKH+4mMZDT3Avo1Nl4ZaAiYz+/LOZh9vLS64XzjjLl
i7PPcgWKENIKofV5foPPBHBwefhYQaIuBf9fmBBSI40cwpDU6O002YGWdLOk3iIZ
tgWS4nVD3OLrmAxGhbr+eMw4M09G487YWuHXLn51CnbKEM4NWaEiQhe0ex8oTgWB
3QuyVcHGKua3XSwG//OGy5TizoYMpCOEHAWFEuJdhNUE/9BVcSMbnOlumOo4zf05
YtOWv0QIk1GE376wWo7GQuZNGhaYpZgrkOvvkKMa0dKZzF4OQqOINSISTuNN/ctJ
eMgsIxNIawGpeO/hqxd6ZQWteUIll4vKu5Og+LLhTVCiByoJwKxh91tUfPIbnLMM
LT3eCYDXMDStcXnXeGQEMNJVbJI+8L09Ro7HCZzN/sKk4euqqcbbN/Eafti62GUo
br4/WKZs0GZAkidZYah/bo1MOwvxX1gjg3w3thy+e+LqBxplILcM9isSNii1bhFb
k6Rr3nJRjcNfS87550JOvfHtpR8gyoI1rQN1vig2Ox4TG/9U4nOhHji961SazSMK
YeioB1Im2QPkt0s4eNfDv8VAb0CTEHIno7F1eylgwb1/kcXkU0y92rW+NFLLqRWC
VrxTxmz7jvcBmXK1Ky5fke4lXE54aMGIwLWyjjWIuEER8taViDFPM6rf3HHAZ7Si
kYoZDISM1IR4FfgI3kDeUwaN62E/MAPERNRVEly5EW5nRwM071osSLK5pye9dyCk
TcnzFEFC8VHBvOjva9jS4RlHZaUCJz35j0B3M7GfBVc6IIKw7RtzbeO1IvtvvAOq
Q13tIDnxNpIlqUjEiw0VOzs6/v4PQwKNfrKxQ/1FXZWP2lEfUS6dR1QRbi/qSLYU
0UUWR+r/xiwAhq+lB65ZV5DbLCwKBH4JYlI+EnR558Smo+YZ3NNTkG2fFv/+oUe2
ixM3PJ4OBfgphN3DAC4z2Gysmct/iy5fFQ//mV7lomwa3wNEWkWW6B2wy5fzVIHS
Yzaiv6fxdnJ0vV+7g540UqyF4vSWZ3vlL+XKs736SRt/Lf/Dm8RKfm7jiNTkP1U8
noVrHV2FaH677j4ShehZhENacnEa3ZgksvIJ1g9ftR1Y1NHBH2bWOSP4Vp+uQWY6
ZpkBwOVlIeRUFsVE4eWxWZDCJsjvCfnHcf/kIQpOQJofx1jg5vzLECKW8/9HE9RG
3aGK4U9OJDEi/l3oEg+JzrmOK3EBnbEe0DKufwLhtp0U50VytG+qP9mGa6DO+Vb/
77bOcgV+ZL7SpOdVX7r/oSThAgsoIBTypGV3JgFu+DczhaEU+rU80vqtMqQhdYGN
5Z/f5UUJI4lJx1POeuTF22CWYzCz1a8B25DxbGZfId9zzGZjAFTDVb5qHZ7rQ+sK
gaRNwFoH9LYk/RUWUrOy7GKnqwnMHCDFLpgTh+5AwJFa//uQOkfo1sxiR5QnBN0A
7g0XhbV+aakc4UEI9WwhP1zDrNX+LwqEO6l8nJHi41w5fUsW+SjXv4BEpOWpAeCH
hTbaIiZx8Qyl7tpP/b8HuNzy9/3PxAXoR3AyV9U3wjomvFuovhV8n7jcFfnKXpcD
iSqfUZAF76cvoqzcviFB6nIKgPaw4Q5oH5H10OGMjWkVYcOYbK9Wj6Y4TibuZb9D
edlQUrhg1hqvvcYYtVEx0+8FmMimpMNDgKAJNsvBnUcFCyigV+56WEpK91B4mvm5
HL29RV3dtJu9ohYGxjv97Zq5+ZMLV9rveJVH//DmVfoC7YqPf9ihhEGeHwkNW2d8
R8VuaRDbqF2CVRnlrdwZmVzK/FnajnEhEw7dKgwjzFfwWKAi+0Mf4pbUv5JXQoRK
PTlmdb1bQwBXVL+Wb5jzHyuKuiJplQMPbrmdcT3qj+nQ58f367eLj5jTn3Zl/qyS
FPCW67Rs/wxIm0zB2E+qSKN0b716TvIMlh6N5pHfi5ow/AXSpwrFeFdt1JzltKAp
IRIAt8N1BIEykavsHqgPwkHtgqz9OyoaVikgeGlXnMgGFT2gLCapfbnXMtiF62h5
KvMzQg29A4bP0Q3iqKy2KSquoa+a1Myb4JQX50vOe8aYxixSUBuLjGhb4NMgggYq
pbdov0LedagwDkRevD0XNyojdqa42QZfOasaFoBsG80hm3OUEAa0YY56dAQV1L0v
HFvuZkEjIvayUh0OJdYTKO+uArPo6tTmpqZ7E2wBEacjSC3Ey4jUSjovBXB21PHG
Z/VQ+KhgJ+IY5sgmLLF9hHXyysJQI9iZczr8FB8CN0pJR1zJ7N9foiUrcKTM+vov
JdQOClhkJ/silM2LtMoIlb3VHH0DlEn2NKJ3x+qh9dO3Xcl++9jcbs0RwTPHALTD
syn+LwvWxnmHfqSXRDzXjOQnO1kYUFzWhzlpevzw1LAhUxT03kT5VpS0QpOXc3Nr
5qVkACNHodZfaZ8zGtwPgU9QDED+7L3nNDgb8hAoy5eykSso5q8Vv0Z4L4h3TA+M
jyt8BBkCMdTEyKz97aaxBefLsooynkl9RzlJ4ZnqCxZc/am4QFR+Q+AGOOj6dWu1
VPJvJatH7n1pX6rEmDXRKjEG17BdJmuID5HiqVlk9ZdARE2grmbx4Ki22WNpWnn5
Y8jKoHkjaEjdLOKKCkOWgq6Q357/Qd4WmUvsK1BEmzEuAwwWlTAoIQBJxAZBsPG2
1ayZDz7RT8jlAccNHLO98vjbm3l1yNq/j1TQXNctvljAbiawawL83RU7R13Tl4SD
VNcaUKOs2Dx7vk5ol3UpIw9QV1tt67T5ZA2vuWvtOwAMudY0AWqomWP8KYvBVLJL
pAh1HT7XB0Kqv4Hp5DdXpGSKu30Jbv3yvnG6sWh3kEZxQiQrD33iPO5kD+Bd5zn4
/76WYxvyIyVFdSKxaTfa42pgVn7x0NtEXCWTIz7sg/kBYZGSathH01AGLMkQ2fO/
xmav2sFr3w4unXWJPT6ip7xrw+dfl+9F/4V9wLb21lEVJNbE6VtWh77YgOHi+F8L
W8wEpXagVVNwO6CFUNayb1LRbFi932EM9LtJoje+7yE+i0aWXL3BDnrMk+kIdUkn
+WJlRwKmd7ujQSQlwta1CfW5U4l5ej9f0iWXRa6EEdy6FfEG4SRwFCQ4DHPz1Bpr
jCg8BGa4MxsXFVCNDxb9cwvOKz4xx3r3rGP79acAvxGO4ebrRj13Z3bfLAiH6V1M
J8mU3ji3a9jIXX1KrYWGQ9xtabvwXCRl0CJ60/U1EXZJLFxftHcebNcZzb+DGjoL
tcy7npEZo1u2VA+UpWa8le6VpHS4QO6SOlG54INOKe/+aZTGNgOnsr+p6f4EcAa2
fwhGg6Yj9miv8C+kcKlOlcFiHru0acuXGlB7xtt2pNqK7nJ9k8+DCdsQ2FmBTzti
8uAsA9Q2oFl9mUqKB8HMvYmZ5TKvk5WWohpL8minYbx7hIRPARem5YGkUWQ5e/7z
OHGQ9Y/OeEjrZtfbKRdC7QnXobRnp8Lp95UNG84O0SEj1khA04NpfyiFND7UI6Wh
w+F1yXaSMp2QAAlutVtvYlNVKn9seicRvdKyYX3+TtpjSI74Pb/ufziQXzf0oJiA
qf8xyeeZawSPK85z5yZruwq7OV2yLfKbdeA4Mk5ozExiXI2BdnUB+r1XsQSZPogl
SnvaFeK2J+fqISklWxBjNnMUzxYYb7F9q5hhf7DEkd/68NBTCdW1bpNwLP1s5X35
fmxRvoPB4qQdf0ROUN+WnAjgV8AJ19geFixs2z1J+Q9TR6Y58BZ6dK3bKC4UVxMX
MpxjMimVE46kIs7CnCgB6cFKdP6mYUQgjVBcm6aOEH/7TjKSLGKQHipB2Uq9kI3a
WEXxt6BhW5S2tpZop4J61pQNKMXVuQestW9h5TzKCIZE3Gi8Wa5GAvQfWT4YoP6w
9D7s/NZDnkzsyMmvQnkkfiQZ9SvDuANjfWSU6tJSOBnIKp/R6XcQLB7AK9n9gKLd
sCv8mGuQCRrNDjOm3JS+4IC6rEBdeaR4uEbmtT9ZHR6wlaNQvIz34e2p5x8tNPcB
pvl2hHetg7RVomlzS15wTdfIYdgQyD3MBx6Pm35dUOedccfWaZCLMQ2tVEAB5k1M
kFdgAJv8igiAKituMGc8O5o8225IvMsTidcgFpynw3JTfwffn9v2JKeQg6LJ8zI1
AnLcQcZlIGG1JY/PePNP8rzJcxEaXkLaJljOU9t7HkodotMMdZvaCGtWulAx5ToZ
2dXu2j6HwNUV6HnSOB+imyNf2Ta3JAAmr7+1DPduFNiNQ1+/AqPD4f/L/3iG14HE
C+chSF9HmtjSeFpkjoG2OAOWqQL6DwRqIGjzyI2S0E9PwkgQ63QSmGUmNQYTElwa
HO6R5X5zZVtJXV+HxbJ3Zdv4WztJteUnZklb1QAsd6tHGLf5tXmPMTS9WZcKucTe
aklugEEVTMdxA8vSlN1/uQDr6eK1KMlG3+2fxyi5eRHtIyFpM1Q23CEVeatJmtqC
6+gWLvXGPDOkDnQmJOaGIangwb53+927cI66DUvIJuu4VvbLkUrtUzqqxzUDW2RV
mPxLQUhljF4bfCmPLQVAkazC1V82LD7ojX/H0yrGGbgLWYyns75crGjdvk44g3Bn
28/mr1UA8zsF8OwmVL1kDBHCb3o1MuLo9cl0rIvSAe5xQkuQaGMse/y3Qq6rqKyZ
+7VjyBIM/WglUsRqToMnieIUQ8ywCpF5T7D8FcCKtGLr8IkYSa4G0aImGwgbQHUD
TQNRDD++qsEVcaZTX5TvfIepLBWrMnAUYtikrvfUhT5KB7uw5Tsox2HtbP4rLx90
boIFKi+Zrodc3+jEpXbjOLRT4XC69KdeCplOTueXhJstWyYkgVmI5tbRpy3XgiLg
HLspDeV+kf0BOC/H+WBiI36P7ueBFfMOUDE9SJ7YMQXAb6BhV3RR16EKkppCdwNP
bgWlkhUPzU0SSQqiNoHUKc+anvPFry/662dj8AZCLjICq0bxmRZQJYk+906FSZvn
GfGu3HDbi94kbsNGFumCNRjrXfTRjLHQcKM4AOuVTUU7HGVsE6V/JGIXbsCHI2bl
QjEn6I7CHBOEhTSstF961kxaavVtH03z0cJc3jiCrSE/jlpFmRe8syP9t7AFS6by
/Qbu2dFm29sXPlo2efqqx5HKU62jd7223SWldtoR1IcW95vX/ffUX75Zy7scgt1U
329/1C0mFx5zZ0TbuPhGikUaZ2FlTbnYitUVaFuy/QKvpVYG4KbWuiyNepLRDWOM
oEblQhCko2TSYqCzDOaHKptSWhi7KOaOILl8cfg4TttsddXf3qSI5hJLi7ccPdwo
vH5jXwrWbSCr192QL9NQSvRRfhdMQssH4hHPKot2OwpQULT/FyH1YSgCyMnYLwfp
dBJv+QN4LMWJh4lF4j/u4RQb8e5BipljL7PwwUOB5H9AnvScSneugMCzr5tiuT5k
uCPpV3Tl6o4OjnD+nGzzegZ0TlmcDhGGVpX/Muv8HrsflrY5BhkC22EzI/zw/NvU
UZ0SGcFzp2qb0rra1AjCnLlUPkLVjw0FyxOIHRV3W3NGn91UIDYDHYKJG/SynqT1
iKhApczayPpl7Y1UuuOko7yQFek3fgVS5Qe5YENtw65BqH7HnyWnhBzllMyc/mLZ
nHCqGdSjQrf9IKR9Isno2tPxBMiK5PwUaM2194qMoU9zcl26u93d1Z2TCa3p8UyD
2qUAzHxqL01hGgYua8KsSmu/y/tRU8abgIu56BqpBC1Zi6FM2iD+MTdcJwYhS7gu
5DMGRZl076BjCTOpxje/gBukJaFAeTuGfA2DtlX+ltDLAZceEjNbqpCUjtCqRCix
kjk1arAWWl0VJh9/Hdb9p5uRLyOsd8zthgLvJQkOfxMCZ+t6UD5lstVRGM0BRhik
onDehCluUQgGkOF2KvihJnhcbfTyBJ4t19RYrR9V/EeWzf09KTpDsGpgTdjzs6xD
XY+F1P4HJLzn4RP9j/Y7DS/HiUEmCaFc2cU+06OmuS6JDnVFTdYpPwdVO0hToR/N
ZhTk5nZKY2eg2BvPXzwHsXIonkaVV5Pj5rtPCsWyg4qKeg6iDre1Xa4KvphYBw31
vmViToj7kLXcr+7jO1YFRHwFRNCoV7jtPLpYTw9iL8Xf/UCgm7fOkqjoZtSo8pql
pK7/ax3ryJGw5K8tJ9baHYsNig7qHOOFONNTHItYRXL+MW72ZchhPhbJIMNqhhTR
hAiPM3X9PdqC4ksAfk8Pu6It/JKrogLtWHH8xL9A/plQhYWKG7N3KlHhizzBNM15
+vzMlgXYxfaLDlcE/l71I8hNSwIHYjWDt4tn3xyJu8XR4u17XIdI9uJukENvh6pV
/9aHDazFZjjBeJAt2jocQAVAaN7n7iZ5nVK/jKkdhfGirF3hs0J73pliuXLncMV/
doWFYRktZ7SjbTkzks0xC7OiJy4vxW45PXUBpF9XNoLThyrQLVhzj+Lgi5zB12RU
jItjyv7LNoL1eUq/OSZTpW8CppFpcQiuxd5HsoHxNs4fGLjC8QDefimUo2ldpM+v
FvKJiA47bmsXJUhrmP5/icqyaKoN/69JmfNKd+bHFF+1maU14FgelblrlEEj+pXz
6jSQpRhaSSz6Kp5MlBAuxfEl/pOQ8aYbkeOPilhsrRcCOiWmTpUDN/JUbE127Po9
CQht9mmXwsQpyjWyVFIFH7DLelxY2MG2go/xl3rL8HhLNDS6xfQr5zVxzQHPco4f
DU6IEgMm541j0vNJcf+hHkO/C3WT8bO4OhJhYIPnzT29Nu9FZriy0x8jlE4s0Sja
L4/dAjHCHk8lEts19T+IqvBgasY4dSSmuDjC2pVhTUvBuR/X1i2duEwyUWCbMMd7
mKYFAnDMjN2JVTUTfxZadhPR7HnoPGYBFI6/fhyggB1mvHjbjcTqGU9NB/HjzgZp
JFJlRlq+CnxLAUPqizJZUYRH1Ikx+Rvm/aQyj2q9rpvAwseiPHGNEW/MwSdM1qkN
eHI2pL/TF9npFPrMSE/6jOIHimC7jCvOPJNFrEbpYSF5mvJ7omLZvdXFqg4Sm26X
DNwtKR5csMWGECZJz0LT8O10KOHQ+lGVDkgSiL+5vt7NvdGNrMzt5dPVYk1uHC0r
9f2MoLfhq6Kmt/HRe8VWXBdqLMMREa8nNPyaV9Up91XzAdkH1gY8SaKpnnaP1Twn
9E2jtx5+Jki9psqXSIJuo5S8CedtiGqQhbgdKFs/N1fH7y7MIvofKJ4TT3lpmuxR
yD8JZSfE4fu7/wkuwFTemTSS9sLwTfhx6PQM3o6f1Vy99Ml9XIWLYmVMebVAZZ8T
3EWwOdR6sZv5In6k1kAT3ghrX5nDZUPTZ2faHjwkmE7sfIKCwmFfhF+oAXN9e/Zd
acewBajT3kxu88Lm7oWfIRn3K73jdlp9XOyU8GZKZgrXmkD9nXEpFzL7/QKNEXHj
2WpcuzafZkALs8r3z5wYBSyfjYHw3dGs0ASwfyiJg+6eHnQ/FqiC98VZq6brdU7A
ODU57R2WFNHuA3M176lEa8Zuz89tDnyPOozHe8094V6wUvkd53IA0CmllrVp3Y6x
NVplBLOyCrpagvhEA5SnDNHhAKvUH4l+RB2/CZHSypj8Ybq3YHqkMtpErUoiWKp8
b18vWJFMGyQadcOM48ZbbI1ej9cRjY26QUUE8b94O+67Aicov4O/58x/7yiPvxzi
TjZh2SYXQkouZY9ssMtsX97Zp1zOQSxsS6K399pPi6HTQAHXPamYboR5bC6hLi6x
UWDL1DCaBn1CHYB1ZWggSYJEqmhRJioQx6p4Qlpb3rRNgjYhYJF0gZoKP8iQuZnW
oxr4YBHjsB2Qm3x07yrlw+VzMqSHYpvI9K+G4pp+ulSi5TR/Tdig/rxVphKXCpAE
CCog/AMURCMNbsaqBiJu3Vkbkbxe23kToDgRWIEDzo6Cp4zQnRSRgOL/j0aIuDrj
Y/pQF6HT0VzA1n+aIGrV91lby4ABqMMGS+SnjffZK5ss4Ln+PZNFxWJqQjih16Eg
/aZ4Kfsi8oiONEDJdixa5Vi54wowxa+JZQf+m2329a/ZgrOqIQVIaIV1mU/FLXS3
hH5V6j39DYqvJLNWCUhENg5R1P3M3G+1eeiNigXVO9r7zpvYDA1PWqyxCzgVP853
VB04zkp8Z441hGZp4ngs+KHckaUaqdTcrFkcUyrADGrcFMtDyp5vcvHt/jZSfI/I
GKIEinyW3hjDSQNXtbRuzYtAnTTyxn2v+YIfBndSngD0TcYlItdMyS0bE0AIyYGU
Nt9UGO+K5d+8/qoUUK8p9a7Wp9i5DW5VzLxm/jqfCdzrSkuDn2zCrUfsJqOm9Svv
05LfYMeYgEcMN+5DTtS6p6/ZN+GzMZqe7JII5A3FcSDCYHnbdZKtpAjxp6w3HxL2
zz70Oxc+vMQyUzhMkiUKNnwR6S6/HGy7EwqmpHUhjfM8Q2eeKpIJP6654cdAzlu7
Z3/hJBts7VuKAPewcFwpooKTuLYQnvNwlHT09B42oYI5MEDfA8bvwz0mZzrOQMPp
WPlg4fTxmt33he7O/Yn8fQTs1HbLzxtX82kJpY8La2V3XoaiO3tdR/W9M48xaO/E
7jB/6hbjYAj1RKUYZlwVZcvvvsnYrksKb7cQw+/lF2hL6xZJNM7OC2YPvxGLd8GO
BxBRvaD/rmkBy3kRZ6XbmPeM972Taf1dsK5i7Dga+IX1lk4PnyCxN+BYxM0uaH3G
/Q0B7YNvRs7WmtTGPqOVW/Ym9al6JPU+DOFfW3VKHemXhBpC8qRcyY8JZgSfOpUi
pGpo/CQVa0eOwKseGnk5nJ2azKUkpXdMn5ktF3TbgCLjWKqT5oxWp4kbJzLAz66u
5UUQ2hUqMBhIvrA5zjBaleIap9odlkWUgYAWYwwoNE707cQL+jUg3sQuiEbz+gWX
B5521QSrjkYIQGgcljJ8M4N+sXPxvT1pDiPkQ8TUtvv855xuJzq8C7JzHMi/wxrN
RVCIdRHe/20ZARryTI4aG7VJwpPb1S2GkIkvcoeuPCNHBQJT6HWsXksmrKlSJ9XI
0eB/IXUke6D8kVSOSoNsAH0OUXWYy0M2t+sk8MAsLb8Mqk4gQ/aRNdb2IwJb1sFE
DAC7Bs6ZWaatfjA/xLOQXEJ8bXn8XxkgiLm67yUmIoSUdroEsGWEJhnVAItJ5f0K
CwDWQYgoUKL+U71y7ZlN+M618VScjh0jkcBoGyuoPuewswGdnRwjz3UnGSctnB2u
HZn8VNiZRcf2veqSM9RkaG9Fu3cuAbVwAzRIF8JC+vIyx2tEgXodgGJXJuFCnmKL
RZ9LfXjxSAH7/Wq5aLk1NDAMEoiO93YVcqZ0yN+nu7WnZ9zKGWM5xVc6OtmmXrGh
V2nESqiILwUY1W40bcG0YC3QsBDkOj2S+SvqBhHiyCj49Kh0YO911DJFbWqhG9P0
CKVGcPy580Rjilhoi+MImgLwK72SE9pRAWafeynWCeQErXnvqRrriRFFuvbEPy2I
u2X80UuOS/txI7ulV7Cg57DPghRKx8OSAPJhH1spWfYtB5ujirEAme9KdGvH4LCj
96TjtP3PoWO5mLyBn0MmCznTB7wSCPmc+h/K4Ymqh+ehmbOroPw5j4EuikCiE63Y
jScwwY956IBFr8TbfVPs+epjzdLOUL0k1AN64y4b8JMvxZhlTtGyji2jwofj0SLt
ZQw2AIM731OjVN9Xy3a+zTRjLKlRQx5JXzHZrXOPd1wjlExycw5DbghNjFRy6APr
BSXbvtULYh7O5Q3zj23Y9XYZlUGfjr3mwVli/Mz1OKta0TalAfEErTJAW5GsxbV2
t5jNg50nE5aPyxvtnD7SWjF00/EfpYJ95aErjluN2JxayIQ1dQ2E5aKe6Y0tRMEi
cVTS/cItrlArOGKE81wIxKIyQySK2UhhtLjBh9Q9EgY2cZJX43UhbG28Zj2uSo1e
B9S8/9Dl439qzXLMTM3Eyo5nBTOxHoTJb1X8Xwy23vNspasQSFuPrKDEW7tzeug4
V+x2USl6w/MpHQmGgO+QPhw2w1HyE23hweBzGt3l9TCi8uTSjTIyHlaEqggVCBG4
LODhEZmNWtNPMrC6M1JQmxytXgeBZSUaUEfwqrGyJaH3bovL44nzvyEvzQ7OB/8Q
9QrDgntX+cdBYlrHysRafntLq9To096rjeEUZwooquxctAktRkEx23ORkFtJSkAY
d0xBjq4UlCtwSQekSRApW6lqVdaH6AwpS4rofkPfuk/YYML6pDAGAxyL3/2oaf1T
Yx3syF3O+LDjgVYJMO7TXAJh6JkKhRDnhyNZlU9tx/QaG1PbQFGYSWwcZcBnZQCr
7/AJ/qSBSjKZexUtEvj1CGJ/hGwNR3c/dwYbnHCdoHOPusu1hi9oGUznoiEMgqQt
UqeuPSCNgPxLIUso5SMTcdUQrjAccTML7ByxRmLSg6yonFxUYZ3ExdrJdVPhQCsW
Rk97iODcbTLYUNOXL/gf9gTJo2La7jcgqNc6L09ipWDoDScZsaQR/PZaTosR6KJs
Qcx5ttj0onkJXzvElBDisqvNmv9iAlqYZ1hzMj3KWflwhIbI+XN5K3/8p++/Ldye
++XGVMIIm1dKhbcqyNnOz1wDGsCCHPfKkwEEQLfobbTnUIRpEPsE+bk3UfcGYVB5
RHdtrsgfbFQQsSDxM6XKYuJpQp61cL06YNPRILo7EbGhi1o+xKWHeK8I4TRovgGT
4E1m8Tc1cyxbMVh+A/nyNfxR7viSQ71lleWEQ/qto2USO2b7h25vrt8JVKOixO7U
DT//zGvU2+Jx8h8l1mWPI6Y4JkrFihgVQv8QAj6i6vDDXkGK/Z+tQjSGeD6DhoIO
yxQU4RMcL5WSDHuyh56NwzxaCVgxzacs509Q8KuEWbRfTUvFpF0Tzx+R01n96lYo
RvX5s/CR+oUkc8wQ5Hgxva1FS2483UpUU1ArRw8UrdEyIEzQ+D8LlPOTjvgcdZ9u
YEedGV3Bj8p5fY/XVC06blmIEDcFf1kDgRWYNHKALBQAE7/KFnTZVBIgbaVsho7c
WLook77m4mvZfWeg2H1WlPwIXj/YFydiZF4DlnajyNRD/F5CgdIgkwgZa6aW7tTW
59ZH+xVqlOiNgR2GQ/RtDzcfwkG6ZrbYvPpnXCMSuKnEkgOFYsEUFeRodgkUq6Ck
U9tFqdUJaAOx1S8Yr8X8ZnLZL5AvhnR0dN7ux5QTLlF+ZgJnlkHTRgJbQL+V98en
Lox6aS+E5KHm4VIVfXb0n7MZXSabbY2I5UZ2zvKmmglp7ChRoTTDZDXF2BQ5sWJ2
07O1hkChbUfPUkwD11QfmRe8oKP7WbAcsxy3IhSc7MH1eyBcxu3PztQYivOXU3Kd
ThN5o1CzFIZIi/LwyjkNqeR0Yjxt5zH0ja3gGyavDfuqcyXt4ST6zzG08S0Zj9uA
huXH9ImCxWK8vKVA5H2OkGJjXa0bCUS9bg/pedRJ5bX5KetWXyDTaBJKKn0BOWlS
6FSEzGM0G6rRMWAyWYCClzJN/kMvX+fYPPbAL6+AE0Hs9AtKKzwfavgZ3NdIvO+0
dhJyfY/8fsDz1JYUGn0Ekw1IpyUd3WqK+srInNc6xkQxWBXGztVaXgMD2Wd+5HT2
xOGeKPe32ycxHrKuktPT72hEmxO5HWpJBh5EQhMqWDMg5NeXHE0k0I1ENbzgIAet
BkQPYFid7ZkcB4HMjEWAxcylFRtQneTZ6rZFJMpX7Lp4Wp8Ve4sWK5jaQD19k7g5
jHXpIsOTJVlXtBXUc1t2Du8KYWFWn/bnn9Hq9jXLUPkbzBKqXvqDsBw8smZVkNkN
a+3MwOqRDxQ+nkwJFhfxP1PEHg5RUEezl8+33Ele5WYrXw3iq4io2yLED6OTZY91
tMYrdkG39DbYajI7Ef3Nmf3hZ0/W+lLPmO+ayqHbDdIJdu5e2BeSoLeK+YPQSi6A
UCBYQmM/I66I4iV9AXLE0X6KJg+EmUQZXcXhGAxIvaTPpJ+F2/WQlThKjUBAfuG3
5JV7O3PXOb7YgFGr5ZtZTsHW7/nZZBnlEvSebXIFgIEuXdzS5hRBdlfWVOir45Ff
Qc+8Wkc6Ja4FWJ+DYZCsbEv3LvOnt0/6PrGiE51GJZnbYVLLvmthrLKM2gMaXcwl
4/uBmwKqvsW0LsI7itqMkOU43sIey8zGnksFHE+6CIi/3eVp1QvuQDkXZRE18yJH
9vcOWCKYvW4w+KP8LgbPOIZdwcfwrTKMHA//clbe0LNSMqPPUn79RusQcjAHvfyy
IawwGzP3/YKczU9LuaKcWfQMu4KqcXEgHcHR3xaXLMrwZYpf2W9wll9zKp7coUkF
eJ2cNYaQ0e4ABZlK/u2vYxKCPhm/gARBl0SYNLjP9jmDqH3nB0D/txLc6So3OlmX
s4/kbDzC6o9e9SyRDLmLbLD6j1hLgCUvp9YJwSJ9VidmNyL0iEQVZZ8nqWoI6+BX
2gUFiYwc31K7iGWnedyrXQtA1ki+xDPB+e5hpPr9t0BpAiTi0Pad9wl0u4T8YRRA
9RkUoyTc2OjJgB+zcMWlGOrGEY8253U0qxoVJGGCLxmukFeFK0ZiEQFd6WfauPNl
4NfPYxh5DH45sA+8IxnpNI+QHqtCUVReeY95SpKW4c6tDqgJEptiHUkQMp8dTMzp
PjExmMnuZ8hoZAL4S0OF9qJuzaHCE4Q8jc0AgGVi8m7Jy0W4LeF3mP2E+FgrDW8e
St9YbLazWuZhrcl6ZMQtqeY9WLHGS7N2KoYB6Y9zzLOCxh84qIhrJTgDqgqTfDIc
2IGiwLGrDwtv/av6JcNBf1TNaLTqnnkxHeti35+uuBD2LfXKU6ix8/m8njE9E+Ol
PF1ffBWaiWHobeEZO3UJGKeLAiks6SZOdPAhFzbPIWzLfdJuSMVGV/AqKn7oeO5A
qAXG6y8yNKHqe3wec7G5ZdX2JbbHLNyfpvndiVATjGTO6Lk7Vbtizm4mQ6miUgCk
iXzD6tjVLVzeWliZyIZKVjd4qSSNQItMJFnRUkeEHaz/ytclBt8S3coIf9RcQc2D
w23r6reMqLgsXRX8I4gsRMCu+ChMvkhO2YRFrK+8JZOrieX7EhHedzh25I7BvNNW
XOBUl1xKa5NJvWGMIwxmuXNpn4rLRLaMGXE5SqXnb6WlCJK7gnw/B6bsOAcIkPU9
rZM9GuYnoOgBfeaBB9x8f6bKxq3RCryZHs8NfYL/YIrsdunVTtPT1Un6PQ0tzt42
gDZKZqa8uYGC4u4Gr8oLGYN0/o/lPBB2yxx7RVKdkBRmsBrk/sCJ9wXrKytjCCUZ
6ptcqgRc06ooFv7i58D+An4ZAYo+AgQ3PnLYb1hOVLuLiafLMjngVMjNWCxnk/h5
d2VPMqDeV/MhJzt2MTo25g+HSDHcHgzcTiuvWeQfaMl8SVZNFqn9nEv7v8LsLMJq
9nSxIrKq/VCE0iFyDEReGBTZgxzc9CmHrQ2Xqr0GswRgeP5uyj2u8gooWFv8IASn
XEsV62JTYeIrWkqvQrdv6GBmGu83NU9w9jDFpSarOi6gXcZ/tJxjgLT+0mE+F5Es
p0erFgy11HCD2Oo3zevuQ7MMXz+u+zBVNZXxAxD6yeY9MH6pO0RzrJDKb3gxs8uF
ejDS0FivFvmWsOwWsav+gOhNDOtHuwAFW18qu6qXbWjxqGMaGnAq9sbkSZDGPz2M
tewRkyAPy9SkLU0+PEO8Hq3EW3SI8lTslk+qkJhdM9FVAgNLGbCbK54l68QKJalt
YnulFW+NGUZvqZxrWk1L1H2Eco6ckpfC97zN9X5WYF6rf9GwLQEIVaBJud8DBC/6
//hZYFXvWNWxKF8i9AuTWVG1G8jS8mLF70cXQnujGXDUq8MKZWlV1AJsNrSob3tO
8u/S2+KOHylgkV1ItNHK5ZCdB4WLOAqXTPi5Hl7Qt4892C0dnxpgTctM/TqPm8kD
v/W+G1+S9jTMMQoJdckRIveSqkYCzPTmbncFzaJLBoZKtD8x0YmHs2WjN8BgRNRG
52z5DhgMYmzV98v2p6Nv1Nkbfmmro1AZVlnwuv6s9J0ygA2snN94MZ5N/zAmov0T
78Fq7ZYoBfltcAVKvFUqFuuV6gt0cXON5qP66XiRbnXBpv01ieMWakq3k+lI+AG/
Ql7JMguHKoXM5I6+oUXuhJXqoYB9Qeyw05zxb4pdvqkJ3zF4Quxxiss6Oklr7uVW
YOlORZg4HdMojJ2315nzVMgTKUuRe41WEu4sni3eX8SN8gn5PBdkuVFbgACsu6vI
ymnONBhEqcarDYWuR4nQIcQs0teWFHpcdMB7fHFMDmPENamGumOJJ8hiZBMpFzBr
+RTX1b06WUg8Ax8Vbk3Mf4QItTjLIfN3MYP9exrvb+DxylK4jSAnU4bzzlaMSt0P
OmKL5ALsxfnm85aihCQYeEomdj758T7yIDCc0K+d1r6NduU5P17ikdh3xwQSoRFm
dtVJAB5rkDOY+a8tnqmZCB9Ejgowk81Gn5nZUiQ9VSH3yGpEWEZsFHShcj3xkh7+
PM/iGPTPDXNOjdjLaD9+rXznwSqX0wMfeX5OS91H6G96YpSC5kyWX3YXKNmbIgkB
6H6HvAtK0/qE6HUlyhzyEnBWrh9n0zmCngBgx2ZehzbSaEjDEmtOGFdnGCIziryl
8T/nxkdI3fwyeTcB+7Da/1yY0YnQJllEbvD8nGddL36dPyEW8zGSd2kXZHvIMn/2
q0Wh8fX6sue6TxP16eFpQgPHg8uibKw/OILY8fv3d7LvNQWF7K16sCZLAYYWIzw2
XTBb8T3gq0JHzHto7lOpXP40Le9OhrBNTVgTfJPNzTJiuLDUNzR/vHjnIVIPlwMJ
DhDMSXPtRPz3q2w5HjKXklYj5PsP3hXRQJDmRBLhRlviCqxWWcDZwqLat/olmRx8
Wlhf4pBNND/M8HKjZ7mf7+5vaXDqtrdyOjT+4hQE4EN4pInkI9swQLpGqJ/mJFqc
2YjLjWNfa8BZGDbnMo6Vo1dY5c0zMHk6bt74BSCagpMzwGbAHstIkiw/tB+ESHzF
H4Mjp4UV0yBK3M6uMapKOod/+5Rj0yLmsKx5RbHZw/t+/RdQXgRfQT/7GjMfsAaG
Wx3ywU3k4qV0tN/ADTbtA2cFcWMb31GAPnnT6I36/SNP8njQ4H71cRDyMbOV+ISq
olH3AhwWJym8VFEElN6TSUEt287/5WbgDrbBHZi6xp/Y8wruU3wIs18NjZSO1TRq
qJM7Xdeq9tf4FqDNPLD32xYqb5t/tWBaoblWYwBdly70xv3lZ7Hq/BZ6RGZ3Z/Og
NGp5v4NPGGvXNvsaYPfklJJ8nHH4dhqFHI9Gc5lmL0Yfc4vWWIrZMspEwkFsQ72h
die3mbirUxz8gcfh6TY9/0N/W/66raEIyz1BL8ezXRyRJC5dldh4bPjWhW0RzG98
hivBV28z2rkP0AhguXuZm5TdzbabSnW75EA4aIWL6c+jeV+g/pzr4P7Oc0Io+iE5
Kk8eXH+1fEhWWpHD2MjyQ1BFdFaL+/c95ap8gweUPooaA4wz51Auf5JiseUUIqG3
tTiSKApDZVhtkFgsrfUzjcRzBdYmUtBXeWwKa5gHWaRF2cyU9aX5svBhDhHaV6D9
U6xDBkZrmHapdfr/rc/uyQgwytJHwvqxzX81xm++ygQOqlK/OIJ/GUzS0Dl+SQ3K
lDkUT5fIHCdXnLNTdthE7NMfz2xTSEVmKKruHlL0ly2Dt0DWB+AWMpLtQKj1ubpN
lMAcfxdF2fuyAfzmRZERuhSm+Odog1K61d16W92kAleeIfnlNrUIs61zI5Ulp1GE
30nJxxIH0HprGh8J+LrCcv3Y9pp/lNohW9oS9sc3NmlYqbx4zbjvReyltRHjYr7t
oZfmFo6noRaxiO8RMJ/MPuwfnoB8q46Bq4IJDX4cOPp5vsIaOrm7cgU47gd4ogqO
NPXUrB1Pm1NdAvGjqQiRfXasWNlojGLh/SwyM2v6vYn0xgZKYIBzSY4qUbHQdSYQ
SBb2QI40H78hX3fb76hl8k14NpkNiXHRhA0FQyW5EOH0a2LkP+ConyASQBuJ4t8J
gGaVZQTzHAj23qPtLW3cObigRanauK73sAHYV01X/cc3u13LZPIxIRROKfTjp50k
8QY7e8zi3xyDT6Rm2xpoNWS/rNLL/ESQk3dJStt7ErmHZzCa5C0I0nIc4uvCfIdX
VFqTel2dmaHbBxJN5aVR2O1YduNf6pQ7M2whptFGTcxH2fAjwwNti4g/zrilulqk
hgCPABdommSX1Nv9mIz95/MAwuY9fJU6xxtXyCVFFea4/Z0aT0Ez7WiubFhq6Fbl
xmE9NjF9x1YTPBJhlipA5aEa6Ob/pU5XAoC4maH6M4m+lYLQkQE4JjKrWuHeD+lI
IVaE8/rorYe/cB4yVSMJ5OI43FQih29CCSg1g2mglrftirHkJiinzKHxvuVUWK21
rJaBXh6iUZc+pMtzGw+5OGIozYvroR1EAnauGI9S1LjrfWTXh00QMbge+nfdaZ+N
1WwcZUVRkT04TKGvBMZcArmnSEEWpL70+fipbOA4B0IJkIbpfRzNeskWbakjjm3I
duAH1wPn+NruMK5hWGcBfbCpOhjP+QL1RbyAmjrQM4DM/hBImfIWVcI+kj+xU8UP
KgKRQjvA8AQe+w8HtFz7AF9YFVBlBwTlbU0KpFmKLxOxBqn3IkCdtBs3Lyl7L/H4
mAwA19oVtJl/IVYVjVTWHYtYoguWNnwK14hzjIyCMfQYaEmt5gwcFHsCn6EO+8X8
QHvUfbWg8rnQHepcfntrBhT7MpnC7K+DL9YEi/yn0DC5Uq0PTwyHoXuYjfCb/A9e
/SQGPx5blzo+1pM5FNMOUVwJZKocyTyZg74zPM12tdxuJb8nRcf3hVZIDpFtmWV3
WRhcpYLxVXqJILESX0UeBlowTE5veWDyq5JhIyoP+IN4OEWPswgJtfT41eTGX7z4
5bQGLTBACEWSYaO1T3o/Desm/E8Y1MwekXwcQbMfL4RJ6UZzzcEFDnFsHKHFiQzW
gE5MnN0vaRt8Oyb7KrJjctjErwqEI0V3CXHKiImxpJ/jLc/pg5CppTyfswsh7tD1
Cx5JHYI1zjHqgg3qazi2MEVLPnFlhQt2Nfcpo6EnIZbD3QYYdmbHezHCCxWNH+pW
I/lLkkA0bvWn8PMb6G+ZgjmEtS6F1Ew4Cq55u/vmkQmjt1Nl/5/I74MX0x+Ya3v4
zz/4CLujT31Wz+BSki1odmhNIOZ7c1gJFe4eI/YcFHo8SguZE2oxvHmalxz0fklh
pugfJesriblTntL2vFclYCJWOUHk5PS5dR3ar0gxN/QM1EuJ7z+eNWcL+ATcv3ZH
qvpAMP5b9JrSe21/jEd64TNThO+ZttYp6p3lix6reUcyqaj4y89XaYoEmTRUDAQQ
ahzY6gkoFFPX+KrsL3FDPZXt5RQcExXmrrQfYSocDhxGRaoUILjrNR6RAEwbjFMn
wSxYu3Nq8yiQukg2jdiN3I1mHmJTMQmUtUaIJdinKXH/USEO1YdG20TUK8inJ3jC
F5zeKFjXwiWEo8DKvjpIkzxeJIB1Pldq4GUqZd4JPjcPyE4swr5sfxMBgdzzyqwC
fHIhQ0Mh8dJkUPaHanqE2oyM6v73oGKFGNkykdYyKW0+OnKUVzlMQf2ra5ylGNjV
4svfY+79YK0hazX+ah09JaGkuE4wQCFtbyIzxYGMfagEPKMj5fIHWeJHgfEbPbGm
MMS5iuFm8RtPY8P8TMOzvHRMQb/KN3P4az4lxogpmqjoHIHsp+zS21Uab8Po2qxF
JweDeFaXazGGWll9RoMMimUOQj6m1eC4hESWRjMyMEywQxvjB7N0fSiNjOKV+ZIm
Vh/et48BG82puxHppOKkqm/36NQJJxNJRPvZVpllxA0xjJs6KB7VuWPZEfgi/fLW
kSZXF0sG87TEcsHUJgkKT3NtYSXM8ZC15kNQ2evUbCh7hgZtvU6Xwio+GIssCpLc
oRdvW0ufF8u6wbG2y0E3+d6D4G9d9kYa9YERZAwoU6J1oHi90bpmd1jBMDpMNP87
JQn4tycDPouHLM21ar94OOomi5YDXL0QZHAad+uf7RdvCO9K0aCG8VkNS8pdtBIJ
IKqZzfWAH8UDj5FedK2nen+lZtld0DNhOMlGQ40AMUvA2QPzaLznoUbkIi7L7RRd
iXVm5r8cMNWitph/ueXNSiDviSowVC7FK1SKdpC7eNmGm3DUn2MXTLjBQg74hqR5
4gwGmqUL1TrkOk7aR0Zbo+RFAqqYjwrvULYrhRwcyPbgfkrfO/a8X2bsGQZ/Qbo3
ldgK7tu6wktgMTVel92AqeFpMB66Iwgb35yuY3Co00cqnerMeb9mirNWkAAiSiF4
FIgLxkH7B/jl89uKpsh4u9SRETECa97i20XX96YBkWCkUXUXgjKw3bunGdBvpg40
pnosC7zV6aDc8swWbq47R0ZWqZFxMGekRDvXeoLVFB0O7ctE4JTXvPzf1WkOPOfQ
9gE7kk9FODGkrfFcY2k+qFYqPrSzgfo+cQ2QtKlnhUoPDDbM0gttMP7uS6P8MgIR
4MR5tU3EESlsZqd8cxcFdTOq61iEAp+F9XVKqYIcFF+Y2cyCNNlXt/WSMzVe8zu/
attivNp6ck1FT7lTwKFrudbL/FwSPK2vT2enFq52k+aySU/NqVMUV0Yx4u/uny1O
UWgfVclS15YOJ4ZcZSFogYgu+ZwJK0uMlHc/KX11+01Ds0nsWGcoUNeBSGlfdXMP
hZ0vsRx8InYuz9VDpocmbbQm+yWuZRLKZGA+g6F8xJ7vR7DpWeCkoWkaovlqT8Sb
75Bb5PlwnAljz74hIJXI00VQyLKXDOVZr/MppGYLV3mIsHcmL9EkMCSbzp1OUNKq
yx0Zdjf7L+LKIHgF9IW+TwIKmw3a5IhprH9Qr2u3tNV9oPSEVmKNQZWBIFOUyYeI
LIGo8BvCpOTdkft7mNDza7aFG9FaG34Qe83X6iNq9Q3lFwX1s5+punZQeUjhEPZm
ecxVcU3/TBX6bCoSzAJrFQ9SXGmkGVKLsdb6FDBi/o0EMiG1bNDnjh9t2uHsmwS/
um32Lmd+HFNCVmuCBK+CzNe6UoY0YMRKXbl2nBBdNDCBDS6Dc6kgoPyQaPWuhPlZ
F2bfyvfb2bsOpavgFtYpBfoPgb0ySKHWTbJVjVp6X7Z+D4KCmjoFfBoy/fCG5+yL
beQbt4wFYNTDFn3sA1329meFZZo5XPWNJU30i7QUL5LDML40nLkixASuwJ2ngcfj
ayVuMPHzLAl3PS8Q/wfx8UWMC1irSx6CkQlum839urfupZHBKuaO/fxCI/HD/FAu
MG/RmGHubuJPvl3AyLA4FYXFQs719HKNK4P1UQLULnk0BWgD54Zai7GDSo++6yzT
firmmb6T+pB2pdhsXQN2NmjeqkAY5W2oQjWSOtSsv2xhMhdo8ADN3+HF8G0FDpTm
7RUMylxwbN5IPDdR9DmoSGZzrBLksVX+jSMwwhunnYlruw8vgYJjqCACUqfAiZi0
y56DzaopQ20e4baWW+1+oLQ8N6fljtebv24kzPMfmMzVhyzXfeiZ9wtI03+/4ggN
EQdLFSqDy+TlE9WRgEwjURs4abNvXo5loBw4JKPeCqkmkL/Gi+RpEqrrSGDvEAai
23zXzcvo6xban3OxujPw+r5+F2KkVf4Y6NR3Xaj1TYCbMn3lnxQmhuLO9iJeYInc
lcw9GvGshPnSIFTW+M+HzxOfC+aABmev0SR0A1atzm4CXtAesIlEu1usfpXllpxm
YdQCytCRR07iynsLEcIW4CRFOeGNQn1x5yM6PcWm3UaMDF9qx1YktjiRGyBY+Rys
OcaZnFcd0czaFVKOvodZ+4LyKmApPep9oVxPVX9hioQrnYwxAGphwlTPwwCzcKBN
bwT+/3tuXItFLbKjVmNJYFPd7w6abXnACxtTmXC5R5KisVDp6f+3wJA+RvapjlVX
bHCV/W+NpVPNuwq/aecz9BTBJesZ+UXtKmI5tHF1z1U6u1CMaqSjUEWmgOMhyQT4
+Hi6MHsJ5hEmjN1EQGnAIz7K+3uK8yfrzBFPolabC3j0GWuJo10iYGG6BQVSlQp7
JPXXIZD/WRT/zjGxS1NN98IeQRbZt1/JYk++05UVsMbjBWw4V+CygR4hV6HYLjeZ
tWHsb+lRL30RXwc/Z/d182EsgxoF4/J28eRP/IBdfpY7GLVEhZO91WJAhK17jlZf
m/bhT5QwXB5L1QFhXd4lo08Dh01owdElHA/F2RD75FHoMu5BmeM7bt43o6Ay47dC
uyGpgR5EQBP4lCALEtrsgRDeLxbhKIJBEgxwzkCp+rV9hgBrcxV3ZrlE6PVsJalx
jtZuxsajvslUzwbRk0aNR4qCx6PUW8hfd3dkmU3BJ6otHTeLp1CDNWhJPXS7UtPe
TXctSeAdFyjZuaqYztCvz4+EgMe8BhbomfKqYIxzBGurn30Lq8jyFngVov21I/f9
tK1IFbWcL4sPkAOhYJ+Ss1PkjKPaqGwFeUuD1SDHnM+jiEy/IYX+YLxPxZr35VIz
EizSH2mPirEJe3iS2GmEKpbCWNEA4X/a1CUoC2aCtoyZnqGIdMfzA1S+sqqGa9ri
FXPXZSlY5iy8Ksk+j6kMTUU3n3fna2cpr2TcYLsF/UG+/uDH1E7qVZh6Y1GFv4vu
tI9ZuMNaMbHhx/v0pwaX5l3Duq/5F4A0Ig3NzoRBfXAvXiEHYR6DLhQp1l+QvQJ3
pe3iUE4WpueeoHYmAzJOLu7uw7rEVJB9rOtoN6LpNGGg7wmQNSpGuU3cGeFCd+cj
aMcKD+eqMni+jCOYTfEaMl2nbOgxRFqj4+dryQfE8orj9TWn+XuBmyU7wztmaISZ
ELKkRlrkd5ictYQ4HCSo41Oncog0CyUN8egf7emzdeI6P6jbTwv8y2EyyoQMXXwA
YZnAVZhB8e4DB9wCNEQ1s1p52bdklRk+RO5Yr1eEw0Ht/oGCzt8LhiFKMfIHlVSD
PqaJ9TVSYCmxRpFBm5J2U/+jQ4MuxYqHh5B9LFovlxTyYcIPM3Mi4aE1cKPRPvZO
3xaEhv6vQWasRG79EMFwf+0M90BPQ+5ZnrTgIXbBafTUkMLq1wnhwJjXIbLUAKPI
7chGXio/3iNdWeITuRuNfVDRRSzocQk33OH//hEHvpfc/mrqYl9lwiWsRLBjs8iv
+Cg/uhXU1GjiLu8HDA8G71GRIzmcsPW9o8qhS7rRMzSpewUQf17I1SbxXJXpvZbn
wI2b4qLPiMPscGVC5ASekUeb495wTqnGiWAFDUpiw4u6e6B83lGNjem5+0T5W1cN
52pEdo/dVj4LpPSzBZCDfuek3p23tG43PijtUvSuu/io3Y9BTSwnIL+An+viIsm4
td4F4Jy8EyUBkiNgHKo38JOlpQiyuuxH68MOWb+A42z1fwTkNGGoUgk/7GxlfKNj
6V3GKFpAvxxNpOxgyhem4p46udHLBPYlhllJk58OemC99lmIgkvEZJb/XIWBkFkn
TOcufxY0op/qDglWtFsOxTQ/qoiyGmLE5p/+OSW4Ietb4wweEp5o/t5g9E2Vxe5o
9Fp4Rx3gmGOAEyAAkQbdMTQFJi2+jaVGwemVN8g/WXHQYtFiJKKw9hG8/OjL0R8l
6+Bdx+TWgimFQRBBtEumTnVWCpeLlNWzhwIyVHErYUKQMVl8nmKNN+9Yvd8+ICPP
pp8DPQ6KdR1s7PeI6rnFx6RVGrlu0CMlTvh/vC5B95nAEVlkJv+i3tFtjtvaqtw8
0Iv891oZ2nQuZkLXDIi0DGyCrUAkWZYkHEz3+QyHbHPSSXhP5G5HiZ3vzpBp1pHu
B9U75QIdrRf+nVd2Ve6BMhO8w+Nkr2JqorkbVTVRD43j4w+U68CAjFoLVk5BCJYi
GemFe+asn+Fr7dCEjyPr5V/bC78vgoMK47BoV+jTg5FeE21Sqlh55hPeZ3Dm2+Jc
848Vhco5QAySdQkWf5hBPqXnSJ8Rc5KKkXRpjjKqsG3D9CiG8Yj2wWv6vuQJRGl2
UXoJATLJDGsvHAq6w0xACS8hvzXoFHmU2SUmD1Mw9uk/S0LbDmgobzE2A/3StXrf
OelWolicypUAN5Rk/5eNWa2+xe8BSExuZ+xN4UORFz7aEWT509MLS/kyTYsUk8we
ySd6bSjmDyDoBMPd7ouO8aYmnpVXCgIUCk0sGVU900w/Mo2dQ61n/pEdkhpl3iNh
xuwS3pWLYzq+sjfAwc6eR1srWPUVZkzum11ylBSOFVVOEUF4ct+5PrHAlwvswlmo
0p/ngXZLWg2s3LiXDbxi3rpfHfQr17JeMnyae8F2o9uywyU15YCn9yRR7pCnnK1N
7nPUDXHusA8WiZ7zOqBBpNjdgkNva6O4lXR85nSV5a1qWI2NZGVo0NNg0s+2xMFv
zXg/lHJwAuAced16XQE2wLqQ2tDyrW/DTxQE2UUXwduXFc9aEeTfgEAbYrtCFKam
gER6JLHR9c32smGTZJ9UqBoXCBNeNWgXj+Bb6ij5Vn/PR7fqD0x/Z1lD+/rS08lF
tNHvxsoOa8DFohgk5YdoIqSt/YsUzW9tV5VaSC2H2p4cSBIeBo4wiUm2EDoBzAM6
qqSUz3MoWg9NRPFctD7JWD+ESl0NNkuRcinU3xEpgGOYfYerlbjz9E3+3NxUbqTF
9DUSNsCwfLJHM/EhU0v7epL4fD5iDgaQDPQSYB7FFOh9JtmSt4JIAC3shFF11cv9
3Nvb2wj23v7l7EkeA/dPXe8MzgaNpqbvvccivD4RNDmBoggMWkJDJPHql4UfEt8x
PB+MJs1APxr3btfXFxHGC09atD2K4HWRk3CM80JqMaezboqJHvHyVrRqeKHxO/t5
HkAyEPFGZmofu+N/r7BVbtU4BK5N/9BfKtfaF3eFM+ODjKWr5SKZq/LKg05vb+fC
K1eZv2zhEKt5Wb7YcINI9iSQV/d457Wk7/2wreVlCyU4G2XDt96+7ximTxrhFS8Y
r6yi+uPs8S+RDiBPzNq6BQzL45l0+HncjmEwK2iexhady7JfGRIIa4pA3yfJ+2mq
DTLmzXrDVIQiULzTkffORDCgMwIit8K4Cnw1SDrfvcYDktJwC5nHOFwYugulO9uq
Wy4pUop4b3DHS9168voMuTsuXmenZxpjp7WRkKQ1LIuUHHOQ02yU4dPyOChPx00M
slO+d5GORGjlJrODqRxirTY+4troJ1tCKYAf/5P48BG2qKOJkQkIBOXa32anApN/
1Sg/pGd0W+B+GozBRc2tgwJVSACYj6hdA91vjzzQ2BocSq5u05ymPHWhe3pbsYGA
JtdwJbu4SVZCbrrflVlpTgCOOlNoYwzCGIY8e0tHGADCV8ZPreKVKunSQlUJi/Wx
zt7huFarYemeE+VblWBM7HE/OMYZ0mA0qRlYFw6bhiLgQyYYTrw99Jz3rti9KDM7
+/AugIkllb4tc1x82hlZtwLgce5WRYJaYBRAJP5oa9UhY+6P6IYFytDIawLcmj3D
0Vx+ztLiikHiTI1L7EmHxzWIa9I4KE7sfVcXshRkC4ntwtoflBE3D/65NTXsUiBJ
LPl+J/tHDWENDANrwlNZkJLgg+KrJJk2ZOQsKu6Y/bEaNy/Ck8LXbhbKKEWJch6I
ktZGpQcyyATtFV45WEB6bBTQrxS2OGPQwmq8piKpOS9AwhfWMWfW819uVl2SfIqx
YS3wNJQTLSQS/OUjSWaDTj9jSQ6ETcxWl1dS4rwxjLg/i2iBIffeyHcxS7PpVxMf
Vq2TwZ2nliY+c0p2jAp4gqWok/YVhELW1cmvImxJgqalYpXw2JJ36noQHppjFMgS
lCaosV3SdwWbn7RDQNb6lTrfVc+1WwV54pBOBmkwwlnFhOTwh/x0KHWsx2uTvEem
OZ7yNaOWNCEoHX62DOUGBkEGuIsFrG7KccKXejUdkLLY76HKVqSeT3WufJxe5iZY
Mh4CvXk7Firuxy4sQAkYJ1hlMshkGhrIiWQl0SGqUsIbdSHchEA6yUJWmXpXyn3w
N7N6+1qXuHhBdzWgl6uiI4ebufa9xPOs6nUfGOlTmhqW+xCeZGKDGN05x9TZIjuP
V4Si54qNGgXuqlZ1AqHoTrQkX+lPcNhcWq8xm5Z73fDORup7KTXyJc97ZmxJ6L6Z
vJX4aCT4MWNfBYsL63+B5gSi/VGgijTGX7ha+uId/MuMjiR7UcNc/rb/VdZEIzYr
qprVn82j6efgeq8ajDkUDc5qo68L7nYoXILttHtVCnzNjDR/PXRsyZgbM5tTQA+W
P2S4N+GG8S3AusN0TJw7Y/4GTBjezREttzEKHNW4naJf2gRh6TqA9HzrfW1Ntcco
0WzPYTECJUOdy+8sxyd2CJUavm+4L6bPHK/ckmRWSm7lFaouzHrMHRyahWvw+hzn
Smq+PTAwMIy46tJJStPLPKTlZFPDr3av/6+g/Ksz9hIhlcW4hV0M7AXXq8xcbzdG
6baMQNzX2SASTGOZ43HHHo7B/5Sf0LVoJ/eTeHtc2uPK3I/cxhOj36qsFNTtAbYY
hCpFfMopqbQpOGjzTba5g7xMptIAB4Aaj8BdiKJiq8n6sUb9yboCotIEWVLw4aA2
NDijE6aqz0KafWir2epgQxvEeFqwyGo5Qy8UwX1Tw5BUJeV9RhYGzYPeXu45JS/h
C2v6F6LMJy6cF+fIbRgK9ki8sdTpDpPbXALyHTVVHM3maOdKVzSz5G97K+NlGZeD
ZbffSpxTn3YkqPAr/3tEXa2dkc3NdQ8eVXoXORm5IZmJyK3zI3l/7e/hLwB/HSrZ
b0DZSFvV8dcRvfDpDjQj1RxE3CuvAaYtCD7ko7eKyksRgjgbbrfihdi6o0txvOz9
VXtVwc+Kb/3pd0MxpFIAudwgrgWSBI+iSjEENixlDuweXljAI57XPFkU7Y9cliBd
LFV9by9aI+aguFdacM7+UlMBSgDjJHD+Aanom+4f4cnyRZK6KRx60/B45dltst6X
VDMTePRkcvj4oIdPm+wR2xMAiv6JRTaQd3C/tismBaKi/aA3lX2NCwSg7RKdYbyA
jzjcDmMt1cnTWdQKu2b9yU0Qt5IJaAEIi5OfOOdYb+USrWdvA0M2YO3MbBmCgnBK
gcXK2df9wSzz4d9lkX84XUcOOgKsGflmam+RLtsWVArj7/voPAonmNKUw9izWg/y
kIyppJpdTskmDAOhNtfe2wvqsDDA5ANUutlYw9ctW5iLia4C00dVenNhI/klNfv7
EsBLz1oMM1HpiqFluFK7jQwwrcL4eS/mAvwQRM7esSWELesc5/WOcvnc7UJjd5A3
m2lOswxL7FlLU6XR5sPGK+koTF/w0IVXjpp8ylA3NtugmOcUrv5yWuiKXR7GvWus
XudoYT5WxWOuM970k/9rsFQp02H83qkDmWoyXkiDgin5ewWhpennaDmpjC7RRro+
X2yWwlOfA+3zGWtK0V4WeDJhaKW96xWTfvcaYSLGPlDtmY+NmB3vRhFPq2yQVd9m
K+r/ZtErxwm2qDmoj3TzhSEJyHYTdrg6E2RE9g6QiagHx3tr69x5h4Z0+EL8PeQn
AjMRkbi+JMJuUsw1Zk7Cl5EsVk5W97wv6nexbJeuaTAOwX2qvfnR6ijjYk6vsXak
WrAsvwV2bl8ej6nyJ0L/CLeKdcargLWBY/ns3Q4md0EoBLFICzshjdORDhDwjWNF
h/v3XCgFwjNhvACh0q3DzGzSQfVKKRUY4nGrx5JLzT1qe1aHXuLHqGYTbhBI15JT
G6Bv2NKOhOWoz8ppMg+hPTrOSbXPoe7YlYcjqSvZ1cOltM5O7HZaZjUdtk7GylH7
6y1Z7fVH15AuyejMtsYeiyUnGajkK2IJk09pQheF8ku8BDbERxsJLQqOm79iKmJ8
5/aG5zqzDn8M2H8JTpojgNpFH9LPGy0BBNxzW8gQFoieIORa920iH++eVh/JTtX8
6eti9gMyZqG4+9+BC9iNaiAodcGfkobUcJsM4SLl86IQIfXICB/wf6PuGuXB2Upk
HIq/uvHi4V0RTAHv5CvhqzQiG9ExwCYJJJJOuGbpLK6KsaTh5NvbFvVFLMb9Mk+g
bQbhVuJRGuQpc3+CP0PlosJWG8do6DCnuJy8o6oG3sqg4PSIoEQ6Fzy9Gv+iMMcu
RsJe5Q9jAhSI1IW2vq84KdUfIlmRfw7eZl+GJfaZ9lpH8vj9LoxtW4a2XdK+yKWp
smDJCUhk+2xbeVs6HyTxfwQa4roW6njWAJKmQEKO8T2+hG1kHoPYg0W9syLAXdJk
vcAwjvWbzmod0Qiaz+7pSDrRv++tbyhZVztp+oohwfD1zKpUKVTkJjkq8PWLLRbo
1Nx8Jyw5cJgKLxjPBOkljx6SBDJ2+mHcL/XFfL5lRNVUOpN+BOuxIkMU7nnZYxwK
6JniWVnm6okq/9Gmpno7Rtyf0uJJs3mZHhbVMQU5cT24ctzyqppuZJb3IJytmLOp
N2zbRWmdYmlk/L9FWcP90zFcOF3oMaIJgMpS1beYzJp6HhALIXU5A/88HHmcfh4K
DKJq7FCAvXPYwiol5Kmjd+MA+i3MxKa7fIAxUzSNuqQH4K1qAnX6xvTmK6y+3CGN
6F7oXjqfvB9eEMFdr5cmSFdH48z5niITgCSZpshIRdk94hg2QrxzJzjeA3w8tPhm
wgFVoHvRsUBt50MWBnQ4r9SdecJBfyCTjSrU9k8tWA3Y3XqhWeQK1/mrM93Ezb4L
FtBTmuX9+Xgu3629ngNvlRTm3lGArcuPLLhvOE1d+0Vs4mac0hfi/0yVUSWzVxcL
LuQu6uCTn6jzxibqR9l0zCrTIUEb8J/LJ6vGxUDAt9v1a7q9jGe19qjrO/b5g/Pc
k1yAsWvdu9uiCt1yTwda6RbvcZQ8ltb+lJ56WWOZN1cZZeaUgXwT7fexUVpA2gtF
2ux1QhZJcoBkPOu0qcjGJLZg2AfRxyZzv+abGKjwBM4gvR9+oGtOciHqt/AgKvp3
LW2OeB9PiEsZ8Z57o8vgwG3SONbWqJ+letL49LPisxia4hDv0i7y8PErGlNAd0yB
MUyNwKD1U4Lou4EeQ+ogHzRykDYd7r93ROInofae3bpC/We0va/35Ir0G+jKW9ec
ycuoWr2mlLiMXmtr62MPt3v8r4vEaPJAlt5QQSvdDxjaBPP5aSGM6WLcVRzLpQCn
FNQ80pMzqW4/YBwQJD3nRaUN08wc9lF18C0eSFaY3eM9HGW/GDpwhxIclsE46Vf8
ag+Bvv0PSzgQNjwAV9+WxhIfizTXtxA8YuXEIiXBwzk+gnxIblaX29gegsv3EuoG
uD3eymvA+vGsENmns2GhW6w7Unp/SK8/ARj+IHl6QsLya01dn3U0SZhr1A8JU4WW
8nWzuEqu5JszAGMjrmtVbD/y3IsqjUTwG/DCcsmkenTs1dxZHyzgxP6kldVwvlds
yMRYJQXzoVg10OSYSEfzBQZgWF4o++uZjgofLvERkH70ElcaVvMg2MiEawE9HRdg
/Eb8NKdzcbgabmfN/Ge7TwYNUQjGO5SM/65IRPlurd7GA+tYwfzOZib3AOdWU+zq
QChr6PNzCvecfrH535rSwzhxwooB5MkMA1A1urs7W5TyeqKoKq5LTZGrif3fkK6D
wdHiVvu23L+iQHq4J/RrvjIDO1di2owJF8TMRV8fNuW6LmMnkaPGXhQQyVQwbzpP
gz4b86r3BA3I/pJhRG5TkRqrftNbMcORSAAaTlPebuMVYBEuJ17xy0mYBOcYARPi
kh6c8zkr/S4tDk/AqJ3TWP+sKRY+MwKlV7P3f4anKe7md84TYQf8ewDX/TnTVTQU
WhM3VkFESSB8BIA2AGaz6MpCIoeEXBBDw4Nppv1pnEWCWWSag0iLGG5eAKS9Ydrc
xJFDcdmOOaYHl4lkfKbZ+XaRPxqJk6tIdtdSvbX0PfZf5CSrhbHkjI0RjCgvjkEV
Hh6SghssRUIXUJvctroG1Wp0+pvDUbQf7Q2KuhghY8xBPbXCRUw02nnQxidNDjPv
aAiz75dsD6zKPMhTUeUb/rfWWWWud6E5+7knALzD4Ff9nysiUwDruRAlcZoppRPC
kfHxIIwIAMwx3t3Y2Y4QvFe4zLB4tgfIfWqGFRSq1c2asaCCVw5tG4WN42gjVn/b
em+rUbDytF9TknDZDf/dWzVjfc4ZZuPI5fdubpaD6DOV+vM1O2Y/LdlYREUC3w46
JA8wZHmNvp5nE6T7x7fSoDfQwq/NL6+Ey3fixsqKmjo2pIo0o47XGmPpBuRGbO3g
62Y2NiVMtEl+DNvFVwORdOmYOl8p0hsJrn52oorUb90+e9bNj1kf+XKhhmcI2naR
NIVHAE3dASi5iC9gBHqWFaHgW5g8z+EJ6c7MFVDP9MgwZUcnIUYi2IR201gNyl2T
7Lf2fw7+udE056uJ+AqDUJ+bsCmBR+xCqBKtOEGzJ7AmqICBbZ0CzDJyVm9WmWve
m9Yuy6xCx9FnZ+DmxmaRojURYrq6gkLSydQlTBhW+raGsqv21tOx1HXxLvuaK9RV
X/hdrvpTOSSZtRFo/7LV1DKubkNHcgEi0SuAkGnZaikbDKgXJnj/WXK5fiUoi+qS
bU0v1cw6u8JxbrL0H++3+oIfF9TMWCXejQxzidozKg2fiAt0jfMyXXNxF8zdyIhh
szD8FgeezomIyxXykIy/jRKtYuU0teiNZLEF9aEMkIvN9IlII6jY+QR1/St5u12o
Mb3ngjYC9PJsVStK8vYatjSd/+ul9lTAGH0ZEyWFaKJOOBeQJzGg3WCgfBWt3sXv
o/kL9BWxNekqEARYBrJ1M6UD5sLNdYnSHobK3PtfLAZ7WUEizMJUAARDcFzw44TW
cqZR1Qp+jKLyk91Jy68vbkdZgqT899R/WY6d1X6Gyk6w5SmD9DSeo5qPPZFesJOh
imKt657ij9iPRXPFUR3ogBf6eB/WPr28UN8bId64AvD7JbKHn8qemRvypNDrWeq/
byHOuTGBrUSUgwkz58hGqnDkPgbzMh7CUllpl/y3NUNlnE/GWCjWaZp6glUgqpL9
Hwv7LdVHZc90dBqCiqvU0qyFKMDNK/Pcfwm/c0jf1HM8Avegj1DKw7mHLJk9NFN9
FVOXWl3GwJMhdBcsoX8/sq2IA3bUXJvGv1fE+3g0s83FIRrH6+slKuLwqvBrcjRa
9Diq4XhSlZExkGYhy6BtgxrhPU5MmoiK/XCQjqR8nEHFdzhwFZu7T8IY4Rw5/6P4
Ajh2OtAiTVFUBgjLh7sbOVEjrCtckBhX2DwaTSffzGvRE5EYGmGg6WsB7wOTJy2o
lbiBsB4uFnzo9WD4XgItQwaAEctTB3Ajm5fxw1eRev+HeFjSzIUqjNtBN7dD358h
nJ0U8N7L5GBMu5KsR1iNsnUv8BvQJgurKiYRQp9SvTrfDSG4j5HurUOZlY4KwzoQ
IiJ77KcEWrv4tvg58aCSHTdLXzdaHqu4+ZhgyyktG7f1iRlQyZbgMLSlW33it9s3
l+baUp5pdJJuZXaCgxigaL1BfOik6ZuDoWsAndTeYLDsjzdKkUtqTom3XgVIBkgQ
iY1aux+zXASAQb89qfQDhm22Dmzh2RkDIbbPJAyjiZj4Y5PfCVzBjfHGaGJD+Tt9
v3CciTxftgKkdqWbS9IzQt77OeGNBTU64aUYfuT/3qb7ayZHfpXia+ObFyh2CpmH
3JH/TzonvKmoJFDw3pVXwPIl3qCmOQEZx2qehQjTJK0El0DVEkZUfk4d3xeKc9AH
JeSPEMWmmi1HNQXlZYuYhxVbxB2hjL+9i80YjSXmVQmrl+oCycZA6+ap8Kad+Qch
hE/AKPg14WPBivkuzBgjTv+tmbB+JJaaMAT307ltGHboLYj4I8obdqUGb9yPo3ez
I1JmL6yQJgtRtgzbjJnIT8eTkt4NLBII/fJAKwFkFqAyTzdHxdsFX071rz1bzXD0
fJy/N/HMfEe8HpzLWRtUSHX3TG+WhEJhMa/tOo5CxZTlz71lu9GtE0TyhQBDqnLq
xhaWkonuVl465HLXSvElsyMhfGIuRGsXa112YmUMGypwnUKfu9Ak4z21UWz1k5SW
XF9ctcAi7WRKX8MekZIqVozsd1O/szP/V8pUFNulDyVnuzKxcZPYDf39N49fSKOw
JtR66ufpGSd48pDdZw5PO+PZSQZlXM/CUlQqalBcHIO7Z+DKREDZkB6rj3LUrtgO
sVptQ1nN8dX7XKLimfK0Tmot0yiIztjzAMI7YsbOhMyOlas44k7XzEH8WV83Zfgs
mCO+wo7/X6/bAgASmCnmnR07OTTGXhfzIvR/A4nC2CpBGfgvZ/pA2yN8jxjsQynA
mxKgI6r6xXfhgoHdddhoTGGkVTy4tVyMASUk2k97/SSII7B3TNLEFzGR6VVDkuCR
ouPC0Bc6XMXCtgYV1mmThv/czOWyPn9Y/nB3vnQi4CIUrIlqJXDdP29fn85KMsuA
c1MJezq0Mrmz5Isiuh3K9I0ZtFuUiwqyZtlC6HzEmlYIU9jBSsJIsvRS3LrnRiN2
yviKqHeNkNM2Yv2l2k8SePAsNXQ7s00y63J/NjgswPu+DqD1icC7fzmTWUVNe2/f
fmQu9oW/NyMpz3SCcA5ztzh86boF9gZB7EwT4IaHZXEP5U1lZE5fegYsCszMnjsZ
mLWSvF2ctEt3LKhcoQn/bY8C4zdQIpEEU/aqgqJ52Grvlj4otemFUfW1jiwzy4Op
2yjVicnkBkytTg2rZ82E5+AVbMOKt8BWUkESFCMVjlHN8YDIhZPfQw8UdtqzgQB2
+N3kqK9nGBx2vjRj8PP/ctfK/G0O04agBjZ/XMhd+eHbk0aSJKfAYC/7iVB5235W
LtEGTx2aQpf3v+qx+NLyMmXSUssptUoZYso5uE3YeKzJITV+pY7+QRCVrZW97K5V
lOqamrCk6L510P0ql59xcGt8nI7Nd4oXwPTyoXzfsp+86ez2z02O1OW4z1Wg8ZMh
zjt+t+CBxLUiYfN8BW+wuHaoBpJSOWdDnNafnPEZBBc23VItKJARVv850qvXLJGE
7XgHb7r76TpR1j1aPbbUcfU2hBTSZSO0PTu1pJs5HAblZqBGXmjEj8DMWWTtPsAN
4mvKta91N8V3pmpGC2YDnbvIs/VZFm3asKM7mg1230sNR2KHq5SKmN6lprtB3qi7
9KWfx9HedCaRlz4cvj/I1rTkeMuAy9Z4PrmzLXebtLlTT0jToGZca+NuQhgaQaVA
GZxiVlxQoaDI+MiVTFa6rzt6SWHiLuQcBvL3S0RCraKM9wFReyM6eOF0hcCIB92N
CpqEyhU1gPKn82bbv7tejl0/1kJ/bn4gzt8Mi5Wa+ZaqMmgbsKS+WwIlpIPcsGYM
O4iUTHWdrMAslJC07bVFjBMOpmjy/DMKyC3c07Ju8mHYzleTgfeXee8qZhUVucxo
4gOybc4F9WVxZGylJp2I923vKbYUql/rinEYNhx7fZxlNaqKR/3cio2k+aJbVeNp
gVx8CfznKvyl/Kpz50oBE3tohY0eS/zdBJ/EGMTN5a4jjC/6cWTPfXjGdPaT/kX/
ZA8W7jQDx1fTvt1tXJ4EqfTs8ZyQhi56jcD9GlJuPztPDYR2ygTNQoR041YfQ5rt
9It/2Bi7tRxrr4qsZne+HhwxCABiha1ramGlxnO7zldQ95MYHmZjS7u5xrWByvVc
RiLQHjaoOd3AUg3c8c2F0DdsDsdoFNZpMnDgEb9PMNoBNkpKHJeBHeLp2ZJc8hHx
z7IDVx/L+lHvut35VI/EU/leLf0QRT2bflVzOVqYk2s8xeu00kKTt5/b6KtBM3xU
rJ56189fB3uUqXR90BWm7HCaueyQowHGqLlYLurI9Yr4qBlSDpunXfcrkthtR3Gp
6WhFjh7L67COVODEgWYBAYgZjVY4qalqdoby6I1KEdW/N+eO1s1Sj+fsEVd0T/4u
r3hfwR7s9N7JtXpRYiSW99+A4UsWNgxA+Vgn1GcLqmuVUIWWHQFst3LeAn9l172r
c1FTPq1OZNdeT/+tkO2l2kyhHOWRcWcO1V1OnqSlIdw4ebZGV69pHjG90wcRpgD/
s2gCvgfhBp26IiKS1RusemfVRqtGKCHf8aRFzKtDSf1k8wvGhuxVBwV7h5QlCqHf
eIyrLEhqw50EpiGhVSaFj+ya2MTKKsh/3BoY6OUQURo/9WD4VM8Hg8zTGIJgGSHU
xANOemUp+7Sa2TdmAlW/Ga/gmQvCRCFFzVK8SC3/yRPhCGwiDsLJikn0sOJcvFko
2LnJ++K0eDBt2h//VmqZMwpdBaSXkNRLOPNZ8zV3GDwYEzuxJwjbFs/lFHTrb1E0
x0sogZDNoFQnICLjsj6PDPIqb+NkLt9LH6ZD09BpRFJRmrj4UAMSLPQ+lgsaGBdf
2J6YeJPUqzlpOXW7iBhJGMBn743nrb2eG7NbLAp4s79UYDoeZYnglNjQYDJFenVF
KBXSFeOzrppE8URtaiRXFTiy2WPmE08ksK5yaPHUQc3zilMUEkU5M1HCt6i342/I
G7bRb/5nFNGP3to4CBbfGuNkARZDiSkjKxMcxDU0maBpPvptch8qmxwJzlzf/Ah9
o+SQ2NS2ZMz0EyW6Ba9d7p/fiOJu0wDA7uf1pulTRpZ9zI60LNeGLf5gV7QXqZN+
7h7vNx4Q2CVhejEQDwzm6xSGgXV46+ojkjjK4RfAXGegrwLfwC8q+ueschgRfXbZ
n7+ZEGRDJyBE3mIT42gQ8dWFluT4WSeK9l/Jj8dJvAwVRvblkfE0DfaHN6pgEw2a
IKIm9AZxdb9GFyS6fgisK+WnOnwU39v76sfVjYqDFEyKrrBPHJlJgO+QKiM+Y8V/
qfWhqZzFaK0pFSaTNIUJ1Bd2Ay9xgwR3p91Hfm8BXR4BriXET/NrYLCHwe1lxucr
qpPZIZP6Masv606RWoMfKPGvtOojBvS791EVCo5IL9sj3w4F0gRLNd+w1EFfLlVx
ZRbjT+feaj3TleVXyXcUAY8T3cKi5cox5vtuQ+65AYwUGOoanPdboPjg5xr/MjCG
kL8A1QpO2ONqrzFm9kx/nABRYD42IIJsoN56m+Hep5V2qiV6s5tjT96sqiYmtCMl
q6H0pbuAAXG09hoR6xEKfJNcepDJKjgwEOq3RRha1lx6SI7rp9GRN5+B5glFcCnU
dzSbml5KriN92BvcKH+3dlvTcIb6oVTnpTDIpuKkfBSEdRXatEQc9xDrRwHAOEHs
YdBXT5QUTIhPpqp9C3ayB4DiPnXFv8jdZ7QRa8fhchcc3pmCm4j5Hyc9RDL02DOX
JyprW/fmYPeOSl0v8m0zhUqKJL0wI3NOizb+x3+Hviepx1b4y1KGt1IrgNwW0mjv
OfX+JGC4BaTI4MtbqfS/aRT380jTgOEsK1DnYvGeMAMP8/ZSNvef0V5++CMaUDRr
BeqJDMVOtdM0cnd2AbKHYVmQlTBWMnATLwa8T2oiWIq3GnMk+6vjMBQ37dnJXNGr
S7E9yDUsiDCECt7Gwm7OU+jBA8dQsZztCvPjTLF/PB2dncp3vSrLlP/7F4J0RY/I
3wY2MG2qtocvrgSk0u7X0vxQsDdMQQo4OrtSXUvbNaxwA+5x5SU2RKwL7/Lx5r3s
/oeY5b6Dha5Q+JKW6gGTklPSz926+L5K/jJJI0MJZcT4LB4t1eRqgGRS3QuS9Zfj
1ZM4KgDy3H8YLpSDzSFw/kfDqWX8YXrTRHJH58KW4r1BODCt2kLmY9/9oP6YDdvq
8xgPJ2Re9UkjgwwhI0dRvTgqd6kYzrobfzq77NVuDiIzRLvrzylgBxi+dF3Q6jwU
9Z82UyAi4xPVZ/WfTW9YaAjMpuMJlqO1eR4WfJXn1tYHpA84MihPVr1m5ZXmu6FJ
6ag9ph4BdsN6xhZNM+EEF8AChZGw2jF54y/BOKJ2dPJcRGt8BKYSr70gRqYBQTfQ
o+rb/dSeMMwn6Z9aRFVmDuDnQeaTOxgShht/KtkgPNLkNFtA/GQNoKHEFVg+EAlq
C11osKpR+3QfQkfx5QD3EF2mRIWT45mm7l8ux0BWnC9W51hH2+D4UqGJamM2la29
H+8pOTWj12zNHoQQUeqFV82KvfBRcY3lRLupgiucodkAow/q6qdRJVxHKpGv55QV
OLhGNCAGgfMwYE1t2oSd3xts/BFVWQa6yiONcnmVPI52ymP6tMLC/08kDHInsxHP
6Nm9HfSmstE2Th6RhBtJnvSHWn/mg+tKdcP1MbbzPVOq2mqJ+IHWeTGs+NFZcqlx
ERQpXM7GJ9wEoUwg1wdr6Ex3yZvMadRH26DBCa4TLMY/oVuAEK0JigYimiV2JxVq
qkYdq9OzsLjYwuawd7CT7omSblFrvB/oW1SC2mvOJarfIg7w8OI9iM9/iYW60QnZ
N92HlkGK7icqyOXU7wMx0yPIwnmBx+UUOgo9nSNUW+fNHP41YsTcmA2ddAy4MtHc
W1bormbs4qKHArmY3BbkpxwGC9ij85T1d6FhSivopSoeXgUqlcePGK/69K6SzkPn
9vyJArf+3a+RotMrVYaXGAqwnDP3m5dMfh/NXKoUPMOTsVgzkNIN9dpY9qIHCSEw
3f/Cqt+2HygQpFGJjfGn34KCpyKx3tzbakBZc7Zl10QmiqlyPD0egrOpS3XLJUrm
0EBv9yN8tqQUe+6q5CgVK8MLII+iMQw9GISogz2mrkrG9aoB7VXPvKyNDV1ykwiQ
gyMqScQRmTujCYeZfnp1TOcFeQFZ2zncJII3qmUSoiwsISvCkaKa5ale6d6sMjgl
4trtqatOGSLqNnNT0l4XtQbRj5rfdbfzA5M6rvkssb7c6NHAw7CBZGWS9xdamUWS
Tb09HnMApooOLisf1Mh7KSdy6vOinDzwuPrtnFcm6xpUWzDi5sjn7quBQ6LlThJi
lzFOJ6yzhtgs6YgDBOHNcoDJu133ao4WWrGAdobnaPumk5kWlHd1GrmVNQyVUQSV
ShhtdzCWB3g7Ugjs5y3RO4iFe0Pv8RnkovBKThhgISv8WvHmD5nXJWPb3SuhqUNJ
uf8mxG7pTXg2inzkUGO3Ornj6+YQM5Rl5JLlLTADFpZZp58zyjl42Ln1lUEtl45L
nqY9IgRMWk1C18IRQw7hCx01VCSvTYy4vo+RtPt9MmV4+UJj04gruRJ7VjvIvmPu
2WP8LFug6Ms8f3k7+vnoIupBI2GtcbY/QCaSGBjQxoGIdrt0C0dPgWaBeYAcIWGw
V2qdLBDPOABYvSfjCBQlOcvTvyuJqL+H1tUKun6ZKtZmqxwg5oflONrOhe1yXjED
q/DKUioLWhEMm6v9KFGu0gdyjOVv7cJwb07O45HNpLbGr1JX0Xj8QhK9jOqnBDgJ
Yz/peKa6I8FAAh8L+QKFQ5lVqh2E8nFqV6P6K58E0/Yp5ao6WznM/jHMEfkRsG+c
r3mA9UtApmzPiafbIw6kfloIWs/O3BfseoMTkUbsl7wO34+vOJgC/jnU6Z+/vk4y
IlfzVlHfEDFLEMJ9TyvcnFnV1lBE+cRWqxXWGx7PBj1C/o4kxDuraxqTnUEoNG2g
CizO15SYls/r0/WdNKefKrx/AUJd+meALBAllZXUiu8EEOdVte8FN4CgyIUSiSx5
QUd2qq+WjaaYLIh0yiVCvW2eH2v0cORsiUiQnKqjtGfpomIjDumKVz6qEqKm7NVy
h28OURr3BZ/Hdt9i6pc6+FRcCBnfdckXN2+JREr6+arFoSdEcUnzT8gQNptoQPBx
q7tTguwBND0xd8/A3Cbwu6dy7+ajFczmVPMg+hKQ3nT2Zxg+/pH0U8zuj7yOUbuT
2iN2KeK8WW7U9oZIpmqPrlY5cSvH6yKhXUX3C9PeKC/Mc6tSHnIp76sEdAqTBcB4
j9oV7n2nOoL4exVXh1WJBdwaTGH+7szJrobWDSrCvLfRFz7VYeewSHRwrtSgEv/F
NTV2NXu/GtIsJlMsphKbS3Nb8cZiGZ6tpAyCBKXrfVsPI1RO0DaDJ00sRXiukMAU
xoLlJOxt8mprXibMuy4BZxFLXT27R4nmbUkyOHyeUE4F9wa97BvNsAyWcnE6WuV+
LB+y4iGycRmfOBsv4CVg1jm6UWUeesmBGszbdFAzVKgAW94WgUwhySUyR1VVu8QG
V4UpUS5N4iyHF5W5yzDs6M5tX4eoV34bcpYOwBts72+MBxW8tGdzlhSj/VsGiHy1
kiVWD4C791+OhO019OcepPZUpnWjhUykZZZ1Uqp7EEwKJ/T/dmC+2ebv+aYN0p5s
QsAaZabfnoV+t8bvkIDQMmv5cMbXsFDKBTp2nAb3wddkbvCBApiMuohlN+r4mioT
IDXyoWBvuAYuhVZO/BCMf82Zue1Wo7Q1ioa11gO8lza7R3WTZVDsza64CBE6FCo/
XC24QexVAVC1LzhaZ4gWgM8W3fAvkoER56T6OfGU7HFin63mRdfsk6T9maD25fIr
oznejgu4Yos/1BwrQbE4AcSvciJSmEbiLVwuD1tFkreG+9YTUs6fu5cN3MnNx5eo
oYeXMkPk2foJ5Y4wxS3jbDLMxAfMQE3yHQc3B/dIBZat1cSpAB/a4cOrpUKUqTj8
pENhyq4wgMV6oy5IinZCh29KaYsAbHl6LQzgZUhpPChETMxAi2NIl049tw6z071F
JqFM3sz/jKRS8U08yB3MlMmjfUtzV99UR8czXaF2LCML815IIpfroegsJ8k++s0d
5fhsqf2267pDNAlKIw7u9UMgfuwTGgUav5JfXaN8xPtM3P7oMPfwZPcnE93YtiW6
aD3L6vLPwEtZu24DioEE0NbC48AJAFROFmS1wZJm919R0CP49REQ7+tPoYQsXTSh
Vf/ubcHNwfpyY3DbaIeVJWdI3pdjRdUzkvUHHiYy/MLLhm3zpdwpLx/DR21fAnX8
`protect END_PROTECTED
