`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a7kjguxmVByDga+wk4n3fM+Xt7RxI/8NDMn3gykZTkBLUs8LpUPjthXNgkncLeW+
25U6PSgPLsYpUqNV2qpTq8B3WuwrnOnt4cNwrei1kIbsPhM5ocgpdIuBLReHMPtt
QRDOtNZBDRBgrRDc5jz0d9XqCJfco+RbCX7O8ehKBY8PrdFguGMqlVynvFc4scQe
Q9yA5VbazKZeMqxpI/5x2iBl6YQ3LdtMHVK78se7w9/8N9eCKoxTRr4HXw/2cLtP
NHQmcWYzT6uaFZCxb4JN0o/Zig6QtCDtcSOKXCD3fwFnLXMEPF7AqskxpQAnLYq/
/LGJ+VyXcxGl646oJ9lGDXXTth902A1akd9fIOcOsAa5rbppaiNsZ+yaa5ENt8+J
e+2kDXWRpU8GE0t6w2R3O8OmUzsq+mH75Nt3ZUSLuTd3vroF3N0keOpRrF7v9vFG
qnOpOjHd1uNwyoFWpDoUNQCgBlH7hPr7g9UHEo2vn/AvEKQp5ZjA0e9DvJptEch7
T7axAIEhH/2lgd0t/AJgn8/KkuVzX2S++/OC8ej2mcIu51XBhE1K1GXzxelSU1S2
IuYgw0hNGPa63G/db0Pm8xO6sO6Pu3gC/LIrV6tAB3pbC2ULOpuasVOtRuzaOA/u
`protect END_PROTECTED
