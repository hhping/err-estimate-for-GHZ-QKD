`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rMRrRby1icRZus+S5aldzJK+YwS2kFFNOpHMT9R4GPZupbeCpzA6eWTS6s2FRDu
gr2vydO0yGFOpODGmVoEeBzugMGeS51+cB4Kc29+2ZOjEaY4S8sG3YrmmSyyK933
LYnoC9T8TXl3eaoOI6VVPEEIjmmLtE4XxCCuOLHDPEtaQt6phRcDTQ1aFR6KVG/b
ZKFHJHFzKnTsfPgKkUSHH4qhjyU4QkJPM5KHdzoeakVYgOcrlLTzrJyhMV5mZQVK
A1skIPEfBEw8KnmhXCA4XQGNQ49oC3dWvWomOtSxbs5uuVVODcyUVNSo9TVjtU+P
AdPsdLl2vdzrfsuHIKVD07Y1e0M6QYqPlZ5KCnHwI2kiuz8Q0vrMTTkob/dUUkPH
A9nx7vv7qnis682LmhfEkOr5Aim/HFV6te+fQnorKa9d4BtDlBnr21osIuZkwrtd
tkwCh+W3qoJtdNzi/7sY10Di8Ag5Xa+mystxmX0dN2W+ymjHhoDofpkTuq7d7tdr
DUJGdvdzUSsFOp9w+sQlm5cQItx6VMnAK2GepDL4BMuq/evOpqek/sOXgMSCDF7u
`protect END_PROTECTED
