`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BN9QQIfo4ANz8EXW6hKHNKkNk1cPv5FQQ53H3CxmgOixc7vGXPx68TqOCBxponP9
ALC0GQUciAToD+i/Z45CzthMg7VCRGMXaiAdwmZ2HXktwIj3MtG2egTinSpkm/fm
XUyYQ3H7nlo86OkMm1Qiuuh3zImgelpVHGRYUeiR0/Rnbfj0J/V6dhLifgb32qoY
kUMHhnQ2XIybWDf61XvbJ8vz1LFpkPzmZNoXXZ4BfsLWOiIPQo3F9pKiigH0lnhe
P6Kro/0iZYsKoyML8ZRDjHBYKc1qEQYXP36HQMjZChq0UtnrQpn4qIcvUJBDHrp7
5D8o5pVe3aKfhxn/jxEJ8ADL3pE9LW0HH3b95C5mZBYfUjZCB1qEWqghwRBjpfr2
aC3QDT8s19LxYN8VFOMN+AOIyHJGyF0qWj+qUJ7zOHjPSzUtfOzEp54/CCRGyBfK
Pf6FbCwrtzXsXFQmZBxEo4ByEtmcDzn7TnrO15W+0JMDKAka2ZJAOtiPJbICEyYH
1m/x4b4GP7LGmCuVEqj6qpmBhmSJUITIH9laCFyAOL91K5vuALpEocrV3H0j9xCv
6+O9ePLogDqpBik3kO3Pv9cKdme/pPa2jqDVp5j/Y8z+phSA5NMoRwdYeXMpbU1b
+J+7GfkqsSGi7bkII1N6YXc0+IGD/AGMxLe+BWxQ83yokdd30HEgYnK1TwZIjp+2
Suoxq0O9j5bfZKbkUpBEJtZgFwzbL+dWmirSZ3M6Zow=
`protect END_PROTECTED
