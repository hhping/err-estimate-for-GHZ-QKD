`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOGhYZv3HUrLPzzioM09t3yccy0eo+WeaNuVGcULbEQM/F4wtBLDRXreWUc9c8yH
Lq/6PewFMOgRljj2d5wzR8ndigXsflwRgDkYnok9NUAcNCXcHhW3UkDE1r9rEr6B
IPSBdji+qDW2X2mRWm5kyGfwwyxKMbJDjPy+RpuC1X/tJs9pz7Y5niC7RpHU6dOt
BONmKWSTRlhMPJr34G0A7K4k4AM9KUS0VqSex/e3lX/TK6Npj1mdHb6SAhNebEC1
a7xsrEaEKybaITf1zOYFJbmFL3uq0JXWCSG0jJLP3Dc9gU0MZQXbL3Pc2gBI09IX
q7XqVB1a4Bl7fSXmOjr67kC8t9N7zws19qoK4AxD7y54cMdvmCMjtG0iLGrl2/cy
RX2qSch3Zngr+hEduFfNpRpSsLPLN2qt9x4A1U9qlNU+LxAive4+fEXd85kiNOuP
g79LGDKbaGU4PJiwIdvN1l5xJWBJUeZ5VlBmPNNp858RHjWUlklSMQrgNh3JXLql
wH62YSe0xl4K1DMuiY4GHmE28O29PZdFRH4Rr2U9Y9EdbpiArxFf38XGckKvoclT
lWdUS5y05pm+9IS7P2ycfC7TY7tejhsey5CV7KyNtQXbaTRzmiGRcTdrXou/QAh0
CB2QI0xMxgtQF+WL7NtaeSVkd/zwfEAu/5OjaPq/8ndpsXLW33H4BaXhG+5JLRuE
+sgXS4H5DCe7UKEiIUxqxhZGHgxuGZecqh6McDgDuRoLxzDlALxb88y5n4HkUa5G
bb0pLbtWe7J0CpKev67sJZSfv4CynCXUVwtYkxJ6CMM1aNVF3mmMl4+Mbmk61zpb
wRzC49rqcztmMsvbCUQ0HcJaej81fviWr/e3IBCgYk8+01BT3gkRQsj80N7J1IRv
gi96sy8FWOY657sBmz5KggQLGN54p8YEuYTxeiJxAVbFf6vhfAS1gTMiS94aYelE
rSJ1wGu2p/8qxCwsN2UM4qjDVzENX4n5Yj5hjbWa0O6LC8kVsu3LIzxzto/p/+mW
QaFeMTm/WHlRV7pdVu3zqU2BXASLAZtxV1wwMTBJFJuSFXUHeIfFOWx+sAzYsMR1
Tnp3W4vXI0fAm0LRZH3+VqL2dLcC3qN9ihhCcXaW9RN6zAl+lRGA/v8Pygd1/k1k
OGrjQh3RGxVxnPVRUhlzd5iI09NTQlVMJOmZrXkQam8ru+agiwobUHGWGRvlXHuW
nJF74xHXSElTJdu3BPMkYAhRD56/bd1xlDT4lASxVGE/uC0Cxlel3N9PkfQRyNgz
RYLCvvFhUTDKBHZ/81NXUEvDGHBJPqJcn1sxqvFSPJA3XiteFThENjiq/66cwy/Y
rS1HBRfK77GokWXpXs9Zre1Aug2cyudqHSXcMayv9ZdySvhsIZzdDBhut0NPCVX/
JyXp9Iwj64glK3qCy2e11sUoKyoTRTDIvR0i25ZCemzeIKopyz57RCeF1Fq3cCLx
QFiqd5UUuJPfEWo4w6fMtLSSI2cTK+emWawkUiVT8R/OfWuRmM46wzuDtBbmC9C2
XhsastSIo1LdmHQGURuWzkrvcaeA8CZzzyWW1tmpfY2Oq2tAfHA538C3T5B2N5Tz
lDp+ZPA4wZWaM55waRwUAt/+ijNcHtpDLnUF2XvJUc4SBucXY3e8ZcUmr5DaGtYE
tqbwli+Syt8IYoJeRgCfIbaF4NZMU+73yGLH07xMhhynDVX8cCqRXC1XDktouM5m
THAjnJc/j6WShtbIXxDEak9p9B/GprQsiI3grFVfWxiTM7zgRm7UCSCc1WKWEBgq
jgFZCAQfy5sTg2Xb1hq1DOPPDJ3DUW+1wfxQwxGuu/EsP5bA5rdvHDaDYZsu1sht
Xw7Oe1l6r6szgASNul8bQcHWeDJS8pc27MgMWhkw/VAW3UNOlElavPAA2w+m+MpD
KbacrdG2Wg5WS5H0CNeTOpVmtOEL6TFLL08dw7/UJBxlYLzpHaxDb2k+ntr1kwSQ
O0ugAt5+UzJWOXHS75ci2FamnIMW2gm2SoCWoQCUi1LCsO1/d/duE81znJwuPfNW
clVL5hljsYUymidM7codAdb5U5RF1aLtfKnU/mFnnBaQa1dDZkgrIfpJ18FGwbGu
yQbTYCjDXG2kcypqTMuwGwZXXsMj605w+2dIfT4qMQ5xrSLFw8Xj1Oc1nhGYzWIE
JdAWe3FNDZeAE9x58kPPdHKORReRYhQuaMhedChfUdGEvqvrxOCxutZrZUPMDvVV
B5beXAlnRsZdcG5mkaASCc6vpPLHAPTbAs9B2N42N03WQX7QShKMUcrVAnv6y0kd
BjR0HJrNmH8O9b+jIWdnZzrgrumfDRAtRRtqnDhpgwisnTS7UMQ3D0RoHKLHBhfN
eY6RQHo/gIeQhhr9psepN3b/FUGjmXSjd42n4U34YFSKRNX9w+TkvDCPBha65dxn
/rYWB+rvH9SwhBstlauk41+nJzl2sGP8EY/ExpT8V0DGWHyzmfUz3cNM47CwnQ14
tEV/sm65H2xeM0KBHQofKj98A2/7WsfASxS/LQiM37eiZLvj1MMdf3XsUBoCo44t
WDxr+cqGpuPzt5bpA1clatCuu4E0Q42k+Vs4NyPIa5H/CrJVlSJJb6tuZrYEMUAh
R9Ohic1Frszy7XNxshci1+EahVQsWQEgsPEWQCNsyuJpBaBZJxN9GyZQTt59Qn8i
N/DzAC2CAeJcc0XBMmrn8A1WBpvok2ZG3e2m/U36+Xya3jA9zDeZa7gE3/6fvRYH
6l5SzOgKTF/Cj1CLu0F06NTgGxxkGMtmKPcRdkZqezYdaFMpqhopi+UX68IbOW6W
hUCQG95Pz3sUnpBhyy1Aqa581Ui53WKqGRAr80yJjQ6ujGHf4MDWtGY2G6exX67H
RhyKaw88xwv5o4Onbg7NLbNfODE6ykjuGj3knZs3itYCG+QkKulO7jwVeY9L26ZT
T/LGs3J9QFNpur3ZHrt82UbHxkpbxRptY1ap0D7j/+46Sj8iTATXuAgyAAV1roKk
BX5OOB/fN6ZMABp65LcgsBG6aVhVg9NRE7HAHfcivSUr8YbOjBCWbIEU+e2mdKUz
Swo6meX68HqyIgJFWclUDYIdzAamexb5hB7UtVD5QBpBkK+K5lZdHXvqeepsXApu
qlIQ5e29sCiEO0VbEMy5KOGO1gdXCNFtyfmes77iVIUp297Yjzk0IbckGJ2SzrvV
viLAvKdMJzQXbRgKHNiXaHjLm2oX1TkuRFCRh+72J3EGKAsvjH1/gH1AT36yFoZw
kxsxIIS641SDT3COrvE0MNX9PC6SLN3IdPmYfm+LYxuT7+66+z022OYcXT6/Y4S1
RDGqifSC1w89eC6I+olBsLe44hPpTIYVcKg+i+7P8XFNfrHdKKuDT9zA/MvrqMve
gJ+FSbsY7nchi5xnyGaV1Hy6SNOHbWl7eHnqiF46Rf47lM8dlki2jKseodeIevmr
BixDRk/dkNhocQIdmtrU4WOnvJugyIm7bBvhka+S7NUa+y/QgQRJqqDUSLaO5d4I
yhKrpvS2fWQL8OFpupVOedWeLqQGkgWmxF+iR1ZT4AKaVS9rJL5mYxkq6I1ar+ew
qr4Q+JrnGc8uRUcfmmsCyzq4vlKWoxMB1RSi7dVs9QvpaJaXvC774i06nstEbfou
YWVMPLZWfALH95pd88D0gnq8QcHlDRV8oQgCtMKS3Q6G9KBXC9vGuoUt82Sr9Txr
Bx5lv28cCDO9q4dnu7wNX7EjErxmVvGlONHGfmgNwbWaiI/ahKSzZ7i3cd+NWZ2Z
zpYoWtOgLhI+f/ysqzlIh9KHb6ZB4oaWTnQrYeW9akVyTec8+MVlvVX76ei5YB1P
RUCeHOHJYVAtrLFXngtT4p3+deQ5jrw+QO95XTSOw9Jq1QqlbvbfsHjphq5ykt1w
3iV0BWrtpqHFRiopeFLXZ0muXafUoVER2hr8O3SNOK4Jir3XUKkYmjT7UhWmrw20
nqPFEqt8dB6FduTGVINW8YkbbkRbxMnkl6NY4d1hXuYpyPvi6NQ5SiQYnFP0mMDa
OuQNyXXQTsdG7PxOIbuSJK8OQaJ/p8KPA3cP3OY/jgZgqSZywRyRQiqjr+OWUZzh
i8TV11VUevBigb0dKDW9deTGWssvRSrTRdSrxA85xh0wqizC/YgNuXeYNoFFBN9Y
b68Fe3xlLZqEk5nCwHsvL78sOiokwwjrgAZDc3IqGyjkSHRfehwK2KVlllQQT/d3
pqTJsXePSH3pPTj2lrCsu62Wd6LrrT5GXDIl84tDXVKcCCQkZeET8Ri11yk95fVn
2SlUv7XmPte4oDFXEtL8Yt1sSkpTT4jtzMElCmdbxLywJmub7KbFFONUarFadsiL
J2sYh7HJiy4WvQnb4zEc8fs1AQ6CW90jsGLwXqHbzPg76AeGooePzyHmViyiGlu4
wa/IPe8qVLx4zydm0tXnLr4ZdUqT24yr0WRfYCrxGQjGUyPs5wQ6+Vg03xLhBisc
zCyDY5c40uawhODVlPgqYk3DIr8UKo0e67E7ognik6nUikuiQQYbY70beTCAOtXu
j6WMxkimc99vd8IdS0YiTFrtsKvh+7LF6bxUjDtfk69+HOeD1YqtM5U+w54OCX5X
m5LThw9N30ByCgzpCgNXl1N/E4GFetjiZyjKri1yCEkCVSI15T0w5jV9f0ZervDI
q0SSvWX6htop4k+m1DYNJqycYiJw4L7LChi9yNnHMtC+F2JjC2EhShz++n/3b1Cr
PdmbSIF8hD61cPVESGHQKce1WDqN0vUdowCI/K2QtZV7iEHDcNPk0/IEGsVBHm15
8Ds3+qUOxVeLeQNT/P9Uv8BOrRb8yAT96wfZvnceKtHR0N6moJNxz6UKeGYfSFEn
7Q8ANmddj6+KiH54BZTBRRo6b0XpDqTdsFuwzn2MWRpV8ySJx8shwgKQX213ITb3
MgR37HOah8ldQcIUID1FSPeea1WQu1odjPPbYLg4KkKSOrRGKeokff2n1o4K3Tk2
CxsLAYi0caJiU76woFBpR2tz77GItYGcUCI4JwneVqHslfCmEvOkjhNB6e2OanMM
HiaQNAq8gx9cVsrxdg5fIiXbiDJKxfPIhc7aeO0uJIj/bEuMqoY84J1tHBKoyRWm
8PdPjJ9VWnjrVL9PPJ6hDxgIA6KE1WpW55/MNq2NmFNSdX+3Di9L2ihpyxo/DHyx
TlbdTq9oGxoe+k9n05nQ8ve3HVHGjcFTKoAeEwRNHHLWTqCc5STcbPgIABf2V1xt
mf5IZf2ZX1/+ERfwyJjxkz4D5jRAZVFd9NeCMGH62H90s5euelQVziUzXRjwWinl
NqiOr/ONtPxxDdxV3OFBQNctvl+YHPH+VuO8o7jgpeGwm2nY0HUUcFHNqZYStnkd
SgywT9KeH+4VGvKBzDTGyswcdlt1kOBb+yPlv7+SaiC+TZ9p/RNZMmQWjGF5UsQJ
Yk1NhldPTUFSnZVyS0YI1BqNZuweuvdOJSbtOPix5YwW920l//8+RCqIL8uUFhok
OuHyNXYATWj6/eofGEmWZA==
`protect END_PROTECTED
