`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aizq4nsx1WipRG5IQICtAFRp+KQohvQr6VUdguZjmNEdrdy4hXM24KeBCXfjjxBf
IAGgEyZtkMCC2nCO3ZkeyQsQ6EjrjDG9nF6Ja2Q38lOqjjIXfYhN8tAvSU+qd+hF
uo5dCRP1yBgwT3nExipZ8jS/LKIbD7oaqmuvt2j2zanM8U8gAaraFCvxCx6bzH+x
HRzpuJ2uGuyfQi3z04upBSyLnTX1sDp6KHw9HBwoc+FdFyKULd37KeJNeio8rvbT
gqnrDvyEmE2/sO4rxTPdAeSPGow9U+5lrGJYsVB1gxLuZ7UAkq09k58aEWqoCPaP
9iLNoCtKC7P2YhS85PuEOaqyXJRKKsOsTxH4k1YZy4k6w6nAVpWTTUNg9GhnMrNV
BML7zwrJCzCA1fBabUYyuG+cE2UWz585nDMneS5bsRA5KuYxcZbSMvT54Fe2YuUf
TcK/WYlQOrQmZVUbx6Eh14vts084tBnaZypC/w+8iE4yxS1sHJerInHQz9MNq1Qc
F3Cx4ln/A3rwy+SpovSsPjb1GZg4lquVL2MFV/1gi9wIbBSZvbLyEuDHjTHyfYV+
O3BV+76y5PMLTrJHl9G5XgNFL41CJhGvdU87nio9H7ZSpshjdM1OmwuvXyGVfdiB
szyD9iEyTMgyU39gXdTg5q9EvfhliZsyhdlNjVnedUw=
`protect END_PROTECTED
