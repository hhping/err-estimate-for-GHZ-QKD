`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jg+EHdYEGQoCQYumxQ7u3KyBlgPfkFvq5b2XPEbk6SoarySEJw1wYvo3A3QLVcZg
RivjiZ/IfbrutdBYf3u3YmvqfsOy5vlDaMjjvMtZd7JJHazDu9Xn7pHCfjS9vhSL
fHh31fGSFwVHEZo60hPoQXfOd+atk0gN7WStQ6AKz2dVbrOt6q3qPla0rLCjVSpA
JncRK5GtFF/DI2hodwO9kD5eZAjBGdVIolYnpPTDNcuCEsz9TCkiAadRcY7fwmvL
I5bWwRZSygKITLLIZnSqJ1slxl147h6HnWtH3h8P5Q326ZfMCrE4UnxbSrj22d0N
NPHY9zVwdwXE39a4IGiPckqLgQ7YaU9d4mCnPZc23kuI0KAXUubBB3ddArFRduy3
v8IRg6wm0V5h43/NRBrDRO26l6jjJLpgzNGQJpWJqhRNjOa6vxff2DeLvzM/befk
t5K73ZDR6HA/gT2XchCHM69NRYFp0P0KLBqK6sCdvfX/sAYByhJauPDr8/8Vu456
7PA19Ojb6BdWj9tOcjXaWQrEuIvXw+PxWP4z/PRkLIS1/GpJKlR3RcY3BSD6ZArM
6XNpMH9+c+37t3I5kICA18Y3I/jaADsmvu/e03NErGEMHxL19bIJn4KnsMMHgdpR
7WUxqqqFjGJR+jrvtAKx/YRlgpklWUW7pitgaoxVrCcvW0dMt0sumcoFxrzb9kXr
UEnbwvkuIP2lE/C/aOPB1vPPfpT3qxly9Jp8Dc8aw6+KVkn/FlTnNjpUofnDgqGH
5HSIbe7JNC6gFFCTLnviOb2bUupc+XJXkyve9v+voe8h0/yyqisK82womPHfrmI7
d2jAzXSDaJf6eMP+JHwxNqXRwe2wqRSCcgDAs/s8H5SjnVwUExkYYOViqDn3YKUT
5ZgzFHj0QqMMO3Gtxiwa3IQAsqh2XEt7+y1jIa6/ra1F8KR8B6txKbyI7oDPoYNM
7fiGUkxm2QzNnIRB3RzJJiuLb7E4fKMB5dq/S79jukfWgJPJAPmYy3xsmYtplGgo
jo5K+shm12xKqFDTclYEZOeAWqL34F/EnOntha+gYkHOV2Zejmhyp2Nzk1LUmBCA
6Qc7kX0rDSFrTRdwpQx3zfPkEpeNhZNkUkBsrrKcx3ePE/J3ltRliW3/MFHzAttE
SBLdbOi4JaJLyVDwdyWSV9hmp+IfLHYN5HKN0oaNFwA59Fyx2SX95S8QPLr7dD4/
p+7vbrHLKlML35F3XS53Ka9jzV3csLfPB+55TldFKs+iSQWZLge//LWTUAsTGiOb
tr71A9tBzn8aPQGOU6ZRciFEo5ApuyA1RjkGisnXJo3yM0T9gM4SKodgdQR2AaAr
75ct5MjpIVqM1s3MlvU5wg==
`protect END_PROTECTED
