`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUzLjgu0UT/9gWZbsT71ANAAJSHDVpN0qizZBUc8p09f833rUlpM0Kdn26HExPC7
rt0M68l/Ch0GVjnAhowyw/lYaEyuR+RJzzXW7h8598nfyzWQwOUYPINJLTlfflgL
WhAXLh92lx0Tp4xEDB6nqPHYzLCGOPIc9CHjaKp7zjOwewXDRDlM/D0DukHuce1N
UdSY8d1hXXndkRpBuvs/fctzn7y4EnjLVtKP2FDhON5NgZQcbK3xIt6kfL+IlgpR
Ul7lZCywyuvNgK9HvyjRMYMido8n0CvqbMDdPDpUp9FIGLA5R9jdtmuwtBec8fpq
WYiKVFg9FQyAomb6BZdzA7RhOpq3Ph6UQGGQBstL2OLhCKdhRBOi4LcGkwyhqA6X
6eBcG1FWBG1BVxMcy03UYn+eZfHHWx9HhIIbCi/fAZ/4IFzohceJYHNP0qzAF2ma
7sJ9t/mDYqJd4YTZfNuSRHG7KHnf2Tk0q+bMyM7Tm44q6iXN2Syn7yypDizRZPkH
Sxj52TkYKTULKNJsj7NBdaCITPfrmwCQ1MhYV9fmWfznugCxckFEW70JBaf7vwlk
Lqtb6/NP3rp6vhfR8yjzTSMNPIq2fNruEhJh5C0q/ktF5or3/NRuXMWPeM2K9Uu5
bOr93Umv5+ESWSclovEU2Pv2wmngmHfgpLXeuOFJpwL3pWQ1ImLTobNl7253pCkg
5/ww1Eyjjm4L4ZxN0i7e2abK8kF5odKc7ZdrHVL4g475TBIk5gUFbo2qKRW/hCpt
Nw5m40EA/x79tTF//T6aB9BkWe5NlhN/VU0iOlKGiCtV6cCm2pHA7pyE8PigeANJ
T4M9OlLgaQZejTpM6l9IB+mD0G18YeCU1Sa0pW7d1vTA/Q/Ktl1mgUYyVAN9rynm
qenzP1KNM3smW3wmbVLlI2wSlZ1DCa9HekU8kvJdy8LwjtZMF3C+VCPFvy/OnTGT
vJXVgs+y8HOEXykcYWV5WaLWhgxBvV/HM5/AJNvcxcBCUCwce+8itrzsTt9PEOsF
s92NML8HLY/pPZ3IsM373vVcSJD1IatwuYVf/BEeAZ0eNCyOySuU1ofJNxzPvFco
Wy0g8OEsZKva9kfUUQxtITuJnL8APkfPPcJJ95/lbhwdAc+90aK/cIkoxm7yxoiQ
Y5stlBHTJO0Afs3DPlm/GvcZCeYhE2xDElqU6XCl0yzYEeFV1yJaDgA3aIe60OAz
NXtqfNYa+5EVPAo4lI1EfHDly3EPuQCph4cLKOTUOIl2bul8TxP2DvOCZxwhlMrt
NPUnIkkXrTPBdhC4XJZf4U+eZkWOH0TfC4wANTDOHsDilSNHyViQRKjMW5YCc5wb
1GBrhBQOy8Rc+Ru/bpsyOUSg9exF8pKgMnILyqG/wdPOUFWeCTH6TkPjhS/Ay2Og
T8qQE3gmLRf3NmMrOVPPgQ==
`protect END_PROTECTED
