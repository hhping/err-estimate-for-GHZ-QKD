`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20aXtgWr7bI/y4SXhJnnAavAB1j9Q4hlxFaScP+iRPgaW2fQSB2WsayeCnHLpd4E
AALmeGnvbBtr+8uS2WY4nrcCaIrZebCPG8FRxsu2p6JKSIu+KSXiymM0Zp1Wcn3n
h2+x/G6px/e/E9JB/EuGARO1uY/LVPpf/aAMXzA0p0XP0uWLFP0cPkLfR3ecM4wk
KnHYhyv7XLuw1fax/xC/tA4V1Sh5FYcLcwiUMHJgbo0ow1LK+CD3PLla1+xOWAEc
in9ONoHREpYKoDH9ocNUfebSrklOnDvz67lpHF/QTvMnRzUWjSkvJFJOfrVlELjL
lUaomNSwCFH6ij5OziJuhlDgVYqzlu6Nu9c8xtvAHsbeG1MChXrh4gDXelwGNT/1
BF572bdk8arGxejSiTJKxEuKQ8lGwNuWUAeaYBDjr0zZ7PoL2ezNCKnSC2fWXuoY
aPIS9DaniCImG9k9if5HrHWXG4WkMdx9cxTtyFdYCzg6vPeagKGSFGp4hsfLpkGt
rUx7b9G3kx5k+d3zg003S+Jhvh6WLEVXkTnOogdGH6Xs+mckWhkFr7eWn7B/O6tb
5RQZI4gHYcULpDpV2uD0EQ==
`protect END_PROTECTED
