`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLWGOAPuRFEeXrXjZZicPMwyyZTTC54dzl79hUjGRj5C2ZOQk9LVp+6otBzB8k+e
BbEC011ncpZCQDjXtAnCI/xhO6hgaAIsa3NcJ2gaH+kiqdd+gKCWOYbwfnKuFJXa
tdEsiwHwEk4mGrGpO0Tbked9cXE9R7b5bmqovSpIzq/qqsu5Kwj+VDlh+o6gz6Gk
k+dWmAREHdYzIb1H23aYmo4osN1wUFBEXm1/Gd+oBslKHgxNu0gQWoSozSIE4dgs
apt5oKnsVHshh1/wVEDqiBH2rCJW+QPxbxkPCqZCgxOiqNb+jZXDsGbJhqP6EoRj
dBbxgg+TDJ3iDC7fHQCNKyecszYaMSMBSAnggCncBjycgiQBDPx7+62VQy5uoY9o
WVt9OCuJ+6j8GKX8rSg5UHrrz3q7ddrgs023Xn8AhtIiE0eqThe6ZKyAz5Jeb0DA
ItiO2gM2AqSizLv2sTzNzrVvmRZLkqUGfeDQxelwVA8RqOZ8swM2umzAE6H5oOh+
ntYAv64V7u2NlIEeTacYRQwPH6DoIWr8eLeReFrKAOYlXx2uVHwo0mzqP9Hbe9aq
O8bkTwwTFmGkVnsVlMb86O7AcxOgbm+5y3pIt67OtuMO+p4qu5Caf3Qn2uEBW4p2
LEr2gINjm5IJ6VBqlYvcVvkJaz891NSoawanUmhOi1M=
`protect END_PROTECTED
