`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPanGBHglBRm9lmA0a9r5Z7DvI8V/0W8+h3CkUrH7TcMDcl2Re1Mr+M6HV9vSJzm
SESd47jfnBAiih+L88Q4mtwF4AfsyMoigQ/k0avKlu4LGJNtHuFatynvEcyS9gWE
LgWKGGqWFmukJ828A0008WIsB0gBq86ryPkLbTAHxFtMeQEKgRJwGMF53sDCOEjM
nHpYTpsSV05m2JNvvYf6hh1vQx196LjzWa/LuJ4KTGgY8jfG/QYHAVPW8qlcA+aQ
VFX+llN83bKij6VFkl0KUWNl4uJCZjUuKU01r7VYGBcFwot/lYRJKayV5ZdRIu3X
96HxMbVI1vRYpxX1N+BVeHmDWqI8+t5xv5HMEinvPy+Opk5i9WOqfZMeM3wGUqD5
ir2ZO+o02booH7N7KFqCrZ1NPcW6j/QooUrxQZr5lDCTx/vxfZqT6qIQAnQ3HpR5
1obs4TDXwwy7+ACgsYPOFfi2c5eFxAVZhzaJDNhsUqgTLa0UFHBRKZgWwJ+hm/R3
HaStJzGxwdja2Y0s88p+gw==
`protect END_PROTECTED
