`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZxKSHVy4cHVfVX3OjhQHsKWrE9h9+N8OryrOcDCzuHQBy/9ujmI2EtPqNZj8SBr
nPDUnlGFQezOzg4d1AyLdWbYr/XimjcskJUj8wiHljifzckFkMX4M1C+AkIHR8Pj
fLijN+J0yBdQrpgIRvDWFrYZ68xJKcIBMsa+v6ZVii24o30uYmWEpvfkRJTnvf/T
F1RUP3uwWTWY07zCnyPz4WMcefMcFfY3EHGvifs2HLHCWEBgQVWCbbzN6R1kmbXj
qvMXtEMQrL0QBb0XovmPaO5feiyfQEG7ZP3syHcmELOlSF9Co1gsWrUrCAC/lwTw
ncA9j/pTcMcDsUQ9oAM/4aF+GvKntHKTEgJ6SXnM47KvoYIctDYdJjYZszLXAeLJ
ASVMXMgwPvlec42fhSe46ECeorWZ1KJ9n5XaXaUeMUo6sqI9xpqT0RV+H4SjKty9
dYOwetFm7OAQ0p4GABOX3PhX/c4lpGrhcdgq0XtkXFpJZm56RV1H626tOHLJ3zfW
WcEi9+Ic2GJYcHdvGFCZW3kQxffHfVP9grTafX4N1E8+8c5KeFcwAcCCcmcUgB2R
Q/FhdLmdJjLyR39AvwaV7ge2ASxs7KwgGJjYHlpkeyNEPbNPeYdoQ1ENHKkSelhp
g8jZVnedNnihF7s7fdso7cCZdGYig5KJ3BR0rtzmXmTVPX46Ljye0bqK+2jVgDcZ
bIz+wFnU7on3B4YugzA1KRx5ERH6FiBamwqNioXK1PJ/g+ZwqjPL10dUzTFE+tWL
/3FGgVODV5ARS5OdYOh3mg==
`protect END_PROTECTED
