`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cmNiSvWRU7vqId5BgEFrPuC1yp6DLlLklg3GNRdGvsivwWDqG70uAkV4GD7K7JaF
DJ8gvchCVpxfogy7giavd4Qqkom1uCq8nz9NQ2Dp3iaxIdhn9kan4o8GiQ9kQjQ1
uE+tUzN9l2zq+IhMFJduqH7IG/0GzR+vIkb0NTyG275d1a/TLkELTLFBkMMfywFl
r0Ct1R2DSSySB654lbna6U4tvZDsFqb6VDfKJ0KgXGcyWGKlFpPjf9yPsZBUx+HY
hOdrKiNedeWsL5ZxdDdgJAjOn3Ph1Wa0cIxMI6Fdt59SyAfqB1vWN7Jqw7S9Bs0b
7IbDsf6PjLmQHxX6l0cFbSWlGDcOC4tbASnITOMGypHn16Cl4PjmVcOoSI6i1i9O
HuTOPdyMH0XWyCSU69ZTGtIsOsXfuAUNdg+8GqcEEFarrWNVK0RNu8Pt6vzu0icD
lJ/JyhNLU+TPI3Tnb8PuatixyAF4CU9uu6jLCtpdjT31noXLer21bsPoZCbuPAPC
isdN0qRzDh3OC0ow7ZPXy7uQJYxm75hImv9A7X49aehlnLgsdsQjv2yFS7huysar
YC2FyReJSmnr9GUDPAVynA==
`protect END_PROTECTED
