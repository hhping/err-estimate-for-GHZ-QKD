`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIXp5gSVDeU+q7JP28N3HjMRUNAFM98lvmbpsFrVb1Owt0NCcDaZLuEwhS/NGCGg
ldOjo1eh7j3BogHleYebY+2CQ2lZ1X54Gsdw2dLnuGfXTm/ahyGeyRtjq/h6McpJ
FD5eNQfikjwkgdJcpK2E2LPrO/w7vhsd7FndnV41OBWMjxMinWbrpV7hjZHvv6zb
SgNk0O1q3bSU/8ssal6eXkZ/je091EItqQJMTW90nIJ5yaBWiMAPloytbFDUKT/i
gOO39wlXJNZsilQpVXPjALhZd5/Ox4X3rwupgQux2kwHbc3wcvcjgWRyNul5HCFB
YNLPJ9M+1szLSForZYa7Q6N6LYQmFoGSbtJLRBPqYy0Vlmpry7kI4Q8RYUVdIqLh
zwM42d4B817OmUFGSmHVZHAoxb6+1aKcLgw+POhf6Vx5XYZ1pO9OEKo42embHa2v
lRw+rpFsPuFvBHkfV5BNqtLWEQDd7lHUkMm4FD0s+fl2jul/wIl3lGkpdP2e+sk7
YOWTc7vkwharkInNHR55+2c3XG+QBA1xXvSPBaSKv9mPJafDSMCAZ/A72MtfU3h6
eyYfgTh/+KyzzXbfHTcqVZ+eR/207EiKYCjsRiWeHr0aJvZoIjWczskuiEoBmpRY
WZDIfCq0G5j4lbHRVloWfgGjXBecS041x0jzPpbeqvAvp23ngaN//hcjDC9f4uro
1OYfLdefl5Hg2cSaG+gVHwgTjcDfvjpQdb2GL3naC1oXb5Rq1IyYWvjqSvRQBrEj
CfZmqb35YHPINlkK9u6RudJrAcaqN4Pr6uuo6z8xSY1GMwf6Ek/x+FqmyLz7G/CA
cJqkd4WrbBTfKAPVlTjiCory2fURQ549rTf7rKbyhG69Wem9f/h0yZqO/adZZMjh
j8GvDmN/1soWkjRSpjX/TI9WmRPcRhp4+a97CIL4zcsF4X2ZD8YlOu90drz+2bLF
hIFW4jEKpXOs/PsDyrYdpYLAz4W+DQXejQNnCb965TgXNdjhF5WkY1LIkdH8ZfLO
e5S++OO99hdEQWRI9N+3Zt/Gd6dCD+KMtWULUTvoDPK7xPG4RnfTSAlFbMfMLfJq
lTX+jJ/fRSrXSFw64pBr+eVM89kesN19xCPVRvN7fTyW6BeJGAaCswTCde16bJJW
Lt1q1E5sKhfMfbFgV79LaWCzNKENOnenQ9zj1hk8XFGu1GV1SAlW3NU8TR/02yw1
Mmq6c5aEq64CZk+FwCsB/K59ZyDVLRqZmoNAnBZhM3I=
`protect END_PROTECTED
