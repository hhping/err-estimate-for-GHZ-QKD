`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9JdTUS6+phfvneaNKYGBV02t3jkMqaAKi2GN/ltiwV1+2SqxnkDX+k4bdKT729Vq
HPOc3tKUnvXKiF0ZjaT3SV2XkRumtgTxlfi0+8IsgAKKfJAvq4IYWQfY16CN3RWI
pJhzJgB3H/nXI9ZP55vEbzA90wIgLdFf3I9GIHIKPJoama6AyWDiJDfjxwqrHfhX
zT6SYRltW/b0Lf/ta4pMxIYDXhNuSu3gDkd+iQ4PKFi5yhVXzISbYyVTJYtxIKJM
CLQ9w4GEJte8JmNNUTQdqZav/WFagq982JL/csoSKxySkhJvZqLVSDKZx0SU4r1s
trzKmnXPXQ5wN2r13360JjkrotElKlWNJJ3ZeZRTaNBT42jPsTIpBs/Iqo9Nin3V
neB0U3k0IpAPA7JmeaZx9Iaov2ChHz5++nzUi+3ufmu3nUCRLJBrYi11yzWuEDN/
JRpNFbDNxGUt6aVpcB8U8lJqFx50d693TtgJLrPZ5i11xabLUx8osqN3YluYEETH
sFnVojrnkr1WkyLOpF8XhxT3RdTNJOnet7IF1qEIiRchSoX7VJwSgkWSI5MlqWbh
eWvRLDmvvuR5TNTzphaJ9JnBlqey5zAG+ntO+N9Bt72S2Q8Azs6WPaCJPksi2gHx
tsjHg6BUEK8Af/8ezxuptbtp0rksRGQ5F2MLO3wF+pchIfgA5Y5dvi2wglTWoC3t
LlNxHxSKX20g3mvlM62sluk5IO+IrOde7XRKgDmS1lMAsF/w1lPWBSwAjgjZEXDO
zD0QIxgGPPG2q7lJeMxKcdknbE0nGu2UYSeRrO2IysuNTYsvgAXkeyvmnJf2qdJ8
BC7m2kOf7FSNpI1rducJ3O6zMpg6QgG4OByumsiLuGlAUkJZRYTKPQIllW3buRRV
/yR41BsvfE07EWR3C86rP95EG1s4b6sSUTxp0HrYKEnZ1jI7g+4FZhZE1DrI2NIi
MQRCmrfqUL1ZuF7oSl/qPRm1dj4TfJ2tB5EMajtv07rjPEfz4cFOBJveJB8x5BWu
pRf4zzguJv3swgSTiMshUM2veKSJuw2EKZDcuJgWR0CUcv9GQRkKCF0m9QjW95xi
yTTCqaZKExQGbsAkgdKu5OJRIAy28CZX1z56QNmPFbhQ/MgVytDeVa1IdW4mc3jD
AC1yRTts75+7RtSqBrrVh+iKhYYsK73JH8+FLecLwwD2d6/s2ZesIBgcWu+XwHV/
ow3fh7xxd0nwqPk31NeyOnXi7+YiPDRTYbskpKDf1RX/Brh6T7QOFaVRXPpWfas7
Mxbeabyxx3BTZU6ve/2QCS+9j1AzS6mTWUhYXM2mVyg=
`protect END_PROTECTED
