`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6InPzVprnFGnFkDC4JNAfDW3DVYxkGW7av6IPm9E5L+7gq8hYIFYHXvdXJ/BGw1C
5ziQN0Y6IldCF0j429Vkc5R6yaMXl7IQGVfH5/xVixDS7jJDCfvjUSNHyP3F3GQ9
t15PMu6khq3d/EO5jcwkeWB1VHTgA8jpUMN1L3T4IF/bzqJgYGMtljlr8wwZGlvV
uBQjL9pgUB/kbd93pbW1ervmnUHbzVv4bR2eq2GOhn+jTc+j2VndgmirnQ0dvRuZ
TXHaQK4bZpKuOlMAj2Q012O8nhxvBgZcQSxMkJ13k7Rv9osk1/JJTrAE5TxPUPPa
HbcC+Ex5ZGmvHwGKpQSU2MH3nH+r0mCez/QEE2eAu1bcOewuhZNZeS0S2oy+iXy1
DBtGmUC4q7P6VUZ+RKEjidEwj6yPXCpN/Ssonm347J4JnKBwXyAD84/M4SQ8F9Rz
QySqqgFlmM8wdXp76RwSyMC0YUNyT6jZXdfpd3i5OZKRnJxH0WostY2vHTJOcesu
95MzRsasAm0ySlb/opj8yVbXtdTg5adYTbrCR7CIRWN5JYADfEQyL5Z2LhP9f+VQ
NAk+RKRmu7d2zI6Pirc6UICNLcYsG/VCL2zgTyMKSfT3edec5E1sqxBVW3SoiXqc
zmKG1ndoDEJhFrMM099ccY919Bys1H5drsx98pY5pKwwhjqZ7Dqxc0ltq0nwi06J
VkZto7sS2Ogo8cXkhyCasn5pJBt9VCnW8uOBOzv/NzxHYVFtgQ1MRS+TWdFjMhPc
TOFQQARVd+IE7I0varXjnGIYVCbu9vlB6jlhxROay2/EYX2w3zrCSm5WqR3I+e+x
`protect END_PROTECTED
