`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RzVrXjmWNaPnyuzCV1CkQ+bXgvCCU3QyIt/zqSE8Xqlx2IzsbK5DZVqsaJu1h3HN
mrg19i2jxU/64qCG36cArVszK0cPCApkxZVJJHtgUI+CK0n9Ji+zvIaJms+CRgWL
6Vv2xvzxINHwTV1kLZmHVV26ZfDKex6UFOpL658CX25kh6uExe23ZgrGZCjB2gbo
PGkpU8udYV4l+y/ITiASxX+tMSIqI4/GP2d/f6MyjXwZ/AbYN/UD/UUa5S3a+qQc
ZIOF5upUYAHhIva7OodEXlTWDssjUYwc17zNrCq8Wblkqv7GjSDADkFY7g02ze2u
Dcc+/vKBV5mSPM4VQqF3FL5wOtfAJtq8A8Dd/A1i6XDvwpvXTuR960dIyF+MGrMN
Vrgy2tPYmVabZOAwuMGCGX6L87RGtYj1gZyGNc0bsE4Olkh4sRodpy17z6LorrH9
ZGoYLxjB2CWKRDEejAoqYNX2NpfOuGJgTn6uiMTOEJV15Ctpwls4hse6KwDQdKu3
EVJi6WNHheu5Loin6KIn9Cwm6pCWZArVIQTl+0ytEKlpee5CbMieGnqZ9WWFO7GC
TAsk/6focxuXJpHf53+zCXfVQlt03REz5RsYeY9ezE6UD8wciuf7PizDWticRvOu
/Pz92ouzNSIK6favQ5KkzKsrcnQDnsklJ0rJRkqPSTGKfGHniDA4lgAnFrX350pQ
r3W1Oq2Mp+//nIyNxZXvMLKpe0L+VD7DUhpR+bxvrcS7jGn24VEfQRFKcJiD8bF7
Cx59WmmyBHFiFE0NBmFcLUa3bTauhBFx4ZPaUFsaLUBA/zWqvraCoykirPovF9RF
8PRXtF7DJUi5IAHq2SADjpOIXNNU8pdqqDZ/mS0bsjLoz2TUzeX7AvMoR2m1mS5p
eu47MPtqb5pQf4CUDDJ0tljRhruFxxa5QnO8fU+g3M3ZGnVZ/5VkMrdt8ToL5L8g
2jY2oLzszKdBQ9dpNJkEs3Cz0tN37GK9QOsc/FGO225QvhlAElsm9foXJ2FiCBIx
OaZPga8O4fehzU+xSa7iUtLlt8jkzUhEnOaMLjjSiiArNnYNJwEUISU45QcTo8du
UFaz57ix8vHSyXRzjC922Ja/WytBf/1+WKXrnp32sLvmUFWKLwfsEOMABTiLkZoz
wBn8IiSZ6OajvA/lyT8t8YQRvtRdBdzmb8g6uHyCxGaSR3w9kaQa4CUbFhRG7RM4
EVhEUPDRd1QTT3c4Iv2xvMrirj0RmJWHTONUQ6XDsKnObWrsdjKOVGuTNlHEFeqX
xplahipTZTzZ8dHgG34H1Ze0z/0xAwX/JvkvX9qed+sHUmzbxsiBCWZoHR/npt6/
pnuc9VPsW/4Gwq3ul5YEURviQ4HJlJj+h7nGpg82ek5QCxHvKiKUu4x2wJv/NqxJ
yy6C/yIKdoaJ9XYAvFd6jYBEv8kcX7cQbiUJObq6n1EdGQT/uZRhVJcMON3CmpKn
tGIC9gutaHwclSUIJInvqoW6VzHIpj9PEC64qxDjff2qyO63OkuQK9q/LGkMDxct
IH16chcHyePiTTunPaLuTEFj8OM9L8i7j+76C/jy+hdAhFI8mGbfvf02bmpT8KNB
ekDocVYmkJFcv6piJpLlANBB3MbEomxRX7bY6zRgjrTgLQL0vdcY9ZZUkoLnM/x8
ltfCSlS5tgsZSUc0EjR/xvPzFoUlp9A8t8jL0Pon4uhwsBtzpkGARmUlvtLHenXU
W7qJ/oDglj5SMBNzz20NvMynIE1wsauD8YxltQv1YOkQ8VhH0/839htT2EePpqQd
PknTnftWDGnv3PqqyUwzHZabwVDoCgBvwxLtw6P7b+O4JwcixC9k2Q2uwZvn0+oS
apYG6HByKEgfi4s4fkobnpsH5He4H7ChAtc80OoOu+MvwEwVAPRXKNeoAqv4cdwQ
+j6qHQogIfAub9Xb58VLlPqZidzSlmTOKKCYiW0Yvi/2XGinr/1K613/0JBffzKY
JKN4C1FqnZYsTGo4pqW9P/K5hK/AlmjL6HY9KfoG/AWQ2iVGz5uM8K2I+6CyuO1X
JSMcTzrSjDKWNXaWDxmr65RxaodcnYD4Yhq34bzjfJLvNwed/0ceCnAZhRxcsK6y
k7XaLH6vlotfxUs/gA4HM4FWjviQF1evt+RGolSUQqwEnN2+aI+wy+u9VVKyZEL6
`protect END_PROTECTED
