`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iT8yIzbsnyR41sn/AepujXFwb90oeq6vxg4eKvkAybzOgmS2X4z8qK6CkMdjxAqR
GahbdBfqcI55GgyDDIK0Rq4yuoZ3M0Fb+nCB49NoE/vm2k0hlxl/1FvxovoWasio
jMazPRMIAj2/s21JPV9vYJG5h3B00ezE5IxId5EDeX62wZEuSQbMllrkxDltdBIZ
SvYl1T9GoeKmGbEb5RvfF7lg4q/kvky35+/+iR33PvyoQlEU5q3UQS7SgwOyrLmG
h+KWPDIx3v9zqlcvcLsMlgG92dpVv8PuUsyqpXSlhAY/qIkpwopiYvrj1g+KBMRD
o5IB3ng6ZD/t07ko1ZeRxyxP5ikkmrg1jCjSjJVWuVKUVSWT8jfLq1fQXhjRro7n
6PxuDWztpps2r8qeX1dvaFWle8mOouVGGoaWews4ddyyoBnDTw8v+35R07+QauoU
yzvQKy4FQADFt3Maq9gOlmWfwmwc3OYr2xf99bg2NxjYW4ecHcSX2xOwhvRqHhhq
xYQjCM10sOQqCuorAm52QjdP9/dGVdHg9HcunuCfqJXvE2rK3fnbsgPspcHgMLMi
gKpoC/jOKtb/zSjLVz6Rz3h7gCGzHnrL3If6nya1RkwApuMcZxTe+7Z9SFybEDuX
U0mg/yhTihyMpOL7frFri4PI06jIrR8FWErnGexzEIBvIw3HG7wA2gXpz7M8eKnK
MFmZE0npExjlfHo8kuTSeMUIwZMyN4HHJDMBd0E6fA0FITErtULni+Fn11CLvNvN
99802D7uqIzm69Vjcyuat97JQGcxvB4Br3CIo2ac41/WdxQjY3O3ETTZTJB+QmXg
QSJj7PQtHALsoNkoes5wOmN2YUzg6ygqq8nz3fFSrP+c0E9QprvS1Mk9Y3lO3lLa
1UbHbpV70e78qPKl/FSpUi1Y6Oepjsy9TgxcUKd6qD0KjOZ3muDONS+4mEZax/E+
TbKHnRBXsgQ7jCvNcFCyYxkJESVSZgOY5+WmANvwYHwGB/u4TwAyLiQLGyePd7Gb
j9JeZDF5gNYlqs4k4zo3kcc7SpHlobvgJCJydR1L1nf4pzZAYxiDMKMlZcuv8y4i
3I2C4arhbH57oPXq7J7PQwa0UhhLZvvaf8khuBkqWFWlxjyPH3q395q5iMQ9/fpD
1DylSd1vysYbzFn+Uem2TiMBNj7mcw6HjTLXOvv50tMns4VcaXae33YxFLa9Dd/G
9Lxo9dXNoqzEssEBhGSSlmEOxjaJYcAHhMrN4ZpWWDz7VVlOlTmOenDa0/KO+rVJ
Q6npHUn4ofCqncmtjBHZXQmS+2LP1uR/815N9FVPvVk03W/1CQ0mUsMVPXAx2qM5
tdk1Eu9ArJxs09L+jxnFkdsd58LLdOC+vBFX3ku1zUBGxXc+nEwmV7Qe5wWrEkl1
y1bszm9F0HRCB/u/GN8jtFFAShG6pCWvwRXGmgDYENsCx3eZ6eDhrX4lqL46s7BQ
sHzXapn4OM32xFpSLStdVprZOSs4+Nm3eptXsPP8Apm1Du+/7czwMK3NoB6E1bDq
Q5hV8wV/4zQliWellznqaokynsdlaNMhyjxD2VKQnXpFLYcGRGP9fn/qaEdOCIiB
IWk6f2F8QKjKi3NjdRriKfcXD8qHsnx/MD2uWcXKf/RUqDpdQ3CtgJkh2hyXEBky
9xRdMzHvjt6haZOaH62jnG0NIsWSR+t//iHY+Y8axWwdhfvwShbeCFxvBT5VYjno
1sgLmmrzmPq4v5+Zg1N+m3XizQwNi7hUtd3WYYKcAcs+rMFQtc+oT6tB0hsWKEGE
yq5c0kLICDSNKvQA9+C9/+iaodOBP24JWvTfpWU7WDH/OWBZcbfTatyXYx1Kr6hH
YowcO+x14oXlE5XIK2e85/t2L10TbMrLVAyocS/Q/Cz1CkiBWwRjZPXc+VI2W6p7
rLlUw7Jsw/v3kw+2hgG/dHVq0LWgc3C3CSQkZhxzeo0xcgAaXfW5x6uqYrJiGuA9
G97Ykyv/U2USqt7wCHfHRXS8xYFylI2T2gD+smgbFQeh5zhaFPPegOnuo8wLfvtK
eiy1qVsHvJ0rym8Vzh0WIwAX6CyLV0WrjxEJvR3zJ2zVxMD0n0BhDqwRUDUhzTaa
W4NeTXp+Wz+BCamPBtVVQkraHFWiIjRnuHWVzhJVbdOyHCuGJ3Umxrbh5tCT/Xp5
/IiGZ4iX9bZbQ8mJ+Bzf34Ck976+/Eg05+8qZZ20ifuw/SOMxdCNQq0exsu0+CPx
rad3fs8zemkp8052L2ABxgMJTWeVU9B2XSfsRUidrFKvz6wGl+BcvzkdTWiqb1fT
IWTXnTM24iHp/qTdUNvU2oX5WrjONY0f7F00EiIx1DlDvxBUKI+KjJECMHxVpOZf
48aNtfnxnUQLoxUPW7F+8nD6hkZPWqgT5WVaTlmYZgMw4Mbo5bXS222ZIXmLGpSI
UGb/dSLblcmOKppBE3yoygbuS/tFYSeUUDGBvBpEvu/rWTtTPYFmiQqCmmVwmOet
u4ljG+mIIUVKo1I+oI/tQJWI04U9nDzzR5fO08nsE6buvJ5zIOJAMR1uT+vKWjHK
HVq23O60VlYEz7EERjapmBmHZDs0o6NDawAl+6x0HCrU1ECdcsFzHmwO9LgtJZtd
YNNG9RS52byMIXdBWz7B2DdUGQaCs8Erdbp2AQIzo25hlpt4xh2w7WZ+omziJsvT
GVVidpww5MF9lmFeuEqyXKmhS2c1X43DSUzwGuXeke3Q/+wlavB7P7NDeXTCATxi
potHEfEHUiPEDyBguk69zpvMyDCRLzSYuAKFJ9Q8xAwAcyqb41rLD+AW1orNEdes
1et1RVXeNap3JA2yTATra62mHZ5OARqtzEX843QuXE9rzSr8bS4YBMSaIivtGTDv
30lflyVVtlZ81dpoPYcl1zV75Gbet+ME8Sd0FZKu7d1tV1osZ8IslmotJ6GL2GY5
ZmoJBxUJzzyKr2+QheFOtRZm4kyXAqI7z2mm35TRd8BpbA9PCyaURi3eDar9CX6e
DwEvxmow1T6wkyCLsey/0RpHH2xnrmTeJ8UURR2ojK5vmqOBS1NFJmBtjtV91Kxm
wM8JvwQ4BkioG7kqtJowuU/3gVwrJ3Gk7GAZe1En+ssvF6IKipsjlmYH62hzpMEF
2Z/x/5UFLJxLeRB7pkQfzTH+t7czBTxNGtjhDTppmxi7aHF2M16O5gl0qVJ/gl7e
rojp6hj9ZIyjJkXBcrqZ9NAZE8P9j2I1e9xC34RYzAdzkmFD6A7cP2GTS8wCq3ZX
Eobz2TLapYy/rf9y/OUjkUlrZlW5n1H6HB1o9ujqodBEDKkNmPW0sloWjD9dq+Ie
VebNS6uXdcki64r8dm5qqNkPbmiJ7PWpW5rIRx+tJo3H9HAX+d7tywxggXnbnPJ1
x68mJvvyW3SXpc5Nyqr8/0pKry3WeaM3iEaPsJnXMd5Jhlv1PYU52t19NtzVHJk4
3TSVu5YW8pn5ju8Wn8eNv7DI66oILU4J08OQDzP4/WgHIcVwJ2G/Pp6LoB5jSpld
GHPE8Kjk/HJdLHR91Y6PcHgUGsenTSTqqQ4HI0ek6uGilTE9yUWo1Dy90dliS2na
5fRp62hxPrdAsTwhPDTQR9rYW3EDlotSXu3XHFaT9ZX6J/ogenD+XZOIzpIz4aSm
wCRLmAScr64eg0R5NwG2RVlQj3fQQut6Ak8Mix2nz3tAHKKPOiMAMZFfKiWCdh6R
qb2R6dzjy/y7uGOU6PWVvIBEFr7oN2scKeLH9VLSSDDteZMFJDFnzjwl3dkO+XCl
cbuyMKo8RP8rU2XYZGEfkvs89pzShgQmXVlpXs76z364sSSuzWf0nV89f07m65/J
PreFDXpnX1xGLwt8p1n8PsyurN9djlv27rVrVj/isRaCFlrHQ8z1hQRSpjWN4cxq
QGISuL41f2xXEB7cI6wd4nPiFtEMe4BmEj4mTQc+qJuV5qD2TapgySlapduVf9T8
wGjyimVTKNquh7dnyf4dVNuHYUOk4pLapiqniaUfSla2jq8lYcNgMnp0+13ZezUM
xTJOl9cr+ZEEtXiUlzr0r43YuYuUMZRz6gEgalhed4mY6M8suOgdI4aTaQUM6BRN
Y+binwi4K4nGBsSDp3U5VmJ0CJGt+EESuj+0aQ4UQnFNSP7rLxo07lcS+o3WeXDe
1m0XMiB3vGhSk2aQKtTettmOfLktk0Q2D2z86Y10XDOZWqfYYvklAqEn1dnxmcYY
AemiyHNAGn8lRclO6Mdn4JcRnAbbCo0a5Dkywt+8L/9iSmLErJZTDZZnUVzGlx4L
JK5VxM97O/5cusu7eQ9zF8XQhcr0fQPDrmL7k528IWZk2vGeL1YgAVMkQ/vH8aHq
OnlFIPcyDdmIowndAK+NmAIJd/KuNplMWOMpS/K2Bmm5iSUiQJ9D0zm1WrAC/mgz
QK4dLfTdvulR8nZ0/LW8Ab3NNnwxhYHhW3zRlO+o3EYnz2Vlo/hduVHEYbgLOBD4
nCu6gY9263majVpp6O6KOl8DFTeglvT+OqP4RMJj+V7PjpIoGHgIC+Km3qt0/R9u
1dvRI6Z/ASjY7TX/oaqFfBgPGDWN9bHOxvy+SJSiS88q/nhoZ7HA2KdUQnfgvf7m
Sg8knbZ9P9ij1q55/n8Fzg+LPLW4lhvgYWH9EJi6Z7b/8a7tuq8rGpAok1M3HNt8
ZfpYeuBWm979+IqVT69Ayx7VbWedoFojwy6Z5V2OjJMjPedRzujcdtLHHXE7m2qa
Bwn++05YHDYtTLlZ4j7cU2qDDOgkPk7bVFvNYGmDrjsXH7j67YXT72lqHGLBHzxo
AC0Zf1MqAgQWc+VtqiuMH6vBEE67mYGHn+IaySsYdak7UAUcJTDhkE1cQHfVooRo
n7j0xoTEs0/kiIqIhk4+im9oIg7BcIZjmVDN0HO0MVNL+34V6GesUXuATNl4ILxH
2Rwff4r6ZxIklykhElsZ/KaiEXntQ2ZvLgFS6ds/2wnQI5u6nWr04rQqX05JAgMl
hRtFKouk8HROJd3DGi9zFj3Dk3lE8hZN64QD/YW3HsKXNmTQSFL2oSoGWlTgkzP3
ky1XpKNJSdyBeozDCoA9jOV5Wm3weIZcT3EOwCILhVGwdPGQ3NVlTWjCGwcZUopK
ixQel+/px6kO59xwuQXq9Fs+O3KvSIHHdyi9AlfMCq/v4RoMTbnCTGnvTv5+zVqg
9D1cNQH8r6rHFwUcUm97eemkRpd/t8YgFO5sMsiU/ZePruppUsExLr6q4Qbn49mC
5GSmyfkfPUIgIARUpO2S6c/gphDQE/HssXcj4/IUKKm1nRRCiCkU1lv0Xy3KABFA
6Plg5VRZIPzsfILybpBSQJURwEt0SozoaVfU3ZVjDq/4+MNU8i9OI9PRDN+pKVJ9
9V4CIjTpmY8XcUX6Nt7rjIMxLAz/GCc64lO/YVuBHT89hYtmh6EBLYz+MOgKJlF5
npSqb9V6dIZQVuXQQmsQZh4OD88l0a5UlULvDy12K96O3NNkvw/wPlcvsXt95o0c
vTxQRe7TaO9GOV8QF3zQpyuQsLb7eYAiLceMjiMzNT0TfCFmMB53kCru1ARGqHBA
cggih78rY7LpPoS7IeslWgFORbYeTYPYBQYxVYzCS3HvFYpjKRUhz3puvhMMQabY
g//2MNL4CDJnRgCz1k25JyXcJL+/3zvrIPq+h7APKu7zKcY4pqIsUd5AO4vDdpCt
ETh1o7i5ZQysPED8s5JXhAovKeImHra2JoXqKY1BzhYswIWJvr7k4Z57C0QU+ip/
lBz9TgHWZvL9QXvj/UHZBWZr8K/x8BGeCBZsL6lQI1h57w5dD60c73MVkAnqadSS
QXKKi4Vtx+6CpU/g1c3lXSB/I1Nk2P4dy2OmEzN+seUMHQiplHPjyooUqo7v8jVp
FpUJdxk8sNQt0TE8cAseqM7vxcgwhnz6rcpy09Dfeo7A0VCZzgst/Hqpl0lT9SZm
zw4ppg+a47YyU1TXLHHKTD/mTVTZ9eubRrXvPt8rkFZpDFD1pwE417U2TION4XZN
4H0CirA3ugodtfxoZkpt8GLDRhs2vS7lgD1kKa7AtVMbAWB5Jzx9xQR63UHB1uxF
I5XF01Z8glQBuftRUgnwsCLOYDVPGpaf+j/WJbdfUAj5oCzBaR/uDSejIy1t5wtP
x7Y6a9d9nn11uHmv7plaN9AYgJtUP3fEq0gPJXGVB6CiAnrXaXoa5IfH2I6KDlDx
mGFEAeOsx32i3gS7YCdBAt0bewx+7iUFpWnXSzu+QZk9ddn0TTcZafpIFSke8Ck0
eNDveU6snCB4sdtmGd3QIMnxLyTqhrWYcPzFstuN4DOhdgRumcy5jcli88cs3oNM
GahpttBUwXdG0wLNj7vcP/j22PjOfOmXT39zI7f1jhLDPT67KIlbS11B9D0HoN0k
vYMzRfbkefqV9x7id+f2JSstIMg4BPndxvwRhc6byui+WWDjqsZoPRwzj2O0ar0T
RCOWNgmcpY0Grt9TdA94Qb8n6fGu+rLVCB6hQD+cYiDSDLKryBj8Pf9nrrSl81MW
FlBC7/e70qs25LxRQxYaTBjA0903f7jILUxSs1S9/Y0Fe+SeYPufV9J8FtNHmwvz
FSzZJzqFOZdex8JEWNJ7FDj/Z705VXWjl61fHKed2Joc95rdWQPr7uqAw6lQ7nNM
bIP0CDxSGl03LK4/Erobw9xwEFqbiINWYsw16Vv8VDFMC3euW3SyKsc/1Y/M/xoD
f1s/CP48gxprvH8alQxM/MXPcFsaxobj0ziKP3a/XE6I4rEIKvtSKX5hAKR4mSm6
XWAJbEzeI++rmfuXn8FhzBZj/6/mLFID7JBhdqrZji7Hz3A5nQlFJKixENwSXjjl
6gDPr4d7kzSFNVqNiw+DgaqwXZdCFL263jbnsjV9NPyu6ivOpfX07oaxw0jSx3Hn
7SlVN5EOA9bFtFljbESlLjT/vLSJ+yDoam8TCpaZac8tsRZLBLnfiH/r1e/nY0C/
Fzo+CdJzh3E9qAQT5PJcIsb0Ro8alvS71btOOm6Gr4iUTdvTHSQ5Ug4jkvms1R2K
oDDnHAWBCuBjOcSYCtyKVcNBSHYIj7l5BrBEfKbQ1XMBzwb+UJcBPsBxvBWOr1zH
ed+Hy/A3IJpEpX4HrQam4ecSpP8ZVHljvALoWHrb3qs8jxVHf14LpUHU4tILIqK/
HodisDOCcHlS3Pt2h4kJAW5/Ac0Bw1IDgkYl7U36wORpvrdOcgIdb2sUT/lhd9OJ
9YNLDUdorQ6wOdF39IRXfBGJD+S8jkFErxLO6dUuHZwfgXv4KjuEXRsGmTkYSS2A
5bdX4RMdpomFXp9oSYWdaiL1Ztl5JigzeyDI3hGYK/kNxWudlRsw21WoiLqa0AkY
8FgyLQ+Xp89tJlb/HMaH/dgjDPxDRlLL378Ot7Nbv/v/AkNu4P75ExvxawFWQvP1
4K2Iwn/VlopaopfnLGeq/5sjMcLuGsPLNEdlHOhmxmWCLpIXSGkSXwFkjaknA2rQ
gFwNxo9mwhIwxNNjMN5s5nKOofxYN7aNIGIyE9Gb4XUNyBwdXerI3zX/dFynIL+g
5nfv4HHaER9gtLfOvgJ2X+N35kLaaUCAR7NSmyJbsn/vztoMKaA/PhAzwB0YSKVJ
4R9G8kurplmqtuqAiBcObVYFkLVxPb73IzX/Dv50h0UE6EgNLEtZUr0mdy8mCWqb
hjN8qE1IqI6vIKUi8/G5OidfSHjRGuZcq80Ru4IeQfO0JGrV7jGOgF4nd+/qRFCz
IRZQ2Xl+5uUGJ1QwvsDDRDstgo6AlattReVboMdslqdmhlJE/Th1SUZd77p8UhGP
a6R0iq6HHGBRlIZiViWgXT93qrewZ6HeI/YclfRPNzeCzmEd3L2pczNrB2npwpDY
BS7+QL35LNmjqu10Q7QIapyLwRNUNp+soihhnwAXz6i++jzxdNwjIQ+tw8UzubOK
yJbS68SA7xlLhsGz7GzBq4zJLQtdbmpntHVU7wAPRqhyOKNy3k/XMS/EaMlBqVsk
YYv7HqEESGCdWA4aUDmkkvslc5qfTu0UfeWHDTjJ1iLgBkp8Wsqz0TXDyD3GSPra
9HgSDmbVK1BYZv+NnMAlYb32gB0rd5TMrakU3t2CZFAyfy7XTRdEB6ak2cAFxycJ
rPldJO5xdgGBoI/9V5oD9JoyKicOO8LyMMbYOOxIHexv9fAk6FrrUbUwnPWu7yVS
E4G8AtN9EVbass/+iWDg6kJun0b+TXTT9o0BnUz5zCYcuF0GCJLZHimzGii6PbtV
zHIvbK+Gmc7ScaMgpVUI2AcyOb4CqlNZWLUk/RwRU3Zo5otTwLYw5gD81faIGegs
8YbVp1wepso7Yb7KWQQfcu6WG0LZqIKLOAmYU6GtxRx2HD8jyTDOl6kW+TGEBiGM
rzmi38yTZ6WGMRuDeZUkDwDp0+uhHneYQH3uspmSUUlftMQivKxmga3u8vz48+79
OiXDb6HJ77pRgcNWI2Ad7+XDcpXGmJxm1IhVm/Sr9z3i3najqnOmcpjv4S8fx9qI
gT+kTcPuJ9xCSv9noOlczV94AwU+sw+HiO+n+BbbGlDjYK66trb07bleunhNNgZ2
bo3fqC36Enfci2Mqp8Mut75SPcaMbs50WibAD80P/X1Z31hMM8FemXQAyk0a5cRv
+UBnZXchX8WbERBEkR9I7tY73FSXyy9RJMP4E0h8aGtA8pcp2KNOUB7S7SnOL/91
iMvjCJkUUNYUkrheslZAcChanb7yB6IcU8Z/crpuQXaMOo/l/hekMFSLoG7MPPv6
mmMPTRhVILoNnOkI8TODzzbM5hEFs7h1R4zN7ojisXhvWXEaJ6EHarv30LZPSNWH
szHUQlJbcFBG8P6MPfuy4hckSS9BHkqeE43fW8VIfY0biI/MNniEwFZTlRwrHH87
RlVpBgxi70CnvW7ZkLENnm+7cKsaLL3JkbE22Artano6BaaBxJwgNSBsXuTI1f5k
jxrN8SBZZJN0PL9L5HqWLGVOH1JMjk3qpR666pgioKFdgpM70UIOjg5JfzUldC+T
P3ktIcIYQEFWKlwDAwYLjwPD9gwynlaf0PvD0s649I76RbmB1vgn1Fvuf4i/WKkH
1CYQNdT4+Buf4zbid1dryv7CkAIldGT8bQn/oOelCFw1XGwBJ3TRZKFdi7iZzY2u
xyPPV3ZXtcq995Tf/TbdPSCZ61R4WJll2c9otqNvchUwU1+R7a5REdjlOp3X3W3J
m8iJVckbW9Dnz0rWhOkvdxy35ezzyxrhn1yeq0oiZrfqR8ly4rG6K+lzyYf6JVgL
wW/63Mg5C6jV1nUd61K2YbS4/CW97RwWLFKJUz2zJILmCwRo9gZieDjyHN9Jyn3N
2hZ3xVKTNftK+7mcHYgjtK/o15VOIReZI/xGz60sgd/YIjC3RmpTVix1Uz82sFI4
/hDZZMqtvefXOw6F+iDK9tkc/mwmqmC/treTb1P12BMRGXMsFWWXXFBRm8oDsv+s
/m8tyNctpdGzyHQzRT6cy6JsnciFBNzgIinq1MVgMIh/HoXabUeTIrMOChGVGVGo
NQOKoOvA5RHGq0uUpWPPP7xtWvsVhk0xvLMWcEk5K8mUiow2gkc3kwtv8qFrjnWh
QRXvdSQHPzwhMcqBzGhzFUHmg8mUEGwqgsOdpaAU+kTmpKrggt582E7djfRUXzOr
QspIwYFVSROr1lLTdF5k5w==
`protect END_PROTECTED
