`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNo2EvNoZ5R0Q4AtlLPNlNoClVWO3D25gZlg+6LC9gnUm+qu0MtOea6YmekDzAN+
utojoYkrnc0w5JTXd7u2LZhMKdcStKNuKFKlP4+QUpkNTJ75UXysHmK1qA7ZeI1l
UQe8bn4BKKn3IbFzvul8/7Xgd29MF3fJ7/Ee3ry6bmNZmq6YKxhDrdX8dy9oc3Sa
OZcYIhZZzxCJiuF4jDt+FoEfMO8jvXQH/sFKeOE/ZaXzE2aF7UeoMoIqZnsw7633
og+TmZoAH3hDc19jz4DSp7WB3Vw0sJcJPVgahWuwdNReVFudVRAJlUtnpaWp7R/b
ngE7ABncgnAZ5wxh5+2OmKOpzP1dT/jWkqs5U7exIew9X4fiT/Wu86ZHin41Tpyz
NVtQLJ3OQDb1oy51v6LgTePlONmLHirJAOglwGJsO/WyZoIStFipwwIsDHByCVHe
+XAQ9IwA20Ow02o5344Fyd0NklVglpKHvsKIymZZhuaTQJLEFHPertZhJEPW5rB5
kd9suFdOa07duu9TeHdX+Q==
`protect END_PROTECTED
