`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1QBqjBvRpa4gCPlfie6ukG9LLyyBgpQlHXsgNU/np0nKjn4kJZ0op/U7rXwvG6B
2TEpl4VgI4aMRxgAYpAxmGX9hrfMlIuTAZGhA39dNXOt1hOxZmqaG0fJ9RZdAV3N
4lrdz1NuAi/SPEjA8ryS9l2rIHuUpFBDTs//cR8QfQzkAxbnmHvZjDQcxCnWXs7V
FFyZdHkcHQkljoXKW5566uoWyXzcBmKOwzXqit/5rEBGPsG7pkUukPnEAkU7o+mu
zxIsaCFdW/WHYnBtAhN254UQxB2il6yBG4nlgN5ZWJlq8pcYmwuckjVVKbbggqA+
WFYKZOGeIonXgJwugHhqsJrQUzIZhqqnd4uYqBYUgQDIZaDzk0DZLEa+69e/Miag
f7SZ1wyzV3SgShx3MzdgRYn5wOuFvSUlUzuJTvm6+6AAU/HbnsWcWCqSO3P8exx5
6a9VdUvwPKCq2QGJf6NXJ2QhyrgGb+05Uq8R3CRBPZNgXo2l84i1CJ1uKBSvYD1o
VUW/Hr6SXEXP4qlH39tyh5AVS2YFNdDpAjgAxT6tnmSx829NFNv95DgOEcpZXpgi
XWbuO478FB5TG/mLvWhhseMggmQ5Tcrup1NT2zwi2cA2pcwwa9JtZ6MDZM15kUDf
yBNtCNGuOn0Kt3M9EPJuA9khqRR+eb8dmaDEaE+daBHmeJoqtGzaCVduaVRI50az
E5Xj7Fm20ZUmh7+O/5KDYlllQgN1WCYMq0GpSSL/o8UX2Ix/nBK/7UeA7KzRK4a8
Fz1uMH9PU9tTgqtPOPWcvDuq8Ou1xxI4/BhBLqkB4Y1wJ1cHpCIViRpCfjZqIjjq
YEeyvIvLFPBQyAZDogStkA==
`protect END_PROTECTED
