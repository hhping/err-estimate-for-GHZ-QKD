`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B96FIBc1XfmkcXNFtzWVaU1kVqr91BMWhtB5rDqexxzZKRztTMMUGZaUD4SQvWsb
bp4T6J/f6qTDx1rW0Cd3T9kXz/4vIFY5Azx824vtV6wmOCCq1axaCXDPcsU9DflV
IjkZ0ZvYV0XVrbziku0Nx9ATqd3z2pM6MK17M8WsF6XxC6J5LK581di/8rHJFtxP
mP5nE1MDUmWMAeYGc0Q/M5B/rQvC2F/g6Nqdg5U6sl2XECutJmQU8SgR9B8ndQ2N
0rn0IbsPgrRNpNHv2BiX0W26SySVG+hnWj7WWLnE/rr3lgWsqTeDxvIRO7ROJiv2
6bVyOMD70gr23g7VPtdySm5ZMuLElq4EP0/aSnRWFRpyk+T5w5Cg7E1/iAvs4VF0
tS3DrhXZ0+Fp0+HI+p3zYeBkIxLyR6en7PP2MJJ/+5oRzxSjT0qYp8vVPV/1u1jW
BKh02HY7QPchgxDlVnXhRb04l0tb9Jwc1FU2cFDULClK+3X7fQOD7tlfhj5ntYvU
KcIU0oXD4e1IjNK4/occopPXvLr5ZQBZBocMs1Cqm2Kxl4T/tE68Ddfimi2wNOg6
LqfKQRByzRfDMIBEQTHmR52Q47XN2dtVeapT9xgoVf/kf4OpQkMDgN0xRCH8Dl8W
Fq7U0iE2QgcZSYMmT8iwZ1FHDXE7lKNofjpw7t0gO20N8SYsgRDBjWOcf8c/2/1B
7i29I5+j45ew/aEJ2HQIs6OlkaRj0USqCx1bzGHoEkdBCjBU+Zk382N4T4ruVt0S
6gC0GhA0xmhxFy3WBRCk5NElJMBPEZn1jXDn0YQkbTgXh2Q5An+OhfX0HvdK6t0r
dqrWRL6DveNlXWb5nTuhDncRTW+G4ev+Ba2peM7Yh9TlmTxooanfm8/Vx5qP8ZZj
KU03mG8bCLf0F7Q0Ya/dXA==
`protect END_PROTECTED
