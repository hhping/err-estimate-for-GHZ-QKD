`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJiRPUHpsVuwBr5ygGlZLANxKf/SgiHitQinu1lBR5iUlpcDBlhP0/0UXZtDDqPI
MuRlfxYcf/nYu81DNUgHZ1rgenGJIVwUk94WgNhwgY0s0yvVo2F85k4RqEYaTicp
6dIYkSD/Iym89g5d2YO95m16mM0wOM1PpdXLSFJ65a3UdVsvXbNY1g6hbS9sTEc5
tckRb8KJK8FqDc7nxLtZ38NwiL/sQiU7oBij2fAqvN5IOC8THpQT6m4uz8sVuwML
c5oDzJvTLlqP+vnnxvwmL/y+M9PEW123k6CgGxEAxIBkyxwbOXraANKFM2Z+6Uhg
mWLBpvKsN8+5d0ZmW4uANkRi7ONQz75mDt3Rnfd8N2GKc1qrdw2NtrL6/9eK4Wp7
A+WxJL2XhjXe4c1JPXMlLnJDEizo2u227kxHor+mpYxPTyz8lSI6GUKr8YK8s8Ep
mj47zkUrF9QYLVEneYi9rLG5GTY9/UPV8/Kx6Rn9YTbGW3Fdr+HAJltD9zJZquej
wSi3IXerHdJwEUJ/or7apVQQmo71fh8bpS/ETj/hOsArhZVrQ+bQOetWZWpyVwnB
gYFEIUN1f1SGmpGO/qgkHMFm8kChkH4HNQbg03DBEbkOs57YumeI+cyMnf+n7iJP
DDsiQhoROHeHM7g9B0JtcjOj379hguSr6n7+uv8/LB4O/Kx7cEd45acuGDrtoj1N
FhIep/9GxyhXC5WmGWsCa7L/ivbTCTdR0UcwIBpGm7AqSP7kE3TPfxmRSYzyKn4c
BQCX9sX6ZhVrsEGGe32M9ea2VAPivzpWrOVgA8fB7wkDOdG/xeoYqrk/NbV1LnY4
i8cfKYTEQCkowPLAt42DnU383FCr0dzPls7iaOAJJrnWvPSCIoJuDk3+i5yNKVci
a91bbRgLJQG9Bl//lBkgqEqe8T+rDzP7/YX6Q1wk1En2xrpKzm048BCRYLU3yGb3
uvWlWcssgG21Hf10Nm3PlCw5anZwZ8huqIxmoan+Aaopmh0WxLfdYzj3zloK6C//
uQ5W+5ONCq9M8QvTS2l8hQ6ML7GBE+FF6VAYmpozMBwx8QwgM2JPhC1bL3BC8OWL
pObCGfC/fBgG6Tz00Ci4pOL+1zTaEh4G5vP2FiPxICtBTZdwDtvr8m3kutEI94qa
i629JX3l2ca9SOUX4pdkJH+RK5Z6KRQOKYTuSsQukMA2vl82t7dvMjcNbwgUZEE+
uj/bn/qec4PdODhtEBLED+NzeP82jbYBrdm1b7jk52x8ef3cOjpXGQwMjmZE8Dd2
xOCa9MUrDmzSsmqhM4r59tL0Or+A6cUJyCQnj1JitpfxO7w5nqSbMt1OD1oXwU5D
19cGcIBS5+9pl2dEwm94fJub0M89jkg0joofPrRbtNN3OTFJgirGn4kurJ4XuaC9
w39RkXD5yrTVx/pmsJIKzq8nHW4FmTxOjuJVkcVrwTCY8KpRjgK2tGhioDy03F9S
MqSJQkfzWpVyyOx+hW466Wg+ogR8sTed0UwO4kXwW+pW0psl7BD6i+P6pJS0oQhE
zWYw7XUHMlTDp9fdPbDnepzm8VMoJMUCdcGNsihLZT8BVB2q/NqV3B61el73QC7Q
NgTgPyqMZ8uqmDLNodE1LDyLU4cPzUbZp500GjtEMaQ+wtcsGLi92tvcbVVKV/9h
ErR6GCnWoF3HNzRkp/tQhAPu5zGghJecEKqyFVfLDig4AorxWzdyZCOm6cxLtCpN
F3YPTNoSpSUGncyr0RvUoBXOijJnaG1tuNldpBmbO1cDMj2B2OxJOq8TnW9XbGBF
FYwLu7/l8ZP9mQdvbCxHAIPCq++01fgrYK4mkJvvif1GO1FBIexLQMTcIYaW6QKc
KKDXTZKDwWW1oM3O8XEbnZkMldz934io8a5W05Va0Wt0TJ4dv3lDy6FJn08YU5vh
V4QllWF9bZtWsRxA/qrUYNGGWoFW4WvWIqxss2MI3JJ5ijw6Ptf024AZML5HP7QK
jGMXKp+9FUYZ5ynHxjBMzmuMJx/Dgkg81Js+WvljbffrPHH6KFspJvTzSOx330eT
dvoZwkMuqoPLf9LLOEOcRY5NstOiEZqLpmIYeZdcOctxP04jHZVc58WR1Rmla6+J
fI/52iqQ4YESiigciDax1nisya9FBySv2LvFDHoxM7lu1f6FGwDonyrw/ABOvRL+
DgjABxnmre/npXRaU31Ie9eSZUMwGLv9FxVXPS6gzz1Wsqd9fI+1tBXbMZy73cae
jlWkVcQROknWcuKO8xAzT6lYuAhdk4YA10xbW6gB06VozAJyAUw/Lex0dzrmcrwm
DTa1itbHZNKCTS0BsSBH4ylqpMIa0BnKdlJtXaGtAl/O5MGsMp5H0+joNqs5RbQs
g9LLmmEBREi/yAvJrnfMFVOmDy3xh3Q/+fY0F+jd3oo036yitizjp0qFoZN8yAnd
A+teYEksdtDWjLi4FeKX4eK36JrvxdsnI+UJ6EwY4u7Dd1KyifGenDABRC4RS12a
z32wZHm2oOZuzwnuKNM1hF9qFSKf2zorQrFTiWcWnqIMrKewp6MXL8eCZjvfpRQj
Obamp0AGeWfLCd1NeGOSh+I03uz8bl0V1pZXu7+QHnqCogHWGG/+95GJy17qWZuc
rlW/3BOZEWoYWRz0keZvQmEwC9EaU8byzKwF+sZn6frw1iQvTP0V1CM62OOAS1M8
Lfl2tnVoHpBiGDy7dJqXbQPHS8cBqh8rAgzVAu6BKLKWWY5ChRLTxV5EIdoMNpBW
TwY74+QehhpndZ2SLVmPOD1WDXBm/80SgKtyqj+6ngCHPIDmNZhjFSkkTNSoEJ9f
9VWed8JwnGndCfKco/+NjM01zeP2Aau2ShN97c/VgpRgADemGBYKJ0CjQ8MzrcOE
KnLaJpuvvrmPHaGkjKV9yFMTZpQyNo3KyzAPf5wlfe1Ga/BENrVLZ3qLIZyjSfPv
coQSTVVQJPMV1DAdXW/Gnm9ZL50sZeFiauA8v+As6gzMuJlMEIs4JoJsC76O2rBw
4LmzVGr0iJfUB3wuMVI50N+rjiDc+3IZLC/F+14GG5QxfRBDD8pyq2vxHypjgJeX
2XmwuixHrHBwbFd287mLAtEJaLc/vYEFrd3IxvqWHwk7GY12Yy2oegz7mzRZ7y4P
N0zRI/ipgpK98A5Utgs7Rh7bJCXx/PcFs6UKbsLGsMxGmh+oZ+72Tjyb9Rwui+vN
hmGLhurxXy8FkDwxbK2eLy6nmHkAxeXceotoD2UAdPkPb5HNxFrkPmc+6GJ/TOIk
gzuLaU6a0xu1wDjSgBRMKKnb7aeDApy0IWczX/gK6zCNA+/Sort5CoHHLGepW56Q
ItScT138NJsGMa9kdATRn3dfZ8MAlv8bB7sBzECJzHE2l1qOq1XGj4ArNLQbLSRq
NBKM6XuS9bBobyAuOFF9GTBd69h9MzobzmZW8pTtwv46Y0kfjilEeK4LF3p+bJNI
TQBYa4Jat+x/udxW6qizFAwDyOq6rJA7mL0Bnojoggd+myEFMkKoDUQsv/JPaBSr
P0GydyqR/aAJodYWceSRQ+/nemC9WGl8Geq10bDIz+ECHczgXP1FlhXDMDH238/6
bOidCfrYSmF/IvTLl/c5wG8O5zY7ZqPbhUkG/KgNz6L68lpQUZU5+2SwCYG6TAxj
JSsMgFzEHLWz1fg6a3RpnPlN+iRvliUzJIFU1RkUlfTLEfdjSj2X0wpKbIAEoN0r
wM+qxaHdwthMnL4mtQmQTvJgJ3KPR/5u0fjgKFSdmSYIoCaLbVn27Z5EMTbGz/PM
4HYjZJmxcX7iCGYvCJniWmG+s9iYlM8/AR8dHMHvzunoQoigTGL/hklU/kJxz3Ka
HH3JbSIU6nfau7BD5Vk0z3vAmQEut4CSZT/iPemkRoING6GSGF9MqiliaD9vRvuq
yVYAva8k2AIQ3JBED4XoSltDbC6dntpl1NcJkAg/aKYBc9Upvvnakcz/C9XfXKeU
B1/WvGPzu+KIRZ5BonLXlqvlak0fptTwLAFtkDNeIOoPyoz12uFFvwbSjMYmw9P8
s/hBPQ50qEQDnOIeTZAlydiJUujz/kAxTDF0xG5Q1Q0Q0pDqHSSSHUhCNO5d62KX
OX/RWa5Qg14OzvMMgYB6c+j4NByTeDOqUF4FuDxA+gchscum7X48iP6jZLbo89CH
8p25O2mg1RYKHvEMgt78M0r/QMgThzKvJAFaaQvgKKZZK18TNMg7gwxbWhi0JWnP
vQ2hKksFvYIG8PtMwVuz4CbF87B88HBPehSlfI67vgJWY2HL4Bk+yQ8zp+mCsk0b
XYOBy4k7dXjew1sDjlKtZM6JGyZhhrR8msSVRfcD7z3I3hU3QbGsEjdrR1kMC2TD
Nb+Guu8vGHNVvPrE/Flh4bnZO9iDFRGN0XvSsxSXHgjmfX/yj7aSx3eWt4KZB+2D
Tj+wUwMp9Bgzt33obVJ/rame4jyUMf34mU3ft4EsO6oTKKG6Gqp8ag2MuPNGlJFv
pVyHSF4V7jZXayvy5VH7EMXYnKYJ1xpdYN1z76YKSk2LFjpTXTYZupNRuHmTZZg2
1ZI+G4IpcltYOaYZv+rSJqWuBL3Ou1jHwuIwWij6e8Vw88AJWbrlK0iY21l0jJ+s
dN6TkGc5XzzMA1PVbYWgV/hEr88yS7W8POih33khyrnWrJ5ovYcbEMNKhThFusHo
9Rw+OCDIiHtMIMtMUBO+dyC42SNLrS9F4CsCS1d678II9ZcPFTEgunbPkfXqXYzg
sVkDa1xVzGmHUFmO/lZe0bxTPXIrLe5lU2Rf5l75axpaM3MptNQVqr84qVxIxwrU
bFtHznMwLqdz+vsua9Cwy61v2Rf1xkCWOlUcrGxpgVMnTwojCO0GyCoVtVf2R+fd
zld/Cwe/SLC/VEkXvNH5MYiZnGq6k8RVhG18blznW0LSWw15/51JZmSPRXeS74LY
7uk1T2ItgPPoQRDyW6WwBcVZd7+ctKzZ47SnDaKPggMec1266oQfj4IU7sMqWK1k
jU+eZDKTCnjiz8FTOS90qW6e3ORyBBiFgZmdx0QwsB5xd1FvolcC3z/sAC9G7Fsk
ZL2W47tsdchDCKxiaoXtQV+cgEpYenIQ9fIK5eiBJ6EuHS1utuYsOIMnfEtm0ks6
gHNaYHbAtdM0+O19TVV5W+efu09UzrjJGctk5sKhOW9KiTxqfGG188oOl4rbt8gS
l4CXHII1JFbtz3gir9+zRWbAJzeSP3mWe69WwPkZfLQrDqsfouR8cN6TTHZU/SUY
8hK26Uyc/2Wea/Tw+6nkidTY2LJiemoD1R67jLVBZmJbwZVacsOJFv4VSHJFv8iy
ZxAHrf6QxktPDAKEIfP1mQ7GtE4//C+d0UNEgmLA6OV0dE4zp5sVGKOlx8I46Vq/
2dHWe6zicnkfFLOp/RtH55qzc+CRVGzdveYqPyFK/0fhICIYh0rEW2gRBwISatGj
87a/V/FsZcnGkaE51g0L7fqACdtRRLldvgVgX4xb1HborKalh80vgX6tY2DqVCav
e15t0aBI7VvUyUG6R11XQGjuCmE/FnqFqkcZEvBKn7DRsrEsfc5w5THtO2Jp87Mj
MperoEv60GihnOlUiMMuvsK6nVVZ238NjQ/6ubbfGSPGjM0cWdPOVeIfXmjAZ4IF
1mOFUFWwwPxVW01jhVgz5nF9ctQfnsusqhEDZI6Xgh/jhD9ldtjzyP6R5gPTEoAL
90N5lWtnCmwLIPLAS7reRcTN81jZRRxb6adrvh8xeTlnrMDC8c/orjuIs75PaF2q
0azuRHRGL8CbpAAdwpAWWVVAEH7d1bIcjplBjZf9cOxxEyt3+Ry88AcV1JLb6piV
Sam0dHPDan71AR3HQu8CZmRLmW1Id7D6JavaC8a2JLbeIisseyXHpOEEA4muTNZ1
XwCR/PpBGGa6dZImGKBSTFStpz6XpwsMwa+8MiZzJ3A8yxIS8iB2btfU8tOBf5Qs
PwgLG69Jk1hG0Ygh6vVGqpJEhlct/L79vxR6POMyORxZaTyZI/RTGQp7h+yXNJhg
ZAma2Yh0D6SMV0jFqTjkuqbKT93QyWYLYKgHhjWLw7ufFsCKyVNb8+n7r/ygwXLu
qVw1w7IihcpsBaaf2AVC4OE5na8kMrCwK6MdJCsNUfVUMjjBFgk9XRJaaaj1PFzd
/EhmgxOq+7T7uagsUdXyGqTCHFuan42C1d9RqAgz2px1YKocDlE84amXZX793JyR
esfKZ4BazFwaNpQYvYvfwunRAvp4XttIe27/H5K6n4iXu+RS1y4F6v0WKgjii4lD
KF82DB1e2Mhbcf3d5FCWBAa7+Erory/D2v0IOdRV5tQqaE4zEpSpBvnDROJX66Yg
jINmsw8f5ojrcvXZzvzfGa/BEDde7ZKuwTVwOI2YGdZ3wHP9EeuzPLLzxLcYNAPV
e/kPJ5d/spiFMenrVtzIFnURQ0E1kMmF0Xkpz/aItBHk6g5ElEp5Rjj5XROKirbc
wTBuQa1uDcJIp8VLoQCFPpMJ7FZ1c8ur1iDv7ExeHbHM7k3olBJ0mtSLhJFlYZ6E
EUaR/F1NdIj9Co4iZC1O0af/Y7O28PZhAUIGJEUPPXCocGcfh/fiI767lg40E73Y
LKBCbX/xQiOM7LH6XfNNgrWp5kEjHdepVB0WEfjFJ4CNJpC1itMyy7sZWjBBAlWj
5/wfrVSbt8O5xfckq/50D5TgxsD6ZB+Fwd9kA+PtfgTiHKMcIInVbetrsLk0/lCb
OhRjsCuzzLInnPrwBLIz+OyJlzkeeebIrUV4VeRn5LKZ7FRLe1sIst56B/z/PTST
phJINtOX82bJHJdzhR5N0EIDzFEtJsRrAvICAqeaXcWlGp61pCdN5thmvtI24hZe
kReZy72a+fLs6Jd3EYPG9aiO4AIiWiz5oHb7ZtFb28nGtNIcrRBFlc9EJeij87Ld
z9m10wnokOreNdiemhLI6hJWmYxza9nLaNfzwbmaq1Dew/RENHhVjpsoKDnynwCE
ajZkQ5v3tGxbmUSFw6pE3lST/X7QYmAQMltQfSk6PI2tLqn1RZds4SfscwpXrpz3
0ABpX7KcwCluIKTSPDu7e9Zpag916GXODrT8p9/nKXn3cSdNr0Bm31ac44Vr0o5G
v8lGg0Ilp3Qfzrbj2qbcvXp3Vd4WtkfgGMIgaQC+7T7a6kiY7lXOAexQCwPkaqUA
v0uWiYQOHZrWeEfSUi+vkKYNQ3P8BUtEXpTdZGajHzqhYM3nm9WrknfzDh2ffrNV
olyFR2wQGmICMGGwu2T82UAQa1FrB5XxeIixvdl2JCo2XZj6eqbfSYVWhK/8Oi3e
QW7tGerHJutENZCw+sfNDOWqBhQyT/QFzYSPOueXyODtElykVyySf57OAA8QnkCn
j5GpKZh22pbKCPiLly217H3z1MvrgVENN7UcbtShMLbQeQBbgw3MKlcBje95/MBg
WZ/PqKyvoqFNE1adle1rPPEI0BA2GrOxXJtMk2bw5HidpQ91xyl2gY5WPkPSyl78
wVCc4EynOVvFD8A/y6RR1V5cY/QUym6Zg2S1V9MmCXn1NqwP8szlVytiaEa79u5b
eYMVkJfL5YJAZdxunSc4BaHnVOLso84hI+mfkI7Qb7WNAPass9q7YHjPCDgilXfS
1+Col8DOCFqQKLEkNq5xi334M3CTM76f+KgG9VQoX0yJliCbcIPv/j3DkBp+2JTP
bgyvV3+BDW8K43c5/QDfkz1uQLSPg7T1xGW0K1QTiIDwOeXLZqFT7zodWQfCtZht
jMl9W5nJpwQlWTcQxBKfOKxv7vWxrM4sn/2/5M0sDzzECi9/fJhNFCYgUlu2PSei
ehMKdb4KSqUVkqnD3lkVZ4vAYBRbgCxADNQUXHMvjuw4oOP9VFZ/mFEgNxrUCiG2
ayhaxqQ6xo1epuMlixJ4C2nkWjyWcQYhAUnXLXg+spZ7D6QLSBnr2Odl9n+Kbz51
8uzrl8bGADOyUISm44lXiZExynPyHMXFd2vHLVl3obG0w4Zts/n9GEtTIlri9J0t
zTtQhjnx+X4OLdkj8ZZCP4BwtBNuC1ttDhtmjha/sZoysHk3rFbDE4sGoNRwzjIw
wqkW8Z7OY8bt3ZQrbUlpEaewKwbraBmw9wmTAIFvo0n6DIJzCUmSBzXoufLnkW3x
kN5dLKR96mcTTKTtZDOMNk/5bZxvweWrMGQTv++SxaJpXXQySSeD1rl//drYfTaz
WpyumePPaPUABLCZClsPZVpGY1T1+j5TzV1HQxZrb7P0KlWzKezpkfjMAo1vd4X8
O14SsZxg7DR4y6RjwvN/Wa53eiADOFwCEyGXhEVTT3HHAi1zVWfea4eKi2czWjpc
nMWQkiQ5UsapVFjuznpD/GsUJypC07yflEEIrlvHXqefB2FQQELfawZx61rs/PGi
2AkzxgqpxA3bj9+e0d2bIh1KfiPDhNlFGecpDsY1ellx2FWwrRULjfLed2x/s3MI
OB4bwPPyOdFoemq2SoPW9+lomEZcyKST/+q0PrcIUDgJzxdsG/0zIr+xYVw+kpp7
I2Bb/npSp3ELvM4FjMRzHyLA8tMOjUf/j7avXt4+C7GFoeTV00EAd2BhedGm6+ik
0RYjoT0TxgbBvjodgigpBEw81vWCD0l4nBy+lgLXaIjXdSTI4NDVKMYhULDSdAPP
XItEG3C1cwGna6NDZ+5uT7PPNF05oRzV4M7Hcptj0mBhgpalwEyA0P7Mc8iHn/V+
VhYOT+VAFTuK2CEGu3WjI3y25aHoWiOQ5kq4zZ6q4vKOEwisodvOIgAcMn48pXho
+vzT/ioyrw/jOftokJAxVqtJwV8z+NKgO9/CfiZVnitYla+L3yLFBEgavi8QIaln
5i3rLxtpwPHKdpjXwXgQFDbERtpEiF0oJ8VCKhLbbK14l+fY32NV1xR93tbjxYso
zobWDctZIr6ofr8d4HObFdAVjdN99KzUxK81YHKOks69p29m6STDTMgQCglTIQAm
sfvpCOPhVk7bRO/nG0cjeW0WNKI28lvCOE7ohEXyNCoXqDc9ARCb1g/LH2BX30Zh
w7LzJXfsZE7oRcLp2ia+ByN7WYZ/in1l9A0Muk6CvJPmJothLmXEF3J5GU5FdbHD
SLvm8NnPvLjhcsiR7ez9s8EqnpDIwn2Dw9To8joBdrChnppqM8m6RA0/V/4OmWaS
WptKsJyLxZXvlSj1i1NnO5t1oc76PLSb4z2FmoOb2bGvEctWcw+rsxy0MDpDKJ/B
OxZYI1GjPBpS3v7xLOy6OxFV9ptSJ+017h30895iMY84ZBFmNcycIH2s3dJ1ZJBS
Rv/3uf+Bf4lwy0yPkBOhSRZoBAntpNNhO6uUiOxZs4Q3IpUxRCHobLNv7nKNIvdI
CuJEX9jjLZxxfMeHii6kI0YTVWwgLdGa4o3e7fHZ2ecU6jdEqm8efn+X/9Hdf5PT
ELgnMHmOpxaptqDqKb4qEOBu2xWs0cmla4eTm+swg1wNRwbpqIbPoEBCrZey53dT
/PD32cML2v1bir2LPuKoiJ+bPZCUc1dyNtzXRGRXJx0ActsP0T54OomPU1SLWYIL
seTuAFhJZsIhyX6fo3cA+y4yY9GEmuiD9BWrOy9mKE8QaZjNZx74qP9z65GP8Wv3
jrLNDKtehx1cEM3STbPfl/E2FOgmX1S6JXGtbxZUsuFURUaxW3S5x+qWg9DKJfYt
U9OwB2DLelcSNcAbrtJ3FExHOweD2FruOt6OdyNp+9wiYQL3WLXIEazSHMpU8vCC
YHgIh+Q5p9u4S8sibfMcbmaFc+0Uk2iV72FrCf5V5I9Y9B17fWxHsfd39Glj/DNP
/t9eUS6SHpLMvN028P/2gfK9EftnScGlqAs/LGDyNmG+Fl9IRQaJLoorwvH79bxB
axCAappEGzs5Cd++lKUXlr5rNAlcDJXljwby7hgRDzAkCMGMgMoWal6p/xalfx/p
CxQzzY9KArTvvfimcNa4hSwc7zcwlVruiQeAqqg0tJ9v8AIR78QosENTjr2Q1dDB
QCENdTwcTeliX6/Fue9ftrpSIEAh45DoV1zAfLSWsclsjV+UXmf4iMiKWQC4HYGJ
P4Sp8YsKJwgwlITBTuy7e8ypPGv+zAKM6aoOJEOVk+lOjiXNCWyViYJr0dM4e8UH
hYzJAK7FpQzJWCKqSZ9SokL0lMLPDroScYPvG/Qt1IHMr0aR4w6n0KuPnD9vVFr7
E/sfTFhIUG0x/CdqVeVPJUN8KS/mlQUNyOCITwyBDwRfwHsfSWmhjLKG9HAb7ExR
Tpd/+MEOGVjDhOiPIBVAS9uSm5mcg+YFHwi7CJSAdSirJcqQNBXhHT/lKEhMdx8x
jFedkWt3RA1+o+qIqZ226Q1anflcUxpA+DtkUkcChHLE5VVAR6sQyVUsPmo/nhAi
suXG5hVwx/7J64cmNbCI4iUUGKEab8O1N8fHvR6FkPYpyUvJZ5CbK7cBTdknsJaa
03VhOZH27Kb+jHJMkmvcfNRJb8MwmLLHmQmdRTfbWtnodLtQQuL3qxzzhrTY2iRs
Kk4vrqJRpqTcukmPWd2G8ai2H8vO1BGOw0J3R0w4J8L7ALvT1UROSwHJP9+bAHKy
oL5a9VGa9VevhAhC+EAyRFMTrl+xyejB8lQOpzyLKZ1ikAkleKi2OOs+T6023Z43
c2wJNBg6ire8kL9HZVNtA3odSZ0sDkaXCBbuyCMlwiG2lZDPS7WXIVIHwH/WYQ7n
L46TXY38aWv0JkZnNiMfTaHJIi6IM0zkIwxN/0gr5x0Hi3ym2Txt912bW0PhqxSV
muoakbsJgrp31IJZILgFTXJoQwSlQkbQwzt7C2Y2sEQuknxNFtW4I5q9NZgY5gZU
twdxFGs3BL4qOeZT8PimxALVf9nl7xdpvV/9MnIGfRzm1F43VJlgmeJfNl2PCCTo
o+Fp99nZJFOBydfrW9LXzlss5p+YxDnbWkC+bvGT7kZ6XtGYuBGVlVGcSPViVnNR
E4gPWetYpzFoBSwua/URWS1mO1tv+bIqqBQPyOmGFxWduPG2lDaoSNE5rnUWir1P
bmSRNONtZ6jbbs16oZ09qtwEV3/omWl+2cmQXz2GmKG3Exe/iDtNTIzuFkEaWrcS
P7qRb6z0zh1gTqvrZNovsSF8+zccTq5mgDtvZd0hPytJo0ko3hfUloYu7wYWS2Da
Bpr3a9Ljh9m1AY20Vgl+4uPKLdQi+l9eKEnH/5EzEn6+Iw4tIYGjE0OrQDfFFSxx
jjKYNwu5YJrWOQ5R9MxooQ5DK6s20hxhtkWa/TcJ2072z6ghamG73a9PxmWgaTnT
ghlBXf/bQrM6DAbt2nONJ/x4MurxOgYRpDIdhRlRXOHcs3RueMMdO5BxsITDXgwy
Otrk2G1sTuCgnds0mjznQGJdJg+788mGaaTjtmqQ5wLG6Ho5Jh54jVYUznVe/AA+
LAkG+16glffdn4IS7wR75FhSMbK6u63HIIWS2YM7Io5Qtk/YQXWAwc0cUed1k2TK
0Bva2YI0OYUAYhPHofr8S1IeFXmkEe1thKVKrBvrPBBzP3QHLY9CJbbkhqp+Jhsh
XS2kSrt7OVL0ld1iRQ96NIFSokm/P6ljKM4gNdJ5yrQJH/87K7G8F8nng5Z+eKJW
mji97qiOyCPL/xotH3PWsSkQkDlbVrDQQ9BiMj/WU5QGaRQV0TvSPJ6Kg3ka1K+5
Miy9/ryfredmgHasX5Ukuduu8tyw3U/AgTtdIGRByGpuIX1P/E0L25es4nVhVR+y
XNIdQbr5ZCZaGlAc5xVsWnqWTA56OMC6k+cXMpq21LOlVVKm1K4wPpNJxyC+DsjI
keuYxbj7sa/bOJW8kYuv5Dex7WPmU9JQJ7lGXLj1h09pTtVHkfvIGsa1S1bmn4H9
LtnOt0PbZYxks3iWhWhDp3oh4Ql98BtaOCTZKYrl9/Yt1WbQDGMV9E/Xc6JH6i8K
9pZc5Q+tDMlu4ASZ/bpwqh3Jd1Hj0eBcnkUrFbDIPQ0ffTjGt3F4Vt/KjCNRmmWV
rZMqL5Ki1Oa3oOhsZKrTfbZmvkR3CCmyEnluLHeieuwlhUmgeTO4sCZlCj3+bcuu
aYi0k64diwFT8ZUDOt1P/OFGTg/wqGIpxnXdbutKP4MEc2i5NAv+f4lCjMnKMUun
p8sZg9/MKcNG4zc3iPJpWFFN37NCUP+PNCKyZB3EoUuSInDXJ5sUPX+LyUUl3wuU
xFjzBuHxGEoE6NzwPmHEKImZIucpqX/trlikbHHO41KXCZs2JVGCBFdxPiycEEBJ
U1pMZP7ithzkI9AcOz+Wo/f1VjtS6YfuecWRBv4h42TDFYsTzXuq76YCp93F+eCr
ftoQouTX9EgcvhwIndGFS5xjI5KGRzA/OxKFQP8cTtnnOR8jWzTlMiOEEzUmN6HK
CF5TIUfVS24TeME+uncOFFdJjAniRDcHIdbINTePOykwxLs5cHX0JnYx/1xx1zq/
qeIsANP2FRAoPI5YWtcomhmC46Hp/62jGqhyJZZD5H031K/O0gtg+P0oIhxa1A/w
BOch1+7pW9jVnsHPKIo13hEHmqaa8oEZ1M/lgAeqWbzJnIPvojcrM5PjHdkwouHv
DQDcLHimF+OQppa1C25/KjnJvtEmn5mpiHzQ5U4iOUlQMMHKlyc0WZmbB/5/H8sg
8yYZa2MCACvppRQVZtqckYgcmzID8/82fjtjwET5ZqB2mtXMNGmKWlsEjxbHwlu4
PlHcEKx1THsEtHcbv7QPWG2ciVnlI4aQIhBb22Gn+okwnqlre1gFk+S2gomhkQ5k
zRpiEuR1EUkBZDr89VoDllagNMZHIQlPEu93wXLwa5JvxnO8WiPiEI2OEHw6G5Su
4ztlf9ZWu+h3VgETF8c0w+0a5ePMd9wYA6nTD+NlOubb7QS0a4vy2w8eDmL4kNwo
CAj9otBPZaWcYvd+hAR6xMbUZr/uxwKYUeVMIw2JST5uITJv5bsrGBYujEThwzW9
mFAISMGaSkPhs7sK3XsGWwON+7s5ReyWMN2amtSXY8YlgcUCgbMJDkvKyl/z0Csy
JJ2Fw2HPN+U2ee7UcnmRES+Sgw+A2WTmeEAxwVcZnukqcvhQn39Ar+hiWH+G5WSm
HTARGUV6vSjMMFKa8cZqgJl/Jf+UATIZtqZ00GwMDEQkHHFF421lhqnKI/emfmzv
AMHHZoOAyaZhtyD3R6nArW4ngBQ0xwQTv1ibz/9qto5grt0GBX5wEOjpw6qaP3yV
tqtH0tfANgFaQriu8IpLSC59QyIY7D94OzNG0Ps2iAy70ZayAEPAudrwmxl0q3jy
FsCnD89Ly97OIAhIX2LmKCLRv1NM9we/7I0PDIrKJQCHbIKJ+AZ7vwuCBo48KGTN
QIZwtd58yh9QneT73jHCf3s4kwGRpoD0RtVSaA8Sz1ZLdqNSTcsW/Np9HZG/6j2L
WWGOmLEHvRz9nFZTEpNH+iek1tEXTAYUvcVE5bb8l1pB4H/Vo+oKPMsbCLTihZvz
gpiu05J8fx6VpRYIWYLQg0Ijn7GKRZyLyscH5iSf93uAZEG/XUjAlzHKhfyZCh72
PaGDWG/73pK0hcY7oI/ysiXCSLhhPalvdeqgYzY+BPzFDecVqx1nv9fSoKVcW3bZ
L1HsftsmXooqb1QU4Z7At4VHvaAdgCdLMY7xAmgg+g34d3XThi5t3DZY2lSkny0q
/INiq2AqUVDSwUgYN99acTKDtVXLmijx7A8OU5cQdztq4AyFS8oqnvwPG/Xd1tuJ
JUvgc3AUg/kXGNUwT+xYgOvKpXCee5KfHz2zfcAMmIKDV0QzCg8mVQ7oYCQOCY2O
q3WkViia4komdI9nr+DcUmTTfBwYLmm6XjORBzEkEGHwFzsHacaJ/KBmT7PsucE9
O7+gggOQaBEN8erJUigUTPbwm0WqfFvMgzuEIfdu8gWi0qO+PdVo7gecrK22D40b
b9oh7f5zNdIhEeoHDTgJgXTd00EtGyroye4o8AjWBFOKjTl91TDCkEtIX58i9Qs8
Qo8ELWDk4xSbyc/wSZv+ne1vvP7ElPVhp3YqnaBqrPZ229pn1V1K5OY16BKz9zL5
8wgU0n/uJohjJHBSmQSD4TbICehRZm3HK5liPAsuTllsPt4Amsl//wp+0lXiwfPF
6SItvqhl38D8FDGXGHCLH7n2fFWCGw0tSKBH6+wahUNb/7LrH6jua6K3vLarMKYZ
O1RhmjhOSrU8j5/sMfo5gE1Zan/NNkAwHluFdK4r0mbcSBb1AkhWJzubGcTL6Ub2
IAPdAHcHIDZah1FW+IbrlQ3wX1Ax4xh62eX+Scv/i0jtG8pYaMNmXXbYzmOOOhfi
VGeGR3s0atNnMisryLYO7++X1njAPDJaoIozUgZZAqbktTyjBv5LFR9NENANvss5
FDrW0khvCJi6ufbSatM3ZRoz2SiEQz3LCbDku+ysczzepUP/KuN6F3CuD22VGlpp
y9LfG60Nod2p2Dk7pDMK8vRQnVLUCnEuFrfoENV3nICsFwSYdcnFkaRWiYtjOlU8
qaIZXjtNhuvfqC9vni8wCd2/L/Lu13vx7XR6NLMO9ZLmsOwmI68Ct/ylgk06ufqM
24lEZbGOt4VVUuzY9Tr7AMcQNwXBvlKGnzrVCes0JoqHrxiT7q8V12CYEbREJB82
uqEQrW3gmzskEcBITXuxFGjolxhUNenOoR15/cVMSpGT+2+Gm76oc4fvxKO8sVEN
/Oq6wp/gNbPCV6A/lPfZnIZAY3i3L+XCmkzhWNUmc7egfhFiOloazWT0b9DXuJs6
/XLlJagOphhJhESBREzlOonimue6IyARfCs+ZmQqVcoxc9P0MPgisQYBbSE0nF0A
/o2OHoI/VAu4Br6BKHVLIRKLSC4FLFZzSclRbEtUp7wdv5mO2SZAfxTHJXtABzW+
eGBbv0uGi6+3urntXUdqFzwbfMRGZyLUBkXe6ajnaqUJIPIF8YFcLBS6rWX8/35n
w5UVtssoqGx2GCIGiLoCJbW61G1C/aOZQqBr3uLwvnbXoEi1i0AieH3kjj7Zls7G
xZs7lA8jGjzLu6lUGSK8Y6JHonbwomDGbTib1bVi0ah0vBzp0KxzJs/PXRzVRiW4
ZTxQJwNs5l6bE/qgqVn9QzYEHOPvO4OUqYvcUZuVsdAaN5jtUDR6DCPzWA+vLucW
Zj7+mg7iX/8Lqy4FHc1Cj5vZq2CJCyk4Zr3W8EXhJryEL2PXUsAb1O+e0eMdxkaa
uP82ZOSam8dhrya7lBC5h8pQ19Ffg441DMjaHf64GsTA5L0lJULiyyseO9C1IxmJ
78+uqUF/LUODMEnfHGelV/xdnuFCAqmW8bsTGWCvCGjBA3vCQzT79BG4LOnkDnEI
s9nAHxwhv9s4tAL1or78vWkm5xYmt2rAT0t+Kbz+5wNG1mDymmUyYpZ3JAU6QD72
Jtjj66BKCUFl69mZoDmDF6swJpYKZP0Xi5Ii2NS+1jkhqg8aIyBSKMiBgTuv4chT
0uIlE9Fi8T/hgO62izkUdcNrAc2kAfeh7+6wCNKOAVw5AZY/pXsutOH/TbrsSOdA
GuTvnPssVXz28JpFz7H5NfZEUTvYFVBK4nIcZdsscTuCX77egdltaF0Qb2YsDPrT
DT53xbvtPenFCODH02hdkAbxf+kEaWTQgvyXPqo1IBkP8oqYK6+iaoQYaNaEsZsp
Fmf+4eXQOsXhj/QB0VwJ9dqDd8hSHCkEMCCBYT4Jml3AJVhnMzGD9PAZz1C9AD4p
1XurXAaOYCbxdx+k+3gRO0zOrfFLzQqkwwJMRF1Adx1vwyOa1oVNoeBT8TxnKc2w
8x1pNbqFiyFIaciNKH8gvfhFciLSQ0+8VkVUKaf5PwslBSyeywUltaJY5HpMdZ0I
H37InHDpuwnxAOzLD/zWQxzLu7HaczXKPTfQvJmhU9SEx9UP6NXdffv7iUfR0SK7
ITbfAgh3t7GbzXrxuxFmLod5sx+gjN8QnvZoKKHBOjS2tvWiaijzuJUYSUbUviN7
0y2hb1/fVMmp6kkAH0+v3YxoCkle5SVBuJIPVH/B/o/JCb28mw1PqVGIQe4uBgKW
UYaErzVet+Ubb5mQIt+l9RjYd4dSOeBL2KpRB7OxJTI=
`protect END_PROTECTED
