`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TH8vUa2Bs+KNbX2XRhAA0wvHDR6Qu9r5oFXej273ifp0T2SloKvBoR02lEDjgzS3
w1FaekI+1p+As3lhaHcijv3bZxWBgQUqnBnUXZHJ4iVcJlu1A6dYzabLAy3T1brp
AhIGjTGoMCZs3HS3xjaR2Em4ag+vULryUgoDTBcCKm4yF4M3gEqploxCEdvyDVb+
IZD9kG2p5muv0Sz7wFyUvy+PKaGP/DGl+uD3th3YL9P/zfRNIBispsVFskCIyc5p
qwjSTe9pCn8q7OWq4Ivdq68j9g6KZin/GOwoi9rnefWg2Bn1YwELlMwqU1Htzrip
K/zwluyf1oqWDUL/x97g4jQRvMKz3AWMr0wLVpHthqLRn6c5V62z2cSDlMUsaPcr
Dtg/+sIocmuZWzgHQoO4/+oFveiCewJ8fMheMucE4PbUilSv1UenplObzuqVo30+
35yTowL7O96sCeErZ+4bwkHk54GtMWNnAqlH2RdeQsslOobmcdPNDAjcVFsEKrWW
XRhHuvhsGdwYgSUEPiuicYdDyds269GHeNg4UAhzfjIcclB9P5teSGvpMYAGIoQ6
O+XxwiIwGD0Iyt4vRcgr0+upFc+16Yx5ozdhyCoSLJnmFqQ7VDtXykUwaeXKlI7I
L1tQf57Tuzq+IG1m+QyWjqAuBuF+j0wm5HomGBKNuc2klFFKaNuUBrIat/eiar9w
nKtRFpvNisLIgvKlS6Zzlhl5hEVfXy4tEQChE09E28dncGn7w6372jjdxR8d2Bni
lbE3XyUAIn/nRCQYMv8lCAEF//+ttul65YUe43SgmIxTfOmvJCNqY5eMGQ/Sgmve
jt9u2FUyjmYeBgvShiBQ5YvnWFyaMNy5GB4T2XHqHOHmlG6iXLclCliGr0Z/PG+t
ztKiSFRo6mXRJaWTzzAUmfGDH6JPK/q/SXaWsaqz4/Fugzm2l/Vx36pBPPjGO9rp
h4+pYJ2tYYNvuCSWVlPAWkhxooIi34YJKzZGWYPj7451wevq6CrmnMislU7+VueF
lBpcAOnkkIHpStHKeUC07GjgUvzgWRLo0KIFvdh2avOx1+Lr9gSVy4+VzKr0n5D5
NVa95JYK3waJ4f0IP5JO5CFo+WMQPS+bUw+3On/+JpWwu3W41uGGBfKenhEumTmq
lj9oLIKDVpUEa2Y0bZBaifT2cGffhUbrOXvgofLNwD01Q6kiVA4lckelpCWHvCO4
QsMaZ8sIV26dE4hXAOEDJ+VqWagdI6EL9godqchnWiCoJRPcFVrQjtLNL/Co5loY
mq96KKGuaSCejdQoe13l1g==
`protect END_PROTECTED
