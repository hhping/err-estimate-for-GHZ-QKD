`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+nnVfg+TriRvQRBAT4AeZ8MMhi7oWqM0LCj3lSxf3s8liO6GFL0Z+68LBDEhu69
RcwsUuJbzuPSjAvRm6zGdIbpN3GyojlLx4hNU+J8oBL6DwyhTIWbtHZzp99y1Etv
RnKqCBaW8XMGWy2clqC/zLJeYRPAex0qUb+MOjRJV/vF13MVrK85wEF9npgfZ2mM
Qnxo1wGbh6PCzArTL/1U8tL6AjvhfK40E/HTq6K3ThlS73HF/fGCIwA0o72pkRBg
oCXcK3WppU5bhuNpW2TgsfIOiNLAbVZtFBvW8wi0/T5SNRF0stUubEn1Owb7IUBh
sgTYShxeI1kjWd8DV8caBlLY9qMur9e33LUg6R6ZwSGwZFAr0GKiM07qzoR+Xy4R
7Z9btC3HG4yF7GJSlR/RCQ7z8iVtZX0wEshpF/Y3kCY5/1Pdpr+nuVRj8O5mjrrN
4k6t6HTltR0s6xiUEFNjzEr0FiePy2EPHTukMOyC/qDZ7izUY684xdCkdvkBtbVV
SZl03gOAm+cHt3XM/7KfehWm0UJ8yqxd1Mel4ZOsgo2PSziT8MzRgoXB4pz8GxaQ
0R96smITf2w3b0Vvgx1qfiSXnizqfrzu1H2frg61UET7cjx2ODnpA7S1ZQqQAAkA
YrOlMU/YsxGVXOwopmLJwng0VVTltgb8aihuYdL0UWM3dqj5hmDPkLye8II4gHh0
`protect END_PROTECTED
