`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RS0qFnuTiiVUDjyIFiksWZs35MO4hbdzwTISUNlSfTkGFBSeB3Qgh4UhLofNrag8
2DybnHbdJS0KU1cxEsqdXo50MXKEWROYrwWz6wmDnKLj/gzy2TU+GAQEH6czLJAO
vrzp1bb30B+QUWsv7VZL9J1n/IR3gEJLEY2FxeJrEudCHdLe2jDM8bqcChY+szur
+WWzZwMF8TgUltoti2SE9KUHdLv60cYGHAWQZ8QbGPWdGquyBd1QXH73VidaKwTX
AinxkaKGzvYYBUw6Vaam2EiJVuwZizgtK2TqYAtK2jTj9WoHQco282Db+kQgzmIR
RpVd0LF+xLh1BrTmdwt/AkeUn6SwXV1aiiqAGy4gYhrWZgQ63K0QcoetyFdjr9Fg
nD/xiOdG6xNIRQTAxA9NSpin77CnVn/jfCRtoFTXp49vLkoV7CMAfJHWtTcrqppg
P2ZBsCe7c3c+eEhdyrcaZr88iOdeky/ADQUoQaGJGNqyAMymj/3onhD6bnJuydum
5M8aKDvql0wN8/dvfEd9DuNdd25dr1Z9kdWWDJTOSA4g2FeViJ4KKrSruHT1OhKc
dQJ753c+AWx+aNvE7ZGRY81s387NTvS0upDuePvZgFjczKDiXLZaqqONeAGStrP3
dbt2W3ZIbr2egOsSOk5l3Sq5+0Pr0g0BDMMnsHZ+p3W6hqeGYd9qgumYRQBVCbJo
LCtc8nAubEPOtYP/T8A2C/d6eQHc/1f58nXdtN8thH7xGAb53CACBIrqwnlCyfxY
YumS3+ZbT2tx5QyzYr438hb1BIDUIwdv4f4HVO+Vs5ax3KGyxop+N1GQNDj9l56g
dPnpoUmnjRrY8Gjcoc6rQ1m44mh6MRXM+K66sdrzGHFBTOxMF/7/ZoJaQb6PaA4s
DTn8L4f9pVHmvYD1gEz3o6J4wLr0ifQ3eP72zSXI0g7/0HByZz22STpr/9+Tw76O
NqJTbVTnqEt3Zr89GZFWSkC05e3IAaseX37tDGOhtYt3bw1aKRO0fNcWgKnQDHoI
Ui/bXLFTStC71lZRvffcCkpR2OQ+MI2v6ws6zcQ6lMYyqjlLFadsSvX4aUsDAqBD
ypw2VCLHxTzZNuJ3Gy8C5F7zzDr2fPum26DUMmcZadUNGYw4bIKf3o2pIJsaaGKt
kXGg+UqYO0bTa+Ifozx4GXmN+S+o9la5lYdTCXE5KEv5ZW7u6MFXmujY1EpR0jrG
PWIGQHNQDTrI1k/G+uIu0Ow8700gfxcowudaZ1Q3BY1gUgksk1F78el/ibU0gAiY
bFGzt0GbUeiUjmo7BAndu3IAzi0bxGuTn4Q7+Iavt332MxzAxDTSgxt7mujkiwDB
I8oxIIX906YXH9yk3zjWms0iZ7hfGYB6UTSqMR59wh32h2hzmWr8Fw/JRnSnNBiV
YmIhk+8/azwc3+7qlyFrg4P/OKUTJtvhRNuEyaA40MO8/SDExzi9sNsDKMTZj3ZR
1BwgArxmYzuxe9RzVDCqw+DJVnQauh81kfemFRdRoSGu/xmKlS4cSz3a/G2vuZjU
hvpM//OulL4xjVAiJK2qrqrpt8NfLvUhVnAoSxs298NDKVn8ZUI23aSGRVF1cvCC
Tjs0olYd1I6qhKEWMFOLpqjY5bHEWm8nu5zO1n9y+WU5r6ij4I0T+8YTLtyfMqfW
3MdnOd3iq64hJy9iaDXvLbjj/8PC+fi4y34VYC4DeiBS0waXD4iUeoCEJPm/0JK6
C4UKgEEkZvUHtn4e9AFOZkEgUIQKCEmC5eTYoBdhXRYiGWZmqRECASpJTTwMsODT
t8FK6cMuf+vxY97q7L6u2ffr5SG7ZTXlYszlefuXWPVPE0BZlVsxEfDJiTYYTbuu
Q+kDA0PLKEkUVxX8dKw2e1DG3GciZYJcjxdgsL/9m1Pv0z8ArcUdeV7EofZvrOnI
MWpgxamyEa9NC200GN3x7Q==
`protect END_PROTECTED
