`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/AvCelwChSx5g8mf1x5/ITDm+G4kuJB48YRVT0E+fzXUfK1OZ69CDfDr+/mciZ3r
0Pont+5NGEM1NEx184UVNZ+ekHZqIsH+sgWCJgvJgPHG9oWOA8kbAxYHDDaszcqD
9TfIleNdw6FSX7kQ9NnZk2YFRdx3n6V81pxULS2+bTw/35jPjwaunx/KA1flcepx
RMEEDDITPOHFdBwVM0O9miHk4tYjSdLJ03M8iPjh6uKtCxB6PPmwI/ymj631XAdN
04Gd8DY76NyP8NUgyfBhKsVEpRMhi1aWy6EQMpiyFDzImeLsRqJepZd8u3qlQJw+
PCHRFTFbfifBJE9yFGIvVxCuSjc3gUIrGHXfpaYXoktOkLsSceNxpA3HWoHPW6R7
LM0+N1qOKRy1TA7cRZMzNOkESoPmUhJGLQQwPNAWMYv6yX1+Fl7V+UObnqM1Wns9
kP96nVaSsECq2UJQ6CHjdWFQ8bTX5Ws1mxZcSqiCJ2YKBDrK6ohJFS6Vqx+Kqq4g
1Oozp1GZxf1Xva3tVhSI8N0nA+Lvtz19+oBYtOTsb+UgslrEpH2jRnS45dU6p0fe
gtKAGjV8jEncqlmnIEghj+NdY6hhsQjsoSAw9m6HNkq0Po7N1d1BJS2uShPlVvHB
AV3/dkw/cFdcRVGxAsKwNrDABr32VAICEynyFKHfJB887ay3VpHDK3j95ZYxA92S
JfSI18UuY4x4N9xbjUyESmsMfYGkMSwq6xaTwhZtwqo6ES6OMdNKgeeJmH0efttq
FUBZv0L3MyVsvcCuemaAH4UJAcIs2KBRHjMHnFFmRlGIc7cyRLtk/OZnhlupHCUj
/Al3nynqERMiC6I7vWgliuuHCUVz6pOah7EKCaexDBjOXybsmwnTVc0h9SCF4omc
0aiBd2VE7I7ywuf50eZlF83/lPWo6D+m8z9W87Ew5r8cKTQbGqfasr7a7J69khtm
M4fIEUNB56D6IJBBwhRmSg==
`protect END_PROTECTED
