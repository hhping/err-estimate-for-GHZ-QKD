`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YKQV3YqnJfgVH4c1atuaBI6AASMVp4HtqChv8EutUHb+KbNlhI52hRa+bYplppaJ
W21O8fjztOj0fMd3JHv1TlI+lItgb54YvB/wTxAr2fqL4ZIPuWHY3chFAK/9oucZ
U2e0561kww1dhiA/VjtBO60y8fYhXXn5fv7vHMgNpiQKuMRLsYgjdv5d4qeoDbhI
ZNe93gCeZddSOijawARImR8jaXBdhw26IASKAHGvld6Uh3/L0xlPnjmFt19NgpSu
jBppVa8RvBFKxgDNHvs286ZLQkTYkfOWzum5bN5LvA5lATCew+3L4/+7hWkbte46
Xnh/UIJFEIg4g+hYt9HC76p7webydwTLWLXEXzPg/x1yjde36QN6uFql+muJfVmu
zDyHwTqkZBEuP6EQRIz+f4kxrEUviEqysLMLq4bjXIKp2kU8+5pg2sBVySn5FzF+
2tPGKPe9LRyFNyVcRal7n4y40rInbh9Bi2Up75GjLprh5OFVe5Fa4D6acBV0Sk0X
`protect END_PROTECTED
