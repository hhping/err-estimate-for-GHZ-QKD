`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7bSmkQw+W1RwM6p/9BJ6IOifG407MjsbBO9q35iqzU+ezXY4Gyteq2gW/mF+7KGf
yGdq3Yr9Z84hMmQ1YqZbDIoS0ONqekv1t+PLgvn/NcpgtIJh+tvta++v9zrW7gJH
LMvXtvNVPuvjOfjrtsbprIVorHHC/YVhK4TqDxMKcfGwx/MPvnYezld9c2wiPiQA
VQyyWwIcdkgQaRcq4XVmVklAfX0CRQcxfdd3b6M4blt9Ke4cwbfWEqLgBKbVk5gi
1emQ0kl/BvFvO8HkmX7WnuTqM/I2gLjhkDhKOxXNvCAfOW/Qx0KHAfFEtj5jtVmj
cxmoWU4Opt25PTECPbC/kR3Vc9KzS27ggBRuXnTY6yIkGGPbt049XxnZdVJCMpi+
l22jkjy3aLQk2uhhBylpNVXiyevbZlQH3cZvprOANO2eys7okWkEU6QjaxQyyErP
d1KtVgCHZZPyEwaz/ZaFZJx79P/b3eXAdsgIk8PJi8VimKU6qdw6H9HrpQRbQGWN
a6oC+qdTr/avM658wfeRXBV9pDzhr+rLaCBm7+iSwRWls5GgNOG5s1Wh6ZFDvF7u
xGnXUjEv2sHRBTxSMRYfs55DvXZzja4Xr1kcTkWh6Om8oyvAlU9Sz9uajJ4JnZop
7aS9vzzul5xAcAbV5dWxQ408WjnD06UYa3hwNxv8qXSYEzpbp417lttWV5YH5/wL
BadSnBQ2Yfu4yI442v/RNt//ltybE0tfBGfwI4YjKFTEhL3+xQqicL3beJKHWhz7
Gm+s2yuKKcUqvXZsLE5ix2znlTqNNkISGWFfeHFJc0C0IOMaXh07Akg3iWqcIf66
nv/ZoNrqLvMz6hk1EWW+d/flN7tsEX7TSrR4AztGlshTKOnsDURMprLrJCvyFa+Y
oWXn2vVgg2ja5dCsuGUu6M/q5+rpuYgD7jVqJUTFyJ7ql+Wfh5dtOa2iP4WJbp4h
LLUaeBz/G7Hin/S7i7rTH4GqCANLmlvyrMUOoP3h0iRm0tEh4H3SL+OB/bLZFeYR
hy5jTHQO4hxBq76CejzrXzY3t1bZ6+ODn7+XyYwFVxodKO4Y/HmrLHhDlJwlbWWO
dNj+wrH4/lunp0qI8QMtJjg0jx3Y7/amUiqEqmLkclbjw4zjSD9M/58p4nBU+E87
UbFaO2THAUMF6u/C9mCmPh3GclrfTakKvQ60zxwmRd8PCcFmAN96ZgJK4hht5g0O
e0Sc3wdPf5GldFHjq0seuwwQYsf22NQ5Dormo9YDk4/GCDn6kxHw33iBMkEdF1YC
jp10MSdK7T3+6LjzeAQWQ9XgphfOr+zI2nIqznrp9g7iWhM5JXNo4a/LPIQopdVi
MgXnvjSv1qfmgE2A01HqUbwAHyHjJ1qSOst2hNmQ8lMLaQgOxU8NdvYA3iQzRA9U
rEvlI9QYfzwDBNEfKg0jW8bZKuww61HyhfQQUV6EPSC1FP2XsaXW7xClyoZf5JR1
GPG86VTs2iCCapgsXwCXDIdVpjV2qZPzPEnnjSQSgsdtNuBi+HGCoUlIscPAVe53
4GhdjWnBLUKX0ImdF8PH6iehFain81BUBKG1cerUbY66nNGTWc6HP+HIH89p6Q/Y
N9hx/E4irmAMr77BxC0A0yDnCSR537KhtlQ5/8XIKGlEXz/PkW0/I52Z7R2wCdzO
uxdkUGATBIoRxNJZytso1n/Ea2BVTCndTcdjCxwGJh7dNfp91T9c611oU/hS+IfM
cJyt2CXkPcAhH+3P26Ab06k4aEdKuADMp2v+BnuXJoapQZGTp84aBq1UyJCud1zd
9HfLVDClo+5686qMAjXBAFfMvS/Kdr9H4D5Q0phrZPUIl8/tMCvRwRiFR/KXURkw
Zz645lLB9ZZFA/T305hLOM20GAY/JiPuA3p00FHzHh8ww/gBXjR1iNIQiKGuLFcj
rp6cbUoiFsZLwNCmozSqewgfseIDPzBH6ZNpatTYiuRIY7WyeUcsEpO7ADatQvAF
hkCXHBY4xvE1gcBIZ4CqrE+GDM7zcj6mLw9+1ngPYgmS+UQwiaEsiGUQSaGO39Xu
aCOYb0E448p7iy3Vy7zQ3Q57W+7/f0msi8caqtd69etpSurU6+JY4IezgeqfaWJw
i9s0aEG9PORtHUKqYJxW0B1J5l/hoy0KikMVGOHAyHZYLk1u64ObKyCvIuWjK91u
yqxihXuqx9S5+MWb6PsJ0dipE6VbbKc85crCN0kCO/YR2GHpjepOQRWWAOkrjJd1
BrdhV9YxyOgfewtFxkwoelZV6LgtduOAV04XH2OUIwRb5hyDq7Zs8PAbUiFXlDED
LEry7brUycYU7FnIvwGAujX8bH6/MTjCgyLNpPat3E7q8PEcPYbYljB4grMFR8mZ
fAh/DMPR3KK5QnTm7ynHe8xS3XWb4hmYDgnsSRK8cV9fIVX4qlrCqQR6zORuY2v3
y6s4GPTfa/18e4Zbu0t8wN5VxApWu7By8tzo7fhcc7RqllAhM9oK5yhbR7deitnP
CR+n+bYWkMqD4N3Ad+jfRChCSGf89m1B937jNcvhj8iAWobDZauuAO8bCd0SfuEA
Jw7hpLYtWD/WH7aIXk/7BiyJx8deMzomYdPYW1Wc7DlWlvUbaMn1pKV49xSAv9XA
Tyjrf+HR9hWe1rEFf67q061TH7hal3KRQmP1CqDmFrjOSa+Iye3zk/oMd6FTr5V0
XyOini+u+15RPXVAABQWhnbeASqQZIq0z6NFLX6ZbVgfvCPkoer8zNsYHKYvfFN2
RI/xqCiBIUSTfSaRxNfx0aUyHbtuK9LR+oQfoFOCVuxra1tHtsXU0NRfw9vaOOed
aMHsLXd8pDjRFtewD1q5FC+MhG/+rtB1XNnT9C4SzMmHiYPR7CXojlAUFej8AeAo
r4iDx27goVbdQYgsKomcbkA7qi/yuDF49Q0BW6tSr8zHxeG/IIYe0p0xwUqNR2hr
+AQwQQ9pr1X3/SxteW1A65zPHWjZM9rnADt3Tux7PfUTQbXUml3HHPmhbsHYXHPf
YHjKWNwZ5HOoW2su1+a/PciPE3zX/JRUtB6fGMeZvajBXQx1GK+homNIaO1L0DiN
gdo4OK+0hHKe5GlXWR9FxBHd8JqfinZBIDy3qNdprJsniIzdyHBSNC82FvUcIFzy
omkzYKU2dUl076SVcfpmH24+O4A+Ya/MiUgN8KkJu0O84Jbzubrjd8M3kod2gLpP
wmJqxqYDaJ/6uKFR7FwSeOqLy1luRPoU+bTZuFM3dgv0C2+eTKGiyU6QnYSYeksy
w7Y0DKVVCExUbBKxofHlx7w68EdP4OQn5W1qgOKXKgttnckGUmYzNetoYh755xEf
rKay8UYIJ/dZZbtLOxccnLM8/rgZC7wRexk4CINKKggFkusP0ThgVMjHIPYMp7IH
aO0hqOW26nObMbBw3fODR/eqVNvElcMhfOF7RVCZ7gzpxbhCZX1Y1xFtPg53kUSN
4um2jlIEjnx5nMVO3mCVcZ7jSd36r7Zx0wvGWkxAVIQskHNGSR4WGPJthV2ALRAH
KncX60r+QYLwMxAlMerQeoQ1oprO7DD63m0M0HHYYGjG6HiuSeoiXMKhRtslEUfa
42rqzIGJ22a9UQ0DJ+MHaDjYzUluNQNf6QvysvAl6O44XWVGzAoKPTtJCXaltT/S
19VlneLcmG/oI6YhCKP6HwBHSMz4hrZB2fVBmFDzDkIGKzQRxZ7DyRgz/EtSg3p9
+l7q8k7lJ9Nkf1CcPlK9hlkGm4bBhwJx0zpjCqcuvDlxlVhOQHEIHhPqYGPWhfOr
WGt4fBO1AwpiwqD8VX4MtF2AVZJdjZnIpXJ2QaN0Y8dyfwLWt7wf9RSDxVPGLzXV
bdL/l41fQFo5WqdaGmbhjQ+v4zYv+PWFrJJP2x5naHpGtnDDL947T6H9lANjt2/0
GeH+Qr7K938ufexxVYTf+pZWZbEi5ZiUF0jx2MMvaIeafECSqCapv0tnd7yGdkwo
hXF1o88HZWw8GLrcnmpy4bbcd6aWOrUL//hmEea66uh8WIwBOepi5WIuVSkBFLuH
oR3qE25XqZbhwHUnu9Mw7elLV8MzfFsakOXh3khaKRSJvkkLGn1HNLxYodPBFxxS
UtaciE20O3r6W4xb9X2HQRnOn+kzFT1B23sy9z6i+NVHjrEWFXgPX9/8gdmQRD9V
taFhqFXIxcTpJmC0fRD+9lLyjXF/JL0atfz1CaG3sl2oH1DwaZPtd+NegeedPt7F
mceMwtLoK1gidNd8NZ7j5ChO5ztiXDP9VUbWlc2i4IZJbX66kuXDMFFxXDJefxyf
aI9qNbjrL/QBB4urUOglYqsq7LdOuaDHli26C70k+jHI481T8R1D38ldm36ninKC
nZJcs185tirGwQy6UkLTBuRhVWsjmQIEk9C87xU/faAHPQoBCsKObTC92DqBHU2f
vP2gKMcw9rLMKdnNmSBvazhwvpxp/0tSL/JHQf7W04PrZlYiQIiWPTQLM2BvK6uU
YKRAcxkCSBRhvtQKutdUxEAkUkYz1kcfmQHXigK4i2y6am0dCySKuICs2rp/kMgz
sPjBNRfFs7TUAV+PixSmImjj8fahilT2CfENVLbWGaf6N4uwfOiiTlgb8Qgey3xx
sYwxEskOsGz1Z+s8hw0Rj1tGzo+grorF36GowYXnzouGKf+oGcBxqsp9zhHU5IoA
LB1ezv0WUHTnF7w+Fa2KniyD0oxPIfyu4NIzOeQ1KxAqL/kDO5rgQofh11a1rndB
rmKi9YuX/YaS22iD9mPnUo4vnbn9GIkqqZnG7RB15wswQsM6ZvFvhXGL6UBMrLaU
INQYVRb+YpB0j8qZcNbsIleoMdmjznkrR3nR13s8RzL5uitzqTRsvhNZUBtyuP3q
ED+NZlbP70oDo//o8z+pRK7KUHfxD+F3jt0kiYlgUXpqW5vIPK1pCa/fL/Yh3Gj8
Gt0gWINb5uug2u08/jSfmk+prNFYDF+09EEI3iPbwlcXnDtrdAn9D/TzEYxviXAl
nPItDcBRhZqPzF7KYSzgfJQNlkShBpz9J3A2G5+YufYJ9od8o+fJxgEjD1PYa1Mj
BSN3LUdTe5mtwkNc/gIZizi0bQfdytqZWpfuAnifGn+T7ToxSmB4Q0iYzeGslbPU
yrQRFv+WFf6nvWtpcQpjrITsDlbX3SrsoDh06fS/YMmtUPizYxbdv40rHoY2j4Bh
l+DlW/RKuCNHFV06Wb904Kz7wTCZBNzV1q9SLDLf/KLWEeMadbPNYwfcG7iLaaC8
hr4GU7eHHROQ5G8sVS1pHmcAcue/k7Jd6mlTb3ODBAVcXwsex5KQdjxy/qvyRJzd
pzUO6Dqvo143/JhRESx7NyNYgaoR5N95JbRFgfJh+uu5/Jw4+FaSfSoK423kIzva
jUiv2NmikmWmAqgNK0/5RSSBvEPKgpreApJacE0mZA6t81iO/7uSQB22g79cIgiz
Z65b5Xta2hclHKq9MHfQEL488l7kHyjHBFg0n126EyGrlitql/ef6U3jigYLgCIv
H31Rh/fTj0chrLGZ5PPe8s6wgTkdZ3PAyN6bFe+IEL3qGkROYUvZTpx2XxC8AgQo
qwGodhMxGrav5pmGtbjXzsyScnTSu223TgmQgkdDqqFA2Sxs3LFKdJxsBGG6fA+D
LwB6LtOu1FYewaJPYlkDNYf9vwDd4dA+0TMwu0gzhC1FGqLa1zTOwQ2W9gH0ilX/
x0Cm/6Zz0A3vl4TAOh/sSX5aK0qfpRGOQ19OJnAGwebTDdiFTneVac5/eHGdTqXH
UP6tDo0IUVmZV9Sze9zg2fXgKod6Bdef1ubkUK/+oS5D6S0mYjPJu0K4hbQbJoCi
vd9eVfwolvASwZfiV4GlrdprWbVM0B98D+OgAc1yebXhaQvIwrAXfbtSQ6L4dxyc
s6L0ty4vcpixwrJj/gjgK6nXu+Lx8Ky/mbT27FcN4hFhqVyiaChGZtxbt30q5wIt
hQ/B+RR6odbouyPrWDbWHRYcNytWb85N1Mkd5FGTRumrzHmxeWNrUBmTd5Yn+ZHk
EJ/y90PYXO4hx5JTz9VU/WKM2GwUqDgK2bGxzDT945qkTr80iSMgkmBY/Qvk+iII
tPRMuSZMRTEhhfv+k7C+ukYaDcE/VSlKVwZM/WyomUPgAkPOQmHuovmcaNSviBj1
96dLBDXuTCP5ZlPaxl3WtPuEiMrt7DOduxCcJyZdQdKa9M5PTCkeA9pVZdZnYmAW
MrX2wZkZWo57Lt5GnwATA8tqFq0wC2Q60cZOdizBhozq2jMzvkqKkwc+82RnV4WM
skyddNgDE4OcmHG4PIkgMtoFDlh7+M9VVqMPhwBqhLE5sdrO2INfuIKVHrbVqnK1
y5rjBn1lvHbNFI0ID+2zzP7PfUAgzhFrB8/r6GIdWZfTXDPhYsyT4bXtmUdzJGnh
CrNi9qEsTn36Gw5/BY1Y5s86t1cA04bErW+IL1ju2q567Q6QrXA3RRsPadaI8nH2
wgbJCjkWcY9XI6rl3kashQyrMthjUlIb6PpKZ5iAESa/OkqiTbRxJbO70WqRNDVQ
jJBRWygkKK7UaSEQmbq0wz9Sh9f1f3HJeaNXf6+jYJPQS5pHgKf5VXGZuqaHybVS
ajinK4pKAQBf1O1UqooVofFfIKvDd2XqywP098MPEfMPbdkjNDwKaFu/U6YbJcZp
V/nMn50Lphn0KvL3Iz08uCitdGB4Q3lZPKfvq/wTLi6cfQZpy/8MtOilcWOb8TPD
sBz11KR16qNzj7AzdGSKGxWtD97n25HKFfAXRCmGmw7LMT7dxlm3hj1IgrW2kObP
/ei/Tt9xCACLA+wLQSFQFwJOLOX454EV3ZAM2xSZF4q41DVslA7+qu98VOATAT08
eKi7YhD/jNr7esMrogyUV7VI3ba0pYS0CzHtMhQiepXxTIn2907XxzKtJqlMrfD1
O4cm9POjXGqqOG3dqTroxclSgWxe+/ImIY7ROguRqvUZj05z2ANmkUnwc077GXB2
O/bw5uaJxkCr7D/HETIw8Y7dEyQlgR6aoyH8JlASuHsq1XV80xguZFmxm5/cTNuj
ALMep2yhGVMcclCqP6sdYAwxN4QNaVy/diNuAVGmZ096tinpVtWjqIkksDs3+eIZ
lAZcbu1GaTITMInNkwI5Q55yWpb1KwtX+Im9wOd6KMLrwzV++u8ouNEx8HbiqNSw
uqcnG3lcV+dLJq5S/NW+efEAnjr1txt+1+ur6INfycz9jtF5QkijdeI8XKOSa0JW
uF9EQKjAiiB89wXlih0OMkmp55pI30WmFsEQ9C+z2pGIiepI6zQwNrkhl52blwEW
HPCILKSNPBn/5oAx5T4cZic+qFD9rVVXk1Vci7xuCrlNqbkuK+aogB5gJ5nyKpQ9
6BE1kQOE90MG6dnjiGetFP5it79O3Qv3nJoh3jWqpmhTi4FXfpLIHN8TGC6BpxBJ
1XmKUe6eoVVhJ6x+O6ltlWxybFDH5AiKOSpw6LFeeoU0duKUHSqaXnBPirOVqBsl
+deT/sjxFoeVrniGITn2WwEGPykonaLrIUgvgJexDEijNWCcUsKqiZ1g8sEObAe+
LVs/w1aJziPu2nq7zRrcU8lny/Vy6qcG7Dfd4idElapzzeUE51hK72bUJNU/DeW9
Bym8M93anFSn6qZnF/hpeX2Za3FvhirIneq6AggMkV2DAK2CGZT+ys4TAYDkuO1a
5RRACxC8HBUl8GhDysA8VOyI6yuBdmfaIalew6h+++5ZsnfeqUUE76o5EVd7WheP
H/J8wopBVJ6dOMAIhUeOhr7OHcuTKfwRNJKE3o5Br0WZ+OO+uxbV3HNUyK59qg8O
uKLK8w9u5eTkuVA1iLfYsBM/+U2PheSDztnt/GFpHmm6Pcgs9inkUEuQJpl4kZFE
WUERZHgexZep56jIeKKPvMIruCWwkBclZBRg0EWKQwAuFIBD0RW4xG57dx37+FDO
Wl0LKRYBxiUhdbu2ug+2UfrRe2FAemIGgL0qak8IlOT5SXxuoW3Gu5KTGBLYPBk/
f+gY3Nf6PCKMj3feZFYhIqbC5Jh9/f6u4KTlfQMWNZAYAyydnHuIpZG7j5zGbPRG
6Mkn7Cp8du9POvzHpAntKdtOM25Md8tjn2HkAFN8xONCOIeFiO4ZAfNzwrEuH/B4
SAcZ3KHLsGGPUnJD6JIjbH3+XawF8gTyyPdiZwMsbCYeSqRomLMURUX26wy7RtAx
mCxYIDEepMwgQE8F1jn2Wscqbu6aRt+HM6RwI4G+xGA1cG1OPoq9uo2k9NfW9GTk
871NuhxGGXPj2OmlmIbSNXFEnca7nX1AZlXvz/Vi4tVmx/PYKYQofb6WjX6jR8dU
wPW6qMAVtsbLWymunDrdE5h5Qnydlb9fqa2j64r4tWE8udpYNT1ffhIqa7UYclW1
ctm7pLqZjkXJ+pNE2WQm7/5mgY9a6jmqn3Hn8OdaTkWENBXRUrS6Y2u5pyeGHDgK
KmpM1rNmlOzo1FympFiI2HTZ13d7xC3yrOjIM8V2aM0tbBHgiSyHmq6NL6VECGLS
f0JE7WWzU+oGxOPf54W0gr2UWi3X1N+x4o/LIhkvMkAwJPhdblmwxusj6MDStb8X
oYKY2Mv57jTAqdHcAftYB2xR68Y2gYNaHNLbd3y1QqpC7tUL7Q4wxOu8Jhf1CzNo
CLMcbU6rNPnVPv5VzRhV2nzs+QMC9so+9lwURAHjsBDmljOcEvHg/13azag0jwir
suueSWjmYsLDSrH8D+XrdcdCepb3ag0nKU9DBaGBWa35uCCvgZ58KH9ns43VWDzI
nq4mXeHCVZ5hvmdsMETC8pScm/a1hZguVI+jQVNEi5L4BYyO7Is2ht8JDSKlvzcf
a2+FUVqAqhZ4HQZsPPZxvpW5BChfhwxRrai+197L4Unw0QN5T4beB8B/oul1TDMb
7hz2cCs3EGC6G7R8PKDQzdx1RQDZ4qp/vdOWb/xKINYoG5fKdXTVe+UlpmnYUQNg
YJ4eTX/gKh3nL9UIjH6Psthlcd0QGCXPh+kz7HydTNBAwdmXbCGF2uW6jPLLeFbV
MkcZUih2UwYIN4GdSl+7bLzRULwGGQfy5c76r4/NOZqhgmiFpmtr9jTXX5ylXs9Z
lDnZ7Z2AE4ay1IWVD05KlcSm08KnKlnoKoRz2Kc23qyIGlktZGuaxbyxFYvv++Q3
k+z2Ws/pBZHss1wN5Wj8iA8iguHq46VN8YIA37dc3Oyzz5PBZv0OyIaWl3bGcdMW
FhPvsgc6w4dYetVGu2Rr5L7dioDw08gFcS5bFsteUvPEMwDt8wao3SM1m1CoUorn
cWvsWl0eNI5EXnfQwC5WJeNN+maQWm7aYsabRyMBAE5t3vAyKwedSXykZIgcveMM
V7ZvCk2mFOptCDqzaqmOn66RRs+hyD6RCSLHPk7zvNzci+/s92spu5Nrx7n2RICM
F6fLb1HHejYFbYzyTCe5f3a/Osgf3LMX30XYqcWL/Gm5QN7liyb2Amextq0xd9Wf
9F9/SGxt6uMh9kvdj3F2TwcaZB/1JVS/nVsx19Pyr7kCLtVdHm6VkLmZGlN0cF29
GGO3szjUPLwcA5yA1GBNbS5N5p2KaHn+o45IzGMbfm8s8eLThzVHN0Qa9FjKzZKB
tbo5kHTdp4Pg2ploLlLTUIrry7/+GGUjRYol1wj7qYiM7pXDtEl/4v2GtSpTIubc
fOXCHs4WOexevll29EEp1Q/vYVjUabaXO4yDGJ99Up6K8gUcTSxqCzg86L2olv0/
j4zwzmtubMr0nb7SPmqwReGXHxhqC68teqoJECwvRoCIM9GNfgY9OoKx81tJFmRW
fPXGFoINV0kGXRNp/EdURkeIcBMkhscxGqc/CAtGeaSxWs4QO8cHL5vul2vdIFXn
8CJyo9w4Zr6ZW820cFi06bSjkG7xY3wFjiitWfmCTX7WyhxcdwBjHNL5mN2sLdWd
FAL4pd/pfqx3qXXUZtfwRIgVNsfr3ujgQyNYT9AuNoMdLnNqrKQgD0jq7m3GO3sl
z2RxirnW7V8bleZzA6ufMAJIU7uQ67ucHgNf8uf30h+2YmFiMpoNVof3iAt+oOun
VcwuGdg6mzZpLWdHN415ROFKMFtzQ6TLW6W/I/o83ql1yrCKha+soE3IQZF45s6w
cV06tZTCgSWd7pY0kxHDfvLpjSr0xu+NHpPJDOXluiLySNq0GWyVo/7Z0BZeqJqI
igZkXvAK+x/DHO4RzQvoRhwDpTm4lnFx0mbogCzx6lox4iLNx0Ev2Qg2KmnVYlP6
ArEiMVwceYUbgK6J360SopclsBDh7alPgxC5tRqcXTmwgrl49D81iha31J0DmQ7L
/3aRznT6jsJiHTmOODb8isaS5X4QeuTTPhHMAQCoqMvmIPqcFVJaGkZSrFXBJgR5
WAsRUDSl50uHZGiBuMlLut1z8DJjrzgrBF/TzLVEJcDWIhlusdlZTZ0jLuvSZIVR
XsbMPfAFAuutkCUkw3NDDCmhyIXGcpBwini/4PnQGmLuXLiSW3ydsS9ZkWPh8tog
oocjnPcngcIVwxFvcaeDj/ZBjsY831fyItOBc05+v9NTvSxNyDKCVm17dZKqqgrc
Jnz3RNuWhtfGMF/hXiZu9Sm0JNpuv13XoVjJelsflMxr/FCyffrwLTJveZcMTxUU
JD+ElbfTiFUj7IgsKyQKSE0Mt9rxJFYgy60acUF4FRw9128uHal3ala34I7Y/W6e
p1nv3v6h+F7JnkYTaeJ2RwAidQmdYFBp3SNHoZCg8eL4xOiusIic7hUpdauvpQPx
pTz12f1rqn0jnmb8v9/lKp6TkI8tNrFjuaX2mg/WkAA=
`protect END_PROTECTED
