`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gzJg5mS/xGl12wYRv+AvM8K+TwUi6k4y+aRHEUtWagkF7uObzYlnM666jAkZ76VY
KmcoLUPpc/Z7bYjX0qdz5QyK5OiJZ9yWjSRRX3Fug62sFXshmZWtr6diuw9Xv0uR
HV+x7hHwxpAlUnpJIsp3vQhgULo0rDdOenjWWOQlox5iH6RDlSnmiZkLoIHCJIYY
ZHchmPo4xUb8YLwO8Z8jZXgojTWnanhuSanmpgUgsbiCSmMo4+mxh7MuJRBbwbW5
HJU5RrpkGEYDaJJ3TuGuXMt9XVHlUX3Z8iUeDAefMT3bzE/Rp3Bu9FkbVAr/Pu9w
ss7B1LvR5YIPFhW+CcvxSjEwOS76p9daMx7HxGbc9nmH9AIvQn+JU8QNtudsTlYT
OtJpG2MbpoT8MRiL/LKMe5eA5UbHIIXp2dlCyh8pTvamDWzpWeVCDujC/KHp6eNy
YmGoIj/UlTXfR7nwKEubU5Skx4i1yMxPqew2AY8JRfTMb+5oumw/EYzPoBnw6xdc
KAdLJhqBD8Q+W5yHDiGDV7FMjWEDARXmvyvgWyfYG32NOL/SDVxMsKu1hzozzWPD
4e7+sGyjyVv2WAKX15QcCoffdqImAnZ6ew1lq1E13kardE+rqba3pR1yEpA3ur3D
W0cCLejIaNbmF7/qzmZS/WDuE2KSWg/h5ybLCws4YSDlnclzXnYCKGjaWwx/ymyS
4aenzmZfz7IY16ZQPeUfkuXWADI9Dc87u2n4xkCqSU9lfKWcFMo2OHJiEF8sTsZ0
I8cjnrgIBI0O0UjUspwtqOYCoGnFKsqO7ThQItY1nUUARNI8LV9ESektBCYx7gSH
+y+MpYma0nAMmQOyg4QHYoLVwU9S1KKqLoPSKxXuvbun5IQdQOVrMMdbFFiyQkGN
6gW63C1gmwm5VyMUa9dq4YpRaGSPSzg3Ha3aLsOAgaOgkiJnpHMbfTv7tOsNR7wO
lNhaXkCAjWOyug0gF6qhdudg7GUSjPfY8zqBqLtxmNTnso7ijmaLaRDw4+0M3ug5
/MV83dMhgOyQwGI8VHtXHLuqswtZ+8SLlOcnCtDFbzFHtEjRPiS4jOSt1ccsDB24
zbLitLYaiXcmZQ35jQqrEwHWu+dUYi1Ta9xVU1ZWVc1Zuy4oGiWGhl9kjcnqpfTT
LCA99QbUPppg6g0aUPYSfniCbZ4F8mb1G6HOg084plGEdkabL55zfnYvHX4160gV
Rw1u/ksVRrhkMLQPU+U6OGxsD4PABwyfhklWOKIkQCQrGiDQOwBM6sTCLQ8ZmtWb
YlE7u82xCnLloIm6KHH+bSVCEJg2TSHfklIFBMVb/+lhQUg2kVVlt/Kz5UB6msrZ
1gsIKoDm1yeA9BiJrOkuGEyuGwkcNRw/mAQQ/A+I3Zzzw51uESWuoeMnfwxOAM9P
F9j3m1LbcS9t1OAGVPBzR6rDfnuuZauGt5SEQ8muFFPrVKuIAERy2h2xQ6i/jRVB
694W80rtOPNk+VTJopHGQDl5lw6Tnr1qRlTp8CR38MABJBsPb9i37SEXEXEpj1qm
ZzMlRneygvEJt/lCQxuoGr1NVvHo2rKjZCd8j5vUJJnlVAPxAVQmkvWEmlEkHtRB
Pfp7jzLn58/aKuG70WZX/I0p6FXbLYbOEnnXHQEclKY6PkEJmO2AHkKdCFYAJmxR
5KnMgEfPel+j/KZX2FdLRYNHkJhHeCoFnigO/oM66hHjaCPlm71JThXvPt/R5Ta0
bLSwgwYx6p1UPmvea9RYsCtO18MiI5zvENc6B6tOpr1ooGBr/PLves1x/jHDe/3O
3jA796/4lWtob01H2hrhKCCSCAKm+YVVp2gMzsj+AUtq6OEl+TE5IgD38h8CyYKS
Ra2I6FglanNWrV+d+cI44NDOwNm6AXsKl/QSWOtCAmDtSylSplnLC9yreroexy2w
+Gxy/gRGuLnstaVY1jnsCme5DRZItxlcxULEm2B9Jca09sJYy10rCnToFySnjuAL
UaBE4GFbZ+WbGuFVZa3db/7B+YKoR59tZV3gYlU9erAiAcwaKdx2G/Xz7aM3yNGz
5aQzgMPQf5r5Dbyy7yOWlQ==
`protect END_PROTECTED
