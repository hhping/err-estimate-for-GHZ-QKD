`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylKwOayryhiAwG9ZA/Pn1Bs4WHAirjT1sOQY9KLFaRoZdB1hRnhK4NoaRZ43lYZY
rmwlVXQGhrc6ytzbT4cKkMueXgl89W92HAdbgPGDPMg0AM9TgcmEbFgV2EOBRQkb
VPAATzfolVj5lBDglhlSuWLpP2lX3CLq86zemiGwtJ6NmPa9+NPQb10hr8zG6WTo
iVojnJBbzIzy8idkdPQWu98c5roFqdHYTeFPQFjVhk34dbEYBKXxL+xehKKAGtAo
bNDJT+iAKDxc2nx1A2p8s9yUmTlMa2fFD8Frgz6MiTKjzE6Fs9G7SWhfzxXwxg3n
gnKu53aHT4cuaLDwuScMUTf2AXWGtDYQ9LSLwxFBmMMJKJO5AK2LftSdO0XKg/kj
Q5OfzzVoKURqfEMFwf6tTLkhdDI16L6tvpTJwO9DlL+c1pJQOkTvoOymKS+pEOEK
KRRrAWFs3arjRjNNuIXWsbQSzSua6eKk1D3gyGGOCB6nS9mmvQ3eqCE/V4Yyr+o/
LeeYbcn3XnwtCz1k8d2gZs1M99uC7uOlrEDrAZyAatFvTmvVHhDrE82UuCU41OuB
jZ1vVZO6NZ2T3u72Ay0G/ClQLjBX1+tZjnMUp2/x51xlapDtcpVYb4qZgUqx1sDo
GvLYHKqRTlx+GN75EjSvCfNTteCRMha4octRr+ucOFaTj89/6iVr+Ad+J2ZtuBGr
TRdWw4ZeYILATmcZdYD2tapnxjtmYhNZdOjAlVvkpgiq8nib85OIjjr2bZ4YWHna
vfVIkJakCI4wfm0VjnJbZqgm+bAopMXX45gWynxrva8ZjNAPx6qApnlfksnBRPal
aP0ZNF2g0h7AUEG/C4NSjHrOnfECVSr+Bs1UUjO1nOsOB41SaGjAp9T07DylLgIS
G749WHI/TXAFPPecS9L7QApY03FIzJhrTrZfvRIL6qpn1amMUMC2JTSEfvzkH6QM
uNd55zDHhRzFKaV2ZaZVm3grJBLZBGx8TlEh4zvokJ/351PlqxZoG9BZM56FwN0a
3dUKOvlZMR7COQwM/lnC0evCQnzzM1Cpr9bYFBHyNsTdZg4S7YSltL7j1YyH6DQM
NzH/8J8olO9xXqtLt39W53JvLe6iA8ZPXpcPQhRGHSBWsnqqbkwO6lYPaTEdawQn
tG8RUPRusBtkHJQwbIe+fglsVp4XFDJiQaANSofgHuBFeQQFIzS8ukVWY7YKRQhu
YDtBjT3oHrUrz2P7jJWlqsBhSri72P27hj755CCOhbamT8/SUeYyC9RKUTlrFqHR
ykvJTGDPWAw8QgsrF4KhpHQqm4ki/AzD6m5vHgtU417PQaTw4Lb9w+KU4j0c4SUa
SUyLD2QG5VxsizL0KpBR+H0gS1JtzAhwztyb2cmINutD0jriMy9UCi+5FJpomxdC
Yb7SAuczgBHNoEJ9H+z4Ng8w+NBAAH13fAEWEN7Y/PtmRLe5AiblfeXcCxrSvBhF
Oxz1uOeEasA6W5SVY59AV6lA1/I8JgZtrHQnj83HOq65/zTmloWlPYrB8L6gTTQt
KUJVz2lDDoBWwJ85WWOFTzUpskrvefNTS9cc30prD1sT8yLNt7KgnmO1+Ijcvjia
pAz1gANE0xf/Zckosqemt9+YyN5G6tTurH2VuMuNus6JsW4CG+aNzXIWoq8M9k8I
LHV/XQXsbXtMFM65TbS3bJhgbvI3JGmny6Nba3fa7+CRsxgbrrTkeMfxcf5DCK3p
fTmJIXXvOQrwwi8Lwa4hIlO4DPIo4daCMUVpOIYYWhUY4WcdP9w8g2sUDWlYYlMn
Z97SOxFOtFPG3D3iAIUcyqJVouQuwnDn11rFhiQn5NMQb8xNI0URmoQwwjh+t8Ak
Nh4thPqDVVl5xsyxuzvb/nIZZm0o0ZIljeHZ9hYKHTbUxBvry/YA4831hqxzb+Fw
w0+bXIeSqyBXv5xeuGSHRmdbIO186jC5N0ZalVTqaZPYa3kRFAZNQv9jaQbVqEvy
fYozkf3YZOfldwo+Yap1cGfGMV7/Fy1UH6eosYO+xHye2RaA8xxttoVRUI7y8T6X
YzUFifkEvzjPInpcNfuXjjmYGwaQYBGWJpHbzYmh29gK05+myc5LlE9XSeHCwxvB
5ED1CstTwL8g7iKUbBezgG2CFaJFshzDSyobfy1paDIvkQMlL4FIlCEbkExUP+iB
gGzzzw7qwgo1ejIkcfBdfCvG6lQL+LA8NGVGFYKiow6D72P0B7vlrjRVH5H5MgL9
5eNSIxO5ZfyEiVIKfFopWLQwcW/UEC70djCh4ZZlCZLHORIBsREKbV0O8tG/S8qt
Es/BcNwmA+yYpKK7sQGh0mEnJhpLIJlqyVC9VCVgupyUdCmeTpQskzoOWAlxn0B5
u+JroFxQG233lERHg/vqvT9rhUZuHcCTLdpVFA55TS27+0kdFq2JRjMfac8mCMXD
3yLp/+Z7GW5JN1MMxa1T5AwllVHTYG/hLcuY8EcCZSRFYuUA+jiiP96ioEJf1b8a
Fx897zPUaRZDeGCeyaGQpGhZ5z7a3m5hvXT0WzFxapied0m/+BpC2lTA/23bObPq
cmJ4fvtIclfGgg7SoDK5y+Gj/RIb0jX4zcQMGO8IG/5A5S8lfPAbon53TX5z5GVy
mgyJQdwpObs7keclMj5dME9cvAmqPNoohdbrcnIu6bXoXs+rY4rPAI3Rt9UKca01
+YlMbJf3kG1RLfWk8NPS5V21ZajphjiVHstK56+AxIROQKFmjbDoWyx5zuJWWr6r
hN71HNNvdPTvBSxWlkXNxbpm7eIuoK68bohp9lgx74GKlnXr1QoFM88lsLJpy2EF
oMv1elX7Ziyye4+ZRITb8O2TAViiZuiR6NZ/N3BsKPsXAqg5hso9Gw/cYQG0JCCV
SYP83xy5RcKSWtLlfxkb47t4B9WuvSEcYMcjQlwZvha68VbRmoVkkkmu5Qvk9yKe
4T73D2BeF/cMHeYtNwTclilSUtZr+SGJGIV7G+hr0eo=
`protect END_PROTECTED
