`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymqDsLFY/eCh1rNqKXMCBWTOxEILb/P/7Tx+hP9CJIGtbBjPVX12Had3WqociCcT
N6X3ZOomPzFJPzi++Rzdkihy00Achk/Om6cJsq+D4AwsGskY+3LyU1BHiNwDB/cK
LE6YBDONakdrWeTwtzEW6SX6p2XeHe1yWpCDZ4xXcR+pHInGuTX3xRPekfPFRHG9
SekKWyloLiiwUyZyMuOFWIPMReKdTp2uE1OBosF7s9pL6tqPfp89Nh2bZbgpv3uT
9Llxb/e+uPNqm+oQiflqOTd01ojRHmbrbfgKn97Or6sYDgZx0DqnAozFuP9e9bMO
GUxOnIr0hbY8YKFfDIPy7eWGpnl5DHXGqsBihnOATj9slSpIQXmrclyF4TzO+2cJ
OqbFstgVaml8YZsbGfq0+G/xaqUyzoaG55+zvF2ZHi5QgkbqACNnTitlGRplik2L
NbiXUx0nWfP4+UmWVcwUBoIWLsImD9jxkScKqVkL4bSUSbr03pmtBnaif1SSV7rk
QYjgvOGLeHhnrAgy3xrwaiPY3vgxc0umx9jlLzSyjqC2vZc0PffWEvZE4ZpJA8QA
Q+PXbpp4NpI77tV89g1YkNRfpkhpATJpIYQ82b7ICWvLbRYics2l3kF65xVEwE2E
JrqrOjeF85AFs0fjLmrQFZ+TdbW+yWRqv0vbxRS1cY755xrUlYLS3sXBpOffHxLh
/85IE8eHNiqzSMjJAuxva8Z23JM16IlEwNDn0eBmIkRDu5kPepfmGdND64D8aS7o
54XD9pK19SDZvdKgbF2++O72Sd9a5wwrUyP8E++e+LAwglBeigcP01RsPmruxDyn
BZVp8w5vX7W6rrggBZtmqZM01R2QgEiGK6qip6hSkgsF25D2bq1L+rMjCgGfl1mM
EqvjqeUNzJPZ9EsYuMT0+7HcIdha0bD3YZLqMX0uB7C3rDh/7LJYP8TIbv0/crjE
B+TLQSOcYrKATWABHpcRj4JOQ9yxqUSXL5iWaymuLyuddTkyuZS/dj8AsbSfgnV/
gb1ZEvnbXvcr9U6tpuClUVWmmwP21lX9KAqydR2JzUB35ggSNDhGoGCfjk66k3hO
nbY8a2157X/H62F+Dh8tfP5IiRhsyg4lXCTfK09/WSKuNrcX/r/F7kAsmMVMYaS1
mxFfxV7q2HuHR36mBnIMkCX41xwRdx5N6XPaE89TW4/RrmOEqmt+swRBI20Zo5GJ
NhNbi3CTBuKIF5gar431fEuLv+qLDqESOz3OOa6KPnJzQ2wYr1Y5HPPBb1izfEcs
W9iLXRNK0hJa6N0LGbcplubKX0EzDt0BHNE4uXAu3/pnh/xqPq6gLVdf9U2vdYjj
oAwe2qFbnH955Ii9Z3Gn6otIomhzzSANlv9Bxc8sp0c+oeKbR5v4CSkGxL23O2KO
7X7GqdDTwoO+KjrYlDTiAFU/uWJtz7wZuy7RZgzYw6gRBsxTZu+ogSXWWPYeXJ2A
EHVAb2e0j9IRo5+vUJGFx4BTjExlYsp9ol6zaZAdS/6sgtU3rkNWxhZ6ehI6UaRe
dh8z3KwqkMaIO2rAiXeGdn+MDe1N+uMLUPs9WIfgHg3Rr/NMbQYPRHaR+9lRSnpd
Wxlw6S9VVFlYye4FZfstHitRpGA53ZDgnyPEkLLUZPOXvpTl5bomnTILxKB2GnJQ
ZxT84PJbfJAGuyOLJQbKKOjkrEIDWhZSCag8KLzsi8B5Y1xhi9TFfjmKBVxcGfRq
ZoqyMypSTgkPnKAHxrAi+mXlCD0qnZeDK/2CQvKOEafXU6TWOse5h6FSOG96onth
IXaKjACdRQhvnL4btEkS+iDk5HQ1YpHv3VEO7OYH9/au2cKNDchNbafP4Fd4teqy
07LUZS7rxC6GuXnw9es4+AjCncEKxE6HxMlo6zCun7GXcSgFP8rEumS8zRlyl3w7
4QpvTXJW7cZIKWJ10RxrHGXuHUYDexh6jY7Q4HCDCoVZORQHCkTaNFljZ+D0YoOx
pe+SVV+w51hhyRBroyOYHf9rjJ331rkR1wxJSaq6j6/nOhUOPSl/A6IGJwpwM79T
O8GW1YwW8gGsRGJQlcttePxyMyeb4fWooUnSO3vFd/WYCGpgy115lOs5nsVa+Gfw
hWhR0CLY+VVDhvQA0weUIWOFJGje85gfDqasjkKQfUDu5ZGV4JbPInrYHqmhzWLD
bUGmMk4OA7LhLrqiYbs+7yskuCBYzxOiDIzYfSKguAXhdFp9ONTqts/fiGC29tOl
lbzc8cXcfSLPEileMK+ngBZLhxPSmDYuQvqcf3lq0i4xut3pg+aanX4FMkB3y0Zq
PSSmH4yhecHYZN+nI+pNdiMz53tEoQrA5bT4ctV0vC0=
`protect END_PROTECTED
