`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxdZm9BIxTVAPG/AiJpTzyG/6Aw+uEcTxYDdqjIzMExrY4UVL79NF6kiGFROWGEX
79YVwJVKcAJ7kjvQ0IHAME4e9fUgalhnM7Et6NOA5mYNUzfaD9/xXypHlhQyHrQD
vFeF4hWWv61oh+qvXtWgVVgTynpkVqfnbTxFFTxYwYBQpXixG/F/IhkWTFx2mzMC
o7jVTUGjj3wtGO+MbIOOuSg3P2beojJrohjdBUgDlv/WLdjp2qA1uB8xkCFaW69t
ge6DbuVOcaAu/yCutq0MWwzM1sPhQZZdZPbIgbU0+R6TK3InFVMTBIRDICV5PliQ
W6N5w4bNW6sGh+9gh3no4v7EUlBX+7Qt1+mCdEmLmnoZAu3rh7RBblDEXBjexc35
QPvPpPde7LlkiZ1lAXFx7KGkdRWH8l+RnxAgWwlHxHtu8FBWcoxnmBzlgVbfsW4U
nOftejVRwwtLPjyVR5J8Lg==
`protect END_PROTECTED
