`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KmxhkNjiDUD8CpQGulrsNkG9pMFuGoFnOrDGhBlX1KNcQVHlbo8EPg3qK/eW9dWD
Bs0jIgOuMjjl3TU2f1wkiXlB9H5MJri/dNmuAkhRqVKMdIi+/+r3PEYGx2O7GM4m
aFapI+/1CvdphnDLkXPn7+GmHqbI7rAl0BHFfNC88b6t8cJ/urKiob1Uyv74ihxp
Y06AVvEN4Q+RwifkwnJ0nnRzbsjR8WICYbEYhf48mx7cVtgswM3hNH1llOJz7p4+
rxGzDXXZFx/YbO8YUJgPd5SMYmuFLzqGu+RgcciDKw9nFPEYGpR8xm/QPxuk91hF
NSO64SCGUcwOpijrmOGdI1JyONe4zXw61T639YxT5718neyWgo7CFy3JGVKCazU7
scHDZzeuzU9fuAwjGvB1uaD4BoBB5IeLFqu7VFwoJA2c8dFbwDUwt+W6xh4+TC0H
yqLCh2JlHMwCpY8bQubED1vOiOMUv5ur8xZrZokIKqLiXvh6ikJdPeaXBGpJoPJS
j2EFD8Gq2v99YHqqIXEF3zVZbp04OaUKqs6lvbeAC+sjEguiQiYsRpE/kzL9nuAp
TIKFNxi043OTvgMOZXd4O7MXhSIXctGAt+1gAug0kEVomCbVDGIfmaIL6TjXoXre
GOje25Dn/DS3rDfvchi5sRQuW1TA73fItqy8yUTr5nxMTIblBwaofmhg5cltL6nH
sKGgg6vGt2M2LdDndJBsJqY8thDOghdcxq4dJHtcKWGHefbTNvQdoPKHQudgJDDy
FSDOwJJaIpgHNJ2n/wTCfkVb/2wgIu/Aaon9OrlWMOaTh9jqPwDrd4sajCPOTKNU
c4rB4naAADl1sQV2qTshIbPi35Z7Jb/GUwgWsiRCBc8j5GSbIb2wV18oCp4HYVzB
`protect END_PROTECTED
