`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UMGYMnFusaLkmf5L2ETrFvk4C6Oi5JjKqDuNTjk7qGiDhOnTci4JHjdqGOSm+K5V
rbNLy/MeAFIsnM5MKvqSOKao05WuZCvjiZc9EJ69xmjXugT8T0RhZhPLZdtzfO20
H6MFSH9gmnMiMe8CYUnEj1sxC2UfuSFoEM+1rrI1xs7a1FpancShYLKs4aR+MJN9
FzWEG7Pu4bVq/NkpjNHYhGvKKVLhVStGuHNzP7KJft3sTK2Po6RnatL9tSXz4iIL
cLHTUsD465pxyE5Y5x+FevlJt99GYMz9iUSBnFSiznGl6iCfIMx10hz9b6z0qjih
Ydt2uxC1UX5l2WfDOZAKSq1zepkKSs+YhnRMTvpeLxhXXvZkjxC6SvZZxsYDEbDO
gcRhmX4ENKGdmG+aQbB+xVhq918wwfRW46gkMk/1AcAz1NEZWD/dAb8bz8Z4+qub
nwPcRjWHR/JwvrOBn5JWBoUt25hOKA1ObazowiSEQ9hRv9rB1H0sTjHdAsGA5JU8
KTftEO+q6Ipk2T/F4BsQh56T5QfcSSQq+yz1EtxXxHA3iM+qZ9bDk9gdG0QN7MBR
d9lMLpopTnuRsg2hFHQ3fUk7Sf1I9w58VKzbzYfz1rwgI0ig1tsmzQHDjOOjxw9b
cc5HfrgltqfZjoOWRrbZo1PgUrE3Sjs21LPO5rYAqB5ifnCoRLqt0fh0OK9CyyFf
Er/IfpMs0CqfLMjjppkC4Dp9y8rBkYhwrSsBruKjzsj97TvW2pGncTAbm2nkhiUx
OxElzTTh/UZSs1fQjftS137BWLzYrJqbhEP0Jy86KxdyabM9O/E7TRuMFR3hj0dP
/3i5DK4mfpw75gU/51TAf4WdoBBJMQoomhmvn0uf/Q2Rd4kjJ9FWCyxO8M1AgGeP
YqL4F5Bpr1maIi9PIEVeXueBadGrG1ESaYulhPinjbnsIP0HF/IfdHCQ9GzDU27X
E+lkwzwNIgn9lm3TQLqMqDlwZv/srPiyCCb5hk7+sh4xoQ7VLu4oIl0H2A7vdwRE
EEMMiGb59+8Gbru+tk1m3T7UPclwFM26DfPLXRZA+V0L61VOCPz8dniQG5tTk9zc
ofBBJH1bmnrdp32FZo4ASCAmc+MMWgF35/MfJj6U65VI/BhzbIC0oIzqhz650KrQ
Dhp3HCarnXzKxCRiUXb9vaBQ0waLsf/5tebLnODgp/lFIMuXHL94h9iGqQRe0iss
K+Dgq/N9z3ce3yKqPA7whNSPJkBqjIhiq9p0vkhGSeph5nw4Un1gL2756JdMTj0X
FfcKmgxOACI7bKJmDKwTDxN1MLiuv9+zKN9RxWvPoyiIrCKZ+kFwgAXXbJDEYHfp
gCQymP9UVvuzRp98hbCkI65TvbWkZCjohdaubK6JrinQOxeJij+sLuy4ogngMiEp
D7hIFKjOrEy48nV2YTHnWRfyjzhqNpnaHrrK5k7dwMJTKUUs+tLrnDpolTUHTKh1
yX/Hh5KcqzNoAY20l6+3vA==
`protect END_PROTECTED
