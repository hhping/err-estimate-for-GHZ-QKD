`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58MSZuBrYrJ3JkHEKGknx0RGmE9H+mt8hY8uLsjTjhRPQxUibxh6BuI27sAkjWZN
pi0/2qHYw/2JmpEabfTNMUTuI2DAw/SraijUa5C0rqy8C3/WlCorQ5BDBcB1hWsm
5CLF7Va+ttTQwoC+IgjmXkU5v26LUkG5gJMLotjOC5aNgv47DZHHnI3Fq5AMcMVI
VTHlDpQ+MQINPy6XU0yKZKGZXqNUze8A453+24NGO388y9Rl3q2oIjHj35+uNE1f
dq+qBlXk4qrwUT6yqnPEuuh7RfGyCdjkjxHIuOr4vJS6csvMLZvMIDVy0IbYAKUu
4094OSay2w2KXvAmbMcgTyxqg1t8enAoGXPSagYgmS/2SkzMtbl4LJNi0rArCLqC
r50GSRz1aAYRjsQcU2AGCfLjr6RFpgpUqqVQNFRwBCKtahYQ18db1KcRSjCjETe+
OxLkAg6Dfsi46GDq/AW8ACK66yqXjqjT+wslUPUzh+MpUWKSplUz5PuGUSAYwjIF
SbU4qoTCNNWT9PcWwXNap3btDxQ1SNVPiIFpB8M5nGDH939EPGUgknFDjM3YkxnP
7SdvcGu39yDWJp0ccEUftyFPe4RS9BC4/K+XMnwcSrnsz8UGlzDqrGhBOMJUo61x
DU87UxJCCL59IWysBZvdCc5YxOygBa9tsH9cfI/EwtD6IErX4JX4zxFuf67v5c+x
HDD1Xeu07brF7JF2uL7/qu24UW5FYcpPY6QUwVRi+iGNbSCXUPdNPq6Jjtas22n6
9GRhbWiRA6owr18ULvdj54LKscPUL+4uTaFIlz9xuqhxUc5xBtQ2oCZ+f7S6EWO/
A4eUVW9cbmS+bmJ8zI+IweD2kU6wykVJRYAXc35hGqlTnnZMqmg3qfSmXRGYduUO
C7dSWjKXwJc+7S+mGOaJyNPb7haF5hFczGhfWX7S3oNZogQ5wPeGDaI95pUx10K1
3TU5QmzIWAMpZQtjipPcCAjEGdIieo101c6HSv/z2W843kLbrBAmjpHQ5dQoCv3J
FT+em1HAE/mRVazf/QhCVK0slk3k90zf6mEBa7HR6kTXTWfojFFMx/NnyMIB7Kot
MDpgdJXUWfKO60xTSAtdok0OYtworlmC3y7HmpGSgikdXnFHFu78wsrlSM63hKZQ
1XTn7H///x5nXuaP7PzWaGfVB2VYEP4jJ2XcCvKnAk+lq/CzRCcNZ6sPYpskwsPd
6GnfDErH5Ptb/3qeU5nX9uWGmptiuD/2tFbHjgmg0lEKYnwzg+xET3G4dZvHZH8i
osQpxZPkjKfFTOKJrdh/dIQy9ECWsbWYoy8bh/3+ZcYgovEEKMskMUh44hNuY9cc
Fvil1X2cTMQ6nn/c+xxcv38SFFli4cpCsg5lKpfojQGsalAA3XrFECwlzm2nbdvx
/plvL99qOpQSisI3fGVW6Fo/GEFJZXHo8e3xjwk7WbbY0dDKXGjXhfg3d5274FEX
IxNru/e5tEwGuFpDLzrS6lkEFpaG2mTuXmQLL0FwTLP7MMhsFqF3hTJ6XFANCpsH
XAVc8WJnp7Fs0lvFvC5VgyqlojUhDCR4aVlGT3LPPzDee/pPbgjOQjEH5kl9rJ/K
CQVCPVq4dvnVD7n5w224XEY9KOKeKdpKx+sF9FMUFNqzRMNipVrCLLPVVCNMCNIn
qZi4Ruj4DX4MTAkhuy3aijR4VEMBCI4MiZllWtlIZTsVZgTB/ajcwOmbpPbgp1SQ
lPu1uqMtXL8P2YuoO7GEEj/9OdiDLG468uZNJsuHu1IepcfQQW5BwnxpvRuqS2tO
gfDAJw3hEeorHgeo30Y+0MgkA01w5dsAOyhs8xSpdh5/fdqzq1c4ZZgVxBBHdtds
CTrWQhmlkfMhOKZUBI4UVAOB06yQTGQGw4B8sz/kglk31m4NgPC9an3pYYnaDvVA
FhpnpXSYJ/+rWCp/euHipG2Ncxq2o7F1EVPWU5ZVrgV3aIrPZRcjTwHdhnJWpdwQ
7bafI6J24T9B3cfcpHKfNkziUf5BkNUw8Uklx8oS6mljDzvInuA6Fp3/E6qsGo8c
nsaCyoqBbLh//Y2jFcBvmGGooqyO5pXSEpUV1U9mqWVCX/VCZoAF55vYHl0MTl9H
UTzBlT0W/tKManW5+TGFCL+zbp/I7v6t8MROxm1V6mUtoIVRJz32hNbZGK6pvT7W
LXQBr+xc9VhbBNFHkXxM+OVqVxQsP90CKk6mCp/v2AIe0FEaf+xEWvLNFkhzqpFp
i9Vr6YjoLFqkHhU5JdiSBElbq33B9hAuJ+dRHBB2e6Z5gd7EIhKt3uIBEQ8PybhL
fmPWtrrNuHqUOjDR7PM2lFfkWsp+mCEp7FWZpWBPqRLC3OhPQ/TbQtnCLvplV6r0
HdUPKCpaPjBvDZmsVzPVVEP3dWrkFu0OJdHv4vXeE53uMpgIVn4U4Ypd1AZCah+9
+PwNAL3my7i8FmLDihTKienpxioXSVb9OFYttjyGX8gcuG7XC+rslsm2uhVaTAgi
ozVE2Pwawc20+IyjKOqVrDTgtIQNsZno6TQdzy1O98cFSoCCS9vMHdAhZVfh1R0r
ogOQ02TiJXkSFsYivLQYoanL5ZUcf1+MamIpMMahL4X0DclrZ32G1ys+lr7vpzVr
uGraNVOyT+WrAsppBBu/ws4jUGt6xZ68y/i9P+3ZyJARuN4WCsH2tGacdNyS2v2G
j3gt0OBdymUxdCkEtdI6EvDUcdsqbbKhgUAr7k6qa2h1DiuYr/pA5E9r7dYMbRtM
bHVjvN8TVnUV4vl3AONI8Yf+z/0TQS7u+zUfydmwBONj+2+G/lae65k1ikLsHnJo
OTjeBXprRkoxi7bpP/B8unaDNEACQMhE14TvIHwpo/TZe6yx6saXhOQpcUfqtXwE
Wot/s0dgLViWrPlmHGKpAnBYv0oufvR+RJS9/KtvDI6lh24JxiebhjrBg0Unbha3
rZSgLeXCTbgohnS4gARgRGOjTS0dDblVIAbm7YIbj1+nNJlQ3oqpM0misKu//wFf
gLrihlCf7xTmkLo7715S9/hfw12gv4mtss7QRjIZxMkqi9fFj0yR1V20KFdeVq4b
MgVIBXGzqlJ9mc+enJl804pDkuOLoKxO7y7Q1lvRE9ZHYV9f1E6feN9HF/FE6YDa
y9wXqOcM269TKoXmusVvqD9LTdCa3hyISrZ3uGhOVobroqBh5XmQKLjmd7lVAPLl
NCIMouN3j/igNoDD9eAvilMYWu25dNpCb4dC9A6YF2EVVZaE+CE27VdxkbmSNUCq
pmkK6cjI6qmMrL+e/isqL2U2lAetg4ebGZg04PzG7ecs5sY2eDjgxrdHRBI76zXB
us85X+1REGvVzzkegak66KrGONRP7MEHnLC/HBT0XXWypAxeh6W9fwoFcKI1PYWw
gnSznY4kVayE7a4QiAaEB3Xl1TjqYmmvNkEc87xVhldCtAAJr/JDPIx1kRPUYvx5
0XuxLXBjGFd7tsDUI7VgVu1PWGc2xvdnc+rhrFTj+H0cMz2OobFL35UAH2KLKntP
VmtGoSaw7cz+RmCPcAZRX/qTpU1FNK00t4mEp3JU/9olvHWvWUStGke8bPcXqaRo
Y2sOhU/z0jRN43B+yOI6uMEn1SOF0I5WLbNPph6ZHoHAOyYSn4PLULK2+ZaP+Feg
pqNL3W1gf/IBVyQp4SztC6Ck+BUEw9PiLuxIkITXqpprkVL0sJkBNLMxQnMTektH
0Ozj5GkadrpbEFwfuKMvagQbkgYxzZYYx1dosup+f2gGSJT2tJVhRWCddvngoy3Y
GJWa5u6iIKQzlaLcfn9niVaBtvy1U4PPpGXV0tK71XJZN+LFyE2AvwOJLCcqD3zl
f2kKJ+QLcE3owIpfRnpF4ffiXNo7RmQdBepRYOi1sP/evTcO6xaGL7q3Se1ZvosO
1RQvPxW8t1t/UOB4bBqyF/8LLt/cCOiaRihV1+6qgEtT8Pc/ZId7KpZrNjSkIyDf
D/u37dvS5BMkS5eU9VX+3MpBFcREpHkN8m09hwKX0wdS2twgj4lEvow8QCtYTk2S
/6mw4af9AVfzQqKDAf2ZWiRXVQIkbgn2OqCeXSpk0W3QblkWnIval0kGxFRPj7qT
2jv+4N4ThGN9DodcfTEQlby15rhTQCu9d7bQYPb+Ixnh1aV5UNQDSCYCp2CRzXXe
xYFfWL64X7oY49GzMpC/vZyyvoKGzWefC9G6LakrMZsC918wcuJB0Jqqmlcg2qq0
ITxCjslBs+e6F3fjphU9+Ra+AcDQ8Sf7lbhIcPgy4V8PTg5Vg+zJl7naS8j5OPIu
kPR7pJVdpgNm3MSl6nJLnbakW+3dDL75JcWTXF+ClxMGRUHoKHxtNzftkCdQtoMK
KmBEBjXu5l/C9qdVPSC0eUxBTBqEIakxuOmBW43sWbTU0gtSLgFcRAFQA1TTrt8G
hP65JibFzzsIVRE4hT5nrISXRAp2S1qX8+qjmvtLE0/RsvAMmMLkoRnKFusXVoSQ
b6a7OLp1/Qh6BhetMWAon2Kr/WOj3S50SR48sCgg9u8jWak+BDP0uqO9Z0CrEyVu
6g7Bb8BS98c8ffG4Z1af/S+lL8fVrR8GW1tzofUEDAu849/qpfSQU6yMrDdwH9Rg
VE7HfltqMMqC+QiGwiCAr8CY1HJryTl88xmmyC0o/lcLo31DFfaTl3Kld/gbeZ6W
F7AkOgUHpxULxQZ8qSjufoFdspk4P/WGaW/x36pN8fR8q+3Hb7akLeKzphk32m+p
sHakws6FIGtPFVy43I0KVCT/y2bkZpzdoZmN6YPt+mUlANkrj96klfUYn5BvTzBy
xPfOr6epNkkutdVqprUoB7LfVSCDrL1ppKPjYbDKYPPRFWTr/JYZIRcQCuWF6A00
vnx8CzNZ7njpBvPjdY6C+ED2b4AeMQuKRX4LTRrihZDjnFQ4i983HitUQcCFdAso
eP4M5yF55d9svLY8QettVUxaB1Qse3CrnqDIr8nqUIOzFvZadtyznnYqkzlKcg7W
F1LUaTVQdeyZROa7M7L3jZXX1lPOdBrCQ0i3KCgQOebEriGSA6CErwG6fB0OvfE1
RLx6coCJbg68+UuZtGeKH8Hegvp4nD7FoqUn1QJhsssvZfsGFc4GHOn4hasAxSsU
JuLB3wlymF4jEfNGatC/pu06U8N+c9Z1fD3o1DnOUkBCSrX7hp0vqqsNHlmpCGNk
VelsKApzdN6x8WIsi12YQz4U/xmvnmlh69Ms9RvXNhC9EcLfsgQV8Vc30a9un5eh
eZNPkhEZ2NeQziaRvGD0MBa8mtyKRyA1Xe0ZjyGcbG03O7U0IIwp9nenEvFQFu6j
9dV8zZ0kexlysHvBTj+f/ge23G/WpinaP5nA1dX6WgUZttOXE5q916EAAYFM1coF
lJyXevy1yNEjzCRGBaVEGPWjzX+NHEqbDdEL7gnPiCtCzIf0NBrPCnLtpRiu6I6N
TxSkqee/s5pMarplFB1JOkRrfwmiR3JiX0++NtnujVBfYhSztDOWbr2/PQkKxVvO
1LgGZlR+BwO2fr1Pdcr18bkMLlAYJqh8hznsMXKX7+xNLrDJ43VTYp7su1oTau1C
DNijT8JFPCHOYS7Hu1Tt2Cp+ZMRD4QBEl+L/tg3knf2LmCjcXyMzGGev/uVH4Mgi
hduRYsntusY6i1eRJ5gOm3YqUxCNvGYC04YPXkqKwJhnru7OU1THOC0KOmCIX5lF
X/m0ojVO18MZD/alVmub9vmAOWzaB23kxIFT8llzmY/uCN+vExxZw9CNbZPu4BRc
zdUEblm3+MZM12UXOpDl/jVXEqUZzLC9SWhWU8VobA686vmfQ2026ddZ9vIwvMvT
x6hY8KiIjjKPNATOhdBrN2Z7Wg4+6n3id2sOjmFdgR0AFLCol6vIO7D4xDjbeUzo
uvzc0Lbgfv6D8IlJmk5GLHgGLUOcWcXdrj8xfBXikJl+NemnAuqjVqsecYSTYUP0
jxEVTFXI1gxrzbHfXy1pTOobJ+MUmCW0Xm4/msrrdJmRMAVOfvp8pkbcRd4Nh0fV
bpRaF9V0ymxPgCXtHviAe3OWrZh5UjFdTPFhT4sJko1iiIjUlrqxV+KHXieEDPeI
5rs78MCiX96MSQGr8OLhj9Oe4F+tZ+sj34yVgYtQaqDAhqrTD6vwGxrbFAmVVyMc
1ACY2C8ca08HcjwAein7Ojp7OHRVQF6sRCJ2kbQ1fon0fngxnmMANw+tX8B/p1sg
EhUISrGRW7wgg70hfOeUMcloJEPr8D5Ti+VJPIlXEXbtnF4ORAohYWstTddeIa4x
2Aw9UGJ3pz+U1mZnMzcn/uWO7nwWqlDKCVAU0wJB0zisMf8SOaQBIFp5DIYVxwnk
P1Y1d9h6o7KOsjf/UGyrv9y2keFW0DCtQ6RDHhve8aL0Snt9pqBpfsHZw3Myv9OM
v4DEHU2EIRkhuc+djmA/yIvQ3Pih3NPN8pScSgtgwTDpE26vGEKnzrGJkN0sI/AU
gSDrh090JRKcwblDghnMnIMnMJ3+BpIuIg4WgUQK0WPvhBWrLOtY0R5n4e9Zemix
Bwfbvyq4gnWiPo5y8XISH7f9P6DcKFsfTe9SFP0LrjJA0gu00RpC9OrGotkBrSML
JWw6BarGulICpVlB+T7KrvVXdwl869aWZ+8rz7jgzAfu/NaO33WyHnAEDXB0qmvD
jQTD0CfHDltGC+cFJVHluhzQ7qJVdbpFlxQrXKQfTbLF0MPJ3jI3mq0JeQ3eMQBK
p/ZOkjWYaSdlKVb+nqNhJj5BJ7TvFI7uIyADE/JIGNlNTcr+mOVjxDTtsz0uavx7
C0XgqkiJLAZj1OVY7RSu4N/A/JUt7nYB/cIA9FZ+MoU+sQk/v5nj9bjdZ0tZUQKW
evqvcjQeX8i53zpNjRDI5zWinfCSTi55cRDnMciiGwDInVVeyV58RtOoqmTdYj17
nCBY7hTWMFL6jljzwtSza8dOMm3XSfslAHYAEc39bWoaJs6lHyi98gpHv82hshA3
/pSMIUIIou+BPz128+SsOeVPFD5W2R3Ve220Olm7HZCUdRkFWNLMfD6rtmurKvkn
CJVZxZjsEFwuJ4tIms2/ZW81UTyqeZd1ab0QJHX9XC4SP5vtpPZU25IVorLLXTb+
VEK8on4K8gJLOyl+UsCI1DFfdww6ydZFpcPmFHcVyzrZS+tHKUWgUO6FYnXkKm3N
6IxOCIK1au+vBnmtoFf8VKkpfzTlfvOEVrH0lb28T0a2Jw6bRKVQrso2BVrIedzH
nFchNxc3pECrkcTzaf7Gme+DC5QNXKPsCBWMxcdCQ3TvhTmHyncqjo+j+bYhDecU
4LVTGLAjerPapelh86MJ7y+6/FkKg+X3UoLjl7vAEXQH8ujOoCydxBVQ6N+uEkVe
e19UT0yK35o7P0G5wje1ccCJxQrpVEaY2t35kUkPnOO/sTV6vSui9uexXwg/29t4
xJVXWsQm8FI50H6PIajM6IPcxG6ed3q8Hfnj6a/7TKC7d5u4MSS6z71NBK0A2z20
Zph3myoMT7mMv/+ZXqVglJJkc7nN/t4Dzz7SC+qGZubhZKJaggSo4h5jtzPC/GVP
6ymTrO3LzdFOFi+8cAOPYONRc+/j5CWfR38hLZlIuX7i6ASc81BCnAsjz7LwG09U
pUjLRSWQ5YeUJzdJIzPa+fwgOX/TfXTo1dkbtXvHEUo3ESars9FUf1/garDCwBOn
z9rV75hPR8pllYoIPoQsY0W3KfQslW2nIXdN9bRRsFe5fGAoXKhExqBJsy6JtGR7
+7nulHbM7zWiPJCvztoYCRlU0qXOWocmHy/dX3WJqCAHDvUA3m3s5Q25aKcD4ZhL
rE/X+oNFNhlYI0yUmiVbgoKLgR+9fShjVFftE4FZ7T+LEnvTdk8Z1N3pk34jjor+
UhiMS26+WKdkqq/rP7vb1xSUK8KJedF6151a/e5XsZQv45OxSokbD6oIpXAsmOq8
JwRlaWcQhez+mgld5IhkzUMEwLIdLC3ckAuf74u3u0EWxcGd4IdfKvv2aGWMjz1u
U36ozBmakK+fe9KJJEK/Os3s5z0Pri/UzG/sjdtBzkrBjfDbWf4PBFLUvZBXx1jW
QyKGymS54+HJNg2fPDBMStxMKpbBz1bpFx7Q4S/NrDMA5PDBitBSUzTbl0i9+G69
lQ0RSXjsAT4Pn+ZG82aOPGtlbnQyONqhDtAuSid8w3JHf8QPkVtcGhEJM0CKed5w
wBfLXAN1E7JuZiwqAPqbAfIUQzXTGa3X10mOWc+LO5bXYNQYA+Y1MSDXZKc8Toc9
VrpQiXXlOp+jlnV0kzDfRX4ArJYVfStPB4qMl+rOHTrZ+zQZ+LtoEzQRtDpY2Zgs
C9ciA+X/zGxLLxWjA1CoCxSuM0hhsp+N41K9uLvuY8rVyi0kgdowb0fg9Wtczjcj
6/x7wC04JTFIo7N7if4KAj9hpiEKie3hjo1aNFkDU+CMl3ZpwXGKnT8v38pVx40b
bgKIHoIrif2DxKIHLjOKJV7+vSr7AX5bOD88w5WTaZC66k0RKaHooTAaIloJZfR7
pYv1z7Ofunpz9XOYntr0VDCYe4xHMWnPSv/ACEzN4Z4skhjjAwj2qbAfeKOoFya7
QQlf1NXaEGGJt6fdEO/NspYlT1WerHkDEui80m/2LYxyY2EzIkT5ov1sTrqoBwup
zTa9QmjTgheof3Zco5ZvPlkpS/G0lWPEH63lasbbUkvWAJgqy9bkKTKaqcmTDRI8
cleqaQlZQaUwTltFPQdUYzPyyprBasosvs85fUegM9G7E7+kO9uGGdNYxa0DsO/u
18qc32o4DGFxPuhNtMENZ3fT6IeG9ox8NSEXhYMLPFfr7gNt/Ze5JrqSOK/sVC1Y
B28rt2kEvPFxlWd0ymumwbft9B9bMFfeCLlipzdITM7Z1M0DyDeYpZ4E3+a263FE
vsvX/DUFio+Wqf24pbBniEZzKdvjSXaL15fQ3nuwJikye3uSWHPuAWAQqhJIKeGa
5R3oKrKAQ3AznJRwLsyDFiiRX+25TN63T0zQyPbRa26IXrMNGrsm9pJHOYytyWqB
yvYKhKDUnJy+zOUfrcbNihIBKXSPvBIghE9YUs/zvwJ7ztTiYmGLhp2/j24b/Wu3
7EUCqdmOa6cUEWQPhrIuSk3e0fZcfAAVzzXN+7Bn/RRiY3px2X8LZYNVbIY4eeTE
nvVyp3cUwB4lpkuoK6B8bOxA4Y1FeRvFJVj2b8QCMNP7cvZshHhKu1sH1PtUIFLS
cpAV2A2/pan64lwADjIBbWjOL+PErDiA8/pJ1t3KgCeIV63t1IsPupqrs3PI11nE
TJ6tCYE9r5Xxvpm83317dUL62sxF36dSO6Yl4BDS1e21syLw3qQUlgj1MAx6kPO9
sO8QgPOykbUQi0WR/ji4w6nNLCoeqW25hbJ9AKrujoYWeiuc1Qcv//bLqgLlxelS
kNkZAnq2KuD5EuFVcswjAF2xHaE/uizYyIDaKX6cn65ylOaWHXOFivNpENMts5Av
bjA6HEOwEfcar1wNSknyjFg3wX6uJOwQ7jODHwAx1zQEin6/jbC90JmG5btUQP8g
jmD7a6ORO90BuHu3pjM/LdgSbFC5OkW7rx8k8PgnE7sCTEKOkCFvGiwnFriaohuy
5qVFvQ//6VqvnKONjfLq1lPcVSxPO6IZ7gLTN+W3/F1dBaxZ9mEPbtHFsRKw5UjD
SMTGmkc+t04t0KfyAnvfrn3TkZWNVj87xbDYCh3ZC5/iBBdqac3Kyo8zvxdTjWh5
JwbiiuM4UJr97nY76g7Kq8IEx3q9qgbfzgXiqrgfRKxtGxn1wfBArxcdpHMsvbz+
7jOVxuHlr+URBtT7je2KiCA9Wk7hDyZJ3XNm9Qst46/Ug5oVs37Saa+3cfkjRYLG
qvE5uf9Yb4OYQ/05GgZ5gdHAbh31/pyG44EKVpket9RQD+/+HGqSLNLu/3WhVIUn
q92EZg+F1tPVapjEMUN+l+P0311T3VvTQ/C9T2cK3s1cWO3C4OvZqgK/CBCxU/r4
v3nsO68nHPbszwWMQquN551ZXV5zVPKbq8TAq8HfFtIa75H7JGihy4baJWo/L4cs
YqYJX60X3BMVFkrBFJfiqXVJsZMg3eSXXEOFAg/sNi0/UL7+eATaLZJIFLxy85ji
rngWoqpPg2sP57iyOVWmm9FvH62ydV9eOwYxWGnZHFO/K261HkhLvRFjD8GWPENO
NHadyeVgs0L0gesBkm70I+mjnV8IaPM33ZvWJFC4py/IJ3QOzgre7gwVXfi1oLGS
7P8rODG5wPxMWnEzdOh3rnakrYr800wfsiRLrgsPTQvZScGyIYhaXbF/ZJiNrqlg
xMftRhh4NTelCoO29Oz9YNL8GEmLwV0PP3nHCbmdEtPxHpeVHASfvxWCv7B3LKkZ
wRjtyAcOdCkVl+ka8kAEcMO84P+/bTA7GaSSpyQMrzEDQ3WXsRsurwLVkEUWxsLp
9xYGnNgY8stYlOjsfHd2+NgsyqEqHmwRrMG0RZ9oM5+wMVg09UOsrl99CvTVbZGF
yvxJVMrVISdvSkNkgLbpkmn6c4w3X6VtLJovwxukoA7KISyBUd3O8Q/BYZ0QPrHg
mYaCgzPujkb6LJ7KBr7XceoRkc6/IR7iJoOw16f58oxHV9S/mbUaLbBJSE8Pzf0S
w9lObrurlIPgbkS3BaNGpTYxtA/2exc+loGS/Mj02BxzVUA+8lgV/k2aE1kAfsz0
LfiuaA4fK7LcWA9YGJsXJJRhNVgUEeBAlfQj7m5iWlD0bkN29JM0Obsc6OcsH/80
gYGZqUESeDAoKmCtNgsMtCymwjidI2dd5m5T/P0IpWOAEOjg6Bpe9UffVl+VryXy
nOYqcRR+Lb5gkrBxVbHd0RON+iDYX2gHn8lR1CG/T2ybClujzd0fznDzKptaHB1Z
PaUp45OYpJvyIb02u+d6Sm4kb3xhdxLryc+58KavaAvZPSnP6iQxm1QPmcfU6faR
sBG8/3Fcpjoqc7l/afrMf1uIBhbDCziTCoc6Snq0WpzqIher3ECnDNiBdSMKSUeP
RTboEUhRCM6n7hYzSAyWWXaQtoJjlBf9PkHfaQXOfWKvRk7lle7V/Dbg8wnoGwvp
UETMzJ7dqOtmdTiR6qcbuHwfLn1AQYAGs0RMGe9BQm9uzgrUZU8AklEMvQUkDlMM
hVDNZrWV3HNyC3wjGiePs48bJQCj8tWIBMlD6TAKYpl3MCiq2z3/daO9LMQgf98e
DYbo+aPhA8ILGOKrFMs7kQTaVzTPeilEouVeUnwYyAdfAvjMvJIWHmawPVcLTFkQ
ADiPBHkxOd7J5PE2adKzTS5DduAaaYm5RZ/itTIehXuccWDbhgp4l+H6Y2YONWBx
PwAxlKForCuFZ1uSUeOLbC2gMW1r1VieJxQdkjwdMpmm24uW8JiVNKT/hPyOmHD4
gnvTwuGSi6yBYS8zLAarEtNsqvHDlSUZ7nZC6KjdlOTiLyIfvZw2F9hSsujEi5vP
nmBojbgPeko5gPKwnFAVyUYzB8cTVrYDaSxQPPPjax8YjQYwGHBzvVaReL9I06eb
AEllCoHOM+zS6pPllJriDa534JRSvSWq23qkbLp+tLe9dIMX5Ih97mcJIlnQqsuF
2WrhEA+Indxy9D/27C+KNktYWHNMY6PFQdD0BQrbcfGDduAoEH2pJOsA6MtIPQMU
cSlKLpR4b6nwu0/w3AFoXooe1uQk2W9tLxZem7yO1aGiooolKSq3SFD+N+ffI9Dr
4JR2KfyM+WeL2atDyBU68nic7exI5EtAwgKr4e9j5s3kAaj8WXhMGP5zXmWYYcev
WXpoWINduax0/2xeuYzKlCV6dCO/KlR3Q+QJ7UTCveG7P/n5yBXP2Sp66pk4jxlL
6cQAOMDoIyTz+o8biUiHH/VUixBA+ECdolBTXD1ssNaQxUZwcFERco/ydqWhztri
FxnkgY8+xH/96p9gqMHWkm6vysBF5qfuluYzW0+hhqgYq7qe2IN9/z3P8kmIEdgn
jt8GT9OkiwePCuB9gkN1UC/XXf9zuZAabuI2MbL5EbeMxcZEz4PSvsfWG4sNF/P7
+RRoMpio9MVwom2FyuKsWiHaeqXkw7iiy8HWQxWliiCC0I2n3oPoRUFWQzOLHkD5
VhlOurWwb4LftMClJvtfyd0/QB3Gb2JUvNoz8p+0NLWMjhHXUucxC4TcSYW/HK4c
46YNf1pMlIM+nqZViJohgfDFxgvX+JyWkRFgJbaymnRo2ikXV1i11gYMs6lXN0Z0
46I+j2wjHWStThmm9vtDO6EqcfEUTb0PCCqb0hNlcyspdodqylitow1HiPzMz2iD
uEQo1JsVpOxMx9aeo+5iAS7+FY+FpLBJIvShKsThO2Mc1LwMMmyALNcapzVkR1zx
OBK3zBECL6s5JciC4tXr+1mi93weld6WQQfQ8Z1XkcQ18tcjaexn3HJ8ILs4UGVX
hWqLc1LyLCtJFuUojHUqAddx6yCakj6PLA7rkoMywbf56U8XX/UFxXeVYTIPTiIY
0PHcdxXYha++lf7ilC12c9dObf/eHTeDsb2DeokPr0Nz3Ee/AUq068OgSIIw1vYu
D8an+POQvWa7zk4J2iVAo6FFpWNm8hXWP3bFEMsL4hRW2MZFJkl5SIGFK56d6GU4
F9Nzl+MPT+lbb+YXZRpH9s/lQ0vDAMgjNo5e/InvOqXP+DK67TnMYZ2oztmx9KH4
20TNzMEJ35MZsPRXbRXikHP1pRvH8hxJFzMlHYE75HDCikv6GopeF9bussfgzQUl
UlC8ikiSEIe4aY+O5OTtfbfgjP/Ebluc673NN+Z+hH0TleBvNZaInCiBqs+FtcJX
WtR4WVo6MdC8oLUwQM3nkY58ETiwJgphpgFB7v3Ah6XstkX4up69pK+WjAIxdjrt
LO0bIpW6TkV3/mH/14+zMwdSHENMgyw/QtPTZvyKnk2PJmDMkSSGY72JfCN28OO5
bTvxYRN/y8BKvlfspFBaXoEQ+fCakZ/B7RWPMl+7Y8t8/NfB1dIHiN3+W1430aWf
Sm6hZ+Wc21zZVx8QXU7jmNTQvUCLkNQCQq1KThRNV4iv5xNaQ99L5FRJ8w9hVWCb
Zbi565XxEXvTrE43GWgShK0wA86g0xEMykZpo83tVvY7U3viQfi19o8eD+CRH8cS
U4UXRkZmSOKgDvd3pgmU9/JRvEy/Uf0Cr4/qfP4rO7QPzhit1+Ow6d0PAHJW1kXl
Suu71Jb8GwJKPmXuvr3JumZNI2xjpRZtH9rEDK3bPUP5lATILq0E/hTyVWUsI0S9
+hNTcfpZvOomZq+OTDNd0iceROFJISCAKO3AF+3fRjsqVF8SStcWyptOdQ81EPSj
0HU1IBxOa+uWtKO371tRCmaQe2zs6kU2tsduD/Q8+FdQ2RBXyZMUMtSQlXrwWeHc
8nwfOVyad29fZc0a9QXkiSwVgIib3S8NtS4ZBBCKx9fGVPUNc6EzdHRvD6JZMrTR
ycY26r6iqblRURkgT/BJl6JY4i84OsyJ8Lr5DoLuYFq1M7PLeCgQ3J+jxV14soI7
qUrmoLbiSY6j/I7+kXsEkhiXoEon8UTwaQuvIOUR9bwWzddBxcxoUvDWj4KDV7vq
/JPdEYW3CSOJSH71lki0qdpjUWfYw0NRyoajjO8T4s7hOIh1+Da81EP5fW7TZvGH
On5Ua04DyuClED/YJJ/4cgt/fUe81lV0oSwmwC/ywp6Tn6KKwbwVuzs4CjXMGt+Z
AiDyrpwe0OlOc5cbcXdshGx/np+khp9eVY6xuI0YhuCx+EzhA/qpyIeX8l6S+f40
XmjPvIkYClWo12z6XcA6lv34+y0spBnP3uwyYpK/rHZ1ZAEtByjyydLi+DaIftgl
N/rd3GENnlXcomrTBmH4bvrdoj7Tdce3s8YUqb8VWK665vudVthnNwsgT/C7PEiB
XR0GO42iYoMPrNHs/xuJJMkaeV7Qp5b0q/wrQRtU8emMr5k5sCByXvXC0fnzT5xs
OVhgclW60MprdE3t1u069m1FENrLTFDg9e8BwF3Ji0m2kaYvyynGA4AN0RvDd6PY
KtnXZYttjcmCJgtyKgBbupwhYxi6QNNfqg6w/neotMN/D5l/j3yu2i5DtVGAhWkE
kH1aT1iRI9Aq3CYpHzza5WZI0E2JCgpEJ0q8Azxd4uE6tjIkxcxbHrWd60IwnCou
He9HEKU6pb5lGq7xWyuLWIOlVGwH9/5OlY/HnhiHfyb5A4MB4HZYBsEYsrWrVQ+H
8eTdm3qKNacyYwgaSw9zM8JT3VSEdxZElZqeP58Xf9Jv9T6VXpfyqJeK4v0EAMsv
ECEw1geMB6o9HBygeGO0totB6/jpiCK0cCTuiDji7gtF+XLBZySgqUVKN8q01NKw
g3Qk1Fw8M2CGYfZKsXd4lJROOP44hE7H3VTcy7Hnr8ajqXudF+w+n5+Uc/YyJIOZ
nySGs0neUhG4fZF34nOoswFanG6haGiq3qW704DBYWyZFx+5saGq59g1P3A6EHzt
aoEBpobf7Bd8w+muL/A1GpXc3iQT6Kw8IT79FGTjLJbFZxIKlIxTVhY2yFRGsRM1
QJtX9W7KHl83VaFwIvqMnA249us+WH2BIv1MCpZx3I6dlCyxx1W1v6jXa+xzvqoz
Woa1TGMn9y+QBKqtFFJ5r3o70afsqU/DAlHapdbGkdB2jyo1daUkyr8v+UhvQK8y
Pr8EijVkGMH+tsepdLnZzX85DFcB8mCmMaN2dA5PXjfTewlG8z7sxT4ub62JipdZ
KGr0jZlz7DBDJ+XBSd1WYeb1ZJRqDQPuRIz3yU9Ce7E5P0pJNHpx8dXNtzadelgg
fc+nwJPWY7X7xa4NlzF5TsEvCLW+FgoCSQzwunqv6bdAugT1NKQE8X0sM5fH/u3E
gHM7VXas3n9iPvNFSTtI6IohO3FUILDToa/J64o8oTYqdCB8VKrwLaJG6qeuKWjm
XBIZZJZnk6uPa9qr5h3HL7nRdSqF/GpNTju4XLll2zougIthOos0w7qiL9Xwc4Yg
aMgE7NX8xOOh+zCZHitcXFH6jLQutpKGJlsHwkWXa7PRs9SHubNmBKgdJ7GsnL1Z
8mGf62yiUCXuN7i8Qb1vDmRjGOpFrSTUv/ToJTQ/duuu78EYcPIXjJLo+0URzPvq
oQXEQlp3nSaR9LxCqjk4OfFLRQhLD1VdMIkqJsL2A1Zki4pG2ahwgzCxOz8d2Lbe
c6PVvI/SDaUlj4AYf2ke5NVGc8aaTnIlB9ihtFT3H5AbjXQtuS8SqtB9eOJhHZTp
eXrDmzP/CtwX6tBKqE5aS8F6YWf+D5UgN3vvUNFsiLeMYGUeEsMFnWnFNO/JBg3e
D2WoEl/PvKkF8F7xXlLvBX7UroPcmd9qeFGRf2WJGJBL8UNhozOwT1ePfbjs/2Fu
go/fU6U8WdfjHq0sDFw4CpXsZ/CkwQcrnlA5VPMSk+DPwNh/gX+6nwfSaff4lFXu
yxLn4dWwN9pUg3Bf90QPQ8BTEFaLtsp0n2/RXr6u9bo0dPMTgZ9YprAzLUYrgtJj
05z1smhN+z/Q7ExXolOsYTqiW5eQSx6277NrJjTCp6dAXp0MyKkA8+K15kDHHSg3
1xaiWOYfHIetYdqBdgU6erlVzTz6/LkO/Dy/VKWb8CQDwkPFjb1Rj5VBFYeWfzRp
kYp67kzvgxd1OrxorADKOw9poNy3E5J+DEF4PDK9nRfQeP7vcAiHSh83R90zZmCo
6vSP2/gzo9E/63FdXXiybNWFfuo3SMcjcdIBTJFKHq/Hn/019hxzUtfxNohaJ7sp
SzZ0tk0tsRd2mKSccGhdQjhynj57kER/s2tuKJP9pIty9D7Ym3dnXUyGXfRRidkq
GJceGE2z1jxBpBF9n8sY4XWnDbsYtRtJ0f3mmtRYGwuu3NcAmF4DL0TFRFEoJmzC
nFD2XMkAMRH6eY2LEAvFecL3hKtGELgNZjFgFYrfjPoxyMNNDjyW6w/h/QSexstd
BydQ8jbxprQvP6nZoN7RuLvw5Yhtj4eFiyp8eCsKoLJwQDltBT1/nMte0Fkq6PtH
04DVUKzmTd5fyYc4BYht8daFPeFyRaIB2TAFEse1viGwapbUWnnCCp5CQ18D2YW7
rg21Nyipu+1nXyt8IgSrpWC0ykWIk7kePwwlP+q1cwSXInA1Bif4WR2llfB7/4vv
5IEGtSSzCf3+XMibPex34fehXTV/iE29vuRfvtTGcNuRSwPQJa5puYMpD9ElzyEM
hDI1DamMSE2Q8ab+RtM0W5BAd/D5m2VEVm5hfvJFwOQN7bMo5nG7nKXhcT6VgTWJ
bdpqICoj5TuVzwWhfzfSIx/l0KIKGg6Aj1IbZKTFi3NZbrFfeVCpIqWVzIl3EnBA
tNzDl+s870ZvPUbkFzVK+K3eFnPqoNyW6qpCPRcWv4HXGQkVfM3sAaT6/23Sq4T6
TjP9zuO150bTHnW1WLg6uNzxYiTD/K+IgAJwYyasEc5V1xE8TAQDGETsHjLrHDS/
9fciEWDLYZCUxByjtbxNAmdyfesSbvVY3hnMeOdLvAPGCfxEQRP1gpEBLaA1Shrd
/4YayleCG+C53lfQmK5BgXfMNsmwnPLU2k4p7xniRkTvj4YlLMNCwVO/oTWEnTu3
4g2BSrm1Sk9LXFRFGl+gXm9UkTxOP9qju6FA04PkC6vepPkf4gh0+NAk1NufuD0z
UywbU5BKkt8m4HmoXPpFv3QJR+OpTkxQM417GkJuRQlCtUWwNct6je96Orpnoogi
pHXwy2Vz6U7zM7vyGRXfRwU7wu/nayHaprgw+TKi68a3uzOmJ3HCskBKHT8tvnfP
rMymz7/eSXG649Zmi6XwL4ThwEIDUdvvlUv+N27+NSw4weHX7oKnyrPNFiTsgQB+
CBKe46ey7wqNGSdE4O4SF//0RK923WjQyFZn5WAuaUQMftrwNlDX/iHjVz5IY90t
cjpcWlMIzawE9B7HjdoTp1U6feVKBmYUO5A/KtvxGb/XeywHSiFr2zW3xQatmM4a
8le4QoNLaER4zBAOIzxAjorCZ+33sL9NmVLVtHXHtMW8yhm2dYNbDYxg9JUyO2/p
oOydsZOP7Wmg4BUu695+WgcHGIE9Gz4QVidDG750cwRRUvWVxBVmo8jK2QSkgly2
5ynECKGkjwtOjYoOV1BJFbM7lgkW5cB2RPpWa1MYVZItf/0KO/5NbujzgNwe+af1
SE6Zx6dFS7FDp+73G+gw4vu0hkvR5suhpRSrDD0TU2uYGFQrH+Dl7l8ymALlqTZK
E85xe5XQ4ZDtuOFVYhtigFqU/rDbixp5HtHNgZACjkBFVvdFiMAivs4yW0tu+G/V
pa0KMPCKXlG39FbhJoUBi3tBltpqgHCyxMbNK9NRXiRpViCdt28YFzeRcXTI9bUz
vKVUQ6g1zdc4HfTd+Fliproem1rX531O8hsBCWIX9ZTh2eeuuWqMbcDn/I7cHYo3
4pgUrEsCgO2UQ1rr8jpaDPslZYo1DePzE+9nLC07Io7hQiOag3MRvKd3JiIwCciT
DT0NLV4WoetK3e8uiyTcGBMVOHDJOi5N9Yp+cnPDKqBRn84OmsNcHAeNhg7HOOx9
44ICCFcnXlvBS8ElQbNj12r/6HTOzkOXzn5oO09FvIQVJFd5SUdgUzPAnSMc/B2i
T+u0YjK9pHSTBGnmqLLRjYjQz376RzNe4g5sAtCfmqINUEfhCAnaGt+LZIKtvOkP
iswg2ofka9yTB6Pi3lvT7LY/W3y421wVm7WEXvl1wyMjMY3i2H7hWPqBGslxmJKk
Pm5llsxrhmisq3QGLwNsxWeVG6yDSXjuP58QSqSX3G2ONj2J++5GsbDpbN/GSAV9
wfbRYKf7HuQRlgN1igMHauu88koTkr2Sv0wH6n2kzEAjO/aCI1aTIgOPX01li/nz
XZ1vmmFWiY/Eilu49BRZYk5dxb0iWTYuKGfxcynvy1RD7SNJ/AOzByHLC3lCRrsp
lvs16WNKhr9ovfV5B1OCDOKSPfEAI4IYSt7YBrFGBSejd90WBfbG4O1VAyQ5bY5f
Kfev8XJuQt305pXCXxChaJETYY+jEYOe+yYPKYUc9jDcVViBI4uMJn7KwB+PwHKL
BUxKRh9a6W62iSrBYXtvSnNjXM+NK73LHeh2yiMAsDMsXdQlBJyNXK+AJLZV3MX1
t2K6RUDS0lhGTFwEP6olWsiR1cZNCzI9YgV4S+LdfNXMZaTGJwx6b/bzjyemZJLQ
zqBzZiBpyKkURpAoIEmmBGsw6wK2uXHvEONjv6L9OuzTpPWo/nFrfLn7y48QLCm3
Hm9oVHLZi2geVJ8iikSp4Yai3Pjg4AKqAHmBhWgHjoPXNN59KjoC4FPIK5xuFwIP
/bsReMX+KUHdNs0dfokPtwbFUc/Z6sFDBC1xOj491nXhKO8yYIYRD/tJwVErlXD3
22x5Da9xYg7fjetxzDqz0a/sMRhkd6tikXqChgbSnrILfyV9S/PYrVgiQ+tILpJH
CejksJmp6c/5X5niYdEOR0I+tVNdZ1Yo6cgtvtFZ4hqp2u7zTCb2Jrf7RXY4MvVm
A1xpmLQyiC/gyqdSUaI3dTVXLdfRjZZs4OKTE5+jpSKfVogeg6RJPrCXcI9m56Ut
UmMkqBsm1VrOESCSdRKP0CthWWhOGXisOeUPwK1A9Uyn+SXUFFokNF27Zyz66Oua
VNRIFr0e7WK/JHjjq80dunOTsnOqgoadZRKIPKkMctyM8LJfmWAifjk2nmFIVaUn
CkqmC2D8NeUlIRIN4RYGc16OsjKKZllxUlMpQ/LGyk+kisGTq31itVISqO4P6j7C
Y580NOPiurj1LOA73b2VtuxVnOgEFHMuoz+jLK5RFoZ1pk3j3t++xnF9s8JFcPKY
Jq6l3Ux5GNcdbNmTRmuFJnhlrwXcUnz20NbNTfnX0peAY440dl47UC+XqwlVEIKm
Fl5LjU+D80rL4wNDaX0Ss5g2lzy2WRl2uDuDxAgZW3TQ8EEvPXrsS94bv2iwYxaq
qITT/GyDYMY2rRZp4fTTSrdQ95hs0qh3FST25ErajEoxU55gcQU9UbX37NhXfun3
0YKIoLKKUlCSuqBzr2E7RfY1V0Z8czwXV6XnBUiEUgJUGvM7Ira1tyi8JCt6nuwd
o+KSdVrp5T6K7OVtlBXzUZx4JOE8LT48s9Zd/kT3V+b/BchgvsLl1Q51MX2tupxv
bENaHvtpOWcuIk8lCnSfeQsD1zmvAZfCR/heIEoLb+C4LVSOcL+BoL7NbNvNsxrS
AuQeOiUnV3PT7Gcb4WYeAdKwlSxXEUY19RgCk5hRdYP1G4f/LhuHLL0OxtzgFRmE
g4FDJPUvyPjXz3Ieyf9+RxJRQhFEEqeaHLaUTOVaFhLpW+zKpj2DtdA9WnfCmFwn
FDRRsba6c9oL62lHRIPMu6XwdTsa+FBKMD1BBODBSZydEdyMptIGfE2ff9FSytYw
o0j1Oyx85ZxRYw/NXREbPo2enwMLF75vdX9NulBtxSdopa0Ayuxj7cVML6RpQ8rr
Y2UI7m+9kkoGRewmhFxFNUnRlqHfzl0Eop7LyE4cFpW7pUfAJLGELcS3NBU4Hm/t
U4GOCqFa/1pVzraRuOLnQnVIw0HR6g9Xpnq+X/6CirQrl1QJmYV3MpkkJRLLzj87
Jxd4T3L7uOKfugGj6Oi/kfz21E+vo0l83JWD6IZG013bzx19cf30QO+gKKJlZZWl
pj/hma1H9KpX0YtrcX8TnHSCh0mJ+vNJZzm5g5MRi57b0VMT8kbsyZJppUZBh1FU
iY6/UMiPRge6pwdtPnYpa9+LEJSS1+ovqYD5zZDCxfrRW+g3b9T78xaFFOfUpm6N
Nd670H1Mxa0itznWi99fegEh12ODcHASN4+h3MV5IB91DE/GWd1qP63F6T2bkFPH
syjq8rNWvxosUl7Hmxq9KccIuzhBsFB3UOIx8+dedd5139/eK4aSMSZAXpVXRP3o
emlIKXAvb3bPaTJzE4LBATK+yYgwGnBENhbfpHkmahKP8OWR+tQHvfXLnDwtkr4R
YyQnHqYlYD3oiBycaTuECHzqzuvqUc/1tJE5XunWI1CFiDWcB3br46ttUXYpIJ9B
Hh2RD2YrnETiNP/agl2ckry3aCor/B3tPl53+WEYNcl65jejeL6ADkEqVdUjo8zR
dI+mpVxJ6Pdrn8CCxIFe6akInBVLXR/NKYy6qSqfykPNxE89wuP+rEH5nW9hfeBS
B3rMrbqEtSpNCqYiM41+cn3UYrfblbpx/vDpSHGKKrLmvjggUSvvYjHIETHF+NfZ
vI8Rbpron5xcvOSROttzt7Hq2tHG9CKqhBNB0O5AycrdPtCvph7QyMlGZwiPUdsk
Oneh0mrC/olOuZjqin7lXUFc8DmqarTg39E/VISeKx/h9HKhFpdBq1N7jvw2a0BD
D8SXbvCCXY/cKFrZJ50ThYC8v/PnE50dW/VS+58zmhwTA6ktUHb/f7bCsABRWyKo
/2UwEW211XMN0opa3U/0ybUUxQ1wRpE4vOFrt8MTVG3IK7YR2qs8HnQLIbL8z+Gl
IdmA7lXmeSI7+UT5gqWWxqCxhVdUD1qu5e6dgH3cJkeciwYAJDaLx1lkU0pcNlhp
2ay6YguDFk9vftFUOBlcGZ6ZXmBSTKYS64QlH9UqnrHcQ2zTAIkV4yrDoCbKjqQJ
NJBZLWlIyg4L2wwbCqSkw5fa6t0zdjEZUxgUON3mUwWqHPz8UVLCSyOFXo3cqnkb
QQzmfmsLOJ6CCig1L8ayQUsGPhkznjxN66XdbZM9sxQnCg/VDjHT22Mj5sQCDmVi
uN+o7Lvfy+oBwQZ5qVD2Dq5/nVsK3PfqEwcLDLcKQbQm2XCNA9nAtVsxG3JPJpdt
jDTsVZxrZv+D5JU/rNiPu/Y9nCPba7sBz47BLqOR7W9Vuln7QV14QPrh0QaV6kAH
PjZUQRsX5i6NZJYGuV2mZm1wq2JqZfo6cd8FFzpci6vy2+fAEHzJFG+5siAwws/n
KwsQ3nuy9WhGXcMwhq+9MNnK3Pp66C03XnchbKBYermlrU3FC4MyytFCn8G3MJWY
1OJqr1TrAHzvHq7fx9uV8p+w+5dTlP+s/3g/yA1rAnsXvmUqVYtFn4lesuKWWgQB
8qM5Hw7rJXgV2TcEadoDM8XvNktE1GD8/UoobmeJHUm2d2rxFrI0hP/HgKUSo2mx
KYNEN5f6p1/ziN39qhURn9BWn4giog5zuB1eNcilTLtEm6K0IUDF+uCg2bVjB76F
cGlHe0IcSiFXX///rIdo5Nc+lzGMV+sKIY7NMASZAWAjvMRvgDoesKhRq9/d6uLm
jILeelUnapG0I7lQ6TL8DhPCJpVB9JDZtBmcWzrMt6g5J90e3H63/n5/pUjNP7nW
GyTFs9Kig0bYLv1pqh+eo3LxRTnZAapNwfplyjESf4p3NIJnZPCE9ZQazK0Rda5D
Oa2JGGSwwX9fzHNap44xPkurnd+ZIfEXKsKUb4evXtUsxvZ9NjobFKviEe73nZVV
UyrXAyLkT9FTccDNgw4TkBYceap8ht65vN9Djm16rrki/aw4bXmwUvHtG2+2RNoz
AgTfCKGSYvQxyEF2Lse5yRD4px/DQp1uurJojZI/VX+GJtk5b3kZEPc0nrbo9k6q
G2omn4nwYFBfX7p3ugjNWifVrFxCFA3PSIugeNOiXSj7+IFs3xljC+Nji2qXSzFX
zR9IOODdQ6cS4e4abrpC1lZC27FrJNjlpzfHJuxD6OB+UlwZJXmNNCl71U5FXCzz
uhsm71CHuDzcXV9opjr7SMamFO0WLKFXZ36VfzKx1k62WHDXQpxaVZYrBHDmLlT4
1Yw7rB/lUkjR8rimDdoFpM4yVGAwML6ARRY5oXSSDBQhq9bJqTfEgqnDh8ZPSKxq
zXZ6mSItToRLA7WUvc6TfuPApmDTP81+b42DKOe7a9Y/imeMpAbqByN7Y+8wx3fz
WJKnyf7a8l9alSSL8lMtelR11dgAxigNZHQeqc5MTOCQ0tdP2aRq3UQ+MKyBGN41
XgE9Pixwuh558xS9BMTyPp6RW74GYZT4CorqSjRQ+Te2Xh32LZtRncjBjCxLzxsc
YzNj0usKXNODhRsQmZCqxj3tRnIPXMI8MUZx/aIzy7AAtIcYwYEObWlQYKRufemu
Gmc4t75FE6Vxk97lhr6/5KrKEmRuyx/r6sqyb1kxkDcyQ2yVOa7txZ3DrZvHILdM
rhNA7REuPy0SvHS+W2KPg4CKc746EDWwlG6d4eV02Q/Oe5FHqwAJSNZmlRrWAJjR
62vdxplzdl4cDxYpIFuNn2Ws+CzB3WruBrsWc9+TtWZ1afJ9ULUf4K2eTUMHHk5B
U1sstqAGUlyTmUnmDfjg1zhgkzp2rQF6NM+K90z4VsesmlVb2XP3//mgc0/uRhCo
h+ghOFr3bk2rH7Ky3StfP73eLRIyowGhO1C6KO4y0Kjeh6MTvQIWBUfzZkxIYImb
dQ9j5t6wYxflVzLQmDBdZtoALzoH/c8M0ty6g2iN7XzvFeDtfi9UnDWozSFaBTQf
QimuFtVUIW25vJ6oAC4BfisUYMNEgih0wgeZAtjvnokUEKD9oIeRekMzK57yzimz
9xs81rOCq/GbV3cNxtMhYvIG5i9VaJsyUorexNRJ2ol3xohlnOvPb34cfn7zDF9w
hscaT3/utYz7/OhG6aP7AKvRGRDobALK6baAN7YGwNH4nfjy5lc1lEecymx/Z4PT
b/TCHSGzNDFnu3Cexk6w10hBe5bvODrdG8mBKdQpK3tl2S8HkZBOUUaE3GSEL38M
73TQuE8ofZOV/MGL9gZjV8FieTXfaPpdAT1nvwfI1AJ/w690o55D5AnXLVPkW5kH
6AELtRYmz+WpEzY8o2TjryP0jmUDsCTrSIPUnhOLSKds7wt4lrkeiR+aEpyPOZlk
4q5JggpyBQI5lDW173Sd0ZHgYLRFw0oB5BxtY1YVrrHkaOPhSmYky0folPEwEsx8
H3MFs0SUciem69NjDi2ykLx14zNJ4fvqUUzVA82YP8tj/N3LFbT/0FTy8TW5EjcO
8jt8v8y2/vdrVEYri1QXVVpn7EkFUKbuH91L9ym+aDjn1Ae3jbaIPhDm/5MBXey4
Jw6ZqIReNgnZz45n1bQLqEUB1RzHSkIgfmsUOlEU/BAc6ik/mqvJ8NO9y8v8vyHG
S3YlHG72MGvH2gbVEKfbjiw9I840VPDsSfNmmbVXt2PFjfabW5fdMpv66oy+UbiI
4gdB/FP70Ojc71EHjTwpVSVHORWi6N4wVAY1PZ/5VrZQq/Mvg57tiTp19191tQ5f
YacxWSXwruny5pmsdmGjs4BT4nV9t3QLQWPlFt6tWfiSLqN5m44Ih+2FjMXxXicE
YeNxzprbRexmraCO8CX4J95tw8uW0XVTc9u2ffp5qRt/uE+7H0iVJVKZ26rf73fx
4HSm6VdHghEA8HIfBrx9uBZLnEAH1JNY2Pz+2LkD31A/FdHo3Lo7d6Ao7iGZ6ewH
KQ8nqYcIOpRZlV+HHePRg0Kf9SLP/SPpqi6l5GbCaAY0p2UrD6dhrjDdXVY0iJ8g
0Eymdj84/6MltT0PpfaeT8K+ggiurmpmJSe+uLq8q61eNjPSFepHUycFRwvXgzmV
sq2rgqVVrMqJSr5h/mqR1Rld3wX9pW1xvJzqbIm52vm3QbCo5nzyKm6rbF6VWs+Y
LIK2AdEGqoywFq5jd3LvCwBMrvzV7M6ke6cdnx3JD7pQ+u72kI1ciQrJbXlA6FWM
4AhBU4glHTfP1fUZxrARNMmCfqcnwSUwaBpCO7Bff256VHcwsna3GRsGJ4rAwJ/B
1GDVZVZqhmNp9nvvHRuOW1Ynb9xqGtT8n7+eciTs+yzz7KOrNT3F/7DMxVdBeWoi
T5oOTdVMgqrlltO7SVFaORuLKUKpEipIioPvLgaZe4LDaSpvefEgPDu3FYK02zY9
b9BwJTeEV6NQ/GriQEqD5hAkTwGhHULEYBOkA2FCG2VxBZZ0pq6AzCeeqAgvH1vK
x0y84t3Qmblay8YyBdyZ+yDXcNV7eHkDLHMUgBrYV6yK+d5yk5+c+u5o4qdMoXLz
bXChimsbb79qSoLYwGtaEOBuBu9G1g3jV6ebljj9n5zy38urygxSg8IvlpNSeB4G
euu3axzP87MS7mYWyVaCkJnYFTZ2h2fD5uYnvuicvYYjioJBs4jMpNM4C6IlGOlO
320DB5SaQgFI+Spd3z8MDpl6IxVhAWMyDT3IgIcFv5aRvJcgk6fY5lGQOmfBqHnu
sa6zTAhEIkeqHBYHxMDtdEC2ryPvHaLzRjRKbo3BULLKwhkgIfzHiglu9aPVXtVe
EDxjqSG5r0iVWkaFx0vcqqrOqVojABRVKQPTlmSi4+Sqb7/Vh6dkzsXpqefIqmUU
PkGhD0e5v747Hl/YY80rdQDzxpxvtIyMUVbJ0yMrNTzJdrqbahp+8fjAByptZDrI
Skpk6kQzAjHOiq2ey9AGiZqACQDZqLNT50DYUbMsC/7n8KOXSR/CMUkdHm9kKM9D
U5xwtv9vDjHWjopLouQGt/S2DtpGywuuKph1cY4jZLcKG1L4WM4fl3aY1eJg1TfF
WBS6nLi9wREGFI3KCVNsCMrTcAzmxsD+Imbs8bQJL8Zp7DvBPHC4Pb05pLD8JNww
boIW/5H0ld5QNKLmplcIBezXMPT6q0n8tu+teNNFL6u/R44qOsxWYEQtU4G0unEf
SHZoU1cN1CJOZMjxs3N1jlONvrzcqz6b+JpLJIAe32EWtu+0N5+ok8EDlMzakNeu
qPrUyEl5bhwS2ukFV4UU8kT/UUwFzWEVwy3Di7MW9fOhUUK+9MRvfIgfPaFx4cIT
feq7dDQMYhe96HITWlmW6WDNrVqx3txq2P2bUJc7QWLSZZZZX9rqP7OzneXRtdaQ
VW7e5/KUljr85WIX0NkgZGy7MFASp3zxtn6KF2vZoxrEBR04Rh8ndE5Nozdf2QH4
v9h+2wm1BMFS8PZ6O3T2fPLsFBmiFEXpxxYtFf/ZtyhkaAQq3Y1Kjxz9KQWDUiui
F+WEMEUe3Ygi0OzTagWxo3MybzD9nAtFmDSliEZjqT1fSurI6ZkL32SwGbozsYKZ
SQQx0RvDNBtt5krOhJSBkehCrYziyCgG0dpb84ZPHk0UmZyM1h/lXezeb5+JmSJs
/vIAWYn5j6B1B7ul5oRHD/keJcvsB6F30WUybtUTi6E1dWDKKOT8uYbYKkG9l3oy
XGvnwnSwuTzZbZLGD/vt2PdONaEK42/XKiWOoe9nLSj9wkHkRWPbeHnEW2PE+/Eq
REmcmDXcR5+KOumvAGdK3sVbmvW8MUKkU6oFl4kq8T9JuZpIiPKgWME/6lZvbAwt
FfKRT48vDTh7zXyq3mpnIjHh/21uRSZohuwX3PiMNCFX6+EXfTMDrM9xVfd0V8Do
Z1KBFYX9zx3412IVZnRt1qCvnR8zbuqYas6TScCepXMxuJ918BunkQ2Y4AbttLt0
wxquAq7eacmvaP52aOVeic6mSj52L+4UJvhvuHeZ5pNh3o9bYUQYXwsaMKciejzx
CMoeRJTTP+6U99fD2wiPe8EeKPFxqN+zWpxAFDtfdn3Y5Y6UW42nIztHhHU4CaOx
h+edeBAjukA2sApT6WuMwyk7xEgcNdjQty7btMR4v1wLSGK2eipd+Rxk8hndmGR5
T0lN3gcb6ffmU4eHrfIEscyPhaxHHdIkqFEjjEiYalux8L96NJuGWbMBxsUS9Vua
MbngBk8gRBdeTBReEr4WBs/i009925kk/wUfsPJty3fi5SNHWEtNnPrcwlxSsxGR
F+jjeyGEO2D1qzmAorRcIzzm9Pc141tz+R51Pi1YprcMgGAIQ9flE3Od136RNaCH
b1a4bIote462OMjtC52JM4njpAjAtqrNKuI3MuC8Cm5e+WajKaEh3waLmAm6icgP
Tb6GLSL4hIAq7lA3J5SfDxQhsXHMNcFCkXhYHY5pf95/CsRiudda2xVtqoASkyT5
1LHnUD0DXXo27wF+f4A//0O7GL2hBLewV6vgx8aaMUE02S9490L56CXTLXAzfKlg
m5I9WMNUaUQkjGld5xHftdTIMSrd/M1AoqOUbOIGRNuguAGeIJpK499TPc6CwKqd
+nv7P0jKaZd8TmDUcQ7Uu9IxsUM7yzcfapEHe8BD1SjDBmFc7ow14iYVarRQsf5e
bX2d2/isW4FKUT3YR4R22ND7vn7iWPcyWG2tpIXwCFkGabJByWIFhAdgcxLb+rKX
tsd5NBfNW9MZbzsmZOr6ym+TBbxAwYaVvCNzriSLNRnrJeFuJRyQjIPaTAvpjK3+
jJXBovdxPWecZt8NuFyVtoSnAoJoOrCEwjA0UzuoM1mB+F9GrDinku0iab49xskg
gl9bHvBKqByB833y76y+6KQRejpyCr1p2+VKOYr1mAoI059lpuPAflGQj1a2FuRb
RSDng1RzuJjKsQqNjf93BMlX7/JGun5b+MxFqnPgvrlP5O1jW0HffEC1qbwshAdz
CAGJc8r1x88LY7ZJsI077ktfXo1D9MMHEXOjldG1ShUBNpwUa+HJRFLXuDazwLHL
XYlS7LjFOeYFlaw9EjBHihusW39PJXtfuPdxzcphc9z2Az2Sbd82MaDg6yYxal4B
yst64CwcraMME6//H8gABma+TaIKqYpQFRrXrWU6gx+D8DlCXoVYaC2u61lHVgRt
4cU6jIFQPxf2f15QykiVG9n+ShAkM8fjn14sNeX8JgQaIoN+4aro7Xqq9wyDwG4r
uH7ucHaDKQCmqJOy1gCRGCrJ3v1+0DTwkdLahY0qoRmpr8N9x/CVRakj0zEM4rJv
h1AmJU7DnjAzbx+AtDNh8+0O8MmLuGPxxOPdlVW15OsAbnq/aU0NE3wTwIVMe9M0
pd906TAMtl+ujs8SIee2X6Y8Qj/vgV7CNakx+vDRcmjrnHkOEJsYVNP4q99WIlYy
RG0xJX24F+yUjSd14S211bY80BnS1Xvu41Wa4wfMnhTWGGx/gnuv3MkqHhXBuYS5
EaNDZvN5uSV2KudkZ3DFJF9Jhh7W3KN4laV2DD5zAOE+znwP/VxJfwKG3/t71UFT
OFovUFcBMBY7Lfx3shzTqzZb8vvIhBiQx2GkKQUSgmxklNz0aU3cMZASXGL6Cws2
NKzqhBXGRBd1BL8sDo0EGY07xQ1eTYOa6Ntqwk2Gbp+ItksKZB7p9ty/di0bArC0
S/xbvhX1p4rGAG8ZA6FmGJovEa7NSA3tIntPiYZ2qcTkI3QdF+15J+SljcYO741w
vSblQ3ax+/herITYDEb83/4LY0A9mqtIk+rQ+/l61df1qyTkvq9/r1iBg8opXBfb
VAk/+YjDsV3qmhZT4NJOXhRSwhrYBWqxdDJn8+5CBaSf2OPr8f7ZXlXKSwAks0ar
Eaztz/oM3pLTNZMc+XmIDd5QPWN/p7aHlrYBS2QL0+9bDt9NIOjFWgBFtpK8QH70
ZW3panOjul2yJrIw2Elh6P/SPPFrnfcvrTuTV9TvyIKwRstqXCRePWmTEQt58eXx
jsJhckuNdtnC5Hkx1L5i7zAwKbLqgEUSIWk6cpjZVq+/x0X69yLC/efm1v2p9z48
sygBIeMvjdTaHJ2vSM5rIuXNIps9UMqE1mzj2KvQCXX1AU7Eaw2x8XLR/L2xixNa
h9vf36ca9v6RApNEwCxYWZcu7731pCKmp9svH+uDwZTUS7RQRInTqW+5MjzAM0Qu
d4Pis7BLimqhRnsrxkQYK5ERBTwsXWFAMzdaRJ+ky/lMn6yu2QVRp7E3oJLv3T5c
M4StN9dPK6fIomZDVwHt83NjBPd3fIv44Hlb6DDb5Pa+E7Ad3JDNHiAacJtk8uqf
NTETVXGsgFjT36+mx9br3mANmTNcNbXzSfLzwy5e2HUQYjmY6ce9rSbRHGv70Kjx
lu9/bs7MXniNRVkqOtGnELCKfvr8BDN3XFlC6pq/wMVUrwSPJcJHLRMnrKFJAkNU
kl1kBfSfTr1X1gqMFrlTIe4+F/PRqOzEG3Wm0jNgfzs0cD6mmuxUsSB5LS/5V4O4
FmmvMBGfNU+Oa3tsPo4RTjbD1anCbb5SksGqxSP3HZL9QXCQ4Tvb1I9MD61YyvAB
fcTcZOTbEQHADMMkEyTx+6BFH7qq9dDr5UdkI5PUxCnboMcAtE50/m0quid2RsuQ
5xty+IFfkpQLRnSEQ+/xf1a8TYgc3J53Ys3eFoztyoV40TscIpFKgjM0talqj6vM
8RWF4Fhx3RhPbcCyuTW3FUwv17IaCrS1UUop/9yeC/nIsy6NGsVHrLLQRkHFpX7u
+DK2/wp/Yq7QomegtqoE35kBk6hHkFcgQFIrIgnKPT0s5s4EbupzrAHv+5tAcfia
Xb0Nf7tq/GMTyGDQ137zMSWgje2RqvIsr1pM0tiK5MOtLfy/ekEqIZN/J1CTPwLG
Au+N3G90e1mk16UzURVXXMELaQNKkU/FW8yyj1FSrSlNLLN1yhloU7BbMT7PtWrk
xUTELwf1QGiAd77Uwpyov6VaGBAh/YiWlDfExbnn5DZli07MZQjSiF9k6GSAH6FN
14QmxrkXj5mqbEmGLyNpLHaO5crbyzczPYngAwXEtxcbUV6igNnjtymq0OyA5jMF
avUNhrYtZ34O0l8PbBjEqfy8ffEwUDQmNL0u+MrBhQmpdxA4/EKiZNHNxqofdXgv
p2vMApFYJ0kQjILc0zxQYnxyZjy7Db2Mz8XilVafeHocqrK/+x7+djGI5/HKZljv
37EW5KLLOCoeHnNMmQTgORudT1n/xQcvV3Gz0MzcExWq7Nv2/XwOe870bbTqZ3wb
VywFwS+FmxQgf3m/YdAR8V+J5Z5MJ620L7vdtnv3aKmwAs50U+8mMo9QqIKlTGmf
usfkCGJqh5D1w1WnhUP9UhrjT3Ttg2txlBOWuvTSn1+WCDIwJ6s3cCXQteelc1+k
qQUSwzWcdsdlxGAiHf6kjEA45YeGWr7Fj3pxaI6a6a2yt/cBa9V3ujuwzPHFRtAj
MoI8SjJ8ayk4pm3SpW/CvezDqH4IOSn8kpcirDiRD6yx7j1xYpm4qB6eDSbYbMD+
GqIsjvMi47A6iyayVy7WzRej+EH5n3zFrpegr0xlbGu480lqRaEYIpsBw0xHI5cS
snDs+dFd+ZQrRKqI9p0iWos3EhA0sdUYewzCZBZwmmdCdL4PFI4M217XGTl8ornF
odCNxvi36KYpkQbafOD12nWbtd4dYjTCa6wdbTDAUwOzMuXZt1Rfux3vSgY1gSY9
eKlergrkjIGVjjn/5ErKFiN51Urkp2hNfu9RStj5stHZsqkc+Cl9XjCZGYMuLy89
r18KhDQAkI+DhLYKO90yS9qQuzhij3yVbqUs7lyMakjFq9ByOouNVY8zyYlWyYJu
/sfBnrS99VcUuuho4gdZRFlzsqb8OGQJYDyBKl3kSa6/+ntcK2h19bpeU/DEhqxz
jR+hObRFxbKVNeEt0BxzQX+hBwJfkAFc9QenXD0uZhi0PTSWC5HCPa374ThWHp+F
bqx0rObbmhaXvQZF1++2UQ15V0oGKcH/nGGMdcbitjwoO2hk4rV7FnSXovhWFF/2
ah2OlBuLjlo04cULc/YGK8YdDvbUXQgMrPYnSXp6W4yz+cbskU/ZvbHTMmLDdwR7
IXh2loljIP5NeNK3cTp/FqXqS5wMSH4lO7aEUo7eGsak2N7D7T0KZ6c1NYp0o0aj
FyuINr+Wxdyiy39Ou5sIywJAKCQdFY8fNuFWFaRgqGkbnIUQnQxF1hn9UktXw9ob
TWmOSgWG+TDT+Orv/GLayT43p77ms4G1oxRZXvIiWPnZKsA6p+7FapRJnQjFPxmm
VyfBGGHArJW5E3WBuJO/h5i999GoVTWyr+zRghu+05nyRjgiJCD8NxRhpBJRbDP4
NrgAWiGMwR/o/Lo16E4LCaYvQtK6QH45PgHTW4Q7HBv/qPtp/s1AjvMzy8zyGcto
fxiT46HQzCRUp5p8hrCXUfb74pQQQYMFmg6mCxsh7i3U3wy3AjbnL9OYoO/uyEr9
6Ko79tkGCF8uVJnmToONEzIo/BYcpMsueo22Uxt9NeBLcECLhTG92pf3tgZZl2Zd
SL475C9vlBl+GEBVQ3ZlBQ/oeChi5IMQ+vGL9hk59HgLVgmzt8GXpiyaVHeQixaI
qKya3p+MD2IRb2SR5UgbWWw3j46PVm/ORBUOv9bHEtPz784B3qTEHVm82mko73ku
Ei9mO6D1JUozGCVvvcWUnxeqZQ9UjGwjJEoIFQajbJnpzxeOfsffxiX1uMxrPdgn
zlHsLVzDPwgjU+HUwlBVe0rehPUSgS9Nscy9hMeXVBxvLTZafWcdLvX4d5KynA8h
WUdDp3re7EGLNcoCUMDS7oiSVOQNvQTI4sBm5QOUn/XJPQcuvBauj8WOBnnJTj4A
dJrgXFowyka3/ardbclZK/AwOXaz+ftgaqotS99vPzXKbPSN7IlvwurDpv2n+BlQ
mpM0HBexJr9pgD1z38w6tUTFHPLdP+ucX8SRdio2fvbo9hoN4E9xk/2Fuv3kaFDG
HeKEUPH94AhFERr+HBy+4pxIEfAd+z4XGLLUdLKNNpMETOholuUowRxDP90/9f4w
RRYtuOpdpqpq5ySJ3X8ME/P9ULhjRWN2d7S06s0C8MN5r7EL6dWTJwF7V39n1wAR
XdcehoaM/aRios28G1b0n3jxwCMDDmcDvb979dRKPIQBOJuHbW3JAzqidynKAPP5
jZ7kDrexjgCvVLSneeZzlDVJOeQw9ovyx8NSf48dXD/o6tQC4hNePy0Q/7ZlRc1r
xPE8FPtb5A9xMW6j1D6o62GsJpqzRtPeRg5S/OD40Dk1g4ueDZ9qYEL9xHJlb5c2
afHhoWxWvikuTY94sq3LL7YNu/s9kSz4Ru1AVjDSrDQrjLZshZaj0CwzuJ8YKl/e
si9Ixw0QeURnQv/TBZHe79OI8I15jNEfQGvFgxoY7buuwpHFE5h0FDv6WUVKhEa1
7B/VnbCxVNqwtEJ3Decieuc0onnJrVL9xavs7tKvBMeHC1zbC8m+n2lLOnqijpTB
3jHK0OboPqrq6DZpn+VltBxlf5M8iahlOVjyITlGD2sr7yarUAggqxcmbV8pzKg7
B9PMCVs2DGv48G3UHFd9cyz64+u+pU94Yk9+hyg5H+v8Uk5z0IXMgI5bAWapZBng
s1dYdlrQhwU3eJrRJbJ51wNYBqb0J31I8of6Nl9aVuKDHJpYjvIv4bl8NaAjsjo9
QPH+tZQIQBb8+jQeqltOd5pkK/5fASRLIaFr1ca3VWsCQwVq91kTa1Swploxk6Lf
zePTGGkkA1W4BqpQyMb1ubXqAQNEW7GyTU2+fdZkG7h6YdMKcTMR++hK3Z1pyX+p
+6UpbGbHsiDBokh/5FMlGuLZomk5QwcT+oD62xg/e0xUB9Ma1nx0BfctK8WUjCJH
4MGQm4p3qw6tvyPJ3YUXDX0Ov3leyMn5xMQfN9ZddEW9jppRRMFu2jm/0Fe8z8Wt
NB8gMCbePooyrUwEyenfliBeTvPr35fMH1GNpQsAuOoKAQ8RO2ZVrCAc4gKjrIws
OSt0fwigwZxtmHvUTmqNUgTwgRpJs5Iadal0I76IN1CbGaeFsPBkOyfHhSRWBpcK
XpFDrOVG9lKezRyU4h31sC10EZ5+uxjO0GI1d8O92d8qikJIjtAGOFOBOV1c2ohB
GtCCm/dR3Lqhx0Au16Inn6t8gKqw58/eOs5DoC/lKF3A9cDRwtifrYf3on2CAQq7
GL4NpL/8tYhS5oxgp8V1shV/lQGjfFrktgw8MFZj6U9ma1mBJTSFJkP8p+vpeow/
TcMxL2o7ipjZFaExLlmNf0BRM5J2SqHv8VN3dLQszf57mu4S4ZNAlH+cawyxvBzh
eU8dOkgeLLs/OqzhDIyW6otpi7reV9T+l8ZmbDPVo5FOZBy5fSO6lRRpUnZGXo3y
OodqgRd5DjO5SmqWqWJsXOI7x3aoTe5c0mi00+q4zfbGO2cej0TG3Oz3qgpYefa7
SNn0aPkVJuj4mt0SehpidbtIwWnXnyrTK231GziMc9T+wNFi+zobKrzLmfs2Yu/X
5sxEP7PYlGZaOW4ZDMr9uP93CehsMjtZDKRFQwMoMbPBHL6mssIqIxm4E6CbcIZW
Bw4wi5iUxfVdjxe+176i2iWGG5kYwXDsoLBFHYly++6YqA2tHhHPO8V7gqXDGdy6
2l+gYfGB9/ySACM8LCLnAnZzHcfdQYPn+mU1CSqtXxnzL3fDt8pX33QCF4A3O36T
x+UhVsHP9ubWWrNS7VOKwUDSOhzbcGlye3LlSPEosxWYVWCqjxHqNv6/evZjJZcG
k6/Hcp17zhCqi+qTgZ2QtuMAmxpf9q35gI7MSH/xP84o4wUSIl63BsJckVqcSFsz
CCvBqIB01KDgh6iSP3nsz5e525k9SpOHWibmiMbbg61KioSbEOJG2zsKFP1e8a/C
34iljtie0lAFrnVxSXwIedvF7BOcwEf1fIifYxS2jg14e/zQuwhy/Llc7AYKt0OA
1Zg4SPD0fY4XD2NmtdLsng+gvVQdkRhb94AoxClfouydJHTv2Pz4kSEjV5SNOE5n
G7rhCbcuiGqV1J0iB10bnapphelgIthqCZ4o7VaZBKiqeIvgNygJJ8RgwArLwQBR
eu14oHa0TqAW3em5dbzNh8EmNfkFghUAZqv8hz2n7LRR5vfTw5e2pJQUvjiXhyzO
fn7Ns/a1ZXFNTE2FkEIcv/Gx/t4wm8V/WWuQimW/yAfQcEdlAEB6vptJt9G/ptNw
ybnPW7UbceMwvlnxfoxEH9PaLckjiKZUZmy0Niz968T8JrESkIxMSerC397itKif
apATx/wZsIGfBlZlQRjUKGh5qBTFXr0WJuwui/cq9idaztZSXdq7EF5TzRWHK1xE
e3Vu5a90HMLAZ3e0L4afqCKg0fFREWbSjOq/LdYjxQaJw2ILQxxTrwi+u3Zq96eh
ehhoFmr9ezJYNnV5na8Fcu3twKlMNPMaVFnJwW2JE31GJd7adbKSlfzYK6eQih1S
/CLO4zfig1mG0DksdC86bR5EtAE74/LnwhzYZJpFCKcZbstfFNPxD9GJGk4Txv/M
hHyGc+pjd7I0zYxP2eYHmZe7SY6XLlK+N+KeO5HkUEI41ZafvnGtMf2+p4RXsA5F
1ExGj9nPGeBqblFSZhBbTSqENNKH3zY3hw3fWrNoQZs7lsUG6hU5e3XnRwFrrQWt
bcOgdyFVRb6Pmx5ISAtmKSXVThLCH12nuIWSco80idGvb+7R5KiHLKWLCCaOnpUh
S81sBFgg4YhDq66zXE7T3GP+oukhTFVxHZQcW9XXd7W9/oEgO23OvFw3gi17/Bnc
SCEuGwsGmB8D63aEu7xCs67a9KUrYJbWLkSuLhy4jFrfuMh4srpKj7sI4R4zKDiD
DFqRg06QYO43xtGAdFq86edimiCSMmXALLoL/VtRupHuwxt3w0qrQ5nIlI171cnq
oQr8ObmejRznoaZ5qNHWQio/+NqkANRcpOdRutNAs1zeIDrXM7gPoAR8+zt41D9n
9l9uX0McwrAvCYBN8/IHYkiSjtjegxj91nmsP0hG1PisO4WsxH1xpFNCzlh/yJEc
OwGoSDkeKcCKh1eJ60zjZ+rmi0tEtDU62rBTGzDTHDaDxw2o8lh/Ka0s310IrZaP
HK4H5xBjHfLDEMfsaXauouFP6Ftahb9YBUNoB4YKeXZyInPN+hiIm3dSHNMzFD9V
Z5mDpCxKWSQDVg24ynSHo8RR54rsJGM4ppvfQKlX2qzmdIHlNTvF1rRpXzhrzRMw
1G8zQCyG1/TzRtYJrmHsqpcyW+C0lWaaSYAw8odbeNN5xAOnusLtmqdyP2e5yffu
36ZVMfw0YQAtb5GPa3wEAo1oWd+aJKGm2DE0e83vP87SiQUBUyd75OD7hp3SxJsG
p9Iqip/bOZJeRYJX8EKI00FqlPoRWYgqE62jv+imkzgdAFLJC33/mD8oVFwvadSm
k5vJs3B7dyg890Angd0+HatJm0Yz7z0Sm44B7Mh2H9U2QUjvkaO0K4irCwOg2w11
kyfBN3PR8r1cNTGLaqpSNY+HRdiP17PrWoMxyPr0MOJW6uqP4HbSZz5gIW1s1gkz
MdPWeQltXoC91n7S2w+jSYJ0SmoXn6+MlWvUUSIKRQPsGwFgKfWmVWeT72BTN0or
MIxdISEXrozcaJDlhDY7ag7+uuMIcX3xlz+j733Pzdz8ByJZCmzkAsoAuSXd5HV1
UzWvTsFJrxuf1R3Mtn3/zhcGJCyr6Tr2C1DDBi2V15lsDtYL2i3LWhnDJHPO8MzD
8sFoKBW7h+IZ1F3febk+CfCv6oZeekm/Q7z/HzhXUEd4n3lbDDVBOvKICRNZRVSv
Q7PjqSbv1Hfe35e357solWbofEtErXiADw6w9eRkCw26sy9iSuzhqLDQ1WmtKPDi
Cq8Xu41Lv2IsOfqp8miLyrpS5JVKi7JT3o8ByjOQTn2Y0vm7iZYcUUHbZURfIT5x
HJHO+a4ayDrIYqT2Trx/DBfOVRsuz675LBeQ0aZaQxUfYpKvCCbQZg7WBqtkFHXP
q+R1FtmrFpFjcmIVUXH/F1YwXVmsN/1lahwpsVODaFejH5KTz1bm5ZncJwB1FGUi
3czmBKDe9iW84uPDfm5bQJWznKIeydzC5wbOHBH7ioifQ44ialwYPzo1mer3y5Nx
29ivvtkB7+QMSBjDU/ZSmvgKiVq53qDiy6gdVgjiQpNjpLOWEmGfJO3AIsiMSrvO
2/5YD+o3pV2SlXw17KLpmRefQWn5vFkXamOPbnHdn9RGD/WV29aoxu0Puix2vbEM
rcQzYNz6F1+gZ8x7dUAxKjNZ1p4k3nRO1ytcOF+wLAsIjPUTaO+G/bGxX73wq87x
/XtN5SCknZtUunBf9lg1XHaFlIVP96WDnXTd7+K/Ogc4jIW/Z+cge3ezIVVCPWZd
oeWUv6b1/b+GB5kKSExV6+cUz2q+Io7xfx57dotBhpOc1nJtAgo5iBUAj1VRzp3i
h1GQsYABhu7cgtxD8Mcbh/9aOo83lv9PGomyucFkKPBQhaVfxGfTXGate6Drqgu9
AV78HihDLo3zFWCDLeZ4udfc9ODtq7ZXGeLX5g1cbF5o4r0JviZxL3u0RB2emeFF
H/GP7k7pd/B40w0gKkyWN+ENU/g0we5DRXP6fCZOXmACLWSjqiWXdzWWiZT82Fjb
TwUusNBsljLHS+vdnixrPwuQK10uS/i3FkMo0qYBXwRZTUBbNpQMp4HUsummtn/+
suRskEkqXAZwk4THUFSAk9rE3f8cMDwbFS95iH0woCQC4IGY3qFkXshElRPsAJ3b
58CTMkHbzaimLzSpQ7QPbIN9h7jgb9AJ8Vb34NvX1skYL+aM+ooFqbjm3egxAKvZ
y138yukVsaMu+dMKjBR1HMOG+1PFxpCwTf4r5tcVfnjtMDNHds7EO6Y5RfRGvO1Z
nZp/7valMhUTDIjtodfQwa0tQLR1p3UJICeWSAWKGRk+PxbDtbrxotTBfsjPGoZ/
5NeYa4czJbBUy0XT9P/kbnW7LdT6E0axRAdpgZ3O/WIlpgkQgbrHKfbDHTtZk1Rr
XmnrGjK3H9N9YSCgzefxmGrWQy/Q3q+QKRLGujALc6bQbxltUJpsxpIcBfRMtCls
Vp2BwUjzBifKWzrD+HNnQmoveF3Rs33BRnhALiFnKO1AwnrPHjtTttCv7N0m5v+5
wrecOSlOrP1o7KX/5YJ7ACzGF32J0XUsyKC7XyhK67AkyA7l09cgyqBeOjMYxokR
Ui6VwbLSQpjwGn8qovuSSA98SQSN/t22u7TD2oEcHsFB5tVTfI4LPQ/11wwU56fg
fQBNewE2Yh32DDgf2mcs+E8bgDnq5Qv8pfo4PDkaX50kZEps9RphrYK3vkVQlRNJ
o4HehQnafRukvBxadTc+xOGTXKy5MPzExwB8g9+QK+dHhqFrG+I7mfNfKPSeyyK4
9GA4P37u1qvHzPdRJXOv6B8Q7N7dUhWd+3Hyru/pL7TMJjh5CUPpxgSPr4nEE9rx
isrBCUf7eIaddCEGvPugVMLI8WR5+vvT6HxoqHCE8L1GnBPHEhHbQ5MvQGSJGpHS
v+wEj80bZzmICbO03UdgmxzzNUW50dVl6/V5ALRLRfX12bSArZCKQo72YUF6x2Vy
dNVUCn9ZOn3+PWpSlIbZxK4ZmYTb4EhDvYrTV+Kq66oG+eAndXeU9cd1DQo2OyyE
Dn2yIpjUGiZaw57tCAg2W+JO0O1DPBehhyT3QvGOfTgStqr36kX+XaJ2mXxQ4/6R
B/CPm/0R5IHH59vMAchBo/qm5MdCFP0aZ3ssj3jURXyqj0M3HwbapL8oE2VGWbbP
/ZRVSJ9Z5Cm0u5NcRoTlUc/MB8rMz+OOwCy9AcSZPJR5QwGR/rIeM2AaGpnDICh9
+MFpAIT8yMgSo4XYph6unrwW9JzYuIEN6WBwVIz1ChLkxNbhb9C6CxAC9jOS4z2u
I1pq+U4AT2ebbuJNBSefAjeGr4f3qc2dss/xbsQUctG2+nwiNG6p8z//FKe1KWO3
hL6HjEpsV8HkWlq582Y7vf9Bw4dhUiN8fpxJ8QZBBTQHhhUWfhoBb5f7nLeX0WfZ
8vU/pVaFwuE5De9e7G/wbMlAFPIeq25w54HItPOW72fls/BJvfkNvB3csGie2nV/
lWDOhp2mV4VPCPHx1x5NLd0qiNrAq18AONopJA0iJ5LPPX4v6PwCZ7xWjtLNnNdP
H1ta8YZ8iBm0QnlKJ4AXuGy9aIxRs5nI/tViC1C2FhNswrWl9JzH8r8Nqgk+FGUS
mU0nCT0pm3qAJLdMlBO58jdsLxRMe116w/XhbfjLOQLXEmMFyFtu2DHo09RdyDij
6ryxgGOkpFi1cpsmGJ7VpVWxsiTzWG5JQIkJfFjnglZDSVEdPrPYLdrO01ocdXdq
YqAsJalxmIWnKlOZDZciPB93xpNsQEHWHvgGKTr7Zx6DPiZyTcEQL7Ky8KVU3sSP
eVchMQpYJOo4eP4EZPVzOIxFd1N3lmfjlPbjJonw/EmM1VpLYPh2Nhr0Nl4/8FV/
xC2tD3e87MrARxQMaFtxYSfpO6txU5ky5t2tlC23G6EfAbyy0BYhxBUo+Avqc4wF
26ym7Fp9BB0qgKt8BYQk9Al+1BvjJAj8H5fEFEcW2Sbq6W0DOjNwEMkg5nDJn5cT
+WdV5zEsOaCMEfMGVZbmrCSZLP0ykTpXoMgtvieIFwIRqfKoHLZXl9CgnC7hf0ed
EdcFi8hsW9Ywx+20p/TEvstp4iy0BYpJGjf/Enolk65EkNU+A1/mlf4+WwutM+sV
y/FPx+vgrqoOpLEj5wxKu2Y2HSYawpyrhT3HCIQxBUVbQ2V203+MlsmPP7MZ5K3i
HxbAz25KeWLbGRIomZnRO8KSXHBKfUmmudL0wTJMafog3CuSWFgCrmd8bLJDse3G
qdALKBmE+c74n0W5ch/z5BmolylV+lltsVcSD33gFsnlz+F2lUJlEbSsoxoFm8Sq
m3p0qtoFcE9LpXyqysNrNJxW8FLhR1ZxZ6EwZY9AOpXdEZ3s5ckj7ndu9CBpvsst
lMDnsztGWfxD5dZrTgZwRdrrJT+39o0OhXgqMvVEhGzpGJCxIhyiBgGfZfYZaR8f
d8Un3opKMvyK6OhMGAi1G5LfnHrDdamu0mIGvJeFwYPcRWkpZ3mWZxRyzEBoOVg4
LPVwqlQep2eZd2RtgNM3dtDcMI4nr4L0Xs4kcn1kQq7HOdETuNqmxH8umsC09TxC
s2kncEjcWvKhK3X7BTBQHS5RmZxq2dop+4Cx2PfL4VNozwDadoJavDFgx2kRVNUh
nfbnAMey1eIOBo4cT3By7QVco1C7Ii+sBC9pOQStOWfPAisREeKscchvsfpZJXNf
BLoBet8cheCCziCMtq+VDpAXrJK0xcPmggY6wdh1j1krpIU160WQe7ZVGaV3ioBr
538EHTra3U/pEjwpzYeOMwekhlhTGH3coJyQlvRTgB/jdUPMGMuPg02Ie8qyF1MI
o+01N6PVnKuWip3jXtw4DTOYAum+DlngCb1YkGd3euLcF+uGqx5qjmOzVMYRmn+l
wRcg820zEFGXL+ixpk2xHtFdBwai2PR+J5EjuoaU8Rok6j9KSiHgUupZ3ifvDV7Z
q40Q+nLBGDoAGF2/sQZHFaR3sPiqJHu5tVYXDFLUDegJguriskEGmaZLkfWTAEIQ
e+1o0AsY2pUDkwDopCllAWQ2Bzgu5GihBBrI0ZEytVOohaTtBldGYcOSSqsHmPv4
DirIO29SsHWoDgP6eRC3KWNxNye6uI8NFPQ+kpyKojZHevUj+f/CH+EMTDMLxCq6
Wa+YeFDOqSPPBm4XScJEtNI8ByfIsd857bv+XlbVHEGXA2dVux1l61/mHUSIfnRb
9cyt4K3gZQSEksPbCIBsXAEyk4nbU2MUFgrhrZCNQpIW5R57VIki66wWhVU7CDPA
Ip9/JAhkTntg7DS4c4AKag+Ob+8nAxfIto5XkdfTOwLS8U+cSXINJgsQnA9/QIqY
wsUnVDbiylH+KAk64xVlkZqy25ldAaY2tXqx6GenYPLAv5/ecRJZ8h58iIwgdvW/
w0qWRmTUQoze98BtbjAuIqrwG9GEC1GYZRUKwLjMF48jWwJNImXIb7FVKf1/C0tH
9ydcO489t6hq5HEdOLOnUIKT05jN21/rsoDiy8YZOflWzfnlSb0rLmD09c1t1r3S
VbMI7mHSvuH5S/GwI7Xo7V83aqb4ADiXoP8OmAsup39l/PNgYDKR/GbdjP5qR6b5
1Erpt5LMjchSNOGyuZlW9TErNPQbfL9eJK6nUd+9VS6wNukmwc7J5d0jEAwSTZjG
98HIr4Hk7U60kTKOBKsIxJwpql1Iz2XR1/WkgQZ7H/6GV8rol+cCCp9AA4yxkKA/
TGTBI58K/JGc4mlb2bXMiq6C8WxPMBGvc2xCgnLCuUm7oY2ilZ/if2uv5o35003a
YjdKbCwlpE8hokw+00D7Lr6d1IoYvoeuLHVNzUELTEmJoYIl/E9L3R9RYvS2JTuz
+7u6GPqMUkMAJvvVFy57rU8gjOLoVXwNUJZBaA60lGnO+ZLwFWuR1Mwcz54d1gC7
hqe++spoFhkgR4pRmnT/7L394Y8a7Ua9OF9+7N3CgZHK/PLWAMFbtNGYfRQrTmvW
HzN/P2EWY0INruIRIQ6iH+9VeZoiDN6kmuRA1FazD14M1Qf/ym3HJGyha4bgTgUq
6VKN1lIeZ2A8z7Xni0tiVbcQ0CL5vMLSGA2GKnOocyJix+rFku6hVWazpQ+jKMhe
U4Ph5ZxPXVM8kpBhccfJCBcJyZLTGBdDTgn/6WnP8IFTG0D4kkAtZuPdB8udHsis
wz5rc+Cv1O8iePK8er4RA48R1xI+QbZlVqe5bsO45Vxucb/JbjQw91WZQdk8vqbz
A9JXaQLkcp5sT2411fbRb4Dm6lM/88qmPjhrfiGuXNR7rXD7+Tax4x4/OMKuj43V
K1c0DrLGrdqUrzI4YKm9R1PcIY+woSeiYCt+pJwJv8AYMpYNI+tdIzZAtH7wwsld
C8hbY/N7BBaS1gJEOc8XmjVj6ROCZWmbG+cPAqzi8qFqmBbIZ2HOGB2W+iiQUWvt
znA1LW1wA/sq/+ipJNp0SpUj1Ma7exVqi/mZ6uAgM4o5J5jjJOoW8vqAxyTKRz4J
sKeeeKsM9tj1RGXK9fLk75wB0UsHwECs1sOvFUn0Qzg6tqHRU+ubq91jKfL+bOsA
Fj3FFsVkwPZXQB+VsVgN1hSl38MgGQ/BnvYnx5Leixqrvshpc+8ovTbncALASYY/
iB2JdeIXkd4ANJCVbQ4R6GEZETk7AaNYvihW+9wWHqXcHSKboJMwRkR1iBloLPyE
tKWT0OdyxDGr22IvWVM7c0NPGa8Jz/QX7SRtOKwAz+nicEqZ6/x28BzR03Abgt58
Q9I4fSBUmafb9J3eU7/JjMeSK0RjMx32bhlyHjZInoYI+YVn1MChc8ai9MO6T8s8
QXUh84XdgdsOMgVDfs+GzbjBCHDFp0mFuhFexrijig2g3Cv8tsTAtDYNiw2UHx/t
1kz1B3jPNUrS1A3M6jAtIXpu8SRIcjmWRj7D84JHyQjN4FkXy7RyqbyKC8tUE5TB
TXGffX1NCEE07+u9eOfiNmp5hg9i2zgYpB2BjZuWDkS9a2w+N+R4/qwpbYhrtDWF
JigNO/60SevnQlMjjq28LghJRvdE0XYw6/iwHeW4paqccOMwzcy2v0HQNQHrmvXD
3OPo/ILYBZcXhJYk2peaA/5tuJPItfhKx4kn6DxTDcu5toA9qNax/V0360dYrpBS
2KNPbEDIfn6qJmJEnyS/UN0U8Yxri+P/7jZsk8RUsl7QGLdKmSDX8TgJjpS75yf3
puGTWHpKLZylar0NTsnZyuuuRsqf3i9IyQQoSenY7TFy+Jx/2/elgNoGlIU7C7XH
/lmBVDaNDOzrugN8kvUGEwCCHMkzyq5/6ydIHNuPToSxf2gJvzcHCvTQmCX18+qw
upGiSGpiBcpRI30fwF4KOF7DfPc0vT/taPq4mEZCEIck3BfxGvvtDzjEsuOZD6DH
A6suyAMLatVv2iEoXb1/MrpvdnCMsbJ811ZFAuCKUWZWBvkw/QOtEvXkJCI+c2go
hByTTybUD9NhAWCk65jPiR6OQkD99h/U8ODceagAwkVTxCYxkElLomoLFM/6MFIe
JdTNVI14vUeWIpo3LAAb1Nl4PgGmOXuQso7yY2yJI+vPE93zjj4rw6r2fOUQJPQ1
mGiuEb/u51jJB65RWWn06lAF/9Y2ovhWAzddVP+PsTdfP85URQbwQjextQyElucD
QSlc0DFJ8/NirK03/iIGA/vJD1LOt6dOq5eKPQrQQcLGYKlJ95/83fW0iiKsoPoW
ZwaaJKQrvMVYmSht1shMSlxEkojwyBXElsG2M0Ii+fHXqGbUW2jaS8sFB47fcHfy
zAgIeoAJU36Cc+UkE8S/cRm39kgmxbKJYSCmRGk/P9I7VW6SO5l1ysYEQYeOhcHj
kXZnJDo6k/4HIawzOnueggEEI3Plpsx2KzU+1P4FZJudQyW13M3oSHejfkuPwgrS
o7WglmbOwm/qqjWusnDD7VbtLoRLFZfprZGTeh3BvK17d3DzHeZEr838btc9XjqZ
OpQmJyFmWU5iWmnoD0Hmq/q2HD2m+gSDPTaekqFw+5xcHiim9fBUHQbGRAjVMAO4
lIMAdIVEpk1xxVDW67O2LPCPXHdpA+9UwYKeuM1VLzSLyG2Yazrg3pDD8RWr/w8W
9PtPo5KZu5p4dEY6X0gwM5/NwjA0PJCC4lW4A5F8785oi7aolCuX6PQ8MtDYmoyQ
aaw8JjFPVCIom2d+IQkDWviS6GDX3x8FG8TjiswefxFAt7xN+EB5KOOXghwZWUq0
VDL5aw8xjqXnk53ZfYkPcAwgIySIBcTCczlAFgFcj2+DBk1pEhVPNU2Qtc8idTxP
frTONOHVnzXc9lr1RYtCy18ttmbsiY9/Pvk3dpctbgDZSqufC0nzvjpZagCzodSm
AkYYQise4HVLzXNGt3zcUmgEk4dTPCoOF6xviGXfqUd856y48b7D66jerZ89Ej8C
volml3VUV9mSDum5Hz8q3fRg5eySFmVrVc8hTMYxt+qxubacqBNlWiDFWQvEhpij
vXhS7QFHRSY99gKklpGjmM1lqQXYvLWZhLZb4bQ5uD9EwDwcaEgVFpMZOL3LNlUf
B/L4LznNOLvI1EPaZgespi6aHUYwYDyJb5JsLntLgqRiQoinA02I4kndWY8BPmhX
aCGVRr9s6fQLEk7kaBmeoEW5P5cVUhxAqB0zXp4v0k0Ne05HfLewDYTWOAhfY+cL
8dU6qD1Qz/6w+ZQWWlVs4pUzwAuqZWo9xJH4AHZ39aNUZuGr2cPQ4WKkAPK6xA4w
douAHLxd0YoMgraffxLKypF+Os5CIDcO1Tlhj+aOKZ9m7HXBTG7HCmD1v6whuswI
8OCzh5Ua8EBdA12jDp6VdaLyeRaeVPn6xs7rSAlEJKaL450uDscnDpjg2Iwo1WCP
Mh8ojOJuZHjs01TyGq1Fdc5zcN+X1x9D7BvepbzzUwFhO7km5gcS4rg3KRntPjhk
zc9LPXjkLRE7e1n4/wCwT4hM47cSD4Dme6dTrfxawI1KLdyvANQ37i9bz9dhY5yw
5TFfFsyewJn9C+ACH+oi8Oc7B1LcaGDrKuNY5RdBsZuzaN5CNkcyqq+ySXr9+9Fg
oui9j2qUL1Wk7Y+p31kddgUmNmVJ0/h4OZn8hkNUT5C9+RHipKLilPOU7st4g7U1
aILeNuBYI5bl+cFjlkQ3qfFbSX5GfmR8BDDUcqRuBTW7heyGwYr+UZLkhxtiqwLK
xNHphy0A8mSoFkwo9MiGwtal9ENOGH5xQphaSLN2d1cT4zSvqxxR12LqgFokEPg2
5EgszqdpgjUZGuGuVdA15UCckKVm05Ul5v6nVEKQpvdX9gVUdUVaHjpxXe1fd7DT
ZM2RbppWoZWw8EE+LGWJ1r1f9zB+3FzAObNjUp+qqH6v8PWIHhRTdN4ffReeToCc
Eib0qwbBsuCSDcOcNkPzYiACQ0Xelfhxb5xXDTpHXj3Ncj59K7r6y3aDAlyAkzvF
GQXRTh0/nlTAaZ77dRnrntk0MhFtKy+QT2s+Qttr/FuCN/A9W/v45IyJ82zAa3KG
NDHnstMQFbD+NoZsPyYwKv2A5YXyd6QrxBL2TlL3MxpCZPkqCNgyNeNxkLMPEMIx
upBxze7JJcp88Zuymc5CpKnw6mLtSpcNOqlUa2eWLH72Q5xoTDyT08eG2OW6NYQX
5jxIfuPTAA62sULYUVGAlMjNlGZmaxBXCZGY39iuinr9LpGX+/+/LPqB8TjMPYrl
L/T54OrzXJSZ8TNyeQ6ObDmhNUnl2lxprghDYZ+2KLjTXQdWpj0EhLOqgJhkgHWw
KEQb7Xkd3VD+qayU0ok2PNpDSG0PGvo5CIGjWYgSpZmNi8Z09eOJucIMZpkF9M7L
PggDACeW3eM6NSmM7aOfevhGLLvW0fYVzx9CIt3rHTsSVq16sKY863j+7U1yzyd0
BWuKwNchhjzdYxuwheToYP+sa3lOsEPw7WIyTIHCjIeZBaCwV6EIGnmbx3PrcAxY
CXQeEFrCW1hO82VBj4NmhxqcjOK7LB76cm/yPiXhLVya9n/K1ChjCLaIgbPYfXfI
WDi/+VMJ9Pn7087ihogBuBG3ppBweW0SOlVfQef8iprdF23U5Yoh+ybHWcSDFC3Y
x3Q1DD8O4RbfyfvirCJeIWZI0sBnAQXNgFC9/CEUh6Z9YPvrcpENKl9XZYTtXLvg
Yg1xnnqmfXd0ebV7Me91TKo4Iieux+pnBJpJKKB7vukZPF3JOymMXHgjjX2owHZ1
rnonQKWUjlMHSEPK9cQ0iUEIBYzKa1Ts2dmVUi/jQyYTaZNWYEuDvdGDawR/TESV
etZ3pynEsRUY0aONyoTgYneGU4j4nggssGjxaf10SAnFeJZui79HTceuNxNo80iO
xxIejzm7bJq5UV1yo6yBfjTx/xXTPH4I72DV3A++SileKkVUQTYWsKTGcLOWsIof
EAPnMRRR/A81zhHvh2+5s22Z7H4hPF1aW0ys9Lc+Yrw5s2Fn1dA6pzFD3xKfeHdk
rRJY5G0xJ+awZjyhAPLoegqfOgNT13qwe5hwvh8KDrJFYdLyRHPw3aQtFPiZSF51
wEfMsCeoZlH+T/DRgJ62cOk5mNEGfINbhMRwrm5oco2VCYys4sTKCMWZy2yFUFk8
ZCp5YuZssXLkUG79uABFMOHXS7uMseJMIQQak9OtsFTsgAN9W5TdOU3chW2dtO4X
3daFCimJ43kkDHAvWgTSx/Z7S5VeSQ8QruZe1ibVGDmOcbK/qj+t054c1y4EJUwW
5lhCcIh1P+Aytp2QSB6lp0J60vTBimrS5ztC53klktl+aGRqyzQ+b4E5i8wVfkKy
dXDBwSw1TmBdELoVfMzvr5Dg5dx5S+ZCeDtiNPD7P55/DFDwQjHfazHCV+VU4x7M
x19PYVamqiBVjFLmYwx1WjXqU9FUPRr3hndDIq2b0MDFHxkAe6jpdYvrpZsjK4qy
lfmOS+O/ahc5hLnEoTvJvRkAI6cnXKX2rp8xHzfGKiV6z3rBUlUYA/NnKTj5Kyqx
Eq8Tj76kpDBzuggf3Hg9zdfyFw97PCTv2XT92fbc5ULBh6UX3PhN2A03kKBee1sj
5+lt44DfdJSMCdgnGGDE/W997oNLFGNN7ztWrkuf4VacuyXWH6IcwKH3evSNLTGH
GDIpUQpN/XwkVeqsw/mYWfGgm6XS1oiPcGCBts6VH+5UQjN9Xl7yUO67O0jfsQH6
iVeYG3tPgwRYXAnZ3p3/xM4WnbR5puO2BSvQDjjn2bsPtT+bOJM1TllPSIckfIQZ
RQFcBDDS8i462s8FVVoMVv/jtMYtQV/RGgNXZUkJkz3rJ6EvfhcLKN2vXDlVcjum
FUmonp+01OBTgGHy+sojH8daHT5UR12h5VJMk3eaWHNq7VHWRZBHVGCoQs7vqkJ7
Hpormn950wfH4xLeb0MJocSaSkasYZkQcLLlumPzHoR7DbQuaQtwH3ZhrZFZH6QB
T1aC6R0B+ifqKSOJ3l53xYTb51Qz08er4HApNXyEx4PCM9BnY1B6rVXYfNO4Enx7
+D3rnSo4Ij4U+c9G7dUWKG62guDD6IzIPStz/0gb0XKxLZYn/JZUFckQaORDYCO3
BTmBObT/HwMzhyElrB49vmR0etWftzElHPQTqULAcKMTv8nTboYXf2tZqXD9amH6
KtavoXePSNcH4Qn5wVO1x88MEC5JGSIW3IvFSoPzU6LLNHu7UWv2yUq5pV8ONOWg
QHktm2ewKN4+Uk+spvNZf0rsohJML+na08Q39S5J4uSvvtTXgM7FcnMfmGtFa/Nm
28YFnfrZV9wFB/Le+uSf7IG41Ul6kk8qIZo/zq5ucB/n8UFHYkieXnCugOljweir
MMgJu9niniqxh4J+GpZuMMcnX0c5qt9nU/KwGipIyulLmGuAna5h/ol6pBGhvgKT
6t9YO67NsSKKNI+/fDaug7z0ir7QS5eEfjyVxYUiM2R22bTmHAaThjB7B+VfQouz
Ht4ISkPBH2F3EGkng9Q6MgbwWM4Y0TnPu2mz1AUCS6CNAYNLaooWf5mCqN6EK7q+
ikZy3HypMBwDRsSioCai1LXOSRPLurqSdRJvsFbOpT55ANZR7eX2gQhtRPTiQuth
8JvP+zssnt4ogfGrq/uYtTIagY7H1bzz70qDSg6YtK6soV+NYJyzuVJBhAx/2sYA
BNoMnF0tZSkwEZvKkSPtFwHpyfqs48FgxmnG+ayCAFqBgZ3d9b+MHb6QxPnu9lr4
UMd9Fy3m3DG7ZIdrj6yGGBxPa4F+EE3qFSfWvGfZZRm6Nq63XHTIEtjgxEBRnZLl
BydMnDJifVp5hy0O8b4DVwFjl4Mdug6o5r6NYkV7wd0rbXJyA0jmB5QHxsLOwAI4
s8jakpthP5pOevbFNDfjVFGGwJK6PMh/IMJKqOA8TrRiVd86l8JvLR7gS+F18hM9
FF83PExwd6iotw+oGPCy+EnR6Ox+9aJZHa4DRxMKRFTQb2Wg4lvIgjx0YTKd1X9q
TeiUDIITHqEsSiFHSOtmcPQXDwUL4J0z1D7Om6DEf3DQjtoBEA9rRfTtXV0waESV
zHM1xysdmmp1p7YbRox2QPXwLN9bsjpy/KZmaOCM86O90j2sJFYpVKTItL4MMJW/
0067FqNOwMqkW1WD+lQ9knPcoXRt9nByMApDBuvvYp4EdYykcWU0dsLYFCpDkMrB
HtIdA3t0SQ5p2ZtTRNWBMVCkiXkUcexSEHJN/wxysXWdLTVlFBwexcxQQXku5G/s
6Co8S35LE+V3TPjDJBU+Ayxgv08kdhXNcfhwOwfwDfpLBFf/E6zfZhuz3ctVFFBi
uF/wzHN9NWaPDoV8JolfD1DQ6APhNbr4CBCs59e+yc5BcqjcK3V/K+yiOag9muKs
AtO/YiQ5x33Ezwe7MRPfemIrTHwfB7OlAhh2kpHTCiT08mHC8N91gTR7lKpcGtBV
z2GyisowKNh87DIktrqXQGxod0AhT/GOyd9q4Jf6cgB8RgZ8PO5ffubGENWh4xvx
thAO/txPCpH9FJWgJ94yxyudFW4IP+IuU6K5mQpkU1E+qybD5O+W1HXBzas2XJ+5
tTPKWfkuFvNXN0kdpQVC/YuCVfVGouDoFPm2KA1Fn7j/tlqBSX5MF6mQlQ3ZB7fm
7Xoahn/iZ+jFKFVc1TxCN0rXOitz9OYOxQWhaHMuy3pgOsZcZQkYm1v+rbj8R9/F
ZysW4KoUo6gkjPJFrH5BlqNuItk3Vhwt7xkrftKaqwLMGjvQhCXLsOBWWVpHYJBK
b6IP0vJVMmNzApPu+OWC4NfOEPYHX1wXqWyDt5MK9Glbpqmgp5euD8aXWmeqGm9j
7AT+KuJ/4xYdUYfV6wb5Ao9fJEE0u+TTUScW3t3aARASHmGb9D/lxJmVEoH04eDm
JHIXkDU6yW4S+1uDPUuWxC4nEh3DWnRJu8/nf20MeEqUivNJQMWTuvHiIKHOtqK3
EjH1tDlcngPF4UzscKjbpJosOn0/1jJBwsDQKifIwk23RBYdF3BKofT7aN/Nabpy
fcX+Rg76tZXXq9ZX1zRe2zRU1kKohJ1m5pei3FSwx/q8n5VB/yD1LT1eevhdD2rG
xDoy0ckGClrKcrOUg7oWk7W/Zu87ij87K01FGqBGMm1cL3MNO9+pCNCrrtDNZ2sn
GkpK0G/awhhEhDd9XaC8DrvNDzBMiG+xbd/HsejGF25t0qd+sKGSAmKZsqsIApQI
KhX1rkJEKSJGbPTCZCFEzfsYSjfMWMGEDYPlYmiVz9jh6EesNcPEPQCTOh1YERBu
wPEoFdVplaFYlTCUu1xCXn3UUUm8bmQI3Or6h+PGPxfel8dbb8CKlRKU3E61jdvq
RFgmMy+lqa1RFBLdTazAifpdLZpkjGlIKgPkHWKjNDUXNkjBh+ZCme+/4O8P7OpJ
ALZT82kqUmbtPZ1msiXJ4wdB816KiAFPKbs6I/W7hz7lZF1kIN8xkbFFXdYdaGyZ
lHki1NDFaH8JpE1sTf8w5IZShuBCzQab7bcZs5V4WrDIIp0k7/tibyte9Lioeo7p
TkxdXfW2XPpHm2e3cS1OI18hxOHNRmOz6BlzoqVDlVil8LNhezFaNCWTpLLrj0+S
6tJlbyaysInwd6uGmsw2CaDnE2onf0tdBbqbNdEU2j6VbjPxDnkCMfcyaMXjES9k
1f8zzgCCYC0x2URYMmFQy8p8T+/dFUxwCCaaqaMy69Htr6R66tk34+gQkzytxY6S
QxKi1vtYxv6nfD9KV1jmBwyS1u3xyMapDf0wjVy9A24PWSPF9KcGpdqGrh/fsdEk
RJ/G872AWUUuoYQzZB60MfkKQkYUmg9B57datv9pZht0QhGGN/0LSRVQ0ENBsZCN
DKwQRiGInra/zi7mhGxU7Ui9f1dlVRX0aXzv7nnsPPlpU6oBDhd7XXIte0N75YZP
w9V3pxuvCEmuSVNBhNbLdq9AiYE+2LuP1bHt0EPZle9R6vNd6E0bTQw8BR5c4RDx
vuNq9kYsWZpCPXKZTYS5vItWMtpfJvoQEq9j4+PrzD86D5QUCys9ji1mHHd/pCyF
vYGZYKfQ4XBCBVFZeds0pkGGjDNm890fK6YPomb+OYizH/nczsHbuiDkAIUCBMf6
yyO/ybZZYiZAcOif3g0asG7R6ghbM/BWZL3fkRqFGthw1neS9E9v8fkpbZdcU8EQ
7QGhi/WlsU+aeu1G73zfydmXxjeszNPxd3FCWttFTfSzEfohl5fCWWmt//GJzPvj
vpmvpQaWxZOB8PLvrurrw2TMSF5xJNkxbYhagML7Zwy2iqHplK4UwlLPPSDt0+t3
4mQtOh5J0vDZfJF0EQnkAKr98UphycQW6JjJBfFAranR/wBT1f+q8sawUycvmOLF
YXUiij6SFXzW8nKYhWNWFUmcxSHcy1L+TJYwPEFPf4fJt3teaRXmoA2Ftw09A/D5
rnMLMFOhW2VbQyasE7FqLhq7hakSnI9WNtGh1YfF6xQAWOCOSzLNj1Hj3mKWdTgC
DwYIDkFnEEw9njVF90YBq9zaAPQkKySE/HrliN9aZE2EElJTOgserd+xu9hRRwjk
5gwjGda09wvXP8wclu7tk88vqpxGdH2znuv+llI2jLyqICYXZSINrrgvhUCtWixv
WG20fk3cTUlUz901okrYWZjvCHuiJGxYEQ46RVbrB4GkSWJdbU95xN1p9owTtLfK
zgwWm5XP9i14Es/pdX6uj+V0AfWv4Ym86qBNOSAizSM4W7ju9ze/N6IRP/kL8H+y
NURpaIDlQtMrbKz5gNTaP44NOg2ptcTnmUqvuNKCt37vUcUjb2di/HOdK7VXJAoB
KmIQreRcTQgxZ3vlTBu752kUxgfOKHVhgODi1BiB+Fea8dCElaFG/DNp0wNeazDA
7DZgSHzspz2wAWFxEYQYxr72aM6EDt9KAZZscbH+hfGqgfZC1eq9yBuFHr0G5JzM
p/0pL4V87GZ4I4pzFqzw7ielo4uN9wHAAbJr5309eTNZ7fmFrLpwEaWUGLPW6+Lh
tSgSvsmo+UVC8PV88aCcBi5Odbty3ZC2V57Y7dYQ5QZ8/Yd2QVa8bket2tusH87S
eu5AwErO+GJejCmsQdzfN3u2pSdB7MTgn8D0boKKU0YLlabLyGNhAZbnHavLA42c
PZfhiE/tjRNswzsZHIkj7scnWXFaX7slvmWYMZkKhoRvX5v1fPJv52esOhyLtIxf
vTJdSTQ4A6Pc88layWnDrNyZEXBJHOvx9zKRIanDCPf37ybqPqrk8UwGa8rPovjj
4QpUtFa0/7WY6rgSsTkhozV4ByXe1sftCGjVaRWvU135LN69CYA6aHAh1DEWMHC1
xoYZdH2S0Kfu7p1xWspo/HnkhalOgAQQ3GneXTB02w+xrtUuPYkwsYL/CO+tTO84
tcdQ7vd349JUdk3jDG7hdlLGRj6qih5mPAxJv3DwYRRG27gjHNzgIaQxusETRmuT
iylcDFPJpL7y4KWTcvjCjb8e5x1nkt3mVKunj/2YlfDh0Xt8jJyLVzwU0T5yuib3
vOF7xNW0uydZjTn03z5JoecqP4/MoxFHthG73a7uQEY8DjDPWjyeV1tJkqaUYKqP
sYFsEATrGhflQhx+YDIl1Ub9ixBEokjR7JkgnB7Af8boB/7ecwzqVGIZQMbGlP6X
ARofR3Baz9qqZaOxxpUrzZv1ytr8wEkH6sqLqp5HBsWI3CKiLQ3lKqERgWAA/aWG
Ag5sc5ukdY+F9YMvfpNFDJuSpCv8QUwH93okSI7wRQkFpeViQtD46BZPvA0EJrmR
sVrcRXdeZ2rThZ6BWVek+/5HBZSFANsWwh46Jnyo+qlNalpMCDf8JjClz15jbsVP
+ibN6EsGxSKsXqafHV33Tnr68uJhS+HLogcfARsg/nSuTrJ2AevE+WU+KChjiWja
+SlIwh2S1292NHIjXyiKj8jXK38E1+nZLMjRqnFIYKO6uDrQejUp0pGpE6wxstOm
5axBndAr697tvSO/n/UrW5aT9IUOsl7Dgo0PfObqvwCd409rhv0zqSkBvKPjRhR4
1lTj6Idh555dGxqu8BeVdSqizXXsqS4ziCdmCoxqse08sUt87ngn7Pp0lQv/n1Ye
EMskNtXBTb3UHMXD6mAX4ElKSa61Gse9Bu5sHXfYnI2OygXka2pvGAVheiee+HBq
ADNE87+ufg2/aCEs8rWs9s3w/1fuhGcTIqySeKcRe5SOKAw/fOxHH0nS9GZIbWvM
Rit/11i8gFm/Eyg4XoLp19Gc1SlddOQMoMk7VhLSsvZf570tVTemP3/soRakTuch
37eVJXHJiuhUss5vkMk0q7UHehmlAZjSkSEFoASPpoRhKeKDPZ+Yh/JXImuhKkIw
8YTOtHBKP83XkzNXnqjUXUuT0H/WPTJnLQjj7itAYtU0NakmYAOotxyl36IV40aV
dXtW8vKeTDjP2tE1Zx3vWBZIjWEvXg09LQAC2LWosTFEmhSwV4mIJglzNno2uVO/
HU+ejaT5dIitWmOW94UpIrR63mguy0jN0KNGIzprGdDYuoITPrxI20aSuhzfAL74
XIZXCY2/mqLXsLKYWo//U8M1qhy7euPa5eGXY7UYPpRUgYSPbVO50K/dl+lB1v4L
oyCezF3I6CGL/fiwPk9qnots/YEwDRTUa9zc9UskMFX4gIGjQsFnchF0JEqylL4F
O4tRneeqoquJorxtCV5XGRz1ctXo5nJwbRd/uhGif+mS2tQRnmKzgOuv4a9dpQXP
yeCiHTbTgYdv2JpshA0Dcl6wtVI5ioRLJqIZ6xXMFtpbpYlhezoSfMmcfTQOJSs8
SFYHdYoPsqF0roaooGTfeVPnhFI6IZgn6YZRoF9GneYfL2EDu/awa/gsA6ygf1m3
3cMmumIWa4l4F0wR43lar8hB2Puuho/BBjE4AhFHpmTFMAbBMHOEZgtq7p7UwemV
BKHmdzUDf9HTG7xAmIF2ww549Javab5Npxbno4dMYQ7Mwr+h3QlyfXde291x2sYV
dbq89aE9EcufDT56F34o6ObN0my4gnxoACNYaQqOA+7hw5jol40dKLaIbg0vdOeD
kwtrYUcNAWIXo4T3ZnwxA7srsPTySgjlyH+424gxmR1MfeUdmGsbdCKjgVi0++GK
zYa7oUwj8rRQVKiUZI5B+QzsuEmIQj+SJPlsaVVi7m1rCwqiaHnWXVr0s4fWVf/U
0LLPwsvJAO2yk4oxtoBUh7+lBD4kIGZzFgqcXCB3ExbkDeHtPkILyaUwFkEBDtgW
LgEQeZ8ZRhfwFQqA/UhUY8zknTrfaSiMNqcx1LaRSdO80CpgEHagqf+pR2BoIBnp
i6MacS6qwPpVWwQ3oRbqDWLg3khO4b1d1faNvkZTyzMf0CZH3M+PY6XFu6nDTldd
0VLMoot5K8nezGYeToLbtxMnLSjC/k2ERT+5eNTnh60ZASw4Zjahu3aUBsii7txV
4pHLRoxr75/F83r4lHm0MkT4Np5JodmEGWcY/vqqCq8IiH6/2ifo57k5PWtJQZur
eAEVO/4mnO6j7Baz8zaXSXPIKEX0p6PUygR0zUQfBLI6j+daTSPkuR7MbSZDk1H2
s6rJaIqOpEa1/9g+GdyBPWPzu/0NeF8sn+Dg09c9ScLaewdWHfUXMywrrjnuHklo
xGfn8Lo9TvR7RXMUb/PUiEGzhLkEQo9NLS236TsPS5fEs5aEp5RMiv+CGu5YSA8w
xBbRX9VR2DkTpFp8DZQDqFhFWw2yzlDRfQVLsiIu8ItgTh/Xa6R8Nox/LhDCrYqh
UT5/h3EKowpWuucv+sM+4Zh1rvQq7pCJYOxNG6NMq2i2hNbPkvspbwHN5BLyOHsL
4a92DUP7b/xXlFoX5cowtWUl/gESM/p0h7MgXeQVY+Uv+fVLTkBqmBTdia7WiePZ
sl8GMqRFNyIpSiLUlEGGtATS8K1ZH3CmQ9Q+k0bzcA03rVIxrL54ILT9qCpyoJb9
0+KHGbGD7frU19TukMsDBXuODXsDiXh6nL1j5YDTvGeW3jRlvdBeNeJM/BkZszKm
t/P9I0usv3dHiWbTqYKdjPYLf55n3W/Ly7VhvAHJ+1FtgcUjG37CxErbjd9qECyY
Y4WiWfgLTmAva0rsMb3ph7sRIGzcZqfc6PHFRrIwcdw18ItD0pR3v6vGeXxlo8e9
555CH3P+C2Wi+fI0viqd3yFRoBJN6WHL+m0qCenmy5yBEdYBz7D9nPqmYVuRj2bL
BqXNdr1VptgLJ1xpdCRpHr2raTuMJpHys0UD1HyprfSXdqhPAEavkT65wPH2h4L3
aevTvoW4LyLdb7FgNks3nTa2k1Z02QvVZWQOi0EyxpizkpiB2FBWsa5AxWCv/s/m
UPzdj0M4OB3GmG0gHY92+tAYTPhB/PW/cLCvCCbcvPXw1gkvsj5o/PvayrWd8VkC
BMuPhpxXi1lgf3+QQKIIa3HMeudG7qKAIF4H+1sID7JlYhSzt2LePkWr4L11vvnm
0M4dtZ1T7GTJCSeSR8e+SLy1ypDl6VvHaqSiwi/Yc25xYZ7Ws4BMaZ2oa3KGFmbd
zJp6EQ+I8YUJWMGN7UuD3qgyRhA5KXoZbz6HRU8WnZ5pGpOnyfJBugaKOoMyVicK
A4bOudFHIXA6UZGkf+EMthgAGCHcdUr7s7kE5Y5giOAs7AJR3xoKuM8m14/OhP+k
HlgMfetOzdt9kP23pVO60cJXCUDxmXi5yoznP8/8ToEDER/RgTkAtVUPMB3+Ybmi
CqgQ6DrqCCy4+cfFtBvFwM2R3rl6DvTEqeNt+jg+3tpsUsiK5UKXH0zCAzCrJ19k
gQ/QVdKOdvvuAAPrQF/GgNYsJtuCAhxJsJDIZltybWvKkid96nShlunBwkLYadN6
orm4gtYKsCWMfZEZeoy1Skhf1X0C6TASy4wN3KXKyYJdz4RH5iMLknukc2BasciE
1UqSDhFw6pzqoGfqeW9+6REtiFCCFG+hsSZvOgvMXLFXcdNpalGwllJEUUVPpzP1
7uB8GPd/S3NkYQYeRve4JHRfVClX0V+qe4kdqIy6r1VnF7bv2K2PIRG83cYlPFtg
nC2tPh5Bg8pxfjFFe2Do9/WUzb+9Q+JJ5HZ+iqIx2ha2yTwtica5jmNtgq0A7vUG
Z87N8wNYn4VEvNdLj8rOZiK4NOI+TlFgMqst/O+weS/Y8uNycG+x5CN7jZOe/dpa
Us+mkhAepM5rrckyR6uOaaKwT9NOMFKd5kY9Ye7ej8rqf2/SpQtHnKGLojDXU/GG
UDI55eSE4oVUysOftR+SGJjthasIrr73zcGeTpOkVYbn0NzGRAeS5t693VLqO+LI
PgvXyIGvelWVhuKmnKdoVP7T0Mv/PWrnm+pR5diXCH98uOZMSHtnbQBbL1QggUlz
w5+tnr3dLppVOMfPAafq20wHy5SeQxETAAlNNMpfc8CvqfN/yqWRBPespxIo0ENd
yW7kK6xMF26cHRSoPV2JTskPYCGrs6d0wgi50Fb5C3IguBXsDEH692+Tiyy0U0ib
ZIKuiNQi5+JLtZ2dR7KplX0HNYL6RXh3fJfz3/cGeS9XOgRiry1wlawQtFR2XJ1Z
0g8kiuhUBAnDe4JP352SMj5b3qbnwAR4JSvZsOFqITXrUhPiqbclxDcMApFvfqYG
yf3kS8eQphJatPYxvdm/8pEWkBnZYw4Aw+7Xorp23d7957L3RRuD5DaJs4d0ip/m
69UTC7gvzKt8GIs1c977xszrnspNxxvpsrKVpLQsbxXPg+r+OpA558cE87UJVAc6
ICQIlou+WJalBEYVcYZfxx9SjZHLp6SeSm9TG8Q69tlzJkmu2DvNidgwgt7/4vWR
zDmP/U6Qi5ki7N86xZpveZ+NaytkwJ2KY8R36ySyWqUvCBRl2ai1YBAiafknz0dR
DuKpYy/5zgnT4R2sbCUCTlMmvZ7XJAfDSdiaZ3Uj4k8tHQGhNvapgRxN0U1v3V+F
80axASMzeodAW6zcd5xGhBAlcr5lMayknWYjECAzH0oeKeQOrY2yavgs+r6N3tRq
xYjokLfDpbAUVOcjoyaD91JR1qvJkRoLXLqIUqGb2VEttsPDMsCzUTcbLbvMq/OV
iNof0cSQEdqX5iEqu0Jfsubym0G/FJWqdvWpH5pKpzshFC4NI+b+6L8NrsqzKERU
Zl4kMQexYDjg8F5+bEWajnr5ORH6xPZbnGhT7wOJFKl/F98C5zZ2khspm9J7+qTN
nkK+oQCLLUrnTUiZgMF5kWgPCeQhm8y+GP6hVFK5eiV9zVgxR/kPwIgmfS+1pPqZ
//xBvUiRjNiYSJZlT4U6sVJEl3q0zRlt+G4Y++yjvQ3aOoHDzU8mEIrlj/ATySj3
x68eybBmjmymym0Oa8VEScLJr5CwubJpDI80+YGQU9qoPGe4fqghErsfm7bDnMpY
YwIj2GcVvqracYprQSOCQ0kreOYEoSGT6lND0JnvtWlwGxuYNpzfk/tngUn9PYdl
Jm4Y+jDHQCXxBJMsd3dn+ayeQOMvybFPXMqIZWPn62+Fw/wFX/e4eZpLi5Lrh7Ov
uc3XokasqOS1ocJ3FZA2ccYv3eXdtQIOP6EyYMR3eYKDKdaKhUdrO29FhPh/4w75
FWT8pIQXE9QeRID4XNX0vX8pb/xCBRbK4MJ7hGCs+f6z78/t0F63HAR/3uXFkdV9
mFBhPUyfcz6Ua3/DjaxbjpMvXM6x5Uu1k5ydE36nwC73uNgRQZsWPfsoxhMZMZiT
nfpAK4kyewkUgYOdZUuPWD+WZ7e3+6UmZo8NmiM4e4jbMjWAJZavfSe08PlrWagT
GlOM/u579vUb7Lf0PT263rpGmVAjXC0AJVUXGXunWHt4LRktcRXqLfWGp8DJVPwk
TJjcPlqMUyOH5H0YC4W+dPeXcW31v09V3oOXHi1PSXh3gUVcxsEtJ0T6d1ITITCU
eZqS0xMNbOPGtkQqtCDt5QH+8TUSSDeVLR6XaHYszjtuEFn3WemHe4N/iPA8Y90G
vN8wY2XjrX+r5AzUBJK+VHTEc4H+bCyhK4EGSbr32QeXIMo59yHk54Q8IMVkoK6P
17A+XFrcoZzwDJdcWh+f7crizBctSPW960DwAz6qECGiZvt6V6nXo0Y/fAglCk34
kJ/IAOK0l/g7ZVSjfVvMvztO57Z7GTztPUYiPAgqjDwQ+Kx3ip7KCRRuEzTz6Zaf
7vu9dCchDADNg9IKBQIbnTGuVH7NiR3hhsbUWRkYTrAsYqYuX8kejDVCPWxyvaza
zuPbcx3rFT9LAz/R/Kj6eXlRfg0zmlM8uJ8QPEwT5otRzBVnXVX3I/EMxnAvB+33
zAl6IV9jZklOrpSvcrXhVudW9QoUe1djzw/cRbwdUcj3NLvXA7Iv4wH49pzCbjlY
xfBJFe5/TQiXF8rQ9/cM1Na2GEWTUckj+Hu12nany2mTwU3YSIaCYM5FIWM4zdPV
ildZ4VdR0W1fYh6Q86/5z0uI/ZaErKgew6+dzdwUZn1GFdQiDK6x5/HWIufqhVQk
3CQBNCQRca8mLauIuzSA6+oHFBJJddiZviXArZgsfo4ndsc/hTo7r9oz6tmGRCph
aPV9fkWjgsKhzX0kb7nsx2IInkWJyW8l06LtKjy9UXiuHuUn5DvtuxjuIYr9Jgl/
OrBioEUwzqvOGgj5CY0LveLyhCKA5qfw58kkSxRMEh++sMWmyBquA8m67o8zOWGH
RoPcnKVGzYVl03HWwaUNWKeJvBDH6pxAadvmIyedHsh4Ozhbk6mzkp8ydFKOMne7
2Ujnn3h1yeykZ0Xr+2S9/XerS/AEu/OsdFVHJ40rU8Tlmnj6pdz8MoF5NobuCKJK
C97z0yXuUXqj5FWI6FhTQqsz7cQR5ogv3eLf9TmNsdRH/57gM2OkNcuo1mNSgTfh
pokmzv7N8QshbPo5Mn5rY18SCKI5Hj5WyZweo98WnjV5KiiLrb7zorRzhcubNPL2
zcSKPMfwOK4+oZWZKKix9HAqoA+JD4k5M9+ugLZ4dxp7Nmw1bd2jALwK8xmoJtjk
Bdkj44Pp671+LJWfhSynH2KdL+3XH9bELTJwI1RhUPbJvp/oAqR/6VCGmb0fh0Cg
rT00L4vY+/Lt/e7it5siTxeIsdLJiSZsiejyMNNY6zwys4JAk7JGkwAaV9sElXDo
3uRrkZAZBSWaFleGs10hqTFogymt1d+N2K3kfhVr8UrU9bszSmFNOEWZvC+Pn/0S
7/4oU0N36u9TjF6b53RSB/vd0KrvG+WdkPov1+ycKSZgkR5tDN/vD0o0AYalck80
D08TKMTKYcjxoK6zpMxYvAWf3azoAlfigXL9uRhOI80XLV/MPqwqxXpEUIbNBRN5
X+FBC3z6F7ObMNrfaYGu4Inh7kWHS3QKoUivTc8PL++klpGHkYFMwugp2OZVt6K5
3xHAwB9d5F3N9inN1cg8bb4oziyqAkg+zsGNac5ViqMG7WP461LiP/RmDQCgb483
fZ4HzFAeWW93j/rYfZdBLswUXvMaWWgMaN+Y1Uu6lofdhylzbhLFiIlz6BkFG9ar
lxImMUcWSm3X3gtQF0TYvXnChSDMCiPnh7LoFXGH7fexObM7siZ1SnGA3i5Cac71
EUzAu/bo5Wvkcdcb67NmgA0ayaLNvMMhbw9c2pLWQ23gP0A/DYrJ5nqqvzb2U2Qw
6Rt7eIdksUVTCeVz35FY86E/HqcJnaE9D/e6lj+ec8ROYUkWdsAUoyzcjCRdeyAE
peR+qLYjVbUGo+cG3fZ8y8pfrnXPd6inpubqcXrwl4ZKpWHrGmL8/OUN33fgRnRx
+A+L5S3xrsUvR94S7YOisAxydQAU9pF5Y9O6eJ4kP1sdZmQR3xx6nssmD2t5tSNz
C45EcEtRVSDKAUfR9MJBBXsabz/kQ4F8HW4XqHbGU4jjEclUjIHwC3WrRBfGF+VM
lwGEU8RIOMb5xWNUCfy9yNY2vlOCJiIulbz8IpvsRQkVCO/iAR8+jj2jApSeKSSP
d5pVfushOof//VVETDluFOpzRer/lijtj0MzocjDMcB6KEVzkZJCoAyWh9QOzfJo
Pa01ZvD3xtNnm0p/7rnsrQc+KE3kaNmkVbeH36FcCym3WbrYcHl5f7cprbRXg9Ot
5MV1lloRuRTB4duT30+AT+OlQJ9j4TL9TWzBrf1KqI11xSWXFdOj452KmhBHyYBu
lpo7BHdeoareSZw4rMvYM2vbTZfIxQUtA2vM0aCrQzPuFK8Pm42WyT2NnAjdPN0F
OAwEMC8Wn4LyyuCVM7ZtkQqlOa3qMe10S50HePxENIffma1m5Lf91+E95FodhzPc
Vjeu9SLLhSrUlFRddAshUFJqa8gxP5LcX8kk1BLZF69XG+VbZSdapcpzJ16OuQhy
cY1icpQ6f6+O7bo/fnB4HJ0Wy5bb9GPlHAt5ZItK/+jcxM4Ynw9mMAWnp3bJxH7a
zEXC2MRpoS8Y1YK0ExNWRQwYFQLPWdegJxcLYimZZflW/quGA1OsgicXD5/lAaGN
EJZJpZ5GPhiy9PwdpnOzWxKJ7F3sxCvsWqHwdyXL+EKlIyJfzfHmia/ulf8wfNvh
m4zb9ReNNP22LvCeDYtf+NhBtFYfXZho8/VYvq8eoMwiJR6ow+KBuQV3p1hfBhDa
qZgXBPlIY7Hu10pTHiYrJ7kDj9SnyrT0CCUxSGSdG8cLAB4b1BugqD+jfvGrT8iT
bqpbWfcyId7JvDPlcBTEEuCLiuovGhWmKN7ZJg8akq4sZKxUYWV31u43AOOhTlxt
Qyw0g422bEgA1VPKPHTvB84yNS+B/GI6bXhLDN5g7ukEnLAAOrAVVLMoI1YFIuri
dsV4swbykSAmpo9161A7WJ4RyR6hvIOD0oABLLLhClBi7FRMLbYW4Ra6IR/1xYfP
5l4dFcAPi9srrDTZMt7a1iZZ6Db/CK7UxVqyBEdzoG8o7XlVBG88HrmUqoQCKw/J
NCcuJbokmbsJBQg0Hu1OGLcTipMs+udtc4WcopzWRyld250D6ksgSaCRbVri5kGA
uhf7g3fFg/NnzMbBYz+/674DG1ck8yySwdMWUPZ02tctjZmF83AjnNYCtwIxIxNt
S+n19xG07sW18i/GgXI7cxE1R5xkDRzAQS0j386LMaL5ymgN3ArYuc887lGklEnz
TtXY65/TtcWuAAjRWd8rurugiWGPbvJyI+aoWPdfaKNUblt7JUh2uJNBb7d6jqlj
aHajvuxUwpz70U9ANwIbv9wYDS2JRc7hQ85m69RFl5s7SNb0zUCftWYeSBxbIluS
3agSYARO3J+qd6zi9QczGhDSYpnu6mw5HDcG6fptKZ8d/NAHuRwu1NvlXNl16htA
JVqFFHEW0rmD9RA/EYSba5wkhnO1vslAjMXjWVHdznPfbb2dxSKHcXAoM0UkNVQD
VNK8hkipRkFc4IcqH+hVqdqtjFrlDqbCcAD1dvE1tpgPQ1lVfZ+GItpV3BZLvOtx
75PtoxV39gxwFUix0GVReliTA/UnxmLqGC6ICWWzRdGvZhxjfRL15iruBfG409kn
9/dByxpbWi9zCyfJqTRxrSvItFUjuaT+YEXQXmsGCbg2scmtsYTxdg3D4oVMSG8n
gCoXc45mI+EcW2Se0LqI0vkpCO47LM87YkZT+eETWT50XbJOtfq9haO1nsD148eH
TJ6K/oqZ8WX6pw+qtAnrd+C1tIGypF7V4ta89B/tOrd/Sv0+ZJKg0vgUIaZTEUmf
L/j5P9GnrVYGAk5peA5x4bgKG4ON2eFlXGBzPdxbBOjaXt0qhtZYvKot3I9oSOGg
C8i3ENRZ7lOswT7jVkYjSyNslzF4vfd1uka6wxknUrFrq5KSGvoiY2U6MkOcE+8w
ZZwcR2KKejVlCoyBaE/a0bL3WRIADsaoP+DLY+/888YHn66k8ENafviTXg/+2r2K
CXPoogqeVUMUneuxPiXPbVR7nitTdUmZpbWaHq95jf6T/UFX7Lldzeth54bcCFOX
2DRV2f+eztdH7QU5nXh/hIT/mdZYN35tSghCcl6fescvZpqW2f2/y47faYShsa0d
C9f9+oxuCXdnxCMH2u4BEjCkkynyQm6TNEL6t3YPysVM7HiFvRf3oiNBGkyoYilt
MBfY997ANaMCLJLKqOok/yiYdCEguYm47t9l1CzILE8EYmUa5yR7AyCIDeeBEjN0
fPuAFMy1n2K3HWZ+v6NDHVOllems5pzaSzDmJc5JPXd5b5upsslogtFFuZDiEtEv
SvSlTwphTMhDE7f7sLqzlAvS0H7KKASHrMA+9CmzI6H6SZL+9soqbxsPK6+sG+TP
TUtS+1XzI7WllIcn9MhBPNvpl9k9f3NWkReyzfjsb42AAerCLlf8yFqNvCkbKarb
Y9BjFiglK7Aihtew6EB+QeBcdQHnVwByFcj251GZaeaVcrfhYxBhZYLepYcWwmFV
RDSzn/f8XpNCW5ItKbT87fDxojLoVaG1yR2QrbMwGO9RYdsLjbAwzt7zsFU9nDWk
X0m+k3LYmt9AimaC+WEWL60xq2AfVYRVk1FpZTRRC2NkQ9ALpyaPKH+lQHQTczpi
fe+hot749e4jQOj+16BgnT/ROmnntb/qNQl5J2jli4Acg7OEooy43eZhCEfUCL7q
f6lziFV0tY5RbY7cEYxaFKa2d0HnYsrkpptFCdCDyc+o/SOeGogaEScwkcWEstar
VqG36ud6tOOF5NAUHuy0nCpTHyxTJ0TxI0PLIE5qCNJRgbpKoDOo1yB0YRZQSrIF
Gt4U9yDtYYtyWIjrzt/yNj5GMBBR/bBKCh6S0vFEQ01gQpjEEnOL5ReGf7eWMM3L
nbKkjmYj50uSr7J2juIIOhhm2F1ccSZgAX7bK05pu0vwfwo/FX1mnybsb42OXPFD
fTQCTiYaCZsQ4osIUDa8kqOPNu34gqei/Cmo1jwPh6Moy753Mlwmt9Ooz3i0EkW/
yQrXpw0xnt7NzWDQxHo4UgR8Q9waa5BBX/VZFBVFK/JsDlCKnPRaBsTsjO8rFyad
q91d10YXJPZt/PNlrTVCzG5vFszP0O4DuxVoM2qlVARY2EuNJr9gTIWr7dau80Bl
ZT0rlivnMNSanfDjc6USqWHkFq+sOCwlHN4iAQYmQn1G/z4riaxkCWcfJRZ6/91C
CzMqq/jZPT4aGANfdZeGzpzJQ7T/djbJrd61lY1SdwevIvAaog6chWrRyVw/4TGi
QMnoNKuGb+bhnDuFxUk+wQGPKjsBprPuqH4jzOjvg1dmBnu5r4nIiT8SKZc8cFOu
Nle/VNfFDU3VkQwzd/7V7nTQg7WWX8g2f9QYsRM8poRgpfaxkHBZvmy3uTrvGU0V
q0VZsRNjRik9eBnPSnm92UDesfbHvftsY8Ef6E/Cked+vljBWQ4OxfyI7phmh2QT
s9gMKIph20GSJ+JE8HIU6vVvpXJAY7XatOrC3hv7EvxQSWvfpu0I+rnS7wtBg8tL
alMCMOFEn6YgfGHMhtKDkJzdecLD0Y0w3XMC+PJ6UXLJx35E7suYSGi7nN54mRkT
hcKtZPxipw222DWqr3B7JFWHRrfB4YYhmosVWP/toqmk0EFPE715N+lrC7OJpwm/
NZ8dedXeKhUJF4bhdpZNEDxvFNnCYxMRpNslFS36Agg4TKA2x+tjWRJK75tK0Ltu
kQebIBPY2DKkrK27ym1aRwdLKh/EWSw2LpCDx2eLB8WhEY5W/Q8oOBoBjZ8m+faz
vbiEPxl4KOlkLP22lffqe3bSh0peR4J1gO4p9hiDrxbZFzgaHfJ75uab2wzePVtr
p1/x/+RfOpX+9DsxQaZrbcZpfI5akheBE+14IC/St6sd5ary/UMOdvcPPAgU98+U
DQ8O7ZKmz4VXc/zpTP6m4l8yqamRi3dmuWDewv2ag0mrgqYmxbQB8+Vgbmp1SJcy
QykiWOnDElkESkbXxPZ7VHr+7Jf0gVrDOHTuzVw1uRz8pQ3uaWy40O3xA3oL/lST
ECBmW1Iic99dzxXTTtluOktgGj8ivsGnwhEpwfB3pfUqir/4iLYg0LfIDyBh3jh7
dNnjfmR8ejVk68PXQSz+u+7cJ7eGp/I//ZmIGkA6P9DA885usmEwXesNDnR9/zVo
cA5bxAv57E8u/AKbAgi64ByfNKKcskYmN+ZoTU6fARQSbNBiJGo51NTBZoA7tJPk
zvBTrYJ8MyEau5QAqw1Dg6C0nsY2LSLHAbDN7rDYvwm9Zx386g+2rcViXOmMJkzX
w8L2R+zlbBxcoPoImnV5PP4BEbY/uUiRA2m4RNdAAz2Y+BfplwMlUFbcWhE+emZh
8Go2H4tWyri3pBGTeudbKEyfHVEJYgKdX6hGRsuzqfVOZraeon7LhWxQFQ+Jm/bg
2rQrcr0IRyo0I01qEpHI2SYEmeMbcXRT5ZMl5qDzQv2hBaE1IRySg2VCLE5fw9SO
/XZZT0vaUdA+syouoP8Y7ZtqOd8zsNutgGd20Xv7Z5qpiBf7aHqxbosn2mec1UkB
lKN/MdW1QJ5Gb1yhH8IaLLxWRaQGZaBes82NgHRRwBSBvhhvhP7Cr2vBFufUy0a2
HJ9tuSf896av42MWgVtl3YtPdA3JXxZBEpsbyK4CzCBPazF/IjyPN6rHcq6pQYDQ
m4zrRszvqI/ePJhWv3VszWfDjvCCgUt0S6nvy138EQBcBWquiv9VJmnd+XRsfoDC
H0iUR1YKM1hpgJN8p1SG3cAxqBWEj4ZR9RXZioEIz1E6nl47cjC+3ipceeLaqevX
lYQkVssVn4hRFPYoaF9ubH0+NTa5gkDp2ECCrL0vnPQ9qUUI1Ld+kyU+L1mVPLdi
IPXmlecqgi78yVYy9ILi1JR+g+E0j3/QgV5J148upk0bq3GG8UkqkyuGUe6lBM+z
/jOu2CM8NRoJrSiOzbeiEpvEwxqNnRZm+IrRM9mGVNBjOi6mEZ07F+6IgaBBS+VH
X/dPuSG+9i+f6StQmkQwCKJt/5htuHcjcMwOsb4HVtIfKvqqYIuK82czEJrFTF2W
H5K1AKxHggYrDlROSOqTP3a29CIFAfYMX7MtBt66I8GwuqnVvOy0brYztBctTq4G
5WxETraa4kvaDCTt1U2rxQcUblNzkRw03Ot0b2ihQ6jd+alNXkalWYA9oFUAJSk+
Ckrba9t/6B+EKbQE4QnQsWClL955jsvPbrkclhZ4IpuM0HukonZYHvG8/tQYryPl
nD1tDv8Ol/GVcpe+6eeIFptSxXMvAF6V8Y0W3mSqmsg2+HBw2dNm1Vis3jznEKYn
OsYah5jijVdxeBbfeE7FVQxczvMjYjZ/nzz9bF7Uj25ovSW4svdkUuroheR2Hn3y
zSEjGXlX0pz+LFLLB4qycDgbFc78jMoA8/VPTmkmAbXwYqpHgtupgzB3/JuD9wi3
NHv9Gro4Sr6KeCjl5QHP4mZ9aNvirA1lPDlE0C5aAZEhs7X+dgXZoWJ/QPWJEaw6
trKiYzfKUyRTyIEjUgYnxn33Lp9TdSmWMRbu9jACbjgzQ8sETYjs0tYZH4ui74/G
YQaehqfAmFBP17bAx8uWkOrba0gljrcotFP+Tn4zOCwVTmt5mlgIVHSer9VJojj7
f0Gz7AEWiIT7qimfA2VGYeLUQH/wHadp2bE4hYz/NO8fCcm7Apdy4AFfbV9Smqhz
nFCcK7LPz7afr9HxBMUOHGZ7vY+gN2b4PKbqQb+V4vZ7gk0vIX/EFkIQDuMW15Ze
XnM1DS/cBdSSrrDjrz47UsDoAy8nkA7mGr9Va0B1RAAJx1U7TB5Z+U0eQn6Tl2lu
OEfPiRPgWhgoChCI4Rcl3M/c3TdO0mnCZBgPYAhCz5oop25fIVmL27uwUKCSHcZX
kKZ77tOD/4rs+gS5dOOAeSkBw70yaUHl+j6OouIoNSAESScfeM0pk58UwtN3JqiE
7Fz6t+7uN+bFkClcBIyndilAlDfo4yXCc8Jylil88uk7kA9hsVzg86cuVzkzQJJ1
BLTSHo1ilRU+Z4b+J6LHshlsBdBf06yEnKbVxlR9gksxIfH/V4qoaaMdBcfZMbhr
45shxXsvDF8Mbx4pZzW+NkT7uK/nGT8DioDo2qK4yi+1RrnJHlB/SsDNwqX1hTT3
SIK4UmpiAKV4xAoQ+fj3dGjXqzs+JR6jpQgqBu5zkDwpmsXW40JhO9et+cCeYkr2
NxKcOPSSgkdGR54LroHZN6lQkOYJkcpPNPemQgD9U6p7015sTWX//rky35u2wV/t
LT13fM7TDz2EfBQk44o0bVIliTgaIOjnWu6D9Neuo13dmUSip9mEVihAzb5Vf1cR
HSsFVEGN6ssOO/v1HEGK+fZcwUo3JndNtZZMjzVQs+fh7Pt5a3OUkq7/odiBI+Mq
yCeO10u9sM83nShKKVdX/zvGfmtQ6Jq6l48fGNuY5bdFAS57KlJ/wlOHXAh7Nhuh
bO86l6Eik//8Cj4yanhSCs+5l6p/PJRxF4PRlWaMNCCNCJPTVVexreXB3oCiFXEw
7sAinvhegp3fuLrL4Al1HTIouAjkThcwO3fFt6c+MCW3hKNv6c3qWZVc1gOVGMxD
rHizB4cBYTwjW+u9A7bW2yCr1Hbt8Br7ALP8L3jsiTEtJC15yuCtJfKcNNiWx0MA
PuhF6L8silXffMxa6ItPyrL3sPGN8EH82wfTQjTgnE4VlD+SzD6LY9LDvmEYrlRr
b6BhtGuKiF/3My/2mn0GGoBtIjStIp70MINN/ylX2vXcIzJn7icNfJ5PK2n4C0K7
q72ZjQanSRW0P+Ki4DuWG1nIUC5Z5bWfpfLqf3HmnZ7h1ay9i89mpy+1rQ6hgnO/
c81grdEI1NNojxf4jgexbSG30YqA8Ewt3rJ9zLbAT96gC8GjAs7ObP/G1Yv+vupR
pN0w6rkSFE120AF4YXF3CtlwSuuTobQXqtvR9wZ2y3hRq2s8IJ3Powhkb5tEiPTt
qNdt34FKcyinKZrNNj4CfK1vJuJHJ/+G20fo6GNJ3mTszPm5+FKplSYdvkQjvXze
HyQaRuZZXcoBIkhlLrwCmOmN83zKx4D3PVFU6U0ecp2Ek/KD6CD9s3QTsI7roCeL
pZuGi8qyljk9Jnf1uubG3+LCU27z/FCXAkKZwh62i/LN78Pa5xcDFUz4MSyJjZcE
caqCcJ/UZxXX7k02JHJBcmg6SJ2YA979gwcb9k0MtfK2HhO1AjO9Kc6OBVi1hZjM
3z9Q14oU8X9DRnQkHnG0hY3dVaNWcQqmGFKIe+0B0hQi3z+dFVpUzSwfEn9IvOvE
ivtv8anuRrqKk2O4rOQG/hWeTATa13trTFIYc6QD8cjeP3wnQfn51lMZIS37zKO7
S9HTvOixOSLAgD4q1YCjG0fNhkHKeSUmFzSFGaJhDxj6CsTvkGAXbzeLFWT2nRcR
06rJ2386q/WUOKLoSjQE5hTH8DPYpP/hzc7CIawUjnSSvakMfl/2NmOUH9W5E6mE
`protect END_PROTECTED
