`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rm57qh/jAf+9vWRP6+nr1UntgcC8NNdCSZUU3F6lzLOoIopjSCsujTqvdkmf8Lh6
EY1GhoPAepW5nhfiuBHx35K8ekIiD/fNWJizjerjwIsmuwkyxl2AlRbXsw1OjiMA
mRI7fCmeHZ2MXFPmHBtlJTVNy9vtEjK8ymCwZ6dHEuq/pvTH3SZ9UJNunnfZmBhw
N1JX6s8SXT3kDKq2d1aqj6P0Ff6oZz8n14mTwdICfdQIe6VJtzagFsiVj4Du0CnB
5m7eVkpAw14+1b2/irheQ2rxuW7w0/jiUDn1O7oUPoSTk5hMmKvTRYVzcHmnVmHv
AcAtW0CXgLwozUg/UlEIlfBksZaRSbXaM5DAH2Y2un9VDG8BjgVWicNiRM0w4ftS
UxOmQvjrPpLuV+3mq06KqDXwLlGAt7MJlo83mB+LB38eECvNygmdX8+40jUuX4AB
kB822Y+5s2q0ILL1+vNzX1IVl5wKm2oVV5rVkwmVF2VKOJ936oQcaD4ccMAxGpKN
Y6AdeL8WOT2pdxOCCemPDWhc+IEUW4ECWtmqZaHrDHL5fEReQG8vXd0QATVomRVk
J1pxtr9SBOaZ7CGceGS/Lo6bO+1RuV2ZZLS6cKmCppZKdLHQeQFwT77f2aWd8/6q
2CEkIecJ0y1mN3dAYGeye/3Lnn+r8ENkokJrB5rjDLum2wOKWs3M5K82CbTzLXJv
3H3Ma/S+LVwqbSK6qcc9pISpZ2FaxRRGvvAvfm/mEw5oMm1R/9k9aJ4pjz1OOxRf
RpPrCN65zZJiEBwzrLYwfNpGTWpuZLd5zkyL187qmsV1wsKrHY04/PNtcKuR5xwh
Kkhh64gmtC1LvqPolQlBB7bVQ6ohoJYLJGOSO29wrPDVSc1kWCKGZgLI9yX7s1/p
ozPty+O5stLyd2Pksqv2P4QDgf0G4OoF0UrP/oiHDFyJECseiIMYyrt6LIf9aNfY
mrghd5SJK8ADtLvza/3rmT4ww+3PVuX7B4fOubxLpzPYdlfZh0Qw5dx67PgwpZrO
W6k/BXvNSvUOHyj5hl94LpFtqlwV3bCeJB3lR8Om1MfBvBL63LWjfY/CN7gmfv7j
xp4qdazuF5G9DuEmCK/4AXncqavqOmVXTejSkBhZ7TqhNt9GQ6f9BPJMgEPWTOsv
og3OymYdwL8/x3+Ec1zpm1Rdw7/MC4SZocMLpbwy6/uTHSStSCNqa2YMuEgYc2VO
KpuZtqbP28kuS8XV/0WoD7lMN/SJaeGcLPPZrxDsZMebS0lrCus7Rf8/VK8Sw8Zv
Y5rO6y4qPSXtPKg9vjlG/m5voHll4AKx9LYpdd43zGIYYrHwZIoLmocZXQLYIE8m
VBd19HH6lKQYbhRHQcnWE/MOw817X3VFNCwDxKzWJlBxY8Synx+T7gVU438PVE66
ypXGc9e4uWjrvzPoqMuUAxiIpTmWeItRmKfPLNMBJyozB9uIERFPNj2Gk+jel5Ph
nmz6F+b5TL85vm5pLwLgKCdaVUXS/CMRzEyAQCOEsMKfGvFXjcsm4o+SifwVxI/s
HZwmjMdrRCcL0rvIO9x4fZj91zapbs88V8uywWCo2GxRAt+gqs6oOZ2nNY8jogO3
AGZRAuN+wqJgAcoRAccPExGfQWnYTF0VSCA4X9EJSaAKraj+fcXEGHXibIxkSifS
`protect END_PROTECTED
