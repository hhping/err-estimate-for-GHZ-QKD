`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPo7tdLbXuScq9JuqEseCwaHPQZqAmcDaQCjky2PDKCtnm8Tk+kHRY5FMOjkYx7m
fDRT4m0QpunUGUciLiODSNQey7vgSIaOj4LLhSEu99Yij+GB5vdGJY0I7kWANAGx
hAXzCeC/3GUT44d0ZG6Y1EXUkIxLeRAL8GFqv7SdmWHgTsmXBhV0fxNSo/KAulNj
igPOZKCZ27G8MkgJCCtoaI3B/yzxX22n2MHS9kbJ5ESYcjbVAmnzCWRs5ubHaa9z
y87oWOixD5M2OT4KLi9ihRXc4TOIoTuMbez3SejJxs4kguZBdWPSWJmQP7mSsAKU
zw6GBwuU/nZZRx4FadCIpp8UNlhH4Zcux3kVSQjVjXd/hybVlFoozh2CHH1k49f7
dBa/9Q8YtKf0HJ/8arMtveR2lqOx/44hx53mh2+2irfpRwFIBIolWOmpvooE1HiT
J3SMYNV4PykKNAcFWAJz4Vd+Tz6iWeVHNrAjh1KkkQfNqzsEuVQlaEPVGoYD8hAv
AL2uxFAmW7ift1lz0YXVzsg1xJLpK2jrRSZUMS+mUx0bCSGdLq1Ujc2wbRIStz8w
HrT7yyyS25blvp0V8K4eLqAy9lBbuDLHjucKDVC0y3b4xO2qPc/sYnOPQGWumfzU
rHre7/WtIAQ7gOtM4+Ojgi2sE232O5RkWX8dhPPYKX9tbDIXsdGUi0IwIbAx1Wbr
89JVK8jaVfkoPpXnmgf05g==
`protect END_PROTECTED
