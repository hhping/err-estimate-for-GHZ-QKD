`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLyB2egXe7n+GPBU35TzlfWkfWTKcLKC7mSxnwDgF8WMLNfjczAXYxkGH0XQp4Z5
/8LZ957vHASlzoNi1pd10Vsxzgvl4FOrXRUyqVGeA934SEsIXH6gsqwMyyWcGUC9
g7wkvkR8wDS5u6dboIsEA8nVgpC7MMbzvpdlzxqU8d6cp6PXSxDHTDIV1IlsxWf/
9SSv+FzmV2dlMhDNgJazK8fVyV9Vx2L5VucfMf9fimJbWqDZr0UjXzjWBXt8LqBJ
Ll7kpI8jvtWV2cXG3GuOVz7WdeJqwnF09I/9qcvuQ7JWnGTr2HEFT+XnrBab1Fli
ScehOCsFvDg2Ex9zvUqHLEQciRiMwaEFDex6Wn1dPeH4wrYtTQzCBmN8loyMiUVf
1O+wUD7YmCvjEVDpZC/5X1Bebhx3RibNhPurZXnWVj6ZJbO6VBD48XgR0G4O1bMH
nq1bzt4F3hLxfwgdKyng26lD7Rn4XKyd21HCUBG4rpG9zMaxqhYyRc/Enb2EIvRQ
eh77zEmgvLFw0XvfUOk+3nr0GYfiFbPz0JRsi6u3xp9n/zYT2Q9i8NgS2zGqTgq/
5FcDVloch196i61gr3PA79N3+/+0f/XT9u5CFfIMfwIqy11sGNVgvm1qr2/n0O3G
sDCQWnnuqwHC7LlSjPzqOTPN5SzxoDINgP7Zhj+um3Vne4Tp8YM3GzewdI9nRLyE
0jhiwFrDiqQF/fhEha9+ffrc/iHZyqULY1fi5emPehk1ckE0CjZ6VpxAwV+Ivlym
nLXlp3nrXyRFeNo3LbEBLuAjOhYAdVIE/+pQ6/bZujEEDjq2U6M7O3wIKWI/UgLq
okDBgC4PpRlB+irL8rT+o/QoL68iylIjyYhx0DY01+V1AgQiCniws/Qd1J33vJz0
0d7yrfgc4yLqhdYnFsUPJ795VCdgQKGb6FML1dJrOxlKEZ0At7FrFkf+nsApjxjc
bvZ/0YurAO1LZbtUxWffsB84LIhQpGttRo/kTAyZdWtF/7XMTyUw3JsvoE6+BOHF
+i0qNrR2yGSmhLVJSQsy875d0iWQ3wOqybvD7+KKD2s33PTSBj9gbwgY56TLc4kh
W6gxD2phv425E9uYpCg0m+bI1c5FS04aoHNzNwzkjF6TRPNlJF9Nn1naZZjwZW2b
dzkLikv4RvIq2rEOwKCQCgeIS3zDf/vUQ7QydgwsWZRkWp0Ulxf36/QPG2SVOLQV
VCf17XcRCC99lg1C33fAU3Fqt90jLgC8d53SkK05//xeKnI3WieRTtHxx7r8C2SR
9QUb4jfXyKEkUrDp2OIQTKY5eXQAds2OcL1BOCf9YPTU30WIDD7gTw6u2p7TlfTG
BIgjvIW66hBtcsI1WAmilzVprbL1Ad+qFWOSoNefoUQnR1Olw5zCEXjSaMvDdjAt
gUGTbj/vEKTN+K8lmRVdQWN5CxN8Tl06NSR57TNvpbND1DFPh/ZhehqAI/LwEaM7
5pO4dlF+7HibCbbvlOXorEGIB/8U1BXz4cvBFRxc3w3HUbMQSEf/P7YXP0GseSbi
mZ70KHJ1HoweOJcOJ9XEcRTOX89imb8+6mvZsTvvTe20fq/2Czjp1sWwiAxYsB0Z
Ok/FdF1ncYeJG6iVPv8Yk/g3mqFwZA1QagBshzD7xgbRpAjx9o76hYtuoDwhH0RR
L+dioIJgohcnEzrtkp3+I6zGygwKGNwpTOo+BhetMuhqW8UOuUBJ9bnpr6S5wlwn
ijhKXRQgbVjdyzapnvXHN1YD5jLR4EVLYqmvEQFoTBUHwB4yV8k/TNkjw7JswR8L
BzanMfgnAIg+kxIMLKWl+mbD+3EzZ9Yd8HOh320XU//V8E1LzNV9UTzJGN+Xbn38
Kr7VyxpYENL3x8P0Hy8vtkdYqiG+9St53uOpRi+ptCXnWKZw5FkjXFn8K+ZPDvTB
gAyZwYH4Cxm6ogln7zbrccPqAOx3Q5o5pIqdBD3oHhiSvv1q5DhJwcgo1dLqXfcO
84ERu9ELZKUt6Nvrgr7f3clYjXVnn3Bs3w0mkmfXBhNnPbB+TKCs+PGZOXXSDj9X
0gGea+84rvgT4o6XXkM+2rR95YPo4Qr+6S5zkAHtxgDnwKRelFVrm3AJc78kzI5y
+5aktZ7QbVJ7n+z6Z55AF8sCJ1COzdN03yIDo8Q5+tU/UH5B00wdlu/5l4j4d2P6
1K5MAy7uNq5ng1ums8ARVSl/QhXhLxf0wwrxJHqKA1EUU5DC2jWjn1lCsxDP9Q2y
yV7SCBlNdA9KFG+SwYQUkdN4jOLbY895WdCAxyDE99UxxneQdYj6NEp7MHu2fin/
kDzG1nACpNi93knqC+tZy+uAV5GtXbZ1KeMsxZvHae8p9XOOR/tOZ/EBRsDw35hf
iDZWfXD4/zVbhrP/jbK95uWOPvNFRuXf2OQp76y+lZ20XgkUE5VFm5m5MHe2lNkl
Dmhhc149IoHLZslfxQqjdXIhIhdxxBvRnmIkn4IRlZej8FnBQ+Nsea09aKypDyx2
Xzk/uQOfn1tRUwUFkj8LU4ev4nweZnQkem80Ykc6INDK9rFvQg1A38t0H0s0J5yD
1jdC+HsBfAhZ9Lk8sK6mtCEZRQbjJSLO/IgOzDLREaFjaVS/I2gPwRran+b7tuQ4
0DMs5ASf3SxW8FsUezA2cnlsHhZvy2fzFMtznyirVzbWmTZ4PdCZ0D6lyp0WiyX5
Qdy0LksO0Nq0Sza/lucJGlOK5KjLBvQGFTcRcTI000x337gEreT+e31poJrcCLxW
5Ljjqh0M46d1K/4N/6VJ2g==
`protect END_PROTECTED
