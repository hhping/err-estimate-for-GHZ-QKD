`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYXC7ZncDrWeuv8q6T2QmtCCzKQY/bMCHvab9/o19R7pNVhFQz9hH4Ao6MLlZS+8
34MRMktZCawnRbttYQsuJvNaTPV2WudivkFG7MWR0adhYxDLu0tgaqWa8rA/Cfsq
HoFiYjJnx1HXyqSw3wwGHfMqmAt9hDoy8z3gz//k9VB6BwdzpIHs+WZTUYq8fFMn
lNY0kYMZrct3Zm1q16Fc9uCea6SGfAbzukN3Sr0KaMACzZSLsveG2Z0s412VZ3NR
UA8Z7ky4XojmYTha7qKH7FrvJvXwQYTDYFRu68E9FPpkcieL6TbJD/HfNP7SCmmm
FRLV5tabKGp0OItUIPPfLGyXtJ+sDatvITZAyuWf04UY7i+h1Cy/sgxkYgsNHP7p
fDQV0JREHTkfuXk4NTJaN0KlFqg+PJwLW36X4EKpd9S7wXir03EBNFe5/vo7TCod
BBkSNpkM2JcyCnzbfXoNRKgOTgffAp1JEoD3Aqztqe1WfAY1XRWv5nTJ3wr0NXI3
TcbHCahkZlXvKZBPf3uC/idmoDt2q0QgIYtNB8Hisz3uCfZtGSK7MoVPu9AhPMY9
6XOlVUKl6MzbXfSvW2X78lBwyhGiqrjvmpOzchOjE0vnfd23ARuYhXIDxYO2OIWU
OVKSSx+RhICdqsxYC69b/TX7GcgJC8KAEa6n5J4XmpwNd0eJjtDgE7T+P7ekQ1sl
8KTjt5bAMvbb1GS7BaZ5YA==
`protect END_PROTECTED
