`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rmVGIDeVYcn5kfbzNvvpToVfgZfKJwAbvNQeKpgzBD4vbHd2o4O825c22Dly2Uq
eum9fB6rJPle+ovBRXexBykPclKyz2lcCD9px9VruY+ukMu1P2KnXSei2Fggcd9A
gjJ49v8On1cB8Dmo24QoAdRDKBRvYpYXo4hzXgX2oJo23KMsKL4sJ0+TVzyxsO3/
pckjIt1VsWq4vCETW4MD8qwif1aPyC8Bin3yPlOcOy44Wq47orXoVWuLmR3o7fqC
zZNF8mqLGTz0Wg+PPY/aPgI40iyeqemD36yfFcQ/vfgR/DzX5ygIpGOjQ41cnNfe
Va9O2xlrzqws5eGeYl9L2K++4PObjtwSMUzolUG0cbTIYSOexhvA3Cdn8uCI5ZfI
z3v9L1gew2zjPklUiFXhwlBYmTbCch2Y6Cl2380/QgHbCMg7O85RsaJyH6pJAOHy
GBc5JadVarA9D8AikjMP/EWr3NnlC50tyrNUUFTkj5XmPURs63REcKMLbESnLIwR
hKkIZHLXKUPhwekGaj74yAbyr4G57mP7VNU/4LwL7LA28srAmQVy851UbAhos22e
`protect END_PROTECTED
