`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrKt6ejtNjaj9b5JVUrpL1+A0jr/MrofhG3e8u0U7ZL63vG+P7yaej6/yuWZlMMT
hb7fTBCz8rRGco3vGKBydsec5dLM7qnbhmkApp9UvFWF7ZibJIE+nS2BOSIi3ch2
skU4nOHErkoaJSYRep1o0LZr/Iu+vLwMxceKoTCGUnc3V87T65GqUEYmlo2iARiV
2j1NQf2a3BSqRjKz0cUDXw118hTZHo1bCy1E8YonCzRQborB3njJOJ8LZRx2eTdy
wloATPT7vWRFTR3bco+8p2f2popJz0XJjQ4MJrESrwkyaDl59DBcMK++9LHKf2Wg
+Cc5SVDH3SPH42neruRF6l6Se3Qrwa3du3sCOOpSlYOJnp9EooAO+28P4tXCRUBv
q3a1OwHfRCEgKJ/ZwCqUeFzjg2t9QRxPlqih0Hop9qqIP5b1MnUBBvGFGQoY4oPc
BlnBYFeEg/HipHJWqTPKaJCsDkCCA6mAw+KtQoTvhm/MibG8yyaS1Of2kIyX+MdI
UdY3YgEeVsFpe5sk7wK1UtsdMrRy8AA9P82xJW2SrEG6TNirjcJjtNW3LWyKsyVQ
3ro74pkGpEOPCWbcDI4qyLCaTBPsuo/5ipLgVi7v1C9sOkrgaaPIGpcXF+SACDgU
OrifraS6qTVlnsoTYveV+uvs/yz2OQjpDnyyUV08vfokOWuFZ06VADvKTm+HVKJ2
Njv5cav28Oym6fwLkcn42QVcgwuT+YJqAlavt80/vqlxJ8wMHoQiTVXK9D7yBzFw
WM3Y0M0n9hNXyUkA2ZBoSOBw8J1nDSJUMbVP9eVbdCX970A7uYQzHN9iE0LHD/nq
tsRE38ER9rrHmDEwrVF0LaNzetQ/vj++Qwq8ukp31xTP6rIv1Wyg2N9vsbC3g/v5
1poHWC5miDhX3cAIPsK5U6fzWXYK8HCj/NBkAISRgvSTQEYGO4/WT6OKHA/qiYWG
UAs2Ce9JEr6/5v17m18wmFwjigqlp9YNxaUu9CIx+N4=
`protect END_PROTECTED
