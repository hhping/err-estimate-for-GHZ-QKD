`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tU6LbhgytkQVudb87fV9NUmbEdATU7UxHy9VcMDzLjjg+0hb7A9q1uKn2qkW+XO
z06f7mgA3HgviGkyndEi0f5JH89sN81LVz7zeE4kA8Y4rG3UcQmBgLNJED/g4/le
fgenEqje+WmIeBZncTo+WphLT7ysZydtLjO1W4lmRKztcaVfs9Z9rgxRfQydULIn
hMjlZrKtgaWhJ5CahZ0Rd0vCURhmRmw8P+gl3qC9A2FVajLiaQ+mQzAtMie9Pz0y
RIF/MxLCXxb1u0KAgz3pVJw1L1R5qaWx50HAwFmJJIpMemNMBhU2LT/yS0zYZagl
lRB5oHMazCiIN5lJzhQ2sQGfSjLTL8JsBqrZ3a9T1c3rJIzSxJd0Ec3aFv2nqrqF
`protect END_PROTECTED
