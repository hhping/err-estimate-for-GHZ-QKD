`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NL+3NqNq9II5uGxpV0VnMO+CtwtSCNzxK3T9Gewkz+KCBvE0kmwiNk1HSjRsDEQh
UAMszUgSkWQUqqw4+s8laO/Kz3vjc7CsqXZCapKZSSidJPDx4Jl3sm8Pgv3K/c8w
oos67bfR3ljTRA4qb7ilGtLa+kndEnGTNZ1xPRIymRbhaY0bM00caeOA7GDhC2Zx
+JjrWraK2X3QpexfzAU0xLdhdv841n+XgVWX7HljbJyClkvAaWBKwfU8KmCqPARi
Evj9scGBEK6IUclxIRtgcrb12rYckFGoPk+b14qZfu23MmMJwy885VCl2uKra9ZW
5uPk+/hgW3xgz4IxyB9/4f0137AusaO6SX7oh4WMEk1h8DgKjjpWYkX6TVPQf+Qm
vT7JifOvcTA+UANQ3GUun2kC2fd7kgFRyMUYUM0w6iTog3oxXeH4STLsiYf1BFRm
4KWGYDE8/XrK4eAqpxBzQQ==
`protect END_PROTECTED
