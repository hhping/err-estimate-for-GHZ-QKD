`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/uBzl3xPHcSTLQVeXfyLqStnhHbI3S9feQ7GQsFhufee+H/w+J3Z86mTUg8Co1f
XCoiAQwrnTKxJXphYZVOuTZTfS69tgl5789a1gRh+pHopboR8D7DtXDdVU9M9g2G
F8y6r9a6MTxa4DVo33REefzyVCSqjSnMJa9IrHUlz68wxENHitpxbJ5aRFphC1oP
tI8JDFebLnEFyjVOseO+58E9QoW+O9A2ZRCw9gxWDycfQ5C/VHFCF/IjBNYI69Yr
qbC+H/SS0bQCeACdAXhWS6eS+9L6jbqmt6x+4oHNGy4uDmLlPZvROoqmnM0KnWFK
AFxGuP6Ciu01mGgt+RTt0e2tKdB7OLRjlY1eBt6g9ljNwNKgLf+dzgqkPQnAB80x
Zxh8uQgT23feE5ZezvaMK4CXYi1FS5m4+AtPLwm9kvwxcbyHgKTzFMBMiMUJIOKL
fZ2E5L/uFg4oy7LeV3Ryy2pdVyOvGt6qXAlDvsS+FhBtEJZIv+eLcHiiATt68P3R
yhld8rNV4V8/Z6Kr1LrMCaIaWR+htLLk9k4J10EA6EThV5cn3TTKjlJLTNte+45L
+8pYwtvn1jFnZ4HOKLUjkUWQ6mxewHuQ7jCbDlRnsiO6TKSYfeRRAyvWD6/CI4sA
wRHfkcoG3IgL31pQ74cjOOo1rwbJ1WdBPx+FVobu1zop+59RoikEqNxyhuP8n+qo
zq1I1pf72F6s+AuVMTZyHtwaCzH05AdReIgJgBNybBYiqIxT4FhJUf+90kY2mXtE
pUHWYsoOloJglhHf4WtlV5ykFQy3jNUrVowkHNjZgAx8Ufq7vuyphU46eucs4d+f
ViJgfb5+vBOT32GdLase+ncTzQt3OeGwHE4OziCViad98OkXhV74Pn3mpvKb4j77
FVqW/IQE2EL1QjyzIXN+D4SoYW096KHnnXu0GpoYmh+hqQV6kQRDagMEB2ik5jEj
sxfYUjk6pjXsawE8pEJoEUhsNCJXqILjBjrJ0gy3kZC9l531TUn8wWUxBuskAo4h
cFzJZuI/nM5wYw0C3GIboXXLkqF+5YUhI6e/q41lh1ZeRRG0lMzRDAF+hXilkTO1
IEAE76fUMPg63N2vYPU87sWLoKDpjyC5vGFFl3tkHlJES61nUKkHWYd33+7iOoZq
hYLEgd0esPYl87SQEZ10fx7FlRP3XaKT4K2mvb4RzbVQoz3nCWIpSNeSOGIDoVa/
aB0xLNIx3JMp0IKZhfdOp+8qhwOfMBlBvl2uGG7xfwLFQZbYL7IjQvTtyRJhbs27
lgnllXIBCigkekzTqYdepOHU/CEZ5zmBDUg4MxEnC8t3jT3++XXM/hMPp9Zr9zUO
TUXSNCkN+c/IYxdMTURnE5zyUaMfoVfKXf/ydD21vKjFv7O547k0jvqtcDDfhBbL
pKmPo6SdCeM+4tehiLmD6fkPjm4SkXr3Np6lCiwfv/SBLYCuExzfc8X2CZbzRPa+
8kvj7g+hbaVukVXe/aL6d/q5/bdEKfxMvO5nY5dmAR2b0/jt4PQiPxecAPB9+Ao3
xOrNRz+4Jgs+fCV2ttAeQslZTYmaF5BFV7jG+pAl0Hi+6njamonkrOEdlYB1jD8o
EPwrnyHYc0TdrEyhQ4ZMHUOlzpVe7Qu6zn3w/DmUu+D/m5P4iWDniryLmjIn9FT4
5ZZ+Q4uhWgYAwuSJhk90VzJqSJafAv5RD0Jm8JVIkVe/FczwfMnJi+Jo/ayGAfcz
51Z7csKu7eYNeHTnRt7WFImZ4uh0LkE0kKrIemNjiKP3cIJLTrn9tWnCq2QEfVLX
PgEVlwW1tyxosSRlIS5RE5V1qPsV/IyM+SuiVMk8VJP0O9Ak/nqzPnLavsRT+pC1
HqoanjNVE6+P6kD+6zxXmNGdAXU/DC9x7ScdzPkh2iV05sT/Q3ygbeIj1vwiXhlK
kg1/Q07or0quW7XG5grdf3sPOpYMJ1Zz2LSDR7umRSy6X1JfqlqlDDuzqMhxEWa8
SyzjUPT5QaVDzawqqbxXDRlRCzDexCjNKwOQH0nD/Kiji21LzI2glWsr+lsfScrO
oQrd/HtJLIkBYUxJ0VFmCTm1k4bxQvMw8uqqDdBjbYwH20XuskuBV/xF5ZVmj19w
qUn7NpK3c94WQDBmqeaYv9A8r9ThQKJzL8SZKxt7NyToTcl6etveS4XOXZKT7Kg+
kMbcAXTymhC+N66+fN7pAGdb4AWWpUnt0tiRGff1MTuF/89Y5/4qGkYGCm7bPs8m
Jr976UiQpJmdenaDOHGOtYNhhRdH+/I2IMy9IOsPWa2SEy4OkTckZUVFCRMQIbGu
og0ydf8Z449o7HjAlesvv00UYvZx7MbhQsIX0yws8fuadeK432u25PFR5DL8/E6e
w6TcSq1XaPBeJ7F6ExsEYyo2sGCUXH2ALF9ueTxMiOdU1HglC1x9A7qnYbMPxlqL
p39+BXALXJ1cc/Yb4v1xYZmWDlBcIUJXBqjvJlrUZuluv2mf6cXn9Zbyixu/3m/e
3fqs87Be472IBOjwpGsiabI0G7q8yqi9cn1a26zdfl2Arzs2wh9FUdtoTokxkH3O
237/0x8NbLGaEPuCCr8WvplD/ovAzBhLKjddvno9pP0urLEHZVjFV+3Zk4ff3owp
e9nEZcdpfwteLYRnuA1EcCQqNeDWP58MvuOgg2gBO6WHPTrrG7tO7fsBmzrf+3fj
sYDQ9/0w2J82A0rv5UD384mHUJyf71nYrO0oa9k4rSTGfNRrxvd4+OBH8CYubmO+
vpxJJMQMKwc1Elaeg/otz6aF0cCd/j1Je+GFHHjiAvH4ikZ9ZBDc6MPE13QoOnNG
zGzcT7LKvFfvjWE0i5SltlCgy0reTOCzAXQOqqTKs61Nm1HAYSrpJCemogI03Ljh
`protect END_PROTECTED
