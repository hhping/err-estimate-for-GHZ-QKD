`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3O0QFSJ1+immgEHxneHfIqM71bDLHsj2mwadXI1VAgPACTL2KpZprHvsr1BWvde
yRdgUUBNeTWBus5WAlIg78vm4WR2I5ZKIGTG3ux7R+Jdxg48avbIxIUsXdhZnMyk
l8XBUgXL01Q3XmkBTHWFhwmw3GuXMZkYoRNBGAqP2VAJffRDKdJrGEXn5l2rWCOf
wwo3pVU7AwF2+A3nWhcRWBVOxrnydD8UM8aQ18nJPr+U2y1E4cRmI7oblEkdDQ4J
DATqyt8sOOkZmLGbYMCXI8qITJPAEb9VVITYrR+d1mxJXQfvSBtDW384hQeWQkx7
zX9yKYKfW9aZvPb1KaIrt0v7DMB7L70xGdqd10RR34Tl5s0Lsia6ZRPtipIlclUu
GVkEN8Kgo1Lwx5pg7ubHkkjSVOwnZhV8WwyHzyt9HX+uJBhpRnmncxfQlQCdWTVQ
2TghYy1LKS8uKwtJIrRFzVuOHrYL3xjzF/nOOL7j3dy1bUsvNC58Db3sD1ozcE0H
AZCnmuUS1oeUbhP7Ar51+IA8IKK14QudDO2qd3L2keADYr8ITIaSGzROKkvYWUPk
ab+rcozXJcW779Wc5+C1NT2sTR83zVFweaqrZK/fuDARzW4VTiZZ5h4/IANErKkL
7g/M1o59+bir3jjhA3kv1LvpkkgbD743OxhBh8IdGDl3C/aTzAeSTLrJZhj1xNNu
d22QA0j+hYEjHZsDyJeIr83QUxqqWuxXY0RCvHR2nbhOiQaHau/IIgllFYmsMS9I
RUK1BvbWhVaTaOiPuQC3HpeJrW/f9mMdutkxhh1Ep7X0ocKXp0Ci6YRUEb+AgT35
Gw3ALOwpGbl1q0dEaQv1235kgOBwhM5vRFaCfDR5h2wMW8yDKUu1CJCDfzjskLPL
9QfTL90xKEHG6TvsxJwi0Y4ItGJ2EWdxcgTovQD5zzfRTMdOkBy9PdgnqxigTUkZ
G3x01PI5+q9DJsRGT74ve371xcx5zc3Ug3rB1M0kfCzGj2iLU9VhLPRHp3lK9+jw
vvc1PY9lx2/2dXP3li0Mqq+AHhjnoQRkQrQK2NQWjxmCdxMO4rRGqaMWHfNb5S9H
mRtlMVV0ZOLsC0QSrgsZa0/Uk5edkcMfrWQhoCFQylrZH3UDVEcmfLlVB0381Eu3
5cjgexWeaoX0pPcOeYM0+Q==
`protect END_PROTECTED
