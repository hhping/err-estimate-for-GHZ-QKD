`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXKRwuLbZIzIOIl9JKtht6QGY1wR+kt2Rr15Wm0CC/B48V/9RAym8K3jdEMafEBs
XM3H3quX0NIgCV/nwZPHGdyny0QCJBnU5OJgYmzYFFdW9DawoEmWMnxhnGEppSrg
Fz37x9E1P1GBH/jmnMHd1Gt3q0ttbQo/W21njUgg4ZlNpMhHS0e/z+TR4YGYH79/
AFOPDVd/i5Q5d2ezdtBg6NJShJCL+yheQdTvXYmlwlYuDu7k/2VIsPfMzoYKL+V6
o80G1xtQ5R8jfjB4auujqOHiN9uht5Ruyt+oT6ervBLZQqxFkGhp8uynybfGo3Wg
yTI1zQ6/FFxjKy2hePCJy/+HfEzG49bBazTwuO9eaRHGfkoT047NfE6Xdf3LpmVf
BW2AGq2/RdgbkQ9F99ChOvUYbY2QNHY2jWof6RSwyaqJEQNBm84tbT/AZNC6Rs+m
l1D7Zc0zsRw2sX3RmbqoeGL5X1iwWbx2AueZRS8HKU+UtpDFa7gVmz2wcYtjGJAm
WRpGZG+LzHhd53/hR1agEbkk4HDlt8Q0btsYN0nn0s7bDyxeVawM7v/rptXT3/fz
GkUWJq+6HlMT+9ZzrCgfd7CB5+yDbmM0mRotce7e4MwQX508hW9BUbpruQ0uJ1YX
AYgh3yrhLd8vE8EDELKwnNzYVnvQWe4A/eeNgsFZFTtl9XJ5D6sGboZGkyvSt7cQ
TreBuKvfQRdyMZxYYu8+kY9U/5gh6+m8y6ErWjeDs0LaGqq6rb5c0illQvn5x7BX
4DPNlKcBGLo5tjGWqLuRjsX6t/8/+F1nByU7Ua7qSxShApGNAQZc5hhKNffml0rk
Wo8lZ+HdD5PtFjsmsCyFTr4F4cS/zulrcoD7eyPoAfWzhgwc47TQmFOGjA3ZPQXi
bWmz0mL8Ad2kxxWccesDmrsLk0rf/Zz/zBkwdl++Ql1CPkr9ifHzSE0ndSrNnuiZ
+wQqn9bLhADuTiLGKtaEHngvF7kYWBO+1fXHYuizk9TWTD1S2s0ItdJjaM8WgqTq
05TPUxbIASP4HBNdNA7B0g5dJ0bfeir10RcLHwlbC7fr4doHDXRJQr4/pMNkkcF4
Xsigek2YnYa3uIU0rw20I7jwcC6KUrqHqsd7p3izdifwTadZP+YxuHjkTutoiZdV
50lY0+6NzqW12ElJbsaHsaKa9pU1OpyK9EokQDH7K0KvIMu0sjnf5SORmfZEfHTN
Bp0GU0wez/+BlplztMvwrCXBpk7alCwn8K/EcgFZtlIEtCImy7Bs8KrVqAONF8oK
+B/HpD7630/e6JfqQhdYb5bMwsx1WOSppv2mCrf8FrCXqqHEIIBlHm47Z+4sh1gw
jns+0Kg5TWMturJpQor3Y+FHTpZvmAu3wpLwJHu72XDxghkTGiqSFd1gZRfha3Hs
zssbyFBLdwfwRWYFCe0gXml0trELXljDmCusk2MdhNLzf6vr9H6gKb73IYvNqgxU
9IzlaFdBuvP0CSh+MDQ9yRGWovygZxbeqLco7SgmjQUKB/udel9ytEMy77dMdZ85
SPGqDhiSU5U1bkVdzWA4K8XEyBM5nhbJD16/LskUWIM3ckFxo+0FpbTZRuALjNI9
KIYVnOxaVdhmkaGrKm1/zdJUo9ZLB4HSGzoe9I/4RwLh490lZ1hI5rBAVpHHNu6n
pBrBFsRb2wStX9Vuj2qN7rJ/ivlxFRYHTJ+Nxf9dlxyMqlvR9ZLEEDS1xpyl9xKo
/eNiUgg3TTSB7KBQ4pILnGM4yRabaNssv1U2Jva+H6Kb+OWH25SoInVzyVodA+y8
XFS5vFUvYyE+u5Aeg4I4FE1j1ETEAPN80l267/j39o/ZO5h16V1vvA3qkSdfduBV
v8fQtOYFaSa1V1Az9MmUaSpqywezvKsemJvUhkkbGs8RWjBUa+KbgpX3s7mgRjkz
Py3i7qFTxi/WhJvmGo12dW2oXhxSLZ3GAkwbdkPqXaTRra0K5n8ygzRPmKQAGV2p
d+XW6yxcCHWdZZRdsO9BYp0NhcW63nXcP3mOWT99oR1O3BZ4znDQB6lCZg3Glc/0
eOouLRrotEJvNTptspxOwJANU/r9tuDbS0EVeYXrz+zELSTpx+88IYMiWiU5vS9/
MP6AjExeHauBNGRAurQMtRJl2P/MWULTyx6/8ReVdJq0rgu1B15kDVycwAil6FPY
lplRywCXnF8u352jsW8yKtzYsPZ5qUPH/U0dAM9QQn1zZJU5YIwdSomv54HNyeG4
dVPvqpwZdvupr7ObK1/sfnN/ek0jbzF86V/tq2pSuKe5iLNLzy4lya9vvc/cViZu
fuybK91mVVjpdlRMETNw1etnVwYbpUdUusEOb2yFEhajPb5pQmiTH3t20IvidHk+
wgLIOP0FzxtQXCbWxvgr7ybIaE/evB1bOTcYwR4FUC9/y1DTehb9c8YPoTp7+OOR
4tIW55I7FEkTqolucAlxpqQHMH9pmahP+dZqD+AiJTjms696i6s9EjZxV0odG+li
PcvbbO7ZATCTtMzQ+bI2/Z366bOCnE8cbP/wY3gCyPRGVNkgEhvoiW6guGVGae5j
+cFG/nAhnBIsEcDwX9c05WfBA6UbaarbHxkSxEHlgdqiFlal9T11IJcqvaJl1U75
l5gJcAnRaja4vquhEl27ZOgmnTdSoq/YpemnZlMjRRGJPSyQcP2CeQs+ZIzMwfek
c2esmDngxyZlgc4Zg4SQS3baoYazfCePQPnAkVRlYTrBFKx4Frxr0X1HINYPLT4d
pb2atj96lNVkeOhW48nDCXtL7l8/6AKjVeZyzq4Va2Hjbi0+bgnzJkbe2Ii1wm8K
UmqtvrmFrHTg3AfbVuG8qsiBIP57Pdo1JIpfSsKGF7fTLBYoBOtiYsNVaNJ9JZkr
qMUpu57GMN4eP/Wmh0i3AQXKtTAW1Idu2lHezXs36GTwIRHSAsDSrDW+jlpKvPpa
EIElEJY0ROJEeztLc6OH7tgl99X/s3502mA/8bLNEG3x6GitD5V8X0IM049vmg6w
6S2xQzPYZp08xbbNljeuW7q7+3byh9PWJ+/O6VlFtdgmngz55apbWcVHC95JLAhW
V8WkN17ul4E3o0b8rmT0Gs+FCfBG/HrIYBgc6ekIAU3+BQD9/4ucLcXe6iQ5JXuC
JtNqZKNKiO57uy6YUR0NFD9ZBqsHdVw/RJ5wFxC1wRVGHza82GeSpOG1/0nUhQom
tsyRfd8jdOt0+7qaj1UQ1kFziQ8bkSnWDBUgULZxIff5kx0R9VASABPQCdgLoTuX
uuQQ5fcOBTuvxuSEgA5La3jQ4QEXQrQjeIHYpuEw1+nrFsK1jo+qN5wkdW46PzTu
T9lYsLc1/SwzZsUZjnb3cSOEUQfm89QccG4MgYtiDr6Pp41Y/zS8+rZrpMW2X3/O
8VB6RWlV23IXPr+EQNzfzZ65U+/2Hh/qiTH5K93bSW+Ryi1lFWzb1k+Jt1mTfGJn
hydpokWTiVyXlYelpSLoD0FYR65lAv3p9pjmAI2xXG5pjM/yX8EU9rK0mtHloue+
AC388JkJurEsnZBPgLfIPQ5eG/pYPVxudXitl/4kthk+0FNd9N6qwVeREPKE/yr7
EOodegMuvD9+/hvONpfrJICexng22Dac9bpm+oiecAVjhCq6sibafYndEpcgvppS
YOHUlJpIfkqNqFcdwjacLOpXwTPLmQ1sl3AB1cA8f4DbspkUl+hYBVMUDV2ioAnW
bucjrfOUzioocex7hfGODtBUs1O+sfi1cKC0cDMNuGJ2AzlpaxBDBiTUxbVv4oq7
2XjSPN0VafntICIbTha3VGIDpdBlTxkHiAHCTVUmeCV3VxahJkvGgkxM5AA4l7S/
AuGxLRfoPhun+tFFz5mQVVyUPCRI5qUVCxxPbx2FvI29MaPlCccbvrBS+mpRkOCb
S46s1S2biBwXE/GnFz7aygNLzQSKt5yI04pmqkejgNmptHshrqTFI2vRptXyt6er
BaQkbBxCPtreDjnEexkmVRXtNjhzWd8xmACqOEmyaRwBo8KYXfIbbQWCigm+iihy
KwZCphm25ozxfLG5cB4N3R8VzpItRlGThx5MTkQqB093FD0VNXpuSIYXfQvjndpx
cZRN23O0zmtlyMQjAMWwSTxleXBIIavNoMxtoEL0EtR9Ybz9k1EuciZxRnIUXwJl
XAJjLLtP/ScA/aj/KWfm8cqVd/aB1JYaVGtjP4BtncfkWkCPCuspr7A6Bbkal6cu
ob0u1LQbsD+zC2CqXEOtjaQhKG6HxKXNAaJFLXTy0Y3AUnI16Z4wzKTvF4sRBObz
CJadlcdfmjwz2SBIP3/ZW7h0/knEsd3IR+wZNG6Pw4oXpi8O2wiTm7rpsenW8oon
g9+Sk8Q8FwZ0uvJL5fSaj4C+BpBQB/lYWpAsKCqF2qG2UIkyTHjfb56tTOhgsTp5
YM23ppeFN2od4Fb+kO0it8oUgZe7omLjx2AgoJvaDMz7LfwZ7645JSXYfdOzCex6
g+5QcEoo5jS8AgltAKhr/575Hj07GeOoGSu73SMiifD1bfEo9VFxN2k47J0IC8xV
zqL2A6zP6hiLCwT8JZ4AK4rzhA8pd1Bup5d3rYUXvX5n524obA2jCwD4nI7ZQNuL
+vPk7U/XfN7ZwklbaJCd5GpOZ4owiI3j+7IGw5PJd82uDK5IQNSMbfsMplhmGblx
+jUz/As5faa1ntfB1NtRmP8Ti7EXcp6SsRG6+vvL0zjoT5C1nNkkqNc+TVy9kHFI
Qpx68pzuK49g+MK4GUGtG72TgUl5y+XNaijmHEW2Cn5NfC/HbH+gcCxRvxq6Pa83
f4dIe+SzHwXVBEU77pChvGQJY0JrbxIr4Y+NDHsotcpbRsbALzeNNJ9V2/u1Gu4j
vGnjXtb+yhXm55rp+B/UGUAsqGlz2j4arUT7VEaJ5V0VmQniNPfv3j4+ldYI2+m2
cYy8QbQ0nVfBtDPkAOWjfwEG0kt1ZxRZolWG/RnR+UhISXODwG61L8b+ruebJ38a
aY/xtI+nkL06y2yRkdEUlM2pLOTaxRbhBbQYbyXSjqNd1MiZWUTgDe424jKLUeQR
k81KrTLH1/oZtO7jEwZO1d/PNtn+4KS9oSlXXNoVyfUfhbQoOi4JZdoyJiQML+pP
XBc+0us5LPifWF3jKjGpxIRNQjDrlMCbnLyJSwrV3LfF+X/Wg6EUDYI0YqUTkcT2
dI3B4o7XQh6HelwFDcuQD8hRun9ZHQ/VqHx69F428M27yh9vQp50tZjbzFde5+1Y
5zd+1KuHiAz5twZ/1cK6XnJZ7uSG1Ovj+QQK0MLGW5wey4irASC3VdmsK8nPB5Zl
IU541z53p+7WEuQBejYO2LsVjXqWlzNJ1QG58aesu3T8/BbSn/YzIw6BX5YksUu0
5z79tQghjZngPKTIcFKnEaaTRdTDqnIyL02OQrqAWABY0h1HkM+HumDLmVb8nqJM
chcjv0LciyerqH47xaIrQcg3wP7qIFdvR5mfBx4kvzI8x/kLa7maOSFB/2jho6SR
78af1LLFbV1k1EzuYIGeQlHij7FkxFlBOM9ZlR8MB1GgrnSDy15pssxIChdKwIFI
vzo8FVXUleDv2aGvHlJmALsjPlqNqRGh4xnYM5ptM16sOHfwGkUQ9GWbGNtTOaId
H4/A1wagkBqqhoaawsoLj/QpYT4tQ4HS+dmqtG5vfu9paHiGdt7kyWwn+3YVXdPy
4jIQRaF4gfHJ39B2dv3sK8TkHVKeNLHT3Ui6/febBzafLcaz1UnfEbw9rElplkrz
n/wLFcQ+FRFqft558vdnCTv4MbK6w27yhPwG3yuTBA380HHThCygP2vZAtIG5us6
sGvvfmbfYOz7B0lBjRzXpvRg5F26S79Ly45GwGI7cWd7wgIdg3OLwskqO44EBw2R
It3jkOGm+c83wr14Zd2SMAa/J5eVS7VZsSMElKMwrKsNTYhYYUUmOo7/f65crguh
Bmug7ynsUofgtv9OJwwOaYoykrt3C2RWXOdlFjAz1/zsZ59PUWdgeV0Dr16Q2fPp
8eliUSkuHih++YJW6nitMUyYJEbUoXD0/xmF5SK3Z/b48QCJXisVuGKNvQw899za
4MtJdsF4QLWwVcUZueiT7VUkNbhltyeTUdViFxE4/O2yFFxy0730qci+HKg9OovZ
zPihHOqhmmP3YwHGeFm6rfakkFIKZ7agR1hRPUhnF+OqBAOELoEw3i5kGt+eNIHY
+Y+nyozSWJcQ86EQkAQxFSICtF1xGfg4v3fVSp4HmVLzbEycSmOc64Vi3ASONO1h
gfGBxCax/xq+j7Ej+RejFO23JdiyChVU6rWdGIZ2RO4a1ABQM1Lwx9gmHbqrjTiE
I+geZQbnsoEGF1rW/qKXHOJs5MryLLnx2lZlOtxDs5Kcj0i9WvbDhvAwAyLxdgmx
mwc9PMnZxmc0+99L62RcaA8uK5Y/yRHUHUXFbcD/7xe5ouTVbQlCxPmQto+O1+Vq
JGbp+JYT2RUEDHGy28fGD4AWcx1+MYToKX3d33xOEEiyw3gWM8gTe5kqPKKNWXiN
DZa+ewbfrf+C6ElvQPdP37qpWgV4AgJ+p6l+gUG44z5ejJ4R6voKjWSjVvkT6pYy
D5snc2BRhF7+Am3z60xynnCpJrHJd0tfsTASPYQ5MnzGPi2DFceQVkXx+n2p8qJh
yEBuZNdntGUZGgr64bsxUf6/XZBlH5+mXNsT6Vv8EFhgqjI9XOh+BrFqCnrQKwmP
eSh881Q9JHWG55HE7VldlipOGXL4fTxCAbpQ1JNyhCBimPz5536s8ek/th0W4Z+x
jf/dnWMlvEDJA3DZUIoZ5Jz6xLiQ8OgnP7K29QccU4CUno87IKS3omcW5FNR9LUR
NCIzYN8CQumEiRX4TeTfgGnaknD+41bQPH/CR0bzWQCyLiYFD4eWdlNVFwl/ciAB
ytZHR7YEzefCAl/w6kFhM8JBqGFQQFsvGiJXyL9cbMTgYhu1JPG3/c4+FvwWPlV7
VIAX0SPpWrdyBkqSH3CcNfExhUsVPkpak0bfsoyfh3L2tYstGWguv/67KiAxJoqk
Vok3GlzuZ5L0V3+lidDpFrPypcyOsjEOArYYLEmje3PdFNq4EMvu4bLhvwgDa/jJ
eHkrJsvsULehBcYOeltrLkzM4Li2bp4WN/z1/ZjX12Z32ilLPRYzVvmabye/0c+f
WtKMHvJvaOWo/ECyblu8Z9Hl99VPWM/OKOXpGC4L63vsCsOGYkJkONnszVecOCXQ
57ALMG5hK4CFQ5HNP2VmZABw9H54vS/jYEfxzvIe3XyqWAEpGvNpmyH/ocQslVK9
BB8grknTg0CzInpuoXu8FOsyG89WWYDqyXJBBzTl2SuxrbG59mkQaUak/pEo1i0I
kEhm23fEyJj7z79yhr59sDk7yTJfr9xxCqSJ0eWg+tCZd/DYO1rxbmh1LQRDUZGh
0zHORjeC8zrNcsU1pYEBM9lYF39mMKtmClTeLILtShBG+6ayCASFX0+aGW4eHtHY
g8z/K490mwgUNsmheMFCwpK4pm1iy/S7AI9iUcC4eaPTRKpiKl1M7Wa2XF0chqlC
9G08z1fNrMdWC4N7bLlqHdI8jEGDIUF8LJvNPbcJrzuS2RpJmwZJODYo7yJSK2nG
SQ1FeIlmMM3k2uqeqkTZQM05ttwawKcDiBHClqxyaPFKBT3Hcg3JkcdfqY++MTCO
AnSfqNWvlVsRDL4xDNm41Avsl3PaxSdWJGav/UjP12fdL9uG/rB2ISglIc2Z/Ifd
ADknPBRnIvZ0VnQR5vBx+dx0vL/Chsfh0ykNoUknMUc+e3v8aCpj5rCFGNXo5oGo
crspuQ+ZPi0XBTb++p7roniTC6eHn8i+HFnvPYES2azBFAlzZyFNqh2lWq+oKxiY
LBYX4bTaZ7yfz3qM57GN7OUqY8SuShQ3emxUvKeePBoF5XB/DBUyJLB7ndZDT+D9
VpizSMJxzpCKHAdsaN8H0TNS7bNUY3HybEKHBI73EifC977PbK8OxmQDKDGjiaE7
P/TylGpIezbebzCysDq3+UwcdPRMLeIkfhZBTHF736KAn/3T2sj0u+zMX/NjPQ7Y
UKR4QCPrChnzbdOR5sI8TRI8WMKojhAF522tRhCLf82OmhyuLLwANMh2ziPx9QQu
dQo1/mLpHShcF4tfulKeJQZ2lk5jdtIN0bJYpixJ21A7GWE8itJ8ECOxd/fOo+Jm
HKHt2gIBVzUMp1FgYVuEVtR9apSiAZRprWTZJ5u2QGZ0FilUl7j+lk6rpcxnypgf
tdaMlrEwSVqaEJDOOwuGaBMAJ34Yf4JM/ej/BjEsetAPw0NrMXQGD2e5tC2v4C6J
vmX0uoMwwZNMdtJ3Q1OASnYRpx0BziSbmWqB40Xpn10G5IF74v9JZhOTpGKitDZu
B8TQYpwV+T5sIGlWJNWXNo41uaSpnniisdaAYqKrbyI0RNhO99diYh6I9I2PbYlt
+FHKJGORD8VzlE7BykF/YYJatnFuSxcM/zVd3zHMq9rScWQ+LxmurdBfDTvw6AOp
q+PI8Clyt4sB25Kmb4fRMUA0DYLVmA8Mw1sogYTHc2ZUG+qiRd9/+qtVAKYeNVI7
7Ka75ZqXSlHE+wJFacxGqt/p4LpstYU5/IeTxcW7XyzT01BehqVhy1UELs1NUO7L
r26626gXCqGJK8BujsRUBmdhMov4sFwGgSZuDkzxvEyeh4XllG3Wyuav37MIVC9Q
+7vIYIbkwHBoYnOSpvvHHZC6eLX/sMJrCuqXYGPxLOhjFebMynlya5KqK5QqSmNM
4krF+5My2jMvjQ6sITttl+5mXgVRuD9fP2JogGUUT0FsmRLeYzEc2N53ZVJA+j6K
GvOudF1XXOr9+CQqtpJy9xix18iaScGt+0ufXULc0iC6BA6uNeS7gsEN5iSrNiik
ps/GD1t2ahykdFAHkprbl6QNhrl1Godv67FBjg5CNjWF7WDdYJ57OXwqzo68z5ng
c7DrOBhPZZhfZyE1dbKdGxoUpBN4oSDFAN143E5EzIY9mXdoY/aX7l7rRHIKIaZc
xGgWZgFgGSObouH3KconLRAFqNfB7+cRvZowYl9e6KrVM7q1j2+/Tf2vSnMBqQkp
NGlgryDqMVkXKn/4KJOH9u7p9P0mZDZS1Pu61zhpXQEyhjmY7d6baUl953Pv32Hr
pen4Zyq1Bnzcl0ADrnmeOwnU+2VKVN6y84/4QvnquZ2PvAR2KUmeuc/GusCIvOiv
Trtk3E8tdKn9Iue39bIxUZIs9reGqURZZbd+B0HpAWThrCIOpAKafBqhvlSZy0LA
2+2Rsrn33Ljml3o7jMuQvnD8m3jPybjRyFuZivCkW3RqefOwIKOShfsEVImryfYu
JJHRdgpQhK3POmjRcQiTFqiWf+z0wHW96IOksRCSFtUAE4ftCrGe3bFugAX9SvUg
uRNf2ljH1vz4q42eM10nf6CYGBiO/vySFB86Xs4lplGvrcwvYJNWAQgttHEMKEeP
pcuIeTHEBf9GNIhr1KApNYWalOFe/mj7Tzp555Bbk84ivalwUwT/MekVrAu6UIU3
JplKoFaroPN2ACDo8cGBF/X9khpUc1r+P8SsOdz66XDjTMcHwaGJ3rM7K/CqB3Wu
5TsfYYkkeuHl3ahMwsKHRDbcP+p0zE3S43CdugJzHHrZkopt+jTttbBhiSt0V4eh
x0mqd7IqsAVcH6ith8/JAJk8vmdY/Y1URyoGNdjT4Z8ahcjX9XxsxjjKPDeTQ7T1
uoBVXOowdMbOhLEHPHKOYpgKIpkDEuV5BFKD2go3LK4sBJB6oBK6MJIPVKiKnTYj
sreCDa9aq26baz+GT5WEbUH6kuH+58CvfNlW9JDW/dMAb1M+RsmjWha9byUMPD5s
v84EPBcDyGAngLmYtaZWJ9FdJjgkGG3oSK3wXCxj/qzVf1Xh5Zoa+wA1O7LIIApL
qcpWAYNipJ9S1OLg5WuzGFd/QzMJP8ZrQqD1vYXgwg6j+PlosyESRk7B3DW3LdK/
PdJCFUOIuk9NHyAirqLLVIm2gju31uAnJEoKbtjy6K8Es2hgttQ4wNS4y4S+nQLZ
+X4Im6BQXvdGHk60ejPY9H6L1MpH7f85obb5naBse5zO3qxAMX1RZS/b/uEIg8nj
+h7vfmXnueD3wSc8bUJDMQMU5vW6X5+J8m74a/H0APdqy8TznFlemir9CipLx+ci
Qe6u78OVuWzxqxSN6In3tv0h0ZILB3uuQmVDK5i+4g9gEbQb9NBhn36w42hxp6YH
NgG45KXh1I4jKMgR/JnkI7qbpTMne8wTX79KlLn5T2fwC+wcPqgj4xH9SGC6sPgD
trtwnOi3SWqtYtHIZj1GOYIm5dgY2xEggxa9cmn6Gpc055CiT/BRo3OAE4QW3dJW
Nv9Y/FJhAnTI0+lLAb12y5LK+0rM7n58Nz5hdF+EHlRr6wzDA3lBMhu9gE+Uw+Pa
FU+sXH8dSNgy5ShyQS26O5whOWwoNFfcjrgifSnEH8CA4EoMV8wYhL60ZDcfbGdS
vNhaBn/8Upy552OxZ1JbmdFgFwW3GO+TNHNJp1pyBikUZcdyMXF/eT9rPohB1tMN
Rb/9cbd6U8WfVi5aXcBar9eu3rvHnihBDyuRYthZqOuHpo7QYn+OhIy3i5rCZ+M4
5gkrVu4g04TboyPygs58Y0wu8Oj2u9wQeQAVBM4NFkaW75r53ZQuZtoBNhLx0kc/
urMM5MZYtKYeRvuPp2TZNQX2VSWubsq6Vl9xStDs7JScf3VYzF1+vFOffhNsn1hN
w6miP6Z8VPqvFrv/QBpHYW/4JSJSwpfXF+NgxBe3FF2rsniBzmyPw86JktT+ksb7
5vK/fstKPxClbXaAXcJH6dSWZcreNc0JaosM9B9DfZ1gpbHMhoyqEzQVyeOKU5mA
ugYXsPLI99lHLbsqgO3X4NIyTvgeZAm8lrCBz2PxvW9cQeuomB5uZp/M70p//IN0
osH4m/tGqZB7bmwhW7E9bZ3MJhkAYykDAyF85f2zQzzeiOA5dQKg7K1YEiRHFRTI
ZW2Y8zHixGJwd8iCn6bo/Opmbpwjda8TZKm+QtUIsXf57NU9C47XjwuP778GF2Lc
kEVUtxJv+xnyjXLv6uAWwkyxpEY33Q3UKSBXGG0vv8yHebsPZnDlbNvxXQvB6MZz
9usivjZvS0bn8fmccgn+BLg/e060NY060usDw1H1iK63zvMtsxjwHmOYnUwNZyJk
Flwmwh5Xv3uhbQ0WsazLr0qMPGXWqNgC5H/JGByXJhn13Bh//sBbyYTddVe6/RTK
mJn9Bx6dXlejV6QYJXBfYtRjlGoSnjxCZYoGiVwhTgCkpMgWIHPAZozl6ikDzrRU
zeiUATK8KL4dKavFTY0iaoLco4Pr9pK1N2xyv8Y5+DSODkLxUICKOUVvK2sHNRAg
iiygYSV9heZg9KOinfq3FtcSncS6PFY9g851oygaY11MZLGF2d8mYKPUnQqSk6tY
CkbRuu4nsod2Zs8GcAP35EcjS8eMMfjTVVBSatgDi4ropfy6WtD/090kFs1hcJ7+
PbTf7PWVV3G7/TpeatPV9y0QIRdwS1atOUhxCtrPR48dfnbH7VQPVkZhsEAKXTi5
`protect END_PROTECTED
