`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/9zaaGIEiBDoVP42X4qe16nOkNhflNO2WVwjA57bgNRoQtMwlxgB5AIV5VTY48l
IsBzT2HE6E1D34pytBi6q+kVs9NpP/ZJBuKKpNLTTYL12natf1b/+EmNuFBP1P8j
P0Ldzv1hxrCGOC2+ZMG5tuiEjarLdDBnU2g7aSExP5CAk6f2IDb2ujxljlQF4tBX
9GsKEF1uaKOuBWY7W/j5IatVw4FdpN/JZqLspuaMd/L4LKtcoB0J8/LHUSCvFHFM
ynfy5PIplSAz6Gtp2S4sBe6bI6fRgp4CR/U6y9QJCUY2zeWJyNwv2QjYY5B89irz
oZN74p6hmDOc8+xB1MK36vtojQVGyh4/IYeLLb3Yc7+iqlaxdN+hLVPw54iT+5er
ZZEMli1a+IcFHYtlQOMkqAavQ06THhsDoLcMRRY4rhmJ+G/LciZu3pXvMdc6glNT
vPX/me+aKhpLK9yvJq/y9fAyLqjU4ELsoR8CcVPkITmnNQZ0w09MT/yuOnLg7Z8u
4zw0cqvbV6j/hDat0w2C0M4c+7t7GuqU1S5I3Fu2YBKksLTlSLFIMl6Pxsl2zDYY
xCEw8qaxPI03DzkDW2Okv8JKAqbi4Ci9skS/wHG873hEjskagRrq40A4GZYltLq4
`protect END_PROTECTED
