`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhXw9uWuuR6JNh8Id9pGM1B5gAIvi8qbFKZjOwpdnE3abnwLlTFqPaJPlNiBrdNI
PePkNPPcg1dBQsq68ON90LG3QqppkTmxkR6qJP8qS9f206VrUzggqa2BfhoWQLx5
fwZErRJmr51KJw5YLGNvMAjD28gxygAzd04VMZaA6NHMvtiBJ55Wa4aid3kJC3XJ
rxKIzhhkF72u5iasbcQVcF5lDCEgiQ3oG8y0sRuSvHyywByn/ZTxOFYVudC1WgeP
/2hDO1EXqc5G42JF/QlQv0DCT2PAdItwiatZ3B3wT0ILI0pAehRtjZ/I02Veypcr
PMhUCrLGk45hUMrS2S6Lchp6mVzdNurVdzYUuIfFcI0T2T6RKtfx00t13HOK9HSS
bfFOaJuiMtuhmxsupQArJRgHCzvFHCcrk4T/UXBei8gkWcbAI6UsRK3r9hk/z9VQ
mvUfCWk9r6h2dxnhNlSYKjTcYkxOZwMpXnnlaT2fdy7qm7UZucYpb4J/LQHv+Zx4
AeyKkuOUkTUAQpTzw7C7MlGGiKscbSsfu0Ii3dxohgrvJ81zMprWcp68H/TqcnvO
tlcKvZHh9mmWbZJr40i3hz1/Xx3joqyYlOR0mSYz0oPVuctcMTGgnHCN8DOKyrO+
x63tFGZDakzRhV/JCb065w==
`protect END_PROTECTED
