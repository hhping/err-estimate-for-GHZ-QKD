`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EN/fKW2yEIMhBqRX1ckekxa8E1Wm96rk5Gka6QFKB9WciTiFAkDSfxkatr05QNu
h09gduhEg9wEFUnXc4miL+xdrXEVGpB0/DqgVPH1uOIMlZLJvA7nHI9K++FRCrks
GSQbeBRuzO0TRKZQMTda/gw0JcCESW4e3l+/csPB+JBAxBd+uWBlOv6wjNZ8pasW
C/fdrpbfqQ5Dn3Gi/8Ka5sMQjvhj95yNkbDxj831RKLeTOCS+5+WpB4pKcerGRyg
wDmIUUo40ZFLvQV7Tk9QGrgVEVKx8mwZfily8gWGPgIZa4rlsb8+Vy0BGPVrwGHc
NguRbIXwarMk4vukpg/CSw7EGA8bNLXz7c6CQ1aclZg48mZLjjfCnBC/jV1K+1Sz
7Udbb+FWi/85cACriNhtvy9e/FLddSVXagMMRdZ0DF4vGzRaKJZCR5gUAsi5rKgH
SnDyMn6PKjxMTsoPpVhqXqFaEwyThdV9W4CTxxImtlqu7nr4EDkx/k9Pow6IaD5Y
qTKj34NT3kLQf0lrpQ+5D+O3LBi2zwo3HU7Ecpb0QHvs+gFpxUMNybogJkTQIBKr
mueL6e5Vsyk6XQg8cVbtbeE+1jq+yBuyt0quQfewLI+duxdIO8DZdMPAvvlBo63B
Pe+wb7d1xGj4IHpmoWeyxexDmhWMkYad0eMQ5I14N2qb7NI8l98cN278pCp/UYm5
rUG9PAntlZ0wEa5myummoyApqeugGEpxA3O2tHwLsj+DrDeBpAoNlptiP7Bd0BJq
DiRKjNut3nkxN2maW5zybBqR9z/P9xuLZlfS1ciM1JBzJs5bNsiwRQ27XAZ9PY07
BFIxn7+AYzo5f8YA0cXdCn/j5jiADKQSY+jErBkD5pyLvzv6BPPr3PMdVRbcDQMf
EjaWnn+Y4R+DLEQ63M1bG3a0qMnIEkOESJW/Sffuk0M2xvk4XNoY7trvt/AaLsSD
9ZNSCu1BwJ24bfEciMleXA==
`protect END_PROTECTED
