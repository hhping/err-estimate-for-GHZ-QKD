`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SEarpHoZWWY8sdAQ4Vr7Tx6WT7UuoAynV4aKcq3pERQ8ykpVwOC7kpz2Jb2eVdkU
wcZOowxJECVCD+IC47ij3rY29jbIqCDnacuUFzreR2qdTHKxdVU4Vtty0BDuRh9P
k62io5VFuZW7z0DbOAtZnXscYysTZJsUP/5Hgbj6CNnO4cLKU3V/IPuKOKiDnUzJ
srT/ThRJvtE66mX8FHWWURigyTiXE/L8X45+jbQqwXrozGHJXseZS/74LaKZzPZ2
sj5EiI4k9yyNZJqchnt621iEqUluLypDKQ83b+zOv7xrwzAl3rkJj5cEdW/tD2vb
QI9Rwa5lyIBG8EdwMGVv3sUrMLZvPTQ7KMPUsuI3RETMCdqH3q6h8fv3mAiokJeZ
O0/cu2Qj51UUsrkD2uDaa+cVGGLLu7bOjKCSMn0tTmkvppbjYDk4Ah/DDwrG85bz
SkD8xCvgxtZHsI15pasX2wXMkBl70yRzzLmb66v5xEvfeeLQPr2s9b7YsnOnCGHQ
lQmQLvILWEx/lUs9TP/imN62JMACHTBz46Ou1Md+xSnhKehKIKMhAoKTmc+rO8qc
Pju6+EcTEeOEZ9tjWJ/s0pZVEUjBfCIPsJQPgfS9wh9QUMt1S8kA9K89aEpBmMfF
2xSTS89xKZ2LHb7NsI9QZGQNiL6+IhisvynUitfLkCh3tNkKNQSNtMSoCNsJTfUL
RW/1tuoKUQfyLqCPyn0sjY1hESY6f3ODNsPL89FKReVrUF27d9vVOVeQaVdYmie/
vBAAF6CNO4+XnCmFIz9SX5WAv0+IznhmeWhJgKVjtGrW3/tap2Frgur5uv/CZtx9
m23TxjKLe1f9YEn8Mh/agPw+hfpFpmZ/f0nuudEmoM4b82IclCuZxVCpvigvg9a2
JZdJxgrOVfErpvkdikfL/5vIqbgpYdK1ERZUj/E4yFOo24YiZibyVtKidV4GrW8B
GBfvKSuZ9gi/TgJN2vnVaF4CcN8+Y0MAqMiOA/SHbSSt/GgTqwWgNKqwRUs9cwO9
t+c+uOo7kk0Srd6fmJCZ4BSw1pjbQtXhP6EXac0q/qTZfGItKnvyczEs26g58M9i
tyl8L1IZyf0517NbyI2lUdSkpbcPNJe6IO3VBv5cTa4hOVRtZpzQoghqC7xF3Ns0
ntWjE/a+ef2M1pwGW9mstbGc74Src83RC61Nu6t5YnEPKVtcANWIQsbfzk2z8Nzl
wqZNMryMA+/rW1T1SPRT023n2+MakuIprhMxk5vy6y3+owjHznwDDcXlGqKhcb7M
CknQF42fhCIvpVB/dzs9mK/BQckqltt42zV14BCxNEgjpsMAiBcfs9aQVJI/Uda2
27yxAr/MtfOASCzR4yuLdEP1ysXk3KxbtOn7GtRt5ki+XlxvxAo8kkfAtg5L5pln
lBoS1a6HhEdPKpEFTetmgsdhi2G4wNna8Ht2FIDtMA7L2jglMvE95XSaRxpUCiax
XQ1x7izosnIGsUYRZMj3NgiQMtvA0l0TsSIyvfXRLeys5dydSncxl4+EdwG5Lw5t
SDCDUNaZbjC7mdgRPvPjj9xAm3OV7+DHQrH+GvfC0EOdvQepxd7sr0/G7sYHBZKH
jHR43oqFeDWsXKa1HlAOFSJ01oGFEBD2d2roBOdlugydrRPdjyplZOAVAZBxDFTR
iTBqjitZrwf4A2OHoyJa1DToHPiz0/dMysOEXJducqw=
`protect END_PROTECTED
