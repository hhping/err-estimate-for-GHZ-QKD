`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0SCrIfFnylic6+IRkE0VJujrKRRsDsJmXpmpujh3d4pII6qb60a4m44TvSVY/Oh
tlHYMWSrlN6P3rFGPikVsPiKab4HvIUz/rC4Wb32B1027iZUaRmyU267/4Id0cy7
rjtAqsODj6reoVyyRZel1mRV4VLBTM/hqnXkjdaA+SbTfgkhROMnjhX/nV3ZAcpG
TtHfXpbz9WlpxYS9QfHMbRi6A8q1tpOoszlkJT1TM30cO+M7ZCO8ZHmlSawbaYI1
as8Nl+LdpkL4CEzKIwJbRWW3g4X0iREOl+0RWPahznpeIBRAX3lCvxPpSFD0oneg
/xl6eJq2AajmzQQsrGNru7ESDcSJIDYR4KtE6HAKJjj43TzAW2JCpfh67RXS8wsF
5OEgYkGLZvW3+0NfVn9JxvrR0YVA+TQVZb8WO9bjo7TUq4Uulv/JUGj57uTUtylD
/qdzgvbETyaWBn/OtXMB4Y/zTxmpp69H7sFPy8N8f4wL5667ehmC7SM+IAksY6L6
cg0kfZaD0/tkhFfpfAHoiZX52/b5P0GkCJPIDzFL5Yl39MFRUs6GN2R6c5OHvMBE
ggUD6x4b06TYYf2qLp9wBW1ABGUbOMQ0HezYR2synG7sybjg9+uExuny7rTvQTBg
RzNVWKkRG0Z1FS1GzVYQW6sbLHil9oTqGJ5iYqdcsegijErx6o76m9OH/gU5gZZ6
J6L2W/fhRxsQ2OThb6CUA0mCjChMUqumRHzFlT8DX7NH+TmVpt0swIYEdE1dAhhe
C7Bjjcghlw9fLpUnVeQeljqS1z9t3UNK1qmtaJkCE9SKxkGYVOgz5UWFTFKzXA6I
uplrv0EoiWMp8rkTeOTC+yHG6f5yS7E0+ww34tvchN8=
`protect END_PROTECTED
