`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrFfsLtznECPSr3rBK6wwDMhnpFDJTnRsGZ+GNkovPp+d0AETCm4Shn7m4PdjsOp
qy+m/CrE9TFJVJsiNotZE8OH0sqIiKYRFJXTkTfTj3EkBVkfzqe8kCDH8pN9MwQb
kGo/1+evyD1zCrz+TGZTJ7TlDVXxd27q3B97Pu8i+e/ocxFXMKRkz32PMw/8yrOC
Uf6MkkDuCCEw+a/gYde+0oW17mnyXZ/wiTurlIVjRcZc5ehFRZ/CGtmmgUJaM+Q0
xPc8hkrs7pWirReUhtOcFzVR2HNrLRLev/jWrrXbklLkPZdA8Bhf+H27WKrPKtFY
Qm8ra62Ruzm9ksXltvxH3V+4vovcHF7JD+OmCIIx3pWX09oQigKD1LLUqSy03cEM
adr8gdvQW41xPQCZGsfZlguolHp0Hc2ocdAHRM5OG/m6Q84Tf20CyFCpcTaPU1Dj
Pz+1jAAnAQm04amjz98FFqC3ks9/7VO3as47fAYVXk9tJOstGXqCCg31ag9E9eg2
X4JmdKD25WrK0YXpzJY1BQ==
`protect END_PROTECTED
