`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlNHuHimEsljHgBscPd6sD0VD0SyDoWMIvl6dkQkPunxWr2mlJpXIah5whxawAQC
pFFZt7JyrZTG4JN61NhTvibGdfDeA/eAqrzlBmyg2o/20Wz/t43IIsyofhAF1auv
hm+PYy62ssbVrfBU+TQUdSYOIaTTRuf9mrJIMGxx7BBcECOpPWuhpLt+PCQTS/QP
UNMUTIaK8ZSd6/l7kBhhL2ophcLW5hScnV1BoGxtL73ubgmnXTd5iRxx7hXUvF2G
o9kmfKfPoDbffVkPM7Wp6Sn0/epprPp1zfq0boTRsl4d8x6T5gGQmXdAZcokiWjY
DsGXBpsxk/Tii0usOq4X7zM92fdQm4fAtcBWpbhp7WpYpOckQ9rJgYFPDk4+hJjw
HtFF8Xvo7gAQIr7wFxhtSqaZDqwPGYbJItldQ1VWiWkq+0e4PveM/H8URlBptJO5
uKKKAl8Xbbb8a9nbDOQ8mdSjV60g6nv0FDxU169MFbS6wFGEJhXT3JkEtT4BLT3z
bUG1qTGzmm/JFsdQF4zfmmqMBC9XRKbAk3GOms2kwEqmk9Mtl8D4JroJGuL6T7/E
FH86PvrWaBkN3n3yDvy48szsGye6WfIlpGxrq6iiVAkf5lotQw1LdswMisRD0Bj9
9eVbFfakcsstDSXaay8tq+9mNDzfnq0IxE1np0/hvOXTtDhZaB0EwK+1nbPFYcGS
a3qD+nZDUieeqHiufahX0or9+VapcW0z1noa5dLCRnY0PtFQkCDcIHr4gRoxEftM
`protect END_PROTECTED
