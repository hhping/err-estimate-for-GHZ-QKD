`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9D17JZXSkW2NuWaUybDobxxQ1RWQoHSUKEovp1qOQdxJjCG2fp4wKiUvaDrLVQS
KMoNx866q9qsXSnMbzs/ljrm7Z07ptfTprA6SdnjQkbFE8xbGElV/h+TzspuM0U0
nScFa0pFP0+QtK/eI6eG1ewGmJLiMvT0ZV8peIEzE3sVa4Odmt0zbXczy/uRcgsg
AACl1AEAls43zwHs0LvnW8CxmZ2U8waO8MBy2ajA+Jkg0Do0D90/rYNIObkysoyi
KDy2sbPBOzgCjIeMGAX9ddNU/GRgcas/0j8dan3IW13Jqsq3t37r5bt3oxb7Of5i
7pwqLEbn/CDumiQPN8j/mAK7EAV2HeesdV3mED/iH1g+/5VXdvZ00I9TpRYHN2p7
dk8yLHMNJiFCRaY4hDp87WkPvUs0j5C8PXIvQoeH5nYZHcISiYJP9OFBDeGtDWo5
0USA41W8Pr4SBKszOcUoecRnQW+LyYrBzkxKDYLL9T62jgKHJFMRG0Nm3p9qvW5g
Ejdyvn0S1paOUFE611ChNqcbdL8B3rjIBJFnmh73ms/o8Fh9rFqI7Vwou/oIX9UP
8/eCXDB9KhWVxhjREeXvmQXEVELCj1GRNFEloNq5QTUN6MwmXVizCHcho97J974g
qeNbT3SSQsGV1frQ5v4dr6/mG0SDBonkSDl6deGThrJUUSvJ+Zm1fLLOgCTFLbt9
NggeoEAfJ2reWTpWioQOALufr+ZXqvE33SHKuTyNxOPKXUd0Rfvv7Wv7wgump2B6
MVyY/QTev7yloegLb9cEgHjazUZIOacogW8geiLkncA=
`protect END_PROTECTED
