`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uN6Ks8jpk0lRZBx9xQAg+yUGusoFz5u1aqtG8T4lkq/s+Z8HEBCBbcpq98vcCrzz
p1GgbGpKLZpwyNYt0jUMuQYvngQxa1WnKmHxxcI26MgRB4BD7DPPRllhpf0RjCmI
PMr97AUglIna9vBx+JZzLPRRHxY8R6rhHtB4tPpkcRxn58PooJRsb0KeFFkoZf9p
m2CNoixq/lrTmBgDZCL/n7JR2ytMAbecmE42uHhWFPrKia7vmNNxhrt2RMTV7OyC
Den4L7gpT+yxZWuuDUDb8MaXZTVkflzFnb/GDdUUUJNErkK3Sg3Q0EwO7Uc1BjOK
IlYMwlRtNmEgS5WkxJm8owqxR+nOWlMFXN1OSM77Lc6/zLuhex72iijEFRd0etRo
z2VczT1oTvJJt8HW1F5XmbLXDFUuxyw27iEf3iAIpFXe0A922OsNMlfZjfODSmZS
2AlmL8KLhtyHHxqnlET2SFhMQ/IrDQ7clDsEPObuKssSkAmFI9aTllEF1l+DkwMx
HbqTxgXumbmEHOhg13r1nq7ldg9yWXzaqxXRTuYlle/oAk0AjiA6U9R/jdce5Ow+
`protect END_PROTECTED
