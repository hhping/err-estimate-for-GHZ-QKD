`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/AuDWSrRjxo2Or1zYWmRE6dgNNHYbTaiUbkhxnFQk5hg5snxFdW3YJ5rQMYO7KKP
LRT7K96mLCOMj7EhlOSBtel9uTvTfoO4fAzRreGoBzOUGk1yYmIXrnf0gl14t1hD
YNljxhoK6I5fZO3eQ2dGe3YQDZ8+6miXhBLcqsob1ytSBQtzaj977ZHyA1hVXMlc
khjUkcI/w18bvg2d8U+FTjrYBoldH2d9ACHlDGLs2NhfTUoj6LJT6D8pBcMCGrvb
SXupZxp66vsNdMRceHIokwtwDcjCBtJKykGIsLIA8LjS9fvv2zuikFoZE6rVprbC
/kfSODel3gfzJq4rx+naaC40NESCsNUxCanRnkFe23VAzqUTyyOx6Vir6NqyBCgZ
oB5ZPZqt56unTkYXqLxwYws7mSnWHOqenuWJcazvxFANBVCuPltnOyFucVyEsr8R
V+3xn4KyYXFW2fWFODAHpbnnydmDdwpL3w8zmm2wWklvKjDXK4go1wGpDlhmayZr
dOTVNlVSyMvpeiIoXDvxQo8004NY0WkDJYSI+gHXYhWrEgO2btWHPMxT6viFkUaf
dwgHSSDRRoSW26eZlgBSMdwLzLjMa8HwoPhSYb1WwMCQLzE7h4reL3Y0dMIkQaZ1
yPHR3Mqm6Hyc2NY4VbxNYmWnvPfUWbm5ZPm6gxawb0WkDz7HE68yqxUPfZIouHKf
84VLO/N32+WoYMPBzDv655VH0ZfuoawQaqwRJlvT5FTU1+GsbdI01ztlCmYJpr6J
x75p+rqyrZTfKEl9s1JxiCK+SlANjPh0pc1Hq5noO5sTCq6huZipJFD8754DGu8P
mjsJR0C3iHpB9FMGdeum36RhMhn3UUjZipK3ZS7YkKO0tg+4ddZ/FBUHlUBC8mmG
ei2Fkzfmp4AFJVihpv4VOUv05RAlwj0cAoLOrRdyKUqtQwmd5BaSufb5u3dWbRwY
ydvdm9auCutBKKAsgXTOsAWkhRYl6DuUmLGa66Yafco=
`protect END_PROTECTED
