`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5F46dwd83cUIMrAxTYXprg6OvfPdnnBK2G/fjFY/Gy4E3lKVySg4gPe4BD6MvsXq
ovxJty2pBhkPF7WpgV2EHMVeGnGYy4867CXeE0F7bjNvXgztj01x8qQ+tBDAqunv
naqgl6FL/tXwPK7YUTc3KygnKd8cNz2mYL/w/hjz4JO2whB4QnAiGpVMLkpLExga
4HBjqK8JP9Y5l38BXpfozqEVwvniNhKriWUcgUaObv52z8ViSR+qEB5iz17DDZuF
lx6q4j+SNx8ASjtVz4bP+Jh2fPYKDrrSKuJhHCNSQox/HviPo2etawnldHP54JYu
IE6OaFH8U3mOoP2SGDhC+/zICrTjxhz4Dj4NMSNUCiI/oZSfqQ4lFBFhjXKggPUF
gtesD8WrizGf/n0KGKQk+JlOm1+/ks5Rgu91HeT5YN+OJi5y3LiwbWChAt06vkak
AwKRlFwzXFuFA5oL6JTdz/3a/VEzHiy5tbhtRaDZd28vu8BpgyKLSt5mfVnza8bw
XYAusoOoBXKRex1z84hazWTn2NfbkE574I+BdTQXk3mPLQLzodbTwq6H1hgRKoNa
CXIbQhefjvkVjLEAbUxJrmxoyBzZvw2YqEUi6h1MI66Osi/eCp7JyHaq881xV6Mg
42RPMfXAG5yZllobZ9YMYZ9NKKcFORG2R+8e1Z/m+9JIwjxt+7XlsELtwG5YnKV0
UQicKJUlgaot/xfCKy4EuZDIzkNwQ0khWPGA1E44HY4zABwVDShuSMMXQAEbFCWm
SKV9m8jmkyBHAAlkVsTqXpdCYh1ba4xKtbnC02mkoXcq6qXAA5KmiuJTpwOPefeU
HtzXlhbmZicwI9i5ykg6qSKcY9Hpq3xDIZoaXfVYA810YCoyFAWc7Bdp1ni7morF
uZxa5H5TDzZ20XUaD2WeTFoYEkLfKOrXRfIo6FrtClg1JnvMKUresgPqMyD0EqDR
AzvYrMsLy21MRiZpVjS0qjaVS6fWKTX8zPLd/z/nzWYAmy8PS0pwdasl+pC4cy5o
xXO6qCzZumsvt0bempuQQpR2dN20eVxWbfMCN5weFE5iQ5LwOGv6algv5ZC39YoB
LHgu7CFR2z3bY7+YdFBX1MK5XJBYAoCn1vjVz8j2iyMxj0vMt5BcB15uNBhs5cwE
WTjNoQxngcfNH3rspfGwUmzFCt1mgfKsrO7kTpwfi7+l9mo0vjMl12KDTXQ4BRK4
Xm8VTc7Tuc0HHIVBLA0H4ufxnSHAL73Mg66c6drjDAWdDD+EmA6Ypr1ptqBCXShC
T7NSLUm7dqlEUe5dWDgfTTIROgq1SQTCz3nIl4yhS71whTpH/MCuasXQroDY5B6E
0R9kZc+J3oxZaglLvw2e1pdy7x/zEqrs+jFAQI5hC+bsvAbCwzrYPt9RM1rWxl6a
aHSwT/nuMyJ56smtZ5g4Wk6vQ37P3fKkIcSuuFgiiLs4paNNHLk6ftoP/j1HkHrr
8Ga2Hzob91BWEIIrZ5K21+oR3rUMcwX0AZEoySJgu0araxfY2N7Px4uvbhDdqcGB
gP6ncVsJ55ifBhv1t7pakM/iFwtGbjVuZ5sBcJpvW3+w+Lip5KkQ8SPslS8lmNkL
ES+wAhBrOHOZn5zSPSKP8AhGRzANbutGiSDBTzT/mDQVV7T9IElQm7HvuhvlTpUX
RI3U0XlnUyAaNZjm4AjECjeeOS+aZITq00d079gutwfwvoGHTAwls57i37RwYHPY
JE2CUSgNwXSY5zKzTPc0URl42PNB4/AlRNqPVsTk+YoxK8JuATvklSAKXzAbE79K
2bFp3gq1Ct6VRoOjze0ULGARgDC6o77UjyzDAri/qlXCb5fK3yLfxYQ/FdHxLqf0
RfFzlN1hJmnn1PwnLBh7vQgRWb+I4I0wH/wceM2dmc8XovB4N+LqCC+bYwTW/DXG
LIPjz/J2Lp605REDUD8mWdUnzeOo0NL34t7RkHdWEwcmhAlVESvrc+min9sWxCdJ
Sy4cL7tz1gRBKopGVSVXaAZIQV5tvhEfvnosjjxXe+7XU2Hr/o1Rr9asq51y5VMX
vPd8Mx6NC/hX3Km6VxCQI+Xuwx2Bi6gPufoa+/4QRVI8vKeG/cm9EMxb5i/E/qa5
bkyIUYTzPW8Y2PgLZperYUeeYAPINtAzqzbBtlJ4fSA870Y1IMOZlI/qDw4mubG/
Wyg5+9MsMSxEiKKJrZjaBz9kvdWQppwF1LJC062ToEauOhNXCGlBEB/WvYUQBLMX
+t8mcovdOeZfh5rmLDrFfskxGhLJcZDHPB1+ToY0H3Kk7VxBSvPGpGf2RXMRugCr
a4Pjr5e7sGp09lQWlheRLmCTx0shjpYyljvGBjcQevaIhIjQjbQo05VEz5UTYV8x
8FpP4ee8/D/0BxQMSMAyC6huOvMyGtPsMRrSGSWr7y+ceIhToX79nwYF5V1BLwgK
FNwQXgGjS5OGnIWmmRA4+Oeb5wXsm4qElORKHbEAAZwmNTi1b7WAL7J+o7s+9pS4
d8Zt0FVXBi5kta6g2jEOFM2OeDEuOxFxaAnoHfk+Icy63mPa63GYzXPa3NEoAryU
uaQQXgJ+qOE34tkDOQNNW5ZtLqOwsMsOrmyC4nFAXazZutXHeSx4ZJWoBzCd+ULB
FeBzTZyt2JOo3T/pPfySnwqkPuqZX6Dt+miFztEiB7Si/t/hnfEtTUoY/dCYGjPz
vO8fxpmC4J9DIQO5V5x/cP7JFNrGXicj+OVe8QW8etNLjrB934D9jncI/R2k22r7
jheDpdjnyINm3HqJB4YDwxsS8kuSlHAonEXbsn2lZez7jeOAhs8lO4bVhzW44gRt
G9Q9vIneIQT7QaplkI1T/5FMzpWe/Nc9NwHu1OSTBUl5jS6Ra74BIx6Pgd6KylER
Qm7u97m3Av8oBwhG1W5ndo4aVkSJ4MJBcgeMEyV5oot9Iphp8tRmLzUZdfygXUQ5
XN8pNxcnAa5BIM+W4lBiwcJ9Rjc6AFW2QIfMqVdhvF8KHJRsZ7xaKtTI3JO/S8UW
x3TWfaBATMfFJPbNpuo+DFNa7aLmn9HAOnN1QzdpYzxPIStk+HWkIhqe9zzxrrWP
q2T1EfdQUAtBmbyObaMiBIQAt/yqWN3kxDvj69fE4FC+Ira0ux6ryMF0dxLL3FJR
WP80ufqCE1BZ8qFCLqCoUfNKF7YzqgNvfsExOBBe9R09+NQJKPmNTuCFsUjb5T+2
GFl46rPNL6ESQnCfUjwKqZaz34zvBP0aj+VG9YtOMJf0M5WkdbhoaaYVoLN6DIkf
KUwgOWZNsXkIHXAIOumHFFkxwyytiy2b+Q3Rt4mwaCViHLAyx9jwSRg1rRVpQ8ec
UvqKtScLsiv6ep7/wEB1a8a3AoHu/NjdHHPho5EDu6xraHEegPbT4sVq5G5b0I1e
lrom7JdygOiKrGj7tAFc5VnqCtQ1xxMxzDYWxkTLU8mV6ah+HYLHvqGovrSdZ6bK
a3FpyzfpmORXM1F1nkgAZxlWyBRe1TWGRPRPOEKoaMQs+3tyV9NjKlSYHilFSTJZ
rQp62ZEhztajpbDCHI4PKeDHlbo5BZY69tRHiKgny5t78nXGK9cHgQIpGe2qB7ev
wrQMsdatrklRofXnHyJABYP2ejOT5L44PReFd5HuXX3ciy+iYLY31QUl9tUxvvAW
Iv8lqhgATxiuIHqiB+rO3AiIFycg48jTdPaETB2ljBAmjMoV8lsEbu8eQ6Cr00x7
H+XOINTubR0OT9QENttcxPP+g8z7kXAabfgf2KlizeK86g6og3S7sjMgwuJ5D3IS
+d2lBUZVSRYuGF+X99WIFb4Q7hkdAlMra71WWqUDwN9mU6u2nnm0vQQYlm5iu6HE
G8klSkuTnsd79qh0g6GYd8/ZvVPh3hR/YYTD2rN/lFVi6aGtpfiefwAAuQMQdq8U
xK6dvWzhYRyKhrQdGg94/nn4YSCo0NTQ+dJafppxwreiA3WnxBJzVG8ME0dSnmnN
IGxNxDsqrJ25UEXCdLB9CzBhux0Q6EXaS/JbryVW1kOpb47WiNXOkhde35PGlGiN
oX47/N98gNXVD7spJeeEVB03gdw/w++fqFALOl1QDqZJML2NX/kKKOByi6yfjnyf
YI7Et+LSic0U2uG49Y2pF9cstCS1/r3j9u0fe3bLHbePZ6GaJWG3TrMrdHaujaJT
0gDktMsayVmTaP2VMkfJe8d9g8Ki791p+vDNgw1wYXswjY+ut7zyjB+fqwR41VlS
M31aezG0hHp1PYX1CszPEOOcIfvMTMLjOjVuhnomgC7nCjRF3H48Ukur4SxgiZkj
DEJ6RIcLNWQ/xEA2UvYhF4GMROYB07PcjAI3ggTRawD1shlejqmUG1mBPr7Gbg9d
dkd+KhgyIK//zQzkx11/Gz9A43WJjuK9px2uKyMVV5KVj+Aro96N8Oomyp2uvfaP
qNUE6e9ieXxi5YQZiuLvdZKfUqL3nQuQLtXZifDqgaJi+QOD8Ku2ZNM+aPYtmw9p
Pav+yFgUHeyqThc0Cn89sHoHvw9JZHLGD4R5uJ45SRkHcKAgK38bk6lDMHriJ+Z4
+A8M3HqtpjhRQC3zpz6whcMekEqxUeX0DrtcEPvmNxfZznVeYv/El3l31/StzBRm
VTlFK7kzl/tdrLflGSsaIMbZke7mAWATiF57k6aq/S4yHwYqqJlY9kHiZGnHtfXZ
Wbc1SCltauYv+rSZFjIGR5Jjj1v29qrJadTiRTMDEaoRqUH+YEofgWeMqqtF5TIb
XV0Z+zLzU5XP2WaYDay23HUBedOj4AMFNdEJ9+JW/ly+WiEXfKDl0CjFPDsyXpBY
d71HsI1Bb6smP5wQhnF0fyAfhLlA4rVVHIKt4iF4fX0ex94Ej7zcB2XxJhG+2+LW
Euyg7x4GOJf1eTwOfGcI06DlElDfTsKQQixIB/5/1CKt7tFfWwyIyfrhP72zoctS
95Wfpu8K9JFuIPgGb7pe5OUeWqDp67ntwM2yKE71vz7/8MdN1cOgXBPQiVLReQ6D
aYlkLaUoXKRMNGDjzX9GTqJjk2JfOe7GE+6Em2Fmu3zJPNC8pE5wRNVHW8uIvPxU
tvgm3PXh0bsw7GjwQNecGLpNRV1fUJplyIsf40m0ZQ0GqSY8ZRhpknYwVvalnywN
liqGBcvuQXf3UyGlgLIPWWdMvuDfe9c2HYbUwKNXzaztl9s3CtpO/6fzDqWnqOf0
siSl5DUimjHBrxc7zXk6GlaGNOlZ6hRVaVr/XN2jYi9csxWoC3+971atJAMDG1O6
BOGD/CUwDMN826jsZNeUCDHAQsPlJ7Pwt8TnyF+K850Z6y4DL0npjTewO4G/2oKI
2csgUYTZ7x4+ZffHnb1AX5nmVsDiTdeNlClKE7ZLr0JW3yp7GJDAki4zJVOeAW/E
G9EhMbgLi3Sfv0ON2i3CoIU/DcwsoJOL9R0L/eRK2Ihg3o3i+Fnkkb0XCZsdcfRs
JqaIyrGNzP7sOpEFBLxWHSkyq0H08Uv7+3bKZ/Om35CLYDcldqMRplRShU5qLjEA
1cGcBgvu1bzZ4zSgyznaEu8jUANiyK9qkCSICizrwOZAYmfE2oPhN8KSwdJZCXKM
FGkbdDEWMTS4gQnQ7PtWigRq9GlbX9s6ZMkbyGRiKjnq3u7mnoinZd3tLP/EQgq+
d1Uk7ynKnOTxZGkxTy/s/mKr/VqIzBpI8NYJGvMiNsk8RhDcEsSbAblvuNWJAAre
+o3uNwP0d9WH2GCLNwlDnz0jw2+PAoJEB3iR034PE1CToV1QJaYwHKcWCkMP8VBr
KPK3GPp5BcZqb75l3uEcM+RRGn8LnAKxTjF82LrTGrObNyQxtqwqu6gTJAuU7o6k
izCPXzT9iYMQE9SCa7XyRNpCf5TThebyEYmNnfnREXXLDB1DaVLkDY69lSloYoUq
v4lRmtMhZKbu0kLDz74t1J4AVFaPDb10HCYA+qKziWHSrPjxhuhzlKPUSmWHnfA3
HG5YYvASCw6eFOCPZHoe+ntnEstxIS17Enl+aUwmc1mUft7LbnsypPRVjYeOPe/8
cF9LTs3VvxwPKYXjY9d2qsRpwOrNMkeamI40fET+mqJv+fUXUrqaQbVgI1AdaRDi
vNUEdCpAlacteF/BID2keTfdQkR2BwH/nBONF8sAVldsWOAxk12/vbiDUYsMLy3q
N8AsJj3iMUxHDryXw/eRVhJzkLkalbvDMgB64PHQhzw/o9aArKR3RWqXUPOOtk9w
`protect END_PROTECTED
