`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kr91xNNtqXEdN4RCVzGELLJJqgmwftFFXj3MmUBPxPtoP9f+XG53ue8v79AbsVCM
idhe0poKOsjQhEeJfxnlhmrfJn/0nZ1ZuAGeIeUqgg9bPCdRdM1ya60zYv3WydZa
FQl+N50GteC5EnAQfcPMjQaknTtW6XIx39ceKd/GG67LoQGhs4G4WteCfBEucsY3
xLwhpbkHCcWQ9vIPVHtVyxoIkYRo32TEWTCLSyYuxLeMbIDJPBcTUyP7/Mx8tEbO
uk5tLlPFyjh0x0FMab1BfjLs1Ix1BZorM3+uDJfLoWyydfl6bZ2ZqnYCutStF7Lz
1TiBLBwBEqadddgiEQyf1j5yNQlXSPXEsR0IsQ6LIg/FI8jGfx+lBJXevwOcBhe1
sj8Q2UCh2/aK6D/K9l5lbbKtac0ne5WfSVRcTXkO9+hnn2rJpsuAYop/B/wPYvc9
hju8Q55+26AxUWn6E3gsxYOkZPSls3PR9+HJCkIkCYQQqOmBT2HbcPM0dv0NmuPi
RMnaV6O5bAupn4UhkO/YvOTtRA+OfGACYxvjFQ01VPLhV2cfunHRJIdslf3IXe0H
ii8gVpmmTlWOBf9B5FiICVpkpE21+6GclyW37f8P7asrCorYADK8gs5fmEJkAE5f
8nMtneE0H9qnzGSSS1L8605YUbCfuJrY+QNeI6yMQTmin/EAq9fEvJVOASg7UYD7
J085zq2SnSAMLshRPwuxBvrzvkNF5MxLvY/X1AaKj6+f5iIeP0yjunbLkmcxx3ve
FNkrNYe0YH4HCtHvYEVHWl/A3mdryddFIzacJHsikUW1TpFVrb3KyUxUL6v9/Ipa
4tMbqjaw0Wf6eHe38dHlld4Nx9OilxB4DVXPIIzcdPHBupE/QXLUdVOecTrJaYfJ
opPUhBcVzkUX10Epo0VEz7PyN5TZNjY8LLVGu5UXSgKeeDRCME5N8oC166SjiRdz
8GMVpAvz5QJkH0oZBz9TSlTnQgmWu3yTVbFT3Yizkbi2optc8joBbMt/cZ2uOH1+
T7mQgrjDz7xqST9gXaptCb2Au9PJRW3isWhRIiKjVj96Yxq5en5ZFWh6Irk7x21j
IsuC7AuPNqFNIn3QhW0YCgOxOK3JqIgK312oYgJpjR6w1pXsvY8tjW2HzjclstT4
jh2EmBNrPfZV/CUenNATgBN3InnDue9gmkW874ZSCQIypDQmZ4VJtHrtfVBXWDLB
D5UsIQ7me13ir03MGjA2SVsIxUVeyA3pZ5k5b/TXJVugB9+0ruyAtpZ1f1PRahTp
3K+blOylUseotn9RQ12p/kowrJYA+gA4HAUJAtnCzsuFWsbduD6MwhgBTuOmtMNU
NDWrZMQlGmCQ36P/1yyz3/P4AozxXotaAYIiqQqpI11KnxYpgQLnRBTyq3bc9sz2
I+yHX91QEDakRf63If6Bi/UFsTROsgpHlBNs6jA7J6PE4XRg7FNYl1gV/j7zI8AW
vbyp7lVU7ilLUXHpcGhLKZq1oGcQbeMXJmNt7VTWgUkKFA/ZDcxNFjGw+Ax1PvkV
xa0ORvAmRwHjSx3wtptCOfe4UowVAes3I8HLxQVcten2zpTTEjsfM18sgKzZBrS/
6T6Z2H5swbf+3tqWGgGQtvqNTkqmxFFSIPzxTd1htZGd3No7fBMaYZqH+L+IrrfG
7ebS1q8l/jIIHSpIsRMMO+8WnGWNsYaD5xuewxK7MM770rrRqxrdk5DAFfqe6Czo
WEBKUrIEOvqWBTvUfm9CavPT/KIh5LymVw1q0kIRqqom3Q7N0Y5tXw6u4+/03q92
NZ8HDwQ2EqDc1H91HNIEHOhop3Eh0pt/p/wIugSm2sOya7mTfnVDdA0xSQ+61R2/
7NRuTqfhzgUPrHNMjMBRg7dWU3CHLKqzteGWWKGFTUOUNrtBqlbke+UXJZrXrHo9
wqmEDwdHziApxb/s8LjOgFlnGiyQ3if8Fb7ls2XV7EjbMorh0e6xju5R7QiAYR81
wu3cGRtYIc2nuYC3gT3c1/UqqwLvNoFPSDyRC04xQE0=
`protect END_PROTECTED
