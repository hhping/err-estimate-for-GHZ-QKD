`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33Qc/CW5n1rIa8qaT3unVX7gNyJzKNpKv/tKDb6Aeaz3B94H7PZ8DUWCtHbKe/8U
UAwRf6q7yqjk40eYOwDGPlIwqPgkT5PB16KTDULmRwTrV8v6keIG55fh75En4rNw
dQJAM1CGYo0q/ynENv0I6A0KCa7gXmr1EteRp7GhsAxO+A0lnayBINhoqQoq3P9b
bXRue1kSx0ON3G61hV9SpDXciw1rsdoSDdS4BvwUnEcEbdDF82kKOia3lKiWng3d
KZQChEkTxtnMwZ/E5LHAMrEdUBqxkVUu7zQFkwkPJ1/BwGIa60221zlAJyvM3Fax
zeoowblCu+13pgI8yixHefzhNyPRMKhT4Ucei5byp0PTb/0r7T1EBFPbEmtIWnFA
CQqsEW0L32cmc1u2uK0CbMo4UeOGCQKCcWis6NE/KANBf6S/57628q6DeZtVWyBO
slcZt/qNPMJNvmGuvB+he8JESQnwNOsf2SImnbSx7RCcGcTUEAw5TkLkZZ9L3XEW
xGxH5cJ86LcQhhQ+g6wNxGnw524e0xGkD/0C8Qf1WuxgYt/fR8LUmyc5efm2GVpB
hII91p8pIPfzvdekuKM9Xwd0t3WyZgyEQlqjZ9VqwFtTVsvgYKxKbhXdCrIJkQmi
i5Y7gWONtYbjK6HpBOoFG1kE9jkBMVWOSd8fbWcmYR5gUM732ZGmPWUlnDmE5E0f
f9RthuXVWCf5WkTN/UZLDKRu0/6LEuxAfZgKqq+sDyFKFQyYHZFbIkB0XLqejymC
Dz1KoW/cwjmURsSAlpIFSUcSIXFqZq3vVoBUCy3UPcBfQDDXIH4RPXYWuQVosbZe
gkp4AbD+UUuZAni3uMpxNnWVAK5muuwOSkKTF288mZRdNfzYzlGyGLLbAs/us7Wy
I0yEovVIoNASCDjITkUJ4SnTLBjF6rzltbSn4F/XgtPDr6tD54mbOs2VvJOgYS+O
DwpP81CDCiAk5rtT4OWJs4A2I8eCYWprS0X/4b01fYY=
`protect END_PROTECTED
