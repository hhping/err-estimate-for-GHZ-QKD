`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XT64HKFyyxxCglFH4ROwdjqWeosu8GTqPrA6vuIF9ozI42dno5THu4ft803xxeX
z2TKjmapnwq9+e+r4KVOHSixXB4az8kKbEyuDozExCyMlAlhXQ5/WZon0OlJEZiN
vSnmVPO80ZRE2+VQKksOJFucfZtYczopZLcCzeJDO+9q24xWrag+BEYGyMzsOeIT
twrrbkDCd7zwe0nbJhzVsUk/1ptenS+Hgkjexs2ywzU4/D226u8QtTtfDcBiiGpV
FKA+d56VRjWnbxsnrnpNhBoXdp5aeoj4s1VyBMS7zCdGn40WRVhQzKqe14ioxiyx
UPtf34X+mRLmdvIX0UW+xXCzcM1fyZ1AHoJYaeHUot72GzOZ1CvFdQhzDSQcws04
ICXAifvco5Y+6OgzLaJaucm5l6vVaR4Vi4OaUTpTeejDPwcz7pY6msbiVoMb/av9
5sWcJQhbJtaNpOkVt8dnEd8hdE8ipxHFZhmwEzv+G0wMcdBzUb84xQYPbsApzLHD
OkcQ/q9HyTnw1mFtS3Ju0v9SD9lO5djxENPIiJHlOaZXILs/Kc5bu/1bDlRWYoFV
Xgd9l27mUAyKLRf1QNypCI5feq0VMjXtWvZ4yU3yGDX02JGd+wife58WeumGwKOq
SheqrLTAp08r0lKHqBDo9aZAfB9W4EV0ZnnEOAvaFkyMY7ToUlG6pXzbPOMBHj9G
tCI309dE7GruK9Xt8MT8OnSXw8eB571yWQ2PLi5Bc8pDnSB4V9ca6vHc20y6B+FZ
NcUgDf87vMoPoscbBJOucXYgO1cT1PD2CDYhjnICS0T4oAJ8QFdLdEsMBYuzsoKf
nARxiduRPQDW23PaYE+U8jz65BKctqb3vCq3w8VeCAvGY+QrzP9/t+rEezMVlobn
+iEBrxiKDMNkOlFANfAoD+xXsp9ZeKcKR9pS8J9pOjAd2C4Cu9vvrWqHJsukdvw8
ULj77ZlHnC3cXQ3GJvaF7PjAcMwtCeIuBZ/V082tAGLKPQlzDKtSii45n2cg0rB1
y9xOyMq/uvtn+MaqX8xNgGlAY5ArYpOVSBfoUQVghT/IzV1brAQBWxttrvBhlF+R
1m6QodVCCoL3MdUBhZ4VlF+o1lDS4dNzqjxR5Si3aZJcCjIWfogifQGHYfeF3GK+
9OhvCu21pvuIhHz8CgwqhQ==
`protect END_PROTECTED
