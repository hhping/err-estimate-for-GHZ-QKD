`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6AXhLXYusNil9+Zijk5dCOTnuc4IuhdHiqiK1ToPYov6njVnoFkd9J1rSDGy4/sw
Nty/qP3dhGnc5RJeOSjYWs+ZXGTUkbVCZH0Z60k7jpuACPLVRKcOI4rJQdSw5aJE
mM8CImPemD3K2fvxj+sVeM1IbulsxcYaY65MRpTFTizxKpfPflZQL7doL4pB9Yfn
gSmVzb5dK8ZBFgY6t+JDqlEYNVXbJ/rpES5vsecNdtrf80c5xQGEUtoY+JjTZQDB
NvTHEFYn8TTTKdiErteya6flOlk+ynH3GlpQa/AHKvzIdYbR5f+nJzbW7mCY9J5F
SCvW2NBK2BNWCWftzQjkZrsDZ3pTUTgfVnkxCqeFw7ImgkIYhAR8dEEo+NL2MlnA
A9YiEybGWswgIH0yBlqFbh5dCwv99neYLS13meBKATxEuaxz1WYgFceRmF0RsP8F
B9zuL0+WRJvcwBT5G/C61gPysdSv+swgtqNZsQycI/7u+4Hbh84Q7jIRmNWSwEwC
qFiG8VGoXYkDkBGa/LPIy5gLsWXpaymGehxLsl6AZ4XsyvU3VmevpITyLJgDcU/5
Y+cHHkrwYfkhfkkBJ5JtkyMC1YAnRNbO6VsXzotVOhM09z2QPsXCg/dYCj4G0aCm
Y5BgbJibkfspkaESZjr8gcZ35UyMAO3DwZGsQh9sR7zr1ZikQtjAsX4qj8XoPge1
Yi0xIITZ38ZhitNmm+Ll/ioH2VNzdTxzhNhGOkTAUZg=
`protect END_PROTECTED
