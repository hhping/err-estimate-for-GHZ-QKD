`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LuXkLEM7WO8YkqLMNY5afPcSKqJcZ8Fdrjuuv2ghJL9tLu4TdCQlJdEDRbRDaGJd
pmPuTf3n03ooEt38/lBuJiTIJ+DTaPvzUPmLGfN6quRERNTjreABr1fKLHRkYFVA
ENFz0djKi+vOLyWyqMknEIKDQcDOlb4g8rQBTrep9LvIvAaqczPp2U/Xa/A8rExL
M6wW8U9OV2FhpbbzcnoBH2nek6xJhAAWCi0vrzQ/3Ll52+f7QnwmR49QzNMrnFLO
0+cE94MGpisHEeF1KGPjsKC3L6jRX2pkBJMwM62j66TYjLaRviDHSecbLq+CFjhq
96LE6F78XmBuf0VupOIuwe9o1JAIQvRp3g69TLgHRsa4JqfLpjtFBevTMiihNfSV
Y4oCH52AGEU4iOBw7gUFUi9wOQ38qBNCCbh4g71Ew6gMUsyuIaS+EQjbUUbgkiAe
BdNx1tt4C3JXWXboZODCn9eOoUr/4ynsWwbkzlE00iPs/6n33VhZOgZAr3swiZfr
lUmeFqzh4QWLCo36XQxeNKDiaO1padKtlBJZyX13Uw13AzsZcToeANtUR3Blg2rX
3EEQGyu4DNM3ZHoxBkO77jtNSiyd6sjuuvZpLpuma2PsFU1P7vj9i+ZohIgMppBp
gZK9BHDCg6boUWjH5sr7hN6SMVC5K+hndpuSTI7XCdOQpN3zbsi4COfjhCvtfx/R
GMcGAAGCRudkXEL2lONXzXsmiiqgHH5/kYlgAqJr+iK+1RovxbIU1RgRFYH+1doH
TJIH3Dg/gf1Mc0o/d3Z3xs0CmctjbzawTkTkHo8tdhro+Iiz4iBHu7M6AiW9GXM+
5mP2WN6A1/NyjaDPCZ6Py4CF90dp2fGoIkYsKlcUXFhF6Mw2oEjQz/5MNV8DXzLB
heO4IAnxtjWJ43Vnkr68GJJJoVn56TKDjBQLIOJGAmZSebFm93B03UeLFX+ZRGqO
Ems4Agk/n/kGcmbibZL/QOq2qCVtX5pu8ktx6nZLuB8kcwTlIlGXgafTL6U8u3AA
IpAiv3+kFEeHnZmmQWR5PQFOmm8UzQGEurlVKqCyLltuSkeMX3RkJpqbUiayi1o8
RfCk1tF81gHHFdrTHYAJ9g0ZQnz/80GGZ0qqC9s6smGIq/s3DDFxd/2lxylH9eM5
sr43QCS0GgBrHm48SAu+Iw1123aJ86xrbY3LU3K79HJqEtN30v1SLz5X3LEEFmGG
gcOrG+7IgpZJyYoADYC5uIbRdDVbr70nsThFG5XkZXKR6XpNAvd/0/KLMKXhxlqB
nwu8KSm/pJil5sWMVbMgCFrbOk2Gfx/j3OoR1NCh+3gx8duyT0ED18FLZJaqYUbr
wXyHjXT0Aav9aD0HyW8b+Sf4pHkVLhEP3x1w9HPJ9XCqLrOoj978JcRxeC8LjjRK
JCiB2NkcOAHT7LcpfZVJtkfLCIbpd0kwhbOCqzrXwhAXHzKfqahK00CxyNwKrAZW
2ihJ9c9vUIXqVnLQV6sR+AlpFrIyv8Vx/xhCIqyUduVeiv809xrV1K219h0rXOJb
gsKY+4XUs+NZzCDRrHxpEJW3WK+pRPXQm9C+2xDdKKe0yT7KrR/UVAp0Eynw03hl
F2+E+1ylfkzaOk0J7k/ZxKZp01k0TborvrzfPXR+Oe+NnrOmZ2hdujNc+IJtL4Tp
JBy2PWcSyVY1kWi0QmaFw7Y+WJSIteRahgwhTU5guuw=
`protect END_PROTECTED
