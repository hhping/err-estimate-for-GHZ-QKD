`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMsh3JxP0v3L3Dw9K9n6ckbqdaZ4ArfdYEai1jSsbD77VhdgJLsCQSFn+viVsSXh
EKo/W+HLfjrUj4FP01/BYJPDOVGYizgbd2+wwFNKTOn9GqdYgvfZZKMYIIF9elfe
aPGQ/VnptyTtyFVHS5H61oGBAqXGTVCrGW5bPcTyIDX2SAVoO8Pol0r+KIQv4+xW
dqUhyKHlZiuYBJQTgd3lL1TGASS3HUNWoOkcEPjVnLdZQXpjM+yCyH8QXyr89gBc
Y7KbHknUjmvudZ+5Xf1vFLRhTT/aYeBiaMrP+BXCDLk49wyKbse0lOZxn2CWJGXM
opYzmKqeBropSH1U8DJDqjqwv+HUa3e27HDKgAMpBYRV0Z1eikC4oQkcdSS3NI3/
7KmDVDEvZLYvoCMPibml1jYaZm68qbedz4EF8grepSw=
`protect END_PROTECTED
