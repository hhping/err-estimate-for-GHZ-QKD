`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6cCkr5drMJ3eiLdIyj00gbIpag9MGuao33iYcCbjl7BBhSoHBktHYUL3O+YruQI
rbN+VfnP7ZesIcuqWF8tWlnpp3/+t2fVGvw6suPS/NNzCeWxvZjN+ZXBKvWpSZQz
omi8jE7Ws1jmhLfAuMVZv147MdS5SvVI/wIAhhAWzXf/N7scuahgCTrzfyAUfheI
Bqu59kT4zG0nqXnlN8RXleUHCrr5zJHjo6WIxGsBxSJukpGrZX+/o4HBx9apvut6
t+qNw6dTPic1hlK1ZVZwUVcDtLxiE8Go8kdA4svGL0Jxr6xZGuUGPRGBs2aKS5c0
h+iR2+ITqvy1YtubgLSgnopUSusNYxDQJSPX3JP8nBFDwsfdJ9kwsBMQ2Zkssr6w
mRwaVGE/h9HkZr1N5I/2Jot2MddPjj6LhM7eNKxwmP0iYRroA+J1jiucqZxTARlK
Ge4aCAtTpKvPi59QOnxQBXw5qONXLOSLj5CS79kzb8ts6KqXThWy9IsNp08d23qW
fb4uyGxhgpIB+Nn4ZFZrKmg63V244ZbW7z4F38yv2NHWpEwwtBbnryWE3nTLLxlK
KmHRwCYDtUIdAkuCdUODilEb6R/4vPNMoOqqIOpEJG8jcxvA2fuoESV0x/NlyNOq
yLJPEthvA0naFdaBL5VUhXnqNpJSHigX+gC6zhIRitw=
`protect END_PROTECTED
