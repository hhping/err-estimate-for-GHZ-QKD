`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/60/243AsXQs3hyAlEXwXWMaIOKDVvpZWadUd53Fko1P1IBp9UwHVWa0g3YSbIZ9
CTPUi4TgftWo++YLdTtedf+VaN9/UbJycrYO1A8hWnh3jDK6Avx2pi/gQZjYBgin
5ln5nl/iZUM7zZuXR3qnN9T6rSx+fwnNVksJJbifFPP8az9Qyn8qC4pysGtY/AgA
Y4fPfIol5mxtDsPQC9gDayWd3L8s8sCEFFAypQPkKfBKQOqZCmWqV8EaAKgfQB9h
5s4xgPS+IzngYGL0S56yFCKKe8KSp80evE+liNf9zlye2LkSejXg9BY4dYlr6QFs
w3srnvA8dghoTB5C931VmrI9fKMEYMHyR+c8ZzCGJjH9NKY4nkGvX3Ln1Tpf0GFI
tQimzGFOwV4xQWF7L3TM6Jk5wVMyFzLSRP6+wCKRfZKFJPg8rinkIPJkPuOBxkvE
poT5iqRUH9aNkufXntDkU8QqgMyonVH6QLKvilzwR4lrKn8NzEWWqVjMP/qSs3P/
qeAsbJB9HEJTmqtDyM6MxUEzr1zq6LvYQz/d9L6wYKaAhA8t1ZMB8QHfxtthP1+u
o+gGJrQYax6s2e+nSHGefuFgLagD3rQRAahY/OXmzyqCm0fuLE9giiP9j4aIOq+I
`protect END_PROTECTED
