`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xp22Kgvo7a/6OBb3ImrSR4flegrMOJ0SyGiAhbshsA0NCNL5YLWzrW5YS3ci4K2W
BuxPT+pYTmp7p1kAv1EXE+pgoqLWNvUMvowMDwYjmF/VlsUCApmAxxjy+/2L+PsF
tm4vx/iA6B97hhEppy7XWoMu95qTW9OXeFlr20KcjltE3hgTCFSxle4BiojITX8M
asTGHvsL+8V3x6ZjP0VtokAVwXE5QyePzTfmjlRRRh0D0lHf4v4DwyUOVMRasUf6
WE6tbbub7xh+BwU5wT7I9SJtKVIFIJnO6aBvT8IQs2jGIyBkHNlTL4kWCQ1qxx5X
pSmBptzDdYmpaQEWAxmAcR+GtMRUxpOhWyUlLkpcFbuGJIteOAlWU9YXhljlaZGG
AGWOq1l5WUf158mmi3jsJ/2XaZCnVCfYutgsOzT4zd+jIt0gKXj54rnYOdVEiMom
pKg1Q3aukDJwHe0/1VkLhOu84ZnfDzdcwRi4pDmo7JaHbe88YMggI+dq+CQnomYY
pfVc61+U15KLJXRwZ++EWjkoWDzuVq1Rhl9vuAEk72lTc/9A82MQFBBoOHiEMxBt
o/AsMjuypErrdj9iSzLXHOOIZOxACLfCcwEnC4snZfRyIObS4CtYKNSpHFn42vq2
Il0Kq5MKlcdgCHNkyC4HcdpESZCDy0cz4tRo6FX/ehSa6gfqkX+o5yxL5PE6bH3a
4IpfcyEaWJ/g/cK29M5anUuCdGAf3E5iG1mzRsFiAWhh2n/F3BeE/iSLRj2fF914
gRWVQtdv5mV4+yhG64e0NSlHEotTc3RRDZMfWMJtv4++Xh81C5TbZV8ykvxTVmKw
Z1KPopyxhJxPUU0MGWMycw/5CQ05qVEosymHgXFeqayWVIecLS6plpge4XLH6vQ0
ZAE7UcgWSUDeJCNXcss4dCs18HC8Q3Qwx+vFL0vG4fVje/CBGXQ5YY3WDLc7jCol
ux3QdaGZHcyeKHaFCicuu6rPJOJTczU8cHfCGv919rB9QDf2U3Fj9UsM1veNohe3
smwDtnkIVdOYNZTpPf4X5ZbBCv3PVpv7X31/xOTv4WuHk+25lmfgvZv0AoGaRNOa
veahPWVX7DpoI05BwKbQXLarAK5UdJaUGzxwUHivqRJOp0IjqEa0ArK8jWKrfYYD
+SAppDNKFtnRiejbtdcEWh/kcfY3DOiBZe4CWjosjAVPdOdmtxidpSs3g5xoLCQf
KDrMUmHPmFZb+i5zTFCwtWZERvNOUTbT372xmjsI2ZCD37W/1LlSLBWrIG6kIh/h
rkbMaV9mPSX3XfX+u8MrRZzee2VQR0ISxeQDTKvrYqiEbhHMpkifEbEvsddx472O
1OSFcXrZB/oeLY6AAm7gZvc4TPHOqXMCvNn716DviEqxJO4gGrOuAdDZUo4zHTo7
Ni6Vt7/XQP4cjbZXzlaA6Gweo/CsZGWrfThwM9YbqmY455kWBgmeEcS9k34PRKyI
hxKDhwcjCn3EZxhU2lz8mc31MZytsQQ9T41zeCpd9aLIgzFbf1LrGdGpKWbGZLZH
oXQfYyEgtMnSdlyajzz7P/zykcEhixzsYztY8iGP4vM0lrGy8jDijZx9HBBoS2FZ
1hVuqb1kz5uV40ngi7b+5QfNsJSoooZ36YsLdl4IEeQbBJ+RzpqkxzSbhG+TwWVW
Ktex1I2YrwgochLa7RVwKwhejl3fnCLxqjeLXa03RbmudIw28D7VbU8TZtCqsm5Y
iU5BA3n3YICSzdF4lrLtyZ3dJDHVlnWr/tYEUbGXH9wWOYFfqpvVz9DCIWU99E84
dnJhRJxe6/HqODWg6Vbvh0wWy0ySetJEXNT8gVCnKrvYmlyBcfr1H1kl/fj9SlY0
i0Kv2h5h+xKhNKuAwmALudk8UOsjKoZVW/MH+C96SCOFsJXRGjfQ6Fm2QL3El0gJ
FAZ8ot41h3wIdhKEOAqZ0tZ42IHA55CdypvhRrtBcjvT6R5pkDkR/TVdaLM8kk/M
r6cH4U8nYVPVtBKILTXYCWxvVowfpy50ldq7fUBtZwYO9MCo63Oo+bA3P10u+CaC
Hy90gPjhbhetSGTOoZJ1Lm3KwWJdiW9VOcomI+Jik5aCt5gjO6qF+VM9zAFN+U1N
PqW0zQeA5YFfHZpG7jjRrf68kne5KcRXFttWZRaZ6E94YOKdTCIEzoD0fIRsyDsG
HwBnBfmSb3EfW4JFXpIZHO1A4w0E7597MjfhF5MBgYD8tUQcIhDnnZRx5tUtJjri
xln5YkkZsTCKBduRRmb8uwcH0UvaZlKSCIJB1gsoKmAfXzYnMVtAlTKk+Spfd2kY
15I2VaT6y3obF9Fq9rRPCCBFfq/sOovAjBcvf/l2Dr+jmH6dnKMflgJLZv8YVlVV
T0awBIglzOmnfyNH44iPvPPAHP8rhmtT6hG5AgUnWWl6pzfjqJFV5W9jf9Af4dg8
yCmETetOt5vhzYGVnlLL1y8fa4AA4IfRph/Iwm0lW85hHlYw1OAcHJ1b+i1ptRTS
GLMd2G/wa2Kkp6VVHJmCyRDyHMudoN9uV0xPV//aNnW3fmL3wvqNarJgox7G55fS
RUO1he19oLyqaQ1tk39khDy7+0316deIEEsepvEd8AJXbtarly0qCanXzxru8Avh
OGQvMQZcfn6pqcUUsCtgJKnHkE/WDozKw9k5kHqS3m3TeWt71aXz7Gn04vRi/8yw
mAxKBnb8H6WBD5sBZd1AVw2mAuQyvlCw2FI8x/DylIEwB/gIpfff67Z/9XQxaeqk
0nMPOI36utZJgCQhyBfLxWU46tqvM7qezqIn0zDZNT64mmr/0pb6yJUJmB3b4kcU
+alOsX0nK6OKzTbwMTBF7/5o+C8n2uVmcrzag+cd+2vT7RNcVZsnOIW6FsvqeBMU
TojbatNLkjS3lRKu3RTFAvm3hOff9X9yFLyZTc+Jntqr80VY4xM6J+6EzORLnIJh
eg0y5m667mbVn5uoP4LQ2m5ebUTvB9U720q5LpJ1xpQ8gSLynHNpGye7e6XlnitE
E00A/KKIed5qmjvpA6GLBHpy6JwSXXRLomdKYWabHd+mPG/93BhrmHmzXUorV9R3
PmR3F7wdxyRE5Vq5Jpazg8j7O6r8U+xhLfTomid9CK0nN3a8JEwT5j6q3/61tdoJ
vP6HebrjwaXcz9nNIPfcoVff0ZUjc0PmIdZbamkTFVvcSkwv52muQZUbQ/18y26C
ugHOw2AqWapGHyLid3mg9kmndOLtFC5RAE88zIDrt1Qq+o8l6haZB+TAH8mGbvMp
/oya2+iSkJTOk9gziEIuxvz8WRcd0CSDFpz8vki+CbCtdjb89eE7TSzqnMhm/WRX
rPm8Px4oxfRpu9Fiwg/aLN47OVSEp9GdohSlLzQP8Lb7jvQSiEuwZmJghzcArnWq
iRATqj5A3z/HHja2UTU4sGLWhlOlZYsGSmx2So5RnxvRMhH6f4DfI4WyVT3N41ba
mOY3b+Ua43oQbRsDDdHCCaB4piGFkEOYfLCw6ZvLBMFvrxUwK7xRqKRYKtgCSM3T
RE2bDt+6PorZqQL1+MqMVq4Kjqo+tiPKtpUTLEY/uHBCMFruqA9NiWGINdR0Yp1E
GIVYfQT184FSAhVV8OkUJ4piUh/DuA1zI4R8jTUBCOX+KAZhM2ynST4qMM/IaHn2
xqHR3MAuT+0Safweg7QchHnxbXgi4rgd90Asbox/I+dXeUmtQHG48KO4Oqp1HfE3
n97nop8gAAq49jxocjhtQpLW6uU5jJYdRg96LtSkimh3HicsCpml3pkXAC+tPUgX
Qr0xYUHf1dx0nwNRUnzIt/U9uUbApz3vLhnIHN3srm3HtWAxr8w1GPQ9ih6E2u0h
WbGw0D4ept+vuPxcP8ndii3tWRQ9TMiPc/4pPN1Tx6yA1uP5YxIp8s9eLyAaNqWM
nYRmEARHdMOTu6ThtxkYPV0ER8LrNmuZlzmUIMrZcbL9fVYSmA3YJYbB4NGqnOOP
Z2RvNjrq1iAkfT/iaD62P4rEm5n+nGMkpWgUxTbVgD//rT78aC+KENls7MR9TOsl
p9eAaydDWqk0kcwLmCElktGh49GOELxrRLI18wzrsBif/8xEJhK8k7lzpL+17YR9
fFh/0AQdf11c8cX5yJrtMP3Y4Xy5+pw+SQgzstB3hKl12Y4EFPXePts18ogR2esQ
X5Ip20m0NAUXjpBz9LfTzuaLz/qZ46Y5ra1WjPfFnBrdps4HgfZVuk0NAVZjofRa
IztMvuuRdhpY4rxAQ1kIaAMolRzET1rii/ZjeW78fGU/wWruzMQGqBOLlvyaiPBp
Rl2BdLBs6k8RvCiv9ci/T1Zunwcz1qrxJ6C/ukK9qkxxji/00yCa6jWLg2739zDk
04mhUXBlxDE6kNjzWj/7T5XjIWwkuHZdqzckSQL8loS2XXOCen3Jvevd7dsAvAuf
JiUFEEElJSGmT8cUXHUZJTff7F7P4X5cAEDbwfEUqUVR0q5Q5Ce5VjLHgeqnYZdR
tumRSVZpFWUTcJ+H535e6C3DkP8mQM5aSR7wO6Dzvm4uj4PUVVQYZKgontddehC4
qg08a88jaxY89h0GHv6LtJoMtMTTk/72k6cj3o7c8cNL6u+o593wbx1vQzqneRMq
Zwog0Wro748SE1+LkzaOchBFcV+YQ9ZnoASLtqUmMkMvSptC5pkA/PWKNrUG4Pab
5iNYsPoWxHCoae4iLCkk07vWUEzYDIV2XlVBJJl5vI9PPA4B8tf56HzebzybpDIJ
Gx8Hqt3vt+/GkX0BY+GMS0owbw6S/+avdtEKolLTYiv42K2KDC4SnLkYiCWcgGPL
TNVeFatRb37sBhE6M/a6yfhyvlAhbA/EGhJAAZQZcQ6o8ZX1yW5WlDcQWWEy59k0
LbaD0xdcu6u7JgfiZcwWIWN5eg3P5lLGIhE+4R3MBKIuuzVRV78MyV7XsjsjcfQj
I13FgtqyULywxvH41YOeBq/HO+MeGsKxAm4ZxMGAo7VOo5AzgnsyMol9GmwPFvcT
F4S1sdb8R00SDrxtA6SoWIEQ1ENrzoQHojzl7ABgt9Tv4EXl7R0llCZ6eE7HPNuw
YSXsQ+ggVPwQ1MmL+F7lBmBMl3robn79Dc1LP2r1zOdfxIfHWIap8Bw4vbfz4GnG
jbybWliK34a8YU+Fgtb8FxOvzB7ef4Zoc5Ys92yyCCSdHhFxy9tuZ88HPX6F8+zw
l6ujkjMK8ySXCf7t8f1OKZgGIxD2ToWwj6wi1+6xJsiV2CRIKlaiQ/jTMkLuRSDT
2MA/F5oN2JsRTHFTPHHhQsGGX7vnTBWbsLc5vumIn/fyiMqJEPcvjlkuoxcjH2U1
C12rcTSD+CMZuKFDTR5gKBP1sNaIZuP/gKPGoTyI4X6bQK7xnqNuxs/5Zex5M9g2
302EVMdQgQ+PRawuEO6EWuW0hge2U+XkomCQ4N87L3fLFRWY7ekAJQA2FgvRihtn
sdpW/tIp8E7/iMngioT+z8mYHPk9JnJwIkDTNtPQtWiNK+NgcDa4ECLNSbygQT7s
TBAR0JyKwoFsY/1mBzwR+5Jd35nQmAa+HL0GITmVa6AD7sE+UeFQHFvZcI8M/taH
JzrKZNZSFzFDqzfWxo29xNU1nYt1pJPXSj6kE81Br7Snt52+KdY10tfoQHZM/0ni
diLA9Yfrz19GayKM7uRF0+Fk4BQ204X38xzqX+XdKEmeSTb6e+4mFgDuUctHgGcQ
WrR298jKNT9CN1wD6gTqe7TDNt0N+uSS74xjzXsimJYMtf9J4O9Htd6ywRP/Z0oB
JohHRuk935ZpdzQAudCkMW2b/ouIxXDOKTay+cbgN6vjvch54YEdUOC75jSZwFWD
EAH9DogBrUWdGIuswYPkDuvKvN/rzkOT3k1c2ESgvfelEBsHqRq61P/MN8g/IFT9
cSX2BPNPrO+TMntkJH7FNjSf2hvWxC6ED0yHI11CCLXd2eaChk6vM951uPYQaXYa
ybv0MfHr2QYBUjzkziKqP4WBvUUeKV5EDSjprQaD5VUQGVeI3Nnfw2KN3vMtmreG
2VHLknn1NE9JXg7CZG2fwoBHBph3fkej5Rv37aKS0DfQAfiKYmRhRBskn+wNY6Bc
MTw6IDh0XIvGOFdiL51YKU63wPYJhfuejuKSDnX1y0OSTG5qGKa7Aphy5dNnd7/r
yL3B/vzYQDN1S8EnHVVoqqNfwD+u2aX5dVWgKpJVATFyQeZkvee9ayIMjxpFycdQ
zry01GEnznauePjMhD+cri9RiSoAokWvvbuqWsVSlvVpS8+b0Xm7cVtDcBMJkOPn
VFL8aeRD69nxXVyvZhc92bKFus/54rP1m/7p+NCePRViCPOYSIWwtxnkedG95v+A
+FjS/txOZ4JlYX6iq1CoQfwtL/Tk/fNbrSLvHyxnXfWclHUwg6McZ+bnAumD2vtZ
Mb3fAIAtJEAMKrBEVDEYPwWmjnDQqixhOR8pqReGZyEj9GAWSN2WFnwgRy2RcXsC
QR25rGbZIB/9OHj+RPTO2Q==
`protect END_PROTECTED
