`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p7RayeZFR0z0Rnw+42OF0P004EojE53HcPqlVmvUqL/8g8TXb6UE8kBul9Y7Zrol
YSvY9Q8NBcoEa9IQDu1DdcEljtz/gjyBw4XZR2Z6g57j1jtWFy1WPTCsKShbDYXg
iln/w1aFSRmd/D6M11i8zEBmHZKjnNovyKoLmSTg8SbxTRyIhNnI3K8uR+ED302U
eC2rPQRtDX3Gv/j1MQeHgEhqnhygr3dDSGlE+dJw6TxauCBEdZQ39xk+BCF9D97x
DqTzXA+GZQ3+vpvQFBbgXSJFAXaAnAnJaYISxmF3cnQ6G24yX6jTeiFZtnApuaFs
tbzz1+H24aVvK+U8dn5wmv1xXpVujEDw3W2F0ssRSy5b6v139Bq8wlalPJuPCp88
NqavttQFgefW++b+qO0lH5L5zh8WefmOaPorcNyqbTIga75zr/ZS9rGPkwSmu/oB
TiSHKmj8CV3K8sgpxPX6AFROvoFWxFvyBc/lUKqsfCza6eBbASGXuUXc97xRhKt5
yuuKZdumdE27HV/6sMJChc0zA6HfISPHaOZEp75JzqvRWJ6lClzhjplvhedY3Gtj
AAHiBf5POdC71La+Lc03z5kGNfljAX4LqJKA91yQoDxgwGJ79PPqMQm9VigZMIkr
tQOJmJnq+i1Hpvot6a6FyZO9fdpp3RPFoTlBsvH5wBA=
`protect END_PROTECTED
