`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rxzi2Foj07PXSoKk7zFr1D8RCS4GXlLr0+jQ0dT6nPAQeOiADYMz4etgXmtnxCYX
y/aUHjOVbTeatoEnEdOFlhWrC7SrL19+iBGopq05SoZ7DCN2xaFlvFCU/kyzhBSW
uh2u9FNHjQHKssKWqTC2vr166yxa47Aqi2NAUk3o1Y4VQYXe0g9klwxT/qmtV8gU
YX2ngf/CVjaaWYykD+LUsyqpEOiJ1tuFcN+jVm+Y9FjhIFDUn15/KEcC5O1ppwXT
jsK5GuxMyxwAwCDNdnAoteyqTg9ifU6nJmYIsQdrcDtudF84/Gbx2IvQDG6Y0k1F
akEZV2IgkDcOKxMeu/5SGQcKhsN+AvyMTmW1RxJOE1bdEg2sW/HYRaxOm1od2VnR
/XILcBXdXsxHYEo7nJm/xjqhKxW9e8NRlR+HEo85bySBsTsUygMfbRBw7VQHP5U7
ej8pUgf8cDvKQIffwbugrAPhj6uWyR6mPZv64Kd4O5OZG1RMM38wTLRWyopVQxLH
dsut8owHDt8Oqw0F0mMDhf40RKbMNepJSc6Sy3HSGEANhFFKkM5k4AbZCkFVSlI3
hj2QnXNNy5EVVB0cSc6Dpm042udyMEWWRrUcw2NV+k1ri7LPl8qPyyc20fXcKbEs
sdnCHBb6wlUCoBCT8cbL0ZVvTJeQhBPEazATzKcJjpXHcEjg5hTi5zEA1fiS/kf7
EaXwAjWZK4qW2WycBRCdQp6J5CBk/eUszi7lJAQbU2EoGlzcaoAWG7Su6t916Eem
DIEnz3n5RxCzNtA6unDciRxXmWa1lW3vnbXsWC0yVOYLjlHtm2+jrQ5HIVALD6Ph
UjM6ENsuUGsTm/BhvFUn4TC4Zq7zWKpda6bkuRObS6h2aJWTl5enRF8XgNILEWBJ
g2uP9M4VZ6+EMqgplpWOIzD0ilqtN47Bd3NSQYkB/aqqubhi8+utIgWgWPKKsg/4
nld2ClWG071pRIIyHxqphA2uSMi7QJDPzTKPGWfx2FjSRPEyyQKWrV97OZWjDJns
/H3DIpblJYP6i2AxvdmWF+Vu8n6BFv3tAEfye6FZWzQbPyHgIzTH+Qky+LpahULv
lRUONVw5fLhihNv2CdH0Z34NxP4mi/+mRnHVmRQl71+PrbSjczEs+46bHNDbYnxX
NYe/7Za1N4w2OdgDHLPgZTMI+jrMa0IXMAuCyUC5uRPmjKMzIturk2tywecNmfwv
jRChm47Si0HFR3kBwJ5rPXgiqGmSRPIsoxCjtkb8FYmkDAyiB7HJldBJs9Sw9BB0
poX+IeyEDJDdhtY0xlF8T1O9VfQqwRlah8ObYcK4q+s2JRwlPIk7kV960h+DlahH
ldEKdRRrZ3B1D5A1GWzrCoRAu7GR3akSpMk5kPnzrA/moPiVqww25+TXv+EWHtYc
AAmm/Cl1Kjkl/sLmMj/Gnalab5LPleWmsWmH7qLiiJSj5UTzgLIxxd8YJI/Ew9kZ
mDBBsmjBaDmq0JMGHpv3+398YNPN7oFgqMuIDltd5beV1antVksugjUeC6ha9Us2
LAZnbtxdBH9iPl9vPQMjqK+wkAEgJ7lsXFuxWiUHDCXgl0Rv3dB56wb2kzr/lYWs
/SRUe9fluH7BcmufiGt1OJDxFI2/XWLswyFnO+bXJ8zirfzsT/mFzlM5u3oqiKY9
ontoYmCMADZnlCG9hXDL2SEkJ7tJlf4w+WfzwQQMoL5OsPQhkIKY/LuAxI3JJoWx
xswJU+ZE2zk3qMXyu2Flk/or5kaXLqoWYltHfSZuVdZr5D7MQmyPkezBEneoIt8S
eGq3jMhmt9316TEPpSyBiQ2Iwq8avkbeqO/ZUbdoPu9TK12BpsSkd0Yp3cnaL6Pn
5c2t/hFFJdWAmxQDfbMcqYghUBlbh9HGXOi8CndkePzxDssLDhzZJjkMR8U6xokd
dfiCs5hevsa3WE8raOuXYHLgULtH8BCurXNwp+9BQbNbcGeUbGvDkiUqFleRMp8j
LnWBtrdY+9W6w++sKxu3hfMZu0RtBwdHV7Jj4WVulw3V2TRPpk9mpQqU9LCC0QG2
5/7juHDN0VFw7Djo4wYmbZWbdimv3+RCXSR3e2u+/IKfohEoxJYvjnQ8vVn0xTZz
3vBxDABlFPZ+xkZNN+ekBMb84ZZ5mKXLkbhNtmap3DF+Yw8o1n9ek9KOTxHBDJH6
s39oSQYUON1bGZhGfdYgfB6lG/j1eoysHbedvBaRQc11tIdoYDebDOcALMqJAaBS
i4f5lqSnTh+DItcO94/Jo2kRwxVZdXIe3FoawB6D/bH9Gk0oXQdyQFJgiroiiKUY
F+LdeJ+RMFTZuORiQzzgJiJfL0N/lyxnL8zvCd3WUYg/+Gr5Xk0IJOtVsGlcnkKQ
4ya8OOx/aQLqjANyFD5olET/Zbip7BMnNSiH+qK2WvxqdCBPkmAARlY4lEdiJvY9
Svmpbu15FUZq1Nqrmcoa4jUDRdkM62b8wuDbiKQCp0t3beyTBL/dzRuc5AeZGdbs
vt0cJWjwfr4PGUZmudrPn9+/8CWfmMr6zeN7+UUE1fwwsk3w6NApQ+gKwN22+ROW
X0suYMQrt4Uf1n4iEVOY41/XWZAfWSY1PL1dcJtupVhgLthjgj1K/QxBNZ1UXEFg
Y5iFAIhN7xCHnfRPE5K98ZKc9X9Ig+s41TnpkgBuFc8Ngx0fBrCzHwYgOVq4KGgm
NAC7PnPN8/JErJlpZdTwsumr66/vuNo4y+F5uo0Y8aoryAfzCgKeNdMykz+YVg3D
7OO8a5+kKnkSMJBO1sy8ExjRByig537E/NRzZ2fujlDE6DvEldSpQwxjmS1yUxyv
zBTLabmyyPmZFSVM6+cR5ixosdMvLiJOl4Fs40+s7TemrbwLgZJc4lijpDswU8xS
OFon6MoaR9HrluIyNmkuDIEjtIBxORf7ktgtgB4IFd6nIq8QyHizU6U6MYfSCCrm
HeGgwtlwJm8S//sA5jlf1+P1FtCsZ6gyzXdF4L6/Abodo9HDJ9yI1m3WRX3UeTEp
uXR5xphG05+51F+vavrgEXA6cHOPv9zbfxtEpY9KUwAKH+YLR+UdZVyLJx0ifetN
Yx7+8RmC9P0XbeLblXwP6F6mO4LRxu7umgBTGJZRkvC9cpiQzytmUC6CmUaWzowJ
i0ysdeXUQ35niB6/KqA+z1CNrWfbuS3yMNy0lDBwOJ5e1RA8zvP/6yHi6hgu3U3W
wSm9HAA+PkXa4MGUmjt7GqnKuCXudkyczSXjKgKWT4NanP9/2dhIlQzj/KJJDasZ
mm8Qbso1u/TYYqxHf0hOgbLICqApGrpctCkrHwYSiLkbgbjWTyivvy+TrGv1k6Lt
IFTzJ+kv7EulFlK6Vqb8rMNxSSx9fMD75MBDKuIUMCRW0b3g5QHz/nIlhqdsL1fl
9lwsdzhbumrQlKMYDS8IN5LYXBv6gxPNgjtBneKg3+mMNQJVbgF+ZzzvZVmqPwwN
pwwPINOgKk45gIyBZLye9itJ4b79IXy7k8ov5EFxMPiTzSQJEp0ncVBFA4j/MmVM
t/QW1+BeeKnHdHPu3LVSDwj1lnLNCRBKErvCFoYa9sibh1jp0k0uCnDeDAcTKCD+
H3MlVhCzI1kMM2H8hYwuc4DDqH6NMzRkdFbMkTgO1yw5D5nEJT1Tixc9HTQnxOpt
I1WVCqsjNselRMtw6QRxWLtriSTofuo0wFxI6P82olNCBCNHScO8Oi1TqKSTUsf+
cZJW5agLcrL1cRldBRgDOrtZVAMgCCgZEpaIdm2/sF1SbSqcsMhrO44SzfwzhbRb
kAGDe/PI05CbnwWpd0raQ+7TYL0HnfFifNLiMAVwHwgj+pXMpK5rGiMV4Fh3+9SN
+UzenYYdLWKvtzW6VtVvfgm5RRzxoDB2IvDnr7290c+FA4/8ZRbDq48fLIaFJiz5
kDNmWRC9fzYJT9QFXlr6ZmDNHAaDTTXNyA2dB3/VpausvIFHNbDMKsuRQ/2Q6j4X
t5+3idaEzhK6GXCZ4j9RXudWT8tg1ctGJdz8/TDueNjIE+0UUGRXtuNgP5zMVFoQ
0JlFlrvhEJbtG9dEqe+k80crxGyJNCZAOiLeqajqVGd2tYyBIdtKuOYTTYrNDdG/
5xlm0VKIOt/S1erjx1ewaby7njI2qtF2uKJv2LdPl5HZWnbl/sBH9bZZuoQKV74O
7SYCAyvX5CbNEPLvu60T2nWURWIDN4dXuJ7mvkTBxouomcQANwVDMkvogIWSg5R1
TLhVwZQgS+crhpzdnESZYQ7KuMHB9t/6xVcq6wxpxsPIRuFx4hqpmLehPSxxUm24
M3HPJ56VkV2PVPxzZun4MMRquh4Nw9ELVQSGDutFuTr9/M6n3fb+Py1yyKqyEm/+
sQ/4OCGQAEuheBvEBRZGW+O6bIHjdu+7096B7pG3+QRLCXPogdrKcHZXlC8ZQS8G
m4a5Z+6aeuGqxWZ1AoGlDfyukIqs15w485cPG6SIUnsLpq90IhCjZ+xXFH8FPK2O
vQSVBidolHkK6bLYgL/3Ju3vARIZ+WzWTWkjzgp7EvwrT0PX/KyP3cjw0aeY1cdz
XZm/r1CxeDd++Dp3B1OZ8ZGCgSwhw6fZGtiEvZL2rKpqbLUh2UWzvPHPnnBFwBdj
0itKe49k9lljT024bY19I/00tYOHfq4qRgSOXax4rhKkGJivK0mbFF31yyvsuALi
sMgMxNIEvzQ1tsX8b1STbqqVTne2i4GHA+HXo7laQgbgZfMnyvQhENpxpa2SuoMB
woDczJlV8A+J+Hy/xMiK5bYWWTQrQAMpBiA95erfBcFHLjoQh4XHiODcByMLKY3K
zDQb4qDE8Myx0pW12lbjGIScHoN9fXSQKWxTaI3e1ENazkssa3EsZJS/xkgzC6yP
UOhzMiGVrFsZCJY5n2Ya2CX5VT6cYvMWBdIN5GgUWAL9GGSDjGLZ9m2iDwzML7Nt
2gVdYHW9k61lPLGsjeZ7NKpnHAbTzrYr+fRXCPDGZTtpGD8wUGoKwJ7WRRIjNoa3
nY3rZqhH0Xsna6mSxdnLdD/hE/k4WY7Z7kYqSGl5t1qQduRJCkzdbBbGGuhh702v
V/ej06uTGHCxcxoySMjvxqjdCOspnJrV+15usgTmWxrD4snhf66pgLQ5kcrvHVKc
jHQWFmmp4CTUt04i+ZzECaW4qA6k81u2aSWyX0Jk30lGq2BYyv/eIURzPwDC7Z0j
orWu3ST6cHGekDulKQ8DXFC4f77/DHEYUQQtO+GI1awzeSnn8xoaSHEARL4FddcZ
wLYzjyzPYU3SvP4cKfvPX9AtQmJ/ZItTNtamVxsM04vEU7QBMxh9k9qCbWri9V7b
WNRp1bjhsC2z2kHRJc6Qx83QcGeHyJFtsbiF0vYuipiNFgqxEXjy5wcEyqCnfDiy
CEQd+loxr7eqSk8Jv5tJw6vMLLGxqScOVu9VsXvQn/oDuARQb0V0ns5XQPkT3Q0x
JP67oUmhAVEYhDem0Upf3bl4DuI30yWYtyDGoR2L9Y2JGukxbSnPSeLx0G+heyP8
iR0u2e5gueEhjWjQPCzZL05rPq0LaVDHDs7nKF4bWUmTW1YAz0M4/zM86doWeG4/
x3hvAUY+SjqMi8WeSkbWXEWsxPQdYeKaRaw2CSe3s3gcfatri4W8C5bOBuVbSl5N
AkiqU7GlzwPxGNA3GOjhCc8WXwQpKyuvhkFJqDrlQaA9xG1AaTJdJ7Rf91M3zZ4X
fNpeAsI0GvWKwVLz6PSIBHAqWjanffvglJcPVtL7b+l6FB9jfyivCJiEXQ6hd3md
tyByI2WnKLkKJuDbxTl/9aoQZsgfCzYPXefdopnlSA2UdR3EssF/RLWz2amt+yfq
qCst+I0gUxe5VMYOGcx/glDmQMn8YtEi0aljJJXmxSn5E52KXD9zCye2famMIFTS
QvMXl9vDyWVoP/Ok2y03DsQcZXTRhMemcRIJF35LfUXdy4tWwU0NPzxwru9zps/4
HNKSbq25oeTmhgxrSm39YQ7Mj7G3ngCToju1HImofHbcTOc5vcjvYNV5CQOtPYVr
/mOQUlk3mSvUgvEGvoyzYe9Hk0SEu5U3MjtvLwOZfPVxKL83ecsNTdOrZBVOE8gQ
hbuxE729tI8QTiyzGMCft4nLDMHlyOQA5I+RGhn6Xb5RqmDAU75n8QRA+dQyEQXu
UlV6kO5JJ8RErkbUDBJebyvAKsdGuWNZW04+5IJdkobqrym7VH8kdcjqbBvvfOHN
ReeYfm1gxEvUwi2GdMftXSXhF0DXlWbkQ5e/6kmFO3gyelFnjbjihEotvyXkgzmS
dpVW5ALObnJ5/sydt1muvB7p5/l1MWNpqngj5QY31iJDbW8NpznKAsVig5wQTPOa
VneV1LGaaQGD76OmFj6pR5WwWKoxqR5UasiJwbnrRS1z5WW7ST/rjdhqyxfyJywB
3PgVaAqPweFguqAS6ft/TGUfWfb3Mu7MGlN4yOVh7f9clnxS7bBiJETuvB6jpfIe
iXKLyh/c7bxRVGcMo47OkMub1Al73kv5+VgiLM+D0GM98XYEfR8jOjbAHiCkDJMW
UbTosIq8DzowKF1kAqtnlBnuMsLjYddkTw4mGBeOXHfPxkotPLtsREpKQf/ojGGU
G63JrMgMrtB+lZEij3awAdiyAtRGfEbHBgHicfbGul3rAbFmIMS5zllhjfzMhRx2
NgA7vT+RmIm00c9KJSp3Kp+CYvoPA4vqunHe1W+XaFD6m3SY2TOuJ8XpyIZXnFQb
l93aVTM0evRj4ViQ+3SKwDEpzhT7k5WN4l4oMwdhYE4JHTAGU3YFxhHlkYQwEZos
bmbAzSULubnHrGnuvuNsdY3PcRwWXaTi2LXK0bWIWJaiWXAL544ph0baTCs1pUTR
qElNoSisd+ll+gCcvfCLrRalwoAcrsEOrY8hkf9B+XZNj/MANrgfYctjDPrlRlPx
vgI3IY/1gUO6tI/wWl0hGaZwolk+/Kw7rrKoD6wlmzRLFnnWgRM1xLbsCJ0OG0Ia
gO3u33iKCj56UPIWqsC/IOx6jZxDRovam7KyIxvbY+4roChoxfZvr8Z8Hp36nYFv
Ro3ZFDS2vtJdXodLEc3nKebzce3Z5Nj8xiAArezU7vrKpyjQiRi76kWKSy6B8M2t
VtZCaGrzeVkV0Pi18ywSh5B7qSu4eLQ2OFuxUrfpsfWS6Oh11LiXhoscfREF10aZ
v63R5gSpRwclK+1srSt9S8/rvmljcnNdfZBhGN7AoO01Awkwbk0AQ9fpkleoJPJW
0msXSHw7OerPKU7dZG7dfPBSDLYWtOoEho+AOIn4A1gJM6AWO4ryT63n/lAiIA2t
fO7QGwa3mbjPdKPOtdGosXB9f4e4juFhA2Mx0dnUK2Kzt9B3kgh7p3gvXAMd/ngg
itzLV42sQn8jFgnVsD857aeKj/JESU3tYWGPe4yxJo07/q7Ew2NXB7dJtFcgc86G
VHSkrgrEek5ZKc4FDgy+KAjKLAhRN3UFsW0f/Fq1Rh+/Z+8yN94nhtzg5wn8JX2j
jUy/Wm/T2uZKTTqJOWv+ym1Gc8Lcg0YEZYm4pB2yJqlA3lFaUwQM9plWgQzFWPmi
SbgTlvMdgfrXoZPPTOhb2fO+e5CEgnlOGHBQ08kauZ8KO9HLuUPhpsE8nTgDzXNl
U+2zRdKv+L0tRFKB3q7yyzVK3XA1Q2XwLfXLhG7pWEqnCk4IqZHdglfO/RuF4eeF
4Alz+PxrSchRVqRg/uCqVpqbEdDFyvrbkRQOM9wwF3uRReUMQJF1LHcjliGEmqRe
ikTSaEeu9+RqrFEF78UEjaBqxSU1RqqyfuDga7dCyehrKrDjVlOaZuMMUk65irDX
72CSeajag7I/mYXfY9VuvlgTf/jcQpCshu0u30pF8ncRojDRA7IR+g9kERwiGA41
RnwFprlqKDGVpodJ9oFqA8+NjnUfrSgcUmBKFYKrkeVjbIDv//ani1d6xJdbepJs
GbpqSvh9uLmm06k8agSM0LwmKQEdgSJbFhKx4T94kX7rPVf2Ls2lRnE7H2hSdHGp
nQfiBA9eeF7Cy16zEZvRdk+35rTFi3rSqk2F+M8PHSvXAzk89p83Jjz5fW1MagrS
kx+kRh5ijgQeGYWbtQtnnBRy9SIFUvcFV/2Wd3Ufgo7HK+lyUMCwDWeW3nKbQNbJ
/0YxqvBkOhZBD5T//c8Sdw6e80moX27iNdKdB2e9UXFK2mlDvo/I508K+5LQv2AI
UsLFCRaxWztSko1mcS2cxxr31xj4rzeWp4CPoJ3WI7cg6d0GMfUnM14g86DgJ7y+
ZWfXiyXdDNYndIonc1CsFUZLeUMZn5+vaIOhAie9g8wqWftqwNG6r4wKK0A7ELWE
FpOb9kxMSVqSjbL/NRKsd2lzIBkfQ0tOyIeZ3dEmhNmRdFY4oDH8K1kaMTgVlU0S
msXlpDx34wwt9qzvdAn71wTSPp2WpkYUv6Zokz/Tnjj4ekE1eECw4fRmFflA8uUi
9PSH1+FLIADDWLvL5NgjmmaNFar+ffKbFDGFmoRCVLs1X8kpiRT9XRFtKbJXbFc3
iXJejEXJacnBEdbXr8KauEFQj0tgoHb/KnortEek0BZt4RW0HuCqQa4Gj/XF7mF1
CowgoLtDXMzmh7/aImfBnisdxTVbkkP8v/IbZk+3NdIrpiQv0t5Kgj9aNv+t7OMc
loeEDcIrNLevZYkpnoAe5NxFLb/i61rG/kQAP/1/CtQM3LlgSI5HraTspgcNZEW8
1vF8aZANzfJ0COLu0drp6VOiZf30iyxbxoDm35O1VKtxZ3gOFwnuIqLix6YsLoJv
efA4LU0veugmrNXXw6Clu/h/S5GZ/rHh/tsxdFo8u0YQ1vkfZavCFesBjwqGFr2q
g761EJQ1eyqHoCuWUSbd6Ocpm+JlNLZ80zkaFudWk+Znfnx2ob1HPAxxGyAlMjpM
Tt0q8Vpty5KnycqqFfIArGCY6DWw4cgMufFBdmbK/+I1xGIoZCmH1yj6O5PnY+GP
jez2rQxWnp75fi9wZKLflgLV9KfowTH/61abT6frFgO1QmM4HxwVbF65WDiIS3VG
LBfsKl97BpvOpVKvrK2UDPFGTbmE2od4xQoPwqBiKpbZnZVh860Sbm1+F2++nqSZ
JoeODVzm97On7meDoXdaycWKaV6MdIm4nrgYqyQsFdyf2IU6OVUeCgTaVwtEPO0k
86NC442RPkMZNQ/IcvZ05KIZXyN2fwo1jv97fbPK/fgNPAXyxXI0a0r3L4cHmGVw
CxcrFJXUjvEdpWR9Qoq9TTG4LrIHyDCmH1cz0hPm9J0BCeiw0ISl9GNb+QKSxC8x
sUTT2a1Xcx/Pxy8jESOdAV5V1kbe12qJNj2lnwbnmpZYwSRKwi1bj5z7I62AJuQu
W1bbiykjXMzdKAbYmsf5d1MewDvHxT4f/Csf++btcwaXhH5uKlMbjc7dTrmrFhTv
Z+YZEwzjx4fGzyyQ+klypcHyAxKfz+wZT0jFn7WFgFzkqJ/BWtokxS3I+D1xmq1u
dQFZuRqZouak0yXWHopgc6vyb/7ihuh+YzDMeYKZ9vN8EUco/Ui+uV1Op+rvDtgL
R2Bj321hcZnxJv41p4na33Z7BdE+tfpGmcFvlGEK6Ng5vGMRt6wP5lIU44RjUBaf
26BGBMZK5Tpz7Ba9QdRteBdna7/gIJj2NotWJiIUceEYByp12Wqrc2CmGIhzkWYd
SuKqMCaOxe2SLChW4NCTVAIfso5jQ8fwptxx57gDjRaNgzzpaHybWqH4Gf0T9sE+
azBP+BPy96y9eoApNOQWluTBae4rMTOGyOi4gl2Bx+uDwliv/18cxN3HWw6O1+17
UJXGl5hbNOCdVvYQNEfb70uiIel+Jo1ddWvFt6guY/0vMgKYMlXrBEwmyyv63aKW
CfJ9PGT59ETnc9b3AqNWyoMCbW0ctcOTl/Ykcd4Nl4VsAvu3lNZ4fR+P6t/DCkff
GAwsUw3vKBK4AcZOaTGR45aCrxNzZqNOieNlsjBYkXimm3tjQYJ3wNzUU9kwSa1o
fim1sSUTS2nvbM/mIEdHIwEb2CP6C4JTYv8oJbz/K9wtdPifzaVnU30z3zhHKg2f
9NEno3AjVTbKHx4gEbJOPKYYdw6VPIym3+4vYhIi4SaXodtNX0e6y8PUs84SFVUx
04x6rxuPRs6wByjNiG33SI53tetUpsQHJgAeHOcLGea2DgVgR+FUD4VccC0uNivu
TevNBB5iU1QgKK3cbBikp+R3nLUQZLV6FDDv6ih7KdyAMs/lCTQ71Puc2euJCp/G
sjajeKHPf70PqGYbW78fuE00DQ0qClD9/lJRMxqhzJAOgUCpeknhwXV8i3o+qJ9e
BPsV4KGeNKwCSvtTjUNELsVYY9BDVUPrSNQ83SQnQgIxkFzMxwH9rTKYMVfjZlu9
77Z4153TtKxgSTT2XSj7PbRfuFohgGxoKXdxniPXqeQ/RGDV2BwvBKtpz6IKrceQ
OyIVaZjdwn+pmDj6rk0Dn83+y7JFblP5TDYFoWrP4Nb1T6EIuNTxl6++UZvYGkXj
aXwPlLjhBqEl6Rdxo8FZ6QJgt5bfILyR6I3wSux+VloOi3HjPJr30UML6zSyJ2Iu
DLWpboQkSgrazLx5CO5dqcvEBUZZRWdQgqozXOwS0FeAoW06pNyt/fGrP/3cHg6H
h4IbDXE7kw4UFsJEa6zwuvoapgW1pbnW84SaqqewUZ5vsyWF9DywGWbhjt26gTSU
GeP3VM/Qc39BU93hUUqvX7jL8GII80nNy0K9J8L9RbEHl+9pNgygQP4NAmEm326J
cxCBaRz0Ct7LAHb8lMowyYUg0OSLbAW6HM5jUmn36Mip/jrLUI6JSebDg6bsmd0Q
o7Ugpzs8LknTJ869+Pui9wcygIo51lvt5hOEqqcTpYeCmTccDD2HNhYWAFuY8JR7
3wmVv1UQC917/rywct2F5YHlm+Y/1CGHW1Sa1kMqyYBAnCP8abjch61K21H82oj7
nWjZy+IATaMHh5Y8UVu5iwRsqEHxp5G/k/Sa5Usx2lpy94PKeIEufmBbzkxVH8Aq
Ye5vHoHktNKY3p4LXqXA/0EuvGguf2QyCASsOcdYRP/cCHlmh5csRP6PGR3p2MGZ
SJ+JVi4zD3lv/pta0t9NvSQZzkXlylcAs1LLSUEX28CWiN6TdiRDzsQxVCarGeSo
NtCrDSmdTyk1AXKey/CooGHRx9+J+bjcyvR41i/DdekWLCNQxvw+oLPfiPg3Ue/P
EEaTLuM+20YUNsHj8y0urGksVcj188Vi9xOSUl2jRgOkvFTWBDA4i3WQ4L8TeU1P
KMslxdlVXt3B2kpi07SB0y4YKgXLeg0p9S9jDl2kBpQi+K79HQV3UNMtsgBkRrIt
/Ko6IdEkfp99w2EMyrxQgQ60CvmdLrq+jg4za0wxWRDh+PlsqCjPlzON7qkrmZhI
mjSmazwRqqhN4o3aW39HQMWuEWrPQSREcg8FGx28NxmZftC6i+fTBnbMLBPRduNi
lf0aAl3HmL2qTwBvDZsJmCPsdpbJ3sRa8awdQv2cofLrjw68rSqUOUkas68Lo2XE
+p9wVKTwi4zj82ngTfsCI/BZsDaDhwvjdXwPuhSJCJz1LnGymx243LiLsDPlv/6o
yyXG7mPkwSDrghOlnQTPjCgudBXd4ewel6EWz2gKEnkFmGFpmI6jJceqIcaFBRtp
+3OAeQAY9p6jzJF2PqrVYsgcS6sGmGlipRWtcJwYCA5hQqn+PYsJKpEIZUFSCXyl
vNFnmoiMhruya0IxVhMMMlejo5XuLDYbksIofuw/+Yp2xOFSqkuyan9qDvAd2Zds
Zt1x+6gFupjiNzkzzq2yNVlSq4ND8ALhLOE2veEHwddEadJQl+rK2wjT29Pn8u7w
fb+dTZV++G9jtr8/UE7VFPpDe4V5rls8PIU+PtbMwTzIEmwhhsI3Unx/ghnzKTuS
E6IrNd/uAMUfEI5c0SqAAMYbYHRXMVuAuYoDC2CO/71vkkUvlfXPrgpu8fJahas6
yuTvA/LJLp7awZBzSPi6sK6gqcZEQRGTd4DLQeO3evek9kZ54fYLhhOolm+QLhgk
yGmE66wFcfCtE4tQx5+3a9us4JoDWlldfXla0TWXxxZ5RGiWNltYFgyLDE1O3i2y
muZDwufCIWliuocaTdfjbEMBLPhnIIa/9zVV4sdfbZNwgFQTU/o8wijdu9u/KIDV
E9fK+yx+PoOB8W9D09+Ji1l0sqFd45daL/FJEW1blpQdS/lnhbx7Ls2kswuZ/kKb
7fMO8DqZC+y6/WTe4i2so1pRUH+aEN61u9+ml/oYNjnr8cIe8NE1lFnvM4cP30cF
B1MyqzqQMfZ/wnTR3xczjA0Eq19f6pO2xpwxD1WLJ1nnTuj+NMTA7VK7Wv5xbP0R
1KFuiUf42apHUk3RjFpvA0V6gXlfr+70Mp4KqA/xo+AhwcXx+DJgvRAK21+M5rP0
0rMVCjNXdu4hCrB19FoAooiQOR3v39r7dEFoQ/wtGPCHxYrX+N/qa8hhWb7WQUqf
DXJqs2xeQJpjqJ1UC0+ha9jB6GPZ4rInByShNw7EgE1cXBCGg8zM05GPx5M5cyvx
cU4qnIk6UBkrpH9eMSvG3K+DbiiAceQGGNQ3eTYAA8vvTwkUffIaJdj5P775AzWH
PgkqSm4khUv6EOowIlkt7LhwFyRyWsFkkJSDCAGRv95r4WJ7/EeP5wuHA3aiBGTs
U6wRwzsE/bP+qn2ahXgqmhGKQm9MzlU15cUL1bo+IQXIyp5ZoYTyft8CM438/Tpv
r0XTGFV/9jtWg20cHyNIr5VZbm+Eha1kI16N6W6I2w0Ow+LwaPc35yZ4I+pITFAJ
rnwR2t8OsApXkSi1FBqa1F14yahRGFT5E5GmnWHyVltSK7JDRwbZ/avICzU10e+j
e2HURml3uEt/vSRHUUT9wbYEn0U2bQO6wKwNvnPgZAl8+J2bqaUOln54r9vzGxS/
lSUuZ40cWIHQKFItAf2URWoJEdjTra6EbJHEw4QbBEVPXOX+BRcH5tN+tCBxPe0F
U33w9br7eZ9wJLoG1+J5FKs7g7OH9UMZfiK4PiL0Sg7wafK8sFgq44qa52e0/jG2
U2TjRa1n89jpF6SmuFLFlOsyyAc2mSEAMGDoP5B8lpBqe7ciHJbqgOKUR7qGwL3n
ewAUEkj8GdqSQKk+oMWcdbuBZiv/gQr2fp/Ed3WbJb/NJnpXRPZYX8XFYK1aabvC
ENQUre+4imybqhOks3crCx/HVD2f8VgAXAcoe8PJycKQLdFxFKIWx9rajvjv75ha
UDlR6GNVHfMegJYgiSuS59fqSqHzBuSqcrAKCZNMVJSYPZpTBJI2zOOqlFg4Usjd
htqYaVNc3WdF6qZEbGL5/BzyYayVsniXsdHWx6DprARB1KNJi5WSxOvPV4Zrq2hV
XQEy/aiD3IqYw8s3qvxQJjvU9IYd4w73zzaFU5NDFOXpHW9aCFpRHxnn5WnW+Jz/
HiEjhE4g3eJNKyurAI3MF7v93+5oqZCYk2cCPJKLFSJesIkTQpcPmcxN72mRFkld
5tJ+goqonLKtGkcPvCIp7YcYsP2gGueKTry14KNP+jUg23AdNq0OMgscpgSSTT7p
wy6cBCZpAq06AtijqVWk8ut/6fY42UWWt9BL21GyxwBUGA+LtTsDie2snKTNb7GR
JAAn61AidC51Qz0Vc423imR/LvWzjTqYUgQB/GOi/agsDStgyIb6FenOXLrbTpX9
eFN8osrjL3wvkYr9oQg7IwKYDAZDVbCVvaZ2zR+54mAImY/gD2JtB/V/NEb+PXV7
4LdhuVe6q4hSPmSX1jVEAcem9Gk34e5pRL53M2aL8PLhi0RaKwoRXMa5yjwULKJQ
jsRNq8sRqhSM0Jhjc1kXVFcnlF74URJGB513qIWEu8U94NPNsCyh6+fNi3P8fcZc
`protect END_PROTECTED
