`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l4y9Cjz6z2Meroq/iPubXhiFmfgzMQvPwvFC0RCiRWpb6XptfH2zWlChn1sjpeSb
aG6oF6KSzKZASjkYxAlN0ae3MXXm+lzJPW26Exq0ythBPH2H4fSdlBWHSFfDMZel
6bUHhnzqWf2DgQVKat34OMIgIg4mSDxeojZ23wpMET4bQHsdZzjH0kj/cGYyLT/E
MywKWY0mTdJNW2lN27D23fd64nX8OtHoRvbj4ld4a4wKYDhTE/7Uu3YXODI9XBzj
yu7niSebW/gLXdhvY20lHnzJVkmt1yuhZoQ9I3xlW/GSXPhkJr/CLez95KT7v0fD
dCstKLQ7EZPQP2f1VP5GTpFyGwSnnCI+oPY4e8poLmeI/CxDT2QvYMc3HRQy+kyx
h6vJphVEBeBUFL1WuzpgeFgXix8oQ8PlUbxm6hh5JDDNJToLUSijiECCVq+ZIot0
96XiTdUl1B17Bys9gaPCZXHZSFyOBuhdGsngU7HXTmE58SER7K2xyQRjICcWPTD4
WkOQ6Kw3mn16eAZt9rb2UOxsleRZ3imVRVddPGlZzHjyfSZqpUxWlipqmhbyWCJT
w/v2Pe9zNy52mMi7nYFXo/2PRiUdvvmmchO1rAi0meCNW6SRFKk1Oor9rOhr1bJq
mAYl0jGXx08p474HXi1EXm14HICdXfxyzyIwKlWbBUeX9AJW08wpWW1H0jiheU5i
SB8jOanGDu3k2t6O/3EfvBHCa7l/x6fWW/BfWkNgniplQRO12F3q/ue8xVGrp733
q1Ap5vchtmT1XkDPqAW0LWuQIzDIxqb10X+ep7ih6XSWg/rxFMixjAHA25Gp9ldF
g/4kBr9p9E2q2YeI6HqatMbYFBpzHLY11ggNTikI7Mcbc2S3F64cgJidPHtW36Yy
XqcxQ3NFV+78RxXrXDw5sumOEAD9bY+JvDiY2B8W+BWDg7ofJf9Y7uVkxg8Gw2qZ
Z6CYDkDxOmppjMXzomv42Cn8VItMaMNqO1E9SqsJXgKOsuk9Obu2vM7ERNu57L/d
UnRmbDmiuQbAIw2B2dxVJ0tvY5pRSDE1kna37uukamJCLk4Fh2qzHz3FCFriNUxb
bTZSrnLO2LZKt+cJrq200S8FjprGCx6DBOh2OQWGmS+jo3NIiX9AF1NZwBE9DLJL
PsH9YIpitgyfddQjSEzgorX4HizBGDAG/55MQ6DBHF8cWXCsawCilDid9toUJVju
uWo1gMXVcKXXAJiV1GvRtvdvXr0TURX1BPg/Zfh+4dft0fGbM7K/9XtYKunwhzDz
`protect END_PROTECTED
