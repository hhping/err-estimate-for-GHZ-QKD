`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a1VToxLxIIiN5JC7Ga0zfXdWQSK9M2Y3X3EPLim4kFi0ozVPAZhrHKEHuorx6D2v
pzNL6kOYGn+ZPj3w/Zal26YvidEJF6C8msF+sAE+tTNfnfy/dEMo4r2mLDiKMOjH
en3SH2cmLut6gZBRsXwQ1XpmwzY4WHXd/BWkCXw2DeKiU3cCehtV2XfC2WyzHfu/
REuJk/YtFeksPpUX/6kq1BQGQJ16glqyWRqOC/CcAxsOAj0Pfva4M78fRTQ0pdxB
ZQ0dVAP1fETNzo39X2w4OcAVj6TZL0znkn/mjhmtJq5V7Xk+5Z15iGgfmorH2WBv
I+sacdfG1PoSp9rvni3ugKBIK89Q3Bi5MdffmPImSf5ofpHLpjNtNwrM5wKgCE/5
VbGkUFRBWanOGzOpLX+eeXzOKqK9XOLowox1JaBqaNmS+RWfPdqYp60uq6qD6ySi
0QCGMbxlZcj2RvthYSS3N3UpTKCQ0eCV9QhlrwyTTeJ1Fn5nwEc0E2u7IdgDIr9T
WwKcHATT4mGHelDVa5NfB/zcTrlV1f69LwrFuTc8YZEPTIHaVy81D9HRC6hkl8Br
FHA8G4MSRq6MuYq6Xk/qTAkhmkploO53nX1VN9G63oAVQNxg16A31HEPgH8G7rJy
V4Uy/vvmZ9OCnVFLi/JnMlx5AS2+lXHdg1+S5PpXvFXm9nDaRbHNsyIPzKpfqAWx
FgaMRw7mxan2ncIXpGyUxEed5DAJDiinf28rGL9E+KzIuytJEF3rh0BVg7iZnjJF
MmfUIPxTMGfH449iMmrBrhoFueeCKqnx5gaPSuh5niD8oljKdKYhMzQwJzSO2Dqq
Txi6fsqoDP9dZ1QUYVvD2arEM6zHlMJscm1m/fbEG7QNBgPUBkVyG8m/r6f9z7j/
N92tbf9nXYphwzhJsg/HzodgMFKa5N3lBQEoxPLtmoBctGx7adMJTxerb9Mnypbg
cmMi0Z8hm3rvYSxK3dHStgQtPjw/gBi+Uyfl4cAgWcADGqWwi0frg1ZDUdtFxCjq
pYUfeNPZuiLl/01wLpcGxP2EwqOHncTowrebgzxDQ4loNNrKLrZma2kXoJWj6GPZ
rvWkz1nkDXELak3SigfVlw8zfj4dCMzqOYdVO0cGhKUxyO/Xo4Hj7cAEgQsk/5Lu
WbsstvDp8wlq0lBQyCef7rMSKKhGOOQJBDX2ydjWWQN1DcV7K/ADqlkAUoOryyHG
VEKqAVcFZpifVP16gK+SXCt39u+IHNYaej2cxORefI4/wfAyKv1I6w8RhrZlQRX2
PTybmiSrB0DrKoc3HPngNF1C0DcTily7PWABQvzanw6FQFQhnYjE9kt7hQAgX+OP
n+/1zL3aHOTdoLLs5/rTIZnbJSRACLPzlCs0KgeKZgq5dxAmEYykNk8p3NuhVVG3
VjzagbS46QSANgL1sK+81r4g6M40Vxh9mHyNibhk7e4ruvrHbDH2ZZcufW5SBgq7
kym7ejku2RSOpB0H2BbsOoUWm0o5hk23LtBqVvfbPc5xSVWVZdtkfeyPg/GZ2Jwv
47t86+O7a61eBonv6Ys9LWvugxodxDuB4oJv+nI25TXo1Eopx/OF/KRVpQXff0f+
CaLnJI8AIZ4/B4lJl4TCttHMYBiKDpm1DJtR1QMgecGtiD9bRqmGWmkGaOFpngrZ
SLMJDpz6KC2xaH0lt5NeVvCHKzOk/WsbOEh7dqkl6Vb8sdnxtlWYXiBJ+SKwOo+L
LVgFHnvMFXcQ6CtEwrKSHbuQZaUrUd1O1FZ3IAGaQJoasubqd+/6oTjzl7HsdQNU
X7Gz57nLTtXDTSUkAD09zMs6tk8RghBFSxnVFt8DGXU2svFaIN7yNiJ26F8bRCEO
6Cp9d3l1iKD1N06DquOGKBHP1eGhUFVcvYCN0YEp8KT0Z1XAXbgkYDHzYQH4YJ+9
LjXdvhKMBhrMDpSyHL9zy7BueBM7u1OodYFHrzEaxLSuHYaHHCZIN2CAG2PJM1Sb
vEIQvwVthyhxzUJSezGdYR/vwF4uaeNEjHLFgB/CokbmLIfscqFC9veeuH4J389p
oap2FEKl0m7jy/kBKqAgvBKtMm+0N59s5YkWF04HdNtEc+7a7VxX4KQvb9lTjmUQ
AYc0E6xume/RRlRXgiuEzYVmCbUj0HmJmNErbEFLLPyGTgUXXpNItAJxwWvqiU7h
A7zz3EfOuuMJ0wIvUnp1tDcYPn1Q0wYRwJnFSw1dlLSJNLOX0tBOH8a+sNSDpLrA
xgIUpGoFbzbcgcggkIEXuti8iB0TfjFTiSfL+ZOOBHrurs9zMxSTy140I6uIu7B/
Z9SCzn9/UWV0Ta1oOvzUPrxy9XP9JdGh8WoCesi/xDMPlSVPyqJ+f2tBpkiO/xHQ
jmE9DDohyGGQ9rOTM1SAK61Z4mgopgrUKrw745Smk0+QkOuVumDMFtgQk+/dBDhO
VOQT+0ryQQ9bjKIvi/mv0utNZw73WofKLXFrBzDPG/KEB7RacVUljGJBiF6UMQew
NiYj6eaYsjTj+W05ePWEHxnOyMQ3D8F2aAvWRX9MoJMz+5SPxjN1wdPr1m1ik9ej
BF7ZrcdHiwMM20dGKIRAy+Day1SPoWwakI9+lhXru0SsrR+RxqD65yBoJ28ziI88
2yjSN7o2PHLf0rDYDdqvPRFpQ9jLWv0nOAYjE8h3LRvHLA11eA8AYAFJS/KWvoYy
FnR+69X4HXneiDdzvWIodM08Pskpog3VyDyXUynkf+dE8Eka0Mx80C+0PtI9Hp3V
8M1Sh6S9P0b5OKdqPmXgMniXNiSZ0sW0WDxixatY39FAOpwifpzCqthjnqkUaHDp
2S/1srC5HHBNS4KSmIN/BO8cKjyHjZ5mYL9DRD8n0SKDKKBngVuI9D2QD1xdtmx5
hEHC7Lu5dqXzGF83wlFpQ0qYCGDsXai6e7EnGJ8iG+daA453iF1DESAuBEtGUOhb
ex85MhtLiN00f4hat7ImtzNUTKZARDXoVL90KmhPUEHEmeFkqLlgLjD1SyvMcb0H
HuFh7b7OU2ciAZopDlVM9DillZdvNAZOeMzTVLuD6b9JLzyygY+j/4Rf7Bq5l5TX
f8cxNUS7BcIonHeb+LUXaz/qoov7wQQ3Xclpvyfo8+WrcpDPR4VZNDx5bnwjnSJl
H4TdQZfLMV5FSlXtyM5qWAtSp0g4CDQl1YO21okiJZpSaGbNTmF01sEMt+/oI2ng
l1SO5gAmIOQs8gdojf9TOc0MLbnDb9KNMTlTTbvvwg4GrcFvsOW+IeZFrtrTrRdE
PtJS+0cf2plFQ6cUU9+xBFIVbdyQcgiV3YrTSbIltZ33jv9P/Q3HXfo2iP1XMXNB
ajR+ZElUhNIC4dW/XdAPTYSm7UvAg1C+BKjrrwL3Mu+wpLkiS5+lCeYAnwrgeGOf
OmWfUCauPPeGSNB8hhK6mlcCXBjRskAJ94Fir6q0SNCZGocuSBIS6A3bqvXsb3/0
iCdBFkpgKNr3VjQ721xmxRHXU7X7xKeI6bt0pK88pWEwjYnOolCzxa/Gp7zZPvBl
S7L47XIri377TmAkScAlZ1lHTsaBSXCLHVoImRdYCJ6FZV4646KmByL8J2TqLYL7
+jVG9lXp0P8W6xS6H821me44XA2MXgkYoexZGR9Qdap8Wf3WUlEIiRx+oxfXDUta
NnCJHkGuU4OoZbtgaW2PDoPAr9p3CjFDgntLDlB+5ltvCqh2HsqsrTsW3SEtRS1l
VpuaeSJdhIjQwDzi2QNg0Gr7dJSFlaDfuc8aqKB3y6UayIlIw4vRkVqxcVrVF/aC
FwVG0SkkF+My34xhd+zjr+jqYhqo4NA/c/iVUiXLknjuHhKVSODr/LBoFln6fjtr
37yocsask7dCAcNLKl7S686A0Su83qsKlWNU2d/2Rh7a1NZuKTudBPkmMb3aSyUA
WNruMrsMxyC1VVCD9tkabVPysQPwUS8yzTeyVKsjnQvK6D37L9UKZimanKAoIuv4
/5Pwf+M0dn5hk8ZieoBGqrqWjD+3r0+7QHwO4yr2xuMQs8xGN1fIl+af98Dk+oQK
3YOQIHAbeasHNzQ7U88GInA06/zadphOXMojgvrR7CzBJDeXGyEn943BCDO7tsYq
1wnBG8CfYj1UNbeeMTjQgwXqaqAqMCqMqFR7zqFmM9PSJweYx82Nh+edAnwsZtkv
3A7KvALS7H0yK5TTE/PwAo08GeVKnv+YrUnzcc1xDBsfXmIfdaEZApREmfQs6C3V
b3O99VvgkuHMEkNgslQVtEVh40ry5zE6lL3ujGVvT0lIpXWKdS04cnzU+T9NiT+d
9DJzxF2+irAvfs+rFEeG3kGsN3KsIOS8QA1SVe5YqWRkTlGBnJLh/U5YyQbEeIeA
B2bCULH84i0pOYGr5cC7CTtZ7HJgbZ6q5b6dIC+F8d2cC+p5PhwykFmI20W8IZN3
k79yDQirLPnLPIWI0p1VpB23G8dY15ulDt8V/lWmkIQ3KlK6CX5nHQT3kfsOJnLt
vUnT2JeZU41sh98/uj55+Vo1CyKMNUflnvIUNu/u6taAbC9wbJyOH+tOdchqIKpu
kyv4M1wiCKIV1HOjskThooS3XtNth2TCNZDRyNluhlofbFYKjkIiP7Kns4kQPleL
xAx8LV1/flmutFn/90FaA+xxUxIU4/d8nLNxgQ+ak2LaJZTr/RlydoOfE2N8NpXO
WgMuTLo1fqBw/kgeeVF5cT8bJpazr/qgZkxYG357IHOhUt/o7MmJq/Zqs8jtIEsv
uLOXB2IxdRDZlLccTJKwfUzG+RFmiNeWyNcbrHlqYBMJDNbutX+7uVYiT9YI5kkr
nVdyIQXy6mMbyOE+481eTkf8IXhaOFG5tN2zVjfvaAH32+H64GXg0uO7Pp397I0Q
pxHMoSckoHpxqBKBVXhap0wQsS4WOo5gPR76EqfCz6+vvdKDG7x2tg38Eww5lJ1K
HhfVWd+WdivdBJnEFoN7G1WBm7KZQvN7q4Ms6Ub9dRj9DY6ipiDVMo6lse/J0WET
MB/MQVkpj0T9exGeFgojbDEFGXO/UG98Kdu3dj5OyXq3vhr+5o68BQDzjjiafqBD
jO8RKARnYEdXQu8jjDqoHY9JLmqonlxGEu3EbhZ7NgrCs73s9XvYF4K5fni3q/dW
fcL/6quKnei6jkMbDgd1bLCf5DEs1a1j8UJ6oDKbQrAMeGNfn+YTFoRLFekTKEz0
ZWM3JuxA9B0ONP72q6+LmtssNc6P5OlLis2hpgJ/H6wTVWtRtKBmC79OVDq4wbyH
xMB6aTTl8BrxDdYoTvsY9V/cVqQvYJgPnixxRA8ojHMlBQruIkcdTRrVbIZyCu/q
SXkkYyPMhg9+bxaUBQhp3XQCZBkl0p8CX6JFb4hCORoSg+z6f/4Dn64pNxEb2u6O
ovnx9y6o8EdjtIk9hh0Blg==
`protect END_PROTECTED
