`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cuaYh6ZNj8lyal2R16RfNgupn5lKGeIM1i31IUkvgSiuiwjS3NyGMQU93VdHrFKV
zFl0AEgQ4njLpkL1ApmbegwKyf0BJdTbAhI8KDd5/eRQjw6+fnBbqxJv9J+Vi5rf
DkbsA5Jf66XYt+cNFDJQNORTkH0sBUAbBAjqIbEVeTPh5wSXL1msmqwv6vgPa3j1
nGAPjIjG9dqj0frTgMceOlc7Byp/+xGsDxN0x7QPH+6KHEsg9/9Q/zGVyUFtZDYD
EjncAqKEumG2VLGKIS1o/mtbibBI4Ck34FmAdhK7aZ+ebMLrbpKM0axq0WQIHuHo
A3QnHneQfedpjyX3AQVKUmCdt+kxavqI7KoX4GAFn7Zl0nA/fPMYcAGO7oXtH7hc
8Xpdc8ALicsxbSJtJBOa97L3NsQas3OugCCj+sWd27KGpJMtrv4yGEn9e26W8sHL
OjJDbka21yPZr965bSTZTkqNIeH+GfCZLi59lsUQVREktjhQ0C25Egu9Snppmq0j
LMmiA+IaCRAciGDO/uKJ5oMLEl6DaiHu7gaSB3sUE3yN57Q9yNUAusma6d3XoxMC
XYxyyHs+foMzjRX7dIOGiACL9bUVyQje9zvXurxeIuQM+UXhQ/AhnRTYJDnpQL+U
cM+2/DVtTezB4skn/cTDn3O5FMYjEzd6or/4t9/reZw=
`protect END_PROTECTED
