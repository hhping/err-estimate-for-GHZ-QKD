`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6CgZDGGUuqIyJhPdp+PMq1zUQMKnK3pMokuECjeXCDOvS3venKPgsJBh1d/XNqv
LaO6mEcn4mL1WRdphdjNvbY7t6vpbKEghRsLN5eN7k4bAMlglUJ4sNMqoP3JagVu
j0O9BDiiPCLtrFe65ZCMo8oC3Lu6HDbzOZ5Q25f4z/eu83jQAZKaEN0+PZ1rmVT6
rUkg3h0lLP1YPOMe487m0db5IVxvxlzdHgcm07DKeqIQwzZgol98zGZ6X/8oOYwt
1USrWlfTAcGjAlq8iYyyPyPN3DFPWSQvKoDl9j1GEHtPF66vPTtgTmYMrCbNsotP
JQCHgFZhFWvZwXcJ0baMZyuevGYyLxmLNzDAAYvm7YtkMyoruPgv1vDu6FCiFycb
0YYaTPMN+wdAAbslEuQ3vbbTw+PtSnqBk+KudJbDoyPwzYmqXIwmClD3tDRaktWS
8pKIQ5GtxFuv4gtsuNZP9cKE8kaHCJByNp563ZUJLwB7VMbtNPHChm5TIqpAwgIE
GDpbousURgfhCVGSmd2Fz8LeMAUHZhmJ5uVQFsCM1F+Z8zQcOvIpCi7UshkJh93a
oz9WFPMwsWgO4ur3ZXQchferp/iHT8OvUZZkDsDYJ+5Xl8wsP2PwmND/G5ByqkjE
x2uCVq4ovA9ArUiSQ+o7cddQLw7CpeGLApQKvDQbTy5/pHOLYPdk12oNdCf9WefG
7yFsaWJD1gC1q3HIBZkbJYoiS509oviJdZtXqCWM9pocLRgOE/JB4EzJL9R+JyTF
QOM4RvT+fctECh3OiXs4UOtpz0d2n/50dqecN/k7UwUJ+YOVsjS/aBkrV39bE5pT
1AErYeNR+LLBp7aAVfJZv+avjCM2UkFs4r6aV8CNNAoQXnQPLc8jFK5NtqYLZFuE
tfyKqEfJ1CfI6VBD65HZj/dHxW9gunT0OTZ9Z6qV0+7EGr5h25eu8acZtKDC7NzA
gzD2i0gcb9lKE2r91koiNjE2Qw95R3692GU9l+lZYpLJ7R5wJy9Rhyhd3hlnL4Ip
NDdZ3Ulh9eyNAuYf1ianJDlgPzfrtbxgkS3vbkgkrQjRkWFdHupfseUguAvwCwBG
gOU7c2bhDRJy+ye606gJN6yIxL+mtZuPck9E50LIYYVl4RhNO7LPk0cLu4p/aYSA
YWA1d5HW7W87y1Y3/KSTj4yYy2n3LIgM+r6lNH2cD1sj+prXBquNwC1jATlLIUX4
USUFRBmFlCVZtNWhBWoBYF4R2VxQAhV9ZjJ7VjFksTZcvp4tFMaS6lqXs3o3J63k
OMTvgodb4EjzYlMs8u4O+Q==
`protect END_PROTECTED
