`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K2ZXtHU1rRzM2qDoa+B/diYp/se3OsnBuR8c6W8n++Q/lR7H4nf1h+sOcr4S/TO+
j4JtWD601HY6CN9z0BNDwR6oOyk0UzjphoZEDvwyELVp0iEHmHwSN00GWuNgMNdR
qMKMK9/xrN1aplZPsJp6q+nDEbt7zmMEJo5Xde5QGZH+46c4jhdoigoj76xlj3Yd
RO3KPNusklyAMTdvMZY4sEhhhxH8dnsuWkX+U0QrajpFkFi3EKXzFQ7UaWNcE0yq
1x3d/VDZRq+Xt/slhzDiqiLNrQ8zqDzE1ZEthc72JP3sbRFeoOuOdzQcAYQxqAcE
gPafo4qNDBs/l9HsTIr6yq7NIMomoM9vJefJfUmDuP/AjbRdswaX+TdYrribrpl1
nhps90HT8ppPN+hG2P8fQs6Alox3Tj/jgKftvqyHZs7rRi3u200JqUBPYWVE6y3z
LxhfeR9TfuZbRjzlFwd0IlnZU4+XEAO4tsJk8Vn4+AmSZXiP79TE+XhHNnF9f4XC
9jsIeG+9Id83lvXtMR+EnsnCBy+cqZ6l5WZ+6jMreGg6V0Jrb3w5wF04uAj/Qa91
I7OYXxD4UouQQL+0L81xWAvKJXWo4YJPRektV0PzsnmcBC7psi/F/MXCbJ4KCDYP
KF4BKaUbJFBBEjh7Olo9ucAcazPYyEoBXVj9hP4bSN8CFdwskjieAjZt0bRgWjLP
cp8A5uHDRIBk32SJc/TaMFbITnkMSqDiYjHD6ldgdfDkmpm9Q/VrI8Mje6waJz53
D/jUPIfZIemUUW4wdLJIZz+BsEe7ISb09GD2rNLmq7YWL4YJK+1WK7O7u25FtE4E
01aUhp4wpmpJ1erWVpj0YgeYFLYZaRWY8q2E617yQPvEztOsuHHgecpnjoi4y/S0
8MUT/drQal7bRUsWuuBMPOFPY4w9pINsE+q1AGiHjL4LHCgWdWcwXseHfOF9EtP8
HpecDPkylXuI6Ds7o8VozILdWakkrcA/VjrkhPBt5PWQtuloCJKCcg4yLK6HuJD1
T39htkIoc7jXkwvftj5lesDgytkgQNDGLyTr5H/lTV8ydqqCFF5FptMtES2tf2N/
ydTh1h0lTUVDonU+h+yHmJXsY06S2c2DrTEcnq+W8XwxpN58G86xRSpai7YIKVYN
5K5HUasVnTaoS58SWK3ArIO4SPGv1T2qUm3j/hJvLWai9UAtTeeFTrEoMoJRRxv9
PvoyX/hUk7QfFu4Xfuyw1gOrv9dC/HDJ2JzGOBKhnyGGjK+0iPPnU0y2hMevDY1X
VHO875tA/aHGSdfLwq3hHm1/1XK5JHPphQmh5EptTjOvKNKOoy301hqzM0a/BA4a
pOUcn/IY9aogH6OAC/bcG/kQZXUJFlzdvErTbIUmrBE=
`protect END_PROTECTED
