`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ckJqNChjTM/VwemWRbWziWzU7BzvPq63srTK4pVyBIvmdoyeltKGU2v8+ySgl7Ye
q5GdRkd/q917Qa4k6Mw/uD4ZBYFWmcDTz9Z9QAQmM0/W7cNPdHpa9iNi1XZ9Ipvt
nEixWLvHmFNKI5fLG1d6FXsjtqhNv7TWNCTh2l3pE9Yd0R9/ciV7B0r0FD67EUsC
Xl74YIZvhp6vIv+Ob9cyqtRMfQBLb0d0dRnAx6UW468ORfUrBGTsy7Aq29M82CGz
18mRbeoy6Be+qFPdfldzTozCvsHek3Roxbmamw0sh4JAq5zlikmsrRrzQNhmNdDU
6hLMGWa2mBygdcI42MOjV/WmZqJ25mhMkN1yPOESizfijxLpLiM0BqgEBfmhhiNO
a2udHVQuKlNcyOfvIQYAKv7bUf3nFRB37dU6sNGupYtsjpl2j3uaJbfPJrI85Al8
Y8F/1wC52NBMi58UeIkbJw==
`protect END_PROTECTED
