`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1YJyM0Fpd1O1twtZ2RPW/bCBtmvO0jRKdvIcyHMO+C5F2CBY3TI/G+hMgDvSZSy
tV9psgOsAwYPFIiAQjVSYJ1G3cMzkbWDqLLIetkfbfjT/llfVvZsFEhG7YvdWDON
/1GcjWfajAXYfLIpWcsxko5wAqGqOas2ykH6dZfF/f1X3OBzR582loojFrda7dME
HSnZCplfZ3VHUKibgiS0wmaJfNx9x9KujZPFHsCuH5kHmJ2u7OfJcnbZXq1DpYfm
e/3Z8dTBXeR6NBA7iiV141nvz5X5nwegFu/7ayOqt2e5A6GFQrEA+HmN7NyRngZ0
YgbyUmLy3DVZ4NRj/WpYuz4OUsCDk+jQKIEwN9/FErivHVxBJmKb3xF1S1Bvkdbw
9YwEVBNNkp1l4eJNGie7D/3G+kGv/j560BkO5Lgv5EDyTz0cz5IdP9I81RCeIOV3
sJ0Ao8wWBsXpgLb8meUX7Zb8aPy17xN2V5KYeF48kr2LhteZHt2Y/yXxo5n9m9jX
lP0u8QO2iS7o6RFrR5hG6xIyj7sRInlSrd/dWBxrbVzqjvRJrSfDJHy0c5+t1a6W
uiGchgo7McTCY33y/+ar9l+mGFaHmkxmNPxvWSO1UIU3gYRwwhF3sYKIzqlX0Iug
LhjT5OBIM7dyYiARODoCvcA34W/AynN6AQtuiDgD/YQ6lIQA8pjo5Q+3pBkRv1Mz
g7LDQmJg0zP0DMhruKVupzKWSUY0XpGPy8A99Bxg26Q=
`protect END_PROTECTED
