`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vb4UGSI97B+jrA3AFqvm563XomJ2H7tAG98/LYxvwYxJjBrYe4rYDpo7VM6OeZLk
fN6+GuFRl5ymOITfm10t2jF96RP6a7iEJtzHeh/qlrXeiPHW2Ce+PziwtNLlixHf
PIfpazxDJdYolkpGKAacLeFah42z1j+uDcVzubYkICbEAo3C0WjZNTUNlGHW21yY
oscOVGAQcednIzYlS1CHfJ7z8dhTAWG3GEqkeLfN9Yh0eFPTOAA+i16jqQds9Hup
9vtNB2jLPb45nagSdGVx2Pv47UFed1ni4ugm2u3AR3wNQIpGrAPECm9k1TP73iCI
assvWGkqBh4hk+CWNalkwq8DuqznGeR/pIFtK21annBAF+uBOUMO7/KId+LQxZtO
1UqIC8KzzhXMI96AT29rz8Aa6Ih9W8CIYi2lFN9mFPpjazNtPneCvtXobUsgp10W
U6LYESy9YA2em10tVi4UsuDJWqOfYGaEvoG3ISIq3p70LC0NONmO1Azi7Dc8baMT
BZc3nVtqnM2xrFSnAEy+Gl9qB99OPsch/kaX5yLasVMXNrhYHrFLSAoxBoVQ92ny
vlKSCDZnWvlK/DxjVAZN+VYIgva9P/M75EjQrF3Spt3H+ndMtA8N0lA5fvXjF+aI
+7Pipzr9BNziVHGbm8jFuTDzF4PGHy/RoSExHL+NmZVpaxqOEUoLwOxjl5V2gDa0
JXiyEc1TZEQ0AtV1K83DtWPuth2x2PYd0lXrj+6TrulMyoYSpPuwzJXFbh38PRkq
2H3E5hZWK/FhrcN7qOD35BKv9l98MHEYD9AunzmwIzTgHOFIX3683+zxqhZbiFS8
t8qw6iLSbEjnYM43xbheIu13r6wC3vMsiL+XbABY8oY=
`protect END_PROTECTED
