`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLrk1mVmGIutBvp+DgPu6LxVtw2XLCPCpvioU89SYji6Jf327jfAPgVwbiM9F1jg
2irrIc5SaLuXph9HccCMcxDSyBQeE8VupeUee+nRrKA4iiHVACQl5h3uhvbvfICa
G2pOPHDP3Kj+NemJtQVKUgjVoPNAQWs5DAeixhM4ZvyiQ+2vN7VgbeF3DqSo8R8s
2EnSSfJyRpkFWLyhBa6nfIcrEs/gqmTn2N55Ibcy3dq8axAdLn6DysRLPedVJxlN
ElKD54oAgUavuKksvq7NzWNSfHd1hn67WUkRTWHOpTTfzCjjAv66UH6R5pGrR9Bx
`protect END_PROTECTED
