`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
keuKoHN5GIlznfHnYzd/7IGPqR2s/rBMyrNOES1bhdUZC65uNpq7tqrzQ6o3Xl0Q
XOOdgMie6KoqFqrApxYUhQKZyi9LbnWbuDcTVsqViDHjpR7tav/Bv+Z3nbBEs0d1
326NsA0WCO3EnMaXcbJ6gBaiz5+c+YCS9/b29cCi1kSD4rFH+LPDUOTgLPk0ZqJh
Ozvknmaw78WZ6djQr5swNQLfkYsaWbuTvA2/E/qnNwoq5fe94BuUWKu8S9xDis/i
z2vtB3mFn6VaMZdZwrq8YrbxHW+VPHR/gdTK5HxWC9CTIxDbjMa4zyOo74d7rtA0
otd7aA74VYcy4YH51P0fb6kZ5f7xaYW+7+wzSQ9T84uhDCxBNA0we7UInjlp7i04
EJ4nDvAzyNo+5TmBBQfLWVbYIJ/XVTaD/4MclKExf84exKNWN1B0e6iCdjTCCLoa
n9vB+9KvFlV72YDvo1uf5bUmEAgnYnpKqkdebGvNPcRf2D8kAMn29YhTPXivXgj5
`protect END_PROTECTED
