`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mbip69Ero/yrTyWxkZB/+y3vJfH9i7rViM3YgKK1Cvgy55i/JsVSg18kW/5gTAau
am4BLmwuguCmTTq7G6bD/E0FF/uCeorOqE7563yinr2Z0IDdB9oCRoVI1E+9oz32
G+oYvuBd2C/zm+N3gfpXECLrpWbGoa0DBDj3n4pC0htpiXIbKeHBfg1CSIHwLxTJ
6xs+83JgLCIuzXq8rBrohMib5Dw2pSVtZtk7beqR/RBDCF9MFMP86qpYAi4Yjpb7
bkUbM1g/4CwPnWQSzq91y3eMqveu2+IgpQSli6ASsE3iivkxG6WQtbUW1az+ec9l
1/b2DdmbRgUnSA5KcQntngv31OsV9HlLdOqTnbau3feSVRypaXXpuc9Sj9mudmvz
TfeXDoL/4FM803Os2rEFSZja+ecqAY9R06G+KxdawEIO29XgGbnJOU3IC6zuVUEJ
E58gVHNHxhWs4vut4yFD26SQmt7izFVNPkhYFEURI8IZlV+8A4PQmrtFif8eQw0X
9w31Xifsos0BHUBhjO73fl2mGH2iLs2kCYNIjMJ85eF1AC+zjeHBgzHRxSIoqNXS
pqFqC1wg/FNgikq9Teu7WsHwe/FEd7lnWuNf7ImbO3nqHVN6d4LW479CVqTbCdWO
m85m9/SMbHD/S733XauF3cUjLFblCmNUpYFKsuD+B4MRG0f47issBzeGNXrqa/AZ
vyyNCOt3e9k8YnF+Q7Y0Mi/MEVwGrauKu2EoZDWj0m3S+lWWNh+PzJyBdGOrsi9n
XDd1y2oeFqquoMrAjZQgLsAOdnimewTHIqdWZhm+10qJXr2vcDUo0AON3RnQigMP
3o1zW7+9J39EmdiM6OsgJXOGaPYxxF9tEL6HbMl7mD/N6VJqymEFVgjh/HZ/Drxs
lDVtrNNr77jFz0QfHCVhRhRswoZ+umwphA65pZQkV/umzfsRG8clo2TuCivbYRnb
e0FydsChI+VhuWAEmKWfKrjvl2ppizNSolLvKAN/g03vL4bBNUXVmLbaoh3S+OQl
YLNWg4s2aWHSzN5ZR7oyTkxXHyuoEg6YAHRU4s+ho/zAu9emcZr/JnhQSGBbixZr
Zw3Ml5z5zYv6NJ3W/2MPciBnzaRagqDj5ZQ6qQAm7gM3/+ogPkYschjBsBeM++Jb
Jexy640O1FEZlEiPgKGtGYcrk4esqjPFPr7O30vWOcNmFYO8htsK93Y07mfrN6t/
7vYq1S0AnBNEE1+9IgA1KH7mwD7MsqMkONv+HLeGc2tNuDfcfDydwF0foWNIZ8Tz
t+jmtv1P+LeE55Ph5yjtemlLOQ4ieAE0GIhP4dHm+m146FeDtWrODf59pvogiEVF
vaDRa1b9Spej7ZvZT9659bdN6cVext9cKNrOPHeBU1JlXPhuoVx0THeYGd6hk4OQ
jQzCMbCuoq6t/ZfX18Pk9w==
`protect END_PROTECTED
