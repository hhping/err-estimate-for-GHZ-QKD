`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PaWmi1VfB8wmyZYFsnSWTjoWqyT/qKyzY9p51qX9+ZNTtgjMCleMZwNPtzxsukmn
B2Yee+o3KJY6Zl4FbyCHhICN0ZLJTNKeXDWD8Qd913/+tsGExox5ZakaTamIcOtX
gH1Fa/oed/06kA+M63oXCr4ncHVFlWZa6dgspBtmvOG7CjMbXZQCLnumra5PIihB
4e9JWaZgpyymP1Z68yOMgteG2Kvhxh9c/W/iqWfKwNP/tJyLrAtp+hqV/CC7ClCE
kRo4VVMMy2gdLzMOlLJGeVyN46W1aAY7pqX9c6wEN9a+RNY9JChERDdbfn/bhRVn
g2SVTl5xAZcDCIz3xdrEhJ46vkT9XBQP7vWpXF33/+BOhgwVTg8IHO6ZOGXny5d6
QmBkh8VrqBo7oOMX/aYxzXF3VUnkbntFJMKV1hk5yEx+qm0xtteitCNu0fE8emFu
6JmpFjkHSKqgElX0NQgQ2sQmWg9fAmXBQkUoOCtT3+b2mV6IgiLvrNKlHQpjMPWc
L2L4h8tpgF6Ybv6mh4bvmsn7kS9kvA/lWzVVdlLBLZ6XC26G0TTbtpHEXmh3GA/q
LP1bMaaFzrcffXPLHvFvVE/HwvkhF7HlePHsxbGuIPRWMcv1dV5PmJYO+0l1ktFQ
+X5QemQoPP+rVNveI39H8lYkRLFqMsu+HJyYVll2KEtcDrWgLmlh1hIy/zZ3kzZK
xYozC30DZk2Swy2q2Rk0jQ==
`protect END_PROTECTED
