`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dCrRQUwRVTUze30zUzIj+CP3M/qS69SJt4RkX4mwSyVhX7yNWiKPsxx5ylOGtC58
wLdawljFmGzxHXRuQ0qQz4glBsJVIjrVMLevJEQWrn0tBrvy3uYfr/wZFW0Ach3i
inLppAnwrfEwB4gGuKqe8Kp069r+79KdiBFYEVTEx5lei98yClUX4KXMqPOA27do
ONlovlbZQzkRaHhvUcwZjuUuwnfHh9eWaTVPoYT9rWzEUieK0DK3cKvvpyUl0UPt
hrKnkhoptNElqRLsQ3UW/TKt1ni/Le5a9elHWFWRty+tOfobDcDNFPceIPPRimkD
UZlCapfeYpPO9Ao1NIPXcWD6k48H8/2ovGs5lUJDXuxAcAIhDH7mE/fW9TxcUVDE
/Tryvv5YGGjnxnenpaYbJVV9CbgE3JA+Hu7e2y7hcdxtYQTgrzbhXi8QUSMIKK4s
vDhfuZVt8SrR1B0FucLkyHL1NSJlqdI65hu+i+GSNSBnsgb8wzxyoduAg1RgyHXd
dlkv6bzfOIfFpAqjVAYj1qPuKQxlBK0UWzrOlHFmV5Q=
`protect END_PROTECTED
