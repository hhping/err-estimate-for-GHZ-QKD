`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C82Bw7vY67kOSCkzl8Yv9rmHNmARuaVEYZXBSHWr2mjF8z7TVcKAUQtdZBr4ESP7
sCHuIse1QxyZ1jWEWZmhCTNsA/b2Wt+kPwH+uMwmbycYznX1P6KA6Xp9duKYGDVU
h1srkDPltNHoTD5P3u/2NWOBnQJj311mjPbISGwe1yZZ7K7QTdlbvbulGJhXAF+m
SQI3aNEk8IcjZIeHbutk9EK6sdh5Zm93sEJDCOHVROpNCBJ+WGPld7vOj8PqVL32
lOdcNRZmgNDQBzQSD40VCsRXT2eyo9Ej/zB0pd1f1iBU+ix4kvqfuQG7Y8A5VhHy
HasZo1m4GyR2qgQZplJUueEAzhYttbCHj4FDxzLnyZ1kcSepSXzY4iBjRuXCcGu1
V0Q0SEuoUNAW0Dsv71T5wcL9vim3NuKjJ9MwCKtZ6z1/FX9wyB1U3R6XXpO5LUSd
uM+cimbOojXX5HVdG3OPc6rZedKOPYwu1ajd6uWDaLgoQWPi/URW6GPMuLbH6QEM
bGGE7GFX48eNv/JXmZ1h1Ti8CIuaykDniSl+j3Vy48zAEN2kfxyFyoU6fO/wjJtP
G041OUgecY6W82LqIvynUORN0pux3V5ndI9gms1AgiShrTgWOLpg3lPUf22hKBac
XbykZk8sHM3YllR+txXMx3UcJSYQEx1V8n1VtFaHtW3S/qSiGjMKriSY6CVUj64L
3/uFRHby5mYSzlBtC4onoaeAdFus2Q/dOlEUSNlqFebWtqudmnwp0ywPn5j8BqnW
rLgCzQMmmH7E0Jrlj19yU6Ks6sbWEeK1DdVq+7jEYgzVI1vi4UYeFABtGDCli5BV
AmNToT67OJowfuLUpK80bpI9K6ZDH3xRX6yLkmyq2HclOgQYqd5J/I1ac17axOMp
hOpQH5DMBhypp9yD0M2dyfCT/EJzzJLsII9WI1x6hJSpGYG6IVML5hw9ULkohwNA
Pw5dQ/2HtbD6lirfaD5vEBf1CytqnwJUx/TijiQMKXXciU3fCWvlhol2DHpdmqCx
Gd4djIBq3E3mieDnK9a+Bv9t+4iMM5L5x7F4vQO0f7CVF6ZUICG5c0RgjQK07ZMq
JRptWQ7cmOW006S5Tb1GOzBeVIw4/Jhd12b4izSF1deia1cTQ7WG1TkitEbYN33y
EC1lW2g4luuez5eYQ8Rkl7/b+/90vGlVxJvVNmWGqxXuHblvsCljlHXMTWypypMM
Pgz1vm9nHxuetjGp01NFmg8f4Y0Vgg8OU5LgUj4BzmqEF+koMKO7ZwBDklszHY4v
pKGBtVf2tXOacI9gHCwU/2zeuSaOY0skxrrvpM8T1NllTjHswbnslKDVucB48CI7
ZeAJ1RWWctXhBvzBu6a79qSnQ2OBUQ0Gc0y1QBOOFGP9Kvu5czMQrmGt2xVs/Wtu
g+0llXMfNFrS3tLScAmdhdEajgJUWse9CqcV+gjTziZg8pLmanMJbu72JkKCLkQX
h0gRNeXpSSiD6HkmYUHa1nbUxCmj10ECEwxjJBZCYKKJdcI4+CjP0AkF1pf6nAKH
2NLyISKCZNv++iddZijpdreAMBVnQRZWUc6cUvDv99WVPcZYOxDUbr2OsVKPPhDl
heFE4RJz7HjwBY/7UM4AIC9Xl5VrBALMg41OB/szX/lokv3LGsJJUlK+oSpDaTzv
IFSRabD9kCEUgeHjrK5AwpuylsuoLvocKrX0v+jwM4f7On/EEr/zA/Ud9tABUj2H
JGVaK8/UIpwk1YuneqaQgZj/TFgoJEh4fKcb6ZT/DZhbEwZxknttDkaKBDmVzP9y
NG4T3l1Tsd+VY6aA7gS1wygK0ajln7FkZvjcGB2O80hNM/2gXAMyUiwFprqwAWN3
Ah9CZ5o28y7cRnTtoKvX7Nd/uW+ynwoY9cUa5D9l6OC3Gcj0nSg26b12J/1+1Vbn
3yJzz0xKkeO1vzeDgEEkn1iVx/rOlG4E5W7IsusEVlXPjEuJGh8N51gSnMUDJM5X
HoTVDGPy75w2lTHdzXNNG7Yxf3f88xEYigBMhflgMxJ0QwDy50GmHB3MbjXwPrOI
DuEPJf2ScJ03VYpZrPE65ChLlhxceAGlfWF6X4w2rQFLHkJToEB6AM7zgCemMRjq
A4h+Vf48pvA+D/qufzHUQ0QpykqulI0RMNpJ5DQSubXR9LUouM5bRCy50/+uT3O6
pQ0p/sti7N32d6AuF5sd+Ghyx73RpjfcYuEhmg84EZ1n+TdOMp77Gs/UuXkntNMf
K+3HDKgda/L76HBI8VUQ+r0Umu5FFogGvuqStasOb02kvaiAmQWUNzN9umRrm0hp
6MXCoYWTomYZ7pjW1eu4nbbhgKOJlZQvxWRTG576jnLrUtzGa+Zi0f6uDLiGXIlC
cJWNrvKKxZtKy1+RuowdOgF4erinFOSEs40k63TJEXRv9ifM4wdZoRlF092Vn++R
wisw3w9FSyW34YUYMXSQ+0rnx9N6HJaCionUVJBWuX0/gUiPh03dKneYHSEJNq5D
QzbuzEqbkYqPmTsOLFBrbxffQBF0Q19OcMOfs6sdqdhpItryYYiikFDEc9H8P81w
A5BFyLGx0mpozLRtkJzxppBMBtRM1S5CCGp/GBvVOFgROmSBatLN7D62Tu6Dh0Hw
gCBoqK+qxW++wSHYel2huwMdfHUCXg3DMLGvIS7dS0uHS+Lwnv9t2KMmF8w9i7Xa
blmZvuYbLaHzahawTRVteHWgrFkEytO5emqY8C6r9AqsutkWr3V6ICDQlRQns6bw
HYzOOEuiworU8PyLrpu//tBzNWCchNxFTa4Hvy89QxkI0ATh6vmrQtYJICbW6btN
Bb/nekqUeytgI1HAiCrCaawpjcaazRU8LRWqeZxGYGR2xId8z/EurZoI7gsIKpET
oBXewt5zphyBG49FQKbaE4R/6xVLSjZhpEtBchJ1mobvq/rQFiEDGUsOF8RGktic
h5H2K+W3BkM+Fr8ja+lOnntFs3NKyCkRPZSwZzkjkvZRGCs+d4KNHOSd0GY25zpB
DBPC0NqX9zvFDulJ5B87+mJCDTNioMhnAMNvQYcnY++bRVpvaeh/VYebBJwgXasx
ZNhCxedxxT47xrOaF/q/Tw21Nn2YWaSQPTrDvr7KSw6HWLDa0WxfLZY8zCBYhmMX
I/1ukJnNWbR613bOf22lgAHlzJNf1NuTRRDZFzcce/yERpow8IopVgxBnrEddnJl
oqH13sC/9Kx/+5sC2kZJM01BfH7Ezj18HGre7xpR+7+XAessALl+JZG1y0CWaUib
8uRKRhRbeQ53hUV+I2NZVEjXr3Jgqurow52U9YFA5sgPm7DfHdq9wfU3Wg0Fruop
m7nQmS2ClivPX3ttURVLAhH3Q3ExQx4UIS/eT90h03q1u++LIiLT4b5vgwDh/P35
FUxB9uM6mCsw034oru2NB0xny3jXjSDBQa25kU3e0Tw9cHRgBBYnWkb9ejKJm/Ql
IL+xKEjsJdojY4L10j8XW2l2cmTzD6HOO4ZogDzih6zJICSR5xUO0LnRWE1d6F/V
tYohN0UaGXuECP421wMtb3rluJbRbQ8B9mONAxwxT1NdpWkX+Pvz+xLXidvmTwro
xMRbyV4wGbzEietJvVCOuOhB0am5Dt2/xoHmxSDx/SI8TLVxl+LMjhM9f37CMZFF
Lg/bc945UZSjRilPq4Q2f6Ko/Pg1OdPxiBUqhB9xiOcRuEnxOUrcsQlNBKsS761H
7pfyJA4tD2OnG9IcqlGgeLQc3NAiS7F1hNGkDsmOT0n0w80/GqjZ3RxXy+ztsQER
UU1DIg1Cu5mjRT6QR5IzYxNgTzFJKWtH0fY2X49y9QhGBzPyKc37TugBwPQtO1nc
tzsrMYaNkife3KjoubYJw7LNtpKBWJs7bJSpAlUfX47cYR98DzjwaRkYrOOFtLfH
tH9ZUxCrcsrhZUK3tQKiURFhFu6ceSURxAfjE7sc52NYzwDSME3ABDWk5zSfrZIL
G3y977LKxuEHLZHM8XrsQg013LlqGo0SwlpJ1Z0dluhuWeW6jNApaLZGkxWBaync
x5ZR2tEjX+4+3q6MwWfgxUYcQBVW4x9bro2BT1/Y8xgd181fQOYkaQvjXR9BeVW5
99ImMlDS2t+Ti4ss4S/b5hGj5MpHFb/QZ4/kTAVRWDawaJD6LxNqYsS512MpOJD3
A3N7ItMlUa8v6YoZFzHdGmQ8cgF5I9cyTFgdxJHoWW1NRmei5mApc/zOKOYo39PX
B9dbjO4YnhZQXF7k4UTResyhvIzDpXpgxcMqM0vZ8jd1BkTNhhIntxHywi3uXfl7
+RT59SKY+ak34fWpIgTS3I3kqN7yd88PhZxtLBKa+eFN/QzNYdmdgrwHAI4vaC/j
5nwdl1ZTDTsy6PiaFvGmOhEJZJEUV4kN7qq5uDY3jXjIHwKi9eViFvfLOZZQ3pI+
Y3XW3sLmil1BU4VSCpaB97gAALW8c823IULc6rF5HX69XIQ4O/RHzSaSbxbAzTYJ
rwcPEqlH496tDsOGv4CoQUWhRR3bm0gTvcYCZrV3E56H9A8vTAkyfrR6MpJJjvAY
FktXFI08q5rmzL1Z6UcbPDDCdxcoi1JovpZJhcve0KxkOR9cpHHAjJEKf2D6e/uZ
6Qh4zYc5gOE0KJtkI5g6d/KT+bWNVy1VHKK9UORfqL1DZdAnkV+sIVsXvnyq2VFW
9cIzW6GCutVOwYQHd0kR6jo5DFHhMo7JcJBGgQ4P24IU4EAkbRr/lVRiTi5+z87d
y0tsiEdS0lY2GqUSfHYK7zhfwH5XJ2ZqOl9NpOxDoThd65UQJEm8YAnjigq+Q+4W
i85dqGtM0ExRQ/i++k6Lgni59TMsZnVyuv97mudv3GZJTXjzpHofFSwJRt8ehFRe
YaAE9T6QWLOqk3BN5jf9IJ63qy0tfxg3FFx1VfhzKbJ3GTcpNnz3qrglwakJCKTr
WIYPF7G/5Gd5qmSKROgAdcekmbmmBNT7VEpAeuTvIVJO5SgtU62XoivvvCvOxPvC
GHHethwW863vKLwu3yVQ78K4Bic7y8tgnGBfVOe6Q51HRjFZx44XnxeUOSK8oJZU
eNpTj/Pt8j7ocNHKZBCEFXzlGTLR4NswLSqhSqljNX17IR6SyYgMUlFkwp0OKWRL
QTE7XnVT82yShp0iyrKvc0Mg5LIfuIdjjPYnVSE1JK8K+C10Cnkzc3y2lbj44rHu
MnwkUyIfX9TnL2EijekMDxe09OrmY7B57ZZjaMK5sqw8ZVms4CX7/hjrw8HozRPB
meswppEaGPWWIUMahd6DylaPl1UGiWU7bLuhppxQP8VP4dupn4ReNvlFZ6CDWJAx
qIFBfFxCWGRkHbUtKXPNj0KDEpqMS9EHAVMMMePdTZUKfao4BsOBmDI/n6gu5c7+
4262ccZeYMTK22xSTrIAZkv+CLY/q3my50/bfshDg8RcqINin0fymGLcT3XFjaZt
dDnktlWuSuNYAxzdz73DmQqcfXP74m0j7CLcCP1Cn6xKFJZivodpCDnLW/BPJ9R7
+3V4a9h3CL1IcTsmeWQU1SeQj0rHTsi1mjpu48MV98xRxCc5yPGCOe3IUHAtCuQJ
oXV2WPQqf5VUrlRWJswnmGVPS+z3AOsdh9NQ7z3SHtl3qba5x1rE8iTl/fYQGXzZ
4OMKxc1ba7e/oKO6/X9k3jO+BPxUCK1Q5EOd69awti6U9IOqlnNl6aLEbArcGZ7I
pUsOp5XjVUW3rkhxxUD62KCJ7T2n7wr8zXw/fU61sK19zqrRkifnswYHqB+J8ZDr
ZkkvpnDp8LW3KPfbsyZ4oq0KIPJqRgswt5QTTsoBzSg7GpUodnr2sEP2Ovdm/4xw
uNhB4Sg+KOBCHhJvMyLo1PPvkMbw1gBN+wNF/qYLHcry+EKmlBwM8n18iY4w2KH6
6IH7VibiJdRILaq1CQpD243KRpBjOl0PbDu3qB4UBsj4Uym+ZFOiFMAXV18pqKuf
NSGdsW8LT93maZY5n2qf1t2kg50eATxVRY+wCsGrwfIj9DcLMCRoomwKI4+gJnqa
qMD/8Tf0MryxSmSPuPbbWVmqFzuJ5N29QQvtXVFU+6JQ2xSt+2g8A6IaAW/w0CMy
dQTrGPQHOnjI9OeaS58WGHsmYqZwicCGcdw7nkYQWWw+BwAGsEiEPCOZ9PsKvjhg
+pIXMDDhBGcQX0YHDSnwO5n6P3hhtL2qGAIb86+PfO33MEynbnT18+xjTBru0Nfj
39t8Z10gQUD2rbHLYGo6rv6ylk6wBrLlVv6yVs1FaOqAkgeLDCKQbm8JHgppv7F3
RF0hEBMA+V02MUKsf0e3xWfb/SmVFe9dwdhzl3bs5OrDejVu40sHvpENhrpt6w/M
3vjdDO+3h9tsu4N8YmPu5R8/p64yNwX9MbcT2OrNrsjoy7ZBSBi2sa1Buju0CcfT
hcAo4XZpzC2XkJsQtFz76TLa81h1BCORlUfM2UqxSQn8JuIZbuXlZuPfRBsD487w
xKjwbP8DM0e/tTkKlIWfdkx8tu5oXMoInewcO2149HFMWfrLokDn1XHH11H+W314
JKLKUMrioImmTH8dxTy6KTPHZ9SkrZxGx9EnEfZu6JJEpCk7PCfjheRwqzFf2UEn
tzhdUqOQNhLLK2baNqjCDW6eJKJdW86Q+b4pq0vdl8dhqmkdAcvczI7olXP4ntEU
88JL6PulK6q4RsHa+jKXvTj38RCOnNpDf4D83nN7vK8ufzwFBb93l5Qh9JpYcpKM
g+tnftVxgP1aSv1DmpG3ytmYuim0cM2F6oJETwh0cMoTEPfLsgrDy10Add38J9qd
9YBgLjsdg/vmDL8q4qGZCKl3uvgISQshv6EKjFqPbia/AiyFxHJVfb50OIbxKdU3
DIlqxZNqOP4WDdh3Jcp8oN4hr8E+G+AVjFT/2VJdQFvWSG8Y9YNv+2JT3i2Gy1Yl
80/QvqPq/33MWyn6+NIfmQ+tHJnPxQPr4sBz0cUsA5D/by3EgT3pGOAPjjbnjnan
4v+wnN5x1k38aihfVeSS4rSYTr1VdsfcvUVH9GKlB3HLmtnvpWdIA/hbmBZm+hGg
TEO8GpehZlOE6LBKSiwVMWpSGK9eEandqWauYavYgtJDTu6NQQrWx8eRe772VFYb
P+T6GILTWU05QRmYRqSs1+TIpt1sEvPBqZ37A55N2dtyVVD5zukPS74U+TAlrWoj
dwxnY3JExQs5elIcIqXbcq5GKgRNIA7RXTS1WFdaJDqhX1qcM0G8ypbEQStxdU30
kmGdG6MUsId/fgn1pWd+YxfP/YcQBf9E2la5PIfpgqFU8013bPEggrL29WIaCztq
skWuGqV0oTdyQA/wbBvjQjQINLYBLOu7nzf0LVeJUrB5INQ57CKYHsqNhugNArYR
fZ4ECx47fKhZjBlEKKb8FCYNr/52O5VCEhJPNtVMC4vbOSm5OIC5fN4z6sYWSqvq
CgGtrNH1T6LsuN1zjwQwK/WXMEWvDkxnSDc//eBWJm4MfyUbaJzm8PhIWsno336r
HzA2M0TxOITxQKRSFVXBjGZp3mpA+31EMJC7yZFXLry3mNyMEjnqPKEvZ43JApR0
u+nkp3AFNWNj8fgMxoMFGAoRlumzNQrPoaTRPSkmRQ77AxIC/wPb0Jc3BHPBqHGx
dXJyqCD/GNLA8kj1rvYKXSoxV/BnKpSvGRhJ6NLtBvxuyFe/I+Zla6VfUhjfO2mJ
gXSempaKjYP+y57OYINr3Fer1Xz05/NQ/NOXHPsudrpaxBZguFXLsLzszGNQfHu5
dn8U1nKKsDZsgAw1Tsg7FIupN0r3Xgh8yTN4aEKWORyV8qn91h3asYD4ZDNALgm2
4MrZCVNsgMBsfy7qvw2MNlcS06Ay8r7Wg2vnhoeeJBvWVPeBviwQ9SQqXguQgNjR
N0ks4H8OF7xShq1M9PBIplOJVnvUbqd93iLdaS8uQGDRsYRtbO2w3JqruK0DeS0L
TpeldXc+/XDlfsg0NGrj6dIoXEh7fqunV0Nsg7k1D7MOXPZIDw30chvvJy677+2x
uI8jg92B0Mte0edg8pYqvZLPukv4AVO4FsNqvMlSlrXZsHmMF+C4khKWskVzLy0l
Oo8lJZwklYKMvfKyhCiENliWGpoDXgB5a/a1RImVzxSW6uvDesScBEaoBFB1S8nx
jSTNdE2fENppLWoBXOdogiGDATZyeVgyih+aG+z3P8qkWBqIDSGr128giohCK5qe
dgLB3Asm4OK/jdpxYGpY3GBsc9e7fHPmNRfOHAOZ/Z/C0PoihoG0pHDCriSGq7eN
sj247Sf5VY3X8DLsHl17NeDc3JqeT8PZaC5OAFUiCJ6YspD/jUrLc+qWxJtJTXWR
EjKGYWW8+TafVDxHRmykbqxaq444A5DF8xRxQJhIyt5olTl12EImfEa28KNU5lNJ
GDv5favrK6A0lSoNZyivOllIwB9Mjik3zHQ5wZNiBl3+5SJT/BN6fhpozKDWIp4g
NJyVaYdLqGytBmGimku2ltkN9HijKtjaJy9jBchcgBmVPE5Nx5dpqlS9SDNDmwDD
bS+C+j+Jhq8f5h3A14NZ/1nvqOcBQqzegR9JNZVYqI3Q2gqAXcRJhDnobup5wRdn
BRzDS8M23LKBXM0gbfxzhBV0+l2so8GxkXtRp5KDQSuNRDkFpW3Hg78gn5U7JaGN
xyYVlZ2y2s16dYEzOXHMOjY8w6/vtbat+SYH/HJQ3evgWHsiGVyIfO3BcT47bS9P
mWlqWsZac7PhlCbFJ0586JY0Ua9NxZUtXbJpcZZaBQ4R3RIvnJcXz+NPPYRbSrhs
iON/2A4DTQjmwpHizlGtbT5BDvgHjGdNwgSgfPtEDJuhhhsDLWkoWluK8oKhPeEX
1keXu4iuvnjTL9/jZ23N4sWcaGj00aPVswQ4qNWH7akE3+ExHGY5nqfqaTuK/G+B
IKKObbILpvZc1cGVcxzJ84nHRjpaXrWMI73co41P2m/beJGH6eOZnPnfiNku2RNP
5dmuIGAjKNlTOtKqq5PvIn+QlV5Urm3LcKo4hFxT5VfKuj0Y3i54u/Inwrz0zx1k
pG+JjgzrPWwpbL4q6rBhrnQa497kcOIE8dx0A8i5MMQKTh7ckDrlyp5KYfFs1geO
YhoWqxnw4kn7KnggLMxOAtQmaowKT1KQUxL8XlsDFT0FHcvlrokMKFDZ15AtmrmL
JJTvQqptaZbWh8vqd/8qwERlBY94XAIJnUFfmQjadoUvAFMvoj82s2URl/ibPVPZ
vhnmk2KGeIU+ae6Y4vMoiXAKXHCBJ88khLqrwIPp3eZ6rUjVKPQI4uXez6lvLnnA
iy4z+X9AxuggqSNWmJwzDY5GqrGkCxZ7QRNLLu0HrKvbzJaX9/Q0ZBPjhY9pBoOp
76WERa8QHfh3NhGo9qTrq84JCLrQFhEO5i4Y0K++kWGqfFXkTxTxsxGppb1HCIPu
iHemHx5o+kgUHUu+60phKgai+KB57AtUmNA/ytDqIPD83ue1bYbltnAvOEakCBIh
feczDUxWJX+UqR4bp0VMLCY3fTqvpIeXC0gMayXV2UhYIFT+cZoTMXq5/XlNrszG
Pey1KsMJlXbuT55+epYrGMshFjZXe+K2sFfKO/XfprTz00YIa26v6ltfJnEOKzZT
GCcDJ0XAeqEzSCOdeT6fqV2rJ694JMsxAmyLTZJic7Dh1/bVxzUa6cVz8s7JKlnV
US9FhaMts93fP8l1DV0CdHffxCzvz5KP5gUEQL0d7WEXlbALdbbylJKVNILC9crU
Zbm1kexf0j+EMjzwFXnDjGiEiimzGVsZAvhwjNlfmjceAw9EuJze5D58moU0wE6f
o+uH7Czk+mXMxwTvDRKFZlS4XB+IDWe4az8nH1PjdaTaP1uBTdSeXTBrt9xdrj8y
o9fqcjwXqMpAgtfsZh/hUMdL/0UQelxJKKOqzH7EfsxdixsEphJ7nGkgjl0/RZ0r
7+RIOyQp72+Zi6cPQTYGU5EPh9iAeOhzPJ2GeQkiRYTFdM8Tmui8hCMXwHH+PXvc
wAaLiluBZza6/rv2/N5d2KfNGGcLaceYPXDWXQIu5llb5GMDrVJ4fWDuPtnrEro9
XYDFtTn6OKEA4CPwCUWlbMG0DjKYICVgBDslYhRM6ytim2+kG71V1tTbQRjWN01x
1H6ScbvGnPcZfOK6w3sEK5g1Pn5eiQxS4ibpHUF/mZTUNK0aykUJca8JWsfwwQSS
lsrZ1tBsZXmDElHXTZvFafWiJJKqVUBkHaBqlvtjPHmhKBuz4SnIrw0iOKH63y0l
wlnHpKx37b1/y/MXmM5Zv/5wT7VtkSIPY5umeELLUAG3ZQXojZE2fFtI/+SFh7/k
UC1Ja+BAC8tjMUkKyT8b7visFiXNbgDEWzFlOTvdM3Khakfi/+hlyDqWjSs5KawG
oR/BvFEJgOVle8LmujUFyQtIycZkpdIt7BAm68baUtvZboXGBfwl8JI1OMoodsz1
SlTi+PpGdJz6M7HLfrDhoA++K3mT5GhZ6MsOVxqkqaswUMOgM/3N0b569j65Mx1b
G4IrBBrECvJ6vdess1vD8L/94czgyZOOyPouWhxWBNmQsMiFKsW0mInZFs+xMzG/
pPnYl2Q8h0S6PT/r2ICqZ9m639ZrF6Hi3g9EwjZhux/szOHlNBr9pJrZH0rFEleb
tv1nDlzr6Bn9Y40KXQ6/F0DIwGfF/JLxjfM/EyOelOAGGo0pAxvrePdX/NjezLgA
zrAz8TPRYhRbsfPln4IFEUBd55/iVswUuIN+mRvli0vFval6UGgEm7Bx7xegCwtp
7EEPyRiW9wHkwPVujoJUAHXXzgGplGPtpbQQcaQvQV0+Mc7V2rKXpWjlB+zzEYKN
PgGMI4kdSkBQ/4NDH3Xw4cOgGecydwa2nrOiluCs2AdpCoe+cdRDdFkKFtRHcLKE
m4H2av+ViBKUzhtY8WYaFLxs1gbMR7/OKrjbUQYVdBe8+NnSiAd/HrJrOmKxR+6k
9g7AEtAb7Ee+Y047R6yfIkP4D0nYkW6/gQagSpmEJF+nXiz2h3qOYVMdADTEQCn8
coA3L36+lLSIHbDhS9REUgsAUK84iOju3tiTsObAymzSYnQMW21wnYwGy85YRllD
K/6HVQvOZFS9mWLy06vRClaS+ro7FESLZdcHLrGOXA8B/Tx5oV0QrflqpxzyJIP6
MRUI74yBHTzURivXzt013UcU2FShXtkcLGhTOStPL0iEP4clEYmDzWFUmmhweXlA
jzNHX0h3p5AvPF2suHuUGnyzizwD7GuCd4oUzqR4kVU94t4TSC8N4SIwUrXYvoDd
0rsPBSVvrMAmF7r8/hQZmvv8GT0fMw8P7cvCvCvZ4TFvk0xE/PrvpoZkX0OXUXSM
STYO5S6N/bOM0b6BIZFLduJHWix2NCoW/rhvTh4qm5+xd9G2Ukr78UZg/EySH7V5
+tyLgxvifVKpd5Q7HmMmP2PYJ8qe+cBcRMFlZv6Q7Tt22CYdEf/DQI+8TQMKq1tn
ajWxoCahYgcveFN8hiNOlaGDRs5qCwHtb5mslD+bnekP/8xGPZN9Kw8LXDf0Q1to
njxwXLtWEYdU4vYW+21Wv5/r4cZ3XmoJUC0y2w3NBOYsKEGn4bRHu7JY5y6KwSRK
UkG9dHilvqyiUEYrQdBBtrfxRD45ViJMJjOESL+CFqP+8p0C9YnnAaYwjUn3QxGy
AVSNF7R9CqLa1lru2FQYjottu+MOc0X2oXXLmG2qFHWDqz/aG1IW9X3Hyw4d+gq5
Ezkg/a4FVEg9rwFWZA9nz5UK/wUBXkOD24wrd4dorfKNQ+rLhHTTZzWLF2T4amFW
zbJbSsGLqsiqQYlepJ10jZL+j9NKhLJs1fEOJNH7VKBlUFKP+SQYpbeIlCRc68Qi
2se2I6bqE6TpaaIpGmIlFRyVtKcYx0rQRm9qEGnC1b24evEAWhM3tsGsM+CCJn9l
KoZCT34qeU5MC8XMHFJT/XdkHcOWGZ4+Styx2kpG69ufMhPGqIQDwsafWa5vBkNk
N5Ygal/GmTr6ovhDiThIblIOF+EABOnn+4fnHdNHEP/oAv7ho/ophFI159gGckaG
mmR1K7sBLRtF9p7ds8Z8xkgk4J/1dHXCE7L1fsbTg++0oMysiaOj/e2EvCh1QYTs
cwLbKlL4DOj2gWMKlZltMPa6BPsM36O+mK3RZRK2r2s7MOQnd06MLv+KAzIVUeKG
OWAD+yanTA/WlmhWJ+yd4XkUdIKqCTFGF+XZo0F/m9V1G+TAYWw0b/LxLqQ3insu
qvZe+4XZutOnOzmZv0oh6Or2N1G8dL41lQwKE6pa5bqf6xdm1st0dAVdN20STXhP
BNgT/jjkcn3jkIaNUlJmTF8dV/2khnkrxzjcqSyixuysym3Hzb2fRYbi2yMKooMu
IrsgeeIl3RSTqGUf/LfnnN2BQzOLPuMCa7uYEUUTBUNBzrfsg7a9CNb7cKpwWV9P
yQN7y+kR8REjBuOqnfeRXspmgCLpWhBzvAOHel9Kk2duiIy4Ac0ZGmYUNZQhi+Ux
eb40MOT9sF1RRVAFmcXXoJxW7Z0mjdt2wBG1MWJWNGEonPkaDWGHSZbqGZVBVTJD
ZEiS92d6w78Cl4BcrJUF9WxPYTjpcCC8TRcE9QJ7bKMIxSKOhBxltSsmZQQ8qROu
1IdeEzByYokekrqSTo/Rr5MT5Str6Y/RU8aIrRhTZd4Inni/1OdUg6BYtGJGdKTW
/+77HQSlFwCkkFsYrtysCKnw5Zoq8HNPsasfhfUjji2PwI4p7P0pMa1+0VBcNbLy
83971pmTOHPvSs1NFOgqnP2+fgfSKGHdx/OeH1LVdj2K6F2lyZVevxtPqnlxZzIA
E6Nc4UOIYcsJXSUVJl+6azm3EXIyhGyuvkkPzpOYDSdPiErqudesHifJtfr4rgnM
iQe32iulZcnO0VxwSgaqKeprmvpOKZP/enANscovTNjdOBVr1PFCoZATelo5zEpC
2nr9t7hZut1bcEHuboqVBfLU+Ym1Kd0KrVoLdps8rABUuRXhJvqydQmeDrBDRkn5
G096Ll8i1qHwOTeQDntMCdwOXKN3Q42tlaRowUUyTvqoNugyxsQakXkH/oc64Zwc
PhHGrIlHlHnH6yZyWgMdOlnFlA9bMjHrY3U+sfvDTfRJuWApg2lK+rF97+OIuRpo
iXcDoBDuO68CVRxxsm2CtHSuGjD+H3a0Ep/ZrHFgm55CEpO+/mtXulf9gKR5yWWs
/B7rNCeaDwnHwNBWnO4DUurkaex7ge08iS+aKXnlSJsr1W+6Bt/gAUZVTRNBHcFe
ul4OLnrXHivA8gPAQlQhe7pKHLnpKywHEotd638bx4luy7aczKsG90C7kCkdpXBx
/D7wCeIWI++5SUAzgH6td7LQCaifUtrrRmQgoyKpyIs1WvnTXO+bN9YnljXMtSmg
G40K/twxAkvwI2YIeC3fCt7qUKM5FMGDcvdvdOJQnhf1ilizmvD47ow0qukXubOF
H1dzgyXHrnUnKEM9rPEdq6m414RMt5QuS7D59tcdIhCk9+L8EZAdUqJp5utlNI5g
VgecVRhZuz5QrZbol23YPvH0r1/1ADt4Qw/htbJNE5lXLTXlqBudHk0W/n3AwdiS
wNyYvtX5B0YOlbkLAIOQ8LjQSHNXooFnGD61pSmtzuCCLKTdX4oeMlc4/hYmeizb
U0hdFQimYCKnOfgKJkvbXiGS7T7BtUftQUGHK5/yOiurHGDG/tu+yuyidN2qKmzZ
PtgRJBHhxef3fFBGwd4LK1iAfPG6v9zP+36IycxOzIhcmBJPoqgmK5evzqH3S3mr
KF6QYVCCAxpM+JrWJHf49hVNQYyHkd2IDpnw44KSJO5TU/ZKtuOdTAocJwkbVrul
SJJXZcEZbfXs+TserjsPsptFp+FtiCd9CTJ+4F7VeBteIvtVElwxqGk5bw4nLXw5
mkF7oritClyDuPFcfkO5f41pa1Dnhq/6FAjs1eqjdmkPJkMD0cJDTwqgadagTqKr
V+iwHWny0XSWhpRZEOdO0vQ+njAP10GnJ5YZWteAg1mJS6SZs6+NxQTxTF7+BoV8
Br6AeHMk0wohMI63BGRGvsdO8LoyG9zSC9qt4RNm1BijFHcHfwrmBugnO2GwF1qN
YYZGXUylJmgSV9A4J7Ty7AzwA2cpilF3pNQNJZwcBERJMMiqU2iKd15wRXJFWVnJ
TSxuqO+O17DzQM6zBIg7KACmwykletnncIg1tIl61s7WF2jF7LtEgujuXy62ZE50
oUcwg+lRA2IsfiblrdsIutlWrEr1uTjcAwPf1rwWufEazOTzv+6kO5N9n7KZj8cT
IVjLcMjM9U4Y5TtFn5pfXAzcIv5ScMgWke7OW6Njbf29vsXCxPIQcAoFTj2czDgw
BugLYPRCLQzaJHnBPBIwj7YU/pUShPNx+FqDAo0Lw8mUFIANw0MhxUbxb8F+Q1S2
qaGzS5l/BSbNrlYgMbj9V2NoaN5Pzn2D7udVlpuPl9WMNj+AGhyALI13RM3reEqA
EcHOG4k5DJ6m0n5zKuIci52SmCFoqbI1JUU4ZNXeegItWLihLbfDyxQBsgTHJCZ3
eye+SfOp9Qf38iwCyvx5P0J2JnnKuZLdMgFCBtDhSfZLWX5y+GT7rLMp4sanyq54
sSYcz0Vi+eOprGv/N3xsOD6tcpNHamzlhj+6S4Xw1P1dZ1JLAZzheH8funjjkPvv
C8t06XelAe/dUzadGMabOV70MngYS+MFFhJP7ZQgh2LA6mwln8/hrjyn1GibzNVN
1V67lLGqPssnk1curgc/E9T9P948lIF8VXF2rDmhqa25gvHEScyV1ZSdQPsDYA+Q
6+LdgRHDo5wdTxhmGc87MTNN26euzTuOKsnwViXVgLJtqL+2fOFT6JzjWecgQmg/
M3M4X5u3mb/0sU2lXtWZOeU82SJtSXNZS7Ba/a9ok/SNbGRqkSKSyic8kLvi9o7p
baY0Z4ngNg4ZJfkUM30FIWh/bHP2px5Y2LcKkl4BhQ2jg2Yb+VCf4v3qqIExqmAD
Z6skkrI7Edfo1kcUCSObD/U1DUuEg++Lb9vhQwI/pSoGV0GHcnaPGrHJqbLHI4bl
sw4B+mqcFO8c3XTOcWKV7VCY/YEtQRRXRT2WZrgI9cjfX7YWCTL0/WdQkzlN29I9
s4YvzIW0iMUOYMKvktsD3u9p80zvJ3abUWB8xh0WT4Cw6vGJPNVNwIpe7mRd4sml
RcBFymRn+o2wB21o7D+DkglyOoHcCzy6Bwmb4N6/zXFaszskW6NS1RLQ6R3mIb6A
PpWw68wD2efYnFtM/3lSDZd16aQ8xKWRy3vbas5BZn8Nd0uYKVhTg0HzC2FTtxli
w/UQ9a0SQPvXTRe0WliqacBf9mYsB6+Q9Vuh9mwjh6LbFIz4r+jRsJKMfFur+wLa
xythnZSogJRf2OXqOreknw8AWs8Vs6w3HpPARjZbbrv3ISK7ydNiDZASL84eZrti
PmxQTfIPl7VDNX5zW0u3RYBTMXMdkmcQD2f1tZu2+d7KdeNjfqf759XwgstfT/U1
L3GHvbDwJYfswcgA1jADmHRdba1W09YF37UDKMHpaxJWx+d4DX/hrZu26C8pymS0
kTUUcuzzgCxa3DyV8auC7L3/zfIfAiBKvWB8hP3GcsZW7pVhDa/w2RJzFOsllu3L
706tUyCq98J4kizeTXaXSZGO+oGRawX5BJ9MwmU6mnepgHXdzkHF6mfrmlFakgRn
cEBdKJHW6bBHt3AZSuwLI+Z1Jy4p8jNRo60IVODAof2xaOsuaa2DzAN5JSTC4qpz
A/tueiOR5SJJu+MVGm0LSU1RDH0YoVdlrQCTzHgsIuLPWYFSHq6cxejA4b0YzHPI
H5DEL6K6OJK7+B1tAIVT01WNXtxOxz5UBIY1UEcRNIYvmJeeiyelZm62lr/+hbXY
3eLKSjgM5ri03clCDV+lFErsCqHOAn44W+NYNv9C18/fRy5igIHPvy0uaAqMSu3P
Uyn1y/BGZotAeJvMtRWPdyTkGM1yLyETyu9f73Fki76E1XAV4zShZ4nvL5rMmP6Q
RsI4W0Iyn4Hcsuy/1PLuvzTtKKBgv9hjwle9rtwEdBZAQ86gxRsiH62AjGZQo6Qe
ThD3Ou1iY0xAn7DX4qhByJ1MNMPcc6g1NIhuBX0Y3uruJu96UP3xOn8pKHczzwiG
VH3mRPmuGQOWzOQHf1s7EvhZDsfhfWC+YrU28sPKW3UD6SFgIr644OY/U294OP5s
XvGX0aTsBNUTyZPglmuZ60CcesVbFUENVbxK4irSfh+8vIXJ5b4lIkPgQp4iB/T2
ejYqThScwBsDhwvdZL495iwCUS7N5Xt6YwEZStgKPyvhQBdMN1FbqCMSpNTCSzcp
ixRhTuVtTOgMvUqpkV6YXzl9FtdYYD2kQ7tgRHCI8xJ4d9E2XuoCp0Cg7hkGM1nO
UDH86hUH3HfK0LfYYqajWWRGWljIQ+0k6ihKvFgxVtdD0/I8hFgnwoj48V4jjRTF
pzzyNIuMw8/EvSDAvkLyYI0CxSPWJWxzLHW4F6dXgY9EGx6bhfBW59dsaa0pgz7q
UwvF1FyCiexSZHNpLohgEf+uMQsA5IkTMkblYAqsSV5VFADGcMQLgReYaz2ivPXA
3yvJ6J3tD1KFfIoBpNUKpBGoBAMmx2RqB9W+tMob1pKmiEFjA8oe1UIY1NtXS/1L
msCxEnLY1zh7V/5ROs7nAKWRskFkqzsLART2Kz8S/B/jIenVAw94U4xzRdO/GJGc
Synw+6/g1qX4LuiS85Byml5lIC3HUwqVk0bQMrC0LoVaHha8PHaNUXfR91zim9ap
yqrK87l8m9LvaAc5j1jurexwFq0yXPaswdP8W0gry2pBy4jZz8m+Fl6xb6D8rGbd
GFLJAqpXVWKjYrS3F4qlDTO7aEh4LkG/rA1ZoKv2HrjZ6TJ+Bx3hcedbMEmWHMAA
utnD/T7h64IksH6aS8L27TgvejG9HmUyxRknI3UwBCMgI0WHYw6D+NIQnFWBX87N
wBJ5yQL6K1AZIMh+oUXAMgtfF8FiNzozZN6Tzi208ihHfIpdQyCZX1Xz2F3+GE4p
KEoG4SnODCmTy6l686A0/HTTBL+AqfJETHgkgVY6UGdljIjJtUXihmIX2XGLvHz5
RbrhXAKDK88IqTONulGcbyBuyO5feG071vK6vQ9q08dKpsNeweOavJIzYj9sN3PY
yModLkccQQZ4gcC5no/ODwbM90vcaAWW5hhvE1VQn9cFYhe77b7uditzRhzqDNz7
JwT3jxdlgRNJimTvkQT71yvLnyAlI8YGE4Pu6AoUUxseL5SL//XMtVH2He/DXN64
HHFfPLh4uuqhyHOy/xq41eGofF5ZW8gkItXqPTCHcf5hpMD3cicgvJW4PcrWIbMb
Vu0gS/Q8pqVNIOaE86KJtAQV/Bj4yORKimfNtpFiITSUUtzBw/iIhTPsk1dYPb1g
+9YfJaDGfYxlpYyWavApmeZEiasLkUagFmM9XndqikCHIdawzyhPh7dDpIomPMxa
Ls2pfYW0NUYF4wQbBpQOT7DvMPc+qy8my4+9M6llo0e24AM5xlHFzkQgLtJHhwZU
xcc7NXkcnEhu0eu4ulyNYNZJ8Ln6ABgJA9zFh9fCApPH5BwqeX6ij4jU+K3BK7fO
uuU+Osazz8l7IsM2zwS7qJ/OqQo4WQl3xmO4e6OusyonJhuu8DTGiLxPjIno9SLq
KnNkDKH6FyuTSSC31eJymImEm30MPeGhj1doSzxeqOJXe9xjha2TnF9Zs13SQndM
flyLeE0MaekZ3FPbBKCP5tM1MVZAGkNThJ/4hdb49fQE5RBpn+Ey0dwdDA9Wiha4
HKeIjlUAWs+BF4Qt7MYCXBPR352bp+9w7uwy9/R3Nwc7XrHtzgrzxpkd1Ssizz1Q
8OGMEnU1hAr/m1VSsM4nhCNE7DaQsivjPKF+0AlhKGKsAG9HpHFfLSHDHjuG49vA
U4jF/MTsVZu6eYXo77bLwAOoGQuwCnZjIh88CpxocirDM0Ru9b/cQzwyIopHABsO
bf3C0X+tXSD29Qc+0e3Krx541X0nCWOjxrWrgPxwPf5tQ58ohnc/yKl81RsbzYUw
P/RM7PBILxqQ6nCbFhfwaF1YshPUNxJF5DJsFLSUrwxp77MZSrMZet5/Uce06uxj
cQx28ZsIB9jd9+CxZHTaE719NBSuxAdtI0eh5vsaqumClRVDbc3xIQQ4mw+Ekzzx
qpTsiUyuSBaKJW7zAQIDmm6Zx6/+PIkxPizaRP2/Rdg1wKtUz9pu50T1aW3O7U13
49KM81HIMiKXLFy3IWASIi9y+G/hgt1sVEIxBnO4rYkFez7e/Nr3aTK9SKn8giSp
h7wWw1c/y00wxjDk3KF0n1071BS7R7oGgMSndLNTYf6L+RJ+4HY5+rIFSDqJeUd6
0Ud0A83f6acSA0quJBU8DxyRrsSUiw6FU8pEK5uolukiASU3288LxufPBlUN/m0F
ioZkvjl2pznXDns5l1aSmZa+RHWwzE9P9P8YhovAOkE6/E7T1isBrFrN0FZHZMYN
dHhFqPCnpPOLsb6U5lCKzNcbFN5oktWjoacouHy2i62ZEutIjpYIvpVuvzTXaJsS
j1Hfoizhd+oJt0sO7z6bvhssD3mXgxNovNLikHuwbta/hLk2wb6Jv/OcyNX61mPO
aZLiwWMxZjGHK7HElZbSAldUj+xizdrWYEHSgMgE+ADCr9IND3YvA3NZ+JTSNU9Q
6F4f72O57a8+lvlF5wMItJQflStTSELeKGTlx5JsbS8Gi7z89koXC1W7tH4Aogh2
cbEqLFkcl6LPjY2WzU3/odI92KzTnWwvOqGaaXTb2Eflr+MZd+fyRHG4TpjnctrZ
UmbyPgKpaBfyqjFxmTO5hvBcqXTIcSOi2cVeoYEzDdIkDR436oAGKJR7fvMQtJ17
qW+QEUnS14rQjM38k/zbQbTqGbNqw/wSIIk6+LLDOwu1KGcN+qJRjm9a1rrddPio
U5Hbg6Y2nGlFx2IdNBmEFsEGqG09WsrD/wC/BJlcqs6aBj81vsq+AJiEJ2bxC7YB
UzFGHa1HHPbG4+4GnAdzEZPgaJTEardmvE2N9waXAcoAUh9wbFopabv2cSl1Tn3j
5ZuRF461caAvmab+KnnN3Xbm1gW/blEsr3YOM4xB5o+Dlf+HN+FPO3wFsSpmk5oi
wIBUWwta/fslrhporr4b6viterihgreCi/P83g0uF/g2aUTc69mINX+boXSvzMNB
LlOAARxUWWUGvpNjI/BonOtsZRcEOvJcR/nvyDgZSnENq9ui4YchyQToZ1ZCq6g9
cwoC6DfmuM3pq5aXgPtXltV/eoWKgBz8w/OizI/GRgUS6vSP8XjyGq8brt3rG+mw
tZRwswhQCOYopyl1qvxY3XnXRJcj9jdGwdZmx2IqvqKiqWVP7A5A8AbOfPqRbUQA
1cpGNZv8fbXQi0UfK99/is/b5XZCv0pgmW45nSP6HLm9JphMB6RbBKYQdw/j8BNp
HGKT415crSDH0nBlsB5CNkH65xKUlxPgFRCfEs0km/nzVQX2uGgZiL99hly30MjA
5ckgRG1sF7QY46rgfgWMULpKAQUqRVL50s4umfqY1OxC81zEjK89NDnrpuhINf0L
JqRAIw4/Izac3dpydUJA/SjCFsph0vCry3/SVI0IimcEHwCtOwLlKmSAzbuMuQ5J
L3GYIFJbIgTePVzz57xkWCvU1b+9nClcKDmS7JcCUf8ayTBdZBYRfgXu244Rh0zo
1WiFBtZ/+7BHUlWuutXzf4P3MAkXvhDX8wtbgqHWh1dyp5R208UMNCgP57DNHw97
NchPi/evNReSNqrjCY/gV4ht5qbRvf3blwY3UrFeh5ePRPC+ftrs23ed0GL8tEYD
j1RCCDoPgp5BA9OVuiliZRBxA13vVNjoUB0GV7D5t/BKdAIN7j844W0lyeOJ942O
8dOfMbTBM63qqNB0p4QE0FMA+l0MhuDOPvQj+WTAy541cfbcesfElkKzzUXURAxl
9+tZrFZaIFj9p0jOR3CguoFJio56s2dgKN5H4G2UJMjnAMCwQZRl3FRqXnDtT6oh
+BLdkud+XITDZbfQXDQoFBAI+Q5GNto/esC/4aojCXQb08qbp8ada4nqcYXc4PHn
aFSWEt/BJQIQTNwXA7HBMZI7rL1tiEJFbjf6lfAEqojhnjnQUWaRTpd7oBV0+pxO
vGUzEOaBOlI3Zq3FGSffmxwD7gzVUELbgdSHOGpoofnSf3pChMDyRGtxKRYStRz0
VMvCkAC0d+O9k/z4PM2Ok8qOUiBLGavnH9rorsUiTUDqT1E3eiyjyeGNyDDxp4kM
9c3Mdvu0BR6kNhlFtbEHgrfBZvwbhxzi8H+h2Nh+YQmtkNaUoL9nTZp1s0RKup0G
dOF67ORR9qFszCtIsWH4yJGWEnsJfVXPbid0HcYpbjLRxvNvM7zRAnXPa1962JAx
alBI7kESOEqVi2YO7RuJ6MkivwclIT1dum88OxqTyNZtQ9gbfkVdkb4Kq8SwfhDO
i1Wz8dDQmvhNV+fjyds3+4axC3eEB5IkM4myxAI6OAvCG79ziWIdxLAm+fUpAczN
MPwzzolVBnKJHeZwZRM1ITHin/Q+ZUXocV6rk90Q8TlqYTznWcK7njpDXEBzr5qE
w2SglFQfgn3uakp4pNK9giTBaO3LICVby450BY4nT5f7swMxyS2O7X45r8uMfiPR
khf3xd8//QHJGrKZ75hvbWEZjETFKEPpz3RBWUjOnDGzLyoPSHtgaANIb6c7sSpO
Md2Y91yDeQTbP5fIg5BP+2yxrc5Uveku/0czAqKRrOqdIwuhU0ebvva0jmmQEJzQ
Zgt+PGP6ugin8srHUuuTVrF5ol1T4G86aoyoc/VjTKpDh5nsaoi+Ga4ZFtDl0Wn9
3UIwQOYgt12vtAwF/M1fAxqBfBhAdn/uXfWupK53Cx8Wuk8WRsowuwiD8gTmvtQS
lct638n+eBOumy09gsQsbHB+MsmG4rI1twIPrQ/RNNuey/1ejtdYmdlSxQVbA3Ym
qGW6nLQDufwAVW/hPB8yvcAyMer5awupL2LZbJ5gliikkNWRNeTDQUjh3AYbd495
fYzUpmQPKlCAJNvBV4FMxJPpermvpXWYOr4yQjW7UBCjTTTON43Zo/DXtfCbbwLS
w4s+S/YcVo3owGyRZPL8f9fpmxi+H4BE6hR2oDEXzseelY5C0q9tGCHHTAwp+1jz
nSgpndfeLwEA4/7haiqLrdcQRj1o9uJLl2XfIsYGSJkXdyZBhh1x1CKhHSG/o0aK
rZzF54ltPRG42URS0bg7Swn9v/i4AYbgT9CkcPNADDu4QSVv/eXEmf5uj4Ks6ogo
AgMOOTKfxAesnm3iz6l3t6Xc5COAf2mlEaEY+/+avnBDmI837NfBmGqucVpBo9Wa
xytBJ3JhPs4WI+GDNyQGaCPBk5fylL7xTF4wxpSvdvJ8WhtWwAbsbVddcK0Z3iXw
/nsJ5NNfSVay2gaiYi8cC17YSjB+VWYmAxVHwMogukBIGGE9dLh8g9hIje9qFMsS
Q2CGD4VYEsPY7qYrMjP6Efct8FnxYGcw6DN9B3Lh1vpP0M+xsQPZ97Psdd2lCDaR
yS/8FbxBdrMX36Z+Z/P+nUBBKnfA8F0i87MZOHBPjpwr/iSDUebWKwidZcHFHaFj
Dc/+GKMqSJcmKc4szdSESRvw//gVsepqR6if515WiBWqhZuZYLp+u4umpIKlyJqK
zsFaI/RJOLwmjWmBhHN2JuKvFTj5mrn//A/At9MPFKOYFj4jwUlO1YnA3LTc/Xsw
vGRpcBOmzr+/X8474XWae/iPSGNAcbuUFmq36o8RnaAqQ2i9K2vJVTga9c8PWjZ2
SI+04ZRslZ24tlIUTx32KyxPHwgCSa1Bs9IeBMtfs1vqtWgaOW24yUJ3+r8mPafK
vTZ3VH5JnQW9zu0Wfk15vqQLwGKVdJXetKXOOnZbm/2iu7zDTpUJNpdz/Z9BPQxj
bQjOnrIc908gsWmojtxnXhuzGLbrFab5LORh8CU+hcwskiFgWArOsc0pVIDjYMHE
eGR6RF8FjEm8i1OKa9cIV5WWsHcKcG4F9lmsFH/pEKvRey7DMzv3vvKnMwJzB4Ht
lLRlXzuhjJaH/sgciqM9jYLa67sEBDrDgJVFGAEKwRLx/16/NOImFd7Bxhkdkxbu
ugHFQzw4gANRns43OIEjSmTSn5j4bUJMT36tr5m5UvZajLnXZeFfyDMy4L6h8mf/
lLl3IOsw18nQBkLHnESTWH8/UoWYQvE1yyDbgPLL8rPsbuKGaN38KHAsog0AtY1G
/HzBfrlMSlZnkcaw0WehFx4/rbecmX9/I9maJVaKWCWfs+r56YefK2rne+72rpPJ
X6DleWKEZ4I1XIcDGP7UASnd63R6ziN8pSZQ5KM9suLFwrEkOY8Icbev+Pkt6LzT
QwQzyNC29V8Q/+uX/Otio+7eoqR3MmJWSkN1kUtXiODYMifJPBS8xzTU9W6x7wrE
dazkqio7r9ryV4vzt96tli5kyz9v3lSAT0qBD1mLccWYh7gwIMM0HmZSHbxGB+bi
NGrnKZnWzOxC/8m85fh2XUGYOrV4VmtMUMwh6nb3TPcXCIz+QZn4GLvDzf4yULnj
T7efswYnj8bTb8ZZjprAr2iwhx6yT45CSuJc0fGW25LdpFSN2d4vi582BNH0cY5C
UvKO3WDLjsT+OPLed1psk8qE+4ZlC679OwMCRbBiZj9OB9CO09llH0w1bQRlRpqz
U0YMtjvAvgckiESI66KPEGUuQKJ0FANLomHWB+FW8W6TwYcF5kvhGVXZcfUJmE2Y
3LPa/hK8ubVI+LEfkwGbWhpheFHf69xeoe2kptSATXlm122LS2WuBcQ8zRgBPKYv
iCjalgOP7rBMDPFt/wH51KPSqzbjIvT2tUyTdPk6GpNryxgbVEAVsBSIk/EkBljs
0MK925j1S4700CQEs8OMhlAak0sV+1hHOBe4oVo0lrx1yjjFIZWQCD3Fjb6meXof
AM1LnjgD8jRlrqqTxRq8HTthmw4r4yQ0W+mnXNL92RyTTWP58jkLGFdJ8z4a84BM
5pAngQ1xAWfIL4JQilICblkLqKaPenB8KvdeYHFII2eIWRJKJGIOs8f2WJN+wd5W
avoN8NFiLXvbKHhT4TzcL5pT7F3/OMy3x3746pcCB2mQLAnu/xrRKPiviorsrCAI
6SeFaqfH3nV1eCQT7kFHX1ewz7gKfiLMVkve8Awjq1ZnpDkt5ChhMJz+LRP//Krc
klFIs4PxbM8MqAFNKS9DACY3b8rsCy4BJrff0lxmmqixGQE+Q6AuDOFPCb3lKDzj
vhgmAMigzAm/eIKI8+VOKh82yTIDtYB1XC/4p4+tdz53MxBH4fSVAxvkXzCtoaZK
+XBEzNeKGzjEv3i8VVQZkeCHOUAvCRIMR6ML7usWiqa4H0I12RBNGZPa1dyjujhE
yzhnTItSLxWUzjBf0w4E2iN8BFg3x/hrKLOKPMIswOaSEj4lz7qmyeohjp6NsuWO
qID2EtZHcy3c21BqcE7NfH0i5zZteVQzbqdEbg3VA8sraetO8HnOVqc+Vaa7Ofvj
zhmrKum1nDUEyVkF7ZYGn2Get2XquZojDrd+fFv6BvbifgWc15KVdFxe/W7mQn4V
A9GJzgVI9AUeupBsLLqcu5YAjunqlarlrZQrn5ZtrxmhN0TwjpSqxG67wbn8oBCt
A1Ug3xuAnIzc1pMJ+qiPNc9Deq7IzvJ1UyW9R7TvLFBVowrlyVxU2m7UtSqRETZ4
ERK2WnrtvF/xpc3cRjfsweHzh1DR9oDqA7iO5DcKmz+QWk1OaSAn5QuOU41AKOHE
odZWZAVnDF9Fiw9fZgepYlNJDG2Ew5s6IOsu5gCZX33cymwWNneibVZy22ynNkUm
zeQ/nwZKbr3GJKKymmkIF4sopH4gLnsqio8SsLlQ0EGhKtRqjDhuwzIsvg/2nc7D
esuF1btOH+4hEm6C/6/WYJXhwYVWpgM4tHh18CV7HPIe34HcrEkSgUk0byQROfLC
7S5vqC34py9Z1w0/Pj4QO2Byu5Mo5othdcFxSf1PF4SHnXEP0uSZRN1Lo/Jx0LhE
605GPtqv31SY2utApL9rEpRuclSO/nklzZ2fkjMx7dFfWhHFmHu2GR77LWKnzsIE
bAtW0RWTSIfs/Fym4Dv1Qrqj8TVHue/5T/6oAOMmNgP+pptKnuUY6Pb/jeT0oOK4
dNoJkXYMrSnvT3Ch6jUOaokp8vFSeHDM8WhKGXVqsHJZm2KVliUOdG28hzTS2edC
RVD3GfZp3MpKsoOxuYpckvbdnyYJqOIyao92rT9j+wAtxVTn8fmdwOgS+o4NkqTF
CGZB4X70YTJqMjwp2csfJXZwXiMe84ZHhAgkLsaGqrEQ4MrAKhFEqpGrSQLxhcoE
yra1oYR8V+CaCmXMJ14xVJoICF40m64O9yzWqIBbfY3tBjNxt7Zbf1SUb7+aYr+Q
bmavWI+hVVHjiFyre/O0TQKHP+U44dXZ/L+EBuKQFISPHcq7BOsBaFmT6CisrWNF
Dgmb3KLXIr7fC5WL/w5BUmNdDY+pe1Vg+C58tMMiQO4=
`protect END_PROTECTED
