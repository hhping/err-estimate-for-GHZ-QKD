`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcX9sjvA2cEdFaSv7DH1G68vGgfQ1UMsHN8plUA54je6+uvV+se+OaddbZjtvvj3
BXCeWU4YdIZIX4FIuXId9tmbpca0braD1z6uaAXD0osydeO1HUvqpL2VrHwvztKG
4Yx0P1xw/nltFvB10++oYI2UM6e4f30OntHefSjz2j+t0y9ymmYa/coiQPeRr7mN
04i7yIRLLa3hCYmneBfgEKotPo1bbPCGh/1mVj1JADm/bMXaR5nfBRUfOWxoz3La
Q0p+4LaeeV3RUEg+jxRAdW9U5HHMNJYx49U6LYH3RbsXNAx0UR8FebSSFuzqJRnD
5hwf8/0AORS5F8a7xOJBXE052kWnMPOCyRk29iXADZTGTFiu9zvpMEakhPGFs3YQ
8o+RSWB68kSuM49Ui608depMducofOK12XZkUMKcnpQkcpILqSG199LV8tkbpMON
F5ufz5lT51qnZOgUejDDXgRbG0AWt2vQjrMx6AH1CimT0NXsAG1BTOdCCj/BaY32
F4XyOE6EznG1L48GRlNUa+finUXLH5MS2sHntBZoKd46/yaVY6VY4Eq+1Fkl3/wF
po+pgSpyqKiGOgKPtoSCjBFTqo6Y8WhbEWcWAJZWzAvYlpnS2ybvztiV0SFfXQAn
IY+u8qnpbGjik3oSqmLtTs4z3BvJ1mPvT2DGNG6h8O5L3K/FCsSxowRtELs5pYxp
ugTHDe2jrAdyk/ve9WXS05NplxjAoc4Mf1sQEi91EBg4ieqlXI1SUA9kNEKZmdJZ
YzjhB2NhVO2FWLIAO5Rtv11XfZBL71zbEPgB04qJOXu7G87dUvRrJN+ibxAA9X+o
Uqnafo988nHa3rF7ONWztsg+gxLagMEDFHrP9HjbsZCNAHs8QmXAnW88KTxZIyLC
boMzop8e836f+fo15njM3ioed7jLEcTRdXn9y1AvJ6rrHuloPGgzp6cTgb/La78W
jexOZPhagurRNQoRwrnv4PqOJx8B6HaP2OAEDgQ2ORDsZKTVK5p0NA0VcKJ73qpD
DVzxkqkYhx55iCaPI2G30/85llcEivLA+omt6ntYtqbOlgqo4Z3uSdR1VVKBEwm8
RSRM7XdW/jmL09x+8xqdnQGGENJs01nyC4q8pH4fl0f4D50t2igglK1e0Z9BiR6H
fAnRQidCGWGA1Nh9Aoi+of4ath1w7zUR0ljyd1BZZXKgycPe0S8HOfpWJ+rGa2IO
5VspSeFrHs7ya4ZwILQkxaYTm7k+mnXrZAN+27d6C4BXWpskYMH1j06rhsjoVVpq
bZZEhNQfKwu3/HHmk1FSCHiXCHv8j3xg3+wFk21a5SR7tfdUtJch35ympQRzUPbA
`protect END_PROTECTED
