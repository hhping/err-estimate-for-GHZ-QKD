`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqm4C4Sduc3xtd3zaYzQGFLjakwWHw46NCzioLKp0IqMEmZXHr7cMtj37K8YuiBY
jPjbXmsvKBOkh6c1Rm4G49ME/ZyTotJD76YmxUyXjUqMT7yZWsrsAjErnLFYRlac
lFB+atTciOkw2D5QUofHEPqXNR3RgUnUGbe5JpXEk391XT8f6YPNjoq2exELXTo1
w13/z3FDLEJ+OVQrJ1w4rwYjgCO22JwdJb7PJJy7oq3hAUuVz4OWFrco4lp6D/SJ
41tIAswHR3h/Amepj5jMSvjInOKHBQRnHfnnVgRkDjW23xHRcD1ND7hP0Ffh57CA
aTKV8Lnz1TAtvdkdpH3/OFACuTWZ5X7DPEsVagnTjGo4+HX8C9GD9k11CFLGqzJt
sW/pS9OFHQeBH/YbQVKgv6y3iFW3w7JL3J1C3W1PgUW4BDRJEvcUOYM2Aod2qWX7
Md4pCnbBC42iFq/p9GjVoOGvqD46azbAstRfRnG2+4Mp/o0qUXKmmqjs+r4WbeqS
REQ53e5LdaH0MEK3Bm6GqgJhmTxhG5goMgjFgPEKIkWdM3N389KJYbujnx8dX+HN
CDGkzH7uMaQCmXuHCnlUZsOtGbhrvWoEe+exnRDIkN+pVWZtU4RhNq5XYp5RurFv
hM0X1OL3UVm24qc+rmZ4GGUISiwm+LebE0OOigvtiRtTHMnZsEKZfot5ye/F4yx2
es+ThzhNGaZTnQQHykW8RHUfz8SlkyG+MVRHnj45gjrLSzbHPDv8EDwjxUQUFclE
L35YHHArV53UYYVHmRSTtNQXfdxJHCswZoDbgoiirSYLods/l4O4hxe27bYkZdut
GRFoDdN2AJRAAxrR1ZM2dSh56FbxdRwRttYhGghIjfFidTI7epw/Z8/MNCXNEsM+
rgexZ791WfV+kAVGaowA7j715Mi4gmls1j6gZu2d3zQYVKiikiA+eEYfLgvk9j2R
m6zOuTAhI3jFQCk0Rkf6Te6SS9lvFtNbYbEDpu3fP5eboeBSi8hed8UEcNYOBmaU
p44pmelGTgcRjuY6f1YpSKY3OJR/SoEVTAIdt+XkAhrdhGDgOVdMYTLRv9b1MfsX
NyD5W0H4V8j54iVh4uo95jn+1x1eFIea8RTnCDiToVO6DXrjTqsZO6IRIE1IeKjs
K+cYpmt3lDR+DhXisw2BO1upnFbQHyC3pfxMDTf/yPrephY/bnINZk60dzB/b3J8
+Jr03dp30/R/FMtq/NtzhxABclqg2mLaK3+MVNjqcSHzz2qxb2Wq2kzdJ7YKhxwo
s6md7KEjNLAi0W6WIHQnTsgFW9PzUn1MFEB53XVp0pA2xXLh15/0Vqj+0e3HLbpA
McIGpzU+3ldOeFeD50QJsysabfgkvyceGl/Hk9n7i2pbJdDIC0vcUg22WhrCsDLO
NgmyWXtAZLELjln4t8URK+V27nU8K/IhR3q/83BR+lo8gk6DYm51hQYXDDvZVcXb
sHYxs3pzEHXnpiSj4JdUqP7av51Ch8tZb1cS3XDfQ6Chd5sVe1QHtJViYK8Gg2ev
WZCxpyB9uNmJOQy1/dUMth/iP4LZwWL/gJjvTZ6O7J7S5LCJt1LhRYtuiwkqFIpb
FXA17r6uhOtthiFJUcmal1NGOvtA0vso9zqFNoZIuvFmNteuj/lKhxmvp7YDzSpb
xXe/ZVI00wkVGID7ybv2YA5PJFGJzmWEyVTBVIMCe/qzBiAKRC2ecqPLGYfiHIH/
yhKcl9wVFHbhNJvma1/Op+Hj6hHCyYG3ec9cFeOlY0YyBUejzEQpr/pRX/ikrnJB
ZKmH4HbFnwHVAP6PXIHEjhiVj8FAmEFssMtroTuxVlYCW+SQuLtoVX+UiiBE7ClY
OI48ccazfZMi0xHlwNdoXtZszqtylUmPupgoEnkmCyyruRl6N8+DdIh0jgbUFHPQ
+hl/Ye8S8ZDh1tjmf99SRS4q7sbq1OyDnnUyOpVrVK6pVXIjNFabvtAC64dkYzP4
w6yJYqhUplwOzEc1YgR2MNQxrANFrN8cciPtpo9AtsA1f4pwkIeirMXOGrqFopLL
cuo0de2VTSFihzqsWOqI9O08d9kPAD+JTRO3/D+oqmriMlMRRCwCjsLDEcaS2Fqf
ETxtwamgySSMxL1A+AfhJaJ9gO1Dhyhnqg3L9NX05IjnQ7OUlgazufnO53mN1DFI
lqhQ+AC+mOWau76MFcGW1sTGs6pE7ebt4ovdIxYfyDCExwN9urwmyxQmT+GkNsPw
KMv2+/Oyw2q+f5jg7vy4Oj3xDRGGF5cjB+95hEZelF2khYFTUi9qQpUsYoEI6ifM
K+cRL9PznoMmV9rVCmvzTQoOxSsQQiZV4BikkionEuw+gx2n56oIs1ITfJ2U7l/D
c14YRQ3LAKs8/9LCu3WoFku9mwtS5Hc1XVasiMGHyVr98C/0NmPI1Hm10odnc/h6
olfKQLuLCSpB1i5ARJx+LEjtjA0K1GZNHEigD6i3gflvUBW1Js0ZncFQM/B0Af9f
9LKHL+F7wTNWazUbn0CThOlgGsK/BpikDb7/bX/vtLIl4dc/AAQL42NflNgB8uBO
aZ1DaXJox5EBIbO9ZeM4VMdUdaUGvyK+272pY3SflQ1p4L/rKMJo4sDwvrUYkgd4
0k1IGxs9fosdcvE3SEHiG80j3G8cfz5Kr1WZRSN1qH+io7ZKMn/32D48hXKcnxV+
ierCY4o++audYuCig9o7qw==
`protect END_PROTECTED
