`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvcHURJBaTfRdFl63K870V+3VWq9rwC2j7LH39jCa/t5Qb4HbmBLtPqjU7+GRtXm
RWgL5om6XI5F/1wIhAMJNcrClk1ozSZoB/moqzg+KYAkO+3sru/pNnzxuZJuq5bZ
fFV5bxFTkfvPh3Ftl98Q1wgC2WfNxWByvzy8bmxuVVWIgwq8l+SYLZxyE2CKogH6
HgU8y/CMcIlJpIDjEbil5prwlBR0gpKOcvJ2hMRmD6pmVEJnC5Tj1iDYS7bweBHE
k9NR337bSSZaqekmWCen4I9oLzAJS8qq5HiuE4Wr60EkHe8GE7cbuU5haH1Ih30U
oduzkF0ePtDKOVxou+koElCnYu/uZO9BUx0L9z5eJbjlp8oHgbf4URdPi6e9SVh7
8cnVZqVZrowIwa3bN2uEmqExNQ/vrH7IfVE/Ix89NkdBv0XhwfcwKR2j5vgT11mO
HHk+9X3MakpRLvjm65ywOXonXhkvP72ICSWfNShCuua4wGpplsOESZVAr2zWHu5M
/zV0ngKisxkSWyfXM4+QGm5QI0g1fENY5vsI735M3588UjKTBjlEujJ/7GV+EWAh
+onB3GWZ6mWXAeimLpXCdsJb6L/xDAo4adrmiznvQO94Scruhot5b5V8i3jO8DIW
IVde6lFhajdfGN38kcNguyuMD0izS0RcSQc5erygb/93M9Y54fkBbtk3AxsBZQaG
9DXctw6xqAwrsUSuM7frjmtv+9AQJPMiEY3HIOtdehhDMwnV+ldywVj0w5pTYZJ3
UNRJGcZOC/mmpA1kw7hLibYJVmGi72xSJhTpjYNw3JOZzzNsr+dbvAMmVX8ZQybD
EMbs8G5z/uxTKmTI/A6aSWDZrdIa3rAj8j4mMtrlQaPaA8L+PejUkqCrpUGeglQb
mIZPKlhFUMnBiAV7IEzwv42L/e2t+Y5yMhwma6YCiQUoWuB5Vj1wxs0N0dgdiCw0
CDNbplXYKc23LZInG93qOFNMTwdr18IN5NvvpDh84Wd9cVil+ys0Ehhd1clnZi0/
j8eS6DhBa26gO9A74eEfn9qz7i0nycYHoC2mJ63mdHr4cXvhGOscLHCEhZl1alb5
tjXYy/RmPgpTyzwGGY+f2ofpgN97DthgQziY44JfkP/io94qBvI+UXTLgQtq+56x
gmx01/CgwIwg1g4JSD3xDPFVHaogUv0lgGFjdBsxF/HKRn/jjfG0zOLjmaQtLsKt
bOZQkFDhQ2pbN35RyX/t9iciUNUy/xy0zlqxLvaxdZTIFrTCZwR2VRTdgH3ypUGo
n40CBs5JsO5okrpckdN+v5cBlA7yzSvdYgZ5XpQOZ5JrfqFIZKaE6k+96v1XEW6/
/DR67E/EEVXx1K+BFgmFADg1d1GwTkzaEIn1aF1rNkVyohloemMDjzA+amqWwkvF
JrLlMjK9zIce+G1KrKYRP6caQ/u0e7OlulJdyjPFddMfw34QF7x5I/RLrDGBLxnu
iroA4pZJG83PsllZA3a64H6UJ3tApMAiik/fR5McYMri6O9mJgWom2/h8rdNfGON
NHJVhMCD/Fs5Iwp4ksDK/uitY5orAxtR2J4+TmMtkDnp4c0N2+SVbgZ2eohHgKzi
dJV3x6K1PypwPSe7ipZ5dcJq9Ia6BL03r6tQFFRwM3ysEhX2tAKWEsjHzuG9tN4K
D7v2FtNQVI7GOPfZNCLPsIP1JZTkqF+PShM+D7MxzTHX6LhkhSEAZA3t6eGE1VXy
mHLLz0hCmmv8g4f46C4CeABTEJ5Tpd8aKetXKqa4QdKxnHZgwn3zOp0w5lVnDAo8
+49Js5nB5p3lnp6FaMkwLlRfko+Bm1iN4HXYhiEVYRKfIkrQNH7SSomr+hSY7Eyx
t4EGG9p6WavSTdvH2H/vDQ==
`protect END_PROTECTED
