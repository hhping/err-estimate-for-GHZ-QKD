`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbA/rqbxrT4xlJqEkuHY4Ye62BjUJ3jE2uDrEgg9H+34k7G387/i7fmNZWfoe3KR
zc5tgeds8YCDuFesn+YZX9JEMwh+HlLAqAcHaI0cz9SMyRKhOyFifnG3xChnOGM8
rg2gzjfUvx37ynnflgHT5qRX454ZYr1xcBXy/4G5a7VSHo9CnfGeXu2f7wgpYYTK
wCjpHEwVGgFiun85E/p8wwyaEvKl5nY9EoND1guvGdwnuBce+B8s5gNPzd4+DxPi
S+VozUDgIHXX8LzNcgtekYRGG9EnEh1efEW2wzXsipnqWC8RUKNH993AAO/JBG2l
GCAdXXeFP5J4lxfS7nZpWzFBh2J3stKlOUhzVSLzZh7sIWHQHQhCEWVWx/qDyzGP
C19z0H1xhS2qKRXWXuKnF6eyeESq/aDWLlorPXw4T3jerI7GX2mJ0Fhj36MgQvjJ
chC86HHwHJFMCRf4XouabZVYX7sc07R5QcftTlTSSXGEqG5Kj6yOc3E4k9ofX5B6
L2ZNVBQBF1/WDNTYr02+7QllYnK7ieTCYWy2p214ZSP3CvfnOcRw+01kRRNrWzaS
`protect END_PROTECTED
