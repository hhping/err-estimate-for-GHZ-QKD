`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
66+IhVG8WKUgZUwlgp406ulC84X0rF11HTrjtc+KEHygKm/oFy9TI9BPQZxiwzOc
pVEyAwi8e0LGhhXHy55jsPWcWDdrA80vky+Dd9zOIdAT6+apW0QW7WhdGbQxGtf0
7+vFglI9NPyk1WQ+OExFe35UEDpK0BTIs0li/sY8wW4xI2GxAxYnB/mWa5RhRNY7
5tkJz7q97KzcndjN2ciIlTPEJcLq2BWhs8UyBYN9RA1hQgq1cf6gnIZrxSIE8uy3
lKVh6E5PU3kT3LNEMLALQVdl5pVYnVxl79LzfsRSdMLkM4ESRoVR9fKarlIKGqLU
MLNYvGgPZCKa7AbOH9tc6zI58tWWcU4+XByEwUSjmvYZrS2HeLiOXIvZXKPCaUxe
ZPAL+VqVeW41Espey+aaaBQZf2rC/4YewkasZ1I5fpd6LzzrRJe5fUXb9ZsZtW6f
CLuWOT+K1cAW7D5f4UW5R8ZD0A1JvUzRGLKBfRdcp26wklyu9tiWC7CQYzAFpccf
g8Yre8mEjJBNJb/pY8fyyauWDWILQW8VH8kJStWBs9BrF2C7H7w16mxMTBoc1/QO
vfHu12BLovoXpNMTLmEaO4jkKvrzrBn2TZVMiqknnkeAD7aef4McOJ83u1HZzaTs
3uqH+Ag+R883P5+a7xLPlhRpX4bKEBngKM1HDo3Js2GS7XNcNnVs7iiba78TQKwF
kxq+M65nJl81DX5qS1TxOFxyfobUiwWWd8gKhRmW03WE9tu5zNYUarEkmMmz+Zaa
7LS/w61BulHrVUMPpFk11+pTVQPx66rkXVqOldIElyrrN6lMPGrQCDaNXAKXg0eI
PpiUZn6M5gMr3ioXPHzah/iPYsX9SD+sbWEGc8jRrMFP0bXkWpFMmyXugKArhVJq
1AiRIUf/zaewwkfXtgScd9ZNn9auZ1QdZ2W6r9j9r7S6HuDbIweXRH8UD0eDo+GP
jwGYPdMmr4BlEDekBrLsbzF3wE93VFBfV/5rYhYcfZZ4PPBRnqCWXyQeL5SwTxPs
ZbKmKgO0xB6O0WXmK/SnI0I4BKaBVErnF3XSrwDpPeEgQcEEWS4os8a7nSXOJIVp
ql4dh6UXl+/Zxr+Ks+rYaunI4OxoM8RVlKxhj+ChdlJ/t6kopuXlSyQtuHNL8FuK
BvDezH3KC4XXE+duA9LeMpnqRGDEccrWK/Wcm9MLFgLGf1GSs3+hDH2Shht/Oc59
TvU6d6g8fPTXOEnqXIsfVQKGiuMa1SlkG8OU3f5I9c2R9W+nN5Ep/alLdjIqMkmj
vmPVrRMvRNw/J91/pSsC2RRtpnK8JtedidUP4xkpmhyAgqVp9WZxA38piwSX+jgH
IzHuClgOWvunUxNyePDOtjZyaEsx2C5VCE0WBVvKiiNQdE51k6ffHJ9/TI73CUR4
kxc1hOxn3rVO59+oYNMilP5HdWST42U1bAuZHzx15yBnXoU3X5pjhQPuzZSAVqUu
U5J97CBAOT8guugJiuPXGDqqaHtBVeLUr7ekPiqKrri8rxrRBxjEslBvJ5zMfyXq
tHOyjtxL9Sh4fvxfyamD4QOJbCAR/0dlfs0Fcpy4URFOtKBHjCbwmjoJ5awVNV0+
DBzglcc8Z/Nl2r87wxwqYbPRfBOzmcZ4rZdWrk7awSmN5xQCioPkGhuL8CkHE3rG
soMZG2bymB9tG1P0jBkRXogfZY2znB0K7Gx2Kb1My0DCE+++aZFL665H5qg6CvWN
gvflPwOMRGVm0kwS7hqYFSzaawwpF40Hp7EM8zVe2hCTaB6PwSuhAwgRNqoeaEld
j5dnp/2FC+RCaEcgbjKWPOyHJZyx4QWWduVnmzDBWUY8LS7J4oeGdkXUimnJbKB3
TX9WloKwgffZF108/lVDNxMTBASogdttqB7nha63vkHJGU/tlMChWJ2kxHGTaGrz
`protect END_PROTECTED
