`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VIbIemKohsV3G4o46wfkV221ewK9T1LXA9+mibbtexi+9d0g+GlVu9ZkYiNgviXW
6aoSDwE6tMh1KpdqzP1ov0Wjn5Q/fxJZVtdXw2kqwIgwAV9AA1ip33LOp2EVqRCi
ZhnBUN/6FF8/VkJHEDa1kE4ruTx7lauLCsZWY/JBkmeyUuOPNtMiS2JnZYLpBZLg
Knp+ysgZGpZyKAss0G2no9igv88W5j5DSRzH4ewR/VWPY81xI38nr+zC+RT/a36u
cI/mXtqjrExEJswhBZrpM2z8WJtBDor6c/0ydoDWNNqvXTCrYha3VaPWng7P+5Rm
4Fjceh5aAExbWg6GlHxkDIDRON6TpJrJXurEEc6yjJ25JvM7577EGXnuXTiBaZXE
oEOOClNa/SkYnJQjCWmieiwrZ3+QaJte/wBlQnNoxsh8e2P4f8CCJ+oh6s7u4gAF
a5UDPVhiIeRhzLbkfLnB6TbtwwiKPnbFJRka5KgrfHU6YYZkfWBQNJem/cnU8GWZ
wg5l4lHXTkNK/pOz2ITNsqcCFrdFRIQsiiWgpIdAc1ZxEYfyogXvqY144B2MCthw
GdYXTDOHHTBC3tfi0bZ1IpLUt9ef/iY8L0Zjs5HmMRbEKZimeVcP8mI8bM1drvxB
HHz77GyFEY72Im54YpoLlA==
`protect END_PROTECTED
