`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3FgitXnV8MnWF7uG1ZpBxP5XnZwlDG8BN5J333hI1rFdROq795+rvrEy3hiMD7N
9ZwVAtdhvpN6d3lsjptA/EA3jHXR0IOs19VEPEkybu2HkOVfVoiGpofO/08PC59w
UUlxHa8pMJkOWUEpyPZpXNFJK90W1PvlkDIP3bcdAOJJP/v8ZPwNeGaEXDt9XY2a
FjEqHmyB194Ba+7IDAHZZkgjRL3jFPl5/sMp+xHAuR5hDztJrJ7Iztctl5yMhcLl
YMaQH/g0f/e6z0jyGQRzCx5fY6PIxDcv2tGyrctSMmBDFoKhug8f0M2w6g8FiRsQ
Xfvy8HWaKuahOx2Sb1rmuVdiYO1yybnkHVG3PrAjOJKxvW6EGxiljYwrejcEvLZn
+ZjRkEoF/cDN5TmEXtzkxXmNHinCdt1Rt9EzQBaF33uq742W2D2AmJ+KXfqZ3niV
pQuzcLgxSkrzMNTkOLNtPjKQsy7CTGlRCggDsI3jTwFy3uLYvYt9wiK/HZETY02B
6gOX75834dg2sM9taadlNVAm6KwsVMm9yOceza8AQjYf1/pkT9OUAVt1ejCI9Vs+
49B3WP4WcrfPpLo548HTiA==
`protect END_PROTECTED
