`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2j5q6E5gpU07S5JsIhHBqTcGjjZjWr1Ac9SkBhuZnSQKPw9YeMdA57S05tXUYFIw
bpgE/6M4f09ujJW2q1kO8umseTfDHl5uUpF3+1xLW+3L4d/MuPZUZ4Ff83nY4tRB
+fW86CImwwYihmUDcy9u8VhtZH3dn9Q0fI3WWyNjwPJdfcz+UIZyjRRDzXZnIQS6
nGvlQ+ssmT44nfbZJqifxYnvS+k47cO/P5OmZK9inWIRmcxXCAClbX+oj/27bR/B
pwaDSSln44lZrpk8eUP6GIgV+zb9CWHGHpT9iMEaXR4dZ/VsreU5uJDbvrhiPaj+
MgvAKi6V4+NtFa8iZ1jLM+Y/L1whyh4S3xlqKWpwc0tXSM5hlfLN8c3ddtY+9o/c
KHQqilK2UdJQCcBDDTtFWVbqbX2QPEOqi8BaapjtMgP2KHlJtzQZ7vd6la5TConW
X1wHAKniNq/zE+oZolvtSfTiSNsytChR8QFdcG/FpCo+JJL1LiFJhxNpTCYy70XS
5cDy2BlZ2REKdxYpm/8bFdlJHqe4yyOpHMYcVqyh4Ax2vDJXefXM/oU36Cuq/8co
UzMPjSLg7+M/SpTj+bjA5iUOBCG73MOfczbcM/zYKznxlRRITUlFIe1SI9H6VDdq
v4Txewzj3mMtSAkv6QTGSPWZg/W+9QsZyNLFoXjwwaJVRpyItomCkoHGKl5yH5T7
ZsYOHMfz++YqlOqbgNgRVyUGRwku9FLC9mYpHMz8igf1Dsd9gcGRXYqZYW29SwHw
bxDAjgh6V4++4SaTUfqpDHKmOc0u7SHeJmqoh7dRmkYbwBSR3VqBUOvLasVRnp42
SHUQ21L6zMeDxOe42xAozdz4y3lxW0fKFc0GXpEY8bbrR/O1LUYxHceHiWM0pQO2
`protect END_PROTECTED
