`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wiVcpy/rjufc7zVCRi2xUg0ZImXAc5Twc4rAtJytlCano16dvyq2T0iKMc2b9hNG
lEEUtW6FweTeYjZ3wslY3pWhtxFF1B/XXRLvWZmHoHkMf828/tin8QkRrzjSC4QO
8L/vECUUdYP4vhS7ZTWHPuOKQ5sU6BqMpzbDVcLWxxnkcPvwMREZCoCuu5KtElAw
YcvFnPmLyXKcYhx77dTUFwN9MyhQht2UVWa2sFSDktpQDvbv652NB0aIuJhWeSP0
pIclBs0KFueuDTfAbRi8qnHHyUKURi9WJBmX6N+7WRWgAuS0s0lgwb7uGLoiCH62
H3pssY98Pq8iGDAj2k+BekWZcgQwYw9YYqgXfMbLTpm17GQ2v8s3QwyWaj3BslKc
KvXfa7gzxThWEjJTzn4ZA9xH2vIicSn+kkRPW2GH+xk=
`protect END_PROTECTED
