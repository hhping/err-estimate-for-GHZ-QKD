`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sN20unffx81Bf5qIDin6gxXklx5BlG1ryYqfloOs8noN7BaWBno3ND0777u8sRrG
HXrpnwuc818r3jP1BhIHtkW/WkbZynwPqRw8NHcjmDNtrRYNdzyw6KdXj6fonTiJ
opJNSHo8LrI4T7durPhWe333jvnAlqgUtM5r6w4+sVoGKpnO6hzfSAyA3//G7lC4
bwIQdTogu7X9/zr7VulJmmw6hMcSL3du1vB55vuLpNMTC4DEigz7hSYwWY6cZrJf
VawdRWzhZZopalyNwO87juKr3mgKKysKcH3HLpCOYGmay1STnQKJfEFTkTMh4D7N
EurJS/qaMq2zs4fLOTdQlunSc9AcQ8L6PcN77ABdISIg7le2adb0wLevIEszvLr7
buHtIsX0wsy7uzfXWpkfJXsPrBpR8ag42i635csz/xOegxpqMjpdKVYjYwjdQSc6
TOCzFW7FNU8xs61FWCUmfgRyptZSROkAhR9b5LAEyFZYgzf8rJih/W6+KbzzgwFY
fcUsfa1jpR+C6wc6LUkASffKxCYiHkZ6t1vHVWlnVKr2VCyLX2zBiW1JZLaEsUM9
HgX3p0Cdo2NjNdSrX0dwGz5Nz/kqvMappb/mc+7Y1S+4kZHNPK5asi0r+pYuDYjq
`protect END_PROTECTED
