`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1vbPJt+4mEf87EksqOOQkoqliDXKG2t1VU4rRbArLQrXn2nFDTyMBn4lNTfIo4+
5aaRXyfJ3lWicoxhdUGwVe3Jpz/78SgVS3IJjNFvQSWge2K2KypLqL/3UUqU5iuX
aGFe8MyywdyV5j10y5HXRbOAbU0x8p/nd+oaiRrlkgmT+Bii/afnhcMVPe3Wrxka
Ll8CSYgQdXdtffmsMbx0sKw8/0PtVQRyEfWb2rDWKREDNOgjg2NE5Hi56vUvkC0E
QNiYlBplev4i7RbrOeDIcsmJGm/0rbyITEViKt7h3Iw4y1QSC7YjF1dOcUsYJ4Vg
ouaI+t+CP/3i+YsCq59PJ5fx1doJhwMmwlm0nLTmiZO0P/LCX8rtaeczj71SlpWy
xGAn5vEaL0IraS3pcK1Lm0iw61HxKsp94ftqaMc2q3Au5OkrtAHbAGUMRJaoQs0C
immOvZ0h+xlUF5wWRFYdWJqD57S1AxctlCkV3c9TDd3eOSkW5D/RAlSp+HtwgpU8
6ujS99VkLzB9/vUWvkJWH7unHpxP60eUMwP9OzGkHWmklODD3OWRYd4hphqeMvlM
vytVO3qeBmV/EAWJv4ZXOSObs5F1dArZ6lpe4UBLTOeLjRmAzGwABKngeef2UL5M
Sh7BGXrFVevPaPOtWprCJ9RhYMuDRB9tcM6l2wiCwpT2okgLwbC0dVF4vMIrrPpV
klkKFrE3MHZByfca1es8H9MbbFGIbYd60DbXgzCpks0WgvNWRSxBSaDx6OIpxumu
ejS+7FtAP0/FC8upYxCgoi5Kl3xpkX2vlcSvbtyjG0+F5luZtXYORv/ZfjltIyEO
2HfRFKJzDA38P2NIYlBvaFfgLV1bhxDuGJHNlhihtVq9NLE+oHW06b2PHqD/9JVY
IIjLvrIBSqHiYyz/OZnPkIvZvXs2r2HpRa1w9cWJNBzTH99VylZmYgnZPI54kjzx
mgNtDY9GjMPIKo21Xm/1leDjM5AgVBSX+sFIbv2XFVut2cFjXauhKjJF1B/tVuYu
vyoPWg9KJG49CWmam5u5FVr37AIUaPr6MPNW95MW10dzYURiZTROkhRaEqByJ2C7
zR1jNl8wP5l4mPJiG+fMSCgb2lx72QVsB4XVZ+Is4a2bti4OQZMl6mGXlHNdxzr4
mkiC5XhB61h2Yty6YDDwCWRIxi2aE6y1sbWAjLlmSZdWS5B+qUerYm43OtSwQoYU
Q3BhYYasYtKgagvA3peI388j5f9ouHA3oz3R01bxEv0z5KJthhxaDVrHBMIwRhz3
qdC7O7OaC0nNgtWf/18y9D7FYBKCPv7z7FPwEYJ/wO+9U7q3kaXHvjFoKxQ2E+LE
ShsZ+p8mKXSra5d2PhV+/gghcz5eQx2HfrsCqrb4VBo1ZXBeQdIRXLMB/j3a51fq
KjT7puyiPJCiK2wB+8tqGXQ9Q89KI6LRiiIPg6DUR9uNhCfQaIUaRBQkxoCH9iKB
R7X7DZXQzeHeu0oIf9wcWg==
`protect END_PROTECTED
