`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCwETR/ZDYfdyYfpQuVVTeWjWZ31h8tjh+p7BsPZEh5bVhd4OylL0Jy/z8iXtqEt
4onPVRmysDs12Gfmwb1pa+Q1RLeuiTmIbMVGlpdNgSVVEvKlJ2FvQI2IfqjQoEAY
tRpnbTtbWhp4q0qlDqtvc9yDdyd7hXuDsNQYylGmn7aDz1LAOnj3sh6lksSaQd4L
n8wHXc/Q8kYxLdQvuvtXppS8jWyV4ntQlM1MxpEWID8FkaUSFeMkDyKpPdV7UqvJ
BZh/AwD4cOZHbSYI4/e5hIMOrbNhrbiHOkiLbFEXMMWNTbexg63XSAaA6g+nUXcg
vPKIAtAJZVUWJHbQec3p9Fg27mn/UjJCfwLO/c7rXxefbCkVTuEhHAiHAotQ5lJz
JWTEUJQUGY/uzmAHx58fIIIXWGJOx+5c576s4q2x5piSU5ApLaPsrS9TJQ1LK5G8
bLuVnYBqRAh2ZsYK+2Z331br+wzp0LsI/bpGC++QaVcXKHY+fxIL0nwquR9v31UQ
MHrdHERPwl1R6/RvpuPtXzprOkoIhzE+0A4Mrnm5NiHHLb/2pjAqolkYJA5zWSPp
gXU4SZvO35zrfJCXMdTqGbCgKeSb+HvMCGYKm12yNLr1AOlML4uPYJbVpKiIIBHJ
dOiCwtH2RBIVuzWHd5ClVN1Auv6iPUc597pBzQ9p/nqbGq1pK7z7EU5twjOc3X+x
rsTE/0PEtUp5sE+efsXjmx/PKu2EGtMzUR361u3dxO0DDslWHkng5hUeUyADJ/KR
d54Vey0bJmExMX/vDv8cp+Dg/8gcbH7wXFyOgUx7l9G4WKxdPPVUn9W9heyIv7Jj
PyhHqZD7mvzZSiPhN0hINZLwp6OJxGNa9p8jLnPs99uipg6HtEZnqecVNwODjiEr
3wB26MXET2d2Dpgc2BM9kHdfVVuS6GBEYqITrUBjx+/4dvhmpj3Vd8Aiz1RpXlR/
ZbilruJrgm7cFdXPm8rwIrDRPyrybENA7CHJvEpgjY6HNQQPaRiLrT1ycSvDFPeY
QFHqA91/PUB1fefgvhaaC0ULJ8Adj3tHSxHjyXO14aJl8RxNlqCyFAb4t1LA+kOU
lGRO8gGAiU6PR0M++vq96P7OKwYRH13eHnDOP9Pcu0FZ7ngmV3NwOBOxr0jLl3nO
bKApFGNpQ6G7/oia9gZ/xeV8mTwITH5EC2RjvSnUPYiWVsdQ94PvelzCdCttyDJ+
+poBHYFdEDCifpRw3uBixYKri//fA6uTTAnlHBeKNzuDibxypLJtjnM6QfW6UtR6
SV5VM10rnG/CJzuq9ugzYjWre0NfHm/9oaQX15kkFBNC9wBmg719oj220ZF+AGwb
rLN4Cqd30EfoBt8w3Sc6SLgUu8BvZQzj4bFjwtM8H0MR0s3ZovWPzifo1+AcYf7y
7UwOJ0Os6Zf3cwOFFx09+W4XN22A9KLoBfc6Xi3B0qJ6LqzhjhWMOMOj2t+T88on
CvZlH8Fm/HhH477ERiUEgbIfd8ygXNOAl3bffVon6KBrSADPNH0sZXU37sGqIZOe
eumM2Jl4phigZSVr6eSHn2kpGC0T+023serGMW5jz1JFhPlIjMwvx5wW4sOOXXSl
XVw00Uu+5Flh3xrVMWbc+tTZpXhBS9q9JjKdJAkk13O1Asxr2kQSbQ2C0Dl8v4b2
dpveSvTdzVaPRc5eX1qbihxx8o0++/b/cSYCdyUxE3O8DF7EGgF1To9pU4Yq1two
f2cMncFfqCPP2P4d4HJeF268XEKXLWz4//TLlgy+dQ9Bo/TGQ6CK0A6opTuIidUP
a4M62NZqMyhzv1dZBzL3Dt8S8ExBApb/QFWrxV322SSBAldOqplUu9EkqmL7BgaP
rloDLX9yq8pKZfCkjmLFfBMuP0zVBZxBAIldtLyPSsme0x3V9psdD4DVyL+7ly/C
OwJsFG3+bpXBr698CmdP27fACLYkZXZnmTRwFH6AckTdSUPugnijMxC0ujo9kBk5
hMbVjgqkXHpPZKd6keD+hDV9b1TO7AcfdbaF9VwzRyYQsTLNxkmkO+cy0NHwHqIv
tdiavcmB1oqHt/f0rSnm9hgY/kHMP3N1bnYzhfNyrIP1oJd+L+AU1Ixe0nUkXWYq
XyvjgLBTC3x6amwwW36X5Utj4oYylf2WEe6ygW//NP283pa5neDghJ9qPFrEVpQ2
lNbaR5fl7ZDactshLadtGPw43x6DMao2k/9UUK9ha6ddiB6edJSJvHNdgjYSPimL
qaP+PbNe5y4ixmVd7yoXbntS/fXXE/b8P+qAVWy0q/Cb/Cn/4BwY2JGQyfjG61XY
9GUvcgMj2HbzcYtG0dL0iU3Y6NdhFmyXiN/VoYZ6S94z+dF0TutQvVHeuZsyJia0
IMzdQG9eJj0TnZhSjfQt7xvwKNlTwwgyxysgJhYlPAj0dX8ZfWgm4G+kOhF+rBQ3
Vykyu4/mQE3uaCPgwWl2PoXvQv5Z8XCq0BDeHGqz+Xt5may5FPHYNf073mFqVXrU
cAx0MNYeg/dUI9KNp6ltJKG6IPouGMLLZdfYn8LPz6+SRGC0Yg6PaQQrIF5NJGx9
zT9xTOq3+yTsQhoOJBLQ2VGZmT3icyKo9Yu9UWOMZj1wqbZkPa8V7hFuA5MiPq2I
yMt46zMgAg5DM2ECXoLH1eY1PjCqcGaRLW5CVkR4HGlmvLmt8JyGkDPOfgK3+FIk
+Ni3oN6jkEH/7qb2yQdRA8PpDunhffkI1glz6iK7xhXFqZhY6WXUyKKpLGUf2ypJ
GDb/Jjqnw56V7Qkwg1oHDir3jVXZKSkDgF+Y5EXHW9l3CmlYr7NzXBObcpQzheCa
2sdXFJXuaVWQzSD9N5YHrnplCpGtW2NJKfjJMeNyl1a4muIZAfACqr84wxkiL2aX
HZzAySvJT4+x+X3UZPUjIZfI3YWZ9nSMFtL0yw6NybuF5jugs9GXAuqY2CCkkZ0O
YpZYr8lrBo/kGQtRsqibnD1WvuEoAOU1cxQtQ8aDNjd+OrJPqNWjM5PpPkrO8p09
Ix3e0y3TgicJaDNgoLKZ/gAzvcgwurFJoXTHaGzgqXKeGytLiL9FHL4IolkD+0sj
IYSV+tgq3QlvoDEKCQ4gtlXVHkVqnQbBVQL3lk1Y5SRGFZYhxZZdDyXLKi4kRPjB
VhmdUErLyu+rS5PhS2eInwPLHCDQHDHBQCTyW18WdXEs1lor7AbFNocSRJ0WPwa/
tX9hLLeDaw20s1oQOefx5ihTOc8sb2bDWUAzs9VvC+Qbo6JczW7k86Qmai8hqKm1
BBfnp5Z5QHI8qgSe3XZIiqUPCPacLOfza0Ao46rbO4Xq7lPg5J3BY9PWxukQuhQt
PByIpOvQq5zfpoqeuuSP27n9M31AHQTxJ36DvHKKTAyw7RICU7W/9LwHlFj5GqhF
8b3NEBQXrncWTQZGBn/o56KMXN7U4RmUgt4AOy+xAHH0QRCYVFUrJc24/0zJCOUW
P674pAkRBE4XqHBTcMedoNa+fNwZQQ55oqldM0BX7gjIl6YiEiw2EDLO54KBl9EV
BJjAqtfXvSmOvs5cQLYoF7wLg3JsMS84Wpnvwrux7BB905xSj7xNMeDJ/NmFJOMk
AGz8fSe+AlYkUc1RoPyzVsMsrHsDTc43EcXuIMLEitr5V5UV5ouaCKMztB6PZ5Z1
lFREo3iO3h1HlPjyz3FtIRWupgKuah6+is89U7fmA1unNEeeN8glnKqWIp5nhUUt
Jl5WbQ6UviOeP7GlVycbTTIbQDGxUByfI+1cCwP8m3OumWLaHBbyQhJXw8IxQPWu
/TfXQCsXch+HDQNFiq11EubGCRZtl7FbMTm2UeCd6lYh5WZaxqmMwhxylPKAFKrP
AZquI9ofwhoPytGaqUfdTXUnGXObnrhjIFHEWoK8qHlD8qrCN08kauHPRhux0VZH
zI/DEm8z75DGRr/qQFRuztrXf3D74HDpg6s7vS5v9FGrLzwPzGqfPWQN9BpNQL1C
VH3ohrgzFw3uL1gTWcBIkEHTT63NH+lre3KpKyp5dCWwSJ37yJV7oRqgiA6Dr9yn
FUq+of1K8ElYp/XEFfVCNBBiie0U+F3TJRQ5K5SKeoA/YdQZxFX7J6BXASMYnHWY
V/05sWQhvaWRpsurv/kJg4GWttmU+8JmKtYvZytmDNrhyv8yYDYR08GcVm0Yrxkz
dgYJ/AHf60uN0TSG9yOtJY3BBiZEOMX7OG0vnQ+5FEk5vPWRinwHdvPUvC+Q4HxE
wr6nolkPjqjk6NArG+Oa4RdKWEN1KTEPrY0P03ysNCTmOpLlHsZqdG/AyAcK8zTy
AQ0ZlHzZxGB8tJX1SCc0aNyeFRbQubXzRzejoMLDkDolZtt/04FSgJR9bj5oif9a
ZbwYwjix6+WfY2KQ9EeNRV81XHN7nD3G0SJ3GNnoEVkvzmcYEYjzM12VD8/mZUsa
fDdQa7sRDBacpVYUAHtVLgjGmrhUAunGbMCctcOLCQhjnqbOrk+fEARnHBdMRV3f
yeQ2abQnuQzJAuQQCC83QnOuOCLmHBk3aqe4b1AZdQxu2LIjAmiXMttW6+IJPfMh
LPpWWnyfefnvKOD9DHmb33T661ob7Vn7Vf99nu38iq+32kW37oNY9jSSZ8p0zLuj
EGH6Ft7kDP5bHfYLVYMKuHWwm/ON3I+wO5pCHzSSrkN0ZQCf2rGDIeqVDWtrg9rh
M2J8aYkMkSdSWvtojjEui7VlQiRS3hWzXSkbWNNLRSevXGUy7qMECIedoZMOBWCj
NVOfQlKVLJPcbs7rbuLrSxfimtxBsO5Xx4kGVWdjSKWDBisK4eGPtyJD8bkNkFvB
Yl8ZA6G9fyFRsEhkJjTit7vaUZ+oTaHrUN2IM4V12yGy/Vjgu/8siHyufeUzCNuQ
f4Wn1ItxVZ9EKvAsc5ZW1Hc1ZB0wUx6PPM7PrN11q6RZzVMLjDjyg6FHu/6SlJx0
JsaZU3AuHE+kteq4n4QWwcL7fsCo7ydcG8al1/0rhVLBhppgGj/+ek4E6AebHnzb
4WfK0vJNICjZX4izZfki7L5LVgxdj4BY03sijdj0MzBO32Fd0FYANFHo4C0QCfMr
gYvzFZ5WA1fZbjtbNshxiHwVKDrPLJPWkVQ/3eas/GbU5jPP06t6Vso7RcxaIahb
CNKpBjzM+NuOaCzP2YJ6jkze8bIiSjahpj1bezqOetHiQj1ocojGOdg0l5BQrn9k
cwjyWQHW5GFhjfCwfKHwj1FZUdKYFPr4igjpbEBOnlbzMYJ4h1jo6lLND2sQcuiC
KhdXX4RmOUwIK4fs6MiWWO3aVBRrdvjjCtFtpVOL0s2cXt0v8ExXQ7u0RW+H58m/
2AibP8+3mHXbXS+o2yCSQNYWarYJAdAjf8hNNDa8gSBYuA7YQAfMGQnqDoZVkEck
qNR1sbN9A+aYe87bHqJW3wZ3sDN1cAwHp6Kbct2uUQ89o5wtl9L8j7ycYWjAKDZd
9XHDtaVBZ+w4yYPCScUt/9JJtXjeLGNcPTKZ641aWa1wqJyKaJbSkuqXssMPi7Jf
bG4yl7us2F2k39kTnShND/X3RzteVgYCKH7vN8uo8bDsNfWKZRkvAvm3pq2I6Dov
4Uhollb20xlClg5K2Blx11GhQxxja3xrpEAUTwWLinzAqn1otcIHv7wvd8DQlcpW
xscgWKXQDnu9zkfbUc6w9hGE22RkIolIPsjLIZiC1rhxxNo06jxEpVKiolFRzf6R
pzWJ0GbdgIm+Mwy8cWfCcD29aVqHiNolpv0iOwLC4SH5leV6IPsKziXuCkAhJ+C+
OB41UxMCuqgU8xBhZF7oAnX97w5Sgau8T8KegVCqq5Wrz5m5T7aYC+NqR530Fzsc
DaCccd3OqInaxRti9ZG6BtyWMJUBf1oPOUS8GbUSXsGRNfUI5h0Gm7V3hd8vaVy5
iemqE8dGCXgFkbts38DrQM+hsz5l93Ef5YhBE+UFM1qP7GCivY5Rs6tZ1qjl8C/O
xcGTx67+o6SIlu0PZaGsNvxGFK+ujtxcoSdNzX9kguaV6kudZT09bB3BqjB1oq/w
tYTK93vNJlMES1q++y34yH2+SIaTxhiUzHrel/1ylvYJVC7vvjM5PG1XyWHLouBd
c3r50BpMOxSv9vqd5fmPvRxK9j4FoF3rIpg7UkmSaicnRFJm7EiVuYz0Q2LmJ+Eb
vb9Q3zqHKKBv/txzSfT/xIqEsnS8hgWaK/kYdYq6FE0dFi6HmTtAaSB1Wa4LLk7b
3Avp+ei5Q1IkE9Hq/7FzVlwx6SmZs7q94Q5yb5fAP4OZG9ybQBNiUouzoHKlBcRv
Mrq4z30Tf2bIfTPJ4qEtU8uUSSRyC2PP4HU2IMvLaFw/iZoxMLLkWN+7pi3iDOU8
1FwVbQYE2LhyJ/ga3Ma1NgXq6taGIN1M2yqx3UTeH4DEAS0caUzK6dtPw0/GrEPO
4eVR/kKTWxG+OMdzXiuDq97DHbtVVYZAk0HddUeLEr2LnTVmOLGZsyi+ndzq5zt6
K2i/Fu5buSix1ccyQJgxOnqga6KjJDHuQY/A1UYHpyCTUN1mtDcRD9hbsXTNDh2d
kFctUFcAdCkHE1j3YqqMVNTrKmlhEAci9/xp9TsAejfIVSAETTc2UR7rHzxniMJU
kAOf14aK7B/jZT5K3UlVqTN3j4amp3tY+k0kxeCjb2fYr//xWP9N8Ffr/X47Z6L3
YDkOVoXd+Pc/o6IAZZsZU8lBomCUdWnfTTyP4MjmnYsRDxSD7uJ3VXEIefptbeAW
+hhy7TZXWwOggQD/OmG6T63L6iJ8Ng7bzg+eMV2ff9wC7HC7la3km3yjV8cfaNdN
ofQsxMW8ALhLaRAF0Her3+cAEFT0VOQ4bxpcPgrsl5msSjJOPbfwM2Mfi9waqllX
mqdOeK7lawEHnhOKRxXWljZposrQUOR1yxf7KdVf5AXDkFDRiniDeU00ok7SVBvH
piF12eLrSCpNYnor1RolZJFFrqZctPL2SjuWWP7h4x7YzrtlYRJU+Rnn9QzJqS9T
R+XCVuw7Ap/dV7niVzpEb/Gir6Yc/FU/6mhQVc+tMudNEH2pjrjUG6Px+49NIrjU
LtJ1YiuOuPxhlFBlv5uGxlcIrwzZtAdYfIRVwbRodwg9gZPGF8Hw4k5je0DdoMbg
ppL69b1Ixlg2CAoUp3LNsHo0uFxI+P+bnyHx6iFTmGKCCon1MR5oEuxaZIgOdaj3
/2+BCYMdKogLNf64bug/LBhnorPekukp3hEJvsEeguqL9l8mv9w9yyvekklYSlCS
TCrXXCd3QYjQj+py1fGtSsEUE2GBXSwHBYb0fnO+uxUaZF3CxSbYkcDnQWB4MfXe
5J6XwWitfcrJYTU11dudqLe/9E5hXc+uSgvEwWh9grQVCAy4qksXujbe9jvK36dY
lz7jQ48ELpc6ygkxHzj4/UkXPeFsEM1s9X9tA1qwnvu79+mAZFiygMLkDvyLSd4b
VZNiw0/pwz5zvRCEEvDyjOorDTKGhF+9+aksPDgo1NtJnjVv1w12A2B143PHDZim
7whrSbqj8JtmDL7tfhvbz+84j5flDAFSWcD0/t3zVN7whf2TI8QgQWtv1TGS+KMY
u/1+pzUwpNG54ViKvxRq0Uwfew0oleSSyAD8E/PCoMDyHQoGjVy8IfQ0iFJ+215B
QDB9oidad7RTGA/T4Gsy4qIHxFQjQ9azkkiGWEztgx7j60A0mNfXwPJfcxfn3wVq
a6fdiKmaO5eBuIq8ZIU+FsBuw5ufpWxGgKm2Qh1LZlFk/jX730hrtICecC6TX8Vx
K0qWLiBNWVakhzqwxOnjAouJbad83txQikhPlec2Y7UB4GWo3Pf9lKRBqgvzA+Nw
UtEz8WRIeto2sWP3s3ctM7nBnN7pvike3YtaHYGviMqXh4tzIg3TY1lWkeBCdw7h
NtJWkRVCbJTlS2DTi6dGoTmgVbO3k+UNOAIus3Kb99g1nrKyaiEHz44VCrfuxImo
8jcZzbe/NAJNXbltdQzqahN2RY8JjnH8w2PYbjkr2Q08rGGQQ4imtxmWhupc+oGH
nO00dGY6yzLbcPEYPDXTkAlXRQwwBHeOclBlReaAxiodPSOFjTBm1Ll4n0u06wkl
AyMkXbeIqtRYVXBU8PddHOSZYfRbW1OOXT1wwZQIqLAkBFaDT3hT+bpwFjDkAaQ6
OHCRX+VssN1sEbLNznKNYylsBY2brZUKpMDb/xBDstLODKb5QomSiyEEKjzDo8XY
ybG/JKMhQPJzJPbFWs7bdmECqEXJUy1EA3soWoveJGTXHrlfpea8SoKl9mmS2+Wr
RqtYTHG/9abk3wr0+7blwBK0Wxs6/HK99U+lb33yVroBoRd4hiWu9KdTmmFSomrL
4eJqcANQow8JMXtUIQ1bVkXwDPB2kICpQ7bPXlCi/B/LCGycWgxg7InV5tMplXpQ
ZRVPi0MAROV+Lx+6X1kEtHn0l+ugXqpwk2Hj4uRo97UICJbThiLrYCpE96Y9A9g7
BBvjZJBfHdsk15E0yIPXUTNqMlQ8ZMKOTClJaQ9kByxsaDjH5v/soo6V4a0l7239
pJeF5lHtlA2x97UdjLhRaQhBfPHR1ik8ODndkxZJERDPxdEhELPcx9LZPj2bXTmV
/Y/dGDqL3APyz3qey2zApK15OKkqRkOM2Pkb9M7Ke8QfrA5OFhJHfdGMHkf+dE8q
BQIZrX8E2V/ssD5quIVl1kKeopyiPYP5prA9PkphLiDRR4eKj4T2OIXkw3e6P/nx
D4h0F1jV7RkbUtYdQIO3ChnD1Sd0Buj+Z+/igy1z98pknLlwcwuX/0bCz5Hm2C+6
XCiirJPMYEBnIJgL8boeC/1oeU5rDkKit6to1c+53LrCT8maaKq7su8OMm9YiS8M
N0UX7HWYcvQ5k2cK0R3C2NX+Lr8Iy0HOR0tG0s5+RHSygn5adiw1Nyycw7oHgp07
zbZk99YcaRF3IMcJh76wDnn1XpwLVJO7iawb4gPJhDxN+2ecbdbFQR5mgVUTXi4J
MNEijSLXcGRjMR2kzbviWrrHwhPXOXFoIIRmUPBBFaVgpiJJyAm9aU0vL5UvLhgB
Yurcfn4rFRA8OrWPhcbbz4LQhwdw0vg7wagdIbWXgH0fZ0U4xaye0ofWU6rU2e8F
79/ukCif5i5oMO5oz/p8wrikzdRyyTpcEGTgYteLcxZFje+ZrL/CC55vGxgCRuEI
2Lo7JAGssHyKDz4Qak05UQ0tEq9a2Xel0G5nSgRfs7PkLbKXNxsYYuv/ym47A0A6
CWvBc7PvaQCjZqjn5/sVafMwmriGwyWlZLFD2YR5gKEeBfE4HiBBFJWn7awIAYy8
kuwiJ8pAy0XL1YvEeawFBqE8OBTBJGEJB9UsH0Mhh3TtQKIMZA4l3rUyUXN8J70O
b7/IsxJ1wyKzR7AsLPhClGIxvdqo7vw6sp02kZ+99uDPmQQCCVWdAKrtzpNUAses
2AVTDNE6r2bXt2XBPQPBFYuUbaHPBazfHgOPZPeukhsRfKhaNs+kUDxRQ590BgkU
JzRA7OzIFZodHUFWCEjNLMDRZ/nyjm6++hAvf9051IxsfbOn+seLICjfw7k1dtO2
2wEKUwDky7PoNWRzL3nMnhVTDLf/GYQDQ5LdL8/pF4QProQPZP5V4SDsSGd3KjN7
mFN+/VCIZJ2zHCKuJPxs8RWA2kntCylmgycTEwObQExcuQmAXlV6RH8Qymx+9Dfp
sBVJ3AjcJD9rru8If9NB0y6aWo44Fp54k0xQxtla2iIemFMn/t8whrDJ1mUh9mVe
ek0C+Xbuth/kW2TaUm/K6mkL161Y1vavXSkkKyLvD3j/c9HBDNhvuqRjMNjRExI5
xzhh8ZzuWzvCFFc3AXCI4vI86xmkcu/l2QILgPie35Hknm7bHfNNgLxTdrmYAlql
d01WSjT3NchPTehO4CpGS9rgyQ1cj/MhrXJDsX0e8icyyf75GIpU8+tJrXpnLMqA
FEaZtAEBbSD6MzdS6CuN7nm9OzSyT6KzkMf+ZFJ3FHb/8oaa2z41M1MG/dnIW0e0
su74x4ofTKqiRiHiDmh6jyL6jgFRdnGg3C16jshT//mm5fqgINoioPTTHan2ClWg
2kmNbk4FTGrcICpgFg9bJmKlT3/bACgMiaQPX5nr7cfFn621jJwErRTgkinOhrIi
vnT5C9WjNt1ph1I8LdqWCau0u/bDytL+CLBVWMG8lLSWISEGwk/4jgnY5oRgqn0d
qg5WZB2/cF8QktnZoMyRBcWnqiYqenuJ5oSIUMW0m0YbIE6fI9VYI7fi0VqkXo8D
oOw7YedQQyPVR1yD1syTencgw0jAGF7yt5za8vRMR5c664MZHWlPyKVmlvqQxXDF
h6HZWUtIAUOYjgWMr9wA9i07dG/KtvdjLHiMbubNIfEr80DWWtRvb4ARhjPztQhU
8rIiLNPL261prk7CbK1w08xDaMdQOQsuTPvKpUIwCkAIFeox/4uZxnrLUmK4h+UY
5aSwZsa1eJuXMhPiaJoZxHE4NfejySfh1Q75yInxt7CmNfr107Q8UFnyH1ZglOko
NTOvg0SCYa3GS+rCEXy5vbX5tqKSxfh5bv8XwPEdIgq9kKpGFNjWFbEbzStskF9f
7CZ3OpWlMTl2EEFUXk3RmDKd6O9fntttkr8YgP28yo+BnKQv5E0LAWHPhCVZif8R
wfyLWpiTvRQVVw9RJNZOkbebO3BfRQQPLDnl10eIIrEuZGx5Xy7uGY9a9OlcIWnt
Wj0hPgXOoV1BcosSFcsmzX+i0dKhyCYGfyERZrUwl0sa0wvSWGPaRM0qWGBIGbgj
022ATlNpMAKgxs/JSgyr8RY5x0ZxzEmo3W4jtfwiITs83I2z+PLqXtQXno1HFAXF
gvjffxhXKRz3FxINNZh5HJ87/X4+B0wy+L1RsfiFKJJmWlydc6NoTGLLv6B1GRj0
NPFLctnilYpfBOR2u+GOmJltuTjTEDvUpT2IEZtDOWwCitgKH4wa15Ede0BKXpX8
ECTOptSBxYpZ7T5veHZxIpBiI7i8F1km4kfJ3cgxwKjTPLbi+JpiJHeFE8p7u3ec
qf278n+C+NHhrJDdgqX5b7Ggvssj8CV9KdpoxBM/gkHJkJq14TxPvIn1I3c7jNj2
lOlYazFeUQ+D2midvUJvdkx9utNiLDRScDW8vyZE8KBFwxSofJwXSdTs8XYUz57L
j4NEb5FSEb+zzBcrvaCNFye9/mcqwmI+fDpIy7nzgXr56/AdBOVsK3MZasc1SGwl
rGi/cbjY356zpbg9aVxbSjLsiEZW1djBZJ3RV81HCTKS4Su4PORHVmzmuoFOVCnY
ZTKx4WNChJXODgDBvdZsTNjpvCxV1+wFQkFHKwwls/+r/zA2N1x4kBvIaUIkAgR0
EHPnYk5FCNx6iAh6KIYBZ5aQ7eJYrMXPZrCpuoogn2r6Lmw+X/5CquA5GvnDNoS8
aUc+KizJA0UL4+A+CBBG2pC6+PVUcu2e5IETYEJdv+yFEREAgUznKsCQrkFG7gw1
LwQ5Pp5cSyscX3yRyepqwa8Q91gTHzXYxH2jbBFolX6AefYKbgFjFdDikyRY92nL
IJH7xGgX3BnuMRffbpjxwIbNPyPXJLI96+jL/9qaSj/YQH5dXM9DnYfdKQ7eoSF2
TrLyBz7pdLESVDj3T1tlxdpONY342/UVX3BEH1AzUXrs+ojll0ESubdRO+igopbB
KD1K8lanEv38bHmMb5wR8kgG1NtpGNhuXDOipcI4Lm0rhmR2bASVMnstVHc4RBXi
LPPxAs0pIm1yoxLrYlkC8u2wEbEaTR8cvtdyCq3aQMawI3TGhlfXQ4KB5PNZ9Rm8
e6KP5Fcw3rRzn80jpyko3jHe1nswlTplDSC5Cru6phirJ9Sn+zYUksvrNmNqvP12
jt6HoayALk81IfJRS6YayHOovcQTBmqUtvqrO7Ip/vNFRQkhGfU4CXtzgYqC2NvE
kDmKWY4yzyV21SllpKtnklxQotorhOlZ5BspcZqvWbBzXUcCci1fVl41VnGL0bn+
VL9xP7a3wN376Bus6kWs6nm+NYftrVixpcbffESrOuUNZFATjh9ioJI/OT2bFXHb
RRCiMkGUYzQRIR46lJTkMd6BGYwSvQ61bfF+cPauT4fbdx78bqAiMgDSvbf4vX4w
UV/bCH26w3hf66fbH9iz0wAKsYJo4o17GOhlBbTuy7xfvfIBiOTLzdHqhl23Zefs
Vax0G0gEg/LBbRoINWovYN4qbW3fOwKGr33a3ig/nam/d8yZUNstw2LoF1G9rCvB
k+H0Hn59cgBVo6zFVTucBhFp+WAFLJRCpUMgwwFqco09WUuGJkFaIINGthvDTkO1
ZGi2is8GFSr6VYEhCzgRKtO1OlgiDOROltSp7yluiCMpS/rt3aEGpr2zdd4/d4Dz
PceCtne7u0tfSPLxcTvTNr1hWZUC4lOwYJAg5qmbYFN7+p0idpABu3YVS8v23fu/
/PKoOh5n8fUEbdCxEqApa85F9BGEf2nm8p5tY3C60IdD0j4pvEuAD7ZBnCebauiL
nEKbgKB1EqbFB35ypvF2EsNX8Pr8c+/TJvDiRwDRfWGfTwP8MXUBZiQkgTAI+HEf
JyrvgfhxZxM0wH/56FlnWnzZUiODDaarvnC0AZv02I4IXvNaWS2aX4+5o87WQrCK
jOMXr5mVrzxzf7SK+KlcXktKD9zAyPGjX+zUwT0gX0M9CuCkL4Zrn+96okOZ6EjV
fZZpwkRBfx8Eb3L/QEbgLTylbYMzZtc+hENzftCEzFW1JbgABIMma8CV69mCvUl/
ofYDvee1eXQIT0jB67+ZAaD/flwd8saaD4Ko/7JD4A6b4Y2zobCfnGzlEEd5Dw+f
XIAW03Pip53udeAw7I/86jJNw3Qhkb9efATSS95kZ/q22wMm9bT10MqCgLNzkgAk
QbXLIOkUkpO+cwE4rA6R2F63oMEcD1o4++nYbf0xNesNG48WNDb3Q4yy52gVJ85m
ODh6H3yzZdGYFrWOCQ2alXcov6FPaQGpWvCBoKHeSEeEmfccXhWq0L3mNP6NrZNS
o7rtZtCcQFawAlN/dUmPP8GWGBj8S3A2BqFRX3L9iXCSgT2qY0dilKQ8sL5lK1Mj
ewBA1Vb2tXkuC72xa7wLjc9r2QS9bKx5VSL7ByNbsEanfvRH+foaasP43QY5n5mU
wdwIuGnpsmrVkJT8bGl2wZf4i4Obde1RH+KF4frhEmFQ0num22fGYgu22kBBlwC/
bZNybuZ82AwJuGo0PiVCvUXuqrS80zN62rHzs9EM9j3lFdSUTUCb0VMpchZg2a7q
nSred5DPZadVuYsh1Ek0/RcpZSaZmucU0cYxDQctp0NLq9AUDtmxAWcMtMXiC/aB
8s8XkbIoVfMEv//TjKBoTSt3sZ2asOOHnNNBXgA/4vj3WFk591n5GJXb1Cetv0Zd
MQL0o3ACaP2eGNWl3+T7LRvJowpXTgTk5nmaJnqR/6MrPrQHeee2y2rtyJtJK9GZ
PiDy2U9VMwXpgCwz8JJgsijtyjrSIOEEZD6EW0Crvce/nuUEt3vFgaq/wV+65oz0
vsRCxj3xwcFrRtmsnRjE+T2HwemikubQZvKcSOa1LnGsAtdAh1JpR1C0QMTyt1He
ak1o8whZZ3afuHUyP5ZcWwYMds1v+pPsdM/0NjCVqqTmHp3BPfqbsDBRrRiniqUv
R9Mp7Fob8yuISK642wkp0AASrg9GmX+T54cascLqBvNGkWU7O13cbmAIgbYDTtC7
UA2+4k7+Gpg5aSFNjW7TFtSiC39AJ+VBn3yfMocYktQ+FcbizZhNxELi9ifmTToZ
M1GaJ5MM4RiNLMMyEvJUeyUZSUaxVenbb9Evd+TqohxTEVebJUaMxh7qR+J+PP0a
1PEb+P/UUkL4o2BVwZh2s1oVzq7vuZWql/o4+oM6R6xpnwq5NnPoAIqgE5ktM2D/
7btpejvd4tTO32BTRSAT3vQBT/ueBsU4jmQa8lh+Dmo6JD1YWC+2hb/9wwolrLlO
lzMyT+yi6A60N1JOIj+QLzSHscOPOOPKQ+NRmQq3zP1IM/3P/cqK6uiU55NGG2HZ
DRcbxJ2Fls3ttA/MiT3HtlDCRlQOM8XaTlI9V+4FXfonl0v7szhfWODSkPI2Lpy9
zbxsKFG/JSHnKFQWqFfo1ZhD3tTHv1V94p/QT5/+Gvh2TcZRhGk4Zb442NKs2Cmb
n0T+g1naICf4esR0SytRbO7fgV/DAuh/ZGZoUPRfTOOofenTIaJC2/AqpqCEH2k0
RP1IDa9/EL59c7GxPggkZWf5FkDUqoNLsdwpxw4Dh9iqDEnUBkJC2bNBLG+iRcCa
EY3bRFQ88+iOpRrto3XhqUHoPcWJWfYPby8r3ZK9o1EQmEAq68bhED61lR02tBcC
BmUDxiXdoIj7pvUh2YTBZbAVRC52FeJBhYd6XT3N8dKIxIYJhhaPQ7Df+MNgWQXs
OM3BC9njSgap9BFt/zV+CUVE25z+MFuUwEelcvSSOI68lfvt1RLUj/Fv1Zc6JILE
mxXuWNZtwTeZMbEldafbkbZU0e8tfhg1tSudkAgh1Nm1edqzzZqNLjEamlaDRDXg
xdSBZWRftZMzn6euR9gdSifwMgBdVpGLGvjeVBOr1BCIgkiDsJhMhxoQHsbho138
dUTzrY1e0wHXIHd9hNS3/R/NspGrj7gHZIXVFglElpLxvMqL0s0+QLJn4DRo2IDj
6asdzsHpnOME4K4iYGPJIayabXdrOT0HtICL3Xzc1q8=
`protect END_PROTECTED
