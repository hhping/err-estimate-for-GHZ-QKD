`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aC3K6d2TTHm/njytJdjSfvByGnI30ie+GB31Pg9ZtEL/2TbnrQLTdND8/8sfRlmj
SBP0HLO+SBweu0T0uAFLpz6rfWIrU7iJN28c1aGy9oTd506VA/mOHhl/2NjyznNN
9Vk8Kncmi/ixeCDC7g7P9cYw4Ttyx+kJwE/66g5W6Ci1BxyUZO3MtmhnkYvlvJoP
wiOsq6L+U37+0roGs37+JqkD9D5zDiPvNjYdhnLhXauBmZjah1K+a6JFab6NYVgL
kuRpFmafmCUFmYGNwvwxZuDjv6umyM1A6aV8PA/ig71mpCAIiTbNyKrjJDgye/mE
9xUNQN1N/CvktCvU22cno9w1uJLLsfqqmxIiKtNcPDf3lLj5u6ox6B01EA1kj1HA
EiSrpm31H+UNaOH+NjxZfiXmEJ3djBoxFQhzk8AskMcRQafr7mju3T/o673oZKhx
m5Fw1UVuH3rCaf3lZWMSnmNbjP1CxIV0/KCUfDMrmwAja4ZF+zfOWpaW3ieBmciP
dqMnRUms6H4Nkc8WrtCjQrAVvXCdMipVU7WME7D04SYyvhZ3gALMD+11PJRKgPhg
a2rphhARfxMkVAIhIIk3p7zFeyNZSJ8NcZiJaDXkLwgsfsfnqQZzg/THKy/Lidqq
u+YuEd0NKIg/zB2tfOuUPkgtimFll9IQcOqoSdp1PnXxwWCzjPpvnP4uKrqo1I1A
Za95+87l3WjYi1AEQuWMLrOSB2TGFmnhz79S2IGB3cnI31x5rElreLLYOLjVeDCU
CexY/9mESlT+JuyNsXJYxGCV1NSLBEzXujwx0VqIoaGMQdxEYMirGiZkYpet7F3r
Btsoy2CIZqEeg89cY50tHNLcEfIMoLZWeVOO3SKJH0kVXqr07ZcMRrF4Tc78ul0q
`protect END_PROTECTED
