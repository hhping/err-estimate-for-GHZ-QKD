`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqJBy1yKT+DpI9vF4e+BBI5M0rpYCJ8/qEtvuCoD0JhXOHce9jEg+XzRA//V1LLu
Qdan3KAZJWrKGFWLhihSqS79TZi+nY1j3iSZ6rwSbPnOHBQBWMKhj1BXaOggqMJ7
eF4aV9j2CCtM6mBUvHBuQ2w4nJfnAMPfRFgyeTnH7QPYugSuitjqZEu86Q25TpVl
KupCgywmCe4VTnjRLCAFpsWK8AoNpF81jZ4hwojHGAi5cM9rVb+So9sMtAJQGpB6
Ocs8I7GZ8dod13fo2NUmS6oyemODSXXgKiWTGA4XmuBj0t42Zey9+SVP3bigpoNv
l3c+jTTjzxHnEJ1XTKeZLZ4LxaPOOVQEEJX1eNRN8Bw5WVNUdow1cZ1S2fOCiJ8Y
cXpRaZOgKgKarSjdvzDAsqeskqatcHpyb438aNtbGV4GSgo6Sg8zh7wA/GH8lFYV
6gdKgTiAhP0jiFJ5KsD1aruNc25lpfzagjC7Jt4XbPunofMpgmeCneoAectQZrzt
mniylqBJewzrN0NAL5I8I2KRuPpYDIkjNa8i08vPIyxwhHkgJ/bMd5+RAnR4N/n9
SFdF1bgU5zZiIyn9ltWyx6RcKuYtn0TBnVXRfepbXK0MxAZhMNqRJWvTTdb5ZQ0y
vccrUVr1rPLDf+OUQF6bfVafTnhrgG7Od6Flcsbsc6TweFJfVzX2ovHyWn9rARf3
DstoH2ShyxvEnlJCdPazuwyjmegb130EzGKMwxEqC4v9bj1Qh8luLSqcDrffRb28
4FBV09SyX5JOix2jOcLksLVf7MqszWBOF/jqrgV+lQM=
`protect END_PROTECTED
