`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gK+wn3KTUwQI3Y2H6NjDQcDXfp/33eURO29rIXHw35r2hxd9NAfiLVWa42qeOayB
hBIGMNFdoazvTbwsOU1RjdCDQSCq1mx44QaHzhCjB5QRFnl1Czn4nL3pCunKTAdh
L8YgcHeD/wyC9fvtjXaFFDUEONR0pCCUnay2jMQQO772DM7rxzWBUOdiFbYgEg4U
mdH5diJPzWFRnnuSb561w94//vmg3WWrvnl9A7TXdgkxO1ZGNNEE8afZO+ZskYUG
yFE2CsKqxcw+gQ91N5HIFm7HChbiuB7q8LN1ue29PIvN+Vp7ApNW8eRjANNdmb15
mdv/E43cev7JkUKtxHWzt6ing9Sj6wk1tZ7+uNNyVvQlk1xXI4N0J5FaK19llxVF
sYFQVTnWJWbNYotyhp8hSpVFY927w8GJAJGvycf4qm3TXRJrkHLWigp3RCQeEsIw
viL27skKVsDCONpSpLvI2kHA4gH8m2zr3y8KT9j8WmukAUvrnHS2u0ZSVSKlmfzn
T61NY9omPtCel3jsny8UyY+Kc3oAtbGA1j+rms29XS3VcN5Pla2qY6qM/3pC2uxo
sHtg7ON7BixFFv4cZ901VxX/+2MpnswVYPx1022mdq8VdENQ7FZIrXF1RvUlOBBb
aEm6DfKvg/GjwVKaO/oFjzDZBZ+WAPAeFfjbPi7KXGI33gBkxPeYMQ9nTPIysze2
rJRRi3wrF1fE2Jbt2MbUQlRPy3pcNYYTx25MQ07CvnNibG8nuKh17Ro/bPS1eAJ/
nhjnGaJWOYEjMsP6fMRQSL0kuBeQknvgTqVXu8tYqmxGcCK0Gq01JBt+lUQRw14k
o/2yVhbx8gsFUyas/OXY19LkQ3Mjm7RS0TrsUKY+HobPSYnsEEGyw6IiUaVbBTMC
1R70qtfh2oDw+1xjCXuaR1rKvHTOock3XnFsIVzAE4g5jfhNY6Ai5/cLm37AGuNL
NSDsaTxh6vcocPfXYVUq3pah2da9fdqNmedPGz0VQb1u2f1rZSzJLb0UWGW4uOIy
keQdoQOLyMqzb8gyuAJDuzLXgZaynsP75oIUUSptXD3sLKjxj3RvQO686lNG66Jg
5f2Fp5GpI3znjPBZDs/t3PC+wnXfTkhTLW2Q6lflKfMbe4Je//hFHhLBymSZqIoW
BSTy2UmkyweJ1LqiDwfUYzbosfpJsOXuAIFooHQAR9omzxd6no4MRFjIJGAgAcQL
BBxzjORNBfBvXJZ+zDLtQ2qXlnOnqrVMvvkGiqKPERh+cuoqZ8dBsnZrNDNrLDDL
k1XoCdZeOqPeaCOcWU7/K8LKwqqS5bpLYoQ1xfSwlWn0E+fxHGgQR5ifq/DnDH36
ZOl92AgPt4eR1CwFthYuK7DjOLJi1Bz1kmMMAWuXkdwc/Nk5XDArd6ZSs5oweWgm
aYr0mHSC34eC2tjZ0fQJYBNNJ2Wel/OtXJNrFqdvaO2oSX293OUkof3b6o3sRp+K
V/pdHl0KotlnW3ck0zooLdUWoqhxbpXN866QiUpn1+H2+k9QKsicxXXAibad0MPF
j6FbaeJjy35psUj6YUrWXN2YoOJ2gQEA05iHVNSmA4h1rPK0s54p+kkk8a/Mmd6w
rmymiysJGB+VJiix5qDO+OpxhTX+CEAMkpyNfyX1jiAxl6FQpustQ24DnnOO/+1d
iMwHTOdrMIYbL7g14sUflyFpa7h7qdZdIjt5stnBpq3vNfAn1YXfPjOgLHJvoesk
TjhAYggz+pP2AQWmL9hM61Ig37a9wDERO0XQ7XWJbiKom6awWqIOTYkIk0gjgyWb
X6Rh/5xXmjGd6Hs0uccb4azu0x1vxPXljA6fL0tdKqJjJ0eYrFQAEUChX38NLvPx
iJ8UCMLFHFphk3Nh2yDFme24L71dHJL6Nt5qvkWgzWgJqFpwb/RHYZWId94gzbGK
n6taOhDzQUKeYJDaTy0JX0IQ89qsF0YqrDx3TiNbWqehCUUU7Vw8FFgqpnbG08cN
UFpcc722uEuWHrkZVzH4iippLC7JTH9KBOuZ8/0SxxcXkw/SbP0oHkZ8cpGoO8bi
7I4CZIE+mkdyRXbKkyxuUBX54Nz/5AnbQvc4WlgrLGSI6uFKL6w3KP9Aro4byVLN
oiCt6r3G75DZNl/50kY2lsGnHpQMzmsNu99CY4AYofQtCiKK6tXd/Ufp/BJKPt6S
axKgrvKvy4u18g6ypUZLSp+xsHCgsnXYwqPgGhd9Xu2yh7oExk2UkJEvtWO806Wu
YJasE7p5sMRrk4xwzO1gRfX7eHbDl1Qf2AOG8HgtlaHliXyA8dSCCrcS1A8qSBwt
82XhRXvTibhLC/yQWLdXpMgOt4YI5Lv4iZXalAt7k9mVvmKXZcISDSzcpcy6hNy+
OgyGkQ1t8VedBXNIzuAdZ55LZy9KNoKw9lr14ZaO1OElLA7rNL7Ck5IhrC/fnzy/
sNSggWIRvI7HX9PLvIRx6gWwFiUB3bf0u/rCGR2myVg7cosR8PwwMQvEw2JzE2fE
zWDaSSKJE2+afCvhnfaRF1kmdcvIv4E1AjfaAATym6e64lef+kiUwlpGnQ55+b77
ufkvxfwfqNbhDsHkloeOahDEygxWfSUViBs8TJ1H0MBT1UTvhRoHzakbTA5kg83N
1Mt+r0VM9R2o8X9e+jfzyB/08krSwlOaGeVZqwtLC1AXpLGWVEcMMXO9ac1fAWf3
iN31EihazkVe/EIRxTFugLPL2rZbDA+MYkwjJZYZzM1NMFo7YxP4pBglVJ86N0HT
oCwn0+/ys2x0iszN/LaAQIu5IrtqloJh6gDU39xRpvmMSA9UM0g/0hroLYfGiLYA
3KhMZ/pHkmUArt7lHVlkfJ62mKSllpapF8T6CNzpW3qKPOfkRcb3+wT6XV4wyegV
rmkHuTR27yQnbpPjsijk33WRScoWdGWKtm8KCzeODwm4/1kAH/5uPLgMB5rDEbqu
WtttBFF4ekF8kpsARCQyCflDl/eExzX6R4pni9P/dYzcR2jAIYMPVvioo+xun/9w
elEyFNys0WIsjw7BY5AkL/ImXR71TZTyPZn9l+r/RJTbZ2ZF/XJg31F+geUhY06j
yBtaqq1pRv0S9pgKnXjo82Rd7ohtBgrkeh50HurBfgg+5NnjsL5/K3TteOjAc91p
INKbnvFtCGIJ4lat6mt+jtDlIk9r0FmmrLdnKS1382SUGQtN4iv4wXv3lGzG0GwZ
rMrLrj6R0Jyck2+hdtmjuN9KeILTTYLLPrPPuT85esuP8p1JE+3GUhvdpf0FEEt+
esfLa1p9g1MOYhRT3SXq2g5vzJnT2roDnNYFLpB6Fm4bhpUcGRLhN15uSuu7h8IR
a3Qlfie6byQg6+pc90cxpMw8kXiD6sMJdnbu7utUGYp4U6VKrh2dBj5eF8dDIYhM
hvKwZsjepWtq8o7/MCo7BcBa+Ww7sv1BTH+h+K7iGQ3g1T6G9SXMtEOS6DYh70eR
7FaFfTCoRIsmxII07j6UAZeohl5jlMiWPPig0HFwSuQRAb+JXJeXW2IofAtXvfl6
nd2qpftvxg9OzgplfHGJ4bsh01cOL+H7lg10FP+FCUdx3+YMJQbd2FZQKzukBz5c
U0AhgtDDp0eLxC1JerfUSW6wtuq7f7YaKeqRwoy5kTMZTcnvvwTKarCvcNz2+FVc
Pqx/fTSCxwtKx55gzvUHncluT1V8JNpwd2eOArakHB3l1kQoSWdENzaagG4niKUG
0sFsCoOoaMEdTAl18Cbccd0E4KxoHRFtn8ykFpHkfLYUOSEwIxS11FSvUQCtSba4
AwM9PXKDWCEf+otbQen6qDxnP0SjHVMZv6XqRupmKRktm9oQdeQCsdyuaSL3TC3G
CkXG5J17yFvMXvT0I03ySigZ4gjbHxWgIYlpyGkzM8oXjBuRZMYIW1dmhuDW0Gaf
axn6a3ELn+yDZ/kc602RaA8LPFwfkmJ1nI8DCPYMDIyXZ0909v83F5K8msY4i51U
t1rAKBXstjisyWyvBChzvNkJiv1GKJZAuIECkBVCtPbt9pGhqaiJ1gMQ/Ezpo83d
erootz7KpMT4GXOSBWhxqR3O5WA8JOQ4JfQFJ1Z1YApmPJ2zSg6il/RWxaoQHU1/
XlrtjuH9AkxDAnfLTIZryMrBsKyxoDLtNr+iatGsVTv72NIL0QtqxwzVSKCQK9z0
IYBrwSEyFeIqu0lUiWX2l/+baEF/3dkFdubC4vtzemXOyxS74k0sLKdw0f3FKEBL
/cejDWPnfz28GUV4xrdnz0vM+yqnygFK6OcKjNEIDs/K6rfaFuESY3CzoggGezF2
8DrLF+b6Eu55hhq4RaDie/oStdY93bEMM4NfUF509nZ3sLTMHOmVU9x6Tv+AWz/2
Bmyu8lPY6CTBsN3k41bdxs7v+5BRyaflF19aojwZzfHmoRx0KVNYlyo30tJv//sK
5B1FQIHTgkC0AOq7A/60iU6wtEzHc2UNDk1EQbf7Hc4oBaqpu6X7jjEISCDJbkT1
0/GiSygELSoAb/Q3QZoKD5kGKpnoamJGrFYqQQ13+o97nWz2bRD0kgHdkF3DTmz1
gX4zL+WYwzOEV65A0ZYqI8y54nZhRLuUyBGMoS9Fqc7R6LPHVktmIuI+DziPGU5x
IMm3DQYTopp/RLTV/NOET9xHGrR+U0iQzuK2/x+js3QZ+3bM9TAXtEgAB3Q7D885
lD7Fbqy+pGnnzGtC+ajjRW1RcIid2JWr1+uqpMz2momkpgS26iQNujyzx+Ci60g9
1PcKBVd6flhatfxeTT6weojlwqCIjyBYyJrvPlrg+tlB9c4H8Jd8cd+PlHzDfaCX
RbjvHfcZrFWzNogQG21R0wdGMess86MglvSjBs0mDJ7ewtVLo5w5iSXEpHfNNQKN
rxNO64YsfoQTTAVodh3E9dwTCNJQDINCE//jeJwtW9XV9imPyX4CJGaNHTwwT2ko
yLsI0Z+ajMFMrjSmEZiQPr1jWjiMJt8ku9xZh14tRRtHtzEcfodEcASAvKFKyS2Q
K5Xk7zYxmifPcwtSD/RXZ4HYX6dniOw7sDTZjtj/BZorMQ+LGwIBLF7p/fF++NOz
cCz/lPTWMnbUSHt1ThoWVeZ9L5s+k9HTt6Q5MB25rgpMxdvxKqFO0ulFxfFswijc
7XmUiURxLGom2d4An9s87zNYBq3uJSVOMIaAPOvjpRmDQQ61nzFAo6oIYbZ2ytvD
afdMshQ4fsa0lLb/OidozZFZ8QS6QYMPF/WmLRlxnSrGVkznKBM55F/bGfR1stTm
OFCAYqhLbs3omOA4ETOGn5ZHguSRZQntB9jF8Ps3Z9Q=
`protect END_PROTECTED
