`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCToBzUwl1VyOQhDNfbK4CUm8iX2XKLTnz9xGhm3OaMIutn+a4mS+uQ96EfXWjf4
sD0uZaxtWtPgh4TUM1hH+o8AhXbudfMqWLU6H8TvxQaPba8P+9O5dutW0GuIDZ2B
HZe0Qs43M3heJ5ts020Pv7V0846yBts5qDRcsqu/3vmdK3Up4j7J/dhNpGrX6yOx
2TKHTnpJ56G4dgnTPiIuQMmFLUGGTpRxpiUcyNVhCDWfITh6M3zg5cDvWuaabGdB
Wv8FVcRirO1D2gCLvHNtEURX6ly9/XQvJHAV9p1Ab+ZlccTz0QHF5Q9pu4QHxtZ4
7WtdOp48b/ZvHWdSiLbkfnS+tZ/ntVfrV4A3aYm4y/dG1o67f4W0PG1Qt+1KZRPL
ZuwU8fagLAZGbt/04J9JpHJkVqBFwYbsFIeEs2jSmdYniJHSkj9iiKFqd4A+MY9k
lnkWQ+98wq/xMRL4wnlpCTpy0ve18rPPS1iISYJjsw+Pr+s/C91NkXcGWjNgRB6M
g0VAjdFLSnyuwIutpHmQiLjeEtAcKRNVx9JndPqoD/hgXPf0jGXTeSA5J0io6vj6
I76xiHbR1cR/yd/XRD5nvMp9k2MYfPMhLRaLKwr7I7zOFfAgb+IPv0nX2zP2Za6/
OwGJUDEjQ4/rUGgx+OdEKSJHm9Mw0ORgkJgIdSSJ3LwDn28mjejFHXTSq2ddE525
PRdwnJNkKf5pjjepLFIRYqvg6+hRa2guZClSZ3tLM7O05jAjOqZkutfTVwWQHM1U
GnMt1D/EgMfMcjzbd1BJBI6Rp54uqz7dAkfSL48tdD3cxdhOiLbK1iiygcqW+3Fi
IOo374TZX4YT4K2eBEReETCspBthyabaPRS6eUPNpZqJpDGxNB7eqUAFRse+kYgF
1vSx0dWnTx5tfq071Auc55jnJv2LPnWdJHz7V66qoK7P64c0U2cC6h7XdWPNd4ib
WBLZiXy9kD7Q0/cMZVEo5Wr9EH1uH6wtTSTZlBNVQj0=
`protect END_PROTECTED
