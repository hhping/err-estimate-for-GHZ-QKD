`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8AQU5mobYCRBqIIuI7HVD958vKXmOST4ARGXlUpHDD8WFv2n3TIvNi7VOhfav9zY
tnwBN+zUvBOZ4fJMjgmxOhL3aQOkaCi1HK0KlvLHghBPIeNjJ+0CJ1Au3zgccsJN
kFjAa1jbYtqMRECj5tPIUJShx23Vlqp0jSYs7+ZQqW9JwIgVCcTsZTZxRLf3qr4h
Gi4HSToYpDRHd/Oy522ZR8o07JkpNMNIbuFtBbIiGdAffK3BcQ2XIXJC1tjbzJqW
xafhKxMdB2wZhCZYXM3xGJpOBvucz0y6gyPykM4T6zfuXt4mAQSv564xQkPkJVsb
EbwGSnpO4eHpKRMqBUIMChJfGkcwl3bugv1i1GhvQCCfun/FoK2stl0DuV1Ojxui
lO3eGz9IxmIUAYglHa2/qtqQvZ09+fSVSPaz+efeTjwHl3iiHpCo2muWNErwO6DF
ulNmTR3Qe+FhMmPA2egyxnzAkTXN9xARXzEbTg0UaeS31qZwu9DhkJPzN/pOZaDX
l9Eh6tyAfB8+2eKLIdz8NHsNkKDUizJVtXReoGPm9AMTC647VsJrPMV5W0tNMTPG
ue7DLKNb2iXPvmavozGIBR1dLSb3HsSOIq2Iw+4KwRvvi83z8hbdIAsTeFNxLFyZ
QVBJPNmj1xBqVXiEy9zzGgKmg6wYoJTV+bdlMOrxQdn5cX3VBsn9fGVqC+PRAqHT
vPJItdL2H/9MEx7E4GirXnR9p9Qcz33b0ujqiR1gBM8XCJixqDrdoP/6wQ2put/4
jc9ZgiyoeWSLPkNsT4WH7ckk/r8Se5fxuT/VyCH2koYrFwP1KEjmD1ZQ9WYBWUnK
AVTVYuNkp3mKufL0ARu9CykYBGaTS1NwdlLkzbb7ph+ir8XOvVNK+XvddmCFbqGa
KcTy0iBU4QKuFu2eF8LKm4Rin/MWjHp385PaDHlISgMi6I+lbQZJ9cSxjbaPjp64
mj70Lv4MvIuDm8cgP86RQdyozzrc9eQBVqRWOoHjtFgh8PlovHEvkAeay94SYi7k
C5lrI0OERff6wu/2RaNvSuBOKJqnrbPAlbV4b0kWnUsXVdFTD2yjtjvfdIW2OFDg
prU3zrgCimV5Dx5myELiPoYH7Onkic0Jw/0/mlXr1JwHi5P/yBPpDBXDY2+rz/3j
0wstkvi1hZ6PDmuK3t5OR4nf8NXFp185eoMCyuADplWFAXQCpGE6UUMDm1g70jHH
e5u9D0lXH1hqlLWZNPeNhKfHknDA/zWjwZKv/1G18WzqbGPJgsUHKaMZygy/N6wY
AQiSSKKr3t3wfYMvIp/tr0O+CirrpBg7yEIi8q0TL+mY2klaZJRj/jhSgOQMNlSj
n92H9Y8WmeuvFkhyXnbHRWFNZQ3LsukGq/r5PaH9WZelCleOohUh2eFhzNHXtS2U
zssdSpl5rT+QowUQ8KLoAxmzW2WEiBmYEBJFUd9ILR5ajiAIlMBypWD4mr7Ty8q9
gg1Fn40b7lwaa2PW8QVV1p7o7hWjaz7XCD6QBAGce+1cGki9N1JaL9tINLz5yVxn
xGfTsgq8rfzMdf4v2DWPHX05oUE3DCWSRYu+wKWMOSsYGIA6HHLr/LtAUxVVfNBe
l9Wqy89BRDVaF9wmQrqjvrh21hOmCggIBRo8W1lvtb9a4Xlu7KZkXxEJbuYXepyk
Od4KMMhLBJqvFieFM+D11xPAiSm75hJxLtwkh0HQaLQNJVyU8wHEiUjRohVbvZGS
PSyjDdxYAijpf/sWQ93EJfIP678D6wtki3TZ7d+G0g+EvKvfwOQ+yX7MrUSo8/tD
lUGocX/huIbdoLpIUYz8R3m9efN3SvS/K23wUDferKpkXfqYbpDWS7aFztums+ge
3/Ly8xluxDuK4VndBQXhqPGzlNqY6Ama8K8a47ICoVWpu4T7BvgoxZHLEi6jq8J9
l3sO/hXweiUIEHohveYwGlQEkNMizcqYe8lVC6vpZq5QwAuBzYwBXiTsbTcTaQfs
790e+LwoYMPOph54oJSnvAnvdFRbbmOHnsQV2oDgizUK4JuyiR1TsZhHKgzA0GdZ
FNAT1gb6rETelrodo2WMDmXJFwglFhMZy0Kh1qj5kxIOO227i6bHW8Ow0JzxkAD9
9FFh/EdeK6K8i/XT07wj/0f+BuDphshvmk0h2NBmSctQqfhEFZhXCdtJ9fOTRNqj
xn9ZbbiuNtiamnWVH/GfB3q8ngaHbiDZ9/ysWhb6GMHbKSkVkZQLZzJc16g/D/af
3JohwvJNU8WIR+mJMBoy2Lm7Qh04qmgXv+KYDwS0wmiOnMATaKal92OBhvZlwsuu
5L0gSrRSL3BWgq5tk18a2+vK5BMdwtyG1e0GNng0O+XQqnY8MzgvuGioMghfUyw5
4pHL4RI55m8axP5MrbEZSXrLKfseO6MAjQSXIeMQ1EWvEk9N3/brvMCa3v/BruO9
2A7XQ7UimDN2iKNIkAdJHqJXNE6QH3kr4x9jEgbFOizKYop7VkgqISUTvw4J2k5d
J81iorMQU5TNLBl58LFjeDSjKtxPD4xAycDNRUIcbnrZIqW9yWvDt9QsCkG+7+BB
iwecgxeIVVKbnwMHahOF1TU9DMgmSSWMFmad3u7G7a9ibou914zCqdW7h7c4+DAe
ojiktf0U1qE8CCz7eMPm6SOtOVpb3QxFVXG27GjgC7jFQcIk7OoYP1ah0zHe0Lbo
s4i1ZHrTGOItZUFhJOf2g+cF6i3fKOB4+YCMKHF11XiMoth41uB+bCk33BpJjt6u
tn0K0Ti6ZMfeb3C4mnWVNf7gcIskN+qyEpVEWfQ00rZ9XAnun9zIN//DaPTFSKn3
k3d5i0On9/bt0bmS4hkf7ePDRdt+5s2jaW8R/1mx5O6h73eD/aBSK05OFvGwaOtg
p9DEXSbXquFELPSz8U3WE8oJfeCV06OZccZc5ppJTS82Fy2vL0QbDSEHEw7X59JB
AlhqcJunSAG5yg6RElDLe0GTY1j76zqNshJUeqP3p75eqGH+lN7oX5ETSV7oIL7I
E825IkEDYGdBFI9qGAY91toEs2y4c1Q8QJIwDu1mtn9wQR5vJX+088/pjc5uOJE6
L1TZdC/t16unBOzD+90/FlHmUtYv/8vnld6HbPcdQMpi3Gc73wzfR2T8Kee6Kq6N
/PY3R3rOVcuk79EptIYW2hAIBHqoeSnKcOil72qvpGZFBa2lANoJ2+LVxyyu/EBg
A5X+ukODYeo/Ll2iKN7ZHYVJ0+WGqTOymetFzvXO7wof+qPcK3Fw2V7R5Z/1te4n
iVcS5Duyycr2WeljT1JCNCfbPVgWh2u5OSJZIXduWP6D7sEYdJFhqKDjZG8SUj1e
4rStTg4cSSIOCYZa0lUfFTda38Edk+bfzjf6xCuPAziySwTN6CoRlZcJ7vCFgur3
LdQQ1SMGlBEVF02jEOEZKDImXrlYohegTEgJ0rOtkfII+wkjQW7++WT7Xs2gy2ge
jcyWAIMx2l2z/3QuSbNaACqIRYOEzxOwzjScegdW6f745ej6r+YTKVWWvDdakBW6
BsrsPjaBLQjMCYBGljvdQEfUV+v7cOd1Vipz5mFMaNw+4024vqP0InQe328PaIf1
d9R5gAYnCGs5LGfFE/M3nnPsD7w1Q99IyIDDfpk7gSjUIsXEZvJd607ikY+oX6sf
M5jsSL8OEmTeJhTL3awBfKA0XeznjmIyR9J87/70FsCfqPtFUu6tKpvHVbIGUJ4p
hrtH1qDy7GV9wGZm7qraoSgh09To75qUiyZwGyFSjJnOgqpyc7VW9DPAjqBA2S9m
KeCuxwv0RgItIDta3M+0G/86BLq6ibSH2aYKy3KeXphUHI/viaitEp0+A8s0tDSU
`protect END_PROTECTED
