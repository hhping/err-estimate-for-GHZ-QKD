library verilog;
use verilog.vl_types.all;
entity ama_chainout_adder_accumulator_function is
    generic(
        width_result    : integer := 1;
        chainout_adder  : string  := "NO";
        chainout_adder_direction: string  := "ADD";
        accumulator     : string  := "NO";
        accum_direction : string  := "ADD";
        loadconst_value : integer := 0;
        accum_sload_register: string  := "UNREGISTERED";
        accum_sload_aclr: string  := "NONE";
        accum_sload_sclr: string  := "NONE";
        double_accum    : string  := "NO";
        use_sload_accum_port: string  := "NO";
        output_register : string  := "UNREGISTERED";
        output_aclr     : string  := "NONE";
        output_sclr     : string  := "NONE";
        latency         : integer := 0;
        accum_sload_latency_clock: string  := "UNREGISTERED";
        accum_sload_latency_aclr: string  := "NONE";
        accum_sload_latency_sclr: string  := "NONE";
        port_negate     : string  := "UNUSED";
        negate_register : string  := "UNREGISTERED";
        negate_aclr     : string  := "NONE";
        negate_sclr     : string  := "NONE";
        negate_latency_clock: string  := "UNREGISTERED";
        negate_latency_aclr: string  := "NONE";
        negate_latency_sclr: string  := "NONE";
        width_result_msb: vl_notype
    );
    port(
        clock           : in     vl_logic_vector(3 downto 0);
        aclr            : in     vl_logic_vector(3 downto 0);
        sclr            : in     vl_logic_vector(3 downto 0);
        ena             : in     vl_logic_vector(3 downto 0);
        accum_sload     : in     vl_logic;
        sload_accum     : in     vl_logic;
        negate          : in     vl_logic;
        data_result     : in     vl_logic_vector;
        prev_result     : in     vl_logic_vector;
        chainin         : in     vl_logic_vector;
        result          : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width_result : constant is 1;
    attribute mti_svvh_generic_type of chainout_adder : constant is 1;
    attribute mti_svvh_generic_type of chainout_adder_direction : constant is 1;
    attribute mti_svvh_generic_type of accumulator : constant is 1;
    attribute mti_svvh_generic_type of accum_direction : constant is 1;
    attribute mti_svvh_generic_type of loadconst_value : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_register : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_sclr : constant is 1;
    attribute mti_svvh_generic_type of double_accum : constant is 1;
    attribute mti_svvh_generic_type of use_sload_accum_port : constant is 1;
    attribute mti_svvh_generic_type of output_register : constant is 1;
    attribute mti_svvh_generic_type of output_aclr : constant is 1;
    attribute mti_svvh_generic_type of output_sclr : constant is 1;
    attribute mti_svvh_generic_type of latency : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_latency_clock : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_latency_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_latency_sclr : constant is 1;
    attribute mti_svvh_generic_type of port_negate : constant is 1;
    attribute mti_svvh_generic_type of negate_register : constant is 1;
    attribute mti_svvh_generic_type of negate_aclr : constant is 1;
    attribute mti_svvh_generic_type of negate_sclr : constant is 1;
    attribute mti_svvh_generic_type of negate_latency_clock : constant is 1;
    attribute mti_svvh_generic_type of negate_latency_aclr : constant is 1;
    attribute mti_svvh_generic_type of negate_latency_sclr : constant is 1;
    attribute mti_svvh_generic_type of width_result_msb : constant is 3;
end ama_chainout_adder_accumulator_function;
