`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjR1x/qHSAYWA9GM2BzEvdxhZ+Cfw0DcbjNbXh1SVh+ZKWSlxBmsHjueOie0cIRN
B8KSKCucjJDyTlvKOYWmVboib6K4C4uhyRa2oqKMHhZSVrZ/ny+V5a9XOLX6gXgM
tjsUVAsON3jLT67nXTJv2i6TAdDX7YHLDhaNYpQfYVZn2sXy6MMDvAeiJ/PBvjD6
pm4c2xdNuJexB3xpZzgI4+QEGt5DyX7OHRlekOJkwC+WR07Fn2zWnbwk/ApJSjgo
h+vPPTAzSG71sgG82VTNA+Fo59s5ibGP56rmOtO9SZrlxiXPdK3T82xUj6qudVcT
pdie8uU0quuYxGKQWyTL/p2ExFd/PN8+1H868B12Zbvx1IFJdVd3DjQ9qltpDYHj
cH4C7VnbHmF2Ppigl57I0Jp6wQZkrQHta1llr1QhENcLge1y4BjQxya8LSMtbgkt
b/TZZBlLgQFgYQ16PsEOF0JggRJPZLoqDdQPVQqLyejQoXXwCQPNZ+sj/D5qvHOK
CTBfhs073Fw1pYk7Rf5khyiEl/13YDl/WyIQPtqPQfy3G3Ahw5E+u9BlqbnEJon9
MktnBiHdBTISEVvCqgHsrtLvJVDkJAmo6QGYh7eS1stdkLeRP25NaPp4v8VKteGp
ac5SfDHSuR7bPImSD9ZghPYp+E+JVbcnvEUmlQv+2hiixZhXpsPIu0/qLhM7u1Bw
kIh2A8eu+eo59JanyP+/aEwMFRhXDoS+eb1bn6vrTqUWFWwf1V661+LvTk/sBXVQ
7IxbUXxfFAJ+FCNVhP8M0i+4jT+GlPDvvVhlmjEUS0A=
`protect END_PROTECTED
