`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohEdjmKH/RNrWMm2sVvrFK+ALwdNmK9l71OmMv3Xtlh4q6JnoVuN5beYqswLG+PP
BXclr6Lmo4+Cw7XwN+BNCJilq1dEmRh1QnwBYt+N1jCTK1iwD8Hh0QnFbWSfT/+x
ZL0SQM863rF7J2U4ieKB+t5tn8CWFBvsFW7hrREYjXO7wvNZWc5kfG9ohIglraZs
8IwNNBMDEZK01wuSvGSbZKlkqaJDS0VKBhGF14Ekcru0u0Zd5y/bih4N6516YJ3+
RiDneoGAaqZ2blNjNyXb4Y+xPLHeStkRC1jt/KnsgYxtiq97bf2GYbzpwSCLABia
cqwtxilWZ2bch8vo6dLIH2av3waTZhKb0Bl5VmcH8fbXi3v5FOUvpnzJjP+cvp1Q
HtYz0DTyA1dmdfjhX/a596/ZWvZV4wx5pply9LdHGFo4zi+DIT9KvmK+n1dnbr1M
GL0smE6MzQUQsvITy6+D2oEOX1iavdD2MnuBQtW1QjK876W1I5i35F/vya1HTZq5
IdlvrJFWlGFAeTRzeZQsUJufpXbboK5s6QHtMarapv0iglmSRHoSbOmA4pFrlJnA
iQTnK418VU/DoyKcLHouTfCp+F1LhIx/RapOgVTw6Eolr0rCd2fdtNOp8kC8ygSZ
jBeqnBgrZKwg6jKw+O3SpChkQa/0ovOcswkzmbONLmo=
`protect END_PROTECTED
