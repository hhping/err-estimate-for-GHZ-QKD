`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uDjcMBjG+FVEyn4HCA8BNYMkewRdzaQrCKSEY1o3j6qQU4L4CbsR/+SBO+GBuCw
plvO82pQtofGnfeuBarH2AQxCwkVbMIhTFU6Di6LaXrQgzWDSIXXdzwBVTFk1nbA
t0/7nUjaBzs/vB71DUyX9w6SGsvcOJSXXCRt5Pg5LKAEjDG31wI7LoQloq0t7m7d
Z08J4er2Ole0GhrkBm52OX3Q6evqqgGl708yrvrfA6avY0QXpQq8xXijEpl42MBS
pQo+e7gpF+k8S35KXQiM4asACkQk1qzNRVYshrBMAlHEZFhyIQrq3Xohb3wPMmyH
HMRzus9PsK7Ng6SqiCgLSZHUq1OdIDARJ3A0S9C6kmtrHEjOXWaIh2LyRXMAShie
`protect END_PROTECTED
