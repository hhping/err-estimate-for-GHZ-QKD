`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+AVjur4kwN+MPSUjg7ziAx5QHwduzrR5OzE6cHmimsfXh77RKotZSlEtjj/hTXn
FRMSj1XXeJnnQYmBfV3supRjQB+Ka/KAuSRxWXwqUZzh0GnOG2ylycAssJemXq+3
qyrYnlM4nC5esXOr3TUjLJ/kEesZKh2xCs/58fa1lwFyk1a/MLxNWvV71egSFmiv
AeFLnSRdek1efXKanKC5yAy3VTb9Ch2hnY2Gu1dfG0q3bxYE8CTgTCAgPZhSgOag
Cw4eiY7OMErR+7T6CfhDyzVyDhsrMA6g1A5Exk4ajvi7f4tRlcUV50uvdzf22Y3z
5y2EH/FmrDvLztE0lYR0LKZh9i7lPDSHbw7spu5MOknVfccjvwd/b97XavGjcCum
DAB9In6zw38EVzarisFmtkljfw1AOG60/2x6qcL52EvfeOub9E8Kb5ZMdwZalM7X
xgOgATHsTNr2xhPNeUtktXlbF1hEDFgOTknT+HrGDIw8V6X94IaCTdm7f35wqTqZ
8c/aDcgYrkKoZC9M+JJ3LuGsGgWy+AHIaH83+MGxHpWymutZmG3hJWHqIjecvQ8e
VWmMk+9GtntY8hJ0gp7WW1JGQrPDXqYAqK5b9Yy4sEg6WrJwFfFyRUcvn8zk2s3+
pNygAR72hL7L+JpygtSGC7fj04MFqy/v9dkhaucZE/jimKauMl5YEJoWBJrE+xCq
2OS+0tUmeNVCDSFeqEEGQPdcmHjEzLBf79RcoiKLzTOSN65YGpfoFYrM3yiWr9ao
7d0gFY26AT0rnr+W2aUB1fl+gE10wXa5bhscuWE1Y4CibMVwuXbVz6UE2RAXFGPC
2p2TtItZCNLJlxNXNTdC7HH17ZoM5noAG8FrjtsSGKE=
`protect END_PROTECTED
