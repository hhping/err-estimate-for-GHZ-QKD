`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GxV1cmkzTeUiPLNA2KAZHyFg8jZs/YPFxYgBI2ltoP1Gjn9jYjwssDF/BD/h0rwT
JTS6hxffW+BoqU+gLjVW5yCy7A4Ralw3NF6EHAo7u2eDR+sv56zBXW6EcxG16yMe
mNoh4fVFEW7rft35Fda05joc9DgEUIav8MfWACQQSN8+6q9/yJ9J3GPVN64iFLl1
oeCMIp10aC+8N0dZQ1n1TsVq4BRuz2/t14/6fGY2EhLMtaitsvbCGyTVaQ49mAvs
DU1WCQSwVROfI7q2GblIm8hJArQlR7ShrPR6edZ2k3lTBKcIsqCd0054zgzn0pJv
rA0sQ1WiJoijQQEKUqZiM8tkO3swdz+/L8Jq59uRhZQV8iR73R0IbHWOFue23KZh
MgSrgO91uV63elEj4Q7nt09xwauLxCmyIiDbEYExQY0WuE3xcILb//zGIx4dxfaj
7AT4+M4OM/UAsYPEiMvF12mUAFshIKUuzh8Opk9N5AXANCo+sBPvKKnNz/Sz87fj
4Q9CpaaydSjIjSGDUwdp84s0DFNUMeixPM1zmuBEkCHouQfH0TtMlYOq+4lHkR9U
QUiOFNhBaosVCHbFSmbbsT52vDMjDmgfbs75vTT9lFUGEc+QlqEjObsQobQ10Svp
WBrS7QEdxZZ1jOpoc/SpsSgjtsbVSew7u7zuCu0R0pP2jqMwECxYH8cDEiZJHXbZ
UIUkUob22hiYurIcb2eLXutPjAfkmO56zfFEX6fY4aAHc1AHmC3QpyXls4ST9CWS
K7j8O3J/8wCytDq6hDufU33QZvHy1TwgZvunkvOic6eC+tO2HSFj+8Lf8pZHOYZe
qnEq23MwEH5WutYa/b/yQNTi3zMqLPOfBtYYW8SgPzKdIPBnOn0NRs9AY3qBqf3/
amxl/kbwK3kIrb+LdzK+8ALnq+7ag8KIXel/q+nDRUgORcr1DMFvQZyLAQyRsB7+
7pZPbkyKMHrHG/oeX5KCrYf2LWvtkZbagmdodC7nDTEpeyQVqEBmJ02uYlWltuoZ
gvew5HNklLpw8lSvpcBMNWwOg9aw4pYrUqZQR8rfm2f9LbAJC3cBZtS3QlTneU5p
wyufdDGITeIGMVVX4eaUaD/y2+27QA3AzxRD1cHhpCcR3JUOu5Okk93cS0mIu83r
y4KjsFo5nFWpKz2Zi76UvixXddnpqyhCGN5rSW5Py0u9lAIuT5Co+u+fATY/eLf0
57p2BIRsPaKFbbqlakqKOdWmyl1k/CL17Uy9JGgq+q9uJSeICm3omrjZ48ruvWHZ
TS71YMPIzQ9z3bGk2QNHhDzbtima3ZTL5c/z3Hms4XR1htohTNccVKLzyb/Givne
mpnFTbjlrcsANDEgj94woIg+xpthQrvBk04SNEvo0VXCo+hMdbgl81zRjQSFD+DW
Y5cbJBa2us3kjgLs0bXXYrTE8w7G6V5qsi+S6rF6RJOUbOgRr6+PUt7LgrG4PGKJ
DxpPdGdRNSwyzpySk0zcb81h+FIMZwgRFzhL9q1G7Z7wJn4E1zWyVGD2dJOy8+4K
no3qrY+Pxxh7pQ9oIRMQFgTAYXYnI9DsjMGiEvkJ8mKXwr52JKSCupxuxt1u3GkR
gv7HQ9hsRXLGUskLALhUyOmsEKuXTlGGDJbpPS2aukGeHr21lk+WC4rKFLV01X2Q
chu4zy7fJE7zAg4tuNSjsoOIY/hfc9fHZy2mBMKzpOVIMWzfWQ9S59qqaFut2lku
jkxUETYCisqS07hCCFtsRzxfe2jJbfhlvTBwyAWt3MdRkHI5drBZhgK0tGxLgpDJ
GXIjyP4z9SjlgKlRlkoaWjQFGLjayWGtxoC/aS/qejwAg7+X4m7f++9HFhjiInsn
kUNfBg/iYLMV39FYqKM5PdMj57DV+KBMj1h14FT3o0GR0yz/rKGKBCZzQu2qSamp
r3IS+74wTlD8aUpGQcWsXfO00SbJ+xEXFGAdSEHdkGxvSltByFoSdMoCKWHWQgl0
yPpQCKH+BCC5VGAUOBh8+mLWQYoNkD26tN+OEHVFQo2rtjGCY+0Sn6HI580550LE
9ZuufFrxbp4UMEL/0NQdUdDM7CjM3c9f11KdwgNb4cet2TS8k8rayK4clyYnEoIA
4vUWqhLLpvZYZm1f43OitqNg3TkTp7jBRMq+K3YBher0sRqzLZR/Cs3SCJQXw7Na
ypi0L7mWw8276uSvxVziQF9y9IydGsAehwKxGwndDLNHKg8f1vaMZY/ygb3U+S+B
p1yy2ViVN7j2MjyLnTRRCl8ZKfjyOtp2m8VAEkG3X1yy2TWeNNk/G5C+tOpIn9Wo
mW3ngDaRky7NXaEMYqojftN7xSGU2452cOhK78CNCe8AFwBH1GtCfAa1WvcR+3xO
oKZsUAcDTit4hDWpOP74nWGLqJ6Ur/Ft5oNvFGxdE4V47sZTpo+QIWJvs021vJ5a
+jL82SAlViDHAn5RwGu6DbkPzzai80NyfhlI4QFEofWxbeMpLMNWhKfIItnS8p/A
t5YqkKtnqTsy+FyH1eldytMcyGdHJZOTO1ropgAOL1RwK0uDxZqHiDr1w/WkHQCs
/6K9SpjXb82JiiM3RGnBDjYSc3WIfmx7zNXHAufU5dqSFVV9JByXtTQrifdfKV2+
6c2nn16guQ3zHeolYle/9pBiN6/kZV83FIGdax+YELhI0rSUJDFX7F7RHmKx1uWf
asr4F/+EE2cWvrRZuD55sXC4o8KawgoAeUM8f2RZBMgRPFEUhqJRN+THDElzbDmO
L5m1GsBcgan6FsoO0agjF/UFWuObBq/VaFRbkd36r8b2DDKExSPzUmuj2Kbmb0vs
QZqDRIWhu3LCrkreI/ZBqi8kmOCPFv0PAZa33r6Ryc9P2oYr1mGejGnHEA0BzdBf
9eMOJIF8c5h7gdjN/j6/oGo07pbbmdHpFZwCHr+/XGxO74i2ryjiEH9AUQ59HMvb
s663EimztV6qV8osvmWqz3uySETZxqqfxjMBD8gq0QlsGOIUjWw4+X7wgQXKLr0C
+RTpWRtY37LYXH+olnx/iTUVtIEEYdyFWMmLbyS138FOJ6mQFsGt4R0a+pHEF/Pz
nmuKO8wWMbYYpGFM9Kumj/JEVpzRxrq3O369jAB+PIIfkzQtTlragvNcvjjVGKk+
VZLSttRva3uO8zF75YI6oP11IxjDE+4W2yCcdydkxDeOHjACAG1ysJ1Gz9qhnoTL
CFHkHwQvhOvYLJHkkndCtj+Y4eB6Nhaobods4sbAo/8ae83qiL+FV9xGPQQDCDA1
rn+q2nFIIlEXRXjRaZJi8S/4S81qwoy50MymoFu1lQ2KcxVSGz8TUhXoAhAPL8wW
QH4osCX010/TIZ9HGvZtrXvkxrrulk6l9zIIsanshUo9VqRLDdgKdF5r4t0lkZdU
ywyynBnvv0b+UuD9iZTYV8ikFj1cbYA2ym487k3F7fjT8rIm/ln37Ev6reaF3QNO
ehPLdnnzDPo7ZqXksFpPtzTpExPD0dY1rk9AVzC8EmTOTYl1HzHcXPElxSAtsiLr
K00ylAOczDLyJcWcB6BWKeGq3L0Y++NnEiQkXINKfIsbKJHJW0T34VVvkPuLPKve
UsW4FM/h6lbZyn7bMTKTISSUrkA0YcZ04LCu8vrclBLoKnwzQ/kJPmH1sHRovz88
7PlERRIlZJlbHXmBNllANCBPEgc6SF2CYt31zxISjHHf67Or/MdVq8ndNkwnHeKR
bjusoEVgB1uQotWf5Ens0V2oEQA4jwkgTDb8QzJ4ujQPaauWO7hZ/sYWwaCcDQKt
q8eK2QLy6T+N6uKm/1L8BOyCZl4MZs/yCBRAc9Go3BB8+J+9B6iKKSSzU7C02Dat
mKisoT593SWIqL+Qq8PU1JoTamC3F7ihxTHCycvOi1SkETrCnxX5njvvjcgQbx6u
HD4Gi39UaTOX+YiYNrA/maeBPEmjBt58ks74EsOKojWfwWF9PGJiMezM+OAXVINe
oicHweRKxRhDgPKZNMk0rCnJrvNx+PHGnPAU2dH3xFT+bUSUtPYhb6KZLkt7ieNL
/tXyZ1I/c/MOvWlBYv7CBDrDgBedNNl2/p2zjVTcCW2Hj0vZ2uiLlyE9auvhx227
MrGhqAS0el7JV+YxMs74VLHOsNmIHF3O+4u6heu/13N6GPzyeO8BkQOBzvfeKtnZ
0BjzuC+Tu2tJ1199U2LJ7UnAmYDQmjK3BENCXlfhjtoQ+rL2xCPlR1mNAxn5XdAQ
D+CM8vTCbs4dGeDA2JA4rv+sIStpV8MbQpuyIopY98jqeMSQv+IL7XcwLERxsolo
twQ6QJadV2tgkGhYOMZmN0NPt9xTNGkTpmXExKrhQHafIibvfeenVD3GK/XusSOf
CHOvPrw5EobLCaNKHeUb+0AmNRRyvkGegvxkip23nkUdDnip2V8T+kUF4qp2/ulQ
lwUaMYgc+8Ygh2jUYgz2Y+0UqZ/yOVHsPlqphtdOrIww6trYAmkpC0gMnBvIqZaJ
aPuxEstlRfxbE98Ev+iAQxsMmxrHyEsaSR1axt2ASy+bWlMz7QbFxqld4CoQCvdf
HgmiACP+DNR0G7fTH61EcjUaxcfH2X1HEHeKHhVp0rgX2JlZK9gDtThw4mcNwjHh
fAj/DnL+/BN8EXPaRcZ4OZmckiM+Uv6IA4eMoONgXoLRIZ9QgMS9/Sp1syL4priL
a7ZZzHaEvzc3IqEwO/4V5PN4EGC8QTlsZ0LUFc2log3Kl51uOIHr9atzteEAKUSW
0V5ho3KQ905Q4h8HK/IoJx39oECuSJXAC3EwX8aGVwpIVaXWQbBD+ilgBpZph4I9
KjOylLqEWw4datIurLA101Tvz5GKEJ7dCdj6h3G5O9xWd3Ha+KcAJ67H0Q/BAynp
FdGPUL94vkXD81PW3CTG1SjEIxYv1pZnhj2/kFQCNOcmru0AuYogg0g+l1gTOj1s
rCLDU7yG+B0P56vB3TtxqHWgxaeed1aQ2/vvM/WuZ1/Lkwpnos6aEqNu4lv5T0Yx
GNjFu8TA2Gm3OTjIzgFWF52g4Aiuta74sctes7uVJfhlwhlDbeM2zlY9NurwbUrA
kL0cJKBFq9/WJ+Z6C7ffZwe4EXBcxkUgMhX+CdGYfpnWjABVxq/Ocf4eBXRcg6gn
l+6jpDtZrHF85fPz9yYTsq8bCGjqVj1Y1IW2tzZ2HBMleMQg0+Nve4CU4hKfnyeR
Cp+2/yDczKjbCC8FIV9whVYPi/qsx79NK6CWmG3DA1KImoK0e0LjTHin2R2X3hhy
JrBaWFnMYhpAPzppD7Rac5vaVDqmotTyG+HE5jWL4pC4xdUTuKC9CK9TNxQxFyp7
t18hLqB00MxUVmhZMDj+ol2sfMOmNT72kNk007aDCtqRRbS2tuDxRtyH3md8BSuB
gCcVixhtn8r1lJ+Zh5UpkIU+BPzo6bn0erugsvoxBLD5NiQKKypcwlvoMkXswssX
lc1Lg80RqI4tOtXgAaiEWT7Sol3ccpORqdy0pAl1SMfc25hGQNlgEIevSkbxwWEj
x+CjqwaVsT1RLXf3DBn/wb6E0mIkbZMT3Nz5B75XMduANbs2Av+hUmT4M3FablZe
y5NOC3Ei15Eiw7XUsacWaVG6fMk+wcKPWxzMsn4wQeh/sWrn6QMnGIsIdQa7Z0i4
Gzbm9NLKlfHjDEbWpXUjk9GvwLZipJwEKiCpzTESixwIikB7aJvRcI5frtegclyZ
ST54z1kc9w7t9K8+oZWooIRIfLUlwiOzYyT7AAqgNon0evQtlW6IONYiS3vHpDmw
7BcWPZpC7MwgJDI5C7ts6hnOx1EbVK08biMJSXp18fpAM+zJNFQDZGnMWkNx0h+O
j18Hz0zIR9VIW31OvzfHh09THFdJgBTjGUVhJGhqfm18jHpL2UxoVbAloLiZoe77
G0pf0nx9cMtj6SMibaypBpF8gZ8m0ehScubbgbQW5dhjm9q1HjUd9r2syuQW7UVw
9Ghs8YvHjCt1q1d8smPQBw+s59nfeDCbkOFBg7OcXsN9Yd0gcuGE6wsJhLKjPzlG
8jRC1NRg4MR/6QlMCTu0vQIUfrUPtQEUcAK3Feg06gelHALuT4Uqu22EHZFxfQWa
/ku3I3enNDfLdKSaYxjvXRlgpijTuZvjS/SAIg+S1H4YgfDJqEMmT8/ewj42+2Dv
pQG2/shs9xQUt7oPFTao9tk+kIQZ+MxGgj62RZB0zEuhghtd+Man9jjPhyOwdFtb
8X2XCfkyKnjTD0Lr8S/mPjpdmomh1bp667sokQjTDIkq7fxQJ/2efr/Z9MoVnKOF
ptk5SIkQXuOj2e0gj/zEw/7n7of0dDaAwOm/JS0PIW/uyZQwORRw4/ku11WGUzqB
3tXcej7xMFrmRS5H1TTMfuMJA+DyI0x8xJjcJgnFlnpLP57QYLiPrFJfDGkMHwEP
qyfvQfTnzSCXEDU1i/yF+QiR2QUGv7TyyfE4sneUkRYTVVNcs6cRZAtpWShBlmEJ
jxyQItnQCaZozyRb6pk3ITymLLWOI6y8kriCrxsqG0076UPECBKNI+9ah7GKSvBX
0AXbKKorTbUmZZ4V8Rdnp1GlIFlejNaUHxCjVfPjXHLXz0VEC5CXhVAhvStghOXA
ZLYieQEb+58w/or+KOuup/IArGT69MtC2Xr6N+Mn4wTEO0psACv+O3p2f3RgcC1P
Z7cuuxu4+9FKBU8BggBr7lmy+519gB0MKVRGxyG17KawrE44eTTqYfQ/RtwMCFtz
5ajzzde7hBtsaXhPMz67OxpNs2N1P1aZsnIHU9vXYkcGqSiIZAfcV8fSv48jDfqO
izutU2r/NJZmFi6yUkFrr9pIgDH8jw+o4sAzNqKq3vHb0UycnNlWjUIFeHxcqtsY
3Y3lgMHqaOJcaWTUwQKVfVbbwisEK1YITsy8QWL9p4uQABtY+yIS8HFrQ71YrKP7
Ifv6D0mIR6Gp6R4iGiOKtC0qThWu5SZjsA8hfO+u6q/NCBGjOhTYIUU6eLUvUX8R
T3bJ71mdGPaaEZPZPDNh27lcK/1KPOowlQ1ScyN93FIQdVKEkPWr5A7p8kP3YZU2
KbJ3VvX/cin7mxAR+BT1xA==
`protect END_PROTECTED
