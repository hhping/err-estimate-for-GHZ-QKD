`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjVGWH9+7mdcYHhigEEcIEdcPwn5o30U0FN7Z8t9uWs1ttQ5IblRkzk3+Ij6cqVX
KIzs5KP4A+g9/BJAPyhatmy39jVDPWqUEe1/UZenGoGQV7jkwSpZR+ZWlRXTxsRC
/7J9DpmXtA/Sfwkp6fdamlKYJF7v9y4+DlBFv3xwyZtun98MwFRC+eZrhfLe9B3H
+d631V/6JH0QBwpc79MPW1quaSWdBLzdHVGU5uP4mbKMpX9HuVJYSZlWp2pLR9Jp
FPqaXZShU6mPgQDDnlV5MZ0vNQ1wOeDTGsDxJMHOg+hzXdPn6c1ujQc4UoUs9k0D
lKeEaerDHltu4hHMi6aYapsBtaRQswzUol+CEocp0ytlvqEoGQz/iNfJe9u7m4m2
D3cXoaqQTOTBnaWKFNhK+pOXJFEkj86lyoTmlwVvlnoGd4rqxROPOHxSs6t/ggbr
yFGBA2h0kiDV3vV3H8NqGZAnzVkAW1t6hju1o8OmB3oO6EBjP5CIZNhxCz5UqZDi
uAJFPWOdiw/scNNxf5mXlM6pWNyc7yftNXx1R6QNug2X4t++TQeG6O1hbF7fnsED
BIWJRS5BL10nOCsEmrlbQ1zuwK9ZSII/fSuJTGwqSAgt/rry+muZEJdlNiGotiuY
jnHmsln99izunX7MfyqwrkFx/lIykkoRKedUZk9aYcdFq80rOnfz9A3I0lmDikCH
31taagD0XrEVSZyo0TlUT3h3PMFyHfpMXJYZ6w1XsevAHt8vFfZaqJUdc6IT5EXP
qmofZ8OQHYdq4EsBxBYbiLwLk2sO0PVA8tnQOWKg8eDjFjLqCf7Iflv5Lswz7fbl
ibiKqy+HpOLUg43xSmSogADyvoLuFvs+qH2/n1sjliYx2nl14jW5CLoaoPhe0hnT
Cd6v6zhKDOE+KN7RlTsxVkBINi/7PZriYqatMIC+eIt95nYeP8qx+BD9ltyJmp4t
1jv7wBvJC4GyRTqfcFijKLtwIw59LFu+rPukvedgkFf9o4PZuOUm2+unjAwzjDoP
5LNqEFvvFZmCz427VaIpI7Z+AyLzX9N8Qs8JJXatjTDkNt5TTF3E+QdP+5waDS8a
1+A071nYQ01fAlOLO4KRQAIWM0xJmEHvqQsWDX9G8jtGz+P95qVOasplJ6lWIhi3
hvSb8n15EHBCRmF36NvystSVyUR58ac0IC6QWEFaKP1viB9RZypn5st0xYkS1W9S
ap6oQyOOMTVFXil8jr1fRCjfhd9ZRmrt1G8jyzvW4bC1sOP16c7WyZl3Em6nO+VP
ZUqyus1AGqyiGhh3EWlimW/w3gvYTYy0dosKSRB4YQlC/49OgAmswHeJRsUY4knr
zMZR/g+AXYBQFydRWxMx7bsULPuEtiexum9Vu7J508bopls+uaBZ9BqsEvKa83bM
OMxpUAICdxaewD6FU/BWAQ==
`protect END_PROTECTED
