`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
APe5AECyhgxms+818PjoMiq/0k5nrPOl5KouDexQvN1yr4y8YZQSVXOYSDD8b/dq
5RqTrMochkek0X/ycNyAdde2JbyROiltrId5JmC23xIciOO1lTZj1rNmFceHGrXN
D/Ob4JONrda0dFQSrJPkVMHqoqkvqiGlm+bng/cv6BSBBCoE9IFO18SVJqO1r99D
uDs7fJAtsEFmbSyZNulK9NgG1y0GcBo5MLKlMGDZU86NzT0AEhCJ/b0hpzTHCCZZ
y57ZTesG6DH61V19TxdXXdaBAZLcnGLqZgdBZkWqDZ2le1INpkd7VNtNXcsvI2tx
lcL4t8UUFQJ8jJ+Y6EnLX/IMDnBrE5g4faC0twqrDFdPGmwmFCTE7g+WshsAWuUn
hJHZv1asK7X/tsqhogoI8ESkOwgjmKIHwsgkeYy150QqirHthUlnHSHgIvvAKA2s
u2NVJArsZQ+nXsFwCyFRpN0ULW6g4PfJByaT9YTKez+W7/sag1Ee054DReII07dG
ty1aNv2jpCbZy4Dkl7WgNYMiHTjf9P87Ga4KWSyuk9dZNIeR37b0/FkKIMR/VEkO
Jl8x29M51QIV7vGXxdRK1y9kJgqsMClfYz+ZBwUMXIdw5t5LDBkMdb1JIc6R/gDg
9MqZcrXFRekmqfg5ZmsX2ZvI/ieQUsEg15yhOfuO7CWz3s8A28YGBGe6lfrwSzmI
GkS8dAjjBF3BKNJ5RPz14ychvWIa7Y2R9tevyhwPTTOcIlHYovSXl3kWSGd++twi
b5INSVvrGh0BnNqJyMNBL57aXu++LXz3RCkQ50Roa75nT1Was9Hg6tg/Lzn/QJlB
h6YtS4N2PDqlHrY1zk6fCpg2sJVTJiAz7NDOF/vaBfYy9k5j8BBBh7OsxFqUe4LG
SxKN5tRHpl9ARec9Gbubgj5e9ZomI5REmQV/ihuz3B0agUxUeJkR5vCby7/SxmyJ
j4ax6WnFwkmWs4wLbGQnGtuJYdeaXCzE47IzCZscPKHCsSkCDd6X80SOpfv2UXh1
X1dONLxU1umgIgnZzVSgPNm7rP7vHFhc37Sm9vTXGs382ebyfYJeKQcaF9DHwLDS
OPTtc3KgjaoHhjuDrSt/Yv47tq2Bn7zY7vwhE7bORzFPWVbtjG/mH9ByaGGxLAbT
2omkc+F8bM1pGu0kiT7FhEsHLYw8vzxpwxxPkLgV1IF37lb5pBVU2OJGL5wKdhWZ
TZ2Qa1F42in4aKS8teBR7m57r5aPGBQUt2piOBrsacylta0pbde9Okoi/qZVmPit
n2claBxLLoYXRy8hGxFGvuMErJvdqVQRVutLWhmxqeVV2mNpQkSOHHx7NC08Mx67
0pzIhMf+C0eODmNCr3/wDPxKyK0rCSD8WFCAU208qD78KtexW7AqpTlkcIHxsbfe
aRkHYC3NfurjmAPIs8knEkg411+G4NhvZXzw4K4fn0/OT30+hUHxhymNwnvAM31E
6fs8bMCA/e7Z5t+M3BmaPvGvdBjs/HXh9qzamCFpUIBYVxZeSi2ZrEzU8SMJa4aV
aZ6Y0joAhZjoSu/TLBFFF9iV3RvSlD5prcrBSAkMqWHF9YpZFI7YZkjO2lpODJWf
xoBkXPmkdcvSmZL7noGOCVKjdIIWNMYO+C9NxLVfQzgGjBfsZeNrav7LKgfahABU
YEw2ZFOZh+9UFqx/M3TPWUf3G4b7SE+VwJgGlFW6HJmHTG6vPcOGqXfpGcWUaCcM
Hih3LzXNlVe0U3NzSTUSxlXDv+P69MXwb5iX6za5zjZgcUlAJAvQlwMK+RLMx/Yb
bjc0VZXXKZCGfAx/MLshFs/OPNtr1tU0xiJ8TkjwwPs54IAYQLf/6W/e1U46/j6p
kIBSOK5SjlN6dAaYfN6rVCEW6qXisQmnlFpI141KMQL9D1AfKTm6WPODk4dVKZst
skZqBsdC3Cvy0zpFpmR5MqI0V2/7g5CcQfGakqVo2nn8Ez5CjhmjtsA2zQZwKQy0
n9oAOwKhzyeKHh5qN4KURYI95dthEgE8UjfTq2Xzx2KJUy//CcaUxshnIg+UQPGf
ZuBeU1Xb8btfTJaSMvEZbTmLJOetTAfPr9m5GM1U/AWIRc0iIAOeGbSPXYfTWn92
GRCpCQ50k8kAvHsBjKRTBgxDN5KMXhsmLWRSkc4tOwW7ZAwBIEgwMaHE4OwtzOHz
RTN+uD+eugj7ekxFfaxbk35f7/9z5Snfwd10WGcNkLFw6+wzE5VpwiyyA598JXk2
TIUe2LkLfQhSoaI6ke86+ixAAZsDap9PBRvqwpX/j31bGGbjmyaJUxx2xsRmD0Fd
N4CFInSy0H/GXh8XHK7VkfUMHrunj1sMZi05ySYLrjkAAHyzbo4EHexq8Y2EOQ+D
IW4npuNP5wUjYE026uwoAoLJ1FWNvHiTki6GeovxB8T2STz20lPwLgmErwEuOOTM
gcq7kJxs/yh5Br/eBkHdrd0xNGHXPcOIof1sixrQlRgVm4qbnJHk5QlosLi29y1r
/paUdK2bL9Rf/4R2TiD8J6fcrWMIQr16pdvFiJBMVmKgAvBkd5FgYIWKeg9OWk5N
Bi1/7GXSPWYJhFuIL/a5yOdMonvLN0VpwmSSjobLiK/xLxyf8nuwE9J2rB80IfC4
DgtgFdXmY27ssGvqa1JgW9vrBypVweIjDH4gXRRNjwPNPeichLzA661eRQ8J1aMd
FRo0Cer4H4Pzlffm7vvHgKtDj+8xX2VJfXvD4NoOha63HKjbpS47HVCWKEsImJdE
BBNJsrxD8MlGXPCUPMuDlnQn2+W8Ysy9yVyAGi1QHKGWf3IoX/zmveVQbxo/tQWd
7rPY0/3xnAXtepAOSRuTDpwDUrimjvzfJJxjhNAo9egTDsoOu/XIFpiBbAz+C7IS
VLZUdNNS8+s+sKj03wNMzeKgxvzqmFfE/N7kybDgbbKxiYVe3ZP/oeS5wpHnkVSB
c2Mo2JF8GbarzUgajUre9JJ6jkvAR0kacF8j+DlwrWMzcPjsgNXgaE+FMHGf/uN2
/pUHe1Mjd4HEOBxRrGAsNyKJgoUCXpVkrjGCSu2cgHuRUELHOAamCqla5L0A29CP
reVlyHUCq8PM8BHDOYHQymG+LBuR7AZnKKad3E3EzOm1BTfDtXfcfptu0YiUGi9b
VNrmPvqIzJq1FoOzWRkkVbbKONC2Ri6hqluJuNrWtFro/kQBd1m37S8RobAqEmXw
txLVhzKtW1bLNNk+Q5OP8Urb9NJj89gQ3JxrbZS9DFGpBROu90y7h9lfst/q9dBu
PT5dPCymsql4MAUM4cP67i/YVKU3wW02Ji63y78okwX8lA2lfriRfHqN7ulZXQqE
jf0zpnTFksahEh9W2jB0guqlBZVPUFA13ypwSxtioOzFJdpNXuk1MLbtnHI4K9r3
e5NeU2ZZODXPnVp75ITpWgcQRUhJ0KKlybrt+TFsFMEbHDl3QDo9POCEbp1Wr6RE
2tcRZe9PVANVtuzIoId/yJ4C1yEBBpx5i3YR5L/kSzaCTYWBh7YoWDNELO2bNewM
Enn9Sn984lRHb0UZJ81ohex0agpTujFTeJK+iSjLYTubFSUL7BUtV3/HlYu8t85L
A3KVMAA5EUKDNRtzS3PBvhjM1lzi239R/rDLyYdysUKSEUBBsxBYNPxzI0scO4Id
8IS3UUXxGFyS2WGPzPnmXBnaH5keEwIM/hbGhcF9/0j+hLhscfJ6WZKl7dcem75H
f8aOQX2UrY8iWs833qer5aAmqxhvdSFGHf0vxPINP9UQdwBnStBAYKRZh/kIvBEl
q92UsG07B4Jg2VyPF+R2LLbFaec23ZtNHRR967e8YfZQv4ZeWnq/tVuOYPieLrNg
H0SF7pOkuQ3QZif6doRBofFzGJ9FrkGCqeB1njCTiH8zLsFqsNVLzuP+RdzPOwET
oEBqSAQQY3gMF7NuVu4eIaiLfz1pKcExJW2DH/zkOC+N3kL+hDIvXs70tAVVYX18
yna9A8/3asUDof8H7X16WdIIkO6zu4kPp5JtZ1M4wsIY0cPgGdVkd1fgppsrYeVc
vRHR+Ix8uG5QSlsDI7oFVza+j+R6YAnAbnqb9A7h19AioazsnrDAPrh5g9fy0IHo
I0pLSnDWx4n7CzHJeA9SGIJqoUJFvNJZNtv3/27zmeeamKuS6/Pi3Kx35b4QyCMH
yBLCtnY90vMCNDEpOjb4Jq9aSWjJ+FBiHp5PBbAmwdNJrlwEVJCN/4HPAlNQ6//U
RC5/z7qINsj7zJz0W5ZuSJ9C9c70zRg8Yi8Qcry1yYbsv8SZ57zqZPAVropD1m2Y
Zl6/LcY5QpRXMA8jZfoxNgkpIUgoegIEZ6YoEipTtNAVJWkLVsuvGSpW5D8Dmvkg
`protect END_PROTECTED
