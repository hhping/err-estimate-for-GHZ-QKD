`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k1AmQOUPcEuiBiXCXCJJQaQsyDpeEq9UtcR3OUJQCm2Bno6DdzTIPJZ4fRutVhLD
8eejcmeYZOuAkP6iv1TDQfqToLQJR7Eei0xuS0lacTELssN2pvzRWt1BOcTY3dkt
A8p2Au+ENBVYGpmdwdKaVghTFuBPtERjeSDk1OdXlV6nZ9oxFbFoIlQv/zuq/vLV
oNmx+RJWotVjpYcn2XrfVsSGFqFa9YVUH05qsl4wrGWLDms/XSsGRReiX1UcazM+
Tshr+kSa8sMfCsU4URMRCOq9rbMqffkwNA/E7fmcmPcahsMJDbX8AvovGtzEBG2H
LGKmJgu7GFc07+9pMs0Wvh81j5JlpDrcCEwlwLQHbUvjxowGl0OOYomBVW8Rw00A
iWOWy7n1IHtcwn309d1/p04v7VH852IqCfaGCCkHdG/sGKVpb1gjuilny1DUTHHl
y//I8ov4HXuQkp/JTOCDHLxKAGtBkiuwS/Ib16ChMxo1sQf0SaP41lk5sezMxpAW
`protect END_PROTECTED
