`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qy01Yvi5nWRU15RjDFnBfo8yrML7if8Zi+VrMhT3UwsRqGRpmIyQlXrRUeEcg1s6
y10pRif7fssX/L0C8eQ07PuiE+Cn8+5179tnwqIUcemtqHYz027XxAcZ/wxljkBE
4yX7vKqun4097vS3wfte5QLaSgKyInvYtXfNY3S57ab0IMnFqDGyiAMVk5UxKsXU
B/3L8ykNP5rOMDdWJDdXv4WqLVMrCefrx7ZZYNWz8DDbKmALMVpZzqyY431l0J0q
2Y6VC3U+6Qx4l3yt1TsTQYKddMS5jctpY0GvUC6fNX5TKVWYadGVlyjO0ezL2f/F
fKPJwH9ivj/dezm3GA8bYLMfxB+seGTOEu102NAdIULyTKIjxZwD8Q+mHUMTT8Bh
c9b9PE1mKY9kbk1XYVw98HdqA6oKgVeO3dZaQtxy6C9okBpDBygUiIyT3SOxl9Du
VDjqhBoT11NVgRCZkIS9zz3006KXV8DjhpL9Rn3MjfT4TAoPtNFqi1cVDnh93myI
Oa43TQUtvrTITKs+yb3h3DRyk7J2pb/9D0LSxBKXw9hUAUkbbx0qdymi33STBH1E
TytT4Ugj4sHHFZ1BaIjfWCUNsOcxMNj4hWKLMSRDDzHDm3DA22pdvC4wsb0g/qlS
j4J/+qJd7/yRODCxwdLx8ThNwARNt5yNIZkIjkIAqRCoyWN3KA8PjG302KpkfHuX
zHwz1VRoLtp2hnUe/1YR/zbqtRlH9uLH7rX+O2vI2jTUnYf63KxEEApO769gcLYf
+TIUgbHayqQB2XBvFb8UbAShXSaIYRwmkPnRF21kQltJt5YCBAtB1sfU4QuZMylK
8VsH03zCLUR9GFJPsPNkBOtVT+djy8u8kKj6fzOV0OuqTB/CejqdgCiUZVc9wn3N
qcKEGIvpjBSTmOyrxhKWS3iDiQBH8/gdBe0XUb48Txj4B28bZoSi2YoRjjzB7h1k
PqhEq5PKv/NRHetPgDEWqIfly0axk2TUnKigiazJP0ddCO+HBD3XsDjYOweYi7Z4
rxWOfm7z0UkNxoPzqTmxoABB/fm8plwEKDFCnoeKdjJOMLSy3ArTNXPMsacDH4Iz
sM8KT7ITv2HKFCZOqXXbnw0OCmH1Oke/kVr01Jk34NhFYcwUCIXx+dbYnyi/cvEi
FhQGFxDsnyHdsIif45TDrQ==
`protect END_PROTECTED
