`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kUaz8FAMjiK6kti3OGaEHQPbHx308rXbVlbiStjTVqSescJq71UlfuvmM+HJ2/VN
15WOmdXvk0nPUWPIto1XpUnfPKhcCHcWBf+UMRh1tK3eKqQl1UU8IOThUYn81nFK
i/zkP+HRhXXWDLMsMvM70X0KRuxQfst1RcYqLf2vuZIPf/1GaojzxZ9IwuYloRXv
bBOl/lW/qFY0AStULV2K07fPjguUM7vVFDYoyTzuDUDUZ5GSO8JS42lmxyzShxAl
oyfsTJryzcdEC6vlRT2BXUBl+sWiRavuGPHqg9DsrFuj3yAkAkIbbMruo/pcu1Nl
UZ3gor79f1Kzg9cSB8AkAN/GvtIIJpCwSMf1GrhcQ1Cmz/AssCknsofBGIN8L07Y
6hAcUDJkijTSPCvM143QrIEzhN0ljfQaV4vw/RcMle17jhlOIgNb4oacxylvzsnY
TKVJnAdm4pa5k/Y2/Cqm5Hqj2FK8h8MbLQ6cbzGGArVv54rlEbPTkd57hJ0Auo1L
VoVQzvp53B0E7cwR8uO7jtQBVydJSXe3pd/ZCWMICjrA6TUNdUwYEXYO7nRXRWbx
QMWczj6en+joH2c0GoVE+/56y5cQ7wTLwQ1ws1nClmgmYKmE5q5x+vuEvFaFUW2n
CJSaDZ65DkZQ+rg2Q7Uf7hXINNnmz3MVIus/nonwEiwZiF0Td2lUumQ7Kx1jqj/3
oQA26Sb0vLEUy1Bcp7FT3L19eNSJwcAgklTOiGiB2aQzIRfkwStMZwJPRQqq2zcR
60oPe4Tj6vDmf+vlPOIUKmEuZ8fkkPxAdpxXse+bU5J0Yh/BAVW0DecJD08WJABC
JQ8/4Ljqll4DOtXO6cUzUmEBMouw/NQ0nNcts3Xio8Btc/QS+gk0Lycoc+NUH514
qGwvzR+/CK8OoKjTyMsIaQklHJaoQ6YyJ4DzJ4hb8u4ISBOeS8HaNS2cBsDDt8ti
7wBohQ0pH4OJ8crdlmSCTU0nYKZ3MFxIldl2ha75gEo412WzCN+gaY04a4Kjg4XA
vAA4HJstW3nnqwOfGSV7BLm1y2xqQcqeXWZs1xeBIVP7WgfQXPp9P8MYPiSbbc1X
GlkImil5CsTicGGg/oshcyY1tv/A4Rw4moeWqIP6hosT1CECr26+2EubBPKxVMCf
meCV7bVI2YzL6MwZHLjc6IDjc5UGPgYjifnDoVBljc8=
`protect END_PROTECTED
