`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cC/+DhLwJPcEtVNGjWHf0kmQWWx7tw7urY1rgFzHl6qGvG5yFroOZvIYvquh5OGk
A7oDXud6sgmxFaIMwpU34ODO7JASDhZVDXlK8Nb9vPAmmAB9cAU2Lx3Q81nDe6el
IG6OduECnUs93uvGxjrRECbBE1neB2TxzmLt8zDA/6qbK1sJ13KtRr9NP5w5DLBZ
Tgd17NBcDTAhl6xNfuXcTOXcj3sPN0mxHSPp+wgKv/1YNj5rJRfnQ92ifLn642Hu
p9thgyTQv7BzJ6Fzm7TOZNaoBRREUZI18riQI43wyz26xc5BDTQ6MXzEqot4Rz9Y
N9OvOJC5hyMNjOijl3JuU0UwWs0WgUvfQDqAs+T7iBhB3pou7twha24YIF8u2D8f
z0n+VrKJvJhJuaD5cUXiPkWGbFd/4lRLj8ekduTzGaExzcXc9QThkZggfJcPrH/Z
Ji2HjMS8vawz4OtN6uWh+g==
`protect END_PROTECTED
