`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3lUxdC7IUjD2eDuhg2TM5cFI9FVvQVLfaegvlQrMlHwWNWhgfnUs3v7o67rtEZS
RRqrHwUhtaKVzDtHMbWEnWwFyVLP18OTIkExHr5OJ9EreHX8fSer2ERND9xFYewM
fx+YspApdyDw4DQp6JvgjdJRHP0nAvkzE5InU/NWnwo7ZatJjSr501ZVwXaIs2aP
R9uhtBlOsJzOvXkBf2Kj7YSCY7u18ND4Fa4B48LfGR3i5LJry8SZ26b1giHx7vrx
EfdP6OdjdoPzrN6UkCailBaX/8CRo5Ot0uBKbLhMl6kRLqvhocKqz566SKxlKiwh
6nwobMvMqI7Ol+bOXNYDcAn4gLCEhj0wZuI8AtN3Qa8XKkFrK7U02N1lby5J4d9f
LV5AJ7gEeDFEeCW47uRN8pQ2dwz46OvAn2D5UcvxfFxqwUXXm4/wkNIlqqBu6Gby
axz3H24lNZGstf701mZ1XBgbhGrKqRLYtxPGeq/CeACkeHJr3lAllXj41qofUzdt
HSjjrydxdToBwRUCz5ItF/vqVxGVgSZ+dQ728etcwptX1d1A+0ehxR3lN4vH2Duk
qBVAXxv9GN6H91TTBU9P5h52OXLKisoE6+sO8kL7KZRHzNug0N8Gbj55glRdyfgy
DSLU2N90gIOy9ZzxYEkI6AiIU32q8clEBeS/cnBOQe0WJaLDA5zyaUalzqr8aFd9
5gCI4t+okOO2MgMvOHIgQQeMETWIHUS3BG6HTeUASynnFFfvU3g869O1e/Dkbxp/
992uF0fO7YGMjORwDqXkeN69WN0sowDVmmpvh1S6l8oK0pMUsFyL2L4z84uxQl6g
6vPa1N9DA9bbIgqou4C/biWFDz/tTLRNISb1KV4cFl7mO8ayvmvlDMv7OujN/BFU
B1AJbGkzzzAlRuNKrJSXmOKCss0WtKXDlgyS1lX1EE7fq1F26Hpcp6+G3ZT4+aXX
ONV1gHRqN7vH9Ybj13rTmyXHCFEca9kUhqor3UL70CyIUHgBia1Y/doak4wpzUo7
B7u2fkzqaTAAPbloum6rrPTFfog9Izw62meuYSaWHvKNm/+aTE+yeMxugH7iPmAz
pvh1ifPp+4vEd7wxgdp78FVJ1kZCOz1qbd+uKQDY3RRA4EDuEuacNDNvh+EaPy0p
6uFdhqXWh4XHH8fuhuersU1NBDzdZVENgLlWureN0h8FWdwpFv4Ov0UCZD9iQ6OF
H1vZKITGto8G/pBrrAJx2sQrS3HGpPtPPSc0Ju9hLicIsaTjHSHRlbDOPrVDC9c6
LvShGDrTxNjiY+HbmygCiF0z0BgZsNq57xd5dk6twkJFxwSyh/RDHVzWng4vCyj0
w/59YyF0jT0Y49vpi+NvWbY+DdAjiLGoSm5W+THJMoQhKc6FTCMVCw2rK6/At3RE
SDGp8pGRuGpoF23L5oVwqv2viCvm4gZrv3r1paZadhKH2kIzCUCFt6rTYBaaa6Ze
ECjwQO3Rng6fpuu3wKQLVe5Q/H2Mhz+2rATwllPFDENFPIurB45dkM4IjHTWVfzm
Sb6MXmFwWxYy/m+Idb2QL4YSJwaLfpd7XIkt1O9vZwHVqKhJ17UOAofDux+TnU4k
QDUjc0jFk0WBJ5mNvo8emkZ+eJ1V6ate6S6jG2vvTz3CXCc+bdF6WbkLtg2ScmS+
i/p1TxfnFhncQeIsr59kHvG1oN6PWWXPDwfRUZ99ClU8eZEzs2CjCSxCBAgRtI27
i403ka4joMG2t7MoaT2eiW5IXCwE6CZReg1oFFx7Gfb2Zlo8Ab3XjKRPbruPSOYy
`protect END_PROTECTED
