`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eoMsUfZ1aw89VpDMczC2uODzlr4uFJ5yXVXHo08UW15Tnmu/EyuNo1wN7NbHP675
khJX85yAaJIAgXBCsixxES2VKyZK1xXr12GLXN1DfhQGAsGliDXp4ojUpdS77xJV
PzdiIf1qw24WD1vaVky39SccSNIvjNO+u6XgT7faouWm2kwSCmGwfYWhjM5WgQTp
E4MmMDL+jMbmwtxlQNtdrjmc5QK3ZGEfFqxiFN2trI6I1H5EUu8egm4MX9UdYonn
xunfKBN+wS5wRtcIuPh1MoFb7WEiethzrQrGnYR3zZRKwcVuqIcCaAPswE3MDwuU
snNheCPRfZ3tjn0As6w1RAX+4d0AG95CSqjlP6SyOW6f4ubeB6rwSsLiDx50LQT3
rY3XkIjN/meHz9JcafjHTeoDWdpl90DAtxZ9Ty6GZB+o11hcISkia2sz/BbDVLCj
MBh4FRLCpza86rbb9vEhjma/E5uO7wTKXgRVUP4ajpfD4yHcabBMPy56eAv1SSjx
ZV2j7qXoawsa1m3OLIacoKYivDA2/nMtLnSQFwGAHgmr5I1zbLSLG1MPABxkwLcm
wlpITrVDSpINSJ9kfrH+JZamhonz0yint2yaK53hos+EPVY4jlF7v1qCf9lCQ/g1
GXKLsHtvATSBaWqXnxqjBhQhDFZz/JhWbThbp4T3bmBgEXC3jP97AkSAr/hQWLJV
7TNMNlfmAFjUW8rXV+NSgrA59V9L0rM1HQynIIxL3woG4BH8S3NDVDMqxzu4d2bA
RU3cdi+Q6auS3/Y7af4UcEdgg06u88JlqkE4ReXfJPzC1VL4Jgvf6KH4Mb5G1ajL
LYG+mEu60qHgVc1ozZkZbt6Dd7u/A5O1M0/4gAWZeWkLZV4eMAsJRp3MNCOoXNru
l5lVzhsDnp+yPvw9soaL4uPFgOHmI0M9rquvOsivLe2gzUouhlDrRyp7E7gp2wzO
TMg5i2HIn96IU9N6IQFo8vo66i8+NOqCFWV7/SxN+FXtHnqBefplOgovWQ+cgVAU
hANpKtsZtOHlxV8+mAZTOBqZr3Gp0hEOCqmGXg/IeLqh6KH5EMifPUsv7tO1oEIn
8ZP/bUiQeKOflVhLUkkd8WCQB4VaHZv8SfOMFm1buf7nd3JTtsEYB/KWIEch6uN7
KruZzyfSWRb1nRPAwZqMM/IAJo3zjHM2MsnwCPQcUSsOd7JIMrBblH5BQ3465kh5
`protect END_PROTECTED
