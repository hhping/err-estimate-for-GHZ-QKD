`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fy6gf7D73SimJFmjaYbuuDcUyisRkqGNL7HiPssTtZFgtLSYDOaWFQ1iggjIKIC
WbfUmFVI4qevVZDGoYT10tMejIcysi7XjjgrV30bjHuG14Knp4Pe9niMiGXKyn/v
TiHd3xZ+rdJWRO0cp0k981oOHrQl5SX7SROK1S7KxVZ8zSqpBbDfrKQJLd72/mo2
PrrvkXbACh4vG2KhEDAmcMaypYGiM/VaX9Ye2PM/L3o6HwLtTjXmvmBOs3knxCUh
lB6Scfv4eMz2CbW9uUEt0ZlC7GTdv5salB8XtnY+1fmsy0Y9HqdaNibsd91T/CG5
wv7PLme55MUJKKepvDlRSuhmTRNHKcIk36G7Gkvk6HrISlA7AlFzyn0xJLWd+gLY
cbGML+TV4KIeAzbPXtdLpRiPI3BtqjDUgpVH4ZvxuHlAN9J2VDTXeA4ZJBHoPzMT
qU1poy9ieXtLIcr4C06h64ktp78Z+hHel8bffBP+h8lWQkCwYuF8NEjCO6ZBlBn8
m00L2gKty0L8m1FxrHnzI5e9ZjQFav/pPf13dVP19hjxlFkfa0FwpXz8GCWyLm5D
gtaYEDHvaqMTtyMWYchss2BDT6LQfLar6TQ9U9pyo3SyXeR5FPWnWw2pjjrjrRUu
wMy5WpdCmao554BXgTlGc8YhRZAReExci9iEuMF9oHEpvMexbw96IRUcnTsNV78z
XDvMO7dNdAzQep4Pe1VOnE1SJ9mZ7DAEKhnjkahZWMxWMLpNG4S9qcCdPZWFvLSR
HMjfXaOinAzr9LHSCIWy71LxAgwo88BpRxwcW3vnkm2ADfFqnCHrUM2YkPXbP/xH
j8x0B1dko0KmZaKz1wBN6oM7/Lxxrq3T12gOI22yDncR1AHkHoY7B710Gc6csT6m
IHdJpexYrRZ6skmmqZj7cB5Ca0vtJyR3XwsH8A32Zao1TEzyYnMLY1nX2KAvz92n
t33C+6vUZd9N+A3j+zji0zbsuNhNwYaHmOX10XfylwNj/lb8AbymQUr1KLPNxmhw
DZRCNuaKCGtJMoJQCihrrjK+LURxwqLfOQRdEhabKnmWH0EBGiW4lAwK6lglOkwP
dWq66Pil+0CBTv4EbsewCIZVVv3lh3WXBAzOvQONOtSUpxBc9tbtBPknOcvHZ0wi
hA00dSCNsXzlqvQroVXSI/aOqvbl7gb0NPrJxmkRGA8IWPCI62kgDpYvWzxAwllb
P6A/enJXDZAQnYeBhLcomfP09y1jenfhP4L3GjWtb/kSMlT30mhAEXJwcQ3WGCFw
Dbrq0OhPGZeL7oJQBwQrEioGJqlB7KJxMGqEkYQP9EvrBWu81TCYCyfVJ6633fr/
S6n70b18j3u04NIQ8PgBY2viZCs2CQLOQ6CiosXBU+BF4Lw3b4Kvks2f0SKEFnVK
Z8BSh9r7vlGSI5eYuHG5UVBMH4ooS9FfRWiMcW7v8+oLQMoHAJv329L97Z4bKkJh
1Aa6fekdJB4/t/oRvrnMvrwFSzwsdJjYDdiunTp/jHEq7jcPeHlL1DAfrqHQWHRQ
AC7e1CeRqRG8CYdk0PqiA3Vz2s9AoxJ3NmfvJGUPbZ0=
`protect END_PROTECTED
