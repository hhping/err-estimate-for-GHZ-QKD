`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9vwY1vYSrYBpsrWrl43d5jjzU/pC1eyFxAVg3Hp5K4ihEODQqIjEkAqPRV2lb1i
uvm+RPREn6jve8TSLUg36Qhl3F/N3afHDLXJKaoL6mj1+ogo6eZxqFj9tA/f0bLR
EehsbrRYY5FDYlc/Z8GWUmmpFV6419yzMfHRGfNZiDvKSs40Aw7sPhPzq+ZwUKKo
6VPI1w2ucd0NQ3/euXNmvMLloqBxEs+c5xvJ0joxFG4=
`protect END_PROTECTED
