`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MfBM3Ook3ct//23/UmlPEgbrFsXkbPQ5WjGSrvbTl9aClAqVEixgl8JPuJe2XGNT
f/+qhX7Ooxi+9OTN/0vu+GYz+BTX3wkxl5i8Vq2tHN47f+ZApjZ1YGnsn0AmRSed
hfXpiuYvQYvh+5xSjqoYnq9D152ruT+sgL75Zu9e1vGbnYoYvCfqOBXPl91eXGnF
IQ1jlp3u3NUXlMf9il1jL25SvoarqHRqoNLzMAJ1LPO4rRvaGIXML7TG3aApqhv6
OgwhsifZj9eUj7Fp+Iw5rNznaySlyULD/78O3mEceTgk0X1tneXoyLlvKzCYE+l9
yOW0FiZkjoLKqll5C0lRatQU2bv3bvcq/au+yvxaKw+EahkuFSR6pdAoAObOilnb
cSODwKVhM+ovHca9QPmblydr1k+ZKd6AjxQdhhZ78TvjBZAmWqMLDXlcAigyplcX
l1UMIyiSlfklrZUc2LbSmd9i8zpCicJbhDDzAtWA9CKZubVoZZ3Cq6WnVv3eVtwA
Q99v/vOp14/mRbOPLBkIQl375Xo+FSwAjc2d6sMLWRgt1fXStp42p0YSkGvbFUoy
oszR5Rj1qWY/LkCshyr1qHIUiSL2plFn5/cxy6qczcjVc4Xl+Xj3iO2J22X4CaNe
cHhYvuqtepTWjugyluL3AQ==
`protect END_PROTECTED
