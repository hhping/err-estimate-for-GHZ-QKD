`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQIPpxdf13vgN412vRMSC1Pjk78wtS5c4GWjG0cdm5l91lZFBbHUUBS73wHAONXt
hrgw3tWUeJ2lbFQnt2u+/5tNlMidewmnGv8EXgTl6+MCqTDxCfuggb43JLpTfY4E
kb0QE4jvS+ighO2qEXaOogNAKOVlEv7EdysbBZm0Q8Ni1FPnZID1vlt/aA8PwX/+
rAybp/b6C84ZOkGYVrcI/642ntqP2dKwo89PW+Ntj0EQQBgPqyQpQf7QOszelcS8
b0GaEgNHN0FSuaDI8+IGbWw1weJykBUDZ7fX9Y/l0SuK702tUJ1RFcE8y9VhvbTR
DwwF/Y+d/SiNmw8ACXWrhnpmxHUW3BqWNdkkGR46RVlUna8/SVhqM8uEHMiDXo5b
EpRSWG30I1LDh41So2xxHD77Wb/2ZMVBJ4cc4GxfIt5c1nuNf/mHia6G9aPDCoiC
hqD/xn0OlJC/c2QYBJYtbT/Dg2kaS6P2M5eut8FK//2/5hZrwiz+O9p0aYMiOB7t
A9Sm14HOrY9i6SKAnhUI4HK3VFNINbQHiwj6Pvb97HJOMc+SDcgKrT1kbcFnAi9T
41T5c7tyKY3sjortwoDHFZz2zI1CSisaZM+4NRqz1FjzpPgKQhFXsIACQvITnXXq
cYi0ukvQ/mwGwiPiFBzGVXAGujpK/a9JYkTaJKEWP0uzlsltutjtPcc7kpitmXk+
VCszd60WWbV1hhwobSa/LUk6PilKTuF3Giaan2hML4kJgqr8n5Pybi5FWIsM+jnq
ruojto6qvr4eAcZti9FnNqluZ8LQ0Fah70DRs0sOFCI=
`protect END_PROTECTED
