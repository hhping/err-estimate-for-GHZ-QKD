`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DrIf88sgrlGGqRyIGTrwFgKQa3Fqs68yBBs5vQcPszpSUKEDj+VRsv1l5+VSPZRZ
kSr3ZBR/nkOfvA3409KNsvlBg9QaPyyCWSCTkpxsq63wgot+V6afDSz2YFx/1PWM
8OcL/9Wlw8HBqp0mwLM2o+Xs6u10kOGlBXYdaelbKTbNcjMK/G8l2hos59j/8PHR
eIsq4HWJ4puJKdeeCNPLBevxc+xrRPjnkTVu3iXvNEFSSdw114LYpYRUFxDOPTb7
Jdd6nvyb+WAQt+K9ui4wntAPsCjDM3mfZSfb17HDtkz3jQfK5gltCT7gThxImw0H
rkSG+pBTwA/BlsSZvYvSWsMNWIVbpmvhJLL6/C9b3T87rmpZrZhU2HH8gQ48DaZZ
MYkfuGSVUhgEv1I+EGhImI+LApYqdP6FktKiiu716mUeN+mi8kpyBmtfiiFf90X1
gg6nUh8HFJKeqFzCPNHzLgluWaXPKrhOxe0w3UyK6mXBqwLpR74kR92iV+0pXaXv
SoGK46xDmNQvdyAKECQzy+GYKTU2wGn9Bu/GEvpNCZI6piSYgdMl/d6BQw0mtBMW
5GREVs//utcUXieZqLB2QM1T1UR1vfLSGnD2aBgKQYzd1aM9PqyFMYQesbtzsn2q
EX5J82kzfLXvI4mqS00DqI7AsDr00ksoQ+JQxFgwMOj4xBG3C/W0embVAH90qbMZ
W1SLb3uXos6rMQLwzhxd7mo2DJuugRuHEIFQlBcbITuLJmRhtz7u+jUFv5ap+aVR
EOdYLCVhiM+n7HOj4UsHgZp5p3F7H7TzaY1mkNwon7PfygHC3/O8w+DvIsYwOhqF
BLVnGy/unKysi6nHLAF7RJ1Q+4l4BBA58fF3RpqQ+7cI9CFaBcV1XAJ5jRicDRdK
vxWJf7izVYz9mzO2Sta9Axsappi1knz0SMWfca44Iwx8oqGB/ApPaMXiHvMy5zwW
VNCb19OEZPZrgWKXK2tKtGGKKPzrF1l635tdzxkQmQBQewBi1WQQBDHJdr0vYEbn
kHVn7lhdJ3oJpd5lDuQ5lI9i/2Qc4C4ShOONin44QYyGq1Y75qu1xLdiKPZ5uOU1
34kf+NEGEhlFvHRv9peA5+Bou8ieb1Vfa6s2QsOGIcF7K+UwwWgv32waFfz7HktK
cEUvphZlZdsJvPu91M7h4pir9MLxWyJ0vjiGePxBWADZhGet8B6SyeU80owe1a6e
iXCzkxL7LsJbX21xHeiBUn5A7nF8Ijefy3Jco6enmkf1JT0sy+tfoE6lbvy7JGsq
HNZnvSHliBQUclN3hq5iAAmwFgHLw7UKlNf4wDpb3a+lHGa7Po4ReBiEu++ue7UL
SUeGMnBVzLYNsYs/IbYwp5HccYjex4LriTByZgeykmQu7xEr78/S7OuP6xbXeNCZ
JKtcAoNOXdaqVdgih+M7L7LO6ovEUbkHQFcEFCKTOMCa9DHaIFAUn2YWJZW/Vxxl
izMAUiImHRTqX0tBcz1Q2ReDnFAJU2urknvD6xmUFrlbqgQPPOFeIjeZcerUXsTg
4lxhjwEY2Di0qDZiLz6UzufmhPD5a+fbG71SVLjDUzcZ10DxGQ1EdjJ0pDw20KCv
`protect END_PROTECTED
