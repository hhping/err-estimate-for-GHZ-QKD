`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDC8gCiGCO0TTsO9yCk21UhYdoF41nX9HVkw2+VBUWFamPaH7+7/BoaX/4hIxBkl
QUfTskAL46T5Paq9bgTcyD4r7MXIl4HOcHuLbFX/xTYEgOSkpSpkcQVt/Ix8bnSS
7d6UgZSKACsZ0k6EGAYlgW7EVIQcjvpEB19GszVJJ0laghNFWc9DXrncVNM3l/ws
PXA7lXegXMt2MD9fMWplQT10H9G34Hp4Hf8nPfdpSngA/SbuEcV7X6x14rFmLQBd
AveejoPAMExKrGSSOhzdzlQb9qKNKwwzF4qqtzRdXBbTyGs21GVIyxb6cTV+a8bz
EUGTZpwgpCmaKGlan+WLjsDRC3hic9511VFAENmQNh4klzRrvOOa6EpFYmE6RDAo
7nE//pfmEoDvfWVzNfM8zSeWcwqi83ZlOdm7YXyb+1gI3HPHzGn/OfxIezYtQKXK
9RWJJWewND8IoVGYclq/Z0ZekvDz8Or6T7HKuxqysWLFLqlgj3xa33UPoR32JguR
8v2Dvf/Y8XyaYx4Ofyt18jI80Uexw4RkJ8P0ZOrVEA+6he9lSjVlEDCcTZ0RxZpT
n6YM0a/4ZlXFhKS3w6NNsjxm8KPqWKyd7lfbc2AqRDSh4a9MAi8NdpRxNWdWQcs5
BTsy2G0cvLDLKDFleXRe+bOPkjOa10KrrSPDjyG44crvY6356I311o4f601bGecy
Qsrdm7VRAIDwA535WTq82hh5FFL20faoThTaiEQgSOIbw3Mbh1SIfSy/SXAkDIb+
Qe3F5AGtB9GSPbZULlHGlJa3KjzZ7f62IT0fzs6JZoU072xL4/4xQgBvfhe9EfBA
48ALVAxMC8TKFg3SgdJ6wA0kffxkVlWIT+fbxJsQ2SyBgY7Q9b9yGTESrTQeARfM
D5iioW4zZC/eElx51kwmS9aOitePmul/2FPEpvCKfb6uBih3tnJzGgRbVYCNxcMz
iid1/beIoGb0f+Reyb+wR2FlGJUgvGLR7IKu4eXoKMrXNtkQYBfd9W1zca3E1Aii
qaoiJevruxhjvh8b5aX0k+ms5Awq/yKvIGzbk5xXadsoZiDe4NnkbRag6xgKeJ3x
CQSaFF5U27m/xVrI2bd/p52IIX6K6tkohG3MHCy+x9ohIZ4lmmpKTlIn9hDr4ayt
5SKcAdDlo5xIaTptf1LA40oZdaomhyN6zY7Q2CjOl2sEkBN+rZxD9f3zhwu3SpCi
rmrYBs+1LzHKp8xiQYQIBiFj3QawhJdUhhEC/xwwWaA+kon0kQbftaZ80NtJTflg
KeznCSUyU17IKojzcjAhJNvApiuoSHA9JN/UwEDWXMIJwTegpsVzuWc8gahjdEce
QS8ZbYrNfCMsvRzykbldDxKt409/bxEh+ZYXGtBFc38yVMh0znVKlhdmWv56acE2
S5Pkhvo5c1FZnUdqdcrf1VYUF22D1J5C3AOxeOxHVgQczHSceR+dj+w8ObNS0330
N46KEQPQNqTB8Un39FjoOtf+/rcSnFwLXJ71i0ZKvmzAMksPPzlt15KG+WInvygQ
yeMLnUiG876W/8chkRZqXEKQaumWee7KNGchJ1+7+4gik+RiwJ3lrJ7+jELhJX1S
kCxWSCx9TpW5Lw1eYbhNoJpxK/mnuZkqyPRlrRyLlxORINvtAzCJea+jg+rNMlim
B1xM8eTkE9OXQimO0xKcQu0N2MD3z9dDP+sVxIMUoGhU6S60uBq+2Bp5q7RlBqd9
tH8DgBbG6o98vwtGIHiMAlAHp74Vaj4qSzM30NaxoykOPozq0u6Rlu6Ipj3KF0Eg
vG0UySV+OcNNEmkBzmvNTbK4rLVmNuqaZUcRhTy/c87RtwRsaCom3y3ZtF0pNSNV
lxBLbFhpyFazeQFxyJ1S29totNRUeU5sPjWfGXr1wRQIFs0lNS1MfN56lVLWF+UG
tLvoqPVBZosGopqZpE32pwiqYYoTl2SEtAXvMI0ObAgNBD/vkAXu1+0Uxm4ryl8M
/184DdunbFCUvxgbFVuqx4ajK7H5ibiSHXZXxyZyFR5JLay3C7/8Rl8GYrZ9LOFP
qequhssZS4morUQhrKnJS3tevNibXTX8DXRTR3yGfS96GKN/SpBGQLb81CMz68qB
r0Tz9RM9OYathcOoj3EOF6+HXTF0kQ5CBpBntWsTIB80pPsmI+1na+KWzQ86sp8a
JFu0+t/ewujkTZuz1gTBPrduGpVDUhgBXqdIOoi7G4QX4aMkIHY9udMo+WUEG+i4
d9JxGJRG85pHOq+bl3wgjz2OK9gpCt1saKGRQjWF+51qLjzHYk/o/6IJ2kRxS3z5
lNS6DzPria/BwLrdNka0PEZSV5IzNHt3jgoDJQ/bjCf+yklCs9C9OEuNGpV54uy7
jrO737wF/N8TC2nkjyUR6ZEEy0FxKcCaOY3jbCYR+UXzQVJjO88yiYi4skpYOFBJ
nqxRCxvgmmrik2bVkjYJ9AWcHLMBm/cDT305jbtmK8/zxaxkWytJv3QYf0E7j53O
CV6EkIoAWPCQ9MtZuCxv6oOt2RnNtZPaKaUdnZe18Do6MsRI0G9yNNJWj3SQat92
vOvqR5YBr0vk3uk+6/CM3Fkw/6REobbHLrPRcBxRaRB2Lgq24hJUQybivMYpRpqC
Dydo0DTXwwjIPjkMUKlyvtDTonZTIu9LBQT4jjKndupMCrRi8Swt+UFGqugbHEXh
j6VUY9WcxXW5Vy9SgndDKxUQ5PVmD/D0EsY4AAJZqoiyMlyZzSoW/EwuSYCiSKve
iY11dd2APNS/ZR35PVTtk2fDjrtuql9U/eMBNxCecsHM2cyeV64TkyPfCO9FyV0T
0MBhJ6HX4DsXUqy/Z5mq74sCsrG55r+ZY5Ilmv1mt8gq2YTyU0draAEhiI0eyPNz
9bNHrtPznuUXEgzOyBdDg4Z85yfx6Y+BTmg6f4067fc8aPZWd9D/ANo1+LQ0JPGx
y18buSFgkRwQ6AsCYCwNFrIuhcZcCkwcERbuDeT4ZGmJtlDjLKvZi8R7AtRMSM3Z
qwCPodJLWmgr4hslQr1phFtxNrnAsZkG1Bx9ckvbt0314y8qUpO69FZpoqpjFx/j
suk8U2VDkt2Klt2kAcHONXHMOFnSn655XtOTx7BQRs/nKj8/fEidKAQkGypNELA9
FcgMxaOasoUu1Tz8nU2KshY4WIgfoJTrrMaYYfFQK9ihqrTS56OQiD5VftA369QW
`protect END_PROTECTED
