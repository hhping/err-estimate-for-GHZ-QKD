`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LZx9t0ueBBLLvWQ29T4tg2yhJaJl3cCKow4rVQZvXT0e/rxB48sseyMgDIYeQ50
I3RQSD3HibTk7S8sDaB/W3ZBAXmYbk1sCQ6PML0usicfX91F/+u4rEE4RHh7ud6P
PX+zQVAfJhroM+F0nmNA16L/sWx/Zr2Sk5MRQJ4rcxbfUZKt6ECjpIB0+bOv0yUe
4TJ2N9xyY5n6BrOtzuwxZ/xqKPvyp+tWvwHUARQpb9Ni/0NfKXAwBM1Xd9/4GB+K
iYVaxbOOO9Sfg33ZZ+C+JiP6sbux6TwHsv7rcZjVe5FbBCjhbhz4KEPg+B8ZaSnR
DDTUwWJTY5vxtom6HtArK08D7EXlOXvtQOtQP9YoXJXPPEuyMEHUX6t90ONiwh2e
IxcGQctllKvH83DyLsyazlk/zLG3Gv4uzIOlJizxJPYSnRpUjKERxyVmrQjExr0a
l3mqSCHrJ0iHN7NVjp9ih2c2hsKQSaw4FPnEIQK5ZT9J197R0ONyl1q3wO0DaS8Q
tBk6viwDt3NIcqQ/FihsS71nh/tQ24HC+UnB9YH1MgXjO543WrLRKYNFPP5dfJDR
2FYTybI98Yx1GA5Obh5T3ETR0r3wrCCh5p2R2ycr5U35UDQeBnOR+/B06LTK/Xbp
DjgCD40vC82koQi9p37g0lZLxFxX0I4wzfmrTFzGgNabipaVtGJCpBsyR2kncLbA
4ArOEzJK9o+1rh7ki7c1ejgJ9oyPj8Q5VKXlABuLR4RBUMQEWX/wK5sLR92Df4ze
J4U/SsCSpjXOcu20+NapPKbdLAbmN6jmi31zR7nxgfsK5z5krhaPTe4NuYDRSKQ2
dLqUkesydOEhQQpee3fVibudxMJfgMVDE/RBXjgVoOKiWgHMqdYpYtege+HmoQYq
O8wLCwslFwUTFxc2jKbNEE8Zpcw+xMCn3/W9CkMe9bel/SGoL39hpbysHxuMlaPY
bZy2bP3rZG4C97dZkG/z/JfhkGH0Gn2ENTtm7j9cV1XAgsJ9kWz+p4iPPwsxVHdq
uxGRrAHTNQO1sui36/za2jDVKeKKituY3ugmUnPneRBIIB1dxg90ijBdOvyY0Chv
AtpJeaTvf+TAwZPGGGPCS7R1liFy8O2LyrnaZQj3h4QRMckimN7nVP6HSXFEZRIR
eJqcLYndW0OzN3sk2s7OYohsiDtSJIxFiqF96tE7Jywawi4UWD+n6qMYFiai1tfe
OeCkPRS+T1ZBlqtgdQiWF+5Xr5FWX0L6ItCFXrx7ll1y70+Srk4knsMByMMWY3Lu
1K48By8ZC9v2rMGqF2HfuFLLkkMSk+1ZhXve6WexV3AHgJw0uW+bpxJ0ewV/nPZ0
bt/XELxa9Ut87pY7npbntMpm2UEoY623WEEZk8rGbuq3/dpk/yGQOt6LpKrJUOxk
LuziFADl71rYGht4zWiQYIGv4z2aM/YACpShnWWSoQmImXUIo4ie9RtnWx4M3so4
WxmhlAYaAEo/JSDBnuBmo79DNechfhyGABExd+HGW6AMFR/XFzSvcoP7hiHsKcgg
YWBrPNnx9xMzMzrENzcADa2v9S7PLeh2kYN7uIOkdFlfmjDy69MNJiqhqpozZZQF
mXKhAjBtmlmIn8GA8HTSfLGQ8Ef7dPbC9fEzOWdYRky6ICWbtks4y8q0OcYs8XoT
+XtwHwW4AKCcjGvkp4v801YrLjXzdficpKHjg8SncmiArUIKbgXSKrzm1K/a8RnV
OfvpgW92QB7ejUuHp9/JvGC11NC2hspMJIGW4qq5fGJLgoxN0gjbhVBwWlwf9o6F
9gjcGiBUitFmfEBUs+CcvBR1se5aISJP5uP/IYJ4vm8vxmb64rbfAlUb1XWD0YMm
28PfGY4QMU2XiVWWdR4NOCvKCfnYPQuc9KoToAjaGbKxzjEhX6LC3O05k/PgduvT
X2jVi9zr9JkqczlxMr77R0OLaXCdlImsUoBrB2zHWUIDOSjq+t0yiX+a21p2J7eJ
lCQ1+wu5kdD86w3iTlfqtfOg66D0PPos79dNK32NBt7AXSm9WeYpuEoEGnNDfq0N
clymRYZ8EjLhEbUUge+HLH8bzHHwW3frysrRr0H3yJHgMdWObFLR5iq0EQYS3tBX
XsJnJrTHe3dyKpIQQlZlJulBYlYrKLOv7N/BFdifex34YOrDfEx2QtKx+QgE1qiP
9FPtAj5ZtHnd6vrzVNi8pTOh+2NtsbO6yr/BPnymWjMABBAaOkk0pW5b0XuCIQPF
b4zPpxxGmOm6NxkDV6X0AHjmRsEYyVKAPdpTQT1P9IeayAcu2tp6vDprRKb76VMi
nWT+Elv/4somSnr6hrr7obSHwkYBvXJXubhqrGGguBFPM86hthZOebLqg5RxfAtP
1zYyel5RHjHUwqkSv6HFZUB1k2RkXtL3PIGJMJ8UsalmZchfFuo/WSW9bkjyWJUB
fB1MJgZGQvZoMeKp0nA6uIb0N/aen6tMhXN/tc6Iv7VwAszvC6lOyxDKfBlql2Wu
oglP27+pAoLPS6vTQ2mW/0ML3MVpgfO3EWzseYa6iM2AMx5dgAeCvKtTgq4CHC1v
YGZCqpDSfZQjGVvv9PbpGGcI7nqt/E/AFL7/9CBUPwig1c6U1/JzhD98yA+q2oj/
AbH47Xmr1VeteJpig4Mg4IL2s1vLf1VR/euyGJU68rfq+7K/GvpiDzrXXXISSlXW
CM5AjCXywetWEix9uHPv814Qtoak3VCbUsxxPrdhVvoQAXyD0bEDrzV1A6swTb0x
RU8fHuXrKQSq1/1ONWe00phXD0Sx5Ka/NZyuMIuQRETW0ldOzDcMK7KTRsfjUTFB
5FnPiIQUCXsXLQlq+E3UWkXm7UCRrtg34rYAztBqLoRQXLJT32ixa6wQEUwokC0t
RdRn3GIlH7Dk9oD5/I+lUZDmu1fsYiohc6rq4wJAZezTreiYkRCgdDEv3qrYmOLQ
VgD7lNjjlbqS9Sl/mbvPUOnqYkeOao+ZqknragoyzhgFRVlN4AAurLRo9lvpKotZ
vJK7ZHGHkwfpqZ2wscIY1gOWq1z31dUgsmaTcAlk6ej9nvcOHdngQnbbnNu7dc2i
4qcowg8xdY92uudY+WGNn158HDNyqHv+aHt/mwRQDDBcmrP2HbLo0guVrKeQAtAi
jv3htFTgN2Lm9g5r5uZO8U8GEGwy7GoG8jCG9a5ObL2TqhSCW3F1hnacMW3NlmFw
edQ2CxoB1Nfzvag+yh4HLLIa/hFNm3I5jz0Xa3WYAa74wiUg1tCjTKybjFchg1da
t2wrGQAcBgTJ4JBv0hmX2o9+nX16saqQHEMdXH4cNDoROwexgUGiYLL14muY4VX/
rW+kJkfmPUoTNTFQ/t4tzR6qST00P401hTIsMPD+6Zwp8ybqurlOhRhY9LJFlw50
Cu12AcCvC3jnLUisPZn3XtpI8WUDd66wjzKDH+lO6hVRxqbRBvOXfk4eDnDjj6To
+vCcuMSWOmk8L4sPuPA/UwbdyrYwc6rUkq8ACxS9UKEDMwwgA1KA4Idninu7NQ5W
aAtI3ExpPeVJZl9hfl7B4c3VUCRWU8xZRZ/kv+R4t1Z5zt+skidhydUPtZebi00p
xUhgp98jR1kA2CdbsF8q5bNsTSRnxx/RBE2iiorUaw/7uo3xs9INc/ZQ80bA7aT/
T5LNTIi7kzu9Gj2HM+/fsa5dSP+lsx5UrzmelHs6HkyiD1SlcnnPypeQOURy8nUf
uJEWXUM4BSupF1PbqCd8ls6BRTk8TS+r5T+eY92XAGbwqDJNySIPZ2M3rM+JIS7U
jKKx7wwflrOYYUtTw5bvf1CycoLEk0r+zIOEs6O71BtpeOG4+6CaoqTYpQr657Bc
zSyHDdNGaDeLt3d+0hzC992lFJ9+XC9SFv6N3NGkAeu+QR1o8nYAMT/EvoYlX/mM
B6tBtZcr1yUJVECU6ErHcozjohi/3UCUI9tgce056CwWuC8/4XrvuZMD+0sYCh9w
aMkX9C1m1SmW6t4uV8ue4twkQnMWPeJDd78+H5nPdWYeFLP9hwNoULckBwOmA01G
wj7myYO14w6DTJVSugSBIYifXISyAFuHdCSPBs58ZqHteJYNwHQcXrAzXtW782fU
Ep2rMo+DjgP9rGsGRFKqOdT8uI2fW2AtbBooCLUZOroJbIaaU8fUCZ0OMi42iQDz
epLmuE96tUJLQAs30V8WIXwvoy45NO6jL4zsSrYyIQYxVVXxFHPbUgqpEKbp+A7V
3N/WvE8NznBFY/mqGnnuSXzVse4rfz+1yuyo/ElkwGzAvLM+P+4FFbI9BpDsbU/Q
wc14Th70NcTQ3K1dbTCm8vKBBnvleb8deAJP/4eVM3M9SPVoucxzO/7xa8+eP6xF
1gQj4RW3KzG7+KGPjSwcrd69ly0xqWd5BeBr88OHIWb7ICN+l3ohSyvTRGXX/x0l
Tji09iTWmjT13J0rBUIhYh0BxgNaAN0TH++hU00rLojX5P0msw9JRiE5gjIxk0h5
quVN+QAm93XS4w/sdFkn3fJdFbeIysYnuPjCBYB07ut5set6qw2MtLIAdqYmbPHq
Hx+pTzZWfSsu/LtpylCVf0cxGgXH0vNllHzWiFXS6e2PV8yZ5z33ZNBlAqNGPCSC
17pV6D5jXOPLBUnYV1KR6v+KOGFKqYnyb0AZKEh638kcfsQuwsqBWsMZ0Bu0VOSw
0D0IUCeimAYajXApKd6yFbIdoGoKCjRAzIIS/7GjPRoKzFFqQ6O8WEUf7/QWVFE/
g2kyNykRU6mN5ptVw0MDPHGKd5YoFznov4U/KC1FQMqd3MPfYvzDIq4AaOBhoNF9
aV78ASyIl4YJDYjSmp1jQQ0f5Bb4xRvbrxPR6yD8WnEzZt+G8SFKJGLdc/T6cIpE
xug76mjbsxagKoozYHy3vs6FrcgTdcbrpf/2yTp2UZoxm5eY/iBJ0ybhHy/5VVf4
qI57Lr3QqCm4Dwunp2Js6Sx8s1OqY+91zOdZr8LIMsc04FfDW7Xdma3J0wpPnFsg
I8Gv6MFqUy3bRM0UuM/lFf4DR9TDpOVDbZl2DcB/x09BVeqbs0Xz15gv4UXyYyFt
6Ikh1nd9Mtb7CAoijpBgX+Atjou9eTQFPn90kxLwx9aPg3aGlSCwUnC8eSZ+z+uo
FVfQ1JrbwO/RCzujo//zwa7pO4jaqQb/vFj8RA7Knzj+553vaR14ssr15L9UDRiO
vWNwfaorsc9ncOOFBrnCwlf/kUcXJJEFupRnsLaOoNTeb609im02+xdGmYDjxdaG
mAFVYGcXiRpWsHc0FyVyBaW1IS6LRMvF+zrwG1R1Y7vM1Kf/kcXRQ67hmlGAqjPU
VfZwcwEERej7Zpy64eL/FKrMWQg0OVZBXWFqZMkZccklb07U+qu5bTiGkg0W/prV
zlKDnRkL1nQ0NywUDfFUb/eajeV+ylaEx9zcvEvWshc50NhQl55VhJiZXERUoYkf
CnxyPImgSCkZz00ynniU6pP63V11+wVhbIfGoFeB7gfMvmA6w75VfNLHD8uZpi/Z
VhFUxPtNWAGQUexOtb9qYa6i0eME+CQUfEA/W9xKaXKDwad8vnj+B2/kw1Ow7wCZ
L6N87WGrlqKLYM1FihedcER5LGIhfQ54bREGHVnBK/pwMZN9ynRSDqo1Yctd7pQZ
5UZgZ/lePxDJBX8af2YdChaTv66krTTziWvPtv32zYE9lZ8g8V9xxGKMvnRgoyMj
ATfceD8Ji/xtZekQPY3mqSckZLgcUyjUmvAWQbZ+CeneIFt6ZAn0gqYfSpfyMCzs
kBf6l3C1Tgu2ORLG6IYfh8xTMGYG2cssdMXiJakGW21TA9LP49OYk8B21LZ+V6VR
0YuYm2cs/f+765Kbt6Hda3hXxG8qMDrAfHQxhgYRgStYc4U79n1YW/CA443ATXCa
hmI5862DqszY5dkmvBaG/UuBM59ZUrMNOloAzumb6CQzYyAapPmWyLER36N1/F5e
N5T0/pncdJkn/VuCY9CfESsRmDPn8v/x8Zrf6PHSGKHAYMeKLSN6hjPzygZcvXZu
oq4BjSygRloknWd1wjkY/0itTTJkS4WT+jNNyvQTq85n+5hMc0BkZz6bNPLBmDqP
4CkRzoakszVeg/zPBt9ZnegLXfH+B2a1CYCyPqAYi+9nLSiPNBMZrNurl8UJjJRt
yFAU7uH72qCcx9JSM4n1M+p02XaUCCNPcaCW2mH4WGE/ITxvjDt/caDy5/0EFiYk
xIuPpI081m7DnlX0mlH/nz6U5gd8MKUpxAGUHNo1HsElgcBcmNFfX4DbpNoudyCH
UbdjheN2f4SftDQvVsfApdVqnL15Ajqcx7sBQtwTN8BSHwUNo0GaSyejYttvPsyz
u8T/fdg+xchbsFG99RGDO3/U42stSkg/G5AvjRroF4ZjLPmaoPiAFDNFAz1Qgwo2
oTW5jvFYeUd99U4fMJPfnaAjQsUdGOxKHp23kPDdNeZm16pAzecsFVGIbPsRnqLU
oav4PtUPC7XHPaao9KNN9huaY0Fjcs8DCh1WyveF4f77HwDhk82zGXV+/9eHWkaG
66DA+fL+Aq01mtuCmZ0I+C0haxPVLWqOOw6oj0hARb+nRNoVoiyuh5TQGBQrJngu
vKB2razO1z2bBvEsajP2re1GL33qt2LpdgxeMrxrvJp+OPywajPF2s4F95hV3r84
SOxGJ+q1evq9uNZ7jOj3EFfDbehLCdVhL2Zjb7M1UJfdB6ta8B35l6poaR6ukWHd
Vuqb4I4az0+/Vz7cIRRHK+QkPQK5cmzMBQGIEw5022/zmw3fvLcHcRT5nst1m/zz
vxIaUAoEzFCv6FmajAOvMrtkcDW67hu6eAOM9qwnve6N9eFDQnSoPjQs+vtdnQrg
cXUIGm0vhvUq3R0TTLx6DxBbH1U6Q++cT1Xgwurj4QdCMGsaGf2jRfkaHmLPDQVK
gmak0qQI7H0jQctvesLKWKBWBoVAY8ZQs+DON5NtsM0vn/px3REr3wW1stYMPNor
iXVI5/OdbCHJWQX22BOSCzJWrPZkulSUUd+5JqLahKahnFA2UG3ne1KnJPiZ4Y4L
UJiISpgfiBfh3rvUxWmnwEEbi+aGd/bqax+lC8gZ3h0wy9tdcCvEWEXMkTSEWMsd
/lj7LPIOqyJ0aLL7lfxxB9la6/EU/0btpNPCltQHf35Xda3TgkCu5lcF+VidZFSV
/vA2TpviY4TDCqPM9VvMx8YS6DMYELbOi+Nhx9kxom+8MNxr+H4Sgt9QwZT8N4hl
PNxXWAj2d5LYcyXYcxS9xcd27zy/VQ+nW7Vr5iG56k1IDjuPD5yP+SsGMH/bGC9o
SZ2tKtmF0UU27tCmjROSUBNhFMTzCB9+jg4g14u1jmFE1OukALlcwIhaujqQsd73
h6mrZ943HHRldORm38a3Y3FoLQEguHA87dA64+RsZ7IS40hUI6RDRz7tu5SvftE1
fMqyKFy2CRceMeR+3in843MsRLgoQ7rw3NPCAz/T5/MNHcMMdJLGHSgU0M7Fhzd0
Wn4oN1f1hzm02NXraf4VVCvd3tAM4+aIIjhpl30egiIuKPXnLdZIlRPuY5StcvHe
Wl7KHFoJPNikdVjRDrSyP87PCLl8J1E4njNR8wRCMG9Oe5eoQrGIwWxXqqPlE5FU
2LFGzrIndmfYrDH1VuT+2xGFDKEOMsgWfx8TtNuupC4BIBSpVRKG3LybQFSAptuL
2ghzAFqD0KINzjNZ7aVyHsqrH+WPKl3BjEBAvCKHxPt5L1Rt2c85hH25GSt9Gdoa
wJ/p+hpAQIP1Y3Oawg3dI3uhPzRN0pUN9980N7703ziEYfacvgE02ITz/0JIMG62
9/zFDhItRS0VVaKMYa3TG3GaHX7PxJLE660twwQK5XtERj+BX15kgc7lEPiyCeDS
XpBzOjNq9GgVuooR/tWOLbH6h5AGgm4uIRafa7wuR0xcndf0yaNB02/88uW41M2A
wDshCWd/JpRYkAAEMCzeyy28sv3eLMuQPO8VDKRQdbZSv0COUL4YUKOADKNyb0kb
7ap5OYAr/+lkvBkplaDDpLf6nhEAFy7y48uvSpC/e6SMKMW/oHxXEyV2pagGBT66
7C4rHiBdsqpQ3ecIYOr2yRDY6lQj9QWvwTk4/crUFRs9qtUfGejVa1jQuOCWqRO2
PmOQTV5pR2lN1QGX0Qals0dy1KkTXyf9W5AqnDsucYhEkpi1hqgIAa1nwzHnmrF5
3WW33CKRYEPhUqV4ZM4GgX2D+aSPElmds80cgKGopWi1uL5JE4EjgWugIbwUXAsQ
d+H7DRBWU78z3ayMIxy6T+RpX176t+RXoh3ksz3Z4v/C3wqV7adOhAVdptew85qa
7+aVe/6oZCtl18HOHeNFCd5xiaP+NGMJLu5miaM2EtasQKSSeTOnkXyrc3H4Nq5Z
K7eFBVgFQ1jN+HHjYzqZwA3gPWfpIfwijadM6L77pv/vjnmV9J19PIkiaM4p0MYY
4rFhVd8oGOBA9gn+9zGC/BOsJVwu6W8igyUQPGav2JQoN8PTeEqMPmmU7Lp0rHNX
J1qyjT/NvziO2aFktlxq9yBVvTZBsgTz8Ga6q853NPK3lurnziegzAJV6SXBzfH/
d05MU78i6AaX4vrMVB0QJqMAGsNsjUmliL7doLWpB8ZsJBYhHpDnZZud6qNVtvQe
1MUfi2KtL/OhhHM3Fpnxht0mWyYYIzHMfAb/15lB4JeW/GnAB91b4sfuDtbWFGPp
H6//Gtf8wXf0ZyOPY304dnB//jHVug91sH9pffG+4E4mOM9ZUPjf+EIwB+9+bt70
e4uTZ6/zVwKWm/ZC7gAie6DjBGlTa/34f6BKAmWmK4DjDGt1e8Vn1HNUKxehTJz9
JHsggdqviJp263bls6cJwaAolfdYKAkuz/eBTeWLyvsOwKbxRskNQNnBStZXvzu4
ZcgZnsqfn9yMLvix5BmM0KS6oG7fMiTjHjExkHnRIRvwUqrpGlkOWVrqJ3qG+RLv
ZdVSM6+RWO0HBlwREuMUtXtmCYzO5IFbtgS2bIkTYd8Em8qYbHGpJAQivpqgHNU9
fMWnlVuEki2GheMVeIyDDf1N5VChMhD9rqqIea95cNIN6jImbL7czsQ1PT2SBELh
5TzpN1azDbInA5OQ9EbxytLLHgwbXskLOiYMu6UvQVGreIU9uDfjxsLeSCQ0sasw
Kv5rKHgIEr6wkJW1RVwa1+p04R0ipII5x1CM6v/UIqAaZDMLYpemliP4H/MIhj0N
aAZjsApo5MlM+ePkvUoy9vc1ad+hsegPxEDg0Giov+gHgAqzZJr65Ao9qN2jG8E3
n5VzT+czFyh9tu9BlQMq+ZnS+a3Z4YilQyPj7R5NCYoVF7E51lAcpvayd6SLhTSJ
tUEmhobDoSoGTdhbJgP6bO2bMsz7dlBJyUyRptFOYRq+N0RZERFV+sa3BevSA3gk
/0dEI1AXRvdC9fQfxMcwbsHwLHVuEIHUVei1bnxc9eNkxQtWmFTrRIRhdKFk6vd/
y91CfLSJx9Xe7e+bxWzluti/eisucPvZti9ioBY7ckOfT45PK2n/PKug60BZpKkI
fZ33PUxcuhqNQCesGKoJDgQfHFpHe3CaHS9J3qnJM/uY9N3tIP590wnxuQuDXtFV
JqqkaPPQkv8jpmzgHS9OEXS1qQ/30bV9oA3l6cE+EvR/iQMjd2dplJvuELNbCZcF
0mh2A+r/bdL+ePy8ZvFH2lMj+rWgYnuPhdgCUDEaOHWkjAIY1NnI1leJD8BZASGn
2PMkYNmtLGIXwwXduHLwgsLVGulsUw3NGLrw8a6fxKSc4rk5IxI59sb+hM8YLPNH
wg4tiVjxwu+zlLy6WprNssPUkAJ8y7+OsOwoG0CWNih1WZ4k9R4dSGmqOsr5gvTa
ZL/FUyPAl/3HthzWRfLmKsEpGh59SzWhh3gQoj2G9uACjmd31dNOvw0Hb/TbmJfO
Vg57a7YorWTUb7UI5+TlJH5bYkxqCsekpBuQYL7cx0Jfdzp9uVj9skmTuw0TWaTl
A7HL6IUbzbJ0cjKW9iNhlYsq5xMaBq90uRuFHJQyYr27xOhI8JBT4v510Lv4BvZB
D6CsXxuvRBaTSy56/zVAv8gFXdW6sAhYjzRsZHg6BdhhuktVkGOl8Y77az22fIyd
9dK2MYtXxY/PgG761lcodqN5cjgAI42SUv3gcbstFvsgycuqK2HND/Ad5KYUyc4T
qY6a4Sj8Cm3QQDwfmY2G84+/MioSMlrFvqTK9lgs2/H9IkQE0dKJYCrZL9pU4xYv
HjVA26o/dst9XehpRiZ4H4HFKcVVd/c4XqLqIX9hjk/CQyin77QtaRlKZLkFfxpP
fgBExkyduMW+djtkAP2uRPrDDdcihSeWIjbxaltWKmPm0SFJVrb5DpEEpgbdHnVO
9mBidm9AISCwZ5gcdVfuNd1eeDMZqwjkEelQ2vlFZsf3Y3rbd4hIevmMvRDsGGyZ
nekiiu8KU9ZFf0m0XukQXgjfmQDrgvHC1peunWeGoiDH9zA4rgEJNPWufAZep5FU
/5voyrqwiE7a+O75zKFIDo49v1SUzEewX9ifmcnPbSvsH7oS7CDS9jL7wJclT+vN
u9cJdh6l1K3aaYRiN8cIJCzPYpYBFoT6Fja4/yrYcHLt2RtOcUNGtXXwXd3QoUOG
yRPDtWTQkLYHUrQjN3pTz+DdX1rOXkGu/W75aOUY+WrWkd2Icuqha4vbXZ4HC/5j
XG96ip2lWtzU0w55nhzdduIHBo78CI/IJ5/31a2XwOLWeXWiE3WCdEY+LyTdd5rf
5bcghEf+BHCax1rPBF1OTqa7PzALb7ZxwqLx8GTidmfpdRXpZuK43b4sXEdcJTeq
hdlvayyBrHg1KcIlnD4z643oPpAiXMDuH3JLM7r+NnYhET86jdp/EJyri6t3NzNL
UYZl9+8Um/PY6Zx0/hUenyQJfV7SGfT7e+0PK6APkDVvLKCFj5nhhsyc1bz/pfxZ
g+cIy+wkUoeH05WWpXy4L+yJkkQv7gx2NLEkQySBQL79dNpHuoULt5FLKS3slOMs
5z1psutWq+HmYW1pZ5WH9MZjXVDJ3qHOCAyyr3lgRxFJMDkY0duFJTzuYu6AzUFe
Ol8B50wj15kl2U8mbxx11DT2+gpHyxVt3ZaKvitKIhwd7a8z0ymcXoZ9tzSgF+o5
d4H4sgrZ/7vCkKEqQwWinfs7klLtMzIG95jf0R5QESEMnLJJO1LVY8Asj0p8H8Bo
dfrKfVwM+ED7Yl2iPbkvuoKLTVJMoouL0IBv+AUrKueQvCebsdHiln1YaBNEL2Em
jL7/hJwFppLfvuofK59g0GZVT7pczO+vXX2CFBwdPMK+DDGOhCxmnik/mPE3cGfl
5D2f99vYJAcm119yMg/xvPFJ9QgdbhOdQNDwRwQ+FZ6aEfInCc/6kziaBcEzwfe8
kQCpby2urG3w765dM889KexsEe4uvHZZMfYtAqBWnG+58mTuy/RHx+Bl6CWVnqUa
o0n8/oIogi+0sFsRtknUJWCV/1zVbjfKYi0TuRCtU5W6RUpxd9YGQmMD5F3sZaQQ
awYDevJiGMZMeTM8IssHvOYCCUaRMAkOnocyhV1XSH9OLK4tV8N1MMkne/NnDNFT
dZhQsCwlf4ZqcFCDeQY2WAaGqDpZOhJcTlYPwZW8Nz/XSTkvQnAjDJ+7+YM4NfXQ
rWj8/flKk+fJvNaZCrQKEpxXTx6Zf0R5VYeIiUHxSHskT7Pavo5Ey5jFPV9JHnlG
J4ubwT7GRfHzdUDqkXMJLxWSsSofAmELeBXByZ7NwRdBhP1zKRfe8JxvUeaCJFnj
6qcl0E/N7sG7I9EEibWBOqUkUzavhsVRJh32UnMRfdZr2LWTJtbhGvtDD5U/ahda
96Tfpnzu6wwpcAUwiMFQM6H/oBDAFiYOfKI4mY+BSDP2PzT+68y8SvAL51lvvzav
ZxgQVRTtxgYWZnbdk1ur4yKHx95p8ztw9jVr1OPejE3wJ9edX2Cq+A7IJ/ltYEXu
voUQoRpuc2gJH2KAdDJvXuR7/rl5WTjyuINIyHlf6TUB+VFIsEDXzp0YUxwgi6AD
dMx8ZZgyEsvvSLGHbNFzGcUgfJjrm0xwlfzV+UJYWe54UQgPxMC6HX9nSlKKdUNv
rnUmhyiSFUlvd8fKn1UZNnHtOgKZ/J4Gvr4YExaNOJXaEzjdB4jn62MY8C8rs81n
6/Q6ugLUYHAxFE0eXbo2N70OGOrL2kYfvuyhQEUfs1jCYATe532xxE6wyVELX+Fw
CyeiktTssRM9+TTarJRsXZb6pDnRSoXu6TuoHJ5MNrgg0GM+XbxBOfQu2zPhx4k4
jVJytl4SYZ5eY4v2gZhCO9+YKx31WlWQbAdhasKlGmna8ITi+9VkgBA387EOV8ld
6nAzUc9N/YbM9qZe9o+O8Uoi71nr57lghaqWRn+7hqzyvz0f9jijnx0oXzsKxrLZ
lnzWN7t0WpKMtQck8wEnWnDQ2TcpFK463xkfQ44LfWp2YREQd6gsZVdIb1KQxEk2
SvU298CrkCmSwXEA5bPrZ2UiUXdAdR2GtxY+n/H/NJr5hI/nqbpdbbVBKitTKKDS
cpgc+G17s1extrVj62mFH5YH5IZfQt8RYOudLdZDs3tGYy3XoMwMvK1i6J4QzJN0
m/9y0C+kQe9OHC7LOLS3kY8wpFP7O7lz99wa3CeZ0E+uWTCbKcG/PtrcUt0YN78c
Jmbr3E2hbDDPfx4PiFKXDWhs7uMBqjhxr0EZXWsS8GPAxWNf0dgl2YbcZwnpZzO0
foOlk1eZ1K+dLg8yKXDzHnBIEso7mxb1LkrlxKqRZ2nQ/jgypPP7NSqPADR3pK5+
c8owjbEAmV8B0Ae+A61tkxkI+70KdxxH37lyP97nvwsEfWxg0vsU7V2v+2K8huM4
ehMnfbVUv+3NU856XRdbiMabMUHInp1gWH/Yr9qqNfHPkkNnjILrYIzHeKIHE+dU
v/VYfUVmpBZSBRpTWu8YUMcG1aDuZ3mcPgztGCK6sQDyfqFZd3Q/af3LCINexC1l
AgioSwa0tKwHA8j6I2vKuPY83N9V1zRNEgPNNapeNcVa1k5c21WWae+BCd+DET+g
yBPP/DQVAT5JtPzZe1zbdNj2D6//12U94Sq27+/iOi38Wog+Y0SYBe9qkxfolWV9
toJ1eWPQAvDCQ5CdLVVqpXJOs0DPqZJ8XGb+AHH3CvA8ZONBh8vh0h16G1DkIf/2
8lB7zR0dgRQ+hQQv6kc+gY023wxiSYP8UDgC/E14+SSIfALjwq3Y+1gJuNFZ5ypv
zKRNfoGk1dtu8cM0zls0BnBzrpcKJwQOJ6eB2icNbI2rRsQc4b/CbPBWCW4Kqp51
GyHbNzPBkkVIlSbVRvjgxAiGRsF4NOBalGu08jDNNis0I+9gXejugOCfCMAOFmgA
PLXOjIsMI7DPSGamVlvztT1jv78VWNyTMn4dtov6GtF7E4P1pA3RsG95AR0LAmbv
Bra28zV0G5zI2WjLfc4aOHkefXGkEGe4/9YFmnNXrMRyOGVuvBSyo6RHDhPN3Xqy
4iFq22J0FsNN+DgkfLTXFKpsGx30vBTOo/AGpEUfdbyNAqRhNi2ZUseD5Gfr7E0Y
XlW1kny7IQKjLb1oJxwlDGNhxROlTYlSYE/DtfIs2OIx6uzYl8Z7qCVs4/C+01sD
MRYzIazV4VFdcQHyhw87p+4XdE9TY5NBgEb2zMxWOHSlGZDgVnovr4U+gQxQgQ/O
5iKgNmgW6PVZIakI9I4NX/aAS/JwNnqQPmj1p3aBFZs2iEjxsOYn2mdnF8+B5HDI
q9+v27MlVvb46UUYDF/Y3bXdHkjlYX/HPCIZbMFRZ76sJ+xlI1d0sAWBjDvNYSg/
gBzN2jFRQKz6K11BWxQ5b4vpJ3wCluWrWX56+cGY14vrueNW9tsWEVbCP1JGUNVR
Fwl0i1cGuymmshl+14e9o6QPPkWusFGCraXSwtVregQ+mLutuo2FlPm8yvu3rEyg
5SX9HkylY0hsYLaFmZxfbLECJ2VsDGSkwcnmScVFZsvG7loiSm/B0r6LbTRSQ4aR
9+AkJZ1WP/8v91+Zor8yE9wRAd5RPKHDSccqNQRE0D9Rj9xb8CyqCLNVxFIlxb+z
QRrZhg4s7pm9qhveLgxpSpSoT9B1CBOa7HH0DhLpmDq+LKGsvgLLxr2W2R4rmMFR
8hIklTq1Wm/Rj+eVUlu0O8UVuR64rcPjVRfSrwRJLTSmmwoYB5tW90WI7l0k3G1V
11kPlLu2FcAQw2LIeno3b5RYMzc444yiJUDU3JIpp4LS4eEe6B+xTUnlXhLzzqJX
UuoHEe0TkBd5N5xXcqj40w4xLrxPACE8jnPkQ7bC7mjbr7aNGWCTkELoi1EI5Akx
8FOv8aazeSCPf3US6rPgmuoXGVm8+IqycOj7rJe8h1o6ndUJkMne7bITqI3aG9WV
Oa43ojE50M9QIdRDGuQfwkTShAbiRKRB6de7EiFfrEubGee/bzADyPxRpvfns3rA
+6tpkKEHwQi19gaLdGQijaQmoOZPCgq+8EAq9bQ2+Le6FYGI3hFdStufggYX7ieS
aO99WOzDp29yezJMwyGaDgR0nDCPr5rsLFhdk2h58YrUBhRXEcftu9tDUgKgbfOI
sHIqKrAePxs6jeIkNZl5ywnYhev18fHNEJxhTtF247IuDU8oxGwFDbh8tHXJXR2T
Xe8KVAdNOw2nrlhmN/SG37mfOKTgSxuy5vfWFs8Q5vwRJy+09RGqC1A4/U0mV+7f
LR1VK/g4/FlHYD83ElSXFVDY7J/P6hzWCF8I8PnPUtbQjMwkZ+NJcbRFMUJnCPXp
LGYPO5jDx7MfBVs37mK001AhgNcc0y9vmVI1pA4pWxGmgNdVRPHx+7xNjIlmdHPg
695YUQmq+Tqas5d0pLHlrwVOX424EWoEeymm1e6SApONd/05B3wQWKCkGfgHShWB
d7sYuKIIjm506lTNh1HyrhP5ubwMLBf3YifPa4afGlBCoKTeekjpdaPaiXCImRYx
G9q4QJ67X5+epowBiAhbNTBYnwxAg1iYcwxXf3sMyhXyVCeiGRvmjIxJhQ7X2uje
lp01wNot9ZrmnE92WSxT2BX22WawOn7tSPM4EMAWuV2iVZwVN8wFdaxk9z1aHyli
02ByH3GugM4VezXPJ6gFHubhz4jSBnhp99Wz7DzxK0Q7AFkKHjBO4OEc+JOqYg+X
yia1YvCUHrmiWlJ80T6s/Xq/+Rnj0XxI2UtySK4igwNqC28S6wktq6M/Ndz8Mfoj
yorNoDdEK/P8XCkqp9+NC/ATF+cpAZXuK1X/OLqU1g2fvOrdwCGepskYQAz7wieT
XwfXz7vT9Romdlzj9roJPB8daQc3JZO9CxisAt9W8qIlxIsat+QwqjXZI32GONmh
fZK4IuOUMI/CYQ+FicZdUaIp+Db9cKYg8v9gJRpc4yDpDe1gkHDSJJXppxrFU3iJ
MwtYqh9QHFo9JEp1DIrFfWCuq9PJfPwlUkXPZX5MBUuTeIjA7HL/taZLQWCA3YwR
LAErvTpYBcOROmLRPc3IxSsna9DdRuUk/jr2b9g35tWArIbjmSpeNKNjm2Elp8bC
yL8kOiMdQdljcHV5NOM5VWVduNGi8YRvVFWJLdAXFkOsigsAJaZ0KophJw52Dtvu
YINb/kTvplHUjQtYXYNayxif9prpUboSPQ/7DIXOskhNuxYcc3tauokWs2y9Mx9k
Fi16tMr2LlLlFCRNT8K57Q29XDG4WtURdBdTDLjCFakhOoyBqSaVnVQMjivEWlHm
Azgq/6IXGNdfWuXB9TNJg81ayBxLBYLtF2xQC+E3G66P1DQfr+QApToI59tZvEPL
nJH3oxNRUC1bueCWPJXl2an4y628y0CKZK5ZbDo1qYvca6KLMRNGDP0gQfkWgwYe
hhz5BaVLBnmspyxhXOzTpVwMCVubhXE6rF/f5esUt2TeRCKitGQMS++DBT9mG35v
ThDSoTbsHtHReJypeAE6sTWwnLV/TEhZqQCK/xKErDJwtGKZ4ZGTiW6R1T9NzzgT
Al0u5BUx3GQrw/YAo+bTdrbJjA6olAUtDFbj/vnbxdsbsKSOrFyi7Hnnrg48r0uT
OnnZxIxu8hPwxs+17/vL3Lyey2zXDunoSueWnu+p/7/OnQnM7jBvbAuwe6esf/9k
iN1kJEVimOK4Bq+JMjI/Y8pYsk/FcF0GZOHhlsQ/lZANowUzIUXaphVvMG+7zdya
Ih6AAnwhCU+xqYzrP1mRU4XCnNXWEi2+T6w1FAAoL3lt0gUYPgr8tog8b295y0hR
zpqhvB6DDofEeI/sYlOYshLg7AU7/GKIqAUpEwk8/ft7VkgvjjrrH9uQD8MsSTZ7
6To6NsN+l3YBI7oI07b0J33syPyQK+qAt+BJo8XgWmjmwLGSZplc1lbosF5rQpGp
RRRRvua61+i3CvTFfSic6jKYQUN7So4c0IDy0VHjx3et6GkobcbZwS2boNrVBEqe
IaPOawVATqsApVzB7rHL9oM3x+VqcJX/e2Ld/hl2efSRsMv5t6dBcZALBKA/3Ev0
lKgxVZ5/dNlqYCKuaU0EQi4dEzerO1KM3/M71lBlvRphSf7pvWIHPyLuhZZyq3VP
noTId1h8aWmhv9Yj5rP5WmmXbSiUevyXRmqNZwNIXWO1PObOSguELh29+JL3BqUh
ZrCtASqbAD9bsa5dinplx2YQlISfQjrD7pbqd1M6XsjBmI9H0BViFNAA2rJKYJj6
31fgAvU61kl/JnarBpJvjP7ZYNu1B6hoUhshvpH+TENja16HJtRzeAg96ElNzI/3
lrlPc1QilOZKZCcxUDRPV1JgoUE1UinE3yOHqWt33RFDBsdmQ57QHg7stZRyvsN8
tOtIJWIQREkVH/cyk1LFW4G8UYEyO7d3c+gzUmJXUV+T4yC1VpqDwhyorVc2wS4u
dWa9jHYatDrbYH80QDi5URhaZc3z2Zy2Dr8nDZhgv7S7tCAq91Ct62yLHTn9N5X1
F6l9FjY9viqHNa+A7z9DTX1aouN+0bP69X9agk/E3kFYcrwcguBqSh2mplDVIoVt
dsjfA4gDWk/vJ0Q6fKrR0Pg8PioGMaO1JGRMwPt8fpo6S1Dm6GFhqw+M9O9ama3d
sxOyCXAyrI6BFdyp7zAzPE/dtSRSVWhmKX+yMjSLK3YnTTr0xldJsyyZpGcMBtst
Yord5WueyYkeNfqGNjxhOLEC2z2ULEQdi1la6RALWo2w0cVgECbQIl2irAs+fW5i
sXdbQWi5gjI30ExPr1Nzga0aIjXoyzmMW/IMTf6d7HhIkfHT0bX/k6XfzLdQwZSC
ZD3FO0nwYQHy8MzJqPdAxEKTKkkuQ3BPZ95X9A/HhnkV6A6LFBXJ83vL7rsStOEB
4Y5yXZUJM2E/APqKpxnwhOrRsSGYkEU6fXZeZ3OozWyYzbT+Myv5FZu2SXv+kCqK
z7ytbKpdHQOsA7A5w26IPnHEzpE3fZADb3eVvwHrp4ieXyxfTIpPUpT9izz3nUC+
chdwyoyAoC2jtTlINwYVSIaQz9eFjoQrk1Q2l0HkRWpKtkmDK3Fnm5ovwtQGIXDj
59JhAZMuGvTd3vFYfnJFlfrHTUcaNzPRstpPfSa2RV05O+ZZ8RlfCuVVQnNaA6sn
A3EU/mqNgtfX8t7ZNkqJVHEwZiiZXIfob5qHDovADQAySTu3CmTk7trSvlGCL0Qk
yCdOINPRI4txtptrLqj5N+Kud3MmpA5/n8wKYWWmHvie6cUEiNMdyMVnkorMUuRl
3zFu0nPAY42rlb1K3kyrlbLC6s+HrzfrIBvyjOIm32KmYGakCOQ7oIS29pK9fp1u
gVpbMFBFoPuzCb0wzKeaDznEZxcES4+Ztc18FRaVMHMpwA8rnKUm2Jkq9XbP7HsC
q0Q7qO/Kc36eyVrb1+edd4VUvjKbMZVZ2AVTrb/y1CYPIKJCQ8flGt53AX6s/F+u
k/Z7XH1WPMCKNd7zA+Nb9rK2QRKmuHPDPYD4sxi3iC/dR1RRJoNL3u7nbmmiPV3S
CcylAw03oxzKnNCrppAKlNXjzlzxYa6sKLv9xnEngTrpOriqh0ywpOGKXn0bb12x
vmYEdjec7+m3wbQTMARhenz4vyqlhyDe2l+R4ZUKIsTvney5brVbbMops3zNKAHY
rJmEqtm+CzOrUYY3jUHZZ/S1NLG2xSRkY0sWdUmALQrKDtbke2qZmspVnNUkP0Wm
caHoskAXS67252H7SIK9hmOZi88S7jLhYZodkO/wVnrYGEuVYd520xRPVXEXu9Cq
Ah/0owVKweg/jeuubR3ez6XyBDtinlHSDhXJm3LWkgETiFXqI8UpuY0k2nQTiYmM
kQYwFqhFewCpQaU+0JwwebY7MIC6MBWwRLcgTrZ+Hz1ecrmWoB5MK0UdZRvrYi0m
MXgylB1b7mmldeni+dJWZ1M4iTeLs9GgynOmdSp299e8UxoThmARlld/L4/LR1BG
kVRR4no30VMIj+9JSMsRXXgpsLIgpOMNU1kK+43htHSUWxuJSEwKNH5I79hVihLP
fDMLXQEdvm4jS6Wb4e6RnhbEX2zRrQ3+55eMtduwPavaN+Hy3yOgY1NXPtuOySxI
FKeLEpkpHdJcbyCMulN1YPzu4TR5/10vrSxq2sxhGG937tBUAK1uYtZLsGYDGQ7X
/ncOoabdgLuW/AI7V/CYQSOKq9cTHb4NJrg01Arpl1dipgzXztFkjaqhIIiTDP5x
ngGiPC+ITTAcJyuKrb/2enozoP1+EpHZAlgEY8bWBt1/nxcsm1AIPaaH5xOjuIVa
TmmCq1kZaaBN1F8sJkWNic2oRWXx2cGOZt9dHiXV/XRhKb9qRn0xodJRa4JLuhRK
mznNRlEh89c94t5oPR9T3r9DUqzFAR5pQ6hd4jxmuq3+t5XOkldwxD8RzRd5n2lb
6BeKvBQaR2MKGFO4A6vpeg2UskgZE0sKIErPR039b6M3G6/NwCLJ+7MZqTPAgOYg
z69Hy7KqwZEm81tsIlP3bZPEgIiimLE5rDJI+lPZfrJGL6vUiYM7W/o+2piLzs36
w1teO9806sMZufLaEc+w+2D11i8obA58QIUqv0RAjIWRfOQRGW0n3HXWeVaUOgJC
9HjJMY4xWENEyGNJu7pgpjDKZMdrKuqukfx3qBVfAPy7hfJ864wO51pzNofB6jpX
ztww1wSk5bxt+W+eJrmPA69mDUW5qWJbcLHqB3wTu8KBk5x6/5DM+D1CLv3P522I
nyI4C7qLoDbiL7JPZaWqo/NicbBZ+2AndLdgK+wS5mt9YctEFs/c7YGtOkRpSTaK
mA8J3Qxqzq71OK/2SJTM5yKsvuHtClfoGBzojz/hd6SZASkT3aWf8YDYsFsYC+yU
bAqzBfqq4moti6D1N2umpkOhuDuVWD+wWiOtwxrKFUO1bij8u1Uea21KNdcUTGLT
TrqTsktQvmMOgYQvB8AkXg/k8KYYVh4Flg2iCqPw9hIRpNvzrNZqGfFzKM7RlSG3
8lLPuUm8Puy6CgFbGUMKIdhwZAHNrZpwPoIjJeDnv4PrpR4OsrGpQOzAhj3hPuGP
5bz7D1U5CHdJJGaCcEEp+X0RwBli5d2EsNMwddWQUtPg/A6wGpeXnJmRbDBPtBu0
+2XoduMd8ZvPzyRMPOFBnK0rab6ym6WcmaUdTveWqRv7j7Gmpm2CqfqT48K+eil1
5foZ4iRaCYIkpKpAx6lAhTakk0c/rIPSQpIdrzDMxAWVVV7bmH66q0u92RmZXgWh
WqknJstWsrBuwvaJROc2jI8NyFREl/dvGmaOzyv+QjLKcTTDaoDkMNH6QsdmVsN0
ts8yrN7Bbh+eLbTTJhJe0nby6T2USoLox+TXn/QpciIAEVVzyrpv5+3Sfm74CSnv
qQAD00zvFU22x1jFvnZ8cuy5AWvS444fxldXbeFVzo9zjku9X020BDyrmj911lJK
icbMnBgeXHOzeA3H2eELbzOaqf6JeDGIEzi2vXpzIILmmWTZccUbw3xvmoPn1hGw
YEXJN3m5Uh0YhqnDuMYLDHfGYAI+mrqfWgWbkpgemv5JmbXyWbWPQIjc0f2pXb1q
d/PglbaBOK4fSaC6FANEAertbY1vwjs2uWblbmkOB4g5DZoo/q/5327nds/4mttX
ToMJ/8Oe+G60uISeBhuMByV5Hb1RqOOK9C7sUC+iD9Q+GrahhzBwmWyjgCemWUVc
NKJFuMeaLzC5JngIXQsAKLP8jWilvL6LvxRDCwzWV9wovqGtxvA98TzitWehyB8/
M/U4j8mNpKdkcLjMurrlgq93b43kv2hMlo0qnCSEc4TcEuEu1EKY84DF6RC6Yyun
W0LJPeQIkeDjETM+119WTHRoZ8P8WTHwyyjt0GctDrWpFYwEdtoBaCHCCh8yFQdL
wEpO0cNDxo0WCa9QaMEPzMAlvVHEP6W6aVPQ5qeqrqeL9JWQKzYuSvT4o52Do8b4
DcvgdWzko+nvjrW1yzcP6Si64IdscuqfxcOhQt1kY0jbI9JOF0M1RRUJ+d5h0UqM
iOkB7lmCgLX+mEzEdDPxS3WmzOsn6ILfDUomIY6W3cs5+fDE/fjr+eva3MWNzkh3
BIsnXVUHsQaYlYLsWg4w92tiRMWz2MiDyLm4aH/l5HQfZT51zxZNpF6I4/idL38V
hCJrpw6NdINUKseD2NkYlfG1zbXYFg3XYE7TSA+YEnRaa7DGlnblIKk7m+Nex0M1
85/4fII8rUgzQhoOBZLpLwbAcCkAiv4KEbi2lKZtPbp7LN1wB2OnXl7B4i7eq891
1yFdR9LZ5Gxp6P0EvGIm18vN50Uvwqay3+yIBMC2bMwRT6yCOoFmu3IZhCWV27LK
4iWKV7Pb0a6BU6xitz4jWh35xS3bqCyzYEMwtxL8rwqqVcarYODFvV8h3S+4/QLR
9ehAfNH/KAnMIeq1YoJZJaZmZVL9S4HTAdNj0B4VVQHEQQhOcKAHlwrM3S5g6spo
wYo7W601iPhVanMZsg4RdDHb8rzSbLEpBVN8ZEnQH87BDeRgkr30/BtEkiJvodtM
LrinA1jmXQZYp2DAIBjTOn4mOiPmZXvPsX9086J79FqVQyT7jgGVmS3jqnVfdb/A
r+jPS6g/t/xvsHN0va72KuISpy4NtT/vSB5xocRvYXmfyvTQljdCk7Y5ae1L2eCM
i1u+9tYpBYwISsUIrlZitump5idLxNXPeasFwFRaXwMCLCB+zjxiLjoZynvSpB7l
r+X8bUphW/pc7CkoeTp/EW3wAQ2xqv5YSBiLXogSIOlDSft05NRX6b1cOKe0Drea
0YSLexkAE4hH5E5x+HNwmcRNBddjuc2yYbKNRF1JXNc0d1xQe57VfbWEJhvnsvk6
ulCPLvFfkCSqithFlIDaNKHYpatxSywNGb7uPLxVZ6TbNfWDyKw4qSwyNQ5zmnG8
LSQ3NHoaQ4Nix2WyVUYGtCdv7lc0hpugYDtfZkbK7FDsdCXWRzlbdhdfJ9qWS2Xc
/BsXCi9JIchGLLvU6ic2vEnn6QXkBm2mOL2NWZldyHBDx96pCPZ3/GUbIPY2jLzS
RUinJDjPppKu/D4x8thWrYqeL2KkMnrPs1CYH19SjAT+/Pt6gLa6cKB7jvwfeEaq
PMSdnwp3ZSmhjp4Z9h8b+MoC0cb2oGPby6PDDipG/Mqscjar5JV2l+sboJYVcXQ8
Rk2d+qePcg/gV75JZ3M1ssZ/MwwIxquAfQOTCSjg9n8LdiVrSJOQA+gZ3LGn9LcS
dLBIQ8iXrY//iLe2bzP5wfryeWio6OntzIb3BkgB/osXm7rKlhuKdHu2kv5bknh6
rHc3ekqSiQnJUppiCY8rZ/adA5tgRAAQpyo8jva4b5Wl8bBG/++vVn5BlvjC/uf7
xWlJ/L+MPIFCEX6P3Oio+uHBcKQtWQywtJNYhVDBuUrGOVaavIiZFIOHDRZH07HB
B49VlbWRPTBa/5Dq3InSILz3hHQR4Qg1smjjjvGo5fpM4qXO2DG+MAv0vOZES2cz
LN3HywQXBHDasohTVTflvpQA3e4hND+RmFklVubUBvIW6ChdvcSWboV+BqFRxHhh
EgzKf8nVlWPcRWsBRZYX6c1rZ6hqZIdmjmv/cuidvVPNFbuQ9u3BzMQATvkonNJT
gUYha/Xu/KhOJo/GVcwzp112T6Hlt7bSzZDPYb1ro5vPzZD7tz8Kn96Kd2hJbqkH
xCNTF4a3MK/XijGa8o/BlHJX7cAqBWHBnjoH51LZEFu9qG6JsMf+XooqlaIqEdM9
2ag9rwDb+TgqHrZMsG5j3QAa7HOdVTm1jExDcPHUhsqZnOtU2Kbr/c0CuIsIky3N
p7alS8IYkh4CA9eLHmOfeVFZfgyqtoh77MN+BU9SOn5d6IzCIgbXwFu8BC5vK2Th
RiofxsBydlbd/Cn3A37vKQmMlVBvuZ0rve+FlQbo5kJx6lvhvzhbqJcYgI6q+aL9
I9nOEVMHUlCgiSFBV0zlA7E77f/RIS5scr52J/Pcp+DVcS8nfmA6kQV8QbDA+UvL
HMr3Uccbuk1woXsd3jjm1Fks/T+WxNr2XtrBKLyT6xdrlttTacpJd2pwP/IrsQCl
fwGxlYdlkuEFvUS72RLkHkByP+6+t992nNEnXZ7NOVAVNKF+3LWhEPhZhBjKPwwG
BeX4O1XM5BUCkrow2Tvpfd/yp/nIAexev6NitXTWXABM4ix/bvW90pJcEdWs4LpY
1NT+NXJ4auqAhIYJ1rmxXCV8AVMjE0t7dUtteCKpAA1LvRI/qCPCoc7ImV2ALOhu
h38jGKrrsK3gcnQKsDQyYTohv5Qd+R4NoTGcofxi8lBpZbf+un+VoyLV+Gr9116I
aGQ4Pst6AreJbm9f0NxGsxGGHRrpCmLN7qvzk5XnzECHhFFhM1sKHgf+1nQSY3jZ
iJIn6RZqpdT77AFTNr4oFaXkhbQTjYmkSwoZcRSAkET1eK8BZRJ4xzHBZG7rFr8+
crZtklLvlGUKm8IxcEiO0vcaj4jYS6soDVJFP6QeM94QoekLvbGHyyfS0Qf9MtY+
vd4dUwGXI+Aaqdtcz/QG9UWHXpuB0mqEbX6+ISQDwSEVVBkjQvCnX+0cLjRUYuUL
HuPuSqWbTBOSLCmg7YjSZpuvAtW7mB2COj+2Lt5rZcdSubmHncB/TU7Br3KPNSZ4
1yhRQz6ioGmGrcSSV4C6CLls4TP0p0LtXJkHCJEDSfV1B11iV5VFswpb1LbLIwsN
KTIOy6q346mPCjcA0CKaJ+WcvxP/GD6H+P6c2wn9r/m8YnmrEZE1F1pkUv17eiP2
T7XDbPlTyVNbn36x7YTFPeW+QHTNXaV4RJUWWdDRZTJmriBKg2CYS3ghtyxtmq02
g8ltQVyMx6fKpE6CbBZwGcxFJORACkaNvcRV77EsQm1OQIM2+oGG9ZQIKqffTJPd
TZKrA+6AirZRHJqf2WH3nTVZbvG7fN+OSH/5dvXm5qCewz4yYYmZDJN8a4T3wJ8n
yQbZ8AUME+9KKwM43PNJj/dsu53Pg6ShYJ/zEGXPK+iNP5fxPKKNkB6WDsW58qVf
9x0LOLhEss0QHJs53ExlV61puG6XvdEV5epXAe/AobfcqkhWdY4j60TECWl32JTF
iP5g++5jIyALsQl04QTsb87fHR7haRGua1H0HQpituWKp2CRqi/t222SxdQ3Tubf
nHmIrLzg6eLJWRFJhB0x9fPV0D9mZeZM4z2ZJW1oqwNumUn51yY9ZCpjXd7ljHwM
W6eT3ogCaeRp6qud4NOod8flTWgU8/vDd9JJhnS10BX+Mgpb2wlc8nHQWQLJNz4J
NuP3yY7y1lECOj36GSO3sN7hunTwAA4hki0APLZSY6zHV2KIU9syRlcaBJm/7w/r
jjxPhCfkAGI3ixqEwcrdgI5oKkGiaxNOfpI8w3HVcTuMGdCydaOOgra+6bykWrqu
JSMVwxw4zJ82g0/KipCu50lRyFEUTGk4tXM7VhFgYDXO9nfSvuuJR+1dZfjef0pa
GxZBjalxvwVXW/zFOrvMEoc/hFY+EdNKBq+HDUv5ZM4218z5y6aku7snBAuGkrSf
WRmo06goX5S8nFwtJIwhfOd5arD/gxDDAjdVjKHStIty7jfHQMst8plIpVGT9McW
XgeTAOfy4U7VjQJVvFORgEI6qj08+3pEx9lc5q8JwybO0JFA9zbNcIRJLR+MiYNV
L38ivKDmxonh00pmJByIIe1KMCjgMWeSN031yvZhqKFI2cKelr0bdjweBn+dyFu6
oxbo+0cZPVD4scWd4Gw92SI7HmjOm6ulffOBc4/eqG55gHBXaCi5YteIRY8Ij49B
TfBcGwwcfcz8w49DZ2zloSP57oxlIyilTjdzyIsEx9h1X3wflMud1j8831g+cHrV
PjKFES8BaZGAGqBbSvtlV10TrQzKWitLZriQz84GWqJhhLlSKG2BgiB2ba93zCFO
tlX7J1tgS9WsdP/6uIMwiSkjj7vSwO2dWvb5Ff8I0K8kpxwpazBz90bDLY8RZygh
C9Uzrqv9PihCVTST6V7Yf9cgtcX4LKIttJwD1pF3IE0GPvGNrRjpdhAMlj8JlWnI
wrjjOE8ydek3PQM3JgkpCBDgiD9JKSFgGAUZfQhEGHJhjsmz8fsQA3GchVidv5+Y
4pMn3QxObqRv4yF4euBZllR35mDVI6IeY8/8/n0zTgnWzv5NIfMKEILcuCW3O4//
9ZXQiYFoYe8Cx+SPAQtmJO2pJ0i/IdwiY3eOf2HE8Vmb65NftR7yvnZk9PEzMZqO
Q3qRf5OrmkmymW/OREH9UrMUvXsui3aQOrNtTW+Sq6GPKbz7HAELkC1mN7ubnj9R
FOPx3tMhvy+Z0OmAxvVnd4iVabeiIWT4DgkY6Pbuvblk/jScz4X+15OCT0qWj0DI
30jTTfNfxZU1W3UYA3HS2UHqvvPAun/dqWorEfqulY3frzK7Bvl2Igv9cNXwHtPA
ZUYidD0iMbYsfWELKdPMJD4Z5lHq5GHb1L6t5w7auHyOZwa+3goPpsEGf6y0PVM5
6Q4n1SbfsqEFm7VA9lqlb3L3N7pIP9SqXPUZs4+84BjF1IObeznpx1LnnntdSvQ0
nE307PgjC38H2aqPW/9aUqtoIqJfSuS/FUGjIQhFM+6BkrnJFZu/0xb+X/Iino3j
wH28+EnlYKp2iOrcVwGbAJqtqniIkpu27152PuA6LvOah5tho5i8UYKrS33xATwR
Etqc+dFyLT7k3n58iQ0/m4vgiLrsuAyaASCDfv11+qVcrb+5ouxqtuT//YhhOuiQ
XQqa0lzQBPAr2++xiLd+XkrT3FSJX5ePH2kWDZWr3+WaahOckbOLh0WoR+p8+EAi
Mvzik8fyKXiYdcCjtkL8xRZrfaIA7UvPXLewXLyTFyk3jxlPGVGTp7xa1oKMhS5l
0kARUQ+dcIrQTX0CqMcwWIEWA4MPwY4ZwaLNPu8zLpcOJGbZiVEriiHUDz/vm/70
kbjfgiIBu35A86gFRIBAJXBxPD2Z871PEK3jm1RUBOzhdEza80jLsJ39zgT58P10
4ddqyw4PDq69AES5nQnT2S00KyKBUBjlqLDWhQtGRZAg4t5AmXEq61nf+eueM3eh
4RP7b57XeeIr9F9BCgtzNy021Jmj4IZJPoQz+zUSlYDo8KbdkWOOGed2NMsAROzw
yD0oW9BFvfHgWHV7giyQlHxAgbl/tG3tWo7KnK/MmKPjhqFhf8UVvQY4oWzvKtkb
D3ioYr3HJugBdJIogrffurHMLtdp87JGQWqt0DuL+T5cEBVvXZlciWQvKsR7klqz
jk5xpSKYM6Eun27VaK+3OwrZu+X8U2nGUHDPyNd2/mvCcYKaEmjClwFR+w0wPfvq
cdO5MmkUiUNl6Imge6CVz4i8YSVJCO0Q6w3jECJis4j50v3JGQPI+UrMyvuzpYud
NZPmbtsPINHdYYomp4YfxMun48fLqbkzbyot64Ec92LiW7WL/iOrbuA0WGERPjKU
sNUv7tfIrxmQOtMQS9PofuHGdynKsCBB86IgI8/58meH8hQ4meMVC99I7aoj0ZGz
GI0QPEpHlggrcVCzeVCVxNsKhNyDR8glaEYd6ce2zyCmU79aghcoHDdBG21rUyzW
7JgIlxMSFD+WlfnxjvJonKf7U/2DCvld/JNRke9dU/R4+aZvFKZdHEfIY1X2Vr+h
BTZx+JKkKPJOuzIT314OLXVPidQxTCQGSGzdq575oFfnEY1E6idnuYKoU6tfoD1b
PZFWa9XJYxxK0Kp+FbUZDU3c9oyLi6PweUDHHGt/4jL9cxlLLgHsuaT8nVQPTEjx
ZpJbRzH/GoCtVPcbgLzw3z9pA9A6qxRlapINNfoEKdrvPr6v6FV/UEyTnPaSmnZM
yoqFnnMfufz/HbXfuAyrJhj3OUtQGrAVYhmD3BlHa/10rtXmsBd/FtUOu3tCYJ9u
HT4eNwbrhA81Mp25FAFWnj7YMOtN6F4zrljfQ0bG7yV3RTwuInqqJ3YT1Lt+AmOB
5ZuQHsR4eeRzYnuFeaSbE8QtRWHndjjU69I/aXNPgLUiqL6qO1zrRji1A83ep5zB
sZQAwGFsYCorfqhHUybTRBIuH+6rz9xa3SVDQB9lEwVl3w2YLyjiShq2WJ1b71nK
l1AoOT7ltb1hzvir1RqDKR7HEC1wJbVaFPQiY8BxhrCSgDQmdkEjJknBFyYUfv2C
DqO97jB6ikMUxyOGJKpohFmTch4oE1QswWXIa2urQ8FVHgx4iRajjMOeHAuWZNh+
p6ZhRRgwy+6BPld1ePI+5z+YISGwe1FxyTkrTOPJ6vgcDsX0Q/PQMSyChjUDL51Z
q3pniSkvv423hCY23lZYlYhi4SbexiMfXi6OeWH1uRZCEkMjg2u6Exs22WUsRuzS
nGWeayA4j8Q6TkBVn09vXwomNFyAvkf/Wr3gt2C3tq5bAK+msjQ5liHTcTUVO31d
aK6+gklHPdEHhRkkBlz7+Ss+I92DWQtzlJ+ELf1TxACSuzbfMShWN0f6AVAL5tk/
qHqu16P+tFcqZOCPoTTY7hs6AtZwHGhllIGzZrUN9gP9qoa0Q/hW49nLkPqInBJ+
EY366H4CLHXHRzbv0a0SQag7COLtFcCtGoeWw8OU8WH9mXv+BgfYclzz8RmGnXca
fzKv8RSk6Zvvwz4OTgtqG+PtwKSWumjvCmtFG2A9fkY42VTvfTYev8PXlOXbA9kV
fRvqAzLeLFoOIiXKgv8Aa6mYFmrIRP7rjeumQO7XutrU5CrzKI5DSp2M2QyVWHFx
LwAZthAL93l3JlkEKIOyhOZI4dXHXMrlxEa/L9f764mB4r8lCqww0KSMErYnzKcp
KHgR6JaF9m4gpAeel+afFStbNLuYjxbisj6gPtbmec2xEvTE9w+sXZ5+hoibUQgA
dfZdN8JdwLKCss98yQzYnyKX/g1/tdy6BoXd1/um8kChoe4IC3cY0IURBPOQMNA5
0kjE6cGKx+6S13CHYFvgZSaFyqUFP5suLf1pEnLGem/vS7M/oGrOJHbCvJ0UyZCN
xyTIEzHIXM8zwpV3xA8Gj2/RpYQJnGPXeo4NxcKGU4yvfNIiBI/vE8f6j7QbPay+
/aUMnTpeTA7YGMrwTin5IBy2gcF76R/5UY03/u8e4GrhCQJGAg3MEfyHdjGODvYB
xDsKMv+e9a2SO0Ekvn6KjUpHQjn2lq5peWHJt2ON8UguXL+yAHR6AmUZNypPQ8Qc
EM+uSYoCov7xSybaehQzB/v+GK3uEqLoJKKXcWhsGDbikl32agkSx+PLJ+meVyVO
/7DqGrPuga8mSmhlZoZ5WMCKTU8OYRrpXk1s0cb3Zg0Ba8D49L5xlY4BITpmaXjQ
gkchzwE6+p8JQ5l3ULwwn6q8/mwK1qUB3VnbBOjpON/Zi+Wp0eHBlJ6mhvj/ibwl
CZ9dLibhkPG4Ttsbv2CjY6dO1OxuXQJEcyezPklxgVoz5u6d79T4mc5HPtYPC+Tt
RbTiv7CJUvx2TsrsLZp1+yf4kSAyjt4y7FDrcuRBHAcwBR8/Ep2ZGlw6fjil0jBa
n8U/e2SUtoZfltMKMG4t1Evi30IQdpHdZ7kUu8wVKWegOmots30DzNUA8hKz92Qq
1LPfbQIe1lL55jwExXT+SPd540bE4anLmuEANPdG/2eYBBYnOO8SsegKtJ4/OSyX
XiAnQ4qX19930IpnD3QsmJxgM9VtqMXn1i00hVDb4/7FREhXHjSPcvdwqk1itnf0
nBNAmdETxFscOZmJGkYrWr/zl0cR1DV6KiQe3loycszZS4F9PB/uVfVeNLe2ld3g
Ncx1tlZhv5g7ERqInXX4HFkYNU80jxdLpaNACEVWaxdd4PUaMRIGaRaLNEZNbMhh
RgOifOTPiV06DY7/V4ennIhwoRocJLh9XILp9TAbe4msdlelI6AjjcXb4iDxCtcP
NeAN9Vk3tj1ae7IdNm0sXULkgHNkZ15UrRb4RqxbREZUxY7IGtYaho4+NyEepJAB
f2YqeMC0e9yBUg3QE3mxblIFmyV07JcfS39HZhTNkv+61QwbL3NptcE4AHhuanwt
hKHcKAqXZ/DNq5TQ80vdRt3wogZydyb5xlAqppUVv4d5kCgVaDX53y9OfdJxHVk4
OJ5B6zZ5g5lmgOUJNrrJCF+uAeCTlJ0/gdwR9Ali6gP+k9RPuzpMxr3Xjtq/CFzp
477LzcDBNslaxhdKEb5fVequHldEWcEHyC8sw3EF/IzM5zWBFaWUfzDSgug701e1
Jvmz8Ms9PR6bFJiI2kpgTnF+wb9wR0agdPlHVp925imMScLG/F+80UorZrFn624b
8socwIK9lH0Ij4AIl6q1IAvqM6Fv5m7nt3XqIjl9khlU8fydpjwnAgPJB3UGR7O1
D1LbrbGRD5DDb8qETiW6v3zfvsndFIdlXe9k1f0e+wA3eq2QY2cuLJYduN+1wGuY
H8pawHN6xjQVsUPLpg8jY/ig6Km4CY7HHwOt+epwkfbkXarIe2RGU7XLo5z8oNS1
yZcb+8DKQb4/OQ6RX9JYYBLdFmjInK+6FcZmgOzD2Jjq5DRjDG/kFZ5/N1tx8/sg
7cgJWFNDtizOIrVL8Kc2hdbXagYHluejI92rnHf3WHvlDlFt2aro20WRsZF8kCJX
TnCTpNZhFw2ezS0ymsWqy6pLDQ3uWg6gaqPhaDe9SXR9jR8e2ZKqm9aSLG1BQhhe
rbNBHI66Bz3f0ycQomwd5CFI+V/C25qD6UBEz1BZb2o1B+AHTWoSMYnpfZfeP4M6
Jw/c3JxtOo7ZCOD7Y7DKFEAZTxpqYtrjDU++AAeBz8uYRSZDHRFxtYyX7qB819P9
x5avfIJPwsYx+GckzzFK84U4Lbcx9HnzQZKIvUBR5nDytnsGEZLFvuqb+o4oxBbD
CCrVPPNChVBs/OyxiIEfmoiqDFxvnxaOLIjn7M0oGyrDtexb6PQaFmL22C3dlqdn
CqKd5QYqasK31U6aA1Cv16noKrdmyzESNF6ThMICCu8QQCsZrbQFgC2zbgYL/bVO
E3cmbXZzLPcHuEAymxZwkvmdc2p20m2e2asVOfftbSR49tshNi3rRg6oyjM4owz8
B8IJmAs6lD+ULE9cf5JBTjlMiGqV+PCByK1nKoyXMM9W8V9GQeYNfUF/ZWjZvrfo
3gf9FNpmm3S9hwz2ROEV3svjdrvYzQ1BxmkMoius5aGDGvtQorTtuTMHgkRAI2Qc
mYteitorNAkuglb8KuSPYyCgMfBqJLusX4V+FGp9DvXNckyxBOeD5jEGBY1rO0Be
VM3BzfMPw+UlrXx0b1+At/v7qNbe50KZhQ5ccOT+Z/73X01DdWdnqIlUCeTspVOw
JA23wXvP2k56RCWGtysnTOQCeMBVC2S9XHcwDgJ6V2/RNV9z68eeVO3kHChWxDIH
tpK+JOnLUfrK6JOej7R0YsMugFJaByCEnzMG01LiYnqd+xJ1LowC9p22uurLmHbJ
mZ8Fez4QPowSjED2WR3f4I2adC7361vOYOflBWM12Lfqrxx8/zlEpajva2xiOzcM
Qs1quUF2JWOuU86XGo1pd8AwjYfTe1Kg/3+l0EieSO7QNKCR+imzDmz0SQa9OCzp
W28aNI2REHyMhLnt1KGTaB9WZTf9KQseeGOLDdWGSHKdncAD50vI9y/VEpPXc39E
CUKMK5UdSXwC1h+0y4L92/1LcqM/ZYzPa2QohTGt8bLcEJIIuo6AYxHBywb3bpHP
+UkAWADVMDHhLTvAwvK+Nsgm+63y32ssKDufQHnEucGEM9eZlG80XfAuzHkVCldO
GdM8KAnFIIbe5gcr3RDwtJOsefmvXJMyAalErl+Gghm/No634972lJG39fD0k3B0
iESE4GCVwRAJn+BK3yCaLEfzu2iIilQZGOsZaBEBlroJ3pL+l+np5dSLISzU0KLH
DZkegcRFDCD9qmYHFgKDqgq8i2IKyTuI6xudXwvfmYllG7kLyfvfSSxuLYwn3HM+
a4CD/S2m2+vIpUGLzBGBNLV50mBb/9YgC/EvyWwr8sk2OEbKHfQdOjjEiowCpEmZ
IUXXViOKMb4FRYcBU46/vzFddc9mL4iF/ej/HUsL59rGw9lnqa0gZZqQcxf+gA3q
DJOo2sEH0MhS9WBj833u4Dp+NPrBVbmAtPTYKMkCR9JpabxRjp1OV+8Ej2pExKZR
yhyw+8skqyH3ANMji9BxICGiO42U3C4a3Ewel23HWw5gDe5en/ntRjA99hvKEPJE
NBxSerJSMxbuGNOuFVZvIw+FvJ/vv8BS3SWw4mhygY8OrYpe0zP9tap/fZhwwM8e
2elvGtFNEaDgX7LxpAvpGhneEWCk84D03DQMQ/hDddWtvCSQg+AWdcxFL4v5LqHm
eS2WN1Y3b+64rw5+6LhlhPeg8gBGXBmhZkjseWxmIhS0toisDNbrltiJZOmXyYM4
TjDeN6iW2OGwhqAApDP5rrmWYyiQgzKhAVrzki7gNnc8Aj5vDidUYvIc1ovc3Maw
hD02eYozdzDMeHDEoA/YD+N2gbIolFzlCh0ulqVcVpWYF4tVABUZXoyzM1YMXkxf
9q4sLzokPZwQo++38GkGBdqCg69te6vYuWAAK5H0alnuU0tdmuNd12MctM1OClEV
9idavaQ2o3CYK26R972N8z24j3XXttDGu3LuchFToKDwReGZOzQ2dhaDsDfwJ6wM
N+ltqJEonGLlzkFjUmFxoF0cZ0SKbQ5VGpuyr7ViTWC/CLOi2YK1YLJmY4zzyYZ3
iNGvnGQu9OwVYrHtuzRqV+adCXkBQ0JVuUxzsuyToDkaNJ80ORFXGxuy64A67R0J
X06fbU/Spp1sJ59Na5HikK9PoQDt3qME/2/kZ9a0PuM+j65cJaI7NaZvvOH8Jwt3
FkD5O8PRRfojANj6NHfcmsrL3wdZIHcz+ONR+wCnaXA4SfTHcxM579PraRimFv8T
06tMbfsn4UgAYud20dZ5Xta531lSMCqFrZvTyzrNYOIHCD2MyyLb2rHhcI3ydbIt
iuaqXg0avGw26xZp9E0By7/wfnlj2CnKPZGPrcd8UwPRkuGe/bqPO9H/f8ZfDKC4
e+PhviiZjuW78CDyAXre+OR3orZkH5MwbN3ekzqp+NtSnHnNhk3LNATM64CLjYbl
n8NeDWdglD5sTqLFZ4o2VCFrZgfMK+lSPodCBPmJCCfldiQWtFfJHfnggrdXXLJu
A/MkmBUzyCe4p14LyA28Fbame1Z2sy3NWUls8OvZ0quTt1/DzpDcBF64NOajmCvj
vTd059+Aq+Ez9SRoVZ7k+ovZ0VfEEVTKFKDXTsh8xpjECdFwN3HTezHP8ghD1zSt
axoWhQJwn9afdfFVRoPr+Yz4w6ssui/PVCXOQWkLX4m5crE5kdjM85jfzlCcp3/v
BVgZ8w24IQgJU7JQdzqTeFyr7GMEBNKz0+gbPvAdCva//EpnwIUh9jBevYqt/J+q
3CsgCxwl+cOSF0q7g++PxJN/sQg7HwrsuXj4DxOtZoDK12mPCA9IfGt9JbyY/wS2
25MxkQoEF9uByEoXWHanKrR/K33D5wsA0FL+ExeW6l5C1rxg3ZbhdW1m/0/O9VgL
75mOdPliLdGLDE0RTcQfuv/9i0e2JmGVHSZ5pozlAXHkTTMPZvJKt/USgiQi7Lsk
KY0/4Zyi1dhvs60vbeom1M2J7MSgtcSYAcdy7/ibNTzXCOvPt6d/q0QDw4Z4yU/H
leUv73i1vNm1lsiGV7FEjvJCW4M7QYtcdhUMNcG+r0+CwUEXGaB6RsnfXJvncgOd
PRmQJZKR/ZnRcuF4deUKEUQMeVA5cNJKXGevSgUUtsXRqSAQsG9lzQbPpVYATmLg
9MiWV9FElqDL9Tb5gpp71cfUnyCmbasvXb4NHYyyazqVR5U6p30ejUNXWvGucj16
iv+WEj4tvhL6PDsb1r7M6M4IQxg4AZBYmxsUVUreH7/q0bLw/J2L+AEtcilQTfbP
HREh2ggRAIhDTASdK9iDPu2h49uijPe+bSXUgpr/fkhN9gwNPAlBNIZaDoWkhSXb
fGP7BabNlqIC6EIW0r4j8bO5Fw7/Ur5xTcG/9c3zWkaGLLve3rBX5M660bf1bwL8
da03jpbBhT3/fgyKEakgyQl5Zsq9aVdYlpJNXva2RoJYfh7fKId6d4S6UiD6Nbz2
sK2+6ma62wmWx17Akag5r3LT69W/9HLMUAEl1gOqB6kDqzJyZpjoLmV0u9vzQ2hv
wwo+cjXVruPN5cp0Bk43aoEl/vDXeVqtgtDlHwc3tW4uYtV2GQxrmRUtD8csTYIm
vHzO9xK2YtAcITCuI+obl+nlV7uuhgHbTliHTF56vH4BebN6/prte9lkiE9Px/hf
Sz6pEaiazlQuMz5CPF400WyRcvNLMnXkDjnrlRPWFgy5GYLyIwEK3nE0QD69SBFw
hlYWiL+1gFeZ4VJY6vL7lZdcxiknKKYIZEgK/VfiFNEZskMRT1G8DAEt6FlHh70b
MDt6mGjFjCZlGDJFLo+Ar2Z/StfqLWtmRh6SC+8MYeCsZxP53PAXS1Jk2wz02tAD
yGkn45NyWETpruOJj79p2IVmgAOFyT7BbQL2+3GCFfS9b5Z530dK/yf0YD9zYBvg
mjSjhU3ipQW4Q9+GNK4tiQCiUXXUAWod5R8drW3AKknn4PCHlgTZ7WOOFnIcUVF6
oFsWvFsCMZ9YbtWett3wRH0oWNewGHTFIWxgvmrVj48WedUjjR0UtR7viRA0ofa9
fbaPNVAYy22Rbzy+yalbvFemMcs0Pj8oD9d4AK7s9uJXRzos1nyA5ukV1O/WIqUu
QMrXqHOiZ7EL+aL4SKE2jI8Wi6Nm40l3Z/CLGE/N7gIGeOWbzNATTgbZ739JBDKT
6pwtabd/vd6pFaylNTAvvM/1Py91IW0AvfiheBialofR1fYf+E29X42EUIxLCEsg
cwbVwIpKAAHEfAsSgwz5KpMZs1gmJ/oMphMXiWuicHOSFWYZ/heICQ0arvnHj0y1
INDgI1crNUFV+xwMug7dqSGd2Pv4CKcgqJ07/noMhl5T6zvJRZpMLycA82j7jNvD
SMEGFjWXOAZPz0Un5knNs2vYr5UbTh1MUCKZOn4N4vlbsi9oJjKIUDW8qjULPQWu
yY++z9Dw0gpOdQxkTpIaW9O784w5SPw2AwevzuLBCGJqcoDnTQvwdcCxP32+tsDU
I1UP+GUPX+AknPOcMN8o9WmFrFDC9lnkOAxMkKfIrTP1VPPA6RRJmzJgNlY8GEO8
ixYtZB3vXMB/RAAATBEEwi1roEPmmbVdZD4yK1j9Mc0AfTDS71wKc7uNmCBpeyXC
vXaOvIAsIH4QeUBOhhf0Nd9r48Mp5PiXinta8UZyNEeI6unX56UPtaGT+xtWwZs+
xhvpMidZCBOlt1hSYcL3vSBrwElaKyyBsaSjeLvMrYQXQ3hPJledSlwM/m+9V3dr
9B/vxxVAO+Vb9czRgQP0kcSenlx0UWb1BZyCFA+lgbB29g5gu1tFYt7YdUHbRW+I
+xl3L+O9PawZbE/OH6/N2YuN6ksBAmWDkrPzrM4zC+Wr2X/vk6MwtBysAxGJtt6M
XkojFNy2ZKvVKvqSlpJjheSVEjSvoeSghm/gmmndshLKyGLf3FAjfOe1qtVdTV9x
Hb+aYqBamfimr6FGV15NhtlhPoPGmtU0eM2m09F01/BGucchtrM2cg4IheDKfVZq
nN4AhCfabuwoWZ4+ahF9fSzY0aFb9WFJLzZbEc/I2MTpEZtA/VIHxkXZLxsnM2il
HeZNKWeJXDKyhrScBkSmZHFtHo5aiToXzFGGoN+RPJHBQp0aumxdJXm46n661w/f
0+w5etFI3VfUWGX/7PYkHL80JYrU4zO1LrXFBej5go5QR84yCCusjld8VY+JZ4Vh
z9l5yIptnXl2fPWUSfVh2iWqjTIWlwwz16qBoNUPMI+6iBoAXfkm/qqSUaNIKB9o
PFuWyfEluyrqlMVU9VYVpi7kozTIknAtRL2h1OopPHW9dA2o4bGbm3rFC5XJcr1Y
pHYGDToGKdpK0JGe6X3lW6iaQuLttq/hJCl1fkZRveo+dtF65/IvFHVn2V8ty/pl
vDLNy4uuaEcQoqQCVg041VCl3wV0+zBYpAKiBM9WsizkSPolFTD97aEWGMRL/RsW
YsHux69cLZ87Vb9QdABtv/YLcKGR/UEJPG9c3leOxpeL6Nl/UTQsgakOh3fGF0Nl
NfVCYUZd3ZQcRoXjvgjjMd0gY1tGhwWPlrp6SI9BgzPVcN2AmlnCvDEK+bwRQ2gi
WBBIXT6cJli4MvbmJYaguIWhyL9ftZJNYIpBSaabCsWXzFU8xy2bkR1noHDoTO3m
iJBWYTVMs7eAWOr2ebQkbDO0ZmUFyRH5Cw/btroa6nfLur6vF9AqThJsS6tLg9wB
n6B6pOxQxOP5Ph9be9yXdmgyd7g395+OJWB8uIZp5RDnBLUzSHqUXH0ZEf86pF03
l3FAnDb6BsCYLGRqqHNovb65qfzkUuVkOY+GgIoyVpiTHUINMd1e3DjPsAj+kIHT
TzjG8rj0O2ZCIyMykJbCma1rOfD78qNAi8upNIJmyX8W689MGpSgaX7i/6ne89VA
YFrFeS+Dk4xK853oufVrZ9hJxysqgTZIm/LAB4tElgjX95H9t2wCe4g8Yb6ncIta
rC4zqSHNnQ+2S98P1V3LzXrNhutQ88a5MhI21vhezP+TB+CJaeyBVUmC7ohcRI2U
6iyWb2XS15gfMx3XyovrKiGF3w4MqZzTB1FamWBJWwZqCeHNViF7vciHOeXKNRnk
P1Nl3g/oS5E5II6+50Wi9kiHJek23SuF0V+o6lXBtDVYS2qcTVfz9lFEhljMhNeI
9i8XnSVHFrcgxqPk7m8ntBfBYNiMaqGP+YMneP5nFV+z3cCNMSoJs/ET1x3iPA1u
QpqleiO7A7r64qZkGNt/f1+j3I3MzG7osE5mJtcKeVF3TA3ZCSbFompdS+agBpnv
A4ptvttA5Thts+DwQdD15U2kevAL1QM4X2BnvGy7D3iJ/vJvUx4mXlHoGMmnLwJk
IjXvi63xrNLI6ubNvBOJ1qPriR1A1NOFS1jITDEoLfE0wypXWCyUkdMVKQhOHVE1
RXNjizZphPXTMyr/aCAdAze0G0cD+8/ZpLUIRY/y9SzrnBg0vxhJBJJEOHfGrqrD
qH4k0ZHugtpZLNt2bFH5wFMzvb4stAfVZwJazzERxjDb3E/OnDtAKtjDeOboslo0
kCdAaWwIQ7Te4LkJxgk0E+NdLfQc66RSqUJ1Ed3byHA+fu+lxUUBTVbXpoI19BX2
aI9+Pxwh+lBWE3VK2XgjXUukyohIJ4qq/4tXfUI8Ge/KbCJ3hZu9IDK1i+KqvcOi
0Qj7u3b1/rpY09EHdCgAmbEu8ZgHKUE03RPJfKMZcXG5L+HB9/6w055EezurtH3l
FYqkcpQd2ljG5JKvnnfErfAHJC/ZqXCv0k0bZaeVGUWl+78qM3iB772JkFZ23tS6
+9hFJDWuNMs+0cxb+wdHRgYs7OebHvHIF7OxOPlsHSG6dKnEicjjQuqncn1BzFFy
ExeoydV3KO19MVD2pB3Rju4tJO9lyENarckGPWth5pRHkZtqhXizJcD9xAHPtdG+
9IghjYdI7jIqCV6NSI8IDZJMgPFP4kd4G5SgSC4qRuv3xR9EKC1bhyNAIyR+Gktn
eWdn5TM4n1MkRl8IHjAXL6kl7SiDX609ixzGPgt676fifGEiJKkbKFMpW94WQvq7
tPy2WeIrUuVpDUYBMFpd63830npGzlpIjPGUkzwM8i6PsEbXxKRhPSMv6uzHYCI3
uYrJaOVbJ52YLQmsY4fvubIdysqGbJ0XjfmNlZ0xns0mwHl5ThlDCCHtX6wZylg5
CYa+I4jypr92y9HcJ15dGVfDofYZUFd13JQsAZLWtnEn5+65C6VgD9q8dALO4lXj
AZsG0XKFfdUK8W3vKsskFk3GQ2um3BNnDJf6aOmpWzyLjEc3gibPtS9IAm90/9mY
xlcFifdnPiEk5o2CrtqXvPtWAQq0oOq5TnessBkGoFZ9kByE2ZttZ3NwteFMAbYr
zUeC7AmtIE/cMJOsR5/Dl80twrU/CUNi4H/uD65jidr9mANfjCn38Lt2rXUXpgIs
/xX/0T+T+dPC6O9xQ8ChCZkdYL/ugbZW4/3GjbpiH5AVv0pzvir1Qr8xcNoX+mJL
9echckZ16LOtGyt/T9xjK1nkzcEOPKX2jKd+JrtZLc+7Ht/ks/9wHCoJCB3Dc6by
AcvF2yHPoh/OleZ63nBuOfhgQuVRPBLJU/7GJRCB4OILih1MRnzKQ94/qxKeFfzC
w/+Kokp/9OdgihdNC8U4y89SFk6uavFfKaX/3iSiYm5FILImbmMibDZs6LmV7Y3v
tPh88EeD48WYOj249fGR81ZctXe40zlFU7inbhN/DFm6mvYQ9CLrogsAnggVISiA
sl1yPy4dmJ0mCW4R86+r73KQaqn1P9iMTpWwtpaAwWBnAzQmlhFnaadhjH3l31Th
Q0yFZO6i+o9FZyQX9r/o7qVM/jq/b9Vb8MkJeZQTQPXt+dEv06XBCdOXSUflnNkf
nWFlbI8IhRtBHxMBeEwQ6cHwW3q5x4yM/fhKbFdWnJzekPK7O5NA5eT4Zr9DEVat
DAedKRGSJvkud1wKP7M4K6I4+UQdhUqrmtxdAYXW6XoiWzStNV+1luZ4AcPUQvhA
eX5Pps0y471q8PHiuYygBOQELL/w0y0YbG6onrPWTfKULByIpWjXeVp2zlykLYFv
WPDu9y8Jpu3qQn4HYOXQFe71IhKp69uZ/U/TK0BVrq8vaPA67uRpFnEzv71nsYGl
Q/PW3n9Lo2vLIcixaRnx5QcMSkb0+srG0i+YFkV0CKGbrWitVGx3Hu2AzRpFEbcy
T92r+r9mZLOQL6bvU9Jr2s5heDS+cDs799GpG4NxfHgUOfGNABevQQzCYNNIbjTj
Vb4CIBI3v4gqH2Zo8/suGZrr/EUS4wEU5L+D9d7Z0Jd9UJ+do/KFAPX57POAkhYL
Zx++Sn7U2x3jjo0SblZeJ43TzDrkrD4kRGAFWeGurdpmwox5ujVwvD63jikaw5q+
gzPrvvHc4LiVIYkh+k3uo5g1+urvjd4YhoEzv9FBoIfMbPCTdYV/6lizXmuhnYuM
mnWBDrVGx4MVy4Ny3AbQ9/XrlDVAtjkXtLZdvjuCmWSTr9MZ2lGIygEHnk32TDsU
/5Kt4bOAVIM1kvbk7VdVy6QawF80OV97pap328eOo/v9pzDl0qSdX0U89wrx1Umb
faFGlcyGepBVG/zIX441/Ml9K8C0Cxut5TVloNHkZuLeUflvBuuMKDKtNydzN7RI
jC0/u2+LGN9H8uRfELSreOyKv13YYiKj/VvvV4WIM5lXeNZe8xGNkCohpx4f+VO9
82f2wSkrhIH68QWcduPLaKPlMsOUjKNdeD6UVNyltv+MCknTOFnBD8T3Kmi7Dbk/
N+wO/jJjWRW3foDxY2Gk2hFdyk1hEIPLhMpJI6tTE+jPBLAal4qcinpdrLAJFSXZ
ngn2k4sv0Q52SDpXH4PfuoPk0YDgp1twbd5kpkE5jlkQQo3MjlMZ36CEJmLFwDO5
kjbmP4r3mSlTX9Ff6Ne1MA1B4iw3JXaE9L39Qz4mStKOkB6KcXhlaU1BC3/NSiyb
lzugh460ASDyu5eA4kuEfaTPNFPS+Kp7OMydG70k14edeHpEcooHIPlHMewkRw4h
ZhZHsurtQiIXmxP8sZ8Sb0vkIjbcKGXMA+VclHWB0pu4QGIxFS2HJoDosZsggBe1
15XYp59UbeCjqznaPE/GszTner5g7JCqLSoEkWogUvvLZUPSLdO0qLh6jvWSbu1J
EiidUPYM7XtB9Vw5RrxkU9ZXnUMDLunkSEyeeUn7Yawn+jCxVYVhy1Fjb3vCMGuP
rQjtfOZMgbnUemCpOxUSkrU4paZkKiA2M5D+4WkIOkz4FFuf5DZvDQCqto/Nj3jZ
/GyNXAhGGoz7Ldo80iUeojOqGAVP129zDOcut6QJcd2BPM2bEtSofKEiv7OSzg31
pjgmz8IvaEbtQkRrKzd8E+syFjQe+amqvIwSk25WGt1jcNBIUZl2ONX0f7UWEDmN
Jq2+8KS33ON5VTFt0cF+XeduIdJbcaQl1BbJQG4HK8/I2qUestOQV/lDI0KuGN8w
ipYBwchkZY4pgTZjsphpENzdOW+njZl4m1D0YIP1mcOf+VJY5zM3v0neyW49T7TM
eed0VlFFCweu7U2C7fnhU5GI/kaW55yqiBCowpjM8MZ9zEhduF95Fam+CxtW29XR
zxq413MBh5MgvtUopTuB9y91+W+6UEbROYtm+ahgb5mjSu7j72ncQpivoCZy2eLy
4LEUhms1JyN6e2+Cui9eX4YVNHz29iZZDCQy3NNEuoARd3n5BkFp7gBuW4Ua/7aQ
K6YaM8E3dMuRLOUdcNVDEickF9RnOD99CQCi4sQDbdErEr19DyPqInOeLjYYBAPI
JCbZPM9CS258OM6fOnXMq8lbzpHKfrO4VaQciaOjbBRBvX7RKFbZ4DUE4ffdxXGm
Dwpo1Nya/zzTlcpJF9nwSxa+bPyMIqR1aJ8eQAfrp9nLNU4sy3/Pq9m/SLLU8ptX
7Bf1CDS6uejg9FS9EbUzxqD42coK2n3rBsL8FjBXvN4mJWYvr5g7mhae2uhEBdBg
XyF+gx3OmC459TVvNYtJY8RqZBi2lrxs1cA3/IuQ063ZkDTFjxe6/0diOEV1z7D7
5jBZv3q8fA2rd2EesRX7pN6tZpShM6OkxRltCixBU6taSjDVBUiH3DNtE37PjuHS
BE6tZECr7tTy8MsIVDzWpvXYmXMwiCwF4x5kWKM95Hf6VZ+yWYAYAwYLeS6LXQLv
3nUa7h/sdu93El3TSELw+ncH+A0m63NCSzRI9HkJ/HiZzLWSaJxbJbPvdlFwjpip
IpnaCR5uuffNd2axzkaRlo5sdAMKURRhS9/N95eekGe7Koufa/KfF1LXtccfU1TF
rxuX1iozzi4PmxTFMCcAV4ZZiIufv7fV+66vN7h8ezJuDHmfx3D5LwH7WW3NJwcU
e9B3LTTmNdVTQdQyGprr8Qz/OmwRIWbGtZ2ypG/0rfe0s1hTozAx4JDdLBIgCMer
A5DNBKbWIQ2Pw0VKuBo+s7B7U/9c5Fj9x9cOuhM0ixJzAtyrMeqEMSGOxKl//PHc
QCOdHsXwyaX0YFIunUTg6ARYDZQy2PR2OiFQAuRPUXc+JYIM4I1B0WMRFzEqMs/u
QDi8y/4mog8WQn3fjSBczgV8r+oq0dDyD0UONC6GJbGmpLnsDR75Pqqjbde+LzLF
tXnuDLavjJGVMC0XssD8zK0Y80uMAY3FzVv7UXTuxkELvoRfCPKMfEO/cd5GbPTU
K+W1uiLhSFCx16GbYOzgJiqdw1c6rnCshzR6k+2Z/N4wMtI72b5hlYFjK0jYUfoW
Inq6t89j6anNHu4DXDIn6nTU7IMpSIVRK+rVbCjzWyciILjDI6E/vRPL29cwy7jN
y3uyQpnx2BMMU+FLcTSuScXRzA0CFu7CyN0Z+4LAc82OO57qHcBfADQz3uYSO/B5
atE09EvsP7yd7NmBJaS8a0yU5cuMYXQu6y/TSjKF/6wQptffAh9qLIQU7O1qiiW+
LLGrUccVKJAgOzMO1kfFMPj4R/DycHjlvbqcdkXWGvT0sfcJD8A8mFYD5Mv0Q2hw
ElU4HW69q3EDinBCIRqgBpVsV2JRG0+6ELeXUWBRIqyv6NXP2C84i26rn9EcLg86
SQnhDcues1r1PrsxTfR3q2HsZjrk+pxMvBeuZNR5BvgKMc5z9fm+k9jMvlP+ulML
fBGK+qR19J1W+KUdFbVytfzEFBZSisFP+mL4ZQ7pBEtGTLwLKAuXgNII74pztoDD
IcV4nAPzulRBlRpgCClC+Baw2YiWZNw2696weCh1ORTCrgek1U+c2AzSUtv2Zme3
3xvyB2sTKCHZEHcU8pLinuJREU4wzO/fJUkpHTHuJzyFdlOZSrKj6mO7ZvUzoSNl
6fFO1fBB4ob08wCDy9iCVfDI/u+FCQn0cYp60r+8oNHPpIR0GwX/QMjJNuZKRLHH
1yi5k2HG6bZ4zoLCUAInQrGxcPjtCgZ1VGsxffg28yPNktlKvf7fbC2wGXPCUMtl
8ID0Qi7MHlbWf69SGObShmwLqOA6HVu89knfMWwpnSPxJh0FGw7YcSC0Tsz01lbc
ziIByAJtesp1s9bZrUkVtbdN7fwWeVpk5ADlc1iwQn+OY1yFFKNRmo/+BDqfB90H
rrL2yCBB1ch+Lx4M9F8U4W2XEHqzsP03pMmfoGNQBRmk8HPdpJ1Hhk3XU4dGcr81
YdYS9Y/KTd8w12aKVNTWCCoQcdhotAbw+odORwMvUriU+3616/dTOY8Uh3P9duV9
NX3waL34S4ZSHoUb5x3OOCHstwvdxaTb1v3hjeCbd8HcjTcrTWda+wF9UhCIt09n
Rcso/BvcHyTqyI1VWQ4Uz94v8Zs6KwxEeBKLpIxroXFfbrgGesXf4Cek1JEGh/ft
AHAuHxprPVt9cBOGOf44FtnOwPZw1LTW9PowqRgSfsmfZIxqZ3zLJ8gPSJpOnTTl
Ep6+jfejM/NIoheY5arQgeLQbnP3E9MfwDUGaZLPFkzXS3Ay2t2551iU5PqcT9/q
OsWoxPIHU//MfQKVAtJHynpOaLBFGhyqqSqDbF70m2yWc+SCd6eILXgj3OerErEa
eN/nR+1X25DpIUjyJ5BHEg5fgS+IWfa0lkKGDeiJiSzU9x5GiE04ovUwBBXfHw3I
LWZGSxO+Xj9xWJU/0oFBIp5nmfVJSI+KZIcX6DfInjdwLUDjKHvsLp7yvQx9yWoj
8FdYvb5+4/7l0xoMSl9W+E+NANHlreD/lidMubHpq2HaeIrUIE/cLNDTohogAQMC
HP1OgLhhOqdp+CHgbIsu59gu+ae6WZ79XmcxIDHMWOc/UW/YvMcg4ihaAtOHwzbv
ukyZihCaz3/z6vBU3DWe1+tCp1PlBdBk0BhUu+M+m8DKU4a8hKg6oxQwMPImZWtL
MYZH4eeiDiKFFjQFpD6ntOB7d7iSoS88y7MeFVReeheMYkZhn2nE+l/thl+Rb/Lf
X/0SkfF2n72Yh1aMOUmpgdMVbB4slrCeL7lE/nI88sHb+/g841m56+6BUlbcTas3
KM0ME1I/XzOXq4sh3GD2GBH9B5gtUiHRluph5OGBjGWV64dhbQ6Vv9P/4H25To0/
diMyeb9nGwj+tAYm4DI6uBaNV0lMhYvKR9bXzvqpasER/wbQplvuugTGOXXhqsDI
FQ+y417RELEvYCQc2LVtHs4PIZSTX3ASNHfLSBdmIOCvrPNf7rgvOXmjvye03G2C
ouxph4DMjIgd9+qCPEuJcFEHgM9AWmRKafO4iMPiunx0FE9NbrSYIsLUpxA22uiw
yGymJNkMaRcwMdDnYlxOGUVuRTm/su5HgDPuYWBk8GG5AgZCwPKd0Vz7PDShPsFz
hGZEITykwMuqYLK8RYret/KCpHBSZT+bpb1nVARL7WNVazdizAbnM5/bILaXNZfq
tBQ/HXMW1zo0GhgLxCeeK6NmfbmQzG9U1axd84hYVcYrEZrsVu0tVSWz1g1q7ubs
bkBlWHFLDZ9uoTob8/ukQzixlb/wI9RwgNlTlqbke6/glp3QQv5LFNSovgFcaM6j
XGiT9iHjEjbqFItqcs77yGeWuln2tVtIjYV/A+59/TGNuSCWjjhxNRnzDoTW3dt3
1ZPKAfwQ9Tl6bRrbC9LcV1Kk3gVh5qGH6WEiB5d0MSDVyMCOkE+OzZH1OkInVQkH
2w4S9VCboq5CLjJc2qRLRQDoSCsn+14yMfyRW2+oGYztzY0n3SNm70zW3mNYGQHN
sDRZxp4fqJcvyx3KAHJnRwsP7PtTijdC39kf7hs/OJvy4KKa7r5o39AvHpDpiTAW
u4eLEAoevtQIGq/9ABZWWEQ5J1nYl7iMrfZDPXbn1lJdvUoH3t9xne+5bzA0/9bx
F/mv0sRrhPurWXbxsX/79aK851YT01w0yhtc6dLGzIWOnH3UdZYDnw8KXFUA5tlc
uhx/KuxVZon6VPsWwBRhdnKefxeAeDH71F66JeQYxhW+xoND5jd0a+yVWfQATKGx
IaGJLuloDXSNf3j8s2mWdXH8n+dq19jtiGEzeCXgMXG3J/djk3pjlIe3RVw6xm8d
9deEuFOlMyrnD7HR2O528Rqj5VzYMacoPiTxYcahrffVU+FdtR1Ex8P6dhuR1EQ8
cWJ20hx7bhtoXQXLBdlBM/VZxBckYTL5tOZgZqRwt9Apf8Ch7BvPNB5sKDO/czmJ
eZU1DRJdPbN/uRuQVChzqJ0TV+LV43GbptRHVDJ/AoL/7tPtva+aSrq+x48iv4AJ
KPa2BoCGEPVeSXOyYZyi0GY8zGb2sWxoG7Rjl4uepRH8wJo/Fs2p2VL/h//qci6F
uppX41kqWemvdJzKVS0DBHGAvRrZcDgpEPz9AuUXJDwRWOG+P5tqD1yBfIQ2zmO8
T0W/h2IDujousz2HNWW/trQDOnqx5yUhCAbF022P+esGOibbpClOiQwTWDTEv0UN
625z3yuloGF5rT8PPy+zuZK1EKHFDH7G2ZWMSvjVOtLIdnM6Ft1PPGL34YmoIzHD
b2G1YbtvqG7DOCdauxTTErzkPJLNvugfVX/6xc13vA7phPBV21AyNAfADQ3iVmej
+kt01w2WpK/V+eeuEJAQZf62125Z18EmpxZWZ9NK2wplrQZ0RxVFwzZdlZLV8OFx
BiYPQ3PU97g6DqDJaEyIQSxp+MpN0ASD4z4EzKwGbczKPo/54zrh1zMSpg4U8KSA
TVP0tjfVaRpIGHsZbC1u0T53Xa8qbYPuZg32xrDkoRa0RIGmVATBdGpCGef2xtBo
YkgCMBwpBtLmNIZHXGXMU5G23knh6D2d0+3creP7afNk4ZG2OteDVbLUCQxJftOG
KODvWSQxYWOB5eD/aDmpjcInPdBxyvugq1Mh7cCvvxFse23aWMVrEPzvts8z4vkL
b9SXZjAMJMiUGQ7PA7/gKks8+hBYvtnhlMkppu2fnaOmFp1wyxL/XDlIjwblNnKM
41Gs0AY7UzkiBK/75U2d+43r7ruNrva3li7i3Jo1/yqb/JcpJZvaXcNJuvLyyfrE
g6wAoXOiWbhQZNH3ZcTom1raxFws4+fiiJIQm0NNY0VvcUcvA5p9ggD3mAoee++H
y/e10hgjin0EN3lh1JxFT7OqZFh8Jt0cuCdWT6S7U+Y/7kixc3XK/B0yJbV5J7Ed
qQOZgJ9gceBeRVVfm0xRg3I4FoRp1GaA2T77Pl1mcropsUJ/Gt0ZmNXFQvl9EST/
ddVQ1umqBC5t4W72IpDCr5V91ytS9YB6Yaypj40subPTSYqmyvtCBBxglFpwWZpS
U7PQ8m/sOfngW1VZ8ShCk4Cvq7mepPKgerzSTO8gw+B4o/lVlU4y/VPEpGspEPtB
Fsdm9s3TnWoUIT0rRbs6Uq1KVC9y8ANECZgT4MUKQ4in85q0T2adeFMV1xN0nXdK
QU4ES7ZcIBm/CWgThvtj/Bo6p27xy4LtcW+GF8bSyBqp+6CkYGqYaieY8Xu0JyF7
/eAP4G8sqkpCs22jOjLF16Ftuaeh2tFN3zbM2OFpY8QTcq9qaLd3dofXqCJesoNf
BXMln3gTkG9BDEpfD+1Fy+wxiPQR11HVhhANqhJzj+Kmn5h3/tAEMpy1awBKPwaz
E4atYkxjh5dns31yZGYwbbHOoXRnc6pU+Kdww9qp+zYv4tjr2FF+nj/THHzQdnbR
KcoMwCg3TwHX79xuL+1N0UTJbsYsoTq90To8lxW6NX9ZSwGHcSatkLiDm5gPz4Ju
q3go/MZY8QCRzScZcdotfe8qBgERglf9J2AqZ2Kciz5gbhGx3CQjZv+cBzm46eLs
9do8KYWQjKNVI8Cu4+c56zAzj61hL3SnjRHPRPBWOMZt6TySXJqqSLX4vpKGoVih
AFGiRSkLRMiuHmYEerggfLtK7PVCuqK70gjyBLAIk5oX7KKCuFu5DOtpE1ZU6pC+
/P4LgLQ2Pmdh+qe8cav80iAKy+s+OZgeWm3VhETrMmmdu0rljurdahBj1rK3btQZ
Bkz97lJYp6uLNH1z+UlPhKww/Kplxi70SACbx4iJkFc1Ksk86579bsm5yc86rDLC
jXwrHn2DGU/tkojy/9DpjiHBMGJEBmw3LCrQmy48VtarobwrKERtE56yciHrlKR2
kC3oxBHd+qHRZWeJdMzXOrHrdKhdde3vVuUh5An9G8uJNG0l4Iv4tFjaLsNVw/NA
wYRGNiDXuDyw0UPiGavXeN57SQRZCOn6OiYLwQn7G9BjEYLBh4tlut4j91ruAjuH
uiMkVV0WXQ+jeVPMcMKx8Oz+P/sET02BP/TeJxE1+w1WpPdVaLkubK8pt6pTIGp+
ELLcIV/UozzSgelNDKuT/trfaOopjVLI+3nOJG0zQVe3T05W6Mt6+pABEU/m9qWV
lZT8cqIwaW1dDVM7uzPT2w5OYs47K+LGkX8VjK2QLcELtUftoxm7nj+6u2copzqp
nDjeI4bjv5sHjp90VugUNMW/KUyawH3PYfx0PY9GCa/gwin6/y1bM8/VWhIuRq7V
epOF9cVRU2ztqfQvruFh4/H6BBmDo7ZjPTfwO0kfYzUbVu8xfszCWsRSJ8WAl4eB
jAPXmWGXYhfWdJvN9/eF/Ds63RwUIxaYtgO3FN3Z/zZOegd50u7c1eu2EwclBHdW
tAfIl9nf4PE/OWyIrnPFmKvHeLqa/qItvasJaFe2uT4PjXV0avr0PvOY4Oz/q53e
eSpy+fsZq3fCcuUjX+ewOaW0mt0NnAeojW60LLqHNdVMnjv2t82XheCP5foRspLi
PYWMe5R7rtUJiFkY5KL5SCrAqwqe6rG9y5zJk4oDOVfg1tciKPrv5WGLjurRdJ3C
hJHmsArmUBzP5IfRz9tUh7g1E2b1RtijJ2SGHRIWvZkesNuG762iWRftLHgOvoPe
BD2xamKtbwpozBOSmrnTjLCQaO1OipE1AACinig1pg63hPIWFAfw42fg+/jZ74L5
XSwkqBBRzITq2la0W/nql8hEG9CoxY6cfm11R7AqtqifLshelubKaGjW4L6+OswZ
9+l+vPyFGuQhSQusV3FGQ7vTnFNd9X8l1snOORICNh6wU/9TmiD1i0FtkhcJkUPD
syr6FL5y5ze8ZACZtmbRXQBaA3aAAkjU9/bbcOGrxh4pqOFnEnOnMYVIcrw6tLMw
pEkzjReOqzi1cUd9kl9Wmu8v9PyRpiNob8OvcHJDKk7qTUTmeqSg902LqvmPiDw9
wwtdYR0L4WfDGEVjbEnTm/U5YfRV/aV8p7r0F+o3sf56L0qKb6/so/sX739OxPnU
ufSjROccHveME+ssSKJgJcZ+tdD6UE9wUPY/iHHWbISNzMAvEm/J2VFCEVY2agyq
EkDYTI9dlpprxtUiR1Sm7G0kXxEQ9QXxkcZMFkv17rkZpsfHaNlrbN6ga1K3yV67
kIJOmBqhuM7sSL5A6LjORJyPY8oDRaWcETL4KkyOyHgjEt+E3e2SHMZv5UFXAllk
PD1dj3yK7+KxsU0NjaQvCgvSZQLeB627Xyj1y2MfLC2W5rwbJpFjoc6mv2Uqyg+Z
yru2ja+BfLo5WpV57oWdH6nLfRU6zTjNH7mLiCv7/Ro4v2MdXMmKwaYTcLjz3vOk
XJESMLlV10XSpyd3Rg1g49VzcQX+K1BkNeWXjQ0/k/WvQaifnlKsopsNlljss1MD
Wu5c4yOnt3jM8QTfKllDOMYFiNwLlk476papsBrwBv/MawVAYujZ1PpXgByGiypf
0dLSgwQxASohKl7Ke9ibyR8lrNYE2tCDqKK6Lo+sh0t3F4j5Zl1YnrFVXh8MPhkj
I8wXFGJm1eMD3McMdwUvJs2fef/YZtoBjQPyeB/svyOalvpq0p8A9L7YFU4aftAu
F4UzOai2itnkzSHgmnz7qLSjCYhF8r9XAyOhc2HB/lIdxgYedPQxawvItpH7vUGI
otCWSM/F2ngiD7d/xP/pXORIT4IxdsoqtbIcjSi+CQnf+TqZfoirbLp9udDyI9En
L/tIiiFw7Ab2fIL2LDjuX26MMwJaGVey0YrSPoe2APCUMUdBSiiRD4QSQXI1wa2I
Hq3WDEbg6vomFXp0JQjWY2DHfHKHd3vlhbhbCG1mlzApBsumWnGRN3jYMQOolPjJ
Hbkuoa9C5XafBbxVaPehq1KxWS4fdIlQ/tq/+oQZ9d/I1uzdlv8JlCNw4cUmFiwA
+YkhnM66AzrZOBbanxsg/3ZQbm4nvpRgZ9+4XPatckwDF7ueQqc39tNpNE+3cHhd
cHLTWmoH1KuB293hTEfpKmsZtDSrHX4Ld5hpFAIljvICUYC/szK4sfHLC2N5GHJw
1Y+8IhOsF0uSQWW5COOc+nob2kYXq6k5rqLR2xGDuYZ0ovzymRURdAs9XW7WGSfP
5xCdsj8m4U+ICUcwwkRoCcCIMu2eE01adiHjumWAlowQLceZGYzPEMCNY5qnmXmH
XzG69QJGSzKpJjUMsb9tRjKoYLVtR8RGFzs4r1+tWVYE5PnAdsA+iLNhBQhC+0Fm
mfVrAS4ufy8yIFKZScTVcwk2gVL/wY2959yT5Vt27cfSLtP+ouweVSxxI4k7E/7J
Vqn1g+yibYJcXGALpzyOyW1DHCnO2g3EH3BRClqqtbPVpKgXtcfqbjDrG6EMTpPj
k1v9ySZWGjvHW7RVQP0TtNMKWlCc4+Kx3YLMYbJXogxYcGfTEwL6kKzZPsskfgtB
cUb7so9QcNwvY4SRW/aeLQhqmw29bNp2+mVJe0pt173xQ+u1WJ2+uHh0a1xl8DTp
iVO2cF2XW1Q4mPt1J+/jC12L0dRSs8sXd560GktE0oayBGdWOdnj+IP0TWehtNjt
fBjnQvhM81De9707WJr/3UizSF2Qmwu2rRNUMdeDTiHuLjjOu+6D6NvWIgufOFFH
TMPi2Mj/gzdF9zHpQM1uSybQNYTN1ltFT3/3TC4+984fu2GsKyWBqA9nXWAq7Pi9
DeXCs3/UVjm1ZaTwfGO1tLtItePcsEgdJjENIeX9l4fwC84H1L0UDehKGWMC1nI/
nuqs08mDc9iMY9zc7I8+Zoo4GzTSoZmFfXKu1QKA025WieKkC1AFRpq3JJXb8tuu
cZax9c3umFKfaHMXQQ4ZJMsf9IFiEUZzsvI1reu71RpUZiPJk8ReD/autnytqsJD
tN4D85zZlBMDn3stauwQa8WvFh7t8arpO6UEHPoEpkxRS5Ndx6AKJ5UWgPn5i5CJ
Wl/foWCkUwv0Y9Act3WUB2580J2TxN/7/RE77YDiQBvbIixtm71XYDHj0sXiEfWY
48uJtXOn5YL/u2fZgZ7Lf0HPlLvf3pCR5ZVjM2zpeEBBYZwPMjJaOZFKA/Z5vW4Z
F/z78NEiwAyqj6EJBhBAENfnuqCkgQW503dXLUSCFcb9Qm218rkyZwhbZE3rI9TY
AviMuh1T9bHNMAoOOLR9KbI9nDsOGIQcaHq1VYx5LyY+ig5SZpZRAYfah8BNyylc
eRcl9iepTQCuLHw5yUF//Y91UBl0GkG5tGRZljoS7teMsPh7A5zLZ8MHtM7DmQW7
hSX0KgabdAWc5bM0oPFWm3BYxMDFuBJpu4D1HUcrQL2vDqXR1a/r2TcnyY0GJU1z
JhUai0e5hV1qWahQxnX3MAX9IOuIVwCLCoyFM7qmR9kyTJrKJf7d1m/+gA+ug+qh
WdYogPB45Hobt3vo8J3UN/G7Qi3ILp3g8H5/HO0foP1sS17LTgy54kQmy6sp1uS5
eW80v+oa6rQE4U9frz4Cinh85RvKjYpj8y7F6G5g2QE88n1JhbPKk1/cKx6sI2pW
aTQxCyrIXUUjOUSk6johhRZljpwzHRGA5ry1f4OIf5LlL+NwXounNOKvoRegVpP0
MafXcTK7sASUL0yMdZTp9nMtDt/n5m2NyNQAJJrHE+UbkkI55m1aO0BRAnf34mCp
VS+B+aLnhvK3G9zy7Y8wkiiH/I/BgYO+ytXX+CgYdA8vhzgZzFV3Ig7mFzj2tl1a
3Z54Gj9dtIiuEdtjHTq/QysjVqtEgibENMUl5v40bl8r96tpaHyvd4z9AFA0jNDG
39itdYPSsSq9v90fOmVldyareWLC90zgpEDu1uEp80lTZzcyPYZdJTU8jYAF3KM5
Q+QFNpZpspTqu2zs2eiC5KLNvP2alCPYUbccizJsHhG5qZW9PhomPGnpsQBxNhkT
cNzXWrdbCAan71j1BG3EGJLmKj8oWKRw/1MoaDiiOmoLSNwxGngY0FOINHLxODyT
6ySJYo9QIyfBYeJKHxmxc61+uxypQ1TiHWWjXyt0rHdurJ7LupqI3VMJoX/tEliG
TkO5CHLvUz2fWyvp5cnLvcmTXSj/KJAq5BrjdwHi15/lkXVdz7SO9bpHYjuSJqSv
FCMo32KI8e3g3y2Xs+GhHv4BBUdXcugbFqLbT2ysvXIK4H1u8s9FPm+0bEL7fmYd
Lcxr+25//k8sCtQaL4rAlg7G571Cmyoe0eCTF3UQT9N1daRnePn+bi06oBPKaipy
SEeFc7HC2lNXSa+ZfqtW29kSCko8awF+VD2le/ErhoUv0n8ZrGr5/S0OZHeE4Sja
wzTfXeA3tyxLiLa97zKOseU8dfNZogk+PAvK9/ny/NsUmNwM5OSzKN8LGPPHSlMj
FjSuIMiDmqO0YFb100NOVnyF4k/j03SMS/Bpqfzn2pX5nWw/DyJM1cG1gEhz4JYT
cJu7WUH3WEo1taZzEm8y/C8W325DDppd5PjN2TmTdjPtkaic+AGOtaUyGQVpL5Kd
Tzsg96soRRpGFj0lDWbqhYFUqT1jP341dGorTRW/il6UH9eWJ/r3m+Swl52ChCnG
EhgY6/0q+IeBm49oSOl3KLELvR69QBK+qa/8ayeI5b0r0aOKbPxXXNNmeLD1tZwN
Ns/YHwkh0I3IsKanAwofP9G9RS7Ll8yVs88lQ2d6jgJEEv68uhfs7MkfrUdD8AHn
kt0/3Rm81MqEkuDOAWPwSUaTJSCo+khii1/Q3wizBza4H1tOkhvqUDssbRRHCkO6
j5RGgKzngwAGeiduGGc3jPeemr8i+pFt7hMgrPHLxozsgm1I88BR1MmpCJe0jUfD
+ldkLIYCRzh6j3tX8GMyMdhbfG+D6AxqgmmkdzVdvMVXHI92U6jZqavWkBPtYwMz
FZ2seg0jvNq13CpWUc8p+lJIWAw5Go5uG+Zy5+dY1nar9Jceroe31Kobtzz9Mwx6
Gtzaux5Px13tgSiPepTjsSXxWvej88B1iC/pDdb5JHlr3XPA76HJ4qrl6FCVmIwQ
zW55xgX86mfWP0w1TVGKRSVWZ8DwePnHVZNh7XlUXGZjHUBDVnnrqh+fCm8EW+CA
UV2z/4COFfEpooSey1LLFYYQ2Jel7I+Hm00DzQmmNR3flfZK+/CoOnd51xBkUz4G
HkUa8CDuDLJFwU2TitUvoJeWiKwBj5ZjGSnNq93//F7c5BgBpfFq0kUwXrSBpC8f
3l4LUJJIbUrrwjuDqELOuT83VnD+sh/Zwsv9IkDXbQaSA0xWSTGXvWzM/lzhXfRz
jPBmxLpmwm64ADka1iVpWwKrSDhHQ1dkWWlmqNz/xaYgcTi2cRrh5GYBMdojTgDf
1j8CjVmjg2EkO8jKRUtO5nqqtzjz7Zs5De786uIidDZwnj86nz/lYE0FQgFfT8aW
eawvDZvBs04Z+cmSlmhOxw6EUybvYhIMYR5FjpaH6yxRIssNy9E3Uab12V9jy36V
Rf6STdXSzv8bc2w9LRYmLBoO/kSwSfP+NFwKG1VTedl3sIxdA+sYvr3Ka/RwjOrr
HgAPs1fihavj3JHPNNiLIQfEktbSlOYNTJPbKLzsgMTPz3V1ZvNFqLntuMMgDYwG
nOeJyIakQDCPLk7VaBOWSgehgBp06jF/L81tHdv8RDzzCrVUaPzuy2WkjGdUiXTA
wcwQaPNy3KMl1RcePgGeH/7wqHjas1t0CCuwYal/pN9TALTXNfZ3cSVzMhly5O3f
lpqPsNI5bWmPGdac+b8wuTitAnIGQnjlImilqTOnbyP6VgxKMX9/yJfQalm0rfC3
4iK529sGqg4sGy2oJFyVKUZSm2UnhA9JFA5KYuF6K7nznhBEV34s1z4ymSdKvNd9
uLzTZcsXVb6+uSAwdcOPJUdSJ+EnO+wLJaaJv4a27DphA7G9OidJNHL31o1o/p0z
LVbjYEtZvcUMTEUb4twZZX+vmIWQhr8FiFZaATwogvZbh56QcUVCdHQjVJ/rm4fb
/l36So3HDuHHZNlH78Ti26sZ7Ru+5VmYRW/zRBzao0pC3ud3JMvxjwyFyWbC3IHs
lqANhklBuFUM/w/Az3tP6vGPLGNpe1bxQsCqxWajTEpmXDG/wEIdKCko2SfiyY8M
5DNNdBTp2n6NiYFdk9d+luGuAmTt4vHkd70OL5lv7b8PvEsZ66XHBmr5ZnPFfd3Y
n6ZTk9y4oFCyqc7TzLpoNFOlhejuTm3oXzAH9g47SkvSynZsKekdrU2K3toDSdAT
8C3Y8FpsFzSNmvVdzPYMgCb0z8uc/5AZnOsdGjBJFKNTgeZB9H+GNvNoeJtJyUmL
/SaqsF8vZ1IUQ/YdKGWQioW4YWc62pKqvFMjCEAeyi8y8MlkyRiYzTREsTUxsT+n
W9qU2BgFn7M5ItqBur6w2XK1hgHay75TCXjE995cSsv5lc9gCZXrAv4QxKoShESp
D4L2EIs/YkwOlThB61q6eREU6y4FEmNAdgvT0vgQH9Sv9Fe45bLhYnO24IHTcUmv
2BWeOlPfRTu3TY2cajROo7q90IsaD5G0Vi5oMChlRbugeh2+BF1T/S4MsdRtNstV
l2K4JsHWH1n/oXq+cMiShkjs8ctRgurtOkoBN9ZC727FEtMe5fJGg4CQjT7CW7cW
wLU1Suv7+cHeHbnSoBOQX5+8PMF1RAqtNNBMUgisdpBRkN1chLPBuN26G0TqE/vx
i74NIsDumy+vrf3c66yy3ZB0H1nlWF0b1Kp9Rb+vXYxPAV/33e1A6E3tAinUrQLT
QonOC2jAsJaLwWNhm2rnta0ZofZfqtrV5WaZQq36SFDFoO6G1NnMoNODfGpeCbei
BhEHWG/wkTXp8EDPp1vQqs3PQ8lK8mcOdhxI+k/lsk6c8WGfyd00gRXEqdi2YkfN
LVhy4tAcNaxMkL4FvBgEs9eXbZQHwx5lP8BvFSMhCTQfxcg4QM6LlTHsJXr96lld
JQc+hYSgB04FI4Rib5GPKWqh6xKxt6ius5wwICicdI8X4xBd/01JKBxewHrEuF1v
sY3es8zP0BO5vqhUkt7/YYQ4QtjrBDbT/6IIJYkrZOhpKhNDbdcWV0k8fUkQIdEK
ZKkD0FLtdFvZRJ3um8P+KCdhYoUyfhHKd3gIwk5V9QxkUmWrwiei+zbMzelzU37O
NWeJS247drjUndjmHozJjUe7ErE+vnntaVmTm12X4J9CpuhykdZbW67I6VMJJ9HC
zPqNmTy3GPT+OvawJVPGGvW/KVBraCJ/O2660eIC65qF80hcC72+pjleBIIsE/Jg
6fptKUQwkLznAALGlUWkepTPK6J6XoqjbLDYva+tkNnD91yNBtVao5IHRnL3DfED
inE4DwN4l2EOssSD9EBlfXZnb8pQRrDRtZy8BFN56DuFuccaZlFE+CKOh58QsPC0
SgNGJ4Xo7WngGe5WGjttxXf8PhsaxAZmtOP9rHuGA9KLFHuM1bLpncL5sLoyqUQY
Z0pc4ZsM3P9ip7ios7NRhYr1rn3ogBkQ/Mj9dedrEv/7TIcgjGOutVQnBSgJOhOX
+ZxIEU1KG4D198CgWZk/NYrpn4UpwHZHwRJtG3+2TJCEmtizkUwIHwVb6TBEeOnN
sYzfrIrxruXBsAPgzHuZt+Jc09NXCipKQQ0OnEuxsGQtYdvIgacvLPj5ptpQMW0F
VEqgouf7ccxy5KGu2ECtfm4gLhKmZxiMx/+t8UStTJs7BCHpDFSLGqrDJnn1rpRS
ePtwoksE31JMWvGEkhyUuJsjeCKHbcOUK+lpNbc74Cc+Fc+XS2NCsg+w6pCEgJiy
U/z2BmIgj7KB+OIOnAWpjhZ+7BGe+J4Tz7J5ixzR5DWAZMytqS1CyR0Ui2c5gXiN
yNjSxANge61Twn/56N1Wos37QzFz+ATAgHyhpg0XOgW6RFYHbcsHxGkWXxN2mcgo
jNiCV4YQep/eDia0XErIL0wqh5FtQkYKnzi+0BV9DxMo4nBEJ4UTreKSIZ8ofMjZ
8gzUL+7QGJ9zU0OpLpZwwpgBdiG0rAAwlgVrcnmilx6gfta+P7LMOxfxp5fmPCHz
L3hVi3y3oOLgp72U7v9FbDOuSFMSm26SZ7K/61xHW+xT8Uh61u0w/WD+nPDGsgfR
1FOZh8i6VoMyIenzwd/akN7xjTSHwvHkqGRE0mPQeBCm+jBLoanOSjiShYJ8Bfuv
6DpHzot7N2Kc+/h0l5t3oGP5K43CxGS2UM+RI+9aOVePALN7riV5NgwIQeUVVLvq
Yw65SmrQet2Gtwzb2gUrv4lnxX35222O1gR7ljhrCJP3UAd+BEEpUi4SzdcR+z3r
UdEoF6y6mrwSnwInR3quih+VNpbN4UIrj6ORIJaTqfYXa/QFnpwjXmXSDS3TVOrb
td23DTiAVErjn/4CM/vKv9e+vx2wkQ6xzIsUdJkTzAatJ40+pR3fXSyVVUt33Lsu
Nbyl/FvH56fIGdBQdXFg2kiLTPkKtNNwEzQKPQPk7KgOKlUyaujj7qhNskAOjhit
iE3vzi/YGYEbVCIlQj17ENO5QalESFxk39LiUgaUmSWvlpVr80exotsgaw0AVuJy
JdCBc/1xYIjrZZf/1X1gpqHGbXzNwceEz3Ml+dPN7/L4kwTvmh41bjSLjPWijc39
VBvZedmN6P0tOg89Nsh4dXSXN5xeTJP5KwhCvj8NCrWeP+9oryzLzV9TWiHqID4O
WQ9TSTtrjd0CkFVxXGqutn43Zpc61DJmHRumg2XQulATCBWAVAq2DaRs+UjUh1mQ
0dcfoQ2acFPgkOhxB8HJ6zDNt1sUFMfIiE9jXm57asMW/6DfO36o92KqZpZTfAdC
yymuuDkfCBJwVn9FXAW71NCbASLMeDwV9Aeonm8br+9lHUAiz9VgpyAVfJRgcSiI
HahgpU7gINLKxMroNlWR9Oi4xvIWzUw91x4wfLkgo4Woxp5P0LLL1wA4vj6ghS8K
UNw111nIrKbKk2wJMXxTe+QDas6woL88vskwp0iNjlhNKptMxwl2gEX9UDHmKb3X
PfHhK1hxX02OWqhySdq5pv8yOHx6VCe1jmBTBTC8gWijUE0oj1yp88vIG1arsog4
jQRmqNQ6i4zgSv+GLY6E3bn1eFANmGHXAhzLIRiAzLXHdMVFMhPKPc9h38BGjBUo
5sSwzPZ0rociumI95ALlf5xvvI7ewDUHdHtdyWE/lwgRDYkFeppausdO3PTE4hnH
wrttURLAmZox3UVma5HbD4DpV7zq+lQn1tyC09CvkBb7IYgwsPwMrsE3ua02Ujf5
sIR6SFPvK3qYuEqWLbr6r6GXRzltdidcR1XattZs2Ubtw7uYmWGMJFNXM1/0Y3zT
AZvkaRlswhxIp/fpa52m7lJ7Tvvm9kTiaJQvNQxhmJ3kJd+X/f++afZybCKiDsQg
zFRlvz5KiKaXMdE0FzWKU5ACmZQrweW8Qb1KLDhu8QrzZ1wKC1NYuH8lQyYGbRwr
7jxDt1FlbqmLtXQ+k+wbhjwalJRJkowTPYY5BsO1T2VxhysdHGqclr1vvjM+WPn+
5oASRIwZ8bGQzv819feGZWMPKQVmoLzJsWF+q+T2+TCi4nPsGeD6xf26gn3e7ld3
xm8FlF8ZvZzGZ6GP/mfUh+oJ719iwsyOTgOUIABsUhNHF1N435z6hkdtMNFVMb5h
/kaI2zh9+4dCcjhOQtXJqIglGOOz1Z5hNb6eH6SWuxgJUe1nVWLvPQp0KALy8iUw
SAvPXjJ9BZl8yVpeE7BxxZ//CthoRi6tWvOYJZ0t4CSOkfoqelROpeNduuF+DG5l
8w1Dexn10sS9foUOlnxfGJqu8eBP1xdthncq40KLdBbkeZbwsVPdD7Hiv1xN0eXg
wKmb1p/WpwtVMcq7OqJifrlhjtvGKFUINQdxopuXh2dl6zcT8u6qY0DNdc7Zp928
/jCN0yIA2MoN73AY1QKuas7clNyyuek1OWwb5h1o2Dnw1amvkTo79iy5rvn1DFC5
0tbvD+kXCc6o/4KwcEUIXqi2gCdAKf6CF8NbgF9ceHkwG4VMjVpAvNMNNYMOhip8
ViUYkcXu9ZQosnhkV606Xlv7DxF9jamuIfcRhnrLilWZIVSaQyRDfla4BSmSA8ln
PFh1dRWMam9msjiFfHiCfdBJTXXE1sKqd8WgHr3JjGOpp0gD1mrmf7AK0exIP17f
OTSjFvH9BU1leITp65oP+X63Cv0RBubOEP1V1ALTeImctV4KdqkK2lfpxrHurlzM
Xljta9pU59LVPSMDTNrQLbMP3wzvXWrVp8IUrnCi3jxkmNXhxnkZsm6HDmJxaMUd
NViTsQuIAYDPdwqU9oHQ9fhoF6pFUyWIRSA/DN7EOJa8z9C+I3Ljb4ZlTZ+2gmQd
7drqqxsYDBaCAKGY1VYI7psL56tnHw1yM6rb+LgowkTYJqf9xPbtlCAL2rAnjGc6
JmzgiOxeICuPY3imhKV6PwuAZUetQXjGWlYU4EB8836XN3vutoI0cRsh4nsRW4gD
eEjHDI9ZVMq8kNA5mx2KRi7AoNrBEIxfyLRCDTwgv7grYIXVaUK5tO9RdJvaEhO8
yoQPQ3jm19PCjV4rbpNZicPcz/MYaenBezXVZQO9781Ly24ZkHODYw2J4W6UqEAm
1jOkYhopzqjo7GbOXG71JzpeuqAsSTQ2kIESU7tEnncS78/jphymLHozYZKATmqA
wgDbfpWpFceJDOZF+XGV/i4ADqK03XP0Pd4f+GWhCPVnl4F8VX2cXPu5v4Az3x9t
MxlRIOUGTHKzrL+u8pRmmqUzZj+4DS4qrsEx78t565C/DFMI3pU4KpM9WuQHifM1
nTh4ZUSNC4ijlEmVH9rghA4oViOuI04JaHhuUmHvxTWtTucSIsCJeoyt0Y2oQ75B
iVxOc0ckJBH5Zuz1CAk1ZKmxi8sBBF9e3/hq7P6UGbvzXnAThn9wt6kDyrSPfI8u
wOpFB0k7HPKJVkeVtJMtp7WG0sQPvXoIiLZnEit5VGXibdwh4ff8OE545Npi59/U
aRhzm6OWCn92QyggFpCdOiyS7FZ8JfhQJcgC4We2IBU8tpL86t8oAj+yKrRUiOPL
igjNVAM1cNwIC0LLZnYwAySSGReku2s3ztOe319tdDyJ7xMPwdJKpSOTdlPlGSL4
jLj4Sq+i0+mSPKMzhNXo8+nG7bUPg3NTM0kqPepnnb0NCPtICBOBHCgd1e6zo4i2
JmFyENH/2Pv/g+zJllAEtw6Wg9WawusThGRRoldw6IU+9nPwfrWY306vBDJbsjqv
Ga0aI154w7UM0NKXTbsvH21rapGVZOqELoQdo0J4S0S7m2hUtbIXv8Q5Zxdf2sCG
URvvUFEkMeXdb/7cqBUB54Gi3mclQTYJKVtMf2mHV9Q4zs3NhJBtFg4BpnVCBhEC
I+pfxLQOGfQd3MMrvrRNK3mUbwZk725aFaCoRQMcs6Xz9m3A0ADa8MY/RDv+zQct
uGUDpXPf6YC6JlYmctEHk3VOZNy89ddSnc0fCt9wMn75CzOZHUcw7taRM3Vxb9X8
Wz+EeH4zCGtSBOZhkAzekE3HCMOqr1w73RvdTioi8dQXyaJ1aGUX/PMlxyyWlAkd
oWg1tSrw8fEopc9XqNsmKOIt/89LO/bCwBv6+E2GvtjtJ1U35CTKXlg0laRODlRv
ipuQS0Vj1UebVv7O/L4QLk7LG+XClFMSWLsch6t/CsVGoB9LVSudJnXGUYug8+SG
tth69MpZ301y0y9JyyaiaH/K/fluGuTdJeSdruzI6eIeqr9N8TO7Ff6tjpiJRtux
9mIa9RDpOtAWohpOHrFbu8iHuBHhI8OuszDwjD96sgXccoTCXnZGwAU3BXvfO8n4
v70ibsLd5gChdg6k3nLq0svlcdmbT+Y4iX+2TtXfDH3+P7GSwT5wxKALm8TIcJkT
OXlqZL8rw6klEW6ZTmAfWsjobvpV6kGE3MhOx/FdJ20P9wzaE2V4TNWjg4Je+ztt
lDPC1zXrlPiGewiSMwhRThn8e3plX37TzISdP+V3U61sWycAiozbQkr4+JxX2jMv
r8rUIgPAz7Xw2H0LM3W42HmbO6vHsygOw4j2RyZmjphD0szOJ1vakk4WcEZs+VBq
I7ecRbVQCnnc2foiN4cpPu8A0teWA5nWdH3s3IOR52xypX71BmOhSoBBzgkQCoSy
qRveHm3QoudJaW+qKMCF/pHawA8mJAiLTj/p+BX+l+lxLeGdkFKkUJ6X541FvX/o
tDyh9fTBLZNPVrPVTHI3EdJRmOCmlVSM00uUZQYctPpIK+qHBKMy9UysDuMmEDny
ofPBru90MWfn1Z6AAaDPKRCAK/RNnZAuXU5cJmmGnL9mojmluEgdUp+iqvJdE8xX
6EZIu78IYt5aa34yL9YgE9eWju5ZoSf7uKC4lgkz3lOmUKk+K+yLy3cSHe0KTRE1
M8nSjIol/ZhPa574Ntin155p90d2rKdmvoXfvTGX4jZGgkowrE8TW4R5IH26nP5P
+sjtK/FT10u9F0zFl7+YLakcJkUK72Xm8l2Ho4wCv0ELAD2pxUVPdcFx4ZDrYteC
TCPowPrG4hxjRXJY7+qNJOYyQzMN5wyhbArVrQb3pP4Lmn5d7IlWA9Vc04rEQFL6
U0gUzDHYfKpitUmSjM+79pEq0WQVWhS6fFwxlpVC0kCBVBxTMQCHKPnrr39rQfpY
Q/Id/9HS/A94XRXSdkB7uw66m8tqolxexcPd9hZdvCn8IP5BjtJvldrJrf9N8S9+
mH1YMvK3dY4OHTp/jlKyvvpZjTMYhCVkQxIW4oQgtVo3jTH7mLG7/uVTl+HQfefe
wBr69T0pvKfhiHvuBE/OWpX3C95MilyYhEaWXmKIqjKZ/TTYA28I7jlSyUxNv7Pj
SSp7Sspffn8aArqZ3uA6b8KR1GboSlRrc3gb4lIKSCfxhyfx5XGPwd5empjyONRj
Lo3+nyXnnzApo+DVzrz/+Xf8Bt5txlbI4OZzdCT6523CJRqclzaPo7pEiDq0DotV
9fx4vy0NABaCmeXbtXJgoJhGo23gsk452vSL828ML+9dtG8Me92cmk4qe5OocuG4
0A7coBqd9/Dh8giZ5SIoqTJhiXcXUXiE3N0N+YO+DRXNAQv+b4kVQF3hcmmH2PoW
IaM32mbiqPpPlXNO/4xFX97gu1iM6/k1jdQXvxoU88gAMM0vK95KcujLP+pOCiGR
30hO31tYu4hO5qAfS9JTc0oTZ8KLL5S5hHvtXSnc0fiOPdA0datA46Ht7Qn+thDU
lI8bxn5Qu2nMIA9kTT9qZpQJtmCI8DW0ReliEjS8DiQztE7jnF5ljlLbU8jfuG8a
M93U5h5pBJYOVUuAnwcgqJLg2CQ4xyEFXx1WJLmiXdSbu2WSjdn9NVIjOLRjtGRg
KvoO7w3EW8wRUfc0RXG51O1wcfIwlIZS7TS8yVpiv4bv+HwBa+8H4E+JVoiYdQfv
PCdp1cfZPOvbpwnshGK397CZx0/tG0VkZ4oY93xdYoVGisjYeTOpqY0LeeXOrqfG
qmjA1GH0yWHn6IDLqnZ9cxZmQwcgVmFOK0sREmm32dtadp/1O5Q3+3U33GlUTzFg
4yFTaxch4nGwemHz+BOUInb+ymtG8fJdhIP4Nzs1mPyHdv2qa93Ma5jSIwOELT6b
wh6gNw0QH7m3FVWJTLOFQrA54MCc6fAowjjXAZSorVoLzhoSN7AdSFAMED2ZrhQa
dm8OlLyBcJYYNA0zVSmvrRuvPjJuzTTy2VZjLiMX1n6wCWC0unBwZwiAwyhAcaVr
2QRA1WGRYGb+XciXkGutAzmS7kYL5Z4e7TuElHFQeRKtvPxflGCGAP3zitw/TLnE
/66VWtk7pPIBssUIO51MLdMxA09vbG/3j+gNzhF7gQqI6zBFmkjAHRGZA+L8i/Dl
g+ciVpJbutzqlMM4UOwzx/Fnl9/96BiycAitddhE4TOaqHruf7G4r/VavyQoDvsI
5YxlAUYNuMbZJFszgEq0cSCTHiqRZwUzOBXlC4sBduKW3XqsyMUOMZcar8kgKHD3
oUhM3vowXOcCc5/z723/Uwdb+YV9x+AFfi0WHcwgpbb8MPvwt+Iz6jx+Qq02Wc7b
itTwhs6dprRTs4cIeC0nDo9T8aJ574t1Ux34x3M+ezA27cA7S33OfaqTqDUZylH1
fMm+yWxncb6fkBNDJIVhlG5awXwjXv/6jzS+nhwunBbb3YJgoLx0MfZ0Svu8cNbC
bzbWMJbd4g63myzbCsaCWiDSmxwHG0nsdtVDqznS1IE/10jeXu5bSfNbPjJxHO9A
47O1v9ia7tl+IrCuq3N4Cm59hnV87bQnmoK4aecl58d/T3ztBfk8IEOO1TwotNh3
Vpj2TkngyapgdJdbxLRwxmr5c/J8DzP/UTrKAg+7YdaQFnEn54k4Lr9AA8HLcDzq
3LDJ0HbrW6w6Ok0DSSWg/t50QyWuiYvTZEloJpfbtWj9x3tgt6Lr362G9yVtET4F
IDVUhK+5R+hRFGmWmEMfpL+BQG7g1VH1LwERQUydo1iqFV8rcKpuewZHKzaCPScM
J6/TUUBfDiBA30V+3ORxdPZpZmsTDSLJlEJaOmPUIbE/OV+E7WK2AqxkTb58UQrM
H7/4KcqBYo7uZrMuWWeWOgj4LyiqOwRE2qf11sU5Y/NrjornV8tU4yruo2CrHLQo
Pf7x1HEnsy6IPqpMK+ohob5UEgs2BgSEuaNwMWuFOYBxp8zcC1TgYvTztt2Svp4t
B9fTTDVro7wcrHHbaqOcZTO2HfNbF+PNfqpj0vd2aJBA6x9PpX0c1KtxvIKVCAMw
imSjY7SDbFswjOjAYWOOxt9ZXLC8lI/Src7fRrEyrwLqNSmLfJCd+tw/JdAX+i6f
0ABHbC6qXOjUsXBpBLqTvIFai3G/k2+Xjkq4JCkwdaPrSBeT9jLUoBv9phfw9gqH
oPgtWBf3uQajsDlBujJwqDH9VADaOXcgN/TGdyH00j/ANlthMptLdXKd+4qWPF0W
VQEYcQoyE6H3QSWXHqtU3W8LBlAeyPHYFQXTGhYgFODX+jZyBDWlQWzf8M/ySM7F
pTJFuLwPFRBmwcNpO0Hh/HLcWKju1B7agL8JK10G/Dqo4hdHD4SybR/4YEnW9b3H
fhXjwUdtOsubhQVTZXdH85Uo7KGexLFUFZZlPI8UnVy6wtgtpDXr6ExAJXr4nzOR
/xz5ZuUd+L2o5gwTS6vcdEi47E6GOjItjE0BwBmpPxmQe1iThRrkeCpgW3YvwKe1
M6gRvp0PLCbdMXrb7SOVOq9WraGX82uv0J1BNWdq5IrLKsC+RIfYXPhLrjA/4n+V
CPt5AtOMoi/l4pQgNrpbyCNqqaaEEC9snFvVcRPdrGjB1oW2pm2lW7SE23As3HiA
ErWAWiQZ9xpmm9nxHYY5bCMHbUZ/MrJDeuP7NC2oyQUsZdqWNO80QlB/Y184QsQV
LjCC1oi8v8W2nRToP5SW7LdHe+3m9fca4MMRFyokCA/HvkAG0X+MkqJmAO1ZRZzi
SKvDp7In3caXdBD6QFWZSryFLFhtwURmjlcMdD7jVs+Nyxxr88/bjj41jWdEdPfZ
pvXDPbn5dknTIbWcXMkxtQ76bTFx3cjOmr0GQbNbsK4KuIoSfWRWBaLn1s6iERe/
lufkVlyQa0WdwBFrdOMQ7s4vSelm+Bntgj1bMQeC+60pN75J62UegieNEliXRY7A
X5fgTs/OGcpZQUbohmllNb7J0JJCw1oP7TfSGY+kwdl8X6Os6PVijxN66J3Gg9h4
r/qRwgv6BrSuD0CapzRdojw6naDPaZZ2XBcIsS7DzWMKclfr5xrXwvQ2rrxRGqQx
mfzMFrUwcu70Qk3TJL2iHeSSzwT+UwEMMtc1M7tBPwVJHkXDwqQC3KsnbAwKjhCw
K0ujBYl6FMw9CquF6ZhrazFDeUhAS5a3E5tHVhGweU3vRcKiAUwTsbosPUQDeozL
JRXTjcydy+y9MFCsgEOuGWxQvIzyQ8LFjil3qjEbegUP4b9h5oW7t3q236UsN6RO
jtLPGCjLzgWYwL4wy2J5uiFK246CbQtl5/4fAkWH/osT0VaxlNE/Mm0/uNgalH3o
mA9mij0glyrAPRcOqLpJ1fc5KbhJf9dC/+X2zun0RdsBwKTsH2x0kOpR9eo8skFq
UbFo9H99+g4YUnaLGv/QFIO0o6v8Qd8APmM9yePmOFA6iku3Jlb4vig/3o3A//C+
WyMre/i9VYiw8iTL3F8iaGWhDXfRckFKxNHWUpP5G73tbdMs+CzXDyswRaYF1jW3
A0NuPH5fjQQGf7cY/YemH7auAkZM3/MU/y84w5Ld0bfzcWSnspSJxrxEnr73UN1e
FR0bmwaXxEs8H1dMNHZri/dmzrNZnEK/SoR6awb+TdKb0FGsTpI9Xsu5SFsDTj4t
fXEpsZKs54KH0I0cquc7oAgHDh/Bl5M/pkPXrniKYPWWYDuow80Ssx3+GUCERgKA
z8KT71l47Wu6qVrVhFQvrLm27n1ij5fY+RiZOT4VyJG18ErBciJBTuIYZRJvq3ZI
qwj0fJcA5tgsN8uEbMVjJyYPx9QkXqzNwqRvx/gVDoJDKE+AgYetYy/nI8E22yrz
2oWP0zaFrtPdJQIbdkL8maNLVZ2DPlEzqIFgfhsYuz7DxrLhx9pbuvk5ZAVzgUqE
8/m1ac7FsKcIpnt2KRN6V5mxP884evT+xdIztYesb/hkicfZEUUEj7No8t30ClX8
JsdxLM/fDBB1mdpHMyL4fjd+nj0Ht+T9RkIh1uUC4yn9Zkv7wTFeB7OJ321IhfXO
i6hIAmqGjXtTi84x6rQyBQx96nKe1NkuOCuAVgQ/rzXE8O0UHzFCmh02HOsN0Rc4
xsHR1Dlije3nI24S7wA9vQ==
`protect END_PROTECTED
