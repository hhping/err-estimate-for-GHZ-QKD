`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kurIXOJ6U0/ggeqsYfkX8MYbrESsS9rueXh92nzBTx0/YFc3tN2GQFwaB83ILAoS
jqA8bQAMr9fW4sPcKuuE2zj0E9BvhU9INjtNjrDXK2rfcBMxLpeR0ShEBUF2v1/R
XoEcVBIGQ7GvD+mBrBreUlZIyYerwkp4WNiM6d5nf2+ka9XPt/cC18gNhcLlylge
svhsrupYVBlm+ADu7K9pzr9AEzlGoTbR9nFuAGyO6LQLADeVQBT/u3g4T0nsdinh
Tb6UNMxu73H8CFD62ILoiV8fa2i/1BiL48b234nPXxY75vNziGRD4E98pH8w2VlW
z1XBz+DPILUcoh93rM/0S6GFulDdIGhgVI9cyCmi07sZy3fSJFf9EOzQFO6l73sy
wwDsH+gHY8Yb16Hul2TVj9XJobxftzo3FfK4bb/yYXEXsSvPHzCdNF1hlghd0pMe
XrcX0L7CQVjFxhLFL3tQS58POB+i/uJ/C0zLSi7Gcq4wB+fbyu2rCCk25Y9Swguw
aalDCykGcycHjGOr2YRCU80dbco/2PYd4+gKrOGSnJfILq4coGSndXspL+Ve/ce2
HAFFH8DwRdMk26MEvdniALw7JKA1jEwf6J4gi6YkOYtkOrVX8XE+6zlFLOh1nxsE
HZbWaP4ReCoGxgrSSTQxPNpalydWas4uURWD2oqVNlSxBU8v+n1aAnTC/SMJ1QxB
X+v89M19qaeS+IwWV4f/d+yw/EuMKLmYOpUxp4XMIR8/EcKmXmhyE2TuhxtJckkQ
P+WVgBo7vPbU+Seikp2illki/BjtKYzli2Z6KGjypQT5sHYNGSIbf/a2EpMBuyti
o96CsGJMe44gecXFx6CO7H6SheI636kLWellMb+SoBcap14kDYHYS170qu5+kwTT
jrTtnjlWlefyrs58e2cHezsG4mPoNN2lYSkQmwp1frV6cPbn76WEqXDAcHYDu45q
HgvVa+2lNLzlcON0u725ikqWTRneQldZ4bg2Y+CL66Ht1ts5e6LE541BkMFgXA0B
wKwgkIjShd6UhIP18nRXrWHvOg5bnfbmgCcy0an5zuPo2OFUjhQCBAJwlb6RMf2B
a9oL/hgftNK493o07HukR6xExDl5DWMF3lHFcaXXWNhOIPfzCmtt/LnKHLv5gabZ
/nfgh/dJDUpCPwmX/LwsdG4eX9w5SU1TTIaNvDztod4/l5xPyrhXFJ6tAggBS0Mp
Sgyv0bCeGdSd0UPjhLau6L6xXdl8qV2fyhGFpIoTEPBvhvUFZ4kAnsO7+IJH4Jav
dERJySGB4wMkUak9uZ+l0HAP3JQaiwWqR4dice/gCT8Bd6pAWwtZxRWw5VO3sdzn
GUufjnf8+7nAiCFMY5hx9/qKn169AtdNBvqGDr+xrboy3qPBQV6x2Sh2mAALtEtJ
t8qfm1B7+TVzImFRk3D4JFuRPNQ/OWB5KbLKxFzO3tso2cvW06JgsmuqdYGQi8Ae
QJ4CXkIVKAZ1YTxB1qU9wXGbOcYZmsjLuyAYgfW+axi0TlwugAU+n7rOdxekgnLH
RRWM3vRJ5w1qdcbcoL//GM1Peuhalj2d6QDZFSmZXbR6DfGGHZCv68AZAELL6OoO
q4/ks0fFfQwZ/EjhWlWzzUEVtQYkB6YtUvPwOwPBgf9Vh5e7uvW+oHgRKVZvvpsX
6Jl9o3qL/E2K3WnD1rW+1ADQVSgJfiVkIGbIM5RaSTu/xZxmDSla6ESoyNTHNzEa
TDpirG71XNoiFne8IdrXnw==
`protect END_PROTECTED
