`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30erHySRruXnZm6W0ljPIbTdEXZ+MPhoj+ezWm2UcwDZ+Q+UyTVh8UJ7HbXsHh3X
S0u5F7XGFzPdSl5pZ2/JoZYXzcNzrIgTe4rNbkpxFlEOOgG/MDECFzIpX6swOm6/
L89dbaPT+jaBcT7AVimO4TBub2qHKgV3KxqDy8nN/FZ0ny2t2otXFfNQC2bFIUgj
PB3s3roiTkF8J7vNPRn9Bu8WwHftI8TLTC3sV/dn1TyhDsyC60vtENVlz5z53VeH
S4Haw0izb/+bWD0YSvMxi05qwS5vq+BkXHXtQs8P21qqftogNUaP7Hec//aPfa8v
0nCPm3qxUos9ZA+jajggzVrHw/5HKzenR+jfQQAwOKLhrv4CCsPQKTdZOMU9hsco
hqVLP1HC7nxb9xrSEi28gMX9eiQl5Cnmg04p0RzRk9UTbjJzSN6jWTFf3AcFLgOD
p2fwQ5ITwpNDoSAb/0E/7ckH8r6JkdPJF5eqMqXdCqR/uhWA2WS3052J5jbnIWx0
jXOgIW8ijSHdLc56u92v/tIjTbyNjeQecdxosTarMNZMCQJLAR+QrOb/V5cZkImY
ExdRBJiuTvGl+p1MGolC3vIv7ZJqHgm2m6ZGstXPL+lES/mlhQPcf2YIiwlLD1J+
qM1RNeEfc0ON+XK9hw/tEbb7HnVmXK32B/vIPtj/9pnmv2y+jxbfsgseCbJgmH72
5tHR0Y0xilY/x9gFB1zzOdLPJFeWnii8Ivi36Pv/Tjvl9huV2FX5Dea7zPJYpfTh
Zr/zSJJnZtJWOUt4bcrPx/DAqF2x+Qx2gfUzVgrFKE9JlGe43yW5BAivYpQTcW/U
RDNYmSdKIGlB1rrX76kw1TZ8Ej6ryaHyvX/luWPkIMEf5L/OpRWmpBJokllsYhF5
B2VTuz++t+R2QsdWhsXg6MM6cvm+DMbwCdDzSfzyMmUydWFnzU5Hdj6MAkm7VtuO
1iB/Nmg1vfXh07f3J3NQdgqBrk8m5uA8iD8SEgnyRkJ4bBtnUe9TWMrVkaZaFFdn
vjjKo/wosIiwZo+Ei0w/XEQPsoqAtW6OA8dy/QWPRzCJnfm7k38wXkXQ8TwP6CzN
Cmby7toxhqX+JwcdOSUz4onfhLXwAvYo+oF4CTYebgfGuyF28m2hmvppfQwyBeRJ
e1ews25rKo4icr6B6eqR1fdkIc95+MT91SIzCwKqvN5MCS8pBbXCd3rjZKoH8gZc
6dHaDGbllruOW3ixQsAi6RATglm0PsV120OuARu7LN7YPVh4Bnv1CK2lvy1jguKw
q5/ng71nf/GSG/9CLJv/pKvGLeId6I9lkD145gnwe6Si92OzcPhARROziUyS8tXC
fTVeiDT7HVpHrL2tLMCuozKpM1yK94biJn+4NwjnNwN77Rfko2rz+BU0zNizntzg
bJe3VI/548oyKFrad7p8rtAnzdqq3Y/MhJZtcOi0INIucUxTDHKaZw0VghtTQWZt
zWAggWKZKmStH9Ip49vnUc+nTN9LdR8jdtvmprfV5YAmCOnh8d5exqnZdDk9gmB3
6NdlQOLGPf+q3xmJj6TrHmdn0t39VMhGm0qYelvONk3k0iEW0i0ZQqb8QNW8QqWG
d13NqeIlK4Aj2+6tMQn4pZMkjXxEiVL9uFPOxfYIRWv3G3E1v7XtNYb+sqFx8t90
K1BTR32mF2CFm84N6d02hYmdrcpCUqre9vY4HB0YAVUv4Ah7bn/KiZ/D6je99aPb
Bj9G0oKOKYhKpyGKEXiSp2qisoaa6n5pqqSktWJMkROY5JqrB5cVPvBNojKzpGlo
5FkXfXdfLtFotkUFcNgme1w6nHzTZuEt2ZzIfflboByReAPGtEpbTGRPUForvJSC
ur6REXeuo448VQdhLTUSFUaB0paMkL2GhyYE0mNyejRG0CaHPCg83QckCotUoM5z
nLNZH3AfOVEdws+m+ZP/Ygvjc4FV9OFsj/KBU8VUo80xZ48kM74OwKVm67v3HKGf
gY+RIKXah4mHdP7r/G841sG3olTKbloSjVnnC1j5gAtR5r+836jvf515rTdXNGQ9
3AYzf+vvgVvm4W+c1dyo9038QpQwc0z8i9uC9jk8fF3UbSkaXO6Bp34vTXGNHzsz
lHqoUMN+xBJTlmxioLYayIbEA9Bx42sF23Q11C4ghHC9LFg3pFTg+Ya/ZRe2sywE
IVFuyJ7ugzRxrKJZG0K3AvOIjbmfbcR9fTlFj4N3ooYZksktTMWpuCx8OzMRPoT9
Hbiw2IifuBy7ZFqQt94SANKQBke7nyHHa6nRRKJuRapT+6RzgU8+KNrRWLQXYcwN
lRFUPXf7dWAV81vjA0f3/Oqpcd0dmu5IYx5/LJSs8uY1OHNLLUrRhzOZrc0tgxx9
JoI/j/yjG+G37vbo2MNVcHhUgPJxb787NMs4lG6WYx0QJfVqEKq/acgMuSocswPi
X4RbIKen7X0c7nLxbXGXo8zM2nI6jW/Ga4D+jhzF2pYaGGSxcx87t/maolBf66Px
KNoy4Pyv0fTHqeltb/VzLXp3eFUjZGmYb6onk5eBj7RmYUPJN4dh6FfRUxiVcWU0
/9xisdFh6U++4kIKHxJQFfYSc7XIghaXYWI5VaqD0jjDZuFGAhO/zznI6IhU+o+9
8BwNtOyPpB2ry6V1t+Zj4IS473Omf3ry/BlB+T/Trc5kUeSlnqbpt5yMc3w9feqe
dgLN9CI1k7UFQqghFl4aV4ejgCy7DaazdEGvCIa6rNMa9juf8FdiaxpBo5tptbhE
4LlIqgDw1v1qB12Y7VuBLO8xAQC6QkTAe8ZcBsJ4pvTLzixgs32MkCHOxWhYFfGV
0RviVR8Cb8zX30Bjw4NCRsOyU5e2C0/z3d+T6tQWWJn+ah6/dDvVAoEqnugtshq+
7fMvTTpop2baHs1JZX1e8GXg1qUsSM2sS+perveA79a1jaGk0fexU8swyzjaZF2A
dASjvu9G8LO6qPT4hPH9StcNI5IMUwNCjqqdVBb7YvIvvFACarlh525ikw7pyEnl
kmGb9UC2X0ZoR/kSL1KXsLCO592a5pszK7+4VEHP2mVG+WfGy6eHFcuXSsYkQ6Vb
swEWK9sWcNCOE3XG6HtuXSGsexcq5XccEmdbiHeeh8iu4qEZ4H8JkuXuOenoeUtS
LKE8fIgiXp+NIn9j6JCHabD2zJ7UdyDGRdgrUygjnPMNmTcZdChKdUeh6IChwF+R
lChAs5OUGQb/C5moeLd+LrCIA14ZTGvLcxBye7TYaZjlHdH76Ck37dP811ajlnr0
rHwJrp0teDlYRo1scWhgtZ2CEy/fdST9Y4FGQqshMs3T4fMiZtNwMVYHO72E+KvD
6Jhk1K4UXNgo4BONN7FQ3Nj5aZAcj2x7/GVYSitFEEgmWxv/XJdUXvHVZWVY5BWP
9c61hebneRlcoYKmMdb9TVZV+WujjTHo4LJnBrYBOB3Wrx9fO7sVztPe9O1JCyXa
9lxpWv0KLg42X8fxaxBiXbL82Dtrw6/BE+GRJ7EBP/BPtCdTZAvM7Tu7lbyMj6zr
ZmCslm2lQiBMoo4I26IMsEJFVEfgujCdEqiByYz+Ckoh2LAIpFRqaW89Iy9ZyGN3
2jCKeayQP1Byw7PBhkWQrw==
`protect END_PROTECTED
