`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lx8X3PO4b6yTiCRhCvidvZdcjNNFex0Ec+RHMdfjc/n3Rgx/qwFy7DCSGqdckW0j
1YHSZgcyvJjXr80dONRBr5f0o1heER7ifiohGXHIQlGiAusgcs5aVznMaEUogGJF
/ZFFVfG3mXkUr5yjcP09z8zVgZbwkYZ0F5vjMdR3bqfM4eKw0yZocWlvXwyIOxhZ
j/T1UrLm79cG83fmjDwfHGDPVkkoylzH9Pp/Lp6sPsVe1zayFlX6Ofm9y7BR5ivl
mMVMU2Tuv9ku6EusKF/uIFN+lrVZhifJRZv0X+E/43c=
`protect END_PROTECTED
