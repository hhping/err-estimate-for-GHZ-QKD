`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/t9z1mxgdaz8HKxK98wJhCPziQ2jshoyCSZ/jbab4oV9G42ocVDL3rXQRd8eIDum
4xY54XglWszzaResWvoMQTJi+ZNhaZHZkUhcLHnsChS+S5ItohUfXz8rO1usmDW2
HOnxwb62ylKPcwYsnI1kveM00c5LXFclAJyemrAsaRpLCEr0QG0Umnwx6yycEbtv
vSc36I3436bP6Y8/KL4AmXkU5zy4FNEJHECEaJZKxcyrcZF1FmuL805sAeOlwqQ8
qZi3eJptxa1g/XXEBdnevghzZ/vRSVjGRO65++RE7vZoasSG9wzxABmfQVP4MYSq
SQF0TCE/LiBqZAC6pYRjj2jeu/BjMD4zcZkMTWCQn/IAhfoTH6Srt8/ylXoxCOsd
ztlmTuP7zdLE8YQcMSv5cAzPXK+zIYtQaqbLoKJ8UNl1HfJLDhbFVeBotiwb9hDm
wYnNIHJDK8xl1+7N55eGbH71xityO3xQi+3Q0gLtnEdxFeSj8VnTCKQJlYzv6hUq
5qBucvmsM9PTWpNUnTbZks695nbj7WgIO9iHQ/p/2BuWZezOcJVK7yWh47U8aj7z
gLiXZKXEm12gjeW+Dn15kglsTL+zfqB1yZvtocLnQYSlHkUdSIT+xTQeUKqh2YsR
Stk/F5fq9vQuX4+xLrRPl+8jNg7Gih7YDxTazcdNetVuS1HmqY7GPsdwki98j5cs
P568+7WXX+hBw9FGqOCNUPv11S6Bfo1/TihQQ0Dv6qwIRFEP/SRX2ewS6t3ONMKb
LAqpCCJo24+pQLAqDROm7bfG0BAMgpcWbMNxOsZlsd6TIBNKgmYh651tmRlyRIBj
nqP/oU9aWx0wP/lVIhQpLArVfAaoGhbuinjnfQrUzOgv4+85pwqAMYMBgTuHSiZa
ZDsB9GjQe/ocnhXhTRW1I8H5ijcc4L+K8WCSuA5kKle/fYgeFnuWxr9oIG/I2C99
gGBlCg5KmXCSiJmDsZ0yT4SzmP52shJqk8s6+M1/G/KZFx4pdQ/tcGZyZYjvC2rP
cPSyOuDeM1BqL76NVU62UZeJ6x1I5yClj4CW47BMoJCnNeB223Di6UHtQl/DEA17
rchUFwpSrPb/ZTl581vfGTcxJquAnVgcLB4l8mgHhaDJSI1PTZnykUZ6Xn4UnXHa
HCOFhpT1iQ0/o/WgLJi6fNS0evDq+gIcabkaAhzdfw8zhlmx4L+Uu5KOBDUzkVmL
Sv1IPaqNcD+6l69zMPRvsjxatqIYoHaeiZKWbGmVI+zi8OxR8NmkPGgxzytPoA0b
m+8EcqzDd+IngvLeS6u3CBxfpINkGWEZ0S5XspVYlMsGDug3QpX7qMEBoXVJJ13g
BcLueg3t+8R8259iW+bfs15gcxCbkVfh8FrHe0RMQsYC2sJb+B2KuxK8WbUhaTiH
C/qhHwWJj2ZdJj3VE71bsN5ec7VCPvsLB9wLzZaurwZHhTcSVNzcm6t3fa6WhTGH
U2DOV4Z97PixvrQhvq2xU9Auu1QT46BVPB9XjZtfVuP8fuuDUQ1+Qsd0MHVE2r24
XN9FOdpn2LD+lMily80YVjQf4dV8XAeMb/rWuKwHvomxNdJN2H6dr/eVDYa6/E+W
SiKa927QWM57b58CxstGm+lrJVlC8cnAUTofGRkD4SaKIibBIIVdGAWSlEuClXzF
v+LR1/bbfQP/TRraMO0sEJue3uAlAOfZqzWWjMwE/bjQR6MPBM234UQbd6rYf8fW
6aX0K90xY5jw7c+cvtQcge/EAwgSAMzPveK30o52mnYcfAjLnEYVOGn2sgFWe370
mMvw8+u47TiXZRyRy2rFXxqPdf8uglvn4WyX9HWn9Nnmfc+4xUcfx0qJx0QnWxFN
nvgiAoedSK33j7cs7lz2TwdhuIpOvCC2mVdbmYX49SBaNampLVWCalnUN5ALdQqz
OBts77Vlss8FzryHBvjt2YKzDe1lNL8YAjv+a2BiKXP/dsjnYWf91QXy8bbR35kN
fDVmj5vTzp/VP2vEUPgXsCuk9YsWGHUoc1ms/Xu072LKg1s0+ae95UODlX8HQ8Eo
Ns6Y7Rlp2C22ikoebPC1MzE7D4A8tizh+1v+yN8AGItYn40F/BWquLsdwok4/VXA
Iz9gnYDLgoF8TKfBZMh0O9WRzk5XGJA8gPaDpoGWAiEt+KrXoYStVWqIAf1tpt//
`protect END_PROTECTED
