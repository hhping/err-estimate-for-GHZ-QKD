`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MQpsohU/Du/1Xof3sMGJSIuWHFrlKOyoyyRjcuWe++uPWwLXzBRj0SJT6J8JXsP4
0wmjEYoAppj2eS1J1kBAyOIw8ko0pW2nkr14MeAfLfW4heAo3Q/p/LxVKYuC8Vek
PpVlZn/x639QdjqYnDBeBZVmM3mgpz9DCR5uNM2ZWLS6B5d0VchFn9JXH78vvQf0
101BCsGL9SR5nt+qfQyjgdK4kku9DpltVI10Lggf/OPQQS0WpLjot006mnMfjYe4
T/lKkKBz2iSx22BuoehN1iT973HldWgwG5Wawkn8EGPYvi9O0lY5YjUZ5r92nh/y
Z+beYE20OFpKvs3H7vxkMY8qLDSN8Ek4m2HkPU3w1A1SIWUo0UCUIfc+xcOX88uv
4x29T6rTAEtOSxP9K8KGSofDW0bhLkmnnWOlJse9m4kFr9YG0WdF7gwHVIhgFq4J
94jgH2iguuv4DTlxhnm0Qkw+c51KrhavkR3pZw82mqSKret1ea6DA4Cj6XGsWwoc
qnmRCt1vEbWJatMF6xU9hjX0OTDv8RUVQtlrVkqAh5N2gk+X8bLtdsoq+wxVq33A
jtWwZ8uXZbpaefEAM9OFwfAsfnaCP4zBkmxk/Ns36GQxPIIBbr9h1tnH5++fjsaB
7xbXSygeQZbZFCQ2q0k3v+0pt2Jic2FYLKVrdgD3UCer+ibov5ybtS6cVKrycAeV
YTcamoXj8d89pd2JzZHcc0qCXLPwRaCuiXrrdmYCCdsIxpaBmqqsfYSX/aBPcaIa
meW8xj97Er5dyudxIbEfpwgqP/Wlnm4Gbb4ux/dhVoVgKC24KRogO2kDugolu33w
T2aw7h7onzMwMh9dmDxeps+dc2/qvEB3p+8xizFUf9jgYWavnDjJ6NW+3orDll9e
uU3KqFl4IHD7kxoh0g7lZ+N+v5/n34CtyLvhpdS9lJNdWQfitf/glZnXkwtSJKH6
Dm56ePIX00QvCs+0XFcGUu6NEIlfJMWoy1b5HoJjwM7Abt/MXeXy1H0A35cwckdt
9iVUL1X6oDjrTApcPkcpwRcFA9bh88SKayOJxAdR0+mOJfQnD9xXpiNXyiw9nQ1j
Zcu3jS80aHToTkDXGgg1W+EANv6ylEThQ0cfl9YFFXqIG++QvqVj9nfJX8111JSQ
5cycY7r0/9FDljOuY5pnJ9fhBUU5GJKa5M8J3UupiBjbwl5myYqMDmnyYEG8KlhD
b3hWGEVX7a05zPfazwT7zgdWD57UzIU+avAtdKLAyheb6ERCgob49HwDWLgaxMd4
GjUYkFgf6/+vAm43x5XEqR89/ci8M3BziMAKt3szvpIAlBazzyuuDNuQbf1Mb1SB
aF9eyf3WEWYoCiSju4+RGGTLFKMZfTyQZybuokyonsZgbOX9nfQIrBymXHkQ7LtV
+vYyflRqyeeuEsBWELE/UZicadtw2DFQ38/592DYYw+4DLFwX0BPLn2d7ZKWwp6V
jb9F5K9Fv4y1IDFMVspsVg6/dd1jvK40hP8ssZLLIrQHI2BL4kdYuaJQLqvM7bZM
wvDatzIHGfA9eYY++2fDDVhcEbRFzhhddwZOVvTBIymgwU962e2NYCQPvVWPDkvY
E6DHAOHvbcog1koVZI2hJOqs4wv9BMyhi3pr8Z3oNjktEibY/dYfbcwAAfTRY3wc
gt7wFKbXQdnn8/Bi6ke+QhHLa3Y9JIz4EsrlsDuDyerp6GU49VBvCFiqrYKixc05
fAGtWEPpKynCelcCd4Z9UoCOT744w+xUNexpZ8XiGVPum9XiA+pSkmRk4eB8yF3s
qJUNuKNYFSPy7ZWHooqa/Fpp0/GMBlOjw2zHRB3IqJ9pgpF/cE1hS1MSm/hji8kW
ZkwMnb5f8jmnSWfC/UhfI/Oqjs+f/z17VTBpuoP1DIIc8K6b/Vrk2Bs2C+PMCISU
/3ZaMnLOPANd0muQgvXSPCt7UZndZ3KTqoJkRtKfYDGo3cdmDTf7d6aQCX2QyFIJ
2UE8X/K8RbPow3yP6msjGc7RbMTDfWYWcA5Hpj00w5JC663PRDnDTKMTG+ov8Rbj
SQv2+DArdOzA0mnYjYnE5tKqPO/nFp+2f5aTHjX73ejjl/PyezLQ3uzUooo6DsyQ
6gWaADhApZJXBqRTh8ZUfOfAMN9bS+ohNrKDav2LxZ5+UVLraLhkjYcUt7L/HAcm
rfo0PfcmpUzkfgumYJkFKiX9fSoNnoe/794/cS956YBPzRjWX07KsmiPmw1gcWxW
14NM6Z4adwb2HEuCYhLBjvhGTikmzLMny3Hc02Qubu0MJePE8ctxwkkYq8goMv1s
M4NKvD9Z7AK5japHhl+7UavKTsVwrIRNDVzC3YpWIgkw9z9EgI3e3JlohBKdQhaH
f28jV9vjbIBurABergTj4U5SVxKMd9An5XAN0EVlonYwDGFqFUNThmme19aGlsTL
DF7UR3ExmK7ggJgsNKbYurT1q96j6gr4KdeumvANkVBSfTXxdSEEYVi28l+2Mm2J
fh1s7iPN/o8FhejJdKApnOscDJ4/mSB074JrexhB5YhrGzF1mUXyvMBXwZzsYJyO
06QsPV929vR8+cC5ywFn9els6CZyikcTZYm0CSm4q2wYBEH1iLD2L/RNizHfE842
RIE8d3jELWQ53avno0vrBA==
`protect END_PROTECTED
