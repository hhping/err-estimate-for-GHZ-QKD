`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsd+MUukS7Bs+BvibpOL9x0dO7TgkZfdc4qPW8HmAsnuqaOb8/sh3w+oHnVZR9ab
IllsWDEOdLLnCUt/IB9VlCg1TDbBZDyisSgP1YhBUMCbkXTyIpqvgtUcriyhXBNW
jHCHCApVX47B7euEKE+ytx8DH8GRO4qVkLzqY0IFYTiIrlHHeEMJazpty5PWXUA8
dfcIZLzvI9BTJM5fJ1mHJwR78mWjEZtj1/WJmRaVKC0cMnWzCoOg/wMH0DtVYhJe
B5tdHaJpsBBd3rWvuGnx72S/7XvT4CctCxAPzzC0JdHTqz8FpwuGFzxtwHH+YxEa
CyG3cjJ+kMKqwrsxaPTw+cWAQv7SrDzsnUXhestNWuRjZZVwjf7GJKZQ5GG90kGX
aDz4vTQjwvKeP1YG7CimvwZ5ZcQYbhkyA0/fOBVRTvb1bDx5E4sX8/g7aP1kPQ//
wn4Gsgck/X2obnMSueOd6o4iI6wjhUGEXXT/A09MOSD2Dm+hVkhBaNq6fpiY0NdH
c14Su40NTEt9/8MlPbQtsKF+4yDvrqUr990n41P+UEb3r5ymr4RfmqYMlbfsGb3K
Yn60/c2iMWyvpY9yY4gOgIiZF48x9V1szkv2hlGZgMLC9tI3sVUsAYSsUrJRNAoq
96exbb5E49oTSma2QehuapUYOcs8SrZFfHtKMzmT1rdzC+bx66bvH/XsCqf+mBYN
LaexukRXkZm4Pb8oHqh9HsMLjBkOeB7Kscenj8h+ylogGJS9SJ2a+JVMEZW5a5Ce
P3VePhHepgu1B1fq3M3vU9Weo4M29AUyy0OYJrIcURJRVt8m3TQfeJgYnopCjIuW
xWRPsmCCZUHc+OL3Q7nys6v+DkWHxAUt3qarJXR3xGPYdKEXrN5LmH6KN6fOWigO
kiQL1e0n2KRK+nlvYpJwLCbt/kKiifN4ydrBKnNwcWteOca0lLve14H6PiauJkt1
4xCyXq9bn6hj5vTCzufaYxljtSaHC2+vluq11vbUlGRIrhACOz+4G94I1c4RBFJ+
vbHOj2BWQ8XF3voC3qpKzODvkD3r2FYDByCOd0CUnKPs0V+Xo4dsFUMxFvUxsYEs
V0EDXGGadqwSqhJN2g0C48VgFgzkz37HMpLxbKQkTUNow7SX7KDHfmgtncvTw3II
PmK0Tb+E8+Aay/hIegBeOzLJ64H/B544odh8m+9zV1JJRZMkVznZyGh5HuFK88t0
K+6Ml7VxvBFfsSDK1BJS+Ps6T9QQhPXDAOO5M3YF1vTV+lgNkrv0+4gQrALcxoB4
`protect END_PROTECTED
