`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
715GTT3vrsMwLEsQhus2+dLaadKk/RcgrNbYcXKym8RL1Gv2BPqDEDQXDg6XXXwY
foPm04SPJBDUr1NdfY9RbQqywfZZtWkL6x7Cq9PYn4B58cXG2IpdoRGOw6c3dXx/
5GEvufAkARhf7Q266g7Dd2+l+jRTV+0rDdeS4p7dBJzHEJYjMAYeFYKwqDs/8AZe
YUuUFL6m6NUbGCgYR1l4+XNEEnxeDz/jbK3ShMgj2hocUMeT8nln6F1r6xGvDqN6
SKbSTV6F4KIOCPb7wXgIujFssBERvu+Y0BzIpQ/isZDFDxfWuMEmSM0Ui2XDKZje
US0BTMNQH2+3jgHYxGopDXwZN7DxtZZyDPM4GaeItJ4MkAcY5gncbMIM35BNrjvE
4xpweESoHWbKZsvy4mhhuNmd829EwDNYnJtdpk8GKev39DkOqNgNXYMShm+WzfjH
YOiE6yb6JFpnRN9Rk3wjXYkrxe6hTBOSIxCHvWJZNMs1+8a+adDTFevCG0ymtwXI
wsfOOsyY8kwboTbxntlxk/cN2Qv8ZBEKe4xDyWypPh7cH+Dn9lUMcQCksjtxXSN/
/lkxIzOIbXpOwR4j5bqZo//4QiOWfhOY0nr8+ivVraI0OjFvu+CH2Lzgosu29tHI
Tu+QZQTy277mgbgR6l345ehu5xSXwZejdd/2wRoreJXX8sAa4QvPJNg1T3nKz0Dw
erZCH1TFWOz0OeUu5tHAGQGxKKgMgh7Nmfe5mwtWUBrVf/gJQfsqMElH3sS1L0yp
XCBHNRU8v/dLhDbAXpDL35TCO2ZZuysnBK58N8jyF1H+R8+Z1DHEP0UxM5eKpXxQ
aBDvgktC6gIpYIxoO9ZSWPcBKJwyiyY6xdZsCO+C3E/PTVmEpkJtooKbnjRTrTiZ
LZTRjV/HHD7ZvEdS0XnW4J3Ne+kHaDlE+3HueF5iKqQRCvfYAmDA9RaadHaxBrMq
QNQ1CYU8dljzm1yAZdEy0tKFBO2yL/aq9J1jRhWKc38ZIcCT9TZ5mr3PHqjvWjXH
kC2FelvIWU92CPie0kaqRXw+Qus9DiVbCxizT3hJQ7w7Mezq6m1z1H3wb7vG7E+U
iugUeN5PmShz1zA3weRG6hcXkDRG6tQ3iodepcRFNSulSQ/r8IcAMPet/wyC+3cH
sn5cZ8/dbNwQL7NIL3iT/geRHzpj4zObk7oNMMQ+iPwDOFYUG3aGw/erxPdVEpbS
MKLv3uK9kiXO9rblOrMb84UOrYbFyVCEAHx31mJlgLGbg5nF3JmjLxbMKMV8jA5R
QTObY66LZn6IAv5SBbv6C23HQaKE/D2PtK84mieQ9p265cWFSpmsVLhGrz9Ef+KV
oJMtCcMSAUTDKg+le6FtqvosXJti3XxWDJvuQi1BbCKRKV8wNuoqKxXr6FV2yQNK
B0n7Bk340vKPgFttKBGs9eBzIBVLuba5LqVJBGd3bwX1BfVpFUB/s+0Mv9sWkjBS
0n8/zKPeMhF3zNOUc9QU8dGRXERsr8+X2qDimZUS0zg5VSs01z6ymKx2xlSb2khv
yrHynDJkSlQhstX0/pb7nQ==
`protect END_PROTECTED
