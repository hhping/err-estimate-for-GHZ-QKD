`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfPSMFkwoMUzQYeRINTQmpvtG/HqZh7VbvbYuBMXkpi5D5bW8X4ft0n3s71IMmnx
i210q5uB1hUwHeu1EphrVb7wiZYlyWhQNAoCuSNodOKkd4EiThXrVUOAhm+BVMW9
MsJPdpcDBB32j3yQ0h1MPnD8YHkKMXDcb54hUnM+zQnix8fFcWqzcmwGp1A4OJie
dRkYVBmK71ymTrW+qOJHzK+8oz+YLXhK3qjnEVFPSdG8SfB4I/4ksEZTeSPCxQHv
dPR2XMqpqKd3YqGFSHNt2HMbw2jHj2UXy7pttLPmRB6NF6jD1+2hhvGZlV0lkbkn
f0XQqkioAu0t3WUOb0dumOarU2+Ff0OYkK6hlpUpf90OndLepZoPPDigsNJRSKZu
/up6Tawq/m+YDAXJiMLb0kWMVYWxoB5ASvGfxumeuT2vizklxFHIkhC74tY3JSTu
Fa4bN/d0JiU4ld3SHF/0jgRD19u1I1orkkO1NB+BygqdLIApeOIJn5Kr3T6oslbO
MdOuYyjOTbPY8e+bQrKF6RGZtCWz0a4OC1yscm4xrbFKjD4Qs++3M75f/PNhzJ6p
FBVThPRUaBD07zTqPXKQmqtITbEoehYcr2P2VoIwNNI=
`protect END_PROTECTED
