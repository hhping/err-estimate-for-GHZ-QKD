`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16QyOoIW0l3PjqIB8JFMVjR+GfQfCA2aKZNKrEL9lAfOmykvthutWhAHVVp+2hIl
QzRVtL/t4/43NBQm+wia+pKDTR9hzAcvZjcbnxj8yXh+sQwUlqTLeOxPFqFF8baO
nW/L77zL2jNCEaXPYZ4W0zP3qffZe30RHuU903ttD5+cEScs839QwEhV3NSO7gjb
HKYx7Rdx9yqG0iexzEKyPMeLKe31n4k0Q6/osMkPZ5ko+mt4hUaOkAZGQTmKeX3t
4JRLYQNeeRu1lmDNSe6bF2Mv+pyZbgIflvZqoDYDPrF2zntTyCavG2k6CrDCd7Hy
7ulpGpoiXDF7jh/DZU01AiB6CVsUwz6Fb6397wUjZwJeuBdnQqK5dc3xqTUUVhzc
vO+NaLJvngYMm/QW8TNVSJyOlvA8iXDJ/bN7IQGfhUMXH2Hhh+6ccsqb5fd2jSOF
8NNKRCI9ag4RWetg6IweIn68a3l5GbE8SI0dSv8FClOPkNOVdDih6JQc8+lHhz/B
k/IbolFf34BL4wRPjT0IJdc4v3KZHdpOhXwfIitTh0N34ViyhqDxy84IawGX5XXV
gGesz0zp0xNlgTSIkwuOUqFF3polwEN5lbQypzYHMtiOubCFsjohAHsFcJq0LksP
8HA4KOfWU/zklcBlFizn9Kt1sIOlogwfkaPkQhnxHFhQ3Phwsv5mqfoovDTj/EMn
DPVfpuktrTdj+JFbbs/NOvD6aLfiQ2uEMBmKX2lt3na4VJWTpxZjz8uxFL34ny2r
8tqwZitcEGlN2VgxyRCoqZNHcKGPUJ1Dvwa73PTKh9ZKMG27/tuZZUuCKnTrM80p
oCXrR+HX7zRTYnPjo3MTAnyCVZ41+j0yCq9dlSe0wYNaQ248/LIbZcqQYpwWLkQx
Fy8dbyxeZBM6ya08FH7XQ4p+JdbFfKs8k/gXz8b7I887xEOjNp+3+PFhopCVe5tT
CCKSDsSuB/227tcAbhCTfEJjgCZUO9gqstdB6iZExIJvSNniTy3upNRadpGz88ho
IBVFvc2fI3Acg6RCIuq2CVuCPRR6CdqYwF3gYP6Jk6tJl0WnEp4Elr7UcBZXjplD
lx23U+g1B/OYEXFFir+ugV7fSh7JdwrejDuYfZpSWi+pKVo+UggUmp5ztMelXEOE
XS/kVyCqaR5ZV0zUp4awSMlDbfg/+aA7rPne63MDG+dyBi5aArV0i9aYQBlBwAm0
qEET0RhqE87VWO7x4d4g/zWgjmkjR63Gvx2bqK4dg3yYX12AwSkWJuycmAOgLUca
yfyaYQ3jBpXEWOjRfXt8Uam6o6wvPXHdnP/2bHcKftd2FYuJtP7QMVHGSv512fXa
gOfG+R4k0DT+tIuyfOoZSsh5ijghhg/mStECCZCAzP7sQLH4UxHU3tWwgETRZJCc
eZfhw0+SFKGVOUyGSVPgA+E6krujx/xzYCYg/j2h207+OJVSAXxoVLZ0eOgmQ29G
xamnfFv5nsez4/1Virr032fv9W63fPsT59W+NYXN/4o61abWiVYlunjeWmKPez2y
d6mBpL3vyblhpD2gpeXlZ2h/HhAiF36xdX25ntoqb7sNQoBqo+Z14+DJ4GpBowyX
T67wzT6cdEg9VzC78npd8bZaDzEzEUfAVlvUnZHYvK+PxPz+ROWYwGYT45YI8E0v
6OMwey8xRZ1L7PClYIgO64agilZ21Pa+1rotNWnU4Mqnshwz1CuOBhaiDxqTx9ex
YXur4Cy9sDTHJSPuLoRhaPkQPmbxX87TuLlvi207HvmUemPq1ZYP+uJn1IWo/O41
7bNpk4czLSqLqpFumdWXlzODm35YoGk8174zOFVuKyKypv0SZ5+rApIXMDqCrRsL
MrlloecISBZm4ORRI8WRhWp1IAnkALWiB7Gss14EMExix1msujkYaZMHV/fcurKL
ynFkgEFCfGmaAYZVPb+97Vh+vKTs+Y/Q+PTcCsjO+uNTTQDCxPl4J9UueF4fKitI
Z0bEgZdiXtcOPo/eLbIieoIVNqhUhNe+VsnkmaUkA163Q+hIKL8/TO3ClCZiAycI
nJsflP0BxTxgGVyyJb2fkSHSTqoR/gz+a206ljh+qM96gV+P9YgTDIimDFZd+gzs
j96mwdjkcN6xZ3DxfFszmMytxCPfjARa4mop/DF/2j6q3KtIwaaD7GFjXzLS4dO4
vB5vq5Lv7JhncYX9uCHJjmEscHQGC3YDhbtU/Sn+ZMOI9pKaNnW/OWnnNfnmDWZ7
KGj+i9Syls3ae8+d24bbus06GJV4PjTjjPrEX52dC4MgJExktImwcAN+27UgteuB
wtZmUCG0DP0uzwMnPwi1DFC21zr+dmYsx+8Hq7ia7nFmDBzGfqQR7XfjpVv8Sea/
XkLmk2Gq80xbE6FLUOxkN/2jJzN57satY32ItCpxNHK49QuXyFONsPuCngNwXmbj
Hng68JvOlCcXc7nNOl4GV22MPBl2hbEm1RuyVsukfXBFt2N7Ar6H1K1PqJ2AxneF
/XF+tR0Gfh+sH2us1nf5O3NtIiYLOPP8nNu1np1riZhgy8U4GlrZgAF/YeioMPSr
wLN8fYN73uwVKiESG7sGhoyLXUKCsBrpfZWdX12rR8vsnOUbTydEO81FjMnVOiJm
ov+YEJPs3e0mCo86Qd228JxPrQs7BBNyVDnngDyH8qqpSd7AzLKrYxVv3EwFVdeI
TMwsvb1wVazWk8XOTddK6xCMzVW47H+UxgMw4diOJOY0ScQumMJXd8CiaNzmlXL/
9hoIkH+U7PcBJak9tpNAcf3Uo7o0W0b2HXwxyvqPnCyB2tU+MpA4u4atMHst8Hot
a1C6Kia9DTlNQfVn1ZXxEM35AacgwLHR1Ia0sUHrNifK3H8EGOtoG93g+N98iboZ
OSxAiu2clH2MXgssS0fVo8uz7wBBu28bOzTedUci+RwvBS7gPcu2W3uZtEN1PV1u
Vzwa5eQxXoet4hGSLkv8shQyhLsz6IlSej/OhPOj0gGVYM4OvuVU+AlPUSQw2gDp
tFmbENYa3xkLk+kJQzCj8lqf9DTZJKK1YAjRAJ9YokxDa3lvjnd2LryrixG9Hzrt
opEEgeHX/VbZldRdAV+QppYiwmDG4FT5UHtZ5FYpJyHcqJKjUZrPhyYZv+cf2oSq
iUPA75q/lMapa5UMchPYftfov5PMmZHnzEDWXdAt43aoHcQfhgWUMXQngV9fJrIm
e+tw4VUT5ye93xNSjZcE6pXsDyQgIq88O15nKByKIEa+iqPcQYCsWl+Ttt0PaYtG
obd0NJaej8oFBTxNEJ3MzHdWVdxA04MuOL/MfW2Np7U4y1OOOeLRJOc/V2xWhLoA
Ts072V5kpMByDvELmBiiZJ4xmQ7E37FHchb3x/cqoTys6zUsuiO3ykHHOldKneqw
QFRqd6SKM5yJg4jzAhtrebFEay754GmjlEo4B2xZqNW+SatNMzqG5w9O6W54C1Xu
oMLkGlEMHdP7GVDirG4wwaJh9wXLgTeF63qQTBWRN6GQL7Vx9EPuopLmnVaioK0g
94i37fY8Igbcw5a2l9vzUwQU8M3DYYKEpMcxHI9vHtyWbnu2yGiduxJKeDI4tnUq
fWzD2gubcIQoSeDHRD/0LDLYCpFtugu+6sIV6lvTBDhISPZD1gfnZ+OLUijXeWb9
n0nDmDUy/K8nW92bmno4NV29wWMTeAjFvZ7oHFeLJOi8B91kWEyl7+/7f1O1+e7k
l/8RMrbRLKeqyo7h/8Gu6FD8W1F+FzO4HC1ldAtEbLqBDdVoWou/RCepT2Iy5W49
O5bZvP97Q4DvuGbzIWL/JIfJMwQztIGi43UQW8WP/4GzVUx+IVwUspFIMF5PutgU
nQzr/Xgyz+G+F9foDctBieXzq+xAve5yJKIhizHU1vUjLC5oiDO18iQg768HHaN6
cxBqJrFa4cz8Q5WtUKvbL9aBbXbH4K1S1jA4Rvvmb3LpH/GRWvutoECFT3l5RLgE
r+4p07ofo7MFK3vL73V5JolasXniqyAngp7XLAXxdKY=
`protect END_PROTECTED
