`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dlwt2NK66P13V1qylXzKJ/1SJQgNBwfAAYeeG1a580jeoJBqlbjxMHOxUAPuaWKc
fa5jAcz05+xDrOUAJMiTPk06wpthlQ0TiIpTJatQJa8XSAP4GUo762X6OF/OEQzP
vqFURuZCsHzMCAk6im5CXhTfykLJenTEqgPSO3haf0b7VA4RlbWlOcIR9unq8Fzx
aDDKgsexuf/UHSVei9Z5VGAYu+B3Y7LOS14IUes0WABHlepoPRC08E1MdNO3QVRy
iJqsnwun1wTqEfidjYf7oSE60KW3yXzgeyDZkTO2qUEndwcgMd4oXYERkJGOTgc6
`protect END_PROTECTED
