`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsW/P5+j6Dc3tZk1ObvpbkAEEUUDqZ18T1c0oNB4qxo9Vfu6FdE7cVw5MVzn8D8I
T80uo4S+q0uTswvg9nEWxvjO0KaacX37c1PRQZ+J3QeUa9zD6HQY+1Ailh0Y4SKv
HOySKut6Q5vHX8qHVjjjt8iYyTkK8IyEq5dPVoMxjd1McgD4SVxZxJY6eMETgshY
xBbTgAZIS3o+70zEd8YlDE7Wx39zFCkyWTkbql/7bBn7W489Z1I7WIAsLGVRfSPE
t8pgjyRRz82kYtWz+qLPJJA4KMsu3eiF1qwWVoMgjYB5boKZfCF0skFb9TVRJkCT
emCC0CLjcIgvDSoKo+o2VOBmiVLv+3iW/UNu3q1em6TVPMiZaAkaTfPgPCbrioGj
i5VV4MZcSeBDftQpDdVk1moyIrd9u03A7/HLkKnxY5PZPwLV7AzV+INzRJReBM6B
siGuKC+ChwCuD9dK/8xmcR46Z4D2klwAjZsG7MoFIO2MzGwG70I9WRSsvbkPtc3N
K0FsW6VY8urshJ7vtzsUSklthoS3J4aqrNeH8p/2LM5hBYLFdzvHUijWqN4u0C0+
U3hXCOaqO+vO6ogoadzR8dHvQ2ZulNgzIXi8yfIaKk9qkT1tz1qa+tW0v8bhS4kC
2JUkz9o1LsnwO3wzWPpKbrL53LdL55uTeekfci+MPN4tVNra22anhAmrTdLJW6pe
oXGiGHnhk0u0VVAz9ysHVYqR2VJyeLWawkaAf7wqZYzFyxoXRyP0AgdgD77zaX2E
5nhCe9dkHGLunqGUZ6GXEfg/FjIfcDdjf0iHkN8xYv6NLyOHHJ+o6TqtFTCOh9B5
c2h5N2aO6Y511ucZ0ID6//nr7Mj23McHgBHWrdjV+MkgCkXL4Lw0pe+CMw6bkYxm
wAawe7UfwTV1FTKtUvlGHZuiDIrEah8aVBYBDi2jAPTaIRul9DuQB1C6cAskBnvY
b3Cc0ceKAgbX1X7pW9an4Q==
`protect END_PROTECTED
