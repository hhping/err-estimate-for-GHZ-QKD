`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6kwxBcDaJdwREBoa3skJFOLkzMDCqZMxLN/9P1mSYIrWmhWCBMKVdelmXHCMGel8
gfNqR7dRlenZz9UP6HfbxMWix/zFFSkRsz5ThEwbJRAxBcNP+UCygvPodChKox0b
vSINhHQBi7uYvvBasjPODSSPIwBlYX7u1fMal6rbc5RHxbFg0V2ounEl264kR0lI
o7jd3riBKPXvmMffDFNUEzgESF6lqeMSNBa72FiAOQNVFsS2kSknPh/74f44t2Fv
caab0vT6uSWPV3y2jZuiGpUl2kMg3EMAIo37ocu4nhgYsRxuFcijapI6t4UsWET+
wTAtAKyOlnbs1Mp9dPG1jiINlBpu9vO37/IIvI6y/Q3ha1/KcPXjoz4V7qEP/jmJ
1yzZaWTQQgwpQgNiNUr0NdwhfYgbGIrRinVeOBBoo+u77ZtLRfM4sbZ9CEEkcT06
uFz+Ghx7/4zmvaniju972kcKlIoWi616x4hrViRqSZ4n2/1qtRzFvzicrUXvS7nQ
Zq0SovQsnEihVmocGLSF0xwnHHMQbYO8+6bav9g/GPHUu8d2oqs6Smij7Vk0Ir80
s4hb8in0spYiC4Jr1WdHRr+Ufb1tEZXBievjk1Pm9hxGnQIS6WuxN+e0/BdLYue8
K9XcD9eXcqA7QdipGT7bccYDB+zq4zqKrBJ7/CqsxXCZ2tXhDeBahCkcP5n680g6
gmwqQtnfX42akypvzJx0dbAU1QMFLYOuQseIta/ihxTR0xxVBUcWtETXN6J/aYpv
atQhKLDRWT9AieOm+imNNT4Lg6WZJBcpwFE1gEmt3w0w8jHgnaJXTEnBkJguD8/b
UzmReSQG1ziYsPReFDf9+51DD+2/ZfJXtsyRX6Cmz3prqBUOfNM+hooDB+1hoJDr
uz35MJ9XTnEGeAufMyf/LEeYRU4kS2u7s4XYpVvEi5D1Ff86BC7mVcy3SDwZwY+8
nxfWU7gmCICqaY4CZTYJ4AT4SWQvnG0DIqyZReUiyiTvLCMhr6EBFRAJPoTG096R
V70S6N65h/XMVrQzdmab9ry4RHsCrU3eGWlxTx8XsDy5aCayKGhpXZ6clSaILZzf
5uceuogzfSKATNLUWrtDyKpXsxh6sqL13bMZ288fs8jpAVileD8DZiw4KYclPIvR
o+PaSn+AmXk0TcRLnVe4hOAUgea1P6D4ysHBHz7Zcl1qP6IAzYVlpkGAk3w2mVF0
Pd6jSHiUb9cxMlUy2POJfg+SdZheGD2o1ZrKc+bMGZA=
`protect END_PROTECTED
