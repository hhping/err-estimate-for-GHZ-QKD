`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZZBhmZb8FHnJRhGE4u9uqos+GnQs6w7408R42GGQj34UevSWRYMZwJ9B3f4np0LE
9F6yz9nDtGOguQ3eMZnAKUEBRggamV04rH3j2NcYBCVh+IhNOCQWx8VYCOX96xNT
I31ck5sdsQZjlw8fX00BLoEegYWh12z6YgEcPH1VYMeJGvxSNBr6v/j3tJz+9piT
J82Zso0oqd8PrUgg+loD//ga+6x+XoLd5Qtp1T+NCPaFl65Ku3g3Tz4+e88z9ZOF
OcHaGud1abjv6mkIXqa802GWpxkmc/6Fsp3tek1ghGJ9Y8zOJZeq/fGUdF9xbUqM
GSe9YPqCrbPhOZD+z0GM9KhfAyby89AtJD75INAC3ntBbWAo8FpOuvKc2BCwOIE4
Gydp6yM0N+NWQRfE2tpe1rq3+iIEOuE/RmxfUjyeF+jkHXWplWwtnXiLRBnLGoG6
gbjpqXUg8aTNM6v3+Xxsi3czjnifjP58/NA1Y8hSNJzrCuxKymUZYrtvGarMXt3o
xTQYJv8rMTyAeY+L3y+Ql9c67rIwxFQHN8skM5d5tXPYBLdruhZFsG5VgsCBYxOM
ioJnQY/HzBwSWvKgQQyCu9NtFO8tR6nTY7PRODqhIxY5vQ2tmCFMc6X0aFqPE55x
X1qs2j5W+2LKxWCmVGcklNq4oZCVQG1Pcw84GOS4aopdPYtC5dX+mmzHV/DyUbab
VJ//CY6kQOyOko6dLk9CZVamWdtIYIhvxQ3jB6HWG0/1LhSc3M9ShS3AaeQWi2Kw
VnhSGoICJg70XvVMS9kuxXdihd+eTB6jfHBIDIDSxm3sqjw7XsLwsSfkkQSFXz1/
rjhXb9cVDMqAf1dHgLYGQH5VwzB0JTxXUMVEr2R/QzAdkt0TVDvz8F+KOacQsCKt
IN1OUArEQ7ZZS4zvHv2JEeB8TuRh/4iFGPmYHOqpAcNv3Y79V46xLMVTx8bs4K89
emnG4K9LE3btYzYrdHEmYji+pCrz+/wwICLPF5zoeLPdv5J5QtYJk9trKXGkL1v2
ZlotWPdJPn4Zr81/DOFjZsBQa1hI60ugYnEqCPoKYEgco6NcDc7QB0F7PIj0fbDk
DlqTbSU62Fa5EU9H8snWbyGlo8HYXcoknAVJDHiMpBrmAQlQtEOLKDim4pFcDs2E
bCzpxfeebnsQr3VWoUk6jRHTGXINO96DkOVub42waeu/86KXMHNcVH7w0RnIVeRw
eYjocMAtylkB1u097MI4zoVeq/Zlf/jwRaTUYj7jekAFIUK9ORFA2o9EPsB4Nagk
e8UjCX747MAuaqCRkhC/CJxbw4V/6ZxYUQNf7PFbYsBBjsg8O19OSYZJVGQtLMna
35FQbElN+KZygFAOcOqxiVBcS9eDGIts08gJcfB5Z6E7rBm7nKvyXmukrofOzDjq
KvLZJPuQKz/zfc8/MbfPvFqHxdDisy9bXquD4gER13xk6WNoajV4m13BQRiec3mX
Qg9cOotX197jqwNr+kT8tOyTH2ditCFIkfJdtoO2Zp4YgtyVfA3LHsugtIPR8h9v
C0ka1nEqsMG3CmVwqRdYrkm6j9AdTwgtgcAlwxNYIfDaHaor8dssK2gVM0j2+VUr
4aQ3epB5C+TBdtShXJGS8t5hdWtTQTUK3TM5prsbHxxV4JpJWPXOBoo3rxlPRpaP
tJiAcjTO9shQFAC/KNCBG/IEBPtEsH5ovLL0JuMf5v0lWpihjEFMIM5engKnbCNi
+AYWrjYr/KYVAWJ7y7TPsvZTYV/joae5h9HXcZI6Hnzbmj7IEXqrsuD8HuQFyS3I
yzQRscmYJd2nqw0SQD/XZO0sX9P6xmk6oe5cHBjmKHuhTOJhLtNdDMrygWw2+50Q
C4n70PktzaFYcvMH69DQVyPJfYH9Ral/K/JNzacqFRtLDw7lZHR6bl7WH8pcYwv1
kaZVY/0LnLm7WOYs57GtzVShFYhGeWVeFduDS56dGWAyN78R87FWHrEFsy6YDcaY
HFctFCqfmPKd1QEBox9A7+ecQ3jW2iG1OXf87zf/5sfbP8iu1VsE8s7i5yVeJ3Oo
0BzAQExpj66awutgcjAW4OOJ5x4N2kYDZHZXrGVurDijc45zwU68h1gP5vlHVsaN
G16QPjDFS+0VcFhZnRXbCz7+TkVeUwD0U5tP6DRH4DaFly00ydoc/MN/Qt0glJ0w
faX1tYaCWsRQRtmESjNWBAbMIl0hQRl/gJBXBQLcJRtVywSmPb2dnO4LpUsNdxQy
ErVII25U+zMMBqJRD6qJ7trRu0VgVyDs1mHcYXWEmZ+KjIV+d5k5MpwLsOwRtbE8
JXhR7+/U/ydn083BiUkUw2jnOgis4noPtmAuL8RooVcZqFBTv/t+eWbJx0QRYJ8P
0FYfreCnpya6cwa5Eu9Fc51K4hKx3s3NMmDANC6FxVfi9ieqVsiKYLIy2PZaChAY
K4TxUczlLdWRl7cq8GcubzErtd8L+PupgCwCyDvWtAY0ANsssCYhQ0JrCFk/4M51
+osWH+Q57WnVMvHpoedTwtKeoB9Ub615baOUXi+yLhy3ZrSvE+Lh6ejjXczdfZgq
LkPrkscWYGNusyXqBvtYEi5mhsKew/e0ZwMCWdEALcP5HlYuHWJgATIi6hprzLon
0GXFh7n73ghxO0qNbpt9UaqJFwFcdUByTTV7eB9JLcvJ1XizkS7ZtYFmMN6PndJW
ajra7y8vCAk3Vh9nHtvvU5S4ae/u84Ed3gJ0XYjCUTKMeluaM6q3lCwc/6YTww5R
3umXnq7tghJ5U4pgqloKSJHVElNVo3EqZkWTtuSbFOHs7MyGdsqQLMd/2C0QEAuE
HyRm2UEiq434Dxa40Q51LhHX9WX9Acr6RftG1U2Rpg+ZbR5saCFww4u4/EG5EFdE
fS4vFmtbqm3+mGdpFCY7nvxrWRJFSekTAYWUrJYzC4D5P0D4rngX4Iabs2Lhnhu5
57HhqwguvSb4v04z2en39lXkSV0jxj6UzcehlVP0wjo4iD7Kz+DdZe7C5zusETAu
SwiiTiMECKuxsDrj3GwTjhvwKhohJhy+ZXzinO+MRh+nUYZkJqKf1T4u9O6m/jr7
fY2IwLu9UKb6xwPYFbdMOVXL/vNGMwIlCb3R7U03R1k0j9i8Pm+IqknyG2zSp6dG
/61ZOZfMmfBFBBj9t5Wc4P9pCNFkm2zSpNIZK3ZNxwDW7bl5rth5mt4hAXXsphwD
`protect END_PROTECTED
