`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hSIdIOlVGZ47kDcFMjqxnXrj8tfX+pbYA2jE+13dnBNreoCi5z6J4iuGK8drr6tg
GMGrJCLu9s9BCkNpFhVL03ryk75xpjSTEbXhLXcWKUhKItSNmgNrNeD3J6CdRb3C
0lZ2hURNqIY+Ua69hJ+RfsfNxhIKSEIjPDc8j0jsO2aMXADQR7zzDioR8RnE5Q8B
VnLTfV5OW4GTYh7bgzcb+e4hCiqw5Y3RwjlTB9gqpa3Hse5BXuxAIDPgjkrCsoDn
c+fG3fdzKjLtJ/dSE4jHAjSvxImyFEpGY997HlCN0hFKPs1EkMJMeRlX2lA4JLz2
gx/aE55i3vCpxcCI8wN1GNWxnJSkzPCIl7WKGSDHQ3Ckhcn2lU4t5Z90KEzt9I1Q
DzHgb/otyM3uBG0Vk+msW3oUixeJJzJYyplwxAMa2KkSxnlfNqSAfVEuHu2z+Rzz
zFoSFX5f5MIhHOwxQkahj48/jtIgkSv46qMwChha58hhQSX580/J5SwbX/oBQecK
BDGwrG4AIAXqOcgEhQ+XcABgeNH8JnIkdwxmfo9A8nAZwAbMJD4miPfURSJLA8yK
8YViHah1dhNhmn8CewdAH5MdGRaiVOgeBUfCyj4qTiB70rXM82k240CUJNrYWsdJ
jrlQfVpO6a8EQgvZIYXNf1uuJdQxx8c+t+uUF7Kc2GaWrxL2It3brWYqsKDlQCKG
ub1P+2wNR8h3GIV/+zZTM6wETEZuB1qsuulaiVZlHswDCZ2hoEtrUS3+vgDN4S1o
vJmekP2CrHlzF/iBQi7cTdTYk1QBqAgiDs2gfUxDCF3hznrS4ImqQTglm67LC0JH
8wCdB+gtLiYDp9hUG89AGBjnf6flPZWq4y+fjbjjOHpcu51WkTpe11llhYw98jXk
tDsrNg48fkz7M52llISTLKo+PyfAaeniVuWid4w6QLuOtIwJ/YVOWkyiI8bfnH5q
H8iN2NsSlvVbpfgWfbYCnl0e8ZcZkyZxmTQt6sprzytCK83nxGf1ss3p5QM7+kPX
ydyYt/pvrovRolc0GHfWGJCE++pFE8A3Xky+BW5PZz/TguiR0950Bwa9Xp/BzDoj
7NII2PRdQAk6swV9/3b0v1/mIHJBn61X3kWy6fOiNWz2IjS7DIDS8SyG2Ce4B22n
`protect END_PROTECTED
