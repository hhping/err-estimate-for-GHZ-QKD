`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sZxr9Uycwnl1KLoRgXsmD1J1dUPR9ZboLO0ZzxZStGttWu7l6nk9UxGQY2Ja5+g9
pMo3bc10iBbGyf8uagM+8MC5f8oY1APRZw3YHJ3rsNuAXMHvkEWn+xfNE1TjqGl6
b7MMddjs0NTsH4VYX2H+9mL8ZROiad+DcvOq1RAYfZ/Ol4jssHjXooDFjfPLVYh/
VgC46IclNErL0Gma+t7KeboaHhf9RVHfnLfYojQg2CVemNGU9t0YxzBwUufSD1Pp
8pdHmz7+TAK0bp/95n93OudeBzSFWKncgKbS6vQ9LfOtFWFS7T0tO3qmc4DwJTco
yJTo6PUQCnYexe8jJZKetyoR6B5LOT9ozx8Kd46fW8sD7b/bvGobmS2VUEpsds5F
aTGRZ9WJR7d0QZVRw41gEJMNhTa8afOWGjMICx8zyB55fGUpNX+The9UMvloJ5IY
ohTGsBq6/uLuNp8FuaZ6f4CTyyvT8jd9VbY6oAMeSJJPnvTRauvB7dmuOXo5d5Id
G7Uo4MAKLONxURtj0/QFTy00ODQwfkg/hWk2VoPdcOJAoynm5ZuXJs6AN2Xpk/xx
HU9PHylX3SB41uNaW4hBS2F18XTENFkwOJZOph15FRqGTfYx4hKTqgKHXIRfauLa
nTcc22PHS0LOS4j+bzEzm9pXXz9tKKpA3E+yL7/IENJMxCLAoESQsjKM9qR2jyn9
gxgO2PhJnKGVbNIhuGavlJsyCA0fHrCWeOdf+ebuOiWoo9Qi5AgEaSy5xAVhWvG1
XLpHYe/1cB5s9iTqlyNdMpDk6ytmpiLI4rFq+zU4OPqzKuANqc6JlFDSvIZjP9LH
2grLzlYCLzeS1ihIuruAy75jkv57Rt66sq2qLE/jQT63yZpnG79sa0OBbKnF5SYW
SJ1hZak/uu/B7Tady8A0692xqgY7JfwFRg5VW1PescPGwO8flwxyinIkTW+5Dic9
H87VbQQluBDIF1so9Lj7updeprudVu+wI81xJJFdefebMxvcIDwgJn1MHWOkZUie
+XqMyG8LlVYAqmtBokZkjQtIqGc+RgN66PAREk6a0QRFHyTS1x7HGflEYjv8r9gO
YXl2FVWSjxelPN7OuKSnILg27rskNPikmtLu2poJ4Lc52jzdjAxEZzhgvykz1ZXr
+kFhhLvRSMzaacoCkMjYFrY0Gzq/znbWuKvnts+xMTI=
`protect END_PROTECTED
