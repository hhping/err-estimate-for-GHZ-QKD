`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2nrLrbqbPIU80/71dno/U+bGGBi2h+QVBKhRWNjjWD6Q6aRyELzUS/QV3XGgT7zU
izuGmZmgLNOFvy4FYNHms0SBCA6iiv/LeNJTYD3sM2wueugpyBWjtoC0kSO7Ayog
MFc0s5N9ZjyboFAh9NqKuYs2c7cTJOygmYTWXY8VvH596jCXAbj52jtqCGYFi25K
ABHTYZ5b80Epp4TvFByeBiYAqw/5e+kXzzpCNxOXGWorpnsSZa5KqVKjGaPrP2xX
mJbjFgkwXKX/u6mOJ2Pv7R8btepJQ2wuA9vJn26YqFpdxEG41yy0h6J9ZoFO3g4p
LnxbbYUI+NloGVEKNUoFIe6o2tfdUVwYaz3vVsSs0paeVVPB081sqURl2FrdBl7Y
J5EZbTB7O1CAUtVvT+Vs5f6Gntdt12uUGo1T2W0CaYCGt3glb9WbdZLLzg9o6/mZ
0tFg48E7ys7DO0lLSRvTIoNu11hBbkvSBDJyIzEX35FIEF5yM2lK3rr2nua6F8Ev
BupTLcNTHlswlXYLLhblfHNOiQ4T2rGCkWfovOZXpqM4AahX6eHNSRLxZ59sZ40b
rIISii3qbmWZMRYTt7aNS74YG2ZZC8UpZuJNbNnL9n7Z2JRds4Olr6lThGaCksu2
`protect END_PROTECTED
