`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/C25d0aIwmiDvbET1ZvL441SNPfHI611AHnDES3mu71b23AyI/j8FBSdgqE4s82V
fjAbOHRy0lbxHYJ7nDFr/1qWcYqlkTzd1EORI5p58SMLztoHTl81mG+gtWFDhN6k
l9ivi7XhmYTiO741YSwUFX2RB9H2YlC5ZpTDJ6AQgCLntaziIOXTwPiEwg1ibU9g
MUCLYl7Qvs1M3BdFhZNqpa1zlQpFnNPpk9tYi8Gc+Dbzf+J+VqS8gfsGG3XJFv+n
v/+qyAcIbXLuDhbLszeedu9eQ0RGuPGxMJBsVxmO/Kq9Kf4Gaw3mn2qaeFanQ0bk
vctXaKR6CthOlhj4NzFXH5Zafb0s/4dckMCpfcEtk2002hudC9ra4QL0VZR7yaNT
xkvDJUR2zPUIoGk4dmqmPnhlrNpKoWU9f6jHwLM92Dve5IlvP8hFlq8jH0f+QzzB
+RB6B9P66Fte6kE2uwImFacjT0UmDuG8EcMaqFQHYP108EOnUprYlAkmUhm/rkuY
l47pDo7q8YugwHHsrN3dzo2pPBUy2HETfyQ3iNGCugGBZP0vR00zNQ1DzBft2GQk
5BOLbD8JmuOtwdWuE+1F44p4B9Eb7FPJHbePwknqzM5m0tPknCDbZOo0i6bHPWXA
fF8LMDvbeCGgvtf6zXej5jw0z8V0iywRgZGd+op39Cz20qB1Nv1sRbyCapJ5/C5u
kZz4cxNgEUuHDe3lNlQyp/0/0+nbuNTpyD6B61iWDiTYHpM09ft+csTyXdVsUbMA
qjgMI7PMsR52ocym3dWXGVDrlEYeo8BjEas1unSVEjxJOb9XRg6UkPW0bLMiqVEU
gSxmV+fmB0w5JYsdLV3Z/9iRXFKjCiFVKiYUGaWIQpDL/lScBWsITHnpCbyQkUNL
7yng+XFHdLJPbemaFhwlw133ZlQ+vgQWNEtVNcWxXjg5Ix22HuLAWWtuCqmRe2bi
YiQKfV6SJqshpMfZTb2D8fzfrELu6tQ9vEliykqD+uZxRoFZdOQCTB6Np7Nq8r1j
N24uhZ/wzB1652Z0JLLGGCPaiAWZCXjaQ2nfRkUB4UBWACwVuFn6oynUv5p5iM1k
U3isQwXrwJrpdH7jMKLADg8zTwceVXDnk1FizHjMBCjYBo8/V2k54YKWl8abHGtl
TrtudIjZAfiB113P1CwxaaUT8z054gTHF8NZ80FKogvqWtVNY2VHG0w8V5d1+WD9
+rap1zc3eht5/sPY6mMNz4/Fv6Ds+IqfojJnXFJ1ynsDFEnuCBgR0NNwJRbhER5a
jaqYmD4nQK/NKNFKQg/YN6tCdSfzQpdWFh2BWVkPZWkwvl3d7OZ94zR6qhaoK95d
e64xwlp0WcQyMh2fOkpg/zVhvtNKVzz+9G6RqPc/DD3F2797taOExXBrKn46Koh2
6X0nhOW/ToRNxqNvKBDhibUaW6+px1nmsE73fmyXoLHPqNUrMWoWcFbSblJQQQD+
Z990B0TgLUE+HFjAosfOeP121RVEQrxNvWpeB0XoOy3/ZYSwHVu1MsBg0gX5Q5/e
E1uGf9betYTSrXUpgQVfEHVPiLqK9IJMwYOHuPZn8BmvTweM1SAywbEiYvMCILLM
W9xlTcge8Nmv/7PVoMtNI58c9oJDqXsV6QFwmuCcicU8j7RWW1zvtlcRI/GBxVd5
b1zfOuG1tkmc9I2d8ltT5WIPOXf4cbijXpFsEfT8PgXn3FlXOBDkT5rO6LJuFJka
6izB/VxaHMuk2qSc20Q7j09MOp0h0dKQymVu1CqXDq7Svzv/vTJb07zggEQRzD4i
m4jSdvM6WUwRK1LO6+Dmejm0PJK6QEQNYy7GBXWpo9MRBxgFmFR8nHJ0uOYGO1/S
pA5jhiF4/+wKZ9/sadiAdz6JT1yIGqr6OJxya0ijF8rpZDIFQxKV7kt+PCYFYqmR
NBOzOXRhmCFg+G57CL7g5+zMWLTBw/SLTXfT2g9mrh8aA58AkXoDeDm6ENhiBYqg
pu31BV7G8fe+vB4PzAPwICnWDRgRhOn91E9yrSv/xKJCVrtAvOZDhRcpHpWMiIGa
58TWZzrlxJEAk57QUzVkzEwGxukHifAhTPqysuodHjL/2CCFNGefzATWmkTzOYt6
ioh5QpCsmLZDJ02kpyGGFrLsn8rpJc6X4jwkbkOGu4dLrRx4diOY6JNFAvE9Weqv
eSeCmug/euYgeONtPZkK4/e4MLqW/n0tudWu9KeQfg5aXfMPLqRF22D0/MF3GP6H
rca8aD2ejF6uSyz7kOZX1vt3fC5J/8mr+/1LTCv92GaoOXYbzaYIL+kPZcehxIiS
zQFQR8nIZGp7yT0DyahQpx0qzZHIv8qSi5lBOiRzVZmze6ca1OT3DlEinI5C4/FO
qjL8tLEg8URU+WKoW7FKvfISD+rADgDX3c4WBPen827BzrA0eeK8DMfI8QdIJX/W
ouDzzAHh2eFTQplT5t/KGl4VfPYd/9cN1ojuLAXHx314x6DGLps+AbfvyXsu6iAL
oOrMgP8BQtkjMflEj9wpUQAs2bVhw1mYhCVc82NTlbeNzUo/qyNxCH+F/NV4dyjq
bkZI/uUyUBJjYC0Q5J6I/B+GmXcG7rgfgAHBMntgF8tLa6RyudiF+LRlwrA4tqhO
dOGQwMvWMD5WgXziMWWCcvdr3CYJHvmZ20ausBWDh+sG33UbFreipZrmRvcAtm0j
nF7gSWqPh/QSRqaZpiXHxCcErvl3z3S5eyYl9Xp3kOQxrmCkrNN8bIxNS2lGdAWT
lrpa/Hh29W7C3tXv/8+KOmOriPlyYpPe5Fj6/26fSJHf76zSwdyteUcd7W8cuCKI
qQFe59RUxgBL0m/tU5Hz6JRczT2XL0PFm1O7Qfhr9joqwCc1querEc81Z5TTbmYs
lv83l4DnZu0RB1fje82jojGhUY/0uQPcY4slm4VIqrnIIJsl6DyTloUvcWh3/6Sm
M/GM7VhvPstquwUlInRTyJ4St+eHjLivwudcJIl3C66zkj7L/35qRrNmabaiNaPS
o0palA0wlK0YIKF6wNEnvB7K+8qVbooBCUjAhq1bnPNmDuYoB9sFX8+KUcp+hyp7
SHtysl5DyOLrbdYRYo3B97C2mabalVYvkJwkdsfZIwLsB2h/cYEh0cbxaSmDZHzJ
bG8HZhQDmTK76chRCJHCNdsPBAGQDtxHhQWP107TovYaFtMhNxj0rQdqj+CTp18z
yiCpC1watFhc53MKbCyUPRC+pB+34ZAHjwkOF0PiSU5MDwJdObUWddqBVQa4RJYr
dIk3CZbGotlAepXsUll0u2pubkt7gsnvibfO9V2wa0r7AD0g35TRG1vJy7xpj1fN
7+vYhNEHCc9/n7CRcld3sdK6l/D5zmPCnYDSs7eflF6NG+vi42OCDhG6Ea9frXW8
c434mJ63hatgQOYy7tWK9iCsnJ7ZIFm918WkiP9AeqB+HW3ud5PaQwhxkBDZb9Rd
Slzuvo7a9wPH4GJ0WosDy75NzUAw0DZUKRnm7v44u2Yw//H6mH0dYWRzxvcdK7u3
IWcA8jjz/dND/LqK/r8RjkYMadnVi6H+wY/q2beKoom1anySfvw7ivLpZPvW1XD/
g8Qcwk1WRy4vZsAQGJw6KDosIy5LQ39vaj5XdU6uR34UKeGmWmbYdn7WAwobig/W
edglRTq6Re04EESK+nlobMlHIsYZ6H3BHi+/hoWpraKr7bpN+lqrggZB3pP21uJC
DG671UwZ+JlrL9zG3751kwCgFEndo1535sjBM0kLxScmflkh0hQqAYD01E2mfUxM
wIFXxaJiszHdQceyAK8IG6ACJ3xKp70xWzDyvGhMGUgCPHPt1x7tbpXVfSMa+9Bu
uN5HFh19+GUwQyJV9r79KHsM/Z14OzSt69EkoGu0xcjA7LYHi/wtEBCoH8hdb9uI
rBIIiCcR7hIvWLn90gnwrMooT2XZGx3NDrmt4L89ER59ksymrOxkERUwsSm2V7nQ
LXDjRrKivH8LO+aaM0XiTET45fPdluzw4ohC+4LqScYOwck3y4B39IdTATvWMclg
wDALe5xjpnjRBzBPi/Cg46e4FWUXNx0QcQaWVxnJg0fkQv42Ze/5NBFmwIcpC7u4
QhfRSSk4sv2zRUcEOkSBctM+zDZDx4hqhONajSz2o3aZjzDolsZrp2DlcHePjHXk
aB0Kfkv+kjOlZow7HOs/vrRKFwWR35R21eNb21mbG/vK/yOtzvxwm0XYwaVMircj
82mx+PsPqKkFKtb2cryiLib0mQlKbGhEBGtMKCwmCpWngSfuwIAZQseygDpuYgh6
EOtrfK9mFB3mlGVtFwc4/4NIAJUKv2KMcqgYMpGSl7DyAomZp18E5FCspVcLcYO5
rTaCyezvy4YJwbgNcjEXcnGLNmCBHzdmuUfMLDN4EpmY3d7N20lMF2M4j2sYEKI1
C6oRCdroS8jwxxD0JgEDEuGfCM8Dja+yrokMdQ9NYH9xNWDVLKYvgkI8rlfRNHkL
QQX1Bu2ih+SO7x3YiszQDNmRHcEv5YcVJCmRxMgwyoRyMOH4FwNtbMiGBbAG27O/
`protect END_PROTECTED
