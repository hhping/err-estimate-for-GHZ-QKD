`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFMP3DUbjQ1rsTVTuSKPtl5kXHp0I5Q7NqAlLn+AHtXvPikRtS4ZfRVk4cqRIHzz
hzyHUJUUWSJpDlnoaaGfesXw6VRecDz8LaGntY/OMupEdXNY0exHOSi7NWVx25BD
CVKGc8C+/Z+78FQpx/IQqBTCWy4XMx44iVgrjI1/PrugGeDiWeRcDonRzHYLQgkm
woTesjfa+Rius0retv1wekIcyxPA/oqrMT6fFTElUAu6smoedwI9Raii7Q5LCRvF
Bxvks5sGmIYDjJnuzEZvZITjsbNTLt7O8g/bB2XQm+ke2t2NEJ5lyHwbuVZ19QpL
6NqX3jpZcRttx104AWZZ+TbrZzHnL0LjrSnIIWItB1IR8ajiOX7kUp3+lwNZTL9E
DniVA8jKmhyRmbZGqmpRvRp7DXEOO4dV2YFossKhr979PnMWPOQKscwC1rNMWOjZ
d+w63q4dqE5I1+7G1KK0XX1GqNKF4b+w51Go3SyU+frtZ8v2IzY+eBLaq5x+rm0u
3DGyffUM/JKmcee/Gxsu2QUfyFyBnfCwgmg/2I3Squ4EQxjkdz4JH8r/bZEeuJGK
sTjLk+tPqsHPACJBMs7XoOEB/8xF1/l2M5r3rXU0RlQRvTnBADbLVLJTGXC+oq7m
LxX0P7bN7OWT1J4u2sK0zNeoM9NoY8f05XDY2Zag0QvAIIvbssbSIjMgTIxOB74j
vSRrFbaZewmyYs3uEvVsJPg8PjOTGb8UmCxc3Q8AzCD+Bj1h1kc6bUJEXM9Qj/N+
y/TxM2QV1cYFS7AUk4nb4GSXhRLxx1ULsXs+jJCVxhBjNaWJzM3Y5Ri678Y5vod7
mZNNHOn0fnDx4OTgSAHhYWIJCqnMDE1INyw2qn6zccYiBtsS8sdvlhnxFm2fKHE1
MYUAexMDDBuiS/YHQ/ksVruExGjJk5iMhIXZwafmmVWMEpYwVHg4Lp/cmUjv2Amp
RjRSZ1DjubAenQGCYKYR7jmLpXONQuPXpW4iyo/J4wAsHZP55rw4ka1aLdd2i9TV
VQTnbj+DrI+doldym5RXGXR2JVtcL4CXupqaSTqx6sY8A9vIzUBObXOKQNYgi56U
JvZqsE4EG9TrLaXlvaZaxvRrpuYT4NiA6dWtkE5+xTLsx5/wP1VuijYgQz4MgpG4
3LIM7DHnkB5kK8snM/2ABmLJMD+RmOgPDftfZ7eZ0q6DX+w/oAPzvNiGX7ZCg5GF
eejxOS40Vbrhv/UXRvQXtFr0r3PwPJluIb9XJD10Ym7mOSvSCMBF/Y/pG5jyNEhf
JuhOXm5c3zmOCmRmssnxTn5VixeMTxm6hy69l/xZFBD4Byh8IeKehiZFTCMuHow6
zv3Z+n9PlIZF21DKX7UXV/CAu6BMpbpyr+l8pHlgA33IxP6PJBqYTcKYaocpTMpB
4rnAw36Trr5lCPknEtEOuyFZycSke2TJlaiA9EpSychfjyeuqXdXEHTuC3I8DOvv
SQwgw6rbmjjVpsR3oITyXXNkFlWoevnathLeQkx5BGxDdCJ4EUOt6HfasfslTUtY
SoruvFLimDo7EC4XqLkK7G56Z7NYbaJ+/dBKxXT/3USf15whpYBOQERhVaPo9WVV
i2uQxH45LgT3wvs5cX2K4x7YTYcIf4v6A/85F9XG2aCXTteiB48YT0r98h3NR/H4
GNGg2VB6T9kPWyhJH5Y5zlo52GufEbkJuaauCpxy2Yut5rXpmkLL7u6WuZorB1k+
UvxZ+nhgbkd3kxUxCNxHKg==
`protect END_PROTECTED
