`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUkZGUcSBBysC5v0sVZ/Xgn/XMVK3Vxov7Cz7CS/omARdtXn4RtZZL6ZIIb6CwJB
5r0AeZthg7cHENUjHJg0arRxBbIzHgCL4aJ6khF+d3Ky4H8KpqZsKDmEKSE2jXTs
oZHmrm3LlnD/ZfVfXjYQbgU+yW91XFHtUJiAjy1VBM6hlNy+1+lcVSxIsPOqjYvA
`protect END_PROTECTED
