`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mlOm7M1b0VvsygC3kSkFHi6Z5gWtmB647Pr/WtZAVwN+jDcqQ5nYT+tw8GmRn0SG
aVUBCC3YiUDuSUK55zl2vKls5qcmGifk/nNOEx2adSA+bacSsK6nRC5EQ8ByDKg6
xwGh8EIN3cJ3JPNBgsdoj5RK3REp/mLpp/l8BO9771CF7ZaadSZ61Lv7BJgsVpS7
qttNKIxm1k8Zad73wT9+vhlPRuwj/EukTvnQhs+4B9vbFyzv9ZYa6PPFoXkxBtvV
aOscQArnR+URAWjWusehhBXG3NVnPT+ogysZ+7RQeflWKFLcjUpqYcodoxDV6ICX
p1XXbyTxORqgw36sbW4oeDFKAvZhc8/HjXMh5hvDTTEqpvlYagdjCOIM17qOD9Q1
fWpoEmwpE2O5mBA3OyIRXoMAm+oKeWtu6oAuB/dWLClEbROb9rX0/046oLZc9juw
SX0yOnVdg4aGR5j4+ANcT/sHcnOB8S6TfO9z+bQDVI55yzV4ote2cdeW9xpUCUuQ
fAO2tuTReg1zJWDbxU5VS57VME8aIESInlyUxmibUklPtkIxwNSu3pGQvSPOcrMq
crmPAkD0XNgyc3TuAttwQF5TGYIdeYwVpry+x249V9LleZFTbCYykKCObvfnWW8e
Jl8WJUvrSSvJBIKtgZhtkvm4rgFSci426PucmVbG92mMurm1JAVDlcuRtF33+GzT
SJ8PpJV30MGTlA36cCKqSQkdzlK5zYpp5rKP+MTsl29Mt7C46DmQoWJxwevpMPhd
UMfP8oaLKSGOJXjtaMazSZgzcV9It1xw/eShEWO1AItetT/uExX9B7/OCFNTd41Z
3wdKkuqXZ+7ZKZHQyCWhLOFRQYlZl9RNAo2tkpU2TE4YrGKra50rU/6r8liwhVh3
EYU00/mW3rdZ021Tb7VFGamDsgzGgCZMMWNeSDLLpmQk0DOLfFgCsbeYd7OF5DUn
c0EEUrfwqrj/G8JnXo90o4keGa+McH98Tg1sWZK/ppb4EOB4jf3Og/aCM2YCBbDw
cInywrz2TQpQO+GjMRLIQFohXtZKNA9xowm9HCnbFfxPECODIRwIydwSHrvon7R/
NEbA/EGMvHb+vO2ETWGdY1ubsD1PBVy8nZI+lwUNtOF0Z6Ie1CrvbHiReHXuyFxV
5SuqAipp42qZRf19/neUwrdjLNvrn1ii9Bsho2T+DQwyyHka+ZzQB2H4m2qVFf0s
`protect END_PROTECTED
