`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ud1TdJ1tYGGnmTZeMFX7MAQVHzagj0l0EIdP6pMH1RgkYwR/fUyy1QtzD/Us5rpX
Ejwk5es7nHo3QT5g9ez3M9xkru074uUYTmCdyeMBbkc2GTMOZno5q5k2mxxji6RB
lgCNn54Dm2QKmQalHSYGLq9G0m8Dcc69hx6nVYuJjKu6MntdMGUuKJ2c0mRa6FOp
aBtKMj8OJbWgXWvJVl/E5soLcmFVhkeMdVzptQ4B7Xi1sG7GfaWVY+JAzMVnKw+8
wJCApXZhH3zbQ2zZVZagSWBs0c3Qy96B86nSi7Hv6GtI7g11rXbGASeY6y3NL53Z
qFnC0qWfeBJ8Ucd4bDplKvaxQ+e1m9w8peWJAUlSyFgLmsYm5jniLmTUtskWot39
1IkkRfKmHmxBwCwlSF380U4Yv0kUTudUdWjo9GWz2lEj2bOrBONkZz4vtwzfPwPn
CClyyRs0j3sNq1P1nKXhj8ZHxyvPDT8RMzGiGV3bIDImChTdHitenw9RqCQBdkxi
UuDMa3ppzmde3ANFr9Jyh8KcnS0mEqf8pF7h/O9BokwM80nr0a2xZtEi7TiIwK/F
ZqfHlvJ0v1pWO6yUMNVQXtV4gNsIbKZnrB1VrdSv2fi7HvRHfRSss4RqxZYXzDzU
MziOz4Ov4Te64e2CIlz4bSOhQc2EkP7Wdx44Wqp5xWTDSLmNElCLI4pUZpAYkJZ4
fTb2hzSfV7sv/nP1rpFaVw2FkbJM3+O38e1swKjNP1uw0+VT495I338WuftU/Fh/
a7v1BZrnkIVVw9uXOujGSCfEXFEhpuw5N9mGlqsUyjBKtI8pPaK8GS8Fz0bu6nci
GwQk3kOmj6h9M+7nH3KLO9YGqnstOvIfajzQCUeV+hmhDVEOrGovgKonQeNu/9Xz
YI27gyCbxGSvONrVQ958no88QDOBhh/oRkN2Z91hPtPInj94bSSlGRD6EG4rdhsF
`protect END_PROTECTED
