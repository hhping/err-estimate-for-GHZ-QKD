`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLN9WERPdzYkAU1ox/QH8ge8z7RUnBmgysLP+NqQIozVTeHnxV7101SoE/8hqufw
9BtgmwVGkpGWP1FQb/nMJ4F3/X8YLjhG4F1S8kna7uZBCnhPNGF/3LozsUVrhamT
Z2YpEgA0WS8S0PtDTRy568YV4hsVCLNKqPMmeVTTgOTH3Ch0tUTwNEoDk51KZ46b
7wlvC7gvFRZBgx7ZIHyIjA1viboSV4xTjehSGL8KU1F2QBIbDIzYNj3u3J2ipI/L
lh2vFKxyRaRe7pnwGuDO/Up83bJx6bjnjDK/TzCVh6NUDLPIuT+238onrOIEQ0+V
9QO64QC7L2zycfuFBNlayTlFNZ0gTqvoWr6M+6BFTIhmhI2cOcNpUtpTS/8gj+82
pAquyLvX0rJym28kE/4TOZ2InllegmtaAPcc5Nw1IDbtznZyZSy7Eu4fh0QqyhX6
XxD8ygkVnuzdsqSzCVODkwbkRWuTSV8bjB94V3byYEVQyBRd9kYJPeFrwrijfUCx
KfOmKJjmHVziiJSV6wEQuQXpANOQ8c5euaQbVyNlrAKp8VQUw2YnQYl0Fc3t5AWk
IBDuPOgq7vjW2Ag4VDnyaSLlxZMxRk6fyvkI8anutnnjp6850rB3d4B6kWTyzPHO
AcT+/DLw6E1VrX7HN9YA7BQ1sX5IH3kwjwHiFLrvKFgO/N9gntnBMc+GbujM0mda
f+9j+qf8rvAuFA3hBxzVE8rl3IN76Ypoa/oVHo7gGx75O80z85Vf+pwGUXdxUNKT
wBpQYDBqb+FfQKn+Oqa4ZqDSwmIBfTBVmRcpwo++jv9qVrcE8BhqNAcI+7vTOP9J
EADIWPPDJtzfLyGH3xVO0Zp/asDlQaTSZkzFv8WnXIzVPdx1SZ/JMqF5w+XAjWxf
ZrSxv8m1iS0GRIS4Ig30XqphqYTMybJA7OKgH6NqDd69EEDq8zhCuMvfVbymGAzf
TcSOQt1kWrEJTIyJLRuJNcwTdPp11nv2Aca8p92HuKTWIGw6WD6Cdsc2uESh5Npi
TJ4ah9ZXibIrfQ0cwmj/oRc2Tc5uOkzOT9kFad9xmcb7V1O8L14eeC1jO+LR5r8m
KSjDaDKm2Pv5w1CtH4JDsr7G81Dmh0OnIynspCVy4PIDCSBpX/+4XpuxM/HGhwzl
bRfq25uHAVkARtP40xDE7hq9D1m1DCMSuWxX6RMdXwPK5Jl1do7P5Yp1HZ28ZiZ7
8A/h2zzmJu4S7WCXV2pL+pHPEL2wLap5OZmoQEI8Dbbv40HgeDrQE70OAWZaD8aC
L94ci8KEB/2fxW8kgCGl1YM9I+3vTGGQBVBMe1hRGSQ0ZnOEfCSZWi3rY9ww9J+Y
XHuKnUAF9PnCISomd/hxxCVv4j4QA1YkU6+kxp+RO31yjgP+p+xI9obb6NxdJGg5
VHo5MOMCZDgFh+d28DCrebpa54QDDcuDdB6lIEoZnuBS13tbKAXb51E+FDZfXgM/
ORxneyQXiZtEn9VPqChts4jHBShSGiR5F4i2OeffbBYpWrA8koMA7ITpKBXKaFYu
X5KEU8H6nGs4MiMNjHPKSSiut39tFqsnSpIYgxRoGpPlzQsekCtF8ZVMwXzPFxuQ
77Szg0OwuDd2WCgYD9Cdxu6gl80S21vGaB+Pdts7TbIONB/uNLofZNVwUCDPsMxq
pPGsA0yE2DqlvV6zgPS2jZJMG8dq4QgrJ07RHASO8ln+ky/ARsi3+XLTvYEwSWXA
Pxdbrtt8uqmbrQcu4HlK4SyprzuYB17+TC9zmDefmY0=
`protect END_PROTECTED
