`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vPiSYG/PBtB2ltPN90x1CTTUvD7gjO5bb9djuIR0WUE+NjVSEnYCCuP5xLPk/5/z
fUb7EHYaibKGeO/2mjCAyp7Om9K+NPvyO+7qzp2bTj/3uLWXm7+xF5QU3TqI5PR9
0MyDWdZNBoSxyoh8YS0SAixEC42FJMSaVF4ctUiWl5qocY39WyEP5jQtfNXYyA3b
6Tic8fb237UTptqo4Z7puFjT8Z782ElXEo1YoHnJccWI8vOgu5PMV/gsiSPYKhuP
TdiwEeUU6cpn9OuuTG13h6inVZQNBPrXgj8qURQrtNVoY87ncmZlcFVH1MUmNKQA
4QL3V2b3iifRu2PsC0MgxsGMMy3pmr0EDILARdk9yr8moJbQQttDpVEnhaC3/eK8
2VO/37PxLhFhyKrh4Sys0LsnrAB0/4XKeULKPcjeip5hSatqx+ASx0mMZMDwxuDN
+ki2yIX8QEgDiav62paBve+MQp9Ekp9L4GmdC9Ytj66JhO8FA1fyzWPrey9sLvJI
qkqUqojdbeVTlOlriHLZ/96VRpMLbKh9Oi1ZWGzD3wMe+0JRzEF57mbLL1VYSKCf
7RVfS0rs0mxfPTSxoSz4+4ewOH/jqy6bOd/bIrLSCoJj5reIUwhNJo7C3k+TrfDn
l5QMVxjepYEwc5qo0quo+UPqrcMTfpURPW43ZHzURESFQ6+oWzjXjWT/sCAVzgC2
PCFI3FKzMU2kXl3KePvdpQ==
`protect END_PROTECTED
