`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dreNzNuflx6sOzkqBo17Kq+PIsfjSkjzng/0R3cbjpO5lEy9ETFXSsqHFgRe1Aq
PQjbifxbt0wjrbIkXh9FQhep31bu8ikLyLuKqhfRH6wbV8Gqmy+E0uqVGSotdkpg
otQjgjLaan8xgfoY8HBZgqjsoJ3CBVj+7QGwrz6zHYSKdYVb+Y7nB4xFwZOGuCCo
5WTOHogZPSHCuvttZzF1cn9w0R1kglhBAV5Ete9a8ijmk6knncUY+scR55iWlgkF
2ws8D3c6gdIIEwyG6pJtBFTCUDjn52LVZsnPrirf5DNsb1pZ0MYhBYqB1uIB7xyt
msb7RGOPyCKodZ5jUzc4SH5T1Nqo0MAKkBd43M/gZkC1UjIF9KckDYWd1svupU+B
ytIg1Qnw2bWg/dZKhurYWYwnduL5JRe9iMTJDWLx3EyfqVmxtRdWo411IVHGUObE
DkliF/5O2ACAI+/IestXG7mM56U+2mIA+CMSM/94ZO8EMO310lEfRC7gaoId0cMV
S7GwA8f+lrTcS//lFsUErtLjv8/V2XhvNQOZxtj+OeYE6djWeERz7PZG3WhtWm+w
xbygmYXbVD1py2cvu8a3DDns6//WY81l1QgQkVlo2lpxAG2tvC1aGD9crcRp/7CF
ZNDLgOXfaXN8Cvbesye0bkS6Tqm4BU105q1JMzk/yQGvVm680/fki52ZkxRV3cXx
mGJBhk30qvq5GynYhO39/p4iUPkyebgCK3sK88w7VYvR41QSTC9wZ9zPhlcfJuc5
lgZmrd+/L7nWJoPaMaJK3t91ZnQLFMELedEoW7F3iRwYPoJm1qcL/SAm3esVJXm1
/VSVdfAhHDm5BsQs0lMhickMi8z7tXr9kpYeZKp3V7J304nYNRTQtc+lhLLfJ6e4
iLl3T8Pumw9B3Eow7w2Zdwqb8hlhdY3B0jZsahawv3nV9Dx3XRWfyUCGvKBEHwTl
aKbVteWbRYoZTt/uGMSgk2kApJPxfiP32UCFPRJHliyYH7PbK3eY8BdHmMehCEoz
`protect END_PROTECTED
