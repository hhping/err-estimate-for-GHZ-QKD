`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/rUQYmbGwf4n0ZU1W0FptpLZuywAQ9tLBBKs0GZgS8MIWXUSAn8pjVGil5JSdwS
sn+spDUKDhlRTdSixzqDSyYWoYyFqNZb0l1pniGz/hx7PKlpD7wghGdirT1RL39p
U1Hh5E6PzKj7r3QTNaqEchFstm/POSmckSIiMrfktyX0I/ucjS+97p1BBI5h6awe
KJ/zmHlL0wcrkdjxIBFXMrwugx0iOuMPVrBQDynPmEbVmngwhpp2zSMOiom0sIhU
h1UgNsTPxcud6WYrAImQSdFwhcdh/pJI5bt65Wv+7iZbb6E4tkNV3bMiVpQxLxlJ
LdQO3iZ7TOwmCSWbLW9wUfzOYCf800b7U/pJzOZrEMy3376QSOFA3eIKMwod8yfb
yOVbVb9EHAYZ4XtDLwLYT3+1KwveQ+MdsFgD6gFLUgdd3S1cIHFVzZ9GuZ2VR/x0
PINBhcEdrkYU2xarZJSP4LUKb6FnXrBzZrtyZdmgN4w=
`protect END_PROTECTED
