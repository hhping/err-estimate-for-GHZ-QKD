`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
coTZoVUnG3XMYK4YcW4Cx2ROxCutFqPsW2fB0H0/7ZB+/UStzX0qi+qcmTHt+n0h
3k6vv2hG6J22DA3mHqNXgD4eRgGhOg8Y1M/UGQiPVrURkHO4axDYi4oT1cNGeAWT
ky+OmfUs5UUYyercAOTywABrzPnSfHGoPIvUYpRSBIUsz+FySJJwoH9XvxYFKGwD
k/dtzluNwYm31pnI401fic/WWN4snNkKuCjmMevXXmntTisSMfzvkzAvfhiUGjEO
xvcTTg0gm7noZkrMj0nRa2s3kKAMGAXQ8b5ZhufOTS3IPaKtMft1Es0M3Xb2mzSM
jvvECTpyD3x09rT/YpSxsjrPHvGwjM5G54EF58qe675t/AtCron69uwuPV7tiZ5I
iRl/qcRElMerlcSyUEJe+2NQL3ifRQEkqP7w5YydUgG6IScjE3j/apSG7UNg7hAA
Uw/AS7oLJi+bwrhoS5h65TkmfKP+hrWxsxmES2nOwtv0j5VSqvPHZon6cEuqYPdI
YXahygZ7PPwAou0+UzbGO6FNUlgFhwYNi54BgwxW/VI=
`protect END_PROTECTED
