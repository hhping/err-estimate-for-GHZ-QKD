`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFKXN7DyLX3LzBe2kB9aDyopsyGOOTd0nZUShFkjVV6eRmI17Si/u3O4VAoRiOnq
FQJnE23TKSX1izww35sPHOYIl0yFzrFNrxiXX5oxurlJy8WTPyWJaNM39LEpkXVy
YRLeP7XBdfAwdy4lBT+ivlklL9fv46CqHDcLm+QZ/sOenxOAkpqG60ZsEGewzElR
655JC3zVGsmcwRQJiDe/fqNLMjs9mjqdDrtmWyvyM4PcCiXhu7gqnEvfTuu4WNj/
9LOApRA9x15/nUpAlsk6l3qls/wQ2qBw7+IOeQwlKjBqvS1senEoPEQWvy1YFjkO
KNYKaRahUL6G+mtXKri+ZWWhBV+o2WUclc7UO60gi/bHkorv4Yuc9lDTyfgqps5T
mH+ELr8Es9cCKAsz7FcgGRYSoS63BaUiR3Hy5ctj9KaIEdcEVbUTTE1BTehmVi67
I3ELbCzThYZywtox/LV/i5+ES6mSCGVSvQHg7iDJjKNj8QwwP1FV1HYpl6/hBp9F
hyTLHcjrc2sRK53zq8BIEh2k5Z6MfVOEFjxBiHj/oOJdIOwKZtZkok+PmhjCdmMJ
sRhf5H/0N4Vj9HoyAFDyuwu/nbSfeyQukbAcE1E/5LdiDBTpehKFfukWEBc4NUQi
`protect END_PROTECTED
