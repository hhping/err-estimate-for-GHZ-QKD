`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppjot5TV9+WQn5ZrtLLls1BalCuxZmTgagByo5LFQ0tu49Ei4hOLj/RtFCbEAyDa
7B14MLiABxkZQvwvs9QAvfiMuTnwo6QSDet4DWu8I7KoLu5LKl4XvXct7EnCQDI4
PUDr1gPaSe96dKIHEX6kLjnHZtX0xlo2IjOCgi9G1lw7JiHpDoRXjbmZHbJeHhV6
EyzOjBYmXpzkemg//aQnk5ar68fR37lO130z1R6vqQ1J5WmY/sZ+aPg6Yf/5FBxE
R+XWHA3IlJfk2XH7cghk0j/P+gQk+wnpH7XpnBeh1+nrXV4vd2LVbTjXeTlOIN9S
IcZNmI1GCo3xCZwNdPVJ1ICqSlBAmGP9wcamh2IlAqtwYiDHzblQ+Ik0GhIsvxFp
dSycW5zsbhzQZD5JnvhJwUO63dTkVZ06aLrQSR5A+S+hxGbkEVggcIGtKr+m9GLq
kPO5p1Fw7X/Ap6SFXPzvCuibjNdAzcN117ZIoKxfmxXk/vHp5N7YpkLuEqSRgoRt
TL5XR3CwEzc8fqjmxvCDKPpMJXsTmcYnLIsyKNmOdFyQsLOdfo9qFEm5jnxpGet3
FkGTDQdfm/jGUG9w9WlndNffLfd72WzzxGAwdHBwyhJ2ShS4OqwcKwC7DW4s04oE
860FuWZqFoRYEMKNKwOXAeoQ0mEUnN+v8RUsn4B7/8DAj6rZV2Y+4+8b31L3pIFP
lPu6NJBA0iUcKyuoDmrYOLuNHQZ9WKw8qskXI4ndbarNDpLDwz9ggXu+u2zO0qCz
Ni9Y8khm2kr/1OX7pt2pxlfpFfSehHXNWTaC2vJVJETSoKinfEy1/j5c6k1srh4I
IFfhNQybi2zHxSp0K+GSojikmzFS38iMg2pmrx/zh/QXk0sFMU+2TjEtlogMW9w/
xEgpOJxi3H9w4SI8VOhIyahVKy2MHkFMTrzXjwvTVbzqVeAIEwxlT6nW77CdFdh4
+sPU6PXCn38vZSNtACqYujba4RLrYOA5i1hVoytBJJhiaB9t2o5qSopf6VlAC4nT
uWxo7zsVcuUizhRBq5sQkk4/n/ct0gEu4+FSuQYSSkQbhtm9Sry+p668JjI9jy/E
SsH9O0qzAteFGSfyvIEacZEYQ0I/lFx5Gd4XqE52J4tABKYKbHnpbBFcNi2sFmI5
sG4276RYvPloZ26k6lgSVC64hU3xv1dgykaRGxLRZEODOfbF8Vcj/Q0kNpdyQ4bQ
ihOs8QGA9iHZdlR6nLrYmMRK12xRGeHAKesGQfeOZQgoiRtNEzx2yG8H/hkQGZ3l
2Nbl8t+8Ogwd29b/dYtHK+8x8TKvMiJc2cN65Sk3pK+7JEjrKb0MhdPJnQtMhmvO
2G60N+qBm+rBzBKcQSOPB8WQ0VZ358Oaz3MlZn/EyBj8rdUhCYhAqbL7nC5bKfsi
kOmc3N8eYTVSvBFIqnkcWuUOtsMe65zDRJdrhe6z2pYqVxui/P5G4YpQWjZPSpCJ
18l1fGEeMQfV6YHMaVS09iVX5o7txDHpc4z4POimZavAjToLs2S9BwVKk9Lp4szO
KXnZ0GiBQ8PG+5YLjNEIciVgEYmbKmZ8SQdTsIO1LJ4uH0Fgc/Qs4G8zJ1fa+1Xs
Z8OAhTimgEjhmWg7X2+BzhJUGvZ/r/zDIwcM5m7MJxBcj/aoDW15QObhJoK4L/wv
EuMSDOtXZD/Nim5Cha3pSu7gfFWkvcgEodmz6RAKa+dHmdnfXuS9KU0LLCpZbGUy
Rty0s8mR3jJmIJqJCyBRNy+plCMFrcilrHVr8PfdSS+8qTV6I4ae2JmUSTyVYH9j
qZyPvPbF9EZa8tCR1LviERnnmmT1M32aVUZe/z6qVToXMVK7CHnIE3DjQGtsx3Q9
iu7KEHeCt+uJeDMERdFalx0RDSIRZ8T6EwQ/qRk/cT2SiW1JU0SBqSvIbohL/oh0
knQJR4sBGNfBG0pNGfmOsMfEcIyUftrHUe3at5zjVojLb+cPsx1A5G7Qhs5rqH9s
Prb1/3fOxyTzH5skuuKPhedtl/m0OCrcH+pvI/Iw+S8523l5R0OsTbr0xZfZO7LY
WoLfDvq48OVEQ4RZ8GI1BQ+RznMxg6nOOSj4inTCUPLPpIjtrPxzGh3vTYOYS7qe
gfAO990/MP/u9KXzB2WhJgfSfy9gRdX7AtHVm7/CvWoPumJ8mNXfs9tLDUuxOlb3
AkPcTUhAZU+8z5/kCejVNm170VqPtQ5ZkfYS4V6r7+S6+dcSh12aJ/EcWPPumO3T
5s2HRrrQb6tQaW1oVSh3TsKeEs0ZBpvcmMLt2/jx1mXUz+5mEbpd6OrhEis2DL4k
9yQ+dmGmgMzkczPBZR123Tu+w2kU6oK0sDZ2rj02Qu2jUpS/n7SWPrfaN9l1spv6
rxEmrcpeGbu2R0d3XcPze+ppFW9MzdDXvgcv9AExIVsc6C24bmSRPi3u65Vj4ojh
ZbLtVeu8A9HdVZQMfa8kLCtumHXsS05yxRp37Saba/uvz+1xdvUpwmjh9TUiCD7T
Vp5Bw3Y4Y404i1NTddor4lzsHDz1UOIXID5PtOoo884TwJ3Ac0AxkS/JRWNzUA56
aBkgKV4O8t/4Gya92iM4vPXlEYw/r8l4Xy+DIALa4pA2rsOYykNE10y9f6GLHruX
R+Uzkt7lc5i+eoxs2ppc1oQqYfez4WzgDxmD4pq8gKJwq+WS098MPCXCZPt/j2bv
/orT0aQllDBC33b/jRSoHOEpDQIJY7hPbQM9boRkZZpRxWr7rFhXGcRx8gWEEGmm
5+PQfpJVHpn+Okk8wS6eaWblFyIq37uDF7SpXr7hLxFGbl52PlrwZoVcNwpziGyG
bP09ZlMT5Sq8kZL7ncw1ZLU3eCxWbn0JdGVcPCOJhxTUscoqXtYcVTdFB4WSxfwk
Qf/4tX1XWsCkd8iN5Zg9RquqrT2rN8hCltXnSfDgF/oCafb+f9qVZGd9ZVgCDhiI
U9LbUOVtDAFVlXhWVpap3QzqujLXK43sa15KmKEV1au+cS43tHwWq5R116W+X6KZ
earbQhIX0K5f3wB2llz4QZcB1dprldjpC0h19VtUnccc8ET3zihYmw/NvdOwVt/M
vvrwQOkLQsiiGCf9kCVgPVMj5rcbQfjllcj+PNNaYvut9auC4fr2CvD7UNQxm2AT
37Qx5ZyUBXsO77seOQ07ixMaZJCdOSmhS3qMCkdlIg/gxEHXB70IAIeEc6nRpRTP
UrSJGuokWiKtW3sv6ct+TMO2t6nez5+MkwYFkNXOt+pcpabuchfMnioAc4KA1DYO
vOc7X9vjYvv8jj2+mzT8etY9TQN++ieUyTvuF9hNFL4=
`protect END_PROTECTED
