`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NVcGMRsjPARZGjmmVcwPRtatZdEcYJMN3GFByWzQJyMOzoMCP1MimLg8ZTvVuJd
X1G6fYQNc3HX2XTvRnEvWeIDxcE8MoHUEHDXaJBQF/lFF2mTTway6+G0Rkgirwms
Lha1ov3/qD0oHV7ewCL/N6I4Id45JxcPlVsXtqgwIa8jx3X6gcxmSTZC71+HwPRw
ENtIDomrnchQoac5KxVNO/wxnctehAwj10gm8nLKrDWhSOKOxioCJWvUjgHDZ/2A
SIJl2W9qfMgTT8VdfprLpy+DlzS/rtAjWUHQwZ/EygWkx3YIayum92XXWcl23wqp
yA1PENPqnAMqM24UGthZFSMj4S446qY/SCNaU/cLyIIJd2UWNYsFGyKXptxh9uJo
CGJNs1OBJitxqKtTxHaI56+EWiC3StlF0+N7E/yndN4xePipZzN1cxs0eLBQKBuX
VjIEv9ns09V7OX5//G+egw==
`protect END_PROTECTED
