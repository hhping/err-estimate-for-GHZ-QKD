`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+PzJcAzFiiJt1ZiqtziJ9YhwT7tytqHe5BhOSZqs2hVbXK2Sd+V2VrOBah1rxcr
qMIzRHs+uGTYKHNbrqh4kQ8/Kuxvz4fZXrKugUedyHrqrj7K5oa88FBnWlJwHYun
i4KQYUYWaCYSObuhGQYvOxAUmD4nCV9cqljgmyXUNkhQaVQqgX20AsxUGez3a8Ht
HPslSjyUUitrCS9kh5krqkDHqBUlNmb7uOC/y99om84sFEk/kTfPO0EsA73cBCAj
JF9MARgkdDIyaZ3DlW3JghAycqKKXwkonwJEMRGW0HfiOJQT0VsNC37ZN8UI3OzI
Hj1iLJzev+uTewjlfSV47eK1TmaaV1tXhmF4ikr4ptl5b4xGkbfTSao4saj+byQ3
OVwQgawCLlFg/QZnO48SqpKxh+V1uSE+sDXZgMpLBphxWzs//jHEHqF65A2uYvCQ
EowG7Imb4iDzqECy0rxHY3VpXh8Sl290lUFH0joiV3w0J/8SXwBonCXNBsKA4pHS
2SRhqDJitpfG5smh3ggx/lZUCFMZWpwDeePVbuRNUjxnHDyOn0TfvPOPFS9/c/bw
NUBvhabz/r5m+QKRhpR6M5XjK9TUGezqnDNMmEci3ZWuUcH7ML/N193FJ/diNBW4
MZZOnYB4sB6PJsM4BWvNAK2ITPqnxHLreS9rOttO/Wc6PqCKUF5O5jjKHo2ehVvC
mBB5W/yn00Xyt7FX7+y7DDn5jsaY+l4ZwS5uOliHjNuRX1i0J5hkLMNWCASplJT9
zkyX/71D8GyVg4Z+5QY099UFTIzWrDC5RPv7/rhh5KajGIEjk9bGbaYpDmKHgDv6
kDIgUmYRmJHKpqB9ujxuJo1y/rd1SGjAsGa0KMETK73AGMSP5uJ/zI2k7Twa5zXH
3CaVoAbq9zaVs96Si9oxL4azOJnl3EC1VffyWlee7Ca9Ak3b+ANirFwHWIFcCXhd
Fz9b6JSWDe9SissD11Q90glvrHpksrXyMkF9NE0Agi0jvpK9Z8bxkzZDqCUaxGHq
9d734zHeoDOZ/aecqJL7uVRcGSM9UHPQVT4wHDwJe2f9lqn0qQ48TdeR2T0Nnef5
P9OsDq0kconqlkgcov52lyeq0DsoJSyPSxeodJ1OQ0LovNXL35bTuOZ7jZWucc2e
Xs3mQAYPPJs6XG9yO3ICAyGwlbHD2IwsbgidXKRmwUa938AYzpVZ97SVVLB5Dpiu
/JqIUDZJNT27KiHpc1wcV8mTnt/WN2qEj95NzXv49ZPk4WeWzJpTSpu8GiiVlNXL
E7viGc3RiX9P9Td0x1t48ZBeA9lrOGH8FOTK3AOw6awJwxjPVyRiVVwwdIWSy3v5
IxU7R/d4VaR6eTc0nysoI/ITqAaB7KDqVVufSLjAuo4zhGgGbWtHDRFLBmPrz932
aR2VopH0AzSg/lNNzNhwt2KNk0tAddQzWzJyN8R5ZX55GKHMd5dLvwDsFIsoo6nu
`protect END_PROTECTED
