`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CwF066LafDnhKu0RKIj9xdxb4wOVQGlb7AHfzkjKX+VukCLGtipVnQgbExTLTziY
YPdeOMlrIlPLRJ7cDbDDe2QBjQYZqMuycqtakdCMZ/8lemEF6+nN89FXR8mfarvm
4uZY7A8VyPntl0Nt+teK5YjdzI4aYhvoWyFAFYFRWJQL1mXO5/2tfgxNwu0HSlZU
tgWaraa3utcvz3qcc4VEgGS9K6bEgWD9F/glujQOFLgusyw4rQ8XyNmpGhHop+5l
AwJJvmTr2tM+SL/ILvOJYmBgGPBR+lJOhSALOHiwCQ5gP0hPgG6msl24kyA42Dnr
fZnB4maDy+ftdl2dIc3s/zWxqzElUT4HhqW1pUiwNGMHOZRXVPhCpSb6neqikzHN
i3xnDRsyU5b5PKvKVXSZI37AxUrHtJkfNLrOA3gKsiwcEn+6WRBNypIury/NLbAf
8piX46b2Z9iLsarCWhiQ6vu/vlN7ebtwlV+FoFe7ESl4NbqFqokP26GbUZqm7wqM
HxvM9CZ8UKQ7s9mN8wcdzP6iPexVI0xCFD/bpNVjra/DeY4O/1CzGzWmAfIJV83s
4TBLjM8jTufBQtuQgDKqAVy2CmpmKudQ9RttCRwdKiQPFIz1VnZj8uzZS7p5nn/4
WDHemJUijmbzuO4XQ4/EdqOJ+TIOgyEwSZdf4blGkZ0+FeWJW1QtHwWxYRQay6z4
aoVu53SWNDLGmEanGYW/3MMnn32jYXstywKtaHDV+P6VrnBQR/nb1+TdhS/WzOK+
VdwXm0HgL21RiiY3ZMQeTsD9TU5u5JtLQAg+yv82v10I/FNziiRl9JRMOK9uk76q
qQPHLUwDZRR1wRafSEH1IQLp96mVu/w23soOp4ajUxJ+XUJlIWAA5nt5OwK1Fsif
s9zUwRVikbcJDEp423cGgA==
`protect END_PROTECTED
