`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5z7CMYhEHBpwKmDM82fhiwz/TWLKdZCXBRygOc9K85KNnJRI0/BgXF9b8qaKNwz
f3qUmJPV1YsKq0mC9buRMIC2kBy9pxugW+mgzChPh999B/9Ez2acJxjILMo7v4MI
5pEj4AG+B41zY6eOx00FcTXoDv0uqlML4hhGllmCuJLMvMu7k4VEyYhjj16Wpd8I
xFlklGr4WPRBWhCn1uVsa4TPX+r3Or0M/V4LVGldyGNZ1Q+dyGkPoik2BBDW9RiY
Q1lhFy2oggpSQqzARhuBkzp6fHmlLAdF+bQyfXJMx558HFSu0NEhvtIfMxyCJzNf
XG0KcXdfihkfiJZR+wLhPkfRDfollOHj2HTVWYdiYjgN+FeObHB4ZHKBgC0cOitk
obk44y1qdAvS1PGGxsX0BCA1skfjC3AaJOaCvqWa6kEo9HdKu7s3kQuCbSiRLEFj
hxioB8mVi/Yp2AEqTMDoILdCWAzYS+bOkX2EPZxxfg2ON0nhJk4ZN7eE4l3lMVeo
8EOPLKNfh0x56Z3ffJrml0GCmTmU0H9KvT/wr5/Tz33zLJnHNcBuFeKmqVeUIgYQ
uU2yGVouhK+KHvkCKrmC2wxtnaABfKoP/Cpu0O1TpXZp9MSBwl3/FIoLp80WKUqk
SVJBoufWfKgrjdNqDIrogk+jr4dQz/lbNX11p68lGwSER0piFnXXWTkLn5QMaknA
GqENXDN3Oy7a3dIbwb7g4SJcBtP3wx82xXGdxTB9Ruvx3AySc2A2XsZ1i9wBlXSd
NhrnrA08dlpJHcOs+/CES1NK/QzDtVlKwyflpGJMTn5DI+pOW+HK9/i58N4x3g2+
ru+J5gC0lwMbN1k+mKDbH9sN4tOTvDPzLIorDA6S3vK7Y4MbbYOJNouPInmdL8nj
FVxwwwPG17rePSF6+tCaJLgRllnnjgAw0+9nvWEgnTrhXmrfBoxs7HHIYs6Dda66
Xn3EoJiLg4YnXKVKoi7FAHdDLa9e0z8dJRNOXSAWWWaUTawXu1Ayt54KKPsb35my
VIyj36X6ov1dSgTyXrM6L2oiYunJJwGB+f8mTBdnEbZ9PfBgdVRUiTT5cThe+cnW
TVNdKvn7VgC0E0zwhEZFtNf3nzZtH0auam4kMy7Hq/L6UTlaq3KvduO+cc6zLrkP
WozbwRZafg9RGodLrAuNY8tS69TGkdfd1Dz+vdwcXx7bmoUt4wOjGOFefPCWgtnn
InIkR8+VpLqmUhiraXCdqARaFusFABLvDfUVouI3WwXaBVRGfqoct9J4L7YvoecP
N0MdDYqzs/mDub9morZbDC0KBXDIeNtJYPyC6ssM6N23K8mgEfMXYTaMrbVtq3hc
QW9JYG2eU4VD3twBsK+ZXbdXfdHSmX0C24HHoaJrd/WbKXbKB1zSLJI2e5DTNh+A
xZHfVtRRmrCBPdXO97lBNWFBCU+nfMLesqrBKhty8UVBL3UO8UdgE18okOLoKmyA
5STEPkz3EsjufsGK8PLCY061yiqdpxHNnMFuo2bc5EAh1bdNU+BhjgxPoa9XuRox
8Fke1WlDCxy61o3IKMVd6/eA/MV/iKYv5kWchiv7DS08HWe5aLCGl+vx08Y15Fkz
b1aJV8Zb/lRiqf+5R9aktS4ioOuPv8VZzBmw1MvtaKa615nzlPY/wwHLDJw+2EbR
wO4HjNwcY4MCpZO/QIOihujHY7DeNd/1Vi5d/V6WlVy332G/53M0D6EUv7JrVoML
gMrMyYosp3sbPbHfd3HHZ+AC4iH44ITDZVOmn84I+40cuD2VglbVlp87nB3oWw6J
mN6Z6oqwvr/FxKQgcnCToNxuMmZZioj80fRZwpi+ksPcGyommPXC91nM0izh/QNA
3ATfyhxotVoqFnefcGeWu61y3IvIwHmKMk3XjBgyNlZqsZuwalOrvAbu62GfhP4Y
MoxdERd0Tb77a/dX+WIThyU+20fkEjm7KccUn1aHRiLnyw8+WzwyQa7BVcty6Lxw
KUDoRrIie1BagK8JqAOzlEcG0YNu6zrf7KI7+yycW0SZS1r7Dk2CG0OJyzQnql3W
90lFjgeLXIP0iNnIn7m9ND5oH3ev7cRvnT46CsP9ns0Bp44K+FHTnolrFnYtAiRC
i/sFqmbBKLPOJRWDQ+3awM9u+2K1IqIBSOBwii1o63XTWSG5TA9kIbXqe+0EU3Nw
T6AYU9YsAUVWtJMnMNZaaHPQ3sUcqiJbTkOzWeGyQZgpv9do/yReZEoJ7pe/r6FF
WItVPiF3K1/youM/HL45UuzA0nivS1xQQqmS9PvRkGpXNpwF5a2JDqnZMs+WqZY/
2hsSLOCMvfH9uDnhpLmgwRr3wR+EpaZ0NI7uZTTEZ7fEADo15piuFzSuhLlGFYB0
pRFvQuj8Ek8x9oWgQ8jlimNMl1W8OC50EzNpGoFeGP5oe1JpTdODEyHbbO1u96Ar
O8hJLZL6yEyKxxIPvNpdpO3iti43hgGgdPVcpR1IKMHp3hSCoBRHZvI0etHOqlED
+Gob3247r43j30m2u+E9QxGnEkSIqG6GdjNY9MchxakLDKQEEachpnQyXwIRhob3
sZjTBrCRuoblXO6bRODaLpgTjEZsx9Dg2AnsQV/DAj74YNYGo9LKDHY3QGWF51ub
ATl3z7y76JMEwmrQjjb9p+3DAomsSTYav1rv2VX4kllPEta0OcpCzqlARoDFcSrp
qkni+6rhUWYohQyWNvyr4DqHOJ+xCmawUG+1COk3HlTEnZ+Wodjp4ZJJe3aFFOPt
at7+k9ioHdKWviiQnrWO4mKwhHXHDkspsnxiA3gRo18i04Y73OhrQdk2pgg5661K
zAvnp0GmZWuS50NTaUiRZJQLUa6BQVuvjtFU0+oqdgap5tPLjFSCOAjz3f1RD0Ej
xbigd7rhLHRR1rT/qMffwLzWVBKfOjRvBKSTfEPN2909mCf1CeMcbP1Xea9NFT1x
930mTT415G8zgh1uudw3TL6pZ6XlBda8ljwN/B6PiZlxVFg+qlw6EGRD8pKTymM3
p9/2Da5wv0D9kUHpSyVyJpFBj9DqEM31kXa4/xM4h397IJNOPohn+HtoJM9uPVKZ
ei92MQKoB4LV4L+NmaONrLYW8VaFKJj5CGNAUwny8VHsIsJsX/IxtMxiYepZgxlk
bGZWj8x4gOURthzjHQEqs+bY4QEO9nYfKcFS/exykLJ/AkqxqkSWGcN6ZYQWgGzK
yJLSyJq1wztNvWuefF+Ef0aOT5WxyKFt3zf8+lI3+UCc8l80yy7t6vJRZyfBlZjg
wGqeyAEcDkRajjyBKH8yUd99zGrnHZn31AT+3IveYPRMS/B/i7HKiE6pzIAJO0zK
OO6wuAXzGg8qtZwhjcHIPDvNNSNnEs1OBVld6VKoKKmMqLzcSFEOpNGHh3BYrwky
5LRr/CBLK2X+vQTpdXsH4lXIZu2Il6kfky3oD4aF2PcQZ1BJ+zSCoYpou6qIpEzJ
qehCWHaASJo4p2lQBst/xTPZFpMB/gxKpWSEgl8YQC/7hPip09SX5zvoGewHhT9a
vHbQgEHf08COE60bTh/I1sRIBez02Ijmc6u+nqxktCsZK+k5ZmZwioaxUv7RP5nd
xayVyeadrWGjdjf6Xcy2nFNPqdRb8z8sEpD8jyU17M1CB3bRGx18/r52HLNCnEOe
rultYjodPOjEJzir9jiDwqJyNhnUwsaeotVVh1zimLXa8v/ZL3K+u0MYk3HNzIl2
D7X7OXFLd9lTcwdN2eSZj9s9cbZVIbELeoAtihoV0IxxYUju4i8rlP18B3N82WP5
KDDDfsyVaPiEgjvtHfCSdl7c6O3cr7zj1v/h2WxkfiE0z7lkxmX/k9Sx4DFNCUHh
2+l25p+4/JjNI59BNEQTt5vi9w+GUFb1utb+vWejGsEl3B64YVLYbZB4yGS3iXjX
1V14hbeW9WLN7d1L9cO95d7hPBV7wUGk3rTOdDz/4MTSpSTDoffvxhkCfz9XzRsY
vv83bGJo4BNg5cd8IKf1Rp0khConbOycZ0qhEyuWu/nqFeoIH7LxfRn0pXEAItdt
bn9PrZ5Y0DNe+QMXYMvDHBi9snHskyj8xq6smb7IjFrsXEh35YGGfVjvoG0l0o56
Wio9y1vS2x429s2apNi/Sj2cYyGw2Xzasaez57qKWltdBP4IPCGFdQM7IiIovBxr
EZh/uxF51wjj78u5Ly3gmM+9WISg3tcmk+TycLaRqUBmvWstvGMmqs40naXGaZdt
WGmurLK8cLIqYUIgtN0JQ70UCAYF9Pf2CWEXPQG4rXXVWn17vWqPuc6V6y38RFV1
`protect END_PROTECTED
