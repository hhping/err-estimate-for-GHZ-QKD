`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJ2RaO0K4+qMXQt0YR3DDITUzldKWHsVbPHiHqJr6rrc8IIttiVemv8vMVAtNVS/
K5+DcMWN9F7o9vAIootkspqdlFxz/VWkg3Lh/c5ftgN4TgiNU5Oh9Hl3K2pgCS+u
9t53h1o6SkjYgNUNQTXu4NsyRepkb/Qb6rtMC7T62Q8DtmMkwabTd7h4o8A20lb1
3Kom7/r9VJY9o0gIKy1Bo/k3Dr4T5Tik1eb66evlV5sAPx7IzDWAEGcX78ED2m16
99n6HbEx1bJvzYZ+3VOKWw0Sqw0tCjHKP/7Qes+YgZ9lbAoDkk6j1dR8fhwBdcuv
n4dquPKgyYiqQ0sWTYsaPV0PaHXeV2uJ9VV2Cq1B0oYfiMNTyO0eEu5hIMuj/1Nb
5u3ZyGpFre/KE+fqpQslFon9VAroh1h3RK/j6Z0dwrE=
`protect END_PROTECTED
