`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWDenP9jW74B+KBNP1DbszDZg/8mDN3ug6naSELegIQ9ZdBsVqjOLh2x4ER1XL40
EVaI4IEVh6QriIdha48X/ZyjyZAG0W1a7VtgMgZBE39Ywr9cJXcsmjFRqKEniUUV
wx4ekvz13NjA2a5by+DsHxybgZmpjM3HM4BzOxcEDoCKBmaakXP0uZHSgu3nGfNv
fmI5ubaFSZBQ9CyfGcHI7iHYuok6F2f/cW1T2YYG557DzMW2CeS4AXkxu9XTTWxU
gJGp9Uw1328n4F+FcNx4lydDTD8eynU5KaJtR+sKBTJ5w0aeyS3i3gJ/+YUlBCz8
ZPTjKpiJdd5e3JDCLAuCNSSAfSbqyZl+9aE5FxEYpnV7Du0B8pLiWx+OUM8NV1u/
a55x/y6qVzlUGB3IsHeCHBNzXPIfrDh9X+TFP1jLXH44m/46hvkJ4vs4we2GXqor
a6a2z0oWToLs2i8LCFHHBFVChpS7H5aRbW85rdDps3YHL2MjGPTW6ydxCo2jvqzW
8cbJVqkasABXabG2Lcv89HVMIE2MwQaVIFh7MnzObQJxHJyH2Nj5II0ykH+2tNpB
ibwDxwV00YVePd1xyAJYDKHQVJvHsBtCxChNqA/N1DdhFTqtHWmX4fpI1FUO9xY5
ret7PDjmWa3+9W/V7MCdjm0FCWPr0xG0RIe24Xx1KGBaDfO7e6wFr0AvQO8pJqm3
fKSXHroV64F8mYLm4br50ErSh8+lnVUyJygx55/oIodumKvnbIBmREn9g0xeO99I
ZpOKVHw6Mq5xOaUxvtMR+o1YUkqMG6fQ/g06mJrCpsO6vSyQAOEPKKexra+wSsN1
0KeAhgeBiFCuiikm1Zp/DYamkbozxwlj6OHDBuH6L2rcBOJTJs2UtsmoB5si3v7v
E1GLyn5Y1s7L+INPiVvo/S97ly9cXRXF4YfZoAH9E14mnJmW2ZeV87npWkaj7WVx
yHUNfcSMv2hDkrjY8vUq88qW/WBwX3LT2rtkfLYyeQIwOU5tkEHc2zDYuGVmiPzJ
`protect END_PROTECTED
