`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E94ZWrMniJ2z9AH+CwYoPgONVo3oru0W2VtB83LMwyW61cNCKU0n0UKj9nFUs2uI
iq4cccEKCz826hExr77F8Ze0hyb/xrcbBoqRNSfYAl1NlmzmCCd0/OLHEQZBu5yh
FwjzKWFflCrDcdivrprnQWTs78x9smVLrnsjrzWP5M/7XHeuIhWh3hP6IHy6Q+KI
Lpn/grs92uGIzn7iXIRcK7KfaLw3NiExx9tvJNtM1I5TIV7WBwh3fYeedK2SMW2w
u+n3/hqsy+3sUbeqWhuL4hZ1NkiyN2+3Ymw74A1qfYEUQyGZIpVk8elsSSVeDaF0
C5b/zwkzjvEVWBAifTxHSUSVBueRp2O8l13zmyCQ7aEe01qfXyoWEkROc3CB7Ps9
/c1F0bpNMYPz9JAy016teikryb/lQn5szvrQDLMikEBqEOa5RGdHjFVciO5VWFu2
tnTzcL9mH+s3QnYQvW+MELU2jNRy1X+B68oLQZUwzm0=
`protect END_PROTECTED
