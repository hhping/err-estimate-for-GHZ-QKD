`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+CDcuCKf3FnJNTSD2KpfmQxcZqdrvVJeHy2gzef3xs6/mB1cUpO9jMLNB0qBI+1
/c1+ANVy9c7MRKyGt80lzUtj28d9prDpKKlHPfxb8/tliMhGMlK/ef7gXmhMN+7q
d4t9eScF2pQ9o6z3L1zoKCkDmamy8pLL7tY+7t7SoAe/+ZPKg58aOXPnCosKF9ln
cuJ9ZqYMpif8IV1ovVRqhAqxOzIJEtW+bDmGo8r4CU52EQzw97g4j2200g0F6+Fa
mA20OADc7XTnjtfhlDuUpcQ7YSLPJsfcknw/xgQBu+wwpbt4pxaO/pYpmXfKieT0
KoYRAN4jCR8Ul6OU7zFrKDN/AVitr0ENlr+7G2gijO42k5MCmvUsWk3zF8tpSzcE
IhLlfDv12gdIoRGyyA1fQdzcnDa1PAq38WHKLcDzGeK8Y/JoZt5aqiCEwKhokVk7
mNgFPOpQn19z/kLeXBb32jKSko5JbtKU2INbsM/DMk3UYjxbayva5Zv2fRAyrhub
WcXuZA3ar3DWlurHSwv//EQIkU5z6MHzOqqQdY5RFJ3/yyj9kgcM0fRuJJBpLJZD
m6psu5Yd2Sbd80Goy8AfxKmZ/4TYieY8BZjv0PHEnlw0wt4ImnQNAD+tPmtzfOej
WkwWFW3p4zIudBBVBqc1SXKBwb+R7+4Ay3SIr/6Fgpc=
`protect END_PROTECTED
