`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sqr6of7nHaUDUE7M0B6EHpDPeOcJvJPyiUaJ92wfk/FsjXqPe4hpA1CV9N/B5ror
BQIfvCrqWaLz0Wnu+nt0AbqE/LzU/agvFXMlf9wMhqrjQgwU8G7jO329iKnGU4n3
46WBgfQNSiuY8o9XWdPtriB6Wydj62Of58p0FnNT+xzsac0T1skaNDRwg32hOPQe
K77E+w/LPQOQDWtkFVy4vhG/LHyLNPwrwTgE3wolbjhFnizIzX7pXafto8YiqxV5
jwXVDTSU9Fx/TbcDsWkO0mAbqWi2Klh/bUEmfiaAQ86MqVyGncaCrPwWyXO6o5fM
fRjSF64inqDtl+LPkC1mY9T9Nq7h2Kwur5GDMY4oK1M/4qs+IrnZZvs1YBCwh9fm
d3xlp+JoJXuOFNfu6uF1fTK/o44cbqwP4w6gi81VDDwW8m62J1trrio0izYg+388
/AjIsOFm9JAWS0OHKULLSzNpZwuwqxkqDLV97Dr5aZ6g2ACvOY1MsHiAXazF5gQ8
IiOfwWFdcATfSWGediKCBUC1cRTCUV14Dg62XMoo7DPsrwjgOV6Hw7dQIKUtGEMT
htCDXGXRsxIwLrsnxZXPpUvh1F2tEKva1BilR688cFx4s95N7eu7YDufFIDLlTRH
THdqmgpysEWNEmvvQML3tg==
`protect END_PROTECTED
