`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6DKcZC31tOtNgD99KB+zMbpw6czYcW1WtBh/y9qARYtO693AlnrFUurDQL/NckFt
DrnRsazBUg+FjJ+uMjmlkgYsVHOZsMlWg0+SR3iLNda99g0F5+T4302mg2S77908
y4/BDup1bw8SNhw4v81t+R5Gw4tQ53zGd30PK7z0TfKKpB6vo6ostatscnI5LQpb
v4/E/66CchxhOTAS7rrESQ/Krn2fGRITVuMPJN+sJXL/ITJxsitPGNExruK1nhvW
yLR7VJduEJS5lhIzbGFj3JQ6/I09HWkFj3FV6yGPcbarovfftGmD/miplebXxFF2
YySxJd3GiYx2Im4rI6njUbVYT20i63nzdL35EdaXQHL5TWksNQf3IixnOELsrKMm
xUDVF45zFw5CQpW8xtYTuvAgkk6Z6mjQ/TzdBGDdCPAF7sZkSUGWxQLS/sqxQ++1
y9GbpegYf1NidiZitqKLeQ==
`protect END_PROTECTED
