`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3DuLndUamPze8dRDaXYSU6oYxkV7Kizil/yQ+Gyr/hp/ogjV20G9ydkcNrYmsQBq
WBxi52ahLuRFN8msDGWELe0kkd9uBUSYB+Uqm2gGSAadpQLm5wFEjd9eKbQD5v+x
3H929g1UYjEFeVIDsBAIST6sU65hqsduSNO8yXUYvnGM9iEh6UrVNPfyMYu2IEUx
8m9xmh3kQcY6hzu6/FkveZkgapE13wmJLZt73r6dLDx0bHtohDXaxP0irykAMQGG
fZf4j0yux1FKtAO+pYeQG4OG+wU0W5WhmPiVvTKD9cJz1PuYHs+2f9KIrXv36epq
EKZe9egUyIABB5g5v977hCfiBaaeQCc4bxDdAg1mF3Fbyuy6KrjLMmHaLigFs53J
gDn10+xwnimqf62mHi6ZMrD5Y8hZHheyZrcymfzGkjrY2s7b+8ca6+96+MHYxtv2
fdYBWhJmnPR7hH0xP5bCcVLXY6SXX6t9slV3aIovuv3rwRFOviQ9PuRRUTEvAiwO
xK+RTS0/mhk+VB1zQ+DGQareB1Blr0YwmNte8SNhgeU=
`protect END_PROTECTED
