`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0rrvBFIKpcXyHVYwM5HBWTj1IRn5MFOnfivO/6HV7ZgaEueTZsVsij0PGoQ1K9k
Eh5YMFL9/4BYLoSnRT/FMvjEg4RaKsazltSwUfTBQaj+deHtfrnJ9E2HMXso+Vx5
e9mQVSJK6+GoO37WogQsFt2opgVTC1PG+yZ5nGmGrx6WG1sh23/CugfaMHvchHi2
AGfnz0FyVP4C5/ZpHdYm6LPPXkUA90y3G7xbnrPI5vqrOxuONM4bfhR4vvZ00pA/
vD/C/uSBwnc7mtC8wXM9VAy/CLT9iUWekNjRaCcvV1w=
`protect END_PROTECTED
