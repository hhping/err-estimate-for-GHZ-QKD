`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
723b7kInFoIwe51YBA5sZu6NX7LEnrStZYQmo+++u7p87TKPlNNlhyVMRGX/pTiY
D4iJbsj/R/qjgJ4d/eYm6ZIYWv7ZuQtlp1atm9lOJ9e3n8snpPEbS0OVkaCJr2Da
de6Ln6/qE0DXRLcfa+WVEdShNY2EHCA6xlf2aW0jT8l8/P9yuPZVpF/nwRXuQcj3
RSepl3+BHF1899bgDww+GUPumWFxyZrsmKcPemChYbilDYnMb6cbtMqMx7UMvz6+
5iDQXZTbxizdjvx14BDQQKGJVfIpFPwxNkZmw8Xzofyxe7HTA9aduBCIAxo5bUfl
AWUU9QueASU4A/XWDQnaWH/EEjvFiIzAeW+KhGORsqBQpfYHvmKrAXLubL80ya1w
kh46WiWQR0je+zfk4WjcubmOmSuE6w9vo2Q8fNE5T4PqYgBW8pqHuK8qstFkMVbi
MrqJwNOs41AZlF+qHo4rZn8LrGRxaT07nni8Ahi8a8JbKFf5RmPkEd2ZfbIP168Y
yIl9kVbMGKoqte7vDFujQZJEDx6r7woGM93vxyoVGO8FLFuWetZpfFEEHHth+vca
7i6IVeLoy/b9CzXJ5GGOjLD2CdHpy/7n9b91oQ2nCN9HCpcyoMOkOg1Lcu/LGDWH
ZPcYDNoNDFX9zOqHFOHKaTwaDTGLIA0Yx7zTyGrsKFFXP3zDJyT0PnkIVzOoOp/C
xQX0m11ZWiQzIffXIldKdqH2qRCo3T+C5ONRxZGGafLyGsI3u30H6Rx+DtQCkaLC
GWcDC5LX+El0uNWAiTYcV7qSDxyzBmLTilg3Yrjy9m40pg55uJLoDBJXglS4WnJ4
2DoZIsScU2mQYyHVmmNhJxsCCUhthC9xUaHwuhHYOP6HG8zNsU49yKYn3rNGEw2z
ukmUdqlBdzKmesS7fDEZ85Sm48wrQY4M1DfyMCiKpa6dGSe2oq23fLgmVzSw2rh/
vkopIvHzhAAao1vEACHfzIjgbePLBN3gi2nLmft3L27Xz/jXbTo3aB6VNZtVPGeP
aLKfSxBxYEKHUzRIghKGIJTXDu4yxHDcJf1UaN5zgoGa+3V9Rs4wzOHfa9VHb7Hs
6ErMSkuEif7tgId037Xjx5/L7OhAVXx90EsM9rDHAOmdc6/Qv2mGef7JJ47/Gie9
XxX2b7eyIJ8N8PbcrAjzZUaNgZEOGY7gSBWPJbeUUZp8u8uajcSWnPRu08mHghK6
`protect END_PROTECTED
