`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSTH6P3md8SeIk+XC22eHJivTb6OEGdSylsatjpqTsfQtc3U0el6HjG5IdH3yh1p
LllvtvGV/f/gL3+QbWeb295lOxIZSkGpG8dXG2FkY38fQa9ElyGbuNgL51hUFB62
3bzgKSlh5y+ZvLN3E/Fl3AhMU7sFdNn3j0pKnOiHLXLP4wWlsEp4B2csXgpQTkjw
hlyVW8IRSORfqsKc+iPt6yEFWIMBtHteOMiWsJCH0+xjRjQrDnsKUQqil9r7nnCm
rZ+kaXc7N1UP2C4YJrPPDVu/lo69/nYMGbFYsiv4nABFbApKiO8Lw6RWXeu1cY3Y
nE5F9ZAUoFkqpg57/QQq5uiAVqCwEFMLTLoZDcXN/UF1oJCvpcH4PUjY1s3YBbI9
R9J45mwUoHZB+rzbCVaeYDhGn+yUz6a0yfWZGNC6LzDf/KyAaWTUEgZAh5Y4HtRt
Sa+o1NIjscrRmIxkSSxzO+dmEBq54f9cn4R1dWyYuInklzT53OfKtuY5asmVRhrr
XzWF1wDQzE1AA/qbeHOww7fCrop9i7bx150qTGiz0RMCdbmBxUjOO07CjYXrUtEk
SXwPt2KFavYfbwynMn+RvKfrc8vjiR7XSwMU41mtyEKD7zVwuoW6to6A+G2M/uYg
anwebFtSpXoKkhqy+oscXA2Ow+q9XSeFF1aLyyYJd6uSUh9NYF0g8g0dl2pwNfLh
8MoXtRRBQ/El6/ERbvGH8jaX7GXOwppPip2wFvsRl8dKUnqmbAjWgp3wBMn3pyZJ
vfGeLOn+IjU12aCk6aRo6MUcFLoMTB62u7Trg4CHazrCz1h4lE9yRbL1jpGSXEV3
UHqsOG5zGiY5nWWcmcrXIaY3YAF2BRe2NlOC4ajQC0X0J8hfxl4g7R351QDczed5
TqhXAIhSJqeXkim8W4flQ1JaEBCcxCAQ4TEoV8Ez+11YNdbLbbmIEUjMShMhoDuj
lk206cbkrWXvrl85VmqEukVI8647zeGBmiBYMKbt5BOxqQxE7pbx4hgMZQdXq5PS
tXk3xKZ/ZK5qzE+0TGJqL6ZTmYRfEm/JWaA8966qjaUPW3prPFllfiM91pvsVyLp
X7jhj87W/VUxhvvbFwdqb57aoCfH0D+4AEOsSi4eGKKIeS8vcCjZ93pGUlYIoEFQ
QSqEiwyYAnmO4AKLNcKk1lhBQBiRKXDVZuqLhMCNLvwwesv//T9PpVeP6lOBNaoV
y7g3CacIUiMm5aT5Zhvg/E5Vrv9YCZC6Vq6mUHjnlbogiD60ahqLqTjwkBKfW7+D
sXKO18/ARorgFL+zWiUVUcLeO5TOihVMPmXtMTNyj9RUWQ+D5lImTus1IPWzRPr6
u8mz49xYCM/meAJN2UVoFCfdhx1MCHD7fHYnyria2ZgTBYGaWJ9vT4ew+fYCmWZT
Tc/G8AGCXjQFhyWGzWyRuYcNe+Ov/AoeMR7TSZYxEMqWPyDOFO5otNP62ts1fVT5
SjpaxNVxgCN5Oci29wXEcHw2Pvku5/JY6zFegMHabZ66RgKmGYuGflgPbN2IyHQw
uev8kch/7AGE2ct21h5P2Kaqa4k4vjt3BMxKpEtNWqPKCSXVK5uKyjACB0ObrTkF
nFa9ozqGSD5YQRjdM2fhOsnOvp0722cyx7PICydVvVp2fy3pKLOjH6GzV5Az6LMc
WLOWE42WVTaqTuVLP1GQt8xnNSKakL3AanSsVbNv2P750AePDiPAsEtgs3ck2Ofu
6jDnoJKQBsYc41EdnZ3k4bqxLJIX7IBgjTQpUvGYCzbPMDiqOAEpTaVuVydhNS3X
mPi6D7hSV2optf8KApiAGYNjL7OkKD6uvh9V8d4AtAk/y8maVIrMYmy8Y1XZXxxA
Ub6xtOlwwdnXyy9U5Z9//FxNYE7XpBMQrog7UNyJa5tYUHnZvS6t8bISzpgpmJMd
laydzyevCAggm0cLbhnNP9lHTOF5KhXoO89jMAxYS/3ym2RF5fiE3MD5UiFq5PsP
V94J0FFefIVqdKgJm3pJwkR8kXwcA6xmNuyETiW2L6PWpPWtbREKeN2AL22QrPrw
WRLUEtatsny7SrdsvhWrgoVy3ukeIi5OFoAdpH2HGmeNFkILfTCGY+8xCKVsiTAx
D8R2Wl+wKDCN5ydbCDqOViwzaLsYv3UH23qJxhb0L6q1qD22xfeHv3g5NFTllu/B
CYgp5Hxhswa/8ZuJhLf2tyNDkQEPLPdRgquc7biZQEK4jsUqtEh1l+RVX9rFpDSX
wQfTPB6q/5TR47Zk/1lrIH9BwQkYQMYIiehZyC1V7TpPuO7qNp0Pgm9tepbhuCLB
rwN1BErOJ+71zz33DKWQ0OvzF2FWx+o7c5xa+0gcvEVU/3u00loV1ZM60ZZPV2pD
TfPXyTSgMPdmfaeMbZbDZDOxIDivt+1qQoFuY4PzeKSTAn6Y1+kfrCNg3RREocBf
u6uwyqsdVfVj1PjM1BTr+Q/H11EZ4sSaSgdpziJQ/KL2sNP8kB1CORCcbatMKlFu
t7TuHzercAaegc1aNGGAzEZVc34sQMk8mndLwXSxgn8gy8D6hRl3U/tv3tIPmlw/
S48MWHD6ULiQlOHy/BBcwWXG0tjbe2Dwro6Vn5pxUgusKBoz8kWixV1jmm/oOyeA
JNBXVmnU5CYgMNmAENBl8Hr7qV5K6/Kzr+iNFI99J8AbEw2jleVQPazuJHZ1JQ7u
8UDCaOa9oBbejKQURNUIsv9WgWuV3YPO1rGa+90OgMTRDpMfuWfuwSoR21g5P1I5
zTMhSL5Ed/aGIQ5xD+TELmQow1xq08L2LyGlSmpE4kW+ucqaRGYdTyqqkW0KUR4p
dV2qQy4hgIq7PpoBfLT9xrRhCXANnp1gaVzdEDlMPwFCztVxdaBuoUVnLkTf3+X1
uvgqXIPPLJihOPSEYopewvIfZIXYXSERXROJK4OH2uGn7nkm5+AxRKWbak9Wpjhi
/mPmr+CVbVF0nlKk47ZyvpnEVrCOWSGeS4+rOvdOG3O569f3g9vdqh41e8sJQImd
ahgATdQ91zy/VlF0bdzxvTI5dcCbhrqI2gUJhvTUmqsJERzVi049zxPJZQLOtRk8
dHh1O853IVu6QoOnIXLboB+XkweFhXyvfS0Gal/ks2FehhW50Hf8drUm8np5rP5/
DcmAr3JhJ/eenPVSy1QbCZGnZBx8r5/ajzpXHgswUVIyTEOtHS4IGnc7C45tJEyB
h87uOLekFe7GZDIPZuzTzof8GKCUbJWWcc24adLb5RLb8SvldG3IN8CcNFMVtb0W
iOMzg8fCAmUHVJeF5jHEnUnnIJHbv1bQPeyzxZeSNvY4WNa0QofAmCdXc8DttZfI
nOw/8Yn6bEQk6G8oM+MNQnoHI+GYY0M0JStkeD0TMFez84U7pvSt79X95F33PE0S
9c6lr72ODFVugSUIVOWq/Wt5vv3FxSi2Ieif2SAGdcORo/korudQKD4rJjd3K1uo
nqZItejDsBQCCnRg0Los5z/pBB+Hq5QEO2nTk+fkIThRczt+5lk53xbInOWM04rc
jqE+HOSWoBZYBjpHmyjOwQ==
`protect END_PROTECTED
