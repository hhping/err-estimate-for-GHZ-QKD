`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q618xIvo3mcP/B1XZZBXCL87m+WOZU6w6ihk2ILwP4xIp25G2wFN9DLY1FegsHBV
w+IoHodednJki89DZPdO5q0LEMEQvp67ND106vpLaBSgjAvis6wBfAQDFS9/rj8N
f50Ux7oSJ5mUv/qj5wRaAg5+LI8DJXZKZ9kHzbKYgu8Zx87+cdU5H8ikOotoeaOu
dBIkVChLB02tM3x6yRsz9NWscarGXCuNiDX5btKWCUOVrFWJpmAymYJ02vXOxRhc
HTtSRmamcmGSQ7p3sLOrOhGSRZ3qPgHYejbWPhnrUhuzSu2Z/RonirFT8PGPr0P0
tgIBo6T43P0VEQtjnKkobgjvtu+aSHrNvzNTA/qKu5uA0gpuyW8l3y/bVKrneQ1j
2T5EYPcYeufoi5/JIMDybeGKlGV0HqGeZkaK5QcUoKq+pVieqhUAh7pM/3h8765r
+WtpRWYOkT41UfFzdfz5OGiQg3nw0EGnPB8bn0X+wUyI+uPkVvlsQ8ob+3NHVPC4
zMmq6AOIpmx8DxBt5Vj5lSb2jEIMIPvt9rB+loWGrR8arwYPw32xn/x+XOL5hDur
HFJq6P51bNikN28EqWt7c/RXAdRvdoLMNjLnn3+fKAtycN7dBZlQ3uTuYb4ZtRXZ
m1KKn39OmmTw85us3TZF5G2IvtYQc6z5FWWQdvTEU/Njntc8cfbjVtjYUQYPlbN9
775qGVZHgFD4QYs7Pd4MRIkgWIHVyQJZG9/0BYc9NORfZ5mOIeFh2ipyvBzdoyoF
JZwT6fotmn0BWjz87sl5f4RWiLatdsr7aoMJBj992/W9tnCL67tpWaQAaPRGyH2z
cxEVqxQcuOf2E10US3k9toesPBTnivutjccCupvXtKdBrOM+QyXlMBIHsXVHcbo1
voVLIU2f/01REOYQsg0pktRwGaGSOW43LYXBKS6WJ4J2VDxQs2fZi/xPfi0Fu/Uz
j/YquYUOhjU26VX82/+gqhwTS7gaHMieJLMzGtYi8fBm0eU9kKNKQyokdOgplUrF
wlTAwo+lugRapWkL6SWAX6RkVdWO9+0en+M55k88wcl0LGAow1714f0Q5cGl3KPi
5YtVqVpAOwOfNiEv9QzeLIMnf4f7XAqJulragAiyEC4bd8zeWRRe2sAlBM9qfp7r
pxb7aU2oWhYCEqaj0WWMDvja480kdmCydD8uiO7C9eexZmImhrM4/F5jdn8X/2pF
ikYuDF91nd5biJ6mU7YcWrCdblcdBbkbvH05Uo1Uy1CTXa+StlD2PrqEUHfrZT0C
qmFevFf8q+Wh+SMzPvrK1h8YNlcsmSO0kQMi6Diwt43dA1JIwILaZu5eivO6S7cY
eGOjISNMgNkUsOdMIbVXrYtyJAIUGoDta5RcMTGpdZ6kSS9PCe7D9OzlW7SfzX0z
cEp2oahvlMDz5a4OfzIF7paiY5qYbQT7T61kXAYahkOQsjDuBw3EWR5I/f803fWO
ssmtSECmPoyFZri1rMWibT1PoBGKed9x3ogbo1pmaY5AIXzr23P6Z85iQ2Z5k5LP
m8umI/BKAd5ORzDprGXb7hHbD/yi5Bd5KQtH2PeiY1d8y874En0LjOywhQihMQLH
`protect END_PROTECTED
