`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oth0ymfsqOTOVsFnOMLN6gfulctjIjeQRgynfBDRzpwhaa+BYykK7ptRkjUdO+s/
PieZmdHk40hlYstAhg5LE/v5PAcC3kop/dCwcwx4xYV8qjGxz4pVUs3h/URat1kS
5zTyZxo9ddRT9H2wsAM7OPH8srGHVaWjLIuc8X/084o0GyH8Zv9EiOKlGMJUx/TY
q9WKdg/ax2+dn0RsFi457BnZT/ESC6y1Y37gM6wfE3o/DhqQtIYkdhiZ9xbZv4KH
wxqurvbJAvJauwwKd1hi7++HYf7n5y2og95j9s9alyLyJCXu3B/222dKoN94by+6
vyB1LLjMo1CQy7+ErpM0NR/R4rWW/j4pkN2/hSHonmY+UYWg2hO3YrYAAa4wVWpQ
Rgp+uiw6xbNn4SUeKyxt5vWbyCCIAp6a5Lr15RL2IWY1PYcY0CzGg7Vf5R6rIOyf
mnboul/+uuho/z3m8nAF+bNYJjSsXC+wBdsgp/SYiv2C7yxdp1JaljNGSxomzB2b
6KxO20Avg0jfypzK1or1VfNDI2qKgAVhJbuW4VtfpAIr+jNDpprtZ59PxeSrH5ik
hHvWP7W1Ac/BSd0kvDlVo345nTv1qZJZujm+0NQjNz8MHkaWQxCz6M01MRtkVIN2
8b90+HlhRUIHgEB7mGF8s/WZ2ECFXXverOXQEpFT7mNiRya42AV7CAGhaYAbKsAQ
hObtwIy6nR8xBD65/QyEsuAfwKYrUxODsOA55d+OSIZfc9eZLpZmqwqGFazL8c0p
z00GDdrsOw85U/hnBszUFYuad3AtF+iUm1shEEhhb7roL6Pa/N3BhmIWrRPIVE5j
BDoKNZmJKDg0gMI+xiWkzQkkYnBMRbHDTWEEFMAoUw2EzgVE9GWeTWb+qaPMSS5M
38kONYsWp9Rno/eN3S79r1/7AsWofQFNU9HNXSlzjJ0MNIUSjvbXtXX2Wml0HHqI
6wpoTIffNdakbityjy4RbcSltoTfJymeBR2BRJG6+Pp+T5yAqkS7YVuUYzhPmqSx
4kZlUjlXTMRpcaTZjx2+YjbWXF/CTetz78/9aGbWe25/jxR2do9bwETaGfaMLRky
h+XAnj+BNKvpHzLY2CaT8yv+B7LIKqrgLvTIjm+w8zdstjo/PDlBFHpgDT8ueZpm
0M117GwLMDQCEAYL7bifEMgmtzSmb1KnaS9rcPwUEAF/+QfNB/GhI8+V0iW52Zxv
T6s8uhRtxg3NDfDyaU70jmeUsQ23vRi2NS716cOlfG4esCSDOxhiTg1j4cOJwNER
bwK68hUulzZVTQ8RKWV5su8Ok+3ymlzqKppMBx+X2zCf1q5rNyYNvredxu1gI13g
QMjobGvqNDzyC7VOq4uufd2GVV7Z1Z0YSngucfaTgFTMCuxqJW6G0Bmqo+pQDxfM
Qx8PRx1CB31cajGrWFogJzli+Nh2InVJaihLqT9A8zhe5YybALTHAU8cHYBEik5n
oKeaJi/pTE5kzEIji1Y3ox66t615jSYM/yc5CB8u9t3mYoXno8NvunA7O8YHY/BN
ymIr944rpCfbdcah1RPldHFRM3hrR55TZhy4NXkfv0ogOo+Iv4K/9lzzIH7Aho5F
NAKd1nhmujE5IBeGC5L+1e/RQWsKuAaJfAabCCX+TJW+CZgrygubHqC1YhjJpPsU
MhweL4W6bKens2yXg7+ELkXOUjJRC4bjtZ7rLaE4qk9Vhfb6Txj4G8omSlBWM7EY
8iK96/Zdv50ETSubh8YEE1WkopNJF2mq909lJUOS5foqOw5iCOMlOHIFBxaGV6/M
GbhdR9b478RHImYIN25I84LGQdgxCL3WHZhATTd2hs2GVjbnlX65KRsRAwJnE0uN
qmpppVzKHr1eO8QqgcNKOtiiNV+MH65F2AKBAzWj0SffzZR6SubgGpuc24QbKd9Y
wtbKYLbqeV6pFre8A6oTPj/OU9TnRjk4kulED67bu+zLtsi6kFS/585sG+UnVYq9
b2Dmcn8vSPLfWI0BwzG7ecaC1pi1yrNqSUv5NwOjlh/n/LRxbgTy38+4WZGSP3If
cwPhy8Kf8sn2tBH4ZxbC3yUg+WRE281WwB8tVR/eijvRwI1asP+JKUZu85s4YQeu
l3eX03TYt/RPufQDHAEQZHzXMsSPbj9LYwYp5X9ydMnefKrJX+YnZHfNhnnDQ5sv
bk819Ue6pYnBPmBseOhOeIcTgOCIIcm58qX0lfv7VJyGZsAW1nblxekpafugquuL
ToMcTo52fGUwZ38WioK5EiiSJxmKDExBYZ696MfbmQy1ntmxlOinhSIcyZQMjKQU
nQFTZG4mlLpXXHNJKBpN68+8MfUAYI4MyDArOfO1qEKNU7OGuqHvwYW5JLD1o82O
3bd+3NgzRcYBlbIHMtZ0vMhnR33A4ZsRyU8ZrLk+ny6I2bMjgylp6toL9OCuAy0i
UmwpEBxs7lYUyqzM+JAmQxXndZ+tQ49FyT6AtEshEpsjdwIn0c52V0WVKzdVsi52
aHaZSncaCN7o+W1ZH+Zk5a+IblUMeGKWawrs1SvVawJrlkO9SxlKLsw4zrEKMO/G
ciCJwidoL2b6Skp/oPdvPcIkSP+vbVX3iOizQ5YUA2KjAGGlK6WOvCoJzkIDRksh
LBvrG3OFyCfHbkpS7GRUpp2yx4OXKRAdTq3tZqUM/UCCmAKZqklVidKnA4bboZgc
RIqQfgAqwsP5hHwqPBMNujwLdNlZOTAYiGz78uvT8O3nsedDZnkvWPcVgobTLvF2
CHf30qmAOhQ1CDQX97f2pQ55eSffMKeab/rg0cbrPr/9+HvUopuiwi/jwNYR9+P/
cH1yr+2KssOwb7qbikKoV3+zZR3nh7As9X2wkCOx8LxnOefKMam0bzY7vqUsZGZm
HyAKb65B38IYajkJbUNfQMxFp2T10oiVuQXXeX3XZRlUtdQ7Su/BP0eCSpYGud3l
3NtJ5cte6qUcnGy/UVSuv5gADQiaqPNs8eFtxaIwv/IJLq5ZNneEPBlhL/09xMi7
pbW6dZzMk2B5Cxyqcxk3bedOjGoQ1JioGmluibrv5XXzsWaqaN/kpiXkqki9K2LP
7dSxnnipeGLOHC0Hq/OaBHO993n99dNhDFC2igGVN8T747nbvj5qg/tFpCxV5q9U
yWsakBTyRZNvJRn+ICsx7ltcs2R58tvbEN1q36XAjemgQFBDJjqD1km//LVeYe6i
ZQYSJeRbf3b/yhelB3CX0ZgUo7hmpkNFdGvKyMz931+3DzD0y+gRUymvM78EcaFi
HhE3SZx8Em+g9gENYOqPMYOeaZenDusN1hN7jpAG29ZE/owrZDnJ3PEhuEkcwzow
IOANUm/pz9J0mM9dWafSX8J9ySyWPQoyPUWNErjdt78kDmcxPOPQFZw4BrSS1Ro1
O9kCyIJwHCeIhI0quUAVKK8Xmv1unFh7h4UIN/QMsBRAekeIKBJyVuJZt9rdECg+
yjfcxIMoBXy10kiussGcObEYjxXXLQ/V1YC1KyZybCeleHddBisAxkrsBI8ve0QY
a0WMUBhMEWV3op9UUdPAUc8Yi0zf/dvKkWngthBkbjWiAnw0Ggvlb5Fjlgvqeweg
CI4P2rhS0uVmXUClXcAv4iRg9C9V+Gz8c9NR+6+gWx3IfDJilv+6A/+eXLeAqbaN
ltt3C/xe/TP+Ixht11ORDV8yJFQm+SFuVX4qnYaOspR+H42i3csQTSri+3NkGhS2
poZExS9qQ9EHgPWiAS6j9i9TE9IAT8/6VYnixMi4CHwzmfT3srjR9SHUeP+yjPTP
Jjfa14njn8SnSKTFBEuVrNOkB4qqU8pHmyZlWLBKeY2kxYHJ6X49oUo3VrACVyKu
PQen94QRnqlSpKWscre7F53jqr7uG1n+eI86ZY29WPNklrdljBo45GxHiTXYWwOF
LkjAdtnz85/vODfTPlqkskFYVikbMs0nti7trgUtaox3yNhLrL89UlO8syz45QuA
PgPsK4d5vEo32x1z1JJHVq9Gau+YvQKQbxHkd6OlaR6ks1XaGYn/kJtbNpzLGOSQ
6V5LCpZ5sWFBp71hMBPI4Hg8C2zHer1d9R5+AHce3MZ1xm32JG8ohbCNIBcvrsgQ
Z6V1vvh2eDAssGmajvPWNXqCtbxgHNtb1sXX92WGydqJQ8ItEb8VAJTNEqLCvH7A
OGJkAAnZk4U08Tt7FmrfRLo4htt6kRQ0b0Y0t7NDE79FAq3i7T79XAHKYeevpKU8
SVDQa/I/XxwtLVUpMNsj/Of9FDOXphaqOk2rrrO21Nu0eTPmDIZ/ut1fAClrFl8j
ZjRGSsZ27ain/8qeuczZ/cEhezXz8RwLl82tUfd5EMAmidWHycFrDCl2XzS7dki0
z6OBVNkg4ua/cF3cW7dogxy3FrckSWQAIdnlCCsdsn4=
`protect END_PROTECTED
