`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1XIUYqli3UiVwm2Oe173GdmHxj9L4SxBMyuqq4VHBM7TDL+SjRQ4D625u7eaZJ+
DAH39q/UaC0rDiJFvDij70qUcbLlbyINMR9ofQ//SHWeO8Ws+RWbC8x2bK95CJ6Q
bLwStxlDn45opQT0AG8J+CglsAoqaSNdCw6gyIjWpJJFCFz9+encki4cuTD8H9dC
YDsi3czhtfhLW6YzsauxclBmHdq9huF1Mky3HS+ibLAjQiec4OCWpbVow5/ypFmb
YGWawqnDcuTdDydPNkLxDJgxmpYI0CoyPFQgU8mg60xHg3OVcS4Wm5qk8uBMIXip
ts/LyBP/zzjawAaH0JIQdnSn6xPCeuINYVja6p0klAhX26FCq5pQpu9nr+isiIPO
FiRj2OaDmrqSFJjT/XfbCv7ECyJozZmW7EF4jrJBDxy0309XHjLkWUUaSJN3IY0e
74hXvrZNrQNelXWsw7sJ8S9pwLd5a+0Rifh+CRC9vz/ZKmDrHPjmH9XY0dYiMiww
MkJCrTVcRT1onLq8+rK9rPsDl8OgWrZzM/KWTKmszXcYvxym+ZsIEDZnLB4zYB94
AgUjkuiUMqVaaKqGY9fJIRXDw3ZOGjaI8nQVLTgrY3xjv2Thfo4tuk6+UQZYibLn
Nv5EVT2SQwzCGfLWRbDSeT3Wd3tf1HQvNCRJ4TxXvVN82m6TYEPM3KAw58tNtKJA
aCxOBmXFA9XseXO3Vyo+EUqZevi9i/yOm1au4Si6QdAkCycvapHZ9Gn+byyAqoDE
oVvHxLOAsOAehDW0kyITtMLtc4DUtVt97dOpxUyA0Wjk97ooP8bsO6tyNC2hQbns
ubDSIan+V1i7jwGj4R/ByyiG17X5oYw7fdQA6oVSqueAwyg6Cm4Rj0BgyLYsepkd
KGVrtcIfJctloIt30L4idcW3lD0gimMrsKMjTYxwvnqmIdstRfAvMzIziD1TVh1q
VfjD9f47AgfTsJQlXlFriSs5r83cZ2OPuDomdpdL9XJ93jCDHN+6toWg6wLBFGCw
X2HoCTxcor6w6wsqtSfriWJwulB+8nPQ9HfoU/JPeVlYK0WLUewuxY/qb4JveAT2
X75Wxan3YeK8r/n9ThZivwafCxUPZSsFx+sqnFDVJKW2+P5iSNX3P1DgbDZgryCz
knaFLkEb5O1ma4FhGgQ1OZKXiUN87S16lbWI6VP7Nac=
`protect END_PROTECTED
