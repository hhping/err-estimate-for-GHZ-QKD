`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V2h1XWCgt260rI9lG7ZIwiIUNCJml+ACvewvzAdCjC9W7rtzXvkceeLyAxphcJy3
GJGMett9yuj3/5J3PRb0e9/uhMR5Gh46YHkKb/Ov6m7miX56tVkFFr6JHZRL1eo4
c61li9DhYQmhDUagaFmvOaGJh4w0MyNhq63+sRDlpA/iuXCwbW9phTJe56xGVL67
ZmM/mLPG0LgP/iq1RFqk/FBzC+aeLkTc7ZEoPJlZUNWcx2muFMIaI2Dy2GTyiwiI
MR3MYL/EJfwXrYo9Y2vomOTyIMkvtvdarKRjRKlXuAx8br9UUceMaioMEZ0qkpkj
M8/vhnjmYBBPyBAFTG4yGaiTIJA+1tm/ONinxJGjekNIZqy5Y2v/qAsX73d7D1ML
26V9u0YCNjcC3pTaJvqKWjuVbK9Ot0Fxw3MGfVlspt2oacz6eyEnZhl5RjXFQjAQ
FCb1MFL0Ssu6HBKzmbF3nf0XGPa0G9CmNH74Z/XfYZJiCC9/o8AWudk8ZGMvHYX/
0xWO2dViOt7UK6spqJEAakPTwB8BLTKuAL9KJFr34P0KEIxE4QXKueRVl0rCgV6S
xbvXqsDoQHgx6q/WlSwj4qQMB3VRhha14TPxWME3QAlbB+Iyy5sx6/739QzSuw1+
e1rxB8qKgucr9jSI1mSVLq1xi7AfvGVSNLyMlldAlezROBEphIWjAF/p6h+eAFdd
S38JCAahOOTyY/XYp7kdKbr1s0EZRE6sJVXS7EV6c2d7ZwAdoUuoqlGDG96vym8y
Vb70PA/IRWa9tTa4vOWnJk5I+lIe8YJIGFT9plscyK8hDEDn7S7smE7zVAKiOeyj
n685wlYp2qL8FgFa5T+Ry21/SCHXPAxNCK2upqgmbwlWeSEuGP+ZrT6hMhgKnenk
5eWnIG7TxxzHh0ZJgUhzFks3anBZt4s9lykjQ3VbRaAvHlaz/ZSxF8Anop+Zq4XZ
`protect END_PROTECTED
