`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwxsAyQLE8UqjUEpTCZWGGoTjLdpXPp4WJBUua6H7yztPnzIXvVWpoeefxZfKH9+
8CP5JE+PVvN+lAiQsUTIteTRkIcm9R65gt5KUDl+U8PiLoXhsCMLLT8PZIvC6jbz
K73JodreIdv7UY14GAhQSizv6z1zZAwpYumerZiiC5Zh90Yfi/xFXrlNumBPudp6
RyFat2cFr0BuScubrAJ7/GKu9533zK9Lx1KSn1czBCOUhgDg7Oxb6t59wHq7LCHX
dK+5HOKaG0xYqKPX/qNWsfc/crdoSvaQDP6/opHQ9eqWVbyy/qjjw0Eoc26MHJxc
ljyfEiVd2O5BNmpwX8KW6bTBZE0GTboOsv1t7BJVA71erF6JQcXOvDjAZSXGsIKi
Zr5NKNnU01x2gICmKYWypWL+LbtFkZwZ+0E90SEWfjG4LCaSIEgfWhjPzr/M2v0V
qGVH1Uqza1dmqvPENfNGILU3iMCWaew71l4wlR94XaUdHN46Pd9lgSUD/Kqrtk/A
N1DwxzvOZQtUNIYdD2tYpGym+8jHiaGTt2LB2U/v44tSj0fC9IGcx4xMfw13iNQ7
yiw65WGdgCK2pbBCyLEQSu7dWpOKriL2B5OEZNparXmDyjjkQy7HHO12dGt0rHjq
sy15YurTF/MVHIOq60Wcc3S5ur6CYAmQXfRtbIm30G9voKXJQ3mGd4LeZKHKS0TI
R9mZBGtFFaY6ZbdRiUCNqd1FLZDgkIXvB/bZ7pVnp+VDcP0An2xQ9b7eon9+qtwe
dg/CvqNLPEakMY6HHKHL3pgzKI6nbfeChRhn1DgspWGZ/fMEPNQaFLC3nKo+opUQ
`protect END_PROTECTED
