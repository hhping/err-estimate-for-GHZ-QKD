`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDURJdiZ79rwChDWImCen4sOlFirVXnby0bB3C/5aezJBRt8vuBZVkzQaT3UoONP
SL7bFj9/98U3bbLc/+PQhxv/VWe+twtRzsrX3WjWAzITIaWRSDvcmFj2hxBLZJ9i
s4vRKHTOYrphi5Ofvt20ZsckS9lrdkUPMmfON7F0gNW2CmwUEEfclNWgy5Ygj3fi
NZqFcZVGko2sSzC0NkPhzLTPw7awyEi5+Abea2scOwq+qwunhExnwKGe289dLOpw
uPRJKueIaKTSnUUOQvEO0aBQVkGGhQC7w9NxlM8OapXDBEVqfxi1XDPzIPPgWWYY
Nm8e6TEqRGhNECK/egtsNgKjtH6z/iLtRf4jTHQTjz2i8ns4ThE5IfHJNu1Swh2V
v+jH79tlcZoyBtT0b0nQjKoD+fGoP3/QFa0qpyZ7MrovQm5gAaWL0QAE9Wy1/UH9
NIvLXvfUiQlCSMbeNf43/NyMudRHGc7dfLpbZ/WXESiloGdiohpUTrbe7UnfTN8v
HyZumBAI42R7ZYHYDkXzAj/gJoWVf3Q8f97U6vBrHXICrO0KxzReVHVX/UWKqI58
U90tY/ttudM84fvCdIyh4l4MIRluPqN+O6toASQLEvF7gq8EJzbR02C0VZbIRKzQ
DKagYYWqSeCZTZZ4Vmz4Xkhpv2qWyLKS1Xf+NNouCXN4ZJW8/slncXn1ICLeCf2H
yfoHKzoYoC2nck6iIFhQ6BeyjAOoWSWeKFB7KMJfdtD44AEv3HguchbY4lMtTaEl
fyM40Xo3aSca45EcOWw8b72XdtItzDdchvXYF+W6pZqFFUREd9UefODlUyjdXy4+
cHINjt8ddbixDxzVf3jIHbOXM2D9iypQnr7z3evb+G+I7sQOGhnE96EUqXWjF6++
fk2FFqZFveOV7u5h4jStqJxLjtoO8bAcg17Zue6nT/4=
`protect END_PROTECTED
