library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_tx_cgb is
    generic(
        enable_debug_info: string  := "true";
        bitslip_enable  : string  := "enable_bitslip";
        bonding_mode    : string  := "x1_non_bonded";
        bonding_reset_enable: string  := "allow_bonding_reset";
        cgb_power_down  : string  := "power_down_cgb";
        datarate        : string  := "0 bps";
        dprio_cgb_vreg_boost: string  := "no_voltage_boost";
        initial_settings: string  := "false";
        input_select_gen3: string  := "unused";
        input_select_x1 : string  := "unused";
        input_select_xn : string  := "unused";
        observe_cgb_clocks: string  := "observe_nothing";
        pcie_gen3_bitwidth: string  := "pciegen3_wide";
        prot_mode       : string  := "basic_tx";
        scratch0_x1_clock_src: string  := "unused";
        scratch1_x1_clock_src: string  := "unused";
        scratch2_x1_clock_src: string  := "unused";
        scratch3_x1_clock_src: string  := "unused";
        select_done_master_or_slave: string  := "choose_slave_pcie_sw_done";
        ser_mode        : string  := "eight_bit";
        ser_powerdown   : string  := "normal_poweron_ser";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        tx_ucontrol_en  : string  := "disable";
        tx_ucontrol_pcie: string  := "gen1";
        tx_ucontrol_reset: string  := "disable";
        vccdreg_output  : string  := "vccdreg_nominal";
        x1_clock_source_sel: string  := "cdr_txpll_t";
        x1_div_m_sel    : string  := "divbypass";
        xn_clock_source_sel: string  := "sel_xn_up"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        ckdccn          : in     vl_logic;
        ckdccp          : in     vl_logic;
        clk_cdr_b       : in     vl_logic;
        clk_cdr_direct  : in     vl_logic;
        clk_cdr_t       : in     vl_logic;
        clk_fpll_b      : in     vl_logic;
        clk_fpll_t      : in     vl_logic;
        clk_lc_b        : in     vl_logic;
        clk_lc_hs       : in     vl_logic;
        clk_lc_t        : in     vl_logic;
        clkb_cdr_b      : in     vl_logic;
        clkb_cdr_direct : in     vl_logic;
        clkb_cdr_t      : in     vl_logic;
        clkb_fpll_b     : in     vl_logic;
        clkb_fpll_t     : in     vl_logic;
        clkb_lc_b       : in     vl_logic;
        clkb_lc_hs      : in     vl_logic;
        clkb_lc_t       : in     vl_logic;
        cpulse_x6_dn_bus: in     vl_logic_vector(5 downto 0);
        cpulse_x6_up_bus: in     vl_logic_vector(5 downto 0);
        cpulse_xn_dn_bus: in     vl_logic_vector(5 downto 0);
        cpulse_xn_up_bus: in     vl_logic_vector(5 downto 0);
        pcie_sw         : in     vl_logic_vector(1 downto 0);
        pcie_sw_done_master: in     vl_logic_vector(1 downto 0);
        tx_bitslip      : in     vl_logic;
        tx_bonding_rstb : in     vl_logic;
        tx_pma_rstb     : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        bitslipstate    : out    vl_logic;
        cpulse_out_bus  : out    vl_logic_vector(5 downto 0);
        div2            : out    vl_logic;
        div4            : out    vl_logic;
        div5            : out    vl_logic;
        hifreqclkn      : out    vl_logic;
        hifreqclkp      : out    vl_logic;
        pcie_sw_done    : out    vl_logic_vector(1 downto 0);
        pcie_sw_master  : out    vl_logic_vector(1 downto 0);
        rstb            : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of bitslip_enable : constant is 1;
    attribute mti_svvh_generic_type of bonding_mode : constant is 1;
    attribute mti_svvh_generic_type of bonding_reset_enable : constant is 1;
    attribute mti_svvh_generic_type of cgb_power_down : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of dprio_cgb_vreg_boost : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of input_select_gen3 : constant is 1;
    attribute mti_svvh_generic_type of input_select_x1 : constant is 1;
    attribute mti_svvh_generic_type of input_select_xn : constant is 1;
    attribute mti_svvh_generic_type of observe_cgb_clocks : constant is 1;
    attribute mti_svvh_generic_type of pcie_gen3_bitwidth : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of scratch0_x1_clock_src : constant is 1;
    attribute mti_svvh_generic_type of scratch1_x1_clock_src : constant is 1;
    attribute mti_svvh_generic_type of scratch2_x1_clock_src : constant is 1;
    attribute mti_svvh_generic_type of scratch3_x1_clock_src : constant is 1;
    attribute mti_svvh_generic_type of select_done_master_or_slave : constant is 1;
    attribute mti_svvh_generic_type of ser_mode : constant is 1;
    attribute mti_svvh_generic_type of ser_powerdown : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of tx_ucontrol_en : constant is 1;
    attribute mti_svvh_generic_type of tx_ucontrol_pcie : constant is 1;
    attribute mti_svvh_generic_type of tx_ucontrol_reset : constant is 1;
    attribute mti_svvh_generic_type of vccdreg_output : constant is 1;
    attribute mti_svvh_generic_type of x1_clock_source_sel : constant is 1;
    attribute mti_svvh_generic_type of x1_div_m_sel : constant is 1;
    attribute mti_svvh_generic_type of xn_clock_source_sel : constant is 1;
end twentynm_hssi_pma_tx_cgb;
