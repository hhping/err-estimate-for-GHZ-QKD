`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhED4ZicuQ5uDyty4Gh5lvS7GTG9Qhe4EjWRX+8X2P4HaARaNdDj/s+RhpTIiThe
H86C59Mevqd25vIa3KreSwhHDO2d6KXc0Ex7HPClGXxxIVj9prBhQiioU2hCB+gJ
RqgrV3RxJ+ecndYbQVCadf2nhdvsV5HrlaRwCOMgo+S4nDL0iad6kphOu90XPpfE
m3DyuwDt1IKbsA9IK5TUM1LfPrso3Flw+vwCtcrNrkgFYqnXVU7tqsnSXd+4tRBZ
c8B30FWpZEBdfLVNtQxp+dS72OFj9XO69gWKNNNs3qG4jFnnSlGyxOYS1wf6yF8k
x6+xKYGkSrCD0QGIj/ANamcGP7zJqbfmtgohOOTyrkgY9tXa6L8a5BizXEIyeqmm
i/+DHt5ttwfR1sP+lAmy+R56DXVgRH2Zqi8Z+IfBMMRmVhtIKlvmOkxKtbBaYygt
t1xNuKTJwO6+hyQKNt4/i3fWSc3loJNNOWXWanmFbxvBb6pEu4YByBLIn+lvOH6D
AvGH5eT5f/XAbtDPJPuqqlLcEYV4hq7VMs7iASbP2GE5hQrRG6GVpSJuEHik7LEn
LvYvp7inaNr7HrQ2JZ5L0GskLnr9EinPYKoqXX94DN1Jqkxz8JCFNinOxjcMmvtZ
h7tVMY8V3QIRsNhlSCqkBuMIw/OevBwHXfZzHblzUtHXRZOGYPEyQwH3ekmB+Hi9
qWaAwqlb6rXNCW54h3vzhR7c+tD24YxxKuNVycflzJ3hvVLHw0O/HgEpqW0Dx5IN
9s2A92m2V7meabJ/0qyCvIE1eE8ROxuKeG6fRd67ewQweAVDmpOA/crnDBckBZtv
1CvLHijaFWaqgPZgSN+YfuZxQIWr/vCJX/GrzauTkWAeOAXp4DbTAKN275tySJbZ
ztGUg7jBgUx+ph38s1uWd7NoXsIhjanTwFg/SAAteyEo4qwU0kvo2IXXBgc5HtjH
XNFCtkBfW6PBjGpASR1CtMCQtiYutp1LcBkTy7qZG5mLuaigBu9D4uvV8UbDZcuT
0uescJD69RP57vpPPPLVYyr5g7+Dkb2nGxZbACKTwZyPEeyf1UszHUJOamKy8tHr
en0LkxpL3F7dCh5RZBPj9OUIOkzVqteO5Verone0VSCRzQ8tdGgYPeesz9DunQKm
vrM9sh+CVkxjluHcGVIF37lpEINsvlH3Qd4+CJ2JB8kZ5WDnMX4V9BgORSIwQdT6
TU+suGj5ccCHCTUOL2LVRSshqWAcxPQR6kjInHQ5EG/lAPLPoiR/jUAQF481pXEZ
J3Pew9uACG9jhLNfAHMhRYCemHTi43WviW7nC0WOB/UlzrBd5m6kna9co6EhiOWj
A7F7WEST/EEpvWerorJhEHChpN75yHHrVLq22rebxy51+MLKqw0PGvZwGPEACcIH
SM/yoOQUPbzDegHeB6B9WMiFWpGTuv/LjUd9oV0G5o9CWX5QHzVDO3/KHjXKfUrB
mVbjNcz3xQUDzaF2tulxJf+bKQCkLLEQGM7HT6lSBaLCd89z48rT6DcKkzyLkwJD
KUoYOxRydUfjszKTzE1qUJ1IDFo7RZhTlPhgnwUoyhCJPbiRWqjKzDhKFHO0XFbA
0sfW//Rmvk01pM/wiHt9rcfChCDJZ5rwoh7pnR1OQmfwo36Z/wr14FoCvqrtK2H1
g857OX9SY9lBONNd2cLEnUtHqsfdfRfxhLtrc8DFqAHtdgNa2ay2GqN+YQipzbxx
YpvwvoykdxmvJdczrTDIjQ3V7MrHIveouqsd4CBhYGx7BpnH/F0TiD4gB6Ya2bIL
nfAzo2Nm7Z1fvclYn+v91euMYeFVGVO05JAi1EfKAwsYZe6vsGEB5r4lnh8UT+84
MZSME5wISodb8UPDbCW+eQ6x9lxDksUI20L9r/lfWLpSyoAujpcvr6jYvOhxsMUT
2cW7/2dD2mYluZc1l5dQe3DivSrMwQFgZHMctCBMqLoXfzkPyKNvkhE3FsFkNgM6
Mf3CfvgP6vi3zTmQ/zR5yjWQGtn7wUOqx2D6JvMwZBnV4aOsbmwtV8OABvgvUsWJ
HjoqqrMl/GISpYRtSTyoLVTqpd0R69jk8gG60X0VNq8iPkPq/Odg899IITi6CGAI
0VBJVqFHt9aEwk1KC9b77QcKM2+MJHOSG2xh+nueDKq7UG2oTpYhM9pbqBw5FXKU
7yMneGKF/l0EyoLapkNRqm9uGQoiuiO4NLYnlwgjhzmAmD8TjLOmTdgw86IxRMjB
PXT1wvts3qjSc22dmOMu1CegHUaSmoDwyO6Pf9JNY5bZbYQXe/6YpJkwKmBt2lJP
4UhH11Wx79biGR+m9Ia5m7oop0rXoO2SxfpNicyUCI9WhrjlA3+QGMnwFbg2E2/2
TImDUgxEJIcXyW6Vkj1lzuB0QVav5sQvUh7bJYr/H38uqUS/jOspPtldql4SXFyd
VK8E4aakanPOJBbXgUfecJvIoU5ak0A+dpPuwVYopOhT/DH3sSuQW6MWvyLW0/TW
zJ8Id1HtJ0nNk2W2a0Xng9Dpfm0JTradev13sGqDIfUq0VF7F8F1i8pEF1uAVtZd
x7yiGvJ8eDhtqt8iCanFkSAlFs7ABQMeG2h3cXm1JWgiENS0YpqCE/TPwbDopJ2+
EPXJo5T7W+CvYqwW/qW6zf7h6nrQo51BA10wlRAV8A1m442fT8fQZL7Hr7aulKNa
Xk9h8Obe7r5qz8OmjYrjg1YhfcNU2rXJtxsaIH2bH7oUlFY+5xcmt7vYNBLlOwX/
/kBHQ8kDXufN+/xC3z14a+wHyVwvIGXpr6I6B6Wbt22ZL1ucdCyZNT2uJLAfAG88
nW6GtYU+Uc20D00dBrzsvmOkYHaxVoOFjY39iPGOeqDluBIh+RGz+Pqjg89dPPmW
h/X3VfiL0HZYyuMQD0kHAzCT9GmVVmyjI0hQaa+xitHE7vI18gcYxXFdklyA8vyv
+HJjFv040zMicMq2x6vIYvETexZq8zoBrFq2LYuo8GwUMXKN6MGKzmkIuTd3wgFJ
+g/702m0GPNvBHoBO8Ky0WCiIdaRF0oYbK4Rr2MHf1FrLWCiPgPN/lETWMJSCoX9
QpylsHbzT26NHvKUYbtRkZzjhtbUd/l1r9K7H+kXKrRrDrLm3j8LY1KUqQ/A+cQi
n5iGPozJWKIJGMOdDTyx6Eva2ls5zR2meVve8VD3FfCQJ2i1cCqip7U1gKiJys+a
PZEMRvVpSIJ4SkLp0YqoOYdLT/gTlKSx2IWWc5Sk4kpNObVY4JhF2gtjzw2HnjQE
ZxR3r4i0EMmBJsvTdvmU8zkO/Yv4dn/s9C4Rldsv5pRnJb2GppKy7nDYxFJaZm6A
CEXytxHscob7p4Nu3jBBzqNbVQLM6cZ/ntlS42jPY+Gh9RNJ++dE6pv11VaqPnGU
MNGXntv77IPGprQHBSRk+z79gUI29MaRt8WcTwaWXZC1tpA20YMVuNx7p7X4hKk6
VIAx70/C/vR0BMX3GHOtDrgZwWYxq72mDSkfCJUWJ2TCLuK7cD4SDtLsyhm/Fbz3
rH1EJaKrpvWffJKeBSYe1E6bVh9l1TbNvqWqpIsfR+KuTlsYtePZwWQGKSXgeHRu
REGicX7Kr1MyY/R8PXO1rQ==
`protect END_PROTECTED
