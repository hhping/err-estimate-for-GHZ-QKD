`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgyaPcqPwC3zRl8pu1ID85Ov9L1WkY0fXK1BacNC8yPGej+Mrx0+XillLwx72VdU
7jGHrRnw6yxgWZJSPSTA85VfXjHSMUoBLTd/tOVCJsqOOSRHrlnbJneAO8MXrhxC
aS8OXETILUGPQflq7pa6a/xREMQ1YOFCtedPkUP6+aDIfoIVAHlbDKNSPQ0/ymD5
2U0J4Jkk/shbx366ww+yo2ofB1PVfOoDoS6BzuJ/kHI3vGMttVX+ah3qw7379fxx
UPCTMJSN+VkcUgL6UVJEHBSD6+onkdvkz1VqWIWBLqX/Sid7IpAgLj3FBUeDeZvb
VzMZGNpIchj+728tQcYo5fNaoc+1ZmyRgZtTbJ3unWDVB0gYCB2gb3xh0wz/LT1W
bioYmxzVDR4vqNfSMsoi5YulqjK/Bu0lPTFaK2uRnBj9fFYBryWv+lXYaUGWLzpw
yDtpe9LELlsN79MqL1n94qpgnFCMFRGou84dBBN6ID8+dF0zNxbUnuXIK1SQfzz/
papgwjy3F5QiBx76Cds1SOlar6pm3HRi4wSOg2ZtXQuK26SRcpZpMOGi59Gjdqmn
7RC3csHcCzg5r8QdyV14ZKGkgwEp/JGqUB2PmPMaiT7gbgKCUsLabjp10Uhakn5e
pTbsNTpIibeP3D8hpujatRvhERNnEhER/O59qRKEnoH19xw5ojtA75ESEPJgi8XO
w9e98hzgUNqgb8wKDJodOgDnvCCfO4w/CQJnskVJP5R8NvumXLrb2So2IsHHnl56
cbGpyP8CVp8BRsbCR8sY+h9CSybQgDu8/9VtsIzF0y373E7MOEOPj5PaUxBYaXZw
P9c6uY2OceurzThCokRGmoszArRKMkhMd01sLVXHYQjzw3zA44XlhBWnUcl4lmhk
8B5FQtDkREuxOK5VtIuppbsurYchdIpSIo+C/LM89ir2lZdTO+AW7Z9e3W19gIE1
c5Wsqx1fQplGcCxMWLI3wUVwBj7VEX6XmC4dam/zocvNswyEmtryYOnRIU+ZX+dq
M03bC5srQT7swAiVRMbBhRwF8ABjjVwpNLUR1I5lMJOjOaua7WIv19Z1C0w0yEz2
DxgNbo6IQ91ypunkFlhHLLROgU6wJVgN8TQyJ94bU2EZsVGb0ZX6Ev7a+2rdHTuy
LvKWErRNddTqC0Mp9IWtFZrLaq/29rigH7fhd7DbfXjvt1UpvU/lsRvPNcVnL3q3
TS96OGerWoD6z9npU6VpDBySqdy6hBI7iguyMTKaqIqntKpevkOXy22fUGuEvS3w
65BMkPh1HmnDWRa+uWC2v1TosRmud0HrpCqlTM6VQzeouEXZ1GTS02yiRjgXY/nP
3vfFNMI8umP1t/GXqLWmj6IcjlYnjMdjzJB37VhCqZKDN04tUnlsVYJuQcR4YHBE
aZe19ir8kX9Ky1Y6KXUDa4eYumgvLfJoesLVIrKRTAcDsxj6/IbSaTLwbkWKHPmv
6lLmjZi7BVKMLCCRFOH+lxcKkFFHSx0bFGkM/PJiAFn/CjqpEXHJhQUOGPgEf3uG
Rt9oX+XjPEQjMVp+XrARvFfcXrBQvqCtDPvqyaUu/TdJZrlHnnZ1hFbpvrGPZQl+
SjEOvO4D1TNr8swONd0ICMSfYOrdbNemHWiGczH90s9PyZhi2anZflEsDGwd4QPF
gmmxhdwRzvbqdOAEG+4zVBnYmkl5yjMINEHdwhUV792KaGdwhLs9fQkNLSo0Qglm
CMcMdYwU7Xoehu4266+7t6lrkXE0TR6YsL7HJRUANUoH3IkA1qHQK0yTVoAEsyOG
UIDhN7ADGgc3hpBQGdJFCw2vCGntZGP75SUFHQUr/KTF1R6pkL2kKQvz2CVftlyW
DvWNKGi74xXe4S0dkp12uMoZIq0hXTmn+MhIcsPWn2o6baGOxl4CNbFf/Ld7uvUe
wiTMDm+yfGdN1dJjg3AXDYMZzyNrhyvhVp+QcrvEfq79iL6cAW5ruJk0K/7Cot+P
/Aio87ATibZrFG8ydeeNX6rzO81/RmaVi4DnFmKyt7MCUUr2xZMZYp6k+jphoNkK
VtLZ2ppoL4IeGb2LfvzdrpgMpZpKRHAoV+FblV4o+/Z7huT77ZJoX/pH5MiVImP9
wFZpUZDrac9fTd6EzjJdP6bWjMb6CEd+BlrRpoxkmpW2sjaT90zLt/A+NNjzMSux
BC7cVUaxejDTYgPd30SUFqlHGuVqNHPjW2mnBDsf1Oev7egywlC69pveDZJSNdia
IY3zOGbjzxA+DcjxcNrnl5eeRm9Dgkvt+4YPpjOV88q9cZq2/u57jyFk1VmH2yLK
mlG/FOQqq0+hFkPHjh9usSErP9akhBj8Cs3wEJCeGL0DkcpQiKQ2esj6+4iB1dSR
+VlqZXAAzGs7smK9CrgNHXpbSRsrfLY2Xj6AQ0oTnZuCa3yvMyNDjIvz9hDP2Wd7
IaTbgMWek6VJCH6S1nRAfXOrHQNtN5IHfSE0utTf/8anpjVTmtPpsWQGL0xXYfl0
DsWGE46jhjezKACw9SUtZKStFYjGqyRSvVQ1xu2TP8Sulh/dmsg4qWnI5WpHIEq4
7Gi7GnWSfPFFW/vxXLlziASrSTmDyjO7hNbfD7oO1UUGbk5AGrjnkEXm2eIoMi8C
dWPVc4phateBXlhJItcDqx0ZcsY709HJJFUNynJgH77YbN4qSj3pT+Bcc9r4HC6o
gifMy3c+zSSZgAOsxYxWqXBSMEHZ6/MvU5B6toO1KhzjTjzT9ukGCKmXgZyTG9kE
S+m8Gu3nH3F+zby/jdW8NgQkpIjhaipmcLZTWy+jrfRCXeCjA6dIbnGFiimE/S1s
7gnbHGifXBjdf0wI6kLwT9P6x2KPACzUGGGddIT31/QAOWiTqMt1rlBk8ZJ9KAKD
iV79S0VdsTQBjTZAlTGXQRCPfpkHqKHUi1AMdmY0gGw7QufkVDMu39ZpDYzgsMsm
YnzXTeyNglKBbjykTT60ITbsty1No7qpLJqdUKBAGjnSya3ePzW6lcRT4A3tgoif
YHidKA88Mz0QR+Myl4mU1GH7qIazBUYHbK5l29hh0ZeQ853q3JZdpsZ7bfNk7Gab
QhJQNxPRmYFOmDO6iZrSX0Ajg8EGzgnluHEPbLjkeU2E7CuU1OyFknaynRaAMVhn
m+YDcyi9n/d4z2YUePpeyp5YD3S7rsRn+0PuOFiA4Z5nvitzrdKlhGaZzCRkOAUV
VQeWjw2iU70rLpL/dXXOEw==
`protect END_PROTECTED
