`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pi4ZyCVSfKUimmnLSpR8KFjlb5KgEL/shZsTJb4jcaQjBHEYhqP/kmqM5l3Ux+Ye
vAuwZiHD70MDQgNY4FXUHLegAvFm5gcbK5gvi2q0nKWKE8IafoXOnAB89lLGWcph
ONeYcW01D+8hQjs1Kp6UFux4rXaEksk0eGjYtfzTd6rlxF22SLEpE0zh7JUDrZVM
BSRfWynU7Vg9UplZEKlmaQxF2xh2BQ3m6RdnHsRY4fXBgIYja9nfGrfE32eW7j97
I2hoOU3us/Iq2FjqGgoF39SnEWcj3es/bYfxVZ/YGWxc+Juqz9k79R/Zmx6Iy3v1
bgKh5a+IEJeBXwEdU2j95jFE7cPVgSatjCA3V7Go83pHAIOs+B7ttbkh5/n+pJPs
r02bSqYCKb0aK3Po90GcxZhM3Krjkch1UYlgC4zk4roIMuv/loLCLCprhrLhcrrp
WEEQMjaS1QkfhULYNLop3xCYxyoQ9sS9NE/N3776A18Tz+ocP7y6qsIxZZt3JG+j
3TAf/85t5urwvuswYP6v3CpP8LuAs3JbIgBkLvQ8F3yj4wb8Mq2ZpvRHozvqFUS+
F9xLcHm6dELKONHsh8iFYlWPY8Rb9x8J58e9BVBlejn5/qh4niWy+5ZzSaZXsGuy
EBD+AYdVzCKXOlXzUyOCpg==
`protect END_PROTECTED
