`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CA991yD7VVdr47J2d2LKWv6/Uuv6oWn4oZLlWwHZV2UxmdH4hj09L56P2+CJ6J+l
gRhPDFm6QqD3gSf1OM1xzsE9Q2PVHVHGVpRrz2d9BID/BBsaEST+l/vPBZIicEaA
KEZxT7Z6Ake//A+KdDh4thAPjMXXwkf9fIuRcLccvoO0lkz4CCfByfTsh7grL+xA
kKoGRFP0nrHFqm9wmsaLs+nBKdo/gLjOAiwUk3faFgkxObWXZAPsdkfgDQYqvuZp
yNUWB11jkG/atRKO+IEQdCbx5x2Hl+CCu2T3hViYm5H7/9EKc+Yi2lhU0OzGPri0
VWWM2EfcYM3u70cy7spJTbM+QLIUzSJOXjqjz1JQnHBAgBBzXUCO4+WhFyjoExBE
vfmsY/E+1N0iV50MY8iauLwRlV3tU3PCRB35rWKogYlyp78M45Li3UYQU1z3+Qq9
Gu6zrNniLc2pLBOJ87zpJ7VH9c0NaBKSsqYDlSSlyl1lZYyZ0by7SN4OSPlUWCHr
QvBvCrxiM7VpLD0nsz1/GNidGL5gncTMcPKN9u1U35JDXLJ9bpJslHJkR2guhzY/
4S9tRM/RfPvcKEokqmNrB10RHcX6sBOomvUdqlmXHQFdQ/dW9VsDFD9Q1tOEcq02
dydrx6hUANTBg93muMo8no2zCHp351NeiJk0Ege/5G5JR/ci0+Xfva432KtvZAiZ
kDzKecpsMfRWRFFMm6/UZBn3u6Xi2ffogDW6fw0Oba1DJ1mFLIkX1ikMIEyo1gdA
CiiISmeb4Y3WEnQqtgwcRF8UaLcNGW7OJyoqWSKOb8JrAkt66K3xC6M5EzD24j6O
xBrVB+Ji1hiPYuQDHyA8BnH0uoiZI0wXD9mkmK2R9vSTii+JtYdbLwClS4HEQYgH
gBiuS9etAm6oOh+7nt+3bTxmTd0w6WHhnOUJPWlQxeWb+PoWrtnsPsNMjj1WbZYa
b88wFc2pn7CpyM7gLOv46w==
`protect END_PROTECTED
