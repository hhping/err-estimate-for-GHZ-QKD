`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nB71QWNv9AnsHQYHYZsSqgJZnnlczGlX0mqAcs8rmXcaU/ncl1FOxQscmwLjUNB
lBLg8Nz9V/03eBq9l6RhN0snLw2ExwseIV4kEEVERhmo6hctZO3JhWTXzQDE+Il9
icoIVx+hy0pwBBQ9iC20Ja3z4qj2loyxaRK5GjxLPMkpZzsxW4A4JyiYOMfIxsFC
WB8WVSuYinskhO01xfqyh7Qvjlcw+k3cxFK+WYUik8nl1FIy9qbV5VdXPFIuR0nK
mFFYgZ+kSja71IBdiEIydPBtMtCz8oLjLoSAiqbI1uWFmGOSk4lgK+6cCNKw8xtR
Yo8hz46KCTrY3nSFOiShWgDKwTgX1qvOxYzLKL/MqipC34Bm7tiQNNPej2BgVriE
dDstaLxmLGtx++I/ahMeX7xHsxXnyrJoTiSSd8LFero=
`protect END_PROTECTED
