`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Fv6i0P5YEW692GqPZ8MrCNWLz4SyzLihPRtt6SVbYGZFN92k6liQW3OZrXSw5qP
C2r9HUOfojZgY+0ffdp6f0SUly/aHn8xtP5qYwGWlw2M1axGxuzwjbUPiLTqu+Qo
VdzAkAgky/yy9zB+fSh8/3fHcaPkrNYtGGP6gznCNUpGF8T7nnDXPtBz0tLdNUnG
Suc/F7j+ROf/mBfdfkzieKB/jVMg47YKPMvx8iRFqGnAPTBFQFx7yaosOZQtpsdr
gnbi8gi/9G6QXn0LbMzwfYbNgUrRMhFPw+/41E7PAXDHFYLkYAHPj9B5X9tXkFlb
m1MOK2YpwlMj7Wzm9SlHsvNWPSyonPMenDPmTMBVQ/dTdc0wMnap1bQ9xISM5sUh
q6EjY93ibfWi1LSVPXavrIsTM7hF0Nr9MmC3agh185JfvytrzSlmnJWbBUG0VjdL
PfotFSvRNwy+LsOLCAYHlHk890B1E3CUsfeMdy/R12u9gQODJCpgHtB2R6rdRwq5
efNqkdlCKoETEGyrCeEm4nHBLeGp77LeomGBuM9gYS9mPJ0/iqZloB6LRUJZCqzs
/PwGyeO9rPN9QxJbCM4xEHx+XCFlOqr1q0K0kBV0nhqN6KHzQTlLeSRU1bYUeWhX
fdJ4vhcjMdrQcrunsjbKP0rzrpVYgOr5iiGc8sowteG9voREyijwPx2sm9ySUG9R
j8K2GwAHS0aCs3Vd8OVkKZcLvunIPvJhr6/5il6fjZXQWRHxB4wQ1qZO2gU+aJ+w
TfI+vQJ6m+ABLpuOauGVEWL0kkjdH/5+9rcRSXxS6XqjEdCW6T5I2AKymohuBb19
hFOYuMJfn+vr3HoU0Ma3IrK+oNfm2PX18cY0lD723MZENzIwUpMMYzXCMQL+lzPr
a6I7ecMGFl1YO5deh3qJ0LV1OX1GUIF7GUsDGvRxL+nWLFghIyo0jGB5s0EjOVH2
kCdMxTjvv9UOM+NfK1JImY63RVFpp122YdMfOMaSayZqrrL+gqdIyIfNKmyv20I2
zdhbOf9dFU4Dpf4cCU7KsnvBM8c0e/5YZd59G6dxEoSZ3/GA3gffW3rz+NAkXSUV
XsidzHs3QiRyOBZ+hTREdPwsnQsfyctMT8pCHq3TfCKM0h3h2xZaE75vdb7/I8Uq
4Wql+1saQRbnem1bxgZowLo/Oe3iTKk1VT4qaeHcgBieN5TIWi55Stj8PvRZBkxm
bg9VAuaMhWc9s0Tr8BkaRQ21R4uP73gfBZB3IYvF9DBZUdQk4NsaGOi0gVVpRDiA
NtuCA4Zu+SSDGzBt3Xsei2uBkAfK9CI/YSK5yN1P9yXW3Aatc4mWoGuJ6jJoGOVw
z3QuaOmlV4qqTen8QddzL5sehxpGW3oFxpPiEj9FaWIBa6jWzQcU614uAxGhrs/a
ariVgSTRTDxrQ4MHG3NaYQ95ApcWHPAPy3idmzmtqOawJ7LOtD8YoRXpc58ECpGM
I36wgsazMA+/4DX5LRBhFp0MJZwTpA8ID/T2KOm34iyj6h98PkfR9ebKQXtzviQG
uX+P4oIA8T9A3O5RwdgHrCixpIQUoZiQKdWUOPVUI3ZNkkt7Zr8/S5Pnbozo22+Z
P12jZk4O0NYm7NACuipED22/nsJeHcAOnqUdqRL8TKSZA7GZLrgzHP0eEw8Rja+M
4pOtlniHz8ytSdVELiw1TQx2V7FFbggoepDOUcpz9yJxVtjGQajEt5XQTTodTAYw
Les04lZMJUMiMVOkDwN/myOgBtENpmlZUr0C7Nbm1Fel4zyGTf/aWMwZG5EquiK3
C/8MdUlLHLzq+UURULjaqG0qTqfAs3b5JreFKX6XTWWJV5ULLi0piSdKrs1L7b1a
X9njqKLK8QqCYupr6FBNP6bmDGPQIrIsEfVtwyzg9WwqdgQ6HItBP49JAkQTf4za
ChGpvXIh+K/0SdyGQJh85iZvDtPOyGHN7PfeU84LLUSq7qsh+8y4AsXIOuoRGDhD
QADleUquqssZehwGJ4b2RHUhmT3YJwtnyyoDAHyBJCePiTwfov0y8g9AdyipvW9r
/jisop4QPiy4UOSoiZakuIthNw5nZYMi9SM3jmLE+tqjASawRNQXZB1ods5JJUHm
`protect END_PROTECTED
