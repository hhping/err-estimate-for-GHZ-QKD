`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzE+7oOnWGjZI/PrpGlpC7nsy4J+MDcRqaM0cTPlKe4c2cVEkQtbaRDmjBDLTjVT
Upu4cplVUqXVTwOWf2aaiYnH561okGeQlmYjsb5XYtS9SsNc7dhG25dYYjYsek25
4eZt8/+tMFuQ6l52sO+yr6uIvJrV7anWmRoCQeufMPAFap/WL901+RQQPntWi1lZ
4jREz43JE52XvDAU8YN3iJWGI4szHkO9+Ie/S/8KDdtIYIOxbcXmlC7vIvnHLsC/
WSZll5HKNJ6Nch28YlVzB4rDPtNxA9Y0mD1THMDNZmodP/MW8tduqoew8xz1DC0j
R4fj4u5t/3tr6ptvQ2DxgtstUKkwtKYenJTrWyR7HoDLutMUZhSAUwq/lu8UuBBb
tn5h00YHjent3nLw/8YD3v/MUvarvfhEla0xqaibaDl12k2ng1ZqgOP2YHTsC5wQ
l8p/vrcCbSGbC46pbEO2JxpB4riIKl4x2wDccj0am9UR+ekjqqQ0cmPLAZfBSUsF
IyM8SRWCaE7P8PN0KOVO5g6DfVIgC+YNvk8vuRVjC4H/l6VfUVHpw23OPh+Suk9S
9wViPDYSRwgsvTUVQJ4IGS5XGRRngz8PCyTgR1pgnWZyF+oPEA7aUg+//WGB/v3w
fgT12dtyF/62xRLg0DJu4aSvp4W1ssy1cK+Hu4tlutYCZDoWKjNwoeVLZG1rhiDe
3dVLfSxhPhcU15Am+rGXbquR0lBFpXNVofAi+SEVMiQ=
`protect END_PROTECTED
