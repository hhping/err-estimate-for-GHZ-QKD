`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
upiy+5qO10VdgbGFCC1WMcNQh+xcEDX+E1kOJ1/+3+tkk2CFPxrthVjq6A9DmMXy
O11tIPeTTQMIUpiOcVndlQkCfvxTP3mOhsAxXOehZHG7z5yJEO92I3LkPXUKyHxt
ylu9HT+xlVyZ6ijgxc98KhgaP0UCZqSaN559Sc29y856VFUbugcS/wrBaXmpzrPR
K5TpUKzQQ1QcdhxImrLGU39GI2FXsSsXxYATxneNDdtDBprDsKANW7TLC/OPVOe+
qz+QNUlzvtZcGBwaC5tmNcAmvj2eZ98w5o5DoRZkKqIHE9UnhpIbl9HfD9L3K4Td
nTioyzWWjFrekevvVIJ33R+WIAxqX+Sfr6mQtbSJlZEru9knVHqnL7PV1Ilb8li8
oBD2Xm2UZVukRVfAx9JoukHaQ2GyflAkBQNVH2ynbrkkN90E80aOQvM9QC4saGPs
UME6VWPcTXhZcSgnNVs9UeBYWivUX+P9Csuhinj/NLtnxYqpy/ZiEI9TMyD7FRBf
CNe2HFOZJYbWQzz42SrDtQJPXj2KPjDw2abgTL4Un4D5Pnj606Qo8RNA+xzIRecP
7sUPBis6fAr7lpARxXomsGmaY2Qozx6NEZpJFD+e9EMWBFjPYM3lmuWh14ivs0tg
TZJpkIifqgUvkQPOgQ9L/x16yMEEnR23feGS8AHgaY3zj3EAP7KYcuExx5e+NNPk
08qWA72rSufYM3gUNohXPUkvYBZqcX+sAQQExkLwE/Fps/96FC2EWPy3F5GzM+sj
XOTXenvtM2akojeVCe5WQc8nIzWdcvQ+ilU2XyMyRca/JEy9qoJdmwvoPQUqB6Ad
8mRGcdsh1+iMfU25/YHKEYFkvLregqZ+sf+ElxntGKA9VuSEnmp1J3iEpXBIRG+T
dSOAUFeKGlOyYTHsKOTFckFFX06b8arlhTB8O1k0Xo7BZsn677DnmcOqhPdxo64r
je6HvJJfA5qXcv1zgCcoFgI1pE4Fz6Ju1NSYlRLOtbauzws6Qvip/yiFa2shaaDM
pr97irpmou9kb0tHNDehcqwZxgz7AkyURyMyFZcEWfIMJnu0BdJMPry//LLEJS27
mgU0A3hzwcJgtDxzli463/bw/N4kecDU8eVn4Rt/cXxc0dpnkx7745HzgrdtMvD/
3vSH8bKd8tTa0QBpIx1FReZxuhYKKwWTdUhPcqSuTfYTZrjDKdHKNZHrp4giPHmd
7s+cA6ET5LS4TSahqK+omZ+hVMPMgrt/xMnMd6YYPotCHhN1s6dUsoeQ0/+mrMep
RVfI8Jtos1meIv3EuTN7oVuXQ0CkKHN45VjxJqO6i7Bk5wCMy3+TDB41t/myQcZ9
B4fO8qJn+ZNAx7MYFKFbdQ==
`protect END_PROTECTED
