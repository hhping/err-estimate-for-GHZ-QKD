`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYiV6k5vEFRT6CkHMA/zIdZt0aA0+HV9wrx7i31fUCHYp5djBbOo4P7DDyBLLI7I
KyM6Cw51ZlJbO1PDoAyGzCIsgbImo3mW8OtXb2or89aEEcKFYyBwMUQJuX4+1al+
v7ZR5M93KXgelQkue7MQNgrnSKJ8TK1LbFpBu1weOPazTG+xVBGRIVgHEfGJ0EW5
MgN8Xgs4+izYgyyHz7+/1ny4xHHiK2pLpxpgOaVHwoY1uilrVbUaMRgmcfDBIHyR
cfmdMs5Y6cyfx8Yd1wLQBXqRwUqtOBDoYem84QuMBzbfxJp4r3PglcC2TcGlT0B7
eJ8O0jFCqqo5stjWnBpR+121bjnYvlM5lZF64jRLSgvxJyjuISL6w/9oHIuGtVil
qqJYe4nPRxroHO7ln2iwBZXdXsf96P16Alx2LrA+Q+KoHHE5+SqKZd7fiTDz9qXi
QgY+YKyYktEZRLUGOMTku5yWvpUH/DNfhwvz8Mxph6pUSNFqpzES9Yzr7DmIcz6A
tyMu863zDtM4NDOUUiCbQmBKPzIE0B5LYl0goGbRBuAMlN89BjscSpuhUaTcpM3C
/IaqapuOnlRNHYHauFrXrbvm14NGoCahEpYSsaV1vZEVfPS+W8tBH5Dpyp5REZ4n
VAtnJ8nFggVZavi1FlBN1Cm+rq9GarkCXUxqfbN19gVpwJ1GHzadg3q93I93TtTQ
fa+8+2DV6NiF7W0SNux5yufmxcOhouD9FNsQW122DGxhwczNCsqUvMjkNHC6hqzC
tjfs1yb58fb0itJ+GXD9yQ7/jYr09iv9uAuxL/YMWgBo5WCOE9XyBjP31pa+AidD
IoSaREIZ81G81lul7DiVH0jOQd3ysGyy04+WbXr8M8vADedOuOdASxehWQPx5+ln
pgPeAKoDbCu0lffV7eHw9bW3X1AWC01qA/F8pGnOmmdkt2Ei3coGWBnjUuru2PeF
/amPUh5UM27zWPSvGF3k6PI9Nt5hBe5aF10QnbyG3OjKq2QDEFXBU4Tw66XnKz2Y
wgyynVqDOE9TYmoiEOnn9rq9ej+O11X+E1V6ArOXtaYyd8bvbuIhQ9kmgpFbIy9i
r0qI2U9flewox4xM4JhJjP8kBs7LJybYEOleDRNrQjyXNCD4ZOHWi5e3+5AtGaMd
NSyuaPtUU8dBgFiYjvTBjY8rxGoyJkCfkhBp+v8OVqgdzKQA/tVgOq216z2WwbV+
Q2vFAHc8vdQ5rPgUYd1/OJq6uo9yLbttZPFZNTTdvCwAuzOaaqdwkT60aet3WwpF
GI7C+NZiwKAi1JrkbigbL0tuH/KNTqjE9YVaEfgBHDHC9eUJDF+ewVycFdkY5hiK
Q34b2u/bUdUNZPDsNjDOiAjanLgQQY8HjHuGSO0SxCMb6O1zILZHjBrP5KCZ4qcC
BkM+0UYmLahDt9Yo2LmMBVVXnXm9vlmmjG1pum3mdwzrDpE4tZPQM/IgoAWCLJ7L
ykvJEc6BOMbV77EBIGWP82R31MOEw3e8qVCfkwlAAKc88qhbkehjL+PpT+Z5aeuY
mmZxOM7OEIbCXjngxP4c/qci/dY4O5keU8O1mq630c6M8x7pArKb2LAAeXq0nYq6
euSowmurDCz81LIv43Zi0k5dZGW74Sl8f3pinxEmkkbzoF88YghAv1BQWY3o0HBq
LmMNpa/3RjmdvYiawZ16/+PSG5pbFqByIJOoLGfeywc80AvLi9DNvOeyeUrCgNCG
eBR6s1d3jnsMri1G0LJ5pG++whDKp+7Gafm+FtdIhNNql9b0jx3q6k/m1C4tkZfF
wcfofMU4qJxg7z9x/Q/5dj2jIdC0bHLd1FU/zFgWXaGeI6e6grspdCQqiQYhMMIH
Ze26kGjzFG0qthD7xeMB2hsD7vh3VDkwNHRdNO4/VCxG91VG3DNW1m8Smo2G//lt
LNu17veR+7+0Taag4HBlA5PoVUxOQtI/fASXyNhIhSA2ty2qcf6XWkSsA6QVLSrm
d4ESxMcwalVxZhHzMoR8hrgm0I+IqBEqCsEYiT7rzmqclr7/UYVrCLrR3eRZd387
1Qq+wFjSzaIYFRgLa1l+rNxKPtQTw6eEN4UexLL8E+4TC9lWIqOo2hAiIXNdwP3l
f3MKnh0q66JUNZWK70SL3lIrgn61e6Mg9rSjek9FlZLtKk38GCmOBtqACFcelDSx
L/gWDTyODMeSEF9S3mFQBYVsRUkMVTPiIlVHBuhsYgPXhxd4xU9xbaBzcMqukZGx
hztAML8hiKFP7te5odHgZ0Hhzq8yglmHsL8OWCB0CWKm/UozXQ5X9w2JJ2rMBlmy
Vx90zKOjPn40azWSAQTm28D7floNZtRzps5TJ3PfdtbBQ1l/llxnqGnhY7OsYX3T
9yf8HlqJyYngzVu/h/+3YNoe3daX/OYIrIzl/bbw7uL2lrw+b3HFWyrYzb63JznU
vVoSQEJpATDcmd91rh6sMVp7iCl3hrADQ68luuYHpyMp+iZr9SjbMev4jwEJqn3a
aQqi41YVMA83yyUZrKvWkuvGfFLlwB6mObGXeQBW/RTyPp8L6rK//iB5XzaWUsW0
CS+ZAGABwvsbjSqNCBa3CiksiMuhB7oDRHR0vx/AnR3jnxOi2yOg8Yuv4XD/goTN
kq85icKWdma/tL8lA6tZzRxK4bCeIKX6KzCEGmFITqsvZnlLSh4+ZLut9X84jAtt
I1w3oNfxT2iotTrwKAzSDbltMRRZS0wzWY2v7KNhxZzd0a8+fign1/6hZtjChabd
kGc1s8EKMYTdHBJ02HqHLvojkHKrtCQtWlWSFno985E7UyvPSut3MKbz1pNsOdIB
rkMhSRgFYBC9Y+FBc+/hbubo6rCcat6il5uR3Nx1qry5poAd07yM0JXlNbP2gX5Q
o7PcSXPeXgQ5pHVBITskQsHHQ99uQHyQ6MGbhAWNLMyUkqj/ca3Xx2IALGhUqNVI
MNX+wQkhx3F/aZa31aX78GbARDWu5jl+D4VyIhD+/5vCLE4+TPp5Bxh1pMp3pYSZ
AvjD4LrJ0N0Ta0o/yW/zWeQebmFn3D7FST2EISrZJ6MTKkVgAZE6Idnwn9KomAif
HsmWt3R6e/GewBzOFZSKl7RZp8aarvTt9bpGA85I0acYNhEDqTRlDFRnMRTejQ3b
Q/KlUjwjSm1QnGWW4gWM2xl2Ju3mWqk2RklYKC0k7D5l6lzgSTn4WCmZEMQkRAI8
wUoaikc9i7GSMngPihamHYTQmSps8SwkqUUBt0GR/YO5ymqPMcONdTL1e4xJ9hfQ
`protect END_PROTECTED
