`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4IMKCNYst1mMIPStcXuk3mPU/xIi79UDwUOoAnp+KxX4XLwOwUSj8UxEH1NQaAHA
cuNx5mkIK5A/TisK5d/QYqLz7viPYz+aX6ohogBc36bqwlF6XDe58b3v5iNzyoov
eSqmYGIhq7N24mHFglDhhLipIfWfr1Pk+lgRIa1fS/OTKrb2zF6mwH6N5ycxpYI7
t9ePLjeWIuRAXMIOpIbOW2CTySWb8CzRcYQ55DVd9cjn1zMsFZJdTrNWw/K6zZZ5
ufrmD9UE+f8WqIighZV8+tlbmii4IRvjdRGRfE5pkJNQP9/nGbjrfm8OwHuSfkCv
uWIIWO4A/GRhEjpcq0p6Q5itYJqEowonkOFhVrpcMEzyz+Jq2HmWOzjroevQxCbF
dmxlE654S371CV1jZ8kWQzlynUy97+5YJBOrWnBjki04ZwTUfiENq493FUo1dpbn
00Cz4Kc3tm09OqDX/s8UIKIcUU9Uu9u3MeeHKIpVE9PK1bkY7ySh9GWG3bUCq3FI
oWxXj58FG0MCYU+1Ve/z7WWSKHqkREb/YBFYIGgrs1106kkWW/qR16zRJ9pWcHqy
k3UbkvCzxK8XCqws5mrXGPOdWLZLaePLi5eTs9pvDZE=
`protect END_PROTECTED
