`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gw0YvO7V4JwgPoHJximoOS/IG2Gi3fMaeF3slu88gucAnH8MsrKWKHWLaBch/7Xk
RPfgXhCBdC9KjQ9+aMfD0Z0rKA/ZC6BuYajTRH2y3dfFwjOiTZKn5fx0ueTHI+05
73j0fN3sqGuHP1YCBfvsr8dS8lXt4ToelXoEpcuuZnRpqdXBTOu3vSvA5rlOyicr
LXTM8NSzc+ifRFWriO5OnJJ6GO5JCMCjxOJAT3s1piVEynpyWY10OJf9edei4ZV1
j/OoUAkJ7eO9R0Hih2me9T9TtVrqe/qyH8VWF3rtqjP8kTcQh6JK1s79fXLYRlkd
hVVwLpr5KAC+fTOpcwL0otsuoYXJnJ4w8/RdcY6FY/Kc9Jr5TMjlyQft5ap+mLq7
n3cig3GhZEebNc1DfICDSlpaEg9eOxXE+28HFYAf3vScplaVnFeCYiQQkgyqcfA0
dGdQ1AmBJ3YZFMTe3lGA0XoWqEgALBzelG/j5loKD6LQqqoporyjcASCZMp3y+Rt
8R+Y7VdRzCmOGnwZD5oW7eNV5UrAMHL140MMMVwlTmdHXVMy9sSSJMiPFCEkIzse
Jb8ZJ5luR1FSh/cDzyUf89EtljHi/Fk4mf55H3Wc3WRrvFhvOhEd7wKlb9EfIQvG
BI+UYebfTI9w81jsMSpdizUW7yuKzvX9ga5wNA/d9aL04vFko41DWXXWoUoQI3hf
kFHJ3HJeh1/0yoBVY5WpxdWnz15EBJsHw+ioc3omfKxO037t23l7f3FzLvkCFldv
uNuBbMckhalkz7v52BWK+uiEWva4JAfgl+sH575b/31fWYU36Trv2hZTqD6dlPdd
VoHvMRyVkWhkSvZbbK+jqINyLyiX0RmUhhsgar1wOwf3pXNqVl0qQFZmEKBGtdSN
W22FgRrZV2ddPxdJoJpJGkGl3SEZqDgP4MYebbikofJ1v+HI8znC5WfgBFS2M/It
exFmG6mrW/Pag+F4gzWuZS02s+h5wuJg44JuJi8W1VcRR5ZaesHesqsv/udcp834
L6N52qfLLI99DWhLAjOEvERbF7aya6gRceERSfi6srsvu/bXH1sJmCHwXvCI7EX+
PwOLLq6FE5qX5Cd7KfzYXN9HDywi4CaNxO8O2rYvCXOipyR5ZuLVZigK8+2HqmhP
0vlS7DLkI9MnEjOjAvLPL6HLvkMHFsEPdSV96evrROm7WMRXtTTEEC7Uj+bHmbgH
+jK5ZWijGQP5XZtlLaWF0QSWa4qbxg2kUBv4aIAsM6QsSP1jCkxJ+WNFg4LQ2rmz
7c/ASNvJVAbnnQi7t5jdUMveFYBn4c2TvB0UeZiwN5pUl6SzSoJWrsYG5CluiQ7b
`protect END_PROTECTED
