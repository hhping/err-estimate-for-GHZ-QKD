`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMWpdVphI5J2uXZodDPyHhVgqwMVIGFhafaSjPnh7lFLa53Sqk5jvr6U29fFjT2x
2XA4yaWGopKP01K0hvDN2XOkiL3ncPSF1t/OL0LpKNieSIIv2pI6jvLuynCVMt2C
HUgeozi76hqZQI8mJytebUQ4FtfveRy2saw8ytz4gdKfisXeMh/Q/0Otdko1mjpU
G/wqeXWH5lu16GjovUVEEQqZeIlrPKC9T7rugMAsbBiox+/dmWFJI4LP0FDRFU2J
D08plkPpEK71j/0Xc+8Ne7R5BalgxY2rfV9WMS+ihu3tdHSVVGMxvfhq/AO1N8wj
xT3UQAb0CgriZoUHtCBRHrwdnaFaItrXnfQhnHXryafOpANd4X8YSelJaikbejzL
ydKWlEqD8KHSgzI1kNUGjanpCoFqIkaqbo/IHok1RntpwqJVU6dOhglgaxv0dSIP
1Il6rf6ClMyxW7EqhO4dsvI8aD9MDL1AkGWCJ8kXJQ/R1JdqKSZQVNP9+LC8nu71
6a9AM5PpIDBbngPvW5q9zBQfQhU0bJdPyh4wClidkumNmfz940+wSvRgnOxQCDD9
z8SkOSRmizNz4jxHrOSw3PtumwK4QmopgHHAtjknq6ZJMAEzgYgw8Okwll1Ig5Y3
b1/6FNGlwgL99T/jrzaIdB4raUgUHSFvLPkjYTNadLzw1r4CbjQxyQIxbYSMSH6H
e6bWwS0+1Ly2EIsEyA+HaG8SlK8sQ1qrtdGfHECRu2EYWWpuehtWmbw1Q24pLucP
crAMq8MVyIhvPn464xzcKR4ec6M9rGJHfdiZuemKmUWZAtF2AG8L5JMFKpZZE7wY
/FamODBiSokKprXxoSujhOjUymxocxgkAeZeK7O7W7TVADVDe8w2W2k9FqORxTub
cITB2z7s89KU1bbOmEi/axdUUhfJYA5E/IkOPSfAlA24xfSyoSpyKaWoDIgvpaQD
kdZjqcta0WKTeRj12iRNQ89YJiD8YuqW6bzqcAmd3jLjepSnbZtge78M8QU5KXyF
KJRLZiB220sKWnrJm7yygasdzzAypLb2Z3l+4MX0nrcoqSY8lqvFORt4nkDBdWY+
+YGk3b4NwLLOS2M5uTjAJGPLQKqQAGSyePIgKmRFJiqWaDnTtAWBlPduDWaKuHXf
RdTlXfBKQy0OtSamh+Xc5E5q4XkLqi/fgilYa/ruhcdJ0Hs2ZcKeNHsy8+num/vI
NqrDhoQMBzAKNFn9KY7htiizoTVtSLfuXniK/TorDD5gTIikiCkp8ptQC4QK7C2q
cez9Z+Xl9SyPculCuyelkFrwNHLcUrpjQ1Huje94aczsPd3uTPOs5JtydWv81tf5
g2L7SWXQXnjpVILa7ZjfM7Gczog7CJlAxtv4PtiNISPhjbSYboLuVPOUmGIf3rTc
`protect END_PROTECTED
