`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k/kwd6Lakcf7bRHYfdT59bhludvxmyL7smDGPBAfjW3+lBdP9Z5YcG6DdUgbTTYt
AckKA1hHv7kSVm0qaxax66cMACODJXgeeJprOK8ip8ia2qcBojyRHw5PG8oqH77e
FkyNyPJWgenLtWVK1Y+2JEHuFe2x5L2LGxYOKZHXWeNineoZ8cQ0+88K3gl55qUI
ivXknQeq0rK1uWtEAtDAeD0uvGemHOSXWecsAciZe7lriW2kYxoGt29wefYe2gHa
ZxMJSMldTtJHO1qIs6kGYK75OoG3b869aEi3nKEdDutGzKUAYhpessMy1jvEnH7x
Mq24o6P2UBM070oJQnlPqOa+b/99jV+NY0QLUPrL+TWvw2azaKFKO+17Mfym3nWC
Nqs0PUDlXoQsmHxPMJuAIkLZn28wUJ6GpN/cUl4AZUgCNKCWmMm27s/rlLKvzT8n
cHVWKB/cSYIYBAkVMKXfUrrBWjbO15Ea8BbNdq91J8+QJuFTILQU5lvRXyrDeDdo
ufSRxcs++7g84oluV8Zy3nn3UG4jdyNvjgL9konQ4std67BTROd81LdpmRzf4dwm
X/1NqMlVcxB/2UfzLFjdf7H98jVbueSTBwSghwjLULTmVTuT3L6gKdGNK9PYYyGO
1pLVybfFnOsV0tL+wtbWfvTwixeCu07W7+EFzkUdyvWtVrGrVO225uid03mcbKPT
QrZehy51WXRyPJ0oC7j6a2cNLVu/1umSXotDppJEY8JDNFsm+QedI//MZ2Fl5mmb
+V7t5KXPRv//zL/ZO8cHd/js6Z2Hp5zzWMB0Qn9QEra5zHRVevEMztmZFysbdbrh
jk3ggTTFJ9vhFFc9kG2KMOiDkkC0kM+1JjVWvsGla5cSWLMiL6qM+nrl6hcxYmgw
tFld1pON3QC9EsmUNipkBqP+ZkgEP6yxeQX8ZaYokeK+PL/PHT87Y/PsFnkqCKfL
q0cxdeuFgdo/WIEuvamTD5EJsZaz5qg8TNYXGOEMf3bW9sKR+1baswzZ+0ar5uqr
N66hTGl016D1RKzswS13Dx95k25GxwE74gTSjj/+547nRc6vXpJL79bMBPIOx7SS
sigDkrWfvavtKNxdrjqYOYU32mmXXb3xPk0tBnUiwgkjtre+nsC36OsHxaDaGa4A
`protect END_PROTECTED
