`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQ+QC3RP9jaW4BGmkU78mq6cjtumcs/1FnRGtUbibAwmEn2UTHEL+HdAooUPaqqc
B+bOsU/TG2dA8C8T7QhNLKyaMsApDCyb5bSO3CHJTATE9dEoW/nzAyRFKlh2+k0a
e/fUkJojKM5rlAQ7lTSTwSKwCv6/pkBJEAoRL4MEiygH64V8DaCUXPyuGdl00mss
B8qLQVCL6l5SMGNJLQCKtMZKL20th/JLMGaGvuTFG/8tUwitUDo/blW5Ja6qktX+
/wxpXqNlRf2PhuaW//05gHvu2FbhN+jAQIaZaHZh4yF53m9MHLKfu5NfyJayyemz
ECrMI7zanxH6rszEE9BHCVNzP7mH79s4PKdf9Uftd+v4MD9tzNpC42OaB23DAu+O
HhkW33RHRmxiPGf6hAlEp2qU8v/iXtm3vveZ4tUdpYcPzbR3lnvoLcPbOMf/LpfJ
YgHV8+XHigI0ZpJha30k+NDdDvTWdv/qtPj6ZKHDCPoiD2n2EqpzKHUwD7S4valf
Ed22IQGxO9A9ckQye4kpQ/UWANLAnUs+f3u57OFD5jb83POv175H9lVBz7lDq4Ug
NL1fbKNRuSj8/SDZ6VEearsjWiKj+/d9aOP67spP2lVjpHLd4/GSaZ9BQDvWYTlb
StdEX2RVK+jb3kgrsdP2zzts2jiGx5scqUy5/UpLrOhyiLaU/vIqKQAfpllnwfp5
BcDdIufOEsB9jBhIuwW8QzkzD8SINOZ8TyNcERcUzscaVNZ6xgydkS2ZBiSotRFs
xbV/05O4bUFyjuGxHbYei3XpNptsbSKyMK2rBvMAaUwKzt9u8aFd5DurCy42MIW8
XbTm3Dac45BqF2wzoMPIxcU9vEtfbaDTMRAaT4CtdghmHZ4aBnhofY2HPy/mUOJL
vA/LxsDmhnazFF9GwVZTnBpnCtjL/tuutLpppghc+BluB4GdwkMb6MqqRXh1T0Oz
fx3CJldizAf4zovE6bg3qQzasPXU64tkDkXe1nmCwqgrvxThCAXhmnIq/48WHpse
4WNf887v7WsQ2BFKNEs7za23UUUyx+6XTIzTBnRn2aaGhCpHPX/teVAbTCd+B1gc
2Iv0KY2nd1L4OikMwsNHzoqR/GV0OnGgBclm+VbdyWP0xfi7z1wHlMWFmNPQk5HL
0LYqdwNfY+wDelmHxHDoSHlkIa3yQU3hvV1Sji+IH9FfhOYQT5kh/nfbtJbXQ4qM
yz8LkKJawmHcxIZet91EeO9h3VDNxM+axAlhVd5Qo0mmDJYBSWVNmrKftGjqk4aj
EnTYkHQ7WG2aDvYe62dheSBq/7P4myaAV1wJxhu9dFxlwL8M0gsf051fTo08UYOY
uYc/bIKLt3wD3nADOGkv+xjZYNdBnWLBZh5tUYcSX+7sEYEr4poakPotQDKkX1Ie
saswXXjgr5j2Cd5uxheV4JzdWZI/CZwdGBvGY0OlO+BVCEQegw+da9Ibs2ncveO8
BaIrd1itAwGpRff+fof/Oku3tKRrTUGz8ZcqiYz9QtppHMr9XKbRGwpi31ynVzDd
kRmuk4mHb3HyI+8645/tqNDVhzFgRHLBGXkEpQ+rQ8FB5MKjlZAicYR6ZkwcLcmR
Nj72qo+OiVdGSyJkYOgK4MPx6WjO4QgBkU9JCXiByQKIPe92thxY5LtepjHsvNBF
uSNTL+8nP/zuD7+cjkt2dD5BxIpjZjD5tvM/+Jls+YBBCmfoYVJpryfi+kUjAXWd
nfrz1Upq39pFp12kn/5nAQ==
`protect END_PROTECTED
