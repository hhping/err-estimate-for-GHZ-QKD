`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97uRGslyy3Hbl/e38YLOv+xZJ85rV8RygE4Mo2hENQzMMAbCm/urSknjvtDsf3XZ
G1iXmec4xPZ2yXbq3YZpjiDHdy5W77eRG4qPTWvOG2QazZNA+mbuTaAKhHAcAs15
sg7QLCoxojxjJ6lGWuI6MVZEgj09o8YMZCKdYYCI9zg844+YgF+gC7o6via3QsPc
NagqIwHHePjo5kg/PApnmf7/3F7H0wU2ndVZDfvjAfX8oPE5aco/S5qvx4Qd4fI2
GhzxXVTaS4j2+1GNWQyT2ZYaH2/zEW8Y3p8ShT8FTWDM9ynrkPXimLn+MKLtnAZL
M3jXzpZ0sTmQdnmhaSvEdGKD0yUUgxwmyM59/AS2EVH2ciUHdSBz3H3VQWyR3g6X
v5Lm587i7fjrgwG93cxnwykHm8uwsTWFeiNUMduXQ8MKvyMLisCemPBUJBrgEx3L
SfMvYKvDdNJhJh0TYqTmT4ADOo6bDyP0FEpuL8hO3JxhL6Fra/kz4P3hVEh3Gh4N
Bz6fyt3DvP/ji12ZTvt5PfJOw9DftVFf5PU3ZBfQO2u6Bf1qJwCSSx7TZelTpux5
wGirr1ktn7MyBYIZXnKCD1RZuoKudcAFbIexWZkL9sTjZLiFk9Gqa4YuCMdZ2tHG
dtqxbk0iXUpMSdNiICoyZQrl3tlVztSTxRdx1lMhawAKQ0AnHWW2PR2FcPTjalMV
uw1MsB28aNpdm84qC/Howtsb13W2iAgHiWvzGnwN+5OAZsuUrVz/JKi5VH+SqYYg
P0mVfzW6IJOkoaOQ6ALwM+EjM2yyYQKaW3oDtPrnKxVQunRBRi99B9RhDqz45a6G
bTVElfNRzpfGFjK9C+PsdKu2Ee9tD2PrGpZrHlFlhvkGSuZjKEU0XVcvmii3mfJx
t8hYpNhNMBV3dEuLJqunE/Qqh2aLnxCmZesCaXDn5UV8V1Mcv2pCMQi/aTa8yqb8
`protect END_PROTECTED
