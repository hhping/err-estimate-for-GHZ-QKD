`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwRELIU8pMkYv+3RyQIle6NvVdBtXoD6LOcikedFjDSo+CPd1JZUrX52NGYuvYVU
q35bG5fQ0c6zTa71AlOdkkD3tYCVXnpfjWnAfgwZevKkiNTj0twd+g7OX8NqczkW
SqWqMNn8HviEMZy5RssgyW8mubYeTvyykwhHmTn+AXZ3EjfR8QVXCQnEAP65AKnI
xF9kaSjn5KT6rXvCGu+xwkeE4URQyA7SW+CZdyJc98C/PEZbxGSi3qYI4llZwNyR
LXNjuus3WdSSKD6PX0WK9Uj2doM+1jS/1dEbdk9evgXp3+ZsMsZAKwauB1jWi2tL
FuAv5eX6dWleJp0jcpWesSh2KY8xheCMoBHkURT8BdppQewaKIuxbf6Wi4vUgDLa
+hS/nPQ4hwCxdbiUZ7xC6kobhkZvvQjQTSzXR8ybrY5f0I3MqmevKFDILBR8nAkj
MOI+/WT7AIsg1xlqv2tixFJvYs8mhW7GxLW4empCNJXEdYwwq35sgwlhQZe9pvIF
c3KmfEjHR/aq6QXo/OZcugf2fqKs6zExvUSJDA1GNMtH8GBk5ky/RudKt/JGwNUo
`protect END_PROTECTED
