`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTetED7LwpEXFfF9X/8TguSHojQpqlJepv7RM2HHl5tCKmTiK0+2gW7CW+ynPskU
k5gxINMnlgi/EF5XSyHayNR4Jx24Sagr/a3/ogOp+1SGzRUAj20keRqw/lBdc4dd
4RPdPs6mLlkvo4JGhNpiedrAov2ZXp9TZbghvHgYOrYXE6tieoqrwR2DlE6uaCEQ
m3mqA49yrJypvuR0JkW3BZj95QtlXDRXy5a1+3Q+2ebGKBd/zC7kqlhzaZt2Ps3w
QpVEui4OP7/AhNKFXlLy+r5L5o05vi8mjbqtcTdKqyNROjHDMxTayXwuXJE0rS1v
5T5+dXuWyROIsHDujLf4O1jW7XTh8C7rdqQMvum0mHMVB6eN+pPE1zobB08BWrdc
z1LzfMhwzPo7b78vJSFe7eHJ9rzFA8QwZgiWQf/pYUsCKzd4NLAXJgwBptFXzjRN
+On67qPEHjVB2nkNP5EhEGeJRC400vJWPiqiEm1WKEPPLSmoXmNTrof5Zy1PZ9Fg
wF17VrsptdfWLQTWIR+SrjcDlVriKwHXGNX0bUydeAXaB+C7dAB0kTkAOsSmZvnS
MkldH+Yelrd+pheOOKd/WptTC8Nco7GZDbkknKnFQ7AU/ji54tCtTfRwjWDi6Zhl
xyNqh3O8MX3Zw/ai0WIw2cozmpAJXP3DqeraAkr/UN2Vv4Pvhwf3wnAeXqYFJ94F
KePX5wOpEY0ioEoCboWQyNAJOOx/WNxvk2XZkWrxu2Dt0JBi8HexpOzd9tKTz/Yz
`protect END_PROTECTED
