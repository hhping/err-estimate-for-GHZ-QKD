`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69zxC/gyv1PB2Hb5maG8+BNzE/B2bAYeKNc0GwNAaPcynUzr8sp69g56pyjiHfW4
KVAY996QOYtvurWHUzBZBprEGXmQPAQRQ437xEVppKVBDPiu1IsNx+DKY1GjiKse
UqIYwD+jWohNetRykMgODeWrxBpRQMTKUCVv6urG6wM7N66rrrwDSYdQ4F2CtH9r
zeYbItEJq/EGJmEr+sVcAdrEcHadZL6LA2ocpsQeVP283RtSshBlMi9jB2p/JogI
cMcj5YWZJZKPY82Ud9ed4Tfo36YOoZkBw7XQH1WBL6GliFbyKcwSjz/F4nx/CKxp
MUpKySrKeJwwPel8GzFu9WJld+kaRl1jPTg3wuUxnWad6sQTEZsDMdWX5A9gGSpv
UUbcicLabOtgWS3slJUHrPv+mT5txuWomee6gclDvPKn+GlVw2na5nGj8HIBT5iF
`protect END_PROTECTED
