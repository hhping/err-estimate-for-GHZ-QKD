`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbZaaV0DfirP7JBzMrO83egZfPNJPdh8jM2vVVyekkTeTA21lo2r7Vfni+Q1XaRq
Pndj0aVloMFkNLSamVdnewOz79IYn2hAmkEAS93qcm2Wx1a8QK6/QiMB/AT9R1Ay
/YsJgu9x/2aXSUdCSuJ5pBvTqeS/MbKhf5bHCISoJ6J/cvbYV4l2iyYU0Sa67PTQ
BH+d/Z1XaHwMxEgdqymNBvpxNRz1L38DnVtSgl861ifRlqCSlAknTmTiiTCz4/ln
7oWkB1pBPWlIgUMMhlihlh8zllWuhcC1E7Ze/Hgi9LGs4qJg/a07J2lxkIiScXHY
S8x2uKffNVa/1W2ZInmtQ4RDXewaczFBBcspFuFgbrHd08GiLET0L9l4vEcTdRsU
kQcEMa6asGC1OMgvDWlNRQpLry/heU1vVATCpHk1mnpb6+C+aV79SZG75mTEdis7
906Y4I/1LL+3zFF0PNWFHwlaOiGhG6LXaB+6oIQD/pU1HTRwiXOqAQWqzhKmoQtB
Vu1GqBk+zurdnhC9aJkwD/kQ/E5LdVUHCUL7VPWmxQ7stj6XtSwc+3MoxMwBe1uZ
EJ+lsHn5Z7IA+AC20PJwg2cY6GsvpCmc/aku2fvSVNh1VsF7phZFMgfw+LRv1V62
57PucEUlgLmOqGRkqYgYEZUVRbN+f3rpUtjDXRAt7CnnkLw9f11g8jph4QqvpE0W
im8jdoLnSfES1oTBIpjyxsSfcrAkCPfD0ZNh+NCYYYZJyF2KiLvbHKt6NA1NiF+8
Dbn+CskbzuKWdAraAjU5FCJ+2sostXiXsczRRHr30P/1OO78L1WBOfo3BKHqRskq
qWOwAtI9VSDJRNMo66wSSceVw91rvxQ0Ljvi1xyY77vfgH1WnpK76eRctFqL5CqT
EXcS986eq3NhTqypgtcHHiPaKknKhL/0/rFx7rHr7bhHz9LehcM6cp+k9DeeWEtc
oXBMQ4kaojSHCb2doNYgK9y/uhhcBfAq7f41IoNT/nzKQFE05RvuBlwRVE8XVeCo
0IC+TpJxi+eAhJVLOjIA0yY1ESWJEhIbHcha+jcQcja+OaCe0vgajY+rDgC9G0O/
CmZcWhDMFEdrdjgQDFaM3rsNNf4R6RGzNxpqEtxvOLBrhzaRfV1L5fSu49x4msUK
AEC5/3aCzydhS5lnMblg/9reWWYn4UsXFUT3B0B5nAKMMgKvMe14D3pevdSreAgX
il9dYZvmfobmUU7RxYQh+Mxs8ac0WQcVNZU+AslXniB6elkmOHRs9mF7rf8zjSMv
lGkTkUoFUxuSBBERQw2nqBdH3VvIKAWLfKomTFWR3FJqCzNfgeDXtTHJZ39KyC/T
r009Ic7DkTcHdPLmsy/iErvhDifP/YZv68n/4A7v5KrnOF0wszhCWWpUjsL8fqbF
9mr+9brMFfdpzuhJChf49hZXhUACmshQCdDnGBTyIQ911+pkr0zOKf9sTJLCUdIm
gBzs/dY+5lGL/jSUgzyF1zyX6BqG0YaB7TWETQ21VwzqSJX7HV/Q+GAt/qJr9GSt
eB+8XczOAZIoF8BOtxrbK5WBToSOL5YKV0iA2ehFKiH/8UtywdFy1oalO5uP31g6
KcGzWZVtnGLyHCVaT0ovzDSexzU7DDpN0dBpCvoXqI4KGn3I67tfAHOXNYfAGYK0
IvJ+PgDDBE7gtlyinyMSo5wPg2G9rbOZfBjP57zmCn+oLo3GH2CDHgy5bWVM0kTp
YvzvJ/EWhRE4hN/B4EvCwJ33A3YTUqZCENclOQsPuRfOaQwoGJVZfDbRO28avaHZ
ZNjxKRFDifXqe2E7BwXaKwzoOiKhy1+Mr6A4cjn0rZa4VcXW/ZGLCsdCZZRjKUu6
DdGNZBbu0Kwm1a0TNRxSrVjAJWyw1p+At0FToY1kBmZy0pvnBebQUNbrqMGHRjla
JNy/8jKim/mcsVQvqu5FStiZypkAYzQCVyw3g2xZuMaO5PdU8UX90Tm+Rwxmv4qr
bYO6+9ox4P47R5zUqd/cegeW0x36lJLBkxINpzIEBoQShKXbM9PD8XAqLahjbjI7
Xr1F6MiuDfYRZ1zUG3TPUhKv2Owy3qoQvj/IhyLMkbdAViB1IMEaayOw+jrNrSUz
6hwy8ni3xT4d4kboAnn4HJ/Ozq4yBHGDdMGgX76txm2iRSp2hn5oKsvhwx8ruumR
KF0m/PBxAqauskFMLp4fCwAxM/HdRroF7XHOQUQqB7z6UlDx9icZvft0VXvgSRce
1odpP7MNGxysWcVgrFg1iI2EJsp5h2lAAdP1xbUf+Q6XrjDKum9SUuHsO3gscNdi
B8t4ryFFdMAW6z6K8CA7Y+wdbJe5i8akyM0hB8zizHc82lYlmzrmcf1wLDSIVWJg
H0LJ0zQJGDP/F+B7D87BoOe8qcyfjmP4jL08WWG/WBM=
`protect END_PROTECTED
