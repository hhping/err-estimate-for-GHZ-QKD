`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vRT70mmBfpYp7SEO/vqeW3NiBkxjbRMgFOx74CvGXdwYKgubk+h4rzmYOO+cipPC
CZOHT81elt6e55usRVxT7534QF+J8mZi6TvoR43na68ztnU/BuX/fRQAcm5g9es9
8qkqz6aBH1j+ma1lZwpvwxt9uIEhJQTIJ9NO35mq5+y6D6l3lFq848BQAMXa+S7X
Yo1hGNghArP1ivjWhbsgMPtGeUAw/brFhsGYf9BbRE83eOnbScYcRK1fAmUXYm3Z
ceM2P7fSk5vgtPEXF4TnvTEj6MKtALIhXvpTMe4auyNkr/a0lTSDsWBiQ+cOAhgI
a7/KtKsg8dsHY+0D/MFxbXRfeqh2Z9Bmi9gQYp9E/jg/CP+SWxjUt6IFK0SjL2w9
hGlD5bf2i4xcgwCAXNLC86pQVFzlrERrkK1DdEgGT3ueQXRHNZV25l5yQeNgHD4/
O7eWaEJpPyr2vBTtzPJDQGzz/c4NRDAyHearySYbUDwqrW493k9nbmJ7qVZmCQuN
x/rEovYgVeBtOGrtgrb30jS7avGPRCj5DgngHnMLVT7pS8fREE0G5ncQXnnP6Z97
LalXJ//LW+DUDdK5metGawW4UZrFfhSANvJQjZKcj39UP7YWRu32dvgqiNAxAVr6
zvVXKmo2UgMxEnJCjoImWg3Hd5NQQQ2Z0qT2kM5B9p9PTuAbNmpiT4uzgYFGoO6e
3tkg/TgjK2ZDzP9y29YwPKGkQ4ZON+SqBE+/HU4RTgwgUHStbCtTPww4Ujcf8CvJ
3NgAd4+P+VqMWQxK2JYAkVQEwonv4PS9rdYQ6YGL4Nhnhv86yIIncJzuYM3rdflI
lajps6Xa+j09owRXKZCll/0N8zGRfEm5YPyzXEJClm/NArivAL2SZlKKoK+sIzzB
I3mmLnGkgXxBx8/2XN5QAug8ZI4ebPC1mHoq+RZ8afhzQo/UknuTEAm3yD8x8kSP
fnaqFaUWuN8mZTxM3sTVmB7aJvNserKXJu/+nWCQHDHhxKOgRHmQP2PeC7ucITPY
c6UP7kE0f3100f3eRYK2pFFaK+RZnARQWuTdD+nZ2E05JTaeJvCIDvxwA2TA9aHR
uP3d6qLg+ZnqQ6QJ3MhjeN9nu8WMmEYtJ+USDF+nZGACFlie3w/Ia1cfXVt+1YZz
5DE+kM9/+IZ453FOzuloVyUKXLTjyLBtSLLFgJwf1QR8j/1yU59lxAUneLVTU4Wj
jHEoBwzQSX74ef3rxko8jugZmIkVL+pmrMruyqW2LPK6urQ6eHeHHjfDMuiXPH3J
MaefHtdL5qXeEyJZ/vetmS4D+OPysDD51yPOJa+149VrBhTAE5np+g0Z6/j/ywP6
W7DB+r7g1I/HmKIAOyPWishOF5GlYnVwUo2nUx3deUrYHcv5TxkD8L/lZWj+DCga
bYm/x/i7awhJl5gzsWdS7nQx2IcjsJ9Bk/PGn392aBv/yIYL2PhHtr3NoW69BMfw
nU3GN2GJJHtpOh4rak3UFxedak+XrpaE3lzv6fcVhiOFSrH0aiI999qwgd3El+F1
wjxVysGuQyJFLXsQLdB87rWJtoyEPP+8lrPYvo6hvyYondFMyCBFJ31vWKMukDB4
sF1iT8Cs8NJYVRu5Z5pxwF93N99knGiGWJkyUX3sl0KfWxDwYsqZRIzoRmcsjn2E
4CjSOocPc+VHCBDCHNipMpQInJHM9YMQltXRgjH22K1uQgwYMlp3Ufr7O6rxWR1P
xlKaA489bVBwMJL7AGV2EPX+mAcqILzWa1jCi9vskniJg32CwdqYjx8IfFHQbN63
MU6TYvEmSDLCtAC8/6TVTXt8x3Ye1NbUznRoWKdr9O2wd2P6vmJeOZcrKkkOU29i
2NKcqFvH0nYgQ0OLOgJJ957IhZHG+v6yARcpc/Tu3Q3gonU43Llr/zRy32yjFC0T
5Krq3LLVlVeTt6CQLh5dT79Sbi0r8VCrs+lxgg0ReAuNDqkAI6kaN6jrBu3Fb7vM
Gb9U9tKABvabgefMFMLD3EIPg8fjAnrVHsiUioIszRZhbcAz0fYul7E40waymg2z
weQv07bL/vl2kHBYGrOY4Rlg1VoWgEA2iXTTUOOUqkTSPlsypqTkC/P9oUaIuP88
qAkkRHRGlNg38dbtByqusHxp0TlGYVy1JOsTAsaFkrpL2b644Wz3AhT2KNZrNIGq
qS9XOiM4J5PzpjR+hifpyMk4tEOliXZKY0snPFQElgi375VVk3ePkpNBlCUH/RoB
kEVYyRFsOednSWLprQRGgRWAoNlaRS7u1Gjo7mfsdqPo06RYIC93ndVtydwBlI2r
7nd9dJNgqxLTtBUl+1TwkXU0u303XxfK4+UH5SFhnPDxUO0bHUUt/qnO9POFZE9r
hyLBT5hr8dKXPGyoASjPxhIQKQsKw4rQcze1qwqYDnlfsIgaIDbL+HZiUSP2y17I
KI4Bh+mSpi8rq9fKMZTCTzpYpLtAVZmosRqzlMGI2yTcK+J3Wz580QFGaaRgVFYI
KH/5jE68/xp8TStLq3x1PGViKzoBVKWepN/ykCtNYBhMDdWrbpV8eukr4l/HyxS3
+vRHAegOKyQi8v+NbSYKDqC5e967fUBOGq1Vt8krWDGfcgnHvUn2ShqNCl/1MsfB
H4DaAJAak17n+dksRkrbiODt06OLK9q51coJ0gJkijc1Z0Ufu5MaWW/dfERxg83Z
VY2T0chYm+Ac8iaWU4uXVNyIc0DL/JMPPFRInhScokcNnsSKgak/7Jj2OCJ3v4S8
ZvJozWEMwHiw18EvJEZ7wV7ai753hGQNmqsJ+ioHgXBM/Gg4BoJx8Uj0sEXHJUEg
vXFfLdVTzjXe/4A6mvyitHooCRnfvBJsF/n5KAzSqgnHVMyMIvx+G0kvO4D1vAOv
922J7yxbVXLC3okzYNziO6HV71YxFO2nwCkPGI8Irybah4lxD9fFvi8V3ZFUVYb/
gNBxQ5ed3ichuD8xjZxX4kxI96eO0m3tgtoPEYuH2Xvt0S4yVhIONmJUa4rtE3uD
BWPxgPYUZNiHtgDODlrO+10rZO/qnT3Rj+1cECbHoEjH0/0b33vnnra+DK2Of53d
OZ6HPDCx2YcwYhlMQtxl7Y8e1x1civbbjkgjRI+4Al8kxQn0ubQG/d9By4SUpoJB
2+dkK2OX+Q+Pk52+a6TRyxbxR98DgMV9Mv3hgsZZcKr465xBDIwSIerEmZeV375I
x7DwWNrRZu/EdA357riQb7ajI02mY2Ulos/aOSURS8Um+B1U25r01/wEFLtM6Q/h
2RSSE3bEcZAA/o0wsVnYw3X5lNoBf3BsPen7zSaSz4HFnoQBXknPn71alyhrrWPC
SdhgPhHB5YAo3NvTRyktaKBUDXvsWFa+OoXUVDkvMStXPGtijKoSiM+yUdKQyv1J
fS059LYW9FYcb/4fKqZq7ZeWFME4uhUCRUdxg2ybjWZmqSQZrUNqWE6q2VRnYZTl
qT7jKuMpl+lOknZgAIc0OhghOz7vr6dGcueHpm3p6GAcfrNe/+/eh3g50lktfoLK
rlWAlUxZk9GOM1HEdtUoJAFzzUcNJiCA/B5OuZ5hERoDpdardzoUCTp4ghu83plh
bVkWkd0ShHQsDaXUkf55X4fmrDvIfQEI5rlXrr5sJgnq5+hIzhFBPbE/Ret0n4pb
JrgfM5jP/I95K4pKrgTVkRP1BXFcepIdArkp77KryxNsk11tA6zSq8gBUR+WcjZY
+AszWtaorwpNf6JE5LFDenQARgLgylyX2dsj9A2E7Ee4HltJsKQqeGLRNBa5VCq5
dMv1TyuLLzab9VXqXK79lqgaZZqcw/BRu0EeOlIJ5xNmjuDKDRQ3Gt5+nESsX+CQ
uBt/4VmAD1Mu44sN29YG3jX0cOchVNmMTWpyyNUKDIOoovI7UlBVzvfLkw6pkpwn
LcyOludr8GxirmqpI2j9iLMplwRzxFGrdzEPUb6xSRyctHcsblNw4IJNp+6YRQ3I
oTkwXHBRx4nA1/l49FAXz9KiR+Css+iLqYhMBbw0gnFZPVntctreW0pA/OIeZFRu
zpNFoxU4vLKNHeAvBhTGGsHVazIOKf8Nn5etZYLWutospc9ZckVvNmbwL989mwTp
0ACn27eBQS5RS6/ibcwtHb/FIsTWlNvLEtBtK0+5TFIyrltyJpcaPOV0K5n2m1+F
s4ACFs1hNyjZT4nLfgdwv55KB8BhUGGdP8CHziJBvOzuEBIX7LaSDA2rBt6OQj4r
VSh+OSC2eyAMosa96Eq0UUVcL2jjeA28sUYDBKmxL8+0Y4nU8FSIdSH8xBYuo1bE
7yxsQLsT5XS+tc+9/U3o7zu4bzZMpm7yC30Jt16eQVd1w+zlx2dmuV6OifTpGOgY
KBdLUuL8HvYC0w3toRNhBJh5dJ2CyFXjNImzXDY1gvUDjwuzddudUGSs/hWZcCL3
kmY5QomPIxkf07JR+sgkH1lYrJUo24f8wuR+Z6pv7BWLU7rBkG31ujgHHC81zNC2
TVrfDwHdeIHKYmamAspm3SSA+/YRhCbb2bsB/pjr0djaaKSEroFmTw3tqcIs188d
iqYoBWuvJ1DUxOVAgGNfx3noh4KpMZRmg5G89/hN1v5YnHgQ9nN2CrI7o+ELLq6J
p/aHj4JpzTWUm9S2jLiWUMsPVRpe34xMr5s4pzGkjbD6tnT/qMa9srVafuh9aclO
LIDKq0QLyP6wYZLm2/LS5AW3B5JxZyADofGh2VbWogACzFc3JSgv15Qy5znOSYUG
U6gbb9R/EC+DMC4gbjM3+OBciaPu/dXzvP6K14Rk65Y3DqkVoG9ck2gmrdXdhoWy
AxEQGQLrGmQbh3lyzP4eRFG9b6heGrhRMrIxcj48KsIdJc1NhSlgtV+kPrJNmwQ4
KYMF+/6kycL1QVRE4yKDHkSF5pMlIcgjYpfJmLUPajXeeqvz1G/czNcxyanieYIf
LgOSPtvhBveQiV9AARWkll/TspizvOYXC9vMdGH9C23vwdJn1ivI+gpUn0tZ8dAE
13XgIUAeUnMhkZ+Br45v/Q+jNOxgy6GMu/QIDOpSt1AO/Jn/Wq9xO7cTtiepEWzz
mZtcL1LU78hz6bwKR+d074v9rUZXqXT6kTgaYHPh0iasdHuFG2z6KUDL97uQIVu0
vp2Sa1jh9M2MWSREfLM8I8iNdq5VAsp6YFqkolXq9bnrtM046mGtTO53n8dSAD4e
a+9443tGc8LApFkAJhpSKiM7dnYvAxZgug4klWDs1qfRbS4Ubf+BLgxF4VaKGLa0
r/hb9wGZIDS2ZHMZLE8l748v/Z3PT40aJjhIHPx+RHk9is9iWUpWz30FvfuQaFPg
KNNAuB2TkC+/Iou/SvuwZivvfdU1TchUbdnQIvCPpdBj5bTc8Z3dt+K4C01E86HF
fc/ibmAjgVs0D5IWJMkdgPTPVcN7OPBI5Rrz2r404Bu4eE+MMYqmIWE+W3V7D9Hc
zOXEEb8c/tkKBQSKZj1mAU4zWsHI9/GmmUSNABvCABVP9ptBHYuO6y6w3YtC0Pa+
hjz6h752cyPIXtYiPSA7WLrxMSR78RfGAINgomXHLbbnZv4QpgZDd8lrJTApPqbg
hybtCwLHp2BS2A+HH7OlPv6GZmS5IoEJMiEtWSsoE7yHDTH2H7a5+3OOnWP5mK7m
4woaOaEu1IELsM/F0lBD9BSdeGkEAD5qgwepdE519Xh+YbpLKweZGYEj+xrdMDpo
WjpOaJcbzcELUFnX08T7fIwnW04QQsxfqIwGElv05DufHaUeh7W/AfOz08ZFIJyH
Ob5ciAF9TTNzexfU2x4FYHzx97MQ14ecHka52V3spnpRyAvw4bs7MZ3U2oYDxNhZ
/oVe4Z+1lPGqFo985/49I/lDGIKQqZYs+4FagDUp9LXGjrmoImlZnTHseg1NYBA6
O8jP1+aBIjFxFLIohHHcYUcs7/DPdTJMGKZKGrM1p/R2AGrJ+kb0JeD39ppGr7fZ
qXkLWK08rmZm2OeJfNd/qXlicmXcmAaKuI2v5d8RZcTEpacTqSqmMIQT86j0S4U5
kRUwD71OJ87d0uxBQOrzNhcTwaahvMoO80t6jtsY4kt1BaCREYZqx4/wGNWwqYs2
i/GXDvjjrSCbQD9CS6HgJGtAVKaxRCXmHYeu/QPF64t28vRDPM/C3xEYht5KyP1Y
nmT1YuJx/QtcUB+m7i2Mp1APwnHN1QQLVMJ4YTBGceb2NXnHZ+KykaNR882Ygu/H
PArPOgZ9qsOcf2w0yicGAAQlxstz+/lRq/c4LkfTfPyyZOeg9YceuCIgzq+Mp3G9
cLCwFvM96sh273W13QrjeqNX7gCf/Ne3KHQvEDeeIdPGGvOCkuoBMLaRgL1gNKH7
LBW9/O3uUu1Whh9HXLOWdHFwasPrLpEcH2mvcyS82rC1riGAn304IaXz24wBvETM
xLPleR0A7oW4yqYkyjvpuHK5nUO5zdEzSND9+kMBfk7Rsp8qlJ7vcWlXr4m0GA4G
WgTcrJX5UhgQVOJf5joa8t04jjKU2Y3+0qE+OBPcIPR62NUCHYiCecE6hLFrV2xn
TZhNaEchqPbNNgQtqXL8Vt0qv5jTmiD6J/dAzhEiF5Fe+OQo5jNs43z5vVIghns+
qNG04JJeHYjTls9STpLkT0URqlwwTYJiVyPiNJEu40FHsFK5NfEexgR7qtTsi64X
reNyg7dQsnaCCxQo8QA3PqFEnx1AKg8W31bWLvVxWgELmAubAn0g+6keZq/ZeNXc
xdDteifjaGxyciSXCMyhybVuj/239kvtZYG+qsqLy5vZVb5u50rOTtLZQaeVKf2t
LdZzhXh6zctJiJumdU6JldG/1NESMCYbQ3iCkVx4igBuDhQLPbAkpd5OmYQIqD7I
`protect END_PROTECTED
