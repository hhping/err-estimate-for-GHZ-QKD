`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wq5co+u2hVOL/uhWV4AP80SqF1EzCJ3lTcg2WIYi8xskMruGYjz02GI+tKVCIDGj
0BxO/BFRg4tvnl2vY+JjlfjMKmFgI2feHYQ2uH4P3LTOYKL8T5rVUvFwsuKhTCT8
R2WEy+ZqavtDZyfxgPs9wdCM39sIuVwIUcELgRmygSLu2jQe2y39zszdb7nC8k+3
vvmW6FR+q8VTuOp7ZYHzw/0wZL71+RYJp+a3HSfnmS5mi6S68sImURCh0dHUsbCO
XmnLW6nhZrB7N6ezhccL+JnhI7YR4leUG2x3C4dZ134qTO7CgvD673p4P/pKvFfA
f8gPJSt5A29WjFhQRIH482h05vtaqCwp1Bi81DYFIKJ4n4wghvZuUzDFqcqbZmQR
tvjlx8VinxPLTTU5etgco4x6LNvK/WfQWCsz3N7aCqtX/7GmVOUEO2KN5O4Cb0Lw
rvQ19x1KvlaxnkkR4imjEj5kmEZ4HrMexo5bf0Mr6uIHtrHDGT6lwPNhlmCuw3pD
YSmxWI6+C0jwNJl8HnhxmFPgrZrxpFSKZogK8WvtMexikjmWPPr4u0xu1rwG2uCI
dImFDzdO1WfnTJNicPYHtA4wAFRHpCMkIfeIvrW4z+vqCMgD85dai83HRhqE79p7
FaWAMBUqj7KoZb/8tvijssuu+bdrAqLXveY9IE18iH10eCSBrK9TJkQ5QS4qZh9F
NcvVy/gncOkEXfoIUdWZ7QH3BkSG1A6bR7YYgvLrqquo3tp79Bykh4S44fj50wwr
SuBRSxYeF6uGrvxa8uW8KsOiSHGVuw5st/oOdJML1dtUzLmSJG6Gu/3x6iWp9EhU
wIUbAAYa4YX0HGl9SrAf/k8lLiW5CkSN7pxrDM8XtUPFjcW3Tk5ueGJI7AC1yoVa
ZpHPWnc7K0LTnF2EhPnnRk+NMO+r2a0kjdZTr0CMKBiXzuq/+MgaeRp6O4AkwTgO
uM3Kz2Xkd5k7SriYKEUzax4sRAlxEBnFkXXmVUA5Otm8+UB++iTx6uG6vXkKZkG0
ZOyFxIa46Icl+hoqf485yiOPckUe/IBptghAaUCu/V8aGPlSwkZYkrJlZhAJ3oXy
E0MlGi6rWU5ebeC2VNzRR47zSx6y7scEeT+JeBL5PFY44Ks2S1OJQUYsr7cH1RVV
Y/n0luY+C/7YDtfHEVNNdDxvhe0WLMQDBeBdd2f5b+R7Sg/cmCx1LGhVJiIVZ9AB
ejKLpDQpgBrjPVy+ApsC6rK9UV+cfkSj8MOXt6DnKxj+4qphnUvj62EW2L2lIOYD
EEcFu7CClXwSDKD6JdPkRIKCCctSCvEAf9wE56lba21npIgFg8xlfhzqGDjArCeT
jfzAs2kv9O+x63H1scDGqrO7cMQ9vRPrrdvly8nOKikb4YSnl8pdCWhxkICbdzZW
/kiwKBqIgCs3lDZAdvDTiECUD8XYdDCbT35n2CsMszyanwJ3jRv7Edc6Dufa2pdS
0vi4AQQrtLXe8BdokWZvXdDkeuarz5DxaelyjKzjGGHbF3pD5d2Y+90ExZOU7opV
MRKG4ua9jmczskottt63qPfrGMx6qNmaq5vCCdWIcT5xLmBrvsPCy97LLejzTDQX
59JrCSs70M2ekVspF1kf43Nlvol5t10UCV/fgtpR9pECH8eWil+a1Nmuv9hYnCZY
SC794KkrWnLteozZqVq5CkmqkO4CBoer4QmEUbZ8JS3hkhcrbZ2e50XWas6SSK8J
WUxGUxs4R/vcsACDKlU5WAtruwV6gy2HKwYRMd6Mlzkasyp2NVKYzObByvtVGUq7
IUv42h35NYVpeHL1aREfVFHptsXQAwQ/GV+WJjMOVU/HvWNgmsTvW09h5e+hxzpD
Su+bhHpgwgN2mUH5GojLez3rtHf3z9QMmMLpTkevYdkWZKHZ/570rCPqC8iaTNsg
S0Do1UvWIU7Xqwu+yHQfZo3FlGSI0SFWkiBaxuQyCECQ+mw8+WjDCwmQpTmqvIHd
8gaFbAeUUz7h4G70MUIG8rv6PmZ0MtS6RHtKq1tdytIY7YLE8tQULlXE9osq88AA
N7RVvI671TlQr31gf7PMUbxUw4iGAUcSy6p0Wc8FsuC/JTkScRlQjlYesIOxp8uu
bZJV51vq//0QPv/I99C0bz/LhQnqwVhPfOVFEw/rENNaR2DIBtalKQqR1MSunTRE
En8F9CTwXpsycJt+2mTcyULL63rLrUUeBZE/lIkfcs6Ub9qhT/Gv8htzmpTw/8p3
bzAtZNBqdwQKZKJlqCVk4WoNrO3JWL7rDE20GCaW4OZ7dk1wS187sf+QWTylVY1k
RfPqPtdjTNGGkGoVWxX5DXtxEokgNHdmvr+J3VzYKDQs/shzyJ5wJswxljp1eoGn
zdRHpvgawgQy8d5NUmVRtNI6+b0sQd+wc+AW/4L5MFIBt/z/X/z4a9cyZw5T4BwT
B8YzbGuqZJq670Wxf4bQUn+peyXnQYY94PEHNe+wKZSy1tiIrQmoOBzO2+p2RZTF
KRfc0o8gzHy5RWozitmQnOtNAKIhZggYoFqkqmS8HdzEaAILLfX0oIPa8vt9QJeQ
JMUjC6mRDyUt7dPfZhRVg6kLCQsZdWJx0E6VXvUeMW43dyl7nI2BwsGKIbfKWbc/
35dfiMdgOXHVK/ORB2cqEm5YigDVu8YUKJfFv6JIF4Az02FwP1iuFQ5jSbf8uN0s
9GHmMxFjjiGMRdsr93q+8H+WUWb2O6I/0kcg5QiDwDpgHMulaONNyWm1mpU+MnU2
zy/1A0U0F88GAoUB9z7WluvBfOijKsQYolyIEF5QUU9ZBhOBlL6C/5n0ko3IN3Dn
8kMEerpJ2xFZlLD8kTvD79MJAJikc1HzFw9KI7p2fFc=
`protect END_PROTECTED
