`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+o+r57xqXe9sWW0eYjQ5oGq3yMccPgB11XdwESgdmHPDD5KYnjIqmzUxEIpd9JSf
IHj/kIR8BhKfbgVfnygMvCTasbNBq6E79S/xkgCrQV8kiZ5NhRHAI3h7nY8WuvMh
VJUwOG3Lr39YYuSrYFNE7wudxvViBg0xHpXd/AT6I+gMso3LKpvI04t+EPqW7HHI
ZjuOX+XECzuw7oLc2ZMI8D3ur9+TjVEJrGjAla6nbdinNQ4A3XZGQKwEP4Cr3oY7
noSpuSVUXQ5LnGx6DLdalGjHBViSTTr77TUlw3TPb9lFQWgXQQva0cOlMV1yF5Xh
CAsq/k7VMmsUr0GwWJFQEiz6/fLQofOR95y3KgFgof/9uJ/jPLJjnsY2PL8rSQpD
DZZBslZV3EWGj8jcI28eq9Qs+Th8D7HeD4yF9vl7DqAV/0ajuEnVRMnTy+gGmf3j
1XOrUJrNrOarjFfVl+PCHbf3nIzloiQnEugehaKdJSa2TOu05PEejddEHhG9qPra
is6DsrZ+lAicCK9gXPrSHS4WQGiycXJiaH7n20uKA+perAwWmEtEuKdrb5DlxPN9
KwBM9A6kHNB2JGMC+mGm+ww5WaypVovejTipg6Hrg/rmSLD8NeRI662Dr8SD6nMo
MOzJgwOaZhrde4bj2FXCHsDPjLHkzXPNKuqxTPQqRChqYrVXdoW0RJWB2q9hYdf2
dV5ibtn2KAF7VCFquGcJlbokZeZvaHEbhqPeOCHF1y6b3D1158x6k4G23J7XBpcb
arLDQJfferuCx/p5thbuLIunT4j+1n9uUw9t2Kr7spn8CRsnqdOMKIFEmgqYlqxl
2WIwy3drly+kFKk3tePWKQ75jtVw22lpCrz5eZMYiKgSMN0SOdNCcnW46HJGjZui
3iLngEV39gfhCC/2F9+HieYQa8nHazDZAtwU9vJEFMVDyuOsqlabBpsPAaZyKETe
ds9N1kYzAVVogkLpJ4s0KoVe2EpCDIKmZCLnXs0dYNNYKK3lw8im7u+MK+zwSN8A
FqjM3dqbudaKVhfyP3sc/t/BJqqjMeyyhC1vSLcvw1eTdJAM+UO/ePrUc3kEr3X3
L4WfFL6pFX5t1iJwaIOy+AQ9g7Rh4MdKP9dx78Lp5VgKVh0wBFXo3W/cWzCNZTca
9WtqqdX2m9dixI08rKnErgvV8wBNFq2IP74xoV9YEWr5ymppLPpxv3QzEQE5S2x0
cquezBlTD8jbvKGROxHDnU0CPfOh83T4cjFrc5W2T33xh277Kj1Kx6fJgKALaee5
gWeY8UEkk12cJl5D63za7k1ycSpdlhNnj/bfCK7J7j5SqHBiZnRFYkf4LgciFYkx
8ABwQgN9s9YL/l7B4fi3eM92lGyrBpZJATbG1NFHBiVk3rYlLmEeiHbzgSLBk5Js
aDOxw9mMfDpv4MSJVZ2Q6Vm0ILnb5dL/HvaoJij0b96q2JxgmQulnqeYvujuQJ1U
/9zSj3ezi9YDufiqlyigMxrQJpuSTAWr659TWUvLZzdSXn/6vS1+EgGFbEUYUJ/S
VXfq9d/Hq71w/YuxPp8EptvIgIVsQmicLQncmufoejZTqGXve2Qu7hTAisG4O3ZC
deWTGB1i2TMYouIqQmqYp2nzPhAc4Ap+ps/qzbx4ARK+gLQZWWQZeNYSsd6R89mi
hCuCt4XfBva4K5hAQZPmVKt9YXkRsql/Forvg5ENnsCoWCPASxC/4KDlTt8WWiOt
IfxzN+KO+j3TIJZppxdtfcBw2bvCZ+5Esa66d2W88X2pK/0uoLWYOkTdfVKZR4D7
EKyABQahWnjksGhgGIGWFFzxx4R6n+c1HH3Y/Nnt3GoQq2xWCImWzMIcOQQBGfze
CEH/dkFa5rY4OHnLe1mXdlT0Pdvd5YVFlTAUv4FjLrXscMh0jfp1vB6Uf6Qqzo9c
RFCxuL6Rmee3SxIl7QLxOLkdicXUo/+eZ/5dLssO90NIrc+3aRiXDbOT9DaOIF+h
jGWXPlCxlbGzNDip74mndzDy7o3qem3gLPUGR048pAvgXRigchWwuhJ/ZHnZaWT/
R0aQjof+FI+PDf1WZ6hU9cnT63r8kof+9oyC1QtXr9ZxUF4vLJhiEQ93Ma2rDFJl
Sgj8i7e8sF66SqMzt+pXxvWFxJ2debHNGKRLoRysjs57k1fjrieGp6VdFv1qsoW+
vlF9nFTmsZ/XlZqp8tiw5l8zrRRUjag5CCA3UEUKwPIQ9DKHIi80bDUIvFqyjKl/
S9BNDVpcD5fk4DLTqelatXuIQv41Gp0D/y+aJ1pz/daewhaDRkklErZRh0hWm+Ji
SKDsWYqBKIiMZrtUKBDd/Cg6SWTVq4k7tdk1JA+3eeQ9YnUpV2fwJ6p6prPnkBce
j3/I6YPsuI6HiIQ8u2EL7npsRvT3qb66VDzgEH0xNd1NCOkqlwuE22U3DZaXlln9
vNoh1AB39pgBA+gQuyjNcTmn/5kJ1oIHW3ZMwAAlxek9Aci/maE5+ghQRL9qTSNw
2oVZKmFetTC0FfKHkYGgs9oWSs7fLV8AsCsN6hsBxd6xvASnv84gpnnuZ8IZVSd/
shGeJGpBwV21qXWdeTKXIW7dEcwcV16R9QX9Q6KnFcCa/tmVOzsKG2ZUmDZcq1Ty
BTu++8A52M3UAm7myrZdRY4MytEV3sy6tupwi+AGsyzzTcac6JvZdqz7hs/GS/QL
jEVFtAa9b3NAOBukv6R2W2qnXLeRs0Z/nJRdrwyVxJWlRH0ykSQ95+jaG4hd9RSa
zxYSsR1V5JGp6o3QsCO/y4J3iO4HMoopAOVy/8M+GWpzM9jv9rmOK8LrmAZGItLg
GcugkUCCaj8FIQL6GLmaYbWFe0URIZUzfp5VhU5UINqxoA61sKF4FYieMnLilzNP
IQWvkVEHFbi91UbWxL8xOYuS6YGg8Pp3oYP4H9jAeJr842vr0psqfvIijsqa358A
VATaAbMKxPPvn/+KTuxUOws56TWGtmVLoFBrgKOANW8BI07/QktQ22OcLCHaOsve
SvcbzOZipEnA+xHsN66jv/SeeGJAiem9u2fxbfSA9IS+fNdFsaaXJeZRFiFGEFWM
MrcUKFldIHI+G6nMC4SporMDRJXcwvcb/AlcLpADLzKLJqEWH1jKTlztH8Ap9DhP
dcWZTPo9utQIf+12sPi0yLndyIJRq0tIiq97R67K3c7GGAqa1MzaJb+X/ODivcSd
U2IFdrjS/TED0OnZfpxKsdmb48SOW13XiCLDaVOeFsjo668+fdbk+0yfbPNBCtRN
fPb3+PCkDXhMDlFwlZRwOSD9GSyLd8GzCkO2l8kFVRc+dlgWfyn9PqSL10hf2IYr
mcXwqNonrePmJFM3aHfxa5s/G3loX1c7179lYfb90wuLb6z/FQgtd3UxGiuglg6c
ssrTXwPN76MOhzx1UAHakqhSyrTpNtBUHKiSWkHanVCpR+Gs/K8Ncq8ZyWoSfw7o
V0VT+k9a8EryEbOTO6OteJefjZRqtMv3yyJUtd7jPPOoecItRPETuiw3N0LQxskA
YQhZdPIEvuVX4q6R/1ko1ephvVZU3pxAre+8cdBvzFRegbldF5jBiei6DKyJFFgM
PfmKE6itaQaupFbPmPaDPe1rq89bO2zJ2w2sXki5XweqUmO+CU5IMdZYTjvW9/P3
tF+WHR851sdNRZAGQsmPTPbkDhIkh3PWksIOyU56PYYaAlIr//aGoJ7aurSeq4l5
FK2vHe9l6o8jRt2PWtqquJsTxzkJrYOeBUOFIwfqHPgrlwHNMKqzpcs1xI4TgSpb
g4kb9R6p+ukc96dtx+DTZd//kOkBeTCVAjs82clG+2R024SwaD+EYbPC+bub5UAQ
+ykB3Qry6xWkhvkKGMJNn49olaVaiVkp0i/un6pgYC2ZZBTUFvNBevZC6aZPho8T
rd9e3vgGzMLs8KzdG8/j7ttGYO99/A9q6+2Yo1CHnAvSj2UZRw9oHE64uUJcxOJR
Aj8OVCeettvzbvK1IERjCj0u7M4pwtjvGhZTnEDbZ0owDcZiPkc53pmFk4kIrmYd
ej/JwaZ6TlqHLNd/wAP4Zh3AKNnykKFbbFhiC7cs1b10t0lugg9gpzosNybyfRme
Hx2OfH/TpIY00oU/EqEXRxXqTqUjrjZ0Y9+GS0h5VEWcJ3aMw0yWc+e8Ck+rgi7E
Xk42iNE6e2tKEs9cf0vflC+TPLDEkh0comDgNy+XVtkyK2no2E/OtjNw2JSJaidI
bYJ31Q+CsSzls7ZJattmSMEAgYiJNv5iBf91sL0+ePVA1FgphsmsrjEPkKEGnqAN
WjhvzSbYIhNl4xJkWmPpx0NoZGEWr6hXDuNuWRVHvQbO336x21YPTe83B7tM5Qm2
FjzM+pgZZVNm/eur3okNeYJyHtEqgpVT9f8l93CdAJfB6QWliv9YGyo/N4ao0ONi
AnK372xm3P49SiJHIbU+C+YkxT36ZbVXbAsJYSwpL/8o2wxryMJoeZtEnpyjs2Us
q9jHl/GF8/Gwd1NUVGZyJzbHqpNs/lJZ7k3bS/S8bS41bVB+5/ovRLuUbUHfKdbC
WIAU718QvDGAG1r4EyGS5t+xUccj5Go85IoHtETh7Cgxb2BZzmBF+pnPezxQQ/Cg
m3GSIJKj5G7UVVYSXPrYwihJ0HTlCCN6puZNM0vOQs2/sY9BgQxDWzEyGp/ws5e7
4Qel6UWTUAr+HFwRUddvhvZLmP1B9iT4f14kYEF9GJaVxP4IxTrt1NQuDRV/Q+aH
yK/DPmgoOH5Oe8iZ+j/YmTMINPBb4LeyGvO7u5fJ8+mnfMbXHhiWoGF8ZQiMJfXu
GTXIkfGGFgF+b1Mrlir536dfXdW6wCtLH27I6CG8BST8TSVIppYg9OzxbASswChd
qiT0/3gCoqTGcwvgVjTwRHbG7YSR9hRxxcikeWC1n93XSpzQSJdt/bOg5hK1u54M
FIZ+wr1Teugaikrt91TecB/nr6/ifFOkoJEaoDV9RzNzPOgqsG4Xjovg7PevDQiR
tSL4rbXc0SddEA8ePRwLijy08IvhwkBLh30q9agoEysGcGU/KBxL7iVn1xBN509T
Ns32BAcJQ5KW3910uzUGoJv5QxLHampLjlIUIm7f0PptZIn6aunmVJrEPVN+EkF2
jRQch6ckh/+0WPbeN4xhxQ9vgag+wlSgos+boSLZgEOmDvgNKJIXazKAMUGOcf+Q
QFUnSbMqyJUZ59Q2Pb7JvREHUVYZqIkobIkOckBYCUMVj8bHlcBCqjB/AEm6t7lU
g2P8EbwRry19+HA0VHqrsoIWoD0BhtZVtCjdTStsJbxxt53QQZxaMl4x4e5xBYiL
fNbXh85dl24ElXtd110gJwtIUfLHsMSOtBrehvpq8KmcgTTdQZEFXo2yC7zI0B4v
f8zrlm5oSnQvcZ5K/gOio1Un0kVYFVSs3LBZq7/T+5icJXgd7NI7BKyllB2TULO+
ULiDIdnJmh3mHM4pR2NO7Jn5ZAT5YN+kS6wQV3avKaPJWlGfGBCcWhJTSyAvWGJR
yYhCCdSxN0wz+rMkRT2pYop30MFWaPNMTYUiYSZ/xGUtsvWCDEJqzI3BXDD5AkBU
1iK84gpgDZfueQhT7/WTJQIyNUWNgbCN4OeaO8fFbD8IBSyUkIX5eMCAxCq71kiq
Aq1J0KV5NVuiqpZdeGxguiPqU46g5apVrJ2seJcp77Kzwb4r6h6/L+WojHOGS0gt
x4RV7Nrm9GKK3YdgEoGT0yEJ1L6SzQ5nsBZMF2XlsYsH4xrDvFX7UYUomDNvWKiC
PnPIyYIUK6XG+rP89huTk1oGHbctvQws4g0gFy7PP+Oe8t2/YAfTMMwbX3qNhy7K
yfwhR2+P9Xp78ZHCRu7g2enjRRMdryzXevElMiSy6RO4Ksnw2SPP9wt44potLYC/
cuAqo8CDN//C8Y996wYxqGHrE8l+9OTsCsDPsDRDHyDwLYmmGnBC9S4S1rj1w1Me
l/lYV9OPz/KKQaBQF+q1a+3BmyvyTBxLyFXMZ37cJNvTPGdS9AiFjbs5hvrnzVxm
//GwQbxHGoVoxzYQyS26xo6GSo51pSo/I50k44g9YnSWiKDcU3cVhIOcdsm/XE2i
ul3IDjcF8NgRXOX1LS5CGEdScPCV+paJZwgycBDAdntPQhOC1TW+UymOpaCEhDRt
+OwFDWdYszE5SVJlj8FPKTxtDN2IfvDRHALhUpi2W0h9bR7OdVbeBi6fGy//GMus
ENW0CicH4zJ7QohKJsrkfxjm4VvR+QyCDkziqRrsftCfOrUwoKUWJUd01F/rjZO4
zL0az+ih9JtzTiSBqY5xoZUJmoQjiRJsfjqFtB0o3XDXcd5nsJtKjhSLqOzhijeK
PnCES6mssCXPb6M3JG6+PjhYoy8muMsrc6MSsVjVkTrivARCPJjn6N6iufrRfULu
C0Ao5eipWhQS5w1jmsM33cG99OEJiOUDjdx+NLn/PkYz2FhroANGZjA2X92Bchs3
rADIO9RszSeIo42FvFuIjsiZ8mSb19mx5mv6R/5uK8df3UjcG48QopkCUO+lzDZX
APxUBqlGQdBHXdB2NeLknF+ay9XzNJQ/tXEkwuMHCCj/A5ZwO9c1JS1+fx/6fA5T
p36/9nXA8cztppluB0LscA6s8rAJle4EW7XsCYgEirCErUooQu3n3YCFTfYFYUs0
1DEtQ34G8I3+CnFwf53Uhy5OUMXgz83ssVFZczt7Yt8QlRETlCx9XEhyME5nV6IX
fJmELUFCVBk6mP0HZ7LciXF4Exeq7PlI/iVu+z8+u5qKTJt/SAl1aStvK1JUpTH4
DbeEE+aDY/00FSWGCRR15F/dki+NsnTvh+knprOJ5WlVv31Jw5oOGtu8IRLlQCjw
AXi9KRW1OzWLPck2/GbZ/c2hHcpTuELQTMZ7tlPqnw8E9FrpjWeALPumAemqRJld
b9KQmvqimMWcP214ROea7MW/oI53A2irWZYB+AF08gOpUMI77jMwUrBpX95Vopjg
YcSPwFweP4GF265l1dZlrrpMdGyMZx9mTWDbWZfQ+4Eg20EhgEwTicVlrwM72Fp/
Q6FYAw9N5fi+KsVZEzPgE1LbnzIy7SWnIpmA/4Ih+So6B5bL7z+ZIdVmcuc5uqnT
x5/JazTkoOIiHuLo5l25jvOT1B8fPL/rA+Vam7nrxaFUBS9HPY36E3ukvVEtLxes
NDtH93T60hwUOuWiUQckC3ubebRxrdW7/AZX1m2VPh1YAHlONbmz0WXq2J9PuY7p
8SNbgH1pVNJQnwO2vMCGkbyq73ySJEMXAq3Mbl7sPUWxRL71R5pW1kI74Ocpnhpo
d8SkqUdC6GHMF33ZHL/FcylUul86RhqrauvomZTBV7r4MxI2eSUFM57Wx7EPj1kO
HT30NcTACM+qSuU3Azy4R/wCB+uTuCYx2QWGB/IRWpQ/rdhBCI1wfo4kBda+i/iv
ArVt5V9WD3nELTcUpRufp5RGh7qib99FdAaahVzDDWGTlmuHZvtNN+vdeAVQBgYC
ClEbQ3JW5hWHnWCnaW6ILPw1MFW3GdzVnpwpmJlBLEYgcTSsvoW4Ntm6jaWcECWC
vkPbJDYzjP68udyBeflEmG8VmNStI3WLtA5GhuJfu729wbec+IPjJO9WV1Crm3BR
SmtH+AHhHEzjW4xX1gF7uFOZCt3rOEb91AyoF9kjntC2AjID+iwfwjjDtshdrUlL
K6LLUmAvJKTFJshWDrHzRt/y+RS+8SLDCBLuI1zwP7n32jjtXXncx6qtL4Cd4AEa
c9PP96zDD3RL4+pvQlr/K6mK86nrlfaaLkdpYolieQRwIvoEs0+MaQ6EdZE2X1S2
zaiswfPJ314h+02U2F39Ph4iyjQxw6MzIqhMIvQIPXfvNpZ2hTywMiMpwclVpN5F
wGUyCMjf0h+emUH/1w31IuGY+mEpv/1A7VdKzUjrhw2SkS7QkWuT/0e7NN1/6wk1
3suLsvByoi6e6X2nSkD+wgWJvgkMhy9wJ30chG5XEunMp/D8JqGry3xMQVKDX9Jx
PyDmByTEO2IrPuMYc3Ia1ODgtcFboMJ2CmZPkbSupQYsrcG0PdWsvqDhlR8Jne04
4MdfNanww7ncisrk0l7XgZjGHT6Zp6v2C9p1H4wsRvbC3h8dyfDOVQI2vaY38QwX
jb01Qvtq8U3unkHs09ju9+MrV+nq3uf4+bTK35vVOBdubS/tWDRHtYw4PEyYpVRR
DnwxCyCXybl0hhAfQZ0g0OSY5wQtSIScJZeiSmSTcAhJBoHvdJzIUm5+56OqEkXc
JwvPQli4Fqn97olE9DtKeZqI4xr+4/2UqrXpTBI0Sje1Rjp4L3Kqz2foXoFrLpix
notcB1MbjVoruiVsWt6Hpg6xqQZkemnCMSD2EdifzexxYqCHphHNcC6eIhLDMoGI
rILSEHKCPEhSownO/Kq+pWqC8AnBxo1xrbVbMtiYpF7egjwg/c742rQO8oRJM9TI
a+v6ZEIRJ1bUry3SxZcMnvlHEU7DUY3b/H0t1Pk47IWvIUCSbtoAJQMPwXvbguMN
FMgENNscryTHpEZCN3mTk2CF2hJgVZL5oxCV6WO+3LH1qK86WPaJrmqRt1ry/Prn
myiITwjIMiC/YojtoHk9rZd/diTdfyzW575WJn7ecdjGWHMl7cGOpnBhcUj9jWZt
FvwpLc7SKeNUzfL+hPpQDuQQF0oqDsbUZOU3IAkK71axfRLvIrHXyzPJiSX7/Tcs
RUj+cO9fHcm2EBUiuxjxuIP6BMIymRDPLalryNfUFClZPW6O3fiyzO6+FZrL31iM
4bDRmjVYxq36zdWHmLCdcZFpWXdTq3HjWD1R29bWQA42uwc49fHVM0j5sLM9iiqm
nV6UcMu9MpIO4jBDeb5WkLMse6AhcVyf7DwwMOy/GvfvYKpTS1CLoVnTmq90Jjih
5cLecjZI8gyVjm5jB8S+Fkz+YASSeINDnc1i4vk4pa7sa3QUeONxKUqgLrAvQVIh
Fw6WJWfB8QxvmA57ZExW0cKAht1W9A4Ul2zrQfxHlT4aU9pEZMEPssfS3ZbtfyID
C93olfeAbYQ8caBSAfk7UUqc7QZhjBDnzXNZJLRpD/EZrklp2+jDo7oHNYR5vKYA
cpdqYuwbh7t4JcQq4hdCzU18De3nWUm+vq5nS2KOMVZNCFe3+NTXSvV0sg1AH+1x
fWQAA66pTkKsxQkSMw7uaHXrXpA87ioHNUJc+cwdVtR0TzRJg25sUyJm5lVvocgc
gclxrGZlqFtHKXvOqMsN1vVIOaVw0kbui8LHGLuHftkfxVgbOAf3LCyqbQfSB+8U
yU5+nuIFeRicJp10zxkDcu4qPqVIE1X60xE2RNax/i37jsvkTdQHzXp0EUe7Fy3Y
v8T71Ybd+oy1cEDqO9VPlJrcAZ9JMkSMohZVJ7thbqGFJd84D5GgEXfkI2n596M7
wIo15ktTLUsPNVSGncNuEQnvixtW5Ne0vzLzDgD30nxut90gMyXm9CZJGwpdrHWc
NZR5KYDNdLSjZQ+/uT9JIM1hfPq7M5YHs2LCLVn0m/anb5E+zRR09NSWs3NfTY8p
dhyuFUHV87s/MzFLsUMg5bRyxo8KIy5RcppyFaS+dTZ2COGCoobBFd1IbWxMNUhs
zOuMXqW6tjiUrxHvV8k7PcaIpaxATBHm/4/J5l8jCZGpreSq98B6fLlNS6NtkSmo
dueZtM8aKccmwHdylvlnZv3enlRExy472mWUE7OYSD/qu71D0xy2qFmY/aaU8Pcw
U6cCxDl/RWGfSZq/V7y+JHr+XQfL77RFQqhqkUKTQFy2Qkhu1X9AEynQRlr8VANG
eM5mmT1QZ+0woyv93TET5awmXrqRduIN7qPFX9NCDLMMxFnV+896fKjqjJmjvaNy
jdN9XSXWP2qYrbhu7XYRd4RmC5VdvS408nZs+XmT7eceCU8uV/ac8771buz9VzQw
vQI1bQT+4bPu4TmNmIFMnKb0hx5rtaOrk6Xd82lwgNjI8KAhn2sLlNQd+SbiJySt
9peNmG/AoMKiYZ6W+XvQ5k02sVPqCLlkp3m8XJ2z8GAKde+Vx9m1r4VdWkByujjP
krY2GBqtQpJ01lLuwUgFr9Zaa/+xiXq/TfoJ9r7NKme2PQJDdJpVQcwBXxCJ65ei
NNeMvsBb8biGoxOM5xYOG5C4nBLYtJYd8sC40ZkR5vYqbYRtXcF7SQwYMD6WeyBO
BkwaDOhWMsocJvxph+xbWm68iP1OERVzjdgnShACHa+Vycd71zAl8HM8TtEVDHlC
t+2joBCweGY6XjZzVTCsWEBySCG9re857P21N687EDgfrbc40MnM8U491MfNDQD/
8gO9NNDlmL3TU8ako/hBaR50mLClcCMZUnw1Tos2A07P56hPgkUltPTkEV6wr7En
J1lqxQ76tPfFoTX/jciVJGEceqXqsic4JRBGAihmfaw0+0/v6KdcLYfigZIs4guG
XKvBYiRtXjM4yGsd+Abfc92MB9/cZq0HQjxd3l5paNmkR814d8mlvfQkil/wW2rc
cBcACThUY3Kpp8S2sSkhCRsJAPCD0D0jQIv/XN0mZ6E5VjvZVwL7M8Y8qMWeLZF4
oWEZeX1Jkomirm/BXnuxoQIAjdJwnFXmi14kv55tk0z2kAl3COeMI4Hbq4vGdw0p
6VJ8ERfSzZ4eaGXniK23pC9FuRLj/9bAZyHEiNbWrUMHA9gri6uVl0/w8L+L9bnu
G8ySX8owDGhsY8tkp4RT2dwiH8rsLCePCyXQqXitFEOHaWZ5BQ8RfxbFMvJuoTt1
bC6E+bxLVbZ0K4+VhbRlvkUiReYsUVV5gqfeqezPnvqWwSgRtrLeXfwYxMg6Kpa1
UO6Bj4PXh5r2/YE80gHsWAtsALdH++s7hsJdtqrwsqYXiXdike/tE0wkspRvTA46
YPu+ldi5+URgaVZT9ABQ5cwj37Cd7PYxORhyIb/3zws8Yl4xwmZCU4ZEtV3YLmCi
rvXGbs3zhxOb7hi/yBdwSq5H9nFsS4LHl6WBKMB7jn4E+wF2FFsE7kI7N79OynOs
o60rmixcVpl7YExsaYWDRN62lDG/zAtqhH++OMMVGqIXdSgO31p4WKGGGLVckCZt
F29hrTdst2psBzNQLYzCOMrPFFgCfmcsy2yZoBLeZMsll2+9aHRxEBHsTmJp0MB3
ZNhP1iT4cMxxw5zK4h8uTe1orqVN1PNMmVctF0mEdeuXVcqrYipV43KDKdxSEtMw
1R045zA8+5MXpPhtcaEfglL3sCPjuiXJ8E72kyePhkdnko7ur2x34Lx9P9mgEL2v
JenVrQ94NvXtnFg/D8GWP6Co3bgjeaVNWNR8hcpvF2jhscopLjykiuvH+Hhyy/4E
qQ74V5FYCX/o4jjhpsP5cmgkK5Cj/eUg0f/umeNruKqx+8vfWQeRDJtZRyCwNqm+
aLEURoLIYg1lxeTERbVOJCDqDB+Ok8PycKUyB/kKRnp73iYwggV6JddAwv9UvdXe
3KJEFZ0fMKEmqHvrnuFVHxaKh+hu0DRd/jX1XENuudqLVbmLj5EyuWF3MdSMJHB3
b7uM0FRYKNg6R3ZktpksTMnRjLjlUTNHYcWj4f6lVFfoqgidT1dRiqQYxu7Sjof+
ywsdCDa56sAFPbGivhGOF0GI7ptKlybuq97xfBIv9eA8RrMho5Ot516IK1zVqqNp
JhFu6YAk2I0KiU1ZTYMq2vrYxAIdNjfHkNpJgNqNhw0Kfl8XA9cDp48BGsi1eyHh
pcO3afhrTw2SMj9QrfGvLBDHGRvLtR4R99gPXNjoBt7FW7Yz0/aPSPIOuixwxvyY
pocrVZ2BcQpWFqT3yPv7j9TZ1mfq89r3Q4S6cAyh8pR6qfPddbbUN9OCmGOW/S3+
blAQEcKSuYq2ws+gDUiHCdcpgYVYyBUoXb1epDvMA/kpaQmxVL/f583x6Gbi0GuN
cCNDhYs1jxzManyw7Knqz40BdxnGEfp2a1L/7Shf6WNEa2a0QLGdylziE88D8Aof
tYvnici7jB6EX0hiTGiUTYh0C39R4sIGW9ekDb8go7tVYE+CcleKvH2vkLcQOt3A
fLLMNgbSaYODEAlxNrxlEa6uul9/HfDGjzlfJoWpP6ecBvU8Rv6u67mxWK4aKV0H
srkMOlRnxvjCvxuvzEpkBPhOePCXY5of6uXSN0q4TEB+YOrHaLGxjfGxMscUdUwY
+8FdBWIx5p9/1cIFCXc2l0YkaXw7A4Nh+jVHetpxYb1nR1QKHCZPmKbm8CRQmcqP
h7qJoxAsVh+fB/voM74ZTPQlcQZjg4g78uZD7SFbvAhYFRpKNp6ksa9oLne5hRoO
wOa1xXDZFd0+m0nYm7uHPucdupnBQgnFCnfrHefo39guee2cF+4tY/g/sVMEwkxS
HoNkLd4Fz16yFPEw5JBQtQm1mveh84TE1Q+G6gSw4FeMVH52g2BWiuPwAQpNc5pQ
vUQ/Nf1m/Mo1EmAW19u8nKCGZux45zNzjKBmTtiXbgYTxZGLn60UG8KGfgncpxLk
q+CJeN8KqppT+24kWZm4ITpD9jP2iL1twIfGmZbE0SDpNLRYkRYw+H70Laf/+3ee
Lyef3Go27yw7KMY6n3Rba6qoYoxvxsth0c8M8JdYv4DvZqUaYri3wx3b1rH9mFbg
dMXItDPcTKCg6dbisrKLNi5d3E4zHAXrQH3ogU3lZ+kA0vfBc5ChdQ4plEVQfvWe
xiPFzQGxfBjhTQRhd/VAunqouvmniB1y56v+GG7Xmy0zRca6AJXJwQ4tGI8uB55z
bAf2ie/Vb8w5BRikeVPxpVvy0ud7mI2S9AuUvEeohJS3g3g3SVxYHy2mAeTEFzDz
CI5Vv/WFHrnizC5fs50lUG9ko5xr43gsI2Y9IsiN75eh9qQGFSGeL22XQFHblu1c
3DvTI6a+YmpAGZ9oua7dMgOY6QR4s1BYJq+41eiuH050v2E8LGbvGujip5f670v+
EAu4wdmsS120Jr9ecp/VMQTP2SdMtGVG/Tkj/rJEzo9AesMrqO0MTFOPHsag7lhc
0iQXF4T5Ss4JPJ72Gxu1n9sECDc2VEFyRfvyLghobT2MV3/gcexfV3zlca312C/1
uv641wmKqohOu/QMDipS7Rv64FhtKd/YUUjkeb5cW2xs1ms3rJTRMtgwCXG+xhGg
zTQ5Nqnwved87zhQJbLec1F1S/turkSLszwFRX+Cq6f6v20PVPhmrPxQv9f8pyKM
rvWxfTZT2iJpLWu7tYdiQI4gHFLTp+toNsSmeMcDvtkuc5vYqna28/gwNlNHQtmT
hJkJHvjVLNMfla0AkQbn7keV77Zflg9ZMTupNEQqmwfotyV0MoqhMRJsq0SDyvTR
O+rL3cT/jUJvTfR6MdQMn/jrfFP/t+jLW5XNtk9tmrdOIPB1dLxbbcB7wFjz+2Sk
0vj4HLObkzVXPWf5B4HiJl+/qmKqmjeV04UG/oKeKJImp44pLKy1tmpifJhVA24m
jtx3vguU4tJYXnuONs8ZJhRCCqUrBGH1jE+z7g3Gv1kXA1S0nKcZko5s8mT1657p
Yieg24aN3JQjq88RMJIHm6RRDuh/jbfKNFygenBFaDX7sEeqYd/uTrvw0j2GRhl9
EnhkY5acXeL/dsJtsR+qh4P4FwGaFsoYKVGfqOgkcVStdpBkrsv7LqUeXByFNl0z
tlMP+z/vNsG4O20voXuEIFL6iI8iVkicID32uCp/aY6IMBGh2aM6OE8Wcbf6TDoI
ndI5P5NfZXIaHg+OjbfA5/lWkVTPW/TEzE7op795D1N7TnYnzVIF8o5GrzFm2+Ev
nWPt0ZrKD0aUKuj3RkDAvh2ud5xU1ZmUSQ5gDZWB3YKz+ExudpbwCSqC3GbjJDvY
kei1lhAQEmn4+drHKvFkkRm7PVTSTdmWJw2qdGhDTaMuG6EmkFc4xR4wz3xKnS0E
dfgs9Y4ZJCSB1/CFgHggJysRUUvbIBjF2NgzbGYfbGKNpAnjAaV1YaA5zNyIkvoY
cBDHLAtmB1rAhAfG29isHN1DDSNqxEHx5cXMjVnDzvM7TMwpKeb6aps2ZfaPFEWc
pFkv1rxsHiOyCHxgm4WVlgeTQ/AD9byTc8ze0UxOc3LP+LCf3qJY/UUXhTXwyfC/
O0G3IohwjVPjlG0OV88OgH9Jkku858uKHpzuQum+ygG4C2Ylig1DwVpeDvzrAQ/x
yj9NHE/lDZwD9yNX5edCu6gOu5HjvcayfE+drdsK0bR2Uv/a/GNozkmisHjGnd2h
sz5OOXr0jN2xxFas2bfChuVrIjE8aztBU7pEpmfDaD6gfY7q4YAS0EPynvaLVS27
2EpUbmZYE1vQ+9p+maVK/+rUFad+LjxCiTdaRuz3lz8JBWgt2u2XPd6P0hH9I1t3
N/7cEhe99g5amqJP07T/vKROw6VwRsE0xtytKDEVu+YJwKJtzK64UL2SZwYy7pHw
idpzHzStJ5khFXhTgPjDjixLt4ej/OZrm74LskqlemAT3bEPYTqubdzaIFCYxcSw
e8zj5SKHM+iirfpKE9truqkismafvSd7+2T2KXa+c0siTQTf3Yf8skLO8U4H+675
ej8ysjSyCjLmv6eKPZ7/N7V7mh9Xd6puRvhUuPbF0pzmhm4RD0QYiWuPnlysZ+e4
NarVp+xw5yOFm3gMeVVBiV2IeXidaLxVGUBizt3vXgofD4qj75pcJRj4sBQiZ2ZD
L0aTTunsAFTflXRqxSp1yzzZ1Xa2fPx/zzOfr71kcIPumG6eketeF/RvbzJu5wRI
ovYbQt0nZcsgsqHJKjEhrMEXgXB+Qew6Z3HrdgMjvELFmDkINIi4hucPWxGsLx9P
iwFtRnlF2bsBd61dRfuNLU1eTtFcTbVKcDPsw0aMOCs5A1KMpzjbE+Y637gaY9Jj
XU0L3+pKUDOwZE2ZN6xAwIBo1lHb/+8Y9qKoINZkXSpFiXUTeKfkJRFPwYWx/SZl
B9AcJTRPPC5+ADx8Cm8ci9MBRIwActD+2Pai5h98liD7YGGmeQCEoH/k+CkZcHim
EcKvWhPsEDBfcL4+jsgN2wAc88wY53bBl6CC0J6nLSsu8pP2ImYhL3WxvsrF+Era
B6a46TWS6Pj6eMd0+IzWhN6N1Xv9S6ljJCB+TEs87az2tyc295/8AtIMJzzhdaDU
DWkxfL6F9JmcFE/tp+K6C6MSoIYNE8xAHzYx+6tlSo8swJztHTuj3FK3zlkKULOE
69lWwREnfUhrOQjQXHjse2aiWOQVGwoKDm01ZIYhA2H4BZZmdJsptt+aQXOQcloA
eZX0atVGvdzbvQv3dUk0BgD8qDvDFi6TbvCooUTHCP0TpCVRMbk/LvdCQh55NmPm
fYjP9qXZS4UgXx0+n+vTeHhOpqu68CYjYAURjmQJ4efoHrrvJeEJ2lpH23ETiChy
IcjtaOy5qcq54adqczjofIdMtkmjtNpRB4qY0t1kcjNPRX5vj/Ob/gnBWglTfMpg
184aDL6weZqGRjWu7rwXhOaM9WL07af8U9cUYHxYLr1dHkUzSYYC5RSEAqaxyg3v
9TsgI+FPRIr466i4faaHkzUVl2r0fLgNep4SwFbA2N292FlcThJZVWLrWWJ5MTJo
4CB/59EYS3dFIHfyiLC4LWX86NaHpKE6wd7XI5NtvuHqg+EZpJplaViC44GDWCc9
hPmLPYFp/DSp47lku7mzo4IDgEs0h4rjB4h1BlImy6N4nieT/Se/FLt7GCcLWKb2
NBhooNWhxA2fwcGJ4yXfwXe91oe1bwaoPi55BoHkLy+t4h+B/rB6fk5O4nnjxXi9
BXv4nYPG9/XYnxS64ZXS8OplTxb1Iww7Hsy2+GSlKy6CEcKqA0F0BGfkVwjeBz2b
EG776COT6UWnCQ5zkPbzJhzl6653Jfb1bMu6+WVUHIUywiFa7sdgFjqaOHfoo9G5
umqd8jUGeek7CnVEWpl8VAaOM2irUT8bnz7+I3LoMsjA4cQKyeahhJlbTE0fKsxF
V5qKoJga6rsqDaGtH0+n68zm0RQkAix2TgaU8igbSnH8s8BjZch1kblUtZFvgb46
NzdaAH0S8LArx79CQbs+ZVRcHNeSj+tfvS5dlheOsy3ERIvyVH3V272FEjOWTsJD
bOcj3WzY5jgpWpKiwYsJCvY/Gu5Jo28+yDQtqzYYRQlaF20IH2aQIYONLi1fi+z4
UumIIhN81TzIVBXzf3E1mBlwTnRlH+VJrrMXI7HHPWcyIZHtHkqcLc2JFfjACyrC
ZV/E1t7hvqWVa28cP0GWccgnuQereaLuojdhHCdZ7Jnl4O/GkPv8Rb8UxWR8g0at
O5uzOkOxhobNHfqsbMJermX1+s4cZ3ObImuiE+fToZtJOySCDmhvvFIhYO4DZf52
dCTB2d+Stmd5aoqDmRWoF9mcEWAAR04oasml3oqmiJckjgJMFD6WW/yMeplsVL2R
DxFa5GEgX/XAc0pZIcmu4lAGchLs+tBxC0vEOkvWoXmOq6IM94B0j562vf8LjbTb
wqUF+//IV/gq28PfrCthbMvPYnsIEVgYwdbKliJsmybgLvhzJEKABa0+JYw6Pu4j
DoV/00mgFMm8WBVaaMZbkC6i9Hj6MUEElVvLZer9BAxwE+Rq9iWe5v6wJv2H3D3m
pmO5EVmtv38jG7wpdNbFCG6BnyoIRBAoJCh0A8LjhOAOMB16BMGVyxPTU6CVrWKz
96uVeUSxw0WobSy/KhW1Scts+RFuVlOX+GwBtH/lublXcLS8OoJLR/Z5ZKbe+eZ8
Ygg5js4/+cIZ0o4zIdFh4Q1f7jLHQKulpPOWs1GCbkvdYpl7LQrCfGDiBiUv3XDa
JtzfaxfUOvXe6pcsLkb2VT4ZOLPgfGitIOMQH0gfzAxbb/iLGtGbYz+uSEsoru9J
PQDOXNp0ZPYXBUY8haaeQ+V7u+y2yqN47qY1rDp/vu/EJfTsDGvDGD+csZK+bVTQ
6JQS26WtFcZVduL65csAve74SExLuG0Do3EzEh7LnG8Csc2L0/NlioHxq9d9xzEy
4+DCoXIhXlUrC9hZ/QP60An232J7yg4ITyoy3DwyJVLr6SFZEavzRxkqlGKVTXwi
qNkPeBpKnkjeA3vXCI5KiHLdG3zxfBPy6gSrZ4mH8JJWpZrsy30p+58CTeL7t6Bp
AcuA3c30CS/nutr7KzLrPnJCOSjLAv1pHoCKL2IoF5NMS4vK0uNgDMQBxvZyxXZL
FJB3JWTj8RSL7ei1F45kBlZMu4IJLFRhTBP3HZMw6GwYylITZkj3kO02ygtsc8sx
T/MtlgqvVVrcNzaa/JRJ6fstfhCQudV24JyoJ+HORRlBD4/GSic9dW/h7O1iaoLz
bfvAvR/8+6165DHu/EvU2GwNFc75YZoOfy5cz9rXsdyjx8L2+kwgKYGuuKJsyYKJ
z+kUVcEV41fyZLwX+hIOmeLxm49bZPfzcJEnlaIsy6TcKclTakMyKkVhvFAJcqcK
DZA8ITMRuA8r0ZylYAuxqUbAeHG9R1uB7+c8XQciQUIjxP08hNE0c3CyIiqxbSdT
f8ZM3Go0OwwadRMsmtgxzb46futSZhIVuJY9C8RG7GkX1hSns4g2r7hbeErzsXz5
C519Xii3AaM4nf0vxDYKi4t8H2HWJDxLxddofYaMQrbPmlJ/7oDLrsNs1koRqAYT
cCuXJyoCvThb/+U9s3O1WrT0qIdwUDC//yPutpddILS8GYXkj/TKuOxUkWagFpPF
tDfJzwYcBzEkSLb+HHqhPkIWPBpjr/GfQ25uQRiMgdOvzBpD5L0L12rE1o5LMg3g
UmS++X9KME1wgQ+ksvvXOyrjKJ6+xjnwFdC0+qc+k0lEgk/VN1RBHOv7vA26V8xE
umqDf902ffWsYSeafHHjN7WuXeC3d8e1Joy5Yc3dcUyDTZw8NmLyf5AuTQLcYhF+
pTKiWDHWH9LJ0wNTijg0Z5NQYB6CuRcomr5VEEd4lKQ5XzNwoA7eOsGkEJBZNLml
ah5n6P+Z0ZcFhu0JI27mf4uKlF+iMU/t6yCXJJ9CQP6wjkeBLdjGASxuCLO/tB3Z
j3Jiow+tftJggx00quKquAn8/C19qKQ2zO1e96XdJE3JmDnwMsJ9zj4ED1kkjMuy
8m7U7gIeyFX7oLl+8m1im1VeEHr6xeEj9aokzr/Zf5vVhJtR/ou/dXncgwCGijU9
9vRWf0fFRyFTIeotmYfWPpnjN/5uzUe0TwuXD8Wnm0qBxvERk+K5seqteHUeLsF9
Ce9nmGgBpNfTVbvUciK6otgdyJ2MRT6z7gqhDZrgIa2ZTKH7w7lYKmXs+d7MBQvj
s9f8QxjO7Ojbw0RNETAY8tkviTGjnAqJ7lU9fhaKvV5AfWQP4PmEgb3NIWkktnOK
Vj2NbfvhK8S6qCHZueA11keIAhQoKarjGrTRiN2PVcI91i2KzDQgMGq5PPjDa5/e
UBrv/IQqJMdJmGTSypQjAbQiyYEvOdvxLt0aSUPuf0DxCbe8lVvG6U27ej3/Sik+
mRRF2urBz75MzdYuG66gmw7eXSxD0709xNbcsMAYlA0StPy6YfQA/6wlMlPmooV5
Z3rZw5opCEOCA7nkMjQMB3j5vLA5feN8WC69H8bUxCnwYBTHkxU1eUqWcLyM0Aj4
kiDAeflgaOKohprSmfBxPPrNOqY2P7yuhjylTn7m8c3gWDf7SWbfyRnGsBLY+oGz
HSZHBXGJPMDORS6/AuPNYvlONEvW90ujtdUMvBiDOTkyKIZeG8JT7awi2CewoesG
AHQpoX5kfJhFuKeZx+IMiu47t0M9MHpC7EoHnxf70EFptaqu+wXwR6DB/Q/IGGjV
egOJi/6Ar91qmova70F6iWOl/JAMif1sLRJzGIVPkFBYTXhPZrWrTH98hpRLOMrz
bOXMxb7tMYUq/Gfs3YOX5qIz8+x+XGidwyd/ArRT9khEFNdQVYo1TlSNRo+7+KbX
KTkw1arh3TN+bsGHTo9ryCJDYsqskwx/Mx9xkxBq8bo979MSvAl3YjZI+ZfUpjs+
Yz3USdXjRxWGIjiHxSJ7i7+ldE473wZyhfKHt+2vMCIMJFkNqt6b/4lPl8rjdtf/
almIJrfPGgBB+cpikraitFMhMS9Gowk6UoD1woMMYrthlWlOWkomADKkuegRcXAz
AK1Sjrsl7ElEXfvA0CAauomINKm7QuqF8s5pRNsJmSGWdQt6uDiwdaxP1kTV0bPN
6XLYHBYvXQcVIf1mili+u85t41efmRp4vYKXV4RBX6bgt35JC7OjxwGWz4hDlqLA
8MvpZHpIzfau4CyjrlqAMD/NnU9yySENo3C1usX0GIXHc56UETc9kal19HpTygtQ
vvzPzwV1iU9tr+O2u/fX0JAMs9O+BlMtA8XhVv3YbaynxbJzXKHOtmF9AY2bDT5f
wu0Ky9VmpseTbzPfN/iVDGCseVMSzr9EhvEhbeVakEtUX60WgryFX/d5IU/hnxq6
9YGnbYINcTyq1HSbleq9G/+LwLaENCenJIvfx4WVjMuPqRMB8CIX6XATIpwKu17m
un6frZkIiaAKzKh+LxdS9sn03ID9lhr/ialxu8LUHBFXskhQky6pPk91M02j1SoF
LB97WWFeC7LYYU+BGD0jCqCJ3DP/u0KQ5iQ2ZJ+ZcZIwhTHRCxDa7cQIoFuHyweg
4iKtfEcoIFL2p0k3VTlttf2M58GBn83Sfa0fKkhVnf2CApCgUeWfdVGpiRhxbK/t
HGLbC5icAZ6T59MpGhXtbmr2egCXlD5LzIHmAlaPKF428MgmUX8TZ7FqhmNBqHjU
QP2UfdltQu8ChypFpKRVQJ8IRoKA0MgrGi0tULcmQSRT4JU/HWc2+HilC2xOV1b0
txUEkXRrb+//7YQs4z2PmgMl4EHspOpUOzG0zezvC714QVDWOUzPDXkNdnE3uvWH
6aZW3YulHhvwHz9e61O84we/gDY7cPfKNnHWBlXOjvxsLr/FZoKAWPBECQu7PV1a
wmedHr9TvS9phXvPbiK7mHsHKViJ606LSmy4twBcZj6RmDUBGOEGPwqdRmllGQ/m
LXRt+n7SkQyQ19RpGSFDtgYQU3MxfYkan/tJsWwqA0RNpKw1I37AHikTAlpVQG3N
UPTasgwW86R5bkoZurhrt/XRnuFDndx2YcaMAZgwyAslSh058RGO+59gAmLmu85h
NzDrSatGUebQQ5xwQs1pP09/Z8vLr96ERc8dB0sb7azObKZRa8q2kgQJDPE+batv
bKnt1ItXL/QCF04nz8MH60EmO6dVCehA6PPDbOtICLxv3Yv7a/vyySrEwenIGKPq
6VGW4j535GdV9G+cjr+yHf8+7n573LlnRoGx62kcdgAKdt0YkhjMME/E8pAzNZF6
vfglNlzpyN1v19QwYA6LwlureUVtVgXxGtXThXng9bX9kqPbDz2ROy7U2ZY47LQC
/cmHN8vUGH+Hw2g7RVDF2tSqidHB9llJ/XaPIVe3QxGgn0FdqsEhlrUyrYyLW4IJ
/MubJOy8MaU93J7zuex8CsgNLCClCyMfV2KqY23jCp79lRSpiRzXTxXq3buXW4Px
VLamokSjl6Y8Gz0kuokO65BbSf6MCJn4xkesdwACLKluuvLkDpgH9r0RwgqUno/f
KmdS1ir8ICCXGn1staQeS9V6w3dFiu33w1VaFP96ziW9A2aVsP6nOtFpqPW8LgkH
WMko7w/E3ZvybUFJxXsLTE3iUOJKqBaGL9/0kNMBtcPbKeKqlUfV9NQKKt5oxnlq
Nd+6vfoFmu/xNYwN2XhykymBY0YgpJXjNzBWSxIou3MnAhDRVUmxs+Tw2sjdwIWC
p686r1creyUZYb1ddpv1xHoq6rA7YZxcSqglpSD4euzFjPTDvsqA5fIVpoY7V+54
vQElCaH3rod+olYTyQxZxEiUbUg58ci874evPWaD/l1Cwxr6CiWL8PVNluC3e0Xi
VKoUZd6fDEPU5LRLRCygaNkZUWG/0gaq2op0Ot0wFWQj6lIkHThaJ1HLPXge5AU+
TvJwcrWHeghfy2tBuGH3oy7LwaVfFodDIUmwDGSQ6P7Z+AS6dfp9LICetHQuV8qZ
24AR0HLeFVfJitV7LbklNJAV4U/mnjQLRKu1P+IPlldz1soynn/yWqEiCPHEz0M6
ANHbTHt33WCa4Ab7hUm3TMAp5V86/lwvUQWA0pUySoS2Tk29wdDPkhG5HKQto5Gh
0t7tYMCLPyIQeE0D0N6h9vhAXqAQuPfYu0ivoY3sA51kj54eUE0uWbeYmVtCcOTf
SI2f3i6eONMn0wvRv2cStHkgXUP06IDrqCc2rqIiag+sJtrXvxGHgGDOXeQ/3jbf
TvVmRnG4aSw1RSTfqo6srXpioRdIo7NXHjsSgtnateig5cuG6GOjAhMOB8SASkTX
KQV3o4HgW1WOFv7tIJm8mH46nB05MxgFwVmMMBCAbqUlao6LpkzmP0H1NEZlXy/s
OU2Jcvv0GK5t33JrhdvZDpTdkj9DOc8wxV3WvSVr+pSMacZWWMPTXKHhkMvjFmwl
0mdPZQ7HLqq2HGQZ31FdsMhx7QGORENonPT/wK90IemhkLwoFxrtRVvPNrBGXhod
caU8aBwon4Fvx48WdbKd/a7Fzm1EGjQ+JJbbMHfUJWriAomJ63gkYjeznbkpPQls
Aa3jBE2T8hIS5iMIUDoiLeWZF3oV2ixB4wAbCqYmWaEXj99neNNB73ILNKcDuwzL
GK67MIipPg3rT1M2F+kbs9q/W60bGoQKJa0cYKaRV7Ue83IsQlNOUfFGGYfHSxz4
mRqskrAx0rLaIMVBhR79lk4s04O4zYQtIHIzg0eHPoLfMY/Zw5VTi9wCwFDAbl++
auZ8QZpmZDwztMh8MlLG6CgYkX/RgoQnoVEJbrH9ANX6jU5KGmUmR1q4RC4rjwau
wOYSW6BRYhfrmkPExdf/6SVOP7dWbk8BW3Z0ymNA4EqV6veaKMI/M2pLcLZji6km
BMf5RxIa7DzNBfZUFcFbJulx6Ig5vZxkIKC1/ucTYU4VPqH5ai+9B6H3chg0S65f
Ursa0bPz1IxUDyTfQgtHg/j7QnMbo28/cW/WPkwIqoYIgXpm68ppz93aKF21Mokl
B/6WzfxWKg+YyVxih72ymGGFjjQP7u6q7//xbNflLmTZmo6Wc0lNODBq62ZIfZYH
zEgiNahfgXxGGib9hTAd/I/4Wh9M92KnN1XrGpectyt1uJvLhdRwxp04Mu01CQEn
OmoVkmwmDIl23ewI6KlnLS9dJEF2YKPe5KT8Rz4rgNIOhbw8Q2+Z4Q7MYdL0F9Rq
kTdXsuKmatP1L5TMEtu6lHZIjjSgyZjHXR1J5AQLOWbdg/GLNLzbu1Bo8zziR4mi
zSi32LRVUmerMUHCp7vJmQHgQUli1YnfCUggcsgd8ooNGTAU7nhM2RUKV913nvcC
v4t6pEaNVW+cWt8vb5XAyMUjLaYDhQYOKAwXovxPSRDHdJZkfCP8HX4lyclTQQ4f
+ezUKuHjDKOXxdDwRRyMZVtAP308hxsZ5QAJvmwA0wSC7h1kQHX9bvQHgeRxUE3y
lSRhfpsDgcNldYav+OaYg8mAxhkpp/8xQloPcJ+a+vJNFf2AGXXfygHDR7KsFDop
tTchjyrIWVvQEaw7Wms2ncg0B0kM9HSXxOWHRGbqZyXadmqoNiGdkvE2idQjDVtV
4CyUNNif2eH/FIMWK7R2p3lw9XbGVNJLCuORFkwVo11irbUb3/FeE/MIiWaGhrh2
OySNsNlzbO4ajJdXwH7gZfPpI5MgtHVD+GHwWa7x3q6Ifl/BOzEqrNPEAdq/XNiC
fKxVudbkYh2mQHTNIIffwnJ55p+bTX4YDU/qxDQU6hZ+rKuMt35d9QgwG7saRU2M
tSpuD/AxgQKyGjCEpGmFVL9hP/CiMfEDHArr7ZxRAPGqmFLGq54LA/GuxT+eroya
Lb3LDM1gAIDvYw0uGtpWIwg7DiDlua2ke73ZvARxRG6w8iykl9iwC9N78/x5l4GE
aWkRZ1B1JPzM/2Sfv0RCbv7GyUMUuiLIX4cZrPnPN2M750hGwLNuG+IGBkNS9CCH
JIfUT8lZeIjdcxZo/jjdqiaVdyFqJJjj4jT9cInwLwoZDDDFhFj9odV592o6B7wO
ONrDfPVOA1f3ukh1j4h4g9XRIQIXKyDh1vBk1eikmWF8lJPJhItBkAYjA0z3/rmd
sWEESGCjF7WBdBk/QdrQOBDmwO4sFoBnGvcJMnBEj42buTulKPYITWpvrS3WHCBh
et9KGrEyDcPLE+txtomu4kQ2ODzOyoYTmFKJ/zwYnQhjHYfE2lh/SeEOnmSZ8syF
KlLP1thyvOC16GAD/TX+Hyu4F+S9E/SUo1dNvCsVC27yYUsn98Bwfc//2ZJc69Pw
ih8+hYGa2Bm/BlFPkQHJ9/fCnwsLp0OIldZ6EttkCSndAcdVXyZI1zfh4M6RbhHD
JxulesbMfud/YB2+7bdd6/NDEYdp9nZb3idXDX+SF+rdeLZQpku9/777O3AtszX2
+DOm9kaGDDpOfhS2AASlKXN1VVYVv55aEcjp2Je3F0YWoMhwIAZ5jtF1JQNob1kJ
wkw4aNXFXkXN+q2ciLmYRsh3WX4DXzi1HuAg7032zJWYUFB10Ijzy5oAzbANhBYD
fuHg4Yy+nLMWolq/PJZZCpb++i2QQIKVzFdn60dqzx0pmpwJ0ZudKg7i36ra/uGD
p/YsC1vn3ufAT7dGPB1Vh+QyvzIMIdEyMgHiJNuyc8B+XZNs1iRcGlDgHFhlTFBw
99K8dIvHpS/NcP6Y9tNpZ9N3Q8SPwO9cLUyMuMTQbTuc+LnuZlLSEyG2yKe04Q0C
0js3wgL0tWABQH7MYC4Arr08Afag3npGdAz9B99gPj7Lm1tHBH63QlcHnczxW4Zd
gDr8V/wZEmEL5IYIbyf95g5AbnaT/tzBwAoh5+y1NYrYl7DlF8TdH029IdWxvLnk
4iBUxVgyavb1UnevSNxX+NPWts7CEZsSedOjfQ4m9b9ZtFpyMWlVeoJsW/Y01sBm
i/94QwRarbQPtQSgSYJxiWFle1OIVp/28BGwSiYUTSIqhAj8xag2yU0sbUN7cg/m
GYx0DYtOototUEm9No+wyr56CZB/3ZJMF0lQfLWevDq4I1fkF3Opz2VQ7OIyQg4K
+CRLYQppn0Dv9sNbLZalzsSduQebU5ttLEYHWI9qgkTRYdcyr3i4WinPyHS0BVub
S8yZXJnoTlISGC2CQaq9OJupfc6m6PeF2cDYL3fBztBy43wTVLr425qKibDEBRYh
3UxLoGZq88OL8R4D3y1p+QbOpvi23YKvtY0e8PU7hONzQHM8ffxEKfwf43LVkf6p
wYghcnqGwXi8A9L7jaSyK5D0fP6xgb20ImsiDc9AYPPXuMNLbTOWvhDpGKZ5VlUX
PAytzkYf9SuR8pchDrAzfNPq4bYuR/tw36h4nZwvqqtxzNxpuTV2f2gzDk48lW1Z
WFxdZJMgaaILhZZ9Pv+K36lHKNlEuiUpJ8lGYKr7AQGcYbV0jJ/E/5E/+8p1j/m2
cewrAruIkEDKDSq61/gI4uUrwY6phNiSy7BWNRhihsTv3vMZExOuH7Geu7GzwjvP
N+IskOlkREw1jFLTAHqkYQpB8LEJtCFig3GTewydBp7sPe1b/9zGMYCzb2VQvyL6
UgvLLfvdOVeqR2BrGiPIv09vKL8ZtCifsd4t3wDrOdMZyoNlT6l2dXQ7CRlcjIPa
EumrCE8CndT6orQaHXUztBAeQCQgqUViyFY/j2ZVCEr1irlWZR+llM/jFEUd5+28
DTtGuHQT5qcZc6vSD+lnMvOR4DM0n3j+DpnaIi5il97OQh1rtciW4qkLee5II05+
s+Hf2qJ87Zm52vc1HG2iH5Jhh/7+S1oSKKAMNIoCOBhTuQ7cRFMWYErRmcxoyeex
J+VGjq1ecXovmnwWjYDWaTPuL028YgHUkwEHzMNKN/YEA0Jx1w7EscP9NFHjBrY8
Tt4yDhQuqdTZogUOit3V8RIaYp47Y0xgd782qPgy/m3pYg50YD+x0JJuCDSkRzDl
FG6SOeK04qroRjx15XD3fDgjX1ag1vUhHWs9wgUnjDiVI3r/Jbxb7a7aqGOXTPlS
dzboCzs2U+z4wZJ901U0PEZoW/OGqJz8WsTk93XHshlfqJsuezMubj8m/Q6VH6JM
ELSE6I9OPH0cV77+3Df/VDMTRv72bSyT0MEbpzqxz4bgvsSKXRclanLYhs5iETxv
bxoMnQ69Fx+Yf45gp+tp0pGXr1TrKUy8WW1oSgkvglmPp/urThLyB0liUSuqaU4d
oPdJ1LM9Z0wqTGAg3oPTxtqjemcvfOZiSpihXmKW3vxBe0pJQ9W8ytQu3bNG+hFy
h5IDPtLqAarKdtlKVYCvDyGK+3YmkG3n9ACX5xWDHGjuvKgObIqlGy0S091kJKAR
nThRXYXBb0fw8MBgR7FkOJjhfOykntNNzb/szdvtXbVGzneoSGEKE6D37DNYVCQ7
Vz0mI2ZqgBmif2rI+5UwtSC7l5nK6pawRUkS10/RqP/jT7M8ppDUk22T+Zl7EdWK
St7pSqV14FRmI+NG3XUswUaVRD8ODd+I0BAs9+jNRPagEIPUGdbHlOfYAXeDl/lV
r1bHJ++byyL50Dr0EpbpfayxRtjjrReiAaqta4zUAYlWue9Ze8ZbdPs6UBcg24v+
Kr2HZoenZ0m7q9nqBo+uTyjjdd9WiBhJlKeSsOb44tYyNUxyVcepzVNbooFkGkRA
0Gl1R/3LlY5ZQamqB93zQj7gxXymQg2LeyXuwSaUv3uPEx4PS+pKvN49NYK2alTq
OHBuZSVXuiMEVkhfbdqTSYMsMQUhS/mMlnT+4Mfsfxb+RIROXZkG51phnNeUmZeu
lq74/awZVDnkeFRwGv+zs8wOCVVYeYY6MxICyqc64x8OlGVmibZTgg8vip9l8wbr
hs4AAdScqm8PSXSRMpKMl8K4t1fTzyX0+fGmz9bQeruAmXkSuvo75zyzGHUcQlIs
cnMCt17zI4+qHDECZ1BQ/lUETWTxcJAS+yum7bl/4bYEO83c4Y6KJSx4FVuLCK5B
NdpYeaFvPFw3eMoSsfaE+7EZNfXUg0M+wdIihm7rtbrgy9O62Td80cDkZcXvWoaW
2yOHzx3VmmkAG/73LHwlqPyA0V91USF5ZdX1NiflE0ME8JJPwYL5nfu3WegZycPf
akvbkKEfcme6LUD89hC/cbZMe+nD5eaqHCvcCENo5AeqlrPsmmg2GKoy8dwPPiRV
5lYa/OUiSwpvEUnq/s9MbZae+Xv0zc38+0H4p+DOfpEAfLNU/apNW4cnva22l0c7
Lie3vdKSwmDuH6QNpGxRMfPB8NH0nlMlhLwSB12eA/TdiUi8/b/UIt8G2YCK475g
g5Le517aglh4A/a20I/BZkE8LX3rL9HO2u/88aTHot7ye0NJYxIBoAR8gz1B2vhu
BxCZ8WYJrGIvznZLswFj2qT2vRdR7iKd2c5iEomu/tcBw0nR1u+wUkdYwaPiFUiP
2hv4zJQMtgIJqwYhuFZDidYHYQ1lHUfqaM1FNKYFRUAyuwFbFCiCJbhU2C1BXqVa
sbZhKj5La+X/yztQjMpdXOVzxNr1L6F5McRviJVaZUq1tSqb0JrPy4P0RAZLtLU8
0zZMPSUS9OPyw/xHP7Yd6ovRdLRb+sxB0WbuxXu1jICoJ2Ss4gsekkcQGdGRDZJh
+JHDFBG4S7j/QwR9uwvTOm/L8O5PWYwlL4BcjRervyUti4Pn4Ji6/enp9s6dOnOO
3qBHM8sM4ku5gIT3HXFlWoX7qXV+S4M39COAR4dvOKUkEWShI7ScZX8mNXGuIAB0
mcbH4mZBQXs6sx5IKZVyL2iI7iSWa/BYtPTXicIoN2DtCF3bRw3uawvjBCFdOW98
Z8t/7cjo2ze9mrX9MnJLqcsA0nLAO3ZfDsksLWxRWcDvoFr6TwRJzpxD0pyZEUv5
axFjq0p3DsJ1P0VN2r6E2+oymbwJDz5TucXX4CwLdG+zffoN9Jc6sKELDDQ4ekVK
hdRSeTGmqimkk4EXdLZEp8RUUmjzyZFDca1OeHJxozcsPryV21mVL+GoeOaMqjrg
bZSyYprbJPiWhnv7SfDgDp90rwAYhz3wA8BSDw9zcXZn34hBTWJxOBMNfATHVDoe
oUtbUyf4K8sEvWbMNkmK11y+nLuG2jVZwaJZz/9xiXRGGo5KNUnRt/LZ8vUG5ey7
t3JjAhb1JQx/6wOtuPSM+WtQdgb1oxMp3u6LtPdb1ZHun3guerxEsuJ7/1DYefYe
yhdBFlVZnPHyN64OXwb/7P53l6zdyl7E31QpenT4L2qqKjQ1C2a4LLIhdJZpM1nl
s+YT4FGl/WcMhmKmXuNTZ15fzgl2JuzaBgJj5pvoizqFLABk+eDM7BKyng8HzR9T
igINZui7FN71ZBvLTyZahBJD6LOAG/0Uc504PsqlUbC80QAu0iD22bKBnHvvNTLb
RcQs1ESRwj6/c2Ar8oSeo7kceOLXgqjs1449kJKvuCcKiWjKaXs/bYajObwyZfEz
0MB0j6JSBNntXUo3XH6NQ64AsG+/fzB8/9Sf3EGd8PvhLU3hFhfvv+lr+5MrcG0/
gz+OfDRRdmfWtT35u/H6RrZ9BCVodxjDGysqnF3yJKM0cwSKY4khQ/E0aWcd+7Tu
fMylf8LDLkopOLy8qDxLqzrcm76J1DRv0s+Z2+yEMAR8pT0KJaaB9ZSIKey0pGPP
BsgKgPX18ncdO0T225VfJ+SR5t8kYENBRJhI27XWhwrD1YYuGJAlzIrU7WwO5h1Q
hIDnSwTbqKxFz9uu+18MOxB4/PO28KNNeADk6zvufSBlFOXsdMsTPZdYXrxvOTNs
KTKqYOwEkV0sPuAwKe/wG4r1mm3GjJAqvcE0DW6j1hY099qbTt0fyDvfCGblm4qM
lSA09gQYchT/8s4brWscMn9ZpErzSnILch+S9P4yEzZaiYTstP2T4gNd58fXN6eS
ayHdoh4zcjkA1ukxoibiM/3PLyMQGrAQvUb9m6hsU6/qHDch2YjxR0CfeO4MQ0dP
5fLx/Hje2DmYHnQ60ik0sKbV++qPZyFTdWfnLQGJJ09EGJ2OvhzstU4OizvJDHY8
6rrTigtAnEsRDZWcEbGmvtd7LlyXHTl+n6kEMShaY419/18V/6NmQyJRzLQ0IgK9
v3hkqB2Y7qOnnMsiKg5roy86+BbsnR2xM3qPbcAR2jORtdX0Rbt9SCZS4fizE11q
PtA9liS3dd94+Tn1bRmdqFp03qsaUidv/VHRscT+7npfaXHdQlz6+A16/mX7Tr5D
QvJDMatdoou5DcwbMaAjmQDbP1Od7RpB0oa/GkhEPkVIXS2eUqwGQSSEbaVGTskT
tY85DCl7di3tcfNAsaGo1t4u9o7bFbqCSj0CjyxJihWjJc7klBNsZTKtIUhE7uoe
8rZKTLwxp6hJDdI85hwb2lAlsam57vVEkTuplNNbC+A7llXmQhjXRl5Aheyqs0gh
xM9iZzgcDBuBY4yrAFzxXJ5ENP63HItzcl6S/PLGpviWMFLbyw+W+AMAbKx5SoVH
g7LOCiW0Y3CLCm4mBy8tJVRFJvZg4QANo2HQLK5YUYPNUJPCxvbjZVBPDL40nOXb
a2KH6pSa3LSU+k+YddjLxSQe2WiprohtLCDypPoq0SHjOXNcVqpToDGDH9LTROX6
0RqClSMZz1Ik/TOOIjefNc30nLO7Y4ZrA3a2qQDPoyJo31db0M8BgmDbw2d16o3Q
0ck3D92kpfX990TyFXFkr7HtqJMtjhtaNOx6Tuwi8gZU4E6XV6Um+YdlDs4+LF6l
cR3s3ZFJsZSTGfAZ3X7hTK0nUSLO2GRyfySSeRSeMMf2qCQY4UmcE3pN3fZFvS+H
AP+IKWEzZAtG91bHgfKfx7hA708Z3JoZ/FgiwWDLx8spjQYcHbkFsNDy6LNDAbCd
e+pCPJAhxhS/9aMwftKlxE8seB+iA5MeF2KLQ9LSi7YBhVUnCcbv93HaTOBKR3xZ
MRQAC/1jC0KxbMr5ewIMkeAl9I/yMsj0oRIMq/4QsERcx7mcbt3aPqYbz3gm7Dv2
1ZgM7acMsmqijUd2eVvYvGlnNCZxv6Y0Z7ZjQm40LOGhgd2OiuOYcnWZ6pqw4EQz
/FeDuXX7XJv7BZ+I0RSp4z5WYUDFqiyGH2OU5jVwwB4r/mTYXn/08pZiJFZlZV12
uPzveV+9WK7UJnO9X9j9KivSjJCnXvW7yGCzXbtTmWs9sdXtTJJMW2mrl9dBQEBE
Ue04+zJz5p9y+jwiligyr9kaXiT85H369F4DZr21MA8XcvzmU4Zw/ui0KhiOd5cx
gfLjlEkXk0WULnHgUbUE5hIZjQQOEsBubde3RG3OhsdFrfqdiw5zpRSK2aiDVvas
/xjU5L5P0jiMjbjmvRa9hoCRZG+lfLwQGhtpx/CiTbRwK1tcvKYLY1B4nBy6nW3/
JFk2D34Z+bF8STryMvylMPwR5Mr7hSS0MLrBThmL3r0xxGy3MaK6jd/8gkBK34Fn
oLVKC1QC5tHWsif7DPt0TUavmbzbiWZ5uAXyBrM3+TtEPUAdn1OTUXRYoi9132Oh
rxCQSBJopssl9tn/RtzGF2eMKrIBQonTTy+2Bq3UtK8jAUOW+AW5NjK7rFohhv0q
AdKXdlgHs2DP194J5WBkRpO4aAEIZ0zEcId4QJVWMYQGM/qJ4IfHkzKF3vKz20Du
3kPVA33wR0z6HkU5v7wk9uU9GHrdKbxA/qNu019xnJbN2pXGJsiF+d3gCpov4NRR
hAvYQ6WKElSy3XOSpiTjgEPlowHvsidZrHw+y6WJoUWYKzy/Q1UuKgaGVCgNiczj
OpdQK7Icp+IhXNopxeTvjMyduQ+oKqZYArwv1yuyTqcO19NWOurvgEj3UbQuSURL
pgdMDqUDgXdPB6XTbgn9Eu/TAQnlnKoHGK/cqAI+Kn1p4SotSew2K6eARRFris1u
rxslAvcvykEq6YM5Ve+izZia81S3TIxDFSbp2XGUV0MQOBBnDBgfdvPYhG5CEDHK
hrCk3/MWgK9YS/pnBqEy0Pk9Ofyo7fS7Qg9JwQfWewyKhdnzH+DQCX2lUFAq7cAK
IekkQTB6PR972YJbu80eMZOcy8EUjTNVA79kgIoS2SnwYZxGy8Pe7sXc9ruj7YMV
ZNi/c4G8Xtbv3SQC0BTq9Eltc4nATrUbLKnvc0UL89phjnbxYh3+5XR60tYHGCvk
GDLq0B08XkQW/24w4KN8u6eTBIfFHK48ZysdKi4aMijLuI3OECze1ijSpmmZVapA
bmqJ3Irj6EyWvkBc/yoHZQpCDXzSXd3iHfFHPDbTaRbYY7zV1M8HnPl/2rgRDZP2
DOvKnS+Jw0den2h+FfCJ4MbNREbWENOeMx/OPYDPdZVvbTyWfhO4ZPWLAQAUsC25
upcDrqoJsTf6tiB8TdTi/3plFvd+gyw6weP9XxunWisGwdbV6Dch2liVXBUsqfR1
xTDdjpbucteDcTbwEtdUo6yulJqXfURkWn/xHcT7ILkHk+d5o8Cw1im2hCBV7aW3
bu1/9fiMzhT8ofxJJ68P7rnPpQDxvy93U1orlwWwq4NmIWhxEvGygU4q4NNsDD70
nYV8AkBuuXFko8AqAInxxr01JeTJmlZk9MPyMOofYohtpgNPg0kCz9pIyEmKHyMP
KMV30q9VN+tZUlKylzfufEotImcVFMdMYDOoNN6656LY5UegNqtO6pqnFmip8l3C
wptk1jO45TfLCA/XjiMEuw/nGPp6GNhCAemWcpTBtD3QhPo2hFrJckaUj2p6sMkF
p+kUCUYvhEjpRPRd4y0r372+upZyEaiGkDUmg6pSqvA7LBJBnXmEcyCm4yKx/zJZ
Qc4VpHh3UOmjiBXqRKuc7ysz4n0eRDDfCdXbJq3Hxr/aofWwncz5pfBO5zRxA6RG
Z4xfUcIkjLpAhtBi4ml9aPokrIz/dmMmMriy6ths+jrKZnlZfUWuBkq/1F8CfkmQ
iJZHRyRM0/tZf95J94Edfhs9Nf51+bhN8mEevvMp4svawjxkHAa5wN5hDaXgIv7U
dDE08ajqQNAIKnreiBNsuDPjPOi4wl0jwLmZyDZN265K32g6HdbWwwIyXeTlEJja
Xm8eGWi7HHDDEtaUuRSclr0lcLQVXKXzPla0pPy6LGkKFvUzjrYcTM9fPVuF/wn4
fb4gplDsMnkHdBpB6PXNNFuKmhpBjan/VOdPrjO5rMSFOmINGSBoMWvpnzQX/eHw
mT6QU6iPoHmpNjrAixvB0gGwwVX9dnkj7voQHhYto3kAljUU0Ak0l0im88G0R+T5
3Kf4AR26fu6qVV4JTRD/RJYZc4yww4/UBx0lNUYKbYSPO4L8X6gvee6ZjaJ9Vwlz
q0+VtNlh2lKfY5tM1aCQSk4pvRoG7Kpwq3t1/4ty4PCgmz1xTpt15+86rbxe4VPJ
lMSikIOHL86NIyTkDzdX9SGuK4RdWUQsyA8Lyce6u2z6RYPRXgDNquVkJIMq86np
fTGPfLbkVPmB8z6dZc54TgX1BZiFD8ifjkq9uxuGyCwRs7ux8c7XTDviJNFK3KrM
DeQK5CXP8JY7nxXgKccSBIqmHVNM3kT/tqp0GFUp9sF91P09BQ2NeUyiwTae090S
zXEzsdLDEzlysu71FB7L/7soPrtNZEsG0+M0nSQ/RPNeYV5aWMko45Dk3DYbnv7S
zzVgrSkzUxDKbDcfK6lXlPXtLeKL2q4Hq1GZEY3BBYYi07uqvYu+VNo3Rwm6jap+
yE/nJIMVyXL5dsr6yHoAZdOUCeV+lxjyN82PWM4gtWkJn6bX4Hf0+AOOsXHu7usZ
ztj0ayowPN2nSRmYP+5CUpv8x5wlMzQxCCfc8X/z0UoGPiEW20uvbCHM/K0LZLGw
e0TbxvIUxSOuzCxRisThoTs4yZpYtUUoLBY5f6bymoOcvJpUBxbd3viqutoeXLkY
AOuWu0hrLPhb089IcAHTaaqyzZCYChJ5IhUd1JiSsEGWBNYdCLVL73m4liOydXTe
K6bTzoJ/cxWwSVvyRcLUi97nrOS5r5VEjqq6OaHgnjJi185iVZPfszVwczomR6AJ
12EiCSkKJLpzsLzLN/Hd+CsZTRwfRhEf7/po0M6OA431yKG7dKz74/0W9D+Ab6dK
uR1d8b8a2xhGLcpkypfPThV0gaxv02EIvKpyCtYrv1k/O9M7igBwHUwabwxJm6zz
wgaLWpnDj2XLduEs3JLnrHnbyrgoTBEt/ScucnrGF5cMBbOat/OnPjadZFoDiex9
5+URe4PsB+QKP2nkDJ6YD25UaETLnqmlvhtaqjhQX4YzDiQEDvYnJJzEg+Ba0Hti
tyqJPXRw+pR7Vgf3bNr1ONSZitPLm1RI+5XF5ea4GxrkPk4Q4sF6GVTxQUEUPh8/
rvB50RYiowHS/90g6YJvJwKNzE2gnAZpO2jxsDlskQHr/VA5a3o/qNFxUTkE34kD
WO1xAvNIS/nDTctOv4jBIusl8pLXTUmbb5QgCQpRWfq7bcZWveYzcHh40gYZyht6
eCN477cIA4r966eaS0kbh8LFWMWjJexXe9HL6d0JR7FpdT15ty5lNndlur99L/Ic
JpDj7TCbhEzM8tAbPO/TvTv0QP3X++A+216CwyaXOPa3B2PtgpH1X3kzqfZgOgQ/
60D8edv0yLYCr8Y7zokB4lYfxUFFwz06vXMC0ZTh+r5tBKFDUwr51Q64zG1mMHU8
rnim32wMCONClF4FKiZHmA/5iGKjnDGvj4NIQZDVX9DxdoGkqUK1xfmDSWKDPTip
/lF9rl/tjy2Tpxe1vbFJy07PUgCBtsuTtLfHrbubT7MjRchNfBRcCyqYCXPxPXV6
xEMuvBL9IwbN/n/Uxu31odAU7FpR3Qy8ACiA/XtTlLCfiCCMhmQAysk/L8ZxnMfO
JGhstljWqlfE91kZt23xnF6zBFkZ5n/CFnl+lRDgC2RF6HFbvMCyxJmwFYbVYsSI
j4yWvSkuVoYUUORl0d8yT8jgqbXUbHocBGI2SlbB5lQbRwSpeuqX5/pI7eRAQyQq
if6PdGxJLlrooq1MZVNiMJD4E4Nfmf6KpzVTj+nE0qaWcdGmvFRSEDWfsGkL895E
TbVRjMeuphLXLc/ZoJBrtJZsvV68684ZEExI7KqzBhfTBI16zDbHnu0zgaCM7Xly
+bMoQO6c/3hPvBlhv5LjbNfn5AAfFRidPcq8gpztNfpQaZnKfMnwS6cviMNOYqBc
2P4UtV1tScjMK+jT2VfYvggfYInM4SQ4jrBpvuY8O4RJx+mz0MPZ9rcv/2Mh01OD
ILTnP9jIUPi9o0ZPLFgnt3TTcMS8+VaVKkYRzSnUImDmMpKeCOkZQrf3NfctyxIq
62NZ9HmjhnfZGO6fbWbqO20EQif6VY6Hu/Rpggz5JQifujRp6OIdTtEY6WmarLk4
AE880L17USSOFsGFCaXxEYsKfP07ujK/faE+CC2OPQ8+FY6YmXupO5u29iIMIQeI
h16HtZc0nyYxIk+/oLtvDlfGxcvAwskFJWimIAYiYYHO3vLoma7dNV4LoKR1xdt+
UD2zLeTVbJJAgI5gK+hYjzmoSHDx/jUeLqBxzs4a0EtY1a9v1FQn1Y28A9mZvsc8
8Rhsmkk4NFhWHoed68fl46KUdU7KHnVxvdtGa1985a5UXwgBci//m1U0+MN4anyQ
To6hFP8Rh9pfqfAZHDKRniJ5t36L2Jr/cpaweAsmhCJSQvrT4GW6Vx1JYNA4Crpk
RJVDI2rjNaWqrIaCUovB5E26/qgQZed9AwiZXhmGOUZAN8Qwiaxp3KwJAc0t0N6f
WmiSr0dufMgGi3g4scQjHFaFwMiJKuiw3znzJJwTxX8wxJeQJWsCvpiTKBaOtkiF
paWlb5q23ypq4QnW2Y+bk7w2pTrAzKkdA5YekAkgEMOHpvVacaKt/ZyEP4wO5Vcv
j/3M6PpW6YXVut5r5zaXwArAu6MBz9hTXImRdoWQx7iHM1r5ZcmdPN/RDPeaDpJP
MH5BgeETMjt7hBJwVq1lPWcDIOYf9NA4Bqav9Uw8f1aVTQ1vo8KOq4lexcA7gCL5
X1WAxK93+bqjX2ikU/vEvkD5+COGAElBGtYMVyE3/959FN5a+QdxVhRuQvWZwNCU
xOa3X2haG/aP3/1n9eVUhTEZmw2RpSvnncz8Jr3EjbeYC9XxroVV6ZehUYqW2Tgs
SjEkfnkjeZ6ePX8IhmhXRwmJLhusHVFSpFThgYgeJXwVts8VWUiO+3AOMLHvTdXa
nZPlvMk7PLlnoQ9rqkJvUiRfTKOvVv7a6uG4W2TUuQYnCpZr81C+iwt+5HbkDIjx
MCZR9XFAS8CUpwqGE9FAuBVMKOt+xbvdPV0S3iopKiqLQ5vHp+jdQD72bcVsr4tG
qqJILlR5wlAXpf+1RYl0Kvl9pZC3oyuPQyJI2gcjHGHkQcvJ10AEpKhlzD3Rsc46
phSGswBQeweJaCMwq9tl4phf51mk2wiKqWTBjyBUSI2RfIzFwzzlHMN6D8Yv25LH
zQw2fi6oPnJ9WVNYGKHGH6e02ZZgErTGa59IZp+6xVbYiGwLIYHouoy0oWJ+Ei8D
S7pjuZAeyqoK58FJQc7U4kPWuIx4B2LPvxaBSuDAzHeovZ7TNw5aLcVGzTxUUoXx
t7wG0InEruOAr9ksL0jtTYBsVocX0c2UhNEt/a7NTvqxF3vfqgwhw1K10C+2THPO
k+cHh9XJiB751HlOy6UdUFEIaELQ9Jrh3wfM4cTDLoWviqeT0su/JBVJlQ38F1qm
EZ0sc4YSXamjwRmB5MjfRLJcPdCM2XvR7d1TICBN3SXVct65jXZbvNLFyVl4oTAA
8uEsxF5TBbHvd37GCGsZPYJJSSz2osYBNSTaatrwNlIuJkkqT4ALibzuBkNPG18e
+HasyORWKcPMGLMCMusn4DQfO9KEOkygsGikNFTFdai8eSMf41kKF/Nwp1oKq28h
7fkr4QLH4FpmGFzD6xmZ5KDejOv6rqdxqQaF1QnOdetaBnfJZkGLuq+/3204+xm7
cK2zQ9lSgTi95nvL0Fkfkwd28qItXmNlWduqleKXhA+LBDF7pd7WueQk6n0C3IqD
R3RKieGqy0nELG07nGATcToKWCGxlr9EUvb4zzC3EeNFQz6Pv6kxkkvtzWMbYhby
5S5iKsg8nsCss7gpHbPbOqrhLRz5TN9ETLR6a85yvmRIrzN+Cnu6uFw1jKGPrmLd
ouOGphZIKajRqwP1y8UrJK/QUG6fyA8fjRp6QcFSTF4bfYFm8dVLBe6qZW77C86u
LsM79ZWJCqtbU14dIDahUoC+XRhBFcsA2rllvs5SW4D8FmKdXKnki7GJuCcywTd5
DXoIB4za6RNFcdfgaGZAuxTjkGmMNDoqOcO3Ov2XLyDgqmI1tfE4JMpKGgiBOArv
PCjYwMDkl1oAa8USaaSksaukv1GnFohOOlFg7jYtXAIrNmz27h10b1tbQ/ZaWBKK
eaUQv/HWZc5KprARLPxfzY5CI/9OXbQvl9QYThB7ik9MWrNZb+q3lgjc/H/XmSF7
EAd3K5BBsgzSAU1xM/1znh4urJYRVo8NQ1JyxpBuRCo4Wsca0vtgpBJyNnNtQeSO
aNv+K1hB7y5vhvMMAzyEY9JctIJNKjUK3fxstX+90f0mpJvT5xzE6sAD4ekcC3bq
3YIb0TrYr5SVjB7tsOjCiknz+6IwbcBecyU5HKsilNI+PxK2mTWG1EIR+nQIpM2B
HK7mttikGhxRQ3mbIwq2bmud9cDHrImU+whFh9ASreSe+TKfGrL5fu0ybrwHARvZ
BbTk04J9P383eDWM8RUFJeQfe/Ey44Kvap1ZSRFnysxa2jDqFUSVkKrLL286Zwse
IV5jvGHHQ1afOt0pdzlQSUSOocKRpF8kF2yr2nPH6Q5oHz7WncbneXLyjerfDkBc
pZ/8P9yN4F3A+NwCzOvyztjqoBkL7LARDBUF7YaeVUlEz0eQFFkJLQIgBDgChRBH
nt8YY82tpcogWnSRgZ8cZxBTTUIBr4BHhdK0Vks8NGjZ4gSkgf/cQmheUAPUsI1X
AjPBx7uR+kZZqcSlwPRaEiND7FIozTOD71tZSQcPv5WoB8Ldl4w7fuPpkbvdRmc7
4nrO7i4yNQOgLRriwAiJqECWSAWfVmaLJvR4oUucS5rZdUqSN1lLb2m5Gxl5WjbD
Wz2DoDt6rkfHBqTzQzF5yfU1xL5/H/mY1QaJSWCtCJg4Hd2QJPmKREpBqfGuLuXI
BAuCeL1oTq7lVKcjWwvFiwETiiTB9TjRz8/GJU7IU6KR5599GX88VgSedK/3bMDT
Ws8cxx3aKgNT9lt3hyE22NKauO4tRpwnQy5xiTk9Nsl5aN/nDD5L4IMf40jzlO4d
PSqxLju5cH9ZLyzUBquOgQ8wE7jz/m6IS9l3p/3pPRguaL4S53d7C3+eewR5SviI
7xEV3JPsHHw/kQExUcKZBmlzEdYglT8L0mgrxmDl1HGitxVt2QQKk46LKQTEj1fg
7VLD0qAy7LelO2b1lBb0IbGi4aiVEhf/QeN+kuDqkJgQbpBhxsxUz0bcFPbLv8A0
mKA0NtJT4srO11aJlDv/kdEQTy9QVx4Gz6zhj9PEI8ssR7kh3eNuqZWpLVa/KEmb
Pr5ofkqoC0SZgj96LBnjJDgYtuUGndn2vYMEVFQC1q0rR6vXIHdr3f/yhaaFu7bp
zE17/9/DTj/6ex/IJjFRCTjp9yoF3JUZj4LcUuW6HypeelNMBK5llY9ZOZ1LZldY
DJbApJ9BV/IEzZ1fovn77xkUV5jy0H9El4KE2GevqFmDgkwxASJlRAsZcEUmz5se
1gGQbaPNxFJZ4hbt53BuEt5h9K6P6TROffi4edrBbAnWNVOwT4fP47MNhJsS28gG
TDwaA+06CSfJ6xWy5QNkKuBhDp9ZciIaMB+vHSP3/bhoe7+XOcxWzqUvm2Wm7NtG
fKK+W45R0Q0JG5CadtHSihftQvmruRyFRISZSRqbDbkvjMaZAuHrihYK9nuN6WgJ
+Evrqc0GEkf6jC3k87jtOG8bAznu3cFqXIOn/li8v6BZg/5UhThZJur4Ww9U2BTP
OPIgvTRwtwgo8YGD3dmcuVh+Lm9DzfZhZpGQb1oyBDSCiZ2rDXzZFWjailSsEMS/
tiit6BYnACciScMZSg4S9GTP4MBtKTGg/LUpfdsXSUO9fH55ABDQhZSy0ef+RdnR
wGPLCIbnnAjR8tGp4chF0wBHXC6gO9vHQvghyW3q8tsVxbSji7Fcx9NEpxDNaQkm
koq02J198vj/5gTDuMc9VQs7pe0UfOeeN9XyXNruNkk+71rEiR1N3pPPPL2rqgqA
zDQQjya+ON3XpL/jGP/0fsrcEopKnonGWrrh+LbsLKgWbwjbaPcKlEh1q72ti1TO
22WzlWnRog17mNyry0imZLQaBZ2ZnlcsWh24HnQOmPLeQS61Nk2vWcflb+PnnoPZ
2PqLDqWBKcIUJuCUoAX6w+q3Co47MGrJx7NhKuQpTFK9roUzLOeYlu6QPYbR/U9V
iIOh00ObzsTA9N9qgbQKO2IRXBJSI5Dy8b5Yjl9lfkEZqadBFG0yGpfG47ueNYHS
e4FaTwUqvEX+Q3k8YpIG5hw5DYuNcCoEvQwYxxT3LUQEoYn0E62bUIy6tNUAVs79
a9cKyYjDIkqIIPIh3mn39RdldwR2/WwHdyC6Xsjq4kHQOf9YFjVkfrE4BZrE68cX
Nr+uCtXGqSacEGJQSBWq1yR+BKaVUM05sUYGipvFi7QhP90a69riLWT0djFKsNd/
4lAoDl4TdkvxBczb26HDY42hCSwjr4ZBGs1L7TEvfAEYtiiql1VZ8f4TQ/WXVvjW
VGQMhh53JjVgwxaGNZy24Ek5sWh8W+VvZ8TQwj5+SYjVqOOuKBHuLYah5FZeXCiL
4EG66W30lNmDhyLL+9uqAUHY0LhFzLvUIzrEz/yvq2cycqMnwe9oUj/24Wjroaiz
guuz0MlNnlPdFEu42ahrP6zb2PskrsnbQLA3Nu5vipuhHyRrl73f9F4p7+geep7a
F81St57qwncgLzIKNcZewIgFeJrbw1hWnTGRb8oTzvm6cNrZ7/xb5MrnKM4kg1wy
nQLFCVnrfaCD4jlWZfDnMd8GbXUu7esYy3/vud7CR+eSExee1G2P8l+iImh5iNFJ
VAnP/PI5kBik89nErcK9LnQKFmtll3+j6J+6CbM94abLEgg+N9J0jrxb18y8aP2j
21ZFe1qUm4Yq8CNk2lo5RTssLS3fbD9rUn0tfIY6TlM8+T+QvC6NSsAx8547ui4Y
FTdRAxp794ED4OCmsjx+CoV5dOOT4DMMxuKqIh24M/sPdCP0eG6ADDMbtGS721h8
lPzgG2okyUole44YpLAGT3xrbwqjNcNFketeDJetG9vAZL38vvKWsteSxpktQz5X
ML6xwmuzJ89Fd+WVmbIF2Lv9eW5z17KkVqymGQvcpl7l+KazTGIhyUVk1AxUUU4Y
1/FYiSogdapMU4X7asp+OfhU+z+KuobER1mIxFhz+R8UhDgGzQhFRNjL7LVzyeWi
EpAdYD7abL87hl6JKNy69YeX2ELKsFKkSRauRJLLLxtneOUtz5yHlOuUnb06BKW0
fasIvBjpM0jpPWk4JWdwRVoif7rpkOkp/6a2aHPHRfhQrwgkho9m/pHkwKlLAG7n
Qep3R+IvQkO3Ttx8r//Nd8CwAUn72hPmwZm+utTNjjTYEd6xv1XnZW0FGAOdSckG
xO3L2OdExL1D9a9wTOZtYcTR4tQeLN2r1LSw3VQPvJSVzdOfWX6xmuGXXSii+usU
xM9g9fiD6JguS38k2av/qFbWrf3dbydevceAUWJHLJsJ7Aidqcqdl30fBuo/4Zz2
gZQZ4Ct+qd/E6GuUlis/WiECIjYdiEGpJLbrwOeYIEudOWm3z7qUFQCMDpFslUKG
3G0YQYOZHlJa3SUhyCJtcFJump24wJ5egNfoQCM4BNeyYq5wXLsApNuoUb+E28Kh
BprLGh0bWCQW7MsunlvJfuinKBliB1DjhJBKbpRKpUXP7Nx3/AtKfqeJTnuZpvQe
BAMH8UNnh033MtB3HseMkB7o4MnJwbkKKxkm4tEoFgB+ZH2ctzsU+Z2E70foFa5O
9XGcAzRDt/UUtb947JJQDj0qVU3f8UODYC8Uhh0cF6exphPcKKVq6H1kHr7sEMxN
m3z2K5IwJsa9c9lLMlzGM8IeUPges9DQMilrrDm3tf9xQnRTCKV6UzExqF074o0q
qzXJ11FhmwJjzZ7M39IoZL+HP7B0kWVzaj6vLOIjmrfmiJODmR4XuvbaVMVg3wMR
waEWmBtVEUoIwmZbv79Uyf42T+zNlZmgaS0QVTJwzSblYqsFC8C22B5IKu9VUwDz
cPp1UW1TEzI3eOMxDvmYZhm/GhB8MpNg6sUEi7CCiNaadTc/xprxyiRElLin9bjf
pPZWe8T76n2UFy5bxzpBA8tgkgWkNKv1VWbhQPil/rRfoyxTweubW/AOLuOr+bD7
0gx5kRLsxOlRSvwmfzAjfo3Y0p57tN6FGoiZaUxJwPga5959yUU4O4QmCwENVFXp
5ZTsJR47CDiECzhx1FXlWwQT0Vuq5IJe2NEcJTFDYaieDmeEXSwsSbvDpMxCyC2X
mCJwsK8mB7DX51p3/RCQd+Di+BiiQjFGtsYRrXapvgdojpmuKGseQt8Hi0pWV8G0
0c/e1Ua3FvDppzpB6vGzr+J3CW/yLO0bdCTUrSsc7zUhijXy5pXhLk90S8TSg3pA
RR+Gwjf9RXCK3vGGVHKjbfez49zqiLXEJvbVlNS67Z4dvzMevh9GTX2E3aapwRj/
Li0nR5ZGI6M0IwQDMuVs32GigXfa1+wMa8dnCAB2tjUBsOiHEpfSr2ze2FUscfO9
ll0bVOTF7IZgLFznlP7YnedIV8ej4nDbKK0HotnhRCwFWN/Yct4ocDjHFzRg1MP/
4/EsgjrCVjsu/J0oHS3X7byBr6wjoURlacGs6JNFj1sxuV01XufdVgjeQGg/N3dh
bZPo2h3NbJ9k/0HuWU6yqZh5PEsQ2kOETX64vsZ2lxzd1VJOJnWqWADxVSlHLbA3
XDjm6IiE0UwNEJAepoEe31Vj9drgvHlkzWC+3aV+dSS5oRndtS6uMh6eEXh1V4dq
q4fCG1eRUmdgbSu7MNFOtaHV3CNb8nElyUjYKEzMXyoakYZaC2goSaHGvSeevhVs
VI/ULUiCksZ143GJR08Av1Gmq6UiN0VV/2L5zdmem7s96ywgjNiek8+oeURNUGD1
KZn2j0Vv0mrPjfLs8Go+E9EwlVoglRxok2ULAR3myuRahBLku7SgK+/aauSrjuEH
GYi/gVpw6BEodG9lwf93YfisKjKUR7oG5aoYiPpOG+kf4A+mIHsqNFO9XWZFyOxw
fjvx1kUY+CjFMd/v2X+OdHoAoB2hSyOoTIZg12M6Q5SMTv1Vl4VzeRWf4hhcG5a1
dqMOxhL336JzicH3oexpKIJQM5YlijxT1sD3//uFvpVR1FTfTZPgVrG8X/76+UTC
VKW+5r3QfvIPUpodGJtTTrZ+aM84YT7IBDFkDkRG+o0gBLmnVUgVkeptYTSTZ/OA
7te/P/Hrjd2epAgGbgnIVyKab9szA1+PrDig1X5Mn1ankM8ZFAb7AwMcE4hHD8FZ
4wlUMzyU7oKRr0Borhuydfqi4J+fyCJRjZN76uSg6TVDpo8G4flIx3pJ/mueXwEu
RylppR43KCLUBKZ+xCDY0YozMRqBV1N5BFfIENdudomXkifXJiwFVAhiRiqMhq0e
R3N+1JgR0adqht/GX9VM0Y2GejG+cpWtx0Hu6u7+gkXscp8J+3IwKTMbsmxFHWlC
kO6+XPgAsy/h5JhJcGEHjTPhlUZWa+s8DCh/6gnslHjDURXzAZGO+39F6RQtqm43
if3KhEQJzX983V9+R0nrENKVJyiwJOT23FR6qF1DQZj2D+bGx9kiZe5HSM/B+Jde
mvcudorXLo20QJ4o60mToXTYgs3gLxfrkvUhzoZSchEx6QVWq6WPxsiFl8MqsOw4
45ftPHL8NP4kM17gBevk9fDMEJ2lSilIhSlcNYHYJKoHiJPBXcv0cmHwLnHLpLsy
7Ql2rGk/elO2VwgkEDRpojtBGaoKGvb9dh4T8HGBUHPpePcOXESul9o/y9akkwAE
zbkoI9apiy5SRRxsQANvVTK+IN/ZkMvAQiDbzDY+VfPWdedi6tt/YBgtuwCa5peR
Q8Q0sbo0yZCa11NfdigZytVKlpw6KjpNLdg9mzk/mFNMG1VWfNmepEW5FXbo7gTG
/3yGWdGplPI3hihM4bfd55Cndmdh9eNlF5t7AvFRYD4faK/Lz0bvr3rG/3vxcgp8
/cpiBYsnve8T2dNWzVBcO0ybRYI1oIL8vpjUuA8teeUhGh6hgYVYMWta+KKLPnQq
vKsOMoKJWrWr9YQsfpZlPKRO4ix08Vy8Py4CYSmBEx5yVqHQgCuKk7Jo4xGAxnq9
MbiQdg0n+1PbiOs/2fVZxwQ5MsbeafAkdP1O9/uBYeH+W0GJTibWniWXbkKxmvHX
4DBqYLw71CH++w4N+Vhg/cuLfOkruSB9FkqsM1NCbsN6HU6y1L63qqqTcqEQ+Pr3
EuYcZ53DDdBVrE9dlLXRMN7AUFo6+hkmlDuLpT9beNGklzv0g2fZzH2gBS/wyMMa
u2U81Di//Af7UCoChEklvDrYEbOf5lNFkIMZ42LlMFsDntsKzhADhhdH7/2sgxUs
Ly/YAasdgddWKa84l8pGEJbiaRTQMXnNWSE3yE2SaZ+aUr8f6rjg84njraR5lXBA
g9j0GrRBX9Jz3Qm4h/6XaR25XxhpuYXn8R8U1TryFpkwklIFe3qHEo+Z7xW5kYAI
ek9fkEIdFWPMieRbpRFO9FEKVic4vH2qoatTDfekJEdaGMpY3f6YN0JQfov6Z4aE
EKIBRMWZZJqspVBVqOkyufgWpd4OYQ7Ubq2jULxe+y1sTCrpmID+NlCSuvxgFnvU
Wjnm+4cSMOYTZfpzmexzgfo06YF964vBUyObaueQT/nn94xl6o9kXoAL58U2kfE8
/Xh52thysH82coC3LyNoopU4caIJ5Xq0hQlou48RVQLQY5TDnF6NhIqjmIeUHI2L
M706dsJeXtMrVVieZcggUm7UJ4/udkYU+g9x28g4nezC6WDQ+z7JeoA1LYMtMlZh
EuZmY48b8zLe/c9ZtcmK2947EfeBeTCSwqVseuiF+z2l2Q1yZ+Mpqkuvw/L8Q1jG
PIae/rgc9t5qxhtvykYY0d5hheFOzEDywFMGpguVF3nB2pqgocF7o8nUVKGvuVTC
lUjvkLan7uj4r0d8vAr1mk2Dtj/J/tJ8tw2xyboSJ1QnrzLJpN2qsaIPltKlULt1
qaLaIga76cSMBEK0+mzb73XsIHD6XT4LZuCw/89knvd5BJad3bscG9YT2GNPYKd1
rdH2VKUWBOdENcP9/1XikohqEjE153MqGtsr17Q6tVfx6LTJ5VjwKKIoa6yqFFJv
a8Mvlp+9ClPQvCPha4f6+H86KRVrarVPtMzUz5Njt2nTc2Hy+W0ymgbBo7IUMQ3d
z6svKkr640Z21CiRR8Th0AAuVmEomPZ1l0aN5tZOgKvZZlJ1UfYFKh470QQv6VKk
xTtyhlY6wuCH4RTQjqqJK7wSvi1TShJ8Gjq4HUraQKbmuFEB/12T9b7nyI4hclQs
H6Tp/kYOs7jXucXOEiK1gZ0SaoH4sdjWLntdZNHlhokrw14+JyXBU/E50BQrxtIt
Nc4Lt9irVNVbJMHzulo2dTsPN475xhvdJnAQVxumg/KqCVa/+eIyoOiYQL9p0AcL
KaZ507bHr9K4gdPTdVfOnlYgNE70cMedYZQNSO7az4McKIQ8EvNiTbbA5usLNDeP
Lr8TtO57RRSg94GWEr6H9LP4F3/9n2Uux6XsJ2C/sG5EEwV7sP9NyLGgLhrjUPKF
6hlXKpBiJ8GMb8p2hkQwHfUfF6atPhNX/5mDUgY7MlD28dcO05hI1ZXk8TKosHcp
3FBdoFY/PE1+V2amWdk5/SW6fIJ1Oy3RSAsH6ETjmUm4ZT2J9oDN6aMNphGDPhaI
+oMYiuZXu3qnAaNe2y4jxWzyTfdHeBgt2CW9jSu9zKXcl4bU7Air58VPek1RUMuQ
3JS3UuP9BnnEljlRcoVzI/d0JQYVitI1xl2AJTLA+4eUt3E2/7bN2SmYRCWQZQyE
FhqrBaT+hbTQa2oWC1BxBHJvcpbXwUoCB6DAmQ+vcASOPSbfCN1j6J2ciQHptgmg
5+wkJ7ooAE+u4toZy3lSqI+IaVwfBwvbkdkyPv4sQ5i3cYRX+jpWmxwfaJ0F0kgG
CvRg2nZ23nstWKRIqCE2Ffv7i9uoIxoqkZcYOpoXrqqEyADwhW+p24cp/3/b/4mO
YgRTa7eEg3DulCW5SZC6XryU3sTLPAVXyzvVHdQg34nXNnRtVobjE0SAwSo2LzLT
gd0zMiVKK8+uE9Nd7cvghwPf8h0DT1/FRksHXLkrpANMi53yVIqBIOizSin7aQp7
MkrbDiWz839+dawb2H91DmXKmZrDrl3Ui/NYmO9JslCP0CQ9DAxce1T5rjCN4oLI
o+4h7UVX727oVw6KzL58FY/htGz12xwuXcPQLEQYrJ0zKJsG+mBhkz94ns2NOIeG
Wamm45kGitTgCePZZMq7BozPpEepFA3PG4UjLjO/mwjDC1VDldH9J0SPirjryj3K
1UKGNzn0sQsVRf8ryXS5X0AQ+lNV3pTAWfp+ocwxV5GVCqd+8u+tuKDxrT+aDbXA
B4dClRkt6uqgzhJ0OXBCXlKLiHG4dEUNo7mwf5n0ocbF1KbK8ZwjhEV3YxRndk1q
bsfG0nfLEeXUh8BhJnnTGu/va2fDF9kliEr/ssBDZ9Ah2mk12BDLrJINLh9XAOME
BlZDArvBm6AoQE30bSyGd7ISVwwhrE6JU8QZZm1/eXT+WN+PmlvrjuvBoKT6psum
LEnCeIHORfU/hl8aUdgISZyuyc0o/QBUMsMiKmeIwIyWjCZhO8mxvHO8AF5ZxLu5
pyM5WTf5FIRode7d48XmKRLuMlWOcz+JacIUXLXIaE3Qhhjy1FAViO5IkcZvhn6h
EK+7xnwaYyl8r8jXlR8eSfXNt5sSPL8Jykd5z5Y/DojNUOVxmZNR25RF6b7cS3ak
IPUiGzdnBnYv2InkcQmmwcNYrIkt8cK9sikIKwXthStnWtg5yzX1KwrRn0yEY0AL
sa++16mv0eSZ18Zc5GgsfvHe8AGKZaB52ehFN7Ldg1io1oVrUsO23FlOnQlTgDlw
t0c7BQIwFaT4vfdvneknBsVo8O0v9BjViLvFvTtC280+rQcNTKdecZFhVGbZBX2i
N/euSygxKChupHkrTr/f+7L3fcUintnQE8FNwI2KTSFF83m86ouIm/TbdftINDTp
kMKV8xL0ZAvEjjv1GnJ5rS+qIthHwxgDeXGGHl44c2r5UIGRP9ctBe/zweeQ3Cbp
BeLgSy+n8hi5rISjRD88LeuwQ7Dana5+tWZXBtgVHH4+rvRuMukYlSMAgEmU7U4H
5uKD55sB2ePpjD+Lm2qcCEzxjKe1MvBx8mR/qGsJkL6l1ylT+qvAralVvIIixced
6Xsk3uM2TRT/NqDltqOFFlWa1UEA6Sdzq9SEvejBbFnAH+eJwynUQ7uWz86GRuO7
KnKMJXBhxFsfMxanFWeFJZ+bbaD1DJwt5PlpAPji/C8HLg9XIvsln/fMVsVYHzvA
Qgdod2QxXABTLw4oi/F3X3wIOxl+LqKfh6udHJORMEAzT1C3rNMXH/8P5eCwa9i0
lBVw06nCeyKaiRGj6nLKto5/len0uqh3+2YxABii2zEV1hR/a/xjP43gdB0EiD2p
kFbGpha7kMT66xFDETjxMpocECu0rQ1gMqCbs7XdhXMGNcP4RflVU4x5h1X8VOEo
lsBHrPOTvMPqax0BSb6w7ANvo2lsukAdC3YyVuJp5+p8dTyeg+Qsj7f9UpsYYQPS
sEkiWxZQ/FRYuTsyfIc8FsAdvyy0vkhDoakU87a+ytnBl4DI60r/1iOdAuaCpNnI
Zp4bYl6CBrETMbkLT0q68EwO1G7kCQVlCDt9yzsSIhD8PktGZmzoqAUh0WqAvKXF
shteZHgESSDJvlLyU1PK+SfsFKLKzpBuPNA+2GqzQhaZC9/hi6wQGcUO9t7rj+x+
NGGORRN8wx6gBWYoBaI0enMmE6lkFIWMWea/2lKPruKAVraVNstQaJuuHMCS9bLg
b7smDlyo+mCSt20KgbRwRpa9QJE1KITrtnXwDI78oomu5WCmQ/qttVukTR5ev622
x5UeTuOJXbctmcAbqfH43W52wD+U1ipwu6807pFg9ymzcCKOWlaN+gyS0plW0j32
KPa0tg1LIuXUH6QFr46OYNmdmXRZS7UMa8Bqf9la2kfeLYsZQ+RzUq32SEgdRiBf
+RFsXauuUpgv18v6PTKxGQfzmLFtO72ZNiReC2/GM5RCKHdzUC8Mxr4BbpuBh7Zs
WOI45HASWbiqCGa/baXn5etVwZTE5J0lqPitfwmXuS4uqzcPqdREPQEhvXyVmL9t
dX2jy5ESGaL3M/HcdN28jlDHL3kt2riTpm26n58Cy8QgEjxk/KzLi5h86EPS+8Qz
kG6Rn8n4B52THYcr7JFLEHU7CMLSGCctY3B19e+WYzd80X2uJTdPjDIXoq/TBo1i
slp7eOU2aQSsjWWRVu9xTUsAV/UrsA5WpE8mQ3MHz1sSOCuWiwzKqRWLkFL4tKa4
y6ZFoNV16cRe7ILDxHrAKVZujaa/LoMx89ZosPhPra1i6qaJWSMePNX377H1Yf9t
I9C671htLcA6S/n8u3OQ/ypoC2qfzfvTZvAyUcv/ytTMDj0gcaP0SdB6B2OqgWUw
StP6cOb4uvDlEPe8B/hcieAWM0XxB1AdZf4lP0jFLEhUFN5khX1fOu9bqLAYwrQ2
krezw93o4hgIWrck2NjOIfSn0bvQv/fLElGP6mvcmHQ2i/nQQe3ZW8tKkhP3Dhhc
0XQg3of4+UX9pECmIgtXNGjehd9AyFLnUNFVXTd/pArtNx1dcVSlDKxeakdo+s9V
M/DIPgV/gkkWxDVK3Am5pn1YkSK90Pys9Ryz+rNV6oFLaWZ70QvzPmDBb76OElFK
8UfEainAPvwnA5K60kXkOpA4o0Bk9bIUwhFcMGgsrkYh0mC51DJ8G0qn1VCB8rj0
pAyu3cqHUCmHCbgbrI/mowfCmE1S7cm43V7MbdPkJz9Ih+gcVCsXUAp33xdvRVc3
3G89G6SLfk9ZmtjAj+Ecdg8zE5EMP1mDgkCYOC07TfBGWTThuuWDnmlsNi49uB5q
B+01dpoFJv8ttgXoQauWS3vMjUnWu0U8oyuUFUj5fmM7/vcN1ZfdzWtqTzoQGM1m
Mai2wRzKzq7nIaVMEYtLc5YBPqNiEbaEidkjtNZkeFfKYI9lRLghp45Eiuer3mDX
FNpaCXZ7NyDc9Jog2SkkZl63TibmtgsKi6TYkr1dNMzJdKqSThM+PUfWa1ORI8Ma
WXDIqvjCOI3NW8LmJZppBmR3eLA/2ivi/fFWpAolIDsyyxiX0zaE7B1JM9KJGGbd
XQ6gdyA1Q36Sdso6mFxZ2YYriJX3qFJRt6s456mmvOO1Q0co1uiK7PKX4VITGGJI
Q1mL1IxbHtqiFEN+hTqZ06XpR+X2p12g0zbyJG4w1RfPNYz72ETeZyT9YzlXRKhK
lkl9bhEgXxCnf/d4nBgZMQTv8Umga1Ha1jBF8KquIGuZNeXaOTr4AdGyWR4M9KTs
kOFIxWZk8BHxQrnzm9CXyz7NnpDRzii3+R5287FzdEUnq2+xUCEYIrBAcxfTPe2J
Sa3pk6uOKUuCV0wfSiZ4lqMMRS21he6lZv7crOujozdr6e0kXNg5pj+wS8Er+zKS
0+yO7X7jg8DCuq/6gbAf2i99kE5Yf+VEME8pF+pqZ65ZAuaLDhYwCoKpcxvA2e3I
ropmOboO9KoUVtQBeIEpdh4IPVw+aiv/sUAH72oiyZ+4ec6dZkls5kyf9PglA69L
9yAI7B9MULtcoE0Eoum/1/tUjocyGRWh58BQPuwtcDz3CpkKIuCgjt3hpKs0Gfpk
BjiABoIEikQITFkb1UKcZAomVdQgsvrDrXlpOsDsxVrboAejSnJn+WDFQeFZpzq2
XYlKTSMT/1/gbZ4jA3JIcxsN0DHCgf+u5lzfIJiTp+EKqcTPjjLGAIy11Lmrlnap
V0ORVsMOo6DmUpuBDaEt1Dl+lgGE7j/Urq8zPByMm5NL7tm1vRhlAkBqbzf46cds
qhRPRgdtOB2jPSDdDi1bCsI1FvSBgdI+uN49CFmR1XX8IB1KGIis27cO2lsMjY4J
JAZMPyg1UXgT+6Bix90pxjUwJl+rKaT/G37IvYemi8uwdmhJeaX+CebDfIIW/KTf
hAWZowxdPHymCk2LpCinjwFHSSS6teeDUxmMQ+mTQBP1g5boX4rEvNAPzf9U92qW
eg4zFqhuJKGvxUk5q8k8f3qF8M7aHmfbWSEdl9oh1/oNYF4u5/5XrqasT1vKqULz
YBkqCX+thvjejlGY7v84+7nvMoQ9A1X0TnOlD6aFXrDY99jhkHxnhQJtcHh1IdaN
6/NDYiw97SmRNOYm6dPm8lhWZzN1352is+7ZFjYgh8in7bceqEb6flnF0h9RxbyT
lU5lyx6kNTZwP7mkvJT3Db/dn6tg35TARn7safBAqIGxLBEc6Xt7GVYmkoKZ4YaZ
JU+RA2SqL797o2V1Mp2eS/7QJxkCvW2L2zDpQLKkrez9MQAF9fNzkdRDAjIWGHr6
O+zi41UfVkftjugLSwnqR02FPiA4YFT834XaYASFjSgrPsPSfbDnqIs//GsXX+Dl
F0HVUR19iVvWj0u8w6sergCN0g04dSb6YMHoL5x7teJA/Cb0v9EehOc254BWVNb+
2aQ6AgOPKk5kBO0KcGrplz9q9h9qw05RJr9xrvmFrdqzi414dCj0n/5HBJ/fzGtR
MKgPrQ/NoG7TYK3bLywBQXC6ZvZsruLg6cwqLTWmwdyHF74zngtF88MRqw7B7MLN
L4g4XfH8Jbbc59e514dESy6fQBftULjXyV3AlaCQ+NF9B3/PsW4bWUJ+9p/QYteA
R4rnu7wek6v9SQQujXZs6rJ+9Rc1ITBasGTDib0VS2XLZRpZrZCejCl/CD4rVd4L
Y71PTp/oExWGhsDuL4C2LY/tnvavm21ltlYIV+3qBkBpjqIaIjCbQEpp0dvrGJ7m
YwepQkHULUl3/vyyrCecnaR3bPDHNfPrjoxQAcpQCtjc5oShS+Ari1wWDjpxxKX9
bxxvPRrs4W2XChXDsNt4hWiiX1wgkkQ+BlJb/RrtRyZmGjSF580H1BwEaHmaSv6S
awarPSE+mRDq9eiymf2gUSDEx0+bo3JFuUAYun/bSjoOl2EiQ6FnssODZnTggQTb
oOKvVg/3VoyJfLfmCMy3O6d1LHIC9zyUxbVkoso9NMsOQgjcAbcktBIgmu1AA/T7
oeiCKZchiCAOTzYCX4TmuEYVOTo9o38N7ad30wuvjIf70rscOxqAco0FZ8/EvFxm
OebcpecLBALV+mTy3BFPzDfphVJesVSitIAon1rgPw2/60VuecigzZdgTlu3jW3G
JOajXcmp/9wGYEW6f8GW8/5eH9F5KeByeW2dja6TyCSG97AknVYGMpV0Eae+DDSM
gGfAtWkRdFUDrjj+YmwQkKixX7vE6+izkZbrk7J7/tuK/ZVLdVp4Jk5pVg5U+klD
zfWxeTlKq6mm6ExeezUo13FKuMzo0VN1HZSQ0HIlyCn6cJ447s6rzVbcYmtF6B+4
q4yu2lfnjmjpZ6Zo/ZnRnwPi6EJs0RjcxGhJ0BDbXfn2qGCfJP7yisa3x8avbptO
CI8/AKk0p1wXLoqNQfImEGg/bi9DfRnHbEQJGbgRjThHtbfVJkO2if9eiutAK6mh
kHskLNPkcEZ8wxSkJQXqxzUkv3m1hqWVshBGeGJYW+jJE4vAH6prtxSJWws7XcuQ
DukXwQWSbRPmPfHRhXf6GzRetrwACOTHdsW6LbK9Rg3B2UNibE1Legs6+INfr4zn
XGvuKeMGYzJg1QMAY3sqd8P/MyHZDOAUL2cLlgHCMK6fNrqzs4ujJaQpngyZtmVP
FrTakP4imJjP55SJrBV7F+9LQ+6y/OLvJTmHleWicSpHByhZB5I25MRS8rJ8OB47
tTKWVplYJk+wnRCyNZkcNWbWvnSlcT8VzIqEjB+gvc9NOxu7E0odm1iOjvnyV+Xk
oVkzaUrXKvV9dky23AC51AnVvOqw/rd76iTPgRqtScgDAzNingqZJk4QWfJWxMb7
mZucqEvV9qfFuT4C1ipwdKQzDxyng/80SuRNZV9/BISKb3oQ3cu2bopb1o/g/fG0
lluQSRwGOb6ISZCeKTRRNTWW25VWB5/HGlcmDNWEVX+OJvS7FvLKADEK+/vpV6tD
retOQmtpDOUG2PE1A8KNuX9d/lTTpDcNWtyaraATEfpvTXOCm5dBNpILjYUI2lTm
CCv5wK3BX3VBuF9UHTbzpWeXmnSzuzPY8xVd3U+I2pOAL8yMd9J8jGX9MJjLtd4H
52gNQmVNM0mCQw1SuGPdRgxNkW5Pm4lYEbWXG7xKOvPLIgEMMFhX5naMIoaOBcQy
kj//89huM/wQ3ahJPzNhlYWESjug1zhnvbtLjlCAApydYWXPIhpbYsxyomz5lGHX
tT8Z7ztpJJcsrLLGOSKs3CoPyc+6MZk0M5heMQyl0lrPoxIQOqeqvVzqFgC7tEUq
lYce3oFn99QP8r8/sEROZA2VTnlPW2EqEr5+9J/ZwVsN1pSdqkDsxwM20k5WiSKj
bQNv+rNfXeiBPmR6P2ClihM+8Gq8FBHxQSYM/5r9eGTA/VtddaVd4NHjJ3t0hb3W
tRQRymmpkWRKS6P/uVlnhQFaBAdHFqrgcFXVma3yd84kduJt1Z6dI9+PbnkH1foX
pePD4+Tk6e2kXX3BBw2wyXhN8dOrivxZPWd4sWXPGGj+sjBonZ6cxbf3WY5wLFPL
IpQlwW/Mb/zE5Pwsid4PrKF6+b9MzZZ3FW/GPGHLsamflnpJ7ae7JSas6U6CfN06
ezugXWEOEg5uHk9wGVuoA5VS4kQ68y3b31Cpi7N1HVtpaCXdV5/KuQXShi89w+AP
JKTqHg8kSVFJXHAsgCFiLMwO2QucefyNDL1nA3FG5aE86FZVohRvHhc2VUzikeVt
phU4cRY6DEHfbMTUKZ/vrIef78xgxv9cYzo9gXODfXI6O/pKVazDgi/UVtKDCCrZ
GtWxsZ1q7i9R2MUc+RGb/5j/7UPRFfeR99+0ZDqiPrqaFzzTWu+D4ZNqJyr5nYYu
qHnQirsHclrv/qez+LUr37oUpte18XJxs7sA1DPjZcbC3f9FoHpWP+6v9eLXyXvK
ogSUpgPxPlk6TdtXMSenZncezR0MMdNrDRYRgLyPrK/8MuT8jmhClgR/73EzOjEE
s8m3k2MHwBuO4vptuj2GpSxz4HtIRVe37U8E1SsXGr9N9jYpUcWbraEXmPFqXlNo
ru2wKz5nasdZMAdn1kACjsglJ8WAA/ME08U8y1ZzTXT0S634Wy4yyjBf9Lb3Ehbg
EGhZlCOE7nYk1xGP7DJ8+pEheDTfzWumLaKoeDh0QM28Wi4d25Ck+hD7KsXmQtVG
x4NjeW3ApU2myUqqFXXnVc7lR2gHsV0MpUHdRriZLRm6Rlb0y1bI3MnSRF29RwUs
23bkF0nHYpP9uCfhbso35sQZozVbELGjdOD3z+xsRG8KlF9tPINiFY/HTFPlHGMy
UJ9zRO31Xssb54UFPe/84hV7clceIcXruAh5uk7CsSHioEBjVCLuZcSrM1i7p6Zc
5ic5TCV/Dh843fEXjbmHZjdG4sJZK6UuECXG4N9fxG3ivfebeJPlzvXA9EZKnzDD
cC0Ywl7lc3NqEaBKLeQO3xOln1ADK6IWZ5paTAdKwb3SxMM/d1wg4ijJ77mfxN5r
Wun7vhB2gr3wDHKW0+Av0EgNXJSzGSO4txbBS54twkdeqqktvVNWSIKRAytIdwme
AJBDg9oiYrFk++SldlPDqMJUF+GgxmLraoEHGlcZuEr6C9PSERUl7xsCirct6rFw
coNhqy4v2220eDvEo0No1WlgFryk1DKztIjkh1wfx+5+DuCtdR6J+LVpasyXyMKK
snWHO9fhaJCG+ztztQk0alLSE6qwMS+vF5n7zCX4i2TyZ4/P6GPJdfNAkqnugfd0
ZDBfjsdujKJQVDc0gPJXTbC6ilxiO1gOds4ojXfHRM+rAmiZxH/KNOo6VUPHg7zr
5plwyoUSZccOQuvW5yGzmZny8eD++cpMpgkRw0eqOAsKpNZacSxtRmVA8i1NlJnV
AYxevviDU+EKgt60LU4ED6mladhV5rz1ZWUH4g8ssMGdVlU9fqo6yBRgBkd5FxMU
5Pd8u8APCeoE5mH9yd/EChhY0yao8B0g/ND4lt9TysN4BSxll3UA7/lkvThk80D2
ZRjL9vNpvrQil7/IUMQ1eQbTdFawhvJ2Uka2uvIFqkNOgvnUV44KLY88NEeT3nO/
+nAh5szBv7SAuST5QpbK8Zxn6NIGNCLHx580H5Jzr0okyghE4GCUMZuxbGG1UVje
wz3tW1mcs9Q1B7sQiGnwLkxRZlHNhziRZHxot4/QTw7lCLa6HKQhwc5HHbqAVrZE
ZhFqqUKfSWRQpxydCW1gkLyLu8upoVC3CO6KboiFyauEB3EPs8hmSTajJi7CT9wG
bfhEYJsl+t695lxuWeCx0dfr6QYAGwjfPPB61RJntiGthcbYTeoAPTw3vw5vppuh
orpnQ+PL/mDyIx/e4EvVUFRC1wbPBYr9IIDJ0TeXC2k2o/caqXKivbZ34Iz2hxNn
5CQwYhvA9LoKPN1qFUejY4AxaPKFrzSX0LyFReYfdq/+G1e7WbqWu3BMOq+2Vl4s
yuLVBxSupmEHGYVHUqFUzQaAPMszLMHPF6GLsbS+4r7yV8hhAOQpt2JwiC6ncA49
P2xrXdVJlj83qktJKmrvDGtCRsketTiM9N7oGTcc6dRIuGtXmGUUk2ZdzmP9hg1q
cAiL71S1wzING56BgJ+cgQz9IIBy/eQ3ra/DX6/2e1yKSv/aLKyqAb8EHpkzgmgt
cCZOfirGrpldZ6nDa0VKsIDR9qUOU4c7EAefS/kJsx+uloEjN8S9PnXxnecYE7wF
XI/kjpakuAMgU5vvPQYip59oepBbbR76H17Pj7JBX/5jnVzYeQaY/qIFySwTFELh
nhXpM/wnm0tFmOx1q/O9aRABMCwOu4lQaS23xUlNt+Y0GR9OH4Mz0ovEOmer+3Pj
5uwCfuT6TOrO1H5GUVde6zY3vm5u5huyvcXDORNtInvnX6qeaJpIZsFPrV5WncnY
J6GYrtrGSerN19Hq2iVOfI5AptZWpuEKTfwvSwB0Ib3NsHROgCxsHqrWcUCBPgr+
brpm2yeBumiTlYxaF+Xa4sawiUZJ86aTpttbqwDpiZecArfDcfYHBVu61FpCdP2D
gvlbxW7ggU8dS44rM5Df7I23a6CQmI3bIG2op18D8OgQBrwpUvocwwfslLk5zuae
46TcZDiIvMMmcMzL62A8aNne1OybSCyW3eB2gFD2KwaC6JBP/fDHlyOqntHUT2xj
O7UGAUK2+s8MTor/J6r8u8Ndwf1yWP8aQzr4oaj5I8ocW6s999egsT7EvWwuIc2h
8P7wU+1iNA8PgA4Qv9kBpbuw4BqUfFtAmNjF4t0wH1KpLR5u7tgvsHS0Yl3p9K2x
bx7lkGOBR2HJtzbx0sMUmgRLkKfeRJXuhOYKvgBp5mg4zuIBPKgVaMJiFHmSfJGs
m640WPy5t8yKy4MOajKlUwkEEPNvhYXTCvZNKKrwoJr7JbFPlqMkDZ5n9oa6VY7B
9GW0JRTsHH1KQzGQLqwiWJxQOgquj/2hUmBEJnN+1/5VWPX9a2rG1d/edKXESKhh
TLoMzSOfxTUNJJ90HtbF9Xdg3Yb5chvF8Wzwr1ECXacveeskmgQ5TnodyX3vnuUu
k90u+sRaMImnyEIxTM3SHSLFByyvfYjdBYRNshrPcWtbMZeWyrKVSHr5p6EI9dbz
mltlaMJPqv+EOH5vVPvtS8UzyqG6nMLJyLcjWPcM1gGPvUp16ZuG9S3VO8ucQQbB
QVohTcIgI6x8Y1AtamdOcPGet1d4gTpcLTbub1iZCu1nH8SwtjhSuHKzQS92lLY5
TQ/gZHDF7aWVA91J7bcbsuSg7HQoqY1Em2DyESF9UcJhIiERw480V/Tteqq09joX
eNwYBtBfJN7DRCBkgWaa5HgzQQ+myD2CotzhbWi3FzPd31MNoh3Em6iQJeS+csrd
+CzIenLbWq3NJQKL4KtycKG1LkzBmhL4rypUFKyycHb0zQVLlk/c6j/vcuVccP1C
ns5OMwrVaH7IUrFVHnikfkGIR1JC6j0s/iJL+bD+G2bPzRaaD5/PBPbEDQVq4+km
MFQ/EvIUKyxMnEVHqq4OUzsSad8GXjTcLoy6poS83mFyubF/KTffe0TWGkOxEGhh
PAhP+KZvfEd0ik/Yg6/ZeBRVaCq90V08ektHQZjqPx0Jou+MXwBIG32LfUFJI9Ez
62+ux/buubuLmxGzN3GlRR8D7aEcLe5PS0gY9x19oJI9MLBZv7/IkKwWo7nsV2eb
bPyT+/O82QtxHArx1kkwxGg416vYG7TKxXcNL6XBXdCbwbikpr3JkGt1JlSTndDs
KAYbmotWLM3h1sjlyCYzMPO8Enjxg75yi6m5X1l3dmTI5FuVi/iududGtHUnuqLw
TPsJmMkIjVx+rB/lyBdR2h8opH2TYTH6TacxzLu018TG0fsjmpuViAtv9teVb35j
NlY2s3d5+VvUFOwfJZjnvn5Yz/aWXgXlaQMzrQbgCRy25x+HHTJBfqFbgGabovxo
QtY7X5RvigQh2XHDY54/oCr5bP5PMouzUpXbSCkAfSkbXdYYBb+oa4S4wi6A+5g9
k/LlLbiAZaKewwov0xc0S+k1YesC6q+s6uibPlleHD8jQkrj2fPAj6f9wV+J0rfu
lwUswcqSs0bfXCc+rS7RjNKhC7f0/FMMJC2xrsx0JTZ/h3/gUKDANz7nZ9J3Lg4L
Ygxwbl/9kDjPIxbnyxr3pBeeU6XLMbO5xw0fJiLSUbuDMIY4RDPJHFzlhtrRFjDb
/7UBbSydi7y8761Daybelx+xpWiSoUXlpnVMnBLypm6luKjx7OfXzlPZOAakSEfV
fmoNp7peYJIIzw7a7KW+PI7ip0fFGZ3ohmC1QwJBl/JdC7mJaITsdFqcVQSrhPBx
Hns370aMNNSPXf8Xf9RTo2trXJIzHztC9aXNGeh9dUA84igj18sgzZO2O9jPW4T+
/fGOkQDwvOlUcmAAxo8tJs4BHl85ODDuMhn5M+5qr9wQniJpaQ12xrhjs6hr3Pyg
I5dNFkRARakRBRgUDmhhsq9wtBiDi2f4FlfipqGgyfRxdacpyCz5Gfxi/wA6rLbd
/1vK9VR7XLA2LxsPpanv6yWjpqrUBGIN4Yw1me4vRoZrHu//wV7LWrOqhGGlyhVf
t9nTR/AB5qrsQOLjbcQ+n+JYxCayh3PEuxkO0qQWOsTUDP7TKmj5ZAlOJXPuie2X
P24BDrLxQboaZ6Vxklf8hV0aRT0YD3hx3isMpk8WtsjLZyNrZL5vW5aqapjzHLT/
JiOAEW2mqF2fZgDgPp0Ay8ScjZcwZ+4iTMpBaPwlKQbZHQJocnbEn48jwZ0YkzSp
KLzj+qajIcOgov1xIRfNvrxkkdV1+0I1i3nuQ7iUQmjLDyPNJjKfrUh5ulWv9mhi
G5AGcsYm7h33hgt4U00JIZgTQY4fVmpnjP58dRE0p90RFxf2M3/95VPZlQS++9de
AN4+EudbvTUVHFDbi+ktmtn+ChR5bD5EQDz0Ws867YhXUt9O1dRGeo8AkXHSCspL
RufXXNsgHnmze4snNyf8fuSOoGezdodfxYmrJ5l7ElJAzfe133idGBr6VZPUCXej
+ERowWUZKLdde6YZ0BvonAfL7InuOPNWzK2+26XE0kdKnKq5f41yPiJc8aPINxtA
7Mw+9Mu2ZIixQOOEcWhd1PemlS/CUTOiLaVtARMAKzoQNirVtFuKFY1ck3YuDeRF
PUjAMd1gJ7Nnj1nE6Tm9gwrsfIpc6NIHK08OOP9bgRmbd+46xy58mQ/MZ5uFIxdH
guUbuAneNTPjfjNixoa7KTCesDvQ0SI8BpHAcCsWxD2o4NqaeBNiWN308xoluhgk
8U23/aTkIAesxzMDxPJitY3nEomp9M/s90uaNs6CJenqiFN3DellL10wfIBQitCV
SZHHSyttKxA6zDhxxWVcDJpYWLSpVhmtb1F3XI3Jc7e8jmSYCpoLVRT3u+7p122R
lHFFPtplz9/ddFPMwyqKlM8yAE/lsc5zOw6jTQ9ZvhLnJReoICilmRnKYcZ8Cahl
+aCTXVCrDyk6lk6e6/Qw44R/QCwCrPQiuRD35I7sC2IBaQJvCq+8HjWfVsOCbD0b
gBaYLlsfro7Ojb0Y+yR6KXbmDwLary3HRoWHey348wj3sFAi0KWvHnjBZ0wz6IaM
jE/CpTRmaRqUe2qgg6ZKPc64cjRXCGhyvhtUfM5bayJcnk6AMMBim4dY9FTuj4n7
h0ZW1CbJNU2UE8EbMjSShMtKLFLdDux8Km5GIwzw0N9w1RkUF0yztk7Ls8cGzujJ
z12mB1CjO/XNAX5dMfpzM0VZd2+Xjb/VS75ub/Qb2L9zvTwaoIpb8RPbEXNAoXlC
0l8sgB5ydAW1emA3V+lJwMhxmbVRj8/6EXOn8lxJSzXwc8ENAKMwluxO9rv60dMH
ViC1hEmbFBpRZVNlrWeyxJJb1O+i/mMTqEMUZY01gCTbJ2GKndAJTLiEtmP5c6Ab
j8kY5KpWYYnIx6o1Cptf5eDereL6xcDI+HHYBZFDs5uVOMhqQ2+W48hN/JRW32C6
XLdrt6G04Lu/N33SSWauvBmS88UezmDRZNa7kvXUACuXxp8WBd2sIgC8T1re026o
jH/57MJGMfpPzDdAK+3heizE/K1XON6+nCZjNwQxAMNpqg70tprue0GzGmIrPGUo
jW2m6KClDn7m8Owogv3WPITo5NCUaHDrJbz3BwJ6yZJeHipFJ7/tdaj8u3C0tAd+
TceAiT4CPxT140seL6oe0Q+P311gzQ+zxUiwkUPb3cES/6Q593GsqQPv2cYajUDY
oGIhxotDb97pRnW4VX6F4uROXcLrSEUwqsikLB4sbCQsyo8zN8VcvgAm/Lys0Mhg
ELVX9v1iokc/XUP3E6VG5PKhK0Ei3G9PZd2+SZ5AThtRe/dic+jy9zVJzBWPephc
ZPywWmDspMPi5Nq05aI7inrLDOL6AfSn2EEBvqv1+D2IWY0+NUrJnKPr2K0oSpce
d9RPKcEyDgozWWT5KRq3hCCZ3QaLKrJ4tfZdWF3ldaTbDhCwhtp3xDMwn1xj4NjE
mafE6OS6Nm6LZFEiciZtgYjoDGXSniDHn2k41iOe0nvT+MRUWgz21M8gyGqeu52M
wI1185SZrryiliH0yToX0UY9wIhuc5m73vROJ8foo15NgDIeswF5c9rGJqQsrrun
28HD7dx8H7zE0dnXeRstShtUJyGt6tEB2yJo/IAl3kIKwPAaKA+qBPhIPlK3tb0b
nOyZh/UkXHYPMc8rQuVUPmNvDgJg+n0LrQxyIXPRZeRcVdheQ53AzdPcGKnIkn7Y
Dw4kmgpCxgee2qm64YEjIJPT9u1UyTPmWcMt/zjv+HlmIYLqqrNcQabIJsgjcojj
CsIIRX9/rbZdEY70lromJkMf1gHtbunZVpfylxFDB3GkGjkTA5XeYaFpxm94vJ8S
NvR3zr9YoaS9ahE6y/u7UUJxCOEEMmCGa+9Kwsd6C/vTvCEtgI6oeGvXMpfpGbZ7
Ek/BtIuqjgxXAqdAJK08Rg==
`protect END_PROTECTED
