`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1iq51e9s3f9T4gjOSSuAQlYzs/6Ke5uhHoFrwJjZGIQNc8wJXV4iZU6fvkU8ZwcH
pUrzbe6A3z/z8N0bcJ/jirrMQtQEw5kARFC5VXrLaQtx+XFYewRxmKKYIDcDlb6a
C5fVE9Xz78Zc9oFP9kqpcx8H5aqdXm+GyS1/JPjC7kmOuIuq6a8jgT51eXraaxGg
6YG9ywUjOzmbuisOHslCqmpPzeBcBalayAYboNAS8ccjdoQ9YWAxl6nsft/DrlNO
`protect END_PROTECTED
