`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zrCvWg9Fh61xbh/krFk5XTWb//h2g4wEMbYH/zhz2QJ21h1Bc1SY3aw2MedIu7Ep
J2y1Lql8OL39g1oNXYhbbt7IbPzEW38SqnPUDCikP+JweFE+7btcNCmCJg1bYins
y7tTR/n6iP8kAkiZTJWRujpaoAhdEUrn0I433UUyHyB+F5vvwb9JKL/fRwBSOFlH
C/hibC+rHK8sPBjYHkbYDXnhhU8PWDF+hs28ma7CmTBMI5EK2oHtQmc+36luQOMy
ZH5zxIx5dNJM7L2I2ifbVPGXrqWO4w/4MOJHfdsYR+VZDaawlcEd5/L2B5ZY7Zuz
UWzum4FZ49OutLEWtMEMCa9Fl3SfPIWthCOn+/BSlyKa7s9/wYqgFKBjvWcM40wX
Yj2aWHjC9yW9XLEXWS8wFGmh3iahImTR3flibhXveO4HOOI8jx8VgX/x+K0bmaQn
DZr7JIVaO7s80dSptLpNQZ6kne+hZQSxqg4Oszb/umxW4oZobmCAuBONK1AIO9xs
f0as0R3gHCHMPAZAqbj9oQ==
`protect END_PROTECTED
