`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72qW6NmauREWKwNcYoLRoWgqAkEuEbiW7CRFo1P+oHZdiZiqQK2ZSa9fWf/3nNNd
nDlfBTNvMyb+ufZCUY70C04qErY2UHWDZSeouvOMiRzwXYapmzH4kz52mZiPFKpt
JOW8ONUUyp27zzQcNyzBwtaOfNHwixmKgXPWeDKcS/q0ehKK5F4TxH+DTUzFO/lW
/74IE0L3QDceEZbj7vyMMgRRYbqsLZwxdnhrJSlSMKd6Zvau47zjWYgm4TXuXdHm
E6sXGMBPLd2gxSljf41WSBUk2xSTc92Sd9m4UZ+kbbtK51W7QLV6SoAwIQoUy2m9
DJIcMIOPMwFkpACMYFw43mDSuxaUwPkTwL3K7abghpLt/FY4ipSniXMLuZnfWb10
EZLfZJwfCXeVYLbPqzqSgTs+Ip4aT6rpCp7cnPNOOUrc0ZLvW7Gsp978i8gD/l+0
dw73+YBPud48qsugJJlzt5bZevAUPoGuOX81Erg/W5nCsbM5hgzJYi2742pF2LBR
xUlMG1T4xDPzBuoNErrl/4VR5lKavC/9TcMgFV3EdIPR84e0kLTyaiKMHf4t6Nvs
nuugHpehK6bN/TXAgmGGU++55Y0tSeXwbTDCPrJCBXv0IkzBLp2eNCaG6m0W8wbW
inTJfLAwW2PhMOChBa55LYRijex3o6h+nBcTjf+SUILzw9ctCDxZrqOofcubHoeZ
2yIiIW9jVpxszRL9l1k+pBtZc+eakVONYC0b6fio5JSxPR0DqucFErO8tgxBBUR2
TA9xLFIR4eNwOxxGQvRyKc6l+jEGMH82S8+LROgxclrwUkfV5VEYgAU9h+KWW4az
PYVrxql4hjkNts6Algnm2hDY8fA3GRc49K6I7mSf3b48+5/VOk6yA0KboUMECt+6
8fP5DuG2IH+BEpAnf7MJVHbooKZbY2znb6YWSyioK8H66U9v4WhvyeKHSwQVXnWo
Ommo5JYS18zPizgMrkOUJngpls1Vc0FViIsSQRtTRaZhBWokOyGVG6agAT3yAUh0
Nww+puvhLPkPzS7HAVjas25/AMGSMok7Fmu0OlNTF+SEvY3DQC25ewY4WWnVg1qF
uXkxS3UOEBWUNqg6boXhLY+NPvBR4M3bhwz3g5I/BwI/VmjojTre8gVrBMfHwjbM
hiW6vKaUjp6SCk3g9jWjqQ0tq41ZP3VOkq+dPXKhKonLnDA2mP1fFXBcxSYaEdCY
ZLPtb8oa6moRDM1gDx19JPBmjGToQaH3DHvOUkfFBM+KQ6J+CjjupJlRqhIsd7I7
AGg4Qx66lIJ7CNp3iYuoAv1UwMmdjcbnIVKa3kTri5vpnm4oDlmcegyS4MMUOH+T
JkHwgb/P170JxamU73R7ROJEN8VlnuvWNaAZKI92OKCTEHw9KMhPcHic83a4r7fo
HHypU0AXxdnlYK8ZUL5Rf3IAoQhlK4pKuTHqbj0GKzD79sas4NyfsLRaR1pTQRYt
r8BoHkRKL3JbOkE1MB9gy0y9lgrj3YxirKWJ+SbKd0Zznm0GpJ6hzzrcRAP1wovN
N4CBTUH7ynkMcEpHJqf7tpXmCPmS6LB8QzEF5bE6DrACrWazCWv0Kn9iBJk/g1kq
xdTaBIlD/GJ5hwqYpqjlhyrLmCVW0cG0wVHdw4vfgH5YyPq14i7phqXAGr2wuHmc
Zgkre4JlTXxzr6iPsQTdjeoFn+YJA45Zt6d8RVnteNYo+ecZJc0fOOoMGwUuInln
P6dMYdasjkiAEKUhZ/w3O8xcOl7EUBxjHhm3EFhEDO2V7mFaenu28VKUArAVWysJ
KJ7BKXdHURqijPTXTlsJvO1TSa4Dbl2GZImFLZDI+MjSCCTEAu7YsY5uMmcPYGrH
G+afqCioiMIdwKE7B73DfGQy8Z9bVjECtDC7sVq17kvVch7xa5e6lINkWSJFehNM
tdmJBoL1G8FPSk5E5Fe6TJl7hNpyANPiukUXG9KWBfpaFf+05+X9MN47TNuHE7sH
lkLwpPorrE6ssfm3DtG/wAMBtot24b3r2kUpaeDKID0wcvdZ/I8HjxCLG+uOX2rX
3fLE6AeBm+QCl0WGMqapSzOLqgAznXK4ir0HBIo9+kSoSsnWTDmCIKfrTBuZl9hy
Vs7/iWIsI2uGxChkc9+DOubFlnk27utCaeRxnPRmXBxrD8lI7RPatb8tUIGgBM1s
xYWlglDvKT5ZfGzqhSYIRk6du4a6yN6OKlZ6QI03MVgq9v5KiqQRjJyB1UEf5RUb
c7F5qf4kFrSNO/8QBafuXojjVSIeRej9kYB0sy8PIimz+lar8sW0CDnuq0JsViF6
R0963ZHIj3DtTQ89aRTDylBfvojFCBHlRv4jQho5F2HUjFZknZinEh3d5V0dXV0X
SozGpi2h48rqQaUZ/E4NgWg3eOlvsaaDSMyW8w5tAClEwlMzgnGd29bfN+g6elVK
zvuewNITMVbqbEp9jsgAoseYdyNHa2LoCo4N+aBzQDI0u4jmIFqTWq9BJKQ1zt8k
rA5Ex7qLZr+DlQ4SS0JZ7AhmHLP++asZ/mM6bfGtEFidW1JcJzzM7i2wVpa3GwEJ
mt+V2bqdygXWal0bl+Erl5cE5hen2+rXcEnmr8ZLDtBxH06yW6DGCb5neg2+5a/O
6YMdIFBZXMB/p8+4Dr3QZfaNCSZqpnKQZuE2gLmAyH7wih4E5U9rAWmXbH9iv71l
HOvQ9eNPpKm5sQpdapogxsUzKuENmC2wscNraS55OczmVfJ33njN6jhAqr/AGOY/
KgbnRjBhUGVSaLp4SAF3Cge87MBbesvAAwOiY69XwiMgc7oHpbDid6qCg1ALa1PI
Hy3WVjDyA0SfGBkhixLMXUpsfAJSiBZHSj9oIgSOVc22QpVjZYfgsg772V/Xuldc
Wcnn4D3FD4JvYRZhJydTCde2/tLF8JTnyskv0MNtWfdXAtQ8dDc1AtCMRVYjdru/
cueG6hw9/mfwFsHoj8RPPHgTHLY6izsmbWBxmkFcWtovIAz1js2T+pc0ta+Yk8UC
if8vQIq5UTE8oVQkEDUx6ancMoqJPE6wCg6j/9jGEyHS0lJBigq6KqKI+VtfE0vF
a7zQorBeNEpF6WgE38yxoqjmsgmGMpS8kMRHE76pXhFdBAmNRqrlryRONj0NdyUh
t/1ux1bD+5cEz+Y0roDV5y7yRRD9l3ILM+28gxbeI3DZmxaG0MoQHTBwPhc17uv6
mijPvOw2INbgeu4LsNm1ynLefxkTedDuMw292HgsVRibJGQojVdsIwryvgJSUQ4+
4jz4UeLtXBcExfegkHj8IeSOu0CoUTP3WlfYlSYXc8+KRh0C/RdRQpSvVKfPp8fg
6zGeUUYgQDcTaJWpcCtyxS+WfwUPXmSH7hCWC6FU8IQICeNvWJ3IxWWOGuPhW1Un
YCmVgiMtB/GN1fB86FJfU/TN0CLDgmlury5LD8p/ojMn7ATr8xyYRYVEVqohOBh5
e3NQXStHjVTEujXZWke5BSpcH1sO1z51CHsxpZDdeeVtfhcqLovac45NkfVa7H6k
MgiZ23UsbdM1z0oPPxdBSg8w3lApon8ZU2cKQ5055t83/A9mYgTBwuNg1Kmp2JF4
SP5M1l6Cybq9XeWINuQbEglJUwvzttdO6si8PZjFA+KXYSVF85qmt79AgATRtRce
1BdxtxawxKvVB1AfzCCYCsUJZaJ1XSjgq5noOy0RrwXZqah7UuZIGHz7dNEXkbQg
jBfKJqp89CacdEyFydkdwQ==
`protect END_PROTECTED
