`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrDVqAydqxWmCIeughaipnsLQDmI3gjbGsiCXQygBkdVq1iDllEtZBZC6Nm2nYxe
4n7eLFMaePmEAPaUa6LISimofx6WAkYxZmy4Aar6eU03FuxMAg+LDJDvDr9IpE/k
RAZmRsSQ5IVs6bQ6KsqigpFs2QgLZkK5dx+fHWBH2aQVHLTpuLVuVHfyK/Elapg9
tY0JwF55BegimRadkGu6XtQwP3t2nkOcPmCZ5Q8RSCfxVqmQJRBlNbPOnyVYbCHJ
FeMKaJhqbFCL3ddPD1I25cCmGoqX82i0g9sAAc0e4WMB7lDn3LBRdTq617of7ZXK
hI7vGjzhSVkeiKbGM7s8Gh+3Zi7F11ByJKYCqmhc0YXgySCZUVO/RRL5CxXnuM7e
cW/XVQvQ1jlIq1qpvkC0ABGXUHq3B/0N0kQ6gNwIKuLOMzlhykjxW/vE3j05LelK
S5GpRslLcDRBn285Tb2tyIcmHYNCzqgpET+v/g6pj69OFNhXsKmB2SfrcQ+agE3+
9R/Yx/aZvEal/X+hCqe3/VHmjZ8mrjZJXj6ghoW/ptiTdG7yteK84TPlaCIHslfy
I6biClUvDeqvVZbNORs/d46FnpCIzd5Rya+PvZvJ3EsFyq2ihrL3HglUosU8td1o
`protect END_PROTECTED
