`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfYCshXHi96hmtGJMmelX9tnO00XkFdc7WyGDOmQ5jKurZJj4EId/kkuFbuJzj5p
5F3z9y8J2WMEZjsJbvXEIfBGeEG8C4vLjOvERiBiIPSrFpKAB4ZErm/CTQK+XFIF
aEDvJysb8VmAyTD71tGB3FszKY8cZIcZUGxA7j2wbgoU/PdltxH+obGX9y2g0OUl
WWBZsdrTbgSyHahVmre494csehdIc9gmTpwdc7n1TC5G2k04IM7BIhOl4wwWvx3u
6rGI72+Wk2KlTo6aWEitQukVdZZCzsk4UXgU9wRM++53NiyxDj1A6EbcidAcukbs
A9B9Xb0QUbKLrwkZ89LUr/soGt9oo1wy0yASpjs7rdsQV14rwgJ4+qLXJFGKkf+m
ijHy9d8N67t/JYWa/jmvWIbYWpGOs9pNx0UqnXA83DW2MnYHyxgRBKmlPFR/aRZE
DIJbW2ZuanLttVCLP7mLVHu5SKm5Aix8gawDkwvEHo1Jb5WCYpryyDG6EL4qEekw
1pRfYmaDWUjcLKNHjc53k+OifUnnFeRdebX18CNn5EWc1a0qAKQlOvCaKo+hndhZ
S1mCSz9I5PmzZL1Zazbj/A==
`protect END_PROTECTED
