`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiCreSt3xk2bhXJhJ96FuNc539gRB4NU65LZao4yQ64f6CDfg85l5CW9AKU+X4Ua
jKjkoBIb+PvnXzawWEVz/U4XbN/F/M4YJEW10mnnywHQ2EAX6iOWX81/y7kOBVw0
DnEpa9mvmfrNyuaEAm3aA8WmdPvjgr/M/y2fk+6rH5iITYkiF9jKeiweBnYTCDqo
FMzTY3loXnlffB0zwWns9lKyegyH+ZZ1TGYEx3wWMmFlS0XHLOvh1tyi+b3iHz7N
E4+xwYtNwPicrIw2RLk6uUTbnMuU0Q12tX7F726Mr5otSUHFWouFHJaTqcQI4nDe
5371R+EtpxCABaO+gZ9CHIRwKK04mrkxk5mukUPDfBjGiJ8Kz0+q55mVhq09Q+8k
j6qrjuKQCiuOJ+ONXI7/rgI4enOul1ljzsAoPaATdQ/26IaKGkiot5pMcHgIYfWd
9fxTVrHKTOqe9PG4ny5QLkqiWADRvb09jc5D2XKdUUZDiF04uP1NvOTRIzurViO9
`protect END_PROTECTED
