`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EjC3nsrBBr0zvtxswmaW11RFyZiNGi7i14/TQEndyUO9pFWnCTow4IfdrKwX4Ro+
6HCavmZWK86rO4VwSwLPEUxshWtvYerYWqFewWG5dnUMnEi4PAimm2q6V812xDzk
iqq85sb37KDP3TZtflvXOCbbmyKwdlXwvxC6dDCmvJqlnH1zNvtgWuQEGr7Sd+px
A1p6TvKF4UelGNkbCMqIlCWWe5S+KHbd6VyNXZ8FCrn9+jki31twxNnb85KRa7as
CKkW2qoVTxKeBr9MTuNfQCv8jkqiPYtX9uk7SEkv7GYaYNumgEV6Vl8KIt8qsOyv
TVxJMhPOmWlJcMm3lKkpuC/K8W3TFYPeRVB8+8u1O2RJCmKTp4i+zUdADBEuwCkW
Pg0FofijaodA4ZVl23Wghzr+eOQ1C4ggBDiXT7rlUilDAcpas1K8Ft96WMJ1FCfh
4mEKZAopzYK4E0Q2pIz3RIqujZ8jPtDtloX4/rHrZnTCHSmUKZ6Ucl/8DltsNcmZ
a8/ayjxmtqww/J0goKfY8glhFzlbzMs35qcgFrHL9DGL6e3Rc4losCX2bWyq0JXz
Rv9umjEkU4xK2+4mr4FD5y0tRe2I5fGIuoWxaPnTiM5mea0KFwQTLhIGjNUljkkh
l56/ZDiQDUUFU6YIKKjKaiS/OlzjmFNDDgRZiANAGtaI0IOoOJ5MAg6CkguFHrML
lPqFHIPgQluLmbz5VZ6nNe1+IbrA771u0C8xRBb0eAefefFiAHEktzFqxcRjzN3H
eep2VqvJuYWQZZwnmWItqAJEJxR8DVrs8dCLdR60haWoTOt7tU6AJE1u17xJL1nb
5DIcNVrhf0iFNWJH38/k8PipzrOaRCEixUMp3SpUSOtos7+lTEhe10vnJYMF0KxS
1dCNelrZUyKJhO/FKrj9UjYowzr8XjGuvMy7Wz/beGA2fEKHJx5Xw/l1Dh8wSoFY
qwT4ai7ezXtukl39nE85sDvOCrZDwIjVBLUS2/Izqn+JesT5PiQZV9QGX/FfV3wz
jRCtexeeI77/Jq/7PJbNwpz8KB+CJVxtLpJ9sq4pIH0G1agNs6BLiTa/RGByOTSR
uIpyR4WQj1DdJJFzaFVL1L0rJQTlZVr8SxktZjaUgxreRn4BJxUecSJNE3xWwvR0
RRyBoI99ZDL9del5G2eaZub3tuPNQbLQys4YL9RMmI3QToBegDwzf6QxR6ZIXqNQ
1ym09qf6mzVUeep0LcM8kN/kafeTNC+5E4LT/zOXZHav4GG0TxuOw5bfE8xM1dfJ
esZ6GA45sKznnmy74QqhmTtE9Mwvelu7+jNhAeOWzCGAhblr/QqRJnjWk3KJl1Xz
7MHa/hfmrfj63nWe4wubpB1MYkjoNC2i+E1JMDGWke3al9MogNz+qEIB1+RRMFfm
rvESv1j70/sDDQnxCq1cRItU6rU07w2yf6g3RuWT5zBkug2J6rbUghdM6BwQyFCy
HlaU66fB7+Evl4dZytmBagJGev4Zs/Lu1nw9ER4zbQkthPY/9b1IKSOYNsgMV3/0
RAcnTKV8aY3G4a3qytk/TiAnvRqJ5dm9QRV0+0I17TATtuGgCGHB3i38+KKQmRAx
l1cQdhusxuWudsRxNqd/W3QMe/v4ded/8T7R8y0929JbOt2MD8c3EdGBLTLWr5BK
fL1Zji5x95cyBwhHm/GiUOp9Z/T9VvZzVmSwDRNLgnWn0V3iNLh8CJnEtQNuRzij
BeVPHdWAeOc+t8CPzu3H3QRy7RdytEbPFpZh1BaXPTrKBY16i0UdyJKL45H+uhOp
v//PFI4x09elwfy6qjzd6uYX/swteDIFZ3WvzIuyit1cCYq5/RgxSFfuVB+nQhGl
BuAc461WW5FM7rSUGFjqcwRkxYAm3nsDRMLYMh+0I0249iBXISPdhaSDNwaGbsKU
R3bDryquOksPvxYFnpQLS872QvfVCmrf4HTY/V56SSJKC4jBXEmzdV1tzXVPBBoV
raaNV4mAQiKxv8uVEdpLiUvs9G5wRUFMxHxpOrUOC6ev51M89YLMjYCvLTcvQGxt
d/MMKo9eRmJUVAu1HWEwbHYeTV33EYS3bFKFz9tj4RU=
`protect END_PROTECTED
