`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lm/EU+IU8OlrQD0jf8t8uEu9DrIr7WN35pvwuEM4CFg6HCDvsCGS0uYkp1mjIl+9
DuNn0MiDe7Fu90lQZs2qW/jYLOxHANKHm40ayJyjCqeUo2BYeVnFFzan/uwoyd0g
dxgs/UWrrltXlghGDy5W3o0hJYW+VrkiAHPzs5UNDxKh+6ssp4zOeWqvCZMQBZQF
tuvQnBOVAo8mZosPtd6ZisdBLsCsAuvDVoRfWG9wxW1KH6ShIiOAglzhT/Vnmlzn
MBSb2wqgf5r/zeeOagX1vEf27wgJGGga7bOPuxfLb6IhGZYkood6Y1LacbQ7tRw1
szof1FFTao9wqaBzxyCilSJOwEx9Oaj+qido96q2Ar6K4+ptx3U5LFPnZK7w6OlW
0HymOiYtKIeGNJTpN8ZPfsvRXgvy8Bud/ECVvlrKPaL8tuhtg0xoxug6OyEyVDvm
Bm49vPNHY46d6uJa1ZrdLV4ZUfq+UWvtTHlyDS21AIey4Ny5aDDwocgdHJnnJmWE
Qq20xB3ERooa8k2b2Sojsd4eC2ciL5ManM8idefj8pAQlaM+A/PAouKNoYbqBJKI
I3NTnHdvQyNpqH55pFf6VWGAiW4eKCQpt5wnArhGdWrQYt8DKZMvwZWiVPjoRlXE
aRlOR6icPN4+Eq1V1snru1+u4jRKE6XSybRE47GKCChzX0uf8k65WuOHv1wcQVMP
j9d2c2MfdSfHkL2V7qyNqXQVgojiMniGEJGxKgVeVrgq9DP3CYByUOg2m/LUZMtd
fYlr/7p1vTYwZXVmDi2+j1Sxi2P3NyGRO6cn3LB0vvvRObicXcQ6m0BORsiq6IUq
yOSTUEMWX3FsKSwc4RPE0FuugTlwbUuggnKhA/OQjz5N096bU3o4wuxSJDbyBwve
OU1SKDrGokiyDtt90InBOGN5bZoJnVUcxZAOP0uOP7wwuWtAIlWNDsBtL1uIbTf1
JkozXptt3x3+mvWlH328MqN2aSnxsy9JatrxbqNW9142ncJiVAZINtBR8rRvx04J
Wbsc/xmI/Bvyz6ZnWvuqKQ0GcMsAN75zK4U09ofXtNOrYMKP0TAxybJHsD34H3+g
/W3w1dhIrh1TbU/Uhj6kwiG+Jz/Cw2bgCD30iDCyET6Cc8ZeQDciFBbmkNVSIS3C
oXrabN/6uaABqYMjUrwq76MrJht7g+FP6SQsRqHjCuZ3fDjVYM5tk+8zmMTqaoyr
ex0yiv19y2Svd2RStxUmO1ZWUAxPOR+UE6hskgAhiZl3b0CX08LWr9XrigcYCnQX
/T2pynXsR74epI02IY/m6+lXzpGS0uNdCE5gCu0Fem6SRqB97qhyGYfUHbYEGFrc
JjyPLxFEhmdSh71qPukkU6kZpsNoK9ZU0mU+nk1pCPUroHiCHeQV5f9JWlC8geJD
CuxTM0iC+qeVEjzvhPCxEhndkpmlRYrCYH9jhMqflIyaqAxsGZjiZ22Vi6+redOb
aehUi+Nl1N9e680SLJwDa7QFbvTx6Y2t189Afb/JjYa5C+uHnKh6hkNz/gVkgiqv
f90uadnDeimec1zI6MnmBcwaRAPdqLo7REWOnWW5q8fqpTpsR/5TpC1ZRrHACi75
IiV2Nc5novM9SkS97K4Mvisss/5VqvYKalGFwpMjSb1XNyokk8GTWbyllLu3cALl
asLgKmdkxhKb8hIADGfbaJNsTzIVH1+flVeUgsKOOoImN0i/UsMABUIBKvny/m8s
mHC3o9WmtircjCQy4N5Voi/GeQIpqGzTDw7UMq9xF2hJh/QZBvWE1EX07NrR/qvt
ir3tKPWpVDvqadG/OO97GmHq8c9irkJi+AaOO+kK2paMTBle4kpW3E2IcyUeZi3h
h5kBnot5+0d51a/hvQgSZKVlqZyVIEO0zJYOI5fjpN6bF6auSfZc21/Z0quYhgRc
qO/1DbUIyCUhRV2hnCMpNw==
`protect END_PROTECTED
