`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGrbV6uSkFCRtLazVtAjs4Cl+Ze6RWt63wChgHfCcFYx8VL/7ZsgOj8twZVziIeQ
paAp6GLfMRU1VordI+hVGXPjCvnoyrQN6VvnIYTJTmoL0xQlzNGI9nKpIb4dZGpL
YJhG3B7PnCW1DMV3xZYViIzRR/x7S+FY8+anNjwfE1p6fwFfeszC5NTvR6LAq9/+
i7aCXFOMSBNJHpqEpUbQSe2B946J4SrBli6aNnj5qr8Fh3uiidijffse0lxD8dtW
gg7aneW91bBJvyxeO9OY0WYlqhwqR6sFE4zgrbji4ZZBrqJmBJ+HpPoSCkCwgoGP
g5EvlJ8WCB5ecodqtzwVfbqiBkdxpNA4+d/8QBtqE6TDPzKe0IiMHg8VWGAMOc1+
YJrAIU1q/U5a2nHk45p/l0keqKMPuTczCceDXjCeEfouGkcoMCpK6HSgG551i9AS
PA1PXlmBfbFvZTAlZD1Ja3E6D9DqepgS01jTWVPtL1Q6/VcOOQwHGC4W2xwxl/gl
TtaLa3lWlIfk25JuIoIMbRW2+HpLhJERbDg3nxYhKh5CkkNr3Raxs+y+HTYvEwbu
qVdlF4f9fK2/YdXWkSnXQsc8zDfEb737JYQV61RdDQU4b/P6wacSbBRhJULWgxJ5
dHVFHN/AQF4XKKAxneCIFVhha4aXKYPH7Jj1tZq86Ol3TCfM0fzCyFIE1fJyXU+p
hBoQfC+kcB3BBEeQTeFM0R+CUI7J3MDUdNitP3AbZ8HSDDAqmRIv3c2P4TiyrWg2
/o8NnkoVLghG8pNjl3jGTqRqRak5lHw1B72iy8qOJyMoZ4CwF39rhkOHgyT23MPQ
/Y/fmM4VOBsQ9I6Peb6EVMAr3xYmWIAffJlMRE3RzgKg9aK5ugWz/IOrkfA7/2/E
Qp9RNYISMbVH309MFi/vpWhQ7e9+XT6Hpiru7qJ6382gQPPR5SXqHkr7SbdJLTzW
hRtlVB8RkqmfcH9ehzcIbnmCvk+WAQzUfsmIVxZuDEN2uwJa6/F9U+4Mvl6YL1ep
lkLmdwp5DxbsVEp5y1K8foKDxOaW1eBOb7DAafHz3xYXrMkr0+wyQu+Khu8LY551
/dbc4sD+ojILLinKDhJaEYajvuBOCacxOfMDR1CDejaOPhcTcEI6JRqfgMUCFTzp
dvmS87lFjrTbfkQdCIArBLgpjGgNH/9hXrxlul+PNlQ3CAVd0V46nud4GqMvNt/c
0a+4b1OftVtAnClxA9avziBvtbzJaW+/UnsXa6Tx1oSoKF0AY2hgw2q0qHh4k6im
2d17UJLiT2RD64+9n8pqMlZD3Myzq73ePq01/IWj7+zxV5DbK8V0W/DYQL2yBhpj
SfbpX/s7V1KXvs/dPGGq8p3m997CIfF+rEtX+PkYrq6J6IjzUy4Z+BbMBY4aLt+h
O6u8WyDg05iH8EjDI9/vWXJptGrXuISYRe3UoaPM/rG93rG1DWwBrgEQDfo+2MCL
zR5sb3SoCs2U1WKAxkRd3QGmIK9e5OqU8vtNqhS5vk+5SutRNUVP2eN652exzPU6
Bq2OGa26d3QAGNPjvj7aSO/Yjg2dosHECKMc682AhOoYd88v5qb1PgbWzJQvg6MH
6JxABUuGVcfBuDujAeFlgTnWI/m/dQ9NEKEl60xHDhOX+W2/EnWPOqApzw2/QqgA
LbaSOCdrdQ/Uegvj0W8FWD4u9Yj4vqDdoLIaxZC+bXju9X5nUwTAbj57obRl35rg
ueQRYnVLZ1ep/I+FmKjk7yO3gU4eklHHTgdv5gd8fJQauWwyeudJEL7yrhwpVogS
57M/Todg6ImiZ4OZBhvdiwymMUHLfP38OhUUI81Myn785ETQRlp5x+tqmNWKHz7u
fWtpYsDR5l/1BbHzCHt98FmtlVvfvjvtScU6vJnrn4hHv/2j00kpbpV9xhmXFG0p
QE7LxMcuyuamrMYturjK4WExPHXXvg+MSVjKGHUpVxA=
`protect END_PROTECTED
