`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
srrR/48YoOvZjkbBPS6TvOU5BXctyS3sPa5jnA2dajYobjYWc62ozgcdpwBPHzuG
cDeUgl4gDezu86lTA+IyCa2DvWAFweD/4N4a17dJ6vflJ+g6HRhw82pIqZs5gKaw
qcwLLriu0tnN8cYSfhzDhlqcTh8MAhGJVO7gCbvStnTCv6RjGn9FlVWts49qrSwB
wICXBs5ALAh1pP8xulPAZVGv3WVTXiFtAwXGTLExVT1j7gQ/Ll2tO5XHzPa04jKR
n0pXI2EP+FrMx9Zh0DI1k8n3ZA6zY78bfVAP7YEW9neImKLqx3H1bee0WdHJnhpK
6twW1Mxq8Yoh0Rc7+6o5dWfoLRW4hVWvD4UAaBj3k6j6AKEAL6FgaANDT84I5v02
pC3CDxjkT4mCRZ3o9plHMQGSP2EfaX72vPs9p0XEHhgOVeq8TbivSKJWVgMPzjPR
LOZic/Hpg82Ly4CBDwD6kXWdIvIAYQK+mzhBvE87IwSuBymUNqkX3IR9BETJOPFe
V96BBr/4aHwFTQ6xsopUIK5/mTPzlky7tP7fY83iOkjCLInaeutHLxOPTOlNFN+c
9IA6d0gGOfr7J8Vu/yDqWIBQa7l2BVG6har/kKk3aW6FQ4xUvsfvKlOZjXWcpXIU
oqfD7C0+gSP3myh75DZMX9LYFUOks9QY3KpwyFL+DSSVI9ngJkBQjZ6qLSCrswXr
7E+C9S4LU9I8emTli6ItgJ4AFvJxrYl1TawOGsICxyCVGFSftEZB/sw2yvg/JwsG
ja/kyUHv/guhHPATzayKlqThgt5mEjizHUfbONCXkpQQgavzLMGq4clqNu5np6SU
Gqw+ojj8VYVEwFfqSMO7jg==
`protect END_PROTECTED
