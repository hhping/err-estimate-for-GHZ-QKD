`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3i3MpKt9HlNCiSLgFnpjMo73Y7S/aPXO8niUWMW7PKfyxkM1cuksCC6Gj6bMu6ad
rgrqdVZ0JJL4vCCZoTtJR0jJNu1rAXj8ARZKz9hE4ibnDLFr1r+WYUak6OpoTgv8
xZrsT4ZeZ3MZkXys29qPoBLuaUQdwubK5qYPVKl8bda2XE5Fo+ZNR3zts9jXKV2R
Z13MN6aoM+RRpc32nS588i4Nw/StfhL2/PNQEmSeeAf/j/UBUwVwfo+eyItmEj82
8T74SRr/shjYeeqdNb0AZhaEmeTTZmXhBl34YM643Far919Ug2ub+Wc2Ac3K9rw6
jMCh1xAp//mVEAMYsVH5uNYyl6GcfI+1WwsLepy2QK0X8vFt0ooDlQyiR3IO/Ke/
DgnoP6ril8ubxxTJaf8Uj7du8cezKLRfHzgJ7XP6uUhmsdg/+7bgTLVfjy2naHEM
Rhfk+nRGSwn/oi+FIwoeOIGpAxwnZG3F2VtioVJnRN5CEZ8ogkobzclUdWZQqHoX
VvRJO9o8sX4AAFLGYjItskWwIgdO1BFYHrT+w05157mTImkck7aa2dhi5J1DrLd0
HPDNCYNgM3csDlf45Lyu+WTNoE8gap2SselGAeYC0lhagRu8SIr4KEUoex7r2IBa
`protect END_PROTECTED
