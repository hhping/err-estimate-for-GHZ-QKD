`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZl08G7JILaC7DkkXQMlloqOmpJnB1Z5rxMJaA1kLJlyErUZIl2kacbsjhQ21T9k
6A5h4lJVkvX1UUIfAWXb1Zu0AFGz0G83+XygkYwkS1aVQQuONGQFam3GCo+N+T9M
mOS2m5BY+SIwg1JAHsVLSsFWHYwhOsAedIDSO7W1+HDVqUQZ2l6y62fAwEFAPHCo
`protect END_PROTECTED
