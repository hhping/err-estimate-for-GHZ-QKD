`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkvFHbhRRYvyEdz9iKWayYRUvElSf77RforYXwnxsaQHQuEoiyxGiORh6Q99F1f7
OM48UoX8Utk14Gi82o9EYTsqLSQwK9xY+s1ijwHFf6SLrAEgquhv1f0JBS/vZSUa
sOOMwvAMags2KOyMxFy37AFRUjnXF6+EFzRncB6ZERTwrNu23UHMA6k6FSdQ7tY6
Ja9cnDa0FzpCRG35aiY6MhQgN/acpzSAORgAYn6zJ+oNDHtcEpmigPcRZPkCwSqf
xfnCct22hUgyCTzaBav1HEuqPbN6nmBHUghXYqJiasaB3w5NYGjox+eaaM5haQKo
0sp65lCgLLB+crfABPGucUyVrBEhk24IThoEmo/AaAsIyd2IppkjlxrgRJUG2lJa
6CRs4fVm9geVqyCchw4gjAPd6p1aK0OUIurR2TFHqxR4874cnBEvFXd5Zr7lWUVx
Ux8iOKkt1hQsoFepRWEGysQcRICIjI+xmGsz67MwsHBVeI19eUU44yiW64APymHm
lD0bzDHj804nIpytKiGI+XCBrBY1HYv2g9xuLG1mDPwfgRv0AnQUBDs5BGzOtjYC
Kdvcko3Ym7TktlOoSwGZ1O6FPuwSD2SUupgfX4NOelL4PhmT6P6tqBVpQZngtMA2
HV4/pWqeeH+39s0CjpAVJ9N2dHyOhdYvlMDmNSQ7fs6peers8itbDdk3R4XxdSLj
CqAjW8cvm21kLX7Lr+oNMHHs5B9t14glp3aOpDD47U8p4I+F78R6JvNWYNoTPyZU
cI9Cq3ZuWl3MftUSJ8LXTDzFT+g2NC/uxfoxj2+B2q/hAaElmxCEnR4M31FU/cCh
wHp2+kdArWi/VqxIOgrktg==
`protect END_PROTECTED
