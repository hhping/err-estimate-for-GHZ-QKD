`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6XaTyOSpp41/WLLJ0WC1BjuqOzb8rzb6OjNQVwD2LEpQ7kG3dDd9q59fXgyqiEB
cHyCEEFAa9I19b0OZsFNJ4Zva8yQkm6wgF+AuhzeGgOrDBVgHjZN1QK/cQ+WdVUx
WHcxCdqGE8is6R+ms7TBJ0q7dgeYo0EeNl4yCesCXdk7anIyTvaf63q/BLXgvvC1
DQy78TsJbpRSfgUTIct2XFLXwPnhC78XbS2eG9Ga270doGIlBuDdUpYCm1g+ROIN
UAUJ+jPw2SeiYv3oLDl4jC9ICNEG5Dvfi3WMOGSVswp01zG7PQAR+meBtyLeHrB8
L4/2E/ZRzAaWYEqTBOynVMoaJWDTnhK38GJ3xOOuXNu3Ckf8ER9jehoZpsMDMLTS
fCX1MjOfv/BIWeAg2phXGQqKbh2dTolms13ho/+Uju+87Rm0Sd75s8k2aThq9Cdv
DpOjGihrsgNPZFGSL+8IsdvbjMpV4bWAhibhFwEXwqbUi6mF9hoMEnU84v16GU73
l83NxfEf+Ew3hVB8tW/R8nQFbI0znoLVXRQgVWEd2yKhJLA3k+g1Y3pGq7hRgyso
G6I7J6wTLEMggno1ljnJHJFA7opV9y3Xo8pE6bfcj30FYTGVk/kzQNdzyBZ+JXEd
+3nuBDQInZ65hKVMK1Ej1mmaxcObnBDnftFfGKKzVBk=
`protect END_PROTECTED
