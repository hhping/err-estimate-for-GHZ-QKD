`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vXlbxXbyucOTPnc7s3CRQZPhOq5pu1ErRMqMdSx9frpK1JBbObfVLaqlfeQ01Cv
CAvUlfNRQ4TBpZl90FnTMHh4qIkkDu4MNBZ7kB90O7CfK35A5gvOr2F3qjEF89q3
q+Aov4CZbaGJ7ME0bkJD84YnQOoX5fDNF7G6m4QVJ8kk/+G/6hCFJOE4Qgvs2pH2
Exv+9sOIiDX/3IGZl4Gd0TiS5BRpZWtDJ0sMcuyTToEWJMs7ohSTZkafOUHnXARH
Q1xjp+QvNDI+IY3byLjrtzWY5JbGwXThuGMJd+lF9a5HsCtOk0MViF2+0qGdckLB
3AsOwCuUELL8vOBV7Jvw2HUUAaeaJXxVOfjeYUDyMpUT7B2nYbqiMRGevCz9vY+r
m3cJXEJCLu/F7itnJ0Wgg/gM8vuy35dpQ6AfYMvUAY5kKWagDmbSkxlPLkmdKO4P
72FlxkQ1ufiXraATWQNj+lSxTfz0VPg12ugsI6p3YUoyaTHeb22B41ZS+thV8ydD
WgQAHsk4o3PhLxAdcC1ehtVLp3icme6JWdBpV9bmWdz78B4W/PN3QmIg9wJzhqJm
pWw0b0HNRarYjfOXiIrumv20FN89uZgb2DvoEhKjdKuLN9Jn2DVUmEd2BA25jvPd
`protect END_PROTECTED
