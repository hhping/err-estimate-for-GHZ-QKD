`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCv2bmXA5OsOHIZv5iRkXDQBpEvuqVfxoEai4qg8baTJCDQW/Tj1M/B1ZPSrY9EN
GP3LzbxPChkkLm7sBBL6sPk3SqazJeQrIEoQeX2dZVSntJ5T/EDNLxMFR1C+oAn+
Qhd5dSzTeSrPlMjE0I8FUY0csnw5iPnf4KxyJJWomAVh8TLtc4lOPH+3zxyJoHgE
zLOZ43nS6TORoUXovgRHEPLDH9Qjfh4Kqe0a5LG9cIKus87/2k7wIfXPEJ+PPsLf
Zi0LJQCqVo/x2vXcTEV9SWG6I161QZyNhqrikXanj4fXWzt7Za/RRIRrASF+Isyg
9HvuNHE0oeC5fSmbxACLyIR9oqvFcb3vyYh+zLm0adPOsDDaslFoIAicL0JTm2fm
C2vaUIv+xPTzQxdLkDR2iEwv8JYmhaEzTwLRhZOyyYXxiRhJ5Hv3uJ7BsL4l+qwU
KFEU+2Gq10+mVmPyIaHmwZNnqGZwNR54NzGR9rpJmEi7Y56zv8r0PM7/rXftbjau
3Y8vBQQ56EIVGGGwvKmivgZsdPILCGRobqFvamiGaofA82jvNpS9iX6k1t5aahSm
Ozv+aiBdlDUkR45zIiGlvSTKIRoqNs33/TCPz7sAALQ9IPeeygG7VfaulJbFW6Jo
nTBY6m0FXjw9fc3ta0CUtz2SbHIx3Zr1k18AWcLWM0jvsXhV67/h3csDQOhzDNeL
7PygE+SqgdBWbF8t9vmuKUvDpwzW+fxOitOo3uVZ2xph10xIBGpNw4JA1TL/slRT
PJQQq6soEZGMjtH/BRFu61Xt8WernZc5pMIibS2qseYVJEDTqtjEAhXYlw//UeqU
8gM7t1CQiSwQs4IQt5z2BmHKqVv4BkmbRl2RirP7MVWCS3ImW3b9+POtA46II/A/
k3JPRGqnJtG8w/2fbja0CNM3ZZdEgZGICEaPHGwUFNPBNSBPNVk2r4Timtf4RKGE
sliQ4sE9bLQzpjUYwfSe5ogKd/DM5KV9N4TTsbmqOdigcypMFUt7/EPkZI4mBbqT
uX0dAWcA8SxBm0mDpHwTmb4jCvfl/f0g0XYOij6jvZ1OqlMhY7KxyfDsopewS0uW
t+WMAjU8YkUeA2IY789m948yXxRVa56S4EVxUHZIZSzUTXfYN67qeniYTGzQfqMT
SYRFI6GNatsIGR7hZMH7BtOYDx/9JzMjZsDwA/hU/TJygdQjpcayzkyLAQ6C7xnL
a6l7Eff5ikoErUL9ri17ZtlGr2QdpmtIl6PmGoNfbSZY3NAZWI4rtZBe0oZ4mY6e
9kQWBevjamqrNJorD4fc4qASAfk0rejxrcX/l9MD0Wl5z37KkiyhyZ679G7xDYq0
2k9zBe2tXLpFrzri1zZ5gjTV0Ruys4UxnVAi22PGPrnC8+SQSwEsWQCKt7mo5WVd
HgYVRRmN8j+ZcrSzcNqnaK6aZN8XY//4p5axxU+gNnW9427BYKOtjEh3PIdDFirL
VYytLpdZgQ/2CcwRBWMwPGLtfhmwGp0E3tDX5V3pu73zzj5ZN0rsr+0tRVuFoiW+
6015/PTkUOXHw0BB/XvlU8oUefYQePpuerXgBpPs+nDm7LytVewpYgyOrZ1wA850
ECtAQfe0hxJXb0PpVgvOshGQpc0uu3LWucn0gaQ4C5JZHigQ1i/TGgi0+Y6YonDi
HJx+lMtXUnv2kbJ0kHLw3Vz4UUm0Ev+gTCDaAf//BEJx6HoSOd4ZqUxKq0nm65sG
Ve1EMId/i1D8fOWL41aZ/KEML1zrxM3hl74OkT4olZEmS3NqwPjJ73IFdgB/aQ+/
YXV2queaF4OrgP9L2vQ67mO8IGDqTBOKPr0lXmLkJBTJjosKML0LyIPJDY/rBGDy
j3oE/lGQwaj+0xh2f3TpHc+Otg8UXis9bx9hsPEafTS5yyQ82MQIGovMFoN1aAZW
kK0eEyYBNdG/aHBOv24y26rIg0zq6bD6Ivf95pnx5FdpsSdvsQPYerbCMlmLYIos
iW99JqzYEgHdj21R0EPXp9jUTAe+Nq8f43mJFQfbbstxvOBcTVL2w07YzJXtlx5E
qToCvtj9g15r5Rel8JdTBrjtWCjQfJWVHIbcBcxq5qjPjgEOkDApC+NvHS+0uQF7
iTUL3yJBh25RvSqreQYlcV+dkNL7Ea9DAssnJ+TWa/vScgd+DXLeM4PFXD6+02bi
jYOS/MVAc+DRAOXlPqXUl0N3PPAgePXyX7ixSHEp2J4f66+2eKR7qXC1hpy9Vj0S
oyntoj3Bs7pE6fd2cDn7vP9KZ+apVdeUehDJ/4sLvdszxqYIeHD9cBZ9QjxZFdDw
rBEtjmzXruCYnIz/gu1M3t4LFKuSv4vfV9Slde7TK56yjq3H3PTr5aeD2Yxq9LLn
iAv4eNYI1m2sfi3r+o0zc25N+QIhzrEkhyPUY29+qIrvmNHIxdzILQ46Dz1oJu9b
RIy/aQwUMjShSDqEBjNNvaMIk53et2wsyc9bD3tq3NqpPBRfSwbyLmpV05YMifqq
UDm6XlixbwCYN6WEvsUR9bUgqHRzflY2T8OyDmaZIhEOkn4w4dZ75loHFgMnIYMV
ElIbwBBu3Exv3nH/dRjvze7hCK7W8fkpl3jAGXVvl9AjZxQS5wur8Zrky/n0WLkQ
eO/dC5y7OYBxBshV9gZnrTZMO/npUFnExcJZ/+QTiLXVzENh5H5Sp4IItlibRmjJ
jsD/VntHO7s9QbwSNcGEI6fschmN4CQtKs63lJkJVfkKW0gq4EzJmJDF98+1dqLi
BYQs3x1s0v51x2n1kJjybwH/chDeHd3QO6udaiAtwlIKC7O1jCE6zBKEi4bHpv94
k9XVxd7Nz9AC0qadc242Nz7aIQfpfCjh/xZy6NWwJPggloYZjdPph5VVZI754XY5
M0Bd2Ke7zCULjGrM/CejayBaQw+SE24dVlgTedYe5pCH/rRm1s/+rn8+S0Qq+hE1
mwMOJKwQVXL9dZXHLPeqe0SAuz2Mm8VIXO7+c8LnmqE4lSVvijsG+1N404pJXj0/
9W9hnlQQzNHIHf4yYs2TFHzlLqiUKw1YJFdWER+5ezUuCppgdIYTeFvEEFfiy2SA
cdB9XkcAWjytgtxvccwlSktdnSONkhvg80f4Kknfh3Vu7L8sIrsHyzxNpxBKrr8w
E5O51Vp9Ic3XeiFrXgvDCYmfu9USb5+VsA6Wf/UQdu2qZ01jiI9dbFt10Q6nr96Z
HoJJ4FYQq6t2GRmz80oK4YNZWg3D17Z2ATOy0Ttr71GAlVs5oAbHiP6/kmUR2sd9
LAjBaDYyoVld8hxdx9twlwX8nuBOW0LnRH77eobTCFc9HBw7BVUxYbJEbFNRS5t4
G2gW2Jhj5ujDGSgiRimkN+umUWgb9yJcCIVPZcBr0RsKPEPX9XULbbJxJx3V5dS2
sVP7A/V+laQ79lW3+ITMbZYVDxYROEjUqu7OkQf/WsPtjimApEI/V4nKdbsjrqDn
1o4iqRuzKpgfIkIEAeKck34kmkYPPq2ch2y7To+9pGzMWrojB6UXQPi8Atw3qmBX
G/2LMKqGBRN1gyYYQcSlJ4IHOROGjCnYqXWJSrjgXvj/lREXPZYvasqaIb/Uni5X
vaz5EmpMYmtwL6CQAsXnces7ACXOxDgr8WG1cL7fVdjvVL9X11TW+gmR7bdpwvcp
8tdJu2/X9xyrz8O1GVOSzekEECoXCZfetlwWSATpnXvMrr7ihjRKNuj5Xx7PwWNI
xt2pyoDckE9Q6PQcQMirEqnxeECRVDpmXEUjCClCB+upSiF7RN7ukgpEVrgxW+ww
6DMo+7MZf5/S+tlKxDlYv9lrnI+i2ExpLAdW60KpTYlVaoBs6VTIuj90CvEsnL24
/eynP88aqmLdmqBRlyz0KmZVQFx8o81OZnxsLnSzRNTQviXkI2fsZ6d58R1AmwyF
OivhMBPUcdBubqShXrSfANgcZ1Vxl0T0q3TwHHCkv06uJ0X/sQr/xhCa41lXBU62
Z3vA+EoEELCf/xgY28k2P8VE6IYU4eKLaWz9KK2+7/HlgrGgZIikL+LzvcEaVnrH
8N5ynjyrjLzdT0wjPPaaXU24Ef4Eifk21wibaxomnl2dpb/M/QkU8jTYghLczt2z
wzBhVtO3k3lhQKbx2ii2Yw0MM3dsbbcQ0I7FNLX4MEmKLDnpCJDjhW3FJa82qwYz
R5IuNagmumDkSqtb/VtqCItqSaM03QEYKWR3rxIBcSqtt7ibgrP340dFbadbQUZh
aMkrOjUuTDTloSbc4AntiN6jzzcMdefZZuE7pmJTeRdbpLjP2Q8DXbA8YMY+IQ4I
Ek1JSQfKE5I6c+XI41qVGSyBSNnbm7vdqVttf1Ut59Ktg51CM4T09Xt+uLC2h7HJ
qpBqM7NCbgmRhhgu+LhnDpCBrCGOiz5b9qKoBIkxYNJFQXOk2dxY0P9rFbCcmkcU
avLrgUIJ94imKvJD1/qig+9nkBG7btqbz8Q0qWQSZU5l0W6gnHiA3XGbPkBYgxKW
RJYg8KUdT6xnQvBX+JJ9eyQyPIDbHMYwqI+DUXQQFRgwv1mozKqPsCnvGs2Te6iY
VnnEYtLMoT5ZtN6H4RaTnaetWaVLC5QqrY/3OAWmrtcTbusBMyZqTIxaSPp0pZRB
Zx8vzbXoc+R7zXXLKII5kBIIKVFtxjG9sT1J7sHVq4NYAUHEvItwfQNjkq1gJrf5
jSuC9hM9g2o9B0A9pUnMPdNK7wQ5Y+0TCrRdln6oz7t8qpJtOLczqUuiXwGcoMXT
Hg1hUx4xbhGgrQNl15tEQCZ+OJBiIXz/qu42sWq9tKT4zAAz+ucU8oJtHuutFLvb
+/fuHndY1lJg/y8dUxTFzX4rPASW31Ye3mBSfNHB8IvYOym4VKjmbaS5eudXBdrv
6ypJsje1AwpjC3lsnEMGwY/y4Fs0vQY1wb4AVWMTFHUZnRDz4c7AgfeJeeY6IaRu
saYy8j5ocTvnSrDyssweBlLid01ORBWxUAy2B17ActsrZFZQq7e76Kk0vHHnyXRP
WejFApKAbD0Dhr3Auv/8z1h4x9L4PtC76ZjbCTkDBXzbrz7aCnM/mE/IOuk9LEDx
ifaMsR6XpUbdiVjs68Qi8I9kWZh43m5OWssYGrUK2LEa1VUMuJ/21XuD6fgOj6NT
uL+uHa3wrpEON2p9fRTGcn/GEQ372ASKuP8ddCID4pJwxZuLL/Lt7z/UGf+i1KWx
LM2xRIgGHiRZpiPJuklevy/GDbVWYeew6myU0PW00xNwtbHAaX5oyypW449RAu20
YZx2KT2ECuvHYd5xuHUvfLQygl/6CX9rAvAmPwVu2zFQA9p17FrjeUpuLZCGB5PA
4T0KkQ/yG64FP7PxtQCWpO1G0D7jOL2crLQWvFD2Q4AQydDh+imlFyYyXTxsnKEU
Fdl2cVt9Hpde5Rq6zsZIeLO2dtwZapigbDsllTWDaiOqhdceNuqt9Er7qS7dNf/m
yrrd4cStQmL80/b2JDii0ljfG2WXEq9OR1kUgZbxKlGO3Ws6ymFr9Jz0JYm6G3B8
zDvty/yCFbhIJ8BpyLwhFxphICoJcbjLUyYlCGi1EBLYhP0b4xkES3iGqcmc0v1o
vpwdQcdTfzundkh7tq/izFaNo/6GAnAxle+rxluuRoViLXykBZ9VBONElX6NyALE
7098yn1mq1NPb5okDyOAXLJkREZD3mLsCtJpT2U7WUZXh4F8zdAys2XAvCX0mmc9
xvJouA6FMy4jvhWklMpHEyBaFcExRu2IioHRagI8K5Cfom7FXpFutmIiLEgFdNaB
hOB/5uftfRh0dwpzI9TQkACv9h9WlAEd+5WjZulHuHERrGoqe/4YUDbPWlbD53oU
paOFX7dyzauc78BWz2/oyfkK+B9IUyqr5z6svMXIhgQ=
`protect END_PROTECTED
