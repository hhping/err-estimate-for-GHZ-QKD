`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1GoEKfevzccFotBaS3G8tSZ64qD6uSxwjx9CMI8skQ//V0Cw8RFcyD2JNF5wLzt8
HKKFXmet11hclBjt+Og4hq5xFP+vWdv7fmt6FoF7i3CsUQbOE37lL8HfXR8Yiub7
OWKUAgLHMl0U1tKAjYGUFOdet8aHfOl+k4cHOylZVnGrDpGBfFpeofrURv6MXTUJ
Zz4ZIB1QSaGHDi/yFZnHMsDoo7HB2tVNt4kfHUvY6PXqJVZtPe0H8+UF5gf6qPcG
C+t5xeDPTTurFDf3HbDP/iBvdCZmvsnCmkpnlXHofZ4IF5pLQGRNgTilk/YxGW1/
tDhvYCbao85o4l7zluSim3OJlxgCX77VPzMyVxVnoiJydSQHP3PdZdR6LSe1U/2h
dKvl3ut9G3Qi9YVtI7L/4ntvL39wIn1Kk8zpPJEa22ACKp0fp5MXTQ0a/9GRwGBH
J7tDK37k0F/G7FkEC/C3BKMfEF6HVHpbVKoQbJmw/azljsfHQr/7U8mYkQyvXmQq
3N/AHRxZHLHPodWSK8jlWdHzf1CHWanVUagh4xyuVNuEbBleTJ/pUo8L9ORbMvBw
tog/9h9YQfVYniUTsaQnjvOhSUVX2OIeYDkMzr85jbpsDSp4MYiWMB8DkZ8uwQoU
WUM+Itdg3MZut1NgZNLQGc3+gH235GKUe/Ft4ytMBBVWyjoEoGhuZrlJjn2TzwrI
BXhHQ0sLxLCpN7dwHlrhrhIliYUNpo3o8RSsGT3a0IFQ2SntVRxmCd4przb3cbJH
0J0RTfbvF0FhnUiAWCarUt3Xlus1AcnBgpsPnwpG1D2/nLshCNbr1qhdEkNrX1Sh
2wgEzmKnzTuNqA1xulPgFY75SR6TAimThGN/X72dLWk4gzV6KrtG52UVMN0gWGqR
Ej4Vp9u/IcmYdS1cbxyUD4kIKz8nFcyyYNLOrYRV6Mu/28DZzBLAXI415iBjl91i
KlY2OAdMDOL41lszhEK0kBxTaZS4Sa+67GVCl/p6EOz4Ad8UUIW4OVsTqzq6C4BU
AUTOMEwaJm5E9BDYBzNzR2sAta1pUFvtvvkiFk0iRuQ4N+r3l+zGVBZzHV/1AIg+
FehqHqEFU8r8GIBlYfsOhQseOZSX5fV2d78ij+rPEcx3qUlhzM41He+9uJjdYMlR
+ETjFF3sKMXjyIIbylGXDCZIJ3WXt/X/idSybSPIWco7B+POKGDCFbXNQwGgGVgX
jxkmTUM5gncS8RA5hKP5EeIaFn2t7izyw6A+5/bDOy5XbQcYoUsbX4PT1VJuicsa
S5nXkmGXBB+Rr+vBJwylzJ8Ll6wUMDfB/Iq8gijHHmVYk6TMOsPpx04mf0Mcm7Q6
y1BSxbdZqblLdb2+/GpZ3hj6+dltyIUAHz1Tpb6tRSLcKWbBD0ZoS/US4ihdhCG6
CauBFK68ouJrjqa6de9FFLOt+F6wXU6OawJcrgE5JPf3Y1LpK+PGSklxEC0GRqKJ
5S7CyslRmqXm9fHTgqCzd94YdKX6dG6/bAbU1HQbN7k=
`protect END_PROTECTED
