`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEHZTGqDhb9g+qm/QD9NFtpqrCZdxcNpCtfs9LTdD7Yu/7V4HEdcY/J3JOmYTwHu
BHnSTbXkT8ESZLiGqi+dhIsu7NAax43vwAEHNzGV5viAIHBXgY4i+f7ec9JGcQM5
35XDgJxRFHDH32Hs1hWiHje2WEUcsfYn+Em0p96rPz4W+9hmlI6KOntS0tXKY7Jg
4WbVWTv/XXYczfTGEaATqX7XE9bNx+6UIcDCSdCJnsRo/g+dYVC0wNzvKUILUwcn
WT/9WrD1IaCAk7MzCB55oS8iMYo2VMI84qoz/RteAmNa1LUPEBUV88R7e6/MSpM3
YK1ZU+CvwOt3Z2xLgfGywsHKHxTDwcLyXNu4qk1zbpaXx7U9Mbvb3nXw7TED1u63
6jBMemBIEr6cyaxU/A2LP2k7L8AwZx5gsiZ2EZ/lzrGiP9EfsiB8OvtZIfZ7pDpr
a+6baJ4votkV4yhs7Z6vEN9d5OJ8rj3kaFeUpf26iumYsU1g4E4Pbe8m1edJgTl0
6odEI9ek77N0Hruj6Dc4cOrvctWNqWuDOcml8a2x5NxmYMQC6fhVDjC4lz+Bfb8P
bqkPTE7bF+Fmxojl+uv3CpTSxa/GYwiz/BN5SmGLIrsbv36m7eOAuoTo+B7MlxLZ
9PLVscD3E/Gr6+hh8p4DGu6EFMT2zyt5+mCfIFegl4QjsjGau0wcAiTUrKzU9SvG
h9WeTrc6UpE9NUYMx/ob8Sy/3wmxxKv7emGXVcyR6RFmECa2RwB4E3BDFP00mSLa
4VnQKxz1AeUDVci99ni7dvMZvqCNPzwqSEXhW3zacKegcXau9OtSPIq5lq5yiW6N
gxleAA5eQdYZ1G1A8HNShdbARs4RGUbt6gaLC5GklbCRRMrvRqrAkw7i+TTUPDta
WRxK5AI8HK/Iz9yUaoMGm2OICSb9qt3NlR2lt9O/Dl87e3GIpL7BTNRraFN6i/HC
`protect END_PROTECTED
