`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zY3xYlCPPNihWMTWGIYkz+6QVZhyAVfrtTQsLjKT/IOVIU/IHzp2vp6wiWMNlt2O
9YY0UQ2m7BITzgWnXgiRz9iEh1JcIvF9M/Fsi2hmHJnS+abXSWQAcXYfOBye9EIP
a/bmX9Bmt44GMP6K5HlqBFo313dOoE4H3VfIB9C2aoksqi+gifbDGAw4NmcQsTxV
lwOv+ZGub4bRyWtRn4LnsBMMR59zmxatMQEohVxGVm9xZ+na1bCuquaZQpxXbo26
JG9abOXc4b5pM1JnDpVEViHBGfMsNVXcOBNb/A54DyP3R/ns4mLQXHzxCuV6/q1U
QG19uu3nGxb05xfg3chwg+HIyBIB67Ii4mXipcDNLaW03vm9RsYskU1OsHjMMey4
8RLJwzXkLuuxZREddc6VnXxle9ixRen76ykBeROEkdU0s35J50JHCeVK02pHb3Rk
k5sy1jwKvN9HdEHrcmEN9UCoaimRk+k6qCDNNJkS1GVaf4kE1ydAhsdxy17iVc4r
0OZloJpLmEbTRIT+TZ7h9TWCUWFaGiitc3rbBlaLKh026IkZU+rbcreVqqyBndCq
h47lFpIAVau90PvLCEEfT2fR3BC3iSX+EArJiBTPgJafp5ThKZtNpFNtK+M3QohG
NpJMMXuHva5UsFPuBAPtz0A57AfSZAv+GwlfwE0uQicXOtnRkXAlYZ5Au9KukBtx
PvYedILYkIWYGmgSqVtBXGmId7eLY7yPHD4im4lyA+i2yIGEuLMDhahJ1AWKEDqX
IKHcah01y/48oGlu5lc/7QMlPpAMlVUqRq36qQzwBv5ppKbuiZmqpZ8EtfSBSlOb
guEZnyES+TixKpi5M/ZhZxkffWLMbkcEmOaO8leCQS9kMyUlzEDL+MWZhheViJBG
j9p6rVFWOV/fTHbp/oDi90oU0s0nj5Zkf7CFkBOHZFMrFX1qTGim0f3QI3zJbkuN
JIicj77/QeAXWpyQgf8/+bG4ROtFitV5nL3pt1cXAj6jZ35bRR5ZZcNdOmEgumFc
zmyj6TVBZPBd6mXRXyzjll3RRgCw+Yo09pwMn64WSbeB36Y44d+sasJ9jOGZvhJn
jWy471TR6V6kiDqJcc/vWUQbNm/8qresL5lb2sN2qYnK5OCYCzKhAaN7BlPKhjAl
h2LB6Wk6i9MZK7PVQUv2FWBwORNW42MG/ryIwboxjOQeohQan59RQhIyjOv7DYCs
AzCyht5eyyAHL3mbYYYkBdMdaER4sLj9HhM6y6ZQgGqffY+e3jCW/n5yYFXCEgrp
RYeVVJemIzxlkzoG8BOuZ1A5L3/pLOWvRpzgVhwYtOLAok1Fr5aWBVI/BfuVYZUi
fyWnjR8q3D8qI5QydAM7ptnnSXFp8EWo+w8pwQj2TD98FCsVKf/s3l2qzP5H5C/Q
ouSWcVaL6GYdpgEeG+BArMQd0VdgwKx4HSvNw3+8ImlG0ffA0Kn/JuHOJfOScYgh
OS/w7SLVk21hj+cmfn5JL8JobKj3zXrW1KfvSZZ22Rv9wFZ9jNx3gUucSQzPHr1u
UAiRCJdVIiSy/fLqtcR2IRPn/OG6GQ9aAOoxmCfZ1KYHmKEJcKpzuXIbSzzJfgcO
co29ZugBOb094xeP7+J5hAxXxV3RptLwPpGERzSqpP8pV3tj50sMfdKd9Rkzl3OW
Hq8/QqrCQmoTMGk9+rozoDw46Rx3q4tqrSwJoXfTjt968lbUPdg8QKMiQ4w6K+JA
CWQhMVGdLboiEydPng6hypgi+QysuTSTdi5a9OkmLOOPdlaklnBdRZMu5ilObK+A
CGZNfFofjpy+GosSEKXw6PCxKVh+ggbv88pqGRUNL8u+yPOC5NqNH8sSxivBkwo+
kEta4GMrceYpgqS1kGItb6RxNWhHjtcR7NvVwXSpWQSqsXzxxijSAF1sIBW53gQH
CPTiuzG8sHjHyirCRoVA7yC8lzXDb/ZoNACJn3M9nR6IpMrWxRHLTgZfLIcsBShQ
pZjoBrfA+XjYT98C4AW7RdRr2Mnlpe9o2ADKrl+tVCmFkhMCloauyvEAJCKblUlb
N2zpIjU6aLyeEaMz264KX4OhiEZUb7DiSe3IsSs7E3Jbg9P1N4exhyC4FT8hTuV7
kQ2wNaj96ZZ/PLrJ0nnDxbUQmFkv8mk/EzJlYMo0AagnDqpikMQhqAwNyDy+T/K3
CW+Z8+vYhGDlXI9XPZEIs1ski9LryJIKoCWVKwEhmoNqIm+K9h+1YLf9IS813tom
s+rGPxyZW4zD6ohMwUW4T+6GpcIQXn54tqKxetqEcoEtMsue71RF0BDeXvUJYWIc
Alu77s/Evv3zN8ZS2tTEtgOohmkF6ziH5dcQkiT5L0t03HGdyQYiNZeaDVzm+Xf/
bhi06Px++7DWmTBcUUmLvGvxSmar1jCOKz5GRPN89nshM+bWp3eI8d/liL6EQSpL
8OVqb8hAqyz/68Lha8Z3bgI3sGeJooW+cBqbmcGQHNIGdy1+1dnIap3pIac/mL/U
HU7tV0RXc5Cg6kuYmARqaYV9j+F7EAKqkSehbrjeJXw2losNvPHvdFVBPOPddlH7
LHJGZJA64INFoWK/h9KSC6nlJa9W1cfGTvzbmfzBLGvI8VjDljCwT8J/K+MVT8XH
nFwVafSvDeB0c+thKu/7Ak8YkRhjxanv5haiGiPPUhyIarZEZempKe3grN5DiuD1
U5x0HP2BQgq4QAC6JklikOVGIoCKRqUWJbHSfS8ca7o6QDgjU0po4LBJGwUrFB4h
nnbD8v88jnSWokvVZnPMNKX+X6J11XpKC/XJ5SR7UnfaMFjvQcyAB+rTtyYJDgRg
fuXTSNhCkgdsrQ4CkzmHu/YYnSuJeV9jyUJU912IA4TKi7oVW0atYNhu25NIjcrJ
kZQtGhPo4D9gsBuiIDUU4nYlWMVW6rqAL9XcPwNODXUZ/Umd8DRzyOxmPSGm1Cp1
6CQWSf4jq/jZY4GoCrtFA47KIzeLkBlNwGeH8rMCnHRguOu9tGWERn3JouDPZlCt
B8VUbF2Yx0JxZBuERaTz/tuhPcXVGXfu83xWgHEyKmarna+UtxAKeD8ZEdb9v4VP
pFa8JFtI3Z9cMQZu2VnM60UURc7OREbr6NxoQcfWnpXSAb6hk+Mw+0FLXbiZL8Rp
gPYodyKTxcveInHclmf40zG5Qi/iawM58k4ioIx2Ezdw/VvN+sPymQA0rJLNuDlI
tjPFRBTjMXz1X0n7+dMokhJK57Hqo1OKxVK1GUABcyPt30arsiWLk6rTLW79Hlwm
LvIFdJ29oLwllbbk/zxdwjHNaMr0eJMtw0fnboM3USumTiS0lKRXsBPai1Rz5ttA
qQW4WZtTKa++0Nsavlao7mXvHHikNSXyxdFt6OwqnOJhRwZyjTOm/H7Clrf/N16v
yF5v+cRCBzvcZpyP0H4jGrxO9XJMe+Uoe9aDsWtk9MHlT2utjoRmWy+PGrPXRwnm
lE0JpCcik6vZ7Ya6HXmBAb6+ByRLrACWzmkFR37ic1DV93TfX8/vkzLRax+qT2ol
N2bcSTXmGlhWEWVwdG/hoblVLH0JsoxbQp8aYfmZ5FF+5l78puQGuoqQ6aVvt1Wa
RflPY47cBnxmqf/do5esSVY3KJrrOakLr23YPpH3hjAriSawAsxF2CSDQ39ult3N
XrgkwDSZK2gf4Lcw57uLQh24Kny1b7LgIKLtf3Lp19tsKOVCH0yDCiHo3c5INkGP
O4Zt2Va9OKXUpnWpgp7Kch3gkLgz+qGMsWkZQTuSJfKtGWetxtGWCKj5nZ3JI4eY
mkNJjLEJdxFCY/2+3m/+Sw==
`protect END_PROTECTED
