`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMvuMtHfsllQ8xanVkJWib0jxbrhCkMv7sLYt+AV40Nxn7EP7fSbVhSISDWB/3DF
U01LkZf7bK6K3YLg/96zEQg2yKZAovlemHdbDEYEmvK4Mmi0XCHa2f8hpr288UYQ
2Fo5yQEjWAnrsnD57FNteXb46mKcXuGwK7cFxPs2RHo545voEfor6FUYEldmq7yj
B95QO/9RhhepPTCAKk1O5MgclDn+VO2kfuWanDGyp6kfjBK1W2jIHW1RDS0vrkdO
PSKtHrRz8IHpkhnWQ+jypFD595xo4qmKALXV3equKjL7OiGfmvYBqzjrZePtTqAQ
stU7F+deoDh+OWi41YHOcJp4iKpfDFow2qGxCdTjQjI3ZXWA5uZ22PC7mYxsIe7I
jpqVPjPE5iszXNRecwUy+s3Bt16L0XgGZELKNvTn3YOhC98jFqYBAENKHae0HXXj
AeiFeLnYm9kKhwv4htj28KyXy5q5eEmoHQ2S3sV5IVf2r9CF70CzkoULs21KvMZM
ExcHVXTLBL6AF4C7OOWxZwgFIH3netvU2Uf7ODkslDEiP/QIKwCOjkhFNkG3rMf5
nbt4OHh5ci0bgCsHmNXhWzoHc4BxGOsKwdeBXTb49OMvCfI6CFousoJbww3ppbc7
2Pr2M9Xg4u1rBPa2+YovoiVT5c9Tgfg+9g52r/YeD5sXR46sKyraYH+n9LyoIHMv
cK5kF36jO4+as+0RvTruxNQ+s8bZhOZxy1QlTnIkQOABsVymUB9QbEzcWUTUg+OK
9O/aXyX8UzR6Sp5dsPYhxeMLAe2sWsrdQpT1l5XrW3mF2IDPSvKhBlr6e6+yV1cC
68Cp9kc80X6NPQC/aFTgoBN9aJ1SdIOodWIl41T40xqSQyYRZ+CBj+0vqZ69ueiD
ohq0aQSdzurCv6C8zTdfXQyyW1WwxeoHENNYO+Wr3IL7ZMZfmN1wvvfA4BGsk4o5
mYNep9EJGYYuScsgU1vnR+kN9iwmUhU2luPmGfRLdlwNBKOf1t+OEysDB8YbpQeu
fVeitNZ2M/Di4WX3NltZBvXDVTwn7QwNd9IJwICuOzQViu1EQNMTIv7AP6rYMGzL
zILz3yc+rfpuyOSXBKx/5KVEOLiD/HKdkaVs+Bfby84wkPGPv2uJodspBTavngo/
gOwRIo1cmma5vAXR8JelezXGsqmyKgelGwR8IbVuUq3nXU2SvEjKmkuDknudqeer
xAFDNRzccegg0Akjb/RxpHdIClaOHkgbYa9WQu35WxyFYAUCUbxDL/qgmkuIB6CV
3fh/t9A/hZLXaX3eE5QpVabbHH0JPNHc3+eHOGaQONzTdhiAbzY40oGCzLBmF1xf
DDyJmfvq+VVwLfXN8Z7U1D55p5NCAeOx2CQwy2eKLPbx4z9YwZ/90qEvypSOJkaI
e0mlzGtfsZN2dB0pWecKr5uxOD4YeKn4CkFUoqlS1wYhJ0rcHLAWz7/5PjIS7Y/Z
cs7Di2pGb4+mJq+WtZQKDZF3fh+keXm0HWq0H61XMHJC9qOyk2tBKgAMBdiu9RBf
19ZwzKY89iEohkroQv3IFGud3ds/Me4aDrCP5y3m1oK/e++3gV5Ea3f7EfahZ5xi
jDBMksHH1YErlvqr9bF3hB2cJmPWZjXNNjfepTub6e1Nzj2C8slnqAB235/XxXUA
X8A8XyqF5+ZlHFC30mddkpVTpJnPVKtCeaH7scegxUXsbisu8gvBBIfyb9GJRdag
We2NupvGXJjnn/Zc00emal+RuwsO4iwWQhHu3nrbqEn4Qg9YQA/WbGejmbz0leXh
3mmzjvnrTysz27/FP8Cq/tMsucrbAqXGxr+OhWJJ3Qh563J3biNEi0mTMmVK/h4C
TiwgYHV/5JctyvbZWYB+9lEQTam2JyKHJayperxsbZxTmDUAjUV9pjeIgXI+NF6U
uQK29ztIyXMmSqFu3FcLUm/s1qMiYGl2a8hrPi97FkQWX/9t4WE8oJPlXFAr/yN9
OXxVvSWXN5csRlhZbLp4dUfPe1e8P+GF7o7bVH2aMlPSf6Gdy9osD7OGtHwkZo3/
4dudpPRaZI2tygMlVfj0/1aJYAFfKpGC2QTLdygcwhOr2zogacVT/51Kzd/ZQk0C
864dN70MgLQBp/+n6Ei27KaJttd3xwe/S+cbfbE56Jf8q1KxzBnQgHZPEI3NhxOE
xdstI8aSIvg7bSNGGnpWqQjitDIuALXcco3UU3bQlQA6K8KDaxM9uglpSyTnFnCD
mX1b47HhYwjF4R3yaDh8/PRLluqyUZwj+i8lDOXHS62Yd0UyHZQbTGVhym9eA2Y/
zOq290+V3TvJrhhs21ullmdEVuQnWRLWHFsPCagyk8rsbSICPZB8WvgZDtG/AQwZ
LIzalzOxL11we2H155IVgXY9It7EuVRKLTx+izDg1nyZ70i+/XecZz4a0HPhejue
LfeWDV+63o0WpLZN+DLcSrWYk5TkR22cR0WPSSOY9ffyVBz7EYK259O5uF2OvTzt
2POoJvioq0vzhbu9qsedGwv+NK/dpEyYpWcdYs11WD3DMuKQ4OjEPxBthtI0v/Gw
zT1STcrK6TRsVDCsdbB0NzdDRhwvmTrgvzZp1BEH8nqYMY6pwHmZ4SN3n5RmYiGM
8fbE8XX+Nk7kfvNd/vHrBdCpc4uHn6qBGO5W9GKfV3Cnh19wPpMPep4QyYSL7PKp
3XJKZnNjc7grVubsHv22+TO4gz2HJ2x+Qhr4fUo9oeysXYMBnSzRfkwpAJVNr6OY
GXShBTmghVJKzWb65t8X1GzTTLX1g1QwXoqckgl7GwHYmtZw9bJxHYbkLr4/tp5d
DKUxiFZf5A/UpdYhqjojuey9RNoQvcae5gX7iKyT/FHhgqGz0Ef291npVpQu0tK0
ibj+GlxBa79p4XUCPuE8m0NbOcCdxNO3mr9AfUDYF7m69gG0uyE2+skk17xuJgYb
oIAUmiLWLkiITZ5gDmPGnxNBejx+j05rKghjC1xtpxNTQKe7qCrz5WtqKqBNnQ7F
dd4fNiG/NBxfaJSbtfRLU4W/junzp0pFdWPotYhtmzZCKhIoyQZYb+1/iJBqmWpT
piZYEmyfxM+TWroYKA5FLBPxLthAgEpfYpqgI5+PQJT/+BiHzqWGPOj53h1qy9ni
gwYCKcJWR3bKoTHhec1uescq3WBirLPTeYXzfM0tcl4=
`protect END_PROTECTED
