`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlOCfWc4b91fVdDa0zAXlP1J3nfu0yadg9cgrvceiMEEYWsgKpJczliJZWMoidpr
Fdrk2AZ9X2T6tWyzZm6rkL9SFBCrGou7abAciaqvnOrjz8iHqiv05RxcujC7AUF+
r17SB+RNCs2u3Owjg5suCT+IJnH6v6732jQW/jLQ5iaSFd/M7shvpsou2RZwcdbt
U+OnMX1IqpJ7SEKny7hKic1O5MFoOoXqoktL8y/QtSO09gEPMBeiEXQUScY2n9RY
X1vToBUAHByYYVb5/J9KYPhsN3P4dir5QG1fDT0rJUNdxuJEPsmX6RQ0raHlL7Vc
8XPycqhh6A/8H8l1fd5feadWisq6326cLk3bYF28O+4HxbIlUnarB50PoP3AH+PK
TAY1nSEj70X9357DIePCtGcLZ3rHcxX28ITW1JYZf2YeGt/wF869OWuqAEAdR31E
6Gis9H50TDEbmq/OSbXnZUBcfLj0mYo1RfsQZhhOqn7Jx4a7/7wlswNm6qMLZCKA
nLUkD3PTVB9MbSirArAytr2cEc+NBlf81xCH2+B/4b8lJaroMZevjjhqSL358CSP
m51G3qGsFJXkIHNP/4V3PrA8jMs8GZczCRrpyrLSLOZQkxabAMYXst3dej+A5jPX
8TPCsLuUTPRCVX+RhqaF7hMgTd9tpu0EGWAWnvoV5Q0=
`protect END_PROTECTED
