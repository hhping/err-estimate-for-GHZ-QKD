`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDqsoEcWAEteuWWd1sRS/YNv+XMeg78lReOIcdSFsTTR4ah1ajs+gVdQjCWfO2TD
lkpgQFp4BbyX0QJMpGEWhTGHRmllpQ69S9Wmx5362wnVKyYX20nIorFLCBprVTml
GDcP28i/1BZ3cQUYi374EDOdLcLUfI1qrd37Msp98OBWMGXHLRlC8Vxb0CQCaPtl
dIrTNwzs5YgvDKgq1sPgRad3q6eu1SAOgviAON8qaX2YK8SFE3uSmu+5w/KSMNQK
IPb7oyYW2P4nzJlnzpu/dzy79nBrmLq0mMLNTVUieOeXbFBnjN1BhltoW5u9INac
q7OUJ0+JCpu/+CW3Cwf2RHBYFQdW+lazo+PQrghThIZ3GYPQdD3Guot6w3P9gQvC
YRh55ku/qIDYffa7WsqiivEDQzDuQEH5WhSrZnms7aGFwgiHm/fL0q5mufvgfQ7A
5dvcdoBrpUrMUQ7HcXw17UpVTULvh3CKh9foNtlBE7clpzDsU+irrHq8M744s7ic
CGm4hSTLfbNtanbyueCHUrG5ngBxukITP6sjstUVqH7t4/TCqI6ftOnhwJf/nVnP
H7lrYBq3Za+PyXuqZgeiLqyjO3V4A7fnPDzOo6Xw8UdxdBBxxfIxIlDd8EaNc7gP
w66eXZ5isgQq41SFf1VYKl7c/q3pBOhhb0IGx5sUC7Aec1jeSTMbkjSnvzpyEJR7
7WgYk7Agik3X76tTKeI0RL4VJrU6JoEEvKurzukh1jp5cSnUbaHbYNEMv/o5XkQe
bTHAWxU1qhOEu4I2oLwHzjnCkcvYO7sGn77fN7jtHMLQWU6NWkM8VIY1p5dUgOyW
x8k7V3031AdOQSDJnoispYusj7jwMlqHliFqZHC8rRsJee22oIBYDujnowd0hdCp
OJcDIfmhI/XWTrxIAQK6hsscYC+Ri1LIzRHH6RnEL/ET0DxzKNzn+3CUTla02xxv
DnJaTICvx6ggGH5yUf4pYHUTZVWup4D/0azs7VajD4R4Mu7kl+ifl+9jMXJOkHOK
FznEXMZINPvYqTuAnlezvEOQXO0dhp91LkCfxXWKjt9hYd/9Xa8ZFnmNu16dn7ou
erB1DsmQ33t6ZJ5Yph6RBPLEvl7d8uEEMpTBUnKtsbz+xWydB7wrxGUdCFhzjzk8
Jhyrwp+LLaRvAq+kX0PtoNR6lDOd6FEsptElkLWf+L/Ry/YLkaW2+1VBlnNQrVSq
IK6huSXtD6CO2MmOl4ropfXuDFgW8LqzHAnlofvPG34767GwSQL34qFNtqkz9CVT
+HYl73pHXHLuyEG2lkWrX4DGtNEgWjf7TQr0+c+yMGUFDh2kNQyX5urpQp/vJBq9
2rkyeS+xvNSHhBMWTnhJVTibx0iaJ9C1NwssXbFE3mFLvRoC1oc3EXBzIC3IVomD
QXdW/2C5AVPmmsf9G4I0iOwAkIQmRx+ezoG09eBtgP2Z80W6aNaRfI6cNWrWTVVb
e84JI3to6WqmjTGIGFTWggW9BNutsaHvTWToN7Titc1vKw8cHX3XP2aOjV1OyrQ/
QHQyy9vIXbARd4LXuECXf7JM8v9xC13T69Wi5nBObD4ArqhnBlJeTNmqjJQ1DXsD
hNJZkkO2ToH/hGy0XUdBjIkAmd9vNdlaM2JnTxxYqigTPy1yPMGJHOEpB5qBG5ZH
e7RAAKd9YWxuiTACxdux+/ZE6y22LasDNic42giQi1hMYnZuP7aqp7FsEAarUhzb
MvQSkHU/wifX/ujXhuM5YbnNKybB4MCqdwMWOAoLkqHuzsOjLHDLxWZgvSUN4cET
ZBsL1ZvFzobKlRb7o+9LavAQTcBsTZW6gHtxk7mpLeSvbO4SRFCanYWtiz41WYAF
Aiqg5mB+2lzqdut/louAa2jRgDlmlTAL5lqpgcqYVC6g3HZLCRYtD1lsOHgx4rES
7UvOSjnVE7Xt6vjbjNtYKEbIeYuIWXe3kISx9hI9UxpXLbZExDi/V6xo+FKaeZGb
03r0CHGr1YnpQTdqpJQmE2ntx8JNjJsrbYooL8w5qaIiHjxbzorZMGqBi7qj8Ogd
p9txSfhzq16wrn2GuhEIcOODwLWuSVb3/n7Y6J3QjZXOuRAQouqBEsh/Za8tSYkR
tduGRifi2FxOg/e2OXdZJzTLPvUotgDz3lgr0bu8zrSZ8vcRkeG6Ii7K3XxAzn7u
wFx8SqycdOQe6wNG4DPYIk3S5/sg5BoBem4OckDTJXjqXFS8cy+2rjf/462XVGBN
N1xRUA5yvezimQ4NgUDrDpdpG1ViuVbBCe2w3EHR3DmRDXL+ABT5oPPBWb9a5rBu
lUe3WhPR9adCNnke9RRzB4pGsvdJo9tIWDhsyDhh2lmSLj7XFbskK8/ACNMTY2f5
WDLrvuPxGcd7PQBYTy9QO/jPiF0UCxMxLu5oCfse2Ma76tNLVrFfj0cKErsFEzBy
9sUiM1mUZFAGVykSzjMB6eJ8C8yrUXFM63ZSIOq5RkqAKDdjekodq8uV/o7PkwFG
PDVasIefJrWYsy50h5ZK1NBgtFTzKom5lWbfYXM30bh6n+02EAThk/of1bBV/eYp
T2mwFczBse4a9rcSJ/Cbw/pWnDyT7++bVytgbtj3TFhkGWJfzadT2K9P7WDUK7AL
nCvO62JewclvkedBuqk6rwzi55Wvr7t5YCNcwiMOMgaex5HJqcvH6Lc5aDY565fq
7scZSpogotjend73IuJQJqJKseo4fLH2E9gEifGg0W5TMeahrmViZG5oioVD4R2I
bz9N3GxtRcZXuG0QIfodvDkKU7qRu2NKUgeltzJVgf8ElTn6TwmyjdIvMFpvlcyX
qAXQwrEXSy1dFc85oNUgoi3I6ke59XJ3fE3Im4o/jeqNLJwh/r6RtASXz05ZIvyR
zw57Fl+9yRFVEEuwimx2fWkR5RGyPqILyjbD89MTI/Z8IWMFPAnKD7hyRzTwWLhn
5jB9JoWe/HP96gdcji+73UccMW/yyQN6xQd99LOm75M=
`protect END_PROTECTED
