`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpGwnDQlQ4xiPsSXvDzvwQxcO75A6OY1/lL2nkkqWNnIyeABj7Y0FGkkq95zhe1P
hDamjGX4kKqep3RAblWzVpcTcUV1S3t90fXjicnvdKqtotFheFt4ZeggKJcj45gv
cV28xipTDtt+laNGIO7RhdF334vIBmDO4VrBpiQHamvxt9tytngfCMQUCKrD0z4S
Tb09TE+qebTNClwlF8/GyIe/SNXy06TJciZeTaBP4YmFHo4XQ3tsTcBBwH2nifku
4L9lPhz4fNpS5iBz5LH1jJzwEduTMJHldohVk8dMJEdi9yXM4OZb36DhRfKfHrAZ
8eyuB865Oc4S+v3RCrPotBdZm52ppFclYqoYJEwIYM/OS4VC5+ZbH3RE6eOv74td
AprrOIjh4NGnjq6/ZC4KdwNwv+UFQmicDrK/Vm7kcuXCPq2A8OHGB/gzXmu+jLsT
vUZRrtiReKQV5TajyI7ZeV1jEbE89eFQMww7w4L5vw4Lcz780/LSIyrBkmcQEWh5
FvvU+ZpDOuhnaWwAT7pfM5du2sZODYCZ+n72nfGQUP5r2847WxYIWX4Sqyix+9ME
ttn+L+hMPRZsWwjqW7nM3V2AbXvPx5EWxplQWu9rqjTgIgn44tIlQ17X8NEEEepi
ZtwPXdUZO757wVyD3dlxuTfk4nQDonISUqTSacQJr+mmaW5PAsRW0Bw17EBkZ/h0
ZxlYRlP7AqjM5PJNJDvDUFgT0iN7YWMIVI4Uau9xKY0uMmw2qN7/C4VwfZYiQ5qb
miYVptCieYAInclDtMomanFnRKw1u+8PZxDvlfMHtmwhTgAaRAE92R3pBv1+hlbg
271oHcqibOjWHO/2eheAUkTrhhPaYvC25ZHurWqirQXpceBu1qjXQxHGVSzf8ZGy
1Lbas/zgxg9sLwJMxCljV1vVbgChDTDBzPtoCketoVk7GQMCMnVDa7DdyF2pC/jr
/Ej7lEgfkufC/QbGBZqRVYLU8FygAPQznVAqDVvLUOwHhBA+0aBN/p/L+4ajw1IV
HM/3f9OWrfipy2dd5EGZOGcFDNzOX4VR//Chsieog7pvzISi8Q9yOIYrJXhP6I5r
mpbKeAeXZzhdpdpw2puz6Mmv/O47/u+e8nbw2xxD2E/S1tE3mgKPBmn0GBZIUaNZ
`protect END_PROTECTED
