`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+ldUtZimhXWUFw0729PbtmxB+W/DLj2uxa70oIFIrviF6UPHvHS6XEVsZfWOX3W
9vYVV3/m4tZwvz60vPmGs5/QdwyXIf2YTyI9qQDNedadvKJF5JQD7YluWwSRUo5H
g6ZoDZRQg4iRVkmiskVeHq07zu2R99IpllaYj5QZnRvZZM0LrKLd6aDHiJkRRxV3
BYXzDqEJX6nH7H2Au12jm3KS2IfpLqRQkk8s5VQiBDsJnM+uH2ouAPUHH3x1oyqK
a9N6WBtT01FIV0baEYxWJRn9eOdnS2CLdzQlwZeJeZJ0/9CbhUWO0Hvo0x/6Evau
PmuqG0cwUwDRH1l2mV6FXt5LzF7QbC67nW6kov2Rq26V1MXPUZvROq1MvYmvABPv
IlTN4dAyiwJyYiU8Ic8j5VR1h8drDCvdTzHmkTaE+P2ZFEWi/s3gL39dkeBcPjd7
pkgfEdfXsac9jBiru2X2CM50jp/kdqMA5k62LOwmoD2K6kBJLdIN30AEmrW/IDVl
RVnE7y1B4YbcyhyPusZVLrDQ1XO6PC9/ceskU+TCWtimTHJkG4zNg5laj2FJX+1J
QjlhIIHgi+Co1Hq/v8uu41p+wHyVjICXwK3QDc04BU93ccCS5v2+D4C0qKfmCelG
z6Olm1qFc3lLv9iaNJAnf1O1jyTTupQt4pbIYL1UZ9dS1ORdZrqgo/AbgCePJ/5Z
hRYa5hN+oiQDqTA8SksPzVUi+cycRE7bVL9jcvZmgdE8EAhDVZ1KvPZPNR9zT58C
XrKlUBQ/Zbj/ju3KDRArP7rPrRHlk9AV7MT+h9PDGfgA6KsQkdKSVCeABJxG8SEZ
pn0h/s6t18K7dvzJ2SKgh+0K5uIvOHGvfsxFfrah6QY1fdok/VgPshrqLURrtbcX
fXR0tTbttytrV3h6mgkDDB5mbf5pSgqcboqrnry4QHqMWKnOdQ4GTrKNNIeEx/M9
mi35s9HDBRQ+zEewIuaYUVbU99XyryQ44vg4Od3/XNKC5wySKXROh8SYIlh6hYp6
tIdPfdF3JHfEpN2KFBNIJAAYuSmepQB3CHyyDw/2S9Aj+PYKP+Jb/upsPD4D7bQM
lgRrBITciYgE/BVPXV6j16sH0/jKVxJOXSt3jVtrONG+M3bJFSffjNSsozbVNU4p
hzW+X1QtGQ6N5QJYr3c0mtPNJd30dspCmOGXgp5nj0d/5O87hFueMOAepeUugD9m
FduY3hPvGYB0+6MvtoZflW1/HWyPu1Cf2n9G8ju8JQsPJguZJvoPcOZQjcBg4TOA
DcvrjVrt57koGrwN6GU6J1tDbBEFFupQQHsfHT7Yyt5isoSylm9QxDhWzLXBRrzJ
7r2dKXRbHZnj4We3XkX4+GPvaB5z3f51K+JvvMyQhrFDfjORfujNQnJPIol88qv/
QS14XtSTc6fmr7FRbCsNLmY5ntHtmn5BTyD3W9qYcayod9HVXkASiEoCw0nokr4y
/X/sKTWrNNFlqDbbOr2raTPrDYEOPRE/QRINGNgU4au5j1DqQtNnegux6211Q3/J
ZsZ93m+blEj3tsZIBgwb3ebd+lUruOJTjIoBsUUULWmkxHPGMZLSsEFepDLC7ojR
rc1YD7dOmf+F4+yhKKAEoLCasJ73WDU/YLOs4l1KZgMv+R6wROHeuAScFLZuWmym
rSSSOPTDztUoPVX3rl0uphd56+OFQVRlV67N1+2fGzfm+dxzF/Np8lAigBfySzT1
GO3LM3+nnM70g2+qQ5dj5je6cA/6TFRceFCggTLfN4I=
`protect END_PROTECTED
