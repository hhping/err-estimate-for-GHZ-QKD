`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxXTprZXE4PKyX8VoRlAnYktjgdv3jSyYnqkMQk6LeUO5juHMUE5OqAForrKXveW
ZDEgsQ9Dtg9lQ/tUCsoq+BMwD2fjLVgsXaTGv5eggtqiGBuIU71UTuuW85NMC4na
i37Yjn7grzTvLtKW4ICu4GnMeY1NFHUOHHYDSSShdINFgjSrWneDuWiH1xgv7t/b
dzwj41k0HXMCCvVqR8yOUT6MwtGLbiSo4OqnDHW9GxPJl4WRzLhuY76zeW0+93yO
zecLCTyXyMQajEb/AUx76vJTyqsQPp+Ry9vqEVm0m/kUtJvXI/6towuiy5IaXdPP
/R0ESaTG4xK6SGZch2AWH+i0sIP+jxLTJzTff8w0ndzUW1Iie76bqMuaDJ27IsXx
0LluBDiLkPO8WAozpxz9F/U+ZqXS1scsa8u350tyx7RsuVb09SHz2OW63A/7CfG6
p/MHYDxaLnnco7yZ9KtV1ndTvV4244bKxSIKM0AzM5/awHcfvVFGxeOBjNd0td5E
EsNil40XOGQs6Ir9awtDtgVy4pA3JA1DtiAY6QnXTsy99z68dFErrLc03uWA3DtN
2HRDu+7nqWWZUMZ4kmaM7cv08noibP9EnaUrJL6LyK57SvIURkbmvE02vp7bLlC4
UQ/svO4gFw20LBn/j+1peWJRSjJ8iIyUFkuA19KJl4gUhInpGMQdVHuKKSEVkY1h
WMY0w5JitgxWyYOsoT1SIDghXqJJX10p/QtEmF/qSJ7ZypB31Ls/GNC9iYlez3VB
wwkDwn/cP/w4hjufoWTnL3wdcrKxC6Lzp9HT8I2Wfc3QIkK42LiqXDPxBh10x1VL
1pzNr/ngarVeA+YYp3/YlI2AFuQSaDsIFlk4zvqnfOpkUWbOuUGQgVzAZYKZU8+G
5MO8qj8gW9GWFeGu/WM4VqjWNVhRJ0jxTetElEWyovkyxc1qWZ+penHCVudlXNJl
SQT2w2SNXgcek1xrvVEZS9p/XYfQ6iYilmrkoUZFhyxD5cobSqj4lbr5KeVIHCRy
RzuVlqotfEaHXlVJMaySNJPkWA+7o1flXxi6tGt/doHVzRlo2OcYuEEY9HTgncQL
YswvawlcaLaid3HdWAuDhtq5azcO0MroKsKZVx6njRhV8wu0GVJXUtHiRTG9u3EY
EXGsVwsVNRVwPEa4CFTV5xf8nkq+wUfdjdawv6Fdy6wGCtDKz+u9Na0PM4q51ZE2
Q348jzC1Hl+uOy+pxVy6CQ+Nhb0YoH6FPvTCjqlMPuY3S59UWW0LT7igjtVP5Wcr
VmtsEwgoxC3LoLKJm6057Q==
`protect END_PROTECTED
