`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAAlMPe6CrCCLyc5keQHnEka3oMmLVk8T/hztYkbA1mxohi9UldoNUdY/yZM5lax
qWhon5S2qdG2QqOdKXhU3cMlRCbDTfCdLe4tqZQBCiINFcarM8cl/R/yeM4vcfKG
Sq31SyTBbFW0/XRtIjTTWkPYvfGu1jJmQFnzix86ZCMeFk6BfNUoJwj3s3jzcfbd
uewGVOCashIqC/L7pIHD8LYkAhID4E9W7kwGHIpaV28QfCJzsILNpenjaM/x+jlb
7xEw6LyJhLdIV1W7NeU/VvzDS29YXreUJk3SOc8GR7uGcDr5XHXddl21IhObKkut
25TvRwd5b2gbdMEsxB3LaQ==
`protect END_PROTECTED
