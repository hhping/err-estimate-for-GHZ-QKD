`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWOD7lDEdC/4etfHCn7VQ3subVyHA/i/GbZWraipPWyznnxoj9CsDE8hAlD/B53g
PdNeoE8QQi7USLUUrw3kYKS3fTNinjC4wTrqzURxHFtZX8xl95Toj9fNfozrKVBZ
kF7VIkXrykcKlapJ3tCHRiipJ+NzvMDNakTt3ut6kdbb3fv5/W/Qc5c4Ns6pDHjM
/zGNJuWlV/6C1/WRABFwBrGSRVypYs0dM7pi0OnhRFKVaKsRNEdKLiSdbc3RR2YL
umEzJp12zdBd87vDVgGroKHlq3QoWY8qFmU37Mb0FcntSmN7FHw0bQzSJW2NsOdA
p4ij0kOvo7sPcQUDCTVTHQYSEJLyZa6PzKqGo8RIZvysNkZMkzJfbO6XCMoSfu0Z
rcobk+RzQ55PBcg//h4B01P0CW36VbM3ib1tSFGxIQraNjiYbs18kQvNVAB9lp/0
QKmETgoTZ17dlN/mZXiz6A==
`protect END_PROTECTED
