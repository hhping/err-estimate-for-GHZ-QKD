`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hsCGXICjQkWxuoPkyUdms3Qhwl4sKczSLk9AozLb/i5PsBVTuKWENrDAZ7KsEZc
vJQjGaIKolPPR+uke01ioST3F5JGktszhJIQ157fcahWbxRkfLxqxSSTUTtJOE1d
AKQsXqaBOe34FUd0WDPDe120ajK6rG6ZgEY2LSdOGPb2RZ70jXSf5qrMbla5g2dJ
Yfq0xBC+uC/wMwUZB1oZTU2J6Dxo95G5wIA6sp8gUORiAJe1cJhor+ZyUxEbVBCA
VjPd8U5o7oFkwtr7033zmZw8r/y0rIATSK4vdJw6YP8YJkJLzxFhvdol6QXa/pSq
/AF34EJ2YBCjj5vHHPltCdz2aBeGSSpxcy2dWOKjaqVwIkOVkwi1vAQsyaCaERyP
blYjdZMOybQXz7I+cerEGESVjOsCVI/jf7DDmdkqDCMDi6439TSdvR9/fBmq7I/e
y1HFVlIqq/mEGUkArLzn6OruPDJ5r8S4f7hOBl/wLiGWpQykggZhsZEglR8jeele
zzazCcgiTUkHLAAkvSM9vX62u565hiz1d9wHWMm5O598WfgvZnqcsJy1xWbFlCAH
xP/OGJrfvNDCUii7AZ4CJSDW5PIAIfRGrBw+D4Kva6I7dkcrZbPOWcYg4t3FeHI9
ywht5xHQVkK253IENlT/7TirxkQXr2IHbNjOuHRbM127D9EXNW1Bxv/2j6nvajcK
1bJgykSFw6J8NMObN2tt6C9kBKc3jKzHN/trrvxtGj92hupeqGf6gMhnVDq7ZCMK
`protect END_PROTECTED
