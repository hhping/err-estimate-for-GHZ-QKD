`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+8nBiPaJcp5aK09vCPzmsNQh4c6JRerASjoEklxuQmqtBwMAHQF8W4739qxDSRpF
/lXDnlRWlUKYT/3cr3Sr0f3J/cU72l7/aE2fBvyYc5tHi9oNyW+A8XHX5APV3kha
0M0V40Sd3Iy55om1UxvliQo6yhEJgCiFZxqg1VeoiUTZ6wMmwPCGjlajF1hl6/ww
V3obb5g63e//WZovWAPVClq9/9uad6YELarmp1rQL+FuFYJJRriyJZUBMZMEsKwm
2OT3Fe7TvC0GPpCPNRaxYAc6J7tZt2uhFH8mWbENj2/w6DUMkwbDvCbeY3nBC8LG
Pk5BXcSso1mDz/hw6mHkmMxxb4W7KmnJALqrsRTngSA2By8pWtsaog0YLaWBDiH+
7GFmj9O+7RFq5k/VgFcC91u4u73zBxf4yorehHDHAybUcrmbIi4wxjqaIQfURJD3
zlBMlZZSDVqCzFcGs1YFlHNPIDpA1kVpo17qIwS8Dou0bjvJmci699X5jM+1AD8C
OCdYnd2DF5OebJ62jMNWDgjTm6sfXPZ+WEwwJHe83auUt34SwFczy9hwGuWWJ3Sr
R6uS9gSmfBWX47miemaaJ5GZXGFQZIAdC4S/ibJeVBhyybeJShAtICvG3wF/UA66
n/SkgTb4jAW1xOvbZNGjyNtsFoxq/31TB4VJTCawE1L5Fp52V8OU3mQV2RLqx0Ch
I9icmz0ZtZoDUteKFKYzVt+GJCxpaqGWDNb06hhR2zkaWD3pp6bUTF1OuidRAKxH
Z/K0W3VEM/IrpO7reUbuxcNq83LuhqsshKhuM4wgJB7XiWg5C+c7FBx2kKtLMUTU
Psvs32312j1aC0Ed7Or6YqA3iN/v9RutDLtjdjJAcbb82SXIs6m6j8l/h+HPGlC2
NWVYkzGaV4nIeUEHnIiaZuH764nW7NRVJpCCkN4/7mQvs7OSN2SKqGijZj1cIwKN
rwM8wqj+6K3bMhZIORxczCUY5mUz2PfD7VpBKKznFYzwY6ThSlDspScmtWPB++C/
DQe2TC2iGMnCzh5wA4uf7lnNJNkMIantwdtbfFR/E9tXVMwfs2c8lxR+vMKDLO8Z
4Kbhuc7cGUZ0fEeo50uYiHq+8J/Em0thfv0FG/5/pw8UHO/m1JBqFS6OEhPvNOY7
u5Ssgn8vb9Iy/qZFWrPKuG8hYCzwW5cvipNIsFzN6GlJRC8VSlk9OUfhcVeJFqsu
JMlsNQ+0t+tirYRN6UZqdVg82jYGvHQM11mHomEVUVGtLaXBWy0zHMEBjYdtErFg
sQK2UycOSqe/d7hdjUfNHjsJFmHKyLv+yi/xCIa5oJZHaU0VUWWEHuoLKzGeKSkj
uirBTQTquwj59ZdWQTjaVA301CM9aXhQuflV68/3RUCxZs2zXwrsjnJq9VZ4a/xD
6P8/cVCd1nLX90GDWd1eT/K/ja+MHdgwK8PNxkCS/bYXyqsKgir6zeDVFuAx94iT
QJIeXfSMWwka0dIwFsvqtayygVBSN75zhuN2mEJ62wNhpsZ89/zGVZpzm1eXI7Py
nUqzb9X/jS93GWEpEBa6kiJ55/UIJ3w1gSCsaNZYr7q1hkaBsH9Hh5+BzE3KwBpe
hmYM4FH7ThpIEa0qQ+zEEF/eDIpBtKAz2k6wY1GfBnnvLpZEkTdgxNhQmCu07jAa
Xu5UYWNzNuuuQks8OD/8hIkMZh69fQ5zktwAJBfqrRmcXiqTFgRyOWB48yMOqlSx
ty/bbrB0M0RK7jaTxOahsgr+cX5Z5Iw89k3m/hSIVu3IxmWYrVM+VJWbhrKafJS9
W21WBCtPcMSfJq7qY5UQhomcqsgHtkyCBMmggl8TXCTt66Uj6aQtEeVdAlapB8fp
GWl/4YwgW9O7ZGZG0AuAbjdy7cVqzzo2ZymcraFw2F9IQzqLOmu+OvjvcjrDbD9S
9M52BNhIeXL5d1JF8eaqV8Kk2kJxl8KF+heB6CK+sKUfnOZY3dG4oV6oQNeqXubE
F+p22Y7ss9HxqyqN5IiKUkLBrklM2M7UfTv1jYmuEO7oJ6ljRspMkKz4m9pegtMX
nBrfcCpfYr1TULLUb4/ZHXul0ti6WGIZN2071QNkemmPMRa01ylZaCD/zlr9eci4
pNC9enH8vED4RHibdlAzR+6xASrRyOcQFPRzWVZj1rM/iHalQPnT1yA6Y7pMbpdH
81KJy5noDAGXEmvCjE3b8Y7P9PzybJCAFE36eAlpi6JPR5iNerlx0Y41AXSDAi4m
SuNg89FAxIsWmaXz+FiXr71SVbuF/EvbrkkYca2dCtzyD4uUTkNhVuGCncTy6VZR
E9aj7moMc8qgjtqB+H3h8bPMZo3V6drE7wcg8z9XKsBk9trM+poiA3qS243Tvib1
QGJwCOXIifJAkH0u1mStHKPAh5veq+8JYn7EpNilZmtWWxSUTuLcRoOvUf0+k34e
s83gPBu9e2XTQ5ZT1AwW/DCN6RUB9kiIAh2tgkMQAfDkncTNW1XxOOFmbheaA9mB
amk/tQm22+uu6dahQqOt8o9wp9s/W8FWTsUtLRthUq/NAy1ZGNIq0Q2kE6edE5Dx
y6P5zfgqLuuagJeeEfOJSgcPP+mpXvU1PLOVQKp2Fty2ip3bvprkc8sxo5oES/qN
ZWwn4GL/urebSsdBGVnSNlhpX008FJDv5FVlnTu1/78esC8Nt3iZhFAoAElxaIPg
iNZoyulPQMIPPrtJ+afB9g5vC6cSEs8MR+V0oBr+l5XmZFFnoIQluR147Rk3PeQ9
Y+wtk6kC41D7p2sio6Z0iiWoeWc5p5dzBmFDr39hZO0rD+noRAuyfbhMec0A2//y
ma579ShWRdzYxDxFC96SMop7RhzOeYfN0IP5UcEhsWgLkLQRz5eVAnmCa1vR8/hy
Din506/k90drKsFiC6Di9oliNVdOfSdMVdHWM7/v0kw971vGga/0yoX0xcWZ/VLF
P88dpAg47uZ+EKspzazyRr6zWYYcrgmFHKY4c0nh3/nIfe1OFN15U6v9UHw6XNxf
SonKvegJnl7uH8OOSdnIN17PElfhdLHN5PO9PJQls416IH/sgKBbDAepdPxr38sP
qjvfoepEaLI5Cs8WylQX2m7vid0T0gZuoqGY6VlG/chPqjo60GnBnrQ7no2FU9Fp
F2T0EOhZ3rDJmLPX89MnbpMpD1VgRcjrp5hw1A6ddvDdfjgbW5M/ZB4FZzp9r9oi
tVL3yeQr3/FJ3G5iaPWavKGq9Rct7+c/mXH2o4KO076E/bJSATvUCPw1idaEq08k
o5L/cMVfinhdKQqW6zh07WH7sltuuVvCzBYB0rau9U9+Wn9LAC5mXCeS9psGI8g1
9BMsymn7Y2fEcz3YZXJvp+3FG0rQgU5RfvpP1KWLhhWjKN23RZrhY9/+9cfEUHNo
WtsMRb9rDxZrXIyi5bQ4H4DyjVz6l0xWvPAdVpXjeAK/wkrll1ZRXJfQQ6mm35lR
W9NghGTBjjM0R8bl2f85dqRjSbM6OKRcoTm2kgWase8lKaIGUNfXlngP1KY/BesQ
zMwsLIFjIgt6qtTK+IZzQkp+Fguyu23KvHTkLsLGMt1IQ3xFcM+IbU3YRUlKBhIa
z38qWO2+0ZRHAINRWtq2FP7o/1bdU53PU6VrSe7DQxOKxPXOJ142zETAdPsEBUH6
Pz7QN/asTPlDWwzuv7jgrNP5V6faMu7Z8XpQNVG4j1yaOW+JhgijR5V76Gm67Z1L
zzJ5Pd5aa4AbT06MBzAY5N12azMsKw0DgBXa3QgPy8bp1BtbqKP3WOfcMHejy5aJ
xUaopcU3LaN2FqqpQudBG78FdJ2k38VoZSUMaBswZT0lRfZVv1kGQ33rV5ZrzLMV
6Fkm3bOB9qOoeUA8FZNiCGHp2so0i7IoG2Hk23LTvlqbg04h6nhbHQ/vP/Bz/zMW
BnBeKCfP82GMDFwZuywrxrgRqbniomJgR8TQdgfZTb4bdui8INDwk6K33Sustaap
IKeJs0Xyo92KDPQa3VHFwRojiOIMO2f83L0VM7/vzSr0O5WlBF26SbmHHnwTTF0b
2LvDr+Up4oiqBvFUjJLQfOvQkZ1cAws4+RipCfbn60OZ0ZegT+5vestUnSxFRHaH
2WJuAh/oucQKO/RBM6hYOwSAsZwlnZZ2bayAZuEx0h0GihMeE9Tx49V6Dk273aZJ
ytWYHTSvvoi7I8V6X0YjZcYZMjoKqiW4zRXWOVvhPDDYUcz8q0TB+tj/Tc8dCIhu
5S70NC81rQKqGUFJuypPuXXO0hV3bkVDVXRjQtUBLEYW8yXD5r8JPAGgi04yVKtP
UV+y2PB4SXS3odjmSJo3LH7JQmSxcmssqcmFrcI4EaUQkk8a1V8aP467Hf15udro
+IkZfSJeOYyqV4+elGonsQ==
`protect END_PROTECTED
