`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdo1/d3SGR8bfllh+LyI6MUtv4QoO6qGBlbkL69fziItfQZ0InR8zoC1dZU6AHVd
9jyRkLTOvS/Usv52YSTKPdflRB37bqCzK4JE3ZMVbesP4hx8PtxisT3Z0y1gG4eB
IuQj30R9pKen49MW/6xcNLTo3jmPyuoQEakSpCRC/kR4RkeIECzZCe8wB6ccqLz7
3fctbjussQmlWrbt8Y3y416q23bmZpj6P/ww08Z/0e1DuEVGFfyB2pKQKzKEzHzN
I4L7IDc4ov10e5YsickvgXtiwqy9i3peIt27sbwFsz+R+31bwCb8ao6PAmAYUfu7
3QoEDYl3eyJrQ0BDU/hbFUmaZPLh1hOr40p5m58SL62xb1s31aNdESFU0H85JCdN
aW8lpFJBZL6SlbwTAD+ngZBJ2D3UAHuxCDdKxi5JK3Cjg2CSZDLx9iPRoKlM55f/
SAAG4gYCzKKf4RjPg9ckuIvrWfcI3B0+VN2t7bzb4a5oGW8fFeonPdVP9l9G7200
GoOqsInYPHO3FKbLbgPb2R8orxjYgc+2nAyTX8263KbWKmmB1VKBhFvUHm5RBt60
XyTTczq2aHdhym5e5l5/neJwhQ8XWkr+GdLQ8htZGLsNKnQdALtUJZrW4U4QseqD
+yKiC+V5fltUH8+Wjk5d/K3thaaU5pnK1PZFpndc+bzULQdx90xoE93xRuITDMb9
nycckPoy99InJdhxPbJ24oqN5WuZ7JynCXlRQW/Hrw4=
`protect END_PROTECTED
