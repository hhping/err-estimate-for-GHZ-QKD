`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
goVx7vxlZFZOlR7tJgkt2o8qZnXdvF69112iup+NUZdErvrwTyMId7tkaFRx/uJV
hfv9jlI70XwdvZQJnymrkX5TJ5eWzq1iLOP14sgDX1MIkuKAa+gCdGkvWnWSMFvT
dUblTOKw9dYgDz8NgcJhnWBVS0q4ZVen0Ysg7OHlJd3sGWneXgGhRwtDZnT2U/cP
WTC0rB6IrBnN431L2QRRtWsHwCdQ9Sifl+ewrGK8aey+zV2zSFfBGg6KwL9ShopV
V05vDZ0eqcHuezAqUZgK3LMndAf8cCIhdQ3eHFrNXiga9EAqcNlOyIyk8QMWUTB1
Trw6Mg2VCFxXrH6/clNEntmXWFN2rZJ7UTChsY4YYAJldVph3xOnSIo3sXD9Pu8K
YB5QsejC7hYQy8FkmkyY2g2PeKI7bFLgIcq8N7/bPRX+zSnmjiFRclpa7FJT8bpM
bmSo4XZichM+wODCkVdzMzCAb4ekqoY3RVyHq8dZMVFdRipzz7001qrbQrZ9NjT3
4Rl29om1+HLu+PFlMjoDZf4/FahubQGMhgPji6p7Iegoc50oP2tPmrTeLK0kj4P2
TI8T/fi/yY8hJG+3AjJstKcN2OnBVslFg04FmFSoRcJZTrbiDfqa8h/OPPK5lkcJ
FBBKPLWR4nrUNewGBksWGln33vb4IXNF5N2RoUeCqEsJh1zAHb/n+zXmE65VI0bp
KuOUnq/J0bjVb7KOFTJJpwm374EK1tlVakZAf9szgwqveyUC2ICELOBrLwsV8QOz
VZBXxz5AZrtaNPQpuEIlAskSqSkpMtSew64DHC4JMt95eezEQjT/7Zfr1lHo3W05
VJN/ed2v7pvU9Rh4WijpnilAq0aWYoLKniLyzeL/7uOvSppAE9iLFd2r6LasUwSM
EHUfgQLTFS5Toirbk7zOy6W3p1Ca4TbaUWLs3XaRxS+FWP7RzmI6exQXt8ZbRQSd
RtqocRSoxl/vu1L6YgpoOaiBoTXZjfrpZVEqvmz/pCvKiQjUr3eaZFA0qAfCTC8A
Zg2iE3d5toDRvlMYF2sARJoWF4d3g8i0O+dzJdimlZ8/OGeJOPkieBYkeVYBfXzY
YP4KOopNJSwS+xHbL+H0qARhU16MYSkk3PxzYUFZV3gF2B1/zmQc+jzHUWWB3/3o
y/2Zo/jHPioek6aJ3s6Ub9wEesuYvaS53XYlLGYukqSMGjQTMWrb13eivOSn6N7P
xqssN6+OeG9/X0QLc84WXwG96ac2HrwmyW8AwK61RZn5d8MmO/vDZLH/Kaaqd0WD
92rn12S86FsqURKDNCqWn4evb4PPsTi63uteg3IUc1aOXnYdhROkG1/qu8VBr3O6
N0MFftSUlevd4hJHpN/pJ2O9ToiY/pkCAKE0O5AJi7jn+EIbt7PJMkYXSsvEIQZ1
3in03Gt4UrjqFm41TfF5j0/qZkoxnEbw3F8egBpg/gLR1GxXZAgjHrMUAi/yqkCA
wD6PpEuZ3MUdvu/oQl9ZQGMcNjKGrRWdztId2dDGNnbGtpV2h6LW5gClvHZVYy+Z
UhIGqbq2xyP8JBNxnheNdmNF6V9xUTiYaNEsLzhuPWoB5X9G2MutNfSqXZr2phhM
RprY+2+OHPYq9Ea8tinjcqK3NlOPs941oa02nQAv3VI+cI+Fs4vPASTWyy0kPxKh
Qyvo4cScDoXSg2+QYriwkDWlF73hMXU5oqbWnN7b8784V4bPVBGfJ4TzhYcirnl+
azjKbkfJvKG68dwd118nnGI1RikjAXtOKOfUFQAkGLxB0gc6639MdpDkB3rJP85p
52mUKCkA0612kWfhzsl8qMuG9in56nYVsgv/xVP2pF7JFRekUHQfOglv6UWIv1XW
Y2Qc9oRDYwwTUkndlJr7fY0amtyabo4EojC5NvMOzWaINJLw0vE+Q90sob9funyn
EuawxO3K1vsokni/UeGSmRaPzS9U8r6c5tRJwsyIv8OBg9qRkgb+1hZorjveTt94
t6sUuIKxk5GrWYBWKLGjhPp/+ECziXEFBFcEQoZzNiL+bbVIo2ySh5BtsMvsPcSB
hDQjKxW9fAeMrp54mkpDgL6EqRVtYUL/iA1Vv5r8XvnMonFEViYUsdrmdRFdvXhP
2DWlABYyk08g15ZRuWBigiFvgivZqwh3ItipkCl/k3EuazvbIPqwSjbxqp4FEkNy
aNl+2HiZR9o3Hqhe56zn8dw1AGhqmBKRPLUeN4HRCvvDwbqKs9l91p1cMPZiujXQ
1c0UEy+hAwJAeE/S+ef25OmKMIRUVbyyUEckVCh2p4H/BQhVw9sKlA3rF1GRhmIe
lidQ7kWhXcQm9V29lilrulre0LGY/Vt9R6be3JQ5JAr3XF/P1hHXuW6oLDHbILAK
ixR9O/eTIxPbe/avcSCb0jML5j/UIEkCqstoYMu8HhtLZduVQvOp0vh01XwaVjJr
LxQnXcTocDs1izXn6UxFFIqnx326+jPdLijqVnxQLPzoaWWh16CPTlwP1uKWT4Hk
s8Sj1kYaw1qkglWCM/UTv/NprA5fTSpd5j5oLZuIpdDvBAf89mIRxRJxXzPHmTLV
9vhV0EuFCSvEySYObr4TBiDhuYSTkQADK77P5uatVFIC4d+gVv0SpjGfFsCoqIIP
ECl8Lq1M/Piav5gWtDzV2tCAUhnlLlb03t/BWwzn1zBdD4efQAER+FR9heufDYPK
Q+fXs6djVGvC5ImdWoUY4llDhq10ABFftSoRSYQNEwg6S1+XHag7LqNrmsMwygWH
EJGFCaLOR0eszWLftdpi3bkSh6vo7zlw9NQnwfBkAf5c4VgF3XvHlglbNnAMH19E
3sHuOPURDbsBuEq95h9e+KyRDhhQk8osO1K+ESaTh052k6a6wCxvPY90N3esxc7q
UWDkhVJtwVH2DZ8T50U25OOy/zxseeFFPRza/rFOeG+agbSu7jRuPg8/SYtYbYJ5
cWnqd+0T7eHpX2p6dPngeIbpvA6FQHcSFA9Jgcx7fMvIDd7wLkq3bCXQAGYsXy9O
Px2fUh853DBYtW4lM7PVJinNQo+xO4A/DMOScoBUXEQb4rMvpEHQajrT4Kj8faDR
2Dfc4pxjFgKLAP3qBOvkjwmvYYaz5JOrhi052TjrlrXQKvSV1zPRhYU8TldIe3wV
Jg0wBKg7IPVJBgShKktkna7Rp07+isnJ+nKfHz9cZ0baB2IT6OTf6K5yYH1MbQ5r
I39KN+pl3gRSNXo+4sjf5sVh9sD/6GquDGa8lH2C0lj9/vH/JjCeHNgZmDrZVpJB
1GPglWxS/aWf1XFQojorKmMIG8mCIKCK/X/PbNSX5QoEI+G+PPr51AVFVGGIXeQ5
UgcZY2PxI75RZPtemJGZhGeL0SuYUWLkQdUtiHOza6EDUkxU3jPwpha35jhb/mwh
y6xZoLsZdjyt0TEB54+ujPpbSUCNHCMTeQ2s2dwHksytTIfmWjyK7BwlILaf7Ec/
mSxc8RvTw3/lYGpzzRqOa2mF00hztDl74TNbwo3JQG51Zu4uI15SeZNdJ6WlP6N4
kFVDbYhc8mSkt5kR2K1F8gnvvFwTDLIWPWP18xOpqjbwjPweoRYcxF+7QkueMzca
oAEnQyje/5jW1holA3ieaB9CWcWGneIRXEC54KlOtt89JnUx2cMeXviH4nU0Smtm
mHOFTCwK0f4PimDw8D7cXrFbfn10QsnUW+KNR1zoQN2g46WlPDAEAL34oxpAYdJa
lc4JfEnfhNcr3sz9LG+EizGFHuFtGlF90S3Df+czzEaTsODCc2ZD1UTYiwA5E9fW
hB+wAM7m5avf8KTm4pIsMH2DmBnd5PCgYOE9fJRvG/LKPdeyVAtHGWKfGOvistn2
y4TOM2VIBM8jdiuGWiIVlvS/nPeGavNkOXlyeIyLB6HZ/fIr4X5VMNIqUnqwqGoM
Tzsyf3K35/lTPA7bXebu+hwNl73Us2D56WXHUR9Z+B/qhrB13+GFUCqOtcJ/6hqe
jRLhGCPCAGdhEupJI6OaaYi5Oa7haRJARsZSfll3zNPMQWX0kjoRaO1NOuzIuHJa
6dLRrkpaHVDoasaaR38XjpPqxUsXuJvlzkgOGPnw/jsqKc6F7a7Cx3LklT1NLGhu
ewDB0nGPR2HPLtM8UikuJAfyaOQOHStasEQYi3qQSrNpqNnAgc4LgkwvN5oV7tdD
nTocNGfm15p4CFwKogAc4tv+DODmUW8U/aE4ySESjztDYvCKXu5AiI4MAe4TRhoM
xbXS+cFnclsUo7vh6R0kG9bEr+i3v5Y7IL4snwXzt+M=
`protect END_PROTECTED
