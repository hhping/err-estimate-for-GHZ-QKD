`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRSHb7BKV3FonvZk6U1Yf/kb8P0B0k9lw45rtGn6NwVR6uoZcomI2vG4YbUK035X
TwlfehKRLVSR6cq8e+Dp8fzMKBEta6WXrqYcpXUiSFjCXKyDjnJo228b6tOMqckT
YYyGzBq3bahcATqhC6aPI+nhJGJxItb3SCAJGMZ44vAXo51dKV5pFfeYVLUCqh+d
FHNVV4VOScibbb/Zhadg1LvxHUBS2Lu5HUpz9Nl8rmBa6xIs3nJPz6wC7rJOGGp7
ox6rii4NDd/n4jlb0LGIS9pZ3AJLRlsBRvpN0MuRmtuJ/vHCDIOGmg9z5wmfadq6
LwqaDvZCrQfzwzpar3Tws+aIZWEQ6nBejRdI1jForKHnnRnZ4I0FFT6MSPfPKBR1
JFEFXb3kgHiHKDZ4ILQNOBjvt+luzH+0jXu1r8nBp70QaFkiwxaZzB5nW5fWieYd
5cCUeJ8ueeaosTH0TQP1m+EgOW3CSRuk6/nmGEGYRbWEz3LAhvDyS+qL4GM8TYKF
VzTS9fiMqBQQ28WXs8hM6ydeah6Ewnl5OAcljgfgqAd7WUrPVX/XOsATk7LmKqTc
zgI3jO7RGbSFJtboya/YeDKzKTRUBdHRMfpPlK4T8np7kv657g3R6bE0O1l6QAfm
TymiXWNuiOWNQArxnCutw62sLt12ayvDTNvdQWmmorqdTJoegnnbr9U7Vs6cqYbq
AsxgSW1F4ujZafVCOX7Yq13M+JxHpOqAITwJ/4ekLjbuliGNeiRCdb6Pq7K0drEj
mzk2wAgrHZWAkfB9SJ2v4L9U06mBm4pWd7gSb+pRGEiIMRvjgnxrb7RFbhcA6fLJ
Jic7sg8sdbliFqJh/Xs7BI01fyPaJi58hvwnUWKBJgmBKBw7d9w49dA0EC3V2PkB
QgENAMj7TQhGn7XIwrXHnRi7SKDKqTPIObTTQcKRkXgciX/Knn+RneLSIHrnTT6b
fJMHjGAFcXINJQbGzMh8Pyez00yMtYRNdWgOsiN5aFDFG4NvU27eXX7Bn0PCOw9J
nLM1uZT5DtDUrPLZspTrZSC0xFXzOl80PchiHxfwHqMP6/XnBktIL3I6C/c+Uh/L
eMuFRrBRiuyp/aieN6+dKag2bhmg5bKqiEIWNoGY34839cwftyuSIUSqdpjxSgb5
FufwLagS++osj/6DtA13zZVw4gjt0s3SKAVttx18umXHHu6h0JYF+r+iFThUJg62
vCJwLf5WL8z4HTqDU1hHZbHP5rAWcmtxuhDCDJBCWNRJxMPgPm6ucTGE6/zy81um
9kUDv+9RseFaLRF0/xMPZoMURTxYTmzCA8PRAu9MqAWTXCKo/hjrBMTA4OXo5PrP
FqgICj4nlS7Q9w7X4yT4G+8UAW5fjR7H95VhXbpIZst4Zltz9RlLFJ+VCyQ9wNoe
br72n9Eg8zs7KN2IBLPdANuNiAVstwGlaeRbYAIDgE01QbyoCNxEXoffEGACdqTD
gCuNZgpHPiDPxqms1egOU5xthLkXiYnEoUbEN2rSQwqqE/0fSukwslLsHVhefYG4
RTQXiWFbephLmR2dS97G6ZQoIVYhhqT78m3btTbFK8U=
`protect END_PROTECTED
