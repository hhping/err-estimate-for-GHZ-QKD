`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kFYRQiqIa8Q2Iv0di49KzESTnuJx9mUu8r7C6i78ui/v3R9UKOprLoMehIwusvM/
gHYvj9++AvdUSgqYyrWoq3B6n/nE9oesLZUyfI1o3WydlAy0zy6U7D/NlUgrRbsN
PcoqSai/iZw9mDNiwaj9W1ZsAzHzVjJsjIqPOoAea4v9t5rjqV+ff7qeYRrbez+L
j5p7EtdjkTuMq4jhxEFCRvodv4zUNQeVCBQ3UHjtoj5XBC18SYHlsIU49sOt/it4
yEzu47BMeKZ3gDZlhcxa7u3DRr3zm6BMvZl9YScI9gXIJ3v4Sod8MxlJpIEesDMy
FP1wcaLGosyeODdimbupJYmmEJ3e+JGOIZq+Hx7AOLDsbPuwvk3nNP94SsoEmPDv
CRtOam+N7DMYnUSGFi205HvQmmBvpU3NsnvaENam/V5gGp3E9CdFpSB090gxylHo
awmD4vMAWUHebSUwZbPeFqLb+6SBEa3iEoiZIOkDJhR3ciEV8jZWJcI8X6GTFKq4
MOfjNODu/o5njwAi2cjsN0xlsAFC55EPJbuzYhBIKEB6PcrJCjEZRdr064lzoOi6
gHDBplAaK4C+CylX8fHylOD5zgeJaOPwQsT4dz+/Q1pPbTuuj1IbUlSlZBz9Tjcs
Oy6jNtAIRqNLyFWrLGy4G6H4CL0HzUaJo1zLl34jIvYK9Zo3ynzsLd/UPwFTaOuj
qAjLzx1gUBuPXJrCYzMaQS4Dx/AufUa3Zcpo0Ivbj8z/s+yHwD+CPFIBTKG7PWO+
QYuYRT6RHzEK67cx9bwy37h8dj9cPL4BmTGwtivx9y+/nOkmgulmYyc2RfQQ/O+I
HZR/y8ZaAogovl38oMKGlfenbLt6a6ZMMym9bvtfynB9VoC+PXIZviRcgy1qiZw1
SET9Ri8aU8Qu79tpNYM8OmWSkbYfALU6s1Mav29ZzSlWj9xzESXZAcHumBwAhsBO
nXqgm/Rru6zoltlbN5nr1NFS7TZ07q0vNQ9qIOOruYh8P9k5AD/77f4eMMWghEFZ
p1DowLP94CHy8f7WLS8snYrvClwQ89M0nDgCgQSYxye6Gr+ISiaKCwecUKSXSsUS
4US5hY7lUb9I/hcb9OCo8ctWz7jGeYjAs0uSioz/EdKCkje7Mg9t3CnWWS4uK4L3
U3oq2NxWNSsFwASLOEdwqMQwvQLf5UK3MQi6czBPTmHvxu78V0p9jL32ln8TVXa4
diUS96MYtl854eFRiKbscgDzBS32AbuzSihk7a/Hbq2pWGjtPOl16vTNBgZHXlFl
Xu1B9G8V0Il0jfNNP2JW1dxBsZ39HJbm5o7fBZu7k+YWAFFvZYUB3nCufQuIv5b5
FZ4n1VxtjkU6lenTvzfb728hbyMYDrnNhxUCELB6A2qNDSZ5HrLBZeysSCzutfA2
Kmnh5qP1qZT1wAnzwugIU8YO/JZ5DXSVNxrkqa2cc/k+MgyDxC3MMdc7RIvR/nen
`protect END_PROTECTED
