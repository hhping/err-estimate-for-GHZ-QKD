`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mj1ZtwMZORduK1ufg3FOqTHTpledx5nAUt2Ri6+a11norCpM67BOAmU6WaXVNLWD
8AUOwzoh4TAO6dQqTIPQIB81YdeLLUxFlVQAWnqwZnjMhckZzmeL8SooN/5BRfkf
8fwPWOYyjlirPvkeIL1cVYzOu+ZNHeR+cT9mBQNctxVlNiqIrkk3HtpGgjGqcRky
MGQmN6KZNmOTM8O4ckhpZFw8MbZ26J0YC0XA4gr3ZLQZLdvSbBTU4xbEHl6Y2sbB
zOKj0X5u7SoxqtaibtXgfzxjn5tFbc1Vcv45ETDWUxaOcDUCX/jcPcPygh+qA0gD
GXpOmQq7Z9baPNWwsaV4/0b7iL3WtbrRGoTFAubtiZPDlhLgFT5bsLX+12X07kB5
bojiqdoVWFtV36CVvuFIanFllDIr4b3k2dFUrLWgLV+ZTXftZV4XxZalmSt80eNB
X28iBrXCJJCy/QPLGwCWjkOuaZlOFskElen8CyEfAru3Gkgk3MENPbopGjyu9tlJ
FJXKmWnXX46EjHtf7LdvRpzYJwQpo0dUU3i1/li62Q56N858uyXRJzmVrYmXCKF2
VDNYvf/QbYEPVgX2VQkV3A==
`protect END_PROTECTED
