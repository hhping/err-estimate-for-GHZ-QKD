`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDVwHU2awD3ikPoSDjiSU1LxNBwVjXTiztqxTtY0Xwgf+JvecdNdYh9PpXjqZBq3
rTN8LGk8NKF7WRP6jBAdUIKKqJvM+ItPtBd3IayeFhAOGttl6LsqbyfQS3oW53AV
S8Xj7iSGhA1VysNH2I7DGNvrCByZ3FGuCmy5AFkfW5MXX7hy9g4lWDaM5f6ACSZo
PQox7I57EYflk5DL2elr39Tyq5cNKVr+D4BNd+TsAEb2MgKv/FP/kcJVHaRLeQbH
AISxe6WNnNCxCbqumx8BT6I4YcOIJ5xHeAadfbgVFa/LqH+ZbzXxWOB1xLaKsffd
0V030Nbign9nesjxsPfpFAI2eKzazmLxbRDQLp6AylmlbtZj9iN8zQ0UE2OSa6wq
LqbLHM7NX1dppCSY73GRIgtDceWdijm5BMslgz1v2MxL3JZg6ZTm4Xnd+nQGAone
4KVjXZOJtyJchxo/E9pR6I0U798vnSicA7DAicKKVOt8q4wKIRAdmiG44tI5DQRx
t/lkja34j0d6DvjuDHQUSFlEAB1fKO3/4Bug5RATbTz4Am1nLJRypn0gdl/p38sE
M4dCdbA3wPITikH+Ovs38GL3idMhK+T/Xuwf6dQ/3YE3FfMZ8tmOKQJc/bahsR09
t/7t/zx0uDFkXRqtTvt+N+5A6BKtOyFxxc2NaSZK2kzWVtVu+YJQPSzhu8uen9Ny
EQFWvnKnBwooK2dxop+ZvQmcxrMUek787wmyDA89XtLhBbafZXTiAkSVqN16mtVu
ZrSxUBPzvVbhvslMEB7/wRP0ZL9gweFTXxN+ERX1sNeHUx7Ce2ANMUF/hYonCpdp
GPuvaTrNJcFxaH0bMpvsSLKXvvXVuE5XrSQd0UI4N8ycjYaxquMIhaOkkhLb6AaS
UkzMTKbTGOuw7ECE74zvPQ4naPFucGKLSrTAuJ94hTWss52rUSOerQqbxqpBwmo5
OGNn4D6tvNJ062/6Cg4SA8NQobuoarVW9pBmTN8rTt3DYh2C9fei8e9O0YAbvFjl
hxSYKRvy5LPMNcDzLyq4ud9UOeIm090AuQLmDSjzABqxl3N62cor34sI1J7fJrNJ
7UtNqKAnGQA+OQ8o3mtL9H6cJ3rmSKQsQWhmqNYcFFrGE074r6FqZj5wCMR5FOEO
mt4/yCW2ndmQcRFta7awMrsLaTwRsRD5jylDSieYOUL3D1NAN4mfa1lf3HRqTF/B
50Z8mjc0gNO/Yj5Zh5L1qB3QEqWEbrLN09S+Tnxt1ndNyByNT/HoSXGIoDDljYWT
Ixrsk75q7IU6FHxYc9dcNNdVmaCpTEuWZol0c5s06pA=
`protect END_PROTECTED
