`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZOo7fqKTBlA2W+EshaPme6MQsuynGQOAH7wSwwlHWMxBd1RBl0Hjrs/LtpK1ESxz
QDByaBiJX4oomwsJoV2ICzy18mbtW9IDkQ7y0HKzirS39X7nPrV/6C3xZr7AACaR
FcKyLUL3FRbbd+qrCMqI7PVF4d4PEu/e09cKxIDGq8XR7TTkkFNTIGy79fzoyfSf
mzvgIYmIroal+UvUdtXSSfEOxaKJsm865WJ0zDs5xe5xE4Rjh0C6iNqln8M3Ki5p
snq8NKjaty8uIowX7IbGNoR0tfla5Ox1dQarni2ra6+bQvMH8nxHJXq1mAqF25bo
AQR54MPTUAhX6r11w3H2sZOmyiyMJcDl7sLLAZm03+xR2KEOcbOXgF3Io0mPtAm8
K5Uz7+aSxqMU9n8s35aHBJo+2XrT/WSnMr4fDR+Lr2WY02nJv11EhW98R/qnXlx+
Tnuah/zvXfzowPYou9Tm/GhICwbOmFbfg0na9Et7ifQmyZQhM8wG+GWIZaMU7ELt
0CA+Pb+XSrfX8GwaEyYgObbEgiUkroaE+HVsJtbUVmR9VzFKz3iOzVNcpwKAX+mc
m/A5zYTloh9yqsJNnPEOVS+POdBw62OMq1vstPrTWzFcATsZszLRhbsIcMl2vUGq
ql49JGyy3MGkxUQ16+PWcS36qECilBu+ecHewsL1ViJ3/2VX5kzgIJDPbwVa2UNL
rk1o9AnyFyRs3Di9M8AK8m0OOEUGEUYK8oUOpC+my2C2ctPLMgbAXmnXJ6Qzv615
ztkcav7aOjiLhng2dOeuTThQy1AUhuX5L4yh7nIDbMG9Uog1k4ig7qdrFx5uTiiZ
72tIV9U/iUUwjnj8+kKltAVcrrY2mBcWy8NLogu3EL1VruBMmrXz8VgCUjhZ+dUe
gxKU6qtU/B4n4g1TIMNuMJfK6OPW/6UgbVDvv+BdPmVcGKlP/G7qNdodG/xkmOd6
fLPZJlc3n4JWSoQiuX0+v5VX/jJbFaq5TodlWfweFJbM3sdd6QtPdfqXfpXAr/nE
1gV9hIzUPGMxxfzruR3ZJl85SnoG3+l2rginPwVUhGPv0woZhvIRAuhbSn+9Gl3n
aLG9s7VhADYDpSAGHaizEs6s0xuvunQ89NDdGS4k21nL03teiWqgAVoIQuQjOj3y
9suKHkNG1EnRAVFgIki4Bhd/KDuAtRnc0hdbQ2KwRsY=
`protect END_PROTECTED
