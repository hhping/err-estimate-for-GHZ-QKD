`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGQ4lIdkUmQSZAWgihh0R+W4jsUNO2ZAERWK19YeDkWcW5l2mzTIjfl3HRBnDuNY
q9lg3ozw14NObMI5eslij1EHDO03s3GvkaA0L/bOXJ4kvrh2HNDMmZ5qWOQTf0HJ
oxbwh/sWE5Kn/IhQJjcVXpGp1LKKFsGW176ummgebD8Zdq3V6AFQWvEd9MbPp7Lm
B9eQBY9CxmBb5BQLtpDNWVJiBZQ6V70RzUhklMkuvZ3r4LoE/VA/eH27IFlcz9Nh
kHLloTNkSU1XcFBT/T+fiBoVg3OdkBmwjHf6x2tJ3hmF31SyqDwg91NbsI1S8+6p
YPdRSgzMTeRW+hKnFeDqYSa+91xe6+oUQAyFmyYTKJl4d9Zy5QMt2XqfGgVhonwJ
1wK69/YThUHzFRNPM45vBxBCnieVG3N0BFmj2WpD75ZatUVZ26mM1dSBGinj1kmq
4AYd45rCnN8PlHKwcEGrrCvkkA6NQh7Qk//P8QjrDGKhpDnHirO1SiQSeRuVaDuR
hyXD4ABLYL08fIqNmZrMubGopY5cbC482h6fJ7BPDDnN7QckosSoIyfsXMJtMXe4
D7L4MeWodM0nlEQ/hpAPwfSOeb1RkAyKyeJ5dJd8DOyjXlrIRePtbhqNRv0dJ2+v
H6nYrbRilhx5yXNudLVlD+G5gJhfSKheQRZ3zpldeDL2hk4/Jmd3aVeQuT0jhbUD
kVgsXz9SmUyZpczXWMLW236W/1tm/8jgnfgAx57feWnLAPq0c7/cVtEYMomO3Q2/
V+O4UFSxJyQEbVRN2MPPT9qPhLLsZey2tyrX1EgKAkZR0m7WJf4v9KZlDhDFyUMe
qPV3CKb1A1+1plaV75gEaspuQe7+dDdNyslz/cZCLuX8iyP9dHnw9++XHxXtb8CH
OEGxE0wpnSH3lDJewvzfROoVgqtwLJjeFcj3ZMkL0dC/qTaYsbTAty/5bmbeeK41
kaMxvhE8UALCuXu6JWIaWc74sBiiwVGn/hFVbm3P7IWCnuCQiY59/UZB7iKrQapP
qA+vsmmPSxYZ2pttzrD6auJXxF2aX69E0DaUoa8tKYGw7hCZMMLV2+yMLFAYYKKw
ytsuY8dX58iBOtT7+omzHzQ4z9rdnNAedZUxWde0r8isXtEmJggkLHAkFeqYYe97
7V7SC/5mR/TfbBhZnm3fmGHlZB23gouAj/M0j7Lo3Sbur15RCJ+HHv0tDvMl3NWj
MtWFcin5OZSvyvkjbXMgVsPm6GxEp6Qvg5mUvoTNpQcMRibWzZoBgG2x3zIcz4Gz
FBEHAJl3eYt+dCkWXSdMf9rmYW9/uiK5GIiJ4xAq9L2rXbLH0ZMlgJlvqMHf2UpF
Ur2uvrfzG25/1Abalu3UyyGPfziw8ieOCHOPHDqwg9gTctTvqST9enW4rXNy2X7+
M2OpbDb8uiWU72TlQLobImsg/VkPGVqK3hEk+8agI1AIkqEh1hmoanyvr/wZfCmE
DsxQC9Y7HYJHLM4L8/szJEMLAc+X3o83Wc9FgWdEDdOE0j+gCscXmFxUYP/1MJk4
YrTiac9Ck+Gg/mHdcNElwvNIoJ+9jJbwiJ6OUy9RW3898+VTwOwk6gSNZTX3Hkel
0xYDYU5ywK/yRKeMcQTarVnL+J0kqeFhNI7ZBADGPUZCQLx2k0VEV3TbxCdIOmld
ajh61GPnu5L2FiZh7lN6aHRv1bTFurvEZ7Kkr6k1eBgHkDoJwnFN0Lyc/cwd3gyw
K3ouSdk/qdsgG+Imv1T9dq3EAwYpi+YpO7iENGiQyO4836FsAK7B0mn3qaxm+KzU
MB2l+9Yuho1SpeGFnJqNvIkx7X/wW37yIiNf+x/vi4BPBmQXDycAXpXa08ntkCN2
Yj6pV0QrppDj2P68jgAZMwKgl23T094Y5D7AvpRwmk1kpnKHCuApooy3LWJdGl1J
lDMjpjUd5T0RhLvK3nafmspveFNdY6itF2lQoi1zkjAMO2AX3XC6zlj3BTVbQeM4
B9/LXmoTxEP4YB+ogULZLZgdta4a29bEQty1O4tn6HTkfsocuySQTpdtLv8RzG7z
CpR1JNFEbbDMhJDHADcJWRbedcfVkUOD6b1EOy4WnEGevl4dbg7+qG4Xa/0RaRaB
TOH1kNGmoS6DzC18FXBQOBUWjsCOjVhl/qNiW+HTbafWMp0G0DTpmnQnIhZCGIoL
56/TIQYVsWLNxjcvLnh69KjmL/bQcQ48ezkuF8DRT4oZ3ljaiLmo+6kwi8OYbb3q
KnfpiEkmiLMep7tHgUdgOMJ/nDAPHsev59g9yPhRoVzillp5TT5ZA8O1GPvDqal/
Lwx2njmK0GaGCYzECsbQKC7KJ/4KPAdQhQ9kFXWu77XSEMiATYEM6NuDxf+1so0F
jLPHsQHL0pxEgl+a4quqS6fqU4hWtQl/RIrxCy4tVr98skKblde9dJ5vprE84SHk
dC2Lsfmv1n5YzToeYaHNg3u/HZMYa2RWa5OvfJ//UbtchLIP58o0LOhXRKomwDSC
H+2yB8mzMg5FrFb1h+G8yP6zuwVu4Syt1dZT3b8T4Ha1UpcRH9OydJx8mM9tQsVB
a4ATrbvxbqYptRwWH5wX6UHQ9tBFaU+epww9K75m3sfI/5AdG+l+W7jKp9Aa9YU8
TMejVXvE6LyABQYoWexIA+jfPrVfzwARixd0g51uXgWfB8oGF56Bich/R9f22YdF
NVxCMM8GS5vA6rYjEZqtS8V+BAdh/Rp+AzcY+MknY+7/PV2t69Iev3BDhDicSzJg
o0KdG5EEA3sPPl5v8JA7lBXJzv2BT/5L+Jn2FUoR+YwTwxhRkmKvU6Yonyj2oTEQ
gQFnoYo0/ul3yCXKPfnUyT4zYheyhbA2fo/eDbSqYr/V8zsvQJDNkSGplTYEGLFY
9PHsWYw+CbCHsE5Daep9M3SmwRh8AVHDG775saPnhF/GU69/cGpZOEpcchlFXoho
LoUuFx7UkCRbcxdIvUNb2myunIK73uGezgDSn47Uc4+3y3bA2GYZoKUVmRZlvW4b
fjltcbWknG59oCQPAW382bJXYOo9Rz9+Af8LJFER0+qUj3hzVM1oGzhNDw0enfKs
oZKbQjSL0K8X8gGtIRVqcVz4Y/BgKE59wAvwPg6nQ7LHYVbWdrNup1TY7+5FUMb/
7i2xNaNPu4xu84u37m7QDzJiNtdQ1Dcgnc2mZVCe4qI0ic21bPQGH1jXDN6QFlpP
+h8AbRR285PhpW9HOVXtn/ohnD7Y0i/ahtENX1LBfmsYBkbI3IKA+wnMwoY4rDFF
vjIL1Q2caiXbKUBaao/lbkTY19s5hpgAW0y0D+kWyQ+zDBfVdzvInCuvZ/IwXHNG
hjWdSRwAQBTwfkBZ80zubrFDK6BwGpIvvBUIUXThqwMeXH4ygWTtqSmVN46eKpF9
lFTIoVffHwvqc/pqcCGxEOVugJmgaR/WbkBDONuDqoefVfYIo3QokB3vRvqzLtdE
hYwZ0mP8KX3HqoabfxoKzOlIu3h3eBF1wIqLsT9P37m9CpIDP76nQcnzA8UN4ack
BobaNM/lU0ceeDlL/ni1Xki7M1hLVzPrC+phJFyZUzpSpsaRyA4t/3c5RIxMsMOT
ovLGzc2DXJOHm5AE3MNvZdkI7smac+AT6DfnzGTH/GCEyvtMQj1oX18fPtR5VSpK
NETeixGyiRMYdzG33UEP9vbavc7CX0NmtOg5jBNLEoQfLC5oV+z/KmMzu08h+tVq
uq1MuO1M028hKvh0hf40aipc4MUFtXN4/xG58OJ9lpIP21y3tc1HwVRZLPbHfzAI
xBvU6sjevPlBhZcVajTSlaegVjcvWHFBbawPfoDe1veRz8q8ieNzwDkRvNzLkY8w
bUd2sCpfno+zvDLEPCImdlMz4gdgVLfSLStnW2BUKI3qoPM9jhxKO/UFtw8zvJ1c
0R+hOiB+Aaly96vDdb7MpBFwTbrMx20uwSgiEqmgH1yNd4F3xP5+cIDLGx05/6Dy
FKafL6XojczsWm+NzXe3i9DKW8OAxMM7MDOWBaGZwYSXyXPFzoTWgKjYq56DsGuT
kRZhn8jCBE8pzpB58uGS9kJz6AH3OmVzeHy3g7mj3MsCEZd2vCAI6JZVlCdAJejE
QKYCse6buK8OIAxjCLY0Xw==
`protect END_PROTECTED
