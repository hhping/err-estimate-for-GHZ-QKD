`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9eGyso/Lv8SYx2KZa18gAlU19ybGGCjilJSOA09uUM0M8pVoX0heVkFq6rSNTcon
y6VvG80NL84S6DsWgLdTQPW3DyZCMB+/VwKSY5IrdFja1eXbU0s5OspIqAb/4MGk
DhGMAcu/ZdWEGZPxqDzC/jIN63WYOil8izqshZcRD8dCml8C3PpAjion3iyWa989
6XnRhJXAj9lZUYUF0ZNGPqL4G5zrOcwHGgz4+IBGIhbIwEwqEpOf14zriGkY/qMV
ExYf5Je98I8sSSFtfmUy/UWAhxGIIOHorcU8NsmslJwchU9SagRiy7u7eGDYUakI
ldQSBJ59k0iIjtjkF5yyzMr5OFbDAIB+DzdpGG11x6+DN0gdPLvjkZVJSnOOnseT
WW9+mpOP8sK3LzMPYO7LHdTWJruRgsRj5j8+4b7pf/o6G4dqY42yu1BilC++M2Xi
uWgEWeRhhGI0OC0BQZc1Pz28pDxyPnXsoGhAB6iigIEXofiA9qqE02xgBsSOJBLQ
QTttODMrAV9l8rv02TkPF2RAKIHi6jC9SFORnnmaf256O1PkmPVmqbF56DdDJPSs
0QNhLGrmNUyb0jAaxBihKZkLfw1j+NJI/5NSnm/EFiKdHuyRTKYdVEu02pf+i44h
eFQ3WBwNz9arMef9EaCpzhOD1ne/KEDo2gIhRPpx6F++BQDocVATs+y6y8p1AIpj
wgLZ5C+He7eH4Bu+A/tM9wuk1QeuHxmVvwkFy8+vfsPFLUZ/G93MKamEASaflKCB
nJ+x6oWkoprUpGAf6vZe+e6HPChf+aox5NTSs/SucUa/qrS7fvgdWNjxOBqIo/kH
4qiam0Ww7Q/PWXAvEFd9nSJO5xxjLt5s5Lp7+tPSU+K80ZPlcPYqNdjj1VKSQDbC
C7hhY/k5ycwssyCWXhAn7TEzEbwf7r+6j2fRDd4wX0rVqO3u/4ND3YdalTODhu+5
BcVnJJQc/Z8JGEH5Fw4P05S/ml5FltVt82bI/NTYTeG/VKyOwFSKU4R3S00r7ZFg
Bg3/47VtsBmi+iZu0kPrwcREppHwLZ/EhuE7nDgscbZSJwPvhpkVMcpikHXPr2Xz
K+GlNdwuMIjB9lFOlF/SED//Y/Io/Rb4MQT1dS0MnPKWFTRI8ddq1dN2JHQlNkwk
kDo8PYhW0WfeOxbP4P/nfieMGDe2cGf5fA42DQZg8d+ziO+4TEacDr3uTGVg7nkE
nQCRMWTFC1Yu5MlmYdEsDpb5gwjfB41HZ4tWcgepUv5g8tHbjr1IHRQOqwk344ys
tI2w7g2uvVjCPhQJmhNsTEsh4TgMKquCg1Fzxw2zyM4eJ3Sc63W3h0sY0SZbDfd8
Zy5bi8llvAK8Pyf13AUE5ezjM6FxSWV8hbfZlFB2Q8ObYs9nzUf00DU0/8ArupWi
Lbuqqpy+luRfHXH7P1q8iMJhmMt/fmWsedf6ukcZokT2dfYCHhuBWTXj1PchQ4f5
dPwHKhEElRceXB0GYrO4RZaJVU73GpjvWm/qQ2VSgXSH/kNvvECe0L13Bsy6gqwy
BxPhKWuwVpc4KTuMmhm1yljlh5o2xKUwk22uo81un0tg8o5G6O6jo3zq2W/CTR/N
`protect END_PROTECTED
