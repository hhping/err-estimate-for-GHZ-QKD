`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oazYwJHOupnqbU6vL4jsVJr2l2gmV+MC8c+plvJZwyJd9+Z4scIqwjvTKz0DLiOX
mC1+RfX3E2SLqv3mOTjlSYbP4tupTpMAB5VdJWPRwJvmQNKx2j8RSnNBoYzA3ggG
V2LUiKwJRWfRW3yVuUd/UzfEHr79K0qMfPUabpmTqJLGyS/l4YH57eaRaYQzbi5P
6MjWWSpLT7ksdCvONQhh54rlfaSPi+VDVHUHkmhXTV5JQPHXutY5iSPmChx3eIKT
4IyP7aI0sQjGucIkbyFgZcr364wZUOEEx/VKJklUWcPznpiZCtBwwAqRm5n13h9u
Pt5kXECsoOmvRytFTMNGxVteWv1pGkQTFQk7R9U57bTI5n7BxRgCO8YPo/T7BjWt
PCBBpQ8yODVPPtsvMI6VNW0DAT4Z9hNiHEo+i5WyR+hjuyPHxpxnAbcK9G1cpOHd
2lucZ1d54LBGpmMnY+z7LZkXqRYouh4zC3rINh+uKV3EsD9oX/Yuld65xv84ywFY
X2KyV4Fy+fe36psvrE8RrFujoKJSc0qaGgHzdFByCZE6pyxxWBWMGOBU8/Ngu779
HXPf0eOT9l3xMNWrHepxAiL2QfSu/7SU3GWnVoTA8ekv01chqvJe+l+LCOLaRMCN
dL4KPQFogQgAdQn0qz8j8sNku4bdR6QzFXdSfAMJLN0lpW0KnIbbSIOu6ulMT2ok
C5MRKs2qdI78opXiqu/eo7GxIrieRZ+CEoYr3e5wCJ6ZwvsWRwUcEUBw3Q/CaV7Y
mkfPIHXqae0VFWO73doH77vKG+ltE+fthz6NK/Rcze9Rs37Gv7qEWxRWclCB3mSs
3gk1IXZyLkX9I5C287OaOexgYmEVkDKmF68F4cxoF5eFhydTTOKZsKMerDWPt5OA
5XmZxyI5kf6sj4R+iUu32ZPj4A3/Jdu+qqtS+IBdvf2yttoAGkBXuBuj82g16WZp
I+j1f9OztNvAXbSzyBWyYbxviQXV2yzwGqiQJ2nzqot7jY2IkBYEogxbpxSL1KZi
N74LpJvbQpQYfFo36SW9zEcXtOT2ndyq7FQcHOhw7CoTQTx0UMozJPs3RSj3OLlb
UEFZ1/BFrDBbODS/uyGubZ4Nz2QTXutXXPGQeO9Lt+JrCtcZ7q1WZfPhdma/wJeP
wbopSQDbE0ofkaogEoFu8P8n1oe5Hd6Wr91pctlWRLA9j9/VXu812cc4NTQtSuS2
xGhDrhBSXbW3gWj0CwEczoun2zDmSMl5e2giKuSZlu4D+WPYpN6aXasC2bLfFHQ/
ikS53beahRH6eWkLHRO8pE0mOTBzVWd6WUH6ykgMfKi09oxfvqMGISTck4ITF8wx
3TtxjDPNk/GMtPZx+NJmR/KgUFgj/q9akNDsJqSB+M5vgXBqiwob7nGxFkSoPg6h
8hx5o4C5m3UOzB0gxl4Miqw67LxoAbh1TrZOmqrgySLWoH8kE8Ek+KqWcpWkhC6V
rVM9bbbZglaTXxaWUgBfY0hGeO46oj2AYNQ6p2a9s9YIN+d+bCo0nCgodD/ms/N6
YJ+dsZw+OvA65XtxcoR4AwqoVQPeMpPFEoR1IG54eWNObvEX0P72Jju+DivoYfsW
qIBA9ED3pdA66alB8VodBGsnbTZQ8/OWAArbPy+BhAWXTfuIKEgjqCYzeaNlpNS8
3yPx+jF0lrtK5zRLfw1+PkQMARRliAV+yId+RDHuhwzz0mNtCdQdl1DUh/ANjRyY
V8qmekobLU9PHffRcO5fSSWalggyuQuGSTmT2yhTF2yo4Hr86m3j8BkfhKgGiZxk
aqTFyYbBWw98MU0ChbCIXH3GNHTmu2JZ7OxG3HBS/ON9nzwwViuKpRYJj6RsalDf
ueLdK8l20y8I9aQjUjFll5ATzHiT+YVDbSAjKBh9hPAzPecs+3V5J5sdQ+oykGjX
jbhBVgoOZk8o4vKn9CXirD7CCi8jF3ZAUMdK2NIEi5bXnTkRgPlDMDLm8kilh/eN
3w9OBEaCKFu2jxPyilpbcZx3mlA78yIF7UjvkNE0Pwv33m/4laHVP5dki5+pixuY
2qGQ2IIA/8s716heWalHstXonzABcIUxMSPSo8idO8OH+Rvr36PauUDGqJwpSarS
/WuiqAVaWHT5nkXEbSLnrVYBmIqxjkTqyGHrfSFMXNF5SK6s4tIrLkP+bLmotuDh
BEeqgPApjSQNPbsIh9mWjx9n76v8C1KHrhH+wCUrcib2/eVh9rONfuCtADFRQ4DM
kTCQAvgaEYRMsMaKzc7ZzpCTTdWvpXxG/q9y/idi4AnYkbiDfV/86+JsT4evDmjW
Icr7VB6L43c2uZSdI2s9zLIBL7WKXh9+/UVPJpGTIhiBGLAyfs8GLezixKfOCtsI
M1t947hZv/wI+9NxF8j/Qg8RrWBcusEuC/coorNyHQWKb+KMy5a2oK0YePJKIID4
Fc7MdMenEAaqg5LSXGCGY7IJarnPcXjtWbZTOHSwPbMRGhgwXksHld3v/5y4IUQo
WTYDu63j4wlkONfYzUtL9KEyljXUqJ76Dx60etWIaQddLw0E5mBnDE+xMhQoM4+N
3t/PrE9seA3S6cz8oP+6XMq+La4Opi3KpNjRMKx0UpTf1To8vj+ud8hcr12PVNzK
XYdCWj7gJt5m3jaNo0Dz7aukVxywl8rfURrd1Xadl33o5/Udj76lUChxQedNAdmi
RCPJNLVlgz0Yh3mKRJX3u43pb92Mfzc3ejrcFqwauvoYfoQVLN00esGW7dl03sy0
fihLKLdU/UI0FMG5C7kjszrV8XW5DTIbuvyanUAdUQ/++pYOHZBJLzBKQz2MAC75
2zzc4rg7rYXrfKe9haaMtDAkdOa4/ovfrKX8LP6SjEU8yfQBWWVfJmczKoyFUkaB
wr9dV+OqqfdjeqVQ6foz2gk08iGvOSHP9+CLWyQFgXj032U6aSpt+aoXNTmvju6f
30PIBadRS8MshxHPAeDhAg==
`protect END_PROTECTED
