`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/OiPSt7Vg0eiUaycmR92ytf8C38ljJuRn3Ntx9+tlvHH+3nhyPG0HFMPu+QF/Yp
HT1HoU53AJMlQIW56/MNJQGoxJ64UKbCCwNgc3dyaS2KlIzMW86jW793TUF4USFy
B6i/K0pMTLcZd5lshQaRuNbItMrmtYrCradhDP441BUnYlGXx7yGCxDKLF6rqdgc
OHdRXMw00MYaM3j9+M3AcqwiUkGmU0URS1erA6a0+0aFHRKOcgXzVsZzfwUsGkQQ
fbqexyxLS6WTTMETI4+WPEYyHlJqu6mHWa3t9nNgRm4XHQupVG3tBWUDgny5exJE
ue8XVgSjtTofD6s5p2/0j7Q3DBIQkq5r00/LwWCCyvUJJ0n9yVJAQBdRRIiE7gRu
wzb9EKcK2sjFAzjZOaAbs98nmQHXOhfc3qIffMM3vsihwxMNjUzWzBjS+GmM/xUn
hS/DbZmOlu68bhojTYPlZJ4WIaujUw/75wBR3aO1ks4oKFhd+6UcoCcohpAgY8vf
ZIDm09sFaSceP//cVR06fMO4ODq2kZmO9qlHnLXWtqzGELs9W3bvGjJ6Z36VtSkn
X7ZFnIMftXrwkWJi7bPR8RRckbeoNxbzsPdRgh3PfT0lu95zEt/3rR6yzIH6bEHq
Wq48drrlTTsev06aLa+Sui+7o5gvZdrL0jzD7QncG/t6ChlfHypkir77NzOL/cCt
yYe5nlR/+nO5ZLO/cDUljdnoSCp7UgpwMD1vpIqrg/Pw8SVgMXwqo2f9LQouXEi1
mzBZ2AEp9zHdjgYRxeLrzEtXIaUDuXms3GKJohdJRjnSQAJe+tbsUY2ls6NSVZpq
m7fh/KnCcVd1ZNRCODkRB6ALBQlFIeTUH1Wo0DCMiXpXXUhTgc+I9MTxOGS9GkQr
w6u2qmlPNnkRyaLsY14qJ5ad2ASiCDqHhogqp5vsJSW6tUB5UdZ/2nG09GUpB1OT
iw9F5XhJV4BcbobYBeI07gio7Astapt944yjcmI78vSHVspseef1uNfN8ba7o9KN
VdCFkEcrlZlB4tD1bfRLVRdN6mD6YnntTOMt8aBerM+outbgAiSccLYMxGO8fsIX
6DO4PrJua/R/PFLtqHH+W0KzqV1j7GTLASpirTtfNX2xgHzrb7aSszJQTLpu7Cxb
H/uy5voG3tuV8Qnt7IvYK6KgP0A4TOetMzDnsdZ+JzJeLfuQGMSxFi6yM6u0DEgY
dx/xDywnnEQjxT8O9xMmIIE1NC7YqukBAWYBWGRIXg6gwfehOtA/RSvBBl2DbSlm
BDxxZPToIDCj/wqc7VAbFGHxs36vZsjc2hFom8eDEsY=
`protect END_PROTECTED
