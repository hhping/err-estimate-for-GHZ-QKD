`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JOrKvRkorHNZnDKMv5ZLGM7jqhSywzuL/rWr0Y05okLO1znbw/lwDQxqNJIPEkvV
NvU1jz+IumEzMiUqDIQRqn3iNPi/a9itQ+4gc9N/cbjXSKZ5/DKF6+Oseu4aAlIE
yZuHPXsOgv8/YBcvp1Lv6ZJT4mo4aWgTe9JUIRwtkjerm2I/VdPIAYq0CW1c/sML
3RX4vA9735jChAEh2wlKtSL4SG7HuwLEVVabXOWCWhLd8egZeRq1ZxIdKIYHzgG+
FgdYkYWiXneqkzJOE7B7rC6MY2VZ9ZbIWV2FscimanS98b5iGorkgGhMMcDXE/EC
n2OngpRRJTzpKVhwakeCjXBcx5pX03Xq5qV82hB858QyyK/OX6BllGkkCO+1hSBJ
lx8hyNA18Rr6LaXElidxUJOa8U7NG4r2+474Jiu3/M0QPtGqAauwZdFc3JuwRSWj
fEWTd/+eFLhzx92Kt8rl9QUbS/5kiEVsVo1g0avUQyZNQWElZguTui9PqtORYQf8
pdbDO5dMvB6+FHq2fYJgdcOaem4aTRq3ce5qTYrUTfPP+apOi0+sUhI6CrqTy/6Q
u4QNt/skjDJoAZxAOULuEExg6VYZwJYYvtpGfNPD8SO4Q5p45Lv3IDtMQ9vR/bwp
dHyLJVpZt4TtCbtzN7Ahh+VBoSjPkxQuft2oXGSWKsf7fjrZsBjOUDQUhxTWgHyC
gwrStV3wbasbnNIML6qpj0TuhDhMBUe/Gg0aFa9zAg96exnLKgN4qQhqE8vzG+in
Iw79N2IDYB00Ywr83n5Bes2TPEyZiQyupwtOKUvOX8t+pKPiu1J028kNfi04vaph
ILdIZzxM8BGqWmTJEGv08KZyiwGvPeyA6HrQngSaho/cTDovNZlfB2zk0tCqRiQI
rRXszmKMvfuAZPNQBwBBzGz8IFCxs1TI3tgAEwpvATvmgvCkllbYliM5E2Vtmbdu
iTUoTFO8QzRyHuezoJwgelm9udxHVncuty4t2TMcx0QDJF/yEkqHarip9+FGZ3hb
K0fFvAPtNai74j0PhNDO5CNkbkay6U65/ZFdBjbFK+kQMDOzMw5rLX4LecKK3JaL
Kgwp6743O6I/frujwRHN7A==
`protect END_PROTECTED
