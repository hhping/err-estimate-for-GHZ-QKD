`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzUjeyJZ4A3MPN3h4YvIpxzdhvVx1eSP/2KfF8JHrspn+V0UUkb4aYA9Z5ab6nu1
d2U1CkpQef7jY0QsJni8avJg4MQ3ze+UjOkfUhts3m2ifo9CFXlW6Zx7WhVQjIaD
wgVdZEDV0ML5UYqCuyo96fyWoPSkBOKs+9+o/4ZQ+uGmlHoVC32B3sbXZ9zKmFtM
1njwgR48cAWsSJHXlw26/w5veNkqUo9l+tUrcjeHWztF8RsF8FEzSmzPPbTTb5Dg
5wzCF8gSasORfK94w/K+e3YrmN5+Gek7XJmOrE3O5Npy7kWiQvo5pkxtnjWDjWbp
qJWFuQEtxn03ZYpBaVOmvm1I4OQUoVQspE3jnZCIpIk/5VXA/5uYZwx6oX6Jls6w
cv3jIrYKRgsAUge3ccwShy+r9oWo10/YR7z3lJxoKMaz8ndCDBx2LP866/abXYjc
Ka/Nm9UqJzj8YF8CGqe+KS9rYVCZIfLEHi5/BThxTT8tA3adyKpNkIsP8JazJmsH
lr0ieXD4tCIeJPatIcg2do3ufplwMU+1XxEh2RgCNAaq+FVldm1GI+5vMkSToznJ
2cLb+woydIwWRlBrN+x7E8G9kelExYa7VF0C3kzIHH2lAA0E3UpYJxrVCg55NvOv
y9gOAwFipMkqc2oNgHGOUduJO6s1nvtfGPEpCAmMiNtiMN/Xlec8Blb1KYRmy08V
2AJQM/1QD/VBYD+p4RA7YhMHNOahXOg+ybpwCdiBE8PcLrt6U4vhKv8dEFsggjCU
TCIZmKXRejF6UPtf6Hqs+3TkTACBFP4Xsv2ZV3kWUsbBx8JakGURQo9AICmnuUr8
vZBhvMp7WAOuwg9hgHyY56aBdJ7e5ewUdN2UNWlyAoKFDhBsZDwl6nQ5m7bQRF9C
fTeZG6kb5rvxg/uBDfBKB5BWwhuWg8M11sd35kJF7U1v+hKAit3LztXv4QIxIM1q
MvaEbRLhDExmIhJMT4kdReN9K6Dwc5MJqI4GfcgirWe6OcINwMg/9VT5+TMdGmpC
TlPnkhXi7CjQXcZfWZInHI6Rh4rHafp9ihAzpIhPjVMOFQ4bq/Eley5ibSmOP49W
5HQiZH0UIZ0caHpXQ/BKY7r/9z0SuqeHeW0lfX/AHyPppUmP3akCfbBrjiQX8Lap
`protect END_PROTECTED
