`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zfLlOqFuGqgV6gFYXHF1/Z93H0LJz8Xe3ab4luxU9bWriV0gMGwFT/rXAPKY/MZU
Vb7smzuiu9dpgo3Y+ji+NOT17c/mhOcqjmEk31j5JDmJfynO6UC+aamGKsgDWtc8
zMsTD61672PanVRtddif9uW2ziMuF+sbhAzERdKA0fn6q8fiI6TfQ8qpNrj9nzUR
mUhxhH9d8D6x3S/nhiDgrFLNiTU93fszXWLlrAggV4/ykhtDIlJHkgy4R5UNV44J
ZT5CTi96J74ogTEhDshbavGYCrmTreJ5JmBoE+5MRvmP+8iDxJUCwQDUrTrJ6xid
8n2zdoLnpzAwI5ne7j9dbQ3t+R4Y5t6TL03IzgPvAbuduTPJEWBaOTJQ5VAIYY3B
NTXR26lTavL2tC3hpB9ybZYFX19yiHA1cTs3jHnXe/HP4U+FHaBApeGAxRNbPAqb
7gtIcnfFJBs6Qvtz+Iw0fFtztctEOoSuBMW8lxQmmTgnuMG7NLHzZfrYI2LAF0pk
U+DktHouR4GIfKG9MGQJhUl3+nOiBvnDCxWHIEx/E5175zttCR8iIA5LWeASSCsD
/LSpqTT+41v9WcWEA/xlGniF9GXS7jmuTpKvvi/B2+/31q+0vqIHpLkTt1YqoigC
WH6MRJpgpxH+JFkjTa+H697axzJsfMDRnyBacUrfjzNH2ABataPEidvsTOwp1Idp
D865B96qB0A9FLzel6i3ZiKUk9fYtBTFr0UFPUieNcGZf1rmqOv36HYbrnw26vNp
TguG1VAoY28Ac2NuP5cgYvp/O7+1iXJUAuRX8Uv+VLt/3YSWr7GvRl12ieI8Lhna
xpz0hS2JCtNl7k25d8Ud7h+OgxvnMEaP49auRCNhi2tSQaSL83/5Ndgx8gPhYslD
jrEkyWOLrFBtMBme0d9BCNpJFsG3Fdrvp/S18nFGvYn5xaHQ1L7nE0SAxb15XM1i
jvgJ5QwBAX/tNA0Za0Ds8KaFK2joQMVvOe8GMwWF5fjtGHUjQot3fukn41CBS9RE
80fIs2MkZLoUyGPK36d2Lg==
`protect END_PROTECTED
