`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFv0o81JgGZjibgTyS2ZtycS0bCQBRdIvuk0GGcmpGt1ZxpPUSn9Jda2wcZbg9gG
VgJ4nq383PPdiTXG0vi5zGOtANA1/QahU+yf0tOCMbOY3G/LSNqplG8cYU9kocSI
S3hp0qcon407CYSmTeGl3WZVedhcJMBfXpkGxqZd/5inbTzRWN73JMv/1gDmUF63
MJ9BG06RzqmImKz98dcr+mU7fate9kTQfTeMOX6npt206Tw1sYHNNzApKQvfE0kF
iFYMD24RdQcuvMvv599+9sNw1TiAzZvxIZ6jLZ24q9GxKeDI3Sm7pTfLApN24bEG
nd9vDE8W5ECMuPE8VQdbiOIBooT6M5dmhaQS/+kOrxhJDhLtIXV6jvRKgUN5WLmm
dFoF1vUJRetdwLdiK/Vi7QmqMFKH3aU5roejl3CYN09b3BGmn7WMnm5DnVVdJleu
/MB2jaypMQDOdSFL1lIVkw==
`protect END_PROTECTED
