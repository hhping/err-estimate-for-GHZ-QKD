`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQx+EJ2xPbEc1f/M/089AQuKqUN6yIRC3XoF/cYU0CtDdeEZJfz4cj9DThGyGvEh
xQHE0m+tGTzLlOzz+fwH1hM6aZOnJCfu7ISJZGhEs+Q3+EXOSzbGiDFdiU5zB69T
9TofWtX56io1yY3uS+5XuXFVP4jHFFkm5+jykjNlJ6YJZntq9hg83Yyctdav/zeA
x7JqWekbtsq2U7wgJbNolIb6wBQ70Whb6xVxTPwKxLrdKQVZ40Vc2OMckUufOcHG
RnH+8J1bhOcymNF8aptDhZBd1DCxErGfxAfKI8JdJIaI3uk0PTwm+26Sy4qw+GWr
Lvqa8pk7oFVM8mliYKqnXfSjSsKSntUHNYPd24OFVyz4qD09E0DP+eJZFm7iHFe5
Ygwo62e4OwdXiXmWOATJRH4678RgmsxaYDnzHAyMNW6bcojHJZDPQGHauYUToh9V
W0YOVdy06ynh3Z21BQWE91naJy4spEB0JgDT2uAMvkqqA4BPFO1lkomar/5MQ+jd
9xP7EDM4HHECBhnN1/fMhREVpWo4FVvDn3qJC+E2YQW/VGireUnERK+P1Q1Jt95t
y8H9T8n/V0+lC3jhV5nx5Zez03mlns1jUfTLcF/YYzaIrdP43yT5gI9Dog8tSsx2
fRBtf41PQLFMPX2G4OUoX3laaeU1jASCiSGehhnIQ0lkl1mb4ftdP7yHQ4l3jayK
LxFW1jMSL0djSKRnMQg39/lBwA4DERA+RWHQH4e8fInGEqLGdxWAkDRAE8mZ3yGK
+AkgTrVDr0nsVjP0B1A3KzrVRPmbhp5iV6E3q9REjNasjcPQgrVmUVbT0EZjm/6P
9yQwBqARw55qdiTboLecdE3elo2FinEdvfuG3ffCaw/4v3KXkDPvBZijTjFNt7gD
GIWiXM7DjgZMDkGDbeW3wOAOUdjLQiqv6w9/kXUM8bIzCzktUwFo0NuctmEMZZ4q
v/B7jqGJ2Kf6lzMSJYqPoc5jk/qGgW8i7aFSRRyyADQPiMuTsiP2q/r3vlUa6U/b
n9jdeYvl36NwdzQCbRzdeinhjQojz0fKOlJP50mG6onE7Htan+dXrdyH0D+X19xp
551Q6XJYmOFzRPWZMGGuctWRUWoLeXM55ZG5wwS/qMzmGTNvQwxb4ABiZ86oKLsk
3CPNH0o4VwDt4ww6dO6IskZ1HbWElMetz82lOMKFOw5YQmvHysL6dV+KSPTVvLg3
76U5Zc0PKBiBt277KQq/CnBL4HrVBFepNqmZw+8mciM=
`protect END_PROTECTED
