`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYbc2uahBbHaj9suz9U1DOQzc2vXclEm0BfDkR0UiPAY8LnRe6QoQ8kBKhb8l92W
BovH+iNSMeZWod5h8FBEUjZMTomspqVp3lA9/kQIjifFspp1kiABlyVmS5xHMojX
54wQrPpFPVKKT0bjIgYym58fCBKVq5rxCLi6DDlAegra9nqGcSph59ldxUk5Yiyb
zQjlHG4Lsu1heKw5OuoV+tBxSIvDULxt6YS+a85OfppeKdqbBqwP6LXK/9hvbNqJ
LBwKXiVL2B7HpOICN9/5pX3GsOocNFh/T+HH9p0P5RhW7j/U2wa+6eZi0vd+iTec
Vs1Pxgj+HVHYNXTiRHHAmLFX4HHp7rkwfwDvJn2zXBTI2PxhtcCGD5C4jqBAq5DQ
2I1EApaWumCECtvGhR4ltSWtvWATBeAVEylZ0NynsnnzCAJtvHpamooDSp0Oxswr
JNideW4NkxQsokxnSdVro6tVWF1qLfxn6xuxPhr+FMA=
`protect END_PROTECTED
