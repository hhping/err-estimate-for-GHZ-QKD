`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXxVZUYmYCRC8QRHFxyjPYmLQPvc+cTMraTN8nqN/5Gz2bvDv5KPW9A1eCwII05e
svOlkJIBqbguUkoljuNeLM6/7qXP1FiW/c63MQtu1dR7n5lAF5p74iVsaLyG+uWv
yJE7zf4CSxan1OMjvpzsg0jqTcw/NyngvQWqYuLHK08w3po57ec/VCbVCe+uh8wk
I1BHSl3Eg3JQ+BVZIYtrO+GfkckEw0gtUO6LZqcdsc+qMsGOYjIOodJsgEtuRXNY
rBgrl3qEcxDk1kVvc/tdpTAuQIiIUSXTXp3FtLLfC5eR+KHjfz4IdKc2gr6s5pZn
bYooZtGKUJ8U0X+WbyiEpAJz08YEFPmiWO72Phq3ox0zSYGtgl+pLQnZ5RPMP3mY
OMl15j8qusA94riB+F4I8Kdh4vnhh8Q8uzie/VTVzcJ37X+R7F71iMSdn8t4JF34
PNb1lAReQewjR2o6eE+WIx7yYrbXkotQoQ3av/ySH3Ae9Gxwbb3Au0xYOMbxOhzw
0tnRpy9ZvJQZKhQ9b+q02OlTg/yTcBtJI4zapHZAzaHEdCjT5bl0b2O/eYYLQLk9
tztfqBC1d8fVTHzY3i9l8u0c9t4HGVgssmlU9sE/SwKw1D+qtDd5M0MBHt/Lxb31
gMMqa2UfeE9p3UJBlqTrJHGX+dmybOhehad7woMn2vBEPXsj5ITrQv3RQl4Mav82
WnE4GI2UfBprLWHZTGc8sklI5TSwlkHC4/V2uX+Mb1qHwUpIN5KrfbiM6qNBTLks
PZXMZY08pjo3P2IlRnxMH4XLSVL6tzl6FqkVGJurdGhszbCWqDIoUINhF6yYutww
s+GiWowHng7h39FC8jxxYjwoaH1u654rCe23Ivr7iA71BUJTLLxzgn9iUQUMbMj9
bZU5HXksuxlW+pDFkvaenpaWS7KruH26eQa/nTYgOIotPMTaQSdhE3fM1BymD0mR
Q/th0VPiGg67SLehn4GmnuJVou1hosN5ku7PXm7f2LB0wOy4RHc+GQEjut8gq86U
CfN8sYOCTU7d5J/xN3OKew6rFjpQxk6WP8lSoE12XNYma1wm+3rXDQceAChB5gep
ZU8V90x5egfpY/sZ92wU7TD0MLMCMZcUSazS/rfzNAJjZclti7z0SNVMyH0kfJvP
Nsin0KcPtd4pHeWUTIDiWSSsEeJp4/qQuQqIqKbCFYR7xqxv+oy41m/4UEgrTp3j
ANnfMrxWgFBelL0DA1fjqiDxqIe74WajrUcWat5ahbdkiGccY031FKzEm9v3SiEW
nPYoKyr9e5oEEi5KpJeoWXmmmBhmYcXNvkEZO16cfa6kwLnegVFZLxc+IrpRakes
E/yE2o94OJtF2/rGExg0mh/dzjn11FKuhIZrutHlQ+F++HOLNZrrSg/Ci9K50Dxz
TpYIKLMeDUUS5u8eO/h6zhLzJk5uWtatF6cGOFLRKqSrzSBPdqBBSOHgjl9E0+Zg
zIGQL1h+mzChmiduLmLgiC2oW4z9LPCKCEJeAFVep2NsUwyZYK5+wJJqUkQNfGS5
2AwOA1EA0VU7JYN/lxforLT3yHlz6rqYxDHTi8wCqnDR9ESYJQJlfgPApqKpU8Wu
vaj4AAUGBZxW1OkMlGU1MW7A+BcYsvlxhHK4X3cHqsJzyjAVQlPR5Gyx5UgdnrOC
l6Moj98kJoFdIzqjCZWsBbLR/x1arSlV9ZnbJ9LGhFkqmo7vk2BrQGWdpFbdyU7J
BiDjU9bWY8kV5emjTJ7dR+nr8WJ7Mb0R78qAIJa6yY4kpsYt3duHK+8F2uqqFJKj
bWX1c+U3jXag6nNLi2WXWFT9X47+hvQVAAQvaaLSfdC4nx2+x7cb6RG8y+kOs9XN
2EWkOYzFSCWbXu6zdNKmCmefQcZ9mTKQn19xbBcJcjQ9W/4q8bckxtCZ2aueddKz
6yH9Gty3fmAGq4mLMbSbGgSVNWn0XWUtGS0pwE6LZKki6piqtWvWkv+CyaFrS1AK
xVcFXn7sWawwE0O+8/q+pDqX7GvPiU+Sig3TtnHYRU99xCj4DZc62Vf0YoeoxFIM
+MPVgtJG3OwqzJQn71G+MXT1d25+mLTGbJISE5XWD4/Elz4gzYQ0et/2csUvMNRk
Z0NqtCXmGqWbMBvdTCG/O61BPHAk+wC2s1XqtsP88j6yKW/e+DsfOEb/cjdP03bU
QehU1ywGh9HqLd9nRjJ7qAHgrz73HmZ5UMqfCM9X9IXYmXNjmYjU8wT98hqDwzVk
aAFMUklHCP3it7mdcOJkia9UcXYZes5Vko7te1ldkD/SipMggX9zMwiPxdG0DVRt
vf5GlkKIAPWUtdB3v07OQubASOMcRPPAc7Q3NAODcGxAX+b22m/NJXuURHB6B/OI
dyh+2QhXtcmEBeb3N6S+uru8s1mSapceQEwqfmHsnikkbEogE2AckRs73RlqdwhV
CmhcvxethL4lW6ufAD/GjLLfpGVQRxEvGpDY9Tg3nUWiKoF7c6MuAscZhPD6PRcp
vfFqzngkZmNSHRXvZvKJy8Y5nHI1wceysSQbZ4o+VIStzBzcdQMNOm+1L30fdYVg
NE/JNcbl1NNlGqzlkqQ2lpYROnJhlJCFMG2TvCB6Niuxe1zd2lqzhnEwVVUviYd3
+lNeKuNMkK2A6oHzaVqNqvg2UPB3NC4aLXuCUYyHtmuY+dt5yagAhU/z0wnkekRH
CiDDVD5by5CBoZTUROhhxs5iWYE5918RRifpepTPGfIZFkWmcuMDQS0rQCBlN38M
DM8AQjz5hFztrMv4QTMUhaxk0wHj+RH2wpaJzkl8+8HCzvkDoiLLJLqQk9DHxwfx
piub87IGADS1l7VjcBYfy4MzMYGQJ1uSgK17FLyIV9cS28SLL+22BEXnV7K3RehM
cYVlALPaxWid1QpH62xrFspJXCmLyWU5/0lR1imkOCJ6kfvBiaatpsUCTFNA1qoM
7wC1NVF0bNbV9Da37Xe+w9JH+7HbAYuqSmp9vldOzbBnS7Oyc+XmP5BnBFT/pOVM
jLDewDDTCB4Zf/pyyBxo29ERe3m7bqg4YQV/VwZqhqJauKfTFal66l8WSbki2B70
ZJE9xM4R3NB/+e/ljGvbw7+V9nlfDvOC0uENlg7GPUrc86Hgolfy25k0QG21n7Z2
hLphAMILe0P943UTVZd4B1Y1fk4HPZbVuXu4H6g8INlDutBZNw2+rSVG/WePXjbv
T4C7kP6sb7V3LNucoX3UrW31TvIOTI0VlNsHsaGbfrFFNrdMqFsCRfoBy/+bDSyi
IEngmcKqbNqjYrz3tGtTGU/+5mOjatlUoiKgziDcZOVYhApMyU6LRWv8b6FzKO/S
0DzqK492V4iJ3hlmM6YB7iZJnJN+d6DuU6nvz39RNvw/KRhWjt8weYZNxW600bEz
syBM7O/ZRadm8PiLBPhKYkoAtjmTPbl3oDpxIGV7gFkdvld48aP7ArlwajyLrJ7v
K+lSJHm7Gm5PVt/fP48RFn2otYtnjC1XEhnhpYVuGO0ukspPw0x7uP+TRvW3m9IT
i7YgKK8AWapUwtApfkbrFtik89rrY9ZFQpZVgh5ZRsfeCqWLY0LdxI80b2NAKrpW
7Mit5tPQeAdbtrPW1QnQ0lGRj6oL31E5VqQwJpjaKtlgLBHPwG4xGU2dlEfdPgI6
m+5Ek2eM3xn1iW5ckiF5e1+3F7zVhB/YLx1eLnL3jn2AG7ctZ18b+Ov6s2hLbhOw
HR9toyzCUCPbKVo2XjmNN6oYWnNixN1JVjenfAhm4X5RTnYm80msvpvdhSJ1dh0M
WER1t+rGGCfQcpLjmF5o+EGVb0QPDlIMxv+N1j0TWbp0nGjOd+yneJVU1lQLwdF3
zmG1AriuqQ00Aewe59233Ge7P8DFU+LJfHz3T/bPBl6unjnpq3oTFbWvFBWLhAHl
tVJXc7yW3Ql5CuI1G6Mm3ksf2cPpUwt/30qG4iM489zzXek+aa09oamijlbHAD1F
HJIMRFklOfH9JnKxNx5dgodcvS2EVnVORH70hGzJoIKdEkAZ2Ce6keicnEknGKFy
N+tQqkZ31WgZrhIUmnf51TPFdVDa1t88kSF2qOf4Pq+3tMytPGFlehPdvI6niJeC
hxvXjdyEr8EGamPmYHjX2yFa3lEasvbtjOcWVL0ATAW3gwOmrrVwLR0lex5UC7AE
JBcXgjhBRp/k5jYk0xikjqTmXTBns07Q8Ql3Ujg0hQLaLGK4NP6D76Lelqt6OIi6
yGlFZ5w2KJM7SuOrPAyyFQvFlVHrnAKlpCtl5aLTXDQ4u5hc/Lvu1Sat9tOvR52p
XiVNtzkalpPkgBdJpe5lCbpo4Hu8WV3pmn51vfcKKM9aQ7WYQRnkD84gdoMIbo7Y
OB+WjdS6iRWEud3HsHhwQQREO+9VcdEeUupXMAYx+0ZK6JWYJxAN1WuJrc0VIvo2
BgqBTzFr23nIlk2gbua4KxjJGOtgLxCX3o55xoTBvjKMuI2jV83WV7qPAj3owRtr
WvGZcVfZh2weNmV524E4Szt+4ZXJYLChDeYi3oqtwKhvwyLAWtzlBAj+imSfB08p
Mq+1pJ/o1lpVPDKNvP9PUIiJkjwI2wk8T413m5WkqMlwZ8kSlnTobed+nFWam8f/
GOmJHgpXydkNezkxztH58UVPgROrEiLbnnH7H6B/cvR6mQzybBmuOZ9W16KLjixG
OmZ1r2cl2JmZH7pi4G/kCZr2rdHXDSoczRGd2VA7sNfq9wDgkDYQjOcJXccRsicO
tvZhsvy3PTQ/cUacNND0911MabsH/V/SNSuci8dvccItD1qMuNYLQzas+oUNv2OT
hiYkuDRjCzm8d4ozPEwVlyYXJFaqVeE1Jb12WanDGQ7bRKMHESV9Bw7tdV8+rHue
pMiZeU2krzRAPnFtihPvAmj3YiJ/LgKcbIarB4xB92c/1EihTbtHh9BjpC2NLm3H
lPwpym8BjHcljvNTz1KmzmKLx0cwRQIT/PoQN6VdqE8i3POB+t4ohNekO0rwqFLf
LxN50nlPMEpdwtHzsXLEIRh3nHjR5pTMiH6ChvPNB1LZVrLpFHT8Yq2VetTNnNJ9
HRUozPBt3z7USoncKMziqnsE1T3tllaIdUA57tZieE+u9h3IYTmPhYhaonrQNZj2
i6+OPafttbQWdovPgIAYRkFiPJqWiAnlB0pLv2PiNRwLnu4qExOQ3KjKhL/tej3n
reIO+zcRlwdbcpaIrCgpdxEibKcG7xn1chMHmW/AIXVXvvsKakCesvpmDh7wPEnb
62tnRkZHObP2u7Nv2wUnjdUUrQ843TODNIkeUMIz8fo0N5HawFOQMWPKrNvKbZKV
CkbrGqkvXja1PAhjqZpnsXuXOgfn1tHjElx7ZVUy0pmVWjenVZW9pV2E0oAXt47K
oi1QEqFZE/Z/qitnBJRH3lD7sCrfbOU3D21ejbqs0BqjfrD4tRdIE3lhyFIvQlow
i1IQOVH5zfzUkYGXC0n5LOYfLXON6QNnUUr77tLx2NH+MUhiGK6DtUqlQcYfDdGh
46xXcUwor4MeylyNy+HUaf4Yt8K2qV+vYE2GsQo6+O7Db7rqnX60EbO6rcpWHiMu
o6BAchkBhR61FOY+kTLTXtVj8dtfHcH9pQveTT4xVwrh3a9Kan22moFIwLRlNFvs
CPp5PkNVDGmawB0I3bkUav2AIFO6evV6OaqqDllI6VaW9cUzcQaolu/D+RtfTX2Y
MKTi7/jaEaKCx4F4wW+YtOfBb97w+z0boqwD+YHnhwh2yvl7D80YPX5mvgppE6re
3ezBLjjAz/EVaSj/HUNLBnyTOvKKu9jPgJcyODfLmLD6qpBb03Rc1T8qYESQEgYY
WIiWllvKOwt8Z9SGVfHo08jME2UGp8bL8pHCzNq+3DdSjIwDOnVIdLh28F8YQE4v
gGQwOur7S1uiOk6aI9rMPLGG9ubANYD9M2r6s1bBtSsqJh54jAy5mIZTJICmb9jt
yE76+6WqYtVQwEojaaBh2wkTDwDxf0hnTFjW6UEZIhbGoWbhX7JSCyJ8T8/m/BKn
lis8L9VAjsgQgsCMPF+KI2El7RGzAyVPBwQ6AuGafg+M0u9gzEbYZeNQTWlJX4GY
pkGdlFx2RZu6khipLadtVC1Dq3kjev+B4hv1CAe4+ieXM9vlSEA+r61EzonY2dDh
HHCmQk03WwriGR1exj1CSD9guwjD2d6WmC6YY+rE7qElL+3P2Mrx8Lh7cyowruGH
RiTFaDeH9w9v5mmsBHbx/eeuL+3soRJiYtZiMR3KMMlDzlItgb9RGxiXQuca4IR1
QFwEeoFOn0vNphf5Eug0ura5vS1ha+CSFa9cnnSCrwcjYUnS7FmhyKXFmZlqat1m
8133W+uIDEna3T76rtdftYdr9melwEI2xs4NpjQYG/pcp//KYMXEZA4RIMdzhxQP
NbhdpnHySHF9NgGN3naSYogSXVV67/0yaJXKyDzKUKn46DbPKOo3KA6r3mY1M2ky
9IIBqQEf+p4C6H2K0IQELYkhnHpI9Vf8nLyjl5zuSPBZYtVlXkwwMKbNXoqQEApn
5mMxUaU2U+HALmmhEFK3JfZcfdsXX55haU2xRUiGg4JwNnZlAJIiFcCm9BRlfGLV
8piSotg9/F/Cq1PIe0jvih335oekoncxdH/2wjK2G9EhQZRaL1KgJpGyw27j45ex
cfwzBvCFf3v0LMzFQ7YhjiW6V9f/8W9hVCWCWLFxuFGuPQV4GDtTAqQkekqCJlLM
nJid4IOJaaZATZWNXwFNBKkm+6Xuf99gEgol0M+77fwP9jEZRBwviPV66FR80jNk
hCVhcg/ebVXiTfZMF29f0mXKGpFNX2yo6LKlMru4C57H3QsNEMJE2p94r0NhQ1la
czG/gH31bc4IpM+Os/vqT1eNdMdTVIc5E0s5rDp2wb5kAmcQ0ubNand90taL5hQD
WTuMQ8UAduZ8YxO52+413VV0shjHJGsZa/HS08bDPqoZGfWEztUKGWPVy5upvJ4s
hEue7qIq+Dc1KSzYBeEThDjs3OCPPWb1xrR5SgfsNKWh1c6q6aDdbMgcsilyYsxs
dJu7mT56DCQy9di57l05hQbmN1RPykONt9TnZOybD4fCebjiLdPtF78LwBDEpXny
DwtgO/Y/2kSajdF/RO+v6o3IwFidZ0Fj4hawpgvTQxK1pxFEU3jipMCnPEFIrO0p
/no1iG0BhabZ7auG/VBqziPvd310gj0tta2Phe3Za1lK0pDu6fFeYEXDMzhm5V3C
iV828X30OKJuhjq1AgxX+oqwvPtUrmrAk070tS9bD/ntVaVlr4AK1mq8F9nYYfVW
N6ZbTVluhqlpV2UOJXTN9gTlPQfe+cMeZ/JBjfyZxI3+hXSDWG9rO/dux2ktw4lO
3LkujD4HDqWNM+3gLsyYhZrXZ1HJFj97gr6LS5GTPlkJL9WHgSfD7wf1NJjcIJsv
AhyDCvy+kuZFIJL4H/c773dMkFYBlXrOSKN8IgpxtIXY9Zg2pWrXSk/dImy0xG5q
8hcgolO3knsUF1fuL5hCo5DoWpo0dvnPVQYnpsgKE/1ux1sHfUqCsS2XPi6YcoZD
pIf2PulcjcU01FEdC8JXQK55O0+As9Mvb58sc2Yc8JdMCgWai4IUDnEkE/DAyJ5r
zrlUBpFLJE9gSicrPrg0Et1rU6+INk6CGeAYIpXuMJiZAtY5ZWodcpMxFCh1fhnd
AVVkFj1oeYzyH1ySM+ezmYqXt3+GDQo1ad9p81I7YynAN665iLJ8lDyfYJJSLa4I
SjnBOqw5d5FQEDYf3s9ZswoLeFNqi8+5EiERCuakm0mBOxJ5RSTwHwB5G6BWEcLt
hfJHaY3V3b6R/uU1M0pc0QQ72IQ7IqW5FCaUZfqZazmZCEUD/9XbpoaqAc6+lZVy
dyjK3nVEpabVQZEA+RZzBou2f9+K3ALY7j3gaK1hldjSakT6BZFpFXqZrzxWiTfL
3Yu/Dokh0hpp5CwSOYto3SzLUaovS4JMtmv1SRd7Gu1b/ZqJX1G+BAomiwzj/LD0
hAiLoQ3Q2swS2hGn1j9cMufpiJgett325cfO9J17UajNEJYfGom7i/cVxUFfDlne
hjLcj6joa6ipcz8Znci2TRcS7qDR9HDR6yed84zgLF9x/HHdnoPt0BQ1OoHZn4KT
QTVxa1O/HhmXU5aZOxwenTbM7YJjGLK/VXuBAnCcMeIqa86aR5FG8hgIuXlXlfzI
diqOzHsrbyTIRcfmItYJYfjmhX9Z5mzC20kaHRlDWAzONKfdBqV+eNbco/VvkzMA
DoRbG4ts5KmeVKLAff0ltNTwQMczovASXSkmu7gh9f89/kIGL3TgOkTCc0oq6XvX
6U/N0mCD61fSKTBnCaWmnNerk4rs9PMNf7ioFeK339q+vrD5xyrykyq9gUUwUg2j
V5f+XvMCWr6I+1lSlGMqiUSwhIB7NWQ6AGipSRiZZdV/UgbsE/rkLtvaCL94c0Tt
DoxiDYSFM63pzgQnz43G+u5mE8XXAPk8ew72I/aaKb4UAxEgZ8sVusvxgyZJ9KJP
Owulors/JQSd2ZP6Yo/yM3MeGSo+f6EsZWJXQdRNurSKCtTclorkWMKw4DFZHVsn
gJlRzfKKG5rWX1FFV/8TnIcug7bWFybPvb8aT/FJ8HyWO6kGEsPKthEhtdVxIpeb
skoBWQj9/1OjKgT2QfmBEZ9+yayjZeuV42blx+b/8yp5jsGqlGuIbzc+8y52sJxc
B0ep/6I+Odbu1s8wKAg/palhfZqrRDTHRsCW+IZ7FgsUng1WsB9G7Mbh73NeYcOo
TwTUGmnbrWS3VLtzQskSNuTRKfU5FsG+uNv8slw3ns8f3zHo5YH4fNU0WsrVyTYZ
fWlc7L6T2v0IPRuT6yJwzVI9z30c4sioaLlhJg7Ik6zcYLk8RIKKSWPcnacb/0AL
hnx0N0+QsmlTfNlwX21aSecOcxMJjVCyavxgpLu/A1f9u4gepA0nrHM3torfYx/K
HV7lj/J/AgVqiZObQ9Ge1Qq3JI5BKrQ/cJpJ8W3Q2n/DUpF01tb9iz8Hw0Xi/aZn
dHQFDuc47F7EVt4IwnTIYnz6t9B/dA+07DG8tWOVuWJ7aVAJQCWnZpHJh0fDnOwe
+bDLpT1prmpFNPwj1cHn5GbMXXJslqTXuiNwdqQGf7nY8Lbs1UfVQhnlBi1ajQ1d
mGX5NYhdKKHeX1jyq1s+RIkA8Joe5jbh78rm85nGKbyxFhogv+0w4DXCEfZ+EIOA
+M3j58CAlVNyJZ2WjYncbt/UKnrg5DyMcIzTbHCVAdxfuzUYd+IDq22vTs4v8FPQ
kME06K7nJXvAAS85FuqhMB+6+ZScL/qfxFVhaMvqYeEGS8fYSMWdJ7u2qlDVFHMd
nRgddvEyiUSLtYL+hCpNiHGfyQyjtPjFmZCqysCa1TJLIMKYl5ZPk831PrVp3C7c
AqR287uVmXYogofg4dqSSV2XHdORzeDwBaqGY5d360MtxPt3H38S9uwBahpZT4L0
H0UGGmdCXIDMaZfQtqHl4lZH1HE0WdoGfHLB7c43Fe9erOquHrnRW4y6jBhee/DM
qCx7FbSX+gXtZOlVGFAxC4vMn1PaiAEPDNSaLt+UnvGHB+qEsDvjP8eDsgcDO1Zq
cuCEqSIuXN4Cr5tbjAg9fX8a2iQliStxvQzX0wPxbTKEt1t3SdF4E2jZMveEhNAa
FkTqG4Jm71z1w4w2BkynPuigvk6rxrQ4eDCI5m0kCn0YYtSIaE0AX4VRgvg3OmfZ
7w2b/92x4aVOq/HBpEqKPeV6fi20tEEXZ1dxYgBkm/+sRayBnKJUkc+sORTvUkT9
4qPus/x4zqgXcIFaX6QU2OWBxOS9Ct/lRiKe5H5y6uqi9qSfvxS63iqa3xrpiCP+
tdxaLuW7lZQY9lycvWhrrnkx/vzw+qacl65Nzsl7JQ3+fXolSErlmISyJEuZ7g1W
Lr2NmjAll35QHZFhMufMzl7W3o3+yO8itjYtuzNy9eNmaovJU0/V2LLET3IUOvqB
3qxlSYU+CmMioZsgzI8X0XP/fKThhYjLcdNLRKdwo86fymHzfOinxkEFIPj16o/W
E5cRKFJr3cM0w2j2O5He4Lf27n4JvSz5icyFRyw49R+H0UQ7R2UbJpkJNAQV/pGq
Sd8BTtrLvt+zVxqk61glH3i7zDCmonUqpofZlQ+JpC1W80FjFnzBUMoo7+u/AMJ8
5y11zvSAE4Z/I87JcOFGeMoNybA/ZX2/VHXtdRrZEBSMYo+GuJ+YVYC7C0jj5k/7
HonHU3W/ZaeVDfm/F/wSBuqQSjYZpvc3DPAlNZPwh077RFyNEMQwtem9TQu4aCEn
FHY1rrhAYeAXcQ4BYGVurtOr5zG8lH8TejkUGG4IoDZ0zdZBLr3fuCV3Fo6FL/fD
EeJWBz8+QcB1NUqeXpnoVUS9b2UrwkMX87Rcc+KD5/EFEFF9rDDfr55R8i7xMlPW
LGKLfuoV9W60mcqy0xURwvvFnWn6WFX2vXPggwZU5jvlzCHdvgPXqT0UCHM5tcJM
Wvr56u06Z5tNV+aVOI01EC4wueggL+/EJyXZUuzOvcUka5AP06ohR52DtdsxQtpl
5+XeRWdVmvbOAgKiXvhujlOHvQunAGtUmzb+9S9R1Mk=
`protect END_PROTECTED
