`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBhH2BENS/j8HfBqCcaOl7Lm+5XZvih+/dfyS3jmGR80ttsEvb/J+Pm265X6eFvV
FitX8PW1CwIP2g+UjSxUfEtKlIV+AAljyW6KSXzF+XOG6hIk0ZvuD4Y76w1J8AhI
QjAkauKxPhgkpEooNzmjuQmJIxdaT87U3wpAvdkHMb2rAL3RFwgCbjr3KMSLhlr/
Zb14klu8Lj+QMHHX3SU3R181m9ZvTVeCrBdnvPEXATz7Z36RqYGdFCYbW+42cdRY
F/mOsU2r0uPxF4CK0O8XEynao5pSp4AhnMu4+HLbk/8=
`protect END_PROTECTED
