`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YkgNvNYfgq0HPB75MwIs65L8x0gInUnOiApNZVCK26SDmvZCJhDrt2Dw8IHlVOpu
OdLTW9yEjWwFoT+MHNCkoReYsOi3BzPkGcwURO4rGhjBHDWmkkIJpHy9pP8SR0jD
vcr/iPK4OSYNQSgFFQ5eheeV0uqpppd58Gn6CDBdkOCnYNSrIaUfL9aC6Jn8LaCV
1I5IuVhSADwnzTUEtqa1+wkSoP2qr1REKFAb+ObXsfsSyhc28rlRlgWbIuWRfzXN
BH405BiL3QwzxmZ4VFfb5Hv7+s8shPYlU+mQdc78YVX3wpvWIYcbwFlJjVoX4khH
Eya7KFwmEjUxr4g3H5nlb+vHyJTbHszs5xYVGMkAlbyH8ysb30GzRfuoXJ3tO29j
kr5bs0W/h3/hYl/G4EvjwarKvJdsffbtDQLPq8bDX/LNpdwJ1460Ipg1JTGJYVna
LeNmlsRdpQTIe8FOJDn8gLQ/FgSe67bWB0gems51a6bmPwywXx9mBTpOdRcVV0F7
9biN4pKbTceZzcYHi4+8jXygvFzVz6QEkurRx4NX9PAFOmvTfRnpNxVXXh4ZbfeY
gbJqfKSN+sl5KR1fmtjVJhXL8h1MvBuHhdvdf1rjF8LzT1RGxObH8aOoMM1paP80
7XApv48QdJxlvSfee/VdwHT+silXq5R05Ze2QhQzmvM=
`protect END_PROTECTED
