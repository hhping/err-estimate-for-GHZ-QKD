`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXvVifqd521i6OiAC7JAYLsOZCs1Y4RcE8o9sv8EKu7fbnsMzoqq4DsrJ5j0l3U+
JTFUKqbm23IX4Y8lWK92Yepz6JH+BaBF3q6vPiuZz08TJ3N2xbw33SFEwAyohrUn
+5Q2vIunPzvro8Q/SDLDs7SBBExyJbutv0j1Xr9c/Jy8wjT86lsdhjABfhABSaUn
ZwSMjeAJ3ncku7lJSQxoObHS9ygkfCDXTBGs6ZECs4U9ErMRVFgPJCjA2zQ0vIaG
xpIqzdiNIYLtqr/gs3wEmL9wtzY4BMkgfmmdKGmRu5kJ/YxRXCM51d5fMMJRBaQR
2LvQ6WEMlGIynFZ6YbQMf1P0orLmHTNCBxZrIEc4AcsITmV/F6uH7aYPt0YXSDpO
jJT9ysuD+kYDeuk3caW61U6zzi4j2amNqhCTZLcVoxJkxQYYLR4j5c+VBgXgGjuU
WviIA0hONxgcBj+w1gj3fisM8NTJSA88kbHDYslA8Ifppn4/socvH06PC/Bpjujh
niAn35qfN5w4VKx1U2k5whtErua6qibWVm1sa90VY45dlrQ8g7IPqinpBidCN4da
3MZQrsoi6R6Lxzv8QyNt5V42J8XgHg3aiNzgDHEUOA8wfN/mKqR1EKpKXFkAZE/r
JWliqOba9z1UkPRgkZaAhsIgZfKv5QJH5Oy6gUPwl1LI2ABCpNhuFSQrhWLJFWkR
+yvvoSjtpVR6zt48sy/mMnyvmjei+dClFjp/991Ay8is8B58cyMlNX7Yj71HGQvr
WdTJIFvwTEl4jqIvJfGis2FpYOcCOIciFYtfLqJ44esc48NP8zZHAU1FPmKprrLY
bCxJQ7jHs0XKBpV7ngC9s0RQjIDIZxEizPT9hsbNsU3TIS6ha+oAW2eFB1s+e/hu
hU7JriW2kD95qe5c3J3yEWHnwZqANpnGwVVVmvfq26xn1EXTJ2D/W1quMp4TW4pA
OGnKRliD2OSb+4SthKMVyZVLsmkEPHszdhTrwIOwCCXk+2Tu0dT5lWaBdPe2TKBV
UDRwbqPyc5XdXTGYsf8tEIFDzFshJSzIlbS6lB8vE+kFZvTdbysQOxRMAsCkrENF
sv4VDdkfNamKnzEdIapePIGR8dCDA4zq8uIJ5/ydIAilm+nz9JSECdfJ0w9ZCYUd
ipoOl/iOj2Cau+LUT1STGr92MzbnuJDTXQeQRc8Kr/bF8mq2o9znQ4Ped0Hr73LU
uSaKyXiqixSMUCSvzIz1gsKYElYoJ/j9Jdt87BieDcZPy+jlmxomxib+WWz4gGFU
mlfff/sl8uWcZPHpvRSO47vYJh/1uN0NM8R5PJAE3GAqK9/8aZfBOXpR+MGjTq+z
aixPHP39Ts6QmGR7tXIn/fFSTxjECighCrDYZZC+a2RAG0U7xAaN1aGytwfzpk03
YP/0Ut86T8MSSDYJR06ZJHyIgKSkHwLatG6F5aOgPE3Gy0IKR3JwGojlITs1E2aX
uqzJOhf3IEHuZoCbp51Y8cTSf7iv8hhylxGAH9KhJXauhAkzBnBzIApc82dnvY3c
SiXh/daduvsYwlXJd9BYITe+jb1Je82ChHlTHUeoshNlxJ+t6KQ6UO+FNYLH8KlR
1FwM8k/TQBhb1AHXm4vFwO0ZvIAMRu7MwmpWBrIqQWpw9Ynu04FYr9M3aFh0m0lD
pI/7PXWhtWz62a9+XRIGaVKGhbHTzXiHlL1+VlLvfr+sgA/tinO/eLqxVymGLLyp
PTu5l5yUZZqw7wv4ATEJCAXlat+ouQgBweyUKoRQBSaB60MzZSOfGzm+lfHfqx8I
JaMM3MvSudRN45RG38iiG15yk3aNZkhoyBSGBHV9akLq3KvASC1z/falSXmq9PNK
Grc9mhBZwmaZMJ9JDGlv6PHxqkaTGAG7M0Y0pFCdoX2xMg4BwUQkC3JZ3BNAszC0
Mc4HG764pQWazmAtmIV9JgGgr0X9EE9WAaOkbkvE9jMCtJ6RM279TIjhVw0Aqf2K
Zwt/6Fx+OzRmYmWB4aRCTBQzTMya3Jb6wXL8bp1Umvrjo8IdQSl3c3+DyUDCapwi
8xEADAF64pTYKjo/s6xLM0JP5Hc+xzu63OdhS06p4cl4mwUJM5aPjhlR04dWqwzN
WeYW+FzKDSmmbbvQIhdk1ya4SH4TxxpPVefz+rnw3PfxhR/cNXpLUZgKXK1rd2WD
IMLsYt4D48dByxLyX02FBdVVGzJHf/Fq08qvCL1HOBLp4QExxxml4+dCYYaD2WMa
+1mR3Wss1uO+Qyd1JuclbXAhJ5x6LmTtDilDuPCTOcmWoBJYQLOMog9OK/TuyAYa
1+qyQKTguFBQAyTpt9T69xWVOQ7U1RdfG9quH1jNY8onFaMb4HiMt0am780YM6n6
3JxQopZtHfEMeURsBRBQeRoxfASMEG1duOBi1YcjMuRsL3P+LynPSNx4lnb8Slz/
KpwQf/NKADob4Fi8PibGmT2I4cllh/4iSYFs4zcC2zIQ3uLtbvYVKlkYCQnFJO6p
Hk8Nu1a8I2/hT+qnYlay707k+/kvNVH0hUAO1O2CnwOwlPLqGJcu91gRvpGr+Ig4
7sgEs9cEBNhb2TcGb84LOT/+VN+4Zr3CIo4DWDY/2KevOLBqCB7SpKlIGInwrdy5
9QPqEt2Sl+fx9KQI1ATDW0XM73tIeW7d/CCxCM1ZlhdJ4YpsBCQXDn5506GtnRsS
RvkAf3hGj+iruX76UiNn2R4ZId1DdHI/pwiOk7vaVjmPB2g0gFam1i8gJ0gEK5we
RQccbXwg/ekMf0mqMc2zUkGUQ7ZNZlqKDFXkj3wblOKnOiykcxxWQU71YHu6d0Pm
u+sgbu1+gjEuQVdLMxCw4yBck3a1gpmKGlDTpnKhKwLLhlCMc3yjlqgeRG3uGGaK
Po3u2ckMbsYgHgZN90MXqlYJ/51gf1Qf3H4U8v16TTagBtw307f289NV8BI+InVZ
UtwYVHVsXvkES09FzkspO2FbYKXIFslfn9QHPY6tr2uTn4IfvGuOWZsCy71Tp9dr
tdarAD5eEKSuy7rdMhdJ1qHC4W3YNvTyLa6rlOlLP54dNHIIwttp1PUpJc4F6CuH
ZjyOvommwDtDyr0g4kP1T3ltvkxgC+f3C6B3l0Taln7T60NkYyvq7uDJO4LMqqn6
KBKWap7HJXv8zxNbMV1Rv5p/3VOuXeFBY7RSQ1Qx0jvVMnBTHUQO1ahpNXh9Jn5g
/SMGScJnLZS7YlCs8He52lBlqicmRYoTVcDaAzMU/LCgcWJfUhPWXZbtodpvOZ7r
uERa/CTzWoGBaXG6jYyktwj49fyc5g+k0ELCbqyHEAfMseMcIpFxG5v1TRor2pSL
j3DdKKNxKj0MOCBTWZn1W8fxrquEIronIxCnAqgKIgr5EoCYMDFA2cMoBFgQIxKn
TBYccunorx6fOUJ+y8d+Ek22937RsLjo4Rh0lJFhe5BDSDx6SeN1fbvynooSvD4a
cNh992x9jY4gUGP62y03Sl6qJ6uEh60dzeBYWvFN7Wq01JfPZMub6W9NgtSVPPMw
s/pFaOsJSu2pfa4V7zNMn00zov87dB1qyWPt/a8flyNXFvyOFWMy4eVRrREAdHDE
t6Z4vt0vNgNxZcXz1ScfhAEUHSRVW4zJEUsZkjvMzrl8k0Vu7kh3kOBYLsSdDFnk
5JUub1n/XDcJvRToLfpqwiF3riO5BMOdZoRH0G//jvLJpgMkw8M8lHzUBCMrR9Mg
jwC7KKPExyRp/eQSaC8Mo5BwkZ2xqfMq/8H9nH+5q67GF18w16wMYECAm/L1NuVV
cyF//7qIlegMqJmvDX7Te+HzyYrRW9MVV7KCeGdEgyXXWr2vCypRzwlxh9aMFqsE
dUIfLOKnP8kg/6EdFUHiZ9pVApnxImicEYxKVEOMRg0YySTQ6y+wqWvyLceDtuE+
weG5waWOGAFx9SDhryh2nQnWodJgHBHeL1hTtyUnJJWEoUdfd/fi7vgCBPf6kM7+
zW1qHLwUJRqrQKykHdKlhHkHB4cJDgxSeQleCxceU+ckB2LPWYPrYPj0H6cjr9Cb
/QUGYjKzVUKPm/CEMF2FyUn/1VSLlnCoADlo8UtWsC8cDGDREt6PTE+heen61rj1
hxUNNcWKZXoOFtnMtZhjd95vNVqwTvM2/g8EPnmdhscslT2VB1HDtqyueEGuPZnF
mc74mSZalTIZ3OCAlK6epLBGPeHLx3QIksucSZYbYv336Shg0d5377wOtRRWtg0w
sPTOugtuCPtlEPwceF8eOEjPT2hsHMyXCzeSe4/aaz2jDA6qt+Wnat79PeLfv6CF
NdPwC5ZQXh5MkL2ge/c/fezmyrwqj+5logCtzwbj4kQiHgNUjN3h/CXANSYTyLID
qQlqy7bQG3/gp0DX3H+be7EmZL4gmzLYL2riGQv6khcepoQ9gYCz3xX8jeGpFpXr
+T87Jo6xKh0Xv/SyuiPvcimiZK/eR4dvBckFoIM9QomgbqJ+hQtB5PDsbDZg/Uto
Go2BoTZPsTJtkQhp/JbcKtthbsWgq3jW0L46cMXQDX2cWlr1wx7zsVgdnV6W4hw2
diUqWaZ3znaY4Mbf1R31LbwaM0PF2zYtbeYZHjvP7vIpWTPyVsuy46VGHgFYlIan
JRXUOo3SDLuGVSQ34skk7xwDkNjr5AY7TyJdhjKlC5lTGNQmJYvNWsy1IdWGbs7a
e2FvbW+ov6sddzF34kaOGS5h1ORclULS1zTqz770brTtToyRSz1WnWpi3zc/ypnT
4VOC/Pd6gzE0KMeHO5/Vibl601MlIVBQ+C3LXkU8NuRHw9FaZ9gMYHfjftlgnljF
HoJ7GiIItXo5QLfMiFBbPi7luKpR8etTgo7FEcTXyNpuVpirsi1QbSqvpnXD28c/
8yZ9STi98mSG8Xcczuo8O6kj/ROY5w9KEstRUHStFjan4TtwKMg8qnxtfvZi4AGn
8tOhyZS/OcMZ5c4gRW1zeoGGXzSkyM3xigW67c0MmVRvkSxlKGFJUPvAGL7dlHn7
eVsWaK7NqF6tzDXgIMUxxIWb65cdz5yefRg74DZGNHbs8V1edlA0hwIjamPd7iCI
Qt4XSStxiBiJrG6+xm6RnU9m5w8wZxnq6xIv10vxOb9TlBybC95YxcXpYghPThOu
Hzc6+8B2yP0F2ZKuN8haMl8BfE8Pk6rSaKTdPZxOOz8God51IECvnBgZa1xYVYDi
ttgx4zBcxEyYbKOCCzZuCU928HJeng3Zpn1P6oFfnCeTLha8GSrzQqan23DVIgGC
wv/8tN6gCMgKq1jt+PIbidDhbW9j3OP4ly9xyWXgtPRiB6C704Af5f/9tdQ0TDe4
RTDVDCI7byFa/Ac8n/zfmEAsGACAwHRKRKPt+2YLTe/W3XHWrn6jXWb3ggkwsEcx
V9uxs+Qn8nDrR92iggjApIkdGvIP2iq6YtcY/+AKdUbSefoYL5m9B13CLvAExmBp
y65zk55sk3MGRduoaZxV+DjnOEqS8cdzoBUHyNzQRaPRSJZf4Oq7YWQEOnEh5hhH
879oPGg41bZcOGMfFTUoK+8wPPMD4plThYa3TCcJENIOuUQ69Yvekj+/1m9Nf3nE
fVDX5mpwX4w2U7P72IbzZFLUnutVHnytfLRQrAIu2wWP0iVS4faM54Y5wQdo8Z4k
5e03kOMPTY2javsK+d5BIcdstTdwNl/1owzGiBVfSbi+HHk2/MYCYK/QaCEdKITy
zKj4Q43ydQOOfOHQX2zwR8Y56ewXOsLpxOFAI5ILTsZXLlx1afGqdvHCXcYUj8L+
tW1aeJeokZx1jWhh9FlgVWhcyInSdqc8qqiRO5rg9hyDR9oJNt5y9XZz+orTCpTz
LYFGKpOld32FAaGOccm5Btllq01vReG9y87+/Tzfn6WFpUiWH4rELE7Lt96HRpxF
q1axjfxk1PNfugZ/SzZzuSRaHUu9upsOolMjxPTm8naQZ/9UY/aJjJ3U4Jy5Cnht
Fs7rGg/z7QKTov8C56Ldf4N+7Y2NnK43WE6SNiwgsbUV7gxPFHAGj4nBiOCAYOIx
DhYXobS7ZHuDKdJ8XBWFYUIIav6xZ5YF8HUQJwgbgvsMxd5oNZag7Sd8FQE3iE8f
Hh/AQh8a2t3Es+w844v6iCsQzGssmaxpFHx5in3zZl0+wArHPBYRCBOAAqYWJ3qW
Z9Dx3fO2btHHp4s2IGeIL7NXNydzQxbzTOMQ5JG7SFXyGWpBEt5f6TJ5vtRoXWXU
XqRSa5FLYkYos6cV7wyTnSdh8/mS61fm2LGyTUUUBuAlEIYDYet3a/iAwizEO9E1
HMijoqWlea7A+AzSJG3Hi4uWLSwCl7TJYoYt/BUOFRn7CbVpQ80LvHIYdr0lvsSj
BgVy1JGeAnWW8bNhuavVXd2gOcV5gS/UeKGNQsx1noiDbQc7Ou3Mw85Sw554TTTR
ACCdf46r8BZEEByNeVB+HKnuCcz45c7HxoTNplDp39dTkaiQOTBjboSAOlXk4wyr
XRfjUWoOeG1GwjvSaxHCrYXNtyz+1OCC/W/h+euvRf9zjzREDpEmfO9tMqM4/AzX
U0ikZrZLY4ejVYZjZpDXdus0n4uEZae0KsfiYI64UNeTF2YK2of27CaF9cwxpa+K
JK2n1gwc8UmFa3XWxezPahudVK4BreJMitzpDRxmMA3Dmuu5R5h2R+i8iDQhfZB6
JOYnVMQ1+0HmqpPAPTGP0bMQnLckORoFYoOmqkkBERCQgdGWTL62xqM0B4ey34rq
6sU6XPJpmpp10pgCT5FfQKjqKCc29XqhnRnT5ODbkbfJep+WZvYTMEbEUjrEuMPm
0w2J/EuVzEoj7llyXNpSzV5ygqjZCmgxkdHEcNf4Dj77K0TwiOyCGL9NakLtqJnb
mwSmkV+pgbZDp3RELcyh68gzP92LAxERufs6Qgo4FJAZgyucdL0tZVL9qMR4zGuv
brFTd3+ZtaPWsrc+GtXx+8vTtT9wC3QLZYOjCJdSyofPf0flK5Zv/ryoqunWBB9o
eq6r4yGKtOzSRB++8jNK2yhG5Tw3f8oNbm5P+JEy3JH1aWw5kBGW6JxuJlpPNvgr
Vbw6J4bbytxksbilQojZCtYVRpl8C08kyuz8OjHXoYJWOzpKJRjehe2GEbgn0okl
sFOAcDd3zmMnlx0srow5e0ElCPmExGNHrVYVdO7beUHps+p3XIDUfqdOrDYzaBx/
WcAVYDAgijoTVoRmDtDeaxCoPZWyEDqIbYjSpJYLeb6zdgyDr7M7j0dXFe4pd8bk
9s78vNHbAfcfO0YTenhhugjiGBits2xJTN1UyFWjNd0=
`protect END_PROTECTED
