`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHscjENPV1znLMcWwaSfZaNfr54ySYPjykWbjRB0VqqPy3XVdE2XOqOT7xbRB8UV
/0+Kalk1how/i6wHIoD6Ag+lFJLbmq1pKdlIwI8tPiHYFZu+itcbtxDhb0KN9xPZ
blu4nW7pzKMBC2d5I8rNS31XmVv7rIR9E1RMpmGW6MjrdjU9WAFqlm3ZiSSRlxEz
tz8rkgbbUn2Ds6VhM5sfCTuzWkko26XbWvQcLLq8Bp1H7VA+p0zmzuTpCMBhLVt5
NPi43Pv986Qcg3xoSdbKyVUZgfuqFuirLk3MhB3294077nJ3oBcd7dPrOu1yCT71
pZjx5xXHeTrxCz8n9x4EaUBIa/ARWYolBWUaT99llQ7ctClthsZrEcTCXUmm/+Y4
oUyGJ9pupr4xCjsnHJNhSjE9M9UkpX15TorkeQ6CS0Tl6lblQm0qdoNtsT4cDmLt
gOK10jNm0s/GN35235//COIExLOMwVL2T3d65uOrsYWUca2//x31fiY+/3+JiEQY
lUa7gcvmFynP/f/DRFhFGtAvEGstupNWw08sMJm/hC15GtBTN24dxXUHylW9RIxt
75pcaqxjktcofHC+TJ7iDPkqJjsx6YRrlNobBnYf10mEFbD6+5xe5DmzfUN9/mtc
aAX9soAiLgHVWpdL/kGjkPwfWDq8cagoj+LcEqVZCvpP5Wtn2Aut7j80rFAnLL2v
gS9XQADDVAYQjH2u+BsempFdrpV0g1f8FL6+7skQDz570LY5BTNc95ADKiuUaz0X
Y6tiHZOTK89UOtPzBm/QLT0bw9yMkVoYYyXkAPIFJvFbX/mdixSXb9u39B5I3uB9
ej6T9OIlSZOla6nkim3i2RBKWKLakG+dj6uXpnHXTsp2biNMA+TV3NPL1ESRWU90
QGMSx9JtTNF6kqTbgiCLM3iDeGpMXqcivrhllOgIp4Oyyf7g+WO3ajjNaTEmvoUz
B8JieTBSRV2JaF3Aj7kEyztxpNE+Tk9tr2PDKbTXkZWQvRsHgQD8fS42E4XIE8Tc
brPAUtJ96zonG8RCfPN+z6wZpsYjPBivd7InVPw0hBH3VZXg3ueb2ORwisr7COw7
/6BpHOtgtuREjxVvcyliVB0VYgigdbCDIcY3xzYeqBsWWGWji1AaZXi4Gzo7dgXq
h477Svfm0QQ32IZFDgCkzCIudAmCiFeGOdZBU7TBZXXXLNqVDP+1h+upaoOVR/MZ
7NGKsBRZyFt00pU715UBhWfG3J5EfZpwNQyC/dLMzth7BnO48zR1QUR8x9l2lqFh
0fMH21RcigbMKF9cGfkhBRX+qwrdXX1z218COR5s95hvBRWleMLhtX9I0Cgx6J9w
+SpsEUwvwO9vIUwSwDQZyPw82xnYj9SvYDw1zHxMj8rlM+n8wbn/flcCQTZvEYOJ
GVbxwIoPbNriVoDtuaYe131NSDv/QpxdY4PeBqBuNaH3IsnRm+O7WJfGXJXiq6sW
8gOXfpqD2N7UJzkwNO7oT/lytAIJL/rLqWJ706jtVLwagQHvAlSjGIljvBXcY/yj
hd7cKCLbOc89g70XDOrnLkWG59euzvOVOaudUFYjkFGdLPX3K/bgSQzoTrY29M8a
zMUc5S1PvsarzqE0o8K9W8e/TAj/D52ACtfJnjuzfWjgXYzgkwMJNl2arw0c3uUF
UDEGctswKsvmwOgzS0S52rIYs9tlVqxyPSMSe8TKmtLK//taQe7C2/J+uq9zQPYr
hLe1ozzEBkjO79cmIsd8sFm3kbc9JxrOcmeRYJBNV30sTqC9ij1qB4AZHqLXbixe
l17xIKi06cyY3RgLa9uNDBq3HoBcVte7AtiQkXwfVg9jxux8eeUPwj+kaD6R50MR
7udjNttsn7EkhpxJe0QrEPgCqk7Xt1SBeT7bI8He3F1E0i4/IVmbkfIqtVVI1vYq
Squsqvuet9NpEE1R8PDy4b8Bl7zcvic5HrJgl816gyNZPTo8Y/QmfXlIGo2S0478
1oI4hEAtZ56TMBhfAZvSPUK9i6BLOzW4bZNWp6CQfCysv4kWfq9Ec384c/zR3jkq
hfRU7rlayyVdQeWddG240dCNpERGW+dwWfDJcwKpKOXNsQ7Tswrf8P0gkzmKdLgP
7JmG6ti04rooz/dYJyxFYMf3kT10VMY019UbHDCV7FUIbzsL7vCMz7KKFUjqQzcS
s77pxBnbdJps5PycKRmhIEtoCb/tguuTh+ucGh8lbIsFUJ+187+YQiqtSut7pAcM
T8XLA3wRMiEi2i+Z5xBKt+LJxWGSysKK8jUMBawF2qkyKUrQpbTJ/4LWF39ipFAf
vA1xDsczZm+B1VM7CJ2SOxLIqEt7wJP9vX2+fE70WHwMMLNrNaCAtrPSKoaXHL6/
EuGBcoJhd41MKAPH8mq3BRkTOesEIJFq6TPNL8X/Ib3znc/l2e0ev3iUQ420HA8/
S68KQgzEmwmBCzq9/GlqxzLSEbgr5VexWYw+xHqEAkjre9azGmqcgB9aQqBXvTvp
WD9MOU10NiXoJCrasPDMXukiqojQ/n+waIXDvhlf3onKE9WNRaSLtlNjoFOHpGin
K2bA8TPgsuniKNdWfNoKiDoAOAkHUo32UlHfP5T0MxjAKUCb8tahSfIV71p8o83O
Y67Q1LEO/e4xVqbxlm9SyTL67/DNiOxEKmSfya0+t2k=
`protect END_PROTECTED
