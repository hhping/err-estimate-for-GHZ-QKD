`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOd+nmb6qeXeoadbC8YKvn6ZmMbOGaK+ChDnkpzpSa3dcxVW/eFnwFRqFUNLYmaJ
BTg4xdqKII+jh5fBtk0P17LcZ23USC+LeOw4YCwH/QCqsbIHjJLc5X3r5W4T2Lp8
KttpJKvsFqW2+rbarZbz1T1U3c4TmllP/uI+gJZYrqUF8ScoD+Ia8qVmKbvCj/p3
ll2PGDCjEfi2oXhgiGZv5e35uamzGPAe+vDRJQVXQL3bUA1swLdvOdZkuVCGY+5P
m1U+UWgyKYDonaoKHAshhuIuIZLKqNUT2Rs838l5gXksgh3XejUYFwPWI478o60U
oOPFEEH90a52ADd/FyykG1J/QP1itKs5mWxt8yLExVMZemCAyoYR2XJA79P+Ja1b
SNZfV9l6ZLVkGBFQJYpsnBv7j7dMNmMmL54DdrpW2/lRXvWdzvRDT5XMbJRInomd
2UuHY/MVwSf2QmkD0vTvMcz8/400q/PGBOFUbJpYwllfzj11//1+4miZExx83yO5
PMMZS64m3oAc0aGx1aCflt+65UCBvlGsNiEPBTjBdUemwk1doRXI8orzCa9mfk/b
EOBWtljXLc6UT83WMXkxOVBApHPZxEKafa3xznIwzfzuflvKHLXafiPjP3iKo7mi
P6aCDA7EclPY51RXVnfppsYbmrwYJ/fRQEZdUNAh9oDX/jstKHVBZImK44KSrOdy
pKJVyQ+Y+iluhDIxqwULPUBDGTSi75u4YDcMDiqrDZmrshSbeBEjuMhpGoaQcRy1
+wivoiFH4h07Q6umQAcEx+cCBdtOMfP/N4TpxrU1efIA0uUFfZI2/3shg5dPhahM
62bZqhbJ4wgvXGVsucuA4txzbXsZ7MsbL/EBkreR6V0Bwu+elmd0hDe0q8MEJFjk
4yOwEbQzmUp7LoTY+W0tfXKNr4cG5lgAT3C/FAD5zBTwXSlI1SqTclI4g9APClsq
WborRzOy7SG2JYOJoIdkiiST2mDkVd4JZPdHLlmxWi9G/AHhO1S0aJe5cMEHH2LF
AsG2I0PWp5GK+uakdu0PKJsdCo0dWz07aiDB0YSS1ChpkWVyJWAx9EhFaQlPH3z5
zqWA6pna0UeMeitYy1OxjxajD36jHsVb8jM+spMckcMKNCQvhwJjQJ89LFIXqVbN
R3r/r7ha/vHXVsh/4hroSvTlrM+r7lAGiA9aEfAgRetD+AYpk7ojVobtiJqL5n3w
SaATmU2pHo8cW/K03sx2jRAS+bzNlQe0MQVpoPL0Pax5YTEHG+LKbWhN/SkHXE3r
28kWnDuDZMQr12yVOc6QvzuabXxvrQd/hSVSXGwHQr2K57kGOECA+LSLI4d7XpMd
7wcLA0Obm+wru8q0fBlkpo5DuUy81IoHDj1lR2wshtVRBeLy/YQ4JAnbjiBrNrR2
PuLm2LeQF1+sHXHegkIXxTPQneduiRaNDfH6VHY58W/GeuyGwAEWlZ2sae6LH23l
F6cYEPZkAi2JBd2Sl4QQncwYCh0ICsEXkMAjLVvYSSwr8sHFWVgZVOL/3VDGJdvD
z6yUzu5m7jM2bdCc/GrnJvOmKD869LRihYxcT2y9pmsiUMFkZ/3zx0UR3KPiDaJE
HAoZrvm9wesXFguxtchIOFvyMuqTdXvYRVGNZZH659KEsNvVpDkGWNwESCFwfJvB
XCY1VLsQ4hfjhwXRqsVwm/0ECGAb8u9Xn5e9SrRlVWA3LM6CA32qmOaZpP9qxiKU
Y1SYYDgTVw5ZcpvvX7b3kkIxlKGq7uBDaxdZfcQcH9saHud6n+P03lkClfXw3rXW
vdmjqj85oPCymwbj80SMO6m4b+AUoMbREsNAMltmXym2bs08XwemJ4yXz3tYbKfP
5xgtefoBvnoHCUhEWOmszh+dorOUdrR7m2Am+h1+cjX5FDqiQ4DT4lXhG8OULt9w
VBzFMZo69MKUbqP0AI+nnoqq5GdIRGD6ZCmxbWMbIc6V21gYq8N72fFPiXLrExw/
z9iJQLId92ATxBdi/XDfBqccFhgr+ZWRB3UvTNllwC8UYrhl8cgopc6cIbq9QHMj
dtZ5+BRnpI3xwaoor5CnHGxiAUa5Pgp2RgNjGJZzSY0ZK1LOinZesbb7HMYtrYxt
LF7NgPsVc2vlD7x6wSub+fO25uVZspAlrnDg68+yGMN1+J+odEohSewPXjtg/4//
FJvQvClfbVWHp4+TxYI/vuQ3e6NQyZCsiGZIQ+accA5Dr4wEYdJsRNs446HFyGKn
SIXV5Yl6OqUELBgWMfn28yThzCcVHuoF0t6LqxcxsKYpD3NDCDmtgFRR7+4DH7GI
O1AK36DuE5J01Y0BnwM03zP+pmE0gE3MhV2occBrZuvQDo2uo/yrDOzytNjbJ3JU
7oTfTrGKqjkUHrtnf2TWvz2lsjstlF024whVbPprhqOWRTKHFl+E9WbFhZu8ObHJ
C9PwzyZ80zU2sS4ArQ60gEF+nMjn4a2ziPbgD3RDtu4V/2AwklDWsuLFmaQQlDG+
aUdft0DVcowLriWWiEzzO4tlomSDw894nkHy3ka7AbVH0ZKJeCbXISLBTFLLrhND
+JoYZJ7bV7bagHNqEXXkJZairl9bxejhraArU1FIli2jdHnnjfONcU7jeCtqwyhh
CNOv4LGIrHGEZklU2bFZ5OUzf0HFr1HJdHhZ++mkFCxZDwbqz8FmueSWUvd3QzrM
dDZyws/RIkErYSns2oywZ9xZ3JIRzomW9bwTaBaXdZzvcE1yfDoLx6X2ji4tkokB
jzcrynNhEp6pqHDHFupuICnMHcxTsRYRggPCTLV9wZGK6L9Dz+Bhaa16kd4lo19N
rmCtfjik4tOiYjo9UDf7kLc2ka8LpTG5bG29//EHjd0dGTkEu7Y9iwPmr+vX6fo1
37XUi3pMY9EJEUbfrEJg5mwa/ygfs7it81yC+jSp7iqwSeyvE6fn4q7U75TQCmob
b1jOX+bWIgRSUtAwkUkWb7KfUNmLq7UJ3y8oaK6qBM2GABZsWEHR1vjLUZvZL6YH
2pnxor46ayog/4P6Z88NMbMGKExEZ8QV3w+/sGyod2ofLrmJHCig6TBe8HfVVkg0
taU6d+e2t+zALm21UTAbbzGfCO+/FJbIvV1sIBLhfHUdnqcOOKb4tnL3NNOVBz9u
zwd9AGJknQN4LFRPjS27qTAH+uO6DFEamswf0/Fjs0Uduwv2p2FlgzO/SGnfIzaH
iMBsTYKAjJwQArCek/vnP453cPPevYQpa8XhDfQ8rHM=
`protect END_PROTECTED
