`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UufimInFihRpuc6yJ4BL7bu5BifbgQk45F+Hwazg4RUbbAVNefuXU62GyWbWqnUu
y/GSN9mBDoBHlVulptxi6KhBvYzL+S5GKRZyi1tmUaiOquQY4UFBL6Lj2e1QjgIh
Jqjwr5DHjScC9G1G0Nf/CYV4itICSjl4NwZTfer6jrqNfHD26dcSXmTdlVtPwN70
ag/HAE6TYnEGFz94ksWI+xMQ4d+WXb56Aqxwi5xrNxwaP6ZAl7tmV2AShcx55uIv
JHG9vEVxFd8BlqFmbV57l2XrUVlOC/3UuPjMFSgUZUHJBSc+3Dru1uNU7M+vDffA
FClA56dccJu4S8zqIBsX36Fud3yVQvP41Ls8Ht1nl3s3bGnpqAvAwgtcuHvpj0uR
OQkvSYOOgpLOnC0S9xm8EbvT+htgYTCfdsMYWG5K9OYj2qudHwioYWK6IyLiLCAK
0Sb3UtWh9ZB/6sbhVHTGlTsIZCyBWyp3u+We7XHVKtGXoQM7j3UsWYPxBNbuDYRp
DwPHo3mw0BzV+wkrRPyMovxV36C/sf+t+X3vPVQ1FhloVOz96A44N/ho5poQjm2x
I8Otxr9QSg4y9O97PaSxh3Tyy92BV2wCP1usmSvHdF9yDQ3b4lJNob/7En9b40XP
TXswNxIEeXpbqKp2b2jSqWHsv2FqSGuHeFwPYGFNb9NbKWhayD3Z8HX7h2nzyWjM
gAfXY3PY6jBr9oUvu2EXzxPws/YhrHPEhxjjdYUtidWI02+Bl5eO0ZJIX0fwQeIH
GGFAnSiAYc+4UBl6CBt4454wryZQuBWCWrWCykHokiXLy5A6LH/40id1ofOD6DIF
80XTbjEjpYJlmYDLEiX8mkvRqwGohN3MQsD3/ZrzSbVpLkGkFnWhTdHvZm6HKyBN
NupzEstHNjqZn8xy31808ONR0YYhaFVWIe4XoC0qmvr1NW7Go9DeMID0tRVYd5VA
CmlT8hCwH9jxbLPKquiR0gy4fijjkovvfyL3dQJiRhFs5RB5sstfl3/FOmldBuZb
IVR75lVNYbHefQWpzsUpAgDEDqQWo077oMrZCJ/q1WlL/GBrRgDv4/KGt9jZ+azx
G2qXMZx0H0fwgsv75u5VL+8xTAA71C2V/HOofvItdyXpSZHWSCMB6g4m9ppYe3gW
+RNPHjisE0xiLCgRdPaeIxS+PzbjbwSH4sMNubvn2nufu7D1efHBOBBFKftz+2ia
wfZUCe6mrAFU8hY9tLYf20Efq74Zab4XgJ+hW1yYsxqmFW5jqpI0J5je6B0UgczP
0h4arP10bIBnY/oSZdhSfnvaORmXuoyW5JpyRdPkEuSz3HvDS1wVLdK2qdXTjr3C
vqEbccrM8ojVGnklQdcaVIIOpp/Mbx4umcp1j+KceuB2qBfzarAZko9W1Yfzq2ZI
YWDDMeJIKmhmCx50AVWu6UeChwKEpzoTnQUx6h+gDu9535XKB4gmd+/zLfD5WmLW
RJjkaS9nUpZnGHnBMd2oXUI3DJn/GXWbI8Mqc7tlp8Gus5tXrDJ6lHIGrxh/rX6Y
7H+ut6HHcNTjLWabwLfxmjzE8VrrsqcW1g5e+XIC6c+8ihgFK1D5rQMwU68u702C
ZgkVtqW+j9DWhsA081Tgv6ApcFCUsrSqJVQDRVTtscsCpqn1wPYw0sP97JQEai/y
8v1LOizzL2w9K/ukgboGDSchN9tN1opQh/hb71DIZjCkoMzRcum1x9rTcJYX0Dxf
hB8vKWNjOjxCgmxlemGZJixHiTl7p3H1hAomH/b+2CxLxPYeKoEfnPcvS1eSmeKg
WqO0H3BLp+LO0LbZ3qMWvdrL48TIvZ40blMJSAYA+D47EuCAJNIAjyriSojwZYDJ
25qWT+D6+tHYg/jspXWMA6H2zuAZnd4zEb6GK07wTGfNOTdGgrHjuUKSlTgOXfja
UbasOpHuVDgAsAY7O3ym6rq0PjEJmaBWZCelQ0HuTAoRYxijn60t527uukoG4hbB
UhRkYXnawx0GMXqCH6uqu1Kf4r/Q1yOZgbDuBjoUKePoed8qRcrQVupympFNdpgZ
lPwLKczX3L+4/J30Ouxj95CjqLcf1BwFEnpWaP4fO/Gp05Trns9oyegu22fUnOQn
UzZWm6rXLiQ4ccgK7oKTfcQqq4x5X3G6MC9CyJ0RIGdlx20ACDWq4SsbcWb7GRgV
gRmnplCDZzrNnZ+mutju+gBUymg32SIBurY3nk7WgTgyLW33r38Yqo4/b7bBPbqp
Ya2FaSJZJF4+ogStR/cHZDLRHSU9/DBRzYIAqIoEHt996QbGA87iw+b1maW6CiJm
/be0Yw69rBeg9dj9Si3pXaaXa6om/KnRjQEOiHHefcDV4Q5S/xHnH+76gUwgjpM+
I2T3QVNYKeslUm/MH6yiygJm0ZZDvWcQHS8R+VQ+WyRAI2UK0oJt9FY47HmH22Pv
RjuzqMddoxOg/jzLrw5gHESzgFlCLn9sDoMAw0FicXi07rrZ/Y8TUMSROfc6jEo1
`protect END_PROTECTED
