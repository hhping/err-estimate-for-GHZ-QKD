`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/w37L52wYc1Xy7wC5+5oNU4KFzE26TrgKT66clPM/AjLlG8zRr/u7a+Fb5CgSmak
v8UqbcVA2sw7VSAi9dN0pFw3irKxF2hgypYgzXXit/1pYDL16YbGzGW6WI1mBV1c
h3NnO+RXtykARLTdS1fqbrNAbQ4RlUImC0gsGP4hErbGH1nM6Ys9XuaUMCZHMbWu
qIQPzLYS16W5JS86jElSMhGQ5LPD0yHKh9X1QtwQobofAl2yNZK7mV3Aj+lOkXIW
JaiprbrF+oyHZJwNwYjTzPgOk3xdVZ/dXt37zF0HjymPlDh3qyGvVKH6kqvwMn9v
5u86h07vuU0I8Jh1pvWpaNYWSIse9dZJ1+vjBlCju+744i9igPoIWW4z7GnReP2r
eDkXg3w/MooVdT1AqiwZyP/qE45XiSgMtf301OTTQa7z9nRgf2tiKOQLXJsEQkRA
q47yc1EfUHQzvWSTJC2CLv9A2CkCd+Fr+59BXbPqVhm7l785ytFEtpJ0xDG1UuHg
`protect END_PROTECTED
