`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTl9sPhymz59sPXXU4pSXiRvmDa7QAnzo/1oLvE6NYi/qq9iTTHg5ujXqtc/1kyT
V1m39hv36Jb1DqcAeuBBT2QKmPXZwWk5cycnoBMiPmEmkXG5YUtluC5EgjhP4uEI
AWR9j0I2TPDGRkUJZa+lnc/G4TwAWseYcJZbn1d2LnOImrkVWFH67f/wWrpm/njP
d86kR70hiR2LMtHqiHEAWGvZm5zCQRiCW6siGkUlLcOG2gilX6Ayj0KtIMfYGqUL
3sQTWnlyg7Lh6zmeDq2hSa2YeyvM0/5DBKaf+OmXAYbt6g3AHGBG4RSAuwGyC7Jy
/xiy2bwzJwIcMloO6s2rgVbjxyZeEfBgEGHbkLsnXdOapMGamFB3xnrl7lNqM5Vs
y1F5CDfldUuFsBdDoxC8JwNNGG9pBHsIIRCZQOiULUArkH/537727Z0XqCqpa2gj
Wgk0T6R8Ka7uxc1LlEZylWNsIR81I1D0PpZD8pJonMGU8R4nt3foMzfG4AJ6k8Oe
NAdj6SDgaeVXfsFSNra48Y/wTDNWq6Yp+CW9mI97MSgV3fz0K+tICO28KQLttIPN
7kT4Hx72mHaIyFlTHR0u32hlJ+I6asi6UylrmevDNRMrPdxkwECNHjUwXtMMsH3T
R/vOV0gwWMo672ay5E80IcocQdyFg7vyEZ5Ir8ret/Se5goHv9g0ZaEfPlqTfKBN
O5IpxD693oQFvbZ08m8xdbxNGy+xxXMro6bqtAd9LXN8AVLPHUV+dZeOElQTe8QA
TlDPyV+i8rxCUwWP3jr8WxECSk9zZVDI93Z6jnM2tWU11vWJiYYVPfdvhgayvQFe
Kbdnmz6m9JIve2vHhc7qlTkkHc5xh9agEPkAipNKD6f25BsgqFoSRdlSGSgOMZQZ
aGncwA8lQvAxI+pCa1WC6ltl3kqgHBCErKorMWBfIpzNJKErnwrFVsYvHbpGUcOo
iQnANdyUOeNFhPYGjv43LY56HuTha+fiJK+AGJgWRHas8q+asMJ3i3MZnqW44PPb
MJ2zCv9hjyF3j8TmiOmjCuA0Vo8B+O1sSROuAQdLSJ6h1u6nWhL0C0gCOEIAqnxs
GSGyLas062YgyNa/ApBn0Il6xBn3zgkbtU3e4jO5oPJVtaY0ZLBpxVO4in0gfKzu
3CpUDi0VgcJ/+JuM1KSBNwvnc921xiiSLYVSPqfEDVQ2MZHp2GyBzVDjFNVXJcge
m80DvS+7hXRIVbrpG+cj2jQ6KaaKDPFWzz9gw00kf2cdzxoCtJ0sBMgwZI3UhiQF
Km20mtFLI/pywDFhD0nBKTDWS5lMo6Hq0kDtyfoRkts4kd4412bH0UoC1nN5pvYf
i2VTnSqdqvZ0vhoS5it1lbP7T0vO6sllPZgfo0mB9RGOZ+SQ34OLE7koTXUy4dvO
918Ne4z5MGQ/ElZ3GB1C52Jt1M7q8B6P4UM1Gc1eG3I=
`protect END_PROTECTED
