`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0a33u6rXk8v9doHVt38dnaFGpuOHc5ghu4GiHT7CHN18mvSuXaI6n1EwUUh8aHcx
mehbJOPYLq2tjKVHN0tO14zzb+///DHpbUVAkPzV4RKDUM8kt7nhqMVcBWkb3Mof
kM8a6gZfeuNZOXRj6TMfmc1VKe/uQ+fa6dzvVSTPjmu49zrNJZhxLdJMH7jjMMbc
wCAs1W7K2HZT1s8jU/tc9My1NeTgxGWabzUx+WPpcgycLgxChCy6tgz7QeEwlvjX
7H1YvuY5tl2G6CDAygd1HbUYNZHyoni9/6PcI6/48EvpaUYG6N9uwby8/BoL+L5T
zAvYdAU90P2MebLaJTmesWUAGFZgrJQqYRCytqt+cyTnykBzc0GsXE/QjZH91+jB
m5y2wvbyLJFq9c3jpYxihVYZHY4LCU+1PvBdlYuEflZ4fJVtQE6kJv5MWUBHUAVC
qpmcLj7gm/8Mp1oTVdLpHumubC2HOjc78KG6PvySbnd6/olqHdfBI+vjFsOaySC8
Bn574lrigTRS4B6Bs+f2e7yTeNNaj9bU8McYIXM1zOULQk/Sb8D+UEY9RxRvC4aH
QtubNC4AhI+rRAsrHB7GbMv6aIaTYfjqPkTxfoZ3bECclkcPPSwMpqkl+BUdsN0E
L8Ye4KIlRrTt//krO28NBIv8R2VRsG9cdkzQjGEZRoX8qfc+6CTa+8U5ZKU+Eud2
p8u+mNBgfklUs7x0350lc9Np921Sy7lOlRq17dV0T9SiL/p0Tt1EcBSxo//sf+6K
VPIXw+QknHDGVjtEYKySFmKwshnl3SVTdgxATZ03OnK3QTuTL/RuLV+nfC5RTIiZ
uviUBCKt/Zk8M3iKJ0W8gks6ZQCuKteVRCgp57T1kv6ZG7NMYyMmv1R2Zne8/yOt
kCPcd3gWAjuOzQb0xyiL3lO7ciNCZN4uso5EyMyZzX1HQV05wcVnZOumN07NnCLX
KuCCy+mG1J1Dd/1eem+DMNx0JC6XIuvPHlsiRKcVgVY=
`protect END_PROTECTED
