`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoSOsykCK3mm4BeOCtq9byi64GV46I3775UFxZl6UP7n/qa1QkihCbjeD3Qo8oPs
ARlHV/e9TBjlx7g5Gjqb20VgDeMBAhEuGt2pOWK363jqqd4Qe68Nyp7VyFZAJKXJ
mhQEis/oHAsMLi/KAkUk70Y7GqGDVkN4uFCbel6tot5UcdxO7nu6cI0aGIB1uBBo
AaC2LK4KBiUPGrZJxvO9k6AlYgvuT5O15qT/fCr7mkcqzaIrGWqPmCUo3kN/bQHB
YaA4d5ggAjB8+qNYyP6l7SuD230t1hZdT9YKyPAWGNyh2ZZvlNyjYStuYbYUT6f6
QUel7SKChrhf2xIyIFADTuv5JkOmU8RqZiuO1COes0QQSVaNPn0j0QaNi3VQlVv2
qbMpiiwhAAZEvjEqrBOPx/ec0vessUZzdz8qEa3wFXEqjJHak0JV//+9r3bhKg2B
CnYYVHoML/vT4sipoBhjdfta3EGptHixHFVyh66D69Th2miHUPDLh+An2nFYiVSC
ouNztZ/jI1nDDHdnd+gJSzhb9emE6yvZeU7iBAzLJg0+3BSICpl+N4n1zDv5nF7m
jce/dkCgU3/XJg7XuST8R3+sORwxmxVw6ur6AUKdUpQkJXxVFM2eZagh77f3JQ2t
412MntMPA9l7wbvQmsl+Ko5fvuDKlwWcpdTpJ7l1lmVlbMlCi/37VsA1QmEXdMef
gmGRmWQ8RW1/CqT/j81ZcA08fmtpnKgO2XbNCC7CbwaCCJ5KbYvWfUXtbxEIYXhm
dwZwe+Zf5QvgYcXAaObBiba5pX7igNUP72sdbqCjw8J33rxarRtaf3pbSgzljrgJ
S86CPCfx0YsnT/Olyox9zgleF6r3oSMCnFZENGHOHvETH8xcLVQNAcFkKRtdmZeF
Er1y5OQIQaKkBb0XOQMFlHkTR2TZtfrjE1y5xQ3+lDKptwvkOFMkpcsXcilZlAK/
iBV9V4pnAJXLBbOxA/avsukN65NLDqbaaO9A6pnJCZB4ogh/F6L/8TioBLYqEAG6
8bKQzuR98WB+zZqjT8GXlfJMwGcCzO5sRNtKmjvOpCI=
`protect END_PROTECTED
