`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BIwlaT7ncU6f5ukLMDqjijbVOXSESMCHR64sz6CQCjsI+6iIPAgww+NhmYmBTQ5E
py+ApSmsndRpNk0BaLcL+dV6XWp3qisJJZDzzM6v/JdDRZMZy8RTCsVIJvQTAYri
pTE6lcIrkmefkAT7wZKtZaz12Pixkrrxsy8cGcU3GTjiFJ/ah2yw7pfWWPd45aGu
AWqxzYM8vGfmDUqh+lS/voweJN2JdVvKTb4HlS/ZyFfWTP/24oUGc7zjXcJs5YNj
WQbVPFlqwjykkMd80JWx8N76N0qkBAMnjt+4FEN0Tx5bzZWfWsuTnp2YVTRd10k/
dx5bE8tikG0xBQeOyyltC/u8ybkeIoWV6vMiZja0HCTleuMRTvkxzweXnpTaQZk/
jAe/4wxvbpJD4WJS2x2mIoyUgYpNViF023ufwy9RNa9C6pksB5wUPXB+Bo87Oauo
h5aazf53BA9FdlkrbONqsaI4KjN/JheqQXYkcHXFh+46ZXkrU8E6YgHy2D8EZ/Wl
kM4DFE7pNOCb11rs3LtvY5Ez8XGCWux8cdzxhNDB7EHOeQ1tcaZfgONNCDwITxXt
vGk49HIddcrJQa/36Z4ifbcbvwsNacsIdx81Q7vgM5+eW3+JyICmfuMxvNaETudB
73gozdpHWZfZ1YTiGGOmPBczJf0u7K3xCkHmpV+fAiUdoxPfMhHWUMDsuH6WwkHb
f6HllZKV06FtSMpnNLoS9a+ZYWhBPVCz9O3I/tddnZreWHWvxjJtjygbIlg4wKXP
071ZSHL+F+J6USbcUABIjYghnW5JLwz9SN4k/Y9zAS9Tl4SeCubxqaQRQ5ct73Qz
EU7RA1/kQdZ5aGjgpb7GoZKxdjCJdbcKIafFuCvgS5e1//dHgSQqz+0Jec9X0kKG
2An7597Dq5OfWihwaN3jQtp+LHh4sNBtxh/zb4TF/3eQ7BvmSlArPsyOEqSfv4BC
oweuNuGzxEaXDc9NMRQ60H1DazRRrEutwJQxj8zJJ4vp5gHC+3054AcIFzRMDA7O
CqKZ/xvN2yDRL6/WcOkDpL2uMcLLK6Vm/hFhARlBhk5BPKiH98nrsTWZIfozM2AG
iOiO/Mtv6MPQLc33sotp0a3klu7Lbb2WSVaOqDJBR1I9TMq+Y+IfnPcmAmeTTy3a
Drf4PykecMiHKy7tF9ccpnvhgtAwg5BZudoMdLbRfcojEDDtYtTmgtyJM/wb0eV+
KXww/1U9BZ0Ot54NthVtqKB4GK/8UgkaXWSerFgv70c6yD2QZnITvJv0e0tS3+hk
2bgo60M4LA2DTUD6WkfrGwef2mu+PC9vYtjLRMPZ6FlR+OCJtID/wFkexUX+8ByO
zd0VVFMjuYDOYiIH5ycKq+Fr4gRIURvuCEXtl0I2KBCEAD9Xo/wNs4vXlEq/T3I9
+A0n4f6XgOTObh+0qC1e7RuS5AnJW05gJX6ZvTbxQU76lo18JKcpDS2/KZIKXBTU
NfjLXZCacp2rBYIwKBPEu5k5o683tLwS94SGKhgK3kqwpMHNrKEVF7ygCI7lpJm5
gNZ8OwmLre6MDlvW07nlobbxIJjV3fcG2sgwkr+KKsMgrrm6JwRcRO19gQ9W4Sqt
6FgIg8DksADV32KhAG/ScfLV1kab6k+J8EYsiR4tV5AXlKR2nM0hYuszwLh8SoI8
/ktyE7O9B6CSUY8cjk4ly0KdpKGVwFuzorgBKfasUQyc3bH7JzdN+uozJU5/Mk5E
wjr06rNomwEX1w29ZY9ageuQqiCTj+sNwVafJ9FCaBLCn4wr27Rcl+1FhZbjTH3s
UXc05DZRthaoeZA5MsYJizVLzUIfFvduWGUuUq0uIrotMw42a5/M+tAyFpabO1yN
XUVvd6K0EF11JEZdIRF5MeZOtBnDNoIR0VeAmbmu+kScfTYsOTnhgpBDWmZC6oKO
czXh+djVJDbDGUsuWTBh981GkJEp0RxefB2xaMwHtb/3Cunt+hJcsx2ObOjbTEYG
kQy20/ct9+uBsVEyt181LyBNuEcYUe2SPNqK7BzVCUZzkrCcL18XgPD3D8CpCSKE
wxX/hoyv8p5jwsX/xiXjuV/61Eg1AYVKmFanGvU44oxe6fvDRC5r5hmmIU0Ey9MR
jlm4Xd3G8L5cb4ijGomFkvebx3UHcuvt8nnl5df4lFgikjkiQ/kEoL+shxO1GJ2Y
6cLZ8PxZbMJk4qAHC9IlRhFScqPcLW+5VMToGW6uFJhoSBnPc+2HOuk/Grs1YWTE
HeVMDU6n3pHskEdq4B4Mpz5Y5BPtDl+flnaRdwUoLc+9Lh1TQLCIfzubG8vCx5Dl
+0j7E98z5t1/WoZcQqhmQMIIR5pGwkLU9qyUGzzRMF8IoPqgur2HXu8Q1dWCoXUX
0TfTmafpFQnFrXw3qWCP0Qbcrejuu/qY1KKGQaeCQo4IRDhuArOGM8WadfLNDIBw
NXiTewJ/4JzACgxW6hrWtbQ/zhSgwpILFuVCCCzeFlFROUt+xiVJ7a9n4KWMJ+P4
iUyU8s4KR4WyWWB+BkcxYY3C9Fwh3u3jTUJ1+fDDriQKti7OGCQZVA77E+FnfcXY
ndH2M2sngBAKqFRfRtZBIqQK8ckQzbdxEDw9qSem1+Q5JwKkwzFkYUX2B445RjfD
7OfDrVWl1HcBlM886UalPuzdAWL6dhzW351ldJtkJrc2cgxXpMGqpPhmxp8wDrIP
9vIMWuifeV383pzBi76tUvhheVBgWmiHSaZk5GgxhSgpUAsfJ1teEP3bLLIBkV3d
/8RUiEE1a7uH6ocmDVWAyvsAsegzjDa7i/Smi+uaKTEKNx2vxZ6yQDLPo7q7qC9E
XV0Iz8Vn6fiFJEY3wOALBj5A64YaPdkBZh5Q4A4znw3fyloyPuEgSWwygh3cGOdi
8VxCU3bRuhd/25pCfCxZ7AbrurZtPc5WiVPnMUgKrF1piBqsL6Te6YpS1yvjXUQL
gqllOg1g0ZTZEgqsjSm8ESe5FrkcT9BVrLm4LJi99fpO6P0l0E2c/0R/Do5Wt6lT
+hnexMGQZmo0wZ/Xcl44uAk1sPpadOOqjq1vYg5jvGkBFa5eAALAJWupb3GWvpqF
6gnelfYSbcCXrYCLX8ey4xK/54ysWDLiN0+8cxLZw6dvlXsTl5x6ujGjSypBbwok
j7I6ZzB6oE63sD0bGwwsk3GuLt3DhzzP4xPpXGdcQN9VwZ20Z9xGCMpWcLcPWS6O
dlJodc+afyk7XB316a/yvVXQWDJ3rbVBbpj4ZiXV101aRICOAsN9IkAD02pNkL9x
Qlxd0lyZHhUA19Fjvivwsd4mUHiP9x5R2h785YalDEjqpOQN8UTLyjE95sXae4vI
C11d86KJGqgkYDcXlYRmGKArhWHTHtLwSLLA45LSNsmYabcNcxjXxH7EPwc8kTlU
SBoI++hjYHL5qQv+tnxbFwRyGue6B7VldYLmnxMywYqyVwnY+/m/tE721COoJfEO
qwxUC8JZb/W53cLIEa6WI9A91qlqECXLQuBeQtiuqChZ9/yLPNLKEa9kvSrZefjw
LNGQzqhsYHRrFfw7ve+FF6a4Fr338pg9PRPdmDFibl9EUM/+Xz/4egmJh9WOSHR9
YbknNib23MVEHsAVs9A3oHRgY0utgVLrF7XoV4iOcW6fAm7LXY/HpxHX3BvjOgn0
9uYGRzhC0XCnY665aSkrBJDRJGqSTc2WvbSFr2wIvGGE7H1JtYWc2YfmIG8xzkfE
2dM0uwk9+0G1SRk798ll2OtJiQu5JiYdApz8ZJolgpdI46eoTY2skBZlo+FqoKOb
HUlFj7e1yjbTPd/MqRhFqdU1ImRgCiDe+Hy6lbRaJABPaUoEgzx8DQZeLvQRAuV/
PGfG05Xhp2xe/xeej/WgLuVpGOiAPWhWTsH3QvndYv0H4tfX/5d09Nd0sogycVnQ
QM2mTqWjJk73h3IPY2EjvGLQ1gDoyQzudoxgUW6uE5QPThX7K8BkIe5+569SHUn6
qtbDUscNFKD897vgu6EGr6fOMg6xAary9b6dCwm53t9FoXWOooizIUDpPCQpN9xR
cMEVuMy1HewH2YXcCo1Z8xGT39j7jZ3sEw7yEYUbgEmJWi/7xIuLSFAgBqlXTqgH
SFIlB0dMHTtcFZdD27HTqvy5Jp7EQNkQOvgvo3LQ+vXylDBITIBWgyO8DDKBQSdZ
O5CSsu/3hd3wTgAyZySTuLTMqJj/bwK2VmkdXfApCKmR+4EQxFqdDJM0mSN9ZUob
YywSrzDYeYYe6HA14Al3cSY8U68G+Engbo50sZCAIPaA1ZO6WKAHibBj3GyQSZer
2Sm1yJRC8oXIcmgiJzKKAcfZIyePv6Py7+HFPV3LELknfEE1GJUEQ+Szzfq9low+
amvos5pkQrlEfs7/KYakb4L2516RbCPFvdsUwkmvo6MrUkQUjfaUrQD+RGLCDcTt
yfwH0ZL527UICx+37AgZC8lsJHMNv46adf6twHj/yYRmDNZ/nrKE4Yw05tp7paov
L64FN+NxngXBcHsgtCAJaiIo8jR6SRRGbLMLd61rC3QAgLWfbIoHJmlfIoWL49wW
BZ5CZ3+f9bk/FDeQ6SRWZR8rti44CXXaMb8U+HaoT9UotZF5X4wINpTiP0Ho5mje
pALEM3wo3wIiAyxosRCqnw+NUs4/3aOUignPOH6DKSPQDASm4pMDjNhC/WGbaof2
HMowpzvo1qh6zhBbiQy0t6TcJdquUbeKwdpV1EKh+ssdW4yFB8vvbL1RY54tujxK
1xGzaLmw7a9xEFW+YpVbHi3XGH4a9iMbURrbN5zhqEKE/yFIz+eBcOjDZjWyTGD/
AtcUyuNz3C8L01zSnHYFxDh2RAuSA7tPmzNKcZLBW1317Iw8FZ2FbMw88MzFbBXM
t3XZJ/xBALK2qNVAGIgezA==
`protect END_PROTECTED
