`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IkNeuDlbw5g5LzHJkfUvd1BXz7kAFikAD0fwIj4teb0cBYIHRmzI26TsQlDKbELH
82eVCZMer7RKWC+EDGcN/z+trwQ9IAOX3lFzhMZ9frBltj8b+h75N1ibWyWUzLrx
KbHGpvI1X2b3dyNFCYIoDPEclRLNAXJ9P55gBLslLw4Dr6/JCAqOEn7XPZhkjJ2M
6pgm7Ma18v32bkS+LSFab5o2XqndcD3MunuzSeL5ahi1ZvMXsRZgN5r/+gJSYg7+
9U4s4GjRHw77eTPv/swVAkZQm8qhhXILvI81RFAp6oo/s++Jp3XjrX4/0a/ly4dQ
z5u/Ywm9MEP3IsymuY5lr+RMXKYmQ4CoTqTG1FU+DAWFQm0N8IjCXgbHFH0O78PC
qxDtVMNLkL652v3vaKtYDf0ZohC1jbZwaQyiWWmfBKlR6mAcAFm6e3VsyDO1/SEl
NqyfZDMeBQoS2t6plMIADHrMzcuLEgnPm7caDNVet3hiedZhNDLulp0txYigwU76
LV6myhXicpfvWj4oJFkWsZojmEY6rqSxSX6M74ODZwGcoMnzwqsLLGm/r9Z2Sn6D
GdmJdwIalYUQB1M4np83vsXxdlVsDBsBtyIFNKEzNlJTo4pT70szGssZYkWTx+9Y
FFXg7hckJD84WKdh4ZO+wQmAPErmhqjC0jpW8XxulrhWQBIjpDhkz3LgvicyY5Ha
m/biZyuPPQUp2OzjJVNzIcHdc1OjE4jCqiei104hC/7vhoNNJuHYz6FHw5he1X8D
4hUvpVuWH9xm4pf1ce4rbR/qtdyY+sxEesZCpcem8FHCMBGpIo4EvCe+P625AQWV
NVkRnaHQiSl5kpylLsw4pJEkWyeMfdeA8pROb3iRAvMT9xPuGj2/Q0t/BKIYGnOB
4VzGO3EI97kHDELfG2MFDe6+GyjtyuXAszDIO8aQ9+u+jNzJY+KAN8tui9dcSDxY
N3A7X59xbvIDjniFHBEamdb51m/c5UrqaazmS4xPkB1+E5lpkCv3nlt9Ss/9Aqii
kQjSDtuF4W11jzLjBZk7KcM7h1V7jXA3huqe3DNUCZgmztNGk+pDywQAC832htQb
d6DWhEVzm0/mKul9xKtBT2k4GgqrIOMDjvBpL0YD+3WvSzHlLUy/dR/m7zYHb6mK
3FgmnWKuyhhYY14nfvXdsT9ZvLnCwzWNQCTXM7Liic+rz0zHDoP68U1+YLUBdrPl
V8YQcfRD/v18XOb4HxzHqoPr3GxIva6yrJn5XW13SnpOl5YETqBl1SOfd7+FRSRf
+bv6qGGWts0zbkNhdgLjWFdziI19Sjve6EvHBPIBV0yt2TEj0BckpnmR08sOSaYk
CZLUK+HM4rtaDhoXfq1O8/FVmT+Wia5pR8X4qcsraTKjglZyUDv8q0z3vwLUYaPG
ICfOnVtTeGAbwRKP3+EbzLxZIXtbht2iuWbaX7Mul40=
`protect END_PROTECTED
