`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wtqZsN9rd/Qg+bNimTGcBzULQiEBvy2hPpxhXUbGEjuaGltI7H1/UhQDvRZPmvQW
lHA795YPczIe3H60uLZcmTx+rxiriV/Yo2KYkNZK/cIBV73RDkhSTKjdIpB9VPnS
f5vWrXNDi8HP8i/tcHt3xEZfFZpji7rvbgmRyR+LZKUY7Jjc6gtNmWtf7V7hTyl0
buhgy9yk9CdEa/WP66t/PIef9Q3MnoxMAwJ6F2xGWA1KwPASwGRSgCnKOUX+mDK9
5EuJoW4LyAFfDH8j8kE0nOcpyRX9lDq7ieINT9//xrNdMR5joHKlMu2P9ZLWl0R9
+pybuhJkJl/z3JR0sMgxW7AB2T8en4G0x9moSvEla/qlAs9fIux3Np8Czvf2fRD6
fkjcN8A+f/XunDS84+KRGSPnnihhQKLKqGwKVh7Qd/klE0lZm9rdsrgxqycwt0GH
hueAtfI9cdf9mEmiE6WMNHFm+occBYZDfox3hrebDKVH0MMhe5/yzdO+szS9AMGu
3sfWg6kGRmP1N8W/utAndzzpZriaJIkqhss1d861B4rHqS/wEoL1Rc/109/xRMWY
d/YD+L2nchbg1OPylXKzvSz/zxMMG+AYCUja/CRTCZgx6P3ly0g/CvuNNEmR81W3
EIZOsVW7PYuJSQSG0xhWE2k7ls5Q/iuMyA11yLN+c75AHQtfN2rfux3bEXAtGi/D
WW/A29M5Dl+/98MVbitcj5Fzyu6jJUUtwz8GhSpHk0l7/zYuJMLyYBdJdaeLpo72
tFeX0AAyVS88exl6VDDN43Dw/GSnINb2jdzxVWRHG9OmZHB9Ke+sKArxussXB7OP
P1GjctI9uVfsG9hqzS/lTIGUD8f+kc5ycngRqqhW1cjl5b8qawe2q5NhKCc8UxJT
wkIepxiZrl1WWhEhBGOfMBI0SpIvoI0wd65hkEKZid3ZtQ69KPdDld08KYTfhIte
7fpg7ZgFx5ZCycALP/YSlJv+9DlHfjfKAIS9mF/Gpd+uMlW/HCl9ea9m4Viitihq
5+QkGVhPUL8DKGMG5a9THjTecDkv6dXmHKif70jQHlfOQ2xTt8QRpAEnBdDrW5ML
UJp2LhYdV0EmvlqqIo333/Y2KoL+PTfHLbI0mY/iCvTd/ARR6WyCqc4F6oPVEi5s
z2YzgLbhX82Ab7A2G67nY/cFNrmvHaPvne1b8hyXCKtVWQGDO61hKkHDHgubpX1u
42qBWITfl2QBAH9FUwMclA5uT/59BdI3rhL4tMK/nmXJw2xdl7Cpi4D7DCUP+6GI
C3xXIqjQyZ4qmVZtUIcWTF39C7Vm35RoHgnF6SwDwYXW/pZ5fUfaDGrT1wE0u2a2
rKz7tsj9fnrGoTHtvz5qFBKjZDio0kxZ2Dt6pxU0IJC+AtFQmnAO8k4WePk2YYqg
BTlJW3bMNxC5u+9PEQ6jthH1SdzIIPipFDVW2ysYYu79mBvBzvE/bdQU8/TqUYNe
QUVq/wTeEpijhksxFCoUJuJUE84UfikCC+uDeEwRJ3CjwKxsup/6Sb8z9S9o2/PU
0CMLv/a3UZF1NEBNXjGLGFfGM2WYMeyL6BZ+UCcydCVLK/7Mgd7R8Np+PipShwCA
e4CjNA1ZAbpQDsxcZ7doqD0VD8RDDBRT/pwasLuMIrKliZC55MO8oKR+beMc0KOP
tSWiFzn2TJQaYCnPafRbl7SAHx/AOZDhQ7vTTTBOhUMUUDzu+TNwbeUdTQ2rpQBu
ULnQQFJerO03KZT2vBNyxqnM4lqMP7qkSAo+EnriihIp1jo9q+aXj0rCau1JYPeT
Eb4qonRlQmzIGFLZwkdLBc01P5S0dhX+qwzMVS+Z5392ufaYzxi0BQkZjf6o/8a7
AMxzgnyw3+So6NetI4Beq3fpdeXq41IbAuAJpTZYlqqdUUmxSvvu1gQQirqHVg+u
YgQYS3tSRPX1PGvGBkP/luDVUw72BDbk7WmXH6670HRMuRFnjw4ntmYoeY3c83s2
zLcxCSacoJaFCVPrDXFHRTp6/uYriNfRWYaYpaY8yvEZcClWJRiLjjC710Q3WqYl
YXGhY5kZufLM4K61pYZYNiwMEApghg/0qVHkD0Ba6ZbteBaNdqihVPiZVW5vBp8f
4d8Er6XLqzl7J/1ofWRiTI+1pVOIIoo5/FsMMdz08mRzO0TWvfvBafnUTBZRWHQP
UqI/owmPtxAXcHCW9t4fi39LDfVByx4eIO1uIZWngJzvOUaJS2MflrTAYwMieg3j
YYPbmq2kvp6up7i2irBWt5iaOha1DJVvjWcUCyHcRsoJJncc1hlQuYr8TChn6x2E
bDQuxpoNns083H6lBq7nJXIA6lYR4pKpXYpH3JdIZEzLyuMi4H5Cx7ctvDWGaVvG
kP+5LpoAWJ0ue0+K6kqrB1MjGn0apNVkSdiN//gwcv498oZ/WuKzCqj4djPcty1n
MUuMwk9tt90UL9VeA7UCLXTbaKS8egbwDN6iy4HJnglJFT3/0Oga0ZJJCWOG6mEC
CSnhOyO2fgkevjAIjp5eL9H8a+KFbtkpBUnB4XaNf3JGTvP9TuOgQujjlDX7jVFA
7WgMp2e2uSREOHEZ7JzxRnl0h13PL0NcuXd9IXj7t1RHXsg7L8oJX0IDE8NjNdsd
Sn57l5rX7osbX05LV2vYQXj7QjP4+t2hMf3M2+6SN/zTzfAV30VfFDkG3MWvHeFr
/B5b/RaztJzLvrPxqC9M4aVvKaUFLECEIN3m4NIc+aQxd63++qi46jb+vU2Ha9RY
Jj4bUPRQjTHyI5KtB/Zro8PsnJBBki8DPruVIn8+7QDnT2PHOeQO86KPhoIhVhn/
CCCU9ZB5COONQTMhxWMfOYR+eU44cLuMLuYdGFDlIGOdpx6bZ/L0tUmgO4D6XVp1
U2HS2K3hpUW8Q3nDeBvFYDn3HLvIhQmrcEznyQRSxlCqlPYLIi6Cy18MWqhSjwzq
ZrK02LoLP7BcDbcUx/IkOSHRWL/4cEhLsFLc4EQZqjervRZl2ZSHVmdSvkrN7deH
IE8ZpSq0Td1eKiVQFPYGTVOoQ6fZOo4cmZ2el4W1XCgm//Fi3C8FaTFAGtC+3NkE
+Cdkl0amX2aMXyOBhgT3Rio0/B4QNlMAjwna6PLvea3PGhOy0oRElec05zaYh/0r
J78kco3lI+eGmU2SdWOoFejdtDzRYJ8kxh7lDWIfZqDT+4rsBR0ZaFZo/8+hKXzK
g8SHLq1ADDpAqk372fEERvhqTASzMLsfv+A8jZzKeCvMI+gRZSlz7WFJ/27CwBIR
PBMHUMFegahDOOibI/AZMOBnIavoeuoAoYOUnK1r4GPAOZ3ryj6VHv6WcjgLQfyN
JpbgS12IoKpl9w1Sayv4XHdHzYymR3YHfUwZ7CCQhBqRsuPX/o4BBkMrxM25bnFN
aQHxJ0JzTjSSjzpqT8XfoOFxbFlCEDfeTeBERpjqhCPtRaknOdJ2NkNdxHfRRXJN
VcV6bm9jASOLmNattorprN5JYAr9p/QqlEoHq4LcW1dE5soiNXVCe7G+IISvctiq
TUISX8iXcyvdF5Ybt99VoH+aih0iKeLmXA0OFrHAl4rubE4acXKHksMnz0T9c8eU
TqL90JDM7H4GzzXH9VEfLJkN9J7g5YYpzsSfrjlR5ljtf5uQNeiH1a7g1D0bLesI
Qs5d9+n3drqE3TNiOg5ouKcG2Mcb+s6cvhstce5+pY0+/WzeI9u1oYCo8YLvCoHr
yr+QH6CHTD6FgEQeRIKt1x0uTJdpJwm35Wp6VUAEQ2ulWGoBGdY8hb1l2UTDvQqm
oWxej/VQINwaEgK6/lHBhhez5HMdp5dTA5+46lAS79uhsQsm//hZnL7VNjm76C5A
FSiGX7rQ0WPywN3tcj2Ly+IRJKLJtR/hD4IXH4VVuDk2q13pUVgBB8aUuxBVtXpG
n8vlSdRTwftX8pjRf2rLBXeyyEOopATcH9h+yPpr4GknW/E/lexdZm/wmCHeo8bI
ZAKVMyVXOePyCDz2KFA16Oq1EX2416gLlreRttmt42bxIN+N2eqX32KxbaGtbmhm
KGOm7mkA+APY3hrg0SS/GmuMsVatFeqGafEi8zsY/RsGyrBELXdwP8/gV5JkV+1E
qsgCiY5oEnQUjKbURZrVKP9R024cKXtGleJw2cXQuomqmqO0SyIP+uHDuF1Gl2kE
dyuEMslVfGW52MOj9SwYRhdCLjTUTbHxQZw6MgIxJmt+mPg0Fkxcx/j2M8W/vY7/
nbY9S7TAYlmCa7jnLygb4V4g3TMA/vb+Ck/DIEm6fEfWDXa4E0ydINj5YGHALKXk
5cS8tInlSyBaBB+ZZb+gnV0m1qE4GIygS1zYEAfOwmHGrX+FHvSvM9PSQcfVK2Rs
DbtnMemtb8QwIUnd/I+UTIh7VBSk+YuG5xQ5aRC/wR/ZIT093wl5unRkcfnaxHLu
7EZZBBQZ/vrLDS721zgi6OjgRj56BeM9fu5XwmbZ9RFmrC1I3FIZmOWQpBIhb+MQ
oMufv5j/bdVkbesrXDxRjGmBk/X+acyP2uSBTRoPNIJ3ORSINMHr4w1nUa/cyFuS
e09VGuQqyVgolaJibqW+6vxy9NqCdWkkSSMfLdg3AY6KeQwKne8eSH7vA9XmXicz
VsggN50svCs9Jpsw+/cxY0RgZ738exrlE0L4bwE9Z8ziAF6ZYOi10ez922ZkKcNE
Z97ogZjvyrMfIEBQfwDUyFGt4qBf8vx0oqbpm8rZXSX26hpHDC52zxA/mNgTKX0e
xBopD6/f1v2nnXX2OO1UIE2wtwNXEiZXZmaIv3pd/vGgL7D1hio0jAubC6V7QqXo
97KQLdkYwVxYDM8St+6xqUE73Ofp386eKYnv6/nDQW9pbJHRoFKcH5tMcIzehkXE
3RxrkYfHL3akF7MaTPaiaDU97oR4IwfIyv32D7OQBpR6VnyrNmAkku6Kbv1ZTNf9
o+XRn41tN07oMiII7YePpAEHmjDaPDeYl7uTZNvMhNduzaQ2bAFvW4tiNse7hLBx
7yPslAR5p0JNzgTxIqdLEBD9sIEKoe/RNAlyM1zLWkwMP31twr5FukHqHIdoMuBZ
xBhpifCwE5+fO2ME2Ws6cvbDLc8ypsf5t3BoQuqqCprxr8M0OmEXHjUskU2zQ1Xw
i2m5NXvDpdXYY00oPDIdaA==
`protect END_PROTECTED
