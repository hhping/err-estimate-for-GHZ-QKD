`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHwEwFGJF1eG8WA0pSsBY8WnR4OIXmPrZBf+T3I6SvlMJMtFHypMD/9+iKVbkvRy
9iypYsU/hqzzQy9beYZ9J3hE9hBj9DV530w/fRZwlLNC44UmXrnpeq5Tg+lrgQ1J
yfJtVlkoQNoILf/MKhKvPyXHHocqIJamPVjriCicE2Yl2yQvZi0RvkWtsLkPsPfI
x+0c/QfXiw/ztBdFFBq1IEX2iRof37OOvZWn3MkRcDMqqt75PWvBXE3HDpCZ42DN
sY1rdarUxuiHrHAzs9MUkaxFOd0qmCIO/xY7mRWbJw/9CJkRSeQLXPe+ddJ4u15P
pm/XBy15SsR9HErd3fAq69Dt7ecBz6p2xWxzhQCV9XL4H9UD0RVX/k26VxzoaH0y
OLalxRdlhwzCF/ay88Nc8riqtytm2AMqDzkRy6/ayL/CB1sDNod7Vx4zrmNfSP1F
6DlfGTDj5TPGALS4vPfRIUVNaVtS93mZEqG7Yfb/C7Dvl+kd1pvdSznSn55jQzSF
u+D5FcLtZ6RBRP2YtyhM7vhWi2WiKmKE4wNCLltcCpJmHaok+9GVCOwnyCRIBDds
X3s3mSG2o5XW/1fSK9u3QoV7tgjWP+ed8di7SUyceasbxo7fjNgw/vY6pQkQrksd
Hgavds9y75IhYbqOXhNKUNjnmpeuraHSAf4cQhCwfK8/l/vDeHN+fUESMswA2vY+
Vcx4aGAQcyQ8/WWDKRGACLcJ3JE2ivdGh2UKyzCScko/dFQ0ZwUYzJTzURL7e8gT
Gfuh3ptbV0cTo6UJftgHKvRW2vV8/G3kxzreX9k8xGeIGy9WIxYvi3Emh0XcvrT3
d4ZYo/uUOxmUaZwtqrtHfOKdhuKjso/rtbQWm+FQGeBeqiNTOBnUJXQgAeya4xxg
OisOL2zEFEHSauF6YiiCzhflBGl9xTdpyb9aK56BAutwctqJEJsHmRmYonJ3jZV+
ZyTAx82Qtg1TdAYeaTGsp67nO/JdkAYcr8c4JSShu1a51Hr7Q6dq+KZewE7XISYo
qbLaV7Ss/OxBz2oze1NfVas4CKmsICE5WFOrFYImAAYKEfgqKtTjmVRIpSse7soQ
5QG+MyLZJcOD+WZNIMhTzRrGJqKwWOl3qsYtwckDJ5Z3Rir7lckQWxfsGtDhPj75
OlRKKUL93V6IjctcRcf9CVq1J20pyJf4/8pHmNbL9fQIruqhcaf2zrcl6KigzCsF
lzngxWB62ZXOkg54Zn638UMsbOUdf/LOsoUPAJLkJyECWpJbWJ5e5lSXL7JByIAr
ODugie9DWTY3I2j30soGbB9roXXS9x+z/VRW18N1Z0oYE3Q7gtoFt7uD2C5XAD+B
h9LiIicvzLnctrhiCzt5UrZtf5YAAqr7l9jShdOcOrU=
`protect END_PROTECTED
