`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IR1J/ahdA5pWQOIWgEPnPccdXbyqXfMv0fCuU0rOuQTvDiiSbmtJprsbXocHTK1p
djkYPYloIl2RI7KBtr3ogXIGGVniifWHTOaFISU26DTXE0AnqLqdpddaQ8jEo+CQ
p5YzGxY0vAHIUNKfnkJ0E7vBYU6cnr1eJfj21JdKYfP2rMrC7/s+keWmWXLXO+Ae
XbVXGY6TdvzyACOtDUXi+CCLICCHjWU2atg1YMrWcxIn6yUXhxpPjM1wE8xOKfFA
ydvyU6z7zccUZHW12OALM9ejvIGApXQgroPNgx/TpIZUgfLhz94tbmM+okjvge07
Y1fJOcxq3wJdBzsAAj2cwQ==
`protect END_PROTECTED
