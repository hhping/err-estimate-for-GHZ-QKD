`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBEACi817DVDLippbMcJ7jinuDFs5COavKe0okfoKr78iCceIYSwAIJUCn0mKG7G
w4DHfZlsq98optcdKdz6cZvkEGWmdKZZfpDBe18S6XdZWv+q5xxwtWTFvm6DVZWH
bOGjL0afvkWDGS/0Ax74FAAvLJtnRalv7tFL2A/QRZqKjXMEHW+d9Gb91/qbWJec
WZGhu3A5zs1teewSNdiafQsRJgDo0m0oWvL39Fd1Ziu26WkUCDwA+uv4kxSms5NP
8KxVUkCQSIxLx1yfvBUG63cNLLteiz/gP7boisJttaiulu1BAn5zTipFJMCuDYaP
UJP3RwX1dW4z/Xj+ANrO8ZqmeG8jq6kQD9gftiRvJQKvSw/EIo/w4u3+1OT236zR
GANK46Z1++hMhFw54CcU0o3UOJAh/dDlLw051aFvxr9jL6U+W5y8KXRe74Ms3dP+
4lfz6vZR7LqARzxoIDADt7a2WIFrA15i+FwkTCc1oPhZI8jnadvIPQ2kdMm05AHx
3Dch9c/ZC1F2968e76VzaPK1oHkwZXEAw0gXsQHM9JWqTOdAZgcA4CPe3iK4tlDY
an/7HpdGmSF352f0dAxc+r7U3jCzQPzJST91CJUG89DMbaWf3ikQm1YbGThJLUHm
EUbnYvTe3eTIA+sGZTXFXAWiSjThxAzXH2vEuD2h5b0eyUk6upV1gF/yiCldluea
bUVWeiniGeA1ptmDQPT842g4w+pCGkbHlhWTawGAMM/JMUjEPwgyoUUIA3oshXyX
/SYen8GQSoJV6O8ldY+C6exv3wofao2a6Fl41xgUnSGMHLm6EfzDVxf2FUTyRh7A
iw7jnignLujl92Wnq5b/lr6twoWcJEjXU83Em2Q24RC+YTtowDdo9M4N2qk5Zwj6
GGQsDv4fcVrehZgwfD4FrC0Ne9X/zXMbZGJZE3Tn2BaiNw0ToOlnpfWiokxfzq7F
XVDlFC7AI2KSzQuCz+I+KwcbEY56BEShAxsj8PKAYnAAMH3HREQ1HvqdEaJHUZur
M3mlSeTw8/oUFvROnabJqBHLOAXBMYruXZRkdyZh/Aa+G8G9O1M7jByRN5RCcFNS
VIBHS9kGv9GcdltjLhpuUiJr4zrNdoYNnLWNgbG4LQMTNhoY4ZuMzm3CagSx0To+
G+7bPcQx2RxJis21GgShUxbo+hKaaotAV+DtakAfL/kzL8IS8sNfkPfaNVNB8Ta5
942ySxuazksfzGFE9Won4COW+QSZev+tgLC6U14vQfBXzH0tdw7GHLxh9lWrRE9z
sFoOVfPw13ihhIQynKe7X+cKNMML1NajtYDLLUkIBg4pQxsxK2ggULHB7BTdr7yZ
HKq7CL6YnpVtnO96FXb083xJQDpl9AWz5lhuCdEcsLOjmEAfqjwcpJB5+fE61lM9
/9wNqCSOdNGSxGEbIGlUbhoRwK1niV9d82iK8J3ByVUEdjk1WeAvbQFDQ5K075f/
7++JZvvSHyhbgGboodi+0f0+EZH6FEdHi9OkVlxOAgs5ApcoIK79ArVpVpGo63Fa
D8ObyQ0iNThkJDwEgqyTWiPPidIIJgm3JPx75SENe9TPPIf3wNEzd3kkNvu0ahT3
kYsJ4HgZ7m3qe3kST/Az1q/buZ0CG/pKa+nnJ8+1HobsH/sDmK5D7fTL6SgnlHFw
7bzw8jGh8Iw3ZVHRZp5NWBCf4ShnD/EndzO59ELj+uBcRZuInf843mTbD7DkDtoB
mvQUv4uD1//rB9XkciZjrI8rFZmfwecG2apukhUj4ReJB0AqdHUlTRmQt4Mx4uqg
QJMwCOcP0kaGcwhwtok9MErnUZR0Zkl9/WRbFSfW0SuHigDbO97BVQ5LVkvb5z4K
KwxJtn5C9Os67REKSav+2gUmjnMMsbO4ki6yD17t/BXIdHFHjr5gfybX5RFY/DDv
De91LXYueDyn6v22BdIOgOmoLE7H72F9YjDajcH7LbM9kETqkBFESpAE8kSXtWOd
HYj5/hpjDYWLIFWd7Vx1+y9tnIlWQJDGGON+gSLOPMHconBZGusA2LJ/uR4DR05Q
e34j8oGYQ4fkTgKykOkxdV7Yx2M5uvp8NnNfpdXK9nJUe6J/cN8YhHcUUg7qDUN2
SdJFvYnv5jolN5xmvySDAf8WZiiIilBv0m7O1TqyXQMQtxpVM4mD2uCZv2erkpZO
VCWNn2NZTJL9Rx65gFm0VixenPN/SIBiDPLfhFiaoEVSOcVNoDbr4915/CAvkxly
QbyGDpScViooAqpznWxLy4l/05MDxitwWUj9miQw2JNgi31EJQdyVEj4nkshP/z8
+e1h05BE7w9nwdHXYEz+/9qrTRTgdifOMsOcSXtKZADkNLwjMEZVpFasxnDxbgKm
YGAyQPXh5ZzKzqz+ukK7NnGHtWSfToYk7USr3v06yELesGHYMNfyCu45A3p9fUuO
JC9toeS/bsTdCra4ZIYQD5itN3PpNEk33lBhxB6WTVhYWgGC3SGTJnXPQnetLv8e
SkZNopDb0UlGG0yVqnVPTvaaifvLo3lDeCZGHCW2+FYLBbx+UspFc2yDL6sm69Zj
Ev4rTeS7dpCRx3v12yUgLEmFf44TUzh6Lcrft88rNSuxwwTubEkMmvigzV6KJkpT
ZtYgXBvOjoFRDDrYToPyi1ioX4dzyKVAEM5vAtjxxqnuzeq4H839CeLzEqL344YT
E67H7bDcZSovuUErh4HuSl2n6B5g7vHIqPTSqyZWj7Ii+sFZ8RE5EGnZmJ7iL/jc
k9vV3U2UgQbxhknxrW/qtYrwrQy3LjE5P4NyPPVLISBHMEuznTHPRdl+IUglFwnR
BgUPAcR5mAU/GpQSPP/utVOZjVM9v6sgbVtRQ8bs8A37vEYpjvbqYyYYkysz+K7e
f1rXbwVxnc+c9tcr5AaoJQ1dSY2oLGIw6al80C7ROX0Vd8OCHlI45OtreVaVeK1g
C6TJdbjQDM4gzSdq5uUP9KQ4oAmJkQQucCAZgv4Rk+ExbeD3U4+2OdZWh1WPWnNb
Zyb0LlWO8onjKNwP1ovs4Nv5hBtBlGf7cm9AIHZgsIDc8+MZytyiRUvY0dxZHeIJ
5p5282NFETr6sYswB3k+efC5DD61ukCEA02YZbUC2OeOnFkPQpK1eptnewyrCiXT
9IQmRxDXb256yDiUW0kd3IsXgQl5yLc8CVddobdjiY85ykNqK0nsH920Osw80TUn
C3cfsqSszad+HkAT1b0S1RE0QnPLq9VtWcwD6Y1Y0A8PFQt1NjvZuXxEbvuR7DuW
fvKKSxagbWno25RzJPN0t1dpDTeGvK2mMuw0lXOYPt/8sWQHbFZRKdQZzPbX9z0u
J7yYHGFqCGKId9jHhx+XqeRPhFFXqG6CTxCALUKYaiMatm6SVv5Xkjp2gMv8cznm
RFcsnRQysbftMNujWbXVPy9gyWLpXBIhF5sqQodyhISvJUWLa7YabBGI938SLeGY
YBrTtdMQg9t+Bqlv7Hmcvd82Tw3+7nLvvlY1c0SfvnbXBEicFLoVD/e5eKGpKQU/
trQzUM8HOSXI6cup9nGCz/VBkV8sYSdIBfIN1SLEXpy3K4VyIexUlblyfZspFXEA
grn6a2zTXFQYOfmNlvuru+XVN1EbeLLOxsnNm/my0Jg4rSOBb31/fKA72jKF3zHK
stYMzPL0BwCEEXNGgcB4Lu1uOl+LVl+e0UENvY3m1xgFstWSqiSBXI6oTJ1q6+Ar
eH1SOVpFgSQ6GigURSEfsuCz5ytk0qXPULq66ZqziXyQ68Mwv5x54PqGXqSOIwvs
uIf0fq6uHzPyeQliNWMPa95WLATF05tMsXq2G523zXgmjbspG9RtwgfkjzA67BqU
GiPA5Ii221Y4NrhVvAeDlDL1RsBhrMBxqnBXe2qCdAE03C5U59PdqdmEYLv3o1eS
AxvAajchEjfi4hmk9d+QYCVS+o+qcpYmVjEtnRPVDpNv2tM2LZnTYxNCwHsr6FS/
YaODJ2yKqrAdwJ3EveUWy7MqVpv0PVy0DQ/e+MH32pdnSCFYY8nH6dcsRVcgJPBK
S5uTrwNhowK1iyTdQDj86wIzR2shYmT9aJSTaLWeukSFGJtjNTBOa5/nDwY2LPgD
ZkGkoRm8KiLi603K61ULg0K0jnPaJ9zsXnQoJYFSg7+rOz/293OerrqdL2swV6VT
1CmGKbNiIMizxzfFg8H121y6zF2lTzvw0//HV5IXQFjKSx5WsjPt3nKXDg9MmzD3
xGsRm+apunVQGft5CB/lzInoYi/lzMqAP9r7y33mhlIFvkI+1CsdEFt12J7ckSc6
vMBtpR3rMcCggIYNFrYdh+8H3iyIYyRYTpUzAtm2Vbw4MpGqRgmUvHdy1vuLjdQS
R0bhKc0Qf3C35IcyAbG9Pr5MxhbnUn6iDp348MYlSW/6F9wexIwIcmxOvFGzisvC
LRhVyNvLe2tgZaSx1WmiGAjFy/L9Rk3buFR6+5OVai92+mH6FnbMN+SmFZGtIpih
i0BxW+aNexRqvr5v/yBqP4bFAy35DJPsQhPd1lV1sZAmyHiwSLC8CY9VBhl67x8/
KIl8G05OCDO5zPwndVsqRMONXxw0e1zcyvtzZANnDovzgRl7bCPIBk3ki55yFff2
deyGjCC35j/N92LZbGnnV3WYWQCzf5bDbIUcJ9fHcPd8ZWTTqPKbTXvh9o9hdggI
WaNwITV/QY5F9OFyd1qLIDD2gkEHXXVu9dM7+4sbqjGash1/ai4Lfeo3PupeCovv
K4ns+UzwMsbsBvYkuHkmk6OcD6kcWYfTXQ5aPSj8zYc+sJdb0IHVZAk2gmjYUMe2
GoVjE7tc4xdupuXP6gzjOKufDP4CskpE1NfuQGxMXd14+GCVDrfdAlpuU2p+EFJt
DZ5M06Z8sWTNKG4Ab41YccDSVNyJOw1gTQ/d6UHA+Ca0nr/MolfW9hN4uGiH65Ob
Xmk5Wmq9B+9dwj9HrMWfvu+0/v0jQJs6O/TpY/M1gh7VhKL79mvaiIT+NN4dZRHf
lbjCKnI/29IyCoz2+sqPK7OoVL9Ocdlj/tWfGFriMJ5a+OmtOtLh7UsFdr4X7YlT
rGSJpvE+Vg71RzY6WqTLX+erB4SGRjASgzQd3CFRVsPdKvUIPXI+kGCwhRGJWZAe
9JGssl9NFblOstf4XxdgKXF9OlUyD+gyF2L+rLPk7uTvsLElhCGCfVpLsPbGviZv
xMhZL8WWAOU11QKXZk8uCTj/e2NcI+kl1IrKtrqiKPBUKI62WdgkyyBoWJt2n7Uo
Hoj1aaFL6gNtsg1dTsB3gKkI6l55tzqk9nwkjlBeJ38Ukh1BjpnMzC5T7pvXwvKd
ywsrHAOSuUWPjRX+yB99QvjhNlRKYhet26V8uhNSL3mySmLocRPSgIQuLtLR8lb9
sThtexKAwhgJ4x0iNYTsuXqswARYjn1QW+vjstY9SrR2zAtQjLGv0DZwp6SjYeAQ
WfSVkdkOMzfNvYKnwf21t/6K/QR2DBsMDUqfZs5FOjDAMrSAxwkYmKIu4Zq6lR1z
R3S4ogLuuiTQa7rM7qKfsM/aAhEx6yKRv7dH609P/nzY/iCyiAneLwKcm8SvOoov
oaS0ezI/SxwtYb8F28NoXvLVo4kNtbT57ousZ3DvsX6D+rulsEnLwQbSgY69IGwO
E6fwP9qaZLTuOjyDMw/D4eGoiZk1Y4Xzwt89Mjd9u8vw8+bKzeUgS3VHUHKxzlav
0ySBZDQFMkrUhwJFbeD66TQqgE04tjHI2FS+rNN0RQE63tQb9xmh5iGBsKFHhn0d
+1mGjwJSLgKQv3mpzdjCdf/21hpLBMFe0tvhSx+4Nv6gRkJji9bpmMNpvmak4S4S
ENmPMrbfC+xKbIO4sOFcyVG6hCG+AXz1aDxd/SjqFQldu0plAc2LBWgMsPVT7PRF
`protect END_PROTECTED
