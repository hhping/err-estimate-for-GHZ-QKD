`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Dr0+jVLdaRdwW4Z9ttj7OTKKUTPPvFTPfnnAUZCyvX6RnyJV9v2mk6pWReXCtNo
vyxiGuGmFhbEqSNSG32mnHKsSOfaWobNTWO1Vm1/W0xXrEAPHOOYdqW3N24CUd6i
8ugNKHkN5JhbLRoQ2x/U1+ejOk6b74QGesvsFs/KYW7udoq8NbUKgRMuyEdcKbzv
w/3MBdL9ipl3p8Ox84Jm3WYktHa+utr9VonLEm6GYkxZaTPqCGAQR25ocy3AlzPc
uzwS25wpothU3shl0mc0N+GqZfxVNnAw9euoFA6Hu953r6qZu/d9wL+ohdNJmfI4
Ur3r1n0+YECatTZdWpsEbSPyrVPVfOB6N7eUsWvrPVyxtPK4pego3lD8OupYoFGQ
10TjpqwZE4f+FHhpTvSRjcE89DpvTdzHxYpMmlTybVAAUbfZnR89YGs+T3SWmr1t
87+mnU27FTDKjLfTIPi/4lj+a4HFwCgJbHgAqggIaJaVhzcn04R5fUkgqgV3pgXO
FekkKDKCCYgoNrVbm78wQ/B2aHQW6UC7ZKNS9Wfp19SFCW47Ao9eKxAiMMV2AKsx
wnQFrlnB37vqs7Yj0wA27OK8HknImsWNzRlJnHe/4sYZ5Xi2RIVSgoJaiYiAmxIZ
mfZKrARnEmnQVi9wotcgVzAl9cPYpdAi16IROKjY5njx5PAbGAKy0Xvz7lLvegCo
6l9VqANorQ1nICBrorf0R5xsJ/KakDEVhgh87W8m3RDSuN/LfLOvqmzRFn4+ZgyC
YT2kRHWQYK5IDbeA/R7knGxmJ8umEhXGeA9xs07HpHHFt86VrPvHTIsIOF5CurZ3
35oO0lh/fQ1sN7nUAV/ItYwZRn4S3Ezbv2UUTV+8n1d+iGz3KQuCLEkoU2N5N4aL
4FtBj1Okfuyvu5NLwCxvi+MekQ9bwwjOi38RIdZ06AifRAQK55lEULYSF9FLWlDE
jM8mcAdWnJsuqcwT9LusipiRMdJd4VGGIP2w7mfTm3/OJrkySGzDTS49B2C1M7P7
`protect END_PROTECTED
