`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wz6uxZedAWIz61g4gW/+k6V/hkMTvUF8mQl66UsajZfnLlZZ81yjmIsHsBkJASFg
jMQTsCv08dT7qjvZHvJ9m0bKySi922BlvZ4o+iuMvbxJGRheiHKrQMFlgIeAHcmr
LWJUkDAySqngyEuFKML9TiYcR2g5+uExVcV5BNc69gBJStFkxYw9MyOgEyTm/ezY
KREvovf3pSw+RFbPGER6BR49TI3iUbfTZ6GQ8d7GiGRoWco5sy14vvv+e1MuVms/
u/DcjmN0Z393TY1LLsxcQ/G+GAGxEPD29LgL7zZsKrhmJ49WkrKJZI1Hz53hxGi1
rHbfZrju4zKSdpx9Q49fp0hWO8Axz5hE+I2766FhO5986aexiJoQCYggtT1TPEVi
XB/rgI0sRPD+etIuvmfXQtqm7YEr6vk1AUBz4TG1XyybAq7gVBDYGKAcS+ocms3z
3SxeAxA3fBL808iVOKGQIWK//THTQUcn7KuzQrAze5hlElANeVMazjwv1dzm5bYI
MnxknsteWz7U31QdaTZJY+rdq4XS1KJ/u7+fP2JRoIM4sP3IdLMw6H2t4hAMPzPc
iJMA+dQ5GVf8IK2SqxOWdYwg/761SVnyrXmKoWkIomzAHur+Id1JlqU+KbVhSQOC
MyL8lpjkTMyoe8+nb1RVXjdinu6WNOhrk5Zsm5p1UQo=
`protect END_PROTECTED
