`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fm2GgU+Zrc5k8JlnAY6MFBae/IcodxgC6por20BGN3V673bdpTvogpipDBvjuRik
4WAWn1Q9qTCcZMw7Ssn4Q9Xrt8nfzfoJBg72KM7XfHV7xLaBR3WU6lOmp9ZAoSDm
inMX5of+yxpkt9za4is4M8YwtlodUBgmzwXvdM+32z6ScL7QCF1tdLnglSRSPOgk
tzegxPmBpnjm9yptXlUxVAsIgSAXQEMrA4jyUEHYrmJQgAoJgWJVSY6uswBHKnE1
7p3XLDB9BxOZgMFtcSFqoD4UBonnzYVu73gZknCraI69RH1fsdWpixJS/N0aJo2E
uCRxTlwGMbQz7KsnjzCDdtQ4RN6g7axq3+a+7QxCVsOSv6m4TA2F7MroeJj3+TXN
gJG+W3yXp0tpflsjc/vYwlNWqezPsLBBAepFt2B7ajHNQNNNmrvWOey+SYucIism
YNWj6sPwSj2SeyVsenAlPMs5UxvoBrh+BWWnBLg9WXEC4PJfEflvAiAgyZOJlRji
3SkTdWgvZFRMRWhH0Sd88IX7Fjr9CidKFJk0d0ANV9KoZyqw8ScyceqX1fxmZlxS
O1GRQx7ofMLpu76Geufd07lQXdwPon2/SafHStb+fu1Uo+bHjzR9cgAPnTt9KsLi
AGQuy0BzsefscyKea1CORT+Vb+0cYRTQPwXN+HDagtTphu7Ud7G1YkiBqQJZUo9M
8hAZklqnnCluL5XcYC/JRXPGIAW8DJaqC9/uLJZUpNq0lsjVes7xyNM/uyOJP+ax
NxaVqd8CcSyulq5/nxi5LW5t+00nalc2ev6M3VIEs3IVuYCyWdXP4aNbNzvAcXIu
c5LUy93Js+cbRKUrmjSYfY7kxACtGSf17nZ5CJeeXUf3Nm3q261YeFiNRrKcY1uz
J5jkgGg0eL4Ch4ZiTiV2hePNY44sV3EU9QQJM2NNtAk/IeBixJUIKG065zjZi2mU
Ak47xTDNSPUBIzOMOQYFT6T4CdYBXdJfLVfHAaTzQPTALPTkZxo4qM7qH6pReljf
tPnPl1jIcdKAgzpgmExP9KHxU03C/LDfMPsdwiwWIotCMRB+tC3gH06xAfVdi4IV
NvnuOy7irtcwfSYMZMUXeY/q9RF1UtTQwW29MGuMAvd0S4mi0k/znDaW781rkIM3
GzGcUZ71jqkvI4b4AGXNnS4fFf5TsIrUMDQ0XQ9XW/HsBfrpRZL4DvMrTLI6iJ0y
/CUad3V5gAtg8kjBfw5YZCf9moVyu4OmvemrsGpkLmjFXs13bkJHjDLRVufC54y+
DqYyOUSNrea2LOmTGwv5clty6gqDkBNKFplYXaPcN7GBaLyEqNBjz8x80CJkOx0I
lZ7OlpeX8ocfTYaggdfyA+fVzsD4EZz/98zxxwoFpMLWJ+0t33pMB2Xs/Yy/h+nn
eaoWrYcPyJQOW1rkAvgEWb9zfc0u5Hhc7sM8Kbe0+tuyuoydwRuVhbaAvJdSre1x
wfNIGQ6bd3Vlqt4MB95IIlpKDcWbbJY1MdOWpAhWnp8SQnIm2gWT0ABZ9JdbOubO
IJBaSqY59w9zkvLth8Q/TgrjgmR2t65c1jxlKPaAmaIjXSaiHnUapWsDfW6cieHr
M7h1uhSJzFFF/DefrUtw6iWmhASx4lSN4IaMbF5el3E=
`protect END_PROTECTED
