`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LMc5U76ejpwiUE53fcza9qX2epWmgRR8l98qYVAD/RqHqj4RkOYoYsBK3V4S9Pgs
GnjMgRRQhZqKwOzPLeLmSEkmKxlYEzd4xIToL/EDofPcc1xsmZ3hQZFWoJ1szhqP
J69jODVImIhmKpZNtglgnwdCyMC16Arr4a9R4a8RqFFbbIpXE0OD2Ob2i+q44mP5
rMqdGx9UZ3u1wHRmTnqmDyEv3/IwOYtqXGaFBbEq2+01UVN3P1Zr/Akn3p3xcneq
B+Xe28VOcuhxFaf3OlmrA/svtzh0LttOtllQGq2/WQsbNXdJa9DUWCUmq3k/28jn
VoM+yoEGt5d4jiLTMrxn3b6mWeGy/dZCO5YCLy/8gub7QSeot74WraQdxv9zV2zO
K50R+Nfnut+RQ4miI+jb1Rqo66Ii4JGwJ1a5P9zLI8rIBQVJKm3iB0NpdGJTgTs4
+h3bbQCadq9qp4vWc1+k89ijNLhFmBb5s54LEV9dWOZa4qW8FAhb+7qzoDRUid07
zcNIjTpnH+c0jRK93cLGVJWlmRmzQouR6xbeHO0y8sEmTvDKDilNOoiSBQbVhuFn
0V5BE8bVsL8LS5X3niB0kgzlBnEZWfur5smawdNa+NsfgiGWMw/oFIoxk0rbEfi6
CfujBL6ZbYXQmwc10SyZu8Y/2QywhU7o/XETgHRhZMY/9NQsEc90Xh5XAEyydVut
XerNow97LJboleiQsdWbwdE0ox6rBw97Q3yrslZ9SUa+GIGuhF7b8FTlZ98aLSfQ
yFbkJq8ZHoEo1D1zdD0ubYKIyxKnI9ihuKiDOHThA7I=
`protect END_PROTECTED
