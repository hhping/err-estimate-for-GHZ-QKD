`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6m4vMEPQulfPr1meMsVYKAbhz5f1QAJoKYLAYDpkmOON4/sfJwH3HrtnHLax+KK
wMyMb/neK/5QgbmryopXZu8UH05uo7IDuVuKnlYcP8DXs0f2vhd89+Id9Chz3QMb
np1JpYhWzyjuK+vNANX6E2m8T9RNx1T3Eax9Aguxyhchgs0cIpAouITOqxLrh009
/8ZvGUE9uOpxTNyv3twrrmDVthq4Eq7D8M7U3t1IvlaXXoW1ncrY/V6aJDAmTKFT
CvJlnSOuu4myoa3RAYd9A3XVty+aGI6cTzApfr6Sqp+qS3kAgGTkcfOT+u/YlxO/
H2K5TjxKAz7kzKrWvdGFKVzpAq5X0E6NRyc2yI08l0jcwCXGMnFdqIb2wbCT4SwI
aYPx1GVZ10TAqhrMHaVb8RbPdpMrcCcKwpbdlEBjCLp0xRBrjCNVP2bQ4hgP6A4P
jf366L7UsaMKsNAl6rQXveZFKkOk4CB4IjexU1djVP9JKDQ3yMOV6MLntyAuwK1/
pQTCiWDg8Hzo693onV3aOf3qllkQ1dmHy8FmpyiZ/Wh0P1iQBz8NPLiQXfKR5kDA
qw/+7qCpliuw26+1D0ThtY07ezR3F3dJXSl0/5qSfNsvU2kHh78c/66WUrhn9syz
6hS4yu2+NoZABIOrE6gOSzQ5UIare+SEdqgtwTQe8o9LGOvNv1bUe0wx0u9bc4Vy
EihZPinAxsWby9z4qS0khMRQuoFIp7ZsDZn32ER6R6vnJdgPvpFMEzEZFr+H9MfW
+IVgdFzvRGJllVpLMoDUch55tUoNN09OPAagdfR7wa73RnTC6XrC36+b0BLrrenc
jlHu6rpdYKAmqa/dzNtAj2sbsgWR4gkl6U3Ot6S30ECxnu/k757zJjOyl+qWHZcP
eFWMEDuTwAkK1dsXGIPpXG4/fFA6RIyM71ee/a1TqZW9pQj8n2DyRKG7gEKv1sGR
AIEK/kI/MUCB/vuZMuR9MXIUWZQM8LpSFotQ+DdNnqrDcuwLUqIPFzO6UHObq/lX
2OLG3DAFmRxH+2CdrkZtjf6LX+e3eVwUP1wqgdYxHZ/pWH+Bl7a77M7wC6yG1U3n
ZTz/Lq16X5dKEMOkrgK58OSOUTZqHSPJYNEshcoMJ5hog7SECm4iIMx8PEQqR5cH
JT1qWBq8lfskW/ibzFh4msbJKYony11YsjelNeY0bo+PPN7wIztFgGKzH+sQAJcu
cv3De2njf2ahkhPVVd2/nxcgZh7GwUHicHIDYXVyQ2OjlkcFNQTLFqfgnmGsxUFC
Fe53VrJnDXuaBOUU6ft01fOUXReWhsEgVw2C5UL+YJUWHfkxuouQiImcRaPrA6yE
QToPX5OljE26c0vqqNsTa6n2Kkxcj5f2yxQOuVrb/SK4UoJJeTbkr7kEXqutpI7S
2XmXdIt/5DjxDrXnp7rUULAj8o4zQyA9LhgiznQfSVaYosEksSc9kpxBYJoFIEZ8
CZJ5VVizD73H+PPBKBJunxBB3gNVBs07foS9Om1y9rTFl70uNF1WFZk8RGJyEj/q
Wl3xs+YRfkt6R3iNcIFsEsKdO6QHBys4CSIEhmwY0Fkbvh9IF++tLAPury+bNLcx
Fo70y6xWfpBxqpejEGCN4gaWTyRHy65gji3BxK14QfNDjVfwKTkrBexvRxMC4g3/
JdlJNC72Pfc/ccc16Yi7TC9XX+igyqCxTzYUTfdDpdmqnKf+jqOVcRWTQFf2bFuv
hqWd+SbL697UaMC1doZNuG7I6S/fX644gho5zLmSi2wQM7PV5tYVAkWmtA9T72eM
QTxctYD3wNe+Av8H3Am4Cw==
`protect END_PROTECTED
