`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rBUDhm9mLZJpPHFOB8cvgFraYkoqOajmLmCmFAdbaMopnzG/ei5GMcIdIVy1i6hU
Nf9b9Oq0GF14OBD53uJwIWCfTzG+KeuQIQhhRPgWZFyE23GmTL4Fx+hSZnOZJSx+
QKPqJLqcJtrZxAF24nd1RLwjgLEm/3UhQNtTX6yHtYDwVd0KlRassl3tUBac2/dq
FpLZvQCrNeR/MOFt6Ptt+kR1lOfdKMudZrUrAfgr5xZHULPi+PREHvX+HXxXHUHk
voQtqvPAuDOsraU5bHJSGoBSDVeL5LE+KEFd/X2zON4ewr6Hi9/lAbnnKcbGSdpj
fBEwHiHGjPXoTWlLylGGiuDHxNDSI/e5xCUU8sF3H8nQU7oRMzEBKV7aWOSSrYoo
yXh4ictFpLfwrEAZpxQHwBS2yP63wuSC/6RKRHUP5sbBS+3gfI/wO6XhHYTypFoI
kD6pBEilbzpow7Do0yTugLDShhFXjIhdQCAgKG1R9cPIgX+xkOqUgMdsueF+z4qU
f61Vq3CXlC8yc3rVye1Pr7vmwgqwrwVfU15Ci2OonGVdxiXuZxo9WJozEZKOjweE
m72ogMPCr6Zi5iw3qI6as2CNDUgdKMcQt8AL9OT76JzGzQmcPlUtU32528na6an7
vu7TabdQtE9AODyi+PbTiRS9oVWIlemSiys+xaSNmLn6m5pROFa+pMVX+UNc6iJM
VGXSUfU0XcolbWotvSl4F7P0wVtedPVgRB3EmZwDbQ5lKoJvJ78YDW0KuybSzQqA
`protect END_PROTECTED
