`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zGmysiy7VlcVpvYRMg7brBkH8qiAjDHth8YsTRL5qMDPKn80RUYBHsYTwdhLXkOa
P36BIx9NA/jQLYB2mV0c0nPJhEsPPwHyZK26CjruxZacJg5943Et5bgDn/ZXgFAr
X9w7leO14xhdl13evjElJrwn8X2C5XwXWL1lhtvQ8DBKDq0G0a+no6RlBfPGj982
CdZt7O+rledHsJORlvEO1krenHoup/QdFPZE9un6xODFSWomQfBpo9CBn6HyZLNb
otVKqmcaAQuOqTwKwLhAy4jRBYMQ39M6T4vSZveoB60iGCJigICWjqz3Z/GHniLT
9HJr/zB6zpuVbjXYobDI/i9oHF3P2Kax67B4/+Kt2KVD5gIr4wkeZkF5b+YZnTDA
euTtn1qWNze8PrzdNe88XNFjkgRMF1jC1eNAzmM4LkwS5oMv9DwgFEYA+RfJNhpb
Hwn9d+aX90HrEBY4BBfn2bH7r89lAeM7/6LEENytmWrI85ens4kamIEcke7YFVtZ
/J9x/v3bwzkjVi0veR7HLzo0+jnd0gOv8Q87r39f1YCdmVIY/nmTY/ztoga+lDsG
EJ0VtfgcRKrAf2XilyqNmORYAYK0C1fP9ERLZg6Yp6Dfi3mi7m93bAGrQyhFjTo9
56/QvLmT6xFjOY2sxbkVB9r4MnanytSN4G5YQC1H/rUz2SDv6vaAeJw5xdaHZFtu
KOAuguFbKFyQrpLvTXbE4H9+68Vrw76dN1oaK7SoHCxjZi5UJ+CQsmNNizJa63zR
wRsuSixQ35zbCjdBoWGBLJ237rY1MUZPitFNZxiAsSbX0WhOnxNgthQpxeFNJX73
ZFVfV3QEf9eSsX2R0OWQ4HEXIAKGz2LeUSW7524OMHASZ4RHF49xe+NsDyTXGECW
/+LURY0bhF8Hq1468Dd9eR/QMCZSWgna/kSvDgmJj7VhKu3qRMjvWK4px8kQXmQi
3hthqtmGosHP2IgdgXQLTqKhHQyLVUrLLyi0i2WIA7Q5q7AsrKy/TuroTjp0Ytxj
tyOs3Yvy1a0Rifga5fP0U7CyyT/srA9QzaKsQe85jiLPG8UzoUzeGPJ2SeuZ/U0d
40nFXNRVu6xfkZ7M3Hnsx4GqYWXAjkrnKyQ2EhfdGcxLoSmyASvWvHFWrUktExZI
D4MpgV/HBZmhS43mikK5B6A+BwaBojggIVR70Mj+X0+GO7+l/CruhK8llvarVQ3+
Hrf7pO+b40OOP1rdaf9X8pmWr1pONcYsB1IJmUHZYRbCDZGyIIJ9P42RYsxXpYR+
uLGn1SIVjlW7y4yjpZiNZCoCLf/d+AX0FWtoBZ1i4T+oLGrhHNnLIMTvq9vnvZqA
xDX25F8E6plBVNbY/AoSRN1ezyo29Zn6zfTpdqmFoiJEsEty5svIHb2Pb12VGuYF
tjTtUnOo3ERxxQWV3AFa0v3nKuhPb749HbsgNHZxBD3s485d2U+MOns8F9q6BwRZ
PnJzUT/7VI3W3tIbQGyR38Ee50C3Lbkbe0aFI/7QeewGHEoaJ8LC178AzF/EdPvF
NjfgyekHWaSwAU6dDc5XaH1u2fVd9i3B6fMqXkS18iDbhuPeUYA+xCjpcYhb50ym
CkyYt++1DPJYNvDKRAGYWUPI11O54rGBAMMQrgEwUALodSi3DjmDjDLqkfjLkuzQ
oJej61FH5cq9dY+KbTEdm2Wn7fI0dwfALGwGiLfyqa4ahn1kDm167w0fUMop/Eae
Qpaea8skIcPRCH2PWioIzdgjEl5IX1syj3+SqMKOTMwINHb6090ga14PENNcb9PJ
59k/I7SlbfHhWaGIQtfGSqL0vQodiG57JMfAxx2p9AuSv6I/v25xnfIQaqCdeiiq
9eh8U8y155xWY8T3CaRrRomapt9TbkHBQ8iXMQbzKwG9V0rWoIY9A2uN8loSsL8D
dko9XfBm3EJO1rIV4xn9jHW0OiAbJW307wBHuDXMQlh0Acd7jvFYfm2ay6B+tyup
bWUnpgo6UyBI8QW2sUq6jOk/4UfcTO7ffkhHfOIhA9iAt+x5uMw0SLOkQk4VHdgP
Nfg7EDAcSMr1YSuo5BEvlAfY1ppiGbNXkGCm5cUD4T7omH9ywbIh7feaNbgso0FM
/GY3Zl+BE0FvVUWohhZJJohrbsQXrpmJYmLb4+CajUJB7fFdUPRCuAukTWRCb72C
7rIvMDSkpX7tRIHqn/AlC3o1u3lRtr4D1BLfCxHo0hLVk4NG570k2G4aLNXzSm7/
TYZaKNM5TnfpvKB8bna/Vi8kK7aCyocbn/p4252VrT8Iwql/Fj54xkCvyl+miV6V
EyWENrZ4ybulJmvCcDYbI1GskpkUe4EK8eW0Om1HRtIiDtHlHUv02Tkcsa8PZ589
lmyQFoD04HcETyf6hEYbtrS+r1L/pxGRDHkicKonC2AUc8T+VgIklwpPrt54ddLb
FYnUBV8V5hlEQy/8IY+GEjheBNW7PlCqD2mGTvIG9V5yJP1U9L72zSvkU1CTdo+9
MAgn5aR9cscOzyJP9zC5Wv7Xa3eOQ0K7AOW42MK8cF9cIAN+DH0odlsdgM0tcTGP
7ctIPzRoiDilEbnmksXWbRgAL0Y3wbn8Xn/o+MYjTQwvvmUJ2to+fxhss4jdHVaT
jz7udXrg47xs7tM1SwgLz/PoMMDQCwBgUNneaxEg4u21lsnsViORthlmBZ39aEqj
QrzL48wnuwwcQ2YZ43k3GgJeV1nC+ce0BitB5FaIhj5p0q5gbGmfIkA5DesLOLTe
ibb2D06foLSxdsMMe6JxyCoJroW3PuLN2JFcjcgrqwg=
`protect END_PROTECTED
