`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gByL+nm3BnJXMB2RHjznnakO8XFlHdOk1ruxpUxvKf8yAcYoTyd5QjTU65L0x/JP
tiXIqV3W1QsazE46IpJu6ap2DoYEQKDQqviDRcBffuvC12iVE3Ef4LTijkcFUOhZ
6ZAwt+9g5sMUTtgYFeylFTun8+dtxryBZrDov6ecboUYNZGnmGwxRj6N9sz1xUDv
4bj1k/uZmcEXPe8mlViH+Wq9agEc1j5jD2boIftb/b7Zib9d0ndH5V9F4goKxPZD
YZN8FhtCUHE3OLcayVGUVGgQVf3ZQH1sSZ8uZm2RUQsrssWmKU/Sp1KTPEN/w0ib
CMu63FfEiZ+aAiOnBVNLoelNqs73xLdmjhTHeyCL/Gv/JRR6lHk12E5EP4eenNSE
j9d2cog857y6CpI29Ge0CcL0lZZY2kOVzm+wJ8i3hYxWiPnrmt65VKquIuOKe8Ak
On8RnITlXjTKlbTNwcLflryz7DPZj/JrmYB7rF8gYEwE+UZFLmutBQzo+MtDJJlr
5QbzrEyL9shtsB5Vo0up0ub/SHBTSoSQUfEE1DliqLSJByIDcVBE6pTkjfK1+m8j
rW/MTb/WsNal6Ov5Chod3j6zwA2UeUyB20LIrKzCUeSQvyifDAzMDOZdtT5xWvmP
sNO0AwSlLSMs7hxibqvf4lTAtMW6UKrd2jXlARlSst9RI9pdfh16GcdxJohIHbmC
ZmS5D8kpvDP3MOkiaeaRyCfyU1aG4OdEFIYr3t5PUigZ2/MQ3pWZ01DZAmTductD
f8zDsNm8jzlgqxMdocAumzDFE6PQTlnUDipnIRrQDlW87hjXcaMVmjKJAEFg7Fgk
UkAtClIcGkhTBMtvUQuTFNXBwDpAQllBZOQKkLL909noPAa+cOxCevwL+2FdwLEM
LbBv0i9RCcXnJNoM9i/PKGE1l/7/fGhefjR+4nnq4MlLtOPdRuv8JJ3ztAflovE7
w1QBm2JAxqXpHn695kZb1N4U97LZpfPlK0wkQ++Mkj5f1LtblykR1kCeCtddPmuo
ddKEt+cpdO4jzIvA5B75pC7IBdgTnP6xi9y2tF5sGCUbOttAVVtp3Po947kGkvtp
t09X63G/uoBMyExoPjikA4XrSeNpRp/HDdTqKfR5DF3DPJ7W06weO1tJiJXhXMwt
PiCtmEXT6cWHaWNmt7EYnagTCE4+Rp+M6Vzdp+BBTHY=
`protect END_PROTECTED
