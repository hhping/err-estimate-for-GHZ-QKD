`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OH2prOdSXyF+ylq4AJ69JBAswfI9ParjGlh8bvcFuYnETFOpaI5ROR6dQ/u9qMjh
dvUV17ld2RBh5SJGo/gCMoyPAqGIZNXmK5IGvzCehCt6YLfF4ezX6Ag912dQk+D6
e6HPEzkhvRwjKNenC4bApN1MmdLYsCEAV9P0kteNaEDL7b051Sjnqyvt32w/v5wd
YgbyWYH2h6qg9rOPx6KN/yEKVH7R3OQY0F05Gxsa5CeR9jnXSNUpgma2QjTnX3gi
rKHgMVGExYLybTaMsoC8TTcxsHL+cTrK3eXLwSJz+//gYExGfLRB40teH7vDmP6d
X5YvuQia1nNKUE84YLmaMClBJcjK86p/fkU/zsDhFMSp6b4jBP9j4CVXOUhJ/11u
2HNARTHATISSb6zF1luSOa0Inwj/gk8gTb66rpVscic3eQYphnWJk0yltK9QJG9t
X8f/pUzjNRO1x59TRnKWdqYK2CrPKASfsvFpUn/wjPyDSVio9XEwrmBxw6CvywPU
nMgeq8tqihb0NDOF+7zixB1MFBo16Ntwu1KAemEKc00=
`protect END_PROTECTED
