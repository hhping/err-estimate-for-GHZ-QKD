`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WQxuAGAuMt3ntDB9z9RLORmS1/pLW/c5AjlHqxBuMO2Qn3hXw34rGoSKniOznyYc
1QjVlxUloJ4PmwQFPOyhx6bI+GGemW8AuDyZcSbh0wIiEc8DjMy832cV6kgX+DZ0
364GdA/MzmaeJSBTA8TyFo/tpgAFpwTVorXif567sOfOtH9AoyDao6Y/UsxifQpv
RnEnOGsumB7ZCEY9AdUIS3iClrArDUcFc6DNflNqRuHqld+f2T87ydiSqvJDGXYI
nodVZD8dsrivVapRRztRzqkyXP8d834tKMVUyjpBNVWj+YSt3+iVnxG8XUh39vHh
vCg2d+xvjw1ZhIBHzftrn7PFpf9mb7W7GNJeW7QvtiiQ27HIa+a+2cDtUPHdwyqp
SCK34Dkx1B+OpZkVZAzr/pYazLC8M3LqsW79eZ9YyyHwPZinN78EhnHxv4ZWeYvo
FO7B3K4EqaESAV+lni0AigwhTFXy254tQeehhXhc1zLjyU/nosiblmGZQALBtqnC
dyBWvzNWHNxr+KuVQp72aYWSh+45r3CP/AAL5hz9chVqrNT/2VpI/voq8jl3R6vP
9vmufbLviGmoVHf1RdVcfpJcE21I0h4AGRYH/efyjJrOlIXZvc0yw4pMQVQizslv
5xcBdn5KbTy7E1w5l8WplAXD7ACJiIO+aHCTaZNbomRgnluoVuiZd4UfhzOuOjXA
492gAqguAmii5e69cQvPRKNiNHX3ALeJIo1fguWUwwOD38VCVGWh1sb1Qab2lRt4
c9OUnXaF3f8zWIqW3TqnziZrOtG4ST9cpmUANvqgYgfKB/IYRnjA3uay0nLpctxQ
7iVxJEGdOFxnk9bfvcTe+/xcZTco8g+DWJsK3McqSEMzM4N/14wpBL/p1mBmJZhe
zoAANZ2ZTbNSfyRx3j2d2EzMc1+o0jgO0n2WpHU2tiCSLXuzF/LCrYVx6ysQeygC
6q1PRDHJSYzuiQDiygEgofXlpAnwrVivGYuFWHfTrBjm3aGn3lnbjuMNtsrS0mX2
2idQ4AZKzEWT4EyVCIfApfW6nySizKgFRlR4DXfa2REP6KPN8JJWJzDJWjT7TQpT
qDgQOeE8SWQlRC0LPhwl9nMUWa11JL98iYgknNuo/DD9CQFXu6V4mVsHROaq5U7l
98FQMZR/YJ3xrhiNPD1omYUoRAMD70n5ervx/0KSTjSm3/TAuAoI5HTfpK2vtFUr
Ln5WDv7MI/Z1HV1mFuEQvk4mkBKFy+IOUlBMeR2Ws7wB0RNBRKHqYXUt8aymbR9A
kPrX3qZ2bl9aIQK4ayKIZWX2ILIYK4tAP0NzrGfhbAotR3ocRGSz4bTFdXZsqP69
jvNMrrDC8/FiOGPEBG69RiUKO36z+JXjbCFsNDNdofZI9yRQBrCRXHn/HPg2YwVS
EHvzE9ViL2GGiJImps+4uVEJdpdUWyg+nouBdD/fluHwwQUtrv8FYkGArPiYXLrL
9ZB2EHyCTmLEy0xB2LBnxMZzgbsyBzAh22cNpRBi+IHJxN+zxsFRph8I6QSjQwGc
OaiTuCog08zBCzyWf56CBuEwTbv1ZgivxONDhqrjUEMjDaspHyvqHALmR5oCHeHe
Knz2fobIbGxeAd/e3fVmGfd2HW7fGy4uyZgIsrwEbInljHPt33MHgKwv8K6Hwv+C
MVNbEhxDyrbZHadJCivXHgs60loorBK4Pfjizuo3kB8/CRdaZv9Volxn/pnXIX9y
`protect END_PROTECTED
