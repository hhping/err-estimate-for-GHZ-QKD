`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vTlhU+CsY3CCfzXY5cxa2QQ25VIA4s1Xo8C2p7h+FgYRTtlnGObDcBymSCp+F5IK
1ZdpuWQodvE1DDaRRUmJFrmC+gGB3LDskvA6yLTbrBjQAmKM4aW6Ect5uuP8cPcs
zociYTOHGIfDf9Pk2EmvxZ5nM0hkgoq86gr9xfWc7CwJoBHedgHTX3KIW0woXNEC
iH1yTX9EAouUddg2s/m6xMW6XLTI/AyM5+eTv6wLNngM2E/LlQAiQ3yf6a/ljP3T
No7mgorYq/nno/w9XItk/zDO6KS1evRxQL0/Ts12GrNBboaPgrvmYzBKYr9htKRS
twFxaYNBuslfUAZ3GG2QZOUxI3p66dln2+68djmZ4fWEXBI/5XEYYKCytI6lPXSt
Nxe7+ImYM/UlXtacd0UJ4S9YiuM7lo65SA+nGzkOvYMjM9x/YZuNlqb9RFWI6KQK
w9k82vd7MneF2tCZelZLJbIwMj+lm72yOXMmuKHpW8YV/Em2rky7OPP4ThWXuE/y
0pZ62UzJbx0N9SdVY+oIfU7+s72CfaQPxZKLf2XOc9tcQJHHd4Xc1ymoF02UW/VM
hMRzJuvA9wexWPNFEjypSJhfUpLFp03fK4kXB77bgL2ujURDqcKt9iJPfgYzV2ck
jNKXgFIBOi6nXEdbj2JAAohY0EjIfD/7wiRcVHxMLb0hUdC4xold2kGhFwIia/TS
hq8sb9V6QRt8k4pu6bWonf6DCZhMd/Urjbn31pGjRQq+725LojQNBj0g4SMm7neP
OPlpC1OFwVf290QT6BzH4xRWLyhtadieXc7vMgXvL6VmKap0kvFbPouNYwQy0pLZ
+komHEy+Uh2XU5NUQXosh1sP73guPfQIer+pBbMuin1IPAe5hiKK/JV95Kwlmvbt
r4EV0qfHHVRRPfh+BzX8GTi31IbGE6yh2BEyeHBp0621bkOzaL8b322Xc6f5KOkZ
G6Ob3smZWvHC4mKsRS+mXxy9y/Qez3a+yX2Vl+Mq86HNpWZ3yWew1T0dCL/gHhGC
zBQcxFTVO/CodUXeoEkZY/+y3SUF+ed80zh6Zx9rZFr2MEJWcMeEx2/GM6pzWC4d
c3CAxZXNJUL/RhL/zjJ+0EEjOZ4ilbdwBkALJJl3UTYkX83fya1R7awJF/mM4/51
TAp0iqRN/2HMhPLufnQUv/IxIktrAICxdP+LnXqT9O9jGaadwz1go3hfGDKjrBJP
Uo/nTcJWT4trmLvNxdUGqV6SQMK5SBuXc2/jF3xO7eVfaaYiQG2aJleZsnTmAuU3
J8OdMUNjtP1OPKGBkqhuSw==
`protect END_PROTECTED
