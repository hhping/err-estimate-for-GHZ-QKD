`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOjyTTCX0rJtp6A3offeAdJDfbt3y7DO6CaXreWySZMaV7pLIF+t/TU1cQ+IqBn3
vUgz/AjWFm/wUfO6by4X3r5g1ACpJnQ4bPGseOpRMx7ObnCRla3QVk5ZSzpgweaV
BJyUT3/TdlJF9Dd24pCzip3ThQ/QAUHx7//UtYDPdpeYSg/Jjz1lHFyuL776A2AH
LSBKMFKXfeeN+H81MZO8nfTptjCs/x6cztpW2wnVBJIrFsnJdzKKVhJRNA2iypWl
Qbr0oDShM1eHI6WzoIhLKC1uywGlYTeM9MjRm0i/JDgLwxq2mfJsi8U7kccDSVgq
hEVfz7BWIo9eIXNFH/sfX8DuNGMD/FUN5xdBhHaolPXNmcVHzp06zvV8Ipd9iHjQ
680zufUrpNPtfuS2rPaDVVMsf+uHWfezC5L2AZUJKnrZhFNcwEZ6aGJcCtFu/AFP
0MFrAbqWqtvTrLluE4CWjXs5Ns7VmIsbXvSBEYFaYLBJ6Wc+J7Mvo4gza3EuvzrW
`protect END_PROTECTED
