`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxeqHI/Ii0KkUSW6PAa8ZMmT7Zy96NI2nMUw1yeOc2xystC62Gp706fI2nGAp8Js
jO/xZGIRSJWOG8TBau/qgrps08IJE5n8OydP4VcqfFVn2wuaC18A8Cxt1h/RqJ8B
/Myv4pjcqTtmk3WPOPmefP+rx/zARN+L2HTy14Lda9ur+E/iIcG4bvZtmSB+Pr1v
aZqUQR8y1NpQR1N8FA4HQR03Ne9PMpdTTrsPjaDpYSny9M9thJtJMaTDNfyf5xf6
czFc/X5zaUn4BqeRq5oXw0MEF7uKkKaMLF464RFyV8919ZWuHvPoXA/bku/jgd1e
7QAuSKISTgPNH/EjJccyCI27BYGYWFksV4Ueu7MKhrQEIFSENQIU1W97luM5cg2l
AA5DaEhxsKrfImqiWu0itjjuKBQgUaZGD9jlHeJyHOrZN0mZaW4005LMzBOOMUHA
kl1hsDF8WVEUhW3yMT5PdA9dPVflydQFAYiQodLPueA6GcsG5DmhRoSKvt764gKf
6ZTWb2hnWs3mlEPRTxbQU4lMJ0ZYp+ZNH0KihMXSD0bGd/VQPUrsYqT3ahYY4tp7
kJdJjhhsdgCByXn8GoPROVtAiA8WPy0K6U7IDiUo8F/+/J0vsyS0XGd90HacdvT5
SOSAb2oyNlLpy1Rrhy8CLsoRFzxsCTbUmcyxgnTGeIgFI+ke7cGusmWv8Xj7zRMA
QGerA4tAlozuGxPoD4fVpfIVtqeRhgriHXxd4zZUVykKco0qgQZvb4+Mi5lTGo2j
Nvpb4Trub/WpgVBJ35x5BSBslW7qXPTfToNam5pGLaAnxur3/L7pfkEdTfAtIP/2
0gHr3hAsnRGHWs1sDpBWalwOkAwNPinxyLu7ekV1+HYz7/XpNE/9p7Hx+0gPRQNV
MEfjNPO6NimJCulwJ3Vo53kwADBrDoABNRB/D1CFrMSqUbOlI7t5d8rEcrarpmvC
blqAC/pDEwN82G+NkzKxnNNED5Iry3yjV3xJaRJKxcNDtu9scJydoOhLcqB2ufBK
/3QV1MIkByaczmJJhKkuvlmt1q4znlbDU9yq4Zet4pk7lEg+74f/A2y1fvHeJEJM
/ppBWIbqbTY/VtXqDxTHZ09wfq74wZ/WKiZVvPVfBhOWUGYa2mYVO4ArFgyAC6vk
PrURj6C/viFiVPJJsmHvITtsA8kh9kucP6ids6PKa7BeQc+BxG5YAAOuvqzuPJ81
sccH+rCTJ4WUdG8l3uZBsQwiGoQCnxauKQgr6gNbQDKtLGe1vjGvrH6qbe/WXVmT
rk+u5V93kqOCNiG3v6hKdJTPrR8JSEAxB2iDA5PYp9xv2ewbzcXGCnGaizbdTgwR
NUrCETDSA0hMViLwaGeuVi02Bc5sfd0GobnsEhlGLg4gGECHx9zMsXQzD7t4hySh
5VyB3RURZ6aHArfBHGBRjnhsbeEq2Q1WZm3KHWCW7GBC1GlFhC0Yj0LG3tvSi7sX
mxRcdXDPPTVopp/Fa/nxsnX3La9ezlzpgOtrY9CnzsOKbIG8WCBMF4XIu+ysVpfF
HYWwl4HonYR+w1xS7tE+T3tWLyChzxSB+PpouZd8qLrCmAZrYubweHNKMNiKXGs/
RpOrL6UOwg7B2NCZPI5/ltF1277eyLbh1f5bJk7QTTUhAEi9pV+90vYRBF7wL13F
kyy8mjxQTsd7wLDdlLpYyq5qvtilTa2T1DO0GnbvMRvLE3fKpkLPAuq4NUOvFjQJ
wNBtXOb6P1hRjtir6fB3b283MzmX/VMMqMjZLGZWqdw/laLozxUfWc2956NPkU3o
tBEPAQCMd5VqT65ggTZLzfqtzds+oGI7swpQCOng6T9Yfpzy/0g3SMEPwOPZdYjq
BjQnVjaPfN2LmQHVxMZfuER4c9b8oyc1SfNnazm/AxWoQHrizIv4UOI8i0rydfcF
afyktZj558eXK9HHWzxcLQrHs7lAnbuClI1kLC+fjOfHlARS3Oz4RpEBTNh1YVCm
USEArq5R3dCuIp8/Lf+h3U/4i2TjTZspyp7Msf3B/wQIFwORv74ApI1LZS8Z9hyZ
lG52eFIqTaeQMjBgzvCBWcbWbzrCdpMozUAElB+N1OwOSx8NviyFH2O8jg7CNER2
CY3oIS8Ln4ttBoHPW4VM0R1vxRZRQ7+9rdUg1jKE4ZGj+ncZM8/QeJIX2fWDRS2j
mIQrpXcEp+41J8Vt9AejLMmbMc4lchw1furm+v/WY/ey/0qBARHO6KuzI/J5I1kB
90AHPY1/Q31vn9zCbDp3CszNvYUiigjCqk8V5+Qb3Hed6RwyFK0HYerjJ8d19AIR
wDmaoY9JNjKQ32FzeKaIBUj2PM5gqVh+nBATtRG8chw6yc0tGOC9mlQxt2jlbHud
dAXUVmZNe49uAolphxcGzhRHUuygCP5X9QO/TQSCgB9Bg4m4nVmfRTCk49yKbNpg
JuaQHt+EC8vxOMHM+WE5VJca5QERF3QcRbccD8nfXF4Or7uXEdznbsDhA+CavjAl
QzhucPHlNF/sMm7tBzSjig==
`protect END_PROTECTED
