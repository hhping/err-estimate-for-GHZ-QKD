`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7GnMoaGqzZxvcatU3nQw6Jro9m7It6LlYxLotea1kGCDeQUt/Sfe0t3vT5h7Hco
S5KPU2bZQC4Juq6zlT7GZhAy+adpkvm2rYGKa5zLrLNd/nY2CkgnNsBgtxVUGSFS
fUwu9TwIN/pi0wnsLd/oB15nr4Vviqq9Clv8rW53TGgY2it5tYsx+YtUolv1JVmQ
YIHGQcJ0VIX8xcFTMsFoZqup3iRd52or8gpWx+A+2FxjHP+BkEDVvLOSzUptjNhl
e3No6auWry1Poile7zZrbk/+37+Sn6W+bgI1NmU0EhV65+xAIViE6UGZW78Egs9i
bksZC5ntAGT7xuv0mVfJt8isut6k55iAVpte+UH6FML0pSgtT1qXH82PgwsrCTrm
WsvXUIeSbkha3PCZkqFbSBrqX1ggJJecDKib2HwVDOLKp97pqNi+g2qaldKe+8kR
vDsNfEHl88KemQFa+fjIyIX+igBVFtpip3F7MWiEoAUAwA5P5kVBMkYbekuPEZJW
8fWsKTvcOwSDtm3rmoohXgHyECPBrAZgzPzKcwfGdqXRrWZ0gL6T+L0v7VAKX20K
R31MdBQS9ePemib0w21ODUNkrOtigikI5wrgU3fqOgAOF+JZmX0Xyijom9pPssy2
foOCBFx/0/vazx3x8WFdf509Kz5yPw/dme7Os/yeTy0bWt5+yjvSP28Bp3MRQ1Je
6hdtr9WoPdOxiuHa598gvj63kpPzCGC90lWdO/wp9K8=
`protect END_PROTECTED
