`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuQbr2gVTGcNzGIcbV96X1f+KYqE3lPqW3YepaiW0M4aXQfMUTwsfXfiQXBolHcb
16aZCs66sErmu93MAYmL+3sEBi/58Unm6Csccdp+LbgzOwkK3tAtBy3238kAYqGG
qlBB3YOZgZHgZI1xyrHP/VmH4JPIrG+qW925oUK/8C8OdbdQMCwRhkPS5sg79N4w
oCtdKc1MMbDlaVbBW23pseIZAYHd7KTyM8ZjS1Vy+ZVNB+oYf57FlQ+QJ9pmsUaE
Y4yNDhrHPN1IwyvcWroYrL2grXE8D4aLKLyaUzrG8WuIJTS38ifeKHAmEIGx2z0A
aYmlRrO+g6bW9hIGCbH6sjG0EuWpJ+cfiAwWqPBQn63LES4M4wlBNG+18J5uy2PD
zALzuJw2PMt9Z8I8eeogA1kbsLVo/fRi3wqqBB+MIo5+4Gs3M41zOb3nHwaz56xC
44rop0n0RYcONDwLnRDVIITp98wyB/6I8AoWiSM2UAayJ+01ciw/B3ZD/altxzt7
dx/tl3dgt6xo6FlEt8YyyPYoXsXY35tyY26tZpgB4dnCQgsuwmIbW5jJSUBloQ2x
pcNqTa9GEwMzZwA8U+J5VQpRT6B4GcGdKLwyxNKGlrqSX35mpBmUi/Mo1+CahQSs
NDGbmumkh/y7iwB57RcmLmYkSzVguCgNV7VdA6Jv2X68vzsaHNk9Zv4+yLdJoKZk
r4tQZAB7fqdNkwgRYkKWpWls+MalcrAVo6fTVOcFj6L5wyeznhymn2miYTVV4kLg
uWANDETjhEQS1Rey1sxLt8iiooGnq6/zgOGe68nR0ue9DRIgXodDyLUbtXQvp6e/
b8d7VlOiYgIKDaQluAwCpE545N8WZ5+1LhGTDftaPGDR9UpUyuduopHzrYRrf2vU
jiYOzbZOl/FvHd3HSXXbbiBtaQB+hmDyM0Ts2vWqZDuBBGm+J7u3u9lbNT8Qq8NP
AITg+vkq3ht18G7rzcC3GeIQ3SekW/drF3umwGQAjonAkEFkP5925fNsVKEbYJuc
kighaa/xCeqoilogV5YIXHxPzK6kuQ1e5bdtBdEp12nDzAOnkq//SnRaLLcR3epc
QmUc0bFPctBG8qh6zkDWgNXhauKp8nbTI2gW2/IHJ0Bo3FrF1iEkuk4ETZpCsbLu
WPzxZ3jSh3FTpp/qbgMrb4l2/Sjo4CMXxqml/8b7fz0oUvUKwGoS97dTeZAj6zpK
x1RrMCfesw55B8H2y1pJusgiWQw9FfjulUyRgL6zMjt+7XFUd2qKwxEm3PtRZYfY
qd9bM30qKraQ07r1VcB2HHX88wlkar/QPB1bUDMr7UAR2/bmSv3K6u7E0m8/zVmh
AIYH+eq1isAj7RxLv2dkfrP5ap9F7qtQrJCQiYGn5HEh1k9UBHsWwM3Ev9DdyICq
A5Sl8+0Ys1AZYq/jeD0wMhNxZju8ytQUJj0kd5yPhIr583obIiOyGmyEcSY0eBTN
ySOvNMwjNeAWO+54deFydoUD2WYTr6TbM5uPMMHZklAKdVsTJStf9lyv9UEo5ttL
i6XMbPkgrUZFW+7CmwmY82gnvQTaqRJuaESoB7AsVPYqXUFEuUJUTazPXwYgivwK
QWD7cSnqTspzgYZ+jTdjCrdsu+0sj90VUQz0FKqm8RjGY4hKhzPqLufN8ndXk2oM
r0GqIHScVjm7AbWKpAsbEhbfuuQYvWKkGvtV9HT9lpSSLUFsGecy07Rd9nM/EwZC
5+M6N5o9pK1sv8VXuM2fDKLnyKXvICbMoYAZLDgZi2hBSkp7B7syqCUnu7W0Ou22
iT2LGAi4UbZ7drW+WYPV423+9AJ+4w+ROCt7L0Oxmy7kb1O0a7SobeqGtoNMYQTg
aNr9nnNKcqm3v8OhGQqHxUSryYImg9Iezo8Fcqeswbge/RHg8T7MY2u9qSnIQH2k
tnIl7SvzJqGwcnCqiLe/44oumJE8kRbuEBRGcLqKdO8K76JN3+w+v3jgQX1eiAhR
Y61XmxvLEHqpwS5cw+mDjHJxUJOngP9JJ1+HM2jWr2r0F5EEzZUH667HNtnH14Uc
y0+Cnwl6UFGIwknhNinlVH1y9Ef2+1vA3b/r6Hg2UEWvZY0f51+5CB9Y5Ycgcmvw
J/aCjlYAJRyDxfI6dhlz7yAZtloQZuDAsyBTwUyeek/7pI9ysuI+YEUhcrcmb171
KCDa+bgdY46f4s3cxdpFKqVa5YhtEetfXBSzaA3zk+b2kYWNgy13JzwtPryWAb2+
84LuHpPOvpO0aXTMVGZNjEmVQIgnnT6akNSPS6+jHyjh561lMQXDB5DGVIhplnNk
8OX0zW2oxRVJvVJPmaLX+k1QQCOhB2jwpOVIcZJvfEfhoWbGJ9aE9pKTikiY7Mu/
RPDDHi7DKeHp+7MFUgu/5J0uwt/a6mGfjPgDBKkZu3PTKhXvOa6dboaw54gJBw3U
d6maPKCj3uCYBccNGdqt0rro5XEOTieZR9QqQICI/frPzdz4vZltLCk64nSmRnXH
TGm0M5ql3R9NjGVC9JlrvG89mPilOGDkFDo1ScBXqtNu3hCgp7DuJ9SNdAn3EgCN
vuFfbGyl8Xg0U6Jwg1IznrjMcjyQ4O1uRsaJDaJOd3qQ4kG15/cT3ETujh+ijcF2
JJ61dHrzGTlsiYM+Mz0iPyMlUgsW8MiepwRSGeAa7GZfLoGObW+UoUmlUbVqqFpH
CCSqWb32YVmWY6Bks41C5ZXHCR/sviF+3PAxwKF0lj2UWCZncLkLjlyQpNeMhAaU
2BLWwVKt456md0OKLQkHjdhIQ75XRqRvh2RcN8r1NaYWEIYsNTnx8pH1aQvfQqZY
OCtcAhuppEc2mI3tzW+2x9kKH/hB4pdtvsDnyxib92Xzw6dJ7susG7as+ULLwyTH
EB2kYMcn6QQtUCfRKCHbYNpofJcD6kVuWY7ozfPwgn9h2DnlAx9a8KP1wozxFJBK
5qO2BOhssmUtO8j/WA94+jLPvqRnLq+nRtYP0JD95dYPbKj7K2sS7eYg0CZ+67U6
Hxm1Laj7cgKvo5rcLxL+Pn0b9ivZh0d4II0sWgue4fId7QiuBAzd9sk+EeXzt8zH
oYjCC26ivCBXJF3SN5fOtdUXhXM2E9IXUfQtc5XSHjcJnmxoN4H+XzyJNbsuF0he
6GirSh3Pv+u0MMe3MHdNrBXHTv948oMDrv/J2Et0bLHjmuRXk6RdF1dMIb6qPvhG
ClcecKcAwVkxWuu4m1SvSQpICuWLX9KeVfG9w8EFZhlfK9BbimREwjJ+nxoArQd1
pNkCTBfSYMw4if+WfZF5eyEwLvdyROCix6Br6rIyNwW3ZA0ThbNTlmIzQQWWE9Ze
MGv/DaWnsPZiqDmLMSLJMETLNusOgUwQueuuJTs1w56PcwQCKWDYLEBVJLK+lsUn
yf71nIX2Z3Og319BYGUyoHJ7TYcB0j8K9CZ+kLIAJ5u7DZNK/EC2+lD6pwCpVfTD
B//7wHRw2/j2vFAzumPSRemwA5+s2tLa306ZBgCGVdmNBrBYviBoKc3mkuNUdSnV
DwbN/ySBrlosVTliK05PK62ZVREfH+OEoUBhJjpBoRfpJEVAAsExZqDy2FC5UWmm
uMaxraq3xfmJcsVgR2xKKCk54WhFklfhKcppr41UizvB778hlIQhNQvi5VWpxY1H
uNVocTPzE0sfk+prURvZtaXZrILZT5n68tu+KoXqRuCPukp3hMW1kJbvpxTIqPfQ
z7Xpxc2NmJbmYuDnLSwXiBpdLP7indfFJuD++kMGi4RUTsAEtwtZOjPDc9Ch1MDt
KwDrVtiujfZTTyOhibGliP3XJAbV4zIgVK6PLBzK2h9K02Mujd4USuQQ2IPWoEV5
x9rEt0x1uj0zhzYAiHUHGYbgblmVNkI6kyLLawtAPk/WII4F8CCf1HR99bKxnxeS
o1nzkr76gGxBHsXtd9gGeRAbbQXd5+7gegbIIDGZ4JiyHKndDMPQwFF6+AN+l3Gf
Wj7ZTcmcjFAV5BWrRjXS8wSu3gXchf0+1XIcxs+XxcLcJy4jZfVIbEATV22ubV4o
U7O1TGakPs6juOciRbfl1NHbqq4PI0eh9iwtJty9OqHHQ35SDbt8AppFYncaX0+B
5eN3KBSmQ2Ejnh9Wugk7Sd0CwIfaaoUzG1MHMZMWAz6awLUoyqaCXsbRuT2f/n75
LFdoIm2/4GVUt+1RM4X6kvUOg6Vbib1nm7rizMy7F+hVznaI/+X7g0OSV2c7APKZ
LL6zNdyE22Qhi7UGWxbQR1f7aA19CD0vX1apEL/7odr5G55vMgzNORFt+GhidQ6/
AcnscH1LvouSPxZxKkrv8BL+kTguGJkj/MaUocWbBbSqqfuOv3OVI6bdFPJtUqLe
YSk1s91Wxql6sbJr1YOM0Fbq8Ls0Ibzjrl/CIN2aDB99ucsHtp3s528PadJAFbTT
29utY1ypmwnly582F86NfaLaLzsImyqMVBQ20yl31K6H8QmnHfT4iiC1ekM5S5Ou
0w3GcP4nb4cLiqCZNqzdDYEeoMAozQ/FrBb8JPyVi6EPdhdXZoez2MSW2qKGyrgv
L5Poy0WwpM+j6hmS9+vIe9mjJbGBRii0twmqXhcpnJe2/I4fmsNhWpJgM1CwW9Q4
d8dfwphOOdRMgCRCQ7HLlK0A+y047GphSbTkuZCbtShr9qNjYS/7xLQyrlvA9COq
i9N8xIwVp0HBoxqKqwpclFq+k9oI3lsIi+Bpbgfr+zDET8qk4c9yl4JWZ3HBocmy
lfPv2hZBGdi3oJtffEwpcuSFrd9abOOOfsOWnYroE4DYFoiwOlQRsLdmDG2Wy/cu
XsFN7uC+UK3aevZkv/ekAGWepVVOrSZ2nA+j6VFnzDMRbZ56qxxxUbTfa4FK+c/F
fhXva1Yd/boIFHwEeaQt2sQdJGMjQZswGZn1u8ISyXWgTmMp4oCiCbIJbSUTIwbA
qjhcuwOdTaw7jlANAn3fFWNyJAQDSm1fyadyITEj8YekuuKAhApWdPVVcXjvnRSO
PKQC84ifV1ZU764w3+1FNXwrKFIlNHzgpTyF26MetSfnednvD15llt4luON64eLK
YX+jypBgz/qNq7MRpJcwhMsR4QtbEcNbflcg11+33ahOEzICoR6zuwkXrcYjDJZ1
9rP3pLcoxdh6+jULkCLTgQ6W1MjgOaB2axUnVIGuLExFxtDZEixcV1NB03NdISnj
fZRkvx0LpnxGHRvvORvLoskmy7cHMuyNO1QygnFs/d3jNYfKWyfe9VAHk0UWV7LO
KPYK9euHwKxdo+fLIPbFI309D+tVj19+pg3qoKSJ83C6Wg+qnZEYwWXAoUxn7xv6
2eibD9Eu8WDApR1GO/VpR4Xfn39s15iZHvzt+unP8d5sloUDJZP6+FK4+ZR9rG3o
ltWZRy29OI7fszWWAP/RpqFn7tdcwfrt1t+uSUarJ75q+PZ7BOO76hpnckzi+Vbe
QvNECWUeuzm4a+UNJbrgSrCtsReAR/HCpLG+rTn/t3M0uknjjjZpQZRlD9IVFe4H
Vmc3eqDN6wpHQzHAbCNDHHwE2zPgT93FdEnSOdgt8Xuvt2wLbnpBktvwjOLEwU/D
9x1W/INWtrtMKfAVYy6C1rT7t0btNAI8A1qGGLwRyWNrGk9iH/Uq9TgOM5QHRpu6
42b0BgnyBwyJryp02MUX3o6f2x/jM8IzCcvbtuXHPVZit+41dfz5r1xLDxtKWlGy
W+wqVwRtgoYUokq60nVyVl72MnqqWD6aE2fH18EkcT0/w+v2z7SMTIn7SJ2c+3HM
ZqHyLgSN6Fqvf/ehECqth/ol6//r/QVuHwM2vgk/xwqA/2Q/TfdD8wczfRKtUkJs
5+KdBEL1bdWH6BezlrgJBEDnrVwmhJlHt5OeU4lKULLAn9vKb7rDk0zTsFlnvJNO
hEXe2kD2RHOpt38F30392RdcecMXGvNE9HLZI+AG/FpN4TVmDsTP7L7VIbw3B13G
b7Om5MOJnO7I2K5MM5wPkvFZjT0h4gkkYcNw3jhOoNPGvLFU3CtTKzYNtTGNHAkQ
dOcuNK1bFVx/XVJsHCsXfsswvAtSV7UU7kkbBctmSA/le5XKvuMou67XE7Baan6B
OujPqv7j3PQ/vnJxqzkmbquFK1A/lO1NSKLibzIZuOe+Q1sIgZiTG0EkU2dy/7sZ
OiL0yF4c7wpTka71Ofq+Ru64BLUGdhi/Vfevst5oSA7D+tzNrtbc+tK2zUEIv/bU
0i/S9kmrvYaC6x0Rt/qxRt39/p0G+SViMfmToxAF4OaDfjJua40TOvYStOGEPRj2
r+x1i1NWmfE+uIevmB5JptR7Zb0PinolTS3Ka6KlhXKP83joJKGxTAu1EVU7cRiQ
6TBwSb+kmSAPYFcDhE7qWump985vDYLwNltgVNM3oBKW3exoxXXLul2fVasBwXcv
BcqcohIGYq7VNQQWc4hI3hs085NkSMUAoYdNeZfmqfOAnnUUeRomnG6DHcrjmH2J
VO9lJp/5gKgbhsqJGWdyzaLYYGSBvkvLTRq5UhZwhLEx9++1wwC3ERjkSG5HsOrs
phpC/imd5EaeEnkzoDHmWv2TcKUWClpMbylXNLUw8yIPfV7kQa3R4fHFMibxwo9z
9Jcgaf2BqMGZaVYB4bT8W+BAs03iy38f/Kn3kFM0qnM/YUU3RWJ/fyXjfwwCY8tr
qoOBmVT8bnINC/sX7vtmXVJcEuMeWcaoJsNocyl8C75QjcFZM+FOsAGru9CoKFUq
kgDbPBLhjFL9hQM3EEVfBJbF1SaufGbETVs8N36lELReaBw3FofF3GPqKYkmL31a
sSDDFLO6Q6YPcVu4//jfuxvjEcvIK3mwkuPpwsomUzPD4gD3xqjuJXBKKgeLOILk
9cOn7fiQKAJQJvvuXIKQD0kluB/DAlbK3Xz2RO2hJjM=
`protect END_PROTECTED
