`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXxE60Jb6ePbe7pwseBhGEZPWtMF4/Lj7D4NnfAp73SmkIXmzda5CKqw4c7OztG8
O7/xdvDm+YyhRm7DCShlLSoU+FOyWlZLLT9giOYxp9Lx2vPHManYCNO11it0VMwQ
s/Zd0FifkiS6/LYWZYyNJL0YwaksbDIJSmiYlRYzDexLGg8XfXhrz5Xc1IWO86s8
pa0UXEsbKRfQRwthlPsDQzTGweXotPEb18EHntwfgBG3mcRW4Z3xsdKe86z8MFfy
2XnTcPfV3ZSYk5dKe+nUfU1nmmiW0nDD2mAsSuO/3qeI8n1CYwpFPRt9qHkCiwLe
pntI1yYgok0yYky6M4a3lggWKq43XBrsREm9I95Z1i42SlDms3kxKyBtBdrHry6C
KzjwHD6SAiuM0Gwd1R9T1tY5uSS7DvxvpewFhYNxiMY4Osl5LAlj2PQco8RbAjU7
Fpgt1199cnbjh+aK8EaRx7IZsX3xejSp8uW/O0gx8ZY=
`protect END_PROTECTED
