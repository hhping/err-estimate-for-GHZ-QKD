`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CflzQXkMUS3nunB54f0fsTKgYHOqQJFZuJjoE73qBKxOlsS2gpsb08Mqe4cwWWMh
2syhxVrTeYzQ6k5xg7C6pRW3qRrEeiKylseG3sb8Mf4WTrTD4lnnx9qz+gwfTurE
yVE88T3Aq7W1RSEGCzQ2U6Jt82rA2Z9e5vNgXyhNm4PaTaUVvG0mLz0wl6GIavkE
CyVXkVmymIKEX1yQQeaNAFoNK1aFUQkUqng1ZxW7iCbzfHhrZr0DhePN0ID51AN+
hPIbXvQBJCpaaSHuTyfZku9Du1w9eQarMohLb1/CM/B+3uBBwQSvch/grqILq5h4
nYNzMKqNACtmt/62bak3cy0kac8YavjzvSi1BGO9OmuJ5yvcnWLOfBFY2/EkvEYX
lm4m9GkUtQg92aN4t/NtuJOeHlNjCoX1d58X6WUkoqY=
`protect END_PROTECTED
