`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSgkPtPZ26gtztxiSodYO1YSVmDqJIZ2SeInoRey+tKafz+/mbo+45zjBPUaI7Oj
N/1dt31vYaHW7nWTheVbskcxnSohqxC8l7WlAB50rP2Ui2bqgUm00M4uvMoWAJ6W
HVMXEoO02SzGm/UAWvOlhNo+vu/yn39CqywP6LdDjYEEEg+SbWmHQNNA7SiJWy4z
YOwNpa6ame7xTO7YAHvhn5MzFLdSE7YQGk+WE2v4HIZYFohSS/Sxa48cgG4khn3Y
QpelPhitQSNlrr/y8vbheZ2v9jVBRbkdrlsGDUpT8eCqKEz0NK5J9Nmy5yEnOzmq
ierpZ9fGwIt2zNULPc+NshEuK+ly4+KK/xUQe9/88PwHTo0vfK5/I7tDRRL2zPlU
9SMytPhn1MZO4WBdUY3uhvcwpcgaHT79EapS84Imw9DBki+w1eNP9FxfOPvbENFw
GOT9JrcqdCdm3sckvw3F7prwjA0t2o3K0C1VqVSb/st8cMLlHoMx0xnb6okmOhq9
4J1pgYTuCm4zLedQqP+t7eic7rDNa4nzBQGS0DrpOFJJe9hM9DdqTcwNSPuplpcy
`protect END_PROTECTED
