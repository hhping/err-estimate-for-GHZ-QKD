`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EvGp3QpLPiICRtbWHg+iFxDzjKF/ivJ2C1Km9EXoVnCflIg+onMkYLHi0YDa2jCn
7PQw8v/KL+NNlGw6ET+IzYmYPgYnbmvdkRv9Vm+5XxrACqQj+vtblLwvW0JqZ31t
7ZyU1WDW3FVrjMjdgf2MaRzvrm0+090kyAlMdF0OBJiRqnK9hP5iJe/dDy3xBwze
2yIqef0/WAsBmikN1BYZlDempV+tJsP9IDDUZGWj5M0rDjgDYXKQyXD2eyLrRMMP
0OPPBB+6dNcyQo9O2jmVhyvPqFA3X3JW5uUIuQfmHgua/nSW3P+mPKAinu1NhBXM
sBknF+q984ON5nOYa8bHc5EtHSVIXcYzapMbWqbCAiC9gLe+A2V6IL5O2oLfi3Dr
7/PHz7VoCYJec40FIUy1fBTc6lsLcYNI6UUxnajE5BAyz6N/uuRKILYp3yLwwUKF
rz3AjdhiiaWo49CPOHA+iuvIqwJQB75pK2FK8k8fPcABjr2qTSphOn3HSUmsNcM4
prIGFOqmpV5pBEhIG3gfBYNhm1W4HYbud8CBQrHeJFVIqtGQUB7w090qDslRyKwY
0OepQ67do/QvMnn6zMqMKFQ32A8aLavfyjP38yOm2Sg=
`protect END_PROTECTED
