`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWbu+sxzJAHZHde+oYgjjVNoWEJbTA5AJCJkAX3l4yvze6a54hNrPvvQ810H7RhA
Y1JD4XESjUy4AEHXwUJRSZcj+HgICDCM3kqM1vkwZmT5ugEWeno7RI6J+jViNDs4
v8aTS28mTd5s5LfvuhJbk8kK6/hHnrsMnAH9w97B8jYk409JDHm7E+7O1EaRfvfI
w7j5R6n2Fz95PB1gnTtfM3Rn2FcomvpKVQ98LXMaEIb+4P9AOGBEqmjj8D1XiyGj
4tbM3gA0D7O8WYl8/0ngwQ5dpLpQfSFBBX1qeLu9YXZN1Ei8U8IQWgZMOK+l6U1U
cQvXVSPVtr4Wy2sf8HQZCED4VhXkLuPoQaIg/l1GoNqkNBTgKWp0IUJYNCD3/Ygl
Q6Ryh+6LqVxHyk5jwDugKDmHRPM/TQaZrhZK6kvrjO54ARmVIIxnTcKaLM+pEIor
K2MzZ7j++xilceaqxmf7tnclXMVTp3ELYKuPd9dTu9auQTYX5Hh/oYWDhwA+R3I5
25qD0hhswsrROcTzkDHyG8eKu9k+CcTcDWrZ00QjReeHhuYe6H/WAT+17qXX1kLd
2OnkRSEQ3E4C7vusVyaMDg3jMTCxtEnGzBX3ZQuglieligtB+g9RaRbTPAwsymDs
82J20DoYFUC5Wi3a9LD2BWpnS/5tiBnKh2RMNh82OytyFW/y1JL37PB+YSSnNaKk
FrCqu1MoTmpz3+0vp6LaPX7xNE0m49XVzrGcB7bpHfGOjQ1nTgdvhKKidkuwRheJ
avBaH6QVHqJoTDRpfCT4JFUhw4wuwVxp9UbX5+9EjdAfrJ1s0FzoFuLvkb/ffYAq
J+8p93cdNCWe1rkJgA8LF+Zs1A9jPoPPNinxZVd5pYcOIm12XzWHbtrdEHlN9CQS
L/ImDtPLTfZfDtfBrd1peNvIoeVu4s7ALRDSEUMiodtll5Hde/D0ZlKmLLW/2ZDf
CziwNy2P4ONQkMVsCjqw9X9rofc5bAcOLzJuTw87qbpJ1l8Er0YssuJgfzR8ZfOk
4986dTgKq2602tqvHWJ7uGOd6jbzHchmgAvJEwBi9qawFxnFQRhj5ABs1OuWlV3J
9+4G4KPZTVZyUePRuJ2DCmt9X7ueHJL0rR5ZcRkr8sP7xyBvsEjcTXu7Hze2PHo5
HI4mQ9tUdKwyxV9+/dcriQXJ0gjrpkGjyZlrG+Ne+4D/XRwhWu/VeqnWbDqeyLQ4
x6Ytue4FGIayvzqvC/AYiViG9rFVZN4rSsK1y+otqckHq2Oz1iMFiUhqpKm0zmu+
C2U3WiwJQ0G9HB22vLerJ/KAa0HkCWTAVllzD3T0WcgZl/KcyJKsUvpTZT2Df+Vm
5f8S3DUxZx7C7SBFj6H60POYOxTcoRpvcQbLbSa5ikBViEXmWWRcfDuf8sdq//0E
ZL9MD25uGK8PHWBCzUf29vOuwnI4pWp6oO9baymyuFKSDjJZpQmqR5GON6yo83c4
+IyBb+NoAtLCtLj7hLpvQ8lyglGkzaqZPjQd4tg0fRvZ2TWEMBNo/LftE8onwe/y
0zmN78o+qERsanA/mV9mVDlAII04NnAdbZdHAp/+bpN/93Izxtlfzi4x95G+E0dR
P8pvyBntglY3Kt3mpdhPACh7w6z71MJJFU1oqP/8PLmIqW2xVynYxIxAS7dYDtfq
t7zptUDgGNrPdtRd3L84cdUmdjF3R21DpKPOZ8MaiuhAZRwesa6pUiNfcaAt1/ON
u8SJSQND5IhoSrdJx5Y5FFdavJnYXCalMM607GULjIPuWgO7y2AOEUNz1MpsKKb9
G1rftDzTpWWWwVrn8KLNDL72e0uE64Jl/y/E500x2lrX8O8D05fs67bT4fLsJLND
B410GswX8vn6jI/COKHzRAD6mOlV9uqaDvLtcSTgZ7P4DU50498/k4M5PBCh0JuR
U9XsJDKSFs2IF/UwgVMSGYtg0Hy5v1TZAnzYa3t7JZwdEKlVupNx1XmisF0WeW9D
y/l1TiulyLhTUIsulAJnJgB2xGuWXas/S9o406yGQAssFZY+t7Fz/o50muwutins
swEu9C6fP49YEc7sXiP5we9alOWvgrqsBGC5HLuWbpbyoC6oeXYtMO21rOLcyYJ0
nj0vJusRRjKQFvG40zfyb1hrVFPDPUplJeeUTOgei61BGlVh7GwxllpuDrzp+Gxb
frHsoc2ZwY/YruLFBEUeaIU8aXuNnt0v4LaDEjGOvMp9k3dRa/oJQNDc8e8iV4Em
0QdG70yE4ctYRrJutiKx/LMZhMDw0CfQAbthkWAVr/RFX4FWfma6SCn6JEYmb+Uw
Xph6Vl0Bkgns68nCkoLwzBiLaaKa4Gv7b6CVM+rQi1ua82P50YdBobkIDKK+yM+C
PtuHz4SFf6jVmDCA8VkJhpLxdc+gGsWgAjZuCGEWnVEZdZqrjKUzwFcRajfTSx9R
EfvwCHsIzoDT3zKpQdntQhbaydM1SAYRCWeO4V0dGupuDyFsSy7dhpVEukKXY3M2
OPj6A78qVKDxnMRmn4B/XkpAhishIGt5LLOCfxlyZeqQcYtNX8AirogTbAwvEg9h
h0hHdWAXCyeZeQ79I1mwQqzG9G57oVOyssaIgqSppLTOq4qmYxfMToB4DUQZaBcM
e8riXf75WS1GwG8hjK7Q6T6CJsF1DL8Mj3dif6PEcSjtDxt9q4quYAn6wGybUX2b
GENQgwfzCcZ8qSaCv5Sp4hZCgEdgzU92QUl8H+DmR9v3FRlvLYYK/p8vbQKrgHEA
+Y/8WBTtcHlVIkYSJnJjCHLHZl/nraoaroATjkPKOU4m69X+ioK750hpZC8XMwOa
892F6aJiV67SK4ig29JNN1XMEPbo34hxJOoslK69lXmn8LLdU0EA+iqwoPcsFE6s
niLFB2swvasg0FhMExMxRSS+El/X/uyGzkAYV79GI4odPqT3aj3hZ6ve7b+hXSFl
NXBmkj0edHoehXW8MpATRvMJn10KD1hh4FFAQZFHMn5oxAO2EFVv4E8MH8bDPydw
mxK+IMOqpIYsAAbjBPrt4++Rsc2ePimHsFazBaPFvHz4kGkvpe7+GTR9fN5Tbwg8
JMeEi/kZMDjAW6BfqwVnUYReP9JYLT0xmqz/3MuySVve6wBdAVP8AUF+KQd6BlDq
UPQbp1XbFnv2QsLsAGPpDcGTnhqWzSfUIFpWYLzeLnafJo8VLtVJel0W5SOHv/w0
6azOSaBvgHgvTV8asdbXL/Z+QgG5siM3gicR1lLfx3I7sKoqCFzbXczG0mHHM3pZ
R7LQq9heLNv2SMQhEpqtqrG1vHslxcr6AACZrEO5FTeZtwKf0yfnbUE+8Ji3pt70
UGXp+YC6hqM7NGF7YtkoqR3RpqT1ojE+mtEeofOSPujYCU8yXRdoY6aoVF9sEMa+
5EwKnZxMa4uw2tQzvfumZtr9K9EEPJuXm3jMM87wx7QSWaugDiBqCCHNQrwn7rpn
p65hY9iQTNTAhaPNAmPrJxSeJKGy1FzddjoMwzhm5Tne/oBC2fzTYiLXKSEobi79
SPOeLLJSqczT5kSp5SoGPttdMh8IaoQnRua9125x4Y6b4DeC1oWwdfY1F0prGRRx
/e2a1P4S/ZmBofQXYobzl/uTlX1YGHBXE67AXWPHe9qeOd7uO6Kkq4y4R7+V0m8f
XFNCzvY7Z5cCUbhzi638eLt4229XPPov44QekbClbcYBx6ObN42D1ANM79ZOFBrN
U5P7YNY5HLK5zjeHVTkgVY5GmfU03dniB07FCkMCElVpPSfRNC67+65vPWNYv8wF
q/aLhG3Jt+AK8hKvLI5qscVRzlMkUAB0ddUfUbDaiX8MjEY0H5Ds3PxjJ3YzU9XM
2Ni+/95f1+1uWU/TDayGuit78WOBznOvQmkX60GnCcWeJLVjnC6ZTnZ0fnb20WNu
z9dCS53RpAAlwMHglpBs3WSixNNC2zPSDX7FuJMnjCG3wb4HlnLYPJ9q8Oiupj0j
qJk6aQ/Y8LhQhVUlEpBeLJNIPiDcLgBxPl79blTzKiDnwDp/bvdNqiNLlQdLztX3
XlQsrNGIu3uBC4DGnxODNOET8rn0Ei3C1KVR3xipkzLxuzHGCJB63IvPR9rg8tEg
gRDvBi0A6wiH7NmGaWUZ8wMQRc3cq6V5a995h1W8pFboD0V3nYxaIbYOu3B70GcV
wNeJPZgK6aua12cYcSipl/0rO+xOrGLbbO14t0FZRsdjdumnC6EXj1sElJRkTy47
KmvTQK0L2QML0m+ym8k26JMlcGsqKBXJVKWj4lHTFh13LncZ8AnSSF22uGhSIzZ4
fZF/8kszV7+uhT0sxgYu/o/++MENkedsa/tjE3gkUR8+WMVRT1bUqd4QwmclJqrz
gxj2YSBPMn/KheE/QwCh3uAaej+3WNFlRobHtpyjURH9UxJQH62HPqW197qSlRdA
NmSTfibLQ95LkylXa2e6s7ES36ZAzd9tiXt5u2AGAsGnwFZZb/a2jrW9AincmaDQ
mB6DwWaT08+iSNKLPZx66m/Puc8DHxeY2HeVRJFT2A+jwOzQF4X4UWnvBS4LBCfg
ZujZ7nz3C0svfF/SSljTQQcNnouH98WPXehqQOt9pu75q0MRW9UFgxc0OF/TMQyr
L8CepCRyLsHZm80NbpnY/RZDCwzbcs0Fyg6FRuYNbcBQltGtkQMf4z50LN0CLYLR
F83LMCvWy/cjcAQmShs144mH9ENk9Dsi90JKzn57jTuFPExqI6eMjmqOW53hw6Dy
UvGgfeCGRovh05mkscmce/KJygpqQCjpf8aZZnfEEzog2v98yXPEGZ0bL4zADUlE
hMySHUansBiISCCKfpEEROfHtdHE0uaaS5DtVbZXCsxeHpbXIscdBvx3BP3qNl5n
LsJoNM5P1ZXMIgXqYOO5BZx4Mp5YoI+r4kolimaD3wFjuGB9U6CJo9WJJlfJtThd
Pe25n7WRUB88u2DSY+rgP0zqo2E8cXZbFariVqHfFQ0usEl1N/219nk1sWBvYynK
8FIVoh3IEkSs/9q8c83Is9DcsMd5wFX4gr/OJr3oy2A0Xgw5RGyCT3yp9Qxx1fjZ
7I21jspP5hAPVd0LW78ZJiG1qa4ZbTdlaOBQf0vOHZe+HbbMiRWphIZZjqpmzTLI
LgR2GTXKd5Bm0c3BlpN80oYeMgL91oQowTFvUnJ4Acw7+mKTGGwXcUO2Heb1ygwe
KulfGWHyehDvsbkuaswfgo3ntbS1sFBgaFYOKuKcP27pUP2tuVxly8WHKLfzZtfi
p72O0Ojo7AHopWCxC1rV5cTKut/Ieaf7M5q7gmMmpqZk4pEexEqVl8Nq8ifpY+EU
oAy619vYyNZgvfSGLx6Msc/eNuL3RiMe5sMLPmkd/2vGRkT6m1xUN8lVmF6aWp7T
DkYSTXwVOfuaFsY8bkRyWizJakXg5s7dGDe7eCSzSdu37xJ4HADgkUzNN/X73vPs
8RhNMfmx9OnDJGgJzgyB/0sGA3X5d5RjywvMktYL2Tlwm0E8V53seD814VuMcG7i
BUlueVZlKm5Lt6PrX4sWpj3GIcxkguI8f6RUuvQi7mhGr80xIy4NDiiFcIPkgMur
BKQmSO105696tCuTuiL3QXLtBf9t4bmhF5Z+3mZqMlpUI9y8ZT2264XfJIhqpbbr
qrA4t6J5gnpJplnEdQJo6wlafsYmBVC91Pge/sUaF9vRnxJeB4kVAqMJcCTXLpwH
z8LGe+jKt7OpHJEpXWxh5T+5wB95eYULhM6h4zrQuZ7uegNuCsIiiA6BW3n5LSMi
RLTbMLOvGBLgT6oALMoGSQ1SzOseyFdwjhju1pv48A7JsJdCttk37VI7sjUj8YF1
ygxM85tCRh1LhwrPKXQpDKgw4lL1VO3pXQzUnSvuCcLd29FrfnuE8584QKOKjpoA
18PZhGA8uboBhEFjmS7sqjYXd5heGxuk20JQm8Yrm1OU9DzMPWzjlz4uSpgicKqf
BHw0ONIOnO27UkUQIf5pmJC7gn6YxkFj/8f2h60Xp7N4BwE789Po38XB+9ITEJzy
8vc2HjARp9xDNrwC4fb3+UdJldttpus91OF+8/Z+lscnUPlBdo0+mK7Z0XXcyTqo
VYQd+c5BK1usrfQlekQ9YozM8ULmSUTqBikmKLbpEfTP5ep6xZtW1/KNj1fbPmWm
quBrBN4TLzhwfcAUiE4RAgGu1MqTKFc0WLcVA24LjV2fUX3wVBmzW/25ej/7I4Br
ZndXdijz/8vXvKS0MOR/bDX3sZWVPshjWwAm0Ee65kh2RXzD48tQeKAo/vPdBR7T
9ObvYOj4567m4ZNHWdAx60fsIm0UGr03qPofwfuJrLCdQo2UIYfS+keac3gGJTVQ
c/ktUTibiuA4ys6h1vHLewUmr4vaPcN95Qmh8x/UHDCau/DlJQUtEEdOvt86vvfi
y/mjijcCCT+5aGZzhDqG4vr6yEyLdFF3+1w6dMfXhp9dc5qpuG1GyOh4B0gp36t/
kBUdOlKHraYyP+TxTVFM0VslGWg0Bzvv7ExQ3G9A8+fSZBibSJzx/XDudPLq6JZF
vx41R0CLQPVxNvx7namOJ7kQOJpapEeMB6Mz/lLzcj4tcHN0NRVJU3HDU5AwPamG
q5mRvecDiqmvWk+TR9MFAI/I/MapwTRXHPadrxRFVGrLcWRoUI4UUEZBmbMH3lr3
70rCgS1jj12zbpXEEE2sRUnv6sqLszKW7vvrqfRcgRP+HZV603xXovJCHblX+k+/
3f1RwWLHgmXAsBbxqTHMjZANVjtY8KYUHc9duW9OFUHI9N+W4I7WmfSiz1y6TY+u
866BVz30KCCcC8bvuJWVC5LPF39JJNvslPGDA2j+BG0Jx0u39M2IL90zIxKUG4g1
qz5LAf7ZNIvHNfJqQSJ1CzIBo3WPF7Pc9uRuTVtQEhokmm7lX9pmdm5P4Y9CrwE7
Pl6w9BvFP2SSROo+UyejP3PbCQE18B0okfoXew/h+PA8WpF1k5JUUKdDbfnnrqmn
uM2cK0ukFhy6nR/OGPiF60E30Q8rnKO4NhNZHRhEdNp/3IJrTjc50/fQucxwY1Po
RhQ7WAVZSBJrYHS+YcdiL2/1ASy1r7gfMtnFrRlk+UAsOHUoGY6qKMB82OlB7OqO
3TDPs3LNs3MIGIPEdUY0s5pyegEzevOKM1MWlc1d/ppEwNtKr6YgoqDOTRMjZI9x
S2hPHoRL2fmCwjew55aZXcQFtSxMH+3E3o9BPDNHoZONcmBJWAz4/DgrmEQjyei6
8FAfGcT7KgGpNvmzexcKmLbUIJxbzizWV9N+T5lLOw/Sdtf0Sdze39IpuOYDUYBx
kbDU95PY1rED3wtxRm1Pw/WGw3hH3R4ObNTwSh5ZW5A8hBw7/fyN+Uc2dwE4Iikb
FLZ1jKp9NSlyZOUtBNMhLDnxYlI31CX4dGrH7d464kD2o6EUNwO35JqX3pL5Hrc7
2brHRdIzKDh8kMmka2tOtbm3t2kCKuF25BbH9x7oPs+m6/PwnPpPjXMlDtg3Szwk
C45Pf2j8dqI/FCFj9YyjppnMoo2z6GIauVikNjJbee2jeBENoFfJpJCsAcE8xd8H
QY5NkV+jdXKiM8Ucnx58o9q1koVw/NWIHo5wZdlVM3aqq29WT5hBQC4GNdOMZHHb
C/8aICsv2CJCt/ceo+Np7Ja1bFi3BC+Y9+nOnYvvzxDllHnS/m2CxEu3/mneNZH4
vSgVCfgmZuInkcA5nPH0IUmuiDZmDluz/Ryssf23wCKCzcgUHLQU6ZRJTbu03UHS
aN5CBbN6hOe5DnW96Oo2RQQkobW5iHysxL6cheeHFxAIO8wHWr7PgFlYNF85bD1q
8tN2vOXiKepn8emxv03pFAO1sVZhVAD43jQJd/YPCagQ5enezzSUehimA8vvGXtV
EbAa+5/1E/GAheA3U3dwvY1YErCA8+CEw+Qjg8cYQbcTE/Ug1PYeBkxUo+QmPg5J
Exlg4bq4pA9jknWakCPPwZJwy9yyAUKYnEsxPhy0mzDnzWaZ1qp1M2o0qZ7VXAr+
FNayfSWoVHwpUhzDZ/1t1bMmvp2ZcJaW0PsiS6t1MHIxIr0aI0sTcibUk64dXlvE
Uo51b55+UnmQQT8mHFCOQaR8ZbzVVXkX1R1y0bqVy+3F0l2gs9NMHQ6nLnCCCvAO
RlhzhbkQOdcq9NWcaPQwdj2RBmaZ1aoqd8zS9TVh8+vyqiQHqCdaaD2wF++DJmFF
35AMyQEAxX8jkLatAwiTF1P1s4Yl4EzvPEzHoQFobaEde+Lkro2JkH7/u1kuZ5dt
HM6SadGAcqlmn4YkJhXFChxOUd1CWf3fT8j8i53YPM0yCPpy2WvBu1ajUwA+seI4
TPW9ZGHTgGTTJLXzPHEaYFL1sKEIHChZG5XTgaFW8Wn98LdTKTN2R3wu7645puq7
nIror+rOl5GF1Kz5CfF4soNkhwkc602bf3xGHKSRk+asTCfs0cR/c3y3X01GlAnH
cP0TE7zlFbxi2KcNdUYFw8EfICoDrdMhVn4bcfhxqKPl2KHiAv4gbdpwSRwjFiQo
VuSsfeLmSdYM3KAZIXGDkRKFZ8mRv7oT5jDibqMc1iZSX0zYsaNJfZY0OwRHQhBf
2OLvmGxKjOEVC4RtqpcICNbAAtqlcMlNUWr6I+XJXqJzCcTN+DQRx6at30VkG0nx
wPfQBfH3wEy/z2siFn2sefCOI3Q8VdZLe6CK2W3PG9lmOgZdKv8t+XhQBIG6Gkmm
cVdE9kZzXmYLCJLTKYMvK4K8rZlF9Jz0QfpU/RaEF61YA8cNMAVlYpFDpDLAiyWb
Mz5aC8EQDl1urRCgihK8kcPWO81ZzA2B45Vswlx9g0u8/LMvrikaz1tRAFisesKV
KTB0XSOa1GqFdpXtadQCVz/G6savMQGnFk5wOafVs2r7xRXgSGwAERt7NL/8E2oP
XEssFZD5CDYJUWVFOKjBq5Dk+kuh+GUAqXHcupH//z6kzUEJwisO9bV3I32cZ/Iv
KAlbh/qzChuEY9xm3zIEt2qGNyaJdrJDz5lv/AeIVqH1mRL+r2JOjcejBt98LtSD
yD9ssdwZSoZrfHx24XqWbQlR3x5maQunxo9ct25mwYnBCBrPMeb98alekcdsJCzm
kLSn63oO6FnAAqOuBDCJe+IEZ+WsvvFxub7aM/oYhxkJ9zxIbN1P75QTbaiA+XtL
ZjKn/mTTZEt/y3iMfmhcbU/OTMnJONis6fjB/5qyGNAHQJXQAW1xAfXvAAYamUTT
abts8sjP8Z75FLyOPGZq8ILQmY1AiTPiAAANSjSqwyab/bb9DjQAYjw72+qWcOxq
eiYQU7PNgfsAgspK0E7eYepRSscanKzXCBg33wPWuYCM3r2sb5YAtYB89wuaWX35
lPWaWqdmVIAd6wXoFok0VkVfrs2lqZ0AH5GhZuywgrAXc+LCgNicSzfP1Ll+pmTr
D10JPh3KMGSYx22S8bAmnqr7wnfO9ZZbr1jT6WELIRmamD+2NwmHTCOMr9kxFIGg
c07in3Vi2ge5WxFsY/lmu9rph07KtHkLavfwkkbwlRKPnkLqo4hnGvyh4LM3qlFK
HKGxaFGw048ee/xktnsVJgDV4kVhv6UJM3gfkXV8K71rQxj6U1kQ9ehy5EsaXq3a
IZH/m/HFnfsz1/KOA/wjbLtV++efmlr9R75cBVmg4dke19efdaoPZMa7YyNeD4a2
dELB2kXkC3zn4A4upzPeNywW6+ulCftuynlUkPCJw2zpKIw6yuZqUESgDq4nJTP3
b/nxNuU7IDv7rr00jlGX5JlMqFEFgPUzfJXDNHBtKSKjYfT3x6scu63vUjQbbVlO
zWP+RItFI10/MikYdGX3JwqMKdnCeVE7dOX+/Vwqomn9n5M6jOIUMDUMfnaVctkB
pwWuoEYThhhxIeZSWv5GdSsQsMs9hFbf6HFwGkfkzJyHKPqYhV0U4SZ27ZlTTEx9
WmAmdXMgoxWQ1ulHCfVkwA+avxLUJoY5x9dP7TnKwl8VrzNXMj03pvkONHrlVBAa
ayWJCwtlqwfOX+FsEHIiSHoluyO+kjPHcLos/tp6WzkWHWmzQGQ/wtDruFYHm3R+
taybtLeiMcoj0uQa+59jJx9dz4oa4U2ow7uIcPwB5QYVaNSS1PFnyxlCh4xFvfq4
TTYi0GgHDfVntfBItWpLmxSjR3AniuRGGdcbYMRPHoWwUANDI+Kc0GzmIixAv4RQ
pEy3FUlhwHCfm+cRrWqRBZ/s7UKY/JTj4KkzsRGQSe9yTRZ4+PJBCGwTpmCaDAWP
zT1E9zh4cZCAc6ps2EG2upyh4dkiaHSr2lzM53sOTg+1jVJuL/G2OpcioMIw5MTX
0zMB+5d2T1HbZS3a0t17DCD7KmzDA3SpMlHtrmK4UzadaT7DmAVibE2Ho5OJBwb/
oOsGZmUEFmpWrv9+DU/3VLB/8HackZ1kJsXV/bA23NiBXss2LP+RJju8N5D1ebjY
RQBEmci6CTYhDXyEfTDJH5Ixr1wrX2Hr9HF2VBsZUqKvNGOAPJ6jfHnObflqWuRc
LMNMtTXEUl2F9TDNDD5udcxYty7+bG8CgFlCj0J2McesyWpgtw9uFXSLDy/1SIKN
SS+pF30Mco8rGInk/CMyUW3B8GBXi2sQ0srej+8WMPBwrOhtg0LvIJxeOwa7xfpd
A3B26SmkcZ9K8J8MQ+cNbSjnbdYUhpT39gHRY/9LODn693XtbcZdKnFs5zik7Rkp
oXf+L9mE7Gx/vdmsE20dCDGDnJlt5z3l/8EC2qxXYZumISxFG3EnoptuliiSvyVb
f9anRB8/04vwfH1uIsAA6ADJQFgAdMF8KbkgRhnsaivhgv72iafZxv8W7MxMLPBr
x7xrZmqc8uJGqO7uk0CeMHiB6Zqv4j/d1Bd0tYllLJg8Q8SG0bjt3yy8gLrVPmBe
211XtVBRS4Km6ZMOF/CWQhOln0hX3+yp7HAxmAvSi9MNQ8u82rIhRZiEJu6/7K+f
HEgJ80973bzvU9wCRMQumibLrx3WJEhvQz891i8QBuh7pmejjYJlEyeF5+GKza2h
kJ2sLyl8VQT3K7KCwrOVcc5LBdS2qANtB7Us//SSH+BBtkzpgExN3f2SYKKOPqW2
p7XeozsWsDEaB14vg5/ujvSFKV8zHD6r6FAv1Xjbrvu9sm89rsFOvrsVHEdcmLiJ
64qVniMn12rb+f1TUeAZ/yKNQ0q48YptClNEFAzBanVGM1xKWtfYUDX1Tx0v8PH2
LJ2Y0hLHff5G8vimw78y0O6vJlureKGXjUyuaM/B6Z/k3oU+LEmKL7khtO4IlPym
GUWFhRLDf48fIg2RusuyYk9NktTgr9Hai8G8NExi1IlbjHbs5bKa99uanqhXfPlW
nzR0zNDLaPUPcJJ0gYs2y9sR+FSodlK7Q0lxJR1JXaz/hcTZOrukRc5//hOqeAuH
RZSTnOWp1bKOg6+9tsTrQwOEv0iedwP6dpnocFh94T+atvNFWQ9y4fJtLEjoZyh3
cglfNyHE721aLUrJiJy9NQqNYywyTCnvrhczMU06HEG6P8uyYcoaLzp09jhWgO1L
AifoA4J5UhWUlA2Imenemq1ua7M1EWXwmI35pEGSW9svMMaphQRNUDuyhVZhSxkt
TAOiM+q8ldOfYNE45ECV4LalGhGbcyMkxsVYtHPVLaFll1c/AKmzk75IbF7ZIqDO
W+ZVAdWvmCVXRFHIsQJatb2hXvpDtLS8/1Ph9va0EeC1vavl4pnUBlyOqAa/JrZs
NHpBcYx5hKQNr57fRaE4z0zmbhswT4eY2po9nutImfGxbs/TkbbQxQ9Yi0mnj4uc
x0WQFtaa3KGihb0+dJff1/TbJdO1V3HU92j33e83N0QZLR6Lq3MZiM/R39x2WNVW
ced1dkqfdmB68ztSXZ7gWmLnKmWonYLBwXwE1N+cAgc0s+wxj+nKhgq9e3uaZnPc
G/erMd8OdZYPiGVDhpF35Gr5yT+CBq9BNPjlvdIAa23hylKn5sNO8wosv1WXgYUo
HOgp3mWA+ZaFwfOCW6aZbd2rbzBQ4PsAZjoaJuttWkkkqLlFAZllp7B7z9e1JmzM
3rRozCObT5UY7BJDXsr4UsVPzRY+Tye7to+RcI44aYztNt9cVplxgIqDmGd+hVNs
CA/TjPrQ6++/MMkETrwHuJFle/q7E7PaKoeOGKxSIGxmR4AW8KSNqLBbY0egkR/n
lgm/D2bCz2ySfwkFf9knFlqICjCqUq5wV8rDh5uBI2sDf5fPVKfAt2kcQT1q6kh8
dybiFfzRvIJkXBRFy3BbR6ewmNiuDQi7m+16PTgwTxmdaxvqqSPSLeHtJSzbPntE
0F/gjXO2EkjxNmVKmBdFYJTJeIBWsid4WIB8w07Ys9FCDchQnQY6l8oYWe/qZzUE
pzrHuXlvCnpgrqR9rO8rJhoqLWWsJds8YMvjx8RXoVz8OVoyvYEM+DLIhCqrgEsm
vFp1Ge9Dbx4HaO362pgQAwHP9W0OsDdDb205nmnF9fr/9mn8nhnJQXSlhyC9/Lay
QaA6EK3SDEnWw7CuGLY9ZDX/ldQg37KaF7BJB4nOBs8rsE38CzKmZaen7lgNs8aj
BFOwf5OqqBdjQgjjePy3KZT7XoqY6IPdETuV7RG5HuWCqiYIWYuc0pMFfMrynnN6
Elmi6Kq26Avw1/wcZCDgAmQ38izCml0WqtUOSsdPYkDwQaYSypHIpNeqqDjqcDER
6NfjowH90vOsYVgVcLUSJDn/aVqiKcMPw4pqbeXTulq798VCxCL0+AnlLgMEmnDO
A4q80gS0/pXyvT1O3D2LteZ6samhyfaZapx3OmkWOjlAM11b5rbTuOiRfWIeTEdb
tBzDnFuFbgK6hh2TUANn5fy1bzmsV8GnPWOqKxgJru4d5jwM7xJ0hQj2csBBnahZ
D/jONvrX7r3Nktgp3ntPYBY49eZ+/mS3JGU+eQT9c635dglFSxwfmyWpxh1Tu4XW
sjWDzX7L2It0wwTwkbdc5nT3ew/NgRh0GDP2LO2qdAfyHSM+iu3Tpc2xNPHCFgsm
p6VIXmrIL2ALkwUV+npYjcKXYuQ9yhv3fs0A2bfMvR0clemc1S59bnZlKOEU/gy0
7lTQxZeAauP7nJYmF33akZK3Lxd5xqpTt4sWPpQ+2w8kkZzZBf863fOBBdVvE9Fd
sg4ARqMs+LrvPwahR+KrceiG+mOkziN5B+WGTEbRcJGDwsyT83AMXQrgKCXRDsro
jbKjou65mgTEMC5xSgwcTkzsfe8maddDaByVYAm5ig0DyCUvNlr5O2D4UEWjUhcN
UVNf7BHxE6VMPo5eFA0WMawEQJXxmotRNnaxZZaKqKPABZw8LxY9Vf2SnJ4m0uSY
DbupNbrgOiI47oq+JFSK+BJKf42BHy5X7XP9A8wtCX53dGEap2TV/XedrV0JSIgo
aL7O6OODMxMzcRbNDakwdJvEGJ5TrHcSyTd47YDu8NLJUSh0gPs86lsHnbLJmZ2F
hQPtBpCYr+tmKTKNt2sNoeiKHCMyKJnqqq//gjcZNWvIjWL2CXvvoWq2aHrSsjSC
tm3/doJaFJRxUT7iHTmBjUAFkkz+auwtAs8/xiJrwzGTEkaWEdy744pjslOrySy4
vvnMBM0kF5QtHNw2fDvzACFCMvwrFD0MzgxVCG3fBMTqLHzYGQ9zBVW5xVoHDBfY
BCtLD6dOouT/mbw1B11cGLbydHWp59aeEMM2xIzVyjLF+8mwjf8Yu8VGBztIP/6f
6NFFgBB+RnD7PpIrOYQ+Uwxb7LWWalVtoE5OSs8tJ0Tca2AgxYdHfvJkX35AvHVD
H9og+uD0Jbh4Mq+/3M2BVPc6l8elaJ7oMwtQ9DL/J5jTK1yArSZiZ2DzulgJdLFl
uDhZR0igL1FAxs0vMyW5XQ47+H04/VUQ6hSZLH1cz15g3y/5Q0zMt0XEN7FmjDiv
+5TCan0cIAqsYYUgvaYT9RIudldr1jjIEc346GrDygWItlw2OLP7gSzDAGXRWMIq
2sCwyf9XgMWq5igHP+Ul4l5C3jnRvI+Nt8suhe46O4Gx3lFdzRAJ9tGDoiw3q+qQ
/0P32x4vCCoFyqmix/YVopp4EUVjF181+AgOb5TkpQeaqZr6ikl9HVSubwjkDeLl
aFNRmPD20DF6sfiVjDtGaq4cRuz/fpwOrzCL224zFBNs6+yap3XnE7dtSR/PBJM/
tbC/sb1PtNclKFbe6g6ByAvJiMJM0xI9gNVi+LtEYFbrIqhQ90MCv5dbg7RWK7j7
f/+mt6Ai/YdXaT75DDP/agzqXl9hqkGE870Oz6AoIllhgXkjnOzjz4khXB24r3ha
5rzjwPUONYvoHgcGa4u2G09Ah/Oj4VCpx6W9q0VDuAW82MRkvl49JFI79UV12QEk
ILYNOK+FKZYMxaTEL7It1dljhl+by2Izduuv+6dXDT5/CRlB6TbRgf7vGK0/eUFk
ncCNLzLBt5lQwuqFHX6//7omdwDTSOONtMAvcRiTL76r3jJbMxPrDceXGh+rUw2I
/HrCo8FIzFh5L+CHITECVB0k/qn7x3Y9dv0+OlfAts37bEhTvynDHvs30EONIzCv
JCtxIAV0/qzGIPkfA5U5nk198ndWoWCZbWMQGaz5bk8zEK/437FGrxUsV0jt0ZOZ
WJOvLH/3yKrWSlSVGnZhO8/ZiVig4V3UqGbmPsyBcklaFAQjeMh23wceUXBuSauB
2LKvMT+Jah+dWAdz4XB6THp+Qc2b28rwYKQQ+4k6z8V1PvJekLAQB+glHxEmZWEs
fqMqsSVFN74iHOdtx7rrCPdtQv8FIs3FNTi33TrCS0XV/CVRyj+8bycEMy3ahHKR
RwbBsU6yRtI47oebmVmC9Htj00BUzyPFUwhYlsm85CK0BuDlsDoUyoIk4yvqLSOO
DONFudAh3e0bl/PrJRrBhRvQHGdnCtDzqU9a4eN9ctViZhJ5eVymeErAwUC3Bny3
mxOUv3faU5OIJ/n3Yw/FrC+4r8fFLfjlr4sO4ws+4j1K8Zaj29KmdD/tBCyy7ei/
1m0jApwP0LagiYVj776TQCTPbjFiAlJ/T509WSLW23JutZ5pSwUM0MhrxoEJ3EHC
g/do3mUF1hLDAvZyoMwWERkuIZbjYPXTXEhJMMTWVoY0zJWOJTrPT8xUGvoaWIf0
Cm+CAdvCUCbhF6QtG/2ggEJXSYNjLVHNG7pFf0iwK+uHXGxzNsflNZH++6TAFN5S
o3MwinwUKFrswn/dYFI6vbbv5wAIcNv5VzvC1sAPmkyBhLYsSitpit/evCRrKcwo
+uvxY2g2pTFU731y1MNVNilRSd4nUEVkctL09zYhxst1Rb1DBATam7Yf0X9z2mXu
CFMEGgc2d2krmpHaluF5ygUmtElEmBRF/G8oiZnZf8NX6usbt/0wTpZWOfh87a1r
dRlHK/aa2DzyyTxkQItL8shNr+UCGwyZJ6V/ewkqNb1bRP61V3jj/HVMUiknXk9d
CXAEIjSuMDnfC3E3GDVdti7z9dSEpnbiIFw8TdspIk3sdWsDLYBVq6JXFh7tQapk
FgGjft6K5gudsDmPUoM3ir4V/dz8+hwqovSh78oWukHd/gSpy7wPh4OB9PDZGI0r
Z77OEo9gjFHOAT2YitQKQvLKDVv7BSvsHcF/Ki86NwR8OYmnRsJUO2sqoG/kCcUH
04XYjNWOwLVKtZQ4xAlcXUJykTAQJIVRBsAOzxt9MHl5HgV5OYNTenmdf8HhJL2s
vm0oKAEP5t9fwsdbQC5WNLjYRNVaiSjmnmCkmnsZATvg8/z64V/lYfcn3x0Uex4U
XQbbeQ4ZRBX29Wcr54el6Uz1ag1sJN9DSiYG8zKQxWhGLR8aSjlwTWcPlgKLC2xv
YLEAlDx6Em6+GXGrqXY4EgP1CxnEfQkILHDxe/ngi7UTPWVVh6NtKWaz6HJDtY5h
aGGEuEb0Djv2Vc9T1Uubq0M/CoxNj1VP2EgmeAxF5Mnh7E6QxvMOykGjho+FdMKe
Fx8pSn6ydLf5spIqSpff3nWTFlpSUo1tHJ6ZcW2s5Xub9HM7FXwGNwC9iHUadhYH
82B5tmj9WRWAKv9LI3v9tJPKPJE7+Vx5B6EpQYtqARu4PYKzLeuljflYIX5xDdVx
4iqLYcraHAlEeCvwvhTbGBsoi5CkUABBxssn2kV1L94Pojopn6O/qavq3ewi/SQj
Gse8/S8Q880ZoGLoqrPwUaVSsLJkoGNokCa6LAt6d8G8nva13dE+YCRSluxBIV+4
imOoK8mP3owpWjYtpaGv/buIQZzZGITzjgI7weIxw1wrWTc5mNBcU2IzAY5+I33m
Pyfy7+c9qfuPV4XnDGhDU4VQ1YpOExcf3I8h0hOeDsXet7TS7BoWVhqTksnOanSg
ZNCjUoR8A3C2oJYeUNvMBsw7j1Xz8kaQAhtIXYPtYMLkfsbo9wRigSpKqp+FEfs9
xX6c7bTH2tXkfOisOFT+of/bgliGKXhMnCxkg5+Tw/VNKlhA7uh1yc2pCwi1q89J
CXXQFmHQjmsXjujLrXvjlTBjIuXTS/vfJnbVbh+572Er2z/t57ALz5cQWLxneH5C
+XJbAyBrvBgVF6JRC9TFkeJ0gXss6SvubgBJPg0rZwlj26OulQeh3lT2OwbLKE9v
+Lz3XshK5W29YWaKBQ283n/WxNuZXXZEvGs17HEByuXZ+/fg1RZ0NjBTBe3KMORq
aI/fJTBEJXbmh9wYskHiZqo7Fywsk0lvDEl24fqQU8RER/sNhRZIdkswRdtcQYP8
czwDdK3mpX7b9r44cNZEl2axE3lBmbldGABj+L0sFkWutacd8GwrVGTD9AHGsx7x
8FtOQ/4agsJgj+Dvt2ZKB6rO+SAhQ7GL6VI9uaTNP8i7qT06/pGYDrR1M08LvZ5N
mW4avCV6yMWRl8RDyXAIsFa5OxM2lfW0n+on3nybVzYKCVAqqgZdZYGYEM1+/Fel
AIsNQyBwdRCqedU+ppySeYQ5srPl27Pr8tXyGj8L9g6P9e+Ti3BrUFuAqHuFyiiU
I6JIUKoHn5/uAzZbJ+bGr5ltYqalcXt7G9vXHedvFdTRQLOrzkvOIwzcCFUbnrv9
U+XQ/g4Jid0Sa8r/DSv8aC2mgRY0dONk0ZrQ5ganQCp/7glmx3vd52hkmofbJs6T
bm//jAIWmk5Ss8PCB4slHGAHPoI9+eXAzZWl8c7Nb7gIZZtRU+DhjwGdlgPDFbA9
PJAoa4hsujdVbwJ0DzvRYHqGAsHER50bH5BtrQAbuVzI3UqCEPXA5FhMIqQo4Pob
+xSj6k8cLF87pRH63Hk6oZEseq9V6yxJ2WbbcvX3myRD7kZW4Ahth8Kp1T2ZCYo6
uk8kS6qMKpKItsyNl/iwMd5PX4+lWyGKe7A/X7eiuesve1cddaC5LO14FDJSZoHx
aInUXjNpnmHnt0hCeZknwEF6JpGMkTb8TwP8ggus9VzKbVQNXEC+3jA5aO4bAJxD
NxwunwvKiB1r4bpCqmt/AssxGBmL5F0STqanfJve1Zahk+ZZGUfV0FZpCAMEYVhq
jivhJGzrtm7sEuBNI5DAAeFajTofA8U2bRHb5aKFIUchNRFxoxPcfVlzBdl0yQ/L
9rONVBKJ//3MT6pZibibqT8WCVD/m52x4K3+aoRtotGBDzDsx0DXTzZaaqDOps3/
YMcJCRLsqsmQ6jgrX6xtn6ccQ3gqmTsRCrqyXhojKT2+Ch5j9ySMhk0w3w0r+yMe
tcugtxVCmP0TXE9f6GMLuqykA6lxs6BM3lO/O6tISznu85VxhCdN1QejVBtjf2Ou
sSw91Sp+bdT9erAQyPzsaHA2Ljj3ov7gPD8c0jArRKr3ehQlo8wM6wEwWBdGv31f
ziMuCV4vpap7D37Y3THwtCZSppy5IE4kgsQwpJ+4aC/r9XEUOG8VUfGAC9/jvbmD
lj8eIDCIU7t0JeyhIRSjgU4/tmOYLbvrb8M+LPLveoPJTDRrQA//UNfpLX8CAPwt
GHiLZNXa0ySfH6zpFFgBnASSdaUHavxc04ZZ2DGqfC3VHWrPCZDrPqPv40gdaNOW
olF7aMcKrbRF4m1psNuPKCxLNQr8oWqK1Ffd1xkhi9Bbgpqb/5tbZpTIDmnPn/lo
7fcmmxSAxmpwyRn+tRTCGXw2qKwrEHvQfS0eUtyAEfbxjQhHSPVT+CnOCN0ouEcE
GnkjCZatkNUYW/yXVfzbYuyu/FAIOWtOSP2cQowr6mFEWhzV72JQDvk1n28Ablze
7Rtbx/QE3Girq76Jthtxgxhi444HO/MndxtNJsi/flQTKEPxpPVB6DErqZiRhNAM
8GjuUEjygc0vmoIYgma5xzXlyZC4giSl6GpI1jm+cp9QS9NnTd/r6VJaCdR1E60k
wedhWOQryL8dJjnjn3niLTcC5iN7VBWuI4laSz6Ve5A8jWiQnuXsChnzlReUiVPQ
glww4L6etuMIVuzXB6ciTpwgv05BNhqGeloUwP8h3WNQcdhCvnsy379Lw4JRse5j
+AQj1r9spPFY/AOcfHf/rTlbdDfgsXldObtSyFcs289ZJ0uzDdN5uKECNef0l4eF
UwY63snpzNkLipiHTJWtGjPviKXlDJGvRkBgDOa7NsGdnCmwzMRh7a8EunG1yxSO
DUaoTfX5KYjy7HdeIxdlGxhb+oWwfZni35sUYU2xZvEezc3TfZYMR9hu2xDI1B9W
uV5QVEJdkL2mrl3BWnFky/ABn6HcmriuiGogKDxUNw/zgoTLs0QB6f1fIp1xNdWK
9fH/kEjx/r1xctk6Queeu24lnR8l6w74mjBs+JkynJF/S0Dc/wFc6aGow6JhZDSN
KcdjjlVJFzJHoYC3wZk6Pn1KDCq7c+rvyhjoXwnCBJo1OZI0qP232Eixy1tQJkS+
TdBqbdKpIZFIEyZ6gwOb5krAXM8Yb1T+23BAMyIlaIgX4pW7wirVszI1Sc4z2B7s
ezEDrr+V2YCDV7uQ9f1JoznxHLTcSPk6/hyM/T/J2FZ1XAxX0pcg+rKSuLJucRJw
tZJlhVxWL5K1at8VSHImi/yxSu4k/4OpJYitcR8AAxvXcWwLHzcZxph+ED4ignsJ
NFZfdFdYf3Rp1/Y/ifHplDZAEste3uF8d9PK+mDkbFWv1JToeaOOhXMLANwc4vLD
79fcK5kllmobLfAQyr36+HR+UhQ0urh4WWjb7vdpJk6K5dLG0DVi17Okeuc5tU+C
qwtBufTLV3YKWjo8PvFdkGXeFRSlfFPngvBUunvqu2LQ4tyocxUwtmm0A2C7UyOk
DyTqDXeP4dZR7KbraDUokMElyPO2b2tXDDLnvVdBb74c/wfO6jUwXBtAgmGCMOpn
8d9lo73QZbpNj881ahLe5ATkDcvW4EsPsNcao/r19wlvWaCCGi3Zl1pIlWfpHyvK
Ajv5VIsKGn+nJM9C/7+dd429DhQMEkaQrWuMEuxN/Hvme8IVP2midlIrfITV6bcI
ZXp6ifa6sI1UC6u4ArVAeXJykZK7CS2E4QPxrw9LfhR/f15XB7Hfeu/UFAAobB96
Kn1kaaiVjiODGATHwKCTw0HTCkKSFoAnX3XbLsOgajVfo3lavp+hWztAqpAE9Rjr
x8lzo2oxhi90Yhqsd6otdP7zLF9LjsBnXjPLiIiwIVAM8hsEE6xPUXSX1vi4zMCt
DheDKbY1nTm8uTLLCaZA2WARyehteWMOCTzeqoUIK89wRdPEGyWZA9dyFmfUlgEr
FnaJtOlxm2a+Igd1JWOzB62AWzcuwnw4lEhDlcLFdPXQFiCfJfUZN5fBXpvba8eX
ONHwCaIrhJHvlVfaBNX7dcG4IyI8DX7YXvc6y5qfhkDwdOV3wBhBNVspnrQjP6PI
BkLU03f4EZf4TR5BJzMD40HgbC2jVF0S7VVlKXUpxDXSwuEuJyLCDWvnQafoyo5F
OLJj4tL1R32nOfN+CL/tNn8lzTzs/a7XCQG/q+hL92WfAccZdK9YzAzaUE9o+tJz
PPftdNJRerCNtexT+eynMMn+OH+altP8f+g6qatQNPZZVUptR1FAGVN2mobxFozl
2idl18IWD6EHr113GaZ3vWOH4Tbw8U+zJaT1HOZ1u6OHqG7N2ir+z3E1wj1K8sOI
/D07uQeW8fD6/ahoLIeQpBK0WtaMuudi4kWM78hVsPPXyRasFFdTGW/n+ujPbelv
oXtOw5KCZpp7ErOaRiBMpO2gfyoAWpi3qcIJe4z2VTRMX6FOaTQYTNE+cM9pA4u8
jSEmtp4q95OgXXzBaL+wtSdT6+6F0X8lG9TdfIp8oB0Ef8PUsQddmJ0D8Ib5DrdV
gi8zfJ+mcFMn3ZfyQjJFX6D9/O2RA3HUjvlRWWC6X3qOaChAeRBkZIr0RuQx/96Q
mvBLRj9LnGq/lmKXmzGByj4l66NCJ1Vqa+1vDSnjypYq5pdL2jJLH1ErJk8YzXhR
D095733nES7oryC9gUl/5thJyedueOGCJKYTX6tWq8TCsFP6zKAfk0nDt9sw1F3M
4jz3yqc7dM+wCL0DFbKBkw0Ehc2Sk32eZ6krAjAHxwdNQjX6odK+6qcCxgqqfSOc
zO/WpsUosXOeU82PfaaMR0aSegrluWxD5sfUuNUZ8xQ=
`protect END_PROTECTED
