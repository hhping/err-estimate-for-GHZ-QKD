`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwOPRKbr/2G/DzfTVIn0LFwr0j7Q0YiX8t5UQthnDzwyKjgD407UObalnqS50nEd
JPyCCybS4SXn4Qq6b1HJFyaBUN3J4LM+nSoViH+P/T1njctXkcBoVrm0jPOpWHAu
Oy+pyTRPFWEF24AqKxcE8w4qVoKeaZ6UPuL1zdanYv5vQNsbCeg+DVwO2XksVyTH
UnDfm7dXjalfSmCunBOAjCvdTTsdWL4CyYheU5T4SbqSRTXGBP7YTdpgpXGa3z+D
C+JOnKEHz1kgvvkK5uLcktVf8WK9rZ6oO4d96pg4QgRvrxrnYY8gnujBxJp8F9Ag
Cks7/ug9emoAB+lbCLfhhIx7NkOANc7E7OsRb5r2ez3fZE/UhWMvoIuUjKzICvLO
Axs9dxUoAyXYjAYJpLSw9lk9fy/FeoGjdLXeMMQCDTMtDr9EGe080DqtBtZSy6eR
xExhuMkVChi1Vku9RBZLlMkMaZfIS/hhx29XsOzTU3qQ7jiFF/taPMHOqogvWcSg
J5Kx80oP2EFTxQvruPcsq8f9nTFmBfi7NsHXYrGyXfkIGVWt5Egiw0ufVYLYLf2S
TrM4ht7qSMpkGQ8J8S1kUo48/1TT/bGWwYi4rzl0gp4kiWJ3efCPIdEkg7jZQXNY
L76RRvEpT0aCoXVN3cm6HGKmahoGabNaS1SCHCdCuE4/6tcAn7UnOUsGMr7ttnrI
dr8qQZHhPBZOGL2ycsiDPj9ZgjZ09pcUoZcNQPv1rHVYiISb8NOMjuHr6pf46SQa
9b3pvqELCieouO5TBAZbIg==
`protect END_PROTECTED
