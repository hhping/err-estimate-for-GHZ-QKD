`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LyLkqdZXpj92e726ddlEnGLJCuifOplYJRphgqx+g4nZP2lEbY4Ux+qFgKJSkA3D
loHl8Q8cKeJ1HQNUbHp3jH3QOt/K5ynu0sWFwd1M+/fGh9r1vCOu+PA6dL2Rtifp
oQbP8esTr2TFxtz+yImbn1feYf0armyFEU+7MvulJ0wAG2r/6DV9xMPovE3N/XEB
vp8S1DXqsEo54N3z07ptA6UCf2L5Yg8uoYLAptRSTZbPaODFi7BGHJjMgHtpW7X8
HWBrsjPhYYNW+QZyqrSZyJvnKlp6lDAnAHAR7KV2CisIGkz0tUP9oUBwE1xsFpWO
HCjxn3Z6Hww4eR+JKmujaQutiMtSty7hte9Ub+17IWwSK8Fx6ZNiKuAXtGzyZeYU
JB66UU9zr0lCDNJ5UQ8FAXWG/dnX6LNK4x1ixoTlyHNbMgWsRWWB8SXb6+7Eq13Q
2gcbfAMmKBwYa7UkeGFTXie0VmrZf9Uj8XWu6dqTZ89rhfARXviDLdDqJ7c/CPHo
Njxa3Kocb+athMxq87Jbd4orpJZmXvV4yC62jocnKULKU9Q9e9YySVu/8tORPPtY
U8stZsGgrkFHvYcEB2S2wPVdBaHeQLwYcvRjZ0fqlkOBLh9RodejUTSE13jV896t
w9i8o008L5qYsmWkpMlMXfEoWLIfMrK4sAbxpWvQjhmgjfXG1WHqEKpybhQi6Jal
gp9CDMIAlvCb1Y9nPTnOOQ==
`protect END_PROTECTED
