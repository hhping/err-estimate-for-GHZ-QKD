`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQsNa74t4wT+fUSIf67JrMZ9PnOOdW4a7SohsseOw9sn2mG4+feFzIImaB6/axHR
uMBtHi+2kBrmxvOgTSWRgPb2GwWs4smPQu9+0il2e2Ne/bym5td5W4zCyBV+9Mko
AxEmzeh7jkD3p3NpIXP6VU7T72K0CrcCza+f52R7KMZVp0/AIk+79sfM/YNUdSz1
B84FQdhFu9Tiv6uIN9Slpd+orzphPiJuE3b59geKeJW5CT41/3gAk7G7dQda+nvB
jSAxlIiPot+6TGZ7k9PGaKGEdjUv9UTSfWcjhH/txzGyJ8Eh9fhMhurWf/JTaxPn
/6QWy/jelHv4ciPSdqDP3yDmMcaH9pzcEcXmYmEnDoUELhmSHlXVNDvNVmAADj8b
IdYmIgEb2BK9NZ3HGguGaHRulMPompirUqfONJ02SrXqsX0Ml2D1vZT5qAWkaDw+
Dxw79IfqZb1kI7I4wYAFyDmQrXkRM7tdgJH/uU5ZSL1Ctis2yKxAite7fcSKtUMj
0/K2LOonlsQNc6ZQMENGTxzb3s1hkV+PiwGZ9ktZTJgVMqdz5UI+pub1vlAwgFjB
V6+cDIpunsDUvON5UZmfSc4dVskOKqrZVewbIA/zGqIoLHxvB5NKfV5b+susPPbh
enZbVWrL8GhdOMWi1tx5iU/sCOC9fBNs8xg//tOVeMisoHyt7dCqDgQ+BC4rh1Vg
uPZlYW3DOoRkWDV1u/J2kapW0jGLmxK5la+YxK2tvw+EPt2Y0ut6ddqSXexhmRRM
35Z+UGdohnIPaZqDNLHsQHWA9DpUKjs3ELV9sqxpAbx07LNAo3MYhU+OfCcKZVFM
50OCsqz+e0U4RmlBv6llslz+LNyKrWo3JtPDdX1JOdV4n9ipd0qnwBpO8WCC7xb7
pCVWqT9vfhKPdvWIwIe8CEO/TtNZXk1PYgX/DxtjRb5ABCIs6voyflYOvYnArs9w
CwoKOm2T5qsfL35H1UT9+0/7WxsSD0HstDH4XmtBwxZMySpmCZlogJoYNp/RsS0E
KiF8C+igU0mXJbv5kycDbA==
`protect END_PROTECTED
