`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KVMj2Kl36cXz0vsOie73msfjZjfY/x5vbeTnShZljd7axBs3yqiBxHL9IdwKUedZ
x5sYWEXS1M+/56HwaIGCy5HvXNRDFcF0RGCId7n02FvVN76m/yeGkIjP6a7SicF9
Vv11TbrrACp453j+Nj69zyBiJRLblgLv8x6W4oR8JWEKeWiJo4fTcErQP0BkCOHN
muutG9Tkie54K6w0VWZb0SPAO8EQMa/+ra00AO0TCyCbazzuYIjXXmLtxFkU0SXC
DGeWqIvX5dPo9fRoLjWpkOkPCfWVxKLDkuvmfqgJE3xySrcNGR8ug4DpQWuWpJ4P
AX1flU0lFzcTNw5o9Q1erPZUfG7FuO+fWiCjTkYX5i2yNiZPO6EJTd0WHUHO50zJ
kHcUf6pMN8G24BuHazERtivgbtldrv9rH8b0hLKsdZWgoT3q/uz8kgAjLv3NL9k0
3QxiRKN0lqGuifCfySTs9barGzogkDUGSJTHd78yQLv0+YRCrNzsWRav0Z0dFYCW
n2QTkCMeL8zDRzE8FD7AZnSBhe83MnI6iu6UnSXjxw/8GAfQBysuWzx+gFdM8owM
/Tv7fYENLnVMGmtHqTpr32W2j1PuAugRvj10p/nC3PMV1Uj4t7pjfgOGwmiZlN0e
dkmAZ2VZ5GCxwxGvxtvP4hi6z3gKAypTqeh/4Z86UDNyd1m9JErg0W0aHoEoOuy3
OT0AfVGx06pCCyhA5zu6yAIL6BxEmRnzxpXsguy5bf/z/x+zlc5SnvctrSiA2hgV
onTWGVsKPKGyCU06vwEsKiM3zZW4iIljzeVp9VIq2cYsIJzUvs3gXygrw+6fOoCC
Bl/+LyU+xTIK24zvtAlDvS3H7Uc8N5GX1f12sJy1iGjkh6X+H0M3AAi6SOMl1DMS
bYIJL2TixiNgH8HT7Nm89/hQXfXNfsL/RXeBboTZI+T0HbeSNzTuYd1tgHf3IxGh
BFygPHOoo2O6F7rfUC7qMqBDIB46JNbKreeyYthcWkrwLDKrRbOey6SUWj3ImivS
tgP4faGJPfa7q5qDms5RfxFekHgpbnnBg/7ONHvNvqYXl32jLXDJTx3Q72uJVN6G
UwNaQZt7YokDHuDt+DUZlVOIAUTRGBr17LaloWOxnL2vEMgpyo0wYyYsIKtm7xAa
HNuMvrZOV7++7I1uxVcYJx/j08iB5JNHejmcAERfJDdgdOX/p9uabHGsmXii3ARr
MPFlv71+a90i7xNNcGXSlSrbZjHB/OxRJ7g1LvJe7h32Qkvy5MlRd7ZHZvr3H4md
I5WWevw13irlHIvV0v6hTnvkKk9uEQLI9nlzkaGX+ppY7zD79Bihh2IHU8jqfeRz
MMesh46mftAqmbUJHo9c9GFxOKmApQKg4JEvVz/Jf4ZPJAA9oh0FQ7VE3NgQ7YqH
x714TptaUBIG66K6CIN5hhaDpRI7BwaSl77qFQ3s//JtEQG6DEzMx5AATHGWX6As
pZZfIec39Yvlu1JOLk6cB0Ew0eQsQz5LI+YptOIxLJiByHd5CcgQFrSPW17/2HST
bjDl0X//qNyWAqnwpJylnHWWVI3KkPRonoyyGBTfdynmWtGXUgv+1MJxp4mO0llu
yrbX1Cm2akDM/xkl+C6l+XquyibPfGgDWzDoaczWnrkOU62FSgP2/x/nwVYMReNp
N5krT+DqinrnLdSMr2RMGwKRnziK9i3rewwmOX2dKmrdF0O8rz9D8ywI7ABS+0/w
biefCOGg/2/AV/YyEjLcPpms+CmAKRbqYbVhD9pd2wesWDBI9ZuXgaJKK/wCXArd
LXVF8or4ueWXnlH63j5sQQVBB25jCCvzmie9xRbWmzG1C+RuqfCqM7YCYSMPPLoJ
sEh+IP2gz/TxPCvtA3lOAiJthoL+d84Td7Y3kRPagsiFWW57MLNR8SCZzqYdZQO1
a8PbXpEWaBJOuyT+/hmtgsArZKcDkbYoR8g6/p3u7D3W2UXtU5Jz8xe5K5POVCnQ
voXBPNhXkLuchs3aZdTmrg7WuRX0LuzYLd9T9DEKMr7iBCXYYz0jdFzyPYgX1MOA
sNfcpSpuyJExbuw6lqKGRtcfnOdaOp/U6JprwRrn2W8RRdmQG25OS1UnRm+Wyk6a
dCGcASdZ7HJzeGQqPFujlg==
`protect END_PROTECTED
