`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LLUob147QRqUUJU6bbGG7ODQmBRV5yy/kASLCL/b422I579sHz30eVHtYZgPaMuH
roriWhkBKS8PqcGrLXoiPgn5qACVy9rIub7VaYeilHzWBYmxELjDd5FSxSl+anBp
57nj98S9tgyLpElIyqDJmcF8yaARS6glBZ+L+zzAD+hcw5nCHdcnb0FJG1HJA9Xv
A6KogRtDxQ5Bo3QkbBoY+b7bhrp/7AN0ReRJIvfmiXOJi0fDJJ4kbn2bQxy0lNeg
1/MAFTCxXBvwYKV7+dOIQmdQprbPRzEESfiyJpJbEQZcjw/gmIBNvkz+Y8yxuo8t
cs9OKYO/ySl4M85DwzTsVxZv0YiO7CpvOcQl66FqtQ8/zghmUNXOUi5tgRg6Au7i
PDSVTiG/uZqDmXsba4bfEXi1W82Z2hahbjLyW96qmA/DQyMxgsVBwn8UYO69DJf9
bfppyQzP9GvAQG2DiMxyrK7bDMFhQeFANEPSzuLGDQMGkbWkloBjNDzVRagaqJK/
uvssVx5jCCjjfa2BCU+a5zDjugxrO2SxnaSVQ8zyG3ySiFe5ebDd2pWCKT+2C88B
tkz31vuAX/VdBJrUvjpOpx1YMiVwG+QO9x4bDdXT6lG+bk1oEwD8GMSG9J4j9XOC
uBc7/nYZDHKVAQBnb9E2aOig39snDLhCnX2NT5m58zKgEVviCNuEDfW1IEv241v2
uwcIb8PnvlEUPf4D0yhVxL1mzE/1dGsrNAuNToL4SN+hDTbFQrIBMpDJP7iP47vJ
WOvJKbXTiO0ltR/vvS9Hv+BLk/ieWkGtCqdUtLQUuY4U8s7CdJ4IJwboLmtmHN+o
kQ1pEtAibpTRPyngKFdW5tG6kcS6iA6l4rFC7MAVCeuqcU136vA2GaFdM444uNdo
5jvAg9B1ziQWqLkIM3DRxzPWJBnYkJCkjUeal2xQpzp2uizbL6qpQpV6+qpjGSY4
omkniV71z2iVzQBc9hKp+NmAPIb2gKEiOxahKVw+/vgU8XHW8LaBa2howRpMMPS9
GNIbS8zqM47m4bjidmBCC8juAJkS8I/Ro2H8VgRnbU1ULMPFnr6Vkuimklewrvee
hBExICHRPNSpzWAlekCHv/p0snVBiS8jf3sMpv582vVz9HJMvGGf82eoEWmBHNA8
ebkYEOeAiFAIJUBwMhoEszjnIccuwiRB9rboC9O/RrKAWUdivTLDvu5yfz5JF9Rx
8G5Cs3OH9l/06vvoHMGv3uNpOVrroiPI2pPrOfCsw9g3Xc+qZx48jWqmi027hviZ
B3PtdwfNHrF1+LKhHUo3MRcLJF0bEDQHMszgXog6+8ivpGAguhpc7QllGGNtZvAq
daQSDwwC8aju0fIPNqpCVOAqv+5GKKBIe6XtkmrYY37gVb3qnUyRabFMh8msKDYo
EfZ+TNeHsPdeb6DF4p2pKtJ8Auqv8gSZMbtR/davt6rnB1AIq61vUBuJ4eCO0XIk
l9E+pEW62yX9ySJNEzJkxi/1LH204h5tDjeN3fQ4LGbTpGMtWb5/3FNgRPlZ7HxD
5wCnc79A10LNZrLxG6Kf4ltiktMQxuDPdLeqM6oO/FMMflyxlpTEBtve9EFnZPHP
Ut0XI3zryhcK7skpJKqjNT95tDKKdUDzt+sReA54JqXSt7wBAorUWzeSNHwW227A
3U3LWUbZBRCcjP4+T8Q6FI299qna53Ag7SmqwbHCOWDmh3yMm1LQJlgJmhnO3mlM
jEu0ifLnPrkaNiADDAErBasL2A1/Ziq8gTuEjPz6wW1VJkQHndqyyofZ5PuGrrXM
rjMoyAyC0r+Fib0MtQ4VHsmhbKJNUupraF3JL/NPUGjTV6CWT5c94Bdc3VG2IoJA
riEKA5NxZWxxQ0TT/trCm8k0KVBPwOWbEEAGfKeviDJwElJks0i4eiWNcP7tyhnT
5KHckze4G9zXxbLRpQDMe5d0RgKiqabmVqQzOgst9kdX8c0wM+R16hWAWlMF72iS
KNkw3xCInxcPFfUBGjXVm3BQFpURuxczG/aFOayRLdKdkfXWFqtNwKNdgXGelw9o
xVaWkpjZoCVHTnhf8kZVL8svgS6fOk9ffE8FTnd1+n0aj8HGZVsafCr5NxXo9dl2
W7r0/BEQprtx6b28hq5WtOcz6QVnMp3k0PnpKWWoe+VxjmjWnmn4bzPFoAQO4X3A
v7YAxpHb7AUytDiOrgBblSEnguLe4nHgEjtnWkg9XuXTwA6x9w2cHdzccFPzQl/Y
qz/mlXfGyvD4sPkCdb10lutN/5CwVuoYYz4LS/qhr8H9p6HPBuY0NqcO3FxHr3uk
+pV3YTQPGLdv/7ShQ134+KhpuqAL6lT2T9WXGqyhtF1/C327Grt6F5Y93RQYogAZ
+ufOSDoo7X9ZMN80BepJ7mLIOiOqN2wsPwjGhFrdh8udoQ8zxACPDWp9e2bxu4mF
ZUKwvxAZVImgbvH/UGjqrJXzbq2+AZ0VkUkcByqgx4HWmrMGnldX2SvnvVcbSJuS
eFAPcz2hUS/nr0pjm5sRn5VXG5+8pCAiDvPALGT5/wz849N3ZKKGhTQumCgPx+wS
jueOkEYNoJPAwuDuIebLs+AXRrPfyYpL7qkVKoIdMLskPK+xaq6t9ADUIqJJVXs4
M1qNAsjzAa4QaoK4XFxfl2My9s//XavKeQD/8Z9DTWGF1nE28A9c7mcYDQZowgpv
VABUGM1C8MlyCQ89bpSeULOoJMOQXMh0ytnZFucSAp4OAlSiCUaFCZf760+i0xBk
KhXPZVHvoh+yO4roDnmglX8aQsJjawxHm/2jyIRBMIOYiTJll3CWaz3bRa9NWHqj
bdkoA+PySrXE0SQ8sWDrhm40gJ1Oxs5zrZQ9cXeYf4DBHksksarqHZK5qZtZ4kR5
aSK7OVmKXfBPOdyTC36J2Mcbh8ceaTJLAMhBOXa/xrOTwTVNNmf0ZglJCE9P6jTA
379EFtLMTS/2B7emT5vF9lj7yVzSfUpCIbFCfqyuEMcJ6xv6mCq9CHyLw0XCpCjd
747yScD5FclK4YXl5TX8EKf3vpvwOYwSMnFXmsuaVBcl8Nuw0bUlydfSGXLkBKj3
eaZzjknrmO1DkunczXB4Iv03jGcC62Rj5FdJKuVQfIKC5jiTZ/KOm1+3ZGkwlITS
uhzOiv7xOBBB14vzcAce2+5lej7dZ4858+eSVUBusESBeCa61e/MU7Bb7ZG05iIY
uPlmcpMLpQuMarZQe6VyucK5NkwTWOG+Vur4zZrDQZBUunfnFlOxMBaeKCjrpzSq
BcMzU7ItKeC9zSwVGte8VSU06PSm1uVBUfcX5DUCNyBbYrMk/5K7ijXmMj2hr8ZK
PsUP7kFTWAIrllQkQkMsK380Lx4h619uaByo6lMWQG3+J3yDiQjuLQrvOe+ojLnG
yWwD9NqYn8QItJZvWcD+w1l3V4XBaOd9vqmiiviDZq23G9oMUqCWXDR958nrYtHL
tsOsvig5KEmFsW+CM65yxsWnbWIoQj6YDjvuMC1/qrdn55kyDck4h/hVk5pqUlSp
Lps5M/pcy+zqG9fv9994xaWTPdtasD6ig1MfGkqDeEL6EyHXZ2FtgH4jK+BwIQXS
CihZomiwKGa65CJ8oR9mo4y0hlvTLy/wUc3/M8rA9AFxdz6u0ghIWwH2Ff2Ol9/d
O4GfPViWo9qUxTJP1kcDxGJmNRFlpYiXVvq8WCGdHuI7M3GmQ0xMAN+Q1d5gcobh
mfmsVRGglUCyMejVbUfaoXQ6dAq4qNwozJglSDcdGMvBoHvEKke40qa06oHe2p1M
B4XoUUZucZwb1yjuOCcKVyBWEMWObA0xlhA0lg+SMVojypsblQREhx4ZULpHzzxG
1olhiShJU6dHzJ5RDm2xRO+WeixJTSv+lSFm+0wYMA26ebq488UPnmTUZX3CUFYB
9YnA21UIR7dev29QmTSr1jDUWXeIIqWnrlhqN/J3HLViFb+9VTgITk5D12tQtmkG
Y5jx0BLXftQoMASrKL1R/Hh+0J4poJ04TRrb2+gUmNowH3JwJROhc2AZEpGoZMjX
Ysaojdj8SD1ppl+Dj8kODbTj1U47xZG4ZS0X6xtj5SOBHH2j7r48Fntsz5oixT3O
hmFLJxEG8ZqJYJeW6nifSi+yrHpuOE1PURdoBKI/emcyIPOFZyiwJWnE+0nG+6As
Ub35WZeUFPnNvpAVoC7MyalNhRtKwE+/jhdJWEpimocyraWY3w6wbzE6ld/FsEhh
RUVsW9dFj53bdxTB85sTJa8x9u5PoAoks3GgUXBt+5uvmelBPjqIoZzkX5f9MQ4v
DVsK2DsREByHzxgHy/hw+uQVM6rJDPobQ5hEHxZSsqewLnuJFlDYKMgWjnxm0y5M
3Au+wU3VscEf0PPypzKJlEk/HOasdVykkaUdSBkpT96OTsR+etmbvunCiv2GD61E
NdFoUmTSlcYOJnkRz4N6tMF8+VIHckdFHF+ZDQUmmG0N+jM+zljcMJG0B3X+AkP4
hEVO3rUUDxGfkiWDIQgRSmY4tspq2c1w9ReU2qADegs53r2y5mdqWVT6w8Ocea6d
Leywre0fDM7YAad4vYPYN3o02OwRsOqQTjpJgZQmbLOiIjx52Cbt9gG7c8FMpz4m
B6hqonD2qryUJKhIjcaYt7sPKaTJooq/LLCpLEfuNuJ5iGNJfsJUfw5exhxiwU2g
KifHxOkIk5jQEc05dkQXNB3282DP02CM9QVba6Mjuz6/0GE1fezVp87h99oaJmkd
INC82inm3Bw8Y4Bs9+5tIesbWqy6iuqO/F/l1FjXYBU72HcecIqrjwLyhvFNStEu
yXQOMIrsjkHeRB5qLNyqNLWK8Vk4Lqa3bclHISaBD0RtaY4KFZ2uLjJDECSh6JQ4
mPxrxVHQDSrRCCHPfHIf+MVg0X4SArB0Uxh+EOjIkW0Y3IT/bQdclFQchdi734Of
caMMvSTRJQ0WeuyvfcgdLPkz8KA0iL2Y44q1hNsPHwbUCRLgHxOIrMb4pfDPCPv+
aE+M7s5OSPrizEJ8XDup20buWObk7GkcWd8TH+IJVlVlNX+CfzI358VREiMWpdA6
sqdbN3Yc4hM2s4MeptjQwvR47G3Eq2FTPjJH+9Q+ekj4RriKcXMnBQY2uujwL8iK
RJ1/TId9rZItbd7mCAb4xLRPwsrfugHHIPMFmIjVPpC/JCOTRNrBhT934xv9jzSq
vvAd2ofhsUhitcKSI3frDg==
`protect END_PROTECTED
