`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fpmnc2Atxly1N53dPpOGIbxWMUxbGSMZ5LOYCiQK+K9WYE0QX0bCAaS5PkPnWVjk
rsm1C5HAkY4n+NKj4kCszBmXWDVIdminv3T4pCnF9pUcwiLYk8lDGUaRCli2/oDj
KG0KbSiOwWbfICs5XBa2sHTEiWXz4YbCcMz1NpbKXhhc2DB3AvrFtpubsLHmr1jh
gezZM4G99KQVdhsTt6FTOrk/hisSpHOxMiip5mrEnDxfzokEhbZkvRpZv7IqT8lD
mXHLWrPQdldlEq5wGe/cbuZA7iJTTiOXNVqOmHMMn59kHumUe4NI2Bwa1BwY+sVc
sXZeiUOD/Mt/1M0410i6cIs4TKyATEYR2eoMFEsC1XBwq4bCTlFT6wZKR6FhoasD
0tLIzlnjkKp4s6LfFyF1lUgN4/2ZxUH/zmx9HZicNSye/lePlFC8Dlzpvr88nFAk
lpr7d+Aqi8deLV8u1r0R5YzeSUj0Jqo4f1YlaujKnBzV4kFwqcmGFA++by/f/9N+
`protect END_PROTECTED
