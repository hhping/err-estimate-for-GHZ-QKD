`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4kYp4FfxK/hlqmz4wTO7fpbACNwLjgrBJEmb+TRp11Xbqs0evfGgORVyKWbYBL1j
nwLrTeRKp0ICj14LrB5+J1b2d7cZXIvSCBjdJaYCYG2HuQT2cfTNuVofP4QNShFv
x3DGz2y3I+Ey8xZqKgfvg1mr0eoZsdVuAcf8xw5XgpnkHOhcPLnKmDlxNZj/wsJ1
4DbuNkDinJEW8gwvMxaKqQV/7rSAgjGZi6SPVBhHfFmka9MEzDSiT96Ti/E+MFIY
4iuNa9YpYOM2gDczAEgotyXq+piRnCj3Gyo6/vwjWLH1M0CYjaQ/oCRO5zP5/k07
jUw21hm+a9UCAp82kQLTqKGlYcPpNYQ1pA8Gpcs2fngwXzOSmaMZ8jgsx4uOtI/A
qi5BPSC/A5mUDWE/dLj2j6wRl1YsdsC216oTGibFpzZ0Sqt+MjF9+SILO3PNqJ96
u+hqUkrmK0W8B65aaUAicg==
`protect END_PROTECTED
