`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JlaM35qCTbhDaATmA1C76dPEvg+9FggurmUw+tTPDE9BlUXuCuRnq+RyxITkGrNy
eNv0eP1VRHDsyrJA7oe2moTjqZ828X2iW5HVRzbcvZ8lftp5bS0paiqfIEB3HG+l
gneKWgN/Zov95jMOQhkXCoLUYX+19yeiBcMf0HuaBkP5NxMdERh8cbL1mPBkZD21
cVwmpykkwYUtvZi00A1qlgh8vzCEvXtz0LxsEA3EzK6e3Ep80AOOhwkwVAsAPE7e
YOxeq4cgeped1j3PPvYJYPD2Ejtg08TIe9oCd6mvxbn7sIzupuS6TDgF10WrneHH
TnVaU+tmXtFqRsXgzK44cqZz+sLg9T7wiLYZWpHX2pFlGd/S6ypaXajJPioJeq6L
NivyJ53gCJlFohKNeWZg914erRGREVNkolnV5ySql2KZwBszbYXZUq4dL97tborK
nJHYB7JbIa/4ghJHZEZdLWparhRTkgFseRvrSRmJ10F2sOAwI0S9v4WdB9eCQuh9
bhtVNoqGO/zkQyTbsgHHre/MDUV/u7iFzqX7AM6y/GXga/lJIUudxOM7vg903xm0
fQSJ84qFMLLDTmZAx08qBAdwBmCfCXFDv/kjw5ObZ86gMPo9Jyw3h7j3qDf8W6vR
ob2y+XG7MuxRv/vqcd8E2O0q4rdHhWg0jgd7kC0+8T57FrAELMwqXhlUNDNHs0oS
Xi3Wem/kdAfCFEkyIk7BXvh4wA0+V+iBSKu7QpPjq+Yjq0AWeEZXN42nt/xRlmd1
78LuA5tClqLHeo0Ih6W3QY4PQBONsJDvjzG29bsDbjIYYVxZ1md6nODU14FaksWd
9LMa1j+w8/YJGS3TyjdQFNMfW9crJBuSv6clq5+5akFFr1YjUyX+E3I7LuyI4Aqh
yuqEpGkLXiI4ry7n5RDzRKLCtSkfzKbLfgubdXAEwbo8paXB8Kkksql+9E/QSZ7a
lKUjY2cIMrDp1V7ucW4YWW2KtvfPdi71+VqlIaebt+0tPU+LH8d6NkfEv3b55Mj4
bpb/wJ0A62t3gfqwhAiy4L5bb1bDvYGzGUhh3VumkTZZpZcwoH+ZNd0h78gF+QFe
5SFQNY7BBEGpOTrS+dxawPM3AIHrziK7dt+T0a2Dv2BZzQofhOOlmpEgO4OSgSg4
u3se4KKE4SOpupjI5KUPQe+jdeKAFo7XETo/TWyvc92I2oSaMzZsOXbfrNK8XoYG
OqaliDR20hZqTUtfXSaIduZeQ8mqBefRWD8ROYEIxysXKsZzlUgmwHXHS1rkupZD
h/pMXPoYi6jtvH/S+dTEXUZnMJyEbqhgqHzMTAAKjmRemuHJSNa/kI0MDKWYFF5C
r41NI5ElfY2EqTMijoc+t1b8z//Efwi1mDy+AyXd0rzSNr05s8d2MbaDLzZftJUq
MqdtmTobpJSxlPlgJJYW8hG2sbCgj56m+67y+5spqnGC6qIMAHKjisCeG+sTTKPJ
sZJOiMF07V3rf2lJ10q0Wqneu9bL16KBAg29wYCSuhGzVXPRvWTQAPQqZ2lkQbAU
d14o8F/TaCmXI0V4WgiHtHVqk4EMjEJ3a2LcLvkaknWzgmG2FbDv6k+957hFKgX2
xQr0IK4Qq2P00aD6qF1L8mPkV8sbVm1Hp7+et+w6bPGL1EJol5NyJkjERRGj7MNu
gNeB4YfaSO92f4OW9f6NcOGIPoQNNN7iLgO0Oup/j6LZuW5eNtWBd2WcCV1Yw7ZC
w+LLDN3I1YZbNrZgEWVHWHyWFJ1hKkcrx++hAKBmj+oEm31nSoZX0Lj4v7Rv/cjC
x25+zelnuaXHUsCGKdAHnA==
`protect END_PROTECTED
