`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3y1EMQzNJmO5R3u23eWvFgpnozVdq4xyyz/4r3MVuojhaw1hNfNoLKzHHfAYpGe8
BaANXe3eKnJfb3bCMMMr6/CNuw4Nn+sQU6YbVhKd5tL4svp2aVBW9QyNOpIMbOYy
X9n6YK+p3mDKCsjWN9lf96eHeHvx4aJH97MpXhcwCkYRgrl4fAgGZlONTeYp3LUx
Jj9nE5ShxX9edYiZ4Ik6uuJGdE5PTgNPm+h5GMUs8ImOcIksL63MFtuJ0u8mVQUQ
QiQ3OqA3L9dI0+l88BvdZWTtPI3yDw8JDeLg2FDLTmv6WA42yum4HnlnSgS8N+yP
76SEYZ1/7LyYja3bsDaJOT4xJkT+YgGJ3CxJ1vrkbxHoFlTOy8G//i9a4JisCrsX
2J0wWrB2QMOFWeU2pIJQ1DNXBjNqLWqnyZzgz1H4vgtDuae1ZopDbxzfTMFQuAd5
QaBECUds2V2rcMz4tzaYyPqf1KzTZkT8xkn/+MUYUnalWO9gp9Dsdx94ismzxcqt
Gdbb3Jiecwav1nshu6iqlw11SOr7SWVnnr3K31Tb7Nc2HY7TnKnMJgjyjRAnJHEo
lkeGgenmCo6Cgsxf3rnrtrq6Yo3keUif4JCEANn/JcKe8ouJB+NWjGGP67o0xwHR
McL1b6ISihuNAr78eIroacFI8qRf88OjUQqM5o1FW8rIIpIwSJveXNsxlqrAZS3W
j5ERuS37+dPpmLrV726dK5oDIVkfVpwX312Hqg3rZCOC++7zQdAEOJ9CZeZdIeyV
02RQVw6/SKuEiiJkxodJcRz83RGoq2ncvIG+o3lhnHc=
`protect END_PROTECTED
