`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vmiXGYnbLk9nL7B6Sm36rWfWznl0Z2V7a0GBQW706Fwd4zfORYdecGosJhllDDDM
FT4px5tlCZedWS0vf/sISR5F3iHOrsLnZp0TxK84e7/nXIvWciBzI8zyl7r/vpQ0
xR56mqM8oKThUwYf0VfJpTIEcIbfI5Uc5tE4H5T7Utc0oHhgXWx8LE2gr6ZRM9Ir
gpwbc7+4OoJXCmqLSkIyslHjbC7IzZqsdun4bZ0kD4YDNbDejg3bLa4QW3KHfktd
bVujzs26xJdfzuEniDv+kHFsCogXAt9jVn3cDOfjoj6zVLQbL6GfUKOYy1GeDl8e
K9+/JkiLfn+yssI4cfSEPIPfQBnHCNwqo7r0XgujJn6DItBMxtI2eMZ2YOAgIB0t
uw5VCsuzTrQTBro6iHppKIsHoaf98NUs3zZoBYC48gKNhUarIABYbuviWxNGWQzk
c8Gu4UaWDuB6x0Oi7hS48jawQ4nbXnx9CIeJLu3lQUTgIuEN68FqeF0jKBqZ3tbZ
jVxyeqbv3SXNKL1IigEThYlQplYzvjNExsg9Ywd2SouL3k8RA5V25m2VRCWsYSCu
CoX0RBFcKUVnmhxFpKksnYuDS1Jns4cRvTCDedFtVa72Nn9YJvI+tJh7Kyyws9Rd
2793sN5vkX6xRh955z8JjTbW1asB5abIWGsjwVTy28wwaKQj1YCmXYD0TdMJiWyU
FyGGuA5sFq92TwP2gd+84oWJeB3rKQz0G9FYCvA4a0MFn8TDklpjg59pgQW+Wwoo
5RHgfN6Zf5csj+t5DBzC3Q==
`protect END_PROTECTED
