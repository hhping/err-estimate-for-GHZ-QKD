`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tiLyNvfmAKNJzcsrZbqFDTDRY3WAIQfcgNsSiTUOrzjWDQAhlOqTaHafKjp5xs2C
QB1XvGs+9z3Jt1yJdjsEEb8UobkE9Kd9JuBN5X6m2bHKhyBrbSG3X5z+pgnkSxaB
cb1HrEe3UaL0szBCPLFtBNbxTOK1r3nSZRiplPHSpMqrKPMfD3jy5pomBSdPaRYg
zeBjE5a40U+0WyDxbZtzG5KzllHnj7d2FPFTv6UuuGSqKcDnl2IIMtj8y3kCjSKy
NLpSU5WE/PQE8rPMGo70rdviu7lIsuxOWt8RkdfsR0/tWVf8UCkv3UyEvYYPIHGG
RK83789LFCrwSwgfRAcvjeRgacJWEBt9axMl/4cMeAvdzHC09jjhFC6hg7RiBx2/
g4LXPzQMINmISZBSE9Xo/QV0Rwi+NSoclwhEkDTaXEbsKXrPujRArf6USQJNDLXv
e79NLp1vp1PPP9gsO1i9wOqFqS64kLRyIgEkQmAbPFK/SgnlUilR5MzLG/R7RVS6
ScqqqN9o2EUNLc+zcY/N3znLxlEGM1EaybmUaBtFs7IE1FouyanN4JtWhxWHq6gd
sQFpwOmCKgYtmn2EvDn1kR2lrz1W0eU1FwGbi7fJfg4okmLUs6DMfQWrDfW8MLX4
DXWRPgtdiZ0y52qs0V8I675Fuj07IB4ybJTNhpyyRRXdU8ND6pV6dsTakJGAyHME
8Izv0MIygF90mRz/r5wN3ZQqKZpJv9e2kmnqaVMvlh/Dts0TbwK61f6XBBrNdC8E
7rdbT99oucHXoOWdweoOtA0ySDzDAXk3Bhf+OVHK8i/pF9FFonfmbS0cp7Xq7JXO
WEqf8vwC6z9GGZM/5mnMjnAhn0AIKLQrfob/ZWZglqoG4YaLu0IKmZglmqJaif+y
OVo6qupsIrOv8oWAFt3G+0W7fSLjKQxvfOABjkwGgvzpUFxgCjmmfL/aazd4ooo4
S62qcmlBlRScbR1JrBdg0JshcdQJMCzhhEX19HkoDwy2IVhclapCudJ6m4lXLGoR
DIULLDNVTiNraqC965u+E6XxkEezIZPqA+DFAQ7D9dMO93RDoNlh1A8Mr46sh4fc
4iK0FLeZSL42sMwM1uNzn2/FEsixVviQHbzTEao/hzCuLssWGUhL40i10jl+yXnz
grvTS0ahpP5x+BwhuyjsS0ngVuEbJadYQ4ae8l6JPColyuHnJXUnLgm9BuA6o6LE
UFPuvJl6MWfoey52R7W8kmYm8GcP2d7Z/JAHsToAVIVwUPK8fd2DtVh1SDqu/ca9
h9FhOE0Epf741zvt+cGLkB2w/KDV9oVMaI8iXFDQWkg1aQyE/6Fx4CVMR0iaeRrV
bNf8W+VRPWbLzzc3PbHvxXExqdVDr4YbzlhsYXI2fQMODLgdv7HcYoBLpkgM64PT
h8hQjzU+r7fY+uL0Omw3jJn+49jzAWzPmyArIPOseKGniL2kqlUyJfiQgJAJc46L
4hOnj2LtVXI/q/d0V+bcq3sTgXdPguh4X6XSd9tfZa01I8afWGhF7KqYz06q+bq9
XqLNduIlTaU7f1WHgAgMzTuU5HDYULvCOWtfHKRQGJHX6ZqpuvGToav9yY2O4vEI
xVte81uI49hjINt6OWUOlS7tknXeeS3CHV93ht+YoZ1118n9D8MkZ0P/MnXk4TkG
DBIX8F+FwFdAuMF/RkHTo5ze3xUfmS6zNSzAguiAs3WTH+uk9Br9O5n2Gg7IFuYu
eLBnsJRqljx66DhFmFL5ApSEcqxeDIHpQdDwHBFyfcElJsknHqm/Oui2clOLCS2a
ai0vQxuJyIjU0wAABL3TX1X4qjOA49+fTOT6pJKc7JYDehmANrxbIQBrWkwolEMe
VLzPjSZA291gEdbj3VNaRPJNT7FgBa7xpmRgOGKxRpwGp4T7qo4oH98ywLE7PMIp
I/rcEjPhl+rKtAhidLoYgEn2RSfCucIP2Yug+oL3++53ilsoH9T5/BNctBOyTuS3
YDH3nVZXwEEcChqmdqJJuot93XpPIGJnPJsyjSlwPmIwz1u+cSS3yBzhot+iVj77
EOIt9cCtz3dmvEazHl5jLZX/messM6t1naPhie49s57LQVgRFqWvdd5k7NW1mEmC
ZSSZIbf48eIxcRW4YeGzbqz9mRgiwnG1PlCs1g0fn0K86+17qYCayCfA9BTmO8dX
mGrTGYsfhNsbpSyFDU2gs0hNgpbEMSqm5RF4lS94sv4bE+c9ZNWV9hivc7hWh6Hh
juk+q2hCJVvnqrvExa9Wae7opTzAJo/kUIu5c2FdBK9yEIFe2xf3hXUXL7pUUQkF
cHnZMabEuDjdGgqWXR3ouVKy+cYK22AICVvdboS92eJL56WTVwOZc64ayr7/NMgJ
Sxkvw29HUUakaCZFsfOggac5vAbVMwGICV/VF00XZZT0ISbsUzXD+0VsFTCIn32r
lGCmZL2XjBr/TDwTgxneJWAcL0z4B3+0aRqP7bqMGZDGE4W/r4QhXwCBOxTJ5oEM
MVsowJqtIn76Tyog8nc/J7ONCImMIy0kpm98cpdaMsGC04SqVSZbRHg9SvNCT2nI
Ix5FOAWAWNLacZCxGnZ8RJtpiXMsxfnbDBAd51jSWV8E+BuHo22lyATRJ4sBMBfT
DR3GFz69klYoj+elm7rKEJNVbXMzwS7XoNJ9NIzrjaTg5+pTFMOqeHgkCcpo5Km/
ZPS2YbzLv9jy7fbCs7ZmaQ==
`protect END_PROTECTED
