`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJrLXHu/epT+9KIUP00xgzyotGoMIhlZ8W4+VeOaD9yrGEBFPWPHNu+HV1fLfXlA
UapAz0AU04C6g/hdP1gl+4h/MIA8B9cdfKvpqr1MHKgK/OlBtoZiTlAI/Qdq0zEn
VW7TsQeJXQBVSTPyS4QdMDw+GkO9ZuxMqGIaVu1/EMwoT56duJUQoqrrCZZjwhIR
rmAjV/9NKIIPNWqgyaj2o5trrimIrLEI66iA8dJAD+qP1EJowabwgLRnu6iXTVES
0vOe9DnxWiaCE7JC7iW4B1H5Ja3Y1IkTW6nNidtp9Si7DoXOj1TN9ArCeNHxbYQk
hStR6ukl+QtBaqr2hXoXGh+r0GLLiErMU2uTGxdfDolGwfWRHEgVZcA5MUvv4+lR
fQGev/T/XhexUBsFpRZPJCZ+YYE+Yau9KsKxO8kDE56K05OhSoYT0bUb4NA7io/q
1/dLjsPugyZsYNcL+fpNHunJJkaAjGz1XUdtXjTJvCXMah2QGoz58rJGEEboiucV
s7eFqe8aUDTx0AOZu5ctUw==
`protect END_PROTECTED
