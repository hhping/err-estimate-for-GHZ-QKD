`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vH5KRQcWfE/ImH/KlLT+5dBMCRTA8fIL2d6nPnCL9SaiCmHSathQUjg3svc0LyRy
7wPYYcI1CtoQFurb6iXIG2OEsLvfbVSNypjKm38vpa55H2n46Bjs10OKnb1sMQfi
IuSoisIKAyk8x+Wp9/f0O+i2eXaPOQnBzKeOhCzxqP+yp4u6ecCDj0jx39m56Amv
b2BbBdCsAdjeUgKY6aAN8vyntQz0Nl+xFpPAT8PmneYfruoHv4shbNGwbvyQg8x9
0X/fPHzNednAz4skQz87uDTnvUVntbkrs3QSbYBCsKfHNY1bTipPRfkmFfhfdTRg
oH3skkK3RhR8/cju18epqRWsA0pmBJoelLSPUeG0Dpi0jWmwwOqjMkj4ieJdxAhn
5/vHhlPTkPfF+QiZRzqmVkr+m6YFp78fyC0qriE0xDt9hbKx92TmBXqTWxlfYuoO
P6RPlstzZo2bH6oigTBS8Xdsv9Cdd5zpATPnv3UlcknQOdZvnmDp9D4mUIYoY7JV
/A/HeHfka2oKn/hulGf2oq+NaATT1xH8s0bPw9c2JnLgYT5f+0XNmRXhNimIeM/k
aRIV42rjpfGVLWsWtrEuU23dIjZMMEi69cxJkv+kEeSYDc+OAlvCQUqbAgL+jWgQ
ICMjmSmCl2/DWr2/Nm3k4NgH/JjA4YBHDgZEw+je+vSJ4w6KlT+QHkndwxIsRy4t
78+SHIdUd8yQ0VyK1zMAmhPYF8EruLAf9s98Qcipr1hYOnQVuKVgxxzwQaSceTGk
Ed8qiD70NAZrghILH68nFShH0ICYr5S3xogcP0AO87009EK3ENgZ2wvtQuybMFjV
CqIiKot4y2sIAPQZUmi7wnfS+bxQR3JMB3ARVS1n+i298SpDt6IdSJ8nwl/w3LO8
oYhYyR1wlD+3oJvwWgqoCyIDCWOH68wF+SZr9za9JQK2sTXeoQeeYSAj5RgEV+0R
unbaA0k/ZKFjiLM1dO4JOVJp/P2dXKUsPPo16wGukeTVEjH2Ozy6Gk0+DawbOMzo
TwAeQfSqjAwC+ey/VTn3Kw==
`protect END_PROTECTED
