`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6aL+JAv9MFwakZQNcYPrjCir5AYsc8nr8tEt5vc1vuYpimJH2qWLJacnVleVlGJ3
1cegT+PAzBDFZAJYWHtgdbCRYb7jNgOCriNjF3TbJY11Yuv8TS2N8aigdlObANrP
ucaKJibI/xw4/Bluy5YTxgr+5jndvA8fTxy1uacbYwtlfYcqgDHCEeeojJ/WIQjl
WTDx9lJdsndad1SikChZTCq53qZJtT1gXZuteURU/Dkcs4vWlxu18xiUMfIbewgj
8V1zNTaX17YEH1c6xl5r0Pr4kfmuucXIotksv8tL+k+frVSqHEJhelPETdkuK8pr
KRSQRYchkobcdtQuSzK2IUGA22iYvas5/N9EwX8MpOYE/xGgfN4/jkILIRYNOl2s
mtU+kNUJl9iuf7P3Sp005GTbAHZLYhVcySaw3WzGTIxNFwt6tk3SIsj7oV/mcdir
TViYf5473SaE+gW4I+NamtjaeAAzAVSil2vM8VLlm4BX8/lSDjv7pU6oDjGhTI3Q
rZtlyGYyBs3HnUIc06KP9QFF9vb0vWd7gqJocLssLFBxmAS8RWAR10iDO9OslAjf
g8P4E3U9sle/CxdpnkWcluasEL2PZyGoKIqM5cj36/kZzKW8ho3cnGRHIou/TY4Z
iBq4yxSOE0yzn+ONtGcB0e93VTAaINcG7oH8d8gyIIbtFNBR0zTCEibp0tIwpsJg
27RppvvX8f+kAvUvRJ77tUW1NuO8xcPALsQ61xncB8YUzL9WJqvMU1UxV+A3uSdG
Hgbjrn/IocAzc7jJ5m60Awj6ftPmb4zoBslabFSb0Nq0OL8mVxuYclkxq134wI1X
UcTZcB9teIkgIybCLMVXio0fY5JU4rIvK+jrVB0P7c/HEtJmQqdBs7b96hkO3Py4
taVIM3yFrBEWdBD2dodaSmdbrRqN5J0WZu2rvw2+ERRXQG8EzTMjmmYLQSDtgB56
5ksf0wkybrxDV/GiholdPxY9KsLkOIbIKngacAzxqIZy440A0qvE929Aq4FhpIjR
m9BbyMQY1h2Agu/XgETjMRyDZ6cNH4CPiH32Mpqd+518scZGD+OXjU0tvjmeF4J8
OCNpEJsvI2djvJjFsq1cOG55iMDANidjMSxsIf/zFS5RzSBIG6emKTd1Q5L0+isP
DaG+4QMN+b8GXacRGDEQiBLaHjodr8jYrcxcuGwZCQ/VetYIz7nsPi7iWUteL9bI
XMy8UoP2KxIYDzFVvUPTU6A7aqKg6/bJO56+L22uZy0c6Pb7bGRfHB5xRzoCdsfF
aI9bXXNv8RsppJc+UZ7cdTSu2EHzAH8pOOyw6bxHZN0WFnZSD9efdG66HA2+5drj
uwyB2/auntjSCV/5//U5tnWn3LHOzoC+rHiXK8eqFxFJs/AfRTkSIjtKsWVtS13j
2dIil1NdIdBffRfFkBpUMMrVbNgkwGBbTa9RtFGk4FRzG9LS3eZp2w+Nt155dPOo
UZr0HcaCgMCu5z6zKmr1BZzOoSrXpmDMkdexyKmM9MSm2rp1X4rBGRzOJj1Y60OI
sz126DOZaxPGpic0GpY/qfmIJXRQS4gjJhRue7JRRW20hW7gL53FerPe9IUiF0jv
YpvGDUbDc+fTvSBYKKlogDTIjd5aHw9Vkntt/oleeUB1/jt8/sUZiBdpoXEdpMjJ
55yYZxVhA949DzKEpOi0k4FgdBaasStrct/G0i9fzkhVuiGxXwNuQy385uGBwxIV
fAp6MggxeDuq1kAsHKzJW6bj/q5Fmejeh1ejbp+bVkcmAz70djFwRBOhiBx+0W4h
I1wsvZGQghy2Yypsbsk4gqxm4NUvjxDLcWZhrZKyk/27ATK6CxVXcI7B5iJhvKli
b3XKKr1dsG+mZlJw9scG0uLMtMlF6cZZoeXyrqqxkTxgOHedQwwAJOzuiKJJU8jj
NhnxQmzNJWq2lqzsoY/Tsv8cCjViE7utlBSIeOhft3EbXDAc5GuCAwcfVfuz6HdV
21GNh7hytJxasqtiud4EQVo5teYvpmQytxVp6VikWsDXfZdYALjoN5JS3QCOEFF5
zHhJgHRGHwf+zIMsgeNpb4WSOGQOIw5PGGwlQFqWrgVOZ3zTG45fjC00WuAv9xei
Qq9x42ROk7fzsEUWSAwEv+M0Rdq9jhzDIyHne1y6c6MkCnbN0A2RHnIWwZg+8DZF
3fyN5me2wtZTsehv2xLdBYlAJJ4flRuH7iBESnhEMfIaSMyS+fHkZMxHFH/gaHGf
xY3e4OKe0LEbGJ/5OVpjCyGMHfudW2htLbzGKVGiN78mSsHd94rxe+6XWI2x7gQ7
+DiXInMLRFge58wnFujYQTw+nUB1ELwPa55Wl347QEecRUf7AS7yf6qCp9DcPKyE
aNcbFW88pUIF9gJ2GT0GDePFVECRfKQmxsG4D4sq8nE2MBhSn++8bfMrOeKd1SWl
9659OxcfnKPEmJ6mkBl8I8LuM3HPYDUiP4et76sVyOG8TzPmPyZzLuwDki4sLkSM
ZDqr3zrlkxcfRUZdBst46fDiRUl/2ZW4g7c9v4fNTyE=
`protect END_PROTECTED
