`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FH4LfroTxcVsgjwgw4PTT9PQzl+HxA51FyH/DIcx9LHQpbEGTjc4Fh/2YJAXyvSB
UHaOOeCPcIPHze5hqb1sYKq9+WfNjjjUUA6mig6hNPscePBj5fj40f9MJwYDcWix
A6Wd4pwmgw1H69LzatrKKMUQMr08QAX3Saell5EgQDrwSw3gWLjW8ia6VD4+ayaX
9yY+orSK9OqFnt/eu1UDD9GK7+OlbZdDfCTIIprnqPRXirCmHn9QO4g0WNaq+IbH
SY7yBNmr0MYgS+bA+G1kbo/jDQ0y/+mhqHVtyGOrbRceOZ2HPFeyP3nkWyL7pfSQ
OlI8RD71DfckfJUd4BW50DtZDvNYXuI19OJcBN464P4i37EyU/9LI+vsFiq2N43H
K8/a1BFkvaU7BaCmd3bZCAhNtV6Xt5H+4e46nSBiroulUhHVH+RZ2PyfqG60xRMy
ynIoGY4UyiBYYMCkJeCAijFLOPRKBed3m/NcVnDet/D70RpsNo4klK03LTTQXsv0
zJgdG8wgXVeNMpJVok2zBAKY+cmOskm7mJPaykQ5eFdvu/dgvG2CNtlgew/YJ8vp
GigL+Dd7ncQEUqrGBimy6D3gKr/Uy+T8laJaCBmIEc1QF1cRO8O/UCDXv/ONxFsK
KXn36et/DUsZIwLJnm0eZSKhnPvE8KPnDD22XBY2a2UtpsxgzKvy2AAMcKIpgDHy
QG5oocbyX3JC7rJmWyYB3vEGw7yAp/vcCGoUfgYoQYM=
`protect END_PROTECTED
