`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdKhRBF/sOF6v64Mru53MSBcJrXQgpMokJUj+8FGt3Sbm9gQXntfDzauVhL3Mwm8
1noKS3VOMdRQsxjSAAJsxsK2iOYw/abKlB8S2pMoRySU07Ee5O6SjqvzLsJHC6db
C/f+9p6e9dUU4Y/2PN+7wHysXS85Fql/NigX34Mu43Nlivz2sb1hu5hODnScIKWV
hb94qNV4EnTvlNa/soCpEMWYEDIt+sCE4WaRRHq6xM2UMXhG4z3cjXuvsd0lv3Gx
lMeuH0LPCGO4zobOHUVZLuAzTT0ruGzFKSuE77KM8F7tLFgfUg8J8+ZoTxMO867S
YkIizvt8l+5GPzniFS4S6bLcyB41WDKxDQWNW1vWw5OnZCtd43dK+7wPPYOmZinx
KD3eLa8XxfYRT/0TOQX2Av+EcDC0tFHc07bI2iwX/E3HoJMYAQK6ms3gAAnooNoS
eYsR8eUH/2IzA8bswhVRefX0Nz68HgCWqz40bB+8byMTrfAW7DcFfSvAkvZ/ZKrf
W60CTYHlnOlgoomQQNAbKOCqNSbQ/bGEQo1048MJZc/79/Ii2Tk1QvuAOGS8XsmN
BsqVafKN2Kaorvzg4T19tikL/GusUpsW3FVEBxUAUegqvrp17Y+dGLPBuIOfgt2P
Uib+dA6SzzRmSBcT6kPXOBShKWh9n8JQmzViAxe7ugLC95qP3Z8mDKEudkZnGQRy
XwMGLyj+V0pvtJLDmoD1D/ZfpJB1YJqPrB3cJtcSp/4zy/tWinG44BVr2tWJXE9O
y7U6gtS9y54+dy0TbWpih3wqiYrJSgP52rHh/hzxbo+o7HjkZs3t0yHQbZA1ShCZ
PK4NSegjlSV1Vl9BFT+I1wWKS5cn72f5eLrYierER5OAiJ8Yn09YLgz9TX+ZQ2RN
8fa878syVlFMtsA9ZLiyH4cYJemgqDMzCUHVhsOc3u+67mCdwg34kS3HlfIQna9E
aSzO7xdMQYdde2HJOhp0MVXsyjnbY7PMX1zsHfkv+tpCWg9IfAkMO9tM9CiQa4Or
Vtw3NQvsY9MxNobn050oBXJ0t7bigLhwAGn4BAKsRMui6l1VESgNTTVCyxLDAd+O
RFvnugq7NxFxLlkImGx2ApiwWD4bqj0uy8o2wVoFEbUzCq9ITN24NwxMYgkl/mkw
drYpi0VUDoMhLcODikSPboH/JCACPL+mYuyi5g7Jivk7eg+DaqsQkF1J/CWLrw3+
mx0pPnVumBJfDxtvhD6eK612d5xrJx+6dXEET0FB6dZJHN7AOpD4ojO19R8PaPMz
`protect END_PROTECTED
