`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U9unOLL4gyeOZoC6BfIoXS11tgb5h61BnhnCiRAPAIAdcd2UB5wCKToQ3Xkso8nY
RY6ssdyE62RdtpCLsWMYUtVR610zz06JCE5YKr/lFGuyhZcWLYmZy7MUrC2LPQGh
7F90KNCojBKa46bncagbRkMV0EYZmJxmV7113c6eSe5lo1DvPfqxh6vyZaEQIUSO
vvDumX/wou3dEITvCcWpqeBg4Jz258rQ8LeejGdkYOgeAFeh3cQ5W7/6MRNJ7j45
RL6C11Lv7PQ247ukkyW3MZrwkehhnEcIT4v6v32wGEQRNtFMOprrMgkiEbvB4vt9
u8ux8ruL7JNWo3cKNByrN6QXhQsDi1PFRzSUZBSRgyUceW6T5n9BP5g6poND01Vf
57h/oEIwPc0puLoH8qHfogVZyt6j9wdH3hlXMAMh39IclD/EFBNNmkG5/Xuw3dRU
ibalDDP0EXclIBQrGbXci2pLQX8Rq8x9odc2GMHkfB5uyWNJgt07iv4GwhZ/mry/
HbQDtN/qiAMYp6WOkJdTRWv/+5WlK4MkzgdT7eY+KAF3F9rnc4fWNuTHIfU7tpx9
tqmQz5ZybzssPTw8pI5IfItvQ9H9oJBduriQbm/1UUQdwHOAkoOaOdPBDC3a/DwB
C7259Y3ROJYkkA7fTxAYlW8wzQlPfRKnLt/423dD4BpO1MOrcQC7ZJSZabgcwZoZ
ZlqiBmYOCAkxLKdlCWH1xyjHlU8SX6WanwudolG68ui5ce6Yq7tgcCeDAzFk4EAJ
NRwE9amq7lDxl9rjBj3AGqIJa4lTJ4UOywR4pD60EVm7WBsj3fl3qMIHD6WsUJwi
d9xbUWsfHkSrMM00zfqzMHR/TxpAdYSwuDQ21ckEwD77kwvFYZ3+OTmSWJ6X33yZ
2GVg1LelXrtzAy+KjGn6m0n7B7foHbzUrsvOYWrFHo1wgGclcuRx4/WWiHSfsdfv
ESHZbDV7gukhUR/o7nEBcCQuZ0p5rLOQ+E0rC7Ip8cRSxh3+gb/f5nw20la3eNU8
FKGDkZCbxOgudFtS53EQRuael7GFN07Xi3Ht1jZwKRGEAa9wOm4S0iCvcEPfwwP0
7q7mmMw5fM9T3cpmKwRUdb/5PcY64z724Gg5xg69LadGGnkCHaFqf/hdFYmIGcDv
dP3RuQhHK6VNpTQxhjUr/1TD6I6w6m+8hGHRgYXgonqGeKuXjM7LzMIpqkgaHk4f
pc8TfMhGl812KE4gv2C9f6A8XEWkvLq9G006cxLCI6qrGfJmA/Pz4pQFlMMJhT/D
lDSDcP9M5PcgMlPJvvW2vqdyhRvj+UCUdYfcJsoYIjvAjnokPL4b/tsYZQriOBE7
rtonB4CIArGrhTif0fbRRCj1ePLyDjQ69KAStrj93hxtewaMt5IywozaizoYRYTY
nkXtzEZQ8PtQYkjXcY/JDN5E80LwBACOXqB1faPHX9drPVI0uKtgndrQ8j74Qz5o
eWSL1PqvwxQGAjNFBb35sJ01usVPBzvvPssFgi6iHLHWlRPI2LMv2pSNT78rEGQ3
QmdvygLeg/uianiBmdXH+LTGuIa+eiIqWipUrjkcVv5laVip/33LHylOL8kTnhzl
EIfwbfLWDdkB55nQjXLLdrLWyqqr3rMVUPoYPAaZ95YExlffTIBgjGMPUUwchU/n
UkkMPLvs9HTa/h7CC8AkCFXBlCbElFQMwQ7fZVz1pViPXHdGCOt8dSheiIof255w
O5SQg1HJRGsO4NcdfjS0Kn9ENBvnbcZ7qmy1YLuntSxnYbzFJyc+wDZP5rMTf2mt
AcjLRnHpdfa+WtOl031ifXVqaB3z9xQxNH86cPkZPoCJSJhlQa3q2cDreFB0LhrT
4gP8ltqkSYA2MEPd7LO2NeQ6tqc9ElJLmsfoLWO6+lesoWEQ0Xc0hiD0LRH4g3Mv
Zap9tuvwx9Fr5VvvWZgFDlXzASZ4srrb8TyDigKAKkmqij9I0khVZ6Je7Nm1Td+I
dPILQwjLYIG+HqfxTUie3CVZ6lV1te7ksxp12C7FnMJknKoWlx3ZDs2GT5K7m2iK
ziLVY8iPTtGqLx36JMQvVQumCZLWZ6HigsK+J06ZMaIRou9R+OpFiHbdJG/N5B5V
Fibx8upqv54xgtQMr2oCgOZMcnW2q2qk6uv0qAZZFqgv+rer0rfkzTZDJIuKBZ/r
ZK84yRGu9F2i+3Y++Yio9qfC/zy2wtsUg7TXo9IprnLpeuixLuA/O6UCaPSJnrnC
OF9GNbiPh5ux7WhezPKzHORHWOMdTAskNeAb3W4z1uVUEGaeiYOx0nKcaHCJ9wHg
Nz3mLawRWkWK1v0O+sooTsohbNJ5GLhOGUHWHJyfblZXBoejVhYyW5URsxjROE6o
oO5pp+xF5uP9VlA7z7EZS/Blm51jB5GGiRvx83Xb/GgTuLe2pV0SXIckpsONn/vk
5BT7u6NdajnEMJV391yTQf9tu+8Qs4hFUfQNiLo7CBSYGsMqyie/z4Ix6t5ehi6d
v6RJe1FLUBZiBB/TrjpbzUdpsBdct5HAJwPrC/jgXGG+aWj3l7R43Nftbiz2l5Fp
17H1zrwcMLeHHrv9p02QmJhlV8M5+6RvtLuVe81ZEtBvdq4kK1GTeXlQC1ChgS7B
OLwB/gVTT3NRpruZbcKAprBWglCpJ15urEfpN5twjnLr+KoLIgVyo2/hLykeoNwv
LD+VaP97TpLBB73rgn86Xm89zpn3/Kc2TE/iOOdzudaZbpyKsNGX/TwY5n1L2spC
FZHPpLSng4z1D8RZ8vieOQu1aXzGk9cKlTDFWeoKewp15psI2g2mWiUr6mm2Q3Q8
KAdo5Zk84rcExAYzPAAuZ8JJOBAzNrLZ9ftBVHfpibkCMND97W07hxagCauvbKPQ
lrT0F6cc15lZDFm7IYt1LbVQeb1lAQuHcsynVzAt9lfdj5DAvZnVzmjRmcAyeAo5
s7AnJYPf2csLtMFrpnhv/4HPfvkQwDlAhrht2AJ744WmvO1b1Byi5VpeO/VSbKMB
d5fPONb0FauOL0urr9zWE4gopr4IaRu4ZLoask2kS2EoGarxCp6g30O9QmPVJqRs
lbqAayVpdwtbyI98vGebZ3Wz/F1+xBI2lMkwnc0/KGkY6Hzjh7RpAZnIYup0bUQy
XX/5NnuFppQ+w7s5H9b6ta8I/c0UR4FC+zTrsKEoFc1ospAaMWv2nwx/d/2LXMUK
`protect END_PROTECTED
