`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qi3iVry9wTrbvoSnZy5JFWEW1JB1O5bjtxzJm/tcIyssrLfJMFdKZVfR3FQraFKm
ivlBqQJXRtvDLT9zy79YCIQV3IvWP3XGcOCvMSVjzsSQIyPzh2V2jaoB7AYVSkRT
LTP/YRD9rIUUldNo9HG6o+DoCuZ10HS2mR15M+reO3NhsAqzrBBwUeSVbUPJlYEf
ujNm2myGt9VaCoo3fBBugMkITSKgOc0mNm+Ic03cv7b2HWJHSgt0GlydxlJTLmnB
QXj2jJSbvjVt3lZx5VMNAYGDTZp2DQ7DkTgaej/UiBxAEb8MO9ihYFwAEC9QlVuo
KrszKy6th2LYdNVnq2lEwTcYpEH+GKz+9dzHl1AalUEcujA8ZyV7myMSo3ds+C7a
8EhReUNPSQpYjEiqh0tpZSLJXq7Mc1jitlxTGqVY17ygogmLJFUQXMoRO+JzI5SV
fofv0nh2P4szDMUf7XMkyQYGZ8pGIjdQdmCaloVU4StXCb6cLbOZjTrGnkTMoBHK
wZBNUyu5gfll3TzMo4o7IYb8hfV6GqxxdQ57YEzlFunlZQTB98VNj6TN6AmLnTlv
Oycx2gptjEEBxDsOz8QOThtuqH90nmyvQnWE+JlVxS2MgJFkauCbIsCtgYoI/SWG
sb/IN8x9WfpsAopXP1hVtHoOSs4duOgNIUdEHFR6wZvP7pdNu0ZdXWH0SEb/pVPg
dBg/WXLH63EExbc/mmayB57io9iUBWcJj/DluHjgGDASHjUOo6mNaILvrLqCRynU
7DCfGSonBelmXddCLhlUKbLYUtS3q0PaQzird7DwNO/AuQh1KziFAJAAo/sac2KM
nZ9RNEaHB1YcUNZUg6n5MdNW9KR2gsKTI7R4wDfOtgWusE3ceisaOKCIa6I55ZRR
JYcYbsn75jyMrylxO+fzgMERPtW0VYA7IFx7K6QCU++1beVXgaiXwXC0XXckcLhu
sN4Wxzy/2ksUyHFM03922wyRsN7kwh6XL3Pb1V1ppXYBajIAo7BjTwZ6aICrI6vX
sbfRbA4MSPVRZ7Eex0eF+tSGn42AUrrTolHsveatVXiXi1UEKDpQOApyS0+S7NIx
dfYnUiVQ3ctmYBo5zbcrb6aX79vcKMFm2mfd/YInHU+iREJOhluHXn+5a/1V3Or3
Vcx1TdX8G+C/M4QOuuv/6FgWmlwPth+8zQ2L8CnNifiAHkYvRoQ+17yJtQQp+QnT
dDsTzke7NwZqcoImhjKOZdBDmi8DUxqwxzYa3FYQQW+wogyBja/peB4w0LSMYSuF
WXeHrSzZCkU4FUJWMl9QAAi0T35APsLvt+ouQVqvscxIKWdFgI6Olz6IH69E4Sgy
x7fEhWSNaHnwswnurDGZuSNYNAG8XSZmc7BEHQQlR3/vCgeLWMBNXNk8Th7r0NOp
Th+OvGjbnkfZzvd3kA1djl7fiyUlHCD2b/ShCadINaIPbymIDy1BQXo+QzEnUNo7
bSWcHEAqFdtSVxZV+jNriR/E+qBrNdA7tNvCbHoCoX3tUY8uiLhSUPotZTJF3FgK
za077U1GWP98/dMKTEsSCyTPtvXdzGeu8XfIc0taVx3yn3Z8zPtxvf+husxRqliV
ORqfT0jU35aVBru48dmPk4kkuLr2wk3t2UD/MD9gqbc5925ISg8z3q+MNP1Fn+BN
SMpR2yKu3dZ3lI3aaWz26ohWM10d9Ga6c4YBDSZtMCJb5TbC7WsO+awopaN0j/Bn
PP1Z30f+48p77q9ANtkKCQoJe8cg2ZPwcB4sg+MQk6uRteBPL9NcCmjxiTRauBSB
bB74VmDGFe/xzeGfVEFiMScaikNz4NZHptARGUUkTOJPAqNyf50ZepOjrq0AHnrv
fo9I16lAwIevpXjqCtk/U7Y66apEQqhQxSXBQ/rRxASITADFCbPP4BgU0MbN9sdS
M7y598bIxbmEaUkSrvog+r7/GWNr2XkFuYqpAed/qUBZsBXli/96aYZXrtvOURgT
nR0IIFKa3R1XN43dsLG6HqKCCAj7Uo5IHIm9Wg3rdTBA0ZtSLHL9TKz2pdN0p5XQ
fgaugAHRA5vrrbj9z9sG3rxjO69s1hiutAWpIIqPmpkozp1pJi3ViAYzSrSTmsPn
9+Ac6RlNOvb/dhY++fSbJfkfBjY87oZCi5MbwmLRQuObN4NL1WrFETlTCN7ZVfrx
ywoYn1gaaidNHiZKNyvn76IQDk6PQg2iY2bqixq2k1bk9S7uxQCCp/AhfIEQs657
SNLToEpWO7AQHN629LkDApkswpvBwfcKKKhcH2GkbENNDBZ13aeUsGRm7Lch8qSI
TFNmiYjt0Rpr7xdzzmFk0Y0xXSZ7UXbG3DksIOD0U4JYS+5rfAk0BxWkWpmhdkmT
H+pcfIqwvDF4nFlgudcNTwhWbWx+4D/Jy+h2OoMVYuvcNfOwuhEi5Ic5eZfy/7rw
md7HtrAsIn9ZQZyb8x9IPF6PF6xAtNeuG0GpTBmi7uPhJXyiREwPplV19mzNUQkS
3sHKbDFp/phdK/aUzxmJpNlwhTJYXRgzgZtJxx0A3R49wP5kUsNL2Cbc9FRUAoQ/
QSbj78tnAdQc/LEvCgcbwr0nBY8ZunRtZHJVljAeRb9gl7WFHtNl7t1VIZyKrd35
Opu4qu0GRz8rCruFKy8MrYPxaef9u4OKBp6ymBxhCsqyRVR6ByfYfiFxJNJd6kr+
tl6nHxGZCWfBwZjH6JjGg5hRrVPBAGrDZX/RaX1vkyw8QaUCV5kBpY8JsJSZ7kt2
CQ0Cxty876kts0HfJhpHmbbuX9lNXuT+OWNdLAFUAzdADG0lyo1GwMp4akhZ61AM
3wm2MxFZ0igMCkFsnA+SFeDdQggOQvioaNt7dVlVM60hYriV5mVJF402vn6OLKAO
eKlYMzZz5t4cWrwbGicc86DwOvpLgAFKdiDbn/Cem2/cJmSJXDld6cVY0gnq08AY
/sUh+s6gK0GiMW0wQkmElCUgRYMqYsXPBaUMrPHMVlSInyGHihSuE8T7dEHKSJGC
7i/ltcWTkv0vs9cW6922daPYovjWZXkF91TkI9LwBhKEmepioMOc2YnPjAAanZOM
jFxrAV/nmBIPdvo4MtyXKFHNEbj1Fa12IF/0bApS3DCKNB/Di6Qdn6C1aHzf5eUd
zYpD9HiQRn9WOJknIi5JRu1a1xG19ilIB/S8zndDAEjoRstVuxkndMQxnMPZ+XIO
7+7al4y5J1IUCsSvRwKZdAnfvC1jF3l/WChDT1shkShk3JbgktuA+0YHKeDfS/7n
f+njTZD2SHBJBU7DrHkyRxQcNQBRyliLt0g5Vtfg+gbyuQSNpKI5h4bwOlOu4uZM
eM6OoMTpkCqFboGIbBi3weqG95XD6Vtjscge3OJpWXsBSv/IbMiTTpqYvFRcOiDo
eSxR1sQv8Jjg789E0rmplP7soWKQ21IgEf9uq8P6B3LfJ3FtkWqnrAD0cPF3HWYT
BO3Z+ibE89+4pMX5elubMkcHvqDPUSOAalAbt+9kSBAl44pVUQSQzW43eUZPhDuB
Wcm4VMeJqlk9qc8ysRtatook/htIzJ7D9lxRjs97YuufbjzDno635YqMT7OUbiiI
dzXmZn/hAo3ixIcxfgxeOBVc05pxKhZ/uGkXnd64u8vd4tEizB16AzNDMAeyzRr2
duzEM981nJQqU3YOuXmmaX07gf/xTGXJ6wQMK9lyRQTHnWJswAzIqzagDvK2TP/S
FJkoFpNf4Xv7jtWBSP0RTHxHM/hdzY/oOdhrVM6sC4tRXxnppR+vodB0R83O8uAg
Ln9lF3ZQ7JiUTRVvYhNSOsC1kwGpNsiGZT4ObpsLUyJU17BvHJcLZZpxK4rqulK4
uw2xv4JlwURNb+oO+9LEiXU6gWHYt9mICc1mp1z/RTuS3sFx9kKK3S8JrLBXKwqV
DHbBkCjzkZDc+omMnx7Oy1wZNQT7xSSLijREUpJgc6SCioMOUa8jlWLBypVRxLdo
6GKWdRQdpKsDiv26wr6+VWNIspHQsnXS9DpoFNMYyWRnlpnrkY0JB5kTLkClQ1BC
pM9wcNJ8doT/wCWLVNmcdWmK7jsf8pDcwyji0clNmlZOYawnzxZIzW/hikc2k0x+
Sr/LzKrje+Pvqwf76TqOsWRc2iC9wNkNNMsAIB54NCMD7829i24JEMXQ8Cj3cIKx
mxUfFuk+YLTTaSmYFRpJpWEfQdxmI7zOu1ErO8FkcaLooI1FCrAwYPaobZKgqFCR
5ppXMNQVIQWuPS3iIOYheOn7eiki9YT+jTvKzxuilh9sVAppIZDYhssq7tQ0+rmI
q6WY2WYFjoP7LA5U8XHkc5s77xEnWGR2Oj4Qj9BSSbDmCPgDvGvJEwUuFwYd2MUR
9kbD+EXs62D//M4fqidPVi+gXQtOM3dn/Gw38Mslicn2bnp7IBdJIMqiekOcYaT3
ce/Vo+2f9D9QiZti4ed+BGL5Uruabfk7MuPPbfaC5CM=
`protect END_PROTECTED
