`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30UCRzmM557Mo00dmEeU43hrF6xZmzUP+Ey2ybmN9ZReEGB5cFIKYmHyXTjvOZHQ
dm/76/MWOXNsKf0LKOXElxntERm3eaTjsj+uhLAIxNMvdgWbxa2dWnpA4AowYSgi
8mrSGVdbAk9jS7SqCE4gYcPOdGOaxMo55hneEOkF2TDwaf00nHZEuwvoE3aw5690
VKCzd9Fvnv0xB5AWK6rBsChF2/cy1HWBfk5wsVuOvBHnuNXaubF5nEg2c0jFvuSL
WZa51Cl+1KW+E37OxepKds1d6sFqjCvI8hPR3fGhXnW+gHmDxPrbJndyp2Yb62rC
8OShzkmhWuEt5OHIXxuWN1y5CXEXUNaIjkI1m5ykVxyJykh2kF8kf0UtveYKCeCR
jtt0IlaZ8uup/Fcoi+ezsi21B8w6pYAB5ZiGtpRuZnkCBRpWe4kK+eHR4NfGB1Ow
ja3VjJMDN+faPM2pSPuipK+w1HfX/5909apgrgk+Fwtvar/XflS+vxx3ncG1Ossc
B6iWj+qGZk6iUoqDQND4DQji4MIFjzquLeEJLQEV6gwdLe0FsCdbVHg2LFY7n7+F
iwxgkuHR0K36k7hD+aoxrEKbYXmQzmh53DyF/k50He6rIBl+151Q+umzb9qmohJm
t2oSsySRV+0EBIgG+TvsEwMNZMUk9BwpuAG83ZH7dy0UstpZgAa7nHf/oGX0fRDJ
B37n0XBN05Xa1jAG24afLU25PK/hK1lp/1D2/DlE4lIGL/+gzfSsgdurghe/EBi2
cxMNfNZ7YtxAjNqLx79KGlHy4BrUNOSccQWgSHT6AvW3Rynn+wU9J5IZWoiDkMBF
Ftn7Vdg8+2KWzZR3D+kJ5j5Caaj8n4OyKq8mmffvGhcdtXl922PSBPWqrjeGSZSw
gtIiNPCfpqJWOKjK4/H/C7i/RSp8GU9Xl1iUuIfH450iM3ALVRKXiXc1wzJFHiKB
jfIHGC9TWASvo3/BTbv10nob1VZFMxbL/9EKBN2r92sknb6mVY99OfqnWPd1CKqF
ZMnnY4efiHZQwO/3SWVW1OsvxYAw4kllaXmBiFIJgcdbpYGKfsVdty4SiGUPgBjo
EOXyK1eW3MpiydeZIQNTM8QnQcEWdGy7MLSqvFtR7IJAIpzU6ntBKEnZkD6J5ghj
Lhk9DUCqcUteg8/m4GydJx6kWgAEqD7WnYDbRryBShMCKh16DB5nJ1D9WP31QWqh
QRIgEk4tRWXmgNWLao35ASsspczcXprBQjbMA04kriqE36+yVIwdn9hmVKCFpoJk
yCvO0MjtngXRtobd/VyKB4YxzwLlbwlTLp7kmMJ8ijTaiOnDXNsLlr6g1HKCpkEO
62A/EBisD73TGLQVL57fJpoZtDJR+fGK5DnKMLn59kvlAKO9Df1zAe+uHktdQDnp
O/2z340JseIncO+uJ+BXmY6xhzVHavHlre+Z1tROVS22BcBfiNb/eCU4+H9+tYeo
kG7U6OzO7NtNIFdjcX8h34ZYenCFKsdxv9/ETBe1DgTUNdZQzWIzax7GxlVbJpPE
AcjBucU45ZKff3TeBsFyy0ZoW0O7kqKjl67elO+vAZIQxZp45LjNRom+G+JhhVTt
vAMTF0YqZGvJLDaN6xkcBfhU86XAunq3Y8ajZeYJV15D1S89AfFMk/os4dTBzZC+
`protect END_PROTECTED
