`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbSAS1KNqCfpuH3Y/NrXQglZ5dLv9jSET9bNMs3pKazGBxdXr0krnpDEYQZ9wm0i
1EIZCAKlHcWkU4FIt9vB9W2Z77SW7yQCHRbblRjLlE+1UPprmpIVSwn+UXpY/hoe
2MlbD4n+EJpESGNAIMu+9cTsUg3h+GLfO6OSIHxA/HbXoOA+IPrB93nbEztMubHG
dtN9hqhVhw78qtaVMIBX6e7w2eKBc0VIpNIYrrAzWnFuhBKcXKCjvG7yCYrF5awc
RbdHMVcSRfbrCH52jwagEHZJVnnDg/0Ep/fpC9DVQr/NkwZ+3RRopJy0O8McZzzr
G8ziHmpgR8iJIAlrOWhCyu/ZI/U/C+RGuu6PN4Gk+Gc026PHs23WP9/O3xm670LS
DHBXqZu/78VhrvONfr18GWVjFgKbjbmvbhInugDcfN7OxTNDC79ooKbSMYL4ZTV3
/kbzWNO5Z6kO02wkqVHNhZAHKMey3/gPQ/12rEXWCtaigP6klUYGTs1p+g6cLCGC
IgSeoeGa6SEyd74yII5dpxG5XWMUe8oR8Z+exghhl7gQzRH5Xr31dTnykFfQoloT
oa/54olXxueTP4Pf8tnX6rUCWKmBltMF2H+xCKjlDn8XRJnT4yrlzRXmEXplJBXc
YSXcNC8KLKB/Q/kWhwBmq74xjD2sinRY2F8sHJzDWD8n7BxPY8cj2W+dXequjShC
GNVrdep0Gk/nAnJhYlw8bfqVAjtzqbQEzMI8KeODzA4RxI54X1QoVtyYyiyuqKlN
hFc5OsJYg9y5Gdy4aLDo4oarmKtohEF0TsZjofmnHP/J6ZNqTK6jks/eyjDLzbBU
MgIKE7+czX1jjA0VYDID2s9q44YFOVCSRwbTx/u2+lg=
`protect END_PROTECTED
