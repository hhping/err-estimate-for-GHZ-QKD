`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2OONLn2qdhPKbCYggeCiCohgCTpHy5vW7fZStw5VN8CNLGotZqRKpx9Rm6fYevgy
+5lN1eI6BqoDEHrihxjvXUfhv+WfkxFUJkapOr5hqv3K020V/1JKyN76YzZ8CYS7
Ome+c0vcFBB6LI/sGLZ6rHHquhOfpwGa2oKXFlWQDSVfTAwAQI+36rUbI72tTfm3
o334+USAhoCeEoprpYePdocX04rHJ1ZdcmzrZebB8B/3ID1F8sozq05kgO4oNbTT
wnwZ+T4ZYDoWKcoARPgp19gGh66rBSVXRBnAJLpOHQUuZUyU0TUwUdt0AEv5aIT0
OzEzDyczitoqporIDCWSHOA4qPsdhpFHfZ1SZOG1PXkVm3PcX1oWQp0PXFKJOKZu
VaMgK9VpHbQE4vRf1yzYkkcNAreGnHiCKEwnkoGBy+J4R4/HsdWqlNV4ncH6IuRE
maxe8UtGaL1r6DBzUSo8+bF4SwEDul7VrXenYq+hABPIC7GcZJTVQaBgP/9TIqUC
DOadvwjarfaSQGrA9lkFKj+ECli+NHRg8IxCgsIVWMEjaN6vjmkPj3gNqxJtUrhb
xTWlB8CGAt3Rx3RebcOSwkZgloLr6UqsxvRpZ/rpH14F7iJGzapYgcX7KBLBBCW+
y4TvgEqJ8/1iF2gyLpPfSVC/IJU8maODxWpJXUB9SDQ=
`protect END_PROTECTED
