`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tu0ogtmOgHQP0RQHzxvKayfhUtXcfG2H4TkXgMe7JJgMtK15UHeonuWIWWmc2gv9
tggNpKlMbxjMwdRZQ+pUvCKEkyKtWt3J3VXf0tmHSiUQMKb62pr4aXEeF04wBUq4
SNEcH7bqgRB2T+052MvJJlxSAqjV+5CQ3wuffZu2ZDry+nyX64nJaDWYzi0i2abT
zE0ZVcHghhIsznOFiNgdSimjMwryGxBtBBOUx8zlnQBIqLGMU9DBL1yKZDeXz2n9
BgbFVV5ljDjHcZi0beBPANr49qGdIEeEuDsn6G6tcZrNDpzECIG1v3gf1KcwH2U0
Bsn2rKrgMRhKD4QRz7jS4u7R9vFopnTjU0Vy456U7lfo/VMDtXVLSzAs7nPt6zmn
7au6VpMSdJknGmmbX3OcR7rRO827LkHcN8Qo007simkFFPP2pKzefyay53/VuY9X
uF60T4O1dUxFkxFPFr0FIZ+BN3eiwf12MEC9Yt1M86AWMPRtt8q2SRMxcWMCFa7P
Dp1exgp82ez/EE9YWH/G8ywmXZRihKhTlBnrBh5yV9lo8a7vqyosWymeZLHkXxK1
HX/W7Y0RAh1rz4Bikx3h8uCmBNA9xESm5l8wmP6AkR9eA/SmkrAFlF1Of3HC9vHq
0EYY+x7JkNgCvtdG9ozfRMA6Q2IG63J+gcW/m/qml97kGEkD08Hu0vsdr+qQq+ZM
`protect END_PROTECTED
