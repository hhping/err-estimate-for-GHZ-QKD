`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7duPRxbiZ/hCTWyvPdLQm07y9OQ4ofvA2ajueEGQhJjHLfmI8ALdUdM+onVhIUz
pc3wfCTeTQN5B8d8YJjHR2rte4n7r1xqAMPQy+AvOrtcAents6hJYsdvvjaerje8
ZBVDCYTiQSMziT8cZJZKCqxNDVZwYL5TJVUXkgEcpEPFQgoL9AhyXAvDxWsc6S/Y
Db9qXzg2LTN3tXex/UtFrrDv5QOU9dGRu4kvPrMh0eMsqSvR3fD5IoxcJQHrADLA
mHvpFJreyrRG552oeM+pBL4nBBfF9lbqQLLN3vAFTAuZpliNzAW+fB5qP7rKqFGQ
z27vFlP+wWYONfkhUMbjA65y26qkOH4/tLVkeVm85lk59/g3F/tdXx9FKDCf357R
uk0yoWM9lhtCqsqVfMTqBDFtvgQJvWWq6/PHDVm5aMcA2mGah2pDNzmH6YeP7Y7u
9H1pbGXJxPtAznovY98BUZOT7H4MrzFA6sMDihhxaa1m2vqYTNLAZ8FdDQdp7Wc/
2xY8SK+xD6DfpNotfnCBxH1dV90RPDmifVA0yCY7BjGgPmzPkHkM96sysdj8h8ZE
0XHYD9wuRllX6owTVY/1sqVy4kKUz+KOUG/roSsJ1uqKl//Yx8KVu/ejr5MGQ0q3
VXtGxoNWdq5v2gt2e18YLCgzTKdDvXdRI8Iv1KospadllymqBYXslF/BlstF+z2o
VaS4652H0SDqn12VFpr6ewgdzWYQi43iwKC3voUOrs8KYFD5xebx/+a1b4NsVcEE
OKY/ze5HXAo41YOCkywM+jpDdZBP3gPX5fFCkOrKweo0or8DN/hVqtfKZQNcuBSi
2ZRKJDZYxS4UepA1Qf+qxkd3wAVtC+wOr7diXZhtxr6KPfJNNo/fQRKJjVW0PC12
w5Viq94ukVwlsim637E1jg7K1UKvuC20ycvv2QmCx4V6Ek6IMDaEAjoj7DckyzZ0
UVuFZBwG1z1dfWDmhYGlaDiMoyRFObm2Nh6EaDDA18/PM71B4VwTkijtBLUPkvob
ZhIQ8CHAjPG9wUCfdQJgYHgV6c41zbKQLcMYASwthVhOP9nGuo3n5g4hSR6oiMY9
pqoR4BaKW+k2cUoXseqXjRiECG+EthHD9/FcDgotOI+v+Lgq93LRMF/uZ1Oan20x
rmy7qyqsbeGWQtfooQMPT8/EQbKSmieccFESlS6HuQR7IPOtGR7nBSqHM6FXpeYO
YWqlEJYJ2Pb3H1Y5Ji/tijYiRvhe0P/u2hbzwaLgZj3RbthQY/Z/wSAxjXtfgznx
sF0Gafdyu4IDjoXLVYj0wN1r+PR9kZ7s4tMZZHz8nu7cee+k0M+MUXbo+ob3YrTh
uZ8qqw5f2+eGI53PEVX9gn5C/GFVYplv1/36QxrccB7PsV5hpuoFpxrX4S6lW94A
cx7/iHi2+RYHrvLsNSY0atw+IhYE5cSHApSYPJ/kwym8BbEUxPO9+JhWZhUFWudT
UMDsRtQD7F9fir2ll22AaotUK/uwnbENgM5zE+DkUjehJacHvTe/cNk99tYMp3ie
7I7q6wVKSX6Ib+GB9EWfvrkZEUi4ZjUb/gOMdlgcr6WqHeVspPtgYwoQz6vIlrEU
XFzGHLYkPwGv4vm9EBC+7g==
`protect END_PROTECTED
