`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rkD7RFT4LrBrmGV7ciIW8vlZKCSUL+2oktQCE6LD3rhl9CZ6qqNxh2qugltFrXjJ
Qg++hV/WgNekSKN0RhcpsGrRrBQMStelL+DgVjJrmpISuX1tmVGUlU7CAzellHVg
/XQT8kMrOjaHCC7pEjjx0EX5iSa4t4MzV/OkseMRpIbBzFiHZp5m+2ynYzXigXCq
13Io0pgeHhhJleAA7yN6Zk0+nh5P81t58zVTczoEY7RXPdZtcWy8hmGxUB6/Xx5s
36g2XAfF2Gmkzz6/NX001r0CN95bPJtuHOoXvpas54EDfYQ3VTUJB+CNmObaPWHJ
rl5NOsUCHWmuUq+URHyJAC7vVeGlIWqLVHPlTmdLxornPyFXfCxyXFNZwWJkKZlH
x2Hn3HVhCI1+5DY+mdIRATElHYWmzTtQAcXJQNEvpN+tBbz5uNd7q1yiXTPQpYNp
dAX0H0T3IfEK+ebZv8r/BIJZG5U+c2Ywpb2ZDUpgrXPvbagPwX2UjmA5lCx1mvKb
Q9pz4s6KN8Ad9HfTEk33lUEWfJXw6Y1JSs5Q21GpwypPrxJvezYaqYv8FVeicKvq
cqurxKC+cWVJn9Yxf7ePqiEzA91mcHUptVNkg2c5VjBRdYwZYatwSu2O5IqcXCb2
BuzlBktIpbjsPDYE0QuRnVhGgQc8CHl1w4qO3JB8QphnBwCjHJThDwjZ3NQrh4rV
YSYF3OywBQsSfERQZ8V7QaGv7vKdZ/ojU4tEOqqujHM1ztNNifDd+Db9Oi1e1LGY
+qU9GjkAxA5JAVSfB3n04g==
`protect END_PROTECTED
