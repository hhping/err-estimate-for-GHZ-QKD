`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJViF2e0OCcO+N0nYWpUkAZjxvSfkCzyXpVUsSJ4r4mWraKbeJu386nRPd5oW/Un
2qT6WWq6oYAOdn7NU9tm5zK6CWv7MH+RfTdjiNpcGXGzgpQj7UzNryHsd7GdAU2u
DUNWIxCS+4dssuYpDkPmNNfxfyi9AUG8Fmzp3MeG8ePpyPhQ+s+4z85sk1QJ3vVN
8gXD01AlVbMk//KmFQuDSxx/082F72XEtxGmK5AvOYO5G/1nUEsf3Tpnfm+Qq/x3
fojkLGGGtZp0UsE5aSWfed25/aHPw+pTzY69MKGhQJxUhFzTnxS8/oA+U7Z2tOTj
Bn+2lOR/3yuaQVm2pgbJBMfygW6uAxgYJYHd6WH4023SxGg0rUsC71YCqxUWP9tX
CVpKNsbPIht1aYRn+9+nQOp6PkPZEb1Y4Hs38kPvjFDDti//pqvB6AvfzQS0YM6K
7o1RNA/ZdDdK11321kAZzU+iccrk/ZoAQy3it8R8TBfnmnvh21Vr01heuSvoWzLX
t2oFsjXzD3ieTh4VlM4XIuhOCO79VCRQdrSyVrrgYPZq54od/vtjCirX5JG9QZto
fh0D40APW6l8P4nt8IyEzMz0v4Gt/bqwnT5PXYXavd1+aTAdEpsK/JmbbIakXSYZ
2aQxqDgxHxf+oeOul7OL6cwSgm5xafDkE494U+D2w9eR6OQ8L+UbWdn5kxS3DWS9
h2mF4pHXx1TvrGSzBLCEPgBfJlW+iBRfK19cFk36gOqm4Y7jQvGimwMULcNvlU8X
nWNOk+i6W3AOlTGXPrCeD98xFbCDOjRCCCXaHSQ9Kb00YsgPk8VtssQ4j8R95aAR
KxmLueUNCZFxxrAK2+cwfTDDbhRvEjqSiwL8E6lNLtA1o3k+yGu8RVQ6cO9G8XS4
53p7IrSb7Udb745oBa0HchMntkWgznzwoeR4wQySyNuOaRU/g26DAQ9RC86Cm6Kf
3flrI65yR0Y51ZMdNnCmnU3ul8qHnnQeslgGMtWkokvtEldlV0kfg7Zyq06w7EJr
sS6PF4qEs2f1eaHDWdBovJtgkzcKtLlCLSVHaDV/wzXQ233a5tG6OM/n0TP5Qcr1
VFNifoHyhI1clkKbGeyGUI61ys4HoZoSfzXOzWYm5Os6k9xbKKMZAU2wNAwqnysl
`protect END_PROTECTED
