`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JqsO9/5180iaD1sKMNSZyyk51Pyk4QMozxyOQw9sq6R+KenVghgVC062GGNeIaW
JpespYKZzlzzJMLiWRAhIhwUS644BWwnvhsFMv1Ng0mWWfJGEl+IPZJnjah08HFo
c1ilE2+vrUyKAEi+oKEesHn1MWsMwLmVHwb9UNg9WEwF3WS7fQeZjzYfUaD/IHAz
1a0hywtatLGSTa0SMj3p2V+UoyS39cgDpwBpH6P2aRhc+V2cvgseOXOQ1dAuvMmO
KR416Smg5RvXSoLc0iY/RTRsd0EZDx4QqXdZqO7ktsMi5znqL/eBpne1hMp1WISO
3xrypcA9dmvBNbxk6dHKnVII00nV9WC77aS+hdF/hHxJwt3LtnIPydlhdOouupml
evq0OpOr2+TAvJ0X+nCVCFwlgprB+TIbqFFkDmNZs+CRqayqwKEYI3T1uczHObE8
840cACjD1zR2R0IzuflysyNI6jxw+WDSlNe790Xrgxbgxxmz30uKJ5N1QMgT72Fw
dOFAPzLAQ32neoouNkzM8/1Tz+nPmvcacwbhyvsfklMv4u1PLx16IBsEQ2NH0PvY
d+5N3Gn+7qH3v5URjyOMR7gz7FAzgqbTLdhj5WKRY/p4d1V4Gyg0vW1X29RkZ1c4
YWgA5vvpk3//5+mk/zcSOmNYcqwYK6v7wUyjyP0m2GOLatRcI8P36hzdz9JlwbWf
f9MiyLvATBU2epG6mDuwsnwYckKCxIWI7UZL0v9jvWfI4pu9r/Ma2k9toslygFSn
xsH53lMJdAHwz8/2/PHRkrl8a/W/PgFQB4zdOw80Pu6dB+aI/Nir+Ld6yiIDVEGD
`protect END_PROTECTED
