`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDaAHSPsH8zXbtckNj9/bAyXmbT8Pv0XEUvY8yJ19RP9KVrzbbGS4xC+x9m1RtYh
cYO7FDC412bhAYZkHjNzIOEdm0tm8Ca3pfnSCEEVczcAgTJ6lDcVtnoLvEGZB1Ur
Ya23qONLqsLp+xDPgvgKo3bsNfU4fLZyX6rbkn0Ta0FfWB2oNSh31Avj8RUKcKlF
LX+dn1JCGseY0Q0hOe97vIAdB3gjj6tlDYG/+teqaaMVmwVE18Tqil1KmKWX5uh3
7ITVadi5Mt2eP8UIF/W0bMidE3I1/qpEPuH3zfvzhz9Lb9h6yzXAffcAT+6YX7W2
kv+10uJWfUgXxJkihbpdpM/o35ApJqxi5vsmB638oWzAAacOae0NGmxLZU/DZ4Yk
5PYmcupiIKpUX6U1V2im7+SlNrm8e8C6GSAGzj/LppENDDZ8yquNgqba5QJFY+Gw
tngfMugS9tHe72zoTiAob5DCnoQsVxYlj14LB3q9N1H14603igNclUzCC5Gycr7T
VKdkjQTTpp9xyqEl2pMQs2oA8/lc8mxDrcomHy4vFBoCYs+p53AC3uq9SqDADdhT
dTMMYCebBBd0O8tJyqSm5K/SG1P8pqVXp+1nbQyV74kyPkuWXBxLoMmeyXUHPNkf
ggd7q7mASkimSiNEY8BZIZ3y2FPLZb9quFqyBbGuiar4UOIlhC6jpNnx7aazSNVS
fN8tmXZmg3OvNPgO9kmbSzYKEUeR8k9Uol1ddm4G7akaVlHbFhni8UGbjzEGS3z9
dH2YvcNXeGeRjZfG2jeat+Rt4jvkWoN5N0NVcHZmysXEGcf7Qsbj5In/6pr1MEKZ
b/dJU8snLDk57gl5GQE0T9y1LKg1586ukZjSi1Pkj9b2+0w04Ts2leLoBVi/MEKG
k8t3cb2jxp9qtwH2TAa7/BxBXcwUWHBB6S9W52NMITM6WXGhy7DxxXqvI1oBI+vO
q725gMQT/FS9r9SG4i33VjO7AhHZ19Twt2djh2oh3REKEHDVgP0HQP4gRqhpja43
Ia7SjMUYbPMgAy0naEEhXAlQVA+2KVUyY0mt7TXaUTo0KGFdHdd1qMuvXIgjRVeE
nhZ49iYTP8bbkboe2IvBg/Qh+G2KqC/Q/8mDtQJZEWWToNEPKYtyCpaq/FZ55cuV
dhnA7wLgGcwwzpQR2Z+5MlLXsWXz2aQq+1A6yB/DfNArmn7Q5siuez9ZhHbh36IX
EvbDAU0/lCgSU9hw5wO5uTg2YjtSGJjHAD57ozB+oMnvMASJ51wTEEW/TH3Cvd3L
Ka4jayW+gL7MmBUYwLfiPWFULtFZUVap7eqzktR56cpvIdqORztyVVitJlKNhVnQ
a7sP22MtwTvU1JfL3M+CwVzl+ZNdKRXxo2s78VLQQahE0rfispsP5tewx+UmLD6J
ovGO6iMHLyLhmWvNj6jfd/PTqoLdmYqUDBHp0phdsQU=
`protect END_PROTECTED
