`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSkzZdm/QrVJQMDEDaN0R9zGJAML6bQBbyLjUlZpJYJGdO9vJD0UNLofl54E9b3i
vOd7RGtQQwc8yLui/67kkJxgl621RvLskxZKmg0oLGXkeqLrJXyT9M5/BLd7fxDc
7UpUUTCdlExQfza6JwOidiETCyR0XjCPVtn18hwlhqg6+6OwF7PVPuuQ8Lp8oyRI
u/S0WCCphKIKLEowadfATXXopXaDZe+0pzLacgXpxedozyPa6CLRnaNzCeVSfnY9
LaCTNwqYshm9FrvwffG7OjsigzYm2yBpK8qomy4/MkAp+Grh9hDPzP4xUEt/1Ivy
u3lDe3ACzThQiPRX2RMz2LbQNROYIbsWmdZO+VKYa1LJQ1UfSpTuML+T7qHR401a
r4oZ08+h4kzLFlCfL7c3+92jvUCqLmfNGBgjqWpkVK1VPrLqBFZR6fXJf/HMHN/r
xqEb1NOIYiagjiQrE0A8eaEmFMyJrA5KYUBvFwuGByV2TxrgtiPqSTiLwSiRr9OF
WDlqFC8RdYUVftPi2N8vQA7TxD/LfO27/OrlRHeffGC8SSuJH4CIutmEdALpWN1v
92WkUMyAqylqRDBrlNGckXFyZIVcR+hNFWU7mTE2BFj5Ekk5njTCsGZIb1JbIkrF
7lgzrb4nSt8YHghpxfmjMAYjDpnvV11Rnext9sWw3zlc1FVRfBcnNI5wF+RB0s+T
HlFak9wkyaoSHZJIG+2Ki7HSLpiy9tYQ8O8DNpTd//kG+R4RFIykM5nbiXhqq+og
tGqSRxMsIm4IEc3iRNn/f5jkiH9xAvdqdVhrk5rJ85yySs7ObT1ETP32X8hKt/Ge
B2gr1S9Gojx/TjyomPbe5/xMO2Et8uyZ2ILpsqEEwVbmG63Fn99f8wXoWqMvXs/4
vZ4yg7i5n9armfukDzLEzf/KQmk/0DrMG0kCiaN67g49tzI3m1YlZeFZsSUib5Q2
hgC3NwYeTv8hadFs/xsybCoMnLQjzDygVk2CrJV7rhqygyP6+swvqt/C8ikwl1dg
IK0b3T3C7nBaUQjqGwsGX4y70QyO4IXWh+UIHDaCcDxF5D27GXQfIPN/e+bbiuJw
UwngIFlVlsgtHv0+i4KpaDgHNtcEtdoh4AVN3ctTKBrjTvn0sDOt/ylxdhIubFTm
Pie7QwV6Dw1nHIsPjcZpPIbBTRwr5q4cpAo1+ulGSB1Elq5gQBv6v0Cx97qvCu4b
Ptt52Lf63RRyDKhOmefH3ohtS0/ucq+RoJJEI7OkVYmpaLtOhvJQ+Oa7lXJiovtC
Lvv8U6HI0+vQhp+75cs6Cl+NZe2pgJckEoGG6jC8hwXPK7r6WKfY7f1MPsA8mSJO
bTOy3zZZVwCtqEsmmnel2fJ6YNzI/xTNKIcqjdN01gr0roe6qA5ZWRhesqY666Ze
cj6VbxiswhZzE/PUE9mDDiqRP0RzyZJbWPO/SK50iK+wgXX4/d63MfHxZ3aOrbwY
cvkD7AY7Yl5cgcznE4UcPC400CCGi6c+2xCJnmPDAFeQ4YXOeya7Jzf9PfLNoakq
sibeQm0NGJkPqC0JnmhO0gVaPcvTcLKbEomiMTNJ1VfwmU0YBtFpzZ6cwd7cPmC0
eO8//aXvitCu9lxsBUiH0ZXRkUYlxuVyLmZDOEBQZUsGooQwo+FCt4WnMIlehhar
4uHfs5csWOmbJjIUqXDbEDqbgwzB8Q1HPW9M4mnJL3QFKKfZHXQWqMBOTtRXeuKh
xh3HhvdKv4icz7uBnP4TG3sA0Gre3QAm8G/Zl3MnTCSVXDwvmCEqh0vOzqzeXYfM
x/RyRvy2BetztWVolWtfLZiMPgzUBjxHUw5dsopuu1s1s2Cs1SjCg0dDRGZCyYs7
q8ZJ8lx05BnWktKpwPuYhYK2VACjrZSUukcSkT3KSc25eqXvZdtn7fEq8DSVcaPm
KMUw1Ql1N91CUyyWgH/KmV2totkN4NXXc06APzr+R7YaI3oBSY0+wRjjWTe8f7pj
1v8GgsRgWvOzYb6EnXZ2SrWkNAbY6lWiJNOwPFxd0XRbfH6qvKa1/jMlMrFm/o7A
oAyEVX2XKyNziGm/FFaijPX0wiboG/dnjl9BNlnNZHyeS8Nhs4excGdiLUvdNLRn
2OBkDg+fOlZM3hb+HLcJ6nvZuMba4f7fIRvdA6L/cxZt3G+rDX5gHaBmGtdSnenn
otgnu8fALQIG8UAS8JnLNqB5iGZzrMoVIKLxSs2QBIdD1aRBli1kdC+n/TlmSMTI
xyvX7woszc5HaxJxZ0RNqb9lQOOYWxVeKynid0Mc7MreFViurY0q1Du4CVjZf06c
bGZehYhe5omZZcTxkjzVBW27ceABAIChD8jlIPz37EHNOkN3i/YYnWiUPdRe9lKM
g6TCUmsc5CPrN1x5TrIp/PMb9ifjuxJthAqqrnTAyA0w3AfhC/K6D3vYxnOjzB04
GjnFcpxI6aTtm7YRqpwvG1E4FbAes1UY7Clc6sbhQPCRVkTWhwkDFGtKHCSaHwTp
RQcG1r7CyNcGqIwR1zHEJdkzRIHpVcztUruVJ7zbTzNEUHbKnSOQlI4XL8fA4xXm
OBWtoBBIDWGfVx//dt0e0B0yIMeumwF0HYT7pQujDCTF5iwOsXDqCDcPVEENUOlw
06YEO3oVljsRTQ+zAJj3+g+WGqHz3gjfpVOpzsAOCNO61n0FfYIPiJZW39nLza3x
uKIw2PPlBNOhE5kBkGxj/17GtLEy6zwRxv32hZJhC0Q3XwslOjnEA9F/XuI0W+fH
IyjvRJktcqznaiN2K467+80SwnxHJ1qGamQ8FrKt6ORj4vsEpeA/Snud2MvZLvYW
k2ZWldBUgkuOIM/LTjJenpmU+Orekj1lnMi50Ma4uAdKF38Rtrrjk37KoUrsvxyn
rttFjxlp9zJFXmHAc5es6i0vC9JDpLk5yFVz1qyFRmsRFPzc2i3sBvr/TvNirhsq
MFJ8ZOUcAnBkT2i7BruaM7JSwLg/l78d9sXJBqBXvuxsZm9cfcTKE88P3gPW7qw2
u93pao0K53sSjCeKnVlV/RbGSIYHo1cphEOV6T8hyXIPdf7MHaPbgiep8LuL29PS
QtgP1mlugE/DCY//ISU9hmO3aHXmkp/KA+VONpF/GAhP8sfBZ2N9nhxzpeVHejTJ
yEHyTPUJ8fz8p2pgu23iVCBWjVcRm2eDzWvtSUAqkcRziGHJDv4k40gMs1Pz1JPN
4XJ1L/8heSFUSO8X5bBjyorYj11s/ncJkPW9R0GIFSJTtFiEhDtDcji/4EMGersg
E4yTo1YWPVdK+FDCUh6NhiksMYrWy1TtLTfYDiTItRJKSpC8pfULX+M0TCwXePQI
eO2xbWQ7zPWgehcga+PTg/dCgyDD5T/cDpdW4n13SSEztpmvQJVNOatuC+A0u7BK
HprzFe4udtHYo/1OgoWh8jpMZpnx/6UD+m/57VwU6XYp6zYsI5TfjzlsztrWQpUh
Ht7GOSOxaZ7Bp8MeVbKIqtAMgPJYDL19ZygDWJmM/RyZXFG/wpPy3cjWn4PRewdb
4rmRpTMPO83MQj6/phclucSxWJa3U5g4eF6StnP6ZcAn1kswLc52YSph/1JjVSiJ
9xYEIFoiv9nHvlA5N6MW3m4cqbbhvIzobnTrxMnQ3o4eUgM6PpKTo9gMf4jS1WCk
0OKCRLmq1rvSO/lEmLV3nxBnnHC66jGBpyNDvQv1USpYBotJf2V/0urqyVxXhCZN
ZFTGnP3RztXF94jtEI/mUqXDTcD43g9Lm0pWooYWIls5Q8XmKbsk/e0gsys8bIub
IBqKE+KFpsKYk2sF6jtF0yWAQfAw6KEO6+NCYTAnXJvvzl3tojyaOXtdpWDJiNQ2
sK7fiSQiWsTBrhLnyc6YuT+n5ub0sIJoG62h6dYoLOX5AG+X5THSCdkrgJWzqvy6
m3Xb9THOgYMzPQTklgiC7fAjz+TC+S6ptrijNjkep7dB6RtQM84qR7/Qj8gjla1g
iFhs24GOV4IEQKuK6TFj5GINLPNHXd1tOw5pfyYk+4ny6VBLmTjHkwig7APqgYWd
XKVLYexDOrNbxr164NrofceNSs9yf5pdG7gMHGS8jL6UcK+FDrScFdrUyuIxrqRQ
nnepGMl+Tv+VrZslKR5OGrEUR6ek8/LYjsSLSolU6ea00MHaDWGs5V2G+bVi2agr
Nsa/hrfEbDzmhXlzhwELbN+BqcWK9Nj8J2wXwKfsc/2GU1IVP5DEq3QSdwRYTZy3
qnNsbDuJQbMMcZ3htgihIsllr0/g2vdJZg2qmXpz4T54KaoOKuwscCjuJx4eKq3C
cSSLmQDLdYEi2XNZZOb/RmT6MKiFl70KuNnoColckVaPIZLN4MdHvhD57XArDhrh
Km3SWZWM98EJskbun0W+Wfk+7RaOYxpnZ28DpOB/7yix2NbmliF3fnVQRiTI1M4D
+HMldxC5H2xx75cBtIX6dSwUu5zlfqwBRoUYlA747eg6YJ+ta8ZvPkn1TaEo3s09
NLCntbNaNvTDeHpdoHkdJHPNCvt1tiqD2cE856R6fdfCTrD/76gqyBt8S3JETakm
46wtBkg4car/Y1UtnazRsE42gckVekmyovD48ILK1HkDwYXmUlv60azjaH1+afvk
U5HWQdbo+2d1gRE3wMEXSMCjlEr9kQAry45tChy6lA82i/nzvo1rwToiPVbhqFRO
3jqghpeaoyVp9KUliNA7SoinqAHxk+Ojb+4FDxht4L7efFIPD9UBs2isntZu6CpT
vcYAg+KNgV3QCbOC+xFaWmqrjH8K7qnEZwYOaszTCsjBRbQQc2oiyiG4JA3+ZbtM
qd+u1ZXHv/Efu0gwk1El4pZOt1aCvNaaIg2s/UP+cxnrBYgAdc9ClXDvksRFmmLf
S8z9udIAs1tNu40coPKJsHowByB0tetXI+TeGtEMljGcSADFpmRK8dPHH+UuBX23
LQnczf9Sve9Ni8uvB9BOYwwR8n+HJxbOHw7eitrYUkY1imEQJLkJFZP3Je/uTaHe
16j/dHT4jYgDgE4Cm9CQwJt9awLorDbF8Fsd6LphxK7Vt+zvspUBYkQcAD9rJGvo
5OGnwrz3zQZJdkf59ZywRiOp5eHomJlz/TQHIOh4gFTlV8TDBHg7Uz6MBgVfg3Nl
UM1Xm9pQ+qySL9XZRqZyNIBGIuPf0q1lILQMdYODOjUN4boAX8VgT+36q2Qo6/57
4GkZduXAaBd9I+IJorMIGrhDmc2NlYDDAvTFvzeqFe3g6EYtxqDlW+6Ksrar7w8a
Dki1rcczwEoIZ0H/B7FkoIRpLGJwRpJa6Ubhx6HlYPm0oZVmUtQN9FEZJTBJEDBx
teYLFFhBdxISli+qpykC33lrqJ9oHIoBXcs8DBNFGdNRVj7T48Ij/NDMEOuWMqR/
fFBqG5bF51rXjzAEtCUl3gHM3bI8Pq4Bi/lphcC7L3aKTyfBr5O042Mcr8lW/rCY
epwnYOZYZ8hf3+K5Etsk+WSVYvGGLOZeKOLF6GYRVyOzg/amqEOsDGGauAPmugIx
qd6yzTEOJTny5MYwyeMRExf8AW2y3NenOAadvEGYuKXAtjMtgMts0fDn/bXCjWgs
ir708GZcj163lAc1MdBOOG6W1Cx0ZRVZ7oYIPCKsOffCjB3fh/T9dt+fhGJFikui
H26ngaqHklgjgfhnhq6glGef7XzMMtpE1BADek33hLF2K3AMURg/2jDjcUdbPAXm
YF8Lc53jkEtcTu5ia3hmdCMR2t44sF9ZijEr1T5I5DeRwNH4KRfByZCICFeSrSbr
Bpbi20YBNOcaCY++1uATvmwXSS6zHunZTX38xXXXj1SPGBFWep50J+WON9Hyklh9
KT/rMZi5Vk+UZ4n9m3cMs2UYex4h1NhHQbm+hGenFc5b331NTxpTHRwobbacnA0g
9GX9jHCY+8M3LvL+gkYHGNdNIxsLj/cu5IpODQJFkkvoO5wOl5Ys4nFOt1jKQJUW
q0ORkVUrKCPOoRDJRyZ4O8QqjMQfBrx5kwQbztos4kAESK18nYw6nReWks/B6BLj
++HH1ajSd2ZgG8ycvD/7NMSqIpSgCkaZxcGpqsFiTlyoI4NoQJi+XwdpSiNyfVBK
otATPKz7M5PgIQaWbYVlE/OAqjVJrL1QsCZyjDiUDXhHArXrSlTAqu7Dd7VYGvKX
lYPwnNg0yM6LRQDXUSukutMCoSqoBduHR6Nwzz409jPjXCcQbHPB+lV0D+G+ac+K
sPsLGaeTGmx6ObhZbH8pXEUFAx2YHsGgRhNo9e8EQEsNmxC8TQi+rGhuZRhkdl0c
FEjQ7g0BpLzCDBZNx+HTJU51MswRcN5NvhHXwGVqriDuT2J7vBvgsaoEyegD28GE
NXdOaLMF28sizfQb1hwQZjunnbeGfWDP885H7WaBBZyaJrgomB/r5f0N7nkFx7Pk
x8ly7+zHxlPv7ZIMFoNwczYOcOFeStVtS4daeKsOirMPlQPspYqBceu6W1gDvZu+
G/JXxkM38PR8nZN4BGsboAdsBi9tZRBlgq6Gz9Q8C73nM0jzEYzn7q5WbRUEIwxY
ll0xbdoNDh46n+J/wAKAA/oMl5mns2E6VfW+E5OoZYmMgB2EAx5aXA/1fjTtVObF
o6qHXjwRiux0g+5jd8TQMr+z9mpWYXqH6wbFDWBXJnd+H5yPcS0LZlD8i989bjkI
tUxP/SVR5tEwvuM3wsp0Vkw7Ommg6KMiwS2AoreSNEOjNMLCcB7HqVJdv6+jgL3T
oMr16SjHLo7RBL2JdRqFs8TFF8IVPylDxL5xXPz1zsIEQUzx5zxOWABr8KPUa1Q0
bg6uzl5CDkin0gmesVwbwjLog520Ab03do4xFX/lQAu+epLpH0ZHnxyxOYjdGBa8
2loGcTAPAxVGRWK1zsavZj7Ynirr73bUdPuY1XD5QKjeK1OT96A5+bDq1GJn5DaG
abe/lKhYjgx5oQPtd2A3y7AQNIZmGQPnYlgramlt4ML7mazgJsFSvqvkSEgqAdZt
xUQ18b15icviy0JkzyHuaR//5hsDHA5CoEahkn3Q6m5S8XNtCE0uRioshaitFqux
05Pz0u7KEIZ9NCq+WJA7Cew/ZD/u2uVtARuskiM44kC9wNEs/q9IPQ/FT/wwpvIz
S/OoNHYX79L5FH/vxenAFb4z3mZfzgrProcB/MXFmYh9t5vkGO2xDzMV3VdH5ko1
cNFyC3yrWISzXTOzcHyjahvkmvXu+nc4RZD4Rjs7ckUfDrPxedLYBRM2ibtHK/zX
Z0GnDW8UBjWe0f6yHKshLw5h4nqHR24vpgOxxJMKRqtukhUWhr9PkXjS9nFlxAvU
M2fmA/KfwdV4rjqHaZVWvQDmzxNLrHaUO+aTnQXKc0smcpB+ChGgYTsRCdVkCZ7s
aO1ECnfaXjExIe50bsK04RK+xInLCmXoLcVIsDmAUuTYhL1up0wN0I+tcLYWuiPZ
cSVK7SaSNNBPFqGkvv/71j2mWbA+7oXzTKwvOGH+rHZVOD1u1osgNLcW62fAnZm8
950HBdSnHZCjXUHndruEAdtkjeHM1zJjgNu9n31QDoyz6POSpuxIBWSZ/UL0JlwI
aRBQUjBFsPGG/DPNrCyQxgCnMSU9iPKWZ6ygheGJ8rMj2mGu7M8E8xdLh2sa7wq9
HLqozi+xxp2qwzeGeVlnd++5G7dcsxTyNKIAA2/XD/h+HF/Ou3Ob0u4aPYfIIUJJ
A1L7teFL2BqMrOyiCTBrur116xu/OLa4CfrLc38sdiyKzMkuyGKaEYR+CVOHa9m9
25V+Jwmd4zv4vM0GtC9DhCV81y5A+q/nhVNdLDI4gTJMUMoD7AYY26cG/XeC037o
4UuR2Uzlyc5DkGWyzJSjKp28bxNQ1H3GsrqyZK5r1iuYDon1XWt/U6xpzvQk+7sQ
yQ7ptq1e2EO+D0k3LNXbxnRD0yV2+GEBR4ZXfoC47CQKFsjYJBNxYn4LPI9EzcLA
sBd8uGlTbmntpq40W6Qvq3V7a4sLKCRfuOgz6/AmlZb+eDAcGRjN/x4AaBBG2WPu
dCXKvWz8k+pT0VpIHz+8TrCxLC9GWR75rv/poC+N0rezw2eUO++A3FM2ygRBANaq
hVOMjj+587fHT1JBa3q4ZN4dTH3MAdUGM9FSYnTVBd94N48UhsZtLQAShsVwn8A5
XFjX/2XZ63F8nL0pTZBMZ4fBlkOQgBoMqkOXls0GCze3l+tlqyop3LZ4jb0oM9Np
0ZBuQcs00eha+6ainFcP5zknyh5ccXc3f8SDhuWW5TipyJ+TcXZMCuNqcrPsiXZY
2lVKlbkE7fL1DgZiuL6gG6IcvUL8XvZu9SK+dADBa6FgQczWCQMLH2EyDj15E4vs
0jkxtSHhV0S4ZIkYDcwONbjrHrg6AkAiU7hf/Ou7VmCOLb/QN76qqttEiPseKmbO
7HiVSOczSn54Gf1UI2clkUG627MovYwZUcATWybEEp3AEmw9GlPPKt1dUdvq0lw3
73vve8/7nt38Zjmj7aYCuaViCBsxuyPjH5jv7UwwbhApE8v4hovUQqkd28ivLLpV
8IKmhaXMxuU6GBz8RUp76KsJVCmORWbdfGMap50m0y5AdoBdD/3b3+PPQV8TiTey
QK6s+l8rvehmTXMftUZ5xYJ+gkyDWg7Iu0Amn24X03gXO+qLBaG2sZs4Dnpob0FF
WWdyaC5kV0PxC8P0aT9NzeT7d1a5SXweswAVf3tT23auzMf2MXa8EuWg8KF8GROU
r/YBIgrWxO0lNJdPCG56Tf2/O4fenZpu7M2PCDSB4Y52FNRhGE4kl0In9XKNZAMM
FWXlYQBrkMSrj78WjcIQgMbk4RQxiv/GpuBhcC3HwxIDuGIPWvmXhdWlmlxC1h5y
2QncdFM/+5l3s3K+AmK9qRMJQcJaULy94Z/1j7PuaSIDvev5UZyqbypaR1asBnD/
VVYNEIWUc8r5r5U0GwQtj9C32wpd1CqDEvCVzjNI5KS/j3tcmU+G47EAKPVcvvJA
5BUp8KXTrSZpHm5UGrS7LprwVnDPhIzAt2mOZiE0WP7uMQWEnucEXf3I4wrI8NdP
JdBCxkrEznU2jIecpzD1VQ4uZJ3jcobbZuFylDvdY45WlcNcToch/P88ojJJUoNw
EXU7Hih2XlmejT4Y7cqK8i5NWemJ88ZS5YJAHe77cH5jKBVdbzcKNjd2y/gU9aTn
7nue47Tmlvx+NPq3ln10DBdxPtt6I9sxmbyjkH8X/cqUGRJJFsE+KTKGDdi5EDZB
BEWerfDOMJvovuYc/ZVvxgZyH3283Bok5qtxedcrKmz/VYrXRXLXiHzc+VWp0Egt
/EIQy1M8WDLwOXtXuBgXcbvo2R/EkG3Hk0MB/8K8uZxSQEUDiGnio1S4x23lUwGr
PcYsa/MJshlGM1QiwmHBQ2R6dF+3nzQktKhJ8J8LtENefn4yxdmixZf34fUGGg+B
bpccV0fGLjt1eoawFW3CQ2Z37AYwC3LuDkU3Mw/pf2kObOSAT7prq5eX8fZpUzRa
aSZdjuKNWAlKSnhezo2kDy/aM9UkVsHF+cU8D+oUSrMUKcMF/5hV2Thu/ZwY4sDm
eNYTdQL2BBgfDBYachQD4d2XUoYi+9loHny6dxKTFzf1MA0e2JULhd83HR/isg9x
QaOwWxV8nRo0aiBSgEOBfqGdFut4RuDGNW6VpOpzjNAi8cvyllpsnTF6LvBAAd/B
50dBBA/xUwy5FO/CqLFkDYK/PurYa/SGtI7QXewmjFw31N9jk+pqIExvkVwBc3cN
HQdeV9DKi6IM1qYsolvQ4WuoGwjBbaJ9kCosv6PPev3jJxUmgInaSxnMGtRvy1oF
hqz33ZrDLEMvtSHfFVGsG1fCFHXKmF2Gb4GPQ3Wq02ntpjX3Ly+s4NcKoksxpIBg
bTKJEUNnlHDijLT/nFfgiAqBNyIufmwvUZubMLfD7U7h1TjBNoTEFeVqRRlxQwWo
T/yl2NVwEYPJbjl874uTEnTDi59QM7wa4voFjk8LmSXStE5Yty13J/3i1m1QXVY9
ARpHzZnh8hC1Ga0Cacqx7DtNiNtMdFyRBkJFEID4j+nhuXEPBQznBE8PLBinWAHZ
8TuZg1w+5Led2d/GPZxxzEUYOCuoMTYVWhgx/mSomQVjiGe1sMxka8wIMZG+mbtu
0JtoHu5Lkts3zIG/PGP2M9yH7A9q7kEOEPaD68JH0fIgchLbH0xQard2fnsirDqz
DN0eC7CqtBqYJWj0ZvJRrHqEVguLZ2Kblx8/EM0O5bz+jyaPICwlAmwU/rMC0ty6
D9Zw/6IdNvC+WXf7PIEoZVn2Z/i+yT3cgKsCkVjp0KHaaoyPRp6wOPeI98M6Ox8r
KG8O9/naJGZoIWke1Tht3XJSJXVuQ7YI8eE8b3C/hpjq63P74h2ap4wwjGoXYLpG
2tg2jwgkoP2nsHh2e2pyCBBHTOGWXNBQDXwPq0ja84jS7oBqEdhoIDkxvv7mphX+
R6dVWnVzhLC2b5Kcc21vlcjOmD1WVWEcWXzc2E4+YGKJFHzn2qzJcvcP88/t+BDH
g17c1vV81zA2rwxthZPIrEj6ohHpIE6fMi1Eg1d0r+dlC7hrFlftl2W4HBi4PhVg
1GZYug/KORV+IT91rq9rxCONZQH04XgCpRTsDc3xLPO96/iTn1LIo4jhFPAqcXnI
xHMY0NEmzS6Frk29YRgEC49fAx2l2k1uCMEkc9jA1XzR57wiGWbmA43mVUvMvFnN
PrihIuuCb/jPvHm5H0StBPHnKD48w7PHhHFPminyp8hn5B07RbpTHncaOKjKFBf+
FWt/teEr32Hqfqy/MuUbeWu21LT/XFixT4W03Nx4jan35sQzumzEwjzAnNz0CKXh
onyw9LlvgAQ8M6Iu5Dn0Jyj4cN/GC1hptktb720JFkjVil8djJbqaOOO94M1G/IE
gpoVzenuZIS5jVlD6chkb7TDx444khrV+ACtT/Tgd0oS/wF3og5y72NeykMNQhoq
SwizqjXn95hTmT7/5uPkQK5pqha1jij4TG1HYYwp5/gRmAIPYhCi+dKeeBoOF4cn
CnRUOQQych05OrVP9YAri+BFT+5M72u4UoMf3xbQUT8ByWKud+UNZfvyp8r68hdf
jKjgdG55UCkAmYxyOrk27YIThdzf85WTi/rGTy/1l0iW5digjTWbjS618TMON9X2
5skc6GlrOue1hUwLRJzBRFdktmckHfGu0egjJQ6O3VqO7o6LnFsxy06lDEGdZ95H
HtIYoBzMaTHhwjTCoY02C3ulK+CwcA7O5LFambwYqAkeYLEYkiQafN3oWkNzcdk+
AFNuKqXJXoPDVhrpm8ML4FqoZg4DWybmSY5vWkpyYUxVG+cICysRzo78aLIc3u+k
8l9D7qvUCJk53Z9TU4cTeD8huD37MyZrOul5SQ4LH7f5E517iecjgsDLcvzenVsj
NDiLi026GUDcRGNa7KSongZbwck2W/tbSn9iNHmcmzbCgc5gwGkBNwGHYsWLqUWQ
8EX2HahPCZ6NF52gl1H5ajrO5feB4dKeBKaa4Rd0D7QkQefdLObJm7dzxyZli7JP
0iw2AnCSc3+LKFA9DTrznAy5DWyA4px5jPFLQfm2/+QBH74a4rtZJd9KCP1AyWNI
nF96szCUMf1DDNDvPT47JMB0vuN/qEVQp04dAG55ZZ0nauSYigCVPX/T8bidUKQD
Y6Mv6A1aTvJ+Oc6Cxr8Cln2IWFbncm0cYTn1QHMSQiflZvzef8Uhq2TqqnKVzwFa
PA/yi5Xx/UucLZdeh4AKxsoj9rq8VyONn+672uKzhWVQMsyV1j1SoTVINgpoQbfA
E+WNYmeU9eHPYSIguBqI6MIZfdksh074yqCeNJoQGSKwildcT686fOVd96GmWphJ
FgixzM9ryzO4XUYEjcLBd7dxoAZcVvDAP1nVCCG107r88d1tFtVfEIpbtBE0EBfg
VKZSAEa5yJj4RdLBK39EOXoWuLKnxSdm6tVmDN4a2zmL5B0wCR+N4BE9c3g5Z08N
VHTDuvj+s29V7Z0GB7MfYscCh2ssTfSCnl1LOUgDk063S0aP8EkM6Swx4N913cvv
aoFfoo6vvGVoWg1g+GTU0dDo5aF8Fd4ikB/jEu40Xip6SQxe9kM29WVLsVyQE1oS
ti22mM8P4qcdXC3pKesk4zb97zWJFmSmNmrsPMJO8afmyPr/835s9B4kYXWIRz9w
fZjSPPssk7nqRGRtEcA0vp1N0vckOku5N1XHtzEm/buiCc0ixoUKK9n4OZfNP7E/
IGlhLsUBRjHWy64F5fQOh9FYhldhb7mp3CWtBm/OC8XU03TOdE/mLN6rrZJJkXeq
OI37DFNRSGtQCZ5LDvb+WA3Q1zfb+LPaeOBzrmjdqsEt8TV6DvrYe5Pv/87fisoB
St/ZYygj4WbFDJOtHsLQWkD4iGWt8rtjNlB1QC5dfIOc1d8RMXtkCajs/uMvMEmC
kdwigsdJ1xFXn7rbIN1OERgH7isR88lOdNsqtakMvPM1HfWDq/yQx51BlOYQdUub
LOqrYhbCi2aObAalqCH+YOCU7gEDwkkV9B11TmGm7TMeu5lUXNbH34haV0SiE4A3
K4BLMMeQFFfGX9OnMo4t1RowNXuczj5S4w//YOxMxSR+uEPTKtFCZz84+RBXXa/G
lpDjK8In/xbcA8i2hdmKKUPUpzbUN8eNNKSxxrXKe36Tpe9k6AwnYHthfrseCPJ4
ulwarMXfEjsGAuY3QBuJjToxvteSOzp5yupvYSwEeMrnl5tMGNrI7tT1QOvJADEy
c+SrKNddVZO4Z+hSWEUGvxRJpwJmjZfjH1Bdy48DEJeTvFHxZlxW2wWsdB/4lgJ0
abstRUP6okisGFZ1Dl7KytbjpnxFK4vSrJaMrEoInWTJ6WgTX5xJatwyuzTja7O9
egGRi7cfOY+8DrOXMSZLkKWstIN9r9Vg3Fg2TBCqFKSGmmBQfCmMTxD2AKgZevrz
aqf9xut0/Q/IgLXYqc6ocrWcaWqIH5GIirnI3dqr9u6C7jdA4PZmE+UG4nZWZXhF
mYJ86EBkcDXw0kSZPbOQr8l8b+uIiHUHaq0l1yAUeGzrgMhrrVx3CKlPO0XW0YKW
HEsPZTJEF7LvDfEQHCso6jUa/J4fYsAACZsjpu5lCspjWjNrZlZ6kl5q6ACexipr
irOnHSMyOsPbjWEUmdUVjZssnpbttk/fUmUrynvRw07cgViHX6oWCHcg7E4ASq7d
NT7AA5ucWDrUO2iFBwNw2UJ++2w7b569Qaauf8nbkFeKNfIo0rroj4+4Bc6JM4ie
n+EHSa5JpbgehgSlNHj+JZc8qUpiFo0XVknOgv6QoBMTlSFCVHTtJqb1rYzakt85
P5+ttFVWXIGkvQw6BiJQTPWEjsTRwxG8sJ5UawRXO2x0DYQX7qji6wCU1CeDs2Ec
Mj9Q3/CneM6qaYF1AO77dkwsw7gNRcokL61DtWHnxvFE9VdJKLWWi1TZUVghpu09
LrMK8SlxbFGKFBLU03ANSEPUv1JlPxsxiBqyGAyfWloqdtXKW0I/7Dq5ZLTvtaIa
dK9RIbTqjlqT7PR8T3Z+Ny1ERRtGSvYIplnNti6fZByU80xgoaPL2adESimlwi+N
wloNo2Np/fOxPrF8qM4Z881X2Ia/JWzx9lRl+LZCz9dx74rtgNq0z/qBEdGRRarg
pK25wH/leyMPGk8U7ec4satxnfx0AZyr/dNiWGzFejkPDqv0sHBkKS9shhhKpODN
tVRq1MwNBslaPRNFWwSiI+sAJH/nkkbcsrzSzgDf9YV6neRdDtKdPRNujYX3XRyA
Bnf1IIYjqFbSBIivc2BuLrA/0zjDIFUeP9tDHh0L9/dAYDRvhwCvhQ4Oah06U8ut
j56GXjPfKrGjBqA6LZOIdTxESxYrYuNLJfI/m9T2WSiFlunRv/Oq6ezrgT6wBXYt
hxkPkO0E63+Ji9XYJfLGVu33yOK0wzoy45WwPsSvmpC//vYYgj+mPs++3xtdLScH
DmmoXSq81P+V4yuRvcogmRd3SeSJ62P9jVm2v6YVkZvBN1VbVbAYDOMcJzJKjeje
opZuZLQ/2mxmlaZfEr6zVO5LRsDPQob70ikvUf4dEb5wmZxtnaKP6idsZyAoUjeL
t2qXJ9xZP9xiJBxShQ80854rtYUNMkOYo0SwzxrkyT5I6a5KdwtxK6irCticFTJy
ifv8S2x/z6mUnEqqyHSqRPlLhHbkXsVdM65x+s5m3pYJLcmjEcXA+Ia+ZyRiIbsh
A5QJJCW5RDQYYfyKLWPCm+o364Dlg178CfZLGDX8A4bH5StKlmBMqn+d1tBFXjr9
oZR94nIxF2ZDqIhVOMo1xCeKaZi9VYiU4yXd3D/cAWrn5mfFuNyTsNbIxHlT3Aab
v4uJFCuO8sJU+j/DpC9nrc51BLvDMeQOAAeDxMGxHdF/h16bnybYsG1jy/eE0qLB
MJiP3JcciW+QYBzA5J0vSoK73aM/9/P9cYxB9m+N2n58Eph5vV14tMWL2rimKWhG
HWOsGZX0Qv+WQBuusx/kGX0wvma1FbZ9hY+jwtUJTY1b8OKOWly/5xqVg2zqdUWW
EJuMvo0fj5RtdLkha5PHkTO25CzzQSUbTVH9KS4WeHhl9n8y1wwG7OCDC0Ijdi+J
Ueh7rdamwG26LnqQSPGhflzu8ub6WvP8abHQFMW+bjJxI3Vsj6d4dT/tETbyk8mb
+8C+Bay0f3lowNHGj4G9TCpjI4PZYH4ETxUyj3hNA8GGIzGNh4+gRRfKXEtaOsPB
gDVf2wuOZTr+C/B8UkI0b+stNdYAcrN4IUgofDV/vQayYOt6uT00ZGB6Sw4J2k+r
bwX0ZrKZEzv5z7C1FC2aGRqUQSKHOOfa5FIzUW9dhBfExKZjMWcXAvp212yt8k2e
8Xdlz2o9NZpnZhioZO9bgNqLgK6tAf0ooNO3qAXimailY2fzE7NEEoz4APp+RPac
W+/vlcpvjUT3rw4gkscRx5zFRfJQdO7t1alAxKj8sq3ru0bfDXVE+cVNGKGjcNh2
3hjFdPf+qGh5gQA8K3zthBge85m5NL8o8PEkDakPSIOlz8KZxrvcgJFWOGEuFel7
Cjpt/a1BWt8HkzYYBhJX2ftg8Hq5NSXSblC5oTAXFTjzyUBAfGq9oImD0UGtXGBo
x7Ya/+tUMNtyJNjt6bo5PcaBR4iCBr1F/svVwEDFfMCmsOmdI8J/M4z7LdaBkHUp
R8rPFnKQM6/9l/wLxX7hmdxrNQ5rKClSHfh12n/JIjEVGO/12gu373YpLSnSTXg7
p1A1IWLaZFkUNFwt8Q+9je7g/aYDY6nZHVj3h2EZRhYn91rgp/zlZBVM0a3+Gu2W
Iix5l9s+3D9JlemMlq22ZTCRJ+eu+Ns4dX8YGQZwuo1523JmAo5RxM2F6jZSBWDF
YBIt+lwamQFl51wtWGGkWuUYqwuI3VoDdfif+X/ndOXnyZYv4ft7vT+6+dz8bOx5
dI6SeQUIVBRKYmtZGkIWHYMGqXu0Q+rcQp4+OeJ5J2Vw1ak5ghLjdhlHRGPjevWN
RFcD7dWXAXUx8C+eUFdz7E87/pRYea5DImPvU7DU+o5oYLt8/l+R9KsE/eev481x
5Ag5UyfR3ar8xR67deOYpUcbXcfAnPqOCJIxOJwi4OzBDMArWJUwfKeIgtbVDUWR
VHyWnniDOtYOzcnJYmL3OpiMvLjAiKf8Hb225wL1niSHMpHeSM+3DL7086ZoUx8q
4dv+GCnm1RiyA3krmsEr6DJywCh2jjiOOOlvCOTES3pcOJK6lJiaiKTAPqLdWCt3
/eBXMIFnqw9c0K9rXr1UmWlrFFGhVF6OcF+kCdcg3fvRvF43t4lKvJNISk8A61Cf
/+feS9RyTd/k9qQg+nzEn5ry3P9cze+1ESf4qshUsqYhsseqs6zUA2UO24qPwEBD
Jssm9xBJctFv3slrgaCRcHsQte9giAosz6kZ8BX0fNvwEDAytbIzTTfo92p+NL0v
AZGx91OXKdL0SYnERBVJRd/CdVLL5MTpZAWylmudgRtjRingu+AklZ2A8mMHIDQg
SIPPxINlF6blghE0htOQSbBTTkGQCxhKD1qlk9yfHUFM22aMHrsubi9qqPH6whqd
THM0y8OFTTlttv07jxIRbhxbyZ8Vjgk/UPsCt7Ugx2FncG4vMOr4ebIfQoUT1ZQP
kdeXXn+0BmumdhcM9F085sjwAbUEjTVcxqTd7MXswfNGQp9jEXImLW+eyeD/kuKS
D+V/dSoTkmcwlbFA5DRKlEHbV3avotLKq2B2yLV+uGKue16YR7a9tfyrqYPpzfWq
6BIrWrpJISW140gkPRKQAGWGPLvwrqpy9ddWxNgxGSPTXIhDn+X21MYiFWTuuJUI
O4+EE+YIXVxGbH8iQpJKuhQv4tBvQLInmOUwkf9Gd4SJxwXv5RCAR1VQmqrulpJ6
Mkx57Td3OD07jy1ZLYzcgnjQq9DAtz6cLC5QqU7WS6aFW8kvh36wwCBhnAH4M898
tIV6ue4vFFymLIJRObbPci/Dvt7rYnMwFRv8aOf6YL2BCloqJlAANnLAq6ZdZ50d
93/GPBqLwlA10hkECuUByOUB42aM5J3G84w1cYqEYdAVxwim07XrgA3JPD2hC71A
lIRfkJhDYqw6SkvBS15f5h8fTzYpJ2u+Hg7Y9H5hXYqFDZtozoTeXVhQhtOUZgV/
uSOs2yh3XDeEvv2s8NTIiXFEn7CVVvcJf7oSPJT8gQPvBiGPzSF08ks7E7Wz5Q8I
pMY6h7mpfRuPdTFiya288BRC2MTLXFDm73sjTYXnh+NTTwa1+uBVlRS+VgVfjl7p
E3qn5XrNksCAC08L1uhovDTLffkaBlhuhPqEX0YOMxmxSIbNH0uBChiyo5GUTbNp
uWMNYJf9dfUuRjWxwRon2eVSjjC9wN5f2do1cmZXFu8xSTCXnX15SBCXanBR6vR8
WOszejhXOGx4kVVb7sJM5QqRL1nkfsHX0W4W25il4rUQczLF1I67/8DwFSbxggcT
Cw6Rug5Wp58oZ3NnSBpXCa52iIxYgCAudEj3pXXtAYjpWmvQ7VI5cnTF9s/+q5cV
EX4dREYdHeekpwFUPw81DiypVfSZdqIXhi5HJVcL8rVxHT9+kmcP4dr9GIa8GrK3
ZRu8Kssnq3LjbIiR7IV8M4M/bhMNUtcXp9vIHYy+ept4mNzN7OaPQ509iQLhNcgI
jT9K+XYNEbGIBVRnYMfvfr8qdMu9d7XMc0Go+9vrb0/Tpjo6tC2FITlLreB6oMpc
SKgKMbQ8ir+mHutVXgAeeqFeA2iPP/aB7CmmLMl7zgYoMzhwYV8aLkLbBtylOutB
NnYu7oYMZsYqtsBfpqVy9PkMTr5oORL10K47SBoyYZUE02mjc1TdKVDu1qBXyvQK
OgT7IazbK4JFic9IUkGay+ixHxU31R1K53HLP6TZh/RLEK81YjUoFDprINk3VkAn
wxpWBYCNut6MPaSGNDmrLuaySFeGU5Laqb32BSfiN++9Llazoe9rEe+a6fDW3vaT
gHiPm6kIkd2ST87EC2qQsOQxn6EDtX/YpVgMN3EW7eF0PFWtU9CsSnzrfoY+Qdyl
zO3AW9LJ+MHWQgwb7tBxAHpspVRdS3vTeJUsGsMdAItUxnqenBWl1LdMrBDRqUzC
/mQxOl+GszAEh3TKX2kUx+AYhWPjFKuMxROwWxKKcnddBib7ErAy2kz/tocUJFH0
9XILJs4VdfWPr6HGooEY9d4Yb9yuD6Ek7stlzkX609ndbY4kBso4X4aJBjpbwOLG
xhhukj8GhHT6/mC2+4QQb/Auj8PLhc3emCIHbIWUgCs/Sqt3CxKPDcUdt1ob7FRn
yCV301hOXRjZ9Kwg6Dj9BqycmAjGJ+FOAve5/Jxx/mahnvtS+MurFmd4YV26Jxqi
eGJzZP5N1rrEKyMLngZVpupy4cDxMx0x9xs3vUMxYwJ5ghZnWJa3Ng9YuWoMHKfm
WxXoAr9x9ikwt6DdKnqZ6NHDV38iW93JuRVJoLYHek7CVy91pPCvVmllmnvGa1WZ
3Zffy9QddS4LOznZtY90MhqdYRggaSZhfrjYBEJ0IPt8txhMiB9PQvD/aVa13lMX
8fX2y9xCdbBIHpA36JqMEUpCv+WDF9nLRic6MJxokUkGHEJuG8Q7f1PsSLBEQXCZ
XzcL1EyXGEclpywTe57V8eiO6z0KXupR+jYu63wuoJAWx0XvZ5I5FwSmEo2QD04F
AH/yO9DyMroyorEJ6rT6R0QANl6mh92G9AHRHqheZW06dndgLGiS9nbYiPtHaPaU
m5aKmw+YYzA3yATgSVinEy/N7m/IzIa6nV+raDyh31ms/LQrYvB8jzHnGpEpcFP9
rWWjXsA8PYdLhoXamWwN2HPf108abdGntYpRHqqa4giAVfes1TBWuvCmOSi+71Iz
yFUjf/4fVx5FcAKWsXbCRev99zDZWq0KoFNDo0w0yMUFa97nfuzGkg+kHU/z2J2q
s2gISw6MNlCbpxKK24lTtFKcLmT17Q9b14N3PPA65+/4s1CecINk/SC07AJgVhTm
aPRup1O1fpUc05baeRBlydwwVy/1WbtN6k1CgcAgRAIVixOPOYOk5GMLgkoXamHG
V6p+lXA4sMytYEgDF4CyiCcS9lDHw185dZzgahlBGM9eD+B+qGwnogOG8+DKKAxN
7SJIWa1N43p5VAyKufo8U0w1GlbE0KAIDZDD+bIuRx/cTmtHhAhKIdIZoDrFrZrH
L/d37H0fjqDh+SNaRacvqqQbjmi56x/WN2LzKraWabBdmbyUYfYDxHM80l6nqKyG
EDDyUDEde6gHSX5WE+8cUoZrQw0eddcf2+N1RA/IZ+6QiDTAPkJyz+xHouauKSDA
qnZ0tPkquIEdzVexjKjTmulILAPxy8tmYV7niKdeSVHJKLlfWm+XMhRsg8rzLDWy
iIx2ZLpasaDwebnClEWMpNO8TfXFtUvgMl1YgCrtfAWBFzgrG3fwgIOgPAkZO92Q
LNHwATuiCcXXl1dn8sUdl8lgMZXEgJpRw+SsV2lWNo1EuqR6oqjXMayQ9SUDYB/J
yGLwp8EIx7j1lVZnp6ejzmnk/myyPGAXASrXnEg8eWqjFkqIeEw5vGcmv+odirfQ
aEXUpsD8ceLTpRB62rm2XEOVDXJZBS7V4lhvpI6FyVe7Fb6uV7GKOPrJ6Bpphwi1
8Xer9fGFUIagvYWU5iyR9MNOU4CmsWalGOj19BxU7rSJbtlq9bI8ngrp/1ZzXmRb
v+k8gTV2EafHouHV7YNGSVr95cvoci9CFemxWLCziVu2oC6bMN/KR3bBbV9H5Tom
8g6iLk7RPyKf3Z5oi1TiOl8TzinFGL5v7YKkVveRjYy2++743rhywa33JaObXy3J
IW3qZPnrbeQ7cUZgOgPU7/QpJjOrSeYYBRJMRfEgyvxBd81lrq9gOFXDgIexzKFG
iyoEPmfFAcy5Oun3cgJU2oVOwlmq2MLKNeOpsTo7A9Y0dVW1jYRCFuXiIWypPvNS
uR7FpDR4q2Az+p5Dy7yEUkkArWfLj6kQG4yi7xoMG93Y1wVLdbQuw3wJ/EDY5Pbp
e6oWlsi/dCPcvrDX4/whygwuhASL98t+DpfKJZixrP//pBmUgh1wTMgl2TntulXA
yz7cVSwreNIoLvZEo4ZgJriDc8o/ariBqXqkIWqHckGfH/F1TcwNgs/UGCAC12M3
zWdqnfuesFLWQvMchneAko5QcGlD9hzD9lX8LX1IseHM0kaQsAwWa3xhBp4fvYHC
eJ0IJllGQK/QBqiDTomVoPdB8ZoMBoc/iB4NeRGtMaiETkSyU+e61XQI+Ic6puM8
nMo2a881WJVBN7uoaP+m/irvU3NP231fyt7kZ2t82adipXynHghp2MnO6uvjoTXn
xLUz/um6u1JeGviPg3Gwb0A55fdLUz3gxOhu9y6oFszaKlJLpQUnJIR9PmadBtoa
DvJA9QxN6KYqsPyiwOG4gRqX/WobNHrF0PSqmXSdFzvnBkKrZ/WJwoTB8DUifGHL
SIqHPT8+fPBN2JNmZ6Sp0XlAnKvMoekkBsjVgNn+P5jMNTb47UemCYg71LAbs+7T
3FbzDx4qBt7fITqdWWOHTlq4I2ZD7UT6e95SK/o3JtQDenLLV3bbakGQJZUlMDL0
FOYSUga+AdyEZHiMaQJ3Ore3S74gkhmQn+Kp0rCQLM8xbBoyg7PVE/sbqG7hP8FR
CPUNkNHCjOv0IEtTXmYWOdWp3dBTttQmQeLON9PRQtiA3KTlj0E0/UTAH9PCWUqa
l7tK9/TAaJNtblgiKa7dA5UP1lhhMwlFxfihzzZAx24nP+NKDl7c599YNhjctMDm
b96h4v9G4GzQhYh5hPzApP9UkeCgGLmEqY2kLKEVVxR9XpuAJArZnlwpSljpkLPg
Komvrmkf5Tg2wHXDTLdq+iu7ERp1i98moyIMeUrItRsJItBWZhtAIS5YzQKTuD+S
kTWogTDOFviprssiBZ9wPmKZG9xJh+xWIMwrb9J+NhITOaaHa4j9ARw7anliCfud
b3xJ+Umdzn6l8NcP1FTMVr34Ov6ZL1Sz3lVxO1b3XJIK4vqbqJNX6i+LPrkeFjgg
KS8/Rc7ev9jx2W3R7Ixh2IlFc7Si+l6kz4r9h1GVg3lAbVzZDSL45bnfotwufWss
46cqvJ+C3uhu+XP/6QfzDSxcRwMEwePJFvCDe18L/0sDG5j9hAwDve7ukEvo3kgI
L0DUOSQw5M/q2coX9/U9WJ7ph6HRgGfh1L2TTkJ1lB47zonVTRLtS8h7vpyF3LD1
DxGV519fq4w6Rpx+XKxoO+q84cCRHze5WimViVNP82WIMj61ZoOX6Vk2NJyYRVdM
AH8IcwpN7q5DnDV9IlMuGZsmjDWTop++whjYHx7axiD7jBrC8ZHUyZc0Gt5ZPAZZ
DAVxxO+YiINOCQWyIAsFw4CG/NrxhfKrpoYtlX4fJttAhvpHfN9rGc3NLJwZ0X8u
43Kah12F2v1R++OKyWDlQahBZ4IkFr143em/SxcX9q9xhjYwBVeJWWiOY4iV4G58
NvnytHGO124Aw6vpbXQAm3IhxcIZUxKqnuRezMGgdEp4WMij0VrnXotjo+JWiVne
kCaKstqv9vl9tL2Rku8jetzVtW7KmmkaCQu7zZs4VpbxSpUebEAN/mwbhyMfSga3
ItYblqCd5I7YVDX+0Efzj30noTa6mDRi6c1QoYayJfv70XS4O4nlIsMP+hN0Fm4b
L1DNUig+PPPAcAkZliH5ilxI07aJqTFejbX+G5MNiRu0by4iGZ5tlKJ++wsgPGXk
8yKgNVk2sUKuxKJp6tUKCk9QoWj2i05XU9nFF4BR2Hyau85fy87KPZP8l2ovceBw
7Bsw8pgCPefydKqCPigRi3reYmCOPDtepIDEtbBzwnP6yr+Gm/qIu09WpfRtbZtp
nvpeLAh5N+oKd3bSTQ+y7URmiti1oiQBWT78duIMGOTxXw70/p8Zze1qx6OavPgu
52w+aQ4ymmSlDvDGX8FZ7JFqM7uYC0qIzqQA77G34epbVD9qngvG0KELOhWPMCqf
OxuVSQZeftJ8vKhGN27zv7EPwyWszhfFcHtO6QyPxuQChcx3njAS9ogzAXslYFEP
cPTwvJL9FTHYE+q63yUhr+HNScg8B+87Rx6pZExOXjEGBcBHVwC+3A3NLI1TyTJ2
IYwd7Wjndj1AxJ5X+3/OewXqbvU0L5OunbtdpdAvUxzFrf+DKuqArdgKuWKHiF5Q
pGABj8eDALDVgpBjFp004x0/NTT4qoByWwjKYCc29EI9MiTKS0TmXtA1/MqRbV27
hKai2vHZiM/DtHTZwwLclVJpaOg78zatdlsdymebTtC69a0clVTB/ngpjPPaQe1K
/sGAqPgxwUfkjh0MA3Opg2nh/o7kAeQyK71/7+mPLC6p/CfWUoTCP8h2ei73hZ/l
ZoVFs7lRgsoAnfn3UWgkyXRVegJ3dJ+e+1ECFxjZb0JlKJywoVhhqjEedmOwLx9M
S7RZ31uCKJdxfKT80vqgJaQTojPlUThtFPRAUieQJEaUF3h5jZ0ICRMj8Bv3TVIO
qZg88KhepDoMOcybknyw453ckUUgCDXeK7Kiis5nRznti3Z2DdsTJToOAJzhmE6r
p797yL3zy7pOmj11XAQW9hrEoxbqEjsRo2/xGoPVEXpZcW3jg/4ZBUF5HbtCHRds
806r5UYfsjCI6sYIS9h7rR88Nt0LbuEKxLuxKGSgk6sRhXYj6r570Klludku7htx
xbWpX9Q+K/8PGD89gpkpYscGCak9mEtJFnqxWT9UUVwyUCzHIOjtvLw3UC0y4mnS
w8GnfGcPpgrjHAO3EGZxSJq5tCCOj+kXN1w8qdqbzmj0RU+cTYkhq/nPuTuwlabx
gwIcbNey+N9dz6tpW8zeZLPqZV1ZoYg3bPnnYS2nUVPf09O32jfl/o1UzmUSicM5
CqjN/Xd6wu4Te2GILaS8e1PQSZ9ul5oaU1WKFoLatluAIqrPOTAV+7V+oCXSCtTY
9/Rv4iKX5RD+M10zBGVGuG3wHzaP39nmFAlWn6o090QyYo7kGNCOPNF5OP3a97vc
d9k4vVd14V79qUrKGIY0Aoy/adMlG88AcVXau3ell90HaskZax0Xc9t+hCxVpZsT
YlGJTNGb7xP9YCSeANtw0CuyuxCPUytVeiBzvv7Xj8TMz1ZBqUlPfZgVEYY6esJn
WL1FrAKkSJAE0iD8NScjo9dYLCiBgks8UzyRijyFIDigHnRXbjQSZeoGyfjOs0Nc
ACyvlfHiOU9LFYqjjzfwFxUvo8d9ZopBhx8MhMKvkgBIcTD0ouvQ+qKrr8CUaCaP
BNclykTZ7dLDIBwF6PMI1uzboEmNCJT+6A2GvhAR0byOskxx8AtfybsC4KJLmghj
zf3xPNi+uZT3cQOutKOCxpbPmjrD9mZXQBhBEpHj/BEM69Sk9ukt+YGCuV3L4J6k
Hi/hO8H+acURaGVkc0qwVjdF6pqF1CF8y01OyqDzS5io1x3SBNiW5zcncCdg8GQz
n8OYL7GMU2KVjF2GKoU15rCvgaB1h67/vMmHhw378Gi7rcWgDOTuBJSRkYg0yKcq
MbzmcUPF2TDpu5gyTxBSVIiyVDBCNN9n6CyAIBGZZUjHZsHugsMl/p0nWX2qNtud
Us+pc2Fn4kt7sJYR+l2SWRb2dWzyJG0mlmkjlySlh5CuaAUrqti8ff+/FfLe5J4e
IDnJuArEwdsrgeaFyqNa4Wj6NISs1ulqGsoToYv2VZtSQXVj/Vq/ryrEXXtSMrqH
mhu6hwkYh1BndYy4A0Ml12YovOLhjyDS6N1W7XOtnUVNyM/PA+C/SAS5CDl9iimU
XKWkZyg2OdNiWtHkRkpabA3x4DpP+rxq+SqSal0wXlkvtl73wNQV8vRmykj4srwC
IJanzWQnVJBEh6j9iNHPUYhkIKwF2dANlE4gy5eJapeECg665NUJzR5SZSjDD+KJ
AyQzamH46Qg4soD+ACCjF3cCiqVf4tIT9pNVgJ/E+FvtlUmHApw/5PN2tdI1W7Ep
wnzSDDd4lYp3IMY74haZAB/TmrL9siJn7EmsGGdIY5M//rqWZlLdsXxfsHS0Pw9K
oD4iz5fyglcPI3/XReD3bFgr9cu5EfxwUtFmi0RnnvuIZbWzzbc4e/aDpMWtXs92
icyA1tNS7qjIl/cnrg5PuHocR70I+VaKhSXIwjxeVR9Ou7aio9G9mHymmoueIKW8
yYc6MkWiL9ymHa1YRw2VV3Ykvuc9cvlmaryXFuGjLBnfN+z5WialPNBYHJq/N7VQ
ISNVCiqD3jfGQ+/++P1WkmdJKLijfeGvNaZBlzuI0qjJggWxTAJeFlU1P8hOU33V
Yw79YmfcddXYqKDzYiyNS19K+wv+k8iXfU7bKYzDDovoujVBqJKJXEotevgH+Whw
O3N9RcRM04djSF07X5NEbx6Nysf3MjSfwT7AAm+03aQFtHMUsEDXB8v5zfut6BLY
yxCves79s+Mwg8VSLwUHjzrOL2hFvEjdo/YKeT3/8SuRZvxGV07lRp601N1/i4vb
mnjLlCWWp5VEQb2xvbXAd+KFOlGSFRnm7jUc7sOsqN96vX/FQmElizZpBkoCJcKj
kNjDcSQlbt8UkteqoaI9adizstgTm6efnPMC/QIs+FoCTaXEEk9CevNkRgbr+6zb
Ha69fkLkyH8wDsGjEDQYK6arEdtt0jiF7O2QewU9gRfYEpq452DiibKAUhlhZemS
p1Ps5KPmKuTOuYLltk0FQsCYYw4OgQgzGkec5ddZegIWnctjaEyhmfWBLZBUt6nZ
lPvMgsc1P5AP5ja8HxUOIEt3ZLNG64AJuUn3OkxemSWm1BiJA3dUI03qiv4ipsuw
MCe13JwKbPh7mKHPgFYHPlyCcLDESCJMMI3eqMcBCGKKwD6Bz6MiQZZgy1tC+tex
ibkDErhpepmoI4omAVOsFkQ+/ihKI3mmr/r3ZBozV+K2NkmDfFM1WhOQt2bQKBZC
TJwtTE4k+lyBnkNINLbtDzJ+nxTlhhs9c699HlJ753hdJnCkGmGfkszc60BiQf0h
kFC1fhHSNQ7LwRYeEgSdNlNDPJWs58TzjTxwC0gYt6VY4F+Ww6sr+y1D4oXHI+u7
UTve72+JH7cxb6U7MlucoJO9UgxgLyzyI8ow3FuJiYoV7YINS2MKJHON/EYt1+BE
7zM1JYHyMvJX4x8COcbC26xToiFbfZWw023+9ppmbI9VLCw5guXS42lYGvScMLb6
sCsoIpY1sJpmbKOhmcBJmX26ksuf/xAHVzYC62ljUzTb3fAcyiToI5t7UDyvtdiY
LKlUERCYujp4r6yy2m95uB3VV90LbM4k034PjKACF8b2XhwYTefEsrgK+TL9mhSN
K/lS37a5sFXaaGtp2cY84qOLj2CXsVzfTTNLgmByA97imm7vn4u7TjmuwaYyJ60F
TWVPnV+O1iQTdzJfwfz5BLPxuWMFrkojge9Lg3eXPMkf2s13xqpoUd4T7gHatpLm
4A4n+h4oBxWIPIFUdo2OmZc5Pj+l3UswkMNDK25Ptq7m+yglJ5+R5CPRTpgfK0c5
UMwQg6tJNjVcF0Oxf2XqJT2zNqoMcrykB2uDBDu2hj/aRJhLsupOsWzxsssexDzU
DaiBxCDlIeEVNkXnonpOE5AhzwaxIaHRmHso5ApB/xcjeIYMOW7J5Sw0wUHFUoqu
+3bDO29VQr+v4pE0i/RW1qIwkuSTBMNDVHTqI6iMzW0Ah9vo8l7h+9yeau6yY7C+
ExzJp0OZEh/Y64JxnB28/OsMYcDYhgZ6RrYVvOB98yzQF8tK1P/JWR8Y7eDALmms
0uo7da+5ZDXuy+SzXPqjtHJqPp+OqMo1HssaCKVIwF574t1ot62em2qW2WFY2iJK
YGZrWO+BYl66njMx3POIboq6vDUD4Mfe/8VTswc1ZPsBTFF7zcoi+/0hhL2oew41
HxmpnGh4QpBnS+7zsyjX16obH8alrRYoJSkgK7T+XlmKU3b/8mLxiNMWFwOxWOUD
G3MDA4aEe4Ieqb+ECAEwQLjGc1P5NYYFbK58T6YQA2k/BLcqlzhCtTZcBwR16WGj
deoDKv6A+jrJE/4t/ZVADEsB/+hy7MzkGV7NaVtDpHd648HrvmE0xIcKYWRn3m3u
u3aXdzG9z5tRtb02D2H0xriXYHjQMklnJcgUQdkeRk7mQGmdOQmfGhpamXpvfV7D
kTYtsDQnOL2FTIVjlTa9TOf2BU3xy7YGl4I862aFTzjnbrNUEjgSyQrO7lfNZmiI
kHsYopsrk8LbREhI2B5Vb80z3iIUSxcYjnQk+GI6Vqi3ZFLxdKUVTFtRhNM2t5sl
vn4ooBgH2JAJ/Uii6l/yBeS6pp1jwa4IuukWL5WzwbGrUfxz9tr6aDgBPSx8fXty
s/LRCWoRy1xpef3ueZue4PpFADbTFtT6Y8WE2r3x1ta4ZwzGUJgcWnJFZKy7M7S5
trthuSv0beCbIXhWaooABkttpzL51pbpr404z0bIZAj6MM/8sJMlMXUhFPbWhdbd
vmhBT/jD+jSip+oVyaYHpEbXsDlyFKYmv9ML/hjW6a0TNPtXyqzSEbmvF6bKOAqk
klZfcqpvjqo5USajIl8Cuxw9I9VPZCHUUyqWRaXq3yyOBde8kLFiEr+JK223gEVP
U/tE/xzRs4BWTWJ63CqcDPawwGV8zaWVFvqZq/InjtV34T7gFxNZXbgRvtyx4JAT
rsAIKzbKtv5B6onNzpnwajp4uYqz3PQ5mTa0cuqCJtsx1V4gim64GmXLg7tqFvAj
qck/RW+ez8FajnnS1c/5J8JeAOt5m+cVTsHsVKRmsACPyjotDLvY7yrbz32p8dft
li+F+GRexRQPBKvouPnPGLD5PRw0uitBsgm4OKOUg5vmsrUvXePBuZN9rMwFd5p+
Jq0kBaEspZx8fTCYvrZ2z/jnS/X10TJmelXMP/7ec9tmVV1uRgfiAmL/m3jK4jJC
KVvvOHjag5WkZnYaGeYkVggWaIWJnkNGVu1atRNrvM4uXk4auAmlwLKnxVBqAIzo
f4iPu8CieKlc9yOIYLw9AXaH8rW0EDfQ8pIGyyqctI2y6/HWTL2r9O/+9IskL4Bd
KyPBkgONqfNH9n9hWq+CrotyCSBpt9L6MK5O3TcOq9RxU/Kp/gZMQ0VwyqlnCyCE
R9fUUIdIVuieDwhMVGgbRdvwTQzQoOPxSBxm6caCiNAfmnNFhmjjWev+n4Jnq9eo
J5guwMTw/EdXRmkXbMl/2BMndbI1ZeL28x6qgiAr2PptXIq8r0ye7hbj0pN5MWQn
BuRDyEMFc2RI/8oFYHs9LbvHz1E7cvpZ+Nh4UXl6E3g8M9HM1vww96fkwUKLVw8R
SVzmvidtK7XmqSfKauhdR1qcNGbBoMuC9woL+PwYR+IRAnSdOBhicdNU+EcSwhUE
38x1sZ1tdKngx2WSHufJvPz1WlzDr59MGnpLy7Gd4bjFP8WQk8xheqoZyhEyArXH
lD0O4FtLQD2zVbGcGuKsLa18xdfxuPgA64EXAP3bBCG2nasE5+EPc9Vg7Zm9PeJr
5birwevPrSlAyfLfz1838d9I0dJJNtg6sjelofC2TufSOlPPhyJ1oCTVv0Loybf5
pnM4Zm2IAhHL8AwZXIPUfO/L1Rrk4kjsEbT+MvxgTfFRKWM0Misj+BJjhG75mZPn
YJaloX2MlINx1l8rXW9oibzOauJSMVEPhVFCUVWCehK/qFKZz3HfPCei0SCheGjV
uOeuSvrq2018ZJV8OkPlPK/mKpBCC7ZkppdqbDL2/oHy7CrJw9aA7TA6nQ3J4FlJ
2fojaAbUB6r9zu7N4t+xYFLcDFajxKfl9wX4qEH84UIMmAE0KEzNbN4KohLLZsAr
fREfpJLmAEL+w3fU8R/yafR23wcu8shJ45dlhgnDns5kJOg0kYxNIfSlTLbdH2AV
ouUX5TEOn2ILBWkQ70CursWZoM9XiwUc0rTwPalYwqInzmt3qRhbofXOGcF4j5p9
TepUu4hg3KAjOuPHZHsmG1X7Wff0oEBsgynQRHwRmYFDwawGm3bQxF3+iLQUchqP
eGp46hKrPD9kdtJXWNlveBOrwji6kanoQ06zN3VkQb79EqYe1Fzz3tc8JF13WPhL
PbMreCzbDBHR7GMDLqd9IgXG97fS6ts9q2C0ARLAVyQjNymM1zQumm2SniWGAt7C
NKX2bszlX3jMoe7vq/9FIkT5sgebizcmDAxHI3H2SDv7Fa7ONx7jOFvN0Yn4VNBJ
DziPC4YpUMk+0mmkkMu6AsMtUxFkIivq2MU99GxLjEol8kqwje2Mppayl4ZsQ+Q6
eCkoTEhRkKAOKpuAvrWdDWgTuOVJ8sskN4u8Rq+1VtIOkNDD726YTh4n2QoT7LtJ
C6IKWBGCdF6NexWyK6dKP8O4cf0KkQlFEgxr/KrfYONNWEgJPY4qPCN7Fc9uZJ8N
mN+fchmHY1vHQnaXFgVIB/2gLwYNkvytjCzQhODu0Ec14p2rE+NXdOLmpoW/cOKp
H5UZxOlf91CjMevYe3yAXo6lz/flRoo6gDYt7u96kNeiIKNiDfDtdNv4UDhJJGIK
lWfoNt/EtD1CtvknVpslTq7wPLozgLyykswOz6i3g3zyfPLlZn7J4qX0EPwumFRJ
0TfrGOWIcJxG8sLHX/e89Kto3rJshm5sHyagMKTS9of3qavm8lZ/XqqCl1ixLUMz
zcn67t+SeI1cfESujru6gKr3d+3rBTryiEM/ypoJm0gnL2kyQkF9iVnFIMHskfNv
Z+7At08n349OGTnOOjhh6t7dC5xlMqohGRi3GvAk7sw5Jx1vuG8tnMZz8cACIpR8
RlsVLtDhkQpNvGSJlVyu+sFW1H3bW7cvYg8AnGaI3OpmxuapqRBTThpj9xZhP31v
OuPVN3DCCTBQEMiP2b3SKA/lgJCBDaBqmw1atrqHQf2QUpoBZqy/i6v53aQs/W6M
1qYZ5/dpGyJm+7SNrTqM8jLweia85MezUq0X6DNA+YolnU8Xoc6UuwRPSW2MhPlu
m/nTBD/nJrYzf5wE/+y+oajWfDux+ns5xkWMe6X7Tw4gp8PUaaZAbo4aQwdr/4s1
sS8c8zLDWDanxFvbgYbMFuZSsUtjpktXf/4RDwOHOsclRe+UPV/GZI6dDATZM+a3
JM6EW7pVFn84p+4WBllxG1oQLWK+DR7dXyTUblOVjPX8EMwAuTQGESC3KtKgn3az
layP62ymX26+7Tr3ldGJ8QWO9/CUEuLJPairAeDhNAH/lFi31GislJdFwvPAtCIT
hqGuKCO97AMn/HFhPTvrk81fuvnvod4Z9oXIkTs6cJAUM+oExCq/8HiFhFRoqtkw
i6YHQ5Ohyx1puWJMmwdIfw8sqnWf+JtK2JtSjLtE7qMO6hJJ1WjgzV//O2q+OUKd
cYbVdUWbez6zrL55zbjNY1Dw3cHk1O3E1r5PH/OB48PM1/Dt1D+0aYKEaO8bcNYe
6ZCY9BeWgzcApY0ZDKEFDbEMb7lp39o9gbDeMFtIOrudityEcg8ku4dXlCqULvuw
iSXNUH56lyzGfG+9I8S+Y1Jea4+B2jaVlsZSX9K/0G7WLAIF/F9pKVBjYWe4MMVx
rD7DFOKQJM3tmAmLUbkN1KQDV/jaFrtT/IG7HJ8huLPwJC9PvWPRgFdnRoLqZYLy
TY30eHMEdOf8zjxwUV9EH2HgAqE5KC3F53GY+7iyCW5JYUTYAL9UBnZ8LnJqwQ1G
XF6rTRfDMCr91we0TMf2bydknzmovfIeaUfdkCLm9DZ4JlfRCMeoUbcPQqo5r/AE
26G9Q4vOO6HRm266PrRtf2w0/Lb191LzwGNZoAFC8aPJOhnExSIfG4qWakc8Mwkl
eVqcQa/SK0zZAQjq3UQA14oT58txOzvaTpDy+TXaIYTOY3KVI5rj+xzGMio5HDU3
0MySp4I09VWcs+8NLqwXlHEABlHPB7sYGm3G1GaXMoNjnhz39mlJJEKwIbGojnYM
kAaoo+0bGhofp/AI58H13hin2EjHPNDj93FQd6a3VERT1NaUQWTZFANL5iqw323h
Kb1QqwDN0ueNBKJsbtCRcQv3NkX3OOnlD2QZzgK8COkmVvwTd6IUpwJQF69qR2tE
YjK6a6BSdLrcnBISASufhxPa3U9xA5NVLbBDpppdRnuqBc9yE1p3Pxw5KqECG8AJ
hirzHywaFzZual7wJjc4pxLZmiCOtTiGuiSjGS3xizjPDSnaqonbng1XiOU6jvUP
R2JPktklBYBFt13wX6U8Bat+WpSBLYKGppBdXxm5EcG1zUYjL/VWugVlhQZ+Bbd0
DInpFiabKsDeC4610zlqT6WRBiTrPa8zdzqR8aiK56n4h58TAiFTuhweAcb7IrQn
HbxUqcOV0sxvznKTcwqezbCXqrSTlyOK0H6S10QH8Y88nCJPdHqXoaiulVKZqsko
8d2RaexdKJ6Bh9qoRZ+9g8GAXiVi+iFXLQbiAb0X+7TtL3TXwxuhhr0gPqVRAot5
N3TSKztrttGBy82GqgLHkXFu4lHdkBjEtkU8j03tIQpR4131BpIZjGfWlVZN1HCN
Ni32hvE200GemXR3rTuMiJxS9ErAPyA25405WLSWQViPUdEvFRNbkM8DCbkVcKFK
DX19TMOLdi9kBVSlo7WFD0ivKaBBx1KMhmU2vfwOH49TghS5Um57frHDcDKuWEMY
UanyGoi3SH5Ru3duP1VOaB442WCkrO4c2QHSU0jEXUeoPEMuIQTrc8KIRaZxt4EO
LhxqJ8y7JuUJ3eLOsFOFy60ujbJC05qhNnoKfenMev5tIpQ+BHrgWApBiZ5bJ5lP
FJcCFaqHAHE3gxozKOxZFUzthBKpqpI7qFEVj16iweVCrdT5wu3xkHTEtPzPCtT8
vFfpe+a820iTIe7qphEj980RMcXPLtAhowkzepxdiZJMoOfUux8O+Uz4HA06RJXH
QqAP6cranVU/IK/BoExFZ0p6SUliqzO+uVrQq0uOgjKMtFqJecq5sVjDtalxWlVa
ZEF4O899rYRfVN0AC2tObJ/koXmegcYTC0+eP2Z4O0qZkY88CxNUK1UMVq/f1ai/
l+okRIhUHEmul9SEUsxK7n5xngnlIFCEczbsdVzDuEhY0Sz3qbbUaQhHqB6XGHnr
r91rdFI1YxhypEF5J8hewHHqsAPfoiVh2MKGajX8cR5UyGOL4Z+MEXuhX4yDq/yh
FnUvq7TZxNuWobaXfcHW3IrzLf+0ohv4+RosYGTr7gTFBptYhPrpLLGSZQ0xE1cV
lxhzMSSSsNfqM0BREHhRafRA85QWegzghQroMJwWKHaofK28uiRlStqHah3DZImM
dKIKWLjulX5ZoR1zKSJxrIVEpUB83+vQQPzx1cb1pSlt+glZFJ0me04bRafXHSt9
b9lO0BWdmaQxQ5X4PwFxBhm/dqSloTFZjbnGI2EpgHXs0IQ1JWqk3FGUBQV9EklZ
G3BOr+JDfnCDj6I0g/22yn4EjfNwrF2tp2Qk3i3k+e1figp2sEL/cFoFnrEUV8fs
LEJka3fgiOgRG4MFtbVm3g600FszhXl48ZLxkJRnWAmMN4zPoEtxMEZgONL5k3+L
El9Jx5h/aKjT9En/NLdE+EApnKyzvvj7Swg5tFq6aUEb5uMrMFUAWIrIUL23GsvO
Akfpw+pMr5JDtD8pQEahjQTQOLmG9DXvPYNIMLBB3TNW+YcZSLS+YjBNZPdtSmmx
wWAdXiTcplfROlPQmiDrnRbYgkpHMR5wvUbXqkoG1I1LLYBXYwHzrok2QJdWaFtf
YuTS8kc1Fw9hU5f2oihEAjfuLkynj2e5XdTNuaQ1s6C6ToHw2BnHLTghFkMe8mFL
+a6oqyc7F1z9wQ9wwJwtASuh3gu45b7In5TkOO75kUPeikgwJk0ZSd1AI+ocenCJ
lBUhJswEmSlPb2YRGdWUQy/Q2CTUwWhlS0fvu4aNMP0EIfGv1zLM/0gM7dX6zZfC
n4mXQusPSNq7nzT4lDjsJ7KWGRBmY8VJVMuHtaKlZJe5pRx+PhMRXw42C78KW9Js
TOSJy8ekLHaSwE/SfbwFiTs1VP9LMNdRIbsth2FhA+1TSkrDrsPtoH9udh9OqlJL
mXrbGfrgLNEM0YyMhbIE1JemeW/5ukwdXgd0S1roCuLA6TLHrzlOVE35CPP5Wadn
8fGTsY1X24uVnEH/i2u3qSU3Y4Lja3OSVzCVv29Ja8Q0bfTYG76BGFJ/FBV1kIWL
rGCD+dAV2/7q6LRyj4uUmBo7+PX9yuaB+f9pEcr23b+0ZuQkPEwzPg+zEsgi7K65
eYH2BmM2arlAOvRMw7P3MGfLppNhESdujyFsPVdDus/Q+gDyXddN8xB4QUgY48Ou
IQOTd5zYeDyqOXH4NovsqvnB1hSCqIuKsr3jsfvte7zSxpciw8PpvWnkWEc755HD
6FrEyg6sF96vJmqAl9NzXpfSGJyLq2wQnLGPvY/SLRmzSxD+qRwj0mkNAhnFTbK4
+ylLNUfMmlK/mb+l+kFkTEW9CQVVK6Z2wNP8saf20EGs50MesfvQFlwH6z89qtPI
nfPQmq1xPdr8LoLormUtuVSLAbECkV0SQQPjqbjjj227fgamYMHdZDWOpyk6d3wM
fa6+Qz4zGWzXQ5FwlBYMEWhZ0bzaAlWvu7X74xnsu3JmvTCbpYyXlXbdPksmlPSt
9woDNqRhJr7odQXB+uUwng37ocgRaFkz4Rc3Q54hbBYZYL39RXa2M/jBmMbyUApD
/4IaARg1F91Vomb9CfRz6NNlaUDEFuJy3B8eMpYiK6Ocqe2gHPy8oFv6OIbG+SFZ
rQGi54gI89EEWgQ19q3Gk80RCUyjeHgFGjXOydsE4mA5MXYbdHKk5uQ3VF3pXA/c
Czf56aOEHjYoYkWtOd0JQ/vGgU06q6YKzK3ZFS7YfQC5TmdUCV4C/nPQmRO0VplR
kTt7kltPPhdmuLVhLFnhPFp+xGKPOyyod8KhryyH50JrZbRW0zPX5ppDuAKrzNjZ
Njg5aMQTRdjhcLnDWrUahAD06/A3gksJpx3tIhCnAj7/m3rRNIXTBI35RmphoAk1
ezKMPg2AOSftwHLxDvLDsxW/Ws1fyaRXa4kM85j43ZIOEY7VihhKmeU0iHNV2wYO
+BQN6Te0/tJqu/S115hyRcEBilK72pAiuHjBA2FqV71XSB4oGx31KumGJZB/WrWR
H1ZT3tlhsXmzJQ9IOiiyncTMHPpb51/qljY78kP8bIiDXGJ9IrBwhibTuO93gPiQ
qImXbEw0PRtVU+/bV2tS68c4IlCTyQ4XzTy0Efi0G2VVBZ2YgD5GC7iTGLcCWyLY
OGcysczBxjGoNd9wo7MC3m19GJvfuaciBdB7QeBtBI/AmHXxaTn6b5vnQ0AO4gjh
X/AGzWtph+JERm9ZnPOE+cGVB66IiWjMcHfkepvh/Ks1Ge2/duZDbWBHU55IgkrE
MAar+3O1IWVTGSmzYb0fjNgcaQ6ilHKEQUsfCxZk4i14IeNbz4nDw9pgZi+C+Q+j
ELKu5gre1Gt9wJyCvxKWEBf4lMNAoAssXYMAuDNcPOM0k93q4QtH44UBsyde6Trm
IFdH3h4ZLRjaWDc6gOQ75wNLLq7O3BDCgdYpvu8JhZKGFVZ0dLnbmhp5yKATO1vs
3qH++x6UO33rNoV/e/IYj/4xwLp1B1hCg9vEx8eCea9M1VgpkbAf2GYg96YEwhw8
mVF3ffDDt9inr2InNcNiK1ARs+IbVZnowOuaIUH/ZA4nHPKUFDaaVefrV9T8WQYG
gzYcrjsfs65dEbs2hU0d4u4MRvkA78T2ZZPYYZMzVMcpyPH02tSP5qJQtGwsty4y
OWGs9hkzYxz5Mm15S5+/fXGrsOLdwNXZ1xXqnznI/3UJARdXrQd0Ccvib4mYzak0
ADq096kxP5WJRNBcivjzwOwIYv5K8isC/fh+gxAiZcQ4LBoCXYGw8v7B2IwkR6DZ
aiBwJYKXGSJSArUOb35mPQ2rX4N43T3mtWqEvMzzZuppYLsKEFhtg2xbtx3qqsEk
PeyZLu00PfSGJZuRrcNJtIuDameezqdEsPEnlapz0ihWERH2uC5G4rrECtw4LVbR
xP0srlH4WveqQ+ZR9pPlzQrjVrU/S0uR8iqfI8VvINh1JgyDDwfsNbkNRPUkd07f
u1zByGEv3vHCfhya4ahNV5B9NL9CwENPsfm6i8kv7DjG8QfZdlZuieBbRvUlNLDc
9reLR/e/CZAp4o44cKSvKeCxni5078CLJxxsQv7ny2f69G3YBgUg62JFkO8DyIy4
w+tdONxNx5zKfVVanWBx0ktworBiVqeXF6XYQyZYUlpJ3KlX3KvFGPla5ng//yUD
zBblJPhNu6oOYW2IhXbiSWuu4Ax52bU32+vUPGtRKx7cu6KV7BCbshO3gmtCglbx
Zr5eHnWbUeRQJDGKn9oa2jKEuClphOhi2a/oeuctI2MdcOQQViAg9/wPBTQ3xXsB
5XP/EtxVl2fm+nIdDe6Fiq5gZw0/NnvrodrsXJDqK+cdsgtifKhchYqhLIS37FEP
RJZuVPlG5ivbvObE5k/f4mTKyVgOeeLlNf9m6qfdnlsNSUZRSEdt9k/Xc5aG14tJ
1mnPNNmrLptTa0UBiGppZBnlRfMTuDM+6WG0RRpni5gKZQPYZDBkp7ud1zcmgn5u
udNvRTSEKg7FWLdpTNU2ODgPx/TRPdM5qnXRphFg16ODX97Ty5u2RbGsP1pX+Gq0
G6lI2Ds7nM3Ne6dE6oXOre1HIXlxQIFnc4PeO4g+y/ray0E4xhCWVUdlK9bq/DyL
S08jEJeS/1GveO+meeZr2j5lPdXnZa18iHpCSniYi20gNNYr7PJ8CdikrAOzEMf/
I0lBPTspJcsmrPiEhsCPWo367HVyRhiAoOmhiLfHQ+3RzqWjdlNH5WN7FLjOJhsE
py+AwAJoKWP4eIiFuVXvTZFlgDOPHVGtOXGKyMdtUkZSz3kLQQz8InJaWzyH+UAY
p8vQ8iv53n8tOK0pdA1eSzBoS+ECRe8sqdmfi6bIEztHdFhu/TkhLk4Ddl7ShVLQ
0EbbqZu3KjqLPU2LCDKlZ2ZQkrGKWTPwH+R1Kl4MkboG8mynmgHayAKBcKb3Wf5o
nS1tZ4G+brZShAjOLwg32mg1qq+8LveIoJrj7OF9gHA3SR2z+6lDGHsZV43Yqz9h
3PmOTSsGCRSPerQvkXWt3kxkYZUJ/Pb0Ew9a8YG1P6tIa1NDe5hOUL827n8V7yHU
sdHh7fCnagAT7LOwzk5Xd6rZXjDL97cNyfoO9CE+ozIWM1X6aalYb4w7MLi4XgBk
6FE4+IVh0C0FgTqCOTUC1myjJQ8/3YVuyL6eWaPwpr5F0icMY8qUpKNiJbjTH63k
ibrySvAvtxS9tJqDNxonwYbtiSyPvpGD/tmgLlP68+vJtCVtOTcb1VQh1irOVcIj
fJ7EvpyBfsTu8mfAYMdw7pI7ey6eX/wxx8iGujs6UC2YzJLEy7NPih6WMhl+kuJF
7MfklddG69wHyqrcolhiXig5KPuHMuRcaRrOOBqvslBd0q1ceMq+3NlJBnghOhlj
qs0kzl9/e7Jigtlg1Yc8/2sr1+i18zLxZb1zy1XHzK0UwhIQBrk4z0JykxbkPqCR
mROpiB6ZJtXXViT5Ea6blV24lCfMC/vdjI9Y2QyA4V/H5PBEiJ/fgW45D5TDjWeN
otSyG1TIH1h6OTUNDmxsu/rvVETz+dXW4JV6+7U+Pzb4vfR+vyPSTwkxiAhaVW0x
yBmHFU6Wi2dRQ5k//lfEHjfOR8U1czXR+dtVDhiXo6YDxoBgkkeJGktJZdv1Mrej
9OpqHmm+j77rr3pRw2KWNmKjlDyIQk7y8QTRkil54vjFWyQmIH+JWzUCd5TpmdgS
BA5PIT4HShqVzsQRZlhhUlgzGeWimGVuA0KlbKUbTpsssNstJFXzYAz0rGMVX4q8
DkU7WsmAjXaqztrF75GXcKraGsSvVqOs4eqVVt+n1JgVJ2ahrMOqCi+3pSgyD5cm
M8Zwsknl19PrRo5kwTVptUM0yptvoC6CB824luT0wakvKu92lWDyqh6HIBqGZoXp
ZGKYvotfV5FWataU0sX4UKtYTN/1/Qdk9/2nYuy1TNnXj4dQSuwa13ZJcWqjCRFX
2VSe8ezuMuionH0SK/47B6cWQqqI5LrEzlarMLDsQS1732CoERNgjzNX8IV7pEeV
OBeB5ncS1FXJnvLN+1GmWl3ARbGlgrKIF4W59wT3PII+NpR/IpsGyj1cAA8tKjnY
IDp5blqxnF0I7f5uDUOjbPe05h75EAFnCFpXqH/iBIthix/3zOomFi74deMtSxed
9yIxlsEinAllB9JVzyODueeacu+uLKGmHWKg736kB17Y8wtAvVddSCnWLwLfTWAh
2Tu4H89OdgcaY42V4wYFMRnZldkQnpvNl8RjYfVscq2wjyJ2CvbHKYTYXyPA1QpN
asksb4yMosaQ+MbFkEtQxy29d6jZUCoXiscFJskaiAStjTchHNakjV51slWxXIy+
FiqXeEO6JCliZziGl+1IJgCtbH/mjdfLqgZGS1DzS5FOE90LbtUwZsud8RL7LpkE
GwCLJiUs8k8WwSx+u26IE+4ommwASmItMhUDz6tl5guJZR72LeI3aDVwfqIXZYj7
EJ4mlshdi/h10ewWWgdyJdh+a7maX8kSC/KlvRlscMQZZ2fL3qo0PelpoLJAhMQY
JaOfo6dD9XfPE8MJLZoo+evnLZuucdiZGlef2tJPj03GR5GPa/yRPbL1QbagVaZB
/x3hMjKpUGqTd6/ctsH9yU9O7SuHbZcI0DkBWIrMdDaiVSnBkRL6hftHZg2hTtUl
vzErIr6T0Rc/d33u9PO0KRfZe7jgzv3+2A3yNk0maBLe9DxRH7yUx6rC3qEZbVg5
dzfH9XmPhQA0mIPNSHEUx5VT116nV05cSUcGcjICgC3UujLuHd1gebT4xkgcVhuX
U7cMsTaOyaMFAaytm/IAxkq0ZzUcOYuVzRCtVPS8vdHumO2EwN0WdpgWPugx3Gu+
lWX55pkRtXtqD3dXcW5tvUI4sbYGYGSWcPn1ANsZL+TN9n7KOKoKtg9pkJUfoZ3x
uncVRYTLbIKLzoOTV57D17lSHmeoqkg95tQsFg4R5ZgGCXjjYLWg5vqeh+098Via
rCUMuWyLm2+6dOa9gTjfOp/JIwAM7oE3iJSEhgAXWU8QYAxIyjKFSMkDzwgOtS57
TvgjAzHAP5uIRMrVkpzVtJea85KJOqxdojr7YNKGSY3Tg6XfSsZ1ljqfxHmN38Yk
UF0ukXNsVukf1Jh09gTWT4Uivv2v/Gy4Rw4hucTkD8Rju5SGK3tQ8z7O2qcn96DL
G2B0r9qMY36L3Vr3GbBVBXxPI8zfMVznCtIQWg7dm/UF/HktDB0UrJY8FL1XhIVf
89fyCdfKspfdw4yJd5Z3uSGfdRDqRNQGpGLI22LXxtwBZ+UPD/hwyUPtxaVIm456
S8Lw9+16TDzmDMiWvkaJpdfqqb5e2N0OeSnk8PVa5XM5w0y/UlTa8LuShDuYbd9a
HR1SAd3ugkMee5eCPGrBzSQaZ1y7ssC7LaSJb219QIKU4hl9Pk30OoOGMX+iTEEk
CWoJl+YU23IvPZgkmHg3w1IPU7o9aUI8el/tDwq//NPjpbEs8TwShRkg8H566/CK
NqWWH4KorSsE5HqPAZ8fgghoycUtzGjdDc9hKlqEgfbhrnkKV3DDdTJqry/j7gIg
nyoAKYWnYwwOG1pDE8m+FiNABP7vWVjDuHefTCdT5/UnLcQTRdgV+8QcxhnykoE0
4Tpdy07lUOmUbW2XdEN1exH9Mvc33eCL9UZq8eY7z2IiQ23Jd92ZTmTcS/74KBiX
Fwizu3Msb5BG4SGdLt7cIQ8GtnUTo5pHZm2C/vrzqCMX1YiZ5vADKd575E42Jmty
JKhM0uhYemamQXxWtUzSBVPTlXpcezoC5yRNXPXpvLYUVTsN3aC28XeVQ1BATyNL
FA20rYJdxyH1zI5LX/DoYj16hUF6hyl4qiQVO9zI7iirAGxw24h/lc6NAXJ8gDRF
3+YBU94jq6JQJfepC9M2OFSSea/g7mTsHYGpYyLwzyhYgt+KlmXj01tHpLQbl1If
TLAfmN+tDHs5S8aUZfn1Hpf9tgEiXhMpK9cnMPafiT+fb/HQC/ztNLixjqMOKEzs
JzkJERGuWZASUJmMicJqlf553ZAmsYjjRHu8mMCjuWcBNuoC1lt1VvKDY3h5vztB
Nq+I2R95ahcSv4UcJtUiT5MqtivI7ETgAqo216AnxUFj4w/Qx7cffBm5nHqDh49h
EDku34I2avwFGUBgpsSqnHvwsrXR9gVnBAjc4kTbGpS1awQ5al3xl9QCDIrwmw/h
2mJvz5WiMJtrBHvbrfR7vHHRMk7koFNXR+G39DG4x+9USM+nJJWYRsUo5Wl8XTYM
ZC6/MpftcEzU9nuflFMj1NhiqnOH8nHy3OVccwXSsk9SIP2Sked69pziBqz4ANyc
tTacV5rYbEVfJI/ZGHm0s9nVE3uTxyISzfi1M0hVrKOs0o8tQoIbF01qbjVdGIWe
JIkDUSiD0k+1k9AahTWjDqrQZPy3bti7eKfedAOHPoEvdmCmeyBOTRpq4GJrjvBT
DtbDFrQcHjoXOgBY6kixpmvub/XzsjFC6WIOob95AX2vBc2dplyGKY/+msARiLJD
BCDab9w3niAu8yh0aq2pZyEc1+PJgE+gG2ViybO3OGdk1M8VvRNNKUpRwivyLEQM
fIkKFjKboZqMs7ZnqMvGFvh2ZiQ4UlOfMnqpoCorTMLxJe8xMn4bADcGszWERGqA
09qg5Gwna+KljbSEYxM2n292vxHJL9kJl+7JlLi3RqyZtiSZrMrgq0oGBybhaxmF
7UCKCbQDvANeGFHHzsBy8Z71B2WxdTig/rEExM8HwOiU4f6ivsLPT0BNsd2ogh59
8sE7QEhhm/It9Im4zBi3WA/fJLXXt5h8Qx+53m7/Z/UJoMzUDNOlpbYmUuyq4eXW
/KH955X7WKkqQctnIGxfdJDuRpa767jTlyYNL9+q/J2T+ZJ/G6s6gTzoMHg3QiDt
lYexVdG8bc9ol0GaNtHL8Y/XSVCAHZNcnjAUum7BcOM6vw6qEvgJPVmDqh084jJ7
unZSidL5+6gmjvBuUGlHHNa39e8XyLTfhj6H7BXkZqjorge68GB8j1lMXxKrAHX/
t1zQAm8e76Uzf7pFt9jaUHf3pM7A+dzMPeN+7HiijnHyujCmxYFIKh2PImP4UlFy
VkWxoOeijqQBleEFdbGjTsXz3MtT7lkFPB4Nm3MWqbz2lrLHGJgiYGXYZVBiwGgA
7KIL1gh2LpaSdtgDpzt9XMF7CwOQU0xCGqBKm/EX3Z0bS1qnXQgHrd4C1UsQgKBD
yAvRhfv2SotRLL7je7umBldsRdXLv5CYYBrKgF/qC7JO6w47Z1zTQj9xKeQ5oSo2
Zo7sjRX78zuogEhSU3d9zShtQqQtK5uk0e33yLzJ1zOleMVHas9JFp7njuXnLO3E
4QNq2VVMJJmqUlbOooXZqH9XKXopwNzF0Yo8iF6aAvzfbKMswXh36c1qep93f7Xd
tP+ebc5ynjiWpFzBtFitvprEehoQ02EFgzWcgZERxbLQ8rIjyAsSezXTewAmFUSD
VKu7vGnG//QKPscyoVJDDYPWTbdqo1qEOJ6kBczeeun8zhs7zbEy37rg4YJc71U8
HSHt595AO4oG2/HY+hcCtKZuhZXV5yt2p/TtjbNVE/yDPi3LpFeVU74EGvzHttO8
uhJucAKRTuoZXDgC6NyGmyK1GEg8VnMaGRWIh0MlqKk7YuJiEMv2X6MN2mdY9NCW
iay8G3eGaf6Hc2kmUhXTmTfBubPXlIYZ4dz5BE6KbUb4VnZfbvh8/MDM22kuYe1S
vn0JfootYkMMOVdz/JQN7yC4FGaCeLY38UXx4c5ammuy+MxHxR4QnSK+tnN6zQnV
NNqYSp2AuTeEfJQUvd4gnpShCCTDN1sXbO84pRIOWUsbXvGK9QpOXjtvFaPb48ZZ
KM2gS4j84PCP1aJKzYEhKRPdFNQkQ6/bxNWXfI+GoMDw7MDwPEn6fxUhI8x8i4IY
/COqSr2gWk+HWhCTtFLM7vz7LL6JV6LDM6v+jq098/HawFtQAlaw6RrZCUadfR2l
nQMitrB+In2XGqmH/IGbeGlygzRX82EHJdsgQ8B148uINvPocYByE/6K0mVLpv3L
c4ssrsIlarZPYbPXGi09eWq5/VARr20zm5ZG978bPVnlp/gl3HCPn44tBnxgmil3
ADhH7dZwN+EpjF4fZ9urK0GqYdv8b44ljKl0q3Gr5zUml4qryrtiPlur0RxAgB+H
7zKiLsJQw/LdZ3qn9+GUAUihMTn+pgwoHBVclI46FH7QTOhTVVMuWvrgWnE+SJk8
Bm9Z2SGrAD7Cr9JZKROiLmndXHNfoFHYIXxxD313StWlMRBrmGhrd7IHoJzP7tuF
3/VGE5ctjHTa6i6gn4qBAUV5fq32qZZCEX2j5YCaJRQA6IVFxQFGU8k/mn7QXFLX
XOjDzQofy2xfz6PvXbqtR6ceb9GPSsdPCgHZkYBOc5V8/cn0qKGZZjk8IbaAPuRs
xeMJ47JFMu6Rp/nfS5LMtrhYIPfxGLPkJQzXhjxN86rksXlFfEjh3wV2At0CXvb3
QnH8NBWSm7jnFaTVH8pzFiBwa6EUKjtPmRMxPo4DhCcwllZJjb5/8kZDM5epxId/
10XjgR14vqKGhhsImoPgGZ5c8AyC9uGOWUNVK8WP+P9Nspx+ZNffIvdGl0eDMYNR
ZR8KxvC6tqpNR/3ptM6UFyYSsDDytjICdTtrwjtysEuN69YfLlmXS+w548mgHZ7e
HgTekgGnrvtg0UsrXZV26mUM1PGDZE9raR8nyFibsMH6KDuQVg9YD9E2vhek05Qi
iCHFf8tI1qIW5TAkTiPxhQ1kILbSrVfX09zzr7XYNFaeWaFW46gvdWPuz+qFxslS
qdnC+yTdtPS5CsNYPfSBQ/lOz9fY9KaEsGXhWYy5MOt2zgfCYx6Q/+R4djF2EMil
TS3hNKFd9QxAB16i6zbVVA2At5ePMHCCKupZSKIjvAKnFAfPZTFMUUpOBsm8MPo9
JHdDVKmBeKi9kLJYe1ri7HsKrD6XsGet6ZRYrRU6t81fjHc6WBoi0xMM11EjaGyz
PCSYs9TmluTdZB5kzGMzg63pfkBp80c1NXok8KHEW7IWDOgkUkao+i91fqjr7v27
Ag5eoChtLJVJ7LEcAH2YfIJ7DCDvn12gnPCeACEOg6/L7QCuNyTe2NFQaD2oo9ab
AbM9elKCBd2cYmryioGmzwFLQ78wNqF49do59dZU9Zh7f3bBWoPn2JpMaEm0liXh
UZ4N61v8bgH8PDgEn+YRL6IvwVGOrzSKTm/BUbFgrA+31ZPmZWzJFm85bmWz150M
WWS17ACCvpmNH+T0A4ta3Gde60pc2Gz0FGj0QHuvkHn7P2TPioyM1+9DpB6SUG/p
zuuTO6FpCXMb/s3Hy7xOfwaJroBrlrJtljcbMHMv6Bsysq7whYrRJowXu9n3agjJ
B7kcZMElrBwGK7BItIjuF2OPs9b2D1judwFKvL0ykjNYQjHdPFT3riwTKpxNttKZ
JRMjTJCYdmDkYg/b1QrcN4ZxJXQ0ZyET8wyHOMaQmgkHsLx+TJvWCF+OI2c78FFT
MgFmgstU9WGXJi2f70jODTgiUhKKazboNZR/LcKc8fUU6NiupLYnAIbu+jnIDtaI
ArEK1KlAuaNDgwubaCG98myu6wYxSyWsmiLVBU2zft6A558AtQ3tiiy/tSZr3Po0
1CkltzBk8bT7x6x6x5wWn5YcshuHdtnxE0A7Bu8U4Hy6ZanUVwCHiyfvqSOn//aZ
o6G+VvFIHDxeIfffMeqRGpsGYUVfZsTLfEFqCQRwOeWyvvmrIpNKhQ15hSdpwgFX
qO42zohkZXsdGT1hNIVoelvHU2H0ZA2kEAZuXVn+YBWFp91Oq/Bg1T/WEBw0w+KA
QRHyHPUKGq4gO5kReT1b4X2vyo7sMSPpyw0iqCo+MmbwTYFhYcEU2zZeLI4cyYX2
mAfPY7ba8PjdQrUSsnAru/cdQxjpxJtoQ0HYBGUA2vxbEF76vC2BBkPrC6i7TrDZ
TWOeCs0LWta+4Cn98d8yDb7UHjNhy0c2FwxfbjLfq6SEtNHxV+vMymrKqW2P1hKj
m10mtRFjVQvmmzYudbffo+dn4EWEKLHiDC32M+s9lDlx3FqFqhDgNSf9Xp6l/UZR
Tys/hGqox8ntIy4XZoqyRarOR9uF2JKNa+WGDPI1LbXjb1KDLR+zZ2MX1e+Ze72Y
KED2B0zo8nVLHBKgJ87eP5pUqmM8SXNbzkYdFo/r8Ga7TrNrgfkdz7w5eJNgCM7v
BMXHiCutEFhV8SFLP3slmirb2DBdRAtQRGERAqaBu89etTqjMJoOwNJXDijcZ1MX
GRd7ou+kuEdiXTLzhs/X/CKU0DZY1Y+FY4e7QFKcQwkm9U/x0yArvxtjmuCCb/9t
+am2nCh7hUMT79FGev87ozodEE8VSylVA6/ah7vHbJjl6wXAsTAcT4xTO7/gZnTL
DMukEmRFzCf3d7JAbUMZr3UQDaSwsYqcFQEO+osk9wruQk9S8OvHWUnHvTMeJNSb
uxFXSexTJjRboo7ny3GYFRfux8hpenfWi9YBoxAw+IjbBwWU5W40qYoFgmP+8ABj
Jq7SQlQIpIyHUMjetE2m+h/tg2h/JmJNMY3MgDoaYchbjcDfpnAtb6cLL7u9jZ+i
i209Bb3abTc11el18xwyUvM6ML/uIdAhTl70HLu8AAUKfucSZ0gfK9U+0jGVD0xE
DYPKHJ1yvaH2lcWQxEhGp60V4nPkBbY1TzDRkajMDZ8iw4sJuYP91XZIGrg7cBFC
A5aQkeqbsSElEGVM/P2+5RHpMRs9YWw9zw+d0zt36AR57VUGzr/MkpTcAz7SfDGh
4PGL94yk9FH0drxQ1Fyc6IuoWikbAYW9B1GbYhOKwBSz+JGBtJF6Ux9EsivyXBa7
PWtCX+ehRBpvop/xdo/kRgnAAkzAdHQHYaWMZDNtwInOguUG5zn6XwnCgnKQSmHD
N5fJNdnZveVsyiUfAnmFMXoHRts4THAQiKtd9GreH29NATCUIfTwGRaPZQn0y5S+
+62uQU57PwetyNcqB/1v0lNOFw6OkIUIPCI+Fsvh8pidt7L2bFAMT3+Y0nZsYZWz
5kHu/bfFOxcw+yiMQ99SuCGhK9ThnQO2b28DKJa3QNicd2NWxBpqVGvu0JdACQ52
t8mN9+8LM66XpBxI0Qw5aOkbrpSl/KjNqjgyJiCzd7mrBdBD8eqfGv8YePyifYf3
hTAKKSynNHKqc2dMneQUZ9BYss2WBnFlfDA+zjnVu5nYhuUhhcb0OJNYLF3Kvhsp
RFLjNK8peqDZHmTVg78PVNnhWv0pGxkj1dm1WYuVEq/9vw853zPjJ6DndzbGJFH6
KQdRUompt33iQ6q7n85S8C5Nxu1BNt8p3pCWC+fqrE+jpsY6I38yBjtbe3fwp9TH
wXuGAlZcASx8BN4lR353Fp2gSHWKjFu7ZAbc3o3QwHDRaaOqxMpqTS7FaiEVb+/K
rhsosq+8R1bsm+uSM4Y+aqx0kk5JlI1urqwuzKy9lPm+0QsFjMuALLYTriJFwcoM
YQqmrFbjtRrcx1IecOfWm/1ZqwWPoVsbuulVe/aGmBE+abPthakL8dAIUcHCbg1o
fcci2PAgwdBfQS1Hu26JWd0by3dUR6FYWUjyWinyRc7Bxo7/0xNJ2xaKnidhZtiz
aCE7NkgW6iegy4x4JTqtqhAUKStOzQXCBjhdpi9K8qHMldfeNSula8tn9UJab183
vCL4+TLblBOx4YOlUGUZ89QeWrtmpbMOkSiCCY2cet12vsCyONbylb6WR6rci0As
BZWvA+HFr/VMeE80LJc68wE+pYIWt250n8ZH3JxOojB0wP9tHuG6wLftuZ+KZetp
SrahQDrCNBU0Q9G6fuxsNoqIgTmJwRaiuR5PEqtA9biHgZX9bUv0IBZOtdgwCaTu
Oa7V7HrmoB1PARgI0n88Bdls0uFC+lUaW/atYiKh8o4FmVNM+fyku9favJEBLlzI
Z+T/MCwLTQSac/sRrIldoFnmIs8VnaTK+dFMdRy+da1/OFklTujCNseFu4fBCYCi
SpBKeKwsazhH58t1wUHnBWRAHq1TzxDb0HLPDreg1XVsXlH36Zv+8MR4GlFHZzPZ
h554o9sdB3oW5LWQ2zYBLG7TX2adZMKRDGEaRM0lAU6rNXy4lSYLrK7EhDAU3+Ah
KYO5U2ZuizGPhI2vP7UBqgTCdnJQNvzbfJrU1cuRrSbh634l3tcETYAY6lbZe715
kkSUDuvL6QmiM2vzUI1ctnd8iNF3n15A2RZ17h+A7upVxpIEE8816thRRUyo89dO
uFKquu8iRhk685sB9c2snwJp0+OFMkTh/JVtgVF4vCpxgYvcZPlJqHuv5wc1uKpJ
xFk7FtvUYe6VMpvzyTDqSXlIVkoxLb5bbexCsyOhRchRaselaFJa/e/yBGUKoe+p
yOhfeBXgiGnYj77r/eBm11Gq7gSKeK462OB/LRxA3iZIJtLbBpm+gVndEiAgokej
ArBhskKoRbW7c+NpKLXkJpErSik3sXhMfsMhxQwGiAUCtBXQ7ETsY79e5J3CcfYC
lM7Qke6qJ8qR4hbycGyA2+kksNyIP8lALhPfd5rcJiitQcEWL2ywNMMJ1I2qJysx
HNMAqzUK7nrg1jAMEglkWOofoK/BxFv+lCwoo4J1u1C1W98ABMPwoGzV3vp4cIBi
3SfvQGVVFpo9PzHse+kQu7qF8ZBzIi0SHitF0dSVJd8iXMgNPaS4M7GHN2KGbF9+
YBR1gZd8P++irKi3ixJwFB+SEpgdg5+/G03m3p4mR2cdy1cqZLRwAJx/46CPkFiO
v23D2NsdBTowiq54Q2x6QWFMDrdX3yLinumfqsiKYECsIafZ72SCLOXUeswHHsr1
3SmaZxyyj2US+8egrWn34NaPigPeFCe5YrgnjYoGy4G5JGSXfz9jAH2RVlUOtZJd
hAtjjtdvy3FtbMxWkOyuzhh1vr3UMcBs/f6AteAIXw5J+sxY3GfcAsfPUBGWa7wP
d6dHU8N7foHZ8QTBSWkREuw2c3i4R5JrVoAOEO6sSdhBfoxLbqnqh+6hySw2b9Cv
Hn/wpKSA+3b1P6RdkiGP1Bynp5Ktry/vJkVoFiYk22f8NqSW6T8LHm9HQAD64oIa
djwIgjmkOfOIuN/7OOZDUrXgar6mE06dlvcQ4vhaSQKIAWSkPDEdCXMCwTdtLIP6
KpucRwVCCBAstnPaL23Iuh4KWaV+s97mZnUhWhSGgBIIdxTvVQpykxBQ9s9Pqqjq
VA8T26ZtUPkZDOLLTVD25hpEpzZiLGDtruG4Bpo684Tdcai57NswJ/QxIAVqP0K3
k9s3o1Gz9XFx8nI9YB0vrPEWZQl3fw0HOV9OEvm0nf1RA6lQ52w/MOKfUnP+7KGu
h4TWIr7Lewe6Cvac9HPHDFGKsk6vJjqV0duTS7AIKhjNTmJZqSW041cM/XkJ5Qhp
/U/oGyt9UIs6CEW/vmmFYMV9N0A+AXuN1Ff7t08knxs+FFHIT3Q6rFfm7Hwho2C+
MwyLlHnn8EJyYe1PRY1tBsDtqBv6YEzHcbv3H+d/gB7PYNv6BuyhICZM0rJbybKI
4MfnhZMC54sh5tyu9t2WC+qJprXI/GKUNdv4bVql/rQfYwSrOrNHenCya7WIyaE7
PC9HvVy2dIUJwHavP0qy9+BD9rWefaH4MlPvrkq+sh9qR8I39ovbZ+TDJOxF77ft
rxx23RZtW5LH9XVhc4LCSFugQYHDKrZpn3Mpwo1vxNQyg4H/wnizv+K4OCQl8Hpq
LAJZ1FFaE3N+l5jRaAB2mTGyX8ZuM06+S5E9xYiyuFYiGPEDaCZa8aTjWz3oZFYy
Romr4yNHkonZ4233knIND1nU4Oie+C6J3F/0b33PAGSof2ZwmiCcCYEVQ5CK2IDU
o9Lbt61fghwbVI/Gu0yYgT4xyW6+/qApQQ8lxIHoYrsKD7dDr6TsrrwONPL0qOro
HK8RdMZsMkbQ3CAosBA28j2qGtn2qLXbwPna1BKzxx5oGUo8uHVuV2RU9perUE80
YERl0VxBbVylCzNuELo8TvVx83qgtgDRDkpE98JYTHZTFmt57fv2wJjdQIilxc8D
gY8mWeelWBnQnHqGeunP4ARHZ62xEgzKKK+2pmt9crDceuK1Cd52g5uHA2+vj1Rm
Mv+rAzMag+qfuwTX7waCBfz2GzGtsQK5mdPJnCFjnxRXuoiLFF6mGh17L9UABAty
QtE40smHtwt/j/l9fVfzMc1Sd9qQc2ikmclfT5ATKNPUuoVzuertlrmv81xfF3EV
xlXQqL+njcMQ3jMP541WsVybVLAx/NEpxZJHrKeZwASqJNF9nR9ogF7SpcWzxm3L
T7ooncRr1q5iAE0oadtnqQfATYUuWdnWacBIHgLjFlaM+o3zGLrP8qcXHcKgCcOy
2JG66CnXp7DbY8gV4GTKhtzqk5kJGegFwgz0tBroeqmfZf0ecNg6dqKRgWHFBt6h
xfG9CEdXDJVVckZL+XWJkVHCE257Z+xxXt6k3v50nl9aTpgKTLHNbySho8KOdY4Y
nIQ16o1F0j4Dvyd4Ck1ckc9Z/GJzZ2KJn4sPG4kwAPWsq1Vjp6xUx1OqtMlMYT6o
/oD9axeHWVEyqSqHdxg6dAfzy+SDgoxZXzGJfuwWypbqaaNbSk8n+Exa8VWJzcX+
bTBsHgQ0S+/6UVham11ifSzXGWRLp2CYMU8AlHiE1yUatXzZ5oRUbZc7mFhSa6jI
5Vy26/GZAeovxDLM195EJE6j0kD5sNPA2mjcyH/6oFU/oBhhfMjTysSTQym88QIy
x7yTNCrLJOD8VfSpbVhlmiKumQ4bENBXiypwiqUSZRX3UpnxFHToJsiGWaGMAnnF
VpZC83qvXNuhWg+nViWHuimwLHpeGpUhcVO5KHF8YAUH2DXZc0Ic0LUVBLytiJVv
1rEDjZnLLJodXTHssLPTTHeFmwOThd6rPI7X2t+Oxha/ltqVCSnRMgOoQBc2j34i
IIkW5x7C4b7bhf7UqAsPc1m+WYAWNZqUzUge2QIUCv2zAwqwiL56MgimWfdgr9St
KrjaEFz4kiSftdhdpGEC03em2OMhcvJyLpKbMYKjgA9dH/RkHMLNR22UHjASsv7d
QtQNpNWqR6lv7SKv1PSoAo2DrG4URQMfi19/rT3E7pXuzthUVKzD1po5qFhS3+iR
SJjcCkHG5m3sD9gdG7CkVzJdBlpL4Yi+XNBL83Y4UtZJlLWotNqEf0USTEoxi9Vp
ygDcmapUXLY755cMkRjT/SX7e/vhk076Cl8J2lHLlgeU1kwuv7tfjNxFpcG2swrF
U1S+4pWIjswHcl+HL+LWYmBm7qNl2pNe5G35N0r0zOYNvFVMfWJRyc5IWWJ+sLUg
lWINVyDdiHEj0WDqzQF9MNTHPFGU3EX28chgdl74Tsnpw1CnLrxnE9awb2Pbq1q2
BZ6xfi95uW37y6P3OwCnrIGDh9h7LrkE7jOPU5O6V6HYcO13b9Nb/yJMddyjvUBp
NrirekFwJ1qnG9nYtVoYFWobJY3vwhg6tX8LEzwofLV9sfy5q4JC0XM0LQg+4WMR
/5M2f1RzRmHsVtvdqMrka8o4ANhP0cJ5CGfe20JYDbn6/SlapbmTJEB1G8x73eRz
0iaMDa5zrqaAIa4igUZNwPtufrFohSdZH5RS204LilUsNXicMkirmq3shn8WAESa
tYOr2NpV5JANgE6TQv1WnndF9LFGgLXfD8kg8fj3XwFSgiZYJCKbTkTT79+y6o3t
W9Fkr7zggzog7fXJvqK25Z37m513mbh8g3M8PUP2UgrOi3/gzFCZFm+lPqD5Nbxs
S6EgAKh2ZLKf01tG9iVxdMRK95VAVnOafqHzSGGzLraIevVq5+QIiRbFs/+pV8H2
bYBPzBizB+UtHFLmZaVRBidy5Iwv8f44D9fCZ9M+nJ+fnb8kzoWDG9HOt3+PexrI
/CLJBFMJidBnRN86Z0JAWyGWLbOtGgTKCTA8oZs3VKxmNXDTEq14ca2NlThpx2wL
WZbZkApMPkcnUdnQqvZw8LjRkFTEXtvRE70yn2WPca/AxtAoi1tRkkgMZHVS/3Oc
xE529oJwp6ta/9aOYr7fApLy+7oZcg2e6h+iXL9Owv5D9cNZQcNYZ4bHYlnq+5rI
wIHv4JGoLgtE4lnmRxhfL1dHJDIHn8FUd+FNa8J4UiK8PlcUvjP+posCgmvkxfMX
EFTjonBmOrCoq/KlUexsn3YjMDkXLG/D3RE6Z7NAQdN5SG73ZLwq4iCsVcHwYKCL
+oJB5vA18/hglDIWaS7u9TtTyRU600AUr6Cxnsr3BHkP5ZIS8Hznd6YjSclxkeI0
2u7YgBDh9tkXdDD8gWB6xbggAGbTP/fAWd80w/zysyxYmNvXf7y/qm+okHodw4Vl
GLyn0vAgkM6gwydhpHA8gEVXgSL3EkiA13xZh6BLwfjsfxsaLebnSBzbvXb84/d0
8XUDtt/W+kerO+CDio4C72hy/ivtMAl3ABaYxcZk2G+nt6c7sYLAwrUqPRH1xnW3
6zh6jizit+CxfIq0q5+BcowsorJQ5djP+mmiKKd4JJRoduuW1j3oZ16A9yqwi0e6
83kEV1bGhHQVhgkgFP61mJNIBfibGiRcmyirGsGskSK1l8vhi8X/D8E14OZhdHie
G8zjqU7hTh/t1D6eIY15bp6Q/Mo4nOgt8RGd4Dpq5fvh+iIZ1cFx6jEPFLtRoYu3
ydOORn6nRM+KbOyJBLjREF8fbjRwm4XfYEJOW/V1F4WbeqAniaaVYl8gxYG5MvTY
+0aobMagGG0D7XT/xXF4aub9T/IHy2H+Z4YIGIb/KuoIiEjbc5Ry7TGY9H9XcN9T
XB/atkZ/3qCInLPu6Hfd6kahcgohUaWHZYpc0AwewNsHPUO8HO78ASai3/QDlBhy
JJEFmWtIpktaMLxAdaIyFngfWVsFyE79y4RzL3qsiFiANBwbGnnHh71ibUlJjNgt
2E8S3kujQzswH5pATX521e4dC0wSjY50nJvaRR6cSSUXJV89FD90de35+tOW2Ry6
x7jJBf9UiLuWCmLLORcm/wBQaFxxCOvOR0hM6XAf6YNbIICDDHjdGSZNKM3YXocS
4TMTATPlgD/iqlTrXi3COOQQ5T7Uearmw968OykXDk8+9xdhgGMkQXCd9A7+uRAW
vGcWB7LjnovfCV57RsRVWnoJADhWGxCm4PYIFJ6YUtzk9fTFIOWUfiLnuriHAe3Q
pQMcqZt4Cxj2jAAhueSMw+u5/1urPraM1ufgcpuqotrG6MFfH9uMBKspPQeOTE62
S0wVkb28c7fcJmODJ0ULXpaNYYrbvMr/Y8rr+5KwT2O+pYaAJA/1Txj00IvUjMqu
zWGNC1M7BS8AgQ/8z8od4WyPmXGKrn1XHwrdLthOqciYLtyLwy7XFbuWnNB//xel
DAaWYQZJx831g82DeOb0seXFtQwwRXNC4YcB5ud/wqTtxEJnZWtl5XkNRmYtt1Ml
d1JinZBXG7CcG/yfMfoTkTHHo3WlsrHD36vBqSggeyaUqi9+03YXabV906xN2boz
lDvpS+1mm8jVpUKQhxoPSylB24At+7pu+pzHsUvWskNoVTvdxzkvgTXtDQRBDZnH
T/k0E3X0Cv1vaKAF0X34JrU+1ZFwhFqePrULyhaAh5fVfWlJ/s43O6zAo4MvGm9X
XSSoBhOkmn6wcOMKL7yv3UNTI1Ux8Ztz53lQ+gcvs+9Q5ZE69MPWFAB82pIGlfmp
E87420bULGJ2gKIFgNxYQrdaChtXGtsdbgbeTiU9sxCJVJbXBVyc1VGXbX7AcGYv
BVrWmVSD3DIOTlwFbPj5JtIaKGF0BnjjoTbeAXy+H/b92vxexwMPeOe5PkTjnLaa
tWBDTKY8sNSEMmVPuSSQSJU1gmu/rA+86faGkcL1hJPVEM6oJwpm0SumhzxWhYur
yr0dseTwdSUG1GVon/5GyGQCRMzs9NY2+XXcURPHpW+PXw7IVRpJTQx5UJW5oXSY
P/V9Cvw10MnU7GZ9Cy5+P40Z9gZhhF9BxQNxOMhnWB3z10Ibcj3sBSvbK4L23uxj
20xZ5AhURPnbng5xOxb/1ZSzRpf7uDDphcJybudX7N8yl9lJ20xcD7BIBfNAgO5E
9rzGkh3Kf/YeP/dG0I+aOkeP08hazKFZ6X63mZpWdXMLvM1kdwKChF6wuf/6YHf5
DHLKw2l0L2iDonlZgyVUUAzBCrcu2gfj4jsvyGm1OYG2HSvzTzrNwv0iHxQYE8Oj
aiIzlQveWpQNujkTPRjAKKNH4huPWBgBTVZYVbo5S9tiPi2+ELrliJs7pTQbV7Rn
E5H5FxPAQKdBYRq8Ys19aDNLAjLqBKmqD9F6P8ZJwPxPlf4fYvqnK23kZ+GSKET1
9C1VP/Ke9y3ZwM9knqnppKXLP7DdBcFrIwM0e/ZYx4Uj29tEQg9wiu0zJBucxHd1
3NoeO7gbs9dpZanw/kihzRGMsD3O9e0Q6SvK26mXeTti4ZUqPf1/8BMZ+0aU/SpL
sttYqgh8EgQDJdZMR3tGmnjUralLQI0DoI/Mz206OVxFLvbsVSXU/x0LkCwnX+Ex
14iKVGRS2dk6nNu/oWr1oTGHEynrbQOhxbQTYsbU1BsIIwIgAXMjbPdVOgTz6HOK
2lH22S/VBrMpyLnsqsTM2KGdAAelqi1a0eojrzVAXSnMMjGmP6uDVIjjibsuQikZ
j/Z64H1Juu1ana2f2fw3VWIOqnvyXU2Q2IaZyMNnvYg0kTs2Nd2thmd0+lTK5V4t
HySckR/WZOFyMo2fQ2ULcg87pzTdmTixO6UDNzNRUoDOxKjfc2aZGJFslgeVxZz1
IToaEtkk3OhpfT34Fvvye6B5Oh31quKu56+mWhy2svsbZsU8S1/lxhOnVm1cM56u
iTO86INXsiHIsRYIyTFJbLeRFzbChKca7BOCsw2wC+Bk94p5Vcva24/c0OpXiuJQ
yTQeaNk9+2BpwY5phHKrINYFZL6D1/m/Xp5Q+5BHuP4amx/XN/6Trtj/EItxaZOC
s7LtbbFqhB+YPlw79aEy2t4poOq+o8XzxfnEyHoiqmZf/5R0F1B4Um5pIYmDIXRC
NsoGEooo5KBQS5nKxssXSgtZp5JwgUexk24bjvMEROMDrJzHNTjNRpPtVNMUSWne
b2MErCNilBHqfg7VSzhFDwgaO/g0dFF7wzOGPRPypBAbk7radpSQ/0DUaFhwV97I
bKXpQ+BUo//LHyNURO5CqHAeTw7UgYC4HLADUqb9/MvusLIdpVzCD+6GhPVG00af
+0cXq42ZQGoGLSRyYqnC9lJpJGqz7XE+TC6w86cUsPL4uAVFFk+t3a6iKBVne1n4
bNS/bdMEyfe5AhUI1KpcXqoBTSGPBZPG0ECtJx5zwxhI4Z/tbIbhvPAMCKAUts55
kcb2TM6+ig+Fp1+PyPLYNp2p+F6xlZyQcj8YRAhNYmNH26HE2lcecG7e3x4bNm9I
yY/nX1Y5WsF20RnzCV+jG80x4Sy5GhFIpi6ViGJXGl7ZqK4zyWaF+Qg+XmXxmAs1
8vykPRExnSahIIF4sbjBHPMxE82PERppm1dUW9jN83gkYMtmf9nAaOz0UBypyCLv
1DnZsRXddmxzIzm3VFoT0hvpddofcJJszCphDOw7kEi1WO6achRa6wlRezTpmO6l
KB7wM6kT6cAC6HC94aPPri8ZGGFggQLjcpRXZZHcWSS2uqvt8pDImGJu7wHg+/9o
vt3v7UZlJFLe8SxWy4rxvi31AbySgbIIzTbCfXdTfNV3cGxb4fhzhgvsk3f8r1ej
1kIoTQoFQ3TEkmf+1PO1mUktM9X8LT6gILV9Y+CDoLyTStYIrN2xkPDlvN4MWqrV
O+JdsoCMLY+BQY/oY8TlrtQF72XdXWa9dF0axjY+T18esHrehB4wPLp/GNJXKhBi
vuGFNI2qfoXBBTMp/EObkec3Hy1XFts03SR3cfzJ0nkHFI0Te5dKc4qPtQDib62Z
eQInN/p73OODx+Y7UJAVV72b78IjOvwDYLy/x6mrRvUnZbkwHU5ZB22AFkZ/Zdac
jOZvbTVmxbc+V5pCjB4aFYi+uMOJXNu9BUUHdYezEno8xgNdbmCP2Dps+jG/YQOz
Qy+TkjoBAZXoH9x5tgJTxFJEXO6nejEkkx7rR6ClvoKS2v44NkEM5xeKmuohyGi9
ljp7Oijtqs3ji5y6YG8mS4SPiuWRdXG8tsjtjLQnIeKYvWszdAjMY7oqfoSgEuGr
nxkowa9bn0bHzZ72t3L7/4b76I+4sQasV6xaSj1dr/dMzM1TwHSy5R/Y7rgOfUAE
gvTKciPHMsuaIgY/p/VVhfqEgyds6Ql5yjS0Ivf1bPBddQwHSe98pMm1u5vLte3v
WJ6X/gsL6BVpky3iQblg2AKa+FDF3/y1IIFoQKlDUtFI2v7sHGpmz5ExHDd/NIbF
mVyT5cIawlJtS2u5B/CQ504Xvt6FiEk+SkBV2+0WTYR8kLmZctEwJApMriSsi9PB
4XiAE0vnopbH/+rjV8fnrCCuiCWCdDxDn2vDYN1nZP/wfHRvalexTLj6g3MnYUwh
Dodc+7JPQXfS4HyrVzswSW/eS2jW9/0MPU6+/R51CoxPRRP5GcBMWOQolIp46aFq
bKbGeLvr2HsQrV0GYr+ig0uXkgEfWpQNuk5xS0hQHtZiuWYLoFW7ZlRL+tniROry
oWbaRGnvwVm/oTNCiCJA+jdVher6+pzuxebnB6bMp/JtvjiC7ZMYJH0NB7lNb4IL
sjHfbXOHBEAI3yFbOiqkCkP9jN8uROd4yDCPFOGJInw6cTJgRMMGzi6cZoHuSn5p
qYh0MD/2AO8F5Uz7CXed7rqvTjG0W+KTrtNe0RSQItgOWdgIPqPUEeKP/PxOP6od
1+vu61K9NsUOIgFoqBh4CI2wqLPFerRV7MhopW4y1KLsAGCG8DtZ9Ksu82Ur+etg
+MGCzSSOsJBVNT/uKoa3ceerZJkkj4JDCYBShc0mlM898P9GLodaBkpbZuoftB/m
+FyK2VTk2RfN7zqWJNWQ3XQ04QGZbgXj0xv4wYrVWI89qGFwE75xuCty9Z9aXQYU
4gyvXsS3T6gHf4yaC36AR2pjVD7msZ/7L5UX1kUPw/MfVlZEgHMoFbzGyA7ag1NO
JOYI3Fo2rO71uZRrT9S19MiUoQafqIScVE4d1ihgwpVrEtz9l7pRzvHaOlZtXz5T
9HdVFgve24Le26F7ml86xJ1M9bVRUhXTMoSYcYdhFtpLdrkeMglh3dBJLUHEquTb
xTMRSTil/WyCDpjS71hNfCLoidRC0mm8VIzohknEatTbshEy3CIkmsMmYMcHin75
W2rVsMvn27fcEQQjUIy/0VBbLi69Hhtji4X0j9IBUQ65MVDi6ImU+gAft89KLAcY
NvtEMciB/dNfnqV5S9eM6W8vvAhxWd6vf+p/eEU2fLqerBBlDqV8do7R2jvnt8f4
3KDLG8+ZRNh0VuqwvMuCZHiKsN8a4ZxF5SiiQSP9iqloWR24tI8SUCAtdsD4DKC1
ByZ9tbKHYdPEu0k+lc3iuW+qfMy0MdUIV6/A2esec11A9FmKAP7KmJOIO0pIxCTv
8/jvJgqiWTJjOAIagb0K+nUOWY5EGv5ut18UqIfDWOv5pDh6HICds/mpcgUN1jNl
0e4C2acLijZKofZY84orkysbFAmJpXMMlPh5cbbzvnSN7Qj/2lP6BlLEeGlmwVp9
dXiqfFQdygq8unaMJlcuUInvWsprPesY58P8YksnC+PJr2Y0+VsSFGZxA4T6FpDv
Pi2DLtfwaAQWlRmTBTywfzWi5vaUq9UryO2tS0Ho786M2l/M2etxSXUaJAEA7YfR
WSK30KeGj643ibE1tQ1mpo+iJ0DJ3kJy7vS0f/80g6iQxKqY6WTg06soF8p7L49g
ymtbC/HKIVWEYrH+98yIGe77tzxxopyEHs5gRv71rfCXlpiP8NR80Ft2qTgWPmHI
u6SKx95hpyVr9MI+V1elIgZI6nK1W1qrrK5lCa0l0txMSfZRkbPPt6ogWViY+T/p
aIxOg/oTDh3H2OnandVAdDq3BNufjyFmSs3ZXUd2NBXokAzMiWjiveLTlpmBXuqc
h4SUpB5Rl5fmO7TAeyn+E/8RL5nYVL/nZ61+Ape+Ra7/QykzEtUp5bzzx/MX6ehx
DpHOImqsuPzGlppCowZaa0TrcDsDRZWr3uTggMPe2ugjqqwXk+Mo7LLHDEdDtzI6
uRQVuzhgJaGq3eon2p2yph3/GKIpsScM/qJulESovJ9t0glhrr9tgHpYNyupKhRE
TqRZt/leyl5E850k9po0C255AKhLq+GIkXH3rDqdvrH0UW2HjK6PHB5mMgZ2XPwz
plPmFyfbuBCAZWLzYN8XxLaJRvL6XDl9DLExXWjzpVHC3HJmO88cBKIPZlkuwsxn
gRLPWPF5ISSYTAPKmSgqgOU7Mkg2lwytiqljP9CnfXi+3jOgyTucDmnK7TTG0HAw
agY33b3jm2pbRA55ZG1LKSn0EKFwE9F/ICLCsZz4DgPhtSLDyuEeBL3OJu5LlsbR
sB5Vw/20VJ0u8PZye+O7t4UbOsdjda93s9FBiNa3KPExP0dJmM6JVDVFlUertPvx
1QQBZxM/k/M4iGPQ38JMks37HdiwAPuyZIew0hhsVpM0x8O72s8F1hQUQGNLJ4qr
Y+u55nH0swdCrHwXQhYpyM/aArFMx/g8cq+MPQ3ooWdr/c9FhPWO8UDoiGOJomnK
/iBzAJIWoR+pJm/nI5PxwQAEkKnBDH5mBgzTnD6zJO573dGtZkPjLc89UEwa65o5
PL0nnZLx3ZaQ9JttonPlgCUDfGH4tPTRxGAB2ZuSWBICMRntFCcXPm89MI9yCOeB
JmzacPTKFcxYvjzitW7tYQf+uR0Zi+6rmD1kQ14dnYBE2A9gJpZIBGnUJl445VVW
mQ3RiBKUirC5R29c64ims6aEYXqvQ2f4a2P6sc8EzocDi1eVbL+P5ZAdVUWildAg
BHbCwUrw5KrmDZeDY/x6fl5NGtKOz9OHszwiT9fn7b1oilOSVWaCA7hy8LZxAt9m
3sxoOjCm7HD+tkKb0GSgtO72D2WDYzJVvK3P+U+1NxMZqXsXPKGw1TOSsh8m6O1m
/0dehGQF0lRJj6I06VZqX2dVRZZtdw5V9e2HJh6+/xKm4KsplLa3d+/KjmyA6LlB
sXNJVUAdi6L67UiT8wOUZQ6avIuat27ihmJH5Bg4LK0Nb+SUv8ni3LHQFBjQz9ar
IQCDRZpCoYk/nekhu2CrvdRgpJhhdeeLS2V0Gja2LX3x+CtAYf/yYdem8q/EhHTb
cmil7mg1BzfwNFrXTFb11KYQdB/qT8dRC9i0RtHVUmrZGElH/RwFcTC7LZOmta++
Ql6HhFY1bhO2c3ljMmmmpzNPOsWdg24KUxdOGSW1VqVVtfP6UoljduEeB7grgN8f
F8MlYdCLcn7u3BFfWW2xYWjITLjI0DMH5VTytl3hdcsMjtNehtEwxFTnHSl6hFri
tAAbxluVJBM8PUmeyivbDLE4CKSO1v/0RXSp0/OL9K/OCxbThrI3mkLcCy5Zsmpl
LB4pO302EGaD9jnrGKqxOTfDOt4IbJr4lcfzT2A/sBDB3Rqsf0pHdSR0o3uKCfqk
VXDBSeaZ88G3zpPUeUqIavldNcCpu66aERBox4bxmuuLPAEqO34ePKrkM5C3dOal
PiUL32gfQz737WzmI1fH65pWnvGjb9Y530OIUI2OH9RANB/4th31ZvwvU0Ov5ot+
CQrsuyURadfdWewS3OXqRsBL/PZw4H5NFESQrhg34DRqWz3f0fNkWmBVMRUjtvUp
RsMiHix8rzNE67UbAneFi8NMsh+SpgJbBV8oWSno5ZrCjiGXgzp/MzHpBLQW36Wf
BEDAYG1L9qb73jmW3oYKTX8Jz0802Dheasc3lNIwTLy0CMlVWTJBbKbVbYO9/s0K
/PFPa8W/Y+algiBgPNP9unz8BYweKTSx1o9FIZNyntaUqf9y7k27CTsT9s7nZulO
QqF2Glxlw38LYFWtihX7jR51c7IQDMP5KVV8zqSYoerQrdDn7xmPEJStKpv7qnd1
jCShNTM4NZ8G6nmY12bR3H7DJ4hiH/XmXTABt9WQkvMnJ1+DFr2EVdhz4hO5GmqY
4XE101fTR4VplTLuMbiJAAdNhArj5QawGs7wsQfWiyBnmpDA3In7kUgTlbqIA5jj
KpX3JSAbHAGApLJjtwaDFn19tImQ9LKDmdHXH61Wtmhn6WDTW5rMQYuZ/WCYJCbo
H84p6LUhfTowiWj1QDQ0mjNP18nAvmgYZXXpvK4IhnP4LkqB6GMuMh/AHVY02eKu
MTwB8T1lQuKGOG8LqBOP7KVN4AQpONDTZ4mbs4RN9bWL4UBS8rIVtUKMkldSD5GZ
VeCDbNo9KkUUgH8m/yQgVmNHkxG4723H99CDtW0ZzHXDSgexBlUKcTpwVCNRfOLv
jASs6P9MhyccGgv7KATHJlI7sgGMgpS5WM/0yY93hdYH5Zz6Hle2ZlJyR9YisWXx
X+8yk7TxeDXrwDhhk0y9kTBqvR9PAuWN9lnyXRN9Tbsonhrj8DTWShsMwK//cXj5
etFcMpI5GtBSFmDx/mudGH03ePxXP6bmQPFiqIiymVRhOZlfhDYWXm+GPHgn/K+2
NYM3PPYpV6c1/0sdebsqcf4ReeE02D1y+I3mQ+pXIi5SD8A8VD3D6EQV+c7tHdh9
GMLpXxOSUT07UW/PrnoB7DxndTvG42C8Sy1s6cJ907OzRyHErSlJrVK7UYDp6rO7
kA34mnPqJtYaLXh4l3F4ulzTjSP+xzwmphXOdlDJ72I53P2Yis5+AevzzXv8eNAm
yrGbtCRQHa247dDl3jwZfR1kK1FUCRwoUfd68Kb22mjfS5GVmSjhcYW4zGYg0A8k
/dixY4oZ3AmlDTBrl3f4JMRWMx6RdvPSYt4vjg7OhLQu3OKp9voNKNGjonRO2Lse
Ye1bk2NSyMlPoP6Q33FJ3nJjuh5GYR+wDkLjFVoQrnlYVMrR0LtU14NslVsuhq+b
yVQUjT9HqmS7Ss+DMA1PXO/KiYDcAygcIG+p/dO2nZLB95mnLhb7+FvxgI4doMvj
iFqA3ybRNX8itaFWW0Xu69cZwtJqj2wzVf36LWJe2A60ZQvpR06aQb3cwD0BVzlS
/QjxPZqogR5fk0ecraifQzoDyUM9li/kNiXI546TEZax901jaEueViNufqIcB431
cJ/pQ1/emCKbfI1xhgX4OaUB4uXFN36u8V9B32TMZgFTENF9JSlszxu5tXQbYrlx
XgPaQvTpcHWTUzd0nwTA/ObT05/YhCo6AN2A3844BLbJRZPNgdIIXzPNMKXJneEo
C548fMJL6e9nvQII2zRUqXaTtASwW9IlzQzNUoNkMzAABGil90zEyy8ZjaJE1mHI
dTeoISaT4AqvQBVuXmoiX2jfgp08ffApztBBbx6q4hX5ZuA2aimfMmUezvve/Svn
kdKdP494Emi9s+35NQijyM6U2wxg8H17cz6OaTaaBZtPA1BP1enk3JMbGqeuOFjM
K6+FHF7r1BSMWlBJH91DyR2dQkJZ4uslk0U0SXDwTJKd3bMaPQNC9ZBizedX1hI+
XxqTRjHQ1pn4h85AwjRXTp7POpE6cjaBPoAP0x++2LWp0vQkPM0HvWKguTunvlgz
BXNjtIImtOiCNTwxz2gtDanlMM0yXqqtBlCs3LmnMwKezbRSyJKtLNrP5xP/oKgi
fiGGVaOILI1HpIVBAGbIFXb+9Em6y9Qf4RhPzVtzBaWynu7iduHgwnsjDahaQdc4
QuNkPFJmxPFnQ7OLbhRc5hXADZpdfYCL3AWH5mDyKPBpG07YLBBQ/VsTXLfAm4nz
NpOxhlPkp7rUT6Cizg6bMtbpyCGQwIZB0iVjqgecYXtDjRYhUl/7X3rmUWMzTZSf
2rOjgNC0VqYyx5vWSVM22PrF/h0at+yytG6ebo9tLvxrisI8AbzQGfd99vPNsrFT
6hXUuPCVSTYJg/GwZJ7lkk+J1Fflmcs3UJ2se7ZqLkjYjQoKKzOEs+Hf7i/FA3lm
HF8YxqLGaIprnOj1thMrzdxWg5iEvILPhifQ3pXTzUN4pC9EAiyDdpDNxg3P8y8y
1RGiJofmzC4jxQAv03MMlJWPEdv27aw9/PnGeqzBWEOmCcnrfmIqhy1CR5oWellf
4zYFq+mUw4M6m3j7ltad2PBRWrKlms73uMzRQ06BkqFoOwqL66rVHMbR/ceLG0N1
cYwoGVomuQJzzVReE+6a0Wgat0AeAsvz7VhGZI9pJS1mNI9xIHMdQ7aQ6NQGJ0Hj
3wpNoqnX0FQ6TKOR+o1VXinOwSqE9F7nm0IEkbD63I8PPT+Fcu0+fspaM93DTJZF
zhd/TxyMioeZBQcyyaRTnzO8LZzpvMd7PWFpuOsRh0ivMmtNOYx/ZbSn4zsoMPJs
AsFl2otiiGdIPVFNBw/1+UWLLif8XekDYYp5aQahI2D+COXRWn4jJQoJLCYrR3U6
ISHzzZWyIJVW7JVqYpyIsHR46yXCkUJJXLlLZYnzBr+mRiCLSDoWhXh7ihzs9uQr
AItxtqw8fqgRQzhyrNmDJ8YH3dfA6/dWmGiOGbvq75TszTV6VXLkZRYDxLe9K0NT
vd+spjl95rYZDCmsCReBl1barciqVfjbkV1gLtgORiRGi6sugSrjz/66OHJOcsRp
nRYCnN/pleD/BEYwAedBOnVhjN22DHEdbQPqXFag8h2EZFBRKkPrgJWoTnpga2aR
tmEPh+/CViUAdWSrnaY2jfWnas3f2XS3KUIn/Wza38J5M1icGRLzqto2fXGvU/qF
UcJz8ypfuQyDaHZj1b6mAa+azjedwJqgOFuZ3L7ecovYpXl4TJk9V3q039vvQ4lV
qMoKdCdR+uTVJ53EtxEnZI4GaliMM5GuAi+SqeHeoEYHvX6OuczinHD2Qm8aSnvg
ySQpm1KZFY3PuHfY+m00rcmRJ7olqApRQag2UvgA5HNk6DTi3lr2zNOPeSjMyHgh
vJfRqotffA7A9Sq2O5YDa/bD+o2SuBMksn3zqM/qsI9W9W12GgXzZPYWN5vS8JKk
6SaMRRIBhlL+jl/u+3MWz6cYnAE37IsagSo/nWGaze63PJgg0JipMCFRQsUUkv7n
P7L2CULdzIqf6hW8ASI2htc6OuAO7ZPVVs6MauAuzGKQbmJjxRE3HYTQo1qNHLMG
hftiJXGFQpRbB0nDFytePSaprKoPDc+F7C7AxFkjtMv3u7e8gHexXuNv4Y1OQdbI
4w7hcWY3rZgkZCDFxMhEz8wXVgnVaDurkzo3RGsQfOFMNYZdiSUhJALAe4KsWfAd
Kd9EDw1CQZLLNVYZG6e8Kz4dIV6pDC/fq1E5xgJEIwRCmZ4PnFffReVI/jBWkKhp
e+8eVCiYF/HJgxPCq1+qdL/UdtUZPQz/jaJTtWgzhN/SiOLsu889YpMajoP+uXko
Pu84r1k57cCcZrA/7LNExhAhDdHW0tQLta8lv8U0XtpGXgwqVfYesyiB7IU/I+sm
0327jaBJOX/QRrZFN8Y9f9em2BHNxy8pwh8veg7Xv+e4xq6N5ILk0fLSGgQq4kIw
cFllDRbg23wIFa9497cO7tF+xIATVywQ7HBEx4HGIoasPyQVsBPsVZfiPRv8ldH4
+qYwqBWVkQrAvqYrMQKsMosoHXpLo+gpwhopnICUqegmu2hQPd0egYHlDdaZKPzu
sM3vGt9nYchV2+rjr9WFg/Jxlu8Gp0ACxD9JR9pJ7Ut/66rbcp6IBl7+w9bmmv4F
JEj6Ry+I7Av3Z71S5jojjFsfrnrFFxr8G0tgeTQ/NO1SddD8s8b4KSS7UA5A+w/k
WP+ybXIz/gXyJe1NPct5YMwghgMiJDs8qWmj76ztJG4fWD3RQfdmk6hbtKZNhW6y
GF2jPgYEv3qf9Hv2yno4HEpYYLwabZf/QfZJ6hn5UApcBRzAZsG1M6j9jlhZHwR7
cmXfAeVL7MqBk8Nz+RI91gxWxdtFHq6zTm1abwS/qJ0pJyClV0wMnvHFQUzaUECx
4X2b+/1VVlr7YGy3+lFtZgWQDQBN5hxbbI4Tc1nqT8Bvm7bwf7lxqPrDZnvJmTvJ
/4MswrNYcN5VKdGvTkXPCeGsYyXROFJi3S7SLROqZueYa+2Z3PVVj9u3e3QM/wnl
fXaXwozTgLfK0EzLg/d6fGnHf8EcxIb7rIAwMtnuIM8T4XVx92WM6t9A56b5QrYo
mVl8MUF4ofmT6oPf8jCGMVlThN+0r3IcRM/GgBQ6RUHVt+nDejzxZp4lo8AnQ6lM
WSaoW8OSmv6xjWKj3HOuaw9bNAGcw+yLBHm7NlBWLrf7QHOuIzeRN2e9i4M+IjGo
QA582jC/6URkxqg4hCRzhyvgitGMTOhcgmhdHl1AusHmFLCQ0RhOwgAyk7CS6UeD
jymVyKp/PhhdpLXN+MDnS4CBq6G/FZZwdDhKfWGoZw6u2IJjf0ODp6YDzlrMLy7o
7UZaxr2YKmjyq0MVn4eHoBF0MTCt2NzDR1Xl051fGF6N7NhJLa/Ab+JSRg7ihKAy
zYCXi5LpviVFUL9RrrH45qKJ9S9g+1SOKFag64ek9NpDfeosp7vFXc00Ur/pPele
ZZprblSjemq7ygleusxRcLvUFc+kwUd+hLuqCbnqVHp8kPWUI0+LQaZ4zn/37pcL
6863bMueAJW/Ja0h0lP4z6EP7cH+fXrwzVCRIsGugwA9MVv95B9jl+UvHmp/wXDK
FF7FE6+w7Xfi1yVZMwatg8tRc4T4tg3ztqEGhNn+U8Gybob4UyPiFfHKgK7q2yRy
8Iuh5Sy9DilfJDjnDorLsJHCnHS/liI8/YNY5iTGK5/35PbpB7PKijymEyi/r4AE
oeeLQerc5fRD6IofFqEfauL4f73RscqbwbjF+I85F6A0xR1BFljkWyoNyhVebCRP
b+18hsRbo/xScBnLYinh/KWY0/Wd3Y0JRADYVPAJZh2OqzUt0gA2MNMayhZxQSGo
S+yAN5z9nMIZ/l/gC9Ch7RyBoeyNwjvtNArZfXFHgjQeMpA2XW7pewKydYvaRFbD
HToe751B7o7RQSZJkQBCpPXx3IANS6J7V6yNfB3zVZ4fkxgM1Mx5Aazg6vF8/3du
zzqH9Ms29/cmpmUSnEPGytqJDNsT6ik/r9K/eu5fhE36iSgEfb9rZR/Z+OwIFIR2
AWOrv/+QPcWza827d3E804MIO735/g0HTpQ3xGxYNKZe/eO7mHvVHfrXK9wONRjO
bc8cSH1EnaMuFAsoZVKZszIKf2pwdlpUtNydzpV0IDarv2iqIHH5u3faV3JKtBa5
5qpIjwk+dFkBLnFjUte0qzfHoZqxHo/O5puB4GNi2rZBVPpjEj/60nyu9Zmc4J8+
cC0QzvY8R1yFEDBfvDWHzHjMwNPpVeMeOIq6CsKFgQsw0rewbm+osJ8TGspdkbPd
n5t7b43tSubz/n+Ca0LLowDAqkKXAEhrWJVH9x+S28Zbww0uu5S4J22SBo6KdEUF
Nr1jHVpT3LnAT3d7QebQqCo1YVMsiwlj610AoZ71HxvkQyA4gGdZP1XxCNkAq8xQ
Qp9hh+9LNA3A1SOO2ixtJ6fdxpNN/COiAf9aUWiLE1fiFOlf7w4o5h+cedFfKYRe
i3rsBRDbB+k8lGKq2UMhbqlIMRAI0yBuJv7rPE8RT721TagSxjs1JyuGkQT0B9qc
WXEB4VVR0xBSgSxeQopTlorz1s28XXI+jnfC+S/3yvbe390+yy7HV2PiP0JGlCbp
SLenlk24C9LF7XWglHOss4yVDzclnA8yZj/+8lqA6odRxqtX648jd8FqI9PEZdbo
uUSBYasdwr4vGdwL54oKUhP5t1Vl4hUQKusYDy/gXOo/J61OrAdYiy1O0b3RpGiO
jdlC4F0HdsfbcwyzcT1TNKFn1GxROKbiTjiKYrMRySFneqfYrEwjxvb4aayMZOLO
G+wSnwcP4FgqNSBxXy5dxTpUceDhP9f7LCj6nfXCGEhY30Yu60e8ssteR1e16u9t
L60eJdukA0riK/39iQXWr9jaPaiYPVaBcIhF9UnMC8W0tZFlOX9H8YpIKDISCSsL
EIVx5v0EylwdRGqy8V2HZOZ2otbnmwp/jjBXtjVlXEqvv1y8o9glbYbsyBhJha9B
kPXFPnM4srGlGj/UXnbF2ptCH8fmaSr5t4KIYzg7pbWNT+T5xNM/dW5SIyDTqf5H
GjIp/g7R99UNL29r8XS6fnhuaMwVfTgms7G+uGx96gwvt/xXbZnPTw61JHQ6TC60
lzZaJQHEH1/pOzEwtkWA/3vlZMhbNzk7z8hLyWazkLZ4ueWClVdGnM9EZNEfXMAH
U8Cd6A4XUBawc2P6c5wFCzojUD4qi4SzA7/Mx9FEsNUEXPvdIeLJCz2IFV3v5smE
rJSa9lQ8/oNnGipogK+eSYty8aH2bkbTKLvp4deM+LKk5XO6g1ldLeA6V6uGAEk7
EIQWEmi2DFU35jxf4HanPA0KOQFZfzf05Uzhws/iqsARgLq1GAMQZ8Hz4uEqAi5D
CCgObT0mn7GcPoMyRZadpBGUG05e3I69WZC9ix/ciVWXRcHeMvmCliq1tlrAtgRt
ZH9JFjzqv3nqydXdl+6pWwsRYuC1Y+wnALQ8Ff8PUso=
`protect END_PROTECTED
