`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvwDzuST9B5dXTYi2kjqcayNawfgxLWL8yINGBSfINWC1Mn2zmJ9wuqGHyy9zMjO
lYOg7ys0hhGKzbu4h5e3ew7uj0aM+SJl+vHZ9YES3SPUnH6LhGul9Vi1HnT5bIG1
ZKtKRF/YHfFicDSoYDtuX3v1fu/4egX77DR8qoAhphStCrSUhtzRnr4yCb+SOiL/
RB8sr0HvqSoqyHsk/b7t/5ZB/CjJpBmUdktCE1Ajy01Xex5G3oPc/VYg6nM9Ppdf
8AlLCPs05+YQuX5ugktpBml5OWKaowkDdj8X5n42+4wnOVM3QnDOJMCkV3y89lJg
cjwjkObthHKZA/U6BheiaKhRt76Ow4e/rQ1eG95SBZYp4asiag4Lo8sji4uAgmp1
eXJfTVBH4ii3l6TZjNDSva7Gkfe7ZxlWqtmhp1bvrNd5nbmWqE5CiMnR2rc6eNhY
mnPZtqxOGePc3RxnZDcj/W93lSYGzYAkMsr7duQlDfMx/0IW1J9SDKigbOZxYuUE
t7w+1S+g5nYhPVMEUBoVXEpSqVwtUByR1bDkAZj3fv604Io3q1Qegt2CMKW4bNcv
RvuauiuwElJRmrwNCf3Sr4VmWm+kF/eloB2iGpXb8vkBa+Q+t+24VufmfP0SCRXN
omqsSwxctQcou8Z/01bxbAX5xwn6hS58WHfQDzF4NiTQsn6XPuhNX+4daR0ITvgT
/o9jZTEa8qqJpp7R5J86m1bu2ZGEOx8AQNJFmr9tf57urp8RIRlKgh8XVMR2p4XO
LXw2/yXlqu4wjePSjZQXlZe73pZm7UPND0DtR10G19yW/7L+4H7SwpUt7zu1vFTN
n0ygH6HBPLcCV/aE02aIJqvLtvfBuVzAJ/rgiBv6SzwXSkPo9KF9M6l/0lbK0SQF
OUE5OBbGcuHb2f/AxA0XYbm9sgcYQvBsScsQw//DYKuYL+35h3c/uKVB+ocs617t
KODaQGMSC6Ujlz2x+JxypvLNxIRufXtOHCOlVm7124pdqIYScBwCzTYTDtD2DeBk
YP4k39ww6d5OsmWYfS0G4dK2uIA8dZymYc7pSnwlESSzWQgeb+rLCo7oBLIHd1bk
0BfgPSyUmCKRJkeYhumPaCSWkioWOpg7H7Uz2aVfM83pHTcJ3ohTtp9dKqvGQejL
vYfCgSKgE9WNX+256IJeODrKIYY0guVMQc5tLaVl43KPUaw2RvuiNkQv2N/Vjfje
udI+9bHh/lwfJIl49Aulw54UZPRjqEwmsKWCgp3+P+6hrocCBam2slmsqAIyDrwJ
v4vrxLme+GAfqIbrsjOgm96849ZfANCJjOhYiXHiEfHcHuQ/1b8sFxTwMjdPYrlV
IBy1wEgRmEQg9Pvyk5XHqYPSMDZ8VnO3wrwo6m7Vl/8nofAPMeq4qkywBevFYa5c
DfOMy6rTQiveMQvC1GLcMJnlB6AkvFy1kqvyuHYdcWfIbKm8IhxmtBp7wjwyU1Ei
oxeKRi5yk6N9oWq0lNySzYaVWH9QEfKR2VkYuX/7WcZ2mIaraVDsXXIm+TVMgtGL
yHqQjvtgNc6pQR5pQq1fJ8LSosUXds7DH373De+UOaB4Pqqo/Neu7ejN5kb4E9YL
UTVWEyvWCwGCjv2yhjIEdf6u015mTvXuZN1qZX8dpx+hQIMLhXrzKFp4Gx6+biuA
JB2Br6WumyvkE6HpNWQ0ucQSdBhM65NpUpXL1fuGd0TMBZFHMGNIJO2HkoOIoD51
+OSiWAlenJdqdMsxtZUqzki7SalRR0IZy452vvqATx4U9xk/mjvbywMFD8ck7dyd
W90RgRwP5L1vbZTOdpiQL0v4y7vpFH/nLWAUVCehuxCVaCvuxjf5xroBkU1uFBzr
Ie2YVv5oCg3IU+FqkQrxqP7Sd1UNvIn3ux9wVqj3H0I8nqbPYsvd0dGztQLkZrm6
7fE9ZYl3wsHYIb+5Du5/IIapdMiLttGMNviFb1x/7JpEBucbdZZzc6WeWtUn7ngh
KkitOTublvcG/C//GOaalSA8sjw2BCrjs3c5hyQSTfz55BfppGod323CxsF8464Q
l4AleAAAXwDh+o0M2pFSNJPsh6N/SjHbWvGiIQl9+TIMqNmirnnV4q8wRBBw7qul
yRtz3xsf+mYfogAQrjChEt/EQhsGp7/HdT7ajmzAAE29zTFkel5BQQPjax6HWkw8
XroPUNdbLkBTL674M575hjzk5lrWRqkiA1wkn2JOn0b3cP8fPQdQhetYZq7ZNqUb
SVID8YAu28W1L0OCqvVeesRYUM3daBJxy4CmOtd/gUwMwLhjePo7EgCBt3ep9JIV
e2loMwaV6xUdfv+DkDOPfTVzWHODdcBSDVWuXBHgFN8Sggg5QLDtjV9D4C4vuuYQ
BLaBSGDrnPotekpk98Zw4EJRz58KzSnyqYlFbW3xbZkT8j5Vq4HBK95tKKaAAbS3
MjEHJOmHgYnClMkS5N4b9+Yvs3zqk8WIXd7BWof/28sCu4YBeOnITFWV1juNmuXH
UAE4nGYuzXMWYfbl9ad9FR5pjoAlFTeVvwWUYg8ZpgEIvRAYndtAU0ld3b1Oj8fc
iihQ1BrBRpCI59OAXddjxmhQ3Yt8i32AcRVL9Zno1i+KiVV8Pd37kuZH3bVRJObL
hpRDX4PUtPRuiHidvNh1UlsUFQXTBAOXEW4d8g64x8CG1twYPc/ZiyG8xcv/KH2p
RVlzrn6CqgXIwFtQHOO/EJzHJh6OMvGTSFDsy2rPpm+P/7mByqVoGH2G6BxGp5MI
ypkfTJljf8hrjZl+g0Msv2PiKK8VBPDiRl0PHJ0bs38E41lqg7OOklSrbJpuiuNk
ZskxnTxnvh++flpTxOi+7ZcODzhnzSkySb7h02brHt4xGcDKtks8QuZWbm1eV647
m/uRKUspM5jB4o/DSwB0MnaZqgchV03vTAZd02OuH+7hURa0wuOIbJRXSj01ksNn
e7M88abQuZ36P8+fS3k8Es5xwJJJnFifkriqmgdQEuCYeqPquKayJT9pYCy/PGjQ
8Ha4i78Ucd+3xe0ziSQtbB2EvUdttY3Egz8GIg/LMxGS4v9ZjOA19cCpb4PsW19n
vQitPDeuLU1wh+mQLjPkVso87XuTaRwPBM+99nLqHkbTGdqU9Qyv39WwHhWeu62a
vK6Ybo0xgAGbA3A1JqCjNM3khqOHyDwNk3Pt9QZUnm181wO53JoqBnOOuSbTcbw9
6Meer/EoSB6Qs/Pl4tX33mi+K8b6DMfATSDUhPzs6SCvfP40hJu4p41ebdPKCZV8
F+Wkw3YINja3316HJsA2iybo5co3Va5EI9tUUyE8LpBf0FdD3R5M4sgE77FfYcdw
aAphDIrnBh/2iX3iga4EwBlnRoMbiCBVypTyG4V+IxYEm5IQAV1XsEUe+dRgtvrn
JPkX0SXMw6f1bzwZGufj3jr1qa6qjI8MkKZarNQhwpBDHCptjOKKO2pMYAMu5gnE
NQY23vd57zUkv5stIbvJXzu0dW0g2ehzvOpwE15W/+Ve8fi8e2CFS6u5ZKQ7pp3R
EL62rdZHLxrUCvNU7OWjek+Luu+xj6Gwnk57xstIim4K/vond4ZgaoKlMQr8/ACP
3h/clP0T1L6OGogw5kDXWRrVGRWkoZ0mzzkwyx6XE+2Ht5lzlQaVEgYr8yCVIbhj
vG4Obc6+QZT/2YC40bHH2MG/gvL0/svqV0FmY4Khnh92KIME9mfFtZOJiTOj66yY
vXtzvayFb/+YcdiXQTUEhw98bHfwvyqovydWtKxgIWwwivt9pJde5/EcyYkrbK16
rsgsIHtJ+LdXKw4CZtvDB25zrbCEzC+pmvfKf1nZJdZwo/58A08qH9RpZ+pSkcr8
oEAIv6P/XDzMIwhzhY4ke6KZ5clNj5mocPgS/YLX+YznP20z5pcvIPJ6OFmkPygc
BkoeS0my0Q8Q1JI1y+OJaK4QmqNSv5XuOF3zRSUcZRGyEGQvbF1+Gd0n+ZoTDFtm
lCvVOOdAXW9SLhlZflYBBRr2CbyEUopx8Ah8TzLMflUYEmgOGBJY/ViCJVFsh4J/
EbrnjBMLTcSQMAZk3AUPGsYePK0WCfEqN+JwdnYVrItJTQir5wVQexOZLWND6stf
jxeg2P3Yw9rz77jF2eK8rrbeGx2TW1hvuS8BaEUw3ifgCyiNqsu0D+DpnYEsWOF6
o2hl4ksukUHKqQI+W54jn/Tq2LhqNbfHWZU7HLAAqMkdlErAFLJg83MofBc5AS4P
2VXbHvOnX+Hn3soDxEG4atH+zAYDZedYq5ogJiFPgPXqhI4Jc12P3VEeyVRCMZQm
3iAeNkRMF5OQvSfpTJ9OqPvUaBtDxnAret6/y1gTPoRvwb4jN3r43LfxZvM38f/v
uPKabRcc/NJBi4H+8KmY4JTFamGORDl65BXveQqwuxNhTmg3k4g6+5EkD02KKBrG
+iqbR27lE1HNXMFZz1ty6exTnXJVOikt/VYG8MGjOnFGXdjfRC3K6E94ignITRdv
ElbsNd5zIHuMKgltfAY6d3lSWhtu5P3Z+CyaEtcOpI7M1y7eNL9GcZBv6ROEg5wt
iqXFtBtAg/AEeyJ4uZgSXIdJyvoBaeQYTJHLJ1rOG3+vNwhhSBnNR2iVvygvJQGL
ZaqeGhQ4Hm9dfebAVq6spHv6iWHHqemIqa5jDviFeYNIR8gJqLlxKLlpKB81I0Wu
/T07RrVzV8zSzuV6kLDxg/ewRF2UME+Gl3wikH4AIwFM6L9rE8wbSFyat6LQU0lq
fnCDBUF0YQzB+8jq69HzCYS4y7MCWMjUodf94ojcC/5Tw75/GbGOZfLdhnU3gC/Q
KzfXRAw1wNNAnaAu7R6tkUijUFs8oQJJLt0lIRjb3Kc1e9ZBVrtH1KA81tnsQyEL
jN4yeFKHweG3wREkvwmcP83gEGQxWQC46Uq4jYgMiyM/zl7RrH1RuJ9220ju5fCa
9YIUVFFmZx22Adxc3su7S6KzctC3A1WuefejwGuN3NIOOYGX12teNbl11gYuL/wF
nMUJJgKePoIDMcOJdOa8vfHKM9/fMhccHCyD3k4pjuzs2dMWkr13JjZ9YTuHW6LG
O7DDOwfvwC/zi7ViW8YZMWh/85XcvN9Bp5pdvzkY6vl4AGm0QWSTM+J4zLsHlR/m
a2PrfjMWRugxl93yZqhO88AZK6XsbxMnUktfsjqFbXVvkm+k+IlYltZoimi/LESJ
bzdy1l4aQ/Lf7jV5Tn8yz6vO5WRWhKawlQsf+V7C3NKqpN9adARsxToUt8euP4D9
xTFGCDsI0BfdRLeRF89PggYCxj0012DyQlL3Gi+PdJYnar0hOqa+Xqf6244xWwz/
PssVZDoOnispDpGuH2DH7Zz2nIKQ6lPbLDed07G30w9cx3L3mscP/VH/HLqoRQRH
c3ZHbKQFnWBp8NZ4egwHr82UCI7/jxP8fSpaxxaSMrn6CVQXh3v7GwxXNHaPzSwI
2cZdmlaV0ngyGSVfRcHlSpbP80HxRzayNTv2pamSOKtLnboWGqGQDqA27cfnzT4/
+nMfOTTKFT7QviJNAYP1RlQb7N/5r3CeIycCspih+uPF2hAGgKIeUxSSuzkEs2YC
1kAYf0+UThidRKjiiLT8EzpUmVSt3fiiX3d5c7E13kAAIHkiJSKMBRyCOYV6Aw0v
P8UmOaxbiTu1vnImWMjGqCSSkQavUNSN/XkFfneT/dvwppsYKMI/zvdoCPcKcEvY
ufnYFfSCglS9+JXyGwpxZex+h8HtCGRCEUttvD/s56mlMDHnnVfMs/FYwA6GVbX1
aBlZNBCtYIT3LICXDxTUPSxBC68qoqJqADb6ZkATZMDkTgxlME1kL9arozkph1oP
y1f2c3WKLvw6xPnzE/+3skZ4ylWGzLgfoCwPeqCajD2B3LhWUqIk1bR+g3gl8HII
09Fydod6S388MQvyRvQrVOTnBo9b4vI8jmhEEJED82lKR0b5fqf89X/qXdnHeo6f
Xk3xjvpH/Tk6T7p6XUN2eGzYSpRu6qBnD0g8nvAvO9v94VoSrWJGDK25078237ap
7+Nz/vpiDn7WbzUPFKZpK+SFBhT0MviwEHb0d+E2Ast/SEdJBnptrjjFPY2xK/1y
dgQCQEdlf4y4Eh4bnvdwEBSqlTvrvQOzf1PD0rh7SaSO3tj4ZYPp+VCJIhvjklbE
L81q1SirPArQs2XJccIrOauRGTN8z/1No76eXu5G3PyWHZbuF0C/PAk9pXfqOyVW
cU2ccT8OVMAUKtqDOdx9IzqZyXInad9cynfl+7EaFCQ6bpnbyDCFDn4+4P4ayw9x
VLMMcHPVHUgxRLFn40qj1baPZh5AN36z9sW4f98ZJzyEw+UtJg1JvXezYeJZukbA
7OQ2ubIXf8a2LjTqFa4COqCqNi/e1h1OM2PgHbjUSXBJYDPMgvQX2QekxzwI8xk2
hyK8pl+4+H9F4e2Cz+CnhoFrs1N7BanVThOPCq956quQaeEK4z3T+Ujqj78h7fhd
FRkG8HHwzCH/nxeYG0jZ5rIFzWRa7wogxOM1ZQcR4CYjKALwSy1LCuQEosf1Wyyw
SrMyrN7gRSWnHGjYzfAH7cJjRvLXLJu3iC3HI3Xero6GFIU7YnZehHJ78QsmzTDc
yUpqQJCFyH4RywbP3OGHRuadWq8Po5kx43heWmA/30r8KjP2m56fb7Uyu6RfUae+
/6aJVOILJGsAG3ZGpqDBDT2GuhtfYxkigPiyjavOy4ufWCnw/P/Km6woERPpk1ft
65az1Ng7/F7SMOi1IGsZAffMRrnzRDGZQ9Xyen5tT95JsCzmR1d2wsgvB2sBnAcT
rW4mVqD+HVqs5KVdz1fPpkszia0pzCFnZ6d3lvDre5DaX6zeIThIxVrU8/tA+k3m
IJ4QtEHXQwg0R+JYw2CfxKOo12OFQkcWI4wuxb5pGVLSJBu/L6SGoK7MOokTr4LY
utR/LnNjEZhxVu3pv1D3TiKmaycwUNubOScxtCMsbvpKkgNcG68+Bmhc8XzPkpf7
Hq9NcVFzNj3reTvpD3r8WTu6hI3c+rbwxEKsyWXmrZzPeNwrQdGXYVbOXkPF4cWe
7ZnzmayWTC+INcFZcOvceiTj6YXyxFb2qYh0dQymJmiNA7Fcw2rvPH587boBuKJ3
uQhQ7WOThWfa7onT12GKmckgPPt7/bnIoL3+Xf4UjCAEpi4rqinxvF17JKr4b060
j7FDHwaD2rxEXjYyW3Tujvsq0wrPlud0et8kRr7szcrQaU1UISUOgPilxyKbP6Ym
fWfQmP3PKnhCerRXF/8aI/2r2OKvA6apAWmYlSpK50Q=
`protect END_PROTECTED
