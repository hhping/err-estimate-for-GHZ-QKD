`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oN7OE7QTQGu7IuVoOGcjjWAqNowpg6wOUGt1ozB6OTlAusOTmPCZNWkxinaOEcXj
Kw7rXouYMQkegzb0iB0D5cojIoFI1dB6lnvECYXRIzJ2oufIA80GhTnnW/GpvyFa
LFpWl/O6+JTrXjYPvfdihlwFwnKBGhmztmetaeUBx/1R+/GJuVdb3bhGtj0C9dxe
F2E+/s+o/vgk/jLIpAqlSt8ft+c92Ox4pfjov92Ql3uF3+BgXUiYEJEFhbgjDolK
GyUDnZPJ/O5X/6qQFb+l2WiM2cofbpMpwfuqEPU3sHL6/Cwgixf1P+/7Kyu1P8HS
TxUxaJ+vxnvpTFrU/MhSHGcIUXc/LiC0g3YuiHLKG6Q5Sf0dSxJlYSNTVWZPWYVg
N6vznOjbh+b08Dx1SBQAGsDw42B39hvbd8HHtfKlrmeet1olxi4cQ764YkjpydDz
helcET4xjCr9jVMbHacCOsWOEefAAwOOCLag5WzQs4uRL7+I5INmp01S5ufO26lS
eZdRBMRd2K1cFNhMkOY2thQlXnrq2vcI39UuqZwUdNzcZ/9i31oFULTXpk3cnxDp
WsK8fEOOju8gyyEZ9lRPaVhSG9MtSIlyrxfde10GucV8OemtIQTFPCBwN4kKBxmZ
WrkL22oeNPP1g3g136oIqgoStmltUxXyfvYkWEB2yOfb8OzNRMnZ4UeuZsrAAEHu
lJ2mQA1ZluMJlVfvxgfA7hoXB9a9FmtNOjiBg2ogipO6XyFfAV+HaniiJl5RBjTW
mFZR5nO6xlDP007zeX5sJ1R5/xUSwMhk9C+iW0tM9E8ptHaKnrLf3Gc8dZNbhSuZ
gg0tV0FVGXqqZtwCYOS92ElNJVggoPz7U+Inf21lNr3Vp0jsIFbwrhKZ689NBAcY
+JZ8oNDhrXSLe0XYgMYyYvvYCt7wcO79WA97BZ5+EvNsw4Mh/xIu9e+YPWuKWNMQ
iK0pbU1jNysMcUurUdt8MYi1hZBiwT/OYqrpih+J4lY=
`protect END_PROTECTED
