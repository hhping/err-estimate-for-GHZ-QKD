`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnPqox/akPuXsk1Jpeh7gMIv+bhde+sXAQNzaL7X9wotoHbBX3yqzkaG7hKsHpCP
LngIT3hzT9UNFZF+d9skwm3Ul4xRKzfKb1ved/EznXZvqTqKDhSKZkz1pQtni5fe
MRU2PRIVrasevGQgqTHS1w402i5MWsjKuh1NWgDujRAq1VtEkQLnZe8Jg6++oKsQ
yxsKmXkdCfxr9M8psfZ8juKjOTwE4lT0HmVlLyP1LGbgO0kAC4dMOz9tm1smUMnS
Bvha0CoKOnwTtE9CZfOB9Mn1bYsmN9OEqtT/DdcZ6qWOXmF2lFT1wSLhy7ViuCCO
/yfvqL7S1TETB0j8nqZTBjAdnA9uyh7h/UruJfUhqwxt+AKl0HTGKFhHkDgRWEb7
y45IWktJBYw7YhuBshgC3+BzzH9q5I7hxUEGIjToayiOPdB2Ho96WO2MlFASmNnI
jNs8KbPlQPtxbNpc3ohaT4NTcwZcq/EXvpdhIgQBvz1l/ZLr9FQnygREYY7fy1pe
+DuOoD292Fy1rPRQAlQNorLLP70G9A/qwmXLgQgW2mFzWMpaQswhzXLd/LPy5ChC
TCWL5u8jyE6cQX2slkVJ24xrC77acYB8oNyE6MfcjpDvorv5ioe2Wx8TDk6eSClN
LMVfIK0SC1TpjE1kL39suENCG9IN+JEGVmTqtBfL0kkl1Ob54m9bS0qhskPRJYJ0
pkXInDi/PNCnnQEIWcDn+g==
`protect END_PROTECTED
