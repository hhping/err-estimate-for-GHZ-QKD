`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ax86G/UydbXKmwAmMB3WvU0xy+sucEFfv7nyCUIsqB5Z+3gyMMWQ2/LI4NK/RSsN
ZSf033HDvySqwPyA9w2TqXhKuGJs+ByYAz9kSU7otAoiuIY8dPgNl2O77sECf0x4
xQP1yMy4wrNrCaG5iV1F7UzKjuxfXHu0BdYZq0gMSsHGOPYlqkoSy6K1Rd/XyfdH
EDuJufU1V4f+DAIbYMqVNhp4xDnbuDIZ5eRRjYFOKZ8Q0TeDuUFmNk2jkFVDCo9d
GHA9vaqYMnkORJ2m9BGlKgTcpFF0QQrrvIaUIsNBrybXx4IxJr1f/cA2nVmcQ+zo
s8to612ZyFDBStE3MKCMwiY3Ynq+a8jUxx81XSogDAcOH/o0J2GojJ2iTgRqyZx4
kU826ith7Pg30RimzirmjqfW5k9nHbW2fZZ9vtnuzP3D6PEDt0qZdPZV0a5p2Oxp
lT1Qnuj0QctmEnEgPOHC5GHtKHhWTVc4UTM4bqVMRDmO7gDVDspjKB3GtLX3isMM
B0ugCtgwCvaSltTROFXRE5XMwiGedCpQPvVE7x8R/tddMDtwRSoXkAdEXRWZ/Zn6
17yG8SMaHW9poszAAa4m3X8D84yS+qxU6Yat+Pw+tmaxRjBa/S4fpMWi4DORKpDN
y0cTSoNGBfl031lvnmOy4d3xyRvQewjPEwrHgRGCtnDMqENau+npqPPOdUEITMrW
nFQVoIJs1uacvvrDGBEhpd2D8qqvZdcx5Zb5oUo1xtGf6XFDRNd+nu+DIfxVmaHW
AUb7r6YFI+8URWsCa3vcjrCWJ0wBM9O3mC2XwMkEtNJq9/EhbaZWhYo2gg9NAvP6
Y/K4MPBUhjdjIk7AZyPLIQhwbcWTL3yvnvpdad1fycnxnC3eIz93tmTTqNXdDFnk
2YNFiIFmLI13nsa2mhbrdfa94qSttDKMU6lpuUYvsG2UIiPppMGnngCGO0SD4Nid
/m+yxHRR9M+vlznkoduDsz80yrnTrYVZ8Fzapo8OJQ+RPhTwIKw+Y/5adk0GneYa
KvNX5h2+XJMy8nvpcYT0v0zaWHuKuRFt3whTF/law7DHNZTF9+8/Y92Qp3PYd7v5
`protect END_PROTECTED
