`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rafVIlwlNYiGo2rIehIUlOSyAGssdPTka9Vw2pnAWEiS2koH3XqouqeMGtR1Yna4
GhIOJRX3ogq8cFjJGF6rR+i24LQSY5syQzpAVDWZUqG/fIlf+VHuuMh0+ilKi9op
ifHV/E45RMlICi27TdN6vxHTVLIGZLsv1FMFkuAR7q4UJc0a0+HYcOpGJ2o8h0XT
Jd6SnTB1Yo1am0HH2hNDE9zSxtZZFkOFUZ/w5/VxnLzT5KOHPbD8KJVROBw6xj1S
GlBebNDQDuOnDZPEdrYzxcNNDx+dBhYg16ubZ70DC1vHtXzzwH9TrvHzX7jX1pIi
B4li/Gce6zlfYO9jG3qsdUSUROuH0kf0jjXpspvbA7LR4Lz3WOlcLNGycQ9c8jUd
J7pT3i3r0xZ9N1BnhZEZJSq0IgvijME0H5d+lXEr7iJr1s12GSHNomV0ieAcw75j
WMoV0Q4spnmWmdaG1bjBUdPTQ6h3tlK4+FIqhZzmjBOmL+UUdMDVR70KnoNipnMw
B3Qhp3a13EKAfom5lHot9JO6lL2XviIqJvSA1ACi9dt8uTSVktM7ntxl1eusT361
VVnCsqgj00E+kVeFXzaSVxn0ModYu2gQtEGnOEcWF9Z6SpMLXa9LHV01x6/pq17I
QpHkLzukwJORy9tPGzjpgAgnGWbg7OWwkdXAs8FWpVpsbMNoH1ghq/rcrP4XVsgu
PzuIlaNwgdqYcQY125Wjag==
`protect END_PROTECTED
