`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DkhiyjsFGginntQTu1I8ZhbbdfGzSeLIlqbS+B8WrYuFH1NBsByD6biSg5A/dEq
CAMP71l0Fynj0xeWzt3b89HOwLX5vrl+rbma4Sh0eep0q9/AEWSIKEJ9pbw3+aSZ
uI2GiJEJjBu30bJilX4ZTuGnDSj2TR0K8/KgzXpOXdusbToA9KOMf0nr8VIxtZ2O
mhNro3ftzarhj7//+v2l7sRoeCgZ95inoDgHdDJDB7U3urg/qlhJyRHfV9QmwoxX
YUqtgyQ4nq8HlyuedLyOQQ8lRnrhhenIpgSUzbCvQ63QdzzMfNmuBzc4uJJVjuCr
UQcjqIBnY1JcoLw+1kjAO/+F8PatwlshcCv/ranPA74V5TQ7EurCiRny2SrA3asp
ev3Fp7UEkCDGP7WgKfFZoCXN+tIEGWtrmKehRmnJuivE5KBXM3RBrJoaPMyvfHvn
guvEKYsFdma/db66aCSAEVZx0Y3uml/No0PLtTSiTjjKfitr/s2LSoZ2mQa91WQy
Mjv+pYMw92rCVxRm4iKTzZLAePeMt6ya55xoP4bRCTRZrlTWZnDLkHphky3jB39j
B0BA6ukkbptkDbFEbNmZZ9fp4UIrMvjXiZz18L33buE=
`protect END_PROTECTED
