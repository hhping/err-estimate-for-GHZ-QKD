`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y2OMjYMBGjKRqYsMpz9oakbm7jkdaajhs0j3Br5H1KGNdjAeWlKNR9plJbdIGuGK
MEMRsntMhseX3VIPNsYUJPj/7LMW2TwVDXutzA6zxudYAueP/Hw1yoIVZAAPqXXx
jV/tlOtWwfT6VgmqjqBIl9SYjLf2CCRcQUhXSwOobhcuyaG0lv7D2lKdV1AWcsvp
nAQ3P+EgIRAcv0OvZhSUkM5mN8lGWrhLKQh4+I1xdYUsmpfAUh3sUPmeVvoQjTqb
XOVvpJC0yhWdj6IwZc7CLpGjFPfVhXCRXkIc049Ds7vcYqzqTN5HkiIpbS1MWAZa
3u4IQVkBlNftYqb/K//tT1XAsUFp2Y7y9yPy1Ij4RTuFC6xobkh9iELtB6D+gtjV
vzJkSDU38M64TlLr69nLWV5KF5njLgILr9IZh2F7HqgtFK/WfLq9x2uSzWCMTgNF
Yk3L2sqH5NaZr7OwJXiCaQ==
`protect END_PROTECTED
