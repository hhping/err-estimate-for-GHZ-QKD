`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7iGsPyYT54EhpvGzOs3x4qeDQeJEfF+4nCl81XlHhRcppuvIckEP8U+6eREWmCtz
86/tS+Yv/PsGWSN8r6911d7vBZqw2KZuAFfhT7pX2QIjUAVsEuHxZcGF6D6jdWz+
yyYhIP9en46+kFnhl70rgCkvPHu2QRmFVxwa8IhSi4pc2MYSN5ee2cgBsLjnD0xB
ADAD0yVUkdpskN2/oL4GP15mnIf4qr+wBavqWqkifADvZWTHFftupNNqazpf5ocv
87smZ/HeeRBaLF6FIzo1MztD1aA9iyPNMqj5ydqB2sdxGNu/WukGMzCEdYb4MvRN
H7LC+4J9CRBTIIeIa8MZrrtK4Lw/JeP0i3H4v5QfhmfPBl6Ldo/77SoR4u7XzqDo
KZiZn+g6NJUXpZXQBvGiu/hqhFgj3HXSMGUfMReGy68KqxuSrPBYHQO6Hmc8xGjO
wSJQkZofhOcEz16maHoSlZ/0Rjc7gpYsfhchDFR4xKPaxWRRNN7LTHIZKRIKsFkN
GuLCztuOmSj+uFJlAPf6V86YqG1Q9KpYbTl3XltlY5P85QQB+tgWc2zy+vXf6uie
mWmuuqFgh+2jbLTiEn4fXIVemSv1EuR4vTjvumCkrZVmt/A7+VqirtDRDl/alqhN
lNKJ1t9TW/qSaTQPqWQFXGTZE5v0wsNRBC5V7JjQJGqUNDKV8HOjI09ntONcMgWd
OOjjO+1CBMPXdRFYOubOiK1A84P9H9W6IKQiQMcLeiCphjmaNluEm+rv0l99ajXl
oaibwt8joVjmiaN1+ZShWFmb0W5e2SL3mXZQzhs29B4oPqdah2RXt8FqaSkVzwex
u0VlbirsHfCRjRGo1YnB7nFkQXAqwf5+YxoTRvd+H3MomwDgzqODGJRPp83Z3YA1
eXD7Kp1KX/sFxYTFZi5OfINEi0QSOFzSsfAAl+8xLUeNEUNCgEzORupOU0AFEoC8
5YbQgYofPGoUZCEub1FrWbLiEvBH98maP8JwEsab1sFOrR8BW4yJJifrVlhl5KKP
N1V+HllbltFKUbhhfzq5cs0G6bcWJUO5czLE2k24TDqWVVIw5t/OTm33TLNi7T3A
VDlIIfAgFakFIEeDfk89KpObKllsxDy9QXZ/HGUFcVWKVpchnHdzbKd/szgvhJxz
Q+B1JMVyPJyrjTAS4PCeBRGo7xu+VKR9wSp3MK3tybRTnxB+frlnulAwaFNp4K1w
vQembZ95+z9smi0GM1nHmiJ4elG7KUS29BJaoL1cR1DCM9qCsJbaRncfoL1I7pbw
6uz+G4ZbL9tq9EPS7ovNu8WUEskXYDJhcx0JXuyjOvYPhMHVgnBQU4kkT3CyFIur
l1L7XlyDodYFmqP2/mqKDvLfVEvrSykRFj9hglfefmv5SerINlNcLa9qcUrx+IJU
BTDFr3CKYzxneIoyvIXzdmL0uTREUPArfnVsANabKSxmfWo9NRRu13+esO1pdCL0
gYchwH8XD4ud2OZ0Mm10k6EZztFk6EdlCK6Uupe4B5k27kH3p3Cj1OktJl6RKSYK
T8u/RLejsgfgMNeP29KJI7TQe3X6RsieeLx/k+diz1cc11Od3g0+YKWJR9TFfYPt
RYmyNPmRxreJTeQ6bzKqfn7goppEvje/hB5vyo7ZkC6Z+1hQoNrDr2dC4zK/MiZB
cUiepphfNPgqQQUQARnYULWIO0EmcUH+tZrvT+pvA/Frulmtme1pa3+xwQQg2JYl
vKKe8kZQ/Q7/MGVQZSqjC+hTrLBGo09I659ubgK4iauolSedzIcPZ+bAIQ4VpQjF
X1ttCP/LDCW09OBHa7QbFbFiDlI7h+H18UcGsWRyqgsdT65A9yhpNMR0HeQEkqEn
UFK6z9RTGD82cB84ElRNCoKk/vXI32MWu3tV+qSuWJ12S2IsXhJh4AoxrxzzcNFG
hQ0jhEKqxQcpq7n8ZUxkvA37oCa3aSdlxhT6KH1gXRAtU8lDbAYjuN/2W8yjBG5e
z2LQItZZynfBx/Lf/vFqQ42MBFW2lwm/8X4TWau41pd6CtXJ60c1HnB4Xpj2HfU4
Srp+oDUU/bgJEvKE3CCN30JIb0sDJhDcWgBbr1YMJWfF6e1+QYTo2nvz7mPr6J/N
33AOOjAnbUXLTTcXVjOnXWlRC6P+5f7VKyYD6vMTTFX4VVQGqK4TURrUgMX5ztVE
AyPn1RXlEEoSHZb1d72fg8q8yEZLllSKnjNwdKc7rq/aPZE7VUTsnwlz7L1rE+Cs
Cg1SSy8PDdgqngxkAv5L38Kbg1Olf7Lu6YKMOo+pkZQwHAI4Kr3Z6gT9VAlEs/9L
oloKOa7lOWK3nnbMkVyRfU9YP9PBZblwXrIl5ToGO/r7Tdkn+YVJaT7dUFKqnQW1
1sXzuMD+/CdKtIxi7fnX9TaJmNG97lrK+TNWKR+shbSLoPnoPCxQJ+xe0shShWh4
FspvfSJbZqyQhk2BCF+lcWGqw/Iv07KMqcCeGaMRAof3s7CweG7k5IO/qAwXyGVW
AYA+2np3+GGVVI/SJzO7pqOPdpwCKjtsKkV2Qi2RQDqS7OJCE2aRgXaRFPkvNnOi
L0Ozxx2fXygj680BYjAfoyr/FgRMV2qFg+vhrsvTOaTfvAzEuJk75sDGnCzTq4/T
FoG0ty7PS4LoBnxfGo6JGvMJZd0iRAjdrdTORp/3UA1RdVjB3zE8uL/tFsz/i5ES
hO/Vbl2L8rsc7yk+W0waGwGzkYtbnRV6akRbFrw3mFxm7jTY6EqVDMXqur17inVm
4mNdDKIWVRdo2eFwxN3MqwpZq4KG17a6kVqWH6ZNcolA0L1fcnVNWqhj6C5yQcsm
w0FsNc0xXrOxeXTAQHbqI5apitUZ1rCLvvzf7MKVdW+qqPY48I1AC4B22KmUgD/z
QBt1pANJLuV/B9dz0iao/YKmAUjPnLxx18zyOWfkJquI9LdCUt84r7etU/gwa4+f
xesgC58xfDpg0+++4emk7jT7q2fjiE8L4qmueJ1igQTVajV5UCURq+IT+giufk6y
WzBQOxzneGlCuPb6oiYr0trM8/hGAdxGn3PTWJ5nhSJFBR5fXEFFq/785PPB8/YZ
i0LcoIqu0PId80zdWGBc1UuQE4bC3S7wDNktTY3gZXa7dQZableSJsauh1FkEmuV
iDvXjltgYVSbcQF/qDHanQHYnRZ/ZS7oR9oGJKa0nIW7LRRrHS6qB/adMdbILUqs
RwprLhJYKerWo+7YEXco2pMjEQkDVdKuzqdNSDvi93m2YIBNfrW804PtvzjGZ2T7
1e4WEZHkcA01S5eCud783dAifLpJN8dWItr5yaKq5Wd6PpyVY/BZKMVftWEoAakK
qbJHMNlblsvL2jEwZ3XguNyuz8HtjePAVmsThshgx5gqDtPDvu3OXXEOYHIuWRPt
lhIFIUyGMZq7LiOUhP5wxGXziiXTX/WJppH1jE/py8RH7LACMWRHNc/oS6AcMr2f
vgIdbxz2wwWI2n+tESH9N9CYdZnfu0mQlN0tcdC4qQlsoOqSf3+ngh0YTeTfo6lF
6HR/P2GqQLepIYPUC+4s1PrZ4QEyqsrZDwlHliQyBtT2g3PMsCvZrIMP+AylGL/v
uKUOwuKxkBznJFTglrESRsq1v5KoAevs9t6/zupecIQH0wsaUggxXfDeThxtW4tn
N8qK521gbcjYuWC+X8E6CEyjN4TtfGFB0G4sKKeDXOwOLNTRS2USWeNoJpnn6a6e
9q0yio09GTzQeZzeTAOFcTsA2gl3TLpuODSncj+9cOazvn4dy1N9+sm9IFzmYvwP
iwXera1e7GL1mdk5WGfhh8u3xWcNmtY3adgCM/sXrFGGLJrD/BXZ43yaJlr4QL7V
F1f5FcpVkERvffFdxlAREcCA4F0TZ6sAFpFM4MhXGqFbzY37F6i3QWhneYtcOCHh
i0fWy/vHAklhBSergFlBwFgJvIziblapFmI36HK4nLpdJRLZd8+jydT5KcErfLgJ
8GDf9dN/xWe+53joaln+SM1bOB3HbHvGviu5O7K8/F1OgGeVc+rERAprxQybQ9VZ
rNBbgiYsbji6NVX1sEK1s9nWQH0PfJ5y4jV//OXD4IVYv0/Ub676vQr1yE7mmYR5
i/OpO435usBJQZReyqG5FyLlIRaOGXb9QTmsGH0OrgQlhse/UCwJThPc4NPtpcWP
WvrUECvGuQ1SuBXQLMLD/QOT95CQSmewEHea4k3QvG14LNTaXBK/euHU+eNBlBZi
79ur2uq7VWFNXmNKiB80fHo1jvfCfpf0zh2MgDJ9z3V0SHLpwoqgae/rFgmnh5IL
bA0ox+4erqVhsPv7es0PMkAAyVKu6MOa9XrmyNLiaKg=
`protect END_PROTECTED
