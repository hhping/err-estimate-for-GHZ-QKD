`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/gYQw15/R5WriZITjB5ptCp3K5JAXUOaT9V4enhYQGTnjV02smVPIqNYQGadzQ3
UMb5yOmpgGFe7FbfNb8a6zbhDQ70MHFgw69RivbMk2c9f6dh0o8OUgQQakIuzxy6
PGYLTRxd1BSQRvuBFAvVfep31qZEsz1DTnndXZm+wspz1EffS8IKIc+o8rdVvMeY
CB0bYDt88FnGb+t4n3sSVqwjH+YE7350dsOflORvri4P8w8ofNBhb3TU8Iju+Nkc
jtOvR0j670AFFtByPdTYXapJrsWQwDKaq93/NzYYq7TLrjs/iZCTGkqwEdc/T3h7
R3S4ytFXzK54EgMKvk4DNBjKzz0Xy8+Mi4MlgtL8dEAMDSAfgnWVgZQuG6B0ZEnX
E+4TVpd0icWGeyBGojMut+O53BRNJpSPnsAd5VKXLt4zgOimgWINKxbSlPlyS+zy
RZFzpPMY39MeorszNdrhMlrolVZRW6PlmICfhhR8qOQ23falIhkXTkafrcSWNq54
pBbNz2fNQRjWgGKAC3JBUOA5gvn+1S8eES/mpM7kzH6bLhF1/LtUDNATO3rxvpbw
j+3GqRieNYQV3rX24zwTuEtGQ6tCzpgmhRHwNSPaqlaNSFbi9SZ95geq/7EiFNmM
+LstehHGAlEwGTsOY89rrc6r93q2WbG898Kd0lvPAbhjz4DouOCmELYkmwyda6dJ
efT282LwMVqSax+CYDFQKyp++NLvDQGepph6vz/JXz0fzl2P5u99R/5LCzbQugKa
TFqptGM2wM6F4i2n4p5H7lvChZar9On9o3TZbVsZN8/wZQwAZSNW6AwYzZc0LHar
JCwuFRkEB+SxORehDZ9F7XeqqvRLvPYSMMmG9aEIYOcv4uOJj/WVBCefCWOq9ThX
eGlN7jyTaKhS/WHl9/k8uZ5iE4YLJKd5ssPIAUU7k11n0NYLGYzBTwgOizsOpyT7
G4xul4hxOG5WkfouLDHSvZJEFweuZOtRZ25Wlnlt4cm4050uPoHXKLCREVg7ezIR
h/RCObucY8glHBIz+f3TJupSHWdZAbFahjRIzJXDgaBoWgJlyhq3tfi9OLBG87D3
cBvZnzJTAqimJvenOco6HNLNI4A5Y9e1zsi2ZCztCn9KlPVrUNRJ48cgfR0hgJCN
9cn87I3f6GCKovfbRplHp4oOybQTSu6B88P/shYge1mUuLkbun/yT9wuHusgITXe
OZgnZ1yniC2SezzdJ0FwX8+zcjeRnnsz0hoCZ2rsE6XQwZSwT9KFSi1b7NjhHqVi
/QgFIc3SJ+emBnAclRVEaTNH9IyWCc/48wesJg+F4VH0lXIUhSTbZPsTKQBuG/QH
JANenmESYZs8dnJJ9NLg6G+CJOZkxPjiqobPOfWBPjM5oo9/5B65Ep4mlNiKbD57
nVpaYieigZcPgDW8sUbj2031iFvxV8TT8eThHjVodXk7xLKm0l5DBflO9m8toPBN
+rQwAqIqGPahvvL67KY0makbjpIZukX74h2MBC+5+gSS/nKyll993QaZWt+5mIbo
6aQ//hy7yrKPG579ResK3luNH8ePufgwfU8UnDivHoYjmhsz5a2lC/aa8x/0/teY
NmYfTqsCE2/GBHEOq8bSIrF/c+HYnHc0iJLqwcv9B4QRlu9u2zoj+pZVqg3v2MSX
v+o0lTzoV81qNoMikRVLxJFWvj3xHb4kBXwiYXy+VG2/TeTIXYdr18HVa9eKwd4I
RgeUE89tVPBJ12qyuu9EMb7qJQJDMBpuflbr26jb75+4aqR1NcAPKj5xHrnbBGtH
mworjRBNgCtY77IffO8FdtATqUAn0AL2LPpIeiaB38YtYYIdfQkyh+1cgIcHvH/e
m4ahHWJVEifZEboXohcko/zgvMsTX1x37MbawpXacMvXHevT4b6XNHNlmXXW94c4
HWYmyBuNf8T5wsBqGV7hiywc/9QmQs1xIR8BOA7hT8qwKLJ4CDnqsfCzd1f2kpBT
X0ctzgAmTIzIeJ1cMQOmvb/HuujI624hwPsClFuGfi3s3worb4HRpTP12Kht9ue2
m7YqwfqM6QTkTaFM72tPx+ZeVKYUyYuxBHCylost+JjuNFc5n2Ljp92fewLaYwak
Vmh/tnOhEMpDGO1tSLNRf0Dn0MfN9Z75aIMqXe4paro=
`protect END_PROTECTED
