`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OMARspv/d6Xp8r2S1NHSntE+3xmQZdxyPbQXrnm+BYCRcB2HKAijAaMfItwhzq3E
tpKtvihjAVI1Z+Obd4y8DumZfgMKgc2XYJJGdRMdHtUEEPXyapLoASXro9zFJRR4
MJW2rEoMw1eo7K2QHnILXw2KU7AujCHLCtAfrrNMu3L92MyzLpR1aXBc4JcUAmMn
1M/ES4ekNX52NMsE1yptDJ0IQhqsU/Mn9M/y0VmIjlFU1tnbYUs5WqSwTIjmTFkA
jE7CADs/B2B2gUB4MSl8YupjH4FBkykEWh6WDFJprAM7O6oWdXxZnHOamDMZaNHx
0GrRawjl1h2nWhhtlGMscj8/JFxqQrczhgn1YUF151Ycya8vw2lEa2kzJE+lNfeq
xBKQMExhuusdC3VYzNyNxoWpoZU8MWM+vUmzQoYLyC5EYtrZFL12Q3CuWaUjNlGM
Y81abFlZi2MHNhVLAk9nriiX+Ikbw8JBGnQUjgw3TfcnkTog/luw+Ia1yYhzQjSr
J1yVtkCpSIxiDZXbw/ZaDBR9JWERKfpc2EBIOWR7lsmrDUB0UQk/UltUzQfeJz7s
GmzSD7YeaaQ/VBkT4B+G3qYk7OttNkf7Oewmcu+ZrBubtV0of+OFDE54o37lnvmB
NyN/CUwsTPMdmUBMB4dKSAKdaoa/XPSUMSuiDQyjiepaHNw5VnuiA69ufgunCaik
kEyDvIBqeGHa2xif01Lm6zpmjx8sp5ecpH0udDIsv/SxAvahmE6pCfBmirSKlWgf
dKVutHKfkaVU9VT4v5pNltPE6ni/MtiU2PB8ig5wQUHf/SkcQjTE4E29eIotLF/x
7X5Gfwn0Sg4nRlS4jxVzWziHTLAoGsxzw34xmyvWR6v1VDE35BhXpwFNlAfSnCoq
nCLJ2fz3yS6rpm5Ep1NsXY9j4kN59kG3zOmbFNuU+utsVaNb6IMZra2nGIeFUsxD
EfLwK2QjnbSmfxxZIsZ2PqQJMl23ypyEgkSIAjomxYHh4PGiZV+/Sys14mHC++hE
2Lke5LW65C+LIQoszCff1F8FwELVRiSfWE7hz5BvQ9X4J2mojQ8CkgLJYtp+t4Ci
V1KOfzwNhzl/zs3QEq+81Vf1G+GEhXY0Nn6drAh33y7tQwO0M/Ya8bMJegQvo8Qx
aqdUryheLVpWzXOzVQJqeiAMJ30tGmHHOo9ecYcL04Q=
`protect END_PROTECTED
