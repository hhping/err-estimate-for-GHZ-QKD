`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXDw7lYsuRhNwb9dH+7wnjU7OggfL57KLBusChtmSc31ryRbaFHkwKWR1DsHIUiu
klYhQkmOnmX19w8Ca3+5yMA5QSnNPR6MsPwrI4bIReQbPaThrARfKLRUkGsT5b15
oVj4066wxbwSBjKejTFjVIH+UrziofaB+DTClcEps/UG7u0ibh6045TD+DDh8DDg
Sr0dFAo5NSKB/1DBjEggs0WuhS3t1NkRBlgB3nKyywZmIWeB/Wg2gxN+BPM77NZP
0+7rCNdKXI9jmP2J9+6AC4Vw3mHu6NbvfuzCSbCUmx9abwxEfiejSE8D4P9+JiL1
kVaJKKSIuAaNLs/J0ant9wVtLK0wfd8Ut8lsAmSP0vea+wd/VmIVIpfkdz3RrrID
fRmoTv+WN64sQi1zIVbztEgO88owwJtlz3/TPcM5c9az3n8jd2ZAzEJKc4u0/LsW
cWYEu6jiRuOcfeW0GpS5fxZtIiCopBxfhE+ya7Z9aUPfYnl0iM8y7ZdgfijZO3DI
Ohp+NJFtkpvdbHZxsWgT3GSUXoHCVNI11gnoXiXJ0LNlDklDdKIaviEVQiqsJiOD
gf29/pPb/X2hDNxshvMGwmYQ1yeN2eoxl6hWVykELnhsZtgK1CBE/dJxfe4mhgM2
1fCpkZ2KRXmAfu3lHex6OFzxZVahxvLdvnBQARRIHdp5xGpeI1+uM8h8g5SXwG4S
4zFWdsfqqdvtHxmIYhYq4ZfdVOhGgFI0BVR+6LpfycXiDIvUthydUw+7c0L0nPAW
MUs02wbl31sEhC/WzNoTud4s9XcHUm3kImYA9OgV7H+mW6QFNfWegsbd6HCWi9wl
Hz7eZzMQQ+2jFUZwbsYaRADC+XLsv74BGxvYBY5yRMo1mZjnvlnnEx1SqCv9iBjz
1UNlY7UCKEGrYCy83SZ03zbSBKAsMTNV8a1qFfVvBVECy43xLYrv6fpu+ecDcb4w
3hHfXDYbPmJk9ItqvMmtLS8eLkemalOpKIVlTH1BqK5uGbei/b6Ram1g4+gO/vPE
i03TdUrVqwJCzzPrPAYsXV6xPLB3o4e8xOcx2IFeuMhFMe4OzS27kMrAEOhx004x
HUp+KziE8tenXq6b5rNHxzSTrJh84Y6z03HQoIcLlUzbBpKGF+ODPhJovBWxI3HB
of5Wx6s8jFzpNNhJmzjbfeEhIiXr9gBt8XFlkLR5ANtn5euoW64N66lkl/ZuqZzN
uiwZOGCotmWDjt5QVQNSHzqHSYT8s8ZawpKZyXAu0vG5mZmeFvrCN1KCOastEw4Y
dFrvpydLngU4boGW6rGQrIqdKpuUnc+ja07AB8wfhpbSxNYreqC/oNw2hAz3WWlA
EEH+8ja+2FymfwiGXaZamDeKoKz3gc3wUspK1wx+VaBBkHJ2U7Wv6KN+SzMCr8l9
PJHLTH/LKUkB5P8detFfP7Um/XvOiMDVMrrYdRWW+e5NwzmqNNxiawa8w+Pke8i+
NUpU+K+puGt12aLq4nbMOJYCviB8cKpUWD6i1Q60YZW/PHZX74gDTLY5WGVGT0E+
QVuDbs63KVoFpC82rcEdCbJ0p4yb+Y0R9a67MKZcpxQyDRgZmG4UBXb5oocuq00L
j49vPgY7uv3xmEKEtXqagr3K/KoNuWSuWeKluqwsyiDInvrxYsI4o0vpQV+4kvt3
Wf9zUzH7IUlXiJrCNRW4qQUbOFXvR9gjuNYjEhzbRNA0tpcPGtP9EvLdT7w2GmgV
sHg0ORsu5G60yM661oHUNElf1Z5GXLMk4jj96xqKXd1nSf9nHfkNVBvhT4s00NzV
AhY48Ve8ZJwJ2KYQEKcdQOm9C5HoEdjEwPvET0LPIQWZwLdDEVCyiVk6E1nfiyrR
TaTKtDDYQjHYLkcARgVt02fpSNXB3bruImROoCSeAaCOLHRn8CnVsXn+f9hjPHvM
aFnGIAcxJuEgqMb5aRR5E3/w5POPaKSnXyLlneYgJEF6ThZ5AuP3ODPDXoKYIHLT
HcUmIhRcxwSvioV6Jq9ywZTkPWtoqEjdIQJcevIwDoSbGtxqEcYjBvP6V0Xd8gul
ueiqFsrx3OCG1cQzRMhdb76ZhJaSJTdqDUJW/4JLwN+y5ROYPzmqgU1soQeDVvy3
3VASV2mAwpaPqKA3x+s4fKBcPE66rN+QL3Xw+z6rbrCm/Gb6oytkPZ2TMdx65/u5
woSiy+zRiXI3OcGw4yJnYz77XZl3ZEAOeiUDwFqKDRSbNplfAS7f2hVif1C8vHbn
uAUEedkFutwmAvAEhjGFWqznIZ6SdNMpspFENPkBqW4M5pWnMeKvvKMEVdi7czCy
vanKtTGkq49CW9y+kBunYzp1RZ7qfYOGft/dVbLNa702N47JqBJgSgs3x+Qzbbud
T9yhySIWpPlgB9HpNDYCZOQNord7O0PoBAt9oUCQ5i1ZVEX7PTBuEzyVIpQab0QM
mgfwM6Z/rf7Xd2viqj9fm/0zZ4F+i9RUl5OxQEEX7/qbD/0IDa6NDR265dESUB4T
edlebvLOp3wdfjVHLCjvBB8ULwqbo7tZkJ0G72gqd3+wF6UjptpXEcQ4C8JgCYSj
2+JVrVmtrCp34MNi7aGRbw6WUH3ueBP4ohZQbo9mWZiLtvCBA1OB0mhYD9D3Oqxv
phLzMgwwt+J+cCIh2BvsyNweHFstV9Dwb/eK20lREpknICQBHv9th/LpBHzfzbr4
Kx6eMnMk4x72gS4a0V/Uj1aJa7WJNz8sAg5plZnorFl/J1VbaltwHAZDC/N3eSv8
OGt5oAW0NNWoztYYnSAdfrHyB7kosFL+9C95hXvraPiVOqiy+YWeCpLXusgzBxDl
MT9X3sb/pyaJg/sVHEkg1QSOqobFFTN+1sS3ApTtrdOwNytbEMcQDJDXe5mXdR+3
pBz+WgScp1SLIlCkdh08NNQWBQA2QnpqgLtRcC76ZR0UcgyE81+6BxAq7ps8rsnB
K5X6wNdeXmdXlcTs+5iw1Bfz7Q/3GTEu86EgS8xCXj8XUL3B3SIuBQ/QEtaK1VEw
N9+QmLwE07p71U+GuFwE3OFXVrESASJ1iuixTDKQeWz/8CRMR6/2Gl9m5U13/cDK
UJ54rWcrlCh67SidmNjqwTCGKt1Jy6CwmqaGqRu2H0Zg2aT2bubYU2vLgNDRYqTX
KUsOsbkM56c9of/VRq8KSqSE2qaK0pNe/a8y/lKXvOgzPmL7xrVxhmtLKEN+60Sy
2RyJaujQIFW4RGxvMfi2C06dCHdwZRPcCslZzR5ZhJwNVSrEjRFhKdmaLRIeqkKF
yYXXWhamdBq1Y8VBAUVS0mfjRbB3os7csdVBMgz+mVf+6u1CixXyVz0DNrr6bns4
BULn+roTDtdxI4IwpZLH/pWXMnzHM7Jwb8hslmVgBzaVlGl4R19iedwRTQNqkRAU
OgcgNaJ244WXxJdElHlx3scfd173Pz5/3JrmPptKFA6BSUmjGz/RqvMQ1Os/F7Yj
c8qHGncIPUt0TzA601sIAIkbgAzmIkUW2yAsuTcKKMciF5DzdeA/QlyKhifsUD+g
ebph5iMiWCpMmIZIO3oc+Fs1EV5u3y9WwCuw2+CEq6jOcLs7wnnTGay9Uy27mE8w
suKlBHkb35nzXnCaJEYKZSe3aEEvT0352Cf4clY9H208zi75roZFAJ9jCFyhl/+0
Bu2Apoi2el4rFZEmfddJnWXI1UM+GO7naFs/eRGBUPf0aYeLQ7HqnrbSSFItD7tF
UiZisY3FphLbMJtiFbyuklO5gtThyDRNiNBvVRp3LI/DYtlqS+l7IGDWAau87gds
LyAwktPJZV4+3c7FWRQnEWuTNQpafP7DwzWnY5br/oWEMmxSkRU+nh5YnXYV6+nu
cvFRTvzAqbnYWE0wYsULUAPlbCe4tdsME0q7qjuDIFK6MF6TLKzCnb1U4URWdSMS
IXBXABRWmkIA4yo01fB5Qgq1wi9DZpbyeYNz1+Agmo7p0wfJ2iJga6lwZaszmVb6
lZHdxRDB4xrTdmA+fqbMGr2gub9zj8J1kdyjEhh6ykJM/rl3Y4TmTjWnjzDAmN8t
eLF3iZOUs1yUL3GxgVlev/ph9ErtZ88r4k64BPQOPIpFDm+guw/uaP+vKTR7S6OA
/LEtfnMds+w3OffeeLpY/yiwTRcoQ68BSGl4eDalQjL6Cj+h5s8ljbboGrlB+zJb
xU5Ciozl2bJE0HhIgNyjGqNFpMUsy3Dh+QpsVZqAKZcDBUYfM4yloRJs5kpsrinB
HVywTp6a1Syenikj54Tb/z32eouFvRE/ObGkpD26cGpLfp8AsE1/7TbBn8OWyuNE
tmIvD2uxxcWwMGRg9g8cZjIN3zAgmOiY0MPr2rgyUinuQBnWlPmBosaMZnZ61pqK
HLFirDHBTQcMy1xLbHyWU1h4/xvmf1qKRR8mft7vUWs8KQEZreMesDrnNDrvKXfp
vlH3T9XaxkdWKF8/Pr2by4hqLqguvyrLCnpYvu2SrJ0pptZnhdpnwMsvI0Ev2Q9s
KT7InNzb4cZsdb6XCUCYCWhgzUPOxunxdquwsjtetzZDy+FUL9Lq4ukOAncjgOaC
vtGXLl+XeTKI1giO3TOby9Moz3iqGjy3HDfY/ZWC85vaJBio0DjokEMmVHucFipN
oS6R0USqCz02rFKjGxZOg5QEhXJppCtYropJBNFn/G9u2i9B75cmaYzszeDRPVPs
HclJ/vVT8LkeEkstC4O+lDywIYstTJ+4SVdy0Ko8KRhyH2J6Mnzhb57bC5jFgm18
odH6iNEawaCd9q38cU1IcI6ZzuJ+8yPinCEaj9Wvf7/0PK626ppXgUeIJ+tlhrni
4YwVVEW+c57eejJZ3OSkiHhBTa1jAWRNnNCzhAeOmcVBO/RQM02EE6xLBWKZ8I5k
CPciGlgwuJMoldfvHgDyCBRZ2aqAU1lBOt1QreSJ5wcPgkQDbQJ6P8BWDCZ4/oNC
nobIx9QO1vNFs9OJCR4wrGtbH2x7jy+NhDwKr7nv0o4xehLVKHbuC7N55KBGHZL+
zMXV1C/L0vXQ/KIHfB/mLJxsI5YF/66AmkHffzc+c++nDSGRJk7ZajI3XhCZy6MQ
ICjYNYqnPAXuVa9Ufki8svmggRjQJKAP6HY2hdrmD/gGNMEVgnfvODRVyjNcGQP+
VgnlFw+1vNmtqhj57fmSW+SSfUSc+EcH/hbSHtuP6SiMUKinwz22nZK75YqRrES3
nKxwpbavIV/bjLxE3Wl3A5cppqu5EjLbIYnMEAEOi+k2IZHZnAdwkQ2pm3m3TvUo
T5e9lQuhGEmVWOz/gjED5rWkHKscK8p2q1pqEQqtMPmUBs9beH11/50vjmDzV51q
Q1Z88Xgr5EGJpBfT0GSdIYYTqX3PuYa/zApw6rucDZbjUra3YuoT4xaWAmnx1SnL
QH82PYJmSvya4nqyzONEgo9cu53QeufCo/+ywxMnBuJgpWLg1P8U8/mk649r3j3G
0CI3fvKFFnZsIpQ8RT4XPY2Que97Lhksguv1TI23GdLY8RKdk/Hd20EV9NUotXcF
5a+PLmCTccgATY5Gtmb/wABs8Pvtt39YPTVRW/sXhOCgEyfT0s3sfQLrFLmjfl4b
Y1kKOTVLCXH3ZvpozynYliyxI7muNtXBYJy7LvPJ220a78z0c5LlM/vEtMyV4pjj
QOphQ3WIZzgCJZaCl5KBFUzkc1ZFYX9pBODyhc7VStMwWejrFK5vA8HEwjqWwv+X
mtHU4wcGVoa2iZfhBw/NyTeZBX+OapVomoBJPK18T1RUEB5gU/YhDyUVsQIdHs9h
kfUiVvdxNbsSnEDTomqDiK0rT5YqRQHrJ8GMGlUBLqHDByNCikIf1UzcS3jHehK3
tYFQdmBW3ST9dpsWpRMFn4/OTykYkY35kORi4DkmjR3qOhcOAyUvvMGHPo25tBun
EhfPXr4smiqbz5hDvGxnTD4Hv8n7jHOo14KCtbYgOe9QRBjVdchkqLsHi+JkhP26
uiQ83kkBIeO5EM3HugwFi+RK77GSZ6WxUsO4pn3aDMt5RJRVCK5QzZRFDeHWjZ2b
Sr0lmolhgNsRWkVCfqmpbLDfuMc8ckzmQtvQD/gUyM5iL/IrwPG+Cd8kguL1Ozk9
m264Ip85FvwLZQnfeNqs4rT5qmg4W5Jrt5pV+Uep8OcK4TZ2A1XtvJpji5QIpnpS
24Yfd36FviGg2c6voIgJcQ03BDoeafbXq1TCyF9l60WFoRJXOe/XIwGQ3cLwl6bz
I119qdZAiAzyGjAV9l9mL5NJAC7leGiWsN+OE5pLrG2O0RppaSl1JjMT02OoDx8t
KnkbHPp9irfYrX83OPULdnkv3ixpzTvDzLjihCycnlAL39OICAtQ0oFaYR3L0j4U
`protect END_PROTECTED
