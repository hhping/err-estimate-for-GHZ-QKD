`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MpKQjByE0lyVsMAZzb4uldruP/hrujOzPUa0mCMbu4HNjkYtf80nWE9tXUgOIbQ8
pr3viy+6B9ofEQM9nv8ev2Lbon+8fI0XDm5rsIDSJVvWUgzzsUJUCKVs97jzFLnE
5y+EQoJfSgReXrmlzAlYt0WIc2idgj6gwMOZEOJBrGL8JVKI36IwCy2JrtV+/Qyd
KLXgmZ3A78rRALKcRWm9wEMu22C0DGg4rsyWLxtRrcCbPi0CzV4ZrEzeheFR7/ut
GWfUUxFbdFDTQ9dv0CcFvvx+r1VGRQeTGtAVvLhE/y8Xq1M4Ve7k+crEimUCu7PV
Cx4xaiSDQAgkIi1Go/6FpcLDXYfeeB9hAZVaLbyn8lYCTCNJ9peANoojR7TCAAbY
M2vgkzKO6I27MUqosXvZ2chgr9RzfiuE+hTpFQ9M4JR+Bca8pgCtBcfp84Q9Ymgp
bqtSJjW18VE8s2Na5BLgSqu1T2dPXf0+XTIi53NQfrrfzsBjKjErL46SiRvSlu+k
1EpVkoc5feUBwqb8f8cYFLwYnWZvBp2dYXH2Hve494B1BqlgRU2tl3/ILkTwsFsX
wU1pmE/hFdvzn73HqDuCVQQeyY9puL16PtDXXMQMB6C9h/MekOlPTr+/7L3qIqx4
DojAu2gjXhEuguNC4obreot5ebPsqi5zCPIlOxDxPrASt6wa2NuYy/KZk4AaMAz7
2CCKMlhRRezLsfnFhaJihndgkVh9PNsxZ3w3/O5JTNB/A9LovG1+WASL12B8iSsp
3+GxDVr3wdt556IYJ0msaA6c3u0G87/Qrs7Gfo/itFGlPd1+aDlEo7D8fqBl6tKj
j+wifYqL/LGnh7y8mUxsizdJ6tK9eNd5HuQ514Jrm1y5dtGFDayFZeMGz2mFF1jq
TeR7JaF/k9/YoqMrkgtGYh+z7PGuOD8S77VGfZuYpTiayisepLMBRqbIrmYLTMRK
jfOQYRKdQCRBhWNhj5hCkliJq9gS8mPuMwPKeVoSt74JiPBMVc4D4dU+BHDKtVZE
t7ESzZbrP2cSrBSeVwvDYREqaKQfjKeKKXhDa7Z7WNPEBAViq4a+Jzb1Mj8twihe
kiI7qAbX1GP3Y5USFZPqK3/a7Ao0dygUeOHWj6GrwHKABigMF4sdru1DAJu+MV5W
jTwSRmnVVq5Nbbwy4N7HX/4Mxx8kksuwxH01O+WqHfemSkjWoD8dDe8o1GJnQn+I
/PdtUU6WIb/pDrJcTrqLY1lp/ukEgw7aBOiFhEnF9uw=
`protect END_PROTECTED
