library verilog;
use verilog.vl_types.all;
entity twentynm_io_12_lane is
    generic(
        phy_clk_phs_freq: integer := 1000;
        mode_rate_in    : string  := "in_rate_1_4";
        mode_rate_out   : string  := "out_rate_full";
        pipe_latency    : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rd_valid_delay  : vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dqs_enable_delay: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        phy_clk_sel     : integer := 0;
        dqs_lgc_dqs_b_en: string  := "false";
        pin_0_initial_out: string  := "initial_out_z";
        pin_0_mode_ddr  : string  := "mode_ddr";
        pin_0_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_0_oct_mode  : string  := "static_off";
        pin_0_data_in_mode: string  := "disabled";
        pin_1_initial_out: string  := "initial_out_z";
        pin_1_mode_ddr  : string  := "mode_ddr";
        pin_1_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_1_oct_mode  : string  := "static_off";
        pin_1_data_in_mode: string  := "disabled";
        pin_2_initial_out: string  := "initial_out_z";
        pin_2_mode_ddr  : string  := "mode_ddr";
        pin_2_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_2_oct_mode  : string  := "static_off";
        pin_2_data_in_mode: string  := "disabled";
        pin_3_initial_out: string  := "initial_out_z";
        pin_3_mode_ddr  : string  := "mode_ddr";
        pin_3_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_3_oct_mode  : string  := "static_off";
        pin_3_data_in_mode: string  := "disabled";
        pin_4_initial_out: string  := "initial_out_z";
        pin_4_mode_ddr  : string  := "mode_ddr";
        pin_4_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_4_oct_mode  : string  := "static_off";
        pin_4_data_in_mode: string  := "disabled";
        pin_5_initial_out: string  := "initial_out_z";
        pin_5_mode_ddr  : string  := "mode_ddr";
        pin_5_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_5_oct_mode  : string  := "static_off";
        pin_5_data_in_mode: string  := "disabled";
        pin_6_initial_out: string  := "initial_out_z";
        pin_6_mode_ddr  : string  := "mode_ddr";
        pin_6_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_6_oct_mode  : string  := "static_off";
        pin_6_data_in_mode: string  := "disabled";
        pin_7_initial_out: string  := "initial_out_z";
        pin_7_mode_ddr  : string  := "mode_ddr";
        pin_7_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_7_oct_mode  : string  := "static_off";
        pin_7_data_in_mode: string  := "disabled";
        pin_8_initial_out: string  := "initial_out_z";
        pin_8_mode_ddr  : string  := "mode_ddr";
        pin_8_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_8_oct_mode  : string  := "static_off";
        pin_8_data_in_mode: string  := "disabled";
        pin_9_initial_out: string  := "initial_out_z";
        pin_9_mode_ddr  : string  := "mode_ddr";
        pin_9_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_9_oct_mode  : string  := "static_off";
        pin_9_data_in_mode: string  := "disabled";
        pin_10_initial_out: string  := "initial_out_z";
        pin_10_mode_ddr : string  := "mode_ddr";
        pin_10_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_10_oct_mode : string  := "static_off";
        pin_10_data_in_mode: string  := "disabled";
        pin_11_initial_out: string  := "initial_out_z";
        pin_11_mode_ddr : string  := "mode_ddr";
        pin_11_output_phase: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pin_11_oct_mode : string  := "static_off";
        pin_11_data_in_mode: string  := "disabled";
        avl_base_addr   : vl_logic_vector(8 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        avl_ena         : string  := "false";
        db_hmc_or_core  : string  := "core";
        db_dbi_sel      : integer := 0;
        db_dbi_wr_en    : string  := "false";
        db_dbi_rd_en    : string  := "false";
        db_crc_dq0      : integer := 0;
        db_crc_dq1      : integer := 0;
        db_crc_dq2      : integer := 0;
        db_crc_dq3      : integer := 0;
        db_crc_dq4      : integer := 0;
        db_crc_dq5      : integer := 0;
        db_crc_dq6      : integer := 0;
        db_crc_dq7      : integer := 0;
        db_crc_dq8      : integer := 0;
        db_crc_x4_or_x8_or_x9: string  := "x8_mode";
        db_crc_en       : string  := "crc_disable";
        db_rwlat_mode   : string  := "csr_vlu";
        db_afi_wlat_vlu : integer := 0;
        db_afi_rlat_vlu : integer := 0;
        db_ptr_pipeline_depth: integer := 0;
        db_preamble_mode: string  := "preamble_one_cycle";
        db_reset_auto_release: string  := "auto_release";
        db_data_alignment_mode: string  := "align_disable";
        db_db2core_registered: string  := "false";
        db_core_or_hmc2db_registered: string  := "false";
        dbc_core_clk_sel: integer := 0;
        db_seq_rd_en_full_pipeline: integer := 0;
        dbc_wb_reserved_entry: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        db_pin_0_ac_hmc_data_override_ena: string  := "false";
        db_pin_0_in_bypass: string  := "true";
        db_pin_0_mode   : string  := "dq_mode";
        db_pin_0_oe_bypass: string  := "true";
        db_pin_0_oe_invert: string  := "false";
        db_pin_0_out_bypass: string  := "true";
        db_pin_0_wr_invert: string  := "false";
        db_pin_1_ac_hmc_data_override_ena: string  := "false";
        db_pin_1_in_bypass: string  := "true";
        db_pin_1_mode   : string  := "dq_mode";
        db_pin_1_oe_bypass: string  := "true";
        db_pin_1_oe_invert: string  := "false";
        db_pin_1_out_bypass: string  := "true";
        db_pin_1_wr_invert: string  := "false";
        db_pin_2_ac_hmc_data_override_ena: string  := "false";
        db_pin_2_in_bypass: string  := "true";
        db_pin_2_mode   : string  := "dq_mode";
        db_pin_2_oe_bypass: string  := "true";
        db_pin_2_oe_invert: string  := "false";
        db_pin_2_out_bypass: string  := "true";
        db_pin_2_wr_invert: string  := "false";
        db_pin_3_ac_hmc_data_override_ena: string  := "false";
        db_pin_3_in_bypass: string  := "true";
        db_pin_3_mode   : string  := "dq_mode";
        db_pin_3_oe_bypass: string  := "true";
        db_pin_3_oe_invert: string  := "false";
        db_pin_3_out_bypass: string  := "true";
        db_pin_3_wr_invert: string  := "false";
        db_pin_4_ac_hmc_data_override_ena: string  := "false";
        db_pin_4_in_bypass: string  := "true";
        db_pin_4_mode   : string  := "dq_mode";
        db_pin_4_oe_bypass: string  := "true";
        db_pin_4_oe_invert: string  := "false";
        db_pin_4_out_bypass: string  := "true";
        db_pin_4_wr_invert: string  := "false";
        db_pin_5_ac_hmc_data_override_ena: string  := "false";
        db_pin_5_in_bypass: string  := "true";
        db_pin_5_mode   : string  := "dq_mode";
        db_pin_5_oe_bypass: string  := "true";
        db_pin_5_oe_invert: string  := "false";
        db_pin_5_out_bypass: string  := "true";
        db_pin_5_wr_invert: string  := "false";
        db_pin_6_ac_hmc_data_override_ena: string  := "false";
        db_pin_6_in_bypass: string  := "true";
        db_pin_6_mode   : string  := "dq_mode";
        db_pin_6_oe_bypass: string  := "true";
        db_pin_6_oe_invert: string  := "false";
        db_pin_6_out_bypass: string  := "true";
        db_pin_6_wr_invert: string  := "false";
        db_pin_7_ac_hmc_data_override_ena: string  := "false";
        db_pin_7_in_bypass: string  := "true";
        db_pin_7_mode   : string  := "dq_mode";
        db_pin_7_oe_bypass: string  := "true";
        db_pin_7_oe_invert: string  := "false";
        db_pin_7_out_bypass: string  := "true";
        db_pin_7_wr_invert: string  := "false";
        db_pin_8_ac_hmc_data_override_ena: string  := "false";
        db_pin_8_in_bypass: string  := "true";
        db_pin_8_mode   : string  := "dq_mode";
        db_pin_8_oe_bypass: string  := "true";
        db_pin_8_oe_invert: string  := "false";
        db_pin_8_out_bypass: string  := "true";
        db_pin_8_wr_invert: string  := "false";
        db_pin_9_ac_hmc_data_override_ena: string  := "false";
        db_pin_9_in_bypass: string  := "true";
        db_pin_9_mode   : string  := "dq_mode";
        db_pin_9_oe_bypass: string  := "true";
        db_pin_9_oe_invert: string  := "false";
        db_pin_9_out_bypass: string  := "true";
        db_pin_9_wr_invert: string  := "false";
        db_pin_10_ac_hmc_data_override_ena: string  := "false";
        db_pin_10_in_bypass: string  := "true";
        db_pin_10_mode  : string  := "dq_mode";
        db_pin_10_oe_bypass: string  := "true";
        db_pin_10_oe_invert: string  := "false";
        db_pin_10_out_bypass: string  := "true";
        db_pin_10_wr_invert: string  := "false";
        db_pin_11_ac_hmc_data_override_ena: string  := "false";
        db_pin_11_in_bypass: string  := "true";
        db_pin_11_mode  : string  := "dq_mode";
        db_pin_11_oe_bypass: string  := "true";
        db_pin_11_oe_invert: string  := "false";
        db_pin_11_out_bypass: string  := "true";
        db_pin_11_wr_invert: string  := "false";
        dll_rst_en      : string  := "dll_rst_dis";
        dll_en          : string  := "dll_dis";
        dll_core_updnen : string  := "core_updn_dis";
        dll_ctlsel      : string  := "ctl_dynamic";
        dll_ctl_static  : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dqs_lgc_swap_dqs_a_b: string  := "false";
        dqs_lgc_dqs_a_interp_en: string  := "false";
        dqs_lgc_dqs_b_interp_en: string  := "false";
        dqs_lgc_pvt_input_delay_a: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dqs_lgc_pvt_input_delay_b: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dqs_lgc_enable_toggler: string  := "preamble_track_dqs_enable";
        dqs_lgc_phase_shift_b: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dqs_lgc_phase_shift_a: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dqs_lgc_pack_mode: string  := "packed";
        dqs_lgc_pst_preamble_mode: string  := "ddr3_preamble";
        dqs_lgc_pst_en_shrink: string  := "shrink_1_0";
        dqs_lgc_broadcast_enable: string  := "disable_broadcast";
        dqs_lgc_burst_length: string  := "burst_length_2";
        dqs_lgc_ddr4_search: string  := "ddr3_search";
        dqs_lgc_count_threshold: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oct_size        : integer := 1;
        hps_ctrl_en     : string  := "false";
        silicon_rev     : string  := "20nm5es";
        pingpong_primary: string  := "false";
        pingpong_secondary: string  := "false";
        pin_0_dqs_x4_mode: vl_notype;
        pin_1_dqs_x4_mode: vl_notype;
        pin_2_dqs_x4_mode: vl_notype;
        pin_3_dqs_x4_mode: vl_notype;
        pin_4_dqs_x4_mode: vl_notype;
        pin_5_dqs_x4_mode: vl_notype;
        pin_6_dqs_x4_mode: vl_notype;
        pin_7_dqs_x4_mode: vl_notype;
        pin_8_dqs_x4_mode: vl_notype;
        pin_9_dqs_x4_mode: vl_notype;
        pin_10_dqs_x4_mode: vl_notype;
        pin_11_dqs_x4_mode: vl_notype;
        pin_0_gpio_or_ddr: string  := "ddr";
        pin_1_gpio_or_ddr: string  := "ddr";
        pin_2_gpio_or_ddr: string  := "ddr";
        pin_3_gpio_or_ddr: string  := "ddr";
        pin_4_gpio_or_ddr: string  := "ddr";
        pin_5_gpio_or_ddr: string  := "ddr";
        pin_6_gpio_or_ddr: string  := "ddr";
        pin_7_gpio_or_ddr: string  := "ddr";
        pin_8_gpio_or_ddr: string  := "ddr";
        pin_9_gpio_or_ddr: string  := "ddr";
        pin_10_gpio_or_ddr: string  := "ddr";
        pin_11_gpio_or_ddr: string  := "ddr";
        fast_interpolator_sim: integer := 0
    );
    port(
        phy_clk         : in     vl_logic_vector(1 downto 0);
        phy_clk_phs     : in     vl_logic_vector(7 downto 0);
        reset_n         : in     vl_logic;
        pll_locked      : in     vl_logic;
        dll_ref_clk     : in     vl_logic;
        ioereg_locked   : out    vl_logic_vector(5 downto 0);
        oe_from_core    : in     vl_logic_vector(47 downto 0);
        data_from_core  : in     vl_logic_vector(95 downto 0);
        data_to_core    : out    vl_logic_vector(95 downto 0);
        mrnk_read_core  : in     vl_logic_vector(15 downto 0);
        mrnk_write_core : in     vl_logic_vector(15 downto 0);
        rdata_en_full_core: in     vl_logic_vector(3 downto 0);
        rdata_valid_core: out    vl_logic_vector(3 downto 0);
        core2dbc_rd_data_rdy: in     vl_logic;
        core2dbc_wr_data_vld0: in     vl_logic;
        core2dbc_wr_data_vld1: in     vl_logic;
        core2dbc_wr_ecc_info: in     vl_logic_vector(12 downto 0);
        dbc2core_rd_data_vld0: out    vl_logic;
        dbc2core_rd_data_vld1: out    vl_logic;
        dbc2core_rd_type: out    vl_logic;
        dbc2core_wb_pointer: out    vl_logic_vector(11 downto 0);
        dbc2core_wr_data_rdy: out    vl_logic;
        ac_hmc          : in     vl_logic_vector(95 downto 0);
        afi_rlat_core   : out    vl_logic_vector(5 downto 0);
        afi_wlat_core   : out    vl_logic_vector(5 downto 0);
        cfg_dbc         : in     vl_logic_vector(16 downto 0);
        ctl2dbc0        : in     vl_logic_vector(50 downto 0);
        ctl2dbc1        : in     vl_logic_vector(50 downto 0);
        dbc2ctl         : out    vl_logic_vector(22 downto 0);
        cal_avl_in      : in     vl_logic_vector(54 downto 0);
        cal_avl_readdata_out: out    vl_logic_vector(31 downto 0);
        cal_avl_out     : out    vl_logic_vector(54 downto 0);
        cal_avl_readdata_in: in     vl_logic_vector(31 downto 0);
        dqs_in          : in     vl_logic_vector(1 downto 0);
        broadcast_in_bot: in     vl_logic;
        broadcast_in_top: in     vl_logic;
        broadcast_out_bot: out    vl_logic;
        broadcast_out_top: out    vl_logic;
        data_in         : in     vl_logic_vector(11 downto 0);
        data_out        : out    vl_logic_vector(11 downto 0);
        data_oe         : out    vl_logic_vector(11 downto 0);
        oct_enable      : out    vl_logic_vector(11 downto 0);
        core_dll        : in     vl_logic_vector(2 downto 0);
        dll_core        : out    vl_logic_vector(12 downto 0);
        sync_clk_bot_in : in     vl_logic;
        sync_clk_bot_out: out    vl_logic;
        sync_clk_top_in : in     vl_logic;
        sync_clk_top_out: out    vl_logic;
        sync_data_bot_in: in     vl_logic;
        sync_data_bot_out: out    vl_logic;
        sync_data_top_in: in     vl_logic;
        sync_data_top_out: out    vl_logic;
        dft_phy_clk     : out    vl_logic_vector(1 downto 0);
        test_clk        : in     vl_logic;
        dft_prbs_ena_n  : in     vl_logic;
        dft_prbs_done   : out    vl_logic;
        dft_prbs_pass   : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of phy_clk_phs_freq : constant is 1;
    attribute mti_svvh_generic_type of mode_rate_in : constant is 1;
    attribute mti_svvh_generic_type of mode_rate_out : constant is 1;
    attribute mti_svvh_generic_type of pipe_latency : constant is 2;
    attribute mti_svvh_generic_type of rd_valid_delay : constant is 2;
    attribute mti_svvh_generic_type of dqs_enable_delay : constant is 2;
    attribute mti_svvh_generic_type of phy_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_dqs_b_en : constant is 1;
    attribute mti_svvh_generic_type of pin_0_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_0_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_0_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_0_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_0_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_1_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_1_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_1_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_1_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_1_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_2_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_2_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_2_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_2_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_2_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_3_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_3_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_3_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_3_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_3_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_4_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_4_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_4_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_4_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_4_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_5_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_5_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_5_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_5_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_5_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_6_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_6_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_6_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_6_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_6_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_7_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_7_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_7_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_7_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_7_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_8_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_8_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_8_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_8_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_8_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_9_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_9_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_9_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_9_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_9_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_10_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_10_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_10_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_10_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_10_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_11_initial_out : constant is 1;
    attribute mti_svvh_generic_type of pin_11_mode_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_11_output_phase : constant is 2;
    attribute mti_svvh_generic_type of pin_11_oct_mode : constant is 1;
    attribute mti_svvh_generic_type of pin_11_data_in_mode : constant is 1;
    attribute mti_svvh_generic_type of avl_base_addr : constant is 2;
    attribute mti_svvh_generic_type of avl_ena : constant is 1;
    attribute mti_svvh_generic_type of db_hmc_or_core : constant is 1;
    attribute mti_svvh_generic_type of db_dbi_sel : constant is 1;
    attribute mti_svvh_generic_type of db_dbi_wr_en : constant is 1;
    attribute mti_svvh_generic_type of db_dbi_rd_en : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq0 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq1 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq2 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq3 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq4 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq5 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq6 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq7 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_dq8 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_x4_or_x8_or_x9 : constant is 1;
    attribute mti_svvh_generic_type of db_crc_en : constant is 1;
    attribute mti_svvh_generic_type of db_rwlat_mode : constant is 1;
    attribute mti_svvh_generic_type of db_afi_wlat_vlu : constant is 1;
    attribute mti_svvh_generic_type of db_afi_rlat_vlu : constant is 1;
    attribute mti_svvh_generic_type of db_ptr_pipeline_depth : constant is 1;
    attribute mti_svvh_generic_type of db_preamble_mode : constant is 1;
    attribute mti_svvh_generic_type of db_reset_auto_release : constant is 1;
    attribute mti_svvh_generic_type of db_data_alignment_mode : constant is 1;
    attribute mti_svvh_generic_type of db_db2core_registered : constant is 1;
    attribute mti_svvh_generic_type of db_core_or_hmc2db_registered : constant is 1;
    attribute mti_svvh_generic_type of dbc_core_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of db_seq_rd_en_full_pipeline : constant is 1;
    attribute mti_svvh_generic_type of dbc_wb_reserved_entry : constant is 2;
    attribute mti_svvh_generic_type of db_pin_0_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_0_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_0_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_0_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_0_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_0_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_0_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_1_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_1_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_1_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_1_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_1_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_1_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_1_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_2_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_2_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_2_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_2_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_2_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_2_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_2_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_3_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_3_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_3_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_3_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_3_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_3_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_3_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_4_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_4_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_4_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_4_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_4_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_4_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_4_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_5_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_5_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_5_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_5_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_5_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_5_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_5_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_6_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_6_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_6_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_6_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_6_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_6_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_6_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_7_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_7_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_7_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_7_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_7_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_7_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_7_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_8_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_8_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_8_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_8_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_8_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_8_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_8_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_9_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_9_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_9_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_9_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_9_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_9_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_9_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_10_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_10_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_10_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_10_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_10_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_10_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_10_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_11_ac_hmc_data_override_ena : constant is 1;
    attribute mti_svvh_generic_type of db_pin_11_in_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_11_mode : constant is 1;
    attribute mti_svvh_generic_type of db_pin_11_oe_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_11_oe_invert : constant is 1;
    attribute mti_svvh_generic_type of db_pin_11_out_bypass : constant is 1;
    attribute mti_svvh_generic_type of db_pin_11_wr_invert : constant is 1;
    attribute mti_svvh_generic_type of dll_rst_en : constant is 1;
    attribute mti_svvh_generic_type of dll_en : constant is 1;
    attribute mti_svvh_generic_type of dll_core_updnen : constant is 1;
    attribute mti_svvh_generic_type of dll_ctlsel : constant is 1;
    attribute mti_svvh_generic_type of dll_ctl_static : constant is 2;
    attribute mti_svvh_generic_type of dqs_lgc_swap_dqs_a_b : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_dqs_a_interp_en : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_dqs_b_interp_en : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_pvt_input_delay_a : constant is 2;
    attribute mti_svvh_generic_type of dqs_lgc_pvt_input_delay_b : constant is 2;
    attribute mti_svvh_generic_type of dqs_lgc_enable_toggler : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_phase_shift_b : constant is 2;
    attribute mti_svvh_generic_type of dqs_lgc_phase_shift_a : constant is 2;
    attribute mti_svvh_generic_type of dqs_lgc_pack_mode : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_pst_preamble_mode : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_pst_en_shrink : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_broadcast_enable : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_burst_length : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_ddr4_search : constant is 1;
    attribute mti_svvh_generic_type of dqs_lgc_count_threshold : constant is 2;
    attribute mti_svvh_generic_type of oct_size : constant is 1;
    attribute mti_svvh_generic_type of hps_ctrl_en : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of pingpong_primary : constant is 1;
    attribute mti_svvh_generic_type of pingpong_secondary : constant is 1;
    attribute mti_svvh_generic_type of pin_0_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_1_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_2_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_3_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_4_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_5_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_6_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_7_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_8_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_9_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_10_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_11_dqs_x4_mode : constant is 3;
    attribute mti_svvh_generic_type of pin_0_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_1_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_2_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_3_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_4_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_5_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_6_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_7_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_8_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_9_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_10_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of pin_11_gpio_or_ddr : constant is 1;
    attribute mti_svvh_generic_type of fast_interpolator_sim : constant is 1;
end twentynm_io_12_lane;
