`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21fc3gV01Fy0xvidTB5rQ3sOuY+EZZjnJX8ZQUdTyoWUw2L43kZmE6+VgH+0CpGD
EA70kTl5pZPFRlGGFP+EhXUoW29bWH9eeEHUb/hGsz/+HH/z9Rrvie6wHxRvkfrw
nkctB/3kIw769LdYe+/jax0Sxv7adPKR8hutheOVvJLTl3JjbkTzncg7Z9tWB82A
SL6xNz/18a5P/kc8LXHLl/Seyg9f6lq3vLGB2+siCckj8ceC50qW0PR8PB/1XkJi
IWD3/HBOFg9mcEDQBUDcYc3q6m/pq4YQP6bDKXojZj538jcy9Sm3CGKUX/KkNzQJ
lFewSULcaFPQk5ULjkLLZ7rF/Us4rS3oex0jFiZ7MA2gMzZCOQRcxrfc6m8mWbot
WmHhBOV6s2SjkClxxmpfJr/s0kjhBYPCe0+qfdXfrxYLzxKAT8pqqP7sWhN0lfmG
vnjeFjeyt7RNQI3iwL+MbvjQomF9i6OzzMfvW5FvMvP90Vuuk6B37ECvTvir9UFA
0Ldu9R/n7ykE5z7pYdhHKo7u2R3+3vTJNAogo5OC2P3WktrH3roP9hpGEgIdQ0CJ
CSGD6wSegXDPnTWQShhNmKBNZxf8ACpCdEVOqZa7fHhJMBwXcyt2tbiZn0ent5H+
AHpwmYjBA5xK6c0nc+uKmAYMX3BERsZorGK4BnMqkfvvyg0pIajSE1aD7gVztjva
EB+kQVoAciWtwpDtog49mO6JmPLBbCF3kuKe5HbolEcgVlin35bY9RnyMrLKgizD
/qoIZqn092vd23PbH9+hFujFlHENWizVXbMl1bNyIHH2EJ913gG7QIPw5QWykk1O
t/gQJ/kojqFFXvYSWb8Wb62w1+9qKLd8lh8blrs/q3zS4l+KfZRKXpKDaVM256Nc
6p3oOInuotSUxWRyRdA1YhWKEdp8iJ383XZjE1yHMcXg3TATyy2wVjIJAwlwdVrj
bOk1fIWaps4nwaofMx27gVrjildVBzQvCR+oJ4n8l2W4rFyKjIWgF6tUhKxvlJaE
ufGMRfVG3uKZmOleGF2fmNq79K9WCi1jg5u4XVN1+9/YMbkHyhoqUKVzegw4Zqec
X65BQlHdnF6c6Kgyv3SGYhhw/Eb+tBpyL045VP0fZj5veS7aOyXXWhXzpoRI4zbQ
+u3zeI6O2ND9pc9ZhqFWaCXMG5/8y+RLsGsMZJd6IJDl8aZGZ1r+WNiInBkBhRMz
gggVa9zvbdrxc+TvUjH7O75+qs7XHjAQex7E/AsaKkxFw7ZpbHHu2/32romJQtpR
J1PLm9TxgfN/R2OnkJyBuqmTdW/DzblaP3VYOAiUPu1wKK7vCLRKlCF63VzxCHkg
BVQBGqYDo8E58U0cA7higQ==
`protect END_PROTECTED
