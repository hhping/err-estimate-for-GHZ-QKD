`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRnhA+BRfGHKXeRul9OkqZRmMVAKvSz97JMWCUa8f4yKh+urykDXAx1cUyZInxuT
QJOnLJBu3h5DHAZoWJoFi+zJvB4iMM6WEin7KBy/qj76/E4OsDKPlOa8/S3INUbX
WET9WcWYw2awSC5GBCmEw8vaB9nslXJRPpa4RuT3exZMrawZVHTqWWnmPQCRTEki
GVPUmJc/N+iljYbCAgB7VrKWfqqcPDo35ibAOjKVMEwRsyE9OodFajVhKDorbw1k
9rNp4AoTGI6lhnhveLbYqhVdguslGYMYNIBF07Gy1IrGNc1SEkRyWkhREq8/eZXs
VEavBKEepJkXigyUzSPMwYQnaqWeWqVwDgZDqg8Es1/0UTuNL3brE/i+lKFUggTW
C9ePonESEPxjoEbsrSQgxbdVkVjkuB8fbL1FvNWy2oR5NguMgnNezLOS5/HbndiQ
h4MnyMSgL9+t3mq4zwQ01q4bJ7G8iYCGQF6HQEazp0+whH0CBeGLN+ESS8OmrQa/
pw7mZYonaxLrCSq52zREPftsxN5kAOmrtADdp+2BfyW1O7kkNnHIUB2+QiL4+EBM
bLQzNmgd/YmDT+n5WH+sWYODOqYjZStPcNxd7mf1Ug8a86o5DNScHxiGiNROC8WS
+3RN7hfKY+GoHMMwLPwTXMzylvCbchaV3dNzAgi5/ttt6wi0W1gVPQT8MXy4IO6a
8DPlvxOG+nCSV8ZZahjGrLex9SDIsofm86LatXM3j/iyXwArGkwjjJgoF2golpKQ
KdBX2ClJ4KSx3UoDEQ4uXboebsWS8y60K1++83P3O+Q0Bpi+hodIcWTtj/wENFAD
MXf8N2Dya58uUVohUMEFCdRjqaRvUkPyRy+0fEQyxfLuDNcuH0Km8dGEAkWjexgG
DWYRF8ZzQcrK9is71teZoYZLhe7oV4KkMmsHFDp5Z3T1C3hEuLQXKQKP+VR0Ry9t
6DvuOrvWbCbs/RjKjNDAV0nJD+fJPou1bHrRi3Z1BGNhABakrIq2fMD889oyGLHj
ovlMmsUIrZiiCQU8re219dbRH9CrZjd/EcO0LGVVlSgHfK/jClQgQAX6YQO1Bls1
ndhM5H4JDEr2b7kK8aA/DKzREt2xJNt98OknxXptR5WHibirJJrGfGaBhuKw4ccW
7wseySqEUOS2xw9SDSxdRdl5Ocj3s3A223aA/Vszfws=
`protect END_PROTECTED
