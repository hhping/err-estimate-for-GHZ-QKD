`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wA7355VxZ4wwMbvYCxMce3ZmLvOtMz+uJyKCehIrphm78oinwQeDcRAo1yNNuHQi
0AuNcbt6VjnK19UT+o6YEgrfR4vWEt/a8+Z753KnpKr7FYReDQ+EWzK/dIkec23m
iuzRh6hVoXUfOvO20qm617RITfbAyRL3tMV0HnbHF1p+Dkqv693hYjdI6Oo2+8UI
6z1nwpFVr0R2zixIvoNk6OVb5U/0xiGOeZjLbOVOa0fCkbsX26LkYcVg8MFMyszt
OGxoPV+s0ZxoWIw9Vzn4KKQWjqMjfaQjvfulyPX1cCY0eClurDYn6Ubl1SvLCBrv
PLGesqNflSCiz4idml38SKtCfODIbRCg1/OUU6rQ4ho=
`protect END_PROTECTED
