`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asy5B9Us9OBervhBl3WaRL+FrtiQ691c+rxWxFKLHJW4KW7LbGYnkdenZLXssJvM
rdGpCBzC0qWBU5E8xNTT/O2uJj94drXeXmK6rt603EqwqlvzIDghNUaocq30RF0r
NtKxK76NNhPSlexnNQ6IeahlKeAvdgR1wdDl2TcWWGRjA1LUC9fEA+A/fX+5Vljn
1EeUW2O4ZogW0WQi4bfyK7zsYvhcDrWzQPCvDwB4IGpJ6nbSxDaDJDn0ePk0KpRV
OCcSGdns/k9RY16pHmUTv6FTCugdjusESio/3BmGovK6HEdr7ZWEAlgXcyyrDBzK
gLYJ+FNHxPj2b/G5lcWTZy54FHO0/8sS2nDTxzXyBWjMi7CZl+Rq/oLZpBEKym5M
XHxvT89z3vpYdnMW/aKhBR1156hKR+R3b4bTI7fFPOG1lwtATHFPdWlhhE9HN7oU
RVT+xwIl28wRgwFbFX1YVvDOE3pWVoAeDuYpXHHIEO4/bgyq5RDhnPfmRjAfcnwT
6lIFa6PdnMjlP0Uskxi3D9tUgFxtHoVC5D/J1zVkNNhoGMqgx2fFx3lP78tRu5g/
dB3lthRO9soSKe0l3qxjWTckIForlv/+jAQuUEAGX7FzK5u8lqf9ZAznIhYqJfXm
ZRpba2enD7uOa+arlykS6qKsBO9gpRIwYQHlcEdBOu6uVGOse/YNll3NMGM5QHSe
+nyClwVz58KNNSZscYSq2Rz5tk+dO/odf0RYDBH2fh9GFOJlob+tsO0F7MwP1OY3
sStokmCsGn6YOG83cURAEiZh4MLqT/5NtCoJk21kz7egi7EYQQOeX/gP+ZYmImrJ
xgfIgjB8+ERHIHWyILtQ+4jelzr5nuOc7YwBFRD4U/CiTD187MKb7GqFh8bObdA3
UYE2OixnVsun01rIRHLIb2ZrIZH+pw3DxnYRdvMd9+QyBTm1IkSJ1knTqr8Sd7Qm
mUBsJdmoVaExAflHu3hMe2n1Vg283vvzpzNuU8EfDB8FpCjOgdum+vFl9f6UBPhM
rHnxNLGEPUZ1s1czcaNf6bpfyzUcCmHGPXohHSvIEXC6ydKga1p0TteA5hhJ+zs5
9OPzqZ1oWqIxCdcc8F3Y9o0EzhHvk0VdTBLUPCuBxl3L0fVYPbxE8vbf2d1psZjR
MaN5lkFrTUYYjpu4OY8D1ElYt5YEXZ7sh9evPePwes9Au9bC/hUJvg7OiWNqIPik
aXTUN55peJPgXmpzJE0HqM3U7WN0mxQ+6nxKrE2bSNapwSsijb0VtKo8M/6sFk6C
bedwNXraZGO0tLaEgh0dG6zIoL6bgFETLPXFhAPT2XuIcO1jIj95TGfJ9IUWVA3V
aeo9w9tHBsGvFjKtm2MhxytsDYQVGzYUDenZrrrhHQUyaafgNv5sS7aK/UzPW4TD
xuaaSzxE2EdBRbEnrrQokRV2RVkh22Bk3QyXZgIcHCXD2jEAmOOBNfhuGuq8U1lV
lRlE6vgCQEEwveRmBJt0x1qZpMgYuj+mHlwUzw/WUGtVl1R9l5Z2zmOtghzfDINO
P6tnlREtxLeNuFoZBpX58PPnkHDCAlYj09FjYn7BQ+wPM3sWuaLio3Gyk8g6/dLN
`protect END_PROTECTED
