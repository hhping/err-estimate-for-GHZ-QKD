`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RhO8/EiEFnVyw7F1nO8SNtTtjW9z4azbtqf1q1bnfoEYAw3gDIVm4T5hEGDY2QC
uE5NJQsROz85dKXLpqeIjN2Fa+dkkbuzeKggSvkyR+g9U3N2XF56Gd2Bj/GtrvwQ
4qU3kcRLboa9vyP09IeOJcMdBld+hLnyCQTRQ1Xz0YFHfBhkf0e/zNuP94LV4E8A
8Vyry/qXoiGfKjRtzo+glr7XxiGSujDKrVIPBgjqkIq4gShlUC1hbA9arjS+8QDt
bdeSfC6Wtg+Dnv9dzqYY+bFFdfow5cTBvSh1NOFIzr78ZNcdFeP3p9vMNdNDJQfZ
S5HHQ0PuFSRIW179I99CLg6QLfQPbWrPg82Cbw9aIIm77l6ct+V3BHKDLJ2TPCQl
fuS4C/exzYltpyEcufhhmk5DE7iC1YwA3Kb7naKg0bQ1BSECj1rjtJosAG99MNsj
pxlaRyzJrTJ6niJdSMFQCWAlsH0V6GgoUB3OAJ7++Q6hSaWZS3XnqjwzU0T/0SiX
AU/GWbnNgyMshp0o1fEOuc7K+M1mKXqAH3cy/zwAIDnTo1fcvZavlrlt2gi84xSg
qri9UsYWsNQMgpP55alx6UUyjBoL9kPHltRicX7WjtK4JrshIKLiNkWuMs55az1M
mWnRyP66AyH2qX+naciVjYj7rTl4kaGw8AM0ueiW5apT6APP5TfxiaWz97Orid9B
ubtST/t5ZktKSytFL0xlu6jS1JmLCIiiTafyRmdeaGamhpa6o8yQXckV9bLK3032
+SIawrq2VsvhLBFrV1TzjY2SUNjncit7bLhSQLkLb1cHsAOxgc4MVcSWJb+kS8fM
hK+b67bGd21tFOSxgmjZ400/rFZ+yzcq91cL+L51z6ZqFOeLqOjfVl5DWcgpep9c
HJnGAqhFzp18ctGbFqxT9mXkjuTnSFVW7KU6naLxv+e/gMUYVMv7AxT/1Fz86M6J
WsKJxuPNghc4zoG0pT/zFHOdbjyv5VX5YRxc8EzjoKD6JU50yuYoULtgmN+SdhOU
Io0vj06tOZpN6Enu+dRnSXwQkCS44TkY4Dtd1t7sybcdUTyec5laoJr8b7GOi183
uF9xXRM7dIpnbgtizLQ+JJanEmIw+TDnb1HvDu/XM3rXagB1wqwEdRbR6HQG71T0
6JAIRLOdeobnXuDzIz+QgkmCABzxtBSeJFcAq6bP0iaPYtLHqlA8Guft0WdGxTF+
vqVnUdA3bfxunv0jO0jQjfLgg30fYUJjjODcXZlNaG01Y3h2Fh0CohaRUyTIIWhn
KnHSqs5eCHvY3L8SDniBx8a/zmZzEi3y7tIBdN78kahZ7B31urMX+/CuJ18ngYvA
XQ1iTkzhu2uvwkorDN2kw63+3US/Z5fBRoj7w9vSTIeJHnwAcU1LKBlFwdL+C22i
AE8SyTpSm3IXdKMCLlC/OiM8b4azHxdCYXii/8n5wEPrTLmR6vCC8iC5wrCQGF0f
inv0SghwiI8m03+aSBYXGupeYlj1lYNqI1FE/L6fmepqNaFxFGvfDbW1wkX6vBIL
FbGGIooMs33tr8pO1JwUnOyQEeqjqiHXwLDiRfG5fz7bBR/ID6ISLzhvjfQZ1fL1
xJhmzBh4yCa4M69o+cb2OVkSZX808fgdvrbTsuVLDPqkeQFom0WywrRhouC0g90N
aB10Svlh8KJPS7Nhy6bjoZTXrbA4cmJgU+FVIY7C6Pj6F5uNTlCoMNJC6+0Rccdp
YmCQC2qcvmwIZamMtpdXBkm2LabA5/ojZAFCMxlek/QhK+3p7dfXUVu8EXyxryRM
Y+1qUoVPUDdt1+aR3GHkkBqX71CRgE4T5cPkH18dQQYk1ykR/UMW5FmzGiQCEPQ4
aVUNd0un7EBRvjbRPTNQxoA36EVgx4vMll08BUdUyVCfNm6f3Daa6heDDSRqGg46
2gUn/sm4ArhnJDr+LaA1OuintVzckRRtqvskjogmZo10tLPR2nWTj7FH2HZUkXUR
ckoFWcVHzGIFjGJKk91NvzQ3AV+YcXJ8Wb2KD9t7zbuX8GFvJ7LhE5Q+QFZ3nQG/
tLKlHN7TQlSfUwvTPJzEink80cNPyZvDl7cSWq+Ce47mI90qrEJo7q0i3aCQJKsT
eNQ7QeaY8nw2k8YobyX+Y8qDDorP/ekXAPq2GAEA4WwZBH/hPwmvBPE8SThcw72+
zmw4UDvS7g/Cnh7YUGsXGK+Bpzr+2/oJiJ96GzY2LXvkwmOm2+n/3fsItszraaX8
N2YiQ/o752GnBFZBZLZTgOkzOTzBtp2XjvbIm6s0LUq6sW3HLV2S91njICptpSA2
IREkbYECwIIWLLGqTWozWRwYVupicGb1/sN5AHIhSn7YSYTrcY3pDL0YRTYm0Pho
nBAKLargNanzyc2NXfJZkfMmBAZ9+tsC5xZS0TVY6jeICumzjLUMC86Hx4GQSNoW
Tq2yRDbh0s8Cdz3lXD6HjBSkUmOx+CUUDySGR7iJISP/lonpEUBqXu/Afz2GKXWa
WgdlheEdJXy4GmL1n4KG/KmpIFA5Z6e3noyGaU16nDoS77ZQDchHMRTE7Q+wjTT1
t/HUmRSn6ZInLScuO65pIjuh+BJbmou3ry6GuAdfmaIQDOmv86VyoywtKLZzOUwU
JAUYCQY4vO7C6ipQaFLagkayFmnqbipM9QcwQixigcLDFBvMwEj00gJcxGnGkNfp
NsakUOVPIH2FPjSowbSebA==
`protect END_PROTECTED
