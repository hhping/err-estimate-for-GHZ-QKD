`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qe7f1PiRUuLEaP4OI5DMNhwJ6XSWuaL8RpHAtEI3EGAeDWU9cSKDKDubFsspNS/i
Ipwcmz4xocCWHHShlzxz3Kuhuwsi28L1DCQRLqO4zUJqm6uhBTMZyk+vHmN0SqpD
5z6D97LUDuNoIlajSa9o98/e1k8gTPpnCHSoiE2zjkdp3yalCM8EnuUaC3Mz68nV
njOpmA76iqbqto5O3BP2B7ahBRROJ4sBMK22AvISr4XHoLLN86y11vzeAqa0PvFU
nCD369J89G7mJM6lyOs4eOiLvxTrkjBH+U4nRN/cx6md5nTiMi2J+c3Uborr/fLH
DMor3ReDuRd10Yl9oRVeQwZbNzX6YLIVhbSQNuXmfs7TTOxaVAP0+TrJSQFL5cw7
QbIKpubC1p4XC9kmjKwcU/ababAI/qGp97rsECQXwyzYxAeomyl/aFOsaWP9EGqa
RcqZPaZMtCyUj/+3zd2UIv0jEersbqkxbdTA4Zs/Zy34l87u0tNhIWaz5nRptoQp
zK3BZg8ezzZirNAuoPCwAZagL/Biw+Iy39Rq7VC8UTMbffSwHeeDuJaw7nuifDLz
8vri85YaZPixhj19qotHsUP0Lsvsy+Y5jHSw7vM8pdS1cM3sH+oibTXs1FoLAF/a
cEdKv80XAAqQvjXpxKT2QlMGeRwHrxzOjcF4UsZ8JHAfH86j9DlVlTKL+U93Rd2w
RXFyVsSCjJ+eszURgQo5Q1ahpHhn+FwZ2u9x0NtPGIwGzK0toYok5qq6qz4hHluH
vY/FUalJyGbzUSw8/zBLPSmLwIP+XAecxF7ZYvyk1/a3EXBnrrOniclEfnuZXhHu
URx5l1mGi998pFIqE4SEk904OFHiLQJtMXg8xd+eWcPeqm7gLhsknHz7s0rR4BPw
z3mmyuPeBw3Q4t2Z7lP059/QFquOWKpUOP03j0iWgKZsKneZxkIeLWr7mf+LX3xD
/EYRUnoP++g1yvXtKCqE8rXPaAm5OGenoKOm3dJvRAp/1SMe+FWNggvEWOmck+Z3
815lpBBJF7oAkO/w7AvnDfg8Oq4EFoOR4glv2/ghZkVXAQcoJQLSqSCAzoAVc4Zp
wQfwIXaydj7LFwi+ZPPHk9MQrN5SxBXkc75y5aH8JlEhaUrT1bAm7nARWiKOMGWk
HRg67CeWOx2CEesAgCdlkhdghVWgq0BO+lMw8Y9D7eyoMuQeu8cDU4NIER592f9t
swnJKQ6/ygzK/nZPCD27q+4Xse3AXUGUl1wPqbgWyXHDPJE1GrBDoY/qVVsunZKh
oREx/+aOoxuW06eNX+wMxw==
`protect END_PROTECTED
