`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8qQTLypQ8qGYEx2bI1S6Fy61ypvOPbmWbjgvA9fbT6sHsvsBCA0J0Z7n9+BXqKp8
Aov6W4CurxSUDMVWQL7eMdAvT9g7GVuY27adBVyq8VE5fdS1yrQxdaAu3sXNES01
W0zKXDr+QLDrOZcjR/BtV2VbXDzYT2GU7/HtnrSBVG58sKUv2+XeyE6cNMtRlQXo
E+tyZ0kH+rAxayEoBSUXXhdsT9/u5v0quCmj+E2vK0qwpuS4kHu5jzvtyuQ66KdB
BBnaLnM4UP2Ceec7Fr+6Ktb2t6j57c/h8AjGmo+h8haZKzLBX0koc8cqHZk+eZUJ
lMDCrjEB6lwTxWR37E7LzUz0tvgiCAJgeh50Q4U88emhYT/6norvRF+KHTl/hMwC
I1dHe5c7YnG8KXagJuTv8o8Bx9IYV9MidnG28V1e29Iu0A8O1e+HaIY2MpX0Cu73
q5rD/vhpqnED4chGmELqL4y0nu2Ipp/MWI+aZSZjrpKii83pAU9xD2wcdo2QyxWu
wHxWbKQl/GwKMwsKDY8YhJi5TB5kB7lCKCQE8FtD52IZ94/9uvlywlMtmhVtfP/X
mA4rgHwHma6FtqnP3cCIrcC8/leR6eZ203RzD04oo7Du+0ibjI2gPVFgIwyVjWnp
HkhH8ROTZgXWpYgdYlB8vEHEzuGK9rp06Xyu2+rBw+YtCe1do+sZ4wdum9iCpu/K
QkSwmi6CIahK/EY91coiATx3nVfcWtD2d2OYTAS0BWdgY7036ehPKITw4B1lKmrv
XpwLDqLE4/LlKe9lpCAHsWlOifVaxXUOIh7RCKOzK9ov+ZZFAXufIsgTYTmz2raC
sQSbQfOWx5nA6RO0+KkjqvM3Nv70ChH/sF/bQc9r0DpY1V3/CU8TZhOZhDwTLWBV
q96sPdNIFL9hd3/C973ducTDDA8J31d35h835FkJXfwB/oZuYIdcU7vIYreCGLN+
dlwVC5vwdlLgg7CxQ/yjJIzVSGVPENWjtY7n849yjcIFyEDYkFhygsM21nVgBAwU
r6Rsut7eq6UFlhHQ6eiy6xrPy23Iw27w6DYRoT14XBis5KJwB4taa2PnfjFWkgMn
zS7p9DFufzX/zfYACaUMAQ==
`protect END_PROTECTED
