`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P8aiAX38z3oW5biF9KNnlJIM5dhp8dbfb5pWpgKYWPxoUjjNThe2+WUuFyrSq1ge
qrUOHpCw76GzQkyiVjHhENQQIVpk/loD8QJKyHs0DW1reP2v8kk9ywxDaQ1Q2/Zx
iKOCea4ryVDckunFc80BjXI+g+BhUy0Wp430pSZ/ZTKKGvRm1LkAovQ0EPsQDp/A
SmHsnDUBqm6pS0wwmZuBApVNSr8cy8QVhjm3vtm6XJuACACWN87lIZnMBmJfzo5/
p6vD2Rt7y3/vRLMfzLa0KYpi+DDSPHcPlGE4wYs3KN3ENIDLGTGjTLW9JoxJ9Mbg
zFf561yK7ckUxZ/hUwiI44Sa9gQddNiWshreFoY5oBMOwP4C1zI938avDCbdEZoX
aPPIIfta4A3uI/RFNsH0yhn0WuxHeX3zwXjJ0rTInf69iQxaUhEZiZkA41trB6fA
YtBiyWfo20rtL0crKYFHGSOroLcEKtORJXzAUZteTMhsBiePtySLuJtsyL41MjMG
c2wKR3Nz2ypXsVaH9fLBcX2Cbp6nMSUkUdhDFnWJsNCdMoMg7V7zf5ueC5S9LkZh
ISrNFWCVbqUkSVgbyr9C9qByGFljS1RlXRJJixSZBpwK7pUR3L5rjT4/d5OQSi86
OktEocffVx6+LVIRXLJrsE/rFUwPxY/fTMduB7Z9nfE5cHU5ikFMrS1A36nxZ/dC
QWg4DsnrZnif8MCL8DTWFX2dlfBMry0atCmy7Ev1dMEzTM5D0hK+ZToTu+HMU1SG
0qnxQgbK1MEJWxZyFsnY4azPE+hIC5tc9E9Qez1FfE5QPKLnd5Za9SrBDqlHNOMW
iyVqanqtRMMNZfoiGuX035rCT2kec0Vc3eQm1tG4odX8JYXU6yk6pbRB7Mp0UCjO
UrSkuOl1GwZyKR5stsnJYqQMF8XkXBwLV1c1UAtbs6A9x4WH70nRHAl+stWRsyGr
xjsrw2ZbAtN8MyCxClWeZfhbOnSY/t5wZFdCc12eIxWfmtn30tq0l9uPkyYJiijx
eTWBT94kFSYSbaCb353DUtnt+gKOz/ume4DhPZx0gOG+E6cfvKUq9Pory/QEziw8
1Ohf2Jb8+rB3mh799xDJrDr4V6GKf976WM4oS8IFlM7T5I8NTtGZ6tDb8LPHmwaE
4TjGh2MCcdny62HYL++VirQNWeaanWXgfsq2161m9PSeB+I9nNTRXOIDqnq49JDy
F0cGnpGPt4OaKXj/Kh6+Hzj3QQz1zv/xNPZ1DU5xpr1O6T/V3gDnhs3++jzaqrYD
GQn0WAR3XgFBf4kj4OR+UQncsAhe7ZCU+mv/hXwo4xylfRFVo1RCXjvlImNaLlUU
Ub7vCqVIEGRPHtblZLq/kUW+eFFW9bAwVh4q/SEbhIFkjNNBwsmO0YCwWME5OaA9
h43SRfGqkYmEO3hEpwpkzwdkL7SHJlWz1UfxSv1SfKumHR/shy+e31euIChx+6um
CPsqzGX4qYFIeHay8xq6JuNooDb2PXusxf/C86K93ZZ8wrIS/A7/jhpYcHtrbZdM
FargevqLO80rNR5PgzOMT6jqv2Nk43LV/oyO5c1PlNE=
`protect END_PROTECTED
