`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOsSAW/JXbxU0G1IYLr00gPgfFXp5kpYFygWpX/XWjhmYpxFp0zLEg8tdBF4JF5U
B3mCs/Hxeo7XYECcFKCaCc6f63RGyU1heiAsUMpsxAgf+LgnQ5KCLzVyuFRfjUYL
572Ed7fbuoawOcrpfYSemeKLie/x+2i2oQX9JJCALGpfA+gWeP4vD0s9MoL8K0rG
Wo+fpz37Ckz1xK6yUgmuAoSgnaXM3CWgTHDnkom8pM7J45kP6sbBedrS4oRDlgOU
Iz4I3FUS14QeH8pGkH4j08AvmxlrGIuw5Wh8V76yekt9PU6poOopYilWKu+zcl1C
GEFe+k8REtc9U/mVK/aImPuVx2K9EwCkQpJ3nVRK+KlShn85krLdUaODC3nbyOyS
HTEC4/MFQT4lPBw3eJIZ7tKTW9b15f3j6Zb6GmGqdsq0AotnOttCebVQZasjM9FG
TNBpUqagKkHqjwofpfqnardf/FFFkBb2P7YRZGtGmMj3Qka6ZnSuTe3lZdPYuhfx
JM3M02aLfwNaILwOx5wEc2VQFkcc/i85r1csxqr0m29E+T2qiEaSkoW27CgoqQoq
Rdq/cyrFjk7yhFrDOO1MRZxkiPeEFQBM+yp7gKoPZoGM1PzBo4/t5f6XdOO6xmUy
bDeK5w3YTmRycTnuQWgYqQ==
`protect END_PROTECTED
