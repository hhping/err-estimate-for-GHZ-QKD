`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Td4V8RpaYAlDwceAE7prwn9UoIuEEMmcWNhib8i/uTba7Ajk1ja0YnIGSjjb7x4E
4Bxtba0koPhoisskuWQP+6vu8jb1U75GB+ZkpNnWo1Y06CD/+tBQuKBgTcB6EZxm
5jKbHTU3Jz2EMbWDkGxl1QHxsvJ5bs0jbIsn7g3+r/+LeOcVseqxHmG03I+XW71t
VBSQtOYBeKW22IgAb9tsHMwbdmqzu2BtL+hL1+omXnJOQaCroL7lihe6vvxas2l1
rGM5j1Km72b7Sg4LT5+HDvgAQRyJz0YD8VQ//CtEmLHFC9HmLugXY2mYChNQ6jzo
6VjX24oMwVYjBkXpSoNT82VFEy6pAXA9YXUyzfqrQTcL6OWCxvRSAh6+cnbMiisa
1GpDi9/yu2aBt3gKsOirqQxStV9EK//Sb3eAxGV7Irv67X85k2Z9qokDDRplAhN8
HEG3ROnvf0nPRDrZaUW8tZnyTM1ABhjp+O8SgIvMX/fFvfU8XRgWAeCNm4sd2Q6U
FWl/gq2fK7escA87XaFW9/AcR73z86iOCLpvok1P1p3HQODeOyPQH+wXlwx2GJIL
gksm/AHxp7Ega439UUz8lJFK+k6THOrZT7DmRjYwBiGNfX9INDbPCnAUGYaUGLVJ
AH2sM0i5HOA6rZtgk/YBoWEBU+fa2aoUkpfFBvQbDtcRA/z+g8nXgMwm2t6q2Ark
MRr0kY4JUOemjvywTdBodRdJ8iQ6lE5mcVDbvMWXPqhllr1eJrR0TZc33o6DWXzN
4690NTPEMOxCTort13rVE6pTZPSeX4Tw09LhGgIMNTH32gpnYsE+d0K0K3GzxVSw
KEJcv4r3cnjXl6QKtBoVbV9lUuiPEcfJXEi3ZAdUwaRKZin8ARRSAe16kw7IeGAy
SZxI6d+gEdMbaovSckznzLdy56/BWFdLLLTys07w8rD0CEKAgUbGgUaNiBFKj3qu
/HDXZUMR2re9ebvOBJ7zuhS+FM2B/zvC49zgCGQKSIIBSddDEbb1mNuHhwTFtOZY
if32oixAQRXsqlZVjEurJVR20S549oG22hCoAN5xA759ORpwpZ+jMGT2TJLoIwWM
SM/rKjTPVtDyu0l1+YVz5b15L0zeAMZASzIVKng97odb+hMF14OcK00PfOK3I0eQ
0Y7MyDNLLP7QxHbskRQa3WQvpZ60gXO0aO0IGuQo1ICZ242pKSyOUfWsVssMAk+k
YvAKSWp21S1updM/Q9WzQhLSkdHFBnzMt5kBICFg7ip2iomKWInoJsuKd34oJsib
q3r+h1RzmZ6QRJuEIFsw6bOaog0bcKct7Dw1/gaCAteNBD2YeX1lRATYk4Z/jghN
+qibxd04C2TJMTJxvdYAunW7dDZ2F1e8uO2Fg0Pzg8+GZrJ663Yow+0MRWfLG1Hk
VgY3CZLkp03kZn7LmKsMykttHogY/GFzjmkOGBwRPyXDAnmxFMIRPLMYesB/njhg
6vH0lrYs00G+KqtNk1BPMsJINZoCAN5X7+a6V9Mwmi6YIm9lCilhqv0IV6GOWz6M
lAhS2whiWpXblCX2ypNOomNIBnKcuLRzX8aDZBXaKGW7YsHaekzoEZF9SL+JUHsm
cVy0MNP2paFqD+2WFNJ5OeGQ0jxFHoYSa7y5qlD/nlyK7IELv7hbB/B/4OtSHaJi
mB30wyBNbdR3HQUHnGWt/x2SqnAuQH3qMsU4Laal3uS//IOX6yb24rJS9N729pYA
TO8HAdsTadcS/e9U7wnyDYmrJQMldtThkaC7rC+yafai7fby0Lu8pPai5k1eqtta
XmsnbePPrIytDb8kXKX1+JDsanCqY/Wk9k7Rd60BC2K1khAZl8W3mmMw15T2lojE
lXAcUzNA6HgFsUX+5TjvrV70vTDeaKTxEWb7Z5pvg89xMHmyn8TM6ApiL2eODNWU
oTAfLyYiPfnIFisAO7keKOuHc9dJkIKZAgIl7F2eYdC3a8rMupsHUGXN+j2PW1Zh
nvf/8TiabBlUfmP6CoL+kcvi8lnCeTTllJ8LVSTUvbZlC/xVXTnXvvRrdZySORdP
LVAhf9W3unuZwa8DPOa5DgI3AlIc7Kcm8yqjYU2VLe/XC3pnptzdONpFn9jMG6yQ
VwCj6RU+q2C5h4tmf0llFpLREePzOVi0AtxJKyp4HfzBOS+NNaXwexf8zBhyarcm
ld3Vq5htRKNc4+XgUqfidWbl+fyahjTUym4eOXI7dNBhjgspwjA2Uh4TkgcI3B3Q
y762+uSDaSrK/8SfID+wBhjpv+pgGl0AxN6/a8VoZxqtDredK0N3BwlJmDmTw9K/
rk706rSjLTphdvkiygIRG7sKYZrpHgNzb+02nF4fTrOXdRz7ZLUlgvSf6MS1Y+VM
EpPcJeIGhEVYrkgNuNu/OSIYjN/qO0uTYXFU/D67FXX05ZvtkBRHfwygr2VWXvM5
hPsy5RzwBmJMRhMWGqLCnANvV/VE4OOLlH7eJr5LcCxWhoFYzVvJ5GOTNruRkW98
4kvVqASWJt6+T3C22CzjFY8euOhZ4IY47PZNKizWAzzOIpQZSk0kEP0qONnkvip6
kR22TIIedQV0EeaMFe3mdqkDJy4OfjC/qd/61/510dvjyjIwhMbJ0uj2Gj+AlHOy
jh2iOljkxKzj86R5r/+OnZ5TRLuh4yd8mi2Lsp9LsAfzysNcnHPV6S3VTkDuT/Mc
A3gYZ2KoTSZB5TvA4z0pevHPqEmJsqFd+Mxi75KkkHuG1hTSwmdZKbibjkYS2FCo
CdJHN2fOCucz7KdcRkqWTimhnm+YiYNsEUVzphDIEBa2XUVuydjr3ZMLZ88WlIjU
KGi3d8//RAwPV8cOqFCwsgBtjoO8IpajvfYwMUapz/uVGvByY/RdftZ4F3ZtZGgM
wIp04HM8P+QndmA/79G3tE/qUs4N1HU0OSh7rHSfxKnsuEHRphRwYjSLy8hzpR9l
bfrNwVb8ELQXGlcQOEVI4z22GjAlOOS4JBaZzc3BSvMHEW6O5CEcDP+FGywA6ZHf
29OJbNlNaD7DzfUUClNCqcW2KdQIGaPWu2rDmsE963Jqp6I6/oZCtIqOSNjzGnyE
+Ah8s30b/zPnnbTfu5+jzrIPzQ/BHWGPf0pXMIUNEWieT4nhr8CcrdT2VA2ff7GX
ruzvzSddqU8t6mRKY2SCb/4O0W54NAay9Amw6DUGdI6JrNzBX6x9vg1dH0UHlsAH
VSlvKLuq1R/BGX9Wuad3gxZoj+VJ7dcqrha7jgIJ+KlxMaJv8TpelxVNFgP+CcYp
sKqkD7bY4rHHg2Eum8uG3FZdxLZLeNcCqgk5kuBy3Q+8jv2v0oGQqZQbCECHG8Mh
bpbB2ij/H618dp9hLpAG5oNz9Y3waiHJNfNtJsiNy2SO2SxTj3OZjgQJzBAjy+Od
iGi+kqFcfzxFNTVzOffJUGTRSCFEr7Q7+fHUDvg3Rua03gLVuP1gmV/g6sS+D2WY
r2bCGv/LV7XohAn3IawCbBK8III8dqFl+jeIyg4noTkZ6cMoP2vT+VuYmXMsffCM
vfjuykz/INqd3dvbFnDu1wsOzGhBnuONRnInQqKGzgH38RhPkfsD+ic1ijKRK8l6
p62VrNYj3xW/vvnmM9VDWlM4GdyUgLSLUgUcrIqTassZKBkPKLogoyRfizopYv6e
QkVKFasJyIOeohoQ4aZaFnpJ7pdqEirzkMUHkCPVn7TYVwE1+5eahwByC0tjD+p7
ZybOJSfBmhsy9RlZx9xy0O9rmPcXYWUYG5jVVzBVeZeRotb1/zhFexEvvtSr7SFp
oi/NlN2wsXdB3isbXbrTc7gn8EA0TuOQkn4aw5erfQF+E0NkZDs+e5vc3N/kiKnB
T6Xa9i/C2gi6v05rBlktdrC7S1mNwcNlJmmd++GpFg3oFEBwXtEXz51y2dE9BM+U
fsLX1eAe7xNmL0atDN6oeAFzlY9Vu5X3O7oVTWcP4vcdtAIy63EF/zGiJpPcdchd
4Od3DhU0LlmMQ3yJCx41xcXlvv/WAsZ8BaKQtSxf8opIAiX6LD73HVAnwBm5YTad
bMdi1TUxqdPcp/b7DLuDfRQYrLIfC7jpfECjbQf676aRHpP7m7b4w6g5i9ZvZSSC
SaUuHa+qML4+sF+SEVe1okzFqvF+hlqr89S6e4XJuWOt4o7vQ2isBLlzdiTQD0kq
pi26pEPbRuedqh5BI4C0Qj1pXkOmReWVDumciOp+EcAzC549yQwBmpIArHgjjXHd
DEiNzTQEXgRpL7IRG3cF2nwu5uYO0WP1Zk11ccrHvjHDRhGdBWJKocMBMxzrklXZ
EInFtUMFWTrPvJfK5g9KVP4Pz+lNWyEh6ukd7AR2Cwy6dTYL6UlF4Ix5zNBL/mMa
1zenqporj9xgBaIx20nPNzsnGR3lCM5qW2X9KnL2BVgoG/OSCt/pGTz2IZo1C8Os
q7m3qgmxvNikDTkf8e5vFViYuYOAhMyW5H2/VmQKvTo=
`protect END_PROTECTED
