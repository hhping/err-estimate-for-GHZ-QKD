`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tIU5Kw+IeWjzNa2XALG1llmRZdaeZp/Z/zZOGGYp2dRxjus0uctU7VuzgDYZniHe
qbXSdBZQw6CnzR/d0deKChLSn2hoj5ieHHJ9wTEVLm5ZJPXQEWdmkCK2SNSinrP/
okpANQ5Np+JQitxpPKGR7YjSK4YL43i9kufnUOouTSKOPTRcwIH3wlJwasbPMU5k
2EmWHFu8beaKN/dDSfgVIqJmSLF274EWwZFCcYFT7IzKbzm7Mg3K3p/y6nQx0ujI
CtOqGsWdVw0P4ZNNPeGz52nQWaWqjRtcz1vvx5ovThuvc2dVDP9T43L0EY5cZSJ2
7bPFEhUvJh+kts0E+C8V34vZz7jdsxzv35d/NGeCO9xZc79Ut2q++5A0IxzD6dwh
pARYBquwGd2k9aGhMMnWhunXq8pwhuTsw9n/2sH3J96bRHc+qHYUUT57MvBth5zy
Et2K6ucntccm5HQz+FcWBBxzILnIr/jvDlfeU5qdXbbV61Oua+BR+Mf3vOei03N3
SvXEJCkbqUJmcx5MJaGCPTGgslRnyKsK6j8T4Dw7o6GJJu1Pr86E0p5eiTQUiuHt
GGnBEkDfSwnzB78lEXTIvFfLrmN577qcdGFioavtiQps4gVXoGGT+DA0yKKemnGG
EAHVPRzD8C7cN4GpMMU5yX05MCRh6kg+Qp6ti4CZatYis1cIbKGaxs2Ty5K0dR2a
AGC5TERJspWk0AJ2Nf6pTl5o2T7ca2YhPULg8fGsGawQaI32HUJQyVK+SWrgf3pr
S0OG6JkBzXnnnFkrRO50nvjkmxdXi3xUScsOr7pEeCfQ8CG7FvRQs5RPRfOhx1Nj
/y7qCSZB3g52ub3uTElJoFJOA5uCyE0PQPCCEYFeAE483pZ/zDFs7yi+3dFqXboU
vWBM+g/GDYI8jrNLGWhl+cDpKL7+7sRGrHQnSmAVHkfMuKNPLmSA/DJwqbUeHIYV
KAqIOQl6oi944l5hp7tEt8053NV0uLhQJWn/b37K0zVLnz6KYLzTTbOKEVC/7ljQ
mZroD/zzQlffweyT3Qgf3bQy7ztvqYRHh9zbkDh86+sO22mqrQZn4w3jIWKvz0o6
pt6MHbRwXHrx4fpEMXBc9orMNrn3O1PFRnhG2Sv2v+RlmjTKYEjMVDM/TT+TBmNY
IE1mGuIvWWnnQXnTyAUxo1UlG8QGsonWgiGMhHd9csbwqtzvoJCi7AXEUnRS/cBN
kcesbnrehpY5zZl7NYNtr/rxvvS+iC9xgmnyrSZQkH/b6SRkoOOt2jBqsnWnsiq5
8Of3qi6ZEoqc9+B5nD2997eFRPz66ql2XpqTyo7gelxPrDtwBlOCrZqg5uWdITmE
gjIMmrZ6BNAGjRB6Rr2e+xHD5ImAU0FwlY6PmoBJXVMQwPF4N9Vw9bOpDjzmrgHU
P2FU/3e4tX+i49EUMTFTDMMkZ3M8DsTElyo9IzepjeJAddMT3V3Uxi6nZMvGDFh7
kRIG0vPpkKkW57lng0+mSCMrRQfOKScdam45Zs2Q0wOvZcghSsL9gPf1sfCEEamr
xBC8PGfC8lOjwUCiIo2wi7shNJ1DIBC/NeGw9rbu1IGgniR1/CRA9qIL4piGxs8A
d3N4J+YtRgz7cx4wV1D1jxwV4+QSAKJmaKWuzv8xqModkNLq3j/2k1YpqGTa4UVF
n+tVv1PAM1H8zVo2HntLxpd5tqF+K9/Ywcqstc1B57/1nvW2KiicTm9cqFAF0R1T
UFg2bq0ABeRwjcuV56TqoJowBICSkiSlwyUGSh4wXpwha5SLrkQOVt5wO3EIGGCG
57owFz0/fHhrnQrF7CHhdpM5+TWUQL3CamIGU+hY7br/dCzMIL7jYdLdrbItuHIV
7xqOGMbv/qkc3HxYl3sf424mzwMytO+PNLyjLeSxZCvRj6B+Y+LXkJ2KcgM00p1l
8orGUbI3oOZi9oS4sGbV83SaThJt7hAEYMTfJD15llmder63/FfX/HkcnBAROX7f
jgBy8/nWZ2t0pIp8OMTEF2dAn/mrd2/5bpJlQ25r/nmKlMNMReedlk+ZGJ6M8Og+
owRZXB9g3RN8fz4Kz6zVttbdTULricgzEEHoO/cG6q53VC+nPV/ESRGaSLgyTs/A
Kvh61RDEzGWxm+Aw0liwCoEX3Nor8PwMDEjgTyuqAcpbIBj2azmF4sB5cx0iH3U7
KONPqy3miPLgfYoPikf/sVB/RoB35vtbrZAxVvB1OqJD8Iw7RV0N/+osdknIBYCB
elMBw0QjUCJ1OTEeatLNQYNQdeZ7Q8rCz6+u3mC1Vm8GwVNUYfS7TGGPoll+9dc9
rlIKh5S4oj7Lv2ii+6kbRaKOmDJlgtCy/vuMUfJG+OsZEXfaw8yVO0+K4MOkGlG7
L1zNCOmeHieAVnyrPJKSImJEngI+pp8YLC0M72VRDin56I3fFfXY5BII6UxdxKhl
wY4FbrhYchyH+gX2FBN3dZulDhX5Svqa/IpqicgDY/M/p4ZX3su2d0GoN3gqG1SB
HI66c/0LtsySncuaW09WGUp3pPulQXzcTWWh0PonnFiNCh7Dxup3Ny81QpKZ/RYT
WR7tqwllTPkId5spg4uvmo6Tc5IvPqw47pUuUdaie5Zq1pvxIshbMPmfXtAEnmmW
iSv5GFY0zC4edAE/tpjtq1zblJ4IqxDCWHQriVeR3ljhQ+ewcm5Or4LLznIhEzQJ
e2a14Om4fCAJVlJdUXDgS+SJujrgxiYZziC5frGJq4eAMNP0sttsuVbBdq5A34l2
Cyv5U9PQmBXcm5se9CNds2sAxkHkS9wZ6BFoFZLre9jC3xM7wGraUHW5myO7nwRg
t+F+dQ7nsMIXERjD2vj04yujUvm704cxsMGhr/Y7fQTsp2BdZxI1GpJPhF7pZS2z
j/auznuFHRqYqZdLzc3RlgSR14SulghTvHENkPdpSpg1BRMTnVmJ8EjU4At01LHm
MaQX4AFtTSbWC9SnC4gnZxASou71xxoHVidm75cZ9Rr/leyCEyrIWqxVQi7cnshL
n1Cw7q/79NmjCrZkG+aIDJH6n49ypgwU0T9Ux7irBcHKv+IdTufsCgIyF6LWGSJD
art5qEFMZb/sldji/m3B/M2QyPdxm19pqQZMXB4TCFvK5jbRXthRB6NhWg1U9BUi
+YrtRdI0g3s+vwIQN0+vSNncmPpvltrj/rtnmnJijREVe6r3xE/jINGds4Gis/BA
2Obj5qdIbVE9sYbbYCW0f77AR4UF/4BusrlWVe0UC9kn6m/FHcn9U0W/al+IY6Z8
K0M+lSlkvTSrCu1PQUhgF+UqUuYwj2pmbOXYYKNODriphxHR93wmOJdqKA1EDu/9
jYygwXIQswyve/7mqx+TZURw7mccOHtymms0crv52TDd9GTWQg+DBMHClT+ajtu2
ogEvLWvNHBJNHE9cw0b3tTpNxamyRNOeX2eToZEVH6YKtFXbGQglLZpfcnZ/VUUg
tCY77kDYZ6T2IHdvfQ6O9Dp4UXaMFm3CdBNTYFubLhIhs9dItbxWAJE6p5QLMtnX
od5GsdzMgZF4bVlOuY6U4AXKqxMQW7oCxzhgsHKERDhz1n1vdG7InNou5PBNuKs+
iisp6gKycnWu4a3bOTAJp6c7DvaGA6lXZO/UJADILOMR9XLICnXYcza/Q4gq4atw
eDJLUhsVnvJNeIKoGRCgN3tC9bzMSWhpakNGhTJOg9IwUPM/TUUh8rX9HMMb05sJ
OoC7OOlGfnhpSHYPf7931aztkgdFsa0QBe85t0IIFQEpEkmt76LqAuVd4mMUJfmE
9Y4nwMDf5Zmuu7hM+OOeH8zd9oOvl3gRupmyLQ6kKC5MJgJh2RtEiU/SNBfRWfXU
bqQpXi9RWfeItvEg6pNwEA2Fv6hbvz0pWoRQNYTKnvuYnIsDkSXO2GLpAHQPCwHR
/O7rWG6+U4ajvh7mtYfUWNPtQMVvVGYaH/GqszJ/YF5Ft1d56gP9eE1nfO0hf/HV
GdDsnmWxKqbPM4OmL4HPCQnKGhZ8reOA+WI3coFcyUKdNecXavmYe/VKvgp+T9yH
v65XQm913lLs5DTl4oBsmhbCsWrhUkDSjvEQgWM74inzogFn7KMJmiO5dGAyy7HU
KNp+rV1GexPH6CD4ost5LfpFwX2gjR2J4hV+AFzhlCju8zmjTq+ag1H4u4auUnri
qzHsYbk10GDea8zkk30Wd6m9F/d8+sHi0boP8LahWru2eA3sKMyQdV1/nnngLnlz
Gs65mG7fv0PnAnTmtVbZMsOorjaRpAcgvAOaA1RfxCMS/BqvMk/SXr11AWcJlNzd
/XWzbBO78ckO7eapibQeFb3SFl/YOyvq/OrtPLGOviKTJp6p3g0nnzOU+Bjp308w
26m9IoJEP5fDY4eJoPgZcvrgQ0tj7AkqqvOsKdWPNiKy+TtOzK5LF7VPoqtoFOv+
McLR+oPqNIiN6cPfJI8u8wGK2rfn5jhMedQkepRaQWuYgWy3KQ4Vh99TACJjdOfi
uNivJFXuOQ2h+Vfrr2ukL9nrzCagHTObQ1cYQrLra1B9/waL11n/TAUOseIvQgOX
h0OTupYh+P3ijWhvBlrIgQ2MEP81cq9YlWSR72TVKoE=
`protect END_PROTECTED
