`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtexEjquo/oVxq6xuJcXX4K/dFHOXhAvxv4aQcSmYg/xdOvwFmDiJe++dxyQ9ktV
nWWtJUu6f4CcmOA4UMYV22VV+4ta3YSbViNrM+/zS5A7lxe322Gh+WJEg6XPuBH1
puE2TUkQ3VXxIDka6H6ITvi8fTyxKqqi2IN4iwdYvmG9wt+2rP0X9BIPzOqLHybU
0FnkYVsD91/nf8qWvPhYxnRWJt+Uwsd6ZwS0eKUkjnczgjYxDsdr63Mds7vgsCo1
yosdNBI4ycsH4Y2OS7qmkUH5i0d1zGMKtnsttYCtUXFJwFI1iLJhT9vaiwzD4hlt
Jy/c2RJJCvkaSdCE+UQ8vPF8asFg9+QvgPbnVWekGFcOVzwTAP4Xy/qnTrCQWoLL
96V4lKk3WlrgQDO94Ui20HRVRfepLhVTkyOXQ8NNoIpomJPHmWwOX4U26eV3jfR5
vBUyVUkXQbGKoxoGDxfCllPm56ziWthDiVH921Rxc2+9/XwCM06J8BlccFOEiFT9
21lbkXoH5w6vc1aF+7xdQIXIBFY/qS/qrHfZr0qLYBLp2twhKGzuNI5Z26NmQyS0
xbeuEamnYhU9PqenVI42OOnEKnK00pADdJpd5SqHQgVrtjK3cN1rXdsAAH6D89BK
REyy8eGvZxYcdbUXBd6gwqiBmOq8mexYPbAFj7JzamoDBL/o7xRKSWX1Mi6BSew4
J2kTIIKdC9rObvVVnnVM+mrryO0rnbkHfCDPeKc1+Vye7CpAdr6feqfB81kffmJR
DgeNDy6xFWMAbCtV92akNSYs2gETfLd9KuxrhP5xWjgKmyhXgmlJexiKmeC3LK7e
23CR9mukgYGlS6En3RpqqiLdcUS19XFpkdWeI4VeY9o6aFvtiDrc0Stpb8ep6x/X
GXnva5JOzxN8GSBqRaRC8EYVwqq/j02yFNYu1mmsPgV0FkH2AbGfU1zi6BoOz2j4
z2n5BceohiAvonlsp5R611m8wC8dNhNrLxPEuhkPBdsth7bomGoWoG7iqZDglMie
mNDjefarp+52deyprBj3rdvN1Txoi1I0lm/SIWWTwzQ01ph7TbfBuhlO32va12oM
ZDBbMEwN1tad0Wn3X6IW7T68PBIuP2To3r8X03oFOgb+FyJS9j0WfvU1hsDb/Xue
Qhe2IPiP3HzGnBdL4oV6VzKfQtGJ3KFcOqTM1BKr2xYr/hzdJunpRjQiZcx3W3SP
CNvm+Cdglne0mnr5UnjxGHi2OiDctOCX3NeVAV6DfhG3xsOec2hqbKB9AWoj007Q
DqRnckelgw/Oo4czh9KjvGVe+glNeWBqf/jMXySa+h3JrxUSGLneo9J7lFepnIJW
NTEMZCyw5MTbckixqv0NZfcaYs5TgnKK1z6zPxIq6GXAqzHe0guswFUoBYlr+8LO
4i8TTk8hOFeBGN/uxpLrD0md/NSXnb/f4Ig/9EZMUZUAOHYPmkMlV3eFD49g0ZUQ
88epvjz6QLW9Cbz/kKWPuv4jK9AQF5QCxhwZxQPL3WQiHLbzL+rDqyvkDIhtaYOD
UtKtGysvlXOX/VPI9KN7tVZoHC6XTm/pF3IZJ1974L9oUpwaMvfNp+OnEBoJhafN
AF5qiQfpE5jfMsS63rqSuxhOgKt5bCXiSh2cyQgJIkdJs5zvNuMF1wARknVmKVs8
foS6iMzdvw5Kg25IsRWwHHl5PcdSCSNi1CJFLhdxXojSdQIU98LHhzgaDtRQKWmH
3Lamv8ehI8WPqcZJ80h48HPMrYfb26d74LD7+woDknB0eYsHVep2WsJf2ahSwJ4s
kGLc2I4wLukeozNl0AAinkroV2Ad828YVl6peco/2jnFIXgnpJXtsBUPjXOZ+8fH
7lBGPBjGEXVRun2zw5HDsVtaslItONaQazwtnvbIrbweSf3MZhE54Fm+SV71WjDe
oR3/RAddr1LoPMJR39v8xOBRpXawH8XaiXzGgVnfjIXOIIfRILfRApQX1zWDrkp9
Vbu9op0c6xqqeokywPuAjq+UJUCJ/1DP8fw03bvUjIAiFWi8HyLq7ubFrlr5uGyD
HcVSBa4xYUO3KQEw3H9SpxKvYRTd/68Pn4xqooNorYrYYfxqrGsA4j6Bu42qCsnZ
AzUBMKebavRyj0vYvvFxKrAj34MNbA0O2xLW00hb8/f4p6mDx2M1z60NbjVgP2XN
YaF1MomfnLwu1X+4yS21Ua2yzqA63k+VF7Rpvwt/8u3J1CiL9p82/uGC07hLW8Fu
EzjbTkPX5bMTNnwZ9AzH8rVPW8Ey73kiWLtzslBpLXorBPYjCeObFiSP0GwpPeqC
2eKNSFf3tMgOndpHih6pybHUBWjhB9tu0fTptR2yMzKHAMKa7cENTeKZT/JtX3oJ
eMRhMixdWBg8l4uoPnfQNCv+HC5pPw3Ks17u+om7zhnhIFsLQeSQBYjBcEyIHkYt
IHYqr684fZewqkGLR7Sah1hnEuAJkKAflUhq+Lgb8CTx6C3t6aPcT3uOg8HpLoBT
me+wRDXxva2dZry53yJ1SDlXyih3FFurwy+YeGB3grVB40+xCTyFGzCpJGye8UP2
kvVvZOW1V0WqyduXT/d//zAslcGYNzzrXTxjTjy5JaYq0IGQp5rbfBvyUwzH6/Ub
WicTKdWQyJAj3uFtVBUMD+AjvM2QnxOeyM6da1dvbGQ2cFga4RUdPceopS8IdQQ6
YG7G0RzvafXfaDUjK8SpVzbk1Kb+vKF56ZKBMGu8zK12a15MQ4niKw+xLzlCc3q1
YTT1X0Q7RFO2v0pS/vWzRTTuCwZN7LEz3qVDRvAmAQNEuuh9Jy9559TjWB7Vjn9f
OaqCsNnQIJgG/j43yLVwwqN72HACXjRUYRHQjgPavh4m/9JHxOhj80IUBq7OLZCC
FbQfZTIo6k79Pyt81X11sIHLNuTu490nPTJ2gKcUyoNTGuiL1P+++RHR9L15nMXB
6R9hJSF3UyaQFIneV6lJY4H94XoqICqldy9DKkLDB1KF0HfxLjc52jjO76uusuuS
nDSAOvV/CCf/m68i+4pDMJX08OGwIfJneszm+uZEOtDBcdgIu68T5muizw9QbJej
K5WJew8EFnslLmyC5Zp6R/36ZwUP7pVsx8NCpofnSvRRElwySWeXxtyZO8LHaV0D
PivFuNwUp/nLuKIkwPABvXHBA52xc7g7wYU9yjHL/b+wIheCbX5fQamBPKUokzvy
jOkxIT/ZWwNQyMYvJaT0HRFiROtQuWvse5PSt5FBM23PpBhqbU+Tq7xk+Plk3jG0
QstYAefTaZfh/wbcbAYmcZAAMSf+iSi+QLUkMmHtgo38uBZFofPaczAs2ZjGZzFH
4kojDTiKDQ0lCYbuY1qkhertEyrF1rOID82zdmtfgFHV0Iur2ouB5ep7i/819DfN
k7S1QuHZy7Ku7Srz9bdj41NjMRuyO8uos1JyDAf9OAASDwVa4VMG3Lf7JjP+C8I4
/w4Nb1d93JX6G3HBZGzoj4xZKOxAOYRDz9oA/CkiH7ZKsKCGs7BOdshjN0loyjlZ
RDNoHPjfOvXlzmbI5zGkTpmUADHp6TM6B0ZU2hya4zlC7/qE6XOT6Pyo9L8YOBzR
AJKrRj5fg0YBCcnfZIEWuAi/CMBGQs2Y+mKVS7rN8q362fS8xlsEOGayoSlKx9N4
pwNXMbk9mIim2YnAsstgF5u0yA/tpC8Uiz26lhtQcVZYa4TNK1wERTPuDo/bBZvp
EIrlK5jMyyM28GW0p6gccrVF59FCzLVSViNB4swNBqf0OPEtoPaI7klWm4XK3iGn
i6WMNIOSOs5ryMMWjdalin0R63O1uO3U10KJQVhP0NGA359wprl0sojDlWgnGWVR
ERo6JtjPsxTfVyLPxaclo1plyfTgNMpWnkfBg4bATFJ1NBovEyUEubPet0GqpyXx
sCEDM6jhkrbwwIBVuKrjAmJmtQ5D9PwVEqPJ392RcRuKY2ldM/GQBkcNWXqahEGE
4W6Id5Hg+VRJR3MYDfDLM/h3lzR8Dion6A9/BaRyVLbR4u49J4YpiGCs5tyBI5mw
9gdMJx4Q4YS1j4aoM1DQPJrIwVmDxSRmXIIgFMUd/EsZ27Z0kKz9RsFl20+cqPv7
`protect END_PROTECTED
