`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SlrNfMRa7CpjJmz1EEAnKzV7oYfhJ+yOX4+nnpYXtE9ylRP/7dudvde8EqrzLTsS
/YQyKbpRa3QSeV9tuce4rAB1rik8nUutyxgAK1nuvVd2wz3KgsHbsJsc/vdz1kkq
f3ZFyJ0Dl1Af+oK/ukflsAda1cX86hTb2Q2VnrU8+n6fOqezz6/Sjy2cUh7ce6rG
PIZ80QOFfKFt5ZJhrOrdbjdqbro3UyD1itHjzVCR6J7Q26gUajOySzRiCFoqF2Yy
Kko+Hi0031thf7s2Kf+AKE6ZWvQhd67mETQ/+ai0ghiignqh/T2WqYI48NjZnKpR
jpZkwSFa7DFA5Nz/TfpvCyu9Sjeo5MD/Glpwt2vtdLhmfEG/UfCk3IB49dZ5nz5f
nt47HyQbkN8ze2T8tTjHKWRhf7pH5UspRhtxAKPXvlp5wvEkFugjxfp5RjHxkCwd
qWR7a6991Iffu0G5O6EEl55EqWGaqcDFMe//86UldYxGHW1UlwjdeGVqeqZpBIsJ
lf1AuS9PxdXEiXz+7mld6FQkxZ30I9iOYaMq6eZrX4iGTOesPN1JXtGAG2Yy5vo3
pkDFEBhRgJIcWm3+jlCOTlhe0LM6rR5uSWSioPp9PDX5W6gYn0PVLJS+a0OMf1wX
23G6f6txo3Ri39ZliV2UR6wY7pKpkUCJjTS9VctcJmWwQOnlfr2NmBpYQ8UWPF4k
wiSltF/wEy622IykovNOFvnFpr5TPlV8ZObjPVHZ5LJu9QGuNUtlqAqhBAtAL058
XtAeMwmRCOy39OiyJyty7D/pVPT6ivQ6DRQ963r7blHzExtreath1dasZJ2dYtuu
wT2DA8kZoLqtZgF2q8JGtrcZD7EiI341ZFBADu11RFEMSQAK3/v+n4CH3pztrLfd
XL9cpgwTtynu4Fvc152Q0kXuJFWxjUavdx5dYlYOMNSMpTrEW9WwOtl85Gmh5+zN
LOTLbMmTnU4qF9oascMUIAyO7d/24MADWialFHPEluh+ykrrVoO0QCsGD+i0sc5d
IHnXLX5kyxoHQfaKOCWVT9Ef5P3R0nSlIY+skQgUtFYyd2eILYkpnalE95vOMmkE
seLqyf0xTjtngIhM5hO0QohxB50DpOWMl6kid523lqBwE3FiVnYhw69rKPNJGVhZ
CXB/c7N0uSY0an21jQAD4OB6hL6Uf7mXV5buPaiblM3HoQf3WJZRjUdrGvrKL+ej
A54exDjZjkbabCmT/+1FkxREXnys1T/swidv/PZEm12in1gsw4tq+dzEilVH3ri8
DPqn5BIOsYzibT4Rgju/qdVI/tWWdi+k0NWcCa6g39CLYddn3dTOlsBNU2SCX3TW
bmVjUzY/AuX5hgI5ptktr+xuRr33LHCO7RcbEfFSwnO7zaAeM6PF1VJnnjOPWLN2
9gcN+L8aPPkryiQv2Pa4QCq5mn8q3g7FgdTRyX9HKodLAhr39mT7zan7z8iNq+jH
6V16TqYgSxVx+X5EdliFdLKnlH+QUikeoq7ON76cwohN4VRWJBV8v7qMdHDG4q5G
WBpMuDVmsFUV30saFW6cKT7JgveNrA1PbYHjB3afyl1paE9PCMeMYdKjbup9gMoV
gb83vMBTb4bCX+ps0g2WipJsyinEDZ7KHoEcr9D7yNomgGuGb7BXGTxthRG2jtki
jIzvbS6nvgq5Rn6KlUlmcbF2DLtBcuNr9AmiubAUbd0=
`protect END_PROTECTED
