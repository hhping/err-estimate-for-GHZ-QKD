`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11mJDexiiZVIV0Jt/pDEXuqcagKmJcpL7a09zl142vZ0fPe3DjkCitcWeQNi81fk
/MmWmQnI98lfzhrkddneGesDxZXcWe2taYrYTID8HfY7Sl6bCcCnb/poG4CgDrtF
KI6OEu927nVOQ9p25ueaVemk5T2y7T8NSTga2b42Djj9bo6lxVvz0Bte+nuwR/6b
4TJDrjnamkcU9Fet23RyHFkA8ubZhU8lLyTGXR0If/a6MlaUb7/lKVVJBC5FG9yw
J1uYehgwkgN+FGOyfj6MaDIknr3xZ0f0wl5jwOh2R1iOEo4Ou9m7pySGq83R43nv
KQIbLUI7YJopshIQb32OvfMsBraC5J5/sSJsrMP9jcidI5BCcpi1Am0TJ4lPAVye
7IpWbpFcu0XNXUoHud8fN7ZrQQ7uJ07PD2MqHVd62tpF63YmBSjn0MBAEdx/+eaQ
q8EG/3lasNXjLC8075qqoK68VgvgbeHlR2iTxgiEeT4kEJ6QZEJma3qO+zZtfByC
f6NhSem7lXQYLBNAfQPTgeLaqwbCZlPOKG823gYBTGn0I6DLB5Jjp2kVandsuWri
pqPkHcoqjAojbrLKJ2RatIyRcxyII05PW7UPKZqqR58dSAwsJa63N/lIO3rJIdsM
znZ6U3HBBYtr4kgOzC1naZ+4DnACTK4ilZ+lNvcxblk=
`protect END_PROTECTED
