`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7YKQPNuLlPAeT2Un4CKP/bEg4Hvi/wWzqL+sS0jt77RZdqgTnjsuztx4Ng9MKyf
9NSlDeeRhAHd/GErEnm51WW+QLlh/m6c3Nr3LgEJFVk3hxum44zcspkhk0TEfKSJ
e6dln5OfMWasbW5hFNL35mQ/gdZeoE4K1s8OWYQ/hFeT6UkTEHXRJ7iRk8yoG72+
mj70agctrDKYBLh3SbT/Zxmog/Ah4PVAl6Xbb9iC7HBiMzhtUrU+wpqSGU++ZR2p
UY3hY35cBUXyilrIt0qL6OphU30qTnjFCQ9ZsUC2/bKJEZ11+76lo/289s3/xTmH
7EU52G7ZJ0mas+RS2fbj9r66onpY4HjC2aJnq6okAhYwpEuuza63G+83dy132LcY
PBxmyh5S491Qpob4YN5rGXdLg49Uhn3XRPPhVqnLPpu5sN0LOSrDOkL7sGho6HCI
jElNwfhUX5IuUSvW2bXUnCn42H2JDDMvvw/s8lLuFP0fsh2Z8aSpSwKWjMtrM69A
JDsMhODvT69eX68Q4nKX4jHHDTLvXkvMS2A0VY+M5t9hrI/eeIsZKPUQq2BdY7x8
T+Bfu+GLDkNCsY9Zmn4309UGe3SuszKXWLqEZPLRKcfyyGJAaqTmMoY34lxDjev3
VlYkG7iOMPeFh2/QoBMzIJ6+1fQUqfpsdUpTZQXpngCDkE0HGCID/Yw7PbNJVsxQ
t9xmu41CySne1kWci4TotFHM9RBNy03BQXnwM+hTfePVPa6NQ6nBjKn0GZO/i6cp
j+iEdeigqGReLYMkKxiwSgRc0i/dxEfehoJYKRtcm1faz7v7cBRpHfcIQ+IQbRDl
4weMFjp8fKuc7ylGqtXqJFQzfFrU86VCh/HgucRXzx8=
`protect END_PROTECTED
