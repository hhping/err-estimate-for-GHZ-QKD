`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MjBdUtLoSNYa3SH2sdE0/7qmhwnPvvbNC0UFVjy++LFFKJXXhvzJa5raUlPlsYNB
toWwkpezGRHlUxvbQanrjmaZHnQ6XubgCG9wvLDFqNgnT7FcRpaBQIqxm3pio2ZD
iQ0ZTtOoj6d5PKNq31B02nBL/ApjVKoWdPoE01oYI/d4D+Rl/D6iKnRouFOjqoct
g7LeUD7VuSD0yl/R0I/Tx2xKDeAResZ1ocAjlCx2XpCY7dVi5TVlWV6e6j7Q0kXe
A4+CXhzETo510koz8LYyjbT3td94sUhVtbWduI3a6r36VDME4BAKj56FCb7sX+1v
19x6+UH55e9GTRoCjGMGLMyZXnio+wITAi5vxioitBse/uGTVEKyYvpZydSvR2z1
aMEGTTkENcP0aU/VvRaGS1tXRascg/vDPAnWkT9i5Tss4YxOKUTbfDrEG29iJ6s7
hJ06OH0WbjG+yYoer3ETVAy2+0oUuYS4/+WCKGg2o3YHnbVbxQF0F5KffONRS0BG
QWzbAQRVrjkgC45t4fTLwB2oicdipss7M8v2v/7sqooy8/XfhD1ByeV8okqFGu/x
//vGKOHERTmBAyDZRNK4vnLVZPxrwrBBPMtoJIywWXjm4zkS2QAdPaQ5baS19w34
ZPqxLZfEiMdJ2KPaGMazbGH12JKWLjdUnjL52T7imyCkyH0b2PaEc572blk8U56Y
`protect END_PROTECTED
