`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DrDtW4kx6jclHE5hhr1+54VjB5auUQvqEiakh38LhDXt+emS9sI5WEx95tXbLKNR
qGaQFEit/EDl30O+4/FIuEA/cuUDWpDRfo0M1iXb7gkTkPSEa0v6NnR89dmdQfx1
bU4km+LL4SG1hMQleRcB7XCz6alQPyFe+f73PwzJuNjNe+JeM00QCDCj2Mn54d5O
fRuoZUXvLj826aKLekC8z8mN8xJ5XwUJL9hF0MS4mtK8SUzEuq2SuRXNVcOrsJgM
hgbZHRNivrJElM9n4LInZgODmBmL/GG94fvY2pr3P2i+V6940Y6LZ8pH6gTFnrCb
xtbRJehp3wTj1s8ylhm0lJa/kCvFRRjkAapxuyeX7idsczV4ivJTGmCp4XPwKsbt
f73vfx0u3Mmj8VmgJ9dBA6AGBCNaCzjsmQkiacVz7ku7fCjV6X+bi/qsrJYC1rFx
Tl7O3HUjZWTTZFmDt7hR6m+Suv8rN5ElYizScgxlB6lEL37qxv+S4kyQutKP/Xle
go1HWyGCk9R6o2PGvEyB8fUeNuopo6RbU9cvVGLrFle7ZMNSR7/U6cOaYv6/jE7u
S5+81GJ/NNhDfI4riaKe2+7+xZNBTD08ZFSasn5k6gjE9zKvuBpr2nwILDWsYbMb
XNun/3Y/0xNu1AJhqSmB6RkDFl5aky354GIrzVYZAQmpGK6OmwxuFAhtX9WNit83
MxlvBT4U+OowojhbFHSiWxitjC4T9LdAnuM+9U9UkfW4IOdI5Pbr7c04LhwRi/nB
4KnOhLLg/Yth/c8Lq/UG0ehlomrUvOJGG5CchQ5h9s6kyHl/Q3uqsE4yxLViQj1f
2m/8J10wfXyAwx7Y7tw893ybCyq0ZHuAsa+CLZpNNagIAThTSO0alPa/6rLLNXjy
0nkmtIQYKGngiIbBqeeBlYzk7wg5x/8M89arj2t9q7rn8OswQvcn2d3CzOnj/+si
HnZ1ZDO8sZzK/T3v8a+KDk3UMaNJ+X1+d4EwoXSmz79C4/Mygv9K/T+2DGy9AL1w
clIXzAArEbVp3YALFcardO9XD4S2ikJkBh4YkQa/ugIaMa+QIq7c8X+v/kBFzdSS
M1Lq/2tXTtXgxd+BN+CZ4F9odlp7DtD1wvfznavSAEArakn0+/H7KKjCRF+LPF8P
f6FXeaZkuK0BIdGEY4LmwS4NnLzSxWO4F46iTCOL4ZTsvtIjwH6uW127TOcNER38
68X/IPjXvGEwaFTyGQW5hhhslCHZb83G3V/Iv7LG21j9y+vxBFIfeAO6KUxQC8Y1
+e6XiBaIa8R+6TA0mtT6zAEdceDMuYIJ9mOD4X02GUX9uwV+k0hjyTDuJ+x9q/Ko
Q4iH5YzRg1FGw6iv/zaKCpqL9kcFNQ4q+0frNjWAjWZi6f2cGDPAtMLbTz5Yvsy3
yXEAAGTFwcvK3aj+d85dBeL4/49kTdP0PFmPDLJLelx40Xq/fo5luOTBLdRQpcIi
lRfcMRMK77btZwPgPwvoIZPheO6veDlM4mLhOfiLGxJN+Cg0wwIE70fp9PtX+AaZ
hrdDq5pi9Ktxo1PRFas2g6iq0QdoianlS/HiNTW4Qq0OV7uoe1renesQmaC303tS
SjXyggQ/PCjD3YEcBf5Hu0/4XuQIX5+rCT7iD4ffPiMxR/2BAkZe4/6YKo8ThEuS
T2V+cP8mqEvGrchK2mmHdunKpuTi2ewO6oH2U8+QAPRXX3gLgkP/J5Y9Hc7FB0mB
3eMpXiLL2V7mnyP3BCxpgliHD5ZVu8sdY0UHJSSUv1h83RVZAmEgIpRDMr7JAOsU
jvD25oJNEyEGRudkdpA3xP+lCwp6jbxng9KgoDayiv+vGr52toCvknkvWkWBAjbU
MTyhMY+lO7SUR5ASgwn/z+OD1MuO00JbYgjnbKcl1CGju/vIGw/rniNMCFL3ir77
0eDPzoo+cdsCq9jQGy1MnEyRtQfIsNaLRGMmlrvHhJQ=
`protect END_PROTECTED
