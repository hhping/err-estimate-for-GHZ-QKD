`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfJOfypHqvyFFT4Q4BgWnvv6w7/94ulqK4IGGikzdT7cuw+zTIrMZdsUwqb3Kv5l
kZgFHT1c82KsoV7dyZSiU2FhoEyuaFtolez/QZ+uQGkyXn8jD8S4KjJGc+Umsh8e
RDEJzV+a5hX7Mc/IMy49s2/94q6Yjm1CP/BJtRkg/+3lhdBoJ4CGI9wJownbPBRd
G/Awa9n4PIb4ce3usiPsNjCYXjNaGnQ+9qjBIA2Y3h/mZL6lFEG13g6sNcmKsdMy
fSl5WOryMjv0UWKEwwcFa6x032bCO5BXbVBthyeqqSZ7IwdIzFzJbGY1cUU9m+Bl
TZgIdBbg9ejKXBthpyT+OV8XwSiN+/V+qSyOkwV7Fn/AFglOZdEIP8c6YWPQ+3wB
QzEJ17qlSqA/pI8JiFKr+Pz06uBIEAMEgLC8ZucNnfmF4wMbh+eB0Uk09t9ID4UK
g8P+CLqgHcH1X72FjcBs1ltVbCCq5MwMSA6WYyxOQbq9ual4zjJB3SzzVusLViG5
zhFEfW44KS5vLceoRLZjCfZZ7wPFV3vriIjGPg1xLZJJPOmSU9hoq0SCyAZJ1dHU
XRTTFlNltQp94U11Jk2+cB8zmqu9Z7ydzu4O4zT/AW4VPAXMQKxG0JxMVAvuCiD0
bm3cYLEvrfvAPhWKfGVhO/xJJthoIQIq5oA3gb31wif9gnVxXKM4zZSENqv/BWbm
9OGURo5h4EaTWqBJuKCOUnQuC2lxj9SeEJ4fs8K75FvdVcF0NkK3iRFbuIV2/7cq
DFxCMV9pTqJ4m1BnnM2aVTsY3WGz6Av0o6m+tXuEtVyOfywvwXJhRqygz0xfeCtg
BhsLCIpiYZd4gO94CZOvWsv3Eb/btI+KjkTPYsAZkNWwe8x71LFXJKTEG4IsLNTl
J36p/iZ08uhf0CdxfAv65j/OTaIJiDWZVzVRPfoutderiZeWo4pE7AVCg3EJ9tBq
mMeinirFn+WoCtqtp6QyJM7WnhCGlnN9rBtuvZKdg706CipgOhzcbalVk9a8qwln
KA4l5HvoghlCuFRujl+j5RrYmonXRl3IVc++nsyDoOzL2RSOxMdlY+RI881zRigz
HGl2bSmVlgBdskrZrvvurNR57EQVYhGYK7pFfRODi14r7q9CK5w+m/qYYW2Jec7K
ZBB5UHcVio/NkmEjgUc4DLmzKD7GNoL5if+XTslkK+4ac2K3lWk3h1R/LoE5Y2fR
V6T8ac5DIx6Wb9O4vMTPF3MlirNVsY4pdwg/LK7Rza1SPi8tJUPDAWLFTfYJKJfG
I166hC8O1XaGnfp3mPU9I8bBbtnC7yYsZnPBuibDu3aCl3hdVJAUHBB6eMbmn99l
MaDaQue7ubRugjYq4Q4ZT6LfEOmR0AxNnj8oNA8RnkE9fTYvL3tlmEIJ29WxhZj8
uvPb0q+1YEDFJ+9f89bbKhwkVh6+eN3a9EP5WzDD0EtSOqMl8imXXVMr1rEpD/MT
LwLGMWTmE8ryPPrOmNBjXpju3DwhxJ+9WZIHuRPFPgFQ5LR2IPOBl4c7sQi2q78X
Sa+HjhatjDbg6PBxdinpNd7qOJjpJNWLax6DIKSj3faZk6Ihd9YR9pf+q9lG78vq
JQ1vEFOApWqKiJbuEpaXHwtLqphSmuBmKF5MdPwlb9IrIUFSJerlnwHLYhC55Mem
toNXhJPR356UkgF2sRPL0i9toXCmE4hprJn4pTKinDLL37OJztNqfMkD0nKQm+Rh
gngnZl8fqOcbT9wUQtG1bZYLxp+YnOBfiqH8NYm074Ws7o3p4T9JHr3nuKDMqJ2o
5KvSDCwHiDRopmGHbYvW3eNBRHsgbmKZWUcMlto1XB7HmmXqbTKaPtonhEapuUBI
M36BCXsc7G4/iIN+eugtoJ5oG99EHTbC0oRUfF6gGlToWJ3wRrlDB60QsK6kQlQl
iCrX1k1ECyKRDRrr+lnKYsKNyjpWTzj2N3svh4drWDM2xFnSFiGGilRzJ+Cr3kmj
q/DguQlKxOpRL5EE7aGwZUgicTDcVqYLWzWrgtuO1qeluplUR9SrE2U7VihT2NXt
m0Zb+bWKL1UgjGRdxYTciF8wpUZ+zOAbnPHp4OQgUg/nakJo+IqZjN9zdW3dRVrw
AiO+q4HRnfAseRcCOiy6RjzPk743vMMZ/hPqFaI6zJOB6RExH6JdoFsHxxRXWmg6
`protect END_PROTECTED
