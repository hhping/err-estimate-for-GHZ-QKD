`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PluqYKARCAcR1+HvxL7sk99jaLG3Gv7gWMyrYfqTYzWYQYYSo8xNeRpxke+XGfd7
qHmU96kN5GGuCdEYwfTBzFxVxjKgaMmp+JQHeHe/IAzd+kJ93nb0q6fELw0qZ24R
rMbI2mf8tcIOEL/jGKSaRXXpqrHBltFLa6gQMmIRU5kQ9GGfx60INWdt3JfCPADz
tgewbDjbXGDCCkPCq6WTTIqOFoG3gd8//aoBC/sWKAubGvzec6WKtTdL5Lt00evt
2WwdNWYm2wyszLW7uJJYYlPnDmFqNli2AfScS1RPZA60R/JtYWyeiS9ki3mMyqDE
BC8HY3qtsbUxf8AG+3AM7MC+tuZq+0v4IL0jFSGzP4DXjNdw7SWFTA5CjN3vQwyi
lmudVafS6gDjTbfla57cg7M6zkaZWsLB0crZouxcUDzTZJluHuuNFvo/pKX5yD6M
ghNo19Yi3MH+0x+PmSNyOd7Q0Kq6o/ScQ3uAvOIzRWC06b2SSxwe0QpC87f4S6Qu
h/DEuBXm02lrCPOhzsweZ5YjrZ8JjioMlpnMVev2QQqKghT4LmCI0VDA21W2oXhH
Ic+s1JCd4gPDqPZULq5opf2ZxGx5iY15FPHdHoQWe13msQYPKL1LTI1NJicKIQGD
gH8MW1TiiepPUZrbAahGricidO6e2ZRdw6Bt6vU3msvLc3oJPGqh3zA3YJKe/jJ6
z+YMVi+arZTKL/ugkkHYnnYyt7Rdsi4Ordt7Fr8DC/1tnJLq8CTUnSz43tJ0Q8Xg
l2XMNKwj0PvusVL/T3+Oj4KRvuINCoyyQ5N3q+nCoskNZZmOzKuCKz7SXOyRinEq
WxkvOLkZ1/6X6OUztISVSXxDenoT8HLROO8YRXPXCoVx66OwbkXycdTeoD90o3mN
IkXD3nSrSyxc5WoTt+ixwFPfk7dUmmDszS6MW1GUehvMq6T/+iqQsOqJKKVgZAv7
EVDmJl0yPJgNi3UwnNRRReoz18KlfbMgs3Gci36nHFcNqCV91MOG7jJbHG9BKPSz
mNStOxJvd5LuOnt6Hb1bAueZGTw2fmgpi/0QuZ87QUPRW8X0I1yUItcSqgLAwM3S
pdMfrmcVDdrpjQud751lM+p3ogB7h1nDV1Cd57+xwbu75pU5SDWLCqobmUKwAQYF
lU8sSwx0zwuUiI1d4ZVEFKFf67jKsLj2F5uy+FUn/CadBH7h9N04/ozuI/W7cqn9
4ybHr0Gfuk3NThUTjLCVy1ep7Z7ySvJXYQ7qYFyZ8Ggnv3RXX44274zyeVMMzzr/
IYpCDn6dHto7EV9s0ekqEccmYY6wYNNzdLI+/LDB3Gryrj6Btn9oYpRiMSggas5y
`protect END_PROTECTED
