`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMo75K5O4Xr14iaIWB7SBqbHkkdYmgRa8KNTPSneFQjGleHRJ4awLNp0hq6wecjT
r5S+wkZ9CyHRZwyz+8u/DXMYdCWXRAT9alvUip6ze+3JBqBn2SegJZV2IxLlOSCJ
vw3ACMMMOF4zxzgS64mgPfjQqbFGvzA66OLAFJFvuKwrPB1BLKivY7PCcA+zn6AU
tPB2OI2oSXYtsuKvjcEhJPcH2w/25lSxN7t4qVmPS0stszvtRHUFBr5yoi7WdvjZ
Xtllh9I43UxgTosVI7XKbqN9EUIgYkUYWbVi75ilvHeFQOtJWwMaQUcynALso2cB
bUqpR1kG2yz5TCEv61InsckDKwJ1Lpwuva8fKKy+ux4xMlcDDB8mK5dxjiP2naIp
GnLx+q00RJhg7igpDv/5Opd1jep08/O8ZCarc+31QZuJaUwjleW3cDHsNAb6SAIY
D2Rs6xdvqdvuu2EhEly8XdLl78qt9VustJYrPqHr/4k=
`protect END_PROTECTED
