`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6p+m19MbPaWLdgBRTqEM2OSH2RB3aBUrOm20F34FftkQbzu8NFhi6WdYKbWCO0qD
1tPpalJMR049KVkVl2K3VcqDp12TTp0RkrpjT0X7rLVKIuv9tE7l8NdsgqL1GU8T
oj1KkwU7NO3LD2J12KuZAFdL4zRiKlcXJuPtex841XzofIJHty8yLd+PDnAlPykI
vv//mT2BVJfkPa0pDeDTq8GPGmmQRXJHWUWMDsbWI2g03yF+e2pJ+vKS6vqhEhtf
AMEjyCL1byGnFl8ODyg/Dg9qKDo4c9B9QEqv746A8uX13lXZp2F70vO5dIbfFzyz
jwdldKQv6E1O1YbleypCEMYoqGVfwezcl8LZyizHeoIseNHa6v/GewYpiRtIqEJh
9Kdb5Hgj5q0yQxJoAuUQHzHldWBLNadthgTM6gRYPisRHCi4lIc4z09aLx5W20Yl
VG9uvtaHD66TJ/HSDpQVZ6vZzy4P26rRMvAWay7LQlyllcPKMB4ayc/DUEVELJdQ
Hg6hhNnqf+7q5m21nynp2qYSg2DY9JyJVrZYfJBIpO5xSu5lC+ZF8ht7kCx3nMaP
9fm5ILSJZwwhGT7uUuW6wKuijUUWeRJK6JglQhlE6O8vm52pY/bRUeBRi5jBHYdJ
/ofc7l75b0wu4lTCbULALBebS0vaoI9Wr/Xqfd4N6ZmyBwKpvYjyoo8OhZx0UTMV
9Vj7NbqbnBLoZ6oMbauXhqIQyjF8jI8dYrWgN+taldtMnxrKIOFiT+bWwgN/LV12
sfmc3QHndzY7dExaz+mJU0MR1CdWIXb9FRI9QpVdDD/KTypcZwQKMDgvFa4dLYXg
snRx9WV3UC1dS2ti805mD+YcwG0BokvmJ1+pQislxwSQ8/dNQ3BS5NyBX4+t7kC7
ldiLpYqHHHYHdwZm4LntVV/bHwKPgiRhhemC3OWaHP7kqANsypCSUzw2kfLVnz6O
OIA1gwAG1ZYZlv9wNfW6ICzFYxFxP7RvjT985zNk2bPst4dmW/ebTSTbJNIkYDiA
QKxSdYIymLjGtx+nYNcnloOTWWzLSUJQw2/KSVqC/8gVfKd8jczGffF8xVyytPlB
iZkSjEB4L2FmbU6raTc1TE9THERFnZz1a37An8rEh+qPk8flXTbxXHkSR9JS0p49
qcAQKa+y2ZCD2SedUnpRHZvvxcUvl0Pg6yEIfXPg3+WvDOPu9eIZwwH5iEE2n0Hf
eg4eE4j5uyeggTrP3d/XIVjY29Bb2zSxcBVDhxS10ZEBG2LxYlGgIvkQ2na4fBdb
Xbda6TWTzZvbRAAaej+dpkKDzNa7lUdllGWsEU7XgZE5Z3z9CZHtGKIZyHyFlp1l
jdyTbhrEH7/kMnAG0Q7v0dILel4x5Q18kERn3S70Dnn0mXVODbFSPczkldYQ0WMB
LC2C3opOoV+fu6VS02FoTB4XFEk0YHL58bAv/qR46D4=
`protect END_PROTECTED
