`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9nxnZv0v1z7d6hPox7Aq3QJwdycn0SOQcm6cqWbSNiSkbhu8yVReK1cy570UrHN
4At4x0bwU2P0JN8fX8E/M3Ej/jVOrBBAXtib0U9uuv8EWzuE+lvky/Pnr/2HycyF
Q1vatYizwSeKUdQAyesJbK31xMlV3DiWYiwxQKfO2u+oRWFQLJnQoFegKImurFTm
I4RMde0hDDmFDelM3pWJ3Z6lwVEErhti0B9VcWPnVpJpnHqV7NZKQ5xHPWjgXzbI
1lM7SG/orQUdXiIpasZb0T42fJXM3KHyDp+o78gDwHSB5BhosZqinToToBgnTTWD
4VZGilFYpzeHZvpNDGqTccHV38VY9mKmYzaCRyp/2eJPnyR9dFMNj7Uk9GR/elYI
6Dq7mdxpfcXhTozWfoQFDbUHDz8eTFquyiFkYxbEoEZz2oWTW7zUIr9ejdqWmgCj
miMvxQM8HuDiia0iM4rGmPZKwrDYk63lPCfoIeZfZD8Whl5po1QjiEmerkFzGgAx
ZHdkwxVqR6OoWzU/286SVdcL3LJW2/1Jfol+v0sNaJxQRKO1rFIcGL0wOJHArIH5
CsTk2kjMw52ejj8b4kQJ0xh9gov/vRmlKDmdic0YfFP2DmrGhC4TEBOktGUrKNTD
NENrEm8lwnrNGFw/2uJUzDJThNzPhvSYYeZIgPiHAbrApWAQkylRgbGQb1y/yBsS
uQ28MyxqeDyIvN5ku+Fl5jfo5SozyBEGlSNkiSu9hPxheh1HUpOX4S5uq0fA8nPK
sKg0Wpm1sHLoP8vF5SI/H0T/BlXUJqdhYXHrS5WaFwECtB6eNlKRk3anuTVHq4F4
Nr1UZuxNAeEnOu877vBe3f/5Bxt8ds1i7C75+qbtjwCk07ZEhBccHvT3VhkdMk30
u/zP7+1nCRJ+k9UE2jCP1ebmaSDq5K+BQ6OBFdujv8pmb/nrQwFcHH78/H5Lu63O
HZILMxy8yfA82KcF0RiVY/L0SCMjCGfMn5it4sLMrjx+1tlOh3HzuQaPLa8MDpRR
752HPTYQ+/gDDg0PBjdkxlN24e83OOkezGtL4RUHK+AUXlRpLE/sqWGSczFl2BJz
WpyTHsdwWCWfSm+3Iq2yVSbAfIlEQbQ6dxnsEpavIo6LLj3teDNYoRA6tfJ+NiiJ
vC91d9L6OgVItxEP1lbp28wnu6GXVgyRMLSw8GftrmfCUcza8wwrT8srbjPR2QyA
nh+LPyrh7eNrhJoqWzYOnpd3MaA8imPhnprUyQqNcHb4IVYW4cwXEyLLCGUklkbO
8izwRZn8ntneUf3f64UYkB2MweqwLatkLRseEgfAz40x7s1Bq6ExvSc0euC9VkUJ
3u4MOlkzE7DezKH8Ftmb702Ls8Y3XmTrLuWtOieCt9qCFYnW++IA01aCrTU3GaTJ
saERlmNAiLv5gg2XFAq0Leoo3PGkbPlhuBZcH43O1WWWy5XOD/CoypLp1mKL60YE
Fm56dvT+VGkaQdfTFLLusoEWsypGg7dYk7uY/k1MLb4T3hF7eEKDVaTeMk200QBQ
vMrPVRMOtqDLWTTmrjGKLMvBGChNv3uZPysGeeivLwQ5lW/BvM6iaWTg93uePDBh
bg0pkQ+s7IOXL0s6p+OWz+y36Y7W95RcL1iA4rJoIPBQTa+kMxqM+XuhVr9+uNTS
qkfNTJ/hByLhZQ4lWNeMfuF7pE44+K/Mz+iDVWqj6fQOK8LbMDnyyxItAbe1PNXq
PK98F4Z1Ob03uQHQtaLVZMXa9JwONpXQ4o5LSkFcOW/kb37dPHwEzC65bT8H74/M
NG+yufchKYoR1tEHYbbr+CrrqbnvND7B4E3jJ2JTtPgmsCO9FqHiEv0Y7JO6UW4Z
Q6DIWk8uIdaHf5/zJUmAA3qCTgQJNuR8v9SfJn/ZlE7kDkzHFcVfukIHuYg68tqz
cNtR6pnmQf1dlbOnmPetKRt6bGY3cYp2H4EJxdU0spW9SVheWqRBA3yuaKV8Jgs8
hgR2ihtlSRFzDVRqPkbRwButRcObUv19mOfDzXaEGInyIax+CpUi2YA10T9ukbM3
QNkIGM8Sw7YiHyK8Nq5zDTDumEjMHgFgEqq+cgNBzuJvkeIQWVMm7vpVnc/XQWpz
Wcdp6gDtYwyfCXRh3n/xYJ7Eh+iYNOJyo5tvYzlbPVEKhlHs5vp5ySdid1PlMdRh
urA/H/lwOu7gIQs3S68Gh0sBs0J/L0CKqbP6ZKIX5dvaXT6eWr/OhK08XQNJYqzq
APyIssS8BUlFgNzTGUGG2R6vs6jzU5BgeJ2YsHDdD6kCgDajsBcKCOAb4dWPdKT8
1SryKwdTtwLbrwvz811tHoWmduqmyy7tI4ceRBXrgECm2y+QNZ2K37/xUph2OZVG
iYjdBKo8cRdtcp1u5BxDg8b3YK7RlsjY3/+3k1NdkvaZYRVGtClpMkPX+GVCsTCe
QRyLv9JngzjbpnTmrKPousyvDmnSqJSJei9lDA9nJJrFu1Q8IYihkqS+2uJ/BEnT
apfvMY1nxLfgS/1ohgP8BmX22CgstEgPAaAd18P5Fo4nMJncnehUAOEjDDiMm6kj
xpSsVJYCvF1383DpKAyV4j06iYcF6EeIAapTkw1KQqiEd9eXhTIEw3F8X2bQqhMI
jWZtAIxPbMg0tqOBz5rhe4lpuFx9HmAiDdcNHwXf090vBptVtb7i6QCltf3sTRhB
FF1WSE7RQdOMCPgoNv+CkAPl1ylneDs6NVZ9catLPkTd2Xcb5N0bgdBSBpC1k6P7
THBsGXFA7avMvQbhw0/n7+WGBYJ3U+gtDP1LolUwSfi99SpLd+JwRgF+B/ltkjhL
jTPYg/X/wF7aS/AJbwTdET55IojFNRJd/zHNILuvFsS/SXAIR9UGlOuzfAvGWCWz
EqeqOxH2N5AZcDpszzDWRHhpRZq97k5JEzB7uIC8OIpASyYZic96R1F+zh41RoWI
46Hn4780NpvwgY7UhpxaSsRGg6udY+wsfJOOuuAe3Czy2BeFwKbcc5x5fJ6d3LWq
QxzsAzLBHvuOnptmnpJ5CvfiKAOADn+YA1z+GK5MrF4Wqg5TMtGR/Xho+9uORvS6
CefksFfd8lX7Lzg+l7WhwgfwX/3zDy1YwsoOWjQRfDiYdYNe5nVFcItgp16jFWAo
n4gDpNkaSSHLMveDmE3ffR5oZFMu5rStKSy4iygAlxEqBOsMkV1kI+wzU/m7B6Te
itouza5e1j088fYrx8uov04Z6ouEhATAMjylocrsRyg3w1pfruvUZkSiymx2Z4Mw
+8Wz9g2a9ufXJOGsNSE4TYKqeeddxdKEGpzQqbcRPxsFNabbx5QjIodm4DL1lDi3
1vBTj+l1JhFT8EktubXAh2YQPq9stnlyhN04C3JSLOdmxfkHL1SVN/Y8uL4qrvCX
1AQ3bABeoxFxy2UIzPx/ia8FAfwp1Lnn//j3GhjTFAwX+ywqJVJbg2X8u+gPSjdv
fVx7Krj0DgjlkxvoYIrZM+rTrc6CJuuRjBdKsWvGj4SdtRZRg6HnzP1xLmZZ0M39
7laQcvDf2pNhWKvYrVS37ZAR+ldVYRT8tBX6QQqz5DHlInn/lw87cQgWUMgMWiJY
+aubgrfs/Ot8UYaG/byTai7gqc/4SQgodVeU9WOlSnqCDBSVlogt8uawrkDrHiyL
zF4NDhesWsylRjFKMfEK0MG+qFb2J6/taquHYUykNzXHWvtk3Nnucsce+s8dESZZ
nRch1xyxHmu9dGvjpqiQEkgm/qybCP8twa1u3x8jnrMlD7TH2jroXK8IHMut2/0v
MgJ/j5CYvax5SMtekBnTGeYXmM2py0qz3bn8PHyNlPcS3eP/tGnbNYm/rcoxjN+U
`protect END_PROTECTED
