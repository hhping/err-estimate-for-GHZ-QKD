`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O5qooOyRdgLKeCGnqiHXPFW6Qkf/GCiypDh5laPcvJeTEut+sc4sMyMylrj5x1QJ
RyOIJQQn+RGlBfsOFtfdz2wZk0l0W0423sW8jov9gYKrihjaqmPWlmbdQjaCJyK2
wi67kHCvInuLgk9nhsw9utXBYD1+wo3W7Btg0PRJabPWlpJI6990I4W+KN330zk7
j3kiS/HGol+JfONS4JQeIjCETaaAxsNOv+8WNQFKjjKEANgacrEcuOXNO5oIZt9b
ATYNi9yUpU/0V2PPlQ1qp14BMDtRKyezlA2HIz2/kTKlRaHBu5fzTqS7Ae/Y/fAp
GocQ6H76eR55K8px/Fkj0mchmOu2Ccr7C357uPxlM2oOtxDfZG2xAyahxg0XFsD9
HA+nDUzOglzj6C10/D5rTn1UnZ/juGCrkJUkp1Yw+ubVWtv9uIJjuDmvSIaDATkG
+xIfxXZELHvlj+C3bf8Sb8YC3LBSU7e9eB0yhR94YjmHcxwCMKhTmJAJzx8DEEyl
cMrcFLy3F1PI/de4BbCx9wTB2xEtwPymwFfJyYOIbyc=
`protect END_PROTECTED
