`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQiv7D5Ae4tRZBsC6dBtHPMCqLJYo5jOnCCHm/Z/4q6p23yJFzWyJ7r2IFS81L74
tWsucT5eFyEp3xJSYOzAR2AtK+MVCDBDoomWLtHgEQsx5jb1ndnu7/cwhTvXXsAa
eewbZ3p/A3JnEegEp6kMoyCcusWS5Ig0juvrrMEhnG8j/9XLcQy+v34FtXHQ4qnu
33rHhU7xMy8vBjiJ/X/i7ZhF2VQTITn2XjghEsS904fbT+15x7MCa8y0dgk6X02i
ArS4ogSvMH+a1FcczHjvySAvrUOsyWKP5Sx6P66nwmUnJ8w4XiETKg78GiG7nAfh
FTjFAt/pziHU96ILc38TA6+heqij0oFD6C+mD6dIwfUZxco34N7XXLzN2TyBNXh7
NccmgjyakCZJBSdKEbYnX/BT5CRK4CVlTWAH7pI4cYqMBb5lYBu1tnCEQ318cjMQ
EEcJJcF0LKS6/VSmZ+7N9KPGbuGCtG5YYIUlHIeI/++OhMoh+9gxBh0h2kTe0CHi
7sc0hBTFF3a+ZeBlqNgLOFoXa8Bd1s7j3o0YMicp4umiOSsRsiZGuHPoE+gAUT4b
`protect END_PROTECTED
