`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDF5CUVIiYDO8LNQ//mnBiyZpibk+ziqGUQhw6nqZVos6/1w8h2iROhxVVRdDGsn
l318slQK3dOFAFwd4KjVEUnjjgGSZ7rGebDxjYm+J//TtyHPgIRrr0MqWbN9WoaH
OpBOmYApfykGN+xblPagubPc1gpF+UO37v5jlpZaSIkvvbLudYsNEbuj8L/t7G+O
ZWXpjUBp9T+ZIwA8qv8LshoNtqezaemF6RqFvVQ2ZbBBXtZ0B/9K8sHIshlyMnTA
fE+gSLDUel3gtKr+34bl9hPDMlN01TRE9O3l+91pVGx80AAomWcnsZnEofQQPlgv
XZHA4GjDCFyOxFpj/n9WC0BRRSSW0JxeCbNoYcvMgT2eK2wIFcU5h1TGvTjay1HC
VHPU6Zvm3Pfw4JHK8cuprVRzEleiXqNVKdBdQjEniAZqLBCdb22yBQg+WuxRgoFM
S/XDISd14d7zv1murMxJc8MmetCQmRnuZ2NKnH9m/2NIHWmDrpKVyCdtW2g4wVTm
sRnTadbunRj588xvLPQmD7WEsr5bHWCzb8qqpOtLkkbXCIO+CTuCRez9tZ8RmedZ
wpOqAnSYTNasutF3Kne9cfP91Ooi25tOw2UURSEYK7apTd7I7WgSlvNXMDt+uirm
BCqMIIBiSNpTWWRBMVNk1bGsD4Wb4EeShwJwxASLgO9oFxlDul1MvKmMoYXB3XT2
F42VstE8pKpWm9VHvQEZi6/w+9QNAGQakPp2BFnrWzQ6XDsISxNFHytm2E51ub9n
zkU6TADjeMMSIu1Xo6Bt/JOX5lDqgWfvIYWi64hqk1rb7dh6S3N7v5sJi3MPeJhV
DOYTDwswKOp4J0F8iIWtN6mBalsj4XEaVvENRCArp3aGtTeXWdZLW7RyKWkv384Z
NzvndFBkO6NEa7ZitjAq4ji7k4PmewHmBdGxqRdJLP2YFkwLVcvnwrUcNIRTIiZY
DQoZEjp8UtUr4l/GuSC4XpFhx9hQPFj4MaSag917FUvk9WK/NxTLmYTXPeGqFku8
RIbppwSIfqHi9o6Wvdb63Mo8eYyftnbV2SWggv1dwaXR3NaiWbF8XDifVucB8SWQ
Yih8evAV8JC57qAqpXEKLOvZNDFbadkjgr6PlgVt7NI=
`protect END_PROTECTED
