`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pk3Mhw5GlkPj7u9JMfsuqBXYhdJ2YQmXvYHP1IIOwSEsc+5G0WRuFS8jkh8Y32/1
yr1Ib1EKD7Zcw2s/w8QoSReua1EWRI2M1CGXx7RKr8i6KqynLBcMhjcU+j571lmk
wv2kBGa2pYcaDNdjEGPWgtX3j9SnlsGEn0+EXXjc+wpKqT3jL53Dh1UdQLLwUN3L
j2eGxq6aTOCI2BdHAdprirNzMFkxo9KYkGww64LpVW1K770cH51kTBG56cxkXLfz
KSk/4vUa+mCRI4mkDc0dix6/5gzjVHZ8Qm22T+q7h3gpu4TIpxmoC0pWpXy1Iwbp
zGd5O1P0aqpzZ7oTLTkLbLDzVj2+hGXu30BRJznXeW5N6yntphA+4a/c3uLMZL/q
qMF4gUAePht7AvUa/sohpJFFwS5X01R9MJObTT2pWIGJ4nrzsccpsdpY7YVwyTVQ
bHp6X68jj1ryrJj5KzIBfBLVdGsjZIHuq/MKcAETVxZwQVFYMP3YzRptBDHQgjV5
5XY3o3MJrO3q7fYuHztyHiv7H6gHDTGEv2vnbPRmLPK5yg/7YrbwrxA5Qv1iOlW0
J8cusnMw1XrwQoYto++6wH2GSiIswpYP/DjbtoQCEqGkCxX7M5CnYgkIzqR2ZZZ+
i/TdEmJtClDoi8bfEHAKUJFXv0hwDCzh50Cejt32kaUhOMcPKX+wtOpOjiNZSfFW
bHzmnUjb0q5MjbUfmrn+lbCocU2YuW9QOXllxNgZGlPh9/moPeXgWP7lF4E95LpC
PJDnAFEGnIjcjwvRZmVD+gG7a9cRORyJzRWYUp2TZqM=
`protect END_PROTECTED
