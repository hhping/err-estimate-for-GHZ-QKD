`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ae5TrBfkn/I1NdDVvh25Fs617czO00kSrzyPiJLS15vnhqGqOVOiLrJaZIY4eZdT
jTl/pkzZkJoGP5CoQK2PfqdL4vbjNwG1LO6QInm4VhB5lo/n0zs+NZYCjhH+OVB2
ETwTTI3sVRyVAMRN6tsQ3gg8N4DcjZuDIvk155drH9N6upKXoBsvQ2ND6yBbG8kk
aBvq9H4WlqQoHn3hhM1L/aqNfUthkkmQgi835Q7fKTRvpa9rft8jk2c/h6vfAKkB
DI4K6EyIZNcI1HVaS3DXkncQptbARWJ8DpHMCWUgfKfCLeE5g0x/z5S3+WPlFYeb
gOQqcvsMq9QTjGNOK5XPbh1bBDjRG/phtIhZMjNi8mdMNpF4VqjVosZc4wbzGCXK
QecPPQRLTLVNDZa+0uYqILZnVS3+KTJkzxmsP0vFqOI=
`protect END_PROTECTED
