`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7kD9SMiMIjIQTNNyCSmuRSKjkVgDU3j064VN2CTzpOxhRwSUDrcP+RWyd4rW71X
4UK3NDojCJGyG9DLthgrbQOFwRCNlBvQUGoVhTRfiWV//Oh3q8Oy7jkI/BB3zOuS
G+OFyA8+fvRq2GQ39HrB/Umdf5m73mEvHqwR07vcyT8TZritt7Rcvip4O0nX1YlE
7/2RjN5d05MWuk8OOELiv2kjiGQWTBSPkWxbOm5EXZOPyE22I4NdxAHw4FrMEFNe
A2s6ZhE972dcteONI+rpTNVwirhh4k8Ty/f3/yIZH8EfknAhaRg8cpG7TE5W8TIo
wh5MmKZOPYDZGtGijI+Z7gVLzH3rYZF1N0exODbTAmXPbLfinyOaiLyD5CsBX/hy
YyWsLIHRcCvL93oEh7RKZ4yDOmFLaSmtn32rm+ho7ujzkcywHl+OIJl+oXj8nPpb
b0Lu3QFh/sk5PY3VkX197VlwBGk7a4jRhSobx8RfZRpOZdQu5uh0Vnjo6+4mGJyG
zhIozv17KYqEzGEKVeHZYsEPGjGuEZDVfVhT17KAtI27ao/xAOY4i23SEqbb63g2
c3vyH+xxiEJqMEoe5I6rWTdE5mI71+1PgW7FLf8SuoMgqAERjW6GA1faBV+u8sDm
zq5BlafD2jtOYplLaVYZzLHceaRJZqhUE4/wqH0sENk4R+HKlHdgU3VCETXYT/7/
Gt/hQpkx/qB7L8YrW18wL0a/d8Umfx8BoQCHmbDYeT+EGOs3osWydbiFtetIFcXm
iKD6aMc9Tzn05m3oxywfbkl6RGUuCN+O8LgETyETsr2KDRx8E5Uw5wFa+MstDVWa
wBXSMmgoHfIiIq4nAXA7OZ1GMpfatogERh1LakseZqVOwHGJWLlzLqCwD7y7PMxs
WYgFKDME3hTWz1LhjJfVrU1/z8idm9NTuiQUX9EaVH8VtQSaBZvB5W9kd5/rtYgT
kZLhhEybih4L3vZaD7iVoLQMIaYzq76KtfPRG6cKHknn9a4b/Voyv/pEvRn5HCaB
DgtuPKUcSR5mBJI9wWmlQuHtdxRJgFZbzc1OyZkJFwk3joWWgni100T0oRlpxQ1n
aoGCNCJoaMczYPo+xJJ40JZtzDOkmJdy9TSpauJ2G2H89gVrzXVPJHohvGDtkL47
R4CHGCK1wag8j9mdWiuHbHrfTeNtxAy7TqqmRubPM7T41vhfBnQoMgQqdsEQN328
UE44ZyqK7VEEECespgXuhOJWJGNJ0pQt89rjELqKKykaPK4YIpdtoCFiD1PmAPRe
OOLhHCwowrIViPW8mVW9OOS4eF2gHfTOOda/sZH/JNrHX0rAx6ruK8b8AWpDyzfV
6EmFOWtXs+qPmfuhwHjwleDULaO1AZ+GSWf0bVX2A9FbQfsuaZuVdvMcXEOL8drf
mxf64qCIDt4rVCzY3V+4iR82TSFE95fKBWxdZAYsiXspbZlYlWJPjNCC3jAaCCyT
79/uiz2vb2JRN6jkIvPtUmLF/y13xKoPMIf8NtyWDVzchBlGRS+yL0Qq9yLFqilf
fd9+OMNLBybgh0Ty3WVF/XVTfiRvedMmwbIe8Ooy6HGFmv7ujIIRyndDB/PQW+o9
Hh8KT/pHWrwX9z3fYzjESmMj98fVwvvMbKe5tqYUkM8=
`protect END_PROTECTED
