`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2don6/qs9M+Z81g0wBMzS5iG9+B7dQkNHx5O0y1E0gOPJwAp6wBIdyCWAbOrsaRq
tlGjARc2VWmL8UqbIWByHy+iLVs8dZVj2yFRvQsyzGJJ4zVxU5pnz76W+g2KmGqP
tiVHYDZZDTfzKoUMOYBTPZ0dOOd6l8XtjPsYoi8C4PeO2+azierhsG88AkuuIwi7
eL+B026f1mbGf7YjnAZkUuEBdDZvFYl1Eys6mJrd0wVQOqoMVXlx+2ftmVRqeVQm
PHlm8RL91bWQHocSoVStKy9m78iDZv8CeRg7ZfjyD7C+c3kNFRpskWGurwio4tKD
sSVi/GboX+aLYM+Eh6AA9/6UaQkYXM3lZdFqb/0ftZUgAfhqkVoZzsfFgJb21sVG
HzolwMEaWMsHiR+rTZqzvA9m49lqktn74ESh9OxX33X+ol0oNEUtCUg86u279UNL
JCsdCsNLjUKVbdIvMmSjVC3ujA5F/G3xjkZaAYY7oHkJoEIDVJ9MDD2ipZQ4usJa
0UcaCWahZ5FxXNnkNuQORQCAr+nDyAOzJh7F5kHjj+SihKSZkXaHfw1m1mdOa2ko
iOBEjH7QCkBzGJvfpbzNWCRIB8gC5ZwfVH/UeQO8i1hiuSeJmlsnjlaWCWMs7/Kd
CbHZ9sna/k795PctEPw+hBFHlCWYGvPPI0z5B/OS2Eo=
`protect END_PROTECTED
