`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jlWO+52y5Or1yMGrGsdCtijrLSkkZ2othhG2CbksOv6IJjn9N5Qjk0sZJU2MzI2F
iOVtj+G2mhyM3rZg9FieA/Q5dS+ijU8drA5tejrsJprrZ4D/sE5bCxtA8QFSO+g4
jvSvhpXahFZDe3ZDmKpMRay4GrY/xuMPyBR+JH1ncSLMY4/XJ1oLdGQxWwXs+Elx
/io8yU6+zNRfxDs0ofvBg/fxuQgCs0zinuPmjc/AVLxMPfah6M3nOX5eU22Ja4lJ
DErU20rHCF+xxPYyoWCDZDVotK6a8e0+84OBM+ON2D4m0C8k5IP91ligxYKHemFm
o3E8RLOQO4MSqpsYM1ymwgYOeGcCq1uoTLxGd/tUA1Mlz2UvC9f6g3/ICqHFDDeI
AUrrsVX3LNDUcBoqYbUuRsoj/w7F+seWSrNtn2tJ2FGFbqswjP5wkoHdJeyTEBtD
zoieaA13l829guFCnAapGjHYK7EaX8pAUnGIB3YHu8h47i/675m44UvpCVuA28X8
M7+E+m128SSsEJum3dD97ypX9dX8wyiymdQ+afluJjJR3TxX4LktqPkih6RLAfUB
IlwtZ7lUdbriQkSDB7DnBA2sAuV8//ZMg4ODpnC/i63rZjcpwanNrvVLomU0MpRu
90Ex7owgAhyLNaSh7XPI9kZt9F1xtocwiyJ0x2Ga/wcP4FjaJwCd8r4Ofsy+LAmZ
PyJDym1Gz3F4CQ22XI9L6u6tj1djIG2gqFJiCRUO6oRNVtRHQQKU5C/FuIsc/Elj
tyP/3ypFN7BB1RvJOYXZdbxk4dalNbCnx9qyLdXu9qiTaBz8TS0T67GIjh6J0i+I
zm4188+98sY3KrqR+KH+36BvSFbQkFY0ot4MOgd8Wu1nRlEjua8AZgNnhX670EzS
lhRerdzgt117UJtahG/v0m0p+4Fz1wtAc7J0JzDox+vnvWqKQYGN1k/ehpAVQznv
2g3UQ/c7k4HBrm41YUlGHFygXgQOnLtvPt6/yofSSjKVwzxcMS09fNxQoppBghSW
TPDfVQNLOzwh7/Ezd/mZXRthrD7QSS2LNm2TdDIjdZ+toHywKWP3lg+Iq1WxZ5S3
LshSi117tKyGHPMCy4YTfCcCccxYZS+s8qw+9f4WndZSXjfTDpXP5cMWw8y7WCI/
LjYhHGarRGHeBFjrZxKaZGfDIudXnkP4169WpDjcJ54w6S5CQzez9S0Y8qbitRdB
3bgIf1LmDey1UaZ8WAJ8GukxSL4jFw3pyj8eKDS+kkpRHp05CexHP0sKzf9XiwSt
RDHg5xS0XSPNQ90z7Sz5Avs9e335XNQ87X3sp7E5pZDKP7cQfKr64ySMnhDf7TQD
+y0Nf/VIqLh1g0f6NLwkoIwkcBkr/w4WnnJ+VOJSM1WCHhUys9tTLNgHdKfHxf9u
ktakb01pZcUbiBUAcnoCUtSpNKtzBc3T6Wqip6S9IB9PQcbGpKEeE96EbIIBrXVG
KNCiv5t6RBijzriLkx3rqjA/IU1RqUTkpsyumC+UdNUoYb7C/dk5rdJv1dXi0Onq
r4aJFwZnF1Oo1hDsKfhOwhydy9vZLa91vD9HuOGhiJt7FtvuMoADuk/rvIm03nhR
Q/SP+CsPARIG2xjNvmlGKMRoO2g9iDhsJlS5jC8cKBrHItE31c5Xeqpx69DtyoQ8
HkV9fnpmvcYdTh1bFCq8/8wXS1k5FvtfzQIhxlKwHlLnVPLY33wYsP3GZNVCPTJt
S+fz3GP79ZfbeFPgIktzjg==
`protect END_PROTECTED
