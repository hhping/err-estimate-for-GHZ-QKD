`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k5oxZo0MBm/hdNvnL25nppTN6uHnOZ3MT4femCuaFjMnWyF83pTGPwOPm/+GT9eN
ukpYlWr3S88bFhH+uIalOiAX7z6bN8LQsEb5aNG5jQuUJSeYCM5r3D4HYTvASnQC
b25e/ckoLumeLb8aBCgr1UuyGkaYt6LsYY/Hqy3X37rL7Q9fw7A5Rtt57tvFSRJ+
T8zODSbAoXN7ZUUtDUAck46MTaC8K6gToZz/M8Jc108rQG26ESYTg2l4hfNl93g9
YrzbIx4R1KnJj2gtjImx7jeBEMS5nzS5Ewyfp9xYGG3Ogj98vOX7+kkvlbHl3vA2
rhpxqf8I+3nKPRf0AXP27ixYr1Of4gfEI9gk575CNtPXJHgiYyPB7zwt1XoCXZkn
xS8ujtrXd1qbfr2mFAqDirXJB7CVXMI1DQNs1IDGLE2W9oOj5SJYSjOEqRp0YoKe
W28MLaqYBsrzQkEcbFKpDLxR3fScTYeq8FBhCQyIg8J+a6EyovdcIKnM0yz+qPGK
RGjnWiHA+trMtn16cbQKKDXvr+V6jeIyJHC4so1cfIX9Tq22DekyDg7KUm2QdbDf
P7cJH3+2dbcqFO9gM1TP5vbaHeo11N/bHY4r8LB/07npFJ2F1fCe0fTJfMIQtJYm
RdFmEkhM4ioqRSbOnCpaLCndqbG4T1TUE4JiNfbyAYRlHutng2m9smrgBao+a88n
dcVTh70SesS3l3p9QNNCW5pqxs0ndYTLoQfmPryeQmohG79jy+KOVG8GBDNLLO0g
wtmHvbTCLmtgyLTzJkpUUh6Dv8fc9ORv4FmOKySe45K3rWqbsIcZM0PbBb9O3TAW
LmfzNAVEmrGRszMXKcmBsA==
`protect END_PROTECTED
