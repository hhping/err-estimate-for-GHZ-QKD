`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1DVZn43KHQfUhL+EFjYbW5+5PRLzhVIFpWVUOH5h0ZzAIGQBMvGZpFC8ov1Mbwl
CCjfpMuFa9yg7CaI43TvbJUp2DjDdoQxtQmaGtJkPtFsIRQCVViGaEuKYFVkSKqS
0hYlImPtVPiwHQXMAH692qCpt30a4YmUL/VHgfbNLPR84+MGTJlBVreZzxXzF+sB
nUS1l9qinTmAdTHfVcrYNiSv4EibYwLWQblN2AR79A9FfzMoLVxYNTECyVp2bu+C
YAvkWHA/ORtp83AZzvLmj4YNfckzKtZo5qzZRtNAI02NJCghSWr7b37fWernKkDv
JxxGhwrJU/CdXvzs7wimQLHkh9KuOkmnCf6C663cR8RKGKKsrEpCvUUYVMYzfKbn
RzfldRK2xVCHPX9PAijnL8qLCXkAWYvfhWc3r8QNlS6SKB8v/3VaLTaIy0JYHdXz
AZ/YzbihhR2swUwAIUkXSul4fbnnla9R3dbiWeArJXra9sdr4jP0dSIfn6wYOuJJ
sSOHr2ze+0Yb3uLgObtbOuP2+1dILf8rbnHa7wzeZ33HWFUYwouIdcnmjyh5ulya
Idy7aNsm7EmQU1FzQa4oxUxZyZXtCjREbDWNQDuCNQ8GJrHvbksp0EJNi0dBbC0y
pVtTgxg26ONC1MwD2DiNk6RiL8Ywk4z7RZb8YSG1i8dMSGCpzigRE9kapcQNsgRL
N4WvlbWj2qZ4kWYWOVwN4Ata6/1Vh9XpJOQ37dks0/6Set5cACgrAEeRtSf4DPVC
WH4wWEMr1K4UslmWdM22r113AbU3gK6hPvRsRiNjOuae7gVdVdET4kdfknTjDYaT
FtDnj8n+91GiW5YtHTFnz9ad/5PoqHN3ghrXaDQK6ulVCRivipkskJb9P/mJVn+t
ggGea/ik9bo3uLJI5uwWFYauFtmHJa9RNoqFE6RSyfJ0w0ON2z534/i2zIVDr54W
Ucj2PnYkjACwwXAggKDI/2AukNHH5fSuwlgHCuEI+cQ7h1xWT0sv0eTTg5Y5uI2e
ATwUzhzyg47lyfHIOOSJBpWhkZeemHrQl/VkV9i0oRYB/rjLTWZd5WgPL4kbsHSW
wixa95+YC8ZrMzMaMcPLhmyTiCZbMdS8v5vPPWs2RQrMYoHQzJEiJJK9/mlCmz0A
unDIpOBPvAn/jsAxYOUQEe1rlDoBoFYe2+Rf6RgSndtlXiEvL3+X7GwWKM5O0HYb
dpNiW3F2QIpuwfKkNt62PIXgtQB13GEl8znatDaKlHEXzBI9y4AZ+1jVFHJHlQNe
+P4bD/RMQKD0WIuW4o471LmilhxaQjeAJLfD7RjkTfP3frSGSdltsYO0Y54US0+H
3oMNLUEnQQNn+vSC+BkOScUSZSrV0q7g1CbkvZv5QnAnUndCsioYaPInMJ9jkjgc
wF/TBbfUsg8TDFgM6/c9VcYA5jVpvQi1tk0yRSKfvCLqvHnCpS1JIKHTlA8kMA/C
mf/yUhW1OI63wSc2yBsaundQ7dDrrk8bpcdrXHomZZaW6Gx2AeKodvA31nGq1dBV
Ow8x3H5NQvuyR7hy1exK4Wicjyg2MYH61jB/1TWvwhRzAMu5L8bULlKST0KqmYn8
8SdbGV7RoTJJAtFhRnt27VN1NsMcljI73FEFVusjzOaDkbufVlDLDg3KTbMA7+m9
IkCaJUwaJ0IEti0CXCqU5Ze4BcHHlCqw7QXhxtZoF6BmKKiFh/xvKRbnyty+/Se9
HXV8aSXF1JvDxDPAVO435G6cxTADkjUgnSyipKq+8O/wInkxK3+SaCO5De0MGTNB
hm3XgH2HDkglBsfIHMOGnoXgb9rxDKCCCpSouOE/fk8YE7P5f+bzklk+PwUfqWQ2
xl7N3cIpEo0mJqmrJMvaMMbWwEpqrVa6HYLXAnFIinKcs9clfnsLbAYlhDWtODdp
mMO3C3I3Cv39NG9+GoMqwNpSDk5Fj0sYDwyjENyBCEH5M+lHkJCxwKMdt1IxRWvz
giE4N+qdYtF6OFgaTidqhf9uHKs9A3O8gdMEjTUDKntUjC7gMtWX6ZmH0Cf5UFPE
QLn1wam5LBi182kooIvXyElYW8gE2pQpuCD83JLDLDe6m66xzS6JRZ8U5BTnrqsF
9dPwvSlL6mwq9WCE2T0qoBWxLDz185eKw7vePLjfgMTxaL2uvONdzO5KGsdUy0ax
/TzKWgm+EhSwle0T9VqWCfEaggZptlHFtfAUQYk7lWmGHVPwDAAe04fc+gOSJKD+
puZrBE2vvfie9L+an4yhCY2BIr3qKeu37yk7Q6PDjDO/KvzfonzjF26Y+o/4t5rA
kfp8TJCZ0iNcjoXU1YLeK3jrJ5QzX5pAZimCnjW7Zb2DpO1FeI3L0pwTH+UB/I4C
4mp6QXN7HFD0ISRxSfEenA==
`protect END_PROTECTED
