`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ThiVcAlE7Law77MxTDTNMZplGRpv7bti8aPuHc1n8ImxMG29zHNmd2mNn8G6baO6
dKWdp8Q3FihtXNkmwdQCaQ9FVftE1P83/ZnSkRrhMCBnZLa1JOQ/bfjEjhArU3Qg
LEzLGsYtMvEaShCWlcaFC6IQXJvAk4P96pdbLbRA59MxFttO3Z0za8mHsZHDib4k
PfIDg5MyURh+F23PMVqzY1kU95aFyg4Pb+b4qIXR/0C3TXFoSQls72KZIFTzdUCY
hAYwyQ2dG7eOB5YKrgVWKyTX+zkx0hDjaTnewLefzHqPproYSE6VVw3QJall3Lbu
oEBaJyWtH+IEicIQGhdNDSG5h/L54QTdp2MPZrUPVVQIE6XcWR4J8AxcYNz7g4cg
dMxhZpItatxhrjigT/ttp2IMJU/t9NMQU/u1WnnwW1+GS69FHkLxf6wT7pJemTVZ
27F293T/PK7e1tvMNqr49Tg9CFsuvjJNyVKJgHeIC1yKGCS+oJmZyWDYZ3HsWgSA
spfmwaVmyasZczzvVCEZ8CwANFIHy4zf+Q7bdL1wpBLW8KGwqCv5fOIobLjLqSvI
7Q7J7z2f8EtypZW2x3RmI6qqvwMhoCFIjbMrD10h5cybLPd1JsGwHrxrH0SqIpgY
MmkpPM46DGH4r233bH8JxUoQURQfXyw7cPnnI7LrTGMeLancY3x2fV9+zhPLgWSF
3XU1GupQp5CXf+DNcxL5lADNcde0iB8EUkY6Kyxx30T+2eWm5za0EShSoxGKQQKk
LOQQKitPimRw8MMze180tOCQ1C/1U8siWyIMWHMOoBW7h8iTovLJOu9Qh/ZmaupY
ViWal+WpKP97lDKrr77/NM4ATdo/sK3vua2jWLADk6xbta8Oyzqr7cOkCvQppnNb
7DH5ikgskTTOiYab76J5K2sgl7cv0RtlG9v58Ys8TkM+RJClQqaAoXJavy7mSFxQ
pvObwHONJgPmaQSgnZx8fvNVUfSrcUPY9CnI5W9FjzZw04qziBm9IHuclBLTy/QG
KCbGUMQbEtg41XswW5h15XzCvHUzA2oUTg/p8l229C04Czc7urCvBlIfnhx0ItHK
OyxiHc0kkiUa0HDj6336wDNY4/a/4+6wG3usbj8noIYmkxk8tcA5QPdMZi99Nz2I
HbcXw88/rmchb7JkW7wYxvAD8JiTHbAkpGy4SM8+Gcb2hpUviVRiJ4VBFwYRaMly
KI1YVa9pa+anKBPtNFfHKMwf4O79hw0zMy0zj7+FpEyxQXwWA/kc+UVA/8uJwSGj
PiXKvATsef/CwAO1hEb3rN7T55DGSKNkBLbFhelXWrpZTzldXptCPcXDRVsGXqkg
zvAw0pSPq9AfCuYdCreQkrmKArb+kXbVJIZdkO49jqz6QjEq9K2H8BRzNhEAxBFU
LiB4ZNKKf1g53bPz6OXmRl2al9tRzJlZy9lMgT5qNIHdDIIgn+A3bBDHSchGW8q6
2XOqz8s8bG/hwWZ9VCKAiLjfILgFdK6XCIYA6DoxbHWNQUJGzAsyyKROuGWwgeSE
a2WlKd4sdblBaeE0pJ5kn82gNUlyZssV5nzAd3d6syQNhiHlMAZnhtmE8jfqoYv/
eydJBp5/D4lQCKhaco3jpQqz9eoSkHplxvf4tl1VQgO5NesDbUTMnJH+Qz9AnNse
n8UuUuLCrUxMgP3VKB0QFl/eFttQacx6nX9xEHH8ELV94oOftpozpOOZiOn3Pha4
Idat9kmxz/hEP/cXWWasiTfCphOImpk+CeBouCcUfvUSFRPKkZdy+QTlDcjaUjbs
oKUlQuicjncvjMwQiXRB+j+ZzvjFDxoUDg/gxr57ckGfmcP+5OkdrQ2pboRJatWF
VPQaRHtW2rM80vYzwGx4nWFAhdDc8oUo+jCW9LNc1eJ8mTA1imrTT1/9pjbr0KlN
/sucNGe1EMDnRxLhDZ8kAQV2d4Ca9UrihDybyMOCoCjAnwRxKWMkTWn1yAZgQD56
ka9+3gB5xvW04tQzdxMoLrt1ZfG45lSlJXf+mC3zeT6USyUMkvH4Z+QLH6Px4Bpx
UUTJ3RMHnQ6U5HZgczrcKTAlf7dEQohiFNpptma9XSt5kMRe7Da9pJZyRh7hGMny
F8InylR8qsrBLRkKnFhdRoZREY7x1V/tcX11NStgfGs5mDSUva5Fue5BQ30YNPdk
Gz74EkU+UbtdKPgsLnSM6Wndgsg/lwvpB7jqmYvRtjrsPJxyabaF8bxldvPSm81n
B+dw4iBiZjDwGXL31+Wjb3cKmgpSm/jinFXNtpYvJvZ/pF32sG16ObWq3i3qGxJ4
0rI6IoZsPaOJCsf1LZiPk7p8iebo7DcpNpmbEUasD+VRbHkymPBDTpwPpvaQA9QF
VJ3612bIjTI1hQeVehxsqDvI2H6Fz7jv9wlyelwkwAKx6gD3bZedNuOwUFD0gDpq
66zn38N0m/OywJHUFz41g8Zkn8Kp3MJMzK+M6htOElYwRB1eiwSCNO2CHT4JDZQY
c2RRg2ksuF7Fa62+uVYKvkZp3gO/IzjdxmsJITXArLBblog4PtwdxuGMfnXAko5M
/0+OK9ALgQHGv/x+0NMQg1JhVAQyTU2JmUq9qkJAjnAVu18SR7xL/XG8jLKTpFrk
0yz6sXGb2PD/FUVLY964pifs3MyXhD/9IYk+2CafffKqsvBR1AijwOHwSoOrjOLj
w0SsAZVCj6ZUj44/pl2C6lQiOtYZq7sAsr+m4tX1XDU/KnoAXTpMRp/AoUsJ+XWD
E6YexX2lz3c81l6rxPI4Xz6Ysqzu7aGaE6S3NyIS2SQJFmX3Jx6ABmatYMVAflLy
5db3w/ZgBbL1PtsVqxiKbemyBUpeYJU1g8GlNwquCwHYZLbph1gGfUVemR/UCSG0
RIqdBtApFO0u5HajIQD2RQ0XhIzQBq0dGLz+Cqbv7aCgJtrhue88hAgNWbG6eA01
PznHuJk9ZSc2P3IM7e3AnQ5YYXUdaM8mx/3kv6KK0iRybB/o7AeCfu90nx9TjkGp
G72wz9r15zrxFsGr/vw0lB2h0VkfvNlA4xvte1pxYJ9WzKAyuNWM1MYDepL0gRc2
U+Xl6UUUR30mRcpu/ZEJlRbow9hb+aLgwp9fdYk4pl29vcpBtz0+rDSUJt/F+HGw
6y9t7azGp02JEUERKgKSsyWLz+x5X2EErcIkRffCpYjsbKby4c3HJI0K4tU64tym
7ceC+DEsCQcO4I3829otWQySSXwiL9WZyj+Dxf3SR6l+o6iLdBrPU0CsHr5yS8aL
Z6lPL+kVcoREIMj+SS5v7XUA47McXt050zJWwpE2/iCIVS2Q6pLYYatTy7tOmJhg
g9OkZAt8bg29zJCZyB6i/ZYGSBC/gbMvlCFzCbeD2Ejt0gkxyWkGU8xHhtUEtAb/
2AQfLpC4cgoei36HnkU33I1vUOAs2y06qtS7NR+BG/tRaqVq7adDhT8T4xYLKoIK
jwHuC3xmAzIoC9S0o0/GQ5zXyyLThBGqj1pYxcyKyPDHiQz5YrtFnajJJfkjPgXG
PA973BfTdCEIYfa1UiyC/NSZcxvQxpS7nj0NrJUOOSctBcfcl05BcWZJiW++MHly
S8GrT2ZtzhFHztNC2IK89vSpr8y8z7pRyCNodpbOzB5Dzo6m8iGoQmo9g9AzOSe3
h2NqVDP69SeRTHt5VlnNxwvmqFm+Jz+1YxXExGaCspIEe64isnUEJpYkwUmrpKp9
gpbzzucDhOCcwVZQfWdzR5+gGuh9mar3uY83CBJUTqXriO/xoN9mHVA0FWcWRjl8
q4fBBwrOzYFfmMyxIQ24I1HFgxzCB72n2gKGm0ZryowwNg5gHxUBm2qfy0J/hbFP
WA6pxLoix6Nr5M6oVUi6TzppJZCJLtqONxpImrUyW0Azn4ZewrGZFS8K0wf2L1QB
qf0TKgrLBCFi9EU/UQaiQKc/NvjMYz9G1kXv1aFeu0tymuZgb/HXJ+w/qQmSP2YY
NBmBJ2f5r4kvIAykAHoVCom0zaFjkezqeMoaFucQxPxKYBslLrZEsb0PPImwYN2n
BQj3NiW6dFgUavx+ugiXZD9Vtv4hN47YK5q4pYLDnhnRE77BynxWMMqtXvJ0rYsK
TRDVSgD2Kdi/TNJeX/EE5iU+TIjSqRe0oU+ua4iuzDMYk839B0PJjyi0Jc4EOiiW
Nc/8YS/O+gSiQ8EXalIGPUK8prAW4ym1FHVy71crcGzD0+9ZD2hXqvgn8JZKcHYB
kgsYzaC+D1gmIw54GRjGaM6XFfA3j6dvuLbI2pJh4nU1OEwU2lUcwmolTxxVkNTY
E14+vX3AeHYxvHj8Ujxx/WHAjCFMG2TaSN8Z2LRs0WOJrYquAyR1zZO+PjsDWjwJ
Mm79RP84Tz0QjONLbuLJ5gyN/JScBsoSFANk9xRy0hr+BtS9sdCAOHiQIaVq7hjz
2h8qdW90WL2kHF7tRCRNZSi2B2mSIgWJuTi3bvVw+uu7jz5QdZCOvckRA9+tDzsJ
S9f2/lzG09OHGG0sHUFKrt0tB952C/eMef82XXNiuAz1A4GmTz8QhvOmB5jJVw94
x/BHGUy2Q3GiycIkRSlZyyo6x7NKn3/bXsk9CxUiSz+JqH5zitxmDhS8pFJU2+fa
cXn2NHN8GDyim/K4+50lY516tPVCDqx6fOqoJapSQsryGHv9D8d0CI1u0UQqgNJi
xYAO2UfgEPfDg41Qt+HWjFT2X3fXE/f+5VGb0Ccf+52BcQ+tg3lGqonZhekHjWke
v+LmDwhNSsuh9JrwbnMu/tIdcRd0UL6BXwqocZ4vFUODj/Y7UQmgc85SmkD8PP8G
9Y4PC71rsIkE65AEpSYDKF4wa/kwwP7VnPzWUEjdBYRZn/uOSD91fSqjPIC/y70c
3HBzu+5zPIC+3wTJt/BIvcwSxWoCv84HAu//+Z5Iu0j6aWeqXDXhIUQYhxYNFTDH
s2doCFrdT1fs+5LmSiruONqVd/w8Z7DU0HxeOqK3XrfcaLq6yCugcsAAL0Nvm9L4
WX2BgDhsRsfs3AI4Cp1eqxt1DNMg7rMFixbaPxGsOkF9MxLCEzXaKMEyv3teImRj
Cs3dvWKRVEPurtRQZ4QnOGiXwIfNVJE6idkLutoKXKt4IC98UGLXw9qY9vbhMGS6
dpZQ70FxeBHKpxVNl9T6J/kSI2JCUBOGkmSbAhZd6uWeYN21Y0Sny63FLsf/ZR/+
hunWvb3IFfJ/eQPbL1G42yFz1fhdX4UoPzr93r6y7Ee4FguRxjgQ3IZFGjXDQ6vs
j/pINwhp31IGiprfobtH+KNy3CZylnb29An159PlXDDIqA5aXNySPZMXfODoiXVD
gW9OUiOD0qngf3NJ2YLofzUnVJK+DsNcWjw/Xibu6hAjhhdM6kuSclNRJ5H08A7+
prPgBS/40aFaJlp/BLNTHzlpyUp6PTHxgEKnvfH4X/wQXbDXgdHoGOEKnUis8txp
gum5rY3rQijEliReHOLsyWL+AwqvNtVoWANbEqvGhJz2ojC7Het8Wu99VAOM6XJt
eiF45ZpGXt73HYIUFMPgi4uifmjsajahsK0/gTkQNOgotXNYQW+JggV4dbPCsKQQ
j2gNbJJfzQI1NVZoRqPudOvpCqyqI+uZxy89jo+Iz8D1L3J5N1qd/vbbNbjPlgl6
dzDP/tX20v7meB+M0MHYtufsaN6/XR3wvoPTgTeBqdFMmZZSBqunR8Vy1sXqDMRK
Ysguquz1YN/EoH2oM7kUerLNcUStwfuUHLrdPXs3UqvzWW6nCnRHRoIu+DTUwEtc
kzHvog6z32V/8OgYCrxzACCGjSAQRWsEML2BLSSJX29PtqaDBotii7tq0fSe0KKQ
afGObYoDqevckW1iP/AVvI+svoOMP3zuMd97OSX0IzlS1s/Bjy97HMmL0CACr7cd
oFT/Cft1yzmHT5HYQx+62lHMQnFNj7KaU+GOxkkCiENLrbpUkVEs013ONGDw2c1S
AMy7IWOcV7/4H6DwYxr+SX83iDZEEi6V2oiXvVGEAfF3R26AvIvN38PuM4vXR6iO
NPKYZP0RJf5FksExN1dQffFqqk4Kb7nrl4Ma4KASSoiV+w+FjedM/3xlPuRsHsA9
CRmtxsH7NFtESlzM0069jLAuhPdCCU2phifA0oVLlthIwMW76d7xV1fy50cYm+Nj
5ngeyUJ6kTEQB1EGIYqUD9TygqVUlVd4VvODQD/YdUgWNNSt6mKtBe7RfFV8ZEob
YsddvmJSbUGuYc6p4SWUMknm+PuvRT7D7EP3i5hkgFYdpxf1gbllnS1m7Ou4aod4
ej8kcmE79g9Ujh+WcpFiBDkumOYwbaehFg0jRGk5kvtDYbHt4f4u8bE4BaEULbNK
plJ3mvS2EbWtFB8qJuxjjCicuyK5pcLrM2T7e2ACzMOHMwHq0BMhf0DkKgy4GEL/
sS8zwZyZTSaKPYwfjwiurylDTPHZ7OFBtQmo4UIP/XtYTyIIs0EEFPJyfyxTKWl9
Nq5ET3/leWZaPSS6pvSCM67TQ5io9BWq67aZYY8t4FObJrS9wYdKHd8+hlYM4Jdv
in5ONelQLGyM/eSi77Jy0MA/YLu5W+n9RRGTaJWfjSiWdNRw/JeW6LRYQHSgF7ZY
tzBd5cIOLs25yp+DVqIo0JnBw5OsGYJ3pVqqAM2v9zo8311f3CykrDiqbkvbhnG+
Xre+qYm2oAyEyEjj6bVqaR+Mqk/wNN0Swx73+UFM2Z2LZINUMp0f8k5AqQc7oUxr
JZmet19AIyKXC4/8x/78MggRq8AP28/4WZZFoHzUE9mFV6fovKaq/2xA6hDNANl3
K0jFLXZuethjA9A0IbcUXGP1v9e2Y+nm4d6104T48U/q7s7Qn78HgcD08Et/63hc
azlVpr13472ktQDWGhEjrw+GMf1oMY0614HU2AsoJ+IiBtoWjvZr5zJSOEwbuSK/
iG+yOoqkcxogNGd9NIakDikE3nrZpoOk7lqB5/WQyGutkp9lfOv7BxUyzO4KC7KS
TvI+kaxaAJKlsdvmQzdLuFx8/r5HkR3jvVj1rePiM2OOJkzvtbhJF80gWk607Ghj
edfpIHxcFlHbvgah2Qb8somxyKglYqPFQjzg0uiLl6JdNj1kE49LhDZS0OFm+Blf
GJGu5qi3CYTDoybmaPCz7oEkNiGo47BSAxumlkJ+8abnS60aM/LgyLGBLIFPps6L
Lu/ho0Xr7GcIX1RRmRiYNk2DNcrnu+YxaCJaTQkc2f4HtwBPwjfPImNTJIxz7+5h
dqU7BWK+S5LDhxQv67TPlEkpLPrbDFjCQCbUChkO0VL+x4SRVb6BuLHudkgK88av
SBMz8tWMqmVS58qvnkPlyyJES8c/ZlJYB2+7rjy6cLD3rALujqUeSZuz0T6QYxBs
KTVaV6agS8avO4KX0S19WUV4kQ2Y5JW4Fwu/2tryar+DbfTt3STE6Spw3WBN+8vy
1tVM9+UEttRWu5cuCMkZEYDMjz3bgGg0OeEQtAsb6NH70ML85CDoXhfybF2lxPhg
f/nHCoeh/RibIgO+vH7uIljS3qWCvrJ8xqZKHBMEBmtWLdkf4uIfOQQnvSgWpSQ+
RHEBsxjFkQGwcdltYOS0E19aTgnG5SXxEeliPlZkMg6uQ1Rpl+/ZzbBP/k0eQJKE
vtlSV9ous8wuOqYaRXTS3rLHOW0Uxcd+RkWuuKm4zx33kdfGu4uhdnm/ses68LBf
PjYTYLOfB+g31Bo/gJdgUztvTwb2OufADtOb8XGve2bOcw3vigckg+cQnERVuLRh
NoPzwY6WO4mo7AxqHjt38Wu7uLYnTknk8zdcVpaLBZz14qBZ2f14nwsgjNuE1nOs
ekDnKHV5wdn5PPyel1FnF0NSiUImzQGrp3+fa19g9v75XObH7G5gAfMiOSdW+hW0
LAKnCAHcPNEViiqv6D6b795poRP3MbvK6/xHsPYU8p12Yr1cPk3zsdd1ARKDwSHZ
05sqXYTwHPeGuJ951eJwbLhzItHIR/kw0AK+pJQ2WfFQj0NFbzw6l8z/fPULxOgP
GCYgE6Lqc8BWWR4lGWw0PiQWmNd/Mn3QXTlzMf79937XsH8BhRjVxiWSJ5VCQBnd
u6I4P65gSo9hD+FVELz7d3QrjF8v+300Mdv4axSLSzRKa5c6iDJpJAelAy5vwAz5
8xM1+y9mRZPlJC9PhLet2CSDhcPO8bCl1Jy4w9MQw6sHl/88QA4Sejn/ZUzINOkS
QwCYjssK455mgHEO2LRwYrO90fkDwX7e5CLgOm8weNx91uqoNCx8B0I7YjMJ1Ky+
1dM0TCyIby+sXp5OdbXKO+VMbNYwnx6P0ucumI0zHgCd9NNbPln9Qvk8ZxCotqdv
lJWyVwGJwBOIIgCfHI8tO7UHCwZpyWQSTi3RSr3XEtSjYmdxRvstHvgXvxUoH7nU
hz123azyHFMJ25iPVLhLYto9EWLLIqPFaW4bJYoWOa3ep5qtUywaplzPdQcJ3R5J
mVVNU8uPSrM4Dpoxx6+VWcYgUDUimF3lUYv1YmiMmtvyezzoryZNh4YiiFdpaqwd
nwnhozyIFZSbV8WyON1g1/2PAqJ7lUBRCwRKkPem8nhlbHSt1WJLk4q54Ovi8XJb
NoVV2V/CxohPaALC4CWgXFmJzaSthDb6ZNNE1PPYSccRtveIbuNndNgf8+QLQ7Tw
ojRN+rR/UMBblXkBaUdXEFfKjknWIKLmCVzgO+1rZg3Mixx/aspqfxG6Anjli2O3
QHd1cQkKNzZ5k/dIyHl1xLAVfLuENF5fYd0Df0qYXYJWaPiffvTb/wiCDcVj23oC
EVtHx5cgUrcp54VbhPBKdnBgndPXapUUzrkrhtOLIdW3oIr7KFc4zxegtGPxwkVc
LakOg819y3wzn8gb/kWOK0RU9cOyIIBpYqBRmdpQBjsYRVqr1EwIj58PgE1hVusX
V9fTSkWCq+6eEQRfsNnFPyUdzymG8xuT5sxAcnhsrnSnrO21TwhM9FRHY/OsZcve
+TLIPTO0bZZJQlaaZe0p+WDlC4pr2A2B9Cd1jcz/YHMah4f6IldxvGFRTFN4VSTe
gh+FlNicTYHLSqezKviMGH7Xnr2k1P2T/GA8vSehF7WWUGZOEVqparjCcHd9L15e
HiALb3fm4HKlgQOCNbZWYns+3+wtk+ojQ98E9TJ0sLacawTx+0Mnw4xJNEq1Uk1+
y9aBNl9FLJTa7goRB3inYlQjfNjHhTJjrxaclY6y2KBVre6+BSFCeu4V1W3111GE
hBR0i/+R1oldPDmngVzfIkN7+7DMUD28I/teArKcazjr0HWdNG5ZnHyrLPL6Vx99
Lh+zY2E8cD44OLlni4IXE/yu2NwVUtKG7wuROe0PW4gkF+6LCF7Cg5exg7nQfssh
SGoD2xLeanVGSyCgL4Ma20s3YRuYGTju0Hu5xabCllrRsWkPgd0c6HHrLUh22OjK
4HiTpuzwIiVdcqpGglC2gp1WMKWja5sqfjrsQjoZf7vexf+yt/TgY+9XSzc3amn4
rjrSyrtpa69am/M3+2e8VMIfsLR4T4aS4XZf9bKScIN1SWEJI6vizqixVbQ/yYUc
lsx5rfyC6JeRzxcfPU8tIXDKHX04auI7eIQqeRCTCXHUcmFFR0Hum0stC+m/GiEx
2N555wIw6vWLAkLFUPq4GtKTt9Bg4UHoETM93y18heFIFsK5tu4uJrmimdMV0/qE
JNWBI/pVK8byT2DgLcej1KIXMpI+Uk6J96XK6Mke0jaokhIgl06DaNKxKKuJba62
BSf44As3cvwoPGy51tbnxPfIewaGXkwBTqtC9gYvSACkY9y2Y4hhfoMFmEaXu9M/
I3l6zLAv95OukejHJQn09mK7ST1yV3x50GPSugw4Wb9+GAsQFvIGgNFVBvqyC0av
DZyAWM55bbeVFogt13qoGu5fp+B5/C+M7qCG+0rwVLQSaZZE0+07CNwNlg4hjBTB
CV6wOVVwRRTFGel/yA4WNACmoWHHdQIUNRqeDVorUh44lTbp3GMKAqJX47OQCZqx
IP6LY5jvryLIgtoIUIRnuYvJGGkVg+nqNK/h09rObLmbN6+K6BMWosPp+Nl3ABnH
5qkDUlIR9V0l2uaSplCO5+e649nPbmiwZveCmR1CTYN19NeLnsYQevEiDAVOhcsk
+7fgyBLtmQElD4KDKsnZ3drdEr98E/kzlnOFJFEcLidzrEHiPmxkt3lFOZ7w6IeW
6KbcIu/x595Wbi8+faTJJ+rime0OQlxl0WvsswhyrLfirVEfcpUh6gCESb9l1sa5
FyZyHWUsSOcExi09c0YM6qExz5Rcn/IEDxCoHEQjNGusaPgSFd0O5r4hAhzR/Jtp
WyT6haK3axkcy79AiSz0I7FlSizfMKpKeqLmpwrEdyO1vqmHkvr+SacaH1dVBfkQ
kAoanOm+fsluYGCPryWtp1cFyL9t8TMpUo81ct3a5QEXGnHvFDc8wkAQiSLqbDwv
kJpr4+8fz2thX1XfnccLu/P5bp0hF0e2UhWBy+47dY60TkI5efq3ziaRdvNGKIrF
+VDD2S+pBT3g+HJOcowoXr6vx2rLfrkzxJAQQPmoW6RiGVievE55r0qV/iCA+nyc
3mB0IH/XB5OchLMvBJMglmIYHRhDFs09lDZW/w/6mCTuYOTbNzFawsrPYgdhEZ2a
mQPKmUaqkgQiHUyDXImKhPTX/htbjOOPyxi0+Sp2pAWANRW2t+4bVf/6ywGX7n3X
fG4u9CjvB/5F1UOt0/S3RcqI/xOwSWtt0LuoqDhfYYBebljESaFN1kbzazvTXlpx
5+vXazwAOWzFoFDlEV17rAUevQ0ACt5sKVFzuuwn/S2D6AYiLhi3ywf1ttXE22BF
hzfWEi5xPuslxVZ/78151tLVKs3AvShTlyEb9TVxO6r31NYRn+n5OXE6d0XiDoX5
Rhhh8oy7Ooj+IBI7EbM9LIKtP3BxhQPoDQ0ZrmhsOPb86iAVhU4K5M4T7UGAK7B7
ZwWptSlfnRshCkCJq4EgsQ/Ymck4QRyrV4CYeJ8vnF38fBJXdKWPeBbJzlef0GxW
90+MB4yg6WhJl8ec2fnbvTdrksEAypiIBoKXB4jK+jlyYneiEdEW14KJiEy7FbGT
1vUhri6pc3GuvKK020QVTEz9LhFwyCRU1ouPK/2qPMpI82iBWy0m16DmckB2cS2m
q3tsrQavIbcyiBKv8XU8m1iFncO8yehUfr7/Fjv591vzrD4lFyo6qb23U6jd8qjo
q5Uej/1qr3zdxdTN9pQwapUar+AxCGCo2TAzPxaoDNUSSQRoNSqAdK/IhlnEmGfl
mYI9j2x4DVfTiC+/rNbvqyiXVymmwdbQSQJy0u2P3o642mSnyT4OMxFrod2/PEXe
iRef5FqA4fzG9hppZhpgPCiZouRceuEoPZCxJaf+/psLSxGzaDLPOKgnaTyT8QGh
9Eob6ITCMCHz4RuRYuDmF/dSFyngbuVu8C98/ElgeZLbtUXj3RCVWkG9z9omAusC
0EarOr+smUyS9w9HzoAFud5ygC58i2yPVWLggZV+Lyat2AkL3oTShyR/VD71Bjs4
XbrWnB1mCZfiSSz+Ykh2phNTvXAMS2rI3URA7bw6h05THd9gVN2dpzrwu5K0q12J
7PywCBs66fD0eyMaqJGWVAl/d0MQpb4pAHox85+WXEApvNH1SUP+dZwExUn6arn0
JnWySmItUUCc+V99hBL1rquJoyv7ddY9KrDTMInQVT6k3PErU+M3+1IcR4DpwCCz
kPto4KqymJ0eI8uiNZkUczozq9f7jJDCM1VyoUB8mg0ox3bGW/6s0RcMfYxXiabj
L8CKPnaTDYGcwxIyc5zQ6SgdcdXNlAintWzJV9qdSI1C3/6JxHgdReAQ+w6tHEmg
s+mvROOs7vwEEa4caFcG7sd34qeJyj5a2QirjBlAQ5MFgP17St8IZ+GOPrh8iZRy
tcRpWcr1lP9Yq+yfwkqVHg+QTyo/0or69sXVw07MFfwkKKI9MNsrCyypIUH3t+Gn
nw68uMbPdLTeww0Mq+WqDD+AzfkrGywy35BJkwWu7AkmkcR2SvneRscjASagyKjp
CGG/3dwmzHR898rYxBiDkjF46DT8xbJZVXkQ7B9DYqP8sqR4eMjGl6Aya0RYPTax
2n//1M8ftaivpAsp/JItY8EPQ1fo9xZtBM6ceMPLNLtNW2dgbT9qQVi+Dh/j2pty
SaJCpGxohPSDvVnTYqco1HmiegJZon4f1TCQnTt1lYpFZwIspK+cfUKIJIm25dyq
uki/TgWYCLsiZUhH2BK7B07LbbE61BHyYVoxpvq235eIF69CUf8Lj6qE/mRp2Pcp
xcrwv2xNSkRtFK7scKVSfl4wgy2ZL5iyx5U+RYDq7JGk18Tqf+BrCxI9xuMhY8GM
8vZwY2drPVkdYcsjgwPNmSs7F98C1IYqQ2FtHUmkN3AhyDWtWCDl/h7JTtA3+X0w
A2mIgJYlAhWJyBiCR8hPPEFGo6AzVlOgAqlnddXsHcRdz7fQEBU3euf3TiV2iouH
1YpO89DzzYVDuaQlqFhBgx+lzo4QDUTON8yQVRiopNmEAXDGbdb5LRDN10g06uDA
c1agdc1bp5SOwoFwUK9Jcc9+/Xivs8ZXcKb/MCobD6HD1KAwgotyrfc42HBJXUJu
/An9XKGiGbYaHXOJ2b/5p4Uut56sUS5PlNf/El84FcQp/LcKn3DJ07waq6l9886g
c6pjnsmSVKZ+52/0meOz/6r6M88RvR3LLmdJkvmQuDKk+GhsBEC7GufufAYZe9SI
LG9HhbkW08yWgqweoTylToCQa1n5PXBKJx1IkvCiAwtSNM23Wt4gEDnVE2ZhUiXE
xYWjDU7LKaq85Swsu/vxj4hjw1LQrnk8JJ5WexOXfaMhY56qXwx5wDnkYFTL7SAi
QaxXUj49cJj9Jl0RBJH0r2MmQuWffhHzvEmupHbxb5/ddI1XqU0BoMC0xahcWueG
BmRRkl45sEBI/Ndtil4O7bsTLjA78IY9EhmoAMYS5BARMxsYEN5dqd9akDgWC8tR
kHwB4luBOWouFFlG9tVuu5LYwkrTVM2QXVlI2IZEGS7jxhTCZCTUkoyrWdbnmv3t
7fcXFxkX6s8eAJto2Atgg6C1WOjFmTM/gk9OTTVmBXLfLFACWG2wCHL3QwKHSZHH
oyoGHHkxsn51IEAxm6fN2Vn3GPPVRibq8XKoVhg147yGEEaHbr1XxmD15VxmQwPV
c9wAUAA+1k7vL8kTam2Nq8UD8/15YXE7MneQcBMvPwu9hbO51kJaZoSMCgP9vnQq
HUxhs/irPAkRBaeqAiqvfBdrrYQ7DcW/a/iT1HOhk0nDno3Ry0ZAHVlH4fXr8pVg
s875lZpLmR/OWHxQnY3PmYIpLnTBWvCmlvpgdgDH1GMyP3Kq6olI5+3qzFR9Nt/W
sF3lo93YtTmCcdPv0s8E55GGnFpKkFtP9x9l0tnnHsN7uG9tvPdIy+v/hgU7xIZJ
kAAHz718TI/klzz47PHvi3iBQmzUZe7li3Z05Kw2TpW0hk3gjfFpqmLljoSpMbGe
sP55VrCoVHxtNbaUexOedRMrUtejZ3zt0ZVT/IEckmReMeHThh0y1WLIOunEDod1
8YPgXh7oyqEQsriYDaZ1aozyCANR7kLj7Woirw+1l8zHK9MU8JZCZQqmbGWvF8Gx
ZYNXz/WSK+Dws1/44BxErRvGe89C25RDvf6vXea+iuVdZrwiJtIPwLYmrQXC+bTr
EGuAGZV0liaoP8wT624uv61r6saj9MraKuqeN4SVl6VayNGK87Y1I4t0dC+PjnhZ
WL94KvM5rFxzpCcaGbeLrBKSHCfyKSQ9FhCtWvX59M4qkMtLjX5wyeErjcySYzNn
SDMuIAuCpLwPZ1YZ6llL7ghPfyvxaFTphPGnmDmhSRF45W90yljEoSO9R4E1QEOa
CRR7wGgymLUYLMEB4Dmu6Noo1u2NVOh+kL0My5QmbFi93Inm2EfiLULvR33qFy8F
3Lfc3VkFVTn4QMAns/HPlw2gfbud3kMTbQSHogNqQvL577UFKXZLoqdO3ThPV2Dc
PjZUhBN7jwznnXPLGov/VMYzrpVhz5LnLzParAls96SpI6hjPLlnUpSzrz7+aa47
NBLpUdFNQ3GGphgVjq+3Z2RhDoSDgieqnZQO6hfuyAlFqNx8Yqm4zydpjBL+3xN+
ny63BIt5kRfMJEBu9Q/Jkt4lFuh5nb4NBsk9MMzAZekpPtC45+NbiBKnViXcbE+J
x6hrRfKmaJW5ZKaYxq/rH8Y/aFjrzTjAEa4AQkYeCGj7F4lldByyu1gDKI/nq8QH
aJQFBl+wcnHwi28bhmsaz+RMQbKHfLOWROWpu8LwgGNxD5s7jySqMZyNVdTwYQ6z
x3WPu8M2GezXscrM8rbSyD3DzHEwvKVMfPZGvt8uU7pgcIUuLCxHt5kInnX07Lt8
U/ELwpeyEAyxkCeVJG1a71ipOS6HOpZdcogtumeK6FXFYaevkMNwi76RCC/1cDmU
lRXFIhcx/oaomIFDkar9VnJTVSPlTdzLxHLAysTOtipolL0FGivKxy3RMko4CcEu
tcJeOBUIy96QXzHVmuIP5oFg3eeroUrJ8rg7ZklTakWISjKrP82R77sR9AGdgcEC
p+xXJBhOutZfEtr5LShgDA0zm8q9LRcvesNFl+w9aUbZTYHsLFkDEZnPE6JDxjkY
mbJJd9/22a541wd9gcAkJsVT9Fne0bgQfdJlh5h6vSGT0KhF9FSQuCZhZX5nJDGe
6CrZKry7G22yfIoqAJst41DN0FO5pZiLF2mRvLq+glaqgGjQkAKAr/CMC/08UEDW
wpzZ9Kc2FlNyppSUeoMD/oPvskOMFuesTz1SNMif5vuDfSdwmboujpuo+iSt9Ngc
A6oT1aiWf7mEcN0Cao7D0SfqVKnWB4ETZO1OkiWfR+ElNNtBvSFe5hFwMpoSdpAu
ZVRby+G5sx3b6rOBgAHc/sibKdXjWr0Y3bksquzKEBPr7WGXD0tKti/Jbn1Kv2sU
ZacHoOAIQLtEjrXd2+MOsNTEVCYb7gtpxoLxNkVn/YD12jCg0MjcIj+MhvZNQqgC
XrhxvLLjiNrxU8RDmoZn/tLeKPOKZB0XJGgwmhIojMnZoXbQW5qlKd80T8sdRZMJ
UUzGKwmAiwubNwe++Zlvn9A6EEiyWFyMcgwU8rLzXE5AvjzMz09SjokMnHqwCKHY
BA2F7JAWKK097qtONfp2Hvp8A2FYw3R2XVfzIK07wnfvs7yUvLgwpqOpiEfJBUdS
RxkzFlL6fItWTnpYV1E+bIeQxTx7yV0xWVkrk86A8LE/zB97QXY5jPa7no7jYyMV
MEMiRlizSrZA0nb36EBebOg1nJ1iknJAb+10bmlr1se7YjNKzIPUyYw/Qs3EfwYV
q50v8jk9/NjEti2VDTONqBSA37j295FIPz5YvUgWjHwFlYjAvOLPX8zO5zgFbd37
uCL9h1G9WwawvW7wKPIHJGKEqJXoE1UzlOSvL+BTfEyuq3hhDMXfpJAIz6xXLY3j
TLrvW/EwwDXbyi3C82pWmagvHtguzLF9Yn4OTWX4aqA27IJKFACSW3MP5e4nkurf
pDZbAZb82atxtCR3fMr7K2s6Boo/fNfAhSjlQIuy89t5ytLviHYHh7QolXjTjvGt
M+2U0rbj4mZCZU6shKNbYGIeXj9YOXocs8a3DTw2Qnh2Hom3aLtHa68CROWwBZZz
jfCdZvmxqvrhazVy1JKM+Yt9qKsbjTFgiQazAtEVaH2qprL5oXrDPAv6doeIPnxW
CiXWWBJFPV2KhryImnYNobuSIgeTEfRk+luuY62opPohcv/td3u6h4daAu7gSI11
CHPqOadUqRzYtqEZOzNVfmoOiwNfx8rG2wdFc2VYT/Wmwt2XoHdQedEK6LktCWQ5
cSkaYlPpfpcGgkduowo1LsDhAEbFJmd8enBbqAGq9KGhvYwKtzHuykCaljl9SNvc
nGwWNMiFnLlEH+FUbr9sSLBqB0OwWU+9Xu6F/RJRqR90bMOec+XhZ2BZ5nHH8Nn/
03ohN8uwKsxgiUFlwa++1oQSYiVxM365iBjZ3K+JCUOsapNX1nbH5u7vQ52kQwQS
0C75YhXc/79Kb4inJUq29TUCqXUhvBHw44LTYOO+XHHRnRL4ZaL4wAkDhV6EyALt
lL6NXK5lzZjVxHNi29lfzSnCiJrZOFfxCsScmj6755OGLuztPPI8SvUZEYixYDpo
mSV8HbAUwd6CIRRIrD5JPnw+UF9yi47ojRR82awUe8AeoKKshPaq1l5dpcwa5XJD
M0JGMSa/0aEnUn4OBIm9vM14TYwy+cELG0KGxk2G+5Dc60gskMQOCD/QfudgM7pF
/VhBtDdXXhg8elCFe796K+8D6S0UrNrmxWL13L2wCd5NEGfETvJijIhVevIzuxJb
DnaC7NuPTJ/D69Zi8t/PQW2/ax5pV9NICJcoerQb8wEgAqK8VTYPiFqsR7ujbai0
qKTKz/fHd/Ork0EXMtXkF8vPsiJv8ZKo4WPxuReIk2vIcm16Ym6Xmj2UZ8T1juJs
upQ41Z9loeXtgv7I3imyWyrPm5oH7KtRpW6iFuRfyWyb1wyU4XB4OZmbqDDLsUJD
XkwZatw8zztuurlRAorBS5BFAwI9KWqqj84HM6SJYqoxhZ0Vuxayg6NTaWga8qPV
h3zECRd1HVXgOMcUZSFCtYfVR/qG4OzqklsqMtikNz3N9SosVtxTqnBH4t5RxYFX
f5kfGLucmRMcNGM6+jo8NDUIW2ouvcIv08eqYR7HuDbkT19p2dBuP3c3fi50dOOp
fDtc/T82hf1FuDReCYnm5r7q/luxvi1TeJ/sziL+oDSAFtdw9LgORQFMCBrDLYZF
c1ZiPp0SQJU9LeF4IM67L4/4wQIPk/cnprJ1KV+8/NeymSnYg02oVKjUc5Qw6c0c
mLOIwb2s8uxDDiFTSpD2DgyQebMQigRDZyK4g+YW1N+te9DKXYRWlnjYhm+q57rD
bdnz8SN6TMqbdBJxKqacfjY0WIvbYdMW02uibYz2NkZjM0kfJOdnE7ZoIqlmwrDM
Rt8OlzgC9CbvqSgfEsRx+k3ty5SJEyWqi/sbKeXxjxnV6LAektFGJg/IQzc1MHmf
kXlGqn3ckgWFKpoi6euv8OSe8jW3cMs1X/ihYUwy1kY3agZsD4afRwo3gqTyf0XN
L4ayHmExreZO++LP3ym52IHrmcDvPQG7ejCMo6sRqXCd5So8usiJSon6t6M2lDRU
eiAnsN1k0Nz5i6fX9wsuG1UPH88E2o45IJNE5HfagPkoGnDmaa+YZm4KAjxmNir5
dZZ9+bfTFTn4WipdA9KxN73IIDUks4Zou/45EBFPpvG674F2j2nT+6TEyIdXHFEh
QK7SuOayOiYvdTEo616Q6f8xjMlWsfcYBhNLUezVNxEOMBdU651iFueq54a8NyrP
Pn/gg1tvsVW9bDqhdvvdVwHEedb5SAObqCoqyWoDQDZCfWzBAA/EyyKx/lUNa2Cf
KWFlODJFw7+upAInB3yx9iEYMA24Qn0w9weSap/PBXi3gCp7GNACw1gOJY4bXay4
w0OJmpYZopXHi8mpNT57COfg6BRdSPA7FqgrF1RhQCcIxjaITULbunzA5ZbJT+VE
MU+cx87qKN+ocRJk1snUOqaLmursv9W2ughMmJKCRPcpm2zh3D+juPoTy6SDl2cu
IKn8saIMUyEx/Fc5pvHFC20ljBlreq9LtpVxV5BtbduhAZGFXJIE9mh2DnAXjnyT
HF6n+ZTK0f11QqktKI2qrUl4GKhdq8eGCBRF2EEDtz/gS+An6rBUmz4oJJ4xc+7t
7lZVxQt7bfEszIUjU/muFNkUuCXgVFa1nFx/5Z9+Nc/HWQTKfB+CC+moPEsJHEZg
Z2v1LRtDuRdZda6y3+hIR+CyvDEcICyVz27izHaR7wDLvqy6GNX0STghq2jVycva
EmkGVTouhwUv/ST77lGW4OgjjOgRakqFZYad9L15GhnxEonTks7LUsZ4hsp8WS4T
l759EpBjShlc1UTQeJM6oV8JDZY3vhsrOgRKIQlNbZHFEnV79MmWjKkYq7KHtFCb
y53D0/G89wrwI0LCpmCUMcm6B21M2QAq7hl88rulBEzdXU+JVXMeqPAL0pGjJ0Tj
27vhSo8euMOHlNGywtGH3X0tsho6q4QznJeu0A//GpH4+dB3EPfP42y6Qx+7F9rn
T/84EKrAbKGUsstuiqvGs+naWow9TvoowWBuQp4bJQg3QuhGiHSx7amhEPYpGA/e
kT2qlaKRLG7mP5KGiDBLgiHZpi2r2nFqME0tkhAfroqIXMbFLv8gznapV8hGrf86
k+Dfy5MniTaOtk0Cw8mL/NgIBRgHpUyKwMHM3slSVTnIPVr2RbFc+LUfq4LtrGka
WgLORb3ddV732+xg+8/JcIeJ+GKfQhJKuNdmQ2LVva7J+nREfktKueilqnYXT5vK
AIK4ggsy5lmIHv8rouHaSWyeVEtoxOWyt003wWQqZfTtTFT06ndQohsRNuRz+Wwe
rj9Rk5vZ2U6XQjm+33mqQf4HFsiZCA4fVsbWrvahGsWnGp2MYSgb2I27ul3MTSfF
9kyFBRr1rzOvf/oYtNCoCh8LNzrm2+sQpRwtwvk5U0zaq6YfMju4Qt2irEzEIF6l
Gga70qvA6jPyM7+3noAzLcY/c+sEkRyrxzVnUnqhu1oeZVqWQQ/blK75VX2Q8mG1
a5SdGDZEdCQ6AXraMw34+9kMiainosIw5kAsitvzswza1EGWBw8CEF9BCNrlF+Np
NBmgMxoZ79rnVIglX3VmMjUIyq6XclX29jVJNRx0tmhwvZcYB9wTkcuYwHpilAel
OeqjUO02WFl++43p6jUCl5Jbto4JQtdXm0z9unDHE6487jhtttNN4oK0HX1Ou2qT
qt1ryCnQqto2qewgEkmofGUD51TJmNItbASTXFYvzKTOpUHKnlT5biKZ28BQc4LZ
SnMT/ZILhERLNjT7ycx+fuYSIitHxjIIQHSKn2GKY5ArVLFR9A61OswTO+Ib25R3
XQmNT9yZWdzQLWwsronQy3OeORChAxLJ6lU12nYSvWWF6/Hs++Y69d9sTeI05Fe1
2GEhZmDQpY4S60dxbW+/94TiGzjv5ZZAiKgHWp/evPKcUYQnWGdK3nupJdHbydJT
LhmPiJKD32wAxzj6m2Bap7HGRDbU+9WwIkTlg7mCrTUxLmJt/I5tMbuNHDF0yHo+
f2y6DH7GvRKRTUXsyBn2uE1P32j+OTiQ/139NZu6L/WL5qDaGOrj58BUawO/ZojS
Mp+FHmXSD6+Q2tTcJklcy0AReX0/4nCjTaHdlFCHvgvlIlgGSQH2wgQ8V9OlCA89
AN89Qi9Mju+s+yRAFO4185FO6cyL09wIZ1NAVSTrQoONJ5Pr//sQyUiVTVb5JdQl
aBB1lgdK6+wUjvvwd5JL5KpHI5B7X46kjtGThLSviqePadHEPapJGYOnoIBNi8bv
oRH6YmO9KsrHpSbslSJ7Kv3Xs6fdMjM6F7hQcQSxbpxitHgBqHnWj3sdIKuFL0hv
61seyZ3z34I+q81SxyxtkfzAGvrEpPD9LqanAMaWHvGEWfgXeNXpUszz1NjkpEAX
7OIUa9hiBMWwoslAuSENmg2XYFdPruue9rDgbbxtGwCsvS7U44HTAPZRYOU5L/iv
0MqEdpsXoWigtPeoWl2cu4IcvHNN5hPAhOvuHO70lw0cOj9gfboPr49ko3OspDWz
XkDQpSRp1Z3gVEFpCYEXzJksPBN6tO/v5nFXRehUeHZR7eFL/XkA0uM/d+wGYQJN
hKYameVz31rU7gNziWO4PKvRCjZhK5pXUgaWUNQO/Cw6nuaHRWlc3tiOJBD74pCH
IKlGF68orsLBpi1A9LqmMLkzMKgZvGxy3z2NF1T3aJZkL9UJhjL5DtZvf/bNQOu4
uqFDnlHiP2t2/aEYL88bRlizEG0PkRJ08XVQtZVfClmED9dAs7wrSN5Ptn6M20q+
aQ9ttQdKtZ3MaUAktoQQt+UFh5SDRN07+5f8qkIETCiSQcDK6v9woxES7H0aA3Dn
FCCcKvk5eSLq+G1WVYZmFiZpTNvpatJ6WTwHRL84lbBYje5plc7obX3QEnezZ8UD
1KsCkuw47qh6Nz+7zZ1ihetWaZXKA7endmc/VlseGBCtPmdd2zXLG62cMyyWUl2Q
fHc4ywJzkFL103N+4r8IoxlOhK5Hm/znUomiIsD5Byf5mMK702P9IhimoJ0mhNGc
EjHVZQ4MwFjetq2GTh9+tLQ5soc+WR7YMVrnkOamxv4O1yZ7x0H25rDqFht2txFp
5zq15WMW39NGgPnAuTf5UKr5ZvRwwQqM/nTK2Zdu4gYYjDOax46xDpPPPAAl6KsX
4IDVxksjGsGlgzAhFNCookQx02Fu5tazHjr8TKV3K8NFEED+w9WtwBQHFDPKldqK
3QM4S7C+kz4DHjtAFemyoj26RlFhB7UASP/RhcAnuByGjzI2TD+j1JDX14z/g7UK
zkxEj7XJ9J0oV8Whyv3jOyks9pSqnkLbKkKFQVsWk24lxO2OzZwvRRyrAnVs5Nne
3bbcdB2w5hq0UWcb/5IYRm+/9kWM8zK9YEtwDrGPEZvjPCbWLZmZ0AYWxdQTujgF
lEejaRA39JhrGz9hi9vS4BJ+5Db/j5y5XzYY5b3V9XIT9IhJlhUUg/UeDPDbrsnt
6o4ldNVJy6x6AerbZV62ZfvCGher7iymweH9UeQGTSA0hs+qQ2sfh0M4rs8Chn3w
6669DQSWwOpFSixDKGn+jbnpmHHzGTbaufJhOZ4z/1oiE/4oVDzHUPQDgd3M0qag
l2j+r60CeMmvCwr7iFk9kLH7fBw5PSUEjP0QLs1Ly/mY8PZfJx90PcDcO9T3fV0u
iP9a0zvxPo9qeFg9ZP2nxcen2/6nQfke4MGRvqd/MzB8HNxBwLq0WZx3e0/goINS
QP5sBRp5whQfxCWH28OGVDV1kz4LzT1IUD2gOgVjz4Rj+fLqh1AnK3HGU9VUBfUE
4AmJ2bi4KDbPyS0e4cRVZuqzkGgX0hnji6amQwSB0XbeTrfIvyRUTS9f2J55CzoZ
95rUNssbqjsJcOn9uafmJEpWKsk5wqg9RIfsfvjlrq6w/AEs8zJ3QsBtMn7uVYof
dtCFr7Pc6Riqp94JUlIrV28DlpJs2j6RXx5qihp2yfKjo8VWDEXBAhKbaicPTwum
KswuhTQEFP0tcQ5Hy3eVgTQWrZ+uzACxI51nEEGrnJB29IixMh4ZxYm3GXlEaqna
2jzcdQ5jju6IdjE1gtXlcMnNI7szKhZ7nZKkdai/g4TvZvaL9h+a/SCGGVgXv7id
jDY7br+qWjd0Rzcx+qwZMtomgtHZqYLElaj+BsNt6Fmg1ve5htrmlugtvSjEg0MT
EtM2hFPiFktVLrdJql+qKsECOZ1DGTHH5QwCmakPz/OoiXT6wuvKyCjEocezBWgL
ONt/8ubPyaQt3e9yNf/2tmyuWY3wbMisKMpK3rhzWiqyS7fzjpHOoLlo8P/EwA8z
lK2VdGIUO52uBbZwkVZ1cykYLXci70bYb0rFrYqWciuT5vgM3JRK0wjYMzb7PRPc
qQNizjdaoXSsCmItCWiGvBWIozvhWFnd2rrOIkNLRFmLMlfxy/F0RAk1M98KhDCD
o7rP7Jt9sjRPLJJTps1tkFNNXBgMpV/uCa2kPbfNumCsGpGs+9sUxcDMkWKiTFKO
FKpqhotQSMaVydQbI33VX82XFkmcuVYWCJmzAF6yXXj6hBYqyvzV3/CDSkY64ODb
mVRo6hRnQXBKVOeGpI1wX+1enocS4bUOm208+iqrlTRI7RcByWwBZA8lT2KZCYHT
wgmtbla/f6fkIRhbT/rK6/5AeFDb8IRxJZgR9TKpmlgt2ZIHiG602FwGtv8ieWfm
JkToX1ubssFWMreza9OuB4vh4BvrhT0cuGpPdYDENn0=
`protect END_PROTECTED
