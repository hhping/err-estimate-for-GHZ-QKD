`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
df0wyQ5GlfjJFvo2cvaiHjuobjr7vutmKyEP5IBFeZwDSSBB1MP5DPa1GdJdRAxk
50ENZGwdBj7etgcYLopxWj8UBj6Ij/sCZjUlcmFQJFujpY3vwZEchqbgsbzqtt+X
9hQw5w41927GATW6DLkBBTw/mSOWZh3BSZIvToGHw0pQyQp4NvyGnaBzruIfg3ZE
3A6Zq2ROeg5PgifepxIxvNQH/+LbBSOj54W7YFw7xnOLNycZoR3/pZjZ+dZHUm/t
sCW4G/fZIgzCH+2reZk/Rf0MQFqpYaDg9hyeLQhcYdml2jIk2d8crXetz+NTzUbC
M48Lh5tvS06ZpBkbIuPgTZw5ztge8HYxe3MH6/Ksd2UV66ELKPp0FgZTKf/N15Tf
GyOZu8PNlunLtfaj5GdqFtkmCMVgVAa0AWCOkh/89RAQu4XJPuythR58mIZoEaoZ
AjSwnilONIKh/GItfDhAGwavy7ep2+fmDOUEfuqiQpEfiqFuL2vFJbZoUUqltBkm
IrnkE8b8HvisleJ+97SnYg==
`protect END_PROTECTED
