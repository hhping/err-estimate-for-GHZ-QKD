`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqY79KsFCLEI1bEHsNqRJkkbXXYXAWZs1U27vk9jZghEvl9xgLnhyj3E2yYDxbtl
DZtyBjUrPDg0rPYtnmxBPlGQE8jC/ezI4PNvrQwj3u3qE+Xq/BG+9REWLg8VMkWk
niR8TE8nOIjfqc+qdp8U+If6xjirfIqoBZhTYFZ8QwlspXIdyjs9cZHS7rRuYw6m
zC6n9mf2XLUIkQc+8OjNeO3zsiQh6qFyVtf3n8fHw1Ksy3+EQ2m2nilVThTXECXJ
US8VNAkZq3Iqao0BBKzvkIgOddTNcQjZE3vMPLGMcqTdR9s4Q0dZeWVxwxYlGvZ4
wTJr9YCeERPSs6/F8zbTHAhOLcGScLFLXeUEcG9Hl0BkUl5eUivdPHKq89/KQtvm
RvvrfC3TD5+AcjCR+WczhgUQEzwO15YjprnuGicNh7EAni+s4dCCLgXxM7XcLgTY
bdpAyVffirxKXwbcfPVCwyyAohXG3KCVWbhbWRAGZNfL23e1Qz66zN74lZE8GZzj
Iy7WOioxUG3UjjF9NlARtGBZtiP4XNXeBC8ppCzf3cl9uaU0VanpVn582XDkW3g8
vUTjMBfLKD5nyr3Y2CCiwd8ia5hE9+1+gctglSzk8uN2AfYLP3TWraDsxaRElHwO
`protect END_PROTECTED
