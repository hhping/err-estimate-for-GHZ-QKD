`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gbd4ZRRp9jFp38ElnX9zr6vEcWRdUi/rUrLJY/sUaKPca0b5clyOSz0SfGSAxAvZ
mn+tNgMR1ulJD6eIKEp0f7XAGZvOpoWir/PocuqbeAsOb/GKdH+KjEnvM2Z+OgFR
ZtGGYA0q1G4X8qjuvT67A70WqXyaSMNCl6iwq7oco5eB+UDTg8Xm08YKzCG3GHd4
WvThYuYfL/VG6Sor6FJ2SnAhikOx8bDzyau8qflwtW7FFRMV9TKKsRr02Bs1SGNF
BDUUYORfxMtXTpaaAL8ZP403YE/MqeC4JuMKyZkf8rBdmoC9votjx5hjFPVltizS
H6bSUGYgpLgz1wQIcerY6L85R0WdI62dNBej8R6ufISUvX+aIf6zwlwKEprxSxd8
rJ/JDCIjRkZpNwqJA46ekk4O7cawIcMCM9kuRVXHdtamb4t7VC3E9MgxV/AfjcLB
jhbuCCB90y7rJv1tGMsnUyP39DCliakQaQjdiLfhpZu2Vv+AOaqxe9rHhlLuwQ4I
MRQ6u6y0l/E6DhepSo7hsquUNAv4c6aLX3xhRyWJjJZfR7dj8V6Sm0812QWYzYtn
G6GzrCK91L7MJiU3EDZ5STWAa+JuU7D/MAO/Kb2UzffyrEdbP9h9cNaTczYIS2Zd
+ZX6jIre8cwhReUfDz051VB9cGQPuM5geEmsbpmW48QSHGLICwjMWyq586SMSMiA
wvVy1g0UrXsDeXD/oBxN0G0nlxieptYcIZw9ZkZ2V0d6Ahv4l9svbcnN/+TpILsS
S8BdRnDQQF1jwOASGhAm3f/SYgvkaJxMoNcfnTvNurCFd5WZ9lNAiLtSVn8PgnMS
JIIJF0pFgH2rPXzvTw4VDkeQPGX7H3qZLZTBYzwghyzRMk/J+mWRcQ2VzB40GlR9
Pui0n1tKf5p123sImr+MVmrthEg7o9gA5AXfbXAAPc3xAQuRpAUnSq1lhJ/PT9h6
cblsdnVSzmj4pcOguPejRsnVGBJPh+YxcI4oW+fUO+xWK2EJGVA8vQNhTh128a6k
`protect END_PROTECTED
