`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogEGBU27dtBgaO33G2htMxzvLtQLBhqfeCVhbGEx/EYBVxbpVMWzLGMj4UjMoBTh
X9+zlPwdzfK4koOyFJRXomzfIOVhp4in9Z4BUyHhs6VPeFTsICRoEy/JdI2zMUy/
rYR9Ht6WVv+TaG5Z2bNk+tZtr9w5u+tfVOEsglq/c3axK+jw1/VWhViO13HmjjvP
71wBviEkBDrjGimePM9Cw6VqkjUfETWZ0FaOpn48sF4WHC20xK52i7hBCj7pLaTZ
1XaNfCV4PabuET2hYIbobIk2ceT+Ctuh6JZAyzq23bGtEHgapvd6OLa/WFUgZtUN
maHf0YJpLv2uXfsXglv9iuhFJmxqc69JcRWr6uL1e53FqxEYNx0ieqQJjy3Ht64H
39uoWucXU9kRVmRrPzsj16gSbaSKbSmTtyFdPlTpWO7FV0sDsFcn50aqJegp4Jz9
M8uLL2H7IqMMBrH4XMSZtLXGQJDDUuX6mKOYDs55p7G9aRfPVB866JlnoQm6bsA/
7xT56pykN9BEhjkcPfDVeDU+DEJb/vyuB7cKIKBJj4LvuXYI5//6Oy7dwoz7P3/m
TV4xSqu7Fh9cvwj7hA7RyZ/nzBe0H9pPAOKsUDZN38feo+E5hyb53K1evzMWuGSj
mTTijP5FNob8XP7hPkVt/TGA996aEbB+7lISLVHOKM/B/IBiQCWWzFgPS4SAhvD1
HCNBx6dlLF54BBcy4YysISdaq+V4uX9KBuCi7Jopk49I5W+wGsNO6qoAUBJ2ELHg
txQHKqzV4FGMYWy4wdIVaQflZ+ibteIbzR8x9fc/pefHOzjER9zjaIukcVG6UcrB
iUNZP42dYE/kcsGKluJ5eCk3e9kfdS/amhPXcQQehwF9/Madn6si3Ndl7GnQbg2i
dqQALGNO72ZW2pYOr0+oFpg3EL8gWN9QLAMiLil0Da9slzkRbK2ga7XUbzmv86HP
hNAHXAnZ351rhPE0J3ktOkJW3e3g6aIB/SMnv1HjpneLgNOhKEy5bplC/pyhsBoZ
ggBnpRWNdVyrOqqC1ePah8nf3awM5LAFzT4BAPzZEnc0D2lDNOiYJ0DX9QwnInYm
6jaLjibxHKLKVLz8kuNcXjbMNUgLh7gi/HQvYKR/UoGED/b9UAb8DMjNkbZzBncN
mtY3yEUhKJtGAsQpG53FxfohpTrwzIBNV/8nr2263rWCrU2QWgqWZSf1gQKvDQpw
`protect END_PROTECTED
