`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJq93xG7h4OZfBPd03pHiTZ25w/BWmnl/nRJ/BLzRlupFru8WNJkL/njwnHV3zQY
iIVYsLmAKvT6c8TCvmG/1Ig/2qiWAeUEUDOKtb0/1rptUUovy3XMF2rcojaD+v+9
CT6KFJ7KBe7YFl/wQWEGP4pjeHDTItbfE7QruedqMEOkr1fYfu/vjLhEzCLwBEFl
1+RWCO6Sl9PNFR8kWZ2AjOsM2Yhgh4ydp0Ow7XYy2QnJmWT9kq6wbvvMKtzz57l1
lYWvU197ZWzbUhIsTaZ0nfhTvWBoLfImQuVsBrZa/+EFjRVySmce/+VUv756xWAq
H5k6hGBEbSUIP+ECcE9V+cZGsoOAe4yOuiOdUR5AicswP8NVZ9gyK9IkfUWriJjr
flpt0ijiHuVl6K0NwFTkxTJTRlwD9tQluH2rSX4d+cNoZ2xOD5Mwt+Rm5YE6wg6Z
2V7uyPjUGXbDPpW42ZeSolcguP1QQSCRU/J4e1G9uuzD/G9byLchhtfZooYWrOjf
19sSwO7zsWeUJaM5E5Dp2yJj5j7KwHBnraTxdWjIOCiUxNoNhvGJusS5M7MfvB/6
Lfx81+s9rZy3df1Q43vF1g==
`protect END_PROTECTED
