`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GD3fS622UwNfvhaIDP5NeadIBqGh00da9t8QZVDPnvin3ch8/yvOTwFwy8ifMYdh
6Id4HCTcGFDef+IG7zL+JeVmWJIjpfwEHR0fCxsGVj+m2gWudQAMVlfKAXelIApS
+41h7/dEHX/Sml5KBrfbrYOB6BKHwgOc/Za4v5fXqggVqDYC4HA5MFqV5MoNPVAt
PZI0tevrwqwNA+fOwta9TvpOdGFLOyclaT1aOOIRe79ilQJ5N3iksbyT2Zh5dRGw
Fykdut9a4kdPJlR3B4iY1B9keZtMz13tyB/QP3ZoiYWuyZnMOKOunU1NJMChTEHY
Euf997noS+gc90Db8jBEuJNeWlfbrmq1Vqktcm65ws89TwAJyTtRnk2XW/HZURmy
jC65q9tK3NZ4XPXC4IKZZ8Wp+bG6qYxbkjsqNCijfD4EGr5HnU2tKcrAXs6DwYbm
u1f5j7laYGWpgdEOPY6BhNieDdZCAMzzcCXizSVlvn16tG5KbOA2I+IauBS7Nerx
MxVChaXFy8zThTDTeYqvCeBZYH3mZicnjkX8pjpvnb2xkVfbp8HdATlExKIX4Xa+
AQKGa9CesnW2vkeV5LtFrMGGDrEDf3mJJbmJjydETheOVS8/uvsvZNKKHhhIJ2/w
G0hYNk3EDaEIaLNeUmCCTYucb/n2aAkFZTKi8EpO1L1HCBIYDVvQeLTLIRHxaX8A
zQV9JLiPQ87N9lzP8QRDf5FWWWrhNG6oYQbhAD4c1eckUbszfvs3MlMQM+Zqcb7q
tEIDsIx3gCqHYQdzoSxb2u3SOgBFc8EpOEznS523LbcaNgqXE23guN+zvoktvN1y
QQec3ofz4R+eEAn00AlEta7uEd5eSxUy+XJgA3kRYGCXfXZKMaN2XIHj+snO4ASu
+BzumbD7I4yXF9pdknpZ8sHqBcq1BF/vPS6ynYpyZmLjW6IMhVPyFa6ZC7AgalRz
6ZyqnLlugvnV21VUqjzs+ZoZbGyRrOstT9gf0IwKSBUDG3BWQZ/Zz+BRr9ht4oVr
V8Vwigv1zYLOMVVTf7ocATvP6mGH4sT+P4766HB4lL71DSDarBXYXuR6tdBcrrqw
jPCsVJe8TyekI8ijlSs64SlPUVZG7oBrHIFT8EkCUGyhiKlh/PUod4PIZcU+zlGA
iMonQ+w1+SqAAMHywzPYsav3FaMyQSAc3Rj6p22l0xEQk0pMrAU9IbQ9S1iJdUyz
n0SrvpyzIJRxVizcR/Kb2TdMrYoRTQHghn6hjIlSkXdHcnhuJoqc5VjxX2i6XGHE
D9CvAA9yIhnXpP4C612LOPAn/FU8Cl1b376uvjiASMZxzbW70tyWatBU30bS1aZl
ZvUZ4F+68TLvWPhkpP237BJoZJTBmqbY4PQUPTiJPhsILO+KubSIrZz6tG+AkRKW
HwgR4/AGoC0uvh8JW/CnbQ==
`protect END_PROTECTED
