`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W5HVzwaCgFM3xm1mg5Kt5yVl+z25qz1PrtUEyNUe3bZTtlsIzpxERLOYpild0+9I
OYFNgwkGikET/CRkPvSE4UZAjacg7GUm9zArmRlg3SEot1cM74JtejjUhEF0KcUv
vglKGkdvQ+axqRVejiAb0bO9SFbURNZr9Y7xXhUAu7G9Pnfq12ap7duHxGYkh2jy
0IxMHuIycgD5U+DhabEHO3r+oLTXQNzXSRV6SWXciNnkWdTScmobx7Yof5jjRu0u
Y3fGucFlybVULJDYVSYCk3/iykRzDClnn2NY9dptoN9JmiXPpoJ93yfxT7uUEw0w
MMV6E6mBIj0z+IUFXJfltyvC2sP4bSfg/I9U/HG5oC04qh2C/y0Ob5WsXIZJPi1J
kg1XstUA/B/1VSvLjvSCfhTPiJdEm43LD/3UhH+kOICOj6nb1o7e5s8Es0k7oSQc
COXw3PCjeafQnP2bXzo2Tf6Pa9m9kImaXhARjSPQK5OcyqhyLP68SRUyel8lnovj
j8CW8f9L6YavBss+hqhCnQXHTTlOHztXZpfBfyejaaafL485zDroFqA959oe422T
Ccoy5amOoVsVJ/D1CQptjwqzaxlo5HHPesqL6D2/RE6/KSUlr92iKfbQB63KZXfV
cmvsYOn10YlHCrSn3ezZMhpjnleVFcDmF9LgIRrjlIHD7b2sFx6EvfYgxcr2LR7V
+NwEleVBDIPZMM9j6KaKGazLaaGRIzR9JhEgnN/1BenrUuppFkWaiOQCKFf7ePk2
NsgojyodgA7GiCKwthZsAdNqwuFkbIad+CdYYRCnp0elP78+CwkyU3zvx5Cl6fH4
SmPjyt8bpMBhc3uB6GMVkMKRKDlMAoa0xWpNWwUtS/oCC3wsp0Intp4MvAteeW+y
QD5akvqfRCg92NAgWfVH6A==
`protect END_PROTECTED
