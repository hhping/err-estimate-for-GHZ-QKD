`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvzYZfykab8rq3Ty3LyoGHgLuOBqjbXIN/rvodV7Km6Dt+KssZWa4gOGlVk9+sQ4
CwTOR8xXhrQGlq9Zo3fFaaEFpeyeI2VZqqzUQJNC/2S/jpmH7JN1g+zQnytapC//
qzZWRrU5E13FnBlD6mKPV22JfKkwG3dMGDrjXWZmjKUe6AQu0ckWCrdUgBYwOHGF
0lTP/ZSPfFWsrYWHKEW+LFkEIB624/ZPtT9h0iiYEuz/FxCwiQlnLNaLaUsJ60rT
sAEvBtHVHK9P+ziurLGB2yU6vCVVBoBo61L6FZvwNdqljnhZTClZxhLXhyD9ZL3T
14G9G/EoeO9WaEGazzLrb02U3vyJkumrp01T7C38f0ZDniA2xXXex1Hp0ERNP5kI
2/WzGVp2RMT0XbqsIgX5zDp95uGd/ntthhI8Id/SaeF2piyORqFQd2nXDB1Hgugc
1myQP3ogTv+oX/NUAcQ4GrEm82ByCWGTOfBPSXpmE4AwhEnAMtbOeWuS5yqPb1Vn
h0jShWpKkeHJifiN1Q3bwWbwIUJpcH5qBmHBUH3rJb6pYKkczMdINrDe31FhxDe9
6xSwDeSFP6sd7hFM0ZnbfM8oTkUDQSA87+/Imj7spLi9950mPcP7Fi/liPA2St16
uHHEqitOr3xNSi+ZKoqWKpsw5yTzFI484Qxd/+UJkWPYQpaZviktk3d5d4qLwPzK
t7XU6FXR+Cv8fcapr4/ZOyd6pIr4iK7hNKWjNaBvHG0YFYTLt60IOskwOrSYSIzN
vEqxtck/Nj12dgeHXI8uNF0MfRT7LWqgIIZXyjJ3+zGvK2YU5VAyK0zMRevbqocT
ycmesz7C8LuxOKdOSf91cGuF48rc/vDl9dFlGFZ7pF7eT2j8M0iF3Ncn5hzIIvwP
RrbiyZVcZw/HMYkqYy7KSy9eC8vq+goiJbop7kPam/esOmrTu52anjdxk6qMoKf1
GUmVJDTJazMaZsrGC23SvWYypws80M2Io+l+jaum3kaCZKG8ZvYeVWyZJe4evjDV
whg/fKG6qe7S9TSKKQhAXw7qZAvkD/lMG3Pi/g4k0bhWbqzyWAelYwVJQKdjls2+
ngpNrYbPZjaiRnvgJ8DcW3KL3YHZKuFwQtdbkHRiluBq4dC6T5b5eqhsHGh5A6uK
vHkNLs9rsfDArSKbLbVrkivbDsnPjTfyahSfDDFCOJjnbto1X5hS9G2FQftlj51x
nc2gzetupTfZkUXQktBFR///a+vj6RI0pXqVpaxM0fD+wpF0b1wJ/fP03+b2zhHG
LOibCq2SNlOsrm6DbGFpLyKHKO1HdBZJAJPGKVl+1mnzpoJV30M1aYOj3d8j2PL5
hVumhnhajRfOZD9hG7tQ2zWB6W8f7FrR5dpqcTh/zppFiIICMFRjOjlX6NmzKiqT
bIteG/zIJed3d3nRPaWPRXpGVBYYEkyUQerlI3UIKU4tZyAwNGT/3g751Ax9poIf
Y5zN+iU0ltTANpqwY7hzCmTi+hKZxS+Btk6Q8y/D1+cYafg7EEBQhsibwKsuNgbV
wYi9OmyB1w/pb8KK2ctPPyuX1mvpel5TkYaJA5JG9+3sDqt8rOQyX6OqKTG/M99e
47OfZxLsNWoqbYmmHsDXu46k2yOWOH0iXcSohEx4QjEIyvEZuaCU2lf9Pb1qfHMJ
82HYRryVRGoE98jKDoRJfoS8DXp4+MgciIJxXJZeSfRD3zuTwAVM9pLzj6+jYqYt
39ZtketQe/WcRm/QboMXoReveaChPV7sYS9UDAG7JG3dSN9U3s4CQpfMEhm7XyLE
8UjqgNS2QrscfCxcrmh1UGE4slFDUFKeDzsfr99sJArlVAWmJONXJJtI0tRSxBBk
QvKcZxIF1O8gukryBGk2zlVUuGOVdrCf2ekIi8T5torEuaCP7MctmCGaZI/7uzFP
GzhTs2fmPJ5Mv0F4kI+Ybuawvux/oQUX+Z1IimB+t09vgrDiD5STNCNgYUxpu8vE
QC6gVPQ/J4q7Q1ZVRsw3lGicvUWbGdgSpWaohIsJENrDnkuOupTyyo2FvTgPCuPA
hqjf0gyEN8R1wI7XGv01wWvZnoHuZ6KGZf0TtQt+6VOeSD8S/fA2aTwQPjAzgc2y
yEEBjVBwk2YhiAnH8VLcUBZR37hajXzF3yI+Qn+nJZFE7b5Rrk32NvgxO+ca2tmg
9dyGjz5LWuBdnHDsBngHkX9KlGJvncwP3Xgfp+6z3tdLChnz6deWT0QE/5oYPAOc
`protect END_PROTECTED
