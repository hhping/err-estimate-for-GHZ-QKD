`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoV/ZfVISTQNQS7sLhYFUvtRRyCOqBo6KCCf1o8ivv4pg8OOHioQNvKQe4iNycEm
mQSnNEIMS5MCihBjrS17hTTvQSCIzP8dIGhp4stXf2Kc1kjowZO8U/fh9bD0j99D
JisQOQ4gG17Ck9f+4GRiy33g/oux6uiVjCKz1pVvnxEtktlw+DlF3zJgvZXH9QgI
dNef7CJMTEJlU9TUj4s1NYerqVJOsYNWtHJ3iySZa1c3KcCdPic2JM0IboiQSc1k
kxsCi+uqDLOkUsNCa8qCGYOAngOwL2ePyioJagqZgeXbnEYRmr4KW7wgESUTPQvi
2fahGV/Ap9ld84CzIBEgdW2myehnLboX0YUg0yIhFH/DwGbvZhyYKziJh2zbPYQ1
0b6n/YBLJ+0aL7ieze8hLPoy0D7USRqUbGX38ijTbbllZgmS+A6hVUvAdyKhF+8A
mtg0CQCE0xpUrnVJ0aKOmvz05xl9daYi/4PCyDshLrO6N//sQCFFTzd4QUHe0NVb
Ve3rwAWu+8f1OUxJ3UhAsIjzgOyqvmclR+kjBMlgGK+XcRKUlhs8JfdYDEhrRTBm
bvlny4+icnOqWGPI8jbRnkvWK51oP1PvUoXn3We9Yf6UB/O+8FkuIoCIRTpJ8xWa
9VDXUTAucT707Vsx4nPm6Qw2H3o7uNcDM9PEAx1U+FeeJ4UGp13Dow3zlYRP5GTb
N3z3GKOZnYZ7E/bhx2Wmujk1NEgfRkttALw4INqqMjQlZr4ZJcsDWdNL5LTz8vak
/LULo9UsnmasBW0e0bL+t9m4F109hItReHlygdiVfDvksTjZleMG2hO7qifZEI2U
`protect END_PROTECTED
