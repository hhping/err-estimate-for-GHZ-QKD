`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeZtMoDaxiHm+ghb+UBwwh+Wk/9ZH511q14OG1wQG50sR4X+P4izN6CMlESkNK5I
RAaou+4OOCRCL1+m2uzY0VPF0mc+DzgiwWeZSaesBrJcggYQxgVpwrb9LqjwfL2p
fqmm16G+6aNli7DVKAznqkagw0NM+M7z2o7AIN0DcBw0nsyiuJ8FVUMPbBOxxIk2
gSoqKmZypZSFSW1HpQk1CMeewQW/EwcajsXBm0Fr+hA7rqijreP7txaLv3XzIK2o
iLoX5kzoMLUQg+DAtiFV1aKEwzj7iWeQwVYKybUSMlzMk0iHpwxb5XDZ3axcgxK6
RUFhx527IHLyLEh5WNLBafDrm48eKPT4FisENhQDINTb4nAtzKYGebBa3CB+L3S1
vz2Pa6JZZKaOJ2CCo6l1yzKrPExoCJsoUW8agh05cqH9roTSJRB/XFPVpXQLPVhV
Kg3F/nGcuiN56c7RJVAdcALijnFdS6vSF2hcQvMRs+XvQ0rdv3JVQx0EEslcpN7R
NxC9WB0IHgYNWW5K6Cbqs1qcn0ZEbJRK1BtzsQXafGO9HJIUw8OGZlv1HuBPlNyC
HG8W8jj5TBmwzkonUQI1524sU1Agnw3rcxFr4468yhFCrIvWPWIQbaOL6bZN20sO
cxQwcz/BJwZ5kLNN3YCvR+HMnzgBwwhdWey0zZbKA8spTcHnPip5ZvDIgNMg/2eE
1MSEk/JhKriTWP+zPUc+PHEjVL21k0nZWAEYpLCyNRdVfB3w4BTTWwWLE7HqGEaM
r6FE9uAyiBQPpO3FcFo8NcQKPb3iU9MqMW01AZyIhrpvePioyzAMlhV2bCGAIIBH
2iaqVqyabLwkByCYY7e46KCKZsfwa3XsiVtC0dbhgU4yy0bfev/ZTaOCgQVltcTP
Oc36oh/pL+tnQno2hjhNcUjM8YllaVIuAi4sBWY79mzm1juw2qie0RRvtdLJ3Vcy
YIGXRBeKUyv06XnCb5ziqw+kp0sfRPmSo3ovWeVC/75KoA+18YgXhMFcr4zbCutU
UA5tV+djQgkywdMGCYysm65zPicTkLZBcuBVKRNXSI7HSQqhy83r8iuNBMvnpQ4b
sDTlGtmH/R1vE3B/TxBDCB9LFGKv/WEwvkPahR9fZRR5JS/5yqbJfEpk3O4Usq81
3hkxrVzHTv2jnnaddWQeMlObIHGJmLpBA0GZz69SjhM9i7uvkJhmwQE2xuytDDot
ZIEzFrSOTgVcWGEYkZIGMpj11+AcI7CHUScc3Tk6IMkeR9mOIjHduDNCSPla+71f
mxk36pveArDKxILt1nxXY1WN/O+bPsuEt+ypKximCWUUJNATYH71Q4aBfZjELfQ1
rK0VDD8yBvclBFKVR0+wekXexYhHGRaDguUp2xxR6TBLrNQLc/HMVGoqnh8qN7sQ
cGBKU0xzh4jFNXGWhGWmZcp+vlJwfxbrwQHhZgt0rrw+1rTqDSH8jS8u/bxL7V43
Ht6ZupKr8ndaMaWJoN6+YV4AltefqsHdmXoXrfrgdnXlXJhkQHAVAav2oZx1MkFg
z+hbMxWOjpIwEXJgAOvDGbgL+QAKJBSwTZH+QaQNWYtX75j/64uldOHWiavZxp3o
vm9dgcutetatCZmjhCNfKwjZAWw5SlfhtBNpAsryLI0=
`protect END_PROTECTED
