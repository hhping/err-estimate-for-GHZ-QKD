`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SPKQQ72VELqTWCKA3smiPL9Hnc1IrDYDBHJLtN8rhrXKkintkeFqSQomxAhbhqXv
GZE8AlyENByp47W3rUaZLPFe6yfqPSILHy/91BoGRaospRyFrpmkeopUOvyQHasI
thOoLVlnYfYNpwy99pavL68S8G9WJhGfZdHUxnQ9IhN5Cb7X7cUHnGlSBYQOi3TL
lKIAc6TdhYBXWiFBcPQ6sqQ0NxEHdeaYPv1Ep6HZ4S6DJ5LSZNR8oz8CUAp2NmXY
`protect END_PROTECTED
