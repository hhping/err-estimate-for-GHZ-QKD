`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kCjBkyZeB9L7s1WMpLw85vxO9Tx6iAgZOUXET/YHMQXO8NWRPbqV2SXgCfwuocd8
MWCt9OSmta6yM5jbi4+XiFhJClyFmk+8uTVbFQW8D4P5sa7JbV3wWwaYiKmt+IZy
boHFu26tYARspv4W6XL3IreSFIEHnEwVH3zbGT/A8zninxHZmbFzx/crMEqBmyYw
+9uRpokowmDVVXfzPc+iLDsNbBkwj5G6ghJdcBfOiMO8dfJosHSKm8TSNwrB3pED
LjkTcnUvti7C+RJohp+rhQOswb1leTC6XRzcoDIDR/9r4kkp/vNbhgERzVBcT3b/
R429w1r/Xc9CcW3UoI0uW7jEUrxHp/1RiYm9okuCI3yI+yEuu8FTmad4TBcTsGCg
FZx/84b4SIszq7PtHOZMaiUxaf4Nu6BpanfoLeTrPhws2ifkcQs40XeD2imUwVud
J315PfkgjdMpz44qwZt+a8/j33NEH+/pwmLmDa22L0gBZRjAWUkUsUZsRHBz1tbs
EKKZ/n+JNDvPuVUH1PXE9MVddANBA7V9FbxUrI/c0snDDUDervGwnrVcikwBTH5X
HtrnjVWzL+4K+ZAWUGre9369/z/RWvG+xNU3Jy7Hetgn6VHUO9XZHv7GB3Xu/QbI
gC4s2z2GaoD8TUL2KUknUQzA59rED2Hd1pMCa9cdALx5ENxZc/Y3zXH0zlD03wgC
rkLYp8GTLgXP2lHnKnYw+PYUqUM71yQq6SnLHdKpWHCUXafUpMVTL3NxWA0ZQ/YR
6uVigbFfapb4SweRfY8tj+nQpL2u8c+GLwaNPxJbfd4agGZ7VxbbZRRKTVxSfr6j
M7ng4phQGiLysj9qZfsktqUOdMwpK09qU+NS0oAXTktdFVhoalVnSmrB2V/a1Bmi
9k/i8/IVinU7NxKOGqpyPOVFaNoHko24CTgnFPlFTGxVLhLqbC8mBPYdH8w5xahP
hYJY/IuwxqqDa3LJtNjqNjnE842SV9wozlcs6rQu59Yv+l2xdq6AVAXoBEHB13PK
2E8fENJ+XZ+YoWhh5G31wgb+0Rz5vjq7gmlA3KqUhqv5DwRXeV/H5x3320i8799y
dQUzX4A8fmY3VL7L7pEFO0/sdNyj8+DEDUcHbJsJvla4bQ+QJ2oH6mjx5qvCuXi1
W/bvqRLter64JICiVHdXz7b38m8yuiTJbf8H5aAkGqSdE+vL6IT0Grq3CrWenlVk
VxHa1RhSoAFt+uomkqf6AC/pjnyc7K7RANa82y0exhfsuUgD0wu2IW3Z6PeT9Rel
zb436RKD9dPuBrnCp76KJL/iW/1Eo9YbvWc5MrlAtFMOwvhd7lA2ufCOLIWacL9F
4GiDlYvGaxvQ+hmj6GNOnH1e/A6hmPQHjCQjmY1OQBT4aZ9CitYo90anklR1WdcV
Hv0QcuPynBxT4RWi3j+3sTMoCr7XPST6ar4lU0AsZA+DE/5jR0ya7jKqnt+ClNW4
dRdtubUKvlun61qkmes6Ciqw10BOuZkKZFTPbust8ub5rVGoQVTrCSAG2VRQHooW
DD3Humhh3dMm5qkpNhsAysk3GtQ/657qw+W6hAoFLFKUSTPmszzyOg/83Uxf8Xfl
WgL3eFimmQ01tCmL1y/wK9SDLJt9q8G4owMseCq3kYCkahkHPUA1HNI6CXtgcxco
E7BdlzFBoWwvamlEuHQNfpbBa55ufdYQUJKchFV1TgkQ5kuaXIIZllTnOutc2jaD
BSRKZiQPH9cGel9frq+eNQa5Qoz6Iyo/OqHuQ8PN6zAaFDw5O2+WR1K94xTx7DI5
dT6u4JKWA6EL3eFp9JExwYx5z6HgXyf5E0utLkrtG48DDA59J/0xOb/Qa8A9g8rD
aDylZuAQbuyRSBvH3B9I2L5XzmwJmY0MrEq14jduL+fJKKkE9Pjk2DJnsSc2Bugu
Kta9pOK4eHH6egsOyiRUSPSWJYjLOIzEX3Zd5CQ8CAnKwL+gzsbLNzUcoHmDwu5I
FnToIZjWIaGqSy9Ut5gJ5ONEBBKeeqyopy3keGhrIOVruHDkEYWZVSYnmEnpJNlt
7H5Gpjxif/Mxoxzo0/+XY3yWb3uw4VEEGxaxwq84aOzJXOwCzDcjrJs6QYxB5jn7
RZeYlMz8qgdzhcqVLF5hLx/SGXGe+gc55+iLNvy9K4DPz7moPBGngVcH5HXyuoeH
CQJcnrVX3YXEVFXdOpyIjY/uHD8Dl73yJgsYZgCe8+04MoVWkRjVF27KbpexUx56
hgjkSzYL1rF9HHykwKsNub5UZmLHalQbojaNHfg6sngJ2Q0/sjEi8y5KZ4vy3uBg
tGXamrjj2acx8iTfQYkEQKA3+FTfvJ2ZLJiYI0X83483QoPiIYkFOl/8VO9U6FQ4
DyTJN+XUDXumd3HOGUZSvRQVLk9cWfXUXRx9mO/Fl4zlcZfan5hxmdq5f4VBzXEu
MxwYKOtLZoSalGrlYrUQjKxSazdr5bcw6Kx5fse3OsmNI0tKDp66pAKQiWH3fn+S
aCaEH9puv29CmO14/lnuPOvXVkT27SSEaQxcMMrnA+VK/rJV3yEvOfOKAQWY8s+E
Ev/66SGS4uZIuzuIILBA0NxL0//O799/sjdCgpJuKmFSzMhllLzYAAl6w7Uw4ys8
g0YJli5nyxPHjf143f9I2PIjn9v28PoeMBk+576HRTD80KwASzRw1xXPJ5QRuqso
6UWTjPBmzScN4sj3li4u/0s+0iYguMMWWkPldUIIolRwn2QpwQAAhiMAJsvpm7RM
aSmlpdfvkxqC7HEeZ/oMG4gBjjSyGdBm5L3rqP3/LyYiN94wVKwtR3Qj1mxaor7C
Zy7OMPHs03qxj1IrM6GaeF9dpPEqRXzLo2ICWxUxgjkm5hkz5b2mMpg+Ytnp0UeT
XP/pC4LnCHo/tkSgRKiNodnMvPN0MZK58yStZV59if7VqWw8uD020l3FG4vugHmL
m67Dzx6RBhIeWpyKhTyaBuOflaf9/q2+oDEjymCmCSVVb4I82sb0X0s2514SYxJf
+nWTVanegw576w77zvQKbh0Vlc53PSOYiQc67VMpcxI=
`protect END_PROTECTED
