`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6larHAoGFItgVT0+h2rc7VGE0PNOmnw019jaE5Aekq0BweBBB3vCHc+XeeLoNApt
OSk97EbmA5YbPIuRi3Sn9sBXns2mqehyipSGSepQe4RrH6vXUvCGAxLKI5LcWVrE
PZGWiQCxUJQm6+8mcSTURnyvtgRylIMvagdKTAkrdJDGRb3F0Jtdq76MzsrIiMM+
QdQzuF7M2yOmOhjzZWlrNMotn71g9ByHmOcS/e90jUIC+S3BqOQB4IwyZ/llh8xY
7kDAjT2jN0Zw9SZMmX675lfgTXqg4z6rzZ2PeGNA1RzlP8cBl6QvFGNo2n4M3sHs
8Vkb/H4r9QitFbU8STUyHb+Xm+sxuBX/Mk1UbbcupZBUWguJidy0WawqMNx9f7o9
bKEzq6eu2I4QNefXnVRb+Hp4fctViR1j8Amsg79qarSbhp63Gw2KA/sqmkkcz3xs
fmwuL5UGL4KS6aAldxT+lTdPihlMpbiwu87urJbsEEcOjW8h1n1euPIwJJQOvYXc
lMIa1SNwNS1LzVL2pZQjsBGskbYQ/LlOhWD79jpavCcXP0HjjwxjGgGcF9jnqE+q
S6+LCGLuq5W7gLhInCDqtISf/t2vc6MG06+mu/NgQJJ8+ScNvGnCsHlji3q0WM7D
O7QJltcorYyEzJLH0PpJbqs11uGUV/Kf/ahS/Gh7eNAZ7mZaOCtDppR4NyrjBnkL
M6f4mneo6c+Wkc4vb+2WCkJRoZpyFtbO0DY95zcgM/FS2dVo55GE3sWUeybVUoYh
`protect END_PROTECTED
