`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fq7W1DM7kapoj1EKeVS8JhfHwv0O/XHvCytQB/zppoHeGg8Lxx5uE8Wkyyqvzd0m
my6rr2WDdLO79ykhsZDDTtK/OdZD8Uj7s/eGXhxU7rxD6bwDZ1W3iB9rBw9fcBZd
JGQ5mTLIZvob0j6J9T1zOAChrUWBCnEV9G+vWJUHpj4pHNTs48TkHaU6BFkPfpea
/RDByxWubWQtvXn6yQNhtgVETZM/il8fwNjTFUSadvWT134kmfu9VA+CmiDls4Q0
8JqqRAiB6b5gTHA/bV0LqAlh0RamaVvD/5z7AiSj7c5AHfQuVBzKCSHjk4t71kjo
ksaDK+E4BMjGBxkSFskrpphXo+VC7U5bQP1sUC7T2F8Yriyl/0ORgIiZF9FXNnkO
Gh5C/FDyDK5CYtObYaW3MCC80aopoujaYFytvd0dfU6vSMrXLCxKsWRR0g71GmLd
p5fR9k7lLPuNen37nAsUN32EoqVhHOygBAvaIaXjxIYlqTrTTk2AsuvoQ89KpNs5
z6SOVxhkubbFFGZ0y+GKNUzYDZUx6kHRP5QdKlumGm8ftdrkYLmIcSGYdPORXd18
4k5oUbo80yrPY00wUcj/yo0Vmdg2a1Fzb97d5/lXnW8Wns95Z5ycxe/YcnnbIjum
T1fSo2NGJ1PvuJ49sdfPx/b1ZidJ6hbzlXM1sx0Mv4QxvZ4XBC02nzaznnMehGkb
3HSLoBQm+E5l6qmEQKOntJ49HF098AeziobovA7z36dD6VtUeU1hHfAy1tDeX4g7
Kc44uklX3vODSIait/xLFHmVDrq7RRGH5rveH8AWxBqxLQ18EbcEF8ewsB9rxFjt
PDjYiGi9TCO0fI2Fsl/EKLFrQ45cgXvobyFPsWfJkhlUVQzZ7gUl7FcTUJ7uML8+
M7LQxf9aH5PfzTmxmxG6TnqHt7aoxPVPGE0g4NvJpzHRZJCOIGOa9fKnEUG7hBWI
Mjw0rxrwQe8cz4GxpFm0kqwvWYqFYWppns8eAyRAvlnGLrETPupSApH0FRR84Uoy
FtWMwBxeXn/mvAhBpyry9XTb7K+R34bCFgbgbWg4L68t0DaiULgD0YKSn7i9m3Sp
YXLnvguncYD4dKKEEQghLVswG1/ZlvpwTroPYBrTb193/NIeBY+NsXlfkvrQRDdj
FVn6bUac+uEDoq7ZDdFTuj+Mr+dc2BOmVU1d3N5byJ0dTfPiH439SX1IAbkdrThJ
zYDBMDAvnx59vKUcBIsVtQOFhvPk1FAw1YEcc6aQpOD0zpUtF55bDyqxszCyeifh
/DWtDYRVHA/3S/oAc4i9XYCyUgj8z+63T7loZ0YUOEUUa6JoVwYGfHJ/3W1JYPK5
oo2IrVzos/ucQslnoCzXWLZD1df3OJU/DjbnqHy95FuhY9wIT8ggGdp00GsMe3U4
YzG8BHzUJe5443P3p8isBFEr6eSF/CAYEYT4dgr+eMDxVQWKL+dwfU8wZWPMnYfx
A94Dcb+wCYtfhq+VveBe2NXQgtFFlAj+ntOWVk5zLnnMveiHJejdwR41BoQU4qOE
KBWGaZJJFPkaGyHqVPqNqMfd0qz8yLamK5kZ2pBExIwz+8pJdIq5Pdk+cNBxydN6
6q2im/OqQWohdqoXXn19j3E4vkfiIztCrkPzD9gJcYsr6LF8C5zqP0EmGIrcF6p8
vKXlncNp9pfashi8nn4N/Gwpwq7i6AolInDWhESU5cdDMPqYbT/NZVqlSwUUj9N6
6JZ2WMNcnQkRPfHHSyoHYFkt6oo3ZsA50GuO7x5yTa/nL11iIAHtp9bmuMOUkbJy
4VHqZ28ffr8AvUWJHG2EvpIjL6SbnqqDA007OlWu/5QREQemZyLiYc7jSJ4OOlxy
GcmTW/naK/iuuI26R1MjbQ9mS+VfN9N5VA2Zur9TDYYkCwOs1u8NBaWYyXyiUbHR
6AUGH+R7a/K6jl4MG+1DxpFbRZH4pfhlKXjy7/cpIE/ASng45OHX32fW4tHjHGo8
AI5qbQzjldhTMFt5nf6Svtqd6N9KV3wIg9nw+GPVH9xdPZZoqsja6RzrsKdadvNy
dRu2rREhfVvVV7ep+e64zMHPYJ61swf+EgvcIT0YT+Fhu13JbSRHUrrqkmPNfvFs
WMCyAh2/MrhRynB7sFAi0a8oxpaEVEhFx8kZx4OhTirN2U6ZnYCCwA/qAaQk/rIC
j1dWax0Kiw0oqXIpXqT5qXhEDsL0VY0LvC3nb2ufQAy4AD90dg708ErPO5Zjz3la
oJjK1ZoF/Rx1meMRuAOvIfoAEUzBAe+3geavw1KP6R1nPzm82o71I2b78bvDoaAl
xQJNn4zkXADUmbCyNDjguG1PDfzZcLStPXeSFOqzR7/oEMRmshRYr+km+w1QLb23
k9V5aF7fEbBPf4rZEdPsOirMOHec7WE/fmXAfW2Pj7PhOceT0OuG1MS8vVZ/qhzI
V9e0QLSRD9L+mKgTnut4NTiATIW7eRWANB6XTi/9q76qWSFIaaEZxPb3alvZcGXP
wMRM+UJ2Lao/xvDL8s3agDPdTel3MZE8uRQaArK4HbuJO0rYktF1THipj8FppIWJ
csW1uXcWnqSBhsWdxMxo6l057isydY8L7jbePK7U8fDibVsO09CEOeFTERdwbqjl
2kipJJdiyBzKSbJGGeKvuWYYXnAjLaIE4dUFJHLNVdfxHKutVwQ1BnajFd3ep5Hq
Fh3mf6eGqCvQok3ON8DmqnYsdyFreslgJb4JRS9KfjiIh4gPS/WtJA9u/mkrIukR
L9/goPqCsihZfQDJ5z9qC4F4PcQ31QAK9ucATg+pGcirpvgvf+Pcm1WKF4tWamFq
RA70qGQ9i1cLCqQXHqFYPSk9Xf2OMOm5lWwvSBCU+JCTre0AaFwVX2vP/hV7JOjI
qe6V61RaF+yBYGTt6xkkJ2QEUFjn1ZGstl+RZG/Aq5xe9whxUgR/PJB13p5pZ+zJ
xFBdlxQSKBxivnLfkj5t1q613776k0HxM8eMCvjLcNQhWNajuHMqUTGnxvJo+Fig
/7udUYLBsEAciXEjQtU5pgWwqZ/MhOQmhZoc1xA5Y8g5VAWmDHgjJwkCqynk5yKi
+zwF741ZX75jAexVE3/Vp1TlQprGkGpyzTriSyZ75JH22SvK8OepZ09FB0AQ9Db9
VKCFP+4f/YwAdGBlX3O3LYW9JZhXVfCyZogcmswVvZ5v/356TosXxamNoxYmJ0aK
1VT3P/PVLKaHRf42O97+DtXSEVA4RJFQrAJPWG8FCRUiUcn8yd4n5JjAy+5quJHN
2rwIc4BdO1dxQ4DjDFYo1PACM7GtM/TU8C0IO2zNx1QmqxZ0vrY3TlY+NSmXH849
aLuQxkEX5W70CDaw+8FgnpXObTr34ENMkOL++awL21vwenE6YEgFzEalgfsslMOA
OV6rQEUJjGwyR5F9HXf8Fx17g+0IhSSQ5dFf66f2C2DbuNxKUo11K4hGsjpdsaaE
jnRJKHuYpyTYWrXA0fGl3KGEws5qt4lfyITkjMNR81jEgOyrX4y97PWgd35CbXQH
GTiZMX44CwODylUoM5D0QeT3Ib0g+N2QTuozbAdpDVDjYJODTbeceiVeaeflxc4Y
npkNAnx4sQYKrV2MtvwsYto14hahTMEtTd94MV0Vnub6FtSKAxWBkTuemC6eAzA3
d9wfGJ+u34l940oqTgo5tIPUwr/i0Zr3oJunqCkk32BiZK+/FFvGlbEKe6cMokGR
qhhwkzKpa5u01pM/69xXAwrRiXjXmB6Wbug7tYY5k1Tjt0RuNxybI4xPQ7GnZA8S
jaM/bh+kyIyPre6Ao3FGS4P+w1k/3qeaGs47ED22m4QO5o5RQHUMp0xQmgA/pa6b
ktCmPRPT4PIvFXvX5NWbZIkcUrID5Mqk5X9Lz0kZ2p8r/FmMIK8Tn70pgkqMmjQ4
KSD835rHor8Y3/9qs2egOdV8/Q7v808s7eC3YwLzHZsFNSYDYBtOLWswbQUATRi3
1ZtFnajrANESk6+trQX/VTSf6ShKI+km/oSaVy+nHO31hiKTk8t8YOYak5aB5+lW
jd62sqf6Ebbz19sBRNwdGMvv+HAUi68N4SUqdWes6BYnylXyavVG9yjOspXIuuDz
IgWf5HJocUX65WJnTMRK3DfJ2XaqSXodAAscGXy3DD0pBbionpMajahJQkZItlhi
o55Rgrcb1jLUVqMC8yP9X8EaRfXvHsmsLUEZbtgy/nHutg17uDcy4brQ1skZaQyN
4sCOSVWO8rwZt1IywLnKzH9NyfKkSENqFJgsP1meLppDeXnn+uLzhFoYXeISeq0G
`protect END_PROTECTED
