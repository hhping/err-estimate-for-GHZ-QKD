`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IVqxF2uSnr4wgE4g7j5uQXjqzdvshnhkwGLnFQrhuzgpuWDHwHntAPXviBVfD9Sz
ONYyYAITSVCkQWQElH9uyO1A0fTNaPyfJ9i8i9TYqFM6jPgyE8TWPJVmBExPBTHP
nvSqIp1YSZmFyhVx1+mCvWGWT0xX59OsmCUKT0/ioIcfyWR9HTS5QqDaW66Yv/dE
kim237Fn/esqUW6N11nA5NfEkfdjndsoTLgSP9VnOyZYpLT1ctUQ2B1dIL7QsGs+
KZ5jeVoNecHrFJHWqtUo70a+KQgIli2PKCR+6pdtJUtC2ghunKcjOMhf1Ps7uyAl
7t8sKyhDZbkfdAY9CJ9j7zuie9yF5v04l4giag8JF67BgM/iOhOViTDj/viHYzsG
uwjXKnetsUkND+dbj3rAq2Cikao3Qqo/YVR0yczRJPmGzHUn3UZ09eG6RcQ+J3hp
dyf7WLzOflGYSOXfaQOlP89S1dyDCI93yF6yseCzW2Xv3Bg9Li+Zla2IdhE7hGLe
HylhZi+mWPobzQeEJMLvtXMVfEtPnQY0yars/IhyY3QxGMuFQtecKikHriMvWfnS
BGc2gRRWjWPv+VafWZvrLcideQ5ZH+W31StLF/lqbPVTHbzlyzgMx5MWiE8hlUCL
hXUFc3tdqpx0g5tjz+ukLCLIRjVhQ/ZLH2ymwO5WXWcgROosdCLianVCdJIS59SE
do4egJKNUGpoMPNHcjb1Eph8yPbzAIRI4cUoVll4ECUj+S4oGkVTpwEeavHHGUFO
GNvtNz7s03Bs+xKLUWLyvcoX/3ESYWOgf8Hm3EvD0eG4Q7tgr9XG7hUKaPVTmk0Q
44l3RtQ09+M3jVI1a42R/Vh0SxjlPXesvQWWx+lxcUv0dEZtEyrKEDBO+OEPbiR4
KMIOaznkX+XvQdg+giFozgsvMB4zIwgXhis6vYkWrEcFocDE1JCDf9xNe9o/a2WL
L30EP+M1NbnlBkqYGUNueZ0pOJv3OZMV7vafCpa6JCmV0zaFuX+i5QdTdVMrDtcu
0RHVZ83M+XY96vlB4oyTPdP1fsWTmCKNTu8cuN+HvTsHnqvpJEV6ZMUx9KgfwoIE
wtKktW5xGW2GHcFIeukJ1sH3OQrjDv0fg7Oz/gR1JMmfS9PeRO0Fao5kI44N3nfC
PrwQd7UmyGgG/XwwYCYK0/IGM8FFxS18nQs8W55eaUKyrlBPS4t9lcEKFC0Ytf2m
oMNgT9/ipZPujPI15bvTgrq8vN+JWkv9MP5iZ5sjm7k7TGR1UZDABWoDJbamGz8n
pVNbwUjatZ99UiGmddfvllyoQkCa4eMiwURzw/mGOrtotheuzwxYmIV46ww9124i
YEJ2XsttJJnZab3pihp8KuMlkahQ98DAKmeTR1eNxgy2Vfijdbx83htgQQZHTlI3
zmglFOdHjgCt1YlqEdTOjd492cGJOOIEbUoz27sY23QniDL3AHYwBOs8feG5p5bb
+gC6lpuAwFjtAQ7K3XBRuzBamhLqvNiKI91CpL4XWXiBBP4LVtNpnGsvEp1iKoT1
S8anpKo9+G7oP8SdXyEU+BfWF2nEBnKU3C37nwzZUIMSJfJm0BlWVlIXZTeOewRq
msgZ69/6fIRd4ZFs6d3dOHT0HomnstPbK0X/M5HG24CgY9ZYU+yM3dOQWZTAd1PH
6PlFvI+Y/xtukO8QdtlTWLbkPQoYesSZ2kR/61ymvco2n2bqKMxi6bfVTvxb6VpS
E/gr4ElQfeeUMoCyT6u4D2F8aH+6rWH0THapBtJTKJSOga77enylSq7nhaJH71/B
qAOq9NtrFWWsjIQyJCepy+8/ZggjBoOgR9iJMDONHU4YJEap52PkqAB5/YMaLOfO
zpI1BKurLNTaMXqd8HXIBC/Ph9viAV1wMkc2tVMazdZFByqxTeQDSWoSOSAdw9d+
z/LW7QsBSv/cTcewkEdZXg==
`protect END_PROTECTED
