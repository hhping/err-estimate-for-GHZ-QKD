`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z+wdYjkmKYhsiH/Hr1qazwV1MaWnfFmdasfWMZACAiehDleBmcBVg4mPZG56L/Ni
qULKBKPC4+HrzUfPnlQSCjjVoZ+k7Bt9xJque31hHSWeXKNhoxjEhTEfNzhSfRJt
/xTm+3ZbBj3Fe5Vw07UAiv57GJn/V2xTbJ/H1aMdZe/YW6Wlvj7hkutHgzkNPQU4
BW4d0MuRN5y1Jwk9acLYygLZpahaNCCwoJEAm5gwtazbHdFzFHrNMb5m+vw5CnMZ
9CFoCuNzggRewSN5/8GI4EHaQ6zX4vXDhe5Te28DIDQl0hcZUOz35bivoSQt1kll
0FcHOhGnmHWHEo0asZGBpGp4AUvN6dosw6VjFRpBeTthujF16rASwXnUOZKM/KcE
KpS2FWXRMx5Gs5ez+DV6Z1QuUhm/VrbZ8lCLhMTw0fWMXt+6NwegCIVpS7RBWJX0
f9IgrVgf/jEBU6EuGtRGDJkGmoEadzRJbDz8DmkpRG5zAvdhnfHLBbdbS13vHMPD
YuOeJFKJSL6EzcWb17e7cZsAWMnk2392KWJNoQS041XM40/BP+cbwZN1LoAhxuUq
kDv7eHxm36ghNxp4HvuL834+3xKzFecc+uK1QDsoybWbvE5NgM+3mvdBkfIKWkMX
LooVRyLtYg6v84etW9EHGY/gy+yGIOHpbPZpm0Kr4bjtFQik3w0VQ/c6xNkd2DK5
gkA84ZPu5zEq4KzHXbPUKyImVUoVze4BeiQSxura8FQkF8jTbLJXoa9HNMIzMbH2
jUCqOdCXFHGjGH5sqdpQsT/vv0xf4FCaXOBeguTUbiQdNuO1oYR3ehy5c7AGvT+V
Ce1ewKlCZ///IizrZa2AbHZjIvJdf3OfNqpUTvhNaN+4aXq6nZfoiAfGj3Hg055c
0SD+rXBEQHjDZzTfV7hN//6vpJdSZcrHeHBl32eAroEXN6nFIJ34pjcONqYDShN1
/7dlg8aQMD7GorolLhGqYLX+hIruCoJdADv6GxJOb0F2mQD0dGnGULWxcGET1z6z
Gpbp9OC72UJEA5a84hHk63sq3t3D2HaKAvNoxS3z9FU=
`protect END_PROTECTED
