`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4C2SIIE6zCaeXuAYpkfeCKGdO43XgxsX1dx9KPnjITHyCB4DOVHosv4wHSNMAXz
VyU5sacXmG1tzWbSNtMUDB08glLDfMGIhbxl4kGx73fSVtX0kLfIud9QolEgRT91
f/rduLAsS8u8BeCkHdFtSIS67r4B78E4qGBDUGcDWwIbd1qFoAabPiWKC2NPue9n
qo2aG9Hpfu9glEepDzKJA+PPby3at5iTfWEZ7the4G+1y21eiTLA4GpEuENCbCLt
ySsCUp+FGLNJg+6HKJxPnmpIym3ym4mrO+W8/FmOX/ECm/qg9aLSjaB5Fl49VJBP
yeG5dqO+0olGx2HZ+T+zxZWC+itVeIYQnqgVTuS3vobGciydUrqIUAeLOTddKhQD
gmXncsnJAOAYvbqpJ3pANfDtwWPEh8iql338mGir1s1LQ1M8aKkYFmyz30OJ9Gd6
4ZW7yTZVDWp59pADS3XpnNDlJUq0goi2kC/wS8gTmHft1NdsV7t5CIkx3S4XaWKh
WEZR4t2PRgdEoXWs8eAIX43LE3e0vTHjwgU+H88BRA6nr5+rdDzQETpcRUYJdcl0
mxfk3TdUzVTAOF5cWl6Opu5lKEwyw6PtPkcilwEhLTeHJeOLZj80GE6CLs+6iHP6
bs02NnbFvSuzWdVN/4MNjJq19wSpxmg/nZ/rEx0WWGI/ELhbD9DaayRPcS34LeSF
cs5l3IV+f6KmOI+gZPPkGZvbGzPPWqVksX+Ev0r8Ov6dFNcKhv5JgqVKfb+wopIS
RuAwMggFmRLhp4BtXsuzxcjFKCYo0/MrFbpcqirXcbo=
`protect END_PROTECTED
