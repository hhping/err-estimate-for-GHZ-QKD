`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZLdPz/ddbXbbabAULCj0HzSYa97PkhYQcwcOjd/Sjx78wA7z/RnugwjfemrjopPz
cRkGdLsej1DfXCOkjWxOy1RaOb5aLcv4MsKYaHQ2dZ9scvq+IKebhca7rV2wTqxN
Rzm81Or1mq8irrKGbGhd9qeZnya29I0ec8dkE4kpEIeZmm/VRxfkRdk+vog9XYjK
j5ifRIhC6kFns+GmUTXuRrhN0oeyOIT77BsVkyKh+coWGQDN2OAPrG2XT6ynE+7Q
6xqzAh57UlyVQzOq5RsiNR3aWln3ibE+cOt5CsQr8ctpkDGhjkKXFZNFoODbiJjt
iPbh8cDeF7qAgu5jnAefc+KdqxcYMkQEBSsIlwSbi6Y2KJj1SS28Kps/J2D8K4X+
zFYDOfE3SyGdsenhXrTB4ln6udhjCIzOXNeImZ8xZ9mdkRfX+x8TwuZygetwFpK6
4UJWNphk6m5ZC1wqvF8usItXXeVgqijVNGiugIw8RMUNMu+m/45i0TUNVqAHrB3j
cxWu0PzQOmG42DkWhJCcnq700vFZ01Imdwu31p0331luqav6FKbg/VV9QzLmfJOz
C5oj2fSYtee7S1rkdZQZbuUJ/93/sNB69RrgO1grnvY=
`protect END_PROTECTED
