`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9421VBKvAe1+hVmVV59qDRHFHvkdLUmA6kDV9gFir+BD0D8Gl67OPujNeOeGwcsC
IL3mIeHMqAczW8i8cx8g1dSWMhnf+CmEofE+wWBbj+/b2Tec0UPNhOeCzA8bu04U
dr9H22Ymec1zmeLFWj4IZ/zEvQUhx3fLK+24V8vjIt+SYfy+FOKd54UNaRG7k3xv
89Hn7S5soJxDuswq0EXGszx3I8BvFEV/3rGVdQihMmAyNdGrWqHxwqcNXbX68Lhh
g8kAnHrEsv3ju4csVFF3HMdzFqtY6SVOmjMG5CKRGplQK/OVVH1Y7WP8Muo7NVWb
b+BOaz8eMRN3HvXMIsaNY1fzztLdpO6IyQuUmByFT6RStU2G/5sWm3kydFTsMYpk
QvLp3qJ+4+sypPisLgcwnicx9VPmClIr6PrAa4ozlXs1y7ClIv/xq470TVsJAuNa
He+nzymMjU1Zz6zFzMzc1ggkaiwLTucwAjHXNC+/jN+4YzLUKu9WJfN8O0frKWtF
EwIGxPzOBwFfJDSUHBuXtqUh5FyWY0PsDqLbR2B2akgI6ALrFeYBhjWpiLX8UXdW
PGUcs/4ivL30B8SAcXJido6aexB3/p2+/acUDXnFMnXpmxL5SYECegWEbgd5HP7a
n4EB1IN/zg+rdtXmX2JCGP+4VaCAZSXdpei8K3g+dgWXtUEZ6tzy0QHlZrOslbvh
dW2FDdp7clNBOWzJHlawES+erwvRF2fiEzbofXkTGDXOBXDxOPL39MZRhASnS59U
T/IZthP2MqExEi3hxBUC6Ah2nmz8Fzd4EjT7FwUJSt5Nujmh76tdu50frX/2d3Md
UaNeWFx03jCfwFVcARZCwJ68G9R8MFgB7N0AubrXmu8HM6XiISNzWhUGzyxQh1vG
MBCUStfLZmkFX+PdKWRXPoGk/5z0356YbvLig0XO9CdIyidkFqQQ6WXhov1DK6M4
eQD9EdUS9RlQFVFvkumlbdiKFXZ06fKjhNN8AenxwIFJhJImX37sfzHV/p2Yo6qM
kV15wVxCh/7bQ6YdoxJ5ULo3m25RceOchNJIEQVwJxdTp+3ENoduIoHi9NlufpIA
EnTm+qfXv19uydPCs+kSfbfgmS9HQZUlD8ZPXzYfb7JlY9Lq23i04ApwyiG39qqJ
aa5jz/UpZ07X4avi2ScKKrI7hdvbeAx84rlGVxr6Hcih+xOY6YKNGVXQPgtkETU3
jRwoJW4kEP5bHvBXpOsbN5psw2SlsIhswTxslohU3Hcb9FDFE2kwrWNbkLpX180N
m9DpJKe9Nsey+1p07rMrv19ySHRGYUFi4hDDvxAdoEC0E3usPLaNaodZITDJvloK
IfIm4cCACe5J3vwmnbv/Uhr0FLrtj0cSDKyhlmW6CqPvF1XJK35TGVSexMMk0kb9
6eeBM9xx1Amj+fO1iuDtOBEYf0C87OQOIyXYoB5Hzo9zbLu+LtzsjCrTWA62Q8iO
N/w835d7dDclm9fl0fASMETGGFtMLNOIf+8fDPXLL6BKLrveunv78c8oCNHHbx4y
yMQg2WRD3X0OdTqOnCGg/YqUHYaUg2tRgzB58/6qNQuqLWTd458eo7XYJtr14sOH
/p7kUvmxvUMrHLUfS9b9NSoFXW1uxvdATiwKslzRNEEIGaBTEYZgyKBFfgp380/e
DgB/6Z18KUsVBrhx35FQfIAVDR78vpIcFE8BXBoq++2IGdthe/qCut2n3yk/obYY
vUbrzKs49IHJk1Zpz7VP3K53t9WjhG+PI6LciYFKtong1AwyvNqcAiPsXSMNdpf0
zu/T4HjVIc6uyHp06oTGh1E5HmcMbz/cQ2SXnhmxbg//OfU+0BWp/7gIB0pkqVag
C6Ezkxpsx1sCHUQxKGHpn4bOKB0KnwuboicP+gbm+4uJuGTGeaIBzWbDELRcVvsU
1504My8cKKRXEhVonmy5iHxIERvaq51sBTVovLPW3HdCEMZ4gtL0VIiGavSxRUN2
IPk7btbomHdE6YjFBPMDgTkvp2rUmx1/bJS/SvffRMpKAw1kV1Ef3x1mFEV4mSOf
/AOOOb5DbaqLSCZ0S9RF0zndjKVVwWpW0L2mCqja57V7nMQExXrYMlyzdmmEstmU
UnyxRfE8sx3xIAqdR1KWhO7+ylHvOgyFMOmD0oFfC9I=
`protect END_PROTECTED
