`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+TSgkCpny6ALQH65mCFsm3ZEnkKGXoNJumD/bSK/+pwdbqR3Xjzd3es3pjjWlSjv
mHxFtd3HejxtdYeimMQ94ENixR+BQxmr/JsCMkSPUGahu5R+CuEoP5cZWqnzmQxO
SVY31+Jyd+ZFuzskMGzVeyyh3ufcnd+qijnRXIVnPO6Qg3KC/HtEiARCkAz2Mcwj
YnTZMqaUb956xn8FF5Al0dKKD/wP5ZR9IrI042mxGRYIv7wUdLzdMWIwlcvB/5NU
jME0xhG3L+jS3dJobIEjbWtwtKz8wE/ifWI59JsPw0r3x+BbE8qUNYaVZambhArI
NWyFuWb0EsoTUJGgC8yNvhxvBtlH2WlmvZgMAKdP3Zo/daHsra+8rDpUsQu88ZLa
Xo4xGpJZC4+4NVY2oznXwA2wwRs9WZ3NNqE6OYEkwCtyghgS/Nik01Cdd4FUjOJQ
YTR5jXlRhNMbGvdxZm2I7YXj1VVT5MOzTq6A/9QZYpw=
`protect END_PROTECTED
