`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
imxxomGqajSLyCECh1XSuwoqOufDWh1A0zq7abvRqmpVO7pNnqHgdNPe3TguRaEQ
xQOtWx2oZaa+Ixeu9x6zyymJ8+bKxJ47XKAFK0ua8FPBxctjdJcUgfUxpSru5yuy
uNZso3TpbmGasJ5aH/A5eMFY/GBFvdXn8amxLd0wVsXHcsXZdAbAgMSvzRbbMwK5
/jWpw3kACh0j91/VStEN3o/OVKFWyRkNRoovVjXp9yEoFhTYBaI5j/b/a6+ufe+Y
YtZMeBWjr1xKMpQiif7G3We83vgK3dgpq2tmPmpwSMOzIpWfZKHNTxT1/ccchqqW
C1NgniXSD/fGTM4s/GHAIce2hhws0lPiNA7vDBynsww8bA3JbUgpE1Wv0Jb/sh2z
Sxsp6To8EkfgvKiYjQonOOcRKZbR0ty3tKu4hPL9aykhAAtvO4jRZ3Cirx/UDgwA
0Dv8Ui5MPyDzN2mbVX35PybFDTj0MvN2cupl3Scl4X7pjW/bNoR/h7PTdqk54DRI
cP7srUEMqihbHHiQjOjhiF9NzdjShtmwuA7g6UCqCFuLP1Us31YS33Xw251im5d6
oN2jyo66q2eCtfxF6Udv1BUjWUo2dsI/ecYZLFltMfuo1iiWLt2+Hwb3tj1kf46Z
Wl5lhlntSIu55azny6YdXmpiECXJPgILziGieoqYXzzrX0jxsYfIO0bhqiVF9tE4
rN+ded/S8GtN81XV2NNQjQH6oZsb25ZCjseNyv8aS1uQpZde3y2QeokBLFk8hCD/
Jxm6m1oHexkPRtahUdv8R7HnDLEzLs9n2qmZENitSVVjlPDuZMt2bgnnPtpezMzp
ZfKlIS5wbde8FBweI3CPBMWWlDwBsTAky3MzjXIy84OkbjhgoAfCCQBYYMkGc8hn
VNHKhoI+haiL7TkEsw5dHFGyS68rgqtKmClaKgOV8g82nW6OV68OeadjSEdwn+b9
YafCzoajJZdpQ2PVFRvFp97ZW+7FOWMORhDKRKQo85JZPXl8phllSe1x9Ta462hZ
ck2cVWUdb/BiasjyWd2xwAV2OSsW6JWkyTsxMuuKwSo=
`protect END_PROTECTED
