`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1/YXYZbpOI3PJqBUIdBe/rB/nNtDiEQXUYlGnJc2oL0RzIbloL0yzRGe5niRcDR
jtkqUxKtpcxaLHs/yoLJSR9ZbYFUm9lwMoRxWiy75j+tR7xiUqL6fNc6XKEY1+7d
JtC9rTu5IQ42MfjBPRlVbyol1lJQ4enHe+YNeSMMpMzvd7OO1PVoPSNJq2NpBBob
WbVhvENueGUDzVcWih8F2x5UeIcUNk36U0zYGPRHZk6pRZeZMPhs/I9CCxCamnmL
cupT2IGa5zHyVPCY0eAJ3F0NgzFTb/gMqgZ2RaWWhxhnUHeKsEbVPJAC43ROMKhD
j5Gzecu9IDoAyll7X56RnbKYKHa/Woe949bk18HXzWhbUdDYwrWpZ20eFRxgkyGp
/LiZhMcCSpEV7ZwwgpJUrYq8Lw0xKDR2rm7uxAcDBIs+9OO2pTDLqRnZmAq9hwCc
MOcrLAbxADMUCGBQPol1NTvYoT5pFQZow/hIvP3jRBba6aarXG9TaD+f85xJUA4S
8n3G7SqbTxw+RFg5JX3DjhDNX1MkQxRPAVt2I/L5p0s3tMSpHu7VVPGnhrgeBQzu
lduUUM7i8ZVVDbI03VVAG0Q7lC+my940qsGM9Jj8JFO/da++QSvX725qfs0MT82f
9EFIZh9c9yPPJRhImV61uedky3eJi8D3xYY/RHRcE7LVSEYrvaBfTC9ZpXv7VVd9
3SuJx+XF2GfreAFQQL32M4lmAFRbiIfWVH4fLGzC64J3T9A/QztymWHAb2Y2etDt
tMTpzSP9Q6zhgtypyB76ZeE52RWVGe9vUflkUBn3WekRvM89kAgOn9QwiPG2ifB8
o4PseLhofsqAYPJeKkZNoT4+wiw14HjxcAXH99ImBSdvunqPvtzQLm4hebETfnqD
9Bo3GM1XW8JVEmB5hFr62SlLAcLQ8xliDtY4/4dKuRYVzWrXvDICncqozZvWiRFV
yImTQYB7hrj1C461P35+gveExG6FrOg9NLXXWjGvgxfp74NTFQZGODyMzX+7HITK
1X55+9kTXiWiuBMsUUvUTPkq/AFPZgH2EDKeSwBYdetvywGEgwFELA3DhG7szvv3
73gfKDP156IljBSJ4z0HDNPJnEWOHz9TvQFFfB3m+grAtRYng3u/Kqm1cfo4FkWH
awBf/96syOBSL67Md5IUcmkZB++a1MU3qJ+KEKeimUyKRSRePFEyVizyIa5w1nr8
OAIO49szJV4DBY3Feio+mVfv1+99Bxt4mp+Zw6goN/eUKYEL9ML9ihsSoW7U5Mjr
x88yIgqhN+HZrG4BAVaW+46LE2BCOx4KeRuSgWVACueLdtLU3348jUGvVN7nTUlq
4ejrq3CRQtV2nffpiTewmv1aOGsgTZ/GiuhEiSnX+8tCOLOfhRM7jHLpU+QrL/Tj
7RD2PGYPNbIdfgQGiiLFzH195f+GM8nEf1tu0s75g1RaaLG0k0K9Znh0WgyIR2Gk
JfswSBFdjiK5xzkR4CMKwNheALmX2oMN2JRoDeXhGAIbH8IYYYdpaCZnSPclkCyN
WcLhh2l8T3EBvIETS2ByKquSo+G8i4Nr/95GblhCBjcprUGdU++lNND+vrmi6Tfy
sY5BrG5oovR3lOFmUw/aOi/DMItOtMpZ0KHoItc+46qtNKwAwzrfx6CMiA6ADl7/
tQ8E/1VQuPW+lIZqaPidE6VQyquBSxJ1BonMUH6HK+rdBfmgcDGMHgxdzZnF/Nys
z53OIXzacBDN+13ma9UkMOEkDYmktE74l49AR5Ctcemq33Q7OFHh7bimH6tsd9kG
eOa+IlkRs+jVINa/WR5vMNLFwHHStVmKRtrYf15J5lpirJTN8cX2BhVLWAJLdm7O
rARQfMJqWcIhP8PkCNS1sWnUvDJjN3d4EpQ5Txltocw=
`protect END_PROTECTED
