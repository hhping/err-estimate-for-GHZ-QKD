`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oE/ind433aFMRN6ONhVVtF42ZlBq0xxgh5QCG7qkjllKftGnShrD7DfvFMFwyeDV
fwmfbyYfvq4YF5+2zOTHzRlVIIJNFzDYequYpjZdYMHwcSqfmXBd+iqDbKD7xfSS
1SLiiK0URih8L8QfWVC7riAleZ0UlkFHxPTZ49HX9ZPic111vCdk0uDvMQRk2gSl
sQTNZbtubcBcNZpuJsBTy4MO68KOLHZvIpoKdi9slvGyLzcYVwPVKY91gpjjFYPF
6qjqIKtHYvim4AkgAQTAR5YbgwCsHTAYZUN4gN1YMcpyCmwKj4Zsq+gziFjr1NkZ
iH2ThS/Waa76QQyDaCNfwmQwOn7NtIyv1NwI7REFu/eJuW9lpHRR8bSRcOS6+VAY
U+sMNc9RFZEz5+jrMca8njONIJrTcylPSrbrRs7HHQkcxS/cCJTytT29qusaESf4
ZeAhl8j5vRq+146ZVOUt9fRfS1D2NAATV3R8bMrxUJailhyYyUq8SSfyP68hMRAv
VM6IRy62lgE3zeLr1WYE8X9u4Qy1ffNkCQAs+V3JC0GNdBavZeh47V3AmV38skhQ
+6UdNmPvsxnWXcVMIQO5R6Ajgn6fgGQ3npGGuptvxVlNzJQJ/Liw52SQPH4/aCSU
r36jnNUZQXwPOJWKGEqg6oY6pHv62j2/YATATU9KCQeZjmcPHTERkRR+kV5p80IS
Tvpcw065/wdDXU1lOPDTiyRkx8jQQFt8D8s2iRwGy4Nr5SVsPxe7rTwiASav5iEx
QBlYFO8OBZ8uehGysg8w9CxZdz0BV+6fW4RBiTEKNfoMi+SX289l3G1ilVWMVDPi
naQyKWTCkZA7y1zn909NrN/1wdQhDH3HY7ut7ojXykGkIJpZX8ABuGSU5Zyfbx/K
5wGWyUH7lJX8QlW2hcqOPvqChGYJ8gca9/aG1Cf6zOGfae6YlSJIRu5r/rOzu/Lg
tvKgzxvAmBPihOQ6LKSAc7yENSwkMID7ntnRqwEHqAdat4ftMKWl9rFhOoo6c3qs
uINjmhPVoZ05Cw8mm+MThxDUyWgDHDeMm9F9g1G6PoRHXJSNoUEDh6O3mhSU9R8y
GRGjxxr22MyDrEyKWoHrGSPRDhz1dRX3FLa7esEEvI8Y+QYzn5Yhf8h8lC8FXdTo
yUWF8jT+9el1LKtGmP/O1Z5bCWfUqVpnG8dVAGxnlXg6MJNf0s/UIjDcEwaTPlPW
LIAkeQ8orqGq9e4fD+yI6YrOchcCRa9UK4EQyW6BOzVl1Fbjf2hESJwVC5pn3suM
RSxG1oUYQOVJCLg2L0Kv/L4sqx041zBP68hIhs62RKRbg/lP+wDsCdgHu1bfFhvP
W3Uh5nku1bWYlNuLpmMcKcx48+LhyiMLNoKWfBwRT/oW+ZtEPzrOUGlH6i5zNMXb
Yt4YsEoU2gBvwdYbqdtIa4eykbe7SZ2Pztxu76Q8Fz+78EwsqRp0gehGuxZDS4r/
C5j+Rm3BK/EhQE3y08RlBmm9gvmKQJo3WHht9OtftbZ77Vudrge2v3JMEQdF1ugN
+iaTx2fOA+AS+TP5Tl2cXThD0LYZ9XZzwxMmHABx4w2/2bTu+FhT7Lf9vpuQN+01
8aY4v7vEhoxwWu+efTjn+28qHykBKoWxfTIm//QHm/hjP+AzqZ4uFYRhB3Tp5hXi
yFcSfn1kU6rlSZEEvBkjxq6FOsbgitewsfcs/KC5QZh/kngbbIM5EiPbpNe2SVQi
MxngxYdwj3mWdhD84TQHTTD4hibAAoYaZDIqa/b2wQvdollO4iXYRHpWe1RaEjnr
i6ew9S9uSVgTr6+vFydy0VmpicrMs5/Y3ZeyH+P3p3pRTnYdw6Ib+9P+d4YS9e85
pm60MjPog753qF7TEgx1nPEJ0DlMQXnIvWBmXTgeg1JjLMDIn+hvAGTefOfvHMmZ
vojioi2eRB/MOzeoyUa3cApoIDsJnh040MkPyFR/R2UT5etc8X9XT+VsoeHC40qy
g/Qa8qOCpEXpeuKC4bACU77etuwmjgSQs00BGzcfblEhREGxzaCaKKSqeTy7c3QV
73NiU6i5LD8PVBDSR/2BW4/wj3sjAjkuefbJUZnG/GJQNWre2aOtJQWo7gi8KDUC
qdoDNlwEHE2VWQn8WcQtcI6eSHrIPwmQtpErl1jJa0aPwTy3Jsa0Il6b3p6+RGDL
eGM8vG8BY5PiHCAxIPUVwN4MQqzN1zutLmxn4irF4DNBJ69xEAvbiTPY8GIrCIwb
vSe6nIaL11mn9wLTFy6LmFrMiamDCRTfEyBKEmWlwhOZn90vLWCH/CXG5+t7zk/v
2HMvyD8UHuL2QK0+iBfU53+qvKxdBJcpwqfR5lpiEc0RCV96VMpq9KnHhJdSDeur
3LW5Gh094/PV3yf67r1ZoAmGq8/tDQoqXjx/ZCrxhZzL54m0t4k7FrjX6nHNSx/r
2NI+rN5XfNOr9cvykDfx6h1yOuXS/6HeTNlrFx4IHRbIIBbbAz0xK7qr+UK0G2YI
ErXLt7Arz7fqUXzxlrgcJof2CQaxbvfs+7XHnVD7Ilp0hads+K5BVivaNqjTZ8Fj
rk6L8jumY5z764wuSp1oa0uDbPCz6BIGZ57fdip/xJDQ3Ylcmc5y112R7LSn1Lfv
sso9VQIFA621MuTCva3/u16EWltIajpcm8kt6PIWYB9UE4ZY43RyGVtz/o1LKWaU
gWn/HT3U/E0zw4WsaCOPj240g1sk+7Xa5BZShp2GS+tfPgu2fMLMi6xJ6Z/DNtgK
ICPfO+jokSIYBBG5CMhMKYxaOCSp2D7BKmZaocsawIL+bJRNXoqe0OhQVoA8B362
7TtDl4PdFkg93RnHkUGMFox/bBgGeSnE7n9komdjFJXwWX30iknAFLUTzpooZGp6
hdiQI0BQIHVoab/waOQioLfCL8GMjQj22Qfq6LhplsUObanJ/iwyYR+7wVPWavkK
rOliCInaKm1U9KjvNA35ODplOUdBGfdW8auDU+KZhyx17rru1V2LUgEqvV/7cBlP
FQgRPAqu4KH+CLXXXqp3j5eJsxW1IOtH859IzXVUO9fmCMmz8c0R+gnRZgLQyPEj
5jxmw95ecCnocBGXEW1MpfYrya1BUhbLgXQQVGrO/7U9HxxC7aj8OdxY/npBUps6
t9/301ftvgWrEXFQTgL8OxiYBVISrV5GAj5q7M3m7kfC+3w7wWaMel8SlXpNNa1S
DVHSFbXLfWWF0ZYbHYNEkzx0H55+lXnLzDQbfZJzsHPXU0QnK9zL1NP7qcd546sI
OtCJsYJNkY7+ikWA1L5lmKer9EJoqQw87i9O1XJN8VQtWmpfLWZ2SjtNA0wutWd2
3lGNhrOwH8Wh7KGcIjUn5eiorttUprqj04R9NnU3ajoERFxN6aNQCEpeADtrQwkb
v22CCOtBEa0THoku8YaiWhoxLG3mqnHrjx2ARckcSsojealJX9q9hoIoBkplJZFr
9woC6Bx+3RNmFhNz9EBaY8lEOInmCR4GlvGZogBofEGZpmhh/4PUhGsxI+SVQier
UohUkfWZryacjCZqud1LG9/Iah+cZ6ysQRs4xE++9E5OKng7ndoWbllxQCXl/HII
dsojKsEaa92+xNf0Q+wqQTeP6MpuCz2wDlkGC4iEhTx2kNUZnpSXwG6wtUoLq8E8
gic/VKSd1Q41FIO5dLlXElyDAB0bv3UMjL9/TQIhp76mFqD2Uz27CQSDNeK5DLbd
M9l6DetjqCMlxLtANm7gsMflpmMfVMP0F3P0qiZ9gra1Pc7pbo5jW0W0jAIJzq1p
F041Sc/b1K7rOhuxSVWaidI1nOIaka6VqQFLPovkP0OCqg8av+YpLr3HC8d4NRy6
GB3eD2yhfgwW3q3WcKlyRPRJ0yO0WLosPZOq3M0b5hCqy79yyieUrKHeFLmPtC2R
GPiteX8x9NZW3ty/6uie2V+kbWPF9tMYUF2DAFVtvPPElZfK8derJxqzrRKvBq8b
O+TMm9h5y81uViwt2WsYR9hLbwQR+/x2LPGuI2sady9Ckbe+qaVXNJTGIVKTyWX8
TSjHbii5N6E6+k5AHQ8Zki+NmEdKNtVX1OPsYcfPFK3V3u1jRCPZV1Z7pg5/pA0X
1WSDU/nKFOsaARqll5SIwYOADKAqqZB6YaQEI0NOZtZsv98X/3kZnKxRWfLeL8w2
gnrk23pBMRTjxnIBq1CzCCrk+gdeRsNFcVj+Ukm3VZNPaKbteeSQF8wfjQxH1eLg
Xr9AXf3G2mtCFHXaglmknqtfNQFOEDkzYG0sCpEUDimi1cviARcxr2yGeJ8v7rrb
AmIAvyRc6Ob+FiHlCBEPkPos8RiC5iuXPAQqYm0QXY4GPPa4RvpgkyK/Gtz4wpNA
uzaMwvwjeVJUP/csVLUFM+ffdQVnsZHRhFX/5rflOHJ6kIHH4JJ/F0QQcPw/fGYb
ZSijX8e7TV3vy8YHt3HMkWOiPEIDnuP4Pjn1rYEX31fXgzruLhziVU0aX+X+Kx2e
n0HdsIIB0Acz4U6nF7mZYk1HgmB25/rXZ0oEuCxcdt//sv5r6pBZyPznLES8HBtP
sdDn7unHsddXrlPW6a0yTY0iAKmCJ8+1ybX8JK4SJtYmB2AhIzp74B9xPF1WyEAo
igdjRfGeLN0Sk9xTn1hhk5Rvp8TtLFY/DvnBCJMezpM4b0uLwy0fAOMPebKk8NFm
ssaWPDx5LxGoGjlzG2ptFLt6918MnI7y6dwS1eAM6kaqBbTKDAeWVTFfy0yua7yL
/+M3jMfU5sfeGssHnx/YRewUKxlnjrfDZnoKu0t9VvZ23btyGgtoFlVBoAq/6P85
z5Z66kId1E2IjJGo0DDO1nWgwgK5RQ/9kuAjQWJIjJYtvdBaeJQGS9f8pXiQJdc2
mfYTwH5i16yekvwDyFfuc8gftheq3DukMDEMZvhY2zppGpmBANRsUreDbs/rtLE0
aGJycVxFQcuYOVpyPFVeHbnX+lNN0O0+MZfsQGMPrt+TGxW3CjuyEdkORPzpdvM4
ChN7UKNNHeoarVMf3S5/+UzMXbgzvWZOOfzSSykzpPa2hzg2+g+9jm36mhfYosWR
msSQAq1Ag8tj9aEYmZ1IkygIvGxthBOf0WpILDmbhB/qUcj4yvGEx8ewNHId5bTb
OXm0POs+bOZ5k+6SAlEY6JVnDr9VdZJPUBohOf82zFXIFSwT7XRnoVdqYcmuMcrU
gLuz+vC3vIEzF6EjaFBQbdH9VhqyLVnnKzAOHlqdxepD7+0gK3Q8MAcDGJn6pfLO
IRVIk/kDT9FpV8Djk0U/DEscxfofKM0M5/fNoh/NKFmxUlAOou3FROAVg0Rs3tYl
n/w5fLBmhQt3gdoab178Q/MEJF99YLVAxCaPMctlBU/GhnmGfL/O3CC2dkDcmjaz
YEAjHgzPdIvMpD3l+sYj3pi8lVAfXrOZk5bEX7MReW2vlxEaUEKIfPf2cDzYHTxt
Kfg82ZN5Hui8/tGGjy89K//9waL8rY/Ny6xHwG7Tb9ubcuS/KEAycSqCgyB0Fjfx
kcjOjXsz2XVYsFxijRZTBXnGNL+bhs0tCu4ka48jM/Y+eimXRwX8iUAgq6tOOzpt
vGEUt3SCBX66DcDk/U9g8XelS/UMgNL6YEns89GRv8ZY3ixMhwbmV294h9xoZ5lm
3DDiuuxdte/sVV8cXZGbstCl9bBU9OYxKmMKOyXm3iCR7+qf0mwF/E1AjrWELW9R
H2+qeKNynIeu0ZJjvEN05fSeLt3fj3Sgc/vhbBFDeu5i6EmTMuLlw6JhVJfBRSQI
MngHtjSiQ7Oijj/c2EtDaoNgPSQlP9bhNVZ5pH67PdR/Ax8wv6sKeX6sC4ETc3gQ
5e3swcOMOtN6Ny2CkFIxNqHe4ZqP7Wm7UBDBfyX+lt2MF5ajKPIHdEy5m7q5ju4M
lPLCiRxsp+3guIyVwiMN+mcv/zGYVvK+TW38t76r9saO3G4YvaDGexuZlj2j7b0k
L3RluqvZ0lZCe2Cg3qr11rVXIz5aqXFAMBzpNUcrtTQe2n7rRCwOp9wpISvJCtwz
O0WEOkM3Vt4GMZ/d2DL/eUe0wliR6u1lmD5xOKUj7wM/+yYIRsxoJ/ywMIpdy1Oj
DYuJEteH/9h7w0q7eS72r3iOeYCiF278SFi6ASSO3s3YBnlHZGIa3bDnIgjIvmES
WYLAEzMtF8wbJRU9IO9L8A70KcpJgY57jL1hGY4wi9tDUbiM+WEpKJ31X5JuPaTO
S4ZhhClORGq65nDvAPomPKGpzLoRe0Uqv+A9YhGPMJfa4/tlLX8uHVvP24Y4Bkem
Qt/b8gdCSQUGc0/ZRX81bMUiBfpbJ95HQGqVnFAtEINhePm178fx5TkVgx6xzr0D
LsE+oCP9Uwq2gWYpUBwl99KNnVak2rH9lRQ3JpZ9DsPPQKjX/Vt3bxsrYH3lm+SK
s9zI0nNfVhaF1C9qE0JChtCuaKwpz83cEJogmhILTOqswPdEcYURGBRMVxLwCnH7
xx7BE3GP7XapldQjXasxk36XH9l7SGL0G1F9XhzB+wHMCzaetJW0yp98aqvCwnj0
6scI2GZ7paOdLetFCz/eWzadzDFZthlY687k6alTjawxUcLPzGGxcOUw4S3L/hbY
4DdE1NZogXWKsgw4bm9vgzVPcey52UDP/ogqbW6Flg+ptxO4jGvITtTDtFujXG+m
26/GxxXPHKxrBBCrQriypQ1LuBbVs1K5tyNsNGD7VX52EZwdKN8L+2cPs/rUyQet
HnUtS8l2z/w8Sig88zAD1MO0tErB6vj0CAsYEcHw537tHxmnc9fK0pcmRZ5C0Uqj
Ohtge/wjwreHOwCSEb6p3k+n4r4Ga7nQWxFgjflbtcI8O/gn+GEJKutHgEJgHVj2
AFMLoiCKNfo1tQJlfpbE5mOJA9bML3j0eHT7nbiJiJMi/3fjmVOlR8McFbRADCvk
D0aHhk0WX7NmVPHbSX8CL30ivXZ+G/9fiTfg9QMlzko0hqhL/+GTGk6BxQOnkv2X
EvzDaK7anjIPKBZKviZRVStYGawdeHnc3UcWzJOpQexxwr9eUHCob0d8ANM7lRd9
xsZCotehlQ1tIo0jBVS3U52YF5mnfsuQmXDWOFzBOlYeMyS8kzUha6on4Gfz0wke
zQm/y5WQESq5E9RS0t6CM1+j7QxYFEx6yUYPzgK9tU2oeZXvDyUJSAWRZ6tn53Qz
7MPJ9SLTN2Hn1/OPZsDqYQfB8UNrNn2Yv2OczUE29LgWuiEQtLPJi8kDgFGbwCkc
ZbMoz7oQ9IqUG7GkSOhFx+i94ykD4d9FbE/uvB+USiS5LhYJ62tyDCzETQapSCnQ
ikYfyM2iMjOv9nAKja4NRJ5OodFtB5avEx3Wpt4aiFdXb1r/hkOX7u+qAbJ6o+oU
ztkfaEQJgZcIAxruUxejtuPxnDcJszHd+UvcqxM6SEnIcGCWZG+Ke5irSWyanbb1
veQjsHLFq8UG1Nqnc6wJ6kLKpHZulsVAMbelYgZtiXL5L3SOmHh9OkvpWhxb9Ywn
yTCnbbcrffEJLUv7jYfERfb36TR+qtq+7L8NCiD/03GscEjQf7R2tE/UhPdl4gJm
D1MzEwtJyPAgJZRFzx/RclWqWT2UPYKkLopILm0+e26ohHyGZV4NziqyQPaQQOKy
XdXTl5oXp3zuTvHiB19b90VVSkoNhR45C3rOtNYONsvtyLWagJcSBi01Kk+nAjiG
xaFviGaCIPHK5qUfebFejQp1MSyLzf71XYe4lkh4P6hdwjcVdqGSCmmLOGj6lBrP
A00pgkBOKevXdAauvG/9ynQDZT09oPzqRNOpBE2ScOxA0TS0Vyu5gy9Xw+cHSDTO
GDL2eqL9j4+TJ1jaA6cfjZY2Qwvm4YXH831bgYISjfBsKlm3tUI6hFIF8v7hY3Bc
fA5aM+seoUVcssRqbHTLS5HmVLjGd5O9nLQ5nuwNMZcO5JEpYrh2R8S8Z4Uho5D5
Se5Mf9Rpopslhwl9cAQFIKN+kO7l6SJefDymGa63kGZzTnBnIldOBsv2qCgBrcpL
sDR749fBG1De4axsMnMbnUoqzlZurMQdVQES0Wt8DHVlLbJMa7RbvbueVkH+5/jZ
o5QlcRLNvzXV4I3OpOiaH5uokJnIhTaPZyLJPTDA5fVOvhXP+K1RbgBMI+l/CG51
Bshr+GKIZJrnrYlcacsShuUwJYLhjdzuLKGr7tkDUNqSa6pUsisk82GtHOG6fqfM
GHN3gsUPDvVPqwTUYKBBEn3z4xjciGXTFbZPOzgV5zVtZ+7Q6ey65h8pMnA2uBBj
86bzziCbce+rIByLQRWJjEibWG0cSMmugybU8eQRFAvx1zQQQmNJoyRRnk6bd7UY
rdum79v7nRyvJcfEqJBxpsw79B9Xo2Yeq+JKniA6WbVdGk6SsltX/r0vU7k0ivns
ft+zk/qYbtQuQPrxwl26b/3fj9gl9iMdpbsqJgllzTxBzua18w6T4Zvej86+PrHl
s/saV/EVzWHJiu9KVwFBvj6FQlRa0IsvTt4vLrvNeyraHVH+OfAhDuowZUvCQe4L
8twteP751noS6D43KwM7ylFfLes/kGcwZBUSmkEtQz6WemRhOU/ROMF36BKJx+OU
A/9SQ+kcSg6m8b94G9kDG1gv52QUTjfiFGEwRfnabfbHnzB5nUN0QMgv3G/AkR40
CZk/yLAtwAYDOEEnqxRUm0P7IsnHCL/UdSksbPOp/+s2DG0NLFA1aGkuQ5NszCYs
qw2LJfj44ZmDrTTPYxh5Ll1GZI6arF0BA3dpnLOVAX7L9cvQAv2Vp15prK1M6XVQ
3kber6esUq2YRg01H3jvCEb83GyHSpBBba6faxCyLpqAJ1MewMNBEcxkFZtURW5u
MZt8y+QEHxyo6yw66vMFiZ6FVHJv+yikwgs65M89rSB4Yc+TNn26H/o3tr2iNoAv
1FKZ4TDZLPI6t59q7coq7sZ45WdpyIPyrFe37K8BvjpW8+LQF6X9wETGHDCt2kvx
zizndUpM6Zxon4L0RhzG4ujiEdaT/+EgZnX/seIeydHMdFCf+MJWg6dJn2SBD9De
Ej+JQrIG4RKzgjTpkxnt/dgGRbxnPNJgC7NCMI3pv0122Wt4NfvTO9b2qr9STYDq
b0OnB1xpun3nmSqtsuNE46IUoJbZdfaWF6tQsysO8MsNk0IAaNpJ4p9PWp7Ts2KU
6dQZOPryQhDy0BYD41m/SFhsmmAseRAxycdGPhDrGrqR467sPLBnMUccumP6bFfY
2oaOHJJ1HlLspsgo/B/CXQ7PF5xqnp1gGCAw8gGhN9OcSRNBvlSBpHylImzOmxXY
gASNAqHes9XQiwekYs9uW0/Lxhq58uQmJLmVGuBl2hAI4YKS8nkHVXwZhr5iIjUW
CmsoZbxwENwI4YdUPonilNxIeOvU2NOBRl7FWWcpIFtBe86uQ/Uz9WHDf656HI1P
0LYwTa/sGY3Nttm5wCGvzT3dTGyJAYcg+GQ6/HvG4kyRaBEIyMh92qH20BneP9wk
qiG0kbG+wqTjk/mpf5+/86UDc7G1T04YAWjYQqqNY1P3Kuslo0ghLxpMhvv3Kw2o
PPDVBSfL/Sd+J6zwdQu+F7ZrY3uibLDFIIvWyT9eLc9STIqQTIYmeRCT0MzomYth
gTF3wiBt6Cc0S1pVEun1MD6epvwmxCwV5oajNV7OqSxCpoHfibfBbP9EDgqtQwv8
HguEKnz03jxdquS7Kk+AXmAY/ntju/GZJ5/OMxzHM0bWBw3q1R2cYnUdGNRAmVYe
e5LjMGqv2CIRzE81JuNEWSlF01kruuXmD+QWYLO/mlJ6tpg+K0l11uVVN0wS9i1N
BxEUMPaEabN8CpByl10t0wJ4N3f8GdnJDdylXOBoqRmznJgahMzCgBHZn4OvyQ41
Mov+11iNGFEeC+5+/el+qItLHVwp6H/TMyLjGvYSx+N6Hdfan45tnTyEmsPRvrK2
kuLAFROXBDlumRicJFYyDoJwz4JbmKV5fGZVu08Hid43HkwgfBmXJhZ/0llGSQWe
xX0TWKTs1deS9sI5KGZfe3lkBN8ZCwzDTBuxi4mRYqIFUGEsn2ovn7VvjeFxB/2g
FDbk+6tTN8jXskvgpt8OLURo5WmODxot1AbiHsVrVz/ZzpSereoiNLdPMt5sjpzf
64u7qDdX67cxYmQOrYJtnJ/U4BhAmLvTgOQscdy3o4h56j/oN0fK4aaLbEDi2s4X
WIf4zZ+WEi2X/emKuiKhTY9SP7bJrjBDOzFeIuYmbxNsPnNsRi8RMNfA3o9OwRAH
+sNqkoGAOI1rDAkmWJ8RTB6KRbPYDDygVCL38BEMcis04Dz3bPRBlZpqIalUqT9f
TCWxyhb3Vvsw7o+EtBgRUCbOuyjZ8LHsr9aEe15/mKtV6A1ak1HsWhTbcLTUnA4V
tQYY+5Ro7AHaCjiTnxCBbS3lvyzB1oNRoB5as8qHcI9/zmAK/3ps5io85hl6gRTF
zTf6Y3kkeJ6NNLfNLOBbdWo9RxJBb1SSGqFJBr8spXIN/tWwfhwXES+GwqMiYpPz
E3Uq2YXRvmhvSrjLB2ahz8mHVNjeeF9cyL2IB/uxqVIPe1V33pUIzwWN3JQ24APp
bpxnSRs24+TLCksw4DU2EYTia0HZJBTDzqIq6bNlSLIN/mMxtJEqZb8CXTATdz7D
E77iJUzbYrad8FC39RPIo211CVomJJYILQD6rwc6lvjw/e1T6dKNo2NiyhlYtyzk
nS0Y+HTlamoxbxEMBSSbn0do18py1N1E0uu4rd+IwtrJJeGPmmbXVfm8ONDkyhep
ks2wX9r2XvN/JPKhxQrAt3OuHdeRr/u8hak2kF1d3NOMY3vj0udV8DpUoqTEzNkk
EFpHMUoByn/M1nHhmE5Comrsv5DwEtSJH5m3oPSJDNaNaz7G+qiTKlfSxupwHa4e
Sr3XPNWaGp+N2HMobHnvI8C4QcwnoO9o8ofLnzAiiftUViNI9ucXScfFNbdrD18f
fpYyegHj2qk2nEk9YH0xXswgVcX/emWdQLD9nTm9XDAsNFpK3e8YC8d+qYEtdoKr
uSAw5a3clD4tq7OHqYoxzVuqbMuM2pmoZdaQyNZx9Oy5+DlHciulIaUjxemadVAl
tdeQEQvrq3bQiwpb6QpEfNYiQK1RsAOZbv6BFaIkPQTEUPk6vUPoX2566wkzbd65
LoiAWRASIx7h+ri/tEnEO7ROZWJHtxCfboWBA5vBJGKcndJsLHfJke1lEx0grUzv
1k1wdRl+sw/uY04sycgyDTKgdk19nyrrGW87Q+GCKM9BZ2quOGuD+yUIM6CbBsXy
fuSgA6OXWg7CbT6thLkAEosmef0LlEYtooj2eb8ZRzmmFrYOuL5D+z2p8vCUwSl6
PiBYS/fCO9DZTOYsCN7HRv6ukH3Coq2P6DSiIrSxYkbT4f/NE5Fb2pXP4CWnw0eL
eqM629n6cpZ+Vgor9vQnv/+jsU+k7jh7limSOJEuuisb1CVDUxeU8oNT+FXUbJv9
jPJJ+BWB21CoAP9zRjXcp9BqoAJJQDkpjeQJYbmQ3exF3htrYesc6gDqIEHUTjJQ
dLugI+dlkM04pQph0a/TARmEGGYFV4rGmtM6b91UdC1rQ8/vPP1m2+JnmP/j2LUS
nTJGwWJ8062/YrYOvyJ4JvfpZYP39t4jtPPQaAvAkrAKZrH8OSUQhyK3kdijRYXC
FzXTv650Wu2XjUBuRr9e6PVPgPK6sFQnpkilZJR7hT+uNA1wCT/DmrVsEMfCy6aQ
EQg2PL/cwwqVLVb87iyIOEjcb0tsMjgEIWt+iRCPIEEaPetBGkO+5BrhM+ydaIVj
nhRhhxagxKT6ZzQh3rv7p1r6d9kfvJY2oEsty6SQcLd75XWeWwbQDL2WXz6FKRJv
5xYFs8pWNR6PgQknDWv4jjrNbR5FyV4MOnZo2VcwFB+ke1CJoRc0mo0BI8KWyGrm
QVzpphuVmyPMjKRdAnfTTDMgafca/bh/cASgmmafBbVVDUnotGjRqhQ9s7LCCxh1
kDoT/bJ6piGjEVKDN/A8eKR+w2rnmGYU2Ky9xymXjJcV5X6eSeE2nsCc8KTHvdSt
QYvutf1qLhgbylxStbOSSkrP0rDR7X7uP8FsVtMDqwqXScWZPk/ht7EzepJasaxr
tNLm7u/B0r6WawObjAZgE3Ky/exTcURa01TibFz91Im3UIZs95eyRRhVw9TrAdmN
AgjwfU1eb1yLPrNvr9SForU3AtM/wpCbhpg0s52ZUv5Q9qcx6B37+HgFx6bz3ajZ
l+kjPDawfbTJKQYf5jbGVGD0XAA15Hm39mkGbYEedn+XstArT36cxZkWxQ3tcHuD
NqvhpTE2NhJyq//+Oh48Kxt3ia0q2wpHaBp6aGjq8584YgA4YxfBz3dQ7IzC6DL8
N6tKcQyAvGsoLEP7dV3rTZs2y/rfgmq6FsaCTn016a+w7r0kLLNXq3SmxAN4PugF
PCFqGFi/Niu2EwAFcIRO2tqM5Nn3d1EqZ4IcR6LQ7gEsD/ZLheVPoVBBscPoG4Dm
pI6y2ksUjmVrAh1Vdv4XSJ4I8GxAWJvT4K5JifF9YFCy6wmwr7qd5KlFFbU36Mfc
I/KUVbzTUHeD/pu5OAGG7Tw1KzgM6/48bm7TnBq9o8QdoEirBA0gUdHFRg8FzOHs
Zk4NrncEovPaWwSXspFYG+0Tyimp7H1gtEdXlm2mJvyOOoEo3TfCNMRKP0opSUAY
/bkT3hhOOLRmKIR/M/efKOQh7dLJCWgLU0DMgWJRatokCaYOVpdHbSfigYJVx0Ud
gkGOOU5nbg5zp9md0eGOUddPwnzx3wKptyQ2HdiwIB3LSRm30IM2xKS6UlBaVt34
Oml9koxTpWrIu4fkuDEH4BWrRez0aj/IrnaEX8Nqy0+i+9Rsfy8X2/Uz0nn/LyLC
krrvaQ3bNnFq8DVfccUgEl+aBd8KBvP5WE8a1rOOWvWVTVilsCChFpldyoO4vkMQ
G2D/0/ob5RCh9GDdf2dbnWx4udQdsM8G+6VMPUIQaKzLOCc/CiWHuuHy3h5gS8PG
nQ3GIoK7moBwYvijTWsxHcwurgd0wOix+jrnA9NfIpoTFZW/K67R8RKqYK7YNUU1
9d0eynRFcMaZWQ9jQZfe+FpnSiRnWs3uEQ/2LG/otc4MrBLLZ+cLQhiaBuSjiq+D
7+QED3Mli6nmQVFMBrSlracmBgmreqgF1Vj9PilhdMw3Gv1h8D0R3CGFFFkfgKIU
c+kAJSM7ju4nHONxmYKUJTbiM/+czZcjsBxA+c9g7qfuzcZOYBLwVS0r7CGXcEl7
2PTXDKWDQ95ejpgnmTXT7FiArqtGiL3g7ajIqujghK7ZE67LGReyGNW41L7TpL0A
xtxZyY/S6vu9XQY4/1DhL1+NA2m7HWL4dg2b0bKIhE1qKeEKNgsPl3FVBZsTXn+d
B9dhnoh5+Q7aF6X93+1UGp9tdd3d9ZRV8Ok32agMWMU9L9YyGCSB/hYQrSv3nAaz
tg5VWuAuIVHQjLZGYZoRGEJqZl9oWq8qTaLss1h76fxydFHi0VUL6IM9EGRA5Eac
eaJOVJquDQH8mOqLrU/v9ShLV70alQDogUuYpALni+ekPP88DCAKCh0tkiLIJ+05
y9ZcBLXYoxCaf4emD10r19ZGVpFuQd65TLwOBjT6ZVw9htmbOqokBwDSjvrqtQ4E
vb1RrCVH/AP00RXcDGg8UPXTyubGaJ2C6ld654ja+nTp+gwOs38kbVmQGg3Ot/PV
qE1HIuLEmu1+zzVCeUzxcyxNRLlu5NzSZRybveQY0uj+qcF26wFbAHgifW2dMQib
XojDEeNFiI/W40SVLAKNjI4S3y6+QwZUd01BAEZqRjx4H7GsD4MGNjU+aBVGAci6
IBsopKSuEJ/zSkrdn/F5oM1Y4g9jTkGcfgxZMuMTparsLfpYuVz12pQHjmjGF4+M
tD/l7ufhWnV8d8isjTQ4AfKM5CL2IY+zz02jxG7Wwk7Wl65ATbFa8a8CNLniGLAK
p6jD6PGmlXFW4keVMfqb/haOPY+bKZbSoFxHKxGeSDgiTt8CcuarzLCElXwaIWGq
z8qjjAbL3TM1MNmPlchgkWVKvDsLbpRRFC74HiSuA+g/Op5m/8cj5cllxCXSMGWE
7zpQe8w45mrC8Uw3rMeBte0nLWAD/kySf4E2xBjUxn5cyVppqtjh/8MowFzNhSFg
xt61tMSluH45z2WxyTdoq0GlpJEcpxIJ2qdDg084Z0m2JD6PngWYGQ79I0wpLKa7
ax9OZMAew0hH1pntKUtyhvrsZcyu8Lld0SBG/CNkvxr/lMvM9Bf6ettPyOAzqN9T
LoE9NvnqxRF6FNktLS04iVRJpKQgsLuZM3nNrISUU4EVDrmnnph5XGJLmViTMgdJ
toLaJm2GQoHLpISyQ9LplH4PDYq8KFj16DnTHE10/naFDAA64AL0mCflkwaSjry0
iAQVy54jJjzD1+GrHChMaPKQ5DeQQ9H2z0WlVWFxw0XibLVPr/f3gRSswm5jwlLZ
PjVwCaOYtRlfgNY/5OsbuJmTbkmf/R8J+SoKE6O0b+fXOU25JCehDSua6jKFfC6U
JUPL2HdKF71fxO89U2zsiteQXQoWfVpSnR4+oXhlFxd3+z1RMLm609J+DDYuJJWU
nR5UfPVasHRkQ04rdthQoFtn4DuNFwJoYp2Vft/35IEK9ZxITT7N2I2Q8LnoqK0w
5ShZqbx5GTXVIp0kvhGVtFVgSlpZVnZedT4h9rLDfxM7BuVr0ccQ8pzIIZ5yDP4W
COBxzd8mFW6m6dstSeQgCnDeLjYWwr6mjU1bSn/qfWEOH1mtEe0xZn0zqQobqD7t
jT0yERz6C2y55YMQX4w0VRHAALLJcC1LeRfZOui++/XHYlin2CiXw6RbdfAVDLIC
w9UZFilN1bepluipvI81IDcaxUonhKJ/giTKznXaGGBWUZntA9YKqYw8gp1k7F99
CCcJsWCU603CFa3Em7rDwioShde9XpB031757Nha3+PguHy4wIHUqGg9Oc4LPCgr
RaJBY2KKFxkoIibNYtzMV3pVhwn1wMcG1QmeHCOa4w6M4uU/Xbsqe1PY040v46gy
LPjBbKi8LsiDRUpUdbQYB0V0iEFc2++SFty1uNc5NXODglP53gOrpfCeZF7ANm+Q
lxjS4QkR3diJiK25RCrwYHaIaXFwxv+n/idFHWoOpZfRtUD4FUrsrDCBDf4JeqqE
yDjqWsIHRwe/KhkVugjBTxCJUCgXIGLf7CHkm6he83u1tfuQ17f5D/agV56g41XG
LTO9Ya/IxBVk1jXqi0ctAGjN9urGNtIysybPBorOpIKnvf/ORYNaTfyc6ZST4xf+
thruzCNAEaTxyQIuB4lWmp97C/dl09hJGLrV0/U537VhSvfvrTsBuXB9Z2SDxbQ1
d2q6r+JicrkejoPgHMTcSnZjADWoCljIzbK4hUVB0I4w3gPJmq3uOV+tY6W9BYj5
RqlzEoTTGfwfzM8vE+RvaeRc2+hsieWHthyNJQDhqUqWPhFzzYCbRFux59o3yzUY
//CYD/f7r25LR8BXnRZkejH08RmDVVC4pU+GnEfy+n70gnQAKguwdEN5yfICuYSf
6o7n+1z9YCpVO3AHewktLcylM7frFSwTNou1CQftMS031ql+gg6esUWD6+KV/Xld
b8cb6IgeaCQ36b/smAOK5xZtCgvZRvsnhwBlYfVBkDIStsN3+88XHRWphXiXQWA8
XVMiXqdLgdKXWyVCUYTTOwkc6CK6e/k5+qwXB3uc7+RtSsugi73LL41Y8nvPvtOm
fvY90L+K+w/pjWFjcTvQTbjl2zzBAg8lulUzfdCXhxH2kkpnuMkS8fg7L581sxHR
qUlp7tgC3AJhgHWlKCTZ7lznovTkRtGZ8sLbHb9YZTVNuaRTNy0OV+hhZYbe9n73
8vUy+Iv9mgHPQ0RdHQeGvZa72wowWePYbZkBUGHoMSUcQE7oGMyf1g0fDrLVm5hR
SUfPzV3L33cJwsUkx2voJ7ZusyCXDfmo/oMuvTcL9b5tBm77Lh8Ix9p/xJWWBH0b
PHW6Hy3FqRg/FNZmBYc5kAv+bNcQFOfdGPRu6hwWIDO9HBpICEbVWfkuZyjxWIMW
glZnT6b5RBqut5PfhYgQUl7zRTNqdghpDW9FJMQQR/YAj7D2k4ftpoWE7WH9ND1y
zr40Vr7KMpJplCmcqvhb4po8VUZj1W/ZyPXJFccvrJ/BOrn7Ksed+NecANiMpjJx
UACm0aCGhZEMP3WMOym5vEldRc4z54taVYa7fGjHxnmFPMvdh2SWrUkybxXCHRxE
wLQJPcVX1+cc0aRM26OfaGwVeAKlVPaoblDkSOBA1pAst2oN/0UNEJgmXBNBRkJc
OFT/GOjcmZRicfBtl/39AmNj83Ikg0T83F4CiEcHzhjIJiJjhG87A1ljo3v6d3u8
A6y1I8oPUuwFA4YOQtZQP2EOLzq9NnIR8+uAHLfyJ0cUuRKkk8AW/Ds8l4uFkQh7
N+JzseZB89vsRZoshUnQDQBkwU0NZeZoC/MM5uXWqvwa8oQHip8yu3G0UnrPhxWD
cyLH1Itfuxj+xnh+7OabkyWE6dLUtmE+AQt/G6vrATxLOS8fpvtUpiBwWEbn3781
QkEk5t/OnyronNbdTa0Q2vUZErfobAlgOR1A3hvuEGqQqLOCInCeKVNLziI4wAfm
+23Tnvp1XCKhcpt+cHvDqoJZeU2Pz0koG9B+ywTBqQBVJCI+EBaVNkXaibSGmbCw
+iuw9EsFpEfXpehZ56b4KtuubCVf6XvquEq/JCTTZjfI7eXhfKMzSp2gjjXxfrM2
mH0Xc6z2vfw/k4sPpycakZZSwdlhSe7s9QOUmRvdr83y5mcfdSw32LMt1Zju4pot
Lxt/3ONHLteUzz948TgoRM0Ssk07BVNY/ZZ7eQsNANN7l4afRS4WXivQyKpEsqjK
PqoOD1OvQMGvHxsnLDo9M1+fppbG0EivhZAKCLeqbJDwYM9B7mxXVvrmUIdMchRU
nA/ykFMcbR1now+gSHmHNLNc37KudcSe6RlRsRohcS5MX8eL182EalUexdeYkSvP
VWHSnMyIV4hSXZOpIeNHVm9QdPagyb/CBhJt3cZm+pjaprmVGImcbGJ0lwUsJJRx
rErFvAWB8qUbRPc2rgo39pT8eEiTogbrocTHNpQxPzH1KQCEVEmdX+rxSUcbXufj
i/156bgzCQWs3q9LV/yXgQO3mQyhejfr5efq1aDdT9b43EYE2MovUg4m/TpSpJQ5
l4kt7vlavraAaZCbNNdIDt+o+PLGYU8gMTl87pdWb56n8+mdSnZQWmegGX6UrsUt
mdFlDnU+a3NWf7+fe9BwIbxxYNrFqJJWbtu4rlO0HhRd0vJ7wcClBbedDWukPvhg
C61NhnSneU+s7ZWQK0Nzh8ipUcrudKWITyIVWN7IaDcYyzB3Ud43AJ5XL1Ljx491
N0BlTNNycOtY/V+499j6SaQKR958GcRfT/qFk/Kw8sMNE0PMAMlm7RENgEAf+GNA
f3rYyGhsveXKxy1PJTScIRrpRRImeetlRMie2HaIy+X/DYk8tCCIOwg2YsBFDkRp
MgMWgVGklAMwc7BXtmRArb20Os7lYenzAzlEjmv6GC5qp55p69P1lQBIQ46UU/wc
kXEDobWF1ICE8kVfM1idZp4W4iBiZITkSnmVgr9nHFjINTihK86YHQudGFcMXE9A
1X1CEY6vHEhMlA8hw2JvzyspH/21x5W58Lgs3zOzCg01SCe+tPdKENga1Ze4/4XU
9WXPQa5+ttjxh7nAshP8iTPxodSFsl7PjAzo+92hKlLi7+Y/H63nlRDRzXB7Q7K6
B08iVNODwpQtHR94oI2cMDiXfQn+94sMkdpvsVB3mwizvewM1mVV2vaWC0qJxQCM
GbiuDAn86A9NteD7Z9aXLLB4UbklcTopjlJCexvpEXtZuTpQcmNavMuLBNmSH2dM
rnCT6wV0i+x1Xb41zJ4KMy+LcoDcgFP8pWzS/ykfjQ0MPfuiAJpng27W6qeouG6X
yLYNu8/kmAE/YUbrSxLZOShJjHWYLHSvFxS8tMFWofMA+8ndCmmf4n9g3+oxTjN9
SFY1rd6mRMtaSMob8so37BuIeKslyzq3EeJKV51cmOghcV2t7tLplnldyWVGxkyn
/M7VjSg4zkNxOD1/Vns6X6DTfPL1lb5ZQAhQlpSrs0jDa0QGqT6Pn99EC6epGsS9
zEtbeIUDvQydmFyQx9kyjz1vX7YlhfWAJ5yDrK/YE7wg/Xh8z22jSuDC3amH04jx
vpr/si4/EVDUPkN+pDC/DVwogDGV41x0ODdGBM7PZ4OJ4AihANnEmcWsuA+qfxIw
qqKnTUHpgea7+f4b+Rz6EV2KBrgmvUOXrZnpX0AtdYNR3haYz9Y4IfyaoKNkwnKF
aJPbqFVA0Dw+Hvoutathnar7GoA9qE+hECwme53CmPRtQyTH7fxO+PxaXbeEdXSE
Govt7JO/tn6opHNz5dYTowWicrNe4Bp4x8jV4aG+0ivDwZXkuxAUGKKhx36rdS6H
ippGGlBgnyu+WG+V2VYQHhsH/3FIsOmuTcV+mkB/5UwtGvhqtZj2n0vh8rZIeJpq
gFhPG+Ut3AvyPCSZlWIaIbncyeT7JCz6CpuBxiIor/iOTKBuyKX1dl1hiLikdYXZ
wCFqQ1J5X9mIrqw2Hi/iLmruEzqWECSVPaDwLL9mnufP1Wc6C4ibiSSVea1UR3ui
Q4hQmsugH21EIdFrq6pRpa2nl2IIMjQv3l8RoGesw5Oklkac6ybHrE4KoPMzVKGB
+Nq7E9h6/SuOhr9vt9MrOC/PeoopAMG3tcSxUo7oV77OpO9I2ThAwj14PN2KfQSs
f0vEkNOdS6McYdALNoTZNmXWRW8855gqzwezIy4+HfGlwgY8gcLpY5+fB+LNlks0
a9jR6+NMjgoCjoH1u5KUHJyUT2zKUnvLdH1iq99a747R9gRJ7xUeb4TnAKmwV8KJ
UfUBFeocIGjmIm3cAndDz0VhXW97nDku3C0yt4v1Nb3dM2FoFgnwscnHtvh3eeP9
RXm7U9mNT2omNwy4Gd65MUImcxEY7Ybbxl85lhlSQp29fugeORrdJiA3e8/3Aw9d
34pcZuVrkQM4J951CR+D5vJTpQyv0sE+8+rF1Tig6INbI5peaMfT+9gMhEUOBo9K
OEdYzUqXGZ/ejuitTTx03fuVcEvuIKweJaVrxVSZHIoP1UtAnRwpb8oxiIBDg5aL
5AdLL2w5DiXlb6zMP9UZYSDJUVT6UD+I2Nw/f/AJr0u3F6goE89aIcp6gMZg+BPd
GcxUAFDpycQQBSE52EboFyNlZl+Q+TX/63yNqWvsSMBKvnvnWH2ZWBoniexGtwLe
8LxV7A3OpMeaHM5qsNB3b+9mKXmv+bjZHzMUsYSWSfyB6UZoqL9KiqOr5vNAaE2M
TMSx/y9XmmtQhfFnDidzH1RfZqKNsCL2zqC+trA41XhCL3P53bQ4BasqVDhJdLiK
DL4KTr6rqGui+D6E/+JpC3n1Eguqo34CdBTak1kxUXxp1CGZd2jIfzJfRMoT5fZw
PplccyswpDYspkpmdN1t3MHZvAZfYM4cHoTbhdtkCq4Jz5RHjQPmMefdp0x2k7gt
7c0RmnA58R7I2IgmOCo7IjT2es8XcPeeWS7+azkMm6jlOAMPGSZF3yXjx2zTdPvb
yJXdYxmtiFUWN9V+PSK/Zhsk8U/LNZWCmhaR95kb9QtOvpJ/t0opSePVNSN4JtaQ
Ey8gEJdQto/Yw7CJ7LzQYoPb3umDlnT4zQFZ801y6qte5GoyduxagABSGq8QNgIr
d7vLJYNT5ikOWlFs04CaGNKxbvffi+exjE/4p1lvBVFhYP/B99nMGo1RT/lqZ24g
PedAepmgWEyyxImQ+JZ/nKvKMwxZVN4AaoqwNzc61QZ/G+9wJUDQGKu1nA/0jLHk
SCX3D5xo6LJQzgdpJIDZ/E9Kn0Qmq+crG1PGrYZPOqQMuMn1wqTkApDHXLUt5HUO
qq9NZgv2IpV3f0npYj/Y1dSqANKP8s1jpzh21QHbOAmWhPho8st3+adY6ZvGgxGo
7WYGMbqSJmw8HOwgPvZTYo3cc+636YtddQ4alGPMLVyyvPyM9J9/bpOlly400ePX
vXVEcJd5NWlnxbYy2cdtGBpx3u8gW+ATxYGEL7mZu09yPR3Bzn67b2BZbdD3HnfA
zruuPdWFJbMR49KwEXJDj2GHYR+u00RpJ1eAuyBYugPjVO84PZ/fuN9WtSrSUjVr
akVkRKJuLRfrTxYkYyZbTe8xLm466AQgXxxp0OvVFX6ITKunCbXH3tr5rEUNz/Qo
ZK0ecF9DqVBgjE1rFimQvtFHA4SG8w/3jQl63QnKVlTVf8NgNWXWYAxIInv9QfoC
rbJTow1JfwI+FJTigjrPDetzRTNA5tqTBPVeYKtPT2rsUleHKnJSlKIwQSKR2oIN
NIi6BOSjVYJLdStSXjzRCCQESPu2ekV3Z1xv9zeYxbgsIQ9nxYTJz1eyL3DeWRX1
cdu3lJpr/cx5frXHMyTYvecRRjD6MFHBEg+TAMbZX6geV/0KkvuV2ETtfEx25KY3
LLfC3p3HjnJR5ufVDt45t3JuOfJg+IlxI4o8LCgYWTAhKKWA50hlBmmvEOEOS207
NaMetPm1k3BdtEY8lhqiw+7twcsKyvAOt855ZC97fCsNzCGWuVNAv3pTkTlsRsCi
RGQlL0tTnXq6vvSJoX6RN0dq5TyroaZrd1wikPphUSKpLpN65BMWAUQirP9Xdnmr
2u8ubLBPidkajAi72tzB7WK3JbwJM+55/7D/+oFy8WBnkoCiP2/x1NWBCARP7RUy
WqD8Lt6Qda+VCYMWEFdzxJQBZ82YmjpPr3WtUFdIv3AZN7K5cTgu2roPHcTq7DoH
+Yx/+gowzS3npGhvRoz7SP2PK2kEUeT8BhZfcxL8W0CT5lliDapBtFGCwDIO+wHW
Y83USDgR9vKg91GP0UwFv9X4F/llEjIkdzK5V9oEw8TgRioFrPvRMxcYDfe03Boi
sAAiMbzxlBz2X40BobmhpnHcovo0DEG8WCYltJOsO1T3+qKAYrtBxLEVpSie4g6/
njHx6bKNeN1k0SRqWSoLuFY9MsNHGSyT6cD2LhhvfI0Q+eU6BYvfwAm5l2Ihhgv8
ozXLKdfGRkh6BTrlTlC2FBE5uy+wJnj2gQDWDgNC4BcezXYlutjXdMeg9hwt4qTy
y8oBAlsIyAmedmYyI+6M1xa6jzFi0yW7g9i1iFBhF3LxMxB7cPQHWKrSq2G43hSS
PVYeVg1cMrEQ9/ybKJdHIa9sNwX1DIu6G/DXBTGwAl0YaSAmTr/WErOBSg5w4wVj
BvC43sS1x8iPuG6MkWoex6WYG3JNHzK+WpcO3u58AVDMFxEBfJ/EtNj7L/lFt1JA
fVoGxGYLbDKWK0DDsmsGveEhCfDDh9Hd3oKSPVDXJqWO+KimdpXLM8N60tZWjSuD
lS3k4h7plFHY4VrxVgP9Y/hgERtt2DPJDpFsWUBZ3qlPuirECMUwA8i8J3WnStEx
ACP+J+gwQ4oyghefjkRzCP22fSDtrEHkgjCZpO0AWLMPDeP1Wdco4sEvVMfFL5HJ
nlL8eV3MZKxp377O+zMJdXD6LQYJ42wYyA5SjqpyfFqX4v+kvWhf3ZI6Zo280IMa
BKj9FNRrn5BuKqgsVf5jo2xHo7ON3giitmCRS/0G+dG5Yh4/e4lMSy8vqLH0GKpt
O4Pdtc9vYaJrWGLfr2Or/46iureJ3QwbemPm83261b+UFFa4yNyIwSqIvuND8W/5
4PWqFX4F9FocDKEvV17Ml36ukxsRYpeM+a0IXoZLgOz9tit3LQE/lJ4yJ2lLHNln
abNGAKta9q55yHJLMrOcSsGz8+dpmSPPihKL075tAA4lxtqM2XpLDaF+hsY4piTq
bHgKzr+wDmbmB055LmJ2dmSvipxVerXu4NTSZ4AYqjHw9UUWV2U9XFtfwRQMbFzU
u9DW3NfAZbQKvv9xzq0xJlkKxPfq3aNW1PkIgE2V2PCfo5qxhgNPgLfo7pKzkn2e
c6K0s4tSiOuh/Qo4Dvibnw1qh6TmNDvE3Eul9kcH942Rcb7nrfTltWn70igfFK74
hyH3A2Tu45v+/6r5rtT2FdZ0bYqeQwbWs0e0xuOSkNxVY2L5U0lzDtTmeSk0YBq6
K1Z9mDEQUlKeeUlkj4KJGkY5amM7sNPRZYWIlymZnXW/q1nRu9PaYDwPTzQxbK+W
PhgGxANkk8CIpGk3zv0jy5fGj5iF4sIJwMpOPdgtUPGviuEYS2NQ0vyOAV6hhjwu
B6vwjQXUoTKFGKuMw+OQ4TbrDpUUrK3QVse7/qMevYlhOSmwu3b404dnMtmMX7i7
VMqr1//3VTjURpZjqS5LQrl+LmgaujuaE/xAps2AwW0NqH0mg/4vIZcpHifAzOaI
And4b89FU6iYSv/S91T6Y+jZnUDWKpVkA3nAIfDiwjQT27E81hxtn+Pl12gqbA4e
t6qAN/OuWcipPCpTsv/vMXtgubVdixC10+vgewMdnFJNlZ5XjZUyFAELjwXNe5Ar
uf6TJlpVKCNuCBNGKWeJ2LHr0GzIrLwGaIBOI9Ugkiik5UDBhAPIxX4QbwhqGLl2
WsBuQNd2QfhaZZxpUmfDxaD+wqvHwz+UikBiM8xHKP6jvyvGs1xEKH0+lZossTT+
om/nG5MmzPJLMq+U5yjFo7jBTj0kQKerSk/kJD5nn+jmjd34GspbrI32tK1fifYG
UN9h2TohLlwvxEiBmb7GIpSUz4lTtgGhR529hvgvV9rEYuUk655y8u5MbjQs2Jm7
gePF69UcKcDY1cNoyDsc4n39RGHuc/sJAS9rtPRRmPIVgwCpjoyPHyJZpngyvNr+
hvxh2DiH48BczhIbb8PyJglRBW8g+Z0gLiOuJcE/dyyQlW8cM/gyrHnmuBlxOVmE
EerIPKzD30e+Ojk+YFGLziw2VGqvcswDKMAXTSUKw6c979xqlj3ql9apTsYxLCNa
vo1lcGtzZcPCn6DQK/kIimkWUBJDbrHKlfCkqcdQkMuRXid4cMyiXf3MAiIY+T9r
T9LeypbNuqX7EA0DmC19yTdNStyj13ow2mro27NI9we3Ol5HSWhs/L4mkaqkHKIE
YL5TBY6WkdEnqaMNXhcb8U14OH0pDBFJEK1FcKVZ5yd3VezWfKeS3Qsv/h/LeuW1
/GUY7JT1u4jQe8WqRbIyd/K4pIZ4OKAx+cziMNEnK8nBoCc5FlaY/nkYNqwsCcD2
agT8krqs0AUjJ4/1XVdxrBxKBlzIMUJ/asE7b6/t/kB87RDutuJrREEaPKmbjCJJ
FTo/5FTLiFN56EdqNsc9z5D439cYKVUeMUXmEFmQ0ONUOwGBTc9GSlnz/VPLvwy7
2cfiztojMvOsMUysm5TMtMMci+8LJQGENy0aAzuFGc0CdRILA3oIsT6vPG7NEFYV
CjEgvr2a9onwG0r+Mbtk2sX89s5I/LuKrE3EWfvVzE9EVSkaBnyWPJm9UF/iJTrl
o1wHCup41Ok1bNNPrQjAXjHwykkLGPlHlJAgHFhXpQr2xtMs3apJDVEK6Gr2D+Pg
WkaN/l9E5E4x4518eHCxSyZiK7cLajw8P608EUxBawsrMoJ1nIPT4Wa46JSGcrno
/EGIOCJ2G3TsuTadenhytVI/21MwrQJFFc1OmWhwHQJCrspeUvJRXM9V1nIaCJPo
/97LufLLGolxNOSE8mh380BPh2CQgClZnITaXA/mQrLOrDX2/4k9/zTHmPz6B7GQ
PobioQSccL7vO1tv4DDk3VP5qLnGA/EVzA4Lzs2IFJ1Bvs9q/t9XHHVd9IQRuU97
90eg+7LPSOOMLSVjPQPO/2vfaNDcG7qzpux8toVSM9u6kcQyQjsE1grnbdf9VGMk
rz6Z1F3ncTv8rQeeNwp6WbNN69TwtrP4H4qUZ9NofRVkczfxxvYyBuyXaK0wXUh5
wtBpolVgmvp7U4hr/unPtyEUW6T9LKWWXusF1OvY4W49sgPiPvxaUhDtpk4P6ilS
YBP9UpqxpVZRxP5ne7MaXHWQwSDIQefm1hrTZhvh3KQ5lPznNp2/CgkL5Ta35Ds+
Wy8Amc+HRH0VHYu821JmdvmndEQ2tjxSdlJzBQ3Yw4zFx/4KhazJIKeTmHXj32qt
WigcQ9LhX7WlLYg5qxg4cKbJ5pUBeCMosLNDCsKc+FiRE0U6tEkd6fwcZMWbzPSu
BokQWF/YI+Rm9KQvVNj4bk1YyeNezn9nBCd/Ixs3zCI9/Pj7S0YDJudVqaPZ+fzw
neyOJlktkjN8ITETO3jc+SaFocT5Mg9gcqqC5kKUjBrpp9N8Pp1/uWaSBiqIslE4
9JtWm8ua8qWmyLshwB9a2uUcgekBCTeAHhQj5XcJSKPXKdEZ3zxq2i+VcrH3zFbI
K5Xv374GXL7tLL9GZqJD9RCWf7UOuDIqiPplEZpph4rJX7aGxHyFgJIgqyX8WGez
HErKSxTSzqgDlv9FKvRCjwr8abn7jMSi0Tzhr1T+wZvcwnttWBOaSZDMV1KcLCb3
PpJNH/nmffB23js5Yk2HRIIdzSR0YfVYJ2NYTtdSYt3Q6eanH7X5HRJgcuCDnMf6
9xQi8OzEirj9klPmXFCt0/FBqLOu0XtNHB5mkg1SYQt/tzJJORnKLGLWsghqoPnS
3YBFnJJcVcm48qORV+Aax1VcE9Yn90T1f0UW4eZvZffgwlsZWnuti6rf24fTv+ag
cdNfCfyW0HdLVdKeRE1bvSd18OfJ43KtSfSxzvka00TCAFxTd9bBwSuHPfW287AQ
ck0Vta1lA5kwEplOI4gCA3N5gOH9eV3e4Bg+nGtleNRg/hEkJRzhI/2b0uTcQnXx
W7/bdFKb9K1YfNTvB9y3aOzSnmoFXzOdXQLucLnvygp35o1A/aFHmG9YgywxtKIj
4i/2oObwIt6xHvnVLddseGQuwwEaiNwFNXwt5Bi+nqrALDuSloHimcSNgKK6cTbH
FnFAraXc4xamRQAdFDL/Xk78VUOS9d0wFdInn0mfHH0Xxg8ZMEeJZVZ8rb0d4+9F
L4Eax2Fevt73tZooVMfv9pyXA6CiY1FWTET00331aJtYSiInyZqt3JkQhHAYML6+
UEoJh6eAkr76AQ4EX6N/3ycO4u8wfaHEMkfWbf80S3jg6zwGq7cjguHsUgBQ6Dm7
fj8wAX8GvjaGwC76DNRRJ3qibWq0AUMMppsmDTmqYOeSmPSjY2ZlPEZBYoLvMCR1
RlPAyg33SfMbNxzhj2jQWeBpcdzV1svIavNKo/p3PSmAMTWlWSxGUVxNLGpbGEqv
kPD1uQ61ryge05sGVrnZrhUpfDZd9b0XUWJWOsfCgU6Z+6Ugb7tmxU0ZhbIUTI4x
90ysLl4DRwuh6hqLTUkt5Hped6xgL8Cof3YdXUENkrv4Q+0Q82Vroge/AxpyFWdc
nF1+RgOEntO/hOajDLKnukVCq07IfY0/CkxHGi9huJ+7dXJSknPCgVENl4G6Mb7T
nlHGrePUCcimyvm0ufzfT0wnKwjpENAD/dcYfqktxsJqriON1jSSWU4ldJ3hgR2g
DflLIUA4qlyroPXZ/CSC5pbgU3ztblIM5q2G8nSatHSAb3zyOy6V65e9FjIlYrqD
MgPiTZ7B7GsvUCT6ny+ftL9+KQIHo7e4hhTzJr89pRo6/37WlnYpS3j3MVjXQZkv
4aZyL+DeOHHirytarlVeeU32zGm2ppVk88YCNSu/3gI6KJ5e3mF7LPWHLoh2/u10
FdOYUSLWNTKhSVNxcP89KadC3jsBzukfMD3h3DodQY63c1l4kZ6mjVSzCBtGkGjv
AYwUOIfLWn1sRQ6sdk3ohh5br/JRYrCLbyRM4egIjQTwxTKTIGLqljc21it/OQ+6
G+W57BZfSYDo3aDuargaOLEwXJXdyJr1bEFmoq2RUCQSGV8iWWv380yMHQxTsBuq
xHXHBLiq9EgLAqRQz/Ea0FUwMOUyXcwnl02agDK8fLOP9wXX/kQWQPFBofEEu+bd
7O9nZ7yeyhpWzzFmjoVywcOtf5MbwWp5cvvXNU0M+Q9RMSkSitI0fXwd0s1MSxXl
DnfDQZgfzC6is5Al2BAJnXpF+H4kmijIzVKAJysHc1u4pgVBxTQvkjT5qTuJCtWP
Sst9Rypj/nF1P1JZJ+kZvqQdjlTZRnEMejK5H1jurrpIvDHecljBOBQ9VVp4fwon
oHJXnZWLb7cDoKurp6ObHvvMaYEkpuFypYq8ZfBnNC9kWTmRfjlNM1HtSfM/wC92
tTLX9VIvPTE3FprB07YQFeBu59rdUbDOu5wBAwg2C5hC10Wr3TZWZxBm1bpEisGp
cGf4JCGG28uzrKvkXBagjQgq7m7ZzpEWehmVYSGOJgmyB2xsw8AO+CxFNO0/JFKV
wlQMju3M1yWhibrypLcidnVCLjpm/QY8wbmN26THbeaYwFW0irJEOZ6h0C90tcim
obOV3+MpM6WnJ3eXHj/UCIlcLQBYIIz4fJpzjDokVTDglvCaqCH+PGqfGHjk96dr
KO9XSyyjaFM03prVU1bvb47GE6hVWSa+9adzuet6P0LKT4qvTtz6SoizjxsPTyMf
Ye1oMgliy3S4nwDG+C25DvLerkefV1WoZrm961sFSSBepwwG6OhI9QqOzgQPoGbR
pXGNLpZO9P35GzsDXsWoSBesT02aNRhFYQRfvYWNAOkpBhltwR0Cq0v0H21rVw2M
XRXOpXTMTLLQ++GlioWoPy9dRDkKww5HaVFOuq+uBQ7VXGjwDDH/sAG/vlGW1Rz/
KMgnhyVfQgoWXQDyGIhxtGOlDkbk00o3PImaQpFcgHoeT60Zy1SFPSkxaiAC3bnE
T8aj20e6dveIUySB+RVxogBrUX42IT1tUgb+3DJe8V15VHlfm01IAIZN7sZ55OYK
hM++9ze3BhAGIWAMzfP1RdSrFRZRNZpX9tWPydaS3+6WwjlaxLd91aea0FCw13tG
SkrOJa8pazgMvmN1rdR+DjzXJGFp4L5AwFcrGHehcOSEmV5LC9yUagUy7AsOFxd+
jriVysFeFqXr3dl87L58jwEWkH2MAH4Q85OrbFEKN1u29sWDwQH7e0pAXrJxW5OF
Pukr/Z6ubJwEGEMdh+vmQtaybSL9i1/ABvgpkwEFHXpjK/bZU/+cIn92/s7040Yi
tA4sV6kD6piZ/cbKvRG35ol+tXEkLC1KQJuoLPH5kKzhoi9qODr8GEVW0iwBIFGx
e2Mr0z3AsOw0dG1SzqqwkUpb2Bw6kbxm6Sbt4yCSXSO9duULddx6QorzUJtrleH5
yl1nA4tZ/GpNKEmRjFUCLaGz6mEUp3iwTVeSlaNeK93A5XfPfwOjOkaw9CQCaPeV
ymieiCSr+WtOHn/ny4BplS24n9Xb37Vfy+pQEMnPmJ9T3azzz80rTK7Bk9g4Pwui
LqUD+25zSFCZqhfr5yEOdKEmkN8KLFRbLMpmaGaG7ZmNp0r/9ED/yG5+2syR5UEu
vY0WwvV9JlWlDP9XwC7UUXm69H4603DYC/y7g+bRfYV/cBcgxaWz8zPpCDW6MW0O
Ekbstc0cxm5wh/0YZGJ95qxco6UHy9mYLRxqyubit21U++gysYNjVVi5WMTemcSP
NqhSIbSYjxqkhvk0WgRkSH78nIZiiQyA1paVgISvOuV+6/AjynGB7oXRL8XQmOE3
vBZH2IySkuehdcxL6aqOZW/aj6TKQJC6KLEygY0YIN0ItqTRYld6l00sUS/QYiAk
Gz9Kwu19a+PJEOIEHsfwDN8etH9cXkSXwtVxP23vhs70BrREXmzixPmagwZIxRXf
3ohwURCeQOTYAxNMhz02qcRFBTuejThaWLfxBIbzCTw0hFllFQolPRKs1ImoL8lR
GE+owO3SWX9hHpK+x7PikYR2t7YczMM3YxgVmiQYWbibiQfuSI0coyvh3uH8p4Ww
1nNXN1ikdxTsDJg4wq24NSfSqF8kzetR2nvPfY5yLs7pr6K16YorTc/rgX+0dWt3
pOHoU3NEMArUmDB3gTfocp9N5A3bIxm76RvS9QJVP6wZPY4DmIAsqQ2NWY0O4OJT
s5D+H80OwddZ4A5nTUaWybNUP95lkuXhtq27bzJssvyaHENLFaBTaWtor9LGw1WC
s35127kMr0ECvfadvYCwNrKb91zrX9APlyEc7TboLZodqTFSL0OF5yAlADic438I
Go0U62vPyYk2Xv8CshJZ7ZY+CQgiE1EmdfNkGb1fV51fNq/mW5xrTkTv1QjK7mML
G4qODzgKYhZWbNrDrpTT3caMQzyl3+4mZxXDVFTj00CXDI5dLZGffMJ8lzKnCQSU
cfmNSNZqFzO3ikX12JjZLXHPMDecPcRA9faPy4mhQN0DywOMingEVGczeFxh9C/9
q3H/ufDhoWxtPUY6WoFrzT/dau0JmhhRFyUE3IYRob3jKOT3h3+VdV1WSziD26+8
kn5qoy/tBjFbfySiUiszBEWnBGUy3Zz3iOantuxIxVQ3Z5E+watNHEpLjwUtXlJo
qpI1XulMwAhiCVMVDUkTGOJ9FYq2muxZPhrTmK2hv44bSjW4R3KtHRI12FOdTPec
ba/5Pdh6UkNPT9xE2CZhNBVwl4UQ/3ZCVaQRRdiS6GTxjC8+YNmKCRkj3HVu1jaX
v3hmH4GjqIMTxXicCx93j+vN/2ksPJIgKQHFmMjedoF51yP/PuEsxzSWI/e93Zal
P0Dy6wHf81oqt6K9qOK2D87PQJaw/Y7BtwvO59xHLX4cGWlcZX1lLAsiZ9Bg6ZAZ
iQKjJQYQ7jwqEp3Uecl/6JMeDlZEl+5WSZLqWZjmjH/GdDrH9dKIOE7hGTEevn8v
igl0TYMWDDh+GfE8R47h5nrryl/0W5kVscQwb8oU4Cp55gi0IqloR5L+aDRSXZAA
1zycd2Xme5qyGAnoFGR9sTGPEZh7gUphTd7kpvgstIMZo0C4+HHkn1CyiB+63A52
rqU1itwp+7kju35aFNavWYV4Y8DPwFJg31+L0Hd6kTkWUQsOhwBJeBgmOPs2j8PX
oVRZ74rzJUIqQG0i4QFAsjNO9pU9nLIRMnuNBTAQJA97PZ5z56R88QPVyM0ghVq1
5kOU8XDDZPuvAg1TknYNlCJ1SlRurLqJbhiiClZkCQjtAeQC1qJxti0I6ncvjXed
4NSrsyrt7Va5VbR3B0VYJTshOgNrkgXXxAJBee5t6w02qdKhg565lYcoqH/uEoCp
0btyGPXcjyrXkDWiz2QW06UwGkjyMOutBsQKEkyMtYeO++vbLl4RLe6Sj0M/b8pg
DF6wJm3cD8qRmxwl48pTRIxQVmea146ed4FPFSkMw+9wDFQbftdILTu48sKBmMV4
5+AvGBRczbCiCtt51Zd7wTLZttt7r0X41sBv6Nbdhx+QStrZoZ39FZufVn8xFSTY
JVBSIhDh840lSlo9jwnZND/dy6MvRSRTNVs//iM3KaipAvj4fBS3JKeqKdFNf65j
/4G1hIgQBtHphLFGxSJSNbmLGQMNhKrTsXI9AP+InMC989WX+CHbDJfmGIhA1R+3
jqgd+L2tiZNgh7lZSrRyOGYXXoyLrEkbIaW8yY81qCTpUl1G2MGSWW+ysAJmBMoE
ijeexl7N301rwbDwF/xtpNiJ4Ih8iBvu+QRvH+7nlFw7QoY9Rplr1JKEb/DQJ0mh
ozZP5BlW1l38sR/a/CyM4T/r2lMS2J9qjwydOxeMCSv1xHCPm9VxipBiLCPcVkGp
KZMrS4cOO+D4uebGv+eJTcLJxsGuOwNBIBEFRviFOId2a/MeULOyyM7Ai9Dm4jbI
RB5FOOuP37LrBE8mzz1TUEdtj+KvEJ0jA1uxMLuTwDNvqgow5bdxrMZQTwCe1QBw
1SOY0gjlUS53Z/ZYhY4qw6SvFk6kb9g0DlVpbA8/ghC7Vfwj75M0CQ9iJ8CVc1b5
SjqEHkpPzfGeo9BXR5Lt/ieuexkaADvkLbIiQHCJJiBaRd1D2Boydx7JzxdK8KLM
9gsbE922gW9EGIv82Z6mhsoU+DL3Ssgn5iWeDqStSy4w1H9a5uH4ZLKnzrj6h91m
KDW+rftFD36U3elAnDTb5uQtZi71y+rjzuay3tWCxUGaUPqd9dBaD+sIFAJfts6F
ideQyxTq8FeAvo5zapHPVBVfR5M1eCVhKjWLYA68+4JqF9hVTx0gUxgewxXa4SKh
zOYuKuhZCYG6kqHHLhuk2JAJWDJiGDRLJabzctoJwUmbX95l0yGTmoRlImO9pBCH
lw8b/9t9B0waByGAC+M5dMPaNl673OyDDtEC4Qqr+K8MwD8pK9yMR9wh2ltINmMO
V8yNrH4L7PH7J6IDjR8CQV+MWVTyZy6QEu8Tvgw5Ql2I761E7WtuQpSVrPHV9c69
O8dDkHA5yEc6M62LdvoHp7IBGEHV7EMucjBRXQtGop+41b9Y2XofZMzs+V85YcFS
gPdu7nQ/LjZ12pPE7/wDYmOQl/az6l6VJ10ndTF/KNif8VI2XI5j/Zi0FG2uxtxV
hyASvjdHKOJzREPWtEPAmfC3bbxRf7GmWGDZnoUHIPSrbUJyiiwNDCvHR0LtJ4Zq
b8WWBOGhGnVwswSADGQJZq5i9y9TmyuTI4CZFx9CmC5B+z4m1XyEeZwS9GerckQY
w4f4KBghp3a2q0xKiHaFvofGYV6EKPf+F9TCTWYW92QVcgSYaEYklbHqvSRj8/JI
DeEbxnQXhWVnFs+ZnY/b/aa6WekxZpf7crQYVGewTN+8QMarFZ2PQPSaoQEBNfYH
UbUTwABQEDYcWlPH5rxxao7rymNAGgfv8MkYsBrUQUaflKJk447xX6Gsy9ngQ/+l
gh3ZCjH2O9H/LGW3u1+tHmPo8Ei8lKtheDLjbQk2MAeeyo74rDZHPC7ZRdc3PLdE
VpmWXAefSY6wYL5QHvBc885iV1rrfblQGNkA5FGBTmUg4ywpDbWYmhYUDbQgkZ3A
gtfurCYbkZqPgsZn3thkAacS6zaUd8Nbah2dvGjWMWY1297jOFHnTnilCdTcJUN5
xiyOStppihk9OX5aRcAEgDS4GUdOx/TpAU4Jrd/Cs36QZ/AKZXEYUX6JTOMocR/X
smnLrm3fL+Jy2TLNrkPA7ypu0i5QzxkL9eauY2018j5xD6x5nDtW5P5JM9joVwAq
8RilNjwDx8chyAVbbN3N4uxYgBZc053aRibAfk9q4yuJtS/OgIsmFSYlY/Xp+N0H
36x+t6w3DTeNjVGrEvZyuIfu/zRZBcFxv/owsrpaXC4TIhOeHyT/GH2Iy/76gOrH
a74dbInE24c39bwfsVrCHhK18jNmZ78NbTu6L1cuYbGLFSQrC3vYMBPtCXARkD6V
NBajxiZLBdIbQgweErQ4hnCIxreu6OJR7YiWK/uJgsrHG1w0omldJT9PLSFnc995
kpvb3amdpS2kpqCscPlC7s6fgUxjJWKxsV3KTmlNUF80/otflmPnZE7DWslava4n
iL7OUHVcKJ0H1fmJ4SJnqYEahcTSISdWiSh4y5prz7ZbDst2gYWB+7TNnFX3buDR
Zn12bnZurGuuHxiMzduGDNy+cRd5GFJdI6qjkaUXZdakodxHKiQ7ywV65dAdapK1
siHvac5peyGvfqgsBln9SpcEBlGJ00Z0tFyktYEInK7PjL13hGAfakUaqUtLUuLo
GFDDte6Z3YkzP28rp7kS6U/IZBsuX43zoJyIB36CsTv4E5Ns4zo7K9nRQRTsrNvI
6rkRyNWgnseg0q0iFEYDoBBt0aMGzDlY/cCSkRPQlH0Log0LrUspxRBDWreM2lvy
Mb+xLDVIZPm0QkYPdkfErNjDa1PE7EPR1VrMuUtI1gqeYOisuAF7uiXD3ibn1RQB
3HymC7lGkx7e0uHTgUlqSkIh+QE65stAjHyc+7e1jBQEBQVzzgeDT2L9ml03PO3e
0+5sz80NBEg4zOk0t+YQyNrNN4cEf73MzkxjPjp07vNMBPW655qVgatKGZ86VY9+
AnQpOre/YtNh6klbGx7t/cyNXGGXo4URHend4tBMY2GuXvtyPBLEYDs+PbmnIRJ3
yvAlajZ7dKC69spx05ht+MiFwSiEEaUer+QnTeVW+2FiFjiEsuSKnVBeO6vph2Fo
01XQxTu3s4cKpwUH2lSt7HIzlfVCJZQLy61YpXVvFxpQwM9ZpWLFj5omkMnYA2KA
k7+oHdh16P13UqD4t2qasdDwxhriXcWsEAGxGCmKvVtaTlUJh8gyV9DJSfrFthKL
PGWBboAui5nPQiGRl4lLZjgWhGXQ50d/xP37Jcc9fl5JLXdgMoQ8dfcGqoBZcdaa
vswPHNFJjVfe+GfjH/uz2ubuUtjRNAIEt5iYYfHUdvB2ynQKT91vB88tF1M0t1Iy
OnYelJkaevTTip9sEaAoH/mSbR1yqTGNOiePxizkB78zTDK7mL6TiFIl6g/kcm+3
cBR7wjAph4f9BTL/AAzzeU4Ww81TmTmFEIwf8jRgrn2Q03FfWvmZVT9dQyD1KWhM
TFz9LuGJRZWZ+HiJFwLn4YoxPTXv3sm4DvY+BQy/dV3d0uDJkGQdxwWLe88zWuGs
eWoQ4yQJoZgbINhga/BQKYsUZKaDgJT/hmPmmCxFMh0ug3D7VrPuJydyqrYxx7Tu
6o+Nv3TXxqanXl0mpp/py59Kk4TaQ2lG6ru57yM3IDdrG9dTJaYeQISTaIfwHKuI
OsVPsFD6PB8Z1EKIOyGyLwUX+ty2Zy53gJkSWy/wG7u4QsdR3WHqlz+3B40fXr+z
053l0RLgQlbhlw3TkzSqpo9Fh84E81MDSOPhx7AWLqSgnfCcmVeeooo7Lm1QaXgb
UTz98Wi5byRS+RryjvWh+6/VezXyJg+TatsLdoRg2y+Yxof2+dWMyFVXWLVO8n0A
Mo+98KbMdDQky5vZYROAwpIPxywkucr1F8FqLr6kcS4Wa4yuzaSB9O3z2RIgogar
b6mvdkEQUZIvfsTUsuOuNiLRGO+IhkAIH2Pe9zfNWH3YIdVscStJk6VqzKlxznuV
KVp2rAbuZpVmyDxI0Al8AqnX/qUfJtDNUlaugFvS73/kuGY42gxXQh9aFy79l6uZ
6sW4Sya+xwia+29OIOoh1rgqCRd79iNb80dLbTzHGdor3ofVbKWXk0tfkTjyswVN
SsniAcSpRBsWYKFQk2IGNIR8qHSibm3I0Bt5mjhoYG+z4t0bScLE46iqtd0Ig8AZ
GjjWSmO+Ai1//p3APzz7D8qxziimrXBa6KJMYkUGrq0eNMuWrDPIegYnbexzYslL
xKu3xu/hUBsPtLgPzuJtBLGN7iktQGaUgP18fx4lUggZ6OWpjgj7C/kagibUAZQm
qMTZth2r5inNKSOnqoYL8Yiy0h4DZsKzy4e0lTL1vsY5JAXIFlrhdpqicCKGFit2
iQO9pWrWET7CWSdgMtJvoguI8dYibH0A/ZQtSU4Ki+X49kqSj/2RDPvZLFIItAkc
8gQO+lpVrXxDPD1amcSkTVx7QaW72QsWzyrrvdrlDB6+8FFCGhcKC+ELdGIPTJW+
zhS9JtibQ3wnAoYxrWx4PmbQzFFwW2NiZzVZdR+epjxb5q8pKQG7/GovZo4Z9oxD
8g0yRQOcTCI6aU3VyVrmqYrrUIMuyOgLdTQKq73xTMc1GbDey2fFxkpwjVBBJ2O5
jnMGXOO3hRlUt3a+gvAV6rlRdnRitx/w5XVSjIwNUCFewTeyxxnvyJThENEH1DOy
Aw6t2OvK3kBXEoekazygVwGlV5bbaL+vWI5DD3h6OqJbWmLPDERBebmO9+dF7lzd
1bSVp5Z3Tywe6pJ5eKJ7ztw74JbjZqo5gRTCm8jh3b9rneZnsFN2FvkyBIGHQYYA
WcmqKh2puMaqo4vdiWn48idxMUX4r+/jo0evddJkG1SxMUikm13CIl7aQyIJjbd7
dRb/gECjY5+/4I8rT/5syqx/wOqdgtz9xiDx+dWgkV7Hd9KGkyMaurSDPmNyaz42
/NE7TGpN4htLVrzMZEpguG0f2OaFnwMw2PKTanIT2rMu8tk5HhcH3vI3xrg7DUOo
/MnH7PXK8ILCAm4V+yKvcolp0KqLwNnIH76wmF3lfQJC2kORDO9+pXAo8ZIhhkWB
LZ6mCuFREEbWx996vmNEg5pMgLJlzhxbva+pOGBWXTvHIte4Ch1uxDiEHk1bhxhh
DZky+PBgEOeXxvA2QhlUs8GtgHG0h05cZGnH+nQYkYprQjUjijQ632QvHpl/Udyp
GSHQoWxeZDqN39AfKjx8ELr4+l5xGTL/nsQmUc05CyiUPoxGZJOGaubKf+NL5bF0
9br+KxUCuwh4wxC1k5lD+wizpQ27Jk42jgtcuo+3J9B15rDMVvxTbfghXKZL4Ws0
0gkezrNfB+y7wl5isYu5lQmobwRe59RbxJDg/+LtBfNMMrRrFtJnfejJ6W3T+gxT
lC1xtAhjMwbD59p+tCSH2eDYLkZufZi8Dfr+14ZkTkw71tz15zJ4UtJI6qr1mi94
HGpPnPROdqZlhiD5XiI3UeJUW3ZhpAxxn01EQ/SGQD79zUIgsHzJ7NpWNHfvvUs0
XvblahyQw4xmbBKiRpcOPPIRHKWkhOZCS9Ee1D4J8W9+XfNJWfrHKUV5trkEYOVr
r+aVwWiUs2Zc9sUhhD/FiQZVS+0XtPxu7Etv7tnAZf0Pp4wtbcHy/F57W1H7a81y
g5RbxCWTwBSkC0SkPcustMkiTwZBBuph7rpS/oc7PLPJACf42mvVDUVG9OO+2o/x
l//HkUwXy/PiA7NRXJGQ3m4FYLRX192gTPba8otQrRR3TmV1zKDufOwLiyP+D/qt
VTwzUupvZObHpzQePqFaIlhI/6qnWB9a+DOIur52PhiHr/E1xsQfZlfZA9YYTR6q
XU0xkJl4Nn74/VOb+3nOQQ1aaVZbECAKvp3mw9nin66/cUC7w8dW2Ha9JpTIdT68
PodVMsbW/zT+9yd5/VH2aQgDxPtDI/C/bz/bILO/dVG6anNnkBB5nfsBYztTLvYG
UgjZsqnOLGuGERgoUTILodKhdUXzRBxKK5WheZUelbbTptHUk9bL3UheOb3QvOiy
i3u0eqBsjJXoE5w53+poj2zmknMQO2mvK9wojOGgFo+cqqTzYcASeZ87Z8PHzgpE
vhp0chw9pba8oIImbJGQvNtnmL1j60J7ntLHKwxGTSpwCkUd4hkaX8yH4wNAcc+M
JUSVx2xQbq5gamPe2Jlfy54vWgXjN4xB1UUFwsBXto42/tdrMfewvheB/Rgb6O03
i25CFlwzlSm82E2eyn1j8C9jGpvDTQgCJBtVKQS4b9EAMaja8+JX8GJ8VO6u3uvX
M39MfDqBVJuqXoZajBnD5sP7jNM0qab2568vavM+/sIs5CwV/M5A6yO6pHbMjJZx
iaHlYgM6AQDr2H3ppJiDEyqY1LoyFcOGgB1KYkG+x65jrol6uRrDoFCKncjnti2H
Q89s2jvpZWU7GVtYiYRC1Vf8GWtNubYUg6SzrM109U+AwBGkV622hQmqNn5/6YIp
qmVOQmVvkZ2DaquQau3JolpqV83tm2PksYrtEp7SR6OAr8qgegYKfKpNvWZGRsm0
eIcjcSaRrOoFMKCVa8PeJw==
`protect END_PROTECTED
