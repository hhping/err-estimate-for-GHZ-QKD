`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZwPWDcRmhvldfYxlPbqbmL4OKxGMxbRNnR7kfWASJSx3sTCsPc6YFJbnqO9VBRhG
uFM4mClxUoOoZFxzKw0BCpep+VWpUIeyMK6AkKvMzvpEEPeH2atrz79a+FIgiP4f
9yaNrr0E03zcxdbVLhKSNxPEWT/kqhipYfGBtmr+spovjBG+CFHBcYm0AfKrx6Tl
qqvMufkjKGYIxElyoFCAAB/H+l8G6+TKJvpreXqB+CLzt44a/Eng6PpJ20T3pttq
n66IbVK1bN+e09rlhf4GoUp8j+nfoGR+rkNTv4ipwRV6itOG3uPC9VZ2YRYRnLsW
TgArgyqnRuKkJ5agsN++n5apU0HkwG8+FxixXAon4SAbhfEuF+XLsPtEd7kcowNy
WAik76yg0U71lLJj4gDudTtf7Cdpq2jCkv85GglVYlA77kGUMluWp0Qx7FlL8weY
x6npVqOYy4/VzJL1lNqfOjR4NOkB163+ab5TmsCYfCwdxf128C9wXxaeYNuFG+ef
gefTU7b6fA4Sp1k2anfoU6t806oOi9udVBSApesdBSScyiCwKrA6JUBYOu6TDETM
ty2QWqB1sqfTCS3GLhkj9l6daCy/2tusR2bWlRA/QnYHgz+2QhJVYQf5PHDQ3BYm
rC5wPPahel96+0v0plH5lX5xkjEDKRvwemG0PJjyIAvIH4fNOMjf9j7CqqMR4FNa
FRzew37XGyJ9URUh4R3V15gRmda9yK0UBPZNwH/e/bNT37WN8YPmP7dnoQgNBnXZ
93dKdEpBi3WI3DyyN+50pPDwdeL3C5jOa2qPjRuLXNHrl7PILVH6EZbWD/mo8nt9
Ik2bdd+bnPti4pxC3D9U7p8gq/Unn9wDkb/nD87wEjgWi9vqKrpN9+udSAvgwW7W
+MTzF4Vcpn8a2akV2FnUkn3OW50zujHbKUMCV/aX4oWbUN2QacBErz2sF++tTiB3
07FQHJpTKq5iM7uOgWJy3AbApvibO96AiXY+YAvopf2uVToa0GeQTO5BevnkfSzA
`protect END_PROTECTED
