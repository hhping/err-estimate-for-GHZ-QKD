`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gXkJcFcdHOFJiPj9NsPY0/H6p3fNr7Mkd6OUarAHI841xViQ3jkW9cj1DKzdg3w
awnPZ0VEs5v77Ud3r2L/fxJ34nwCQ2KhEg7FK/BsAK+N7ZECFK9Z8PsR3VsQsqH5
fpItWUlaivPjLvIEl3O3E6j/aZOQMew3bllAHaWnxxXRQOQFz/6lY9TLkEvuB7Em
jpfIYFCAZFBMSgg3PX3DSd4ZXyOX2HF3OzO3jeaz3uz1go7pT3Wq1jBuGeXTiCtt
VnwR18jvAFgM94HZvrdu65nXAzhzkeNvdh4BndAtHmfvpMfIXl/+s1SYzZQpDPSE
uOWeg72TZqTPu8QMn9y5jNgyv+TDkxXeXN0pSS0qM0p5Lvf+0AvU30zFzDtIoJ/+
ycXp3YemNJuHg3hFB6Sv4uaG05bXlCz24Dwzje/0108jMldVsf1474CK5UqIKTT9
ar9h1udC2ywNVsd0D7q4mNYKk7Kiu827Ao0c+2gIB3mER8tgaNFJ6vf0CnGKBPe3
490hHDuEGdqOgEx7jBX8vLujWgwuFNrn9d4uIztry1Q=
`protect END_PROTECTED
