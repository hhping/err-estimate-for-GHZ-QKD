`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7rxqJQuZTfXF0frN1QaRjBcv2EkeWF2E+AFG3OaizM/5CIDTcCoNOkpzpc9vFape
3+C3qjzLGAbyfbTa+6U/gVwdoS1y/+lDEQqLi4gtnTV8Yn4JYBTkq1JpFIbOeVv6
vAyjfUsIFprsjjMyLTaL+rDDtivA71NsNYyDZX03yatCPe7n5UCYQl8iXIlM7V5o
fcCbvOMvBibiPtaBAbg0utlvJ3Z5K3lLreVLn+H5siz0db1wxy2qT4yzRMnEVvNS
MIFQFu1PF6Xq7gtqCAFXtbtAkX0YmWNYMW/eL4CKjowMVnuPJj9Vu31Vkv4eH1Bu
u+SiXLj+1rLiDsOEQg+gg3WmV7Qd9IXhXVGmMjxckD4Zmlk7LPVWHgqVoTBcPa4Y
ejNVhKL5PAbnTUWbOPioGFsW/6GHcdu+VYoqj9iBPIUyMQMzWZLQKvZLbVClDZju
iHutC5v0jx+AOET2OIekJO5FrbjgocVIbnW18o1zDGQTO3RUUALasQBAATsygvJF
oBpKY35sR/tV+ALipn6/Q6YLaRp9RT1eiaPvagbjfbbRtV+WJS3/1HlDXwNI0aO9
yEdJXm84h/5CoVgezmp7QLSvc6RKEKS9PBTAO9qznnJYyoXTXA/4zZTfICULz4ML
xNSiCFLP+iEp3G3MhNUi4jLcmsPfAuCRRuU33TozgBbkOlzWp0wiNthbFiJGcG8G
1EoP47n05EQUE29t5a/tdYNBnQM83dkKDlbaHDbwd8UNAuZTGB8mUyNOk+e7g2JX
kNeKDrCkQ78T1AN8Nqh89KxQP21DKxwNaXdyT921mYkbBY/sZy/e7w45Q5pC1P0n
8QJ6ytE6lonvkT96HN2U/QvuNAu2HiIIt10p+LiQppOlEMOQ9I+msYl4fsMcdIPl
rMaCEqxKMIF7JLHe4vQj5QlrALmAFXKiPqahtG5YXktaJc2OEj4O6WGUniRTDto1
x3Fe45F2uYaQFqwHrFcTk7n8DZvMcVo/0o+UJj84Pw8PYERXCi0XSB9T54MC8tDs
iUKKfn98js7gDbuXkMrfJlXpqjKFB9NG2VQKUVben8BBUam+ku7l4QcPIX9myV4l
Z5g7aYegKgSSBLKniQOh72bYWXgJWnQgX5sSgxTGClAupmh2OnvratgEyhn/S2AH
FfycpCOq1SHBLUKGtlb/jN7YHAYmuEZ55pZXdtzdpDHFt7qwfQZkJE5GfZGDA+/N
g8aTqqM0xvlLM4AQkGL6RI2ayLbu/1oAIrhGlQNhQ9l9/3fQ7UkYtD1nLe5JJO5p
QTlqXV2QklQcwPf8WNB3hvKTzHhfo7ZBHSR5fdrCCq2wQJbSW+iYyIMlFNaS1PBa
zaM7fe1Y4YwVjN7oDzSzMAfyQ0H6NcZ+2PAVKgPYeNk=
`protect END_PROTECTED
