`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lhFDHYkCzjqLygn0g02/hn6H4XUM1o3aNFQjuSnogao7biU6ktY5Pz7PSsJVzCT0
UNqLm560WJ9CLkXfeEi/8se0+BXPizmQ5634+ZgEplvF99DcspDn6iLo05YoXTp0
lW5/jxUiVI1Wo1vVUfgDRz514G3u3Yv6s8a1unWdAViy4IEsLOAx4FdnEcxuwzIG
+uzbuvA8IA5/iNIkoAscTshJv9JjiHGnLpVKaa/Xj0Q8WctHjEKOvhIazikqx74V
ToycW3LYsWumHkwZUAjCmp/dlXu76aNFo6vrkVlnOodZUwItjhixWZtE2x/wbHLG
I9zBLd47zWIl7SsMY27fBLqFVio4/4VKQ3wtdFoHi6fg8R6qHzl7EBqKoM0NrxrD
QdcA9rsWns4jaYKlrIxQfbh2RhlU55+TBZk/hqIrHXzW+mQ4lM7MzZXQyxXD0PfJ
A32ULfK7nFc55mteB/7AqlUJpF2EwF5l2FVTIurTZAkikpAWgLJHBLgtg//qn+Pz
wPx1dQ5tAFdjt9z9EkR4VmZ58y04TyMWoJLUpC87mmQxoU/A8SHx8Sf9LftVGP4i
67Nouh5MZcmeePhYVOFr+Y+l0EfjYbJbZ7Cwmned9YcQCddy9GDYNawtSIiFobBG
TOwg8l2nRcwqiGhxQlxQ9pN7ayye5iS/8QbZpGsdt8VdTZ38ZXS5cn492ThankFN
JFmKvV/XJOb98N3aeLTRNiMQUnuwFCsKCOwignzxGsPTLvKswTreXdSsgbgAONdZ
J4YktPcJFMwSflNOiuJSs+sTe65iUlGO3Nr+MR0M83+BA25flpKLx64pnreQ7aQj
M+xaPXquGz4FiTdYeRsWIRkN6eEo1wzTsCUh4XNoqhoqfNOpRlN1AtqG0+SR9/B5
BJAd1pBV11jTG3HihWbXeXL/k9GupPFKBAFotgC35WXx6qglaym29Q/OCmKw+i8U
M3Je4jkN4PEjMAqxOMv8RL4XpzX384mmgSuVtnKHTGUFhipCwP0Yxj8dR0XRZB6y
r4OEKsJwSaEUbeUdFd54PkU23HZR4XCbYSNoTPUPaABuSMEKQKIqTBxOA0HZtJnT
RYWsg86Yh2ToR+2mLoHreV0emGJyVAlkcC+QCJs7z3i78M/2wDaUrTZ6ZlbxA/Cb
4j4+YIPBowVaafi3MXyUBx1YOlfD/KjSpa3eXs4yHrznKNuO56UZBntuFkOMUCwr
AsS1RCgygVxSBLSpl4DMggZcb7R40OXEyF8X7eTgsyToMle6IeBR67BN24XvVoob
MX+B1qPsn0Y+P3CmS3IkiCuph5mTE70q7+GY8xSHnfVkLjW5qmX7P1AKJHQaOG6J
AM6ywKMy6uFRcMBeVJRNuleOTp/EW7w2Ax3MlD0EP7y47eoozfVABtHH91Qewyrh
Cstz4s7HQs97VnesbSogoJ49gEdss3ld/w8ucI1sbcqGk+zON0b7LGKRgydDJ7O2
u7A+DPRc9c1UY2cPLmLKbDeRUVy5vMRhqzduqRUnXlM=
`protect END_PROTECTED
