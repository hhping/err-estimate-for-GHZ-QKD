`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zI/MgnONUMlf6LP6pi0odjOJariLeVM/Dc5v8ozmVVoxU4GIM64cpd5ZcP8MFBPR
IoSTDdxn5SkJxLxK3rrgQDZQHZpBXguga/kmxbAJsHTy0TM45YmHjAx0zxHjPyuM
HExdaKiE4cpbqKHUPLzS3k2ecJgA5wd66v96cEEnWLZ8hnfZSBqle9ecFHMoGv9Q
5Sb/41SVtIqL9le+Cy019yJhKkITWc/4WBSaQ6RvsolSe1UziaJH4dmEAdWlTjz7
0eeOuZFZrj/2M510KID2XJ2Gigs226je85IAZq8kcV1D/gzWNmFb2lBlSW7mGu/p
SR1sqpOl5kR9zhBZwIZX4unhP0lZcenUUXnFnP8AXq/8auxJjgp9/aDxlwaY09HD
HZ1YEgijbD0/OAHl9SsBdP99fnLdZ/fMYQ7wOtMGuZzNQtUxL85GkB7eft3SXzK3
94DNHMhaQMAnr2Ur1XqXo8uQcdc23LTODGx5/PKIhY5chJ0TctgAWvqTickKxHds
Kli9MQFyHQo3ll6eSK4m6C/6HFDRPp7o2+KnPZy9HWg1mBwjFloimtlXN32/Q9VT
6dXuwJd9oGmdrkAl6LPFNFMdS9mekrZ+rz5o9EwtvpQDXxoYkAAKv98kTBrxKZrP
SXL+r/o57/sQpjYebNRpnO8ggP1QgbKE/Z2Mq7luXDiZ+cQYyWHkFMd093UI4SuN
s/WVPbkbk4jJzSuPTt7PiJ+exoav3+QRkadLSYeDqZpICB2Y0ka72jxX1Kl/+YTK
`protect END_PROTECTED
