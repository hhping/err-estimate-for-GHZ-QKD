`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ze+27vR/mh+J0zgII4B1chMgJeQ9TTn7cKme0frVS6D/3DBjX+CBZQc9jTs3ZgmR
9k2nqpPKl9G/TKzottjwjSwfBRbg7OZ65XixbKUSWqxH/TK8XRD9V3KsTtyuRKnc
Na6EzQxaKU8QJQMQC7FMycte3T1liUMFmUvH03H2//dEhz3AqiXdxIyaysCCmjLS
XCillR14e2LQ0wuruCdyl3GYvT//5xnllKDQyrVMSsICD7Zun1AJF3a/2ddsLEiT
xIruGrYPtaFferQuTW/UpK/zufsBgvNRlA+xMZhjzTop3YMCLbkEQHYWdOiuJdJr
JaaiL4UBAUKsoXa6w9CD5LtFxxrXVp/g79ecA26Odaccu70NPpwutZ14MXzNF8Br
jOR/fjyzn2pvdj65cbZ9B+rybqDvpgCzb+nrk/26s4QXdxJUYeTRjSCyhulBQobi
2KD+WiB5TvAjY5635I1pt9ADtoIT99IvWAdSwXVEa9nqApgD8VzFJ5Tu+n0zwqac
E2FeUjPmIkhKv6wjFNyC5c80AELErVlhc6sjzP+2l0ztfTYEU450j/r12y65wwoH
s7SgyKLaY5hSA2uxmDFNg4XCqcXlA4z7/cpWAgNyrK/9H4PySrItCl+Sbp1kY1HC
fLXiMVODZMlbdwYMueDzdVdjKnK48QG+AR3UXqrCoy8xTp2pERGpsCNblt373Y3X
WVytDgqNvX20X6wqAcsZ09L8XbE+grcW3j38rdrgOqJEewI8/qvpujkoprqHc1DY
un2pX9QquosJxueBwM0CeXgf/P5pJYhfn8lmTelGTdhLFKD4Vr1vBPTD583hQBoW
SOhSCgOnF65cNKe/d9hldw==
`protect END_PROTECTED
