`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EK42BSPoZReQc+bxaQaV+nL4gh0yZEn7agAsY5koQn42LE/t45QPg5sBY3jArfed
qxADfp0UehPhQy5gYFLi9XJt116tkIrURegTdWOp+K+tXKZk7pPaHbQcLymffZt4
FY82Wgi78eKQ1lD2Yk8XsbRFIaxANhwY2MKzZFI5RgU3ZM8dTYQdDbJJpUyGUJw7
GL/GRWkbTdLBe5ZAm4zIXPw32FxUE0yVxVOlC07X0cXnRHbo4WWeVUtsN5OOEeIG
XEEuJwtnLsZBXF/OxAPxe9LBtyYCfy4YdbJDOgFKYy0UypW8btVhkewnlv9b+zzh
UZwqa2MG0joZ2EeiDh6Ue7cCVYQRqkIhK6Xo5WLwWLRBF6Q232TzCEPoUuKTP1Zf
tkglg7KkkvNRsttlyRpyD44aX5BDon0gaqIrifSzYicx4Pv1RJWXsD92yv5ctdX/
9KXUw0AArRLczZXqklCFCWbGpG2y6JfA/qH6HdmowNyxmbOC/74TWFwXPkYlyhv5
WXK/ANtg1Qx2QQnuodUch4sV2jlm7Op3wJ7pgNeusU4r4PPnZXs74IDgbcoElm3D
`protect END_PROTECTED
