`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
azIeNoO2fhC48ePFPyOmqV35ugLzSkQtpi6pa8CQjWE3RJFfnt9sZihKnPumXW6B
1JCHxqHYBW/8mNEczJ1bJ23u9qEbxWDHtpAEIq+cAcgoNegr6l3718+vJh1o4C37
s+rCW7ZODRyP6MD8eAFSGAky5a13M7CUd3w/GW4nxpNmUpL68DErsLFNXxKvlSJe
Mho7YzD9hUmfvsDSEssYw/QdgNHXWoiraougRDyP4XCgoEg7iZONlvu8VD6Ie8Eu
Btv7docKh9lb5NelM7v/mOO77kCT3We9tH6GgZQkTihi4IxQs7FV3YVLLQ+W9oXr
KoXR+rWSuFmpoCZKFN2SIJZbRoWXBKVX82hCssw/F26Vu9ME9rPASt3hkppP4gX8
BWrZ3kcX6lT5RPgU6MeFXmsHy1CeQDSgprUMMM8pattOi3NNL++S5FyKQXvhWqwK
lRk0s5/8XVMaMSmAb41XjamN9/tf9HrUscKNMSgkL6sp0bwCD4gfS6K5WHKqO014
3Tz2Dg/4dEfyQGuMHznYgGRTC4XT7WpzKAgJ9rU1XX24d4XkJAjxDT14MA69QoPI
SHJgzy2favfiSnc2TH+T6LZmcNHpgoPHwrHMRQenhyaOzlI/LycbItjNi29oIfrG
gLW/igw2PsphoYbGC3c/hNjo+Fdjmc4kJSFZvKsAiAoSM9UyqYeiKxQFEiEnoZ0K
/w1S8DhUd+1Np4Sxkq9/ZJraqYabF36959rL33hk941wqXbsMzYvDMeSAC/kx/ut
mKG6qOuC0uC4jOLZrNzG/hsIp+oFTfP7ReEHX+qQkw/UKZd/dLpoJIIS8+ElKsDP
RFWMqcEwDtPeQgFO6d0rSk4AaX8t3FOJ4BkXoEFe7wz8bre55LS1C1Nav15DF5qj
EHw4TAtQ+Iq/z0RrTR1uvo4v8DEbDfITnKP63it5JmgO20F6E8z+cZM/5UnIIajB
eq23+J4/SUY5arbbcaSd1zqHFp1ngpQE7oH47ogYnokrn8hGt3rXzYNejtS2atXa
aKQ9USOlZHM0SbMEi1urTF/HRpQCTyZqaywrnRKx3pMuFq4zsJI1UzqYxGe+M8AQ
e5IVpvPVDGjNpzkFOAbpCvwu1t5k9eveYXP5yYeNRp9fRhOQxMHogHqMBIjRwUbF
hlrkDnVGCDVJm8N7IFuybRC2hqpVE1hjeClxZjRxTc7HG1EDbARp+LqlGN1IYYfD
5nS6H8o7wGNkj7nrnnqY9dFslUnF1NQFtEQRSWCvrRBK38l1p0qAVv95RG/rdzgb
apPIzzA95IYUikbcfcxASeiunE4Ft8zFkNBsYxXdKq/WC6nEL8YpKe8QNqXBee7S
hS73zmihGSJPJG+F9atSvbBPqITeRQiDFSmQjsjCrbn3S5U5HE0bkkPl7330r4nQ
NRcqbS68eX0DE+lWQ2XcQOLMGRuxIfwoqycP8PtPqw9kP8wHXqUxF0KLoqyZ0h/Z
0mkjOICG0MmWiQK9d3ZEOhGYd5S9/gJ2xUYfgKTAo+AyD6j77gNPR0+8qlaqAhV8
lhn301tvu5PWl2cbfEybWSTfewg1HWl0o++LZhXCjMwZ6SWDji+gESa5q4gvGyQP
7cKhWpR/MZ0P8vsNTi0ldlCrV/E+pCI3GuBqAVxHKoRN0z9TXsTKwK+RrrQw9QoT
bv+Ei8y6/WSraxh+fpIPVF2g4trQ/adAyFspZezIHEv7IUhvM62Ve+0P/YN6v5LU
xKbwChyk2htQVMhHbZ0sH1QqctV9xxXcHJW6SFvfNeNpf02yJzAJn8CdQVuZUpIx
SstnQSQpG+/u2uIyrbhKy008A1VBg7Z7Q4n9Aq5QdzTSz4kW28BtBKHeMP/pgh6c
WjH79o9CBAtOsc5lN5lNH/5NKUCvnLgpizGZ2DWq+FMwxDzlKMgjRvixfSxvBCH4
hL3fezy/BBaB8J1YemQlb6A8/I+INLJyJk+F70axP0VUmxZ8+lgUFvemoy+QIqfk
FgYnYibO7/CBbAPIUSnicGZKUlEuzk2GKmPbnFEvWVK/NgwvX9XBbmGjGMQfaBKU
cuGdbH8eOD/dy1O2t0Hb9BMnJ8lLs0939iyJ4u/e9bQQXxPxdtlFeZn+L4xse5IL
KogAvYSNJrqPYp1lKCUIbCA/DFBW1x5iJfcTyxh3dhDnUnRvX0Hzbu5jkKmi3F2H
uugYygycwliKmBLWRUsjjA==
`protect END_PROTECTED
