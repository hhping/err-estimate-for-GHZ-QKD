`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H082Avtgp8TrIgao8Bm+osDkKtpmsmEHIpRpL7DjlUYDHFZM7u5wPLM80sWTv3CU
A9e5KwM1ewmtEHksFEwiTkUePtD7ECxwgeOq+CVrEIgpENkLzOmiHdKuoVXB6OMi
SRBgyMxL++kPf3KM+1wefgvopkLCdY7OPihf2rH+/yOxH+hOiPPOMCDRixaxq5xe
hfO+CqedlXf47F76zO5gdTpDZzNT3XQjC8tcHGsfs3BPgK035XvTECCwi7BD0XDS
BNpn2HYDdOq/5qxCdraFZiGcFUlJWVw2sboehqQyuEVpojjI1DAqHNNmxMlMAtHd
mK5I1aw+tHWjuge/49pnn4Xs2VgoFNck4KTfG8GU0jDU7/NvDVmqL4iEXLV20Y7U
5qgOGEiYFN7koY3TZsIlKvGtdH3zwJswMrkQbe1fNfyiV8m7MRzWg33QJ8mcsKcw
r1ipRhmIc7m5tpIOsGx/dzM/+4mOHan5Uikck6fozSjJEG3OT0Rc0VEwfIFqdiSa
TS8VnHdNhzDDKhIEumaq3egGCIzziPKIMchhtnBY1Hc2scD69zbGIxQxmBWmuLV7
YWAUrdGIoM/gOd6CvYCvgKaoL0T4+pQ1qZf4xa453xenAAdJ1c1w03NpJr6YurfP
lCthgsjqD+Mu9/MiUho/Wb8/CZItD+svCba+z5pu6fBgi4L6QjF0yzMSUQD/aPqv
AWBcP/qfGUt1hc9MlWy66O3u3X6iMCvKBXMW0Bx7TIyzFFZsMvcH/rB/uLrvtmH0
qiR0FRx0kHqaNQKwdzkaPTueYXvwOJG8pfb4bPpGqHZ6X+FXgdSfYsEDIpBiuiaI
+YKUlhh6sasgW5JijLmDQYaP0a09hKXmVcgF5Ry0tIWrIWjcT9yjHUgFnQjVSeEh
waXHQPX/e20Nl7M5uuEMBrIKxxbz9+oKilLWSWwvWpRmGTGo+dSUTgLFR2g8gX3a
djxfGcAYzh/EF+gn9f6tZcuXP0Ju3Enm9Q+twEhYxAUJwAV6Yc2FfSJL4Mt/2XXe
e9gRhYg6a95VtVcGm4DENWdBquxFfDDY2Jg42320IJZfvJbHYzKcE7sid3jEf9r2
QQ3z6cpXZ0FefUgboZ22eMrKE6ZvslfKA+cUZQLa4BODgcRLb4nbiywE3JRgENie
lPARErdaCcB58ZWildFFmqjHc3msVaSInoQ+HNhI+A0BXJaor0Wv8yLuzPlOC2fF
GtiALRJTWBRH5nqJCVSdkf4aB1TxYDNP912mMRfirraHSXZClCtlhRKC2OFQnAJ+
srTOTtyYXp6/fmneZhYGRPJLqnGccBwS65hAK0uXJcir85FbIwjiqtJA7yo6WuT2
9BL/ENGO72AZXlBupUfHqECTsXFXCJNfQrqcphBRcvKe3MUSCWLUib2KVAzglSCn
WzgEhoT1F1k2sJm+y3764UMmQI9AoiKwM5zzldCdn2ZREij/q16sykEUk7SvRrVN
rI+/NRbtIkfhTQesAVPX7UaAlo8SCQ9BzOBDCnwS2CFHH8bGeMm5tDuThaRvpfMC
SDwvvYyFCDOpsop6TxwCw2Euks/Rqn29zZo1/wBOR/gHMTitYcYDXVjL5QOosBT0
pM1wk6+9BR9IXMtK5xste/gkFmvIz7q/za+YDOix1rH/vobI8pQkx3BGjlc3cQla
Ng5N3IQAq3myxH0wOGc9jBROHThYN+a1xbZYzF9q4ykrILdd0Evk159BKbT/xaFx
`protect END_PROTECTED
