`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qs1W4CO3qcxNIF4taPC1cTYzYv/vq3qfFqK29/ohgTxKuCoqwyfV6/bbjYfxjkgd
xk7EP4fr8Pt6RT4ac/Drepq3CBIj81hbrpa87T73Y9WQXkHq7nL9iEYXSFdtKpQz
5eHxgk0m/9Mvm2cY9pP1kyB4coA85u+OX3Lryywnucojk7ZVa1p6d5PbQMN+vmyU
c4DtnGheC07tHBqxmReZpsAh8EbJOMibv43EYkx/J+/iYLUaVV22tcb3MCzaLkCK
h2RrPaIQPLaqM6sI7Ln0jT+hfX7vo7c7mAmJFvQRgM8e3Ndbcohc1iITJAnpvI6T
cS5TAu1ZdJCFR5yBB4N+bteoCNs0fSuYvsGKtL00DIejlEDZOKkLfUEe6IOAQfoX
13sWEiAaDEFKVhHgh9cXfPbdb02cVfH8ZOtvl+iOFB0KANgpIQi/L3A4Xv/t44/7
FLr+3bEVPikv+YNtdUsdKklqkT9ymeeBYa1IO0e6XyTwNdhL/jjskZ61fSFKhAVZ
JziPbVJec+7w+W9y+n7AfQ2flp0S9mZP+o+TmALDqUZPjaenvgbZvhwCZf3NN+OT
HOqYOJESGzoQICrtSgATVhOrkU2QfqrV7EvUdQVegrRjBvdWI2lehsUEH+YUQLrw
+sJEZSjA57cU45tQyYvCLVVURmdVd4TQa7atk52D10DLeZhmLVc6UDPEmwYiSbJa
6CjekJDdRxlfeHUd0myLmxUIvYqqdqvCQ/og1YizPdDbrNQ42dM3OUS/VpXA7aY/
mIosAqDhQpOxBR1O27YoL6KaEPZ+d8oaCpL8hVJ50TVTawobyAxps8iNWfWvi5A7
1z5uTxsTwQN9XVFKi6WUO0wzCB1BLlE57SFNY0eJl5O0w5gIRsxBgwglsQi4tYzq
tPt1hTXJWISyhbu0At0zFBP9Bu6yCTFM05yYRGgdoBBpEx1rVHejSciYIqKA3oKc
`protect END_PROTECTED
