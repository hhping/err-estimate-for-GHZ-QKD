`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EwSV3Yivrn4Scfb54bebYv0SIK6xYsDND/k0SsVaXvfYDOU5uyfJov1K9/ZIAKJ9
SFwR/Ab+w9VV6rNyBxcTZMPIuAB76BHOv37TC9nGsr/MBwGAsmDXukfkQ3D6Lk5H
ucUe0lKtY7gflJPEfgfCzzkoEDwxG4d6D15RkmGccfUTYioMkgBsTgw+51nt1tyf
WkDiwnaX6UKN0MK500mNh9Orkoq1MQPPWsXRa8Q5lHH7Z8HbkRutBbdidDFcCCt5
3KpifsSi8QUZZBrgKwDrdLlpi+Q9gierL8mqANBD2ldW9LH9ANr3LlKGFqMFQM/R
VvMz2hF76D47/InU6Co5Vb45Tav5AjsmnUtnW3RULTlFRGCJvQbGtuaPG+ajCqPL
g8rUNyzq/ipCrYnxAxOBlHmBdDF0Z06V+ijkqo5BjgAI4GGZoYI9JpaHSIwmHmas
CIls00RG3bwxczM3XBOOX6cPpB0BhrCFy1Jz+CPaPaElwoxTPq8vZRGOH4sa3HkC
kIHtQXzSsPemQaTyZwkGN3p8uXKY5DsQ8BTDp32+rNiTkHagrIoR0hdm29VGLNpq
hoglVtmjMkWuwxckS+Wm9+WaMH4o8vrxOHOOPnOyELM4MFQmDsrLjXRUFl/7ojVg
`protect END_PROTECTED
