`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97YZunzrclDa0Gpl4lbwaIiji6GCIbpTOlA4azE7VcsvSpUPDtqlNM8K+SDaB0O8
G5+GdJgW2BOu/HysrumlY8o4Z/HgeVSi6399elo3Fc1zCIJa0dU7WTF1cNAhrUFQ
OR9m37Y7kaVEGOkYEtZbt89NjnT2krhBkdONoAgJu6I9bc+yWRJfWlSR2YlsFyu0
/uChbCisYjoGsmLjm4v6YQ5cIyt/4GzepYA/NuCxYauKDshJlMDqBICwt7MY7POi
EC/F5ndW8ApVxugUi2FiFk9YdWQAF+nXr4wKi49gZZHCNvfQ/dOv1iaIAabRpzCI
cmrp6qhrRgtEaFzn1Lysp2gciGovA4t3vIn+vJTKGO0FL9gFEjDVFtGRoIIywex7
SiwmrE8Ke/gUiZwRAorZDdrjokNtlHMXlXrk7Ju+RP5ebcnFS7gsljJVZ3DHXJbj
Bd7oEBjsY4jSu2M2/U1jis46H4ug2Y1QGxB12LPwF0eq9+jWikIDtUa3e4kNRdSV
9TZ5yd+J9dK5/8beZ/1U0YApOfEqBIcYSBSm6CgVXI0cUPTDBn2smFEXndnzfB5M
`protect END_PROTECTED
