`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+qud3hl1c1WKKLJ4ZW0PlYEP+j6AyaC20v1ncaipkqlJu1zQ0MU1A/MtsuNTvHbw
AnAWRKJU+fRunI+lSHwmxnxe7fdrTLU4se8cqfPKqZRbKI+AHrAD39nIn1olxwwD
FG16Tf8LvMXevDVUY/gcZoioHrDNrE13MmTI1ifzvrlMEGouHQ6qaC7XKiFpDu3l
vXju5S8T9BiVJAYk8XYPPdQU1J4Ma8zMgX70zAzNIUHTKwOdo73skDKglT5tvf+F
E+Xfqzi2HlBcn1m7AbajsNWcF3lY+CcMXDzvQGc8GeHeTPbg/kwnNDiZw5iWGkpe
lyvQ3E/5eJqqS9Isb5ox4jNNnbQHLvUIbcoWkFXo/ZSAB8rShcAh9rz0qWBzwsvl
cjLdw1AXvnbBRcy7dmRuMbsjmL8rtKYUPmmfXjD1DfvkOntB/HdQBQJ4r4UADkQI
TvNQJZ1RTij3v/MsgW+MXov7i92Nu5vnqNrnFXXLHtQH4Org4srNooqlBIFs9feZ
nVRWZL4OmjD6xgnlqrVs2ToSCmpCEeiwzQ2rH60BRmYPWKmwoeoqTi6T2KV2Hhi+
nv3y1D0nxCjagLGTnDOPA4MAe+bHPmWlyeOWlBry5ArYwEJiW9BDUbopiK4PKrP5
8I+JiPqr4rzc9pnbBvaYWMGv7A7ZI28sFo63BZ5MyitdLiL5TM8M00H/oVFHaOIn
rS2Vb0LmP87nXtA8WnMiionuOox/LWxdm++donOIXiffNm4UOJAU1hwTRp/qdgZy
tQCh+CKWd3cmY9GIwKlDYThM55GoeMeRNGkH/H0AXCFC0k/RZ+9XHpqKCKAyBx8l
1b58AmgUHR7S1sPceQG2fw==
`protect END_PROTECTED
