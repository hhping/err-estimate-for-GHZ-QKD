`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+A/rpxDw93h+nKL8EK5rx7hyQkV136jRPklBXH2katG+s3kjsyp432M5ccVsSpCb
injfsyECTRIJcGt8d6X+bjUoUpCU+2BkeqE7tWU9nCQ+ZT0HBN9gqaoQGuSjwK/1
Fq1vYHKiPq07GrmYZxrRtdNwhZx3VwmqZzFgCxLkxEf/r2A3wiauW181aiZ07Fws
ot/5YfNITH0lnCD0hLICaNB3K2bpD6Viklo3InorNLsvfErgdiqWyGcWlr5H7afQ
hKJ2+9T+kqb7AXWSFji28Xka39gFnYbmVZ2GiOKhFAW1qpKiiZ0Bp5274YqmuiHT
h+tCszasveyUFOwxLQ0Kd28aG/pte1QflofsS9S3lt4xuS3TeDZNZDCJl8yDgNKa
yM875qPC/MnBZKoSS5lAaWQ8LBaBPBTVqgzft2ZMdmfEifSts44GXijibLYg3CCq
Th2UYW9kUZ1nrTBpEmbdp6l4rJAbqbxMNEdiWiNAKxXCYxsIbi6ZKPfx+pYCgqas
kwNwCxCorWSY2EQBeUqI1S5e1bhu0jflNSJgma/mnNY=
`protect END_PROTECTED
