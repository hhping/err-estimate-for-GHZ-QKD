`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kjx8xJPksxc3tbHg7WaYBedSVjZ64h2IdjxAMl4b8jG8Nc1miB4R8HekWNEbA+cQ
Grv29jy1QnjQ/BhZyVKGM9SIx/EQBdoEhBr6lX6IX64bGNByoKZP0tJmIoV2pF+B
Vz+JVBkg9zzwPAUrh9GQlsko0gFmk4viDuSANkUaeFBytVXnRVyoE8SZvGGgaBac
3lyFGpGQ+MH4IdUU3qjPdGzx8B43xCzxWnwzURx6Ux3w2rhwuXzDD9iTDs38yGq7
zarXlsbGh1rU06M5LeE2YixV12GRILFWU6mtTC9VFvzEfxY98aK0HguDDUjEDDv/
2LXTIBbDGnNbNhjIlK5WBsyUBxJNSGRtkuVbm9EbSJMD4kUUnMJIZ3f0dS09gg9i
x38r7E3vX7XxJ9gp6gZL8i6SGvloffJCH0E4/g5zIODH7VWkCZEIJ7iKgeGxYSPa
52bwYj57eNXlUqp7kKALs2PoLA7WTh2kZ0RrquEQgU0YoOeU1wsGmnhDWIcRUs2J
UYaisG1q/E4gOHOQN/1UNfDTHMaX9AluVDl3rAjjOQfpHAnel93FIRrtiL0Crfy3
66ptKbb2zuBWo+5tD58NKiidkJ6JrmzJyUQDT5mh+G7FJUjX2s12Q8ueuWiXshph
CFevK1z7/brn6r17cqSinvDSeNP28/4oaQxUw1phekbDYl+5IQ6Sf23+ly+nKDgd
eEQEUuv3jSTxWQy9hy8K4NTQxYWtcTbWppEDbQT7Q9UdppKmvJn/+LytoMBiaxw5
MBhTOFzEwoyfV6WzEFbY+ExJ8oo5wi0cZSWGOUMEfD5Jl25BN0Qt4MgInTpKHopE
O9fVU2OWakf20ccJ6JyfpLthkbZxE3jNFoz7Dr2Svc5PlbdljKM8GkYcTku71yak
vZTDS/K8j7lHP5KTVvyPk8MLfpI9jDEHRM3tpZMkIgSP8m/h3q+F6kB2vyyEaRx8
OZj4WKk2pds0Kd3v+U25nW28gv1Ze6D+K2s6mlMnMMY8wh3BFjv5WL7aSEFW2Lv9
ZpgIk/wLTS/YZTc+XUlnDvKR42q2TDxfD010BZ1ccgU6EP6/ifg6bQs766G1LCTx
5pTK6TN3TQWwUWtuO7dUPpPOShpyu2AMLaVyjNEiFNluMaVS55aJmN4xMsu9bwyh
0BaUc/McIAjEy5LQ3AqD4qqwbJYlrDO5HTeyP3K8fxeLau99JankeppeZUwgR+/K
Q1XxCW2NqucR8fub+8QWF1Ixo0JlPQ9LnSiJHGoUKEr1Y/YrsKf5PaNTQ/B+/FXy
Xu+/3YXT4Tj/pbkAuU5i9ABcHDHrBGUZhnI0vz3LdMw9xbnk2GUDUMa8wT5fMAIv
2eAlPvLnWuX1g43tRqJ+dQCUeGj7Taiu+FxCcDJ6d8wTpvfvmHeZJ4YxFXpzWsar
pp58Vgi6ezqNfDSob4qa11bYQMovSQNIpeTWDRLOqmkur5vtKji3A/70bbfgHbpn
sNUHnifDsN++fsA4ovrOGgUnXD8ijkCYwlUzSNAofkWmAgo4t08Kq34N1JKYDN5q
GMlwevbdO2BHst1Y5veW33ws/f5rvWAHIUsrmD/35tVHT/yJzJhcmWxfECN1se6o
1gW+mTMd8IsNm0+sQFtLs0Ku1FFzc7BE4SewToznrAeMcQp9NhTHOIAlMamSCxnN
eHoS5H8sCyaog3y74r1cdZF8YlZjCRmFOFb7HmHP2HTqvIZoKv3Tz++3RoHHFuvG
e6BOzTPQQ3ctWB0/jQFt40Gk7Bn+6Y7NhslZVdQWWx3dj193zdo+mbksMU3WK1tJ
4yNrtDVkuTW/Vnb0AQukhbXfiG6w6mG/PVW+9sBRy6upZ9yzj+X9xH+DVfaAGcDF
LLS9iJaGas4RrRPrzSXU01O1ul05GqjCY4sgovES5Yo=
`protect END_PROTECTED
