`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3sA+zMdWQ0qZlz488G7C6wP7b1oyUZRbG8slfNBwPa19H3E6nAbNsBDucLIFHdN
IcZaGu6Ono2tGLRUjn4gSsjAA6W6aCxyYBn4MdrzLyUH0eqNxS/L6chMKci7V5fF
jAnWsMoUkB6LyUCZVbg8KyHVNuRj8yOD9MpUsVl2z6s3+e0oGipJ79jDDxlURuM0
rvFRXsLEwfHHv3F6zGmknLnoiXqqoq0Wl+2oOkov4piWdpopSq+1SIilNB2a0N6i
9kid8NNrAOsYRMQBbQ70uartfN0JOpXcx4LRMgvWQmcyDB89GeEDLgJbGX6mCvCq
aQGtsc4Hm2fEobgKkizW/iE4T/VChtDEheB4rWIxl4xnAzxBjuoDrrrU9LroJEGb
KyXQIRnHyS6Wj+28LkGOCnN/baIstpc7lYxJ6WQh235GrnxvKjjQyNmVlS4K3oaE
HQJTCEqPjBFDjZjUoNpRSvKh3SpjZ4XCxzdmPiqTlfoGbz4LBd88x+eX+FUqhvEl
RzODCXP03uOIrD2bPbV7rHumZElD2T7hNDnYFEyRaGoYm3XJkmkRXX71/q6kFUSx
YN7VkAa+048EeZSjYVcjVQ/B5Mdm3+B+9KUUENZux1vcXT8RrGUE766EJgbkv91L
gvUhY+ganw9aIkLpzXAScW5qglP7q0ZAx2YqYOxR47kDsFgMBwN+CcGR4JAOYUSr
ojxBd4ICiMkjjwL5DrUu4hcmzza8LfqGv8muYfHQk9mz1IznWngaLOQeMHy3ji3Z
Gfopr7fm99WGqQbNimJkhMNP/k/ki//yaM++j3DmUvwluHsJSgvtB4hPwp1SbFAS
Qmwc4NWri8+gbIdtczzg+PnCbXe30nvtreHtsK3CYMWX+Oegokj1QjFYJJ6M5VVS
bJLCrq8w8KAB3kCMgz6v9Bc4L122fiJbz+cU6l2DjPMMkQXCAYPC9AKuSi45jM4X
PxiOR/1OcTANdFOl1GOszGSOv/BFZ53m5j0fV30TND1DmMQERn9q4+hklpEFKx0b
rANHgtV3BMMF8Poh5o5xKN0tkl4NczWleQEW1T8wbOdllwKIPrmzUzM9FqC9g8ZX
TKlsjJAPe+Ki0UOC26a25XjILu9uwM32aWV/IyuZymk7zjsBl5On+LQOnsp5p8M2
htbnvKGd8ijEyeUgYWc7PWmYc8pI8GEM20yPxg4VuE9x3SLF1cuhrmDSugINW7L5
HW/tOKld4Ti/D1/dJGddjhSdO267Ro9Zec7TofFEPkcg3pEM+DURuF+Q+WEIaoSY
1sa+xiw3dJWCN6MVRfQIA9HHz6j/VrQJLhlE6kAsI068lBPI3s39F0JRK3kFgYib
+hOskLGkoGcFdA0WsUT+wgSa4pbklgQFFkg7FIaP31z9TQKB0IWUO1cBtmcpYpPZ
Lpv7qHgy0CTbLTgNSfKCylHpwBAgNJZ6qIDALAFK83KQ6spd+btWA73SOB0OyDKf
NFlMyGBjAfA9fEnLfKCK/UjyDQHS8+SQDoW0ZC1NZLtw/EITUXqv3a+7XUXUTHFU
fdz2U8manRZCZ9UAujXCJIpfkW/w+R+ySlyDITNkJeV5ax/MqWXO4TilaMPkoTTt
zBUDbczrhS7cQdz0X/HPd/F9muX7XO6OZRTKWBOYJbN9zYn+R6KGy1UlKHzc1U0I
dOq/q2GhP95ORYUzN8cYpirwSNcbVBmjWxiASp9mRgDe2hpWqot6U3kBRcIdz4ZX
xwd8Lkg6P14kxb92LFnH7rfOIwI3O2t2cWOYHxs1ff/eZffox1zXc1LvtQ00rsTI
k2gLXputtqWNK5H84v9qce14cjdEUujR7GdHOOD/FGhknncXbckkVkQztcGV7NJD
yO3WhyVeh+LTgfOwNQpmsIvgafMVIrH0ToxqOzERKET2mWryMdWtxl+nZC+inQwl
TISozIRMWh8ErY2tCnu5YxJwL5PfSIZ0Hq1IE/DZ5HtVPXwJVypPL6L+fxbKtHex
J40t0ZqEQz2Kf/Cw7OdZehFRvaaotHn177KS04tG4y3uH3AdaiJhuk6ujZCkO6f5
hqj6YkWFE4nOGHa9KjApvku+8cKbI6WlEiOFEnLLqcxjqQCBosn56y83E6kV1IhE
1Jj5v+6bwuyX2u/dlAoyYVVVojew8U4Dqxk0JM1wkeojBI+bX9BsG+1GkX0jAMoD
5Ex0k50UdXdqYswVw1cJ2e2VtsOSoKuAXjNIBPZ/Bt6sKDvpKFHt1e9dalzwUz2f
wiN4yXDjvc4baHNHwdXrE7t8TEN5nwH0l3WHewELaREfWfCcWDBv0IuU97qkzNcs
zK3FuGXP2AyIZF6/eAjnWgaRWXWhLX4OW2G1Cc9FMGi5szNttFwqifREfPAJfD6M
hXuBlWVnYulXTN61NyNeIZ9pIyj7jDaDv6Qs0L5bQHBPYKWPjb9PaDRlkEHj4p7H
wlFde8zxyzhhwHAjNjHshEckX2GEfuuhxhP5PoSC4SN+R2pcPXTHXmofuKoCZF/z
11kWxvx8zZm/P8omoFq5wssvgIOkNMU4fMpxNlBG8bO7ZMa7Dd0iyHpPqzlMtlqB
yCOmVSP1ittgX0Hj87k0+92PVr60MEySNxjRNEsebAO4qbPyqCTK86LwynpGB0SB
Y3RTOgAqYS8W7ju6Ux9TaDlew0bnEO/VQMCV1eWKTOvNob8nhASgwLvnnwNa2bBW
PS/FzDw3YNA6gPF8vW0xLr7y7w3BBp6hwN0/a4ncRfN5rlC6VwBGWvtiETFZnodN
cnEHZaapiJCRDCf3aFSw539F9rVHeRLT6DVDSp3MwPwhFS99n/i+OWjZHCqwkFYm
9s3rkDTNS1lnXhRZepwvuAGU9xIvwSCh1Iihw8Sjogk5P8Z5xcW9jmumjq7QwN7I
9mn4NJJ+KdXBRmIZIYiD1NCxYYj8Nu1eRZkcCTYsACZw0f33GRnhvO6AzdzlNM4r
SRGng4s+FWWz0lVtdDbBC4s9KxVT/+pcbn+FG6AZsGDgtJgkdR2SD1lo4vz/CwMb
9hhTho9tBwRLw6nyAIQZqBiMhiM83gEG0FdTZElU6lkvvBd2tpTiuhTMjn590Eri
X0j+dCgqc7d3RI8jcDd9YpyXIHOSkuAB2KpExsus+/OV+umdUoNdgFORZ8fp9yBD
OByxtN6twv2vi6Bqyps8+E7DJWZARtAEnK9MtSzYyahmn6uVZBeM0cnUAFLXHVQp
KX6Uz06HjNp7DJqNtxpipkjGNeUEBEYjcftz2Ajw7M7bXXiQ9Dtqc8PFv7g4eMR9
ethWmt1Zuj9bfuKJurB9CcJVa1CD1Nq9Jz5eDwNynQsMXwlO3g4LMTfKAlqA7y1i
5xsIU3J04CX4XHb/wwF4qDltPrq7uaED8qmt8c5rF8Pau/2XWvDzGney5ldj/XOX
8YJX5nP0CZdnmGeH/idWwKfhmCy8+dVWag21QKo+bRl05uQpK3CSNUhcctJigEhi
zhYn6bci+d3jrUjsClagug==
`protect END_PROTECTED
