`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3ZcpaIdnU1X08PsKFu7TP3jf4sqBF68pdvrR4/lKoTF4JkVf3bBxr7TcYWJyoPx
FNBIj6fB4OzeTX1walmOBAjMQpHJtH1LWnzExOh7Ihm0/+C9hqZhG6tlUuOjuc/I
v9QZNEoGUHReq1DkcDEAw4GjlXHa4nXGgSx1w9S4AEa323AqI71Bmq2hTZu0eplm
Z9CDAKNU7ng1FuPnGsQMvv3F10kL/QGdI8Iveb+3gu0ARgNF8xnjYoXc4tHgUfNV
vv4mFjl3y9D7jb+sJujxpXovicSiIjGQOMCsaw90ibHmTIC0r5GIhuR0ekpmKv7k
FuGg95xlgs1GsM7d6Bq3c0P7vskrSxenz+TshjIeyWSavC8BLo2E7YvrYlGT1LOV
2z+jG+bWlYnknBDHW92hM/V91qRDc+0durpuyqdJipMcSeO6P03gpwDerF6ZPGXB
fT/WtUIhzO2oT/tQdJMgoE0/HSogawciF+y2zBo08yb1IIy2/ioJmfYIR4LwgTyW
KR69AjbiRIsSpsFhr6ez3ZC8EfbraeTjryqJ3XJy9gpGzBiMnwTCWnanp33cTfZz
0OEgJhuHss8z8Usp6IoNk0ZaxqZADpQsNC42RYKPTogO/vO8hl5kAaWBtV5seBsO
Zi2Kn2PN58Tz5WOkphgKFUBxjH620r9sOUoMrYsOnJiH9w9FQd+vmxPmu9Tk0l8X
1a8j4o+ovAuXeDERkJ5S5Dg2UR9WJvIAvJQbK9xPe75BxioLaUXg3aLoEx6nuEoC
OfPUrwVZAj2tC88CmAIMg6wvmnCBjCjnaWtyOH5QMkr4ZnI44BZqEqEf0pUAuDB6
dJd0sCxYYw3wWIb2TGzeemyWlTu4F5nE5XsxD3nQQldgnPk0Y9NSZyJKBJ1/Mcol
JtQ75dRR9nXBxhk9NIyAb9qzhxJ7j3gorBRWS1+5rFDzrR0oKcC85qfaifgcKF8M
URbj4czX4O0Xi7M6AxXkxfxlsYdOzfnTF1azWUhHNJsbrQbWofGh3GnBA88xIE0u
vl7jWmGJpKZpufZ+WbVwz4Syt+1SLeGVnjagZA5ROQP8hB7+e29m+unMXsWgDvNh
k/+DuDbKbhpHrxPhvUY4XbLC7iPRLWHl0rWPraMOC3GmC7IMIgqAxocH8fx4sXP9
pGjL8QY8OBCukHToMF3hA5lh7xidPpmdvgyWkpBTT70TmOpUK3sFGOR5l9COSdWU
4RGcmdayZFduLdek7275d3JiYQyenvb0hEH9LpkkjofTE9jMQg+3YwzEq3Safmct
Ywf7i3ttrFr7PWya7R48BUfIZTpA1PaFwYDYSYfwtiJbDYLOD1y5jQ31F94cnJAE
wy0w0CIe8td53V6kpBIlHORtCRruxkCIAJu/U7mhPLZzQo242BYlHz4DsYw4x7Q8
tAaHIOcJO49LEQ0HLkZqyxYDkZsYFHaFXdB870WEelNVNDHkGJRS5oNV09eKdnC8
0uDVCVJp7pierMmm+Qe5ZmIwQAstwm9OpF1X6XZJnCHsM2dDOdA7NQt6yP0lgv/g
lQ2eX9D4y71nKbRDXYiH8nmUGFD9eWnx0bPmva1cUFxmzxEPaAiA9dz1zN9WMd6P
CVYwz+0wZiwT+Wysp+n1wbHhXgtqVmQJJqS+NBwxTOY0W8rAmgxHHflYuZZd1eze
wIgmN9uFuNcOE8PcCXrqBcoi/URa8escrLUuprv0BbQbD8xCyAD9X0Y0/7MzO/Dz
w+y9f6HhVkZY9J4Ib2yPknVGyajn8nf93+IY4R+MfYt6Uz5+NYyd3XDP0D3Txf4g
1PrxbTeMf1uK+nPgpFo+Rxw5hylibngTlD6hbZr/Hxif39ZEewNOStbjH4NFlpeE
lZTi62O9p+bfWeazdvIYpOtcf12uFlCd8GSuPE1emWbLwWW/G9/9X/thNBaEpIKn
Xy890ef9mMGp7+OsSLTJYG3c2R4ZSwBGbbtiIbqvH1cioLuSeNeA9HQ884oQqKLH
fZ4SvsobgIsHh1I9pLCTWFqFZXJn8NRIeJcb05FQzuqsUa2U36VyCwCLA3rbPn8h
qhgz8Dzrc9QaD4X/BlNCFbN3RNlCsaUpT/AV8JF4ASnk5959Zb9Dwo7h41GwwPq9
pTIqys+YszdZ8kSXdqYMu3JwW+Kg0p4em5LmHz9GQot0ibL1auUOrnqpRlC6ojK/
GOn4IVJEDpFFb1u/X0AU35UAwT0fJ7Z3vUg1JYRwajxLWZnh4LPlkKUD88avhVFj
sKioT5nc/+igEi9tX4Ha+g3u3PV+uEzhvZdyBdsx/qLKHjsJNmxlNsoEbIMo3Km4
96hX0MMhmnE9lYE+12TcqpzTAePygkHEiZ/UCKqTqUj6jBrsQkpnUH1VuJBgknyq
IQKWLqTh90bKMdAvanDRIUFhpxg2g058ZEh3GtTRGDoMttq0/0hnYId9sz9nS3kP
//uedzR+jLUipneO2T5u/FWgbE/1e6nd6u6rNDrkcBsyMlrmBNls4n1+F5ft9PiY
lwrZ4CqHfRm3TSs1Vah2UNU3Wz/uyjELnN/zLHE03y7P8vrnGkaT0qz+wBYujK95
ofrN8birB/sqRG1xvpmVxbTd7UasqvrkMEHJtcCH6ptutovpkunbPoVOcDytd9TM
q0/QC6aT56jVIFb60TYqbgEzynwQhb7QZhj8kUe3hGu3z+uD5/V/PthRf43EAf6B
ZNUe52vQRNjFhpyN5qedj/nuD7/gdlgri9nXj1o3XW3nGZ+bc6/ADvHt7Yy6Aiit
H2EiqOCutMVkgUABdKo3L9hufi3bvw8CQVeByUNuhnYVqZAI9aFhETAG07z6LdOW
ieKu0VdjlseF5pkMdeJNsr8Tt8XyjY+y3Z/SvvCnAHAMnoez17i9fYp4OeYY9rhw
l7CmVSmEBlfidV8FmtWdJcAs3sYhccGwrZCW57YraGlQTQQN+wrIWcJPAtX+rvMZ
UxhsX00s1Uhp5e1+44iDtateDi8J7yLDMjoTdRvJ+4YoxZMUDwolF2LPP2xLv5sQ
e+n9t3m7CZ36nktnHj0J02WhG2En84ouxGFaCDzTgI52dFIGiqw0SFzHdW7QzQQd
4a4A58fQU22N7QEPeHBasKtbOaZq54IuOdPQJfJEhzmOHaAOSz7n1hSCQEOBDhJh
mmfXVCW8hOyYZtCsTCeukaDGhuBKMRS1s6PdBm+CmF56cNrTnvsN+mXwBlt8OlEZ
AhyckZsudHNw/qG4V81E0md2wLg9yVoyaLotqbNvFu+ccUTkEc0s8pxDvYSHasp6
6l78vE9j2CDXGpsNGyYhE9C0BOSj9HTB5fUP+6ECNo7POrWnX6NMtNU/AhiYcPFD
`protect END_PROTECTED
