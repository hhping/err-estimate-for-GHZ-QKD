`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcVRqU0u5WQfzArMvnntyNx4atf3B0+Y9jStJglEEYRous9jhrQz5rfoMcj7jDt3
qzsxEto5GEEueqwcK9CfBbzPyxMWvqz+ZGqF32xM7PcIfIY+J15+QMxSgi74Zx3v
MvxjZZe995q1+RdnxOKbERCxYbjaXQoivf8ok6ACNNd0GsoiYmWFNst5fbFpqh4l
RrNuVjSYLAn1XWGWEyibm4o7PmnrDyokH7SCoZf75Lot4L6zosdLfaW6/n63aU5Q
Oq94sEYqzOuLCsAZcwDB4vRJHUlWgw8wlrWPRpMlqKPLZeFIbsQ9jI+RqhPC9tVZ
v3Q2ptw5zfgf88vJAoG07Pwo5P5m4OX0sOfN4bG+4HCK+0wrmBwE2o0UeX1asVkN
kETofGUCF6f+mBxhrJvOfX4I2/fCx0vnPbsTcGRKKO9KBjZrUe42WbT9sRUqL+cM
J2BteCYj7FA9Wq0Jx/kOlB5oblAxqUHVfT9BEQRscnwRs4PK7IHxtRT8xcnvcNAn
bZaX8dYbyKpJnrdch9NTpg4+sMsDnToVMtnSvQ0IGC7bt1vc3kxdGPKJbox6CRAt
JD8cS6LpAZdc/e1z4GFIpOImHV4Z9KUIWzsfLqGQQLZOv3FbBLTbnK3jUTYWjFPD
n5e28t1KUenVZ4gqLHb1At5coToqiIGMSA5t1pPjPGdaDsUDpWGB6s6en9lPYyYR
gcOZvTyVGHIOtESL3c0LtRHtN4Gkr8rOH4C9tuvn7AXxJhaowBe2XUSxxprTtd9m
TE3fcKWkk/yT574ExgqIc0RTOr9WZxu7yqitgEMLMUQS0knH5GGz6k4zoowbrPfN
p0eT8opljNl1niCtKlZdENenmQ0yMHO8PJp3KIqnvV5/l4C8fPJflIIcRUrIPsrV
+4um6BzYsHZDUpQYv57nky1o2CpRCNsfeWJKk8xsqcyS9VpK5M0b3zXJyPuFTJrs
DHV5N9zXhEbbYiscD9Z2xw56DrRQMWQGZdiZkdONFM8OODcJMnwA0PpyYFLZ4azD
O+F8RT39k9Bbd9KDutp4HrZdHS7r1nz4xz/4bI9ccMUkZhBNbaF+rDT3vbae30hV
UqtpClfKSSZQDIjo1hjQGzisv8NN+4khCGr4jwRpj+dOuci+Io4HT7SQfTC2m3lq
iMEShxftGlW3NPi+byG6xXpw9vTMF19mOS7u45Y288RhPE1Oza3n6uHxcqbdkVuR
eO63GYQcBRd1YYVBaEaCnC3415fA9RQCRgJqHi7/mWjR7dm0Yhz6Dg/2oPq36rQP
UI11s3Ux8nsHCvfu+w4CAg==
`protect END_PROTECTED
