`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ikc8+F4ksGHzvPWDWD//29N6tG75lFY5axdR4zIdWwthDj7cEvB1GbcqAQ7KiXQD
BNwnQAh1Xj868rAjjgLAevIEtTn774aYW28kXf94FKGGWG/oH0SVKcwKOmI25SKk
CSBXwVsewnIFUjyEiGb4CGH6ayIixosDL0FpRnVdM6MighUvL2+CG1v1ZBzz8t1t
ocGEmYyyhNfyhqVopAcV1CY3W/+86PHhisbRP2XE61OZJIV3NNxCpoyzUvOXy3yP
Lk4j89zHLb0roqzT8nnz1h2JMPOIPGsoh4vsWI9fyte6yvXprxl1R+h6yyOnP9Kx
skWQu5bhtbxIHmXUL4mY5AWXkwd+BGLIuZAhO4xZ4XzIZ4ZpbLnq5lMpCtMoABlH
mZ8CMDLzEktN7i1Gy/CLt7zhFxeTJvLtVHt4smbPDx8=
`protect END_PROTECTED
