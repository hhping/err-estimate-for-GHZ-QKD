`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktEKc037LspGlAYFZPrekR/OCglfJhbLX7aDOJst/6A/Vo5ye8SrVnbzKumFcxQ7
JpxepI9SMVabR8xBzqj04kBFgiO1ipzY6bjiU1kNfph4Q3W6w1OKs4S0qzu93bHI
Zjr5YUrcZz8Ys8NhWxT9J7Qh550z4t8T0YZ5RBjNu7xFxaoJNUJSX6uqi2cH5CTS
lrXEAumo391OHUdLx8tvFgHEKIVhaUi2Woc5v1ZMO9lNR+zftpS8mHV09PsGdeQB
JL3Op2Ct7yyPMnd26+iG9Xu7JmJCfB26tRz5ORqipwlZUKO8k61SDDvvTkZwYV7d
Xb8d0+45MYi5YB/P69R6IzVKfFhA//4tUuQ8xn/oK263FSFKg6sDHt5HJ/qDMWIc
U2WS+vxOmjRyqG9CuBWLNIIhQFMF+7o5Cqql0dMhXy5J58RHHDNAY8UClCuPeOZ+
HGMoaAYkAtbR90b0SeHycSLz/tIzPqTvTD93K3Th46HI18ytr153ernUT5E/daqc
P8jS6thhLkYBt8bpF6Gt+jD7NfZ/m4RPnf8E17ywTA+OvC+/bZoHY//P/Gwrvk4l
5TgJ3prxvr9PRhhFssMDuHVXYSJTqgmRmtQGeC8UKIPBP3dnRyWFBUzajB/hBEz/
aMkz1XabQO1DF1P8UGp0nlmqUQalHDCdyWFFK09P5vEmsg8N9CpiwDy+AesYyWO5
Wd8pVk08sIYZdZEb0Tln5SWhMUDHSktyD6CXxfWzCOVXZR9EJjeeOkHJ5n29NlLW
KosMNcXZJuwN52LPccxeoTy7CZGG/ZkGNuHsiBTZT2gRMsViZqQCsPVH+OC31E02
Gso/aFqho4WpluVdGxjY9Z8VAcQ70m+lrKBBCKXczQRgmW+apOBisOQnBd1OowPv
lp3D5aoCn3DfsaPhYFjjPfijn7x4dQXK89COXxIHISyORj4baWdLtNBRA0UiOWOG
GnPPhhWOR2vuamA4m0eq+8sxQfbMNkDzCDaj18rBZMa/DpCmSbdLKrnhL/QMx3iD
QJTejzO/QEWLCyzl/gVCyH86WS1X3UpnKzQV4ta7vd8Qf3hHaN+EQwFzY/iRiAq1
S/qzXEYhxP8kQXGdDRULYsK0zTwbpE0sG/HsGL+TVWLgl1FZ4ztOq4HKuvMalmUt
ZgaVZhgZUpKqrNjLT/jtD0CSAttiu/8+OKSxM0rAyIdZhtVeUNZ+eEuMPBR911V7
ApGuOEnnEZcxGUqfF9/xs2lia4jIgDw67JZoKdDZBWA3FpF9GxXwiUVtV/PkvYsl
zV0YVGHDkNCt06WB602M7e/xcgXdHDT/vO9EIzdtNeYttbAFWU2FBO6Q56M+7FJs
KARVuwWnrS11qMd5vFkIJe2qJ/ySfZbvLlySperG3Cg/u+eIkSyy/jSxrNwj+2Ur
XgYy2pBDu7e2ZcAg9wHqfO3tHzXQ9sTWCZmtP96CJKz0jk0iLWr/cuK/HwlC7bI6
+lwrHWk6AREVLInZNSMejUwA5OHJTIXzWO/Pv9CMpv2nLy2iQFR1MNFIvKTs9IS9
7fOLLws4SWP398skoIJCIkSHhH8ibWQYxkTsOu1yobGHAChb0gMhkxtOjG5i+F8N
9gw9v0UdAHDExfA3haQwId56sRxBoxr8SK/H+aeQYdvzdu4vFofSEygzrIROeXM2
nCLIh+4rwRjQlupbDrdtpxjaH9snh7zUap0lPJ0xN3XxWBjf2zgqSG9DUmbjimzS
AKIqYoX5Y5Y3z9O5cMXm+qCiOOm8gFDssNzVjA9sw1GuTEgXLuyySsMjLegjZOOq
uS0WSMyoxU2OSo2Z2MP0ZE2M7mxmUh5aawm9eRUHAvyiDbm3fY8dLZFiuteTiKeo
7zpSyPkKDDn5cyG+aKsVDOqQThKtE8ZSDh8doZXJScuDzTjqoTWS/Hs3T1aiZIri
ZmdpxsrIcdycdHjlPkQInKDtuAG5qp2H1bBxkIZsuyCJPL57HoTMVWs7RQRuCY2x
accm3VwQfAz3+hEiuRIrYd+I5YnqmEAKy1JssSIvSIQyLt1gL+5WzdS/bq0iVkcO
mPDtftTjhW+HvuFoqcdRaOfo8H0Y7SCIVfi6tyxbMSLuYSZ0vA0qatD1zFA2VTFZ
QXhlFjUoQaeeyLyMoe7r2ItTcPJzgtFR9YfOanDugzeW3di2x50lp6J3B0TRQX3C
3mjkcV0S36ZsKyPDeW4/YcyrPVPqh9tXrobEUwtS8aHBQv8cocMahZQu61w2cil2
VJ9mfCRATwiVGfaFCaUlQSugk/gjjbknKrRajsAIixK4YowyUCKq5p9QSdI+n+bb
DgEzTm4uG5jViaW5pA3AmgOJoeFdComP1R7z9RJjLnh8A724orZzeuzWpH3U9MNz
MNT/MdNzp348eZYsiVTl4Up1EorHteP4rG6GAisAwZK3yqcDIXS3dxLnOB82rZnf
a4I45ON9tk3AJKScB5SujwHOttnJVWYFGAolu7rkGx4BpbXilruorI1coxM1Zpl8
GWwSVZ08xvVP54AyUaZbj5UnH8Sg7nEqFycto06JofbD40MJnhcnoVx1ns+cY0no
mKs3UAQDcYdSNbwbujFDDNNtG8MR0JOS/G/yJX2ommOYJU305JDfGcPgllFkdKcM
/6Khq1YXH+GZhgUTVsE8bcme/cO+yC/fPp7ua2CfNoMSxiviNJ3m4lUOia3Lb90h
b0a3k0Ml4CVH9Q7TOGD5agoKE/+KLBTmzbd76jETIoXnfX6Jxa7QES5cDHtFGYoq
rPfmxiiKwahbFOyBSxFH2GmLqKR/i3FbRy5D2JHebMWX04HVJG/MF0ZCO7HNYEAQ
iuvN86j9nrTUF3pSbHzrPzraF8szXrdzZZO0u9e5ABdEaLf86TCvxca9rUARXWaD
65JO6hSCMFP0xOBnt3a1EquIHXpdwFeAgknN+79kWkHDI+S1ftBxTGWj+WvCBjMy
xL/TDIUy2m4SCD3/M1xhIuIaCKO8RY1vcub0BJdjkkLEyAovQcXn4ReWGrCHFzys
LUEd+DESIb1bDk4kL9qTto3BdF7eJIgdC4u300sOH0zI8RIlOHpUpZNXLpM5CmPR
KkI+T82yy9h5L9BxU4/U7QMXj/yoKPR8rvKNFhO5r2Vij8ZBQ+CjRFBB8hZjIi2a
4lJNdXZ2QYXGPqfwA0Qzd26YzTo3Gee61VHYsw/yG34dtEOvphFZWV+5R1MzBa9q
Ma18b+Fvrxrc3NNtE535yQB+bcD76YNHjJt5yX1Q8wmhmug7luYodi/pXSZcgBxY
2DHA8Wh76Urg0FYdx9uQSnYuuD9HSr2QZ7VS3kCuXfuBkL1RFDLJw0t/+UxXc5Tw
mBD0SN94MCzNzSc45cBfl+vUCh53bkRINp7iZkX7eDB872u1BWfbtAxWCtIVDOCm
+9UVR77gEBpBgC54oZE1Ve4aoOy2NW2xBN12NO+gM9LLUkWLrboNemTbEXe+Ja49
RO9bjZDSSJTvg5FKJ6OKOs85sgoeOX24EfZ1k33+jO4KuWMbbm+BvgTNW2UIQKuD
9JCnfTcaZogNWW54Kx2y/4z4W4qL1eCvcw84bHk1PvbbMhfogxTXhUVnvOehEaNq
IkFuWbdCrWjm+VCDCkICv7pSZZAnbPBwgdKMLjV489cAlzmdrqzlm8vtT8wX2xSJ
vcw0kp3hisRsjE9TC+L3NYbOf4SVpo3tvgJN3dK5YGEATx1Ngn82FwvBCeHfSzDf
oU1ihc4RTzxQN+nW4sXtk9cwtiskXMhIhpsGfTQ+7Q5SruRWah9oX0UgIXvRJmgz
o/rRA6+NQoJls1s4kvdBUlhwjewpd7RMbZEuOJnl/YA6iMJf/8IjB0327/PtwXnf
8A7hNMP79qAixrdb9AEjeCnT/1PVAcBaChX9RtH7+SOYLxOEcM3+Cp8bUD4pYwYm
TFdbR9xN3kgjMeB/tLXmAR/69hHafNhP55h2AfkKljlQhRfwTBXO5BVu+6tIA99s
VPFe1UGtkY6BH5j71izDHp6OqB1mxzyaveVKd7Xz6xuG/b42Q5jwktm2nHmYWzbl
SWvEjNvQotirYXnsXxyuxyFXpPtO9hM65vhZujNpPon/jh2/8J9+T7v4pyPyoNrZ
ybXy89CfJ0cMsEJChagkopNZplAV+5mgDQz/j4C4ssO+i8JRc79oUk1rCbnD8g09
lls86XatHouretxbiaYKBJ8wBJqLYIAciYFLgJcJwnAEI4uHKE8Xz3eLUku661vm
Q/xKROABPh200xAkGbwTaEKLBgo84ExGiphttbNMtvBIwSngf73yVsIGo9pwfj9F
WYzBrD7i58KSSBXEtFK0SvL/yp61T+i42+IJiOicT3+sLUW3CcvZ9TYFNS1O5F8x
h8fK1sfL3t4P9Nl0Py89GQ4hcTmdeXs2YICWIkeyjlCZJd0njSkhTpGERP0GVqQK
Tv+VQXxJYcm3XYV/lvGpUDRFpcSkUEDoOQZv4X2tWapD/3pVcpUBKU4F5+qmdoHF
a7jqFcCvXbGzgxXf/J3+mTP03OvbtKBWS/5UvO3TwuHJ5C0jf7rR7kQHL0txEzC4
VQeXRwMOsJqZLazcREZl8QBQpgtTNHSr8WENYvrEXVAT9aNq4AYdQklAWRX23Acw
55edH6QIg0adj53jndyuTOpSjjwzsQpqm9mv2ck4l3USFu/8+mqxkl89m+HX5kRS
X9bghY2ilHpHlJESgBofbydLx/Yg3R5yyLICuOYcKjORfXeCf4vGipt0mDgzsU7t
IzcPBN0h9jKMY/LqXq/6a7PMv5BCt1TNVU9AdnBonsklOa5DFzPHnXpQBM3SqqvX
s8Jc9J/+z0XuCJR9bX9tg7GTt4zh3yMgtSydOaCsTmcaRpD1a4TU45IiGOKAeLNv
23xDv5eO0tH60JQ0z4BAmQ==
`protect END_PROTECTED
