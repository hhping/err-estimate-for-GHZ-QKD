`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ijQb5KtGkDjA/0H7T8xPfKjAKxxOrrPHy1h+s60ERRL/DQrmXtD5OjXA336uyrxa
SwIoNkCReTqayCnF4nKvmN9JotQtfUMSosgeQWA8NLdCfXMH3fJvy/hLlvJEAy1l
NP5IH69xKYo8Ixl1Rig7Wnq97ai1+zRtsPBozXChgiX9YyghpcmfU/IdncOPZ9Cj
lFQMwPt01hExIbn/6jE+lsRk62dUFFgCj9A1OXyOVRF/eIgpCnAi97Lg18SagM0i
5RL1aN2CNbc2stqjAt8e4vfjFYTjo32A0xcTw+SKQZyP73cT0prrRKPNGNl4zKl4
sa50YJ5UD3qcyCjUW/W/HwF2w/ySSx+98hFu77vdYlI/1iN272A/APnFzaE7FWbu
JY72IGeiSjVVObqOjCrecQ==
`protect END_PROTECTED
