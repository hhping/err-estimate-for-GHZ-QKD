`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MrLkeLZ+K22a4HfOZErLa+Sm/KZtcLYCWrFiLu9XTYKa51mLvSB/BrRCzlvADONm
oxa/0TeH2DYJjJUVluz9Zl3Zd5Bs2ygue/SGlimAFyyllJIP9Nzd7S1Lnso/IlkD
hRh6d58y7mo8N56QqOAcq8XO77NkRDdRG2qqAH2jFCzJUALGPRS8vDJasf7MJi8V
y17L04JgU52m5be7s4rmja368g9WmqhijTvQt/mwRBiJ6F4kMTpgKRZIW+kSzUJD
BvRkHq9gBrNU0xIVIlU3aZ3tmr7oSsHynz4fjmdC2kA1T/KrfkBHcqnUwKmwDkPb
v2aO0T1BSPs4/Hy6DrEJRXIUuXIObDFnnwaTAl5OzdiA/uAQ7pF7b2VZqmFbuoBV
S1PbdoPl02pABLo7PWkCFdC5fjrFdtZ+UBk0uFYvZ37TOz+cE87i9E+MiXVeewST
bPppQFgLZrVt/PKY132SyQUkqxTENGzy0FKDpWq0OXrZiQkfqOG4PG6mJ22h8kA5
BRTak+600369QaiQ+0WzLwds/h+1HVZ918kSOe5gh/5V9vAqGaeClBykCwoU81Vv
wrpyAaVWwlD4ijp0MZfiBf4reHHKWpgSyZxu3g4ZWyoOea6aqnBllObNKp8uUdYL
dHtmXRAw0o7vs9BQmj8M63IzVWYL7y/eOrBciPUSZUWe3O8o40OpZh9Wha0yicg8
vDis3AOxeuKw4nCEkOFBgK2aP6SP+7gK5XVE8yva9P4t97FYOi5qfvGuK4v8NiZF
D1cNZ9ngtSx0pDc+8EPwztdajW6Ik5N3Ndc6kpyX8w8=
`protect END_PROTECTED
