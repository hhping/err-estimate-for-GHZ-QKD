`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xo7BXyZF8iLREPqCwzloiVMiQAw9dWUCnm3QrQ035llMXUbqDJTMh3nBpVM3oI+x
1PnXMIDVGUfY0pC9muTgsT8Aw6qy7iLIFL15ZdHqLfTX0M+7L64x0VR7zh1oJEzb
B5FO5kw6QnM5Gy/yX+A5bYx+H8B/xu6PzrCYiVUqoxC0BRcx0foNw++pZeR1d2h8
zfsgamsEVar+EzODux+VnE+Q6gyL3JWg5Uw/jsIG/cYeFpSRsy9MyzBZY8kg6amr
8V9pi43hQq06jqFuCOGtgQ0qrCtNhLS9ebfgkFOD2UE2dWRcayBwOCWMylIpHFmt
QUpwcTw0CP9rKFx9nn2nzGTagDu+ZTlSGSeR0O1gad+Mz2qUaBXH+F904AufGU/0
blucwSWBLEvY+Zf/6bc9clgk6mEaA30r4AWxrgDMiLnyhJAoXn/1cjrfZT0UfcwM
LCQ+TtuqT2wxemmaHh4SNgFdxeILXECQZWPufK69HaFul8og9e/YHeR1ioj0nDXG
nA7LUjyTlfDxoYJxOjftHlQGgvKrlSInGxMz3JERZJxG5anx3dttz3rNtQphHCQo
pFAjuyPGhn2t701jlKYrgOmAgXutBdr6S3vWCFkpM9R9KOuyX4fqWqMu2wo35W65
DYEOgEz+UV5AGCF0z14ofOdPa2htiSAeF28dv8a/z3l3ko2bdzzUm18FPV1oHY1o
xzfw9woDVIdJ3H5fuV8+KRyCWdQO0vJinOS58++xPKN4ga8VqMMllqx4fYOtCt7R
0PcLxYX2oq/0Uou/GG+/00Z2r6ZwZpatLQdYsBmz/sfln4Q6SXBV/aSqphxYvE9G
R2VD2cCLPmjPng53YXF51z5wzbemKqupFXTFHLM/RPRVNeGUxZmEyQ33vVS6BSNf
nbhBBZWrvVDvZlsAQ5JGNQ==
`protect END_PROTECTED
