`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iEDdtwG9QWIFcG2e4eNqmEUMdagrw0X3W9qY046fwqnlKMe9SJJawq4ZOoVplJpQ
v4MFKf/EXsNYvee4Uh2UFCQII5qJWiLphxBW8RcGAn4RMQM5T3PJDgdlMtvAs2wD
YoIp8XEqqsSRq4SgbV/n0Yx6z1Qxjt32JiXR9llLFM4eDuxO5GE9Th7RCaBqdTGu
32k/9//75RhrxMi9/X9wq0wGyPyJSngUru8esu0kEgfVah+OsgXJh+WnGXNB8gHq
M5gEV0cLTb4GGwFT9iuPX8OsGS78RlYPdfF63T46vjtEpDnIK16POjGY5Tc5gQjT
4XTdawXGitqAUVPZfY2IpHzhKLytjsjZgCLPaptRAcT9wMlhEYH/GMJ9pVu11/2X
iA6Aak4UQk+f+KuOkf1nuxB1yqykCtyFYv7ZcIulicDRN82LWanFvDuAv3i5nfqH
egFmOSPojwy223lmqMcyAeoG91LY4lcNeGG+6Zw5XRNqB0rqZeKVwPnqSVJ9HEVU
VagORntFIFZi/Vci4MIL5q28wSAj6iKVRg8SWDjAsHnyJqXlB7SUnGlKQ82SRYdl
hHSKxqjrTXUpZIiueuUaUoWlqDu7Y9lWuqK29AkVxQEybivGYr6W8UwJzWSgcU9l
bu0rB0E1X7dPDmjBbByGCH3XITJbsJ3hnE31UcmOdfAUblzetZ/lDhBdJ/4l0xzS
x1m/5AqaS+HLz5pIk1quRmYnwQOKnqwoAcjqs5x1gsgtazRQjn+OXNVxb4mJO4UH
IxXnStPVxY3Ed3blWtxkL71du+f7po89HqO200xPf2mFbV38Xo16ujHTKmKnP6lE
3g81C+zU8rPxrxU97UvPMg8MPvXkIgwzBpUnMJ6ffXNzRbrTMrC4NEWgcF1A615m
CVd61waCxg5SIgE1WoSZ3GVB+YVDE7VpqLE4JOcxY3JgkFdHmY6meSwNyd9WckFx
eQt4M/S1CtoZriVciSDoCQQGNSnDE6fiI0P2NAGWND73cyicFyg+RGAQkhxlMFFb
LB5wTDJUgUZU8+xYxsABDqjOOeAK2mMEiYjsx9uH54xe2qfGt9WmQrghnuIglHy+
DFZKsiCft9b7nm4c4uQxCa8op10Z9y4ut5/qcrP5JsX3B6Kn/JG6WvTNLqIGtsOQ
K2IOjyVWigF0bikRlEImscv6doH5zKMe1NeOC3+0rYLR7Ao7qpxjgHQ+5uno47XA
2ccKwK5pqIcevtyJqLPNe3Tsi9lp+IU+4fsqGt6u5VA=
`protect END_PROTECTED
