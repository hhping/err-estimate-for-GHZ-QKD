`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
45rd7kzQS/9Sm6S6HWuZ8yHwS6OLkDw9N1F6LNSrnE86XPUG+YvHFWSVMbUHd7yf
lPz9wRfunDc/Tk7LfxGdxJQ7erYyEpkmRXixGGfRjRP6kQQVwbJmalAoRt2etavy
xmNoctvq0P2oOTpzLWVoWe6C1lmxoKHgJ0FBl6IAcB9ONDtKJH2/ntQfFm6OW4M/
hq22YYXKSNz1HuMu/LrMseW8+j3vAIjougq1hd2LFBnyHWHy4QUC5+PZIjWnX5Xi
8DuiV+nhns99V/gS74ZfswWBJYqEi1THnR1yjWWSFXPobwjvaTIvrV8B2DdTqlpF
tgwbJ8GNrmzcbrHhRozCFzQgg0gJkMBIyMSFF4WNB14bOa9hfrX/QsTBBebMG/AR
gNykCb5xgK6YNwyx3R/8MNf9cz+szCN5KZpXUklGPzGEsQxm2K/ZfE6wuWyB4r0B
avExWmLPereJSwYk8aymz+jbSN9rBNVipq7iH7DBiHYGRKJ9efG8b5gk+hoVnkqq
nlo4pMn51A3hMN+TbivyZSLLedzKZaWTR1yiFDwrmQ/JEBMGCkWUC63PhaPl2uhP
BmWg4mKhgwaGYME33qryuneVWC2UJpuY7c5AcC/ak6M6wFIkrsvHlwPYLzjqgGei
TY4gTmz9oSKYImtwjBWiD6z37bUvQJbO84L+5+ZkBTPaGlpAohxbyGhnlfy30fZf
B88U48zkbsMBFTiHACRiatowymeppLeGmVL0VBqr5CAoboJae6Luk657loE9Pt73
hUxsmoDOyA/aEuuZ8HA9iWKc5OEHHPTIdHdU/qOFKNcKyxGP0CobTWp5k2XhSUE8
AtGH9uFzxTNNJR1lrEIyvTXwcAPPC5mR8Jw9QUuRbLqC9NuwcnOwEC+M588cwq+p
BfE5vtSgRPypF9UpcxwHVUdLwOXCS1zI29kY2jypVlel0R0+d4UXZBRZfNy7U5lp
gNg70DQzG5JVXKW2sLXPQv7pvviuRErkVXDovNizXJfhz8svJ/EB50xEHBXV3NM1
+c4AUp9OST3TKjEgtSi15V11R5BFGE0/rci0HvZ2tl5Qywc6vpiW7Bx/jMxdCRRR
1rBDx6noICFhjj+gqGCtI2m6HJjhMZTf7SHaGoU/1bjiDZL+RRPQl0wH2tf21B0h
LYbusCHCHXAuwMSH3jZnCnz0B7GuKErOW7QNzS0et7kjwgxkA3WIf77sIZ2gWdWb
tqCnPDl/VH4GIxcvkwfkWUxKV1Vtrb7T+l8Q9lx5kSdEZJGFTE1N3UubPqvl+RAN
EFDSkZ1kuz7+/RzsAADpi3L7hCGM6uxySRo0yJhT65/vklwD+6+abQlniMCeAsX3
lrbeAqavb0tTaLgm8ghgkpAfDy3OBocDPQ9ft9XbD6DYBDRMjEu1MloXpLgN9jim
grCu1PLUgLc+XCtiHawFM6ByRbGvLsRauoPeYnz+FOtrQfV/vVhtakUAfYbKkcXd
b8j0JZshqNWiRnjVk/3Vwjzg202HLbNLRvHZ0RW0tlHCDBZx7UJ6ZEcJQWqmtvrQ
E/sopi2xJGIbXzpyelVuWKtVdkkjFAvm55KCnfSn85D2iCcd5gJMzS7S8elFKnvp
SNazMAank1za4uOaJBguSHrR8eozJhbbKr1B49ct7Vyf5DR3N105cbTAoC8vhAoa
7oVO1s+5AP3rstAUgWtEJI5+ExHHAIgoTXJPwYX8JjrUbKFsWsj2dnyoWCTk1/Ym
7yqc+v9oE3Kc7mzAMqhEChVvTXaoM7lU+izPIPL6diUIro62N+eAer7GWu7eUh1R
ZSxyR4sQ5nRyzSANgRmZQnunBYsjMg7cVArEjr0ZJun6bfvukpKMZ0ubjC6ul/GL
LqwlV3chf2AnciIPnaw37qanNXQqXvi3edn7FlFX9T5y8E+/CGVKI/sDJooyPNBS
4ZeU/cDlQ2BKcXyv0BEErsVr2AWRGo36d6EJ6RCB/wmNuP/dH6Bz3L8XlVZiSrGs
JhDgA6QEun9PnsR/EEtDD2xUpZlAFvzwjY9L8sc7BZnL38GRk62li821gBIy3BS1
HWEU7rS6xfzFX8iJlG2Mcr1/Oz7bmvEeuOGQPYDE0wMSuHYlAAurlBqMhs4YTCEF
VIaxzkWMPV2nRn3taN78jVHcRSQ+0dVgZT5NN+aUqFP5NaAqVvoKTgeUZ38BaIU9
X9PBOm1kzFFdYuRPKetd0whm5ByidkZWYjTkJc/6aiRQm/Rexn8k8X/u9pejRz1k
ER3V2+/aUnmqzruSvYV7d2WpB4M6ivZzOvEGlP39p4GsOPhnvc2CQ6bZUClujIfG
zpWY2yW/n70w/cbWolrrO2+E0CRNbWLtU8TNhZ2pqpru9ZJtbpRiMC6cb35iY4bO
cO6f6y7UtYL4QA48tovsP4pGUkoJ83WS/Gxyq/I7MzMtkb9ox29lw17puy6NzAQh
xJC0GsOvM/ZRpkuQBi5Cgf5gLdZvS0Oj7YWK5SnaB//XYyN8D/icbPKcoLbDWvyk
ex+GKhLlok2oo5mq11Z1nFYoIz/Tx7lQwfljLMlvT1IxcJpItI4bI62c3Medr1oi
rcJ8xe3PbSM9uHOLdwETtnRhxFomBE630721hIQeUUy9SyXGr2F8rC1aIK2NAIV+
XHLBd66s7QHFDy3ZcmOAj5Ik8RGj/JpeSOv8BsYl9e1FOm8tLpeV/CFra18XG6Zq
IX/uXdcAP4+rz9/92VS133KmZ2OH2lQSY2dya/BGW3FX/xR5EEoju+mzECvSa91b
p/JPTvTbqx3SF6PsEi1uPBpu3Ww/JF3G+Zsiq/atX2+0IWMiRc+zkJ5Sp9YFburd
0KLQt3jXVnG/DeJz9QtLCBDg1ixzMHXTKw8BvMwtiRG2nd9M6E/qPPBuwfClBJHo
8Gxdh5erK7733tlWoyeLYZmiO2fz85X3ZdG0QSLODScBhHUtugzVjxJeiby2K8QS
n2LYu7Vj0kspb2nl4BwCCBXXxfbRpp4IALQFpsmJRACxfjJB7TSl0AGE0I8uZsPY
WPE+pgYp78/bXBOO3RiQWpj7/+oOtU+SehmrhOmGiZ3D532tt0m8zncdRWsc+mtq
pYmdlU8cCqKfq230wb8GqWTZ/KwD/ZuyEpOvNYC9YF4qABDDrW7Kc3h/nLVAmHVd
8DriKB+P05GE+ob9ZbPL5/hyVwKZOXqYAfdGDWHdbemfIImVdGs993CsEZNtYaxz
Krsbhn3AYGNDx4TqgKtLG9kkRITwerli6wRv5b+J/U3fOn4QruOvwckhOMRIctBz
qJud404wQNS0W0Q37RqLX5kkrPWXfp/lsshISubP5mDo7cgsxIXSkzLL6uRes+Ia
BoqOAEQbKl6xyKsuE8ImxkSs/zIqK4qfOEmNngqwIK3UMlIPGJ9k1YgcIiE/rS7+
2jS6Pog9JSOOCug7GRgINPL20gTtT93qlKxvWlCw1XM34ITheAJEkMKfp/ECLLCO
l8yOcNnozrs1uTG3JQWIvL6rvjMC5WDKvKErFe7o/dECCYgsKvE6bPtH0YY8VMf4
T+0OocHOaPL/wkPodAKR2JUVwfkxgiiLlsTz2cyqlMG65z9bdXXqyhpldaTXJZMM
Z47CwUsM+84NAF8it/K4LHPGZca7hUz6n4NoULw8wnYcmVroAmPcy9+3sHBe1WkL
6pZDFfce3UaNQGbE7DK1VXh8ct6EbjPr4Yx3F/ZQZ6PAoV0+e3trXaJ6QvorJg1b
EnXSMZ7WkEpohbQD2FBtxdK1opQw+mCT/LW/iIp1XfZtrmlULgrtZ85g0vtwhTgY
SaV0nuQt0JBPgiv2k+KxunyJmNp02lW+OP98BFhYpVbfjT8i3av27D0wNGqjISy9
+oaaiqLzaG6ek+ZYwIKCAOyqY+iWFFtLb2ckj2bAHYbDZdHabukgR9CP0qdNtbp8
v4fm99XMt/oZeDtU+EtQoivrVJr4IneBub8qZnQtOfnHZyIxUeAiGx7vGUT91vWR
N4BrVfhwYvMI2DX8FCOs7fCwO8lK8z55cZ7+RO8xdY4UjI4wcruPNYHE7TX4hnPE
nTVyrAUuMwR9jSc3lXB10rmfzVwi2mKDbNoavVbfKxcVWpk78fqj5h9pROtMge+O
krxlncOmz89fdt3YCc8neA9Ya6hWezbE4y2Rrcs3xg1pE9X+YE45LLOwgy7cyB2T
rEcQ7bEs4jpwSRnkRFYPvZ27/cyuEi/mlPppZ/d2jrM1ozEArZwyFKa5avn14kKG
ofrlN7cL0X/hFSYCtEmZ7KyB1M7WKhmyR5MDd2zo+e2u3FONYMKkdf/MYLxIsV/5
Cm0df/iGf32mrK+YxAiL2yF4Dut3CjSY+fNz12u9jp6JfgvmI324IW2DQnupYJxM
K2wkTIcci3yja8wZUK3qdOXgFnXfZ9Xhi1+TXHUYda3R16tdFK4PrQeqpGoU+JAw
7m7sTEN6gEkxdeo21X4ohuplJO8s/aJPYPCcw7y61ejfR2x44k648FUAdjS3iSdD
xUeySiX6I0aHzUVM7MT0qjN5uFKCtvgqnGWNLMehAOlf8oJZQMnmDc1u5wztfLkx
CSHclQE0pjx8utfRH20KpQJdN+BbHPv3cclDfLms8DqzuBp+i+TMwK63Eb/wgzrr
nK8t5AC5gBAamVgA+A02vu45GhPiaTuDQnUVDTHTsuzyJ/396sgb4ME5FobZpF8F
5u5GMgNGkYfAjC3HhVrCraRUfVHELrRSYLJm8/DQtuJK8kmVumZXxpol+UpF0baW
yNIHkQcKZLhnTND4Qu2y/BBX6TwVZMbVQiW4wDH7HxTQoo2UqeOPS9qT42XzEnck
k5nu3X+nCRxHKtIvwbbNQO7UoWfkrz/rT5FxDFSDO/uuZ+ptmeo7+EbfuWqj7s68
ZwcEToeql8oZErfAnUSUzTbG4zqAvS6TLMHmuPwXA3EK72o+PnoKRTbqa+A/OgLb
Snc5jmoBVMdS+ZX5dh+oG9kD7tN0pnr/OKtUUjUK76gl78JS+7jaYFdLWfsJxGyC
kGDrkWG9lYjGCXlF4YHBW7Az22Gf+af1JGZ9Dj0XfPRnPD2OOCEbh1EDQ0Xi+RGN
zrMagrNSH3TGkCkoh6PkHPMT82bVo1q3MopseKdI3hSFT7ifsNqY0akTadI3g5nG
GoCWs1FfdSBd0Lniz92ChTDZBbTtrbXYhhUv0ehahlxsSj/4ISFubyqXPEvk8SRV
murOXijFtAfjCaxhM2CN3tIrIwJeKSlY8R+cQelBK+66z8X4Ulaw7rV//52vTBFM
RwM1VVTHC0mdQTSGhD+T2ZSCLbaUwP9zcu2tUxZpI4vzzTIAnzNZMdhceAl+guqP
d9dzIm5fKYQHC1YqMfW4jZGBijq28dkWhaz9TlS2K+1N2koA8xU8nB9Wu64nudUQ
UDrYUW9rbNb/3NwHK0EjSEu1lcMw6SR6NilH6PU1TomUoqbUQDu7C8bhgnLZrBU9
540/2m+7NzVvrxCVPCVCNzCZjS8LfBuKbhRHAXSyAZ+tt2+fWyLd0/UBRJtUh2Rt
Oj+mtwO8HB0EjfwUbBQ7A9Ik851QbcmrmKbM/QYtBgYe+/yLHbCXKJYJnGRm56fC
RsBpXmmvDCUhnbCvMFU/a/Mvd3UNK8SXW21OX1eUCoZNT9o6T7AzbywLLmxqc3KS
LODZuQiPBiUqKagBSm4b7V89qkqoikgFZ0BTaTpuIqR61pv5BO0WUf723ThS1yBN
Th+vDm4hFlFSU8jEuZ76VGYEnsnlJLzBY+c1elQK5IRiOCQ9I/JJxA9bIX79Fmae
46pO4HcOOISO7mpeHTkVNMQgL0ncG5UL+eDDSA/vQu4vxbqAK/CLl2bV+MW+F5Jw
jDJMkZ4y4kd8GDvxm+nPCdsBDndWx+AqBrSnngeQiO0KGRFjDcyS9mRBoEscP/LM
jYiKkQsmAaXVXxufb9+MAFYgp9cN3LGIm1fNTq8bhuFkf1YLqGpSiXoiBwHCjuNn
yg0S+xbAHwnasj5RezktvOByYq7VffD4ynzBPMA8eeDceB8MLwDoTI1ULF2xGOmg
bu1YN13fE7T3lUc+8hZSW6+tmpSH8ONCd8chlLZIzSbICIIP1rqgOmj3UCNj13mc
jYzQbbsACElnpkQkYRjVPlea6UOHvCCrSHe0QRFresVQOhsSHsFWQPIZR4+RAp4N
Xuq3Swz1V6GeUn5oT4JrvnkNkFnDpVYDV5AA92wGAZ2YFZfuTKbcOzvcjjBYFx7Q
7wthqJ4Ch+GQfcRHdr+HvT76H/H6EEWCBMNcsxD0uvU7/aeLzufXbUYeyss2Necw
0JQnEsrbtbJLY9p+GMbgfco3DpWPRBu5pYGFpGhPFA04YppDm9zxGOED/OffDvCx
tkNxyYUeWNUTXKS6A1xcHNcViiM0nMil+czStCkOQ6kJ/gZLxE/vSaXWqQ2b252y
69qwH2/XSQcWCpFEkMAAU/78vvi3mSMgfVgvFWLLZEqU8M+xR0HhQdu4Ox/oN+jz
2zvKMV1sROcf19v+x3n1T8ZNty0BqnEMusYlFMNBWcfo9BPBLSWcyef/PkgyUif8
EcAtDxXWxmNQJ6MYhscPGEav1Sb9gp+QkE4kZbTJutXY2A42ccokV3rECvYLxFhD
DLD0K459aBSXXJym9aHukuXG02GQm7pBuPSdTXRaLNGqoRPqR7lGUVO3fpU185Xf
bbTeo2gY4JtxXMybXmZu0wqPwUrSU3gv9JAgzMJISwl7PbrpZAzJ/rHFw0QWLXuD
oJJBooi7xrtTZTaacLjQKLOrhnI5H7OX8SM3h1G/9wWIqQsLdhQl190BRCC7SHL6
2YgZVwVjVtbKyKg+TAU6DL0nYVzBOVUZhlU9AeqTLSE84O4PeVjZMWhnyHFJReF1
o1aVz4j7eokSHE/483ESdTFMESuheLyWxfXcIkOWSlJdbNlxrZt+8ctvb7e/YaVY
sSiz8jNgGpW0vDtGJ8yiI/YtRhTcXTdvm8W2L3OMCY+16HZPqTcbWot4oaMRkNnI
C+1wrANm/z44J60T3iobrXdr0oc1uCaskh7WiQQfXBwXLkBoounuQ+//OOj12IhD
WYqVEX+pl2dx7cBYRKJ17KVK+R5E9QOu2j8IDo0px//yaC5iOnc/x17B1jLDFZhg
DmJFMf4UAi2U7DQmMIGa2VSMCuwlv3mj91d/aY74TKEKTxfxNppQ2uBFeHrIPP+r
7WRz05rttjWFKmYjpQFE0h7a2jcJoRD8B0PqcF/xpq0yKbzJrcOHxM7Q2pjPfADR
rrwKiMnAWIOjJvO6Ov9dy7Q25AkI0MnV1tjOYEder6Rhm0SRZW7EJ7WknqWFI8PC
N0ex2Fioy/OgcaB6NqKtpR7mrvdI7Ac0EflAFwODSu8UfsC+ntAUFqk0KO+yemgM
ocXkeacape8hIKFXPg2Fz87HaAbUQiK3syk9udfL4uDikMB+4jRu5wAB9C1pCK3G
E3tqFDm6sfsUyM0pEXWSke8umTxXY9TSg3QQdEjNrFYT7M5koe3DzHkDXkFyeeur
pctDlPa4r9fB4pQMxhZeEcV8TWFnh1jlU+wlyxIQMkqJIFoIL2/w4+zk6xYcDUqF
Sn8KBI78aSmUoYqWshf6s0n5nixKCpReAQrs/V8wiizsGfQPL2BiU0VspjUkJt8n
KKOVu/v9St8zBMFBr317ueL1Pc6nShA6qmv8y4Q96tpeVF//dGGSXF6mbMuTmTZt
5Cyk7Q0fTuaKUzM/yIuY7Knc2i7ce+3S//zTDda9piCkCaPF8qh3g1ecNovhw3dM
aNdWSN7GK9AzyCM/QtDbn79QN9OXk5HL0DFOqkQJbyVgXXTlMOlM7S8gSh96plSq
vecN0+RtDrDeGlLr1RlG9XmxWrcu2RyhL98pDOArzkwMl7XOQ+dJ2jsRvxGaqruQ
Fv7oFm9IJePnnDxzuVsNkFfO85QmfLJBYq0fx1MZ+6aid+sHJTWqjTxPXgE+2apI
8AJj9nC/g2LfZ+LsBSr/aB0Tg1oHM9EXyPVuDk5m9qFINZz+J+eNU6bjwWVIOTIc
SxCKehlP99vnag598lihT4QfEi7snSgoj1T3Fg+EStFD5Ckt/nHwa56Chhceafx0
gMXD8OZsVY9NDP2E05IBTaLhiBIhj/2A/w5ldb2Ah6eLW1F919tZDKjdj7SOISip
PQA6nkBpo4C+yV+DQHcCk73stD9eldEbT/M5BMNvQ+eddNN8t/MdmFz0gQHhZ4NL
tI1lpMzhBDIrCfuXyhiIN4au5al20ABNPK4ikpKdL18I5CzLIfwPIYmFYGVzJuR4
Ghg4vpPAjnS7zs7WLumGu23JtBk35fSjiQk6hy1AoVs0wy+emEzZv9/EblAPFDJL
BhUELG4+IMBZoHNtOdViQ7TLrmh6DORxBgRcUNXj6svvxl2uwh5Xr60beeYlCg99
mxBb7vVe3c4CD50unMYmcC98+c/6ePLnQ6q1bqAni+4sjTu9/GeNELH339gQ0HK9
AkKW0XkrBMwb3ox2egb/oWCtTkWmzwvDW2OwEwlcvVeJgK3/5LY2hDV1P2WBNG80
aqis2qO96qgris52bFMHrrk03onNpPqcq7WhgUFvqnBs3w5M6xaKD6UUHrZtGzhe
oSQU13F1rI0lq6eplZ60Kmr7TzJYybYt9AP4I94Yh276FNJYDFsllvoTLpGr17h4
SW+Iah38qIslFcLZf/P3I2PgWbATq2S1VC/cCJGLBiK2Mxb1DRvY/rC9kfEWBu8I
ZkMBlTUu+dRCg/MdjxdLlo2sP8OU6mXwdfCvYqqbxcOJMY3m7WAWxmdX4M81qCZn
zHjOavLbnzZBt30yaamadXHVz+sGk0B2v1J0T26cpfyuydYKvoDCKFJ8k2vsApuZ
Z6YsHk6A1yIT1UtR6pNfAw4MyhpuglfFtHM03ZLhevQBzZJJRnvooU67iCX3vhbi
ehtIfNH6J6a+iXWE/NNSo8JeR4YKOJlMamEYfNJ01JfOGMe+XxZ+7kdgXzFrBzxI
n2NEcT5Ms+61o6E/BxUdDPKlJkUDzmaaZptR7Q3UUuYWU374NLlwYCIbZuSj5tFb
9wiHnBnt+gNgq5SIZ8JSoyPKzEEQuRUVWLt7CuNwFqVUdYQ8h/KikF3x4u5I7D7F
FcDhqbEP87qMcDVVoTcsLgjHijEQtXcANff0qrIN54VngD0grt/Zbd16TL+Xc9D/
vmgo9KezZBtdAOStzdv4fgxBsB+65bpxblOSwdcbNjpu2pkFXa4B9GZau3t9LcvB
6FinuG1rUugWHToOGr7bLpSyBgPN5adIH6aMUdUzwgKEFxrAKnKe/7XLxCMUv9xR
ALqNSmUsfLR21xUPYYMxzT60FuUphJKDD6VyMd9fm2bnadQbjzDB5lA9mfRyQo3V
vrMUhR/Rm1NSFvgdXEjPgSdXizgudGt3QfZwTfogn2KHDDdnHiWDygGqvc5qQjaY
UiTM8KfolCxCSRbEWSosFmJdizxSiXnhzKX4ugrz2qqF2pLnIsSZjm/sRbaH543n
r3nKGmLtuaZ5wOAXyGUY1mwFdRgFNtjdZAEMLzvAHIEWBwvCK0h+9mw0cyLXbfef
odFtTWAgc7iBbeW/6thj42bcCvUZshVyn02zhbWbVA5ikjUAH6H5F7g7/Ks03goY
6IXINkdQfUqSUaFlM1drRof4cwEvPchjnsxIdW8gpL1EZ5b3BtXJoVSDlZVKTiWD
ZW9eytABrhV2JeQT92aQW7xaqkJEVtpQ1rh/xrgWGo74lM3rwiAZIF6EhOJYr6hh
54yRs3TkA5/wV0H2u4jSO6A1ta9QJBEGTqYBHoygwSHUmn1eb7BGPkcTgle9r8L3
L07ecB8vPLPHlYNZ6i1sO/grw4xFk28F9P6Nk6QSIfsLGlMh+YjTBKloMtVVuT3q
ClWg636xTomhGePhXkdwm0WM7SI4GXmOTGUnN5eTy04L6wKg1FIwk9fr+Fp2VGj9
BCo13VYNV9Kl631GWshN0O7Q5f/O9j+GZZDwIk8geASMGQA/CFb9YNcwdCsTQBCy
Cet+BpsyxrdJuh729KxB2fGOXew5Zts+aDzdSBVK9y+xGVRZQpF/6jwpdo6n2LKD
njkYc3QnGwWYG5pvmYhGf7n+/DFjlrR0ut2wPus+FdeZIjd4X7lba+5Us1O1K473
m6uy1AoR+lmsn5/ygbfbxa42e2v7pndeLB6fKfJLT2yQXMJyG499XZ/b2Gbks3oZ
VIOaL3fBJ7bvo7yEeiso1rYEJ+MKplBDnomsQyUPrk7LVMe1CbezmKabjEhtBId+
psIuWmu9AgErbo5EZdM9xVA3KcUyCLXeuGFJakkCym5+xk+TL31TX6N10K/5Oso0
M+Wk1H3XzmIJotOGlk5AW4PACgV/uFWbs26HhZwqN6SX2kJyGLbKHDcVzHg9lKZR
61IGqapn3CD2fX58H7u/kssdSzBEdNqg2jhaWxRYFdC1wId40lmKD0CzG6RAXZNg
OTP2+rB9mb1RLSc3YHj1QUT92vF07FDIjJdrQBcBm9BpcV5ITBdiq+3WVJJHUaAF
SvNYwxt5UCRZmKrp6OsF2YQBbnQsZdLENUnJEFYtRvfRYaYBPaTEGuPRtpM1DHLj
cnD48dAh66BCPHT1nYzmZMLlRt9rszs22KDIqqpt1IfQq1tl8lqraKHVM0Hm/nN0
DI1Scj8yQVzkSP3ielx0Ybho4+zQBeKffdaEXiYaJKdU38KJ45l+ha78BDAPdaNs
8fp7yFlA/aLc5VmvB9UkEKpmsZvQppN/nZo8f7hPK321UvWSynzbeTvG+UV9cJj+
eJXX/ICIqL4eFbrf9yYDR42YbxWSOOqUi4OAwqrGXrk+Od8VV2eTl/TqxLpidNlr
6huNDGpXOKFb+eH+5CXUwzWxLmTMGqyFOk+B9iQmAkJ+471QF++OGRpqU/42Di/J
ihZufCpXaz5XmPoMIxL5fZg1lwH61IEoCLYjqRjoqrfGxkgLHnSU8Ntn7CerW/ND
FRFsbJtTz8OM5n98XAxi/RJQ25lGYuFHnEmjw6GjMojZbUBJ9CxHSZVYGvnC/3l9
I3yKED4JJglEr+jPIwhlqDoSxdxkkHPRBm7AowBC7vxQYK4sHdMIkjcCo/47uymH
RbEDECk2AKOyRLv+QOm2iMcdEu2HREX8SUZZkyotwE84PWutWKdwubtASAjB8DO3
qPVnAwbFq3bUXbkmEMYuzH3MedTrIjlWx3xXcCaEUf2HfcB2XOYqanjYoYGXtRtD
xpJo4eyy2fVBXlVVTbZSr3vom5Atb8IXp1UKCIhh+IbTauQvOV+zpI48T9jb1ePi
SdQuKQzD6RGV6Kts7017/EAvI6cADRZQsin9ZSQfhLypi0jl3qw7Wwps7fOyYw5q
RDu4nvL8UnIbQsE19Z3HJpyVgKjF1kfKz5Do/28HgwrpNOh5gkQf1JpoNeYKvD3u
5bxu2GvQxIm8q+Xw0xs+HxvSdZNcM/v6NWrJUfKZKoYX8WZ/kfuAgUWl9NUGXGOd
z6ATP4i0TlKfPiMGVw7IZfEPBZA/6vlg58UAzQCOkw0WrafGPET4xlkKP2xFv0K1
e81BangiXIbvO5kO16tMmM9h/Z1j0ShPMriZtCeixdJ8vsuN0BlzaMA64sdssBt3
eN81wluUenV7/s442bqG4hVTWj1iRgAzcYC+5kC8DmStKbc+oCxeRR4NsFIy45ol
9nEKrZE0C0eeyudFpkCemGuXIR3Hd9evm80uzelL/NOjx9UkdzxwU8YrSKd45NM3
B4wuaUxBp0xAVw2CNkThyMa1yQ+iFA5ydu9WO+vRGJYFLMsDJt7jsHYm3YsIo8fO
nnOYRzoT3ImmYIJcJmUWDJMotmz5OH3SPRMNQlUaZoY1gbQW2FXDzTU7uK8/B1BK
DNrYSXUF266lLo6+ppF5iRdRFC5HDU1QnG0jSZKwbu/mA7NCOoMSRkBeOYcE1cAQ
GhgN0XzL6HstkjzmArOZM42ldz+0ew3pgqWUwuPW0TaYVgkFOkxP25DAXqiph7x1
0+cxPLgwrAEhQ4w1v3SRtJk64PnvOMTvOogpTck5c8+/kYTVSkRNcTcKuhc53Baz
P9pUAT/8KWtR+v8CSr7DnIRDzArcG6Pf/EyM90S6CKYmQ7SIDNSBKJJtB3ukd4ks
F7wKmnJfgIH5ptmQd5DuU+YKVQU1ziwnRTGNal709+nL2sOjlWNaIQOyARntpq7s
YUoDfYM4GvHo3F+MaRGTwDtJ6B8r4XkHE+aLO69hlOtCDEXD2fgsr3PHntwx7+ZG
CuviZDq5nEYVlubrEGqeGNsDh67nz43R78F3BgPEb4TglkCFtnBYIO3Gzd/s92su
0CqZjPtpIAOvwpP8oye0Fz8rY4Ycsb7Jcch0CFPbXWoTdP0WmEsp4VpzUaR7TrVt
aMQnPsSPMbNIt6MJe7IBXgVGlWlqTz1OUjpmk6/9oDBkvY1Crgy2IpaMNSw4W+FB
ZTV44DjNG1KlKEK2Vj2YkcgY55CDiODntxmIr4ahVgQdiWWxeiY67f9YjADZ+YNY
hZuY/x8p9ogl32EQwLxR3I9prXn5S1SI8yeqW7W/FqANqo6mIqUaIYLNval4Hex4
iteUiUlo1v97nIQNBU8RLMVYfNz+qowRILqw/X9YASJMt8Wxs5Qxza1PcM2Jtd4B
qaRtU8tLEJtp+cVLt4+ndiqqv0XHp4Vywd3DQeLttPjKSxh+J0ExwdmI80jGiKto
kaG5gJbiYGL1HtKs+rZvg5kpXnQU4uDc5Eq5g4HHFfAZslpvG2oDmh/wKgQ1TW9J
KVglZyS1E3fHP3SQ+V1K6zjXAF+K4GMO7F3g15s3VjIDpIbcpzpfVxyZFm8eyFYh
WUo8vIYXGR0zOQW/Ca9cppromcU9ky1qxaEX15BbtjTVF6d/XtMvEi01xFqHRtES
q6XaZRzqFkoY4WpVRcHQ5FrI+BX9k5TnBcU8enFJ8uK+vbeDf3d//yh8y9ZuE1c1
rz083nn5S64ao/YZux7wzTkU2JrCTAQqqVfFBv2pC5+acXsu7B4pBzZrDcyiM952
GVp4dWBPjgVAs2BKHkQHQG7lkmhaUw9y7fmt6d36DQaCxNxMOvx3lftgnVr4WGy0
ZfaPcX0YReq88hXEMA1idSG2xnExNr7v/YuUvA1+BV5YS1rbiirq9CmRSWXGUcSZ
oYpqNVo4cJms0Yu1CWs4LeZ8bxMS+O8pIEw9kLorH7w4XJg1BySFHtEUU9JT4GZI
bWNrqTZRcpazzxGz0nTeOhhLC7zsw/27hdhH/yz2pM4rMU/vZp37feX12btCbNh5
qsGoeZfefA5g0Bl9OWO1RYO8u6xmictrHEe4ig57t+Kl678hnrqzetRXfwg1iWWY
k3ixiIvChZyiTA+HXBLY/0aRCqTjRLjnSe+viXSRIR9Q38UAOUhnAnh+6GVO94jU
AUHkbr0l99EpnU2bDEPM1nHUtYDjQPswEL8HROW4fVYuyC9VUHnLWTvwBRQfFYfB
2tv5+WGVCZ50aY0pDDtC2RuY/lsswDHS0TdqQVQZccQ3tpNEIOvOHrvtMrdup6BO
8MTIrHBVvT5ZUWF+B/c8iY7GRYsEFIAQaIEXi6iA1kEsHEOn6vLq9aN1gTBe0rU3
Er20VL0Z+T/QIvSFHGMlq2L65XeEpfEH13nEJWeBnt3XI8rD+qcNTC7Ua89KWa2L
0ulT7CVSR2PCQRLaFOmvWEKKMF97CFaAJ7RSKYnV/91KCfcTxZ59VceyjGTF6ata
UJoOQI1HkQLFQ/VCoJBzrcuTrBNoSKIOpbBTO2WVPsCbgj8Ef3V8f73F1ghUtavv
jGVnLevlJlBI01s1mi7gQGu946yH7VE+y4WSQhOw07Qs3jfSP7Qb3G82s6a+j/nq
UGvevzERrvsBqqncO7H/MdRbwrCW0AFGhf7UW8C3nuWt6YlobPIbtPpO6v+NAShU
hAPkDXFv96rR8YnEy55A6N4h4yZhBbtO8QmSFrd1cNu0keOrOHilPgOOes6Hs7Yf
qyhJ9sXVAZvu/5lJNmLVWoEgolfe3yTc/5UVC9YemHcee7MTwGPq5/TsnODfzH2I
YFt63QWBLsK+96Qq79oIBPUDUj6+VwkX8EBaGZCqjPI1dFs+F3WFIrptNzvDiTPw
4fPqopGLwHiynOmjVoB7oXwVA+ugyraBINQp1lvbHZN5SGe2hB4aviIouP+F4LPA
WtlBAlO0CeFntzclAkSjguaWbCu8y6utJRbbOH4aZr3MW3a9dfdSqO5HVLC25sGn
lbju9hHCHqRedboNRG8/nf5IgiknXv8ro1H3bpPiEEG9rrFo/OUC+QuecxlE+TDf
6Hyq4IbFNLd/VGzdYKwWOoXeADANmths3Awa19ShsiELpqwU5f800wJHFoRvLsgH
Tw4U1nEOfgcgHVPk40lde6ksm+B3dyRzzNEq761UrOTktkNCzYFZS3J8/F/NY9dx
OLF7EbKMztAlWLmCAnX6PpLpBisIGlt6xZlhz3OgBK8i9keGNEdUbdRsFZ0vFgYI
lHDeTPQ/9e9fZiIOTwwzB1SSldZMh0QwYNDOqHbwr8xS60TuNGkMfC1L8MpZuhvX
8+ylvmojf0Y40/fVenUpivy7AXGUnBdE/FZ4U0kRC06mKLUwegbIHJcs4nlkV5YP
8sgI8pSrcZjXolHC/E999CcfHoHDAYp3QaoE0W+B4x1tnPwrZGyq62GyFj7WNGeg
Zu0fKMaFyUXcJOCNc6Yh3lssOWyZl+W+HNW8fDB40POjzP96ba1pMRR3yN/e8yPx
xLaplNvQFepXkJ1ppoZvfLvdecSBbfzrKuFaLqIGGtpIFNpdrMHN+xFny7Op3GAh
nza3n9nrM+BSUj2mIURyGy4tlOxcKqAwE3Ckj8cqChOyFAlam20Dnku9V89k4pSl
ib0SS38yE+WBZl48xuC4jsjpc/0fSSguxAWeXjEzjh6xCxTQWGLwdTk6YTCwCu11
Uc78EVyjcmqpSS0Iz6YQXXPHqYebW+GVlmma43LZXvY7NNgjzupEaDMcE+q0Wuj7
QK0D0+JbtWRy3KV1bCHBWErIcJfy3HueXjE4tppaxjfuzzyBiKR7731KAi9ccyyd
4CbshklTfMIDUdT9tBKrDI+OEZmph+dxTK2O9syYHCTiW0qGPdhtIXTi6PoD3m3p
z46+P/QZRlUb87WT3wh1aY1c3c6vW1ME9O1in8y9IV2rmcxzn7WfaJ1DWuD2iPzr
a7/9DSQN6dkbCYCyiUEekdLmukok3RL3C5Ks9yxBl3LNa2huPgvAIS7BMGbCZkRH
k6PMHlSru69BS2K9S8Hv1LHEa0fdKoPdy1Iu5k6D7SuCshnfEyWkk8gbaEPgQHYI
JsK4YRbm6q8/kPbrK9JfHn8r/+3UBNvDkXgi0PHBWRiXvSAxYFYLVryFdCDVYgmZ
8AeIj2MQoHhUUDcoGGkU3+ZYrx7ghkAmY1g23gaRUyAPBtuuVh1YsC6uAjhF2FRr
KIRkGELy97pFKQ0zL38qXeJUq/Mq9Vc41+kIZbV9Oo8hqJbdLIGJ+JracVXCBWdW
eOtHX0lYcWTc/no3hlnp9Q8lDzoA2R1J0DNBy/tygG/DvDs1UfsQFRBQVizN72Xr
QPLvDDyoYBGQ4DqD0gdsbIyT6/71X3/Y6mmte2ULTNPOGgCRtnFFkza9i5z235uE
e01Qt2EJbnR4pIRPffC0X5mCewugUx55RAzdIO8sQ1dr6g4gf5XOEgZA3mEOz7RP
WRhUjTQ7HZIFsm+nXETDKqGbyu59q+Bdk3Y/ab1cL8Po467LjGU9pbwqNwcySLop
xFROkjIZ11A+9aEvAofqmKz+MQBN//km9ikHvT0ogWxpijHIv9+7f9GbB53Vzkdd
QzFDDoJYqDqX3015Tar2siEafM2GSB3huwAI4cQXHuumZeAW/6TSigN8sHvU6mLB
8d1qyrXaimoz/A/dRKEEzj7i+V1UKC0WxRqO57xbctRinAczcIGyT9AEy6PETN3U
oaeRryTw4s5HtVzo5i/JDBPUut1b9ci6HrwG4zae8TnG0R7jai9+CsIJE+qqzl9Q
RqYA186axwiG9EGnUgodxTxc36dlLsU8HPGj27ImA0JYeCI9GX6AEG+G6YaqYb6t
JVSgvALH4zP5ceg7OmgUtE3Ujrvyos0IWvQu2BQQpnOS03PtWtXT26B/g06dxJgz
EhAhSvU6TeRplSRCv2AZpiXfHCK4sxalTVc7fdDDpsAIoNXsVzBqbmrKRqxYHIB1
mbCN/mU91QKVo1cCuorqeq48iClJko8UAHixDLp23C/gbwd0Sy1ODoIrD8axzNck
CPB3OFDS3QTUpJehuBM/WhcwjcbU50wY87dRgy7c8WjJ/lfUOmS6AoQTPb5XL4ue
tL7the7Pefwv+UNJulhyM/0bTY6E0BTiBTohr5e+Yaa0xEYVisn8zi7fIYNGshIR
EJ05dO9IFLlNbn9C0FbCwYZE3IiLGxffGRZOMBgDE7WZvFRUNV96DJzl9AWTa2pb
y2gZy1g5FQeB5B/Qf2IvyUKedjc7dZtoAySHff6l8dKihuKuoeGRtSJGzXmEag70
FUi5gQJwblA1p8SdyRcldYxs5/o5c9k3ejtfAYrO4SPsgic71Q3rnRKi0assKLA7
CCYFV+R7loQdWs03inf0I8txAYPL46vM88+UVWLY8jVbX73j9TnmtxcRqhRIJ6rR
JgOwjNCjjKErfq3ps7DZhVulXhtr4kIwnxn8keOVwaGC5l0qHbk0wRsmZhs1ZcYe
4zToXkH77NXRa/Lk27iDQ4FdGFyEo30Olh2sc/8aSE0pv0DAoOUJbmvw6pqxRTJw
TeXPmIjnfCia6MeLf6daVLUADM/tcwbULmMkbM3JjkHPh4tu6JOm1WixhJ5I7/Wx
fflj6jMtdteEcg5ok26ZxBXf4f/hicBjQ8Y07tlZXMt9HiPzAZ3OtQu3HnLW8Ywr
rkfj1DvntlAFiYjFKRyWZJBOQ4W1G4Hfc+5bTsQRV3IEf9aHBfOF6NgzLuKxV6nN
3gS3R+xICDXnYo04KJ9wnM+B+dWWINOth11pS73c4+nPG5x2/zwCYyj7/KiM+iY4
BmzpmYymbWKPmjUY0jJjn//W44RC4BEbjXnpYALBKGK+XBLxYz1m5StcSYtIweQC
fA5kMVZs8i4k3RBydLFclIwxc6sHi94cH5qq9V4QsMIFXrfkXwA4tVMtpCtVOBCo
bdr6OAcWzZ8+D447j6yuiFDF3V4OXmbg19ne/xCrhn3uAHaKqbtritemggBCxFtj
7ppaXWTX2NKG65CN9JV7OJiti44rQyKs0Xh5QLw3m75a/uHw9xs8bJC2om8HcBbn
CS+AGc64SHJ2MCbTrAtSXHj9q9Obf+c0Qzg0dz2gruFzmFSQdnYVgRVQmuSVDFVj
tQTwMR2NUDRKOF3cIhH/I1DEyh/JwvYsBeSfU6ERhMgS2rtbNgKq5qyoxhpmunlZ
AcNtP7V5uKa7cMjdJpLC+//jb+QZcJHJ/kxxgdgoCQ0FJidtImjR669OL1+EB3h5
hzRIIJIbN490M0ZEFN2NnXvfQArobTcVJoH9Pjfx2E+u3Nu3l5GqQCkI0tX1gRgZ
OAi7XVvxsHsP8trN6LYsOCv4+MlMeZxE0g4v46KP2dIWj84zhm+voYc2JPTGYx1c
h7NZGf5NypByEEkmDmE0js2oxWZmlnLISqyudgg4Ixa784NmHoJiYcr5gg12J+Dm
gk34f7iXDEzymKmCp2x/4xHeiLr0geEQ0G0/uxL7zNlQA5WE+DoH5F4+qUwwUazx
CQl/Z7ksoqZV7YdPeOsdWDi9BCYpy9GLAc0TgaVhEpwMmL9G3F1SWkVHoWhfXTBi
cD48glhxe49lJe2oUMDFRMto64qfASRyotdPFwSvxQa88ItBiCnX5p+KONOUx5eJ
LZt06kfSWf0jyYPGGktRg7w0sYzOQeaRlekWZWP8kCeOPvwVgpAim6caWsEedfC+
KlAn/5Bc8X7kGa53+AQcl4lCx5f1E0G9vyaCcL6V0A+0LhiXWW+ZUTtWZS0PJNbR
e38KQJOhZUR9z9+ho0qdtTlWZFFgSrh6RHF81TEXIK5HeBD2X0o/FB7Xt4OBsV7R
3foLEQIgmYLIrDoMQEBF59BpDOkrjjOF5e48ZOEr4rrCIa/QHPQojnuNON8jrB2A
67wzhP71Dl4nr5VejWjWzw6J/kj0ARJRQ4Y5n5C7e3VK8jjT+0G4Ng1c8VBrj/UL
rrkm8Fgu6TdgA68I0vtdG86gl68bOj0EjHWp1bHaCUxXqRlE0UkeW3pZBW15S5fh
CQAIkxVwtX9CrnxtNf9QLdKPbN7ayAETeun1s+SMGiLKVy22/KXOt4L4d7PZcrs9
eh1AIXIYSWfzXUs9G7/JRIHI9QXb+FaQVv6IT9MqWM3jxmBa7K6+8d+40a90L4IP
34yJwpjNMycYm+aAyhy4sB9CtKTM8LXDAK2+oGmYpXpxA+NQTtWvQyxd2nLtVL1u
+5f4P91xK1IKXYqQ1b6r0Tyfuxz1C9lj3wvLFP2tEdqv7KW7qA8UErYIIbnJwhAa
C03ekBLXFUlR9PTfXeAJHt/4ryaR8yyzoV0oajlTog2kMvBRfdwGYVtCei/rG5mE
sdO0q+COWn4mCBEIIrzfwOEGalgyg4JYXpZ3Q500u/7TNoQqL6ZhDzBIY7Vxuxgj
E8DwthKNuIm/YUB1ZSSfkKieECxzKw5VZgofn5J0q/D4KmSJT/egcQcfn/VQ/XBl
v+VPUs0jCDle/ETLadYyeGViqqTmQyr4UIVq1DOOk9Lypg1qZeWnUH0sSUCGFVhv
FAwBsSFY7Rh8k+br6K4/SH8oRAdm7lNEJXTUOuE208EU80G3ZpP7YZO/UJDrWfO8
k5sI44Ji0eM1+SJ+gM0c9LFW3sj2Xj2WtmdrpqQGbyffJ0HL+cVpKo0TgE2A/fRh
GS4Iuj38BD8l8ZUUZ0ot6/Mv1VszBmpo4/J3XmDonxojDeb08HqimZVcA5vzLCnZ
2lfOovb8aEKyKmtj9MpJP3duOnXnxhupCLCZjDWdEQOW2lbDFx6zlmyBWlCU7qul
l/fPH3gj0EUdB1cbpgmLJldwKTqU1B3bZxGzZd31Uu0pil49hpKKhd9G5IaGmPW3
e1WX+fQNUKIfBBAvDkVQSuAd82LByTyZpzKoE2ymifOLUYvn/h+QOIoNAWr5imf6
GkXHb2Cruq4e1bptLkIAykmomz6iyUFwivItKXueqqJMyt7apGAptn5LFevZK4wC
tg6OeZeSP5KtOVpR+ZHZHogGuoJYmzkb6nnBuSBfblyjwq9NrmSC0BUYfo5I796L
j6IQy5lKH/rvwrjLdtd0Y1XhGbJtlLX3aNr6raE3Oy06/xoL1lhreyficHIGY3Tl
X20QlNZ5h2ywDr71zpeL01xBnTVqA4AKQW8Sq/nT5TNz4fqItTv4CIa6cUn1aiT0
sQPtdUneeFbvVuqqwk2bgvLjmlTMhwrj6N6SbvCD0orBczvd4eJP6a9dWQN1wKO2
5lHUeRcGDUOGJpVpHqjxbZDqdXcffNEXYtzpAmMRwybH0/A5OUsIaPQeA7FxFUjo
SHUYbzXNUJySdseXbd4PBQRoFSQfhss/QJgMPf7PdWLIDnfvNMH+zLV1vj7Kh9hH
OGZm3XcZspMcto5SPG5xBvEyM/7VJh3MkKY0Alg42420hHhlavwwCsl+af2Hdp1L
Ly5XENqHr7WCM7XwinWEU/RzvYDrMjN7Vwxp66j1TbW23meOlxiBqMXoZkor9mIf
8B8QcnQaIdBrECVK1iXZOUy5LfdO3AqlkWoaVu774VwbpcsUKB8UoQuR7DbZl4SH
xOOeem2yp2FMVV1kWjwfwb2mSvp0q4EBit4g6+ylblIlU63YfARNILn40/ssAsyu
8OsT6F1kfM8txOPgxCaOlRU7X/3XBHe4cejF3AyLnTJHG/mQVRqFDAdV/FyiDyB4
/HxJNMJap19/sMIkvwS3BoYkyd3BRM0cmo4r+O8DEMvxA3xvC8hqvQKWna2zAnop
ScDGhiXKvA8FRHGFnDAlgrrdk5Pxs4qovrNDrS4U+1ac2P+KyLu9Zo6efb41U97I
L1kw512R0/Pjdi5VCqV+nQied4Av3dVQOashmNapOWJ//CAbSB2qWcBV0Bhn5w6x
Sg9RgZ1f/9w0gFVri22u0KM/L5aNWZwYjlm2c9Gdk60/Y8vdesM+xm1YJul6EvQy
Ajo5Fgv/cqRaksZ27F0nNivO7ATCo+q0ZaoCxSmIUFnVPX6F7nqW2XxELzrc0zox
`protect END_PROTECTED
