`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
89J1+cKf8DGUYfWn9AzJIAJrDw0VqcycIBcw3HPMATS9yTRyZ5LIh4MOGc56HgNI
QRcOaYbj6JmUr6scJjfOHteAKcCqrJNw2laMcIfdPXoGm1k4ipJ7W4SqXnK+Kc5a
Yqf3ApFpXFDxnv4/qqksfHRdt4uBc5e2CDGam3GrdW467viJrHC7NTJQWGiOPCyY
uDst5IoSEt7TOJ+xNijONLQonyJGoqhQhvaCwDLUW6vQApY2lnlPPge/zSZpA6ye
tAYH91/IQV76cCjcyqBLGxKoPk9TXjOwGLVj7l8B3ESvCDk8OKnBebu6sIZmRmsG
uqKG/LevPJN4sa0Mf8o/EoDytk7aocuTCTmh35rtVrg7K+jZngeFxn2hjNKgC3Fv
jVz5pt/TjBHcOJqbSYpmAKnRKEPBKA7b0Zf254Dx++bUQ8wQU0mIM2L9QBrmutqs
tntCWx5s5iE6MwSluWicAQiIHt5CmQn3G9Nsg94uVuzOSo+w4rqyyu65DEhkIzNA
4GHFRLdB1mxItrw7ufxlE8pvVlSb/8hFstgK5JL6YJv15hY9Q4XhRTmWu1zDraO7
5rijK4pMPg3+Q9kvCx+pyl+s7aHQvUXjqSpCRUTUagMZ5I1dvuwERsK3d71Q7xrs
31gRRXydyPnmu5gRvwOqsoU7iI//+q87/4YsU8Bh7Locqh0f8vf3IyOdajt/xKRm
JOaMdrYQkE/uZdFAP6giqmrFpo0kZ5DyTuodZNS2gPcGS01I/KrhD7W61TmSGzqj
kSwi07W2TXjMap7XnRVkdsdAVltM8qpRF7jwPEFjw/ZyA5qm/rIO17vaDf6BwPqT
j16MP9Yc3eQoVS9bqV3GzV9effx3X9hlIKwHTeBaNIL1r5LPjMkhjkj54DZtfJjN
OQlIbkc91++TFwgbPipY/sp2B55JiOKJsB3OMl6fQ7ExVljK9KgLT3szjild2N1r
UwEua3bzIaPkmrl1iJzFAyd2xH8ejcmcAD1tSCd7wHm6is0Ex6zoq9pUBh1F+14E
g9l24BMLSI1cHWQbXX5UTqhgM9HnlePDLFkNiEv9oEDhiAK40yK5AmTo3osSz9/E
5IJgbls3VOXyppdKai8Tmly3c6DtP1bp5zjo/RQ4s+WR94DhksFeoWCLWwqyqtOf
DopbcE2KNy5CgJXhdLTxxLNG7AyWI7XIbwx80dgPmsIisiieM1ZOsnAzf8lLE50X
NitMP/85LruWkFELdFuSHOGRl/yT7DO0sIISGf1YtpQZ565JMXUAUI41+b1RI9Nd
OTho9cLKemdYbml9D8hu8vUVlSP+XfrhvbQl6zVHreaqupXLQ/m/KtjRTCwnJH8D
UwbdUOhwlqvPBSisrpBpydeL7vgBRq+9GS0lZUL7mwTmsipCJIPHi2D7/qlhijZ4
9k37xPT6KNCs2gIyg48KkjlOGdsnyVOlIruUoJ09L/Nmez+GGU/MlDIdZ8yN1ttP
HCHzagCW5eb4QEReRLZa2HWmtqqtMNeIWd8Tkmq9gZKvqttiFJtPp+kSzWjevwqk
oFl1nVv6l+Vyo8JLurtTx7xLkLnAMpl7ybXKovUkcMreHsbATT8+7ryVHmbVPgZ5
rm0ugwxxzLA7S8EwP0R3UNx+dUE8a1dHZUFyKOjvXZ3FDu/VmVN1UgLRCg1bDm8E
XzvxGKkX9JswSUCfxP0NGb1WgnmnywzAtHNndJdHxV/t3xh6ciK8Ps8BPZPXe2Fv
5yc+eS1n51JkX8V754xbK9ePGDlDqjlOTeEu7Q/H+Dav1sErM2PtL9lgzLcLUCmI
8ujPnRRkPvn0SsRoYpiz6qrF2hCiBwxGsgMQCsy6pSi7valxPC4JyObnP1WqVouU
9DfOY+zTovoEMomaRZR8Ubs9lS3sDSxEiznclJEqUCnM35SS05U+x27uYy81bflG
Bzu5LgyOgXgWKiMlrY4VBOFz70W9CGw13m5phXOOG4rRpInKyHPVAfUSjFjhSbmf
dJJSw0MUM5bmgsL/F0gx9FBjrwX+lgJPkClahmmx5aviNg45dym4/nQ+UNYfWLzB
UMcQn317LYNXNGkIinAJaqC3Ue7amLPaVQBCpWYegWloKuW2x3sZ2Dz2g9SmHihr
ExKiwnWSmwX6Ly19qEx0mpzG06vvRybLuCs7dF6hN5DkQkUBJFVTWYQhwtZUvXio
1SPru7JZ4R3G+y0qqui+XW5PbNIKFOy+f3A36iGKEawAG5Lf7ki3VRQg/7K4qR7W
ECbFr+a5Nj/Xa0OYrWAkcedC1ILFddaPyUFNaWU1wUJpH7DMeYhTTnOEEXzlSwkU
2Y14pI77ahUXy/uFlpeOUBOiPwbAPNAIo2+1XNYsliMWKqW3+IZUoDxkw7ouSX6M
7yRDx2qpy0Mbma+z5yGTSewquf5zYvR9qdl74q++9E3SPWijODiEMFudcHpJMzXR
eSZ0tmwy4MfuUIhKy+leDEpsFpjhW0jdDtp1FUduFWLvl9dKh9yRgV1rbkGYIVqZ
gVrIzygja8San491xkXN5grKAUENEsgT3GOY3ddDRblgO9s7mAqf4QXXBgmo19QT
LCkcOPvGtounIFTYsR+pXRGreazkTlJxkIHRWkWPTJ6YrXLEKPDgdgSzaBcXP2zi
LU4uLOwwMDR26aOBGr2vVkZ9SvA9A2HNryTKplxj3W4XbgCZdNHxO9cDIYk7wI59
/FRGjW8sjUA12cE3U2mURfGTJ4q2G41O6fVk00K2I6JzU8J3LSplhyQ5j+bKiV3z
HpZvcLfTd9OPN1NnKh9TvN/eWJbZgjbZs5K0JYfn3pXr34VzbOFldhV32B7KEP6R
DkL1IjAJ2RIilYusHtZquAV9O+PD+d7XcMG8DqeaA1Az6geqWCLFZVBP9Yarn/jP
6A8sFiit3J277R8WJjkXMn2TBfCifP6syH8A3Yo00wr4NEEysNxSWwPU+gzV+NBK
m8Zo4YTTP7lKbqYEBwJV1ENNqEd77HS+cDOH+POy/ADpH9q/xCEawtNdUBF7AbpY
PFcxk9rk78jJjPdmuHZhZyfUtXZ3WDF4HoLQ6UkJH5ak1+r/GSTC7uXro8x91Q+M
2t4DLltODeogrhpyxeZk1PTSxsVMYRCQ6oklWc7QarM51CZtoE1hw3DpuqMdjQJG
bRYvImYn1+zYT0DDH5++EEd+ogJbg5LIR+hylkhFcMWIwiqZgy3nYKMdHe8fRzN4
EI9PqG1RALVaqOqIRera1r7qq4kteVraM0Mk9jUcb9S8EAEUtzs5B6Ak1lsCl63i
nSx1Bm4TY+0MZYL/QUUFZ767wS8pJOSy9zYAQhRFIPB7mTwZFps4BckKfVmhipol
wIvVhKyiBUX09f+Lj9Niwbh7jvDkRYS8LQbDGC+j4eTGkFFjZ4JsqjLpIw6F9HpL
OonYlqL2L2HVOaFUUhta2PSPnf2VGTNBSrg5Tw2vROtbP/6MUZ5JTM98kJ5ZZJ8a
BdEO1HW5hrCOHh8C2BkraCIArxzfwKpzbpJJdFVNo/axaBbil95grqUBK4S4Nw3F
/jNsQKQ2rJ+vlgDj0Wn4ZIyEkGa5kj5pKJelUk27mALFANuD+M3Nu3roppstel2d
A8/TQkAJ9Ilb2XP8DOfIBYHiVxMHPBMPcT9YRI07zvQeqf4/R6bsfFetqX3tqn5D
dLUEFHfCVW+s6afmmwC7VXcQb1vkPeMBCz80rhWbeeWjmV3mUeaP+hR9fXilzS91
TNJHQsKkPofUoolI2lrc3MWODNX/NYDe0auhzGM6c4xYXaCZQ5/ojjChwvdovLi4
IXfrCJjN119+L7nNqxW8fgJt+rJhtSS1fboK/z1dwSpCLy1MpMSo8g07yo6wIz5Z
L5pW5sC3n5ArGZJ8TDFnhvcpXuYMbBwMU5khfMwbZRYvUrdYcJOJDTYA7c3hBThk
vpwlRszz8ki5vhVpCs+ecVyesTVcJ3/q9KpUieyrL/Vw00qaoFiEyjkDUE0Z1APO
pg+Uc7hg3eToYMU430fvSUv+sfSWi5TjH2Y9qoCF616X70+vNFw6dmlbm3j4u9w3
Q8i+tYzpSa5KMyJkV+nkpGO7kU5MJ7IW87nPXJp9TgesPaFiNMl6nltG3D/DN++Q
qd1xWFJIHLwPsczu0lxt1XwLFM0I41o0Mg92hoNtUBrQZF7e/EvdIVCqlSy04eE6
01ipTM2kfICaw3cG/ZQvf4WAz79yL1+bWWjc4k8uNv+DEk5Q1i098cDx1NFTtFC3
Evi0wocDc4nIS2hRD8pVXyZ/BLmWcDydnOvWfHz2GI+B12Wf77iUEptPeAGy+g+X
51AzeQvZQ6OUAoAbXFgi+zEb3X/p8noOfj8iDrYVdW7ApUDQTdJrv92i8MIvafBf
NjXeoFdedIcqkTHCotyFUBF5ZC9XVoXAnhLMrBs+cSkEPpaYEeCzEtLHQ7rLsGDd
zmd6FZyJ5Cd2Awcjj+cSrX63qowhN2DzJRCDs5umtEXG/zxkMtBv1k4VjPY4e3KE
A0biGP8aIAw8yjqzZf5THDjgJX8qmvwIQlJGV2nohTMYjCmKSwtk1Xgi8Zz46R+Q
gfEJq9Vd0AIkSsGbo+a+8WqbEiCr9Zh4cfotyCAkcejz64LY8uBkgSwdv34Y5Y7J
j8Kdib5T5U5Ic/6/4/H1WcJaM7fDb7rxJcvgILQFvRcpH5nM6CCUHaLWITtLCSVR
SbHsMBTTYqRkmTnv5S9/9yyG+dvPwWGYgMAi52byTTt1Y1kARwzOdd1A/O/mDEwm
NMWL7UGRuRtUVJmqh0gSN+RQGNip1q+1yu9xaivWPVXxBj0C8y/bsE+f3EmzLLeE
ZJtuzodQvsvG2pWSd74H/Sow/pHDawfk5OidkKOrkcCaYSo/6yz8imrIRtgOntUO
rufUGvbJDSYBvRkwnpiyhfqm46viel+GvG/gx4A1RbxCFZgXJaQrCK8wasNBmTKT
WkY2+QxSM8dO0fBn576T4ZiMIwlNBIbHkykHB6JamHi/8ud1SAR127k9TVeme3Lu
eA7PZDJfEnVL3EcNg2dG2Rzvr+epXa/lO4z365HGDVjarIIrVfqW5Tm+uSkI16pn
TTKi8+yRnNBFKyyU02nKbHBUIx843jLE29nVheR5dcZZLLPtu+yDtA3opraGQQv9
umcpJNkwA1RnbqD9A+C8OoVTQTdrXzn1JooDgESCDpyhBGNtoaPavtSen+VKd2RJ
HrqI3QSN+ThqWFjBbvTPw+4BCZQFauxcU0+20r5hipogWqB68SXPotig2GsITEzM
llfwFHRPBS068gwDlfhBt/bIkZZwql+Z5WkGsI28NAKy/SbqEuSOL9Pv3Bd1Fy6f
Tq8/vtbBfJVChXhhv3y71VxOApFoownCoOlmULpMDp71hvJ5/jdTd1NYzRrzHals
o1SB2YytaDqaV+DjtbVNIqXBXcqQo0DxJVBs0Xm8Nvw2kPrcpASSX94q9Ltj+/js
AK0oFEIAYxbuOVTOC/IHjrWsDKT5zaisbA62gyuONZel9Gl5CdMdA1AQQ8P+ysLh
z8fYpfAx28ziLxBD8WWZz0sqJ/yb6Yc86RQKChbDQ6v51pSjs+SlRXahRA110uT1
b5cTgJi7nIjcw+bhEjj3Aix1V5sRob1nmTh8u60E/Of7n8QlPBhOskszsubutYxR
agv7Z5NtQH2GzSL9nRv6NtcxsNqWMTrZr1t+zH1HGKZhWyEYyoU9zAq+TV/QEg6v
eeJ1rHh0yRNy8D5MJqGAeLTQy+LsRIiF5nVt1MKxu+x3LXojxoTLjQiiVTr0NKTK
SEzlz6/n4bljVqbOEx4/MWrYyhXM1ifDCtK+2GzmLO3CKsGNLSv1q3oMhEx4VvyW
knM5zfmTXlj9EveBzxBo+goMO98s1elg8KRlky9woqwgGgvTtDoFfPfXnBrDEJtY
xJUJOzHzCSHIvJ7xMs5038PZ0ZIevYlpGs4mWt/18pRvXAtk5es1IBmLdZkopLa/
FusTtKS0RFibAPtNErmZdnxcpnq7abJZExloChfuKnV8EI48jrw6eAN50SJpiJT0
5o2JobGy+IybiQX/O7FdSAyVzAUlYBtQqBMIB/ovpLr3kL43Y2rI0LOGRMm/nxwG
pmNV8zkHyCSOLXbdPD8d5a5Y4LjBnWPtfU7POGhALseFzUjMOlCzwBsj5WmaUV6w
lpMqQ6UKuS/+lDg+YN3iDvz4DUf1WOO5BqQamhR3gNos7CVDCVuCqpncOYyfFJ2L
ZGjJwCo4VEsKVz9wZ2CfOIKQ4eAhjLVuGgn1pB/hOP2NdKekrrN+g29EHhDlRwcg
hBpdxWWzX4TEet0LKHXVRklTmHSNStPOKFmO/CY2CrSaxcFgn7QH/e7nTuGeUfBo
rYz/NBUX4R4tK4poo+LVsHs4sCMtM3ii5ekGNjMMzF5RsYlFRtInrHj4mA8ylvKb
xsLEPVNIIEZ/ZqSakhVRG1wU4JxjmBFM6H+4ylT7107fWx6hxDX6X6bgPopJ24tg
ubKn66p6E8vdZ7R08RNl8C62vLBkner2cJtKs6cio1LtMTVNaHMlFRmO3XIEwBt/
4FmY03KVtB1jb1wvi1vC80T9sGQd5hfV6vFTY21Re+0QkTlRcDmm9vUiXKJ5dMwi
9IC9I2k4YLAdpCTfzL+IoaUUN8+24whcJAGPpYdeTBlFpXCavti1oOEHtPPMlRep
V3260tvhZ9+HgJBriUXK3EgafsLq78Y8FZdLR//WwcAmN6XnERGrvvIuxoITrxjE
10nG5TNWGUbqatcEeLT1D2AZU0eygSziwNJzLwWeXL9pRP4t+5/qqzbFBnSqrfUe
jPBNQpk6/ImjuMjyhTwfADhCv01DJX56hiSgeQNOckvLQ0yLVAioTn/BQ/7SOUhM
0aMkAa0aKBLOs77yygbryexOc3Y8yl7YFi/u5HZpcM6s44D433NelHZ5vWmWzLXr
LNa9bhncP0RW6sXiuSTu2/x/284qDqR31ObzJos//sZbivDozH3iwmOuyhUmSxpI
zRd/cJ1o6gPMdAEdQGhVP87rUjWhclAi2H0vYi9dkm4qSG5nZlEgp8F7+ibRSZ4D
jcernEf64tu5CbrsXrD5mObPAtrClC38L+KKAd6KonUTf7swbSek2SYspkCX5JpF
dJSVNyiVAXwfFgVKwV4ONtYbbC5VNpuoFS030XdX7cuRuMpW/6w+SZz80bR69dtp
crED9YIaYglwDPyvHwGmLDCc67WmMcDpThnaj2txjYsJh3NN1YnjH6Gh9BjxMf6f
0Y5HQ49xIVd9seEOEnWdkE0MopXSrqJg2/HkxBt1g+v/08tcFiLUA4GyFrGWjf06
xBXKgv/o5qJz/MCDyMWNbf9eunuAvrP/CjUguxJPPX6TZX5IKVCix5J/2pcFQlm7
ArA3hPWVlwngwFNt8vlZoc9QVhNwhDpoYBGXlLNBePVaEdurAM7fGOGcotEkGB6r
swCWPu7mtgkgOMkrmCZzaIKmcwfftPS1QFpmWvKFSJNnwjVFnGizN0fZSsk7VYfB
8mU02gPpYJSosK9Use1f6iHxHqHJ9ZISsS5+X+RsnWR5lTxK74z5/ZDLrGimJ7W3
6qsz+VQNNoH/4uvUzczYMomn65xfbJ3H/7O7KCM791p8CbTv+ktZkALZPC8LSJRK
xVHRWkQEzvZcKt1dXnYRyhFm3nERs1AfntOXCAP1sH5yaD0GhGb2D/t9JbDQikKA
HNudHRQcMvxhmV7bCXkftKEuk67VzP7G3oxJLt5mVfc6a5+KVoV+sqMq00SlsU1P
ME6Rvq7gDjsnbaFN8uyf0kcDUFuKO9XZlV5Pl1qRU8mrGZy2SJrJvydTd1PcXI/H
sMLET0Y3CosryvVVtsnhVUkCmmpZ6hUfUQiJpq3jbQg9xlqTDbXKjRQxJ4c3QMso
B72iYcveKHDXMskfLdoyJANcTOCu3Bl/5Fl0VN0sGtcXRSyPPb7ONvJ995y4g+/V
nep+85MeCqCv162prNgTGspUAUrMtxye6oyyYsXWC0ZPfZGHr9TK0tXz7GEmYekg
BM6i0vsVwjBt1MXHMC0HHTDUJ4o2cUEbJp6KZ5WO4SttB8sZnxkErCcv31/CjcBR
JjnGM6zlgVLL4wCAHH3+FoEJklY0APp3n/pDQ4+o6o6uhMu32Y9+6CEHy+zgwCLH
uO986zdb9VIgsPdzs0CeTfXIz1aOZ3XuoW1+pJZX7wBCYrxWQyX8VarnLM3jFmE7
peRPRzi9vrS44RTjiH9rqom1jINSXJp8GkzwM4JHWb5hFixI26Asc1vQTideh5Mv
FqEKVXbY3Vmr3Z7n+/JYbL4EchXFnXYXRZSYITPb0dpyGqXj1ddcEnHx7q++DO9T
szne2QviQMK+u1g7ayT2PgGh62KDHMS05qP8DeRYH/NPxso+V3lRrDFMcL2BPnES
p8BcBfXKKgGmWgbtxRgcPIywwpQEPN3ThBowGHXbForXp23Vv2QmLR8dzS3InZtM
Aiu7o/OBSkqQ3PStJYWj62DT1GwdeaqVS0U4o10ctM76efmVy0ETgaHGCxRjtkJ4
OTtBIeXFYxFn4T395tk3tbe/U05neN7Avd5PyBDyvfU/WXc/DFANtwfxLGRDnuqh
Ar8Hc1LSeOMMVpdQ39XxTAxbINZeLIz8Z1S3Rt6DQIhuD08QluBgjDT3cF4YN3EV
MdwgZebtsBxFVIaZE6VbTtchBsZrp8aQzzYcQbnZB66DXhuR+Sv7LVMMamxXF53s
/SEN1kQzzRzQFS+DWhPbA6y5N/yOXHRuD0UQfPK2LLJFXYvD3gUr2eLi5dqW8stg
WBSQNDHl2pWy31a64VnrsyJl8QGilDES7hxthXx2mRiJ2CXjqFewtmMvsOGdZhBb
ZoMs92wwMvnFOR0Tj3gaUfywropXXZq908gN+FPrEV1aBkJUvPH86HcQJJ9NDTjP
6WbqtNbOnYyaVHefaMHMayLtW8kG+w15te+3cDeGrDMEDiRQ0J681h7beYjkOuGq
Ni5dhiECaj9rHNyP26poRQrDE2ONmYFje0X9G1QbPK/uqEsV/ClGzVZnpXRHFtSt
0/QKYzZBV367DkUHAmTBsIKWLPNptM2e5b/89g36HMGILAHvJQsuad28rTxjl+7l
+9I7a6EYQJ14+pmsAQ+ZkIKzsRnoYT3vswhXNKY69JDgANgttBO0zuGDjVyGInl/
xkZuxI8A1zGtWr0EIkhCMJt1kkCrhsPoYqT52QODoO2juCiAu77TGnkVWh94N1LZ
ZD/vmAfZ4jxhxMJohfpbtXBDEs0TDSi7ifwxOth5W5E4109JCLwLVCWxzEMYiQf6
Uk0jizdJyqYcsuuz/j7kTbqUO7FItPtwsuLmO+WX0lu5pGyCEEOGQSwV/97xdcah
v+y6RSZJ0odrIb+tq0KpNoI665+nbtymPHS6SZyyitKUC1Mssp2JASFn4Ws2yyd/
qxKiW2uNA1UoZDHoGFmLKSMokNHF9sHmUXaRDPd+iZILWQ2c5W1v+WW8k4uVHgRE
6RKU/Lg/1lKsfwwLx/0yEq4CY9iXgwCt5AOlA7vk/PqP6Gv48S5M7OwyURNhbEZX
UHJOyTpby+WT3vq24y5/lMqWxS0PiWgLUPHvj1zeB8/fqq8M1uIC+eQjxIwvsbqL
KL1A5jtYOwEONab4APizC11sVgPkCXxpFQfoXZ7M14YiMv9Yu4vCXKq1ApEp8UHj
Sx9DLIsp2HFOmjsG7xxg+yGL+vN8gdLwHrKJPfsI0OCz8g2eOAmc85mKdoNsO3XJ
dfxmmQW957gtsjiWvr3s5RwhVcJIjzhFux9eOrw/4tatBsHenuthCoPjNOdAxcwe
5tbYAIrQ3SyQk6WoARzrWc2CKXF8khVLnT6dtEht+PGx3zLC7PLZY6a/2j9vRhzJ
BbdB4XhEMpMVyB6nwqKPhexIDOpBESCF5dez3aWJiOb5khI5GDHuHBUz5EqQFo+x
9n09Z5/DYvh/MEklxXEnbypJWyGhIyKE2BJxom2+hjBTo6Zz5XxqYaYmuVWilAc0
lQCcGj89kdq7mWm32MtKAqmpaTsbUxwzuL3EQThRqPW7HrSMMIZa50YYMSTX52iu
/D1LeMWS/z4/tAhFyPyR91aQrzHMLwbZTIt/u3ewykT+hK6wMM1YpC99k5XDxVXq
xFVfgIiPTURfUghCLrtzAm4yeWnMCDMhMF5PrjCddGNgSwUKmUsp4baTr86+F7uk
Qxuey7uSWMRB1c85BDgHX/NzVVHDDys9e7yfGMXulBzzXAf5Trg7Gp4L2/PZcpyE
kMXNVUsZ5zxTMC62lf/G+htQRmIgMwDQ8RrEDJHWBwZxIqnLu/0BtjOezUSlYJJW
AC92PQMZJO4L3wNufCZOO5bQ2HzsHCuH2/yO72MpXywWzU083YNycFPxX1IOQso9
RhOCYEWU8SP9ddekjHkq0oJxWR0JAJGas7GrzHMaNtlkxbX+fQ1EtYSKouacBZmG
3Ub18iw1DBnkQzUqPJwuEAiddrwcu3Bj1n8gIHKckj36wcDJESBgsISdVO/vt1PD
x8itUXwGPuMa12rb4lICz7QM/meWzruLzytBCD8BuXSyALoATUFx6md35hAOgH8l
dG6yA5O29oZDtXVkjKE7AQ==
`protect END_PROTECTED
