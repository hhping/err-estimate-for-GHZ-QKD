`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3oevlUzUcf68Isx/1K3hH9X2YWfznco8ksFMNzC0l7YnMx56pvs9QFncp0OWaYGL
QhwaHuUzlGOF3nPbQOuFJRO4TXfu7wxQC8THU1iflmJhv7qbRrvNQ8+O0et5YMI5
DG5++MNqda5TN0os0Wd/fMxxwjhuG0ivvgA/NAWag+m3piE+WKSrZYDka868jTEk
WjO+dJHGXYN/7Q+s7oEPinuWsB4sMs8f65p85blwsfHkgqUeiO21/lR9ci1+vlDJ
x1LG8XgQghXxrgYFa/+joJzXKbYCv3ZMHLfLGP1kb7hAbdIzLHnZnBnn5Qg3nyqa
+g0Yw/Qw99GuzkdNOrtLMv7IRnfeXCHYUf5dXmwlq+FTeCjOn1gHS7Ix62YyeddO
HGgdDtYxTGR3y2rpYZLfAvhzZ37WSgAqdsY0FNISXFYTieo9fQaX9bPWXp0yjQDD
JtBkmIw/5TzY7CLu2knI8b5UCNRpdSz1vYUbF006F0o=
`protect END_PROTECTED
