`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyINGaaAcj5rbUZP5I73gaEjclHQgxD+cf7DBcVIP1VV3y/GVdTPa2u1X1e5EDUN
PxnRifhZ32vLULcfU2yvDGALsGjwl9ckI5/VO+b5a5ZLZnIkWtubHTvQiuRUCQRN
Ce5q0SSTBJPOz9Mskj/RYoIpuiRMgHRycL0ctlQWotjYedaFFS4p/7KPfhMsjTtm
N6IVa40BR0Ci5OEJ5Yo2CjcdPIrelSVsn21955XY3XfEvV0LwUUDs5keJuXjVP81
0evU3Z0Qt0UROo8ryVi9PeKOgOPEKAQufp+JOUQHS2/Smt2zNDPRwLivDIQoD2ac
EVGAIdxdz10UbeOjNqINdC+aHPg+7V4cRY/svumB4eotAL1Rf52f9cVQesCuFf5N
chCDCFz260NjHJhxTMmDgJbb65qhN/BvFzmuFE/bWksFaFYpLGpnGCflbDf9yEMv
X0o6GE79H4/K24ldt5rvMabictrGGf0XCqYX0GzMJFPjE9EQ1vb06cRiRYzfT6cd
FWItJwP2eIvhCGH9Il3tdV9z0Xvjv1JX2CBVGNk6N7i06zm2xl41ZhCT8ICwmRbs
LeoH5i8PitP5X6RrbzT4HatoldHXj5Q5T0/M+xMCg8TcyTgtL5HHPgwdjei6kGtN
v4LOwCRX1O5ojshVcacbv/+DYP4J4ck6hkA6xvsVrfv0T+8rxmA1+kMMBK/Irm9o
dAxzRm5+vWCS4liCY6AE7r6FldcIPMrllTAsGaDDpjfF40tvqbu9Asp99q40Q8x6
wAes7xC6eIbhrCTkb4ZFGWhhq1YHACF770uQ+m+EFbyRAoUDRbGHNEG6kDp/mel7
rrFAoPjpsg9arPsPe/vpDDaNYNprLcBgFwdBgfHMusRuw7H3XMoyYI3/soekfUmz
gBN41Y9ZJrO1qPwizkBA8Ci8r1X5wF6I9JoVslKibub3d3YZkiAFjkDdkDdC8WP5
ZYezEDweP2fHX6c0fhRdlJvZ7vhQpt58DJyanPSYa/Y=
`protect END_PROTECTED
