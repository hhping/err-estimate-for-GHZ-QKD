`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhaE6r4lWbKoue5jwgxJ68HY9cGRcJSftpWU6Pvtye1HAZQc1YRQ8AUyF/VE5KrK
FCgcwHCJH2iFo/E4ve0dOxw52q6ufgt42RLqQIDtjS571boUrSNhRUG8rt0JCbXZ
UiSu6nsDno+NPVwvhdjBmULrv5jZX1ITCttgEOvPoZhWrVGIOEG1J78gALt+Iyb5
4+EM6Lyr4idxBS5ZOxEZqXWTKROZaYCCAqUfrVd+3SlvNZGKGP4EPtzbl0uKn6su
oSUtTB9VmJIANiTLoOEQYju8VXYIG38BWZZyEqgf/+b7JO/Clv5dIQUSY/gZD9NG
M3C06S530w9aYkouJ4Cli4pj8HoGE8PxzE7tLH1P/OfogF27htvE8nuPDmSprpg7
D5LqBedDVxTfWG/fczWe1PlKmZQ5eBKaas99XMZznZQd2rHht5Epm4JkY8rd1WIK
tuZWrLN+wfziiqCx1kWrdiB6Mm3OKmuZ7JA+dyS0Q9FaTeE9TOIXMioP6t004RlI
IImf/pNmpRE5gQZ89WDuWTGhCdfNSHo7v+ZfAaJFjYJCH+nStY/Tkpcm60X94y6M
cAe44yxBR5nV4HBzq4SVzW0SSQ6ryxWG06GB8ebyvlaNO2HHN8hvz3xMPTyJSKF9
71VkCcxDGdhVWSnYPew0aYimf/x/vd2X4ZdGmv37b4fng3R5f3YCkarmxLEObGR+
DB06Z091GV5O5T9p//EQE/kG7Am0ObwjWUxZle/HiywO6PBaj+AtDeSLAnzZAM2i
umBZz1BQAsALYBn30Nvx9ZUw+pxfr6VPg1bufyJsijuFnKzJsRCU9RgsEWgB5f42
/AEybGE3Dw0lKi+9UoTUJA==
`protect END_PROTECTED
