`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNq/VtbsS+uvMmxnqOf7XJRiKGjDR6HM/Ya1qV2bf/+fXbHsx41oPLI49K0gKDKg
1u9l8NPmPu85DwNPk0TcBFJO5ZKRFvjaixyuL5I3l181j26FPXmvfgDYOOvZVTyw
BZNxatxymVQv1fCMXXPNpHRa7m3oFQPzUaVRl32aThOjL3wxIkgf0OvKnwr79gMv
MsvJqHeKIp9jSXMpcyFPVwGZ2GdMCu4gm1rF7QEAebZJFVd/FALlW2KFUGXMcQJm
ktfrLrgDZHg57bRFfjHUPmn9SO3n/9oWsQlTIvh+9vKWomyo42BX65/YBZ/qRdX2
1s7q3JTxbzhadBdEtsfHUTnTR1fZFb1nfnrhCC9B3emGz9keJRqVcvKg+WjkFWTr
33i6JSX90t3PEG80vhvcg39t6yR6MFOStlVVG7ejtCSruisuqK6TonS+ifuytWGh
MA6sDQiAMwobF6rL4dmEA6IZoE72d6Bgd9n7gaN4jsY=
`protect END_PROTECTED
