`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ln5L3QeXcRuscs8XufhxWctJxSEGRxD1REUcP5Wp2EyK4g6rmP3IirWb+MFqwaR7
sCgxIpB2iq+M59X+AlVlQ8jr6cMnaNWmwZL/J427GOfMHcz/EuHCNizgl/2WpQCC
W5PKEuBV8JWPnBdemDwkkDHFRGpFgWs0kFbCs7E9opbvobM95MGw7jBvQhVehztD
vpb4XEaGFtwDTlqnFL8ZzqBqqLI/eFSA86lqj2l1GpMyUIFzwxokDrdheBYN3+aQ
LO8VFtfUcYNDx79nfJ90NCyq1DChDPHb11GMSFw+WS0zajF4PgnBlwTtD16uDpaA
OJZ8iblJFwgHhPAywaq/FH+A7jnVmdW2Gv69vuT4lMUiirAcq4I60IsXbVb91QCN
LZmo9mgFLeQIraZnSYFsRF2IodK7eYWoJ295UukN7RFtcK/odLQG1QQx3uHi2n+M
qTU5/wtj7M87NkGnJwG1ALw65ly+BKGfUmVFeyPga2iQBo3yG3M6l7xzJKrg6/z2
e7hp0pam6y6L5UZcpXcyAgin2xPaCU5vHX5paUPRbq0IIPEnTnSskWZ/XJuqMNMk
/Mt8MBjHmpB8FEL5Lr91aDvS9tBqyRqHwXOlX2WmLPf4scxFxKa4Uv524MUbqRyc
sKuB5DCbP2s7a0SjgG3m6jimzGyWqSjpqT4h924f90d+GsrWUNBGLLCA1TsCwHpJ
tsOIIjCgg2fWcPWpmh56i/srGXJy1etNdc9cS/fCMrynfubcXnXO2SSNAASHn3WW
mCrPofzKnhrtPLwU9H5fXrbzOpKlsvOO8XkYyhDa8yVqGO5oWF4hvGdlvpWIySbT
1vc3Wkc0M4o9ARso3dHuE0CbID+wnEPQspDSuTfu33CeuQZQXIgnUYreEIkeWKcU
WO85tUt+G2/POWZbbmgHbdoGQwaDD7Xi2a0JbaeL1PwA59Cn33ry7LVnaODeg6Pq
Akshv6yzZRLjOqf0BQe7dj749+0JqS9X//b33JPmtYFtoma4xnTQaA/PXyc8WX7Y
0ozXkBKRZ82cYnyBx8IVBo6Sjt0U13lkMXWeT+7lMz9X6hGQ+BMosSOP5FcbWlRC
OJ/Ut6bJQ2STtAhMsWQO9k4mF1lChzipjRCbmbnNNd5YCm9D5kbyQxzwl8D/OM8Q
sJN0/jFYQpldD/xr1LtRIhiWC0jbBoPO3vxiB8cgNBow57Kn+1ygYr7wePo9jJ0t
XDc0KJk54opVtpkoG9BTWiIF+nPaYLOcHQP2drwRqv6aW3S6fyjgtN04b1MaFZ5y
6sF8id++QzTw91X3f6hA6Z0rAEpxbsT/upQtXKEJjMp0UntxBfaPCbHJ63q1vl0A
f28rawOCVVgm3b50XtIW4yzluvuZ5LfIWea1o88yyob04LXcy++bpEANimC7NFRD
/MLQyJoRaOJt4eRXIb6bFgut2/KcyBmHUyQBZPOqVfEL7e5F8UYacKbgxvGJ6pLW
0pn/NIoE2hssqqP10zfvt6X2ep2jVND4M+beCl9ZPmdVd2TZyH/ao2BOiExEBDbY
WLRi3BgCXehMxYQGZkY8i6xJeRPK7B+xTw3o9WbjIxSJkN3U3B9NAg/jEutqOH/J
8JkQjMLPaSTmAvULitkx62pY2ePA7WbrM0lN81Cx0syRR2oQaPmHADg2wvPnB8jG
7n2skYmxDuYHQpw0Td84bUlRp8IzJLOw8k7bwNAKEHcNp2XijAryX/2GCaZGPEny
sqqVA24DeNzYw6k5ZoyT1Lpd8CQBPAwjDNGtRErtuD+ljLJ0q3e9tAJxW83P/4it
fYe5emLnn9d29vZfnQ429syvN07dqzj45kkfJwgxI5MYEUTkopALHhH/LbpdKqxr
BMepp5tLhaj5FNRaN/IUsILu1mJ1B6D9tB9eyRnafrt5xrVoBWPteJzArouYuSsQ
hEpBAu6Gd7eaKLUeRblSerOoNP4sZVbxIEObcsG/TntJymZbEJZ8lEnTici+oY/5
`protect END_PROTECTED
