`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OWxdqmXCUe58L+nXX+D/yfnFzUAOG+Cfrliy1bsF27v83Km4tATqduXCYsVYzf6c
YZFKbcOi5LFopMn1w3Mk1ui8dQ4RG/nhaen3Z7Z/jlL1Qyq3QIqC6iQM2eINHznP
b0bBRg03Oy48Eb6l0RkI2BG7xpMrnI6k94dkhCyEwHN8H6vKA2Y4qxscUcPQU9jP
faH3tQo+MJ3ZsB62e6LJTfRagT7+Q1WxidpkT5+n+hymLBdhfC7ow1QUsB7fDnV4
klHBCFptCGgjC6aowPTGWWqKEhq1WjiISGOPH+0dFBCVfjH6DEx1e/cN4/+ixEBE
YwTJrRxAeEW+TSEO65jdfDH2q0jXuHxZqyK5qPFv/V2rLexTZ4ju9OOzF5z4K5dz
kEuiivwoYhUtgtxphelnK546J6nWVtNpvj4wK0yK/hxJohZt+I64ff1mKdusF8PU
dtv66thdVYoDXvu0DvVEpe6zeoBYt6DLBZIAmFK5BCPbtz+CTwJd4+FuFsr3N2QF
uZH1DdoPwGxKaq31LvwDqkgZPZHC0ELC3GMfj/1/Wz8f9+z083e8ykqCWPxivmg8
cP2sh/ydZLqFSMh7TZMl1kkIKipGdGlWnSTeg4p1AstzUj7loO7jg54naFeT12jc
LPO8Ms+RxdtjseNEIuOqrqA8iIj16rtu/Yhhc3FEHzcMal8yJRT6xyu6Zgoy4saa
9/2Q5DJbIDKNZhzTFC7CrYSI+lEzmTwIwc1y2ePNzlCvtxZ2+LysPPyyuK65QArP
WApyONPlPi3qQNs/DB9uiXABjggIziWwgxqXRFkp1K7uwFADlJ40q1azmDPRakRn
aMEuepv/lmXIjm6oP8R5TNXn/x6THfOTpln3+q7sBljf+sGG/foCUm3HwfzhjujH
Na/dUxb60nr80P5DPx/QL20sdD7eW0Z/mqSizOTKLEmGATQlLtQTOKpOYK7DyBpd
VW8ZfnwoD8Ef1VC/lXpR8B/p7RIOgsUn2xyy80pAc5JIgxj2v5UIlsOBeo4IiAzV
H1Gf+aYAkhtg2tOE/3qoqjGk4waiw8BetzIX3nNMofPXs3leth02c9X4J5i3FtxX
FtgTr5STdBQbh2Efps/eCLjMFMFiwf8DypIIFREhn+99KQk14boXRLJY06Dq3Ghp
d2DjkZipJ2zaqdbd6Sf5n2Fy+4Sj2/E2o/LWsPvic4pzNI3Bzj4Lmnv3JAH5/Zf2
RTiVaZ4nr7psK/zuMEvsOk6lUddL0jYNQrYN46+plti/aSozIKoyK53xZK+mk5bE
l7yUzHhjl+Uez70RPKg0pivyQUuATsr+a4eh9+CvvtAWw3U5ivhW3WKk8k9Dsey0
ECGHhLt+GWkN6OOBftxHll2U6Ayl8Od2V0Px2HTq4DSRiB5cWUD7fS+1siOkSE5c
t3dED8f3eKW2/3fcbu5odeQqrUhI0vafePv+WjJ8ynIA1U3kUw2Fl5YozAVO0KOv
D+5e31d8LhIFNGuxIx2A5NyX3weCkINznvOJUVSE+tNtUtoNo6sY9pBlKukp66zp
+6MSw1Ej94JWACPzonEt3wEUwmVrxDCMT49VqCyBxjvTymnVYsQ2NCY009T8whya
hwDYfgbBJGHWBfS231C3ST8DwNnv5rbGtSO5BdcSh6pnQs6a3rHOHrTBQDgdJaq4
spVHPvifCav274a5kQB88OX11EHDgVwUcAoNgjBidZmZXOhdbo+uAqCIthWRREPh
bl+B/T2AbIXDhUEld4/O+1Ts34GLUp5w+OxIMZv8zZsBl+twXskUbhEZnsQTWvvX
JHybrvVDV9+PAQsTQkzt1v6PFQuKw7CaLLaih2AifcAOAyOJlFmOv8OtSV8IjgNW
1Tg4k4KmrW9YXvfcwHgPDUrrTqZDiWap/gRT2nQpBQhem/J8pKQIbeLzVN/GVrnd
44TGDu3HJcyHW9uLU1S1b8Lmxk7FipOfcRxNDQh3Vrk5JsaA8kiA3yFP4UorV9O5
4FHvhLy8wraEf6STDcnMjoqL3izKZ03HAQz4VuwcLXvitv3LPPqqnqnungQs0qEG
BO+ampakfRUk0HMrSOkz4q2vBA6znsaWBM4feHcTwbE=
`protect END_PROTECTED
