`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zq/NVP//Gl2uxIODG0aV4mDfmRmNaw/akLmpOD/5FzXls+4w5xzqodjiMvZZVMl
hAFWVDd89Ukkm5keYxLXMf8Q9I5ZffWESX++nC0wTsohha1FxM+aretxFcHcLlxe
J5mCCIsbhRjuwWAC/Cjs3tjciRkwYpll4KApqdwceA/23II+RCXTqYcp476koTI/
olweG4YKdVWd/4k2v3JEtq708gw4oWRlTGCM/cEuf4Ujll+io62td43CTN5VppNC
8/YnBqftbdqlwQNjMT0B7M7Xfe81zy6lHL/LpPGqyz6J2dh9OvXoqfI0h0W8R4ZW
MRV0OkYaLZ1U7sqrjNcrTdxLiLQtk6b9T6umfmTPQC06Rz65+Wawgzj58Mc6Evq7
mFU7AWBHfwF9bqFMI72UsxiQ6SVlesX0uMIAhcHVv/Zw+f4hUrNZ7MhtSAuXN9r4
n+y5+dJ4QVZuACrKki8ronLqdPWGIuhGtPKNt+JiQM4RD9MeLBZMo7kzZkqm1wVc
RcoDMf71MM5SeUsUegf+GGHJ54J34Hz8zYNdxVj0BULP1JOKtcqpm/s2U06fxk3j
`protect END_PROTECTED
