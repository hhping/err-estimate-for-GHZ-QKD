`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9J8bBjNJcXmdJxu0mGJIh+jKidQyp1l7h51OePSy6w2RrLVEZ2ln7on49w/tSOK
t34S5NXo0EDY8h01NOx50BIfEhjfTbHOArc3SMPMdTQNkrLa5LAHe16ORLOFxpXP
dTJnTMNC9pdmIb+T7RxbgrapJ1RmLxqAipVWRX5SthuJYCRioHG+sX4l2OQuHF/G
5FOSLF8CVHLWFq7dp8vItzYy/Yx4Hs0QVVFH2oE37nDXW+Kcv0ScbPrjR7SPH2Rv
jX6iI4ayVy7c24/AVTnnyOQad53Cw6jHVAyIkwI0ifOxgteyi6xCNUE8sBiMpRIb
CeV9zJ2vrJ5DuvM2YmWtGbwdBdNL9z/UpQ9WwjM7fWLUmgmbx/3vDkybTes9j5fi
p5X3AamQv9i2kOgM6yjyINqdV6bllEFzeId72otTtykYqSwm17+8hRuYRZ80aovJ
c1vNQS5AZ0eq3142BGqWig/EGU3gH1uxl+zwXAUdADBmcQdqWNBobqG9MyKNtgcW
KiTKRZ6knzuQjSIAg/Tvr2vFNKkakeSM6mSj40gkSDCvLEM9V1+BlyxaK6icXQoS
4IP0cwZWltOSsQycL9A3vZ2c9L1j1WXfNJKkoAAzMnh1z+OYuuG+NSWtQwIfLiGB
PvxM+4VdIKrZJLwfM3ZH+y9ECwOBhHH1OVbD7+3ll+y1hWVGgrqkqrQ0YRBOWwYM
4HxTZAyIiPvjM+2rKjy4xfj8zhqpWxCx+CN7XAk5Oqw7hxMU+pc2aCB+T9L55Z8h
T4RAnZzB7r8f/ZDsNFpxFbSSvO+IysJNDkKXIT2YDQ/yunXU5BHIk0ScO2wsurm9
jAXp4vBmHep526MP5e+PfJx+CtepCw/LPMS7IGJBXWPtFni8sLvaOBpaibkkksym
OHo066GiNuSugAID4ZIJK1KzcGVhK3d6Bllis+CRq+iWV7jDdHa/QDVUJoKN3vM7
DVn0EXRzQsO4sdP/d3eh4mHq8dTaeysCZgRm8Up4sWZJQtbvGJAFbx6kyUMvsrzZ
ECUgdKgXt5HXiZDWuwfxovLmPhpw+6YJYYYwufYlpppedWLq2BxDymW2Ch/uK+jb
j95Tk0e53Egs0x5uyO7u9S2YqvPRnWb/pMVwv2W2BDDyglZAMKMJFYJySZkaZ/89
7UIOWY7ls0/O+ZMfMhzxnDhJ47N99yhfnz0cIS41m9IGLlBx/nHV7wIZI71Oli7a
gfpERFb1xY+QbWV5glwUPEPzoR5LJWB6qJH9zgQV45s6XhhblIyaju8d/dSgtApY
YMgt6WPjcDnMlLHTBRsJ3YwD7ngY6Ndv5q9gzgrXR/QoyRBmB/95sxr37Qvz1VY0
Jsho351A208htD3pjglmqkGCCaet1YNYuUJLWh2cILoymQAYAplpmUEMguo1dmzA
TKTg6a+TJFwSSWUcjIvXCWpcMBwiw7q52Gcd+BYoFt3UOH26EpkVX5EhrkuTBh2I
hQaEN4DrSMRJTo64d8EUDi2WSW2ZIh+VjgZcXJlrewU=
`protect END_PROTECTED
