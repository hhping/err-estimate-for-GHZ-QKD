`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0sIdemcVhlizBqbbVWuby4tik2G/vZ6o2eUSwZE+rAuXx3SqoWmsAbzMLV/F0wZ
3pgFdU7yYCcteWStXOAjFs/WBE7DL87UHxDeZ9SIFjMchlwYSatmHg+ZeYuQjKWx
3kK1SpKiVTL+/vc7GG2/RQX1AIOcbVhbvF50My4VyCGx+CwdbAIMYBzj5BbZ3Jvv
8lCJfPGGmyAB3CbI9KyXB8rVwCfVINl116FvSE0vls44oJ66PtqgLUtR/w8KoCno
8ll/Ptqsq1BTnCn69GHSyRwfj2DUg7it4zPm3hmH8ojgB3mefHHnehDiJQh9dNvr
YaDCotZSnTrLhW/OhOpVRSwknV8wxWpfiz6njRMqVRrJgPItL93knd+d2M73tuG/
bHYGwJjYvKUOri68g3OtFGgVs3+lV/R52kUIjtWUJQVEOLK06sdWGWupKoDrokkS
x7gF3qpkAEIuMWJ/DJ6lj/GwCGlxh+W3wwMJrRxJEmveNCvGgm0MaLM2gaWDARnq
BxulYIqLqZZweOHCVOtPDy4lCu4G/n16wOxsFDOfZfjIGoKv379ZQtxM5dlRtvhr
9g3uwGv+zBKftPWwGk8WsOUD9T3cL1lGdGPrmX6i/a8jX+qCUrshvPBaTh4Dpuid
TxfkJFr1I9Sv1lCyBL4zF/5enGqY4wZdfRUg8Fz0R8y8QxXNF2KrJRWRMZ+OwaxG
soOZLtN1gEc9zrUy9fKxRlRyQe4824tL7QJZnVHB9ABGBgb/eNsXttcAr9LF9v/V
i9uG/pvm35eNPuhf4NyRizBNbp0vkBZmeP2qqAWGYNajOKVEU03DYJp5eAj6sxFS
ILEA2SxYK0Xwe1+2y+J5b5vTD3UPvH7zPG4oQtreqb+k6h8eRZ/YbY/Md1pA4i20
NMI0Lor41ig27J25puld23RUbrJtjqR+mA4WkHXMNX1bQLF8/t9jpzOydhgkpKsv
NyCsj+8egdfXw0pNF1DdTT7lFVF5rywcGp/OXoYgpqxqMGu5lHycvXqnW6UogGFg
87voBzcSh4iTGbB35OmW4t+v4AKdbbcLgALN8DP0bAqIbLNfYtQbPEbSWs0vcDui
ikaRh5GT4TijBRKmjuHea16xNJ3L97KP6F+I3QKTtLhpC5l0bpWcqiElb2OLTXxv
4OCmi527lGUBHoJS1D4rNWWIdniRjUzu89atWlkNngniyDuustb7x74Cc/f17DQu
kvG1bFLISPjiKUex33J4xn9HblaIoB1eqBfcb2qYnPpNQaJzVfCorHLfbpr0fFAO
vFyV19z7Eot7KqHy01JKJYOy0W7+/BiGFfUo172R1bn+e2PRNxtWmVd5OLpoTCUB
m19snMqj+zL+2ps9CNb1Jm3AlAC2kX1pny9sqORc6tWxZf2gReEAU8qnNk5W5e/Z
hNiGWDDW1ijvfeQ2WkfLjEi10xv32fmw3J269bpj9LLCX8Y8KdGvi7ACKJltaG+q
ytTn+BJF6Pd4qR+BsQb25gSWlQlxbDS+8DK4vA5SZDe5jHclUchlNoccbqp9ZFsw
VMc/QfeaegV7UHkleL//L6KWRNEz8jFZshcny724x8NMXOom04X1sWV9ldzrOhQ0
m7QGhVXrGoJB353EoEj/zczGkqu+xCm1ZbF9IW4VkMR0dnpMkXJYgna9IUCDDlJc
OC2+k6/9mFV6BmydhgSaKZWKS2pktZsyJi0F/UoWsDCRT8Bqdl/T77bc0dndiXYR
QgsagzKxvEs3qH8r46vQTivTepxvRJ0DU6KRYwZbpxRmgetSU9iBxgkKGJ63QnLs
am1SAd7m+FXnASH3nEPNidUJXu+KODFmBArYDEzr/sg5bRWQNDhXyq/sm4P63+Wg
ev28QyyRa6emKzIfz9CPgF2x32/iOa1KU412ZXmpXAvAvlTHyCSIXSt21dqzgbhK
7sXwfUsw4RTORCdifle2Auh1cRqleYydp4U+YmpASCu1Ig/hDYaCf1LJlV7WUXvP
Zr52/jzJrl14WVanyhIJBw6AK20flIIOfX0Jx9naLOY0TbLKyl5y4qhLa+RykK28
AIcEEYRD6wooIbtEFepChJFh8QX+eYDheL+Lbys3/+br4a8YqoWjdRivrFAY5t0R
qgNbLD+rC3Y+M7H8fvGdeEJ5wJzMDS7CUizrwa8U3O3hQPTJeKHe5Q+vwlwKNCVv
hxjBl9Xh03SmciLZjiwkQXW+Ge37k3asCNFFvLqfBexatnYdGXlHoVSiER4+aLPg
hb66FVtt4Up2vuueonKIyvcMt+k4UE5aszgD7F6qvVABOfhQReZRGYcOzk78FKiB
TA2w4vhtf4md1s62a6ASCQryOD4zwT48eDrOAcFj+gBrsmbQQWOS5j42xK12u5Z1
QSIpnFYkwejoJReanBHxS/xM9gy24Seq8M3Fw3AqOO8vy5tE7/dkLcYL0WfbMXXv
VQBjndSAStnrYesmItHziM0eXkLZuK1C7Z2NnhrxhOO1V/iJhaxOUtQ9Pnczc/cS
ganVytWI0NMWP0Dvo7o9zKxK9K+vQQe8qkUoI15lVT3N6S1bckqmpvwLFFpxG3iO
zU7DBKRoieS1RP8FWd7JmcWqTI9Do5mUru0BM++F0EI4++yBEdnn9Q478mrGsDR5
g2WFFP+mDOEhxmCIEyN9BJ22uUpedtT3Nk6vXfNqpeU0oCsWoawzOY4VceXJhEVE
2oH2QFYLujtEmJiErvqxb1EF3/NyfSN7H7/UttU1O9aUp+9BiwoF9WDqqHoubNP7
KjTPmrZnZjhOd8OhT5VcGxsvq/WcP+XmMtNJe/RstabGKpweiFwz6mKsfRsELMZX
LCINFa4Kl69HqUlBV6fiEhB6CM1KGvHFXX6lgdQ/rSvn+wPD7VgNQML/jFZlo31J
ScNkr1/3l4LdidXB2YaRsaqceENxHZdOPpUdHMESRxSIUu0f2Ld1rE2iVbZWNVc9
CUIZymBtaB1VaEz1MkzhsR7d7ZAGmrraVlNtq4qtSXwb7VMXIPfkzMUrR7dB/RHk
0TEBo2+4Jbgapp8fLl15vZE/bOjnpf6U0VwcVAXo5FM+NztNocXNN8l11hWuRhQ2
Y4XK4M+2RbQFe4Bvc8q5p18gcMgUSLq1XXZZP7mwNqe6+jwxwv8/ALOSdggaJDkM
Jlydcx74L6KA+mokx1iktcrOQtpZp88Sl2Qdt+/RSCQsQlt3o+XR0+AsjXXQEx2j
Eo2RlINzDc1AbT9VQDrjIwjzSMRnRvI5DXphgWUeYCoZp57MEQUoeP9yVZMiqZsq
EC/GWlfhM6QilZrdOVgpGnK01mwwq9LgPa3rAxffXR8v1aMDeTjThELzvBJYGsfX
EcmcBVT1gWIZKCTtkGxH2vfnd/Y0zanI8lA0CFoVaMtlaoPqrKnGL9ZKG4/PG2df
Ntrz/qo6+zqRDvBnGXgxn4OQApN9jsPDSbO0/FB92S1j1DECQymderbgyrxGatG6
AtmbiuOf5swySAgjWQQmjhbZ2nYeL4rWvXZjXRQM++kIHA2fmWeJlWG+9tg9cpw3
YSdMXba/FMHXcJ06X6ZTkVfZ3JYiT0Iq+2x2qR0LWzxDg9rLvskJbTV0s/J2MaCV
0CpPW2om9ePEmOF2u/q8oFKUhSH6Ss2Q9ktyuvIp1bPEehDGXr9e8vxojly1wtsO
GXano6YMiNheoFHVeBtrWiu+x/QKkGd1zH5av5jTi+IwrrdL+xkkm5zlfhg01jOP
cVdr1LwTJDguxe3M4ReM8KNKv5rFgR6Uvs8cRnhlIT1Om24nM1SuLEF6gkHwKmSu
yV4a569DNtLnQN8RzFzuhHVE4FE+z1134ScisfcGRHjQmMKT2n4MfqTM0I2iUDk9
p6RmcwBd9nrdYkoEixEHMyfGG8h/rTjPrAxwmhbnrrlFKsQJAGeaTv6IlX7rz2+E
UpJkgIlnX45AfUXGyUotkgzfEcARLE6aEjmZ/iXEcGSgMqQotSBz96+8JqZXv4sa
Mkf3FYIpP34mdL4QrdmwtMeNZ3KW6fVcURPvIh+BHBBXCS2xiaCY7tbEKveXt6Uw
JZoA1Dz3rBvMsmPdaczEztSnBTzmD7imQBAIjdghQy1ZKD5BdLmeNU0nLMnuG8Ez
fF30nbINL4vfLb2RyZ02x7qO5kirSvl1lISEx+p9thQm0N03fYpdWBch0nKPks/h
CRR1/ZcfS4urgyNt2Fqxf42Bzqhe+oKEp0oIEJZolzAFQ+4IF1I7zLOANXsQxbEf
fLhXswUNvmHDQaZDOUaoCftM+/mpXjlXgxKPxmmPV4nfwuBXK4rQk+yGZ2kbGjTO
xCcWBLXNLJcsY6iDXNST0vWWER58d/5eSNGsX1JmywSiQmjqt1xJUtZDAVQbCGsL
q7itM02MhAi5zmjIcPm7efzMOpOhB/NpBcOZ8Ig3N8f9oL47REqu9lAX8xpBlAal
a/JE+jctQkTr4ylPizqcQ4zz0FajDtaiA08AnOZT87stFZY8TxtcA/A2NIwT0TyB
k/tUHFMZLK+PAeoz8LQB6kYZHm9XFSxXtZlSaoHgIkU2EhLPyZYzI30Rs2BQFthj
/z0S+4ZAPCglLDbPB84NGVvVASk2ACBei10YgYy4mDKqOv3jNOWTk4mLaDy0BEWU
cw3ttLoXJUlo6RPhyDMcrtGioeOvHrPF86JTuIezNYvqTWGO7cnwARbUFCkV9681
0iPLU3IML8RVLOi0W3EyVrqRTysAQ3kJ9QS1otiyRfxlsHIpxi3+RwEEdB2iFYhU
isD1JLROAVNDTv6Ond5kxuHXjGmYAFHe0g39cCblbwVrQksmDULOcufp5eYVpdqy
JCZDRWiBn9f8xty1lfm4DNeJyL/ehbjwPtd1OBZotTMhHmNBRO2MHuKxCEJ4ubyi
PcOvQBDVIANbRn+IvTiAO4VL6gSDgA7zQl9c5FoInw86x/UfRpmbju9ROQXyyxIS
bPtZWlhqbkqH1IZKnk4O+65QXFldAG9mIAqDSoNXdIHU4vklsr91gXcmFOmTZTNO
sBmo1/GhTmoDsAtiZIRl5INoc7NXTqJkVrFk+Pi+jj90+DA4Q17E4/4XWpKOJx+h
0pXM/l0EvqYh3izT3gDVvjldVe3xJu6dVAkdkMukWO0EV3Vi3oxpE3ODK/USeH/o
LsRwG844wtJNuQCxAamDxHsu3TjjwtMiXGIiA+m+CEnF3mF0coObLawMNO+WPXoH
lsBMFyp1cYU3Z79AxrI+dAwXcsHkBiLXQsl5oQYf5g3dQrwjyF55OR00qhBNNko6
rYbJdnqeqWmPFHQWjXWm6CMyd0/ay7Xezmv41XukLcvTLd2pP+YXylLQK9J7d1zR
3MZKpHy3yFCJh+h02WDQV7HaRGfK68JbWmxG2jlkswWb1Ykd4jg9wZq/jvTeZMmn
uy0ytJzWrRtMCHqLUGAPnDsW0i24nQAKda9ygXTnQhJLZgZmEQAiXGxbU/ULOaVz
casNBPTqD9Wg0A+l6eaSYbYfBnqMezB0Kr9Wa+TDPM3yQZEjyeI7B+ILz/MJ6ODg
n6dHpqtCYXuUIKFg+tNtll2XrldtJnj03QujoG4wyrfguQLI4suWB8VilugY6Nh8
jm3+Hmpv4aG4TrsBRN58iiakDvlUxSQClzpKwhHSsP2p8j4237EhsaSt8unXVy/w
bXqD1DyflC9/G3GTP8EZDfJTb4Z3jEgk9cXRG7KFn3s2wteTx0umq2xaDb5FK6AI
p/T6HX+eraaAFO26BKTIgHrjQq41vCDAALgvrxoaVH9i6TSQOIHiMFly+Z4h5nH3
Vr2DrSSTIHauZwfdzxGxVxNUVmYuElVsjP4ruxcDJVQdHVk3liEwCTPs5qBaDnJT
Wq1y4KPOXxSUoeGqKamw7RCVDQYdgI+8jbVXOg1A3ajAqGLWALB5wxDDgaiMOUHx
PDn6FUzXeTHzdQ1KqMEvp/m6lqGwVrG95fB2U/pjoVTzmk2LA9e15CVlm5uY3ah2
MOvytwMqf+ggeB6dkWAnOjLM0VVer5anBY8bIru9bqUt9CIpzPejNny5rWgMp/LJ
pUYsuVCHwI3iCpq3IMmZewKp47BG4/8OMZTLp8WpHdAoQsE3TYJeZMGJYdnuKqQF
n5aaqDPRyicvKWog+sHR3wxLPu+9rTBc0B4g/3SGi1Z5odJ9lSOePs+oG18T5h7Z
WJjOdLEgpXq0DlpqJOvo5+iQG+4YmGfsPyXw+cAc06oTHqJiZwGB4SSHN9jSzTU0
0kL1zX2Mef7Qgi/IAD0Xpte5dUo5TrpejUI2r/q03wmdDXdB2QYK3NI4on83A5ja
QiRA/gkUgD83zpBkvmBt7La/eMeIoOqPEJmk9gaRnGgCJ7gzcexgxXm5joQWtTPd
za4kTo3/fH3AKYIzfWvJpFiDNMLMoVeCh5lH79TW9U14/Icew2u0nD80Fxvz36k6
Wr3QRkvYKuf4EjJ7Dlg2EwA8TtHud53vAnyF7BEI9JYGGJ1psxHpjD4/mFvSDreO
TbhFmqiYCyboi7gcms9kCy2pOVS3D6BeHmbq5TodLTJQmJz97367IOKOZ38FUpX+
mjy4pqOU4SsOx5ngEm1BL1+U+jPn6+ZjQDvVnCO5cKhSkb/U1gJRRrs68GTJq0Jc
TgRXK8cSIR0QF5K6GBO/JvykLQ980ktGTBomiN05ROpDuQRwUccf8NbBzUP0SMQ9
pDd+Wxd35Ybs5ewxua18I69JPIXsTlFcYjaC7wVvhmxwUqfEqFkBQyrzZb4iXCKG
SaFVXHB1LmZwvE12aOV8eZP0AoCSfCbhK2kqrvwgGq7Ct7cu1kBYX2uGfqXV0Afi
wu0NJJnqUqijHzrOjmZlY6taJz/kIJAd2MmnubQuwiPMEsaMXOXkr8+Dr1GPJ/sJ
P/eRaEFp3kR5Zz/Xj9xfzvxbpGm3I/dGRQkbJ4A2viKRG3vcj2+g677pGkaoeuFS
+j7HMB1ov+9eHCShT6d7EP0l7XlvFmny/mQ9sy+KW7rouKVinOyQHQ32fr96+1jq
699PH1l//F/4Mr4Wn/5zluOrMEqLlqjI9WQO8A9purwqai2NlEyaYPOPhjwITPdU
8Hu0HjtYr1velqljwdYldcu7LKkWrPR+RcgYV62brtIz84VXwnAdUvzwnctak8/i
sD8lYze/OYBTGh/yq49aoRH4pbA7OtCVZbpOVZkn5U9DdXHdoaCRApEAxu/YjBBi
jPh8zTftUGEarEvAraRGAgltiY0y2qWcpEOMW9+DO2hpdIalhmuGcnxhnFZZ4Zga
f73t37puBclIYdS2UltKfO/Nfk+WdK1by1XxzXvd9KjyB557D8Fk+sc0Zv8oHuPm
eBG5hT5yim1R2HMmPv0IBK9U2BABU06iskhqPl6B/uBaGhdj+QPTzn7/yAMSCzqz
2C0xqU3CGthbNbHjDCxvOPb4mTVRupLy3lc7TARqvVSBMGbWO7UA48Na7/8EBSh8
soqR9A94mRNYAUjhDDcncSSPsVgGb/ZrQxNkeEPB3kGPxBarQgdk910QpQDWq7aT
C5gziU6sbSBG2Tw45Kfl8Sn5MJR1psMixSNWtBBag6xVlTJKQ3uICAjJ4L9cdJ+I
eQUoomMt4elohX4tWC++Y7NfJLgJ7Q9luz1SfmUQC+TkX4teNq2ZG2ZmlhEd6suY
aWctqiwgu16K5xUn7hbrQlSWY3uaBVZOdRWOmQSw4fMEwNnHwx7a84BlvaaaX3yA
lhc82r1w0vj3ZBi+HsFNgoYb0I5PljT+VmFha4GciBBQ3KWabtwSIGwEo7gqefGq
1La4/oK8l7eBTBSYbeXvO7F/qh/VAAC8Gd/KJaMzvHMTlfqkvbmmtJm/vHEPZ7KY
gxYn2Xd2Bfboihli/b8Qh7KNpinE0UJLS4kq2vnMZfzzDgRoCl1fjCF0tQJvu8HK
Ut5sZoRSt3jQ43j5rg10Fg+0v5LdhHy0kByuFJk8pzKKSUG1UJP9g5F1TtoT2td4
GDj+1PpbGLuSvI7iSYXfJwKEP/67Bfoh5+knpUnlq1fRvCuQ+2mbqdcStfhV896t
+i4W17H2g57UYRW7WmEN6il0s5ZWTiw5yZW/qO7ST/09zr0Y+f+hzESetOWVJf37
DSxMkr8BFf1eC1y21WyJOCEd5V2QaHaWwQcp7SY3d1h9ydLU/Gnqd2oCFNVWiSex
gA0pa33A+ezBzn4l0eh2PUo4zse3u0iSenka6eRJfk4TORGKNacOf9GAuWq2GQpT
A0I7sG4xyuuc/LFHbdJtmDx6hBk82rasIl/NEKulodfHTf+kLlB82mzvl603vDP7
rxukJNp9hrSigKxUr/+zsB2pVu637wc0Gm+j/ELGCw6zDtBmk+0e1+RLh11LoWZG
6XU6H1b4xhNJo3MiwVD8+BmpfBYo0xKExXkLeu7w4H0HVLR55b9mCtS0t5TkOf1T
ZO/ZyBl0Z2miLAQ8TBbnBQ1ip82Im8sqYUgcrQeAQXw67h8P3+u0aK/xLec+buno
l4Bv5g2xHMNkYUcwIcsLdAsgydqU9MpDD5ZIhgY75QWcp+6t1DvYzELztysFmB03
+VOjB+LOJ+flaLrubo8CailoivZlMa2njkFvsdiwMUQZjZTQCCtp2Haidki6kPdm
9XERMSVXPSfvqbSEhQpPglnMw2ktkrOol+UjLyWYK5HZeMfTUadli8CYgzl74IUu
Zn2Wu9lSULoqBkzLW5Eef5oSUXsjjNwTlYFI+03HvT8D6VH1rlC1qIWIRiH56RjI
53TWNISsYiUAfFaPLXy1wxhT2hykfNo+8bxHpph35faQd1CSdldGsWRjY5py3eTJ
oo6zhZL/aRXKJvfx+0rKibhR04VYFvzi/6AArLcvIzVV/pJGmZbNWRUza23gSwiY
UD4q1qJhhwVg+jN5x66Xt+0Vax/lBRml1k5JLepPYn7ABM4hJ/eYKZ7cX7/OTYdc
jcrKDeY5vCRGgR9TupY8zgI6x6Q5qjkNGeJqBkE7Ne311AFpRIeSMRLQvC00CuH3
M1gweuAvrXj/+rhCCUdiRXv5cUk21KUEZj0zMHmMp8o8FcOfMjwyasMPlta/Sr+4
7MLrDxbdQUNnqSKx7ajD7GVRi8Xjh3F8YEGYw64MrJM1cV3mmhGJ99XwmYAJ6z6s
b/L6EwahEpNuOY1uhrBOKHDNdi8WfqOJGvMyDO9L1UADT4ANng6KFibcrP4kM4zU
3y7LMNRLJ0mM2lorrKpEJj7mLDZDJ5ZvebYA9qeubDX7K7bZE4QBA7WTxoepN1Ba
GNn0jMDUY4DEie/DKq2MHzpNT/6xy1vBBLq0/BT6V2VaDwDbdeba6J6fQJOtd9EG
EFO5tNBLZTOB2Q61iBc6YAA9vHH7y2fPRSsE9z43GvIZuFjnZA6lSrt5Qa6u+I1F
fTl8TKNPONFcZAY9LHXyYwAeGS88z3jq3xpa9iY0U+aq6EYzPmzvFjTta5BoQ7GU
DJhWvW6wSRCezFGR3Y3M4E/u/8B7fe4W8cXIHTdfeL+YGAs/aQFYzPRX+klbqNLL
STM5owVWTFnE+oHw5943RbMIaHgowQZ7PkSLU+WbZ95xWCwtcEZNclqoH1OUQz8x
aZBYFeRrqJgtq+En0ysi5obzcJwDswfQ+gYqDj2mHc+GijrzbCaKhRHQiI1wRrYq
ZH5nqvsrWTxLU4GebzB+yzh5/fcGiiWXT6hAXkjJwquMkE5cIANh0y/XAaOv9ale
v6WITV5vsImfOnGAWvw7fT29N+oQvdp2atEPxrr0a66wI86hzEfHfdxX1yaH4wWx
fj4OyyU2zGQJdd4pB2fXdkUZPyEIp55EAI1z+LQ5cfDyG+tnS3uHRt8/aPlwn1AF
K+9CrBmFILP4xuC0bkvckqHYqQKFSCInazg+VcUpelP2/Mz1fyRulbwoamS5eWb9
xYyAJTAo81Ae2nGHqQ+7BRHVGK+V0X8XUrHitQMnH+VeVm62RwQm2zjAol1hjA0r
7JgQ1bLQYHyhA3oDXAKD2Ej4J4gZwbt+V3D9FZ5HKzfXBo0tiKbPmI2mxDEFlJjh
x1sHvMxZrDs6a4oYhgcpGwbtX5YywT5ebkY5dIaqr/eOA42k7FxUg0ybFmId847P
hCiHhX1UPq2jPxweygFBMrJZAEF+mpmMdtjFMIUKJdwJ8Vnx/P3CwJMZ/Xbj0pFI
9kfkkGha4uk5jSsD23Y5vm2z6NfvCOb/QSRxXKgnH2NTvrl+OwlFpYmp/V5/D93R
+s08dgRqz308g33urOWcToqwM/+Sj2PoLfYVeLnOanIzJXJ92W5grWKdxHTtIeOW
Y/OW7hlZ3i+YcNw01zkMhgphcVT31g+a1/6EHDlCqJpSNf8otEn18wTpj/YzYLRe
qsUweFDXYsCxWxa96BABTtMYUGYO5d8whdVa64qeRogkHAxWJXwr/kCcdfFiA7Tj
kADMdfuc1oc95mU9xz9CRk95dspDltMd5635lh2qhx4UL5auWI7xESAIy4SZE4m5
AwLin40uZZ/0z1Vb/klJXH3I+NEjK4m6OVdRCny8VidR5usjoMWt/lPhhYV4FEA0
iH9MMpw8MnfWLANt+1yGaFB+nXC+Ycygvgnv53CMP4PR5X4RPABw6faGJ2+PluRK
tPf782u9P73+Uuk901S0ZJtVZN5bps9zRls4+rn5iqxhHXfOccx10o4uTZxfafKQ
YmGGGZ0ZT24avYdLssYj2j8kWK7g7eX4luftRBLrYsuN3CcriGvhqrihhuOeL6B2
aVaHkU9sSVE5TkGOm9P6tTAve3bluJW+3tfTjEAg7BLKdTp7KR1abJh7TeGM/o6x
N4/IbU+PFNeFe9k9tX7L5uSG0+8ANKQEz916Vfi6lnqBv72cw3MaMSa8RTKZiVUq
blhFUQM2UHs8QbFOXCByK5PfsUlllrl4LYxMjOhR9Zi4SDUVJ1BH0RZ1unLgU2Uo
amoatJjpNt+z5c64XBriUvMbdpSGnSaE8ks1x387y8TrOtMniJM1fnfuVccozSkd
7MAbhiKe7RVUbeqQbg6v07O7Z5vlX56Fd404+zX/EYTnjnkqrw8u2gMhRS7Qh36Q
12d9ztGjCtPxWA5Tk4fQlS0fuA4EPOU4wD3xK0f3B9TSwyb+makamIo71seVLEnG
fgCtPhGfytSEP8TY1LvBZldLV7bRXBJkW5slRlhP20g/f21gB98qnz1bK7pGMowm
PUY77Od55VkGZiU3nM30ZRuh7sS92lw26pECBxXQF8IhJQOlAgYq+eloCs4y8+CE
Eo6hb0+KxwIN/juh7vThFqa29eiZOiDdrW+sArdgQdJEBr7p0mS39vvUEFxWhy48
koXxh/e0HIEcAkerW0E6BLewz0USS4TPG5iVVNFB7UkgA23JyTvx4OYTLlNrdn73
g0CaSHso/Axz3FdG9IMWhRqUruWPmtvDuNbE8AC0X69+7XTjdYN6GboAglo1DfkD
46y8gxKR+ukEinhoVRYcNcvM5CKqPUyqmeqCTghAjHlDPJ59ttSKYBp+0NUTxcdF
5qXE7T5sm/ZuV/Z4jfjaeyzgPm+XoaZn5wd5I83b8ykMVLR9RhJE3/aTq7mb7gR0
suQ3SXb609LcT+DrH+nT0n2C45tZC4ZY8U0h63+HBFHGakKpE98cZsk7yyZJKCbH
G3+sYuMobO6m8h2ceqPU7gN3PubSRjG5waNHbQMftzFR2k9I5RSaIeUbpnNjtDXa
iGlaeOr5jeNizE5GU7bYstThgQcGqfX5ZVVcA0u/yYtdjnMcCSDn0kqSr8bVtZ6N
u+zRk04i/CfuGGZGkr5SGZhoYiEQbfcbk9TgOUQO9VWqzaaFeyDTwGIylRU1VDN+
HfQRoCwPbYbA95p/TXtaCUgyC0O7opBaXwQjHX4dPrmd68e38VlIPbCNh75YPHgU
v8V9yqqVxDCjfn1bjxNP2m9J3WORAGx3OZ89+SydjQsZOdI4l/NG9sGLhLGXoagN
WaB6oJb+cB3B0mXbWwP/jhOd7RKFHwh/xnDsc41mD5y5S+KEJlQsfPiyZt/y4Xug
6HsyawVnpgdAZSZe3j3t9Alm9ZJDNMwjBnA/xjJQ7XeY++U3gDHJYRMPNNEhggk9
yx/OSrqRoqgymBV9FhHHeD3L1UKuw98O8HvgStV9qQr8i2AyFGv0bCiwpFIDWzUe
3ECtSstn77hPcxSDgnh6pTQyRnRZVMk5pSoOgdh9zAo1D1f6tlXZ6B2h6aA8HyK5
i17wYl+kOOcmV1nQFHBkPgabTmreAFdUSpJpUWDW4KdCvJZzejCkcK2HuJAmV9/i
wns+TNOBqaK3uHEO/OhmjnSaq6xOk0yHJUdjEz8RqygqumL8eI5CrDNOQS0AaOYJ
dKdb+2qerADu8AmYI2OasWTmSth/aQADy+PuRQSLuEG0nniyWLm8n9GtJBZztzs3
GxnUX1AkPirviEiMd12c/W9B0mjoHCCnagEKyDpQsqStK6XroT/vbsRVJ3iwz5bG
zO7Rb1lV4UJd24wQunLMfFMNUqP9vOJwtlk/CakYiVMXS/VmNNh+tL7q8YbOPylb
0NCk9hX/1zy3dGk0AuwdS+EeVGe8xRI1gFx9lM8CBfpFJ6jE2iT63/RKEw8MgAJT
JbVhZ/oj2rxYjixREEdrWl2xOlhO3zLtA//tAF+I8pFfGmMo7nLKSYBo7r4h03NH
k95UJVRjg0AOxe0uqtxU4r8Azqhk2URg2ZQscYlApenBeR1d25UgCpiYQRTNlKmu
rhYJe20GKPoVixK6E5RbqopHLlh7XLEc4c9EPlW1C7kDmCkSuHzgQ1+oq2As7yqE
JFCVplk7CaXB9prj2IUhgkX8L8h6qqwyAr8HsHJSbl4I5MJ+kTXE6IY8RtUUGXbG
F0Xt8fJgdoOdG5tNqZVXi3MK++FK8emT5yhD6LL7siNDfU66ii1ZRywEwuDSCvU4
/dZOkVanAnt38AhjKKlefw/EtY8rO7XnURFDY1WUL+3snR/qng8O+ZLXu/Gee+g9
qYAtOL+emxb6DoBHGwdLQuasK+LLxfJ6XXkLr0hGqslWRdx9XTQja7qmCelTNCl6
UbJrsX9kdY/ZegqogFDPM2bcwP6no6m8+EwyMRuQAtd/z6RqijHPt1XRJA0D3umP
wcMthySusKMRDfSfx48EkGztbzLA17y8mAC3VxZLsv12V3LF/Mq2B8S2wRoK3IY7
C6l8egvqiQpDiQZ0WTi5TxnEaJIEjMCbr7HF7V4DfTk1Byl/ZNy9/kkzmYAvMQK8
zbZyOsc1/dzmvMjGFrmYYtQlI5U060FBvw3nVGVWIt0215yg1N8j5xL+RZa7jz+n
zCQ0SZrf5yCDINsmE64WsLGqfghrHGwkwa/z7v6XkGOLOR9gUE7gcQscl1CncM6H
9bomKuS2ZwFiDXAZq8BLndPG7V+wjTn9FTC2Ddioie9a7xsPgkcFMcNH1ta18ZmT
`protect END_PROTECTED
