`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EeHC+zt7VqlnZXu6TNtJBnhLg4X1a+M7PL2K9ufGjGBPwwOEjFcj9T8N6URDL/1I
MIIBLhWYUhVeCJAtsoCA+WGz2Nr2bU4d2ixrvSnm9W6kjrttZA3clEpooKMCoP48
dL9n6MKoxfdcv7gegO5gQ57cED2SSDg7IUczJVRdQPq8S6GA97Ms/UcoFUJyGOME
gSXH4HjP0c/gIGVYymSdlfm6yY3WX+g2V19hya8uF2uq/iXJn9ZXAscDT2pBf+4f
1cIpvyrDF82omnf9oDnfQv1qwGAjeIAJU9VHcmCBDkmFQU+W/Vlyg+cMLGVvXKT7
AqH55fsRGkXp1WCbTMF9N9BJYnkrDabtZJFB2ez4mSymGrVd2k9YC5S7ecodVEm5
HXNsL7HyfKkmW5jaJTBBSZiEYRt4bOgnGOsBnQj49SPQy3h0eg7/A9zXezUnWS1j
4Uir1M7IR53YzITfKwwbmNJmUM7HmbRfkPbRdVpl2/1UEna0opKh7DU2S6umQl2Y
9e6QmiqniiLh2Tcrtm17EKA2i+cWYs3X8xUQAKn1MssBW+zpqdJq291jKKGLP0GB
CfGxgCPPKJVKVQ73Sr65SQPPZ+AUlSjPJyRTNXvwvQZVvtaM7sIAbJvqCCds6u1u
7m0BvSoDh964NVz3fuJL3yXeDu1j5Nq/x3eBF4PBrohdHh64TQab1ppzE7QqGDxH
v82ReEdGOIv+WtK3jok1DN2orbVxbB8tutKXf9pVVu4mfHttn/FNYGyS8A/0lZ8Z
onA60e5HrboTFvH4lXx36Yy4vc2nw9ZzZh8FhZWk/SLF5kSvG/GwjMRiKy1tPdtU
nOUJ/bzo3ZQiIRflN8LftTDmFYWiGp+vk3Q5hUz6zkcO/Y08sgvehlu3rI/eLNFK
ywAm992s4mfLqjROsIHOY1dgMfxOOHC/XHyRacmnCpO0gr5qCG/5IMCgvsWWJLAP
7ZfcjWhQB7FOUQkkeR1GFwiMXHgDTFSAZFARPJxyjNy3ER1pSVfxjJvG5ay8j63H
xCHfEZoMGOeGVvh0vogrxW06JLwykhw/YyoyQ/lSMyaGkHfCgWupvjBQWfMDYAUG
/ZxkR7lOfq7cZGP3UYMm1L8LqGA5Ae9V5Mc7QInw/Lj+v4tS7Xw/AefNg8JwUx03
gD9DOBr2ZXGHZypOA7WYymZb+RjaPk/gMiJhcUcRZQ1Y/hHtmp/bceSiS+Aeoo63
L8PFusovFXNbsVlFqfxqO4f46GeofMoatD5CCRZZFh4J8GNmq6xElx+qkVdaZ96k
oCayxMKSs+etgOBQc8/qrVdVNy+nvinn7ZCv5deB9QJ1X+Oomb58e5YJjplReFzY
ZKBtwrL7u/wHMHZ4sApVy3/7aMdHq0v+29zNuesITGhx/6Hb4h83Vv7VFsNlSnVk
JvNYcNg3q+qk0xM3m88ajkNV+11BWTdoWkgOfqOu6n4/n3GORH280I4vDwpN4L7I
0kB6i2Lm74+Jvgaowrh0eIucVBPFhW69fYP0f3i4rfkvTg94LCo7uFndaz0ZXrNg
5UEq0puz9KO9hqTClpDlssxu3hxNB/0lJa5QgNw6D1cQIU/1ynbeoaUQSuHMaQVI
okfMDSH07IoOoPQUs/6eKCFLQ4qHx6GfijaqOVZmMpndMuaDZQLBhv/YesM6eZDa
60UJWPj2wN5iAqNwsSI25TQZMpAhkwmlhwEq01m46FDKiAJEwSQIuwRhSuVrmdtw
8QyNJD0LKYeTDXQMxU2Zrkog7LESBB0v1UQ2ONwcN2I8yhoWDcENqmnLt73NW/ij
7GJNjE61VCoKML8fDBAZSHdIioRSrZPY6vIPwwu51KinBAZlzZW8WGNksUt9fCK3
QO5mHIen9CBPlZkPMf24viL062gw27fZwsP6sfrL4FEcNoKLJVnnqeU+3qN5r+EZ
is2F7uuXnGYKDfI83d5Lk9XeTkRyMRPzM62BX6sSuhAjtq9n3zlVmyJmEsSYBXvu
rFI5Me1c2PAsak8CXe5RsXdI0MJIQqWMw8CQ/ikxVP/PhoJ+OBfS7u1A2g1on+Be
9SS3XKvT3YyYWMSfcEU6LKb6QdhCBlyNrSxtP53RPZ9uGrZhR/Auj1NVX1v8b0ID
LMLsTRjq8f9D6knTQvqAeQ==
`protect END_PROTECTED
