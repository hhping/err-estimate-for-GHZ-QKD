`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cndScJQ/75CEOjhugEjufLVhVqyOusxxP1XplWxbZYohjQWD6jz2B9BLJUySfwm
CQdcW5xZu5RzdUlQ4FwJWlK9VZtfwOMWJvC5LvCP7uJwK8lcgygIP6Gmdldu52xb
Sh3Jno7pbX/ZARVKvlxX1kb4qBJvntxYe+N4Js/u+MV+j7l8v4O9HyTbbNakQbIN
gBA9yJGLhoVSX8X6b+2juBAL8KV+vNK/+3voDnqgp3rvP5+vlOk+LmbAmmrOBA9P
HSemIxUGJiKaMN3P27hA28eviJUhg3VlxPCqfbeOsHXu3KK1JIfExaAgm01vGZMB
vnX+8rfn/8AudcqMizgucqsRhNlGL+6IGdugYuMGvRaGT7kN+lef+7MF/3PtgMqs
9bOLZOs0zDVcH1UwzdFceE9S9oJHLV2SbMWX1Rq0B4tZJ58xyxPXjHMVWxMZGtD7
/vxwvBjlNq03C3fz4yeVWJcRbAPgTFkeCE9OdxTSeDBS5zqSj8vXh9/n30Lg/zn5
BppNLP4qGq/o+dBJu/1WL3vGZZv8GOvqKI+SdGGGEaK7Q6JmdW4x7s3snqfd72mJ
c6FaDJ2b09UAVohvoO2f0nuvXTraKiqB+wx6sftkiEQVM30zwCoGcxJre//9wm1l
vjnuKPUr0TFh1kl79PHJgQed+6ZsCYZT5fQjbr0RbiedGPOneik/wl+VRg4MVUBv
siuD4QqqzNNgRhCWNgqB4Y83ulSuFrLuYxFuzeG5PgPdFxKVTCbGBsa5Pok7sqlp
b4upF7lQVVskm3GtC8Zzvyh7Tv6ShwgZa1oZbua5W4MRHaOwz/R30HK2WQcdruzJ
e8iYau2h6M8fnPMfTkHp6LOg4uFdHefKxDZJRJkK9/GWZFvk89dQ8ipm4enacE8R
qh1aiempkmsLRaA7yqrEruXsXOhM5vK5A4Fs3wD7IPLJQtTmMUg7sqbJyX4iJZCK
T7brFsVK8BQ/Qyt6IgWNR3tRPV30oQqVDWdoALWmEAhVP4k8mEhzS85Jx63CZCVP
gUdeh/6+LQdEiONN67euTH7SOkkSfi6j8X2WvSxbWYXBVo0nQXq0+5mKjnRRWhDf
Y2nA1bYoeF7YzThkJfOb7LsxxySBL8aY1dP7JiyQ8xmBZ+CEpC0iz6eE+Xi+yKmp
/kmubhQ4IAAv7FXGT4lhUpH4AaBqJXfPj9ycmjG9Ppr95fInyxBEdguJMWGZx4Bf
zeTGgTyIbmhQ0YyQfEGmsZ8m85jS+QvfPdNPjnepda4jiHgvTuAaY3gi9g3n0203
GLbtOdEuBcFj40W+xsmzmsjYMae6k5bH6Pxfd8kKVwSCe+WI3V6BZOqMgh85FeTw
n22dS0vIhbhgwRA47LbN8u/4GTY1nzUZwqmysx9v2lnP70zbSi5YJOKjx3tysmiy
P1UoHAVKJZzPlr8/3iB7euBSa2giiXIPeRDCUizPaTHL6Gmh6WSrJBr0zVSuylvD
D5SEkkzUtvY2LFQ9OwcSKc95JiSdZBdMg/z24+BwBJTywDD7n7i7ZpFfRy+v0eHr
0xIjbRhq0vQ64ZdgqNhyyM31gz0fxtF6FYzfU6o7G0sKaRdK5y9TeXQi6IwN5hPL
Q8dGnGZN7nVar3DxD1xGV3mz87npKeEJ5gH0dWGFMz+50mdo4lQeN4cetJ5hE2p3
z96k3IHupYhCXLyuDxiWspWMiKsrSJ3DlKebXy4ziczzDfK91ynMe9Ei9XBCOFqo
aUKtYF8Oi9o5cWUS+vCO+HY4OIOsiBnx6HMpkxmbllVHLEyrtI+R/r4L9TwVt7+t
xJ+/dUqZUjKWqPSSPQCSzw==
`protect END_PROTECTED
