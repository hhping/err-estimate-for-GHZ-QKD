`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zH97vmCGGY5IPo7/kRzBcu6zMR49yGY8CDKhMkMAxPZBE9ierpt15y97K9hxP/8k
rVjp1VjkEN4dvvE7P//7sMbc+KFUsbA3mvoRd95BJ31i7UNg/Dptw7rcMESpc+re
ewICmgiOP1qz88EKfcijgDANe3uDDLVwFvtassgs+VKB7906MopvuZYT/p5t+fnw
SBbeDmuYw0Of4Y3rx3IJOxuvFbQO5ArnFqp76h5USCAy42c9A+Thj27Fk9378mh8
B2Fxdmdon5ysBAr+4rdg9EhSelUYHZFwktMNfH2RGtB9absmkVqoSTXa3xEQTKSB
ehGjnXQn5i/7Bsvd2PeHGfCA03IjHUiguyCXaFGOHNeVVNnGKx3Kx258SK8r0phj
dDiuf1j7SaRun0T/ailB/f21uxMiHLzfdCHZmIXhZD9KS8Mvr7KohaRJ7vM1w6hq
CWe5XQN9uvEU/bCiW894V3MXlfKmACPgNXz4CHqXWDIcTOFEU4QazdfzUgpMRmHz
cG1zN8LTVQfOVu09FLIPpuWjECEReX/GPcwpB9tzhpjhi/jRxANAP1q8lfSi0N3h
gwQpWDtB7k8SK261qZZS2JYcUVV3AMIRMbl1g04UAneM3cKIhbkhw0fUKlnZOZqh
ojZe3aYjcKoD38i5LETBFxre1+9HYINH+0Rvu1JqsHGqM9f6aGDbosFGetSBErW+
I39MAwfjHTjXQSGKqrYtqDbHCjE6SWEZEbu2vXi3/50Zqt652ABnpf2/eVC3u1c7
7cgixYuaEGNPPAggpB2wAWjgyKIqZKRb0Wi2zrr8zrVHKb9puCHFBw0x8ZcUCSNx
GniaAcXSN8v4ih9N3+mHzgJznAPInj2advgv00KJCMFxnK2/TmDMjrMOvQQRNeRt
eKM5MjuJLdiyIg2SIQjAnWK0I79D10qiprdzsoNtIBPVVb+HC0geumG4zhnycb2U
1UZSTfByx9Vi+07TOl2sS7H07HIR3SD2t/vWLccLovOuhBjzMF7YOatAFGzeNf1A
a1HFo7qL7dyePxcAQIYHhOXm0WDrTuIiVgTWEBgXOVvLKl6T3BGyCtw08NDP/xb6
1jV5ok4ySmPSDDgWKBBj9kQVvBE3iT/scp8IWM27YdEkvRecgLGypKv7D3YZ9diR
TIrAlCOWB6pbFrLgpj++ZByXY1i+zLv7i/hP2ubFe0f1A/aT3K/fW6tpuNkhrIvE
YzjTAnuVLq9XCfJHl+IEzFplHv3vj0t1eg70l4cBhfbWIyydkCM7eSuOO25MRHN0
/YqB8Jk9dYMFiRL4JQPiDg3Xu88Tq6JUcDxyOm3AgQWcjdLLY9nyOlGB9oLdadj+
FQgL6gDY+X2HbqT2ADXxM3124Ag6n7EDt+tUbpXp38l4G6pxmzCd7UFYZ72HvYv9
1nGVNtXQL5KlSHpaxwV3ODopr3EUEpDJ7xtf+XIbjT7dkmcvHKjVbjV8dccX6/0E
uatKiORGSiOB5kmVpewxcFW07dXAvVuDOyiNecVtUjokYhqiG+beTWJT//phPewX
1EDMtspCLeX0VjvE3b+0C9IjPCA/gtNWRV+b3bAfAB8ABAK6QPA9s0jK26mLwWYG
JwYp8AxS2TnB/1ks1roETCShOF+g0bnpqLNtnXNsFaWqABYbDy/NCVXQJDIIpix9
oFGL68FHTSvOZJM+4KCkatuuGgcUv7M2su0U29Vn29JMM7tupUxMl/02FmvkFCFR
0jPe1KrllRAbbWS8WeFszhadIgWgN5Jp23f63ofNFwzpP3A7y/N3CoFxFqY0Q7a0
bDpBpghGv0PgL7yVV7XYmFyuTXxzGHl/3xuJ5dLZwJ2ATBpiMdKfAAKKztzpXcU5
fI0wuYNZVGgaiVTyn5QxUp9su+72vg7Tp/xgmIHu7EDLWlD1/HL6eJZTeMSNU9eH
KWDfzUpJjwOVdauN9SfVqxcCt3xt+d1hOuDK5W2oTaCuIkuHxsum1y45mL/pcGqo
nNkZiDvNG/ZIMXD2N+aZaLxw9vGHAhHVqCMaINnlhEbXK9j1ySc7pJRj8uy0wN5F
aVti5A9L5lEevDIn7GbPWzY9//ZtdyFTb3+fw4N6oHNChbEoAPqmhaq/ZRAWHtwy
3FUDy/UGsVtecADyty6HKYzGCwO8tEPxoHjwgIy9bX9sfV+zRKaEX+8NYGbAQ+i4
sK/Jds8rxlDEc5ff876oBFgzUWYfvM89FwywBmwdgHgncPdxBhpc96Ca3074e5j7
vG2UOSGSERgYNMpXJwi/I2991XZ8ayOLVnFnH9o2K7ifQiLpCI6jUAvhH5ihBU4Y
9lno82tkqBtYuthlYRfLlVht8M7Nsp4nSXqDrc6hm3y0wskgLo1PeXalvEcskmvZ
t1JZuiiAD+f9M0uwE4z9raGYg6C6ukJHLMJLFwwwRc3ila1DRd40WrwbGBZ+cjGV
GEGs3Jud7zfTGPXWRYFeDUOU34Z9iJoSqiZCvPkqGIQbKbLYJrb3oje911hUxM2T
kmVoUITg7R/mwa/ZpeEm/VZKrI2Z7wnR09Szb1CRdPJvMsd0Ah0MjP9D26hVVDaL
Yw4H9GWofJ2obQ7vE8cy9ni4owJlLhUZDHuFEPfUSKCk1/UGfRnmWh1cqQK5PmsD
bwAXnK75h9mspVKPPTWAsnbwA29fYv4J6ZW3UZGcSbfROh+07joJ78l/x159qI/G
FFC5KiUse0r1hUXm4Aai0D2LktQDWMv7+k3GZi3d8fPerychhkTImr2DYtDVP83A
hLtthorIBTFX/ZETwgUahZfEjvwMmBc3G4IJz4Ra532IH+HVCaRJRPOQN6Bge6HJ
ELKZf+2SN+33Ww4ABFJG+JkwAS+5Of57yFW8lYv9mhaGELZ87ulpYRqoD57F+tdP
q68mdg9/m9BoGuXx36HGgenF/F5xPiTHv/T6cFUri/wMZsj5VkQ/W+m8IsN7vHPb
Sf/4wtAh8chNgbZNHmfTmX4bfHwWRuGoCS/a2ha3+1c2UqWDyCZOUWaVvMH3JAs7
PlFGfFsBB26DyAfeICJ0dxAkCgSiOXL3IWbUuPqmWM1fkEey1muJA2n9JBF8y2ys
Cpp4Az0wlId/90w6tUGyENtt51Y6eLW5wzvT2ooFct4KXX8rIEYP5QjImVrtcBs0
UmZwkSsFY04KqjmTVRtFOv4/Pkpy67Lz0DNmDmeORXUX+qckFm/E1DdiKUkqyUiq
gikRo5xj+WnQKOpW1gPALDjaa5Om8oJxpCApS0mwt6NDICw/ddNE4MYwxl0e/hSt
8O2bOB2kMY+5mBxHHMbL0OJCd247CV82SV6n08SkIuJ5mWkYpkV50YKGKW+Lu7By
so4/+8XrqX1xWP98Hb+/nhHKEMSqRCeiXVne2JXaDvDzqAS+B6JBeGjdLhPTPwAR
fZJBqhC2E+70r6hg+ot5zoMyNhU1rju0j3hF3LlMd7W7hK59p/7cO0nANnG+ST+T
Y8mJNgTvOy5Pjye7pPyI1ArFVdAelZjPfj6iucjOswzGSQB5BnMVuksrQRH5PiA7
pR0S8Fwpa0d8xOkKs2KUzpmPcfsS7g0wYbLTzxsh+i1cv23gNTnid5ujgR24ZYF5
n8jGlRTJPufcCEBdLyd4+wMZ6moK2wEpkZPT6aSvm4KyNWyyfv1zM7vZyUHzvX4D
ndIjaJhOIFtfpFsfusYQ7M3eKdAfUWyfNG6lNbOlFIY08BdEAAesaEc1pIQpQrEY
hDeuA6o+9lXR5nsIfxj20QzlEb+A09FWH8iGA2m6VALv7ooUSHDe7ieEkxLl1/ul
Ntlj4kDdjcm6DdihPo2O+eLOsFO6ONfU8OIRprqkKmRG00zBL3ChwJ4yr3EuYGtL
t9UOObdxx9CBRXQoXLDBqKE9TpAXoUKMGVq/enWNRx1UqUrehy9uRp/ZT9/RLcbz
meAEaj/RiWpT68qp5yFV3uALCm1mAscvWyYhWpwTeelJulQBr//l0SDTwbJstnPQ
RWW2uxhadfN58a7CjLmPI+xF68hI6/vw5cLLO3HGSU3r2Pko3J+m4fL8cSgpwOKw
KagjFLPwJPrh6seA/Ebalxs7OhCPimGTo/1SVHNJpybbzwQmS+oNRwT8SFBu5g4H
9n6ITr5Yem+kMp1YDeNQvuL4NTxjzsnJRr2fKPrKCkL2YH/Wjy6sZz9PRQz1fq0l
0+742bmk1iZQOQNxUtjKQOLMPaOuAGvvdvnoSF0E9KRWHnTtYsyGDQ4q0+IR+ncb
AUJwVy2T20X571DYtzeAhsXkcnmX6oKBaCcNdnU6xplDp1J/KCCDDh/l472ADhvc
GVF5N3qQNtnnKBximTBA8QJ69vkNM/4A8z0+NmN7qtmNMbxfF2thob9CzwK6gaY/
O3qoXLf/TrPHepLT+Gi+Evf+6+cV4FCHYygtx745JVaOLw660lGALSL4fv9V0rqS
9dESJZpJj7uyL9mM12SyCIDZOZ5gAhJuHtT2GQYj61QolRTMuF3MKnbRIPCzezjx
SheT2CX4WmJ2wY/UAzxwRIfKwj4pezObDTYB6+5fvaMm20Cso75/59itwXv5z4hh
6OL9eN3zNPXEJfkAIht+9y1UbKDHdUhLocrKEkHLsIbEDc99qhfHmwkUCebEepb5
OoxThC8+sHhxxHkgf6IqSK9KInSyZf72rmxN08fZ6xJxLk+0w+9saN4w1PtlfK65
fFzYHKIB6bNop2Vc5IcfPL+KSAqZiYRGymMzuuYFoS+Z/PXIxy2cAAqVsyF4vzAU
1HzUndikOZe7vLcTM9+no78h9QVsVBMxXjUIqcggG56UPooy5fEenklx/9G8r0+k
Gr/Hyfvepr4Br8v2QINfGYYzVZygDovs2uy3L2j2LBDGABXfCEeVn5Q996U9BhJb
c7XeF3rAqtww7cJnVEWVadyoWMEC1hIuuwrZwb0jkQHzFSOutPIDQpaBGdCgqZux
M8EJsuX5KwMPPpSjLIG1pm3Vwk4PYMjE6mykGJwVY7kzzITyrrmRrjIs4MLvkhCX
Gps+ZUTBnii1eJFR/H+v6qPdOZPXP1MKLGeKG4qDqwnMsse1xL4VykQy614Oms46
BH4Dm0HydZ0Bh8UTaqJeJxBVsmBIZFJ8VGpeb8UlGiqsEDT7nOyv0xsh7ASgV6QI
TdxUDlsgDUF68V7mXVicZ/F3nTcwdMW5jnsQ7cNhPPcRTs3A4ynWKNRY1qozQIma
GUyo5Ja8pYvaeZ+41NZwaAzyq1myx/ygeVsgJabK6/woEmXGVZtbqd8xFPSs7w0j
LLKl1bIediZYVCH1Kuq7WCr39aMcIYtsfJStT0ElG5wvScxHLZ/LwMQJeIxEfMKq
PcdzQvC/VgU2CUhJ765IEtRQeZxZHmYws7UcACZHR+dsBmsbsp3jczgQ/JpX5Xsh
KKe1FDWg4sjXgMNAT/IJL42WRhiDxbIa/wejKJbZ/pwP/RvfYTynQzhG7ry3jela
qR0kdrWZ+ITZN2BfBL/HsCTIrNacUdyXB5fX26xAT1WBZLBs2KrOiGDTHZeB7YDL
rp/Dk3AQKWMa15R4kBbpzwy6ryyRV4JHuRjinr9sLy8VF+zxj9JmxM8oYGUqLKg5
bbx4g5sAEJ5Hz1j09KEEnvtHwjEu8ZskaqugC0JwNSB3s+qMxxorIgp9+VmhZz4W
FXLfj2wChpTBVs11crvhrnr8WJt/SHZAR7/VcHPE5cdrbnN8APmB7PU/48lzwq6w
DkixmkT75foulfYSI+dkofqoUr0LU5prDRTR6b4Vo0fvgXhpwaDzTOCmreHMAdFk
61F6YhgsCDbD79JSiQYtbZ6V27i0RT3pvrec/eOf9/cZw2wSszSKtOVMGm7JqQwD
uA5ePLw2sO2dgd/DJQGrDoSTvE9jJ4tRX5ZsE7ooiwa/cXaEvYFHchazDd2Dq1Ld
hmbbQpqR90+LFDY93FtnR7gcoJrV+fwbJdHjPWNUieO1DNmz89VJdImOdmBy7iW0
nU6vjn3w2AtJ/bOAkSSp1bEHhiTFdSHmNNXVp9yC8eCWxRgyVl5Z8EVfuFA+OSUL
tiaLXBWVSjPtcLbVwaQnxGn1lcZRCuYVHykPcTZPKqjziKkgIAAKQwc/6bq9GOWZ
2bfihJKji3oXDrKf5MsxXf9ehTO/getBE6uBCWUkDoEvrSH6abP00XOO3NeD+BKc
OKmDNWd8kish8N450Z2hrGyYRQJWiFwwh0Bc+cuZ2YiHYzVgIYROuQ4gfXYHnQCA
ZEzphbo9Kdf1J4ZqPbq08YXGiXv7FDTE00VrvUc4Oz79CjAuY0vaxPIc4/bnG3u5
Xtb9VxDLoRiYrt2vH3RO5tVI1TchCAcKt0v2zLY81FaINPntkQDVhijpN0qUM4c2
CmFD/0pDJVV9e7Xw6f1neQ2emigty5j5BWoCa5dkTdfzbZQZ3D3Fr4IklGniPWpJ
53EpjXhdX1K8CeH1TU0pNyf1+4j5DxePRrxxm6cJdlmfUFBEs4vFc0N53i+KT/02
KJeZfPXawbWO2lLFZpV86DqhJiBafRPPFZkbwo++kAn2rJbSPbZCLKURg9SFnYne
IRF5TcR+30AQwfxnD1mMFEORqGXtwHAoyCoWlLMDy2Dy14cAOkPvMxAvSqGqhjD6
8C5xqvQIcNi3QybgoVpU+spfAuvnYtGPS8UUUe3P2uWP0c1ftZpvTAt5An4qEvLm
70AcI92QlS7H58FdHuOaOXWiDl6YbTIeEiurF3o3qIyadLFTDexii8tDahRSAxwN
kkskJ90QRz3IgamB/8GB32xnmdxoFTsctTZwWZ8QEI3/ifUNY0WNSjIt4OwdNT1/
6wYlx/NQ6feAVRWeuwu5OZ2c5dJzfDgKag2Y/s6rkQkga1BwAqLehzuMIGTJqPXo
nTwjZjRB+JQcZphnFth8Pam2tDjbuE2ZWSptt8seCi/2WDpxG4grPC+RPtT/N25Z
9mDNwfpIdAR9nikJWUvFwXRS3YEBbnSOD74KZHb09MY3iTR8nb2h3SghcaCHAxjv
kmwl7ECJJYoOLcOZCq1fgjcISD8hJJEIqBTeeghQ6QXICvMHLph5yUI49a8f97DB
nNOZuUAq0A/M3v6OLxG1AdA4aOvMb/7nPXsZKLfEry5F8yeonPnU6673OPzJb2N0
SmALpglQKj9gVh10PP4XNMKoFdHEfA00xe0/exltEbWzg+2nt76aF+uPO3aHCZ5g
zfk6In6/y22/ooG5GqTpdKEI+WnBGTQI4EWL1mWE3I3vnTsHLLUKuh6ZyQdd2IbC
Q3hDeLYGHdWd+ALu4RLcYxqqRQ4WXAsLITQ8TvIIQ9r/kPXF4EaZ+994VTFu9h+9
ySSCtk/+gxBH/Fp1/qObfRq09NVs3nJTB9dMCQ6dKHEfLHR1g4ezZczH9EZXwnQS
NeEolg7bMytZ56gvoj916ZNwC8XTvQtP478lTvSu8HNJXUZ4J7PXP+H3cV5tibLU
ke3IeKU/Feznm26uX6JIwALbj3b6rPFV/DzAICzja1AP/xYziiCQqvae+AiFAfi4
J9LnF1jQkKpSKOfTFgKKJt+jWZI0xzHKzgUarCajSasRnNalZv6CcnOKovXgaXco
AFLBpAZ4du1lZiiEtRhv/RMZD6Ql1IPnTkCV/tAjaaZh6PWdezu1Qgd6Y2Dcmsj2
26BkpGrewqLtuEzw72xi+3xztQSVoYE5RB0BCNZMUKoIYFd61c+Tr90N1Sj4dPna
UTLmedQfk5hrCMq9HjG3Iv9gHL4JyKX06gloqZNFoO2WEhhYSQR2WcPu+p6DmmHi
AvbD8fpFwA7elXg8IrIetD0RLWUM4HBBQ4B9uxk1hDW/wLhlyZFyVabx/27V6dJ7
PeONlDn+HhzIXI28Ed0bgw9EqovPc01tNzORg4GxbJMUQth+/YMfOqJ0JDq8KPTe
MJZAOrjmfkj0QDW0FrpOaJGJ9kwBx9ixUM7lF1HmkchPl8N23IXqF4lKPG1zJihJ
USAbEN7SCgMyaXYHiA5vunjJHf2gqhNslIAWEfyEvVIpcvy8fZTq1q/pgklvFjps
WksJr0eNBM+0+N0WqwUvlBNdI/aaq0ysbfQclq0dCq9Qij/u10BoNfQEi30magu7
jgiX7NRltXjNQn5JIEkr4HBSOHve81lDL6JZtKAJBunmwTGGHQPKMXP+FxHywycG
ZAoNmKkfzlDt8hAerzWa3QSpvqFZoOFCiDOiANhRX7jbaSlOb2/vkehb9Hk431L3
8oD/QftD5bQbLu+E2lDhrnr7pIXjHg3sEsvevYj9Q4HXvwxMQaX7eBRF4HhHF54o
vYdulh10bYPEkoqXnxqPXXzSIJQJjlMLygG6NEFnbmY14PK5YnKVFfcGAjL4XIHS
oRU+lBp1QavqnfaNLtAipQF12bsNIeeXhHSjehVYD9+1/vJfLz2fnRqEbgOBSuzQ
o34irg5GJh7iKOWx2Sae6Ws4wWZw0+L8Lojo7dygRmmPlLvpa/yXqt1iDKkDEIaU
Q+Qt05yOtlG/ErQYhy//c6sAeN2uJ8Ap9MIMNf4qHvb3nffr6Q8T2mvbu+4qs7Q+
qEWUdrlE1xBf0eFkk1roJFH84zrT+4elpsukbOTS8FCVt6u44wI8boVGSqu5uf/D
F4VuJKIIJt3rUyW0WtDp7UepILE6hhjwONhitTTGwAmIp/7OBUaLW7RF8XgzBI/u
E/095Lzd1HYhtnT+g2Iir4iCL2QNdVeSyzLWDADre4Akzt/iPtnJyWNdOqG4p7R8
WePn593/H98udoaLNUH2Vm1+amQqfXY+vyZvelHpxWAIbmL6t5R2CgGfQ98gtLsf
VbNBIgkwjD4iS9Pftoh60hbAYAim9HxJO3enu2PGnO5Xlvo1E9TCV8dfS4ozrLC2
3yf9+Z7Ddg1d/W3+y+mBVXvtUPB4ysbyKE4e9xiu5Yq9udniMXcXBu4EH2ia2yQl
u8vty0UIw9ZF03obdMRMOAAFQSS1ypJLh1uG4VmtdDcs51rO6QQ+PEKLBxI0g09E
49Yz5WgnZ2aagSL4vPbcvVv7mbHtu/Hg0OZyjUad3YKCkFrrtzwQi3pRwp6VLJcW
W+mXCuVmpIDNpQImsdALV1UMe2tRFkubrk+Ht2b8nW8uioagniiRi3lIHz+3edMZ
6h7uOYPYvzN9v/HbDiK6GMegQxOkyP+JQKP24JcWHoxGqya14Fb0es4V5k80xOV3
dg+HpStzxT905kVhrfBHNAcD/wJbOOkjJit94bIur6T0nwRV2/sMR8GmnBoh+BJy
2ajqnVeUMVhvn6n+OvyktQT5zm/4v8EoaUN8yxD4WBseOs15glh5+OwVfOrKjXQz
chqHodW/i1G/OUG8ovBwrCf5YTKO0GclesSa69QVHrMob1EzAIKEwX/sNZPmSaB5
FTtjw5TYBUkR9gDnn5rwb4/E1DgBXY4y0HInnAM5TBNUMkcGSqchQTRwgThgy7Kp
R125vgAo2qong3X8MCle0JuihqshWPX+xRpKlraJ9iHntcfZqRnVZ76YYUzoQl6M
aDLV3qaXnx73q2kUAvpcxkQZzk/g7A0Csx4xCofiz1VmrVpvs77hQsNaJeRXERXw
JGRJnUG4iDoEwcry+OARiWbRinKt/FEIx7Xcs+EixEsEC9jZq16mEW+P3n/eh6jS
0hzFiQT3jZ37K+rSIU7j59JIc96kptfEraywomczgJLFdqMVXyUyi/FZG3E9E2UK
UjF1jmsTq6T/tIO+TC5yAIV/MSSG8p80STP/gniaB36QR14oEr/QPsTgW6PqXqM5
Lfm+BkZzmmsYWVQlNp46FqvGS+ghhNo7M5zNlOPf7/AO8+OAqYdyRApGPoRzy84z
ZDQP2S7p+CTaNfbYnxMB+IakX7DZ4hICvGUQi6ui+IGw1mHEHlFZZeuQNOr8taVE
p09f42ouzWa89ztx/NFNRV+J7udQH6KhhIqNnTS58Z13kLwiJXLKTKBU5pfIdmF9
qQpqhXqxS7aDBuA+2AJGvqKd/t0Bje8EV/JZRn4pbN7txi71qLZXDslPo9Q9zWlT
PcA9XHfoYjjnab2wun+yT+xBGppn1fpXEkU2HgzSEdImI3vsT/7K8tg3W6N5B93n
xwmxa+rBaRhb8VG1ia29KM4WRUTDF2HL/dpPCJDgIaz6v3JSKtsvj8vkjolZD6sc
xROT/Eh8O2g9TtD2RsaGZkTo+PIU5MUJQcCwo2JdsQlelZYNKQGBZ8Mn4Lb57l64
DYiZbdf4h91QiNsn0M8dTrITHGzUjX0RCoYSbfShmrq98YlwnUhx+i3HWvvGGLxE
yp9FNbxjz1lZPlKl4TZLr879c8YNbT8k3DvzY3NYQ+aLnexjXOgOku1p2/6dzApI
KAwRikyWpMdh3HsosN1cue/jcUsQIT+A89zXj2l5zpFlxwdtSQ6AM96T1SKsueq3
jf2mMhP6ptNt9XnlGelODSYTbcSE53/3UU9KshhOQGiHRXJj4dxu3z6ZpMBypavo
lfgOLrrYyW3KtTyNoBM1qnrybBtq7dJtjbLBOYH7LnkDh+RmPFi+qJKgjao/VBaX
h/0Z4c7nJxaWpHq+iVpddZ1nuWuJV3Bj5Fh713dopreojhdqMNN4ocYkDjTIwRkC
SZrHMc6wV26VISrlqCiE9w3WWmsXeujtGzlE6YS95OD4UPb5F/DtqE2926zS/yYK
yR3d5Zx0Ui+WA/CHI9VXK6VkNH9UiGnaAsDBRPioQZBq/TYB/5gj1+SYLftDYj8f
/rMI/zf4+/I9MBDMOMFa47z+FPDHAHOLSzvPZi4JX+TPPeZwzRvoLxr48fSSYow0
eWm1VXiGUTXqXW7SEmRiN97Iq+YRl7Wktg/tCI9nbDTABLym46symPFlQJ0weoYQ
iMCpaPasGd5uO20suRamQYBNUmtGH/zVB1egErvAn1UlnkW7dUWW8H5YFvM7bvW5
LzDbCHW2H76J2q7asJSlckgqMeKReuvx53X82rd4Fdd+meV3r0VK4QeH5WRXqJ0J
VfXYPZxJwzKR++OczEMz9XYMtWZPTQlTZhqTfBbd/iTYTgZD7L4p9S47vti4pMQa
wjwjuukokcZNs6fX7DxdrxfLf2J8PHl/xk8ZkKzgI7wcy4vtRpUlRzAjycLmEd9k
7jxlM+IY35O8Na+evzVUWxcP5uaWSrrVtp2G7Ye8c12tu2NK2KWfhn76fFzghszC
1r35VoL+ou40kVLhCv4TGMnvS/0qhYG8vRy3W6ViNUZfAy4JESrxtuKAr636qwFf
0mqtPVQfZSReIJ6A9hR6amo96L2LZLIn6Es9eVBSrCVKEOzYRTy4bVB4xqdQA88X
eCI18CEN4CmxLc8xSqO5NBYkaRjfEfj0m7eaouFpPQIQ5AiDgb0M3DsLIhzKqQCc
H7Lin+lszB2bHkbVsvGOfjLpEtVY0qyCVpZKMX2ZwstOq26o07ASYbYvpjHyrXuG
e+im26HO/Meeaf4noHqfGrSwGk9DM8er/y9mOxsHJYUoAuDSo5TpL334UO/bIH/u
bac7SnrzkbWU9frnwCUXTy1lv1V/RvV5Fnhcmfr6I7ETpPcV7MbXU+f5cci6dek5
Yw/wcinq9Xr+CK8mXeSqQ2Ml9dTMHRdvknZOrnYRqoFyaSsAEQNkVOn/vBHlKFXS
ZdlO8pFgYDF+eTf5gapCnUJ4FC0HHUZsBaQ4Xpmy7ERWWv18LoO1F86CIz6zHgPW
upzjMQdmo0wWjBsnm8m4pW7cBqWSyXsTuM4mIjC4A6bUCMprf6ONuZwSVcq9sEdt
R3ondXBs0xZzseYC9exEjVsMqbWSH+etPy3QqY9Q+XcVKdq84eQMYoJIsGmC3ifq
njwbnNpRR5Yw7tab/vouSUqZP0a0jJWyk2Xlu9qNwMoQLZTmB0pqTafDZPPLfxZS
Els2Hpi3R0Ym1CnSS9yiyg8n6+ASQMj9ssjW0FI76s5ki7elzygvmNC3K7GnP6Gx
LbvxrjoYEatViSIRoZrs4E2WSOCdjeoZXK5VaY4go22GnORh6PZOf0VwMKTJ8ulm
MyiHuak5fjDub5Z4LLkW87OCPA2JKR9CTK2zwO05NDx435erPTDWE7olOZA4ZXCA
vNa3QWIJXBSiqGcF3yVEux2lfxeOlulE7OWlsccmwmwYVPFIKBiTWfgXTJrWnSAs
YXKuvYBrUEnlP80z8qbJBZDV4hQAbQMMeuPysZRJHQ5caNGKUjou9RnnxtRYJwbB
ggaWVexMq7R8cj3ffcKvjbYe4VhFW/MwNr2F6Ox2/Y6DtcQyV35lzeMDuyFNofCA
pmJNQXYjADk+/huTMJFxmsDwX4omo3ntTTm7ChN2lWDbixs/F24dcBgPBZ0xt9kj
FkMVWCjsdxiW5Tf7OkmPCDLpIlL/+Y5BUVG2pfrfO+l+AFEhG4CLssy71RFrpH2R
6F3Le/XmDsuC5EiWdNrUEx9Q0pHhjwGznsbffelocXmdmOhPCyRzuaPkndEV9kmK
lLuvFdyQ1JjcXpSF+lYVz955myP0ecp1fUxwHWR9yaKDDAwXG084hv/DBnVuw8tE
EaOnAzBARnZ40VfWimRSvz4OLraDFPRmCGit6q1ZAYAmjwQSTWLMZ6kuydw7FYjZ
39SsiU/irInu4Qo7XzMcRX7gNNnNQ90fkLZ78ILWoJuZqJmZhqRKw6dZqetWvb60
pHfYh82jeVL/JOnD/7wxwiYmN7XkwF8Lt+SBmFpmfcFJ4eIvcNvH3luTrt+gIIQB
xG0HYEujUDEyMQqxGrCQjxXuNqBxCKRBKbxiw9UnGKzlbQj/JRbxWwPh4s7ePUjx
kLA0uMG6AEyblpu7fJeeWdFUV2CaYAV2s9J3ccMkFzm8Ct9forpwv/Xcqtt5QMIb
RexzVsBGvhQz4XBfI216ViHNqJPXzTD7aL/7SIwl3kHgPDr3VBctDxxwZ1hiUwoU
fEJs/KNOztCluhDJGCmZCh5K31GCszITGmB5nGRoPju5KnorY2L2lNtzWFNbTHJF
BRSDeip/fF4gMkrFCo27Zqq5Qk3IWb7DWbr6/wwGHPTVTj1EVNzLaTUg9IInDM7k
vfoCDrfO8neW2BZP35Ix8g+hm+b978Pvjkrsh40N4R59w8vYb3BPcsebfgJpbOJd
QdJAjK2nrXpzzAXeIU86HUYbqp8usN12Vdu+7ju+F+TcwHlWvPc0KpVvV1BXwJn+
bjNJgOozJyEbidjX2lT3SZhlMeEi0V+sz5UAkPpDxEoX7Y7WmhyciihacNgw4C/b
ksAxd8oIojAePLUiGwT52PRxvq+1cdjxcJL3a20uALB8WRbSMzIt1RgBcNL1//ZG
jfB5HKame7NeMuqlf2HOn2SXFSr4yRyi80snV+TcXqQM2tc+5VQ4RGUkeDjVXTPw
to7olIiIMcsO4Fy3zbDXAdsFsy46oQeVLAPKOmFz4De2k6kzlFWJtcQW0Ayr03Kn
TeCQGtXl2ihivSg5o5ocggPtE0bDJE47MMJnh+Ww67hafhj2Q3bakjJmg2acTPQh
hJP7bvjFeOivGZrg8+7iCa6kHQxQlYHeqtwNeiIgpOy+lJQL2t+z7heEN8l3LMqJ
bEumBhJM3OtGcf0Dn0+Rx4N11eGZBHr2Akp4X0CCyz49o/wZ0rJiiHrlHEX49ASQ
VT+8kgpr+lcL1k7YfW+oR5GnoUDCo0ZcW5z0o/31taFoQQ8lW+kmmGKQQ+oxwf18
QiROp0U1299aZW3Hku06vi4M4EEt4eLESgcP9/Ua6QZIx8NcfeTImaswtvQgRB9C
N5E4vXaABE8vwxwtmxFouI8oY0XvfwUkQy+CafSceqYMqD4kO9OUc8/qchb4gnVh
i0DmS+sUx9Y4hh7mxTXUp8sCiAyFTuSL3ZhI+BRteTmurao3hPGqfmNi/KOI9sGq
XPaqATnJtPFfdpcFSjKWcYYQGqEXvzlkWzOTWXp2MUCNtj7zBOCb0qst4BzJvN+Q
YEf76VRdcdOTyjYLQqTJqgZ3WKgr1rOkfgZ4Tu3va2lf9bbUVZKqjWw+W6M4VdNo
Qs9EYSQxS6kgkgBYhZtAOwz9nuvzCWddzd60Azzqqvy71xS9bmQUB0dvlvca9C+u
H/2drmes31T/2YEyHvAwXuMjs5Jzw8tbd5dzG/CJZZsvgBXOLCvuMpyQXhjgoMrS
KUr92Iqoy/7jiIjShd73rp+7KGG8QYfdqFV2iHD48RnCcIV0PCuhaUoxO1cJAiBe
1tzCxMbO7xuCjrj9uj9gnOhkMCHcTF27VaGPTQ3x49lafPxDqD4M1lkvgncy6Bag
GdtrykMqqTCOtF9gm0dG2PiWc4ZEHB09EzJOhiDaLCf17ptUSOXFi4JSomvFD7Ud
8Zx9n4YNrT4Tm3hNOPPHMc7eXPLYra2qF0mXbefP+9wRChhqysVTHNR1EI4mY9tF
NLxfOne+6dBfZobNotNju0or18fJopiOkH3zF0qLniN0lWEBXpQLjlE1nWLPr3+o
wcjiejF9NXbkcSCH2i6GdsW5gzi0xBvXU//rF/sHfWVycsL4MDeF8c8EUHT+vMwb
hd9175fjTePlQ8K8RLkgPiXwc+0B2JjYJplmpqGkpc9fXRRhlagc42a3AJZ1a3hT
9gsPI0UZAGaXcrB0F6KqmqXZUEeCKdG+HRC3SFDJWEm3t9ilAs1uGsnVJulpL2Xj
YZoP+tuhsKm+XADmYm+ekp1Zwoc085ucFuBA0rqVHOlIwdg6gA8Z9fzE3RgO+IX3
07E4Lgo2xVtY7E3E5Ud+OuAoTKaSYv5UbsQ6ZkdAc8yPdrR6lXMX62w5JO184hqM
D8JA9mdLfdDZxGpW9/6cXGLYezgf/1yeQS1C9PaXD2GEDIYBVr3GY7HqvpWZpnXV
EKHomtCpU44sg+O/zRsSJdcHwnLNxMGzsZnEVYl/aDrHooT84Br+7E1afMFKz4oJ
7JBOBgjxNGvbO1lIaVT/xBc388Xahku/UU+Pbahuj5frpn5qDJZFwoMja3XMNgYl
05f8FS0FyT5nVzJe+1VVSK3VXD9OF+ats9a9smVyX2SGzdxmdhr7BixP/OTWh8V8
JbH55OxBuDA2qsGhwvAcYH2YeAQ9Izfp3J8SlnJPA81W5D4yAHhmrwD2ZEh8sEL4
+ty2rmr8Ay/1tCB6lXLvzEy1SdXMwiIP+5Wugi2vnvTVK7UsqHA07lzgU4cEyDsY
+aVlrEM7C1wzTImmuqINE1/EwP0rbgtMSSBVfmvLG3x+80M8F3jnV5Cxh9LzQk+V
Ce7RrcqB/btn9V7bBBxYHjn0Bw1Vic2ayxdpgiLmfYWW8oGbL+U5BYj2+L4VFKaz
ra3dyilPo80Q2lwz5U80Oo/Zk4opOMITY8UH00QFXbYL1pnOM0ydN1Soy62FSxoF
nPx24vKjXLKwtOOa6Z/FeheqyS1PClS2qPmXAfUfPsgyyMAEcCS+1mq28dHQZh9q
2We7U8q4HlXOnUBNOwOmXNGmNIEoSdJdtH7z/nQ24JYfLHqfCRQar70alkZ5v1BB
2wwgysaYdiOHxWyvs8152o0d4GgBpSyBot9XVYy18JqVK/82N1wwnHjEJbsDXqlm
8rE36/gTt0fqWo8fmCv5SQLn7Yu4gkdfjtu1Vwh938LjtPpcQgCh0AVX5fsD5eDt
8Ss/CEUFbQWnhTJDJztM7Pb/d0n7RM+vsym83wVQajNALRiBi2WIVjKdaA/OyGti
drjc8l3gz49L343cRY3bLTLV93AqVaJAWzZKsVs3VbnuENANhSDicOrvWZJo1O+K
WyxzMWMd+u2cxJNYhVpTE6HiUpUWEkWmyxTHN1XCLlKRc5a74+phuB1XGbNectXb
B5GhqYGajMWHBynWyzSsMR2+YjEWXHdODtsN9Zb+bRpvbbbSxU6L90sFLo4JD1aB
LDfrDRjnDUIGMM9fGmCxM7J4eyP9RZHIIY3xcTZ7xOUyqOSedXZCfkDvLQG4esGQ
33ehBJiV4uqLyD7TcTyCM0i1ixrdWXypKqqUH/j0gJ9/bp9EcFDSXgFR3083YYZs
e+Da85tcLtn4yZcFv4uA4b1EN+NUENAYFyxm4L8r1wImXj0MbuUuCa7bZP1nv5UN
bURXnzPUbswGODtN9X0awxCEiENVWQi7AHM7IlCmIV0VDWQRJO1OlqJE1bL0eUST
Vd8HzzMm3YzrW6Bg60XNSag0Lo15DBCtUva4N/4NcKO09L1snzi9kDgMYaQZ3oz9
+KTj4TllZu45FIPQnklk9pSJjuimruEOT0RLfnv/mJGWq/NjjzMSW9ipKPuzrXU+
6pB+n02UwGqUlu3XB/ncvG+SXVAV4R9Pp/eq9AZfsx7vHNeyqPJRt90uV7yqdLAN
OM1/kFN9+IaSNn20zl1FPcuTMibZzkNN0ZzcYQHUh0uBZyegdQemiVgBJbyRGKlt
+Xd1opTi9VFZ9wPQkM7qpi5anE9mbJtq0adNn4RfU2AEVyHJ0aNbCOWIuZuWqCQ9
9AEKKwTNamZgd1MgJ6hvN17HxhhUfljgN60kNLhtSqy6/r5f7/L5cbc/KbyEPN+9
31vXBFtTJRt00Uj8CrY3PQFUQ+Rn6om59HxvlwMONdR/VF/5KSsAtpnJHsZc6+IK
/B4Rp8BJzgG3uGllFLR6F/xJjNIGPyUPirjvFT9mBgv1AcR2g8WBXrylpGcPX/d5
2XsAxW5qghC5fQwnamZl86V1Hk38v7mOxL8sBEx/CFbfQgk/6Mp0o0X8jdrQuFRG
4UG63ixEDhbR6C9uY1dMxVNXDhi+Bis7AtL/iZuXub0/Y3DYge/P+3rhgBz4StWe
n2rrOL6jrKWLLqV+yEQJ3HMtzJYHtGaatQ/qd3C9T2q/2OzPQG/6r0KTsY8UDZKT
kzGK/kqySp7ZOrAD9E4i0qi/mmjRO6upnH4jqDEQiHlH5vSgyPdwyV5z5/GGoG/R
J7CIS3M9TnGljoaEutANKTGEC1WBxqMW1YiJdV31UMBWoY5/zK6/Qf9QH44R4a4Y
2hoSgs1I+W1S084Kl8mZlXMKtEHVDXgXc9MC6WC8egbiliHXxhcYvuupF2KyJwdb
izhFjbG+P/0Ls7dE1cVlPhoBep4lmX2H+vqV2ZgutYhaZZ5FGAFRwRGJk5w8WuvT
jHc+HAs5wNYYNh86Mkw3O1/Vh2ozh8E+gMgfXwGxetSARFJfZNaJ1qzLls9J12Iq
As26V3Dbj268AbntmQCwfqSGuQiqpMw6x+xjF3fDthEd419nPuEIHkCynQy13Y76
aIgr9KOHTgGq+WK+tS47W487MxZ28VaMSr61Q+Zrutkz1fi1g1IZdFRE95/Goe5z
gMAmXg+XgegLcVLmYsvmmhvThaVm8nNIMZNYbxkERFnoTuzztV/ilihJzhpm92QK
/Cw8OzXVBoqersLBD+PvpmE+80ADFABwRr+pZXt/5WFzcKuobNlzE2+O7bWaPprB
5NYNfp9zz7Eq+TInINpEMhBhDprtjbi7exaTTaXMjQwrC7QqQIzqVlrQxlH3GAxX
pZRdkcgIC5d/lft8Eg0AgX0vesYtt/n9I+vMBQdydbA+aKn6QuB9SfFovZJbSoD0
K3LcsRqqnfMKcshs0KpPbnI7O5Pc+GXPmUawLnblbvqf70puXHfUnNegI07ILSqf
9JLvjxoaDmKDrgnVU6RLHfv2+tTwts5ZUlMHVI7yFGYCol9clEJjSjRAZUoeFTCl
55x3bGSdWDuoXtjdqqsBi80rnftRSlVpqDGSAHKakReSGe/12Pq0AmvlkjjvSY0T
m1sK/FMNadyoBJ8nrZyvjslWsaiBWte1w2WV9xENTPq8wnEj1sTOwZzXFuSFJEju
oqqEtAYCNfWPNidYvSjmTrhw7z6/mIAgs9s36UAxYrsdozfNVJZb/9N4L7TyVgOj
DT9t3dpHckUsAWR6tCNjTh2SjeveAw5DYS5O4++I7Fy/AYguk6k/BtcX2u4cjVul
a8Spm3eM2ndvq3jH0ekHGkdRSm+hVASAP4jb52qxGcEUMCLH/d6HReyCIf1OgmES
0d6GCP9KTZrGTZNNoy24EeKYELA82pkBUpysG3dyU2XO27Rb/QNwwCEGkaZPtDJU
EdTwpW34h4ehibsI0OFcaszWtPN1+W8iGPAtH0+qeVNJQRtk64aypDjSWs5mTfY4
yEEwVRGr3VudPjg7kMBXz2qSLoQ/6AObGeD2gqTDQIxdQffF2+0FQjYHuGcAO089
CM09wehPrZZDwEOU7P48Ys47sYLS2Cp2OhGpZG7qfxtRB5ukBYQNuA1JTQxkGQgY
Tj0GpIZoFDgTro30YaV74z0IgiDz5utnawImcnX91vSbrE7pzEeiGcmA4eu5nqp7
0zFa74I4r+55Axs/2xF3JflEF9WvyNvCWxCFKjBnT09Z61e0WhDAb129JEBxtF17
ImXLquKSzjhhByjttI5ZbtjG2eyvsSIgoR+cbgDUPQrQ1cS+ZvYDevlnRvfIM6oR
3p86xhmwiT+EN6h41CGlnLOlnUbtvfW6KIDN+S3QGCr98rhyf8PUWG2CkfK39FIZ
kw6uAFGTBn5g2K5KbRCOoPIXKKMfOKe1w+FBafLt/7OdYK1N3m88GpDgPujJE5sR
kP6SPBRbZee5QMvsU2TgmnTQsRDBmifef3q032FCIx9hXYJVi2KjMqccemQ7K1fe
uSUXTtagtKB73Jnc640d3eicNEMEik2qZEIiOqaVa/5KSX8+2VAwtxYSVhBXibRt
JWc9IpL51d/rGScDguzok6gTQF/jcY8FuF19zyJwcwsiT3n6qTkqGcRGp2Gt0QL8
cmuO1cV5of4H6cKZkf3pQWx81kOy0scYVUteDgcHi56gCzAlw7LPt/BtoX3OdOnB
cgIG9SD1IY9MJyoRFCHdG08ZoCC0FytGkH8Ep4BeavMHdn9vONLHgD1Q8npOr/jd
c0fFs06oZDV1vrciH0KslGtPbG+9DExYIvjrcLeU8fpSXsL0Jl04zGHx7+lBnOIO
5qzZBSXgMYulXv27SjiyAVXJ4DxCUSrIsMNHdHqrp+F1MQpVfstZNE+DdzyedYyr
zRuQ8ybPJQUD0RnwSlQU8PsJ7gtzgm08Tju1uChV75nLLElXIrueruhqlW3lrCBi
08krXywdtpKhJiZiWcx02Z16g1KK/1eY+6b2gxV0vQWa0ikQzW+DfmQ/HK8pj8uu
EHFOoPev4YzSyZYRNOJE+UuoDALax67LKRKDrztP7qgWYgB4HgRUSaNWc2zrk1nB
TDG0rVFQgoJP3sTLX+DVEg98keVYX7+J+6XPNu2jOdqLx9oG9BR4KpgCfRf9DkXt
VuRDX8OGOAhp345j+bEqpbPzhWWmipN2rYLZ+W8udN7xQbfjHjYB/llDi1HLv3/D
4CZLbMJ7btzwaeabOXOxFHwRDI2fRLNvI5QcP5USX/UgGBiZJCuRwklDJw2IZwP3
LaE62r+bwGXUbCDX/Eg+sfh1Blh7FcyHDe1mEuHM/IEw/OdoICp8hUE3pzwirdwZ
KtTTv7y429C9uqVinQd98Am6nwasObm7NjjSev24xujbHv3263D81HEUm6IuZiyg
APJw9GZ8c5pHej9F7hn1U1J0ArkcNHGUpxRSx5kRdlIkAoxEKgLhYlD0DL/kyEB1
wmJaG5JmLRjbsGRSc64f7LFBAxH1tJTbxSrvoXnpikG4y5GZDkAeNAWO8ROKYzGX
hDjZ9FiwUbSI01CNAotRElftZosuko5NO6vAyCNgzZBOACxLrQzeCPpDJZwRqYaR
7JwOA5/OD3OdlpdDQrkldFDah0tB5/Pm8p9Kiu2Q9/OmQkDxB4a3LbNg05xUlHSt
N28dSZRrggZnA/eTPHm6XcnSvsBHPLliyFWBcn/Lpt/1dT8WULkQfSzE9WSX7PU2
w6sB0a0GRX224nxdPM+YbJd0+uBFJCSnFIzvXg9EpSJDwpXGeP50jE/e7bLZo3Rq
PjcqDW/FErPCQvkdVCE3wA67AULZMBrCi5/CYAbaI0Q/SoHyLsJaNmswot1fBKBi
bJuVVU4fEvXWnDFQjIf0Xj/YOdmA8Z45Lz2Ix3S9bGioYvMnO4AG8wxHJe2czHmf
GAGKjKsqMHpNg42vgHAHCTesCKY5Q9xdESDjAJyUzHCmvXgc3bdNpRpYEYMU6nGR
Xlrt34xeyg9vqjgQXAkm4OSRPhUk5+1MYAvAcLIDcoByCBIcpFPNZqKIGyfAz5oQ
2jNTyP4G+FCWoCzS9R6bHvF0cfCl58mJgOl6ACq5+Ve4N7Jvp+nf/kBZTCz7GgWW
mRrXK7HVbdlxOBe/BzzbUW/BeA4Zfe4S5E2qqkHU/ug/OFBHKgaFSpfaJnRbVEKO
2SLbT/cyDu/3debA2eQhydksoqdHJ6Wk1YpSrlzuhVnCd9TYfQ+zbXefCW7DjvR6
STDfhfcHKC2QhQgw0wwJ9OgoiyYAu13raLeDVO/MUR5w/4UzTjOd8uuWs3JG68I3
zmq0uznrbnGRO2M8Nf+coqBNKIYJCOGknso/0EPDZutGOO8fwjpmqn42TKHQ61qA
RmNFBGqcMU5J+571mV8sc+a3TM9M5SWgNNkiFpKadvpqbHT9qR75G+aeDbZbcpSC
p2IHmRQVaNmOXNftKR+B3X6pHNw5jhexukb9cYcfFoPGlQSoYkngGbjmDW684iGp
B4OWqdj338SfjQmcZpSWdYLF7ZjJMeS3UfKRYcmO7J2QGikD3ciHJokrzNo6LtOC
lPanoN6RTCXGfF8I2/4E08oCE7ZgT1Ho4bCfSEoBRBtkVXe9S0YGRz+Wp/dE/15A
KlJA1nPlNMKfYMCKoqqJ3dP48NvxnpSHcBag40qfGPI71RO5G/WMOWPtzWLHRKUh
54RSp0PhyowFfWWk2cmdl4PXEJ/hEr8sa6spEoP4bPaSL6gMd6A0eX9nFsU5lma8
1fqLrE911By3iU1duae2SToaLyw3jVrUQoacAu0/VFdf6dxcqXPioO1nIKSTcU9y
EOoHLOTexZpbnVIFj5zyxLxUBz7KWSFS5WEKeFVlCHj1YbF+mRFTmORiaJegNAWT
juvV7iS0LFY8Q/RyufF2bh5aej+zw7n1X5m4yfBZLjMBILOTSXi7YDgtv1QWSlvk
6wDYoRGQ60+Amw6i1j27eVck1+IUu99kKOyusBLNnfaNoY2Wv8Sof5wtdMy1QXRJ
WxMQAk7vZrE9vb14HS7MIL/hNTUsFDrUf7XAUGUlQs1TqUK1J1D5WB4YMhXweBkm
yjpKG77cTc5vs/9BCouPN26pfZONRik6D7+pUw3WMtyvW2ojHg6hpnlfVmriysMq
AWRBGZsLZpVu6oHqIpSTGMlbVQrappXksJy4RcafizdLCzAfDo7R3HVRAg6XSp/M
QWj07o0c/7zXoNFFroFSyvGWmaOU0gR2M6/lDibuYwLhnLRv2vZQGoQd9D2IQqKr
DYpyTEXvDzL+RhECv+diqPP9HGnfka9Yzqhe2WTKzxkSR89kTSy8+c7WH+BYSwnC
7RRPKM07DRxl6dGI/ii9CgLf0Zbl2fG7pn+8Y3NTa8eGm0ObihgfUhCEVWNRqCFk
NeRo1y5P2a1MgoSVjIm3gyIuODoivmjBzfhmS9kCqgAUSP60Oj2kb6/f13BBmdGz
tIfvLN3SU1xxB/sKNQyEcO/Su+bkfYJNvg9B4WUzCf/gz/mW13+6hINRceSqv6oc
06TO1gJZrsxRU/l7p+/wjTe4ibrcUI+54/U2GJLKN1e4J7QsYmujO5NeJufl84ii
I7MbXQWgkzxgGsYN2N0ybnpGUXvN6PhVeZaG+c+W2v81fja9IazKDIKcWzftk2j4
RcMEgggO6KDol2wGauAJVHXtdKogWvvpl9jWIEg+GGXVvbbbmzCCQ5R0ola5+xo6
Mf5o/Gyj9VU94CV19eruWajLnREf8FWbxXM8T/oNPRid0yGXj9Rv2R2aBSQKcd02
cHIH+qln7dxOfp9RjMS6b2ehsB104whaRNHySRbzQSdQA+UrXk0IGI3slbzMPREf
Xn4vL1FfIUedlEh8GdUvhSE3wxoCdDKstX+wqWaSu+cuDrA0HnEmIrwMxy6rHJjG
//0pUShOS5w+rThJB9ytJaaLvYoqBBWhdLphdd9UZZOpZ52hnXODMig2/7A2DOR6
fuSlWlwvvvurAVUXNCOg5Y7JrT2lsYp8XfHalCiwGWxZD8znZ4E3Cu7HLH1p1CRq
ydXaEO0jNwt15BQeBl+6zBl2wAATSLi5evfeuohjyMDcnaKSLde72dDyR5iKBubF
wcJUDj8Rp2pfmB1eqT15Rp/mwcoqts13E/pXoHUYwdmY0+cZEeA9Te2yp94LaPJo
Y85vMHSA4ym1o/pNgoO0ZQoM1NJLTKZ5ZmTBslmtsSFtiZKPBnOfDiTefJeG370X
V5+ns9U6Rc9tfH3GuJZ36WtfhwkN+P10vk7S+h2Y5c8lm2yq1XZY6oBtrsXuTa2A
2O2GXoTGsMFzJcp/hMLpb3/z1tK7UKmOsRxjoSP3quP6EgXc8goie/2aGKjZi5ad
qGwpmcNd6zo9Bv/jg7/Mjp8RkWtjt7Ohcyjz3PwmThYHJXHYW8b57QqnmdnBo1k3
CadPOtZ+UdTHG6wlx6HSdL3Cdc3tmRTnfuqi/Qe6jBiAfZgmx7adIHWo4CRvKhhp
kpTHQyPl+QV2c3rc0I9DR/ZjFBrrUL+Bgsmjo/atFxDykTH1M5kZ5JC2P61jOnPp
MDO1kdTBBix8ziJ+gCWF9ow2MFkABhc1tb8w3YGqE117o77lUH9L9WHvqnvOy6ay
DoFcSZE4Zq6GzRVAMDnbMTnkZdTl+kPNNyq9JafA0qHlJpu2vR+E1jE+1pfFu0Ne
GajkNpQTf7ZSsaNssbzq4145opRdLbUcGHnjaAHEfrQ4VpAwLAMAk6/iBdnWqV2D
NmsNozOTNAB/357WC4BwRZ2TDYXC9yuFmWeFofUYDxXwaBUDuHBQps31BVHJ7tyL
z7Dzsa45c1eB7Bs0+bATxueF2UHujLwM6NjsrpffsqASBmOZ+rGnS0VCScCl6O6i
XT4CKXREcS0uJ2gP8W50QCG+EwA7/6GoW/vcmuGz1zLAvhOmxQRihQLf03UMj9wm
ZNduAgRkxIsA5kVke5wEcD3nrr8irSfBLf+ihp0yvKK24QPcgQZx3Gl0iCZh4+o8
ZJsdfMIcoK06/pET7UkLlY+WjM1fOznGlT4FYjGmMAo+5BFGfPkdgMS+JBe3zOzZ
tnqE6TUiO6ap/wL6TwY3c0mBlDx6nkOgQTmzO/42Pi6blD9C9lGCytPjQR+6D7P6
emXFFBAMkwUPMAVuf4spnfgd8U0I2rdUjwIjSW5R1ZjEhdPgGgfD4/GHXlurcPHR
BQD6ZRYtoi3F2bD93yPBp+lxUNItqLi93S3CAAeuS3cyZu3/Aw78PZbSJSlJpmm3
JzIaD2TGAJetk/xF3X/ANbxLlhulOh+Jf20fBJjav5SmAFaMcK+ZB77visSFlGc2
sXOASeWdW6+XdiCt3A9jTcI181sCjlopuPYoSaUXMGAMh4rJEmMkdNzdCrAZ3cXa
/Lix1hQJ+936NoKx7QVGaaIwV+qu2JM4aM3qXrnE4yzrMCUEZb5QwkFLVpQ0YIol
d8MYclvRbLPTefP+eHX8+GiKiMYCIZmVa0Cx5N3UYlBhwJ3f7qq7TbljZZ+CAvEv
BdFhP2ZZ72u1nRwYPwxtq47/+GFB5ur9/48VemUZwh/yUeDl67g4cjj++Min1cPI
wyEdwvuvE7exedsPNaU6MME79kiquYGJOWF/+HRO+KrNuDh7j6o10NEKzW4Sr2xI
0AmUkjXmS8FM0NJqE4QSDbYYXbCSPn0Z6b7SNTEx+Sjd7dXAr6+GYGEdXqN5IKAc
5nHiqFe68SEqM1hRAx8UZD22Ftw/XRo9fR1hIwP+VVFsc2jR/IAl76ougIj3HG7D
oxK/MiyA+oPxX8pLeyLGcqg1JEPuCYfoInIELTcdT4r292KTVLVnKOtgkeMypgqK
QuRcvRNooDNTBYBJGK6zEDlyTFP3VhKSEUbLEW/x2dTWWmAJi+nDjf0OpSZRpuhb
YEYwGdP4gVdVmfiMAKYj30UCcMQasS6PPHvsqyT9ivuRbU4zVvVlZ1AEVtVP/EqY
KhNUW8prT0wSokUsfYhEBL3zlPS0HmVJT1A4mri4BLgXN6lXmlxwpLW20vDrsgjR
5cfhrzL+0psDQfIjMh+1ry8iUh+G6oB4nk3mQY7fkfM5uQH5jHBCgfa7zg0Gn3Lq
Nw+olQR2f8BwXL24hkaisNbSrAW1voob/7l1ZLXmaKRdn4IjfrxCgFMjZYBYEmpr
sn65uI9dgMUtn3sdJgioeK8LazR2gBBHsdPVyYXu76olGHFbegxUk+fgGO1Hnstw
OroOUei2SXm9WmwK16YiCsG6Q7zl1xREYJPDbQXQEqZ3W5iM98/7HyF8rg+94C+1
yPlTgrQyKaOg0tTkxM7yxTEzZY5MmtLqZ91lunTUZJfLZEFt+NBwa7Jpx83Fo089
CeBO+1yLaqkbtJ6ULMKbJiJQ9N/s52IK3aXY8QGet4330xpE4CQJFE6SJkTe4YaM
JVYHpWGIQGojf5vs5hPbf53bargEgRMZVY8XF8nGZBr5qWBQMlvU9bSlZJLZIGNw
ijDzx8zWwAYocccgGzlhGOPDbM9VDGlZKZAdf2gn+x9xicS7++NCCL4VcpAGnQlL
kYS0S/DShITMEUD3HNdEGCtKC6zS++o7w5EtnjgUTXF1gM/4M7Xb74yfM5QFkiQY
rX5g1d5GdXZ0QuI7WWhDkmssZFOJDVa6tGVdt6FL/zDajMvSJpcrdsOF8eEM0sMA
7Et5V4OeVWGGIzC6t+6RMlGJyoA/AnRP5hEWPv/cSGbdFM0lrVr7cDIcDS4HSELt
0ZCw6Q1KUmZo4jNfoy9bk1mPvuOR8lCPuacI3MUcESwkHzVeLwHUgmEAAqoDxo9C
2iO5N9OLNUMFE4CA1JkJlLup7nP+pH9GjHzKLVUeH1O42KERVSDjR50MzsVMB7b/
OhVfKrS9SMLCyPATnAbR8Izu2Zjq1B/flpH1X1WadyER7JPv+1XGcv3KQbdkS+Ej
HsKEo4T0BfAOFbZAychdqYeaHvftKIbD1SXQLM0QYusidf1hOXm/GmT9S0mUw1lI
DqcREPB9VzbuSftNQy6bNRmahL/1I35Ujbw23rfoz20NED2aIw/RkvAwzKPIAuGd
xv0soYTuFGkE13e5gFe1ZfvqgwDtmqmanDhHfDhu/h/mSZsY9HWzlDLAZ+xCZcmX
BF2Buh2GovpFIM4v4MtearRt8LeA7KsEyCXvLJtC2zSxYR8FL2FFBvumNNRMyU8v
thRP2zD8j0NfXaDePd1AOM1IaJkisuH9mXqaMVF7NQ065geHsfFrNLUzHtrIFH/M
TQv2FBLWAjkEabfQ54HuvSgl6KsNcvaIUQGn9OY8pMAKzKXG/2OfHEw6gQuLAdLJ
Xea3BmfUHAtegTP6xieb8nCjueuaVAmDHEsNxd+mSPrmuP68Q1m5lso1Nv+pSDEi
nFPUU03X3H4lhnDacBOU7IIdJUQ8E4alcNW+YqXpGgnFEoTOibzBX56U5peMj97m
hePl0lGcb45aNJN0kVb+2hgN7xfDxm0TDgWcLFI91MFRk4u22kg/1fkiplkD9k6s
6svga6bDLggDknavekZoTXRx7jKqiHewHPTYczWBmYEgOHz7dO6iRU1C2w2qXI7f
gkT07aPV+dybBnekMl9CTQbodSyDSmpf0wqyOy1GqYCI9tIHv9MJfPBZq+h93Ug0
g4wFhWEH7uoSuqL358ORmAb6AkdIfOWYwU0bwCT6MdTiDmKbdrUJ7Mu+WmXkm30w
7rnisPU+OBWcU3lO8sMbFpR49j82CoKHJLV9iPbReOpp2HjHYWaBIQNlqNkYUv2N
V9YR7IxptagH3xMoHU8uWC/WGjIX8QiNIsRFN+3AFkoKQMfWPFkqb10cfJ8EQ3F9
2/yQ8q2/inP+FNfDvY/NixMDPYJtVBA5K9P8fjktmGivynwuIZIU+4CUD1PgWqL6
mgkNvmaLvTFJ/QnJHu105qnn26UejHT1ogucxNYAb/wwy6ON86sMxR/r34iWQUG9
S95m4aATYYhrxRomqpFH+a9mgmEjAalRm2sPzg32UdDdoqmX0y+MSjANBaYvieiG
5Jf8rFC2zljRf8bgEwA5kVvVPkRx/zOVi5PNJVLI5LE6qi7UZ4mqct6My0s9zhiw
ocrRO05CNF3sJjbBvp6kIZEqzown8B64FrAfLavJEPpppq64JqnOu3RfkOLFuJie
u16EPRWGHCtlIT1KNENvxh+jPkuwEHUuExjfk+GZpyG8fcFOeH8XsJuMn2hKsy6o
6AmbToWvH2Mq6aQsiVJ4Wao5I/T0g2WT0HJLSBElRI1qvfE5t2ncfOXlj1UILUj3
+w6Vz4yXhLxKIL0O4fEPM6GWjhM0E/8zecVcZJZ+l6Up0uxVeN/76gvXolfviDW+
Okwv0Im1Q99/6LF889ycLeW/QXQ/j4PsJkNrwdrqQTy4YOPSqYtcz/r1d3Igp05z
J9EeuGNMdFgyixDr6J011J9oHQmasHyfqBhopeBEEWuGGkq0gWk+waVKgkpMcn+p
ZvbWSVe9VgjmUaPAIQ87mxNgBazHC1uPz3V4zL1xewMIERLzsLBMJNxOlyUjy3+H
8WMUZAic9BKZXWKy9ESiCiAFnq6aJDTV/ihZik1M6NBROLEAd560/7azITloi01u
2kZb7zmY0bsW9c/K6C4GhS747QUm8DHLjW2v7flhV47pO0hzeEamVQ22rsaEuwn+
mpD98M3E4IkQ2Q8L/XGgAbsMl0eUfozeK+wYIqdcsKN1z70Xjz1Jv/AGWgbR8bDR
3C6xkd5a6KqSMiY0vzCjWmmDJ7SLFvmMJhSV5NHjwDp29yEFTPJXjEePXg5q+Ci1
Q0NXwaddXLO6L5Nm9ZMJ5vpOl+0+l6oVW82OshGzeJWrWJuBXWHIrWUVx4pn+0Yo
zn9aajBDHYrjXfk0ZtlDnLBv8uLCW1BSfCxN5vf09oT4tp0lMnbT4yL1StCH6x71
bVwEeN5pVtapEHskOJIopExpVmJGKzhlcpUQlJT8aQHAeYI3WDlolwJESs+ldwim
4KT1iDJTRoQXChzKpNtP+43Y9IFLL3CYJk0MZwCSUqVkF/Cd85qQKWxVfbPQt+6/
pGnQxfhZxMIlethMRk+lVOaY3eOja4INWHNYitmHEmVsd1b3RmjG15J+5YkZmZ6v
q808BYYKOc3xs1DO56kz4/71e38x1eHPOU+TfO7NDt9SN2YjmH6yxDmPWVnwwKtp
QQSIMI5ejLzAnOIujxdra7/ajPpEG9tU+Or+bcjz7KbUEfnov3vpyoyPD/bZXn9A
JVeFtEeRN1H5ndyk41j9JlyXjolKwtaqRK7xL2yRrdifmMGk6xhwT1KoUmVcthuE
2kCEVuIy3aeQs0A5HpIM9EwRx/X6VP9Q2w+cCAB0P4ik+tIMr1e6ulGJpULt2bbK
DAyw3Nq/IzfU46eb+RKLUq/sQKna5I/yMxXM9+AIbfamPgtk6i3aVY3DHWThD+b2
cRj/+BDHJZFb5ig0Gx7RU7ZUJVBmHJPhXN1Rczhhac12inVZfy755ZATnQ7G4wKA
LikxHajPVDEgNLgC8t/6bwok48JcY7C5pZu3EOzRaiJo+KBJjnajNo+LXfPZd4Mx
bZ0lwCN3tYtUkwFv/p4SsM2ZoL29F3lLIenR1JeqZz5tnR6HDH4mDbncJjSpQApq
6BN/8Y92fTUFsP0r8SNU1PpDa64sWl55M7OIQ9NaYVOqcKca8ZpE7cQdOyUG3Igj
Y5eWywxgQ75uWBQKYaXDuR+tORyy24+u9SmsTCPYIq0lEb7qYSSPhmeurdT/PTtu
CTABOm5yq3iscbegkkHDHyIxizym1CbBhOMaENl3Lp6YJpk5gsdDNSyEi4yPH1KG
rNVVH/nrdIhhTyEorXcQMLvcVQuqAUFLqq+FzXCgY27FFnbxNCOpe8CD7tXgTecd
wmdAmE92eMIUHHM/AADGXVTox0yU4GIDL9dMCqDL6nolHrkEaa9hZT84LdweRjDB
IX7g108dYZSBNuubgcW0nOIrsznCoZTlKZeuH6sx3z7Fnqfdxx6YGg85drbu7bD8
dxLb/r3TLJT/R0rDRC0LguYKrCsvMrDeeoY/W2FwuiM+i+BAjTK1UkZj7fbiiZkr
fBX6BkBQ5TrqpeC3PryP5iP/78/LD2MlYdXibM7PiKzy0lJXCqr9cBEfswFROz5R
hobooe1XCtAdj092vvXQmrudRRlb4mk4BVdCmZuwExmY+qH8T/faLhJlwn5xFxVc
RnSBUdK/nbvoAucCwVTr3R/l8JvZz2/h0ik1zXx45Ci5xPZ0vAHO7sTBDtAerIXH
URrMVu09D2YH3c2+izrNNLkf+dO3dRJlXhMIO7whFmFJfsWYzlMErCrx8lDvenR6
MBxhkEhBN1pet/TiT0JEz2jhefr3kqZno/7Kd7iGqa8vX/A4cV38NGxx0P/W/dLk
V8vExT2DQPGCGaciYSS1aI1z8V/v05RMQuMAWxwQzWvOVBYTiKw0A4vkrX/QItu8
bSQrd2LBQyibJUPH2+TK0mc2Vlg0Z+p1uQACQCnX/8f7IXr8iAiTuqubbfbAKYsG
98WLbRtKE0+Opl1pMa2NOdeIUmsH9rlENl7cl04NMNr4W6w1cMquxFmxkOF4WnZz
4VQTxiCHJaWOhidArFpe7nxTtyJ8zOwzs4YFJPnVCn2SNyMGWzX/yjFrbWaq1xzX
2tvpiCLyD+V3SII5DfXXzHaix8Vyr7CXTflrPPd7g6uERtcmQve/+dmxKgx3El/A
i6H9bYjWZpN8/zj4f5VV90w1pkwLVjKdddryfjdrBmRJ1k+clOnK6M8h40sz+rFP
N/KE8cyfJeza9lMxEqDCUa9xrfz+tc2uZ4uXhI4iwEBqLDDYr2DieYJlUqqqBKma
rPeynKgmk10c1SSuRuMF2IseT0SCRgPdiQ8543+MYPCJJrb9d1qUuCOqYQBxnnOM
r/yzk2BCvyfYkURdh9lYkbw/TWs5n/Omtr6m9yL5Jm0AL8lXqCRkkU2T6XtEgfW5
nUf5Cg4MMW309LZBqvYt/eSlI/6Jduxwn0WIxnw9HyrJ+nVhpdYKuB+7LhrNzgvi
WwVzEJzoBkHXiudj9kSl4hKSKFK8xV96hmPM+eTgkStslSEFtUZJy3v3dPj4kGgq
YSoB0XoXhj25SuYlpj862a1B/TYBf6zl/Ym/mg1CEOJJj/qIX5u6c5D9xOt+fLIL
nFGLUbiGGwM1rUrnsPxTu4eSsCCLE+TEuOs3uaKFURYiZOjEDpAbUI43WJYUH4Ae
ttOG8twTPzZsApiYEhIgyrPzKsCxQZ3gUJ2uRlUDLA0Y7942IE42NVFHwIk9QzHA
zQMfsnJtAD0xuhOoO5xA2Ee7pC+nKT+5Y5YAuev92K4/52PP80d1r/ZgRLRW/7Nh
TVvqiikDtQLDNNcnwR0Hk5oxJiGRyhmu35E1cAwBA9fXZvpryZCSa52bVY/r0R88
LZKsVd8Omv7WL98vLOHmKu+HKbk9ayRuUnULn+MCMElyvVFQXyGNn/GDHkbMXC99
EGODev6PWvZxFWxtL6MjAx2ph59yugMYWS3i/Jnolny74MFrC/hteAEuatvz2V/Y
wJsc16ONuKkoU1VD2/81eAUjsqejuuKCckrFrAoU0RYDa//uHHISMku2h/CvqyVJ
1CSGxJUX5W+XKDneQLWjzAmT7BLkHbeaVNRQe9rmQHBn6Sk/XwiaECkkd5Njvtzb
cfFZg45AT+s3EEUKnH/1QOsY5atRKckNzuA2QrKHQtfnwDEyNzyq/xaKtueQRXzq
hR/ZDg6BKFPfT3xTvz336qq55FmGz5xgMsRTV/cgibl1PFcRtUaPh3aFE2GzX+Dn
ptMwog7fG1P/eVza8/y7ISVz0BcyZ+hYqDOK+75VnXrXH8JhtDHn0ra/QMKb8F3O
fbsxZ42Iq5pIFW72wImEXmv6n89VpMf1iATy4zE9xRBer1F6h8HERWR5VutQlX+a
4ubeMvKOkzb+04BZfkx98BMZh4/rBOh02/7UJFNjGFGlXtN4Z0KOs+CjiSLtfN2Z
BMDmlOmnxvpbwA7mrFVW2lK2012Qg90hga/t6ueQWg/F8lHpj9lXpHdfn7ZCQlL+
Rf6OZTZqy2ZE5MDR13Wgtg9FjWKBxnkZncVH0UH+KdEVomqayjD++g8BBSj3357K
qoG0uLImYWtsjsFQSDPSM7fng1aL1hqdnS+9nmgN/rhGjD15dHRE93UWtl7//UDq
f2w5tu0UQ8cQfr+zzu56db8cw9QDmPQoY9BZmnCgcny/TSRr1OGYHD0a32wwfBWR
ZeDKO1zXMT1eacohpEjDf+OIqKsZSdvUCv29WkXnT6zkZEVCLZwGujXbem+qAh2r
qK+F3afqVGHVgCh0NkuI12WLsjSge7ZqQi2LBkrqFsxaxz2heobAI1ZAAEe2FcRO
WuPPyoHxb1kU6o6MHw0gEQahxSpBK0qpKvgNFx68FRR6nMz/qLg9rFnT06lLqeHY
oT9IQdln42+4Ji56m4W9IXuvZlyGH7bvT7OWLpv1nZ8AidaRAmwUt20kQOodvVGM
yZsXvogrpIp9BVvHNpJvq/kTTwKLQTYryccwmnsuhgx4NQn8+oCrf4cXvCC4mqny
7teREkGUk/7dGWjgaBnNxe8CjbbaskH0Dy8HB/5sa3MAirAnJonpIYKqszSWV3yn
2/qfBlVNxOWJVTrNzvtRZx484r7ro9dzW9YftDaEMLemN4ZQLfi5/buZzxaEjIZS
Zw7lKCOrZwRj5+u8hF1gsHzNjZNOHVPfgogbIFH4HAd8JEiGsm1Hs1YFMunYfGaP
u5LnHBMlwsDRwPeBbKB8Z7OfTtqRy2vjHg+z0Qvu+rcQYfxibAv86GSW6pCJOd1r
LYFvN5zIwjkPwQih+78i8+knRwkHLHnoh+BC/N0hpmZPYWLpVOSNkARjwK6lh2NY
LDzKhs8t/Bkpr+yJoiiK76goHSi0MEliI8AokY3FfKiKFwFBGCgfltGSbIB1S80B
Gr9LPkvnNjn/9r/JvOxx+gmclBbq7rSW3MJhjLhywV5evQuoCRPw4ekGfCZWPD/J
1O0+aSWAt80o4T/cw+jvw/WD8b9xT5U/3Pesh2Rt93iPxdUd332nWm87SYZpWgfT
E6YkkZWNYvXyk+w+Q3Lkm90jv7nGIXQY7egWnMv6RzITfK6nWw8EcjoKX7DdaHgp
ledU6ZgEA6NsBiuj95H3qA9VbMgzVPbDU68Bh4aoCVANVjowRa1P6Py4nx8TtFlU
ZxmviyLsjweFqzJ7SFSHIz8TnxALk4zVjlvBfWhc2SW9eMRqeKsBhhbwyddtMy30
Un+OiksUcyWJtgHG7b6bZsMDHykLhPfkFTX3N82OfnXxoh/Ji0h9oC+DKRW9o2FX
lm3/CBDDVw/pu/kllKW2yNPDL3Z8QHGQgVkHkVKdP7Xvay4km9Qhd8L5jHdkMs/U
hXDVUg73SJEA/KacazT3nKpndWZ2eqwLoHhSKWOeA35bAY+lO29/b8HkVyQun6+L
2w0o8ExDbnTI/5rtO10b5EZTLDX+KI09tCyuwvNlZGQCOH1F5vKxbWkowoMTvxjf
WEPajhqceafT18WaxzPl5Qx6Nv2am+IbwVcczOV0wNeIufZR/XwzmRlZUSTJbne2
tf7+HKeWbzjRWuR0hnUStALRgDYiulJyshTKGRyL2JyiieLUTN+hnz7+4MYEvgK+
esPR5hl3rN7iECWqdoJTVVv1K4OLi1TXgoCYovV1QlVXpYm/RV1Vpx0rVs0f7sOV
ype+a61OW0f+v2IWJhv6eni1/zgv3HI0J4ddFYaM5/z4qAk5VqII/BdRiGQjsdYy
3s+ysFnoYCdkY/ND7k9bvjhwDMkRNmfbGcVmq3jmq6NGVYWqqc1slGxmwQ03nUoY
ST+W8zFouyfidJL8quWw8Wdmdfu3Dek4yQtm/6bpz/rSkJ8YgCi2zWQqa5N1B9qM
auDsSc4XfjLvGkZ1Ldu49eguiTdYTGfOTTfN+Mnaw1mCRj8xTd6OptwZbXKxuGHs
dntJkfVeXdWXWw3qkLfjmN4iLYgB9dwmkC8fJEAeTcyuHvh8BAGW1e40oir53awn
sHnp0SRuZodyBaQMV4hhra2RGHW0BhXrMl5PhLC8DcQc3teE1iRJYfUEsY8VFXDA
CUG5MNt2c11YxtWzdUn5TZ3TUW0SpDJWG7HIfvuEGfgBMKNvY+sPJgbTHD/xXKxG
NCJvp8Uj7ienqQCt+NAXTQQBSf5mkhMeeczdjAfM3GdQ9zStx6m4azW8W65kzXhf
DQXEpZtGLYhvtGYY6d5fWdYurAiv8tryD1ZRE4mu67yjK8Zb/2pd4rPwq9Ofo5/r
dHXCYc8hT4V35094U3fHuChBtEIXP3Z1WJ0r5ZNcez4lldc1y4CWhcllZvyYK+dC
R7SuFVNM3WrndSngl+1/MTTol52sRs2fmePm3rARJ3DgDoSPabkBFsb/OMBBazcG
fjPkRygoZgnAI/xvzb2UIsU1v6EdjjieMxiZpYDTpMSOebkYL6nY0fw1joED72Jg
ylLrJDy02Qv3PKTAWvHrKDFc69F8ayG54S78fGoRtlNtvcKOcBBEbKzYrSuOasM8
X0wjYnlA2S1TV+CJbvJIeQ5EoCIDcWLwRapHjEow16dTokTWv7UserKWAqqwUKMX
h82VnglRXFmFNH+qb6eG/stMaNjsXWYHdSkBXn29QKFATfyGBCvdq2yfCK1iJGAu
VCTwyY/ODCip0fA4OgP3+e2Nxoe6j37APanfBdE9/wMxjAcqJYNujnmxyaFpsoND
GLGZztF3y8Fk6mMwhqMrnwgZJOZSQMgqdNbpU7Xs37CWIXuD1RUNggn56jzeQqqS
gMKLB1EnSj+etg5hHJKH0EpiqNzkn5MusTt/kMUQMq3ogT6B+aDcWAXaLdrgHdrX
uSxql0HnsTnRt9HUKsb5lqvf8+G6e3jr1yG429a8mC1EPvT7Fe3fDr+wcVpGUH4j
2vnSc+v+9VxQTdAzom8eL8IJq9ZjtcWcq5zd43y5R+3w31ec1gOjcdt5ObrSFoRS
edjSWm3t4IXUuEODGdHtQgVpg8xg0DrI+oghY2sqbRLI2RJTHOEX8JyjToKVacQJ
/XNQzUHWz47gGAx50k1VtQ9+2NrhvlX/A5X4bvv8A0OB9jTfi0bB6z0kCnw4S0bL
ZhmkdE8thvJg7nR9xKqAINRyfhtA0J+rB+FHVZ8trjbWvn5b8PrAwJTsQ7dH9Y8h
KJzQCF508FONOqzIzZkgEgXojoeAdvzP2R/TG0jsw9eBmPfzMLnzAqpDAuLaH6m2
513DvZRu2YKUBSLr6N2Fzw6WK1X1zD1lvbElRqcsYZJealJ/LJdcM9+SmEu2l0XW
OZ+muqszsml2f3ZJ2E+wq9ERNxvGlfCdlKg9OesCMVhFlt/qF9+h8Swn2VxUDiAK
uQd5t2QlSUZ0srJplnja4VeW1WgoFgGkeZYaGXoQ6UrzvKydtgqoR7E/aLyEseNG
7J2/PVUjHHihusOHo1kPj7mtPwSAYOU6DRrlbMymCK5oJajI2tOxcqOVG/5nrhRv
Xhz7m5ivL+K+O3+Z9s9uS7yx0LNSrc9NmExTnzvtRiz6SbCFxafzFujAf8WRmn+N
VCDZp40kWX19Fk4k0Wbm5AdizxMwjnt9+gexKwex2FzBmqQAOVxjKKlxaz5FibBU
sVKGJjHy/DBZc9314aae8vRuwzRcnYs+EvvMCNUDhsrxPtH3Hx83rDgIde3Q3vbH
Urv3LrH1ynOdVX8kL1550BE1k4j7PlAzxRkGZywH+X1pPWrWmteNz2pNinijquyl
GJHzTG7QLGbxM2rt/i9Cr7qNJQWr89vy87wZvOSPucQQCf6pO8NpZogLgN+iKIX0
uclTI7BESyOGMitUGxfaaN5pK6ywYciGKETXy2LUw9JAP+udf7n0pWowRSGxauSZ
v44Ndj5ZBfiR5fvJwXENbWI0wEb5lUjw1zvKQcrWWUa91EwysD6lPyOi2xCy7oPu
u5drlsVmTG/798jrtQMZ7hhtQkKEROk5XoUCRLdSgX3ua1qz2vjminnNwUmXRztv
adJ6nlN61yJpqyrPk44KvraAlP8MV51/Nio/dxtrlTCPodX/gwmCIGKdj68v+ke5
ucnB4m3wYZgdEvLLI6z0pGZTvDBueW+r0vGl85nG8M0RnbBsTTgyBUSjFDBIVnZV
/JE0nW/ByefcT12XLLvEY1yERKj6pWtOPMW/+N0lKUzclBu+VXzMUrJD2ZE7UEDz
7JePVAi9S4zu6avCL/rVIenbMBrgMJj3HC5nStsoz8IDuSBhCa/EB9P/RB5TXACq
j39eVF3PabZnMapaena4LCAk1slYB352EI45OAkLnBBV0tDPFd3kJkJUoK5ZiJUe
hfCxb/iQTR2k05PvBUZzC+yDTdrfyRRRa1Sx4dLJpNRZ/4pWuTrm6+5EUvnDSNIN
61Z4AXXuZ/5GZ4KfpjRy+VeZLU7axzkeobdBxjg6qYDFg2fGfPJNNNqnFX07sDm6
uGzQUHFaQclEz69V7AuBtGkbXKY0Rxgux94OayTJ4ACx4N8SRbeQhlSv9baETgvf
29m6yJotVOMMOQyi0QdfK6ffNdzxIkCXnrIwNXGwdLdM0qoFNjWUu4KqG8+9fTWD
hSLA6e1GpdVWovxRkxYHbEbyosELVEicISFE7N9DaKvfoJViVeRVTvskfS3ONPXb
ccNmFeJF1hyB0/pbMWYhmoMrgJGP/lLZl//yuSDAdaZdVRGykgwy7vcR+4t+eaVD
G8JB6GXM8Dx9cTlE+b2v4FNQpcvYBfieqCblS3FTcMy6g0L1v7N/GdGnOwylbGik
6UCfznv6nEOo79//AmxDFDxZ3l4EaiQC4E5/YHr3oYPpiXQp5C3vDgSWeDm3bxHN
EPYnvK6fJkaNax/Vu804oFLP18Td9K8MMFJ1Bsg23EmAVFnCql8N1LulTuFn7T+1
8DEyueTE0inAv4rPzKj7/Vp4J4vqTd8DlqeLgDnIqj4LnoJa+5frjCaSFpUhMXWF
pK+Zk5s6ZZlETWXU3LxFOdKdH5w+1lOJnaJqK9OWm4Pl0ywrcoC5jT9zNTi6gfRM
3l+SaUhkVXMkVWa5JFqT+VW9O89efSq9fajJnb3naGJ2fqmyiZYVXUjvwIKwoTa3
ejZMnjw962+X/PxdMqIiBFgbHcVawPRwrBgk5h5zh0ud4BNmNCBaEte5c2YVRBXr
T7QA/EqFbu43/V1lXziB+KcpiEcIeepVf831tnoaQ6mRWDFzBf+KeY0hVzzLVVp3
95HWkpMAi0NRaC6gvsR7135CCwyl9XOk/BKcNZgmZWHmmyuQUz/AST2GIZuAhjDO
mRTjsqpgruETxIZUJtclkDvU/VMXgwqnBALNcBG6EUuxQee4GJ079TkKmmdkmIDO
N3DjFKb4Ao+ba9qpMGvVWWaNfNivDHLqTSrGmQYbLpWtS5l4T3ovpRsRmICAYR6Q
gSCdQpv1asK97S744+8Nw8gvKoU4wyzq0ZgGYlTPqT4Ub+N/oD4RxQ4vpNQAaLDo
xS7B3YkKIAxNOW08H8ICo4rTi96rHhKzxLto5t/l25DLzJSlE2jkzz7Vub4Dm7QF
pY9d9ym/nVhcv8pYwrng+PGybslAnlupdze1YdoYpfk2ESsjaEE3Dhl5dMgh8Sa/
fqt77vKFZrLnyT5OPxxV1mRuSRzOPGJP+wUos1A7RvA40NmfhoJrPR0Xwr6Md67p
8N1+9eaqPImzLhSCVcBVe90YhFWw4p8ziqJoElZTTNl+eKcR2KrodmM50cJfe9pw
5gjd2G0+lKlhpEmPBPu8fhFRuOgZJPUxEoEviaoLPaFVC8Xm3Za4sY0l7RbzWezY
Dv80NJTaRpPQJOeRotMbukzTZPsYo12vcQTXrmJHMmgrfZjP3f7DbmjklwyyIrpH
S/oPhM4a5qeYxmLT/rNUUeFAnMu0dxeeJAvFH9CvGBVTzR3cjyohK/HdMVCMrviF
1CIYVYdnBSZIvI75fCFfZegHT/yDj6urzyXQlHglmGg6lP5mhemzrU3CtVJeiq1a
mCOP0TAHy2BB3ppwkaNgzizWHzsEz9trZLDtXsq6NZAX80RSg407zZgeAe/Ml9xH
RfOarpcQZCdLP4IULfuxOqOsFP00rgzvj3gIusMk1+2Mi8oVocHxKmtgViU9jeQQ
TDM1NmyaeAJhhlNXZ/wsgiXAc0x5KCxcKWZeti0+hTuJP8Kg5Cvgb9SSiFCwUr3g
eN+LncJ7kpy0yFJHm3/NgKC07SMxa85Lp2uWdPhicjfAjScFyw0d4lkOjISLTnrG
3quY60kCYdmiCQ3qgZYBJe4w97AQO/QTSYbwjDnW7uIP+qwmh7lf/yI3L40XRut3
znLMvsCYAbMk2O5aS2bbDKvds6sAhXIZFaKs6u1tAcRBUxO5hq2ceEbtSKKxSqs8
t7vGQn+T69GnacSV7n1JJ5xnKmfFwa5Mhw3BlTzDfELKA42jAqWEqpQblgT6ysuc
737rgWnwiHyrZk21K1hQ8Qufja3IcZmeziUFoaypd06ZVSl0hGmxUHLhOipMLGPl
9jkkWZ3+r9qh6Uo83oHJ7N9mGKNd1hE5/ZrBUO0EFrcHM4Vil4+NEU/HR++kndbo
Gf73QOzyUDY8tYN5DFNoh3bJ8Bzdcm0pOnQLD0Hf0FC6w7+jpBNklN1/gHiwfEbQ
sgHtk+oecjOsA7sPCx4BkMu8HHZU7cyq1/LV8gxMuB+pc4ZTdBQcUuT1B+jLG/VG
NBLkmOVI9so9CsB3OupiPZ/KJk8AVx98/L0TteY4cEZdJ+TEDck7BUZBek8iL04Z
6sGbKTEYsCVI66QuTxogqeUc5LCOrjPbEJiP0/ZDNAPyzPem6wM3mGG9fmUdlhw/
p7RaNfg59SKZ5hGrTQ5serO09HseXTBlS5iZH+aFDOy4ITWi8IEczJZl4c2MF8sC
HJoHme3LXFqN8aO9BstisvLre/+HEfe7uUsLy4o53F5QFyGV9196imqmnay8IDgx
Eb0rgigOHMpm/oReCPIoTeQzgNDRpPZ/pu52/AR6RuVFCHlPTBMDPDDEEpM7+492
3py4Xwo0qlDBmMrzn5pUtdp10G/rZHfzf58LeMXZQiu5y3uPLFOCURJyVMOdMHIs
GkKR8Z0b4sQ6mG6DPafZUcuKHqzU4xELVkPTmUcdr+dJDlS9Z+d1D0g15lcrbAQK
vmQVtl8uN5N1IulG0fIBeu21AjA+X54v2qa3LR/dqe2jYkaB7aAr+PmFLJlsXI0c
Z1xsR3dqEIl/8KOJzlgFUVjPWgQeDrtsPhHb1/ngwO07BzJEmFNWaYA2pHkI0GzY
gtfGrXJL3peh4QD5QghZhj4Arzc/bRWmm2tZBbZjTWqTZuSOHe6Lz+A1ICIf9gvV
tHI5DN58pSgyXkjP3XWC7aG6OrM/J1LnGRD1aIOpleeZGhY9sxLPXIl7xFb3HYXN
r6gwz1wYBye3k8F2tCMLxWOc2rjsMrQsHjJBJGPtaGjx/o82Fsyp3bCyD8ikZkKV
jg6uupYNXf33AcG1lCTkYwIRp1QRbEGgZQIO/S5lbklNiXQErxYO6LraSA38LE9Q
KSCNCbSY2ZtvAqKLP3ECaEaWJZRr+93zG7yfQL9irimbAiYznDiL6dWk5DgzWqBp
kllQKCKbkRgpZrx4qyC+E5CHPQBs0MlbK41V2pMy090GoosfN2yDpfX4OljXEuj3
Kxm5pYvqL/pA1ZuQIC/pLbFiqyWUUXtq5fL5KhQssIlMrN+oGyAfJzOLJ+bPqPnw
+soN6xKuMCWIcrZAayu6L4yqIjh7YpmJAIhpOOws8nGh0xzT/AeyQPSfHXDPst45
7km00xe29nPBkL9Z0G5CBF0FFjN2GNvijVVSrAtbTNW2brh+//m8AU+LHZXCajj2
ijK8pEnIkOQ8uyLVJkbO+OX/1vw079Aab6uaKqVZ20rKlALFHOoGPvqjZwDFbzdQ
V+6j0+EaPa+mJutnKeKd+qaolTMsXgCg6k0GULsZjUVyZpzvdxioWOwOafWBivEM
JVvOgPN0N5jRWrMdEeaeh4CRdKhp0OnqjtHsgs6vMiMNab88IlTdINI7gY8GLYG0
YHMANv+LmENdoi+vbXQYFzyKbi++sfh8t4Y2mfJxZAbTemS6elMo6XUPN4DWBgn6
3ezD1A/I6vzbM4PWoXKjgNRbna9EXXIOshiPuJY/5SHQ2JienVQqpvkuNpR3TCrg
jP1ymj5n6mteeMJMl+73LWOglyaWcLCaprm3T/l5D3Txb4SqFbEZCLyDtRHeUgvn
d7ZBSt3FYCxsE4BR0XIrWWNjChVmFo85hIYhCGHS1TjFfT4KjImvbygu/UibPSOe
/3ix94TyMvmLEa5BIuAvmogjfc0btgKRLdmJl95TjyVucEyOINVqRaSxzxyTSr3Q
rSrCAxZU8PpsMuMPv9rftJYHJXP0n6Juqovp8Vupt6kn2mQbYdC1kRn38ZDzTmIc
d5DMegsXjLEmRzf58oiiK+8FA6G9ZE2AiLllgUCRbnLKt0/Rp7ehLxMsgxkLEN4A
u2XdTDYQqNSRf4AmF0u60f9VPuEr6P4tO1LDOEuDwiSR8RPW7MIkwdOnnP9TwWAA
QrwFOTKZfxLy1fIcOjtG1LmAJJoH+KoxQDns1B1uCNqcH/7nqYDE8bylN30EsjkV
GcNhYSfxAZenUH3zMBkAJQT1MoeIx1AM1Rmpx1QsJcRBxfgLymqktV4H94y4Eahy
5WTG8inNB3eouAZIXxk2eA59KeMMHzcQAQtCF4AF607yXzFfsWJoDUgeQbaZzC6/
vYUxh1J0RKw9qeT+JY/zDkMvpqk3iDtNfKLiXhh9A7ez+j34zqOZ/p+FIh1yOOzS
ixlF5Hen/blFPF7E4qxAPgNV1mYUmDobMee9d0mlgylb8rcgJW8IjP4ZDnxzVNdi
Y5Vj5abGVU3rQbDavSiAwa/I8ML1/RK2NsSMbqKVVcqb9p1/lUcgdcJ/ZBZpJF+9
cUYix0A4092rj0n/9XKPynEnSy1tUdsrbkyQSn7VHVhRo/mdhDQakH00L5STNhgG
+AiUkw71qiydbqruazpfmZ+QywNPyPOAe7sUZlZ8po++nF5FVJGDUOgaIpJcRBE9
cKinkeS4q7MqdNkRmKWANCYR0hgm6klGV3ak4hz2clX6/RTu3I0BtsRWDuiab1Ne
rUM1eFwl9yp7WZOVg9N93fBoxrCp1zm52iA7RR3KkiCpvuK7iQUq1BPU5FJSjgHd
r9wgPH3zrtAERHc1QyatypAYdse19fEgJq3tJcU+yNVkRJ7ZRR+GWqFhJM3R8k/A
4KQmsOoo+xP2R7m7mRVKej6Jq5a3CGlmMHiLOD+fqqs0Pmy6ybYIQy31yW+pg8KX
Plj3+tA91SnlcZXZxoftltKS6gtQXx5MOrgwGbQSl2yrZS4/YmczH+PQcjEppEeP
Prdx5G2Q3+6PvkFRJBa7Sqg6QxVIYFXDKs+msMHt+opy5xXoV1YyqXhNveUeTzk9
qdn2GbyupUwFTEvhdP6Ts73o2TWL8otuzYjfEKtAvVpX1l/PZo2q/ZXPrfseE6TW
D9lSCAgpPX+3g/XW5cEkBw7kJ6rfJ1hBxuJrg5snNU+FWX6YmPjRHXLdWV2gbXnh
A3rmg5zc0cNwSP0TtMY5DKhgRS084JH2rrxF8XMGoEomt7QYXSoSRaYxC754XNIj
E9wfgKVYsMKu7wwWAhxKp8C5iKPCEL/pBAeKMtqmCm3A9b7iT1+WQpGLvQDMKR2D
Lldtx2O5S5ago0Al/2T4Y9VrI4qj0CnIexi60L2xUKh5Hh09MdLMAnFXruJCqt8q
q3dRFQsfhLBApGV9ctdb0A0jQjg/cG4p7MmYrpJRBmB9hvn3ueL1GMF0XX3O9Idl
4goLrqDVJ8c0TU5ElhQqnlGDtb8lw9Uygs8ehkOJNfBT7cZ8TEbKsWF2UhjvrUYY
WE9lw2AznNwVaMQYCeh2lsXapiISNfXcXvd7LZTmXsGB6FA/f1dsG5ONr7yMHJPX
Z8Lu5S9fNxwkP4IMEzygCBw1CYPkTBXED5dFtF4je1/wgbROa/tG2CuBMl8BTx4z
HSGhlKdFdw/GZllrwmZdSjKo+eY1xBJE0OPB5UCjhrqivBP02QkUDM86C96yz0cv
65IlL4gmZePvyAfAzA1m28y6pH9lnzbEnwlFxfehC7KrOZLlWNu9VszLm77BvcbA
2r1dlM3zGNFcsmDv7G/dH1Ss2MkkIoFlGzJJy8ce+aQP/PXYcZom3L0Z5tCSaVIh
G4oIit3nTqPV2h1FsCj7IwTuKT7j2QdkuSq12glgOAQpR68omVoZSw5fAHthTjae
Yx3BE4hClBAP2bfP8e+KQESYdT2wtOx7GQJuiBwW/Qsk1+lrbIqJuopB3VlmGK7h
I9Ky0mikXlXfoakQ56NzFUVUbNkLHNra/bGsB7Dj2iAznumg0NG1B+NwJSMJ5iUD
hsGDqBMupjqr/KP3baBouOxWk63lrDcIJsrg4paTJz2RB5h+VNBQgWmsrnC8iZ4g
53mhIsgDkTkg2fvJzq2w+9KPMyaFQaDK5B/7G1REEJWKzzNuOgbaKcwj6/T4xGWA
y83vKRlzfDIpgFJvJkMALjhdVQyd5ctQ82x2qP14MFMLkdnBTQa9pWvLrYWdLqxx
hzrQtt9RnjxCyoYWh7xfTaVeGadrg3PTLrwaREbvhpkgXseKfd075EcEQEVlEMjX
/ak9rTllP6IdU2ziuDRTlwO45sxSWfJpSOaoCdwJTyg6+se4sbD/RfpBxoFK53EM
R4P/hod377ghtccgN1b2FEjRchKroCoHRRfZMJPXhBOntPjS4FchEXNIt36i/nWE
3UcOJhA9ZLbNRcqlaNP+uZq+46QhX1fowv9GcYrNalxI+tHBROb6XRIPV6cQ55OK
xnBmwzKb9QktRYbB3b77Z3pFif4u0sm6Yl8ZbDxFrhlNQYB0YLul/M4dlCDLK6Hk
o2nZQT+6j73ZQ5SJtoSwLjUIMn1ATzFrdhmVXcLFnlJDUrGwSjwJimt77C8FLdS/
5oZYJOVdb7RCpwpZKhqRtSYCF2LpfbASquG66GTf3E0Og7bSli+dik99loe/8uH1
gT94bCpUYSjAe4K1EyXu6Zm9XLodg9OyJlIpOj+h5I+Ob1UcsH5kpZukULsJlhvJ
pa/jNzP1pbuG95Is2LRMXW3mr5GxTKl3Y/nvqlyMUIN0udAuC4uajuCABEQCxe+G
Mup9GCQNiKpcgpxX9cZGEjFKpPBJapqGhzAV7y77+z/pl2EGxDT778ltWzmDugY0
ly4pOINzrd1oxrr8foRir4w4tv907Tahz4nngYhzW8J9gFlKrm8aEdRFrLTDCKmx
L3AO7T42zVljzXUY0UVfBhQ9I8YTgXY7Tyxe5l6xkiaSY2eec/H7pxwE4mQlq1Uu
2sQ0bb345ou7K0pi6g7FRBeWOd2xPcFAtT03o6IEOeh+OFM/TiMqHaGU+XHcF9tM
XVlQ3MI0bHoMaTzYyKZxKUTACEvZhd9drWOR4XXjkAq7m63JF8Xsf0ZJFyyJFLz2
RFlLHo5Pizdp6s2xaxkyvNOqYFXa5Nb8GslBEVU4f3GJfoDMdnpX9lHPa/DDbeX8
I5bqAhmfwqPPOdv8OUijBIlKMsL4HXriB0eiUzbYcbavLMXpNvstZnWGFrImBXkh
QQM1HQQEO3087Bz8OywWgI69VyiuiZsb3Xg0jPmBiTGEkQXCrfg7b93Lc7J/+ONA
VksSd46/tZbkDs8PUHO2bWk11HNz7MMiS8utaACoMIxhDbFqeoWQeFA6W82XfBqv
rwZrAq0CRSiTSdI/Q+cbupbaURBJf4ziLOvh1vqAZ1Tl6BwZetZ5/sxjZPhlAbSX
xdoIqu+1tthZbQeey0mSGoVA+AxiF3eM+FoBmfUC/SIEytM1X/4zS53Kyt+A4RZT
Ptk32JpR5ptX3+1DDHeDqQA+UCki3bRCqUmx/GggWvYWIKQVcTRIG3LB8HLkxW1U
RJDhun3tz1X3nRtZKp5v1wqFqruE21F6PRy3AKjnbzFrfr/Irblr2bLyqI7ekRGW
laoB7Pf9O0wGKfpApyJaMGhAdAvS57Cmn9RNnbV2KSpJSD8e5obhnO2wka21I8vJ
YQEEp9ffv6tFJZ/4crgnppRxLHoUFtKvoH/ndt8ARvHzbXsxAA48N1xpLdLdEZLX
sOHqMSqegZHrPJUgO3GXS8lxN9EySY45I2TE9HD95+jnDXjLgoQUm9QV2TX60+k2
WQqx9Qea+YhPOE//2uFVsTdha844YTZx7qiAoTGSSuCpHzGE6yJObSiO4rDrQTTT
YUct2vwUmQKb/z3PD/i84PbSetGxKsO9BlWgfjjwoCSVYz2eBCAKOMpvZD9YFiOi
OSHWGAhI3858AOHW1+wFZVrPZ/j/FKZhjZrvfVh9mUEe6nSPc8JGquZwxlDgfxMB
uWL/YrcDDK15y400Jk5Ni4KGwjLUnqYpNp2cBaZSuzZm1VyZLEWvLY8ie8YngpDe
DAv7Klbc+n+w/iE43RSXPYkuT7Eed9gUESc8OMy4E1ojwVKZ3k1ss2EndFhjVPOc
yn+qQIyYN6Lacyi2bvwZ18qc97KvrohHVOyVV/xpgso570J0iE5NS7IS9Djc+nJT
zPHPpgWzNsLBhhs0wMw96/saiaIDD2CBFa1CTmYFcugf7h40eETi4UOxL5x/P5AK
YBYM9LesaII025VQ47My+CzhG/1XZQmJQArqxZgsm4Fe0Ap27IJ3ND8FF0KpAQxt
o9v2QAeDhByl1qoRgKWl474aTynOxCykMceRnUvA+MZDBSkG1hBpjK+uyl6MiJsK
xXWA+k6BrV2L88p46vE9r8EBsgQUoTBlFKtPaYZK4g5u6F37J5CDWBbb8K0Ur0ZC
SCKtSAyi1M1xFHGuiRxj/jI57hxacDltim0dJmYdPh6M6Mv+DPMdOGmxvxzGGdbN
kEQKD1sE+AKqGdXSBEskCyD6y+uV0zYISbemFwen3uTQbIAoYXz+zRym+ofdiIXg
7W32Tg9W76EK8e2NqNTRAWmqyC6bkkWUfBwcoyN4y7Z9d0CRpWhFBBmY9xvi9Hil
Ye+N9NDdxOtaSIf/UL9opZGYTp51Y42iNw+O16vZCHhJfEwz+FMc5lGwo7MZ+6pp
J3hhV0KXlymJhbjZ5/bDBmX2i1D2RdcXLUhdqyd8ia12z8aq0iv1FV6zF4/278ND
+XmgvvsMTRQva7eouCzdetQculAf3H1K+7e8DwJ0RuEhUi12KPpsSJphivSFgiyE
qryB3Nu4ASYbbicqPx7PN6EnpRDeq7ynp+qsomI6nE+kqBI54fvqNJtF3dntgJUH
yNPpQdYkfF1I8xvPJ1/euRxt4frdaaiPC8GlSLIMaOAmTSPv9AG0jAsXj6gyZmY8
DZehOtgWr/LzqdE9LMbW0ya1cP0uOFs45LrsOrENfboIh9r5U5Kmef6yl5t/1CXw
cT0rttg4hNgUNrpkMyFVsU3xXep8YZXg2j/bgDNrNnc6wHPYgvf639TOIIcsrYeS
DvFd9YVFLZgdufXTAJKIOC4h1yVm2qLhzVa9t3Xg/4oPcLURF1zK9k/B9jLIVWdK
sMkp9hheNgZg07izOJYOzR6hS1MZEhDeF5n+Cc7QykvOaDVqyNeb3JkAwSFWQWUo
X6TM2hpGTQ3TZuJ8c1xfPcrEWq9wHvI2Q7deDPutd8gw5HV6wK5S2tmMSyHjBKmt
Byt9NL6ns/HIwZE9e2NGg9yRkY6p19IyzNb5oculwwQJfvbR5jRbtBNWW52oknf0
Zyk0u8ejPPSmxeA+UZsfshbihDrh0CbAsTFjUjxuMpAfLPv57faxshN7p+LS8iZ4
aMtgCrs1ZBaq7QNn3QYGZQwkE0EXShRlWRaludDYwihAKKlBeZ3ivhf1AoqMIJhb
VYaPBxj9RdIt7S9oOEjBruG0HjRaJv+GtpMo79a+OvcxIcDT/5oWYk42MAQ+SaPY
FLwZmCeU+uc1nUIAYSgjnErIHKsKfEk/FR0WhDsJNUaSF9IMTEpUZzqyNbjmFWbj
hVbFSYvd1wHxmr9JNN2siHrofHDN024zevSnioUCgTlw2cU33ICOHmRD567IOnuB
C9CCfMuJyh/thwU3TRNRJQSIJftEGqkAGH4P4GwXC7Tu4/PUKje+MYSwKDkIx6tV
x4eKnfmEIyS+os5zVMbboWx/RtnkkMnPEffMxAcP84bgMzHeU7a8zU8XYOx7t8kP
YaWE1WpfZ1i62HtDlamNQmXCpE7BKQ1Zar3/v29KhGSooe4O4ZBQ0wn7p9Q6wBqv
BebTrQC5Vb3r5/0L09HWtK8YL8xuYa8+JR9Zv15JEDHO2BWabtnIwlvT4d63RvPJ
tzhaw2RPLGGwDD0NUD65GZrIyYJYgD2kzb2jCfW7/haiy8o+0uEFo9co0NR6Pp8B
/wN5ikHaXy3HtS/oz+FAiDe66tCKSKIvw4xJfZBm/JHet6uHhWHhzNAjJ0cekVxX
Jnf/z5HhNUOxXTaUw9/IxiYAJZ958Ft9HWybYy8tmgAcsYnOxUzF8AzuDASHrHYm
kGycF/fiOdCj5A/xL0fW1YWibFNaxa7ORbfzhmJkklKmRFNfuRC+oXlVgTnJya+q
nypvVC9PV7+NjhV52Br6B4wQU0XKnJfVJlFuW7OCvOuWNhwYpNhR9tbrgDHh/0x+
aBmkS8bL4E9paEGD+ExLGZF4lL9ma1JZ3YA+/wTxRTxz+C36cF/zzEw6UKY1zH2y
6AzWhZ8+/PUO0vUyTkyffQIJT1VpdRas9Dt+Vk0aTjZNrcVaVD9tTmpJv5cjrmcT
9lFxcNSIBQKSjDaQIyjBQ0rH2jHymGrMl7JE2lHypL5YpilN7Ru8kurQTBWjIU1I
W+u5nO1ZVXpIvOpKyWIhjz6+eVnG0n8lMuolhEf9U/0dhBnKUk+pwkt6LT1U6YR7
w+ybnCCW63MYFSOVYNbQBgqsGPropyoXjSh/gYYBcHDE6Ci+Uvgu/RYqPazf5/qT
cl2Iovo0KvO17QhWlYOG+koUlWr+um/nn6ejZkOOA78DmWOhnBbfqv/P4oZb42/0
LOD5XHczc+DBakkERaNiKwKVRIW8vGClNJOYmpC32Asoe7QoPR+Vgg3E/M5S+36v
8lZqwe5XrYy+xssA4fxy/XJVvv31TiLXLvNV3XxOOPa168kWE4SZm3utoMKyZyo+
3VEmRyI03oDMvP070mWHvToGQ3jF8eb3pdWkfT2HiDn4ncYxUmvJYt+AbuzWXF/U
EL/hAm90+PgWyipEEnsQtQHP2TALlq9QbblaDY8DrQWvSGyb6PLmoRv9tomDZlwI
lQCAQo77Hdudt2eJhDCSurh2908Y1jsKPBfGpctdme/++RICxzQ2+Mr3Jm68rsHx
m6jcxjPlB60fu4/HrMWt6bHt9340aX2J95xYmO1zA4VA+kOxt6Qw7bGXJu3fE+Lz
MlBMsTyeJ57dId9Ajm/+7uaVtQp8qskm+lnKc4iRdPiUOr3iW9Q2i26jGnOIqFJ5
xrZKZib3cL0XsO0+zZFctMk6D4fIoM3xcZUZ7DRodVlJpOuWvRK0ANfflLdAoQGV
Szk2V4F8MaxDCOLGfuaifRVmVYFUfR/Vg7apE0MtNH4qpeNfGyJB16peqCDg/Zwh
g0aZpirA5UBv4RGAZOZ+sWWreLhtuJhlBH+Ww0v5WFMM5m7DoKlKR3vDSOGfH/GB
u1SlzMBN+qLA1gA57avTgVmxNyowNm2bDaIssRTmgV/Ih53o6LgXOtQxPCWd7oLj
1UlaEzYKSUWqU88Oep4Qa8derOGNIPPql5HKA/WWgDFh7TG3gfb/BDyGxPYtuDo2
TwS8IJQPA2hPj75NulT/AD7dGqKy2FgN8yLSL4ey6u35F56PlH361mJrgqg56PL9
IfjT31BS8a/yfHee5dJs5FsZuWTPdeQXogkbde7jGAbece+9PkB43pmc/ydjg4hp
rfAERC9kXAS1gJE5B0PsXoyKVlAQUCu/mEnsd0VKHD4WnvhfSHP+Gkrnocjn8OgU
3D6cdCa9Po/aLhNI10vZ50iS76uAAzOln/NCLmtTXNsVT85VF+8h0gtPCJF+5Rnr
9SZS9ZxyB2D4Vw/egfvs6L7L0IB5BdNg8g4uPJiVrLAktNjOPnFEsHYeLbp2LUly
G/FygJAAzvXcLClMHrA1jsTimubynLO3xwnucFlmqn+ryC+0pnFcB2SY/d3Awki7
oCjSQdg6OzS6L6Y4lHvmgYcpd244tTcgZFV9PfobZXfANOR9IEWhKC9SnmPUb604
uMd8/pQYlPFxprg85Y70I02fGpSbo8bX17zRp47AkFCR8Xs1z0lm3+HU0JHZfNeo
/qfGvG16fDOjYThSFowqv/+vBGKDQgi6XpyqWod5yIiPedL/f+BfLqmlrTx4FcSQ
fA++oM6hrYC6LkQoYDfzWs7gjZfM0siEwcq8mPon7YSPrDSCX6CrehH67RJ9jIoy
N/r3VgLun9HDXouj6jHtfRQn9LhWiRPBMdcWV3L+qAL+qQXczH4QUAxO2pcpsikB
Shw/m6y0aU8V/QTgLAgi0YxvcpdtgEUuzfoecF7P8KGZKodiqblBpS3CP2VieDzY
ppjG0P+9rpvCraNtX60VOQKT4J5X231ROAJVA0zSGgOZTaj5CQ7sX+UXSLTS30ri
oebJG2HeSiwMVYYG5zDRRqoB0A5lu2Zr9IzBuduEJGSuuAYeBxNCbJJUxp7m1th6
ZE6hu2vRARaY4nfzKjUWd2+aG7JqhuselvGqeXbKWn0KWGXX5V3oBUhn2Iw8iFew
MAMy8LWYFhN5AVUR9nd9viNK0Ynpf70+PKMjoEF8XEIYIzKO7FiTQvpaHTMvnhck
OqUna5MhJ8s8MZVLs8Ayo+wrALfSZKwIUKdjy+8gKoEC3VANSNnKZBeo5rqD7cGx
DctVmn2J4KeQPQUAxZk6H5e6yJNtBofonOK0KbSZ0OGV1EYoVMolOWuDamcRiyMx
NjGI3+RHc4jq2eus/9L13ahru3ccmHOhwjestyrxUOsO928JrfLqchs0DXbIfxmp
QTceGFW21BpVxxNzMZ7CDbZmIGK0pMV2Af9WOvvlo3AGjv4MhrVh+aSkNW+N/8qx
HAB5HIQkB53P4PwP4VVdB5UJf6Uzy4KE37Z3zEA8+qUgxWey2GBr7a720GE1qBS4
FsMjjo9EOQcBdEBDQPAYZKSpLB+POXcIiUKgzJ4dXZ7xUsrWdjjEVKs9g/rDgeNS
1zHCRpr5thG0wM0MLXncZzHWAgb3gFtSzu5DtYa8Rc3c21XK1zcyWXDmfIMrT988
aodJ/mfEIGQpI7YlnsV4mUTLNHZFdv3Jx2AK71vFSrKhERD2d/I5WW9zzxY+kuvV
aucwci4yk8HIoKIrVbG4g1avbVNRgm9kD1ilgXoCYF3Gb9wz3vQb+mrZdmDszkrv
FsKWf39V69BNf/0u9vMOXFNDZGiLdbb7mmXaDOH+jGwKa7w04pRTxTGKSo9NFYes
HVGwKmGlWNCWSoc6sq830ArfaY+fq1CUlXwT1dW90ikU1vBZ26yF/DZHhYFBRSlr
rbQ4EYUCQLkiW2hZ2CYDLn4Pepalt78viI2Y3EiTRNvz39AGY4yzjOXIPuXA2ZaX
HKmhTiiZcpsWzAzK+Ak5Q+v/W8e1qwt0uhzpP4lo+SuBrXu3nlfC34yu30kMc4zz
IaH185nkoUKJa7/hnyWTsHkdkewjDGYmq9tOgTq+5az/m6G2lr3LIHdYGE934YJn
Qz6xoKnqZEbIF5vsAs4FQ59feljJPbdCLJsD9R2kRcqyBst5n9MdiRR72Ta2kV8B
+lBRr7UFpV0EVCs5CQ2AuUGeWcMtADs+Yugt9VGROBHeVtb5bzLmffD0ClzU8tKl
YuA3MfXwrfaYJohyMNnANDqnpzVKIWAVqrg7ILy3r07TCEBBtijcT9KMIlIi/DDv
0HhD6KAVJQMc2gnjLHco/wrwjTkKZmSwMh6AGUoI8kDQq3q1NT4fzBad4dicwEYt
P8Odsb/YOWs8D+bz6R6jlmnFbMRJOTJgE9vmmcinvFinPR+ftC8NcRPMAU5Sw35I
JI4dol2E3JqD5QtbnbkJDIS39xE9Xa0VrNWCHSyjxFWUm0YC69iD5/br/42UlN+c
yTQF6ZvGW9M9i7OpOo+ul7D10kaFObqOubOgVKwrJKhoziW9aDR8ITi4EispmTYb
kg7qXgqNz4BqzwHR5F3pCPLlntVgj3O/AgRhzLw8+xPn5NBuDiAcDh8z1QdYjN8Q
FpjvUpnRolOwJzMTLkt5B9CyLsBbeq9vx+hEjxQsP5ZVxZG7waGRGESSBhINbWNu
P+G0KuSZYsVl+lni/+YQllvL0W6F3Wi1m57iQe4EfTyY0Cz4HEkF9MvL/56aw5C3
tfMiflwLpeWB7mCkBUBumqPOdARmdmN2RC96MCoOQwEPwSGHewnC8wdGI/HrJJfD
i4GxGCsfAAljvFcxvXlsngkM79PtR70DNWHsbtlcgoBNgsUm9IIhy/n760Tir4sc
OpV62esjetIcyhoIXWS+9gjB6+jyB51ZkL3qNp/0qVEWC0Fa2+npxvfeVtc5/zrZ
OiB3/EnpnPmqb7ILrTb/N79uUmuQv6vBgruImSOUbQKhM4RAnTVVmVjqlhY6SSbT
lBQk5dPlEVrRwbYJitmlLcrOOspqQ+4PzKoFX+MYeXC3DtSS02wMWJLTEhDS8Uc9
vyz354vd9YfStvFb0HVAjeBzBvN8zyr63iHbMtuOkKA/S+/twY1kiISV8zuZr0wb
Qn9xDV2VEPEN4Xp25AekD2NwrSYs0gwy5wbj/KWj4KBhQr2vFBHOiESn/TWsFACq
ioNAfXajXftnBAgn/VJRtQ2D1qo6a0PSRO4D9FJ1ekvDRIXB7V9PGTh8lOue19pd
Lv73+zCkyFdibiEjCTjDKTA75av1cE4wMt0Yi7G328qUvzxjiWKzkIZExMjbMW80
LZGaZGL/5ARMB2SoYJUJAAGgwgM4nPJPUoJz9/2bHlrZm8UYfDsraZv6w5T3+cZt
1saYB+avZWHFGgxZZXWvsWM8kSG0iGnR7ScrU3KnJlwEZZeTgTT4b1XytiTnbHe3
pk0RiEq5y0Cu2JXl3WGJrFFJu+elJP7eACZ2p/JeqWKU2aFtYgyKvjNamiOauP/8
RK9pU4XWL6m0DMVmx6rGZexsGEsQG90dB0+4Rt8Hpsb0fAGtIzOGqV/yMibwFXsg
mqNGOtqN0WgdAbtnmHvlCAEG1lxfS2K3ugy0qWwr1V26BND940BwJ3vcn/FtOsIA
OIW9i9hZFYoE4yqbgwedFw7Cdf9z+UP1Q+itbZ/TLvPHVmDr1VjWDiVYrGFccq6l
NhJvZVkHIXa8F2exH692yql5qch+pq/qusJ0LPoWSrc1ELUtB0Cbqv67C5qt37jg
jgtTsNRqeJ/gjMGvRxoICBTi5PJ7hTMckkUE3jDECaMG7xuPQ9ocOyr1os2y0VK5
mGJ89zQkgohFe5CwJ+nwPhC4v5kzVUBfwFjKrq/+W7BVSp2FKnMtwRg6NrOhTuan
DwwjJVXN7oGkIZc1V6/e+P/yjqCnHKDvNHrrRk+JJkUN7JRQFU8+C79b2AsRvYEI
IXu9yCdmdOphPk7B9tgKJHPakjlezQvcP3Zq1BMUeZSTzQDLf3Zvz5/MUrBl5XTa
bi/+yPF01BTNNlr2MgzoBpX1+ZHoo3nYNT3sKEmb9H0GIApdjkFnCssgf17Edc65
SoCIPSD6kvYy88vHBGBxumtXlZdlxaotlYjGeCVlbPIBuKiYHEhTMwWtxbRdt3FJ
MlEdZMQritXiRkLis6ktk5osPg4X57slEVx/rN4/zVAqLWEdt9YdxP0H3loZYfno
iTnW5JOWfDO9VcwehJ5fbescvS5kKesnxQIMT+Yp5JS3Qw3dn6in4uE0LVnJlf+N
ko0PZrRDZH7M2rPF0hLPpUv2lw/9EQ744BbaH0EiZnU6biwUqm3lavmuHeouRc/V
0B1myvNRdSVHnfp1loGws/CL7Ae/rP3/1H4gx8MZkkvx/6sB4RQXLbUrl4I5hsCP
b4aWnPqF8e6sifJVbtA0j+Vzh5O4A3lNJWxoGC/dMlyNDZTzQ+R1d/E9Z2u4BKzX
t2APhbd4B7YFyfD6Gk6XOmnKs7+UH7qJ1lVnpstGNe/llmOwl2AzEACaR8pIezAk
RQnAm/yw70UlXkyaH9i69dUBVDMpMEwnH+dn6ySAv8WbhtK+bZbiLfaTH+t9KkH9
XmUX6k5ugC/j+mof6RjG1/NSPmy8OT84HQOyvSMQkChDCgHZVCvx2NdzLSUV0I2v
JJlEppW94fFVRCk1qCjXP/YU27cc5zLMGmItSW1Wc15P76AxqWZbZTPJd+twh8Mt
of0p9E7NuHBtro5wgVrLGzuB+FiM/CrQtxv3dJh/YYDUOUEzPtvAtQ3lrRsA7j+I
jwNalQ8FiVBJN46Jkx2aK5ZY9cWiTFJDR+VXA96Zb31qDy3865hKPFaY6nN32zIo
KHKlmWaG9LNOyh8ShIrxMHXf8jrY8M9fgvz3mqbcO27PlFxPnlS4BHMYRUiR9uS2
rSikbZRr0H4hwWJa9Uyog7qWzsIJVsFoyXYGgY8CSrOV1nmiSAwQ6EoOAKHoW0Lp
sDuyGE1CB5PLCsLvqMcD8yHZ5umvzLHD07VnA/CsHYiW0rkm8x5jVLaMmkQGNQDS
UkwfIXf7CqwcLFfdsHSwkB4ZuBb65OvzBzYhM68nn+Fcbpuenkl4BXH6XPC5gEHc
KiPzbS43At4T3v025v9rZRz4bGoC8ccM6MiT9oM006jCti/H7Eio9trDIk0IBU15
jpz+t2cXRW6W0RNHZ/iIGZGH2hjkCCsYj5bauHxmNEIlxxU6KA8C0Q8CvvB8qMfl
tVVaucC39gClOuiGWhEMrEiCLUlxM/sF/cdpJdiOyKkzNr7nOVbBsRFTbr9PKpI9
iKWQH/YE5unVluvKtWV1eSViiDai3u19HyeohoVQ2HNkt0krHEYhJCbW3RB/fPES
LdNznozcB/2Zpfmi8deraQF8Q+/y9UAJvhi7YgbPkCmnlzf91zO6GDcfAj9feeX1
zFc9id5wNT5uw/sJ6zOkJrWYiQD9orv4qSlCzp9H2KHp/hM4T1FALCWu9eYrV8Au
hITvvfEVogYd9fSO3ge1tZm4wKN9XfW8cgX0l0LVqm+KnGfQbR3IPf8D1QuueATb
zVhHbb7flW4Ho66dkC+h0PZuT9g+rfYNx1FS8D7gnLp6E0nI3ehXwTM/gJzTINM+
e8WoliKFKDzx+HUT/Ewlar18Q1I0GxZhIBPZ01Fy0GOswSvlBrivqx5EI9+fakc9
bUa6zIv2aa00WhTQmcWLBVNFDS42KSo9T0dNCBi9b4pGSJSeQv1nhc1DNt5M9+yY
qtXgq6l7O25aXgU0vJjh5DBlrZJjJwroB3G1rhI1S8uEI0DrapD8yOOB87On+6Q3
vqZyDMWyrJxraygsTB8H2KfxKKUAyrdn+/OVisWsBAqvlQKPEPvby4lHJf+Zdg2j
UM58dCQ+1cv/DMe8PXM30SFNFTDU5Aa8vRr5aFhjTsRcvKFFuiGiHvFBVWXH1FzG
5prHvuYORcz+nBkdG761WTcmVb1mD7YDqwnVu97gqDL7IjzIS8xhJQdQAbyOT5RV
rqkr7Otf7pZnIRRnWBg6BV4JaBmwCD9ijit8+XdUwvkXtovdRO6Wj14z8FxPHtQE
SwdriJhCxCE5ke6JxdMVlAOymeMxDwNPaSk0k043sY+DFA9VLi7fPOQzMph8O13e
zo1z+kdkg7PUpG/apr8c23/EbW/GQzq8P0c0ASKoaGOmo3MQW+pCeOgNWqrEPsik
rOWxWOxFLiOtaumKA4afV5q7b3Hm+z/rPaykw+i6MynHjyML8MvJhUATQj9C8gFC
Hv4vfFfEUyFoKmldeofBao3IBjllZNWlEmyEB0r5Z6ONgLKk4IoS97fBOjMiBr6m
mWOke5B9CzSJhDo3ZbQBfdoGZNT4/m5mMSwDjUv8p/rZrxPvMVHcCbrgpTRtHPB7
PXKK6MdT0e+nmE5itrhirzuKL4PgRb5RoJJBx8ZT2hsenhiIgFvHl6vaaxS74WgA
6DB/BcylT1aqu69hcCKB9npicowrupOs+lDIdzDl1HHZ61c2ml8Ijr2b+qbENO6E
G2/7Um8SMU6ZhjepxKqtsg==
`protect END_PROTECTED
