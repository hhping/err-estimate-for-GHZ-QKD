`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cKHGNbGYzdmGOE2HsM1MJbeE89Ys/4HhM/MvDPgazQjao7w0p/hjk1ULOjMeHdYq
CjQ+uu4OjnSd/ijJXf3UKEaX79sW+VJy+VySq/ljw3KMPsd2LtMt8zmpHLDmM4Jy
+9HfAOphuuLaHplaOoIRQTnH0Qg9FU1rHj60cfwpYbSSbYD+W9ps/S8o9TlneVKC
ckA4y5n3Kr6Sw0WiXzxam0z9NoSRLyn+xwAmVeZRLMBsF2z0z+wmjYHr64pNZRv/
XTLef7K+Y7BySCHSmoUvauBQURZkpXoILYla0b8Bvl6K33VSa3GrCbNh+RgdbwH5
4pJ8EeXDMA+sWcK9azgiV4YzENJ/m3DQJuo/A0e8U2T+X+xvGhL4mXUOnWSu5GrI
FoWqYMSZUdxBgqPbI5luN3PRnVp1Qe6Usw99L74HlijzI441s//mZ5F/fO7yFsQ5
4mVvK95UvUYP3xbr260fRNYlSbfFQn+aLj1MPvbmKAkTMa3KxMeF4WafjJITQRuT
M46peI/k5mwaCnyWYjpTFwDvYvBiW8NMA9DcDsfypWdbBQo1xeZTBP8o8XTeFk1m
MMjHlT3DQGOrCJvQfP9tyqT/HUyDg9nDZigeEULeM1ac58jrJt4IOxwahe/1JTxX
R45UY+uVSgMHv6KuhIAvwa7yEsdPsN7iIC+ZXdP22bFJ6bdNVBh7co9nlGw6DScf
ItbhevgFuRGmiwmdmDrz8T91/kKvV3xYVF13cAaKcltqmwcKCMbLs7GGKeE8DklL
iAOg8WZkts+SWXJut05aflDQvpdTnEy2MIzOli8soSeR1NIOmCzgbTHvhX1zqSbr
Fgule1KjF4mC55M/Y0ncE9QAMOI7HAuZGr3HZLA1+h7dQRsCdOaga/55ojjJCtzV
bOe9k4YbPOCeXGCqNIUU3qu8RWEquS15MGmqpG5jRGXDKHhCR/7xDCXOwCeUihZp
UhNoBu2SmNXPaiFJ3AbH+BaMQEhyL6sjk2Rpi60kyyV2qyFrUSOqbsODKun0pdNF
tAGhLlVm3qlNw0kahLiIqBe+IwE/KCh9yfS/PuLp18NmSMRTM4K0MGJo1YcRIEcF
uxIFGsVRlJXx0xYs9G+EN4HeEVkDT8uSSyJp9mYkGUmNvffSgzBIiVNpKJDn4kGe
vxMjqOa1hATbpt53BCVWgUW/1qAXpQFDWKGGFSt1TiL6TWSk/GWAkSnBIziEgzT8
Y9GZ1i11ypW4B6myrQqjMstLdawdZufyXFN625Yb8cO1Y9W2DxbnXgyosj4qkWCi
KNXiYE1WZR43nmqD1ECu9m/3LoELiGysFgETiLXxfx7zpolirZSac2MnAxfiByoG
CkqylPMZtwbmoBjlFpwN6fzPtnK4WixzSkQQkIs6rpZtjsMgnJYDThdpf4amXTgc
8IjRqqZzEPbWMyZaGUJ8Wwh+pgZMf213qOuSKKMdOJ57BpQba+6HoBbOM//6uNRB
vfp9prWWOmNHxlscO1OUy75TX9SDBYBoxwlubvJmnBGv5ZWBknmijL9WD7KX+g5t
XjW+1LxEJdUYgifn082J3We9ryrOJvRejeLDzTSoaNIdUjQPXdkzT0sHyzXNxScd
uYEGZ2Ml1TKEJ3nyRK18fxlJXRhOoZAFYyv9wZkmesxwI9ZCK21N/3wmTebjdvF5
wrDDWzCqRO+qnPFZAEnUn16xZYUYDhQhSEe6ipxOaU1ivrhvE/7KDfrVgaMAWxAJ
0Q47asdO6qtcBMIGA3jiFPzwZH/BjZC31QHyNW+iQ86F0J13WA9ZycwkxM5q9rVe
AZCbev0dnvUXbwKhbwfg/M0mW7Z/RaQ9rPV2vhvyUlyP8EsxpRHqJcB2OQ2k5+ng
jBk7o4R9Vp3cq3lA+efGNOYUbXcASBO2BlrKe/5ABadtKdNp3aVn3SsEejasxUjD
i4ogEWxs1kB9JZYgltMnV6wOR5rHUlla3WKDT3GVsvY8/Pqnj4CWhzWbmNgaG2XF
v5VekKujvR4F1fva5puSs7mPv9qQUpz2gQiSmyPRTuxrgLbDnModPJJuJ6s7IC0B
DcPelxXb/ppJDM3RYzrRzh8cgGMtMzV9vOwryrstZ/NA5CRCmKZrIZ8DMtlsY4RP
+SKJm4iERJQuGgk5J31CDI45ZGaypo3+IjU31vEg7guOg93doMC3qRA1B0hwSCin
JGA0fKtziTk5of3phwfpdKsFPTJ8soCLDSI2Vvnux3/3OcpgIRMoT9R+z+9xthhR
7lkMJU/zuPMjio7t4mybhN2vMeOeA1ejGbxsZpjU+fxsHK84T277BdDkjCOPjr5A
KiNoO+EKaHYJqKsQ03A/wED8KMwLXW1Hz6vM32tqNY+I49yJhQYEsQtD0TGe572+
C/2/QsTrn9aQuhLCoAh+biCVAju97oEAOzD37/3xvYZBwkeM0ySleNx5CG2GBikj
sZWQzlW2UztH11RazHNeMWBSKQAPPZTZiHFUaokpS1Z2ibhAU7btWi2bm1VDce0R
vZrwkO6mjGkxlCmmr7AK0a65QNgMcdHXURbtCAT6N5/zoCu+D/VBsxfFFVBf4nOV
nqak1GeKnw0BwdqpQyzq8CUzsRhfmsue2zFIem2kKwn8gD5VwdIcST1w49RlsfPZ
DG/rVHXqpaexAOjP434aC5Y5nloUXKo4TGkbgCF8ot0jBqcoGTW3loJKFun8lIpM
slhpuRWntDr1dNjhck6ogn4q6ljwQml5F9UzAJI49gbkq4Iis/BYYRt1ROa0MxGr
vT5ExTqhPW8NZL332olcfCcLnbmS9M7NTbUbZSxoUBSFVd5l0bSK5p7xNRlnFCbk
roe/okZX4HlVC8RsmpDjYcwr3rQzCupgAv8qc2RncZa4IvQTr5INsJ14zZSFovgY
qrePlup9Tty+MJw40ayB6DF3esEBh1eZzP7e2Jp2VFVG6wDj50hOE2/CaLhU6nf/
LDC7PM88xKosycqeeifXAf3DHi4IRybVPNaGZwqLbB4qrm4txcdVFwoEoPrliR8X
izDm7HfkebgsR24jFdBEkJLK9yjaR7uC5t3YbKT1S7qR4aOs53ohWNk4+hH2bmtd
CFKSEJmBOu9MzWI5SnSowzx4q6OnBlMn74fxsRBijjUmuJW8LArMH81dDbnNENQ6
TPtG5PBBOZCkN1QlITbnZdLu0WROGsOJzanqb0ogj3GGiPiTj+px4nKVbRoTX8Xf
teQInkItVfucZnn6rK40awbl7ePw2e5nvdHhcnAF03Vcl+Myo0qsdzql/YxmMBJS
UWiKbRtHCh55fHqZfS+nvg/AM4NYzqz/61Em7kSYNAYk6ooSKNVcJRBqE7yCVG8o
SV3u5NZYYnVLsu2XneGRNU74qIqbt1i6LqEvvWMklrRhSVhYQTQWW+ZCGnWKYftH
NxMkN7WHrmT7WuWTMNULMl+wRW0UVeoNkov3dJVkrHYTWiY7SxG+TFDpFGBFn+/S
K9PbfuClupkW3pvH2ZeePARpIhb6kcleyGlNIFGVHZedIi4K69gL+ZbOtEw1UT0V
jNJ43oE9yWbcxNHRHt2OvOHa1XWAM+VY5VZ00rYS7RwU5X2IPdszPXCls15zg6rZ
VwcT2tgaBZV+ZCBHXavhA3U3MgY4nTh5pIw/xmROTWfgPKq81KnhUICmK2hKBz8t
`protect END_PROTECTED
