`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P73D7/SEA1vad3Z7iXl+McbLVBnYUMODK/1Ny3gn/YB8Cp0vdqKC5Hlns2HfadjZ
ilEDDRhGZHjchC8k5JmD+gHKwh56hAtoEUzJhEn4uLxqWlccTpnxZYISPzdKOnzm
2VpxFcliV24xhvNcUu5DecmYSjDFPVYt7jIrpPYXALEp4gUaX66Qe48hEnxXlWd7
Xyq+Xiy+jh5kuDdMeVThu8LW5nhPyu6rf0uaOfzywP6zEbx4CqlsmN0U8EtWylFZ
Yn+90Qj06xMCTdfUyLJYlcpXrlXN3SG88GfGb1TWSYgNhpQgoe3/zGjSTUtqaB01
a7tnyjLH0gDpRqgJKVwvgU1GjQAF+hH3L5SgXXEx8ZP1ivdruwhBs8fCpsbRjS9U
sFlV9spIDa4xKml7F2NIkzNPIR0KESl7WCLS+i5C+27ig5TWMnWV1Z3DXU5xORUF
4YrwuVJMPgSZkuqClXzlOFbp7bU1mqYrX2okETOu2KNtxgyha8yoqCpE0S5pKpTB
jx9+LQbD1xR4NCNvLefzLiAWcy0XsGNKxiTlyysQv4UasU/wPM4k+yKD0uwxjZO2
RJ5h7ygdfYeaXNfONHLZvOnus8jDhQ4yCuxMK/bpQYGBWfIj6Y/HIJofuCgcUW+8
/twa1bLuAc5xvdQ5djJ250UdrOm3xCqg6FAaUNqua/DfAqq/jsqCgBNWCxh7gpcB
7qYaP8dhjno23xaqt4skzfKvM4cjhOqDW+wFZndFY7IxsPY8p09aoS6nuHO9I1AY
RUhWy/65EwHL8TgjRLeorePqpGDLfmqnXY24rw6+nERStghUo0M9OqIV+cKF0eKY
bhWZITIYM2BAw+HPRlpQpo0LLWSIyo5twi4SjPWVn4TjJCJHV90rGMA9oRihiv5Z
F/fkyRSPDVlimE1Rl99JV6GZTkvvtGJiOw7GaVbZgFjc8frbaeF7ySu4bFGJRcgk
2yH2vB6enFPadVMmgrg3sRS/KV0WJZkGZqOFOhJ68i1qooMlhkDqU6KeKD7BpI7x
FGpfZIM0qstNyNHQ0s7RAhidhUbldfPcKSWi6YiVsJ2SE7yAxoiRt9fQqZEoPUMT
`protect END_PROTECTED
