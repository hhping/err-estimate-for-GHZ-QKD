`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ImkbDrJBrGisGP6XSQhkOdiIAsZT/lm3nQysSf7rbxQr3KR61rPs/pmCTczN/AAU
Qe0do9M6DQnWEET6AlTHG1P0OZPOWv2G8tZ8OVPDPo6H+l3cTvs6VEm8XP841guw
iYXhZXL8t2MKEtc6kAi7dLrxS3kJ2uUdhKDbs21kdXvksACM+0yWwKGDF5xm7mzW
6s+wcj1C43W1/IFB8WWNuDn+kVhla/hhHyjq3FCig3XFlWi4TC/vfqO50NWNhnjR
A6TlB2MXwnedNUJRRn2QIVBH3HawuhSL/hlkLnIDpq4Ev/dQCVx8B8m/xrg6aBq3
3vH5g61VrLaasOAmeiI01ETg+NQpQmVnOBWo/7wHqgUdmYKkeuveDOyCxNkmg51R
jQZx14Y9w1lcfcF6ekhkAPB+LF7rLAlL1yuKS8PutrOrIQXSAeFnCZ6SdoLCLUBD
YoBEWyt+HfrlLkG6RzYeHB9SVZ2AamSmckLgyOu5wniFpmq7OZX+m/amH25pIdVw
+flQtEeL1Ms38JLnNqTKN800Wj0pNwZsq9jcRhvnlFQDqqOG6RBHvLA01NBDQnXh
9vj/3ZOjN2jfkfrfXazTUknwT9DDgfUjSdnrIY1TrqblPXfmK02fNFoqjILISkCF
5F7vHaWaEIVDdP3b8TBVy5kmxBZcPaVhfEaC8e9tZX0UYcZ3rC49ttvdQfuvbNCR
cpD2DEOuP26t8R8S3hU7OU3oX8kV8ijFHehM1/Mc/urTzdL19XiPAlnbxW6Hnfby
edLMEfRfBvmbn0tv1dW1Y7eZZKe14luhiSr8Ql0iWzPQMCWZhGpwSaghyEICJwOC
koKEd/MwRb36PsPS206n1i7sUumOEVzd/NBBMsQZ4thBqT9YAs1RchRZjT2k9U6V
O2t4GgdUqpflSRG5q0ErIOC7WcdJ0dl+hee6jV3Qxf2ZrnYT0Fc9n3F9Txv2mlJO
qu/5WZTASWEsCSV5NyGxX99FgW6NkdphurJqpNZc8ZHei714b2KJe6QhjU5g7ztd
0hzUMQkr8DdkQl2/ice9az7b3tMhW7cKLIBerAERMRYshNP3BW4ZySHw+bngQSWf
rF1y4ICbDC5+GNcW6PQ2ZTMshrlk1PrPsHZhQzAY6jufe/da/jAS+89EzsV2VSep
Adrap5AnUxTV38JeYvTyLpC1uiHrihmxfX6x9hFgmmojX18ND+Swjby7O7FtBIfN
vrXiaXqZijA7bzb2ynXCXN+DdXJ+tBzXGAQo1ficoXOQ3Uv6QRZh9IY1P9LPm0eS
0bpuMQ2kN8yg2MQ061C9aAoBXiklBDnrQNWMIdnSKOpnvnveXXMBrye9/9C3Puu7
BF5Gbl8brEdPimIRAwEl0epmkpvtevggrd+NU/lwhtEVqRq1BD/Agh1RUwxOQbRw
TS0uyDW6TrnsbMvuhxYHI3d7iqg7mNvDqIJC1gRltvMM/1sHOrclCcLcttVfRzGq
+fSnTtqSDNLupvxxAxPhalENQx0YBpzNfzCwGO++5AjWKtlZVEC7RpkRhpCbzBXP
xyDhEVHabINuMzn0Bb6G4w/R1SLV1k9li83/87+sIgCZ/o1aa2RnrCh4DvaGRdh9
X5YREPeXPepQpGa0+ze17FKlFAtnFdkPL4/JEpEdorbh3eclCcZYKLiN/TRxfr7g
dAIr03Uy/uY5nadZy05h3GwoCFsafDuTrZG/lJMfPOtGmpnJ+ofl4EGc/QCfr457
z64U9I8pSzYUEZcGvP4gtrmA0pedZuP7CFXd0LIWRslAQjzMeCStJPnjwTYRrPuB
yO/cCrmOAn2MBZlvnksIyDJYXye1kIGCXTHPoQl8ww11wfk6DfAxdJ/e2dZaABv0
pGHoDBxkTpOXP7eL1mDro/BO/i+4jUXvtdhjpBePzvOeQi8ZXK9oEpU4fTf58ryt
JdBbgnGgfoD8GUsR1vcKAQosa0Cp43HlKe81pOcuqPA6njZxE31OHvrwfLdLtaXp
Fnim/JiyPk4JkOhHjgQ2AUCYLgV4NyeTGDtoVv5/WVpYwEWNIHYKlf1uOwW+S2Qt
eL2CJuL8USEq8lV36RYP4y0nC2w59iSh8Q+tz6mI/JsAmzkXP++kSV278SECXneh
bimj/gd4igt9OG5WMGdbEuzB0kk6R7jgFqcOpz8XEmSc7a4eqUhTZ957hg9ViiVH
Bgf1NvyRWRWs6MC0fQayb95JYlKwQwHk4IN6vT9984EAHzTGWL3gbKMvsEthtA9M
W55/zgJP1coueaVBVwFzbWqKQe0aQyRZh2pis8gY25RhZEbyaRSBgmtQhxABGgqy
aJlDJP0CVqv34sTVo1wJ3oHaFuJX8a8to/zIRCKu64p29O4k26tfF8JRD/mzvCWz
ZSlZjCCPfia7NjwmcsdzxO7ZlJg2dUWLOnl0a9Rl/BitblJf/5q8Lr5eKNzXMJW6
TrvkOhschPdcPh7gMO892m5KfVY+CxmqpYR42saZO2TjmpkVHnsxy4rBmSMLUKUe
GmCTPJfMX6tXdABCnXzXetBGs87+67/TMt9iIm+lLQSeOhLZPGoLnhCuoe5OYxAM
ItAU1L36Z2ecjWSnVGxt0Kpn8Gh4SCizL4DyhP+YI9Qdi0fmNJxWvKnZEAn3OMDN
5HjjZnB/bieEEH5M6tSxlHO+H644BYxOYOj8xieeoepZY5FDjmN4SvodllBHk1RM
E/bRWxJZ9B/y86sfUUjxCTKrG5MaH1e/a1dZBeqYG4oXI3cCXa583f77p7q88pXw
noD1JLGMbS6NrAtybD54mDvxGqM9V7GvSf9QBa/i+P0WsxcJXhnEE7yPcpWuwbHy
+1mqXdT6lfcj38s0xL+XfbwrSie56/8kc1/6ZUgACe+lxl/epd5GbZ02c27UNuW9
0fyT6KW7qyO1qL6vYjaAbXuh6cG7oDIE4RUYgMBJWDFjfcBq6bIA2fvtE+liCcxu
56F7KHFlzqKeu1PApD44u4zYJ779i5hX0vA+jt4QhTxqCJOw/h1bSlcWK5XNJyg8
KJI8BRjUI23C2J6ikJwRCbznAOePI+3q25xxMikk6CK8LBUcrXLXxS3EfvvdoWa7
CQ63gftUqZFNyWY1CJ4seCkMZMt3UXhPj2P0j3BeewNkzXlhw0Tn2uOPtvOnE+Qp
+kxUWjjrpUarAFb8lRZwpZr2nh2mbBTiQYy/m7sV0SgRfG+s0DXTxO0WLX9+FdW4
t0y79Uc6w/1p3e7JRoaDicjM/cP2Zeg0vv8VKcrB3P0jDvJ4Ag2LrXDtucYLPStI
Hs49j4ELX2iEWc9bsrOvqg==
`protect END_PROTECTED
