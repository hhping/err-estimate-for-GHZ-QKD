`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8TOU3wO7G8uTQGHva9xuYfCo37xvyg4hUpry0KD1XoalVm3DK+SN7T7/LFJW0cI
6F0hlQO1nP/i1HSLfTR4dk4FfAfdE5xRA/dzvzxmQy293q+wDv87P5yQu+J7eaJO
juOHv1soI1I36hsk30PHInzuk7N2ObnyKb0qibIDwzRbfVLbZhT3rfK17rXDJI/G
SVGafEJw5EPAvZ0cVJw7gEy8shs8zYUmRyTUm7naoDwrGSwUKZlBM028nj6dZtrF
l1sd6ga7VA27bGr9O5ZgEPNHV/ozjk/CSl44RO+EVYhFEG4E+ZNSR2xnUYTuv2sd
5bqM2Z9MAFsLEFhsIQtvpwzCMPZg0VFTD+D/2Qs2jHzUW/IVnAPdGr4r2M+FeEfh
EpNZmUEvC+GF84LZ/COje8ePui4qUmjtGJgUWLQF2nZKpTQytOrQ8JP7RhsRvjrR
04ohM792YgTDDpCYq4rPLFbX6aEcIATQuDx5ZAOlRVQdCROkBNVxdjjjeN1c7Vfl
USOn+7HRm0CFAA+lDn+02i7oL+0uuOVArpTqxjreYZarbvMIrXFg8oMJNDQOtxnB
zsNTb/jG3U3vkgoswigdJ+lxeUZicR5zQ3Tqv3IKKJyHKq6NU2WztX1OJgDb1BJ0
9yqrcC9kp1sY8GCdgYBj3n6Rfgs0f6GrN+SnW7wgQ5gvAErI1iAy7imelA46nGVU
G/7ub5wkGfGfzEfWVyzbgnFv1CSTmDQLWDCVtCnoaL8cvpGnWxRh2cSGhjYlN/ik
LkbjBdEoH4LA8Koni/hIC8fLgitq81xk9bkDMnktz75hf3e8SeAXVJtQGgUL0A2T
sOfxVffqKpQMmqGs0xgbBLVIqWrAOsa4mWgnaz3biDbdG3FO+XCamC7SFqj3L+FO
9h0rucDzY0laRCy/WvsbH36oNatvQFDvJ1pVo7jSrTKqgu41b82r+IOgM5cMBu9+
TZl1tqcYbTdhDKjvPaN87e9V0I5QA++bl+OqMc1F+vMAPT5I1gk6PVrYhtIWXXHz
kXyECuT4c9PwDYTiTlsYEi2WOMxXaT+oArLSLppwevdVpL2S1gXG78WsfLTmB70w
0y+7kmQKnBKO8JoC7De8MYa2giEsdhBOMbaQjzGO8JdYyTlxxM0/djeLhtQGaf+c
0rtmdsZfzz4iD8Fr7irJSIzJ6rDnezy2xRBFUSjvztPYl6TfysLfgjqaJT5e2A1f
04K9CKAb8XDog2ENqDny2+w4v2AVRp1+1ITi6P/dKcWIY1IkOJDretrjXKibBw6X
ErVnR72KosLcgba4LwieK6+h8KD3t5e+C2pTcAxik3oaehBCsB1t/5BdETRM+/EZ
cxCn26zjVSov66wvQmcBwos2QlYye5C/wwuF72+ml7V8BOVJbBjCp+xTLe/+w6Yg
Xiur4t8BNWoSpsJiRx/65ygwv9tCWzpA1NLcG2N1MGXsZ1Pxr28evjW4lcn57Zno
hI6ayaBMydYn3zLgL0LG3b3DG+ppwhsXUUkAR1XKaG9biLx5oqZdyafpJAmEQZNB
Z9rZH18PMA/XquoprGogt4yYBDYEJJ1UjvoKMV9BVSdFXgTkTsCkfVYIfm/G/RHl
Yq1nZ5FrEnQLTuHRj8umLgSVNYWk9DGp0JjanHzMfBOR+Glpe6HYTk8A3rwlbhrs
n4pY5wWUQm/VtP0jNMQOCN6SehNTjDvz7yfYt4LChN1cWXNgevYWj61j4EvFT6zU
oNIuIwlGj12Scv0MEIwYvVqBYGM5B7NtgjyJjX3HMyKqSzx2DKmkItJLAcXkHLX2
dyCQ89xO89E8dTboDxjxRD/Hw+2FsNYly4enjsnEpak+0LtLW/V+Vbahq2QAkXkw
S5hfJPRCMjW44YvZUwmgxmW2r++GA9t+CNDqPBXA2G/+fHxZvLJpiBcNQ5vwgh5U
gNflyC5EDpvNonuLGKlLCWETB4ljQCpITMG7EGkhICE1gMVA1MV6Hv8BtWwOCA+B
GE6vUJyE0Dv3qv4w9erVZc+C6jROKqqw6LjpRs1V3OeXdEOtkfImF5Fqd+cBRwvW
JsM+lmLFTCCh5/lJuVmNwlbMgVpAv+0qhM4SyERvhgPH9PAO8HNIzElLjZaoMEcE
g3j/6ClrjH2lVpFMFUTfYz6MriohxmRKkYlvNsYnjom5WYTSNX2MMdWXp9h4yezd
6fZ0i6w/7c60NxCWGcf1Zb+CfC+lwlVfSQ3MK4mFohiGM71qvEYAfUvIDLaBwdDW
yMtidcpj82tuucJnEum4WewZxHMMxj0Mzx1MRNbBHAi3kM+C6Y5x5rUts0mt6MO8
jmHpz6Yj4uHq9AqlPnuogyrdWTlVmDAN7HDH5KiD9vx6S2p7MRx7+pX1BSmqy1XF
bkUXqR2DI8X7imPX3ZKguQ63DwDQMj6y/oNkzQhfUBR3PdJjZgvpPNH4KJpsvKUE
QyqFKNFR+tdxzHJX+WSIcM2y0Y/imDb5Qp1Y4Zwd4jwe+rM9PysGccNfpYYWhvp2
Pl/G97bwJXzM0rPlGn+qRQ73aIfmrjlkGQCZm4x42QfnkckQ7FzyzWg8eKSTNlbl
PTamq5ecO5+IiX+X7Arh2koeaxxvsR+Y2criLm0AgpxQL5XkXgEggNhu6J3GEdzX
YXAPtn/Q5NDTKw39YPX99MIHNNjIE/Ssg0O9/vVwnpKcuipSCheyEEpKllZb1tCh
zMMg9Msl60jTtx1G7D5TepXVckpfuLnEh3Evr/CMwbFfdjvarMf1nIi036ZGI4Oq
2V2UVW3krAL5k/QSwvPPKC7UcMgT4x+FWAnbGzNWSRNpb8BdwcxXkxaNZaelNk7I
4YNSlC3El0iukNqfnSnrAhBTf1b4hsRzRtCwNjG6VTk0+XSlSUBFFBZy1msuzj/p
lOzGxpyATn4RkYizzOYQlB+zXric56dZVtZHh0pkGLXfurzJ9Goo66sevbf/abqH
zSIzLj9ybualyjLHAPErOfV6s+w4uDIoP2uVMXeTASKc5HRjlziNO5k+AU9cU4/l
qQKcqSTmcfeAoHkRe0hst4zw51cJTdLZwnaffdKLSMiRmoL5Dnh+t0OXsvbYENoL
V4yEsSBiTj0vFm3HSaVAXv9Tj6olRhuhhbI3b+YldvmT8nkyw3TOA0MtsAvv13Y9
maeClXHYR1ICMtyiwbmeRTfsu1FyDuZQe4eJFUdF4yITV0h2OWaTIyfSoeFW8g/W
vRuQ6VNxBeeLv0FpoM+XrdNreSPvMviwjTB6x3w5zgGW5gFYd1ckxLVqbgH/6kXJ
KZWQqu6LXQZu771Apq8b66tML7y7cUzcf3zsXzCnftRjpCk8SktR8VJFe4XiTenm
RDz50N6BwbZ4DlFrbhFpEDY90t/rBMKe+dmfNJLs0azOCCevTjqAxntKQdh8kfTu
CiD9uGGLGEVIFAZWC/svUq0/WgVD2RkTx6/lj0IAjoQ=
`protect END_PROTECTED
