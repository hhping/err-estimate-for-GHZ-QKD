`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DSib4l/pLEWFaNs2PhsZijzvAaTUcWAp/rTfKGF5RVfCXuuGM8K0Mf5vo0QOJ6KV
PIOW5VFsXf3y7ZZ32Nodd7yCuOx3D8Mj9/8gHqOTPz4fTm2uFZRdtXQbGShHFlgs
SbE8vi5YzxPiq2l7ne2WrEVu0winsXwrj3QUBArQUAkVo7CiSQPZpJyqWcn9enOG
rrBe7088aCPcOAPrNdz3RHWZ1sjf/2SGt08iV1md32mRypE9abyO0R6rKlDUv8MM
g3ksAjo1Q/ktcsnY2A9QmwhAzwBhm+AIr631j8uc1OxddQ06dZ6+exyqYT+UgowY
7Dyy7rg9PXKKr5+VcpGBC0MfaNGuN9GNocClemZ1Y7Fl6f1UH2gC5+GRAW6gc20w
CJ2Sqw9m6OVO0yShySaP6FbtfLRLu3jrRN6E2Fy6kdvRwwk3rJBPyCs8qIj5A0Cs
nqopCCsETprnD88XvJDYLCu0e/LeTeSKtu1YVNoQc4uRckq2WL/vTfTwzXiR8XZy
4V/clwOCjBimDIZX+G8Qegeq/BVqw154LH1Y3VIRWbluuEAF5IdhkHVf0fyV5gBD
YpNJ7goX+XMYUzLd2HKzsOGsKP8OUciBmjzN8RqAckfydbhc2rU560Dk5cZLebjk
RuTmrgWadRdfeN8t28KeXyM1bCQIqSdHLSNp6WVZriphYbVzV/gOqtSy9kigqHDF
uJmjRkRhMNtyo8m50ZYHniNqqUsLboZ/C2a7fb0hoCPmxiH3O4FNtLwdNlxnd0d4
e5J88s1TyPcy005936Yr0vAVsE7YM9yXppft3m6vzQAbbwzvMSMNdJcwtcPdMKmU
AKOnI6Ff+Dr+dlvSzYHdzBqPXHHjClzY4PzD5v8iqDX7V6EgpPx8/48fyTnX/cEH
/jUHnWp7VfSkNSk/uiCz2fS3q0owqml+QAG9xUE2GpayaNJDQAIOUrtDFjV16y8z
9bLgr41geekVfFbwevDrz0/WDqU9FCIK/KN4fgpvgG4YxtVR8a9jzZkVpJSQCVUq
2ySImnhzH34idvwezdRl/C+JyiNO6oVHQ3OTlkquPUIisaeS1SSPvhkPUY7aBVtt
GORKu14/ujCyzdTeo+PjM5od4b6zW4A6MOJ4zE0/h5wUVAi36BUwpLNwQ327z30U
KprOVB/xLZ/2U3asrBV33JAXIW0D+pZhyGx3UpNZI6fonkDos2fFKFabZ5M/rimM
QU3rX6j1mcbRqqYetHq9BwPfUItSIGRNTq57lC98/51hpkXyHU/6rgFq+eE+Y40H
CY9oyzrSiqtyjFiy4Y1OIhgiMvTmsg/b2DndqqCS3kiJEblkHpCoExHcqIj2q0TG
R2V4/xltf2QNMuQkWchPt2PFSGEiJRwGidIp9gLOQtu4/KKHPgKnmdEDDswNbUTq
eza28uwmIrXbzCFmkt4EOowVIUuLWR8uKSBcjiEpUr8R4VHH4VsynYjWSFJsm24d
L02WaZOTyBUiPZ61gL45DfIImVCcwqa+9tA6SthJgK5rVah0xAo84/d0qt0t3wXE
giAX2iGbU+pSM8tb1dlIRftfq/iC2pNarLllBVtPYmE=
`protect END_PROTECTED
