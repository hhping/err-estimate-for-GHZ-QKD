`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SGlmu8w3xhl7xdTTGF+VvtQ99ojXiHf2/qv2lsYLq6lfKzGlBoPi89rp/45iamff
JDNiCU35VqCxm4GWl6IM8HRTcm28M2Rb0Rh1wKuBFYT8WRxNPOWnjI4thF68sD5I
+O0OFLQ7d+RVyIrMsunJOzE3htfTw1N8sdf/IteR3uGiIuEvX3fIKE1R99y4LeJk
uysPIckIGY/v4rTBc0JotdN0PTiDoFJTEhaAVeTz1RQS69cNcBUXEZEuaXSYHRP6
L+HulVN2djVavJpPTiTqEdWp5nfHbFUvKbRoZrXeRrredA7kuSXTtllRT/eQHYAM
ETfn58Tu0lqgBSYYTLzz8XzoCMzb/JuRP4g6MmlPwlY24xWR0ZqWX/FpbtS+oxbV
wxhK76sceRnmIj7vCm9HLFW+R5ucqam7dN+0HFCHWLSxDvUya0bQPxsFXlLPK5U+
ULt9bQ7bFLogk6E25mfBZf5WhyEm3Kz7xLpczLTBiGnzYqw3cAXUOX/DEVTysLQE
shPwCWcB5rsrvpwQBoRwcCROt5O5GEnxdydshhRXw8gOPG/hmNaE8tAO4ChvqStL
BrO9ouvDXyrc2IIwqZFlvE96FcBaEeJsfPTDHUnu8CuMOj+k9D44KHTWq0by6Nr2
C+0991g1pZN1+0XxXh6kP6eI6pZwZJBm+PxPseSdidqXPvlfiHjF92FwPAOQ8JfO
+qjQsWkPx4aK9UlibsJeNVXgDtWp6zPFkT5UWHCGwJ4Y7IhFPuOo1XDwWpYXEBKJ
6NbSYLcxpF5TOXXbf32/l9i9D0Zh7ye62vwc5DVdOyhlB9diFpJOlCyLzOlc+x/c
eu+h2R0+LwUKdhl6NgxHfLYP+Nr6d/XxN1GiZw82U2vMcZk+pEym2TOam7M80mAL
SKmzFA5zPn4p/InBzSj3xulKcHbErMJPlZp04e/68xaZxG2yoaB4A9tM52bVFwtj
Lt+jweArhLyg1A1Tx1x0Ex//SfBZGaEZInG47QasLaA=
`protect END_PROTECTED
