`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
80HHuhDSGRcJLrbDO7wd5BT0TyGncZfwUl7+2kTfG2C9C6gZAPnQh1R2yWjBcUiP
ltFVhEf9H0l16LpSS4SMjsnEnCkipcue0i671ok5Y881WviZ6XKb5ddxZzo9t88R
HZjFyHBAH9zJ7An0DFtb3UQRVp1ZNgyncO+C4g24RiTuW9AIL+AK/Ml3MxjW1jAS
dAXklBYeWbVm81LL10qZ+IMZzOQaaQqIk0yG7pPABt1AdTtrg3pnycHeaSASbexp
Cyse41tma85gKSHs67lTmF0WOA3vyvOZpaJsqbt1r1YSVzu49N6qz6dIynWz8ZWI
UWskuvZJhaNwr4cUJUKcbUhTmyLBh6bWD+7gTT1Nv+8l6g2HsQemdAj8jLH1Ngvk
4qBzGuatbIY3UHxLXuC6u2O6FhWvghgWomUKopoWJCK9DW5TMvM6r60J6bPGwcoI
iTlEcbVHKjbWHBv1FG11tTeUMzK32R4EMGIJpiFNXkYualhs1A+7px/RZwArNYyt
K9eQ/7jfmW+qetVS8ErTRrzrApM1W/x/udHrNX3biMWWtpMx4Mpb+CA58INEtx7/
G0fInDy/1844FyPzH7fpXQy1Jl59u87Rr/tTLzWmG/110cj70mfrwH0y4FHpT7mn
2Ys924CiF6viQkyIZA6N8l42ZKpvx1ba0WUodc3o/Q3PTnimUBaCg8DersGElfjr
Qg2J8xf6fdLyv4diMz7JgkNCca0ZlrB/xeuDXaCxHp5SWagmt6c3nzvpC0l4J6NP
lwcDZfnCDYSj6Ulg5wB3KAM1BLSS4O/4BOTuvYOhJO8Yauq9fC59d3jYGZjnJyru
/YFb4H8NwyPRJBE3rDd0rg1j6VwqYMegvpP8FwN+sSN6b2X5KnS1AYSR4X1f7mqB
bBhlnbIQsXixR6IoJp76kQAN1WjBEXfy726Yd3xJx4EZCLle60V53pRPiweARil4
KmaBBGR42yBLduaVdpDSBQvANNjILEzn+0w/7tNzWAGQY4q8ogwFXQV4sHGR11Ao
JyJc9qc8QLUHWngL6taq7Yi55bsVVPSvKfs2Lgg4r02GD7zNrmr17d1taomumMpl
8V6U6awsBfFCeKwGNwU62A==
`protect END_PROTECTED
