`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XrtNBKOiGZ7Ch+yz5UIneS9Vn31ymsisminHXGaS4LlU/A2lnUdCtxIoI2j++sF
r2UNpqUFskieUO6BXdlyngKJl1hfGsZ9nJQA7iivZH/zaRZOxbDThD2QSvzMm5L9
KQydQlhF8fFtVafQhIY6oFpqQoseKyVf99qhAQLt6aHWavnajFYHfiYkKW/k2BsG
ie7RFZ7+nQ2spxo5/b1+Ui5BG5hqgfUopxj1MtIs/7F7IHUb5L4AXBiQbZgX+Hdi
V0gkc1PmkyD8y8EzuuFix0D9oEMJxWPMWVYxITwumJhN1OqbucU8o/ufFDE3OJPK
iLBvYPToyoOeTpVTLALMvItDJWQg8rpt/AedhXVd7kqPJ3nmry40jrUHZc1Asc6S
MF0/MtR0yYhOhpmm5Aq4lTaazh4QQC2XrOqMIXNHkPXP9V+Q2DXC4CsAKR2hY786
Bd930NyE6iSuEhaT/S6PgXS0d9gnJvVSYXC9pU9XkVi28ZsRLI95FclsO7ENnvYl
6hHdIZ1lfI4r/N9TTtwvQezyZMSkUn17YhPx1KQgf3ybYFmVtYhFzW3jfE55ck4A
Wzvvge8A7MvmuDvk8TyxaP1kEi6JMM8TvJsyNWebncS3IJq3Tdr2UdBQukXO0bUW
bC4WIKjo3FTrLZHNKSESPfCewZ/3TZlK/6cKFiL2ijWShPFeKayzAq1a1iwwceg3
iSYrlh31h0hm0rRRmBErSgn0UzOiJEEq/6zZ68LmSy+1s5MzsMw1u5qdDk8G8Sas
bEvXjCKGp5Euf9jGMtxkEbzZf1Pt2hF/I3NbfMRhj8rLaXYoLM7cxb2Tno2kUpzO
J0bnCRpYjpJ+kP0cI6xGvzaEwRsJvwebiqwdcLbmv+yv/XmCodntfJqx5kCkMwC0
AR+AyhkTiEmWIz8yvFRhmocTIeW0KS23M5L+J7d+E/Y+2opj2C7yKlMmdbX+A+m1
y/icVvCGIxHvuqqDjZBzkwciD/tGdVETsb6v5lnPemk2aX+kQpGsW11fegIFNyVI
pGACR0oWjbn42t0pMRb+qMI86AMwM+Q41mOXkfUjwQr/xHVcOQfOSWEBPkSbYV+D
bqEpfwZymGp3qRaXE7jrTSf12oaVRySLt6l1zXX4FH0rZpARyGxHvdBaI9u92D6K
w0UKSxPEc3KLQuey3iyOoPUswHyQFrlnAdAoAAkL3UiVBpp2zTWKPUs2H8pwAm1+
O5wfjoDzz5YUhQgRC+A8z2qh6qV5iOnUf4TCvbskkIgq1E4xvS/9+dDhHqmpoKR5
yGiLLzaSnXZyCHto4QBj3A1A/exBgxwO9+0k33UP4gag7cg9yZwXP+Xmw34HC48e
K8EVOdQe1gQKash7+EPWGyeMRfuunbEob1whWnrn45Tsl152xKHunHb26DYZQuFf
ClVB5GAubX4xm3snJSCKjgpNHDxrobTwQH5mn9cfG4s=
`protect END_PROTECTED
