`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvf1QvHWmmde7OdanoxpHh0KJJFvQI7ymRWRS0Ul0Lbx9dVev8HR1dMoUHGKkBZg
Da410JgIqr1tFv6WRG6r2nPQkgwwpt6wqUQt27AGsQsHey5WVJq5VyJdc/Un9KvE
1pLc3QCyyfpaLav5gniddpC8Ura5jKwVZcRf/RBvJJT/OronC4qudR03ojqiqcsO
frorAFYTNN78EDgg3zVwjFcwLZOjosyN35oUf0oN6+UsKcDTfXKwSbLhKYX5ogdi
oQu1NCx2tn+GBwTSLQmebaC5tAWhQs2Mm9dw9MPgZDTITvWaHDjvg5/+uHpppkRm
u1Ljja2VGKDqKCiVods9Cdr8K1Ynj2zoQFGP9YwFc0KVKFWq9JqAI5rtsp0O7sOO
mSr4khFGcvH2QTWvwVbfjV5w6l250i9rgHeBYySCi2+SSRjbNfUpsP89Z8crbQtc
nmcE/4S4bsdJyHLbsmUt2NLb5/m5ogj0xkclRbpxVMqMCtfoOw2fSbL4d6PCg/mj
82/mLC64a7Qvcl9I9xFjnGqC+hNrI1VxtUuBG8uFYZ8/mrfDSxzIqRfnUMA8gKJu
Wr27AyTFDfLngps/VCv3NNNQEttN33zTQFlA9Vx8LBFBWJaXqoWmKDii2rPS3dWG
q2Y3riQqGFMJQdBAnjbFS/V3IaGFG5nF4kINaA8XMedIfE48RYTknLzpDlQKJMiV
M5gWoAeJTwMGerxLjhVXWB2n7H+OmYZzBO/auUBAMkdZ04di92JOMrm09y7QMhJY
ijhgVoZoPzXriHYU14VGx5kE8Pmekeh0tHzft9gumhPVmy0jBCkRNeBdJsAWbIdf
2XNmZdaAGpXERL3P4tSGNq2nwoSMgxNjOvBmRFNAb9SGndNbdcyFSEPNZqUvLgUp
orwec/0w3LmZGPTWk0xBS8UdRgSbVhfFY28N+8bOenpnGzh9txpg33Ps5bOFGU+b
5ELY4WrfDEDsMYe1pper6OBQzN853Tz/kSdYOMM8X6Z7Meo7blaZmAWfS1PZisme
7YtIdSOnG2TaDzsHe+pCuregNB8+KOpuShPKW8XHnV8oSTwb0xUR8xiE6pmPUoDR
/5Loz+ZikpdzW7EEDUlSJP5Oor90zCLcitefv9qFaGlFFAYLBA8Nx6yvz6tUOc7b
4d+tmLyufCzAF9dtTxhWm0nv18LSBvhYwwgnEfqxsuT1yTJm5UHHhWexsazNBHIJ
WB2ll8B4ErN0lmV+wgAZxVfc6Y0odO7lR63F6mjW/MkOpXQAEeMqQ3TGkYuOWLJH
m2DiATf7n/n+1LD21jG4T7j+PzDFDA9QMI6wDOFZx8a21PeIYu28uDR4CwDqyyzr
JIMIZDeJUsxBrG9HXW+mGH/mZhMs5kHCmnpZGBvY3RIwRhG8RInUdHMSeYRAzFKC
wX8YOD+97D/RNfAitV2DUAubeV3u2pFHimibjVIcJbvRuSY2UjBDI3+Oi38LlXFf
00dSp51Kvm9XaysdwrAaSb1hGSzkhjvHMkmCmBs5TXIfdsRuFIUrGVeiYR6xANnp
kRHR09HdHcHjjZ11LujAHtWAjP7KLpdg6dKe6JOTNJt4+8RHAVwxYy4rhtQ5ppU1
GPi96tRUz46QBsUxasSU8Gou0K6985FRj7dOgYLk7ir9UqExxzb1VSZeC0EMWBTO
q3ggMRodvAYiaz7aIsh0OpbCWVfa88wyWMD2CsnmopnGt8Yt/j6uHTc51f48zfih
oPF8ViQIQGCkadS3nRDGhrehii9qONcidepue9EyiWj5gBAm7SwvdvCrek8OM/EJ
ukLg2CJW3YeH2bWRQWiKukRtOCCHJHPSNKC4veO9tke7OnUjbFxQ4wAfILXo2aa6
cHvexWM4kNJ9eyiAWULsLktxGwOFONolapTqIbm2W3ppwFMeX+Vv4/kRDIqdakdm
zDwMbkqoVGez/EcfWs58uGlqxhOWNFb2STmEJMvIpnkRQ9IA+qLbhJj09pnS4oxd
o7wJrnYWbLcoL6UdeXjLaoqOce1ifjXo95swuFQOxrIAAUgD8vQCsRgggiv90uf0
tthd+HZ/LRSgsVZi9gWCVM6WbgShbAbhxLalOdf8w5FNfRKYDKgb2jk+SnsMMz/l
`protect END_PROTECTED
