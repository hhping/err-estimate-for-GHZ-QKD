`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3WAb4+TNk8+t3SoBmxYtxOR3DbrmBiK6/4FjaqX5kXpYmztCU33dytKVvLCzrnv
P9wKOpuYiOI3y0R+K+iQxH0ecMW4bXsFCNtKaHpE7M+/rWfs5auoCmexCRj86roU
EtPNrMmMaTs1blttSGjc3WIPBtSsiRThVuFuuaDcak8+FSk+s0r9VdQaRY4ohKT5
TFH8YExtEf6+ptcLDhUTwRdZruE5NqBIoUYMQD4sZZZC65JOeU0wOeZJUkdJZLFa
Co1cEyKLMRunvq4XtYiB111opHKA6BY89XG/BiHi4x+ardOhr/wj/qD5C3/vUZtV
UwMwF5lqIXxz+LIVeBaRyR3C3fsSyQxT42bXF1I854vH/j2FaN+cdHMjC1q+wR5c
yf4nt5tLnQdRkRQ+GcKQWHR+yiDYLQ8Frq6lzGZwYK/QD0018VMIZ8LKTXd6cKK6
/BcBZB1bjcW7ZCqLyFJJWOEC32ozlt5d/XMPw9tAPwp/4wyYZbYW+gzHQpw/vhoa
77QDKay4OjVC6A85ux3gzaHP//e6QpugMXLHOaRS8rWigE3b6D04eu+/nVvW7AVN
Ycq0JlHNBSYfVGyzHOjdS6BArmfu9ZYxRVBFf5Amle48iipW+bUrJ8HKLiOy+5uW
s0qhnMCR1znlnHT6FshD9w+eWwXiBJPz0RehrtPw1rgFgWdgXNOFYuiyLqLEDNhd
F59pQvtC+OQN3G03cPZ05VPykIG1XgPeEU5NLNSq/8+I9jlXHImy7oL1DJceOxTz
YOQU1P5cKWYQfS5BpcC4Ut9KO9lFxI0qT1lxAmoDTBk6k9NTHwjDFja7U2kFCwri
ih1qweLqwZrv9KXkUM6rg1lA8CWagtXiNjFKP8XjGSlFQX93EysLXAHp15NEKGjW
mAL4JO5TImpVe0Tg5kUE685gxWIutamb2LQ5MPS6XTrd/LA5N7zaNBb/2tjkPKEX
o3XYoSWb1cEoZIAlp+UNT/uMdpMd9bFn8ccHIje84l8RkEXlH0eOT5KaYse//4FW
g8ehEcLwY1kOrQBHVDdpOlurR02SXxIFK5vwt535KlUGZF/8QHq7YJiSm/0qMDUZ
35CN9Kb63bT6iEPa+N4KoVErbd5McpYbbELp4I1G7X9boxvQWlSLFwrS+3tPUPIT
HR3qCALuZc3mwhefnljSrE7bg6ZepZdwj/jxgPQUy7zZj3XkxP0Wfu5/DZmQX0SQ
dI6TyhmLI9i23sAtYGA7aZV6V82udbarE4Auh7Ea0xBOw2ZMbEt02buQfBGXzcO5
kyMpSV14UaHecAxSDJvTxAVSdhi25uA4nTh5kBo3fWdXw2uZ1e7PKL9YKrGswWMV
x/xrNGDh8Uqk4ESudsZQLSJVGYvafuDF1KliSPfw38DHsAibbNJtOcCx+AsK2wnV
OrtrcGlZWpmGtwjjANwjsOJmyf8j/VsdhxSeyqZs+zqacg4VY8iuaO0YhAXIef5z
3Srbbea5PPKSnWihNbawvWLsrwaLhfSWPBIfGLfvGKnqARbmSvOGtMK1l9w4+flV
H+cktN5u9/cUrcFJnhZcIab68xIMAFlfPeFB7GKXeTJtJH06jRFRbdYIwHLj0pJf
6wseSgL7OIu77S2kWuascDdQ9J27H9KifAL/s52Gh4ZhZLi+HP3PXS4D+fK4VG+6
g48aopkMvQEqwhQDOMdg8zhWQ3vr/oySgcz7xyMPJ9Wj43DPlN1SK4N6uI1x1eph
6yaggnE/OS0ubqE3Hbs7Q5L9XFeGo+4d8Fce/7UCNADET6DzAxGxc0ut+nh2d6VU
ly6STODK3KiSPszFfNXfz1pLmLuiUoElmzs5LyziPrRk2QNg3vzJRMj3ajCAWSRw
+UueQZuEvQO8O48JZygl5GRj9hWbveTELcG3zIPud1m+qf6ViIF/xRPAyDDYVrKY
d9BE85HqwUlwYMtSeSfWTzqjVcUtsmujl3kWQSEg9YTVR3Agqpihx+7yLtQhWz1x
V1fHHdQOKDiM97Ckutfa2c/1PhYcslOzJZLuaJBXNhNpatfWbZbQEnCugjbyw6da
9nF0Gj4QSSsQJXAA5c7oPV/8qVIzLq4FWAmmZpReVRL8GWbiSPI6SuSL4Cc7oRF3
t4mM1iqel5/hwvcjKbsNHp1PnBMbp2nOS55NyXZ61aNJC34BDW+86oEElydRJ4fQ
Cm42kSmi+8bj5l3WTQQ0kdBIHfO9zSqtv2dIr9aGI/r+LoD+iXYwgF5+N1hkq7jR
H3FcwGZOvVr1AiK/uZlkCnxnMmWpEUIe/6jxyMvod+OCBaUKKCYZfhBoxtxnB76g
p6hBsEKF8cA1tCoUz0+Yh+mcAUuL896A3YEdjcHXmWyl+ee8/yIfprr+Gwo/F+CZ
YtLNA50/3bhpR1sa1Xs8YEAiD7Nl4huhn8S+6dXQrl5Q21n1k32jmanxrKkTPUjW
8OQAeD3nhCkZKNbqvT+YdmnhrJKldq4ay1JwN7PxATndfbWPnxYALNughod9Ihue
F6+SQgE5mR4NQ6CSA3Jerb3xM8Tyc3EITB0pVfzaNDuSUwUHXQBpe70mBebh5Hdm
Vv8hIdx1Zrlk00kPPAezf807jn+87cU76fQUlrGVb6iz4Cw+op2pvbbL9/jAlrow
5Ktntwtg3KAIBiHw9LqXX8w4qT4Kz/zK7Pag2OZgCY4ox4hltnzMKHpzq1dSHtmd
iqT1JDHe6moqb26Efkx1jj1UZNMQFj+IxJHUOLqE446Z0WSLsYrtIVKWiY5p7Xd7
KLt7LXK8lxQ9gUT6FFg01l9MWjD/hKDQ70Oc1ZrTcUVfiIyB2oeaGpbsIvI9lEVv
ZtyGcwQsOOrVMCHUMJkrNVK+CtXlAgmRZDW/AZuE9l6vb2GPmsq25cSq315UlW65
ZQtLDjaaPjyzdBje4pve2NkH1/3SgoUIBiUsHWNdC8c12FlWQjz8zwSNGV67NFZl
Q00ojtHKod6YKOz0jRiMAw5kcc+0gFaodnEiQImMfv9LBzEA0CihRWH2C+9BSs/9
KfAuN2Git13+hWbMj/ruQl5M20Erw0nPee48VRf5t7+PE1UC2hFHBD2O9Os7FlbS
`protect END_PROTECTED
