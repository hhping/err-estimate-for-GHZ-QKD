`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPbJgBRBs7uNVAiyuMDbyERULwNiCwWLVh71lvaSEDa2eqi6zwrYKG2DnZtbWgqt
xrJ2pVCMfBUrrrkWDqe/tVqWjQBjkN69plLMhg0Mo6UJwu4iaAGNOTQi1J46Plf8
2vgsZAQyvoBRgLx8Gn547poBcr0TfLGswiSAUOss5QsisquLA3R+jHipsAvQ+6vI
U0Fp3FKF3xHtQePS2bXDeqjifUmD+xxUXKTyAf/aREKCjhvyYUdezToRUbPymndb
JI116pIgaDVgxXVMHreL0XglVA0otJhEYCnWuJDJJQUYJxLiAyqbASmu1JcxXtL8
fIV7eH0ShiojJf4KbMngWm7nVgvaXb3KaSdMUFQSHyZXWdghE7Ms7camx8jUkqU0
SNVuYQ1NoyMMMXw5gKWWud5rOlPRuFZ8F/+uuPKdgzGXgVPzstqoIGdHEW7cRmUj
jksJRcrCXQZJ/5ojA6NNMnY5M8c0ZZgBL370zM196mEPkcTqc9Uz2T08W0Y/Yz/C
x9Bt6qKH8+3foyosw+nskU1RK1AmA83qIZ+L57MmuccyEH03UE86yWmxJsSjopNc
45x3IaEJ6Y/W3rll2vgR5VRHEanJciaOxibNhgqL0MzLPEPh0aGnwfGPv8U1C0Lu
jpQaLrunn0eAzssgM9Dx4YjP68A1BP/Lz/Uv1OhoX4nIZv1Qpx7QqxiCwY5XoN9c
3yS4/Ef5krfI5FUjr6ouFQ9ABsTDHfqMaPLq50dQxN9jNssPOWK4VSfFVg8y59D9
kQw4PkqpgsZh/R3rdRw7+FHbObmdwg2uKbVepC2z9yBZBy6X4G4NNU/3i6ComboA
6Z9i15yQUHIBOXE0wBlSCHrLkLNEgTE89ze1VMK1ykhBBESzfa25HvEDLlpr7mtg
cbZ3kylOFype72l6fIdFwpPytRMh8CHbxaAxt2F8NEFTdekt8cQyRWmZOTL84mvh
wL8ZR4odLsZzNkQ71Y7UWQEuxUJiK6RWJuqoRsIrq8tE+6MzEUrYxGGN0TEyjl4k
CUA14+gR1n3p0kkKeIjP1nWALgDW5lEGzH5T2g2lZsHSfavLufpLOkJ0coI4WfoE
O17l5z48vVTkpblNbQvHm4a0220gsGnr5lj0J1QYa9VlzwiT/ZlR8hutRzs6K9YP
9aVLSojEk+2umVI6EYGGCMxNNE59qspNqZeD0Z3201HJNAx7xUJFMNZI1hYKhHA/
`protect END_PROTECTED
