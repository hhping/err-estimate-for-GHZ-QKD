`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34Mi7QpfiR/wjUtTAGmn0YnqpFF6x5p+RkuD8eM/0UkYG+7fTU6OrRL0f5VVw8nO
BQocmz4PVILxCZBYOkUOWEwsvmcPhQbtMJA3yYZEwLk9bovx3GijcpJCBnFxdjQB
C8g+BTPNKEDmkzshtRb5taMkKKFn2IK+qhwnewQDL+RQoPjcQRMlxU/RTAtNe/dp
hloc93E/obxfDKG5s4dNxaQ2BH+Qbu5xLvwDBsNZf2zuLxudB/YcKIXebHbvsm8L
f6cKtir1tcMMY+cKAONuD++9sEalIpzKkaScuTyUL5Vr2z1tDWTUm+OEf+ZW45tS
dxgFs7NtmZOEe0seMrU7FxWkA5tu0qPbPFcNyD3Ymq8KsvxZ+NRVmDqUPW67YSN0
LZ2HbWz2Fr5DjvS/5tb2fEg8JoFF9ops0uhg2bV5JfEDZk4vdUyRYGQWdpjyT84/
44fHO4HtdK2jOvPGzWwheYKSvtmHfzf9JMEGp4JBYx4=
`protect END_PROTECTED
