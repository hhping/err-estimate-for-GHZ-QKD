`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZPyJCxIzpYUsnBMCwpSYyA6xsaEzYX3h69LFCCq+zhycUnu6AcTWk/3nSL0Smr5s
yq88UXgHjmsUveIWaHP55+BeWfZ0nsbAzcjA/DJGBebdEQwBuFnJAG+rU06MxDWQ
4SO/ftCVcElEFcV+H1Jo2x2EeZQC5EPMqoaQI3DieDot0gjVc/a0XMQL1+7P1rz0
SLu6V0JH9UJCzxs2aHRjie7WTcoLh9lQ5yQJmxS7o1Unb5+SfYGPOtTQajtK3EOk
UYdzp3woCD8PcW6q+5AdTcZwLtRtgw3SM2mV5YuWbVdFsNUPPUAbUq/IJJsMnrt5
Dxi5Tg0j2IfCUzgThTDAZcE0yJECDuJ0jGsqDFxI4tIPw7ZKLE4L7UK5qHBsZ5T1
MoMBU6kcCBNLWsADZ4oe0bx7Ye/DefbA9mgizgDlv3r+jaXPJymkSDuh/xr2+80W
C1xsrDHN5M7haFTnrnZDb1geaq1J8Zpf+IyzCB4Ddam9E4n3ObNPGRU9Z5YF0dTb
F7D362gkM3/XWFdMW7hcDTBIGy35pSJUuKH9wlLWb3pZACz1iwGLX8Ax00hbJj0U
ZtVWrAfemPH6cmbWTXwzxkpyhQIYNoRapDc3J5sz7VEOvn3LaghNaIzEoQ9FAEMW
57ehYPaHYC5GdT3O1bc3XHsARFRvTNUimopDYtcjYivb33h7Y6aVWyvoEtXKKGSp
7ziiHqn0Ht8ienWCk+sdkZX83pQ+JbOLr9SofHYhafWb+RNMuqLSXTu2NeD8tomx
ZW4oTOClQhZnzL7Nkz7FiI7SAzrcmi5nbKcjPwlEcmmJneE6m3Zdf/AhVcYPbh7O
qL+yeiANhmD2V48il+N1Sf5iQjqmdK1j4xGnVUUMK4p5wlVrIMKqtMK/D1Kr6JVZ
HHZK0UGzTIPNOnRT06i0QCvDU7M+MyR8anmQfMNBaT9QEGkE47EybsZ8whihU9QZ
6JAdC1BhRqIeEbgsaNQ4x2Zzzeb3DYDQq5uAswDX+bgOQ18bgHVXpmJ7wPvTvfTd
S6qeGclI3APkcJoTtCLv271kQniDrDZXzdQNFNvZEN/Biggp94791n+HC5CtBb4E
UTjKCorXsjvi9g3//9S5eUWbij59o8hWk0X0Oyv9rWph7vQZHRJUXTb9T4dMbris
YwQXy7X9g5hZ37MSBPC3Bfd6YW8VomorexP8iJzvjblL8oz2B3SdehVSHQP4GFTi
kUAL0/SAa0LD7+AWjkfDQHF2jF+f7FCTWj/fL2+wGxW60MDDR1JUNm8UmXPNtXNY
GtJXDr1D5seqlsSS9IjMLUy8o1Wx1wn5kEi+pk9Yhoepd1+m1ylltuYVEhE7zqAC
Idlbm0OgNwSd8OKbJ9cNzUwc41yvz3VAvA9gqROUMRGDTInvyyioml2s+YAwR004
ODeoPGNJraEtL3Bh6DPYMRFBDvsZuteE8HJdIdgcVm/3gYuVvw6VmAb+qWIOTfvz
yGzz47XOC7X8tBhi7Rj9Zm4N0fOoDulvq7wnj8V0JBK39iPkW7wlitF1NrSjdl1z
1diNtdFNgNRU3MXB7UeMRrZCvzhZc/qKEcU2VRQtPRw/IDaIgpdqCgyrHT/KRbIk
11yWsPRe8hw/Q2PZ1/TLPQWso9Qobnl8l7cTsUVZ2yABRl8wzklk76/Oue2MSZuM
ryNqMOGI1Ps7e3fQK/dzu7xmpqnceM48lq6ZVdqriovy7eixPPHRzejW6VEULj53
Gf2brm+ETkV096m8acYqZGwZ3pEZuBjq+LJ89GiO2jt+rUfQJ+aMZLf2hxLLrdM/
UvKuZmPbxvvb8I74Dz923VsY5wQllch/JD4wDh2WJTYRUh7tH/St5e9oAX86ZoPu
229eV3C0FIksGoYMKv759jTi515VS6IKNDOLfe+yGVKP0LyBeUTtMKeM6WQXozGM
gU7wIVAAFerxjedzxAdD5DDoDiU8723dU4u/dx1QIk+qn/0dDYYI8IYA3yRvvb8E
ccndeqcBdc3mBG4BN+ssPzFqgTZmlQpyx9cogdiQ14RJ0mmETSrG4rwutk8cCT50
T6ql/gZj5l4QaAIFCWeP/WKOMIcjRpCVlEPH4I0JYed7hXy1LCz+iF3/ZSXhFcR8
6kAzAtb93Gu31bNjU4f6JzMeID0sJS6GsZDjm+9hww1y0wzczx2BdT/cnfKUpiAj
J4jfkuPS5QTzoN65ljAYTxK24epyFM2/pUQe1U58WDgYnVtebqNo8kAI0BTgWKXF
RU1zwG1mIlQdLCYK1uFQSATRAGNJ0L+TcghnOj8wqkCC0UizDUVPKxVG+goC84k7
B1d/buYv5iga3hjwX4cPG3v/+MSARaKw1RQHORRDm22UteiL++LrEssxjd6o04cU
NrKx9HwexqGx8K3R1OOVHhiO0OlRQrPm2RfCwqvwmavqpL5tiMpTCNSXGZo6+vLt
nFxhJAaFd+F1ntExHgkHU2I5FDjDAXUXpO+KuVYo0urEO2NtdkuFDl1uWXCxJVkf
horJaHUBWXLMIjG8LaOOAmF9X/erelZTpwA1SbdY6+vCuSnfdynyUKGPcxPp/BRh
3HVOQYyJ9mdU8OXnD78LjFGD5v11284kUo6L9N1x7BciVB9tFLOr4P0ommcv7/dg
9V1Bj6x702AtBWGuQD2R9u5duKh3p/KFhk/UccIfdrK3PbqWOX8UnEmSbV3OkFkP
+kVfouIOjorJ/XhjK99Eqju5TodjRWDED3ltQyDa82tELsSngcHFWVLnBxeRmMDj
XNbKxyLX42Rh04R/KRt1v8nrvQYiUMeFZn6OmBJmYqLvId/FtOTZ8oy4Goup905j
e3x9/x82N9sKqIR7ZVsErOcrkHutcnFK1PY97o4w+mP+CHMVNJx0W6oh1aokraXA
SEp5e0AKDMV2xWSEeOPpXO6IM3U+GYUe3PZSYKS/vUgkwQb3j+lhDu5DaI1/eDLz
2bXg69yrX+A9qGOLi7m+gqtPlESQi+svHfkQJHOntxvXeov93cJXuS/xUrTPEyul
ODcW3ezmcPBtfQ6rRKH3U0r2NJb3hx+cJKpN0A96gcsaHtcj4jWJplrSNj58iBEf
3lKBWksCcESZeCzRHIYvmmqhc+RbuyrHcihVphr73s9yLSO8I36cBoM5H2dh8arp
5LKpFFobbgu3AbJN7UyQ82u1yMa5OPO5TSBGbqWlupCafyFy+belWwPkSlbck/3T
Amzs0BHEbobFPBVgKUwU1efxW4ahALAh9yfg5+PtrPUGbWvX/h483uZsL1CrnN7w
TdbU3KVyvQ8Y3EMaIub4Kdzix+v96HbP3RoiVHO7bDwy0ApD/nL/JPu7UUHURDAZ
wxapBZm8v5YLysNE2dX4dz51nbQ1ML2lnP7PTlwKV2rocKPa0uqZLyVnl4Ombe5E
UnMPYUL+kUNeR9YeD/RosYJEiccMeGkddrkpswFOdhf5b17Qj3hhuSqDGgFkUmT4
V8J8vZNVc4qnPm9n8ywtIMABFKQasnDUCcv2jMNugEK+ecYBvSslJG1l35VrDI8J
eog/XIaWwlzQkiWTpo6bVoY73SIfJKqp0l3uiZisqXPSGKCIF5Z+VeXTcJT9p88P
YB1bdUbf5dEZGkbmln6c5Gy+lc18wbX5Vq/yOQp1C2e74sU/pyHRZ1DLUKCs3A9A
4d1aGG/qGluj+AhfXaEbnlfHxQf+FSFKAE+XQUpHUDl56bisSvYranZJUamwQJ+x
uLcOTebxhx7wl9ef3VrqOnjW1wqLfgEzmxxQDEXNS2MBtviHxJ3owmlPZGUCb3h5
tuyShAKlpn1hpEJKbFjE4pU0ObmDMgsFTI8ZrH/L/dnu0mvUgyraQp4JvbUx5YJA
aNXZ/UbcU8pXiYS5CxzAlcMMybuHD88bDT1fjmFf5VsfrdecbHqdSWsyuw+X8XGP
yIztaufsOp9/ObjCeb+EjLr69i9yKo82VAbhlQJ+KpJ+XRlO/flcvKnQsiSWg0aU
e25LPpGlxhacz2NEHEByOovFBqDmM4SD9O7Dsatec2ofIKe3ac1KJdBEemfY8Qij
qA2bsdyJEOs4z2U5yY5Y2KhiSHW/oU+DRPi6/WB6VTPeuEIVLkKAToQGpa+xU/hE
s5HF74Zzl4BJE3Jd4vFLCeDAz0dEQPlNvQEUo2jm6ouWjy3SCuZoSN1d2fa/g8z0
jOni6w7GOAG4sybPh0D+I5Cbb07NFhGTPgGAdZIte2N8yEued7BinKIm7qE/ljL7
l/UxGfYyLnFIXL3q/DMWlNHzBzvVdJf5HwutBmhKFi3EaW40QFE3sK0YR9dHdD5f
XRPrTe2wYd4WwjiDdhFhS5UO4vdCcng+RKarICedoapFc9PI4Fv9P2/yTztENKsj
ck8A0hMdX4nhHpNDBAoG1KZYA05hIjJIDlbiFcMTnd0IMWP/63VZ6RY0M7nLzY1D
x05CbVR255IyNQI+6ynhXVPE5DE6S4vt5LNNKytmy4sCAui7CCPoUdPuwByP7wIU
b+100GSdkL2TUpuefjJ+AOA5vUULhHFngg5ck/pmE2wVQoBm6niQ6epQpl+1/grX
BN/+8RVNXmXgktQusuIE8CifGWIGb3YhjPOt92K80l/p5Ojf4sXqopsSXaNl8wwH
zPRCkV+Yxf/oI9+tf/lPjGf2aJTIAEtWnxh17qWFfXj9ZQ5gqeazwSf2b2BQbKVM
SDlWK6EvaDhJqH77x9bzcbIinWOhkT1SOOlxIL8TjawxIHneRoUtSbj9F7mkesU2
cpfgzOaZUUtkNQjPPxVfBrN+yg0mBz/8o28As+HQxMOMilqXNmCnx/bts5vTVmQm
jGUaw4Whies7kcl/jimp5KyBhZkFy8C88UzIZROS6Ss4aTJpI8n3W7jKrIcBnM+q
J8dG8chCNLz4VEyc3rO+vpIuNWUxBPwKZf18LUmkd6CTOy2qiVV3VmnLzdKMR9Vc
5tqY2isPn72rs6hzlzhxROuNM3VSLGNogo0gX5MDRUWWvxgjWPdGVqvckqOymCP/
uMjuHFUjOIzlykAIbP7V9VYIgsOemrZT6ieOLZt2Itz3PWz2/N4EsYEBuK8C2drw
cCxfzHzxQxwgolJubeA0qHrZ3jpvYxy6+iiqwdEkvakjedrV7vyJGHTL8PrLhOhR
7hftnk603C5iLSPB0fONXcjcvyuMLzFlMqu8dmvqU0fLJLw+VG0bZt11dmJwScwB
c1AIXv1wDPlO1JFHTK7IQAXOF9LzBvs7C/ajRiA3CQjqP31Gh5LnGnkTF5PCrnf9
wuG0swe3LVTo5wPWEIWAZHwS1OuUwLkAF5OWSin+eIkMBmFfvaOl+cChbb9lVvMS
BnONAhFJ+2P7ghXbXmlfJeIlDr9aMjCvnOTnjZyLHNDEsc/fYQ+lYpC9Vchz/jA/
lDEFd0s/iuHgVT8V/L/pv0ajaP2DPzufoE3TkS9T9F+dIHQmPf/j+XKybVd0W1cO
bHsxOZx9n46je++Ex6xzL9LxS9y8Sb9eYjEtREAFv9QId2xwzj1oMMaYpY/IjR25
xoI6kh9lBPyLev7XgSYYJRRgin8/WwbMBhhAjKkiJ0sWy6bcXuqLQA8c4L/JweEa
ov4eHAAEX66bNrUZWUtqWgEkmX3k2Lt6IvpTSTGj3KHsx1rOtchL/9/7erozM7ur
hTIOSF46iUFiEdzPSCOPNkiCsAHZpn8zCe4Wo4WpPtk7DEA8UhAqrQktED3GX1Kb
j99l6xKg2JzbKRgrlQIeIkHJTptf1gDyRFj2ux1Ite+Rxx6ba1FAH4j3OJAwDUQk
OcX5Mqrvy1v53Nv42Z7Fre1lUeTJOkeL/8iqV1LEJhVCQ8BdCwmcWTC6Mnd9hWew
2pUMMHp6S+HmzdBHISXuLbmcGGHJqwhjrh+CmZK6lDgQ8qlZm7QSl0AIjPOSroAt
AE5bfJlax5AZ4a2XVPVLz0xD1jdT9qpA+u5SvyduNdOct+4J6Ku05DiPKwLoaXJb
iJVhUfhGbnjVrGSw7jBGm1hI8nHhl63eSLN4LB+BhGzw7NKpqSlbgvlxdXbqsp/T
uGG66pz7bgr79YIKSdiaMC6VjJ2DSLVbGN0Azv7TNjrLpoyqXE1aa+5Y6rLxQC+U
DkGbIJaa2LIXcbRirNiaX5MUzxNZ+3chEF5OF7Pj4lBGy8P735OPFSP/K0xxsHsE
f0tLr4yFKHrTDPpx7fhSfjuXTadQ/pWIiOIcuEnINxKc32bKXhpfC6kNOh5dUTr3
NdRNCIboEBHBJMYpau4AZ2Kr9ytS4xqMnPXVUQK5y5hR9Pup/znMFUpA+csglgWg
YhI7SIo0rNehCIOaRBSKhb9hYngnMSnQQa6p1eZSSsqHA6uom1w/LNlY64wUYVy0
E2XfPvBOy2mkSU2RmFG1LXaf6M6UdSMDn5xTM2S2De3ylibNG1XVOjzLIeDZyYr/
/tcznPQ58L09VCkMB0ObCOoaoVgUgCBpaHX5pt7LnEEbsK5FFOZ+5LfnsVSYkLCF
DvOMbt4bpX1EOFo9Q0p1TCPNmpjrujvrx0woIHq1ieAiEBmbFg8NNlSUj/h5oUls
ueDWd2tieieDIP3+PXi3WOXtnHT6Tyk4W24eo3ACvPexOiqZZMmz47j4GaoW1jcD
9IHGp8ApJv+2+Geogma+kKNNqjeQ3ya6FaD8WuTHwsSooqJpPnzjjdyd8R3FepqT
EOQ9IhvL5TIKvS2H8wKSvNvm0M/f4r45QLSWIrL0V9ll7TpH4YO/RfcnmWD6pkk7
m9t+kw6gTDQE+OaDdCbiLLog3fSo2AkzXiawaBwsGZ4c+M8put5mxwkF/J0mJ2nq
Yj9muIpwnPTSiUhI5UOSIPKXMd3nPbX40F/0Dym91VyIyXK9mCQD1I5uwmornOK+
Ib7yjhogy6iUIvHx/XeXTCh1Wh6nCBLoJJ57ypUSw2wNEUhKlGoi5TVniz4BLdA/
R+c2NTCzUP3l5/GrZTO13n4M/IM1YPZ1FCsV04QDD8ZvVWEFbgft7OWUT3Sq20ZL
yZloWa2yIQz65IIiahgwgSzuwCMJxSAtQBd2KeM7fKO7stR1VMb7VkYvlGU2I0rQ
6Fkpu5wXI+ZxBLomCiKzhnFMu5Y6QrNqDmFTB5DHQK8daw/QRKuVQ/Nag6dKZexm
YO/ZT3k6AOVp/3Bfnj7dUJQ/dYt8c/sfdyRIK0pdaXB9L2flLgYd+LDA3SS2ndHT
ax0Mm/Q1Oq9N1oxgWy3H0fgZbAVk1vrwVqsX0BSVyT17LkRV/p4Fc93B2XHCd2OJ
g+tX+YAQC4UvhmFp7lvNNt/Vm5gA0be1gHoH2Zj1LLmAIiopA4HuTJoJVoq+bYXr
NbB1tzfDZ1uDvRUot+J9isviI1bLlVPW0TjrcwU7EWQWYbrTC84xweSiC4IZ2Z+U
+TU5SQk3wQ6qoKoU8WpSow==
`protect END_PROTECTED
