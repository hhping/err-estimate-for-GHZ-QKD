`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1xvMIHDFGU78tpzVM1e1TMVIyzl0Pa3capW6ZS3929tE4rEX4lOzH57zeDOtN8z
Ym/Aw2DrzHu32yYoIyxxtK+YfQQcRXVhvEvJHiY7h/EbMwSzso5bdD4ud68XwGGS
Qbf4nB/9t1sETZHKowAJMTIjmOyHwOFTjDm1gMIHcqErhqOHwJk1gTuBxGpawX2g
Zw5FoCArRCEumwC+yXXgDbwhvGAA21SVOTIjMp9SmeE7hsh9hCmoI9VMI9Ke/tV6
Uy5v2WGa4hro+Yet8Az/tTEz/TZRQC9QqXBOtMzu6MdCYh0IFQqW5mOyUYCxO19g
se5vcYFWSN2YL3sBu80BCw==
`protect END_PROTECTED
