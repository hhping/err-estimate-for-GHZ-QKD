`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NSJlaonAoR1fWLNZiE8t6t8ctTHDOtI7VpROT/TIq+KEOcehPo6eEs//0tJZ59MR
vsk0+/NnDonQKTIGXf/m23riZsvqb9GeFBuQ1Jgvxdx50YU8d9Xz3LhjhbhJ/mYW
NW6fRwCPEAwJWZLLM2Q10L4M89viowPGVXPtn2wmqxkke9ZBQFTMA20lLWqHEb8e
swuT/h8uAsKT01o4AElgU1azC+XYmXB3WEZfbdxOFa6HAzmX2OOHfy8DsyzuAsVr
+I/wvvEhMbsxNXcIzEExxF5EY1yn0OWEhd95NCGCHCqccCtB9c2lZgBFI3GCr4uZ
3om+uirsm7vJN8BKoTagsMf4+RMR2lv1ySLAhhh0WRiIhMX7A/mMmqeuWrzH1HP3
pWu7cr2Cg+FmZTspVb72OX+VWCEjpsmc7NWeXk6MlB+IifqdK1seNQb6LFFP8tTA
ReAPko+Yyjcqn39h0Y8atrvKmgVDXU6vGpZbdXY+JiiezwhF2nMfnr3u4Vg5dFc6
QUJnlK/CxxTmG/2Ahagg/suC4QjsA/byKPTgnLtphdFdYJlawBTbvya6nUDypZig
GwjkcJQTV1j/Pt3M05fcuZ0P9wflmo6QDYldlio2o6a67AdIN27CyFVkdlzgPklh
QqU+eiOZKikv6V4M3YEJfYJpmfLEtEqam7j4fGDFERU=
`protect END_PROTECTED
