`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yazW1k0s1x4Fa/Ny+XZHQgAuGyuRLlC5PtIYr5JnBTl8tHXPVhssZKWulPmRA42e
6L4R+Ufd/BmfDdjciznKNegeaToLeQwPV+6Zs3antVNfkCqRWk8dTCiNrFpajzpG
avi7PfKoMwWavm6z/6795XTr3kbtGTdzh3whyvn+ERY04UE0wszpM8m+gQg7Dpjv
utPHU1Gl/Tepm8QB6e6c1VppN3Uh4g9Ggo+YeRmrAT4FpSu2Gm1CO/W44Qp1/o/7
MoGemATFkf2Li1cnVwz/Edjy8u0dnvPG+kvYH5KN2HDRLg3mD6L+y2xFboF4IZjf
1lWP/k0rxlloZw12KKQ5c/457ub7S6dO0holUZI2Pczxn3VMMWWS8eOPQhsxIxa6
+1OSLKpQhVYSilNivdxPBtWPSXFcIQtooJfuVbFoDilREzfV9F8n0IHLK+bf3u9t
Ao8ryIIKrQritRX9F/Iz3Yd8tra0iZ6ZOc2Q0ttP5Ddc5gxnWUDGhqGdtX3uxJmb
DvmrRLNbMwmNhYmfYb1KwnpzBga4fLVBKJJF0dV5S2vCmeXDKlJTjWnyQS65+Jlj
MZr1Dg2P112nbAsYK2pAp3PgWxzO8A5zEzoUXUrE5fZicDQm0NDDtPQbeXYWrlQl
oToI65maUy15/KZRLhjtWjmhhQ/WEHFZClWiF1FKtgoDbvDqAAKJIFN6m2fPq+sA
SNXgwGjkDZ6GlrHWxl20M+cqSaE2kjdM6ywg20Ai6Uf1G2/j/QP4InwgxplM6QKm
fAUdLJOin4542B4ZbevXqmL1Lmmi7tfJfFExothixcEhIu0kObJQlxeWTmsCJVF2
VKdaRgTjOS21QgLmPQ80CQBwDljA9ImYAUoOD+1gmj+dSm5LYgwwHwBMUZAVCBCY
9PK5ZAbLBqGXBvdXYablBm/rZS4xILWCvLD62OvVceoBxGHV089OIv5gKhy2TDzv
BdbK31d39vAGdAkx6dmgdR6DjaCLZKuCL32Pegh51QOfjQX3DTuUYCOi8FtIAzeZ
RLRyz4/jClMhExamDPwEZjB5lCgUIVGP3rH4FYlrLumhvE5dkmMB4TsMYXm2YNH2
IaRzFhJtSlCf29cgodC985As7qK4s0qJ+giwLaKgUuiF0Tw1hsBxp4UMb+3x2qMo
OQ7WUIBjoHnAtP0MZ/ZEit+4QmgL26qRb5dw8YkC3HqaCCGYF7ZyEubIJmd4iS37
wwfqaZkGUy5s3sxw5B4IZuW8qNaiN8jvndCz+wdMefbibSIILGXhq7w7+uLdGQFB
i6yjkeiU3ClVMparEXzJq1sYpI8l8SAJKVBPYZfN9i4P5w401sAA3vUDudMHEZZ+
`protect END_PROTECTED
