`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2M7GeZiPCTS3kfc2mgpK3peV6EwatMtro9gX78ZOmD4XAAaXSOBJhR6YPsH9kycl
JJ+4ptYGBcrJey15jDUpYXDuFvHNZ5aw4D3r6qIcxAs2U+JMpf+3SMNGTpxIn6k5
m7zES5wwzeIMB08TZYMA+EQwqb9W/Wn9dwrYPQCd3e0QQBVFI+BM8EvYyV4ZqRsV
oIcRF58ai95FYWEshN0SksgW+PqXNCAeuGSZZkmw59eGUgvTQ03LfFuABJVQ7CN/
gyADoFEWLeE1E+FJzbswhL98gD/sK0QOG3djF93R4TFQsxIgI6rvCKxD8MQGXG7/
HaLIGXs6VCF2nkOU23MUejQlW0NOzHfL5y87h9i5QS8DxL1x0WPNAM+zsBtLV0xf
DKOt54FW3XPCBE28Yjgg4f8IopkZGoxBJ8NTgy4czYlLJ0/GupFOeN6cBdAlWyFM
k1wZ763CjjXWyWEFwnUbolUbKAm6Jq49R40gcYJS98JZGOgGXjslOhSxOGXPhZ9E
lYtejwdkOCyROn/qWcBYntgsqak1EYysBRSab+U6vI6dyPEbAFJ+eS6LbvJsfYrr
diIZLXTx1fJWBYN7vT9RtVVCAZfBWpURMQjmqIDQtfUmq6KdM+SMyrKjVSTunw8B
ALfIT6fSJnQfeOwBAFazmTSpMcD4bajMHvxl9xSQZdlven18yI1EfAyqRlhmuJ+q
0lEYf/ABdS7ViT5GLKh/4cdex8PXJc+QTNt+R0xxryBFWOlMyMT+++OIGkwI5bev
oxNyhTB+naiByUBytJZJ0JVff0hdy9raARo619BdjVuhy68b7LUfm0ov1GKKAZdg
gSct/5w4YnhJaN2oLnJRriuMxxWxg9Ur2hArgtZX8VTkvoKp6ca/YjKy0noi+SfV
iKuF43Fw0gPeYnuDJszCzupls1SX8SireuRrNijLyjzSsuFM/gN1C/SZD7n4Xq+t
DUM+VXpsWcleHZxaUexG8kFAudrirhklOLLtrBomsIC3m2WAKYZqaFHxthZ7dxy/
M0XNJEbcbOhTLIzG5TE1Dji1PqFJ2h0hdNhr+KCs7+Ag+z4/nO4xkL+kHqWqcvHT
uJYW++G8Z/SAoIPObfS7juC5cMM3gwRIIjmd97yfPihUJkOVI9zMPLOmAPFNNzlj
HnpZcRzbJ7WJCBCI7M7aMxDrS1/pvS46Fd+f1qn1/aZ1X27QxJpcNMdxXJ3Jyk5K
J0s6cD62piXxG3aYJCU7Xtz90GJqCGZpY1fgS+W66fid5rZKv6LaGwx23dw0eUGd
5hkiA5nMJL9UInKGc38VQ8M/BQWKv7E+UuIzx2cc28I49dVmhXMGHtrrs4xSdgFL
oQ6RRAoRYqdDeDDm6tUn1A9IrvH37WSVxUl2M53ee4ttfFb1kK71giqR+yYVNh4B
CTQv8E8YGWpkv1CoY42dnBvmUYGGe2ep4mwer1XJdsH6XPOCWmvvb073AQAs9Hbx
D6AHh81phR7Xkb2gR4EDVn0Tv0gch0GRPMloZA5sPvB2lzGigg/T2qRN2dfUvyYs
9wsBzWxYrzhOcsN3Lbw/baJIgspu8fADB5StHJrJAZPr6pnJ1SuImrG4HSgz1Dqa
npm6dic5PPNyBgNjV1By0iT9O+8iCTHJKp441/bKJLiWhpptrf61auuX3egS/VVn
l3piE4RLeXvSYUycaUHma1aSGNrTqjczGDSV/EE06aIVpzegUncQ66s9BdgnUbMP
rN00dPb2n3hKPRzIzFXr845kh+a5mI3nq6bZwToCvQAmoKTiKtAXYJU/rCeyWXkq
OV4pfdr3O+DpSOLRdMRzPi+XdzQG0SPvU78oRTLcG8K4xs/30rTqx8kBfmbupTrp
iPk2t4re1NlwU+RxJ/W+5YHvsAJ78XENft6fqYlOKpseN6vk5T4HS7wEyqHHgGdP
ZVCslIab6fKB1wrmTeuGzbrlbXBF1sQTLfuBgth+J6yDfsSF/NVTdgX45sCAyjoR
J/f0zoizkJeBDnTKc7ywlRoheSR+z2BIEDHk1+pWt+jXIN0m+L0ubZjopNlgDYey
ekpIA/kMzHoMBTu3QDj6UKS1KdrMJQRV49Ha1fMIvOhouHmZv60W0eqFdnLZcL8g
iuvSKenRxj2LGxDc7i+KniV3KIsVWJ4IpGRwLErp9q/GiWx8xcStW03QLWlv5JXx
/h2NWlWCj91sS9XFk08kvf3TQm/kPlPnPhGySjtrIms2LwrWjgxoW8DIrGtjH2C8
JjI2rGDyDqEG0ez2Z2zPSFJ5DivJdsxwIVkwLH9I2q9ifbREboQWrEk+uaT3f9lq
lypixrn7tocmWsU13vG8ATVQqkrOK2CmDx7G7A8/25R/zsOAqUWyb3ST7RjHbnor
N4+YqqVry4XtgexHxe0SIpkL0LddxV0vUkru3TPbbwAVJGD08CaHWgFALhr1z0jo
dIVb4Syhbl9w2Dna4E3pgJ4f+tFTnThvSWBT0MgH33dr68XQk7JjW0gPs/tr+pbP
uYXtR90z/5sGN3ElBPAOA7WQiTZg9mHRHoGqQf6kaxouA93ue7g0CMRfSPSTy8m7
99j/06sey5tv/lVKGQQJsogfU2vnvRXKaq3waIlgW7SYeCMGm+ZoenFJP0jodqdq
y0H37PHXIPONLxm7dDOwlahRrm8szntrqWN2rKsr+MMUIPF9p0CuQoAB25ZYHjS6
6taFrYkrUp/WmHoGSNkUpVaHUQxVXQIgChoFvCrHP0aoS71NioVhxMmfUM5HBpjJ
8H2EiwBoEUhonqQm9CBoOzMIiW6qfdN+3VOO57gqS+vjaBRA4OtVnT6DGd2EhhAE
UTH7PTHsvJRB8OBlCQACKdufbLt+ZhEM/vb8e9U9l1WHXU0R0RwtRGkjk5FeW6kV
LyGd8kngf0qHGLoLf4+gNh+E3BYhAhbXbiRGwqZiovg4CqMgI1s4fKd3Oh9mrm/j
BTbmqcmzX6TOkJkbEMB5p3o5LiggIMnxI52ZYR7tV5mj87ercb0W/+H8hpSvGu3X
DaSkAxVnO9PHuGjqJw16URRlhE4ZMp2pie2CabWsztU3QuWcN6U5Adgrt1hmEePI
`protect END_PROTECTED
