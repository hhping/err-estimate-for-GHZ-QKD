`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AIZ+z9kexTXtxMXjW9CHbI2ugKSF2CAQgyT1ApQIthnZnOCS6agTy3MNou+cTceM
+5aqM3vLxYetxcivLf1qwl8JmuYA546OfmOKdUktEcBuPoFli8+BOvCxjK4lpc4E
d1nPYasSXeenlJSFGDXpn5rSle1zhnS7Ec2woOmMlS1lazjCL8R6KsBzj2t4XxsB
Fexkn72tOqnQjUOqVS99n0rOCfu9cEIvwKE60Br5iMjwBt8S60xCZ3XzPILyegTd
x47RA4K1cCLOQ8d/yFB7qv97IGuISVzUJEFalH5VgL0bTakS/WQf/1oszJMUefG5
J7AkLD3+Tll9iOGKHA60er0BGv1wkxEsq6xgvAfsIQq9vyRMZro1IDxN3a4tVa9h
nSrmhmZeWVittZ+Tiqnk0enqyk8/tewndNWHqlpCc+Y3dpVjQ8duYqOJQ1oqedLs
vhQYY6JQ2KnqzBv60sa6GqadX2ZHFj7C+Bm05q5EBWZo21uyQ91KCg/TVy5y4d3n
b02h7O2pB0A5SBLySGlKIFc34NO4RzFx2k5rzQupfh27WGFXFEEMu11X7YFBhi3T
HRQnYs4MQD/qMTT5CDQYB4SR2RSpVREvOTFpRiHF7Gxnnb8YDDNtMI7gU8lwrSY6
rQ6BbeQHcAa2SmtdYsVcqMiXX7ggOH5qrKBsR6gyUgS6WckRsfir94b38fiXzQQP
i5kBlZDWkySew2gQRuz7hSKvXge8lf/TaK+I6LlQ+ZFehs8qXqXzugAkOmQT/gId
Jpj0VboZgFRofXS1vHkVsji4V+eD3yC2AeiOAXB8jAJ8mRZayb83l0r3Xvy2lSRJ
bWC6rnILC3nlkinZ2+JanMl96U9omC11oWrCwUt1xbMBt24hdoHqKoF2eZDVoYE2
LACZiuALNFZ3sG7o1eqtGicgwnl9n481tbk1NeyFFrR5zAPFE41Gpf9b+HLhga3p
JfoaaPUh9+w95ej5We9j1xpLCDb+znENh3zp0wEjLNO/EPFlBxY00cuN7H+Y2jSr
1hudxgalNI4AQddbqSjq86H08FVL9lhX3n77W4PyErZCjsNVfl/wTSP0yPye0JeP
puFjxutsrJStbIVfovrDLTnFPKjE0wzz00z4hUoIiux/2ErUaVwH/KXcGU2k9z6P
E2DArn6+Tf5b8s7ppChoVKBCHkleqH85IOX7WvbGpRfnTUIhUH7I7BEwpbFhdsmC
nItSnvgXaRaKoGdOddypjXWCjk4TXGy1HldyFVYo/M13kD15TFt6artydfriptEd
KdAp3TZJcy7r/je+7rVRkZaWnmmDZK+EvuUaQtfnMMYbCMnn/WYWZys66xGJkMz0
ODynA/2ZwoQhTDnGhnDSYCuLIdx/yzmQHRQJk7zgbcw4rRpVjOov33oUsB9w9FSL
FEhMXIoZjnMUY2axMzdA+7Xs++/dBjk+KKsTySqZ6jUoFp8RHpaEtyiXJuVmfo5N
ujilDg8g8pph1nSk1slM+uqZdErpGFukGuikpNj37xMXnaO+w6c382VMhgpm+1ZM
6i3IMjID6QUaVXvzZUQUF2y8b2MITtRwg8vJO+hogcPrxQh/sOQpjjT/WpsG4bUK
Yawv7jF4RDokUyE8syigVaQAvXchASCcM8hSjb3vY7D1IZ5bJ1NEFHDPTQxjmtbV
NNYy3rlyvnClL2qfkFea2Cs/elaVvcX0cNfCaq90a4SXJhnnWY374FiCn77t0xoa
Atml4S7XiupBesI5PGR5cmp2fsHyGMvuUi1bzjb01xkiIsA84QkroIp3DhZf36G4
XUyNv+5WyJCwB4ooYCJuQ8c8ICfKsuQmxoTdzSFKy8QlGpxcRqcwLfUYwxUygFhy
GqO81ba1fHMJ/rMdKrNC+lCUilA+16AAQVVddzhcXG9uBfWyVglrN3CoFK1vX9I0
4YU9lUyUVzOx0agmXLtuff/XVPxyYoc9l7QLMTa3DhEkFB8XFb7ubRmvLOiPoRo1
PAjz/wv94S2vUDCJ5niiDrSC3L2PeqNPI1kWs+pFNVzQrk/ZGGHHv85tomvMMtvJ
GbJBKCaSCMlUjk/LkVDB3uCBnaN6DIo6A2OzMUH8CNs4SpmhImHFe8gIH/T0In2m
Vl8O4WiFnkvGpzY1+Vm0IE125n5X2x4SQS9mmEQ++qYUTnrkNvEc/Dkt9fzihhQw
TA6+rKbWgljWGB5IKlImS9qhXecWl755o9U4W0+J1uKQZzJkWI55P0of9i0hweJz
yyC1/Tv8XINNMGjxl4YkK4hN9JsaJ1GmznepA+SfUrQf90i66z71jvPU/zbilz/9
n8yRRXb/PRFSp7CGNmNQS7kI2iFkgydESW6uWxeCPP/gIw3pyG2Nvf94nBnJe+hf
9Df4Yo5eutPcIqdV9nV7iwcqkdnefF56TedXHkugz+nrdf5Ahm7KXkQpxGkBu0BD
2cSQbf1LRtIH0khE5sXzIRgxvGKP+lXUKIEM+G3pBCkJehpf5mxq8ZNnvZMkc2ch
8cffPskOXtJEiZrhB4GZUau79VBkMEPHvYDODwJWD0qPdxxuuNT1XEi1kYuvCnhF
McHe+Vs/FhlJ029ZA+PsuIQj0bpFEgtSl8guVkFRb1Tal9vuI4Ta750X1Tg8g+CP
9QO1FviKEoE1p+tqq9ODb+VAeTTifeYpzB6RAu6d6oL3KPtHMDiHuV3SXGozo7uE
f+UEFF1EC6tZRaOYI2FGMlD71nxvRW0xy1FitjjNHfOdV+2htpTJghz4rbFGkEou
V7NOTTiqtj+mY6luXvlwCyI4I4eCBniEVYs1Q7erIgHxbp+UrQqLA76phK/F73Xh
CiYJ6mfNszydQ6+aA2qWoNP/mD6DDg3+CifUu2ZNXBgWoGnmFIkh4BWiJyo9mqn2
H5fij+X0gVmcXcriGgXII8CQQJp29VApJYkbSU3LnTQwG1rtKAhWrqot+ixnASEv
8TI+IoKXDbpnPd9gaWIBxD6sLjn2OmEgQqRJsNJFYsA0e7/m5MGAkQL29Zu2IKAy
hS9wKLJCX62Rn3Y/nJagAx3xWgystiBdgsIfCY2OuUsEzp82U+aCrygGv0UPPD+q
ZX4KbVO2amV/t0y+W1YQvHLUdr9+OnNbI0WX6c54qOU+MuRS8cDJ22wsIChLXGEj
TPFrPL20xEQ4nGddg9nVbt6LinavXqyqel7qw2OFYYRZsJ1VD9YA3nxrh5Il/HR2
Au4PYcGp09gyAZWUNzH60l07mr1RJ5oA4a6ZSh5lOFQEBQHOoViAB6LQrSRYddvF
IfKubcJ8m6YwvpoMOXVPTOVAXTLd64rmV0KKrHCMz8IGQM4KdQzuCPjix9rOPIhM
2jDIkJaRs888yMxYh1unVF8Gks+jNWpthq2a7MIdw606dYoWFRt8hWmI6sGoNh/E
Jx7hVwyoZ5ZHsBWHajrB4wsvAr5edNZJWBrndH4/s3ODiKRyfn0kblUhGWbHyTau
PKYyM3q4MfeWVlRAyZ6gp6R5wgJak+Y7bPD5i0XIaPDKvlLlxMkISBtLhV6OrgBJ
g0kCZ0+n5ldwbfwEzuwSf5ngzjWP+lRDMi25T2jmiADgwtbQAZoyqqJ9xqRiPl/q
tgvzojb2fKNjslokMXy5SwGl2h1ZJ2JV1KhMeh85UXwVLEOborhszPLswg7qLdwk
9J1J5TleWxmJSohSCpimoDzNRZ+1uKi9zwVrsAlo2fwsoaAwJgtqU0j7Y3y6NMt0
d99BY37GSNaQ0Q8BoMtMPM9+X8RCgutv086kioDPM5tdGXMMCh27x7l8ngcj5o/H
ThEzIH4FIInaiLDZYfxJfvrlP/iOAbpcWVCk9Ys+bbgM8skSMWUg2O04oW+dgy22
x0rhNJ+WB57djkSFCPACFbR1wVsci0PV7w/zInmTP2mLZzmEgLFPEBRwbee3sLv6
aZUyCN33Ptor22zE6gl2jWZG8aawbAtRoj8X9JUs6yfVW498TIN9Dvejen6RxJxw
PUUygRKV7jBiIWCqfiic+FyySUobslribAKPoRHUBnW9B4lbfNlfUBs8E4ltBORl
nTCWip5q9YqbcN6pNEDBUO63zHjANpc9g8eZFdeNJWf4CylJsZHmA1JHG9v4clmn
LfK99LM32r3G+p1YBfdkEdIg0YyJ88lr3lHJ6wPZICERIpTSjoofNIVoh0+Bukl3
boe2ZqaCmfUsvEheQImY6/iqL70dAfIdWUubjIlkhmh7E61z/cUbyUZO8gfrblol
pBzDZMYENOOoEIVeFoFqVRnWfCsb5WxD0W9dEaC0vz2XZIH0aTmHszHkL0UhODNq
t2UgTLcyRzwWVIp/3U6aJvHBCZOz4LPT4WDQaP/3XLpfELvJNBZRYrE12lZK1TI0
TA2hv8tISG2u83ytOxeAZBukpPnNNVl66x1qxHU4fN6DoUrOWboKNwyfL56S8N0O
YETc1aKj8fKNcHVgqpS85SCE7Kx/t5qDHbPiRv02RcNT+D6WjoSAUJHWgQnD9joX
ZCdvE1hdE3VCCisFk7dji84wS9lW/sPthkrIc1Qhp1LA5gxwnZrlchg/ANNT0upt
aHdqAo+i2nZC1XaWlvW+4wZ5QktF4SyePdOnSVa9YEzBy4MtRx2MNKwWQl/gSGcs
Ev6hjgdNpn8oX5CCH1St/ZRsqmRFWK1F5mXti3Q8woBDK/uLH7qvHwYFYmpp6Vkq
dHsx2xL7LNGci6ASZJCle4t7W9KxzDhYwdajob6we7LAsVycL4KeOS6R4iJtnit7
5tSIGWjZ1aDHXcsLOkR1QpoD2MdC9mzHtsPhwSy/OMZsU74RCTzldu8wJze+hyQX
ge9JvuHw7uzunqw8ME/Q68CbmY+4b23wIYI+Kfdryk4hwiD3UBLUYv3aj9Meyq/x
hhO46iD+3To2TBCX2y2P91ah1ey8UYEmgnopqXj/H2Rcxa1Z5kn0IHgaqCvz/R8P
lrbDcyZSqgxHnDaczQl5HPloHbteE4arXWpnl9TZRNMsw4ySREDHCiRHvu0CzJMn
QEW5HFHgLIxpVbPcZTDbwPQ4iLUXkvS70RznoJ30jxFSoRI3BUiAXDWI7LTsq3hZ
LOEQpAx6S11MidCpRcUXBnbv8tu/wbRQMG9QFwyHHRmUqC5mdbfzOlROePLh+Sml
EbyJnfJ7aJ98bO1YLMvTxF+BHyFsQuYDwrdEsCx975cdleFH+px7JjoCOxQxtf2l
bmamNz2b8YOAFzPRH4OYGgO/KQLocYg4bix976zQAVcDKDfQDrYbwBGtRazI/wnd
9mKuTPAI0olFZCkuKu9srhHDAjQ+1JXHo5mdYoUz7cGq03N8NBPDN86EYSdJhG81
6hONQIZZJVbQdh1jb3PE/+mTTTbjxY36vfacksrSEdHKjXWAVQY1f1FOB13klz28
eIGIze0K1xJek7drnCGKFTxLm9F39EO4fNO0PovCKtziDtfTIrGG3S2QMkeJHDC4
Gj9R1R5sDpubpZE9Z2TNUG7K9TpLqOCvm3Xv8wUVZZs028FaJtZOTON53F0GQriX
RLQuN4qMZScIVQi9yRy+EXoymkYCz7xN1reetrGdqJ+uWYW1Exed3rVvp7OwH6+6
IJmPGxxamzgcmYArmM3qQ0BFN0AJ5qRVgPIbKPHMIcqusnxmbx6wZ6KGiI+EYoFK
Hh7Nx6ZErMrtrvQPw2XEuMfcW2qDGP3vx7zfksPEtv5t/hfEJWbg+XD9WhvjM34n
/rfJKYPPCYziK7qf62KuyAhTsGpbqV3T8Q4KPV6rSTJWdfxvmFHxeEvTTDzm+wwE
yuW/vCPXyAyKUGc9Y0Fwvw41Mj1/LhwNYw/HLi+WlM2bGgGCdr0Y31Upkp7fWii5
zNw+oaISnnW43m1RVwB1jbGR/nPGfX4A0K0fTPAd3sU90tkO06FPoeUWonAGQnLi
duP4gnIoRt0JdjGazhcIqTl1YSKkc2UEAmA4NjkarxMvXXPuoYvZJKmfGBMGp1XK
BAhCXzUDr7sViZG9qbnBsKcXH/Iq/d/9bM4dRIzwYZBdU52YVqDASfHKZYunUlib
moEz4gP1AE6/WPOPZf6NNWCFfkF3MqUdPOB+bk9rebMnhx5RkVDTwmMylIyY/pSo
joZOPMwf0imoBZgsVeLL2hweghx5MGKxRdQ92eyiM6tfLiZCymS9295EC2lp3jMz
jIpyz5pBzZAoe6qygx7JsBPYLb2QU0nGPn9ydzlblgXg84rb9iz7iH2hQ74HVYEq
NU98XK8ByBiup2uzyBsS+jbIl2gJ3vj5qYTb8Nr7QjNnpARqs5pdvmmKzUzErmQh
0vWBg+fQ8H9XRIsv6oLr1F76G/ecUrpOYaIdjDkWNTw975gsLRlQknltN5IlvYBw
0q17ceQnoH6ZYxmTrcUhhpCTBFPb/U1WVNSSqj3rITAgunZeG4sBayYd+W5Ml7f+
uMEHQVQVbTqOFrc7T2lgUsMNQAqX9e4nqvPyZQxk7E9sKRgz+gXtGcmqaQ+/DPLM
QyTn8yo3gm3L53Pt/mYn/EJAShfsgFj65XGO/mu92ZSD4ujv5YFmKwf7UOSr71B8
cmf6nVjgN3W1v46toNUUxuBA5paqR95T8g4+x0uUyr9W1pmgJqAvvcP0huQUrplt
9YnBdi3I+1T4eSrAPwIeupmhqnJ8i0f+vG1X2EEtRsmvOp8c5l13ujh/PAQID9xt
bDJ5s1tmKgsK53d4vTFbf2HEJD5ZEf92vkCOlTRYsKSh5sxdviIJqMFnUtE810MA
XRcqVg8drXAJLVIG9dO5Zs3tBjREJNGMhdt1VJjOg5Oljyg/SrXysgfyau+OPrZz
i2g3CTHx75NKxq6ml0aGbGAm9pGAXZUvgGInWb0u0mYYsJDr3UF1zQW3FTtDc5Ya
/y+nd3iYGwlrc7tbhdpf5ImbDhxrPxhL4Ttk7qV1jzCeEQPsOieQPVcO85ZXhCbc
f4pk9+zO8ka/V0waU1fTiQnX/W5yuEwwoIU3y4QChtHL+jZjvf/kgLZvS3uRcExV
C5OexWNI5zTC5KFA5r5WYXlffi95csGdgEjTHBXVzBwoQ2YwleYoDQyugCHNyZNX
Y3vrxM5SVMZ2hvnLg2ni7EhQUC7naK7aHz62Yk+xhyTShgDhSv6hk1Q16rzyh99j
8oyqlgffp4z9G6Rnn+KvmSarvse0hKuWQxYcSUUs4JkMeL5jGm0Q8e6Q/SzmrAba
b39Van6b2OHAga2YAGpG4z2V8WVJou7mN9KT7AgV50vkSXGiZJSa4HMsm5qabW82
kVeT6jnsK94ooVEsLXTSR1bV922f6qUb8mMrUs2ZHNJJi7M3+h0USpn+ov3C+L5s
2YQxfnafKn8RvR/5vpdM6eLWRH/e147Rt5gk1sfhleVqxdSoBOpwLgB+G8755m/7
5ygZag6VZtx9BUiYh4fKLa19fO+JBUFOnNpc4COBRSybP/6cp6j3r+hY635/GLlY
rJKoo/6BAzdI6Dl3441yCsx/hfwhbGGhz5YxBMW+/wpbWpj7w7cLsnkhxVQEQ2RL
a8I8QKgc9zsIK/Ui1cxO2DxGfMXaGCZGQBlzZsbB9EqcfUncK3wdGwTYfJPSEbZa
sGrlH1gJ0OuvppiN67gAHzj9wW3j90duCg2ftvRmyt88bH+DZQozykAvAj2cdNy/
bzVMLol8W2MB58nM+rMt/CNoqFYuthcnEeQ1gWxhREOWcFGsqG6B/AAS9go10o8d
eu21idhKhNKDdy8bmvxdLvrg2OeqDylpb7MfFPsA7hkDxClh9BfIEjYtyJDvqy5a
DfMmDaop1NZh2EqKaQnKeRw2Yk6PLRntDPyRmVGv7jqGPK4UBRQZswvLh+783yyq
tPoCKGO5tJ5Ky9S1Nj9ZXnQxTiZUYJzvlJQpSQ45VTBeKuvmPPMSXbaebv+YmXtq
tK0sf23fLHA+AnFZfmUZTt9wdo34Bk4OmVUHEsMY1Y/KlK6rL7YvTYxXBxDTHoXE
6dHCkTte/PwA7MIAgKFksBFrUer1f8abobSSa/CWNYgfOv+C8uNbPMmnfs0kIiIA
NDMNoYLP6ttZwiJGng6TQuuZoierYkqNBjwLlXK1F3QYigQ5CY79NkelxEnAGHTP
pOiNH816ADQ7vpUxwJm9qkWxCMK3dZxMEjkeWQiwF1bttynQXEnVLSCvyScHAD/f
B7UWBrA30qC7c99okHurWy8JbfdlG6q4tFOc69YZ22Duuxn1MYjCTqLkHdkwTlv7
GCAdrVu+Ew8VgDgJ156wNgm29ArOQOG4Ggy4JvImXDVUdnFS+jUp36tk9sRIF8on
XnN3rXPtNqbWEBe3fl1TsYPcmm1y0lJ18xXQSPQn2j70sHhby1RUQCXo2O6N9SjF
VDtwJ8Bv56kgvKzhGZH1GOK0+7vMnFaBC5B6MhG8y0Lze2LbiN1UL/IUEJGwHMel
D8s5LZA9G3HfZKAhH/hkqOKhy0ODZ+RHvCc2yauYgu6wcUA1qc8vPzN07HwmHGIe
Ai6O71pEgDdsni4Waw3AKRVI2JUmMgqCkpYZevNjtfjEV8vhY2cdIp9TK+0QjriT
Y6ML/IIKMxKAlHYG+HUFSgjmxvZNJ2tmALaZdiOpHvNvDnjNGfcZYS+U3b+m7ea/
vM/j9tURxAK88bsICbL0a0aSrwNr3PksbJpDaZLYOAeih++bWXhjevodSiFnLE85
ogOHeutFpD5/lx7ozZEtY4AvABIgHNAkGZxfYhN7RP7kTQwMmok1czkgi1KO0Gvu
RKvUebT5rUyWJ0Oi+EVj8WgGBomTe+wd0KtS7TZGXHuX2g/cnW6MPBLM8EQA9RPK
O1fBDHCJtBLQ3Jl0r3FqVVPqR9X/PXjstWQrAvW04Hc=
`protect END_PROTECTED
