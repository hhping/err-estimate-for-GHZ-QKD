`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOUbUG3GU/rBuTt0MCQoBzinJhmCDmUswMnCdtrG6Dy8P7+9c7jCnJA6WpDSrwDN
nuTg1cZRduelakdS8R/dlId7I8GHRfazojPvZCEW/vMvlmkNySc3tOgapfRaQblO
SOlkpBuyTvsdzjE+egIql4ZJls0yZdkFGuPLCpqZPzvAZIEnMRpeUBG0g+1Iff2R
gHz1Lk/wLNyX/sq/MYwOVZeFeL6n4/saHdj3+x+ONGwd4+DJ6uvlT2hm8NEQ7rBg
7O3og25v8AWQJ51lJX1LzP4SNSa6tU/9BEV0W6Bfowwc7CQxpBgoSoMoprOtgKCc
rLaLc14rOY6Ai2q3pKxf0Qu72n3+czz4YyU9KjrqX62ScTw9nP++M5mgt2GeTnwD
JBNRb8RMNdkVBXMvsBddG5Bz429FZcM5DrxwCPwYeOPG/fTZuHkOGhyDR/MLvyZ8
J6dTlY2hmud1XjL6i2Z37J2Zmy6uonJLMIFITBKAuDQ=
`protect END_PROTECTED
