`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+apVXggEsbSjkyoDVjx26shQr7zx/Ko4Ya1VZB2VNkYDbw30/T9Nm6eh/y4I/gaS
VLh7SKEEqSfUN1VJ+2DJsRp7Ir1+CvFDOEA/A134YUrEoHRjt4B53LfZIFQLIm+p
fkZaYbJJwPYGEsP40c2P0vpd86jKl8f0pr21kX6PqfJzZv1ch+AedlZa93PKddsm
ORg2Ac/VbsSPYP8nk0Nk/2MoG2sKZM7DWPcM5AFpO49mmTfh+mQH6gUr0Yx4OAsz
dozw2CSrEEO2MFiVIef4CIgyhUdZV0jNDIZc4Sn9qwgA4wAQKSpPn6d0L6AXXj8b
ykRwk9Z6NEW1dczKAtxJf93xYfdIvlAZB/GA+Ohfzk+VLnHSUPTWZnRy+WE3g0Qp
8UAIPOO2BOXooQaPn5Z305lGnTYrtN8qg7r2jIHJKbq+RjQgmz1YxqwjmTjx6Qam
3NSBe+ps3gZxKwBUnOF0AJKaNZXsxuMhq+FaNHF3oQ1aSgGhypt/c6pnU577PQOz
6nWHL4DDq3nOlml5S8CdyWwDlyE+MEefce3ts4yRDIsn0EJEcfG31fhPyHg6If8j
/xjzuaL3hfuZMKKUaBuIvEQTKU5Kb1xYbKdj+vY6RndQ8H8k15ov3k3ulJGIpMUP
/jJXuJAZVmCiTCOYHuJdJ6/gAd00sMVV19WAWsrtuzZ9Ize+g61QCmpE7Hs8ZREo
vJSJU+V/EjavxMoAoF5giruWRmwfk8SrgptpQ0HF4eXL6le6JKdZ5heC7fnbhSgh
EPRtHVBK6EFFS4f0pvleFzHaWHClzJxAPOlAKH344OcHk1FdyMaVdQS0wpoyeyM+
FxbTLb29hAxLYcMdwijDjTP/blPsTaHCE+HOdg8Q6zJuIBhxJp9cV+1DzEVS+B0p
lXrbrlJuTPSpALZuJ/+1sK988+ADndi9i1UB3B3cP15eP9BAM0I0gSkHkAZliJ9T
64yjY1dhgH1ROpLL6I8mSGnWkLndnjbepXA85oIg8IbIv3cWz2oBsyKXyhPq9kWS
QryacjFS6/nwWT1zSj62/Js5/Un6bWulSCgRp+H0hyXv7IsqOK6PVgg3X/tLX2Nb
p2qKx2/tmghVnIRmX7UtZVfxmq1+mGbuEtmuKBjMi9bBNNFmfPOdlfVsWQMT3qTb
/G0ZqqixiTQq2Zbx/mKxzPHzJPgMfbLr2v/2vXckoXvO+0JrLeAK1EnlD1NOTwCs
k/XUZKBuPuHvTJXTjf2clqDLClRXHnrKGjnl1+dAsblQNg2YDMDPz6CXipsgWYOM
teFlyW57wlE9AsFEYpR/DL6kc/3yNtL/Cdg38t5h3cyO7Vhb5Kv668TrWSIbeEG9
Q2+QQd/Yf40wdgKySJviPd9PUxu12Q+9r4d+EgVXosbltysR6IRI3XbXBKwbmc6r
LMRrYC+gkglgxdJ3XxZqag==
`protect END_PROTECTED
