`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWkWyif1mYYpsG9ew9Kz7iXsUgjvz0Uas5JTx/UAfXX25bviLL09frDVGv+QPOgD
agYxVoZLN/ry44TYdZbAFQaf4PqXA2loMkFTNUrVflz6ffZ/lHW54kTDyL5+4A5q
a2tqbmzQCHxLQ/CIgbuSokVpwXUu7RO+SOf5byBfQSs+uIlhTVGcT4jPMo8JV43J
MIpnD2PZlW5m4/3YDcQkaMonikyPrieaWGUqCforsa1hWJw54WyN8fKrHTPXdbly
yZYohMIUi+/yXsqDDPmAG8pNaQRgQ5jplMiLX4EXaZTCWtKrCvLw8EUIQs39uBBT
eP8IecWEfDy57sud6xeuIt7yigHDSbYq6WTSKSgSIRP22jl0aV6zI5lDwgBhCv0r
AFe5LWKDAOnkZEfOdBugb0EzgOAaM6xBkIUYYHSSrwnnb+OyJplCZD3ZD0YvG6sz
iM0gThrVDl2eNjZvcnzHPpYJDS3B1tTFs88alfmUj/tTaxRPKQpau0oDqQznAyWJ
4sxF3sac4By+ImNapwIPmu8iP2IpYRrfWEP16i3mPkGCYeEJvIqrZjsPHv5AC1J0
ny+cedC26jJszZqFLyQewjpOLZI3v1wOKz2ZUM1/UkAjt4Umz/D3EW4WJpsvhITC
YEJfxfzEDLMWOzt8NB9TFtmh9qjTi/Nro0PnSSR3LZAlh81u1EXGogSJsZna5qpA
G1Y0Tlg6Y5SOSTRT3HjCcTakpCEgJQDThhXWvkaSillZSsyMC4JxMFnOh4JZNAA/
4n4Bo2btpiOTvEoFyZuq1sj3R3GAt/FJexHii3gXwfskXJDFz24EqI8v+KkUH/B8
I4Ou96ON9pke0aVeV8UPGc9yCOZ8ilGxUMhzQZLjp0ePXBs/2PwM0dwLHAYJHOP7
Vn/Uzt4NZ+pebOH7N9v5DujWj+juI+NAFbJ0xkkRhyK9hXUnl3c8zYUKeXAdLUSv
3OMNuKkogKiG8Sw7WrYl0fMTns30nXsp3/135M3uVnQVJ+duZL5Ax7+CS72hkcyY
YU99KCBvs9LytvHKPBGF1E1MFPjCeQj2DDKDSFru51HKvWcXn4iHl8oVbyQmdBAV
ns2U5beBTmmhiw3vOcoURTVqNrZ6rhYTgULWB5EiYZgnrWUDzwtTjpAptcfKhIua
2ErERMPyQ4Q7dSvDtWMOS64Tzb6HBvqIgOp2i9ZLlZX3TGBmadUC4xlieDmFYSek
51hEl1/tljpV9BbQ2U5BCgNrZzAlgoaU02H+T0h9GoU73liiD2UIY1VI4HdXpw9Y
zon7J9OFAuztiycH6oTJCiUCtS2EYkM/+XXE4/HQoBIFQqYyly85EO6SaUS6Zwkc
AoafPTv98IvIUoC0DmvYZJDofZJ3V56gqOLcO/1o1i6LuCxnNTpM1NbN8mkBrkwm
8s/OkqSK7mDo7kXFsCJQntVIGgFMI35RkVBEgMFAKpZlm4eKVVjdWkXpGYKa3c61
iHnI3h0t+ItQB4/ga0ZYWQhYJYvbvaZd7S48W0tjklTtTMUbX9cUAWlwdCqv9KzF
5fSy+H+N2aR0unEpxzH2OZ4bFbTM1yh4/K/M87wfPktB3XKNV4OCEETcjiLJZiG5
4sPcfhuwF3rmUoEydfnE7YG+zXuTzgmrgG16hfCShw6M02/qsFgVyiw8kuuzbZxg
8HGsN7m7+g6WVCYwEHhCiZYfYPx7SLwkKAKYZ1Qez1wtt256nwVqCF6k+RerzNVZ
xAAvdcQHsqDaiEZXKqzpozfc4FWr57xt3Wpok7c45/JaIGci3lSnld022yvfpOI2
zVwKqLDBiYqGlsc5QhXshLkzJFRZdhvajuAMLxybAtKsY/REFUNzdXqVQOTMezmO
e9GeI17cUk9BlCNR7AlKEZ7OUxt7y7JC+fR8N21BRdsT1okfylYdGYyJ17VC6HJ8
dt/UbbUUutkDxKY2f7Djx1CCf6BNrHuLUudlaB6NAtFpTYzkHhIVQCabtsvdWTbY
mbKnF4lpS5D3kVnonBr8V3leh2rUB6QVOS0qMZBXORg3c9QBdU3Vjl34jutK0Jwm
sP40Q1HE8TkmPU0zrf95wOWswrn2to9CcL13q6UlVZLVB2iqp+jmz+k0NlPgvxEk
7SDVmS+sTPzNXoyZ0A4r0GAvNLMd7+TxsrKSHUgK99+sDhiIvFnS5GrZ4r2G1rJA
/WwiaGALx8RDklAiIP5oKr+KZEAMQPWcGVuCCVKh2rryIrCYrncT9Cwq08/e19SQ
mPEK2sfHYMm9WkYvfqwAsq1/xezEZJgh9GITTCFsDhzTV4Sef575mkRNPlOaEl/v
W8j8+SqQzjRETkAfwRfDngWqikWsgmS8ykToChwiWZMjFVfoOesDXG3ThoCsOczD
+S3urLZQdkNfxj+0PKoQ9ociWTiXRvN4zVE/Lni2eAk/651OI8BsMe1coOblbacs
cIT8Qufa54++ki15Msch0Biqq3dvFu0WWYkOAcsen70/RNAjbVZQ3fBTkFwKRVcd
IAPrN9R1zNARwiLfHKKFjPnPzMBDrS9lYs4Q5QGx2aOpIT9lCg4+OdCVJThXPjPC
3VTvDIPhclBCBOGVTjfLI3L9BeLuZ4MrVRnbhxlge+MbyEp0ynhajhjq9hke9TO0
f9UaIfFDlVgKm1RMyYt/PO+rOPlClR/xdxJUbwDb+7oxcbH5fMOVjDBHiIQstHlQ
Z58R2N5mBf/jflD7uxCBbQEktMlKo/sAcPo3r/gAU/HThe4A1hZku5gF8C47C/uy
6S0kM6WHeKfvBGtcnGLU61ss7J3LUzniTYz4y7qrk1l+J+JemhccT+3Mzs+GTddL
Xai+fxhURoVyOOWsNi1mOK5FZyU3PiIrBJA7uYsFLJLXXTX0bBt4EGDSkn7kHgBM
CF2aT1PwW0icizPHs1aimW2DZY1T4JPMM2hnZVzxitOF7ewWo5/Ei7kh8V/ohJ3m
Spfyh7G5oO/FEo5BBc2xI4bQl5bxo2pghhJw9gt6tInr/BStR1kaqi7QyA7SxEj6
BIE7unsNLQ28ShaBf3HW5YBn7MuqdNzrdcuXOtl8TYZ6jsSOldHwBjUXttwL2SXt
UcJmp9aAfVKo/Jtg3dkIhlwPZY2LyLxbL/DrMxvzZN2uHcdGTyXzdUJ7CnKRGkby
rlU3uEj/IuNvMDV7SlulyFf2OxJtsSnubz1lemd/mQFQayjG0AB+YbE6S7lwrMpb
Pbi9vvDe9kWFpSHgJB4UXVeKCU8gRhC+7RO0ZjyyyE3q4sMRk6e9iRLfwzMqn53j
JRwl9FWJkjs3xJR7U8KjZ/ml8v/EKcFXgBGdsbMmpzBrTLZ56ioVuIwizmHLwTwA
jWWaDgamh8rUA5Tm1QDhdzob+bd057L2AOTfj1SbD3Xqq/50/FoevCj9huDs3th8
GZCWYbXpVuB3iwMEdQnrGUAZNM+43tD9CxMViV4ADbpyCPApMuogg8EpsfE8Ymz1
vjZIRShzKaEqHOafA8o4Y52bynfT75yLXs9Z9WnrdRp51ueM9pqDmKPTFy9ZtsIK
G7aAnyusVyVbgGW7cnclFWxXabzipYb9xUjzHmIwga8GpiQLlUAxjeGTQV881QGb
YDETAA4596ULJorTS9Hj7WrznvJm4hpV5IRLGqE3oV7X7L4fvo6AWETlOkqBp2Zb
+0lu+LdBUYQGK7DuV0laNZOttMsF5F+MPBw2rVI3iOf4YugdELgq9JrUiSGmatbY
hcGLNTSaLQbT1JahvbsmVp393D6nAxlgAasjALUfcM7oQ2/Suz2kXCxpb+LG92qp
d32XUaWZvRMYroQ6PGZeORoMp9cvfuOq0TKfMuhrIIqAeOGLXN4wv2Iu46GSuaEE
Ui9eUDJEwlPq9vUUfycPUZKBTpXbtP7dpVnY+qEc8trZ7WeBDUknsPEYkLbR4AZb
6SQ+qvqcpgmP7ewIqTb9FlPWwk/b8737yI4hgZt3e4x3mkM+BS+bBpIojxGowvqD
tn76IHmaJsr8jBLpmTjWgwykB9f5+frI2+WJv8q82MA/eUqrMjD4/ioAKlXHKFJ3
E/ap75UgV87Qnu0B665Zbg==
`protect END_PROTECTED
