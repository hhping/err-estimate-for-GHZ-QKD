`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWUkHNsQKvpX01O7h9/v6wKYwPPC5WSNH+OIxPU0QfVIUMZ+h5GYUJcuNt2f3AAI
8pbWufJ9ooVq8ltyS668IYgdSXYR6K/i8/HwEuaKmuG91a0bHdsWqj5dVBgyroUZ
5Uzd+8OOQzVwrTy696Y2NW3+Ac99KSshnfnEl13L0aKJ7lql3r9JYO03/RI6lAuw
f+/SgXXDb879b9AsLR6EykY7ZDGdv6hFnlKJtvRTKKIRjfo4JQzkMZz+6FYvsKDW
l62PIEooBwoKPC0ZYh7gijnGGRUggp97Sr+Hp8GRlnTgGPql0ekBj3GTZUfgTHlu
VZ3Gr0c6+xawNkvhNbCuPv2uO3o1Q5LJ4BE9vdxvdqQnTFntfl4Brs3hkWHf30ms
dM7uASBBuhl5J1/8YV7wrqgcTHyYBS2ndCBt01uYflzQ3wIYKEbMPM8fbyLQlF4K
SluDtybr3Byv4knC+OCh5Zptc7L6hOgjZBsS/q4Ir4fgmEI4TNUj4P+FZdaooqem
cQa6LY11KtwXttaOJ6jF0vuR65xOVZGIr0bDn7kVEl1IbYTH3Ai5+oGikQL8xk2W
kNai6CS30ULrEzScbq0A/8yConQqbBcYgAs0NdbvXO3z14T2QE1bTSlxP1sFVZwa
u18V19AlUT3MjFjIT78Au/ySMwWzwKwNZkNc25tc6pQWqeCPPrYVaqcc3eEZMCbr
9sNUYum51fc58Q5IdP3rl8Hdbu63mU35ZbZ5XGclSiBtuNNnDOagnalDN0WEOFAE
GU14bGK55ZR3/Cr2OBKKCyfac/WNwKQCu2VBnS2MLsmciiEzwtqnaHzCjNm9ZYs5
8rhMrjYUf9wk8DfweKP1IISIIdNrw0txOJviEBpwIHQmTfcHW/HMt/136Jx0eEIw
/vSQ+gWVxhaoQBDp/hCKm2A5j5WkYzGpBNeT59BbsU8AlOaPSh1kGVFls3wwg98x
pGtWZjX5J9UBxBqWN8WhK4CB22u4xrGRgUjq6ev4bwryt/BHW/11n2ZzL4RvFceQ
IpMMFJvrDTtvy4usqyd0m//SrzSOVLOw8PKUm5tNhFq0H26KYh/9jjxUxm8I7hjw
n3Tkfu0oRoFdsFcvnuWMgw==
`protect END_PROTECTED
