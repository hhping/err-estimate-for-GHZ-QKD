`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gps/ackvT9FeZzepk7PopipvIQyMAGMw+h4lsaxUpwUeTwu/0vVJkhzxKYuormKN
cFMyaBRIvVbTbEZh7JCrVx0GgGQ3jQKOV2t4CbAIZyVqXiM+B/1ukUjUe7N/+16b
Rbuzle8rrx8lB6J/0jpe0yZ3yiM6u90ttS1jdVo7tAq5+RxGA0VrGSExN2zbLhlE
b0ict2c6qcJlICkKIvimtgcPcCivwfQQ7/lUDl8b68NX+VVGsfkmdgoDKjFltaHy
Gyn0IuzsAUgL4tnTdSc/Mz34Btk6n9je37iRd8TDbH9qbFWKXiNg1kpykPLIJzwp
waVinjDlTuewpuB7rEUE3bgpBAtMkj2JqOV3pBweHbklZYG7qiJCFc42Qnfs69Wq
Jqv1vmMYFiKl0eBu6SLeRQzy3d20x40ryoUvtfVnGx3VMACJUX5A+9TVuA5oaTKk
mKIJfHhqNAsEh5PPzpAQBDFHH/KjN3rx3/gRTaD1vw9CpoRHHRf+tc9fCyXk4blm
R+LDA2Ljv/NvDgd9b8PYsHfPhVzHAQVWNrwCtDVypp6d8mQDkLI65ekg0BEulCHg
UjLheKxZhIShdz3pdoaA6w==
`protect END_PROTECTED
