`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x8DmvhBA/YPMBr1bl1/kk8mbPldH5evYkRGwL8zsBQ2gSSF5nipazzaWvnqrDQ8t
zGXI3iJ3xe8ZTc+ebcLRGnZoxzAkX2NBkGol8u2dPWsbhAyy1pSAb56b/G8SsJZb
qC4AaqoMTJwsOehEOifCxzp2TjtrTFSrGqLvSX7JelhIrwN0lrxNnSRzF1H479/q
JSffbJnVxZLYEtDm4kzf25Hm879tvIV4dQ9X7+tjTXxhD8IGTHu8Xaw0iXH9GOUL
l4c00zp22KBFZil/2mYvD9xudtopHgp7Uggs+eBNuf8XLmpkjF+tukomMoyiL7ZC
sJOMcbPRc9nr+3BoxkSunDm6lOhwPU79HgkoE9ks7H7/Zlozd7/RrV87DBkGqlnN
fASQGk3hItap1qdILHMsnRQY9YhwEkTcOaGwn36dLCi90UA2fDlwdpGeF4Hr3SCt
mu+mwNZgv0gq0+hnq0R5PMoP+V/GDwgoIp2ODsfIWxoyYXJOV6WaRmXRePcQZHfW
HBS7RG5htwUdPZwbgggAEEe7ArO3xquGrKNNRbd6pcausc/olREZS/rnaUVCQOLm
Jll8wyu/y4MWMmGL84fSc0h0fmfhzm6xgCXXQy68OrmVv5IhYDA4HtW9H/3xjmUs
slDStEbmhqFFHU2XnISj2wZRP5b/esMx78hxaaIhVYDpGsc5JBLmS78acAdwrlU3
H1GNF+uKJogSOVvYXSYX14m0Ys3JSZ+lnd/I4VAlPHdviePaVJr62+ZOJZh/HfpX
qEN2qh1azOK4x/mvo3MgOQACA5TqFHVjeewTc/30e07HQr2WZ8DOnFJEx28hyp1s
br0TrvMvv7j/Vs1tRpPpPqUXHU5cHvTg3G92tH2jRvCwtUa1yh0qC7ZI/B8dhMVB
TxoLTAaEKkjeEuRpniUXLgFOV46emM83oLE7OPTdWU33kIe9PnmM2y1g2HRv9T9+
QBQr4Lhgj0uCZISX1ZyTadiZGkZMT2PvFJ/AQm5jvucVTAYx2hpfcXR6dE8xe8Ow
BR3WXnburSUJZ6w7nXgac2BQK1QuT2HrMF0kpTxTjygzbnxAoLPSBAK2W2u3dmis
n3gUcftv9LCUzBrACiLZ8YJntz8iAhxbV6mynDvQ5MuzrmeVxLlLlVSyAKFcGd0b
B/EDO69FZXxyz2Shl1Bmwe5Dgkw3m4eRuksbiv/uWdDWu2q3mCcPUNoA/NqSrWbi
7rViBDavgaC6ta9GdAOGt4Idp/nierGnfFc7Cv1zdP1ZEvUwOyLVIxNF+R4ymWHa
B5kYjfaQTxKCT53ZM9ov0tt4oz83EZJ7ykdX9lG8iUWd4QJE9YmegyIgiNkbwnhp
UEkb8Ddx0Z2W4Ap42t5/26wqbBMuHOinmMJR24TH5LotoG7m0sw/cfJbTHYtkBie
pTc9zbHk+iUgwo8huvlIXePnZwKGyXxNIoUvYZOiX2iS6FCRML9z9xu6Xa27FTHW
WAOvCfeqB03odK8Q7tcAysOgvVh6pds9KbxFSDkUs58owA0K/PknBchVDSjCBboy
o9EJ4ylRFcNtkHwuBtkG7+D/4XG0DztginbEXOqlv0AlWE2uVBT/cs6o/W8Yj+H0
jSD8VUWFEd8FEktKal2lbj0zCcNqRpLA/j6OO2T42veL3YCI32HRc4iVj2oZoshU
ipXKmW9n4Nu0VVjMOsfF2z0p7bn/wwt5Z6dRoN0aKlBUEYf2S59SwiV/pyyIfSy4
+PkpiTaDRXZljTM7zQD22fnUiYV4YEwTijN4OV/Hh0a8wbJrQ4HtIK+KuZZV9ryD
lXqzwHZQqQbHDdoZ9lxp3Yt0Pyu8YAt1A1xP01NmHFulPGtozOOfJndaMc70YonE
XMXI6N4Y+5f4U/HTSxJt0ZtyOZpJ7mAEQI0Cyop6D+ZNO3JFP9Tb4/aMav0Pp6q0
T0Ev24+nzMNJGfaOPOXrJoSuqNJF+6PKqP2l1O4S8aZnLY7rloHbFrHLBn9rtgAe
iFBOaCVCKQk18jAxalx7csoC87tXY9DVCLQUZ8R8amSEHjN3Uj/8NH2YMxkhkUGW
2Jw60mcZl2c1CxFQ+xomWAF4MpuEY6yYrfjsT9kzPiF2t2TBAim8r5rLXHwatsVc
+mjqQA8ANd2p3ojuKciS8fT7oqlpye820IBzRneF4rlGupTTg0VXrdYCH2gpZlZh
x+Chf02sDRYe/BxKhCluLdWw5uTtVPXQbRN2RzIeeHyTDvINWXmNpvuQWT6d4l2o
KGyyZz/IACkJlSlyCIS5Uq9jM/F9LLL+Yj1Y2PUs311qtMm/kkwPTXfBmqmPFn/A
0/7QLV/h8mmAVGn2PddA/RbDo1tTfHFzD0+Z/uOjlsaQ+lCPJkdcoM/044denL4c
RweTGMzdJ5oIC6RoAj5skyoyCVWxDroZefClcFj/HJpRgQJ6HhdAf7x4pumwzEXH
xwpiQYFa5fRStcqXRqaG7a1H/+dk55Gpy6Dh9RuNc5GYx1sjZ1WDFdxTi++aYQYL
`protect END_PROTECTED
