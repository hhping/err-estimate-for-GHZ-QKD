`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjendlaGdJO/k5hiB1aD32IdOmaULkWhNkFAL+eF7MCawSEr1EJXcNK7tBEhsL5z
N45YbncHZxkL2IroSBQRgjcZOwmWE6iQ9iRM+Uvc5AMthpX0sKXzsdi+leb8uWCL
wdioCPva2RQrOSfqQnALeaCdMBRlP/aN/cf9Fh5gyheA4ZYXPWQKW3q38Vc4NLVv
vD22kgWe4VRHc9l9e16WTpW7imT0DMwNMHBdJVynRA05PmaZTIHxlIF94DB6+phF
1ybHZW2nQoZmaALxnibDnXyG8yQy0Ezcwx3MryjThDxF/r1a3pfNOYqWSoOBIzYx
y4EYApSMpVR5I+AignujLIS7Nty1tqvRdo6NAykEuJw5JVbnRx2O2F6n9AUPcPKq
QtZ+z1l2TzIJjtNW6OnrtCPC6CORtqslh39zCr09e9feTgBP+lhyjo0uZzfqeFKd
twvX1IU10/3uTt7V4sOvGeFcGYKTvXCJfhHtYEua7C/DnfzDNfFlsaRR0WCrAJW2
EYw+W+0+mHytp0AATsJePFCvyaNWTA3PhQ+GquI9hVK4ZjBis/JS+eTjmOkmLxJV
cSo4An1vL5UYmgyoN4Yp7/kD/eN1O86HaCAEu0VueVlL3SUu5xHdGThwZ6Y+MwWD
Q/LdXPWpgphqnhuqM3SfXUQT4PdjvXC/bQT5e34wcUtuFQGv4OaEGXw1M4Y3NwYa
Kx35mArWw6T+8zR21/XsAK77npv3st+YoDwOvjFGA9v/NjhZXm4YAgEGwRJABgDW
QzwjlGLzYCP/DHy51KB2TKxeGYSO2wADXLT3zA0e9r+FmMeBz41nEYDW3b4VwUxZ
VxR/xTAT82ubyqkZ9wtGqztPkzyfbtKKa/UG7wkJVRP/wuztTxUsrNxNz41VmjXu
tl8tBDz5GbNrrxRXQ9pWfS7dBzHVZImPmfauj7BLYpvk8ptVkE5L/tEtYDnmAJ5i
H40zSqZlSukXyagpvJ20nuke3jImYyx0ltZr7tcyWjJFXlQNTSC0JybnB3BacGHC
wd+faB+2X5XTJMo42OCzg/D8Ly5qNyJPP3099ohQg26g7FD5pndsvSs71tlnYEm0
r9j4ytCYZ27wH0LAwqKWavfnf6hr6BEdT+4c6qKSrOP0OBfzU2bPI8uKeej9wpM/
bP0peVBHMcPXpRCHKfkYThgs4RHboBGmErfdRmd3pIGgOEae3m+LMIQJJ1gEsCGJ
prWtnln9cVQCuxP4BBIk99TslpXE81wnj/uDzIim9Ek/BKVvvp2n+UxnnYFk6s5j
KRwDMOIv0XKaD5Uq1S06BLe3pfJtr0wwbVRepwMpJR/sGfFWM1cXJwX8d330xh+q
Al5OhBpJdIXQCrCn97r/sMFaZhbnpF2STnc8X3tFhtjrS18IBWpjBrf0Ec4y0JbY
wGgWCXgYzOF4wQNWG5tSu4EafeOeTSgla5TxV7gV1T55CAF3Sy9lP8XEUtXZrGkE
FUbN9lr6HrdcUexz66Iwns05MlH7BTWmnbBS+yYkjBCWUolbgxxfxzGA5iJ/e+PG
1xWD0R8CyoKABYor6u/31b3aqo0+d1kjyNK1PzP3PvdHtD/mIAoRi4mDF/bQGxX0
AVWo3BegiXvXT0T/blRDGs+9yCoBPyiesXpQzNr2xa78X3C1OETR4Kl6aO2lpAsJ
t9FgGkdmmsKQF7wSR1D6ALO3dxQBRHlej/GIO8WHjxvk5KC+HSB46bX4ETlEDODc
OruuVYK9t1V9QX0RZ+plU9+ur+1Ens+Vs8MUZHrlDS3B6hmnS8EyfcEMtbV00KGa
2MIzVdzKKzCdH+eG1tVBVixX3UcXmbPAK7ruAqwEWwcwIIqg/HsOMh471WrUltPy
oSoMGG4M6eQ6ZkIIxYxbRg1VbLXyQNRBeX+I5nNn3Gi7BF1rc8BLKX1E8goMM+JI
j6v++DHAPq5X0C7ssYKajyy2xQaOs7arQtYmfj0NGsUvfXxl6PjXifq3JZ/5M++2
fAhFSFNsjkh6UBDy8+K/y887RzbrDJU0zK07eoyVXxAXkW0GQeXbr9fVGYRaHL3Z
AFcQL+tPL/O/X5LRbOmM+j9l8kBtOCjvhwyA2SurmrRzG2D0FHLA6LbKGC0qVP6i
o2Oi9qdVuo25jCisLs7CSaSH+yF7K6fy9t7hFtin0qQkjiT4bhPdOlHkSjG9PuSs
ZB7vImAAg9L21Ak8kTaIZ5JlcBrnuDQAWggIxEB498Xaq2VisldxkWk78gH/Q9X3
VW4WbO4/s9PSqaLaDPCgdB8togHRDyBsdxHh9O3iUtv9QZB6Xd+plPRQMRHO9Tgp
em1FKMjgC1UsNgWYiOXb5Ox9HDYIk31Fh7R6mD5R/HckwLQJp1JP5bvaq3IweX0b
pTXrzHB2I7cMj07l50D/sDl6KQFBhlMMIxGbLPAxDANy8EUM7CQ5JizGuHVaCNpU
fX9TGnjuj8U2TDT/qSxnikaVoeric/ITSC+zTSyZkw/+R16f4Hbhka07lqwma2k+
C7riGFKIxkUyT+kSTcpndO7u2je/Jo99XPzMBKOaLhNSDW/B0uEVwAvIa/DQZu0d
Y2z5hhqrJATKckTNh/E6unKN5AFolF7OGYXd9CC3l5ltRQQrR8k46o8Id21ii99y
4dyq2ul7XsXrVEQ8HGY7+RaBVT9DM5uHtXfv+NFR+WG2Ab/qgQIiMqc8NFGsX59N
E5F6O/aC50tR0urqBow9QOQLrUgg2kbN176oHjIw0cKJkBuDK1NN2wCExRrW7a1F
JbM/HafCMzWvq5D1AiyQc+wtXvoqfZSgFsexa2eEBjqmImsu62mV/zX6H7rK093r
Aiy7LGdPsq4vS3Hz/AxIVu6at/TJzG2ZRa+Fd6X8v7RI0RmCZBY/2ML9daCDFLtY
gg38lWKL2D50BEqfu54+dZpqlpDVTWTBt+112UOMaZqImysg6eNjQg7CdLTRg1c0
69G/uKJNaTA/uO9BVl16p1EngCs/qkB2cZPnXNgHTAwJS4eq2cP1l8g1CDHPtA1s
HSRVT/oprXtCE9/O4D6uG4O8bliq5G59dToh0M889ExLA7bS/yG1VvYzuqAL15ER
bcuoFmQAgA6DBq9RnNGtLGFT881IFFLVzU4Gq3+IhM3/NkUEhBpnzh/6ajgJkUNG
k17ZKnWorbYWwwIpjmEGF9aX0lHSA4hwp/BqQOwZDDaW2xmgnavb+BXXECLH61Bf
`protect END_PROTECTED
