`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wMMuHchTtvn1s/cE8Dz4v0iEFfPwcEN3D95x+B4ld+aZZkAdQyGu5q1kn6vuUSsD
tNCS2a/VI3smoF4lisd8VipVOeuHWaEFfXJkyjXta8DUwWeC4jLqpffMfEB0JH9W
Cst76z0P//J3s5N6zBOf9C2iO3UOTVeM361S1XDPwpblkE/QTa0aUn0jSJDmQnzD
S39OBqs007DS7bIXiyLEFuypVxJky8/GCxwxKyI1eLZjeThZr5nGDpIZ3ENEqWrx
f94rl/gsu1tS7f84Z5t75HXFSYKOdgHa4bzB9mxBp30R6GVvQIdzAzdRw9YqPxT7
vb8o+Tt1xU1U7CYgEtco7jVgcd9QYGu+jDhuJHOM6+hCUQWUfYtiK/woGjYJVoY/
zdXqa7Wtu4gCNFZVxAx1Ysvq5J/EN6vWXm6dtt8Kjo5DAm2AkTsdHdm6l4kmtfcq
x/XQR06y4rQmtMqvwutdH/1hgMTp5LIJzAzo0wjUHTezYW216E6r+1SZFl4IRIt0
2GvBRZSQXypyzOmydPjbiOpPDT2QvEzG967irV7ZD6gqhio/vgSlq6miDQC0X1MS
c24QdcwsFMKpJGfx2p6HoFb3fkYyc84utGIAds91RwpImkEuWf5vmbg+6kGEhQzp
T7fJ4fCjbHv9RDbBfQCQp1utcEmBiomp1Yq7qORee6RIRKJW5NKE2HeVX9D9ujOf
2WHD4vmCqoqBL5RK4Ym8ioUONpiZb7tLSceohe2t3oTZWi8WzDCLW7DavTrU0cKn
NhiRSLFwTZMU538QwYS2eiWQjv2kE6ZQSzw50WI6j7/nUlrX5O12B/AHawbq+SjX
RMChyploZWfa6OHa2IlCG1AoPKis0q4VTOqRtAQ7jl2dgUPYgTVWMta3VkkvoLnt
iYC3ZVgcPZ6BL8L2r4BFCsVfd5mDNk/tzt/xNJwasOFhkrsFHDlVTBtIGnm0TEvX
RLFCe0mCe+NwO7tTAAXU3gT6LbWDF8jHon/TE50fgtGAOEhstHm/yNnntv7YhYD3
hRTEwNrX4F1+3Bn9K6ABlWLPrE43CsK/VbRxwJOlLi9tYv/M+T5QAc9LIxLLGMzs
auNvNKJfNmRCEPFAMR08af3GjvII7jxOKkyPbSTFLwLDmusPoLisYe4PVgDBWb4W
/Z3luL0bmh0sTefTlCLNDD5ow/9ICnBSdnfdpTydoRLiG6wltYf8LveFoldkxZqy
odYufq80Ga31BdxiwXgok1ymm2k40Pax6gzx3ICJ6eAf4WsPDRNhmUlW/gIXUoJO
mbbLe13kum5s13DtLiz+IZsigxcCPJNXi1ONXyyv6Qoih5CHkB4q55dAwdewOawn
I3bASMUSjxffX69jCDwwBO7NnVZwThTZi7X77SjRgKvqOMqqBT8S9mYVIDOnV2TY
tmh10cSi1CF6J+QdnA2/xOv3XX5UjHLRZl66xmZJG0zApohkomSXh2Q217NlG7AP
3/8KHkBZJNqP8AMAmaVzWlvIBeyuoCypl1+OyOEwbUSnBc+vrSmpUCIeUrw1/9RI
6c6COOQCUsv2NB7AzB16hkPp6N4R36dAzHrL4/83X7H0VKb6Wjryy+1aCXeV9cto
G408fpGWkf+wRVVzJ67c84m/fWPyDcXenHEylc6zfst0ygd+/cx1t5j424vW6vFc
dos5TZf6xpu5SHgjcqDsSuW74mhJduuQywsaTO336mE/kkXkXiYCsnfY+YDjYVjg
d52ClSX+Ptd09CahnK++A8xcrSXGUjy2Hsxh2+sa9ftanRpSYIyi4xhYo0ovq+Oe
ym7WDstvlddhPvmdqniFjcnz/Qx+7CBd1QSL6qnXTSI=
`protect END_PROTECTED
