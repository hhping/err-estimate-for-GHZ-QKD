`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Ygw6Xozbr90OE6MqzCjFTKY8BMajO3M6R2Xfy4Tibi564RXj4FPlwbZ9+617f/R
6oXw+ZHtX/KcArlitcOIKmMJFbRDpfA7sIBN1YL2brIpvN21WiC7+V5GogwbiDwI
6rFNOgmnRgrTaK+Z3TjK8TyK+SctmAZw5tVMmORW+aGvdu2xKAopq64lWfuRkbHp
eyd5wMg5po9/2GelUlNHJrn49sHA4J+AUmT6/gKGQ9VIxgTmOAhVFfjewyZKx4kP
0BhI/SqLQRQwDC18dFrshVfwAxRFqxl/DP5BGjVQDtBoSvWqwik8wLOw/ITFfUee
Wq9e0/L9EZxhzs3jqfuCTFlK8AWdkTytwKNuB1WKrg3epF5eQzlor5nvEWESnXYm
639KI/UMuM9giJIhC9IvtX1dEA8MwZ2HoCMbnCRiL9NlwkNTiNhArOHOoDDGZOTz
zlwi2bgf3v+hvwm2QLsT1/lySua5RI7GaiOi0l/t3vPOFrdEV5N2EAgGGsUnJ3ho
vQ2tgATU47EJj+HAiTWKGHIE4Hdkx0DULBH9QUVuXVOIetWla56SVE2f7Q24a7lA
4cRgpd+ZP0XXjCCdqbJuMUGB9bG8XAaTKSRXMi1IRRk/IXRx6/GAL2jWo9x1zcyd
BbMwPfqaAIlY50fUvWZ+DdtrTkc4AtyLPa91ppdG3xhUHi0znDR1eJCdiKE7sO47
Q963rwmmyYlzVOeen/jPm3Qdijv0Clb6XpuNH3OPHeZaoimmzIFcfQIYotB8YTdr
+yVfTgEyPH/3S9VIFF1kZNAVnLPrCs1pwmir5anatuJ9FqBGRsKAnNN+NhEvM3Kj
WSSdvJG9AEm1wweMYESumWP8IomdcXNqPniDqrEg26vvezMXyQ6zPHhr6wlLrWRF
sC4puSfltRCzzSYqP2hIeQFk/CBa6P6fToySvX4bjVY=
`protect END_PROTECTED
