`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pR/5YraB1/CRtMPo2Zlm2kgyV4DKkpOaxHd0zsaIPr0mgWHL7urJnclriPNhiGad
l7wQOEH8TzfVGtB4qkn6X7s9Cy2G8N7KaGXBYMG87An9bgfRhIQhB41AtFl1wAec
w1z6oxcJ9dx2NJzibXqaPJllwlFbUYxL7DmCDElPoKmJUxfyCAGNHU0/fesrZOrX
r2M4yCK087rA9FNP1oYpj1iHareDCfBrcgxFPQd1J0pMekGXgCiTc09cYPbghWqn
MPVL0SKP7gPdt+xNMtnAf1fZTr4TBnmoNJD/HUzpcEdOo8qMq8Xcv5je8j0CHL/Q
OYRufht3H7gvBquL9UiSi1an1x1vbsXJYxL3bFlSneh8hBC2yAapp6dn4uD15uza
gtlAZD1o5+MdgD0V4zQYy/MevTlJLxrOxVHflvxwKZ7tUfbcFZCVCsQzyXgiDkdN
mCCjyBtSDLfH4EJZ3zthmdk7NxoBtt4jI9+iCfqjO1+KNNrPnPMC2p7bb1zV8PP5
uzat9WgWYZ0VGM/OYwHvn7YKNMJKJzlxfidYwohmYzvhEkhg+LRlAz/TOGd9a4kb
uTjd+1kUX6bHcBYrxWMzG9ZKamAR3WOSwcVRjb0A1/EJBVu7mDKBxLjE4g4iyO9O
mBCVvGb+zyHgbV83jzmYQrJkW2J4J08DHzmYf+LMqcya4DxfaToTBaf/zfm2+Io5
7vOHUbGp9HM0U4wAL+d0Yg==
`protect END_PROTECTED
