`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5alfqBbaArNqrVChV/Wy7cIMEqZCfHoolGpwAEnC5tP2EpXt4LHaT/k+d8wsWWSO
sl6K+FOHTaAIIWRlaWJ/t3KSH9HPMzUUpPicqm6kOQRbx/iSwNMdBAs2gx+5bvJD
rWupJVFungB6ub8yTE+Nz6JwZ9xxbU404YNFpjb+uYB2EytnZkW0y0QkmEprOqCr
rI1O939JIdRUSR0oHsoH98/LKf18KQZXaE6IX20xBSuHgLzObsqqbMmGz25EOzyg
LIF6Wiv2ZpndWERtwZ2gESe3qSbkyZU0ZG3jtefeCLr5ptZRqL0xAfH8pNV3yCGN
T2op61lOoOTwfnkDmkkDSxNHn3CfSQcdAZZjC0qfJlwprq1t1W/36xRBjRm2Qe7L
Ax1j1mgZG/1jishM0WuBzAgCThRB4amQIG1bhWp4QyC8AMb0oSYJmHGQtDZg9/EK
MZWtprWxWrG2dZCQmpyUSOC1IxstmUj7qSX/AtNZig/WdlYJk1QqWWBu/IWi2f76
MGawZyvuk0CyS0ZIFn3oZjgsYLSQAzploVaJYU7P3kHK0RmDr0SpK88agm5Iqeln
uWO0f+0FGKVVfUi1dxj82EXJ+H3EplMReFst5jLqSSpIomWWn74YleThebY3Px9L
Q0UIi/JqwNClowRKiT8jZfNwC1Rl0wuB7asBO47aLNUF2Ls5CxpIn9OFVmpiPRY3
nYPHACwSc6KlCngaU5mXcVHg+mg6+CxwEm/5XjqiQMwfMbok9m5Eh4l1az/OM+dn
1wzqFwfxO8wIDSoUnoagxlP73AFxCBfdaIV1/b1YU9l1hgj/m8avPj/DFHmHmWGO
iOURYdu4OLSMNdfbpGM8IgIfioRAeOLeJWBdLRVKdnOwXCxWXmZTMtl/ws8sqRfG
mOLCk+E7ViRGKgTFAIkruT8bsqc5+0LPdNjsvNShQLHSECntaePzvl9CJamm0rxo
SY7WJ4NOqsoHs1uKnnFXfA==
`protect END_PROTECTED
