`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2DS06cEMqhxYf+5nOjVBObVg3ugyE+qJXjI3Y2PT84mxOeCZUz6hXU0ibC0GDCz+
dmIlsgfYgXqYpaHbfkbF/icj4Sn8nomgsP784+0UzbPkgz2t3H3j0UJKUcTK6cR3
+RWsb21FjAEso85ci1/JUe2i0CoUu8NnwpB/ri1eN4U+RySdJY10fWnPGuyB5gCo
GeQSLUgrtbs9Sb1y36Os457jTmBaKQEBR8e5+0ZuH1/ynw+0OfJTwi6Nx9B4V4IR
z9sdDrICTY2LgexpK3h3hOkHXOVgtwFxWAK3I5FplAO/wq4cthCKZnAmCmS73eOP
+S5vQnITHQcdcQcDEOPvWPCwQ+kk/iFqlvFVwD5Gh+g6o9LbLbrUkMtFrlGysEYa
t6k6M+eIVT/Uy5mFJ5nL/Y3EyEGXK35WPZbgkPmFFcCnHFfCqDVrHQ3079Q7ylig
GeQ6l1L+9rY2Ps05LFNPADXpnjO2ybvZRebUNxhQipo24q9KjWORiX3zKHQ0VRTT
GUpjRDrugpiXII8+7tIxRpLNvi/1U8SnZCCPeSRu/N1IUvu7JiZ8mL10VMjJZgaF
kBAVxNnhxtQfvXGP9k6uta0+lVi9wWxceJCvk0prkalA/S7qkhOj2eOoDQ72I79S
`protect END_PROTECTED
