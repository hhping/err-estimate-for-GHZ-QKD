`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iF4UPEV4snCRdkqIdP9V+NCYcSuvNovW+d8yCrjX2z1z652zqL72iwLCbALbfUag
yjW1GoSUfWg1ZMSvrARCYMhN0cA5Fphq+aCWkIXIvIV+3mDy3uiuLBlSOOZJvT2p
6YaujC/N1eHbB3dr7kCh/EMtNWpOoKyF530Mcg2n4WHfSEzYxEwEU2o5tYRfh3vY
TJ8iuMP5HJqfcFlXwySF0w5T3jmOY8eMYx0qlycaP3IWHoKZ4a0p0zVN4D2ue3fM
IWB4+AGZH2k3g1oBBQR+LTrTHo0mmoC+PfgkQNS6/fcNUKjl7RneN6KxtwyjvU5z
xbSnZutIBaUoFLmVArF/+cpiOf43OaPWv0wvyiQafWaHM6Ct+nLPnFExg7OHBdGP
5yeqTBJROh5M5eE/+jtaTLBP2jch0R0Bv4Qu8UewdPF3seOPpIw/3cTyIlNmk+ga
FedbPl+mgip7uAEu+CU8hyDeqcuk46KAOtScI9QROLkWd7SnB1Icifv3sLpc6Ndd
G8xrcrh905dZQDqNvFB0r90i3T2E+n6I31XiNSJIaUXk0FGDuE/gINMdZOvN/b2Q
1gNrZVaEzlNl+BLigAuBxT0XlgWd1MCqZSlFP3SIZYb0gYdZlHy5M1jMy/bTzYR+
aZkBu9cg/vH11ThTBBnG2ciE4dQ1B+YFsrXn35NCoGXUWaSShjIOkuRz8FcUShQ6
beHxO6b5ilW45vO9WpC3sICza7oAAY10vGIvkvs10CVeR52Vqw1zb/h5K4VXhLTP
bKRn/+XhRiyGM0ZgA0CSQlPrYyvAH+8O0w4NHKim90gE0rEfeUBKZChsh24rUfBG
0fe0XklrJFanOc2s27Hro0aX0WYZXwZEQr2cM2Vus1j1kAmIrYILLEsN2WwO0nTQ
ao/YrlE3FICjsT00woM7eu4hcojHdK9TAog6AVKSHda+Vf2r01YtwB62CBXvzUMC
K0gVJpSZ8S788lRN7Sj2fk1sCdUzuXI4pvfBJbYWq4Mu6WjbEQIuLRm8uZ53ABJB
6/OhxGCcDRwjsz8LfIT8KlmblubEk1CR7cwvEBDgL+DRWslcADMDO2a0fizC3jqj
oEFhZskiwgQjPKk/mthi2j+WaPnqtX3wdBcUiyzidqPhubMoweJNa5IyVC52JDle
jBmAIi1E8Wjc1zTDD1yGhvttKkEdz/DaoXhp6CbvIzgwKGv0a1C3TkAvAIiohElB
W7nxTDGonojNbfqUIDZkJCmHW5okhAItEVkopj8POaJi7vesGcViuU/ALSsKkW5h
`protect END_PROTECTED
