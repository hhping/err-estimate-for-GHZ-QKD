`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kXq7I9qiC8+p93/JVrJBLdU07bACpB7cztQSj/YLhlg/j2iV6euL9LZnILorPeqc
3idsYNPfCxwhq+DSP703GpsllhIxhGQL9Sqa+yyn/Nh7CiNe1rteRCF7IpxKR2Zg
dQy/779h5ERRnPkawICWlVt/jUYf0vLHgs9VfBRUGOXmDtJAqI2mFDtwNUJAqL+N
xabf9Kx/qhXDx+yBfSqrSLm5fqUqn0gCiYuFNYluoDwmX55Pq34JOrRAMGDuWCiB
w/y+lTFr5XnqnVVXP1lScg3U/8IT91AXU83PA3jtOOUEFW8+pkWXJTYD4bOn6w38
jT8RmQTV+Vei33Rair7eX8argYPAAncfhiEhPSXT2QXhwQ8iWhggoqc43d12p6MI
yIZ3sCXFX4w6ITB+9AcrzEMvSBkehA2HMIUK2XEvNJcosOXbiulFZEspkGHQRRq0
3btlItbhGpTOV1SOITIvC22JgDXNFaiDXk2EeY+nK4Q+8sX/KdxybVg791PJknIa
+Wb8PEpmQznO29igBNx/hp4tJ9DtTUXUD5nhj5JYsPiKjb3qu7Wn/9vfJkweMauV
iko1GKwf8mrm5h6bX9AX3M35LkLzdI6nnUMJdUDn8ajAjjLn0BE9uLa0R25nhyhY
siPuxDqesoaNLw4swqFaDpVVs7ieinh2CwD189GmE5Up857SgL6Le7rO4ltjLU8L
hH1nnYtGvfQnBnjCuR3RP6FtD76IW0nGSxhPQuRE8Cl8xC4153gLKHKW52UrOoOI
LPlw0crBbZ5mjJdebODVCz4ccb4Qi2h9/RVI9OHAsPdnpBpisioua+MuDnU0tpaA
xgqQ29Dnuife2tw5mJXdf3djtlNnfXUphdYXIEw+lY4WHi4rovVOa3jL3vrDOrBu
qcmUwcaOPvbAm4BjPkcc/4BrHzMeciZ5pSJLPAaqCuklAMcisQ9in3YO7SV+VIpY
VamI1pPueuGMLHiD7wwgyJabUHH7LiXfS097jEcFcUjbPLC9S+6MWMMsE/wsRpsO
iUIK5oddnpJVdQy/frV5KiTNAgiWSLnic4zg1pZ8DQ4=
`protect END_PROTECTED
