`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2yyP+nakEd609AQcy94zso/lYvmsifYAf2xSfpNLRz5picOpKkSUiVN4vosAiqoD
ccuorinY05cOMXnhl84HVJ80SNkIsqJtosS79ar3i8jrGT/ePmS+2Q5J2dSJqgVA
jNmoqTXPreadVOXAKZcgi8QjoH2D7DjLnp/mJp9Gx0ODQh7pzXpb8uuHQGcpqpIa
xruBYg3vR3TnZsPXU9LP59eqxoHTAIdXf/rIG3ariNgCpPVFsaLUKvGVyaIQjwrf
NddSlnlZ0hHavcLxINmPKkOL10ZV9jRpjvDG+j9tx30pZSiRFqw2Rlt8VuAflmf2
j9wrdGDsXoWp6yMHKK+TesPGka1pmizk8w4wu0lMXUaAI6fdtygFcKgOr954/Zgp
HA5QoLq6gqB9WgRpgahPZKKX+Qv/Z+sMqFALihvK5ni5G7mtYlWxxhkwRzHkCBBh
TGN2Tw4ErjIXYnDGOB/L7lE7kD4u+Pi+8Lv47C+M+xFWlfFr6OohSP+6jAjNDEy4
871USYKvb7V0xsP/vi9Z67ngJuy0Gtq/ZK46pyW8bCLIfDbqGxDOMmNO4r0K1qJ/
TVghQ0dTnBk5Eg82z7NkbZGvl9StLuTGf6BlzxD//QdOP3u7/Mg4mXZf33Ss281b
MI0c5ddL3qXFqlt/COaCKngDJJXqaQKdB8Jgh2Tb/3h46rzB4rJdYrPRA/ar561B
tVqpjc3PxxiK7lORGeH3e7WMt7YKcv9D18OWZ8WxE9eOuu3wvK3XrAZEANohWUCB
mqvI3ewDY8oB1W7PPiWf1aelXMLZ/f/8/bMy5WZ+eJTNYyGhya+dSNzfk8vpjD09
r6r5YfrTMdcItPAQPcQ33CC6MFVmtVn0kCHNXHoulQ9aLdii6dY+WwnBCa5tgnjr
N82/C6nOvD5c1tRmmQe9NzK6YCSllYhoDe9xuCyszaMyfcq9nAnE3Gw0/2QGz0Ae
fmImi1FLQUn+xcv7XT6r+D/rT0fOlScsdNEUI/+vTimNz2XS5op7vgtpktpWV2qQ
nGfheggLL4yLMKFdKybzfOVRmi9p+qX25XbX5VWB8ByTrFa24pypW0fKChvsto5F
aM/YrO0+kpS3AFy8+r+AbkzDPAxELn7dDKyWF0EdUMWO2aISPiaa+fjg5dFtJdrf
dx6azHdB9YSI6tMCsqG2Kzh8ZN/xWN3zPzq/fKgoMt3KICHR8KcdaZQinDZHvPC6
SHEfs+3b38OCLpZu7wCdwsG41F9UgVB+0dhIquHd3gnTZKqOZkmzsv4KwM4A0kQl
qz3s+3xaBIB7cvWKnu0E1lsHNwsRtpOuNZplrH1+HnAQXX9G2EQWBfHSxK+gVC0G
spQfkv8YaXqAomwlBOx05YgMZwUhMRIL6eCLuh4uJuoHGkm0XA44CJh1ldE5Ah0b
KCIX2qIDNh/lrjiUE0BcR5EM6Cl3Cm9KgkVMP6O8EFc/iDfL8yxZ3Cgw0MjOjlA8
e2u+V/2/XOquFddLK//PcmgAIfel6eM/ZbFRdFE3F37wr6yP5dmOmh4SwHOcphF8
JwQZf4bXSPvxE/C2mpPJYPW5DU4hyXvqs+0lCOpim6oGgIB7zaO5HUBKjTA2BouE
vVaA0seRBJNjM+7fY9fN1n6+oksFALn1+iHd1+s0Urk4GGEFYLySCtxAGgnDEgei
W71vo9sH80OCeq4Fq8RptjYo/Wi1G1Na990fzrAwGQHa3lrBzdvE5Y/7imnPU316
BQYb8HXKIKtYhl6M0L/u6bTIMce7dGMbfCLZ3wvee+7411jFSZByCpBlnu/WoeDp
uQSGMujfbR9OWRixS8TkE3hyUh/8WRL1UlzED7qGmX2Ca2rfepzeH7uH1dlG/IdA
WzBkv0oUhdv+PAkR6mqZG7QhPzFh2VuK+YP5D7iaK7s8IXkX1enckNdW0cDKeFpk
vvMWKKSqGvtACedsYZSK6uyB60WgewMGz0QCRVilLyKJ54QuPcGyf/5JeAWEKXkb
1pCgx09lOENjNzFaDuwUvgfaVaKacYqRXUPVGZ8CwObBUzN3U76Nswe3pKFh4HfP
khfPmCJ6pbY+kbXIqZZwnTNx5dtw9dYyVBoGrHKHDzhZ3IhZrQl7Fl4kqIu02Gfz
NxVesOGddi+d/lDf5WgAuQoSqf7M0Fw5avOVfhXxyFpXV8/8Ig2cA/XooU49/Qpy
GN1p7pNppPk7niG8qJBOffwyk/Ul6cotsFlHCllHDtlJOjd21UfdPkm61syGXYes
ShAI2mYxsh+1YCTeQFQyd10uTAnHGstXJEHHFhGTXXCl0gvAhAcHbH8P8HCLpvC0
aZxVTIaP66dzE0jsSZ/OWwHgwZvsfcWIW4zHnKBz2G+jAGNkv9VWi/cjlQA0CLK1
LFfLFV3lPkQvKOAXL232W7KDvIr7xlhslqL1r9xvyrCspEzhpxmVi+P5/d2ovTgE
8rXQSVAkiZT+bNred2mC02mqePUPtf+6ILs5Lm50ubKyyVHoJ4Ysg4unsLwaeeOd
g5KNBG6Yw1CIi5lUqzdLxs1Tus93xPsnX60Lb/KZWtadEuNKQppxhKiZG6DfVDdX
cyxCsJ2cFepY2HhSfLTd4aTv33P4ptqPOAY1im+eQ6ShBBUnlOUIZLoM7V9n76UP
utf7F/q54f4FMPLvya0SudRoeQfzfcVHMNyVeD/wIg0NOk3dwVEqb/Yvsg022Fvd
oCY772r5kBN+U8ELvaqNXe854Pu9BBu3kkB9OKN61m7g8W9E1U8amBHoYxaVr+dl
in/KE/chNj6bNb7DwYunoCSP8JoD47pO4mmyT6W3TJM77fssVKiYL3CIq3FUL5FR
GHb9lelfBpRUsNm8GoeN0BKCrFMAlk9tMEZqNeBGc/3rntw8b3+PJkcZhKht8qXY
I6aMngGv6gS1V72mftBoA2elGEUdjcc0plz+VGMZ03rYR9eNAXotJGG72kSulMmh
1MMiPpvggMpjBYvJ0FM8Uip+ae3RjaDVyuQjUHJPTxTbQSvFoYwsM5XnQtJ7/sa7
EmchBolwHPBHB0yQGW4XmOPDWclfjMqsH7p8cGl6BxhYrO8DtcWskAq5SRsnVC7J
/xtAVyS8hLFeZC8LQlH/H0ubT5Wbrku/VKcv8I2Gg+T6mZ2GujEOhvakrO5xXPbf
7UpMEqOpqBjerocVuR4tPRJhQSIH1SjiSTXDDJLQsVguFIk3QrUIg0v/fI2qAeh6
jAEUtmdpViHIMnz0cHSYtwzfRzYixs3RKSbjsmOw44Fy2XvkIHpCiBdZYvY+H+h0
1EvIZyPo2pP7SU4UcniRTgtEDeGmRorFxEtiaVZJFUpN9k8D2BJXy+UGx10jBGli
pznXpUP1ikyGE+Bj9acQKYe5EJO1hhsskMi6veAWnMZyx7m+r0NTsSsYy3sjcRJW
+lvZhsrD8E+eQKhwg3cPq43C9W5T0EGX2pY29MmQIPVymLYrxZjHoFBeRbh6MdwD
yX5Qna2qadOWFnpr+78233MNqxgpjz7ar/VdI3Ast4uouYH2EFWSQUfGOcCxvDki
Mbn/JCHGHVcJ0OSqxvS8DazTA32QGMOvJ37BVX4GrcdBkSRoLg+yLE8ewuvvtRE6
Xk+P0E73oHYs8ME/dG3H1ATfYFJ7mj3Sd8LS/QnsNl0qUbDM+T6Q5HF2FUcAgZJR
9NK1t4pOh4oNFFVZxOUcbcDKTku6fKOt8Ozr/eJr9ux78LtEAHZcqGLSaTnOTVW4
go6X1fOlJN9pY4XB99T/7vhrfaY/ir+lbkEsDGl5A7/kcvn2GUkY8qulhJRh/7wY
`protect END_PROTECTED
