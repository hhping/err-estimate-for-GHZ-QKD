library verilog;
use verilog.vl_types.all;
entity twentynm_cmu_fpll_refclk_select is
    generic(
        enable_debug_info: string  := "true";
        mux0_inclk0_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux0_inclk1_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux0_inclk2_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux0_inclk3_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux0_inclk4_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux1_inclk0_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux1_inclk1_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux1_inclk2_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux1_inclk3_logical_to_physical_mapping: string  := "ref_iqclk0";
        mux1_inclk4_logical_to_physical_mapping: string  := "ref_iqclk0";
        pll_auto_clk_sw_en: string  := "false";
        pll_clk_loss_edge: string  := "pll_clk_loss_both_edges";
        pll_clk_loss_sw_en: string  := "false";
        pll_clk_sel_override: string  := "normal";
        pll_clk_sel_override_value: string  := "select_clk0";
        pll_clk_sw_dly  : integer := 0;
        pll_clkin_0_scratch0_src: string  := "pll_clkin_0_scratch0_src_vss";
        pll_clkin_0_scratch1_src: string  := "pll_clkin_0_scratch1_src_vss";
        pll_clkin_0_scratch2_src: string  := "pll_clkin_0_scratch2_src_vss";
        pll_clkin_0_scratch3_src: string  := "pll_clkin_0_scratch3_src_vss";
        pll_clkin_0_scratch4_src: string  := "pll_clkin_0_scratch4_src_vss";
        pll_clkin_0_src : string  := "pll_clkin_0_src_vss";
        pll_clkin_1_scratch0_src: string  := "pll_clkin_1_scratch0_src_vss";
        pll_clkin_1_scratch1_src: string  := "pll_clkin_1_scratch1_src_vss";
        pll_clkin_1_scratch2_src: string  := "pll_clkin_1_scratch2_src_vss";
        pll_clkin_1_scratch3_src: string  := "pll_clkin_1_scratch3_src_vss";
        pll_clkin_1_scratch4_src: string  := "pll_clkin_1_scratch4_src_vss";
        pll_clkin_1_src : string  := "pll_clkin_1_src_vss";
        pll_manu_clk_sw_en: string  := "false";
        pll_powerdown_mode: string  := "false";
        pll_sup_mode    : string  := "user_mode";
        pll_sw_refclk_src: string  := "pll_sw_refclk_src_clk_0";
        refclk_select0  : string  := "ref_iqclk0";
        refclk_select1  : string  := "ref_iqclk0";
        silicon_rev     : string  := "20nm5es";
        xpm_iqref_mux0_iqclk_sel: string  := "power_down";
        xpm_iqref_mux0_scratch0_src: string  := "scratch0_power_down";
        xpm_iqref_mux0_scratch1_src: string  := "scratch1_power_down";
        xpm_iqref_mux0_scratch2_src: string  := "scratch2_power_down";
        xpm_iqref_mux0_scratch3_src: string  := "scratch3_power_down";
        xpm_iqref_mux0_scratch4_src: string  := "scratch4_power_down";
        xpm_iqref_mux1_iqclk_sel: string  := "power_down";
        xpm_iqref_mux1_scratch0_src: string  := "scratch0_power_down";
        xpm_iqref_mux1_scratch1_src: string  := "scratch1_power_down";
        xpm_iqref_mux1_scratch2_src: string  := "scratch2_power_down";
        xpm_iqref_mux1_scratch3_src: string  := "scratch3_power_down";
        xpm_iqref_mux1_scratch4_src: string  := "scratch4_power_down"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        core_refclk     : in     vl_logic;
        extswitch       : in     vl_logic;
        fpll_cr_pllen   : in     vl_logic;
        iqtxrxclk       : in     vl_logic_vector(5 downto 0);
        refclk          : in     vl_logic;
        pll_cascade_in  : in     vl_logic;
        ref_iqclk       : in     vl_logic_vector(11 downto 0);
        tx_rx_core_refclk: in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        clk_src         : out    vl_logic_vector(1 downto 0);
        clk0bad         : out    vl_logic;
        clk1bad         : out    vl_logic;
        outclk          : out    vl_logic;
        extswitch_buf   : out    vl_logic;
        pllclksel       : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of mux0_inclk0_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux0_inclk1_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux0_inclk2_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux0_inclk3_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux0_inclk4_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux1_inclk0_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux1_inclk1_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux1_inclk2_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux1_inclk3_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of mux1_inclk4_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of pll_auto_clk_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_loss_edge : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_loss_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_sel_override : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_sel_override_value : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_sw_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_scratch0_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_scratch1_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_scratch2_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_scratch3_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_scratch4_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_scratch0_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_scratch1_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_scratch2_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_scratch3_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_scratch4_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_src : constant is 1;
    attribute mti_svvh_generic_type of pll_manu_clk_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_powerdown_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_sw_refclk_src : constant is 1;
    attribute mti_svvh_generic_type of refclk_select0 : constant is 1;
    attribute mti_svvh_generic_type of refclk_select1 : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux0_iqclk_sel : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux0_scratch0_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux0_scratch1_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux0_scratch2_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux0_scratch3_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux0_scratch4_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux1_iqclk_sel : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux1_scratch0_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux1_scratch1_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux1_scratch2_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux1_scratch3_src : constant is 1;
    attribute mti_svvh_generic_type of xpm_iqref_mux1_scratch4_src : constant is 1;
end twentynm_cmu_fpll_refclk_select;
