`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5GnKbJK9x91XoeT4IhEmslMbHTxQajlO6gN8q9FlYjIgjvtLCIt0zwiGZd0z1bMk
YLl5lepwifPda8WEZXGxicIj6gldMpcnGM2oHdwsYcXQfsa0s64EOwFNRk/yA7ai
v4OuzVdtszxaw2S5DKCKvyjxKBfWHlxdsOnUrCZsZpzbq68dHqdqukljzXn+6x0C
HSFSWZdSPy/0Oo/GkXLyLT8GOCbIFoNb7BCpI50++AaZpN8kbxTmtFjjL1ia7SsC
Q/NmlXHKBaCmojknHHsvPo17gpG2PDtO3ECDUGMdlKlCC8t4pCJoRk9TQoJ3Zdmi
Ey8Hh4Hrx+ZlPsY7/XmTw0ajzFMB69rFxwtUxSQJN6AR8LFvp6ZF/hYyksCH5WHl
vt89bkH6zFHDrxpPJLLXgZr0sqV9nl6HTeUGt3MMBh5NE148K3jjKwU/FSOgfFmd
YkaYohsBPL5hfiE0UumFtnPRuc3s7sTK1E+VeebBTU62ldmw/7B12R1dax4sBU9V
op3Tne+5SKwkqJI6dPvELDMNHry2eiDrISa9c7IhTZec76CM0z+8LlZ50+Af0lOZ
PpaSOFpgjRKIwiDYv8ghl0qFoXwGl/7RldvU7kPyOrjkP/Y73nw/3C97eKOepLdm
GS0ueDUHbdzSLJY6r2LeGyhE8dugh0QBc4ex9vUsX1dcgp4xJQBpCRchlPHxnuk2
SXwaAebBECNFvWgqJM71oqbN6oUKxglxJYiWHSq0NF+KqTHS7pgph6bF8IoQKlVw
dhSUR7yqkJqL+CVLK3dL2em48d2BNMFn0G2AGa9pPt2X8lmQliC+yeTSWlA+y7t8
2TLb/Oi9JsjviiRzAD/SldbJ3o+a5UVuebVj2LnqSJD2dmOFMk9Wwlu65F2vIWGy
/HZfx+jpY21BwIeiRYrdAMpOBeycpyl63+108jtQQgNxSsILTqsHMulJXdh2pL7p
48uryZVwvjtC/Bnog2kR7fDcvQeuBdoAYeu2BM7xhGVX0rT4IwHGqwTzKc4udG3G
wSqDTrnnzLRmMxZjGuV+h3n3ywEaVNspNy3531pcCqvgepLXNqLEQVGQECZYLDPs
S7EJ3Air9Dm9HxoyytK8abCIvNbA1WiGOOcBiCC7NphIywv8fk9flTtI+3XLCFpX
CDHbRFSsEyrQCCyfo2SD057WHbz2Ex3Pa31CFvjGZSMUefcxqNGKTHqGTRDrP28p
qr9WI18P/pyheMAPWKInjzvFs/NKZwOxxdZaXo18gZF/ziKQetuI+/9MyQzjG1Lu
memi0vAGq9K0JEvVAw9iu9kwLZq55pt8hNGUwWivtUCUS/pVrZ1WvGY3R65YgNfH
CO8cIrMv8Qw7QubJuqW6FFgH9X1CrSU6PfltzgSLc6fWrsPntqJcalXCPCktBsgD
ps03SSNKVysK7rVQSqamoBumG3pQ++ZuHyH4sWRHyx4=
`protect END_PROTECTED
