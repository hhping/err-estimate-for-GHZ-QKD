`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+a/5ZQ+bHF3brm6EEbOlVsTTO9W4YlWKbURVCnane0lfyhJSHqQVcMf1N+CE+I4
9tYA3WUfUolJafdmbdcE9yRyqRbDGt40jEHKpmWOgQAOuYzwgPN5hGXbE4i+3+gO
9BGILAQ3EfxGYUeCBZ4qaNYqt15ltPo7rWVS0jPBZo+5vGHs1GpX3CdnRSQ/AQi2
b8a/sToeTTMiQRrwcSnWTM6L4k88BKH/Hed9kG1qY3Q1+kbgsbgiIg83DdeOS8Ec
fHY7/hxq79fY13qe0M5tlcUNi/eIeHeC9QXOJR8NQysZ3dpYEvnDNlN23uJ1o7lj
LZGM6GdjCLvmjEVNwn4KgUxk6qxoYnhWo6OTArUm2lFwF988bHSfFGKnlQHic12L
IGyQpFlTG3SYg5ENpsE1jPo1UvNfQ+MbWI2P6alqsTJUWf5uESBfezJV7EbDFWX2
bAq+S8ughMvy9ncbz4Ysmpb674yPl5T791FNYTyY394ZFgbFMRWfMqfXuY9hCssx
Gvf+ioDtYlgkW+rmZnoCP10utAb7Zte/tXcnLpSaqPqx1kGKJLGMzZ481nIM5+vu
JUMer6Aq3kFkiGvjEDNcyPtbTrDblz0/eP1jVn+o5lafzflPRgFPIPMlRwJqzW1Z
c/TcXowiN70iIZD7L2iuBMZ9onMBt9zVUz2IJNJHiubKQckiPee8UN0lrApZpu4X
KWUWZnvAwwjYcdzfkc785ie8M8Q1pSVAYSvlKhCxbrlBbzRmCI2DLncxihzBGHO2
C7Wdc3fknVGd07yOUmMzD8so/7sgiKdl6CRuK6/v+asQi2LsHNrvfGIt7elBXFXh
zqXm3kr5wWbKKuHUdFe9ce443Y7GOsN4ZpBaiRyFqwcvz5DdjEXas7BZ3mO45Dw/
rBrlcF9a4RL+xEvbs0qZwufCMWoJLD96MMPtmZP+zz9ntzPWccScSKp5iAsal6cm
jIZfq+yccBuohrO3tfisFtohXVRVxAF+8DvNclwR6PGg17pggrP5WUY9+rvfNqso
MfBnvXZbEWFK5EjuPppg0P9H/Hxzdq7YnnkTI1G0ncHAY7knbTi37HnsZrRWtrYF
mMeg/Nmcz3bfeUtnFBzFRcsKZuPYSsiZjmyCIeXJmcp43Sks6M9i2Iwucy0ItGpz
VYuGP48hfeD3ERV/rhfGuCR4cLyem5pv5eSWvJpsQtIjrx+i/RnGLZam3U2O9ftQ
QDOIKgaQtDccKn+GOXNEu2a/CnDc042tbBs1YeC6e1dwlltGlI7yCr54AulCyNNi
T4xZtr1oppVE0dy7YEg2vyE8FBeiQaFY+vi03wdCzoz1dFIFBczvRMcFQ+ymF5pE
YHIxZ7Ip0RZ2qv2DwWrNQtqZuZtAO3pTcckdpkJVYb+mvZk/N6CDMrTYE4RTeqai
/uE5RVMKbB94yIcqYfH98LDv7gRuUoxRkcQrATe/4PN0Tn3v0YlE/RnjXICig4+9
5qTUsaW2Tmojlyuc9ZurjOVH9CO0lOlk1kmQL/WDnzo+FZ6gFqhFwVDqzOacQ6+3
8X+384LVTlpJC3VxVnI154tKy271UQI3W6lLKx9YRiP6mYT35YNtcL28G94HowoP
D4TFrvtLWWx4+57BTrxpMD5+Dc9DSV/UIopzQgDBo59Td53umG1IeaCNwL02pYa+
QiSfbQ+DhVjpQrM9aKTIkEGbvmhnWQRhqNMG8qB7Vk0q7mOZW6SicjJlMM3i+UqH
iU8rzTpJvpMtnvx9yjzd49dNdZm7SL6pEU1/FBVu3oZaOmGTJXZEJ3LWS/72ZvJ7
WC86MDyd5zAN/S7BWdzjAUQlxWFGNtAXp6Ifqbs90q6Wtam65tuKVWancyjQd/9S
QF8yP/CUy6WpqFFf+DEFh9wfjr3xxI8tzJeSM+IEWUNDGhoMRCMINh4rvhbKLhyL
hvX5KZXg+OSuoDYzxJpnVycbYF4+oqUAap8tDuBOlxlj19E9c0w9Kf8Eq/j29xtX
1ozGuWBNr7kJZOT4lGRM9ha+XsdePcGQGBZUKlEEvndRvm5LgYw9Z9bqeVO1gRbl
S/A0O3lsnLiaUvK7W/u0aUgc4UNJdvJm1Xa1uZDTUZkEWcenVIWGU3wZP4Lp0sEj
vSE7cfvLAW695Ijqn6YegMvNwObDEZfcLx2FXQdYTgWVRSdkCVwnKwmjsmJGI+x7
pfWfBXR9OrSrLg+p4kba+nzgdBFZAWftfdMWLlmz8RBhy0NvbdKn1PYYTRUnbXyC
hnnl88vhasQ0GovY8HOQjzpSXLK2StzTClFS5DDFVqTFpSCku1ocQod7xXaqvbf6
YOBW5uC96Waee7TZir1d7+ZU7b8vvsqEtYYKHaB1/YzGmLtCr4pusKvX4FVcpQxE
UfBKgRp65mmpxVYd1AXGqgbXQGxvnHrWL42/7cWu3CD8lKTGlVzeJ1oGdhYHYzkK
hodsN+GsGq3typNGs3n2UfenGHnYxhJzcnOMZjbUebyGDAnOSydeiebEjzh4ZJY1
Dm/wOtA492f18pXDnMc21GJtWOlTm7e7dViTbvNcDuJ4iRXEhttLTfbaOVU+TqJN
toLVY3Ae7XLSniZLhoXnJjroFJErRmlblz3Kurw1Rp4AJavLDSIKPf0/aGL2bbiW
pymhbQPCcZWggEmnFElGShVNUIF67JF7TZDSIf9+Ow1lz+pD81Y0q5NJdchhqrfo
xQgsNyJnPgpVYVS81+/rlmdqQIme6q2RHsCN3jgy0CncFXFDnz5XfNKkFrd3ZOS/
QadmJIKTCSsXNnt1YH/o4C3BtXoE3SQU0s/fxr2dsjFobAeTBWylK2oK5gQ1EGUG
G1Syfcn9dXVEhH+oahJRJe8kV4brFiA0KMgv4IPIzc1CxE+HML8Uh8hgSJ63cJmX
m+yFX0W0p6omgkUuSG1V+nshv08W64shxL6ByZwzsP/hwhA0wsRHK68TzpnZfMkg
ptSa8cd+deu4C8ttg8dqLe1EBVZVLfOk4YQGcKxWjiQRxN1jprXWtpvoG4gTYcvg
F6UvLV1vz0yxewLHCbsILShZCe0cWEPshQiDlCqUtvdr0sCXqDQuruTsmYIhbFOU
rq6UqbqsCDXpNEnSXKrDO4sAdI/4tA37pUHgTvHxk0SJDySFH2W0KsWVpGExO95t
w3OO5ykufDuwYIvK+s1bwxRi/XvSRNrtwUfmDsUEOD04S+KwxBc/+YpAksXqesJI
cV6Pl7840Y3sr+jfaq/A28wKiNWAwfTowixHKGBLSe4TRd2mSS/WftqaI8rTF9so
3Jwm3UvoYt1lTSPllee3I62Ve0QNpMYiy/aOjSCpkkBuloOcK9y311qs4M4kjrKb
dB5oGZoLZm7qCAaqKq4vhedWCpZej3qVhBRFDfKExY0q7211Iqur5cDjz0h3VysO
Xb75IVMAxrCBuzSsL1+IYk6tomJdLCdSBU8ZCDBk2nZTmB5tYH+yMnWpuHrQEjs7
ikRMVxwfyiI7EkqiEDNeUmnJt9mlD3UQWUNl+YGU9j+oloPnIgEC0wNI9x/ZVTfp
DBl8UoiXkXGnRAiJsGMeRi7KdJ0O1F/RguyKcSu+YzhUxTcQhHzUUf4XsVu99vua
zhFhZUCOTALaKG7KL++SkUmN3OhN8SSW62QfZTuKNBQv0tS5c3no+MkSaPMX9s71
VavOc3fM58jgbruf8g7rSt5+ksVgQD/ovwQuA4ijJyDTJcEfUILsoqDeSHFtDLiJ
AOchnhOo61tEklGi58JSfcfpMmpUvKBvGXQb8blDVcy4bD/bDdOsCLvZLgQZxs3l
pA/ye2w/tmIxISlqxCMjLDvfUMymDSNrpxi3tbZtFq7GldXqoipLj6JTd/64lhu1
QTb8+oXnsjrDBF/ZnDf1g6HPLZUGWj0Tsw6fDuGjnddgW0Z/6x4YkMFpZLNqx1P4
penSeklgC5t6BsD6wTwvhXL1bgy2kx+0k1tOmcdrizHV1/+MekyfqcvU+SrtlQqG
8bZjGYnoDbdwQlRR5Z1lbsBfKYY3Ic8roFMmvhV8JSAFh5+rrGDxD5lHjRaCAmeK
efKY1ZgdFwD77MT1MOiE42DDFV0LXIzJPjyUwnM1Ea+6lR6b6D5MrQwVtGL8isVU
3+PsIGku+KTrPQ0uhh2cWkTa1wSphYJKCsgqO5nLDjuTR1p4ymXh5n2ee126yL+O
twCB8n3sXeU602O3BCCKeA/jEAuFlRqPc3o61+ZUpLlXLIsNpxYX/191DSw7Fl6h
24+iKIL9lS4dUpbbuqFYOmqasRyXNU88B9is7LAlef/opce8z5i2yjEwVrQJlGuG
quGUK4tpX5aT3Zv9D/KS2ygZu9ZRJCvcAuf9drl2xSMAaPm9hoB5p/yuYaFDUg2o
+8dMVwo60UBbeTHJs2RB9gyG9TRWykZJTDv5LhkncsuxJUOWdojqe8A2MQI6xB9w
tEDAvAkdxg5UcSpPUglIrjNsrRWKuE0EOZOc2wTDIHClo42KwE0ZHxPPsODa0Ntj
nKJhCwgXuF1AQnvhoN02Slz7s3dijQij/kJaFR/oUw6JGdQ1kYBC8stnSzSR1sR0
baHMg7W6P4FtpxWABsBlkDMSxRwnEtS3pOtCC0Ca0lKQniPHSs91XM7PfxIjMtyd
wNReUuLRN8s4OZWX050L9ey2Mo+i6DVMYtYFdo34VlupRr6CtG09tYi2R309J8vT
wsGZXVxO3d6tw52GlxvOf7WnRwSTFFDgsO/+vXvKv3y8sHj8HBnVI+rZ5vfG9BO+
h6jRblbdTgJdCu7Ds1sDUieWUhxI5p4A9pzUUvB7OsqeSOecPtflPmJ9xGTTOZrr
BaPV1vmdfIKmL9IIv/I4VeUhbBRJuuXCdznWwuX3OAZ+/opbi3rx7FDVTWjS/7sW
O8NUGTgha9ZUMd7zGwfduR4WzU/YRkbu44H0xdgnysCDPLZR63zfXm/CIVHGbd0L
dlUa3KJdnTNS70evwgalVaGWduhf4duXcaYuZWfO1/5MwOYqogTwEl5pwHPnDqgZ
/HPJHU8U7iIdy4hcUTQ6vSHMDxYcx+XG7BZpf0aoPQHML1egkUUapiKxnb7lMUjv
tL2u8F6lxIfOANLhpFlZth51irhvST/FOSzp0LONMn7vxnaBJGbumoIBQzTsLOv6
0Yq5JF3uvM6yleviS9sOJnxoBfXHbJBlQmQM27+MWefxHagh6wDV7dVQHPWDsnzM
SLFqc4zAMolN8uadffApby+OsRjTA6tNiHBGyozplk0JuMYbwSC6viX+eHwgfpKI
CEsJs/d8FYt4rl58Dm8DkmRpUkpi9CmsNiszHqUAKed3fn0Y4V5tHuzV6Stbea7S
kdBs1EbdI77V+XqAWjLuPHYS1GFIqkyHM0ZRtYOkdgiGZEQxgm6uS4DY2J38qwU4
82KV7m55Rxve1kfAwK2B2YYPTHDa4KAvNvghXLcgTgxniomk3/6n01qx7OwIz7H+
kNpMU7tVR9IEYz5VdkVpm3EjWSYbKyXNhd6sG3qTvkkCftwhgy/qchc+8YzW0LtW
R2OSS47JXlDCvckwUwByu7k3pCzOvJjkdKhXVQSjo5BI/G8b8YyZ0Vumbznnp2Ug
701ssVT3ZNS2hsayHM2uwuBB7dxJVer6a6iX3Adx0dM/r6VCQCRlwedyzKbwIA/1
zwwkhfmfYs3oqLVy/vwI3jKk6xfTKYoYocEq9VCk0/hGPgPcjdoYf3W4S1E4nZR/
w36jZVTLBbiNQp2NvorVFGbhNKFTipfHOJrvrE+FjZ8ek/+HwdLJn9lLIwjmjX4D
CQnwrrKb+sne9LfinES0DyY3SnlH3KX9i8pwwf+qyZBszP4P1ejrQdFvba3eJF8E
GJ+s5jdzlueN47r2A+JXYQ+kkQ+f6COJ0flXg8v7VspEG+OFoZtgyhMq3A0ND2ke
yRzsBX8yi5rFxLpzaE/pdIx7+0GKRJpynW1s34IVc7NAb93AKSttJtunntSwq4Hf
ry77NH2hCb906UPoVpAvqfet+At/wTMRA5U+5nhLkYfqxwNa+9IVLCheLUPpMVN3
AfQkj9gWwfuEqzP6utQLd5o9KXjlPgvD0Z2YniVciBj9URIWfqRbz38+RuZFGKQ5
yIrMXLyzekYQo5HsiALudacpft+Q/Ce/AYZMuGtOd8khL/HEX7LPWWtZ5tKystME
b4OyRHly7H9075XZvg8eUhRFVpjknb6bOdgQbTZT+5bLUc5fdsCIROhL3532DX9+
EtouvytEaqDu35SO+jVOmUGIO+ANStNfpAOlqimLAMtUiakgMBxyXLGnXduA/Xd2
HaA97OCpw3biI1+0X8crDXLJnuT8UcnoCGftxm74lF+n/7IFxB0jb6Yx97bqrzCC
qGHN/bLmgr/TI23c50LouoFY1+yqnxyxsnFgyZXJaTeT/ZCP+PAbYjZp5MJQ/vRd
qqrGm3O/tai3vxAfSDBjLpLbj/ou2i39H1VL6dHirBkruzpJQoungXcqAjSYs8i5
GBqy7bxNpsdRZPMttIX6+cMXObldb/E2SS2FzUb1a0YbM0rgpu/reFeg5C7rvxjD
cQtXddQVEjG1USrvoXQiE7HQVAeBslGavOq4CElkAJqOD5y1jMmVXn28iSpBRc1g
cmQT0i1h34q0qunRxd7SGvubRpTg2k00QW1lm1EMa14XQV70WSrKxpP/IeqMSTaB
eDABEt50EZYimJvreeZZPfdzMhJLrBTJ7x7XHSbnghvOsWx5rlQZxfpedjBZlKdX
aHiQZXOMbfaQt23mnQtL/7idzutubENRl/rnzg+hruMbUOFe4FmWWN5kisVb3Fsm
ubwb+lS4mF8U+ty6B9/OWWkhF/MyFAdRYeMJOhCwvTueQBRlo14asm2z1M+r6bOS
TMCMEI0a/NPaFJB924PsNuDkpkY0eqgwHNZ8pTyyTAC5cq+eYDL+CBvaQEDJDsus
rXS49AlgPao2bo02YX6zPl4KLiizD8PoWWbH5C+xDGpmdqxpxKGtk7glVvoDdbX7
Ti132F0+kbn77jPBqaO79Q97dKfDfMCUs1KvFYrfKbQA3j6B4k3X/9mL5i97qmN1
AAMicIyJib8nZ7Vo/kPW60aXiMMQkrworlqLZYJq3x4cAXQcaEkvl2poL5nthDTh
RfRC7BtBrOyEcQbIWQsvdFwA0GpmaNwFkK0AzdZm+9SMFvv55NX0A5ldv0Rjt7nn
U2dfO5jvIYjSvVzh3SzMKyT8eX6xGwx4pkxR90svb1woKWB7lBY/dGzlYS0LvxHm
hmvh8rsyuZ9ZbfI+ILbYVb475yZyhgLNcikfNcibeA8wFEY+AbxSGHm7JydL0Us5
S5JQXtEyjORZjhA+83guAEr6PFW19BN/2ga2AAGPbfCbB1BURCaa4LG/i1DBpJMx
sDxu/9/e/lHHGkOZ8KCANBdTSKcS7fmRd/FRGT0ET5ylHBYmB88bzK8nksWJZbnY
H7Pu/EAOpCAt6/yflv6ZPPCiyDIDtZgikn9Xk0pQn2ZunpP8y3i8wLG2MF3xsRM7
uQV8vteKhwFJokn0h3EjLW5Of5TK7QLX+z7pz5Hmhuqh21w5vXahoRNQIfhUAjPV
BCukRnIvX/C1lkA+QefHlI2CgeXGTCzSXZd8sq19wNAAZz0/xBecsf07ELYYqtO3
lZMuXumOKWQkh6OXvhMUISIY8jYxcfvuyJz7yUC2KObn6PTxiRkxjFru6bTfX0y2
y9EbqbarWxh/Zns9a50cvxVxDrT6hBy3g1cZaYLcsGyeub9E+wkadzNoBPjXV5I3
Q8mB7jR2jT6bCiJRf/ScKI17Y5Cavn5M2SdXj5FtdK1pnU+8XAZauRTtzc31Us9g
ahmQ6VLxXmUfde4eJn1kvnoy0kM/ejsIyJgnkrocze8buSB3Epvs+FkWB/ehdKWe
deV3bfSguISO9EEQIXJI7eweL7QvoE135DhvMFGSYDaKO/IIxMv9gD+0QxzIWwRM
kCW32kACJOvO/7wNjZMHN/SzGmGvTmk6kZpe/xVEcYEV741I/H1CIwqLs4biUzi3
ntLZ7BHwZzLu3pS0QO7x1JPYUglsKdiGRgCcz8mPE5CVk2q4GDK4D0BiYkcAnPJT
WVQXpgFmqMxe1hsufzQx9aY0LkamVTYeP/o7X0ohv7gXPaCITV/TvpWikOfTT0qQ
G32e81okpxK+6l/lrSim+j5lx1Rx1Ja3Ows4VkRihuboHYgaF3TC30xW1D2s8PYF
XzZRI5E43iRub6FJbzVFycxif+fvpjgai7FspKJ3edoS/+i+IhYjAleD8SPPvOlG
1kuT0yumPt21qouWKMnGs8ThSmKJrG3YheQ45+COO/YRL60Z33X7CxXJIc2lGFQc
QGyNkM392lwoqlFNDRYT2v4zFJDrpNwLqQylaExCLbOlb26eZYtcKkON+EC27I6P
Nb7BTKaHLq+dOjX8E2qtd8ZEyQKChMyrzBhmqHCchnzCG1AIeeoJdg8ESqfYhi9+
6DsqK0h52y0JRK585XpIaZMxX9J95qm0zpYvPYdbHtE9ovAKcXnxGp+3aQ83tq2q
5vjUMIB3/2NsYKoO5kpCYZ6iOMZtLbQXEqRz4SmwUp6JNmy29JYaGen+06XM8BpV
`protect END_PROTECTED
