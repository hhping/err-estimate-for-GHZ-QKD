`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iN/szS1YKCARj2Fp3VErrNT0tYCYv0HBCLJ0OrdTuNNOJDWaJt8XnVFjrYZVZugx
Awi/Fi97MU8I5Z5xDOf2MuhIP9aaBhosWafFOX56blKal2RKbC9AwqsOp8zpfaG3
k4xe+vtLFmJeRWduQQ5l8mBS+rT9MeDHekoOc6Ly3/aA4HMmwrYo0FPw7AsHpO76
mjLDtzd5TvCuyoA5iV4knIhVEHvdABTeGU0CimmlIATDd4tt1F8bhmCD83ssxL+B
IrGfwUEqg7cQFBaY/G6j6xHzK5hsWdSaY6GvxWvHAOFUPgIHqH0fIBrUV0tUDsJo
zEVnYt1NZl/BWPuhbyj8yxvlu6BMhM6cT7Ti4QsAVZ091xH6puUQKsuzA82g5cKq
FYNC3q6DewwHphxFWj3qDUYWMNvfntVXOyI4bxrJL4uSmJnz+AcnXf2nDSdnMfn2
6fjlS/JBa+xbjaK7P1wBKrTILkLnoR28aQILZlR7M+SEDi3ugnxSCYsHaUICFJ/l
BDqwlUKv4LFigP61SgAA2mA4ZmWn3XSdY5BDSYw4WQkd1RsEG2n2Qm0WgGGl0c2n
jagjvXhDCFMHQL4MsmfUtyKrFuX9sdpDUlI8fVviDex8J9CHr9Rg4mIWPzvou1jB
3fDmxfqUm2d5mgGqNLoXfSqqrqxKe4mpJ2wbqA4Uw5fjAjQ3bMvCZld3wFy8lfzP
K7226r9O8wVIk1R38hK9uYL5lNT1kP+sO7SZfuDsXsmRXMzkjWJpJT8hh6lJ+ZsP
CzAd9SWL1qVrp5wuL9u/h9z2QjjFVH2nd81H2/2qD2m73NA8ejZNNVX2mgChp1Ql
QikBxcuKA71bG3jbR7xkT5urm6JuZ00frq6x9/+8IbBvpfOhshYROzvh0ktOyUlW
2X/SsDeZbanY3caCVKkyTA==
`protect END_PROTECTED
