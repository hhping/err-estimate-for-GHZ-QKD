`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJfTap9gafh4K5Qdbi2g9KPHIot0resJwLuzwKjzLTD4EBxWwG5rE3eC61Hykz5Z
Mz/65YCY2DjUCLYXLTwtM0N37OtrjpSec/dm4OQNL4XKJR8ym1664rZ2aGnHjmZh
7ntpZhXB6lMxUztJLIWiF3FXsDKMOyboKTKFHO/Y20NlHWh0XLz5PQMLWjpfMeyW
OjGV6aZEd8LTJdlsltRAJ+2sPTxA5jND+7nWxD91F4q3vBrTgf/3KG36YOiudVA4
nMmbCTkOhXTQt1KAyhPDGCefC+3jE5ZYSG70D8OD+ADr4tMUvI2j288ujv9KBEF3
nd2HdcBTfe5lGRqgEGIpv5x7zsFWH0soqABRB4AwSPA+sFDifl54xCbBkRjTvGsi
zE5tzFWxl2RzAtC1obRoPMyyjgel8WP+6wFzrRLS0vH4qYbXFKdnUelKzlbLMaoa
CUOHIBkAAQEguamvxHFeifZD0seenMf390J0BOAHUIdgNV1FQpuuZ3bK0l+QAWeq
qH5bfDW9wh5XY/a3qHxh3YKd4uDQTnL7Bvt7hTU5+Xov0leWWz03WK4Jk0T6K/+6
irdhDaj1GeQj0GgTiYQvi0/HRi2DkrXBjc5zEuIfDCqpwebSoqifxK5OiRbdHOzH
uzN1OyUHYtnX23H6TmBIWblbxW5T//hJqqQ1O1PumWUJblocG4eQzVHxMiYqWAgW
K5e0mH9kSCGI2TeHkgsrr0y6Zq6FhzFa+lhHl//we1/UToquzKRqux/Hzfn67JAz
yYN4PiFMSE4oeD20WymqvF7INFlLBwNVdqtpXtmugfJcli9GF3K2OV3fS61j57cF
EIqhW+x02AlMum5j9xNqN4sOAiWpZudslUdh2FVnLc93szVEOiz9AGvnYuHhopGQ
cthejAfZq7+aWQQ/qaid6NQbGFyootbwzH04Ep6BbluGemcK3NK+y10LuSiwPNgC
jIpihHtYQwAOa5Ehwdu2nRF0lc+zHD2rdCNpxjNekDXKgqQjSCOhHTKhbSWN6faq
mAclwG4MFgyeDvZi3IwJLEOgxkOYo0wLbPe8KwWnDMPdLTMI//zcegSxTHa4GKjH
cjp0nRF8wMrkVvmsG5VVf5t9WYb26m1H20THo1sUANqxC3EhyJuoFQ3FdSYJLWFf
lTH4v0bfQLqK0IeEj2s667N9XTzH7fNnUnU3KyE2QElplgZlW24UFxiCR2pXS4re
D3V6pbhSkHR3Ux4rpOY2pl57oi56Mo88lXL41XqKF9Fr3FR3AWB39YhXgVFJTIqC
N4LI6eSXHEk9k27RP2KOL1rAAi8USqYyM8Qyc+VYQwrU36RRxoK9XQNon6vHjaDK
`protect END_PROTECTED
