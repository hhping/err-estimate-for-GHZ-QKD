`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HOia8iDnsEgLLPlXUyIbxVFlMD96pfo51Wm1DbKe/5qfM7Hax8zutlwG6mxFO6R
3fNl4B8+IZSOp3Akwin64hzVN9rQsGH80gW4H3KgtixY/HpmtK+RKAVpqzzOr4aj
2w6HqHWd8sxirl0in8cUehZCYIAasSoVcwOSzlD+KwvP6XCZP7TVbf0Nh5peCz0r
/S2gU9FhI8oPzrZFZKNwdS/AgjC5CnfWUAiqvlKt1192MCFkTcUbV0+yRzz1uhGB
cX4ACkLs/HzRGfdF/Js4XnEdxHGpcgT8TyRVV8VRlzOnAbcpgifgmuBcvKMTFkWB
qs04mnCbDmJfBB2unXH89e8F31dw7g05Vi7yJqJpIDyQU2Bg0t8T2A+aJUL8WB36
Qi5AQUXcwG+vUKrOtSOGB5wsQRSTC3R0UkFASf85GSmfcXzuN+gwJVvzUZnK8myY
txRGShc32MDlQrkNm+0QxwHx3q7ndsTKRIDKEdkPRVpS6kbkFfLpHFpdX36p9hoH
4k2W+VUv1XcbFrkcGve3JT7r/L8vSO+7Z1einpmMB+SnyXtFIAJ+42+bk8brY9nS
J0LtLJgT82sJxdUHLY6UqTWeb/ZinW9r613uIaMxs34lYQk2YGIoc1YL7G/qQb8s
2c3KBS013KvvO6T0AUDd/MLD2weENs1+szp6quFQbrz/v3kBzUFc6Jwg7oDg/RjU
bf8+z90Nm75qEqDEjR6gBNIsGkwOWEuabBgMaQH15LCu9XdsNbaet11odKM/5nVt
NyylDF0CkKsgjT5MFWNYqAHYxvbFSRQEgJulxEG6qSnXmA/ofhaXuhCTrXJbx0eW
xseTB7D89AcLwai0BVbRNUgRZ4jouA7FUE9D1TpX/Z9m2C/4w9D3DEm/+INjc64x
V9ybsGo0TbSySWe3ghtPkAnx9gOsabMTvzYg42/WG73A41dGwS6ksMDBFCYeRxbs
Z+jghu3yYpTnf2oMQPsHqty4QV4uAp0GjBoGAWKHgCY=
`protect END_PROTECTED
