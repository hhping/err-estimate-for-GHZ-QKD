`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDe03LIvLMSkAmjNdyDX35+296+gFvMtqJ1InL5HWVVoU5/OA04R1qpwg1snbkcr
t3ujHaKP990zcrAdHwSuQC6EA+Ejewwo19Kh/o/NqM0dOBtiUFh0ffcbIdBYAO89
cwdDmHmMWlf7UZq3Qi83owmi9RNmu44xkku0Xegi/cIrff6uqnCYIkAnUPXcKYaG
oinnD6tUwN89CkNdzTcH9f/cv1kEPL3D4CjWc50wfRUKEtfYMDvEN34DSv9ZLzPn
ezUPrpxAuQm4H7HZyJfSiXCkHJDPAScAC6e83H6Q4Fh+P8Q2g1ZPzzvRddQ5/lax
XpPEC968rjqZD/ga4g400SLzUjCtJTye7LNY1gCvnR2j71f7CvYPzRhxnlDiDTgS
2jUeaIKEB9IKUEFSzRgJVabwzOG7Uoxstv7D97q+5P+DlyH7llF1MTP70PN+sCaU
20xGjaepz/+TycO+AWMaA244t1sCY8kY6fpzqOIJkCiUw5A7rW/Vrmblqiyt7SzA
V6y0ImhX5MVNTC6mkZ2bHmi+dZySq2KWHCcP6NEUmnxcsnGFFMoY0Zt0tso4he1m
lkupZ29XjpJIgqv/SEP74x4ojDsLagp6wIG9pRkMzUFuM1jKLniCdebNV5IQuC31
fWMzZXXlRD94LNk27gqhIPGjI3UlVt7Hm+GFjW/ugUNAtfbtoJ3Dt0CNwW1i3UYg
ndxtANufnv/kzt6P0BtH2evjEwvWQFyf6AZ3RbscRG50qltQgrXkgJY5DABG9AQy
7qb43lZ2RV8IwknFsSWHZllBqqzMMUq0OCtV/Q4qLZ4v6bZGdPWoQp0Xn3ieTpmJ
kcTCQZbYx2rPKfoWaXcToM6wpwCZhUC0BEnONMLVHA7gqMkICOmSZRxSl8nhI+8W
PR4cE2VRlM/k6INhLiywEqGokCRpbaDrm1UOQzT1N+TlXMAiiNEYTGgfN64zsFQd
Ew9ZFuXG4B0zZRdtyJaYzn9olnfN6Uf2FRQAIord1FbuWkcf6NNHpmAbGhOCiF88
XBXIClkotQrwQBFr3Az0bVqEYIo+ZfFH9jzLNauEm7LdD5bTG9AF+505RMDprsDw
YQIUVOOHcJ2yUOvw/nvaRgqFLLMZRwkD4Q7LQxKcC2amCuhF5g2irRm3LAUS39TH
q4wS5ptS+RG7esPQdq7npPcA1otw+6A6kX38IvgevarVOxrSxPOfCPEOAdmh7uOQ
SMrKNE3P4HvjhNRclqKUD8x4ExzbWsL0sP4z4ooNyEZUEqMpznqtjZzck1dzCtLh
NvrXQeol8+JiWlcnomiCXvHOZR13ZucQAYSm41E3a+H56VVy9MbxxKcwmGt7DAYR
dV8S7zOWXCB6/e/Akt6SHYyN3KqgvrLHipIQE9pQL+5kruoNd/mE5rMG4D7tQMSz
R9WVzxeISzW5dspqLwajOs45m95F7sEDgUVPVAJmfEQMgF5xZbdS8CynmfmkEbyK
tWH2+E42vGdfHekfRazv03xvIsaN4DmLfW3pB7XaNdAyd26cxc6v56dxefevAGoZ
SPbthKx7pjNUr2mHqGi2SCszM6ChKb0vxep8tJ5zfypGhpAgfra4QhkC/sD/c9yz
RWLx1aMbY2EP7s3TRDVeEKTmaAXkAvyGrSgOVU57UfszUZokvoNxiSzdvWIoDOni
kMia+FFR+WshMM4paEN0QNmEDbdYsVC1wGXQPXLxQMMQOsvHCyw8BXa23NRlWSBW
6sRQEWdUwHUMs7cFN6o330eq8TfV2ogF/ZieirXe91WGAyjx7c9SbK9dvyOsIbyz
rdgqHVJGPZ4htJ3TpskIn6qvQ+rGjh4274Fouz9FLMTdB6hY9NURgUm0HBbPKGPq
kx+f57uIxYaB+t4QjqlyScSHOloJLjzWh+eCj7bvLNc=
`protect END_PROTECTED
