`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RL3gUE3rXtktL9L/rtTUD73M2DFiB6xARFyxxs3ka6Rz/ZXgGc0bP5psaP7HOl6s
bQm10nJGfynyuh+EElfPvTb9X52z/1sFxaVfE2Pww3B/bhSGXNQ5LlTyirGBs/4o
aMoXfdNEt71xa0d5ndaUYrfMYLAmS6Ms8rY+lBFVFf6k22K0kqkTbgBq2gl6Vuga
p9DCGQ8W0OmJMMnhopyyAOJuQtCAVPiMErXvNVNHIiu/rz5Z+rpGxdRWilAGg1Tr
G7qBRQQd94jeQVkDZzR5sm/hIcRe/GJw1PR0xyM5r1Pcskde4luMze4LkFv34rWd
YLTG9UIEd3EMv+5L2PUqcCvkqQM8lQEHWtfUZvS9QsfPy6PGtIaqDL2z1/zYLE8l
1/7a6UduRCTXhQT0VwG71cIciTY6wPg+LMwVypMG7Vhhb9SkK8QGPO1iQu8JBAGB
FVcKOvxZrecsLQyseKKPthn4bRGfdKjFid8hyYL6cueH7B+VVxRzbuKBhaw+Fdgy
UVNeQQCUO2kig19Fj8RF/heHQHjUeIM4vKern3CPGxdSCFcHaQmlq8mOhasM5Tj0
lnBUP2ZD5IMGkFPqc1e0EfuURjZYvaSF2jXaPsBsJH1GLeGiTXNGQlLXnVyc1HJd
hv5M0jCPPyfaxpvcvDr+3aK2+WvTgFzo5PsiGFMV+FAZDOVfLZIGg4GUcs6lmpFa
cm8WBKIpyCdPOgjq0Zp/RGgFTGrdJVSC6pKVLL4keuLMjMYahxKtXyxmdOBGzpBW
GsyaLx+IoLkc8iLug2j88BTyUaUrMowURBaqBeQPPCH+5j59G9zLMYWneMI6zOwp
mJQaoQcNTEgSHrt24ezNSb/5+WLbke/oRhdKY3flR/R+Y7HutZ5Rd2URsxLX3jnG
fTCLfFoo/aivv/NxYzHEbj01SuETp/eQa9I+uTR+fyrIm8puHQt2cbvrVQ8NQyXV
MNT3joqxPGujuQvldmn0Bwbdlu+n6nTnWesrd8tHBndNeGJf70fKP7mqg2NDrfpy
CUOfDQ7PTk/oKA/RD/xyUw/RpxvdPkS8D1NL5fVHYFxQScpADfh0c9wbgCsQId3U
WMATh/Z1ntD18Zl2v3lzyJ9BCcAIYagTsnNtqJiemqYyiWLt34v0qxIHYHTbR+dj
MIr0eQvrmxE67TuGJN4WI5undcPGbRIhATaYSx4fry/ol3RfhsjdekXlAxIhCBYS
nQsSsbnjYXYRjj9AqShYXOy3PI3HwyZsAagsTtjeyrgda7RIut5W2PIhLPh7iPXx
Js4b6AgcblAt9Aaju5hyvAp1efJ9uTqvp0m7zgBQvjzlKs3RvIanr3dYmRBfjkbv
y04NNbMZLm1x9URgE5AudwMm7VOBgTY8fVTA/EyrEKFH+pCBC+7I8EQwdkyejKLs
pDtCTOWV8ENlF4fIibz9FXXgjROaMMx308Et4F8sWIxfxGhG6Iq4c0wtaFysOgtY
6LkAwPPb7B4hfiDEGlPz7BdcReoaqOsTdvai81fu7LiyojdQtJ641saabH+8zO/X
h7ujoQfu2mGoOknQqq+yOjXrsLGIBe8UKUMy9lMChSD4JTWYRPYzkmYtn8rnsuTZ
7oT6zz1IiLrLETKKuYphOxRItHvYhkRWNmAu3ik7W8j2a/duXDRKNj+NcmOr0d1Z
L1HoHv6s38dd7YJRfncjjCjOG05m5CEtEZ+dvObrgbov3KmpyzSQfKfQHInWTQGX
Ut+rm7GHISyTrw27F0eY3Wfx0vuq8MUI1DS9mdeOJbPNW2kfk3YsnYGFZbPG/yvH
wmYXzR6R3nMM+v79V9xwx5g4MNbhhacKqn8APLByzdpgMPrh/eofKGQtoXXQFtCT
s7DLCmxV6ZQTGAaPMHJJoN17riPSAfJLenHdlzTs+EtsH3gS8LDF+jCavodimsZv
7iCD6g8j33XZIJZKhsaBpsLrV4WxGDyQR0rKosv/lgvQcipLnN0PWG3Zry4Vn+Am
X1ocXoNnzzzIhaELidgGLrr3SBXk59ojhtjz4QiZSY6JF+nKgs9q7cpkhJG7ecGn
`protect END_PROTECTED
