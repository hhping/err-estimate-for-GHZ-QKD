`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiBj2CVIByTDAyiWmTHmx4xTeYou6wlHCiEsuRuPgS/k8AALas+eA+lCCTgpRSZe
6jp0DDtzAKJBJnxV5lA/NrcmDv+hCg6WfQ80p2m1/w0Rqc3fdJCdB6HsdHpVpNsT
wb68ItE3ohqjMhW7pKiyGu248iJOS8mfprUkQ/zIVv63T5+phEbeN7ANUXT53uJK
MMqTRtIrnehc94qxuRRFftXo81gOUhesnbhB0NJJ86qxIeg4lb9BTYbGqI4vOZ9/
MmubfJYBZ+ONy4v9za1FAlOWdHZ66UdkRxeM+1PFCO6szoI5zdG3lBbDDEY2mFrU
vpGM6pkQZvoqHyNNVm0/LD4cVodVhX0zaw0p6iiOTqD1jfFE2Gt5d4ww2eJhMsdN
v3RSNRSG1XJBSdAHMNjJXAVQS29xeyL0Ao1YTMhPuNJsvVCxeTzSB4K7i1aX2NuN
7ZfJHTLtsRWopiicH9kgVhsNu7HngAHcjydI+6qxjxA2mEBA68corcvv554UWuFf
dVMKXeCtq9J91KUyTgAEqh7kaantyU6ySMpDrHQIip3fNdfckDxXfoaok/rOuL6t
fCBL6BtUF57AN4oKQeoBF4itZkE2U5LxWz13qPFkT3UAreB83WWkJ8rTL42QCqdl
7ccRfj4j/u35TfDGSa7ULx5UHgjy7M5MAjX+UWxM634IMQmS3caq/u0nECLc4kCX
LExBdMRza5I7fzUL95iyXNAJLaUQ69BEus7hzavawm+CKWnXpCUEZaXp/SqxKhBL
nLiFKrILU4MHtAQfSFCLwKxIYT/OqBo0lGXQy3PHXGya6Ov6oCY7xwloignPmzvr
oesDz3SzA8ylnE37UJ+lqw==
`protect END_PROTECTED
