`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lHUMMK+hA0Y5Y4xrFfJUSqzUa+Bds1QZ3rPoh38oIn0g5J995KAypgsQfYUULAT
EGPtFRSz6Yjxd31DtYJFAjpOIuu+MP3sPr5iM7DRg00AHay4tR/DGXaF8RuvT0MU
snmv25bDIVOmm4rtcOovG0IVbzUUj/TN7RXgxokxC46bRNCkFf1DvdkFbW8z+FlY
RJO4dWXkgh9lO008umh3+yToMIyjp28EKg3Y9jwPKwF9bVl3DsABgmvZdoijVSTS
WfOv/OEg5N3ljl/AfoJv9z4GB0JcCqG6JQhOJb3qMPUU4oVOWWaMP82BMo4HjW7X
AE0KCdoYMFZbR2Q1cfeExneDHZAjO1rVx+QIA58sIY3VkePK7GjMwRV1QpmBMGFm
ly3x+g7E5dd+cymFdiEZVUF5vglI3impc6f2gVGPQRjM55TtTxq94WXMsioG+6a3
hm/oFcitP7HPO0QaTtp011QQRfei117afzYa+nDvNw8XAW9RwnlpM5ZTGcJVqQWC
oMkVH0VhB07GOk7fq2G8GPP+KFDijyzp+dDnC79iek0pFcCtQLyqhgpQE178bNk5
YgIOMbvZ6mCFriUxtjuGZKvaEvvWK/YymAxxPs2xezZGEZQsxiuWWnEex6/lzfGT
IsCDMxmPKVuGLkfNOf3sxpLgYcz9qftbTtiKVZElqBipNvMw+MWooUmjrc9iDC9R
1nOU0JLoZVCj4H4pQR684SAc3kPgkmYRyxCAewkagkRCedYVt5irFB7ijansUnEb
9r0IthN7sZhIPjks4pul9V/H++N/z2pwkgnSAcBjmUTYJ5TZo21Lh0k2D3i6DqxI
DNWQuvrsIyI2tA4gofg5XFpiG3cfOHk4z7ShViCSo+N0wm1lkXxRtkj7Dt2pLtj7
wA1eBJKXOrtDVsir8GoWU90W2Sh6is0Rcy4wW9UwWbGw36I7m1YsgS9/sunELS2u
8uzJIjofMb/GcYBpHrOOHQPvaMbVXr+D7DCHp4GDaDdZRjD327DkhTuozAaOdlzy
Y9ALz9mgUAAHcQUTslXZwxkSaMAbcLGIrv3EzGlRElt6XNjf0LY/25JAqB5d7kql
RM0UsZD1lB8/e0xGH0nWhQpPIAcvH1DdZ+YWPCAHX/uONx2gLCLMUWuv8ELI5+Kl
ocFg/jFoEHzRfBdxk6B/lIhxFdd7hvjOdv6RHPbAHZvzM6ldA1iBRbcUiugTDVe6
/hUvAFWDHItE7Cf1Tn5C7qH032+XVO2oChfByc1wfAPc3RqMsQSWzbLo/TXTiluH
/ts965m92Do5S/1z9b1GQJTMsQtXn1ax2wli99TCdVOdos9MWZIK6Lhm2jSLSJXx
MNWCf99cFa1AcMwehhl10ozC7Nmsb8Vkr2LCIKip2Ly6kEqYVcNYTAEqvi4FYkyU
qHHj025ZQW/AUcVIuHA90PLRahs969bKopdm6yeR6WNqoNiz2BzWERsINhupSwHb
MdGVW/DTRfI1ldKBzpq4QA==
`protect END_PROTECTED
