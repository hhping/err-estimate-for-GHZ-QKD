`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0M7MhOpMFRlGrlKiqwsvdxxhVgmnDxfSQB8NZz4eycelseX9DavmApm5lmCN24I
VJwOylL01H3Q4o1mi2WW9YtTFrojEZGLa8+qLhcC3f9Gi6qSZB0UdBQsI6zkiIa7
9tb35JkkC6xTe+GorYalWYSy4dA8RWZuX4mx3b6055IeISQeTlysJtE6ko1xUiao
kvuFos7c8PocFQmk2oE8xItmcqoaTXYr3VZq+BR7qpy/na7m9aULIVh9Bzh552Ct
gFA7XBESVKhtvc8pkpFkqvhiSWwglX4bhySdlwmw8oW4R6R2c4bjJ/2gzl8A+yze
cQ7NCCFR0EtvmmxSsNg17TikzmZ6p6oiS74xgpkTPpTB0Awu+KkgfBCWsqJCuD8P
/NinhSP0/dUiukoVRnoXrVRDO+DzhouK1g/iQcxPNz7aRc5hza/dhmjoA5QHc2nd
b6wubo1GWtkgLag1Ow4WvIoAmB5NdWgQu2+ldOXNWOz/syIe9Pu+uez5DcTucTzd
xP1UIZFTJqe7L0nffmOq4gnfdF1Z+KRk9hyQ58/IWzqDZpbb4HhYec/w5Qc8i6kM
alSpt7F0ckg2ed9dq3eDjERW9RnXdkis1Ch/6/WWahe9EV961oAbtWcvVIiXh2e5
L417DNn3JYcaOG+EQMs6bJ/IsqlALvGO5Vt9hTj1YNFpP7MC/PxsRPFF8EApBAsX
2o2iSkqJth/o2goC7USZTXHJZc69GIFOw66mfAFVN65TLWjMomQ8deruJphbR1SC
2SF+UM3Sg/8cT3g/BUo96g==
`protect END_PROTECTED
