`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Id3ZXg/9bf83uUmmdgAizNTNr+t8Lmyk9pHzQB4UvUkoxErrobcRXh5BWjKmNMQH
XsbgCOFfTfNJlVnS7a6SLRY5xwoWXZMb1LBDfzESkaTTIPJigfw7N2rYulc02WHA
Wl5LPIRvUISl/z7tH5taoDnH1yr/HYsFogtORGrye5ItPSr932Cpx0L2bM32O1KL
yHsozuDvV2aKu0vtp2h8l/A5t596Y1Ob7n8wZBw6NIqOTD7QjPyzcDvOLrZn2zIZ
13E91FNvdPTzUbJtY0EexDhJnzne53tASp7s8Pc5awKuPO6Xny/lx0FO/aaK5fEI
qNsmfhnhMENz4Fz9TP7JR2T4yfWTnlzYeiSIC/n/2vWk0zX+cjI7eXEYOEawY7pl
l2siT7OTJPcH3tyCq2TJJffZkK8mmc/yqsKStHNmxNuyDtDLQzEP1K4+VTHpbGtg
IS0koahSJswCTwhIzPpUawDwV5e2sDbXs1nLMXdizTUoaz12xBTxsfCWk42T0WVD
+a0mNCZzmm/K/xub4/gmcHWKPu9HgtCswWRb1JwkzzJsAsZOZ4eESqVhE0XOHkch
hUIMH1+8KB3jh9gCOdG7dXKhbKqEcvP0mUOQ7S2pA0GObDX0g4ytZPzpoOBCNmDg
TVb588+d03hwWVbMpNieM3QvTVcp4hHnoQuvkrBdHdvv3MPOZOcQw+bPO3FZFoFX
bGm5Q7S9hlWabVtgxB0q5o+WizgwZAuaPub81ud/ohhXhRqDty+NK/ji9mkUMOyD
I7j0sY6zcCbW+SI1n4M4m4sbfHly/jO9+onx4k+LpLnUuo/aTljJHNRhPlu74i69
dP7TG+AfxNsqtsxq3P/yRYRUZLYu6QvRUABgheZUDQz07EjlM4ezMlZlQS9alU5a
PMbEEjCy03u8X6aw2G27YHPfa3KizpPZhV1LiJUKl2WO5qK4HmcA+1tlwFQgVIJt
J7GFZyjjvkdN6VHR+huMjFxc0nXkP83oC+RX19Y1wml9NJBGp+L11eqXIKueMM3W
zWFJnAvHC0K+BxJKKu68VuaDIDHPPxV56L9Fm2mkh8TIWPPIAHfTlzRh7XhfzKUB
0xLkioW1rNmupnVlpHTeBJSbgKxWMcxMAOdqTDDfdQCddI8alkzE+HCu5cWzQBh2
h6ZZ9pkyKI30afgB2qQ3AiWp3WuiyJHv82d3qopuCIrxfV2KN8a6Pi6wskDLUqbs
nTVXl4NsXPuRJL1HCciVr5T5dolYcKBdUXQoaUjOBw7vlnhxldefRnWM5D6GOTDA
K9FJDbPY2i2Kg1IOu8NBO/0s0H+ExnjllacWjYllTR1+HtK37orAXMTb/lgqhWfY
hBMy4vZcZyd4j4w2Wr0KGsacHtYuP7XGnWkiP1vzM4s66D03GF7jwrnog4GSrb81
YaAABG2rJeyJJhnb6ZIuo2RB9iMeqBiMpvOIsfTVKwH1CuT7jGnwOFjeDiMYCurb
XCl5RfigtAwYGKyDS6rDSx/ScqLlhE+AxayFyKlWZqPtTMy39f6ALKNm99RRyHAL
SwU7BzsC8uzdzYV39wqsSqwUeAHgtpLyJYSeAMUTBawaSJ+n791WypoYq5eH78kc
tHeD0Op/AH5M2GeXcsumkwEl7lTOeOcL5DZzpZxCluZGAoY/cFx6uz0wqZchH5Da
Owxfq/RLeu4TZogGwTHrIIhMp6bU6xxBaogioqAqQtgef9i9h7xi3cTUsHqQeA3l
`protect END_PROTECTED
