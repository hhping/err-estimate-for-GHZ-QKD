`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mm8HsZ+npyo0jfi/MgcIFNnZDTYELc7byU7kJjVhd/l1zv98Pgtem56eZKYnOb1
Knk5DuYaSPgqSlRa8Mh+m318e/tfHQvNM2ZoHr9/wrTB2r82xKqLcPqG3Src7Drn
iRIoN8YXdaRlsNiWMpG0Rz+NEK0KbyJlnM71lTjfqY8QjjYwqdELKRHdg5qCZOuW
nP7yGasL/9HnenQ6yl/T8eYoBtttdCN9NG6bSdasxxdBKY70z1atPYEmPY74AYT+
yF93QkD+VowDpXmLKgznwRfHSQl8IFKfqp0gP+cGTHIMhRWIKytUWJDI6ZlFRw7u
VKNShJsIC085MFT85F/7ajyvAkui/bA1cO2Xm5+8fXuHfGiqXC9tpChKvB/a++B4
XCDXIrnMRpRoKxkFA6n3LONn0GDgsJi7BOi3yYNVDo7jErSeIQ4DtchTNwecB4Pe
/3Xqr0Z/h375z+bU69osuGvbi717bICmzPhCpT96JGBOsEXATNmgpvDL5PGQCtJR
WOH1pzBBcxWlLz3phLAJqZ9C/rG4rZCWN0VQMkFSIgET/CZNjJfGwX4g0Lxgxa8s
heY4ORsQ8k9JniwuZyG1+gn26tdt6KiLrUXiQ+pPEx8rzh8v20rit3NjKu4d9sze
x6k5nwHF1urJyWyO6bOELXTldOeYR9b8pP1UYsuQXtgHMf2coUSkWYoEKSVPDQiM
GcXf9vLWlXZWd5DiVxk7p9Oojytgzyv3SPYcv6TwYIP5XAOnd1ew1sTGcFqs9ax6
XbEK0y+g4lWpWq30NgX2vcqMOUpsD0UO82F3HTXVqDsJoW86ClkTX0JW0I5lyzKs
s20fYjzFwBF7kE5oaIVBeg==
`protect END_PROTECTED
