`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3EOUMu7GURVrXCKh9GUQv9fV3PuDH6uYv43w5+wk06ipJbgQivpu1vn2QTerweP
tXP2R/vGtdpCEK5AFl9trty9NdRk2wJlcGReIgZkSkuvVbHifJi6T0BRszYpCVPx
uGolLijBce+HAivL7mFC6mcALwvkPpNCcw0IAPQNhLDBTYZi2h5wShiq++oTEf+L
RVyUBX180Vh8cav87pTlg7Wh9Pe5FIkY2ziDrAZLqr8A9wpCoN7qT0NkBn5xls+D
QI0PgkAsJtXH5lI5ynVcu0JRAvydgWWUBwggYbK85NmkE0m6TDR4NkdwoWBEhm1l
Ah8ZL61hJQ0AVHZe3tY7J5SPGUA3+RRsN9cyEowGb2HHeyx8R4qWpBGpfZO+n2AK
QS9oVVQhLhIH7CNsmAV8M8j1yjtoeciqoH2chGxHb+6YuQ5cAKUBZBb9HrLsfip0
XX/LG4IKj2Hkf6ElEvQSOaRDp0Ymc2ZqvK5+m/LHYvhae82H0Dr8bZZ2R/lAJe//
0lf+r26N8BSe/lT8a62iicdt4+VDV+3OoAb1Ai5KHEmX9d96aSuETB7PLmRILwvP
gypTWhiXNX2E/Xa8Izai8lPslyOxzyv/Buyr6bZkd5KbLM2uKtqcxzBJHUZXvqAC
iGdviQc2ZDzo41NggaRmaZZmmaG0SNDcPPY3KlOYPuvckBvLN/hMXY0eytIJtZYB
Yxnt5Pq1AQwQ2lmZM8T+0FcjOIENmJDZgu+rVimhOFSlybX7zWPQ3oMeHT3b/YlK
vJW588O6MsnO5YE9JvWbCF99Z1o0b5FmuFE6ftMCB7uFsEAYpDVAT1Aqd1JOSOrC
izFDVqYmKGLwsyO/JZJaNx1OdPjVi/jX/m8S3ypNEUci5iZ+YzwQDiNS6jEiGH6v
9zfNEW10vJVKGc4lCmiF5b7zWwN0Bt9uZaSDNrJKbGmPLV8IS0Q33beBUJJjsr23
32HimFjtCf9QhuWU118uTL7ZTSTZ/+QoUdw9Jeb1UnZR/NvM7xTbnzVSbiaJZXpd
T1Gt+BEyPo3uSHSg0FjC/pGFu5MKyLrE9ImUv5KTZd/yb7exRZwofvgmk5Tx3g0S
Nr2hIWsedBzAICzFzzW2FZi+xRE25+q6PEiVc2PWQBfIUiNz/ueOWQD6F642tCn6
p7eml3G9JG3VduIGFGRdBdfjFu3cMmEJMzFT2nfudo3//z7Hkba5C9qrI7xQmIvt
I5YF7LVgV8LM5l/RmBZfuv8ZE6t2V5mEHX+n02zq0OSQD/5jjCDIwOavqfdz7qYE
bwgyOXvKzb7QL7/+PQLoHYfNZrfSEuVqtoC43TPNLGHLDNRzDuk5QwY/hewMYLQD
QMVOb2oPUpOVpnie2SlcEqtoscge8dR0X/WMciwh9vrDxtkrTJCk0O7kVOTcLbhX
wq0YEhbcZiuBcimMQPcTwvBrGpulb/vg0hW4gPPBYeXrlahgisJlgSGvPoFrVRcD
BOb5DG12oHJ/6D6gh7phPmgyoYAIamq06s/HW1mk2kl24p8I6GZoFDYDgcbN0UBZ
LDOZ6YhFoj/3Ldv0Bgpv82E1XS+cv/O9hiqJ9fdhbWKZP0D1DTjlpy2D1iGzPmd0
ggueDSBx7tYmsVeT6TQWIXayw4W5rT1Ao5pEiuXvIiyOPNt7jiZzD5xtg85onJNc
M2ZBRpqFqMNlWogPgYkBaGBdMgc/zZnb/Fphu8fOhWOaM70VWH2r8pWjFcGon68C
tVX4T5+kY1GOsFkSDpjB1hoSz/sGs05TCd18XVkRL82E+Yxl8yEu5pIPYXwOYmFt
STyAnKv8GLbykiGNU/nBP1eAFaRtTQxS4tRuxGlvxEuboBuNV4UQgGprrIsbspPl
lI4ziwpmHd1spmlRKMHJf/+mp9zuhSx9CYIQ2m9AQT5KmC9wVNboJt5h32AXNo9V
HWIvNnyRTUjMeTniwknRfAJ1+xYgFb53C2YAb3390T1gCNkPtjRT7iwEru9SXwYd
SroO8tOucFRC7f+6Jcv1MA/eALOOG/VylyL7g39h/l6BOs031/nk+vLxxSG+lo6q
UMTCOG7Ao5KVYAAZDpsmhx7kyk6ZYxn+7HVorar2oUSpFMaTI1SO/4LR9c4lAjYS
K7j3JK1NHxV7y2+fgClm/OliBtF1wuvIxekFFAuFt5fGXdhSwx3uW6OzI+zq4bsE
R84A1UVIquR7IhlU6ZlPCgGFHlvpPivXtBxbCjsvzP6K2ZrucvtH9CUaMaV2aImm
IpM+TYaDcK/C13oGLpTMWqD0TDQmDZRT0KV4N5bboJlbG8Ihl5VOZTzoW/CpIwqr
Y2oaOinZ8HFIws9sEg57cP/jBmvxtRpV7m7T4DJY3woJ1ZrO5QN0pGgy5x2NlNpD
BCVzg4a4C1PsQ5kSQziQ3RIfp8p3lFZ41ZoDsNKvLfbO1aKPjdjiAw9noOPdwJhd
LTKil28C7DzdQK1VJ8n7anT7CWLStec5+l+Y2PCGJFbYUhbLDKkuAuq/KKEAQpPL
WMW81gdDL7kTu7C6OKhdWPNt5mcaAx2ho9/ygcGPiqI80NlVvgfLASw+XBaKVwfD
EB3gGBFOBsT5kf7o0O3nCksZYBJhXU5k/noZqmWWE6Faz1ZloUMWzPyB88c30j8Q
J3fC6HYZyKLc2XFqMljW9W1jY7a1Y5OCTJF3fsTtUs5Eawzaq2j9pX4CWaaGrUwS
9uj7Ao8LoZSj7SflNsRcivJnTdx0BTf9YPpmf3qCpHjApsApcFnjBKk3oFlMz+k/
Ndt38rWVFRiMbiLoAxeD7R7WI6Qej2+uLizfAsD30gXWg5lW94XqIjtlWbviM3CU
v+P8+TyDSsQPS9pb5IRnC7cChyJeb5c3YasuqzQrc5ILh7uyEllgNoNJTCgtFqSw
YJPcabkYKQs6sNN9naeq6vWWauMa4lT2hk+ZIC/SOaCU+4UCIHUKUWEDqlE6kfQm
FL+ZzjHESfjhAi/AVApiPwgH07o2MvE4p5H0pgoU3jH7V12D1Gi0r5h57EHak/3t
vQu0wnO+UUuF/NCSo2FWgA+hzFkwxIH3Q3z54o4m1n0wuwqbXuBjvy/8Q3xvj5v+
22KsSbPumSiwOf48RBxA/e3nI+VZtoFYEam1IVhTGFHst79sI51xAYxrPIv/Ke/R
KgL0USPZ3NnbSG/IV3z1zBIzFXNAXIE6yC7uEmf66mNKtzohvlebdkUDFO0nzQiw
6Q6bmBOLtGVJBGY0ob5em/GmDUi0xUzIRE8hGkvOa1KTZUbYzNGrXO2kNrDzzhPV
0lr1Uisv8NV+70+xkv5vyVWwO3TRzFBZAb+4ExcMNFwj/BcLw+AAST6XduERMS3l
4W7Qo3E+SW64IdO24++RFuRJsVtktRRvEjZaRSEN30p+Ltfm4GmfxaTzWcUDWYSv
7DisZCNSjTWDjR58FWR87zqGjjdHkPvmLAHUe7L9K7FfR1fdoyfYVuSXdyMdN7u+
OR6AsRDhJ+6RIfnqrUkua+Ut6InDBhWKKROSop/OhAUbSXMqoxIPfxadwfwtCEH5
6ppGFJEZsO9ufUSgFALWf9aV7tTJXXklq7cht6Qxd5xP45ZnR04JpPx8a/CUQzfY
+HaN/tsVC63nETlqHBBA+0bGMNxg7jKq121xGRhRJN46RvDjebOv0RApeFoBFGBB
eWwcd0yE6bMEgvhZ0OO1vwnpqCFNVO+I0KqrKVc5sdsxrcgtkIH+Vtbp7KifAXGE
lsrKVyGoYhhYH0AYxYJpjFnVgfww0dkt7oHAeuvKv3vm1w7R66mcJlKaIL1y6MG2
ZOGnBJXrsrzBfUqTbrx2jGiimle0h2G1RttGfw+5YPKP+RKTMiGlSuH1Qe/HjRlm
UQbjjrzIWcG0pD3yrVIOur2sVMCT5JEToyJFEa/espLwXsOX5P/SwS4Sppsybwxv
4s9B7zTgQDmWEEaQgjNcqar73vsrRaVjN2MNwj3hrm0XXOcaZ9rCYNpQqkLJAT7/
EkewB8DcxByMqTZXt9rSq0E3zFrAmhPZcOdj3K9XriMWVoIbvaCKjLJqWdzOsgoF
kMIoz9WcXK+5YlXORPBugPPNu9i7afvXOmG+/Dv8m0I7rRQOuLm0ovN/uUIRsBaB
zCcl8sKQlENYz5SFvjwW2LDwJG7ZW8tgx6y3l36ynTryfhiLLPZSX2xhPOoAMN78
Zu2TBuZJ6vudQQUjtybGY8g0bi12QzBWXTURpsMECCflQfjRwDEzXiYa2HNkreXf
P55DBwvSyfrsACXNBqC4g2IBwpQjoNw0t6ie9V/IpUPg4YpNRnLehZzQUBpmJGYz
AB6uOaWyRLse54/AkU/UImtOm/79+IbnjGzCSXa4YpFkkEe85d9b6U2HVJu+bJ6M
DGSD73rgDIDHya8SbtCwHjefmbilN53C5RcKHWcP8qetC+0zer5o5TK9QLMPwFms
XzVFFV9sw7H0ZQX7m+ISn2OAwVupxTi8HNOOmu8cD8H7Vkp/XgRSyru9PCs/3kmJ
HaQJw5ZcF3jcOj4cAvideFfk//5i7p2ddoEg7xUYD0Yte8Sma2avuUfNEJaIkYHq
G9dHuRkYIxkkoTXQfmVGYPZUYOh2IEsXtBJG8fsnerkwlI5qcBFoW6IZNMik7EXB
pmT7Iiuew2lssXuQdj9cWYJw8D3L13tKWyNh5SIrJUtjGH/ULkqXDujnulbBNuj3
KIQx1qHFosLqCF95e8X6LbvVCAamNL1/cq0DNcRFSgKyeY8Uq/MwrmZ4iSg56xya
fassKPUX3rpNVn8tiBcLrcZzfshYrWjwra4pWdEtamq9QP0YADsT3NUQMVGGh4aU
du9sCtLUYzicSb4goGl7LMkmEuOyTmr1M7vn88To23GbXT0/XaL6bJ7zQqEtrqXJ
14jyc38CK30EwOVfzLfrUwUgQ8aoNoTdv/gSStuBju6Wt93mB6u72jiSkUbevYHO
VA3L1y5RwsM40uwRCM68XeMLqGuz74AGysFIb183dPb4xSVpb61L2pQNWh3kKLPv
Vu1+jG4MHkbjgJO3h4fQ/BARMyh8PUwmoHyDNHz4ay5j+TwKV3F8ZKdsxfNdv8EX
o56y4vjRJ8QlvqOq953twERp8GkyIxytINa5n2jLKWyFZ0+Ee5Fn9SEJ0wfCSTGA
nSZAYDViUouZwjYf3GEIMrmqnJmVgvobKCkwoiCEw/4u0JJ2nMVTmxu0XneaHatT
agfYefjtWxOpscMHD57oy6FzFEonkJ5i1LrT0vMsngtEfKR1WcpFP0k/gZZcAGSB
rtUunRE8x2sOUuaJxAIuKjA+viV2gN8IeR5VrRm1Qttibqg845C9oDvUmzNdcW2O
yfJC3AcyStsU3WzvMjr08GSCp4yMYHy9pizkTLZu10WQHlKmKYeKxkkWhbT1kxH6
WboX2clT7Xo263FvdLGge0ML5ftNwIHIZSkLjDXRY8EVTkC6sjsCcvBItNN8JaQl
X7l5GLoVW+WKCHINDbT4X6L09JkB7NgOETU82rFBBnirb4XEWegjcCn4cVJ5le+o
M5+W86OeczDSmff+vBsl2i/KcitaCrei/iLRCgT2FvubN8E1uhbcykzKHVFvMhjT
JYdGIayc8PRI8K8/vPUP6U+dFu8rB5VU+ykwm9qx8I9ZfKONOvopmQvS1op/O56U
`protect END_PROTECTED
