`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
amO2kvxqQxc+RafA6AhRElRston7PEcrNHrir4gwOFkqN7EX6cMBGJIb5qVzxRwA
eribU0kN62uoEnokt+g/vJOlaigv2MpMXJscF9HR7CIhW4wWBNh9GrfRXBIQvSj3
JUwBVgrfdmxRYcDvstnBFXh8LopXsgdJrSaNlhXg6cWVaNb863rGDXZlIOFBKfsO
fDAnYjldWgFPU1NMp9qB02/T19OgFAB2Xwfek47U+qH2s2bzBdgxGv0nlDeeaZi5
g+0KX4WmG2onQMRz3zLaN52AXDqOSmk5GAavh+hdVjMwN9V2nWa30zYj+Xim9jrT
eOquEzhQmkTF+O3bglx4xngnZo4dg86ipP1+opFP6Fr9UiGxnHjHsNJPNvXqJc1F
5dJHylkcvyIhhwTk29D4lBb1tRZBiBSPve6/ZJekxBgacUpPYllwP6xcuGGs7v3W
+6C4TxkvkQgFCWj26lBDdHe7OcTguZg+RriLsCcALcUx48QJu5fHIHX3sRh+FnK9
hRxJE2aMTUqFjEx+hxnNs+dtIq1FVMoHnMq7/iKd5QmUBpcbWHqvSC5BlURtIf6h
AdKPcp4UB34UQ8B6pOyThF0gBnIoS3s2DMoKvetavlYhDJ/Gm9ZMX3/WlxZrDI28
czZFIXGazsqrzjjLSiJPiSc5s5a+nuN+L1ubUp11iFGeqlMOF7xlBY0451Qa1FMh
1dSNJvbIiUdgfXuHkSxqu9B7etoys3DHpgwW7lPRTlEvb8wR148dO2wh/sUie8nC
o+XqvdimoEB/TE2eOc8I25SU1HYnfzgpgTVXlhqE0O+1Aj4UI4+kIEWOCfx9So1F
bdPJJ2G66fME9Al7t4J6bvCEeksS25VL+25sdbEkAVCo+WqDItzqStV/DWw9Ohak
nlEhtcvdr43Iva+ZPSme4hW45314zUUydNDXDhqYrNyDXGeU9Ox7i5fj8YDE8SyE
0O7fb1J/G+eQVZ3lEgJNw3c+pMOh7sCL9M2B4NzMAT3/A1F8yUpAOGgum/B0jQ8L
DbyBmb+C6Y0zeulAT0sQ2Z7YVbCyjbf7lDF6ksCUneLC6k8XTxEDbyVazmqMBJus
`protect END_PROTECTED
