`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uxDhaH70pLBatKP11nNKe/ICj+wC/SCIA2bxncdAzu1QPNaquoyvnqK4cF+rKpOF
wOJUKoqf3ZDEW2mOTpI5bDU4DHxVXnz23mfpC6MzN6vhaj3EwhlonlLciCZg615y
yfEMXzhyZUcFcT895RtucSlPC6Jm/FRZo/X1OZw3hsSRLAYik/s8nZq+F6nnsEBU
3rNnEFtlZbNVPYcfZ2lAERanXet3vJ9VPY9KhNW4QbWd1XFgKtnE7msZOYyUiIoa
DDz/5COOSyW3bIq/D/TQhuVJa/5Gr6nSz+Lz8BtDAhBkbv2wFmxw4MTWgI7Sx6wG
7hCKOIEPhte+aO2+MmsMzdaP6ZGVbNpzTldI6kk5VXioRK8X0QQpjlBEzqSY8pSF
`protect END_PROTECTED
