`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/rd1NOmdO9BQNqaj0TGIukTQPtPwE2fVCSx+xPy7N7VKq4RhPd9hSdzErje0vXp/
GNA2j+h7Z3yP5PJK/gQkvWXGMvgs2fD9cSlT2syr1cTOB4/LblSWZvUePzd4Ze7Z
Kw4IXmNZPnEDTBVCUnHIqVDbIXKSqK9+kXODbXID2FKKPBmsDJ6Cc0qgEq9oD+C2
FV8AOfBvka0ghEv5HtMDL7nNblb4hyRq0FONuo2zxmm1yGZGIMr/EQ/lxDHBRg7A
kw7ptOoq+NiWGuHK0SqJPcS/w7VQQXqVx/jK7yB0HXKzbkBHcyLYn+1zsUBEzGe8
46Kij+xSwrxftgJoUz+Z8ByBZru2mVW/5zjAU1d5CAYnbK10yxEH+cBzni1QavqT
6PowF2GP4/q3n+bjWfZMyYUfl7lVkY4PPOXrTkjlZwBE85Hpi1l1cDtMv6ODUybB
8rqYSvl31V5S0wn3KEKTDIqnnUCMhBInG3EYqLCSPwUKSr7s3wN050/1F7uYQKG3
kFyixZBvN3E1CXD6hmCogSbASEEK6u59+DCZyQ4LFlB3GQaDrUUKJyiDFx2BClnq
`protect END_PROTECTED
