`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0TaW9IqVVAG839442HtN0e/A6KSsxnPldPh8hvevhzj6KQasYt0y8U2XSoNz1ZTb
bFDg00qYRFSMmA9QFa7/76yrXBiNEX+0Bv006tHW+yO+Z2MJijL2Piak3QQNkyWs
25s3UdrXa6Q7Ql4fbQq1+4+CQ5JN2jwWEirCnQU/E+LNqo+2I2f1Rs0Fx347/aeZ
eWYz+U0A2q6yHTzRhSggd0kZL5temHfi/DojzxZcFEoFY/y1xxBoIgjbl0280uyp
7Ql7OfH9gZegXczNjzhxxEz9BfZtmXQZEOA8d35mVposMMPSmcBRs9lvyy5eEBoX
5AqkrkPVtsPu1aViSYd3dS+Jy1kIMtxHIakO0TneN6UzDXIywLOi4Gshx9vv/f31
KUMafNLLG/H6rk3/yFI2HA==
`protect END_PROTECTED
