`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VttKVn4itDnD8XB/KGgFNfPbq9TwEPPXJHB8FMV/mR06pHDhf2U74zDDTZ4VG5jq
wQ/H5Uj36ISPf5u+g4rCwB6w8h5kx0XwN3RRxFOMVOzUTV9bViRInlsYde68pcdQ
d1JMHpFTL2Aktdeo/twZU3GUgDmIy9Sa9mk3/OpEgAXphKrsijlvUNpNVAP32GzW
u0Ioi2k3qk3cRmKq89U723oRvhLLpckhS2Zof4S0wpYmmzchdkK4G3qNPzbsBy41
cxfMltgqsz3JnTrWzDUfYLBhFBNQ0qJG4mKbYLGx4Iynw+CFli7p93f3096I2YiT
Io2hFN1ZtTaMCE7/+P07kzYNX8MEZcLcdW3tIlbuTK5w9opmQ8FJ0wc8k89woYG4
CCIK6hOTUk15tptMuku+bGIxHQ0zWIOsTEtjihsu7HdimHZax9z+lCQq5lPhED/8
EtC0xrIg8Y4GtwVIpNoG10Qt4Arxu6/4PACxTyfkthNX6VICxmxEskzXjSaMRZgH
hevS+OC111T7nfJgywb6rJH7Sfx/o2nqXu1RlcXjFeXM3Av7NqdNLoSLJ0Xfj19E
k+Pr5v9z8diB+xgqUwkeCKiaZ0nzs4I7+yaHx/MbJXafTXzK9wK4pzpUuTNSv3i8
XJdsI5JHmQx4C/lA4eypYiB+0FXr1bOu4Vr320rzNZ8=
`protect END_PROTECTED
