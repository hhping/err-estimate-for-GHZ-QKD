`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mQw/foTctF0FMyQ50MURv11ZzmtCKSiF0ey4mtyQFyFkrBO/xvGVinYXP3RDlXs
KJmGND+ytLc8yMZNPnCkNJZeLeG4jK/NB106XUpHVPTx5gC75isVyaYwq7l9jiTm
/LAzA4TvXrG0gQdzn1j6QohjwQnePbdBAPwtOEjrUZek8gkdHh6ZrGhG/d5ZilGN
9S0Mvb1bZLb13Ntb3OUVqrFFySm6w5zfLkUaD0na9qb9G3M2tyQd6CBHxW2v/i8B
DP8gzdz0VQ4lHdI4/7zLjZbfW8sJjotbUyBZZH9TTCqZ4tmLPGFGjp7LVmihIavp
kckk2SKmfjpJBJr1OOnu4J4h4xRgBLMml9DmC2l6NIuOHsbERvyDWCQKXg46kPdL
bPzz9uZu+hgsFOTA0qsL9PhWDxLn4UbAOow4pgXkWMvMjf8O+0soBa3F9Jcq6X74
Fz3WQjDbEQgg4OJFrk4vn0DWumobA/+Xhzmu7oP5nMim8R5lq2vk1jkd5bYLvS4k
YKTL2XeLVjXvY9jRgdnPQgYpnYyCyrOgezHjpIxmsN/NHAJKc0/fgPqRa/80B5xt
maVwYa9iCDWaVS7bcfPIqDTKoJRwbIa3F2ZbvDfntbZoRhTPdm1wv2gGGtN76a7N
arW2z76V5ahJnE+tU5PUjKMPBdMZOa7GOrYffG/TCYQQ1mMIVq3hM5+iOYrhAHNy
cgWAngYN7hcV514AAVuJ1jf8J2R68RMmc+3bSWSdRJL2yeS3Ev0Q3AfXsltt00v4
rahbcCPp2oBSmhE/bKaoO2bqtDeYrV7cWaF9Me+dc02ulYiw1tOLjsH3QRoC71UH
kgjuf67f/HkdKg3PHnV22S3ubls45TJxa+WEwj+gm1Bg7EEXcLWFfSGafI7Z/CKc
Rl+UMXjU1N4VhDC9bidLYX6Cjdch3I9MJeRthcBMP7WqhjqhR/AKPA/WGlI8oeR4
OkHMNd1dslUJbd3P81SvKvh+FyUzkL+1s4CJaA4SbZ20fcC8khNl9c+tJeJXGMYu
7DXSkAiNPnaJuqF0Kbc+IFUixU/HD1TOg6EfbNHWBVZQ0Zm/eGq66fwxkQcGGI8u
IRZn61VXd+gpksYdK3skLzJy/BTIJE1Nifsr2aKGAY+uV3yDwhtbU1b8uMV7lhpf
95Gyx6MxM9nskhsUwVWk6zNJCwhtk9d8/7VXdJWNsq4GIhVuqJbZbgT4DReBP/bk
edxjQzd+OzwLqG3UxewvWoXbLZS9G19cOWONwUWy6hp1uIHkzSG+BsSZnR3aEmFO
wP46Hge7a832Aq9pzrv9lEb/kz5IVFBNmVYWCXXbcBrqMf/5K4RGMZekQSKGodkp
i5xJar0a84Q20DH9VCNFP/DtUgBlwFfAVzMcx6qNzmns9JSYQDMsJwZgFabja1gE
P28eInEGZWyxbm7/bpmXwkNuLhDRyy9YC/kjXzvwARzf8pyZTBNJUUx0qK0XVCLQ
hdnZPClcp60ZqNJWYwfPXSgXzT+RIfJLroIfFgbP0BVqxHzjZy+IXIEiApr/D4//
G67LlnNtCfoF8xZuYM1rKbpQrjmK6srQlYRISA9i9n9tqAs8uVoTwmromqBA6pgI
037LcwLg3FxXvv5tRTs6PyOOUO7a+Cyvk5sJu6FPTwhbw1VwjEe/aYBWHrkTK4G8
L6j4A3UqL1PXSO7YqnQ5X03BzfgXsfxn9FARluh8cgDpSLHAoRCCVIUtyW6MoQel
sdUOV/ihHGJ3RvhAy+Eb+TxEo+7TH0ljw7oRFJ6aDg2i4o8HeaoA4OSNCYlpTOj2
fVCGgjARGoPf43PMuDI7elvW/N5TJvWRkTqOcnd21M0DkEPAfbuHSI2S+eRGKWMn
A7FXkTBTnnHXpR3bwoO+0/tVRpq6RWczBaPPi0AC0GsOeayeVenHFJl1koYj4rs0
FnSo+4HEC802dw6rkx6iLZ3DWPqbqoTszOTnrki6wpkf504iy803Ia/Az3k/IUAM
D0uEvUEs8sYti3mcMAj3RwSCd0hE37GG+YFTFcAviRp5gnz5VtJguDmoEEYUkbBJ
XcNlUBCxGkOyl1dYAtewvN/uOPZF6JHkpuPsfJCj61IjLuv6bNeMsODVOJDzuFUa
3t2b4JtBw/FGas7v9kONR2440LiG9f0jxscr2NDXzJHjGaCbnA//3kVIhB/+E1dI
S3tCwSSogXaDUU/9s2NyudQ4Ad5StGXfMeIyeh/hfsvlhr3EwvWqEmuwWEMqw9v8
QIeDZEzOHgzz97S5iqmAq31vaLeDUHYF2c4h+o1iRH05naO7ok1TPGGAFMCtPTVY
KSVGElpz6NQm1pj5wxB1yDBWQjLgGrGpIofeNdOSXSLU1PGvJmJiD7Sv/6FomgOt
Q05LmxqO+UTvzU+A6LjtayFuvZ8Wjvi1hHUbUzb3q0Q4eOxhW35zpx90AzCAhkgd
PBIxnGppPf8Adk7GoB6aILcD7qnCK0dNQ6oyNDN7Hn7qgSAFKnkNyoDcxFoOLWTK
dr4+vJrTHmzo5WG8k/pxI2Prh9UwJhBcMnxBwNdDXHmlM8CL1/Tw+3vMCtxKzfwC
YecKVNo9nw47R4niwPgYePxImIEGpt0K4rpwWpqrPg2qy4aAcYyqMYRnJSBxBLV7
ejyBmzObv+WCZPqFzC5y2WFwuaVIyzb0HsCDTff7PXqwLb9MuP8YjP4bROntq15j
NaS+x893x+FtFD4LCYXzZiD3TJlqtKSYGZt7HgF5LpbleZsvZP/+ph9xxWf8Q7u4
PJKbN0JsIgTjM2ivVjcXhDFSfV9xdDOxhThVwU83kIVv6H8Cso4DAVHfBMgSKkdi
ouq9cGVWQzSwj+SLU7fvkghOF3aPtQl+8GtdVn7Pv3mhh2+N5jnPv0uIF+JvNPPH
Sw+Dr1HXoLyk2zeb5W98AZr9bfJJpONTOfDHlK7LNMQhqgcnbMj2A7Emj/0Aie5+
9iXI+1ZtjufeTZ6kO9Il8r8HyhSWIZTcq/6uDmjHQTwwwWQZlO1Yke6SwAjgcp2x
lhj1wIEuDTebc2aiWEilpwPC2fxxgNFJhr5+FmF0X6Nw1T/PHiA8pq63V/GIuiNx
SWmHECpXwnZ8FCaddKS1ePAj6xTMSyffKDoN54Js+7XGb0TlfI2lTtpS+joH/nZk
HXy9p59OQW+lGcVdgBehMWs0ZU5p6z5unjlJX5hRVIycvmaJ/wIyXScFvwo+xgsY
uCRz7/R4rtEQx8fAo7mYTEcwwGcKf5riPV67BLDBBQvJkKewnA43yAMLEGxnt7Vt
ehUenoDnWsIAc+sU72iv3abSfNjw4qNJJ+SB2IWwH3RJqr9YfipxNHrCdT6DsaHj
RGBG5UqP8fn/3wICdn7SWJcSBGspS8dQo8MGWT2iTe7vZ0UuqBD8UrAe4mpeDNpP
6jNCRlnmPq2B3EiqWmrEb2dLi2fY/wuKjbofEEYaHrqpYSxPhQB6G6w9xmzcH4nF
DCuzoGhBUd5sMSkC7h2gOq03Xmt3G0xxet0rYDiDPLaQRajVFzFYT75XGbMPIOM9
lKFpi5ldOU4H+s6CUu7StjOVlv0olx5OUWquPeBySN8Y2muKaTwbFE6MJjahJ+4x
AATf+/O2EIx/yXHbnyWdi1M10q1+uWcDQpStWQvC8XeIdExbq1RZVN7Dz4Wb0ISd
rgABqLcifo/AjDXOrFubIPaJktA9pZAc3L7ot7+S4pCE9mUqs7zcDIE/fH6mJcvd
rL5HSGZXhmH5I2DcqXiFquZ2xpaRo1XpfWwfEZar30OFDTUJ4EPLmi51JOhTJAqd
wo66jc2ebvCczW7PIw//c7Oala0wDf+RnZJN0kc6MwOSTDuubUwmwxz5dhugsGJU
GuCWsRQDEIaHhzS/eNE3thfWfsRWSczPkcVdy7JK1H+gIxKRo5GnrfnX6+DTHY1u
iboKW3peucvLxxugWgsbagDsEbb87hsZ4Ed9vKV2vWwtO27sdK+A5RSBc3nlHTXZ
/z9IWJS0UvSGKTfM+9ckXP8Sbx8776PobdbljKrH7vu0JFkZRrNdS9hg/Svwao3J
XP6APiGV7TNThD3LTtniPoqfkpNAHbVy0kDSIytkaSXLODp4kEHtGFgbM4r6YWeR
srrgMm5YB/DeIz0fBM27keA73xhJOK60Ju/Gpyknrm9agH9+7xG269rjkinq/03Q
Yd4Ej8ZATUMiZX83G8/EQDVpIyw3jHFTJYwgazs0XY+1BAy/OWxUeWl1sAlxLsNl
lDHjk1n9vGWO03mLNmMq+Co5UrLO1hzZSCfrBaZ5iFEu37kRtFC3R02Zk8PaBbi1
os/9NrZ3ljfRjlebSsurZ/7Kepo6uKyJag7KfiQaLpdfgiv3mcd9YxEv5SK5QZDY
NGDjKR22xqjKHeh/PzxFq8yI5JZfn25utogZzR05PAsiQPo6vD5NE9GY0xpwKU1C
P9QoPCoia0MK5qhnf8UPTeQ3s5o9P48lqP1xH6YSBKKkdNWhU3GOWB4ETx99K5Yo
H3RzXaXy5FeuOS5exEpJpon8ExmWrLgT7PjK5sgQk9djS2NwCPgaW0QROzTiWwQh
qHzg2nzeVLtumtJDyZHXz/2K2TZhkG4sNDJgvQnsgOPdwg4DyxVl2ERBmlGdI1Dl
dFo+rWWH8/D6DO0UkEMvqSexUeCVdJ+ESlCdJuj9SLO5I0RAqpACPkNo7tqGsseL
4VAim6czFUelTcbipBXGTAZlA4HnVbjtpDIDSdPqA2mBG67/Fumxz8nxGG2ifWem
VoSlsFieoR8w/P7nz5Ki3xxCBpW8j7t2EaeBk1pfTcWXOAqc5M6cgLTFoadJD569
W30aIomyqpiq98No8zmy+gm5LuK82qxM9d3sw3iqolDxyQ6ii6RqxrD+Co/912SE
//eDnZIAdEqk8HpKYbOAgF2Nre+vj805/CiSEIdV57G65RE4xMnTQd7GmmkdKF7i
sQrZ7KkDnpTOVYkAB6Ekulb7m8D9SkDdT6pYMZ6Fppb+FTjF8800rQrV8cGLF2/3
9ei3kYWE/rPZOCXhYlql6oH3yBTfl+yWbQCdYCt6N08KKGbCipO3PsjLkcodeero
J+dzpRK3+U6ErICCgiCCoAgIyIeNySPd+ecBxticZ2OwW+mPiakg2LA5uTzYd+8Q
mXcfpGkfBA8lPgfGamutGuBIrhOKqOJl5dEWgXrh437YPQ8MjauXaLQBcjpwnkBH
W0Y54XmFZWL8cygZ11NWaOdpIk3Uk3PAgWqKKjqe9A6o02xTYLrmrt84vVLu62o4
LiPTUBFofPxhXmsDH1M1rXhEpegk512FwMIjhDD9iHAeIsRAdxvTL9nxlvr0TQlj
RPnoKZXUEFjWjR9yxQBr14YMAH9Hd4AOQ+iyjmfefn1d91qn+AeHHfWWCE9IlQ88
rRVGDcZlUv/Nya/61CL/t4JGolttdSa9M5vseCHnZItaJv5QycPaq3qGIF+Ji4A/
tdOLoq5yngjPfV+v0fKY8Yt3g+q+FM6VeKApcoREooU6U8XgkK1SSrnnIX8XeFqm
QRI3egSkoFwNoHRB2D3vxixw5LkxwMZErrf4htY/SBMG8nBdDVvGVWPlBdSNNYER
Z1ACxDuC0MLLzUVBr12+fOk+by/v0B2wAFz/sIwlxpILVAmsP6aGGdi/rIHid6cK
opSS2T+GdZ+5Yd3qdf3D3xGMNVrdLhPNrzkjIuYMkUZf6Zcu6uuIAUG1LZzqu7Zr
zG524Vo6aKsmAhA7eyCjUgm54xK6baKLSAvvyDAuPZNk7wXgXWfZsqhhXt3sJrnT
pSa5GChiPS5j1Rc0jz2h2zaN/k9SXpBacvc3+gG3OmGzC09jxzDAzx1FpD9r+eoZ
0sxOSoWE/ghb/njO/SkZJ9BqtD7N7obEYtV5yjpB4ncJxSig/uKCkVC7M5iiPUSu
GbwqGax1VT75WXiRMZnI+/3C4lDojgkqU+AI7HTA+3yzO7OMi2gxdXFSDSUhr13O
WDzBlR4GUyMP6aMIfBiiTsRc5EJc53O35OvJMLBbijxqfp7CwD+/jV5Z263cuaTp
8THkMTYZ4v6zUlVVoYj4ZJapcvcRc+tZqBMT1/Z8i01lml4GVzWjC/sopJhNo6Oa
ZeZS9yFL3pNcsex6vkCUUY6lhdJBprooErs9BtM1LZ7XheudJmiEopc3FO5IRqrr
A4wTbZzsA/zgTjQCWXxE5QAkqANVY3Foj9iSdPL6r2GlsIc1pcBLAM0+s1QKrH+w
HHZnlfYyD6TkW0PGN2WxVl+fSNdmDWUdNYbM7/hot66WdeO7DERaer7B19r6s85y
uM8gVr2i7h1oOzu2a+rBZm9ETrMeyVwKMwdu94SuubEmZ3thloXwfxpc0NlxmrfR
kJbRMcw50kGjoCSrBl+JMOgyM7OKthDYBTaGt5TrlB9JHyW74aOO1QimlmQ7/LJy
XpGLqBIw9wOTxRohq6bNMPuNqADnRnlKRIK1IahLBMXmmRpGWNpMiMlr8jBKY+vo
DgA0eWoD5Q0KlTvz5LexZ299U/fbkVuKNgQDT/ErgVAiWgtMXy0hT+LAGTxFNFKt
9cI4X010SZSWxe9i9BQFjGqnxcbzCXSBYqhj8PiveG7rW6fgCyxj2hxPZeoxtih5
fRKAjjbi+75pBRe8LbFpSIt0b9iLVSBPiGLio0MzWLfWU3h+reSVMKN0+rEJqUCV
NxllrjG7+MzKyfCD8aLp4Ne+jE/HN+dhqkr0IxnkKJBamwknW8g0PdqjXvSIES/s
/qclVdC8Q1YUp+OAexUs6HTbwc/ybte+hkvltMmwvQo3pNfcFSmnMv4KnEUJQCoR
7qNvZq4pIMHAqZb9n2KZaO8bbB1f/+AhggR1oOmSGDSVbqzybxyUSpHhRD4to9HF
aSyRQptQPXNSeB7vnyaER3+yetSn2dTdJE7GBY/gnt/X+SdNRkdbJtWCefElSGMN
mKM/o2Lp5g8EqwyHeo9y95uDUwNyXiJ6RY+dGVz1KSALx5Yf/TVauhhsz8hY79DH
LFvZDzyWHAgIFGG408NlC8UGAsp55CvyMkFLEXoWmY8bhYclBfep65GthX5tRpyu
opj8+NzWuyd8c5xBhJfRT7Yj0+ikKuza3Y/DIo8GhRH0rUtN6hmgeGccEk27SJOF
i7Muq/CEbj4BS4k4yauFypixZOIW/Z0FMEvxc1B417ZGeI8IjT+3ts0+6dYWxuFN
MSYPWRCoEFwi+t/JxvemxVAnwVk+LeddAVdNo0I+Tn7FbeLreUp4cj2iEcZklk11
OuV3qVpj+m/SAR/4JK/jFTklTSlcY0ji5j5xJ826SWSQAcc25dFHwa/Z47kxTGwI
WZodHNlCwmHjL0FCTZVjBEVJPDnM9Uwwb3jl3VwBeXvI0nTv8Pt3/0FNDadz/fb3
bwqM0GrFlaAhPmCESWRxxrHj3kgUzaK2NLaKQJNhFX54xLsOVDi0GowOKHk297EO
3AKsvBARY2cxOnXRcr4j+2YnV7vPpA1PNNwiCvVnxQWZ+UKXnPL5Nbym3WOsq1uM
xKpCxjaB27gSoUtzvqXGki+ZWTg+kXYwawJHq2Fd5ggPiKPh38LKcLyD3MKSEDTO
sXFdTyMzwhTza9lOmF4eF3R4y7PUewi2NNxRbo0Tig/niofWSF63okrMtzyUyC2X
A8y/FiPygXtoMriP4GAOW2Gp0MDjv/k6WPq0RmIiB4hcp1lm9fe5RbqK1dD7NDt6
TKzn+4Th5NROzz3zSTJI3DWfmCWrojMdeNEWBJBbSI0U8gvfw0FdaeU+Rg3MlymQ
IcL1Q/s0udnD/9MwHAQ3EGsfi+2Iwn7jckhMoMwhcCXY7E+SgDZvg1RroQhUSyM9
9lE1nhZVC6IPe6NSEXf5uSJwzT0nRkcbIcQW5IxaVXvcTSdIw+IWC+96r7LaIBMo
VXYgRttJF7vTRtl57gvlm3XwPuwP0u4zkNgnbUaxWo+OcKwCqNeOXH+5kKIDUkfM
N3TD8mZxmRsyV4e8XUf8D15yM+lrmGgKHazfMf6z22VmoiAG3YWDUckYqazaqxP2
/22f5oDeWXPGu9UrsFKDUPZCjQo3N4kw+9ZaNQjiaQT0fFtWqSFv4/l/KzxY1itc
XQYN6o3KV2E+UF15EwNCvaKzHDWusMRWwoybBW1HEK1EeRbZ36sLXCVfmLhZJ/iz
kfX8RSMsGAy4zfp4f9+Hg5Wt4buNHwh4smObFI3jvvmBC6tX8U0rirToYrqUc9Z2
iSF0OnMkevqGqQw1VrYiL+Fen6xktnGpFqpATrVOSOo5TVEQXjVDEMvInH8t7VCh
eT8jnhMGhaAvH1zgWjGJ5FKKkGUtfZV4LXWTIyWCvyVrrbFcC3KiqIr8WRNf0N9S
IMYwYDbrVK5vCtaXVjbkeBLZVJpGDzHMQ4pHJpaHU6FRfBMHMqcpblNE5ZoDaz2X
VPodphmv7iFTwUwhyNwGWFQrJjxzuHpsUzVzM+Avhbt7MgBFE9Sj1Zo1N23RtsS5
L4TfV79LQzB1z/gk+dZzy7P9k/LKyxwAslkMnUdsTRB3vIOH13qd1c3t03hQfD9E
f5+NOpz6fMKGyjIucj59YPd+7hvI+t6pK/+0WcS0n6ZJ3lMR+B57jnwHmGql+HwR
Vi2HO8kcb1T4bQ0cX0HwPlPu8PrIU7aYfwijVfsjy4y7bff8/0cHrlQO33i+3b4X
nxjtajPXuH04K9pO67mMSQ8EK3+ThIm0Na4gJH+oNC2V93Pim/eaVqYdRj5w8p/T
QyOQQMKbIwPbNc1hQr29+SVNcZ6QTmcN7Pa0nV3xQldmQdFBPRyYVmN2482LRUAx
S8om7DPHH+lHoD/8ytA/W9IkKYWuC8NosIJUaXURXxQzmsBLQP8mHvrLOxXm01Rk
GaXlHHRvWSturIhAA/xMRhzgTmeMq73bHaC1VEbQUThH+Pb+gHVz4+DSRBGo4ZyP
ODSeys9iv/Xujb9IO339tjnZHhGHRyLy7F5itvMvaYYOx7DqoamKPvhh42fXbxNm
6k0Jv0C6T1kEimeQsmrXoSgBvg6vGkhSTepdSkIfHNRinNHqYwxIHKFtDFXBFEjl
5qLnHxMEVQTyjMiBPMQtib+eOZb9PHTfYKohFT3rvszZcvQhUAqo2ZyyEusA4rF9
W74Iaijeya7L+d9PUt14U8lAT8gvQqs7aTgB4fC+dR5zrIIAAb/+EdsXSHu3sVQr
z61plz7Ejiy9mC8Eyq3QwzojE0LOY/TGlptn0q8Ydpcowz7DcGPMCK1Ou4JzGB0k
ox8r1WpGOhK2GKIDIQyPRbqXqftKswp9MeOJWfqiG3JIQzHr7DMxP0a4DOPSLmtZ
jMQOrB8JUR4g3zuN2P/m1k5HZcZju91ZwaHCoNQmjJkI1R8RHyhfwQX0OcPNpX+4
RKPnKJmVLwDcGAzDuInmHYPOJUng/aE8NTub0JPNU6AhByn4xJ1ZNH/g75OMsyqp
QoJZjP7bf6qoBoYhYOwpnpX7pf79schZyEfEthdwXk6aVrbeTPLdrjbZp9ZjKeil
H+ivd95piFPSN8gs/hO+/WmHoMTwyOXPJT002I71gnseK2xaBy+H0Reji+TXZG4U
QWHk5Na0RFxKJDNotVQvwx1MdFOvmTmq2Mc6+4wyjHQhcGVuOIRUVAJpk3keZSy1
tQG7vBtp6dwwdFfTQ4ekBEdMC/xqdwtvipWhMgObnIyaEfi9ji7+jUWx7eszDTCN
5T1dRAnmNblt0oJhJCJKENtnjs3svntGuMNBIkGZP6+SYTV/4KYG1L897wy4xyHW
f3IJmCelkkRR9wNQE8SmMAsJciQc7l9znWJkH6SehtzXa6E40tY7Dxb6BJSlXSPR
tgxEWO71WP2NuWUZ5moiKpVebG2YM53bblaS6h9qHPRucri/0HNwpsxqazjbHmhe
SpccMZdLL0uOl7chunoeL5yHsN4+0ZSIQLsCU5Ta/2V4hVZkGg+bwWO1PXAN4ak3
OYWyKWvHKnh4FFgXk55aeq7NK+ctBs+qou+AzIJs/txCy1Kz3MMAua0H9MbK5BYA
vJMBA5A6AVVuHCe2Gfm7ql/4XaUVBSsDdeIR2XaTv/ckINsRtmnxHe0GeE+yvCwV
AX1bFgm+Gil/Gz5qE+8CHS4OWekkoe3BZhlvEK48KuZyohLOaiVU6+mo3rsv8SWB
xw0l1suvMyqjfQ2CV9/krcJN7enS8AJNpmLyFOt/yicUorAraFu10JRVfyxlXUB6
bprdeUFHX+W5dKp7xFsDpz6T1J85jYd0dp4DTRmUoLQ9eyKb4BEdpM2D+jnFSuDN
MbSXR9WWlcui+F5K98loU/if3aSnkI6O4J1MNjK3EWOcet/20XgcMZW8c81Dvl1f
HoJyt3+VQMojuac6LwfnublxzZWL4qsvRW0C7acTubFGZ51xwADhHf2xY0012+N/
DPFUwtGkGo/B+h8tl7qpHI7j5AkfZqlzkA69dQu99Io6BaFDLzqFSaQt7A9NSz/z
9agBle6CjNR6vvRnptvNCpdPpmd2cwb73SmRK7SAtBM/czbmB3tqzTY9d5AdcKfn
YW45gV9n5UMBQ0xnGdAJGKuYFae+VS5H+mA6POnLfMY0gDvDFgCb8L3AaAVmN47H
8JIIhwe57vdoGbV8mh+V7Erb1CoEBDD0DpgSZ7C0PlumCknZ4AlzzHnTWb7j2ZGc
ruEg1m9WXPJ8WgtXZ6hrNsmHIBKJ8QMP+N11GIAB20dMLudwzBW/VIvCVDP3lXw0
M1UHmU3FljtwPP2TQ8tJAflyv//uf3o1iZmqVvPTKKWiUIGhQuUuMff+K4Xg7vWX
HcCrL5ml2su4IKjVUmnTuvhmYIPLV2/x7cP/e76CDrHE38gmF8DidH/7UUBH5hN9
kTYy5E1nwetzZyaHXuhCFpUqXBmeBnidyfe6YdqBrox5mFeBqW0jN7wQAnzdi5sK
tGydANvZh4QxA45FAzN6CnBbS0fOCbd13Cawax6ajiKCyu5mCJFpM1LiaeEd1Fc8
Feef8w3iEYxOmDvUAXZbwVT3Gst71LLQKnA08cJrh++XfOpSlCD/L+ax5auiaBuK
rjrKS9VwllrZP6mJa/JD+RCWCcCttbU8nza/exg22e4HYn7bHGN8MFJJDWCGbU7A
o6iIQ1Yew5WsEyvzXpzbqMAUUwqTpcM3Bme5PqwdN6Bw1Cltwz5HkgOxF/sU1Znx
Qw+TJmgyt/pwsAX5MVhE0DuYzsQcI13SWMvFMWskHcsu0reFCGQaF+AytmuN57fO
We4VA1oZpqH/Ob5+PqX2zqg4YUPqvfvSbFCWR1GWLbsinpSBbpN60We1dTcs/MDY
AZo2fvpYUcjscy8iO8RvcE9wMvbMIibBmkL1TPmyvuaIDs49k7LYpNQS56LbHMis
r+TIoMw/I13rute23Y+IXiSb8iNQqh5WHyu/fo89UL8Kuy55PwUf+imMHECcJvcs
IiYIatjDRMpGwT8uiivfHlmeE+ZB21mUZp8ampjdZv1nKohJurexfTtzUBrpG6/M
Mn5iYrCg/VFACrGlAGkWKVAQMbZIq2M6HeopkDzhorsWrJ7jLg2ti4d25NxGnki9
QzEW4qxxu8/epOYuEt+zni3ZgS/GakKjIdrhFGdMyisQz9AYJ/xdQRkOf3/+/qcP
2vnyNKazoYFmVxWrODVY26HYvNK1IbObjNMxM5JCqUtqKi6UpwmkCBnMv9lG2olE
+4zQnQYfk1XeiEGbwLAlvXv7hxjCrF/UdJq2lZN9oy/DEu2iHFQWW71XlCCYGiZJ
VQjvK3x6NsWJf5AQQjtYRv0yTyKxT7Dnq1GEmvz1HWCX6YYz5nCtLzxBPCE7tHLn
Lznr5b6sUQrSdq//2SCoeBP8epANpxP3XEMsd58iaqYr/GKlv7cbEkPZa9xnPMQZ
73aDRYSIz6rpEI/sKVxOcTqbzJMU07epe49lMhcXIWtMqcOSKr7ExPUh4W27XDDe
6S/w3b/JVhRLsNYGFWXUiJ1SEBraRgx5BMbeqyFQc63CJitw5crdnmN6nFcQ5bLV
BqH22b9ze8Yn+XmtBet2dbiMnwmh03yWon0FQ+tcwX0pmMiNXIsJPy5Ug9B/hGnf
pB46LaKV92ZpSNuwgQr3HGSQE6G7fgbBa0etIseEwRQ/DcQaTfsya5U+E1JXUzCK
Ki2MY9Ia/l8/UczllzKqrjieAWWCzgXRLphWLD/RW0afo0oktN2u4xAHPqAds4sR
BkECD4GFp6c8g+4pBmi1lJKbGMFhjcw/uxFXVx/8lAosRBGJBbvn9/IiSNCDhi0d
9gjsYUEzuG2CyWswW7L6hbWc/53nmP3xVfl7uLmHNRhNmcVQHt0xWzsJd3COHBfA
RlTwz2ZNHRPTo1mXOo53pzz5a2laBoKuK1y6x0xOgRHUMvDokrPPaEaDTxebg3b4
KS50EdT55BsOnr7FwBYdJWuzncP9XY4KxNTKKkdHy03jeYd4jJtHqLM9LjW83SgA
dk9ie7Xuq34BrqakB3ovMYSfHkyuhhT+c74KVdlyILq9/b1BTUuR96n74c+eWy5L
p5uXpR1TbO6WDD8p1DmbEuDilZuE5OI8omiKUE7TRjpkd0mtuhrAPGNMPDFpxjgf
0yxZ8+vyC7T15ka4O4s9BU3EwiE+2ijWNQhCtmzjQ2VNbdPwYofHUVLiwWYbghr7
hMgjoE38ZC6zlpo90FOGRWBg4NPmnCTmcDOvMUZ0cZXMx3nYw/Bmgrw0i0sd3ekl
11JTqSKikCTiEo/sQ7wU4j4nZQ2t+Kmo1hjNe4qPBagUYJO3RWJT3/mPMzvFRC7F
gyDwbPn+IlkpeCWF+us05CtyU/4hQ+tRhBVMlwUxKLy5KiDUxoNASLZGl8brDyK2
56gpc0jRBaBz58E6wxgkTlukrnHlb+9dIvVRhJTYma1E13WZh7IbSZtFJ19mELwx
46hn6fEHLTCR9VLUWfbaKGa0G/amdev+KbOd2YEKtiU00OkpU9d4qZ4VNqgbi47D
TCoD8Lws6XD76USDb2tqGWPK1O7hndpzUEFmdIrCma9kfJ5NxKaL+ZGHxZV8SV58
Vz+6DBUxKbL3yNWzHM6+KGqIiEpolLiPSPznDJ6LTdFZW4Htw4VqsvWLY00pMRaf
LiVnZfDb57/XOnf/e8TdCmyKiGuCfmXeZUP50y4pWcGH3nHj+AM2Axl2LUU73da1
VUUqSHHkAyfVcobt/gogQPo+XOv6LE6PtX5C4jXWTIsxGdHkwNI4GozmttxljllQ
IFaOr/6puRyP1loH8HODLMof6BSgi1bYxHZJ/No+xd3FROYIaocdrezv2xc4XZxF
UaO3YAJUrSM/D7LQXV3uXj7XqDCli2qZz0gJkzT5z4A/Mh0hj3qJj/vVU0pX4O6/
+ILl45vb6RRI9KSEFih2sr7umDSlVMY7mbZpeYWqxMwYzSqpsllap8uOKn3lTjQr
ng7dKDenCFOwAtJBTzKygF7TofzwRKjdPtIiUIPFtQmZ6+K2iWqgab019m60jTPq
zIyskjsrqd3OEWEIF7mg+bzmf8tesHiwReRgNEKGvgJI5/G8epcFO/f9sRW9g7xo
sWaojp23GwxAUPXQ9VEf5rdHMm4hrCL1D8iWhaKnhK7AeFGiMuvDKSgW0StdnMmb
GgqcJIRSlnHVB6yXRl5FjARi83bqV+My7LYRfwvZasnTf4drzYWIJmt4Hs5zLvbx
gSomYsD6YKHQSI2Oj4deGwjCzjjnjYNz/inmeY+DeOtcZx0Tgcl+9NMiVbNnwc2d
U3EmZ5Vp2pJ4wm+jgeNCBimzsttC8sr/f3bEA/9x2l5iLV0n6fCCUjiPgY1grh7P
ZxrZysZXoq1JtI0DVNLpceI8JSq9UfCil5ZAO9sRdamlAdaVk14Zxs/GF/IGsrAZ
A3mMiNHCyPlOn9Kg0Qe7/d0iG90rZTaj7TYDB0OpxYA1RGqXpL+Egk3X1BkvYO+M
F9GxDyDnua7x2re5I6RSyB+VytfrBELA3cZdQgGW80kesbCYuM2lxdlaDyR8UZRJ
V2eG0wK8WBvGsjcDGbhzJm758leI5hUyi5EgwMz8JloxTYoclOvJdmajiebcmx+p
QDqQYpaGiogr4XFDsnXj4YHNjQg7xqlzHmsPPsntWrnQa9kkIcuG6b6GoFoAV9qU
V8enWFuIrUvfPu6vdgaTqKH2OzlmCbwH8eLcCe0syqkNiTCKhMehIMWAK+lyeI2z
jWULdunQtaikdChllLlflGuiYurf9s6023bUbQa1xL9x93/x/6TOs5pIEx6caXyn
LSu7fSarrXlrmVt2secH9+WcbWIjVuk49XokpHX+rLO41y4ssHG2dSBh+BI4uaBs
JEjw/pvR4vwcmn6lay89mrG34XFuNbHAmUU0fgb7nbRIix7djOUr6Y75XQPj7RqM
aRD4XzkI7jIL25jxCg0l4LfbHaazXgeFFOJGy0LkAYRmjOGglS5/vGj6dZae1p6x
RVvoApocskoPdo/0L/Htympz2W97pvJYyhbtnmIpu6eTq0xn4RahhCPaiHtB8BwQ
l9oUpuXMevmkXhR93pDoBPbSXc0SzTh7Co1sm5XCrGjQIx2fP0XftfJFQlSNQPpc
kiRhDUBFTbWqtuVisfP477dNLLdVl8Yp7lOuvLs0IH/5YgYHfHNPFc45xRl/sVyW
MkQiCiM6I7AIFBNsGGfINU4QKh0diIQV+gOv1Fe/10lpqY+UxCMy1T9NvH3MraI0
eNSVhT7uRQh88pTynFpaN40O/+ZLOvfAViYxdBU0FH58m7VdbQzuTL/n+Zt2s4kh
Hnx5BV1+RW0W0utXv9HbUn4dMEul+RWItovYb3qNI+1fJb5sj2xnUgU+S+E1Peen
31eVdoWsQPvZ+PKi8OrrvsQIqSGUl2YCYTz2PaaJuhcw0k9msK4egYC02ZTHou/i
ihFqm+PdV3DmaxbCGkNAJWmSt7kayX2UykUOTZEfDKPnwSBE4/7fbWcLZ5ElYIbg
DngEhiiQI3GIDBKgL5fffh+dtXrO8lqO6dyf8KIWG0meEtAtC8Sbf9wVA7/ZDsRh
ht/StoR8Pmi5u7QsJWGl+sBJjknVBXNnWqmR9hn4Jhl1R3aZnjI3oHDCWM5a0Qa5
492jVj9WdLgbgVUoxE1DM79QC+Vvb9E2WuKWcB6eejuKq3FM3Ekt1/pvGG6iroO4
khIoN9O+QH/7OHbQ0Lcs+70UI5r4YCgkH6xj2SyjUgdD3AwFgQhJLGFW7wtXV3CC
pV69W4EQJhtWubd6gNOguk0DF3vDGlwhzUyZKvqJlKb9zgqNuw7x869Eenv2vfc4
H+OUHEI+GTAHL8t9APdLzRR7E1roEz5THN7jc4K2MRi0sNpIuf423IkjAYV26tsF
529Wug9QjB3iErdLYpHbgQiytfVVdR1opTp0SgNR18YbVhkQ5/x8HVHqF7YFo+Fg
MU+KPwZ9gDtuX1i8Cb5V8+1ogP9VYJKKXGNQx8A511tAjs+wzNUkYFEXyJIr5H4G
HZXFpjl6UtO9yOSWagVG2vtvzb6Vrl3eaZcdf9bZY7vSm0vBlfoYdbtLkvk4aWGz
9repryMqgb9Qi2vVFnjsygH3EsowqThpDu4SaiJ78f1zP6AR445QFGXPu4viQuRi
2eql6Ts5WB+tprApHegY3G3Vym515JzOVV830F0K3xNfLqznA9HeE5K/ZCb70OvV
z4U7GlN63uce9cAnl9fdbKcHHxyEB+0ss8s0vo8VmNeqlR7EvQEI7TZXtrAvqo2V
DVXgegZg/Z6ut6ecCsWhCqgKI5Z1v1Tjvb8bFq1NvpXCXdUzAU7IWbnnWLv4p9II
3dIENzQaugBqN2fyh4SUxUL3tvBXCCL9BNPDjj8LcbzHXxQv1dNFwfUnpFSPiE09
9kEHU08JIZSrcVFcONQ0OTR5l6o+xpOXZllwz1hjbbHSpomDF+v08BkEr9uNWTBM
v3+0snQKusHBBhzbRq06SFFTLo6ow8Z9ROsrg4KHGzqKuATrVJliG7co4pw3jnYh
n+6+/2wOkk8/7NDOvld0szY4ofz2G54I4VWHoMrdKkVyRjbVCcCenMb9VxXUVXHP
XtKpxR0ciIWLPOWCGzo+/os7rIli3ug0c/0Pb/9Je+6hu3b5r4eS/u5/Rg/zBQkS
OS3uEHlzZTkXesFesnokPpuyqvVydH1dBa8lnTe1rVMUBk+VB+PT9AtJBbXyBhBn
9IFc0Ptwp6tw4/NKbS+8XK9baN8I9SVWbYJ0W+hjhQ8Ow7p92K6TdeWDiVw72F59
uP8iNj2QpE4g1Xo2OIiBbTk/dK5P6MKEnmmEFKP/HLLxCgczHYbT6Atb5i2l8i3l
V3aiNTM8Nut5YYLVmAdl2bc+iDZ+KOrtJsXLrsba57Jf1+6rPhVG+IbkhePRDr1c
kYRKe1y0RNQGWwYgkn9dFjRyquw/2zUWgMxoFwQL+90ZDYNFG5Uy/Kg4NBitAFlm
UoZxaHZehImwFev+KBuJOExcgZv6njPbYhpwHonRxYKRVNXn4FJVeQIB7SDn49yj
HTeq5j5zlyG9h2v4wup05ydGx2OehMOzTZ3C2ZycOncv4BNi4UZqGdvZbmYtbqxg
nVBYR16Uzjf9HiiRFjvucyoqYdDGMUH9jbjR6bwQbclA3DKe2nVCuUo0mY3OAeqB
CuOoZLzQUhZQJcNhh9a+88in4CF5q2Cm/roYj3RYIQrnIa2y2hEbxy3lMYNSnC5x
oOtcJC/Xw9R8vbUo0G2zMyK6OmusCwih3vx/TpyP0Vr+gdELCzNb//J3A0JH4nsh
mWeFq7mQWcL5+OnrjwiAGuj7FdCSAi9AyTLlyWa1ZjxLdDAdlqMzn+ll50Giqj+A
TBffSRSDG4P41DYi8fsVOSpB1c2vvjJlQfN57qlgAbrLCo3Yxqh0NEUkMt5N2VXw
g6LrveOzaGYOcpDb3yf/zHp/us8gC0KhA4RaiXT62/xLEM/lb7s4Koxyv6sOrraY
X6W0TblIVyNcUwNTbUUgZhJHymCoVOUGMEZMNmaPL1YXexI+/CEolqnhIvEjXoSy
CoyoBvh6PsjcdbdIQdYxDgtqe8AWOsOXJz8uhS4i/cznUHeawrHP8T1JRp9BiPAD
/Hbf+I3mLAzZ526M16eepf/djbYlIGkTCxu4931u1plR7r7WU1tQUt0gNBNiju+F
DA60PnOI5nM4EEK/KFP2FwXqL2Zvgx6pE40Utmc5Yaai1S1iyQgE6C0tFHcMsgNP
03pcCZ3vWKGmwMusldEweRLYGeft9xJu94MqBUamTVF7kqcPW9lBeffvEQa9s5tM
y0gziBT5Uxmu+btydU9U24Bitw5BESotRBUQUvWgZ1UNTsl5oIg/mlPS+YmM/+Ju
CGmNbmjC5j5v2ZALjout0Moe5KvCMgJPF/ECK6KU9FNbwmwLQRN89s+zSMoZjax5
fgvE3fWy8bdIsRPepMS7Um1Zc/q58HzGZkyogBj+EhbO2I/3UH78qTwlStL/7qVr
C7misf8x/Htr6m5nt8VOU/Egp3ULbjcREGvwrH3BsazsWdcXf9f/hrgfVqdbwXXg
V00pG8TKLYH8MDo1fRG2BXk3jZ+eRfiBx8Oibec6eDz93NiLFiS05igUxjzEmtza
WfdwjC4PhgkpVZGeLTR30Xrw+HuFKvMDJpJmJHDHVT2uaW0QALcETDD+JgXyec28
6RU3GuxF26a1wkKB4HZqP9BPfST8ZfAhdLD6Tq9mDc6z/ZaFezlxpn8IV5Z28UBI
PXpK+LMV8V5QiSJexMgUK8g99Rgm3fFphy7ljhdbxFOhzQ3TNptc5laaF8f/ooCB
//4+retnlFo4evCbTy4rIrTqrxFCn+DA+6O0NmCIYZ2dQGo5aHwZUspBOfDrkadE
kYkYqHhWPS/jp9x07VVmYG1oKcugGtOe4aHymQW7bcxN4p0lXkkVwSkiu6bLAqmL
CIi6ZEc5vRzG6akZAg8lFXbaPmC8tz2NhTqu3Sr0oWG3BXufyHu0wpflnTH3I3Dp
Zue2B9jC1KW6fFSo4lX4LmjPGg8EHtLyBpBIyGdDGopmx8kJYiIRe4FZHaMm94jW
Xv++gDlxJ4gXeLknpx0wCMBB5Ie4KW8f3zheEwlLaL6Xx+LnLyArG/lkk5X3FzLe
fozh9xhvhnKlrvEnqQEAgu35qUnYtDglDmpbWfeLCrn6V+4x9GOXyN8asQ5vZlpn
H3jc9whJ7b9cezARcdrrmmRWGDG60hCJ473rr9YCYnNWjEA3TPKHOaAom0oyAYZm
1TonlNMbETNMbOMwkhGinRZ6ERsTfQSuJq3KM18kXRB53VSkaeixosfjSu+AOai9
4S8EMUWyzNuxuq6KzdvuFXdGrMXW4hZhIi75bt3DQw58AsOPBvejVoLMSPrctzpg
o4NtEhjMTFtV/NPDHEGzQtf3LAi0jVyLqMIq8+WbKcde88AP25kn+vlutGU8X5Dv
TGQ+rgpWbNJ+qyGLl1URITZcoerg95a2+gmUsueuK6W/QHruKSHBo/Pht0jyU1oT
DaSEVS0fGH9W8yTJz8AWdvCPmEpm5AHcNp0NCE86B8ujS1/JnhiAJ0vJ1n1ycdEr
JJnEyrygHdIiOnP8YAyGWpr0+9tnghCJ0EKp8LKMlVl7ZxgJSaYjPYGw2QNK/agN
uF/vmroreEqYaSK+/nIVCFf8GIe0YQt5NFnnomDV7n13XgUgX3VvoLt+D+9n/hY5
KURKxUhlJZDXv9ToDnT2rBziZ4Kdp9mlrCa67cUO4tVKbued7f8ObVWkkhGYHV7N
Phv0VhsEBphpupZ7ZPNzs3Fh1+kTnQEqYTh2fJCOwT9EsUFpOoBbgiJAdgLcY5Fo
+YH2ncOHXTPENBaOleXG2uvsWidUYk8QZ9yPoUR5PbsWDUHRV+KYCyUYd+NF73OP
aF/R2lAa5tkdN4LN27LB1q15dQsirThCSyYGBxwobQBvcjOKJwM1XKbIBYnTLZwk
itjjA88cgPG5Q6TccDz8l7byqjhN2AY9nDf5raI8CfrRKiB2wT4QttAgtbZrHdR9
63NFbEsZHDQam98wWQ/52ejCIvMR/SI3C4seUJEQ5EA=
`protect END_PROTECTED
