`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+INARJgfUzhYfqFrNMzku6ov19hBzS+Entpi0Ar00hS0KCHvNGO2KdlonD7Ueq70
mc3tRU4gglKFL7NjjSKKayA0sUowAKfvF25Pc3wxLoxwyk19PwynwZo/rJURaV2s
O7leU63dVgQPKIsJxFxbCKWOMqERimP19RSvgHqmDvs6RW7FqO4oXAm4g+Rm58It
MTB15lgEGM1vfd+JEx4dR+5cyNJ1qaD60R7CdQGWtAikysWfs63DUvkHH1pr/oQH
eJI3coXiChcikuS8jau5q/4OBy+SZoz45Qu2NwfbIOqJHURmI64ffWPTJkchweSZ
TsL0TlAQJUjb4A2cu6JRwj02gjnRZ8NqZ7Q2dYSnX/cHzGgcy8iNeFIOZm7713Yg
3+d0m4hVi72A077BplVviW5PW8jSh9cRAE89ASSMp473zWOFfkjgzwcesALTAKa/
urw990xBA9wvoVtDj3L5/sIF1TD6mNPfBg1sLBLU+lTMTLeQd3q6lYR5hyR1Y17t
YRXh1UsOPXt8a7OXnlVzM6tAlf5fmS4JTZIPhuaUuYJsEGJ4QXdS3vaX2BK7EipK
gWvp0Dxw9lMnnZJxJ8IoizEsXKqU302IIpD7yOEkLWCZECGdGn3nqlfHOVfEZinU
15FZRuCmnjyo8gUVk7Wv/SeGQt79SzPy9hGRyzT+0z+8b4of84mXqpSdv6UCU1Vx
jK5f2SIrmE1uK3aVr7IepxBDxC5PW1kxD0TFMFDGHr2BV7QhFhA80SZlYTBAI/20
`protect END_PROTECTED
