`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1q5dSKa2VVf5coTrK6zjMjCkrG6QvvfdGDzMn2n41x0fvkBZOFAyEwMslrDIssnQ
fB/Djwuet13hZSF1MgJCu+3Re3Jov0vXEqkdix9UO8HLaif9JxOMhZ55p93Uwz3T
A4c7PVDJ6KTUN0hsGdsxpUbWNtmqlM6ONEecxBLn7ZsuxsuJxSnj1S+ItX628kkT
VLDqMGge9FvQRLZ5kxEMc0BpatlDNVkQPz+VPZuwo/u+x3N3M3WP0tZlTWH99ugf
5CqL2xgEkBsJZkP13qdEBP8YDniWgaz5Sl2rvDlp0R3yqO78mX8fYLjadBOiUB70
fXL08T62vPrYaVIIw8h+r/GMDsCXaiUvKimEcU+CPYOOhocpddmWhjDgrJiCuS8n
XODe/jhmi7fdw3rTtH8kPOlyr0exzH2PzmjPqk8WnwUoj2SnJiOa+SeG9sKFBto/
ZdNdxEaV8KS/jHeV4VriDEMwICIA6dtLB2aDzHTHhZ0DYLF5nKghPlPXipVh/If+
QgiFvbDhZaigjuS88FPnsEWFVcP0UlR2nCyiXNIRNzfNjWWXX52yeRaooS5LRoAl
DWctAQq4yzOA1uwXEEGDzwajBkVq+s9R7zmznO45P1b2YHNNTWncCwW8QkN4VEKm
N8Nh+jyeY9BQfMb2YRpC1ERC+ju3TuRUk1TdXYQR9Z/6K5NdQAD/PLL8Ib941yUQ
gZ37qD+gdtbgpcudjxyYHdxSx6qfUs12pjx4zf8f9U8S9f9YQ6jfFzLJ/E94ZwTf
KGtVaPSGpEnJIaeEqkpRPcS4zMV9/JEOMw0H3ks8jXO+Cj2GRU2lrD8bhmkVW2k8
GXjOY0eF630uWToRD1ZJSVVCc2MHSgX071T2T6JcgE5IibdyG/VGrbguaNQP/vj6
nvILMPdWjrIhPLc6C7uvqWVgBFzcPIJnPva4AoS8l8SfYbMr1L0PduKMd29pV0HX
/xjKya3ORooRmyrZinwk1QqJpCI3wMJ4PZ1CBXtnRnXK9oc2we0EwIrn1rVsX2xP
LLRk1NaW3iT+wGa18hBpKMS+8mumUidj6g2quiEqFAqbh6/+Bdr4uk2YZdXOZymM
fQA/r0KB0IWDQqndKmOagl0nHLUkc8iD4RaOhOrLVVmfPtDwtVrjE00gDFvQQbUc
KdlZKib57Pfk5tFMDIRN/zArxSE2WD2VW5MIWcMWxE/5c8tG2uuHzA5G3F79AO/f
pC14L1284J8e+q7PmCQHtavdW4/tUiLRs0kEUYeO0C7kpVLW1aQRSEeJ1KVuGeO6
RVgOHJtWbERxnHsyTVWy01DZ75W/BVEXWKf4us20MdjeiFjloWsX1PcLBorwKwb7
A+N5fJXY1HtPcqiplI2c2WokCL0+QMcKtJdnA04AQXO6VnhxeU7b2MHZ9/YKmyPG
FUaoTHK5tdwdBJXJnBFI5Cx7Q1MwVLkYfPQlcVddSir7w0GQNicWfhlfz51zCRTc
J2b0QOUeK025FG4MLsX/ETNKi0s474/aiPt1AWTk/OtTmLlOrQMtL+431qw4f13A
bGXbcmgIMaDcq1pcXvhTw+8sRExtgd4t1P1DTQf2qqN9GZyLKyG0B4YWzrg6huTi
v+4AEaxIZE4MJq2Yut/bhCAcc9kL7Y8dcTwxq+nuqSQsUa6bEC+Fz8UkfBR/jsvQ
P04mVe4MV0TkpfB/lqxrkTzLsJ0IFM9gWnnfxKsUy8W6z1GhtElyDSYTstHmzfIH
FARMhwPRK/rr5bBEcP7PGNRYPfECS8TIR/GpxKwQ1t+5ZGfoPX4yKJkfWCqNE30m
J8XrLxPF9cHrwXA5hL0Lcu15IcfAMfIDMA72eFD1QH3AppLga+mNQXiuLCkGTfi6
/hCnUxYcieaXoJ+pqwxWMHnpIeTH1BhyNQTjPXmMCIREcYr+u0AhxEIAXaYyTBLN
V09orZWkLHqpoSipW9dLoY2uTCdPV+QVnHTBgdOaE9TbfJNub+cfR6XdJiCE9K4R
SsYEqFY7grAMk3BFOjB4wDRtVqjM/jxXgZdUNhKJVc5FOsNngQyVEIwLnuYPnRpB
CaAAddUsqoLeB0B1LKde04wi3UqrBp1SmBRYyV3U1vC3xfKCJ6x+Ba7XAn6Cl3o/
stfdDIF8AV6yJzMkbBblYFYhtoKXahZ7i0ndNdq1k+l+T5CwEG82GYNdjh4jv+mQ
p4EmmMom5jzwMeKr4XUoXxaNiEl5hTPOlc0+mK7ruKVh3lS5cPnzirAQNHFBsG8G
bsDAjTROaQb4GxJGbMqY0NdHBBP/VosIFNU0No2//o2L15H7bIcJVONuE3XUelA3
6erJkrP8fC+RiUYI+45nIp4TwU3ytZ74D4ZBvgAIJ0Ot+yoj5KgTJYTfKzCd6hOL
f5GictHsdV/7qaCxD8sJBikK25gL2zFVQgy+bF9FaUUxB8QK5BYW89FlQxbBvuyy
kZJXvnZATVRMgmpV1yGrV/DFRMtckdomYCaPcJJUXep9OMRiKDWlEwWGamUXD9E0
bY/gSwdRwtJIz/de0mdHro45LrDVVLwaErFYYuKJYYRgte+DgbYipNNVUti4RscE
M5hWp6SLp4+qEfeqfdeVcDPdy0taEjCftE8LiJhOIVM4PJFyRWRrs+E0NBGDnMxl
XBMA5iJHvVeH8xB+MvzOmHP1zEXxDVK9FZQLdjQqVAtPZ9CwRi6q26zJ144PhBWE
vO3qWlf4Z+Y4jlneYfTkUA==
`protect END_PROTECTED
