`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBXymptHNzqppx8279hixljZnqfGJ1r0soxp6zygUd7Oumz1wU6lqBXSmlq6Y9ed
UpPZbUaeZ40+Tbphnhgcl6+5VHcL9PMDUTW+iOz4XKR5FmxpExh5vsFSiHIqeMuz
KykEQPWKx+xCBIb4yZ7E0i6ausc7DpjTVUZm8/+VtjCVxvSGGZXGU5EbMIOo3GLQ
mJRNc1Ge8P7rGdthgZdVNjYKdFLPScEov9US1Uini/yMJ87TzlFrq9HxxcDJKD8L
eLurZfqdd9VgxF8fEoiXuGur5hKHTmonqJUqd6K/aoEzLOoHK5lwvmW7BGgIhZQP
OtioTVdtCznfjUG+8S1/FIZrt7Jr+M0KS/N5AuDpvojgUco29iKJcIyELH4leVdH
OvgYBw29TlBXuv/Lj5vJFwmBN6gXTEZQ8T60iPyl8+7xqFydvuuN9JIfo8a/3a8S
cmlOSOCu0JjK7GC93CbC3hmJaj+MrHpzvQqCd/rEzD7TN2/I6jHkp6xqGM2FL05z
8pZsdJz9MfmlGNqaH/jrG5y2YqWtNmlVFWWdi/syMSyxKj6Q+FLlGa7+0JPBdbO9
H7PIdMZManlSdgHmShLBpk4IIVd+b5gjg4TqToSFqP4J9JmXmWoSF5Lln+3RKV+e
Lu1MZaVNoIusWi+tvnrVJHRo8r1arOzqvnz42tcOhofXxdEJ9MfLKgLy84RfZDTI
tCCqeQRvv3A8AMA4pN3GDETfwUxypU73m2bXMyIxQkvlnNOzjjpQjXxaOpjMMsTX
mnRnz8nOP/W28G+ik8SqOmZTfQXcLQOsuSwFr8l5mwBbic+lckDNUE0Lp4cmP2fI
94XKixPRDt8xIcKY47apHeVWoj1LVBljIn5SVFUrNiqucyxyjCDK/qfVnkrBIRNG
u4/gNoZYBAB+hplHB+NvNsGV2FTd3UOTLZHnZYkGRYQORfUmI1voLvPqrYPqntYO
L1VRAmKwlAjPXoGHvjQr/poXG+3paui2e5Q50kDFFrsj3TDBNFzMqq2c4TVqF4Tj
CfHDdxrr1UQ0fPWHFS4V6dE9wljHjQXZzHVn8D/i/5Nft8wVLOiq7ndECzBvBFzR
uVsbzzcN0LD5swQDyW6iiQ==
`protect END_PROTECTED
