`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ky8Hvfg18H252AFCRl2WYOz6jZStYJ9jjSfaYUjIPguEhJHvQDqlxTc9WkPttiY
R9REH57OoYPC9OPtxHjaS13pgoqewd7kjN01RcViIWge5pNJdDymgvIhpbTyLG4R
A2R7lQlmfoEugZDWC4epEWqkAeuhVmczTwSJ4r4SK61TfK462fSilSY0qv9pxwup
NgxJdbx/9zLFfDDIBevLXx1laQDZPTJh0Hkst5mRXv6LvH/+h5xYMhz+gb+FXLVJ
Nocy9NVrhDNarGYQ4APydu9GT/JZOG8bvnQDcOBvfqAEIevx/b8BqdXzcpbnDfbB
veRtTh9di9d+wKs6O9pOQPcuJAgX/Tg6FPnYBhhPHmy3dbPFMEGowrmy+XWvL5BS
mScpL4ktFkk7OhQNIpXulvFCOXd+Y8BwRr4BvBeu7SFTyMXjcKXMghhMayfG0MxR
BEQb+osJ4yU6sejJbiyi7qX0i0cnAfMztGp9IdCKh5LBm6l4SSYXWNDurn6YO29Y
phxW+rOtJ15H6CC9a+AuufOm7UGrSlpwU3ph/wSCDEuxDTZcvr9i6B9fNlkX6X+t
Y969K/Ax3cpwCpWIyKN0oQU36VyVLXGGED/o1q5ofcK8be/BzX2Y6u0Xnlhr6T0Q
5tBcVFFztk3T3rHNWcJwe6hwR4znr0bzmudqd9Wnb/8UZeYqtVCBgUlxI3BEQ9qe
kW1YiNHa3tsYbq5gKcY7lpWc2VtPbuYi77DpW7jwOGtd7d5vyqa3nRN3DbEqoVVA
fsB6OBJKb6ByHJgezhVZlAR/cqcsWNJxyUNO4jQCG51hoI+QwWz1gsWzEP/G5cgA
lnfI23qZNpVAwqACQ1YRXiHlrGpzAAa7DhKTvThYVI7q68v/g/gq0NimHB+P8j5p
BMoZqIKs0+7vinuYSt9qpC4p+TGkzrJJRPQTFwB6Hx9hNUrTitGu9tI6HqsmsO1F
35oEra20Wj+DQe03uNOmpHotLqARYQEBMWr9WdaZ0z2ZvNvSOl7pejLhzz1+Z98b
G+aH9V9XU4F6y+/KAbPmRg/7uno1l0FyZqZQmBGawWiHIs3+cnjG4WMG8PUzqmFu
M1Kkckyu7aPpQ8q4kHvgOq8KZ/epLClSnXXpSAekaz6GwdbKZFOY+0A/+XICPQAp
hGuNw0Cscu2sOADHMlO7Hcf2nKwsvkXRJQoVR+1HPhG5WJdHR1J9PsCUwJnUJQ5Y
sOwsN0B73WNdVlB61D5XOgjIZX4ySkglmOwNafEZ5Fwz14nxOYwUo8Ae8Xym6yzu
9y+3/kaFbd9XyA3Ps8DVPykIE4LLxRG87EF/EJ1ueXCSqI4+PaSiNSCf6TDXJ0Xt
nnOmVE9hlh/JZcjwYKm0g+eO8owYKmCGqdyEVl8zMJElrLooMMg7PV2rQ8OTzopB
7PwpGJ+y9wW57qOrRdPdJE3IOLKT8Ow0sCnwxo1XtuW/IWsKlMa7eK7WPbH1HF+c
GqnqWqjCz7BwJqd/UvmozVlRjlNvunTYrkVueeFOvQjRA21PQXyIukwpAFL+ed+x
h7IN9Dz2QnazEcDzavQHKK8nnmMJgbcR6aABUBPd+DaqwIdbbosw7jJUqHvmolBY
KzeTnGqpVhaC33EurL9KXY9kiuhk2DzPx7GAoYzPyDvuTKYk5ZtWDqCK9Kkey7Sx
DHvOVeU1JUwQ1PiiZ7RoiXqMbAJV43fQuYV5Nfg13lYyRIMIqeeBmZOUjt+UExhl
Zmp5BXx3RCpZ38Si/waoXvofcFLzFy79LM+1ieUJ8TWVHycsviIMV9CxARZORhKo
8BE9VCAU9OaG93I+7ULgiSfnYVKvScFDmFQ6lqsjROR2Tzxe3iziRkaRjsY36VT8
Oq1q91iL/DCi7WBj6+uC+LGBQozQtuSRHNs+mUIDN4FixYbdRSMsYDJZu47J+JRm
EDkGp+xOF1ndhNdLo0pcvQcjLQ+V7njKhIEpFMEKkFmXLGdgaUg9fIRCC8vyLMt2
ZvX/wEqtixngfwlxPG6wtBbxGiMKbNR9cG6LwQOjB8cdRhgDkleXgybVayABjtRG
SkWXTQqNJcTinXuZgI85ww1XTMmCCOck05KH4lwiweGKSlS1sG1kLbeMhsTTLyIS
+qQljK2A6W1uc6TsSGJUkdulRW7PvkdUBGqkPVj+oEqjCn8l/qqd2aLQndt5H2BG
9mVf4gIOwK3OitWYs7z3EWWpFzbiTi9mRdEzEZQsQYeWnvn0GT6zvi9YD5jGuvKZ
`protect END_PROTECTED
