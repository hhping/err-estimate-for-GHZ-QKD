`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Ts2NM0aKDWvMSOsSN0cTONEMKfo2dDo6tyglCZ9sY5/umYWXSYKWSCiD8zr3vjO
usvfcpPu4mQxfdeIvMQdx0QkMzsF51jCFnOt5rp/DgcIurY4vE7eWMeM9VshvcGP
0AeB2krOxO5iEbXvYcznT3CMtzGD5p5h2y3e/YMlVkP8xyb9oal6k66IxhxRe0lB
vN9ymXyPfqsOIFhpya0MPk+1BI27CwZzCzZRWSkLp3XY6pncVWB+idakQMK0Ob8Z
+ZjVYlETTWR3JG2E+bCo5kP8Jmozj9YVmo4sD/X1XK704XcHwFbhSAqDwRJ05FP4
orClOOWpmHXERSqQfHjj6rxGRSa5e4tL0+TxuiKeJ9clTlm0GsXXLIADLPTSG0tF
10BY+NNG3glbvHk56JxN9DVx5HopCA1WXL22xJZt+ctJBRiUXLM1jKxMUM3MUnGg
0F8jlxmTyXxvIcPd4EAXdgattiIy8bq4KVDMC7BRAFmCA4ol86HSSIQzChXxlNii
FWXTXJy+Oot9Qtab9GpS9HnKCtrmybP5R34/0gMcS1pVGLISx0+Xoop8uOwLd5e6
wNVq/eVR93jVgtFGZjAySNCBVJBe1r1Z62OSahHhcOu8tPiNCi/7xC/74othxvJ0
RN3VTGYCvVNPC7EkHRx7sTTe7rylK8qZhzeFW2eMzUpq0oWlc7Sg1qV2r0U5Pg3M
5iWodffRDq+AF8j0LXaJRSzVqUBdy08exqmY5BRkFaN9225WyFF8+3HmBGTpGY++
YqI718OPkpsQkP18Evkr4ZeaaO+VBPmeWQmRznyPCPesnZM38LTjq5rYCps13MNH
6DNiAjLz2A8TvOE3MK6vc5KHM1rmvTiw2au8Jr+M7xfpXBYMp7PLSXY0wf1TnKtu
v8uz5259E6xFi1J02b6grh0z7WVm/wxs794vKKK+G/JEmWc+/LacQhkIWCh5XxXW
U39IdKQeGT7c1JlVsNX5iVgqfCybZbCEkyiystvby0c=
`protect END_PROTECTED
