`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYiLrECd2QlJMmnaDqQNyeqylOtNmgiLxhqT64ytnbOfHphr6Dqv2K8a2BP7ZbqT
iCYZFYInv/6cyLvNZI7oDOpscjocVZCW7zs/HoMLDjUaGabmySkbnYPuzopyPq4r
MV6yYtoPn4hGifAfFv4xWt1GGwOIhIRWYfSMQ0LfS/clNbqyrCfOSuVg7b0G8vyW
KTz1687K25kJAKu4xFUINOjf6B+qxxZMk6d2dxv2qdhu0h1znQ0tMydEGEQnl6GA
qNu6HCGItozt5EpQAKvgCAvdosJrsByYdpSdgW9NCO1NoX7d50a8jJskhVZnMEpI
A8jniLT2IWFBUtRoTBdga11DdQHlBpIzzuT0nNH/onyJ95ReKZ9fc+Ot7aBgZ0lD
PpJTRGtJnFmNEFGXwwH0z7/lxFSpLqdsCOPovEa7+GtRVgEX21ZTolEUIfC6G5Xa
63rLbTrLBdX/pHLsYXGK0dIJPDSNYDqt5Yn/oLVs6KidIQpzH8CtyHVfWcZzabps
cz1K9JbPZsd96tUjwb4r034dQk+qSfa71MMxBNPSqkNXMcfcDEbt4kCuHGZfy0jr
Vsfvd2KcTpCjZDzKHR7zhciCQRD+MM5h1fFZjOP+l31HpP/DFRONoFJI9d9F2oI/
yrvxtRqngQOxUEb8j8NZ07VLVsXdmIue6ptoXFznN7k0aJaz0W9MgeTFOZW6TC7g
1bfa5k3RJSU4Tm+q2QUhtAUmgpJyODW7WHRwLmiT68NvVh2VXFlUeYV+jxf/2MXK
eSHypD3gmeYKNTSufY0s9ijYvEeh+9FDDo/aqvBLw8X/j4S6d7+UiiIjLYkvmlPi
6Zvp6Sabm4s3d9RppIw+1RG2kb+OGK3UJUBc95D7EpEdKqrMhlHqFy9WB3B/OFbI
uPxidME7qHQkQC+AsjmKnYLDr81R5WmrUGo9TKQ40K0bx1Qlg6Oxmeh8sFfrqxmX
yD4XYgqo3YjlRfOexYA+cetMPvOWWArpDr0MB7e8qc4JLugXZP/njuHR2FYVh+77
bX69J1m3wP0f/k70nnV/IMo4cEG4OPiS1cGmXX3xRi07OxTsmjmg/G9f9D7XLY/w
zFWqsbJ9aMj/cRbdB32vKShf7lAH/PQwuOWcVPQ0R+rx3jzG9rz6XPw1wACPj4rR
qOOr/qY+BXixp3jqZtF/6zLoOgz1tgn4OIIFjcTiMtaeNK5Sryf4TpLX5wslEvt+
dOBIxCDIXtFeGyrPHDZRvzL8UK7Sg/chPjf6AgxPrBJ9pZ/NTTf9AXL7Uc574C6J
p+vWBVAJLpNq2WY6Fw9dbgwiWAMaMkqq8URnwDsn+1gIki3PI5ew3TIe2jncde8F
OpGKMy/oJSvJLL+ttPB49nARe330/iY+4L+7mETYz2/gZQPOexR9sDLB4svnQ7Jm
626fY9l5KTkV9a9RTf4hfp+Us1yyBGGRX/0QhmOcGMMjzXW5ToGfhPIfCcLm3T6g
LpcZt0Vhj7noSqLuYYalGhAgoo6qIz/HrP3PCS7R2Y8E0CE5f5K1og9CTwxluQK9
1qpYrWZCKjtdb9dR8Sd/9jUT1zo1aa6K4XH/z07ZuEo4rLKUIzPv/PzXUChV/ZTc
X0tao9t7iqFfiY1RuEeLyUdYm0yF5koaXEkTxkz6srgcXZelyfH7m/RY2YLvCQ3C
CcvBgx2xyj6PLFqLIK3UTsMGyiIbtnEKRaj4cjq0e1SC4wwSIKLJDwQt4AM2Zr7P
DG8S3B6fyB/3rmCRrxxXcOh6GMaCsDldZel03X+haq9MF1Vf3wHjRIXUoN9EMHn8
pF/adydi1kiJ+kUJ1mSpYIS+4RNtW0tBnsIJnm25BUeZBIZwDh5MYPMkq43OJRSx
LoqHMqfoZVcIXAVqxRG6qzeDzQx0aQmOjd51NwrD+5AzUUgPxT7oeUyfwN6q0Yy5
CL+u9acCkaQcRbvVy5nhKXO76NnM2SlXiJOPxtDYt0CNR8uZ1/L8jg+8Kf/4VwfU
Neo2bU7074i8rq16X7kCM3QA1Sf3ChXddncgkEbMKw6+kh1yNh0VQzLXyW4xRrF4
/JoO4uUcd5+ufVCy6yREhuZiIobEu6fBeB684eaSCzqVGRqmCIReiPjI3YI8fl+i
L4pPCT6ZCyBVRvdOQxMoZSrB5wtT12Yy1MoD9f5k9IExhHFCLgD8b/bgaFsgMP/B
OPLwiiTU5JDPV7OB4/kuvzabsy9Ca9foOv16/tbtyG0htWMotR4jjpv7h4cMlbCZ
GiHAdQbl+xmz8IL5Z2+bl970w+esfSDYiLZr3xxG5BbiSMk57+L3eYGwW6GNvblw
cyCXl3yhrYmDrS8sU+8hjQWKPRmaBptPiwMs6nKHr9a0O6j12AScbfgUXlDg1OIo
zb/v8CIQd9/WRym9VEwhZKtokhVSSNWgG1tzxC2Elk2FL6gPI1rvoxM8ek4+Vf2S
J6qqwjZaMvaV722rbtS9BnxLQwkJY2F9GAS1c+VcwvSHIKveeeWqGTULjZS8UoW0
VdrBZzPf4naM9Yz4jqV4BM6AQsqFpkG9Y315lcHPKb6yNgtU41wBqG3cAagxmXZ3
M+NAztwgr17KfSOsfZw6qucycVxms8XOTMZ5W6+H9DJA3qJlcOxZl1cCBWM5v9On
+HWjA+upssgowGFKDv1Pa/PoasVW/+5r+rAl/4Jo6kqCjXpLAEnAA37d17WmfFYt
bD1XT5eJrsdJccfiFZx/iZuY9tqK4EiQUWIXV39gMiEs+MmmzU5KRN0fnM3hWJiN
ThcBcGosMFMK9nTVr9xEWu+Nb24Mw2sEs6nN1NUQvybDG+hg2jLkyYPWP86wsBaS
3ZTATHZnSmLX+QgxEWuC7eyXGPlAvNVwLeL8ab+cjq1Lg7da9yqg0/h3AWTfs/Q9
mTvDzmhhh3s/knGgMVPd9IcuyXmSBAi2g9cHRmVwnkPfzln7awBvB8EqQZiF3SPg
lWGYY8h2qbWMwpNPOzhaZS4Ka+sU9uK3EG1sCIctXY8g6YCGAeJk1AJhW1T7jjqj
0ZcE6L9vi156ed01R+AjByKbWxk9OcZako+VLdt+3vI4/RsUd9mnB74l0kNOZQo7
yOV3cSzTThfmNh4t+EjGjfS9ijrH0lea8a1sPlBB/VkX3mQpW1luL4vtg85ZDZVx
eBJwTjqvLbWDM9z7NzNLYUFdW8clQYKWv3VvcVjtg3WP95/c7eTRZOIhArLj8uFi
2WOKmYXpWGAFmREmORDSN+J5d18GML4V0/ijg3I87lfeJ4a+1NFkesE9urNkawn8
50JzPULXym9Ontzt6u1r+BV/d1M6w3+4rKWuPQVaTvBDxyQ8CtNRRMnScfgKnVn9
JZAbor4RMJLQ6Bw9Bn4AeszmUnMSd+OmyGfb8yRYYyiS6KrqayRHnaN27xwiC8rs
C8PkjnPdFeWFG3v//dlnUw==
`protect END_PROTECTED
