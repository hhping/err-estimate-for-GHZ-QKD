`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEBx/8ScHhR4xGd44ICWSZW8fR4gzl7rUgv6TlHBzgsfytW+xV4VB/YxtgTcJrPu
NB0J8kTJwFBYcYDS4CIwwyyeMFWC7uQcSn4Lm4qi7DAaj8XK0YMVaxEIr9ftUjJO
ST02c6cAWBPIdJ3Hb4NpHI3K6jwUwCrQmMufV4sTyJTZnZY6biYtixCcOxptTu90
fdg+nvI/z4K7mpSblfewl/S9OUiooJ6XMateDEi7BO6hn5zk7m75UmAF33a8IdtS
ZXo9BMfScbtWT4EucwrBykJAGcxxuRCR1IhvkW8GRo7n2//bg18/icpInAD+61AN
u+G+IulVwqKJe5MxqcIyMDxqlE/621AOjy+yVu0OLlNbRM/ual73oRkp2YPJ32Ps
eoAg12Vw9kluruBejY6pQMv/+q37fy52UMbVJMXZY840scpmUzunBDAoapYJ2Bqa
tZcUSwnVIWlCf4RmTiKblylm4JEPWtM1I4rQ6V2dC6JLeRO9BJLV5BE2EO1Obine
avOSLDdJBXQTrd3bxXP3nTBqlgs0aEeHScDiJsweHtE5kFyidiL1eACV8j59hyZb
Wy03Y+oUPooNyL7Hhu5gi/G9p6ecitqd8cnAFva9eag/udXSR/PNpDCw1s2bAyV1
2xdNlV7BW8XO57q6GAgkbCKvaipcBiS1Z4PfruSMNc0KXjgNznBVidgZ+sNH94VY
/mt3S/F3oJyZG33bsbMY0ULGrYw0dpmKDaHeVOSrPuDdI4Z9dlYqbSexKZMiSjqD
EqNWXZ0ZnyiIW2Xb5VAvlPdTC/daMujkdnl1ULusJ5ZKDM6eplbsEAqeRWTjgMUN
Gi33vRSSBIKtWmu3pUgHn2Pndz4H5rk2o3BVnsfsJ2H+kN9qhdplBQ4iddDsE0vZ
4moovUqP5HvfgTnnydTH2rahLK/hEIn/E6EYx3QgCkcV9v/d5wD3uvTG5JWRxx3S
Xo+p+kZmvIt7L+Qn7Umw0HJnIujfERguhBLrU8kl2a47fSTYrMvgX1MOd7jkoMRm
7qRFVvw4FRjVnyPv5gHCmATteIm/PTj6jtoADq7yM1LzqTtFgdu8fUvbrbwpJEu+
eOp8w4F4cQ9RBkVdIvuZZKtYZ4s96xuUAg6XO0rtpI8zfyop52ppwPfIK4gFhtb8
bUhhEYMOHTNdIg//7tuP03ClnZDZk1veP0XgNEWGgm9TBs7WvFXaYCcsZmXeGS68
J+rWzTZSdGvYujKpI7kjNpq58z+m2GrAaNWyNCo7AgUmj2RmHrSDeO6Zk3727+PS
Juud/SNblyRzXX6P0qrsLhoMfBtMIIOzHkj1lkSx+Y5CWqTzms2sablGogug1jn4
f0pH2lu2psbtf0Xi1jWUPLv0Xj3P+maJ3emK0OCkK+CCl1rZLWBSjC63xOEFbUxn
rZjxHO/92n/ze9nzX/uF2emgfJSitFrwWce2BU7LiZ7vlAlKt6WJwGFG7QAqMY3p
hdU6l3UurHNpw9zczZGgwLCUDI2eSgGq4qcTn15PfON+8/Iv+CcafLFwxxXZJAM/
dY6B6DmsaNRgPJN7z+XlZo9gcwyJqyH804ob+V0KKUVpietU84+huIYUOmuJpOcx
pNtdWAXDPb4AmwfENex/TPFMY6X5GSbY1ieXORuOgS426DJwIUdoGltDUJKhhuSk
DAsFLSJ/rQ9hfECVNsST/FUD6jF1UEirNBmflonmdF08iLy3CT9kjRHMxbxpHUzd
VVu6vloLsq8b8UZEA+P4eA1EtejDorxi38iOWQlGv2FgIfrXMcBzD7fZMsHg41m+
+ZgFANI367yyd70L6IdWhqryZd+utma/LoY9YzJBjcx+XpSXEZnOzce1yTWrtbrH
KkpMEZhk8PqtpV2MQB9/YfSbaTX7M00ikKZ06WVK32iPIiYGLSJSsW0AZjifzI79
/8/LshhsCe8UroqIh5rcGu+D44zCOg2bE6b385fnanvDJbeeKcPBkS914vT/16MY
p0C5eVMeupXmKPQhln1ODdfBSHZDCJVrISap4bsPVFVcPcX43NLSLCpON6ppSPrd
g56x4za82ZCxjKlGUsmHelL+g8aP+AvzrflM86Et5DeFi5cflR8mc5n/5xRvIhHe
bj5d+HmcBU4tj9fxX5Q4A2ttk+cjodtdOnSGcN0bawGo2hwPxkcSLmVRhDgmXMpb
ZQLvzfkPU/U3E8acp3G7Uzl8Jteim2ByD6jyQtH1blw7vP9kfV3xGWcLK9O/ujWq
EanYINxtzzq2Obp/ldc0ooT9G2CVGD2CUyt1tuYBIJ81bygifoFFvI1ruKBeXhHO
7GS7USkoBye7DkCYkHTY81ccfuzZZZGX6inaGm7zpD3eVC0md8eSmttFzu/siasG
Cnlkdv0HD211m07h/i92VsIdvVtqt7XwpVI0OLxXXU1ISrm0VNfJ6Ut2P+A2s4la
Bu1O+NwcGMHgelUFByvj0qATzjwdS/TmiX1u6clJLp7twDxKSANz4qFWzMJog4v9
siMU4CxsyyZKm7awljGK0eLlSJjfjtuSzEa2SjpJ6ecSC7SHjl9m7XyxgF1yiiX9
e7x3P8TYjKpY+4nNcXpCqPrcYw84CYzIjDD4MEYPFKm561vLEv4MVXcuH3LQbwLY
CPxVRpuXyoKGKNA9hh8MMbh0vlKevNxI5OK/80PYYbGVbei6oL4ZuOUcJua2J7zI
HdkhNus4l4mdKAp1QoGatrUy/SfGYTmAzflgtXzHHdJrZZPL16vlfBvJPgJ7x3tU
smG/9hqEsp+jnBOrstQixT1BeH43/C8o6GfojyiPFmKu01v+b9H+qFG640vHavij
YeI2KOq4HC2DChibs5O7c0/c7e5QB8TsVfstGOD1gaBAahNMwJiiPS8afTNT/2dO
Jrw+Yh6ozx3bxQX/0omrRwSvhA/Jypbzk4J9xSMWaURgP1a46lhTmAFi2H8ucZ22
wjjIYNE4GbaWaHDcLPJdRodsDYq0s87aIT5jY6JmOYMWTc70NgjokuAd4+ra/bUY
eONCsi8O8wwemCeAlkstHi2Bx5w45w9+ZpofbM0Pk0XwXnQLmvLDS87R/VkZZpEj
8TTfPAEtL7mNMcFPD7zG3HKF9h23nUh0J60LQVCt740L6m5sGPiNcZmb47UFZHzB
LfjF10Ab2aLsKCyCe/RdKT655jEk8Ht49hoYAuyUyVHvPb0fc+N60I+y/iQ3qLL7
6vJa38+SCm7qo30QS0CSjdpOUdJme0/v73CAoBh0F4dFoUp8yeCm24qhs47yPr4p
hUAv1/zsMjRu+BGjlYt8JxobboEtW7aznoxvfEeldQGEaO81IZakskOhreV/RgoO
+kmn4HXY9ElNTWD02qGKHS5N/o4oyOiKEzr67bvPObs4S9+YWBCNpDiOEpHVz2M0
nVcpj97ohPgf/3oHlIw6Ibc763IleH1hU361xtmXYbIKsn6Sj6AcwREz3DJRyttm
DS1HswcTzwQy9gUozQf/674vW54MAWqv5lUE3DjVN9eIREnRa/K4bkYEL7HtEqR3
3vn6l4+uUIZ5qAYA2ZETC46sfT9faKSGXEq/0XgzYAuc493iVg1IdWX2QJ+ddIKn
36zc9D96dsluuDXUb+9Ms4T4MVf8RxdjBSX6H6MZY3fwY/FbIsfwwla38GSMImYa
xRptvO1AwkNFzjhr++EPSIVY+3O6iJ8+sEEz1F31Sq6HgNaiFkRjTtTNHdJpgOUd
Nc5c/1cphG2WdISeBFqJSI1OM6fmrdzSmBo9SzTHqsEjQL7GmRRXayUKpWfrpvca
8oPppNupziFcfrvO7qzcMCH5FgfM9PChriGLBx+eWZz8zpbHeuUYopPA8gG4Ob3C
noxXuC0zX4GgiSqL/zXMbpxAmb7vizjaGU3z96SYK9u4sCMP0q3oiW9+U1dpuGGI
zvjl7FLWvf92NmAIybqsLC9qyhGaIeUpfTxh0UZGGY/fIHjphJ4I3Q5TgNd8JrjI
z98oCu3zm4PcGuZeXzDDcErC2r8v+1R0k9/ThQbzKv8zlwD3jwlfssSO0XirSR3b
3Q5piNzxB5lN5QLjmuC/Kcuac2I+xDfd9QFtD6c8+5J5BJAgJg1wabf2N5Y67IjW
IfXjstkghSbjAXuIPyse9gLEs7ikSX3nMMuUs9QyPG9zef6djsfLfTJHed3xjF3j
BaxynwA8rvWiRvKcP1Niw5Dt0Hf0k1cq1FH96EcA6W+NSlqz2myCyXtkGr0ajGgc
0tVew7QcNlfB095+yngitbJqFujJ+iVy425e07Kc7U0hG24Bohb6u4on1wMgCzwP
ofSDDx5uvKEsednIdt68Lj1Sa9AdwUkgWeOcP7wmxEWfTOyPZKj4iVjMn08wuZkQ
npBThRFZMd42Lml68fzpkjjUlq809ZgB0nuP6bnbrw/FUWNXB9zMmWFXF+8t20vi
/1zV/IO3R9u8cUXbZFZeanrGNtl9q0GJ5ncGDIyNworMyvhryIAPtznB4iyxKWwn
JxFF+07FDRpe8/0Z7tLXJmq/RP8odMnpYK62igrqLmgMnCmuvzS3mDNSIP8x1CqN
Z2mmj8g9dQBOEu0Xp4uS0i9/o6tgHsglixmK+L2DuWMoHoYEYrS69bTgiVHFQFmp
kxswlXOzTYUNW3BbrREeNJUSooW/W9NSE12D1qg6U4Kl7e1xxIjpp5PAUnzuqYT1
jvUUz+W1dKtqWrjklBTfdWEdSZ0tmukf/c1FpZF82jHGJEVqaO/UIvzREo4c8SiW
3y5GhLjLRpxk1uqlNEY4U1Tw/DcQ7AKVpuHQUT7PKSJfpmTr2J2lJtKuHbD9bb2q
rkuFFNnaTQnaYy3eraOiCjD1QP7Pz9/wnMEAWfjNBPcxqVigVpTn1hcLBN5eWJ4u
3x4N0LmqGsnWb2ZuylURYzEER6RHERzKxKty74Uo43FWSVZHXljglNVjYLC53G9O
cw33J8GiNtzQlewNOFJj1yVqOMVg/z/2fwLOmwDYBrBaBwRbI42bX6GAgLEpYnvL
hVOXXZIKSVVhD6FPbk7SwKWGJICa+Lqao3w8O4Ie9SwQyQHTxhdaH9I7JjKG6x30
3qntYp51YXSx//ZPL7gVtnHGMaMM58UDdNQeJEA0cn1Q+MkdjjBq48iv1WNja98s
sdpA902Bp0MeALJAuAPgaalVsFOC4890Fi6RwjWC3OvLrcRONsHz5ZqV1zn5Q74N
+mOvX19EHI1xVDsOHK+kgPOpBPKF0DrQiOcnvXMcg2G02RT9o9iDiAuJBz7AAF7G
7KNRRf56AlmThK9/mYFpyps1/4qHaJ3LbHGfT41rpM2nQr6kou+NyimaSxA85Uf5
ForDek7IUzbLRpiP2hVxtx0N0IPGOpAbQMPGzgI3t4JfokWL4EK/7eYfO74KxvDb
+TDsjEYfmMPfRedr7ChdudgotSybz6rssfOYt4HIPZ0z5KRmMcTKWmEIAu/rp3Ys
+cO0vxEiKPzEClQ+Cc8UBaic5g2nwRW6YKeBaS+yEJXLBbjwmjd8Bqk98FFjlfhW
mL87J0BIpYsIpBwgcsxJmjBQ0LQ5CFytPKF5DgB/hZBYic2xt52pvHLcQ9Ntikck
DuqUH50q4YP+5AYQ8ldRbn/bSoUUQzNhBmMO/gDRSJIiTBm6hcnZ4Eo0ySnZmSlE
dqYVxZZUeaqLezB3rAiLhDZunJF2IDrBVTvW/tbB6av6A5x/dPxXT3SNe5UgHin1
dVNn9sGLDKkE9yRTjbpQu5uOVSCnooec0BCg30rUAxIvlo6mHORDKH1HLm59UFSi
j89fAsE2tjH+mP8we/sRVoUnwgjgkoCN3u015VNBn/oaXo/LzfmBYmWmPqfx0lHA
QPCormxO6VH/AMolnGgQrYIoE3fHKWhxNiIl0QoMqk2fcuukrGohQBAzv1YYPZYN
t90jvwOoRrbER7hW73IDlo9cHcP/S+4ESHvYtGI3D3wzFk6j5ef3Jn1gi6EEdxDr
emVAKrSvNjuiGaIL2RMcYT1th/NQ6LwY1O/bvGbXNkM15Jr/py+kzqNM2BWIZ94Q
5RVjsRf9k0XSzdqJx+T8ZjnGMSAIvHo7KAvdDYE/o3V1RFVbjnjWSJn38ovjQlLa
dJWa5U9BzwwY5lP1wQsHhLHeJgZXxWNv+wZNQJdBBnBQx+F6j7P9GE9R4vds2mYg
ERQZeVOP7MvXI7AEGmrYheBy5U7mpE5uoDJ/UEGcfdKNqS37G8acXBjSv1r0xeUI
DxsQ9i5qae8E31noFvIW93eTf25cql/8Y8eWQDuadYK19KH2GGCQXRJLn7rt2u8L
fOLUJalJSrZYp0OqTbLUwsieYA20GycxYFVovYSxB0W7js7GXDYu9TE+6ZwJAM+S
wmo4KvtBhtwE5tu7djfBhsIH1LSAdfahtQCVWTQz6DjJM7Z7foGxvUXIgwcVo36S
kMInzmdsPv8vn3eED0RafeXA/uX6jXMoNIJKYfMEuO0YZgcjUfpizAaoLHMXaHsx
kTjDfey2HjXjgqxQiQra6UWL04OR3tH1n8K0XXuWdX2nA9QX0AJ9nCK/Ov3heOa2
C/0boipVQw4JQbgeRC6xwQeKTmd/1Inw8EDpstdOSIgL90XC+ul65bnmmrdzjxNf
tqmq7GRa3jJDjzHPYnkDOJ75pab9a9/zGP/kAz3OknvGULrwGMbPG/Og5m06HE2E
7S3/vGy5lmG3dg+K7d/8BW0Ar/44/FqrzrBfOmQ4yYNtjOPSBRpfOO1KaVt5Hd5V
ubcBbND2CSOfJKBk0hyKy+DU4bTc1tQC6ewo5LsrNMlnnoFZgOV+xhuS275+q1cM
VvN5oHtS0ixvyAtRLZzvJNo9NILPj+D5/m4z2/pW/z/CmJpRE3Qo2sA1N64drJn6
Q1qhWPQ7gIDXJWP3ZR6oso/vfqj4wfrAjsRc8KIOnuR5zdF7tDFlQeeX0iVrFmse
FwswNMJvbMp/kIcRHpxogmEXUh3yuBFKXH7Q23C397Nj9u2ID5yC8W1yQjDg7nPN
VZUxc/RWKlfDj1V0IdazHL1fvTeqiCtN1SYU58EQKcqC6JMJ6a053ICG0tN6HS9/
k+L6LoKWTwCh9gUmYkIyiegthly9zM/B58MnfXqdL5UuyY6/i39ZVDM2CFzYDWDn
Hf4DPMw+L4N8b+lSPeXBzWJgDSnQ4D+8HAV7VO1Uol7N6WRM4wcSJoTIDFpWM26w
fGOlAVfGC2AtS90TR+9Bwr9i21fG331ROCSpE7oBqWghWiZjYuxOEpR/uRXt8W5n
C6vk7TwTMDre4aAcoMlPQJ/moZ+5LXrT5ABBzAWIaz2zeoWSHM3r+x7NQpzqVNn4
lZbn5KqaXmY2rXF1Ng13wYK82zzRhJCoMY7oMPb5uREllpMT362AkfHndmv4oBFn
HZJnwfDK8JnoeFQkvNkK1UOQSC/F6yhB+7Scu/ztE06qSkTTMeyXeCIpWQv/OgaX
PULqutAuF1jAPPvOznTGt/CApq5cE8OYGRdBl+0LMfZT4ShlCCC8fRtFtOgO4uwm
fD0TiQE5E4foppRcWUrL22jG/B+1NOyt7fxWfKMawOPOi6i+xXPlVlcEcTh2LHDV
c+EsQhdaKSWgz6TX/PKSCEiKqcJmlhyCJiQaiRSqlS5CCzD0cuKrwM9gtmmYKP4M
BBREoCX5TZgGFRcZ1hSOAVHbTvlRVEhIOHnlNjPMynNTiFz2Dz9MPAMamDAByflW
DT2kqTNkiveHD5EZnPwZTTdJpAf6o9KYcMCz2GLEzLK248fUwEieKimK++b6Guaj
zIbZrUaZuBa1YjMuKJ0Ad5wcsGhF4RB9RIa/Px49VTPTkDQtLm9Iqya/EdJV4ifW
ooxLCu1TXhlbSk17fs+lgYyaqGNfJQjF6a1aTMucxUDxqolByo25WtUl0OToXSwc
IYyaeYylfcIwPNkP1kXWGEBvaOTyWoioSyNexoW1gPidSbv6oBXeqm4Zpl/5KaIE
d2vr454x7y+YGvcCQ5ASJB3p3P9oWx7+ehV+sN0Iy8FdMyIhsefddi/WtyKvn+2O
1Hb6xRxyWVt9CVV+rdGgmYE1PM+UGFYLlSzVB6JKnIJCgezvVFGm2513+t2G2WIC
8nMdh4b2+fttTHRivYl0ZSciwAMnTg+jJxNz4Y728IO/pca0KgiR/zD4UJMksEuX
JANSwEs+HaYD99vFHmNSU48LahkgHVrgYaxeMT0F6RSq6cFuH1Fr7CSAwhSd6cKY
LAN4Gc5oSTUiknEvRAa8EF9NJ9N2wwRintTWoljDqr5k5CVEDVezcpGqVTe8oo03
rpHOLvApDLRh917g/u3T5o20uSmjXmaRBoeHgEkJgTR6DOnO2SJ1addAX741ojer
flaHeZ+S0zvQu0bsCJp5SOX7ozMpbg7riCrCgp7VuiRe2c7RyBKmBko0gGEEtaMb
/oPfAubHhVn7/WLmILrZ4ZOrleTWRV4uZRE7gSJFXJXTNG0SdarmuO/MH+fv1GrB
IGB/97296yUvLXc67QEdnovtdCQ5z0/qMH14p6HDUVLdMulLPuzMLDuFEzNENqzx
EgcKeF6x6m9SVMNVCmSu2EHvJodzzrKtwW/MaaGeMP4CCMXc7DAE2pt8eH6eq5ms
BKYA85tAUGjCVgFJHyBi2XKaVQTxlUV/zzjh3IGe07A8zKZXYfjWY0KemtTpuduU
B2Jc1saumWp0iXdgrTAeBYENRxf3tRYYorW5IYJvE0cCnel3rl1ONz0xK05KMKQi
6NqJ2uJnPrxSn1oNw/eM4I/zRlLiihfsGg757Ti3zbpAPlvjLRQ2oSMKAaI6W+zu
ZhtQAaLr8lXmqTLoHAMHns9n9sNcGc30MK9yqe8rt2aRVpncBUY8elJGKGmz9HGg
eczMNmAANrW/AK/RX725axoQswS8ZtwvK8SnXl7XKZXKtu8PwkwPm5OgYkFeI+vD
/8meRoa0cKcmzDPZDpnE9B3Q4ZqaXv1m3MMp1LjptNfLf+2v6RxT9GqLTruBLyPt
tfkyXbR6SscYG9Ne8WAJqEu1C+laURf5AgFmPSHJuj1nVq4eg3LkzuVluUTeNKVk
qTBPVgMrL6U05JIHgDuJaNvbKmkq0jUlSOK7Gj40V/kLVpFWWBJzfuvtWu+yPdr2
1jRTDgNRiCISJceuMAI454eXfqVO2+gn/mBU44eL63vU90fmevbt3GFelaq2+fHf
dDlJf1/oc4ppJQfVjNhLyWBvf+sVMBvqAbW0xkzeL3Ep8em4jXsIuBjZaLnjELmN
eHHMDZS1HGQcoyBEsSxoIlqFzzVVLJQspf6NmxmLNmhXGfFsCMvLwne/4CQlpplQ
q+eq0+jQW3bqFJTOnmcHuTd4WS2uqer61YU7cLFiwZ4GoTeMJ85AyG595bBdzW5h
+KjkhNhItFSvcVR6l5kHWiBKlG2NrsA3ql93DpMTDf5HslnKppdqWJXkvLkZma0Q
8OfMh8rZIpPa9mswjK/q4Z7u4bb3YLG/Mc9+VFnunHOWKn2heZMWfEf6dTKLz1lD
h4x3XVYNWuG54S1oZaipWSvEEikolfGOu7d4LeUXIb1twRBFXz9KJQq0m1Zkt4++
zSpbBPA0ffJCwWm0wjvPyHo5b7z86NQbdpQKahZQM+J62bp2OLO9Ks/GDapxrTZR
oU1XToqGWcqNu7S53AZdiPkR/IqAuG5ho/C490fZ+t1o3glztfQUcuIGlS+1ebCE
XFtPgwlWUFZP9cNr0+PKALl2V2T2XnjDtAv3qysZHQ1d2Xn2g6/N5cWDcSFUsZ+p
EzxqqjhVmFBo4jy2z825Ew6CGUwRGUqwjIW9DNtNkA0Ln88bndfZF1QgqoLITIe6
IfOZ3ofHuvf/gXwSB3a6VivJZpvjTCuZA7s1hkzc+nwKkfqxH6y8JQ7ZrisePm44
wkVwGfYzi+w7VwnMjQU9nyND2WB0ym1WTpOMwjtCH+/BBja5kNbTxXlU1EtINWDp
EEcDtkRvLxg/s6YN0LvV80l04v59jprPntqie70TbRV4CmwUOIDmB+RjZK9MDjTm
qyqijaLDNzJPbs23KQWo+Txd0DAHNxbrE9PIcyNdBbL/NqEd7l2h+h0jpsEF3SBD
nRSLCi6fvpiHuErwYNzmz/qWDP1sp8Cr2vOJ278Y28uG7E1RTmSoDNdDO0j7VPMk
WoyrQERCvQyaGp9bYNB7cAw/V2lkVZN1cNjipXvLG+bIE4beBRF1BpAiS+CrS1WE
TIiDX28540GVJNNyKxDAqyTf0cH+zQbNRP3xHzQLwcfLqLkRs4uFpAy9riWMnIQN
iumX8p5TpEuN4bBLVdROlar3E5i8LSwvDqV/GsTE7uN6iSmIcz7FzmVg6xc9utJN
8IdOGCmCkBCDE770/1ye8ll3zmCiutl/VwBKN4ydavltNMqrtJHi3QIUQ4ep8ts6
3qAEptPaOXKpRPYPs1GZkXSY/5r8yOa2Yar7KbMjyW3jtvWycrcTOskWI9ii6EgP
lMIQVp/rXo/SHvMvuesz7vLSrc8p0ZkmFOgd85eqL8+0gEAlj1u0RhJp/IRBGIy4
7D8Ha2MASvuifAKOXBkUQ/ck/btde3uOeIgslr1CuMW2SdT9LpTnTe34qDFQU+M6
MG72jgUiioUKKrYOAWkI6GgvDnjiExn8Zi6ceTEoueYmwpxvCEoTXepo46ghXDgz
tg9whIopFx1qpyaU5t6HsJF+1IOU1f5zomtEQf0ZwNh/O3KKlDxDup0D0VDcMRJG
alZC7tiqifOxXufBrsPnJbwdY6C83b6jPGEP/LSeYQJYcIBPy25AQ1tnJ8tDvU1k
smGrVP1y42aHSkbB+/eClEd6DXbQb4lCdD/u2KEbSlcvJ9RpTjs+Z8JTKc4uzugr
SN2S6IVk8cBhd3orefeTuw+kYjWPqul/AhG3pQuJbmW7VTS+GpOzPlrpgDPC68Px
yRS+PxyQXhD4THOZ2l6XnQ0I9Oz+/hj13zL7nxrVhUWCisT1IFrIIxL4OdM1zBow
5qa3VlHnPeH3dwbGNl+LcYlUfExM5DdpdRmqiyLsLnoL4bSfKUgs2Me6PzJIT5XQ
Zv14abX3RgeXsX/q1eRfii+pP37GWATzHNc2YR6hdX1TAIp+g6BUyOICu0Edsguy
ZiskPD4HK77aTLZsYRDe22OdJv+urvRLqP65ytX+SsPOQD6r7rE7OYMSGlBXD3t/
Mu36ffvGLQ4gc+fK5Yhc0M6e51vAKwlosm8Q8Q8ccE/azLcyXLqijzdZ8FANaXfG
hgG3FmUjE1/dNNcC0cSrGMOgxdeouc1sf2EjrKQqPxrKyExqUDv4fZ699mIXjC05
rKzP23A0syNCGW68/df7un2VT7pnBYrgPWrKU4f3JHyr2NEPxkak92UCngXckrBI
mO3umZaiZIOMWa6zTPaug1d6xN6xVMXos0mGeM+98QYLC9qMvh6mN4HHLPNexIBe
aBb8q698yjHXkkCLmzz5swetZSxl6WL/lOHASDF3j41DsgDrC8W8TpihVIsY8hV7
bvvB53p9VWQlg2lNeRaMRNcGSYC4e7F8En04jv0uabJO5CKYQKZ5uKYcZs5JWIeG
l7mdQe6F9G0e/hJZDKjrMMrAkbMoxxQZy8wJFpTfAX9L+MPaovyqUOxxK5bJyAgf
NBonX49CGmrVoWibBfHcC56GPmUin2sNTXDBU2tDbAzsv8/eiZPBt9Fn/MBqRIf/
+x8YbGueibOh+1fflwF123mo9Z3bWKUGM0ECIbimV6QlrywQhx7n3w7v0+D3+KH7
/vno4NnVUgBXOVHx280GNLsNSRHIWgw5FGqSfwyknFOpDfYEUVQoiDK+U+w6dCXz
LBgYJ9PJbZApm/taEXySpEMblGjDiCKzLydAtgZruMjA0JJ2Q7kdNTnxaoF/3g72
o/H5bsIgQK/DDwUZ3CTxGdKXxWQaUABuEVo4df5Xyc2rM1kcXxRhHAgXbtarXO+D
t6yjjXp9ytEFJDjso8SCxJiFE/hS063ZEhS2rF3VyZYxMTRPRw1i4TSU0OZzU+cI
J/Lc9a2h0mvD6sJToG8J5ABh+LNEJvtvx4q1I7Zvmq8Dx++qufzzJ0UTJgE5a3rZ
CaWHtHIB3lQxIDpCKG+N+C7nX++N8suXIPe63Y8A3f958ScnhzL8pyH9PMDeEGy3
R8HchKLpxBRx3ExWKes1zGsyXRe9kLZsKuDp/I7EYbyu1uO98P3Z8Wk+bmVpDd5o
5QX3pL3jsjcGttsgLBPj37jBby1mNiydHF2q7bG4Tbx8czdm8BwLzONGXh8wYjNS
go72EQDcDkk7QMT5GwOvOGh1SwUhi3JfMf0ce51FCaOIs23OFprXMo5Rlyoj2YTG
FhISI204BqZ2LTevRgdLNlLVR5iJ22QSEFugGtGgwP23HB9wmt85ePNF8yxp5Tk3
4bbNbG3h0X55uxk17ht9tJWpF+syCpU81XTgCAg+dzYk3I4fh7EDCVpLNiYPvhCy
DC/Z5VZqvvQuvoHib/1bHegpo7KlfEQi+uaziOY4pYK/ZhfBCbDhZTFayy9g8D38
4nplvgJw0+zfGNeSqJngTZnyKi+UJwZ6v+3Aa1th1wAn5z7AJqfzXpIRtdI4RM0U
0gHRLxdS3H9wRTVnngZfD1m/vagzBGmz2w7YFSQgP0VUvzJOdarnDFCcpEXW/d+V
hGMZ9eY87f/vqMLbWGnrhe8QputR5bRcuGT0Ehj5jwyPH0khwunRYH8TxU87QLoS
phQ775DIckow8aPWb3M/xx6m4t/dlTqI/olwvb+ldJtlhR27cyjlToHrBXxwcMYz
jAIHN9uWHgCZp1gMyACMcVKMXeYni4LmtNh7aGodoGbRQAd5w8AFLYaWoga2Ryzf
mBn60qwtDKOVfsxXbtgk6BpTSqHsn22Ub3W6JtvzwAMUjFA6BUlaDmRfTJlsN9YA
n6vssWgA2XmeI04WJjPOlAuJLzcVas18ZdTTE8JdFEUx0+nmZlf0ujSsxfa77KGS
3CWMWhHi6VtjvVpuozFL08o7xhz4NTyLcbu5MDEycoWb0/wdtmsKdLYs0D0wA2oX
aV/YAZ3aL4IhGJQJiaj2OcRcc67p7ZGALHNECqalzfBlfNBWfClPaag5GaZPs9W/
i2L6N7iRtsbeTzFvPlURGvlawZpqWGwXmqf250MU2QDvZbArlHxQVQgK6wyNkSRr
q31ITjjcSq4AS9Oc35rhNeYLtAauQS2wVE0kc3QWWd8gy93TCYeI4YofQHFMO9BN
tGxgCicAUoRg5G8BOXIcDgHDcJ97o9O0klF7U4FiHfg0eSNu0XJCwF8fCKJqPsmC
TrFtngSDqFEqNdA/hSQi2wdKSJ8zxRJBQ1II/KH5qMf+735Xs5I3hZLYyAnzngtS
0yl1jBxWakTI/MP9SURN7e9qKGaI8FStvKOw2DJkmOWV8xiHWudM71iPjLTvYiYL
GeW+iF881akm3HWOxqrNUiN1OldkCthzz3eyG0ZZJXlGmjpnPSIMyfJbOevdltUY
0M8X17hgk91GVXgXm93HxK48wPkpuiWUc7WOU8bOf+GzjlOLwEwdSkTDaiEXlhYn
aLGGumovfxukoXCVy06ZzouoWrfkYWBwXh9xSCXCoW2ax3JEVjuu1iu4zoeIUfoL
/8JPohxO3Qlvgs16jpGPTZwXwWc5eJ4iD8H60Jn97S/e6D4RMAbRHd8jTOXlcYf/
Z1atdOkxSiOve2P1L8NV2cTm5f7EB/UyTpJV43sxZ6Wywi42+ONGolT1FNrPkMaQ
urxwKRM1rs5rJc1N9pg069b2VEFl3Vq1SJBbGgM+7qfyggxBpDMiFnA23324/Af7
fQcTTfWQtDv5tRaNEVRdcmtnqHa8T4dYr51OaygbGt1F7bwrKyRYLTur1eRc5z8w
lebwfw0AOu0ImvmPV3twg5lyzddwpgfAwvCJrNxYa2UMKG+rBMljT0dZt2dqc7RW
NPiO8gS8YCz7Q9pM3+Mx+yGRjxhmm0OcSyXki34oOeY5dPIAUWwl7H3Q2iDFxleu
LQ+Vcp14eTC/FkLUa6DPAWKwTpbbG3ruazjbGBCo4Pp29PIM4hTfc0jKQt2dO/xK
Abkug8Z9jluiCoAzVmmpJRUErDiYOd4OyD3GqkO3RRYSzD8sy1y7kmIFbKbLNKBP
GGngZsS/KNPAraJCgIThABl5O2McQkKlG0IfIJpuaQsPteyrEj2P3gt+EvDM3SXn
jjrXx4olyDZGjYKf8W2AovVKb4m3Bs+D1s8od2p6hzMFJeCTQv/ByfQeVrPrqDoj
y7yz3wiS8Q/Tcv3oISQIpr8tA+qHUIxwYXiFo+xOH6MlItuS14MIXI4FAqHA7QHd
x+xpuVohUZbZjlhvNQ+CM+9Kohs0hIFFCF4XYtNtl4pwspbiytuAwXV2vcZAsgQw
Nj5ORTu1TozUOW4Ws04t62Pijog+SCdMi/rtOZozq2yGHXF4Y4+kfswaSenkFTjP
MCP+lmjM1Z69D4A2EZ7HTiaHlsl/apkj7V/ZZYIPgYn9doPfAej1ns11Y7zIwyUE
/uosfPnWpZ/1Na+6kzQWtWtWeC1kg/m57mJ5EaZTAWy62R3Hfxaf+eKa4XoMZFhs
hYujfw6Lj6buwahfZHkrszpMqzBIVdS/LpBZQL0l5UnclN0s7D6NVSrqDANykJ+u
wFXlDq9DROmlSSPuSfvI7p8iNDV44VFVydLk7zvhBE1Xs3WdDuS8lO1A64hUUc92
0INFsGWL5K4zxrUOlHKOSHnzcX5KjbAO36CVJex3XbwrPWvlY+ikCSpHdtbE8ARK
uBFt9dEq5V5gEnjZX1batKfRKwPRx5yhXdWwAH9+MKDYgzlSDs7/Een1L3exDZ7J
UXNY1QSy739/ic2jXhhQCrTJ8HYSAC5VKqn2XzqQCh5lrtRAIFGHycU0XahMJSun
ZOnJhj9+zbNS/YfmpCIKTaMkYgHr7Xnl9VA+MsJtImlDceZk/8TxC8AJSLb76rBG
E2amJh0k41IdQKKHb+FlqJJV8gX2nF1Im5yo1eCPjbA+OnXANO6z50YqrmiedBMU
UzoZ/1DgMJdMGCMS+MZ42MdN7CRM0/4XA2s/qo4eqQI8plQ/rtkyn49avCJzk0gk
fH+ijmyj2uK445YEIGnBvyINaPOpqrBXZuWlg+1nPSH64GyAFW5MsOlgFQWS9yy6
tRYifbm2OBtGisBeydykroxGYGUiTSokO+ZkDFZvgihrbFw+vy2NuCzSIK/nFvTl
lR7ufKgOm2WpkOUAFg+hGbPlz2n8yitY0q/Sshfu0qOW+mAlMxyCSSTfXUiZqeD/
vvGvWtLhRHQkmBTRKsRha/Okzksa1w6ZBckG3IHCE9RWBJXxuP+Tls16yuWz4ote
NKInLNx89221C+xzKMfCUKTdE6MWgcazl4eMnHYSkaJNVG0sKhrF+sU+MLgYoGUw
ZVEMAS0aYK2BpnQeS3tzs97iEX/W+282/0bRLrudxCrBK/Ulamgg4UpkCWg6hs7i
9TSGbSxyHd1fDNjeh48MTcdcExSFvKS1maXg/NnGxmO2/lmuIZPbwnzkIkkZZE7D
ZEibWjmuD+C7i0VaZurlH0gsdCpAe/fvYpJ2GXkk3V22+zdYI/SOESNZRGtv6oSr
kC4LCvt9cnHaW86k8bW79ne17I5k3vlCbPAh8At4slIL9OavXZxcNRPOMq85XXdK
CmNTIJlnZq48aYERBlOlEq4KqThssHdPiadjCJTO6ze5nx4Ycfh8hqLFL2PxVJIy
6ulWmtmIH4yEsrg11j4C9flnK6tb/3H2DzVlwSvuC99kWjqCdqCF1CD48gnjWC3v
vA4sjfp9G1yuKGCjmZFpqsR6L72cFor8hbwbtMieFZ29zYNp0f/t0gR+56wmq0X1
fSAxTtP3qowkxSNMQ11FMwj1cqRxyVGPRbz+SImszB7VN9hbosltD+kVjBWcXXeB
Zh4sG98Z3J6Nlucd2I38W9Wdv0Uzm34bT/mNWzHpX+KCfNqfq4ptVtcu4fjvAEvs
QSdzCtGXdTcGVLSPAOmlTWZPlI/z3h95EUd8UicKqC/C0kfRARXnhtsqe+709I/Z
kzPFOGYecmIp5WK12thtyyWAkFs/K3REIeEvvOy712O507WF4aJJZq13AEtVXSc+
jPkraEoE8YUY9+1/EIGf36p2AQcgD4KduCJCUCWcnXUxVqGeq/U+kwR1gsAFjO8j
dQl98owOHoj11Ggns7kZtqb498agV4O4l8jRLCv/97cFZKqklcRTptr7+sJ6/nqo
o6WtlRgFxK409nIDezMQHZQuSpQyrybAI9GfYnu8Dra62kWrUfwhPFSOQpeCXCgm
IBjK6qIUdFVGZV0binudSLj71e+sn/9NZqeWpsn1e59GqJ3ajIK7lCWsJDaWQjho
tc5S7gcv6ZovVnsXGhwNq6EukiMxwxVxWdKAm7+MxlgS37GC54PErva2FwkJSWID
xME4UTzbPatzqg8rFyiFenit3DbZInz8zr79Jp7LVRpy2mRcOaVvNXO+YQ4U8K1z
O8iDWBa8rlGuj2GOtIpgeV3wcmmSSVPZhwoPOCCnwwKs4J0Vi4Vxp4iu/OTZLo14
Ai4IZdL9sI83VJSfRduXsJ3Dl0olsTOvbTAmPuL2gESQslgtKKu2VmteEJ3RUDlX
zBU9OjIjwKbpA0V2BydfmEuRMePGMAw+IlD43AeFx7BGLqUb8EF5zyZvBu5HSPrQ
eYFBJJiAipr7u3zq7i6gFNXc1mvHekLD1JHlo8iVNTms96Bhm/tnTto4vCyAQ2BU
qlrIYvTMNJaVtazahdSZZUjQEncqiHs0AG56SS1RG8pNjQXN63Pi1yHukzQ/uo+X
sCww929bjilRTV2vHB3dB3x8RTxVbZPceeV/D5buTNcTQFtKYN5vXF1Ded/jFoel
K6B9u3vIv/kLVxyn5Us70djx7dYHtzy3j8HCK11A0ljhvWKmkh3kDzycHQm5X0D0
ji4PUILtrKwA4gEUp1EXyf2kqkc+w9rNJTpTujtWEQpdKMy54b5PJzTtGd4r2FsW
TnexT41gsTRHaxWkzcLdgtGQBfZmnVu6wd6YBZ6CxfOtCnisy2TveNdjc8y/QrU5
oCGqYO7+A9VZdSg4QWmGoCFPTCBX5+fYqMklY1DZSYDO4poYtDuFfMvcxxe+Z9fi
JKrLQAttD9QUrdff1/pD5HFFV5Tzw+vDUPQ41m0CaUcrtw0jxARFH682IhcBZexL
2hNCkzkxPuCAkn2y55miVzzyDum69tzfhicsg3Zt7xmpCKjemADbSz1LXZencXDS
MTNOu5IKyekNonLHXHjWqU6pbyUdDhBoz+vFx3gmieDuGcB97uzoxU3lM54dLyvc
DBRBOVh+OlaaU3XqCS0lrPPELIl4GkMeY01d86tacsCsEZtFjmz6pZk5ItNvLZN2
QYP+3oG0Aky9aKuaNmjZBSXNG/LrHXa1iPI5vygTqNVvmpy9TBAOZkYNkT1AlRNV
XJ/fX6VOGIodk/5NdizAvKsoDnF6DcApuOtNLWMEaxkB8OkrwUmcTrp9lHenjINj
Hjl0BEZ5tmCJlYiZ6ZPR3nG0g0n/z0MvE4RsfAXT9pUIVeGvrGKt81dMSSSgcB5p
gFVWuyYbsdGLoOZ5lILtRjNEigRsh2n2zSrUH4vIjIjasXvWYAPyRRejhECS/K1v
Ycv2D5MuLztMOYK1bVKmriFUtCvo4WwFbSp+RRUSCEmWW+fdGMobnQhIA6wGsNcn
IY02g3QAIJPighGbgkCGedqUnCu8/VUblcRWq33MtLJf4laWQPAHiW/vVm5qEnav
/WpuXB2rIfOns6hEzqXLwzjiSDIXzlfzvX5MOfIF4MhBuQvTg5eRkV0BYaXRnj7r
wVzkzlLWBODBuGorE2FX+tvilTI1xtx61J5juvECkbtJhy/n5M3mSEbnrGdCnedk
USUm1XBqd5rw3Kjs9Pp1Bekq7bKauEKZRYqRp1mVEk8hTYILbymIyoUD8lTUX5a4
UN8KErZ6Ohgi+K+FYCs+unP/A5lLSj/lAXahaIION27l8dADhHZp6wkaKUKwcqhl
/UOIahxUzPWFBdfMsYK/xOYhgfc8SOlR4D6qxz8gvApHmPVRCGEhagrIK4DmXGp1
9C4SNjjvA0+h8ZnBe+Hwr+KDXbX8ra+WfQin/1GiPvZrFWYsVl6HE1gKatI/gRJj
xH+wT8YNwyNH7+x0ZYdCvNPCvJ5LBJfiuW/iFLqIKDZdg0xQSdDvqmKmUoSJ5cAh
KFL77rtX/0ILRfHRSYK8BAF2EjWYTcgca/XIqzcRFLa6DdT5tyUwZRdX8fbiseVB
fTeJbohmzcqweGqDQfd6Aj0bialnzq6xn4ufcnE42YZRBhRZKfbL+RzNHWn693HS
BUNI2Jm7Dmr9JfG+tW92R3V2KaEo66cTmXJoVw6isfma7aRFXYzyVBcxDQ9WyjjJ
cpvVqjLMc8u+njT8YB7CTaQ0oaZu/XJgi7ygYDfh49RJBXC7vTjYdgQmERJKtLMq
LNJVOF6qvAJk6CUfQWkSaBSe82e6KatDShT0RJTexwHSl+VaOkZQBKEBt0CnBGJj
L7ZZIsiwBFn0hUu+6sHD1CQCzNxfqgmdaa9473U7JzSO4z9zJ4xrNqU+S+xYh0+c
nGTpZhPw4eyg5+QBhr3IKzSxjg/YPZLE7e7BkCyEkRmtRRGk4Vf4W27kUTA9GCUD
FctloWgDSi76ca4BZkXXO0BCFekygLLJ8cogQrDpUZmqyzHXXRXq8CH49JzpRjNw
yVxlFY4y1nUHIUtMI4rgJ+qQxSVVZqTgQo7ckYVJiT2bG034npZzRdulAowkVgNB
XVwF5Rr0m7vcp0tVLT5nyuFNGNSQXop1thIE/0Y2Ck4vFR/xAP079VKhxwyP5CN7
0qSawHomTSIdTviNrdekoLBTfDumW8DewHqa0ZsiJxKM32kgvmJNsKWQYbBDP12i
AUlJhWOdH1sAat/0zFENG6C44AC1tWFhAkuCDKaYBouIOBdHcKhuJbo5QsEvZbfk
/1MMjvb+gAd8/7Gbr5X4nxWQq8ht4OYCU5jQa/x134yHof/zRw/zi1tnbCf+e39o
ddX24d0c8FAovb7pY7oa+Fo9/9hmheYnR57tH8WUHxbGCqt8818zuXGZDM8jvqh5
h8mYt9jdDSKziqoCMwZENlAI46rv7mLeQlzH7UAmWdrDBsXJjzGVx2W6S2eSoOr6
kRc052iuO+GREZnqiKy1WUykLCPg/PCJtByPr/0hJmYLde+ctr7kiCWzesyaiyRs
FpTbnBnYt+RNpCoV/dS1jZVN3H0d0K1FOdCyYxJ83lVZVVN0kYs40oCUapNXd1Bi
YmXl3pUQABt5PHVqvAywcaQLpf1o5UydDFdAHqgjeMyFG8zxglS5kZvldPFnNI4Q
zyAqTQILN5AlwjqX+Fo+h3RuT3HQPmAyER5vF/BJbX+5AiNqZz5laOVRXMynjIuE
cHQJw6AhlJaSPFn/ccRknvwlOFZtM5ZUMIIZN/6AJ/svM4CBtK2ZEequmHqpb4+A
8S92huvWurIMNAi3TUEL+KR/CKpcIa7RexEPd5yOReXwt8LEZh0kPZXyvFdpD2EG
5L8+nE1LtC+9hUEJKD1zgIx8llpZpwu1QJoTnJoQwlHBQqHnhKM1XykimdDb/5gG
k0tUVmq7zVDiiVTgMErHy6hMoDwx5Yi767ln5qJgafiYwQEvJdv7yjXhLE5y1icR
NVji+4XFCsSdmdfkTz+BJRX468F8c3bd/xWZ6kw26OJ+REbd53/rNuNG5Mjr2wkS
A9tNJ4+shq8t6EzJD1GKKOn6cBreQydCmAPU7c4IkGH4d/OGw5nh/qkZ/tlx0O1K
NS4GeuB4ayERg+v/7dMg69JEzKTapT8ryKKGogs8A9vRLuXM61kX4VMvG/js7rjr
JQJcpTA0Tbt61Pnayxv+18avG4CC2+1SX60GYABp9Kxb52K6DyB++XzHIh0DiZOV
iEYyeX3E7N9kls/SfIiOLYE0uTkdwaSxccjEBks5qGFABa0v3crL7dUeer6bGW7x
A9B7qVdquooBSUdpzdPopXVq8SWlkkgU9C8JatNNv0Ete2RPo+v6x8pwn7deK+cv
rz5Mz7ZROqy9Lg1FLbymB9paeZrWHcUztjb7iR+n2870b6jif+JAFEuReshzu5aP
3EN2ey/CvIwdZt7T+EnejZvdcQKlaZVxaHgGbCUiww2t+mdSZKDM79zqRNULyhAh
qtmZcQNG/kKI3bAt1lsaQQ9ogxC17nHRy2hsk2hsPlxRnnd5Ysvw7I2sRZagsirK
ZBG5DChxQeuxIt3Y5dTahFEjW0X8Fk8a4CITPkRdH2dbmigOK5Afmrd6a1vf2stT
Ib3MVl9RzT9oyADsywOKuM7D3M2jHbNlKZ8po5hdLIsOX7WQjiZB8vyAHbWHEjD+
TsBGMirJWOg+odzL0lkWbbpT1UaIPz9Wa3cwDsBMWzrvJa7sXWDseYj9VFDc5hOs
VXLBQ6cOEWTQ4u/Ce7YVSCFX71nUFWXYgtIa0KisF1c5srl0LZPViYM2cEkbkvnm
Kh8BKxEfxvFvo6rY+BxahORZAYfNcq4vwxr9KajqpghPRb6R6N81ZsKQ0PNopLhL
uaN9q7p39MClsdhc8i4XyXf8eJagkrEwxBlap6a08y0g0tQmqfTrYCIKreTOstwe
H6oYXoHH7/bKcnQLhKyZX1x2eR2Q1xEGA3y6Sn8xNwPV1lm9ug9SiGcX8TyCUlIB
0GkpunrCO2Kfj0bVVUgUBpb5SNQGR2iUVHEtkTEQRzw/+dxX9s3AnnxaChVSlQ4w
HnUHJIviv6W7/EaPQQQVv1grrCWp5KES6elQ7oegdbhNrwGQm08yVaoBXIlu27ct
AE8hjkYADzv+2JjDZw3A54YzRoi7eOR/1E7tl+I56Kcb+7DyK2ebXoSErQl0JFGf
wDzGET1kaxOfV4tVoKKgONk3mAx7DbBirgW8OPLrgIFaHKSmaExsMFiDz8CKts3r
pHW0ZgW5glVR2CsIJj9zoeG9J1lU3Phy33BY0bZl0McWhwJI23ZuTbqnLm38JX+i
aVe7HvfQMvLu9mxcPG6fNCBAK2UvSjaveVsSrLAxTmxxbWtNhpnfZglITny9msAH
woZA5zzOR9LlKDxv+e8amSM74Jql+Kcim2gd3qHNUWxRLlYgsOpB73BaDrZJWo+O
5L4M+S92qkCDtgHnGCYN2Yx0g+S5VcRVcXbTEWsv/mi64Co2o47Pmp2araLkUYwX
KdZIGg9zP/X2+oTXdBccMfz8x5o/0r6oEl/Pvf5G+z5B6hw8TL7nSyKgYtjQZcCp
YRksjGh2o1ZCfE9NKe57BMOvo5NzfQX+FwrixRMOuN4NCLQRtDTE99k4UU7iJDAb
aUmGQ1gICcIo+12I6cvbPHBemvyn4VK1p0b+GSQj3vhvtgKlnLeTLd65JCRZe+7V
gT/tZgr/0fqvZV9gq0voPasGoPs/VBL3+HIl8HwCpVvRaQVNtYDWBiAVgFGQj0Gw
CbDqrixow5mgwjNgryBGtWnouofo7N7MlSkYFJNkoGDhrbhk3LBnza749/ElfrYZ
XTjlbujjjY90EhUeWgQTy7GR4k8qvO7QmhOAw15evkwq6YL83y0uHJNQxpS/cb+n
S4JHs1lhW3JvQWBcpDa0pyyrXZ7lR80FaxTAtr+xgt3Iv5wEx/aDaVdUIq8xv8nr
+6VL0Q5e4xA+oQ/NvNTFSc7wyf0bG1MxveuWjfCttFiSAlIZW0TEV7qrsg4mXbLV
ClsfCQF3hdyzp4cQTCf+o3n5pwVlN935OaFQ/g/M3E77iRhZG0P/Uoy1XxSOdwiO
eqvZsQKN2WWaxWIu64C3V9AACGRrqr/h5rWRNnUHcn4GS38fdYNDICITXcQPP4Nd
qufku88fmDqjGmj9y2enacqOIaTqdRjjaZIWO0JZgFlZ95xZdjzStzUrkAFjobC6
iikeYIm1Spv/ZcWiDudduHj+bRB7/3m4NqyHSxj7WldgUGEgKqlFhHgIUtj8y2Kx
nTfdeVEfmgNHIXIWhZ0ssg2yGr5+tUmt/JJTvVyb+LnULZ7Cy16h+XEbQ4HoC7SY
VyGX5ErLCpIacLfNghgjk5PhhsLDZGdvITiJo+F4xoWSEu5eQJkp4NpzdSuH1XFF
VmBalEMLXsudfFjFTxDjjpnqJSlfpO4/nr4c2+971DuP1clkB+stM0Fgv30cgelp
4XahlUMzLepjxjNp0gBDEXqAbZY5lA0F/LFHYbQZ/uXrdtBg3IeKrmiRVHSDDNtj
IbD4Y5faWTcruIrnnZrWOff5jPd+/gAsquPIzuD1vSyhcwLkmjiNr/lCFQwiLLWL
e/NKPGGhhBneXCNNKlxZNjyBVyJwzIhLt8cWdqpwH3k6yuYfPhENxYSJ0ztLSJRq
PJeYJweElDkbe0jhCSboqCsNIKyTyfEOhogzUCpLlo8uuv2VfeWvZd0nMAXzvpWJ
gnQ37lla9qXwBHxIsYU9NBdL1BDuFPXeRHeGhUq+COACEKHCqEWQGFphjDvX9a0F
hw8KACUpJBo1IQpSHxfeMH9qEm/wsTVczWU8zBSrs+YUgNH/5PBjdnjcli47YwW/
SgsiS3Z4HWw7LIknmfKqm4qbBEilLWtGI1bCr6uhMTRnCZNymJZ0RjrHYR0ib+PA
d1m5kS9DolVITT+BuQuVuttUX3uvp5P99UHIyr9J0Q8XgiTypK7VwAk5Wr5kMMS6
FNFfKtox5hcBqQWYNWTX3opHNYv6JE4Hj6t1Ei/+GJKpuBWE7LhgjVEjhFqKMg3v
EUNHdEcCFCYmZHfNAPgziHjMDNQDXaad/C14UAfvHrLsHtuwpWsuKKAi5O/krKkC
Nz5wS4K+UmHQ8U73oxh1iJ+4h8DMwvh4yjhIX6BA4inJZjOdPw1axEV1HoZ5mN2P
lUVEEXaYaGFVDUze05i4C6PK3+H4zy4hEoLabWyzxPqHPTN1mO9X5Uu1g6V6WtEi
o+boxkSrWCtH0biGWimYkBVoae3Prt5575O9cYsTYB6eShq4UeYA0DD2T7A8d04O
D7JcWiu1VqaIZloV8S2ppCjnhnAoV61Lh3/aqDjfAnNjF/ohXCXFXXoDLs5T0pZz
WAhYBwi5WkfYptA9VQLF+/A7g2MtlKWA1Jav1LtxwZBthwOJ/yHN56DZDoONvSCD
87wUQW1LdO722GCf6lbinDZTmsehF27k5dmQL96hPxxhnd//tfoEjI6oxdzWsic7
88Vs4NOB8nuVol4XDxWxYxXW6ZyMnSQkfNorZq2LQUFIWA2Jkgm3Bha356LLpT1f
Ldo9xZUb96OtpDarp00iIc4QymbbIn+0Mbdq2KLiHd1hTL1u1cEl9szOi8T+VlKi
H9FQn7tJn76+D/KgBOtsh/+B6GNGthuSdBSkpZ7Xyj9OVnikV0sLs5YYm1GuSsvI
M51IzHucUO3Lb3zkeV4NYruxwd4gmqmj5pl65a6YMLDOewm2901syiiYuj8rNWjA
SbAnPFgVEL5O4iPDuyXsq0ezmDvMsSOG2QpT1bvVTO6JTK8eEvFBvsE4Yffc7nUs
iXoNF1RDG7eAVn+VfrXBaHR76EMp2O4ctgBazDzbxFmc88fZEJ5mTwh78C35nXQ4
+80+x+hXWVTlz/sQF1TI4xeJgc7x3pzFHxobSSUlur2+CzCwmmyAmsv669KVITKt
2xPCfVpMazdo2+khqI6NlTQZjl9NDwmZJBhjAZC+icCQRHXhn7BNv2jvhB/yLQgw
OhzOuvBk8z6cgPIl5pP6SPtarkrg6r57zy7HhHOhyasu5MS0uYeYpF4IF0fro6EC
vRZYIRFhjme5rNy5gwNfxU6Ja7HQAPczR2cFnvx5dcMNKltQC5Qg3jjlMFjPWj3o
kLocwNsBvEIdIxyjzckXrOq1vhf/0WR2HA3v1HhOP2FMg9LMR3kGX3QNfdcByNM3
2l3LmKdN9D570FWgqJ64Pi7Pyf3kV/Tju8/UqaTdi2MLcJTsXmRCVuSEHZclSaYq
2mDDrP4xdvP32KHWu/C0nFgSDNJnCEvVK6922BuhbYak2Ak4o9hd5p+jCOV55lnU
GWET0/hw+oEEs6iCmjc1wwib1BfoVt9qK8JzN9Qar1XVgV3LBbZxohIMs1SnRyyy
pplc7idPsGAnSA/E+ePNwyTGuQMA8QK6+rkhqF4p8ka3IMqoK+WVyQiy7VpdGsLx
tgURZbFhXCbGXrafMyYaB/FpqXiqJvtgehpBDezvhAAVtBFoicNBZChXwrX6saCo
ojnT0F+/oBcBUuXyrj55onDUxwOrsxP7wrcZMGhRzeg8+xrc+nG8qu+GV3E/BFs3
wQTD0yHkhvwHupYwET0iLF6q4A4gueKtxChnUoq7bNXBiXpxfwCnZZ3B39iIUjE2
/oAnDe6ud0NrpxAYb+uSR3ZYHlAQ2daQ84hJcV7Lwk2qVQlIBNq/tBC7zg5R0oNL
cB7oLwZ+sKW2PlJsWxFXTQxbxmgOV8SV+WrFXyiXbbCqRbNkJoyqtfWHyo5/MTZe
TZx9j3uyLVGk8215mzFsV7pguOAY0P729KilJTl+PX+oTBdz2Y/UbHlCAwhur43N
ky5Dze1SHN0kEVsIZOQ4LJGutMgXN8kfkNDrtsMdfCKNrmS3XKrEcS2Vvi1JYtH+
bhyhb+wxfI6KCfyHpcHMx1DymNfeXCzyiYrD60VQEQczXz+VafO/SMZlVdl8vPDJ
uysMJjn0r7wqrBAeGOKpDHNMmhlLsNECG5KOxP1gMcnjrMc2b9q4Q/gknW8gW5QK
QpxjSa6n3yMg7vEDYmyKIBWdFfJFtlcsUruFgJ/9kJj55FCr9gtOhDbLGuiy0JHu
TSBXEzDHFdfViKFvG4PUcOgQ+Vb82xowy7RfCjCRnUOfdOC4EzmDFNBtzHFIhUYT
7zhOc8SzCEEXpYZ4c9Ix3YNp4n+EP0IFPxgCzUSEYR8TzKQodAvaHhYBsHu60R2/
5hPLk7SSFFVw5dDqUDJIgVc0DXn37OwXCVrdBAv8iIsZePbYFxDI5+0DP/acPPWc
x8qPrw10rHCWLwrVGJt1az3tF9ckPBSIc8TMG+tQJsXV6r87QKjpEFSs3uH60Amo
vN8ImHvfQHhzAYMUffDdOjYkc710sJeDByKO/3mWc2bG7VWGzAErHFLYhWJi5kfG
8SovLjZv6yGg8T0g2AEQ6Gs6BbfLjgWMlQdeIEGHJF+8AzdXYCX1Iu54nknk5M6V
RuwzW8/Nsptv4KjgkDO5Wybn6L2u+b1xPLpZjP0jREe8JnR8TmTG9hBKM51Po05z
J7+SVzd7Lqpp+54Qk6D0c+0L4RnSLz01E87pLLuBq+0ak/Yrl1sbUfuuxYZ+Ly8Y
NQsqYJZcVOM4pd5ELaRyOIgIiDPXqdB+Prbev9X75ADbXKShM+89uB76YaQH2Opj
fOB1PViajnp0IaWJ5K+43xjE4vCpCJWTxXbbGSMoqn2YiVwUT+DDNSfLzBSIUh72
bvNPbTPmqhH6mhtySnkYkT0Aw8geHOBYXleS11xwmSS+sx9hWqEXT1dJukS5Jsg5
3Edks4xVA20xeK2JjS22tDTKDG0xQpbxnJ937gsWZEva9pehSzlrMI/sP9ww9Ybg
nmbZagSZf5YaNvJCQ0dJync6+IhnewS0vO8CNqSatgOWRgO/jCfvW4BQyg5DOSoP
vTf3pmgbY4a4pEqIbirKPIxXVsOXmf9DAVsSNxo0oqbjxoMKwfcYxBgPGgQpc4i9
TzyVdT/BW6JBQztKGIigtysC9T4TNG5u4MmRpGnE/Z38quDukJDTadjeurnQ97Mp
svOhM3oZdi1DL1rRb2ueTm6MbVav6V0tvhB4+cuvSBVK9+ywmvZnUNYQxA8wK2F+
0Og8Qcjc5rONA7eQiaj9oS3xq7njcxuBW1zXPuHRBzQd2u/UeHL4O/Hlc4bbmaSs
DwVlu2d32ezIwqESKkeYu9leVInLv7yNRNpWjy4TxJSWlcUKrUOcbj+bRLooTbBa
dnBObVaWk4NxBpSqgglIx9gsZATJ1QcJDOzeiQ20qHPI1SSvwwTJTu9rQNZvZo+E
CLoe4zuP7zV5MUK/FcXVlrxqGxuJJLO8+Y0I/bs2MzLC1lB+dAWy/SHyrEWqCBzo
z7+p5L3cJQ1QP7c5sWed22bhBquWz8gqvS9dEmqMNQyVG2elO7KI2I11jrwXH5uz
74qyQMAE/MqfRUoA/wxTWYOq6Ub09QhjAk8TUBbICn9XSNdItvcpK9SZ0cUPJGHt
hnxpMNnNtrsIgUIf2j+jKBhB7cZLG9Gb7x3ig0vwkaSejLvUQ+AHomEb/tBnV8Xv
cltBwaEKM5FMyM51WRTmzDBB12IcMDY4trlT0UqBufAbuDS4znVgJhZd8MSiTwV4
bUJV0TIXaueFnrx2Ajn4k7AfAbPnqZu0CbbKKo2WGzx1FTwAK+kGFP0XWSIeJnnZ
pKiW8LOWR57oNwMTpJVU2gBvua1WwK8EPNxbl/MfgdTybj6KAf5Ump6c29X4YlDG
tfKnj4A7MpeDfgpSe5iqDWQ8WfEcQpXVkla9LTGM3CCdufQJ4cWPtpTy5IkM38lP
wzxdylVzRSVugG1W06sisVP9PNsNFRZYMvjPDZTnkFOtMsFyOmPqrkyNLkRGe/T7
1z5xWoqvoc09Sjaimy0zt2XrpOW6z7T0OVmgi8yOkXdZFk6ykl3qFMt8MMFrLgwn
y+rVggAulwqaaGs9lTUvOSaW3g06wCCGwmM7AHChthMzHYNqwN3EyRZc2UH1POBr
9QolG5TxTGOvMX9k/QEvyj5mh5Ju1ji2CVibCZinPhUlEPUySSiXvydUBTNXtvc+
wNgSbvgseHnKR09bnD2deknPq5WbYBireUD9fjnU9pqP1aXpOKkW2HEPHHofnJbl
IOxDFa2H+deKGBoQgMsokRTRJZpw2K2nDaGDBviFha7NRq7ED6ZUL4XNzn8XxDkT
Qp5Jf74F03sMgRRpMkIia1+RX0QIbjMnpwVVUuT0U4+sBbJjtS7mpAD6uLMThtZj
NzynTM6JCdwgU3vGq2iyT/9IjX0npO99f7RLDegSVZ5nA7GUJjMWmq1GFjcLyhP5
qY9S1+0J8TybOdQ80aqPX3wO2dfVVW7DZvWg5qf2eRlSUihJbMqptrNVIOgE9mDU
XZoFQoTkh2Y5qs6pgV9c/fZaufcuBUot0cenz7Pj8P5nWVa90IsTFsHDCJTJPpZ9
gNo3AZ9uqXPdh/bDAS8aqF3HahpLEJPBKA2uKsqxrt/etZGZx/+iHI+gvE9Dy7QS
CetV+83rhgQbfBmPVPGEYMqHZbMntGgu4YH1R6M0z+gpBYrx6lobU52H4BgpPP6i
9tks6nTsC5iGDJa1f7U6+ebOMAqOMQ3vaK4yEPSv/iIHY0I4bZt/S1S37Mbl0WOR
48tNPNDxG44jEwQS6AgY7fh+JKo1M3Y6KD1T3phuGwM5U8veaAD/FAn7WKq/EIMB
P5GYgrUffIlsCW2eylv1yJWWTlLrNedTRJYe9lKGa5rlJRmc6FzEOO4H+ICaBkZ5
deFR0VAV1BwC0kfWeNhNsnTeJiz7fl13JK1tVikg18mUeqHV1VEnlu4fr7JwYmvs
LzqDdnWueaO4xt5VjKV3nXaQaxthV6Iuh9q2hUnPwTCNx/GCU5Rs/ta6dNa8AEuO
uH6+8PFacGFSFXZxYJZLRcWUOP9Kdmnztw/QarK95zfFLSInhMIIj0NlExHIwns4
VPN9onI+aRq34lMwS6LwEiYbyBU/85VipcrIg0ZXbYBBCcK/G9pkBhODYXWQLg1l
6UItnHikk1+N7zev2ulnVwlf4lAhngKZ7XhqsLvMrGGsLBsx4mTGmVwgJrlqI+qL
KY/GXwY8kZNxBmjPVqc/lhNPUj/8tMp2YCZRXTKvAf6GWT9DZiXSeCMBdA8CkUhh
ofuf0NLuBRk6C+tmBp33ckxnSgF0asinjjKJmFXowFpg0HdtvQJyrE9SN4VnyrHd
egCx+zxE7FjDVncCpCy6E/T4SJPEIIP+ycsAPBFb1iR+fCeAbtmYEQSpgxyI16SC
ZXMY29zAQSe/AoqrC8rCN8IvA88O1lPuvtHwhfOmPAa0U/qCTtyp2WYbIAMIB8M3
ijEkk4x9+yrD/L7MQJhMpkIBBNCAamXmCKxX5B4kYRYaQtaPDc9YyInCpZvci8FZ
gwh/Y+Wrm0JhWmShEXnhN6UQTPv3gcasIQXv0e4jiaVPn9jmGraooe9kCYjQ92cV
ydmtbKs3tGInnmMZqYym9b+zK6Zyr3xXFi7B91rkkYVfxieUew2q246inFmVwnHt
NwAvOezZSU0atc5FcCvEh5R3X1pjQy1wf16H6ro6Smr0HSRol0fzjwFKLu4yVVWS
Wx1m0Y963ZjQdHGz8myUmse/SCStaUYt7sCUClKtYR7+aizKW3GbOPOI/bFGV7av
aWYhFPQ+skSXz2bqZP09PbbtHDhFikgSld+E7gQdO2o2VRHOJ54TpSarAlENuhAU
KcO4r/IxGPUOnczW+9OK9tkWw7/gOnqU0B37EZ4Gt2gm9VnKP3X/4XtsPr9KzBJA
b8mw8OcN5XME5SjB5fj4DNaelyws1Ar/OePrL9qHePNCi92+qlYxSyLapu12NVDb
9ejCfoDxynqWIylVj5OOAAs7FmGsLqbUlF11N3jZVV/wR9m6V7eN9moplKd2VmEl
BkGWZTP24BptzTjvrlsnRd+0nuwa+NmK6lUJSFKAaUkN+NCSJ/HrP+6qXM1Xc/x4
3YG13hrZXirewRHVCQV3zIrez+634N2Iq8Fdt6pKzqDG+2OGIy81ODhMXs+jBthb
7hhLkzfz1lePHv25Z4imWxINt1c1aeF7lLcTzTYHc+KXcCi6Err7ELa8/6SaxFkf
0Arur21QI+zF2acVNPcQ0TWAg/i5yDZEk5pVXOvq0tPZyUHB0UIszheXHJly9zQl
DpZ1kuNWa+Kbc2GqQLHaphFJji9cV3DNExig8vVOV43Q4wVbCs3S/ZlK6HUX+FfF
G7b90mynDVGIU66pb5xI7yObO0ayJKUmjdSzxvixw6pZpzRIF6p3VeajA1caDUXJ
gB1oeJGHx8KSATb5cVjK4BUgw69FjO71FS/kTF3tzjZfItzDnkO/CScJCFBNSKMZ
cQRv86MRfKAwHuMrRTKKi373kG0hqpnaNR5sVdz5dAp8/xOnfOCykYXSs44tzNR/
Z3HlegVaYXWqoR4z8Zb1z7dbsptiTuBJ5FzhdGLLepGCG+Z61EeHAN+DYiq9/9oZ
ndjvdRR402c+JfsLDr4a9s74K0kJevta45/yH3etxaRj0RDBEu5sUvPF5QMUBFnz
N0IAgv1L+C2CVj9+23eiJKhCt0bycPo7kTS/2UMXdnZJzCoUz0lesxOOYCLF25ep
ZJ6IN1m015cS51ML9tOpZ5vjH9lpiEP12jLF0xpMb5qrRTWrCuVJXr0a8nXdkZqx
sZpciqgaww44FsV8hswMJgxfQFK1L7KYwJJE8WOPoHJO5yibu7KbxktjlBdeDw7A
unLjzKF0qXJyiYXh4KqotxjQsYzhZL8Oo9cQORb6CroVSG1t03RGTS4fqkGc9YFZ
SpLcmTVg4tzoN31dKa7AcoX1gBtPdL2N0I/c1vhrwL+NiHf4L/4sE94OQOQsO9ek
tExSZozAAVPDHjl5wrHj1XSqCsZ7wTNU0B5Pw+nFbfSdNz4/KU+SYkWEmr03k8Il
gB7iXFJr3OpDBUXvvPhoUtwT7dtrE+e+feILZuRR1uvh4H0bc+a/RQBYqDR7tySH
LQ/+17zkXdHlh2JdnrmbaN+z0+76Mart3BwPzJw+4db1cbEgQRjQcyyWonK7URgS
UyesyDbQFdy/BEL2GlUgqPwM1cHcMkjQg4IjGKgA/Hc5/FV/zzztneySRb3hsMhh
qxI9A1wrPV1Muta/Fe+kEIrvnTQf7UtAzxBNviD9oKoQ1UNw3U0FCuj4bZXbmFI9
U011BN6jZ8ZOZNhvAF+RTvvODuaHbXmsua3jWnHhgnEocnuSJ0gGnaESDGfKdMY/
Qg3RShthUZUU/mGS3MtB5oy2QOtCSU5o/7QsY/AUeTNzv5yJh9uVMmmOiwfF/Ozs
XWf5IJwJXeNIXoJdX69ZpqW4qDDlVcdXR1VDovlsx0ExThSvpX9Du0f2PkMCV7GW
XPM742I9+BZW0OtVKF4w2koszXJr5nKeSn3E0LvqV2MFIQEkBhlpsFl8OBKgwhck
zFyhpyohpJ6sjxsc3ITteh6q9x1bAMkIL5KXmxpgLbcaZCDqABvzvtPlfhVjSFY3
3tDq/O2tz7S1/pWOyuNdRv0iAgEPXW17w3BBTRC0V5V5TfcPQ7LPi3F8Xxz/2CHE
8kirXA0G/WaX9bxdG1CjWaXu4pCcfYTNQTEjwId6L3Ei4G0Sp+J+/SltbD1afyuG
pfxtbu7QnO9MwzF16iDb5AshT+tF6eHDdWFj+ZAAkFKxHTz00veZ60gbjmj6UmWV
csjb+E8BbOlZsEhT96d0jJTKbrfpXt3bGGZayINK89MSodlRaQzcxkRHmzLL4SKF
tHldSplCBfiPVWfNClbn+kYKsU6SGPs9/WQ14XuGuwr9HC92o3sZlhm3eJi+iyNq
SJ7+hrIoBsdIGWbyRc9BPT5VucKPYIGXi7FaZ8t7SonzCbkrbULNwzZz2rxi+n81
gBERWQyr0Pw7THcyX16W3ZYoxx2kvHRCVgPqQYgoIdud1GZNeeoK6/MpxNtifzlW
XyPUWOrFjXNMkxrXp9dhnwDPK72lQRn8VJCBpOBHdr8ELVQdSx6jREnDmZa0BkS2
AnHMVxrR2Z+FNsPAeWZB8YvAsv8dMG7q+7EzYNWQB+kJ50gvzaRcE358L/dMgPlN
50f+qaU/gKkfV7PoFaLvzgMRR4jWalOurCmjzcP3dOQLoiuI/BILItGGvKuIew5K
MzH/+21k3+fUuy9noH95L8wv632lppVio3xhelarzw0d4fJHozL3TaoeZ55S/QLu
j19M66iFhu1AUbzO73utbX9S6jyQ8buktEVAolPo/Ai7D50q02RnJzd6TPcUqS6q
1tnoKQezq30eGCzxOB2R8Gh9QXDl4qh/5fcRJY5d26VDOA8sDfKOOhUUFNErrUrq
ySurnVURylY9KR/NXABT/zjdrehEpBkUJabCHjIVcJb/vD8IckNamFmJumyC5Gam
8QFd6rhBgJX4VjngfM4pBKJW3X499fP5ilCV7Yin24RIib5XjK2WfF+qbPTBZeEG
y+fYreU79JOe83k2ND9z5NPnJtMNPWuZE5CFgjT99XIwkRMVnDIWfhGBnyYp8clA
ie0ApMMdQlZ0ZwIzdXPsN7H5pX1Z+Pfo4jDfeJ7/KlRuNP7mXGPXCwi8Yg/ppgYl
0caGz7PlsZ5bQNUcgjTzgvRcyiu/kBU9IznyyZeVnsMp8rDgUUyKseFCQkmC3RfZ
Mnroc2Eh4WZHI3ualE9d1aiAkdz71AwSFg3C8BBYrduNpBE8fKy+HvBsSfwAMI6S
pxoEJHd+H9H4l0nFk8wWufI1blZex5v37KsLlOupBnUBSPD+QZb0qZCFXQFznhN8
r2ByEkYBIuI3vSYPD7xqLd9cTMlYDqmfUaQJ0RPgI9WKbPuNEvkq/ws1lWjqsszC
qKrAqyC8KnhWQUeVNTjKI9Xzvalc5RK7gjc5IS/urBOpaw9do+eZ5AO7ZjWTIw4i
YRJnbysIcnlZ41KXeviipkaU40QutW25IPZJ2c2KRlxARtr4BlEZL31FHfMayeKD
4gYfg645Duh/TW9QK7lpHFVXq0zTjHWMy80C45WdjPpxm/CZOYUt8gvhTY0LKwsW
XhLHRX0BVCX5CItfnR8or8/yM90h02aXwLfKUzD/zG0M/Jf2B6DMTHdq+grJOJCM
G5rEjH9KqQOC1GO5ydTVbl1kNTpAc1A4Ns1h7RNDJyyrQ3cCQ4ksuTt/aF/K/4N8
HGagi6+aEt6ESjREK5x8ChifcKY5A2V5M2Ekt/n0WK/NLYLxaU5+z6L9KXUUAze6
0Y0wWMFngnzT6kwu+UKBQPI9T4TE99L4RZ06FUavf/Lq5LUMqdWNSmu3Cvp/yTGT
z3xQBR4HdES85qjqpOcNJHkVeHSgtswHPlkIxxND3/NnrcWvVa1tTZcMQ/A7tl2E
+iVLYjyn9bsEYcI0bN78StX/HerQVrgWTT0w/NonoXu4tvQIIdQTgJDNKBOHKr3+
9AaQxMv6bLknXyBkJVHJJTLihQNlWOJRGYJL+JRbAGPb7excZ5aIKu9WDG+PZqkH
aYGjqbn0ayw/SHefZ5vprVssEFRKxDmPzUCOGelBdrVRA93/hT60Hv1StGzHOYNh
OP6YwvV4P+lyIpB3izMWkQ8zIEAvHwQWuSKlqAfyJBVlceX1e7LnffudIm+LA/Un
B9/q2Rsq0A7pxmcOR/oX4Hugu99KLUB9uHnX5kRp+rls8R2VmO1XOrJoVTEocg0m
4PbhyYrW9TD2VauSKcGn2WKkXdNoWG5VpdTirJIQie1MQfGAeVVFb1OewbYtlrZM
X/3SI126ZgGgQ2IAVClZ3jMEhwBInbRk0Tx9/Z6F3FeffhAETVnb51uy1PS7PCZ0
7yh/pA+X1b9bZ68NgpHNbIU3mz8HxWyZo99qu/PSDYQISo7PlR+M+NuqMsAFSNH1
0ZsITFxL/aiaLdXa/G7jYf58gi9F5j6jBs4L3BUevNg1tIy64dZzwIUUsI9YKBXz
CmJluRXrBfAxu7CysivTub73ACTeX46zh/x8lzBxWqjtKgngl9IlbWeBIgHjG4Tt
oMIA8i6DRy+E8gUljtM6n1YZ1UXrO0KTL/4peykGLHlM0PlvW8cRZSZeKaqgJ/1O
4EqKmV+cGKD1UHOrMZy8UDOR0WLyNSMRclQh+Tb0ZnwrrnjWuvWQyAzbDvoZfhfB
6LmUDD5klJ9v7bPMPSV2TGWGS5qx9197M/mkn/ukss2TwBZ3ebmyYPJ76CjvzOql
Su4fY5SQ+LIGTlU08QNpNMJ+9QqaneS4TywjAZc/kvbrrPMtgRQbO58sF9naYfTE
wREFoKqGwlib5m7scgSqJahHNSZiU8TVz0Q/AYtlIKI6NeizHtgdGKw1s+cciB5W
vSvm4tDnxWVxEL5cub+CHgiFEGgim/bjIj9Xf/ZaevJbeyWouHFla45KslHWGH3y
Fco385TkNb6GTBkXealvw/XacsfgTRt/Z2Bm0Iho/7JvF/oSpgJjYzA9Mn130vGU
57DyTNcfF294JDKH/f+hbzI1MPq2aG41COJbpJ/ft1ftdXi8ItDWjto5PFd/ynYy
bVmAM2rUQK9ue5ZZiMGxwWFfL98D0F8iM7winJEAoORu1KiIvB91s2N7bOW1Y0gb
MkOV5KaMs4B5NVTAhn/iDjPOXZLLROI1fDy38WmOfgiTy4PuF+/aLH40WoqynOJp
RvGFhTT7Or0FyJyo8M6J5lrkN4JdBlCAfbD/jYWnLZMqAI+lRiexOYivZTqRa7e3
a31tWe+iPoI7q2PfF8yvKlDi033AHex4uO7Z2Ce33AbRf4gVPhUvGoj5G+OMg/kK
a2BvtGnef0tNwFft2LAwAfAqqh/MxR7yDLG3rVax4YmDc/Xh3F/L67Sk6CC17iz+
mKRhVELbcL5UFd2xkKjdECBgN+ecxY/8yn4QnAe1XZR5e1BAM0kjTSf8UHK+cSNS
0OnkqECyaWJJOZuP3VLD4H3Th3h6Htf1hBICPPGvGJA9JBiWxKXbZ9Y9Ac3niOV/
eQnBpi981rLf5EALUpXwLomZ1PH3iM7cq5qunL/YFJLzz65uyiyqauPqOlYKZrb2
pB+RKOFv5cNrKosKgPi7rG+oC/Hspl/Wslt5DLeyo2KygaYhO9IrsdAAFDH2tFLe
KLj5cekHKY3NiP5kA49uRtSTUXE46tQWCo9PsyyfuGqAdMPW6j0QNt6P1briXm3P
yYhZ9DAuy4pLadD2n7E1jNpG5mwx9X9INiShvVlBquKtmgjLWQBjHb2n11/AY+ij
nigwoHiTJy/FlFxFXpF45UC9bnbiGUhxCy5S3n+wODyIf+/WRVJDs/UNNoYIDMbG
0jgDehCnm/POAZ/LRfXOOExTpTkEWEjebsdWbWmtxQ2wHPLd7XJPB7XM9KUH1rQ9
SGdKehqBMJmor519ldl4R2UsxNFTRvdhA8o3BFuFj7s9iDnwoIN308Q3n/ps3ziF
fCfjF7hFioWRY0SGVTKlHrTr9MgQBEbAICqTS2DRkTWUVX+4QtPzWXp/1xOxniBO
93cIvwU8cCeXGEA0QKjuaNQumGQls689aj7AlAbA83HLQCOT5A0V9SHS5JlyHui5
ezPvzihZz/DXbXirgJtABolBAx9wJDoyoq+mF+l1ey0IOZ9v4AMDUAfITilc0FYh
UOCSrzlKp2oSWnybLVgx6emB2SzNTdg0kFyDPBqY/H3EAjddQOBAWtvAgMH0+/pW
LzzEaB9eRJcmjBonT0w5taJBxv7f7OAvj3dM3qrUqAu5gjWpHenZof4vudmMYN8f
Cn5iB1Tdrt+Xrhe8AgFK8OpbDbSVrL/FDNwDv2Ry4x3KjZp1cXav8ipSWiyzFSxb
CqiIKhQbY4yiX5hC2GvNl+y74tY+TdWJkrY6bl+GTHo8W+VC7g3/yGxSvFEKqyM+
q6vs9E77zjsSvQOzFr40vPcCFN7NcsIK9LKauN1BbfrSP6D5j8DBBwqFrcDXb9qG
q65dw9rwDr1NShrGjaR70r9x7KQKUEMI4XIcvQvJ2PP2JRWYLwHrgsXNIv432vuu
GTyDBpRITb5HSLVCAZRG6tXJjcXyjo7uugzbXkUPeCZQbk+jYBBmYOXwFLPJCB1C
Hz5uG3ocvufxv+CyQJSbyxlulSSdLHLwKKkeWcN/WJkMNy7VFCMi7GGW64MmVsgh
eZIAIrZutUVR9+93DOQnfYS94qu/o2A7+PYP7VgAFgzUP6F0JhKcey07J+JlpUTw
nJKtHJ1assnyiHerfz4l/NV9c1zNncY1pNkiBOCwzgd4PQt3wzB2yH/SUziYr5dR
jH2cbuY49yXywc4rD1hT/qM4T9K3QRPgMIRFwuTqrxG8XWe/csEcwlBpExo5VguQ
tW2gqj1RDhnzHG3fjm0hDqzC6BMHwU9AsW1wxWAaYjVuDlvRY72mQQn5sDFBtqZY
pH6lpk2T6xm6IwU9Cu+CT6oQ7WTLUIVOEIUzxxxslN+wR8NVgL3EXEqEwNVIzHI/
RQmr1r0Qg+jVbQqlN+toFk4mT8FcKhwERwGWCo5gk36EQ0BL2QJ/5TSy9AlywUmh
ECgxhol1rbjSJDMlQ27HtySx2a5ZSibKsozPOSnV+2Aofqi7ta6kFpLgv9tw1RrL
hMVZU8DRugXFupyNg2gtvCUjBe6Qu41r1QSqP+zEAUFdT4eBOuroF4NPd4AMeJjF
NXxPUJ14S5HOn58Y7O4N5tp66iJMZpZzhXbhGgcF0ueSonJMRa+v3VO1r/RGvlkV
rnGNCQU+rNC6bDiXGcLiIGfwUMEQQyEheu1Q7vNWkhDth4SxA7v4ejk6qqnxmiF8
ic00GigNDIgZgvfkhd4BIe9fmxIK2Ez0UaRDnEa4LS11mBd6A7/n/aqiFfj5/UCu
s6QHz2s3MbLdA4hhuzgSa3hwYE+xZ/j6wZLImPwsrcg/wtzNGy6jftVuBFxAaHN2
8MsvjTl4WkZXvgx75AWuJESRdnPr0XcF0CUzDIo/C+uUm5eirCKuYWadcElv1LgV
ABcTOUNMAFMlkrkZDYj5FOsHGNKWmYuTBbRaqW76KlR0QK7GO0tpWHxJ893Dg2aO
wX1UTRLpJNM0VCVg1/g718FgEMolll2jRrrwxCGLjO7Sx/WP9s6eYuPKnhJPpQ6I
QZ8s3d7KTjwFtOuq+ekRbcGAbX/j2vNvwEEOVoAlWJ6KbW1L+M11vP2ywmMdVx9+
MHIDI+tZ61A9w6fgIwCt8U1TH+EI6O4Kb//Osvs94yp/wnUT0w0Y05GlO20qQ0kp
hBHXY149DoJ4uabFHjPsLzobEG8c6Om1o03QbCcUc2UCgHd6K/YXcIGgbV0xB5zC
SAs3vsofBeojZvrfikoHKaBgAcLuWuYFhWM3OO2yHn0O2ED2NDsJzDQd9cE+O6Pd
I6w0RqnqUrU+2k/JIc0/7pycgC0++/J4CiBRrUzRk1FLtw78+mGRpkQMniu34Xlh
HoN7i19zq6DdtgSuZ/cHeaX6vSGFKJEs11pYux9G3qaOsV2+ULX/188Z76aJzM2c
DtOdZ9SLqkhgxVWvEMUXaR7xHiTIvbhvFnn4Q6jcNQoWr5be5Q5dWF7dy0OTbgPs
+H2f8kwW6IevvFkhQg0/nP3RLuc16Kai095UZ695Qm6DQDDVW1oVS4E42exuxR8Y
Wwd+n/ivvpgz9ITDuzJYNPVenG/LvL3LudDvHSLGHWKnME/kA3lLMcLQg/mzx/rm
thrhIBPBYlMNPahyVjI7RKw+Zp2gkY/y1QjURteLvCKWgTXcm+k3fZc3wsP21ePx
eiF+1/3ivW3dr/R+Q0drxOkCkK+l8pOaIYJG1pvqE00T4vucmn33iGywqW4ToIwT
14HNXFu8DgC6JvPnykyD6RhIcntfQ/Waqq2amRFRwEWydkK56Tnarfy/MtUH4I+a
yVBCXs3FX+WELhSdD3NFzUZRZg/k4q8FOkrMkwRQuQjD/yjOCOHXSfsDow+xbmg8
XhwsgtEl9Fr/zXWitNudxs4fk4jFhzpm2y5aHSa8+3CtbwPlFjSMo6Bn35apiws2
y0W/x3KggVtVA36ok7xZV+SqKRMkLVkebs4bC9GY13ssTnwcFQ0cNdA30N6DYrii
tewPAAXa0JfKzoXZsgSU2UWWWPtY6FTkBS7m1BAksQ8qy84UiuWXw27fuOkfyXdN
KvUjGWz2Embd2duW9LTB0xbfs/lu7YpcmQW4axR8fwrP3lF2feGcblE1yOLC8ok7
rx8RXOeSyjq82y75CDiQVwukMtb+K5zjHSDnpvBG8yUPsTgJ6YJy7viRpcmmFM0K
2CcczvcxZqZFOTuLnyd/DetEhTj0tyF4gL85og8E27g4weGTbTPmvMb790BoeSWv
1+kHBwkv5rPQbVE9mk59hG1GHeX3obL0N9qfurZJ0tIv4CcV7CUUQNYufiUIoEFo
LIccib+aN4HJQHN+N3ekxS+LTq0LSUtGB2nM3tGmR3XGvE2oraSlMhy/iFVMAKfn
sdW+GI0Ga/y4N8RHzvUVIKzeGL1CPgGE9rfNTCReY4w0xSeeUf+kCkmmyEYR8VjV
vjvbdKUUtqNo0Yep2+QI2H4C49xJL4ddSuereb2MsFaRwn27/jG+zl5jKoAQK5Os
C5QfMcAHa+CnCkhmVkH0Iiz21EupE8DyZQSjmM84UotYalRp0Zq3G1JaHXulgIpR
aN+lxl70RitCYS2H8xQ0now3bfCEarW0gBunH/gZQzdqUN6ZIQCsG654qsUZSQae
M9vGLUcpTEH5BxlZdm57/MiIBOUMydfo7of2LJHnJ8w0iGk+gH6VLHKiZPo0w6jz
JLIEvh0FzsNi1ODE0Qwi7PPd7iReZHuGlxOEmgADC2HpTHc/yzkxZ94mKo75Qw3S
rUjAbu4d760Lgj6ZpHJI4WSdSqjVywY0uOc0EwX0/KF20GNr7WiJqedNOwzdt/2b
P8Y0xwbTNlNbPtSje5DDADWl+zxqODhCrLgKMrw4MHm7s1/YmpOUmhH1t5NLyFKT
B2+E1uPHWj82s8CqhJpInmS0Hk2TfAot1FdYe3ecpHj9PuMWaL5rO5tcoply16/m
ChMAgAKo5VUtWWoZMgCxM51QEFitIJJHwQqvbKKNBeIxWHGe5JOAIwtaH3FCoR6f
PB0PYT8Q9e5HB2DTwNbnPSiRaKSAOT8JkS3eIXRYR/sP/9d1GNqcLLrCR/8QG6D7
ZCAgo21eCX8nyTzoiPV/M/gJ3323bFC5aixn55rVoUbGYWNCMdd3+yvh107G4718
GLQntIW/AJq3QEE/ispcxacyD1hDyni5D4DcrOBC2xvAbCETxkXBOfoEPsqQ5BEb
v7MOh+lrb7v46A5j6aK02RedZDzwQKJQ/URVTSeiCMSZk2Y9gUwArH3LlDuOuezc
xkyVmsa1Hhd+slArQYveg1f0G+eyzunh2HnnaubfRZ/lDWvKq3mYzpZsS2n1MpXp
74tGOttJEopw547RgN2asnc7chBPEAQDFyVObYUFsOjBPQZ6dxpXk/QgyFLIbiVs
gpnuuksbinknmH5g9+PRloMejhTXtu6/UDtYe6o7jxxqMQ82IBb7irurOO2D5B9U
SZ41aWKxsZFkMRNZh9iKVWOC3B63bgoi84sq9tcbwvgESWIIMTZErOKZ7/0UJ6dV
ce29Olv+/8chsYWjbo75Ec3Llus2RE+4RN62ZpoYhxhPJsOCcJPy021bd4PgvXVa
eSQiwV+U0kS5TaRK+bgWfAzYrnzOHgMGlDeqCldl3NTp4iKmwCGsnJRKK2BV4iJ3
MJFMxtB4OuxSQ3Hfdoj5+nbDKe8gzyVq7x3b7yDrjoupryHkx+mpPMwjLIozh5Lr
aMrkIK3lRAKQDPhrubjJ43bIXzwiOSPEPXCLWzc9kma//OJnZKrtmApfJhzQf9a2
EIM4mPYk3HnPzXYu3Ly6C5X9M3IgQX70v3LcV9Vp1h3PlkuwjEJ5iBuJljncjR/S
BgGqOTP8uIw+HY1o8nHI/3NxcnycwoLLaP+zuiEU0IpDQFCDHYeFQJilMykwgpIy
RznFyutc0wwJllUulIMffpdqaKVnfm1jKZ7XsBkSPljW7QGKg4V1PQEJYBF/+iTT
X9eaB3YAI9yZrXGBh1nJJEhONKgQmNH/rL5Oc3pMD2NiA6828jBE7E9j9CA5BGt4
yQ4iI702ErNzx70OdP+JKIb/aNgdZT6Y8210REe2u97mjnRjUTkA2qOmOb4LTCue
Xzic3Dsw/eaRoKOIvYV6AyAmpAFOjvQOEiT5sPtXX+WfmsYDKibD2Fomj2+8kcBu
9dIn0/PaUNYib4XbhvY2ZkP1PtUa0y33qMe38SJ57utu2IRU4lu9CaPAD0rkkCM5
M6TGT5Qqbu4J5E+rxG+wQHRJlCv3ow32D1VdttSk3wBPjTFr5RHNVHMEFp3pYtP8
G+36NZo4/1kIhLTW/sPCyKo6TJWr4C6phy4fiiKeFJi1L18bgWtXLDpiw5f9H0Kr
qgqBO1fBzjiHAOog0axb5zWFJdXBTf2vOER0kiGQcfk1UzR5Jb+O621Lxv/O3b00
Wvy8m9bfq6t9+QypjSDHsCBQ/adlncs+akqbD7yyz2/HzAi2fe5rKA6OCj0sQ2gN
Sox+mSz5b3p0zxWGhycgit9x6/WzDy2oKhIAJrxUfhOZRmlKfqh6YvuL3i8lw3hA
2ivpZM8IpPGsVNY4vnVNniOat5dF+OUyeOx3SYoh7GL8xvtwRw4xoAtRU2rwfcHD
1/rb7N1FUUuQRecVGh2Aq/k8R1qp79NVCk+nHGvPdgJulbGjDcmcCJEGxhcCggiJ
8z7CaaosT/x32qF8GywKrZaXcRC4cN3mWnHWgjrjivcTZOcQy1V6V17UfwrQR2HC
n/qaLT6S737hQDB6dt2PWDNhsNzzPGpeUO6d7omWMEO/CIt2ljAwt2JpEcor+R4t
jI/vg8zdky/KMs3XQwlli4kD/KdQg522jftgMzep8gnH7VCQk66GcbB+zJq8QiFI
ApDG9jkPpdql3lLp2TKsO0kzQtxI3dmC1e79iza+FFnbpmj1UB9Ip/FiErA+JSDy
URvJt1qSVBPmeAUQPJuhLHnVFYiSxrdUZTs39kbkc1kGjQjo4l1PQZ/CQTh0U9eY
uPhTImnbEyeinIXIUmfJgHmzPAbc9ZlnnAo2cLkgsOrgimr2D3IxdTlodUvuGPq6
tADnFlouQj5VrI0/iEI1hN/AmU/KtGzxnZYF4xWKYE4tlvdF/pDn7YuQdND7zmjf
GXNCdzTf1GojWK8tjlgL4QeXkoNoswggnqyyInXnxtwsoRA3HNfo3Mrz0v/iQOiE
TVCqWp3SK1nbfkyqFPB3AK5Wn2ilGNAxi8rzT0VEX6LaazFu8wGpIMox+q0x4jnd
ZZ/asojknK6434fpjCEM4zoF6jHLO9Pa7hEM10TVH9E6Dp5d5fNf1u+StmBL23h6
/kd7HatD2ScvwGbnlWRSEhOhTyHtBseAE0hUtwWtsEMHwItd+oJfyCvbr9kNIOGe
c4wtCHBVyFiY/W/oBqE44L1k+W/lU/+m2CG+cI9M1YaSbbgLI+n/AARrDsZH2ygy
U35Kxs2AlgvQf2MlCTIPvxnokC8flOBL9h5SsjaKIRyNR7mVIc0F5FitiPdOgj0l
z6tRI4KRDko5GymXBAXUCy3c2QyH40TyOo1isASAE9Es5udWdkO8UU3sUIVoECdC
BZnRltaQY3Kb4Vv5o5gWxqla5wCZq0sbD5wG71HPB8716CJ6m6E/Uo6SPfAT6Ss9
EWeRFxqQBZcj4mHljchQD69MhZsKijBd+hBdZCSPMfR/pgtN7r9BMRZOm3CwQo8P
2wQw7uwYVm91V80j2bXnanrJo+hQ6/XTZFzNeIizz54gTKG99PujkHaicRbZv6xs
dHDfjTGA/kgPx8anJ6pHtIwpCuea+UlB2TkdYoEukWUkOnn+Sb+ogTQbVIHczilh
3kMK7ZPG8o92Ef3yseeIEJyqSniNGw3YQ7IMorjmN+jJaYUwn4W4NHLvJmfEGrxb
rEcg9TjINcEtuepLd1aoujfPGntp2/b4u/F5DYnv4rRp0llYdcXraJWmeduvbw7c
uFRKUFuSWD3a0SLQ56TUmNyO45fimlqVST8dtqecofc3OaF59TE/PJwqhhDxKVsd
H4wpZ/3qWkVk5WJEEB09nvdQd5uId+vmmz4nNvf24y05Vj5Emq1V9lQppwdRZahx
iHpo0zli0qfI0shOCmZMs5tYcBL9QhdVmHWWFvcF3O97sWnd4pigphf9cC6cUazd
WK7d5NjDTMpsgHRMUySJPJE3UwDSjDKlGVWrh6kfSp0upRKIm9e6J2G0bPlCcikc
jXQDqJlSdjr1pjyLPR6wJ6HPNx8Kp3WCaSOw+HACz+0GMtYj7cqyFa7A0Sqsn1mI
nnZv9IEfLQaMPLeSaRugJvp2HKT0WNzEgafkkwUPZh/z7ccZFv8B5k6pa0KaeXPn
FGsEfc3gO2zUQdC11CHNPUk78yD+hTLhOAOr3kKXErk6wu5ZIwZBgBdxPTH+NKxG
E5TvLoxKgkXn5ssh2GbV3YOp9/4MZhGBx+25bIz8aoTZfhrYn5XfT2t1M18AAeSD
dXNtcFu9uL7CN7D+MXFgAeIw9rLDyW+FCHbPZ2Tz8QJ4elMjanl7lRNCF9csdJqd
sKyPr/VYnVNT/Qwx3TX3g9k81qKIxcIbt6NpCeD0Ecdwe0EaDZWVMzH04PJEmbEw
56XytQO21GSEJxktRcVcNHweMpt7TNnYPys4hHFC6tKsZ1YiRqDBiwBrlYi4vgRQ
k3uDLkS5RNjU+UGZUHM1u2lh6X2VckhMQqAWbGKHbrwIQnRs+oOHusvyislTqmL7
rxiFNvkxSoBHoxJj0i97StP7B4GJbQexvisLqeN+yAdpGtvWajEWmIyY4a2OGS6V
Ovq0qq2XYNqEPBVhX98qcgWNoX0i7qR1aaPkiSdj+cuuLZLW9BlQcj9WUvpT7Ioe
PP+wPfGReSdKlelsCEAs4KnJFlquNYc0LxE4YcTuGoPke/Q7SIr6EdAZ4QmX9drG
FCmh7msXq3TJIp3N/mlyliSXjIzvQzHyncDB8+K9156DTHnD3Pe72aB+q3nVrblF
th4eJtCPE2ULdAlHXIsKF7uN+EbWxRFcb9EMccE1pH1veAxhcV3lpnUsyP4jkriA
hCuISGjjXY51W5xrBlGSxeSKYJVUYHvmSYEd2p/zfudVU93qGolfWBe1rBE7YlXn
ndL1Ih4F5NnZcB3RpR2nEPGoIPIgtMnFHoPSBtyL5BgTiTd2BSgcRkzSJT4PArJG
E5L/KLGTCXvldxqvj4SorYNNu9vMU2uYeYkxu7Jshmi1kL+UsH4FsdZP3lNLiLSP
wq0E1fxHziG63OZweYjhb6+D/clleACrHB9vxHWzijKM5RZGYQGKflpYohciVA2D
uxjilpYBfOkDbJhziU9V2/k+3vMzn8Ebv7z9pO/2x4TJloy6usYLkwjEsrDAqLuC
wwgdjTV9UMEoAOfPlfWQjTFeYILY4PGfCNd7I8FAQpMJ8j+fA0hM8qenw+ZJ1prn
fZ7tUvK1VDAqvXkVP1YBn2SU9ssbM7D+eCdhCO/odElnL9dA5iXvelq3o8Djwbn4
x7joP2ZLB4Dpjqdh/GhwnBK2cfMRSbtk2LHZ+H20hAUhkaVMAtqOr1frRLPVaooI
WEqwgsPS0+fpP1r3XuZRR/Zx8YvQp4+A9yGEexxnNmIhsV0P9jXTGAzyhm9pGKvP
YB9xz/lg0Wa1d4464QfpSQC3mYxE1XwGdmmratiw6w/mdYhwC2U/7x8YhoPTKmkJ
/OpZ9HJo8ns/UjbGnBbg6DxbkRVWoF8ppfpn3QFKRDyZtrzfOomhRcoTvWCBNiCo
IC8+pqxyHEijlzfQIPYN8EaMiNh7h7Fs7ri4Rx4d3Fp7EW/JbBVcOIjNRgVhLB72
Vr4jgbiioBxf4liOVDSHlz4eJC3a8MpIJZ/v3s1F2OHV4pPMpF8oTx6wvZEEq3kq
n+kOHqsGZNBET/miL5J/nTD+jw01d9T4Kj4AOpXp/WMdYnQxaKDtmNxKuRgfbwaI
YY2wwFUIsU8Oqls8GS9w1GQ9I8IWpqbN2/SDpZO26czfnRPNlzp6Rv30u1v1BrA1
/FqGLnZ8vbErOK65RHKcCkzae17Z21LsJaGe2V0mrRU0Xur3RBi2fiUuav5im++E
ZJLmETyzxwCZJB6ETFSpPIr9NQzOfC2ZUQ4AVTXZRnzpJQpXuCA1NUb4o4S9w1an
KxNpXyBSeJR+MubE+3tMW2YUDp2lknNDOuQgmvuESucErvzAuqhVDmb36q+b42cP
Go4/1yP8Ankt08GlgAtC53Z4p6daE0TUlP2Frf+0EvxfQtn8MizT9eYGIth0bUMa
i0vymARjgg2Vx4XMii4fZkNT8AyoFL8ke23WHnNzWOm9evaoSNCj7cw2DprMixlD
pFPBjhUrla3WVWJkYtLK9frItbK4J3A25wfgQzMVG7W0QMlJk0A1TgeRzbCJMrDJ
PmPk85nu4ehsQCppO99ZNNaJqsx3Yw0Lqnsdgo7UQd8CMEYxXahFALztSTeUCKtC
ODIfYm1MNt85vu/TwQpHxLM8wsSoDmIwlTk4OiJQrLWJseECngyUkncIiHWNDwGq
R//6GqSzRRQ+camz6pi9auXdHWNlvxPKN1/cbrMxSeeLklHEKfJQHONAzHmCefp3
OtKVZrjvIeRZMFFhGZvIQOe1RLSXoc9gKmfFLG8eHELAwSmHeZX+A6naz2xE4SOt
WXTLfoEMI7O6y46KH1bbseQEfS3A/C45+E0oD7leeroAY11WB1zl4b6qXiREZa4W
6nWqKSi884Dq6pmbEAKJZXDTOm0OMRUc0JjAevTm0SIV2BP3PQK+Zu6BmFqNUz2X
uNw2KGsSvXLdfziaDmQvzP95E4W4St4sSc7T0T0TVqmGsN+ij2Wc7PuOfrYbn1r0
m7ddJT0Q4ixR7hUGxsJ/eOMJxuyS9sy8Y+cN3TkFfcYcClq5qNfTAxxwJ5DnQWo8
4yuw7xIU7yNW5P3hR+UDCR1jp9SlOg+R26ifOMRCCI8cYfWYO1bvTOcO2IQsT3PQ
UZbz6aB25/sb2oUZ5UeIkC20lborTsO0F3wVVaK9LHUNlodb08f0+OiJi/Cm7XIS
7x9vHdDBRXHql008ClRGdmpcEiKY8NgOPPSvnKIEcAamMVz1mrrqVYhdjHGKRW9Q
GEiq3u9kwlpigTLYVshML4cLmQDo0tRIk0R1nblYxQmJKQJ9kHSSdDCVAdcPg9vo
2HQuaMx2SeyvG57JEPdKjFZ3NKTQMumD50MSdRKbK42DUFUp+QChQebziikXAqNj
WMaUBWqMh3dfF3axh29/cKVUXJo90OhvNdh0bvQMzWFkNYtRVOErOWLw+mnItxaN
1MKl7Xa6gPTCq21B4tvuZAnC4RoP8sTjpK0beQuxHoasOlT4diqPWHkC2KnDUg+j
BsT5ep0a/gGcEoLM2dEqTE6S5pRsjA9tay1lrDg7OAjmx9+t4eOGjvs6tpIwP1jQ
4l/Z0PCVRcRNtfjsjuu5UTuXA9uOtqdtMJQT+A/Dn0TreHynW+YE6NgoU7LK4fF1
C3MajXS0zvc0hUMlk0SQo2ZCElvNR8LRdHFSz1S9kVHvU5xIpEu7A7p69fh+1ZQW
Lhn3c3HNvVJoWQY2dy45jY4ygX1OYCS6uHLFEbmd6F4CjclUyKJhjm2U6Fw2wPtM
E5Yqn4fUklQBHmQddmYrVEEgqLQF+JfmoBFcwy+0Xpak7fptyZiKRppGQMKnq/H2
vnG8izDRsOny4tb56562f8JKLKYs5NjwU/AEck1Lbi31thLFTcVriC3xFHQQCSvb
it2bv1bToWa1PkieWn7Spwnljf7x9O9fb+YbUfj31CdHEOdVauoCzLQ4Bo3pW39/
r7//6ZhkBJaU/EwNSWwcp4cY9W3apWcEHxOMaim/sMrsvIPS4D29at4q1DPg1LGe
O2eNAbf6+MOWzzfdL63OEy7O5WCRj75aNSBp7q2JTEbZ1EoIeJjWiL4CnDEcuGaJ
UOjDJkDZM5bRUErgxkV9MLyGr/liQ5S++/3fGNxztBp2HuLZGLCwTV6F7nRyLBqJ
N+3Ql8pthfRma/bTY69Q1blQzqX+mC+l6Hxytus7FqPhMsvHegLVXxcGLMp/W6zO
6DCEJVviiKXqJrPoirFV0VIoZogRXrttW5eJRfiyprAjMIiFoUBDeaCVd51ABExt
nUPATPfEs8z5VDR4ilSmItJbD4K6Wauf4dkt9EkLSI4hyp/bTOn9i90ivICkCOxd
TkZ8zJ6w2hvsSfCd9bn5ayxcYqOY0J12T7FuBAxSbDAoEOUwIoSj/YdxQ0X9DEon
/pY4mbw465Fx4sY1J7H+ueSe3x35T9Cz/2boutO1SfqfaW0qhZc5gYSvEt663tdJ
OkozAi0+Y85Xnpt0r034EQlDayyVpDcM+KreJh/lvwjbtDggBF6183VmCLGwrNHj
CsRd9ZQNuy49jjuJ8lruLemFTLn+BLvI8MFxN8PZPoIJTBeW2EhjlgnYqzmRvQgO
bRPllES6pWfxay8Pak/gVwyDQw+qtATbOp73yJ1ZpEl28BVX7uysJY0zUNQsZ7Ep
fQCljWu3E7qjJ/IJTHckqUeNbAu8MEm5KyAv/wJG+lPenIVD0XVtfwdekC6SzPel
Sqq6MYjJzBCskUVtWZHzx42wgBuuoj0kFQgpwBzfeIh9fXyqX6zYkrgS8+WAfC/1
a0/3RKU+WGTDze21w2FfegxMHqsmXgVTbPoy5wyxBazIHZpILV4vIerQWAt6uJkp
hiqkiRSaG+LyP5nTFQev01lJRGI30jHc14+Kmm78hVBqyTcFTHavUw+SDLUMVXtc
zkQuqpdPedRJh1d2UBs5rS/eqWXfQCHNyJbdK+6H/Jx2SCm0AO6H7XKaTN/O+bzA
AI6uuQuQM/9TX7IQANdJrQbZn3+8x5mls1TwOtqiz52so8rX4cfu6+bqrBMSLmnN
8BdXVK6Nk6aHxixc/ZrnUMcPbmC7Gz3mswNYD0i2RCPYz81l74rM4447M54k25Ty
ItFn9DL33yJWc2/jpHbl4Phuv9H2n3juruNGqeE2vRkYneUgfRKouF/S+1urRjkj
PDPWCmM4+TaJYJCFh20JM5z9Dny8uCAmryNwM+4MG3DVSsRAhgqSlYEux49WeVGO
6MeALT0O0xsfdSpxn09aeRT0TeEs8kgDoSmUtvpeP6znYd26ejkdPw2hbNti4LfT
LcK4VATaE96po3Sdvcv+xQiQ1i8X70oKbVsXMR0xi+FSDhRmBDygbXdPIWyQh3OB
fO4hhIm9Y7C9MK9XQVL8D1xBab6jWAWv6j9rcyZV+p1q4BMTU5ex6JjSEnwUmonf
re6ZWz4wgdr760ve1w4Nx4vs/67o3wmmoQlhGbU1BU8kmvVmfeUHuPiUZYJuWlnS
7OxBOrPc8N0XpsKKF8BfyrV8VSzMxkqIaMfVGLO10kmk0mbdi3z9g5aZxE1jKv7l
vIi+Aln8GYwbffRBD3MZks1AdlozLtE/eaFS6TKsWMmR+fTZah3LpiLrKMqgVkac
rIPhhfKn+KJ7xdodI5oOjj4dG5kDZgjnZtqNzVPnyRBg2dgJoeoAIgDY46fFU6p5
ZiSlRabrd5gCh0v9A2QXoWMj4h36nAuITJkQVOb1FKuYFsYZ4HC2nUQXHGQ8XwTK
2iyBBO0/i9wTOT0bzft7pGp3nK91U9zxksf3jPozeFEQWKhjZC4tbxXUExxF3Cer
Wos1LhExOoKgkEi15Wga4u5KQPbBDLBjxlqJ8CYBHb00tQIcKsf1GxrxYOUEhmNN
+d/CyEAZFHr5cOK8/ow7vkE5oqdJ5nQOFG4J1/q5JsOxw15EauEmtnC1clZO/gWy
/tJmQWJUoflOY0JGrVWdZVxCUiqPp4imA0iDZwIfVYWWyEnnt2a43XSZl/0oZqtM
ELmhVVrZkp+krFrg7m/1nydereTtVFaBTXSNPECZHHBada/zFqBdXw9A0zAuaWwZ
cOp6IkLbVptkJpk2zE8KE3BlHXfZU/K6cyBez9kmLWum/mpxESErO8ZP17mEEbpc
LDDnM4VFWut8LOXTkypUEulEUrGWZU1HZXhrKXg5bNqusYP7ArChNHAFxKFYXl5t
QCgYIxZhBbro262qQVpqPeQ7lJTSCNDI5yR77U+kh+51oPTZWL8nNNql2bpGUeoH
nI3bhdTRdN/wAUsZ5IIshFOH4Ecm/jRmBSC6dVTJtJLbMBmuh8w98Nm49NQUfMim
gtIWxJ0/q3NpV5TjMJhfuJAxu4dXpBCupoFbZLTbkVMAyqCLc9oc3UNPXVzFqRYe
Gxy4LEdNPSxFAmGNgF05TdCCSe9GuDGmeXUZxc6tOM9TT/JrBvWIa3jJGZXxT+vP
ayDrUVEFvAtjXq1MsvS4W0qAWx5fpTJwEgN2be1TnJKsCaFuTt2LII4olG2QD7Th
f2mscp+pIYRlMKDsBr4GzYejA1pL13HctgkKDLPOPG11i5ICvWnz/59KqJ1s/jfU
W2FOb+fWRevJ8jhCOyJbMLoHsL0QX48eATwPrHDlPbyFUggItNw6r/uRX7LXlMVj
4E5D4H28wt3y5EYztLkRBRTueWynOQbnWGJZT/1xtXPm/DmMFSeCLszQczAKr20W
WF5nKqsybRmdtSoGKKqJo5Z+BJMJKm6O+saDEmC5Z4lscTH2+lXCh3j8ZaLPprUv
iEZcAjOMCB1LAuLGu6uFzgAuBuILywmRc6jTAi6ZzdXLX7RDfjrSNl/M4AkdlM0u
u196y2TbTmh0On77Zu93HSGOpWHKBThUW+cR0cKKURQHWvN2zc22kQHBwRGU6b+a
tJEJ8t93UT2NbF4/DltSjGAwg3kxXMOgLtO11olOyn6MPfjJAr+ezcipA9fIE3/7
0Z86uLGe7KCD6vYgvmDwz2dxhlJoOOKQjUypQjKwx1GwJFzEus+FLuFjuoBpjVTH
wMqcr+rXcqg1VcE3/vABrQ7n6fLjRS4UHCCEFeBAuOASjIczDLYMLM+eJTjFUhBn
wRz+h/HfuN4PdV+pGmzBinABeh7zdpeF5T14wsU/XBqUF+BxbuprVRuGB7nh0FcA
3AIGFLRz/Mr2CJ12RSe2XtC8hztukfM13EIxgUSjnpYkR/D1rG4mlyt0bFrudhNJ
7Iq0L+PSP5XdHty1dWG+NCLep+UNbpPYHgFQU8p0gs5qmvkyF7qiKdTbaPGv93Mr
exRoS3v3+RZajAm12ypxM0tFcSM5a6GKp1XW6UhqJnj2Rhoi9LWwn1ejXMWgnIfa
SQkzGleUhzz15dmcQ1mpTqUmxr3MgHd+yPHg2Fh0hrPRk3kSSPj25/qQh4AMsTqy
3NG3I6vpDbz3V4pr17PwsPiJFXNkKu+h7DZpvU1JDEqr5tpFJTeJKltj1Kqog+Gw
Kq8YZzrdmP8Kr5sYEja2WFjEcPd/+1N+TyJt0hAgPHGibTp6NnmBhDtbvh9Ee//u
eJlZnZgt7miqmz8XA6LpvObSQ5NPRIqXfZoCL/kwXAWHHOj29YHr3k5mkag4eesM
Ev/PpE+4IEstDrNs0k6MgqG6dRpUyd25hXvNI79ZvpZ5VbFZ3afeE8vsKCPiq9oF
2SG1Ywahei1N+VQlmV30jmzJV76IeL7byLcNkvKpOKjhtJKS60ddN0zVaD4dBjcz
63ClD3O2Kv9eTduwccC9iXzzP7IYSJd30twFYvROiPLpRM0SmqaWCxoPzD6xJEot
2mtrXhpwI5/IpzHDcY8g+AY3YBtxzvjkrHyeBYOgXae+mj+JTwmIREct7fgxMyHs
eJCkBVrfmbUIeH5aHl8s9Gn61z9y/ud+iQP+MnywzW5NM8zcI+ADZTpUKDinhvDi
iGPvV3fZu4vUE1u9eouqtV1GvYDK21Ih1nOgjvEAplTm/Ud12ZybVPuOzBHXleko
AHKJ5sxyif3wKseM4N/huqlPhUBtu8eB8EgrWJLKdmDe4eeWzxYHy0NPRscruja0
eA4v0OE140ZXBAvx0L1PDwyN7cb+AVkzyL/S/KJh3qYYW+b/zI1XH/nmXOj6XQ+Y
2xX+ftMXSfTtVbAhF4v1qsqJQZqCG69CunawfCrhS21oPKdesf0C8qLySr9NaUGc
ROocW829p2AwECX6fHFVDrUHhhLRSrTgQ+HDOCeMvuP48B0cOB1+RvmcDIrZIFvC
e30LvA/dh3n07b2Z9fAqPecf/o4alH0dGqCNSZe93l+fYY77Q/ua5HEtxWixlzsI
NJ494zkm26mi2C8bdjTzQPWkSv8s+0pJtTJDv47iT+Jt4sOINY7Gk2k4YIfy78n1
40q6AQ1tvrnMcL6tfzxSfI4L7VchFyHv7u7XMBXcd4jjRzYDCIQ/XlpilUEeKs3i
+KtbriRx6AukLLmg7TmLjoFOEFbbW085OWdqwJE/HK9ZytHGqyEpMZaN+Xu5jTRq
4uzdivWI/6y6y7shhLk5PiBAV5tDVgqDZW6PA7g8k5s1yP0Y1J9N2brDfEp5RR6Y
LnGV3jb83bSQIg/R2+PZI2HZqgze4aRQkAaZJzsNa5hu6D1tDWHINbBri2QXh4gO
90sQ7CzWiXrf5yzE2dP4g9FIKqAV3tuW1XpcjYmCWUb+CChqVV1tidHfbvdj4wr/
k/OMXUWtw4/p/0Bb2uK19QtZ4nduEBXHD7wwqrtQ/e+HG5gfTWhwYALc5U7asunf
rJ4vzvFCMmXcTjkXfECBBtnov/WwZK4nrtKF7QNfwoD25uMgHNfX7mgM+SIl60NR
cng+ycZFdsX/9oTiGJhb+ypmWTcp/LFB23+T2oYAhaigSHFiFS9utbFvoUm/JBMs
UWaOAJMNDDEuJgGRHGEHpEHhN/tpES/cmIpn4zwL3AGPUy4pMT5nZK5WGWiCi1g4
l7z5CiEB6vnLmb04PkbvSZ+jPUkLzoDX9PqpC4DajfpJLyhUP4nxFnWu6k6k/fBm
32FUYRp4hD+iYJQ0OMwFKt1js1NwTS9B/kUUhK9nB0D9xnRijZik5XbQaBfzuMt4
+vGfj4uXz3vHlOAfn11HFLd8HavZeUQLSnqRPe691zkH95cmyd1XrXO1R1tHa9+J
uHj5A7E//Ixu/k/x20rnv1EMBZNvKSmmajLAnAfOg3uBZ+ZQKK5M2GpMinqqELcC
0c9WtL4MJw9RklgxoJo1mufIAvwgI6sXhcKWuU96szVZF8U1DVwpkCT61j0GAn6M
MqCXxydQVARiLTnWxCVBtVoDY+gTPM5i6vLPgUiYnNRI/Tnl9lp9z6o9V9k087NX
G5BezYepPqBsrKvb5uLgb+sUk8obweT+DpJIMZ7rqxmynmSWhQj0Kxu4hZYjtyZc
TyDk3sMofhvVQz80Vk4FeDWK3CmtlZ4n29SuVXr79bfzYBh3yhl6a+U82SL5UZ8m
fAaR1pnxCrsxi8S5WuLRFoNm1ZeJw8aRSg+jSqPa9YajarahtxKBujNga2mbvPIF
XqKi3PjPL1uSUpNY9p3v9PZK4X4Ozakye348vxxG7fGNh8domtwxXFNm6WAj/etU
ZKUvcX0bwmzzRbqtFn9OiF6yT7nFHEgYM9YGEjgbGapugdoxEtWGKE3C3/nqmVVM
hzts/Fau52Xz1hHQxm9yPECRBfTBuGLpjQ26VpKPC7RMdyj4bkoTPdUUMUcwLeJR
iRLuoXdOH43bO8l//MymTe31cj7ITFJA1UBb0r0J4K3aPaTJu6WJtZqR63JMJmyt
ciTaeEtm5/Fr9PMM3+Su79vuj3HxfH7jmo/Lu7pDeyL5LaL4AUVIDjxE/Suvoavy
UJzU3DODQOzbN65gllN8gssF2XQksL9hODRoiXzO0pyiJjtAbPFv1dWSQbufk40o
F/Ba0iZLYGzSfr80BW4UALPptWfW1KaKETwW9yOBJG/1+SHC6/X1hgq/Vz03L46v
2Y4nURMyuGwi9dGzy+9q9M5kvSz+chku2wmnaqZQfGFH/Ptxet3FISb+xRGgDY3j
6CIc/7Fcv3zgPTlMqyC8e556W2cbNBk3IHbAbOfYLW7iDDnegAxO5qqpDZkC70+K
hiyKWeFz+F+RexKRqYBcYvKXUkt0MkEXD+SRP92Epz52esZv76jjZoEOk28Oht6f
axyhq8b4+CXjiOfK4U35OZHeOCSvO5/BCskJuWCalhZ372ChQv3mWw7HQoS6pEr3
jFAQByexGp/2PtrioGfE1FChuE+IFOeAvZIqYoBxWOvWdFbNXUVqSvGxQ5GgHzHK
zthfqoflo7lbwbEG96OkQ7NRpwbaOTAQazb8QGIa3ogkkoErcZZpujmC8kZOFhUg
VxDCUXDKgYhy8xBbrg2sm4bmrILDVhOA2IzASHx/xlhR/0S4DnNdbQFSU3ywTnE0
Oas7yR/TdfVMw21/gUn3ZweYteqIP8Nqmb9V2yoeu2Vq7RXwG7FDgd7hyzDmbHj5
Eyy6Z8xWaoisFT/cmVSHhbwivQmfAOxOajc09FXZnFquOVD4BoYelnm1t9ek0hT3
qoA2kQCXwHXCwJEGb+tiJhGuKjRFAw9eLDXLX1DDDXw29S3K/paIgq3n8n3U7Wte
gzDTfo/X/PL5pwHwxJQB+yuRAYePGcW82jwig6boAwTQYAMyzNysE3dKttKYQEF6
ibPWpN3kVIGsJGEHWrPxHVprSioMoNOUYMuuEIkNgCZs/2dmVebbMkAkuKSpKHk5
r1CtXArHPEGawQ0gFGZBzhaI/pUsKbtAiQ0VEbWCXqLLxZce2IDvtEN9LSNzNBY0
SDLDC0WEvTn0vePBewOyEelIqxqQyXw/Ya8GKXTckWHrWwS42xzypNrPFI8fWhJZ
Uvaeid2ePw9WZhsDlqXCxIxgLoo/RHLHHjCLVcVlY574Ooww+0445aMGpB8OGOZZ
HT8hKVUVStOJkyVBwVt2/H5JCZ6PJcuvfK9tmYTkXtr/zl0uLnFMzFrqhUqBavNW
bNQxNkNiw4hUjzX6EgCpeZeQBg71d2QxH1tZ4NTKTtpPcc17/Mz/u/h485kS2mY8
YLYOKK8KpOs7s8w9E4OhVeFO1oAwfhB2O/4uBZyHiFEC6ppXduw1DhTSmrT3bLcq
SjnGICyFEA5tEg6j5uzeMimojRThvBB2C0kt1UAfOGQZ9ePdGTty6mkudhl+7RhN
q7XNwnB+imKuXRJ6oupP80PxOq+9Ue7VIy7kM+KNUcNryxEWnZcTd/vcQSjjlPHm
91D5NlKH63F+yTV5wVm1b2GovCE1JviJSny9ziYGIlsmlMF9x3qEqD2TO32T60we
yZXcEFOt0ck/ldMkaFupRJ9XF6nNztXS1pYC25SMUGADxh7LG8yxInyJFbsABVmB
fdopE7IEHNXQRMGzapJVjiNFb6qCt5HwKH5nxKOKLk0rfrIZJC9hPKHa6xLZXAQZ
1YHrvoT14cWjUUqKgx5D4ID0obox7O5grH7jPB6PmEOJS3w78Ff0iob6lWOE+Hch
PNBZkp8FZl85jbIQv1AbYLQ5yjY4IFg+8Xs/eh9BHSlF9usVCsK0zmmSEuzvlGJW
t6npoXoELEuGPNz5EvcCZVwqAoz9DIsrJXhiZRKV5sgeVDqMq9t8B0ryUDwTu1zq
1n/nBPqCNU11xWQ750NoEbU6l1f+GPsNMbNbhxtxL7ErXjcnhptCTkhCX9Py+yAc
qV4bh7y9/bxUHLZZ+kJvKwb+I5h4g8QYWvsep82kEv8Lm1x6cFmqR6fFP09gLN8m
VQRiC/RHWdWwH06JHIzHdVbhtu30GoyvA+ublG6eyjM10+OmjEllsH1z3ErJVDwy
l6tZ1Vxgf3kCePppetsegnc2O0AOK+u0RHZlLmZYqjjTljcfsU84rzH8/tAk1jqT
k4Q3w7uqLNy72Zl8O2acZ8OuZ66Pk3F8uDBTVdXiFcyvqASUR2ja+N0Z4Xztvq2z
zBL2WeBkgPbTCUt03sHlMBzoqAFq+JfXjn3GkAMVuOY0sVZCt6xFNxAqQXhJ8qvB
y/njkis/8HW+DJ+JaE0MFwfvzQ6TlaY6ITWsxsbiFpMDZsK7TE4q11Q44eyzq30/
Zxp+n2seT84ZXLqDjIkx9zU+d1kIzvpLBGzVhYnOGj/dM1itw7dNoVwTF1BLlVCX
cviPKB04V6fuPNuy2531FoWQDiR8w/RBzU5/a7gYpoXX/tdTDY7hnTCJyTH5ijyz
TBJjfJ3dgV1NBQAY48SWiE1KisVhvQuS7xaEa64X/M5MrqOxGCQbPWREttu2IOsq
IF+wifetZTsnLuLAG+GJyXmuY1lQHAWHfgz7dzIUv423p8OQl9FFF8n/b8bJodCt
b6z4zPbhwm4d5E1Zsxzik4dbvDmooOn5NsZENKkBnRoxvJ+mcuXFclkVWj/82xbc
weQXDu0d6zZswMCeDRlyoefzxOxarmImXSiMWp/ByPKJa4wfXYcNoAfFgpA9P0p0
W8TJhodpgZKDmqgfi6KCILUs4uHysfD1ijQYBXQAmsf8aZyCxCjP4phux5ZRG/mb
/Rx159sMqqZLLfUIqCyC7Ohdk3tUGTqfCflmA2WU+jnkZnIxS8f21YCfMPtqSlGB
ql80NcmnMrTx75FLIWnjVn8sHb7IwwP418eZ7W7h5atbzqFFbWFwYCPuyTiATcN+
4xuX97ndHkVS55yyCios4IFim0h6zHjZLdgHMp4WoEYtg/KI1yDH6rfpBtHp+D6M
ex9qWx72RDJPNVKNfwHX7j+fiKuTH2WqL1PVnYtJ2PB9nBJbrBHd3e6ZCITupLzu
Qxcyf390NIawELpFrmqQkUjBfQZdFxQmPOoNZgt9ruiRJZTnR+e0pYVD/46Y7GzB
fTc/jxjs4rK8BH3HUfXZ/l/hJXkM7all1um16ho8vCEB1aiemHVo9kkAERklnG3+
AtMj41t2nv+9cIM11lkKw3ewvbWam2FnmUHafi5zNQlryOw8e9/f81dg89BPNdJT
WSg9Elh3ydMofKA1Nr8EWvafpPhNU/e3nVwaye74Wu/zybXTYePoss26WvGijEeQ
BPvnb7Y4PObSa/P38JUwtujdvtAr9P+rcSAkSfAtu8oWqyisKf5NBJ+Ma/iBcKpm
O1iHJgGNCGLI9rs0c5fzDC1hA+4XVd7Haq3M6QBhc2WjNS7gXzVZhdJiSYIz4Hsu
KuMOKzC4PBymF8yDG3LgwhWHrdvnYvZrXTW8v0rYkagPw4QrBfNCZJmFn5LK3Kw6
qPhqss47YgF4q1UsBWH8PCV26vrx7Z7n2VJ+C5mIazx+EHrayHK0atsyQ7HP5Duv
yImHmFJn1ba/7xaq0Q5kr8hsBrppJuKoHR5EPFwMt9lufVtRC5ZUx7+ZpT7KYYkL
0DBwXWcC90ggXRlnsDJUBQAS+50sMEbp82rxj/UHM8PjJMWqPBnAjt6u5PBzmlSP
tioehdEZTUdFjw7vDN6fFzRJ1UyDvGaeINQ01YeziHcwA1d2W9pNStWLWIdEPbmF
RZqaaczV3rAIRqJrPVFNH+MHUURDT1ZINPg25b4aMV32cJfQWPnIzo+MyMgn3C7B
Sy2YzhfkLbqM3Od641TKLKLQG5Zq1HdT/UnUu5EwDC0tGBJLb7oBdBIHbcfVP8Aq
rMkepl9q6jnIsrEVPW6227czAACNIFi/819kwjRu3iu+hgFss7KeM+fowXgam6Wb
jGt06WjwC2g7Wq3htSRuA3vYbndqUfLbeVVBJoek/5qFJMhvsOAd5tNFI1ECd0vn
D16PpCTMN/gVcUAGb9c7cS2VW2AV/R4E4qk7ck6ZqtTNTxeKhEx6wz23+WbUoJz7
o/WgAQAe877vjrw17DpsXd4+lMmZMNOcFcrnlwqiUR9xqwxRSu+H316Qph/alOCw
uOBWDSNjucMhAFc8Z91IEQoF4rCBtXuItzWRPf1jDw1j0mg01sbN+MScT7OWEh5A
xHZPIS+1OqrA8l6avxCacWH0ZyH4X33PoMjElyYnrbtcyQlu8Dedk8o9WdTH5ffJ
ixOAW+V+Esnv8eHvyVqhnVxVkKERm2SniKoBtKvCkzAs3oMK56lke1lPOsuCQL5Z
PHuB7pDXs2d4/b0iKSPOjNKHlCtNtLe6JpdAgRvvH++ftXAUbm7Fzscj+REYCiOp
qXg3mon1kYbsq1fP38d8fadlNmq0hAlqYvfhZP1+feZr8DhJoRcXF4tkyYAVC1zx
MgHdQV4p+W/VUDhIiSsguR6rvolwEr28goJndIlHUGd+hvovLO8un7YK5yFkDPKD
CYZDBujD4rG4uIkbeJDf3P/E1S5Wb/yW+CUQGAEDek91hVRx9lZnLbeO0UAjJjlE
w0R/UVOlzH0uojbDBfE2+HoX5vtS5zw8DhPBeQdwP54v6yzsgA5SARzIhygFTan7
ZZGk6Q12ZiwvYjSrQuQPuxzheOGGhF0DybW3QyLkRQSSklIIKeuoYeQ+JDgZUfRj
3GqPbhLoQ3TJrSIg1IVwYOINaudXKt1FWzjV+Tv1gE/3n4ZZsetJawLSDJ6ZBPRO
5OFg7o96T8ztew7ELZ8yPGdEo3I6gV3ZmYsaes+WciuvOy8Vlra+AWo2D+UbWtpK
R9HlhNjelp+xWYbpoAKa4E0voeCxhB+xJPm33ZMwNmR/jFk4SHLh1bBNULhP2YEW
ppzDVipqOnp/tglnhSQHrq0N8w5BAXQyaPMyOpBAnIaObeNkTqKiT7E3Hm8veoBX
H97LSC9/s+Vn4eIa0jbH6lsartnNHH0DB6cpgwLS9lOFVzVjoO6ecL69rmMSdv3D
LH+XEDMPp/k2W+KMIO6Y2SXVzREKkRCL7BH+Acy8/e+Z2fHJiwO0XKZ4+iH6WEJO
n0drGF1priTM4taB9fM8x0HCKbEy/K2sLieEY+IZtvRneuqMgoFoMtPhfgXydfE9
thrPS16fh4uBG3r3xH1z8jAHsex2xx8IUyNQpXc/jVbbgzJkx9reomE7pFoAxqeZ
EkC6m3zCB5OIHB232ciuJDLl99qAhZQrKFAkDejypGdoEyyLXJaDsvA1KVPbh2/L
9HKkYh+X1b6PdFPbkvRmI5wDoh1MvprZW7FE1xXCg/qWqyz7PZAyBof3K5zPBSii
TjzHlABTr/dYA3npLY/JLujXcQODqc74LpJrE4lyfGQZq56XnN1C7p2llT047ZXf
AVIsgn78aPfjZyE3F/kgNwjoT9g5QYH8q1LjCqcRxi2kRN9rYXc+je3zPC8bgnlf
//VeENeQvIc0N+SCDeAN6WlHiQq9T+IuOe0KiH926OtVfYXTx4ebXDUNM+Qq9xdB
uklk/UhNDmm4LWr3z9YcvLhus7E5mz4BEmK7PrduGYLTISFdJMvnyLFnW/6171S6
Kqh0kyBskupbdteSswohsHcb4qIu3gS8CJ4T5JOYmLYgVrCAOVgE9Wi1WosE/Kuy
hacPAySNXLwnx/JfOdAcpzJVnHt70eqfaVp4COqse2f0PeMaqu4CrCsnt4D7P+gy
v1bRRvyPqVCKicc4nyXF9FVh1TC2iEqkGwA50TRMD0FPCE7he9e43RCwKhUKhXT4
qPU7pQ3Oe7SxA2my3pgUKFlSBn1GujUXOdWOU6F5iWF4gJKfBsZuaX3nkxuydmSi
BQbw6SK4g1ZoSShrHsUrxwzqW22N6au55r2adrfBKQQWHykBPJpO6mmsB8PXJMz2
evLDHxDfsy4sFYhTqRRLPFwjlFLve37sK2mLdUdw3BleDlFEGxha+GPGK4UbU42g
rLvQancWhvm/btJmVUIHCu1OUseW3x6wk8B32GKnyAv7XM5xJzpuiLoPcKnaA1YQ
cNUdkqWUIqTYfRy9MA1dJiStT410KpTI8MyGjkMrtk1aTRjAkkadI0/Kw6HneBIc
Xur8tnneNNyXdAgDDz2m+aKsa5yonZSpL6f8b1255SR5K3yLQis4ftv8JFPBDKEr
zxLeiJNBXqQnO1UaMYpyjRo53zvd7/NBDtudkkNKxSIeUfBFIk3H8Uyt7E1fJPgK
XNGxxUTJCxPA6uXOcORQ9IXnPJmw1B+N/1uP+qz/D1VlSVPqkKaRc1t7O94IStEA
0PY+zqxigX4aiF40qroki3chJJacRsd4D744KnHq5gUl6iPnAHahtLHsDAgDHhU6
gTWX5Ol8eS7EVZeA1tp8JF4YPj32Zii2hlwXoVcW28E9fEf5H+Twz6N3joW3Z/OP
RszpWNiYWGestJP1+H34obcP728IICdTs3njdnXX2b+QE0ZBMiEtuMs/CH7dQykg
JXaSUJBfQlhRjiNcXWMiqEF64L4GOlx6KEGk0u8IhRjCj9tOWzsyTmFkBSd3cRV4
BHk6lMINwbYhH8ps17c+AXkMxJxRUJ7EVsdBElCjP08DBPnXsq8cGW1v9zUV89mj
3ncZK9tMTiTGP8GSreVsNEkrBs+dzmqAgiQXxJAcZRl+7mZaY7I0iPPjxCJtsfra
6M8AOwPZrvvxMX7QqLQ+tni4uTF/t5YIL+1NUzeLGgOHC5OZyPP064nRVMKt1rY+
U1bW6j4jrBOwqlBr80cm/9imasHe+QClHpdCzVNQRUTTcs9gTNsIoBBDpGkSq6eS
s9y15izEDtxNb5yY5qVsQoCVE2SYXqa6rU/gPVE++M3BsYcff8iEndG/fMK/Txsh
6VTgpOmne94L9xmmTbjtlDXKtDtHPG3C4nmYgt2+9r9R9SLqaQEMh22UN6oo7BiF
6z1WQniLFH9BFMozsV4Pmdf4ffdjWBQEf/nBStXbWnkvdeoopg+rWp5vMlAd6YqO
yrI9Hh/xZqfa5SegioiyJUBa7uxFFegGNS6D8heG0V9UGC4jjvrCfgGsXMvCG+/g
F8+LOmeO3ubtzoHw87yV1dXX2m/ygGyXpPm6uNeCs+ADo4Bb8jGN9SNJgv5f+k9z
QqEfwSyaG+CnJvIpLggzS7Q9sV0izcHGfl5V7tpDUvpKuugvRJJqt7R4BF4oA9rU
YSQ30Z6SX10ZSEMw52ZKtms7QNkCpLBChhkuH2KHq+9u6KC6iBRfUCo3nY4UwEDK
spl4CcbXak4eG9WZxmmjx7aCWXDSdoOp2UxsLB3OJGiYNqwIiHFv0XmODm26xJTq
VhQHLWCUzYAtSz1Hz5BxyDy8UQ/l3dsoWffDrQkNHlOpKAkbFXVNT6ZH1C6kKnDC
m8P6kH2u1Ui+84IN/c7ZizF7C6F5NbsD5+HHEQNWNTBtx469csS1vMKebv5IxhnC
w8biUuOvtS8aD+qVNRHmnopm8GxFPAjUr7kWdjqa0icJQP2ITg9nlRskN/hj9qKx
Yd+qtmQ7MGcDRt2qD7aTDEgNj+S7tUSqkHlA1HYOYgcAZD3XMd8Q38B4J+s3YNgn
7UFhwMEP3VVd0oLQQpofRVfuK7tk3KUZxzQNXrsFENyLom+A06JaRLALHgJwR1vt
ahgX7tj3g697FYOMa7pOq9QmhW/GjSfjiyqFz89C0ebsuv4gm24s/u8DOH2RLPVS
lJJ9JgI1w092Ya7tvQhj7W3LawNwwPjSG/Mi61WnBoBfmRhsKqScIEEZHI9Ac0Pt
LGD6WhkmgZ8VKxW+l9PrklyhGAwLbUX+9Qd4cspvYc/zx3z2go4DWJZVgciKZa1V
8nNPef9qT9v4xjI96UMV3yysCKL4EAdO4rBOFogL6UofpZQ92Y+MruRuJ+9PA+ur
mwSQZG78aE16sIlsVOZu9Ukdp2YNVIpQSlDrvX/FdpN07BCUvd4+TzPeD/YBretG
IJX0u/Wl8RWkrlEiG0lTk+opj808lmZ/Gfnf2sKD1r/umY5oBS7QQcmF3lOmhiJ7
hvXvqyITrK9h/51BUOm2NWq+vM04ESkcXQjZnLXDTX952T4zr5TAmnTwiIDWB+u7
5PHj+f5kjsy1Wc0HcDsKnoEWsqjEqCYPmTuld9AdvHJeDe5miwC4gLu1Y6wtmbIU
qUJphFoJhPzOZC1p9yB2Y1k2JV3hgymiqQ3xdKavc4o/rxI+gc0VFu+Hn8CsMe+5
iKnI3cC3UEeyBf6ZuYFI/6JIebis50dTVSdVXRqihkEjT58sG6FEaZhwjqtF0qPv
wGf5Zih1331Ej3VEYWcdJjL3J749WSosMQ8tJYKhPyFX2YDzV1u7ZlFQ/bWKP/BT
NXw99oBdoPzxXhLNa1U5Fnl7mbkns4D61pOh0xCalPC/za0JTiB2J1YcUq7gbMF0
F8tK8ZCbMLblFPRraS+F6QESKsmsog5yWKxi2SsO0pRpBM2lmxYwsWfHlqtjQ8Ut
b7mXbzjb9RsnOWCnEG3ftgPdYIPn+HNUixewRNPSbuHV8wqL2tkArdDjC+E0W9/n
S2J4pdGfsbSAk5nzNOOupD4eD/ptOBKaJkJyvrgtgTIEKz9+tkHWWg/MMoNC/s5u
IiVxb5whqoNLn/P3SGNAiwbfNbzrkLMGfDGxH7C6xgl0zQR8rONuPblbcp1PGWPf
Bx4DSddWP/reDjFEkWoaEvFY4FgP1fSADMSiIHm0T9QrVy/sJVfSTfcsOoNFtOk6
XjBtNHd+yOG/7t3Q7MsO7FQio5x/zhMhpwacAD6FVWSMNXYanMPbxNYglXGIOG46
4yjEFGaDQs8B/C52iDnf0uaCmf7vtgYsHqY60Ttvb724xNij35J1zJEsYdGFTY1Q
LcgUDLIHqCoZ2577AXub7+2XZ72/Uhyk3KjC/mb1BEJsGfPsFlwc7xczF1x+N8co
yLKsRAlHwpS3tzFU1F4fBwIV1OHL8Ao691nClEpYBlnqekltu+uvArX7I4qryIJj
N+UH0VNCh4mSoRnE4Cw6rRjjx1GObFs5bQGeUDYntqIWeh/pq9QLkUQVnAriJ0wG
j2FlKEYKlAD1gVEUm5nrpRwG03o7EOv/HLdZ4MdL9Xj3nbw28qbgspdXXqdJyhGG
QFOP+G43vIARLTh6y01hOXMiznH+EcfCAnsv/+KaTHL+vpix4UBe89bXDG8OqSKk
TKre1JtvcoHEVkVoHEnibBCScqn6ahm1n5ANn5iVruZch93GoclyRKagN/KdCNP1
3Gb9R74iCcZgTEoHp6WkkPcDWWzfOfgWsYXdvSt64nJZ9JGgoX/yz8ZvPz76EzRX
H3Xwj9tSRbhhP0RTAV8Bb5zRJmysPJOO1puBQXA0V/AsuSMWulmKngIc9olLEDMN
4pmblcxOhU7oecCD3TKY4wdICR3GMhW5q5oNt8msM/LytIDSq5o98Ia+HneZ/MQo
sPMcnIoKHoUlDA0P9a8NA7T7J/6Mt2Lfi+ibhAVZp0pWbsVVos5ZYfoeOmOG4I8T
efyqOmRq/hFDqSkg2LggzQ45+LH97KwWWPFiL8KnITmAMj7AUBpYF7gaQMSM/7XQ
xuHkFPOsmfAB0UZOOqW/a2tySbXfbVxba8+Zd9y9p5yGVGflz91K+64QXpm32taL
OEnIRg97L2HM5OK9WDsH1xL2sloM6DtevJefpxW1Dr11qMiw4eDy/G73caz154gT
FkNS/BjTQxUSOlKxZn5M5q42c6s4EG5uI12sALjipJ9zM8/T2tL1fXk95Ay/8XyG
9SyFg2CwOmGeMUK7MY4+CsTBwtGpulLjlhbjRxx9rzPsFbQMlCWR4xedfKV65QQ8
hc4oS/YV0Y0CME3TjZRlx+iqlRarn+zTsYobg7AAMMTL55QjoHI67DKtX8Yp7G5h
1/BCphv3r9u3f1QCnv2/VuxjPdJ8f6QuIcf3wUaeSHiDjWCPlfagzqLD4sY1jqk2
sBdFSzWDH/46YLzNDsrfQVKJ6DFM5beT66THSVtjUp6KvXOXglG8pVOripB9gGCe
HWRK4HdYQ6qewVZ3yqBF09aWBbn9YWlyCB74Hb43xwUbJmcFzFzqCwUAMDFIL9le
ldeYYqws9BDkTEc50pvH4/+aiIynFkwwwm0i45bhKz5V4If2hS2HbUfm2RkEkFwy
A2oL5jPUXh5LA0d72oHGwuJLrLNxbJ1r0t6fjq4O+gsNLn2E4B4z+0ytHy4tFTKl
jsggWTA23+tkJlxsjsOVRid3pGzUyb36Pv9YQI4wP4NQ7ogPOHk3cfGVbfWDyySc
aKx2YX1xUwGWoNGizUteiTD27m15GAI4uDVAwWpMLVd4NGgrf6eZrNCVQFDot6pL
+IXC/9e0y2F/wGdMvCCJmVDtOgBohHa1im7HF4CRFNsBcaoWnSTfQmZ7KIuKif/f
mlCRloB/kPY67fN4VkKAyRGwIdCutF+bvU1MaBtZqajnSbEUdpsoRYSeH4GuSfLw
JpfOpVa6vM8sqS4x3QlBQ2ou7/X10fi+T0tCpnBklmvI1mDPDiLP7sp0gGlAPeVp
q/qSXWEt2L5T8Em2Vn/6VpBw+pgS30zVnfpwiqs+q2lQ9AwopnB5D+1qqYId2LIW
7mIbejdhP1PDJgt1Mq7D2SM3EeQjWBLepYMavapwKeGnsl133HHnFpn+EYOzGpWy
gY9VSx4U1h91U5ZTAQ3xr+BXgKCJZ6htqqYwS8lQma3+5dmkt1HlxBdhwZf53W6E
nizEQauJN7QUJG/KyWz/rZusK1l7uhZ8dmbRd6vz0XvfGl+9dqc6MK3MDDzN2Umf
Fnr0j5VJn7tfbNS1UClghSRW+xfjWjPbNsrXWFZlUArbb7XbwfEuIEW29kVaf/nG
8kWrdoW/rzXa3W8BqQK6HRBWHBMggle2AjJEfRiF2WAkOkqca25N2AzxyWO1awoO
mnvhUQxldZD196YHVGCQUsZ6KDbsNJd9DwNUfudB9vse+2r6cu/fIJ8Re31CnnyI
DGPo5I50T6aP6G4MdMWxLc/ow1VoU0hSTKZx3T5HB8+t1UP95zVRNKyiRZN/528S
uSO6g8P8/qdDU7Aohihqox/aY+8W1+7SKPQiQrpKuOgGcO6aRAZhza0gR5LD+1UG
3BoEnQ3rQXPx4H+2Iy7i5wTCxondSTiEnfeQBORDjAfSYdBxeAOptvsd/DKpjjUl
3hjylPyYUoW1WTKhELHRNGS3Ouw7LNKBq2Ayc3JdALtCWxvWel0pMMxz5xtlsf4H
3elWOHjJy7uG5yVu1siTgkrx6l9D+mU12hPJYPN9PKeNoeAmzGiYa8aqmxy60/58
fPOO+p1M74DhWX33NS6ZGkIKx8bPQqGbvt/1sP+06mOgeHYJXH1YhhBgRaNp8BtV
XGr8uWGcXGQmB2UObFghS/UpB4uQZsnuvm0QxAVU8C/2xxPv2prRr+oDWwcQgYvQ
Ut+hBk0Pti6ia/mHmrMuaLLqzYoXxjCs9TL6ReafwHh04PuI/8VqWgBaLsW9QQ5i
AX8yXFQsZfnATH+/jEKXBDb34ujrnxoZqicwav4WEfoVOohADpRSXbfM0dcjdPb1
W3AvEl0zYWVJmhRbfVvkmi//Yv7cAx0gVITfhYu2Ux8MhVHpYvCBPo6ULX6h6O6Q
rNmQoGpF99ictJ23zOdiiQjZTHQt+fGR3Q4FkmMyZGj1rVCs8igzlOyqizXCqOAe
BOQV73cesY6JrxCLLXdHJA8fGcEKWOz6vP6i3oe5czeGx3t5qyAtFEgeWjkVhtme
f9/PWAFV5NZWgCNqLjHtrJVANO9RwAI1WauDXCqwm3kSiITRJ7TdQmJZqmgjGMAc
TUdsuw0ZiVyRswVxreCBsVrvUWS9JEpeF/O4WOfwdylvoOrxv5up/DzgxN+UFFp9
zJkUKzntNn+tDIYusq2yGh2h/jkDroKlPjoLRq3rmcKUe9ql70T+3NHnAllzy6Gn
UFTOS4gUR4Kzbz8qowCZnzoCSRNuvwd6ou3VDof2gvscTds/dnsjQ/HqXJ4PyE2p
ns75keHoCeWP+PFpiGurm0JgAi8SfzHp/um2vOaab4BzWeD6YxBC0w3fKgcmy0sZ
EAUSx+8qPycWL2X/dxxRTzdxisUfyTo7ewVWkqVeZWgbk/UB3IYiVQRw3PFfS7Vt
fyadroE/Z/YoSIt2ItuzJ8el3St5uIWRcMZqDVlGgVWpGXQpDkXoX4zJRF1YCBHL
+MkxESbZfYIvMq0uNVarf1Ju79EfPSUDZpRjRg9UsRbnS4Hxt0k/iJmaBeTTWzAM
/+fMPw88y2s0ofh1nzyS6jsnqj2adiMI/A1VR3R9fvZJvbKGzvLCGtf++ex4rhSc
ObYUmnd9Ai3eIE8XZo4gjtyBWZkoldkBqn4pfFSSe1v70XZjROwLj2tQu4vP95SD
jtLaIFsuvcPSEsFkQ+s66LE3zdB19IOhh7clhYaQGlg+K85tfRNkEJipKeCBDUZo
pZyngBVyQqEq/EFg/sYdq7q2TkHyMbuu76bPb0+wnd5gia+HudsJSUvZX40ZxO/G
u2ORAtaCi+rNIfJ9ns0NgPuRB968ubBbB7y2120nTgVDhvGN1KFl90fHnc0oEgdo
58CuHvQ9cT8v/WUKU3/rrO6ysREUGyTrYnYi0TUS8clE1EqKq8hdXUGRaAkmQdtu
tBYAxa/X5JvrOCQufneRz2ADMFycDzzqONn09xAqgZ8SfT3B2mMkzfWLKXKTCX/u
7ag8RYOm+LBLgfwl6gxXEmxzXlw8ke7CfU7nqNvhGEksrbEGSRVsLmmSOMePNElG
QVACXuQqA5vH5uKSYIbtzc08LNdC3wBIX47U+Ev+PZCz76GGaJWcyxH/6GszyJ8C
RHXBj4ei5UAXO2zgY7cb7RQG9HtdyCjn98G2fyXiyMw9rJ5p9vPLAXd9LPOg158A
mxngzkjd8vWBrUq2e9dIhTaDpK9i76vtE1IjJivmW/zM+NxOBUPCm9fRSopn4biq
4aDscU9srJHUc4kGQtVmxZXFwvEnO5fd+0li2k0NbVOjsm7jpae2RBJ+dnjm8pEq
0VYJvDdTgaMjzL/JwJS0xvZg1twAFGW/trs/Bvbxt3UHJeDWuVQT1XmzZL2r8vz0
RRLeq8RnPotAEpPwgLPx4E5G8fJvBn9/JQ1VArJyrikoT0VkXEFrkUihfT+/mAOd
JMRqdkyIK0AZhMQnfnpMmiZqEsOTWWpR3PUoMTOkqofeGukVroA7hmrO6H7mVOWl
+dvtLbahkTQ0SJlLa0cr1NOTj5Li2shX1RbJKRpEf4dm5/N16QLQVNSsJnTSwF6R
BLIVGFeYZgYkXiCLQu0OzR8dqmJblMeyABxJ+nl/tsAnjEmGXdRscA86AgTUuauk
q6v2uXRlscVY1O0JiCIQaWOYIhHBk3ou6R09ZG358Dz95YQNIC/g3VlNxTPyUELj
WtJ5tjBwIGjMzIwM0qfiF1wgNRQYXfn1/I+kYCyfJwam44t5fwOBDjEzsOjbqy3Y
FT2ikYLGm8C5KoG7eg/pAPWy5sjIhgYi+41uqB50KjX2vjkk1C3iAcl34VeMk5Ah
YijC5I9/3BL83AHso/ZcaYIYG7HGOO5HnYw4bOe2mTYKWEPqmfoleJWnUSwbm+XF
uyjvpfRnqClld8pNnI7/xLs7+hgndFur283oanIQjO46zqjCSDM9HhAsQWH8ypzo
mLFYkjT/adG2thkt59Jzd4pcf7bVRPxxEYwiWRnWYzVNgLiqPMt6AivKhCSsBWBv
3oOeCxhCDuoApDGIFmVP750qqd5EPm4js8/EquW5Q0ONkBssrN2zhGiWAySERTVD
r0RHNDMkNArrinjedUQXQmr4IERH9winKspHBJ+hEw9aGPQDxuKutW1N62OKIlFS
RzdxG4ece7hkuo3PM7cj0hj2PKN6i9QBMaNE9hy/s7yn8J3WJNZT8kK8+jykbBTq
gRuyPtpCMrv9V5UUGqI16qyInEvPhsa77sxM077lawYcINsniHrjtFCU78/elGju
vOr+1tceibzEJn6yqoqntzG/vHztL3q+wQ755mYUK5Lr3Bd39qDhz9o53r8zChyA
+VHxXyxBhWGF5FD1F1WmxLuvpnu7X1GlLN+ptTRzjhRnlNWx9RfFDrhtfUSQVewj
wEre8x8Dy5HuFJttn/ce0YIqSWIfJqxy8Q80tiBA8uMYzEQ4l4dHAU10oTHeL/ik
pn+bUQBxEk7zv0pe6ovg+f7BGP4ItK8syieVXwBlbJ1UjEvcToXVqCd93u2G/F4K
+wXmWHqTj4vqghT8bN6YA5JO3KMkY3GH7y+EUKGwNoUUlNit1hIZcZ/42OB7FXmj
CTR5XvWNFmNvGiGsvLGSIUQpJj0CsAV35RbqHRU+3Kn+/TidPl1r2aZVdl52HAxk
FVFk1GL0KHHlQLwT92LrlrA3HtbxTJN9bUiQZ5383SzfAgLL8H5PLRTKtdSwmFEO
0eCV26tqC+47ydeHTGY7EbemiKRG3IpzT/n2my5h9FLaow7hxzLs+kI1zfBMlpVd
Wod1ASz94lPYuEd80uOM2dIGwqzHQqzr4e/O+uA3OrLhDmKJIt9zeFDWmNlFA0kZ
CO4bJS4iUsGpvDJcCcSSi0YO4w/KBUypR+Z1N32oXDIt+XPuri3YG5t2tR0PzoKo
R3J0gxUS4o3wlJcR5AqYd394d1K2ahohA5OwH3hIt0aXUkJZO39nEtwlb1gABZfZ
4aPIibXCeT6fYaQ8ORZ5q0uF4PCVkdRLoZ2nzLW2uqQz3FGKInUn6qys+ujKPMzU
A1X/Lsg90raqz3P25AvJuv2+fqTDzlv3hjra2eNhL0a70gCe6DnBGptd/UNIqYgN
eN87oA4TqQPBqy42XfTznbsfMWBH44/Zuwyb7pf6IUy1+dZazNynAulJlJGbKZPO
kfW5pVf5GhRwmhGNyrq5weBaCnXpnzrCOXn/DCa+/jUlAVbuYlQPveis7zMFFRav
VIygBwYNwWUlZeLxfnVC+I6j25eU+lVE1jHIw6LWHbGP70TdASpbZRisYmFc6nWB
Q/BxWFpNkd8il1rI6F7J8uSM1/Woh9AXG7NUaLxfzCrzYdXcZF3SnZdIYrnKHPZ4
h0CYyI749NtztZfejxQtzEkBdq7E9qCuaZjquRQ6U/t7pSKMLAx1IMZuPOjLMzKg
oSDKV2ay6e55UnIQEcpIfbNOJjs25tvNj7GEn6DoRozF9MiF1lD4heppLZHyHlSx
q0Q3kD2onesE9dOXBaB1drdOssCbJZyk1+gOwtcIyYM+Wrw9shmcXDnric1dTVdN
bRyQGZe6w/6yJeEgZy0KNuyRPKvR7qtRUl+ly0iluHwo1uJSP8asqi4r04T+TiP0
B1aN/CNTOPt/UIWsYCJIJ1NWEsdzCDgF6YLw58F2kQ7l/K8orOeYJg9R3AuNaCiD
U9OGKpgg9Wltgzq+9mtNz+hTnf8BnQWBwuWMm+z/IzT1UfoJHdPlhSwSoYEmnV3W
BQagerZF506fOXuKFCIN0x2LpFGmsiPcUBUKJUmwJvpo6mPBOcmhuEbcMdW21mF/
hqLqDEL8qaxbTCrv0/9+lZ0wKsKUXwLqdse6KPXV58CpWoNIjMCez5FATYpMLhQn
zOaCPTvxfS8krgw7paBXD3zP6Kh13Yck6vwJjwq6tsYKH3ZA9ih+5sml/sfeaBMp
eAbpTrXyvzPqITRoBarb8576Zu1HgpCuOwIOlzHzNEJrTYQOYOWXJqt+HiBvpw2Z
he7JUoQOPOEBzPNdkSFxYhZi4oV2Mzxm4I/hBSJ2072naEVrfjT48erwa1+ArdtR
ZmjZF0PE0tRXniM6BchQGyrhdRiPALLA0fYtviZi/Pf3RO12cppTgx98l4WHiIN1
SriBAPfDqJwr3WKrXNRXN9K9M59jREznMNwH34GmgY1HK2V0UFwdpKzsyMGFOE7v
UrEobjwb9fGbN9BryR+5bI8Yas7TcM+IQvt3BiUxomX3+rgBmuzsHyB14hsP9PHI
g7ZfuFHYYhqygFVa38Ngdm9I3tKfJqp4eAoBcH9KJO3sXFmNtDfmwb9jIsBS4LSm
WBti0m/Le0jHAGZEBxYigSl8rNjPai6+DCGJFtY5WMF8x0ozdO77CqYtyoJCKOe+
KKabJ+liiAOL6gyjnEEk6tA1BwmFBuPfHvqJT1XrBd1MWg/UNEGLijLn8SDfycya
22g7ZjY5oAyVnE6SS+KQ4B5fl+ATYX+4sO25PR6c3F6CWH3l8RtpbJsU5eF7xghh
I+DZNBveb0qtBxZgvOLxYofZNXHiRuSXq4Ndup1nsq+kWOrZadqhxAoFTVvCzjbR
d2+H4x8joc8Tqql9WENeRDfNESWn6wHE0pZOs/yJ3KnhP+eW9OqetcIeBo7uIrfA
hOYVcg8+aDk0THRxZFd6fnkJ2Y4erXO9bN7NHMrpRk2Xy61e4HEkfPeGMXsCTyXA
4RT/OkjD2afmwywM9/lqSC8wBhXhpAX5SuUgpANjXuYiR9HNUDB5tUCneFi+CSg9
XD19m4U2FnhtJLfh8seZJrpSWRUdRR5y4qLckTyazNqM3v7K7PwljmXKIacRSOD7
hVj/ZqPR5J9iuwuhlW6SCX1wp7J9z/HSez/E6GNoO7E5w0nQCiyqc/LWXw4nNuZW
bEn2rRjpqduLLgD/p0LSBOmumVhUOkKZ9s9nZPd43VKuV8RP/PJSBjxzUTCTbKLJ
8ucez/iJQb6V10BAozxr6nyWdCFDZAr8ZfRpGD/4H88uF+u5Pt73kamsT/Smx0DT
JRlyfp7scFFWOVhUq9qc83l5WBbMeSuQq4ilpxO5WGD23nbf7R1/cwNtYd6uJiV+
RLfHpSe2DebCdDSteyTyLgdwCk/BhgewgkTeUTUz8g1R+a7neOXq1pU6/wTwKGQs
eVZGpjTwPFb56/YUzBtPfmOCSQB/ci3WuRIp5GmABzKT7is5Zs3OstpuR+ayaY2D
Amj+MDoYfetHV+fSe2w/E/xcsAK9EcWomgi3MY0/a2nU0f2T3H98fG+a78HMjmGZ
2Zk+W9B1tjwwLbz0rKmNnvfTg41UOnJ1h548RVGeO9mnq5065QmCtp6djGXXIDCz
5pSZGkSRiyHnLo+lHRoGt08YxFOZgOTgDPEYp7uGcA0CnMQD+wjFGKIBpNoPcD3g
PRcjAmkyrI0Xbb+KfGJvEz1AzXBQ6cpHIsyzDVXytTk9HVGL7StPB9mLc4SAx6JO
1GdZwzasfgcnd6K+XGhNGFdCW9UrtYjXNU+mntxoHG0uEzHtlywKRq7HB2KQ9BrH
h2YqBEJnU3IU4ap0WxLHKW8SlzG1W6zdBBYYvZQOhu2OVTeHmmz8rk15QeZfXQ6P
J0AeGzGMu7Yr3sM3GWFi8r8NIDz9hrvgt33boCvNQ9hTQ401r7DDgAvr0CdO96Ng
t0QtBLODUW0KQMi20maOf9vVQ3x3X4ybH0+FIA1mOGE/1q/1wPdfdcIcxa+jjjLp
+xVjeYnAD9Zz12WHVUIniJcxQK4Y8erxfYi+bcm5b50Z2FYHtYT0kNmWDPCOGvY6
r3ok47OKj+NpXsWUs/H+Ludm7Y710nOexEoCXm35V5/6E4vF6T9L9E2KHHQ90dyp
xa26I++lYnKeuoVT3O8zYS0qA2kmsnV97boEG73MTnQNzmOT4Mf8rj9lcEQfNc3h
t8RNoXJ03CvhLLCRN/4qYSoyaYWbp49xp9cBhzFqheeChs2tS+aGPO0bQ3t2Aysr
7J659hNwH83J1H9k0S+BA9oz8IuLwE4o5CtWWcOn6mVvqOZtQ0C/V0P8q5M1cA5j
GQ4e4xTIFNPIUs8bWvrMO3I8mpRm6DJvH25NNMQOW5MygsIEzunHzEhJ+BujXMra
fbhiAo3KXUIp3lnkIiZLL9OdC2rEEzEreVa0jTAYBbiY/EEaxLLhRx59nS9nKowd
fiV/MIlUynnCflXyfvzcsv+or7ajlfrxMaFx26AIA8NtTw69aXmr93DfUIVz94Ti
LjKVrtfqqEJj9vCPGhymEV+ycuwS/UoGM69o3nzACX7wGcLeyG0FSDvisHQID+1q
RbdxYFXbjPCgHW5Ym+eeZ15PJx1MrffplPkr+dw3DckUJLvc3CY6nkWq08qc0iEN
XWhpPEPvukg+R9CrmiOBKCTLVGeV2dYpF1kKxEx0t2H4mfNhYf3ngyd11H0yymoM
SH1zfcCTB/a/hgHZya8knn/u68CDK/3NCv7oiGlC16LeCtBrbpVgmPx97A8IkifG
ZzxHAPYAg/qDR0cWka21yJbMj8mqvfzTyNhJpmxqpAv3C2xlITpZZs3C/BpY5B3K
EDhzEM1GFKw/esk4bVCPu8Mpkoe5Zf9JpWcaHhHVE/ankam+Luew6tkw32BZUNHo
8rv70bOVn2g32HJ0OqwhqbHE+nmuoqTFMgwy0fuFzooxSg2xl+NGwhUsxylzLZ4r
IzU/mGDYIJ5AJsYp/v4ZjJk9Xr1tsAJKfPozFFiDaoWoQher9lJy/VIEu8pwE5Fj
5AZfJ8iadL+2Rb0RwRz6pqG2znoaqZNCk+nldoeFDbvk+6gjajIT02gHuV0CG2Bs
IyY6kgbHj7sd7pIr3Zkj93Ep3MejSwSvXnkx4c8YdMt5ENk7NyBoXSwNZcC3EiSV
fDeSpxOKUnwwIoR/A6Nqq9WGio2eyfexBJcJLNJstoJYeBy9G/QCYAoaqc/zaG2E
FvxWifRN1154fDIcYTNCyribJwvARqgOjvza6FTKEZ/0NPxJAWrhUg1BRD1OpdZ5
BcJk8uihKIuEFChJAxbrbOjlW5v1DEzmoYxtQgufyy1+ObgzcMaqPtkY0nZws8pw
2954NeQ7/FMLswPeQ+5xkkovJtPKJXxeqglBq89RCL0b+szkj0UDwV8sjmPGewyE
35tJSJFrgIoSZoJEVe2Nl65XYEqdfBZmQNwE1oFCZux5TYmLUwHV5omE0o8oLfcf
qMgpcauRz7dFCpg+qRbnnlKDz9oHP+bxeCpA9gqUxPNiVM7VBnQsfjaC8+rAD7G8
MHnYlt9k+mKEFcimNb0OR7543cnwxFb3Xe8xt+rSHlBkgFPpI8ZTwP8ztmzAp4Hm
dTFnEL9Welw/owjcQRnpVJ4kHQd29w/KhunRZAZ6134/Ft2mUFOaoqIpUAOlRnF2
7UPIxcoRc73Kin0PtUSkK7UbhhfCXWUK/Q9uljIRqQiq+GO+B7UmfwEA0rVub6r/
nyGiMBe/5173m47GReGiqfdVLfVRV+PE+KY8QbR9PorPDRQcH+Y2N03CoSVHQZrm
WC9LzWaOuu3L1xx2MS2wYjxhfDp1ZhbTf4zNhNnjBMPc4M4jTDgwyfgTNxXFHmXq
RMPXEJDS+magG6AldEVJHVD5cclDX1HHMSad3h7ZsCdNsDt/qs8cK41FeEKNftwt
qE3/yGEON721hpkrxZZd3hSdaoOOo18NUfjfPUCAliwTLIMPkb+mm4S5fCouptp0
bPDAiHw2I3Nq7ONTs2PBk+whWfbsbX30YjVL/yS9w3JxeHH1mZpA4U+yO2C42oTz
UrOv0kOug0S7sZ298o0+xyXM4rryPl2C5xuSbvskjV0XTm+7ZtSus+DCNUNd1r0R
bibtH+8sXyqKS5rPtwZ5XgPohl/uVcloL/moE2ESCJ4lW9dF03E/PP9ER4+OHh/9
bNzgjOHaQLXQN+tCift/B75LFjHnDvL00UZaWS0yu+yjLUtQjQZYvAXKAGXpSjqy
VMgc/HMRlp6zn5nG2jacQ9HRQ/psq46Q0erwM0NJg/AsOssCM17+lYPsiqec50Lf
7+4RIDJcjJ/9A7N6GG/C4G86keh4pEKnCe+G8oFtx9Im9OkUDYuzmUY1+ad0PFpm
yd3YoeVxNcFJG2eLw+8x6GIL0XMI/Sx077J/e2Hnrn/Y5WFqCYQzvxHaZ44Wh7oC
L1mExvhuP47R5Rny4twPJGO8KSkS5q0NxwCfJFzrnVygbxziJyTAFLkdncq/c2Md
3nd9gbSFhEaR7nQOtItjcsz1CDvCtC2b5VdbJFL+djm+7macMMSqotInBmLnRS5Z
zlRs41q1JOC5drWTczLSTAKKVlyqJY6S6C7bBXHgL9/mwHgqdQhwgomBnZxSR4pE
1BRpccqm4tdVVxK5wTZTjwA4j63dIxATuACU7pR3sX7jscLvAsyEAmiLnxE3vq1N
s9bUyehdNcAGoi7RaDPHQNrotMZ9ACx3DiO4Vf+bCYusQlXhqCzv2qy8UBKyt/aG
sDp62G8tSwjlOCv9pn6zPTAshJhcT9RFlbrIAnPQxBM3M4wkoGtoS4srw709mefA
B6Xj2y9PrhY00MrSYn5XPZzj3lzDHzK9UJ8tjFkrWY9+XJt6pnL3np6T5OjfWA9l
WlCfQrZmck1hHsBJwuQBcm7qZZX8EfPQpk8eA8pHIyZmiSk//baZikJunq3MQ+8Q
VtUadwB6doAIaTFah0aiZamPgHHAEOPFrxaiBJ46+h4n62wYx7IZqcTlNoUvRX3P
4nXUuqdCYX95wPjgfn5DRYHc9GoskfGkxxMWTQkEZPT1g8hp2FX7JIOBuXAr+PqO
cQ+6ZSR1WQ4CGD6LYDRXbDdz2v4miwBDgoWudNiWwDrkMVY5ze7lZ6iQKJFdT7k2
neccp9vAotE3EkBaWi60glv0TEc/R5IWPwfPJ90oESNlTaXjMGB8sTPBLg7RWcGX
xN/rBEAk0k4x+rvgec5S6kFSTLn+ek8CmaEd2FXC+fWKgraHqHrqdDYPrHoS0RF2
hip+Yq4WXpc5maDUH32sDDL+hZHEgySfMKQxpfIGaakj2z2EixEfQHCjjOh2j3Pz
pGRrW1DQMKJTR3fxsBcavzX5pnB5b8X1Gvi+A0SaUlPo6q17GP2jxtz7HMrYQvJm
OrZAuNy+Cl3WXqACMEZhxid2MdiR5v3CwSpZOAlbyFkxPeh79GexTC3JVgTi1wmz
n2E4ObIBGc/myL3fGtTDt8xiUG2fqo3ZWGYeWvPSOYvf4IsRsQdfFrKvhdOzY9uD
GXqqJEW13ZwHQrGLWj+rtd+TtFpkfRw2cQMaPn7gAqcykKRTuunmfw3v6fSMy6WP
T0yu/6EOomlrHGDAaXmTjBLmHAzRoWv+laJsmsXI+pYAvoDhG8rY+GYxn0FLCpRg
IO9UW7OtD6rJegYHn7xbgrXun/AR2JKu/zLO7Y9umVOhhGTWie+FsagnKkMlriPN
iReYoqoUxEzzrhKflyEErNZYLVMoJkOeDpBmkqmhVecMw0djA11Y/Xtrx2WFnVGE
3P9IQClTcV4FLnTIvmr+VTLqxIWfR8mZlZU9VhUy8zoTFaqISe/JYmqNjdO1xcXO
/uMEszaTlwVqrXRLOAlNpO5IgYvr23yuzm+P9YwTbHp2RWDfIVnO1UhAwjVCp70J
EHPH0EdNkgQs5+zZRwU/Mq9xIpiRukgDQo5PEdh0R3O8Q8MEdNX4l26pOeNR7jnT
0YsrY2ZBzuFOy0QXNsfNpeJ08GmfpntrFmER6ref75+wHN/Kdkf1H0jtupP8iU+A
CyrgBCNYgOoQlqQpYM6Yf76r1bN3S1OgMtJ1p+nVLiZTQZjKf8bxUpQfWqF6h9JZ
SaLIEQQVQYVJzuJJW+lfYAGVvOHBmST6ntZU9PLsiUQru8pyvwPXW/CMYx7nBQ1N
Ulb0KlXc0jWGjknK8P1TuXgp2RJOlKPxhwWq5vsVLl1J25RFAeVl3rsNojOmBiOk
iavovcLD/KgUtQAne1YKK65oYN4/H4+cZI2RGh9ioFsxR8LNOvqtObvTzfvjCZnc
ymlZpZk4x4g2g1t9dWz+6v5l/oGyA5YnQoj0aEFzn4Je4kruQyPSkW/aZfh74bKM
seXduynTMApSlNydcY8GW4Y5qK63aDTlnVEX1zNgljy7OYxNW2L7N3IMLiYU48At
zDxvRqbkLpr4aiwaL54gz1wRyixOGt33wm1LlMT5R1LyBzO+1EEcGn52x2+0SDAk
d3p64XxiCjqF3pxSrh5KfwQ8i5wm63nEAHyW23szws+Gv2PI5AS7FPBsgMGdsuor
OA5JYzpKAh4q56KrIEFbmxYxhKJZl1F2stzpQg+TgAd9nPCt65/2D/ZpXdEbMHZq
S8rsGVxx1+J4WAc1iyVr+ms5DVexW6aU9414jWop0bSzXN6/YpXq1koBP37O893i
E69aEmG8QQoHZZSwzZ4kEpOZ7E9dlvgWkKgqn8pe4tX7DGfxdLjCD4Jk2j0pXWAg
9vYVO+lf5LtcX0DAI6ya4HBJH9p0mBDPG3qmV+A/b3FB/aBjDyS9p/I2hlPYwE0A
gq0g6PAy54y/M2VC+oJpy56Cyx76BryVM7c7vwmvY2UNaMaAUrDvWNjEjN88669K
tN1hGnZg1t0b95pobWYh9d2okQCCiWgvZALpqL+ys9/jROJu83vMSYQHKZy5tsGS
rG0WMi65+8W5nH5EuGsC6rd4vu6uw77LSrLzk9TP2ljjah7w06baM/d7Y0Xr60Cp
WzI0l4x6rTH9KrsN1ZFTzYE88OKLkKPit+GuURxVwkZ/gr0APmSynIVJcvoZpo9o
rHyNZNioMEds7T2NfdDt9RoETy9pU1mN216o3G4/iJb4u4JgMM869q9LzdNwrrL8
R/Mj7a3ZxI4icBI5AMgAdwroAv+dWAqmISFgdVWGtgYaSi3i59Of++EDHpBN7c+q
vBvP3gR+upt+snmziRkNykg2e/zSNsZcPAfM79QormFM1eOp7mfkTRQoRrEMIaMS
FGgmWVwESAy2li0d/Eu/f6XOX4o83eHZUUKTnJg7ueHRRu8Dez9nBWe1YJzAQICB
t4YCFAXYoaQVU5kuGjygrvFM58JEt5ONkXtd76kyY8x2iGeDgX1dtxt4YrtAZlnm
hMYp/JpKVRaGLEvMEnlREFT16vDmJfrA6a42B3cja6/h57fv3pZXAoRZ8pV2qvhn
XQs+HrzJqoZPBdB1u3oGoRKGVWD4IYIcn+yF4bK/9oUWwT+rsRcG/a4YsLZpCM1j
nxv4O6w4csY+FIeq597dVDgmWX+xG4PmZCaQ0vVeVKrfUGG1kmVhx/Ax8BXc5H4V
rEXk2z0Z+FIxDjHMDjSJbsHFlEfp9dXcINmQnDQUWheRL1AvY7z6nKsrBFkUWs1U
1jvxpv2dOH64BJl85uCk+17BWYMUnoRkrFkrXOmZSRET9z/8GHwmCp4ESfoAbe7D
7bZkJB9LCo5SS5rPgWX/MQqxR17Y5L7TYkNloe1x0pUxQw8Iyo1zw8OhHJC94cr8
peKaZzjuzm0RxQzMSiEN9ENOXgkaN4F0lw8aMSihibx0d1OhMNy9u96W2ZRweXTU
BRi2LHRTTTs5+cj/QQM5foHYGdClDSXAN57fkZnToSB3wY4i3kSVy4UPW8abJ8Q2
DXJyqdZ2xt21fHuP8PR6cKmOC2kYL3kGLChlNm6qBK8DBVcZJak3GYaB78ppCHwW
bY8OdUhNOA+CrIn7Zvycz0oMUpwkVZw3A31JZSkVsVhqXUKhZzPAtXVQjubN/7cq
0eQuJRIyLBnjepKSsmHBqEDBC0/Qv8Xk+9eWkExvJ8UqvkKrrD3TnL0TnSASlTWo
3Gwcwoo3lmzyXD67XpqJDtxHvM38g1zbBXEhMs3kagyd4iqUuJBqjG3N9fG/6lEu
bELFa2p/ezkGVLgGuue4LRwH7CaHNULTEP6R1Hn9eoiaZDGjrjRa+E7Z1KOo44l7
jq4qReKcnIMOf+pdepscBJOvmmv2hpsrAmiD1YRBQ3+8SB1H+ZguAyLJUsQy4pI1
Nr4AdJLTad/WU9z4ibfC/rn0zi5IRKP8PNDzP8JopBNotvV7z+28b6/ySwsz+SMM
xILMeXDoqzpIxwj7gtEd9iqTb+5ebZ+Bi43ZByFxtjyKQ/t9Tw8LYiHebHNRX9ps
GBxugItwlGgFrPAWb8oqp33iyrp/+vJLk5k3U+0RFfeiSG3ZIN9dz2XO6AVainBE
NY6VEDxgr4M8ZDby3vS8kasJvBNwzxjnRJepJOS8oeprBdbI1yyDYnJSKXgIT1ZT
HLNc3MW8qoQ2i3FRfKZ9yBksvWGJozPaQGp1ZdMUWMUV5EK6DLjI9PN7lyHjfeOz
eI+BhEnu9y0QkIRZJSCAA57NPuQvn1DoqruNEMEE6P2HJXW5Vd8FZbffL/e1b0rA
fa43Ip0KOesd9sCIMHhLLQqYJ9OI8HxyZ6fOGd0d6LIJyFut27IrhpSZ4EEJVKt4
P1uA4jZz9z/U5q48RynElULwh1RjPT/Irx7NCK1Y+rt2n0nRZVglFlZPu8Ez2C/f
Til6+m0PN1oo/yVVJ3nrKE+5bvSdHQQFsYdXVZnFSobLpik0HXjiFJwvsai+wJcw
5jv3fJBk39dyVdpMC2TpxbIcAt4XKuMEu02rjR3Jd6+ZdvSAP+B4+bjywLOBwFsY
nwdUbzeyXpFWwfENjzl8DUjMao/BB1Nb7jsCAXH65CLM8PFQC52rqf0X1/yHojg4
29p3cMt4uO2jbn8wHMHBdpbqmuxH3F8fbdq4+vemolLoomBekJrEt0KaitiAIcAd
eSh7kIF1X4K+/KWjsMvKMmtaveZop7TjUcm8gX599rvK8VxdYTm9pQ4pQdY7fkT7
a67x4bjWqngM9oPwXEvM+1iqM8lr2wv1Ivzy7nygQalbf7u9tDcbQqiXzXpAOgjp
9J8pRznnuc6X5i5n7dMhwwWrYNaB5BZqumblkntNfjjB7eLotiu+EGAs8YkNAOm+
qzgKzGivkF7IqpwdDqLDNEY55DAJIV+bizYGOfDBYz5TXedQfB+uolsU95tGaGKi
pbiKoHcKwP/IYvXIA9FgzhUDoNlrzR2L8R6DEiVR7upgPr0kua6+VGjpxq/vDuD2
jz/w+o7OWxPkzPlCKYyGX8nBoikmBnCx3Jqj7wmnPgiqQkURzIutYS5s88A/Em0E
TyCcClwhxiwXzIrvuUyFxNDVEqSjFP69iy0EkNZ5rttYyJcKQP7v5C18DR+E/9i7
JzFRizX3ylH67U0FgS4DzXEjTaH2qNdM3djR2YguMyKPG75ywoKunGpOkJ2UwuTv
fLCBi8rC72xks0asasjYxuK5nJPf3D+BLD69Gp3Drru1DfNVhuelToagbHh2F5ZI
hbLC490ZdYo6IAmPmLbrMTK0NUBmuIYKnci+JZrc7R84keGLgd8Rir3LXiNIqVJB
p14eQ2xaIFse01CjqIfOj8APwcPx9ANTg1gf9waOjsDkI8R923TuU8iHlJ8kuAzJ
OXql83b4xXaxVJ3LuVmpqncqtBMBVoAYK732zUdcEfuAMJr2uGFBIMqUzPw9dNST
7Y34j+tV4kO1tIwltnYJetJITWEsp5zs0qcx2BTd9H9z+xqMzRarDme07CwVp1vd
5H1O1YLHQx/HxLpa37P38Mlrf/Pt0DLMSChKDDe4wgd6roXRgJIDufGzglLmVVFL
3YbiTxQJslmU9xSL40+Vc35FO3oEP+fdR5O0oSAs7tevmtCeQfjh7IHSxZHM9Fo6
cDCXyP/nBsTgUf27p82khparxEyWb12k/88lk4wG7fePVQQkkwclmeVg2QtXt9QW
oUDEs42HqU6q8G9HgGT4MnwAadG3RxzZLxk5L2bbwOLIVj3+gVCLrmw2WD5lkCnQ
2Xc/B5CaaIKmqqojoBZPKTCvbXURdsg5gdjU4wLmmlXYjLL4TW2dJs8LRwZefv01
1c58eSQhcGLLD5RTSOkvnuElImjIPNbjIWhctrETfhCxFlSTmUA/uSK9JrTI8fxi
2EnLW4CoTm/R0E0RsSDP7qSFxxBBka7bN41ch0lVBRFVV2a1ZCbclLbsjxOlHHVJ
Xn5Rr8yfIQANwbO/bswpoBy5EEGQEzUPhG9GbpmsKT7awa48Yn08Vn3vTMcI7FYc
6M03rO/ukapSVgTDZ9TUkZlQe8nLg4sg6vxpfCeXPAjUMYROSJIU/EKvRUAZI3og
fIYKPVS707OE+QaWGVsCNNhJVmJzJA9qfwpAXa/hO65WhnfmIqqIzUg24osCMUFM
suPG89x/ZwcphIqNoKwm+SS4rQRhOOWjjqnv4ySbqCxu+n6FfZHgGEzQlPm3orTp
DAWGz9KvPvDdpNY4RHHbdtHJ1OJzMfyMJ/u0Lg12Tpy+iS1ODmsRG1WAE7IHgjXj
+pLzD4sT5CpEoEexyMjL6N/qsVBiQsKX0WnedJhahcztZpXt4mGkrl38M8R3nHsI
JDT6hoqmEwMD0H6jgbLKBVl2BZ+g5X/wKtE+whF8EEsUGt3QwrVMLoHoxkIKYlto
vwGWA0laFpzXKCwVPeGVCtf5L4koABMJs0xmEbtIe15OpIkAXZQlr0u/eEHG6AtJ
vKmMGPhN8QnrqpEZf+/BlbZQaA5bH0w6VIj/6hzfBklvbb80ilG7f1kYJoAg6Hwo
oIJBoJO3+mACiE3WhUQOsSrG1bvOlMqd6K28HJllKjAAlfurikFdE+8QTR8OSNLq
IkK7qFHc8/VE1GRKYopsvgA0ZUEq5tM0gpGFvsA+HGoOHXxZYEq8/fobRialpm3B
UQxTEuBN/htTOCenOVE6yojVfI5eAsw2AGwjjq9c5I1XsmQO4Ps8V8MTaJv9JV6l
dJUDpRgGERRpI8umt2WbibwS007Rb24R9L7isT2eFfLBruMNg7EsrCWIERS+iEE3
ce2MMemus+6dd64FpqOqIMLsp2MqpxelBYxNlgaLcRTMFGSZMH4bVLedXPasgSTA
ka/M6kh6OCc3R8pcId0IMoCGs5cflIACjs9TyoAl1unCXGSSYJHBBaMVTSJoHmZS
ldttyWRuLBM3z/bU7qM4wXt2nhXgQmEyv2cxO/KIZfVwEZqMHYLPCt0g/f24ysqh
7JSFEK/afjLejT9USVM9jEADh0WgnDGLufr2qPRKu5EvYXg4+xjX5mzeZ4pS9DYl
DZ54yZPuLAKmllKuWFrWzy8Kxg1hoiz2wFVBaOxUWCQZAGjdItyPzvy2sBvzCj4j
aXUX68FzR+lgGkt7Ua9R78HdJN3wjz1KR/zin1mtUosSg6EIDlWoXC/O/5TK+wAd
PWK/Gibzewlvir8VBFyrpF//zxryb4BulxYsBktyDbVfefqnVm4rjYiAZhYaWqMl
uTXpARv8Y3EGyVdQ8Ufj88AuMa1KZVk011P/MEQQiN2qwKY9kWkg6GAwWscSII/h
dqhEJVYiupz9kGKe8cxC7F0PF1h3TlLqWr0d0IzQ2FZOL8nAEr13yUI/0inCUlJs
pDrOUmPXLq5PUu3IQ3dTYAqQ2ovVYX1vEqMtKHmlaM/HdWN17Dmz+1gd/msIUr9E
cES0xdYFbDC1n7xx28/D4JZXagBUaIpAigP5zA/p1Fg07mtSiBZOuyoTSVqkh5HM
M5eF9kuryuXqxjepXtkc3xAL49UPkVpPigkh8hYR4C58cuDUIgFzqOEGuqJN72U9
nsrMVA9/6XG6vlMUb6jEkan+ITFTMM69ZwTzj/sUOfZkodAjGAAY8hDlq/0rBkz+
5ML2Sq/mmBsnRTwbInpAL2nIbCpds63fftqRXJRaXMHQqFAbhC9wwIUiyrpaRVls
wUKBmXYAPxCWccqv0n4VCnoMOQyYThoGuCg9UKsATN0Nus2xQY6sUUHgpeqYfga0
71qRjPqBccY/hOGdeFacbcovmCwEpx7i+LSpMCcH3mjkJlMwB0qZwgmpgxNUD4nV
WGAVsd8A2oDJ3SvNC5Pt9i1vBG3Tn+wEKrKXjlQeM3IWV584VeU3yN+JdbLQ8SjE
xWKDafrnPu+a666u4thF6B3rpw+1xnJ7ajVl3YZa4hAa6xXeqDmZ/QmXIZ4YrrIO
hd/EVzYwmhbx9EaFY03NppYCMkMsnCC/g8dLmfhDkhLX5cvywwO1pdGRYqbzJ7/l
k2kGod48SVk3IAkKs7HhDeWSj48Prnb5s8dU+3vxtOudqJxNTswWFiSnuWWfHSVN
W8KK25wI3Eh9O78I4yQIX6DeGpEwb1YA/FK2A66qVN7ke35c/2FgCc2vejm7qm9u
DVNJ8jxtlYX3zU/6rMTJkhSMV4Wb/7vz/idN/Ql11103X1i+hyeGkKPKCE/YWHhP
iBrjVCs3WDXYDIkbspgwO341wUT5Of2TgyheVhysmpNpsWsunY6N8RkA1I1PyaFQ
cxpzqUtZktJph6WTm9Wv50h963FL5gcCjRdAKdVyLBpvOiPPJiuP1aOTDbppuWKm
Eqnw1b62mLnzqS1jyqqtMIrKdMK/rvOcAIxSMLK/j8MHgaRElzSUMX5Q+czVU33/
eIWERIEazXLhS5w8cDEACARkBc/UMljyfYO3h55GDQ2Vz2cBAQjKaomKuWg6ydm0
uprjhHFYUuZjaBpJheVic7bN/8Mn6ZKKgwaTOxtqm+dUQrtMnz6Xfms1qWaeNC/M
w+MsacYKlKqhynFv7O5voSTx5hTKdKADMvBITNmvJfkrrdCgyn8Uo9R8MHjMvWFu
kWS2SEV3xDqgp11dJeWXxz94PQpNvRkC2xujhWmkib9WyyTijogQiRkdc5UO6Hph
4mpzmWY3hTi7w7eanpRBF34Z4L5NgZoFs6u9xRSV6i+qY9kPVpsn/EcpBjjpJ3WO
YjkQvGwXv129Gzixwib26fI9pGFdjBPEK9tKNhpClWo4AgURVMbS4PsbLiAHIJkm
YVbVxgFFXlaxY6ihR1pSGFZZvNG+CnKul62APo83lwbEtCdhibzaX0iN9HPtWQjN
BNNmpIOIGh4fRdh6rDpRJ+lqXG9lISQf8/VXOJslNhU+qX9vniOevw2O2PQdh1LD
6E3JaFfy6LhMx/VdXPuqrumxozRvlGU/vH2rZrAn0Vf14CjCshcKXkRCqY40pgfa
vVKWL4IHzI96oRhYh8WQNkJ8UYJSAPjgpif4RJkQF3tSGE/W+1BOYUmzdhqjjwJL
teRt9wci/dqh7rPmo4m9u+Tj+BC5fueovkOtbQ7FxpwAj7lBN7Ih2dWURRyHvop8
bQagNyWuSnmWiwThmUdJsYLAHx0j3Q0fGr5s8BeJ/9IcltxWnDjskC9tPdPcnx0Y
ylr2hFYb0zh+W7dob9TlmsgPLsZ2zISR2X0Hs6W9hbjw0Lt6J8FWd/OmIAiCJM4v
Buhrw6Pi5n7eH8srqahFTODVCZgTDAv2neThPVeTOMlrPj8wbeCZfyO6Xr2mT23R
N5jZL7iSmBAS+K1i9+W6dmfvXNPY4OvyKsHqmZRc3AjInxJLo95tvRFu8+XXezy0
dzpPilu8DjiwPBjYkum6Du4MQfs69WPbgwAJYW9eLQKRw+TiQvwalex7pt5Cb3BP
ip4UJTBjigDGuKc5u2kkdn/zLpimsaYk8jDRseGae9GCZW5+nClun9rRkkkdqTCl
cUPRTNRDPAi/+GN78KW6aBUHJSIkNly7CaD1QRnR8zLn6x1XpS3IOoDZJaDYXWln
Jd3vwmQLMm9NJpU5bVkw1NzdUucBQWmL2cq5TpxCVTfRS8wC0AurYpuJV1i2iN+H
lAWn9pfl1vmYSmSP39ZZwqXFg0RHnYJ705742i64PT1Ib2omxuzLlOC5iAbnyJl+
BIQQpTg08ER43A1qF5z0PnMTIE9Lq72464vdoqb9Dr9UKWdKkwTrzNtjXjoJNJWj
BxupJ8uQ/vQKSdRK6Be05N9ydhBD+6NtNcBXYnUoebbSjXFnQE+45NUC7g8Ob1MZ
IXgBfrqUjBVl9Q31EFmSkXMCCVM7iTlNNOv69DQnKeRUp7otxeKe7U6eNj5Qj8Vg
usjwkWgiJ57DZtWdwERQCOtPECHFq0OD9uNHOnlTk9g9Jg6EeqxNT8rdqKjCDKSI
FnKQQ3GN96ibGorRpsFLSerIWuAlZPnt+5jsVqiweXgRQkace+5v5ixMx5BK2YHe
sIgSdSL/8+a9co6VwYDGugXztMb4JrCpaMO1O9XRb0xRHcfNnG79b1U3J9d3cMma
RDJV1j6Kv36igEZ9jF0UfVJu/EDDMhJF2ffIWJta9PefyuRUG4F8tPbTn89RddQ1
Hix/vv+pJBsbFUwIVucoo+CgTMQhS1FUzu5BSzFQjOc8wSN1xm8/AT92K/3czIJO
JDWuUGffAKhdv3ZIbjPMbKHdeIGddyzhOd2t+QNAUF+5xDOQU43YemXY+lHEbZV/
gvEtYf4/D6tZApbXwqhKI7PwTuzuANTeER0lTWCWCwlOwBaNug+TaPlC3oVfBMix
0VJf72MK5BIFP1q9rvlmj6xRLC2RRPquixUhWiu3X+tdxa+PsnMVxJbBKOrr5J27
IRv0HgEeIusR/PFrtrFepTey5i9iu8Hj77Wn+Fwnwf7eL9eIaLsq5WUl0jYRwPTG
11Z3U8Z12w0v/nWsHu64dixc6e1vg7aAMIXU66YnyqyDCzx3N36A6SzbBUzQ28xN
aXEvgWMZ67Ge3+DkOacdbDPH8QB8c7qQjse0uch81z5QPH4y+cQyI8a8Nb8p/RS7
uDOKd7IZersn/n7NdU6LIJtQB89EUYEDWp7ap4dkz965Nkl3Wzz+aqIBodsHUYF0
iP1IiR0wNBjMHxe05x2SqGpIQ4+lF54OZp020aj9QzFR08OROpgZZlccJ5iSTxmP
qgrfGbwYp541jqjiAn7BBnv2ZI5/qix6UIIEXLY3Fhp6jmJcKQYATh1u4trzXK+E
OY+Xu1UbE0x81HZhJ3dZW7UOkUxQx02d/qbyOqZPi+U0hh2Fnz0YFx1OhB0Isevu
8R4M0CDV8xLYPxDNi28cqQdnlCWlx57K/FIUsEyHnExoSQwO0OlsK8JtTiaYtXDs
2fqoxoUf7MuNUfL9/1J9xuN0jsyJ+ZH9TtPXDHaXuqoqU0tR+LBHwJIsKwDaaXL4
OKeuoIDCF1z91l94UfNbyQRRosn9EVX3AkBTgDHyDimpHDZqs2AOQ+ORDhu/zwwM
jcGjQZ/on9wEyl7VZTmqlj4UTR/DwR3M7leqO1bJli8106tgV5lMyZEM24qoWdY0
GO8XqOU3xxNTRcBcD10R8/4OheHFqgnd0nSZ8MMmC1kXUERkZRw5ZkwU0ARYYLbV
6jB9faTv6WIMgJ9cf5LZ/rTO0Qfk2hu9Jvz2D7W6o8qh8LAF0WCHUcL/JgPmdjcm
J8IaiCrjl4rkldYb4VI92TBW0dTAKBME47JCWOerxd2UQ5a5nIbWzzfJld9v2qig
RAZ+yFV+DflXXC0nEHsmoo6wXuEYBemd/v/hCZ2exPvj0Fm9bFOxqO5uDGMUkwc6
Zk0xaJa3lZsIt2krmuJTT32ZrDgEGFOLQLfSklHhglWzhu0UuM23GvNDn897UGiO
dGPtgdjwCBYj/PWCbFDa8udoQQyzg6C/8iNErmfmq5jE3qxMhF35z49mTi1hzs3J
9+DdU45H9NbvLhJMTj+0tLLi6JH8DB/y23jWIK12XU0IV1dmGxV9T2wwUps7tzsk
nzAD0mA1zIu5SUzNogS9/JyolGyVj2kpwLgRTMym6wfJkS53J1h/OhMoHM8xlXNm
oIgW3QgSOVN63qxKVMha1c7vHnqNOwBMObgW1mdtTWYKH8OqmZst3H2zkbgbb+NB
a2DmxbHz5ZEgMXWc7QL1EhzfTxdOjvmmUYV6EKuTUxL31kkl7f03vSvAQTUicG7U
6bQ9kjEuJnD8xdv38+Lz7IpW/msVMmCBWsuIbO050K3S2EkIhJ4SkB40APH5HKJe
0beWsJS0Smg6LWZv92048uwbRnZRTjsnQNRMZjFInU8nvtWOLEFs3S2uNAux/1Mv
8z0vg7jiEeKl0Jrt6r3ickLI+k2IbU41gvdZH7vOjwyMgDrGonhRCDXgnZV5sNJA
OU8cm9zTWivC9t59y1uvynuN8SDK5BHmJojBp6QBAMu2MSyzq8rMj2MckU83IkRg
bWWdZ4jBGCXch3hWkZ3+rSbPL4t+NenYufJICjbB3kBYcb2s8UOyn8Tnb16rHT8m
/BHhDrZvR7A7n+Twqcuph5slRvVo7bPr3/+I0WaYsIql/Rcg1XrumjpRX6389CaN
sxHHJmXRIWKX0M2p27acij7oYQJYRONv12hzDPRVKQC2EavbzlWRqWc5g5/Ge+CE
kIQ7TPU8NPj56ry3L38gS/4xV6Wyf6BMOdSkTPBefg+AFgoKgDd7KK5/O16hYN/V
f/Hh08nAsOd9M/fchrgVI7FxYDISzZycN2J1j39e370HKICk5hzAUVDmyV35KTz6
ollXj21K9fCrNQdh+xZaG4hVRYETuhnis5lyU/jNtcBIM6C9e3w9Qc27RJwzX/bv
a6sxiHBqKpaG8AsqVPUnTD4AS3wNf68gbkP158IsBmZeIub/dUuvCYKB47Gz4Qkw
nYYxeLHQTf0+z8OIVvpT2E91OSA1vy5VEX7oLSjkkHibiCQyv/VwRs5RHzHUysID
FmX9ojlVu7Z1gNyDjuOWOt1tsyosB7dPqZh/PLgJogtLuZaqHVzgjxzs/g26cJZ0
YxlVmpdi0uZipunj6pQczxUV5lWk7YXH9jYH3+inpFkJkc79mF0P89VmpNhL/UnK
SPvlZPf15m1aJMUdZFhUY2QYjdkTbKTHJvT2TO0C74UNWLoqRZ28IHqygsbC12+Y
3kw0QWKKtslv17pJkwjfajfX1a/OMVP8BlxofLkgkLpl58X/ORtAqsoeOvJXr0WF
U7t9zU7ZZG7AIIknSVKXLEuv87bFe4UnpJUQ/MppguaLe7rgqGJJOWSqDkH3ArrZ
niAXIr7LpEPnSEnw33G+4LPVGXzCG4/Nhwi8ErJNYgOftX5b1VjP/+BC3Zpiff0v
E4GMCz/Vqo4b1U3+ZEdteCaVufBoS7lDPh4NprTJ2XqSx6VFl9LAiWLVI4bqYxgO
o6kBjX1huEar/rTpjRQ24rLpMTl4LMf66BPDe6hOj+PYPosPc/z2ZE+hAuwDO+rv
Ay6+RfyeXRa2+svfBacwPd9cmVYhhH1Wg/+xPCesiIWwTBSjmwdK1JTiHt5GYHWo
OtQt0JgUbdeJiHy55SvnD07q83ll3Lm+aCfZ+8Q/oYwkHY83+RktWsjjCU71CTgX
i2CVV2fa1+Cb4IVA+6x4dUgkpuh8iSH4cfhbaMr9ob71+xphY7O7x7o4mLRr3cJf
XLnmdmVzYiMSdGa7r5imHAnDfThYOFnFnMgfMJw4NZdYOh/AyUfWKfUf1KbKESmc
VcACYA5juKRDix67ox84WASrzGiBSRjnxNTgehCD6OaYcp5duMhaIN7Y0vki8vBe
03WfpnJLUoW0mIsi3HDOGuTNtrYmqo6F4XixSk6WrfTFr6MO9mCvae0HN6t8P7xQ
J1Ey6xcseskncVyaVYgvJOFghe4+K4SQvyka3TArwQi3NrvK1LCxnZ1aN41nx94k
23WvfeYvPgLGMgwHkA8/Cx4RWqxYqjEVJX/WB/VL90zygTOGZrqfLBdTKvGLiq+x
gO4h72judX0UoKlSXlMcFg/87b0jkLDXr+Z7hgvpzXxiZXt9jeD/GQF+LVpPhzsB
D74bigqz3uz/ZGkfx+e6KILNNuQm7Ki5eSSRS70LrxvtQpxADXILil/ZY4MGz6dP
KjqFtrExYbHtE9FO5qk80MxAa6Jet/17K6GikV6e4F2u3UTJY2gLIEl2E99/OZ7M
NETO4LDbU/Q3zXzjmHk9mcSUZVgarSmYrblDaBSNhRyZDzYrvA5DmZKsTsi+zEFU
ACW+yQ8R2G14KzgkKqFnhmb5fCW0Qk+JVM/1VvV9O4NEUmNinisIqScVG8lnvb4F
bMDBHGR+XR/f8zfFJSCscR+DNqQM93Rl0rGTnbjEvFqG5t5OqqNSOrKT8RLAUeW4
X9OSLZMZaM84nsVXMyxpI8tDDibwOdePP00dQ8/j3SeyuSnVWAEp7zFHMG52PQUZ
2eV7Dojc/+AHPhGHMmN0ajkX7AKmd3gkdTgljGn8JmIh+f6JfKIYaO2a20xUgr8G
I016NkpVPKQXZ6jvwUvWrwNAxDqWO5wZoeIGjysn37OntlNVy4DkheYkvdecZ8VZ
kYAvlPIxfFisyNN5BK6+0kKcw8QMLYKyoZqZD9/SdvhGIs3mfZFnFsgXMZhjU4fQ
PDyBiRCf8zmiXJObEH8+6lot37zYxPpOVkNFKK4UspWHDFoqo8Vo3zeKhDeh/8+I
pknKqDnad22b5DamSJrb7DTkwCQup5oMDCWDxJP+vESZdTuZkM5WXtGghhJuXGI1
rnLHb2qTfuHjeGTTkvS7ffJcFE24UVcWrkgQp+3lnY8zkC7ToVAXJoRvBqO3MO4p
AF3in5tSrQ3yt20G4e9uEVCabos8rxco+tHcMdErE8y/vFWUBBFOp37iiWuTJXiF
2AJX3JAczFDToKvLB6kPJc3lxemFccUstEs19LXoJK0R0oNIW0x5BVFxhTA5VCIG
wpPzDIsSp95Q7pYHGkJBpwdQC6L94kDjkzmOUeJQc1IM0Um2AxEjJf/KVfd4MGyM
e5gC+X76Oln169LQMGObK/lZC3c4qG56yMT5tu6PG0oju9VlfLwc2NaL1VtYI5XY
J6dc25UKITk82bYB6kSrmK5J2NUJ+ztaLebthZVJmyvIY3uQ65K9lj5nmwE633po
0m2WQnOSagBVXYEO/Q1OUAUOr2U/AbgoY1yoowtdrdWYyBG4JVZU1NP1B9GL2pT9
vKaQ6dSajJxIW+tbOZ8FuAiLReWnkkoYRUMR2uwSR7+YswmfSFO1XOsHBeU7MNRi
eSqjFVGpjMxRECnlhSoEkp/XvdBv9JIwj+iBl/ihq4If2PQXT2GvBnyR9UYZf5Mn
WRa8BEJGAEbhsv1uieaETYQlopNpLJ2te/kMGXtffMHkensvjmO4CelUScD37aJb
jz+AFD1975ZzULW7DptWWJNUA3MuKefxolvnhzLgIXFW//RhkpE6zkBf+WY5hOVa
vK5TdHQ/NypLflyzgYB/rnqFT67IAOG/ACetfYdFDtZB/k3mjslal8wMnXmO5Vp1
TTOTSXo/DXBPIjwaVExG7UXH8ESxtLpwe/9rIi7qz9nzO5va3eQzELFteropcFCf
PImW2PEC5WU33XHwp+TQJM6p/ZIlM1Cij09OVxPBI18Bq/hQqnQsLI8mcIMtSS8U
17fpnqTyOQZolBYQyN4IlkTC2OBK85aTixyVQQ8C8lv9jBHLvUPWbZmtaw6jXo6j
ouufsoSBs29QJEdlCjtqwpOXwQLz/sYabdlUr9luMEz+R35vLtxTxVYCwoUzsK9f
ERMAMShpjUVpQ7U4lbfU1/w6WS+DkCJY/4Z4tTnwQEUX85cBrAguBe6x/JwFH+9d
U7r40giCUq9/uot67LZiNEOGbsF7Gz+YVsNeCdRdqsph16bxVqNxT1xfAlsArQHj
/sCgwveFhUuAZuEKGPhLmhxgs6ge7kw2kXg4ZeizcNQ8q9jKdryU1JW8YKK/x3X5
dQr7aiYJ5LpSWrLu8WH67nV+0OQySu/A+MV6IWxfhy80aDGXz1RGO6Z929NemIgk
ojjSIcvYV+QnLiOvIfLXRS55GxyDEw0Qzjqo9M88hdNt+ctF2YxTZ06hCApZWTIq
Fh81GuVl3AQ96u+84pDoEqSpDeU2tn3UGek/qbePt8F1Lf0/wLNkyBirKi21jYr5
Yy/trJrXYAbOZqV8zC5XqEQ7D25cEhUYsgKpkIYIHXsKI3/U8BQ/KHIIQhKC3RoE
6X1jBEBRfN3n/F+GhlawN8l7tb5g/aYg1Ccrp7ZI+6Q9DkYKgaMhSpOyfjwJUFBR
XobW9ZrvUxzlFtcpo+p9pXUZrtmt/NY6iY7Fn3kgHDHoPAEFZWMYHeQ9NuAC81g7
iEioQIJgsEPAHPRoA/pGMhRhn4pggEQV2CQsc0emlkEKWTWtDM/6Kad842xaA1KP
Z7V6WDotlLoFcIhefSnQ7FkdyI+9Wp05XCCjJBAlXZ0OeAJGyN2hret64K7r1DH3
6wAQImpVQDDUuWoVh2WS4fyM0wLzGHNWsLBJsniz6q4gnGlncetM9uhaMuvDEZ4h
7nQGaaDQi3jTtFWRGQn+GXqduznexcbLWDB9XKlNOKnC9Y95YUcP2CYwf513XUZU
5n9s6RHL98Fml3SRsMZh/xv2PX9dC6gRKEDpk+dCMGk4zWxgGYSze1NhJPH/+AWc
7a0rqFJSc7+gRJX7WzAw3/CTS91T5WaLvVOq4Ilo4OmvQlGZbdPw4c0EXw++ez7d
NuNw+OuPZWJrzEbnhtWeaHsQv0wletYCHZ4WNw6hP5GDPO/N5EKFBAkNrezGnwG3
RamR+FV1thdoxYlnD+SSfUlfS5vTOlFvOtl6wqV54fwfL+7UlXQ2Yr0JqN58Qpo+
AMkbQhCiyIM+G1HPFk0OC4mwp8Jh8JVOL8BMOGfltrzgIMHK+vfYpOCnojD9y5HK
A/6mqqCcD4ojVJZYQsdvgIgtycmUSDf9rpJvMexrfY9DRgOFSS0DXRNwCng5SQSK
lJLHqL5D4Qunm3/74IWLBXK7FlJwjxiIUgrjNhyDdoUOgv14p8vpPCbI5LubQRDP
a4yF/wgeyGIC7Fht6+8Gy5oKsR2dEyWI9v7tVOnD3Y2eeuiIQSXYaNi6e4wR4CIx
9tmDtqGU383P5HrD+5vdqvnWWJC+f1WozIdqM7ecJ7IdLgSu+Lgeqzdt/vobyhd2
X4uc8k1RiJyfmqKzgVOMywOoVczjKLLFcnepWQJ+qXmyUxUV6EMzkKHA4vHB0eAp
dRRF62EyLjpv9NpgAZ5YBotvblp6bH+gl0ffULawbZV2l3jHeA0dAKkjriPPood6
jwFYHzq3uaSelle6+EYOT01wMGpjUbkgW6YlmSZ7JukfBKEyf0pN+XDlgmieNG2D
ecsod9uIANQ+3sawLvqyWdvEg6WZNXqPYinVtmjAKTQJWfKizqXLJzUdc55HTNo3
kBFVUyXdImsbRNMLWgm/H0vF30rLpbN24QpLR4O06hxJprGXwzxzBVlNZHJHRL5H
fEl6O/OaiXqqmZdmN4RG5EDwq+q/kHulTnYAbKlaYDDDlNZOxJFQULFO0CIyh0Qo
oXuwkjgVyBpTDn8F5FI6s6viav/GJwAId15rrMq9M2u64HIL5252eci2a0JT/F5X
8hcFhPgEcvT0he1OsiDSLQe4nGCrrEUwLON4wV1A59Pl6yh1tQNBYNZKN7JGjniU
RKQ0FxKv6ynjMe7SoT48Jye1J12uQSrq4BOYPfH3svIaUNHRiSVCOs5q96dUC0Cz
xkeDebQulI5y3DZBt4ROZNqfang48H9v0ujAP1WBXT93zC3f2Q+wwI8kL9bF4zFh
/XBuxrzWZSGcLKb/9IsR1udVpXw6f6tV6sa9DOaKov795WseEoaST1H1nf+sJPiw
yvyoWp1ctbfyYTuT0E1XKx6zuXF8QY42MvfPYVj89t1K72McBMw9AU9dvOE2txKu
CrdaymiBPXxwlZj1NxtYzRAlWhbCedHuLwe5CODw9OQMkblLHgBE/fGrWa5TfZW4
eyuGpD8jWQPUDMmV068vffFr/E9BdIKSAj9mSBqSHjgCtpQ+7M+jxy8wZu7VyaAu
ZsIiS+EFMr+cGJgMiVTFPzgro67wfxHJPKGQZzo8U0FtuoL/D2o+G4mavo/243xB
8vEdSYlHsJwRbVpHzbTLO+ZKKAk18HLyVRHl11/HwFja4QOh1D2deoPyT/d4mItz
lAG64waso2zl/P5P1BgP0mL5I609gkOUBCCjRvx80ttDqlp72d14su4Gqevx/pc9
0928PWDlXYnJwIquIub4DIhmZC4+FtddqoiGjKjFGL4pyre5sDEqBAJUo0NSyrIS
AUIFh+Bp6TY0WQHg8EdqjnR6yu14+rcpMEIV0h1aUMSm/4Bn4g6vC8toa5aYzB1h
1IwPGyDY0/MTQ6fXQMHuG0ktm130XHxWwISv0uGEP4JDv+GI8RgPD3+LXylTyiLW
BFy6CdSrm8ghamgDZUeC8NExz2BY3TJFxEoolb/JvjnbnzfcttSogdROjFM7L9DT
pEdejO52CBau2nnYKPJnaLH5wPHd0FTb6ymt/lqv1QYMdwhaLJDC3G+bIHTf8fSS
jHpaTFoIv4k9uRYDSMB+LwcArfUEG+kDAXnGEcWKdrkjNMYRJeTkgjyjf2ORUgPY
CBVRZN8VN3XL/61IZcRJk/jQFi2O4RTDotYla8Tk1xzerR4754KpCoW7CLgD8a+p
vI7p/GcdcGM/O6JoPYAlLK/07T3MZSWSiJYHmWCwY6hIs5/dej+sJo+luGAMDwXD
xLKou80eQnUKaXR0XpYlnRy+N5akIgxKWtN5U5s/fqlVrk7gjlrwhTYSMS8bItf3
oYwuaj/teRiwUYaJRFxEAnVcBbpBvC9km4T19WreMBWG6nDAUDEvgK/6wyj0fVLI
TKlCs92R5cvq9FwDCHaAuAhod590uObP4zIHU2zvpaq3xwH2zv/cX58x6hhZPZJz
sqS0myI9fUE4ZHFCvxpjkUrdKpkUzvtSa25yvvuDIvO4MPmTSLwcrWgSaNrfCwnH
95xrL5DWuDX53AkKdhMrLpCLpju9SyWUizWjuEnjacMwA5CnasObcrP+wD9vv/Ct
tc8/5EDFRqgn8RlYc8ncA3ci7nBsvV7rMZpyXLyEce3LAKJ3Nq2HNSW6zyd3gWQc
lEGTPBjT3MFBLSn4dYGnltFyBIzf1rg5CpQfnka6ExFqm5kXE5YedMWW2uphcPd2
qpGAdi1UuOk4J1HbRKey6SDdXzjnP6/eRpQTAbBx0dIIFZOdbDAsaDtUE6OViNIM
sSlpZ26Rvb6vf2nNSdAS0YFyMf15pIxfIpwI9+1SIO2MLgHFLKVDqJ23qAmgXGm5
/hkoLZesXW/IiZsnYDixoSf3Wlxi31xDkJ8iIJtq3V0LErxEKt4misU31xf2zwcD
h8+qcDUt97dGmv7b0wEvmWRk78HaT5uI2KROBUGXMU3EVP2pm+TSeIHN585ApEAE
S3Sbv/2MugHmF/d3/WjF990AUeGmOF4w7QfBmEEuwaMMIvDPCIt0jc9VnWm9L/6s
0M58qSrCrDBo9Bq4qwLrB2H7avnb3FsLtms7w8/7jOpiC3OWdV9GrtNeRWvtBjUw
nY1XAB5ll4iPy+wERCOB/Fa+oeSuOZ+pFi6JGu0HbaIytNi1+zUgOxQf1a78K4E9
13FwxkedST1WLeObcViB8XrQU0aMWjiBe/Yz/2+kcTpIRcxMx82dbCFtokJ4INnk
ZxhcW34TAzeWBxc4n9h0Vol+cRM1yohH8q61d6hPy9d+ly2C9tlVJlp17mPQlVYJ
iQ/p5/xH8zaxT6LhhNygvMqHuysmJrhJWpwNajpHxa+gEd4kSEFMhpv1e5bWpOPU
r+JBEx1Xm5eA2Ij6fDrTTmaeKL1old8qSYfW8eMj7tYmDZujolhcJZLQE2HtEYcb
8y84uy5iprUG85UR3ochtMuCH0QPpiuzX4R3w7K/gnj1Zze5pB78hUBnnFjRiRtn
5Ta+iPFaI5G+pG+Eye0Bv/pf/YDG0KqIK33RmmtPPFmxHT3M8cIwytquUNTflcC3
+3FIeflqbc+dGTZm8yzLRKa9DhkZiz80OtMlNOjKYh+tBYdJkpeXPmyNey7YdOO8
REZp/7WXn93XlMyS+EtsRP9TuWVW61avNFvYHcf1u3U3YBsdPH3lH7qP6Y2ofag7
jfYFmKtJ0lBCyh6rAybYfuxXHEwfSFmqjqApakT3oViSB9v8qfwZHCfn8usHcW+G
QJ+pAWPlCN3RIHBzIDsVgwF2ERmoEoUA6WoD7JD8HJM1eCRma1kefRsx4uUMgURL
Xxgvqj8kAfyPp12iBWvf8vVcQn0e5Oql5MDT/GZiiXTPhK86xq6Suw8PFhGpt8Eh
vYvWRli7v5RROSuu9z11zaZ+rL/mpeP5hvTKOythHN5R+YM8Hb/HRvjG8kIJtnRv
yxjikcBGTwOEjcJX8/9egzav2vZ/nsC6GsNZlNhfrTJtqDynDUvfFH355TiUppZO
c7QQEPuHRbFvB+Z1srlW8dHzySb0RPBgDDj6i5I2eM/5ShmWKnQB6j3wTJ6PLOS6
zLGwT9+X7DUH0fChUjEV6VzKhTrrIKU92xuenCrzjS4akVbdTTjSpN8gFgQNZl+v
QrBstx/1KDcdgYb20omZYRcRDZyQ2eFQKJFUefrLeT3UyPyV+lzSD5k50wqgm5Yr
VzJO1z9B+pV74o9MQyDBvZMOP3KZ6ZzrgiR+Mf/G8LXpHxZjBYH29DA/hdyCuQ2A
APYBQCMfcQKtFTTFLylFEyXfgpF4aLc1vAJ6MO5m0SUHoUuWR19OERCQV6JYhDzP
OBIEmxQXJr5bl3aAJKtFO8QuUX/TgQMlLKdyPmmJPV2fsPuh/ek83wvaun0GZmVI
nz3JQlKrjz0jYIwUxmk5cCiy33jMpVzu0HiMnHZyO+4laNb1McW2IYGRuxav0EZ6
kOHCk1Pzj3/C6rDEW1AaqqAN6D7HW78sywzUM/tEZyKzeWd8CwNpXJH9Vc8K13bK
W4o06pX2FSA2q/HrL8HLGOaPMSVbd0rK4R3Sjw/ISEFLI7XQNmtwgADh5tGyGFu4
0XmTrpAH9TBAJXA7h3Codl58OfER5LodKjLFd782VeliqV3WIaFEzsaDmXRyocT+
5zPfRQGWP8RaYMIapTvHcUCWA9NJqXKtExZ/FgtAQIwaa5rqFN+ceGgnmxju5eEA
AvbuzNDRGYq/4TZ32TTmFrjmKDZ68Mcd23hvnjTHsmrlKFIETQsLxeatoVMRHaAh
4CPkvd+6UQoYjVPY9kSLzg8wUtgCGpwiSWhipzgO9/VNCCsMi+kZ1U58ztLTHeeI
LF8xiaPkM+upoJPfIDpCqNJpybWQpLZhmiN1UPXgVgn5fJ45DyH5AjDrblztqq6U
0UgTdUNaOMCtjjHij2sx0mQwoH3YVvpnrghym8Q135cGRcX+TxQ2jHUhwdU/4wdO
OkYakqr4ltOv6MW8leWV9BIY/3qSDODu+qhesaVMmlFiSsq/rYDvdW/yqpufk1Ge
SGBsXozXYgNeLYGbnWxOyuEnesuenzYFT2Q17oxgHTXrDQqL5+ynH3I80GDT2L7o
BVaNc8djxwhcw05f7DTJtVGlWMfcd99jrmoWGZVfRPt56d10W2gB+AlmjgS2zPLw
bQepkqJx7JWzZTrO7ZSfLVG5p+AA94twj+q2DZs6+92ORPd3KRfAsodLcnhC5A8v
FVUZzshPUV8IWWkkxPWozMHvGTt1SmoQkWUUv0KFI9Kjtt9Z357vEuSLxGqZC2sJ
TsnW1dtjQHzG/vPS7fBw/eGsjp8WxWnyQvyaQVVkQ6v68Cs6HjcPDT4Ks5Z7bnW5
ovphRZmNYTJwATN0wIoOon90TlhzOM8XgxW0/4vJ1xP3ciLCCdIy/Hqh4IsAXh0q
ycqnL40yNdRm7Fr+2UKOnfFzcd/YQ4JoK+6LvKPMTkLSAtpC3tTBzvOS/5Ww6FSB
2ghGn8dge+IW9FP5JCppaxDobDgLN5rS5MswW+I/1j7SpE/jqlABNWPR+Y0NkXU/
s3VQ+vv6iC4rgCrMwRhBuVydQ/PdM0czLyJISjrjG3ZnsP3MCOS9ztPeIsXEnrM2
csTtRusDXTEG1HKFq/tP69e0mXx6Pzks7BL6sUAtPhQ7ldDnRrKGUM1veDr2NWgi
euPiahNNBJ9DhVHDzt0STuc8wNYTO0EO0wk5GzpBbYCp7NBgkwQ/Fxh6OfzpabpR
BLdwwvN55QmAJzOmFsknOym0ek3sl0DEv+i336IUyrpeYWicQLw9QQyPwl+cPIOJ
Rc381bLciLgUwD63Ho5OLtE8uqljfAw/Dx+Z4aWAXvV0aibuEyWP3LSotE28CBYz
m6zjM9OeZT3AQx6yuYKNovQadslbRoP8Lss24I0Ci7xL0Fil0kE32o6ZT4sT5pyY
xnfROA8gVZPMjsSPFxhywQUl1Crb2hijaefwJezegDvweuTZRMIoqKWrSygJYTMB
49zjHdWW9DvQYbMU++9/LTgvZ7iqn+FAg0XQeaa/n7FXvDnr+hhv06DVeYyFacKY
U/bPqrTdcHsq8MG9zmkWUGt4t215XfRoh2DTYoxRbRoF8Q6gBbSk5XXRdrsQnkMm
pLEIYAbs6xYX4iWtGcSFnpMWhiJoZskHV/5wfto3y0l/UFRtgN2Xio/mW7M+N0Qn
MyUntdfkzCxgK7AavjHXjt1bxPoYhDXj1OeVqDt4LjZdPN6y+lOJH7LEDiKvjbmY
dhRGpdK+Qu6g/0Jhi7boNSDBcXrN7ar/uuX5CFMTn/nz6k1kKVAIduOVd915yKsu
ML5OSE53l5Ms+ZjM0IknEXjmZnFVdkeqlBZGA18wXPB/GZkp9KjNwx/7H4ST87BE
eR7tl/n/DoRI+pVZmwDm2fPhNPfyXDCL8nmN0yrxJYgFebwYXmQrnkTDLP3Lspxt
Ry8qzIhxPC+cqbx4a6uPtri0vynytuZIIgkevjnluy/oqiNiMO9AAa3BhJuc07v4
UZqF8NB3yoecrwBcdANkgppXKFZgQCkih48X5KCCVn7intJKzJmADKD0Zz6jXygt
nfzOBh5ZbCe9lnWlWXmZ9loJF/UNueQ389izYiUG5t8fu6lF7K2DmU7qw04zHSfO
/aYAa8vHDzuox/9P28VONQMimEubac8KlSksHyCfE1POYjzlV4oHDRhriRXnl/TQ
dJGgCSe39WlvbhMMymU4XliR0ECK3xNnt/yRBBjzDpv0fbmAntPocdoVaSmoossZ
Nmx+bpLs8lvgd2U+khcHL/ksrmsuB97JLFopEbR3t4hCS4DC2B3cmxm27KPdt0SD
59tum330NLDy1YRRVjkQ28Hg22BU9K4pAlx5V4fiR1u9amxf3ZNUlavX6KpB3SXA
C9EfReA9FPnqnIJ94KrDzAjLxYZ7VbSfywsY+qkZ55bJ6B9M+yucRgif6wGvsucV
LmS1JGOe2j2kuqC5ybZG114SaPWHg2hMG2URpkymFhpaJ1e7w9fyWPkvehe3XGW3
W8yKkoN1M0HZroKQq2Z12jjbuAVMTbpbmit8wD1CExHbrZci7rA53LD9QjgAC0wZ
87kkT4hcl5YP894uRY0+NW5xwH4Zoz6a5T1fJhwgUWbuFIKgGkTS3cOSaheZrxnE
1Fs7zi+f19reqmip0gE0i5s8raN90SufCy+3Ie3FccK7it0L3+T0w7OhlIja8sW5
JRL+4XVkGVWxzZ41SoQbsmgkJNDTLmsc3Du5xV/k1atGM0AMr3OjJLGH8V7h3Yry
OBFq6OPoQ0c4vsOq+Vt4Lf8/AegEWNPU4e4byszwtxn+JZWmz8270Gr2Do8tfto7
9bmfGsHGP4j64pIrqKyF5PzRYV06VgbMA1TW4e/ycwbCuF/WolhxUsGIGIMI+jig
pH7X/bxmT9s1/qjdNExYiBOjHBdCOHJW+TvrunE0xNfKQhKgYz1LljCd0oCJnWCU
rmId5YQJ146FTsxvkD/jepkalmDuGnMav0TzR3A7J4DDj/jlrGcL13CNBI6fL6ko
/Q+LLOWsfpgaHfNtrrYd3nPCu6M00lRzsodIRA6/9HQLAFSjyAz8h1rHuq/KGCgq
9kEDqExN8nl+NGOfUNVVu0jGqLDeDSq2pul4T25lISK8Jg1F9BzDQj+0M7G+wCvo
VsUhN90JkKGImCa8muuwO6mpU5IfdYOU47JnEc1kQ8raq5ml3bfQwPPj0rKTyMDQ
xYJXNMZxr+CBPaXD6azoCDdmUHAVmpE+bxM3BdAsvDW+w6NsGHscwiG0nApx2ypl
aBqRv1ViNK2H7vK7AG+khyoUbGKs4vf76nSPXg77sH9ygsijufNLXvRHrrB8rdAJ
U9abVYRfyk09eezgr80N1abFihljyMf+5jxfcwblxYtrK73nk+3ETutHN6lR4Ojl
eLZfBgBAWa1Aff9JQuEPfwH4YlCgl0/LkFP++U8iBJgbP2bassVUEqAvyUJqEauN
1b11+Oz1fD81hBiURFQ2aaM9/5G4XwPOfhbswyL6XPJEfBKVZk4FQmw2lcqKgUw+
YDlRXGRQ9jDfurLPMxwhrC51KsoEGrwzLUdRCJJYeb/8xNg+T3li4dp4WMQ4ggWk
DxJf5UT+T/TXeFD0lGEN/CvF+88vRq3Dj8T5lRrm2j+6E42XS45lPUa9I2ZlRmJf
aBHWfCZSmI2vobyyXNRufAm0OZDwQ3X2CYrKbLCUt+MOaU/0A6+Y8EiqWQ90pwR2
N/tuaKCrISSYspvV/0zNvnXAFHi/ih2qYJdirOfoFLFSoGbU2Qg3oMbrucAlsHFY
sfxjcnAf/QVEG8pgyIUKzEKnPNe7g3XdLnvySHO323a/49Duuv2P3X8MM9Lf2Wrn
LMTpXOEULJRIo3ct+epdEtT9ry2XBD4YhC58nkfCc87NXZYZ+6RLOkD8HON+ktFT
40SlYUIpCH2oNvWjWQ3TMIG+f1usEW4H4ohpD2rO4ClFLGFtSO10/A+CbT6OIn/Y
5xCmd/kESCnRNnbmUMT0EjnWu7dBlpzR0iC0/PoNaAcOJ3M1A8l6JN7Hq64OSHx3
PC1iM5OSIYsqjv+HS2Z6C8+7BdgXTV5hNISVIESmElLyy7N5c8O4TK3ddxJFQDBF
I3C4wOPBe55EDzLVdfeWnkmF2uL98rJ0b94oZi9iIjlxK04+fcGy/dsL/ZTHucWN
nO6g6ExNprUSGFbS1ImOfrZVncNIFqeyISVRivG0bQ5ad9BiWw47SDxfBudJnMIo
pad95Feoktad0Rbg0A0V2NYB6/Z4G1G4THh/6KpXIdDya+iTB10rfA8tc6EYnFvh
yaKG0O5+aMcSzHnJHZAb9OEJcTKUVcgaxNRK0DtXNiArBg7wEQQVy7DmENoTQf4O
7TkdJ88ToJojTtjWC84NpoE7qOvHesjwmjx3p+YK4U7EkrNNFEd0cI9jzPhrAObD
ga1o0s5UT8g3C+gNfYep1gmO+hZD8LHs1clU4a3sp5LuzHsM+Ir2iVUzxRcCpja0
dLFEk6Ma1LghbzaDvmEela1q0bgoeZdJqendHMrM74t3i0pBcGmz9kJ7i5ETTbsw
IJkqjDkHVz8Fwj7L8uIiEcK09Fwxu7pR8wxw7uXWKOcNC5R5NMLBzHcGSYEuAaGo
PK3D848f3xr5IYEw8lIFP6Lc20BO6J5floW/h0s3CLLBuiECKA1gsDzLcBQFhmUB
icNGFXd2PfwGHSRI4injzGsIxTr7C/tUDlwHXMtbsUdh+u5C0sA1DS6sbjiTTOyG
UQ8y7ToODhPYmPkb2W5sMpm4mWg0H4U+aHrJnhyKcRQvciSX74fPPp6u8NepMCny
DEFIVSzM7F1Oxiuv1mVwdU+9avYSCNF8yI55VCWQa5gTfqTAnfmU/EUBA/dl0HXT
KauG2206vvB9EZSHjZCHXsUQfA4czfyH18HA5S3yI/M832vgP2ovcGZ8AnWti7o8
dTeGQctuuCH19k++eyVc+76eQNOri59OGC46QENkDj1E7clNQvCw/Rm7Fj1FuLnP
X8obfIL3icqw8QjjrSgHTi6RYABRUzsPPfVlaxV0qYBheR+MPLcpC5nErAaQnpP2
pGMN+G26LowTXZAzp56j5eCAaGmoZ6IuYR3VsIzcoYkRE5UCxYpVHXVGn6UojUPl
M2/1JfPLZv/R6Gjek3ejU7tu6jL2Qd5zkSsQOPWYuwD+ZWdnIah1F26FFzuniPom
/l9IGAaQ9NSmC5FQNHTKGdKhnAvvd2uI6VnHDc7XrG+6cNwJziKamPEmY3rdO67t
WbOmlMpjKn+8f434HsPpKayqP0edA2inEpq5ucGfGfANOeHcfXil5kS/gcH6DRZ/
IX3Pw23q8yMOHeVc+6YmcZj5GrhiL7EMcmYoHhgF6kx/qIOYn8cyu+pcAL3YdDOO
XDPPTxT8pDpovwsMRPYnf7TQmBOsirpNkOMWLHUKDmO5i3I0DNI6/U7z9SksFTUm
cljdkK1t4nSZnEG//sIkr39GTtCwyxLGpfubbPQI1EPr1meSPbvtdN5r2ZTyNhew
P205M6391gdt8cJlrdbdZ0Hh5g+Z5H1vN1mdo25h0HNNnnLjW3Shz+4G0BIkqvJT
9D24dDd4m+IfQTQhUcuosKUgFHM1R+fE+5eaiXO0fj+IbmYc1yB/gRH/FVjFTUNO
bIQKJ2SAYP/+vymtBUejWZRVGFU+WCAGvTOna+bJeVnlIms0dv5mhg/Omq05/cXE
Fdw24wobpHpFK8R1axPy4Pry5Ya0yu2JcdOMEF3MQ7cBxpPYr6dPbCzoBdjDImY/
Sdr+2eAuz02kQOUsUCA02FeKgCyKx0IyuNhjC3C3kqpdT0aN4W21ACbwenRW69Gh
ZzGHPQqpX4Bgwn0PMU1W7JPN4GHzQiOkX2wOoGz14i1RMAio4ZNyVGAvnOheg874
y3JJEH65VkhrWPYFUGRzvjOOECLaSJ2wBBOgbbtKIuXtaiSCjOjettuRggNGTMbL
49wwiruJZPra1mb6NeRcf6litAlSxISnsJgN9cBJEw6bsbCdhJAR07lez+uCSKlL
LY+Ix5Z6QV+F66k9g9JX2Bc/6IZxDjuBHhX6TioqYTNhnA7OhJuI7lP9dkBNuvd7
bwIKilqavtkOWPZT0NRTjdfn8uI/al2yJsBh512XX0eZIRz4SQnLMLojFqBDxYfr
kIR/6ZSZtgzimzis/k2T0nwuFwY83aycEvYBhSs/RaHuIjXCKwEaTNiSBsm47hQ3
g9cyD0fePrjxY33O6XeLCPPYf8Fog/C3UHssfF8qMUXT0A3VoPVDmSrgWVhBGjtu
WFH206BID0omTAphcLu1jPh6hl1/EiOddhpmpLzZZHLZeI975MPC2M9F8YR47mdQ
pk2FKjWEw/Dh2+UhOZiLrhbxXoN+9NF8tREeHaT1G9eMj4hNbcve0FXhk9VsUetI
CZzqSTzOBQZVLfm3J9mJMcTZ7ax5JY4KRbc5G4w36oCdsHvWD7fLZDU6OQj+W0A4
VgAoQDdr3VzvMY2gKSTw0YsYXpdUcGpqjMwJ/M7rm1bfAMyt2MFOcWo3NdXOJu/o
8KMIRexivkJheVNIDDJsnDm3RD8gcXyowLMwgt1Ew0yV6wbnWEiZUAHtC9m1+tLr
cuqXyzHI5rkVFpOsIoRzjv+izH5KyHaCvJpzDuKbvD1bjHifxe5/NarglHiHBKJ+
mj7knPJ3ZkX+K4wmLInulyvYLcldZmaMA39nKhjrngKcHkZwqtQAI+u9kiFfVLXV
Zn+ujruFQhrHtw3ZY+WibXdCDXV92UmeFwuT/1VbtZV5k2t2a/IIFZL9o5Vj9imA
qsFxM2KK5nJh2e9y02x7uHSE4j0Q5M04VJz/Bzse147XywvSg9DOuJbIkZxvkEE0
Zh8AkmnT0unZ7PwAZnmUjOx0LPDBKcUNDBvN6STBB1uOQvZbBvyooHzbtCENjNyv
EVIM7blyK2JzfdCJL2dkhY0MXaqwRrQ4OHayXgmrDwU87jVMx3iPYxMHcTmWJtI8
7u4ImspaGGaHjl/WfySTLEKzTLRdfvJvwhLMMpG5OAtqbnQTIw4AOh1uomhUnTRL
bnND6PjgpGb9akPHKyuhNomv/lCTmgzFOe7oKQXHW2HfqavD5KyNB/DgKje9djkC
7nT7qZlMWkcLXiHMhr1IKXguXb97bkX61yKGifVf/mKR7FLXbaU682NfqEI8u9Y3
zBlOhKMANGYJ++suLU4/IhNgqGnZwfpTFLKkeeDGNoLnMjdcKxo680VhCR8//xvD
1YKl65c+fT8ODIsm0SQqXyPTiazuGQMLmDMxJu+xjqfacv5ypd8WhOgpE1WOVfEO
Nxa23u0Zp5tZ55qjKhntvs4fLbfmrrre7ONZHJtThpN2Kb5uFlY4BbfyFIBORkkU
DClFIGGn6rtaFwKBg2WIJOP1N3TZRQmN6X0mW0tWGwMtGM2v6Ad5+/W//arDUBG8
eFlybpjsgxJGja/y+WndduYBFw8wy8h/4XdbZQdpUw1ohz0oV5RyPQU8F8HPMNW+
wZZfd+eho9YUvXuSPpsj8KxEBBuVdCDHEQf+GXA6bcbvVxNQd8Yv/sazsAHfzq4n
ZHmobM13zkrFzP3XhUJrJicVmo9p2YIApefKCbaG6cQA5lrTI0N1ZDvAENyfXbs1
20gehWX7bcZ/pTQlhQTSxx5ejHz7ShjMsijU8HL+zoP4gj3oudLd/5vtaP+FEtyi
xqSuc3cSRatSCTQ03bI3+okZkgTKL8sabRsyWNIue8qDsQKmUi4ijQFrhVM5i2JZ
TTOh7X0gr/YX4EVU0/dl+qHVCYMwEL0CtoCxQiAqVOp7l58ATHRaYnWWi5jfFTtB
YNKtwZmqMliqIMvrTU6mtJkdP8JTEn2TiiNbEF6fTA0Pj157iOAlhdyoyXJFBSDX
Ae50y7ITE/HFJAoabqX5p+nLBsCxO/VCwyWmC0f2Cf+fZiHUsgoDDIvqbFF9ESSP
qnUgoAZPkQH3Le4ENqNE9e9bplp+L/TrQqXiv0AGS6NMM4d3R+B3mt1Yyhz8Eh6Y
MgrPHIBh38/ggIVkfB6IrQ9o7aRdmmzeRwG1Sjl/6w+pZEDhQ8G1gqq2Mj2Sc5dU
n4zYrVNld88SFTAerwfq2mljin1ftVL06H5YDPApu94ibTfzk3zKhpflVBDCCWne
fmqifQjUTcb9d1NsQmlxWYoQATzpBTkJ3SMIvBb8QD3lCaTIm7JUXQvN/7VFeHAu
TSfQjeN3Cvi3nib4uF1zkkL6h5THiwWD8DQoxLPblT2lDoGFNf/1zKwGLi1jlgji
5J6dEJzXSheMp8DCkmEbzbjkN/+Fvt3oFetJ6is7I1uTcYb15WpS1rhLbIzXOYaP
mOgxw9FdvrdKdXvyRLXZBLWzkoBysLlMKGdfYpjmrlLZXgQEocQl38YzHoVoHZuQ
aT6tapl6pmT+ptziyMx5aMmPDmABgzUHr/K8L/axgaNtEyq4h1AiBXnUMEHXC89k
R/meG3xW8nm9fT9oXkR8zz4qtyKuxwUlM+yIo7Q0LZcZbeW6j2S7pV0kvPKKKprC
DS7XeWRVo5MZjRA58nt3MZvMiwJG0s9GTExg3y/rL0e8/GXQkg+mra4UmG3qGOzK
opFfQHAg1SqlsMmjZo3If7cjjONPAFEgWWkrFa4HvsYeyW3JFhfihThhVI6JjTpc
TvvbzZClbdDSM8TBCaNeNPefJPNLe4WNGqrygsKvD0MUvKmsYyyV5/6pXjUDjzv6
2VtTzarKJLphxZ3WKBVuC8VlK58dRERYQrY3oAGMmCgZlMR2fCevaiXcFocgD+NV
agR6j0MQa0Av32X6qUExyZiPZiVkrFf1gYmcMWd3xVdffA1/RcDoYrJWQvzoQ7EU
KwHW40kd/ax9iNUcmLrkdJ6whDDVQZjKDwpGV5Oo268hh5lpEpvgY9y15tZld6/I
ZZhZSf+nOfjm/P2RF2mmKC6tvKeocDJU29U9AEMQM6B3HG25DjLn0NOwCq9okPM/
Eh5jdpo4yLiqS9FcC2Ubxg1I6mEQ6OMXNUNuiEWCtlFwSLgfB0yRZW3sDakloX05
FlKfFFu7u7cWukBMAxENzRaEYhXQSbjanoqr7nFUpluku1HNFwa9BV3DoSdvB429
fUlUqVLSM7y6ECHJ+/qeX1Wr9Ny9QBoRYO4WAi7ZfBJukGk8KQPShlWOThzPLqQa
g+F4GKE0/pFZRUQaySLuP6V3MzbUYxvhIdAvoo+P/YX7MoZbmYcEHjKePV+eG1eP
h8lAcY0OPb+IOug5hZz2dUivkeMGSWPsSqH+63fpldIcW1qJ6NeI2Y9tNh1FHK5k
DP9qJVMoLz2tsCSZ1EH02+sl/zTUt4GjUHnSf5oP0wz6d5tiwiMXKhUGlTgyWDF2
lHBwNyk/DAG4V2kDEAnNG9UzdHoWlcYHT8ssU0M5Zih10f29Noeh/Cdv7VEyfyjJ
KwTGECW8AbN+PggLclez4DdQUdKDB+ZGyeAvaE9BL8Yqe3DJpyeBmGD4GGwJpvpg
VxLoG315wKMLW7v0Y3Xd7No6ixuzD27vWzGBnHJsq0R/B3cPHgMcLyASkI9nqsqX
KsQk/3eK+wiJL7KUvQSAM58Q7EYQHv06ji781LGXXPcCSqVbifbA/Zc7KlOsN5JT
g0PQtS9WfxUAoa5Il/RvY68AyGtKRMESHQeNpcoF71cmClJqeiV1k6G+VTjYIXZY
fG0Jp7hdCE8CAGPeXnTH0zL+xqZtvujdGeYPBJbAbz62HsmeZqASsbvIpbfhOGWh
niEDZnYk4JqjubX9G+07IF4THu7HMCeT1zECnOICeDxdpUxUgqCItLpJjQc9VRKI
MUf/fp/Gn8kHHjlMsTdYoRzEyFxS7GKzsKE4c1rnhP9MEBhVChwoRtPu47HX/ile
2xz5tl5NXP/r+8+6MgaujvHkOQ5KoNwAh/TFfCphQQu2LuvQ8O3+DBrnxyxKTZfF
AITI4ChWHQ6tRooO+EXOkXytBmudlUEY+ah+QZElZ1g0aniOiRGhpKPm87fgJ/iT
azMxtlQAX2ORLx4GXTGQ5LrwJzRMKYkOnQdZxrPwPMQ5cYVTHycRF19zvLq43L+m
PVy8P3wBkuAZOaUZTY+bIPp8p8S3eIVTqZuf8J1hbZUCzVH0wdLtZqRRIuOp3BEy
R8lkriFosBMK3cxV7+yI2UygjXnyO6H+7GWikfZgqnv5Pv2XLHVnvobaQpEVGQy9
YwgPQUkKpSpPfP/q/MQSy4b0B/ptTSR8feDkijvMmG2x+E3U7otWTHunGF0haIZu
Y/A87+A3KarugmUPIcynUeMFQQF646+NpRTBuv1k3+C3yshi8RO6TZ42VMOJFvh+
N4anLlFWG481942ufCtZVyAMsyRIItYC7/cHJuEkHH4j7JZ46vsuzO4W5COAxn0+
eautVVoP5cW0dxoh2eBkpvG1lU5tEasUFS+UvvfMP7nH4y09G1quBdtdhWRWX/EF
cbrpQvfzlE1SHoLa7efaZrxrOwWGTptXfWBcOTn5pOUX9Z4ZeCqlKXWcZXjwouRY
E30qDm6Sv2yyEPuGWJVwkE4hyDk8PvVaO3c2KPkIS2xs9fObZyeRIJ0f2Lr8HPAf
q9RRw16wZAo+7Tgy+5WeCncB7eBUnDIbkkMUy1RdnRgBn0pzyOKxIgNMmv+sYBRS
ALDMrNzrgPAn2HCA8iuurNAK43LjKKxDOM0mkRO1vC2bwWRzWY3JmX7O1S0J5Dfr
Rzt8XMFvFIK3h8zX6XvX5uUZE9Z/ziuBNVNmhW0Gcty2dYRgjYebR6D8FLhM9OVB
I/Nc9HHpb2S16lNjloP+RotWeYyu9o2oy6aKteuLaUfZQ/fVgY1r34VLbeOqZ6Gn
BngNhjJj2KGWRN9TA1kriLdXmLVCqc/OiNB59yTYsxpRT2kGvNtcZS8OajFZssIz
z+qtLwBXSJcva/cYLnOak301S5rGhXtBxdySuQ9Bnc2ACSrcF6TdCLsCIsvI0mgY
SG846Ey5F+8P5P/i1+4N16W7NZrP6QOqXc/XdQ83wexBpJvyrwdQibcdxSWVnIvo
Wz3crpvHlxhBmqepAF6OpDi56KgW1n7u9byO4XRN7GxKk+1o9m8Jmm4sW2Re3I4I
0udyH6QCS2/1ovmbDpeNDZP0FDSrzvG7USnJWyjD1p3s2Hw4qjmuiN9aE/R8C4LT
YyTxauMDANoRNoF2/+WfsoCZab47LWEJa66oW1lf+76NAZLSjQm72evkjKU9VyZK
okWIYGQ1vk4mrf2/MlzQe7EVAE4ucalrF/WPTH2bTZIdH8stqXbMaZr1+KyzKTuC
4K2BIRRUHW2KqZmUK16jCYmpvWyl9/LvGfj4QdkechvXr3YYDIlTuG1kHJaa2qfc
HJGj87km/cI23THuoCzS0g4ijHysXHhhg6oRYTfDzLd3jCH3fspsdGEQ9Ivsug4d
EvOtlzpYA/aIrJdNl59NQJmswUqRora0riIssjEEwdUPODTE/ids3pzTLgk8JBOo
sjgG5XVb0P0oX2EugpAAe3e4SxKzgO/Wo9U7eW7W/cgQf2I2EGoQ9SDBw2tAlaIc
XJncinlFuDpOJ4FoG8mIweBg87GOAZ4BCYd0sIvRyTGVtw5cmi8Hmb8Kgf+9MHW6
fxfI3L0KQqkNn34zUtcGJgcpg0M548ReB+RcZtthUqlK7qnJwcy7/H+KXC0tdiFT
KubM6CXDkOadlrg6A8yfdS9B2t/OU0PSqULPOVgP/MmYt9/lgE0C2tSs6Stq1zXy
PUwG1BHjFo0MetsSB07DxGrslcxLRqaU/1W1fVoZdStabH8YYp7FfdAfkWZeZ+fg
Hb8FTe9RG2xKL8HV0pa8bEDsw3yT98YfVtmJFoOXWQTQtYocb18vD0fppqGJWZv9
RklBj0RLPgN59RmqeraEGfShY4mcOLiZMgIyPDdCLci6g0c3e3kpYHfrLZ9brCyd
8xgDDfuPdrYrjUhGTOXgOHTXbtDgd1DmY835l1ma6w3e7/RXaq/JHXpUDd5JhX7Q
H8v/h8kOHdygWUNjpl5qNyLZGCJS2HPbeACim/AcwB8EXs5SHw5AZCK9vZ1KKzjU
c+5wTAcTas+fKzyURVmL7d6bZPPFaxjQUgYClyXGD6SfAljJRL9sL78EuCBnTLwy
Z95GDk7bgAccvj6pHcBWroioL8wPchDYxGJm8xldg8ok2GcLGraHZfqxI8dVFx/y
tOXM12hRWY+Tmysp9Z6qFQ2R3TrEMwWQ1KaPUBCo178jFX4AeSeq3DKWnqXqLb9L
PBPZ0HcMIEIQZEQAGKdNCm5nYi1tyyHl5Y0xQp/vbaXTdG1ho/ePgiy9GOHIx5js
HFbqkBQM+OQJBkvFBMAGotP843N/4ujo1f5ImHYIGs4fxFrRwn/IM9S2yZCV3/tN
JNB7snJhATQlmOnxVCneDCcbWPcE0XhPoUSzlvdq+DLtwLJJZAFh34yMVCZzvf2M
bAAiKwMNDnw5xNWkiZ0xqjRmtHLwJuzkczYt14saGTBbvQQL+5SzYqMlOIm0AZJc
CAHqjQnWQW3p/u8xlgtEbASDEOY7uFOdNYlGQe6OlkkiS0QMaLeyxw4Nhm/v/M1I
pKk+dBCnjcl3KnMG11sTNbq7rqXVKDf3FQu4ZJ8KtnGnpz3BEyRLRo7KLZSIEOcZ
bd3GoZmIfs1sD8R5KMvApuadWVzGoOY87r845MOmVV3TJn7tIzlDUSa6zto40xjW
H+NWqHSG5Fd/g63Y1+IcVC/QBc/0/zmTqcQtXv7p9Xn2YVk1ii910oATSMA7bgym
TFBT1hjWty12taAZoSmDTD3+rIbrOaGAHp0YUbSDRG0uZAuBqSWwqqt7RdOHRZ/G
L4Sg0xFtpLK6B3fO0xLzaeAbvFpcYexdgFWQ9Y+xupzisc9UOv8W27GhKOcM6c5T
WBVBNY/WWEu3U8qm79QAZmHgrwxi8Gzeze27ZGsuiFwEONupqp6LkpOB5b4rkyjZ
GDhF4neGDHiaDStpvGRgfu4JsSrX2g6gfNDPHN2443eHpnCnx2tEU/AfiaCjnWQi
5umKwSD5FyF9/fs26rYuTKmh4VVa8QsTq+DDhN+dJEKFANAsqRZ3dLoN+kDITV4G
AuDHZnUUz4NcI8jKyNNSDh0ch6dPyH+i/+GJAlpWtzlviizUVTOt+VTp1NmqIaus
bGI97+GoKykIzHlXZXKzPPi6N0IVygUG9WNr3Sj0lcJ5/7fDlWItx4SYbe37sre3
BxoN3id7Z7DKZ7fiWGAd7VlI8KmALvnj0/xxkVjIMU/1iOGXsEPaho0dTrPbTDij
KFadw6eVIkNlcWcnSNThqSCBNlCpm6Hdav8WGa4fwSJdOPEhKuy4/24UCxBN0Aei
ICAooWL8fVPcjXHH5z7rTJOlx6/8ZG4XR4cwPhhPL76CGUWOnhUQ+n15Xpa+lD4F
rU9oZvbgBPwYoF7MXH+uAB6/GvN+knwABnpAFbXo3d3HAlFi6V8XtSYTUkFha1p/
PWRnBb5v7sYNU4ClJZIbT6XCaDuOxkHMvj3ipfODFdxlw0sU+ARCu0aeX8b0lYik
t1K6DohBsNrlfJRyiRd0eJdx1lVPMfK3Uy48Kj/6B4C/VhX9B6X1si6g23+IrcZP
xas2q0mQNSON/6+E6FnlfH8fpVxzBFPwXsQz67Eqxtvor5/Wf4afS543EyChQSbr
zMn4PwgpJwGtvgrsj3EeQY5+jqNWol2i+50yg3nMprZUk73iHYXhe94gSkLzbSmd
wgfD2ZFsZ9wH+wNR1MUnZGszrSrJLmzN0OEziBrn+GYVowDPOGGcF2xHc0BOK4Wm
o7FgxtxV/pZXVznecifeaWJVCtmvP+1jaNZM26YkO7HNC2T2yJl0A4ZVbYeTdcDe
OGy/PBcNbV7UHs+M3CANdp5VwRLG1Gkr9lKMPDDwnDqzTimft6HcDsp/3cDEAWxc
4S9q8+2TaGFBg+kXOLn37pQ3INf+YnCbLxTcgydboPdGcmSQ4FpOuQzggyUPZHCB
59zpfX50Qpq+SLreujLuHrQjkuyLv8x+I0LBarcB8PxJL7VCTgoDjTy0ahzHcGVv
Qb8JVPxWo89AV7JzWn9eJHPHXmOU5bBfVBymIqgMlKE6iYUgdfNoVaMj4jyUmWC/
hs6iB6RDR7PKBXroF9FyM527eBZKXY0BVGzEWe31D6yom8cXezQ+1B+s/nSoXPQM
sEOkcw24pyV7uZMFMg1dkQybJO7szXIDWwCF3XX0XvDPmMcvQtx/KPauQeuCy1Ru
4313Bq189SpI1C9sH28/XrG8MVdJrfWaROVmsnDTmzOtlDyc3d+aQP5LPJOzwT80
KF7/oq1bDj/IQ9tibs0pvyyHB3QkRUiRQ9nL2RH1sLzhzJBPrQ82DzxKOcDnwXY6
tWQ1Kjvxz/KyZx/18gpGgPpcQ97yRTp7OMTVicEi/FZtDK8+LUNO9xePGyU+re0p
0J1M1w8+pIU4I9URufVZGRSNCe7DmfMYv9oJWESbxAzS8Zj/yj5qZuJl9bZYsGjO
jJJ/lhfEzwOlUFmYY2LIs+i+2x53iWFtMeKiC7/ztoEtuBVNYQpkNVaEQ5vyIDD8
hOENwVSujvr5ZaQxXLMfIyHr2o/pB4ibIIk2GgUp7CoECw7mi5LB2HPOkgL86j3R
MtewIdAwKuSknyJudpZQCGtxVV9H/jfHh6KhY2FI4H+9E/tGoIr+M01Vt7o9wc82
zuXYxG4oNkYANzbdmJ4HAphYDjELNqm0E/VrSg7hA3AOCbjzkI6Kfgr4ii9WV5xg
TC+A68XKLMPIvOjagYNLSnPuF02Lz39DrCEDLL4zFGEv4AXu37gVUwoYSKxI5qKN
azJtFsL6tBXN1wAku9VjzA3d9c96lnyeCsw46X6VGNLiCxbrywnS8kRJgPhJy4Mw
CA5HlxMgFvmIBham6kFx5TI/WVnzKy5C4jJFaG6jizxtuCq8kTquJtv0KzUUnBoH
aV9c8MxTKCWDdQE/pqzFHDTpgsJXWCx+mJgeaYYUETfSZy0K3pywCe8IySuFbgOI
a3yT5lM5qCLF6lVRvTRml/XWgMd+APTQSD56/JTTYVXQ1B+4lwEql6orX3A4QCHF
QA1EQ5Xy8CUjMl/ct8vlzQuwi4US9tbxxT7C1i+nz1UmjGNNACQ1L3oX9205ym5B
R81dNspvhya9U1PU47JoNhPgPcybLwSPmrbSfQnnKPu9HUkPo4FS/UY7pyd58IP8
ROWE0eDldVcRlEqa2KNwes0fLO8lvvi64KGkM9jLJT9qqibHUhkzEi1T9WoWCIj4
0XPNns5BEFf6lf63otIEAWfraHhTMj9HcX+C5dVi2JWhOJSUO2DR/eTsUlimrL5U
BPX4JCOEvJGmSRZdJ2hVrgdQAOMmRwT1S65IUU90hcGNGBwwKPRoN1ojoF7Q0/G4
6W/ddT+mg0IaJf33iqsa8nniTHsV7HGerNDL1B5Ic1xJd4zQ5C8bIsJzeG8AJHpc
icayPjAwNASTNKjvPBRZqleAPSXeQgeUIY/VfVHloROExGizuRd6FeJVi7jnSjf/
ru52BQzMXwGDN7oXXm02kWjihEMXL7v/pcxMuBbn3ToEHEx1lNaCCkKzas1oFSUX
YC2s8+NVfW+XD4pcHW0qOjNDWIUqovB3krmb7YJntCQweZxIqrU6D2mwmV5EGgL/
cEdxQ2qRMAYcoPdj3bUfxgF4ENdzNYqkoiakGCJeXbzCPzYV7HcjUqBSZ3vCwBjS
6+orWHMvZoK1uSMisb5kn7eNSNcQHlwa/Qru2qZLwUMgh46rE3E8dxdVlJ4XxhOg
aJxUPla5WWBZ4tknhjpc80gJ/WtuYWv/V6ft6UdLd60loaX8EkiqoUOdUg6SKvc2
iaBhds5c4qkjcBl0Vk4/xxDerED2On7X5VNqaH7R9aUM98HCu9LUOUvP1bB4Jyzg
ewFmT0TwenEb2TbrOJKcHEoqfo2i0jBn4ZcChzscodECJAZGHrkP+BVvRZSGWTUV
231y9Z6Ii9vknxNTknN4RmC7iPirxxCDzTGf0F3fiOB2nT7teCpUrLXNhUUrx154
p7Vqx0me2flBzcVIk+6oJgRtPWKe7t+Xt/XpLAd2KAvEQlAhV6UfvM3Jqff7uAhS
mDUJDpAG6SATwWnYiySZ10ol0aIWv/Y6RPt8cybfSUuIDoOYakV6aJ9Ds5AcIj1h
xJHVRHdAGvGJvD4ElI1vX4gUHb1LZa6DISwYoqb0mhVaoWBj+Sn7k5+pTPix027c
YN1sQ+3N3imfaqqm9qIIfofjyaVhs9PHt5VvxmAfZT0m1BDkqvkMOa+jcOOkYmhm
v8NzSqzKITbv81qX1FswgD97MmV5/vM9j/vB9RHzG7bCANLPgbjnv3NWdAPHKXUo
I21PrApswFy2hlWZhV9tqfqNaSc1x3QRY95Q2V1thFRgybP/4IpikJEGCJ76gc9s
8QLayo/PT9196++DT6mfHFJwv2muU4T5y9Kcnh5bj2oBPOTzF95fI/4By3r08QR8
Zo0nv6qDncARIuKsEYjmhMHCJPJfFu6TPnUcBgRSbYGzoaYXQ9YKQ2MhOuLmV2mx
1GWuX4GsNkx2POq3bBvrGhKjjNLwuFBi6ZqgsW3LWhtv4ZJ1R2qeDMZrRPlv4oFb
fmLHQE5rGBJV08cvOadbQamzhPmU3gO3DVmWpn3QLyhEJMx8yUDmeyd4Vyp5T/Kk
CVLanFzOfFm/LSMCn4boMzDTnd/TeS1MfSLf9tBtHlx/LeaogZnYv4FYuNSx0QDs
S08tC8dkndgiePBryzElN54TR6XXfTBxvJK+Vv7bSirZJFIzi8wUdjr/q9o5rR/x
Ht4B2A9AeDjXuAfY7OrvACRBJoxgl8FZpocujC08j28g1RmU/sS+DFitRx1gswax
CbZyHZN48CugE6+t3tc6JCuXUW8iYNRWumGxoSX8/zJUQP3xvTPrNmbLANXmCE3Z
CBO3XysAxzbUwIImJ/QLsnitpFb9PzYJtG2wi+2KXlurkdUxHL7uFeNw/vpT1n2o
XWczIO1KbbPeIjOQzQWqdFkZtKqmnZA3hce+lKAXozQ6liCY4w2AmDDbMJ9ac8yZ
MtI1wfyOXTs7sg8Hjmdppt49nnWsMurIgQDlwTojUfNhMH992fIzb7cqCo8G7QfE
b0VKNBM/UBh6MC3mndFLEMith86MM/gzTOY/+GsKK+7mUbEMYaIELF4OKraDzx/+
QbG+e6IDR7fEJmIrm6NODV3ZqvbS+3rJdhrXmFOTXcDc+H7SA9K6tk+XqFVnFSWK
ajOGTzwmq00c4yxTusKlJhUhkohr5TDo/I0pht+I5wtI//o8dU87NlrDIqT1HaB7
IZTTvdgzHTOKwb3TrON+HrVhKy8/IxnvFpz30hsh1KeWqvv26MEh3k47rt9SmKDt
Erkgnj1BiX7yGltF3MdSJ/1ETU/dAT8rHUnYwGexPGMlCS6epBuYy1Iznb/QxtU+
TvnLJQiGkXzhwRZTCXKhu1F9GuvEsSaOTBIXsgiCzUixg6H+UTA8rZTa/TYk36rL
prVxE4BqrqNsMdiaqeqMbsC1uubfLUYu0WCmNJAfl2jC28zYUd0LI6EDGx1wfiOE
nH5sXs0yRaN9ESfzAvf3BGyntOcla39bO4/fr+vLB0YX0gvigyStFYPysdVdwd0d
GHe34WLM81FKlrbX0eKwx0rXxXcX+T9wbukchWUtIEtsi5tywFt+1qqgGPdnC2Wo
vRR6YX6JaN51AkwcT/SSePz2oVN5v2EZ3+XEvOwgsC7EScf2A0NrPFi8PgDmdvnM
46KB3uPEnt1cG/hRLyhYJUS9DPSSA2USxjCWyMS5k5ReESWdIKoLlzSSDQ9AEkQJ
XEdA8DVefjIR/R/aNekASKg3mDz1D24vgI/JeqwQOb5MtLaqKOT10Frq4tB/bapL
Xtoo8VvBlo0R7JMk84AG0spBGqB3oMS8h2Ih2fcwrZpdEDUsKY0zf36cHIUCPLXK
OjZolPWHuROTzoKbdEI0/4bNfCM2FIKtfpXIhQMnj3B5mT2X6hPiCTedGiL4sJUk
a1PiNLt5v1fY7MDs9ZKvcDBpiaaxoUJx2nUvoAgRvNOzYZM/oYqG14iQdeVno7Ek
hf2gV3HqQK+w5rbuPE49Q2C0Od5I23yBhoDmPrX9gZK2y/ASVq9Vy+Tvt0AEEO9O
B9oJZK2jmGZcyVVY2va5HnavEsH75K0L2n47zz4FC032VhqIbASlkn/ayXgjgjSV
XyvtggRooZnfQj98TCWNuowgJf9JYz5LKYGql6m/umNlmOefNRVnh1Xy/3fABP9v
hqkvQeZK942GeBx4fSVXAKbZHnXRoMdrtgIt/pMPjJnMIqe/fUp32Xwj+mMZfDSz
LGUTIbZ5bJvJnB7CUPepLqnLPE455J3VPfsTbweQbiiNY/cOm6DVjCpWm7JqIWRb
VeU9MXWfCBHaZfbaVQhQp8ZbfEeFLYhSVXCzscZATJ7RnrV02G/COPezBgzhR7lH
WzmttOqkJwE4KFwayuGTRHoA3Gl06HAhNjQIRc8nec8nj9olnPrWWcduBdx2yqux
w/WP9Wgx37nNDkPXuCesH10RS4PrLBCETGUB6nSv5NyECc+DEVvWuX75Q1ddB2SA
KjP/mrBqYes0R4OzETJuKc3uf0oSA0qRm8N0q6iq6AEpR3QOluR2ZVipAA3UDqDM
RYeE0XS0584WA4kwwlC3+XZWS1ER0vJNiKp72KUA1BOnxJSaDSopCp5zZkhVtf+g
M+P4mvgh3S1jQ5kogDUPWu4OpVqRE+nPpeTYNABDXkisza72d5oz9Bt4XqDHBDmN
KxrUtc2wFPWF1/4zyhW/flJuN4+AdLj2ZAPxWsbzKjri51UQV802Yc6FNqw9MFBY
HczsuCYRsG8w9ZhvuNrfc8rsQhjloHKYd9YaBH9Hlj1uHzqId+FHofRSAK+pkOPC
XBj/iA9kP9teADX5ikN2WOQJYo+RC5HUYlQ2fE284kVc0dhf9Wwgy2G4i3BQyyWx
V2PgYh8EblK4TQuEJNLJSkWYhWr6qPE4tb14U/+BLboCkYloMgE5TcV5lGqNzWzR
2AR9oRm3Ce0uAHM1peWdI96Q21fzBlQ2CPxRxLFJReGmDZ3Gt/3Ikys6FUQDiMJY
3sAkn3elPZ6kpdNbtLBJnHbLgS2fili8dY5/iBfLA3zRanLbUUfJgwWzcVAMQpgn
JJsCuJL55II8yDTifidickd2fHv/3Gb1yQeBT2xGPeuNBsngAm1eTDZ0HtIwrIBh
+yh4mAsJ98c6B8+Zj8EcHICOrCmDQPO1iA9JYyuzEPJIZkOUvTR5qAeZQGLyS1S4
7wINWWtdU1q44upNcRFaULpEXj2/Ye5c/2IhZq/LuBZOhzNVUZdR7oa/AgdLvPSU
U0T3Uby7B+3RIEcbox4AjDtO/TRi+2D3AVJDGqWnpmU5gY1ATCBAXkQRkJpak6oJ
XwcqJBRaTSCtHziHNUoUi9OvQoTmF+cp0iicFXuO1kQfwjtjhR+WbWpVNkFNLoLZ
2Dia7ELIPW9J2FYwV78XcurfF0/r5mDxJdV4XMW0V0HdTRkPijq3xjS8mi42rSCP
rcxgoBo8c84hw2Op5cOrEUkxPMAdplJzL8VZBgCiJKYIxKM/4ElMny7Vlid+htB3
BWKSta+GAWiZUDhUv3tj4Cqsv4n5nO//PVrig8KWj6cHiX18yl7GH8G/4ONAQCRh
hkbDm05oekM96i3/nQ/uq4+g8G0NsNFHjw57Hgj90G9TMi1OBdqxr5zLTkVn3ES6
k2mxZsKyeNaonwvkBGuAJ7z6Ps9i6/zZVRBzQ0PwL0f/PBzg+W4gbZSh+qScd479
PXyMAUjaI2RkbPeIV5fhWRl5yregcxh0ISyG9HYjCmKAtaG1+hqG+UGs5vdDw+xL
jvSlGOPf0qIIOjpoY00LvTL/wJKnoLjC7WRKVdLoPTojbw2hGWzVx8kkIvp6lTGd
z8pIwnfh7TMXviOwHD8ESzZZc2dAZuTXxN+j7pI/vavoY9Qvh6BcrguJFxnB6Xrm
q6AWklniMgajh3Xgi9XEaQfJc/7Ci/7bpe6wy4w13O2pj7NgPwxQDzvXQckmnewY
yFmR4PeOErUnEMYo0SEFbyC0vjiehFrU66Xy4hvBFDYJGo8sQ481yufCnu07ArDI
TGnjspszepzJl0w65uty2caEWMSHq7PEskG9iL9YXj/IP/2grjn+kq7GJxlj88h7
GdZCHca2CbRLcYxPbcHUJnBuYG2fnZndhX7jiYhsioQQjPN1CGxAHMQ363mLPqrq
yPQlxGAF2eReZSA0jMpRfn7nLIjJT8FtzWQ3IuAoyZPrTpXdRtthlvAUv2Il6Qqb
2onIWP/T1GSRLJYAkDCR/RDyq0fBSo/blOhjMgJnFrqgo99q7My9Ft5qH8aqjKSF
OuiARUyMVhmZUWBUz6UKFwi+F/4iYx2eSmvmNVRUnV0F6Z9OF1XySGsFtyeE2+i2
vXtsCPGB+UA44veBiJv+5FLsMwwuGCQJoyJ95gCKO3FkTP3oxrNfZc0S9YHkntNW
QLMAHQ2Pq6vgXum7xm76Ye2rrfyN9LUi1ENxkuj+D7FM+xcUg4OjooXhzOugYYoH
cX1vd5PAoEr8uhneR8kxtVMR9rZUPGaNucldJtCRRZKqd4RB190C2HWGiTuP6Qvo
rQGNq9xizzo7glcTraWzdUzKFagBVtHt9H7Wwl2T9j3CZ50ZBHDLXrQOOiBV3Oa4
UxnfQvlFiELYqukCD9yfX48qijpVP160xsMpbq5g2DooOLRMcvkwqpN7HBWl0XdH
uvJ7ZaWYZJ+5qkqWxFW1sJ4BzIIIpi/J27kwMYHN1x/rncfurklejOaGBqMdAQjL
Y+lzXy5Y4SnANqky+eAyXr+72MlVAr0NYHgn4iuF39iSOfyP9mqhIJZXfK5XlSwW
I0DzXciA+9IQkx2JOnOA88PiIoYCMCuS8EClHPjQ6Hh9AfBYDXe98VtEnUB+MUUg
JJKoMltLNxVf+NMP03fKy7LzqQGt+YThsO/Ysx+pDoWAyt6R8JA8tpocGHnV15B/
JqM6lAg2niEYqfOlhUiZrFcwuz38+4DQj/313zAUhtfKkf1Nsw0i1ZoYrd1BVhmi
i0Lt8WJg6B7xl9UXStTyfeKVkyDdo+acUBDQZRJ1AQhIIh5ls7CHv8evCAQrOcWS
7SbTrVcmGyxR4DB0Amkn40OtrlwqpJO/znnNJ4rxIBkyKltlFAXusS775qI+ArhL
XGJGe7We+qhH9+8fp7UbcSUQ8mTqbM+L83csyxe/CAFaYLa4kHRZZ9RvWFJ/Fj+g
hvUgea+aRKYG0graBX8dQ2pOtTcX1TTKgd5tfep4vqCM73tlKLKhkmYUCMiiMMwW
CEYbYFyoze29j1QDT3AmsPiBXO490ItbeXNS+HrnXtHY/MWnT8g5aa/VKyYF7FyG
49xYOBkPA9CucZVxThC0wEgvstaEY1Mputcn1by31TUlXSdglGvpO9TR0y/0PZut
CN6hIsZSaRjAamgHnb91792h7V/idGxsduOP1TKUsWTQGyy0mI8zH+uxAkHUtMEG
qLNXMKSkEAz+/0Z5yXy+jaSUnFsz0Ur41cIIA9GJZm1EaioMU875+x5g6CLQ7L8M
p9bcncD09vGp+/z6tqQsxgBkKJqdlByfRdArSaM1iZ+KOCMHtTNE9HiKJLhfC9ds
BbKVh/vlgBK4ht0p6ycf9n5oSv/TgO+hJMJMp/OBrWTgSVQ0pmFCc6/4XGcVuRKV
tpeWDz6gp4HPBt9s1+a5GmBU6vYYglMBcyLUcdDsAfXVnOklaPnlOT8lYbC6+zIJ
0dRnYLy+NJ5jrvbR+J+ftiPoK/oOIuGwQtCySh8pFhnw7aqfY8eLnWdaeWNJsmhj
kxi2uLEHTV7bgz+au4pa4uVRiNvA3faFFOgup4l8WmX0rOXppc3hNnwlZj7tQiFi
dyLYXjpj7aVGvsWToH9URWwZvsYnb9JanufmnTW7PFwUq4lhFAsTOOiynpJj0EVG
x009uxUSpoFvZfvLDbGq96vJBmc8yCltMADdDEMWxcGFIYgJogaBOs/MK3HYQDwl
fksG41K/OWXZREbkhBuMIGBujN03a9L09XJkMClPV8QgL6+S+u8jnYYRZBUHFleV
9wayYIuU2luwJa5A/FOK4Q3xJP02V3rYBIK+iGaA8lrtiME4kBMeWm5tfUSLo7ke
AlLAo3anQEJjI7+7V/6p5UVz1N0Q/e8LSlRKHufHki+7tzvDhNpz+aLvJQf64+7h
KIExa8pnbg8X9AYtb4S4x9H/eU9hucWFBddDpxEtchHat9miwPVuXHcB4ugfTryY
w2WA/hCoiTztqW47vn+FRVtLByDjvRpS5sym1CZphfqtZ0d2xnfxj9M/hmS51T1j
mESia/e90HAtgskkg70vcxq03WEXfT4/lNBeChsSGDb3JfYpCjr3LzF6GmOhQWHw
wOu32LKmpNfTQa/zyNXhcABYYga34z4dxpkKhkushqh1ZThly8DGJgkkeIO/r+Kw
255yYbKoEe7VqT13C5/CohCym7YiW/02jNH1DKSDhsp7fd6n8NSZebhBoZysRDS7
0mt+6TProMSkip0lSdR/snpAuKeY5aKxqODAnYmOlsy8m7yvYRgkvQSungP4R2d7
Jw8momdzbI5Bq49mdAOIA0/aySzue/mB19sn0OyPxFccRSMqI5X6tjpEmTWGNofm
k771IB787kRX0LPrD6x+CaUoY3hsXrp0/YM9nTxiMOMhmV+vICkKWPIfP5N+vXp5
jeJxaU4zXDuzfGda23haDK4Ac9i4DnCT2pMb6DHqFAlwHr3PKggyuQD/E3xpiMbG
C7AOoRlCgNxrbSVaAEHjIcFiO34TxzCPER+k/cPb/hbNf37lsrKzDliYi4Fvltr7
zUKPtWxBPeyMsepVpZHRcSjnsRYChY6dO47/PMP3nZZuquobP6g0owb+e3K2FN88
ZSDtu+Bl//JVtzszSSzJ3WY5YnRSp+cm1aymAb6p4+85mN0PT+NzKyjunf9JHVdb
8/4sfEquDuOfIadD73t3jGowJV02vGn08IYkUbZKf+8bcvz7plTzNfiip80dX00q
ITx6Fa8GRwMnJPT/zN0BLl2+8gY2yFpQtcjLq+seJ4tegCKjDVw3dJqGjayaoBGD
F7ZbhBHBUgJACZ8NqAIhWTFo2Ru6jJsWzvblGVdASNiOkGx494nfnW0Ce4gze9O8
WpFVu35LJ8Q7iBF2/Ndty9SA+nT0gwsWPrBDHtRN0dY7YfjZxD66F8w1NXIsph3j
ZCAJzsm3OYOKmytlkpevShG2qmzwT0G9tUxMRlz+05+8NpC3is93oHiksuu9DN3e
WGOg4WzTnfAG9rz/pcMYtKsqdp9Y8HF2432vMOVR3JolrHPjeC8uMX9Xh33ciqf7
IA7lRMFVXDz5VQivwLOhAWBQfWAmtTXpQx1OCGYEtNZpafUQLynrjzda883sHITZ
bDvExWYXHb2l9ZynS0D115pl03kDz8Sm35WJGYf/z148sBo3g5OeDgo9tiNuapHD
yitRVH/uuIhxzwzFHNueKSvnPPaVOpyMPZ1zKUtxp0C+fWA+lg9/gdkAcrusU6QJ
hOp4rsQGQZwSSLVHOewmRZMjn4ix5jkiqTZlMowCFMFqgrQvjo/TvVn2VoonUv2N
KQGazoqGxNEEFH0RYS/f+Z6PYsyqK23biOjF3fGKcvrcebsozgmNT9b/HLtL8Ivd
A8IzrJTA9wBrMnooLDrG7EiCPci6mLGZDVdbB836pGYXQHklp5FDWuBRY9+JtjHa
3S131xz0Larz/PdAsPdWaq6zYDt+YUpNAxrTFpGCfx9wXAi3FRrrg8+r7pU/t+9B
wESLd57A1Y51FzIM+FaD0kEcCWBQXLAprcWHMrKF332xBcbiNt384692w9C+ba9i
Bz319SCg8C7Dgul7UPdUgqPlLSXYKm7lqje2aIgvggUAW3Kguf2t5ppUExp1USNO
2xGBXDf5TuPIs19es7VTArpVR9UhJDY3BBMhRzObu3NbWiVn2Qd0boRxvK352KDO
BU3FHWvnrBI3GhTsOCHkzWMVHUz7RL75KinZinP6tH0VAOVBMoHZk2SKbG4ZfFrK
J0m7IdBAfIxfbU4MQJKIsikEEmH0GQltuYWjUjFy4YhP2PaRtmhb/JOZmMUKYYIp
RQx9m1csiq8gdLJbGUkKR+oXczUx9/FxfuPKuENwkyKcPbSH3+IZJgp6ScM1SJu5
j3KW1tq0KldsRF0Vc6nLc56QTdJSmiUb8QdFv0sfjnM7T1SIQoWRtsuN7TdKcmCT
W+kWxtMdRmf4IwZR+cLU/nLN3aup2iCLjqXxmrLfUMZscQRitKUnC1Zm+qlZ/wTr
sLreW/y/vAtpZxDwjGTaKLtjaVR1f9Un/9E/qDccOKFNoXTPpcyxLFo5o8glV5mN
Iu+1oMk65vXy9/QiUno1CNKGVv71deXaJfxSro7QhXzeD3XGtW6KKVhq93979MCe
zA2EIQtDB/XyywJp6d5624MtPelHq3IRV01N1PmQsM6VVcX1YuSuq1TPLZjS10DY
8WuHwdhGZVWSqcQjlfK2Lt7+8+7Lmp0vx4dmUi8CtciKpKBhEkqnjMVNn+DVqtoI
FslIIQwhvXthXblWJOg35KS7CvQpAsUcRv9TfR/jnY0lhY8mTVwbbKk7B/PqQM9g
ZoTkAArz8hixrgGRSC5L+MnFAwiiMKjuE4soAJzR7CHw93pdeAlfJ42BIArVrLI1
ceQx7PYQ+L/KB4X+oZSFxyROLOI6jH8o6ZG801Ze3UT0UNQ9/LUhc4Go68p1xu6U
Rzte6r+s6XolptaHnXGgjiJMFHe1dv4RAriPYkrm+uc2VNrJU27XZ0QdS8baI5FB
RKAY9HWOQ+EHr9VrE7IFn2zROhKE+iW7CF+EEqJ5hU9zpN5EPokvcdh6VwIxPL41
kRPHl0Vg+JL11Yn1A5LBP50JDhXU2tq/UD1UBwTQ3f0N4eITJHf+XT77ATR1dIhT
yMhPVDD66+X8gmihWtjAEuvZWAvtgKk1gM56y3P89osFcxOs093dFlEaMNTVMJv0
KkGzaBwuBWoLqzuQUyd+GlrEuySGU58jTpd4HGwhshNWH4Go4LcdpzIJPfj/O9Zc
WSTGLP4lqKveAGkb6MWv0MU7xe0xLZvaUoML+VANPH2C3ZVtvUoKR4ubaeYwx0lo
bSR/SOuAswZVA236sTDCBp9XhVxwyJ1f8dwiM+Dut7fW64XVY4JkfA2yWE8KLdtI
FkL2PbfIH+uAA/wCQf0fZQT8UUwPtQpRF6joq+K2WPnMrKVpFGVGIkuoYw3fMzTx
p+5H8zxVUsair7gHhDPwb5X9JN17QI4i6pQT8XJvCla4szlS32s2ou+iKoMRC9hV
0hoAXlcD+W97KNXRfikhy7ReK5jzp5O0Hp1TdnqRMfu8NDxODjQQQsYsoYvNu6In
I7577ftNp6yiCUDMErvblPPK5CbwWdfxl122T9l/qIRIDcvjtCju8nY69p1augcj
0mRCfw3J69w4mOPmZtvhicvba1/skzmFBd7JewGvc588ac4bgEthpZims9XS2nKn
u1cgaD0+AvA6cnqIPajuJYqdxIVYUwTF8PUIioE5ffDXNHMgoskmG5ANVOxNl8xn
6z1ENFXDXNgkcp2LFVCxI+nZJIb1SSTrnks+fqAUFgOXr5x84sOzhfb0H+ZEjih7
VtWIt5y2T67d8qoeg1+iHkdPCG+Ha7cn4UAti44QhCG8pADXx8JGde17ZGJZcnln
FPtAd2fZ0F57RoLKpVfZXYZxuFknkjtbR9KEr7thJvj21mMUtAtttIaTABpcZu09
Ds1y1oaaIAXdGcberbmDGpd2dZ5IBFj71X8MZNOyHKBTsolv1hrG6NaE8lpquKjh
2OytcF4n4JQ2o5ES2GHs4ExwWwy97Jahbdn50W2zjLrG1NzQVZA5LLFtgmurvS6w
8j6P61N4aGaPlzbjQWMVSAzqd4T3cF6oOVAvOw0OHO28IACWc0NmzlstIJPxe9p2
37kSdqbibB7yj18Ib1oX33hs4E1vdx0qMYOb/JKImI7h8OH0SJsVszcscKMahwGk
e2tNli2W1/VruW3ribsJOG87fkKR/oozp0o6deS7oNvFxh2P3/ckDR8sxRmDixQk
p7msXYZLFxQrBc+7C+NeZByApVqWUSq0LFyDn25R3t+SUSN53T1OhRL/PxqHhR26
ihSdVaZa5cR+/MNi5smFNNKe1JrmTSH8lf8oM5lWOMaDCAS/GyjcLONaNVEc4hTA
ONdN/3CNH0vIlEQXSorO1J+8eWLHhXK7P9mBeEZvdR0Fnv9G8bk3MGkOk7A3+g0+
IObVns4JNLPzaE5Bn1aC4NQI6wAnqwOVVePhzpp8tGt+bniQNaHF+5hB2RT8Vudb
HkxssZLOiTDQHIMdkbTMhv1deueYVcinpJuuA/nW0PTEIugVbTHN/oHnxev78xp9
4rJyBHrgPHjgXUrBJqvcP6dprpyCz324olh+b7To99Cs7CTg8IgDRhTwK4PXaPZd
hTL+rBE4VOS0wrx35esjR/xJK2aEgl+CQzdOlUQ8iHEO0DyRV32vMdSrYpLfzYjT
/gpkAli/9IM5DgyvtJXm/Xo9h4dakV49d5KvsFt3r3PWlieiBsrysLYajEKtluc/
2p1m8CJkp4VihcB4v7wjGsgQGqRpNCrwndKbOAUZTrNIhf5E1eCpdIgAgxDnfzbj
J11Z2gNYxto/TZwCIwWtHT3zl/G/VEksn1hVPew4EV1VH98V0mygXRC4olA0S8Qw
qCb5FNzwJ8lNA+5/sC+LPcyG6lodp+TIoLXHDiNhLLYkjdGjkcnEE941h7u6pACw
TSW64ZK68BjG67LTBX+KcKFaprR2MAHuVM6ofsnyb7m3cUlicQ6C3HriUoc+TIKO
tmMyIDL8Lydi/hL5NOZAJSXwP+AM13zH8yqLv5O0KTfFPkQz5AwEuYO6wPXY8cFR
mc8X/mewEV9UmAhUsZ5rYW/i7bX7dx5OTpnQHR5X+6Y4pJG+sdTRB46ydS1CuMYY
pIw7pliI04HCfRVK6vYbhGTJj9afcuGiU5Mt+kNYYysDHyAC35q/8fbljlXmjLDk
GP6X4KRN5m0CSQh5jMfJBtPPvFvpirjIKq5qPJZ7kvUTqEbTJzZQmj6pMlO+stQ7
TyrH4iV7bZm6peuTYKSSCn8czTzrxROw0kgwrCyS+wwEFJoXcDpr6LuUTAZ4A38s
9+p5j/SQhonZCqOziiPK/bYkTP9axInoWBzJAZ0/uG3KLgNR24Tr6ib4c5agucVW
mNA4fh1QHph+MKmfeup+vLCZ/JXJoW/jV82vneeUq7CZ3evmKtorLEpbVx7t4oz5
S9uZTP+8XvHJrFp6QCYf9j853T0Yu0k+KFMSMVtS0sWIQH20hYyT7pisWNYzL3bX
K3YAlykaJkxCb+wA4J2tceZRmN+U+bMY44W/VkvrFRjbXB89PrYm9NR/HcGHC/Gc
fEe1jfyS2KoBoi74D0squcHzkEFC0RcwLWPrTJojkT7LwPItQE7Pc8UhZ51LZ/5U
vMyeYX+lq8sno0Q3YC7/8C7tqgLLYzz+s9CtQ1tdnhvcEdEG21kj5rKImYEMwans
jNIz5mJxFRvtjAwI2OPhXO30mq0/cAA75PTmGAks7/CmE188xmgV3drqBD0LxXbW
7tcnxKuvfWlUonrbqFDMXe73qlsZ6UwC0Y44MNgLNtZvOspagGBZ098LmsgtEslA
QRZZ/jE0rrt4yjtfpkrhNc9q7EeiMgPWs9qFNsJkB6HrKJFqvBerm1SDhLBfmdjM
WyjVP4Ow0u8Z9aGfvpdVcQQSVswynfiM/CcpIFd5zD+CVzEbD2YEvGJ7TG09xYRo
yU1jxbxPsPTVNJ9PP3YzAqcNQKnDmgIlDd766cd1OoUyKauxIOtQRF65rYV9/Lqv
LuLWON6GLAocDw+wswOaSol6US2jyHQqo4uxxRw3QmiPGGJA88TavWYlh1C3Gtuw
ZCuVU9DYKi4JWrx+pBb/ZTdM0nRJTPJbs+v5Fr+/DGeQsWdmwDT8CCRy4yKh+2V6
h0EyYgxo/UXaaOU5N/3UdXWdd6Xr6qtAFHRJ/uvAQ/jpvH2XR+3HfLFsR5rXNv0E
PvHgnHMzxDMLKzkz8UktrmUiuw5BPDsivXzxDScIxcW2MC5svMtJXgAUsfaR6UhN
L1whg4UgxYZQ32mC/J6d+aXW38v2YfmO7U4s+APgJwBo2zrkahGHfF8QSLXmAT3y
9BgV4qyNzOfxDRyrnFReDorcctLHfRH01ZfSjpedTP2HqPT6HcMxyGLzR4piKoLA
WZkMwdvig1/Dsl4y42MxOjWUJEGhfvQuF/NXF7jhykFfQbGdSMQitj+0vajR8UUI
9feMahIvToUwIj533pOZqIljvX5dtsRJ5SS/X2x2T5aKgdjJ1ULbTZ5HFyFVvjW6
WPmRov5ev+Xc/UIY/A3LEJUzoO25bs4liHpy1nkV9oMeay20TO/v1sVyronnryUs
mYSJjlrlj2FqLZh9rUnTKMSjmpNciYSKZSI0DJHkPhCU4xBBB3mF1Ic4UUFh2/zd
fOvpv6Rn69q969HmJ2wpSKRITHErfyyOPo9rnR/vnd5pFVQOcHMKxbmJKO4l4Ziu
gYgyem8l+ugqSWf+mom/5aas+1GVKJUlJHGrAfKceTWcZlrL+/kCPYXeubeeORJR
WQ8bLR48JQgvSW6Ktz+7cpf1BQOvil1sPjNhxRPNeExJNjKKWiBKqLEFWlFwTmaf
+OQ52MpkJSZk3zg/j2JKdi0JOlU7nMYD+x2ztR5K80lQ3ySfWcQdSvJ4RXQ30ZYi
ExQ/hZMDtJ5EO0YgukHXuJxM4ncqjil9oMM5kv6Pi+CJAwDYBkOhVc2N4ym+vrGz
XgL7VZMCpZDGnP0UmnZuOZfzT6ILbRGdX2r34v1lLkW6dh9upDdFfalF9LyhVdTA
lDWI3pBkUJKibYgPX+7xMAqUYIW1ynJQQ0KxwRFs26skKlYKagNB/wai9zL43CE7
s5Nrv2O5qiK5HNzRJJtg+Shwbj9l063+N5sk3TWNJAIOPsTOF0JZzk25621EtS6H
ZHimilZdvgvw2/sAOOWwERa2La8syfoiS6O34v4x5aLHmQNtr92WG4FayXwbUmKL
NSuBrd9SUVSHt6YLLm8LZhkgcaysLFozRUc+mrVvjSxTEswBcn/Ufko16LJVTlo7
cRPnh9yrYGdrs+wiOuqjTbnniqxa2TFmSrZlGIEHQu6g9D6UgWXB8XDwhnqPhbHx
phl4NhMhqhI4oNoESPm0sTXlqklbkfDQ9TMVrawDOe4gHmgOumGEPLwP2AWS7hua
oy13gPv9nPZDiVZCKGuWHeHDfR97MiD6ocaKFEUVKj1310e+67zokRokx5G4UC0r
DHc+1p4c3ZRDjtHUczDSQQA4jQ+9B6r5woagOSnf2pp+bZYr6qkEWnKpimi1yfEL
yzqlDzQPjIjMpwmDLUE3j53alLSOPqLyLlQMV0duLYKK7Ml+xki+RbCjjizwAE4S
bG3BS3f1cI70yedONNL/PiJnWyWNz3ApDJKeBpVRswed3hJWgpUGEkdj8VxWVWLP
Bnlg3FW0n1p2MHEhGlLnxEmYEzn57ldqAinIRnv8P1wCWmRziomS8KpOWY5mVkiI
gpfLTzTxaG9dOJEQNSYf9OBn76i4WIlxIjNKhx1NiMjONIQPiohIf/sj6nD0SxkW
FJv+93Fhl0+41vnOqBbK7GlLJ1fhusfMyzEuE692/saUD6NcQUeOurPO/wEBNzU5
cJlPUe/bytzxa2JX5O9K2oSWsuhV1sMl3L58ikt9+q0bU3Z5PBf9b8cWQFDt9snJ
Fa6IKsuiVe9ezmDURMoP3Ci1hrhZfvFp/fuz8D0h0KETpyF/qTC/kbJ0wegko+SP
tH+BEF2Bzrf6U+ruz/XdZkUC9l8vkKzU87ExvTl2d3TAiMt79ryV7PiG9+9fzvzH
sUWa/QVe2feCWodRTkv5RisrDSWXhmrXk3D7eoh1uY5Pub/ZePCPZSWlD2PJz80Z
BnRroDmVSNYgDYVGjEoObfyeBCbzX3VwoUx5lMmnuBQzi+TQvDX0byhd671v0/Pq
BP4oVCcrDofrrDOMUqOSk1R9+PE8MhJfGM4MY6Xmj05A0m15byIzkFDhYvpjsKni
l9+BlYXunY/ZEMaxAh7aPyHwc6/9sotKt64Q6bdFBau9rHJKClSakMoetK57JDpH
GNUkhj7q8pnI2oHA9pFtr+IG9sjSz6lAG7+WK8wgH5MVEVIQ9GIk+lGcwAFUlpqr
GC+LsWdYK0+jKo+Zj+QZuvSo8KoX8EnX1qXqV0G9+EWDXy9eM11dHfP5bwfpmOoq
u3rqrxVjqpg7FIgOUazHQqLo5nsxPABqRYc1KWQRKJEDgBOiOjt3RalKxeF2i5rl
hbuqbgYyBlfrRV8ludS2Hzn+tJFJuN9TLx5bQWtbdTQCAyJjTNFS9ZKFgoYvW1Xm
lF/82SOSQ3NT0HHpETk/7m3+/TX3iiQwjfEe+IBWNaqqKsdWZVf7AJUr8PxkS5N2
aTnpjEU2e6h8Q5TWFWsnwVshhZ+F/OemhMFQOSZpLv5CVPviv+Dmj8eyVw/KKV2y
iAsVzZMRBpwGZl8YsAkK01ga4TZaDT2PKvHs/4MtiNmicTzj8UQP/nGcFLNAXApw
vvirAbTkpTAlm8gZaBVSUfcKOdRhb5h90mXiwSe8GfzCngmeYFUY06SUdVGZ5wo8
jUeutXz1DxSZiqjikWGAhDTjBL2058PEYDIG73Lv1xq265ePKAfWVA03ngoSIOyv
GHLq6KiF3wqh0jchvLIcByCJecUQHCwJwfTG0MTt62VhWIUTI1c6Agc4yAKnuyDe
QSeokNsu9hr5YwxUzcHRLr58NsdAlBA8Qa/gG97zb5y4VgjhE6tpGIXobauM24Dp
YUoe0jQmBRKLfxhd0EJelJBmOgzhdK/nKv7i6/0dCZWFXg2iAJVK9Qmyjjr04Jex
DRUT79FkeTrzfYopgO8Mg/RPk85owx4FiNE0f7Zw4/CZ/UV0iLR2Zs3V4nKcje0x
mxygh+RKpLFTSjWlTTsucpwu3fRbCLmiXi93OPZhBOIwwuueR8gYF2V3ejqL59UJ
YEGEvlPDckDVQUeFj9oSB292kD4paO3sn2FCoDWslGS+Q2Pd7opzy0W1m+z9nj36
52TG7etGBKWXOc8S0inV+PqzkGAXDngdg1ksIA7NttQ5oNg0HfWfAO1KW56WJqFE
KqnYfYe+jyuek8kpbqvY8D9NyR2hzKkEQmb+WvSlHW3ZKDZ0LyZ+2ajdJiHOFqhn
LBG3oR+oMu7pM0tV5J5Ydv7r1PIhGbVUo+4cGSqTm6BvCY8+/4j7Y6lMw/MJFbjF
P2MlpwpUQ20IY5Pmd/wWpxYmpSpT7i/6X/uJQadS2ZIW6Whsp1mtrfTtkBVglznD
W5AtW0RGdp3BYf9s0V9U37877BedihWz7HE3tlF9rq7mKthuRvBPRTBy74AylHkg
V3N+cPVoNsjfXDmFjEDRSmNKcdeNf7WGRqZ2aDj05FN/FnNdZS+ezpfX8t80/q3A
umr7UfTvHgT9S/9yMKIr0FfzuCD5RGcpopNfutqVdfz2WCKSeftzGf+xMI+LbPaz
ZuJL7Amj5mcuaYnmmCYWFvTAGklbp+nkxqn5yoZZyQoF4A/Pz3aLk/GCIB3hZHu+
2iyLv0lxkjmCFTwitMLbtbbtocG/YxgHrjvTYKPOJuqpxk6AJCwq1s4GmnOjIqKy
1IDEOjtP3JlDkg+3JXc+MYQPXT3m5xJXB46YPKWrHIG8AiSNFevMvAVk8t0AidHG
elcPa7DJMfPIW4s53JNMENz/I8AKcRqltmPEcMxlwndbYpqm0CYDLw8sDVJTGqcO
VLj2hewn5qIGE5/o7cYByf2tUU5Kust7UttRlN8+pQ5PBDF5AxY93R92gs+dD5+I
rbXlN6TztCD2oHJObbH5xiuMg9iQAXXweZmsEXnsUsfmrFOGhFmBCV82HVdBeE+t
z8VhUHHJ+xx6xZIMCWMjx/QwvV3Hq2pIihN3cWZHSWiPAXkrcdxC5rBqi9oo2AGN
GyJ5VsWmZgYafQCVAagDWTi1xaae14NTSiUHpp94meZf6seQss5Oc3UgGBmcyNxB
Ic2b8A11KDFRVMROPPSR4nAEDAEDPExQC7PAw2fInYzewV+lBYOsuvvvt5S+5Ypz
f4cjnRFCvUjnHfcY3ev3YReeUPykSZhscwkfy+QM7Ztm90jwWqgMwY+PZnToCGxg
DXt6kUrUCZ9aniiTyVKk3NfM8PKXDdh+UYifyHXvtGuayxUkcSR0mA4/QrfZQfoU
3wk2QkITNbVfvp/v3dvDV1Z1+ma46eYPb9QfIiWl0VXWrAnsEQRKwG/BuSgdDtqT
RG/sZZQtgQ9zTdRmoS0hXcJjXFSgVGzZdYmvtMYjTKUK9ZFZGc8GWnbROLApYkLN
qTt8mgAxb3bvaM9Q5vkSvZSZ4DTNQRCpT28N58AKIWJAm/ARfGG0oaMeGhNraV8I
NJgDHevq9awgHm9TqBx2K9MEvSu5VNWJnl7sdMaUHuK3bbMxCw7eINoQlIbl/MsG
aSbZLSmF/g8sYU89uHulJdiwB8nhlbfaIG/3PuwaAqfYAfnTT8h+j3V9Fp2+dcHZ
uzS9jYcIFiLRaHYrcK3zKJUX3CYyTw1K4b5kRlekBtLV82YTVzh+FLom7ojNl0U/
i/PPIEoUGV/L1jQUllc8g+aPr/XlUjAJQgDvPqQbs+NTwNq4L5JhBZxvkWIZiBH3
A+DjpGssJSAgreSDfSSVAcHoVFtxko1v/LU6Z555RZDu6p9NkSjrVYGJDMRUeXDA
t2C89Stj0hZg/RffLdQOGaKMluIF6CAlTJ2z/SlSQZcD7Khjb7C9Klrx78zqHQB7
iqbudPrRpc+MznrnkmN+eD9CNs16S9DQ/sYpOickKQ0DVzYpK2ozYBnOoezjYL+p
y2Co86ZMYXOqxfxrAYRtTl/vRueP5nzxQE8Oy9OntsRfO/D8Cb/A4Aa1J8MrF8Mm
IW3bvYlUI9u7+co4CrJarpbWYgLqnFqq++D2jjEQ8XPV7jOKa87IYy11ZRECHZQW
10UyfxPUWpoQvBezJmaLpwtBN4fXrFUTFEz/dmXXAiDReo8/ICXvznQlxTwtT8UB
8s8iCBwwswacBiWBTIcLSVd/YqGacGdCXczYK0w0ELgTkvyhhra/WgIRNMyeuDoB
d7bnLp8PbezywBjDakCXAtuxMZKOM9HCwvVHEd5xoxpWTKBj6LY0HMZE+FyRjfSL
FScqSyqxC4I+fb94flr3uaph0Arg+OWiDD9CR1tTCNJ1Nxptcczhf23F+H4RsBEo
bYdUXT7VX29PvFnqllkVi7IaclVn2HkieKJc233B7QxrecURw7c7i7QV+HLcK0PO
sN7TA69NOZMyYsEqWbyCXqzrI8YD+TTNPAjIk5zNlBnQsvCUmIqe8DsHmDTs8w8Z
Rt0r2MDDJlWptrGCjQ5cySYrrlxS+HQmDqIwU9O3ZHCwHHfQ+efIak7TitUnL+OC
WuzVERu3pw/90xC4lKXRmSwwX0hznrO0+YLL47u/N4J1JHNqbh/YvTldzqx9ccjP
8HzsZeE1bDv9zE2OD/wIR6KdpBFfLbTcKw+vIqAaKMOCPRELCA7Pjz/fssygfCGM
W8f3AdOSx+VoiggCUd4EOUUEYPkjoexthrboQI6+pNWjjK8CLVi7V2gTFgpGppJX
jqGVRcyHjuU9yYUMJDxeDwjEe3w/bGmS8hDNJgOyYGBcS5re7Q5IpghINPfRhai/
sd5Vle9bc8w+ywT6EfPz6xAWhZ/k9PZZ45aW2mDtm8VZm1qMIWuIfMh8mlAqD1ug
42+J21UUz0lwxNO8V1rsCg4+h6b0hkDX9vdO41McfVlSSAFyITMrxnvKXzjotk2l
4YwKE+cNvgB5GBLwT2Hfeksk2bQ6ktx1i5DmNItXWGxhz0z+3k9ijniOKYMw0mjZ
dO4OrbAxnj4iKdJIsMOLwyFZNbx1xjnI/J+tQoMpvi3vAemSQRNy//TPDLSIR7wX
hxwwUQVXnpRzq+5qXhUmvSh1rGxHFRtYW/JOlnIyyE07AaHjGaq9aa/nKctIuIAB
d5STPy1q/hR/cU1AI4HmYu1d4u4rWLfellmYsSKTyJlo2e6BJv8X+EiefGbFcD8X
UWnYlI5Fr2wPL2xNfit/7Awm4Wz25Q/+QYR3L70l3APSqXnNGpc0/QPTXG1k85qC
NqiZsZnBzBHXqaJcffG+QPPbcY+sAwfsH1dHHmzqUJ4HSgYoSfZ9x5ArCx7dGe/Z
MCWeaxSKV+8PTnBNgkbB4CEWueHGc+r8ExDq1dB+9wp9qiW+1mnkzZNWWq7w9UxP
01rIVAfKb3S0Uzj5bqZ7h8v7NsiYl94rXKr4gvfV6hJz5aBibanBorPnuYvu17pb
X8x5+FTGLyrsUKFqvs3/pJyJKjrigDAozi2fBj2q8Ri4wAwN9KK3J/6X7V9AK7UO
MOED4mWs4A91pFW30KCTrNLlzvfjCKaKg7uSjbK7BE7XMSgikABKrjYwzejmbIkd
7Juaa8Kn7XvqXiOmP2+d1Tr3tksxjaYLYeOCWV9/vGSOi3VQwk/A7jfXaitZoA/K
HSaeRAqiLDOg3cApd401hmXLOtUklSIsZykeOFZ9YBklcA/7bNHYrpd++zxUmWPH
Oqg1cs21wCTmgwyzQ0gpof4HN3Nl61GdpF83rOKyRiWPumnfWxDTp9W1Cruw4EHK
WV0wd+OEE4xvjLJCoLtHra3WTyjv1lE536C1IZq/H6t19vV/92e8qgCAPxuOZvW4
i8dK+f77PIfckDHsYrNY1ypelALtGy8EJdO6ES40zNUHGndqZiOtUU4Rduh2zo/3
MFNQzyEpdcZRMIF/2kW4K6TW9gOE3I6BJ6N/JkuPVUjlu1wKlaWKzI2Uvpv5qVAE
R6nicg+SdzepIn1tiKaAodlwRN4bbaAHyri+NFNhWExOvGpaUy93B367tKLnzStR
MZ5TLwkHVRMioyK9N8h18XlcwxbBYpyNKPtDka/SLqBqP4Ah5RS55l1wREg891dd
9p8eikSDTRblp3BhcS7yqKx6e0mmWkwD6TtUb6TNZ5qHgt3ZNcBa5LJ1PBmkQ1sw
i2PmDh5J/4Elc+Fc0lSuShLQLsrK/okr9XJa4yD/LJ1V3pkHW04gPPDN3PXzadoA
awg2wy5IXCIzAoQWV6940aacPAd93ZE+MiMkgyZ6o23OE2aTeTnpeMc0tYodUDc8
jjTeX9Oas+2iW3L6tv1GbRNn0XxIxf0KZquGsuprcY0x34BEO7BQORKe3IQXLdAP
2TfrIGw8Fca8xKtVMBEhbaFKvwqCct6LqNSWrIufBEzxHl0GDLJTQZECFRHpukuT
D1mcd561w7UkbCoTHJ5ENIy462yPoqClY1TjbozYLbxyaEj8GKSis1/ELkr2THPc
ctrqBbDwLlcTb68D50XKlqOFjw0OSk8Fmj6JAx4ZO720wMRVM3DtePhJTEohaIWU
zJbGwV0k+w3vD8HKnnkm8b7B4RWRuhfbtnGeBc76KFWrdzBWiMl4sMBqsdr8FjsG
BnFr2U89w9l8F3j+jW+CA7mMvAgDUFk2gcB2EWC3Swsa2XUTLHZsjw9cIftxA/Z6
KMIFpQi1eMwfLhmysm5S3M1gCgPGIDdTBBpsW0eL9xbwIBrc1tOA/QCgm07bwxCO
ctFo2tRF341SEo7oH61PNkWIgDeySp67w6VvyjwMhF0+0af1eanBSv0a2g73Rett
fA5cQ7Way9YyY+8HJ/J+BnTS9VqSSfvtAqx/wGHjG7cWigIx8OCrEySW+AgENGhF
5HJsIxhCTjN0QEKmOklk4KGjKn/P8KTMBP0JVeqcD5mWmG3GrqMxbeMH7EB3c/pS
jR1JmrcuzethmMTd4mvDT6rwUAn4NZM/V5DuN8SGAzuo5nfb7GO1vUq2o/tZrMaE
MuKA3C7hw8/xgt8wtIC8E63KIhRPpMNofRVM7ZClm9p6k4gynBiXBOD6TwcAfsBe
8cuLId8KALmRO7TleptiKPpfdIBXCOat/CB6q5WhVXf9bMDjxeupW8SLwHnexEBD
jeN/tIVrbF6evMOgPLAk3wTJJA3Ss1iIGTpETJLbOO0/7RMxPOvpYJ0pITrQAFGz
npqxmrpVVvwSnx4gKreunDR6xN+XyonPQI3t2CWgwFVRm7w9WRS3L7t1zCZsgAVC
i+zTgMlxnrwB7hMRF2UN1XGO2MaGwb0Ty/IWaEyTuApLiP57gY1C6OdONs37U9+o
EyP1WxGX6ra4T6F8JiYpXe8WTVigtpHAgi5SS/bxxcNRAKdSSDPwahCSppn4Vx74
1AQxCesDahJ4QKdeBf5nVxqVh+VqhGi5/zPmlIJ4dnfNGvLE0+6Pfy9Hi5iOAZdS
IpetathmjCNI2K5K1IKP2+tY9tIUSWG27eojfwcGrbu0tvNGd35Rc5KFoptSPe88
/7f/SVk+ONtjcdVfNjR8hRqKMNjoDz5jOLgCKw5TaJVJWNJXXfU5Vcmww7NaAG27
hmHcjFDrGT253fusbTC+zDXxIeqYN3PGKHIckKdF9NjJfvonxDwLS0B0rRmzLmRH
PnsFNgGaKSpnP1zUGNhfoRlhINJF8M4YSK4sKo7rn+Yk3wYWf4JasS+0rKNxF7qp
4Ow06gZEMSzWk0C9Dj1ze+ISgiC23panFhEzbaKJ2ND9M3OTOquEJiRzXUNm3bEU
c2FaEwJ/eBDAoP9FJ2UpRJkVJp38SwNTDjNg9FdzJweNbaaqy5Dfy0mXZUnAgzyl
gNsoHnUjpC97Xs3k5ZFzmhEJb2pjU5jYS4syq2A+prNCvgBgWL0VAtsXM/WB5Qfl
A+W2EKxbl8XIjhx7++stfmzUkOLzydTLtOAT+tXBHhN614C60XjqpE/K3px4dP2j
OX0kNZu3iD7zUNFIdPzCMVPomv98HrVADjEDMrxbRegZ2T9MT2vyXQ7vWXoy4RoM
eSMGNl+7eibgPupfKmSE5LO415n6CsRq3/PjWEw5JrwJkn7TYtem4GLWUHT00Vf8
nARDRpaLcET6Tg0P7rei8aV3RKkPbC7H5LXYCgiNp8okie7XfdHzRUUnGH5f93bD
eeItpI7vSgh0KtplyKfqm9IG642F0U0YU/Ks5vn6shiS6gPqbO85kvi+uAyzo0aO
hj7zwINpfd8AxHj2V1JWXIyK64N/6RTyI/9aovtgwBs7isb1aH2HhaNkcj5tttqM
i8SNkHjStffEtvUW6WCmsNSDKojDaVgiUcg6xkLgeixfTvMpAl9aPGE03Nmzt6dq
kC6YQdiiUs+8z1ARHgFJomJRDEEChy9sbWGIaBMI+h0xUxtOnaAgSMl6eFRNUMba
Ip0Wr4NrjXpVK7YD9FXtjTRd1c0Mb2kKB3nYckz9WPMU17SEPMo6NhT9dc2G493t
lFWAifq5oVoMB+97QEt8aZMlUiFnM1KDxOBIa5B+y5pHiFJ+/docBXflUGFRyLwV
8UAezKIy8/0ppuxS0N1pxHnHQx1SNqFf7bQorkvfKTQlqWFdrVjIuMNIP0fy1tKH
1oSeRI7b2GwreYLSry/JIICOXQ3B4ntN2/2Q8gC2Nv2RnEKQMaEtZqjTIY4rVKpR
mmBgb1H7jhLLqR0ZXt9mbEBTIFjj3nONshaA7ReplJ/kU+3i0dx7fgUQXI4kt0Ma
aWwbZvVeyIVAWiMvH6RZZEAEdBXWgdCBoPcbP4xbjPXYAnFPmtF2gEULManB+8xQ
2RgQNKjU9u/GUqe2GogJ9LTBd8YtQVz88M45wAvTZ4SRTL4gweLF4CRb4Yp2WAVF
VpTA20DNFjs3DYw8mKXs6CUg0DwkLr8yAZSKbrNo2TdVwTO90Lke5AfNDytadsVI
Ho0HV8hU3pfES/9Cm1aCcrvYNT1LRTadMZG4cEYXB+uB1w0eZxlEi1zsy48VjHwD
KpXinjAOwaNiJcQcq9FFyORWAshBaGHGHqi203PGRDmBVWHw9X663T7tn39W1r4v
Z/+wOFBWADChTrjlL9q0lgHsVvLj//buP62hqhGpRpRyZ5xXK5fJ0DjVGPtKP54v
Aku6V2KrMkH1626+BuXdtXEQShqrcQaFNweoU9NtsV6NDv7xZ/V/KYDD6Q0Q8xet
S3Sukp6BR605+xx1Fxq9gtMnmqzdKn3s2crj0XgLw1VUa00DlluGww9OvilQ6IAg
9yQHDPCXAaD+XPeze3pLxYtdnN1aYjPLX5kPUAcn8fxEclsjGREPo7WOi+cx0ivr
8CzjmeATAtOQnqNNiNKcGw+NNL8Ss9FEjEPINRM1uQL+o84Jw4U/9awzCgGu/dtc
GD8vZXwImq0ZJtOxFOt/rVJ+uw3E5N5xMWcERyngKP8G6XTH1P1rnDloLLwNbsP3
iGhwd/mwuGcujdN1LSsFIW6DfJE+kOkocKG5n5K7EPkg7EwaUouGAIMyQGSOdjIs
fxlYyy9A+AD+T9nD5je6RPIBU1Mrzz/WSxqqPC9tNjMdBdkHjMt4PbLgszg8AtcR
1ZfONq+mZ1sXga+YFZU8kF0ldm16Mh5ftlPGtxj4XMJRwpn5IOujps/8JFapixUU
zMQTOQw5IvMjQdEA4w1bV3J3tX1ff4UjlTtSnsSOkJ5R9mP5WXz2F1kNC12CqNHy
WGcOLcgno7w5Pgvj+uuwTQNHNZqqa2zclElcgHP/FQR+oCh1X8lROt7SwK/yg8sz
PATwLQdSiepvx4mzXu2VHuxttO2ywnUdjlUETKzMYLiSxa9N2r1VoErgyj6h6nNc
Fph3CwR8rbulN562WzOXt0dS8BqbIf6fQ1l+Yl48c0Qid6nEXZPCxrpAvy4A0Bha
prC9Z5SbkvRkUw5b/kFi1gF5etL848zAgJ1+ny8zoDag7ZQU0uwR1KlUHExDY7FW
/wByuafZZkh1eRT2TRwXtUNbzSKU1K3w16tsJ34TMXruPMcu+mH/FswyiBKCsQpZ
J44ViihqIWg/UHdUk4K14tmQjD01PvV3IZ94G8ShPjHMa6yWEUqBw4VzPiLCTHOV
Ttf/wPnTyRYg99yPI9SYP4mZ0lJStsyegWDLATk3qGTP+zgPmcLawBROYFa7SU0u
JYAg8EoATCnsS3L35scUHCNiH9wqCpDyfUZvC+iqVY1vdWsd8tkCex1/TBt5Q8m+
C5JykXzMHx/U0aNvlNx2z4XWsmazhfv1U98iDy3aq66qz4Oh1YSEv/y/mscvniJa
vWlH/VsQK/UBZixK450YT1dZwjD4eRaEgO27Ksq0hTBxY385yJlFtnSvLr6MOuuk
HUs0094GmMgp7Q1azDiXmOOdH+LmXUf+FP+qNW829cfRoIgLfc8X5tWROmiOOmip
F/rSRxPWlKKHf9j82IZT+T+A+jsOrYstgm4aNCmXDXXKQFVymthUMYg+GJOwwV7G
HGm337U6vyFkoGAa9AEKw4Z11xoJNsXfG0SzXYf+aE6bm4t0X876Zn2mqgkLBkiY
WZeJMc9Ovus449IBE6/NOTS/KcxPDlOof0JiSi3UV9kAmO6zqL0KA3Ef5BohJv0N
uQc5vJs6VFK78bkuDCfvXgq6kayYB7Rafxtu9Axfhjg8v0cP9ERO3kzF2lq/yQz1
upb/wcn59fE7Jt7LarCbMO5m3UFnrfkLtOi/g7j9Mdr2e7kHdMl9C6h3ekrE5knD
GN8b/0sksHPaihSW+THrLSLM6su1qknX+/K5+QZtqU0F/VfHMlrw+i4XO63xRjH5
Xa6vg276ykyl7H//1XUlPukb3lpUOD9r8s58L6wkYLwI9ZyAE8o1YgmOZ17CI19r
679q7baeGAOeXeqT1vLCr2DOOx2mEVgexlDsAifoWsjXYMVBL3CfTFjcOhGFnRKg
Q64D3naAzIWUsqxMpyaKdqUuWWd7t1CQGe3NoCsdPAijLf3n+REYAf8fa7hjgkN0
y1rsSqYo8b9SmZiUBhDnRmbPpav+uEeqjYnnPuncTl0Mz2CQxvkyr/Cv6/t80gfD
9aIEL7cprcGrm+zZvkPb0W3LMwrSVH50kUwLBwvt2csc0QU709AqKJlFOR7R8hH/
1p+JMbFi5lJQRJB3mKjhJYS9TLQ4Mj821RwwaETsGBCtDjGwXbuA3qgCCDnqG/Bq
fHK6hIlm8RDCN4zL9Jk9wHbH8xYegv+f1fNHsP/Vf6l+AnFGGn+Yg66Ff9h236q4
+ib3Ky66HlpgeANaUyLP+CYSTcjaNOsG8HzCUSlk4oFfqGL3PB8vYSA4O2ASWAa5
4++vgLlHFcCAPaRpORaVTIwSSdmnLbBAsWoln0nzFvOp/9oHw7c8VmF32FCUBMHw
rNwMhjVQH10syIm+Vnq8Y3OSnH73XRnArXW0auyphe6e+bNNlt5s92pMWiLNDTdS
zVGpagX1nwrMq5VSxPyBuDxAQ0anOaoBHzknsi7JUjF0Mp2Lyz6gJjhFwpw8QRiB
NmK4FJmhrLWIgPZYLRLnbU6IO3DKn0QzsiFVe0NC1XKTXEFI+F6i1Nwc6RsGhW83
rzsAHxwxPUtwukBdLwWOZgNGc8FKD/7EiWy81qFm2vLpABcncpA9orA48mPzrlrr
mpGzYH3LaJrC+PQZR/a3NPxg47AdFHdc82TvAEuygtPMDUgmSVMuHKaYpAyGxIek
N6Jqqpn/7U9hdZr7ytTenOAwiupuYnVpMgJf28VbY/q/+/t9P69GPdd7LHxO1y62
AWK1TrnDmXtx2ChPI3IGIgE/92m8G8lyruVd8A3pF/Cte6xCUD/LAHrxTRCzDGSB
pUc/pgUQdqnqEI5rYP7p7BOxKQDviqBSYmnze/THy1fdzJnm6ieQbjFfoNhN0Zf/
OJL4scv/aQRBNqnubs0jGrgtcQGc2hBaxqyqgh9wWeWXYxkt5wOKQiaRRqC1WZP0
xeQS2806+cj5JkZgq4ofkUmTIJnqdZNCVW8PTRmiYUDyO+SbS0plJL/+j+IL1cB/
HDokJMguUuQbg70o/hlBgzYc76yLhnwljRCtbsS+Vx4Nq97KKTr/i8UFm7QRmGgz
nYgUEiRMQjCfBk3A+1HtcujpoFjUc+mGhRKGCqKCiFD8kuXMF4e0ASdlL1P8C1Rs
7md2j9b+hZfsUPENku9Ba3ZFV1yi3FubHz0UA3mxiDJtQsl+SSutA9CoKPj5+35A
UOV11YUFDO3GXmitXC5Xau/xmd3hPAoDCQmgYRe5Oc2ntyumOOvqqBp9W5MY8Ebq
CyD/HKbp3h3G/QpM4XA8uztoYOXcTawGRaVnaG8sg8vVSQ8zmklXKLdtSx4+vGvn
Dw5EUp3jt8BhxD+6j8d72Mfffe5wTUPsR9DFjW3YR1mI5BO7GHTHAAv6gQo6TAxq
O4hJNAme77ioftMCjosS9ux0knEcFw9o7dpZlgHkLLAt+n7IBeFwLsVVG6AaUnnn
doK0wHbG1wghAiVILGC189puT8XZKHzH9+DPwL5mmkow6vvuB0Bc3vXnvuvPXAwr
A4/t+Icxg+lQEQ2fm5E6yOhCzYLMxLMT6P+Ucbu/Adkw3kI2dBdGG8HzulF22BmK
k/Rv0WbZJMHC1H2aq3YTdUefA/TI3F8s+hbx+XJYRuG2KClHkXDnCigOkOY2SOPj
prhMZghn0zGGLwtEFVVqThWW57t2fa7+0JFsCjbs6fl0FBdUM0Qed10b89d4iECH
Wfk6J8hh7JF6cVcKnhpc2M1zpiD7MUIuDd/21I94fWXfRyguE20+97YIsZ2T7/i7
nsyPcOC0Yguot9b1RHSV4q0dFcmW9LQPVJgU/1bnscRxCEoMY9lT6FmhQzPm7CSK
33zM7CPPOyBLvcaL83QO7tIC/N081T+hJjbbCzw+/BydfemHwka5Earo47sNEwMg
7AFQHdnW2RqN/AcyYIJwfViYdxkCd8vFh1/IiM6NE90ZpGQXxJ2RDkfc1QIkUIRl
2en+FnxbPrYE78Y3xkWKpGTzk/c6ylm34LPcsjWS2rFg/Xr24MVLuvDl+VpOnhcY
GzrV46RN575boow5ON0ShbGByEo68Si2lvAER/8Oy3bKQIRTY6yZQPI6FW43mPgJ
lXD8mFvUrnWj/+/wkhcofhiLSvmfBB/DE+w20IWaKNGnYFmi/v3jo4NVOteelmHU
IJfPI57b0W7saSFcAoDHPdV8R7LZpUk+gFwg6EZidU5lePC6qrb449QWFRRR5gNT
mCgBx6yPpTJi7FQNX6E/7HBFhhdptGoWop62qNg2uTbq2BkLtN8hGLFVztk4mKkl
g3mdcE/sH6kbZZHlDYWIJY1JYEmf0dVifJx7KSJ1k3hGqFdW+BezaJkHDXxrC+8H
wB2ghvVbJZl5eV520lzxz7Ot0bx4JblUKQquzyWtgvWtY2F4AqjVzYCgdvIA/Ixr
bDKeBTe2AOmKSV8s5ILHD9wA37UUfbipgleFxwqRcavp3HkWM2vwq1/eTIaeSwMj
jh0t7f/OzEe5WtzVH3DVAGpqsp+bRBfAhTMTagxg9cLYQR1SK9A+DjBBEoLaUrdB
2F/SLAMAw9hykdtUQQJS5hN7/EhA9Cvtas+7JtG25jMd9Zdt9XA4CgCVBaM8LMi+
ZoUbbBVOLUhX53COjWcs2Cirw2Ciguf4GV8M1LMuCn7OhDl7i5v2gsFIfRlGdEcb
IlHgvCEN/D8hnqVJgm0p9DQftdi0eZdhoZfI9JuKPMpfrMsJxe7gCeLR6Atlii6r
VbEzpSJycaT7zOEzE6KoEfiM6TYZTv22XXRQVgJTmUhhPYxhmvZPX8J/M3uL8MJg
2iWP8IYuztW+U09Ogr1nInNFWVVJMWDbzpyh/zHMBE1v5cvyyLPbk82tLHiPT1Wt
j2YifWWvi0w7z/EO76z5kTnRpJLAkkYFv3668oDW5aUIUGSEMp7klOLef1Qxhyqe
jY6Ymzy35p3vTgXM23EurznsfuHrt0YRri2hxAC8IDpHOMWr3XYwj6XkRfcls8MP
IHR329yigGnAYcVK5Bm/rh9QP3u7Sl/TIq/WE1f/Or4UmNplckzcts1wZLzTwgur
SHnRaNz5FXwi6Vn0ZWXZpA2iE2FnItolUTTS7TeucysRG+GQROEl/rbUWEtLzeMH
HGMOt1zUYc0MhDhMUcifh26leFTdBJww675hNZ63z2hO31mK5MGiJ7yKv5cotFfd
SPX4qe3dD+BEbWVBiWf1QLrvT7LPM+vgmQADK6Ss/6AokHnmYx5gSy2jnnyg85ob
zqKY3baZUb/Qv8ckQT7Dwzq5/D2P7kDlqsavYVODxPKrXiiMDiwz6ghVyEMJnHrP
45+qm48Ug1kEgKx7DZNbZZspQjIrd19/unsIBUhQm6xAdzWQCV6HRScye2pa7/uV
LR3SqTFpQh+FsWDdQWfr6O/02ZoTnBL6ntMBz/IsI1GCxjjziq55vijpJF6CmOC3
tnX/BTecrB+BnitobeaVJlEgFjbg14/yksNw7IKopdKrEMOEMLNOVXK6R7clX4Fw
Dvvbo+Ce8Px1sV1ayfnqVkMM1HLqQ1yH0A7Cr6jJdMP7IrJmPdgl0pIKJlTg0QyG
6HYJ/lrLQyT3jv0zA6hPbIn3ETmLINXMK5BJf4CWlHri89F6O5K6ihPH+MebbQTK
pX6D5DvG/tT8o9BvKQEGQeoM0RyowP1wESSrc7iMDqTMD4W0aHp0LFcZmY6C1krT
JKevTu9ZY5pDV6sS8haYqumCgMAs5xBEdE6ob6mWpAdyNbfa5JvQMbCp1/D6VDen
VrrBzzrkTJddtZ5Fq5awN1/XrH+AdlYj5e9CLubhCX+ZVNPbH8zhtT2aYxIHhObf
KpUXyKnasVu2pLUuqOIy+uhIAuZ65+XTbaEHfEbE7JEo2HkKlQeOg2lLmCoTzymA
khkveY/QHVWLDx3kKWSXiiU2kLlgLknAzpasLbgjQY8MMYw7Q5D94MPEgX+lGo5z
FZkNxb2t2GZUwdXac1LIZLAoa4wHJd4zmJ+POUAKZ4dGGdDxR7zwiIbIehQdhOxc
JkBUmslDgtkLtvKQbzm/MPc+kquef4Q/bD3zfkAw45iXSQ39T+igK87kfyRlrUaQ
lFUD0ABkZTR9BoevEHpYVYx8xe/ksS4OHCb3OFUDTv2oBVcNSfrP8LLAtqFE6mM3
iSGSBtbevEsRuIREMj4Y8t33dKoGVqaEnLiMapPtMS7Btkg9dIKeoeKEThhuhBPy
kH3fJCLhkvc2NeNsgg/4s/s6UjuVCySWVS3yYquoi3HswhWNu2ERcqZzBAt//7xI
VbZlCjWO5MBHnBUOhGcldFJpn1QtG9t8fkEfK9hxPf9obMrgVOW7oQl9bVmphmSh
ukHHOrUwS5IINbGNDALBy06zx8MS+E2pp4MNLGdCsADPAa0ZJlo6Ah1zWRm8r2ov
Ow3s6WzBGhR0PpA0exT3qtPLiPVMgvMXbK7wcWBQ21mW5Q2Pz65l0m9g8lSt03s7
A+s6h1v/51YZKE1eI/UnpSzjebfoAyUSXKIij9JihnMG8bMM8HcXMqHUz3FANgbD
l8dgYFWzS5FUkq3DVu7iKNTcCGnPCfGSzQSCGLCDIyR0o59Cbw2rrKjPA0zKgbI1
jJdKBueS6wD6jOzbtfleemD4XMGVd2S0e4dm04IN0k8+0+Ug5pztj+HDVapo9hNB
rKV0mnR6A4Dz+E17ovmxT8FaKKX1QypcQDYVjE4djJw90CW8BO+VQhZrWmMYRmoC
NoALe8t9wkZys+6eKSPV8ec2ODFypGvJv+hFOLSQXkaG2/uBra0giqJoSFxxp2m8
JYi6E58j0cRqUngp3/vGtmeT7pal2dr5g0iI0zqXOhKkpTAgqdfMglSYzePF5EXq
oBi7xtDgXZvp/5D/oQFYFmDG51+opJh6T/T6e6GqAd8IIRdO8eISrmBT3o7hDKSn
Dt4L5WaADgVEBlD9Vo0U/jVSroazveVhkFRpY/GYBgzEZTzh69sPdzNn8FwmmiTe
iZe58uV8Tt29GhkSopQ4QRLIWHzF1mNYcyRLdRzFC8j68/LpiBbsoWzo4eOgftyt
vhTeMD2SWzVF6s9hFUG8X90P88zV75ld84umVMKUyRqeV0qt2lb5ZBO++vGMomEh
oavA5hH9tNV1C7OQ3qNGfrAXf6jnrlDj63v2W6RqeiEXZHqaxjc/twKVchEU+iTJ
1W7GGHpDej28Q4NcRqNi6KMRrQ2lmWOG8u8mRv7yeOS99tLrmLhsZ8bGUrFVZRVV
BbZR6umWJdx4D11VKK7vVIIAOCJet3rU7aDUDIat0gGk0NMzzt1CxX/ZpWwiRn6C
vPh9xE0qch7zKznOPLTQQY9tob77+eVBdknp/Rgg7FLmzsyc2PPkDjqPh61GsNF5
QgfKciAI+WIHa0HAXHwz2rJquh36GJSbcWItHSyX5SEg0vjutnV/hjeZxvvagcXO
ccm4dMpaauWPX7ll3N030kLdjN5baJV/358TcYijpaSu27WDSkCozMwQhSqcrO3y
VN2QUU2WxS4pS1uvx8bYFk4S3O2daOfvjsIqaR9/GT1x+A7sOzDVs2KI3X9pbjF9
03mKoSZdOWuTh72oPIXguwV4LUx5iyVvRnUbE+mHRfSPcjxuSFKtlzmB0pDBub5P
UDHi8MEBYQ30g5aXNyeHh8erOIUrOKVr99SQ4f4PV6ofg5SrKKrzMtKGmq0+HvpM
B9Z/jcbeGvEtmpxCQk5F4kyzSHjbE98vq11ReMioDHOkymss8N0NHDIUZUcT06nL
15JjpNPGoU/OSXW3Inkrjv8NuGRPX+PMzUZTHOxPfL9UKMzqz3RQZ403OMFE8rLN
ty57yr0cvq2x0mLIwq2JKQiIIWpe4CrFsjrnVhHv9tA41DoTmVhYumUsEYWXHCpE
TvxLxArQ2/XpA6yykf2vIsBZeSzJyLK7cpOeH/110Q9PHjnxBGuHQW4I5kUCg77s
RWoitNv4NC7ZHlG5dqdtT5TVLHuueZO48ChSMd12ky23m/wrxOdkU7ljwiIgoWFd
dOi+qrI7tGkCyhmP1Rqgos9caDkpDIuPy5WxlLrJ96r11LNgk4/QpYi38JKnd31+
1TnxdzodCaVQNddqgMAx+DrqfqGzSSCel1oU6EXpbSSEwF+K7MWd9tnK08lOMLa4
gT5wyqYUR+w74JyCQtvIuU1KY5Z91vuHE3npqWCl/XdiZ0LWM5Reia2agT6BzeVJ
E/KxzmD90Ub/Uw/vjH7QVCtXsbRll/qeyN6UKvPXb6Xt8P20Ls2Q6jCWLKDGeCPl
7/dFRKLdn+c6ExeJ7N6oedMJEF6bgwCGIXlXH9buk2sHxH21iXHss1EqRg25Ly8l
YYNMUSgk0q/UQITtfeNUgvPacY/9tjGEODx9X09RavU6wQ3cZKpWzgtYLvuYaD7i
XukyXyZF8lLP4BDsr4mrrToKIyfER5qu+C6y33i1L4ZiqoekhaxvIiVuh8wWgXB8
UhkFfmJhqEQKPPaQ34EfcwWPb6h66KYd6tScJoCuHnPnTP2NpYnhd4Y/bY5taZEb
JCXM/CoMcn9dvWArNUiOGUELSQcian3f8sNb9mbU2maw/pWRmFClv25rX2lWpkrv
/7HgJgQdXxHhw4HSXK42qtRWakLAoaEbITC1EJiZOnOHtbikxKrpVyhFTA+HAGqe
U4Dt3C0dUoVxP/5kcvfeVa1qUW2JoyMHNr/+TtH1aXF98o9QRAErZRIKnKlII3j3
zkxHklbvy9Yd5saQ5glaL36h9bCtTobB5LBW5HKrDWApVknux4Wfx2fJjvP69VH4
B2u+61hofQuPTLxsRbmm6E4jMxauMeo6chqOysUEEsbjdTEc4DojcWyssOPY8vkp
2UHzOwETLw8vkmeuHwC1CXoYZD42SRhXYcVpX05j9ZPKa2NwYIJULAjY7F7maE90
2Ezqgyc1FY1aohAlK+97bfZIDeq1C9L/3xaSwj/0UlKlEx8gcm54C9mXAhmYdo8J
BuMhKMmD+l6VyGlHxm3s+s/PKX/tUqbZOqFE7lvcnFC/iei6rBXYr9PRZmPk0BaT
uNBfh0RJ5WCaNzacHVJfQglIF9kZua0h/D4drmOY9FJkF4p9FC957PWuA9X/+lUh
GfHKTJSsGN5wtg7W0SQbLG6hQhfWevItmhUCH+UM3GEtQR0ZU+ZTWd3TDjN+HVuw
fl2QibXZlWF/BEmCexRg5ddFVF8cnXrbDMp3NPe556tKgfdtm7N0XcrQYx1wXbmz
NBNiitf6GNIqyopzCVDNw1k6MkCHMz783hNnFv2xq+8D1zQob1/UmR/bmxJf1dAB
PrLRkHJZQY+3cQ73Lv/Y9ZsJ8ew9OAn6hO7hU1Hf0q4xJE+2Eq1ol720Lwy/OBkd
g47K1GkDJbjutkllob4w9jfrzR9xRfMHTs0ZkdOI2MqNQc3SDPA3plpff/qptmAV
eWbnGpZFB9Yo88s2+cPnHjR+JXfk2hCJWf2Q5kL5DM8htwdm8Jf+9GcGRLPjmwvu
FjZEdihY3RhrTImZ5s/X3WObtzA5Q/o29wrv7mdIfAd8rytyVfRS4yLPJBWzURQW
mT3EH4fTen0pX9xk/TBizEAB4dzt3116s5d+DFYzzgvTk1ocelZLCj7a4NtAAk+D
TzGG/6sI+tKcOu29lleHtTixDAyL4Rkag3hDQjsPia0vfTmaHla4CfK9LnHxpwmC
oIYFM1Qkqz3pRD7JQUQHZH5S8TvgYiO8ND7uF9IZBNRz57oIsD0TwEouyob0AFYf
VojOMsPjtcp2OdfAJ+mEGzcU81ceAVZ1XVBOdVeECK9X4skDvR8hzOCWx4KDOokA
g4pCmvI4JiA+rTFQQ7wdqjniFgdgW1w/tN36skjWcyWK8uhXu5r+qI5/TSVKIKJZ
KJ/PuJBRVRV2DIo8/e5ZmBotOoZ8O7i/gEvEfZksgesQ++YgocB+/GCPOquDgyRP
0CK2ywfa1pSeujY6tIPtcUKQOxjH28wCDn23u7IWLKwy6hViCGEEMshUDtn3RjbI
+8gSCUcbfdfjQtVr6oGqOqHgFL8IcDJrYhcU3BQ1NBw7TLOovXIxaVJLEHfOrm2e
2/XXh3otlocmEmvMI+BDZ+fcETYQgvY2L8dAKEyk+oaEDlefhAkAGC7DLNLfOt1b
6+rkNzFlpEBKj88ehIWp0xyyFhn9JRyMNiFqBOAsWwR1Bpjkz/z++Mx7eXJaC5qo
EEUmgwgvO+Gpc7gRU/AMqfIXI2+fXXbFP891IyaK+MvylKR9Qp149M36QGfGiTy2
jn5aK0JtOpfOkbA0RZ7D5QV97k9APJ6yVfuj9ALwr1RoHW3YsYYsOw5B0KipjB4e
1Ky1Wfl1kP8a5wAHP+7VxVMcy3WzRLbPZ0oL0O/Fcmf+y0vRlR7onBqsRxbdvkie
2tLYo3tusDSgybcZNg7ybHbvGVOPRl+xBUBz+0JbhT1OzJBIK/IHsfURCtrNegQD
bxGounwZXUXlxVFdsgq7pNDPneMxopg+Wrssrv1GpQiP8ifKzc+SuPzIFJyeXqeE
+MorbypdnAdRgzoexVR7l6dnxPKP/j12IF2hZdmgmkebO2I/AQdyAD4npHhP8L2d
0RiitVefYXthqzvtA7DyZJVbO1e1oCf+Rqy9k/zh8+Oy3yNfb5BenNkTAQkW2FYx
CDecJM2E94+10elMkOVixD3x9OLC8PRE5mI/B+R4WI9rr7nqxduijC3P2Kvtx8tX
A8QPxLXx9EV0lvuSO+LeiFAVNK1pLYJWuTqhnxoPfVOZResxIwnYoZ4rt4kfvDMa
7mATNraGPDmJ5Bc202HSaRZZuapYefJeN9FVc/i5JlhCX7VvDOjAfYyZqVnqfKr7
A4J86LmZSnDBeWhF1gwDK2ACyYQ9ACtVUtQAaSYF02u2LQsm+DahWM7/z9F8lEDQ
wM7esHgUqlcdgw4wJU30zvcHWXdoMr5FJEwrRr1WegJlGM/SCDVobjxpmOq6SAV4
2TxcWPXnaC4LBU2j0IYjKBn0IjChLbQOgI8NFH6O/wIHl4sk/AF86ll2LBzW02DO
e0tiJue/nPgqXVMrCR9P5cYt6572Y+x8yMr4gz6u8zZ9s80l16x53zvDtIBs776v
AOu858lrkA8061uDFRlcBZnKCjP3uRKeLpMq48GrohZwgwtj4C8U5V6MMADLTGtT
yjXu2Et/l1Cgp1EpbOdf/Gf042JJ/HSbLtT3J0zuAGz0MEx2yzu3Yi1yMjvHdivF
jwBwcA9WM5eH/UnBNYiDV+8Z2sdI/8X32TyGk+LdXHkN7s0Fk/nBqwJ+vRNIPTYf
5qeArph0EZatQPZUG6hnEqUH9l0uXPYGDuSTwoT7MCgquLDcsfBEaIc78xa598HE
KJgG1FjFi7y+JV06QCSV32a4eHucHcnHV/nNRq5vYGoXrmLKOEzCkd4nhvLiDMCI
skaHFswcqLdte87sTtucjpxwYgTUaB4NjMGhlLsSa/periBEX+mvnVRjhS15CI6i
GH31ohduQCaMxkr2W21oMt35mvevCH3Ufr5J2o6WmPIQ9MT1KTl3nDqGhoyU3EpW
LnuBHJfztnKpUAtPGZj0HJPh/mNgUeKqIwbx9sr9RMCmcuIP7sosl9JvqrKDZ7M0
fHJVrdT3ridU/B6LjYczIWSK0sbAcX3e1Isht49ozcVaBQPZ27mrq6XTU3J2Sk+e
PEOEwTXdfv1zS7q6+phX6zbaexh0pZAb9FnPdMFM/mPD/kK6B0bdaRgehpgOmMH0
j5vNMizOOPftZsqy6S/Df6AlsV/AHTlCdNcsdAfz1prd2V+ZL2U6B5Cxcxzt3Ki1
LL/ktAI/9YTo8hItjszuSPosqZnQPMAIPParPD3Dmpr054HHLZvoCO4F3UMrMby7
m58z29IyYtnM34el44LegafwFtjbmeMxKrsmHgjDse5HmeyCbhA6+sBlbo4v+2b/
b60PFNFRjhe3ENfTo4438vM9qsdtldeiNHYXmjahCh422tICCCd+HPuGmUTHDiPE
PgUUre9toczpJNVtRra29IbKFBMQdYoh6sTAhoFnG9m+0RFO2yS2AZWvkkJ8+yBS
TYXEHCU5nfGzukhL/jGrh7a9abbsJWRrpIHjAOVZnoHq5Hkwm/JHNJpk87Mb+Vsn
leX3wJH9GkhnDKC0qmI5u+z6Jojp4wccY+tet7+g4iZzb3DnNflORF7m722/rVxL
ZoyHNjnzvHKuey0EHcbIuMl+qVr38rZE2MKGB/eCRTBJZSsa2wEePj8StGl8ItY2
x955bcH56BOdesQq9/DMQOlSR+5YlItmTfhmn3tJjSOOGX6627hdAbZJ34VZMUcs
bF6BF2i+HKr9bJn/KFSl7QWzwz8nLrzMZSBHfuZwwz2MmsrAG2Io9ViBeMqbf8V7
U3XnX1zA7b0Yh7OZFVQg2NfHLXIoDkf4SwBOFY0Fh9d1aTWHIQ9pGlyXI1JKaEqE
jzRSztKmzHQP9iwONEwfydTPLOTxo636L+kJuGr3SKXxURazMPC75nJKNeQStWHl
oLiTwEoKfpr4tznhpt5zNBW9IgTG41nprF3IyK3ALfqbd5Clo2lnpT06ABSWo2n1
B8MbbVeikl4QNkP86V4oeXlRQGXrD2YtzAOyC6svWz0YK7PpfOmSLabsf6n/5juh
9Mo8NDOvjG0jUz0JrWLLCOfuzoALZm3vlBXuYu0cYjswvNgrvYNHXlSiZMl6QWc2
r5JkosDertZV0nK/vIOaIoQoFX9L0p/3gBDDzk2cbkc5heHkq0lptpYBQdsB08iN
l4P/wESDnycXVg7rUNqQrnzoA99sVJkAuIwiYaiHz4LjjLiwySczh9IOeTujROkb
6HH/Im4fCL5BCT/P+febAirEqM8NGoWCMPAMoJqljIz195pyIOGCyqAalZYnKNn5
6UYtBV/5lPxNYMBLVtuRfSPVwH+CGTaytkCBqfm1LlfK01Ri0ejHSIXLg2dcB/pU
LcAfJnL3MlBn4kG9oGHYniyU1nmwRC0Nubl/JtMMG62JQ+qWTIgiDVX83TaBdkNg
FRLDUUf5gmTXrIkL0QIu7XFJFEVezzFAP2TC8JXf19q112jut9/opVed5kvtiwvC
oyGdhi0CzHQJHGJdqfK739bJfLzKEU5NIjtDr1per3PsC9HZGzvDjKbTrUDMYYGM
siidmXIeSEH/PvRFTJG7U2yTsniXmpP+VT6Z3A907+kJmp9Wn5joWA4mGPtp150s
1mj+gGwyR/H9y6UqqHYqIQ+iAV5D1UbC3I3+o3WgcXlN0e0lMkAPJmumRih/gbKq
s1toACNCNxj73MgMmRtRpi++QaXyYfenPZmLmt67vXlCUidsvFZVm+1u1RVChzhL
v+Cz4bhear9hUUBIPyhDw8bSw0PkDzIu0loxdqfrYARuOw3r7M5HjH+0thpHymfM
1lu6n/Y6r1KZ78RFgz9fUj5H/ArfsVj06LI5N0+/hVVTmGfIhwp55v02h5mTPn69
n3/LT8Z1XHIIrrS5NFPRCscKelp68Wx7Fx77f3N0qMa8EnFAs7vM6P5Ed2HzZx56
RN4cKnTw/+YUilNE/2AdfyUmzedHdbXil/7GiGIsyEeskET44NzvxwBOrvYByCfG
xiCk8s/ho14J50mWXTNHZ/KIYzi5aj5uRkOG2W2k4z7/KFi06VFn5UihYFpOTW6x
PAMcR94jpHfHL+AfMND5AFWdkLxwXlYA9qScZ9hMSpG2UPNllzhPKzblabIqQx+/
XEwBM8oySUyo3vxnfaspmvUfNJlNKvpb4aCzkzGK5FnrQMLi3Ay7asrL3Vd1J90k
Z73u8T1G0opyM1wZT44Sb+6u4l6XdHOOiPtov8qvYQS/7oHcMU++nkyNFiXzSCWa
2V8UH6TDJ9Bbd2Pope6iLcMzBw0thl5sDt/KFdii/vPnVViNFVKwha1ZkpRpVcR7
w0MHW+TncO8nZc1/Yo//9ciGly/ZCoZQZE8ofl1XNs5hOIEBkJca2u8DQg/RFvPX
xjBuhuzkr1m5TSMPPgsGK6qYilW71X26lgKwzz+CxFQE5HvW6iqKUpMXZrxg64Q/
TYuA7J9jmrP2pWoLwiKY8FhWrG2P/4AQNIcJShz5dJ2YzPfPnIUk9mVMrGAMxKP/
v2AxrIAmF9Daa7N8CXFSO6zBGMCxCUVVYUa+t78vaq2peghAB8fCHv6esn7L8Jer
4uDY6+fygWjPQ3P7KyM0ThNbhzBoJ4mjHhy85sWHTfCijHXSVHsoRH5fldZZ2HXx
ix7wkR7Y4MYGbxBCjREX2eNaE7Ny8HKfRHiQT+BbW3nWoCCpuzZ7zz+hZu8j/KAg
zmyXzTQDc9SFsyHs9F7MnnF7G7ibs7VvL6Jr5h8Xm0Fj9PI8ljP9pQ2Hzm0pnjrW
quAMPqtgmfh6Z8ZhTnYKIrDhcw81PYap897I98jvTxt58udCxf2Cg+Hnsv2WcHhi
OBgbC37n0KHAWLg0M9aJPifK6ulxjh2g+hkCQGLdQR27WDZnWo94zzMwLy9986NN
oaJ0yI+XAdAvkIo5WKN6OcTgH4N7K1yb+LpIDrpIq39yjAy4s00WAgn99KbAcPDD
Uw1oc0cp5SGcwEi8+Wh1FuT45QutN2BrnLKwUFKhtEteGxGLfcc2xGi7vK97K4bw
FiDYsfF/PfTlO6sTBTQDuhznoPZqceJCtNJ/mboWUIFckb84tMxIWnihCSsRwtkY
CI9t+7MvsSjjPPp8Lsw2l0EkVSiwp39liEVOPEuRp7aC7Tj/6/WIoRtpBmBdkLfp
WRQUvcPy4ALqDuzGWQOdf1Ki7pM8Sgrixw1b21SP6WVw9qdflC5/M56qXuAOXt8f
xxSjKq+2L2BCLfcNHYT+RSL3UHUkVN9rReGcd2JBXMINnZF1h7zTB5li51oLEmit
zKrdCJG89VLs4mVXmH+HpThP6SiqMrrlpwJ5e21wcwldrnnaLFOnUhxkk0LAwCHc
LPYAoYAbW1YhHOR8PZMaJk3rClJY+5NCgG2wselUw1DLgMT9rafjKAqnKLLlq9AH
cG1uSygQ8IcHN8eSwD0UN7srGyVP8Z9OsWCko1YlD2cEN/+5N98M2JYsWZhCnTBE
4vuB4m37fP50yIJ1+ZEEl3QfrSBLWTFHfNAEGqRbfSJ7HspAY1HaN//57ULxiNFl
CHvU0YhbJrBOyktCbp3J2qEczKJEXXkbawJZIpgWNZHWgeRpoQCYa4h0EJa4lkfv
+lNEa2a7d7IcrfkqNiEHg3iZsEWpmMNel180XfLNhXj9rvQK/yUlLgz09Rk4vqZ6
HgbZHTvRHMGmSHm4+xcUqNxDA+PAGecaPZjoEiZUcIRlFA7hH4EZQ7Tp05RE0kKV
t3Fgd6oJ8V7UBT1o73Jd/4PyF4u62qheW7kxrd71vsTXteJDlQG7lJDF7HTE8mdz
nutcl02Lj09mVa74iGsMAcIPioRc2of2LCcbdW0UxCW7HOk6eHlT+3fQNBMIOZ2O
iPDrxrz6/wl8yFuZDPfWIAAyxm5wEnKOuYPfbSIKSNWw6hWiJwAmO4HZaVSPHm+l
FO+0ihHsAOXNxvhSnddQsElhUCAsQP6DF8Qb8ShzokAGN0oa5VauyBIFT5GnqMo4
+4n1YMJ7FulWMwJb3WYBbS3ApQtCqTg31rQPwUO6Q4lBGdWln+KSlKRqsjaLoUag
q51IxsE4hVuhPxSt0yu9zEL7FkC5svI9EE83gWS8iVBFE39QQrws2hqqHZQ74/2K
bI3zF2S13KTwd/ZCz4ttPQ0JU/IC6QbM9j05ciL/U3M7QBagnlRNZ/9NIuhECmwk
8n6M0YQcIwmfHdQWlrbJb1aUkgaWgC79BskrD44wXqOk0Z6rg0kL2qOo6ZUpH+jk
J5GRh0Lab6o8N+RxigMfk6Z+udE19PQaYR+LkURArrXazEvrD7WEmkv9aRaK/LOd
VdepwgidR9U7s1QgIVLQQPygokpyvyWZ2Nt1jipT6kasbhj4sB068cmEKqYjquRW
HhyK/TfrkgF0S9iiIT3KS8hXC3zCEey+9lATg9E0s9hyGbnWccYsSSvaLACY/PqU
FpWsLcyNZdTiyfGBzUBw5BAS1mtqOX+LDoi6JcYbAURb8KsAa/YudGlubHp1p10S
6XJ/hbTbYk5uU5tiB9lkXn6n1HUU1x8bl/7eiKF9eV5jPc7HY6HJYoLH305kZEst
b80HWOQpMSApb+Mi1WGpSccE5LLK/qKUEJI3mIuj3ozNQ5IrCakuyemoXFhonxiG
Po3cZ40IDxb9UcVyaQB9/JYGtOBmpGmPFQgQinL5IBTDs3g+AhRFYQLodsiMsDUO
iy8hQquuwXT1F6azQqJbWrLPpuk17w4pkQfZVflq6oPzwFsAN8r3c4FD6GHcS5QV
l/klbrHvJ8MGBu7N/edu4nHyJiwwB/Zc0gj431LLHys3ncVIembNvmW2MEQ534P5
jqrEwS/raNWjAfVhk/Ks3w27Rbno9zHmJxqeonzJNq9O+D/r/cPuMjKxfblM1rEt
8G1p3id/8o+A2TcTW10UhB8m7HBqsId/VSQR/KfOTAd+oT58V75RpUatVMb5vf/N
E6iRWzomTPn/KZnIhvDT+69bTOKLtZ31d1M8w1dUygX4W4kz2iuNkK0P42XCFVe/
1LCY+7PUw7MAdHOAZlmwevAHlPsxyQL2kTZv+vlxVYXHzdkraEVrVuhJY84gxSHf
20PWi06vQB6XapyL7rvxYci2cQvQjeTxad7tZyMabXj/06XdWXKuU0uExrqgwPHs
Jx3D5/z0gjWRdUPgYe2JxUDfJo9Ex6ThzBCopZMt6p6k4vsFFwlWCd9Vmin5ba1W
1fgmbHZQBQq6Dwikh/moWWMexYbf3pLe5v/YqfouAZm8BNkDGOJ8cJJ+0sER8Z4Z
ijdF+z6m/0capuaoZ3HLKX4tLQ1Zvu3y7fl6U0PBlZghwKj2ToZoKxJARhunHa1m
p1vAr6zozeNVQToIg/VVytwOFe4abM237SWq9TAg+RHn28QEdXGp/H5n3u+sAGwp
Y3sKHDzVLhdWTOuB3b069XDHwjMw5qfJYuz0USfV3z0HR5d9MwDUo1tAYoTp7/Ys
qLq0MrJzeTf2LyY9nw+5wBQ0t8ZDnVtw8jGS+j9RPWWCwL0FFXK48SQCNc9qNnHJ
KX27/sQAih5IAbaL9QKry9BGgHnKZ14xzsJ60jHkAarQUU1Sn0muXZ66rOJPKYij
ExGsvO7f/WXEIvvQsqgZSMF+Bm9kM3bOxKcPfVEGEAJFWXjFFkfLSh0qg1rFlUXP
2oUqXqWRLTXpCnK0zWfhEtojgE2NUUPO0oikd0tQqtcq9oviaADVWKtH6bK8+9us
PRqPWGg6iAMxfez0YujtgpiTIhC7FtWWPsQ1jrRBXn5jE7tTTqZRtF+giNLl46rq
/y0WzIPzoMifhXuLC5p7xu369aQqGq/w0cd+4VhlLtkoxVUzZOfmAMJ54NtVzE+L
hQSMcsb7NDEBRJJDaMLbEbzFEeMdhAVQqwHZTPQt5PryBzIgNSTp3ui6t1Uwy19U
Kbsn9GbzBQGQi9Kc/VFLhs6NaRL+csGOZ/Q5M737nF52z5SUlXprQaPE3dSZQIxn
vwa91lodwqNLcRx9f2sfNws7uzkoQFpeR0j0PKv5MCEqEHtzAUcAgpTAOk6EjPrC
scK8B7O9dhC/N3HX/TPqQ7ixy/UvN9PHhB/fB1SUJ3RBqRFErpVUBxVQGAes11az
3qsWftX51pV78NBxXYtDB53vLFcMGgHHKd/gxHpU8KMtVimc6AY+zQV+ZmRrZP5j
xs9R16sSgv7QWvD9lq/GH0XEoshwZkCRXPK2jS5Fw3Jwq1VXxKSBJprvmO8CQILI
OefOt0EfVcBop/F6IEusbkco0k6DMyOjVt3Dj0OB9W8F9pxzqXWiqf676/FcOKkU
gOcTDgKk/bEol2GDcLSYj6Xc919T6VnTwO+WPoYILgnwy7xKyMW1AhIGCcIekliO
WBtK+ChITm71iVjVXyXrkskUuHTCeEBVafI36O21pnP7r0u4QjLPErKUa5S3CwlL
1pWAMXtohKYGvVb2OAKSRDlnQlvPo1WCfgTNmzP8Tu7iMkttnw8Q23Gfs6CMUjgx
b/GURpuzwK5HS1iqhA6RKtKa7d9u7sCrtyidltRK0ArwDrSGGvyJZz0JQRiVA5vV
0X563PVuU/HDy95fKu8WVaG+/ZZ5vTLSHBHRsrkQhGkjZNvCgR9VuExgG3Q6nQD7
4W3AxMCkT5fp5uFQzmuIArukLtm93SvKCWWzQb6y82bH/U1xVCp30DdjpbDQaNFG
mhDjp4b2L7bii4J2ctjC0TZIMYzYLANij0fRxxXDrcGZCF0AXShr9mKF0Au0bKMd
wx1T6S1Vko2otREoh1EmAqDiq8jej5EZ9NXEgoAMjssQ1N9292Jk4QH1ejmTJXqk
UQAg0JYi2FuR9+xPfdui6U3qhboAG8N8D+KbL27uzb+maqIpoTrK9vOk+ryM48Hv
+Oy/xZ/mzfs9XjChAz61PiOQ9CF1EH5AE55uuVCFHqX55YJZ2mxg7+6X7jmjaGIk
xUAj2HiSeXSGbGz22+mbAYPie3bL4fFMkzDaDKxBWRZDcDETonyqqsuafzb78dwI
bk6t7PUU3xRG01SoClpn9kMCXaorJwEXsyd6pmp35NyL957v+g5EojnIsljKUoUQ
uMvbej21W3q8dKiRWffIIrmfdocHf/D6TrKQPdYRphscOwX5vI9IX25x3QcuL1Ih
MsQSs49DbIxZqLqotmNHJnfRET/6Suq9D8IYotwzAo0IB15xZNXjhd/hwtLgMIqb
BdiHo9qml5yysg/gXBW1PNSYbpKPFweDwnaaGCO6MvWvcJTud5VEARdo8yfgb+I5
lh/ko+Ajn0SMenWVMUNcX+nRXJLxo8hW+zxBp2OfFdZH+E77vXzoy5fsgyfte8n9
hxgUwWSIOI3Q6NiRdG+mXDsjpdCD362PDI4c2c37HLcRGTzCh9/Pj4ence6CglmD
lptm94BEDEQJ4aGQJI+x1F+F3fcxdyu4ZkWFRvOend0I7mSRFGJSKd0JyPx/YE/B
cZeKOemvB7MoQc9sGKLVwI1Df+BuGJmaO2VK7aLPmHVOj1mx9HC6uQ8k5OE/D1bU
tZhWfVxIwEEAbwIQEbuL2jdPAxkPac4k3S+suLMAelCn4hNTPSBmG6EDkCI1MGBr
5ll//yU0Q447l2+tN5FWkT9Jr7U/YbYKAHaBNIhtFTNmB+bI4JpElWoTzyeNX/Ls
G04wA3S4e8sRnMtADnG1FGekWOBLjH0XcoDHoAOLD1jv3eH3XuRvMHWTdMtBZhg2
14NXYzlLDF9dT2o9QwRjYlBRSFPdeJDnwV6zEFDJyIbJs/Cakh/n3RJ33nYksiln
qpxavqKsLGpGMbmeMLPi215UpAyvK53ArdeJnAohvcLRYVLEos3J8wdXRpesFny9
i/k81q8RdGpMn80xarkWiDoIU/8FWiwedSr4TXzK5PJDv0KQ+ncgexUis1kuAMkv
GdS4OY+nNJRDR40lBMa8iKvWexTnfz4FDT17YZqsv+F/Pp6KEgRSLooF/IsTfm8w
Yo6kSPIIOugb2zWLrXDYH2/x1z0yXD4yDawOsMV4lhzJ5pgo9Mkp8bl7iE+68nwB
Jds4I5TrFNaIwu+4WmOosQjQBNH5IxJQFTeIR9GTv57pyXu8butC8pk5VGXYIs4A
w53HugqqRvGfjVtlA2dRgXFwR8LYDXyrHrrOJDil4tJGJYujpl/ZYaU1o95sEAIU
8OstBe/6thHrTmNno2dnpf2Oy6xqdHfxF+4Zp6anSa+OhmTs+VA8YhPtPqvDBYn5
p109Ih3l7yu+mcPlLHtr3wQ7o5dEHwzgRoLg5/6/Lq6R8YBotVYZoMBWKPxza+/i
1Vn4aZ9E0TLDC24/LESCnun+G0SCcK8Y4isl3jevjTi7tajyaSnf/DEQtH3QcSMI
A4X0b7sh35xTadTafoSnC9eGITRoNDnK8Py7Os5WnqJE4yfFG7N14qDwKDKHxMPv
OyIS1dZdCZaQksWqWL62HrslU0V86r+mW6ooMlJVf8mgyrmC7yiHJrQOkX5Z0ydM
rHqye7YqDDo61DYiqn3C1XkubMRtm91USig7KP1PKECktgOvvIsjJMM7yVs/1Z1r
RuVHSaHzF65YlkJTTLAlD+2vTakuSzEuU0kOZtB48YCDfDyEi4JVj8UFKxSGZTJj
X1lVkAb/3c+XWTYRnd+hSBNy/8dwZc9Wv0CcMml+iedM6hjmsL3Frnu3POpcZHzU
1HAym/bCKBDl19w1lV+n8OLz43NHcJ+IUx8y7jwaY3mLPpKmsuiaPfyMQUzOlMpc
a/m1dS8m3T1sKjZHD4n+tIKk4RVjxtY3nP529pzQpPgiEOOGIxGu667WLAze8x2Q
bLhrPcUkpWo4wC5vS9ItYHWbgki6Tl42HlU/9HMk/km2DXgC3aEDUDODejPL6iYK
/Tpi7gsWsuQEaODNB5mWQxGQoyGetgvGplBoK4BtZv3WXdpe3Doq0l5fOCjnCpoy
pkqzr3XjFe3g+WMTLNaGrFhYQi/tqWfIDcPgxo44hYcqj70WDlGecBzCYjCEaUl8
LCVpjyWNY3PXwk2ngbF537pPtxItnS8OsXBKZv0QgdWDk4qvyEtfs59jf+7ASCgL
pQLKqaMYXIxMDFV1El0OEFJ2HnSg84Vcvaq+8utJnkuO2VMkZlQv2ETe7TzNfmsR
naw2woXdP5LyCsGBY0YXN82w8MLX/aK28x5EHRWnqoRQxIy91cZt1kLVqK2xQGsb
lhzhE+bC0eBREjw3mwEwqPqsBBSh4KPc6hiqv0wETujNJPI8Dm8omrsHGEMRUs1C
2WCeDvROrWt5ICg4RKieazekGHC8kyk4e7Ju9AfynsTVCFZ9SVAqVmSx4pytHrBB
QMfEyqPc0RZcUbn9Qpt2SglZjA+mudJCzpw2p3ybFXUWhC24WETMK/AiVW/CYCv8
nXgIMPk/fnGRDPDShQEBq3+KjkQbuPmTzDgFUeb6ITCflCYXoOlRsVd5h0KVUjnK
hbRERP+SVZ7V8layZMAGph7wbRBy+YsZPLYzVQBeKW5i80NWyYLu++I96yO/+SIn
qnApqDQVyIg5GMvTD6e9jZjIzVeza3Pv/srfPnb0xsraq9KHRiPxZbyQg6pyccjL
EbI1Rs3zw7xDF9D6afywF4swhS7ZoEOMxc9YwpPCBbWjvB1heHCxZPlH3L8SuZiL
NfvmHHc66sf9t/TxeQfC6+ZKGUAYQH4CLYXsRgkDk7U4Co+6mYHv7RXDjmQBBr0a
rBKRDH/RPMIHWDqlt2HQQyW5Ywf7xT/JLYuHZlnzRuLMOnfB/6k3mrnYFxToIcFa
F7Wajfj4qh1eIY4CiqEXFaGm2GiS2btUg1yc4X6Db2coqU8bnda6IVMhXQ/seg61
AxXlfEDgCwdGyRmvGYkoVUZSjV3udZIWzJjJYGhwfCULVViHg6U0XSCde7DGWSU/
sh7xfqa4zAuP+az50VKLI4jTD1ZJgWHzpoukSblObQkUZF0vDPwBzeC3UwPli3JC
VO3C6s0QLFsHKqL8PL3aqglim+2vfkRQNvNR0FDLKKAUM1kFBAcOBjBbTjxK/WsT
rX2b9FSNIH/hTNeV3maN51gHDu3z8Y3i8K3K1vmJWBv8UKgxYZj9wNCJ+bzd0VIo
UmnmImwqSzzRm0ChABcREJDeVNgspRWiAQHZvDWbSHs827Pts/t3thYk2PSGqCoc
V5JjdqDavSrzjcVV0Hlf8gd80dJ00qcDFfMVuOdXC3nird9euTM3jx8eIcE+7v4T
UHLOY6oC0XcwT6rlNmwXMJ2dTdSYJLQvXldbk+6+bA8AUiowgntFZurNKa/bjjUF
JmJ8r3lYx37iYByes37M2Yb31j6kg012t/Ez3e/S9XJNrSO8idCihBNqQnGkfGnc
nuxUVdYMl4I75UKUuP9BKRbOwBZ25NI9a1mltupQtw03epBzhDRLGwUTgTMLqMbE
sxVWt9YuVpQj/QpD/8DKEADuBkd64/xUf5hgNikqH12L+e8yz8HcbrX/Z5Q2c3Z0
T8nvOwYCQVSDcXy0Z8jYTcDV1Zh8dvX2weHdw5awOFpYCoxneWR/VN2GxlwzhwQC
KIDOOK0rR7QSms3a84ppQ9Xh0cFdlE7hxiTYbse463p/EMd20ntSaRvCrLG8Y5M/
3UHeT/qC5jxL5ew7fDkURYpD3nJVDrzGz+vJS5AKb04XNwFZ0dmFTPbNvwjmYo73
EoDVBmYDirXMHg4a5Q7RW752rG6nyzbGrVD4AKFZKJEq5DcSn9qdetqr2aW/0J17
0/vjP3lVX3F1xgWqGkFqwZk1NsIRjwHvz7QtJwOsC6V/bb8t1hOnJLnTqe6EgCSs
IwDCvu/bfwiJKHH6wzLoWov7O/ERnZXHy+gjjF4EtevfcqicTBmIu1ZDzQdT4sBv
Kn5+vOAXKjfqCHulWv0iNN3OBMwA1Mb+9tnS1UZUzMIJu+kE2hXOpmt1qhbzevss
nBZUnaSwAbHX+sMZYDr1Gzuk6Y6MxrhjdeSYNnEsSjGdD4zDM+5QJSe2L1nT4dL4
b66HDPCA7wN1bdE9rYav1zSRRM6giTkEhhLouIJYb1m0xjBtbpscIr32ynYKyMeg
GWmPy+MSz8m+kY3lltH1yFtUXrdOHgS55XgxZ/a8/ogfYuoCFTF+PeHS4J76F22R
89TK15clgUZ7zVvEXY5weJTbm6bv02ih9NqyVALHQUrayThOo2xPQ7RAL8UK2vtu
KZ8TDKsyE2xEaiOo2fG0nhCQ5b1+QlK/KzUKo2zWmFQ+GlFWviFEd4VY2Ggahrj4
WlxMCFfYYCUauVBlp5nJuB/dCGQIEdaNtNr/bShzg5tUUDMMhrJW9KTRx52JY+WF
R93bZiBA/nclA5qmrKPR4vHOgpR1ra0Ya0DjyO3/MHWO3mIODMIdF75mPdBr1GYY
PbjT8OwKF1MAG7nx9h6dDvkSn51eFxPBfQ9dHR+QW3aTUcsfXqliRiQhDENOZSaD
kQZQH/9tmWE/dKlQYZGs3Pc8WgUY1jR1ukV7kOPZHrRTGWKp9NqNxKJdMUHcuk5K
f2xLybONOfETOJldoDd4CfmvVoxY3DWyF3WIpT/j6KLmygIdqc6LZ6M9n6W/Fl2e
H0Osi2X/h0m2rIXsBIpTYrHMNHmjx2HTgJK5//zY7l7jM1ygn3Qb45J+wAQkC/bD
1ww5BBZGppuihStFWeuPT77VCYezwaiQYthV4eU3Y/x1a4aU2VL9FtCmOuaPT48h
y2TPpBIF4NZE9LNqnmIYIx3bCe78avhUEHET8F72du1laFcERjybWWnVs5lOHmzY
EFTRWar5fj7Ze9Mg2m+TJTZD58diUorO1HeiF/ZZyypVD9cZipIUu5GsCL2jSpt0
a7FelwlMdRrgm19sI6aM3QXXRQLSk+QT+BToYj/Qs2xZXkua10RPC57whEBQPlOe
TwNRxovxRM9pOjMY4+HNsYDntPHyxh/mX4H+01dIXmIHCI8hheBXbomtH9hAeTAN
QqlZMbV9bkRJAKpk+vU7ZElnZLQ76Hbh6HnzewGpQXpd7F3taG2fv32xj+zZjhC9
/xZPKLSx0dDd3s2wuz2p7vUdp1sKTXLoEvbwVne6cHWo5Obr6mGYEXpGYhrLL16e
nz9Gzi1aZCUKam9MwU26Ftx8kjUMM8wgg/qwP1V7ba0s8zG3yJFa2UqY+kNvH//s
4ZZwfAgRpGO3y8oX94/IHuID0EA+ZhKRAdoP04BVOvN0uz+r8ReI9qdGZh33pWLw
I3fiu73AOjzHd3w+LFiEusSvJZez9F8usxnUKz6ZE135TzX8z3KQHb3mAYlkf5ql
NB2heG1h5QibZ6d4XI30QcUtlyl9aXAMqN8J6JdH+ZOHj8oqql3w+sSOc0xOlhg3
XLPckCrqBhDXTTAGFtAMQbdPjlQs7dAzv7kovWxkaAfYnYk185G2fWvOa6vv3Bfx
buhm6xNLykXfN5ub9eStaODqHycprHdYl2NK9WoyH75+8Y1cTwnyQ1b7IjC3KCHN
cPIZekDvXc/N8lI2mzzIdpqS7SZ7pF2201tIfkR9b8jr3vycnRJxtfV7szOQNvyp
wAwrP1Yp8esQk40DGc9Y4mt9LiUGWkjeQ9So/poYKIKXdPKbLI4xRcRDK2Z9JJjF
0bMaExKsFm/PQCXlEufZgG4q5b8TPabu8eq1uHFHhtAIEE0ALO7uk3cx31sEkniJ
jaJf+E82H5lpjIB+j0vqEPdrDEzAlcFSmDlwA0LqDQR8kwIl8Auwar0GQEF7aFwC
N5AihAHnMrZnzc1HUR0aqLcdyiomDwNx6SAb6RWP3YKr8ixbfVwc20vIjRkA9Goj
YgxI60BWX4FVohW9V7ZNRDouOStjCmn+iQDDKJUXYO3GYiAvPIPpifirXtq0Sc5x
SyqOKCmHduNcecT2oRM/TLMFfBZ+JOOduID04YXW1/kas8rnJRddGmjkkp413pMf
ewklKFWZBnCZAGbQkZTAVSsmyuXuLyg4bZIyhaiISNxulEPd0AheBg/LAOYBS79t
f7GaHB0NIViyQhEs0uApQ41dwcXq3GtiqDfTMytStUMP0zlrsQFI8wb6M/N7TrQn
8pRNSk5AdT9p+IRciaky3oeZz6SYLUYOYB9ARIhGYg4dFKO346y0r03YUr8wnY2J
lMhNP88o/Si0FimySqasEfNhci0KXdKkOfRDUcg78lsIvv/LCtnD2huiqNkOCBBN
1JF1vMvoaOGHm1Yl9dkivOZneOXI8uJ+4LhuRwbe0VtNdziSDYTTtlsP5o5c6mB1
kY1u3Vc5w48hYCdz3Vb15YAYC/mPttiUkdRx6hBrq3eSTgbej6NZxHGPPgdwx1/Y
o3BXfecHsN/NRQRyoBr90zGrBpplmuawiVBz36xeT+qJmH80uJuzLoz7anyATVPK
iaW8URTPfwJz3Vu5yVxZSpibFQ6EMbBBH557KCJOu2lNcLO+sQFqCIQ3gCD8/PM9
1q17QG8+/O2wjMvg+IGE9YoCOYhoNAGr8Sg7TTyapCKtib4l5r7vW6F1ligyrJk3
njaxEIQeglw0vGqQ+Q+/lYUp1/n0ShB5EfXw40pauqDJMOYxcCow9bZq+cLMjSMQ
uaZdiNjLK9EPPZmXTmsN5lTSL3/5Th7Pf15SglMng2WeTj9V5uv8Pbk1WWIaDnAm
ZpKJ7Byyj+TrMGCcrDcsI6PZxCnD/8lW9UxFrH7if97QC/mjitJ+xZQcJ6D4bliz
lZO/nqL8DL2Ygrx5wqStaUU5iCocotXfdnrEOTe7a0OKXQGbqYNvC4eUQ6TfNEbq
GyDDO7MzGSJtvXUjzsAw7UMSNRSi0YwW+X4uiKgzbFDbN5ISLHW2ubjvds81L37r
zx0crYg4Q9iW3o8L92i6weipwVj2ulH9OzlKraC3GM09nVUdmdUkorxn2g+xNpSW
zRMyXxGz/l4y5ABDppkWbqsMDYVoZZoxDSpIYzfsalI5y6WsVM+auNit1bbhc52b
lynT7Bkh6RkEGiXaAwLEq5FcKdOyB6+3cjB3Qpkpps4YZmF/ZZmA/MQov5645AHj
S46NH0qxpIuZmn0jCd0bndHjE15v4mBg/163hrEZEkf7c/cKGEYilAF0z3iQwr+m
jwUk6AcF83BxELN+26ex+5CogyjlTHwl+uur8tbW7kg/T75WWPxkWJtjvFsWEKn0
wnat5JioXW64y2msmeMKRNYEl+4d3H0dbcXiqMlHw3LEcrmqWEU5tgunN45ICT0n
6ATnu+mdo6ji8g+z9KFEJuR7dTnke0oxMHv6qHoOjhDrrq46ezK3yjA1GhH3bk1D
k80WoZp8rkDa5V4+BXjb0FMuHoG/vL1HTFJFXrp3VFWSGFRl7Sftlr8VVlJFsIiv
Er8EDN4U1SuQDthBjpPPmsdGlP8z0F/RjwVdICTzRP0hnK2SCR1WoSmqaUYFoqFx
mP2GLK+KTcjLDwwIY9a9JPuhssV4IisM6n58Cp8RrxfKYoqNdtJuOemC/eY0PQxF
7yK4lA16B0+sgSezPkYLVG69K54IqFG6FNTXb8QfitVGVWV0GtDM5SWz9dRCSM9j
HPSORyMxENVfiK4twUZync3V2xvJRNWc1UrTE34Ouhw72KeiEwf67a2ro7z7NkGB
DINap8uuVVWaZxVVEnncT1B3nzZheS2JMSAXE9HpefHGIjbfJED3IeX3C9+wHFf3
S3SNGje9QMmb01fziO97DV5WdvmhZ3/EF2JXCWdkLXCi1IO8XC5cP2DX4KhIQM10
FF1+5enTKWxQNSDLzjR6Qm0TtVJbmr2xO0erFTb5yr0+8ivz5vKVYqlXv6EvwDFc
ChHIdGjerime9SQ18ghSto/tu3SoR5CkD88W2fXLbBqIiPidUrUEEVOYSy/v9sfC
mQF/1l2rEQOQLywRLbuY0CjJCRxA0dklIiOTXyvE8ARNb5jVeZLPIFgFYB9nzOSR
YaSFbe1Wj9CYmZhBONHEByvztfNaBbqUyTvG+gPlwUKdC94EvmnQH1urQbppBKxN
JOGFW/ZZup/Wt7TCCt6S3s4M9H7a46uCCad297tk80njU4Dm1ON58ce5bNTZYVuv
6vl8Cc+HekYJMoRX2Uq7dH4chN6GiWH69J6l5nSigTeR+YwY4GcE40WKToSJJLzW
M+HaigRyh+D2sYMOnYO7HYsQ1p0+tjrMxNWFZUtCI3iZ4TYkz5O4lPkuJ6yJpN+l
rfxt8QeJ20l2wqJYlz5r7c/jZs+IU4UHsjzE7cw0CNA2k4nPV6NkJzgqAX4IcO5n
eU6AkVz/oz5dl6Jmwi8fHwYeT1tIrnWjYbwFUOAivVcDLJqD1SZ73Ck5R9yeY6tz
SBQh7SLMVf1w5aLYY6kWbjK58ntonpAxRGioUkk5FDKmSXn0UzWJsFzPxUtPygAp
amSvJ5j5ko0A0PMzgsXkAJQReg+7cKIttBl2NBKgQRWviS4bqP3jdhiC5SPh/SDB
B406F23wbh6PjSYaimEFEoVrbKDgAmFAz0Ng5BQ5swtmjPYMLqP5CNEZJehyLXBf
vlDvfEvtL0tfeUag7OY3VcdGhvvt7hq2awUcojywtnPSmI7M0SojX7gnUrzvXsJ6
yRq1F8xEMfWXQTynhQ3jOkuN68JPB5FndtT3LRihvcvMY9xQcT+SjHBWTp8SaRXX
0rAczm7vWuSy/b4TGcK+51dwxU8z1DHK136hwcjJiAu9fVutLiUCkL0QN50cFNZv
J7kAcf8Ots+6mhvNczY4fbqZjN+KJjYeTfVHesy5ZEkGbPI3lBgwTeq4kNfumj9I
z0OYZ64z1RreH0rl9hDskHoP7OZQTPahQyt7Kk3piaAdjWhGC76sShN0m+WU3eRX
TJ2EwGGoBIDlQ1PzXg67+Sw9La6S9pEFbIn7nbpcgx3f+73u9G5dcggPfb9/1U9+
SOoPcr4ftnDHk1JdrQBpdiWrL8qPLt39BKKvc5iaWDpyniqRdH7eQ7W2vT/slHcB
2MRe2W3/BbgVw5HME2h39+cYdABUKhX3Y7PBdR/b9nwxp+HzkfBo2gGLK7Qec00Y
dY9pKEkTeKE2c91DpRnVaY13xoHZTOT/PFighApgwBmuJOn84TZXVId68pnIlYrW
jDQAwDPv6Aw/PJsrnVdpsRocC6OFsW/OTK+74AFV6TnJ0dPVPA25oaLspqXoL6Bp
w5cj1HSOPYxTf/16eZxmSz4Icv1GyiZ1cL5hU1zbeQ0kw7eN22t8nX74YkiZSthl
3sIVFYff7ynrlxeXvczz2NPxZ/bYe2rm3dQZcVWpseJAYXT4NFiiv1xLR3hKxwSy
CSOMNzAG6hgj3hkLLCFGYAUT5lieMVI5rrbhd8y0Qnr3ycWQjWIa8fdd9r5NFpMK
oOdsBa+IqqIeAooGgujN5O3AJB9oqEjTzi+Icqm3ukIyhmgqTRYsxAzmnIM9tznH
hQuJP0Rin19ZDHwEga/fKaKhjtQBKf/TUVbcypJTeI5kMJZGfEacc6nCAnzzrMIB
KOKgXebRFk5QS8Kqhg/YYDT9nQb8djXSTHbrMVB7Vnz6bpgSwvS0pgdek0IRe/3M
PyPow3gkVCxGjSYCa/kW1KMbWxFnGEiiEyR275ILzZ1gjac3aaKI3Q1kTV3n11JJ
6ABWGVgc0o+cIUyFxuhI2G9yEXYspR3E0cHow1dKLvLlSb4dptw5WUR9B2q2gIGY
fWatguMwsKH5waNYbh/1vEBmGYtRRn8HCqUUV/E2aXlR3lUg1ABaBFZFT6K0EOm5
xL+1AH2mjMm/+Qmwj1BqUpgbP49XXnAJ6xAbPO18ePIcwWjfTTYcEeBffdaFLR7N
D1uDQkcy5MKJ7g+NSdiEwaR8Mqkp2GDy4wHo5O1PnC8DBl8fIv5Rrb/WbIYW7dlz
vfP/TYKJJtYZTlgKt8ZFXov61X/rDLdVj24Re1/EJ8OKYRyeHGv7fHuWdDXqRfWw
fmGpUljQYf4h/ztrROEJZWXkHorpkJBDYJUmzJ6Nl5BpEnhEmB9KN565aq2b9qPP
aWkAbEYc6zw93/tsQkIf3SEaaUyzTLbGhiGKifg8FlYaHv9GNmYKLQrk81MRPGCC
7Mc0sSSCeom5w3fNk4Wv8CQKJDvPkiXJUBU+iujtcJiYpPmEFVEwrDTWlOWuLLWr
3EpFZ+N6La5Kcg38uaYgzHHHhVoQ8xZMdP+o4KAlR+MCTNFdY/xHi05XvSTuYuJk
quCBWzV7UqxyUJhBYTifOZ1XB95c4ut5CACUDcEvtWWzYrId1gZHZXVMgHdTXCFF
WPaN5L8usLLxc4gpxj6fZg9rnBOMx2FbUXYdso5jJcPEFmbra9uoDWL+JYo5n2FE
FWVxlGBEYT2Nb30Vxiz0UnNxKDsRlodU2sNU3qlpzLjUP9lQ9Lx9VG6exTwyhaUA
7GEXlvckSpPZK0fkZHM4eDPXTa1iKQ9ml7DfSsZb400UoAxMmf7pvQJJe5SN3dQj
lNpe8aQCwWw4c8Bv55DyyMH3zAMB69q8Gc0pc8ftWnzq3SlNyoar9ZvnMPImP5Ey
GhNa4cbi7wmN3gGtOtKnudLm3k8MrFwB0T/Igou++bEzONLyz2bciQ4AUK8xE+PH
dJK/060K1OeSk6x59j5R+Bn2zMAJz0pUhZd611UYHgwIjJOq0+b3CRf/NkFh1j1o
VmkQv1T4KYqS/MfiRzZ6uN5hxXd7Y8pjJiQIk/ezS8+Np1ZYNJ8nqORif3srtDtt
dmPOShqwWQtF6x1tbiYRaTQVIvMq758bcyMJb6FegSxk2yQxuoxTUlsm8Lc12fHg
O6UZ4J8S5uZojblboOLJsqxfo28+YvK+1PnUrJiwfgjBdsMNQZ1MMCuubx6vmoRd
d8ARpl5GGRTsyudXbY3AuAZCoozfGdqN7XHO6soRCw68QCLFcIwp4n3NY0V2iBGC
L+lXxhO993E8zUnMBg1189foaQyZd1De73f/763J5ivikxGZfnCCkGWB2QL6Apg1
VNLhraOwjpNfkN8/f+I2KBxMOKOrTba8dYdxI5ObinAMjYxyo9CQnSKYlxoLDfnN
Jv0WMJN6svAtVswdjUKk58jqxHlnDf7xG6RoX+rfXzqsjphEv5jef0mBZUpFeuDF
JmkGyyYYDkjXV/qivtNyiWS67Au+irzo8HyJReMJOU9x/bahJOT3jLu+u1BRGc3C
QDZ4Kigkjm4xDCM+va0zOaVh4UDm1gLQ++v13z0bS3ZJeT2yeGUYyihKLhEdWpdR
Wlhondpl6FPQaNlRve+d/zmMUQBhTEdBkVmXwEqH/iwxeEKaAHynK0mm6yngN/Se
V67WHYVjFwEsnuJl1JuL8RV0MPEFT1kBbXW05PsiA/5WCC0d2G27O0tAhlR10gCJ
6eRyoDpYM3dpRdDzGxWKWZJKSmjRKf7MnVneWgnnZ/7KPqqq3IqNft2N2hNUWtvS
obK2iGPvS1tC52lSY82ze3IkRglIom3Y/L9Pet7uzJPpoU05NULCOsEtm4bSeJ/u
R3YIL+0nkKqF0daL0TGKsNznW45fvdvkbQcs21ETxlrGqeL2oWseCC5S6zOUEZWe
S2M2LerTkB1ggg2r4cM2TjbK4nlC0WBl/BnPt9VEAs9yK1sV/EUyymOWvoWSoVPE
uHyZJFJE3pLM0p5LTYSMvAKRn0j1kgFG92FPGY4pyPUzUxHnaH43bXhuT/bB+twB
ZqGVzvNf/wmehL1rHPlpSHoJeGb9jacYzWxauGvRwo/sZEWKxC3S1n6g93dBSpMW
w8ItJdCB9mtMkgjlrUmfvIEKw3GqeNnbApKuN5kOb5qhtx4PMuHRUYhmpbpHF2K0
OjXg8E8FiRZ2qWI/oBGLbH5S+OuiXYXpuduKthHnx7CMbhw+fLhZT7bYdOIYb6i4
XiKRZU1GdTyhd/nRN8FgZZvqR7p2KgpB6gb87w44iQhki+TALS1Tdy7owQFb0teo
8+mUv+LqvrGyjo+0qUqDdV9D1rzVYoJgDssbktz7DSNbkkSZST33LkfWQaqfvUjh
te3DgUggaiNyfw6JbN2fAlKRBjDpxlAumCPTD9/bY/pfDNy2rGSmmIk4zu5GrTDm
UHIpRNc6EvbbqUlyGorY166t5mB5l2FPj97QCSXIVAmSiaaxYJkW+PV/kSFEiV2t
Ah9weEd0EBSVbwqJucd97p2OF9I4O4OIwAs6UdPgZqyEej1PByl1R8z48Y7Zha3S
CriPSAFeCtzyR5HDNChdnesUrDxFNrSxDm14t8X1c8x/eVP07IDOuiyWsH7BvYuu
UB1IkZJgnh/ZTIHmsnFJwjjXMAyxjUO6jlIOBtNl60MOpq4xc6bgCTnDONBLKFJa
WPkDcJbUWRLNDVIphSydcIO81/b2iMF18q101rnOb8XVyz/O8Kmm84OMWPY2e82a
+LToi1CoF1tAPP1ZwYzF5h0acQZB83uEFl5k/OGE0yK81NfDsfu4mOY0A9rcb4Ec
2kAUsQ14Ld8Ps3y9UnwKd28ZOO9cfCn2GziIJB8GK7erhAWQSq0cjGT7q7sx141T
Rq44AsqI/90IK8TuFDHVBBuU6rBkrVlDLT+4Xl3si5l6CArA5FEj0u9rsQQnNh7T
dukuV+5T63F+6TSK4UkbxspGwX7pbbfFdo0vcT0l+lceYjA5hdLZu+70w8Jkxv72
ylhQjG6WWfu7z5GnPBcabe19mwCK1/Cc9jv21LMvGY2nlZ33/E2aR9mlh6VnbuWY
ab9Zt4hWK2IEi25TZysh24zZo6HwKhmYCPZ1YVRq+6kiPdTnAGmQSji1ORgBNUkG
rubsmMfE2xllj6DBtfxrD2d67aYc9UTVQpYnnjm9RqeJgnNpvMOuz83lAu5oZjdZ
jR7a/H+JXsnRhgUxVhH0e6xvrWY9hSayYoHm4KdIhLV8wKA/u2fvVqJ6QQybEcMW
GZUnKR/i7OzTNEAz1oNaAKgGHv/Xypnh016WUAwrv8bZ7fFU1lQGQPz6oicdTIyg
KNo9iYASrR3zZpIvsrMfkERdf+DodGfossRKjn3d96Qs04uSdi78kiuI9CmDKXqy
se/VwxPtOFvdylMR1XOJNFEE+FoAOR+WfFITwpddAmg9zEr6oqKAcc1/7198+z3f
gRfOZkVEPypBe4Fu3ElaQIvf+eD1S1E1Ha/NmYu4jQNsB0n1MELTuf4C6nGOyCuE
+5RuUf0PLlV8vun1TAVhgXWS5aZANtzY6eoY8UnnrpjvWyqyqgyKU11L2Ls4ZP0X
8FtMyJjRAGz4foBPmzbZ8AvDvEwqnmeu5JKLzMEhvGDgrC2zUIvcYZBjB10oX5sY
As3Lef0UkWqjCXrvv2zPn1Y8NUpL4wGoUZaLe8Euox6kE1oRmIEeMzwnzYs1yHR8
VqZy4dvVmM3F3Ay698pdBGU8hYeynazIm1HCSDg3TugFfjNyVDdD9bZpzM3GcpsN
owBo3LBJSED7ikRQAxc91A+8B5wrnurvWmbLwK6Efspdipzr52Uuqdq+CvS+4mHz
2mvcAdhYLI1cCpdLSKOigYf2Qkl2WjJVA0xYaWvz2I3PZFD2K2XAwXfuZkfUA74g
j/ITxmVK2gQJrASikIcnQ1+KaO+vjljsWH+iAa07RBp2Qya/XKz7RpTb0kWiT8yp
G4FWICfczkIBcDc6wc2ETQ+xsq+6/tvcjSl37eP1gcYVaITaMBI3Sfi+mOXQ00CA
ySat4c0rrixbheoHewUoQXSid+fD8fY4hI377indbUw55ts5Ql+P4rLckBJgwSrz
D5byIKygbwyxeeXpzFllzaw5FRFotloOsHqVZvBjpFgaDCbYPeOBVyO7esT3EaYZ
j+/dFjSoJAEleKfxSprJJiUSUWtUwdTSPytdieX5QPWnaFdvJ8UkO0YhxB0SKSmC
wjSLR4ao/UuA+0pncZaNtO6doX4mp9KhV8f3tYOZgFfMugQ9/iHaajI5H3gQ6wJr
s3hIQ/KDTbI8jDS+fWULS0BWrG2Uuu26wt5Bf51GB2/6hSSQYYWPls0OVNvphDGR
o9ILZP2J2hl6ccQpjEpWoyQf8ll0AkPJ3Y7jGwYpGUCaSqE8PekyxE5O2Hig4vqb
u+6QVHUceBvh4UeZFuddUy9AGKlOCRgMdwCGcbUl+OqzKP8yPFB1zb7lmGpz/Jmw
GIv00UUGbg9UYIZjM0NATyqRUFjrivi3mKQz6HSDNdt446H1WONscDVcBdXvnhCf
7jUuaM3CCNZVTPWi+H7gV1sXJDm51+bH2i14laywyepRmSKr9TtpDUXJOXp3YlTP
Z7u962x8yXUxZ7C0T45KC3L+1XyxAWltCrEYBhpE6ZE8Nvf0pIB+LLvHPwtFFa8O
WwBBeAgTerkh7mPAzgg6RN5e1iHHjX13h/v/c7AfhFZjUIPPOunfDHkgsfo1+qT6
aEYmTe5dVOkuncvRikgbGttAIXHS1riY6HjQ3G1Xb9AyQfBqOuYbNY2EKqns6BlK
6iEfoD2336l2Cz/vR36bbwyxav5+A2/O4voe8LACvgQLamDW4A4oaJPbSBI4Rogb
3ZXjG7zJeg+mp7LMozLh6B6wScVQoUsbKTWxeBIKZ7F7YrkdwETGo0kTiuVH8IuH
QtqIveTVzIgMZPL8mJPSNyMvK7jC/NZWDdVFXTyKRHTR0Mzrhv3I50OUdVPVz1EX
0P5KRC4GvgS56+dkkM/883+UEUBv5tk1OxlETIyUEpyDrk2npe0zS/ZtbHMn+S0s
HihZrhm3X+SoqGAoueGNuiQGwXCKvh21++gOy2nEwpX9EbYQ7LgkvqoY77c93w2B
+Hc69zbfxhuUseOcu/ABrRlUSHZ+M4XYp+x0xdjch5rH2oaTGyBXGZwcgobSJdBc
ECozglZZD+a8qIWpFhFZbXipulY0NAkWxs4s/iTTUJpv2NUqygPtnU5qCZHcVPML
w14YacPtgzf0ztKfM+Gu0zpdNH01f5p1zgg2+azPbARNWSziJQPrqUZ55jX8NtwR
3pprsEH5lQpJqyEXgMeMBzMigdf/1pJdKqfK6R/oUg+VX+Vsv+onmoVTTByGiis5
JCQMWAdip1O1SHvm0XqBgaNkmZ48UblSoR13qgDg0nw5z5YGDT28l/q5qvySKCiX
sAij5DweY+ONmtm3qVqSNMzFjdHKwCcP7/MU0BpQjNBMv+VVLb/ZQVaBEpzya08M
ik2Vf3Iha66DjJfKq61H6RQZUj2+AwZCcw45Ufq7C+pyFsQlKY8+IByex8ENR18g
IrRVdHofAE76TIOY1zS8mxgWBXbvsLtcZCX0nhpm0GHkiWWjYYOSq8gN4psCQVRn
wmngm891kGajb59swYwnidifBm7vnEM3cQ5mDMyXOV+Vj0Ud47xRfw6q+kyzQI0i
UCOiP3X/NOt/2eHRupT30sL3blwav2exL+gBEiGcYifLuS4K92s9iJzUsmVs5Nqj
HytXlO1DAD3lx9DPiVb1pYnrfvjh8ievgGyZrZfVH2Y5+lfBSTVOvZUZiYO3OTMU
oumYICY6aTmAvS3ZGp0AZkeGJTwEY1WeNVccUXCKb6C6/7xKfuVTC/tTLHM/ygBi
jtgTuhDq9RdP/a6U2KKoTi5ceFHw8MRYtcjzlvsGZ4yYrAILdHjv5AJWDpdfrf7V
yGvYz1pWfdY/Isi7qyOAMVKcBUHMBogfVn6f1tHulfC61TtuVR/434p+CsD8Z+LH
L8D4p+IOJkCjZeQEUumi1iUDHMmJSnfN9XdC7nZvGg6vfs6k6gj131Iu4XbpQdDJ
rIBCST4L62lmipixJbbSHeLINfHP+fTzU4W7lVLRUq4Nuq+GCIpgIatNObPz7jfM
g/LXchH8k9ZI+dEAxqks7LeO7XBA1xNV6vHzNBg01TL1AwU9nOlDM9tNvXo4GU7R
Ccb7278gCykhWsng1fJb1Dxjh75j4ycbFyBTc+eYIBnH3eM6BMKkDjlhpYvpVxES
BriqT6RrqcQ0LcQSQvchf13eKLNRFwOtrEiZ8KXUPAI980kugXpg//v6nVbRTvbK
1V4QJE86P4KjMG+JrZxHte1Rewjjic65u85LEqfKd7GewviD5Dx8UdIZeKMPdFj/
16RaHVMi6gKaX1KRwUL3BxrpssRCdq8PwiQT2CrMdrW9z+WO4EBGEJfyGhV4SX7S
nZOl2x7Z3tl334HUwA5GSyiJ8TJj7+lqEJdo+YQP16YVO8eK0pzG7uR4OEDONGxs
1V2NxD4Jgu/Sw44M73RwqdD9MxbP9Rz15q+1lfqg3cg+Bm7NW6WHw2EDcVqo+W7d
Hw8OtHXHSY0bSYf4qa4xzSC7Ntz8Jv4Bfw7HHzRJIJ6MPGEDO+1wrTyD6VOfyUWm
bRvnW7EJGkIYcu2Yo3i6e5yoQoIPjMe+kxpH3VJAK4n8IITA2VNwDVtfZj9+B54/
kkEhFOosCFl0ey3GO1i585n8ocXU2vAz6Vc0P/hRdF8iAauge6avRMEakJqETL1J
rc6i40KJnCaEQpgZ+iVHxgzcMj3qXzNAGpXufZZNOcD+2ZBwkWcez7teX7EjbHPX
Gpxr3OeAxvfSgli7IwNsF5sq/NcavshPuF6udTEyd5lJhQ5rF6PyUFTeOQPpku5v
MkYZr9QesFS2q3VJi3HQh+DecephvOnKnCvIeOVlMTFd/LrDTiSEKKvpKvPv6rq7
B7UxNr9pHKuo5NRKgN1Q3kovdiFvO0qId9AH7k9maBH/9VSu741zioU+q142wf/6
dm2ipFs+FNzIdYgck1boK4YZ7mku0PK0ZJA2JBUTYqnVKRckl/8DWS+V/thiIEVd
sGdA1xvUeeDJT6FtxKnc4xNv+CirP0mtRABIkW7cjg45wkMalPW8MU+PnrueFjYw
iMPyb+C9F9HSTe4QsdTSrI724m1mDyJuE3nO6TyGY1KZ82RdUKaSBr/k5vJhlEeI
loFm5C4PtLk0G+UWs+8NCEX5oH0KAs1dwF55CesvbgoxMHLdlF9KJjtsWlqw2CXE
LCtZBEFpo5m4CmI7eKfAiBJa++Ki97xZSuIAFuIO1fUms/nj/imiC/rzTg6FMXKY
XoLaGWGIrnIHKcSeE0uQ9sDAruZbdTxq/TD4f45V1XAUNyP0u1L5Xw5ueP5pWPjP
fvmZzzx+zshzQWsCwdZMZ5g+Tnjf/+y9OSiJQHyV8slVsYRKpJ/0Dee7X9rc7eNF
0OBea3jhx/NPY8hf3BCwhdUnxuSMz2o8TUX5qigjrjtKsjFfn1GiXtly1LBV4ech
tDhuJW7r9V+5/Vd9z2F58n+DqUnAj8v33yluNbBBGYG7x0GX0YT6PMRgEcb82zxC
/jt+LdqEKRba00fW/kwZU2y/2FPBVQ3JFIE6nRhiKAa8iBREt1FScLf2tQV4voOR
TagLh3UpXVVAMawQaUZpfhTP1Rp0Pa2Qlaw1gxQI8xfpUu4MjUSGsgaznlyetxYv
74FumtgcWyOZbbJIqkLcsWIV1NjLm5y8/BMyu7IQpY1yx5/Viw54bUkxeqw9GHxT
RsOnhLaBH6Mfg69z1oIDCGtIo8rWMrMK2cifIOJIuBcUIdgHGtRL53DT3AqUBpct
tpCXt+aQYzhgfyudQDpb9ngk9/IajJqsHFMZCRJ7Mgg9ojiAsz+y0E0tAj7uvuUa
V1HcM8r8TOaNTCUgh5R132dPPZVJ3a1Y4J8q3JmyLKF+tjR3sc71kBZ1QH6hSOMJ
q9ZWeT1AR7mM/tHH9B+ukDGz1u2Qj3EwlFxHr+BAKnTCFceZAnGVqJ+6VMTWdl8a
9fEiviIJI/89tT5fXII1CafIGZftmZ8Zv6vSc0G9PF7K26GmtfKzG9m8JZI4LcdE
ksv08Ont+HnMYDB88OzhQ6zXqguaVt61X7LZVtVLxFVw4C9Kh14tdl0zIeJj0ey5
3tVm+eP4cPnfllwylkIdGFcuOSzGwgR+3Kg3bp5j1hD0JnjvaNW0CpNInJOCInbW
OM7cpuZSClmM51ycWuFIVQtR7RAmVwU5Jobb5HEngTokkiqvuiS/MGsWb/FMGBOg
BYUixRVY/F/NTYo5J5d5e5nup4dl0+s+bGOV/9EicBB9ZPybKvR2o4qloRR7vhj6
F95AMxhF1aL/QF6YWFzPW9vCgSCd/Z2yViufqNO+D5K/5lbc71cH5UfVv44+OKCc
Im8tfCF1xjClVoyAR9bOPjSzNMoeSHBTUgkbTRi1FOwQLZttFeMLQ2xFCdwbJ4Iu
eEdb1JwZEwKWLSKm7sqSxUJB04r1DWNA61T5Z77aMqrAqI78jJVR/HnnJw0BV3vf
nuWVPRHOy7EYG0IJYzqbPRQCWOdHKRbJGTFnebLp3YJqAhYEaHYtgCHYZQRUqiDO
kB9WXiTp3u9F8jm/xt0FwMx59JXZQNYhATEk/+iMUwXvfSf3QdrZkksr10KgdIIV
8ozqJiFAHfQViPKsmO6GiVm+6UNp1KoBa5jJNyTDvEZLCN0oH1Y4+DWHZUWiHQ5t
v3o1Az1v6TIYfi0xzNM/X5cnqwyJytzjYtSFWQIl5o9JGAcH6xgcDNS1KXrmdVYV
IOziSeqnq9yAZkvXoOtWBXDmYjTwX7hX2zWjh6a1k+5g80ZhlL9Tq7vYAipVX33U
/ejZe1gJX5IeL2NHLN3K9qG8+iMY1qXHLYUl2Q631f97YCrF3uwVpPSy+ks8Jgw5
ZmyM9OtnzOUYiJXcoEeo4+XQSRvXG+DLrnJhiz3qI9W74pdhvIcAO0ximYZWs4w/
20XH/aDS5VgZZyQt4sPVpZU9jyiuHi4ghJCiK09e59YrrQ+3SlPrqoafL0lIawNG
5xYWODXbk3c3Wlapi9rXufzVgM8sXlhXl+6HR3W8FuL/2DpO6zaPU3WAEqXQmZ0N
quBLXHlP1XMeS93UJid+xuZTaTeY+VWfhZ7uZygS0sobz7bSVmk4D7bz1FvM3RH0
jHflu+zepBovrm6I7vm1FW8QnbDHJ0Xxa6oZeDIKH3lF2cDRpB9GYwBwAXQuhAYy
aa63IQ9elf2EN3/LXIWGj9JX+zH5R1cXzK4fdxjNFFPW9n+bY711dUWY5/Yir3dy
Tel2lpFzutaYAxRIkmERefujyfyZATD3sulmtrDz0VZRF5jlFV76Y9/DftoRFIiB
GqMufPSXLSdhXJ2OLP3ZbsHAP/GCF6KxDjwWUrpwUUHQIbpnrNZAUKW0FyjwJcjF
L6M4rHnHlxymUZs8W8fdHFivrW6CeZ8XyLjQqScfm51W7SCjQzxq9wUwJTQcLBF8
/UiyImclVn7lc9/aD42Ju61NBmrub5eLW6cO/GrVzXoKPyA4iFxjUj1THPHuTARX
WF6ABYydZejPXinOUP+P0Goxqkw7vT5e1wIL/PuZmEbGJOxGFZRRK7JWFWNtxcL2
n40EhuH6sct4YaCf/JimoYU/eacQwCzgaT6MtD0PygMHsu0F1IopxWtqPgI9/3/E
0LoZ82roxj1z03RXYNe/rXz2aKkOOiTgoxxfgtxuRKj1dwWwKVBj8E3CCYj/yZDm
O7BZxr257Bn8Hi2QckYASKMAcaVGBORx7wBSDT12JdkvqCOimQlNX8zR7TVM3OAp
KFhn68iFf+l4Ezln9gQjeu1MyU7k3k/9BMZqsgCa5RcW1YokHpEF962HjgzG72J+
MdfzQTmZu84OG660Nkep6qAQy5irgbaFkrP4zoqshtNoUmZQBiJggbOgtshGSb/R
hFJn5aiPxqJay3rwuRoebRLSwKuhPduZAVApUtU9jW60wJLbp3kRs+lX2mDB3qZl
7qo5m5P2ul+LOwfAIygg7UEDjIv8vD9F0rc7YjF8NtVzto+gEb1nNRf9ftQ/9+ey
28esAd6WghkVzfosUhmFfv/ItcfpMv8pL6KgrB4ebxxWjEUf7Ug1tA2fVVuCJ1iV
qDbdKMXabhHE0GTtr2MMYkbkQ6u692VDq0CR9g8nHvuzH0Jy7h6kTnoEzsvjkp7E
gxSt9BLRsv5W+rj+KSLW3t/3iFZYDQAO6C9PEWgzJ/KZVJ6JzJ9MYGzNc1cWIn5t
hwla264NbacaWBYMH5GhUGsCLjya0kmiUmtu4Y8ao1YxXisEa61HS/02SY0tLLm1
azS1S79UyUvQ9ur95iRd7wdMuS3VsOoOcHk+65bbfzz7+oMYz438ZX4wK2K5mecM
JyPaOtHjY5gaUFa9vTsgdGs58sqpjCzk9SAA9QrtVpM7OSln0f6VtDuJ5LYR3vZp
fDawEpV11oLpyEUJ7tuyaWbueVgdfCmfOvbQGR8srGPaM2jBc64OMN6v4wmzl7/w
Q3wMn0MsznCVKdyjvzvotJ9iO0kK8sybVtdsWtOh2FmRRb69UMh82Rcd/jvT7Pa8
KoN50oppT2cqYN8ZsA05+BWlAvLECptNZgJoGQaB3uVBJ66xhUngYOFUxGoHWZme
K9yCMCwfk/So3iHCh3ltUatYlKd4GskvVL2Bp92N0a4t7klAyyAT1seH7MfZPtRs
akWwaPqCjDjgCr7GEjgArRjkuhOmn3HWiwawjVc/iojTeUODqsswC45cPd4Er78+
6FfSz8hUGdEu2AqHlXOtPaMAvNGtndtxKoAaKeE+YMvkpc0ktzCR0+GPMIcAbfov
2+fFr/a7qsUh0HqN1lR8pyeBpeoxPdW+ECsXj6CdMhTWpmFry/NrRRwxY1XrDodt
Xoz1Es62/BJIiZaHKprNY9K1QZi5Appu4F14TUUclhwBIXeS0gSNONMiYwqH7qn3
2jmtHnQJFDk2zSSjVpklFwG6tWv6qicDzAjvAo23jmzlC+2A5Zn5ZVX9mDrLSfEj
ToZLAvuvJjBX5/9D3EQUb4ktTyY9kg6KH4ZJLPSz7p161spoXoNVD2ARGTUhRmjr
sF1su3+4O1mS7yGiMbi0zy+rMEisJ5vTG6mcn9R1WgWeKpNx+klBkORDydHYryJl
8iaO9XotWWr94Bedbr2WQIypRtjx1t/4uZXrqsbUz3Yvrc4ge2Fd8JN0KuLBmyAx
dwG5Ukt2I5sQmB05c7q7Ku+KtMYp7XzIo54QMldT6asE7OESlxGDcSs4b4QxJFUI
DihxjDcFt1KTqLsUS8FrdYPxbzCWh6mpshB6vuTqJIIJ2GbE9C3klK/b5x8E0DeG
vB0m4I1BpJjMtzL5DUlZDnw9kN1JbWh0sfRrzsz4bDaToGudywsUmznPjTLN/knh
QU2XjTkLOkHLLKsAiOhpCPKgJ74RA3pmb7Y6g6zcEgZlCfDwQr3Lfu5rTXBTrZKr
f5cr0S9PrcTL2w4uIOf6Rqtok7uO6QAVlTTI68xFYyGsOmzGe5DHtaXPwVdNs4WK
WTR3sV4zmQuBhvmbz3Z+nVH+BjWW1zHemilxOubWhH/gXiWak6/tw0lfpP31Ooc+
SEL1ze1TTKuqFFKkJQCQiVcPVEV93+dPjut7mQNyo9Zk/7IyoWTxYTIruuAKdknM
e0EG0QjEVWUKiJXj4BcddmhQTnfR5vDy7gpaGJmF9KFnHylgaEL2W9n1HRxMAzeO
oKbD8DxQ3AJkP/SxDUfNffzGlflq+ViG+m/rvhFODt3W8g6R1Vy03ckIXlkg4BBd
h6MGjl0sKxNKnCEgAAmHaBDd31XPd9DR90h9UJgqd2GIPxPR0ekOVlieZp1nZArS
DRsfvI4k+KJUBTL4QhGeych41p+jAmDZrbkkjKb1s6+EIR1JF9KWDh+YnWVsZtM2
Sg0hvNavnXuJnnC/OvxvXqthDhbfDOAKn0lqUP0Q41C5wXo32tyLnZThZRsRTDxK
RUcSgwB9aV0V8ajialrh0R8Tw+/1f14bjstVfV6dhczpMHFfbH6nJR3vHFqvpcQx
GO5wwUSH1taFaVpikobCN5wNHW6ZQztYzhwLRute4yM+8dcJC8vWzoFxzdO6FYQ4
pT1LCaMI/tpt4hvmQBHDdIlXsUX4eW1hPWzNqSh/c8J3wtX2sUoFJD26xhlKJSdH
F2XiXy9wmyKhbk4EL6WWvyoYmzVKLm8WNXVCEs0RKb0ZBCCA0ICUAN79U9BR3tom
zKZmaEJ99EHddknxFpYL9QvESGU0a10O2kofqNMLxDjAY6LldXCdTmbLpFeke4jL
A/ZnPoWe/g9yGwwvo0HdmQOdotjQW93BPSAYuTSdNULfeoPCoUZK+zk57z/yB3h9
wKnH3BXVmsdzCTnv+UR1BiRizUa+Pe/57s5WIEzC4+AA1tzhuNAX74oFqgt0tpZy
U2Wmx2ysD21NMq0oisbRYIwRRjM1LeC/jogMOtC69dQzr6Y5N/vk4dMbyGO+0hd2
5/AlzD1BybsL25LjVTAKkp5HDVVLHLAORfvVONs3LOGechqdNITF3VYETWl0U+nh
0wJiNFSvQor9fn/imeZRjVsklr15b/Qkf3eVYUo7IKaJwGNgV3NsTiNi2yGsRpwR
czusTRVuvFBiJL6mv2DgJqyIrZd74nxNRAyBPKXyc5PillPU45WW+50irDWBOrJ6
d3Vb8CDj77Sir43xAgb9ohFTTqITCqXC4k/KeamRadzyKE3hCh9xOpYEhjGC6RKe
poVCzUvheQHSB2fgU9RA9wibfx4gBQyDSut9BatzbzfTiO62G0NulJd4BkNKy6BL
Y6N37PyhAADg0R3MlPGDjPwKGmmK2RkINXdzYcgi9/WYwVtd9uRxduBg/HCZN81l
G6oFo4g15jfVr6shuwP2WZ/l1fZgSY0bhN52hY93uhdHWIAnkXeA6UNROXfEFHMI
NE9V8od5v682x/4lOvIX0NjhM9xMjo4gvKfpe6tpp5AU9CPOEz3VkaoKejiPtE6V
TtxIKvEO6JgluQ6gtju4A+kgf756v4BbEqJeN6gPGmzpMkP7nbyHBrNSvP/ASlvg
l7J/zNAZHhWzT8NhvTmrBA4/0mgU1Zah+6rQcQ5H6mko6ZWh2O9V6U3tDDe1WWuL
4N/lQ5ZMpSuoKyyC3rg4gauoF8fr5FwOVaKs61jLD3sW9hFYhTueOKjyZNXY03Dy
dZvt1V/XbczVz8j/e2wMJlyG+b4aFRuKyY4a+MSpQVAQt/7KGqGKlLUoX5qzfr97
+Opa1z4Rfvoz4KdG+euYuZisgMzo72VID+DqS8Z0cPpsDxelQAmnta6yZsng1x6O
aeoMDA5jpSoncG0OO+nLDFPUUXyrEPovX2SmC8ppY03mgB9JDSByEhi8EPKazgFi
wE1pKC1O+ou4AMo1p/3BTgMHqeOuhT5WpFkALNY4PpPEl0uolt5YhxiXRHczC9HX
Ct7KPFSEZ1eFP5ExJmYqTlyHf9kpTb/9yJf9Rr2GBYHtY6P8sArzj2ue5hkjL52j
50ddmYffGIE4ECuz9rVM/g1yoWe+qJ04/iwFlBbXfnVPEIF6SDvIAuQbJvIXaSVQ
nJZ3tLNa1wBVnJ1jk5mTmbhKUTPBn3UNdDnb88DHl0XY7NaoSwhjSDjaXgwUo0ql
NTHuw50bbInY/ndEq7DMllCv0BHIKj+w5q98t1yjrKecLkBrYPoBj11pynXTrvOW
PfpRDJzqUBsS/Gf+B0ZkbmRmwZ9CDv2I8ZgIF41Nt09NLigCA3+6XFMnhUxUYoaA
NPXbl2USK0bcQoBtkTA/BtKmp0vuDSpFZ531nkPX7AujTDwTHx4RDyiyzveHZg2A
anVUx6GC37R4zOnYRuP14iQjudDPCN9h9u9eIP0DSohJzeTncqz9PQM5KevTFH74
/aGq+NFUGD/W/MMVVLKstQqnEk6FBvjAESjy6/w/e/xP4eUdj0SaKDJMlbtvtgYl
4vI/oupbxAQq12S/ZpNUr3ordTCtsb9NvYbLJGWGQquKVK9JfTfk30c0rWMcaxgA
9EzPZrAwlrPMla3JZocqhx+kjs+PElmT0++FS2pkSDbWrMxMI5giTDGunO94W6zX
e50N+memoAWxAv1oisbgBoyFVyrrjrBq+8TbC9tkZldD2tvrifrkaShBMyevXLW8
sLG+JU4lGbq4PyVJJjnacVEWCCJB54Kaa6EJ3vCi7zODKCcluxB2pfTVRJw9Y0Ax
3h/F8vLG+RKSHBiteP2ZnvKSN1lwIVkXJ8FgmfMI3rba3Qn7bSOoKA3cZTFvh1mK
PU/LfO86ZGCYz1eGrNZ8ETu8+CKqUMCiTStFk2KW3fTeeoNvskj0XKNw3YEbnR8d
gnEB5X5Vy/4T21xGx8c6Xud/v7KQyjGj82a8QXdbMM9gDHECgyzhqXt3/VmFOI0G
o6A0uGftmzBdN0hqGujI6o0DHbwmFlds3KBkpKfYLZczpXn03N+iLyvSMzW+S4zi
ax7K5xC+f0n/qiAOes10oCVpYgvSXa0lMzMPsOKSoMHq5SyqgnJ8whfdFToHWjxV
d8F+va6koJFv+TxaroWVYdrLr+E5Us/HscgHnQGSq+E4Fy/jYMJ8JlTnCseDPe7y
b6EZl/aGxgVH1Go5HT7me6IXBAUDXKB23Oz7CPUGOw6T+AkTTa2+ROvrzpoyXibm
+1t+mPbJq2RyrHuH4zXqRI+LmhNSk/Lfz7ZKDLu7BVkrYEVgu7ODcC3YP0Y44uxE
2d8Au8S1wubuYvmUU/o2Iv2QLHL4eb91wBicLZvezUYDaILLFQNG4GJ/yn0j3FpU
cfhRlgP8D06YNMAaXeblon3bKGCF32e/ADS5VSKWrg6BKPaI2RQu/mIyF0/Zbcbi
UGeTGGuUVFgAW8OLF7YKBW6mK8j4yMMx/P9WlcSLCLp7y7lKd2PyoWsenYbD8QG1
OCSiJdmmZ4iAr0I21mrq1raQ887E21Wfj01L80ZrP6CnOf2ptPoDB3U0fCJzfw32
S7OrMCJKG3T5PxrlJA9Ojp/nFXSvmWkFCX/1jcikDACjUI93XPq91L0LCji7UcT+
lnqH/QDSRvvNJ2QlBv/mDyu2WaF0RpDcAaTdyjgmHX2h+WMAuufeBFVUvULVOqi7
0dSaZu+f98DIxB1LYiJULdGEQrGVs2Z1Po9ATLdTUiKxkEuCTD6h7o/CVFZaunUT
dptLvJb+j55qM0qTRq0zfWwAn+1ztjx6S9Pu5nfD5WlBVXq/3Icwzfis4ybYg7uu
Y7KEQSCZ6lrjD5hmqlzmMif0NK4yJC1DAhws2ywFQhyeRiXFVy6AjhFHnqvrU2sy
fQB1d420Zg1CWLEjZWZUrJjvUz7SaKZ4PJaEvptooPiKKtnLf2kKG8LG8v2iBwHS
Z+CHAw56b8iIwJVtoUIMOUmi73ILioP8Hl4R0dauEIYZcXSUUT2iKlpxOK5qbUxz
o81Rc97KJLOPnRIvXNoP5O2eSlbK8plp2ItuQ5zhI4DempPKrU53Uxr0rxJXEANt
LuTu7e4UtS/8dOoDaeRmsRLgzgunfwABBCFmZPo0dgJRvzcyAFFKvxR6/nptLfEZ
wokONZOFxE9UhLZKqlmruoVYhIe7G0YCXk0dDFgHVYjY7bzxOQ8e6aBkc5Wm3qO6
7JIqmiQfAJP3IprmK2oFYUelv0/tr321tGmfdYJYpACpUvI9oAKUDVIL8Pn36yb/
ZSO6TSk9XdriF3K2CDVUfaso3nqlDgAGj7FdpVsSp1G3L39J2tGwLdHqDMAAASD8
7WNqcc9ZbxPmnRf4xyt9A+WDhZDfZExDP0KCGqYzGuSi5SlvJF4Yqv/n34oExwqm
VL0jSD7gF+1PGve7qVJsBq/zC/6rMVgFLJ4hSp4f8K4O5g6G62kTDHyjHSsswVfz
uMhXsHZFUfrt77QwTUpNqLPKBUuwVAbYfKe59xTFAEamwXbOFhEmwzUahpCOxD/6
3VaLDxKXvyUI2ksCyOJz9ixGKSaXScwKjUWimO6qZp7z4IfZ7gdoLn8n8QX511HQ
8COfnOd7VAgpJYuQVSOZXVKAjMOnHRm28x0cbOgr4tCV7+P/zQ7qveEAUfzsnm/Q
/wAIZhRcZwGYmaC1XF1FMnEDVfIAPpQ1YoeyesLiXAvVInPn0sqZ793zAqRXbdFs
cXKC8GfLJHnoHYbxHNmqDt/RtXO7dgQum+GEqIRUdsNWao8jcuXFRFccOvge1MCH
TkFfwBx08M2kL1ZrORSxYIeaD8R4158omwFXe0kwgjAReVFhJ62hydX9C/2TRYRr
6rpKprSHyJGWbUkcBj6YpQLbUgEoJB750iJUtjoX/n8syuPd8J0X6TjjPp+vup1V
tklxj+YFkSSSt3Sf1W1zxXhEWrsXeqgCHCVU5Y3HjVcfDJ7JtEiZDq5uw5CjvXSb
mixG7A51JondeeDuf+ED89nuIbymcCQKm1qUr4zjlN2YTSSHnyLt8mPZklWLMldl
M3R8Wh+5BvoFb2hoBZ7m1Zhn24anuLIUzLvtp9BEDMtGy+bUICFZ406S77uQZXKk
EcrWtX/tWJUiVmEcPNpUrWknpQFHBu/D+/67EPuMZUvfZfz04YV7vOLPRRVaUVqH
w9bcytq+VqVPrsDs2J//oLgLgmyW3cL0u9s1N25HFIBjzssGKGUT+5ZZ9azlwsac
z/IHEKAXBilBqEyrYl6BNH2upOFc7y+3C4oNgvz7m0dnSp4Yx4c3unfJWCHiuDNK
s4P5iSHlL+1eS/f58BfnG1Qx0SKzbotv906Dm4RCSd2v8/jqlgi/a1CB9OigfTVv
X7a4WwXqmwAbFlzK7k9l8eg3ITFznggn58u7LdEa+lOePQNexwvoyYcO0gtumjtC
VVxyxWpokf5vrGM1PrlAd0GERPV/3oe664BXwZbEP6rX1QCnIIQAHzm+zEzzl9T3
zmU9BIqHo54vfU5Ge6cytjLIl+EYagAmty0e2KdiEMTr5Yz2prprLo5FKb2Vmq/m
6+WCzg0HcRUhgEnm2DCc3AJjUXxNHNb4Yp3cDGam2S+TPLceMQibg23U8XI1/IE5
xpng7VL4QuoKqLaY48y7+bBKb48FYDe/UBbn29kkbte5NSN1XLdlziOWeq3YKX9P
t9aY8GlB3N/dV5BYCmjO8d++x+VZtdTRSNf9f49nHUmO4asaxkJsQqXy1utE2EYi
yCQt0go/oqnDSjFKLrSpbGZWVAOrcGWGzYFsvTgTFnkK5kD34P+vYoaoyhpeKY4w
PfNP6t4eTZfclsBnRgVv7cadrtibzenF6oQZcFy3Zz+YAdCiXKN5Nz/ge9eveHUs
MwdgVUAZKZrY2R8FQqx9uOvJSyqAZeBKgYEgKKt+px73nYo7w9GfLGiecCQzrjTQ
rBnvTHwvMALasPWBcida8xII99J85EkIEpeWX9RQb1ERnkJ+hSG2OaO73rmH1RZs
v8TyOH1unYDvG5Q+7uXVdV4YO+9zmSbG5GTQm2HHPU5hzck1WLs+ZbvaL6kxDgPl
dabG6pGX+HTVGUBlkpEtbn0sWDAuc5ynTQeiNjVUnusw8ufeejFhQLtFhCAR3mJy
hmv95yRv2bTJljDvxy8Q9U9SxB0qE0abfXlydSHoIenn+L5ZlQXSmwDcPJcM/eoD
87/i7WteqJvzY5AffP+HSuy+Q2Np54Z6VExMzk06+tCqj54TzacTgOCQ86aCjoP7
Bz/QCSv/jl6sY5YVsoMUqFSRypuOnStYycTYKcyANkoenpqYHkgxb7X+Pl4nA4jL
b8yCxCXQg9UjLwK4ftfGxB60wsKQLwlpuJEaSOvyTYJOfFWPQcysNFosh5ZcCYBd
CAgJQAdY7gGLldURkFqfN36bSZMp0KH9KK19dq2CXHWcSvTjr0yWe5hLRPTNpfdq
GzjiI3IXkdlG5XoiZX6M2CWz0uywQZelN9bS+cpk9JxyFecDBpLY4YERBvU8h6kB
pkropfOGgEZTIQiCf+WEjxmX8MF6McnRGw1VWmcA4QMNEddU5zKtkmgSUr+Ac3ro
Wbb60MOul0B1j+JFYb/t8lce0Motti2ZBmMBmnN3txf4Kaeg0xb66wni4uabxUNF
rVAUKf29QQie3xQVrY2Kqj6PG05iVkhK4/E2cKZ/zFxKRDWGFTbLa8+yEkmCmS1V
mE1xZfnYjv7pIPt7/qrmI4HEvmBJaedBpe4XctrAJ2ufmjVEW1WDRuojMy21PPi9
HTSMkBC1BEYl89/D6f4aQu11/2lSlXKfldzCpOaly9fbj0uIRvkS3dmTJZnSluXg
4Hzjnsu/bIOGKk15uZ5OYh+bF43/DOjHWRokHLS7ziqAHWDloDWmv0EwbaIr1cvI
pa67W3t6MMnS/ne0mZidD9cQoTwIqILOgtcarYeTPmmc2n9wMi6qfTYRo+G/1jhL
x55FAHZoVtRf1Yr73wgbjZKQFeRqJM9vKQ5afc0fNF45WV/Bd0XBExjPb7OCTAL9
l4Akhix8CVkJKF27azg3D5xKRTwGUT1YJOedFOt8MY/9mRyuPRZ63fvfvtsUuHjt
9rVfFu4uA59ivV+n1/qT2I2yWjqc3tue0iZP/PZVu6tvXnt/xH9pSrPJgyyHBDJ1
891X3PFT3MBzkA7x0D9BU6Wf9WYZrIBJFgf0Vp3ckF2B1/MUeGWGogWadHN/iDKY
Rph0glJe4rNjRjanTzNmdD+x916blu0PCuj4/8BEhO1NXDnIn5CM6Sz1dzyA/cd2
cYCgLhXWt3FaKvYuRbEB6HwpvG4AP+JP2WrWtSOr8dd5yU0OQsEeC7ftUO2exDR9
UgH+PQOyzFvxZzWdf8dOgmFT8AAe2S9DcdGJ3Ut79dibfWu4kEVK3QjUH2h/U5dm
OjItOLxIV8eqFiapgjo5tI52My9+d2VF2GVSz4/IkEQ7EPOpbJemdXBMVbodl1Zw
TelpT9NZIA+XBUd9fg9lOQ7megoixDl6ZyAOp24cDuyMJXaIZ9dO1pPadRDWo5xi
J1gsdpqud8Io3MYaTYx/TXgw1j9jka/EVVLDPUAXS2xrgWO/UL6Lh9lbkxTC4PdX
09Xj9/yS8eChGP3XNxUeHQu8zH8CyWpyxmmx2nk0BDwY++pqzDOG6CItZvBRo+hq
Lk+hBdeC8QY2JG22p815gXmfCknjgbUXhjqN6LUt93S6qjFYm/gYuNkjLgGUK3p/
XFAM/c76w3ElQfgFwq2GOwCFWAulMPLt/SCBMS3ibztrAT7wmS3WFWcTPJXezGl6
aT3Or52UPY5naPXioVdAF/a21hjzDj+8kBBMMAOUZSdHMQXvDeODGSEpM4gRakM9
Jy1EyTnC/sMYfSgVYUWKz01NOduLnzn6GD1lafNDCNfZfQ8BYCao6cA6EEXmMfYC
I+TJpF1u2u/EjmAS1EuOJGRsOmfRWzfBQx6QgqZEhhN9k4YmEOn/MU5KAUCH+Kzf
37jlcpgIvhQmzb+96xz91m4r6CcoTPfFLKYRsDx/7sYwkGH/TjZiK7HL5nJ5DYTS
dCcsL7WNu4hP0vzasCvYudUubTjPBa5a7xqrFMAXDyfK8b3h6AjHsg8X+6dKxRrQ
ccqfOITvE80erPB5Qx1OQaecK7N3hyqJC6/FHTNfzKe9T81kTjF0SvTaq7718vVi
8BHwFXQCR8EPnDFxj34737XS5i95FkGqD/hIdcAIYycG++Lp2sbqdHK2x3NWEbOL
KZ0bN3J5vJLp26sKKGnAp2blxyk4KeiTT8ZTpGFeN4c7FKZNV35hAQiOe5823Voz
3qXKFnNAPX5K0ZCaHEcVqSplhXZztEvhX18pADPjOA8LEizpjqHhPV2KEgDm3JxO
K4ULp+bDNcIjChoUSOWYKRejCR85dQq68JSO0eeWOHZIsyheyYfPruj/vHc9uy5M
JLK0imo3lyiIe8GKe5kUh0PQgVe7DhmU7eHvb0GWMcCNisPmd0Gf0dCfVF+ckV6R
PiwJPrlMHInnBw1YA2xnlJte9oSJJEk0NzP6m03sfU2HHFe7nO34kUA0HDz6ZxEQ
YBNM0bDxVBCUgI343F7Lm/emj5YNpIm94vex6CdBakn1OMujkLFX2UbQJvzX4BNi
+3SYBnJvwKtWbZVAn34rHCgoXaxfpkC5EoNxe2Bea2TmpWpSpf5rqLGAoav2VZYj
7H1bwOVbU4RlaLsW7KB5s1ph8LMOLKGbo3FGN+cHZ8ZIc+HXmd8uBLWPKCMdqWaA
QL0j8B9YpYhd/KOJgL95FxS4zRB/JXzYU0c6+caQjxDgjHY7U8864xbihSFr7N1W
oMBJNxT9jO+jcvhF37167XSAUO8z3OhLc+h5zeNcHeE64PwYPydxSPhaVtmouHzC
lxP4Qn3To2wFauR85dwFnodv8wYvJ8yXldfsFs612QYFKxo9z5PS9uzF1QdtyvfX
Fo0wMqnbx1y2Jpgz+khXpvZsx5Nzzy/yW2lxV4kHS0hWr/5UyAZrE8fEAbtKxERf
UUUZMozZLvoP14A8UnCjIxJdSMLL94fvSKKzYu3iP/ZSyGgkzkSGhG4PFUpEiXsX
A5lHoRPBqZgQ+HMjyOBul+qBoB0ycA4kEApP3tJCYCvcey2OfOmEdifqetIo4zx6
y/xQHMa5zXrOsAxsOVLowXeKN3w9oi76xeITRu5XZgC8mkNAAlcLqgUqdNyHcWDp
5Ac8c1lzH+SObFukDr5kyywUCp5Vy6mrmPjsINo8GoshKzJjSaHSFV778Cox/R5K
4lXkLwngqbwLNmYrW4JtejrXh0q9EgqN5E4ot5gGyrFJ9wKO0nEWx9KLlFjCkbLI
MRlf53kt7d5dRZldUD/6hynruH7Jtp7dL8mlfme4hOTJxLaysCFnOXdRtF9IPPgG
kkgcN6U9m8tdtzL+O3FS1ejbaZn/dGzFYShizvxLkEsnWz0nsLpGW2R7UAR4A9+T
+L41jzFmFwHXVYvyg2wAVG4/oOq6/o5CDfiowkTiwvuN4pyrF0lI+Ls4LHK6BXld
gg1Q5kiUR6aQRhKdvtzfjbAGzDmkeSNYKhJ6uBo7wLdFKamn3oawOAMer2Qie1Li
QoOpsam2MfreQbbDU8bBFQnRZAq/f7ft1Dpo014rl0CdaKcnuEoY2pMTYRprFUJm
QbioKPYyE4Lsd1VZGtzSYJuY4HK4BBzZj98+O2LksoTWxI2dE03N90TngJVoFabh
RUJYptME84xRR1J+jIJ1R1oFxeGlT20KCg7uZj75KuMIxobsB9t1qjXLTyx3C3g+
jWjzstyA78zu4nDa+bIduZyINkfCW5eSMtAD5VZEnw2xOpsO6xA12v1fIVT3H+Ru
UR6+raqzsPmJz6+ZmwYJnYZbQPdkrv02ILWZptTwgjhcWRlYGtkcDE6jBxG3ttgv
s04pjObZmKvMsTUxxE8BFMZrsB675wTZysEh8LEtszfduwx+dVXUQQ54kEIzTkdh
gTZVn7dH7taFG8mrSUI/8x/A4rC5gHp46iF0DUa48Xzw+XI7GZuTx9H7xnMjzUbN
RjEby1BKFJhvLxTBvvGPNelJCAWJoKgRaQK8D5L7zdYWnRBY9pqgvbmnRcVbFcC0
RAF5DpXBWlNiavD5wVUDrdkX1808OxW+2/HQo1PnYFMoLNZp8lmZ8W9x1gNLBvIS
MaUyajci7jjs/jxh/V437O+BPWcCtrpD98vZJ2r2iU+/K0fK1CfVJMfp3OQl2oCX
A6vD4gaHTHfiNtMkqmFFygXAXMnDM7nps0MccJGzQ4WEiKPZSt5PMM7Xdg5ajkgW
uw3JlBQ4rlGvoFfheTwdP6c6oJfy83JXhuAChRjp+oKj4DKsfkkxuH5KxuO1fTnw
Cj7fMAQS2RmbGJBne2d9lr1hy7DXqwo1s2oidspiRNl5xzUR8y+Pwl00mXr+Okox
ihrUpzhZovFduX08hXPWCteKruXjO9l3O21y/AHr7aou2RwARI798HSQAiUQ2Qdu
WZy4pyQDHs0aGvNTcalGdTum8b6B4JAGoorRKCUJSBe5TMka2CE1xcdR8FNYUktV
p4CB1VWGDCFkXq4JUs24tV0TzT0s/x/5rbvLV/85VuI4qz44bWPefpHf7jpOOkrC
tmgA231C2S/YR+Ve6mDXI0MsGTiV3mHrjEHDeSM0mgjY2BZfHGdvRiHVoazQzIZO
iQoGxV+IZ1eHsfyjJ8AmgmMOHjK+w4Kq7Wbt/NQ4ZEaPy1RpAtLs+ges2H0naADD
AMKXZzcBi6g9XnDwwv4t5tTQmtwhu8bVrYjO4bDc0+tH5kgUIDmV5NM/2qVAXVJR
wr9zsorTG7vQxpGjJDBbW9Gjj3gKf8OSDne7jKE7RYDYhnjl+o0GdLRgFqhEanj9
6ReNYlqfnOsZLNPzTKlqKFpUYujaXUpblVK3+4ItkXIMC4hVBuqBblJV+xL0aie9
udTUv+2yFoIQCqAeT8v7QmAnK4RT1Q0X/uw5jZCVKv2mXX2uAGbGyoFgk1hholeG
afWc0Ew6IB5nHVOvqZrHpYef0yna4uAI4DEqmmnb7q6NMn3PyOv+zjXCJMl2o7WW
kZlzqiPQGlUbJjomFNaIU+R7ie4CTD1vXlIOroRYRFyPeODScv0loQJ5FSPptw/4
ZamD+rWazgBLrj8CYgcs9G1+/7UOOhg7AyZ+xxVXciy7Anqe8PKP6DsLNdtm3JKg
y/+DChQzdza6frPnUs+Dtz8ZxvgOgd1dJsCAQ1Ta9lSBXtT+4PjjCJLCdjXWXk+7
lYbhVlRIF4OFFrXYZHh5dsiR+GzyKBV1V4Pq6N/Aqh48hp8uIxShQcdbnzYapPyH
YVLJ82hAo4hRZznPWjSWas7lDdbBGsx7IfNxZhnVdgWuu84hCEoCRZWzPVV2t5rP
WfCqDrCzRhBccTYVQnGxqxU1umaLe/EQEGTuQgdQW//fz7FjnyfOvXNjtGwrgzbu
UuQLy3A9qtcYk4igKQfg1aq8Ytobc5MfBuMML8YiIFJIGcmHh3F0Gax52Z5BnmDJ
TmzxineYpgHeuY2+pHQIUL+9V18jcKXj0xs/xQuWiwaSUNVRjpfGPFS7xP06cYil
rrOCoeUn47dyccQTrWKP4IxBnMJRRsMdWqlQTtNgdlqegiV9NDudJmK/DVHEf1sw
zD2aXVKW/2RUs/Bsz/LukvrPnYFIL5w3PFwTi/No/1+KVhUABoVsXdSOX3cnftq4
VINxHE9VK1tl4zsQORRzHf807YV7ipZIVQBSvuCyK5myCt6+AmQLLLjYwwGSfxxo
D8OvgfHTWR76LeyIqiCU2eDD6Bbk77czLWKsNjrIBIWMNnGc/7kPLJaTxCPIg32b
/i52m0sEhsTN8DH9cUZtO8rUaLSZGAfwDQSOfNU/Nmg1OZXuBsWvHGRuwLvwR0JR
VjdyUI32vIY2kx11XPJp/BfJthbyvUKSDr47X9Px5FxXf0lq6no5w2w1nWdts2/k
uCtlYvMRbl+F4GArMkUtduGqkIMPQrIz2I4QGV5SvxUt/RJek/34YlrmAdJ4ksLw
wsA7S6WdvFGUxVUQIfuQpPbrrYU/OVrf8SQpvRilrKf5R362AYQX75sWCtcqvLy5
m5Gufr/s9puD9DA7awfFsDI683EYd2hM/7cssHiQ3/E1hlZYZQCErwZkfwr1CqMV
oAH5l3BXNmWTOL8ssCZ148ImkV3hQ5e5t08f5wWRzM50HBaMkTByU0vxNgu+BKx3
yLDOgTm72qqMQKrkAXfcBkXwimbG6UszwsOupnhfmrFry6SXuJEikri2aLk7aRlm
dh14+iPz6G4GehhMzA+0Pto9i06JEKjN999HfN2bjtEYMXOuccyML8CKQJexNK1K
+Q26nWu6CZc8hOydz8XR88C/f2DgKC+xnACRiy+ODoczzvxI3thUwn+Zbd26ZLdE
6ZUo3y2OYy9fyl5EMJpW4gdmt1RV8kzDwnLiO43/NolD4DTmyKUhy9BfHWQd553M
/jXkASYmgsBcsjupr8B1GXb2pC4ttV9FyKf7aCXy4XdkfDDcRHYLK2IT0yogv18E
/sxw3OFCc0zMj4ilbYQB7vtctBpH9w6vAbkKQgD9klKVE4jchS5uwVqaDaK/Lt2l
wrGLiRT8bNtick0g2BmrSMwuQWYhm8noM91maIeZy7IzM9nMVUFwBUT7VWk/wm69
sZPsxrlu5KuYQ2sg+3u2ji0PqBm4OSq+B/Qmu80NmW9e+U2W/auRR+aypeU3HeN9
oYNBRQ0AfCL532A0TWAH667/1CHyaUZvKyRPb3GMPBHPUUimbmPhxZEnQMPA1Cz2
FI/813s1gWgVTjTU33MI6k+FNwXQpsQ3z/do9pg2Tsff55ho2LPqogyKEXsN9s2X
u7ZgcqCbJYOAOzyo3iyLAxW0S34C3qJ1GK0ASAOfLnDbBKAvTEmYiWXOscG5tWjJ
JruyTxw4Z8ObUpJ8WTRsi2xk+x3jRhpbY7UAZnBjMof7ID79thpDmSt40PmsG+P+
ux4YHzvnmziUXkmqtLQStfWQJuUzGZD10G3M5Atj90FFtxVc5ZFNxk74W/inglur
iS5NL2icjgbauoekKI6otq21FUG0eIv6PRa/I+UJxRsMCk4B7RNy6B2g9J3o8HpI
3SW9i68JXOU/sfgHBMr5SRDBVJA24wFMdqlumb3cKTlwQ132+OoTU5M9gCi9IGT4
6hdhlmoYIhimR55T5PZflF3v1OjJkTXc7tXTtzCqeURp3tCCHhGva8bI8ZY1GZoG
pZD/pzLnboofEW5RWiJ1P6yITynozqIFydhFIjP3kQr/jjziPvebAYuGxatlgqMZ
y4XbQV10Zbglvk/owxrW/sj/fKRt1cZUQIfN4X4j/jsSk6SOZP1Z+Jf/oeMZGj81
Goomj1NNp6gDmP+vIyahmg9nMbMqHIypgoXydjGDv/TO6uPvk9gJmLzZVtMsedTO
SnPmVkjEXQg3v1J2zqbmnxBcD8DwlXlXWr0kiAwJo7gv4vMr3y+MVBJgYTXzmjm+
07GjETHjY1+l9570VFaKTTkq7O8e7Nq//AOe+3y7+pjfkGuXZZsbu3g+KhIJJbIE
zJ2ptzAuND58hos1kpij3RV5Xs3oQW7+99Rsw8oMQZ5Dj7KgC99WgQgswShcfe5Z
0y6Wf3aXRKm9svOpDd5bX3E0+JDDB8AtrTjVbDonfWvxfnaAKyTZDIZ5uC/Kqs80
gzk/uwGWuVjqd0NZLWbVTA4xgl2HMWUJf8g9c0+ng8AaYCWIfbhjsETGxJDBQhDL
u0t51ORoe9/IwrPQfu07/8LcicvfN4hUgM+YinNMCEBdKBOIuFdkkZE3fFIdmujs
IenkF9Is1A0xzt3kJZMH9tM21KHMZ9KpV/ZDU2w99FTKz1YN/eSdt3RCA3PRntck
yZFzm6eVSrtbpP8Wk5vSh5oPHlqu0Zf6v6Wg9uX6sVr0m7qRkVuANiR6AbEXGCOh
OA9zGVXkp97XwCkIloweJEqjMammA6L+WsR1JytEzvboxIVWNORQmRofJuaQ0yVA
s823aTsjbkwXjtbFNdi0SVV7FJOQx+9Ps8oMMYYqaHdSBKhkvl/cXASl1sXajID8
ISnKvMPm7SxsWu1ro/WZEaXEipck5GvRyfcFYkJjgtqQ03rK1x3HegoRZOlaSiPL
2v79uvy+bHlxsyPLH95Qc/ngfD9iWmTIhe0aaUkuSLvBkjl8TxequNKGJ5RS1ORW
l3EF/Fcp0OQi2N8HX6F83pwYnFkuSFvixZGij4AR0W7WKh1EtfwYHeMdNoKuCkRL
LHO1u1X77L/d+vzooVw3QbhJHYHf3G2Ai84rkt6qIWa8C1SvnHtLXhOsK9S2m3ol
K8zRsYJNdqSbrFFImpUyAfq1I4ZoFOwj2mywwb5SgCdHNnodCrItg8YXEvOKEHgW
y3iRX9g0xVujFfUp9QOhLwSLV0xLZZH9yW/wRo+yGhnED5K6Z5veigzI0vLuxUYa
67RhdxSWMRyp9nkoyFcg26Tjc2DZqvEMXFV2V5ugd48Lhxu+LCTfVRCyVIl0II8h
ILBGW/2Oq8ODEvqx/G0dLFlg7oOnyCSN83vsDlQqWyM43Gi/fL6Ki/gli0HFgMs4
Ds+lGiivxPbM8WWpRqXricQHCXyPBX+tEzz5mQCYLP7ucwQMcW2HkB3JRK2iTodh
QMvvYXCeHLHJ7xo6d1m5sb9LoO6zUvLWTubhDY6yTKxvoKVvPGQCazJTu1alKh/e
Eac4gGn61TC6X2VTGdvGkULPkoW5zzAeIpnNVxd6SGMSZWSi9UKQEP5T0NOQSEvu
Dzll1z+20dJFpYIxkXKSwSt61A9mbGpuW/zWtRELboLFXVQxet5VqhvJxS8fs0z4
K4gtcwUz7tM0xeheUhn7T900sun8KZjpQCL+kZUyDiKzZNxEtpk26/iimT1ExJpp
r8+4ivrtBdLZeiF1Ron9prn8NXgBwAgqqWSztpp7bdgxbLCmc7P3kMeTKsWtFLBZ
jPu8GxqICwFfTPERjETs+IcShFQdIMmi3GcziadWg8AdU75xseSI1lYxbOfddZFH
7xn/r8Z8C/8CBqhXDit632tXdhtcDKfblKftMDJPV0ELHf3pubUAJZnH+jwGxKd0
sPl3+/yuUSVfDUQWKPjhByu+0nrPdHzCW2IqNdKad6/zAZXqKozgRlyCDy4Wv0xF
0aGNh5AqPFxTlI/Zl3tanVaKUB7zJRmf3Ihy8pgn0LHGkmJJEYcXp3ijm9f0JWVr
rdxbCgHD2L0A4T94zl/90HY1AS1iFYRAxQMv4qxeQuyxu1hJJngmAGxUQblSRSEq
Nx2HcTv/OEYlmX5yVqaXe1rccaYOVjDjSZ2MJCaMOupeXNXavLQR5TvmkbrX62bF
DIHDThvuO87MHWmnEOizStJWSkFC/uvkKooY/USKSUEACvzO87ia6NyxA/Sdkpo0
LGnQ3G6sohfDFgz3DtHSE8uP73tFpTO6+eE/ptRPgZ158+dcVxEt7EvHQP6M07IR
z9eTxAZBPDdHFX4sFo0xXHC84fsl9Fi29Gv6DKOxz9U+vqy8ZDx5rZ2QnS0ZOJU5
vBAt8p7ddlDU6u9CEltmjqsvYW1kM+QfissFCFJrjKtO6AcDq8yYIcV2Q1szjLxS
ufhtt0GvBT81NlzXXxePxbpz9INTxKLKSwn+D/RJvKr3s2JOGfh1yRND5AOlFjF0
NMmlBb6W2qTPiec+wAvSJnk/QkIToh8qczntpfdU4PL2GYs/XztkRvvkthq+nDnX
2HOO9l+JBIlBB/5IW1gsjWyzeC0G0jmo198EIkrpfJhq7/+Fyw+eSR7jk6OH17MF
pgElZcmmRW77m+WqFt4CBg5T+1mtJvZbjzWNSd9W1b2F9S0ydr5YabYfG2O2/do2
Y+Y8AghJ+icebbOpUkA0ztq2wCtCxrhAAYbXCUPB0rUBK7twqczlIh5SwEnRBlM5
DocfAHBLHkvWDvbBAMkkcVR9fH810vN7msky9rgvEvuWn8tIPsJ1Aazl/4/oBiLf
zyXcz/cQEjw3A57AhJCc0D/mCv5OVTVS/68O5p7FDx03cHFxJUveDldpl2LfH7HK
GYqN2RL5+3ZXGXF4GkoUNvaiZfVYmyChLN1T03AF6YowgHc3YdQMXIGBwjyS9wsr
1+LKjgN+nnv9DEl03nZKkx4p6I9ORvdyZeU3j1IHI58f0uVO0LfWo8vSCJ3CeXde
CIeyW+2oagf0Soxr2LBLWobVOnycLz6otOqOaHLLWJJWdJ4Ovb5Yv+70dXZUQfip
lE5d0It8XsT8ocOHRjcRgnL/3zUSSvuoOBf1CmjFZChS7AEE0ConQ1vgcVy7KO7Q
plx807s8rPjK/qaGKc8rBqEziRgkRigTBw0BJvmOerwW9gYNY7h6KpPMZchrpCUq
iteHrWVpgE5R1x/w2vGO1xPGRQNHDRLTzQF816IZIYiz7C0PbZTpYOdwDuItFJ5W
eVMs/k3VoXoCFlI1NDbKRLADiyIH/aCAdnMmJvvmuB7v6SpCXsCZHCrhHWDqncvI
88LvkoSuxQ3u3LdomX10LzMd0QgJCgct/JMn8ct550oi14Mk7lNHUu4n9y8eeVbX
Ss9jlLhSVC1NmU6BnGtpelHdIWlCqJZJDVA6UDlkd2B+YJIZHdzdsCiMEYccbNsV
wcBqLQEI70BqG6IFRD3xVdHY9tyXoauRl82b9fIxZkSUvnzTByVjgZx6lGM4vayq
Y1EHVgvy2EIrmMdthFS4ckjRQL++ir5mWCMOhCToygaZQZ28BcywSeSVWFvBBkHA
y0SyLk7mpHHshAfXzN0pM6jZrDio2pkd0itqBBw2hPD8a38+Ok7rfiUg6YLftqBy
y6vjvXyKRHDFtj+LcUH9LgK1GiRICqMOeX+0E2RkXN8KE+Mm0WFqjufrUNLpsZFT
TTZ/BqNdwNnjOShVjx9GIt4t/UOBDEQaqVjF2UJGcmP3YIJhd8WWg3JjXWKBjoba
TyCuXRiqYoPjmVO3Nqi9ZMaOm2YehZhGxE9MFzZPNZ4+EUvZYrI5zSrZXYqBuUjc
wYTeqHU0GrBwPxV/tCdPg36Ku5XmobNYjDU+ensUAjLod6YWoqP5g8ttUsI3Wnij
c9qSP+GtZeffuXgCLo9nq/e/B89gUvrq7dNMhbyB7r48Z9HUZRCheplw0a11DISj
VMfCG5p4FQJfyFaKueEFGheETytORv8I5yyhGGurh6H9e6oY1bqWaW7Mxlw8LJNX
xwgevVg1r1zJ4hRma7OO0vM2+1VoTakVvxhMbfTEE7eKJwxm+RGaTtmTSILzgfbF
HZP51UYquZudj2LEMmOG0vcM64a4D07km0SoQ+SLywYkzfaciQ/OizqRGxRyC7RC
gQuS3pXiF3xmfr3YW+A6iSQutf4ANbkiONSTPC6pd942H58fOPacO64th6pn8lBL
95l3+3gr08z9F4+Wwgx9o2+9oJXh0/k1J7dkDXCMCfqj7hqmbs6Is/3H2xnbYiuK
dbsQNFIKJTLieZkR0pLMdNpKPWCnGGwnTzl/oY2xnoXtfiiuGpFRGUFZJyEagipk
a9UXcQfg79kAp/Cx0msvQ/7sVpMy5ZvKubYpM6XqKFf5dV8ljsD3dILUf8tJc6q1
vFnH5vil5O1JQUpxIuwqSR+r1GthuiXEM4Bff/zQovj/aNQKMwMt3KmaiRNc8VOX
K6jCpSpjCGdZnEr1PVAXoyo4hFOkdfk+2lm1ze/yJpP1TTMb1fCILWyUOG7g7NTZ
25/qSs/9Ha0OKgL4bbSAc41kVYW8vA78sUvKcYkLFcPTdXWQmT5gKco0IADp3eGC
VD5FTM2idjao/QjJK8ptXPxYVypn1dOKhswWTdSOU4jgCAD1pmSxO3U3w3eQ0O0e
gfi76oIA4SnG7nzEHta4XWuZYrpMaUT+VyxYJtw1hsaVWMRkA96DMsZIngcU2IU/
XPazfS4EUeGv1+0Lq5nnpuvD9PCgNKVMsSh/AXYmGW2Dg4TKn6BUUBET1RrW9zIJ
TlAPA992lAb4EyyqXrv/qpJRYTM8TSRtCcRDGIVlkjpn+NQs/SaZjzDNZOIhd3un
mTns+nGIhaL8dr7+kEHmm1m8YkL4i5XuCcotxMpyueviSX5tun9M6+EC/GVNBTgv
JUF05/Z9Nq1KbhF7xOzBqM895ulJDjXHhLFeE8ZL11X0ZNLgIL1LOJ5iuMZd+2rt
Zqyzx2R9vhfcgaiCcadErrQqgV3g7Ot0nNywzBxJ48bmjSCBRicTFWJYkQgNqR8S
NHtFuUxfBWnkxf6DD16xi1e2RJ4m5/pLuRUPw4D7X/A5X1980GcnFKdA3cLuqL4c
XRw7NweY7/6r7p+jUvokkN9LpHgTTV2kfy3c8TjpA0cafPj33A2jIxpg+e/vAbGT
MuahVv4/cDyfcH0j5Pjh2m2i9c52+lhh9gTEcgVZDlf3bzDusan+yGq6kTQP6YFP
OioAxHedAzGmJPBbxlsP17apYmzl1iIpSUOuuXHUG2OlJT02nhadr6S5fFXhni/J
O0fVhoS2LdDsEbVTzltTTp8U7HzVFbFBZrKaiAQgMVbLMD3OzYcbzwDTCyRNEX1A
WmG6kzBJo4UhBv64WB2qYdePPAE6rwfSLMANKJ/vVJuE3Pl9uX4Mv5sgkzyQsVIQ
NuxBrDajjN78YMGDSxYL2H+qDv5nQWyaV5KVbMR30eS0/YmoqlBQ6Y3kG9xlNOY/
fLQd23Wvq7ByzHxiYL1DhldQ6FKX2GOUrE/Ox5b1gMdbuOojJSXOzpwQgY5aNbBp
R7w6PEJRNmzLAS+cHU/VnfsvLr3YTrZ3ECACpnPPmNKq/UOUuZjmUqwvBlssI5K9
ZoRZqbpO7vfT3bJNEKgRR+5EcYBpsvA7dp3XLjxj4sFO7AtAsPRB+fdjRfFornht
Hn18n36aStXXT1U/rFQQebhPA/ET9VXwQ1GXQ82rkWk//K+YRMTWj7rJWvnBBhoa
5V62aVeckgyrVB7IjhQcmwanzKURJIRO4j3Yh85kAtjzWpHOxcnVkcNRMXstM/I5
deHphizXFVCP3iED172ovKRI9WKkKTiswk844vfk0O0U5UT0R1wZkP1v49sl0xf0
AlEtGF+KcKARzkc4uL2iNLMK6L67LD0A/K3npz3tvd8pFqdwODIVEiDkdH3Y5Nwj
BYTHgcTkcFhkIHTK7GBHljPt+Z1tfQzoRn5csafNgBFTMGPPUHlzeB8FG59WFRag
IQn8pIyWg/hl7a+5dKrYl5ClfMXOdzc2WAQ1dzhpy/jAD25HSPIaFQ6FvSAUfsjx
yeusjSiN/ip5PL2+bYWdM1ClQ7fFLD8NeJgZJFjXxYYY34PVt4APKHTqAygSNTtS
waoDdtbdzaX54XoS2y6c6spwuEZHkiZh5WeLFpWLM7wa8qon2NrnKm/V1jBsJAu/
lloHihkOUskqBKYESI+Fj3sqoWPNTlWA3L/IdLRvo7+/1/8snC+8QLP5qhNeDSfS
8Qo1ZNs8YL7aHSi9/kZ3GR/dzXGz4F+tV53F2m5Mitl6N/Hhm70vREK2ezA9INh8
ZbGRmpQtHO6yDKXSwJ3++wSXFHcq1MnuQeq+RlLGgxZMzysXVhjQfo7KYqY8FEOm
GXXVgsZvBISGj5zMIdniblH/WINxzgua8Ezn+GkgHeGDi31wi6ZJBPGKUalUpili
kmKc4d4+quLknVshHx4tuq6D1s6L9W6HU90fIdEFdkDeMd+slOG1UQoqlUW+la4X
tPkhg93tuvZ9NHvNoiZV1VXJD98IIa32rU0O/+/KDmqUGzjQeIJ83x0+j59cqKvS
jOUX6Bh9VsXxbHWHqCeP5/ky8xLQfoWtuDtwG3DOZHSwJdwG0tNG9POJIn0vH2YJ
uSV/ExxwbShs/fENvuLkPgG/zBpz0csK5hthndl/6UCtSi6fAeBLsGmYD7WoAJ1V
+yQp5pU04lc7Zxe5A7shGcoBB2Oxunk2ESvvkr9G4l0ADU4tmiVQH4bx3AyyPX2L
LytJp8YNttthqtHrLioc3VlxCfk5c0OQRU7IOW86D5chqssRaz4QuwgT+SKWnQp9
t00ClR6KvBwkONDzm9YF+iVpzLFcHxfLxI08P0K7ef9PNPK+2l255y9kHBNr559x
X0IK2x8mcTytoyfzLuhBc82SEkZNLcNEBOImqRmtYe18cPbCqYnNqtHhCtyF5rH9
kwX3DdGUhiSiSl61hNqgkbBJ0h6jo9ngkdMJG/IRf7OkkAHokXX6j0aHNDwKOena
72jh2aXGAicdxy97z2VQ5SXPaWm6hcinw8CEqLnhYybIaCHI6xWMJiT3woIMMSBf
FmHClnDvs5DsptW6XBtyWEa9PAKGKqz5NkPl4QrcD6PwAWAQlaXqaPJDnW3uSiFo
Aklmc23qfSCyx6wh+yFBTkdaGyDpXt/gPy79pBKDye/LEK0UEWd6TYVx9KCthCyx
umWZoATeXCC8gbNqADgM0FYgizjjpl9h7SwED+rPmW9WOsQVfZew3f3bEaxuE2AO
32rkLA+1U6XfHwFo/5sruJOWMJnyN7L6ZmFENQWFXCAAz/NnE46EWgfhU3pXi/BL
/Kwdvi7YYnzLeMFdk9xDjG5AAPmyNcJCHXE7HHTHSeutQyJftHmGQqAkls9NeMjA
The9zn+FSA1xhVSlEU4PcJEIiAkXZ3kxw1eDc2y1WFwNi1Y8Vfoghx4MtWHNIq3T
EppZZJJt+PVqmnGTNFN2UIDHtxKq0Y84VSsPBN5Jxkhv3sHBJpn9e4DJpTtYxl/c
fjBjfAuEPgyzpmGPpI5m3d1ewqDHjAnW4zzYnWNIW12YIo+0nOq05mo683ddap7P
r9PPPQCflWiyh8b/IOuQSe6RWIdbVyaoQJd5vZd07pTkQoz5dGyoO3cy4/DxOvXA
vkHH690wmvP7kEPRGcx+v+PefgKvaG0L4/QR3fvXPOqPqiUEVy99f69iLrqi1QSp
DBxzXW4wKnj+KsEtb6UWaOoIUN7lgfjEyFe7us9xxEAaxPP02zVb6dVKlp3Z7r1w
tMLHJAdedFwUorT/paaok8PluSFcCv13e17y1UAxTx4fBlpighICF3osiFU9acoM
57628ttGPI6vqEhgOt1EU6MgpLcOptMJw3d6LBIxF153jTytnLCTkUQIMUJfbWbG
RMDDUEQGHmDtRI6ZYK6c9NZlWvpx6xZVoL+jtwfwcxmoljQK3mU32wHwbz/7ja0R
LhLHwydT99HV8aYV23J3sGX3SPosyixHIcdVQK5g0Bo1Iy6XaXWlkCqblBtrPov9
6rMKfWecbzIRJ0MmzKCi9Xj6g/veEIqeR1MlWkY9Mabtw46qf3XpvybH0eQ5vPU9
ztCdeM/Za5X7JbD/ukuVwWiyYDITY0DwQQJ9DQ8g4sUcQBGg5ilKCwj8sGU6hhKo
Dm3H/4XEOSknN1Vrjn0KToONnMK6JmNYAUxIP6+FS7MA6Z+ulNm8s03vqH3aJmDw
qIoDkt8Hj6M876QeOOB9RmeOGn1RtBt2yIm3BuoaKwDGJwvU8woL78ioVVAgyaZa
hD9Wi4l0R7EhgqjDgDbG6RgBe+5qU/a/XA+a2jKV2fxLjnSGsn2idf0aDV6DC43a
397Gdxgs+v5nwkadSouaFMvplpAD+dZNHM1Fbhr7xi9N3kG1Vioxndh9blY8lHec
X9VTAh/aFvd+KcJMSCFng+TILBWalJriYqRp6gzsDA1BAGi/zWJKkwY0NeB3fdwa
g6vkw2IRFToQEnvzbzY+YV0GcWelhxolfUQbVLglH1JSmq84B4efFVfwKwMqKjQV
JiFNc7ycuJQOB0lX/pytvdkPQb32ULjRtd5sYP0V5pQg7oYJODvyAn6/TEZL3vbe
mCndfLc6QiiC2jq3VuBpcqSEbZmhKFfldrn3VpbL2rd4kkvhsILkaWnbkhfi8mtW
PhAge2xhfBlVAtWIAd7VJ9S6fH2nB0QxOgKpfS2TCOfj3aAQynDPgnMbgZljGhVa
hdeW9KR51QvpLkT4hQvHCot8kv5u6MOXKOJGTXt1S7+T0WGziBvR6iJ7ihu+ZBQK
ycPOW4SFvsqA2+lFFWTqANHInJ6SNHcNzbeTlQr9LNWZ48CWvJc3Yb18uvzMxwrz
0RCYz0aMrYAbge1U8bw6JTHodx+MhnlDdJIHwB34s+BwHhiq91JZp/U3Aa8ASo7M
d6sdPO8gfyz/3mDhdOKW5b/xZswOqwdgBkRGE5mNDHvKsTVrk82XCzgFrp9mNfYR
EqZCrW3kWMULYIGnnWXVOEpAwKJr4Mvnydu6levMOxCl63awu5jKlsWC9Os+5wPR
9kdQNsBzfhcPhoaaT5VkeKxrEh14tZGfWJYjViHBq3tFPiuoNyWVqmUaSCerE95/
4Waq9DYszULEh/Ul28hqjXEsbuzo0cd3ocP18H/fkY3AbsdVxcKG9tcd6BnkT9qE
2lOPLsQTFosdkXZUXDBk8PEvOyLzMPWQ1rvJcDj/9iQskP6lipwJ6v6nJ5bnH82P
yIzAYUPm4yC4wHeHgzrvA3D+066PPwaYhkmw7eJA+bCeQowds5esYjYlkS5cXt1y
OAtYtMIZtYiu7NDbC116qgv9h1JbNy5a2HB1CJD3DnmQq0sMhQpALxM1o9EsiIiU
28k9oNwZfZgu/ae8oB3v3Ss1dmLuH+b8MT2hFH+uQHLSzhjPMJB4zAx/TAA+e1PF
OoSqRmUVZCcBzRUMo2U7CdLj31Q96Js73X4fFyk76qETgmOmX4Z1PKJlbHDHVk1F
GDR5FJf7TRyZXOzK4+SqfAOV6BdOAw5QP5uPOk2pl8JzYlTcZvaXRU+nnvakfXeY
nRqmuxpxdLxSGIulzy0O9xS0xys0ScLKcb45/aJFWU3Wvfz8joe6Eo59Kh5IJhqT
BxDL71UlOmSMd2lsxQCxHnyKpEGoZN7+3oTa/a/CWuzySx/3K2rdsL1r8jJixBj+
buE2GeDSQpXj4DxXpRp2VXE55i8scdVgDH1uc2xXnZ7qNxOLTB0zHBvnxxFydGRe
bVzm4HmacwzXfUMDgCEfZbA180bzLPJq2pMs5Juj04RWbO6VZd8HO3gx+mMVAbyo
mT8QiYAUF2BqP5Tu+56SjWOZDmFnT9luJOoeTok9AKFjKQXtIyv8Lc30TTI69T/Q
IzHMDKQzLMXXDzptfBB5FEx+7AjKA+8LxoFWvAijEdxtd1v4RoSFq7HfDw61eVVI
EI7v8PsDubukqNcN0ycduTggccbmumNNv0/Q7+6l00plyy/Yy7afIe4n+J8qSzd8
djKx2fa7Wlpn34TU+CTZNooBfQHWKbn5SI42Yax9FbSXHwnMy9n0j1ESsi9WLV47
N2cUyygh/CQjW0LsfC4VYmKYrTW3wrUIE9OUxwNJRQFC7JD4D9OVPbwYTTcZteK/
L5TlbAGhJCUcr0Q4SoaThenetnrFwlzmyr6AnomtLR28PlIwhic9zdfMX32DH4eF
GaIrOkAfwxMdtZ/TEFE5aR4I5h9Q4VWKRykmJx/xLCDZF/q4S7txdloH/xbepUrz
L63+vTnIiyuaMnIvtu+fLgXowMKRCLwAX2DF6KsDBHBhxmWYDBoNb5qIdWq7Gd4Z
ZpGtPVciVZUZqXXdA2bmokJV7gz8Bwg3NNG3SqC4Lt5yiJlDg83YsLfkWWC0yGbB
qYzSZIHTz4oHcXM08t5j6jD9vpFAtGwwk2DH/zA6YHV7qfEtsmJerL0izdHRYrIJ
wrOPcdGVBc3hZcKkslOVGVnl8oUKhA7aZCS2lOuvlgOhH5QQqpjKOziCQudES9O1
EXcWDO0KulUl5zMeRJrp9Xmfyd/kCIZ0KN7cvQ5TzhdWWSpQGAKWYR4A6MG16bDz
pyYY5K8xlGYE4yu6aoTYyJ4+K7r1NPrbeloMSywL3G8Lnkv2lJAyTSRO6NjyLh24
ou9KyaKCbDGKIyX7fYHADyoKRk6ciAWzN7+GRG3zlBrPhl+70vEk8uvNoZKiKldT
UCJ4pschHBD66c6zBEkD8uOMa0LGit6SFhGPyXinZB4k8a6LCZOJNzj7BHiZOm4k
Mvl7Xvge7inOQIxwjDNZxuNEhZznNbAFmMrshlgAXT5uob8nDbteFf+0CFEKy+4M
sCQ1eMOlBB2JRmpZueyJ8REUT/OfpB+qiB7BTtd7CRhGqGpzm+kCosOEtQEQ7r1C
BKmOReEYHzktoz/j/022Wrx0ueMsHoQEtemiIgZ5L+rN5qFiWH9LyfY+5s3JKkuw
xSjvVbc3UHeWMfbehZP/QW2OmrFwJzSREUAfjc5LZ/oLFc+fpFsDiOUFCLeT+nDv
pvI3A+i5ozRpdt8rBgDbQ/yT+spGoYAlOWiVFVt0fU8J4+esUAC+Xrr9kVdDmnni
6XwclcsXkEW56YdFrBqJ3AABp0nB26WuvsrksXlNxZHEPq6ZtRBC2LQlXBrfYhg8
V4/KGG/tg/Sgpv6x5wf/nMueFuNZs2dLq6Oqxpk6NUBKagJtqwSDqXlcqHMeUnPN
/LO7ygR6SWa9R8gnIjNDwabGp7Z1d4YKysojvA6+1sxEBvSP6PDlBVAzziqqTlbI
hn+za3nAaeSLjIhB6sSlNT6uGsrLPaZjVaMDlqLF8gVvEyS1GzfwikdiJ4oDIwfC
Wi+JYldRWGmxpoKpDn83leisxW5wjkBdIJeg60CJSexos2RqlvjBjFKJ4wBl6loz
oriajCMc/I18z9lRM9OV1ZNdxwDv1F/lzKbV+ZpUzWU0R4b9dVLgk54C4EZdULeE
GAyGbk/3Ch9+BlZQCqFaHpv+CUbk4iTo/orWA40qZ/yEpTUnILgSXc9RS5mGQXUh
vHPgE/g11A0RTZw/loYjvNk9NljmdRIQ0Yy2mT8PQnV9Vb/UIT1PlwRSDV9+J9G1
iKHkIgLaHaOtXpcBY7CHiFRYOkIz+PvGOg0WUDvO3AS6TniHWE2Ne5k4JJI4R6zY
i1Psf3yp4OF1jt9l+3xtes6px7SkcQhZr0N6KTiWp5KX4fYC+q3GFq9630VQR2Em
PZZip3WHKGZuP6fRVtJwHJCEU0aM9P6vh2uTSYcnLYU8f3MXcy36OATER7O4ctGh
yEyhYkakCoJHvRjpqouRcFLJTg/8wvOQH5apbNNtzAlV8fBii922gcdr1amSqnWM
HZcznqju6GNGTCsLjnUIA8liNTULT9e8wpN6DzD36IX/noSHHSwjYM42Kcl5j+BN
wG7mbqu3poSavx7p7ABon3xNgt6N0ZNXxUS1ploPN3HFkQ8quLxVy3gdVdFrV/xD
YrgNZed+5yAdO+8gkG20UCHwdlZoc8AAJXI6hu4gLGV6r5sip+RtFoxe6KJvmzQA
nonHyLsHnz11T5potT5dZsDg8qqWmU2FyFzqUQUeML5YSSTRmQzbbjxzK0LPm3pz
uTw8Qws3KSTbid6hcC0rI6gQX1/0ZMuzmKDZ9C9Jjw5guKm+t+e11QOe03Sb27TV
bhG6vquzHbEJ5kA1EbarQNB2p2Z58RbMZ8/KL3yMvhYMu86+KaiZw/cCahzJZ2wE
otLh9Wcjr6mScir7I3SStgLzTCLiqXV+dugQDL/s00eIzKBobNeAlNBiTO5hC5xd
wJXVUw4+qsBfIjwFEfL0cn9fpNa1cIDl+6CQIEfoWs2HxAJmTGPbLIp2AZuX7xyY
qI6lDQ2b0ki90Sum4ZGZMdoMipbSrYuwhuB6KynGqB48V7QU5sz/CJkbAjadUHFO
AFygWNkhRiQ8kCYhiBCEqVwbBDztDlEXiZDzzZSnacc38VZZGI3srP6U1Xx28LOd
9Hvx82rOl34ZmebO7sYcHPHdZ6cfZNAxa/E+GelskoqZi4FAQQQcai9QUs5km/og
m+gdQzQil66NYqtrnMdXsjEosqsRkS/4mdKyRop2i/UF0yAaYsl47BWOwqypjVvX
H/ZwsRGWGD97VB/NSYLweYRfDh5pGpJ4HNTA5yaa8/UZVjugJ93bzLPWHflGcthx
dL8MHCwPOgYc+pWYZ+ny3l7LpybgbjLbcckS1PxYmsBAgJ+B4vX9fC+yUmabrW6N
JUZwxNGLTB6hJFLWrCRgdhgdYdszIVWnjd7Gadlj6P6vj0Jr6RYW4YhflWaKWauW
O+TzQ6HyvckaTkBM3OfxJWDH79XlWUcJI+01h1b/43WmPssciIemjyJ8g4+bmhky
p7bN5i/5pZpUeUPcYFxBsQ15OpZ0KHfshMNxoLFZyk0JU50OEuCU3OOu66U47gWA
4JU8o4zhXc7LM9q0v0B76IAmYklfjkmb0sI5hjGnuc+QiHlZJbWgToZMVMckbHu/
RyO3BZn5z17R58GEJz2CV2a7wFym9/6QSdVUzx35vCyagnEuONaCwXzmS7zA66M4
eaKcmXoU4P5hPROhRh450YWhzjauNR5QAM5zgssZAp375LgpdZ6k4l+9boitfBHk
mjz3LTy5dBVFoK+mWZnluKzUvItm6UMv3GBxA6LrJXTXDC/A7K6VjCXmLrclyvgp
NfwVB7KiDS6fMdpcYv1U3/l6904+ZWAYVo9Um//bn4/7Y7Ru9mMy2+KkZCqLEM9P
gg8xkEPDAu6KzntVSRETbhkYITvCK2LoilZOKEnItd358QFYxRtahVknk36RCxg6
4VffouDHcs/eLzx4K4016OxX1G4kRRPuv5VIwglXoGu5CyENi3E4LIuAmbLGYQlY
aWSNP1nkQI18MNai1ij1uDqGqVCBi/vombxYgl3ojv6BrFCvK+X+MYXYQDP5OXQc
+OdUFaWonXHosg+KIsRtokT3L3iAuBW3xA6r1+bg5+vAef3nEVQ+aao37rExt0q5
fyE9Fich1XBF5UQPQR2Sjwh+7xzs/qDN+N0ImP72ur3myvRnoO32EbYXhVwb1P2Q
OCtWiWqIY7zKaDRdH1Qtwsp7SxJ6lR9r1kwmLbLd5+1xAsplDSsNQRb/5NCP+EHw
tD06qJtferDoPNVJNg03DHTJYwLS/gd0DVvCIxaKg9QUHy2zXVHH9CrUtcPiL3Xk
Y17FDe+rPGe2Se52beYGFxdSfM66jwU2dEh2MBsBBwpll5UAzc0tdrvt7B/u8ifr
k4h/YNSjtV997GyI4BFYKgpOLzLZHN4bR/xXP9AKE1QEX3gyoaL7opc9S2j1Nhrm
eXuwxbOce+74VsQZ5O2pwWxW097eTnTdQV9LQc9g4znplFmaphldeVMIFLpnbTou
SpqT/e86mgkiZaXQstO7fj8wqSerRScK9JE0wb3dF4zQyyuxgBhQKlN828sgw/93
ZbO/mFkwN5UxM6ehqb6DxYV424Gjvkhr0xZtvIvjNGqHLiMaKcgQql/+b1HhVrTk
qGZy4L0Y2Wuav3d4UZH+wdhIFXNT6d5jIlcCBC3gPsDsn8dyUt2v2zQbBGK2I+u1
egkpEX+RH7HAZ3FuBoaajkvpidLUaJpxEFvwDskhWCh5/b8dTNagFDhFZuwnR8d3
yPNg7wqLArJCrKp2/8zKaJYlxAA1cEQnYZ3x6b1H8y5bzQ4J3xsnlewSijK4tQP+
5zKPAX7/QwWKaVjWLcG4IrKHALX3n4nkXpdf9AC/y2tTOP77uOe/LNJW0BqhxvMO
lmqdENk3fYjs9hCsMAVWv7n5nfqy1hOZ0SZluq+BTYervRz2Q44y8KZE/KlRWf40
jmm4zSVgM3j07q9D7MJdjuGSqoPQvXt/fpQ5ZDJd2vrrvsp5oHg0+QCPaRrMvHLn
bmgl8l2P8HTKRPavK18vbuCObOOJIvPST6jC9LYlexNRcJBDCEZwfxEVkaYyLUAB
atKpCsDrooFOv6EDVSqEg0/o68ezN3VOlaJMI/82VQXHTbUvInAXjYmGnb3yj9YL
1w2uVtHgG1N+t08ZQhV/JIcimxUk6KxVqVN63F5bJdjMroMevehc5xu3aawW1s6z
0GO+/8nSqYeVSxACjxjSDUbCbYIxk6eSUf9wMX4k9CP9ozxdjiOfLN5woc+Xfugy
XpM1zyXgS+pqOQC20XzDOzwL4vuwXOdVYOBB5mnn16dxOlkWBGyGV7thom7flLzM
707jMIjHSFiDTpwUeKHvBlmUlYMfRXIuTp2k02z837GeDwTv15Dx8c8hcgmq8pE6
Ffrp0PkIseF0M99zhx8H4vepDKkwuA52MP1PH9/cVZt4gqcJXisEBJd3dKkqAYvz
sDOMEGOwb/GBMG1Mg5Qw+0bBFwlGovQ5Ihvec+K6DfYMGxsZJVdgVoJzvmdxbBsn
b+wAonL3iDf1qUpEFXTpd4+rSVHIXeC/9dd6LdeKp2itjedXcQriWErf15JtOosX
skIdwjGBbEvSqGtdMFsC/j2lK9iMZFb+E4BljxZ9zbaIIlowHt3d2jfreCrLZ0FB
dJW8e4YpWsZDi/hLmbep8uEpjl0Cg6rJL8GepJQmyhahYXvW86prF5+69fVUgB2P
FqTKtZ/RSE0ccK5PcQYv3MqXaL0hszwNsihBD79aorAq7wt/ucMOugvQCwaj0+hU
RkpRB2P8d0Ux3mah8NrCj0kYvdMWc6dM0xT38tDaFLy4rlKbDl1x+4lZM/X0UOzy
C6SKMlyngonqYOQL3ap1V+b1sFeBwyd2gPg+8NuZ+22Ry4Pa5ccKzgQIFZSB7Mro
8FatFN+2+/vt9VVrr1xuiNBqolT/m54n/QKBUxTRoCFmgxo928K/ILt0O+KW6XzX
UrAPUQhnyJ86XHpQUth/So8uuv/iETb7v+ok8tysp2+6AjOjDrxLaKfL3MWXy9nj
PXvi8nuHeqIJWmOi6IclSI7X3MJosBMzgmq0g6VGDEZWO4E/j78WRg+XUCieGk1s
s/+kHNdrFcNkP1XFfP658oVX1nKE2U/qhVpg3AtBuQt9YBhnmIL7kZg8904voZXJ
9O/7z3xwT2tTlfyfuknW5sbgNAdZJFOzSMFNt65wCW9r4YG/s4zcFGaRKe+YTWum
rnSUQotNzdbkNh8JdPbjCT7BGN0+vN6uEbkM0NNDV8EdPxl/u82aU4g2aBmImUdH
SZMyFLEHrFUUAovoVG5LcrC8gsu4PB9CNZw03/TVd5WQZhij9TT7v1HO9W8HA8eZ
m6dvrPoeO3s0iUWCboVFSBcK27Ygi1YgPKLCnK0OOxsij/Oaj587hRwyiCvMTgW8
zYgj4GcZDLV5mATgEiy3tH7IEUwZNgjSJFmG7hrGP8h/W75fPSXtwABuKyv7oDJy
KjQI5CMZDzoKbqCmPprtbRZfl0BOO2jsTtLOnxKinoD1XnZathQvXglNu10yLrbs
fkLjplSvydZMnXZUmeuIFLPWDX7y+vz3GoML5XYouigyN6MG6pkissiCJQNEaOoG
0+6CoGm5WJOOUVa9CNNTLjTYUsnkSey367yRyrWNB2SvpzjfmsR1JbfB0e2QIdRV
N9e/uJ418LQ72pjWKHlBFfQxww3aV1Cc+UixaxMb3uXwk9WullQpshMW1VBXlk1a
w8IN0SfPNtjN+JrhNQSO4476S99PzJEffo8sEO5NXM7XDt3F0EE9qK10bOj0WSTz
HMn0QatN/bBykt/5ptiKtmgRt+v1v6iICk/UblgVKr1fMi0AHPnfcgssKBkMlNMc
+54hIVZhttEJ+l0rZaJjN5QY7YSe083JIwIR9eXL+koa/yS1wdH/3+UOw0Rc296q
8IhG0YbPKTGLcYVTOnOv5TQRMmGVxdk2KICKPQW13OuPGkSPnqgKUsN5mlxvheVq
chtJoG7qdssCg8uB7EfHcDnfSg9K71dUQizJJnMDA5Nq/Bn0htBuQ5PxlExzN5bd
r8rshTlqvS90us4917HD0eXRGAkPkJ2PHoOlcOkUhKrldBSLuv0c6SpGPSLrxtsM
3TpWGXkOHZ4M5LvHYXtZVy3EKsuk5pW4PfsZ+wPAAbIDXiasb8UobNzk4LCn/kys
3UcQ1W5FTKhfHnHLVpTu0ULaCer6DgwP43S+KlAcVkqfiLdvdJ3BZYIhOa3VRNlv
zvRzC8AXHklF70hlMwLZo8xzVGlKB1BBQBTwq/yswsDEjcpeNxjzMMvPgyza6fYM
DE4o0cptDoLfFf6FApjNqQpTIfh3ZgFx9LTD+JwrXleIcLT8MLqLFepmNboGvAyr
hrkOhNe2PilHjTrgq6TsrIG2PQhg6CoWCedZTOjB0KjQmoe39n8GnhsIc5AlOPOs
MzLdTMk8aMap7e2UBMVyRbH7AUfue/fWwgyELxdpj2Tx6SIgoaCMt/Xcbn4KR55j
j9tNYtThEpWgUuESUf3ArmESuHTjJdcmb1Rc+BWtsulEH78g1vqkTrmAOtTpgvVW
lf6LQcPP7SRrtahSxO98lFLBq6eF40VZozpGvn910uCWqG9xsjxTmRyRfC0R+P1i
iPeujMAPI31tgF6pjaJ8L7A0OSp7XxOQZvRsHgcrHatKrQelfMYd34kon6VHmTP+
hwOx4EYDq24l4/+zHDpqCjH9jyOvpeLka9XRzSw8GVgpegKKRfdaUIaCNZtvtyf4
iiXKVNOttD3M00IJnmNHfBn+OXAr7+zh/3vtJj0tyk8oxkBALlzu278iNta86OGd
YkWhkuN0nWwnBjhRw6KDKYrpiXwRmEJ8pAUFX2MZw50mIirYw6W5kL+5kjEdy7C7
g1XbS5qsqDPSr4RD7KENVX4l7Jvw4tIEiM0VZBN+lSUXgbLyQKsHB7VOvCTodZxo
6dl6yO7vAkndR56KTEstViJglUmRbHXeQzhaGzDZTi9rkHNrtNaEuF1y2vAtrFDB
h27IybongoIJzFJEoRoIp7BXgas3SXPaRQXQfb6f7VVzSF1QRS2VvVTfAronMiY2
5x2Sl/TmyHXXODSTxsqI2Wpfq4coKpsXqXJKktuVukDLzI45vy5+1AkER5NeM605
RzNpWHaWnHxIa4xU3Fk1U1tYseTVpqF3WlOYfFqFYUYT3UG+2O0iffWAG59PWvKT
6rAczCyWgf5H9tJ3LT+ggDFRyFo86XKYxci5XQT8VeGhEVlHjALgi/RkQ7kESL47
ZeoJmKh1TNyyG+R2qsh6gvBcttEvKAmL1qHX1x8Fp2xt6nb7ehvQkXpoFETqLJsj
zUZOsFS7qspCPWUDAfWmBQ57eMwRU1gYhKn8t6CtT8EAPEfhmIhO0oRWBP9rIgnu
GbtAh1A50oh9OoM1xW2+Lk+4CVTaHEKwoaETqWfD8bi0gdIq9ao45a6JjALiynOk
QptZTrYcMdHAmucrRg0qzwQm4HKY1gsGmADrTBHMcDPt8Ja+/kCYgJDZfw9CyMu0
EhPXEBGfSjNAbDa0uTxBX8N8prvYRW4Wc/Uovat1MhB1yJKB6p8cSy7/mF3eJDBM
KgcJvFVWMFEXrFx8DfsL2vx5X6VWRrYRzXF8UtKMvb8vBaB6AskICXjVMukp0WKF
hLrOvAgsLHR7XHst7Lq5gBGMPr5oyhzeGdJLjb0UInQF2GIJbwdcgjXj5XkQ3mNf
XUY1YwPSyVl1x5NdcmnUaE1CnzM9M5F/Grq9sRy44Ez2BfWgOzK801O4x8iTcaba
pJpmtsYiUB0ur4z5xrXfU/X8fukvlPd77rRsxHYq0H2HsSIYuLp3aqDAmFn6w1Yz
e3O1Bi/rqSq8cVnPaRLOgwpe//kw+M5j9QMChZtWOYoN/r6mdD4Gx/qd2BVPpIHZ
GKQY2uqXbUkBUvOIaSLktjBCTZQAzXRoHhNxj27H+tXt/b+0fHkbxTMbjeRYnU7s
ZD8w4ksMBABAav9Zv/j52USVcfyAjnUAezI/6qPiHWxP/upNe5Jsozq+NTarruDa
ntNv7SGMCR+En7MYyOlczz8DMDwIXPhG4YPntA0XrzfA2fv2ei3nHvjHvG9wYddm
uQmDExRqWKQCJeyLr7YOdBYo2pz7HFncEFibopjvG6C4exYBZVTN9k9FQU7jasrI
vNQQ8pRv0KHcs9CJMX31j6AB1FYQOr9elZifcWoatbaIK/AWZxt7Ud2qLjwP+TEM
YrFAwxhK/F1w1lFIltUJIk1r3KqRzfOEHekYTjYmVDacb7KYvsl0Q5rWjLZIe3c1
aGxQGJEGs2BvX9SXTh8k6V8h4Age5npNkg5KlPcUgCQ9hoKo6GqQO25M9YoGxCnV
T0aViugKZzgPNO4eXTWG64Ff6+fCdAutO3rB6C1zjxwbDQN5495Q12EzEuJ5CZFf
13KMZ8/HVzmVxMpqQn2foEsArHtUhhiFMzuUw037ZfIVMD5qLe1VG37hKj4osv/H
ESuzxjPZRy/5h8svuIodpIy3Vqy+FO2ib7z7nfL3sTGwgZgZYlBe7o8PH36UqyRM
Q4hA5xNa0MNnXCrDfQVbOOXulOW9Dd+81AnoLNc+2UxMGt3QxkSP6pxQzTTfbQnN
v+CUVbu/J8lEv55tWMH5TG1ap+JTdO8oNmYUrXa7Ivxnn3C9rvEsOb4xjTwsrH6R
7VWpasKvU6JGXTJaiuuZT72jmcPhg8p/9ralV5EMWfhyMaCfTFvMc/wJL8M8lI1L
rQhEBoWuWQxSeXQDxpdTq0AAfF9rcXwqqPzvvCaAXDRDuNuPToaIFTeEDHqxZFFn
lyRYVvtR8v3cRhmWuSCJQNmm0tnOSy21YPz4qgJE8t0EqlI9Fi/eQc7n12Dnv1Zl
ST9fRMBdnO3XcMRntIjCgkiTbiMKR9eg3JlwbrkNq6JDGJTtupopyeAAsJlnQ/pr
3OzpzfFi6kIihohSQ2vXLuC9S6OKJY8Bx2iEekeEWrSS18KnSZeVPpbyvXLsjuk9
M36YMBbu2F9Bo7Hjf3KTDPLnerojCWWnA+RayKtXA6iNbv++9CYquT7EGDm5cXNf
UDy2xVmh13LxD0bTfsr45AXXXnDT7I82OpMy5lxnQz3ukYorA5HULUEhwtzGTQtE
aWyIK3HWMbZgGnwZRIjgy37nzIrd/0uvASVa7iD7RfiScHm+n27XWGUr6dLhttLf
UxVsEhYR31qMdedyzuktGgASatVZJUzfrA5RKiWz50OvRN9aUDzsztuOtOpE8xKJ
0abJW9J+fwsc5SlDTxl+2aYRp/yOwpAKOl8HOU+snGB0IRl2fMRbRgnDU0piR9Gi
8j6QWLG0FzTwwnFZoLH5q1iAjXz6yC3P0OZJfM8V2WQ06qG7Yux4J2lEkLyAgkaH
ulTIgaqTA/CA3GAwDi1zXsIdDuo9But2Yj8MYIWm2rXaKwH8nUHTGZ84HfWHnSFT
z/ybEyGuQ/E59HCVTfTcZDY3Vgp9XNB78R/lhcybg/Q3H3XkiEE/ueEKhD3RMscg
0R3D77OhktUI2rNdQhtCVAi+hL5D8C1EH2JycTcpyW9NmyWeJ1pM1nZUCJOpyOy2
DsILVVT+A/fUGmEY5/USk2IRVOdh2tOtgdfaQMzcCXY/3Kh/AroLf8G+Yugpbxuq
I7Af3l9zswbnIdzoQILaVNpUBiTTHDNsGTvVF2k3SYLVcYopIJya5dqw6ZQ0q1Sf
HBpeePkEG1AfyplD6CPkGNYb64l63jYRvD+j3XINgzCaZYbf7XiAKixduZ9U+qAo
ORS3kflonqStJ7RQiEZ/zs86KWvXLyldinL+xKwnTwI4qrXq+PaHEjIOA8OGZanv
W7ZMOe0yoCHnSBV9T3gFBFcZ/atWDPBsiBvipOcU4ZRMX3Y2jqzpLQHvTtSZ8uB/
+6eD7pMSEcbzOhVqyRcRnvzM/VTjPfX/Y52WrZLOTShtknOVcLF++KyNvmBvHm1n
D641FaHxLExr7wy8N3NzC7KuVnr9KbzrjyivthMhfGHZDAiJMXsQmXsfJr5qdBma
BXB+buOBzZEowIjKaval6cjAceDyflQiskA6bWEfEsJdsLED1nn2UaPw6GMTrX6r
EsX0mEIJUBxwlKHr1mQomv5AVV5If+ZiIIynqohzytuZ8fkJfRw/Pk02ZEOf4XwK
enQJQu0nIZRqN5qLuhUKcbTvG4UZXo909mqW76C93zTBZt8U5yPxpqW3WZfgiG6E
a7GYfkbfjalXz4qrMoRj/iYKWIp6Kqgtr/DOsvdApHv0fNnlo6rRhMuTqWWF6s5+
nISlHbODcATq+dvkX/PMwHAPVGKUZfHI5pzRMYfy+jI4BJ7MMsuqLDA1MXQMdU2g
10kp8SbjJGdd1kOOw3fN+Sn2Cpxpa1YwHrwgT0hknKHY+WDX2HQvqdpLUNa820CF
87GHt5RCtopGR9WjUBbiKwSdCCrsMEICfLp0YlAenA3rLluseulZbM+kdaEK28F6
q/ZEo3AjDAi+wo/Gk+92ZTOf6VihXcOAESsnpn6M4o7KD6xxpXj1l6s3vz8KbZbV
O5+fvoCZYsHMaQ7atAn6bIugDnv005AkXOiEGLPNbyHowZCum0U0fvrjatXUk6hf
p3vZlHn6lUEQUfdW0aRRy+iF4X/ljYHVADXidudkiP1TeUiyaA8hhYDijXZfK/c5
xe/ishof78z3OBtC671xnfyyH+qyluJHhRteXNxxKdEabwuOQZaYu88IRk1VGVIT
4nG2+2DTkdZwRf7GG0hMIpRNka6j9ktbQNEhPEUhBTusjooCaVO9cI0tdnngzG3L
z7Bv46xeBwq8gMnRx1+sifMNqOpf2d8N9ZVWv19ouildszpqEN4cX+gZ9IHemupj
QY5tmhVmtW69YC8ubcsSRPY2wXO/dre8h/hlp+4FBNhXOupmpewcBVr5Qu0B1EXD
Uyp4vrGqfY0AioGlw15wXsVo5nvL7UZEoJAIAYKySY+iRBV4fdhwYSkAjkgjnQzW
hZJtkyxQASXworyeWl6jgp6aQUZIrsk4FMGAC9WjI2ymXhH6yUrau/yUJ+xNRVQG
dDcNUYz949H/sohFNBW1E9MqWRzK5p5Aa/cEPa8C7e3QXw7LqFqTk7Qm8suwFKOq
CtJ2fx1Ye74AEDFTPLxsNIDBGP9Iu9W4LpRwMj85KHl/NhFGGbxyMIRvPQ5MmpXK
d3aQEFHi8Sde6lCMy2t/PMgsiYd6XSLP9Gwl4EHOf0ZhkWxXwHjJGVgZGrV8GYsq
3Zdks2GWW8dPSXX1WGby20jJlc4AErgi1A0o4gNMfcTVGAOZPDktmK7mZ0CFkopw
DNDGIzRRqFuhFgdJxwKnkeeziexHHhgqW9avcQ15L0adF+BcYeJfcaq9UGB7f9sh
7PqdEVvbSwNAZHG9BBpiwFXg2kh9rRi7G8B6T1pRVk9/1crtOz8JJD9YnJzWO+oY
RCGImWafI3KU1u00ZtD6xQcgpL5/UtAZOKM0PjcZANs3nZmkARCHDjH1XDcQFizJ
UjY20Dqlpv0hl+efOVAHQrrPR+S09lZBKJblhq9Pyam5tA6pXsobC8VgrRqKeh0O
n8y9F5lG+pNxB7tRxh+dBW0ZGQhDyhJ6/rkV6NSBqq9Id77PTVl4Xqsci8vMJcCj
qWlC9INsBmZypqhGZn9jTs4ZNTkhp4cm8zYfWy+snukJQ4rTA7DIZykyNrxsbZAG
P9zBRsML5eE8bqg20bpN5RHDAbH9pHr5oQqUZLYLXU8W+I4SGDxZeXGJAmhVF8m8
Gy8CMcbkgyVk1XPxtzYq/9nxqrdRP9TkuW5AC7pBjOQEj2D7kcU1yYrARQQtpiAZ
cyahA2F9bkHQ54i7kNRoh0C3OgaWw9udiga2hxEMl6oh6GWDkj4Q+2bcQefJ4iSy
Ux+gSAwtKpPM70ii5JPPFOkWbpjFsP7tIJbE0jXgYoJoOjo+JZq2WuIvkTPHlJJv
k3TjTfk6yrxdPY9c0yIYq3Oi2KoREortFvpXUIm1Ywp8FtgVNChZRhoQj2y1t2mk
KHh4SArFen9UVGYmf4H8bXvK7d9ktvXKwcR6LpfyH4hA+Fn2TSkG456ihbDv1+Sy
Dv8/wl6OSVq9yuDfnjfgG7ktrkvlCaPD7T+PQ179Wsbo21jipjcxiwrDF/M1zThX
gMCf/XQi8gz0pQZpYpLXA1iZgnADidT5wveluUh4oJf0DELlCUIDCKG/gp9w7bQa
oDpQD7cZ7Phe8fT9Od7HwitKQmv7mBLTaQTFEHyRRT+6knigApc4vdzQLdtQiquZ
imezmnCgyN22pIOeWtze7eD4QlboSsxSbT8OII0Q/CvPrxHOdRFCMOlQXjK8+aoO
/+w5K2LkXlYo4anYVKrBp57Rr1fjFmqvb+MllczqvLkz2lKgO333jyKRR36uahx9
IeaDgkidIenfZgmuR0iDeQbwenNEeTXsp9GJh5FSl/aWD200hGA8aWmLri4oov6b
5PozOYg5TIGc1Ev5FY5Yprp/D6tm5nCBZwfPUqr2zc1SvDeXjR8FnoUb6MMtZNXf
vlLuG3lpLxlrXVw5AGGOCpvkKD5kERhcxM8Im8tA2sKXubdVfbL8aKuef4lKxqiy
YiWKZ3JYYqsz/WiE2zRh+J7sXY7fHxK6cOw2XeYlRRibRbxWP9l8sQZiCKcaOvvx
9WQUjUCsH+9ALHoqZxgFN0Asv4k7uMW3XPh9DcN+XeMTCJpyfjKXXoJf98oZzEpD
3MRbTCz6ScUwifyaN1QOkYOfA9AUg7MfMH026nZdSDAO3fPqtzY3xLymBGvd0yRp
LWzgSjd0vHY2vBOyxOwWIBh0Yipsw3Ni9NBgfFCAiWslIgFYtkXfHEMKAxWtTHHL
Q5RVyaD1kbpo/vqUtH76jLJOR9cPDjb/rShpi4Mwo75nq57RQFLmcipFaaGJ0f6g
v/UMMK94rJPZpvMFZiU9HgSM+jsM3XoHO5Y8kpHwQVTpo6eNE7py5l3UbrrBckkt
pZs1MD0yRChslg03QPGx5cUKcqLCPtsgzppyXQSBdzITIHmr1HnS2v4TPGL0BMds
pg26gmtBnjG8setDDEzFfgy3Cu8mfn4vk2yWgoVTIIJNbNivd44q4CZsaOOnb5JX
fjFRkJfGYR1XIAf9tosej/6p9DprjTtMOzZuUv5kKrrmRbaJSa7sB7kKGyfRUzar
IgXnciFa0VmfyaW8zftpXpnt6w9VpM4d9E/YOHd7BitEWu+GE/hCugB8BubBhGNP
/EODsaaIelj9IYvX27GQn2csar9DWSZy1GkeXvXGb9QnhFwBcCotFs2biKwTjkti
6D9kY/uXvMQJ+qhKc5sc7XQ7Pc/kDPMnmDTSEF7P/HoO/s2xY3Xq7yF3ge0QTt28
1/b4rmiNq1qO5FEGjS0ZrWu8ePVSufIAlkwhc7uoAeS658JEx6LPM0CqbhJ++Onk
76OBW+kinwzdPftEO4GR+TLMxv6vQZSXd9/ajOUFZJ+p59/caKB6UNs+mZzBb2L2
/7T/PzpXiG+MZzhDuOm/R6S+LA8sM9ziZpLItp6M3ULoR+bRkNZhQDPD077ox9ya
aUNDUV7U+eIbWRwh+DliQdZlEfobKgZbdb11NoPDMHMHSQthPjulptdkeYnOc2yk
C114D/0YFt5xwaWVLqOUWR7JJdcxOx1p8bNl9AtLU+G5A9hToGwcjjV7CkPVyYkx
Bt5dIgrOnwunK2dg1R0hV5n1OWoZpPwn7QEDROc5PS5es2c0agR+UtxWyXuTnas7
lLEzBhB5MjdYtfXIZTgj78lJLDm0Xs5QVj0ujwH9X1X+vLC/QqaVJlUJXLhk+50u
E5UqaqbXLyp40HIPDErVRY9ae/2Pz1N/VfgOmGkdDBRuWCcRQE1h1M8QLyDpuB2A
GXYH3uyF04C4TDp0QkGWwOXCysFnohtp/IZRwZ59uW3HoMVhYIPu25Uhdnhltsp4
XsIx8mVUvFnroaGE/1KXR8H11R23v8A8CX8GDAAdezXiO+YHMD6jvIt1OC+2U7s2
8cbrguRSF/4/lMJIqIK9LXFafKTwjuxR7lqaOVcDnwHPhQJSNi3EE2bgilhwMs0G
s9FBHksqSWRE35YmwwGKUST6bhQ4EOHtkU22HXppvec4h1rIBOTkYb7/kPAyKGng
tpqkyKpOsJxvyQZn5o+sidyn49sS6vyFUen6yQ2KlJlHBh8u8x/RJhyVNf94knsy
nade0zdvYHoYN9NOcOASkskp7eo1M3EDEXCovUjF64CWheClLZsKVk8pDaYvKYNM
Eb7hgp+53oOY2p9q7OU1bHpGkHrWt0NX9BJNmELrKh29wpSb8iJAMrQI0uTSIpvf
GB63BNYZ0RnDEIYyzF32TNgD2cMeS8ZGrhPMEgcHXoZHkXVCv7fXIjKDDTv9plAf
WMp9z68UMjW56XYl560MeHXdEjfhSPk9yQhDms6uHhPyxKxvnvFODCUzyl5rfQEs
mYEPXPxaue2DY7v3j+Js87JkFEkilO/by2XcR9JaTlpkyuTeamStqEAYn+tlYK0L
2sz8L83JEl0a3oiAXiN+e1nOiQEfjBqd65DbOPs/qdVpJqkDbBuH3Z0orRaAk7f4
CopF1TWTa+lFBdJSlBL80UENkDW6bh13T8S6e9R2JHyznVyiv/5znD5UI9wTs/I2
W+6wB55TJYMaqzqOWf2AR5I5ezCdvK5JRDcTrHCn/89OxbP3GtYBYTbhoQQALief
vjuNgVo/ZtvaYdAqquzX57AhGkFfZieTZKIm7mPRx1ovh3Dlbgk5WNx9KBrh086i
L1/irVUQSrANBcvCuiTT/A2jurbSwDaNFq5Vqc6MJt+rsgfeko5wr5qvje4pQ+EV
ostwnmAemzhU4P+146Pego48acCqSg3203EkVZUL62YoCmZW4zQ54P7QTSq+xbGz
xOOYwCv9n/ZVndhLFTd8gmRYrDgm72uUFHvL0pGtkVSqGr90Qd88s+YKjQFNJa8i
s5++cFq2hDcGGcumOVjVpj+qSe/3b3nQo2rdUaKcmeWG3VljThoYiNOZ0V7wL8Ct
2ATjIm1cTrnisjDIJyZUwY1d7/hB6G0/Kr712vPKKIlvRQ87Fq5iHIH9PQYAo58g
lk8n5WaI6F0UsDYTEYZf/6cnunbwuMXYGj/Tp8H8fhqaY0d1pzY3tFfYyk8pL/GP
aH2EYXz5x/A6lHLw9sUr1Y76p5ov/ZSeSGpG0EMx/lp/Nw1xDv+GsgqaT59/RchE
ZMXoVELpZR1nZbR6Dqm+kkjKDUi2zdZ1l8vjPW1EKU3P10CGtwYBvfravNVnQfdQ
ZiQ2T4qpmRRECvdkmaYMNOqkL6QF5qcTRWf2bH2Chzj33lOdF/hnWW6887yCCww8
vR5HcOnTuzyd62mnS9oZeNAYe6xfCRRLK7dUJPXdkMZQ0AEWVYaryZE6GU8B4PwM
Hu8X3Lis9W38tD327WQlTR3VJjuJVHhZ6Y70DzG4kNX47LS4EjpUHYXFZComPZPs
6W7HdbkhcD1BgCYyfsVFNcn5BS8Ih6okeSXG0NLLALKLGE5qmUYrRjzaTpmNqizk
UBOSaLENsScg7zo86jgJuGPzf9vz8wc1Fstl20xgDyDDhY+UQZqOuEo2votfGJwI
PDY1VG08kDr6WUpjeCWRp9n7AifD6Z/GnX8LqftBqcCntr47SHklbk6h1CoAuVvP
O0h4+6GsV92zBbQ4MYjnDfgA1t5eJr0jrli3V/t9R0Ubj/y0QW0IgEazSaa4tF7P
Fvf3I5PQSN8+HdWWo9XoJtoUuvWjOIXmiDydEJ5P3euYjzFBDXjBeOQGOIBQuLpK
wTyIJmeA11RdhoDvXwL8DyEYHoPC5/gBn/Bo4TBj5uM/sIVh9P2U1jsRGgnWeChI
GZAx0y6XKzNgs+Pk1RtEJFw+mXYswBWq//U0B+eqYsZTC2vGiQoZyOJV5hdSLy1D
JOzKeT9+SxXXV6R4F/B7txyXv6So+LHM4D4ib1rRv+ABX72XDGTpoMfjhf5Es3Gq
+KXo1lu6Ivbos9ZqDtfnsS8IceB0heqVO5B8RWxG1ZACGGkx7Esp5mxRHz/gllUg
yQ+qmi7/6OLDyai1aABR/BrGxiGZ6K+dERkQYQvmX3wx/esr5ANv1wcggX/APo9y
dz0vdej97qo8tnm1JONxnStb5Zgx4q0jLWM83aHYD7BYHYBOWocSxONQJt9Fuyv9
9Ou47FA0Im/QdJdeG7aE23bgz8A2p4XdW8lgaU7ukqct87/A6Ri/csPqDzMiiRCk
MVITZxQeh+xrCZmUvtbR6be33Uu46KSrDa27jCz/Ilq+JmdykUoqJ6fLT50cOW/C
0+LRFaqgEycoL0GPBXI5SOjza2+fsg+tyvTlUHlp6Ku0iLb6B7OFQHcd51keDh1/
1lpq1Z7j/L2DaILSIjZOnUCfaIkPwTtJQob0+jujGj76PJOyIE/Odth8EMF7i/od
QbfnnJifSozFQLbknW/rSG2HuC8I+Rc+3/AaNV3gIfrWJxPCkl4pajonFKkGV64+
iTg/tEYXiMzoZg3e1cSBnozFv/KOCjHZva4+Pav99k8GZ2XmJxSju31MFmnoL3JA
fubI3Lvx3jYssGberSM8/jebs43Aeao5td8BKUWi5aYmlBAZ1rEJPwB1tGkD4b3/
+UhXg/s71phTig+aOC+JbL3F3praRFx1a3STqM5fHdXgDNfZA9y0GH9ChUbaaW7L
3NQ629UkEDDHHOgtDb2YPzAZ+Bt+MwSRs57eG4TaGIxbVSpgroNezP9Ed4gQyYz5
j/JQbh3gVTg50DrdWXECgdiZzz2dYvV6rQoCB7raT9yZNHJIGIUNyD28OQ1Z11gg
DT9tp/hu9+AsFqeRDMeAY1i3+SpAbfVcOKsKWuypCKwEeSwoV4IMySUbV9vFjoTJ
PRoPhzAaNfMqXc+tp/I4WqTrOPtyxSmlc1lx1Zl1gk64Ngi+7P2DRNCHEolQANSB
iJJUGTlptMYMhgj/sv+sNx+SgyDVd7zivhfqo6AIoivdKMISuV1nLQNSOOOXaubS
kCdBnfWDhpUHDqEGqrogCQMcPTR2TsQm59XQ2gay7tdMHq1S6MR1eWzjAW+60U7O
OTzeUuVtrT+2xJUR0UUKpJNOmIAY4uapkzWkU4gJdicrSRwU0jyCjb1F8RgtGKXf
qFOUKk0TrMiXw7Q7yrlx03LdCRZKXG6i/P0JbN5aSe67SCKtkTeAYEtdQDM3jKTU
m0rv/3MoEx609xwYez8h1yw7ZyJHQlOIGc2NsmNzSeTFasgtQrTYZdUlU4JIwPkW
hg/hxrt/A8l2xZUtqr6ibArO5rzJVlILTF6erGSEFSxckBLihW5M4fQMoBwDK8at
rJkW5vVxqOsaOzSmpQv9izWuCqo3x7prfWS14yjRsNBMayjozhmrd5pUwjKz1koH
mvFjdmdcLwy4mB/Ynd61SvWJWXFn8Zh7/H0uJ46L8AgtR5lScd2gYrq8lccZsq87
qIUOPaBV/svoOrjdWrRupXh7+nsz+bWZlkmBvq+UqI9Gza0MQ80LQ8Aa3fhoZnof
L4hgY8JMJh0DrmuSotJyqI4P3bGPZzuucthjdxmJDLPeTFtdxJopgOn9iybCu5+2
ZdOhG7s4N7Fo5fsTCO/1knmBIhCDTRqVwobfAvIkCnCxvWqyjVj+hU4Cra9TqMVI
QEF341v6Qv9KAqgWQEfvElavhTZkkYUlvCfwi2FkklgDRc8KT0rhAwyrJKv25ErX
jqykJrwQJ5/nV61d0NiX5tbF6uDJCW9NvvPl+66cYJx2R9pGVSzfpln3yDXnn1ng
j/mYstuubzxVMcud90EfHc7PS1qqnFoQp6+DS6smmqaXXeC2H4Wfpzo1GN6aK+ev
OyyTQ3hwuzJySwVjWALeyprjoMytQYA48nroEHioj9XslA6CLcw6qYntPjJFtYiV
4EACYK5z12UYWOQg1AESv+i4c163jRkgA0/v/uxarxt25Shvb/tK6ZGM6RDWNoA8
xe6U5yhurehOqCaUXTXsrFp5bwGAxspmyY6yxaN4yk4tKY4/lhQC0Iqt02OtiS7N
rZXAVM8aE01GNaH78CPMGx1RuGp2QUIsXPu4GWG6DKAK0mGGJQI5wSAIx4Twuu+d
4O9dhqRwDW6yVxOxHU5hMfvNuEEeu9aVNmZGTvZ6pADgeWv/R2DI9vjHybqfpdv4
hj7kePE6/AZ5fMcDnufWmQcYE9GPqU+UJN/PREi1O7hbihKsqBoIZ4+P+9ZzH1in
p2QWTQJS3Y5gsHlz3/zFNIy478e9M+CE1JhL8x/oU+DDXr3/VazD20/tyOJg6z3n
Xf3ReRH0cuedcL2SQIt4GzOrJZVRCf22VO+FpMVbAJ5Jli0x6OESRp8UL6ka3ncI
kHaTrUDbcJrxGYUUa9pD8+5uEoccQx7StCA3wnibNd2GnLKEa201QaUJ19C2fkBc
35yC4teXPEBmDkCiS4xzcJm3OuW3w/0bNWF1BJB6cm8e7JStwxm1tTdnxq2uhAW3
jIUiwqDM8IARlfx/4eBOmKfCs/60p27sOVzFpgorANGuXHrk+lRPOmSnXaQVNv3a
Klfpz7RLdX2YO/rKmlI6pSHLxQEwrObKTvP5cxzkKmfKQPNLSJtvULSnoMYfiQUg
QQd2z1sRMKn6RVVzYgNbKp2YICxcEJO2WxTydNVhOx+v1guWjI781NOP8wt4MUxC
NsuVx7DK+8AqJbdlAujsZs4eTkCLezJmFSmJMDvh28E/2p7GECHqfD9KQUGzPAYs
+72zBDxieQV4fUMd9c4B6AKjY/b4BE7xsOde9HGnqAyhNwGdDi0vS8yjCqAK0FTX
R4STAFPTZNu8yedMadDH/aSsV32sh4+LG40XIYoJxHGmqrVetCWHmhiiGGXuEkBT
R8fgVMuHKQSmKCmNTJV790tfiP/goFdAWMd3vVFn8hcJm6h70InCl7xQWmEeF3qA
Yf1K8DnhPgnaTnm5qHvNtQBapUHBebaR58vumk3GEQaa5zVNrFhrMX6ey/FeTr9H
UcpZ0SdoWvvZK9mEuH6e3hzelEHtYTTzJlfTDxk7bA9NEMPICv7YYj+YIQmEs9Bw
rob13Q77hywmv+NZsR60MJU1yTn+FXVUMWhPjy5q4LlFPJ363fkCXOMAimV1Yhse
7c1RdYFyBzAi+RhMZl8t7YeXDU5N7JD5ff0xcFRJqAu+C6a8S22nF5bIgtd/MlFz
ZyqJ99nZAEKVSfuVNMczLr5H2p8MIj1+e1TiyZjwgPuu5BNZHbtH0hUcdRKisxmw
GgSMZgz9g5trD4sKmyRrtCEzTK9kauGlWWtVQ0SW5IGbLkqTEoRm3qZaplMwmXM+
fY6o4gSgpeeMoToNv3xE631DZxqoJ9sPfYZH+44t/kESn2zgqBnPZaesddwyKTcC
fVHMjusG4y4+V3AEUlLOkOUekCgmF6UVLL+oT6oti6TPOTIg1a0IQkrhSzisFeDA
+IzBZWrboDc50Jcv8WpjZieTwMh8OHThxrTPJpMi8YNTd/BGaMEQsQ3vS17upt/R
K1lbEBGXeDKKv96TimRTN7VgWwjdlqkT/EkCQj6Sm+CriOt+mR1AEMfiLBHJNdta
ANTCIuSpRlVbh4iU8LTq9OUFOsNaH9BgiTQUlcM13o0kzIs0tGR36wdHlxwE4zzl
rHLK4+o80legB14oJgAzb9JtKDJul3REyZSCt0e4b0YYwy+jrR7SA8h7IkcW6kxV
Q/Jnx4qzIViwSfPKVbTNkwZZdnk5Rl83qnp6OQtxJjmpMLIzdy983FLiGzrY0TKl
R2zb7XxjuAH4HDVTUIhQe/IpeF5xlUq8MDPLnXHSrR/QFuxlDdpE9jKpR/sQjYiT
YorMLY6G4fwxaAuUQvAbRoRqLmWGdafBmnaUemhbdO1U+mTnaNyUYNbp00ebPWSE
ttwD1kFYJo4R0cbmjmeR9BmSc2ovLLR1n3uJ/Gj4ouQf02P4LCoaiQD5gmhjm6K1
vscRe/PdzD3Ye9fFqLQL22zkODWvcKpC1LDYk8WHCl06y3Ky6XNsIpISM7/wXy2Y
eEliP87fN0BeUvIPDhG87b/fJHfcJ2eGrsEOlJeib7tgMHpZRSGRSUAgQ43Lh4Er
u2zt9b5toBPbgnTD9rbe/wDaA7NkdrMi5paz5ZArQlRcUriMgWRiYtM02Oxm5ZNh
xzFwts3BIz6EgM78to6sVCxq0ZFZJ23Mk2gERAigvOdjXjRJyicBMf7+m7tHpib9
uBrrerZkvB9OHppPf6QTH3O2jUTehJ4HCclr7sWn7h5GF1whJkDxwchO/o66Z8Ip
x02dkVlZidz9RDRmegX7KQoUJkJZU3Kf8+01YXnVkhLadMFfuN1HhhF4h8/7rYEq
vlxlbpL6unJ3NWU0A7b0xD5GfYQd/z/iMSAXKUma9KtAhYzOwQMkN1UiPt4c8nJv
PwFq+vzsWuoGA7dzZvHNDxq2twpkOORjwDXE7iWeRdeMzZq4rQravpO3RJABpcx3
cZ4jRsHMAUTceDOoizEDPpu21M9Pc5O39Hq23WQcnxLRKr3eqoabRvAVaM7FkoOZ
bvuGxP452zwT64q7+mhN7sEju5sy0cOuV+YiyXWUUexvb3uRY8iaXIA7V0Uq7b7s
fx1fSfs5lPDyNN73JJ/irTgk+zLSJBAzu7zUVJBsbQazUWkq13/6qaWyLuP3CsLh
bStOjOTNb88eDtMTiP1ZbGCJa4qd7493rbG1qHjAoYRuu0EYzErPa1p1EJoV0LaG
ndy52soIwSsb9AFDRLDhPitLohIDq+3ZJ23bqTi3ZOjQeUkTLhrM+R+YZ7abok6S
3bdOUEmxioMrLUhNoBDX4K+/KAXgUN4qNAJiNXYJzUNqeencXsHr9qGAUJ2ZWPHm
5bMVRsyZOAuFJaTYJUiDZxNlxTPm/Ah1/cPzeS8oQZaAbGZ2E5ZG8BUmJBK+ku6D
8KA8Mr5p0jhz4QHkafuFVUPTnTExNBclimT+mLxkwNR/T3aK4+0jeuJ3FyN8Qw1Y
65Hao3BVHmLz96jxq4DlYvW8xsEHTxRtpnszWP5CCLMcrLHSgAmbXaYd+eB2BbQS
7LNzASfBKRZ3muTOFg/amYiBOzKKRJHvZTPuQ1KPNNk9FhHa1gCWl3waRLYA+pwV
tT0d64Ta5PJJl28TIbUKYdJI6y5/KybQQ0PDMRDsdP2l1c89+mQzTyfHg+kNeTI1
j/TpgtHH8p4Byp9eexE7kS1nb5gL1N2CukznjI9OXYy43eN+apH1SyG7H+OBXauD
9HDREcjzkYtg56VFAVpEUsgSLWQ1Fs+iQK394EkM4DsapDTnpN2jUbIjG26zHow6
BXW+ymRRqkkeUBSDbjXrsGh7SDi+PYUGYHL7erfEpeyGaJ+9JoGQ2iswf0XZiqhN
yfxymYPoCZoD0brOnZimFqsEokRzz7mLruwFVmlGBdcM1h291hc9oMB1dp7CV9nU
qUjKB5X6bx44tz5yVZXD3/9qdpWkRmhyMtFHOm5fcSNjWk7ObRht9PrZiHpA4l+E
q6wdddOsKkHfltCmlqvEDmB02a5jqYXTq5/zf5WwZI7yAbkal9Z6lqONe+yPBSTo
QpJU8mG4UHulLZutnA2TXqzjz5JYYT2ewIHVazlucCYV6xER/c62B0VWK7+ir+P2
qgsifKJ7GcoYL1iLjK+jdvXaUc079L272gThRCs7KPBtoZ14KirhYkJZmi882BdL
So+KgzFCWo8/XrJ8VKyycZ+gw0nztaLUcfMWPC163ZylIYANgLN5YS1V6ehsJAu2
x0yM+CqzPj5LMRjA0n4tG1BSz6cW51bGw79fSxdI+tZukHN6DuQA0yPjOP+6hS+R
3hGy4wGSr7exQ48Qz0Vy65UJUYiBbEgBFKIQzW86uMAWftIRhRZl8zWcrsllamPo
clUsjjQJwlzC0Bj0FQz74JcTvrQc1wGDcZ6Ha2TlsMy2lzxMJ1Pquxm25imjLC+8
r74f3YfmqGy41AZ8DI96V3zKG5CicysDCcGTiCkrt4eq1bxgREFb9vHjtW3jx4IQ
pOGBqhRDSR5KSk5STYP/a+e1prc7pV/vy24q827hX2KPVpqcIFSTUT2e2UqcIbOP
O5d1csS0a4ZI9srmYIK8F1oqC//JMYEaBZko0TJ4c/2aFJ/XMkFqo6fTuu6LbPb5
PWTxyddmjQ4s2SlBS1N7VXeR+3XoKi5NkGdQaMOGtPsal2jcshKQ37+P9G2eauwk
unWynrvpcxCcZ0BTs+vRrlsD5dB8RRJt9RYhxMOWwgPYW+v/6vAV9VRrFA82g0tb
q4cD2YUB4DUcO9+MwCtFS/ns2EculjGJA11ZB3sYmZHzYTwX2ka/cAFFxuaYWDvQ
g3wG///Pn1hr3OUrn29a6x8XyKlnABuqQpJxfdpZjHtY2+RZmULrOneVQ+mnzmhh
1Ph1q9eBgI0vVlAVMYhlePoh5C37GUKKRrbzD1uSYz2hk/F4TiWAVeZXayOo33O4
RhJjNpmGLvMvkoEVrlCP+On2iZkEi9mxljO3aLKf8G+CSAojRRg8dBV9Ocly/0LA
Qe4zvHGzJeWTe3JuPTGCON6qqypd2cj2DWC/ReNqMhGOU4K/ToDlL0UYwd5GAH1C
zuPrTunzGcXsEFxicAK4hnhAVqxKWPc0uOjjqzzst4/S6HZi9OieKsurpaS/MrQU
wPJv6Y8nXUoCFAuUv0rF0Q3KJxa7ce5KkoRCZeu4/LKYW56tRkLp0gt2qQ375cBG
TKj7IE824ztTsqzvEn+2UKnGXava6K00tGdWBay9JRjyk7SDpgYgvveso/uiaM6+
aU893J61u16cIarnsmP9wU4Dc+2XlK13YpFQu3/J5lMoaDeaVAZDmX4toSXKcgfU
UPrmGDM+81dsLjQt2X2llAiJVV2oTIkPwpXoTtmonZi95Eo1Wto7aPEv0K4q7yCx
x0T0fn9Ge2RKaQpv7K+79crhxMtdfkPjyIGPosxaswDDnLm8U/vJoDZK9tSNvBlw
35y1BEbr3e03RjfMQlLaH7ihUSdgIUOJcft38Bzfd5WYHCD1oCLruIQbDiHKNKcy
dqjr2vk4ctkHL9FelGpK5od0KT5Oz6t489K24KlUiNras71ettMoAT89Ca8UYgY7
qx2Xzal95n+EG9tD59t05ZFgPlCifiwKDIQvdEtp5mVXPfdyI1ro2HqHtOFUpASs
gGbmDaUNUl6GnHCDP80WZrnwvGl/TBP6dFG/eHqc3Rgd1eCEOmN3GeUR5HvFyCfL
Vg1ycWMrvsi0mdIu81DxXS1P+iToRpQHfEFaIJ3mqxdOPpZnRdC3XP2qI7DTlLkD
n1APTEP8OVVKPk9uM8CWc7MClvhHkmkWv46XTUi4vxIB1cLcEkg4PGN/B/1ueDMy
5vD12asWVvojlgi8w9MpAbjBRmcze83qRbwf5ry8pblvuV/SCrOEDrvrc455/wW1
ynuIVZCsYuOwtT8WhMRI+wdZvv4C9El7ys2JlW4G5afVipyea/zhwf/4ObkUQBkI
eH46RNXQ6IkOJ/1S4CxzlCSXew4M6jbG3qFWgPQHYdIxZe1tRQa4frffwuCIqFaP
mI4pLIalzR4oM7lvHPLRhwRDWlsT59VOQLnyabxLRNt36X4fMIDNj4pLRgl2+1cr
9MLXb75Ks8bUEjbFuD9xlGnLRyErXUvY3yNT3CfY/CyT/aeIkJinm5PaES7MGBB0
seV4OZRlsjMxR7e0n81HozdeIFOgylrlprWzBN1mUHGNJ1Rpt+wo0ULcGPOGm20u
GP5VUnqeRV781rJ9VUVjJTqlhnPSi3mPmo0u6KWpbZXyTTKIfktfgM/6dfbmZSid
PDj07liaxdK03Glj4IXRtsKEa86qtmQwZG7UFvgXMsN35W6niRIP3ZVY/xbwcqGk
NqlMBcZgYVt4jDDXr7DXEJzFihFzR0EYIUZRV9mfHwc75xs6DgoAyTShnvmx3agX
f//I+UBhBXvr7dYUyKP0DeyHrytIog1ZFRSvkl00ZKiHv832FFRJSHiQOk8z5WOQ
BVR1bS9hnAoebFKgUJznRZi9w9FtLLwVnbUBKdEwKpqGk2yQM0vsVlty9UCfMIHS
ZUL3fm7S8uWZ/uXNrVtvfj170Ru5OIlKBfHCdrJKc0WiBV+a7HR+ThHYTIOmnVuY
fNGCv8uAJSU1OgBcJ5D+nFw65iMs0l7x9PKaQXqn3tw+rpRmSfUqoia5TQJHrycp
nabqdxSWMWUGIUOKSs7QCkgrFdKyZIEvLCxRF7ft8yeFrB1InYHfzHrt6I2URtTg
URuDk7Y7QkTvoZ31Nl9PGLwfyW0TDj70hzhpg2RWYv8KRmZu3ScE90ZrTQQRNvJG
llEHjX5mcUXD0No+8OC+HtUGRZVl1NrXAOeuRWwFLkcKk4OlHQ17tdwH/D0JUgvw
tM0HeRlkUgNWD5FzeVqYadQeGhCB5dmRMyWgMtLsXIEFZouY4BLxCCwTfzwKXEPE
HH43pfvnLd8VmQPNYQ3Ezth6p4cHmn78kvBf4C/jWrD6eOFpkHymMBcoTGw8tzLk
O/k5pRQ6qR4z9ZYfpnxFjc6Jmul7zQLtLUfBaEJn5YR7Z+8kOTLpVvc+w0qhw72A
1v/ghTYeBzLnjoMCJr6bANntyV9zyFCxKhLsbfcZ36HcHWJ2m+C2/JH/yvOKgkJn
etyjWWSty/uMIln5OKUwOCRl3OKaj3KebujTpHIqUpephtiYCSWyghphv9PcW9Gc
gpxxwqObauwDF6Le/LmRDhJ13JK0x0lOakShInQl+RDpUM7JoaLjpsAYnLgEhMW+
Z4ucKuAwUGrXxdXPsa/1iT5F8V0fJnheEfgPEWpldrPukCVsfi075qz1/jOTeEE1
NZRNd8IT7cWsO1pTLmFnWuE6QAJhl5rtIWwYfFYjTklaqyHw52cGpCygKlKu86cV
wlIJ+rbMH+YqHcoAm9tMg7xXnUfGYL9M//RUdZjgxHkdit2sd9hMk6BHGFMTkQIU
3g3+oo8XQNPf4QYBeuFONVUoNXrLjnsX0CrMc24fVpycl83+iQWiDJYP1wBL1ql3
jbgqUIdUOr613SPp1O8E1C+CSXTDVkZbsIZhnSi9A20PrTXftmC5sCb0XT3gRplO
mC3k+q9aWXghyCOmOlA5ODgW7BzQD62j9WHAN2xqRfK82YvG1AJCoIsiyBgHl2Sr
FBJsaG0+zdS+LPZ6AtmNoA+PL9DCfFU1NXj+4M+1WkH1xV6mIicwG2nijITT4xGh
FWKP/tTRJuqeIcvMmw19tTNRz6H5wROGvhrpFXPNLgKq3GirBAkg55FvhDcZfXLc
2WvALeq8/dvZfdH45RV9hSvxwWjyr/ySU9CeU63P0vBeIIR9A8XACQYfJNVM4T6J
vpcBLk6OEorosVmp5miGZpaeSGAVf78xA1pW+bu7vFvBAcW1ZYcPvdpzSMXf5hx4
ceCWnoMWC6zux8SZF6D6osDMapQBvSxxNfw+lrSd6XxbsVlHJLD+t6LXTdq4oiC7
Dng88Jne/7japPLys1SwFBN5IFNK/jge3Ilthlrz+80+/Ig0EcI4Tw+fiP+aO05/
+sMMWlFnAuExoGLZivY2J8Iyp18zTJV5WxN6QsgZXrJHo8dolUmBljUY9XxQLp14
S1l41RW3g9kA4envpZmI/vfLJNRcA6NZv/MXzhFcR5xMdwrNCOFTZUuEzx5NTH5B
PA/08ViwPINXAafXf9qb7xuczMHfCKMlnj/Txl7VtTXYqo+WOYYqtOVJA6MKNPlC
B/xTh8h1oUammeMeZzHDIQWv8VCzvuk6S8D+XY/sAeIuNu7ImbXWo6sd7U7q1cai
uJbMsC3WP9gKhHD1mNl5YBL9DxIspRWjl7LDHF/j9gZgjcDcCBgMExp6lodaatWr
upGcl9J6qFGBKl2NQttGVUwNlx5z1HZ4Cb3vo59d9K+nvTom9fsGugyegaqcmvCs
7WeObRhNpPCTDFEJzU6x/1SknIivBark7ZNKhQAJBuxn1RXz/SfoZBscHWwSxPKx
+fQVv/XwowCLTgK+Xn5cbCzS+kyEhVsZCtDgEI2x37C7Tlfkhkn/PXK888s07JLp
uHlPJqXx21LoBx8HBgVPSamJ7Gc0cFSlDTw8nwct6p77Q+Huw3IMf9z+MLfR6V16
Mu5dL9cF5d+bsZHSpN0aW7Gztec5b/cf/tPlf76OK3KBvQEjMMwdglGPzVt0NyAi
7xcxYqUKJsTMYGRqrPDMDcAlrODdJid+BsB60LaQdJrtL5nwbS1QRcoTL74PFCCv
8WMPJ/Hm213Ssgnn7cnGHlES6eT+3ZDYB0v0DdvcecqeUJmWyMQf5ynxSh6waavY
iQTS0jWxmUNaArthW7u3M3s5ASw6YePo4rzi2PMd2NOM18bj0zJpEcQpCCSDpwSo
Q5aD8uYxX4vORN2g6qUdC5n+TSKZcUOZ56r2MSOy72FUClVXc9IWwX8VlC6Y6ppE
2uq1CKz/cHOVUH/KwXcqjTJrtbOnf0rNY1O9kLlwzuMsqw+7KmoRodnuRVT/YxGX
q+aB/WiV42LD3+zA01og4FJz6GUf/WbP/SPijykMp6+urkjSyPux/fPlbFuRUv4z
Ce33vYGlBZH5aKZAdzVGB8Pb8x6/DvA50HEyIwV3oWyHrzRYw3P/ds4Me60qvGcn
BpEX0RqC9oAQQI/TqYuS1ZSEXd8RukCFHiVRfz6h9ehblq5GjnNMHMuwlQK5xVD3
0VhP+SJNirMMxq/cL73750CpxZE61kuOI8Y722CwhSPLA5/ZBwNIn+SLs7tsV2m4
XlddEFDeOoxqm5ccy377qgH1cWvrHKGKRzX+NmmOglfNV62EWBdFGfcmwg1rJTGQ
Vyq1gDyh6OB5FCkGf32q7QbrwCwpE24y85h3OpcuxW2BPgeKWkz05YGR60V47Faa
u4xFQhogARuBMNW+8+AmolbbmoiB7fY8dGe3tKPL+4La2uvSrM/cTmqTBo9Q5nFr
4EokqeqaP2ms9GeaZqpNkxFaNJGt6BXaXAnI6u5kyJ/sY+fwN0s9Bvcva/kq1j5G
J2Mw1M8lc0tKHZ8Shltdn70y4dKUSufTIhXs2NmU8ItrY+zLaaj4ViQGCcinq4JK
bDA8zmpWdQ+EdrQAspsLd6F/RP4Cgt7yhtU6bDahWiRD9f54N1XvxvTMpmbD1B+D
WkSkfJuxRfCjjXoyb/p6haAImQ9Etml9jBM6lmBe4Ub1K7r8bxWQXP5S3yy1YVIR
tT0dVVVPS/gtUIw9YWGEH2LgjZiBjYfMrMz66o95UbvabxXWTlsOya8mGVOEi3g1
V6wYi0p5IUrjGl5kzDFnNpIn5tu2V+Us2Ln1Shw8IUN0faPjX7pSLME7jy8EfFVf
c4Fm8INa6IuWfzmVgTPq5cXZPUFUg+iQP8pCVxL8eF/qBDI/kTwJVl8s48cIV+mi
GpWshh2uOnBehX59SJt8ZRkcUydb+36vn3pvhvD0Q5OQSwG2KZeHF4t7lSTm2Vvt
K4eD3UgjrSk/AW+0LV2BV3151BEXvu8VFT9T15v+IUQq+1DYdv4X0pZ6XDwpt3uD
DLIYtT1xSqE9zNzrpShQfByJxRUtlFw1IorQ9GJJ/WZYlzygKiOI93aO5tBWeaDR
ftSktgrQLAG8PB6g4jJBsU0VLERtKcjlmfufes1kVSE4rpcjrPo+A3UBnkDX5S61
vuGdp3il3JGlbEIc2wzZSi6+AuPPo0AfnpxuyeSWSvTH3WJX7oArsHXHWLy0huKk
8JIAYhXmv+fytqV4tQfyIXs1nW7Kxr3CqewoLKSkIfutmVAujX/4lzs7LGKJErWt
E2Rlkrx35Jxl2kqpubjZ8u0wZDEf5ZKaRNeM9S04T9eCpNAcvvzITA9h4B+konXE
eSB4h3pfRm9Bv1oBWZ3/C7sl48H2Hkq5MVMQYQY2AH2V046JY3TZXvAf4sFms/ph
Tc/R+8h/QnJUJOtwaqJn6dYYGQnrwqrxMvDaAiYegP8RJLM9Ggr/Qo6aGv8FyLUs
vaigOG7B/cYYAz5ncaz7C7fODcW2jWzrjjHrCdJvCnrH+UrJeIkITl+d5/1Qo8Dh
1+eqMGl1gPBDh756HSpwrw3lJ0v4RzeSi8FFoV5uafggF97qKrLxZ660ncPBIexz
evBCqbT5BOPJZe4QIoCi3GI1UHsKY7AK9cZrHQOIlWzrEt68ZH22n+dVX+q+5fXB
BqDBszmP3B89ntRLvYYUk5iJCYzrHctyUoqrLAcGfvy3PgiSKTSi83Ihlb93hRBk
TuOx1ffd0U/XaLbdMOr9pMr/hYXEOt0gXAsuX5/YIEQMPdHiWds6dcuResA3YXlp
aX2FjgrWpY0AtGGBJv8Q0PhGx9FONe/hZfpETdmbd83DYUNUnOT39dGA9MZMQOWc
7oYg9QstTgd3V28W5OV/bgWH3CNvIKcDjJM+IKix183chBnYpiV7Ei3tVGLtLPCG
1Syx9SQt1zcpNlWuSNUTJtf2NTc8df1wpmYf1IBQySXBjO6gYgqwb1GupcCrSDj0
ZUe3xrQMek4/w7AK1CcYG4Ls2F3NoxyCrVPpYRKaIgYKES3vafyHtUfjrUPqUh/8
pG0BxOzUy/p0/qtFw9Wb1vfv8/WYAtgbT1J2rw8l4onQKZVOi6q0aVRLHlNWWedS
YJQllPyuzElSjehjLbtIkwM74mvIXUtaxNqAG0oGokTfwl/9CbJpNa1IIlFtDfXq
XQBEyld8rPL2ZDpdy7Gqsl1pgEnUGLFg96WvJ7dl+ypAXHM+/v7/zBPU56zFva65
hfHLhbtyi4x11o71dI5P9m7PNlE8hyJPdFGE3rpzV8tcn48XoBntHKgV/dcYRSSY
+J+l5GHQXFFWhOYk+aThlze2+DRUYyBHpkgiC5lyD3O26WNalV2GnTyOL3LF1pjL
GmyRyoUO8p6KeHLGsl60EjLCqfFO2tvm5uQjYhZUbuvimKetzvCNHUyyQBht1g2k
KI3Vw0wruUlvPUWZ19lMd+sNySHv3bIyKjfRCg65LWXsM3VwS2H0N+6HPPDF9oWd
63GD0xdWuxr/b5qXxaMP9+WAlMkfYxGM8Q9PjYjX96Zlg/wxBewEZTEEinEA105W
ouL2JhP+kEauFoyxNOzMTCqUJLQYe1ifEFg5824ntKgtZFXZKJbJkN+AOrMrfs22
Vi2EVWzlsIXxkAGVq0wUhfdosbB9B12fjsVTycGetAVNen60eVP7xOkQTasOWL69
whX/VIk9LuE8RZs/RWUosTkRzeJ2HoE2gro5Kw3beqVQ0YYvHrlyfJOJ0PGp6kEC
gTleOfEYOEINWvPScYPxVHLkVjzVcPiqOHExIW03NuiEjiTNvhS0z6a7vIczEpoQ
gAwta8pgTiMmKKXobwY86EoKKLPHtYB4hSFKGBErIlWlYiYqnFU4QUmwQSy/CtwH
QMOuATQMsl/BZmjI5LxGGtXBZ6bacXEPtgibSaeSZQgWFDdsM2GSni1yuI8/D2nI
jQeZ72bOs5OF5zjZvZEyPIAV2+bJWniMSQfyX32MnSZe1zTdX7Y9qBabLR+xl0Jh
PteLx14hEMcJEdqxfy3XFXU7LJrUzU3lsu2ulkmzNsLF/+cWZWxaIfZp+wI2fGUv
LUMR4gJMCyNJjOvCgKVlM5O1GOM+93jihHTlWqHErUMUGQEN5Bh0Y/347FR4HWzb
T3JEfx/wjVPe0YJuAdvXF1mR/K0Q/2f2aD7UkCDKa/E+XmXwtaVQsy1SOFBjyZcM
l9qoSi1109obaTomfPHkz1cFpWd5f/53o9diSxWsbllIPaw9asrGAqkzuABpHnEy
lhZ+reJYpHhh0RNE+M0E8Vqoy4PwKIRxjKKNohjZ+P6aaVV5R4qZoK5Q5xL27mnC
pKYW56dewyA3zooMGlOYUYG4m3giU7FDQm44gYUuMtYDgti8vfF0AFx6Lzjz2+1u
mO2PX3hhTGnMX2fK/5bmD84feSS+Ygf7+EI0YUSFEUe8gzB+yaZ4m0eqr+LyyPir
+RP0Y3hoPn9IHPrUBPHf6R++Bbrz60tkAw2zEiudsvGsn+ZANF47Snvy7mZRo+qH
F5yif4cigOUoBNYMZxFGhuQrrX9k2xAA4jPph9FJpDJ+9AnvMYl/mgLmxAukRsUY
SLayVoTyXPbNBYRqjdej6ij6AXTroJ9XT9ERucClwtF1+mibZwFipXbORBBGPdKY
YfhN7SQ/z9rgTmiQowz77put+9T79y/OjknwyqTIk1UP2kgBQPdVMpNuSkVz31m/
clZdoTwbIy3KWFyeHihDh+B7qZmvXVH3JD5JxADNijldTXUBP84/xByztmGOLbmV
c3ioP6reisQgYAZB7AoDOahCzDfmaG+TJQADMI4PZheNRGLMzU4BBKMDYz2bD0Y/
lZpdjPk+17hI3oPc31UayOs4G7+BikHjTrpcHaI/mYNTzHRXmXO+0dJXlIFz13+0
CwQNwL7hC9pJzfQab/lwlgmg2wOGTCAI+pbFOMIBY6fkkOKwQh+AZSliczeO+Ck6
xe2OOzgtPCfwsOKzZE3fJZYNgGTJKpDsFBrnS/zv3JGJU4xbGm4ctIxAKc1+oORn
0Qa7TKYRS2ztaf91Q0zSFXiJcF8UN66pb8jvS5lVy1qyS2jdKjsR7B+R6HNc/f/W
TzTYnIao9EV2zyMwcNa1PcufpJxhfAUpg9tsODjbAC4H947CkDrOXHSFtnEGIZ0O
D+pmIwZiE40byhfviKNbmw8bP7wohsKs1R1611HN+CRNZprEnmnfmOvDmLrcbb29
hd+nrtArx6lyWSKUEMU4GvVcyY390aLdI/QVzShfIs/M3y6f0tCSR9QZtQrhi7zJ
JHIZk1EP4ABvOZVZQUXwBmDkPOx9ruvzd9ySiRMjxfVXea+P+ZmsBwJMPgZcGZDr
4xYYluB7k2o9jXyYTbLKjn7W7F2XssaCnKkSzZnI9Z6ApDmf9oXRSyww9X4IueMk
cKDcyl/QVFqIb8X/tIpCCIP5yO04YuMF3nCNtlM2KlvGg1QmkkI1shXkiYFBiMmp
Jkg+pctFZW2VX7a5OZCLkOHHA0zOrDK83iLqIDfKK8T1BbpE8d4s0UycKj1GZHuA
ULJw1CCHQDNNhuySkD6qtetbjFyNRus3P/aOaE+pT9bx4ai99bFGq1dg6zNpXvgQ
visDLjpdj8rOKQOb/9qUNj9R9OyfDdIw2WLhIpWW05QCzsZd+oMWmBIQYddveLq+
iUFH2mBIFHI44qVV1BE0YEhXzxysVPBLZgA9NMSJiPp71PCwongeDrs01LKLfNjA
5/B9qTYys5VM7UM7XdHOKfvJW34hXVCpxs3L6+aOBXkZXmqwezYsdlCYgl7itHlp
XrT1DL6vkljQj4YJ9pEh5+BVL5GyFaWzpdo22XI4Oh/qCMXJH5ZfiP93HJwV4v5D
HBDWrdDk2CM4mBX94KVK9kh9OW1ssFu6Klp/RZ1jQBYW3WZn7KCL4q2TQ0MDca3Y
AGOGIE8AP2HhDPPhQkvZBU82FAoav+wO+etOfb76K8Cl2gIywdrhG7MxhB5s0v6P
4uwx1HOKWYYUYoE4iR2tsiv0mNAl2kCZ9eqfxWyDenEJJpAC7TKlpym8DSY5tMP5
R8Yx5gOjFq7n5RnTPaEMQQ8AWqGqTRDeH12MZ51ycp3D8Jf35P3fv4UkeJl3WBDY
eFo38pTkCeyC1RoFMttmEBjfBtAMDYcgaSpLRXwtyfeVZCOBKbcOdLLXEIkot202
UpqItaw8SmKJxl7bl4Km4BORsNqWKm+pMH48kCDf70Tu04t1VxmAz/73PMkPhw6m
2m+aFZqkGczNn55LRhP8cjVqx8vWaTlfKBUd+EMYbLFznYRqInDGyy6aYIexSPRi
mY/O3OoLWg82TWZ6dGTqsw1qJXvLLJ9e2ucaKBh02T8QWj925PPGfS1XU5wHttoo
fXZehnwDaK1+gzBClEvz4ywmQpdd8w4IPLcFhHvJ5PuP2HMdC7OGVOg/x7eAsArX
LF0wAVOhBSGwHQyOe9pRcreGgv7maiI+HJYfFWjfV4eCtdQDVvEVDtSH9f18A6s2
scGXOVPAH9OloLjBDrJu3bBgmuicmIovIlbbcpzTrcYhk/euo5lOPucGGhTHuibF
LP1OekU57pdoSxXtzq576WzaBZhnDV/9RcqoZ1kZbia8rmO+YCeHTGO8E1U23Elv
gy8AfpkvgjFjdm5W8e4GxLI+YbSpKyWlQsj0bPiiczvBDM90z60q7xpGW6g42KZp
LNRJ/ZUC5Dqp2+nRJVVyVSHV2rzepPzgQSuZAatsVHXJoftCIYyS4XjEoEioOfNW
/HWjWysmxFZjCoORntsxmcM9QMDJPXD3oZ3FuY+3wSLKrRHPQZfzkCItrdEEW6hW
7z9XPp03cxJn5EVDhwtJ3+tt1AHprgY/XFHhgFV9XnySbVvDxs2xvzswUORMKGhV
nMhHbtc4crPRNBapjLA5MybctQV3iEsbD1T63JbjeEaqrA9XD8sTs9gQS6K1lniE
cIB92YQUdRbgJV4twJkBSJovxIJsIng5vdVRY2DKiRlaXfhlwcwQVa+tZQIrtvC+
BMHDkbzWkPpK3gFEAVSxl6fMechy5BIQBSVSDWpw8hZdmO+G5xVSlIMk2CmU7wnf
pqAyy4IhidG5ui8KyQr3XnOOwdH8un+wu1KkFap4R6NQalit+7JfgBsXYQ7mZrjj
iBGlDAcME1iRgrgPlKEAEmUU7miCtDbepmJQYAD0zHwA/aqDVm5r/XfkqxpV5nW0
042JJhgFPV6eQATLdYpaADDEFgEkOYpBmRKWpYDbWOZMWQgiGs6hbVuwzpwCG0mW
clsHZtHss6HhV1wbhc6Uy6Fjguy4WXu5DUKivDoBBVjkqa0sZGmz/WQukC+s9Q5s
8p1KJdygorXHkg5dVL/zNnTFpd7aMkHLdr4uChyNgXsyt0zOXBfxKHcQPc1oWSPF
h9UGHeGsE2RQiocUEdI4kn8g28Y2TY7UDCGfaKm0ler8hgMcYRBE6s3B3YzpElWb
D3yqewHlXHA3qEHK8v7LtjfnMaMuirX+9KHShbeqEOEPmDixhhfTGX44imzHmUbA
raKvZ1aUAnGsnD0LXIoozx/1akeUGozDttF3W7sXmhB8MXoKkcNQGi9Chm0XhW5L
kNxSZLcx1eW2Dc4ymiz3oOsA0QgKjZI1ogVbbyBBxL4rNNdhtmfeFuHjYZM4yxf6
LcPPuBNIu7Ku4ogxnaUWst1iUg6MS4qdd3N12Fcd3O9h7A2jlIFtD/ySgtD+wMKF
7CawWOY2OcJ9IawAPi1Q0sko9zjS2nAc1RNTuAq+ECFeRsw27skMKiguHidlGazG
L2WRWrioxI4wK5dYag6xQd9+rHank3nS2muRAiC5r/bxlgCBm3PmznU1aScKekad
Tl7H9WO/Te3I4Eba/OOkgPg3ju0i5w89xAu2jIBFsXUt6DfJDZ26kP9JaELIFddU
yN5GKRGwLaa1YTqaqRIcmOzualQIGfVY7nPv1T2G22TGAm2bbpVSqmGv9kWEv/Xi
+zq9vP7vfa0rLSrbwzQE/nrFPrgl2LMQ4ZXJCjS90CpE34lOctc9gN/LDN7KBV0I
5Eoo4hsjvSQcapx99d0eugg78DMijdh/GFmG7e/7AL2YeXq8ZZKP1LB5qgBzEqxg
9GQF+nJ6dHQuIBfiLY7RVHyjTnRTgRd79JqlSw6MOcmPmE7E3rj4kECUb41iO9O2
gljuQQ0RV1z6AMB5Cvf9VIOtaZ3woBIHkltJGwtFyaalZsMrxiPeErFa7n79S+bM
KgYoeB14Vt6f+MeHTYXa0gh28Sv0pJD4AcNyPKvEq5OthyJmmCLjn4RsC9WrOX1t
qIyIQ+LCoRLNcGHan7FUsC8cIQTDAhEm3upSgM4gMs59YsjL5f5K96JMxkHsfF9b
7+Z6RvIqbbz4wdHrG8WDqpmDa0hfjWASSQjwl2+TgtoLMIoiWTmXgpTYUSI4XHsO
/wP7XCRwWgv5KgOXVwiZwdHeb1zUHCMczzRcH8G/zX+yWWZs73vliENzp2m4TDPB
0xbDMTUJDEpqgSCyvaXBmHRh0zGKo1lKqduxbOU+1ou2xFtJIrZY8KCnKhB8AbJD
fykp+sLIasSFnUZKAs9ijAyxUF1gxiqPqmjhp5OognWXaPbls1zMRwb7It0IfpkZ
ldV2XcDETglHWFRGaVtpqMEawbCkgDDOTCRK/9/nEvnDX+XDCIRQj0YWbmD6IZp4
kEWbYXoDqsrMQC0WYo28uIaRTzPYiLzzu57jByZDS0atUgkQ3zGp04vzwPyPu+dT
1/3FHNoLIyvztf91nrZfDAY7kJpSSJ3B9N47jb7etIsLP/qbTaghM/cvBQiWjx3c
hjhYIgaE3wDcOVgDpU5PRyEbI++vPVqgDTY1GQsoG6zgfZEVcvEm6Af/c5wkb6mq
RCfQ2FmT1IEpCQGXToD+3r2El5cojslGd7CbFXXFuqeGvQlTub+2O0Wu2BGTkZEX
Vk7p534QNuR1xA6GHuCyIyTErj4Be2EMycOZQjbBZJz1FjMrod7rxmZ/PIrXSXxd
TwOCc7nJHUy2gh2Bg6GqUwYCrQPFhALvCnrNrTI+nMFFpctiR/xAb79UuplAJeTi
1vHKjHMWDilqNKGGw8RwMAf1mDg1lsi9YD6bQ6qxDXzqj1f/i6WOLLVIv44DJ7Wu
NSF4c/q7WvJsDu/Rfheyg8XEI605l65J3+0tP+TdQJSrNQCjDVCXf0j15sixjJba
5Aq7/p7D+JmYdhzbGy4qX7wPxr8ITb2eIOzqKYY7o0phD2lKmH3Gm7r2UATfj5FG
7TlDRVhJ0fF6/sXltgJV+NyK7XIvgn5TzdUMSsRuzNnfDuHqHDGnxfpioB5Zycdt
bzZOzASJCeWtmR6ulpg1MjdBNWJ9yPJR2StRl6dlSe8RLZJv0Lpbyt8Mvu3w8RHN
ygjHfa4d4/kC79nlgZX4K3x/SWAma4is/+NGy3nVlVWMh92X7Qnf6Z3hsWAlIKeI
SYVpeiNLGwMdcO726r50INz8TKTrPp6zvhyhD3+vWb2L2hk0v+oI5pkI9OsIs8TL
fQT+WNcoClDaXHxDpepD37tPUjQjSU0qanym/teVCZkJNudeISAqwzl2eTbNCAgt
lh1cMsTXWvrbWHZIdZXgXV5mXyM5oTDBNZNPP9/w8UeapvDhAKOKKaF/3Ig9rt4B
JBfGPfXx29KheWnBHo5SSKKq0E1iLqwXI0syZrdkWbsAb+Hh7uymu7lbpQjbzU0h
N6YKCtc26wCyZkMGzjNGrWPDU5cSjyFDtNA84lOTK1Km2z+a+IE68/3SyR50yEsJ
3xxstPo7Qr3YjoXaHx6WU2z/pFQgm+cs4bOATEefnNyFfqAmTYypFlIJyOGzkV0Z
JBQQ2lIjMVShyjlxtAHtLHC37rd2F0/1SzilEDbEqHoozocieYxRK0qWeKp7/PXI
qNUhXyxpdTFFQ9wWP/B2sTuSLjrARPibMrxPkubQH0aEIxxMkzTDXXgbEolKFUqO
SPDPqH2Dqco/8cL1oTXZ0AlU3MGhFUT7EO30byJhOoObz4tpdXx3D2xdlh1ZnkLD
5LvHS768HGzTbeQD68ZJ6UslubnbXGbULKFOV5fcXzOUXmYchftH2kmOkXCrR0cV
uyaE/kPRUzKjILVIhodMu3rWl/BaAWDmHV3uRHkyNtQHK0R8fzq8Q8ygItWVgyjR
/5k6RyizEfNLv2inmSJPmL3cFjsmNMaIl7djGaOc+VPAuSRFh4E2TjMZcZyDWK05
DxtIaQ4Gy5TAiaKOpENAMLpbVeQABU+6BEd1B+Vjx+iys3JwbZwcCbWVzpF2rdNw
jMuZTSuSmc/dqXrGstAkZP25dhy7r7G6MNXb45bbS+bbkGK1c8z7BRtw8N0YxfAS
+JUn8Fgj3/eIfNqhFkG/jRjRifc+9k9UyqHJtNx/384xX4jKOI9K5SMC08DlwvSn
1iHjm0MzhNsYJkMf9nCD5cmRUSCJNJjO3qfB4IHSCFVCeB8YjFr/eGHPmL1DCeRY
XsjaOr2xD5OK3/YzDq6tqiTrJDlBg+UbdIRsoY7Ox5xrcj6ycO8roZiSid7/hDjR
7sQc1jOi0QDToRGEF63ty63NnZMHv011fSrCvuJ84tYi25TUnZcNj5yFtbxTd5yl
iaKlhAnz1/qZl7JqPf3tf8+Pv8+MEC0TlqEM7Xrcg3E6oBlPkuOH46pn0oM/SXOU
IDQsVuIDCyLVC83dUfVotBLaQLFQZGCIoLBBcV7qDQrLTwBdXUjIGWUiI6h6TL2w
2BAuwSN3iVu2R0+WmD+y+LQeFU43PxfgmhY1QmO/0fmTr9XGo82XZsaR3xUkpp/K
iHhoNPBkBoPdm2BaAsAlJ1WimXigu0LlOD6zE3cQi2KIsxwCcrOlBpbnP5VyVpXB
+dWb2WMmgjJmW/TH9dbILZTCDgg+9nX3hYI5eLUnOMH6uSo8G1GMKtbtIO1WLLUw
9Y3xX7Ib/DR6nP2HuDWFvlvIErvTxjcAnHW//geiL3zOLbxcLmghyG0gMYDTqkx0
B4RB3jccBqVspFGGKbOYRzI6iUO9/NOko27wHlSob8fO5wVZ4d1xmeR4N9AS6vCm
Krzhk872hxXzhBE7CHbEUMd38kCOEn3dlswp6KFhn8UnCzKjD7qcqHc3yt7SetNl
pcqOu5riR5Ob611o2xMtnf9mnJ4IzaeX+qXf21Kh8XBHdXFFoxn/YjwIzoOuInz6
16nBIDCphtKM9HgK9/ir50TcRR0Ro946t7ZMJo5bP6sdFyKPTI1YBClEe8Bj0rrs
eyxsc3L4Q3LcaIMTerXnhdY9wAQ7V3xyHp/8bmP7eZZZWhGA6YW23DH1kQzhtq5H
RKBvoRKBuS/QifHT86/Rzk5hcM4RCUKP8sDoaSi73K2Gd27rLnlF/SRcM1kqjhp3
AhGocY4Rp8KFYv0P9CKZJwMXSizAkGpEpqBl26fQqx9+Du+XfTjB99JYMNFrkJxX
hRb/EWFX/drE6gxlrsXVrNZ71XB8uSxmfg56eyttEITK3bhwniR/w86PCDBBgOcC
sNX+MayGOtZFJTOi0+F08HkRHSNzz+RLg0KeybRL9khXzdC7zG4NEEUlQf7tB6hX
qW5TIczThhslvtqURM1jg7n0LTxmMdXpVd+35VXooiOEnWuv+2d9Wt3Z92A2elmM
gt8SBfsZj2K9WNnvB4hF3KGamwIBzLGMUGGO5kT4mYm1ey0LcMI7lpPMCmzwylyN
2Q3k1ea871aNGqU7T6Rx/hEAjFrSYiuq/Ph35Uo8pH320Yd2tieWP5ukHEeU/Mm6
2CNfDKWAq1JYvq9gQHJ4s0FfDo0+7CK8IFGBFWR8spT7gZLK24Fs08m0XJdzQk3C
5Fs/kfmW1r32Rz4W8hELqZRTpnLbWnq4Koq3Aolh6KwTA9EKfQZjUe88Eut3KgvH
381wi+8YX9ylfh5YaOyRquIZIEWx6RsDmyLhqgmBbeuaLLycOtglZiMM/MvPMidu
ArYK4RWtjlkDz0zXGucfyHgnQ5oUY0Kz3VVdwF9cj3My4naZCrJib2sBX1NnYm7b
r/r68uI3UHaid3/Rv+Br4gfKSOJ4cURahf1XbwFRY2PYyb7gx4epJN/19rJxzgxJ
P5JsLz0Wb/9NAPU0mlg3LohAiPIwKTicU/6F3z+/k57eYbn8RY+PelOdl8ClEnah
FiFLKPPZ+wMNcafl4znEYV/YFEl21J4YRm+2uti6YQ76Wlua76yiNllhYztqbj6N
0stgBMeIOp5F98UiJV2oQmLt42hcqZ7uHkvPMkMYgoEW+QUIqWBoFGrEFZWCs9kg
iOZ0YxAoRpvr4iuH+w8U12nWnwd4gnriUi4MBusyOeaM3QJwrD7CmS40YYCQhEAL
EZiScf8IWnttnC401xew8/cEZnmEz5J+lq2BC+vvFsWg26HliJP67zfBQpD85cR2
ZIg/cIbCyQlsaMZ3g+J/w85pWDqFUsLpjtEgvqrQmOhV+Wha1mocYNWofiwCFjly
lYt9Wzj71NG/ipiDNJgozFXne1HiwwfaNI4rtMtJABUM1OU2rHSdte5mrNS8LWJC
Xly/mmSnlFDQL9z3mqeES+6dLdqo7tTwHzcivh8mC+zuKMYUdrNJz50Sp/IDotqI
Y7/PRlrhVd6HVhYF+eX6EKod8OLC5T8O2i9FaSI68TJ2otQxslnyhuyFzPdze2k+
uzG7fugw0SMEuXlyHn4M+73yftq8JKByaUm3BRjqEUZX8dRYNMCsB41roq95m4qC
pnu9dgr4dnEDsJTnxrggQIBp5RnA2e7k+EWggIZ46y5xmwSxzhmUVxm/FnzmuEPY
ORqPVjCQl0Mq3YILg1B+EwPi5IZBeRi05SoictP3JsRGCYtLLia021QuspCIkfcn
cnMJsdlzTQIfn5rIB2V8nxG7z3elwyVbqKv8XvNoDCDwpoUtgW1cpb/KlBSNcwvI
JT8Wzx9oZ2BWY9ZHymlnC/JmgoA2tHB7pRT4FkfHYHeZSSsZ4VOLXwR7zNyxZgKQ
PaYYSBeiVXloyNJPQ38YBKvVvRK8v8mUQ0yoDrNie9SPhTHYl2Z2tFRhl7WYWi6N
r2ai7uz4UjiifkgyOnPaGPF1Sqzo1CK1oZ8JeELskVLrX5bslL1inotihK9N+y98
N5gxbKIsDBFDoLXEtEYA/3QVzaVabYCAbqzA9e5WGknfzqea85tPLN8PqalnXQM4
v3tRjz+KTaATOB1rStUE5/4rRFrNQjBLwsTUENIpmqy1FEihxEcSIiScctvTko1x
RogehEv4DXSKEsM/VuUouB9i+Kth6Gw0+8o7yTiQFKpnMyFgR354l+Ex+NmKRfJt
gF/PMyAj3IKoxZk81nUqJAnHW0PHs/ZuEOEaiIsbyz8R9MDjP9hVy+UXpgXu2VFC
RKA17aQQ716EVPU5yMDWMZgu2/NjRzf5mRyxSzsEBjmRABQ6kFz2qqb90K2kUfoZ
nkCJ26riFho7sYX/KH0c1AT5eEpUP4UNX+I0wjodRAWHLTxN6i9Dlu3l/A38VNFn
41fSEgZpSg0x3SiwSSRC8JRzdTd5+nQN8zdcmrvO9LVR9uIrfMUPr0pP0hUIKR7w
fZf2ZHF85dvHHRUhO1u1UXpTKIqSNklpd34E2EdAIhNa1HVBaNjILcw2hAVMNtgf
8cilAvzah3JJTL2lDEKPSTUIqvBr5mear4aYBT7nQst6xj/BsoiPkm6I8egKquoq
AXMBNtnbHjXEjFEDvDwH8HCjXJ77RHMc066cRYkCp5U2r61akzEkfauLtakCOMy9
sRRtwGT+yAoOgA9CzSijyFZbuOv7KcI4Vy2sBckcXBwIa2OoTdg+EaxHQ+l3IHy5
vgMUucLA9p8fPnovQ8j5wcV4sdaN6GGpbWvkWSM/UFlB3wk2tH26sX6wKBW7tSds
J4/j9c++rPj2i3N+4ccCgKtuf9KWCHNCFvZCVAVrcGNJYY3VJQkdVe0k44iQdN4b
MjBBGIN9OMPejZK1Bods68v11rMU2cKjN+sXIpFTHmhcBhwL0mpamNGsWL77JQda
ELgDGO/3F1q4iji1Ep4PrqyzesyCHLXjJXVcOkgfXl51G1i+ztvaNgi5Kuz+m4pC
Exa3bJk3BS4b7wjNxWJVixh4sxzRaxEcEXnu/+IldmclDIAjBpHpxvQHN0jRSngT
tUkac0WUGIFlZ8Wa7bqseJ+Kw3GF71bjpSCG6jqmkYN7NlKn1y84wPu3AO1kpzRV
mvfAG+jAFFwCUoUZ8MM/UEk3lPzEKPTyf4C0H6H42csy3eNfujJEoE67tK9890h5
NzWjVMYa4dryrE4ku5l9cmLRhEUO1LbCjnShDNTM1S4Ea+9QcburFuHMVaVn7qjK
8s7OkOSgPrHlFohnaewMdpRmXPdowflVk5n7gJZOwSYvSjcw2xmxef17Vhbgq30y
6nK4vuFdFXQumR1caJONHi4Wt5CWIEnOai1eyigrshrDj0QxNsSVI/r4fuFAreSB
/kMqqpNNq5CHIeQN1d9aRuExFuI/829pTUkljQbl6Qt/ZKaVSNFWOJrvKXEsfXzT
YdmjSXhNG7dYGyxFvh800CBkWQD0gQtUpCdykInWPv38ukEMZniJEfsNEZYK+LHe
7SJCoxKLPmkL4hCeqEFShkl0lAeSf5/GHyXVXBvUBfgHQLZVhuelxeNrsPZDlDmU
1wZyRsTxtgCiVPTVl8wY8cVNHfoxA5ULZpPL+AFX6LtVaFMjsWWMHnIpmmo6Khuj
LVFzhn4cmSM3/5KypiupQQDL0LJEcR+OZxzVZdCd7Bv6ecKBRjTALTD12CqXXJY4
mwBvvc/zN4wReOz+2EWy8zo1mpGwd2RSAdj1yYT+iZuQOo7/OtO5meSWXNLgYiRI
mx2VkzCzp25rthnUvDONs1bDPfUpb9JrzPvLojrdGtgU2TPYNVmicnSB/iaa2sEb
nRl931nEfwt7g35AnFRlvCNt7WE48UEyXiaD/AhPIODDeKmPcZfwhZco9baTQLVh
Pd5JJBKSl5Hby7F2kuHy+kPTUyRXIVr2wY9IvrQX3tyeY3YhYHazWvJ9zozN19Yz
NRJ3wzeFr2qnQ1pfj9v6hvRRk3WBC4pT3i/HvoK4dmIsYS5lhfXVSKgNX//8eJ0g
dJUGyuoVmx2QF3FnrVzrz/8dPDdHTzppst88GTbw4nyFe+CpX5Q89OxiYj6OFs2P
UVhCCeh92roWkH3qHKWCg0H8ySijWKoWnuvtA7sIyOs6h4zj7tP9oqYgbBfau6Gp
2OLR97W4QBiGnI/cKdVRr47obv6kw6xL9lKD/WLXDYVbn1frXTf808pAsSXzI9tn
QOS4JAoCIQ5zjke22uFW88YRcqv8SNHugkyQtx+dlhsCYHF5yf8JHCNLjS7cEtOd
6l8gpyO92bvbcVDOHRlCqsKpDUa4OfbrPJBz/e4wTpPasJnkDUWTU0vpap+TmvJA
tKbk5Dk2FwnnxKmx26rpKJDrK7HzkLIS2Kf3Hng+7NnoXJWHtKC1XkltULzq5Sid
rjQrfFLgaiL4X6xA6CCNCqjytZdmrzlSzRZKd7zwC14jG/sFgc4jAdAQ9gHtfUI9
tlbVV6Eac1LNganw8CS/y9nl9HvVanet288zlMFw+GHLgOOg53q6hhDDxUATsz0c
E/z1oN2QPwjoHXXpSbsUtbBD3H/mGn1BleuUOvlFmr0AewOyDNPat7XeI1qUVJYS
s5ENFgz3R6fCRRJEmk+FdCaQFIFU9+lYke/AkM8lATYs6gUZNirBBapDHSHl/t5Z
4X6dGtDVmTgWpYItDjI1akI4w+OUvRYC7TSFM1fiLqt20CazRxWolojAc+nbILxA
3SEVUKwKDzNthpTjfFhIuMoAREvk0grxiKtYGcBmQjP7bPvjFdkgp14aMg7JRSyc
KGTMDq5tvEiBE/lEwhBQ1hQULY0j7oGeBkMClDus2MC8JpS2kC2QBcz+o3JXRG+K
hrvledJ0/08FPJWOeFynxe8BDDsgBsHTtgeYT30FCdc9QQ50HPThvopROg+oOhjL
UlLHqOBU7s1WZ2iwFEr1G+5pPgVaAEeaIw+4KaAYtCYafD8LGhRgjikBLcaCjGyh
VCzHvaGPd3nhSPxeIHpki7ax7ZeQ3zZzT8NjU2HKFJTK7M2pRk8pyRV36UiHXWiD
x23jp1vhjBbOILo762aUUINA2wcAf0780OnpXnC/vJOFqYY0c25+nyTmsJ6uThZz
O+33bxI9UIo915WLZ3JHd5CRwz65SdS9mdYR/1Gnaot7Q7pXVT+LQyqG0PAtknjF
MJQjJmrrDoVaJz6OtYnRQkmp3gV/senNuuyV/97fOpFGoncoA1pgKenBsxa1Cr/D
LUHMn3aqG+nPcCueZ6zQm1+HSSEmazTuJ2kDATvubhaq0KrXWtV0jzGkaJDMw4hg
YetnhY4l/m4JEBkSOdjxgD2c6ur16NDyeAV2ozYQ0fZ4fpum8qOt029xK8SGAHcE
acCOXD0/6eHg7SMd8vWWd7yhvHMLLZkQ24GakWqnEXQ1L65Jc9rG7EMOoulKJPYY
BHdIN4IHhL3OQ+WXkA2+mQvMvKGWTY4ibMnwbROEas/TGRDI3YprwDy2I11Oqofk
8N4gQxfx/B+g3Ifv2j9txfQjGqFB2FHcDRCWu0V8hEH8jBDlwY0vcGnYNYsypP+/
6ekljMFkN2Pxt+c2MyZwh+CtPPotP7PKUl37nk19YjT3bh+5u1FbH80T3n3ZzMmZ
hXGabUqdJ0PHcaYCrgjtAZZUBMTm7AOijW3wAVpufAm87E7ImflBjMy9Ugb0Xm5R
P7AmiWm2J8Jw9xVdziV03IITpfNYfMIf9I09ENixeTwUsRIwTd8bdfBFvD5NjFS2
QtjJ1wjJTh5ZKf4ofdfUmdQIAkiNEt6+LlHLvlbtNVaMQ6ska8I2JzFfC6UIrzQX
MvNsakl5hrC3rDOXpymM1rQC9WybSN+wRATzmvqYDuRiOOdRXey9vyU7ZcRIIgfE
Cuw/f9eSIk3qnoXVnAJcbOz0ZHf+vqLLGDCfHpxif72F9x0nVJobTE1ME0ZUEj0I
/qJC9IWtC3G2yoz0I9htCSBgpEPDhJrnKLJONrM1L/yKnm7YaeOnpT2Weq1ltZ2C
7XY6O0yziaDaegJDgWIsyaHpQRiYm1WZS9ZuWdJBkYFhZQX2haGuDiERounwq9Nu
GdLlfJczAou2x24+kYGBS5zLwpTuVrR90Cc4Hhn+v+1AkFNTNpB5vg3LMuwt2LWU
t7j0aFy+silk8FMgAPbOFwJE7WN8g+xvotMjvZalg3lFc7nWAHibryiI7Np76xoI
1yBk26EhbTCrnWrsA4OS/r690Lik/XkN4lMXuEBdQ+PT0g9vkHn2zBKlMKezbW51
xmdRHD07Ogq/Nf2FYW3S2FUYUov20HxJdulTB2or7eyNKTw6cnnaoWzBNKo2jsfq
Tgq5b9zH6FppEOWsQoaQdnQbsBGhRzJSP8tcVRgWqkWSwxU1nr7CeZzPheqCgHGi
OqFjZ9BEAlaG361kf4QOKkUPFsEjgYbGZNXVf+dHT3wgC+es6TtJl7TvxPh6M7Jm
ffp20NHIZSxi/iATMqDiiGnpgK7Cj/qtJnLY6SinDY/Eitcd3ZMbf+5+odqPaRGn
pm6KM4ldxITmXq3t8KZno/MAFtWhdnlEY8r2oX5VN19s+gNY0RtmNX4L8/R9n/Sc
z1jSzcJUtM1H5gdFY0EmGzxSmp2qFAd3bEzbaCpAnwdv9TKx0/VwpnLDDXpqSf0g
O2sD05WrIacU/CWmnuoVLADBWvqvMkGUJ4EEcZyFbLohL7OBGkYquPOjZbtBeNcn
nJKuvWs5UAn4tY++FuTJkysa2ZV87xDz6k+4r87f0Icu9QWZ2SMVdIxo2NyyFfhc
r3QiS0twOjW1zaBvdQJFnDGvqFMp4oepE+SPGuz9j8MbpuQXVlpeZTOjnoq7i/eX
6ofSRlhjZmyl7HsJnDyvivpCrRUcy14MjFJHkS4SwemjvZu4LJM6kPN0yC/F6wJP
+J+Ohh5nvLNCjLy8qhrazfIBLuJLCqa2vILw+FzngraBdBi9rMi2iGIfAN4Xhr/4
ncOjzp3bLizFcvjm48rt2UrzY7h0pfVkozuDs3PZ04ucBfSrDiOpk1u9pTIiARnu
dRbwm4Kn8G4fbCiOViHigjcsNTSKDPepCYxiyh6I98A6okgWxlqIk4kdQzQXfEbp
pKRo3kxOhp29DRiwmIxVnRsrdGTYyRbfOUlg9+S3xZGTJymax3FXYfAGk24pFGZR
raW8tfTUulzevxTc6ByEHgs5rktsGMjC2v9dgO3evY88/kyBAzZ30dlQvMMWD/R9
IiuelGncm0Wq5TTUaR5ZFT1z4H+ggR21mMDUHRPkofm+iyn0qiVCz4j9HE4tlf97
uygEX4ZLptM7uU8sKZTtM4E0xEg9xcZy+5I86rTnKV6Rz/161Sv1yIAQ/7fqLKC6
hBNYOblk3kn7mWTADT1FlQDjzPw10ukavi0K7bBRPzbtj8VeX7gP1oq4gC3s5B+V
kjlN506ppchYmITs8th9VHgx/iNUqHNgpTI+Y4pUAedNobItnL1/Bs+gAabpUl/6
h0+ubcruXQaxnFKxxxuSY2X4Lso0OJpyyVcULXQZM2QOL+pBTKVecrM3ZvFHOHNs
MuYN9YxsV+NfQuHQAqI3pU9rTgoQtFz3RaNdOvlRHrhsPj2ebeKpCAIDwSAwMggT
gbUWPiWg2K3Of3Q5ZO9mWZOG37J1pK18+jiAjTIqS3FVvUz8lmNDLzU6+3JNw6s/
2ZZidzw0vcPOQdIxQ8oeTeKXV/Ws/qOv3CKpzLYBUI1SkVLVpVHssdX8PMphZO3L
49X+BkcUq9L9bmwegKPZAVhCbF1ZAdlSOFbMETKEJ/NSGNvbukWBXCgCydy0Rrc6
ukxKrFHpcqyDna7kwkYNTxfN7hIT7ifyt9E2V7iXJpDjQYuBzJuAZIhmx9p7jFlk
6ARVkbwFCU8kY5ysHOSPGGOi9xLwMeIoDQJdnMw3iaNndDv47hSlGjC71KvtwHPP
Jdwb50HOY4UPdlkb5YerESYoBtyqvb+nne1Mv+1oBGo4iASL2Pdyn5L/tMJVzEBZ
TOuzpPZUn7ydcSsHOZ9+DUOC3DESvpriBUGFsWK3VgZSLGWVXH3NMgyecSQATNEf
7qHuamJMK3jzvAHsDtHtGihw2QEr9dpazm/j9aDaWMEt305n60pLuNzlNVi8RGY0
AvBPneL1+kJrc0NQJyWA0p+SZZGJ29iVVeqv1biryQcxYLozR89biC3CGOdfvQCw
BfZbYWLDEnPSzwcTZTZUDUVX9TiPJPtPMKVMKR6wEbHwwfv1we3+gJLxVUAyx0j8
dYblnBtCjaNsMo+sVj1aVUVAQTpBNnh+RbwsG3aau8r7XBHwhzvGorqmgaJzNyXn
YfG9Aiu5TBUaEk1HRbDcRNdwiMi5cCWCgkAnUdJdAtfM6w0ztv96knPBe/X3AlTT
UFJ4TlhxkRx1f3mRVfrUYZlbNacqEwTMZ56enGkQXGx1M4/sEzZE/CDrsw2KV4ct
ksBSKkSuF1CtPXDJtoaZJTqGgGThSjumkmbDuFE6goHV26PAGDwET3hUXamEaLZi
mJy2OkOEa26x/6uT3CbICnkLqEYr6+Z3SX3Wwi2K3H/F6B1/S+AEh4z06UpzgK9m
Dj53u/BiH2CurhmFJ3MpTVPac6Re/cpimwkiS4QR5Jp9cfOZF32xiwfqjHgdiESO
3BbZwj4akC4okG5sYMbZItTKIYcqHY1ak7P9A2QTC3x+lCNluweQ0x+6qMPEGF0z
7yDhxvyc3WnvMyDM+ztzCzD4ypxEZNc+LRwoJO7dzbWIZlUuOFQyGBZwMFtRzyh5
vF3QSIZJOI6BGnoo3gR3dsI14C1G/qGWGCK3Zld+M7gjc+xjZs77vo+gh+HXNmjO
Igb/G3VZGTCt5Xtq6AtZKVLBi7ZHQlF7oDGbm3lVqkbKud/H+9B6DFgV2EtMvUce
fKdqfwQExZSy/WBCiVayFMpqUgKKPlT0dbCBaE4U//af8Zfl7gK4vilKhfa+88+M
HD3xvfhqTQFgRr3x2Q+sC3E7qgIEZt9K61UctmpciPqtX8+P5hr7V72hipz4e9Sn
S9p+fn9SH7Wa8YLQURu3bAGHZy+Na4Ps3UwrOIVE5MeGGq2QWE0LPzKb12fMYIfI
Br3btvDKYFVHsiHQxBKDXX6SdkQV1SeaC/RpcIvSMoqsdEALCxJTy0dfSbg+3kuS
/rJ0Qnpw5cr3hDh/MOIa5Rqz75WZrDKRkV0Ix6fFml0urDGeLMUngCOrVvY6iF/L
y9aj+5dbdo/eAitTkUhbzAUJpAZRIL3eG3ZJ9R0d7WosK8x7zDIFzMepLpjPcPuQ
S3u+tgvgh91jpUF0cG5mPWtJ2S8nZ4YqVfwu6AElKDU77RXU5jniraZa5x3JsWvO
q1PS4VcGbTQVEaONtwht5sl5LUm6EuMjhAWW9L256qaGvXWaoQLNSIvAH9teWNlR
BOZIgWzSar3zD0oh+itnTKUk0TZsFyZJ09XU4bNfPM3vIevan/tJPHoW59woF8nx
6XUr5aIpTvPRmNLKNpukU7xt8Xnyncnv9T3WZ49zKegw9h1esARDW2blMADAfSwt
n0AqvRVae3nOiDnF+aMTb+zER1C99+SZCnXj31cvVW4H4wgBi4t0uJfbZxKTThbe
S/bRG+VtPSrXbitaxC25R8U6heerZOCpnSh2f+xzady7beH+ir4fIuz9Jvb7KsZq
2qeGrbdOlFUvccPV6LGiE2JZfr6m0KS0P7dVLV0WtvUPMc/k6oty9wtBg+7FoPXc
sRkG7VtZSI/dR/jlfXs/Q3lkSkA8DulakIKYEJNYI6fv6fBAHxWbfiuT5X1b2MYW
g/lWcvOHgfYWTsiDlL5Zy7MLk+tRjnacByA1KCxvfPvoAJPkzXGbJ2dfTWgUTxA/
+t+9j0FI7A+9wCnk+T+gU8g8ORYSpCmCg03eH01/3DNnHWwBcKYXU4YH2oEqJ3rm
kDbjeljGLOovVttBH5lopIjTBLczn/HEV7W/UDP/VbfUiQ3MhmmeRg4Mk105Wa6j
x77d2q3SxWNd4NO2iSMiduRdzwJthfHp/KaVILwfC8zb4uLNHOmzqPbIQzLOwf1N
ygbZZ1/6oJtSVjHQKh9LqjOyD+bHgxHF4bWRK705nP0gNSE9KpPXzYH/JuuKvpcq
kk5SFQy9dqn8NeZxvlZLRVBmSDphk60lJa2yNX3caLU0mVe9edCoe6Yq6AxhKZLM
+xpfLekfabHudXS70o47lRoGtoanoeJWXz4IAohu00+l8SqnXZzlLwoQNabO2Dmf
djhOoSeuyvXhUorNx7j0jNsnFr+0DtUaKWSrqzuM90ISkC7AO7b3Qm4OTGQpfTTy
LCG+FhunQW90RDOsfBO7TGCBBkftswmS9d2vgFDa2jF+hFlOFUM51MdDfG1pmgrQ
A3EyCTLZEUZRXCiS0dWXj1m38qRA9QnzlKSiZwWFVOOmMVdCyMKhZyTobxRkcwKw
mtGAjjV1m7ptn9FfPad2PLU/inCXQsqazBZS0Dy9Jn16aX/Xk9hOSGKu9Z3MyOyx
fndShU3E26g3xkHMBkuIww+3eaozgvv6MswIK0uQheGXQ3PVsWK5X+V67IDEWwEp
jbpbQvzHe8G6U+zjskXtkR1d4V0O+M8dB6gUZ0pG+DRhspkPvn1y69EtbDo7F16L
n4jnOewtAf8j/GfoBXUpBhaRheuqpT925JcD/Hd/KhxYO2A3YhmFD9i8VFdNILQU
YBi3TP1z9/Go8fvheuHaG2vk07qChTi6eHtp19bmY0u0lGpm3dWWNIBrQBbJkQvw
FW+IKK4iIj8s+SVfdOkV/nNBfX6V485fGYx77J+tjixsEV9ww/NgvWxOrsEkimo0
gOhHN2b8yMEo7e8je3r37g88QCKcOsh5nriBTfhHRBE2xkDWi1oAZ8eZqg3ef6JU
hiXQO/rXJbe+JODVH3uqxzLtj82Sq1fK1vxlygGGjH9uUlhe+wcYpTHnN94RsEgs
vqgHEMjpc63MQMWd6805d+GN741+UjCwi+Yiz1HTkmQjaTttMQJrRra6ZZU1hzeh
28nZYSejwqUVOg00cbMeRMZyMmDSEWPu3X9imx8EOoQZXvjCUtc8Sge3AhuXGMqc
2ZuZHr3/FJluvSIqQ2TsXgUpjYyDu5g4CvLzRsc7IZT2sC4lFgenBMu21lJvxMO3
m5GgNJqXcMKBAv9GaTvdPS3VSLrzxc5j9B2TCsGQdkFEvqPe5aIKLp5vP4ADhtZu
ftKUYHp/sBFwTqGdMSWpMfNFivZaHCvx2v3SeKvdBvo2YERY5NMmBRd5RCqIEYew
ii0+5ygOKXmuHRjZvCOoXTHe6UtOKlf/OvxR8j6gzgHZp1wKVNZiF19ZNLATEcgD
4s7VdI2N4yKjGSOZXnU4dvvCzB7V30GKJQHeqva2N162QTnP6YZg2bdmL+Mvcm6q
NCvXe0LTyoXG6TPTWOjfs4FPJNxRA0xO4wGu+2vIKyxvKRpX3FLNZhekSaA0/Sa0
53c6WoHrAsYfa6vBsfMtkB+CQv3AjmUbZHluC6H9+O++52AqlRNxLVNmMitoxOik
2W60joliqfXXWg2Yuu97CodXG6CWUKCr7w9G9znXD1SeI/NK/xQj558NdyM/AwWi
4eCekj0TvYLTOQLddiZCXtdQLnpvmIDD4btt9gp7IPzg7xkxxxfudic0xjQ+4D8G
C+jOEdgtM8lB8RYwWqEVtp0Z6qveb+qiJWQWOmFF7Q4qP4tBC++CnUe/jOs/MV6P
WohtdqEz7gmz3Spe7WvWzA7MyYQ4tGGUtBRwWlDp5v9NdUQHbTDNpHdtPwtHoM/n
Uwr3IeFDWnKNGRh+Aquut+GLC8ek/K6ixRbkbithxKn8iIHVt0oqk2H1kPwmRwYm
2m6QogvnaaMuBx5asMgpDBEsPazG+xVGpPXXxQK48INchSrSWeOMAGgoOgM6pWh7
7u1sPfMFLQcmwHhDyVF77MfFpftglTw8jTxieFXX9E7+JtWtPcJDzWQAXZ1N3NHh
XL40qv2Dv/z0wJaGdDS1XQzaks2Fn1ECQDTik+5odlIa65M0u+y4YbDH6Z4M59uD
QIdOjvi3HAtuJhkTSpqD/IYTd4gAWbEYpFy5tPFK1w/jB+Y15Xo8O1OeTWs3B6MD
C9oWVy9wU1ffNgSGzxRsBhzjRL08qsFAGneiQm5GUFpzehlCe+tvj99cNWEXuyZJ
uDIyh0TkjIGv/WLOYFuRcYg0Fdon4YZ5KGHWFTJ6EthmaOpE51clxXx1zjccpsEs
7x91if0VQd0cBEZwo2OhiS/A3c92dSh8REoZDt4txPmexRIvt5+PW5E7StELnMAr
21K9HH6IFBiPvbgzcJYtEc1yGcKSUKl221L0M0FZtBSPEVnTIQZuaJb0QJgj/cbo
XeCZgoiN/oHw+D1blZU6va6mSZD7XfIbJ/uj7VnaZJyKm0YFwBWReGLlx2OeMvb/
kdtT2dlpfFKm0C2PPt4C0deIzqX4S6EW0s5L0YeSrLU1UpYVLO2/HWmFlqyxr02t
Z/jmzFm52OTX0umah2y74/Ohq/CRp2vDbuUZZkhtve7y4iSd0A0km0hoaQuougao
eRQI1Ntp7l1AwLazL2MkdvmyB8cloS4a/fhBFXF19TMNYdTLcSZNNC0jp0S/k3JP
fqyPvT3P2T4crDOXHmW+PkuIZ6fRgtKxcDhjUBULeR9eIBIj21OQoHZMyaIq0MmS
N7mgg+9yP92u9JVlVDKOhyIEKYQzMe8MFG/E6rTvVOFSCu2C8OZNHc7sAtsnf4SP
YPyx67kHOXrdxV7ryuR4Y05XVRWosl2/pCaAKiG8u1V701eCl5vvjxtd39/dwXKb
DSov7eqSWq4ueRavmsotNNHTUUCL9aYEt5bh2aXjq1jjlvJVRJgvPmBKMMdF2YKz
N3xaoAXVdOFAAJY+uIUNxDR5UGZsSTLBXqGqrtY4fnuGrGL/BfgPSVDrz83HB+t0
TnOrf+YEP54mlE5oFBWws9GyC46bFKeZDhbUfIzfcKoAN6fwZJtl+s06y2daheel
XetBmFkM7u5jwVHhV6D7l8zreV0K262/4TqWELywGUtH3R+mpmNYO4Zx2I8E5KxJ
tIYZlG2XGf5QqaFSfk2mUJx+NCh4J5vClYIqH59cUoSxqlQUXR7kWi8xO153f9sT
9jpP1UCd4uxtPS6zPCKUM3E5EZhad1/bIh7uXFcVUlOY84H1dviW9s9/pr/y1hyA
rIMQq45nNGlWv5iwfjuwtcX2s2b93G3tsLhvk44zZ4FJVLvXISM8JnAVplMESY6f
LL2jKBDwhSbfaHJrfOgXmZkaDFRiWlSuK8h67Y8CX6Phscy5uT5Khm376C6IX2vV
MNYPtmQXHuL2mfxvEhxdW4drBEhH1CwIUj0O8VmjynEoQDm0tezsBD0R8uMIgCwi
TNoRFsOp7RbE6JuuVOTUgY7m0HlTUMaNvgu6ez1bjW0RumZOza7k0d9Wg5jAkk8u
WmWWg3vzCLVE3WYFiiQIx0uGlb8hMET2CxKHe2AL8mcaIPoWOarN02Cepxbk1pDP
YqNo4gmO8G95r5pBCY6x7+mIYGIUYhYijjNXtNJmWRPJgiDzupvxSM65Y8JB/7Nw
zCE+zugmTVgV8iQNWQp7aiL74xVdn0aOMGQggyv8YTXsM3T/cAo18eCNVrTR1Ucc
x1rqmedIYr/7aiW9vQl4Iwfin8sVktE1amlPVsJifWtWLV0GzOsSo1/bJI0miLjR
+YFieKDA5ownOAkYyrW7YfEHr7CIX3cfryYQNcSDNIXL/+UgF/j1gCKyJBDRr6St
jJFfe5/Z2Z/mqlpvAsUgkg8LHqnfDqRJ86QCinGZccS91V9f+SuBBCBhEB8BtrUX
qCWFXYgjhiyF2lWeZsxUzTYbm+RgQ6BM+5cEXKgkfBJOnUpe1N5l2D3qKgTLmGBf
YLLFX+iy00LTStIeYSJxQxvIApXnsY/1ILXVOGSHAt4B+VjiNmR3LUNuH8d8QypB
UbKmvdqXYTxybsd+tVeR4sk/mlmuCALztOnFj7a2wWL+y34zdQpgPggu6zpWDX2k
fDXu60vKhcpcIaXhQWA17/9VY3nArVTFem/uPEtXBMYXaOgIgu/ed9JVca8+vWXA
VQ9RqrlJA0P1li9/rSzesiMBbXxUN+n7D/dmmCwNYHnEcxMTV910zfgwT2B2Hg9w
8y44SVm2pp7ok2fuAeg1+OIjAXEn3oph9Qhg07xnQQD5kEJfBdkPNYi9zcu9Guqx
Bgcm573/4FCWuSTxmvPqZ1R2NakeoUedbzY2OuBrSqt/JMiTI6+z/jl//4UMCFwY
QK5rMvLAFwDiaYes7GTXMXWN3685U1uR26Mh2yyOc+/tcYWRCG1wrIBGNyPM2ljz
AHCocBvqG308EnlSr8xOhhjj9joH1+hS5pziV8PvSDzQuhB4+lq/DntQo4qglb92
wIsWfyfzrkc5nlKA7nmgxq9jgCDAyEh33e2d90POZU9KiAYWU4AZ6a9MQKuwFSG6
ggp8ktcvrBN6XhJ+TkimqRlXcw52Y8kdrjXzcqCVeYO7EIcHHPu9dDMbY7NMK/iL
ImuRgSPATe2g++uXB34rZJ0SvPTceBfpUTrxpuJRkUNLvXAS1xksHLS81DszJfil
Xy2g7h3MYXoDD9xUOO7nr3HdPf7G285jqxy4FKBE/HyYC1B1tgFlgHz1f1d+dTxD
aP7duZJk5hoFzeKSoxeywmHlwNmT4JH0zulfYwvHonPAZAyEQImylxWmuGiST4/a
zRw3MzCblk6pbfDQxZd5XKqQWclBiMDtyNHw7EKUepPUVv73DcVYgNKw4IilDlzp
dctCQutJ9eCz8GUO/Hp2eDDEToxdEyn7VPDBw6wY6ISxpA6BKclloZwL/4atjfYP
X0uCj1x8YPC2PJfRXb9VWYh/uECdP8ucIeQVgcdKRe9MehD4Vm9QZM97OaOJ9ds1
6tf5AV8jPkyKj3OA8i15KNeTWf2OJT7xfKYoii3nhJKNydt3YpJtK9LiGaFfDHH1
ybBReNnNGMrbAV5iG1zR+tnKELNawbP5fc1i770f/Wum9qMGeBHMa/jJisGPW+jg
Uk0pll9FUwe5JX2soeuD9p3vybPDkY33s25jYF4KuiCs3x2nwB2UBuv7svSGT/Ab
jf5OFev4GPBZWLIAZaxtXAIlMS+LYDpvayZgrlES3hf4qnWcopkmsuA7Si5FkaJx
jd5W6ISDYZS9Sd2zVh/FiOA6nzxUquM0Ye1TtT1sF5iWis8EkIAqZmgCgkM+W7mg
7dNRq9+YeaXkUj76tknKryhGLl8j38XVZsBWG1Km/RV2LaXydUR6JJytJLfebPYK
E9T8pOWnDU3+Y5d058pZNFK030wZz29OgM2fqBFQ0s8NNRAyrzp3iSm1AyPCaqpP
5OiraEYe9XyG+sad0FZdavx6uTL+dGFtPZide1sKroT8q2zagugRaF3AgEP4NLTT
sv74oAq/BKWijhtut7OSBhtjSyrJjz9gYlE5TPZhGs2tgumBs4hNCDkECLWvr3A8
V//+xjeA6at32Fr3RcEJmcbeN11WJks2dAiDRijuV4Aguc2L7Mr1fm5rM5U+ogO4
onYpi/XF5jvbgzxXbCxvwdt820PFvTipv9mslnpjQAMabA6mUpClpRI9EtC5ibRD
PYasQl11JYBIWwfEE5SbPrbThlokSAhgSkxZyTXwjrb4CHxwUlz74KKZPjd3Lz1x
GDGrX1XHr8Al9HlPRfEHP9qL2Enidv7O8i8iZPQdY6BoRiIIrjHUWLls8ADVcRAS
2HrHQSJEVrxmBra2touKMR3osNgFHkHP15Wd3K37NUNwP6yLq+cw8wE9qsdIp1Be
0lnWLaiAjX0VwAIWa0DRcz7HbwZcADgROiLWR8OYGd44MfpRa8YvEUvkSRwdkGYZ
VGMiZiwJrtnbE1cMqR5sEN9U6Y+ZBTIyCGCt9uB/hHY+28+jBqLRaKnwVN5BbHNL
W2KyLqr0gnSC3WsPpsCjgkwoYOgZbCeJQI3DHb4pOkmGltVdCbN0L2ulS1Ntq34e
wQduw7EaDsZ2eh3G2VTdvq+S8KhBIU4u1xQKaj0kM9oN5nkuu81WHcAcWajYZuo7
C6wwaAXoNjmNFwJQV/sAjpkqkv8MqYje8ueZhxSITPPngYoXHcAbPpGou55VMvkW
QED3i1e/TXfgOBFVxC6JxxH5T/w9i8+6je307xpHJURDq5X4eXJaqhE1+Sa8ZntV
IGC3y7ld1qccSNaa6lk8DKef4uKOmCXKcQuseD4Wp2AKH1hpUaqrwtWhnfM8K4U4
ZFx/zWQKCn9vjudcByCgPrl6IuQXHb7kAO6jNm4oZzoEN5VcXVeNK+WJLFNUsq1+
nP2LOzPX7I59qv3Js8aMI+FvgBfkWiPeDSwJda+cnaW1js1W5YNo5dpip/WUo2By
rEGeDLuUj4TUoug08qPCe5X8jptBNnC60/E9SooQzqXnUywWLUjzwMptUcnpy6br
lUsHvA/WMFFl2hqmTdwgFw215jepM0BVgjjOSGOt9Cf3yCJjcOR+aJZUSQTY10ky
l46R9jFg5CB+xa+wWQAUeXRZ+4Qzri4pa3wX+bYvhmb6kKduhkl6t9Pxg17uVyL5
gGYf9aIJaentJT2lQ7sQBdY1fNv8cLgQST5Cq7w/hTGM5oNjstQbE/bWh1SC4BbS
QTNWegUSt0IU+VsodCAA9Qs92t8M3CfFIib74nBHLBt2kLhVcTJ9um8QbnY3aach
FniWL9h5XFrMyH3zMvIyAvGGQf9YG+Zw8kpUuXpoY4/E5UOBpYVewr+WW1+H0dVr
Gg80d8jUTh8dufn93JbbWyiW83Bm0gyNiAOYvrPKBvRIBXaSwrMrUP8lPfsEkYYf
YrzqE8fwT0j+zONvzqjtveJRajmKIfLkNYeUecH2Ne4lkMcRnmKyGdCCpGezzrwK
fdZqrTWbzXfut7lc1cbowLHejXsIxItjQMS3eGEjRN7/uTqfRWOWvU4eOMj/HEPg
ddYbdV+NnJxWDpA8vMUpLMfApWQg7Vtt71NyN29xgQH6dX7e5pSYx6yh2/KH32MT
DtMNm/H9zd2TXK285eTrXFmz8iImxN6fCFkfzvCc0TqouJRvHVUQJBxVzq0MoIYu
8ZCrDqCTF+3AfSsivfKjFi600LOQxptvB6JB3JyatKE=
`protect END_PROTECTED
