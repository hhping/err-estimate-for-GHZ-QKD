`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r1h2FnkKK0ByIJfG3voVgLOOtOBRO7h2xcHMf8OJOHgz5U2OtOvwz2uwuYNcFxtA
F63D9LJifViKu/6Dub6G2ByxyTtrNaZqnlWxJX+Ls7n2rHZ57YNsakqZUWT5untB
b2cDPB5JyVcFSwyYLniGic+ft7TnXF9zz/uRWRRhHbC8SxdkLn0DtMxdKlBlxgvV
d62y+rl4IlVJkkQID/QPWVj6f39PE8lAhfYb8fAIfYDCZyxSvILOdYMtQ1YwPypY
sQgPALTB45gsS+FzrNQxb524wN12J065OMl84HJC/877O3vI+8Jgo2cV/VrevMRr
dUXgMPVufCuJLxQ0cQcoL/wSiUfG/2JJ+IT6HLwjlk/l+OBczoCmK+txVBvGyM0U
GQOmnY4BfxqmCpB3lSOnC087qQHQ0Gvae54TB9CV4/kxQ+td+eNgXUvavPkr9grb
nSZIsL0KvdlJzUYpZbgG8mh8/YZg9eCetFES+ZYInCnQz0tEdPKOpNhkXPcBkPJW
8X4Oq6T2j7FhhZNq8UIsJ4n7eWPRGtj3AqKGQCgLlhQ6xqA+R6rMpMB9w90J4u5V
mbLENV0lJBs4Xes5FbrAG+jowN4FUEcBWmdFpZxCSXADZG+w7QJNsJ/0nVmTWWpS
he3uhL7UT2J1uVbSp5nVme/SW9r0NweC8FUaEFyRuuWOJ4iWN+KR8/oiFpViNJpd
LOsT70wsD5o/hAnv8Xa6x8PtTsK2uTJrbZe7u3LP7xMw/1uc7Z56Qe8vaCQVo0HC
3QcFireJfl+/k/8R8EMB3chsSE51+tl150Cqu7YyUaTr50evB+uUPhsfQmeVcZPH
7WuM0JR5Eoah3DBOI0yv5vY4/ubKH0pO4kQ3u8J+MPFS8HW7mrqQreE4TfCfdaSd
Wh2VBVKDkhuLIMxlmj7H6SqeGQTJKhkZcEAOXZAw2k0ErBOPGZWCeqzbRKud7JlM
Gwyycip7gXDoHvRFMC8PPAlYpDEgIosqhY5XU2fQHkb6XLgvoCzinX/zrtn6KE6+
DLM+RDhzMlybsYVYqDxwlq8eQhgBfWuOx2OejR5DMeq/VpNzvbAIgXV/13NaYMVU
cVXxwPPtd9L/0KPAnhIp85Akmve6OxWRF4n/7yfTpnFbp1HWMlkjKJT4XH8IYjxY
ViHWuIhLLDv9ag6KD9KmCZlQIUQc6fhO2YM5eRpLy3agBlxH7J3AJ2Lp+e/Tw1xZ
blCsYCCM20N1X/HLF+d1DWEfOIdqrlDj9fJbMpGJyn5NlxO9j7G/iz95pDmr+mxt
t3X5C1oaAhUQ5u8PGRKeZ++yd3Og++pEF5A11I/ZP3xyAZDd+Wtsff4y2Lh4wNeB
Hc9rv8107zTMrf2zLJqmqLyqjdzoRKMHMQIINyb/gsoHdRx5tvbI9H2qVPXO53gP
C0/TRJfKpRAc70lKbDppWmFcYCgi0420onGfHgBA9zKEm0smIn03hwhh3F/7UGv3
eTMkyKWbettJ8mx5ZmIacgeryn43S/aet0QZjUthSAeuDDHjjjFMIuFb436XSAcn
px6dNbZ8pbNeV2P7QOD2Dx3PQgtj8WHmLUBffH1NwZ3kNIKTqUQ/e6UlYh/PlAv7
6d/omKjUBnla5g105dD0XD1MjfQcf8dod8uJEZiJf4ueCNe20POInht+JxKdt70w
F2xKS24boR73hCAAA4V8Ddka1Ol99aoE/kMZ808UJ2XlrKIiNo0jiPvb8maROUT7
X+kCgMQK6WYEBRzzstWBVaYxZdLgSOXULU78WE0EcIMLhHQJQL7tmQvL0vSXkf3O
tdMJCb1T94eQ/uf6lBKuMTO7AN3ldbQisOnRtgQf2Hsq3aWONOW6AP2+hOUF8UXI
+rJ2XjHnLqQlnSgQ7W21m+IFkqdC7Sghqj3agdOx4CHwiJuTl4w+LX033whht1W3
+oHAX0hJ/rRimAvVbJyNR5SrjU83eBoAJxIxSdD2vb7CkBrzW8aZ19zN1+fJR40j
CglpJ1ByYb8W2fGVmOqp44LLdTe1ZKOIILgt8eXk2QJbwfzlh6JKgBgi9AQP7wZR
NwN3YDBKcKvv7ZpDIxh9PDer7IknegPOsgL1GQQmV9Ye29BoAFqlcxLJyg3XXkxc
7ul2MAILELWBVRqfczj+Z/1JdDIaEeKpCToA2hq1mwJ/KjwgPDzJ3KkLjpL7BlVe
ucRuPnqk33NmLoHrqi0LjdmQF8V3jnrAyzuIbuqilKx8vmQVD3uMU2Xe014pfyRP
uYEkCqoK6KRZQm64XW4pk5Bs2iviMLllfG2aBgNxG4HwMSEIfoYg6VVXUIBM04R9
5IZGM9LrGFOdT9FsPqCxEAUSfCe24CbRHGNsndirE6p360UG5nGAiglq5vRMYDTE
zJm8JFuXnjjeDLOagavHQM3i1VoZhZCvHzY78zcr5jY2E3QdCyiIfNGBAOZxV5iK
SKFV1RQK8eQM4Yp77gfIu9624FMeonAxG89/F4bagGn4zVSyiqwEwOJYcSF39b57
rYJWFm7T7F1wrHcoY3MyrRUKSEsVdHDnHqFzEEAzcy0lig+BMN/dTMh2g9Sz2LJq
6P0kX0A+ic6JOuQC+2kQ+oeS2wFSlLt79tuO4ATYq3TOB+69JYIrBCfTNpuAIIhU
Jd1xcEcs44M3ge/9bjwDwVfYn3a3kVS2mJf3Jlnxa6tSxYVe36v/3xTnbIsoq+r2
02lnEZADDTy/X5vU6IaLlMtFp6Gy8m2PDDalxhP8leK/wJtI6ASR0S074trHeP1Z
OSwS6ulfGzNeFzg+eg1DuQf6a2VDpdUSCR7VdO6g/kXWOs5yqIf2gL6Tg97YdHP9
76DobUEzlbCVy5W3jC+kqS42+zykB9+uznt5RitROB1w5X1cXaoV2RlGYArDdKf/
p4V6re0a8Bm6A7GJbvTvz6x/GgjnbOS+V4o/vaO6cZ1LIRWnf3lxmemF4dn91J5/
xzhnqPgWX+WthN1r2L1trStJ+9uSSGTUze3yPL7czfr1OYGTCcanYlutdiGyrKou
IfjkBmpS3tGgp33/R3HRLvhwMWtW0Jv/e7plft27LRn6Zx1Ncx+vXfqkmtNNu/Hi
bXE6GKYgP2Nmup53nLmXIuXMKq9cWQbOCToIYInbWUzH7qRbJ2ilGe3VBhAmHCKU
phRotXduUl+Hs2FKswLibeI4CCFWif/pfDQyPM0BOPJiHg55EMFD6W/oV6NK3f0m
HYPqIb1JohmSCwuuE5UnM3K5U3JmNeKZO+YnokzOivsTOx2t9OImmqz7gfUjg+5L
N+pz4yWkGSBBgfMYN8/k+tFrLxFEt6EQhscpjccDc8GwCoKhQZJYVIS0aAUWkNjT
XYEJklOOnuxx4g9DIIUSmUEzRB6DxUXbv0MSNdeDAhAqxcQ0qLSeBR27zPLM30W7
u+PTj4ZnWUf6V4h4eB+Fwtfk1h9yPQHmBLgAfrNPpOLLCCSfDt14AlAYefH67g9I
bgHEi/SevOf6OBj8O5tWI20FNkbV28TAKFxY2A4JRxI5UMvw9hOopa/LBtIQEd2k
Sp9pLTwq0jt9FbqZy6exxy8Vt5He4DHL4fDJO3lOyguEik4hKIhiYsFzoY1vsxB9
JdktvptueZZNyxJle+3K1JgGCdWVpmH0Q9TE2kcw4+tEhFZQ62eqkZBFGxcPqHiB
s+0T9220c29wDHI5x4LX4eCjJx1SUKiaAG9eAcBaLVD53Z7a2TYUoO9R3tgEuTlt
C2z9pxFMF2SzbYz9GUB5r3Y0JK3VAxbzEV344kr7JlymCOAllr7M3UXnzlYHbvk4
pMeJ1hG/TMjbgJ7f0e4iA6XZL/MhFyhYXFcR/hADuOxwz9T7dEEguWgVnmYnXd0+
wawgeOapsV2ZWsa7b14alK5L9gbI3Lj++97/LWV+yOaHqtEtusho8Sew9Hn23A6X
a0grLaayrszuL2jaWaS62t88zulLNmc3om6ZYBYi8MOPJ1O+y5gVc0f/Z8g7L7wT
C6RAQwwrpdRod0D/aNYe681Lbs7cRCmY2s52B4plpGyR8lC/n3qGXvoUHE6pXxfV
+I/Qaeuwbbk45huEnnjQ7REfveDzC+KNgYcW4uG4JJsgBWk/Vqik0FmERRySFBPO
wr28K6R+jI8PsVQ7fCQqCRekeBZ1WyCB2rTfzEDRhThWOXL4GWSRdsbSejclOHNl
ccvfIqFInpUvsJ+M2Cg5MWDDR5GtATf165ZNeS4Ts6VIZORsBZVe2jJ6VZ6sgxkD
bD6RyACLy/zF1dTQ/jmIucb0XnjhRkjamEyvDqZ1O1CeSAw6q+nuvDJau0NUc7rj
TRO6M5g8cujc9Vc/hU5HNj/DmwUBqtufglKjvRFIsHM5Jdz/kGBViDjkQYxnWZpO
NShx74BhpxsVwVoSkkCW5ninIB+zlgjM0OKyXTHC96di7+RmQHsTn22i/6+3mGN1
Om9ymdeu3C7msX6zjV9BOY5R+myOuSiBjyf8P3kBseHBsHAcuroRieqzFRQq8pr1
5yySL51dsenoEpw6KkvGSwuK+msOSaG1SXlPY9NyCYurvmvsniPHgC46JhVxnI+l
RmMt2NDG58ui2jBHZeYSq3TaZSSIz8AfHLAHZMzX13g5VYEDMoL9NWirPiWTDkcQ
x23zByGRSBhMA/AY8Ue6R0N3qx035G63hb1Qs121nJFL9+b+dzXRCLLY6m1/k+Cc
aSt0A/+1vvgzM/iwLZ0FaIadDhtIfk7KaXsXy/zjCeSGgxvqfxIudUd9x/u3ZaMS
ea0I0ymGLFJrx/m/YpW51nQWAzMsdotYN8+B3YTk3tSPP8N3IqsZE1+VR0LS5Iyq
ijDzyxyGzZ865rvpGE+OeFOPUcAmYOxxiE3EcjoNG49fl+x3CK6Wo/Jtk/UquJMf
+kZPWgStkYaJWkbaE8k5V0jnE+sNg7m0VyD2tk8P6lg+I6PJAeYQts1iw8b8Cxt5
PM+K353SIo6ypK1gHBZv9sNUNOlb3GZav0iIch3EQ2yKHYqhm2Shx/YVBTKuIZgr
H0ffwn5WthhRYNci/gueKCgYEz7XkAXVeJUu1ZnTYpQ5fvP8iuF+BQjnPf+BPG6X
hPOc6m8ZhmOC+25eyBTzOijffUej4JL9zzsrKEohv6Wsyx+KMPeeDfs4PDdXiY7/
Pa86rbBJUZleiejjIRB6AZ2rBptU2Pr7CGIBki9jV1lDk7J3XIou12ds+uo35pqw
l21F5UJC88O8WwSYfGcQBY9Af5bKqcAKzexFvFu18IZn8BcI39/wd1cIt9Kcv1ix
nhOkM88a2g1oBhD1PGzWVXGZPUYmV0DIHi9PKw6wm5OukH51/1dsDTFgaymTtShx
bW+8bcUkKdZa5ei7d7aUGhtwysPDx+DjK3e1gccwa3Iv1TQgOA0lANp9nBnQWwzV
pjzIZmx4txz0SwM1+Y7g+0GsiJViAzMU9qH0wEDlBUmLN0i+84K64URx6WsR8KOb
YHW8T1WPTL+y2ROszfQFynhogtoFhvzR2c1Oe9++Vmfzwcxtdw1R3o+pfQl9jXKt
CGPnegqRSmzWQeuGnMI93RRNV+CaFGg5GE1LAMi67IN3CYmqKpJiEb1B/BhNUa+4
eo9bZ6A/lglcPu9PC/vjR3ayXrjE+oDbTaocsk58QoGFSpQF6rcAU6SYxh1fVDT4
wAnUjNbn/m4C0BtXGlFW6Nun709ztzoyW1CjIM/uwspLnRdclamC5edxbuWkj73V
EeOKHC3xk7tMMZgpN2qiOw44Ts4jntGL2oLq+5K14LhSXvszqB6cvRhk+13TjFRd
OxiH5Tyunyi5xsgzXFGDu9SYyBAox1UV0izr4Wc+2wRJ2W2ZSuoJlmwtQ4SVRgLj
jNH9H5Zp0x1meT4wS4t5wcNIipBes7pwfHtC5rZlJRm86j0HFLW/TQj85+87tJpP
Jx/maVDRnrPB/l6oB8xhq9cA1ypwwLpduDOw+EEkmCYgMiuFEnyu16dShrJMfvSr
3Non/sQoZ5MHcXTKV4rZJcbtiwLVcgU6A1uw4KamguC8dGGSnJJv2KuQZgc+j/Fc
d4VqnCbp4dmHiw+3aqI8YzaCLvAGM8xl3ZKgNlnqQBTvtRZrvwgFzVgPG8lN2XXK
3opXrzD86bYX4Zakzno+w/BLFkPJYnCP4wzXVcIMton9DmPy6riRCl/W4URftjvo
R9FmH8mrKOcW25994MvIJCxcwXc1/WhzeSWr+MDfE6PAvzIyUddu3MmRiu9DZHrV
fZno7NnQxnON1wnl5Ty7576IID30KNACfXGQ9RQ8pa5IvuZbeWmMUoUnXhUKDyM7
+r6dZn/IEohQ/xqOTbwMX4L5SBR7Nxqzxsv4g/njbZKb/ENPKvnQJvFmmViXeOT3
bi0ZIO4vMJ/EYMEi4RfvgfJv0i70bw6kOMH0Mh9L2uRnQvuUt0ZHpOUIUM9dK7H3
9zqMcLUwH6aR8Kk5DQBaMh++iyPafWyVQG/TKI+IeT5DvrYWHTMI8kCEJSN3ckfW
A67x4PSe3Hj1oeyEYD9zazERzftS656Y7d+eEbyIZ8KUmVFGcm++POZFtK6TxD5C
AMIFTRWyka9Fo7aJUVw198zKmN6M5jgaebVGoFzMKp2oKXPn9UhLJqCWWU/lKLdt
fjLGpwhgbH4lJTVwC5saTYBFWwbj45JPbTT1zyz46G/nSGfFk04DKOFS+yUMir1R
qikcCYnSfIVWa9H1M/555UKXWUj2yiA+AxxWDEdRmnc+/as+MLtqljVsKm5m8UOH
wwan0YdgiPXA4hPT87WZ57paOkhiB9Xoxcmjk0y50J837fYTwhvLrd4hQhgi7QhH
zSqnONzQM0EnquNfC059nQAe3KiXsgDo+nnlImSEUI6hQ7WdAPikB3sdJX+2tTUE
UnuKtGxizPijw2XIADfNwaUYTvQSYZ9IYQTfJcVQip5/fKoLNM5L3t5Y9ebOhnYB
TT/eJZLS0TDSM0YmaTMLUUOCFBqfmMrotBWHWr4HGPE87cYQVWMMEeSFQR3s2QFN
Xx3mut0W1x6wEf1iyL+QCkpksPGsgQYvqRcaUSDHReTevw814aYliLphiWpBR0g6
uSwrKT6aNwJscinDtYu922k33jnX4FryVV1wLxmDQc/ocXFADqIDQpdc1VmI7bBF
nSVPViwQyvSWtaFq3mz3jdOWMVSGUmmDs6HxTQD+EVntxH7+438n4zl/WJV4BFx1
Qws8ixYVIjKFxCTQHVkPSA+KnbW8spm5ygAMpjM07IQ7u1yBqEo0bK4Odv2I3ZS0
+OfnRjLKfsXQG/Gxl/SOsOTfJBWmzygOdUFUhqf70A8QlA1++OGlFkDwulvW/Y7P
Ut4pgy3HsVCoCseJV7orFioUXMIHo3Nlh9rwWB3z2SD4Y2dUEpQh46kFE9X7sKdF
8zE0eqT8Qre3vRMUShHbu7xOBZND7A8yflebe+qUg/q+qukLHMpG/uHM098AvZBu
X++PDR/1+v8Q6vbg3F38jmhVowWFj8PjpOPlLxP0aKEYETaoCdk+o/Ky1ikyW/9V
zy26iPNycXThVeyxGagKAZzJaFzjak83gb5QluHbVyWutQ7eIhMCbIeVzXFxi0p8
E0RcIO8tiV6CfIxkFnGPzGE3Mj1oJZF0KWrQkz1McZUzQ9IhxfwLod/6mxb6Y0z9
6nqF77WyaAYgbjJcE+qDK3d+UVCDh6DTkbikBq7JIZ1Wn/WsBEqPRvZfRxcpcbVZ
/ROPEocmBX5RToXOMaiZf+7A1/ghiv5w1azDafo6/lqBjuv2FMhaotO7Xh991ntO
X6bHVcfe/XMOA2Jf0Q/LbqgfjrqquKHfBSqjgT4hu3AFcqQRKvrfkftJcMKQmOED
xbP2syN3HFkY5EbMJ5AL+3Qtih9sx4kgnbV/15Bq6Tyi2M1jyp1cuBcTgIKUOtjV
ZT+q3ZhZ6Z13ci+gQTtVQEaYtT75wVwReeOk1B111XNetYH5xFJD7x/yVTvYHmpd
ZZraCr0zprSoLemCVW2DqTBYELgHbJ84OwpgkXYI4+wPvnunF1AOmBykZAU4XVKj
8XY2K9pxBRr2x6HH3eCUUsxNQg9YkZ1nfSEALs6tA+n5D//JfikNrnKq3tYLEkPC
bstnWmW/eoRryb/Zfj0ADr7XIgmjuBMdGMYoB0gguxt9ckABtICPxcfFe8cwyriT
IoiCiwlckrsgr+l6MK1nnqa9Hsg29om9azZE7ZIibiAtIcODrAm0aj9NE9xGNMKd
hDXj4/WlPqIdqZSdsDq8u0LdH364SesLbUOTa7thqI7L58FqkLkAxVmHHICkpIw7
T44LvWNaCC8ERzopSqq3j8DbL2kQvdIKOiwIuBhNo3eIt3mitKpkR/FZgikNVzso
ICoeQZKXwom7fetD0vD64EyQ2A8vTsMWbWuAdGGVO1s5sJoB4RZckxICfOWZKDyt
NN34Sf0o+Guk8wOLnJKIau1kuoRF4hp2azZxwf5l0YkNtT3AFG9Oym4EwpTcr0Fq
Fwykh/BjSRhaxY6X8Kk9SRiokMJir9EjBkWlnzlWb6X5ILqCTKIqvHJL6dS11riN
+JCLayBgcczn3CQs1mAvuV4pAYGAzzV5z49vyYIM0+oPJG0UtHpq5FIEWQ0dzyv3
KQjnBgHnmheejUUMBkXY7MP/nF4ZmixXJJCfRRQpzU+JPozjHIym29xoSzRv63RF
klc7kfcm9L2rCgAfp/wJKCxs+FV4ICH0yyBkKATx0QGNtOfichUjCxn6YS/+PO/e
OJC7jOYdkOanwJxEAuouXsc4FF0XBNE+QONdsdP23kKECkiH4Ef5bALyL6PDa3DZ
AdDE1TxclmWuRmNK0i+dI12/PzySwLjqKURbshIaf2/9KSRAGjbhCCXxERcyYKBL
3xUzuSqxjHVoNSX4GmwEnxe22QhoKlxGHijEv4fSM9FlDpcIBiKyonc32NL5LBtk
u/o5GbqD+Sy98P6Oi9XMmHg5GPZ/zliM8q9WBIQp86leMPmxH2unPupVQYhcczx5
+TdU4uZRUErYVEiGBWG8CMlH7R1LXpwwE95Z1MJWvLblByx1k8QFQBxoan6WNkxA
XhL+cD08zkkEe424cVSybdTaA7HCQfAZZT1oSCrc4cYXxCp1RpPs6XLbyONYwvoH
RKOLbeSbLOXnAQrksmQxMOY3o5vDUcwC9P4Ls9C1s08SgCmHNf8EooLVvMEB8/8w
eezzhs18MktBQfA/42vNC1Iks/AhsheavydCXi/NCZHLaVtKSdkAMp64C1uQWL7b
yOvXMoemSsupKUqzqS2VJZA7gmcYbPj6VOkY9ezTNUVqVjUT2WiBaR/s5GzLBl/B
AIU//dE3cYeURtyM8x1NCRZQZi7fPHbJe72ONqZO3EKWM8Kb+ynlsMGmVXBlXYG8
fG1+vc8VOGcAHl6OqbbzdM5pd76llMIFRmSNkjFWCK6+ooCFg+eC3LESXyaQRqrO
RDcawpRhKZugNxjuheBh7UUZdjv0ab2Uy3TTnepiDlmPzdTRiQGNJbRchSBAA1wD
r8N9SM/uMVxxnECgYHfVp8E9xWXGhT2WD2Gh/Epr04/jb6LpYnQcJ0hRvJZaYZqp
HDf7LU3/kTtph+HOs6xOtfJ2ubNvr+hkIGWvrIOLdpji1gzF1G20uY6s17ATj/em
BZAMFsmX+iVizoBLoOxI2aX8VI/Cbyf71YRSEDF1wX9xF4ZkMQsRHP00g0hkpHlX
kpIb9eZrOv3mlzAekmrw9QFrnvwBQYDBADSZIR/txuhCQKn0y5XzNBP0chK3VMxp
riAV0B9FtPxsjBHgnjanTzvFPgh1xAf/SewQCvCO67wwZoTh87ntsJMVbHMFOsrx
Z6v4duM9sr4EFak4qylHq7CWSqNd+YzIhSFOPGlJrD3oFdSlm7aWM9xBE1rot/at
UtSk3FA+x+A4oIsJG4fIVXX1azsjilFq5A5sEvC7Af5drup4UkvY6CeTxsS4rSXF
Am85f5IHbrW8FGw/WyDQLVySiJBIH7PKRR2b0uGQQ2M59lpJ28DvtAvUAfk5+pmk
hQp5pysT/12/U0frOMKNR+xSpIzuBHWKL4fw8xrMPrCyolSzPQ8gaJqG8wUu3zoH
k/r14rI1yXKnbCZkphVrANXdfUnEFHU40EZf2Wa1IY3BULclevM3TOLlzmGJSo2t
w7G6Ujy8Ejt7mAfoarVWyaLuhF7emTMSeRFytyg5ywwJjlL0kjidwTFHzWHKAu/G
KFn4kiH8NixURJmump5lwBqq9usI7fn+rzTo/PiMfe9EnwrEoeuJtFqnJQe20ZoF
2kxFUYqKZVHkEaYkKT2IVvFrT9Sw/6kdqVCpug1mivMyUp/RAUrIXRRejoXLMrmc
mUDkws24ybVNxMFW6vD0Llsv9Gef1zStYhpF3bswLZg3avQGmzCdItUrtMDGaHo2
D6l3dFcZlHHAxpnzKIfvzY3on6PsA/oK+ernhspGakgiUVVGQwqoyRelRLORwIVV
malsOtqzrSjfajASyj1IHp6AjnVSqwQWdrCw+eyjjNKd3G3ejDWupkyQ2HS87PWb
QTaRXlh4Phx56fIKYgZp1skvKG8BO3JgxA075pQSazOsM7H/dVggKJPYg4uqluFV
gHfFfxFMAO7cTHs1Inltj0xCqjccaXOr9xfy8LOFkHvHZTIKG8Fb+MKfMnmzidkA
V3MGDNkAkh6sPyPft8lKS3uDLLM5J5zBWLwJJfBQlANpg+NIvUvC77gm6pmYA0ww
vpnhDhBuU+WX0s8r9LyNJXitGwWBgEQgGdcDvbeETVQ600nrcbygtC3s9DQ22nNd
9Ma4MkH/GZEv/hCTB5OrjkMDiIvQiZdfuHBFpM3v+k7AKfU3z7Q5g0FhhO4TmqBj
ZfsKySTprNHcRh2F9a07vuXXSCL44Su4TYjKqx6T0Hpj/kSPb8ZN0+4391/pSvhl
xjhmPzlid3xEsP9hOXq5xVNbpcTCzBlPJmGrJnNSV73jAsBjWvIhqsj+P+LfOphv
/YyyA2/0yg3kCa6RF8ipwKKxEhuZq+x71s1cv+5aEqmI5rdJjouypblvxRaPmdam
maNZzoRI8cFWdzS2YkNBPuIIpX5uvappcF4fc9wWOU0bZUMCKBSgIVce+TNhefzW
o1aziaBQcUcbPhxoAM8yVe2uhMLMRnrPbPHWuGF3xdPH262gOMsjc6YjF/wBfHhi
YwkJZJpaFsgox8YuKQmFhdceZjxrHONoLy12qEfteT3wwZzbJhSPM1PT4EYCsJd5
axlLgOm2IxULvpv82T3z+Gsfv2IyBh5AU6bbRkAvxfeTEyc8jXM1Fhm7NFG38Ptf
tq6Ns5pt8xamJz21lngczrVUSNPXer0Kam2Gs+gN4wst4tZkJyiRtzjtWnorzOSI
9DLu3T/lHcb1hKdvT6C6EZzi/g7eHaFYMznLs2GiZ5B4IsikGDR4NwDsi0aaleEP
FGK+ZYGJZeQWV5qYKlAMdne+YahKkCelYDQ0FtO3HYw6xLKRCndCLmnwn7wY3+Ex
Go5m3JU6RJgbfJuZpzzFZUQGgo9FSt/KOITMw1F6/KwZgjmxusG2F9ZbtZ3UaJAR
9+8Y1JCw80vB4j1V1dzyuhTq0tB056yhee505GXqEuQQRHgwRxtDyn536K8rb10X
gvE7PiEx4w7suu5sOnzQ0hE+XNQRARuiEOTXmbjsfjYYSWLJ0Z6AwbyaVN6MySmN
Tz2neeGmowhfzNyhi8ehCZwm35BKgopLdM++fiylgZVVqHkr0XrcYLfcaEZeKlMM
Bsf+tdvNpdC66/0Gu1gumMK0WcVre20UrAgbS61wTVyzYW8ysAnicyd1nccQsaPw
xh6YU7RTHyMGgaBIcrCmPXkLJQZMdoDkTrmSgdUPrHcC1QdSGf3VNjklthZi+T+J
pggtDP+01E1FM9piKA6EzBu/gJJRqdTl0cx1xW/DRWA1/nmvZ2lm9Swg1QTTsZ/U
rO5QyG76+BxesdqYzrYQwax6WpW5bEDwrIN9whfQo6IykgV4L3HRdFDYkZGpgPTF
fb+sqOhHOxgxt5I546/Pe2Jp7WOpXDWufHWiA+TccYqUmlSL8cPazntZIkBfS0S1
On/7SZb5UdHxyrbxxzpCxMkO/2CYzSkIj7L9vB4QV7E0QJ69SiZEYvHD5rTMk5PB
ywtEEK4eztsS4YCYx/8cNtGAc6+zvq3RVIJdxNdNpWCOhiQkC0/xheUo1+Nm9JQP
0OW9CyE0e0S6AoVwE3Q/3Up5X/h9b8h1bJUJgyJvferaXRr/tOL071LwoiWfB19q
HAgiPfN1Nl6AZsc1W+5w6hsBwnl0GYBGF/SW5SXKJ06Pk0bKIxs0lkmjp/VXKXwQ
p67QTIsXyLrhMhnid0WRl/xZTOeFJ2BZFO4CDNj++Pwc045gBCL6QsFfOTHAqq9L
0rsEYkHIXGOKrBq08I2EJH+QofT5vwvDmMXW3md2XvHFdMZHvyWGeOv3GTJKsbJn
rTHg+dX7Tkn7d+DzVoiZyHjA1P57Zm+sPARBzgAHYwOSkQ4sZlVtsPrErO5brsYN
ewtfhgCznUxeO7CNowur98FvfDxHZtxRvlZNXBNGSGy+5GxC7XgRWYfZqMUER4kJ
Al2rLlC9OOsAo+jkcXohpN8cynbrdXVxtDe3z10ZOE6m5g5Y/aZeP5miNGp9QG6O
Yw3PdraED38PIfmKB8ImahJ02cB6q31UpF3YzXrR+z2x8KP0VRjrkTvyD+X+XNUO
vbeRcy+5gzmc2XMgZwvEs59shr1sDFREdsXdhNsTqbiThzW+AwDN6F+aflEAFegv
/3U9l/smqbAhTr8hF9FREGxMYM10Lg94OHphw7GV25O0JFJ1zwTMiXeOYRc7aQ5g
a2+yGkSujh7qgntv1Y83QNBBaWLXCvJCT4v6xqbuF8DaaH5kownoixDcgD2eW1ju
O/lcb2xRc2lAdSiiiIuqHGQbLV26ZKShjXcbIJDWhXCc2iGU2xK7fdxCc1Ks0EN0
E2NUHpRc4uaKk0Fu549g9r2NuaqrV6sosnxu3ovpkcAVCl3bkBkgY9T6Oa4BtW4g
PtuoMWQLiWOV6/uDqEKSN9REwtKqOvMAbqgjshi8U1jMQ3gs2zp/mJPiojhIDiQk
xFO+nnGClTokl50xkNrAtv4jbsXrru24H3SjunCvBySrSZLYd4ey2x4dhlw/uJg2
6Kg7CaT/5W0NpUxbuhPADuW03mJ1wXYOoqzanP6r6VthMw9wuWpdD7HotOZG4vg7
iE86y4E7NRWhfxulSDa77ogxXDPiceSsMenGx/YVCKWDEA81E0qBeAmdM3m1XkGM
oUuaZOLdAOlDrw72vfise5ytDgi8GKkzLZsJN42Jon0NJJMJvjIwc6xjrO03Xkwv
g0GpJfNokMltb1gyNjQ8+ygzVkmUlxCZUqYLxXMcSosKa7+M8pX94AcZk92dZzhB
CKbqmTG68nVEQ7eHC/0S8Eloctuy7ZooVPUthr/5iqR/w+Ml+xwTKQOGEcg3Pk0f
/ubSq7YmljrBuR/tp7/FcR7EfWTokcTXIVXXqTONv10YDzJjavd+noA/Ge3HPM2p
MoXi/bAEMHZvSAhpV1GVgvzEF2ISj4zCrBez2iG4GKWv7ZmciT6EY/X+mW46qCAe
dVjbEJFMcslOWx3xK43SN1bgsux5FnvcwEcuh6xgySC9r3tCN91+YcBiGGtz+JGu
5NGOcgXNRX6G3KBOoNXlEGHzwAbptcp9A3F5MfB20MYhNEPLaBHSP1lOQk3UM/2B
8sMglRCYBt5zUUUDiHiQvzeD6yiEGgbfbkrd1EoLGdzZ1E0Et/GhfH5XTGhWIVjt
+lDvmQAJ5dVFbNrl8xUYI9ge27den+kqLPu0bMGvhSy6NFWBhTeEMCKGjyDGR9fK
uq2tZLTzPJPcQtGE5awNW8oODe8ij9ru9EfDZFGPzhAPQPVxg3wvPBIVQVPTJpdi
rMZSa4iZFNpsiMJzB7apThdVVpQTLGeO5Q49Qsjiwtq3hXbTgKYm0eqsjLi41+F3
d7h8FClxQF6B0LsXaEQy/2PajnYYYmWMGGk8JcTW73fro4yKQNBo38I8B/VX+dtt
9zpOz5bxqSdtPZYMuzi3Fgty5C4KNi84TnlVOA/KARn6ILgOU1pBcQzeNbQlxVz2
KIWNyUETMVWua5AmJQgFNtM3eSZhXrWSF5OiBSs7on6OHEmMwEvEPGzJ2eBRxveR
+LJgsFT0XG9YUSihUq04n4emRtN7pEROPe8lnevGW8Y3e8no30ySUkRNQ9ibQiFl
f73e4MdBBSs1j2NvbfDP9Smczm36quaAhObuk19s4GwLZkVrGWUe7kLDCzt+PqKM
0hK2fNe+USCvv8RmyIInDfHTW/6yMVAeiR1va+b7bztd4Rj1hj7KYE+NfUGOdev7
WwTBu63BvlmzmbJF3HvqYdZiyBU4cNZjZ2T3Riw2QV88duW76+4dTromH/hy+b8f
qgTiyAzwJNkZ5+rz2xCVfqTe59+lFKSYGoY1jlw1wI6GZ/Sw2uv6HE4Aw9P0Fm1H
yxqA46YyoN0LX2F3dkpEs25uPf2p+v6YWT7LzBkr1OYPnB0sWiPvE92QTDV3BgRS
Ide+AW2n9nbFuwSQdI29s0L6Qw7G2ObM8WRkdKSLX4FpjKbOO2jXvATr0vtOkPJP
VKFnBvGBJpdGYF3+WWkJbGnhXcLeRErdpnrFemxsOd/n+D5GTCptv/RWZK+iuQKp
AQLgWoqXQRxnE77gQWyCdlz16jbzVmjzOlyRXltBqnBQSX3uW3eQGFWVZj7Zx/In
pefsLYNGB9yXSrI4HYk9GqEYoTDS6VdQ/Kgqxe7hLZy10pbcZaW+AixvrHlBvF/q
uZd8nXSE51RAK/BkF8SKAhEEsm/JzHZoOsHl+ONrEixl4Zc+qNVfrrt+Ii1AKwQ6
Ep+ci2ksAXgLg7UklGvChh9GVGtJHpM7EW8p7p/m15qLKqvHkK7x2EG5FxuVNQ0a
5ezGB//c6zVnaGs7lvgH2gCl/ZS6/irMnMEPWFIJzRqdgfI4tGfA1l9/zrRMjZpJ
d09OBCVt40AMSm6WDZ+RL3+qM5XMjF8+eqmBaUcO+ig2lrf4JKeauFMoQHBhCNE4
mrvNnTqHI6gUVP6dwHIT0npGpu2ZHYWSIGl0OsmYGbFhNf06JMAXP4WyvqoZsqA6
IFv2V3N5nfjKCNeOavDb96ChvJAsljRp4r9QfnWg8oGqlJS+q9mpy/y4HVj9ZJNc
digLU5e+Z2vkaCxx24BtrrvSHMcr+E+oU+t4JrbxMDqW1Ti1AwoliLuNYo7vtXRU
kTHngWqrW2OyCR/G3YyVi6hoY+YgFyz/f1YAorIfwKNrAa8VSt3T8ViWwVsRvtcF
/P1jzZloBoiNVtMFDwScWtYpyuir3HrtGxzXjIwXxFF5CmDoI8xQTDoisDSe0pm+
Mo5g9ofsVbHjrfYPYDCJiimnphjnxhtZoPGvZlUuOTB6TLigMYbT4eEqQv+AZFNC
zDCRlKsTYus3QmPYmZZVmrMf/lMpKI+ShCqgGuUtQR8+V+Qa+6xjHOaxWlmCUoFq
aJSiFIlfJGN74tCUCzn6PD7e7t5XIiLZGqtRa0eOUDJ2g5JXJ8pB2YB3a7jxxnTF
9XGNS1Nki4oTyL4XJxZS6lwzgTE0ObIlXV48fYc6kzbFMCk+JbFjeCT37rSe8O4T
S6WscvDkfYlUk4DfyziDUyw1BobjG7YTegeLsQ1NyUmj/nS0Y4hWu8lBflDWUXqL
TDe05NII5RvoycjFUvMingg1orwhOqRQtK2/C8PpdJbcdlGeulZ9f3PQTagx7q4B
O1AaK/EuSkEhQUJ/1z067U0W16SPcFk4kOelXFKV6Gr/jxzUy2fbZfNiWg/sB1cC
DTvuayGND/ROXldZ1pp34XYs0IkUFRCDisZkNZwm/yLBQxbY2kEuO6eGeg5GIVHH
pK1v4ueHtQG1IcXsfhu1UNoRZID991iHSmJ0kotZ4EtCwHAJCH73TZPelN6trGMa
9Lw3hmCcKBmDuwm9BQeULbxykQOhWBplRAJauU2EePdyjL+CNbPxJ0ig6ZKKPQf6
nXL7R4sNfBD7pLWhu17g4CgbgZx5PgIJFuUj3fOnLnrLmDeYAq2Q7SubGbmZAGZN
uoeHNlhRXTLjSuICQrcyIbhAkcv8yBaq3Ax8EyC7dFNhMY+qrjxUO2AnURjSQeIU
vtvNBu3znwPffoDzl5BDborCMMWxS3CC2VQTEbxcET11X+jvWBPB3F5F2SIENZls
kgOafT6HK3G1UM2sdZv1mlzIQC/UbqXASuS7sKeg/i/4TuFXieVRoRbdSeHGxB71
pY+Kk6KtPGE9aAoIeee/eWgdY9BfC2DCKuXskokSQ9yEG9Ncvnk8OhCVMcuNbQqm
R1hJam79ingwv+pFOA4O/IH5T/W471VHFbzxR5wdexjKQeMgAtWFtm8gOEwh03cX
YCi81+9Lsw9Slk8DgApcZ6i+uss3fs2EViisRUns5ChwnKXHvAN4o5+jH3nyj4el
oeS98uK1b+hL4y2TCLWqIlWf4+dN9zk4QgRRCq8PtTT9b+DVWyvXQPvPb7xhOB81
Hty7HuUcu9w88cOYXycLt/4LWdNJ6NQFgKMuZwpMEbmbxaZxfh4pxXZok57tqFXg
48aghvOVnX+r9vCnHC2WsDl9w7vUOXnDR94+OoZE5CbVKTAzJQPRmQfh44VvBeRz
JIILiut0XktTUJqtBjylhAesuCbRgzcKOy3MJGAGtw2fnnmXKkuAGo4ifHaryZRC
N0w0LcwkC9KMqf1816LDSRnL3WnNJxUw84X/K23tTGnV3NgIzKCSwHybwhnM0sMQ
7JDbTsYYiEPGKjC3zov3JEGcPSHj1iguCK1CmyuW1iQSGI9dkMYQjXfNOQ5AsxFR
pqvhR2+/PHpfb6Qisr2P/inAOmeeHM4YJnH66wxwisk+QOGxJ1IU581k8ypd7SYf
jxZJZauz8nEAowPpi/RGDmkC5SuJdZkRJloFfaaYsYcDcHPVbG+xTAiO2WZyVgtE
dcvwgthBZzeMLNk+v01D9aq++DWFyVgzkIIEwwCS9zQHDIOFiygceMjNz5unLCul
Npxynm2BsG1leMjssp2/fK3xd6hl70p13e57AijCLf+Ivkd3+vrnwmbScqS38ftQ
MnSnsmyRMqp7/8YilHoGKWXvIclMAF/zOz/G8oexBa9spqbtRHSH23aiEp1WbxMG
NAxQVmVtvwMrLqQUeF4cNuC/sCnMlqII6jt6yBYxYjlD0nFzHCrkhdyJoDOnrdYw
gXUWvUFzqnVheqDzn6bMHjiCYimcPzGTD0HQ3xQkMHxg4GBBIsbEjaXypliF5HZF
iR40gxBWoXFrgXY9ZH7/OGA7FGRt5e53GW6IxZEQPVp/OsZ7KMAmo9PkFhV+5Hf2
yod2rjG+47kmF/Yy+EnrTIY0ErDag30uAB65+IyxTUr7dqBfbp5H0zwrce04PVae
FMwkIxkNfPKvtqrhsjVUJLtklBZLctC7nrDrOOOywiK9FC/E0km6hP7PuOorwPbP
V3drNl7M+Ak6UiNd2UVqyTHXMkpmTtlpCcNxd9Mgo4OIk0y1hdaR2ki2byCnbyjL
PVNjGVmz285GMezZZOA62sHnPqfPhlZ7VfMd3x2QsD6NxEYE87YGEDRK9nhKLJ3i
0ciB502vSvRbyHusAiboKEiDnUtHQSikRLNS+bfdR11UGPE8bRJURSRkmMMDqJHi
TfcGZUIv6aU9GXHuXhO+4A5V3kvWhV1fglFyXaltkfSW9uUWl6Hv55MUCFwlFPR1
rw8jmBiObt5xQLgazXVgO0cFrSihr9hxI8eDNIP8Ayuve4Hhjz4X22+2tm6eLaOB
JPhW1TcZGP18PB02kKRUxOlHpB7xa57yfmj0vaBi38MjTyt/jUjwIz09Y6kiZkCt
tZFuktMociGQKr5bsYlgtgz2ifLCy1ocCIPRoBZSHQGwak2oTDDf6xOw069xmBTs
5hVfm1gDtdMwXXywZcmveW7ijzOdNxTZeKr7JxD7IodY+dNViUiFFQ72R1K50dLo
leJ2T5ZaZkRh3fMAM93NPtLbLJkIj0qKQIV1w8/SKw5UOc8Kwyd2RKmxWBgqazFG
eSq53B9KSa86NbYkmLP/SPCeBSzD82jkJY3W9MXGBPFzGq2Ae8ZzvH13H+z2U9la
igw+UMvdRFqaGYd/1cjZS9DeObfYErOd1Nuicb19Q/kdxnYFAM4uxhuQyJBuBqTl
5u4Xe6ze8ZiA61Y+aBVwU6W0dYuM54NUpID1pZB1YakrjrTMjf0JnfmrQQ5ZxWRe
4rsglPjZhf5rIqgdpDWF9ELHZHaxybBFdiFM2QuCkOzyzUfTnB9pdWnb929nsibD
/JefO7I0P4O4826xwi3T+c5uJ7aH1Ue/JImlagLObm2E+iMz/Q+qE6kec9DK4I/d
Y39cNARfPjpZ3NnTEzzm7Wpbs0Xq5aX3fAPVQN/8Z91ZTDHIPC08c18vmfwmE77W
uSGFNd9qHT5m3NWaTRtLAZGbQwZPIWO08IFCvYB3eoIHcMlz8or2MjFvP9ySIlGN
AK2K0KfmQIi5sT+JbOkhA/dciTYqFTyLRY/6NUcIxi1CLcsmP2ekKJuUjhom8n6/
vC0McpDuK6F7FpdPVX4LkcHHUk2vp9+D3sTA2CAgPNs+FNtXpkYGENtLe7WM94Wd
N1lyImAUQ744kf8cwB/Uf0/8CdhtkiCSJvRsg5PuPEPX8HyaHGmwx2dt3FcGh4d0
bS4j4Za6Y28lOdQfJdf57YUcHXE6zJaohNYfC5vtvigfDEpbPg0bjg00FkfS0ui9
SLlVUWbBhioT23CY2RouN4xwyioBI8RuoZsKrloZc/yAC+6QS2Y6zPUq++f5FvU8
WvrmHv+U6uCLQgAtpkBdm04TDG4G7YGVm/Nupe/RcxIPwUmrk+1R/vh8YSFAMnLd
+4Fy+buXRZrkLF1kg1RJqQ6AfVvdtCSIMGxenvRXy7MCIxfngTAdBQM1MHCCyPyS
mcwummKddmWdiXtmbK3ymwg5l+GPIuLEk7ysaP54HxuyzBblosGcIC4jy23cezgW
78lbY8PVguB7tKe/M4lfdkZqeP89C/pjeV4E/Wzw21VzwfFmaVvxHG5EFc2AAgc1
kIeAFOTesH74VFLmPITiUTJaS4mv6v+4AYb45sLzGcMQkj/41T0BTkmzxh8tAvAr
RLmzJ8ODajYBDadP/HnlXQs5bjTLu+wh3/RtWrm24lNoQlI5useljtrbhDMqPGDs
4H6WPEMlrsrX9a8vLKk5mgG3Fu1Hg7PYs2bwcjCyPnsSiPgTdYTNTAM2pvv9gQAa
zm4LAvION2dYiLxaUl0yRDPFk1fPNj9g4JBkC1d5fER5YZyd1DDsMV8XrJT8wAf5
hO7yGN/z5vA2HGdkHl+bzjmxi+wm8syNfdYNqho2QwSk2Bp0M4H+3cPVELD4XaAs
LvBQDvsU1u42l/RAw1GyywItALisd6e/9NANnxSInkgr81ksJIyHw+59ceoDPHxU
AV8uU/NctVbexpGqQu52Shm/lHUUz8KuRII8XnRvdGJtg7syTYYf86V3faVAogqu
pLjd8FiX2PykZcENHlHWQRHB67+kJUNBz9mclQ7kMNWf4WrbGyMW4mpHlzsclazF
ovK9N9uaHhn3PUXOz0XQcksS29/hYAbFy9MiFgeSzbQ4y1yqyqUXKXiPwQ8zonZy
cmB2eHwo/oYBpkWVVu8pm+y231g7ozOrs9upHRoHmxS/VKrx8bNj1aJKfp8VwK7Q
8JHKcqyAJGpHm7PjE/lp6KLOJamuMzB1eTyro41c3GuP6MwMC+wa08Lbf9rc0RfF
ZzhrQBJ22Mw1va7FJe07e6jnVkgGOGBjE2k0ADNL8aVp2PMsfgvdctYqeY7+c8IY
4JJP/ZbT3qLJ18UQfXLkcQs+YU1w/jgAxNsiLqgTwcqkykEmUjoB6EEUtqupQxBo
U5fvLmzgEFU5MiLKXSs5HuT5IHvNxoxTMvW/f2KUUNh/MC6ZCez/KcE0ClRke3Lb
TP3ODCUQUtWsOwEpFallI39MC1mrv4wBia3S722rw/czoZOfR4LsU44K4tvQ/D1C
jvz1t5lWVMt+QfPevaq9tQS4mvnABUEx0pBKA9CIlEhSg89SxT5lxja30GA8Dnz1
qtKq3+8If6IEzkO3H49yBIMZDgNyg0zrFhk74nSdUIXV9z+xsPNcyFLZe4JKT1jR
kbeKZfs8h4z2NrEb0HaqX7ISIuiqJJyj+b4EOQRgyGFFw7jiX74/SkUHWy3T0SDw
MU42U8DL1dIsG6lJSpDDx04vJBofwMb4GKRIr9JCYa66+M2atqBGeradZtOa+sKG
fHyHcE74VmJJ4gFrvkdJ7QVdYqosrULtXZzOWQXh4bL1fxmfOCNuQInb9U0pxZlj
jEsjvRCJ4HVJeZ+1+xIOpsfcWgIHCJlqa+o4QYuELjtQC0pA2h4uyGu79EpfUe26
4Gz9h903UNYZwkxa43BPnvvu0xIJnmTFqhrVZHg5wSRZz/dgRNkm6k3HiuUn6Em1
a4u/ecCS4XcwyRGq6MMnfTBy2S1sFREwbvnL0L8lN4PqLau/VrXYpb0xF1k1OyuC
D2yCDAOO2rNN0eBVtrqEoS8JfhZf+Twi+oBqUnVAAsC3uh0zpfOKXGWBzSTsLDsr
H/pAu2h8qmhlyBJie99OeyqFLf2Q0G2y9nggb9LPunZpbjJdnSk7zVJGbHo3dUhN
wRo+/koQz4vlxK5PGbQbXfBjufadf+wpELyLjBIB2OgKf3FJAla1A2mupOmAUAYo
1XG+QtmFa4FUgfeucpP3M6XiYW5clr0qGvsa4mtFyg3Z2RcE2lxHBeEzlH+VU5Gp
AZPdzzFPNRNEfCpjyvtT+uM2YgGl1WLi69osA1t8qfbN1TQnY4CVlR1mewL6F/lu
HtYUmraD9HeBCe/dJHAgsia0fxTKha4SmGI4bbyLeQZmGDdY02JmKHk5WYIgrKmo
Uwvfn7N05wfJmniX0PLtYNvBzls/mpVxZ5yluYGmPxBWuz9iVjk0u8p7YkMRsh+z
r0zIZvWPY8rquFh7iypOaW4Aub2w4pARx2MB9iGvFQfJGYc0eG4vHwa55mbuxJd3
hTJ1AfuCGlpgfQP9f/3fwO20f4LQ3eRiUad0R+8nuxqm+hkKuxazI54Gk9yYtKbZ
Z73c7yD+Owcj7MT/5fJ/GCxO6TZeIyIulTtkAc8RZv/qDUjt2sSV8z9hW9yKD0q8
J4FWkbAED+2hGXpiNDaFfZ0TUORD1h6hhsicElS1Hfr/buIi6v47ZBMUTu1AteqB
an3aZtVM2BIEa2owwkSbNbK/oof5DXNQb0qXR/YO2UKdsZazBngqIyFccQLG2+4G
6b5ur3aPG0fjS3n5gR/UGivWzEfr5p26ZOnJ8KL8OIfIoYRBqOYUPvlm003L9lnk
qnKWqGkgjBw+MnU3jFMnGmPh8VPU199Brm6HVzWjH3m2TidlXZ+57ZOOrIP55YKU
YGqrxd/9w9Mp3AA3M4pTpYWmck20F44Wx5c9bEjPCUiHRK/icLJYegBm8OYLINaD
3yu0Dnw2U3rVy1bWfk5SMzmwl+6vvA0JOnMs8Ghpu1r58fVy7mhCEZI9iVi9Pzki
Z8PoCkAlRTj+QcQji9IUqxMntf7zYhn6Suqx1sFZ7T0zaCGx0+bjWaAipDjPIe+k
WMeM6+dALJv40702p1yU0871NFgwvc6oCkTW8IpMTpd1lQGbIqzqp7CK5dXWi8Xp
Q5zfsI4TYuk2oSKtu914sr0FC6ckLwXSJYeNpUExwSy1rAO9Fa7QTNw1+isl1Ao2
sKVKMviKlgAu+UIodrIktplbf9PvG/8qvCZQ62+JOM0F6nCHBLApe9ZVId47exPw
TbP70WEo1IuXja0EKZrAj/bS/61aiLvzfvhXj7z7CaImKmLqjB+0ZL/4bElx+NbF
UMw29db4ZEc37sR8Gk+iEcKcv3quVVwJErQvPYLZ3b1yvGh4nsMcrL5JC0ZsiZZ7
kn5xn+xY+IzTkJknQgq3QMI97MmVNAHgWubOSMf1IeWDDl9GGWhDGVQzF2ZUEK8j
mMDXSoXZXxjC/TE/S6PxpQYLX3GGgwylMKHwpOg7hLE4faF36UJTd1mXywGk0NUh
X5CgMy3B2F1iQ1yX03Vge9SGIruCrgD9g6r4hvwEKi98TAFDbdNz1JDfrLN3pHCZ
6sBitrQh5I58NA2tu0TgYKdWfyaeMXulcFOmuroYH3u2pSp3J66Xdvuxj+KoWlLN
qFURjGfXk3/TXUYoM7DHd0MnrVWOc5V8SKwhnzgTv8sQELmw1cLNk2TrW2s/NN68
AVs3o7iKClUj6B2LzXiO/vRKqBvdWTZ6U688w6XXwUwKQ9Ga0zpQa6CLqZ/sNvN/
XCrf/UN9siYlz0h82brZIL4JAo1AjMS6U6DzOklgLj6SamcWkOYXWbUf5QQOV2t2
P42i0qVDVh3Ez1uBrhYu9JGeMbk0KXi3hjKDW70RQu7ItIRVPQGlhVb4K1OZjhKt
b+Jb3Q2UUYxAwB4PbWW1Dp5pR0LIJOb9BwEBiX6M2M+vkg1gjgRdbUMttEMumqWX
zPcAB5aXEVzLOit2GI4Trx/df/KlQz4uRoAa55CoG/kRPsh2HTWE4hYNfIaacfG4
mCsj3hJXNx7SVtCcB2cpo+TP6Zo8T56MLIVyTzrs6MJ7OLodjmAoWVa/uvhAPuE6
XYJTsagiyeAFhZzrOWdyOg7ingLqga3g6qQqdDbb5Y7Lpmkw4iZv29zwlw5Lp4AJ
JDN8CqhA5HTSboW9TtMlk9HKQi6/XUtmB8TlgOw9kdsgEExOSQNf8v65z7SCNFz8
wlnpemchP4W79KPtNkMfiENkry8x+apFkAO6/Qbs1MHhoyX7O4cm3AKu6+aPJZkp
c0PLldy7cQEr2SzuQgDsLMHu7UB8HCuBeHqaPBoOoZw0rTTpDN3PwcGrG94J4Sv+
Ru2wKxBXZiUJnFRHx+qKTRRYy6e/3/9rOPpLSK4RWwy2JSjqzSuS31DN6GObsmPt
arxBjTqkaDvPilYng7QA+WRHZez34a3zb6m1sOe8TT3GNd6sNfvj9JqtDX3J/7Q9
BRkxAHOjXi8D2xVTKZFL42F0qYFz/TSl/MSawRyp5Ih6gI6e39Wdwf7ZiXZqkmRT
lDNQ4PDGHhWOgLChBboN5gDaJuHFc9pznZwpSMMkXS7Ib1mACFOhcbog+CLQS+rD
W2CKdfs7jZzLo9xnvdyGCsUU1e7zo2mD46xqfqTSVJM9afMk2We8znfTQTFxklia
IgtP+cUC/PfxZXWAZWkEAT45CpPdkVhVmTaDko3Nt/MalUUR1tZVhhf7Dkxxf/lb
7WaKZzcVPXtdeClrSK6R+MDPzXuY+LHhMkwJMYUOUjjmioQgsFJYZs9gcLgudKAY
VIVOnvzHI8IdJVCml5NtLQGmTqfe5qOX/jmCCRRyfiuHrCi9j5+SEfjliV/Cyp54
cyqhhHMx+pYbgDEpPWUJqUCe+lU6GeknTfQM72PmNuFXd2SjtiUfofSpjyTPqPXb
5kY1ZIOqLq0vx3BBHU3xGa4bcZdHQN135Yn3P/eMsHo19YdfXsRwB2/2BNpHFXvQ
M6OAXktdppTQtjsrCMD1p0IhEGdLvXf7/W8iTBTMIjayy92mUMref8FxLbSlju3K
LWIlogqwBgCd+3SzNagmYqIsznSJs5EXcWJfL7nipeJthXThQS+NQR3b7980n7KS
MpK2I+v3xBQB8Gx/kIca2uEyqNy1kmw/nxzBd9lrqX6w60x6zAgq0BrDvD1nQ2hx
rpV3l3ST3RkuWyhskqK9p+rP/OCIp/eC7677aqIbaX+DptKUz2Pd67rbJ2/8BmBM
TF/OL6ElORTBP2L4sU+XmKSeXi7fPM0EKYQ/EbJCUgoF2y2tBMDR2BMujjtm3Y/G
6yiVJh8xegy1eDUPeDtCZiNlra0cWhcWvdnBRIceRZ2AYZZWqFB94JcUYAffBGIg
1vGmMGLW8VMX9jr7T20Eb4YrjQOssIHsStHZzrEXO8PhylQZK3EsnxmqJXdZhjWO
8Cey9wrvrxylt1m/7GDkTzrIjFUzXEHKGamGZvV8ZpYyVNFNGZvMaOqxD4WftBlC
Ql7EPrlvYsoa8ex90bTLZHrHpbBB5Z2rWVkn7Mng7ehi8pjh1YuPXEtQhBaUo5t4
hO2D4DHrm3UfK596NSRelXfJtYqm4HujrRqplkfF1/k3s/pNyPuWP+bnZ0xG2Z8T
YBDXy75gXGYewzC0lCGypSIsXunN95UCeynCs9nLLT6CnLPv0KzhieJxX3h38X2v
EiNbJjnVPyXb0H3bCEPSo67Jd0EhuDxcjBU292nDfE/gDnyM9UkuHnS1APg1mRcp
GNU3pYqbaT55eTHmQGSuHuZ2N5/8yxukxJGFPfI97iCLHpctdu3n4+duj0B0RYkH
XOnEc5e9PRoXXgoYgPlgxeXj24A93i+xYkDmOQm7iEndu1E6WpFjFbwNyuooLOdy
xrL3XAfOp1s/FSct3A18TR3QQnqNZwadq6rCYKi7rNwKQuRDt6pgeyWCCissjuoj
OjXCY8pj6S8PN23CL2X4bHnAYlQLzW7gLmkjQxKX5GNvrMBeRtl00WcUbyRSoixD
OTMN9W6upIwYoafQQrX29F4EtTSmR9VbySkkWN2HHltGvOQOdalo5N8gBt+jYbB5
RzCEgZCinOm7Nw31J2JzFX4FZvssFt3fh9GkU4xiyQPLI+P6rZFKETE1ouEWDJJB
MuwmR0uMNNGf3QKJ9lexzJucK6OSbl0Xw9jwNO3gv0RtEwAU4mz4l5GqxQ6Bi5cw
Ojt/brRMM+qZoo8UD6TbpdkicP96EAZWSBHXrdz6eqk94mk5LFSqQUOPaUfWd2fz
6BFg7yC/KSd0J1BYOxgEHLtkK8yj95PrxjE2YB5UjINeXHeatqa6lGTT2wSqTbbV
m/CZ4LZNDbTSfV3w8jZjY21Jn0UTADgmrvvN6UVYA7ebtsh8FIKXacWPft1Fwo31
cuBcxndkEcCt2U2Q6EkhTtgb2LVLjO0yE/Sk7kgEMGfkxjowKPDAwt9TE6gfD/kU
kHirRbLfnoxdjq/5oSQnHiiWr+f8iPsbRIdJ/FRsmTFiriC39gI5yolrDnSuUkDW
6bJLMrVJyAgT2KUB537G+ycuD4du9EHMubd+y/BDpp3rS80iGj/6V8F63CRKLCxY
Q6h5pxJfiK301hyeN607dUw16mqA15sKaTcqqc0nWaPuxsewAseTRQjPQpOC2bUv
/CJgV3lb5Lzof4MX7uvIyuRHg0HZ6XqQPGvD2/94EeMN4Dk0VXyLD+SNGxx4PRO1
Lkbsyfy+kBXUDUqHLzyFspfT942fsq8Exp8HaHXmnXtbS9NGce40VsrVozXMSzAB
4/cdSbdIiNPCEBkiS0Ea6aRoUy1rpqmGjrG6/ctrrYyPgmQKYO5wuc1dI82G/MKH
bnwFgP7SlDefwEUU8wndWmkQu0iwAh5UtBai5JmqNjxKrz7xJDr3R2J7Pnsz/fT4
FKjaTXwOA1i6cs3eqAjRzenK2tmVV2tQtJZggxXttaOFUlkf74mttH5JrMuMMVPI
wYT9iUsEH4nlhDENX5JSENwj+GJMnrrQYVI3OfAwFmupndek9TUJ3OQ4cV8qTfu+
+RtGkLOPWEx/fvyd93jFkyKXjNQyY75nCCskcz97O6dzBZ5C3JLA+H+EYkncHTko
6VhCfjdevyceJgKl/kUW75Cuf4fsjQrU1gt06LAODMIRVBHGsfA28ForNMKqSiH6
7Hyh0Dvs+bvo+YEb1jcD24PJjb89Zr/+ikm+Xu3WZFeh+mKWG+vpYm9YiUJGmItN
TNwa2SiiUOhOuLskI9YvoaX9KSlvmunMrroHcw2CoZEEvXP6YQkEVcbXYIG/7oTu
Ikx/lgIaA1LfB3UZAjpeRlFsKAbyZR1lSVhWBslL0uvfuLnf1KxMR7o/+1a3O9/X
VwGh652fqqBNTZdPgQD9Y+3mqsxmkROfZecWH0nAqDUznqqzLkBlROF8IevXewPX
Cv3MrR76Q8fdMc2YTvGgdQo4ddNQ7QbgxExUZqYRjzyQHT7PRtsP1scNO1RdaQAR
kAzGlhKkoHFUDutJtasslI7YynriJMkWTvi7TyXZchMzbSwd+FeXvim+Mx3aGZyi
f/oFczLnkHte/+dwjt1HHq8mNi+ofBYMLNZsAhLxKjpzmoBIsMo5pq53w2bzumSf
J4Wo/shkhJrxUEohKOAVLWn3Rzq/SanUpIkDG55hoNL2mt/V2CFvlTrlHEa2OWBo
Uq+50/EXrihBwHKxmeN6n5iryRN+9JXyeXVFVTtn4E9yXBcqwpd9mkTCoG1IPNz/
xXmNj4bOz70IHuyxb6KlsCjBKr3FVDDyjLxFpMmXKOYWaRF+616sVLg8i+CxSuOL
SysDg/0AeOWhqOQ1J/rm0FOd0LPecw4EcO0bza1HXWn0Zmnfuj+KPNk77rTaougt
dj2BcGDE6vXwxxFIwGYUOxII4nQBVtUuqtMosSPtA+LyPZEUJ2ecrYRbxcu5iicN
gpXagGuc9NESg4A3vvQzIr+G5S6pptijV/ueiboQs07MUPhCGjOeXKR92/y6wgI6
4bRYV10Ka5jUH80BIUbGG3EOxXf6TxKX3Ndr3W/a2GtF842O1n+hV+1h3OwZ7vtY
oRno+9xDAKyHAa8x7IjsB74LElcvd74imP7VzxKV4VUszLwsnWxJDf9NEIz4z21g
K0IIOQ08wjaQfnRKIgSPv4cqHnSSgmPsfS5xSQ/RXB4RxmuFfwGQffO/oRJhzgSB
gty95AGeTALz7KgT5Z/tT2TxlebkLjy6nOXr3TjrhrbyCqJ9Oxzuh07I+p9o85FS
FF2Wa8U5vAygeMXmJishtQBCg3eCXON7F4cit56+4JCscs+A9Ud1WjR3+vzscGZG
VpxSVJnFQb7Xg9G197qTyc0xfWwYwcRUJXhy5tyA227qOmdkMqnkTgwsOUiQu/sh
9Nh2EyMbsZQstNpciukLNAiNerqeeABWpjzF9YLkNApnt99FTRsxZbCyMFsn7w1c
xeC57s92Z4Iba+E63rG1Tvi0xjP0p8GYxQGAS1pZDHSVgY4OIaTCiwFCXENObMH7
nRYtBzxq9+RllFNVw8jkVXk6fRwrGgS0iDqSoTHGExaTkdkdny+V57DVS2+hzMYo
LAIw789RTFwnbV9kmzPGfo2tbAC71GHAaGECdivFZz9EMKL9YDgLDK1vN/Wh8Tid
4W/lOOZ+cdj0mwxGLaZORpB46hA24u2rGDP8cDD58J+/lsI+IYQ40uIK4Xbii4b4
zerTC1DQKDTfYQRmKGd4bOEIWCyJw6L26y98Uvb6OY6zlC60R6i7lb2UE+swKD/f
46gcPC/RV+hyQg4NBGjEpMqOiqftjo0ZGMbsDdirftyK4SvN0sjGzxWWjtnWCgUk
bJuUYGgH6PJoo7+On17yvoBW7QxoldIaTChPDzcnOWAHbE9qIt3IbgKAA8xyDWP6
9/0foCyfVa0lhjXfgpXJicci/0gQq44q6uKXvb8hNAiVk3Rp//We//vlnGlfcKjo
PcUTfM5alIiChmIRYX5IddRzEJFBWLMpKiDKz3z67EFlQKRl0B76GbpEePsCce5H
w0rFZJTcxIXsCJt5b0hfNpcG/Dmj9fuEiJcgewApsX/1QorVl81iv+pL7MoH53tO
I9tcODrtVAaWTRtdo9NID+M37w06DGsPEYzxy3iFqdByGbRv/fARR1NJjjfLyl4b
YU/kADMHv08LC3AkmL2N/CFNLbadVKyYArJFm0PvObqCWU4qBwHCIflrXVCSnWno
PuKZ1eZpS0soJm94y8e91ASBMZyhJZuzSAL0MYhIaEk1anJ0Svu3r/hpTbOmAv8r
il4XHFUVFU4M1o0EwrcGkmFlMF1TS0HopAEgilI7Wip9aJVk0U/9p0kRFhuDqzXs
ceNSUqg5AbrppDSqpoFrii5hEOammwy/BcYokk28AqePwj/i+BP8sh4/dRE2S19Q
JAe2Y7DcSxwM+bc71SWK+NZ22qFwyUubpYZcTUNBK2VuBt2DSl4H29ZyWgsJgz8U
/f/vR0/fBuEP7QD+GpQNYhGEgwUcScz5t3Z2YbgPq6QpcJmx8MimeiZQUSSEIIYM
ct+vffUR72kt7b3vfAA8dI3hpjI4aQtZn71XMV1Ai3GqSZgRQG/XPPnK2zD+g3LH
tSu9v2b1kYx3MnFe+1ypprwfgKX3zoHfzpX0TrxeWFpJrB6WmY6Rw2ahh6+n8ImK
V9Lh1Y0QVdluwc4tX0lfSyxNCPMYNfX/L1HTBm6K9slRIVS+6S/Fr80rouyTheuL
5tHq9wTpwTDPCgSjSti+dYRZrBgDlSv6+BU7FGX64kX+6f85x/JziUK4drj/1zUR
ax0u8ul/tz+oGcMT2EAUu/u0CRHNcCbOXaaVjHDdv511uwsBm5MTRmOcN2mRUpfl
GxBUiGa8mKjGdM/hSye0Ed79Jz3YRY7R78nNY3jd10a5azoZ1mAvsjah9spPKrqQ
qVd0n0nWRf55YUqg4gHV/S/EW6gyaXT9JA0NXFsCgPzQT+XQtvU8kfJBhy5LwZVT
0fSB03TF+UFtH5gGDThNghPJdNUdtjHWUJ8AnHeEENuiZqicX8J6ZnCDvCvySxNM
zTEJjlbnGFAbcv8TtXVc9uqNrl0Krf6ACAixbdDUmwNeKfzVGYtcBgaOJ8YxkE3B
YHnOmX1SKKWDv95Ut/BLW4U1Tlrd0QmnRetNs8tuZuqaU5jui4NYW1jNZW4VqNsh
Ssxv91qXTyZDUGSCEMkGCfw3sHg+/V5yuajp0FIzA5qMK6qKMImOOoWBjg7vP7Fg
zk+cz5Kz9gUTP1c+J/WrgM1EnQZwwSzeKeyCDLrnVHVgZkAdgsEek4n+AYR87MjM
JtMXus/acKOtOfTS19YwwmmOIRXsLiJXn+/QCwMkqkImgmEV4FuvDTmgCXYaQipP
Oh46tibeB4FF4mIXosemtXkaQ9KOfl65RMRTuhRHVX3IURqjW449yVCOSHVdRMOR
Tr0qqgeYBH7K8XJ6pXrGpmyL2BkgDsB5kVdu+T4Ms1DIOs1DbW+pTFqe3oaogJON
XubdkSta1cwFWlGvz12kSMc4G4+D+wd17w6wYawnWY137ZQz603NtrBwG1ZQfC9p
tOYWhiWqCBzqkcEmOFO81T9NoD767rE+7J2GdndurdgooedE9GP7RhE4NKSOVoz1
7zV3aoH11/8op179RkyA42CMybD8fMH/EqWGRyzYtXydYEzKhmteDmCQxJ3T3OEB
f+lsB2sMfU3jYXoi1xIH5p5U3LWdJuZcTxij1q359SScjjhbZKkepJTA+0r4n1n0
qc6bdvJHyuDuix+W/wGlWVc0ldbOgqKXh2DnVSQCWjyCCNr4NvM/+fBBZXfF/kSl
3QCYt83ya9EQfKz3K6PukVLryfQLHoLCAhxPB5jemEA4BPsCt3MkyjvaoZVsN5AS
eOkydnS2pFD4Nvl9k+BUsnX91jlIQsoHX3Cjb8A6UqwOjNS30MsfDirwJ4FRtRSY
jVNtCnjaVdH8a7DvHz4cdLLxQ6KoZ+0axDTK9xFb92ctzr5GayOZ7zSBWVWOVylo
0aXSBlUmlk5ncVBf13ceJ9wTn7xnMzOoHL1d1EGpIOG89Bk6SOF5m9vDAjtA2uZK
mZWNR3rc6nsHMd5RypW//YlJEqIsZBpxlB+HXDtHJETycHSW2k+t8ud2nJHdAv4h
3mBVcABrA9l5iaj5+YKs52Z/x02djXdsbkDK40fKhazhppFsvorxx0q4nua+lhbA
H1+TMPnwJrgsYt9pX3N00xabYfGCtIdGdASOz+/7J8P0zS0V+NejvCI4Yv+XeCMI
HUBuSRx7EmH7JIkrMX2EUsIyFmMyZy2YaSu9ruqP8BBcHb2mHsDZvdPCbeRaPAtX
AoK2cvzsiZLedhQPMFtbvO+VApYKKdaoXvnZmEWe+edSf+Q519TQWWncfs6f5QD0
+LsbKfrFyagvMv/U7q2rn8oCW/cdMO0CO4LpDQAwSvpNUxCHwm6X4dt3tgmK33yb
Hm7aIQfReDo9pOUN7CMWQAsuwm0QvW7rARnMLZEbKkSYOMChXlmjZgT053NzI9oX
+XiJc4RvzsJesuwTAw5beSWX0SOK7Ku6s17DNPQPKUTT+MwyErdRW+ggZJ3bfrd/
Cx3jCmq2Se8XWb9/+9oIwPmDditAcvIKppcBCatGjZXb6phZxoKvJoJH8OetDLMI
PW2t+fGSa7AXCG8AEs3u1oWGu7+JXD1YYXgTPmBXx6A8qiyTGTW2JkT6i4zMBzIC
NTuFxbd8SDbKSL5/jGmKBPX9mvTvfz9oBd5ymfQgUBKunJqr8RSwUBxg+JeEH7rw
+I5aOjr8WgBEEKTPcN8znBWygpjB+pzc/GlKDyZFYBMo5Z9jscCO0/HUQN32Q5ne
vhJddAwdVUKuStl9ZWr6birEcXuFJCCGeCrvIphM7swSr8sVba50kNMHZjvYF+xl
w6qR+3oEQki3v4P47Rmiqc7gXD8UOIkrG/s7z7XZpVqvENSLMNZB0HYEVgMQYnnE
sFjbqoq1OoKnWlB5iHmVbEheUwQZ9qRnkfAg2/jmmzA/fG5Ekr8D0v2OpZfX6r/C
zKfZJdxZcOvi1oqZF9qMve30xmv0OnTXRqv3sW64qe4GZlkoMUfACB/PVt7KMUwl
fGIQS7fKK1PUp8EECGZ4EAmLGDj70fbeZbwc9s8sttud/EN9wiDL8p+EnNMPCFFX
/EUKFfsXZoiE7VlugqFxe7OsJhw12QrBSG+YqPcOQad4RLi6kDKDvSxMNwr/GM/q
++0yQBz5HqywJ4Fh8SBr7L98qy8DhWyrDHBVyeRNHERGVX3crgZsw9SNFfGwFl4P
e5CTs7TpGpgB55eL2ADdB5pldI/hQvyMHg2svu5nNprd925Zg5zAv1lHtiK5y4X2
2VW8GW8tshUNOSQvDiUnr/q4x9xz55PQY4UkEmd5QgNAm6UI7tykUQUfm3z0NkcH
b1Wm+NJf9ghfoW5KZs9XAe+HxMONtySa7sI5JJ1camKGHNn7s+K+6KLW1go8U7Uh
Zc9M74gm55xpyjU3kST1StmBL//hFtvMRkxz4QgIkFNO+e/n2XWBK875Su/NwpeT
uyXsfh6aYlN/2uzUh2bQwRZA5bFJlWSJxaHJQQIlGr1JVoqWATOqkHBeM0+nudCS
PUY6TnPTIk5fZDvWh/Nhea55t5UtaDxAqfHDOavYTBnEHcu0fnBz0kBcKKtd1F4j
Pm07okqiu780rD1oCsfGhnE1FRniqTerxhyWVnRMdCWkCzi2acPlSCeE9JSAqPqj
4gKTvEhAzGC+lc6NDgQmUScglGYHORn9jL7fGMWAlHnkzmwZ7VsMM+PeefBypSCp
Z2BnmDpNYKoaSTwndZ+JiglyeDvh1o5dPUlpD8lPUtbowNsWZQZIOYJIh5DsPp3T
eblXndQwIKdmICkEw9ubEXKgcxFYRB7UKvI5ZKF09nx5RRcQvtnTb/gEB4ylouIz
2SUU1lnOLpZFeYQ/bQxigpnaTrw6RFSFvStZoQ1H2iLrxkSSwUtLafKCmYIDzmd3
YDtdFU9whrplaFncyasygOCcLvk3LJZxKIvC8pIT9nx24twgiQBF2GEHQrTBfa7B
8ySzHKuv+9Jqsbccl8rpkCTW5naMjmaT1j/Xfk875/j/ixBFAzFoX9EuQezTIOTk
gvM/4l8zWZSmLCHL7PF6XuDxC+a25Y13dgFxYvp9EwQ5wMN768T3baxMGGicp9a/
bHaTiBkPr5Dr2Capy/vD+pIm/GvTbX0etkY/yf5t6wKwUkItH0xHs8hryS/Szahn
C8dFmLgu/uARrL9swFHvlKjYeLaRGFrGOBZB7cM4W2d9Sz01tuoUN8kRjyBIb0MN
JTMQ8FMxaPLQGGdy9n9WantlGFsyRdtCIeWDBGCpB8bXy9X576TFNKSk2Slnx6xa
aM15Xgp5LLWqtaGGkhmsnK0MzzGFjmkxLnd9FIdgU3wgdR8NXx1E4IBsbffQmVaW
lgfZdhIWE3bCODZBEdKviuei3UTMWa7MMqTdXuTqpvC7Wu/YnmZ7rbkM8wlRhNwM
6WKFWu5cA1IQ95whLwBtGerk3sHMCCnv1YjXEc/LXSkeiiOFBYbtxdimzz9CGeTF
cujfVHGsboKDL6nKRKAW67kRE9d9VyeAkoii8bklUM6WUpcDEKpp0xdp1rKPwfHl
xeyq69rRKC6vweE3BKiaIUuzkJ45JCiGvyNnDeGscAmwtqWuv2dc4CFpOpERgLF5
LqejGyjfne588LvU4eMz+QmK7ktR1ZqkOh59P5PIkw/GLF8Wtk8o/dlvnGkP03/f
2GcvLL2D9oUmRrw/MgmQLoTRg47UASwToQzlYKwXf5lKi7NqkUirssnOxqiH6nSF
tPXr5wk/5xu9qRbEDJOBJW2G9jmnCpLxsnzC+zHmH7VZ+H0LwaC0hmaXkNF3fBfY
nCKG3+79wkp6PC6iEtZuyjpHanuceWNae6LxPZl1A4Lh7QRokGXmdoFHomzDdPNn
xaHFQoEDNtH6XipBLLpO9we2UMrtrxFYadxR2FyT4MScNx0vFbnP963rueET1/Op
9Szj8h3+/cfZwcrahkD0YmkaHFalBGvYX7YlKyAr6jem5H5zCWtzfebve9IxQi8C
86ABARKWRbvN1jeyzjnNqR9iTSvem5em6ltFydJCMc66CZVEXm5TWhRbD6o5ngJV
7w02VlQdFEKIyYFd6F10kQN0laNwLhyP5BYI1jXhnzAA/M3ltsxMxPoJNMBDmmYh
anF512mSSgBbUGzCAYFVLA9VZ8/vibnGRUFB8Jgdasm5F7ky2WYiIUcUobyZJJuC
16QnN01BZAsycd5X/MypWJNWBCnFrgdETMkavaizMuZrLBUxOyQUntycdNY37UDH
xNpiqdw2Ak24ElnLu8sdgjJNlruZ16n8hHjDD7v46dAOHuT9qoCfX4LnGxlfmpIf
nV6yLxQnSlmY4y6PJOwt9dgJjYafgTg7HX6uUOFvcSj0b42kElCtmnyhv1g5Irat
BjzkkyLvpx/nlpbgLljgH5NmilhhICqdVe1xgJZwFvRV4ofu7NtQ+Ff7/3tLShqN
SO3LsUHQphFdbwYboy5G/EsnAZmYftPTTKsZbXUnobvURMiRAhHQ/LVWyAdYTBFP
uKHKfhO/Z4wrHphP5MKCHW1TkeLgWVFDVifQ80TLTDmiwWJD2HLM8qpkOYimbNEu
5mAgv1GcopHS09+LPs0BX2TeeF2TNsCEbBWGmXOD4HwOYJVUHFEVlF1Gi4ZVuPr3
FzQ0+5tARVY29LZv0NcOr5j1gTwEpuXccioCf7n15tSRFNmCANU2toQ+pDUrSqPY
6HeSBjEdYTadVBo8/2lf7tTTHmb31J5uGzdorHnihJtUakCPvPhvYBLPoiJe9FJ/
FQRVp6xqmiaGG6UDHTfuR78xH0vrPSx+Jzburo8j4oWwnvN26egyi+DiwMZC1XKt
2W+Z8O78+pobB9a5OzyMr8E6it25jVb1QN4E3YBduxJCerzJEkDm3IEUKX/pXLgC
+ifS0zq/2FpyEZw4re+TJKnd0cuDmH5QoNZqDX6qld2SB1krBy/P42F3sZvTfhch
rSPLUkhLtl3tVz80Gv5ONS1J2wl/ZeNYZOWlfJkw6LLHi99YjePrHUEyVtm70Sz7
3XO0B3ITJd1PuS+XhUEC2Cz3NQc3+bYTMtXszUsOrJmwsFLZvJyVjeVjGNbvAA+9
MFGCd8R9e50DgEiknWwx5+5oVhVeh5JavoH2ob0Gj2M1g7PW6cryG6RugovMb7it
ZlfUUo0LUSsO/gNQWCG9E5/MfY+XXYOuJiBc0NOoZiGwAzMEkUulLRnJyWBtltJD
27Kc82UKGgKhTW2YNlxtqHVPBYIUPkaY1RT3d4b2ymb6slGYeG6WrGE0sjI6JErw
++V26ggoLdlfTFscAarJWwBPvXyPKBRELVFFffS/KIWW/xuVaZ4Jsv8lmqV0NeBx
AIvthgQujwxZnQ799xsnuXD8qA2iPHD1ENNrtj6xw4Dwt0GUSQdHXjm9P/ntt5On
H+ea0x1U5R/cQSsBo3IIbOimCokuNE32HZzka1/d//JPnKja5M54/a/5U9pC7OWr
UMxtFSviDuYnQF3JXV5L4IZ0MnAous6V9xTFUXoJwJ0+aYNsh6DiCSSfPuebRkrO
AG3+pJvDLqiA4JSAl43jJcu1iXa4iHSbzW3beC0v5hFu0QM4gkb6YcBexviH5olu
JJgUiHrCBrI1Ww/03c2wk9WcO9hc5Cy3pUz5+LdA0pv/oj4jscXa4dSRJt3N/Bf2
+vXEYjmrw1soS8lbyQ23Imo8Pr5C0JbYz277kw9cRjUlTCkX2jcv8G+4qpu+HIKq
GJcete3MTCQ7C+sO1PcfbRfW0zF1XnKsYUNFUO5n0KNpGYRKx2TAYgxHvbvhajhz
DaNRXbFsyWuSZseKeL7iRKkqtqSV44E+GQf5U8VuY14gAIvzV/N7vhR6MU8II0O2
ct1oxZgHGiQ6AXHWZ3f9K7leWA2EXJ0P3nIGo2A4yxWv+H2bzpRD6PBH2ohgYI68
xTDC1Ze5lKujkyUi/9llHUdMinylOeRWsSkISfHtFxTaA1HARr5WrIhGpaAbPYx5
z6FXFTqHtqxIHts5qWK45uD9QWTDebEGu1t3dYCcA6i+7vrV2AiHzhgKQ1Z9Bjjb
c0YD0jCpe/MB56BTb2cdEEUe1cSVmEys4ljkBwKUPuZnB2ZpGUijiQM8cEWriTKF
srikuwsA2GGqrI3g66Rnb3m+c+cyKcFTSbDi5qsPt2rn55CswK26HfD6cjFa1USo
QogK6dnL0OET/FwLdy0FVwjq9OsMxaUbKY97rIy3QONpYClUsZRib5u1dJOTWnRN
qJZ2hkLUxncPP2q+U7hL03OyVg/HOiI61j0+GpSGihj8y3E4hKhgZcBV1GF9kX5P
6GWIGjBul2CDz3SLN7YhFEIYCaTeJwsyVzK3hY2mzqYH0SptdiR1pcoIjDu+TE48
aAx/MGvXjEzfL7ECyXHsbx0Ki+UyzAYPgpBCbeTzFjRciGuEsbSbjOV3RLXKOSqW
n5O+ES4S4BkPryCbCoIqDCHUMD9QVqZaLYKKTbWHkqvBPudLU6Lf1AJ5jhRgFYwF
pNj1Op1LTueJxaofeL5q+BCSWHKDkLuydLI9ZSt24umm6r4xp6CUkYN1SbW4UbW0
LTqKvYGBdSWUylzX3caFX43tJOFg5sAy0z9H3z+w9J0SOlVIy1wD+MxNuJf72Va0
C3btG3fYrj7QvK3XB1IMy7HbOPz+akOggs9hC5dobHz/Y/lWEgdFXMibtC/gWuXh
Jr0ee/GpTFcghtCN/6/ve605r043+0EPgzyXqL9gCz9Z2xqUWyX4InbDqh/dBxcc
Rd9ZJz/ZOnUPrUutwJ7hEY6lZU8If+hX7QsrCDiKybwbHSZLV4ol4Llg0yv8yn61
v5LuuqHSwM2Msonj9HZadsMqp2xacWVL8tm2SeYcfjrGAxIfVBDZN4y3lbi4Azat
Wm6dj7zoNc+WwsjWngov86Hwp6cld5/tTkfrS800d+ImF+jhBwlIr2DEEwxs+VBi
FgUYZZ81P1/SX4hZW79A0kY1jX67QcSznVfi9A9KKvPpKwUFL6W7+Rm4cK3WltXu
8UkWdHhSG7m2xRq983aT5WXWl5JoSXJPqaEAgzRhBYf7+UjWzNDOD+EOstXloudO
ZvEUcnmVy8Tp5aY6eQs4bkkhA1CgeSaVhhF/7Z/W2jfqB5Wd74xfwy//ux7jFgi2
cuWAId8lxMpxecam0Kf4DLmfrZe6g7zltK+bJQLicKz6EUBacYxUTZKfppdTqZ3G
zEhoTyL/GaEFpvKDXr8PRBusk/FgpesYfP5GSCSNw+p409czY/djluP4Ulx35c+9
peRgmzRGOG3FWiF+GPoqDyT9WyjUAY8ZTxqzaBDk/j2qxxRzrE4xA1aK9ZoOXW0L
/hnAt+fiNuzCNdHvjwnS7wfu+WleFPSV9y55WuP4oplhkuyd2X/BbiqzZNHNPDHN
X5wnCKVVsNkmqWyoegNmvYgrs2LJNoGPdDi21c8xdz/+NOVCwN/RQ+q7QLF0+sZ/
JOyn8vjCJ2oThfgms3MNEZi2XGr0fQbJX4wi9mW7VURXxrFWjbMUrF3q6PGMYTS5
oUQxSAgf5AgxcslWGYhkP5JnTW0Bogtr8++kHkLRIZQ12GflYrvI3aXYPxyY8dad
/6nOsGbahMIj/vLa4hzBnnXIQ/5ArogQQ818mUKHG5AQZ75KF6cvMbs+Up/xGyYT
1RVb8j2iZ1p9rIFh92lQYjFBvqR4R9CHeKv9yyZu5tGlHf/CHsSEKF0CHRzZIlMo
1ncDGB3vxDdx9asQejFSCLAHl3oVxVV2oLvl9XS2iRbDwYYbbDSZ78vBkmpdB+SV
a1DtjFeIurZelTv7VkBJEOxyCmU9IjCVQKJ5Thx2/+W3+P2g1kvdwaxHk3/078Xd
1+ZEeYOVWTK3P3La1hUmqgn7jylw8/iKIrJd8Fw8D3gRVJKkrstVVF5VYGloAEnA
RF9V10zNpJBF5hwvrVcFkExdfWLK1I/J0half6qKSOzYYnyVRmTc/gVCP/5bQ19K
cCJUNADppvxXHR8wXs773jwCW42jbnikse3E03IG71RABCIztui7Wmeoddx5KDHm
3j3CXJk7aH7mZwLDSw7BJo9Ju6L06N8IaFic8ky7ZM+Ca9e6NLORTMRrXJKwz6Vo
NQBAsC+b7wSyJVn1azCMe46EqU5jQtpNMdNC/I+jx/b+M7VX8iJ5yYM7JA6eweuC
RcS08Tk/Tcjtu1sKhsQvuNHRpAS1QfMysf1HftfDAAx1fq/ImSvRNfwin2BClBBc
PGp90c0y//FX+bYUV0UjxbNP5ez9pZi/RAvkK+1QpEoUbPbutNzwra2oPt5xQaAR
O/SMsorYSLEbQu7qx1Nhro9gaFhFN4lZu+Ik2Xu/L4NWonPx21Kv6jNHg1lSVNAQ
L1Kr9brcAMBxrypLWsS3cf3eZ5ZkOmYSPlTptwLJhglQoVFJ0C6TFrlopsP3WkLh
O8S/FviKs/EeZgCS+cahsT+1hoIZ0DRcH0aauu4bUETxr15cKMMaTF/nz8+gsGby
pVm9ZCJa/65ypjptwYwBIg34OPsZcS4qdq6LF9Cb9IG+9IU3RNcXXruAQOxKJ8Tm
DzSwVeqP9z17tjhRDOm/ouS5FzByfUqLtNx2wZpDgCW+VZQTqRFwSOdETrrD5pml
NSwP5E3kEdQ8cEd7uiUf62Zz/8UGACtDoCKmzHp4sLgQiFhjS70W9faMjxdqHM+Z
xIoBADXsBsBWiFewgmmJEuy7VnLUYSfuTrvc4MMiLlaztNhIo3htbq6ru5WmBtDD
OLq4bofslkSTdRN8e4PVu3Hi0Ixgpmjd7ZQ6dh16Y6s5kGIn6r1jsTWlcFsNrjfW
mdy3hYSlyQV6OEGpciuHAn9BTNJ/PlF9zEBFd7KOYukwcS/4pWMpVFnZk7V/Rlhy
x3Bos/ci55xl7ciAgex8NwLp7j7IcGeIDTTYe4MK7OIA+YOrpqLuFBiemCyb9gXa
oqqfDn9u1EHJM0/VopQ+zUmLZvH9qU0MB5opsDfBXsa2zr+vG65wiCI6Kud30naz
dOvOtA1hrHQMjzEPSQYin+INyfKKVEfYnYWEZ1/kPY8ES11bM2AOphQlB2TOF3DI
rlsXM8Xvi+AIwEEXcfW9J79ScAfH/IgThcOjHhZZHttUsVZKUNxHb0aIFvyGFdCx
wTv1GQADSiX9Bd7a7sYT5C9OXTXhgEHbBDBiUiuPfE3cnDz23KmZZRtDYKJLTR++
jHPw9JttHnOgH26S+Yf50e0Yk+FJptxzpcRkBkzI7KWgnRIODpmg1PVWFDd5ZkWU
7crKo9ch+Yh2vZrnnlWgjWqZhQ+EaTBbp34D2ZqAjF/hOpqlSLhKt0Vd4UrEwAP1
uQfwSgs6ao2qB1YEcnA6bJMdI/Iwh7neldjx17irHNYIBr/1MI5flCf7E0OoWsr6
P+/3ZvyUKUqd6NkFX9UwNM/4qvWTUUvviiTC2kpxiPNZ2Zn9g4XK+X3NT9fnDqPb
lRMv5KpBCSYnE49qTzdIa2QnMVHtJ+WE5ejp0w6rMYTMuPRwlfAlX4m/wpUmZsI6
T+zdlrG63CBLQcw4LHQ/KhqidqeAIokBF4gpd8zmLOVwQbiiKY1T5qAAIhZx60jg
yHiG9UHKu53URzQz+5Dh6oUPczwYGGczf1kA8aS9b8iSE6sr01lvkGx8fgbMamk/
QSHDmXsXSz7zQvjf5rhTQ+rJhsr/FpvJe+pquwa4HMxkpM2J6lLUc0XGMecHA9oJ
dmFvBez6cPgN26IyFGaDG1bgFn4bBQprqzixNyc6aU3xh3nSzqhUG3xeOaGGGBRw
WDYbV9uciGseNmACgF+ja8jUNYWbhhn382etVoLCdD3f/YZuVWYo35sFB2QLjqhY
+EZda7r+hhpRKvbtvXeXYEDUI4YPTEF9XZEkLaWr2niz0dWeOBQ+OobKosK5M/ro
7QF8d3mZomc36bQP5nXgngqkb3e7NdDKdfjW4Zn6nPWWh0zF+rEsaOW0IhpGyyUM
xeUSVwunudUXrodKuDXCtM54byPAnRN/HHUfIXWBouUHxUHBZGwbMmz3RCsQdIq/
V9Uw2x/z8z6A5q3pQ9rErrkSArpYptAXFspfU0TRk5AEdMqscEI3JhGOzWbijtTX
6onjBe6f5iOfRjpte0SuF40LHKs3aQC4u4Li8SrmVNHJ2q/mJgC4wABr8cAhD82d
SME0xEUOlhnoUCzSDhIPhb8Ps5VK21LFrLpJd3B1HhJtPlnIhcXq/JNECbJuWWet
daHu6Giff/CN6CqkgzEhS9KjNzhJu7JJIdV9XBSN25D1nCOcRQmcCaK252owP/ec
g1OumSevMjTm2OEBknJGy3Pue2mRcBpWIuewDayICicNh+JjImWU5uSFb1zTrf7Y
9vMcXLAoy07uzisnzJnIapFY6P1xo7nR7jDbDlyxGMF7rUySvKZmECICdH0G6F6B
plDejYQYi00Rrt3O+S0jNUf3P2ahf4lT9+pOzilNBU5EVhl7A7tgiaG3xA5MRu5m
/3N7GczzogDPc5oCofyRtLcNyghghzrMOshqg9yVRd0CzQSoI6u+006gFEeiy0F0
EaArTzQpiJQX6mCkKSZDhEofd2rGblaxgsNmtFUlCMQmUi64vFrnTaU/N/2em6M6
wFA1TEdfWet8HNfxsgLK5odZybx/KvFbz0iOJM1WdgzdK3sFE5l6jsiUy+4VzraE
ExkjqoW3f4LjILCQE2SKWDEGiv+vkU/E+fKe0DBEiXBp95sqqBgbZZArFO9zeGQ1
pUbHkqNFtvF+LG5o1snN3wsU51N5lx/D2S8LN4mINxAmOBQJ9ieKkbkBXN2bobrQ
Y5ATaxe8NOGeGXAGtUAcVF86Kq6yDsDv0GdLo4M1omvOP8ltr/vkZ41/v9Wj5zrA
sWtuAxy99DyxTENUS8Hsl6OxbTNJBlclOGQorNN4I9DnXDwqg1ulthkat32/BP4I
4983FwmJKlRaIislDeGu72IJ1w8hYAGEQxBGK8GCOFGkhQdistUSOEvfRYDYS74z
npISzgXcwArRRilbcbINZ6ffEbCO5eqgyTwVpeUMs9XoGtULG3xrPR01bom7K0Gd
nJd0jybZr8Py4DkUMYQTSf6pqfu4HL76bhdINryoaCiG7vGDZfUsn+7Cx0xZpXoI
AwMigz9ZadtaUBT9kICuFkC4joEnGvl9bQvTRTDmP5OlC4Gv2ry5EnaZWiHaFKrC
EfoTMCdd1WpqjBf0RiEtl8p6U2vT3QgulKGpiak5oG0djj3tucqrDYpy5NyzPbLs
I4eqAk/m0HKK2GkWVrpkbqNLJNyuQVh3qPWj3klmY5KblBx3ctk1hZXXMPL/uZBh
/yrq8Mv7bQ9b3WmlRwZbLajdO8dq4ET/s2sTXx6pD9Pu8gHp/3Ik42rpijqYVNBd
qQE868j52bWeP5ZymK8q3WBcdbLk912arNsYXNGE/+itoRtfA0MvuV2KH+FvNhD3
v0T4+R6397iBqS3tMZW9/QVwfLcOxr8gXDvmIyIf8JUVHM0Lz9HlDHRTawfd0dm/
a0Zyz55XCo+TZqZU6/d0bXe22z5VOoR4BIxobHjbOMcGBJG5iyjGd+l/V18+w8Qw
TDt93gOuLyyejjSee1LhYFdQj9wHoeqdFO6o2u3YgVQE0NIQROYnecs+5z28qahu
38+H4s+fPXG9ls9HtNb3OnlHSptyHLL8JGHuY0ehGn16H9ZQES+B64F8r46TRVXe
lDouCy7MgVLCoS+wG1ioQ3iOSlGG0dbHMTczxmoyE6bwTLS9HoN6uhVqj8tsseTc
vIE2e0Npl5F4fN2JU3p8GTcljZRuSxWd3lBIQf6JWlUIoVNgx2/0pfQVWLh0/06r
BLteKTTaIycoyxbw4/6KwrkNsl0zLTp+3Nb7N42cWigHMq0ZOJo3nE87ShmoDK84
eQ5qC675xZmpUpT6v1BaJxyAyPEVbhM0KNu45t5Y9qPlLaKU//UjiD2KKE1hC2mu
ZKL0wQyk84k1XZm/Wz7r7gzPB0vqLlNFi8B2k8sYAfJvVHFl5+3rMgoPYn83acQh
3EfO6VmGPS0O9HvcbXW5g9X6UVModty8KvG7G3EVnYXNzoDU89cY0X90tasgT5Yq
znPwnJG3xQ8agPswKyGhaS6QycGvP8lXmA3dcth6eTW5v0/xK6Omi4IQkGcwj3va
sNNd6ARlyG2zM4ln3LGsieJsjRurznhklZpnGNSe85zWMLAcaFSOBkLMJAS8OOhb
U3A3M2ghhc9Wd23Kmqf8HkUAwNLZfZpdnTWVrrL1WVta9nWNrIRsDC2jc24hkDIN
3Lzc9PF/iZQ+p6xpgZKMWxdlEfQd56L5qThxl/zm0ebVZ1EXO1wRe/zTz+vXVd8/
Rho26PWoKKnOBdaYnB1BKuTrSgM33fChtoJeQiYszqJqhHtXA0tpxCF8S1b6r12n
33I8IvTJ9RgUo9hdGtaVjjCbyZpHW4t4+8JslBD0kKN9PVgzABY1MYZyUoeCGuBx
bGEfFjz2ogDHNzFD6Pq6lumdBEsvDHkFUYsR4/nGOwDuAWHZB76nxiz4xTqgHOZV
4tld0owCoAZ2PhMXoByMosGVFiL8GOz/zhOSWHVBNcLc6wsAMzC2mLLJbejfcZ1o
CZ3+sTaUS2hE+D6XrwiF47cKQ1o6oilPT2eh4WnoP1HSVxYUMla2U8sLRw+zK1Hl
NTSrJXjfIoQ3Q/5mFXIGgxhePHMY6l6OCbFaogDi7PQqqbno5WX0h+azZNQXZUFc
O36S2IIRPaMTjmm1/P3zmI5NO00flawHKctrUwOJ2qQFu4Y5Ut3ojyFnd7kiviMd
ddDqDhD95aOfc+VD1fdRb+S+G0TKB3Tn1eyv0ovzWb7z2PlRxVO21FrWxdI+dQL3
0FB0A1ZEdIDKMOm2/SEClfBGR2SssCgQIfQJjEagQ6JThHGmhjfwdncIXRclPQaP
UptXq+r4adIYnDhhzQdD2HdFkqNh8lp7gLrrLXpQ9rQWhJ2D9L3xlvgP0ROmdQp4
R+tTjiU2tFsZzmJiQtMdqPgDPNjnOyJJeZXxAHo7gPrCTB2EkC9BW4Jm0eY4MBe0
VqWxKsgOupV/uSuwGyhSa9MRfC4GBBbHDDpMMVSpmEg+YZN/uWpwBkGcPuKb0DyJ
4I/wgNidxgMSG6XzyXDSPCVL+f3gGBmhxCSh/l9ksp/fYCZRyrhzHLtHq8v+f8/Z
/D5lhvKoVuQ2t4u3kjMLDBo8MXs9KsIgQbrhVgHL45Oc0NKtLpuhyP+6Etck2h0u
56/vkZL84bAqUmLjYivExfIlnM82t1Kd/SKPHzuP5pl7Bq5WaW0q4zmjUwOfKRo5
XU0AuGjV/At/3r+j6VZmXnNNIYhT2VEDG4lu7tHy7kdtChrosYTyMo4vp2chAdcb
HBnbmb9OWqwrvhjOLCA7uybelPexF7YjC67SgBajvFjA9+h4cIbeXMGF8jyD4Tqr
Y5IMoV0o9gR+lQL8Eugd+kZ48vLleTioCQ97ljWHZ3m5wrexfYrb4oWn3TMB7Nbk
XvRpMLlHRxWEco18fMxSXRLZTFk6X7KKfv/pc4DYSlXnD8f130Y47XkxqhwOo/aW
O9MTFpqpfgEVSVYjd22CrAlEove/heb6y+iNtWVyYWv9Oc00N6z2cmBCuvq4lc+L
q8qycmQDqUkITlNmdk2I5XT+JPZTnAf3oCs++k2e/rzEec8md8yI8ZW8DTYiyfz5
BXc6GRg4IwYJVfDRmIbC7JNa6O2bhG70xc3WnUrDYT9rxRUy0E0HOz04o2ROTxt3
MnR06qD1YVoHiyKyEAyYTYnPP90qqyF4U9LFCebzapuZDYOcVOJhs0TFpalJwPK5
AhTK6vQTeg5hz5PPTWRwFRpdgnhV0ZfSN/Kb68QIdc2aaeDYImyIy0+ZBTfTApjT
cjJ2cDS6WZB2VC+ShErFLagA+XN9JhY7X8U9BuFwLL7ASd7ZY26b8mO25P/6pzqr
BURoQOFggSS0ahGbArv8DrL5xsvBSlbZuyab5qhLxVa/iaqU5duQgglnWZ+MSoSS
/Xr3FhOc3rLWaj+/T05dDTvwJFxjhp7KXvlrAJ+HGA+haooe+UZyzrHs7Hu88Q6h
Ae41DtPi27+oq7/a4EeWKW/ADh4UkMqr0lRxdYjUO6O7g9KsPU2wnxe6XxnQpzBg
/JVeUJpO920BMKlg7gp10bq0EoZGgoLz2ozxUqmI3D1QXFmVBOwwskMUERWqPjIH
u6gkCbzS9mk9PQfHrbn6cO/feHiJtw8cNfB1PmrvubNe3WJAk1LluPv459NfT8K9
YY1Ij2zKauSIC8f1H+Nj7NPT01B4UyUSenDoaS98qy9dCWzh6qRf3tUx802aPCrr
MjuxCFggDm37fTMkxsaUWjGGwMeFn4px3Geg3kfsfaVWpp29Pb8TJzstGJ0MMPP9
WgcnuTGCQI/37F6F4BgluKZFnytElmIUP+31d6mBiLtPfK0zqOXRnwC2yopuXJ3H
6zzvRFTOxnGqt/61X+cL9CXMqtysR4oJ/b7+cY+Qk9x+0I/JvQdCLl9KHpsAzn9n
Kjd3oGipV1PXhqchLgVw93FXgTTNyGo4pkk16Yxia2sSjX97WmP5jKSjYVNoAbV+
SGv4kPNnahW83necJphsHETOAoUYaLiBPVhtWC6ZJZTdmhxmZR4ptRza99/Fg1en
3v2pC5kp4JXLyU1pW0x27NGU3eqdU+bKYxe4zs67Fcrb49m6XC7rjG6EHMo1UMFF
fUOkW5ehSXORiB7soM8L/OaBQ/1Tn76KBVjxMPXm3tjAny6ExSzyCJ3JM2B5wdod
R5GUs/itJLYulX8dKrQYr+2qU/37nPRomkh/2gpV7T00MTtvjqnGJ9QeyXNz5VnQ
Ts5spSiOamuMPFdw50dRtW03y08Vgxja6X5l7D/Y97HNgcvEv4ykOJgnKfuzfKDj
IQDeLJXqgI0JaPEe/chjTL3b+JcE6765eYNiE4cEf2fjSvEA53XwXQonv8ZM/1kJ
C0BwUs+jANkclUDf+9JJ8EZa/woZZ+0i4DgFZ777vikduGjxezYkEcBp4nYfZHkM
k6qm4JoEevumb/exNuorGojbzpbr51J3PJTr0j7fnRjUvxq8bx9dS0B7V0Wkaa2v
IwkYWXX1weaCarcQvE6aPM7CYmvDSaHxzLXxF/fv9HiZkfCYGTsNZeXeaubutshh
prhriSYIidCWH2qlZr2AIH3jTjmxLakQChk8+T6xEGZ9P9q8HXX3wGLnIRvS3L4r
YzKTPBb9eIl5cNlCA1lq12WwBbVmCZeVrzJ0RCGh4hd7za6g5WpSxsNXq+NBgpDo
QDiGq+NrtQWDIz4yaW0R/tpmpBu6XrfUJFZ7va1dINtw+IAQqCEHGM8VBwDjJ9Uv
8/cemcJgjmSA/V2w9Y21QsTi68rwMn6jaFmvzb5F7RT0cOhO9EozeCHPd/ylPCcR
YJ6cGq8mA61qkrq4e45g6rA0K4dQGglw7DHD9VkmBLaysRS6oNyIPtz8iYKDmqhN
zn8ScTxDGd0xT40BOlEddTYZH2pyY+SmCQIZfJNTGSmlokE9zfs+icxGhjSwCJ2l
jaeMIaOqX86j1Bj+Awf65wfMr7zTLfXUnnYATtEws9ajbvrHy28MkfhRz8oPFqSn
DpZoEq4CkPDjLdWISCGW2xiTmHyGkDPEf4FN3BxNUbgmo/mPdP9st4ROzZdTy8yr
kcuUSsYVQ0HStqE90MvwcU9knXz579xIVcaaT3n3WgCjqM4ID20M2wpYqfSZ5foC
KyWM2uHEwILrGgUJAeMJYipcYghVz7O1gVAz2JJHUQy+qpnJ5i/iYvvAJnxIHPgD
lEJ/L0PV0+GnYAcm5wxIYMOOW+GjKBsIDccH3jc4HeHfMEkCPFGocYxc8d8f5R6e
BxTNAi7vlkHQ8e+nCGbhu6RssHz0V5rW0lt9ywmyJLtJptmLQtRbwouMPvCa+gR6
impHhx3p67m7ETyF9kb8UZ8mDNMdMXndwx3KTwv1utgyO9H4CAD1b2Oy2Vghdm8s
ESHVjcMcm5NBDoQc2Qq0ktu2RNcLb9hLJntJzQjloGOsJl9xHWLAtFGk0gwjuJA4
cNyoBjZwRYOaA4/PgUmdQhiqOQ53pZNf86ZLC4ZcTDs1msPiu80L0RuaQXMSwZGO
/L+aaL32nDcUgqbIgdPqBOscMAktn5HaMH/VcddiNzE7MIU0zWJ/Z5rA4SLSfaae
tVEZ8oRfHfQKS0OfS95VeZCnkjKOEEO21nBanlAFHauTjKsYEbozn0m+WMRZB49u
FasoyqtU5j0JcyGg9nAnt2cwnSkdGwnHXZKFi1gQ4ZIMmGBJEYbUwB5Grx2kEtWo
/5nna14FWk0fYuunQ2utPHn5YL+xeVDa9A/szJ+vGj8dRVBCc7d9l4gfbVSfj8xl
Y36RQI8k93UFIDfhihHDXin1ry4FTFEggn5wRdGtvnQYe+YoaU2TFBMkKOeyXPbT
sZK91Lm0eU1xrXSe+YD8RLSVuQrnnexsD7OOKlN5OOdOALIpu+HffNYFHw+yt3XE
N9vixbEoO2uHWpVQeaAhERxPHqsRE2Z9H6izgGxjmp37wrdefQqaK+x6hGUD3j5a
/vTsR176PJsmL+UoahCl9+X/VPyOGOTKKM0HrrWf8iBuGkysPk0xmoZmu9znfTrs
ZUCibbaEfiObBA30wxXuTtyX5zVOsJLteqy1bUMzcuatPiLjYOJHKbzX0yU/GbYa
vMQMe+MJw448jQ9YrezIgzBvvDnXhSTXp7PyG00bOctKbba4wjeP/ZyUHZRA7+ez
k/NhRw1i+EeHjf+GG/wK+wWFpS6MeheX6j2AIMXLmjV9yGgr8dOyjHMpCkfmATms
azOvlWJ/QwIZR+97GpMoPxFohs9WRPnVwIjj1VghDcbP75e9/rllIUw9OyJF/EOG
pVO/I8sySR6wYADpBbKjtfZofrYKGP/B5OmlROoXF+Gdf/pU8MP2YS4nx4N07i1L
OpEaBCv6FzHp7aUUhcvVbDbMoK+iOIeTJAXYHmAnzmszT9Waxph1UrwaYicUpieN
T6cCou/C1GPQkyPjOW5RunCqWKr/5zTalVxNC+ke5V5z4pKMKUA7O6wBWhCNVGzA
TWRKfRSIeor9rZvSEfgFQ7OFhJJdjQKDS7wWKMeKt270u1xavCKYIOTrAzFI0vH7
nfccHYPetdxXf1okPZIpgeq9LF6aTaqRBVZ8MaZ0QIZUtybX6if8UQptp+xYU9+B
jD2qk+y6IqNQzjs2VS10mr1oQ/EXGLMbrmfjswktHgeE4pfbYmWMcZD1NEVLgque
a6YM0UBD46ELFRnFXmJhRRsBu/rVg/J+9CoN8SYH377nuk+/bBlkJ15+PrEHKO0F
m4nQa3BNKTa1UX1qHnQIphGtnuZvOLpZYmuA/5cHLHtljKIFRwV5+XwS+aTMiZG/
gVUe6YF3Z145vbJR1UHwuY7V4qso1E8nFEGzK/Rqpxp28KTnxLwExdCnxFaKGARj
qg7LlZ6gN439i9zAOeSBgs4VYV8Ab2WNkq407l0v4UQhe3iZBwKoqRF96Al5cnYq
NYPYLa6MWsq7VPE8bS7VGfO+WQuz7aLnnZxv3uN54mwOD4GgXwVxrjnx3KjYZchx
P5SAIrxu3oA523Ht4/6JXB8hHfWzTwxLvrRSAsodTS2bIpIphul6sehj2Vll7M+3
4aRzIA6KHhJAHJnQPrdXPaOQ6oArwlEKRNhTTKfHp62rLvYtfPYXlVRs6dRPvlRc
TeZuufKBSuYQufV6oFBhFoLaBQGXCEF9tI1j8HjIKqWQ68W7UnlyO9LXtdOuUNfF
1DxdHaioKx3nrMiu6FdsLIxeePpoRGhv0YpE2egpdmgIRidQ85VyrU71+449J5hY
2jJ20jdc69Q6QceJ73+q57XbhmTrvXAi68EM962incdHJVRVNAJerRvD+oosPxAp
l/K73pgDzXc99aq61UD4txycbNzxwLNJSd6OUHTnk03m+CLXfrmSBRe2Cfx0o9p8
mE1520Y3p6bUTiLVuoADu0ujH4VHDzacau3DQKetdXHWVX9PzGzdXXhuZZop0t9u
V9zzVQERDvDMYz7ubddRUxajFkccz/CcKjv1Ipo+jhS6+uzratvtovofZwIPlRMr
JnxNPGXh5AcgKe0Fbsn24Y9pH3DvvFl4Kwv8xnyFD/60+8oFDnl9d5358WgG3qD5
SMMKy5bOtj0e5eBURd4HbwNTbfcXN3n6JpWAGpJEqhvBBY3eXNDNoumjhiNYRNyx
nPOq/CT2Z0b2y8tGMreeoClhoo6+nend5YH1jVzEcteoogkGRDmJGi1GGBS6IcIu
o9ThBXcqZLidAkvE60IW57jEiHZdj5MLDiR5Rc8wr8tsAchO45Kse1HF4aUKCw47
M6oH6Wc/jrXi5zqH4fjbE4vjFbqvOwTvWQSToBfNij8LDmwwO8Z4ehuPG8T7in5U
Rk2DETH9Ynp5P5rNbUM/vFItrimbl93P4fLfvxtErs2znYTYypP0HP7kcnFrr7bB
mC4eu4eFxm6HW4nNUmN4/bTBXZqvXYVg99y1c6lO0CdASipfD41uNjNztZ6IyQS9
Y5LP6uB7oUXUHtlXBd/YDjkABgT6kMG5eO50WM/pXmgHuB5k0Fnaff8Cke60gxti
x9PE1oCrwAB2958bs0SAaChVeB6wPclBO+UJsEMkC6S8fhUikadrRznCgXXIBZ+R
HT8cNOe7JldGOxiX5EUnJT8zbFW/Z51G9LauOcuA5CELicYwk3Zhnxk/pJ24Kqha
qurK/P3o7KR7A6wb6RmeynZsMbn2AFo5PDJLP0Fj61zbOZ1MfLqRXDwMHpNN2aTY
JFwLSXf/YtFN+63o2+hbbQ+ddghyDs82r/P6PIdKHzNyyYabFkjeN8qy0K1LTJhP
JhiSOvvFVPYm9RJi9o1Y/a5G5+nucR5d8XdaWe2LOLkMZx7BzdnrzKRNIFoTTIug
kDer9lV2x+QCIn0l+teXehyMUvr9xv+yoc/6Vjw5jzbeOKdLisHWIsAxzaKGNZj/
ClKBYqvpNMHW/p999DMxZzufhBnRjCa9onj3RpuLzvSSgYPRSwELGh5X7Z9jZPwf
CnHAdd0Vo/QxdbwOxRM7PJW5jpECJEEwvedBbNcfrHurflDC9+3fEOhLcD/gZS6G
ym1m8x83xo4126695TE/k9EcFaeztQTj/4m1O5h0p0Tb11qCw0NLg1AKT30b3urr
7JNUsHviYpYdUPGB9Tq0DjnTAM22o53Jc4pbri5823Cys2NwrGZiRV16WiHK8gFZ
meW3xq5mgJc0gc5asI/bT11tH67BM2BWsERyPuEXi3ZsYMcpmdHPGYjqv5NZblsA
1hebS0iXLADU3A7+bQkjWufz1AUBU+Pe+DQIxw0z9t7bbR3xUNqER67j539OggWL
Bu1zp/TLcB2x+o32FabViJFss7PEfUYhdBkUfgWnkL+jcMgJwYhvA47NdZ/7UxOz
VniX4uNCyOKbpXbt2E4gU3KAz8dshxgfaGsn46G5ECWmLcP6Bm1CBLP2ZsYiRVLN
ZAQjGnTunBDcl1e7TFFB67UTVD1hkrgXiTFczpwyCjUbgxb6clqs2wlPcaFo32DY
vLEgZkzYQGTWsHoF03RorgA3TREIjMZmKHApvLY/u2zNcTFSxN70MbUYQHivabAM
VshuaMkH9TipuOJ1JXGVqZF7RaYyCD8/U5XfU+9kV4oktF+AZvQzf8rWJDBidNf9
VftsCZQyDCQX/mHZ6smwjnYGO5M7znUxvy3ieFxeZEEVv4kpKzilCBXTKquefXAs
cU3iiXVDITjNegY1wP3eWzuntY1Ij51nEOVeWszeaX637a3Zqojdv26jzZPdpdP9
sWuN23OBQlksJRzDB62kuUmGHYqeyDO3c44ZW05RJDYQBFI5SP+F1BDQcgKnargM
IDzVhAWdRddnJuKlC3MmpEH4PGIGG9YV6TAu4hi/J0+xkiCVFYBZAasJyRPH3VwZ
5tqZGyhl6H17HjdHrKo1l50D3e2SernIzquKaQHfiFCGNGYrAqzmsrwhK0I/uDOX
IKyeyedJFSFZ52RrzLsAPgLgUabQmA8AAzhutfRQHQ3cKFw1tzybczvWPTXintlQ
5H72NQL3cUJ6RzsAI/I7qmAAItF7Ht/+mqreOsIK7+1DTehq5hPeH0v2PKiSemkG
WI0gGXVaXOyiL8DT0q6nHTTt8bGfxm/OeIRIE+kXkG8FFBXf3DGz/Cdc3F8q1nh9
/JbS8iUmUM9Vr258C8se4lrG1gXdoO5Rd4KhJwI0e6f+FpMT2rs6xUmkir5diYC9
FrtVdrFPCpcz+2BMjKH38ZZaHIT4zfSszdnMzBZz4XMNUjtClduwSufIVp82jksW
CeN8RoLvngKdIGdAAQb1KyN3VwGwGGXtXeotnYSmcs/71B6AYxHv3WjUxGNDrfJ0
leNnZu9PbsolHBq3bwh4waNJGfqO9PCUkK9nmEpYft2PW0X7bH2ebVmHH/j6JjRe
ZLBn1bLWlk2wxH1FXEgAq4dWKOvlCbV19Z4EaZBg2gOSKjYzo3E2kXRBvo6UOB8h
7zzAOxhKcL8E0bUWRWZJpESalcP0dKmxLcLV29Q5shpYI3U6KMrbUgb1im8ZGmp+
TlEXos0Pm8gasHhZG9Lpj1uNRbenAlXzncUMgP9orlNNuV63JUFkzMTbI7eLWTq2
djkYz9MO9wOL40TC52vupfBUWpHDMsq2Rz6vluJuJ9a2qML0FcQ6IcZOiDMlvUCm
KdiRX/i+4O3vBRNtYtvV7UhrLAbQako6ZIqfb2mq5IGtjzEN22ChHXVqzPN4pOpp
FSzvlJpEDPC33G5NLE0FPHp2tNFTRJmkF8RL4iJuBksUmB3oP8hR5AEW7fLotLb9
XrY+CUKXyV7BeXz4H0y77uUsyhyV/aWLDAF+adT7imMGFpyNMO38f07Jd54Ln2NP
O36B1QZFR6zWu+3FbEjsTaM+hcdtV/3vUl9cY6z49ePeKTCm8B/0ZwP682gQYTsL
8LoSdkEKvnGXfLsUc67G3gEDPvllWk3midsDrOg83+fQGQIM3I+HS0u18tSLM07r
SdTycd9KSF7zxnZTlGpqvjeH3r8i1RMkhWB+T80fIF2WiFmMikYizNfAyemg+rRI
KuqauMnAGh+LSiD2pzEziviOOUcufkElyyPEde9enb5EUbwCUQS00ydAOk2WALCb
/r8K2wVo2Q9/u7nht9JR6stGTVtxZeKs7KiVtXISnZBfbhFJIJeacTxAesEooGuk
X05kE6IghJDlA6t0ZXFwIG1D1pp9vqjFMbf900R4rD+iLn9GPaMoTXkgu0l3i2Qb
UL1xQ+rgynpHLC/BHE+FMOF5yQaga/3knfbyESlGqZ9gW1YJhQZcau1CYlTv9j1n
n0+jNlCRVvlDnC2DCKkqc1ZCbShPY2/cQvB3sJOvBHQrz9GOWhm0kHQ23eKuHAW5
BY2N6voWp6LgBy0Qz6WnWuzjYgWLBx/iRb5F3Vtk1R0yK0Ze0bXF51ZOJs9382Dk
nRldIgR5Mk/URJQIGu4WHVs6XsirZZic9vZgobpCYKDrimlxB5oFh9Nr5JzmrTg/
fQdyiH9OAdJpDrrTd0CDCVwMdGyLof2s5BJlPRfv/jllaGEuZco5aun//2Ntm7Vo
kb3H9OrPqkWsHk5zA6RT9+bVV/QB+aZfwu6WBud9O//sJTToLydYMm985pdOJdsW
rhp+h/MIuHrqUe9bj6deyx+/ufs2hK23xQDyqkL89i1bmrPvkkyJu2iCbKz1Juzn
b5U3HNCmM+0kNJMNQ/2gIO0YHagJz3fBXE2gA77GOoH+V2DkhHTs897BGR4AJaYY
8fseG0k/F6/IvXERA//3kpbEeLuba8bjwzBVbVzjPH6BNI68eV00xgE2yucjVll0
rzuzAmrkI/cH6MpmbqZwRMhRsgZmaqMfNbVgc6zkbmhKFS7wAuUzhsWa7qAyqwvV
u0niukkQEXYtNROd07mUvHjIC9faVkTEptB5wQ7JXD7+Yqug+BeZQT2jt5McaNWW
MItrD0jz0EKscW5CRvYH2ZAkR9J9OzfxU1B2u5xRjKpPItGgm2JdjznxpXPbqHbb
h2zUv+DMnfRX4uUrH8MpBCgAyehaIisU5M/y2uhMk3uPheKZ9qH2L2Ykt072mIh6
9JVoxeeY1KIwGUeAHhaHHaktMDVTWkw5OZe2Cpc/nuHKZ1EOvv4Je5QXIIXmLHuH
/UdRpLQx0RIzPcqxdxkwBgBHH/SZZhKASMFXj2YE4T3BeUNHps7q+9JhJf8OL4wa
LRMjXRV5ER0PeEnrVJnTppGEBfBSMyo3K7n2TECa1wqC4xiTn5r/JnZhHBvFgB+/
IO8WLnfQoZ2mAb3v4aHNUMCKibPbBwIv+Bnd/sAEDtwR1QpHC1OGbx7BK6evZv2S
wJz1OK7MQcdbGBsnu1Nn5lUp7Kqaj6k9c/S2RE+oUki7VBZJ4WYD8cb3LVe+QnM/
/vDoWP4XVoFDo4GHHVvBGKLqm56Q1mSyaL5HaKUaNGfQrVjIIfLZsGxgmLCM8h3Y
OdFugXsuNZlAGpz/c8YM+bY2CQm/V7Ulg1ndX/EbgoNWnYIlZaqKK67UWhIWkgsx
goCacJJ1rdAdD5FfsxFiK+IPfKRPFfnP3KstGYn+AHuM4nUckK8BWb1EA83wQ++1
Fb4+D0TerrBmEtmW9lWzCoMhMjot9WtGJGAtkx0/kZMiOuT7AGDWBbu+CM39SAG/
6nlZzsQEiAuAR0XA4rwJx/ifGFjF4iERokI0+YeUzFU24rm6XJA+naDBI4viwKBy
vo1TWr+2vtipZCsss/Cznp9jh/JZ1CyBqYAMWDcHEmMJf2705hT6AC/8WvmkHpTM
MDcsql6mQTGSxth2qjfNtU3rjVi28oqoWLNPKvmGfqCHZ1Tj2t2lIp+Id6ym7/rz
/Lm1ANNLF0/xs8oge1FjKDf0QiHMMD5u/uySl9rj4WGq/qc9Lr4dNZclss+wLwag
Rts8fnb9lb61d0Ajbr5pc/OTAGlrBwofxHL8oePBfNgTGmS3c9Y9ySEQ8qiTYcAo
TNRzSbNfQRTCHL/xD5trgJPQgHF105JB3KTaM6XQ8OnTps5DV90Q/XJzhObwo06c
jYfvTGmBtumOexlID55QNyJNOAAwaUJjix2hEQfYuA6RqjpYHTRkjjh4GlMVVRuH
jn0YG7TMpWTcmbJJgAMgSFpVN5Ik3oqtsNFryyqgfgVjnHVmIwFBB6k4LALJuKFE
KRWuVhSgGFlnlJwkl74wT/8vBDEhDy8fCdQlbxxLwH9QH3JV6oRidTDfA45kXYWZ
pOVWYYhBT3OZ2IriniuNxGcoIOkdlsyfWeo/S23jwuAacQfKeuQwg7yMrqDClpd+
zma1j9EQweIC05GQK+FuKbfdy+MUJKAg509ggxZypugxLoq3IXwvNbI+dc2H+nqy
pin8LGubjv0kLRTMjDcwJRyDrwEPJhDCwIHIOwjHyCEFU4h8eESQNLyh6U/3P85E
z/+ANmUSfWM7qn9W1PzvHAFJkZySxR2dW85GeKI4LDHQMlYyrY3v51LRBdqEb5Xu
gwkyA8lmaHotV7pefuLsahrOR8oAdtVa0OPzeYW6mgMNWREELRZcvLOwEL7eE8wT
A1SNvkpG+5c9Y1d9exDyluL/+ynFV7M42mVSbT7ffF9AcWj/0pBcjnh1jh+vr0Rh
1TLyhCBwN6LBDcM7YaCUHTMLhmkno954GOKxKLyg0WsOUeTJEvbUaF9NnZKdWICP
8pii/dkb1Hh6VX8TEm3Pcrh6hm/t+jik/dEKCv+zIpT2I+YbkJ1S2bYj6cH6apwl
VLpaROM7KOYU9Mk57Gveu1iH9I0cVXdQySK65IHr26bTiwrBrYH1kuPSocujIlVk
S7nFBTKkY2shoeYKTZK5FCSiC+BFUgixDpI1tA9Q/efgEs3CkegfYEj3FzuD+vvj
i86wrOxL+YtgUCxT5pNYRLPtVVjr3jmrsC2VTtKGEGImFkagkueykHfCddBlxveR
7VlIo/WJVNGbhA4qTZW+rcnvoXb0xPkjrDpLpgzLfxa9g00h/SodgsYfGH8ML9lO
i2ZCpHZutBnqnTBXQYKxW5ufp/atOtbBKLv9zBdyNCuqwFzxjwaqldbmEUuBVrTr
EUoF2XrN3z+PR3bTVd++ZCJAUvH3SRxe+4DCy3koNj2yOtGOvH5Uk5+SFHqgiGsc
qkqf91QRt8E6N8wb7tUja1TzJ+1lFnWfnqZPSnsUWbunxxjo0BXIBrpC0F6X+v5N
JGstBQ+0MAgce+Y94TsIVm8S8n8k750KTHEfIs+KHD0YxwDGPxZBIeyw16ewvNwG
hcRickepvczkFqNtlab+3cfL+EZMSO5VctGkRRF0QRChC0VZ/1iTYqji+w3WVupv
N6IOrukmmc2kvm/ql4EQf3X6NvUuPkR6qDYVpHXuRKl+EiOYQ4Xb6ACTwsTQqAb8
HnMskovteZ4cc2mcBEGqVanYqjEUl65UIHJ67tfA6cjK9p++T/fO+42gAatv3liK
brjLEd3ddzkjBZEW8mSfVxZ+MT6r/teHloyxdTnmeGu2fW2MlMk+0at4t9yGoit6
t3yUHzT6Glr/TN3jt8ehFzdCeZXKWk2r6gzngF1rLPuMKx43OazghXhDEa1kF1a9
8Oh7bxXEBdwyy/6qqPTx2SPq8FfH+16gsrxd+JN/G9o6FfwChBxmESegj8yDz597
dWzcSy9yzaU6i8KzTJDAi9Q3NIo2O3mEHU91UuoT8krCiz6gmzeReXmA34cBzLoz
l77VTY2MxMNY//a9ttZZMls6P3MDH+McnZyDUmecJrunsyKQHPTYQHF54L+ik21D
/BYS4Sd0wFA1iwRU6eR6pjsSQAUn7CtQgdlxjd2vDTjJ3et4Fe/vQkCJ7XgVLYCl
awolObG9T1/lnQSkc3i0OCrDvS6CpeI4RGLxcaH68gcvH56vq3eBw3VVNVQAJUAA
itD7usAYAvqDlKghqXK2Ek14FEyWRKv7j8DU9z3TDOmcPkUXsxgKKw0jlTJeFhLw
stF8ej8vIzZxDHz4JdEXsUa5T+sP+AfMqkm71agPXzAynEa3vGo+CtEPAPkTJxbR
FVpGiGl+LYYcOWJ9swtxC/85kGwiiHf0JomIjhFAO/iw1MiW5+PAxWCYC76KqyWW
sbtFJpoerlNqcLNkO+FSRtG+uLcMMI4SeSog4aPXAz1+xl9fBwnVa7FrBTQogpvz
DvnLxrGbAuQksnKy1t1RlxvU0ExvWrjIdu1B8oFFHjY7J48X9F5crzV3wWIhTRdA
DSYTzyArerJlza9O3/xTSUsrP6JbvpGdHrVOrobPQn2IkN2vxbjqLnsE+3CRYB1M
OKTGpDarBSv5PhZMO2kgC0eTfSpqBZRTb5mWtSqb5mpkY0NvWEcBHJG6jO9Htl2+
lDK/76yuo33YY2nI1IB5ToVDj3Sin3mMFElyrhnnAR3waTwLgN8wEIyPCVlL1LCp
okZ2Vl5ZUhDBGkl2BbQZZGZg9pBdWFMu6vyjIm7EVWXvWdwZt3uf6zn+cZoW35xD
kILzsKvZuxOzIv5ToKsNXbJjTJUoNBQotRjnhKfsqNb6GrPQz1bSw3aMWJaLJ1Hn
qsIT0G0pPmNAnrLOTvjNu6Eg7U/x3iW/3xHKyD6I7N6bMKLyG43MGmt3ppKiGVGP
QnTd61oh9uzJMCJiQKYpxcN3FA/PHL/BTanL/EgXvcwXhqtCAz89FHHnGCqNgS/F
SNWvLpXePddyoimLI1DV5ifQCs2ZqYBuRmRzyMkxQA5lYFepepJjdmX1j1zd3iJa
WKSDWOzPAmjRYMns0tdSO+5ne69i1j0R7jX4X0m17Wx9fK6Ij4Yw2ueFMWCnHlwd
IoVzynWOtZxQRyVvDsenhhhrLU+A2RIrZvbyAcJZmY5D8eT4r/CSdtQDrjKh9Afn
eUbMWo7/aV34/ZAWaEltWRUEozbfxlp/o9OV/6UWnh8T3A5Oc2Z1wg64X8kPvrJl
Pb05t5kRhygLX3GBV0a9enFmcdoTDTrmKyzo1x/4rH6Pk3DEINonAETORSvlrc/4
O2CguutRqEUyo4qjtIDoJ2+9mX4JzDZLlfqZWW9bOD+XMbx63ka5LrhXZF4oCsF1
CNfDyJP4KJAiv2+eYv3/aGxVRxbSpvfWniK/s57KD3+hZ/uuS9v0shzMs71lLGgh
RKOsaiy9uKVS2yMT5nYVAyMLXRrDaDcTnnuRvlg38T0JtWIcfY2hrxXZUNVyXOJq
LwdflmNz129rX4z3gLaOgDojB2i+GBU/fjKnsgOB3ruwEdcFcrpYZ/catHXi9oft
GAy5VM8T1KMZ5I9K8BBYpPgSoFtidwHzNcgMQ86jM7p7Dy2dLwJi+A7w5n74bdey
vjuwaJJqEZdJ/xE9ZT6UXckHSP5C0oJewMUNOf/eO0bLjYeHY6kmO8VCy9grb+/X
S6lX2GOe494Dw3UGZzA1+13qPz0OCZWoX2NileirUeRcPR2rDjhCIHR4dPaLA2eM
uBiCxGa7BddYZsNAjPTtDD2T5XXGKLS9+kCGb1Gm/uRmBH/CHNC0jl4MRK5PC8Zf
0wHa838OEEPPJzSADSWv2LIJ/1vs0iz2yYf0nM3eS9AYywV3ZAMHILvHG9+66yeH
nDmW6bWDFQnRQLTaaF8xLtP785h8xM4Pb/smNh6KPM7Q+jm6BwClnn8i/yn5LJn8
VX3l7/YqXUeTp1DV4PivkjLGSHRfMbOoh//GU4nLXoskwo2Si8OrUrS7XsmXbcCW
`protect END_PROTECTED
