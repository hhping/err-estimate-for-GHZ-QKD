`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2NMKsd1fwULenzhxZflp/LzH+zUcnhxzKvQxqgfaCccT1KGLX17Q5o9yHxjCMliR
d8F+5dnDJQQjw2pHiVsbEhd6a5RrB8+fqyVsGnlScCXPOwMgQFZi9NR0iK5hc99b
7kmwim4yeUo3nJJ9Pjrrw7vzu6GA7ZOPySzqz9b3KgNKqJ96lagOg5CWERjE0/ro
+Lt6agbBGdJiBQYyyW3RqBsxdZt0eb4OQmTLPR8L2Txer3GLdBIQSRC6qZ5g4eAa
XhyLBa+k/Azr/88CUjbFtXLDyOrIXORG8TReEI2jRXTalzj0nApKrAC6At06WjJw
o19pg0XKNZwLhmGqJMVB0YPkLDEz39wikaovcMaSWK/8apmNoa5ahawXaTVSoc9D
/CWbB2ePxojt+TeAtAxNGgb3cYjDqPOqSH/7Qxxu3LrYHunFQNt08eFzCpafHH6T
BOPGfI/eyP1IspK608eoqs8kN2/gmtYBiaWNMxi0mwlj5iWErNYQ/O3UZ3xy8yYq
NT/Tu0sOOQmbBDIU0Ol5JwZrorwXrc91ZIlwwcQ19oGdWUxKxQKj93AjwJ+a7Ud2
u5nR3lYOjtkBKkV8/CRJ2kX6Y2lSxS8WBiXRTqJrmmD1hNLSAQbl9RsFDiSZ/E2a
X6mrc6qi8SSRojbHc9MmABLxxwcgk+IsK8+cdAd3xocmSq3+TaaDlOhsg6qGIRFV
hs2h7JjXQL04UtMsu2O4MOe2equsUTutymve6TSSdBk61i6OZKQgeQFdAqi5mK6Z
n8vZLXftvI7HFRjhXr/49LvUIx9nMnLXZjv9e7YgJsTcsLs5twdB+sqlL4ZmStb0
MNgG6QqMRYVRMjev+QUlJOFYAG0RZjVq7iZeWG8qhLwftoveDTt7ynaMm1IjwK9S
YuafG321aIj2fm1QVe7Yg5YjWWGHehgnmE3lg4ZlAvfZvLyqV/de2jEuBA6tP+zT
sdmqQN0pBoI3MnMJkqe/atnE5HOZJ8PMNLJ4Nc1k5xuIBx9dWSNPUDV9sTdJ2510
NVs4/QMGRHsZHplAOxjxvEV600SHuXnL5JedcTcry4RQMPS4br7WKQY3t4Z1Pvjv
ya4eYNCXRALXcbOQqiK0aC3S/rx+k+SvNB1dwhkVle0pj6xSyCyUf+GsZndG3Fvw
3eYZvSxkmaeyFotVDCoXDcByJHLNPIbxFWiHcpIxANYLLnbQ5ANI2k987lcwj1BH
4t9xZVXjbKeEhS7yxq3RpVOINdKefXp09tnz+FVW6X04S0gn3caL4D4mVoQiwH+d
3u9dX9OLCAkDMEC6GcuJPOkPtYcQXKsTXImvMr099GoB0CzGmAFeqwZ+sEDI63Ro
MnsTZF7NLJVOvEzhmugq9Na+DEEdOMhjo1oS6J5x4dTf40AMHFz4fOOSGaSAEljU
ezI10uHF0mN15rkZW6pAKKOza2kf6GC06OjtQBSB8+NVSOw5579my6zLiczIZbl7
pMMDrcFbtrY6AmZLaxHgMwtflxaUbcTPLv5/z+XWoQuIGnREpXOcyWgTnEsK1PKe
Kvts+S8Yks89pCitHdvobHnyXt5dawZ9W7oj9d/z6HqKu/l559qHJB6IT9AW4Dk5
dnmZfgQW3ZR29IpTPKOiJGBMxDS9fzuVMcXjTZDoOFjtAxCDj8SsSn7I3YLpzYKF
SK3xfpllagPpPWD8IB67bq/XwR7R1R9vUKeq7SahBE/110HMdQUZZ9ZAVncrcEtN
ERp8MeFbz/KdgXst1TQA6mezHI+Udul9wtggEdtWtkpB0pPRpUv5zbmzKCG3FP0w
ssQB8B+JQzYId0L/llG3vYPCs7V2rjcGE6EEFd61GxycVRpFYqndI4NiwkTS/Iky
BwxCvTGLPMflceQ3NkbVK5I9tE2pi0yDFqfRWPAyIViOnOOOz0/qETiY6RhMnYJW
5HeSvy9VVldo2M92Yc53qBrM6+Ytvk0YORaQZ6UtTUBhHeXalw0NtanAiKrnX8oj
yE2eVOxV/blOP+SA23Rw/6TPMV9Tv+j6kdbUobHVEw1riasoP24/DFgMBE/k2Nt1
+KyXvQqVfDANKCgRN7yaCFnwH4uNwi7AvZD8evd/XxbUb7hJvTmVDki8UTHPaijg
2hYzs9tnriHE3svQ5PBDsTjbGhwf4GhDxrWPL1lfVAGVJoTwgBqn/ls4loywMLKU
+nMLNqFL1E+O9S6Q6PgYuVd3crOuTKPhbG3OjyjqUaG4qFraOAPc1PSTP22VpzRs
jf8XLJ2PWwbnE1GwZf1kQus8Ht8VSN/yg/lQI6KFYYZpak+2rMcZZYgBkR4zqPC2
E0WL6LlmYUeAVz7ZuqkqS2UFa5QR/xs3/h3f4nQRXs077CajL0UPHlt3TOftIZBo
noov//jvF3AJl+UWyOTgq+lsokqc6mzgFt3s/6OgZYg89vL40gq+hmaIQvS8LNNz
oTG0mEFRBzVA90/V9C82+3jyhB8JDAOZoN32lZ1EGZIAGhJSgRTE1tIqrHIND7LD
LiOPdlZ0YsHK5XFb8LrOcMMYO+NgdRZGGcH4NPwgilCJmyG67fyT47ULmILOxupl
GPouep0iC4PUSQ5cIQJPLEgBvtKe2Xv/cDJXmwDfw3t4bULMu3VganCMRibjbtzY
h9SnpVc2w5r9tluNDVHdua2dGQQtKhZcvdsKv4TGojP2KGtI0GbTTZXJH9zsahZA
robhHliNZK9pn83Sh0wn61APHWZAkfeI7o5Lm2slP21hi+L8/9j4Q8QSXdp4Fxrf
ius0Xf9XNpfvouxk7Z/wq8rbMqBxmVNZJN6MiZa/5eNkgf5Z3P7B/FjKUzs1mMTK
ue+zT6Y/Dpl074Qt2xbBDfMGL9NPVclU45WgdoVzLh4IACSkeAxowuHthdIJhygZ
078mpWU98lVBDPwt9kjv3iX4kEUDaMH8buI0lv84dFJCOfGOEAG6wLA0o9eVSJxJ
NnhZRWd3J4C0Swyjl/S6WAQu6UU9PKtZQaXWDggcgZSV6lmTJPipcCxMEyWS4twL
1H5dEeYYAG0fCHRdCdln3B1IW+2P9jUPrWQULU6AicqVF1asBg8Bj+eApWIXvPFG
FLXBrqURiR+GPNz19roqV8PMjtnqTovpUtQBGjP3ea/FhzgxSicJHpnkCz2vXf6+
wW1JPr313BIX/Qut6JYmcHpbTN6IUGm7woILOLvgkPUnA0TMCDl/T2kd8hHFCyWV
tki+LzWDSnu1kzkyHNG9HXrVBHDxvlEdxPYGX/5nBEuZPhLXI9ElDuYREe3x5Uvi
RtfbuUswNnONDbSqmDORPrfrx5V9Yo+HXx3Xcdp/t/Xqiwpno6ZSGFzakT5CpXu3
WGrH2sJEx4Jt5kc6Z6HgKycXHJTfqgyy38U3RLhyFm9XlH6HEFutgzVztakv1VA5
2UogDi1SwPbRoj60AGrbAv9TIN4ZikWhvk8v4qAZGIBbHjeW29yhsRFl9jlku2X2
V7tsKFThuOWeQal/BZmm2ABfoQvlcibdXGMYc3fC1xrRDdvhijsMnR5pWKJAq/te
5PKCL0En7f/gLsnLDcSPeOc0/zgwbAJlz2cfMlL2BVYlRrR+B6jF5r2TwpKFlACo
JnQRDqSdz/DRlAUERWyVIIc7BfrD2gXMHwtwOrsdN6iLz/3ZHMGEuC8yrqLHOew6
xq6Hom4Q8sPcRVI1IOrkmMF/d8d490vj0VAJoahlnPuZkrjUGuY9A6GhyE7Qj/8P
b8wvQHl2TqzD9xqZipdN2i8n4R3JRy2P+YjIAb8j58GyAxT/JNnb4fSSvbm9w3Z+
7//GNkGtsieq1SND9dYNjCaY4NH5YqFf0IkyKo/Q3XCtZXWy5JqZk5dq99E6iRmp
BHlSapCFgt2WpA0NcaEuuPEciXZaHV3Xy3iRRh2KjdIKnmDbzR+2TwRXHGj6MZ0D
8j5ud8Vg3IiStA2WGlS25wf+YnS3ug21MeQNyLc+ldR0DdgDCv/mzYDsWZuj4ZLI
hifZf/2rsuw4cE0ebt5ApGNNcoWhzTR5Oi4mgbbf/UGZa4kG5sQX6EgWnalpNi0/
pt9GI69ajSsooN/nAvS89etjcMpwi3rNauWbImuMz7ricu7h9/kAN4SrxuoaHmkZ
36NvW3GgZs+0HS126qKWTGycE2faH8hVSSfym0GvUki5INw2nKgSr7Gd5BooitYB
fYC2XXkfllMwXwbNYZQvvAB5N3rsIpNNePKgCek55u7rvEdGSsXAD+Jj5o+fCpE5
WN13v4Q2QM3eUi9NvHp44S5RchuB+3nFTqb75ikcVgIYNdw58FR3MeZbS4pvIU9e
Z7D5Q7EC9xrYGwSZ0Z4Vlf6BRfofsC2fTCk4WFdRBVUrPvIp+2UNlvUj03U8+OFH
9u9C3iVc3XxOriQek1oOUDdYLUYA4+ayjkXVL6taDVlFnISdlZBCrGNk6i8Y/C2B
JKP8ee1I8ffUtDcNPeXdMBt50k4X0JTgC4flIL7/VNyYV35o/Ctuty4pTG+qeWnu
Ir4uxOuNYRngOESY9z53VgpykMHt4grFSyfxpCMueawXfRsr1K4IU3BXWm6ObHcJ
VZbF32rPQ3Iq+vyImSpFWqEJvF0I5n1qd96xlFZLQzzxuCKavyy2n3Xms+PlJS+D
I6JS506ZD3GC9ijCqKFli7Xr9XNGIK7cztbqVCUXW8QmzzzMXpzFLjy0woylE1pr
jLkJ8FAYOK/g48I14QDm/aMnG92dQ1g/zk31OGzBWgCHKd5fEK2lJqKRR+U6GQWW
0o7FEp6N7tCBU71+azJ7SogfxQ7RMKelCQ+nxHSRJqGncD37fScHnP2fI34AkPuE
vPsqNELA7vX/MG/PHw8BQdab59CJ0TBW7t2RnpgQOy7ye/Z6Vqz9HcVCxQY7V+Io
UzUFnxkBAwCA3VwRDpiQ+JCvSmTxpBX7UdXnGvVBgVw+9HMyFiSoaBVgLIMZMjZC
0UbErh8bJcFKGeQmPp+VnnLBC7OxLbCQw3H1R6Nvjy/gur65u1Uf3pngtfWR5H1c
Ykt7JJUTN7/eZ27EgFIiH7365y1N0bgcN2la2tFB1d87c5bF8B1PuGEgrQ6RnvQ0
junnmcmv8VQn/TKZAD4x8pfvya3ZBhwSA+7am+9qpOr+xmNiuBb3+Yo5xDD5r4aL
3KjV4FVf+h3us6muXLBfveDINRZUIkCU/yoYk2UV1HVRpvKwte/hBjX39E9ddiU+
6wrrbJKT1GHjIUnRaqAMmjW7N3k5USfSFj9g1l931V+IkSZVdbKbxKX/qnb2spCC
aGKhGW1d4FbzJeR2QJRRNfjgISzekRiZK4HKufq9NOUZzxhP7o29uYOFVl4Ffdcu
N4WxWcKnswxHGktC0DV3i8bNdg/gh5M/CRZOY1v3OcRJoVKjUO0r6xn7InGRjBDg
UMW0LEfqVYhfwW/VSAaGFRd5buyE2oz8NfiVt/5HvAJhu/ZmYhrbuXXKUpn54ZKk
peOTyI7Rhg16bFFZLEs3hQf29NIC5AwGnSGqW5zM2f0/DaI9/yTOMeapHLWTfGxw
kN9h6/Erjn99lb04DRAFUgagi4rHoCB8sQvvvdXwZDx4BEwjo3fJ326fezofeeoS
Sg+VLC+6ZtXQpQvYC6xY9bDYlveLaDvNE/QNOK2ZQxwLZXnmCa9c4RP/1DtpHgFz
SY0E73NHHM3pIuf2VVVvyoZSdsySY59MkJK3qcl+1Pg1kS1QFL3YGEhs6UPjNTNN
xSWVtTBLtFj8wfuSP5ORSHD7UftWegcdTXEpj0fbXKSxB7czdJD7vor8DPCwlZpj
jQPSUnvQe6W8tCBXgMFNcvvEhXUIEuFdHbmXHrFmZrQuULa/8GBl1jwHP/jMn2Nl
9UrqAgfpTak+vUlvtXF/KGJX9yJz/g9Q0VzKyPOiHaxroI19uF0beGVuS3TjAIpX
BCVav91W5Bh9UtWAZ31DZR79uRBK9dIDIXFBAyn7x7b26EnOxpPBVFYnc8WAx5t9
cuIIWIs7eciSy7wg7R6ZEuXlQh9O7wifjjM03KAt3IWHXdwcJ0fvV5JpMUIJWIAE
8CUChTkqPhNgf3X0+z29VL0E+SXs3NEvs2jaaBisOS11HL+TR09HJGJX1k1SjRyN
a4l3d7eTahbgecoG1p9K59kdKeDpnkYiBmq2mJb28HsSAonpUmQZ6A7UTkeUBqiN
S9LsByaGq7lWujAjWFmIOxaefCImPbslGUJ+KzEi7ZOsShCO74VCkLRqcmJjPqTz
iIKmRzQ2fGrLXNR+/YitgVy5ph5JIMHEVY6oLr4b/nB/hMJHenJ/G+c0/bNok3ZG
sgiMuL7jsBCbo/AG81ykc9hHykC/4QJrjyBHibzprc/Ha81y5tGZ61YDVw++uxBc
8eHrJnRs3YJqz/dh7900cZfWSITo03/EGY4FDjof6Agh8CmrOrvrdo1VW0XN8ILe
X+ISQ1+YX1aJaaTe+A4YDibRaDhpmNyS78BwtxExVCvmHw/pPzuXm5OD8na1B6WA
E2aQTlCxQ633Nx7RP5AaqemGjFkQvFXJaWKV/K6xjkVa3AzxjtwjRif8F+B66YRm
DwBbS/C+FcCsFKH81+QpcgUA7XQMcO6i3gw5XGFppukWmoVCEjs5Qj96clVHN87U
keDoMMkOOjEs0TOF27zKHijgecCD2oBB1mXLnplFfi841mirOSGIOG0OfJrH6es4
pqUkGqmtVxqg5NmW4LeY/0xt29FvXQQzSgwxvc3WLXXamnyhXS5FyZpSVubsyAK5
FKQliYbkIzlsQ6iUbkCqE6iZ43N4nCc9535IPupL15nkGXsmlcx7JvDZN0RlAMNT
v4G8/VvKWmk2X8CIiImaUs0M7pkvBd4+MNdQwxfd0Q0EW0s1y+K4CaegY+YiPb82
K9+OyEDe6ufm9YQZdgDZQ5+W6mXArXuepD8bQSaC1DOLJgsdnynHwxB7GEwtAyIU
+RAa+s2V+aBk0ed0GI58mkNjuH0Yjla3myVi2oL2HjClAEWoJl/wbqCvE/dIOxCK
at9ypMF3PCVBXok9ZTb2KRF1Z9cO7g9NhPogIEl0ADs13YuDRuYKXBkGy0kx/2lK
GpmM6bu4GVB14OtMcARGdJzNyMnt2wjDVYtWKav1L5yIt8X7qDVzPkX0Kso4rwfg
QxkDSG1PAkAQqljkK4m9Vdo1kzX118+Igknvx3GuX5kM3agun5Jqrsb2lt6xp1n1
MEpEvVlo+2KvgFTDiwBshkuKFNdcM+3U7whdx+w1gQKjuEW4zC/dMBn4bJFPtVv1
un8nbU3p79ml/OlwyhCTP6pdAyOu5QIYEuTO2o89LzYeKes5lCV1c8v+MjnEY1Wd
5jPHpUpP+UT5ItPans10BMY9ETkLNlXPnhk4hF2Y57Cnr7ucFXK/o05+llFCuqBD
eoSX1K1drNfo0TxP9AiJdenU2LP/ZA+45KCfoiaS4x25EXlhFbaElYagTCFZKr4M
v0NYqf+qoLZKrGODcItrqMzXtDjek9cdvprNcdbabCsCk4QhsyhTZnjIO9CmRNkA
bgiXgSeNX66ZF2uaDpmc1PlPzn19jUzJmosHvxbZrEzDUJkMJtsOZb4isabMQ5MS
HiNPAjFLnx0jb8E6Ami9129DO7IzDtpDWcINsFG4Ludc/y5XygYzEcvA201NpFuH
QD+jMix3mPIQkd9LDIO/u9Wt4Ea0im14fNRjodD4KupuLoS3ut4vBh0mpr5aVY6x
u8NjQJ+bkvuMmNFZJefHVlXOSFpS4XyR04EKvzHepqtYK/Z0H9fookwmFZ1mVKMH
/Niy+hT/a2ZZhQ/LJhJmsXCC5i7HgTM9ym/YD4DTzH+gGDN3LGrmS6dEWur/yQiZ
wx4zhvqT4YQFkzMxGzz2lVb6rAlcs0q5S3EUFMaKcoaKQqzljin+29FZvnTF14w4
t8bdyFWIBCzBfKvunDraHUqIdu0W00VuZZzH1Ud1RtTcF6e4ana4awqcXWp4KVHv
lKH5ZPEARWCNlVub+WQl0hzposhf9phbCK1JTDX4YrQ+7EsuKQ8F+z5lKBnIXeil
2ifWodc41/LrauBvIImTnY3BNvCBBDPqV/fJkrmexfDyAjQ1SsA4MYVFh8yGFFDc
SrUT2tt/pPW97Z1nQUwDT45OCWIEU4LPp3jsrsGgy8ohBKUPmsGy9py4zccyKX8Y
oR0aQgqf42eV9foGDPPmY6fV3ErjESTHsKZuCIuMIl7vAbVM7lWiZhiHCHuakL0H
rRsiLqMEQYKS/5fRr3cix/OWl1+/adUREvk/WT06LeyEH1PLcZ34dbC1JPyZ98MY
6KPjozRL8s4Ig3QtoiVkzI3TG1iJBbCDhE0l39uYCkCMh1bPEy20ULZTo99A9NUu
eYigtYxAVnp3ftzb4bR9+qAMCHGpV55hYabkGrqCgjrOLwxUxWS2iOtyBhUwDu9/
WORgBiGbYyua3vCfyuZz3A5xV7cCtDfeQM1oxIXWUXBBqg1sPmzM+2p4C5fUgr4l
BJEIqeVYCVBL/vj/9bGzbU5yRkd3iUyOK1auT7nN0aymqmNGgc8UL7Hmf/mmTKVa
jN5k2RDyMaGuJbrbvocpkG2JdS1IMShYuHIm4KsuG0pEVNa2IXdTZOXC3UYkWA6C
hJd74jzbBcBPMEJWyINlFmrN3IjRXHUFi6uH3eFmQDlZjok+w5TKwVnCCRPBGqL3
BPjzTJADFrEQg1i00IhYAusOB0HRwm8eB4uzm4x3HAt88u+q+alMubJjmIgp/zZt
zcsCcpxRX2HNeOMsoGpNII8JL+gmY96Ecpz9uehXFEqlbcc0xHpIqb9vigG7BKg7
ybK4oCMvdQ+NHbrTir2g+OKMMJMWNDs4lCFITnUe2EifphqDLj5bRafC8QpCjYpo
CQhbRtCc3z31aOl5c6ab+POHiUtVg11SOxQ6E06SDzxUOzBd/Hb+2h8+xN/Yibv9
hpmlIu0iwkHNHvSk/m6QdDV/Gc1MQl7DeYKdiKhAHMcGqhO3zwqpP+2aygSFquI6
YNDHiFIWMaZrLyvEygBH39TRUEzGQMye5F8QjroX97MAkw6meGa76Wx/0wVqCs0M
Ogn4TviuMlrJPS75va461TzNrxAidDvqIXda1sb8X26j9mPgCqxB9hkrn5scBGbO
C7UPCWFW2qX/FMq6wGtwK+lXaUgm0q1fyu80RkXmS2q1sUvHm97Yik+LFEEPR3VH
1/T4dC9AjhNcOQs5NL7eBTyoZon8jJR7+WulK8bw+GvoL1JI+oaadnzNb+jTAb5l
jUF5QjWBUpZ47ozJ3d6b+tH2lKMgUevO63m2vc2+P67F1DVJ/M4dic7iscTaL/CQ
WHowYDY9JqFR7BmJYX6REQUujIIxeBE0Dl10vRlDnugpnrKOY97Q6/KlAR6vCyaN
spagmcrBPSpKQzkX9puR1VdwATpJiP9Ki5NpWPq4eh/o3IiiGn3IrVUmyNBxGlxe
0ZmdWrfXjFlbcv/gLz10uzRvwAh4J93TeXgRedX56gAGZA2iQDg6d568RUZ4ghQy
/YQtON9qyydAzRHWllt87S2GlN4/7J491p+LYHCn0LMCKJEmxnhEVgKQSmAdCQZz
72Iq3tIUyaN4i3QA26kFuSOjxayhtxET9uAWhIC61Rx/vafxX4X/WNe2bxLAHivT
p530otXE5MAMWwvsdbYSynZ5V77lotKdpUY3CubuTuBMyvhycBhx6xpZnvl5piWx
2YOnpJHX3W6RNY5p4GqLC2vGQDEAxwtpYWez/a+tqzN9tVBTINhfDcvWzuWtBY9/
nr3Dh+GSiwFXJoJWaBYpJrmo4M8GOVWNGNGN5PI3HSovPFHD3EyEQu5oUF0BSLGN
fTy/op10yuo5IsXL5Gp2yLwN+TB5P6Ffv1nKK6pWp+ber00Bn1yIyKfMZpWqwCw0
tIEM18GXeYnVE9bGtlkfSM8xf2KU5BHsEmzle4ckKxIh40toRBn/5eJlfZTQL65Z
15I3wXGZ94eW6ZXdM9tSyYj0lr+l0rfOSwjLoAf2QHrVhYt/KOfxL5jMfCh/xnur
DrF7PwHo49/SfzEaPPyf4ATQRuA/KKsmFXonlZyMKdaGfUTZajDvrOycZCGbhVgu
3+QhkgELG9muPYHU3QgEGPYauiK4orFP73ez6k8Q+UQMItpr/BXZ6Pr4MT1Q9730
XkAtLlzmttev3KnCFij/01Q/WE2v746IRFbVirjgrCXCfFOF/ipN0mG8MPY+LQ/X
9l6Ccgx2EUqgTmwWYrEGnE2eplegWndtrvo9OCSPq7dXJ9O1Q6GhS8pOJKYt71km
uqwQNNTDNExhi3Y89R208Ejn10DeimMghLdguPTDFmGEsQmu0l79n2pSdmC+DqGe
EHiRqjczchksH6dYoCsYrUJEiti/ijt6iI2zGHH9vqwMB6DW/Z/jqk4ZUAorMr2l
ylkxlCWTnYe9kYNJfkoaAo+ni4A3aGm7LeHmfCrSNAdPDejpAMVY+moUmi6W7Mdx
69M741eNJSNyN/XDjYX+c8sottZLjsdtCt2HNgQayh9S155dNfkI+DFBLqv1FM7q
GKDCBS9FIXNwF/O3qIrvAdqp0HbgD5DcbTFWm40UgEf0EsOJC/p+p/8NLw9v1riV
kGa0rlFp1J/LCS0uhHcfub8vXIQFI17hiE0f9oApNnxYp8jRr3EOFTLmGiXSiu/Q
EGprciVs/Lpig1onG6khWflGkInEaCLGgJhZgGbNpiBCV2CKE4EOPCR9SA8QM8Pf
jPiRKJSmE2cfIOvXaQcUVlFYN2nQJPDva8q25M+cm1iMpCmu9NxS8EK5msE+Tvtd
h1k8kGw+2dInWwoXwvVX9MV+PFnwhz/NOX0GJhbltEN2EtI+otAEQL4XP44ouWRT
pRcuy/SFuX5Hd9SlP4tckjKHp4mqeOAsqUy7XrOgeJFI9bkiPjRwv41ZK4n+Xj7L
OqjVHEsvRkz5MNtgli3NoJj+4VHFKs8UPM0W7jGfN2cqhor1RHw992tCT13Y/RVw
6Nv4/2AS4ynjcB9mEqFt/dWAGgjdSJvgQK4+HSZ1xk/Qf6kuwv9Q2+lAgewJyHT7
JR4GKnGLAmtU9HVykNiXOJ9SVewLEpC+6Hl0/HciSs1RRsf00vmzk6mIMZTh+m/U
tP79hRVK2C4mDWwdqYuN7+gI7WiH7xstqFSJuHJnYKdJj7c61YbswyJ2kTQCrNA/
IncFDzyeA6jiL4DFk5mUSmMxiMCMIMtDHwYSrsF9XY6Ivxlrg9O8tGFi5BvPFZ6R
Vhv6qpTpOfgeVPkbQ9QzG9gM4nDypUVLwF3H5RyVbU/+ckUWMBXucVCRROHbsP2V
5J7gB+TluGMyJ5nNpjat9VK4fcJ/mq7byW1wAb60YZkH3m6tqxycUFi/kb+qdyb/
2R0ExBrpXzxsU3DgMc9saZhWrhIzGfhuz3rNUVF3jlIKtdDi5HZv5H9rSV/Ezpcy
sWxEQtTfh3vTb16FMK3L1pjAoTIL3cEaj8krgfDvJjzWRwGbS+VH33vuL/LxqqGJ
YKlz9hdZbdvXHcSYZWIfkcMayZPaH++HjW2Zf/J99UeUjBRIFNngkiqp2zJa02XS
eF9rRcMGGbCjokqf6YdAEAnHU/K5xJCKfBKLLEMH4fTNf9LJrIMBjdFvLkFTwB5d
EF/GpMg2Evz5RSt4Nu/QgKrx2x8p5e1auzTdFrKnis2gUSZqlxZeJnxi8k0TbgWv
kuwUC5gcew3Mej6tC8XkeoZNhV8+kpbuylCr/G63JZk64dQAo4G5GyErbh7T9xPi
rGOcWWbhAISStkHAhvZ0Iedraun8/N4DOs6/KCdmHsyLUe/mRfv7+w9lXjSeMefM
xeMz0NiI3+VkVYMcPwI7HmxCVWkxgHLFodmN1OJ3sfQvhFATu3ricn6Jp951WFvJ
zk9aqbI9ztnut/+q8Mni4PZO9fS1crScmB61yNhDT6YkIBqBOLnVZWIKVLD3EYYr
DGNlHQ7CGw2/12CBhAGD8o+pMt8GtvJHeuG1EdlUcD5mCtlBfftQ90vIPB7ZsG49
1oaTeJaIBnXaF15EnYL7d72Pebit73e/qrgKHNyd68bx5R0QZc7rAVKFFus92Nn9
N4yC/ux/6YuxWuS5qPV0qpB4ytATtRuIO3ZFbsE05jLnGrsKqpY/0RqbXFz6FLRT
To52tWQIHLaNZd/+q9jabItWSFkNzr5Y4MSnMOW2ibqu5Hjdv8Hntw4TF6ELSAxl
15D2BaBdKxYv/n7srYdHeh28FjRVntoNicVZZwNdgxFH0w1jiNwTKS6w8pWpPW5D
Ui124BPbJMdE6yi4XZ/+6qGxXURYXdihSIz4zSXJcO+XXEKMP9i8dybqQ532aNMZ
mjcxS0KMqapG/HElymc7Y6JWJ3/fGJHTytmtBqpIDoCyQjCX1Rf6qSqxvfuPjPi/
DvrWsorBxCnfj/AmPDuR3RzibCT2DnAT+NmBgD7EMNnouILjriInB+dpObr8cWYW
4QUdk27Lt3VxwyfHbUDLHVTRyWlU7NlHxzcbxqzb+2HhxRzVvcKu6X3SIou8VICp
SXhhC/4o4wPw0zsH6xobsjZPmAIwsDlKDqN96+1DPiJbmHUWD/i1UrMbaNe+9uUe
CJU/deOJWF0qRvj+afETYR1girJEMZRKF27002ekew65Svea1XujcBDR1nfqpu3F
9snV8CP0LlCn4zURo1dFdXA3vmpPOz7/LaHR0UunivGBh7wShvGZ+1s6V3DjkUXC
dmbuRSG6ydnJgcMzHY569qH+bhkYI2pbDy6e0pYNIFj5qsM1hFdNTpoN1cn0hzrc
3vWZB2/3nBpnoSgy3wTYHnTxTtHxb4YCUb7FCXEOOkQ9y3ZdY4pS9ntWS357eA1S
Ynt2O3bGzYSnWkdsIhOva2Y5qZMMxIOn+kbqoNyRk3RIHcBV8xXD9Yb8zNXmZH9v
rAwIP78l2Tws365jIlyEulMDpKNTgx5rjkZgIDrbsYLEtsfDK03WlicG40RqzzC2
wTsdEOUmT1jxmBEVO8/q4v4b5H0e+b3PuqIqZ1aEqbvQdm4AUxcAqBSQv4welkvs
X5E7xpqTcm9VKW/Kz2YrhSjGTXHDVdMgRt4kgJJYt8E+CsE8mRiYqUggAkq8wCr/
25B9BELQ1vkEGYxz1qC/l8yxP5ExZHY9u2GBVwPTmVx7h6T8RJZg8Sk4YJCQDyKz
sBhl5x2YGVVQl3Y24/p2Au80Y6APKOQFXlxM+PMzt2s9AUcIjLHL9LGGkQ7ganGZ
uFNIYmtgN+4Ti7VbVzx9lfwVGSyX4mnmwEW+j8xenxlIIs2cd0C6JTioiZVK5zuT
oiAuTTBNQw84PtO47IK2jPNeIkAxd7Qr0F0A5RUXCDte1dx+HLPRcyPM8rEYw8QQ
Zfcptd6B0lOGOA+HwcQlDRq3TVG9hWvQY3uuXLyTaODFX8lFA7H6FWsuaLm5RwpE
VDRO6NZ3xQDesK6gI19WK8CAc016EGS9CSLt8j7RexV0tYewXhrO1q5gDcVaBGxV
9H5LKUNAnDU0b5hx3kFGWFU6zt/ZpYRA5ee7/MphwYqICikuW6/MW/u6MjuymQbY
DfhVuPj6KZJip3tUjfbNbr+NxSVsbyuKzq1BQxADX4Pgggms6MzTbkdF9AZf6s7j
KSYQM94ZHhFfHeoVcskQLHW8T0UeYYDYFBMuGZYOBT61AUca+nLXjd3Fsb5VXMcp
JP/LScjOSu92yGKPcJB+ASp0MhhjT2QDkvo0CjkYlYAaZ9kCLw2QuflywiHY+XzT
7u0qRF86t263oH343BPLjTXKtjxJjrp+9bCmIvgzEzKxznVJdfpwyVE1kedX7pEY
JeGNoopj/+e5ZuQnkK7ta/4D+1PDulTO/2+uuF4vZR3gt/iX+GLnwR2qY+BbRf/T
UD8fSQjZmPqmDB5cBnDHLwfzTNsbOHhcgKooykJKIdqsc5awHXC84EGIL/oW/c4w
y2F8LRVKPtyTl+XtGz8F9ddppjw2e5Z7SiHP3hnhIytnOgwt6K5DS4BhYR9M6SyM
qNHD5pEKWY7DBj0A9GM6wBL4aJ0HwxMTKUcSomQEpZVL1oAa+8jeG/yT5QBfwNoY
7V3wEoYto2r2enFhVDQHG3lWU4SFQZXNqYvC4X+6Q2JLs0lBQ+txc6HHZtvHFweH
xgJiVW8HQUaOhM64EZ0mY2v+eXJOUwFiqIE6EKsCMIJ8o06ghjWLhaiu+UfG3V52
L/KpmmQpRnuwvtOWCaZ0h8XH/X8lA00/IHXOv3u7mW+z8hPd2LMEND/CyUGCz1Jl
mpTH9UlO3xn0GzW9UFggKYNIHkpUGvnhM71zoJH5eheXGnMx1YT/09L4nV3nwPv9
npBJkvdgmS+u8IwBw0EsefvpCg7p5akFpLaM3l2IakQdr4X0HVKw30avkX1EnMIn
kyeG8mHZnUR30PHqr4ZUmQ6G1xJf/OHG8MgT2CN/4xatqnrOvdv3oUrKQo0DmNSp
fyecVUMjub9WsIwoO4rcAL/oFhaNoMUnmgpRFKz1DLR3RLoplfvJnPB0MAZLF5Sb
57U3AYaJQVZt7jansMlcY2TBzK52IgbsKeCt7q7A4YudDMAKYz6dlEM8hNcUE5gx
6hUeM7npe3MwCZkIOr5Kto6nP5T1ZkWjrL5zvlGUWEuowS1pFUY1vWpi/4BgVzY3
6xZ3FLG5nymd4KMvKO5yZUo8LcZHKHo/Hlr2iZlcZPgFBMynUYQtOsJ6JUlMhFva
5OV33YsgTCiLM3YyUM0R1klWSL1T8/t9WvukOlXk3RYmqEBzXyoOV3WNLKFTMnzJ
fTRxfhQsZMnO+XTpj895uVrs5m+CeEj6Ud26u9c4nlE6JfdrJyr2Srz5KHuP31UY
DT7uXxe2xC1svtJrtOvRLRF3n3GW3T7Ioau32/qT1tLGk2v8GWHzeXvPhcWF8+Ek
1CO+ruZWvQMg+9e+IYFZmI5kpwRDvy7W5YlAlhV6t6JJJ4C5ztSG2qISO5eYhN7T
0JBhI2M//1O5M/hCECuCPJu96FzF5ak+7v8S7LFUhEUBVq7K46ycWrbhivwRGDBu
UAr/wIN/puKiNLq3wd/sDLuKgs4TKIqqZy+WGH1H6HPuk9xDtkobm3UDljE4NZAF
pZzeH5V/nCqYFI4+DpAZq4H2tkQuFXFNItj4fcnu/hpm27SV5O/CuXlB2zhkn4K2
mfwAQomyO3EgOFe2fAkGzBUR3lATkBQsp17ye6lILW2hCuPoohBjJJBx3ns6YLdJ
Y+4DvKX1dmtR78Fsh77TsoFyK3h8tUsIgF1UBsdNTrjaUiXEXjD0ib0SxQ9v7YeT
QJsylcl7VKQswOnpE8z/FkVP8RLMygd6d87YOLFQqTJZk3P8lz6iLVWbiTxvRX4J
U35ANBcuWitQuluWISjDntb0P5FhV6E7UutU/guqUHhld8VWBLKZUoAP0hvnlHXo
0XC/pCTMfI0xu96YyLXvEOea9RT/3AH9upgGz3E36fKY92RPxGAFjci4+EC+WUfa
L5MX+ZTFecsKIPLegLRl0TUw4gBUfWTMSFxX6KjTcojO1qDWWptrrPzjcyEpoQ0p
91C/7bBphN+sgRk45xq771DymvuPQYbvhXYmfUiOhXOSWNcZgyB8aqbSVPMoRF5R
orgLk3XT8eP62BeVUHL3jvu/1BE4d+hqKK7rixNKMuQK5YMGFyb+ScNxFsBauedQ
gTbgVn3zx3/i5wJGv0jhpsm1vbbU0eRKfneDCYK6uWDNCOvx0tLugoHDuLOOR6Us
VkES+cPX2mOAdm1oEEeVCxpbgttgSirbOXvXLmJ8DS3H/LDn4HRlX4udshrlUue8
L79vJOCz2ttBDmdhZ42Arvs2O6dS9gGBhtW93JhiUWo5E4NrFWkK9nb4AwWS8hbB
o60XfCTTfq+CVH5A3tP6ExeQkc1BJU9bMDqkbO/+2nFpKzc8DxpuoIpMd2flw7PC
WnE+haGOPSXfGaO4m8gFgle1QkQJ8EV3snP7ZZAeBWkgYjg3At1DTbHa/vCbLijj
cGlQrHiHfnQypR1ryLf3oZjELvYLKw+NSPTPklm9AqbhqIpHgSdVb409S4CwuU2I
1+qOonOJX3sj58HNq98C/DOkbn8ue7ywEjzhOXwRLEkIpEuc+H/tBd7eXLRFimBj
+c+OosT//DusxZwtjiClSnh2wKXTYQOz2IhDa5GhiTXRplk4lJm4+/fYjQx+neiU
ao3CcxBDOgSgobe92tveBq+Ryng5l5K5xTWrDIfzqSdxTagN8IMmaBgDlLE6svCP
45xKD+llOFuGuPS0kp6q7etiRsmSnRluQN4SsRLP1HX1M89QT4sJ7gVTR42ByFgC
wV+H4KksGQGSV9FyNB/GWAHf6JnEkGP+pNRXV/fUfbJPY19uvTY+miZ0Um1PDGmv
E8yZonre1iJLQGrVf94Dh4iguvDbYzsZGSHOGPvR2O7czffbv+0IY5mciwSU01i7
OQRn+IF04SWYbavytWj964l/2vfQN24+sMDkbRF1EkWgHawDtWv4/EgkEaIm2p6i
cXZHWR22BxGj7t8KeZT6M5XOlogQLXl+K02br3eLhY7a2i4S5MPXJqoO164H72WV
9hB6U8g4tf/Q4rVLFp5PBI8IvUS9S5uG0XIPQWaEzSVSrlmBCtRNUGXSwv/kXZY4
vlZCbdtkZzR0j2SSJ2qVno35MAT7rKHYJvv9mslcxqjha4fFysDCWLnd4u4uQ8Us
5qDtDBZsofvIcGKJ4mmp/8HacEx98sbwysLcSD+HtUiDA6zudkkmGJdCrpywAd6p
KjngqHRZNrR512s/x+REu4riVJwvJyO67xD+XDdXoYwRV9QZ9IE2l6lEwQdtPT1e
5ZUwHbFydAWftna1LDbkIWcKq+ShVQHLtTlipdLj2iaZmvCioeSNW5Lb4FS1jMx1
KRY4OmQHUS2DYKQO2+vVJK13UsIPrpyZXxQXra4gQoMLVBhzjNgzKxGlhmb8TmDF
ukKuYisXaucpZy3z7K7lZliANwX3EbV9gp3UTSj7Ywuk0UZrqU63vDb9YtgLcC1U
qSN9MpF1r8zkO11e+TBVW0dwge1OLhUi+kNTQ1Sunc+zM0OmXwPBK3Cz6V4+ndjs
bY66bYLRRKf2aIbZHC1dJb1mBTid/DrCvvqYa8tJwMVYYCjopd42PYxF8JG7iQzB
W1mRGHJoOB7a4WoeWpkn9HyaSS9/lEUDOtFlkM8Noi/XoMMOs1DfL9MDtvoOMPnM
yMN27pim8QfOiw4CUIDP3CwkIw2ohlz1gHirMUl+XyEMrI91kcYSSDg+sbxK09x3
tbsY6bIYX7cyJMnNFR/a+Wpoyvqdz1QtarMd+D7Ou9ssDmv+edheLIifBZVj/KdH
JrAXieeevTJyEqK0ByGXrM1KueZbHZ9rCDM3OmQM4X0OGHh8wgIiXhUw+0QFcyGu
gC0aDy4SOzQAHymQ468JkVWFICA28SEHVi1w07jxEvgQay4iWKkM03HAZ2EHHg+/
ct2Xd+q9ga2jzN2Ur5iDrQJ+CivTfBd4jCmT1b5yasuBxuy1yXahWX89R4Yg3KNn
L5COQv7Hk8AYALI2SUOP1wMq3+fgDHTk/oaMTAGTWILhgSnLYEpVE4gItN19tbb0
OvndrfZRFRp9ppL7OVG+MzhPaXiPgDmx8wZffxpSAYnswmedy+DXpAZ4RaB2B/KA
lkPZjPx+taRDuW+jv4dlcOTo90gM/VowV96d453usyMvnTy4qsbuO988m6YC0G79
oZwah3lYfC0a3MW0D85Gcy66GTs1xbALA71Wg16bg6hV0Pnppr5kxulDsphUeUou
acPkSjifALsXg+wY0T7fhC20gdufbrZMDvz2coa/X/ZB3EgOkDo1g9Wg3MVd+sFk
qEa1i5n9IYY/Xrv2brAiobiD+jf68p1KDf2u8dXlXmZ/KYZJhFwH8mFxfS47IMjj
7t45Gw3p8Sr6EtFWP9E/lxG7hIcAj5prEKrqqD9V93aNw/JoTrVA/X5l/zZ35g5n
K8ih9JxfoHLDUK07gULdWTmtSl6e9IBL6uehGqgdJXhz/FQH2Y1lxBFRrcCkVo7M
l5oaNxFBtFo2ZVcWoRsi1kPWtP47ttcV71rdGXytKsnN0PMnPPLQCRpwg8UQujt3
oXY1c2hzAiNHmFj9key4G9M535YGEAgkTVRHVStSMbwmdQrlHg4yV7A3UwtOTBYQ
AhCvF9XMsMIkes3B5MavyXyYV2P1RuUxFgzMFxhFTv2VW/dQK7Mf+PMjbLYjGq3w
n1C4QrDs/Hk0McfWOlavfA68vsqeH9tyOSy7Dd3FLWw2UaClHg8U1sc7XTfVWWN6
iNMk6X5f8Lovh4WXQBxXEF1kknGd8o5yDGxK0nbw0BXVlNY86vYkVpR1XmrA9KKf
e5Xtvm5oAg+2eQaals8S1hMxKNenLPK2nS+i/AO2sbPhrt3B7nR7RdtOsHG9H35K
fr4c1GwWpi9M86svhJTjmeLVvoDTWQ7O1aXIphx1kgYbbgqzvDb1iao6kXEoyGA2
Xd1kQb/naNoVnZcqpIMjyVWjTVfdgnfjJLnBR3qgZK1vanJhFW0iUj3a/oVhmNFD
nz1bZpIwqoX4ShRN1o5/4o3pXFTfIXyQ0L3Q9/PHq+11FvInuspLaxcT+v66YEo8
XswE659PCpoWGUqwdsOv5NEUEFwhA+NZQ/MzVoFkNuNU2uP3jsxgAKN8+co8aDuJ
OU2YTUV0Uaf8oYGmteVP8NGczT/gh8vE9diPz1GDdvvdtBGuXky+QPAujjnX5zQH
fLb/6bDVZXs7R+gRsIHawzNlDfFjMd2+UEEk1KqFLBExqe9OV9rrG5rPElQ0F1zB
PkPM/PZG+iAAXHNF1T/J7a0Jk1MmzO4uC0HbVEZCfmgPvOX4r7f8m+rSNAvjvruk
F57n3EXxTG3vVS9SrRA+972CVW9rJPasrWaaVysRdJtF6qKmMZi1wk/pRV20JR8F
UdltZY4K4ooSL+/gY83XpmETqDlN9CLGATP7SozHVLlQM1vKPCzmQ0JAKeEav8iq
uv3uzcUt9N0jqsUdfbcasP1wqNo8KumS7vuUOzmD/zYhB+NfuzlzOtyFQJRIyWx8
dvMVWVuIUnS1HPRIQJdfXl+K6LTXopBd7QmMgB11byYQcicjzmmpN9stakF8etHR
izLM7KQyZuIb6Cwq6godgekwxMmzD0LueLL9m5zNpoa62MxZVoL57SabBYr24z35
nUaRL5/i/RlzTEuDDxKmOhWx/j7lln/ZKybSo1Qr2WVKW+m4HNx+Qf4sFhgQKXDE
dDdchOr7LLHw0F3HkudBk8MdsIIqlKbJkkVcQR78I3cgmMrGo830bseoE4zZSxN6
GLSVF/P2gRE0ZQUOrS59MlGOn8aENgu/1OHvS+V+ZQj2nPH/vIyMntGXoWy1P8xY
i9GVLMpJaK99ake4v4DLqqnHVzg9bSrwZCK1K4xJlqmqc++tCmpm6BEZQ4R1lZMn
MEZun+6zEvxRStM6SUWQdsgQpJ/pazg+wrtuCMpl54xhT3iPa0KKu1d+6A+Cxso6
+js7NkjSxrp33MxvsTVHSjkLpowgyM5b3sTrhyRXSo9FE21aP+ARB1Xa3f9nXi8y
qxFGpAch69MKsGFW9lvkqVDDPfyo4VPb/1lAuB7gX7bZea2HS5rkaqntrWN+2o+7
E7PJXcSHMe43PoEdygbPUUnW7euHx81zkg0oPemeR2e7v2xHi5epu1LY8Rhghqug
byTYB1U9K8jYsevHHVYewKarAfyi5IQuDWO75GXVWbGvXElA2JBW7nPAy/pxNTsj
FglaYGfS9pqy8Z6vRomfQTmwTubaqZN59NueFcnidUsoGOjGt49VPg5kopzI3hp7
DYr4k4YOOI1/cgw4RG12vH684QLpa07EzWNFhPMNWTuDOKW2PJfy45MzsM78sId/
xZ2/OEY2pa9ZTRnxkFxmiQjImRhwc9lObEpxfzal/9cd64sIXsik7mbbWfJHKL0m
90iOrSDriLALrzqIytQvVEh4Dtb2SYYzc4KPCef6Z837Sj8EB9glr51HbYw/oSv5
aIYL+FY7rcKfVyJUDFvzJZ604jOy5rn8N4BqzMIYkUTXWE3mUKsEqVlTNVAaWFDn
oVXh99KrhEpCmFvZt+VsM1/BB2G76Flxt76U5HbGpQX67jhVhfPmAnNCHG4bESZC
E14WWzyHdB+Tx25jSmagdq9+VcNacCORW2qUaSz1qLIGpUuNHEIrklTQ9J0yaNTz
3arUQGQsvYWxlbisAPBAnCUVjw/chc3RLQb4uunQUOFlg7BkjReljs8X7eUvLmx2
fe3ItdqLxzbJUivUStJJbXpt6sts7TCyRKuWEGx6Pkq22cpLsRF+drjs2iQvF5cb
pwkemH0nb9aSqWcQYhnXnYE/kFuzq14KGuLKGc+VN0Rq5xGaZRO0J01uXmDfXWvL
CF1x85FWlHn9UB8wz8uB9xi4qj5LNny71zZVmSXZ1m6chhpEHgOuC+8OGarRX2xN
oCjahIJzvGDK+xfutpcCRkDPBX74yQ8qSGjZkrTeVQcbuG94ImUfcwnNWE+mBT1W
KkyrCD9MWt3zPqkjQqa3wBr6RJmDumZHiP6ZmA3WG+d/MVtveytlvCl+tZW+LleI
vqdOimkYvi6YYbf9F7rH6TBZc2r6TwDCjIIISdYG4A0RtNmiawKi1CvD0LLi10M8
CX5DOhR4eozU8gwX/yhRfterttiVpGUZlf+BUuOj3Br5X+LHQwYNQqhnCOzeyvOW
KIuD9MbrBlxcQMMgcDUWHD66eDPG+DnLo8l/J03LFTMqHOSuktjdNVmtnqFsG3op
LH++Fn5aljA09Dq1KiYfFCBkU6gKFrlrqrV2q56pvqA6ZSt3Z0fVm4kZnj/TIjrC
merkeZLwgxAgVzadBDjunfKUhfYK0kRTpDPk3FBwgubo+v4rXDiHrVzV9/uDfPuP
/+Yxr0i6i/cCsYJYTWSmqd6HsrahfZ14B/o/Kb1xoApAP7c+LPsjd71oIq5SyFuo
LcLz9PKRlKcP/Jb5DmNnCNl88uxfmLi2Mm9TF5PdrsNYgtqIKWDaInbUFFpcSYhO
R85RvSe1jBywS93TS4iHjTgI/9Ie4NgCr2lrrW0RYTNSyWbwO6wnkg+d8jYjoRXQ
urO1Yrl8ijDCXUN3YjpJsmC+i+wINihT2EIl6hkMbrMKMpIddMFU909QIM9HeHBf
40RJXrulOc1sFfiqVU18SWzh72/dQWE04+78PJ4kGmlQfj5iSrFcZsHybUsc8Agj
2j5rV3Jck1dpidFefX2ZQ/3VuODOuL6S06l2J0JqS2eStlvpmGN2YJ6n/QCVzzmx
P30x9I35RFCiHK6vK0fCSJbKK3VES777kskaRduCUx3BqLhuOSO9kRZGok2WCGyS
10mMTPhJC4PdLoYMpepjYPreWbItu2cB4njSbCD+8njthoXYcjJxSm0u6xshWkZI
cVkBQ1wSmGwTSVppC0Pq4BrtcrqzjZPJGFWRiZBKnN0R4elDIHQIx/FIFVexXaQX
SKMg+lyBETeEtPIpk2bvytFlLG+t1PLcMC5f0bMOw2KxuuIx3pxtol7p16n4MWTS
eSWfbzixZACXKBBkNnRCyqiQpubF9M6Rn8kqSNJnWv814et8Pe3sy9l9tibha04L
lTmcdCA4leTBItvvNCW+cR9XHZtwG8tRcBRZYgc8sox0VpgTvZE/BeqCFOmE+6LR
fqsQzqVT7Ra2HuZKiU3rQ3vtkuoydFqyHJM2dsYT2x0T0t9VoVJVuaBoQ4pyvaAK
XOlH9/mRslunwn0w5Dh6muRURTGYRLz00ZaHhi9JIFvrVFZlGHQFcaxhgKRl0/dE
FOqXup4h/ub38oAHJlu5z4PE9/BLahKTkeTT3qDRST1bFs7BeAo3tyL46xM2HZXc
beSiQ7+qZx/Ti6wgGrgqgIAIOqDNJyI+F2YIIx6EYkMh5akieB3CRBrj8G12sem4
v1fdBumvhWG7olq6+U3FHyBTbVvVQVUuS3njhx+xskYsSYR0HJ2LOziiajmL/7I2
TXoSD4gK2K0JFw7p1t/0pWmopAnL2wvGMRc4iAZfJxdWf+zcsbaJPpzPNLq7tma+
9X02xjP4VOabzBopplOlBkuOfkZJcGmf7BdGeFVD7mlPtU+l1jQ8iCsGmvUvglVX
NIDAk9SbGwYyehbXZjfpugb5WWQWUhJHx3/cQaoFmfvV25qKxHJuLzXBFvDFEnsM
YGooIuljop5b0+YjchsEKMpPyhH/4oYVikbImmhw9NyzaMmpI467VEjqc0cAkyoO
0WK8FsZ0FBDNr3qtevgv7u2o8VFSeJwHOxByMrF7+ZNB6mfMafWt/4qDuuQx0I8q
LfatYKLFTgpEfiZ4WviT0QwdA2JWsDmHep/dwgcT0BKKlCBBTsXC9AdqOA0ID2E7
mIsc5ZBGPQQupCyOqWylphJfESlOeoSGWoMmZ3OAC/yG+M3k2PXtqUD5T/rDsg8h
nSEL5IxutaQa7W7AbOYAOSm9h0KgTUHiTp6h7r95EfgRA0rBBk/vSR6JDeP8g+fm
YGp+V3ENk7dz9+EEPPOyx1Om9FsWW7GiUXQKOBppoadL5vH6nlHZSfCwYLTdaH2d
OyNofh2iqi8UKpDc9fwc9/aqNU3zn/7FeFu5ylPj003KjkZL/6xOl3Tq8Ycpd18K
SD5aY2Cuzd3BMEEmNd6Nfl4UEpxX6jJdpWnuRX8N89Jwu443Vwu9HpEiepcGKSxW
BHn+m86XnrVr2/DNz7soGhyJ5QKwFzOYrNokaMNdGegLTAbGUVkdTR+gPFrO9zll
12kOyIi7qbOMl6GtfYcOkbaDbkKFmZgHPLdOitTdFL3GlR/5KWfKLVTY5i0gYmF4
hhyi0dNpSAOG+HBt0V2l39H3IJ4ske33fJmYmTfc5kAYHxSjQtefzSTKkwc8bGR3
7wGRyEaquCMULYBfck02kC7lXHohyeg9InaYUEOkKvQGXr2BaNt89rxTbrEdLp5t
ENkT4p+lFf4F9ASLqnL9c/DkxYW9WtcsmVYihVUfpCO8I7YXcQrlNoJo6fOWiF7F
N2XYZELbgTdNaJ1dorObgqkUgBXB8lnUCY1J47bjaOkc5miEBar5a8qWPYFG9sW0
u2F5nb5be+ddvblb+mPya2vUF+7yqGczYvFMvaeF1HkTJvas3pnHUN8wGsO15/WO
11lGnRqw5N0piqrgoud+HSI9ax9hGTaF4RfBAUVjxGFZiDR2lnIeiX9/1lsrHdFX
KgDPm04GJwhUuyakGAVl5u2/eF6gOTCAXfq94QHcrvf0tvo7XeThcGKQce6pFDf5
eBDnsC3g4Ik21ZEGIB5OMUEnzlDN0N/C0H6yOIlhmgJ9BO9PfedY4Q4vLlWg+F8y
E6Zowi8D1IaZiv9o6xcUzNm4QjaoPayY+TMX69B7S20U0zzE9JAEiX2mybQ2qo42
jU2NX3fYylyRDCDDgtYt1YKqX+ivsYk1zydngBjugtrt/Q3ljxcyYBWIZTvbxkwo
uoJf4c/yTpO0MjcxGD62sGbTzxYPNX5+YEq/z2GHflivDJAwn5PPxDd1pE8nWTmZ
KCoqQvH9mVnjL58vDjDvoKZ3WxQzOjssX6/aR7dFRUuun51+NJyWr8FAKs1ClEwH
WyB2SOQhq0a4UwqoTXMXGUoMmDXAaB+oRPgZ14I6Ldt8ycpVwZwglFvgE29qhKBo
f9pJzV7EDBCzwHTQH0/ztTfERb3iZ80+ZElRoRQbKmn9OkPSvW8l8kAxfWnUekMQ
mgNmVs3fdZ6mIlZqr4BDVfU324y/y5RbvSyaqMbbpj8ga7lAEXbaTY/C6ZNnBsuT
uTDqkeARQDtUBqUw8ZQs525yPWP3PJ6LzkCu0DVqamLCR3wC1cl2r424gZXLOEt2
qGvOqZ4FyXXIZjZxNhxOjzBnvlkk9MndPe7a9p+FV9CxAYR8RPvMobNawTUSuZjE
0xjkMO7656CK9Pc47xyKXtoGINMJ/Iso3qbtEW0IQ1Mu7kIQ7xEjEn51NSH6tg+3
h4FH9BL21ClGnQJY0kGzc92Zo0zZCC83SRnteHQLX8VuXhDGp1FV8559zSNro61z
N+itinc6HhBcqckWudg9JOPU0D6cywWFUUp+o59Ekw66axPulvhOxAhf1pnJ7KPJ
ugPFW/ESZDc753VCQjNRtZ7CcKNOwMekcz58oua9351pC9gTrLvbudcMc6sH4a6B
TwA4BGpJZryO5/I3YbojurDoV5xw6m3hYRTkTMuFSc/f3YNaoKnS+IZte3Q/6FTm
EKin5xyH/l5q/EMcqNKT1mPb4YkwUtf5BWJggsCPjtdKg6VCJD3tqCL2UhlbNGLV
KIWQeIf7gLfKtyY3Ut8qJjQZp1ePd6iHhD4jTCQfL3Kw9PTnbdoGMhPIkFtGohos
tZVdp60elQfGyiNX7jdQxblALvFPE3t2gTUYxQMlcVoAH/X5Aq+exZAlIBPoVO6n
PA3ustlstw8rkDMV28oMGKeEZUxADytdLPaB0IP9wRULc5WIZlrjXHQIE7GzprlA
e1qkdP1Rp7gJlcXsjEjM1AfpzZNyjqLojcLmiig/bwyD6kxF/6u3OsrFbKsY7Vmn
7C1w4cXyeoJuaqhxdHzUWgOscdUw/2YtAzYcS+n455muSJY2m5BjMVfPPw8pAwrD
psSy7x0i/eccX/gzUJ0RPN9Mqib+OW0YwpGjDCNhLrf3ieLG1wBXfAA1JkWgQnkm
xU2PnNGucpeQGMv5rDO0xqcqvMk3GJcF7DX0D/1gXO4mFhiLaFWn84RIjQJCWeLX
Kow25inq6ltHm5Yx1D9VLjkamcd5VZWv8DRmCtv8EU4gWGCtOtN3b8vTusnvgDeT
e0BmBlT4UtNu8oNZxYDsJaVQr7KLtRYhNGY5x/5gWMRf3+tBRq23gYV0h8nNOn2I
vML8+m7q9oeDuzOzDJb41rZLOoMCUl7kYRq4Zx2AlX7aJf5Sxy37m96f7bX0Gahb
EEod9pS8E2i8cz92WLJKDzcCRYkYJ4Dbd35aZsYe0RK4BjzCw0AlZwc9QPOlJTzc
2abaULotqEZBziwP2VxvrJKGYI8Y68n7i3onrAYsFobuINWMpZsn1sM5YwRaBi1L
ZOxh49Ku6jvBc/uKOtRjoc6qxbc6TZ2/KUOpRX7GM+l2D9ccE//QBkNC4o/p95lE
zKVGUf8+BEjuY/aPvGjlxvVT1fIhTvzxw1so30scUI/1kbP+9oJ14Q447NzSnArl
BcxwKdk22NUBptJR1gPjthXrNbh2LaWVV70PVKwpIblHLDVMAjDiyApkyqMqDWpO
tacYmR0GJd++/B34u2P7ecp0JIbXI4zlI/nWtjjtzNbrpZsdxCDXCHOw2NyQ3uLP
+Sh5sEBh4j64wlc10410tVV8Up8SN7vmsrUZWk0dODTkMLumMA/AmGTmwGd3PJuX
RjedmPYkL+MWKay5REnQppPtebTxBydVcafRF2yWd4jHZruDBhkswctQeKQYW9rk
rm0D8p66GNigAzYvTjhsuVr7T3eLJwg1/JQMZLu20qQbkX9Ie/6zOUrUq3hThMzb
MatF2+3rKBo4saob7eg6oA8iEPtFVIe8v33lPB4rXb7osPorWP9HQ6m7jFFW9Gif
G6wFArxbV+ll5qtOqgIGyOlNnmMWTkP61591JIx/k4IxwhIeEHUEY61qPK8HOSsv
p4+VuYyiYjHN7PHFNgHHHEjxS4vz08Fbf4HeiYDPhDDldZ218WgdTQz26tmdKhsX
9fSj2HgTKp1xyhfqWlzaLSyZAfhUrcUGnme4JEjFHT57xKLygUWxYkEHVnL9Rh/o
zb7xSYTz1E96z8Xdgo/QHSAnE9ossjX0KOf0AiI/FJa7N1Wnl4N3NeY7ZHT/SUx3
03TENaqwX0hENK0MTbKVgXAMs9dadm1GbdceTh656NCEaSth7AZnZ/XMBO5zYH9L
oIB6GHthU+4GLIowJPr71xM+grYeLCaOfD9Y0eC1AVbVXUfie50g9gmdKls7M5gV
1RQwCW1HY3Uu+4Ka7O3dXPqdaqOxPhvQFamhVXxs+36oEEpD4ytCazEcRuvG7y4V
/48OEV6FwpzJO/i8SS1crZrRerP99w6HKTG5wc2NvSMCNSAD02dL6pxTVZP3eYPd
slAWoe2S0+3oFk9QWiJupGSo70XoFIAnf/ZbnMTP3fJuOvAb+LoBgK53dNAalUg5
resoWxe1hhEE+q7LrOpA2nPMRWKUlbzagzBjVRsM+b7PVTgHVpdPpNsMGhXqq9Do
0htstPh6ojbMlUSR8MU41nwdE86QYKikG3GoFx757+eIFFCoGptslRORT0lVTxA3
9JXluDcCL2XMu05jCwJGBDdDf0Fy85BXPhESr0Aa+UW7ROgX3DnWzdbNbCx8qVk9
MYL7isSGNm9qTNMroK9iWWn0l4PhYlXWR1k1Gcw6INTA0SmgU6fY4KuiVh2OKmeS
oSM8UhI4WtAXEhJzrmvnygAImA3Hp50ski9R/XxcGTA8ZhxWgc23ibjMucH8qPns
VtOpQ3jX4cqwLoXfrV98vO7nJrNSeJzZ+tQy8DOFBJgx7cp6KZh+yirrpqOpMHy5
Sp8spQ3BAyGW10KI/hOYlQRjMoSLBaGJqQDBc4jADK6ftqAV/qmvBWxxH/a8FKN3
tVXJ/gyqKl4CaRWKeoSQXJKHjr8ahNZJqTWS2tHKJjoYhxfwP5Rp/OsgEAUdZ2+x
LToCXhzfjgSIYfUxaLKBObaVNLR5XC6UubjvRcq4TsqwCX+UOqSXQZDWVni2FrdE
kmWCqxJG2Iu/xUxJtJMfu6IPsA4r0oVqr2ObdRMVe32HPswnY8o0lwCDwUkTN0XJ
7Pj2fI74R3CGDzbYW8h8vBW5PUpqyGR50dYLRymZE5FHjQJ0YcJDp76iNpTNqj16
tpCHHo5ZWWquyTptKFk+60pg/FiYEr6DoHRWhZYJgXu7ZUFbSAXjCRFZfZTBOQ8R
N0hTBlT2m1K6qZWoCU5CKbfC02yYOHlPGvw6d9yWY0nzpA7L76ubruTsQneNeYDB
IMIKAmI6uTQAiPzQyTWlmgDRkCZEoeQqzaJPdM8csmK+qU+ckK96eS+INmfkBBQu
mykKOuJkQCNRSJ/3JRYcvYSj0YIrPYF++B8qwB5x63Ii/hJhTweytFwt32fdxFqg
W0yXNCX15HBs9zr222Kne3854EHdV9eTG/D0CElL+4SfyCn/fAPgGvPOAM+BOuGB
XC8PPia7bEWq/Zptu+I2r9GY8H0+fEBI1gW4PGwL+noqSoTrPQQp0qCTGnE106p2
9eBdR3i8u5JjpiAsFkP05lJabIu7aFYBXuaINJyU+L+lLK3dUHX7d6BJFxOa5LxZ
ou8mKtnpkaGFrEKWH0SRjlzBbcAu72ikUO6rEqZNtB8u9l0oYI4ABez1o38GdGHi
x1FYoPL6jWG/mecKXqTRidYsQgf97pDSUgvpG2ts/nuMUtPCF3OgkNq3hw1zYoMK
l3JDHsxVs2tPYbdICSCTr2MgZqPzrSv8gXIvBwMDofHvQ4McmAWzWc74jXN55BZp
PlvybRbg3KfYiX0g1HvJ8mLwVHnZk2AGiX/YfYqx9uEs7GMn6QBNaZmgl3dR67+0
5yuH9nKGjkvt/W7ytUQQoYYSh+pL9aioDL9JcJwYD+5pMLta/dZaZI2vCtMHzMSb
CBeajcoenidDbli8j0S4hQKABcu9KVI6RJqV83vefaF8LSsytAMviyuzm3/8pfqh
G/O+aSjDS0fvXxn9TYsHHxTXkSu/zTIOLd51lqVEstC9TpyfUs11Yr6PQh70S0lM
35wXbc2nG/L9iYAVCtE1P3VGC5MDsVG9xfF6SZX9MOa+8gOcypyjWpz6jJi+vjNU
UyrHrST9oi7WhK4JPuXrLBIhpSpOairGyX2sdWl6Me9FIY2Y3rpUzzxmrzp4rP7T
cmO44AOlB/QLxYu/8uw59bVFkHtpjm6I8HqmyBWCsFtp6M3laC1QFrTkPyfsPmQ5
mROd5TjHWugwC1N1ZtcfKxp495z4AZpBWx5EOwiXjAggU20yGinkHQfzo+WR0tsh
2M1fSomSB7/JVNl4Fpi2NuC6nxvf8YRWaqC6A20qOs2sGDJqOGgTXqg97cMPrLki
jFB0n7zRRZKlxLy+vfGoDv1GtZGeg2bXZNkIlyBjXpHDfD+KN4klrq2eHLLDlf0T
MxskaFAvesTYCWx60rOoOmvV1jGzCy9/woIv+zZ5/KE0OqjOFXl0GDP9Id2H8uHZ
Q20afh6PbEyXD4Avrd9OwqbZo9GDdKxWBxMGhH5irmITHoiTamLYpbQ/sQ+HZIq2
ux/iSZu9UEW9XUu6lkTomVrYcYN4Y/Baal/iBPOiHWCoN0bs7x7OW9q1FXkTBnNE
9sHvG4J5FCMXG/ICp+Y9H9zVv58HxlRf06NPgnPZZ9106lqJwEcJluWLc+aqQheo
sJNbi71KK8oVeCM78ztrR3WFNxzyJT8R/ywIRY46ydM2DVufK9cwYdE6B3qRCEx3
FDK2b/zt4g9AgpQ+t0EQDoItfiMJNjbbCKXe23Lv4RkNjOPuKCGeBUrHoLSMs2QG
sAj6vbFoRM7lSf43BZA1hZXEcu1diq7Kc7+s+UKPzPW+o0TY6yLQQhD0mrlXMFuS
PAoeoRLx+QeygWbD9ToTvLvd5mfpgavbKUpzvRhW6/zcH0fMkPLFT76jVZLvfR5H
A8ex+rFooNp1iBgMX/A0KkaBtqBlyC+B5PeqVB1kKdBomrOujgdPtxBhZgSnTjkv
gVKV24jP4I0fqYAr+f7DTia5jTnyglHZBGVvOPwcJjabS24NvpZ0uLgvir4iZ+Iy
lG+CU9/uDYKk+SLM55MdXCLstrkyr3EApVIMkioWcMkK0eVdA7yQiG44jKHA+Ncj
RCpvzk+c8Fj/Hnq9ixaW+nZGPV5o97jHbWePDmqR1IMSKfmh5YO8LCmcdU1emjSg
p1Svwn+XbGqxZODbEPx6I+5UR1A3qvoQLXnHIR1Zmk+eLnYEgofV5cTKTPdT2P4g
W3kuZmrhqUaOu9LBrJbk+jf8GSdnofXsqxYTOoElKfsusnQwbKGLKLbddfQWE/no
F6rpKQjFVOL0GM5kzFFBiJHbpdhr3iPDfyx2Z1HcqtgKmBAXHZ7aaY4FpEDuPi9C
cBnujSU4+MmqEWqZU0/ydQBuS9aXB3VkF2eojxJDiaan9eur2o6WNS3tiAzQOWiB
6K31nopNuKlcUQfRkjv5FjeNB5471fNpWIUI7SvCtQoHo9GYzKPVtVpEovtCv+H2
XLMyX88qio9KC9Yj1IYpaddrtGlOEEbTJUN124TYjKCktFgeZtkJ63eA2dYW7Y8k
PvPLC7wr8SAJlsOu4E5Y3WipvsFoGbvsMXhQiQzsFuFwrIOk8jD7s4mktVsLMel6
1UtcIeqLnss0zYnu3Rezfmv42ZqZ4jytn2lAVNX3c+kpX+IlYKukBUmltcEfQs/y
uzYeMzHXqhOcrne8CVk3L0zw6LPhfwOMAtMW6v48wl3moi0s655yPfbCja47OA8g
cQS35mpnYWXKYc3rw8jL53LKEPPKoTrpdem0TGwjX/RFZf4XtUmMeFDeH7PzM+1l
O9UyTIgqdeEw0kteD7iCvlt/3a+lsG2pBH8fLpHvIRh4QkOJL/VhtE6EtGGbZMo5
bp7di96gnGJd1/dmklVriKySLoR42F4sLouSSPtl2Toav7hY18pGVS2kOyQqJ4b/
bJqnNdrSvR0m0l/KjmB5V31eTwZ1dd9FLpBwATDXlq4gLS2+5tEG/IcFq12O3CeO
OX+rqYhWAtvVWBzcPZ+U8BwD4oyZ8epbLGySXfRyS94wizynE1CR/hW376OnvDev
2X9gOVn2/Er69F6F8BRiuN0kB9UPsQV5yTbJh+31uCFmCLXllBWtLv0OQ18AsAfz
O7G6rZbzma+odsc6Jk5Q1uFSRu933scl4G9J2NOWoWNQvYmr8FxvttKH9ZH1pacB
a6VYYDC0mu0lVzUh6sVccL6vwO8dREZktnu1Qr6FwTydbLVt2aC+dttnihZ40puM
CJWyDDKkjwJs3tutk5BZDLFjkMby/LOlDuRMrKupfXViZ6q8hSd+NZntFDh6tfsG
1egykd+4MimD7iWp0pYJw4k9dPiW9Nzkp0ZR0BzBb0T/5PtnWQOXc6B4jdr8id+a
0fgyewLfJWb6ZmVfSoOtPyMKtO+Euxb2HJlW6zJaNVq5yNFw1b3QDZxpYkayeRsS
Q9A97EXJ/ux0XgoQZkXGqZ7QWIN/MjuUIOqA+AuGzs2ZeNBwjx921SU+oQ2HjkcY
/AqshfivkvzUNIj9CzZzSZ717mqKJjO/mPfXDCB71uKmpPIhRLi4MtU33S3HMCxD
ualiISivdiOu6x3r4nAmihSaiExdSjcyAwa0wzPwpaBfWj+fQNYz05avCC4R/OOB
CbFSqemEywSBxNfYT8R/poqSilGu1IeEE9PDnQaCCeR7gAUg5/DZ/zWrARnypBB0
hhYjQtl9SnrSrIRwkxSY903Z8pUVc/Ip1n0bxUtdOLMyQLzJklO1bPFNUDSR2Crs
KAJiL6L3th5BiMjDV+PL1uE+zUEMve8mk0kQs9p1DesS0JTq+MpuHRZgDdlKk12I
d6O6chcPJA/l6MpDuzpPCOvV/IpEQQsjVXPa7DVhO61a92BhJpG9y1+UJaPS95RF
CbVPlOrow/2j6KVtH8hX0eISiDwQvJWK4vhp0HtxKHuuyDL+SfsODvgX06H6GT9h
ue8Gw4JOz7OOLo4sdXQK1GTOQeYu1Lb5E2IyOmjDD8GajGE3CWkLJeJbJqb90lgM
5xZuIF/fwJJc1PBtPjXMn5aT3Alygwnrn1VfojddWDx7upighP3BOPqXiaF+f6aO
Kyu7pWV+UspcgNJF0lnH6OG9kBMlVIbt8g/eg/387exqEIIw9lcqy3K3cryguJLx
f175Llt7cgyhsgYinsQq4ZbIJ/3UarjIE7zbxycr/mXrU4zXl44F0XoZ4l6YoJJX
zS7MyfECKgRadL55SXOA/FEkwr3demlAcAMWvfKNyHeu5kQU9+/xuFvbmkyPFB/a
e4XK9LgGWBKOpLl3RYf1xBeG1ouTpkbF9ovynWD2RJFotAsLKMIrWEsx1bAjChYA
9dB/tOEsvdMXAFXBCdN/Iu08MHy72uv9acH5TtjstleKr2p+ZXiDfqNWcvsiybVl
zqMZMj+3/WXa8iBRRKED2zl0s9VQBP1JNl3RBb2XvJlPYblLEjwl/XbEP7YfBCAX
hBrXGentaQCc28iUUp09vueIvcwA1X9wYA/c9kyL5lP2uUCyKDC2FWsUMHAVkwC+
FM6w9CborJcqa2a4B7od5nhlhWGfDcoeJBX+LoWdQDa6kLjiSS75kTC0IU+cMCc8
KcWV/5OiHvffagW5Ti99VxtY3vntaSDm2agzQTeqisbjF45spozmFXISxBgZwN66
ZnX53qdSOU43ynqc4dAi6OVsPvtPJXNk0NGl5vUX2P6zk1Kc8H9OpfRpFF0gGpbK
VjtmJfrs048aLZXHi60pswHCTAuj7/WbXSkqNw7M83nAdKy6XJWexFBMX/LyA4uW
DWUpmE0MaQzGd313hRTrfOMHBsLbJtI+5dswnax6nWiiKkCUfBRsDD0M1ikC9fdm
jiz/UWD1dZcgw7PEm3Q6qoKVEuddl/ArHw2imqGzGnhKfovSgy27jfEoNcFhgvBx
wb72pDvgXBNEOVTMK6tWciFxaL5yHbn2y94iZA/JdTMvtXwp9AOVn2weCT4hONTb
g9TO9ZkikhjuCE5dTg0Wss3CvyOc16QWC/yc5Nsve/jucwJVIAggQekZTVG3dHpd
R7ka7nVqQJTIq6D/0d/rXEfircpBsnPY/gQr6FX/ydBgWgtRWT1VzyI/U2Up4U8y
Ei2o8hiRSscskRx4t8ykm+cMRI+oCkYSOWuatTsa5FX9g5n3hDB1wrhSfbhXmRWs
uzTeIPFfYEhzqe1+plrT2DMTjZnSYbi0lgfhznJ3yRoqrb+guqmCQPbPW9XNS5Ky
CONC24vYrDAOU10axJs/JVyjydEsLXh3fCOMdwGJ2WUH0Xy07AV8hntzyR6oCACk
XjUt8gwpE4T75UN1NB0qC/AiCfAlUyYJVUijVfJpytXlnXSS3GEzIYeh34J3qNn3
/WYAV98EKLxGF/LAS5G63hOOAaDJdPj1qvs+TZdcSTqw0IdpuTZkYf0rvyJcXm7W
B2flJDgp3LQiSZRGrn9BcDdTy78OtJuQ0ip9V+IfzO6Lpcm1N8Zd9N94ZwrXnWK9
FKfpkesDZ+Zd2lcuYmhxFwqen9YOhoyVKA/cruaNeynQ+Hoz5Lpyvpw4P3Z+vmtC
dPttr0Z/QLuQGdNvuW19j2PXNg25zWUQzbRYPlq+TuIr59O+1fblX24/qfWmlJPL
j7zMddq1XwwoozJ9+gNjPffUa0re5d8MubC5cxJMn1N2qgb9UheMHhN3jezJsIM+
7WPYEKwbYyZ3KA/Pw+Y9TFRY/8zfykMEshai4Dwd6fKs9kjSCU71ufko8RjM2VSz
WsASNVNyaNoDa7WLZ+QsT9D2WmB7RhzBUn4/k5UvnJ4ccgX1bRq0wjRAjDsQ5681
hxTnKxsIKj4LS1zm29cq2yb0zglPFPlOkFIaz4bcc/BirPlpUK6VE3DrecEueFuM
Wx0hKXUnDQnbbGbW2Hmpr+MtMCciLjeUIqPi7ob1jma7s+L26XY4w/fw17e83cam
LTxvfSh+5BHYAY8InkBL7PJzyALCiX3qCiNBxdk1M9FgYJ6lhmMtywzoog153vZh
hLSx72pjVH8Sa5xR7Sp9o86awj0BZPboKmpzTrcjYHvkx0i9AOBBUMHEzF83Q3O4
60fQhvlmwRxqC75rcQUIba26w15P/vVd0nzfYJsNxJ4u/cWNRSZxF4TDV5CoBWfX
JPRa/wAFGBd8C0/I57VD0k8x0szkGDE+pZehRlBZK9HeP7d7bBZTDG3KszMyGqql
MoYiAFkP2mLlDOoib929DFKPdEQ/uJ7xxHwGKr3DpnWG59FA3mK3l6pp3wIsEUfw
KqVqs/bJ2f0wxEOWCj97BW7l9gs/GJxurXoi5W6RliFNzcDnIypNwXllfpROFLEf
iSGynww3HCOg+yTnvbfD/nlG6vwTHxPJdmZC1J7VQF7yHzkEshhMJ+CyE9fXxuNK
s/FdhM/TMFcElN1N0T2TfJU2pUSxhzf328ZFeeGL1yQdC0YdbKZY96za0Bjy1ikd
N7uiaDFHOWGxvoU3SBLIt3AiOMBcZ5yeIPRqNtiE+hnxeTy0+r4Oy3pWA47dC/zH
/BAQ3zi5Xrjpf98qOO0J6wPxtUDIpRrYwOOjunUwbfaelCKfkLsniF8Z8jaU0cYe
+H2bU7ZVwHx9a7y6sUfql1YYv+cH1EnZPldYuWUlm59O3iOMP9OJ/kWCSvs+iCzG
EQ3hYyZQer2t8AtbYRif+sR9qcKpRm1FKN1Xz+DgFxN8bpOzpCh3S2oqvsYcrSxw
GOihPZ1w/LzgrMMJZfV4khzqo5cib4FtnmyaqE1q0qjzi4k7HIqShIhsVOtKJKZ3
QIztiuVYxzom3WqJ5b3b/wbN4pkK3HGOWiiULZd+ZJT4pyEts6Ir8M37aEGQxtN/
VbuF3AZ1qr4Qg21cAxOMAPeb0TO1ku3KLeEoED/U4ExqmqmDRJ/bGczgToR15XJ6
53eMVOL6PLIzQGI1vTOs/ulAEAm7E4ymY89/JEIzO24338UYLZ1Ylj/S0jJvEOLG
/rlHSHqe9M2vYM4m5waT7ALvIUhEdK9XZ2305UTiLzDWuHepkxvWm66ZA3e74u4Q
kkP79FncPNcL/eTR3nQvXLUbVH/UnmrOzMLvKQD1sUimzlcyFuXZckh0WNbeqRDo
OlLdZZM79t35UMcS0SyDVYRFJwEJPl7TcaaPik3oOraRm7du6CBum5Q1NVtH/6I0
VdZM2Dl27SFAJ8L0/6cVkkDAektutm0hOhBnpZ+KNro4oN7lwhgGYQdUjTsCtJ3W
3r16H/YoZCJklcKIwmGWdngoXTY46LmYz4YcueXjNtYNy3nu8AYTRVNfZ/8sBi9j
FDcdjVmCFC9TN4MBiFanguehQkchexsxeANWPwH8Ai09lH4xVGIgEHwEZHFf97Tq
2z3pAiX4kEpdvQsUfBl4NQMOwbA842hxX/vYpTk90fg13tbMIj6r6FW1acC3+XkW
cVWHEfAuPA+HQxgv/T6AuL63NNEBDdKYu/VQ7ribo6VThrwfb4oyPve4tDPGnF/k
Bc2kiLCI8EjabxlDNJ4fp6h2PSJxiQeV9a7642TvftQAEkvmG1bZYCVZxcdskFxY
J0RNIcCU59g/BRJ5Vn4fgZJ3aa4LR4B6PeA1c3VdntBdQW0Tj7VG8JBd7EPg37+t
m4Fsd7iMwLerwOp2bkPp1goz6jZRWf/qkthqchMoE3kC/bQtORlUL4UjDeBfwFbH
Gudd7XrHFTqRfNqKVdA9D1k5aZJl5q3MTDtvjZ0HSzXQboB9UHaN0jvrMetfvewW
JL/TEw/7UUBfMAMy6nli/GHnSEjnWqqQ2+FuEfBixCie1D3Xc9EmI5xg6ukv53uU
icgznrzoFiIOnMQdaV9uBGGsVLNdt306fvBgdPnhNI0/YTPT2GBo1tb54jP+oyV3
JhFRwNET8LokkUbDaiHYIebVVVn9Wqr6N2+N9qIhkuERbFv8U0t0liAnyAT4QfYo
KUhMFHoMYJ2VHCtQb/rNL4Iqo1kHkyYPsrhBzk8F45vTl/AxDeozM/ySeX804MZA
BLhBsc5DQU5wQkVTHXRRSFJpwgkrkyT3RH1uNayoO3CeoSISBbaxF1FufR3cYsy5
8T5SVpgGm0DGFoLPNtsn6yL86MqKMVU7BSF+IRop3PXzSSAS/WhlNabj/ocT87/O
D6XR1DOOkDUZe9v1jdOYyyPDTnUVm9jIw1yNQjB9mS+SQHL/s6QjLoRVTuP9eSpZ
6YeLP5EbADwjubwd4vQ3DiU1Hu6bmruRwOUbZI319mwqeSvn0FIKjuLP28hE091M
BUaKDt0XRK4NsgLMHYYSkAteL2l1EylbEFFjZZDeBYdS2B03byD6VcVXF/+h2tPF
D700H3Chkr2qyjOItnp6wwC5Mv3NoWAoMikd0g3CMuhTRgAyYoOcFH5PYu5akJBg
/gEsuxYz37Vn8Q673jpjPOlr8kYrq6nqAOhqqwtYdsooJ6/YI3BltSblQJj5Nj5h
rxdoeiCVObAqHuCsSXI5GzC/lEtKfa8i/jjCBbTUxi9DPN9aiSDPu68eksBE/oVe
JgSaF4xQyEfTSERqWoUnRhjcY/xYdkrGpbNxdGrL9AzWy99ZH+iCVjjQTZrPmQ+8
eBUeqGSo6CRH5CNvgFxyicU1lbX0iiHgOLWqLfx5xn0Uot1hx9GKAZFVWVqEbaOJ
B+qX5fI6tgnpB6f8XxAi3e3n3y0AZTEJUQb5nC6jWlGOjtgEza+CqOoXi3BAnPUj
Hs8koAF0hp7EXkWL8XPo7VMM0wluhE7wGTSfp0pEZyynkOjaLWCWwj24DIvamz9D
EYuaBU1SomaxEQJcEU/HRBR0epWHfJNkeqa6kWPVnhKDazQk8Zwtp+Taxxg5uGwW
sh3fnW0c08ixBgyC6TShsOLjpLHbWLlfmWKr2eBj4klHSP3bQh5CqS+ja9ZhdmQN
scSb9KEkDBJspbtQyqwm8qpf+4mqYDH0kkLENgpZyIpBzGaxWFD18Qg4LfrIK7sk
qBr2+a9C5xZ+sMyoRSiENz1+/W98wXNvxH40K9IqyJZrcEfpixoIRStitRSJgHHd
kPo2G6M5Vfp1yj7yivzOo5ZuTNqnmk/ZQFzrXC0cMfU+eJ6UVbA3Idxt8xMx6P+N
FoquT2BNzbmmob4++6PVxGL5RIWGZXCl6uu9ouhdqStgc+BEu/h1Bt0p/vMnBM/r
ZwSGoZqYiM7omdiV0zx7aw+4DqdLKrr4tv0XnGybNibyjwYViHJq6CqqlLh5kE8j
R6lGm1bsl+If+1qxW4pL29Z8SHeienwBoUSSWcphbxNhNS7I1xO6T+/0WQ4ix7DK
jS7gt9GSH+woFYgeHpIM65EjR8A/uLev1wk2NsymdKySgFkZmXObdrFiN0AOOUGy
KDHvV+thaaynzbowRmEbTZ8Lg4nD9cuaJMxSe3SnuUQbuIOgO5txIqbp0xDlMdrL
JDaV4vBCEbAxpeqfewgL5kS8PxsdNKEDkJGB9T86zdc+Onbb35yaDKM3rDFqB/Ei
HLiaOB6mD5M5uXqC3GWjikNmFp6f6F+JJ4AgJNzPI+JvJbAR4YqlH79I7flMEq1m
2aEyQreXiWFna39eQKJuwwss1VREhdtGo2/DVb/ONX5GU2XaLOlrDU/PahOCUCMs
eyaR+hcz5grQpkR9I0eW5bV8VcOIp1dPTAsWf429D+Pk/fEbQ7mKEUrHxgjDEYfk
nIwy6ir20MfHmoEhfDW04NSWmRChtv2avKXdxX5jB/i830+KKcmXbQTQwVZStNd1
y4qZtlmgZq4khRsEUlta2S8Uiv0EGu5OmAwL9SpKlxQCgCt+ukVGGIJxISgxHRlV
cjktbAT3sxvoSRKzO3xNBJSCzsfCMSG2IA3Y1N4W2G1xVujU+QPmjdEop4/0+1nT
Ggl4ld2cy83+svtlx1zEfdbS9X+F9NFSeIG+w3+1QfYJ2mFn8m1b2wnZOmJw3fuU
S30a9yQdfvstIYwKHqdOIpkrguhkPc0o/7Z7NxUt/kWMskM3fTOt+Say9+SegQE5
NKS+/EYrPqYitOj/LYhabpPflsTbIuFfjDl8AwaZP8VbzUYvw0BzWY5l0U7qNCL9
KCBkPbnCLhJinf4aqWRe3dI1B7EfOcl7XqGkQayiSCuOSXqkG25F2ORkIVMWfCHh
PdJ7EmISj8Pfo4CVXoJbCTVboP16DpTyotmyh5D+z8jbPQOnlT2obQJpdIIpyjIM
hZSdAHp+RtnaA4jtWDaou+LAmDR4hQggvehXOzIQVlJ+hztsWhzzJmtVtwsiBhah
+ZuNbV+pO7fWvcc4kcsrapUGm+yxeaTXSMKnFAI81QIbo8ZtQxSHh8c8tQE22rL/
EP5s6BzDq+HXUShUnYIYx5PlwnvYfmawEvACy0CV4JzQ6Z6GxTnvFny86YyuEH6Y
JiUgfjtWj51vlGIMBrauKtOwmUgt453EvvgdDGOGof+LqPJNoBrgHEj6O/nsmHuE
CuaiZl2hnCdJJfvxmr7rPiDfL1/SxuHQZdfD4SK8KHjgMuxxdwQMlEVxRm3Ke0A1
lmSktuHJAhtC62ZM8jgvi/Gf14jJclC/SnjqeXVNPtyb1beCBiZXhh+r/cwqvN6h
R+NvROEdsAJ2Bz/w/tnhh4erKe9u6mBxdKiNk1PmdbOP9H1c1LchhtWCc0m7GoVR
a/NjuSo+EIH6pFqASLaLhBxx+GOxX7PEz2raLLXv//Qawt8YQngvjNmqGkqTc5mQ
aBOaWNyQFBCcmYZczdLk8JDSaUK1cKVUan0V8f8cSKFlgsKV9G1fYj8Afz1Hnot+
ePWlFKmytxrCL3l86x967+Ddv+AuGRI3Y+D5Qtn+wPmQ8XMJyHp1yNQ7uD4STkGu
Ig8/QCXEMn5Co7z0BgunLDnnMrE6ZXnpG8PkK2g4IR4+Rs9LSwwJeVatbVTiZpzc
Kty82W9S9GQplPxtac4SjQkiJXmaX6dG3b1uZO4xOFOmV1v0UIvF0P0SzxFw6Pxv
vlq85vM/ADu8FrRz9ZOMoTrt3T3LxRQlx9L4dzwJr9+4WYZAymI/NXfPUpG9gS/k
VerFaQP+xhhQnrene+NMRuplvBFVL2ojFMEWrdEUZPdWldcixNFWhdEd1D1O/NT+
wzZ33kgW3J7ZKSpxsyoHiVG/j04io9POu3Bb3/oMGHa8hewj0qhQlNvSLHdLst0L
HDPKA8QxlyxM2U35nY2qrut5M8zFOasxP5Zg4bXN9sWg3ZyrY4Sp+NQPjXohbn5g
SYzT9Hd9MdG4add+pZbyZ8iriscw9CKmDEcKsaj4Lqs9X9quJzXgUbMBtBrzeHEt
iz3o4lvZDLT6kqoCruVfTdg6DO4/3Rp8ohd2MCe6i8BVdWXQnSqhaLfqd/dPy9NO
X2n1lB7eMs6GN5qq/MHrBxmBGf0I0Oc8zRIZZLRZ+OixDetybAWPZ6VfE1Wq8UmV
dx+mK18rbXkB0TVBrW+NVHThZxK9pEjzOT/ObqzsfuXdzg6o1FtBa/LYguF5TNoK
52xZMWU+cqfsRBDhD/+w/qPaMDaAlVi1XtgfGyh6hsch66Kq9E2puEtQQxhyp9gY
V6QmVMv5i4q3a+OVafWcO+d7eszsDD4v8+J5Ubptwh5GQKSsdViDmvNKNgxnjlOv
1WHyqR8py3shcgrBQT1lhwpKbGgUTLLJzJsR+3Bgx5WQAYIJohDX0zZV1IL34q0p
kRsf/ELgVF+G4LkWvXjqvkopvwXQSl72LZdcDlgb8r5wB/5crGi68BL5ABg1jRyr
EYh464d+FTPdOdxXpGkYGjwLkEg0IJPM5QhSg+HBiabXabNmYbg+tQu4wmSSrTng
Ht436z0kFxB5+0ga/AxSF8Xk3gl50n0o5kjyrigq2RV1JQbo/ln6DM5vxSPNr/4g
A+zdznwNiKSmovC/wMbnv84L/4lKtuC1mBN7c0kL2CjCqfZclA/4/vIJYxi1pV3Y
PnvouMZBqEWuJ51E4qFL52gKvunNof7l5AGSIAD9rQ8R63MUf9QUfcp+L6etvcQo
MKWP+3Y/6LQKvqEeR4w4Bimry2rqSi0DvYNtnmPIDBymk03Ld+pjRdGHGBvY80iQ
iLtSTqwnMxINeLr9fG8RgBZwRIYUDKha8FPpUAGnddOWv1MxyuYdzb0fHQimPoky
AbQYCtVidd/wWGpcZg/YFUmMO7HhFyNZ/ukCWG2svGreONliV5d+cmXUD0MeEkoE
zjkIazgb/TxTwAUYoDKWLkECwjhA2C18j5Cl0Ddx1j7orIQNPUKGmraUWbd55yi9
Mb/XGnJi0f2hXk87PPwSMxFz5HwrcEqiOIWmmez/5JezNW2RPApwtiQx3a4AS4ry
I14QVaHP8GTaUocr1/AyHS0US92sEB1ZeubWxCaSiMLpajGSUM2yEg1/J+mhHF1J
CPotEoWRdPtqN8PCPM0LeN5QHmSQ330+97wOeUR22O8AXqi/EN4VqLkC+ekVRW0M
1njMnQCLcyNQVZvvNhiJma41IHD+y5/QU3OiiBBS75trow96LnDnqNTTNJx4b6m3
BckMJ2PyqjlHy8fvmD6fN7BsNER2MUpCghWaQqpsiHl2sZj1SyliSeot8ivWuaRn
Aovpwtznt5B6FsZmHzq0OgNpr5TqoEYbTvMBNlEY0bSayPFrd3NkNxqXEIEJ9JQD
gdYxNbBaY2J/UcY5I9DfJYJLQLP6Tvhc0fjREUYrJzU7AqsEUNjzXlQ5pqCFm6K5
aQ6Oex504ibGz6YsWLR/uJ79j+bdq08TBu5msgDPv5d2oXwq395+vCbnwlSsL++V
BOA8xEXNgKkkDYBU99ueK0nDJVjVj4DYdGXAPS/P/KTgdTQiB83eGtaRP3b2lnBI
O7QmiuLornnqNZj25OEBmfAZqUMCfiiNFvP3mptW7UzbuQhoVtTV3vveAAQh27FS
diL5PoeZ3wUHz3cRWU6wdVW62a/hUTlfXc72asmoEcRDLXt161fBULjJ4c0AvTPl
iJYwtEA4IFcH3fvd08el1gHGHNC5ohZQm9QWmRt+SuaOErYtAkUhXB8mFqv/2Cev
JTWf0aQ4v2DQHtf569DFbb7/vkA7Jdx0w+yx9yhayapzsy3N/mZTFJid2O4Hclvm
cljVoelToEkHpeAcnl5Dq7KjG5vsSr6qLd69zQUayR0AiyX14Lx0ViVr2W9IisVy
yPAxLeWk0pDqkbzd+lcrG25g5dFn2gbANSkaUYVx1D1GQV6QjHobs+akdMHXGbjY
CoXUrVuGMmhZakwKIZum4A8YypdH8P9TxcnQuhQiFs6E7PWKF5TEeWnuz3F9q0B4
ILNWJVTgvjlCpEpNjd/WET06sK0oKjgzLMARjbX03CpYKatx5AcXhEsmN6SHf9Kz
KJXzb7ceqg2OYGJFP/em0WDChzqgY2QjjWxvqISLeDCU6J5gJLzn6ggl14XOIovZ
zmodbGjF3PL0mdxmnZWwlLf6yU4qmTPjSznFKkoipCPvp6VZQ7y0N9h/lOc6RdR3
A2XXMVKmxHdtNObQQ1ORFcviNXemCV20ICbILRGy5mAdaFsGb9H554DRy8qa43zP
Zt1qPAaqpUCpIm2Pvdf3ibp1AOm/WtP2bRR4TuEO1iLSPekFdMrSvsQPOU8Md4Oz
dcc29JelgGLJtd5/jXzv3K6y2T4kBAEb3ZD4Z8AlrXgJz02Ub4LtzKAEzv+yasZd
P9PPiLLP6xhrWoyeqbx5rMRjeHERRSzJwLS+jgP3aTT2Jqk9ORxAuhG5qCccj5CI
eZvbRTeE090M0N1ZSC8Uc662ZkjHRIqsb9Oc6ey/qyjL0Kuh4One2dYyh2gLFzNM
ZCUD7SL3jObU5Lzz1CJlQVt6siz8Ip9mvUu+k3NkbP7zgO/c0NsRa92934jbxE7D
uoMKmUnLqVw2UYAgDHqRBN4ZlImFh9J+q//iLVLUcZWBLO90pezsR+k2fwyQ1NUh
8IPITysTFFXeVGr9NPbVInrNMF6cSFaUTnCeIQdkbw4eiwWjd52qX0HKCwKxPvk5
KDTwCKlFP1zAqsAF8n0kjeBPqkqfZJwqHFol2kmwwsq+FJSq9cbpxnArlWvSd6dv
Du0AQ8O3MII9QOuxXJo5mPBgGdO9Gb1UVHdRyz/hFtw5zm76UjWy4lnduT5mh+Wv
wW2WqnBApS+4efZBvmQfzEqvSTQqjW8RBvCnc/2HLSBxcwP719zFEZefAa5iRq3K
FFXd24e0ejL/8IKa4quE142t4LMor/4su+/2aRjrLt5LphNL3L0oljXjURj+BGPj
BXr2s2cTDo+GltOtAyShZQb7nZ1iHQSxC48L+BhIVVeHBVy1s9n3+plRO/4NJffD
w+kXEsmrto5RdSS8bPLBWfbnngLAQhPBkGATJ4RER2K5HEoijz2yx2s0Ar+WhR9S
X2l0cnb2neZVp3m143cKJSuKnBEq/j4L89O0KxbByfu9BW38dssbRCE65a4YMyGu
gEUA9ltFrBqKtbp2sBGyCBTCDxU83DxRTN1HWWKwwSKz9tYXRQbu6/PWopn/YJ+u
VU5ikCfbqTEI8Son0gj08ZsrNZO3nG6ZBEZm7zenBfziQDaf2jdgb2JuAlT3KqPP
YL6Mylb0+zx8fd3kXVdFImad01AxitkrRiEm7fk9J+mp2tSvN+uB8DTlqUt7Hf2L
CkiR9GEGjtgZFviS+YDN9f1VzQc73BP/qzcEX1cx4EgyRSgJ4xz+Bf9XypbGC2xH
IYE0BEFE/cuZjxyiVNIHjqp96oKILwzmQmwpES46tdLRwQtWVh5j0RrgWPMxjxdr
8M7ny8VMfpD8TSUF+ALiPxwVYKok+YJIabcmwNSFlw024DU8RoPQWfs8OBJ0DKxH
H5GZLHF/XLiGRPxwmVvsvYxKbnriiiX/8MUQFi13RnUpLJlJuDu8b+rIyEvAXCYj
kZ9yrKTfzxMia2nTTas18YE3AChBG9dUWAOTA4pbuTypliXpFndmVM9ArUpzSSUO
AKZ8n52Pfat24Y1X0kNCJtw1FUgcJ4i/euHPXoOlFuagvuPLI5Rpe3tz1urs+lao
uHMF0h5k90zeg2Vc5MJAlb3/L26B96vK2/5KsgQnD13ggC1l0DWrkn3MnVsaPQxA
knj0J51++9PbqqAm+Oa/YhKzRMbKNyz6ssFtjo09D1LMWu0AY2Ozpl2qtLaCHtzL
lL0mnfPRK7C4nj8vtd0rID4KcAQvlRelfecDlvs+Ij6TtAvV3qDb7V+sQhCKtIjZ
uVxoP+Tdn+5ZFlbvoU3WuTD6IPUX5oNgW079C7UURh5M0OaLIT5m7bqPz2jaxTWK
6xvGD8MfE2usN5KlvSN3/RWqQqbhHeLRIQyOlJe17mIBOYaOQ4Y+MXQwnYLaPj3X
SSZI7uA4K+/gGTKaxP8Ukx/8d+T9DD4ySIRiXig7oXWRew9vFNznLenS+GKvZNW3
HsFaopvTG+ypCyc/uCkWLvmxceqKXy7J2UdhWjt0hNV03DXFuSUa3TJ389Vp7E+b
oNHnsAhhF4x2xTM8KugVWAGK2BAeDK/EfFnu19UHEOC9fEB0TucQTV3qEEfvYNVC
7NhNR2ZqcgV1NX8VriGCyqWF7eB/GGCcPDY2G3cwXaJwFyjEfoENZdyZzJyhJTiu
mT1wN6UL+NBhalX/BOTgBVko27dBLiuywt0ASpcAWCnXFDHogZ9jq39KXGwwquhJ
euwz4oDnhUI8bAS9xBpQGsMwFUhH8sfTnK1eDYXCBzbzpA1PZWqc/EVmg4D5W3ci
EiSUt2vc8X81OWTk+QDn33GI0kOIlsjfaP+SfAFFnEHrn3ISvc2ZZCXZ85y0KlK0
0jsSLeU2jvMJEMQFiatiGglUDEl9b6yiFeIp94LosQIHKe11i3TN5qiv0ZOVhCfq
KwQAnaB5vgvZkGavd2dAGxLgEeJl08JinwqaF3CoDMMIGRT3+8r580ZpJTt1XwP+
4eQ+Mkb7HB4bpQyhzBJ9bLq8nQlEWgtJSih/CQNZg/UhKYYubsl3pSPc3xUdSo55
UtNhNkRUVOpO7n9BbHoHuBzqOUU72Ml6Licpqg7q17HgbqsW2CrFxwK4w5ObLKz+
p5WV1ceQcxokccHFO6Uq6C/j9z76GPoNF6zM5RA0+IVtbeFs6buYn8ovM5Vr5V0y
Lvnbb39GHvnUEae8s6WmoyBzjCxt+6LTSe4qAEYFp4D5mH+gMzmv4KL2kdFNUKcu
E01Gg/w2rV5i2hZsvf4EKDclYyfrCL5iSTcDwt+EF467b86IyT7rrUJowxffkNUz
YZP6tQ0tAp3BnGXmTHf6DQ8QxGfkWLws1dvBh2vnyFY2KO/o6JrrAf4TOwWVHhvc
R2V8Idd1LDoFOo0ffCVRKKauX3ihNEtJjd6M9RJ+N5jwFPsz13emZlhhR3YC1lmz
3WBxo0BZoITem7CcKGmvzbfKFmgITJHJVUxakNtv8a0jzTB1yga43jC31VutFrPP
AnMmKZ8/fOdYRfiJchztSDXm+WcB4JFNh805ojWRmCW7IYCs3Q10NlxiG+M+bH4j
wW3fzrYgSgM0vheS7Ao5tCWdYyYpjLWikh6EjYIRuN4zWpSgGBrT7RTtrV2wstlX
GOYctG74sz3iUKp8xill2v1AgF+KMD59TiszSWbzoEh+SyodM7IcUxJythwEjgiR
PVFp3B/YtQiH79bAYB2wYFvOPHqhK7yudXl+bMRsGBpGgtRlpGgAxkrbX3ONXkyw
ggq7lfiVlzML302/fLnXDBMQo2SbWiMTb8Gns8RRf/G7h4fAknBgKohSPB7FU8Iy
DMEhpS1LV6BjkrvP9h1cJI66Sg0UY5YEjYj9YtvpgcB9jSyx7XPM/HDKDvfFFglj
ALTG3CdsKz/G/flvTUPlyL7790jaP0/8dPcwIVVTnwgB8hfqIFoAJ8sBGO7P3QRV
1AXDgw7kM/tUpV4EMuhrw3Ytyskd8i+M2cS46nqO67mKuxm46eFZ7qsR7uWXhj76
2HWG9+rd8Vazn15Q5CeYqLgT9Iz5eNAGUFradlD7fUHv1mfbWAaxZrCF2aDPrF/B
8ueEihuVJSBicBMkPZT2jPRBZz9qTB7sqXkLPb6YKWNO9wfJO7JY/zfDYF5pY2/d
nc+Ku6D7tr8qSCcZzbE8IY6pVS9lX6rO/EVTXy1TPzQpB8X9JEKcqsGce7txX3G+
pFP4kBghkYXx6uM7cawV0Qfh5Y6Vov+/7bFL5kM2mGlS3l16wzmO3ToDds8BbRwA
4Y6bRc3wwvpKbDLKs+x3vuCiTB/XX9Krak2y1+cirjpWW60zx+a1iYFGmrBfhq68
s6Haxx9ZN4sA9VFJpd/vErkoAb1HJWyT5aGofesIINwg/aFfCNJE+upmEawfYf6V
ulu7GW3mwgXsioTi3SuiqVsn7qx9+3VRymP/qFm6Pe2mjhYzod3GwRvkold8nIC6
fEI1YTB51oMybNJncoytenSFHpdkWpPlSb/x2vrkWehZ9oYQQfyixhB0pvLTNS4e
I6xlqhYRI7Njhmj4ehjbbNjm/dh24FineOLdLgNaAakC71AcaW44PGEka6iRUdqQ
lZvXb84olw6y61gMill1A30I9PTyHG083ZGAiulcfZkkKp3gQ5qXkMFvwGErQpgJ
hqo7YFa1vEiicuXA3RdtRMyaOgcBXwXJQezqFvsG14pdQ+XAsikrzppRxCIeTKI1
87suPiCuc+S9qGif6cHUP2FIANk7KJWjSvv5x6s+t3bbbK+51RvqEraqPkKGYa+G
kc/65dXEUyie9/kUn0qSdsU52NHVW19tQzNIQon/347QTW18e+8JpdZxZoMxusoV
dHwZE1p2VeF81AakJTamMW8DIHKTGMuelKx4Df3IMznZ45EWI0WTjVEvJo9f1ELU
bZBsdYya5l/+0OD53vosdXVZUDqBvj2bAXJWQRVCEhdjZb3CD1Cf4dTtqfhNhsu5
zRVqanae+UXVlNSZy39zxA86HEMnpNECM+g6qaDMRmNhnM0VarV4V10jhYZZ7AQX
4Q1cNdyCTwlyX5DNtyEGR2TsqKJLuaLI54hIIfPal/tsL0WIXJyuV7z6PbQrMv12
2DG3gA+5MWscNjN/cESxzyeI3rTkFgGw+rBlOgNC2A/1RDu8pip0sSZVb6bF+/r9
QItJ2ZiN7ciMkZq2xJ9ODNZNm6AC0XFkP1dZ5XcyIbbGvavTUTrHcfZfYxJ2DwTV
/indpKKj0vKu4PPu0N5Q6IJkLduTH1NBSlfVYdR/atCyqwiHf0JWc/JyVwbK5qh7
6HDGSAAyj4IE44Xh63wIN2oxRKfSCCvVDhDRwRqCj9YrKu+W0Pmb1+n+lmI7gJ8d
q8gK0+ChswzBolUrQjaq37OFuz5iVDIru6rtjXDaZMMpBpWDIuBO02qOEoFojo9M
kE9+nOcfIyLrSIwbLb+N2e0dDRkM23rDdTIvrxvghx15Tdf2s5nI7/gstIUCkgRC
lRoWt6U9XqoXI66mdMtzg5IbS+80Zo7N7V9knxLV/iqvQ6EjPCxaIhSmaEKnXkTD
1BTkxlIWKLUqd1V6YI4HUSO64ShPxcqPpGfXO6sqN6RRWRlMZ5/SNGsSm+5RqDLi
MFdIVvV4CJdC916DSYcwFdbB80bjaPKtJS/+tjICJYVGpB+hezn9PjeFqTZ8Uxk3
3JYJ5skZjJtFWUqaCbhXBC2Qs6lq/8SX4VStythpp4zR0UFlgYsYRld0gO01dyDM
jUPJ9xG/6Em9VOe3J4HgwpkSJ7zZFMXbJprUtQ9swQmfQgVtaW7de8BWQY5dAw42
xW7ZnziMMif6dnpoKtNeEB1BrC5voUC90A/1t/0bWrHjA250xzGPdqrjFBoOIvip
8CbM5PMKDTkjeDDEIIdN/EZcTYVoVAbU0BosiskN+4F1bgyM9/GnN0XWieki34ar
ybBAfQPNwnAQNqcEqGPhl2T1HgEAuteRI6p0tQhcAzPpOtsY6Z6rbcMlC+0PUzex
hgjf1Z1Mb58C7zlxxBkowFoUqcHfv0v7RtXXhvygwl9xWheHbT73CsJ/db4bPobo
2AaXdnoA7gEjJAKMPTEjQuP6s+8dIbyvcdlznqgLLObPcrhSW5yumnZUVWJMPXB1
RqoxqBD6WAZKFtI45WGsV+I0QKNbgkbhRA9e1zxMIJ0JGXQF5pwtJ3obqMrkRqbG
4xkqP34cqMVz9hntSiJ7tTV0kc4Lxz1CRo1gQ3WeGa+j0DXoDQ1QHdE61nq8sYCM
qYS3wBuxUGzgffExT+Ws5SwgWrtpuqB4YynaNpt8dsRD87ntu2e2LMUsAvqK0CEP
YSiwnTvVCinYsZuBStMBfkY/SPAwPpmQVCVxBxcNP3pqDHVaPXSQcEy7YRrAFwKG
ok+ypCiFTPZQPN5NkeWWL8ywKYM5L/w9ocwRecLzb9exZng+3l9Uwci7eb66S9jR
PxhjvDqMEua1YizRduMRe4RLu/G6lVDO7YRYTnCdVBvM3pu65JA4OAYBdGrX2/M9
ac7aiKQwMkwtotSaVgIynzpjnOVIzO+mWf1Kbhv2BIz1ZlAwnaXwVfIfe/sdPu3Q
CPOy/XD9Dk9jD7KBefBbA53XjL5isoCOKJAs8gmuKJ4HoAc83de5WVvZTyTH0I/s
0SxHydD1yOm8KeWFWRDnqSJCfWA5/t0TRfzFhH0T+AVnOTcIVxcjEXmBuRYepSYi
PBKd+e0ZKYTX0AtjE8ULmxgPLKgXqLkvYp9WKky+zgxzjzdVpYXyv7wypgHLkapN
1noNOiPOSDGhszeBxBc0qlK6R6bl8ekwEg0uUAfyY4i04m2V4jSiSpeHLgkZxiCk
0ryidpW9GqjSTUXC85AQpe4cJktd85iNTfVz3kDj1hsHlUbWg2WzVjNGP4rJTbs4
rGEzgk3b1uYvrSdAucm4Bz6vDfcdULzu4yJQ0/AAxDGpzdsTxQatPANWvCdznY7H
lwVzobxLtPa0h8whFrsAIbPow17UgcaMpbkOBPd0xgLMXISVF+UvOxlP3UJfinzv
TDpGIBpzDHjuvOUWIsatSj4A2Gbpk0o+EC0it9PM324jhsl6F3TdoOAaRLui0BIZ
g8HuWvjt4ZojTewTj2J/V9/lC/ASHx4DK6YxpDBlnpV+pxEEemNK4RAru66ssY4a
ENOYxPQ4vD3DNioOcpMfP/BrvkgwCAmf9TNDhA+Ch8Nve0ozYmo6pKm0hvUwTyY6
u85o32y/k/WNZH4yTzwAkWahyGXzAjK9hs7hYWoUkBTSQAVkINxsTocFMsJb/epX
+U/x4zK/+Cpz9/s8P+BszhUE82soogCnPiX5wUCbpaHhnaD+wPpf+7cTYeEhrcEa
Ig9VdGHkAVqAD9Bl32yMNO6dhNAeea791wN/5G+RjW5s/Lm9e+i9EmrHcUxqk4h+
66561X+lbGIkEDrJhDhN82BYd88KyjeZovP2J9ml0B3lFpREfGivb4NRtuPHZEMl
zhAudmzQJJ3EedehUz9PGBmOX7PE/NbR2AZzpXjFS7fENXjgK0YFjyqST1+o+LIu
M+fX686iWwr2IUx7agLoQaEhcwzMSVXBkt0dfnxcg7ih2BZdKrspqyvoNIUJHfNQ
h2axqe5rkyQ2fU6U/wvcWpw/dJzo0EeN1adBaP9aILruw2V5ePsUk5cCkUFquMi1
jjcTsl8u3JsQmXvKsnbZDrJoxGQHm6AcZCTAqM/Sq9SwC7IU3E3RXMs0bpDG5lIj
Ov+iE3A5Oocfhbb2nzOI0+FQT/4bRMSu4wlKb8CtP25LV9BBxq/KjClMYEkMZbjs
3Y1f9+4ce152QyF+fmFQqcGpt9b5F+zMd9FryTYZhGEOx/5KvxjxmbksAky/4hjG
Ilrd8AqJ+9VhiYFFsnuYVKYTQlJm+evjjGm4YGo4DLisrHlUiPgU2NAhnuPTPTUw
tibFm8lyuqpM/v2w+3HhLVep3cHjS8L6jLPWp3mOCKA9bf1lMUBeu7wIbVtOl0oQ
2t/YcWaBFD5fX9m2x5U1QqwbKZNiI6BMbXrZ8unuUwUH7IsKn3toClX5zaLzi4io
M/Jm22APTHlwuWrqrYe62aACHYk1BTSGx1M5TSJto1W9OK6i49I0oPJNG+2aFaSg
yzGKWX7KTxIBvKpXrJCc2OIQz5zwFVKb5zLx3h3ikByKSg+7P2hdJySaiySPIWVz
/M+x0g8qmTce1Kmgae21H4ZFbbyTzW0+DMQWi1j4lRq+I6MpI/ar7KE6g2LTY7H6
SLnpihxMuYRzESZfkeD/Gu2ZseC9tzK5R6VwKX6SnhBpQAFcAgAKr79DsBvmoqbM
OJA/0YW/3pioCv7GH7DswA7tyM4MVO44Y4v38ESK86ISY7+UH3Cva4h8Vjfjymiq
n7ULJuvx4YM1qGyNER0O5jxh0FKrg+9awZAz17nvKJfST7z1l5DSJQfCRZpZ5Co2
IE9IIwJnHLJVmQ77LI7Kegr4Dc3RKNuI+TXVIoq9lXZ40JuVpDZumfJzi9XpsbCs
pzzsN4H1RNtBDHM81LyrATDavFkAz8afESwTliLfrcGEuSVaSKSU2WGTfQ70VQTQ
tu2sR0YAtmoZYPhSAviye3bMIH1YeLA8jmKhqwBn/cOGxRNYV4SX7giIaOvYT+BR
LvZPgsUBvytG8mTvkP48nY/0QKpgLlwIdW9Pqybx84qfq4ehJ4P8fTEBFgl6ztQi
P4S0g3YxwxkP70NLQkTE/goBdC7uGu9MpO3pi0TuYkxOZ6JLbeweygshv0LWr5GD
22Q+f0lSdY3C8k1aOuhbX/50yow9wh15yLDXdNZhtoBo6J0/UX3nAdgsbLcEq18L
sUw0XvwkyggkZ0M8tM8Gbppk9cRQQRhruZME+4j3VhmpJicv+l+0Dtc5lTtMWQI1
AqITzJsjH/JjCDTnMOQCP+uS/nSwK8FjADfMEw/6iakpaEIfRKhDrARhNFJHBByf
wcmmsunARI9kTyoXAwVYgiINTcavD7Zo++ZfyzAaqMEkchJxXYZSOxeDja8gefA1
t/qbHonSjsmQgZBR/NK10BADsfb/nCuLMn7U/9hsBEsYhzm2hbRHI2fHxBwvp/Zt
YrEELQoVMmD427zGDOYhHSy9KnAaT/Cit/7oTpaxfJN/LbDXZ5KGjQm+gsioC1Mh
Kn9RGH7UiH+6vBVlx5mvqU1OcT/ID8QQ1MxRo9TyErvQjzQwKbVCfEjzUsdQMach
Sy1vkh8bYmfZdse+SH+XyuBFH4iaCUFy27eYhmSqCx358eUGA8y62UokcwuLtBKF
GcyJmi1hZLKy4TNSOFgMs0JfKIlD0+gJ6V244snup5cxmFawsUIWmvFV9kTBcv6T
81hexEW6HN8DIVo0HQa1QbQaZ5O4EOIxhAEpRAAcWfGPzcnHuNhAKkM1jWrGH3Qo
heUs1McAT5SRktxlLdEiYim2T+AlahpZbtiGKIlhgUJCWvoMUtPcQV7gMOKu7rJw
aezrGM2U3C/yxgKVIF55h9c0MUnT3R1iI1ywvLkCEBAjRUl6tSdf4P/H1mhRIudV
2rWOHmERudgnlpfSAJMU2Loo4n3nsxScJz0hdkxKeJyHubcKDkTXlecltQdWThC0
zsXwUL1kiU1sHSdC3VX3msUxLTTCpR9E3pXZSkxxsYpTiPWxapYUjnCE9t7jPcfe
qUJ+tox/Cc6HW3GY+2v8BD3Va+3foXrXROzs3p+XQXCjLqMH4KaQmGTq5btJDSbT
CpCdCkaPOnvLjHZ+xa3aHa+cKnwY6jjPSDH139r5i8U21qofjy2cNuPe33Q01T7N
bHZSALXYmKYN2BNuTovnhz+FMpTj2/IVzY9B4tdPsd4E+GwzrdGnhOswkGrPwwb4
6+IIKB3g9YL8xdwyLPknngtz7Z5oAkfzV9bSPxHlKNzzmotvkHrdX6suacZM3rkA
0UU+Pf5xvFnV59NSKHCoCGtGI5nmgZwMkaYgJWjHK967gsX00O18F2MN06AWRYZZ
JYAfqo7trOs/YUiAF59ldD7T1GFuVU4HyU9WgKgbVv+jes2HE9PW1Za1OW5NAkvi
zBV5JEXd7Aios/0rPTskOJoNOO1NBn8LYMZQeoFhLYS+tVkikA16GkjkPKNxTNeH
DXBfkzipPFNhAHqOHrzIyWjDDy3ZuzaEBdmDO9HUljROUIot0PyLQDPAapQCH++e
E6f6Jw3aC7ee5ID4MdXaPQaTc203lf2bbYyiOdE8fCyhc4olBBrvcTp9ckBux+f0
R4ZOmSigfuadTmXbT7crd7psBCCuUJKOTHB3aL4PNFSyex3ruG1ywrQV77/UDWsq
YeNRLFdZ5QXTK/JbN1CHBTXAiRaL9K0IwtpBRDR5amCRBir+9YJraolXOXL+IHme
Nd/QUKv7riorTNXDjWNKtyht5VSAjIiSdffojZMvVa6zx189dwv5+f+/JcEOeHuE
iPQU4ogbfLPWRIvxV5f01hGbnI9iUHWIdWb2l2w0WoMzsqR9+RaJG4080LUvRuO8
L0ef9A6jHrE9fmLpGWcjiwJKhn9Z6aiDjPrbz7CVZ/awSP2Prh94QiCjCACo8962
ZJ3Qfr6t9jMeA77MyXCRvN0HDjeYHFiMFvT8UWPGRAmYy0t0HS+lG/ayzcJoczSR
K6hK2/vzG7R++ghsh97YU6gVegmqpoN5qEt902yUXqsXFPwz89lA9k+nPnQsZnGP
tyboVtAR3Tz9+nSLBZcVdlG4BdMhTdB1sD3/Toyv6Xm7YaEH1dgOiM7Jh0E+R004
HLaAaHdYkRU2CPCLtSZBhi2P3TTOEvGbYyepEKAlH7Q5CKBqNQpxtgx/6IO5GXVJ
aUqN6gqQ4t5wiF9AszndI8iX5+HYKDKBeBYvR/wTY/ainaRgAVBpdOMkGKsQBEDd
iH92WA+t+1F+cFjCpMlKwuchL4Y23cyIxcZ/kd3TpRMBnH8ZhuRdHeSORn0QdgPm
WIpPRS5iuFy6hSXXsBL/tr/E1JhoOhypxmv3u5jJ2AHQ2aw2J1vYjjNdtehR1onv
bfkNdlYOgcZW8STJr8AmIN4bk83XFoe6PJ+782aXtIm+SPZyEdb+6Qkyu1XnJu6A
y56W59U78jMJtqTQapSimtjtQ7W606gBXxH8ptOa3SyZDAiSOkpESVZf+YjizYv+
nPOXXQdyqTjMwO3SGoq6QfcW7pwrtzFFkX/GkEfVz99Ang6X4dyiNFHOE1V8nsIP
A/2jtDQXjOB98wQLRg+y/cEYoxLXRBsOnTO/EIZGBqwqG0B6faYCtHVpFPg4G9NN
6wiBGmbF5hOyRTeSnY/HDKXNIToWfulG/h3DJeK9kjd502A9ndZK0SQXZEUwbXzK
zk6QbFDlbQy1cWS0pFuUKiUp+BmUiWqpHluXFz6bhqoyk5/4rQvi3f39lj7nOPr5
Xxws7KTX6ox8jJmoI8Md9IltEqmEQsrzTZTuwRQAtNAzsfPIoa4Q0/nhD1cZYO7z
ZcL7LhvBE207SwP7O8Xl8ZJlSfeJfV6ajfvAA815186rmKZvvbOcOmFfIaczKbmC
9TuayCneptBpm6ffdEGptG3Nmdvmp1PY/3aTInBlFEXtPIRjVWPI3ydbUzliAspz
x9Q1E7zQBGEyowZ+B/PfRl/gsv0gjjrANpAOa7eTVz5cEIzTrhqs8OPKeM6W8+2A
6lrB5+9nitWpxcKdwPsM2YCruoFLJ8S/EQCp5eUWdNym+F/XJxNiYzDEBl/u4ulr
gU57n1wwlHYPqnNlyxo/cnQ9Dg36qZedLWIjvboUxDBtbpSsk/cCkFrsTjNxdTqc
Be/eTW87zRihOa6jEU449Z/4+CVG5IWT5vJCCWDiN9U1tAkO7WWwnW7hwld0NE/V
gtIyVaotbT5htS91hpVYdYrEvHYLgXPnUJ36ZtTz4VbbPGOyT+jPyWKNpgHjYgE9
i7vR0ewUpLt33+AAP5eQdd1fNZV6IUUvPi0IXyYCVYp4issZks4XAA2V+9bO8IAB
utimcVt2JcLPoWm4KfgNlrzKF4ciE+U1YaPQHW6D7QnITeTvPVImNSHCZt5Izx9U
NsCZLn0gqa1iwAhY0zsXUr3OzoxR+9pGLUjwJS7qcd7APC+wV64OKmiJbI5MFV8F
C3kLrRtzn1OV6niYa0qJ2gIcBY54+hOy9C5jnC5g1Bu7dvTRqyIe/6eD6/XrTRew
juKbiEnL6kSmXrmpyApmYYc8As+EKHssb612z2UGpN2MW/ANVFdG8mVpphQkcFOZ
YuW3ONH9u/agnIbjGmQVV60oVC1EP8QIB76odg7ipeyP7HCqmnLUaROeSufDfdIM
rsQvcJOPhD2oA0HdhvM7Y3ZEmV9H1scnMfBNqLxZMtZRiN9M3vKDBL1LftXxfkqj
+TxNelHu0XLIXgYbRpbJARBHSxoC6lWN5hUDbxHE4NnLtf6knEMIaofEVfQvkdmV
YFLiMP/rO2rvHEoWggZFDQOyTYK4vBTmsaF+c0XN/AF4+TAbqxnXCBZDLE0rSZSk
qed7P6YcNHWVLK+T9p0NOF/iTOJrD4s0Z4b3ujN1HEXEOaHwxiEiULDartwAvYmX
0lYt8mg7loWn6l9j60PUlk3M4d0AYC4rRKNB1z9B83ae6+z/22jlwSFKRcaSklLP
EchocujRMeiYRHMoNbMLKI2nKwz1njhNSqxPpAThJV8y4OwYfa3vJGADw+38pJVw
JledQSPOCNntVNaagOkdNlcLDhNA6eAEM2IOFLVUQwL1BpaW9wvZns99gv3i9MTY
BDESmvEmZAkaq2bYepMBF0D8qgWzIwkWbcCFFT7oE9yg32AjgiVLfGwDLJDPWO5z
o3O6TzTp0t1vI+An6I3SQT2dksnYNkcC9gPpy0Hk3mysAY5teOfCLT2FmOHUidOT
FFSsFEo7fxUNBOInjA8PSF5E26pfB3dniu+0w6Evc9+WDYJ0/rO7KrJvMC94JQX4
PDDw99Fht+ZuEaYEA0JYelcM2cW72+UlzKaDUY37G3jc/rmLqOGbiwWB8K5vbgSD
Yp1NoKuPqHCzsgycSfV2ufKZX51HL+ZA+AZc+ij6SahO63j3Lv5ZEMJduyjzza07
Ymg1A7zC0AHcBrRoE001DMOs9KZnug06DyTCNPlDcfUbJfcL1KzthmofgXruH5ZH
52Dyxi2s+XIarSvybLZm5+2nZ+Wh2fe9YNCyG3rGjXFVQbFjRLaYwwFalByq9/lj
sXCukhUigUu8ytym1k/0GXPvVFGC2O9mU8IWA9KJfv7FDUe22DTfjd+3m06+Dslb
yJH6Vzt35/mcKbnRF7GDdjaquOVGQ7LWQDbuIggyPVAbrCsYrJ7BYgJ595KTT74f
WroIYWe8GfLUIuolufgIyBIX67cHw2OLBY4btcTtl2GbOi29xXFbb6ZECe0hEHmB
RRV0xrc3keLT7TT51/rsGxDk/XM/2UAXS/Kfovl6S4FtmLg8FVzxRLrsn0kArC4v
sj6ze4S8N1IHifPfNGR16ceBAu6EfbaxcsQEzH32h8Kl9A5CdDTy4dLuhropVKsc
o7g7JLJJce4hvoBSlcV4W6EdO3niNbiH7phEfEMc9EY4mXbYrszbIq045BzoyCHB
Fj9gnfYUa8MeKKvTp4+mI/9VVyQ54C9mN8oNH6r5uXSmMjM8utatbOjdFBsInv5i
6Kcc92GJ8Ladu9725uIf9T2kQyEcdSOeOJzqJYGme7F+TjCzXVNBjwEMKX7fSPvQ
XfB7MKFgnP0/44puC2w/1LNP3r+yquHBKbFcKl1s7YN/oB7iIxsV4bQtSIOB6n8y
MykKhqtXJd31a+W4BoSyXHsFiweWCwULehhK1wMV7xNDPuqy19Dy7gKx29AH6OkT
CkPVu+a596yjQdtXmSM+DPhrzC208/Y1Ls6iAzIJLcwhLMAipQqdKocUJEc7WjlC
E3uCEHnuFa/hwaMGt5zBqk/uBgHn99H3OWdQvZGF8MkhYbJLKnTtHS1bwM19koze
nE4sJBYd/v+ntBIo8Dg26Xzg3Vkc4UFU5tswut/7EcXP94+1IAOe8Mh2YPl0fw0Z
FKG43vgVSk7zErf/hPTliI5AMUN99lepTdqpU5Ko4ocwNZAvZOKQq1u1QswHQlTy
bg76ggjYEyCb76TyYaAa8EZJlFot8ErUzTkejhGYLCzYWUB7h630W9nKiUrkR2wU
udfdmICYZzEtBaafj/VEl0ZDePZ0TaeOTDXUVnhRoHo8aM9vh5+tvEgq/C2uhk37
rXLmYnqyiKu3WjWHtnMMwLXjv2+Tsd66Ak+MXCsWhRCFJ6GMA1hG+cbIn8aORi4Q
aBTUJvx7TLAF7vtiofBNaoTkv3ge91CTwKGZnev9p0kcprN4t1xBZjxuaHeFhf+Y
Tj/InkZhT70t+1cU9fCuD0qV+HND691zmXqvBngTChSGnkgDzrZFCS1MiwdH3dMU
3YQrRrFBj6kY1slMdbjyOC+qbMdWf9U5tegUl9K+pzdPILUCeOuV6TmkHpqNB2Ig
MPyTQYv+WVqJXcCaPRHkjpaV/56737W8b8uGhu8VvsnJ3N/qzBgBP+TC9yL8RYmP
Fyk58EyykYNKspGjCmy8iV7XJs96xPaj55b9Gus7F10yHQ8/1xCJ+wAEnLB3SbfB
GPfH69587J/aomzosgpdQpsXGXP+bpEts46PD//1PWDuIZLgJsKyp4V/rhgP7gy0
ey3mmxgpHQnudXD6U00jwavphwvURRILcAaWLwG3kPQoWzMH/c2KYuLm+UYHCk3u
jjFnTBpXXT3C/+76E7Y0elyNVQel8uAoKywTShb8gMdS8oheEbqoDZUUBZBz+jjr
C7UurpYbekGyBZVM6Mwq9TQQU2TOUr4gpU0jymzhW+t1ByxOFByeEd4eCtlDG7pZ
nAd1XfdcGiEmYO2hzEW+Nt3JHvLXJ/oFT/b11n4YOprTOamiv+ajMh5ScX8crrYf
+Pa8alInI2qK9mvjSZDJNRRZ4e1bCobR7M6T66dzI1FAnbYRY8KkDCMt/60cSuaw
HRJczOMgPaK/X66Pw9O05w8+685IKx6bc3k5yTF0u+Esygbdv1nExVMk4TZBIfVm
DIE7b/0Fxj3F07jwiZhXZMaXXbBJ+xcVm4qwiAIsCzlPUmP8B5ms8vXC2fjWpI9n
Rk3cPnmh0K+HPfMdYs+XrO5hjyKKar1l6Nn9v1eKZqZk9lvb2r78PRuStPmfXyZi
VotPeFIt9AgEzQtY9C6SKorT5zEm6pd5sOClB3m3XSag4MFjKK6QER1JbWAY9oU1
YLD/uxIS8FDQY6cLxxyoeNY1dyUvoSzSz+FKY8OOH/zAliUd2h0zMRQnFv9//9Ju
WNT9dyf3AMEyk15fPffCDp7I1DzqIQkYrhy70ood3J3Wh/IqwHKRt/ENchmQBywc
K0Gm/lrNqNr61bX3/EMw94vAxPR+fWBzSvP7d5HG/yBkJg+SqnccsChZvsTna47J
QF0tz0r5Ir82EDNZ1GcAbEhVuFKncZ8y87CvhfoAOudnFah8SaJXyI3aisqhS3Kt
Gal8tZGu8RH4FLK78LavqRt/moPmeiuM/JM3SmwsWmZMTivlIVGsWHiATFd1UYAr
ftoQFFhWpVScOOiOes80dS7cI7qNWDgTMVIYWhGSxqqCI6Wpl+z7I5jPCT4cmPJe
ridb+5crg0+efduggVMNeRMveptHf829HalZq2w/EWkjee+ZrkaUn68tnQvF14To
9A5Bns6lygthStT/YyExRzW2HaCvyHu/rueuYMvDDBZUdTWJPcrrSGcL+RAT9cOu
yhpudyOkKqejpa7rZllPzouSz61RvpVxnx+wLZ1DVAFkDXDQ3ou/Wz7x1/vzdege
3ea86K9OnfVSmQUDQMC/cJ0nfNgxDrKLl7OVxOnX7v4Wju3yrGZXeUJWrrVAq5t5
SqTlWSw+TrCL2sxfK5BMkMoazSiM++T5KWOINjNEM1uEAbuzZYTlMoz2nd1hEsmg
SLblx2vIwgX8Jl8OP3OBAYE6y6AJigSHCcFX7JA0EcWf4sXFp9VxzJSKbGeIKEuh
TRCB+T/3xxfss+vBNDaTwS/qrll0DRmykgxqcc99gLvHxwIIvcC4ry/e/kU3XWNP
5ijFfrdKab1hv3P+S/3VGn2dJQ4tOxjkhF6P+SDDF3xNFDeprX24iFX3pms7veQD
x0aHSj+SiG3qIOHWEnVhDd9a5vygth6zn3zu44gOOG5HRrczJ0mHk2g0Og1GLMqs
oMtP2dmn8jWtGT9KaiOW8KOVN5wcFAE5BZEa5/tF1LlloDIjB3+1qR6yW4A6VWPI
YVDcuwYHMPI7jLsgzsG0UhEQKNx2iEd4B0KLjtG1RXNQimP5P6Eh5A8Z3MVDttY1
/kowhgWnIb7z44bU1sXyQ060RG/AsNvUNbZnGbjw0CkDhtQOvz4cVjSpLTSEHD+R
XS+hZVI6Gk3/Ykv9Ql2qWsIbewiDANvL55qOhfhv1wjm6WOcGnRNKJoSyqoNRN6u
D8h+Lpz4ZH8UY/TOD6qT/2kDdE3D0lN/0B9yjGs9YU4gW0Btn6h5jK81d51Ey1lD
1CnHLLH7f+CqIyuscn34R3OyZJuWlTKoJNT3MoBmySjsFHda60BtrRr64iMMcLTJ
2PhThKaXwbByW2czb4SWmFTy0/Hc8gPpJivRERsqU4J3HEtiqlAU9q1HpPiHrKO1
QdId0JW1CbwDBD3tOpCojLL4Xyarq9jTT0uctPqrOdYDsIFCJZC25i10wajQZRmZ
okWuJXh7ujIMRlB49BQOA20iP5gV2IPrWV0dfNvtuV97ZEq3ZuR22/phVa814U9g
vUsWbAxCm81EYvQUMxfjMD7jmFbEqCxYxRSVWuBTleb+s871rzxZS/LqmaSgA/TE
nS9UsrSdTm6f05XzJKEouR4FunUnNdsW6r+axRXJzZekAumd92hBAAOIMgKnU6Mv
ycqybJJo+O8jaU3LD0Mp34VLEYQGxBlN2FK3qWWvLjWG0bjIIQTDGWVRYqopruCG
YRwYv7LxAzcds++0Pqawndsy1Pf3c8B7+keKsNQyBMCLsJYLKMEhuANgdr5nKavI
LDctaV0W671g9SekzFFuR3GuI/bSN5wUA4cgOMUcioEZYrvVHOGbBYxO2ZUvpjUy
GQ0SrhBgkxBsEgoP18187Wg9rBOGm/d2S27EoyVATZ3rRMF9mBaMJjn1DmoVPxtY
kXMEWGlH+pw04DTbFlX0klLKi5jydrfXZFjWeh0mJHXWZRLhuWKettj+PWsZO3/R
IA6C/gyg1Yc92mIl2Og7wBbhs1xJBKO2vRIcWnFqk7pmn6xge7d1Ll5fDV48NBPz
8uc4hIeY5/uZlCal5e13JDjjcXYD88KZcFuyKJ0HnmqSzMRNQ9UNVhV4uSDsImab
YECD3eH1BoXcVm6AIDpPiOi7A6hQHRGBmEvVjJLLVXWy53gKhITRSj8A0fU9Lpul
7AxswCbsNviVOvETt5IfBL0BQFQcfUMpgWdJv5/dGulsTXrEEjydUWq+r4qCyp/q
KZPo3J6tQDNvOOaWWfH44bTaE0OuNjlJoL1GmxTBs9YKv7XqQP/z1sQ23JIuWEBT
gllGtEgJc7Whwm0hE35jIhVDDJNOZPgCrOEvDCJYdkli5tKiJ/kP1gAG6dadgVUI
cZGzJ8Buzkez2JHHqqlMmv29aaITUHw3Og4KhM8YWsJ4vcneoqYvoWHTO2dSttrV
jczBnCLrxJBbLqPgXl2L0hGK8G6Jl5mYb79qgSdXNnN9fpWpeX/45QddVr1Sdrlu
ymY8DPdHIvOBc+09WbZe6Yg+eGn2eWudTwzq6HChW7AkYcQ7qBVs3q2ZwOJi285K
goaRFNUnnPxuZp+1uVhN5NbxbjLKQjKZOOdLKp9ejrq44HB2+Q/hHRoagNqppm9T
eauC2ISwkmGilVqNdsszigKaTjt9PXi5m1/Hgacq4zo=
`protect END_PROTECTED
