`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agnnRL64O9kWHjdW3NCMVWsp9yhC+dZ8Islk803cKwGQXN43RrLzSEAovBVWzufw
+GHvM1wVElCgykg1nzGP9Dw+ptV0KoNrnm5vEq20bHboh3z/1b8DcVeVeQBnwnqM
rKh6XYnTG7G4igF5VzOYT9Je1IghANfOJsCtUDzhAEcTkWjbXSOrhR+mogw7kGAJ
GNk2Z+2o5OjdwIOaTsLbRR07F6hFWGLerERNh/VDzQe1mP0DiCONOseRSXT1dBUe
qLEqh+8y9FZrYfzc0o3jfRwzCWd0xkutEiQA5OLlAwVEczORE/QKLm/gOiHpBcv8
Tas16NLTmht3ApST7YiWO5lNBkzXT5vf7XFmoRqyUk+9c+HEGhUVUZGDhGOr98dx
8P96YWZLC2NId+8hmsS6LbbdVqdhknSB9L/NntEjY3lMo3x1RB+JRM+4uU+DjWgB
ByAIZEewczpzCnL2ckm297P/XcfQUl8Ky1iR0g+ryvEHIRbodO420GWossgXspMx
wbzSFv/2mAP/Sq0ME5yYKmiq0OS1BO6sH1fs4Y0Pqma9zU8F6GTiAaYCq8idDNuF
FgHZ9JLhOrTfSZYKPlVOnNszYmnazLi40IrkFNQCcw2bWMIBUzWfDtdJ54Cuj6wA
abw8/SB3uYTq/UawDS10xxgOeepNHswd683PJFdXNnq6ak75uykRXovumsmYwMzK
jm5r+F5XPyhB8QX0WVM0CFEqU2dXvW0icnvt/NPCyylNkW3B/2M1Q5eJO5uqSc9V
mT6grXZnZk+WxwMSmyBPrPc8UyntrqIrd6XV/gLQRa61Ey7igc5GG2ZVcugs9d7U
VURKEdcyTs0nYn1KkjsuYM/FdKA2DcAYFdNcHYnypkQ1Bis0aR+I/rWO8s/q57zr
peT5I642P2Ss2YSSrE3PkM8bzZ41biusHL54G8/NljMRJ4GZypZgqsZwCJp0GFsP
E6TXeqnfbB05KsDKHJ6mh8DYlpTDsjl58tgTFs4p3i3ujDIoHTlleeUWV28sLTjj
zkwOrD2/3hvdSZ3ZbW3Tyzg9g7a540Gl9DkSHv8TmBc8PXCJZYGDwb7Fvg9W96ye
o1XJcV+IL10uPRDYzyVpVt1TFzuOx7O4Xe1tfZtaQCL0i7z1lFTVr6fCXEv5AjHf
F/qCDAXrY1v10hi1hgGhCcuP0fZe7MW2ykcH7ZEk5HMkOVjCs/ybqCiSTh9WT5rE
5uO4twl5PmiAI/Ewd/15lNIrk39v/Ygz6pn9rsgomZiH6rIMYOjc2Rnj37V9k9zS
8ASX0GEHEvA/7Uwcv38zhLtklLjeZJ4QEztydhZeX5wuAFlHARUoksCKLieJ+fzs
yfFlFHT19pMB7OkNub+TjDRgF75+5413eq2Oe4QTi/1QZtMNr7E8bxZUvZ1U3XzT
+XPQTDlcyo6aiGwPk/bVpUYvlAicvL8UGAm1cIVj9E+lQgxerVj2XgijZgTkYelg
J/U3e3pqezE/Ix0LvGuq7FGSvm+qo02W5q9HjOfTa/TqF4JDDtvrOVg0EFlNVw1t
2VMeofdtGTuAfrKeHPzZScf4TJXNV8WS3gTaPvK0WXuf7C0taWNJCWrxzzQPZqQj
3QWpljdbnHO2wpAGxx/6NmqNc4wni6bHv1oCkOirQwTPogus/VIz/nFgVa1+vPYL
xFfM6XUpSx6PIKHiMXiOC9Ny7DFIzAI+tBb6xuXMYppBsfgNq3ZW3LpYpWLeNeC+
n+wiCMhipQjKC0Ich3scv+3S5S9f87N/qXQYRGaKlHi/M+5QtCa5wciuBCA4QbIW
spzt4BYFGJNDxjCujaNh4uepAhssGtCq++p9zVXZf6AVspq/3X/sJfgyLP0U1Bj/
s06pyYtmui+pjtWLSp1tA988XAisR8u9EkPapxc29u/A+KucZBcTGe1VbdxZaceX
J6qLNh2zpW10qYxaB3I8IC7eoQeybWXjiu6135Sq8HOT3L05EEkm5hPyM9rEK7Sq
ofTz8n6zpPqO6q9ZqPfE3vDDN5izj2kj0Ccu+8srYCCuUK1bnI6q5Lntolv0Bfuq
En10zFCFZGkIh8FLUdws7X4qIrGm+zJ6U6WShex5SYiPVV9XgC3/ZCs9Gc6G7k90
L25Ianx+8w7VYSfGJvNZitVLyghwsowFfHwWkPZMvO17vYB98a3cTZEOodlraXp+
XRGmX1xBjJYKx8nXBQsg+7XEjv+ZobMuzA2qtmdxGHgepbpNDtPwozccwKtqqPPM
Z7AzIXAJbE/saagG2ur7uuTDGT+wcHpkkGBiXL9csNoPONoAH48E/cmPhxOPMv2q
3Z/JC1hz3K1k+Fqj9+3ae8XboPr4vf13/q0bmFAHHP1UqjTYwVXlzmTEQNsLNGor
kR71QlWu89cq+W9waSvatdG3sG5bXLci76bXBsefBMq9YmpWfMpfRNRAS2B90J5+
fjMWPLHQC3Rd8mKBFoQvCNyTMwmQceooEoM0Kv/2tWMENvmnxXszha07BS0K77/e
fDEk5YGRA3zQKSZSYaPV2B7JVSAv0H+UR/FrBjoEzSy1mxTJFlSxVODzE0kjAsus
zEBab+yzehokOvvi6G8Vzkj2DpmeGYarPLZNJmEg9//riZ7tdTa4H7YSwPnaALTO
s8+kOlW6yRAkc7ux5jLuBh/e9qzCzfEWZCczKqcQG52WSwWjqRv2yXLV+Ey0Z5W+
V2ABd13M7/E3dCcOLN5a68FxM4xFW2PRP/zodGSiEMyaN/59IOqoYXaU4Dvd0PC5
381GpmIddtza2T2etB8sWtiN9HpKN4bzromotZqZbwP2f/Hm+e2spuSO3GOkgW8g
3f3F8/EFYl/iSbQJiXAG7iwNudrXop/thjMS7NeMnq2lFdIbBmhiYXhRjemkyHjt
u6YqkdFyw9p/u1awHKdVqzzFjUZ2kXim2giHjY6cqjOtMGU6BFEVbAIzOsWqzUw0
FFI4qyLsiNjcnOoUac4KbIClyc+xbrVQznb6Vu1KsMkJaBc+uYiKG9BPc6rJmah0
g0/2qFf/daDTTwOtiwGst4l2OXF9OzKdaQYVaiP1eskO0TFCAAQQsPjB/T62WxUF
Gu8NxFG9YetDhZSkD9EZPz2rwAz6aGf4W9nndZPBOG/aMiP0ygeS43N57rm8GUoS
FWHtrZON+6m74qVt2exPwxn/VqDYj4elVNw3jPSpranXFbwdsZ3JcuCTFx+bZvhM
mHli65gRnTJVfIE/nCk1qBSlvzfohMVW2R+QhAYvUfjvfTOwtcYeGSq0LU1Vo8BG
4T32psjcInuFzous3hwQQwonWhjcLC7y0fGzQrEKfA7gfaZa93mseUOY5cN+a9DO
mJcQE15TQIPoNcL1uoZExN7FyRr6FvPIe9tTt2grRsZ7Oz8dkbFpcWpMEY5Xpxxb
Ep8dirOGd5Xny9B5ruXd6CSucLNIkgvmc6+Ln/oK73q0nqVbFRCLXTod0nrQsY4W
oNyDl9d5D95SzZqCUQHW/8fBswL0n+a6oxwyxbhwGj15V7bd8pAtY3/ilT8b7ayF
7xFes4He3WeM+hJmlik9M3em46HbzfVxUGpZmhfoHJnVvH604hCv+tc/EorJQoK8
+K4fD/wl0J4F6jPA4dNT59ucx9EWHQtOHjXENxhGB7JEKaL7iqwd6Fa5JsANshcx
JsPpl6P6OyqqB8dlZurgKyFwwhYDkGhEQoXBUv685nh0emFVKr70YXRUbEPyIe2S
OF/Kar1L2HlbC2qYDUD9fOwJ2eEIdHbt7hou84id/jnu4CtSgSq1JTq3h1M5gvb/
PnxgtTQvmrul5+2rfC/oypVBPd189GsJ4L8cV32K9/FRx+TbZgPfnVF+p2NAYyDG
XZTFnq8QYT+/FWE8VKT2zVEWixbYCuy0c9/doG5+2m1jbaKlT1AvGe5wuZ55eHNE
xzHs2lsJi/sNRjJgFj5QOMJL4bdgGYuxkz4NJAeA3wqFehzdcjoacyKm9lkxxpsv
AU60mF5VIP9tFnC9BvTHIwvwj4f6Oi11h4HrLk0O1FZX4dkadtDfLoWPOBt9k2Za
wOChtbZjJuw6/K0uhkERoegujqd9VDy0d/5EVKX8yh5wnDeNZzlp7MyiceEqJx2s
xbxnI9dU6ImzX0yGMVjVjuu4uB/7qUXM+iy2yjtySSFUDTq/sOl05Db1Gk0W3Ufa
VaR8U4dzcrDeDY4I+AU5IGWGPCN7XjB0lo0r+bqKceGBlGenl3pCxgMsGTPGV/N5
miaMjrS2UxpFF37CFjTlvWZ6N/6WTufv1k5bWetAzpUYcXAzwVZUzhLItRwse2Ee
Kb85fiNylKTgh9vS5k8sTDPspkpuf7/B6w7pHUlFFynlX2geDSc/V1PMkJXVouf4
tn/dqW9H12PbBWRf+6hSbYVNx5m6ssMuC2NL5/9WptEojDLxC3JgD2GPVOZtcFGO
WKmDz2P/WP9987E6562uWiFbZCw4uKUEmKnAS7moL/ZMkZxkla8Bi48pXwynsslP
S01UvuFqYoje4xbLcd4V1IQ+vpOkc66cXbrl1zEn+p1v+1hwf8xcOakbrPP0nde0
TFo57HCQG09lG4bBsHjQbz1WC+qqe1DHnUG439DFO6kkTRJ82VruesNJm1FveDsM
+VT4C3wTD6+49KtEiv+MU5I6l1Xr/g1BOT45aoesGrcNnXYnfR2KHLm0q7RIGOnK
fgLbXDT06UmbfO+AKb1L+J18FPNgKa4+hDQ+lC/tFagiuyWfzEcfsoqiChzDwPfH
nrdWoinWJ+WaDco6WkhOo+cyaqh8e68QhZSo3fqULKYtMKWtMzGPtp5MXNTZcWy9
4pQP/dbNw94hpoteRIKVH0puDqAfXLOl86o0Kz1Jm+Oa0RtQ+ncr1s9W6vZ74u9b
dlYyfJ43bEeJ5278iOuLy36fUAhKLyXCTk/aeLwsaPyP3YEbaM51XbFY85QAqTHo
Q5BKmdWFMfmwpCvFyJR3Uk0/zHd3rnAXiifdToWdCKLh1HpXwR7nG7u2aprr/o8q
c6D8GwDUf/UEfy++7sCEkMW7ctcbwDxFBwuj8JHo3QF5Imhid+g/6TCNb2r9ITFN
uqrL/a1Wd8whPRDzheFzvQ6mH6do0bcutT093fzYcWieePWoq6q9Tret562sTQwx
8KAss4DLPWd6rwsfarYpuX7tQgAdRT6Mn8dtKWpN5MDIhHKBMlx867HR0Na4v7eY
7YwsazSn/tlK0S7QW9sKEqvXASBen7vPEVzpwCgTUEGchPsN685dGTstjgi+zVof
NYRxWho0WnI9Th4jn40GLlqyhz3qgdsDFGZqQB7tuq5DmAY2diMaipNJmadHnjqX
1fezehdlcaueqkDY2uVsOrf0vCEQxELsjiQHVPruyZfXDwKcuiYTk0MM+dJ9WYMr
jdTjBJPBbJ+TfxToPwnxPfsbgaGf5zv4watOqAjtUnCrODXS0Q6V1o4K93+OcMFy
TkHBRHFu3gyYk6E72Di7heDhJr3Ci0/3fr0OTGMTcvgxKpWmMNI72+V03ysWetsN
iktTGrKS7PSSsaSqGvu1XHIG3Qrsqa7LDFSjJPlSmuuW/qikFlVYAnVr+Z1FXtJ7
x/+smVK/LxMPdEYMKWnBSJ4S6FywUadxsTJDGZoZ94U4UpIANibLgRaYUpB0HmVo
NdcUdXk93ryakGUlp7/hS4GU8p3+6KBR4yAD0KPZ5juMIhW9tBtyt1RUCINaioDK
cPOjgxDjLBLBEHb6nYak1gfkVHU9b1528+sH5hdA5isiwvpYoyweSZZTNSAqYVzz
BNuCEkaC/6eqtpqVXsYuMJMzCUYzGWEzTSUv5vy5foLh8RJPdhFOtndirxdRELAL
VgzruWWuio7ajfynANb6uCDeOQeLDmRVSUqQayFv6pa4bT2V2pofn5Y27bhHn+JV
2xeG1FcPmyodcyY7sJ5AobBiH/eAiUwn3b1+rkw2k5HmGVRNb2evOdAAe8Ofk0pn
c5hG4/3Db9CPAd8vPu3yVDGTyosbYwhqCxZdGOWKFa7GXzrVTHVr3wIIY3yOdOgp
yRrnSglxhRe5gy1obOewfT+NGv8Bk0Yc+JPHq/BJ6wnSOCoqtSZbfHxf2DEX8buH
bP0SyCRq7zZHtE1fe2bUVFoR6Tma3LJ/ySTAT4PnDag2+qsQj9P4tyBdkjUOAun7
AYp10y32W8gkD101PIjwC0CLO3e5O+vBqxWcbnin2KK0ZfRSRnZCcRDfovg7mANY
zXkXAnWdRtqRYa0hSteFe4YEgoskfm6+xzQrO4JwPi/JX2u6NAMRJP97div4rntQ
gA02lSqmkYr6b9FHhn2IrYZgH8xvfl35ZOCLGBButacis13Jck2okPKOtgbEj9wg
F/DoY48rAHsztUqHuDLbW6x8S9H6Yl93IIx0BYOTOesduVmfMBIuCDT/ZiPfewCK
1DVXDK/uQ5fJCEWItlcy7MRMVw+cSd8x6iRtZcUlr8ZJ624Tsrt2duI96sVQmi/x
JG5x2ShOTGkplk0eSvtWmI1zPJzBg1uPGrXJ3dggGb4TYs1ztwnoU0QG3nLkjgcN
DPNS402HY3ClccYMrUyLsMLBp9kWUjLx+2g/naA/l4L/uzh/KQiJOdtQT3PWVpW2
pCGmsbr0ue5K5jefvOqtttFMcaKb0gPPI2eNzju40LCTvmrilMXE8kgB1NMlPs0e
k8ThMxUPIFW9XiGJFLmwcb+Ca4hHZ2JE9mhWi7NIX/F3rOk3lUou0DIZ+4p4Ttgm
pgvfPPajsFPUKlG4MMCYVqdbe0o6qMLDyVqeRd0jmopocKQxY8fk6x77JNJYrlvt
mw9nVn8GbhnvvmwfPHgmfgzv4KMJFxXsmuh14AP0Vqqs82iBv/rV+rxocfz6GNBA
VZ4brFPy21okj8ikaOpeixT0BbOE7Wz2+mNxy4qINgQ6ZeWjHtUkhG79NzDduvMM
cFOIXce6hbBprZOALVIz60I1vRcx/a6pZ4u6g5TWIjbbYGl7gKyu7+Dlox0Feofp
T9lWUAGJXBkbIW0zdae6k+C9oHcs5liPyOPGu66YfeUYQ4IbD3fO4awNYsokc+B/
J1UgDDVhEa2ce+KZ/8Und0/xMMIqPprq8ZCbXUf1gh5+Tfo3DdRYgHMkZY8j2y7g
qeSfujH1Wp7u+S4FKMBOD+ScO6RgH+WzpDgW7w2PWn9czLlb/o9Ew1M9wK65q1qr
vKVpMgo2wBLISNtzp5TFAUXe1urxQYhbc0zXZywSeJ9tXj3KhcMGcg8oZp5arg2Y
qacbwZtSt4p/JxhXwZYa1FCA0VO4SqTT0+gT97JiBNd7XRRzX+mv76Wja/LMwWBK
BzRt2p9P76Zs8bjCc9vJU6yZ9H+l+8rrIIELBWoNFjeD1MAG13yj4XLvfiTujWUA
36VJLPRpNLUEqEY4Evfzuj37XdsSw8oNUGPty6fDIdGXh4mmKHMiUru2IbOy0cDr
4CcyppmsqF1yBlA0PwDcGc4M8w6VSfddmdFGIOHmwNyWNVOFeY2N5JgbS2uBAVgR
i0VCHd+Dor2N/DFRIcmFcv/1LuWIqjQd+vfONoQ1ylFILo1/63Ll8SaCZ1DY0TVZ
OJrc+tVbBNhwmOifC+RwKEVzJG9I/lSLtnpP8ExBo4olgm7T2z2tyrStYZVTH1MZ
2h95QsW5wNes4F4nMBUWPRDI3gMtjlaYfY2s9y6GN9Rf0P8IZmlVi+FGChijHBFG
jfbXUjVVG9/7VlhAggtxaZJpQkXuYwI51sAGB53KzX135VGc90NXqspbgsO6ziTs
2aF18kifwajDEpS2ffY0n46DXwDveXh/KoPZd0qWCVab3BKllwgjlv3V7LUNdJvf
sR5vZjTJYa8ekmOo3zyyb+qL14r5DU2FJyBGOBeOyCGpzdB2gfiYCs8Cfppp0iuQ
EnVUJR+ZaXg1I1AmFOWT1hdXE7L1oEEhIdx6fIusta1sNWvQrwhjyFhLRZx9SLHF
DqJiNZATYb9K6WiGyqskJgodQSJELoJMW2RsmBWsHTwWWNNgkUgyrjuqfgEKM8SY
xItyPR02SQ6nde4zErtYdRxQXawWWCFga5yeXjZUijTpQl/p+Sz6MtAUs6m+ifB0
/LDzjgIIUcuUtJGnp7lF5+9YOxaL4RMuk7Hp75NGt4isA1g3txBcb27XVHfFJn5G
J1+QOCGgVYYJTMrLls4m+dQCPayzTOvMbMZzI0Yr7isf9pX0e4LWHyjX9hmOi/VM
d6c3egobZYbrGyqDlX5ospeujgkCT9K/7jiHd9HqjcIl+3omgQeEVynjH4BLO87R
cNESbV7DlwizeTrpdvE1zzUvk7D5Yu7TaAO5QjkWvcD7F2KmKFql2YJbHQ1UEVfY
mrqWgpfxfwwyMVHV5CN3mhTHtoFoBuf04Nuq3Dsr9HJvQACsE40yAOh1p5V7IFvk
ZFSXVGixW2+zorFEkb5kpXWAcPxIsxMyKxTPGpBUwFN6DCcZOVq0svAOHZbNkkeM
EFQdMxI7bML+q/kUzeYMrN1ChinztEEsvc8kYxNLl5MVfmXFE1a9kTbKbBdsYBxE
ULPv8+zy8wbS0LLrZqMf5vjlk/TOaJXvSZlteN0yZ3OQfy9CGkY3pnqvir/Vp5YF
Fyw9Y7yltIG3AqSGcD08mQALsQvu/eDKjQxOiVFfSF2gcJRfNeKbRGb6WPTGNIkQ
ir1IIQPMi8F6Z/cEy9TvY2owbT6xmMqPgWcQwjMF2MsaT31zmjImE0O/vFMbt7lJ
r8ykOJwOO7p/XkUIf6zEm3FvYMXfj9n4mCjzkwmzflhyS5yuUx7KssOMPOvyDvCH
mMyRmUkMQFgX91KyPNNYD5rr8Q2VhDlTpycgXw8shzvPPM1ojbba165CrPFhtVNi
Ercak7/o1yR2D/g8qAYCr4+vqpXPAthxqO63AqOCfoIKC1BBEacyP3l64oWh8JZy
Q7Z1Ye7c0aZftJyZ0UirswDcLGe3MXuqWSYcfe9BTx1lxh37azQH8GX5FY8ISmao
BWsG9fBasKwVwGjviUQMKaJqSmZyNbbkUkx459fphR5qSijsAwXBebhVQe0qVs9C
tIfrTrnxHxo7ypyrH2K5e4cNo8SSqCcJJ3qvbCGRV2sOss5GyrMRK4voyKUfy+Z/
EDt1lNCh/hkZGQ4jreIMMNSvtnLPm4BDyfwGaXmoBkPx8o3EMwN0WxIfO1sITGuV
37NzBDmpZVv1vkRtFmsDWi0evkhwtBjU6r9ze6Fii4DGGBgwB7keIn4ddk9zkVCA
+BrmZBJHFNSz+ZcoPOuGo09DKkVjqz6cLGS4jlVSzdsDLvwWb31UZsPiwVgoJ0bS
JsOenlMH0rqS+5ADdNdgCXFdMyAXQfB2yeaAwTlx1YbtrejQl4+IysscXrKfl1ok
/4Ibq/qi0m3nHmAcFwYMyBslzMc1LuwfeQ8hiYJRmi2Q8cIIZN/mDHvy/uqM/wML
xsks34SN3L7OYvte1iqrjAOyEAhrypJcEMXOyCfP3pgHOKhIjz/wOofNNxW470FD
wVulTHap/fItqy/RvllmtZK+c2dmSQWRoapjIiNzuCvP5TbxrYolfW0HYrkft6Ch
sAblTU77sdhBFUp8Jda34Nb27THbVxOJpTNZaR5w0Ef/HuBfFV7IgyjQMPBPf54g
EhTJc3PWWhDgmKQa8ElRhdv9UtC/wMo1qCef5sGqbESO4nCQtaHQB/AYJoTFHk6F
zPy2KTm7EKd7SNTaG7KGpoY/1wQgsbpvMftzuieNiwuXZa+5r0ssdN1FALfbht+B
NPpzCNocduXCfwRbKsOydXWPMF9JFyEXjds9HdReWO49nbpSosY1Sfj2woO/dpJY
3JF7YBvmaBN4uJUZtuX0w82wX69nxnK4G2Ds1AiM3sGlutCRKa09rTZhSMU9GquR
UhNeFLcg5sKMQsD52EebFbhKmVKm5BcAqNChuUarAsPbuEm3v5QmDZDTAHIcZwXO
muC388EPpV0VrrLj+UbqQRb5+IqOL0Ujy1+exz0xPKWhFIA8Ui0bYdufxDlBPYeL
tqe94v+DEXORP+fbrJR97xt81yudoKXGvCz3ejhwrBop+MKbfxo2wGjYnHNA3EhD
i4ZXTm8VQ1eLA6/wCg7ub1irSvaNHwGv/BR8Dfe+akmVl9dBd73JD88S8gIOvQDH
QtVYxn+0yYMf14DIoSVZi1ieSqZuQAYtO2/NMU968PKLMzIZUnWKbmsPZCAThSt2
Prg6AW2bhnPLLWDcH/pjOfUliD1ocaK+Lf12MAQ3YfbRB4BkRUB55WmxaFRLI0kh
soPIM6/QVd9X3toz7CcLc0E2AQDtd9kPTIuq7Jn8u77u7n1WhN6dmKEq88ZEMejt
QhFU7OiZ6FzKM/WlxjyTzbi2TVeJW3mQWX6y/H08oPu6PgRxzIQ+4bhr8uux/jxy
qyIVZgew2orW82jQp48QV+MVl+7xqWzB1cdRU2YItvDU8ObhGwGxxsMdLXBNdk9n
a7UK/HTbsFer3Uo8yhXLpN27nEFg0nZm17gf0npqrL5hsqKgleYb0JCrXqh85Cd7
FGGXiLKihgJaNAl8YzUdpX6s+dl8+PJVf7LZBQ+vMfTRvhWmEgwiM6wRrmOjx+si
yYLaahFQlHorJWL7U8JkkcOCI9VaWDxr/6EzuEXz9DsExWt62tKY8JQcNqG60Yqo
2ZMbdW6quJNujOuSrn9hjIYOImpBm34yMQ/adRI5hoAqRhzX/G7QptxIaBNZHksR
385ym0gWaZ/k8zodHzOzgC5jl6BNKefcEojloDnAlSAqtuN+y/m7yhov95LdD2ck
/xFOS8uJTa6yx6gJxjpOaKOiltBajELcZb0QyPCFbUrWM1M5Sp3BM3gKAeOwP0jY
+SRxrq0cwRBHEGJJs4qujHMmQiefO+KkCbS2rKj9cmA/tN31iSWfIxwpfRuNPFQS
5VyFVYHcbg0XWizCr9NSNwFmmsYnLZ7MqPqhwf6iZ7wBJRoh5OYcS+QxrHZiNyKT
FObtMgPH+JmyZLGyd4+s8PpA7y6zKFN44RDm46gHpj/K0ngM4Iq70CiBKYCHDIA0
vNuY8K5dlsV1A535ujUJQ+Ynn0w7H+9HqKtKEIVfgX8Qv8JmUg1gj6qEImVf9z3d
YuOZEDsmU3zvaDGaKWEf9+bowzsH/D76SR2YAg3art2nAyBxIRZJY8pUOHj+cOp8
+ySDIel0R9zdU1l3V6H2s0Jpw/v1lPhUjxPprddIDPl7sxAqEVyRGaIDtZnV48oX
yb4yXOvgAPALYBUrw38mlG4KasrFZSiHCN5S8KdDnYG2G2LdfLD+hHnCEHND58Lj
HcEZdrui+JDRJsfKHJu8cxcPkjQR5d5T5NJQ+mklaar65i6xOSor1lCi+uphjI5F
srf9wHjdAOb4ndfJcX0GX5Q+nvP37aLVOjjEVK/wsTLgmyeygZ6FL8O5QJ07Lztb
GsftTIBIPb9TqtLpP8lg/PoITH8P378mCkX53PWy8aXPsuIPqFb6g442OuGC8Udp
vM1osv5VQJ4fEMbdNybRqJ2tPU88qsi3o2Tvm2SE11qOz12BmFpIUFXHPLJo8yJm
PSsBrmFIh3C0/d3VF7Yma3YS0j3u7zLO5JQu8AiQUM1DJEq6rMQ/7SZtqKe92+1Q
rZrGm2ffqX+sACVD+oGaRyTeQyjnb8HQwQ098yfHj/QKHAFFv/g0ERZFw7WiwKO4
xtKfVk/aqrgqW5Q13XK0XLc2AQ9jFo44VTwNZzkHNmToNiVzALeLT1FsGevi2bCL
TEOLgkCjW90YHZ/z130qCBaZ1lI97yh9VlMuDKcB/MOHe1E2HF7PRVCt7jGLxRU4
makX1VvyCU6lbLumbPbAJ7RueDo9MvHB46X9YhyJm24zvHlWWRuOmPR9FR0FXbp/
YT+oeWX/eEyb10KjpjvOw2/hQzSkjSyi+cQjCpdAN+JLHdt4Em2DjONul5x7LkhF
PMwI/hjdYnhhW5DjjehfVNbc3DxqUCIUFk7D+3S7cPUGYQ9CH0x4GLJ+b1/aiwzk
x2gM+1IXd3112je54lyCD4suM06oir78yw0mVS8o7PacZ2mMj+2TOTSgLERWPyBr
VnYmmH104R6y4CxjoV8AKjvGa5bGDo/USi9yTJTA0PwJiiORCI2RKq668eD8kKeV
4iVEcy+gyWOrEgFVvO4eLGbDr5dRwpL1I66d7BRo3uaFYaZm35hon0qLkoRYozxF
MgLVNU2u/0XsQfCeOkU4jucaRlvflrLVfxr/gbCohg00SNbEVnVpo0ceL2buB178
P2L4MENH3AXVQf7Gqh7THIy1PvMyE/zOI35u3Y+UT8NXi55DYWCc9xqlp/2trMLn
Cw4Cxvcr291g/IsyrwD1cdPLdoOKvw+XG6VEVM8tx+bdXQcdMqSuVoDC40NBC2zq
diN3GjpRBqtMygAaodGP3qIGTIMa+O9WXEahh2ZuDGLEy03aQbQqLf3QCmhckVh+
AYzCcZ6rgADdtPmZn68dLTRIl4z2bQMTwdKiC2PItMnvHH8fj/iv664HYkc1YK6W
3H+jjXqMnQSPd2ebISbenEy8oIbAdf0bNboqnToBLnCx2c1N46/ounTa+HGOrHF+
CrR78FuMdDeSf0BMDClbxdZaN7rCZ/9KklOnTh7NhAQ2ZyTQA5rhlnNDFcDz8WUX
fW3W25GEVuzr/qBWULOg8Oc6cGIQb7kEYSyvWM/rdpS+rGcDCMIf/PRPe7LrAXmK
FAVknWbgO/SDj9lkrVYJtJQbWfN8OSpVRTRufntDisrhxKTUs6sBQucs1r9WV+gQ
DZ0mVyddbs/5pdwweILPe6mujYwqpSvXVjfsh7yUrwDPLXjx2qHCjTneb0v3t4ZV
Pc8Th0AwMw1BFkZ7EcV5s06RbxUuAXQ/qroog5u2KaHx2dSC8HYFu0ZK0SWfiUbM
Zbk3L/JH5r278qSYeC5wRJuiqxRuClvwHNcWztRBB4rvNb3QB8dmZAr0afz0ikqw
SlR957RSrwftP0FRTlDm1mBVIkqXvIq4uLWlN6rVUT3VQomedSpn/aKaF6cy0Hi5
7XxQpxNluuMDUV/Wu8kxKGiRKGDh4z8zQAuBAb0jkbyluUA5tSfAb2F4LRWNrmn+
XYT1c15OlIcMFNG8ng988XD2thq6/miL44pxZ5q79utJ9gnU2FESk5KEINpRoI+7
z7PyZIOqYpSYhKHqSMpd2wceIyDt2vsw2rEJA5JFWMIJS1iMNwXTyShdOImsh4RS
FyPY5R7WVjwjnfio/Z5btM9jf3YgWauVMgykBdJFjwUbm29IbYe9Pgc54eNsew4b
K9ZvIbmGXZfKv6Frl5vEIEylXwNOaZ4R7sOfuNL+uWkXw+s+907dCaWRi1y9j00J
PF4g9LxZEFc5gk+JvOfavb68yuxENGE/SUrJgaJIyQiRiVe//9gQv76GYQztptEv
p/RCjS5n62H3hdANjo5AvHXDBbBNDjmxziaopXtCwGzh2Jr39oH5v1gdWmaBYBJp
jYx4IaegCOV5sk36WuOynU5iEevkMqCftMdH+TToTmOVPweV5n0aO1dNjdtMq8vP
5HoShM+GmGOuXvlS26EHwsKloO6/xrRYvsYw1VWlGLmQJgHPCRgHUM7Cws+cdkCt
yO65siHs/LulNGiC8tuXM/iDY3oOAjBbHizPpRonyMChjqz6hhspKCnM5Dtu2jXb
ueh/i1GunDf73dnuxl3vNxE7f7Qyg2FMxzcgZ/W3oDKrHD/uj+zElXPf9LLJ/myr
t0gGv/iJyK012HeICFBLfGIml12wAc9bHWXaADjMRvFlUiYYM49xLgQvEOViCQ2P
Wh848TAyzYxWOTtOzo7IPI03RzP6qc60Ue8JU7RVyzz8iWI2oiEjILpz17aINzGc
zZY8D4Fa7G9IkGl/wP6Fi2cZkpICMeg4REespDX4Bx96sYXflYY7Kwgu8pE6x3g8
RfdoyALlyivS5cQP28uR04ekWqjo9kv5a9dDfGZoeog8kJxJnFhQjCXsDMrbaxmQ
30yuQDuwxDAQeucfenqDKg9O043xhEIrvozPbKZZ6fZdviLguTO3WlhqoBSOHDWp
Wh9xZj3DeF0oJbqBwmcXyNWH89U84uvQcrBuTot6ZWh4v6DT9QCyl1+pi2Sx3nCR
AWrDsDH7r3hpTLU5MxiQ5sBduxpJxOoxKSyhHIDPr9uIOQkmi3AQQI2xi42cMQWc
NccRAFMVaTrgcWZQSFymOGNpUmj28JtSwTHVV5cOeLmDONxOEUfzdBV/7QtGpY7f
hJ91/YvJujdzI7f8jbjQowW0QQIu+JqpmonEJ00iFo6j6QedHTiJVJq3wvbsOyE1
47dnLtDUW7kmq0ecFhJ97nG3f3tSPTY6WcqgMjV/DZLL6/TLX71jPB4UJPzrjjsn
6kXt8QGbcB8utobYuFl1s4R4RmUTccBU/oXOCE/n+YJMZvpaQ+Ga6fUSXJj1ZATi
iXCOOJYkPJTV3aQk5AibUgFYS8rjG04W0GEvplxHB467tQJYjdN9Kf39aYeD7OnV
L4EsHMoM6sucrodjC8wKfZ9LAEj0NGFkaXD3aNlb/BPv84WqF/t8W2UZbP6VnqoW
1E2xUhOWmL5dR/Q0AuhZCYtgqdDBwgr4WXNCb6eG6KbIaM787RYAPAgsS2RPicdT
phKWgFJUos2iJWSpfwprN3f4Qgruz1kSUZa1SDn5Rs1j/pMg/CQaHGkHoDrfCKMv
wlSOX69aCfSQoA9EYTmOrp7WC75O6VJLvqj7qVfPZm0eiZZ7IKAMmC+WlML8YYhq
/40qZW7Yk7+gW2qHlvKmBEwsy+smhRzPN0d+CBGtkltKG1NUxWzjE9MbHYmSFi71
OlHF4zqu7vys+d7CxBe1AY4isj0SIvmW63u6cXDVyZefI61V/uIbsCWibldlt8QZ
4501N/r1QF5b2aDKoMv32a5vr9TridK1mkhhXLfcuSGFj9RVDbo/PK62E3YycTX0
JYHrx8nvn5ZW+18n4R2SRPOyftl4l+JhQmwthaVJJ2lLfUVJTnFOpOGQ0jnFiMDK
hPm/sI2maQtaIuGoaV2dsS4NF02BTG67REAo8lQW/Y1sdtbFpw7Kp5WWNP/njUXP
mCnAOOsubJvGbHwHolT/7ziHloQ8ZhEq2iSIKl1BRJbLX0YP1xiKtaBKs232Pwrg
wTXxRxxi/HamwSRmVZcHQMUo+1FJEAiJXwhQBo9taiYfGzt4xvi4nhWGLUUFjgZ5
4H9oiTPKJf5IFjvHh6hkZJoeu/Yv2E1JRK1e+NOWlRllQQb15ORbG0uUeN+Zm3Yt
jKiqmwjLI0J3AcJDWXNE0LNAiiXZR7zLIW/I4vHNsaUIoyrOILvd3ZJeV1WeIBkE
kL76m9a2/+Quz/TjehIZxF18cDTYYcz+5DtuK5fRIjm+62U/SxL6nnYHcJSEtmFg
320Chkbd1vUxtwksXb630MUN++KNaQxghvZ9lWcmP1qgJqE1LfuWkrhUYqqTvGDZ
TQ3WkTxf95vwcmwfJmsk8Xym5lVy+m0RY/ovJCBQNaFILruHYMywAaiNhBpmb8SZ
YgYkCTt9ugm9mICtZNchSEDj6JeirL6u4vw7QJgn25Uz5A+tNjGqyNC3Hf7Kt989
37WxNF+9T2GkwILhZsohFxv7bBtw3PeUml1txzermBtQ1KleTScXGOPTRf3mdQmp
BooRy39QUPT+f0PLB72e+k9HirgWDoGGgWbZpyEAOzXi//t0eboyfGls2BzKekZ3
UaONZOiU891BmeW9IoXVfoU8yH4oCEqlswYCdUmn98aSJv+rs64q0uGqKyruve0G
EEBRZ3Zz6U32KXtM/TmA9jEMOrRl0qg+7RydRb+fpn0zGHM7wISorhFJQdYNMDbK
ht8GhX8itXIoTNgmDV/C1TaUC6c6G1XghfV6mYQ1VQS0rGY/X8wgrIeXIjb4Cyhm
5LYf7fuGDGD39vp4drhxXdFcub5Uv7kBsZYW+CwjQWh7yhb98UFUj7tQhViLtGZz
+OWrWfSotrGu8KjVIY1ya5gvsz/0CMderw77NUx78zTac3twXQbQJEfEpYucAtqp
lYDlwmRhRFzdjMzkNlUIZurH3TsvYv7imQgyc2zKc9jcZZGWp+v156JcxGzlo9r0
/6HpA3svcnTlYw0veoehUFR+xlzkstBeAo8L0kx1kfU9qQhJFaLFHZOZ7lgaqV2/
tTbCVuiuuOtiTM7T/JgHeuYLyW91UL8sW9RPbbkjTeCrCP7+7kJLrbw0cHpqflUC
D9YaBlEwoM2tA+ZUQW7xKv0CQJoTxxJtYXdtIhtihI+yTOcQpt1Zsrb/TK7/RXb9
gDaNQk4jnI/DSClGWQT6oJm5sZwuL+X7vgFZhevz2nLJ6R/RdJHAJCMlkgjvzIou
7Ga1Zm3IKYPhGeRTdRevFyi5P6Wqk2iSDZ/NlhhJsS3AYvz/K6a9Nuzy6QjhagYO
tXhpKIYMDvj1Sn/aquPjIEZ2edIfpg6suPVV0KbaSc1f2HvrB4K/ySOk24WvLkqo
jVu9ETH5t71EhBmMexVkug8HwLXg9XBj0Zrf+hJKT55anYftNqZSv/xlnTWGY/hV
KvVnRGKyt0iHyvB/t4mWAZt42dEAevnT9CagQ1U+X49d9wuo+8BsaGkNWnmZr+Sd
sA5OU5Qtk7q9sJ2YCR/c6A9qZ37Gxc7Yy3GgImZ0YudLlB5mohvcW21WbOhyZZWQ
yqfs7mR9AisoScbCu0eczpiJC356G/o2DlBKYd063NQLTNCnmvBS7cRbGZ5qnOdH
FpcwIfwjP0ysdg4m4oxaCOcXRNHjshGUkd80DgzWmEzQh3ZoRcg/7Ti5ewYgeMTm
gK65r4XOOwqx1rWXI8+LOcBiLYUnOqiD1H2em4jOZnb/L7XFh5E1/hDaXnTcOF7e
5sljYVZUb5+3qV0Tqx6HaTZ/JNE9vntyz2QOQULGCyq+X5xD/EPknPcFekniala0
ywZsNSJcR15YJ5ApuHQ3Z0sF9qWNzl95yxiWvUBzUrIoTA7M+L048wMLokxMI5+e
0N3OxIEnN59DBVP3p+aaY8oI37GmpX/2/46i0/FD6V8b5boxtmoUAMQGIqqDNa4d
wGvgrEpmb3bs3GwCUKzNsdApBaYH66nsD1LOe36XKIaUdl4OuftXnMbjesXEj5Sl
X/q5WAVBvpRstYFFBCcsNcBf68jv7G7/iLSzm2YNBHVknADcOpVYnOqwb6TFvFd9
Rals5gxZ1SHMi4BzzkIedJ/0corbKieg9CUaRebxRXhg3FianiJ0fjrJP32PNq8Z
jUSuONALkDKzINq2hU7+NDd829Gcbs9PN1wHGCnUacakn4LvZ3J/2Iu8CDBtzMB0
8kNo+0B77LHg+pisLVwscL7m9kSlTHGrkYrkiLTx31QilXPgZYQF6Gu0w+dkOyEi
V91waHFfCiAhUte36ZEAVa+YRCvqk6R97OBZZs/Oo4U/KJY4p40wu/GZIJRl9q6L
Hu5jPo5NRu0GrL5LsnXdIjjouBVPgGav3eYA3cXPI2c4vMoubAxjQs8b+baWkoXc
9NLwtUpvNrwdCf52yyzLVSvQph8ZZ2V/tSwBhFqjEpSGMlEWgk9C1w74HWcGbRR/
uq/kzwzSlwn+UAStY63pUAnan7j8hpRqlSTDfrDWs3WqbIhh7yle/PV861xsV/+q
XjlGhx/1TcNi5C1W/Uu6vmr4IUKjCLgzBO4Xt8kcxs5BgLBY/vEnQPmfGoxl9H+0
oFVv8qpH4GY7nZR0n7ZgqPLsTB/s+unsuHiU0v8+NPageqIRouSuOG08EEUVAvw6
a9k5lh4SkoRU3eWttKEAqNhmrihpAzE9sWF+ViqtCsV6UfgQ1G1OJoNfKMMarRxC
62iuV7ZjNQzsNBMoa/LlsNdJYBorIDp09/RK6PzCCNvX53QOQKCTntNWYHu9841j
Nh3Dm+wjr5Xx+hia+taintdBio3HZAvYBQPUsO52Chg/iHJhE4ifjGboXqbZi1h8
aILT3bqYG5G82gCCxGpjJbsQ45Z06DIIGb+L67Kg6NtUVTg1/+Scs+Kz3WdIKGug
qSi3swdtUchTfHcCJhYbVN1psuY7iJmH8dumssDRdptgv3tEEalfU6ir0MH4IOyK
/XH7LbN0pzyWdyV9B8rH5qSxJw7ap5VjwvWwO6GeddJf5VQUQhEMbC/nG49ZFsPE
izQ3TCNJwH+xzNLTXg2TEc64xDyGEMMscsCx3IjrYGjj7Azaya16Z8bQGpYlMsKX
ILP+06byJxKvAxcKCIW4S1BDzwrnEGY0v96rC7L2a3w92WYAIodSzMZOu40nPjB4
mYK2GTO1IvI6xvKBVSoSPMM/gDJnAUeuQnmrTffgjhtDvYKYn8Aje4/ZtTOFCUIv
Fh47KLOV79JbY+UyYNul+VaDCsb1DgHlXToGGZlAUaA9rvhL9h6D7VSh3XGyrJqY
bFOSLxKwFeroQblQIrFwaB5OAmHPUURPpuFrvRy8yZpATOANt/j+gqKGrXiq/Rrf
1HwcnBaBb3/eveScawbEV0RZ0RuEU85+ZfmntxGV1Jv60zOKm1pWOx+qC0G1l+jQ
FpmqhSRotdphemUnamk9h+AQmRBQCODBOE74PhmRRceWFUkorAWuh3Ai+Zk9BR9o
wj0kUG4c1s0oltwq1kQ24HEFKvxSx2QZ2jRoI8ER+ri+bhArQRPbFzkYDBACScmW
0wgsJvegUgir1jHf3Mv3wCZy1q/6HR2PWCOLJFgAKXTGXh7cK4G69WdAPKnVQ5tp
8HXeledgtIx89o214FRCUVSgaPkf/iFQh6qzxMNsnmwkQk/HyKhRaNiaBp2AeZtl
yfb4BJ0L8JTMjN+2FTMSa4rtF8yZULtPAUEX7aoU6Lzzhnxrme7yeVb2ykOA+mhX
xca8SJMykCQ6d+Vyx2w8uQLxEZdRByccQuXkdVnvHihqSYhuVVWy+1gNjMJaKyPy
PE2UQhxjt0SB/PI5qzVJcCUTl1BOzfgG2NywpxRAt/rhqkrD39CwSAHiXRw3m1iq
sbErBFCuIRLYef9LK23kWYlUMdDL/03t9dSvx95hYu8Eph8f1FgLHZCD7q3kaDa7
Uz93pmNvcVHeqqQA+XtvrO4tjZJtrRWpM3BtXCi6amqTOBtS267vs67BdKwLqLqp
dZefqz8Wk+h6KSVjv0VrLUY2C+AMmOpAYaiSGke/vN4f6Ylx6sJDpbkkRgbA6hRs
/md85wze3yiFQxY57pqE4NKil67nqLcYk5l+B4N5uxW+pdwJWTtaNGGOuzcV+RzA
hmAUcFDRI9QTMlWCpsyUxLOx1u84gVljPAHVuHPMsZBnE8UNXuLgouPNMAy187s3
C+4AHtw2QvbXGEKrpG0vDS0YZp1NFtn4t79YfwdwBZoJN5HBo6QiUc4xggAt0+Vz
IVKTY0kv/nKXmqvbIeJkRFajHlBGgw45+UdS9Nn3ZvEGt6szQoZcoEmdBtnQ508c
l0MrS6Sf3JjNt0ELpDejgUSxx32UwoAokh+10JOvHjzJydFEfYjdkQ7ljDsUb8ul
rftP6nsgKFNnlqoBygBDbEKYtKxOqaWrrqa9+xq26gSajGeHtVQ5sIQVqBG0IaMa
dKcOma1YY7Urg036PXxF24jo6hjTOzAeDrkkV7tnod516i+c+QY1sept6UkAhS6/
1Rgcxen6v3EK9Z9tCnXigd/sJ4WswLRpiW/z9esq2ivqE9XwLGHc/94MlegmxTHi
u951zbv90nHvBTiwq03We/WlvBv8jzaT4slLcObCP0ZLM5Ep7RSqI11qcJM8RSa5
D+Kf19WoNismtCNmhbBZMZINjMCc/iBdGItr8R+Mz31K9sftWykUPXdTMBMtUxqN
61e3pl7VSRW/qSt9RGu6khILaGr9KyTyWewZjbbw6OznOn4NFO/I7qhw/R4Uxqw6
MMzDTrL1waL9slhoo5UADnp/2ZpsOjdxRz9KKpijKrCT4OVEzn8dorBQPpgimswx
4hpV14P1Qr9q5SQNGuFHE7GoeZSDGWLLvRVniwJuU05urQ8najuXpmW3NaIuoFTY
cGIz/ddzoAk8re6idd6GYQrwOjZyL9j4bLWBDDQmbGI0+kHiwm0vZ8vVfM7EsJtT
489cnR1xZNBhCftbBJrlH54TZcwEyEcBG7s4Jfl9x6cXqYwL80GL07JdQPjnJnx5
lYItoDCWQh7W/p6k6Ym402ONld3B3I2pXrpN9XHNbVKNz8tUztr2H6WGuFC88Pgs
qh/PvFOqQZ30hLhgvhr6Sm7orXlbO8s7ZljQziuTtRvR3y3B01OlotJ1AVRFN4cr
OYQwFhzSMeadbIRrsIiKXYJUroQG01efJZCoMIb1lrfWIx7KQtmWepSVpczsbxSc
gEgyOt4ncPvvCXidXD4dExo3cxZKfeWq/2J2YFBJH5GKCRGHryFgFpnC+zBB2FgS
DbYdnAN9jYqIKQDkozL7YLQMKT4Sz6Q46CCPL+Fmx10NFcakgBebdxQptd7X2A6D
OLGSAF4ywotUAdLY9s2YHntnjzpML/6JwH7vnh9s36y+9lOOmafIpZLrpHxzwd/R
9aJu0NG0HbXCKRX3Sb45y1PKkJ9L7uHlk0MMx2tdfkeaj5WoxefiOOaty86NYmEw
S3uwIy96ZZ7ElP6kGgzYHTk6rGrh5k8C700OyKcX12+uuDFnvV3zp1HVSR+fbjnp
2JV/jiNgImd0bcXndzW3utzbEbekX0YSZ1Zv383P5Dvxm6OvrRR9aOTuZGhyab/q
6yuYuE51AKS4SuVZpM2m6IswzH8O24aC52ZwhNfbv0j+XX5DHmkbOccpBgNb8os4
Hc+Me0c0BI1nNL/QiovIxlq2jHRWC4B34JBZaX7LP88L1z2FtHoNfbVrsTV3Ekq8
EKf8wL2bjQh56KQAvuZWuM3Rn+CMygo2B0/firFBewsyALzgqk9fQIs6Cm5dLy7H
Do31lTf7M3RJkcro3Y5p6JRfxyai8qWGw4FEzt32N/CkHIIm7h8GcMt0Z983pvUj
3x/ErDCRdBrhznB5vRheVhs8RiNrHZ7UiJ/VmYnXki9+vpFWtmJFqC6HukETtMlD
DFjt5siSdh4XKQSzF4vz09XvQWD2D44JThUm1szb1kgCAIEifelnbsl88okoodDk
rprHnyPZBQMOBPvJ/hlKVJVA7GoEZWyCDHrv+7s+yrzKQooQ4I5FrWebyXgj8bc6
l1u+UNjYNZYtyF9FThC5DJv1nsiRZHsQaEIpK5m98J4f6XPs5dZsbpxR4spSN0DA
rYpyRYVFVTnA1OKiS5OHNrBQd+OwigVIpRvNc9L5vm9z0RrlRjwe/PFQyfolS65R
fpH7fxoN8K3J0UmeaRryXVlamxWvVqniA/P3gqx1LPBk8vhQJgUhS4Q+swaNB64W
9JI/CUl1nq3IVD5NSnW7Bkz1bA/SO9OdD/TaHCkm/F4SaJLL/PaafpF28qsN1/le
GHLuCIE1sfNtIn/LHPJMm1Jt9k4nBUTTW97rqp4PQS9iJ7kgQ2RSsAttkL+h/uFE
gQAa/dPOKUwfCh1GNYS04rlUvzQRdPHRagBwLSBHsjOefSvEk5vIiDwfk6BxsE40
A2bNWZvEXOEfKnGcQ7ZR87mSJEJgom/m8W6r1DD6Lh05QfYkuscaLcL3ElG0T7qe
H8l6X0U2BdafV026Qaq2nsJIjbET/RabFFfDl1L+3e7HHHLb1V8v4qcWIxF9rJiL
/2ueibhJ0wS81GT+NoCVMY1xAqiuSMlKBQui8txs1mEdp8hV8e3BAe17Ops9bMPX
RlYsXWSA9mRy5BFltwsby6F4nPIl3bVtC7IoQQLs0E617cEC8olMnZCIfXHdgmWa
9XBkaXvfKFQC4GlHIxWhXKL1lMAwd7wvWY5VnIi8gU2GqoivGtvtMD2q36uwldnq
F2tOEK4j8Tdxf/awpqKXp+9t6qHmBiprHEAt95lNlIcvvy9cXsxoVi0HT7zehPvn
Sw1J5UYccdkgkybUn5o4ui0ZPERdxDPeF6vt8M71HeWavIz/Ylfjx3pHySt8dfKO
q0lI6WsN4qZgDDhF8f8s8cxlXk4b5Fu25xS8DbdTF3JX++XF3b5PGshO74PfYP0T
7EAbzynF1PI3mAWNDD4p1dq1u9272gRP9PrQiwwxRmFYMAtW4zxJQ0blV0bw2TPP
Br/Yntv60BcLiPBQasEzgWWP/hzq/toAUrqfhOWOFl4wr+DVkdQvQ7h/rZo9LCBP
ZO3IjWuwqW4bCgbZEF3KLuLdrSqzaWYXmEEPc7kFJdKa1mLbQ6qwOv/5a3jx7DbF
5unPUDeUFSgUqAsgfgdO2kCh28KVqCOMCUsrm4+A3RA9wulsCqz8OAkGXtGBmXmc
itEGXNGu/NWm6iGLlVTgm6z9/qZw7Zz7wLKWri/XqnKs7mIhXJgC3ZI2Myj7ci/6
Oh3wwN5+23Ppc8DiBy+7HwEla4ZitjPdYiWeW8dh06PS9rUWW0X4jelH4yR1YOHy
qPtumlI4/pSmvUPS7susRa7P2cOkvhHG9yr1XZk2Pun/m5IO3V15+H9c+JeCzL0y
CG/ltye+nOrWoOE2GdK1V81FPepwk14PVxJioXgUoarRJGalwdVVTQ+z1aV/IOCs
O2UR/SISa0r1/KHFcJzP6J6lOJ7sLdLxfKypI4Q42EtLkJ7dKXz3w4GT8IPnlewl
2+C4V8EvQ6hSZQUXf8mXZq0mxFOr5bs/+64K3z+EzzUVSScBLqHYNFyNtw0yGiNM
Uaq5cW7UtdtHUoyIuHhzdWGZn1kWEZFTvV15PwObFHTKGyroHixl0ZzLoWTCQJr0
xgP7OTRYnYti9hz8SrUSFVOWZ50mNtkzIvUMoHg5b5WrzzRP5OS4rC9BCqXRpTgC
DH4q5m+tWyH+zepvfP+LbwG4mob9J5fNbpoDopMljtdEdwzmvOMWBkqpUyk5+W0o
BmxqwndVv15cZ+j+6QArajGbSll8KFRWxnCyrEd6M3XAhatNc2DRyqfPLPc0KyIX
phmkOdAqe3ejzpcjxr+hhSikYSxk+d0M4B0rcg2x9DoBGHjFwx4MdIIheE2FKkz0
MN0dniCGI5LbGItYUMrxvW+e+eTj04eLCFcb93dwg6Xve7d1mXKzEBC+zpvmJvpu
PuYsNyCCEklR+UwZlcVX0QWXxg5H459XvXcyZmaduv1x6LDwmxRbH5LiR7PZEkx4
uXfe15MpGt4kD56Gs8KlsiRorG8WdYv+HkOirbFDyt3I2Z+iY7eqBwtArGyVjwKI
b33uLlc9jV2TmP+Ndd0eNsY3DCGfJ3bvcfQYKmnZ/4AzLNB2iqhCIPQ/tn7SMqvc
6RjCfXP+2lzEn9MZdggGMixKUA9Ksal/WSt8eQcv/k4qmLVMkWUSibOrUwivJm2d
lKHPk61crf2r8NUF1fBlhMQn0Zm04OnfwU77/nMVRkxxjAfzZ/DxpQz5WY4612RY
oKnHqGVCWHxpJxNU+cXbEYxU46X2ebL3IXoJTF+m+5Jzh83o6sZE771OmLFwSRem
c4LA/nBF40QSi/8maXk57mfGJUDbCBg/5WN8wABYrZFQdvB9GaqvBgFYn/UbzyL1
naYpWKUVCN/dP7b1NZ1sN3j8SM2dqdTF/EJ+HKO4BmTfaop16pOsvIvO+mLwPXl0
7AttKQnfts0TTVm+Uf4Ef82PM2lXL6Opkwsv5XQJlchNv8ylQqP4waYQbOthIjG3
wWhIznoiBCjIPxyNMGRprzQC/P7x8EHKyKDhFRu+aUs/4RPWxDu9rLOjf1UKfX70
/J8lzb+6ywc8mawWGTX3BVXRZaf9Pw1MUJA5OODd+dojiI6d0sO/w8A8ivgpIjTZ
IO/jtG3MGGG+yhdbv1mZBiTWsv7cJP3u2qMmvUdzQAfPrPdMq6qzmrXHQVwR8/zS
si9uYwTdBjOtNNoEiHeLWUgriifO/uNaZBdYHtSJoorZoDR6GJe5w/f4XBuCmn9j
yYK1D3C+6ngz7GmItPfA8pLp8Pry9EPfxCt3cErxgTd/wvB46JTEeTTH332vn+8l
GO14LpTAd/UbQ//BrPqeNAtRp+hTGHUArlK0GZzE3WC4p0j8ovkBQmmJ6wdC1sMF
n6RV8v9TMalud3wdRRpyIfKqy5ReRjRDz6PDDaG6/mov5FKEKC+/VrRX/Mq8ApAE
Blw94txLipDg4uiZ1kQtf1zIDBJnEqRnIP4v3abFHaWq8K7yHSvSLB+t8vDsCKPT
fbT2p5tDUP4OG/7Elv9ILojSmnFbqDz6dxsHtAhzlYiv+++F1jwhZHac9aJ3cRxm
UIpvE3BNIcEtXTFIICoofrFx/I0UU3QkYms1kFJ5IKq0h5Gm7XIzXYzxE8c5GXa7
eEsNyZE7RdJbU5Ndguxsqv6YbDC0qALQPgak6VwkgI8izHTEo4UIZIV/ULJCTdZ0
XLDc/Z52UxsF8rnQOKB7Rq5OUpXz5mIWVccPVxgyYm9fQKMTxFWXehNdnomdiU5o
YKK17QFAHyCz98wPsv46DOIQ01UBLC+2VMBxsuw8Bnvvm97JY3ISdR46Pd2MCZeL
/96IpBsLBIWnrLHGDE128qIEXj/g0hs1IuWJbU6xtN//1GAkfk+vaPYqNMrDjylH
2PUuOkRXBh0UshHIyNV74rV4HkpeqoermXGLlCD0AVL5VhiDKbKGotJOoHtFt/om
dyqYJBe2s0poITcVSddGIh4B3gAxpby9vMUXjCDYhUxO3nT92xSmws3lim9uc6as
yqgQ1t4bmcTc2Ib1mv9bIAS951Uwq+cCPBbW403x1lnksCOvEEDLYg0xBZkaE4+T
Caqi5SMzrXQ7QYhhxM+8HrWd2PSul18tJeq/pe4Uc3IrZhwAaw5O8csUcpasCsGw
s7yeYEmN4fN7z6o3S1JUCcJeSVzhUkdkvpffZpbH3rOjUFRzNuyRBGe84UxsRlaW
t7j2ipBVR/cNKy3IHeGOZpvkAF5T8mirkVy3Xft1woJBYpJYaEGnNHx7a5v8YBS6
gnKvZszCTIUbd+5xbvANnm58foNCPl2jjphyaPD5ywQ0iHcF3K/DMxUHSLM+oE0g
gxE6qrWA4PdXquFlCyDYz3L3yR6xwQi75TbNz7cxZWaB6Y88SpWs9kChLWIpqbLR
SizY5zmSBCdbY1cEbnoW1hsfKIAb9UCQ9Yy/3VyY4yDGAuY3CZcsJNmQCO2celYP
uBWmWluR4qQGLw4ilUtuzhhtwDFnrBn+WcnIGnwvIp6CjUue6fzrd6jdfYbri83R
0E52nLEgq7Di7404li/pUXXZNIaAO/E+PLF3yRJLk3Mk08L/YH15c6jk4F8dCH92
JqjtLmWoesBigu2+IL3fC8MQH7aLkrH6XT+vPCKvHuZHiMkdA9LbD3z5GWo6/tUz
LyidMm0VJ+b/RnbucpCIPv4HFbHcgL9/6RLaAzKcqI9imPN6rsB/B6+UbhtxL+g4
lduIvsMXoG2tYDSikBFHkidjkt05QK+5vkRJErJj8mUutzuJOFCQ8ZA45je3jVSm
3iRGJ/fs4X4sQuMVOYqcHLfWXYj3e/N3P7nKsO1uITx1eH4s8UtMKoyuJwRZMk1X
rW640joNqbjZOZojeNOrr6pC/ojxYolPgJl7yljiXGyjetrJHqlRWSN1TQmYhUXZ
qK5OOYGOJ13OEtZM1+tRGDm2bwYvk6m73luifn1iPUYeOrGGSNnec5KiVeEu14YK
8GapiNj2T1CzC4mOjl47TZRBk543K0hlaLMD7O3zOzMuEUEAoP+agvSTBYlyUAem
q6cywf8qLGivbci2cGl8Qxl1idtSwVv409fDOetVwCV8V5oQA4TcGZqPKqvkJPIc
PVpPkjjXbW/6WgRA1ItHZjGeqCTn0BmxpzQk5VR6kNCkiXE9+99y+pxRrZDcFqfz
fbMlpKYjG7GIGvgwSuwXswb90RJn6Ebi+AqQnZCk2t8jy9a2NbD7JhvwWuM3pBdV
zO1yzUcsyvusHCsdRfy4+/r5LBti0UVndzj3R8h9tgekt24p0ECBjERIndcITNV1
gWHqNfVLy+4in12Vf1Ywig08XTRTNT3t/FlvqHLFa2efdTLC1KdlAmQ4VmaJLKW3
/mrHHNyp1El0BeGFux/Bnh1oVXv+xCPf2iUkfUxhc2t62ijHlvC9BJoWoTWlz0W5
h+PVSeRKkYC/CGXPVJhe6+AIO1ybzg7X2RlFZxmpf1hvcutNbimK3uwkvyt7EaKl
BzO+OgDKJBwKQs/IbmRiDYs5Aq0aCMFzlcVXPu/yi4Cgoo/vcsRyIeSZRnfWlM5Q
7xM55fLE5BpDU0CyPH5cnRvQuCTO4bOPw3iaoLjSH5QhS3AXtns+vKX14I8tXlwt
ZI1+ANGJhf31/qCB2wtcZhTRtB2DRfPhbU9JsQwcgPaHlJtxF7rOp/tTQrQFxPu8
b9Sm0jaGw1UiaC4NlS+y98FnVZQFeVFjGmBiLzP+PlVBXhxkcYW0sbPsQDU0x4cO
8yim8ZJDTEaEQFPXU6TQLC37qSv2+pgPOMyVzm+m26lgdmQSoUMoctc9LM3G9mcN
p+1IIEBbtmeAwpUBYZxwyEDclcP4CNM5p9zbjfGraexXJbA+ru15wOgF/cEhDn8W
WwN9EjIsianOl5A5qGqJ6/KPp8GW4Htcx/Hz4jP9BHgB0ryF2LrNwh3ga+VYnLh9
s9YxNvF4bu0E5h5cpeICbjgxrzJKAa1sCmfp6ZBDz7zaS+ly7yDJJbn1hZERoKnE
yhD1YMs9ipwlSB4PkdyPCpZ5mfnN6L4lPDTNcEcCw9cqiTfCCaqbZtiy0R53PX+9
3AZ+PxuKx1r83HMco2A9FzDHu2tVwCamL+TLU8SSmIQYTOg8jK/XbhCp0Z6blkMq
/JNSryd+ESjndbaL5vO4lcDzJqJoAhYuNYPVEeX/yI5uc8PYkvjx9PcCZ9rHrE1R
1dfjiiQs6PagfyV3SqGpCeEHDsObkg9CzV+8M3OMHtd+AQPWgBYp0NrI9/IWpuFl
R2jwhnwQ7LOnsa1DGOyKxw2cGxFu56e01lwxkgoyqDzjC1xzpgzaocacGzl0TuYr
d8DMTWpAD5pt4a5rUQBpKv47nqkbYb8H5pCP9RGGRc5REHoPUrzEwYigpCgr6YiL
6dDaIY0cmZ/pxPl5hWJYLIoE23I73ot8eUreu+DIafHOG80i719x2j5LymtZQ0Qt
/FcNriL0hUBbwrilrFsWse1XCUQ8428jKzvypfs2YaGugB6HrJ7CleW8zmRfbuVi
k1gbtuACqKyZm+bfM9190sb93JG9HMqkKs8mLfN180wmVy+lq9Llpob3BBZj9+SO
LyW7qEFQ8Wps0I/ODfW0ienIydU2NnvQ9nloyb0ks0LFPhbidOjK5Wezg2nu3AoX
DFs0uT6Jz75lC3Ak5LnzmhW51PmTdjfiMMVFccZPal/TE8Hum2xjSTA16wrHj1z0
9mqPhLSnCmDlRgWSrWkliEZhcs9ZjUqZVBNI0Y8ZtzqPe5jE35uvLEo3ULbzPv/X
fKHjhQnwO5KZxxMTdeH7yWVmvNvLe2bRpuw8vmaPs+EEOqNavKbM6BzLZ4VQmM9x
oI/F6+SkuvAH8zryjKZCKkQ3z7Qa5uWt+3mxnvKwOr+p9hjVyxc2YcNfKCs6PIb0
JrzaRkF0U8HwlxajjnmlE4L9b2U45nx116Gkc/thfcAAT+6N/8P/Nm2aHa1fQwwx
9ye1U3TskT1s2PWlzaACC2bJkQO3A6rS7MVWDtupNm8HJdzI9mCfV0O0xSIYBfRj
OBGHxjf7q8SIv2CPL8Pwx9TxlTIpzi3XQ5dvtBuBOt+gH4eJJDhO7zOrofTw1u3d
qbkfcYWaXjTNwCsHI63Gs+ooKlHi8JrCBSNzncxNw+FFyuNaaWg0XVJbalu2lbRc
zb71n7rvKPZUHB3WbehzivHgsxuXTDXCe0Yalt6uamO44xWUT3Rz6dEUcG67ur7B
gtLIfk2UZScXfMqUyrbBr2xznH+ceugdB6pHz1nDljMFHUxnzYA49Xuu0KN+gBUV
CL9ElNrXEnTcOdLsEsvsII62H8ZYIfKXOlyt6YRzDl0opmngyLwnv9/IjSOzS8+h
bTaVSAg2T9HriQhlEV7elWHtWcddzEfxn0fDGCICStqJGZXSX2AS04Hlt0DV17s2
aK3CL0WkEkiU4zlAg6pDttPaigF4R4/ig3tX6jmdq5U0QCnLOahEmupIPe86fuMs
gYXhvTQOenZrad/0j6Pht+0oygp8qleuze6EckhacuiTdCVx7cnHo09XEtuYvGO5
q3c6t21dYfla229KPBsEczIM11Xyxl45qT0qkkXgr/8sfAvMlDNEuBXGG1gOJwou
4ngupt/hwXn5ODJo6KASnjK6xC448ZK2mImtpbSQQq3OsqAKnQBqqEXf0yPMtz7C
i20xMm7lUtgD7q5OR+wIrurxjw2Sh+QpyotRWE4WM9QyXLeJidhFepn1RH6LhMBT
8moBpsCZpoG/6gjnjyqTw9dhCncOMtT2maVq/PVF/y7cKhTMys3Fu9lb1wT6XxLD
u9XxCspRhP9e5604PW/metuu6CrW3tFJ+VvQxpsMn0BCcbG5MC77JzAkhuRl9bmp
OT15GdY7H77N3lszMn09lGspOgLeFgBTq6Fz5WA8XoLjgKul5TITX4JWjFb1r46e
51+yiq3e+cTjn3oMgyWd7bQ8pZRtoldAf4f1fCgmQMnIB9wAJ54SA2ICL8VVODgb
QT3b/jhyvLRne+Ro5pDb08I0AHBrTA1836Q1AmxOXvabFmIcas8cX3T9xeOUUe8H
NB90QimNulQCa9GI55Hi4KICYNAkFEqwxEKwQtK+wUGYZrEX1Waoz7WAkW8jKgPV
uxeFeiQdesICUwhy1fvEPIRle1UMV7wSeQhnJZAAHQ4EqRkIKD+LAaIEsAOpd8uT
vDL/3Vi+DzqLjrRt5mpFwue5foolvnFtaipRjGsQjOMu2cUmWhl3hhEfoybtdMU8
jAyA0q2u7Ftu3As3ggB/izkAhUbsaoCQb9MV6qHYljPYMPgVRjKbcP3vANBo1teZ
zyLl+xiRjyHu0se4GKQLbT0ALqtt2MbAcebvh2Bo8kJYADaUB9p6gPdq/pq+eXpK
bxc8EpWm2oW1thsj093PfXSX8ONOaF2OGUG3Nz2FUVwD1T70yoq/dl4XsR0Yu74h
uKGWDltEsGB6owHy7ygOkjvpRhZOdCOMLf1L10EMCo+C8fjYNHfTHVQfBj4sVZbJ
+9RZcFfYp+3w6IObJmc9vBt1PL2bWsnNz+cp2lp8NdCFc1rm6JfWBYBvjrsyF6rv
IgygflVxlKTT8TLKWSQnVehLhetTI80Vrtm4sEatB+68X3mA2f3iKtYjfKQ/aIex
SPuvAitKKRXZGNya0vhgmJavse5XlYW5wVGtfGlNC+YIQWXnE4UFX6lLuSaEBUwC
EyAakVT+Ntd2p3GpHhPcZuOWRpZnbqWo6nDLD5ygTDLP5uy8mdcsdRQC6aU3ST/N
OEPvXhfPKso0q3BhUufcGCT4KwnVJosyQ37Qi2uyUmK+BvOt5UMygio7bPD3vjd9
n5yzWPezW6bq2ScW00n8lxa5F6TcgPR4ZZ1v0G/h+KYWjlcSaOLnuyXD01zkm6Yt
0Q3mAiODOtLnYqOFJ/Q+8TmOsT5GHADxgish6tDJLgEEa5zlRAya8xeqyyoZEdNJ
lGWGt5vcMWy1RXbHItZMin88wFq9Wz8uwPh1I6L6oWC158SNg2LUjgMYRcvusyYL
/kYCqrUp+vvavLEwmbrgftjkiVNCFtcVDL04PUIfzPNIIsIIPk9pp1KHsisSrjUL
xAyv0jCpaSubqHsqWQ5SqgNj4X4h3spuny+SNCDWP4cAuIEgKVp+BIWk5KmFj+vt
7WuC6jpReqIG68adVePjAxl86HfUA2Vw4gCx/UpC8aFScyshaSo5383qWxjnJ+vO
eIXqF6K/0oKS6SYuazgNYMoxyezeVQLBdBislqwoxBO4j03rP0Aw9IeBO1OOY1Zi
TFfiyNyYCJmjZWTd8QvTvVizChow8m9XAU6VTtrnAe4ew8YNApM8ybpRWhiotnW2
zEEsfZliqHzDjI3mwM13MLu0tiHUDB4T/wixiSf3FXHde9PqswlcGf/P/kkSu0a1
usow5LcANIYtVsxuM15NedLITComKdiwfRbM4tJ/u1Wk7o7Jkfb+aFi92hbLmK6/
RLHRvEhnj7Gka/34zpFCB9aZjpeU4G5TfaNM+vUtax5El0iwfH/p7Ch21B6KLQa5
yExFz04TONwWzq7/0ZWcVtgLtDtzSZSboN6yXhcLGx3FnRDtSLVlNUoWawkc7uET
z3HnVUAScKwUwuXLrGhjJMxisS0WReKcL2MMw54yfJkzuk11enCoHRplZLwFD4f3
O0J6slEptKLaGkFwu45BCVYe7WkI5AXsC2nvxrBt4ufjz5jidhAKG81LQthrJGVK
3rFIr0oE7SDyYIAP32ym/KfNwKj3wBU3QoFVS0ub8ZOcDdI6tGR9snn8WxeXfypF
erCfLgIw3MMv3puP2npPHFj4wUnbJayhxnkjBu2Ma6HcgVbOAXCno/I+HFWHZ5tI
lYzfcae6c6gWvr6c6zbiIfu3jMutl+WWsQfJ3BCbntobTz2NbW9ZezDuaRh816qd
RUU6aroktIw8VV0L4Fhcobx70TCU/OCG+I3BtH8k5Zmc6Fdw4d2h2jqVP8aZ+QqX
GxiiImsVdRliu00uPdApVFwqu5Y3fdkmmhHLUwHkYQv27krrGqXuGT+UpRy5dPL6
rgb5J0ZPIjnN4xc6XQHDEYN1GvyuK6aXHG0z7vwRGYYoaanj2E2yUncLEzta6SAJ
oOl52DNeuSZUUsb5Tg2XHKyYKSrWgoZy5zVtn6qMIYW15w6CoZsc6zJ3GsKpHoj2
m8mJIosILcOBG/a45dQ4yg6cSlt6kb6DCP95LgSiGF6IeLjfEU+TDL1+HpRjl7K8
YqZggHF5HOer9YnZu0N5UQSkmgjgwsFMNQALq6jlYtgTBYYN0gwkTDbK/pFs8tkR
eJURjvFQFvkZK+VXoM/qXZZDBeQ7zwgfQprIFV5BmR+9FKozZdFZf9C5ROg9ACSa
iqoo6oUDtkaHiEe31rNWNwPJNWjYy8a1NMTS+FSSaJe2oOZ+789+nhSKqKtz/Yk+
1r7eJGq1I2NLHvt+NvVLISyC+57FIC32X/Nx+67Iy7XdA9BVDfOKc7qvvsfPhm77
gjzVWp17DL//29S5gi4+y/jUNZXcec2zmfyga/MpvlIIXiHUqAwR8osPJxqc/UqF
cYsx4FWtaaX6IojE51+oxinprZCQU6lNAGKbOigKxo3q9ruqIeQbTWc46wtOPlq3
mKqYzKnWlWl1cXE5kTS/iP8Ae/jiFuTDMIv3cHZTeigmors+uHkSmYorcpiRHDWd
mfcSOm+aWTXrwSqoqF2BX/YeTFB2NktPpJ4fOwpR5AItu5gMu2+ZknYsb90RWRB5
KqoIr316JaAJ22BrgbC16RCoviSPn7y80Pvv+v6N59n9xWWBfNY/YcUSEZY3esIa
TTv78LXbf5kLnt+TvaRnKTntkQjY4uyGKi7lKZ3uly9ieVlMI8xw3b2oG39boJev
KrIGTP9SgNkAxJuWsoPfmXajH7W06Jkpf6j0sY78as14y/3Cp2ujArq89A+KTlTi
YlTeqNAcfz6Be61e9Er7zYctaabOsT5Ck2QYH9CQVLWD2+Ig+/cUS3lfdQsutuh5
XxzNwKg6OtsaX/4InMDYbyJbJwW65EzeZgdDt/FVeC6ZNieM3EPOLBTC3gV03fP0
5J09Uj9RcTbG/HinhL2Y90nG6FMPWErum86iM9C9AZgXS9tcB7Q17mE2Fv4kClYp
dX67bxMF1N/MwRvuu/cnaJV63+NTgFWFZMo7wG3ND20C1tvkFyHV02n7PzTikq9/
pwHblghIIGn4GKIiFs+XsvFj6GyzzgwMa/O5PkCko6GbGBML52tYOzcdvMFVqbDM
bONyd/m7R5P1E4SQUehyzpWmswyG6GjEvln+9uD6wH52AuCXOBQ4ltZcbHVJxggw
HUgL6KPuS26XIZma6Aci23mwQ+FuKWjCYVgyPtWV8VyDyA3rfe3xEMx7GsznEikn
bovkb3I5gST1WDYVNkKJZwRMAs3B3M/UyDTdnJJj758drkX5mrB4o30uNSSEmp2U
leneyrQbgkgnxMpbiRtefRNvlQaD0ouOBSkgEYJWLniDQasaX3ntYyJ9sqDgjNdO
GBZ9jJiNwQ1s8+Dmy4Xd8C9yAFu2zKt5WYCjrzVdkKaNq3asa9sTODIzG1vAZkSd
KFBcXdIAGEqW0zAE9V7tGwvOzjN2C7t6+aNG8Bflec3HVVAY0AC9LGBri9Hehlam
SUi17F5slZeb9F2nGmaTBR/HTI08WZ4jWztgnt+sfXo0APZb3ecLYnZ0ATleX7qN
sdME8RmgBU1whrLfWbSW2NB5n8QB+tdBDsR6Qve3exXrdHzTC5346bY2gwIZFW+8
msBVVHL9PchWEqR3O1rJA4wXFQQq6h0sunGCsr6W+vP1hYoDYgGbCeGhRs9zd7OQ
2QA+oU+xYyengVsewCSsxeNuweqb62GxpSNiYPA7chzFC9XNHdT7ru9cXGW0H34E
WaIXw9aXNeyA2tZPSu7fhnKueRQ0ZWzd0/gtXoCWz7fDdAvXxwsEKzaQKPFdihtB
n0dhvBohQk8mFHRjfqDdvHWHn460hQ2GsB5lGVrLBT4f11IfSlxWX96/N6u/ci4s
huPKQ27/jgMhFbbl3UjElZmsVepRIAwEtudm11j+GkczSVx1+A+yVh7F89lta3jg
V/cDN9p6QRH6d+BsNNNIX6X3XYP9P+hkNhVJ7Y6QXAo+SIjdFz1lP3nTLJJlaZZs
d4/TOp71kl7XhgZG9VD0desu9l+1EJXRKpMlHt5lG8D1LjtOIj2k3dPWrJlZ7eqb
Z9BWe0QjH0se6fNcEGYDp618VIfYJLDIlrS/0l+XxMLpeKrpQw0bfeL0yay0P6Rc
7bZc/Jh85n7/TCb00ss4j/e1Esur6U1brS5qsGImzWSxzr7e4IuYy0y1zRFrwb6P
3QOyFzMlD9yRNGX15YITjkH5I+D/d28khoDzMl7yuf3fZgqaeMtTUl/88Wh/bW/D
BaXtm6cwmQHpi849VyS8riv5wr+9by8N/l0r0M3usy5NgRqdyaHHzVLndibxGrYM
RTtb1H3M7aqbeIgaN5hrPkjbwhO55v4GD6i2MR9Gg4YwvrJYpfi5S9+Lzrd6/9KB
XLcXbSTlAd5WmenKC/NwEyriPLX2NFlgb/NwqW/mUh61Uck45rSfwVUka8rV6pVQ
YyhqKnA3b+EZggSHQsV2kM2bP8Et+uL9uT71l9WjNENcRSOIJJ28bH6ymTv0y9ZB
ljl/WOxopCiF7wEmsXxtQgnWawuQ6RzUAZvA65k8D0zF0hgsWaPzTHSVJAwsBeuQ
r2z/FTe4gIQLWvm1ahAZHjXyYyYVXhsJX1Z9QhYyz1mY8gtTzM9CaFfGD2IkXnia
aDKt5YZH1PMqx6kPmodA5pk9jnnoeCBpRTfnuFIku1LxLLoEyaJeIIDyGozkgPMx
TtvtA7sOJKDjDHVG6G5WdqvqKVwkif0GZ30Q2zMf8gKbCnIA44GurGE4brTMeJhy
CNzRB7PiOX2Yqc/whUYy7Jssrt2EV+3j23IL2WbcS4Nwyk/AKAPir8Snr8coMt8d
Ks5D8BwJPe0sodjBwSqhQ/y70e4o0LfCnN6CY7fRKSCYm6uUPbnB5FudaKoCmVAC
g+INyP3FZiHSmXyZGvMPrS3xh0vIfKjeOdUT0Cqpti6ke4PQZAUTw0VXVFjfCJKB
xhdR9oWshN/PUWv2cqKHZD40GSuNZD0juY07OmNxirPYAnKnZ6Bw/VNBubQWaGlo
u7Cqdk5kbf4eZ7S4eX3BkyogcLRJSuPmoiPB667u2P4IFN9Ba3Vn7W3yDIaC6Spc
LDO61g5dHV1CN6OTedEzdw10ZodOfXrTR7YQEc3HBm3XSV1aFHXaech6vH3MH+2I
G+njW8ohyM9mKQGzns5s5ajm2LvAk8GOkdVDGJSGbpX4FhFQNjx0ry5ETF1lwk7S
e8QoIKDr6L9GKg8q0o92Zf+N/ECLxayv3fZOeFRve442kDRJfSuse6VuUBqW2rJv
3AxyhWsh7q6MVyCo33tSgeTZA69Emk0hzX7NiVp3QoVQf2EhYOky0HkwCWW1KNKv
kDgqoOKYiI6wZT5rLXVrtU7lNmFwNUnxneZhX9i26c4bBbBKB1A+UwGREpPrwRHe
Kbe7dbc/N4jAMmgWBuZ1suQRBl6X9Sj3Oq8+YfugsWtiLjL++/uwXGZGBHK+mOGH
rHcPOz+0ICBewxxOFcQeIZl3UnWvPzt2cyd0ZSISwYH1R1bSi7rMbGxW+zeWfg1u
o5E3Szv3+LB5ozS4R33ocj9Dn9y8E7ktkM7tEmsEUEhvLAvQ0lrJFLiVH+yL0yau
zGZ8OUO3FG7e1gjqm6CecPPLsdk3pubXbw/OSdI5ZdQrMYcsmNrjiVg0E9SFJ/qW
vvntssTDevkTLWhzSAzlT0tdx8rzzos72IOMR8Kq3iKRziZabJhDJJvYKP3BlSrz
s31b7lnz3I61A9jNiwRI4tOgg+0voE7ccyDFMggYcQ0d3wTez9/RDHQSJiS3zJT5
OtE3M3vrZMfQpZQgUfojlgXo6usSmYxn7o6lwMcKOGk8OGjZlSbGR1jvv7wWJjqt
jOeEnVVKGS9Vt/KrrSpbitRE+jYk8d4vyOcBlw4YS/vfQa9yC9Zry44xGBVmg9cV
BH/b04xnRAIHPwNat/k7Jp5RsPtxmeE41Qxi0gltZxkvqAnKQd3vQsnh2sGv9w+Y
QSCDSJCZ2o2YC0Wl62lp/mcFIAleZc0P/zP6794ueL8YGzGgD6AZ+9TPEUhrEXKL
Ow/3ySVdOTHFVwk9Vw+D1oewjBPg42489OpEnabSbJe+zCun9+EUX/ZqQRdsorpZ
GA6aaoUv/4b19Eyl+JssKQK/lQ+UkEyQF96fwFgsoEDlsN1amhuuB1bJIZDIN0zj
fSRf5Yazs9j6W8rZHfmDCFi289zjkeypSuLT0li/gGNvJ3uEqXEN73X2Kdwhgt2U
q5h/8FsB74d13TD6mXNpqvHja1GmCFfU+LHE8lZCnfN3LkQL0lfhFVNjzSo4KdKQ
MmhJ+pUlz3rqTjelqI7LIqUIf/iUiboNHM5lB1Fx5feo1e04FVNg/1sSpg81giY2
3UVUQvk66oUxiTH9ba0fjbYH8Fa1AcTINAEZ9j9fIMoFHqCLK3eRDjC/2Yq/WDxY
JDdamPSb9Rw1/ezBKjfinfr1jxn69vA3dgld8Q9crIX0rZ/ZTFcBJrpxMnm2oxb3
pYh7pXsLV2r/UIvkY+0qL6gBiTUPuL+i4FIwyOBiHrCWT/8uKYQDMHqHuxleQHgE
kU+AfE7vfYgusre91j9SMpJcQYK/P5Ctjq/wDdf+ArtZAAkSHBCaIrFhBTisQuqQ
lp+rWQV9yYvcvgT10ncmYjtZ8D5lWS/KX6iE6q2cxGtfNxH/ftEPR47+OtTshH51
Vt2eF75+IteY6huFXChncl2kVBz0lvoXu3yYGN9oUDtCvxlBg2DaeF22KEOV5zSR
NwvBeSBpxAyoRypAC8fdxnIidhnZB3AjmokDV9oTyRB6C4rymVJfD+0PW/852SDy
IaZ0WEYLes4btdoDBR27jktj6f62TzgrmnpTUPa5sW4atcamJW2EvLba/9yu9WbR
1xs/+eq3L9bVxMm3BkZVrdY2Oop7SKV0kjv/LSbI8pmVSCh7QlL0oY4UAL2CBTV8
atnPWFY1CK3cdwZ+aLtiVdf5ehtyQhovb9DnU4jVygd3TuFzejBJ9F7bm4gjsGdT
0Lvaf8rrdeBVkybWl26SXG4hcOda8r+X406SvPvh4qWRfxL2YuOiyhesJL/Lanh6
tp3YOzO1Yd6dHr4p8G+utEF8+DHuqOqSb5R0kDb8gO08pwywaUDStIRvoCleF5ir
u/+0HGTS9rjqQWEh2QrUGAL3t+v4u9LRsRZwjv6LkdEJ+vedpRGbuetyw3/m8sP1
A7N0PUK7WO7sabQu/sLQrE9ctgCF5zcUgOzq5Vj69f1co7/30+pz8AOUuuerG5pi
HUKkyS+wckVhhEQCRQ1EplJ6sjcGx6xX5dvNRIbpZwsH8E0b8FyVFFgYafzFYBK2
af4alq9pnqGwwe9XzZrssSeocwdU6xhjBYVe2ZE1Yk9Zn+9GFiXYjJqSPUcyI3EL
f6y5gZTwP0wAs1wckldEhHnIEESq/c5QEYOCns5c0HBZ9WfayKfK1mjg4TL8bOX8
tJUmHWEVoo0phdOknxN4+pjaVPX8JRTlDkiyOEa4greuDz4W//JO/J9DPq2lLTEu
ve4RnhuvZn2J8l8JpEbdzHku0zJmww7olUaVYi7IMKjkGvkvI2Hna8ssWeS+1859
06ybFWpm7+4ewVsQYCdEHC4QLYQgbTXxSzjOU/JkHgLqR6cNu8uSBxxtkdffnV0j
CB3t9iYWyeyxb4IUd2y8wWy3TEQo7F6j3ADQcr3iIVPmlg8hMsiH5M8AD6uub8bh
DA6hBdiawAdRTx0JHmmKj7fsg0oHzoIsiJ6df1/PfrTP/lpnmNJ3yjyRdyBTM5ks
rZ4sJ/sCuGIOtqpzLBuYLoAiRF0xcJ6i0pdGDZDOm2xgDKIIwygt9jSdPHG2+gWD
6nk91t4uW/eEHdlmf49U6zNWBpShaTEsbp9kf8jIIxwmXvE07d7aD5o2/qaheWGi
0vs0rus3WBxVR02JBntaC8b4NeNHnrFVtm7nxPooDtzD+6/zANd59K5GVYttrqZV
XLi7vjQYRP4FtHc0yc39O+Bq/8kF+qwRRTRxFEVVzvcdDUc/Jn7j2XojwIqBNO38
5RgMYkf1GeGPSh3N4iUK9Mwr6ta46nof+YKAtx6o137E687mUu3Gnor5j63HaClS
EtX+fRl+z0pYvymzfF2UISF5pm92ny97yjhoLtIyv3uodMVFVHs1w54ijWu3F1sH
+1jGD0n3YbvhW9Qkd2dQ3MTjEROZRZ23xHGWzSvmQjRJ1RCHJxOkJkUxyPTL4zNK
aJIIq2HDWWNY3vgrjLGEcY7lLOUM33LwVsKoUzZ+jK8OYfG4zGcYQ7u5fauKQ/Ol
qxY1P33nogfB/YCBWl8kVY8VLq299KwfYRYJ1CHp185aP+Rz+cPT+8Qf9InaNj8n
tyHSKtF9Eff/MM02Qh8AaYK01Z9dV8AIbhIDtoQQEG2x4xHzB7LeoSC7qf2aJy1w
2C2wIAGO2bTp+e/TkpSbYnr07gdJCT2G8xvdGAjI6OAok2KGJ4qUFPBTrJczn/AK
EX+FkMkrLE4trtA5WT0TDAx48+UkAj9tXZYSV8COAHZ3UlvJbBJXHnyJhJX+fgLe
WHlOXG9uKJk8A4SO8tF1AvQS7A1Cq+N9KHVj2VTf2aeWLzvL+dWO/W8ZbARz3y0w
R1u3GEfLRLeR5wAacET5t3dYoRu9s0gbVPXfVMYm97j5LVPrID9qT5iUeONaVydP
XAHw85IeUZwupWMDX5qly6kGrQMYd/qMarXqll1D0CSRqXJOcio2Fjgd13QhiO4T
iZ8rm+n9DcwzTBmGi04H8cNX5btNyr+mppdDz4ctEnqW0NlrRaHbQ0snmhT5r68x
cBqOuAHuF9ojAhYhsDFda1MkAEfa8dLfg93ys6KiJOxd9gqDR9t4Foz0uHTmfljD
6O0tnYdMK/RMoph31zPzfxKHfTZgneFuiZ0bklvha3B0OI6bJTcFtgpRfzUxNRJJ
0mpMfR45Xq9sYF1HqPQMVSYy35vJfIYIeUI6NlBbe1eBuLHKZhHnWhL5g1KsqYT3
Hu891tr61H2lfIn5x+XB0ytYKAIc9hQryYO9sFtSdg0a454tanzDfSjh6dHBWihk
1nOTAUeAwBDTxLEmDMHxQbTkXcqznx1xlpqwkhCjXycgvdztQOoHCzElwTo9PPli
6ltv6olFKYYj2iEY6V4qzMoWrOwD94H0lSHPgRLalQeGe3tCjQeMwpipuX9yGOYm
HuCek7Xhf9N2fcJiLtAlcM+P63BtC3k6moTsuv3nyE7xHNZWeYb0hSBmKdl0Tqpt
1y7UG7sgBE6v7oVHS8MEa4mS98b9lPyzTEAxjdJWVXiwJiukAzbK62kc1zB7JH5G
NGXYg1KlS1+POgoL3A+1dxx8JlBmPzthwv1j7V11SgEfp9hjWTYfxLxNVieBex2D
mcNMxOsFFA8JvS5lsV7pJpV+wOlD7+4j+CIu1B0tsiOec9HOsURjjT/HKBxijIpJ
NH6KsII5kLi7iMW2CQ2rlMzk4ox4dwcMVR+gKQTgYhCXCSGHfnVBaUVQqAnXigEs
ySIMkzbCQuxc8vxyAkE/ra+FrV6OWp6XNVztsjIcGEojBsRWUSj/NP/rJYx/9e/V
GY4hJriFQiAve+8Hc3AfAAOj/YeYUA7Jqtlh31y1rE5bpOS+j7K+ga6WWD6Em5eG
GN11tCO4NhpS+kD18erdQy6t4eW+FFEJLRaoSl128NZbxyR9uHeOYPWJgJ4iMdY5
twuBygt5yKuGEC98vRVv98n2tD4adLIVUrMnjCUL4y5mS/q8XPaWCl/aVRHBovMI
6aDZt1Ze0UMrYNGERvONvEi8/h2501LFIjLBRsMnftWIgAoxo0de74iCjD6mvB6L
1K8FHUoQU9XzPunvqHiX6bSVz120BHJrb/XlMYpm0FrxBVmREMYOXx4pBZCEOTUm
vPFhywBh6Orp4dJePwtQh+dLW7HC4Mq4YyayP9oP9v3C7az5sfoQULku3bVoMdUc
SuFwXk8khjFZXgMwjn2r82/H44qhBzlzu67tHf2bMi0Lr/enbtany5hmoW8YLO9G
53FoYPL+hNFd8TiWJjIfU4LPPgGLjYAf4J6FgbKGXw7VUHoXDqNjrcxLro0jUXTy
Mw0yrqKA8qa4GtSQTT98txrc3lhLfL4qO9gy6g+BNokjMgseNrj+ydUciqBjdiy0
+2e8Ikiub4CjQ8yB0fcZ0+T++N4U8e8BgDQmEmKMiFu9MrQGDw4vH5LfW9Ql6CsW
pfapu/SpfXzLz6x4q5Hpfyo5oDjp1tWZ6wOY4fFEdqxVi9cAU0pDJKfaWXsKFDvG
2659zDx8H9VPFThnQfHhByW1/L8P+RkKyx98DApoz69TvrnFVXD3vxJdQDTH1M7g
Myk4z/lBxf6RUgY++F+aFlokh6zoVPo72kWnlPAjjits8S9WX/Nc5iQgRVcysKFr
sl1ZfOGyV1TgN5crlDDXwm2IlbNjLGeznLsr0aZFfR95CPi7GBNe96K7Ncf1G1dU
uy+gKgwMgRhCbJbqhjAM1MtkKwzm3cwFseyDI+mlv+NOPZfLmIzTETB3Jxu+S3m4
RQ3unVq/EHt5+QAqYWiqBLCx7BNnWkZOtWBj6PzQa5uITwRldtNVlTaA9yDbXibg
KdnryIcsny0zg0/SlR/jWRCX6Se8XKLhc25mO9xrxbvCsUjcf2RbQf4Ai4r3ffdr
IKj5lxPf+/9NlgVYGM+ALknhD2sWxn84V7IoC4vtiWpD+70m5o3LVfuiafNvxWBX
d6+QKaiEoEpD+rVXSWwvhqV3XYEDhCAAGXl4K0LbXkgmKEKTLo6CftK/56WQUN4q
1ANT3ks1M4jFC0HZVF1P8XyOVK69ltuSESLpooEV5q87uAbb65ylNssaSlc96CXv
kXyNT7czlnA7BAO2vbeIv70AeUPj1WVN5CyPy5biNtVsRJ4UB5iQ7r1iDMqrooX8
s709qT4kKulYL0yxV/j/tiDGkXfcwnkrtDbFhbW1ad8HS9GeZBY13/5RALRq+9Tx
9yZDbmn5vhmqADqVj0XUuJ30DT+V2tJG6IN0bFQr8b3SlRFW5YvO6k8tFjZ1fNb/
EVH1quLeX1yDjZhowSM9QddiiCoq7wF2CJaMZNuE7Gk7+1fAEVgCRS1pSOK/0slg
QMXeoplrS3UV9R4naVGYchdQjPZbCp/n53bW9E/sU1w8YAyvr1ionV6qNWttatzr
OQXNXrOH7L+2rZFpruMgyNHeQ8TAjOuIHtruiS1mPdtQ70HaLisig0uQl3Zd34kN
17sfPDoIoCOOVr/mpq7VjsNoSd5bIbvFHbnGwhbVjtDqEC2Sb9j77nQCkz7/pVX8
Yt7DSk1d+Fh90hoUKzbVm8lyhNyuubGT6TeG70NXmtVI97AFGOvUKafMONL3hf9w
MrxDcjJYAPRvoKgK2+p9Va77EcSZHNO+eFsCqr2d3ZANrzO6yP6COXfzIaAnAxz9
v6YvE2PcvoYHIiUhiLdyLLDFc6Yr0/03s6lmkc/3BD/OVHANdlwvdfIk17ktTR1a
NAPSh9HwlTgCdtOx0UwsRET6yU0Nlo/vs2vdiFkL9hm8cPpXNfpR/qJ2Wgv8b6kE
3QD1uk/LMT9yU5ej8Gh+PT5Otw9mxHNrC++izoQkmJ9tTeZ3LHR2SCc3gjZROim1
pUKKrEUkO6Dzn+UrrSGn6bClBRhDFiVNhes0fXgmUnzdsJRBAjYL8WzsPaIYZGSG
PTolQmXBxdpgg2yojX45/z57Z8+qZjM3EopN4R7bePAzo6XnplQY/YNWs0I1x4Bx
2+lyuscgtUSg77vBR2Nlxyb7+KkEGNYWmFksMshVc0l8HFTi1SvP0OmLAeHHyoW5
0P0i2PxzOiIfXBxznyH5qpQTYSQe8mamfLF/0SKSO/+QWWh97m+EoOyX8AxBoaNr
7Qw9yVGoEs+EXYvxjC87g5QYCkIn0bZtzsIMUKpY5i0rmpNbJvuIYPifOfLfsNEH
gb6EKzfp1l67ZavdK2BWihatdjvVYTWr2a0iLCmYCpKDcgDeCoFVuenRcVFPSMvr
jQRAwjxOpDi6dFtLCaLJgRkxv3PDq9XETI3vlUTeqGJzEWZtAd7EE20/wOI3TN2L
28JMnZE3iXcC4krzNGFw6NZI9PuscI3dqw9NXHWLDCcGwCcUMQudLPX0oVjbAvvw
rMzffTDkIqunyu+puSLo4pX9Sm60DY16GFryyrt3M2mJPvmptQBYOrKo2sNhze5m
0mANku53k1rwu6nl5NxcJFqDalQ7wG9aesru8dSWA1oDBgnl9PQw9c1sxDkDzIPn
psSVynpa1GBG+nlBVeL4MSFNRf6BOc9oOlpaa8MIDCb1ZpooF/FWiMgHj1cLzabq
+pN93wIfitu0VlB7Wg6D3tV2ScHmnjY8DS3E0+CNotRtIOERaD//3wxf5dCWNmii
H5BJyVuzFEGvs4jwIhhsPsj41CRrhj7PsgqVjds8d3DMpMnM3UCa8eK9qHbLs0Ym
GgxMXFXInf3yeV+NHKQhI4Zk/OzOG5JB79DDUofieMIN9xS+sq4JHPpRltncfiG0
wMEsXjQY+bW3kbSU6mjj6ikHDaANWAGKKaCLTNuELD0DaHFZ7xNWJPE3ssWU9pXM
tfTTW1xWPe1M9TKIJJG5iEDXJuj95n70i+xQlRFZnyXjb7fTrCTBO8rMqWJ4eYkM
AM32ltKitoe/DkcfNlEWZI3BPtE/agxbP2Jbi5MlJYYmEBDspBF57hcT0iUjMAG1
RWjOrRwV8ARMStH78bGtRX+86QY4tc7iClDVveH0xsBaLEYO/jTp9nHgPxUbWqDU
qQeEyCM2/6JcHam5l/h7WeVZG4juWIKrmv4O6PkMWdCmUSxeU6QLJ6HpwlYIqK3B
RV2mg/1DBSYjg24wRWL2aBqk4sQ0AOHJBI96gjsvfxqWXh/hHvLFQUCux0J+Ndm1
4APBBN7mEZFYUCl9PQjhCYphwZgjyOUdIsbFUX/VtEPCn/vH9kTjVFzda708/Tz8
75fuw6CyzTtC+SAHRIfFbbZ3Zdv5hQeIhv3iTZnh0eDhkfHh0KYkaUK44MikEKzr
Z62w85KQK0J5RH2Xkhh3IiE/WmNVF40mrGzTh3DGsYqmp3en8yIrZbUYsJiJ1QIq
sLaoou5sd3uCwv+5iVq9uRYvxH8UmKgbRZFS36YeCpiLLImpSGjjmxsbEhHXLqAL
abo0b8yk1FtVF1WJdZq8r3P45QdtouLSyKtrW2R7GE/SsB+CC/P5mHs7xYzmoH22
agvE35kKSAKCuulgsPRgx6bE+czuOTCv7XPqm08gSLHa3FEahx4VI9CQ5EuVnLYb
dIHH2MteJXkNNVq0SjtmyIW9NNdWWo7Ydt15XTiDPqclfWKS/rBaow/HxX0zo71G
30pOp9XKR21DFf89jXHwUDY5YIfMKuINud3l5MLgyl03E7q2SI9yPS5lf7Fk7lCr
x2Wpp8JL1UpBqKQxplTrp9oP+wjYWeau/ZAwQPtTadjnsPnSFRpTZdcPcldAPm4v
9+jO0OEKkfJ3kTYtMOc7Xzdzc6Vv5meM2Gaf244yurZ5iarndjY3Br9gPOKLRDAA
oeFDZeJCPyKI3LKg3vjW9iQnxtKTfPXlqmVKLZNMgL0L37wHCCTqtRKiy5v5Cp5b
r+e5x+knXmeKuzq1LTexmz1JSotT4+pHmXV7hiW7CBkPfPxSEc/r+TeQ0qtMhTx3
2i7zsJuymjujtagVW7ZALmwXkF/tidFHaGo1j43VbBkzr3l7mXvZcrUVnjyCOUv2
SA9EtpdOt0fOB13/nnZm6lwjw67IV1dSDGVf6+C4PowKijSJyTAIbqvI4ahn4BAz
wizJX+sa88pMnrMrs8+Qjqv9U/QmUjzsOpeTn2CiREJn3Re+rCEAAKnnE9Ls0xWU
QMi2djmng/cOvsjt3VnQKYM6kGNIiqzX9gLLNQlbyTq2SxMhDdpHFctjDvnZbwl9
gErZkv/jT7gHI9lfVS+MAngtr8KuIujj33hKG4Rh9QLhVyuOsCXl0R4JZQ+qIduc
Uz6lv2pb1KVGdb4123IYd4AihJca1nDsX5ipUUsmFyJoyL8tdlMW7I6VUAde8Jht
PMuR2PM51Dv6obNgrqxgWFBvOHOvLDBVD3A3O2arcDaoFGuSKbCrGlTVXbkI2n65
Bqhrzw9BgJj8APeoTBIewAZEIrBDnLwzYf1Rv8HcGtiCrSWmtWTiQ/2kTyPZN5QU
8vQQLzhyGi1w96Sb81iKsoU5MHub494fvQXt95ObiEL8tvBy05h7rXJCHgDG+Jkm
fU+9elJwhktRSTZjiwvQdJBXXbK7k+kmYPFU1TOCsVpflFPCg4C52jj9dtI5150r
bFhK9nRfQnkijejR6MeG3qruvmRob1Mnig+AOQuBYoIUrbeyfeyw2paT51apU3yT
FNyfQVHxbaJLAwxH5zmF0E50Gbab9uyGWlNACxlhAM+mp1ZesZ4zZs/oMkeg3SE1
5ARuslA388se2NWkYrcdSYhFVsVa0uhPIZaRNpy005mlahyzIVaMIALSzILsCsME
bb8p/YtHlggYbDm1L0/lPbVYULwlx+D5u1MYFWBR8ICyBN6a9jz0DpWfjJeAKVbQ
3LpVc8qDZX0rpYWPwR9pzs3oH4FtgFQzTJrjp4+lNocy5f+OvEgYdroOLC0Ay3SV
wSQg9avVcMgtg9aa6Zaj09NGEg1RWU6evNy4qGJW7pQDbYCmVuxWcfwp1BrN/HYV
y3WSBp/3YjARpPijz07bO2d21vc/sKM3ZmCH7KUCkwTnnO4Thn/EEAYXPw2xFhiI
r1truarZ+bVkV/8MCe7s307ck6JD7NeJsuYVd4u6PCyfYKGnakjKDfVIVXyEJN2M
arLpd/q+5+MZlurshAvPB3laL2m1/ZNyqRjfhSnkbCHrQfodxIpxTus0ulQaatih
+LULG4AVYONSQIR6XQ80Ww5p9CDCDIWZUMGcO9Vn40V8So239h2rX6MbX6mUj6MI
nZRY8CdgS4XksGWDP0rwOyWAYt+O2TNS3nUhWFVerGkD4w6qcnaYI31s4YolMf/b
UwzX2FCDuRW5tQEDhPuNPDwsIiqlG9lmzd6LvFYD9L35JXFLeCqmGBimWeNznn+O
cqsbhVDn1eTFtUIQ7SQPtzjmA2cLbD/YYSmYs2zR96PkGS/6HRP5vEeaOiDLNkvr
7E9fCi8STeELfyvITaXEE1hWGSk/c9YTVti8j1ORCF9ThN0uzHdzNLgq97iGpbkE
NjV067axJ9Ocw011ACGk5Ndt9hlY5RkUF0rnemdxjMahJCY3mSwXR1SuSxmz4rNG
jIsJMN7Gbp6PCUDSY99r+ZVOtIul/9YXZOe8nd81Nk8AR7p2i+sLGBxTFNeTkaEI
DTxR7gh8qJFQMZeJygPxcrPJXWs8RrERsXh+1XXuHOWICtwrlgFPgKyu9l2TDwRr
Rq34jSQD+ipatSTvJsnZrCki7MnPH10QnpGoJVBJopwI28U6RnJuF779U+HuN+A8
8urDHn5pvMsySkxEMnEmLa90val9KEsFS5TZxHez+yKfJ8vmOOr8u1m5wQx+bd29
QVw4Q1y7Wose2ZZwsHolE2LxdiNhNtQcMkdrrqbq/CzXBzShMKG2dyqL/HnOF+0y
cHsoiNvGMxvw3ixY00DzKZjzD/lE5Of11U6zPexG8MTuVp9mHA81dZrWN/QmtJib
Ah0OoFq306jZjE2/MsbAOVKohv2wzfbu3bX1dNuU94v+tDdnIvcBGMCmpQpSLZEv
acy6ArY2QT4dltYoo1VzlqacdK85gbrsFewUGDj5OOjJU79ftisrqq1keB/WfpZO
M9QpU08ty5vCeyaO5dNydESY61l2inEwIUXWp4tUtFs3tnI7T4mi00YoVFrvCVjH
xZLCV4s3PamkC9OdMAMQaFAi94G6LnItOSygb7Sus8XifXAklZDhX6WxjJrZ+9RW
86jDAZt+RAWebR9VpVsY2vAOQFd57rS/iv41vFhRW1msdEK84nIeRH+/sa1et6Ws
ii94lFd9uGZQcEn+FFlJ/9RSbH2bZN7b7hx+f5FTpHrhHG0XL4PQCtvm3KZ7m9H0
oEU6MjVp2cjtp7abg1vxPazNBdi+kn9l1lKf9MYwzEVUxcN1dod7XBL3FVAK4JOe
RwKLc85usuY6sI3W5Gb2qdEY2RYLg3XPpZNPe5Va/ZQb2uMz/z/BVUI35KcZ0DWm
PPS6VeEUV4iN5Jjh0Apb5rpdSpfgvFW3+9i+/n49WvulhUPRJODCD0V8eeSUl7pq
6nfNFiQbnm+i1STuf5t8JgQF7XfhrrteoXoPmKN79kAmVDuRb3X6WZ04gTLSgK0v
4SbKUpUdyYALHMLgg9JYGSt7MFuWXojF9AIswaHyEOk+zxjTTbFMNCujaXgt1TNV
7RT79ocjsFO4RA8o4Kel4U/+YgBacCUmklg7TU5NRERnqqgzODQvS6bDTKt1nD7k
jaxK+Wq23rDh0IS067oysfDzR5weKfy7+Rv+PXGVhVLlOkiJtR9gf5YTMdYqAqdj
rX9qpjPh8NzkVU3QoD81QvkeWA+uYywb8U0HFmpN87gMwEIQKfg9CbDyjmcH5mZd
+/QlRHhJ+FVXGISMbFqI0mxJtAx1fiXSZLBRCBn4yWKNabJv1IZfoUlW+V1MNcjx
cqPAeRSWtmGO8kuDzZRjdYqEY3W/hU6sscLwy7VgobQrO5Nz43BjFldjZGCO6EnJ
M3FssbBv1bmKePC1BR/Tb/3fMQxc8t2vm4OUeni9NpMBlC31y8nkoMnUBVk6iV2g
egqi2Yo9dEtPpHbChrO24t11pBUGF8XvV6csM6iDMtAYjzHYCQiGl2Kq9y9zYYJ+
jOawIAUtsP9KcwYr1DwxWovWDzX0jXlvZbmyEB1DyVm3CoTlDCgJSCfWEFx0IfB6
Apy3S5tTrRRx4INMTRGVNA5Y6xAFEcK1S3IpYJQ6t9Q5iUb4h7BDYWuvg6xj3uBr
hde8B59gvT73Qp0bOIL2NGRK2M2QrQ0r3r32Qfc57EBXBAW5Ah2T6s4qoemhdw8Y
ra6+h+h73aQUNswDJrFtfg2E/Uwe5jD5yr8P7C7dgMkR8cnwLl+ES6QtDtypamRG
f6zLGZBaR1FCbKwkF05ip217GymCxshNHssVmFhJaqaGYsquPkOTD08qplDfsBFe
AEjWlYok3ZYril1PURMFazdCoIN09+g1KkXqYz2afvrTH1DsuXb+P++fFIK4P2Nj
EYwvwqJLAhH9GvXD/86LcK0hxf0QMCgnSwXHc2jJMfIX6/omeiuSA/OprLLQbKlk
zHE6/3b9/ZWNEW0ZFF9EfNsgNCv9jmT9PhCP3FUGLWNdghQwz4ssnRfbXJQvHOLp
815Hl/Zyo3c7xYZQ68lE9xseHf7Rn09Wm2JyOU3vH8j0TIAzLFO0OckhqBQtQBqU
lYsSmmcWhqBE3zIswx9ZmR1zYBuHUhxjkG7vosfbHNoZhR9QekYG+1lGGgAkduDS
kEQhsav4rTns2v7AApYUmZc/KZ6FOiswdEV7BqryMvED1qQmpOoEK/NGg0Mve0bY
ojueqM2w5V/maU/Rx5/zspBJ95NC45M+8mGPL3iyvpaPOyeFOgAf/gPAPhwx8qN5
Do1MfWT/FOyaC/OaB/1PHdY4KSSLRZcpwhOFG8LlMlkQIvrUtjdjXINr6vDsFn7b
B66dfpWKtH7VFMYp5wGK+qP+KXUqqBHkm4uar5zHhG2gmJHWFFfBsqdJDyJr6saW
EqHHerx6CmsuD+3xoHWyR6M+sUPYA5k5UWFrT9EhCmt56vRHEgRHZjjiWvfJbCCO
dwce2c61bFECjySKT9rfRc1wuLzWFKvaDlcEqVV811qXjWICFAM5rhyM2+1OxGnF
rKxIe10ISZRB0j63zaNHetF0Bg1L8cD8oCCNUW9gbB8Ryvg/eYdsy+sWH7GS+1kD
rs0x6q28e+xQu3Xh2zhS/18vfOtPUTJjpO4PKBOUmkLaSIuIH4Y8vP2e/W/8RioS
hqzoCkxL2ubyOOlcH1uaB2m0akIz++dCt36UKr6uBJ4f6vmV2QzsSZ8+R3gKo1Cm
tUDmQJKaKIfdUZKd76Td5E5YYRKhemswPieO29tlG21/NAxYDDMxBWAzTh2ZEFvz
V/7qQ4GpMIbVMQ8uZbcQmDdChqFhB2SB5E7xs3MC7ovWhdV/RUFQnPZUp6//8J5B
xvQ3UMpoaiBeW1yWzdZvbnKdbQRc9auJMphf9iu4DC7Vk3kyr3yjoLr5a6DyWyLR
xsok2jt/xODxnhii7Ae7O6gBF9eCGqeshkhlth0g8RTjtY3cEv8EaWH3iTp4GeyO
2D+/OBpwy/Q4HLCBiRq4X4dyR3H5pi8iPEBm8PfBMa76KjpJ2hR0mi6arI4BcaC3
cZfKO9xOT/oFEx/aKyqqAJF92ssYyefySGbKSnKNiGyXrmuUzTViCLGNbTqtBFor
e1UbqJmu6pHhRGkHfphOQM1KFVZ20dn7djyd1uGMuhkL271MvyisBQe3Rvw52wPS
jCkan8mnw7wW/RY4Vo0dcG6iHu/u8WabQAgd3eugiTMFNrfsMECOKiQgAA7R4xJf
tXPB+qJNJ0Zc3mNxhHnsOPaLtxhBNKC6zOEGZT8bjR6L/lq4KN6SrFvRZWlaSomN
gKbRSJTqXyUQjEG7lzJr9yyhCEM6xgSFbJ23fAldB4uUs0KCofiwWZcbkjd30nyN
IpjfAEB91tcLLyC6PNGy3Gyt+LTl6SN2j3Enkbt2hSZh25d4KQ7a2gLUrl9ie6It
vN/a+f/zXgySpUc5MJ1+QijlDTir9tAM2Wkzw4R4vXjgxZ5BSbO18miKK6PTAcbS
v1At2ZLjsIgAEg2ngJHqYtKfYe7W4J7Bplya/LQ0Sx1v2ORWfESyxrN6YUkF/pj9
1NDADXLuVaQARm/h1zNC3Yhb5L8nR4EGT44Aln0nZx+0kyxl5icH6lXIa67kkmFr
lQ8mbdao8ryPe9PcUmuhbAGvG7Zkwp6Km++v4FNFKNpuD2TQhH4IMd9p+fncUh6A
vyhRp7LfZ0qjtpNumxhoO9yYEIdXPbCYrLTPxsTvAjMO7htRJYw8LBihpPg5A19h
fearz6XGO2/mypIdTW5AtI2S9pSsV1E6fCjgR1khaQBuDG73U6UOTN0dBAIfHZaf
4Vvf/3z4vrFzyRvTSLGAcUpLS0Ewh1l/QXvQNo8+KNc7Gc2/YT+K4+T38zDnziCX
k1Y/ER/wdOMpcQfXisdM8JTNO8A0nk/JxBZc/cBlcNdGhMrkyMKH9vqqzsESW9Kg
evaqv0CP5SBBHO4QF2s4VxXXRyahOCGf98fNwNfyqs9QHzmrPW+ewhAE2GaIa4fh
r+wGNjR7GSxjp8ZHstFFnKI/l1rZoC2P4U3PrXhM+InQVJRZeGHR4uSQZLkcFrzz
Phpz2m1PTyBXzKt238WEu37eQfxbX2gCC5yBoWbbtxJY0Ht6YakTgelEifkGV+iL
gGW0MhkYssjieu0yIfFlt6v9KPAikddrlIkyJmF6ZKtruhJinXc6HpagiIdrycbY
RIKClXnHQzqf5zDqFj2l6DH7sOZ9CbHzzcJnNrlwjIKja96zb27pNjRRs9mtlEg4
QOUZb3nUmzvE3OMGrYypKbdJozagk3Gre+siVZKmcAbwFLBZjrGftSox4p9qGM7z
2MmlRobCXtqIbv2RZKZwqWu/epnH76648xrUMBs+x5+oTZ+7XC0BEtJBSvZd/PUX
B8+CfU3EeQmRAj4LPUhg01PUuSoaFGl7rZpm9Vy84r6F3CaEcawL05t6DNZyeL8a
r4+hbrZ7oQE0au2bWZZHgN0K5ph0C+REAwqrIoCZo/iTRksE/J/yt1HFEoJfxyEE
c/Mep8DeyaoZ4t2cNAofJmWbKTsXLUMq6GaDvgahRsJujTUEylxVZqe2Z1kihEH3
i5ZIImHZfISKITmlpl4xUBKbI+xoftlDpoBnq6NVxrHXHnD5CcECXT9Dxy1R6kh5
5uSSwwcDJYaxXmC5momNz+vn0Z3psOPMaSHRkd2w1oERG1g6AQmF0r58unJrY4Pq
nCUxm/e+WZeJEdW3ZgAbsyQYPei/gCtirlIh5mk4Fm4sRHZvOy8JTWvvmYCmKdlR
WKgyNLL/TvXzxMY2Sji7tk8EfDxxGZ6HtNJ5/AXGs13VTMilBYjRN30mp+SfIUrt
PX6apAXYHdfnk08ENRfARo3aCkUOYgcuPNQazbbUHjNkRnzqrVzWLjULi0tws5G5
qfjbghyzTJzQot49KkZUWxWg+jTx8ZqM8Mvm4sdkSGJ28NpqESl6uz79r/twDygY
sWHYy+Uc1jjeixRLBkF7uxrxddfrApFO2785eAZ0c58sjwZCimn4TTGbYLJN+4o4
cHIDJ4RUeO00lx3USOtmLs2rzpa/CGaYcMkbwm3Mm8t7l/lbXl2ewut+Swltux/+
pvPlI1Hb0leMavITrPBEavzX5zmSCkK5ODdHx+7ekbC8DgMXXtEJte8hkudVpqWz
YbKvWyUpZWQSFbhwbQn4clm7E/Mr9Othcr3Xhilt/6ibchjRfodoGity2rUcwO9t
iOThH+cVGB3mIaMAUl4cu/OvG17TIbPVj0fSt3yu4yoE3CIY9PDQul3rypH2kqTy
ETzFo/RAvVLH0gGcZjXyLOmD7M5gYt19mCnJwMb8nrpJE3LrTcl7H6Zw1dH0yvoo
DP1fO/Gp7teC0bgkVOBv4YEqAK5szi4S6G4yLhiOcKGDG8mqpyr19QIZdlA6ttuA
730egu0ZABsA2PLX2xop1sB4SqTq/KfO+aPqT93/FNZo5anHENVCGZjEB0hKdl2u
tf8laoH+xRGYsRCv8lOiwuuneztoXTMblpd50IwyPsqQv6jBTDsLHCu9rKv41qJ0
mq4ECwg+hqnDgTQydIrV/+RemR4qYVCPwAMCCukqtr6TJlbNW+Whav81TMTIRMpl
eZ85bj4iOa09Qx8kisr+SX5DVJtZMRXlAu15oEpLtm8EG8/e9sxVVqn/N6tsbu0e
Eve//IrKHhC7D4MsTl3LC2iGJPOlU+QaznhUN2r2B4ojERR/8UltAp8nnaC1M1qH
dAcG8FAgZbNgxXdyW+U4/qJ6HSr6ecgVYd0YlkMf5RdTUsNZ2dMzsYCdNrhdQEty
blOO69nquqow9hMtFADn9yiS1GKObo1tNBErZMrWgOGzo3xshsCbkDRGnV7bk/qc
YrOS+V+PT+xkjqHdpu3lGIdMFwBzabUmzMvCSwSxYphTegOChSusXtD0fZv3xGp5
hAywoo1+LSr7Q0tCLd9lu+cysWPCo8Yz13GNZhjb8dT8JjEtNbNOhIWBMjyssu8O
WEG6Q7xNJOPfQHLWcI5p6v2gdmhyc2lBnLlvUhV0B4uLS2bx8rurWdUpDHP8UiKG
S8Zk6vYa/psSmOhbTXaDrGV/e99EmiTvV5R09NtFzU+JCdavjpaZzcAQby+SlCKU
tEdxEtPFPEnDFQiD6sOxnaTaU5hZiijxxy6ogZa0hosKwMSIIWWXBmgSA2FUix0l
xjVBMDhyhieCHoxVwwmNfJ8QrLo3DMaPqQ4VNMVGwZVufAUkZ/t9mcZv+HS8EAN6
7ToNMuscJ6TPku0P3tb1OGR7vv2i+xkEp4xcFnt5NtPnA+vgQX+Fm/7/oT5yXDkB
ppAzV4TNyPkF/viQWufSz5iySnDwxFNn/Aquo2lSUXcMGXB1bA1aGyUa0xqrIIvb
qnxwQlcXssFYtSHnmo73tjbCSrb0aaLE5rqWFuQPChh/4UvFzHT6sUsXpoMWtVby
qL73P1VNIYORcejSYWw9do7Gx+RCkBbTfwPuh3qJHqPivEllOcUSTQNOJyOLj012
aJfKGLPWcuX4WX9gNEHgAcggEsXsRiFf21Esv3PJ9Yg3O22sxaXedLMCNu+HgesZ
I+ic4vjiYWFviIJgcvN3vvhHJDzdwtURoxMGdVvFae42tDE6begMh/5iQG+zh2b5
dGtxp+HeU0AThM9v2f2R7+RMESt0Sf+Hna2JwA5r+OgVGVnYK3a5/HbaEfgIthf1
iFXcDiKYhixJ8JRRJnsO8vIOirHaZmZ5Q4MCPnhgjsLOXANxBjbIrCAnGvIaetcs
WaVyvwB7/05v073l2qWOdNLQZDBCp7C/+TyeafOpewZCFNAAGHv6WqU1NimbMoX3
+lkShzP0lzU/dZbtrBe1qsbiX9g00qTl+7On53/kwy39bGhG8Yx4gUUvvm2D9XuL
Z16HbMrC9t4zzCZwuxsv52o2/uqBe/HwCk0wnFMbC1iLxEvoQ4cjdeY7e0mmNFkA
aqKWMGjYwOAO+dMJGWwCBTQMOMyyWHHp9DLfLfEpHibmLq50I9ob/GBc7xu8ywak
8gEg6OYF+Y5pgc3jqtqXu/RITzDuUIRhkCjQm0EJwhufkzCDHDfjqPy7cgMDQHBY
9GKP3oMMaetLQNQwFPqmi4K54t2K5UIA9ALkWGo7QjUNCHEW279hbkJJkJVv52T1
GYnHj8b6lhxZhePlhcXSsYtcasM8g+7EHXB5V/4gWe4ZVQ6SoJAhbT5B0M6QFhJ8
3AveV/UCn+eTCtytTEIyaX7WrgLdd0354bz+XSQYsQ3UHHoK8YJiYV6R0I/Ty+yV
mpv+Wpoixice54ooEIzgWf/m6PCZlhe5mi+OkhuLgOwGe13m0U8A8KPM5Jg+tDIp
zQISLClJz2LctBrexcHQ2MTkO8oPF94FxoEQ5STpkT7/fIaY+VZBgqFrh/1RYMQR
R4AIIfnh9X+83ZtLTlzF0fg/pS82KXhDZEX5wwsJvewN7ASxCNPIzNoCThnu44ds
LpFbEpCIxqc4eAuMji/yLsYBO7VRt0UuuRcJiqW8J++2oN1aZIQjhT9yynhrfmmx
62rpw46LgAKHvP7vODlesu31UzHv1m3c1Yd6RzCmv6fRN5lHYXSjNmezt0534cao
PKdFXqBorSzVgWCZqGg2y0q7QgknrLKto9LRfUPLruYcacYAXERw+Xa7Wot3IXEd
DghZak/j/cflIfPMTx9f8hzhd4ePV/CcYWTUGtzHyo+EJtlhvDW+ynXPzvM6KBiP
pAh5rOiSHlRRAxZxbKM5aTaOHY1PNrGRaSFA1+NRGezo112MCW5D5Ytiri9YRkeF
x1nWKL/CSse7VMh7pxGW223885ssLyAgEHrAdcJ5kPigLRIzTIyf+Vth2gAma5Xw
rJfQVKyoGfZVkQ1iNqfSQoc21o9T8B1n+wrRsB65ahRdgC/rcBIyZ+SQop1Cn7dn
ghC4reuRd5nZw/ytvf3epG5e+rwWt10vFgAhoFjX1pv5OZEAz4TdaRDcq/mQmDj3
C5N90vFYY5Do3E6TYkukd0C+tv9SWAF4jsy2CJbNnJWkZxOBul/I7NAGWd1kAx5R
xElZTf0oTFgPOrol73zvTrZVoCZKLvJjsNPWn4WKZiW/P5JaKpcO5IG+WVtCHxBE
mvyqqgrr21hzX3nV83fDrIPfWZ+WMKmylbW2vb74AxlgtAp8ExxYsLTWYwgpmsOi
pC7wWcQnFiS0EqJ7rNNlcnCzMQMZrlb39KfB9eirWi/LMIAq2C3bkAyR3bGYHOH8
MNkAvgZn5rKRIsPh27qfy9GEc1OT/nTMAwuAYuJgZXJu+qTEUWFNf3hHGsLZs3VV
vLitKB56VlryyX4VAPSqLeCTM0YlAe+pfajAY/PxaDM9+SXRm8dh2XLxyKfO+YAR
MWy2t8Tl60FvxCMp66ByI1Yksms0ksG2jJz5bTEgiJSS4vq3t9xn8GpQEWbr2/77
lG/KcT83+Hah/36TdZr3BuVZqHpgBNU1VEg2Tng8HHetFWLMZqI3M7AcpSz2xRhz
TZdD9Del7e7apWCwILUjYdNRlczd4az1KjO2BPPcG3xq2PTn2TF6d3jTO+493ck8
/+RmD1r4MdocyEMzmDnWgxGRfhJtKYlRY3reCauniG/DKqyx7sW6uberfh6D5ZKR
rMUGlLq4DYmd4TaEvwcGhElLC+NeQuOowed2P6zX5BACae89rMFZgv1+pmjCJ9QK
W3YvZv2H/juzRVPLC9Jqy3djkSfESbTU1Hnt0GQbNNlC0/PCIKZQXOpAqh0UFr0b
VOfwJNumTTVPWH0hHivGLZ/l/3SaGCy+nEUsod1SOhe9NQnxxDNtzzFpIP03KDDH
ols5v0rhCsxb53ocf6ukUPZ/Wd5UlkocIY7oI9byMb04kV2YvbuX80xamFhUR+Cy
E+lRRNk/amQuF5qH1QHXl48Alw6Tb+AgZGMjFylN0ImUcBS1LxZhwv/kfx6TabNU
vSHbcMigpe47zZ89jZ58EAA4KO0ibXCqt2BRR/aR8UxZlkBU3JxaketDB5quAXyj
W+vv4q8MBX6Je8OQaULoHQf6UZrapFOD/fFn0FpPRadp+eOsFX3Gyk33pbl5Z6R6
x7wSH+Qo0kwLMouvk01SDjKV/kJUt9JVQSFcIKJRSmu+SdBD8dm6twvi/ltPc08f
WlAIR93OEBjm3pa8CjkLOeCXofwxeE4I7jIuKb3vYEXG3/gfyzze3RihiapmXQ0t
zrvrbvIrVdex2fY6PBACB4Rn1i63RBoYMa9xbfyj7PNYJGpTB96NdoqKK/rOIBM9
0W7cocjb85cuqX0EVnR8tiwfSg6sFlKmIVrTTZJWDUWLLfI47jaXohF0V7BYCqcp
sP0mkBxgdXpVJ0lr/F4bGTcSuatmT6auuPAY9glkWFLNBd9wwqTyZvyxoz0DutbU
MK4BuoG3+1cx2FhFvkfPx4svOjElnWWjAPGXVB5Lar+jsblmluDBBmM00hW98pgk
BIrrolvgEYo2I5wc/mnb3yTZucaZIL9nW9J4bEb97tm4h9nwZor3KAeOG5xSPo+h
MffBGXFpqKNQIodMhNdWm90J7uingdvc26a5qozuyBsdodwxF1Q53mTTaaF2PK0F
haGQKjqe2Fc40h6ccj65gZrNj2nVV1nf0YgPp9jtavuEy+fm1q6GeH+qe0Fr7L8U
AtbnlWberr+D8ad+3wK2+lSE1oARhH+GErcQz+nNEa0E7UYzck+jY0lzP6Ak3V41
CW4SEjvBzYPJI6AIRMRYxM870JoQzOWQnsXWkFeHkIYzVjmqyymd/ShCW+fnpky0
iSA+SKaoVORxGln0Jyl4RvCK0OHJBK4d54zVcrkQxXhDoRTnWB1L8IGt6fFWkWDp
a8M2bQ3JfMWYydrEIjnbOmQ3FT4CCdhkMX6UZDFkdCkH+uaRW+P1HW6c8VpnCnZK
7xzusOp49Enk7S1ICh8ca7X69N784nrXob49XwCd9TllvyeTfupJ09YABU2BZdqn
yHJTvBFk8vuOgaorH9yBV9UaQ1GMo7TUmTwjj9o85HYJZCIzhkWMjUfYWcnArElx
OKs4Aawk8ygbDmamxcH7pYs7ejvtWEjs/kX6Ahw4NteKCRMHe7W+gQq4q+lhLP7Q
z3PQhCZmYzwRJ1EBNmf7GnN06FoFbl7Gz3OxBLsUmtEQbpUKTl/t7tUPBFRsfsoF
M+xyEDHcdAXJd2m4M0fjMmrtmNuVhvOyMM8c7rJlN1/GIEmmY1SR0wuV92wnSgU4
vAqCGutOsNmuLPqrQvWcMAmyOCgu66LioqCvxxSuop0M8yggzjX8Vm1MP+O4pb8L
P8TiS0zmKCECi4NN7Yix4ZwQ+f2tq2RJT7dG/nWLkwX/rPIlEFum6eKvQX+/hqzE
z29QsasaOf81wu+ODZ186M7BXJHOBtYvOjaDbopfSXhfBBJxwclpw1qTFWcyjStB
srO5P0g8sOLkMjF8ZZmeKAvUZrpvTcicpvs3jd0ycwu4QaJVi+Z6b/7NT9rVUrHn
CcyTCmmaieOJJLsC9Whe0MRS03VSNji5wfbWqrS7xBU/68oZnjVARfNfuuyky5V4
wspmSM+DQN4ri2pjMjdDs8yJEqj+UCBW/Q6kg6B2W5vqvWp5OyeHfDn6dLVtMQ+z
fVB6a66/It2N5e/PbUV7+HdxInTWbqtLVHgKzZP2dnSfP7DWNdIBUQHVvAbEGmBH
URJWvQ2HkuyFftm8BFxl60vd6FxeGpUQxrf2JSA+0wLa9OLFYX/+IgRjniVq48sP
fKLe/f3BKDXk81NeJ9il6ZATuzTqUOM2xDdZNOXpOVXVo8yCrZquk4tg3CxzE6D2
FyFsIuxhJnaQTYRfTAKSQNNO6yV04HQtL6/1IAp7W9pW3ILdrZ7O2XDukLDH7qKC
rYzW8kAFFmGfNM4dY8ic5cf8VkJ7OeAK/vwjLaUHfcmyNArEUNPxQ5enNbrv/0C6
iqbyce7H4286+zAw1C5NNkcBwO2OPSgZLn132DdoJc8P/WL7Ovv6ucShSL3xiixt
af28t8ALiSINkwgItkEK9qZrFbgdFUghVtatH9mxegSsMaalr46nd9W0ueeO/Q1I
0tG9OMWvj1sNuuqAOchUCtMfRF+b7bvKB4QUJb2ZVj2hyNs/EQtbzcltlvL+sV62
BtmshvyCXMhKpsWZKs+OsbUO+Ocrqj1jL7PxPlV6aphd15qVcFh52IEt/Duij1rC
u+uXAkBdBZ160RfIuPAOWK8srQZRJQUmFigOHDe5KjC3Xl9Cin9AN3/4tO1GoQLx
otpeE/8QzNZVq398vVVH2ucsywij/hDaaQ01FODWKrHd5bp+7WuvxdNr13v0OdvQ
WxNwVlaOaogyxMl0u6fuFZLjWe0R1NkYCjYdBBi30mGLvx3gIuxDAO2r/A7OnYIR
x9slBmabjwQc4wiUqId27uA17UvBx9ZXn2zsovI4NEa6zWPxMOeVqhcNkJH8QSUG
eyRyxHR5ynTJa1SGSLo5YCfR6CaNokFrSvqTJmRpr6KbrnWzIHEAxnvWvutEsGUz
jm2M6JFl+Ho99DDhFBfP/nuWZcO3cJuY9khzwn2vMqwamSyzv4N0ctGZ4YjcKsiY
2mfyXElbvPyHRW4gUr5sM4+1jbJ/VUFo4DxpaA/HGIO8EGNsgpCqFqvDiHEK1eXQ
xjsLV/uRmopYfgmnBdLy5q4M1IhVTU82o1RYKVAhPJsdAgn3Fi4Sap3vxANszCqM
mWYCZAtU93EuYzticu7UMepKza4iomgMQ1ePxNfVR4u7BA0FfnC2uzYjA9KuQFnO
Kkld6WN65OO8C92VCk6Pj2WEEbMf91YDMoz/UQKXox1sgPL4PZH09Tz8DvDZxRhG
asbpTrqmtRz0sEl4lPFcK+kxDxuPqbvq4woFXtErNK33NdWfBrsMtwnH8VMFXJi9
fDsQuvuer8Q2SapzMRf/fpoOOjvHtAsGm23uDdbaWV8idQ+Gtg1xsSCZwUgw7j10
N6vWTjzZakb5HG+rKtbCPkOaJyKbR1ylrAXGDRNTMrqgH8tDdbdyUKvvDAnRToIX
U/HeYktCWfbQAjhnIFRH0gwDfWS6GQVxmX6swGMQI4YAgHK+UA3qaHZO86h+pO5/
iI8VWIIhp7l8ZXRaf6BLWB174Fau1HHf7jYfbCUXrTwA6tJVutVojSW94OVWY0O2
H0+i6seHEFd2whiQQQ2SYlVRdfvB9v1i7QUFN0TV8LYzGGSCjaUY4Q4Wc9VVWC+I
m7z+GSoFLenEb2W6A2UvPJMqlEDxPxBYax+ybTTGsrOUF4oCYvk0oveD15lePMWv
0qSNf3fkmVgPdRe/Ls03QqFkE5QGr8HneFTyPmMRPYjy35kM8WxmYwOeyMFGTgXJ
YZc06Vw710xlnrt0G+hrUbnpzFV6RjBrju4AuBHV3H0xwE+1PKY2KZXBp9M/Ziwx
ZTp2HDFZsU09LDpJ6GMrvgQJUrfkh9l5MV0wS54oJ+pve+vUKJ+ybs1CfazGQ/Yu
WdS+jed6qmkj7+lYLj+3PgYxec5QazUZqJCLp4XtZXffAYpP6V1dCcrwc+tn4xCB
YBF7SSimMvbBhyCC74NyHVghA8gR8AUWVuUeBtJL4DYdRAlYG9ry9z82gz7XhtGz
vhtMqKGrKM3xBKluAXdLV5KJqh4xFx/3oDCCvn72WjxAbq2NOQmAGH+rVoDu7qg+
AVMfrHv5psm5UWnyRVRZsla6y2IhRohDegrOUeiqcgaDqZTlh3RwuhmkkPaLuj+r
OM7/v9CCDT+U60NTbNXlYwgpHBPAq4lPt9Gd+RDiURHvcwKMQZLvIuuwsVsKpTDf
BwWr/7XnrePWCQSbxNvDDVOEaRc5kLffhD0Ggy94Q2ZSe3KcivzXi6fPcdy8Wqwh
Sm97EEWgkCpKAq9Y4+fyQTGIcLR3YE9QY3CzApH78EyjWHwfvu+gbC7ioZ7hCDdB
8EYodEJHAawvQsnYlv8y+ZwalzJwUkbTYgxqTpLSp1LbmR/gSjmq7AWlEn+awL6J
CTuCsv45xUv+qVX2rbUtfPQ5gYerlYmIImikiVyHThcfFmQZzrcBi+e0VhJuARsy
LjfghD8WRcJgdQwCDvDA07ARmgA4j3f2HhpVlpEohJiYk1w7JerzDy56HaQH2tcK
TtEREtEhBAzZ89ui4fGUD7ntVchdyvKdvKD3ugFkfD5uSTl8qJMldZPYUnU6f0to
8E6vfnpfrJ1KP8lOqfk0tyQlpogOqSMaPa1+7je9SFLMTRJDvUgEiooug5GU2g+v
qrtp1hSg/hMH1rXJEMyP89RJ1rxP6FdxDcxHH5N2Ca4K+3iBNLecoMCg8sMXBWHD
Z9t7Ev0iAiAu0RcxHh/o4EYrlTzJ706Vr3q/6NsSqCIzdG3EWPtSOR/t4FOutFaL
0pZRkzpvrTlK0ktG42vOaIrdDb0ePwoFR5VqQF+4EkHlyolL97PnD53m6uL+vxYp
wSTowYs9Bk3ll9km1vN2odwknTuOogFrzyz+ZuiTyyKIeMj9zpeIQXX58KyuImc2
q1lbcyWgHft9Ol8CMM0PL4dk7ab1SrHXx10Dffl44N/XvARbqZIO+8xaWcPit/Rq
mYvpDfdfBmgwH+d5OL+Vvvq+6sEGpMXQy0vt9sqC5aZMKJ6oTmRMHxJ99QKuO9wc
+aLb2hcIqy86zqD6nqBbqF8Vypd859y8ELQgKIvYXd6uiG1CJGqDGhq8lt4M0V3q
qoGYiATR+sPex1TeBcdYJT1s1lGM0vFvIGzHB06xD9Bo6Zbfw+dSp5GTNaQwq90l
Om8jnWtP4K1veJkhL1miNbZYjLY6rpunHncHYH6kcL2E3XrSUNHllY2glItnetZR
VDMgmkUZ30Lrdn7lWkFy4rRpanLG/6vK2pyrzODUB/qSUHRVM6V0vRuzT8ZYKNu3
h453WHm2pLhPGjS6vfBJDnt8/lUrsyZ5j8Lf+3Dl+HKN4qM+8bTpJ0bsCZHKqj86
VminZvlkr3Am+7GFrTKeGYdM1r8bi+stzMgN7mJKH+9dXXbftC1FlaEuU+ruF6xx
SdfdGDXbWwVymqtr5jYCW/JzGlMrqXl0BioNSrbL5FxJiB3pS8GUo7H40QWxjnZk
dBX3NHEth+00SNyoyobsqOVHC43Z8phjgsR0DGNluc1Zkcr7A6lfUZThZ31d5IGT
Y8RcPFjc8EuOVNaITwW/YHQJCDbFvA4rlOGxwD1GD7IylqZuj21r9t03gZeE8b/C
RswcT222OKGJ0yUzEWXkdRnTiff5yxl3IiyJgbYH7wkYRj0vhMrTKVwLnKrfslrP
uLcT4NqKuHhk2WrKCNdEaOCvqnv/zhJwVjeJAsaJnOm69ufm0scTh/C6LjihNi++
lkCqVPJ7O6W7u86j3o04G+lSXEeuslbkxooxHiXdN1aSSp/dnorSa8kkXPY+DRn9
0JSA+qY5iXGngwF/KRhYfucOA4e2U5QuDseVZm2wB3LexBI+JLhImwAiRhUVRGsA
wnBbuN0CAEqtDW4C00RztpPWiGC0NEb/QPzktejxeDAyk7nXGhHdTnzUfDdxlWaF
GTn09gfAB0VNatqFoUj8/byAus3trJ+S1Eihj5QbK4Gxxv4YXhBndYxH0Oud1rpF
UQWjD1pZ77LE43gn9cop8j3driB3Ctt1jaeVJP1gPhLQCmh3nzG76+lHTtcp/F1e
3NeSasCRw//ABT2zNglH07GzNqqTSTt15mn5XVnZqqD7RkQSyxzKop+OjexpnIHG
TeBqKulX9mmYRyGVm0d81HWs4FcgbeiWhYCYMqOH9idYWRpyzi7Lu8uZUJkBlgek
IhDJJ+IZPQaXik2YwSl6VKWol2xF0NGPpZFnvYiriCG6IL5cn+UprILnJHRL8xkt
IcbV7XhPh81qUa8rsQJM65fn7dcN52n+WcWSyygpznFqCGTyQmeSwPrLnqBt2oi7
UMT5/pz37bWRfdlK/NQgF1Mr+0uFyQ2hLMX9YkfIfYK64K4sOBVd0sOjWauQDUuo
v/gidlYUNgsLWY9dDVKO3j0BHjA6byNXi1ULvK6EfWoY9weBL5rFhZ82S6Fvfvg3
9fCnka8N6RaZCSFoib9PHHWES59YCm4+snAkYeOn4ErV3lfQyfzm3hSOtEYMW2Sr
Q9ROBiHySZwTLhPYMNWMpM/ijueRX8VtuN8bDJsVDAtsVlkWxz5SWfYCjw+Jf7wM
As+57zOO2xKm4p3pXJ/Ymwtj2AggvTorBs+gMFW0EpFOyeX6dzziYVnGKoWzkTuI
SUFjN0Wgfayv+PRGi+KverUdlAWZKUo4LBxLNq9R9PtFf/JjsTayX0iAJtN0kHmj
3/peJK7fLHrCuQ5/rWwIhGu8HN1DxJRTL2PiR7JLYpB95Qsj1VZ7egWhc9BtGPlr
7WmVXCHNUyl42AIosmNYuYeyHUv05hVePVTxy5ChOf21iNgQ/3uKToyhN6ZY+EKf
ZhMJFQ493rzj9qK+vQ9yyEZqbPUKudxhP5xLMksCZ7Rah0eRBh9ltvH3oisfgzIR
J1R1E+qQY961vHoV97jCd5TaEzNc/tyrAprFH5EXsEmfdmeLgmoSEN7ujNZFW9Cm
NTSVuMLpTHnaQ9ow+2NsiNOH/LYJa+a5wePlaSlX/8N3Wb5OsVjwWB5KskSHhG7Q
zZNtwg1vP28ErPtv7rRCv8IZWI1dlfD8yBK06iAQK+s+AfYirfveFuZG4COhi16w
sPXSUu1/CYNC4aC2iaBNRfWZrKms4Qr3yaYisQA/+DST2TheVT2nh9r8ag5OnmR9
u1Mpyz40WkGaOSKIYt4DwUT1sxLxSw+/qUUZUTpVzE5B1loNaeOzoma/9h75zJWp
qLF5WInCLBue8zmU2kQDr3XJFP4VthL2K9CbXY2qBIUXtVqDT2vwaoGIHNBbmqok
+nvl5dHaaAcoZST9dWZ7MHP8NDdM+3GfJpIAVdiUSfwokDhV5u35tvhunXdPnqbH
gNq+xzY0f32kxWSssf771NdiRrZUiEn4lp6PTgDyinjKbsB5u/kDhxsovB7GRZfP
eMxs1SS3HVIXDxHg7SNMG/sHh8lsAGj3xK/3mWj2FSwPIREjOdzoQbyoTI5f7PWc
f/e0ChOSySHDPLEDubMleDhFvQxVH0fEuwhbCVjc0VADNwDGvDruL4Y9qpl7QJXY
Id6GkuMb/zEsKoTpxyujqcIkqLiS+5IuAJJPiQqL408h0dED4LZOMF53P/clTX+J
WWvtjK7QhMsdEIvu3yCpKOmdP0vi2mEhqGy80ck/7+TO2JnY79io3pxZpkiqf3t8
IbCAPY3gfWJHpzvOgmEvzMYNy9/gfK/VVN0Laa6ZcYO/kxgD8+E+GXQdaqUH8eaw
wUlpASudmZjV6w9woYf0SYlxiJu5uhHRy9AbK5WKD4AqOPPeVI+05lQCKQlBhHps
jwTET4rqBgcoqBFx0SWbRTERpACwV46MZUeuK7SQxA2KM1nv5FnVND8sU7puReiM
LMW5X7Cnqtm/06nt++koZxB9WrdONWq9L3sEXltBL6ghGNdNVM+T95J5J4YyEsoH
YgUNR3aiwyOqaRFwvNLSd/x8D/+IVNPKnKMApQQjZfNhlokgo0BBL40Fw01+NjVU
mkKj5/OFiJFmPCd4mUOtxGTJuFUmJh9rUaqlkCteVsEGTUWZ4eraJCqIXvwkD3os
0WUeH5ReKo66MVZ+xRZ51FXFakwWZmMM6Cvuxa3sfIrChdTLAbyRY+LZSjDRr7JQ
FrxqEYfZXgS355Fy1hu+OCZyDkn+6aI7WkQDqc3I2irJY7EvX1e/nwKAyKy2Rbb5
0T/22X7c+ElCMoTn4ENx/HMb7zv9CGgeRqSg8K+tGAGGnquJu17dFhFvTl1z4y4e
y86/fS9ltZdPLAB6EhSj3e+wO/gBiTd/PTNAB/m9ghLDiCzlrts9aFD7S4Sr57nP
vYA0RhEOEAdxFSiDJ5H1SLGZQ0iGOERhVPDsJ3aSnJGkLIo7Gm8j2SVy5Jdjb4Fp
32koHWLU2foUIqvGDhsG3Wdoov1WP3nKD022sjXOkh7lfpKyt4zZ7hvASPVxWbR2
M7qsXCeMJa6/CWlE2OVP7IcxVa9RtrPUH+E3S06fZSxTiEpi+pRxjNX2MuGymlqV
XTgwXKIhG5f8+Arly//wTp29bGIP3EqqE2frz/lC+ljoS8yFtLAyp+88OWeqMifC
IvMAOHEOdKmwVxtBsUesIsGQ3khl9wrKOPeWgEh0AT8AfYRP9KSCm3JTBpxUkO3R
Ygf+s7XkdPs3mwLU5jgH0qMaHaeOZgK5EGIyUOjZr0lu7X+2GUj1RQw/9DDOzPe+
Se5iPsmg98G22Ne92wikJqKrMKUo3SBUonBVL7xCV/WT0XqVNwRglPLVIp+62IPN
6BXRQ8JbkYLej0TifWN18nvdlOjhwDAssuGWX3aK1FQc2faGSTq9YsuJns9YgSko
YtgqkYK97PXSurvRYiXd10+POw3AEr5ztoXfyRPyDZE8qttK1NIKNMszQ64VLXo1
h87mKo9NjAH0xthiAACrA6lp6jwysn7QxJaBfNjjmo4IzKx+gcXec+tlXrUJFdhr
T/WId0y1JaBiHKhcRq3CZsgzlUkI10uBxjgEvIEZKUMQftlQre4aksDn2DW+N+qV
E6ncXvyx/3QkT0yiwdEIAIgUcTmzrdTC8TxloaG8bHx8SHMhXzqlAuglFmsVjdOt
uT4z7wD3gOpWMMWjDW2WyIe0nMbTAEaQJ6Knqr/NqZHAKTam0+rZS0mTHKx/qtEN
s8c/Adi9btONJMFzXohTVmRNI/tO8aVYG7qulg64Dv4ueLgIs/SpmrTBPzug8E95
GiLmyIL1ySxAGCjGMfBYfgwYhwyVqEuzl7JthuhHnat+zRXsSDR9NnH2ZZ3a64Te
amjm23vOuOmZy6PR7cu0cz8+rwogamqWgidGMUcIjy2TfDISoZr/a9BF86skpuMt
6SzQes2BEsVK8lyTw5PeXV8FhN+cDZKjyDhXMJwn0Ty1SvSDQEuZ/5/TuIzmGPPt
GSlruc2SRLcbLQrGm0EENh+vAQOI+wp2slyLTVr+GePfV4YSrkbbty5wdmIzcytd
E6ioeN8KO0SNvuHHR6jDaAGeFTccVFo6ALyBN9HqkDVLt7KCmF7M0KRvXAx0Tb3n
TqL07/Vp7lvnVRtC5RmPtgUc3+NbiHcBaMt+q42FjOn5m/XfFg6U758Vc7InBUZL
WizcT/UoS6mvOa+al6SkkCGjZalHdwzx0ZPUgehVHwvMAuCKJLoM3y/IV0omc3WP
dfqcgX8rkNKb0BblEK0bYcGAhAIVwxFOwpfA3fo98Qvf7n8tIHmLCF0pmRidslUf
QQAk0fWCTGKibUOX9cIfNRrn2FpaGYRr7RdJDQ0/EouxSJVyQeAXE3UNpllzb0+u
GeZyVFd7KneZydKupvAKhldzNOF5EWdiQkipa2Zu4r8IsX8Mg3STdy3ZXD4oCUBT
tGgUEcjMFki5AWWpzxHrJgxZlCFLGPCp2qjoOrybcx2rgU7XBQW7MrHCzjIHBCAn
4YcCnNliB49H15t4uBMoh3BJPKQX5SpVnpIrc4cwRTpXMZebWat77gD+S4pNHfjR
6AUiBGVvt+/IC/4zRsHRrltQqFijpUupw9cdw+5NkGO4df/9pyDmAYIdn6nL93jl
uEdQedwr9VnBloKMdt24NcERam6NuKE/ZU+4dZl7g5uwM3wAeDRRu5CUF7wY2J4L
ek7t+BqzxE70PhlBF/wJwDKQhFJRPzBjotKio+EfjZolSzqcjsv87DtawcRgtK/2
Jt9JhgyhHQNGj4f77in7BLoeEkQkOv2XF9E+58ryAsJ75o3uzoiORCLvVlg4A/ul
zF1jGNL5Gz9iwvp7DXQNbLjUzaoJgFQNIrWVRBRgMSqeFNKGV95yflMWWPFCo6FT
MkYI9zPFNGnB7oHfo1XunCFXFh8ftyadomgN5ZCQ//8idoQdTdp75PxC4oTMbTpZ
1mwDvF1ci4Gz0FYdHf9VDrKkQZ9uh4kH/OpjjFMxa2JW1DCbioaK01xAm1NPRayc
WEpDTWVhbUqicMQXCO6iO6+sLZPMR/4bDClTbRgy/7IxLOicbRFz1kblg9SN+L2j
a/+j+Abul4+mqoPWihWmuYpSTupSqQud0m5S4xhp3E5sijPX9q3UdvBWP7pFaHrr
1/OsmTXKSK1xaCMjptoSApjf+dSDoB4ROjDw/nBwJ1ntP2J0BatRNMcZGq/jIb8R
OJa9I4M+49aheUE4COBx9GThIbi7mUnzSBUn1yV4joC0nBlTtJG/IVM4JI5FiooS
vi0nLCW+9hDX0lWvqsYxhyLZCHyqVZUt/zZF3FfO5aI+TyXlUw8c3l6tIwkrBduq
Zy139WGLExL0TODNeveQdPF0qeD6+6uewlkM3f/lFryl4ahD75hW8cBIgm9WRwzM
S2l7ml+RuzQ0Pab4D9C5UHZjl8INrv17vIER1KiRKDk8HfINar8FVj53aUfwK/t+
9H5ZfPlGfFg4WCCKwdM8YxT9rDAIAEjSBOXj20CPtKyrOUgvGOj/WezUyR+gq9GQ
9SC2wwdd/jLqmUzD+PwKQtx9NEiy/ETck2bM1f6FqCuIIDA54vfFP20XjAwASla5
mNuYkmVptZ+DVz5R05ZOFEh61NKB6Yv1IuvjNtL62GvGO7I246Ay2yunpZVrkMqm
CgQcmSOuOdB0drsQ4Z2AUYDT4JHLKx/Yx8IU22QjpXX/ZEME6M5HFb6SxT/WNQ2C
buh7Kq7f7jBm53oGAaJmrC1DQBBTkwPW6QoSiFOdSa0Jfo5q8+fSA3LKE9ul8AG3
Z5WjqW/r0Hc88X/EaMKLluxj8mf5aLtNdaRFvAiFL/jjHZbSRL6tKcpraZdI+s82
cTaQBwGfoqmW7z/mp83JiwVcBGERTKczshQg0Nvbxl+L9bYExSCDDZkZ9ls7Qa/P
3CXG8iRVHMcNm2GrBHd68lAumvQ0jpioI5jyI/7kWIxSj2avE8ZINLhPjtvzz0o5
2q/3qVaqD9AML0nRWwmMnry/LG0lfqt19EpiB9xnYmnzgPbtCBPe/IL1ipOwps77
/Wk+Lq19rws36IJsBXT75olOXbr/tA8hK8vJhxczBGXgegk4B5+MQnce1EWIhirK
du6CurExBzgZF5dyeCgHLXA7hSeVRATFnbTTMCSYPQlADsmPf9Vi9axJm3IvbpYY
PUVov9zU6u6fsDgD+7IvrmZd0NTmnlgmDQGzh/cWImaQmGLFEqAIIXMkBLJTjpIo
mvdha/XktrHMwCJJcvjsnhd+Fnl47UgH8knRC8Y8c2twFNeSAjit3KxzjEMdbg9T
jpOqylLS+YmB/sm4pHv0evEAAn0dYYe9PNIN7M1gDXk=
`protect END_PROTECTED
