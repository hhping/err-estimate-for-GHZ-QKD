`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FWGZTwzxI9GwRsEabMBP3wbmEqrElO3CK9chTRnVE1SzuQHg9PRBUEtddFsPLym4
PbKxVSNzrcGQtbfQsQyh2Zut0J/eICdarQnwzjSZz2OdO6eBaFnN/LQyUxj0I6kz
KbJg80wK6xD/AAkZw17ygFqfoshX605TWCXekTqpBSPqo9Xu1BcCifcMkM76+OIF
/Mx7ItyVxLZ+8Bld3yjyLU0ymfaVFAgDvEHkLfP9w/cUJdZlDVZwrbQNS6ygCHXM
jnbXDivMN6WqwiOnvRk/J2J7Vxz0e45SmkhwWxb2AazS1fYgLizkGIUFeC0LoSIO
3VhJOiWEIOsKxGK0b3+vvuplyCukNgkMP7YKrlLEJDdBDf18UXfn+8ECW3Xnr7+3
Enuq5jELIKQDlHiuMOfU3nPND8yN7ZFuZnB5OFtKk/jgiBzXfhloksp8GRyW53g+
nM3l5G6qMDKiQxZpNX5HNOuAIattiNB3K/ZwaJGVm9p5o/5YoDRstDLqE473xlZB
8/zHsEdz1VOWkHmwDqjVuWUMCQB0W3ylB5IjG2TPbIlZsbNExJiNCQBAoXzCd9DJ
nRasYJR0aUUpkzgrn1Q+fcOxGZhX71rbFBjEOo91UfKp0g2LnlHtVCglK87juhiL
P6AcO4crw/J8NEX1H1ByM45kHUfqBMx0RtI75wsM6RrKMQK5D/WNR8H7BFOWNTml
lyTQYiSfURD6CqLf2amwl6V/Ay/y7mtEL5dVed6+CAtJmvv2lRi1c5QelG/GI/i0
7Yy4ddRXqTrvEqoPYpP2WFQYZdg1LG/VdSRzwCL9S0iud0sBcF68R4jOmYsEDx5L
GyYZnq9mcat11OCpOij2ew==
`protect END_PROTECTED
