`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEy7LGVYPg1K2+gE8oGpJk8VsgTTl5UoGrxImqz5gvG/aoids+cBEAuv+IOz1iPh
okm0UVUsgeqiw5EX1tT437ekaYaJbnJ9+7Ob4+/mkS+RWMFZqd2z3cAvubifCG8l
RfRZF0Sitohu1bhaMJ0CZoNJx8Rn87vZnPAxoCUb9Lr1Tmk3l9zNdWahHBOw5/z5
2rGCykfx0fcFZttCOq5ys+tA50TN1VTptEVdmIOOTrfxtfkSEa3b1PCmFuU+xMjx
ROte0T5UAR/uzS7bFQAGp+rR9HZugndzh46duI0w9gS91fOLzrEB+xDtP0ljTKV2
Ln5PthX+y3q9THr9IE9j8KBEW167ZIIpTY7870yF9Ee9m4GF+z6QVIMn4JNMF+/o
X/cUgmXo10KiZsdZ49f6gjwc9SDu1AhUBsilGXtTICduc0lm1QTd62LFBqQ9Qk4c
zmSVNV2CbB8AFRtw/77gopb+q1xD3njhKuhtwCB2dDaIO1uhhc8S4lyBsoA4HRkm
RQapwHnsQzSwo4c/xSZInohijdUhOxhZUXCBH5HRI9yUACRfHp2rVtMPo1l2JHo9
Kjw9veQZODvZFhrrjjyRjNL5Qa6d8FacbVhUxsScaU15eAqh+oKM+sXPwkNiJbgJ
6TJQU/3mTp6d6/DMJXZoAyTQjzNg1HcVfdO0N4TY4X5yJkE53ezWqRiBoxd3t758
VYIwQ/7RR/1UFR3bgCpT1/xtrP+lzx1pG1Vzz0yT3LL+q++VsKoCI0BvBJcYW9dS
kUMF1A/Ia3XtdM8FIRjnHruWae9lEvGVb5L423Guz6E2ewl6XLgLOd/W43uVIb/O
nTtIs6867vz9UL1UU/8ts1qXEKwDJNdR1NEQfR8gvsHgZtn6MFOOzGzMVNoKkpHo
dv/RK4ZZJuz8575wGRUPCJ0HLonVlx++xdDQMoEXpCWtTdqOzsBSeL8faWeNkuD9
cJ1qXdwtUJvD1k6NnMyY81QsOoupgjG9SpN9+Cy52qNC2Oyh9EJB53HjuCVRUYR7
CVUKVnEzxB81+tJNeU3ujBXV9WSSF+rYGpLoGrkkcdvfwI6ivy+ZbslALhr+MQon
0RlqAhBaO1VahHSwoascRad2eIpxV7MRFjMRLhLmsTlXEQeoi7aryDwgxa/MDwDd
zGReNewN2KZr3N6u6jAQQESStCm0sAk4cpfFeZGAi1tFpCqRshUecvzKKnEfdTz1
y9HpVR0+cVhNFO9lHlFw6pVen6Ne6Ypa70AB+1DxJdxJJkFp623OtgcbAfTu2FRc
cIipeNs/qViqrdZKOzaf+Q7oca4DLDiDWWGe/Tms+LKTJHuViej0Jz3htT6gil7h
VDV0bJb+rzae42NsAV0lUPBaqeab1FEAwtAUqWYLL1KCrgJ7136+ftKUXtdT1012
rz7dTFX83ZbMb/LYfZENcB1olQtHpp/DTzyTPL1+taAfSh3wvFgFJjd3oHE14qwG
E973KrYjNXNrEfPy6BfmMtQ2OjMc3cxjmCXrrQHOFvtCSdW+SMwfnMq7Q2rTK1QY
qW0xCrspWjIPXYweLKq2YJt8s5lGbpHOLedYpglQKXvLn3LGp/hiu+o9sI2ZihBT
LoTbh0HNN+XZ04mQcx+BrQFhTgIPcgDl7OqUcwP2wBrE3pVbWtnD8Sz1lKqSQdQW
GXAE+C3/CO4zuvMKGsNvHwjpVWHHGsSRZWhkgROtEBL4WGufr2UrXioopFjshplq
WV1kRJRW3bb/37zIf3aWZoCsLkOv7SQg/zJlPvC4hpwt1Dlxn6IzTHvUsthXkklC
6zya3kFsY7GSvWm0+UldjHqNpyHtsuDhc0cStxFRnmssAC4kjiNRRMtKm1IW332H
6/gqvNihh5YkCAtcGGEJEy5YaY22xLfQN+HBYXgfyomScbbWQS8xpxTAnxGANWJd
o29FUyEkb89ZUgFjrl0vhpbGv5SqPhqShNcwkWDGJexLac2i8yOLEsP7F8wqHdmt
jkA1EaNGkXB18KLuxk3sAlKrOW0QVNkweLFqFoxCTMZ+y+N3Rui9NNofzREOJ7gj
`protect END_PROTECTED
