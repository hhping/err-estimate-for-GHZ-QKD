`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Znvw4d5B14KhPLSqhwOZwFn5JOly2wnmggB2VAGz4UGKziHcW/CFgShTGkq6gDwp
q5VVPXZBBiKa8UlyWnXNvvyRikD9xREqVs0mxQPyV9OsP6tqwEgcOlcdC5V6qTcL
01XoLH77CyYdzTVv7UxXuee8Ia0+Iey+8Y91C8ZnmtC//DKr+uJZ8lLB6e55AGUg
xDOl05GuNDSk3V3URUhsSuPzj/N3FLxlXTTQUATXl/KO6DXKc9LfvK158FrNacZN
qnJA0vqvsB12JLyn7svZ7OCTtbsarreLyDx79TPReqa42H8F3O5WrrLKGAwQh1CL
pL4lcmwyoNuESXonvGyiOehaVVyuQNeKAQfdcAtvmd3rqgnwTtpA1iJTcc4/CmUG
Tj9HlawU7xPkgM8+rjsOHvdczlYnEyejMf34vYGRqLXHFD0ei14pH/+hHGjFeNvP
FbGfFYPnwFzEil1JKO6gBFzTyYIwb6h44WISUDUFnHwkP1wgOnxYMeD3VBQYDFll
wE/uwP257OxqJUn5uHNDR3RU4XxbGD3/LjJ0SfesnIpBgVlXqjj9xUorZ/FI9BHo
ZyZEFIHCofY4QevjOJ6CdpPP5Vkpd6jAkUmgG9zwH4mBJ00wcxgA+Kkv/h6Sdw+h
HV0LKYsnajQfkwN/Lup7WsEftiVcCqm/kqT1fVe6io34F1P2ulTLXFljaJOYqgEc
i0j1rwI2UDCLfoWnPatiH7ONRkdFQ8foBOvZ2Muh2Pjhxo2ONSZ2w5CQN7jAI7UN
+pNetI/IWCyEd1RIipV02L5HW6IqdifRUIzfVZY088EOwTLhnDqwdSyq3Sxq0Fiq
2jN/Rq3m5cQCqt1dNZGKICD7mbdnbhh+CZgxP9LUjrmOd+sbGjgBvyHOQS/RCl0H
398/9cQTf2mGY2T1GHOmxXuLGrQq0VGOnM9OQB5ReZnMAASxjGU4D9QQH+Rre4/u
rIZjeUoX3vikIiMzt5YcpFCwbvNhhXGY44gY4xRDjMRvgpYVRt+obm/LpdWzVzje
DJSbxJCyUAZyF/njQTe8mN5Xf58pOLSFjYCsBmIBMEU=
`protect END_PROTECTED
