`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2Sq+VmQEsCRb0TY8EBEsDZ9POUltT0hHmB3agto4RcWKeB2OrBDs9WF9KHRGknC
AGkh2T8c3ITQCoyOq+seBQkl62JsHVE8M7FZBwRugWT8D5xPECvO0RhIfOsh+QCT
T3xPnc1gk/MGDfEqlIl4qwyZ+ACqa3qECKdAhmWj667U1tM/bgYJcS7JCDCTUZMP
Cxr3u0IBSWRium/KksuAzMFtg2K2ugQC3iwGSKbAPjp59CBdlBW9gDa6viw8elFu
PeZvnhda0XrfxKojGvYdWZPh7NARM8AwI3G5Bc7dPblJ1TrSXukElpdsfg9pKlSb
cbCSXpqanBJFh0WXxko+PEMmiqMSwbhBbpMFbtYr9KWW5qJcLnwxs71MIYfEWyOf
iZJ/WTC1tdGuJaBlMN9ndZn1yw0wAaL1RsQLvKMqxssoc7EiCVIxmbgvLcET3vAK
vi5cJaK3ULJya8L68Tv3cG2+pIGas2Vi8dlO6rshZwOae4l2d3tVeSr3Ar4HYZXr
au0Eu3ypaxWyMRGDyRuZ9OxFhqI8GJEzgz2o09lxgx7Q0eqQ280dihtCar3/r6r1
gafkNMnx6ZizpJRw9Rp4CBavkN9nwkfmrncMJg7JH3gv4iD/tl+QKxw+OwJJVRE2
nf7wqNNqwViGp3A1sxWw+Pe4YofhFLzEXST3tud6xj27XmlECa2xwLov7oitZJ1H
tkP/0iVWNos2bz/SJ7ssQA/B/SqcGLC6w/dBLSK4WfxLnLoQcBKN6wlcrHmw4bl0
7EEYFV0XAnm6QmCwI4m4o52S9W1rxfJRU4+PF5UZ34YwxCH7IxrIIL+OeV9YMJST
rf4PfbKAJANTZlWu8SZrT9UBayXOLiyPflsOHBYjfClE9P9364j1iPLhsU/BgsoW
qMLWh+xrcKCg2dkKH7qdNxs+tiv+zlRWhCz/mRSEuOKkXr+6d37VjiDEVth0s9Xe
TwD8h7rDsb0rj1CyaOLZrZwBe0xC0ZgqOoGbVAWgPzmEJm2LRUIMSqT2+PzQEjML
jByZR3yC+zkoAVrIJytTlun+464onjzdZcKzbAUjeMuE0KPj5w3aqgKutnq/Ua0Z
AtBBpjyjRXfv+PNBGq/NYOtKChLFEiekumzoVNeEHfr7ovb8MXjQGhCtOlhelNRw
7/AIKFQORbpHMwXSCs1+hCJX0eSl/MRg5+HQ9kll6SNdKKQ8q5AvBXgcx+lXuspU
ivPJ6mGt+FpyzXjMoI+RMl72U7TTMqS5pIa1XSuM6chvDqheC+om5oHGPzZ5BZkg
5oUUNApqv8V3/risKFSD+DNGo4Oq2SxROVPW0dKZtO8wX2d/+JSd0x9vbcZiIFYQ
mOEmiDBeS9/IY0ChK3I6OvrNRHUF0A7+CYHLfOPEoE29r7Ic29uD5mfXZXR6Uk2z
w0Y/N2/E9g41CAEYqJYII8DpeG/L9fk360cmQEaj2JVPt3fOQqeGPHH1X8kvi6aa
0e3kRhZPEbdbBOsQjmZ55D+/OoVsE7l+b3k7TURXltJGAfd0T8xI5w5BY8Nyu51R
GM762trLIx557355sIi1pV/iOU6EpZIJmY0lawY0273QQ3frEP++EbjmpSmy+lzD
0ueKZZDGX9zbm44hhzG3TfR53HB0Ath3hAlBG9gmAbuW4Lhmq1oOLCeNCfcQ6/b0
GQACXOi0DmTwIAzKlpMrrwXWQG4Es7zdgJ5/vGdvh9RyiSmWdFDVZ6VuOQkdIqFt
3z5seDtpwyuX+3/7jdRNoUCyjt2TBy9XRHnwSz0JoFoNoIcgTCcS6kwQIAIEcIiA
hsCgQ29amOdI+JcWS3NwbuMQCpgdHFzSgbk7xr6Fi7pjyw1VqQMJGsQwoKihbJfn
FKNNCjfznp1qu6cQf1qoG+JkpVpmhC9uV9eLST3kqhcYgM4QTW40KsFrx2ZM98jy
bLGQIGvYZhRtuPVcogUaI8JY5XSj8XugcZYcQMe5oEt7lKhgBN++TNvOqjP9vIC1
ZJtetJt1ZyitSwgBkoimFi69mUbFJTheex6NB1/cDfe8e4NikoseAsFJbgbGNQcD
kMMoqOUb1+tyyH4aRI6koI1IzkQ60bCaayTS6daJddj/fqGRM8WqHp1OvMt/4+YM
yx2QVzh/44rNn1stOFPGtGoEkz6x/F4bNlO9udaSbeyEPnM+qAXpeRXk9rkqDBUa
bMlDMSoW+QtIUsv/Jz480wtkL8uan5dlMAKkGRmSsSKsS64hxMrwlZrfLNyAPvm4
XlHwTrUgEx/lY5cuT8rq4Ay7WQY3Vxd+jSXN5Ap0cD2vd3IVR2pDlO0Sa0AsVsNS
dnTIt7x7tovMxuNtRPJMg1zSYOtwkJShYnptitHmtHdQrn8dDVFLIfktlWUdd1RX
33jHhnHTD77n1uRddd14Jo11u/oFNaQV8ZaypxeEwhWGQ2vlrkt1EAv7/sOW+A8b
sFP1GEIzQLTrjK8jlk+tEwvnBepmMo/6CqdngJS4oi9abqd9IvCjDUEmAN66+g7u
7CVNbSQI/p6MAKgqQe+5lLJiX0CFtoCpzLkatQa1XnVrpROQMJUPoqsk39JwK8cV
mZU7W0cNeFglzZ0OqGlL7xHJOjXWqM2p696HjcpuOCyfF9DW2uOwqdaviDBEgOdQ
/JDw1jMFwxiPcHKgdOK7rgqK5Ww4IgF4DDaG3b59a0sGJ7xlrFcPJkHacpUuJw6U
QNWjU6GAK1J2fDL566lWFe/RvHW4v1UK9L2gL9sDLdJhml/8BCqIAkr4SZwj7ddW
y35or6UchWlWMQSyqXeIqsM7vdIQ422vAVDFv0MHUycw2QR58ETRT0Hat8RhTen2
OZzNvHJayn1yE4RxehFE/kPTeESulFTJyzVr82VcAUt7B/KVd2P1p0opi3XDEOfq
yRZ1trAIMaoZJguurx1ZmuV0r91AV3LpNgGZKwNAo6p+ylkIDML4GMjzdoFPbbhs
LqYG4nvwG0eRk9OPV+fx9GE+CgvNdXYzNKnPDJ6V4RP3Iq8YP3Od15dhTE0VNERf
dZc/DQbkDJsOztZ1j/ePWsqBgx8PDObKkhJPzQSFZJjwMfcGnnPPZBV7vbqELViA
oo2+quzR7n0WScPJHVgrnbo9/hH0qKVh72Iag2vzCjPBgQOS2buK18zF8CBcidWN
EZo04ZmF7S4XaTE915cdCuAgBRPaGwl6wjmJI7gB/r50eo2qKhDJ9xkw8MQ3GswM
F+bkyltM4uGGlcGO1N7BBdOpQIxFJdVAlFIxjQ7qdxrr/OtRellgOrTQr0dqtkuj
coC5LWPe1loqR1Trj+XjwUlrHZKhUEzQB6TG4G7F8/KGu0fW5HY61iazrc/FTt0M
ZtRKX68cN53CQZSppQoaPQVgr1bAWPMAghfXqzDeLL+bEqGGEM8nazCQ89KJ3eFH
FEc3KgFL2aALTjWR8Pm8fNUNShkfkN+MKtloRZyeX7L54AuyfbJ6FNs07IiTdveQ
zwhliB0zzFTB4/IpNMUFrUquh2C05VoYwUcgLG9PeWeTK/jfkNZ1VFfJkiX/K/mz
e516pvaoTlAZLsOvlcFeiFybDFZO0OTtQlBQeZSbPsqqhsrlhDA539vFPYxBjzm/
9EGgvgXZ2yyw23BS2UGRl1OclN+B96XJyFqwoQor98+POGW79s6ZkKjlsiZ+TRZ6
TN8r8dE97Bg3KKDOaRfudKbSm5Ksld8hMI1R7XlOc5CaF/m+03FUt+ORVzoHRApN
wLsG2N6Su6ORsEcMu7J9H4SYqBGn7M15IpquDTwdrMNzKU1I/S/UDmfTzF8m7swo
gT5zkCSkzPiP0jp6EhfNiTCK2/Krbb0MewVARtwjUlqBakRcLFCvzKccI75fw/O/
T4Jt2azY2wKsPY6JAI/6O628UaVK/03L4vQ72rImnJJDRtkYt491IKQH2cw23JDr
d2u2FlX/SyEi2eMWpUxPUc2oGv1nbhAj465pmRDsEVxd3MA/dS92dUtWAdn7sy3V
m13haKYHizkXJY1g78mdYOKOl5ukikuhYjVhWVxB1yBhYA4x6HByPdOxzzG1oIlR
TVLVKBpO4QC5BxeTipdRd4FKCtRRYGIhE2CIAdG70+y5sBohHGHvDU+MjZ/Pr8E4
VaJZq1zrU4rfrT/cC7ApdLis5OOpBxHHBbxIUF1L0e0B+eBh+ijBtZHroS8kcr2/
HINde63MzI2+GfsouV2aj9UEO0OVEETxYUNrQT3ebaPHiZEateNPqsRv6rfRzfnS
lSD3+thggtKABYRSpjSQQUTSqOZMsb54ZD5/Ik+WpjAG2BRa8kMjDe8XdvKX54FR
zna3UBbq0ofx4CiWZZ/IqgpY7ltY+pxWb4/fe4uaHCdh4HuNYpSI9E2FkgK/KhbS
Hq59cbya3C+ajjL779NHjKlKPmN6wvW540UBUDQHU4D/51iqJkRrlPwCh6Jn+s2x
6g3sR4Vi5437YgWK0RPb4sdO/SAzZGy2TFNzCvYrizhM7JOnWfkUI5NgchhvT4u1
vEvZr11Jbb1u8kqZmDebP830/Gqs714Pjh+WI5oDBjTaLWEUsERj1gh7B9g/D7AN
gohrDPRjWsEXK3xQuzjI7NxaIdvnmDnghGqPPbTs85HQjlmTRNwSYZHokdx5kjd0
Jjl3FV/hEYils7SqfrNIhDEbXPY89NH+C/m7SlS/ivnjN0oY+NKDHxHa9G0bOzPC
CcYAgD/bamM9z5qwSTa9sheotMBlXISRhb32fWdtTP5/WLOp7qXPEWPslporQgjW
cX2ansKx3gScUHuUOR9AIRSgtSLFbTuDtEcxZn4WgewlgYL0oCaOzuw+L/HwNxja
CVxZOCoJcK1nH2OVEnNOB0FFBPySiYppsFpazlJsv2yAFgXLrHkP89lYdyTGH1ZU
hGAWCrEXgD9pZ+vsQvCMpe+n/Pc3oVS0u6gYTOjCPKwzh1sj23uUqcqwCZhyKsOP
wgbFrgFIg9w3sy3oLtvyS1nf9hMR7YRdn5WixMJsKRGuWDIQhjAZj+ss2OLixh5h
y6g9d5Pu6JDcatdmOfYzx1A6CQLqUXkw27zqqPJOWyF2v9wGqgEkkq4rZh5hhBrV
GnlMANBoVztMPxdxEUyrMfZHV8t04faYZHJ29b6LAGtbQ1b+5Pzttvad+N6+MWdA
CWykicKu+gNQYB5AJJpRh1AIZIu8lJbhXx81VWJ5BKWFQ4eZMUPi9I8QzNFmGkoV
0L7RXQ3V8GxRAI2kSYlHBPM7BzB7y5Y93ZAfHLiglW35QtPNZ24abR2pdTI/dV6z
7NquCqjZC7McJPFRwK406cjrVVdYRclaHhRU+LnpHoihqR0/arwinNUmdoDvm4ow
d76SBd53b5sK/KCvboX2+i1z95QpE90xoF7P4Uuq6xz2oMxuxMU8NtYc2fp8cJN+
r5yeLlEAuzWxpW18ijJlcm9U/2DTO44l774+ZVe82GBNjnpqn8OiO5IqGZf8BoeA
MxNWYHWbbSeP2d61gkH03yGkNctcn7a3KIiopS/QiBm134fTr5A3ur1mbez6PvIv
TeQN/De+CbyPlmCVlKS53ZMODFxOXSCCJKkm78hYkyw2GLHgXjd+GZAgHiM5lg76
2bctdOoWzR1bFKuhHOT7xCLBclA/bti+YTyXAoD4g7ErPgwDKn/dOTxhrGGU7BR6
Xee4AxtRez3JCFBo3ncoDhBZzYjzWwkamxgB6ij9R9U2G8LhsdyVcNRneWav6n4a
4DXxdMhZkrVVtmTcpI0CHcGbU3UlvJZZkaY3S1qdb44ghD/Sf0ytNGLkeasv4Gz8
epoNF6wg5hQE45fFnCRypfTcj5lm14QlnCW2WSCgTTGSPzRtPF0wzcOYJJ35g7NK
u4+B+0/0nW4ePYaOtMZQ5yCKl6+vtMdZr9lTf4F//xg48DanTnVC4CnuZ624zSOz
LxWZHVPBFxNLhDtJbV2XrTWRZ6eUOS66QoU+KjW3H2IVfCdWQ71FKrgqGudOTVPD
WNwSbKFgBquCmeVbzOAnJK63/GJfmtqwp4LoUEOKzKvcn8Yh8T+BuNPSTrznIhak
4B2kh2Zk63bzsBaUHW3I12OHTvHHnaStWJfCtyykV2KfTccsXTJod0vy3+fm8tm3
KA/KzvW4D8483E6GmwUb1aPRbuK0YU55X3+WqX8TxDLl97L0aZunyk8kVOotT9nh
XvCE+99y6rgOLg7sgFHDmZh6l6+xD8VqHS2JUuaxPHgWGFTK3jF7blrMnJYsO3z7
M6rVXSfMw2ZTzFNK1DDLiKY19XZ4EMhftOYG5qP3cS/XtmfdHHBxbj9xJS7RN5Af
eMGPirqzS8wEFaVExi7aHbxirNbHU+rp+ypKCOkaXa9vZMLAfU/h6lqgLWAqJDOH
E5fbIfNhqmUiFFn5OHNuLoHWqrh8fYBwtpIRVA1+G5O310qDL31ldZnv/BJKwn0Y
06iHZhMM89eSmAGRlcQhy81XQxBXvzLtJ/T5KAXnhfChGJjfSApqEd4K/WnepoR4
8NACENJOs6OiOHLD9Rd66OEFqINco1f27ozwMIPoj0K/xmAUmmyOJHEanLelsXGE
/K+aQ0pA3gkkVCnC/q9mRM/FRsyJpfM69/OLC4Ipk/pBNhsVgf7FBZQ1oMV33/CR
uhlWeQJ69HwDt71qYdinwkoCYGn1NuSxW4gDat/7XvD7CIq2JJRkDS6Uc/Lqx9Nd
WshkMCrALTQXncNRFz4PG2J/FeTItczkPFfW7R3rhOYy6lciNDXvR25WJE0mnIqj
C7zpg8RlLAaASMeV1xGlmljzplYkDjzUaPE7/GrDlFhKv4jy2Ij8NYoNqubNtfHy
+YJC1kEHJ70mjAFN9e29N+ypl/pZGX6nCKf4J1plCw6SUURbCp7sddFHbbUDT0NB
QmzyoEHnMvxB2VtwuxPa750bxZp5toN1udWvnSdjhO2q7WIBaRKKz9TeAUh5yRuc
1WFqWf52swSpp5HD5NDTAyV3UB59rlNJbkFX9LSqB3sh3taJrBw/3O+pfyOfiFXy
Tx0Gq6uJL1lR8gg7FVbwwWuFfwwJ+9uY3Zwlpz42zk6EFTqZ26KlmWt9JIE/Ys2w
sLZJ+kw9F6JyTVBtIKfo/Xxd1/3koKeNoe9zz7k/+GMP0W3pvgPJWQqp4/kesDp/
9EmjAA+XECgi4/ThY0kSh4Y76Ec1KkIufH2/63hrncLZ+SUtUEhY9Fe6rsw6IwDP
g4zidjmgowK6BDKzQV7ZVpLe4Zgf8E60EaaHkXJDaoOcJaaf8koH+spOqBINlRVA
i3eRSmE/9FRY/OKSDHWg0IS1W3hevOEfcy94lImCESPYzf7DrbBZ71yuBRdQzQ46
UzM7cwtruMHMy9y3l3JGUqtTFz5pQWgywcXWnWzNqRyDTLTVwQKihyCwWM136GTt
zCjjuPDqeXdqo9UEFIkCPYu/orKbib3z6nu1U7OCNDQbFvFJYL0768p2/b9U/pFq
gb70V6gMXWcJ5Y2oCEjDmjoNqkJQVTcFZ0/CtQdLQ+fDDPFNw2OjnBnbY8ZVD14u
Kg5TqCWQA+g3x9x8NO1WGz96Mnlx/HrFUPXYgzJ/zal12a5WBPvWdVItCFO3Smia
zQodnHlX9KUe54odOmZWmsh/fNajU65113OtMMwhfa6meYa0xlSiC0NMh2H4GdSz
wj5JfHtUpW+yOhzA00gPskfhvgwCEupllj9ZucZsic98Wg+ZzOsnPCYpXgC60uy5
tL4GEjSEk1qm9KImV6h5PSrJCnHjQT+5MSX0uQPKZnsSYUzZOSZEqkBPll+L8osr
SnS/QlXiEMdhcmZYTtaxmf9rGm2K/7XKsl9Y6QorQVmrbbsHlIz+GNlVr6rrUvdq
2ed7Q4riUb8AdpQEJ4uFnOaKyHkeYUZNQ9eA+YUSdrVucod+XBGSDcrwJi3i8Jau
Z+UP2zWL0EMfF8yQ8x362ucDvQHAMXSa+2/9PrWfmMlIXu6SWhaXq3HcWNYSr6+o
RW7ZvbR3xSvBBe+l1+BDYhrPYqWRt2wyxO32vy41VokMq3HmUMoYDCJ/o98LYB0y
xLXr+NZdvTS4OyDoisXkDs22oImb7/5QRmQ5YVSwGhRalOFeSNNxj5bIB5p4ZvUZ
iaMdiMx9KfLlpwXE+FhcRMQMnYdcUmbiGxjh+wHwPnk3X6h2hcI6usm/7TBZRg29
vxZk5vXSPPLPBVXKJls2tszRRVXxOQPG5UXi6ZzPBU6UvLx8aCCSO3pP1fsonJIZ
5fKMS07ZrHZwumSDgLl9YRCdzaELC4dap133WnVRnJ+MksiG43STVp178vu8NVKi
ZA8WvXiD9xP+unItDfBxFANppPicXQzA2dLbhU3hkL9pwLxiblBmMMZxS7WMVe2p
2y+zSMYm2qN7Q6ZxJpRN7kYD2d7HcPqoneYKLI6jFS6/e71wYvhm2+lo72zbFxNC
KrzJmxclPZsBpdqWV2znXU2rN33W41HDjjZhPl7tucMvirRodfHRsnHcCHuWjIXR
w2p8xbCKqgqc+u8u38zrIF7fhe4jR9sBKlEUHWbeUJB0l0qRgnvHKXQnde0Z4NLo
Ij6m0L8A+4MNNe2IsmA8J3EP0DWyz6XUAc1c4aRup9GGV/V8jmDPbH5Rvux9FKYv
6kQgxHKc9w8ra5JKH7Gzke0UCJtfZYKVc/lldPGd/dUjQ9dy9xyBKWfubmvCN6+T
HzzaKKC0sJ3ns8BXzwBp6ROdPisJLEC/N9FkSRK/8adHBwouzglcXK1BDDoL6UPd
4vfCP7aiq/0vIxJp3LWV/4BvgATGUfAsiue8iuZnimp2grl6Y76FDeFncqY5EAF4
eegTUlP8SP+O7aeOXup/OZ2CsSNk/nff0E6IiNac0fl24IUK+3kI+dhZjE9H/cpK
6645bww79TuAKbJysILdP+DyavFtM1RGsjqqtoKaHQtMOk14CVqStdWUCSJ4JT1E
ncaJuxzyJvFtXfbp1Wk4KkqA+/oUu0tbXIY8n9IuCcQnBaY8g2e0LRroxKk+MM6Z
7P85Cs1x6CpOitLIO/1ZsQvBeNAs65dqCbYC5+sA1gPVuzVibN2YXQY8KnKDWfUF
vVFHEGFLNEUUe2Bq5Dzc+QcMDb9gv+JoW6bms5eU7UeGLB5xvIFHeLERFOA+rBw0
lyryy4xAzGAq4bjzeTcm1AT4bSUOAAKFRtomcKi+EL/MG19gIC4vwwMaNuh/pwPR
DAeHNIZkBT1PjeRxvSRl4Bgvigfhg6Ie8iwu6x/g7KlJrYJkY2LFqKj2gr3FxO/1
n9K4ck3T6T1Cu7dnO2wNQyrdmPZnPvKxBjjs+YJ2FCYXmEKf3Us+2x1GTUgaJFuz
Ns1qWc7JB/sfMJegIIf+1bIEQvcTcp04/cMugQmRGsJqWFElKQB5RV3s4JQxQDbI
1z0UmINtwK674dhBD1ux12vLYnMjdbtQOzBbnaioLsrDPKHax7xwXOkqw/sNjXLN
fgu+5ogYRG10QXn6RUmeBxo9fJiT8uhh0HLKQe+G9efcstJqRL6blqXwHRu6N6lA
LewMUellc5G2EsK6mMivnfSFmhX/djCIXOWyxxJN/zedoyZWTUxUI+DNv6y2PqX2
Y6G3ODKLprYxRibbTDJNBHC/jYESo1dqfHUw6A7LSTjze0zpO61j+Qzo8EO2qhjl
T0xfRXe2n70+udRC3GZ/0lnPKZMSdGm2wSK9mbhV6Cl3bzwQlfgvjLmYz/hsGa69
tq3iO2Vyph1Tx8Vhn9txGzfgSkyPiLOLd8OCNwvbT/WFs0plG10rocoh8dWzxA8h
LMRX/eaeRq+SmnT0098Xsn6vixumC+iIRotcMY/PR1LNUd0demehBKwwV+xKaLnY
edtz61XCmb29YERALd8jJE+KH4NWYo0Kuq3p2zFtpB4wEUNpNrEmGp4o9woE5ib0
eOPZhRhT+IO+twRX570bkQqXtrcRU+iuGIhuGaX39u7J1Z7ZDGvFLgL2XJ8/htUD
lgHvKsAXdRdP8mP/W9cjNxCsqXaHHmQMp2UkVq+UHBsFwfWpTxGTFuyDPpF2RbJ1
+7EjrXr8kK1yPp0kaVdB9Azr7+IUBAeMPqIP7gu/8PeRr86JeFTJuvla1Zec4XCW
RhwO0qCoEJ94APygRQ3Tv02ON8zl6E+QbzWL9b8igQQ8QbXay6xBYS58eGpqi9aY
DvNyTTvbx0fJWmnQg9dwnLboWWJ9YRjCGbXR4lHiKqyLkRUHzvUNM0dDI8HAuxxz
0iwMtE6+79q/0eoI3XMbDFvi2Ijn+VxZVK0fgMzVk6BoGegfMzevF20viihvKDu7
ReMx1Qji7OwynsMrIyKjBHmjWaRseqMiFmYnkrZKMO6pTzIwvPFktUTn8BkTeCLM
qJ3FtAk5mu+HdZjkz3wxwh4N7ZNOOwYVVAMp8/Py+98I8ABx6AXLGUxHqpNenH84
2/Mik7uXxAPd7o7uV3f8heaq9h+S25tlExPHzc7ywMFyDtwvkcBqFpby9rLOp296
Dy5p9f3EtFbgGLhXUiX+kWCPRQW8Wl9sW9spxjY45Shp8FQmPAxva0n/nvy8LMku
oygEa+WtyM9rkt7tzAjNLtotNOvIzWVKuK5mXK+tNYR0QWncCSBkh1j3YQIt+wAk
TKKU/DmF8FJvpDnUHjZlBkEWwKd+MgTZnVCP/5jvL6AYCJWK05UpXZa3bQ42SfGs
r/HH5hFKhUOlqZr5XKO2eUJFUDIR6GcijlW2WT4FeJxnV+ucKBYRP98uV8rJe+yE
C1vPiRQcp7KOkqmoO5HSv1/R4ZCtTwyzp9k1FaYqIAe9GDx+sdaOAjvISHrrnbo2
z5M8Nx0k5vLGWOl1ZpZEpTBXJ4Zf3MX1cY/zIO96KkJRbenclClau7W+5ssOFJgn
eTDu/z4AYdv4XWXV8AEFyM7nfpK9Jqmkkv+zSOFNHBe3y/uSdHdvIMatGcAnoklT
waKmdTk+9p86udRLNZ/JP8UUBidky2ax1GoPkuT2Bt5MjnfxDV0BCo5AQEu7XK4r
EcLF9IcX3VUuVTAcqthlr2GYNZOGElcGNBjaDJelOZnZ8HlFAr7e0KrxyVPthh5N
ETVDgy7HssIOgvAAaEmcAbsg0rwmZl1CmngDI5k/VRHwDcbMM00RzWJ/qY98rIQJ
5Ut8e38xUWIuZNXIAWb3+DnNYXB8tLdbScKfuEIBqmM0KOpGAJsVkssqPx3vmEJf
ZPvF2jERh5SLyiZSztCv0IMFSjcs2Bz2LPt7mOrPnI0rSgr4BMzbptWTaiuZn7Ow
ZmznemMexkIuA71fJbeKguVjI5RJBL7aRei3BvagkD/UVxr8Xa6hKrXE3qJQCD68
o2kwuRenzF3xZr0o5MluDiNjDus4/uykg3ZT6knSLZ+zYJRiw8LRc34beAQ+CcLW
f8g1EGHIKsDseOLK5spzgmX64xq8NFFBKrHT2SNuUlVVnKe6V6SIV9wehpDSr1Wp
IF6Tir/FxhP41kaSnMc54vyIb5d5qR3aDhF6BTkX77QSAbPdHTbmSprvSyHqfbkR
tqKUDf4pJae0zKzWBXs6mxDWJHFWkcC/s9Qt+WaUJGxsF5SZH12TDc1Sozed1N89
2FcenWOW030dv4LPM2LH6yat0nOHQuG+W7Uk7Ee1sFQEMcFukcNnDkbfNt8a60eR
jQ5tVkJh7y10ZjjgtOHHFYt6F5hs0KtE6Le5Ccd+kO6XNx180QQGYZ0cDe5uD2wg
2MfanO1HPaW33KpLJNe1buY2YLAkIsyOSkIEpfrUcgpzzy8b/bMO2YgtsZ597iii
AEipl9LEqNgT7g9phC8pnqiqNAti5IYq33fCQDwD2li7jP+JroDhUVAP5C+7L+aN
PXAsDKl96/0MNGjpq/KuoDxHGaMnnxEngvNYPnNPEausGw51N3DpcW8hfYT/SWPg
KmOrNdZ8X1KxiC/aLYINzHZcSYMo3ZEbIy/dFiulCo3V3sNMVdDRPwjc4qBIVFi6
nE3WBPZ37weh2SyeSUBABvMUk5W9u/oQJzHh0Qb2aRrviNe0MIbW4d4JxFknpYmi
5lF1Ill8sX4FwR1C/fNGXd70C3ihRaFrdEy8dMCY0uiLEpFsJT+0cYjc1ADjA7yU
N1bdAc3E2TbsGt1oxgFiGiK94B2/uLHVGARsHmZWIdt7bVDypDbDh59F3IjgEaGq
Fs/53jpyMTIDaxi1s17Vpsu9sLtJL6aum7KP66iwdQXxTtYcw4sjWpQdUp/F9tb5
8w2YjgnvgPAkla8mieUEED57789t893R/7c3UUFg+KxfqXkLB0k/0SdGAriQb1O+
0bbrAf460FqMRzek+N8RtmZPqxHsGRyVa3e25B9WNWCsRRew/C3+ZFnCGHwqe4sD
sYYAEFctyfC/OUw1cApJLjC1ycSDBRqoLQq1JVv4Sw6gV45lugpIoY8y5smOKDGT
ueWDuCgPbszqW+PyTrqRu5ZoNGaQhQz7LwFLuUnn09fq1dBwQngsZo0s75q8nYG7
irMApInAbgo4oWuqD++yiRnVf2YgOCc6oCTauZ/4qMmhZZvSEKcVMo4awwOOC/8Z
fe83foIZmNPmkhDfFbFfEqQM+CM0fFrcugzRN4lw7MeoO+KurD1gft2+YJ+JlmDC
Unb3CUla6uYDCve2yVGduzkrhddgk/p6iOj23rKnbC6d825Th4wHkMaFibjzo9+X
hqU/adGQh8KrLjCOLKO+SzTVuegaypzOcp3jDgy2GpjMLolt+tkt7XXj8FDM92ON
rKG129+wNBlpuJMKZBXQWHG9tseWl53mpMXIYhfKyvhZAPHsnjzplhoOUBANKpyF
QVlghyc6q9vT/oaNQ9FKD2kdgGBUqeGHFwCJrnrayKs8VP+hArZW0bnNBZ/mEbrZ
O9RCQmN9tuHTUFt+cfr2pUJzKcIZDEnVamUgQ18X2UU6XGOksSkHCN78LPXiBgv6
6isFzR8QVd1mIlQOm1EUVBaLrHW1wEDi8/GKZUtx775GXMm4gu3x4/9y/svZsKDd
KPd92kGcWBKHU4U6x5CAO0B35oPNtxcwux7wAjAUZ2Ul5KTsQk2Pqr2Dh4RXG5BC
AB+788HuyKo0i7ltOJb+SavuAb264DzuF92XIb3gQXTL3fvbB5g7Uagtnl9/LcXj
mbuc33li+FQ74mmrJQfAkRE+NmMT2aLGe6eWXzuCI9+/HzB4Imx+Wnt+vx29bEyB
9iWmucnAlP8VR2JmiKOLe6xGEBGn6eZKtAfHGcs2fl4s1zAUCH+onYG8gJrbpMzC
hrPWvCVt8AzDp1X6gJT1KeMhbw32qfTytwqiCIa8cToujWOOP071/H27pqBV1GXp
Ekf3nyX7zoQqRDQ1C9AfPtVh1o/A1nl/EqSdI0QliIwdRbZQdSW6HxSIrk5uND7k
1H0utydeZPEeirAThB+WM5sgtY6Be3y1Jfp3yK3Ps4IqyexxQvZoZGhE1mDWWQrY
3juFVzezIYdOfLAQ+KaFdiVv5Y8odaIXwd//YQTAsRKPmngMhL3MB6w8uNLSUheh
fC8Jm6YfKsiWEk3DU/BJQli0XEo5JWp93+Km8sQm/ejKvxKXJ06q26yfouPFCekR
8u27fNKsPJkOm9wm6mj1IyNBF/gyeRdBkjucOdM19lBqCMEP7ZXAcgV03ME7q9jQ
sYH2eMOkWiwM/WDWtKCNhDsC/KPRDkofbhQD7le/eroo83BnIBQJEVmsqC3pznQY
4e6LNNqm5AhRaRwKg5QI4InFE122oyirCNgVyD6AwgWD4O41YUS2ZftRJBg2XYoR
/hGU8ucDTP4ewpoT+bPYXx7VOfM/dbziXrigvtR7bk2axJhVn7KqOeiNr4f8VITr
4wpPSYSw4XlzXNTRiGRWGagfNFdytoqs+PnyRCG4uoJqdYll0FAjDuM/xyFB87rh
l187yYpfrZNqiaDtZcgqHdRDOd/xx3XRW4nxtO1Iwd6pi6n1xoYl8cZ0Mbfz98uG
XBAThdm7ejqX54ChZqgKu+/DMhto+n0xRxp5U2l6XjJOAQBQE6ezINiGOrpHwIsm
5Z4Kd2J+dogK25Ml9qJtq8YnUO3kuNOKFdx6ZGXeOM57bTROqVqqLh7RMuRR5WeB
fS/5U+J4p80SF4vyBPqplVJCxsiQg1njwlV5sbGQ0XLbe463B4dkrsqDUXcMiHrC
mRJNaDEi9IESMUqe9MSyNDLg9a0V1JZLj9NteeC3/ewAR/X0KuA8Rn2YK8axNgHI
NOXx85Cs5V4CftfClm65eRKZJ0T9xDtGSnRscjiOEcqrIa81H9NKBBHBcKpbcWVg
Ezir+A9FR0PacQMmFjz8ItNdKNNgFDic0uMQcL/kZYHcl137IAgm3bY+bygMZqBn
kTxh/dOy3NaqCyIfYd7Nrdtq3XEdfMnbjNrmnJn4U5p7wA8A66eK0TyYdhe7icHg
omRHht5NfsK2fpzxYgtRiH5mnoBFgHKfMukV3gazW6yAbHWGjaRkOS1RcHstIBUg
djXdqUipXpcH0Acb/QyHHyKx0138oltd1NTE2D9V8JYH+f5xN5lC86dNSvoiBOwT
RU0dRGjws37G6UhCjYVCDItXoxwfEXXoI8vKIUxH9NWbp0XugialzC/+oSqF7Db/
lnmXdsU2x93/nYuQYmE3sAc5i01d+im4nZTAoFfED2mYss+AWBezWwE3RsvdktoL
z2S8OsxYqYJntrmTsdVamUj/7BsW3jDHzo+fVl0hV6aSCTzQUHyIESwMSBlOsXJj
fpNSEoKC3UATG17KfHEGONSGUnuLTVMQW+kQjbKycFfN+1OjI/dZCflkZGTYmuj3
iG7pjcbCPvWVt9y5qPjeLJpTcNFkueHjZV8fZ/t/4QEC6WBwOLWYzf/m0y99TRpA
ymO4oozkzKP9sLQxGmgRRaqfFFIt9agDLEyoYt2vJxtfO1n/A8y9zD4CV4uj6dyg
XJP0SgOrdZz8Rl2pqaYbvKCgxQBCqwDzUn8vGOoAfAEk1rzntCkBobZtpjNUg0yN
IaB1WCGJnynkoCKvMRmv8lPCstOKKR7q1I0oaf1c/Xm/l7C7+m+ain+EPov/yn4R
OwOXq8YOQBLOsUpT/CZjlb35Ei9looV/GWJ4X6UKEUb20RTK6K60cvR9XaAfkmy0
sqSQW45y/gjgiG3nnpoB5+wvtMME37eZAjBQ/rgImpb6RCgOJFVj+nnsguMmVzYJ
4VwPGaa9nfE547ybMed7izBWnydkP0K838Oa0AB+pnEuKeRM9dlzwk091flBVuxa
ejj/C3qxyPM7Sv/ojCkEQY8o1XmKZOFXyb/4jSEnPAvC8TWTWnqwWz446q8k1cRE
LXEFnycP0kxo8hCUyNKcRvT46WziUBiv+nFl2RaMO0a8gvDvF2EsooOLLULcxSCA
nnBbD2adHFCXtw/39JKfGrTH8J7fsOexkk8etbmhYC+/C7dlZDltH8zo4I1i0oL+
/j4DDJLyMkaFp3/Rnr60Cx0e+/m8TEvM7qakOMKrJsUzbunXusJQ802zarOV4R7I
pIVkSekKjcXUprc1gzumOVzVkfAbZLxHvp7UAFpYTyOQA407RYpOqNFanYvI1ZJ5
MSGozwMy3xJGrAQj5Qw9qzftM5L0lnavvsajFplTpP+nEBe0mHPS0c7dUXFwGMg8
RbnhrlAxXJKqG4GT0FUt7g==
`protect END_PROTECTED
