`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R3KOjX15HEoqx7PNu81OiL0mLs6t7N1o8g5fVN8zzYtveXPZoH/e+ZabhK63RxR/
BqdqacaYXVhprQMOd/7z0fPDquWIi7QY6nSkKy4o3OpRgbAw4glgIzpCKjPWfll2
Pzh4pVbCe5df5v5lvE12epR6sicq7z/St2p3z6hGC8O8r15TvEq3ZYfGTL9ChP6F
sCW1VyQkS76rZb4BDYV8SKlT3K0BYnTx4FzOk6TRcpIV+Duiqx7GYxSYD6H0Rbjp
pO2Fm2GG4t8j/y1WtuYRyZ8naDf4t3b7YU4MN6xadYLKQoEDBzlJFng5TZYr2rbp
/gjpy3iZe5nxmA1fSWqWX7+9TpyAoV2aHJx0rJ+IXskHIfqkgGPAhpjw3brOYdwP
6l4PrZHCK6Eb8esXV0drTkjJ5c2XEmW3IvgAWuj28KU/1wVw9joMc5le93HA1ktZ
8mfeU3iQCm1Gi3S3KakoQ18xCy8srNG9mac0of73aOTpUnoRN/aTYbFlYO9ZcvE6
a91LFGmSbhUzo7fJLmdqZA6XVBd1nYiRTC6VSoB5iSv1U0M6skgToPMOa/KgGzIX
oU8yLyraadPc+KxajRGPtn2231uXsITj4sZ65wMjn/2FiFgIoc3x1S1WRM7HsfKb
cF9fs0kIhIBBID+tXj8YEm/THkB/fZj/5QME/Us+ilV57QnDX+RhjN6ipPdvoTP9
idCpNfAmF4Fxp6GnQuwlAZg+EDxcENzDGtR5AgeCTRM7TS/e/kWkx/8oZvwdlLgn
TJ2cx7S7RsxdTfHlZ0TSR032cWlnlKqyvqAQGmpxyOQ/Oxi4FuL/OIK65WYZc976
6LeiUBfTKtqgaBTpxdIvUpZlCvV041RTVSnBKnIjrc7KksjmY3RB3prkDANLUAWD
SYDcQTm5z6e+Tt/aTPT5dDV9ApThOukNcBOvrXyRDjYzYhWLNRcezhfHD5KnU1/M
yPsH56bTe5COyxe2+k4u4AUlMPiA6sN7/JdqY8ojTgq3FsUlCtcjLMJ1jmxHS1WR
MVs40/GQtSohnr1EIFI8srkWcxbrTDEGnTSZEQjrgOZK4DmAPsJusST9uxQCzD0V
yZOVlvbeDQcxtNoawJBULnpxfTaoS/tHilG8OWN5hVIohl/JaakXX/E+paX/IzLh
iC452ip7h8t1EsJTo46TVxFXd1CLxkreTFLfuR8cRdRNDyppAr9faWKU3FqLQMMC
KRkVnn3pvqnDXBQpiD+P/1JPO2+7tR5EGxjpnAOgWmLJEBDldxUxwREh1WR2RCnI
ei2W/eOPFyJn8aukeemUdfZH0iVOJsmZrR81cfaLIcqDn8D224TnPBni79TgCNbx
6Tf5V10V9lgs9uWkn7PgXhumrc5VcPIChD69BUuE9XdON9+AOYYga1iT2nvF99nI
GnBcwc9GCem7o9dlwHB+PnSPfsSDLFdYDchTgf56a3z78cfEu2/JFnqZ5u7TNBCH
2GN6/fWJPdM62mRaBuVDCw4KOU1BN6WJB1L84Ym21DDSml1teusvRQ1zmq1hvOOA
rQXb4JJbKL38XWrpxjbxRHE9VABv+dh0IHq7ua3lirR6b+eR+NJgfb7DUvm4uYfc
Ez6v5dq9jbCl9fsgyVTxIg==
`protect END_PROTECTED
