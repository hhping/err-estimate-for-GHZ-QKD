`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWD4PByUEtYJHtLD3z/PAn80o2kzOD4qELqKnaA33nVQLTUIBcJds/5o7KATCvmD
VP6CEmtTTjeBGACA5RSzGlNa66DZSdDCoQGSTbNu9CTdTz8LJKGfAX/J2AKXOB3u
OBxTHjwzcdnTLhV9lBQXIvQbhVEhkchPFKa26tZVj/SuFG7mnjfc+GSYBgQPqRBS
1f1GKEpm9/qJ9lb0e269LshDCaGVhTBeVtP5iiNkRgXhrB4JIKiy8NgXaUS/YhjC
h7dnM2vq/xW6zws9xh2tn+Vav9GmSzqzR0AKTC3yQQ4DpUIdVBWhu4DjFEaRN5Nm
X2HEBPRj+mBd0vQHYxd+6076B6I5VaIOUfIZs/ErAR0E4hCLYrCoVMKXX9QZ+QqP
tJpLVbYTlo8y3Hlr15muA7/hRyZny+sKjRu/i0v6v0kNBLT3kIlcxOWwQZe1Eqsx
pTEOSg+a3ZY02Qm7V/tXVAD7dmNUTxwXShvCT0u2yUurLO6zsA9XjZTMNAH237SM
tIPem43aGMHKHD+Yse0cBMXEw+76zgcxptQ5IDJdiecYuA4QzWbgQfb/6JSCd6Ot
doz4WHHcN25e1cbwUGqVIffjwp0tOjsUyJcA6+wG4EMhV5lU/qBg9QkZ7aS5eL6i
t6PUXeeWP9Rw7GE3pOzj32Gb0N1EU5+W103/kfHXpowVuoKmibZiMzbfALkds9Lz
shWRC/Taidy93jwNqb94v2r8TGJ5mMq4DjbuAYk+F9dS//D4f1v3CAkfXVrCeU8S
Rzdylk3lr0ntm02OVBxSo+FKS+vQRLEJWw0dqBj3p38gppWCMWE1JNG2jpWj1D8s
xuIR82sOXBzHvxPE4v+dDptO71mhOlLrjec4/vAiahYUMCxEUuBMHR4LLwAgBpgr
KNc4FghwmgrI1FTzgpZ4QxyMrQSygP29aS0ZQ2I8jjlexQK6rZTTEgmZ9uxixczx
jiK68I0pF/6859dsVc9zVRFQxabDYl61nKWb8D1mQHzS43A0iEFWCKTFJKYkDW87
A0TElBcQ0GsBPAbynNCg07nRpEVjrY2hawou7CMlMwhTWLzB3NC+iWHBG5IvJVCz
BKBC2WrIioAfcd2/fGNBzYThhPlANp0cdto3IPiQONQ7hkKzByE64x8M5h7h2hed
hw2hQLtVER7b5hk4+l8z/YjrBUOel39xdI+8HvWhMONE/TwDYjjtXgCGOMuX16Qa
ngHeDaP5WPwHOqqSXdGglmehwwBP3XYEJxXljcryO/AGEy+TJw5U4GSS9GROl1V5
KwFE6kNdf0Ug4plr+LKdXuyVXnQa8LSKDCpMBAtYqgxxz8y6VKFLRDe1SLKyGsFW
lqrwctkPHG9cCFh/yIq38Igf9f/GmhidzpTYnouiyhv/P51QVgqvy3QbM++9+Xlq
GOfjy5+zmNGNgkZBbSuk0pKidX31F13F/39uz9swhtDqTZqTf9+82p7EpHbkrI2T
IujTPOHurVeC5rt2lWjMyvhtWG6iKR1TokEObWBY0vIQIDblQ4pc+JE1e9qFf+UR
wCNF+FQrQ23gb7qwSAIjpGIYNhZlCWl4KSS65+SuSs9I5uBdGWFDVmH3cbqqCqZV
E2BEE8IiqFHp8P3+fe7FkFNk4nZlm6PzIb18AgiImnWtnYTA0yQ9+beVbEJ4pq+5
eDFL322++GadpINjeTBNug==
`protect END_PROTECTED
