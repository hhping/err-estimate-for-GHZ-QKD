`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2LV7J2CJh3Ih+MxxGNY2AeGErIK3zIkcRPaAjIXxg+bV307uDYSaTxX7Yo2ywBe/
ZsVeSML77Nk9sDC4phjWG+yAuTNlupJ2uGdu+z4pLs0kRhQA3XQAuymZnvdry7Ff
EK2ksHlOqtxWF5AnPtjetkSo+K2/xGQb/ncr91E+mEYn+Q7xu8OJSuvsxY2V36PE
0v1zB5xft0QWB2R8nKn3wbivQ7ydytEhh+z43LKcoptN3w4mVw5YQzRMSknqqIcF
+z8lb2GA5gv07L1dv93bKQpvm2kxs+HxQRrOQQFkpeQZjEkRFBJ91AGMsz5V9RPl
acgENH/N891OH6QdiuAABGYIkUZGYQjRt7LU/s0+V4d1uErQ8yuny3yAxDDQRR3J
IBO0e8daHulI8q3/qEf9wd8N2n3EVjGZ0f5kzguaR+9XAbKygGyZzLFEHm1hyM8D
gfFvpdnly73AapUV6YRpPEXdvyHJZL+AwqyH72Ijl2ySMOkBpkAJIqEshhrJKnuf
5UICOv5+7Lghb3s/Whp25fuyyo3dnzpMYmSQSmih/mWO2gf84T86vuNA+Ge5GMJF
jZD2ioUTvJbltzMb9xNg0WJPQoTQ7ZZjQvdyzaazoN8C0sgDhO+Rt4kNYpNOn8wc
/bKb5OKs1S5jkez1TpFdWXeJvSwa/w1hx3aBaNC0f2pMlpY6Pk2Fia2AolEL47+c
i5f3OHc/Vf1oaQ1vxEvY3Vjoi8PXnGpsr6iGzxEbQ1nVBXdg5f+PCkuhJJrr4ZFv
5yh+9xSOWcKmqDZ93xDSPwLOJHdjHoxlA8K1Q5yFFg3WTO1nw/gbbXXP71XIMiXH
d81M8TQ3c3Asf/mFmMpEH4AmXvwrJrZ7q1rEHFrDy/0HSXPT5tlNhXgIqS2h1Bot
YL8oz3CdnkbY8xQo4igjKaOx82C83GCw95NXTnmwYJi7c4G9U7jgSbvw6wwZbNXe
kpFZQ4F9H5HfxTR6Z9Maxs4XKpQCtccULCZnBrsUWv7/RWTLbJ94/0FNYE+wB/Qs
KtfuhxMWzs/bAvIxtw2Qmi0m/SUnXJyMXzdy4HF33NVbLyH7Jtbvye1A0oLgix3v
CSzqBf4F6oXWI1zemO1s7jXh5y0di6CYepVatfl5aKeEqNFXDfPKW126ceF9Uxd1
/H8/FlCE5tyW7pFa2F+egoN06+FB9N7jwzAurPtePomFJDQmscCMps0HK7K+2lVU
twl+Qzhyf/emZu7W2gkhDiqAk36xrZI7i6MqYgVF6mc9m02Fe6tLpD/LooNSP5A3
tLkbxvI16dYfdUNDCKVMargAje8r7c4LFu7GN1TzrP5aDb3YGEQ8vmTg/QYuvpt4
lW5n57mkA/gSop5IvRilof9SJ96vZY3/B00Q5Znb/va3NnVvPQ+YJqXN+RkEJaeY
DLv6nyl4yueBdP1Ooy4kriKKexRGguSJYJnkN0874lnMON+njrvtFmqopxMSItT+
r4/hkE06ipS8PJ1pOAeSr0L8h37p3VJSR+u4MFtgNEAJajWjE324AeRSwztQ12oE
Ah0HQzhEzcUJYWcIfRAghVlfhTLmV4PMLpHLgXyjcK4+lUhtJflRSoxDcDkmdmGB
1CBLneSx1wMwoPGiVFBrYSFaCZ/Rfgv6dMHkEBP8RlriZEOME8suPTdFCdzygEGH
sqPNCRmPrm8yPVBoMoUJAeSq8CHkPnJrSjWFvHnthoOvNekQW71fb6iJM5Rz6E+z
PDq0g+/YPEdmnxAVai1ShT2/VQg4Fa7eE5DIhqvid4DZYe5oBu9sNSLLEh2eXJnN
AxqWfvLMVx0U23nqWTjmHePF13wjr2E+AuAhne8xWaT/MSQnkDaY/1k8EwGWRtCn
UyYnMJB8CgDcCzUR3NrcLG02isFtUT2vB5q7OY/vAM2msMo/I0sxn41hCfltZBO6
n8qe7N6gmpX9KPogJs34DB73qSPHSrwXFeUyT6rjMgNS3AJZ1JV4slVcRgn/ud6Y
3UdtO9mbUAfb3X7tWMo/5nusYlWyCTZlcbpJvgf+NUi9XC6oRnvH0PMcIqZMsoED
y2gLTYa/qREG8cllQvwwM91H3pexas6ItycmZpe2WRGZ84zvbke5ysuEhxoy+jxg
c1sfJjaKi+oQ/JILR6JZ9RIwSYKc2uazCjHKsr+7vv5GTg8O8fxcMcYQCrVW4VZC
WBvZZYeyKG/Q1YuKpJszFX1e7XgZjfM9iCZe7xP/yA1Zp7o5Tn53R8s9dPZkoRX0
wUzxBVbRfa9F+Qeg2/nC5LBshaLUGa5KI9MM0A/WN9zd9vl8hSauEUgxX2zb0Mkr
b3xEVRcOrWkuslzwXzeGJjew6LmkWiWAsWk2Kfu80sVtiToJD+6Gzh2uqcCfrRWW
SV10SKSdSCdcEOtZU9r/sPDgP3paj7N1bHL9MRCG1hJPywtKxZG57YSud3JJBE+k
zlifJBVmJEnwsz/NZRQjBpBEQBDcaJJ/x28bHu6rjqhRa+wmQS0aYH3eq+7h6t9/
9AAsTgmBI51ogyz84vE8fcgYgB2B+burU/QEumDvTeY1zuS4Ukz5CwuOA5h4lWWM
mWTrfrfvxYO0SXRXPxmFj+8JN88/JCepXHg5Uv6Hd43eEUG85IHH5ksyHRnJbrma
59aowyR0j7DdMyRymTZ0rYq3gQck8wsUWXMP+phj9e3AxCPwjq7A4pDIz5axiHi9
Kaur5UUqezsVsA4NmejYxasPknC8hGTOMbRIofyCSWTfouEaXpxguMPd+o09fzaY
XRnWDrd7IYANXRqj8CvGTScp0AtfH4pPvw4aZGmmRSHXZ94CcHbpj4IjZgJFqLdO
AtdK2EDISmbn/wll7kqOZxAk9qHUnjCYh240DZfRFCy0tTQoyUG7el5/5zL+d//i
PIBV9WE9+VI4LGNlXQUKtt9WKBgThQ6Pwcrmruf0ZK6Om259GpiFLV21E8WrkCG2
lZMZ2thrmgA767XywZUbZx7Ks3E4B0WP8tLGrAbvK39+S8lUP74Kkxxobfzvra4F
fzJCGsxKAiwF/p1yGLWd731yT7DrDInu21h8cTBFoxTMnolX/xBIO5I4LfrvEA9R
FZz5G+93K+h0Rjdigh4SL+Ur2+AAZcGYIVMvPafCiZ46DMcmT5/uPgGOyOLIpOYB
/118ugN/S05GKz6gZsOmKzOaYZ5dLj8LI6IFtklfoI9X9n+ZNZZomZUSOcLxUhoN
B2sWCkBDbfQ4RzR8JuVlUqK76ROK9+96VEqdO0kzRUg+qd+Rhu2p0zc3gOyzBqQu
H9GQthPFDwrjzHR0Ek61zhw2K+haWtNKprFtXKmGxGindoLHRZO9P8dDSRE6IxRg
AUQiFfQ02qLVYYWB8fsumB0hsMq5jvE5Jpwyfz9JpUQ0hfWNOVu2K50pVR7bPwz/
ANjZgdnk/l0X/2Sj52csjM67eHsYsPUslCdEDKm3pt/OGJhTXP0NrfTMRmnFZiAU
9soX5QDTM8dka7gGCvsbt/tjXE2wrYuSWXhWU/NjSalR/4Umfy15E5rHn0ouigJn
PE7lXeEUaNeObaLpvS3XK30vg6+BXmueLRDefbAYMvO5b6rrDP6eLv/+wIJ1xFET
Vn4QLufNVOYTgC+9NcZO7c+pffVVWO/eqTk9ttrSX8AojbxcSRRywCX7AM2Wwl7H
G+lI+D1D8SnFABDEfQYru6EgmOnmyoRjK06Zy1zsfeKDogq0lrCj/Jg59LFbXA11
Nl9f/CrVGtDkrUbfUEy7ZIdFEeZHiHl+XiAaddDpN41GUwTaXbjCj2MOUoQs2PVw
bEg9ora/9Iym+rBpOdy0iaOHrEcXkuwE/whqXDqoLpgL+0AmBaNjvUzhXBU7Sllu
Bj1LmRRZOjopEJH9e7NIJEmVuZxZ5pSbDc811gBPmldr3z0mQaPr8QlTbhajrXEE
XDuBcpU3GlDqlFpH4ll2qjvpk1e2D3g7ysB3AE8SKDIBSjlUq4Uul8sp0Qr3J1Uh
oKhGfk7keK3t9Oxt20TL8IDVce2HIlm2wfQ1+Xh2XEbJlxM6GRaoFE5NJBrVm4rT
FPHS2fJLtKs+toFEub7ovIXDwxOeSdaEjJU4QgIYrRB/xEQ6GYtoUDD8mArJqMxZ
OJ4X2fFUIuqEDl0pr5Pdy3PQwJrge3FhzqSo58Te2cow8J7zz483PCATR6/SnzhQ
VoiFwn2/k8sfVQUSz04LlXJhqf93pC7fOGrBT9U3buRZOxeRFBSx27PUSNNmJdZb
1EmHrjgY8LOvp65q+0LmqqLxtxvfDTkrEedUb2Dv0DHL57SXyGQaXc3m3bTi6mxi
rkLNIImBybPf/WT4sw9tfnNgud6yQoNCDqKGv4+yrL5VZoqF9InwWlr9rNTGRphT
bV1cTuLjanl+sBG4+SToz0HHhDmaVfG74vT5xAqueBBEE8vF9l1gVa4XXko2b0t4
YaHMyVzVpwg0fVBAJWU49Thv39pGxOi5GH6RcRIh/tIMAdJGkQSZpW8idubrJoeD
LJpzAZccF3amnAOoiyXBxd04dqlm/vPLsNU6jnLdTEL3wuAARmwdElRTb4qmDkB+
q/izvMDwymBUBNyJFDfgNrWDWmYTyY+qwT9ViKBX6/1HuBS5odUnHzfais4E3HVb
1M6BU7N6jMIhELDPSBArdJ+tWIaeGXEeg+gRuU7HsQQu0a4DZhKRnOhZYBJ7t9M7
7lvmz5z+d2SXFHKM1stLnDXh/vyV+jXtD/+lUx7A57LalqErHBjEUKOXUPYbHvIb
BjZZAGW03ByU+FA2Z7ju5vQeqgwhln1oeNX/cXpmKeq440hBsJdZXmM3APXIwF/0
MEndcTjiu2/Sn0Z5Xerz/e4WwI7wRc22uWL176RVt1sNTL1FZYsDXOJUcPo9a94x
A4NB6r9PaRy89SAUk6A5qL1E5jvkd/9ryEtnVvGNoPxwwSCL0Uc3lZYuqPqRfSxm
Pff156uFbVrtWlt5AroUQDy404PLuqPkr7xxEeSCdOadIIMbEgSjDcSVUQ2zI/u7
qinBTobt7vm+evwPYZg8KcXMCwxPZmral466CHNu55NZToytqOOpH50024B6XVWa
U/mA2+vyKUj5pxohfXxByVCUEPVMOXPpj2mBxBpV1MeLwpOxk4iHemsKpt7NQpbl
escOwkIjVGy4+8nFs1UvclLRtXsFU1SrV8Qo6PD/HXeBpXLA8crbw/BWM1uU12Gj
jQtRfSp8nR4sAR8BUIDnRtRnEUrp0FZQaw5a7uJYpBJWPB7PrJ2atBqHXkdDo7ug
/AxXkIb1Y74wu3C6yttHBcw2d0RqiXba4dNDCb8zJcsuxVZHa5QzZokb+zOL72oC
yG22fatSHACFrO0F5rZxO5AAGCmPwTocHOatlBGwU1/BUPzqvyWnWRNuZxD3kFYP
kBlQTLfFNWG2DbgCKa51IG/TneRxe1SryjVXgeU/NeMjsFB5wmTRhiQH1noIkgnR
bpov3UI/iVb2recewa+f9QbIOUyePP1lArN4hP5Hf1Oj46tcA5qBcYb2Ek3Cabg8
pE7aIW6x+5aPyltdoCk/uE9ZXrZfMyzBlvywdrln0uF7cuHokejipdh7+/FiykF4
166yAtAZGOku5AACIvi6SNe0yb3WVRRWjkf1cNlCI5mXVDxCNPO4ArQPtHkHm262
retkMC8Ble1Zd3tPpTNg00I7LaH6tnd3Yz4vjO7KSY4pO4Ndr5Et7s3hS3AK6hZY
TmHtFJJD8vDsKW2P+g0KZfAOqUwieXC8xJbo5vo2TST2rye9aGvjiMyakDwqkfIO
mFqzzZTpM9vT2ms8aONqmj4OkXX3+ZtKJZZpThjofCqXqEGK88vP8mN/2TPCVU0q
F84sNKDxJzHyy6BNrjop9674GyBtYpFRyzQixX3xuhpe51o28E8VvkusF37GpCAy
y8eDedlDzv0+ojdBda/aOyEVQg3NaR3cYrEvVpSZrF1uP0W/F16KAen94X7EN5AW
jC0+Yaa7PjJSgAkkxFvBaMBNlVnbLwMQdEv3Hp2jlz6Ko6L6RgtW2Beyf773p9r8
vTkZSZh/9hXVVWYo/a/kE5go6+g5o1j5znEQIPqR2lvMAzP5e0SJwfuRyTk/nG1I
hO8jWpJqcyIC+MwuhfndR9UIwKfJItDxUKFNiWse4GrKok7UxRxj+ROtocDdieGR
KlD3bGwgtOhUjKLBk+OJTkdKp2JQIe7Tqp3gsBinOlyBguhddnwvCN8YSJmpmDDn
9sppkmyClpiFACBGka6XhFudR5bfVTodYMIfEr04ysvG0exgHVYWq8gPC6cJpVgI
MkP/v+TsAXXlFgingTy5x7XQO/KrcG1q4uWss3gMjF0WM2raAF09+PtyG976qQRe
rW9hC3JnbpUCVXG+uC8uF2frrVZrI/EYe1XDJXw5F3o5DeZXsbej4o48tscYFwqp
6NdfhfMmRzzKfzWTCRy6DX6R07RAPWRPFtK+NgC4JVJNo07PNZb4/4ElwEz2f7WR
NLngTAF9Vt6uaYgtov1SG1UrkMtNy+Df10mmLhE+UKIGMT/tm3oGVXZKPhCoYpXC
kCqxRrFgQSyfowUpeszNy5YWHh9o8XRH6kNnIQaH+K/V3ckPCoz2t/juW19J1tdi
drt0o+WmhC43YxHbK5UJW+5sRWRUgP8ysc3QohTnTmWu2fv+vtDE64hsU6HdBAsL
bA/DdflAjq5+N/NNR1VQ7g6oNMUNwXqhcTGDoQN4rNyXLHStXwYw8ZFFJSGwruAf
w0frmJ32RY1u7BTrXs9d9yY8tRAhUpNAbHEm8A2MJsI8uIVczSVld/yqHkhh1rLh
vsph9reRrgn89WVVXl0Jyb7hgO8wiS0apJcaEtsW8WEjh536/gcDTmDJxUNLiY7h
MfuQ13lyX4WboRZAbbqTEbMREQWLYU/MMbkKeoJdn+PjsgcXXPdutvVoL7PR1DK9
RdXbPdXulfYmjiu6A1+KdVT0BVlUA55uZbKy68GJvZBdqNgUl1YrJMWGe2rSzPzd
9rLiSiU5/wUPPuS2CmTXBUZSqmuatQl+rzS+G8DpSauStVYXiUM6lpy3mhWCaK85
UTXGPzGVfH++Tl79iP/bSM8HGs3a64v7ndfkXih9BGeFhirVuQbvanQRKpJEre/C
agRjgSMpicSuOnGsX+BBVKTUdUTZg2WW4PM015Sb0KbxNT+pQCrN7lrPddoVX2mb
KF4kioU8SYAbUS80eMp9ieNlTFEL8HERqTkgMsOSFspqjD7m6M3TzBaGbCfdqPRv
+yFOvwjUbdunIuo5dVdr0Sr8OixFzcQtBnTUrzeXIp34vg++3nGLiYFYKrdBjPBK
4MT8FisxD909ke8I2mbqhsXOjgWJn1+XD/O3r3FY+LSbs+L75LquxkN3D8k5j11c
qxIlTeiv62iy2J1Ez0LSe0fXZCDQnEWCP/KGMbG1BK5mJj1PqDF+u3RFGlXqd5/0
JFWaXzidAZZLHavwI0EAILwIF2H7i2MCif8Xzo17ZmSckdSMZ4rSVSbbCEPv72Ke
dqh6+hRUGjx1wp4UJ6z9C3fleK5oEbuVFlvn/s8IqnvH/01gI5FgTY6N1lEwQ/DF
TzVGM5QcPFN5Vopvzp8Z3IUw7Ku6i/Oqir8rAK0oY2EONjEfr4sMvgzEa6xAIEKo
SzCinqY5cf8onNZT6FKUT/2d0PLNc/s+3hJkfAZQSTOUmBpiMABUi0oO13pJRqD/
/Rzw+MrQujFvxZpB0jUYYbwDwxdjxDn+h66iOrPCPqP/Wy9Umc1oS9wK4X9QVZM0
ym0MTWVe2xl56ickhfCxW3Tc8PIFt0U8x4I4mme5hbJSa6rrE+d+EkK8Bxi7x2oz
TTdgGPJvCGh878+xCP5igzDkHQVmqg3xCX2mybP2QTItFPjyM7XLBj0Kh2ggE7eS
aXdYEC/KPDmbyZAjzRp6o82PDPRjdJziHgJLkvTE1IF3cXHmaC4gB9Xiqc28heb8
TadNuyXLGOfyJ76wBJmVYyEbXnipz+QwuWXkRwM9u0AMaw5hauuaSHu1y12JKCMI
/I3dBiZJvIP61jVpTHtMjQXK6sCvua7p3Tf0GfJiqPKlL+opKgsQDsjvLevWOGQi
o4DeGfpru5SGrHvOW+5zYtYkVwiG0Qj4b8VEAL+3pRAdyIpE5JLddT7riK5UYGFl
e5tRYJRXbOwHgn7CrFi23FPT6sSLLib2p8K/Vsi+WxjEExr1InCQ8dlLA3IQeH8s
oT/+1JKJoDNJd7f/06JFnN3hJx1Evn6VgzljrIYCKhtSKA3bnzCNiqYdRh54c8FP
LHBBjCu39KjuTYTV8sz3nOsAgCN0AvZs32gZr8SaXeqN6zjp1JhTYwO0nCCJeJBV
FdRAeaT5wVhaFoiQcRtTnpyzLsQRQiLSNFixDoK5OKnOxb9k6pooxZtDEZ/f7aHV
3TCwM3wbUwKq6/YsyGGgl2T308ZljqODYedXje3YSM1jHF76yjpjceQvVJ2yGzs9
08iddJ8xhTYYq/J/TZeyIAh+qqrAlOXcNd11pfEpC1lgHR672iI0XpbmM8QpCfZ2
7r/CX6R0HrQCJvbSQa46dRlbhL1pYnVl6NYOIiyN+f3E1T48mEsnBxkG7tG9sEvJ
BVaGP1uJqjgcfnasuyQm/+rJQ4u2qD5fQ7mtGFM/75913t14LCmtKB2xSPnjLZ4J
3GHIafN18TBM5aYpwYKhgLFUG2ZAvRrl04dDPEYuO/HVlsfDlnyjvgJu6/rH2Vyf
uelgYVg3JEcr1f9RLN4vOLM7Uw7auypdqn+Jux34RW8/7prKN2SdrLPMjWG+UQoM
nKAzkfkOp5aSs+W1aez2Krwm799p9HABWRgRf5kRJtrGz/z50d2sdTfib0g7EuGu
TcEGGfFRCIIsvy3yc3Wfbx70X3VjiNJlJJiAEjr9WIOwUDI9kC4VSNBWTrXjmmNU
KaRzr+P+QZVIrDhvdPB0XVfP7VJlW8rnmfWAPH084cPVJLt/KAprJ0/IDTKfRQu2
vjsJ3YPXTe3XCX4+MrV75fdArQcCYd1CdwGwTsZk9BAzOOl4CnVQT2aV4nS0ZUzj
YVQWpmRgwgz/Jpis+nk1TkFAQInelDfmb5PXClvHnEtq7Tiqr0h/6sqyB+lJXoIC
UEqO6ZW97PuEAEbvI0oNBWeuu1XkkNl7T15OUSFLqoyj0IgHmubenhzWf4iSPD0/
PWt1Tl/u7OKfPJZStEavBG6L0rcYiTFnvX++GKe/a7LYqTvOcNPBv7olBz9oO3/j
UpVA0bD76vID8aIkL/kp7WVTkZWuIz5ZVDRwpnSOIQPt01l6R4VoAM/8Wlx9BIp2
CxjzoBnju37xL3qkDAXkkuN66ENH5ppkKAKiXJEazU1peT8CA9VUs7tSPec+gS+k
5+uw6VWfHs+50PLd4oHhzzSxRNrkL0/WuzzAW0KGh8KLpEFrx2UY2hEyW1xErFgc
dK+GVRnyhHyRofraGw+cKVEsGJHiHDx4oH6TN6ujVe1rw0Osmx16xF9qImvydWGk
1ofHC5QfnN0J5zKoj5Ba/vw2JAZ5fCX2nnNi/BHlK8RkUdzNxCWIAh8BJXAm2Byq
gGvSztYTxZJ/O85lETtznYkmEDbv7H6VCzDIXKp0+Q8QEyXnwYZJfGETnMdaYVGK
J0KSx+G5HnFKl8WFccfIydk7GR/d9t+cukEILt7whbTqK1CXE37AfBwBC1nafYBd
ZWxxmzfueLWAdBwwu7v3YJGrzOtFCauv261sR8/Y/nSOfbftXJg0qOOvPkbUvrTH
ztA+luVOh1kWRl87eX4hzlxSJJvftFFihAgFboLMdC8++dgnf5I6Aebtxbrz0TCN
6/Ia+kdk2j+cB9syqPvbv/rVBztdO+LRpM9xRauIuS3lpwTzuSGGFVz1gX0SODGV
nBQPYGVIvZaoIV/ViDwsyqeFmqWUlJCkTXx3A35bk2Kno9zvxCKY5q2qasLcTwwP
A3pvzRAIJRJXN51abbrpbv+Jnz8TFGphRhDFpMcelg0hP8kjYuwHtNoi61w8AMR9
fzMdPmye658acayGXlAlFWaWW1umGj8Z0UgICrRAQdGuAMp/HTEJuLKBD+cvgrbn
db1MAq+AIWzY8mJxJ+ViGkgaFd92TKVHxWEkEKgZozlPIznplLEhwWKwITxOZp0+
f249Lm0dfakDc34/gTT+QOKRM71Rc0tICFel0jMWRqzMQL8SCrgRTqkpZvRTH15e
XK/IwAcWq1qQDJ4awh6UFO8V0xZvmztz3JYpfar3sOzd1K63MOCyIlfLdPZNdlx/
R72Av0JM5azZ8arAyl2iNMHqSKJFXGXswS3W8z2mZZ4F9uARZZJSsPYiYAIY9Kpo
ZTtHj9bastUSHpZUJ6s1uEsfhR6Q95nU6L+VeENtvL2HpX6HpyhxTlEM6OjwaKL4
MhMP94BL4tkn6n/4vDSl6rEebdUJ4GRwi1TY4QVngxUvBwT7FpxzlKJUx/XM2mrn
KN2mfD23LtPbNxofyGf5dLhn9ogZq4fZofMths6hjTkyeIwbYPVB4zGzK2K1ycWs
s7DTtN0MAxb5nAxtHvZft5WVSrkjQlc6shQRbNYiKaUTig9enOiTpzx9Wim3PSF2
eMX3JXX3W3OIgr0n8voHK5iFa7l1YoYuHLW9qTCB1Q+XgNwZTDBDSpdbUdgxDAsj
yVEpXwr3kNGOZ+ywL5BfLuqBeq9MMAz32vgIMd+ELFLTgXXHKN+D3AsQHGzKXFJp
8UC8Udj+KKhRNGFu7MRBYYk9zCGxV+tFMoyYmLoD8xbN0kWxygrXY0qDgF6riX/f
8GbRvomZNCY27lslZGQx668btteIFXcZVQ3JtN5+SvcnvBc7HZ3Y1l9UY22fi6KQ
6je8zA8jiPlpdGf3jvAPNkzvNKV4l/7CgXOiX5+oDUlxQ0K5ZoK0EAjGFtJYexTd
TX+54nKHntKQYJzDAwdUA2kIkl3p1okrK/boB9V5WP0gCjToNxnyZel3eRi+lQ2K
SAAOjUF410sr1c0PIuWx7Hbj7xSUYCw8TPr3JUtF0XjU5RdSziHODWLnu2CdET/C
jldztenkofcagmecis+B/t1B37ko4noNJUF419QS4XXhJXvR8poZ1tlbC2gZ12GU
dA1G/Ob5c2yjJNCkXZ1HANOk2pnd4yWgqZdH4w+wMGDE3rO+Z68XzSSMk2vFe/Rd
AZgtiryBcwE1PS8HutGr6pO1BJ/grSRDrONR/fue44znBUsBUQ+1noatULOgTU7Y
VThCWovH4d6HoacMDQBcjtENVd1L2gdDPT7CRPIdGAuWxGKrEjg4qOctSnuEYobp
2PmsMKyTtAzEJecavu/m5MqB0k5VCvj8nAowpk6a3ibidp5h0ki8SysKDk++0KXm
yuE6aHLrCO6ssOnt24VfTpPnoFlJG6RqxMBmUJIH/3SfLK/96X8jzPaFrI/33dr5
M5aUlUlkmptYU+WV+0HW8XMfYt7Gv5aZmOzMl6wX660iS5jQ/rSEhnG9rZDrrAMg
Wbzef7JJxhD33zd9DseCBqYPG7rZyoQKxEvC1Is5WatTMVBBSwSL+4pGyd9g9jOB
wKkm2f4cXAsOpBCZ0euTNg2STjypZ9FrV1Uh+69WAE7n56+zFOAbxOEjElNJlVzk
g+odNiLJAnorr5ZxOjh/wX3E9k2OQz67otyXRGJeXjsQ/8zHImCi5t103xmGzKi3
3tOQTu+z+8JvnSabZ7ECssXdivbSfA/9HBNZSvaLs+WXNpEVUZphXg4PGwL6ns53
PqaCGKq0aKikCSnLpp2SfXpyoHXZGLdqT2ve4C8TN4lB+QyJRNzxAPXNcNa3oFl7
nwCShbpykjRLkqZvqT70XS5A97aDWGQUmqQSYZIZDIF4Q3wc6evXBlagVXm64mK3
v6bIBaDzcocLZ71n+wb6xEkz3x3iOg/xZgJjhlaj5p8eDLimzDUDbttCnY6/ILKG
ihU934mjpPSbNpztr5k0wYBtc8av1gDWSFHZ/KbFegp6UqipjZRZ86BJK8v2freR
ytVd1t97Ys85sbD8ce7sxTq5SvJUUrRInR2KFR8aNCFgEsOvr9uJxEjUsg3aLsdj
zkKAC1j+BKI6KI/cEFr0Es/mhzLJoR7PZGlstg8SLVPXMN4qAaGLhHQwJxlRz4bx
a8rdC4AwZcEUumBCGXusu11hUEi9/GAEvk2BkWYIbayFuvlxeH+xWxdsxcoIu1Tr
ZD87qkGcyRNDUN5EOh45MLwTFnZ6FG2asANjJlvJ71kgZipx2htQyQkyJEb/MfVX
59KagexvIHrskgVgZVhyLe3ZLGPKMEpTUbsQnTCGFwg5ohafiJfEbMu+ewmk/ws9
4awksE5iis4MiNnf4al21wIJyRskgIAJJreHtH7driw7T+gM3qUY70e+QEDBBDMZ
ThSJoCw+FA5v6ImFcq0u+bw86PXJeuhqj3mnpQUA8rvAwf8XRIfFl5YbtVnJU/wK
1q5997NyM1Edq+RV5SBzqw5JD4k8cZSTzNUjUvo9R3iJrIGq7PI0EpKzR+q45GcB
ICsP1qDyK4pPuCLUZYjL2DI9+YsuN5sZUFay8cJCMFB3SNqAGGSEwNr4Mdck+heS
u8YO3dcyCBE7tGlGAxFHkECexMaFluPAZJuJIq8K809w1vn/QKpZtFzQ1kcm4Gpc
awtf5kgp6yCLeFI+6Ndqh2s3dcMsk2pKmvvythYdEICfM2Q4Aj+n2+2s3Fdtphi1
3A4zit39sZ2UQUOSijoI5jYPQ8eLuTJTyrjcghxf7vrsoSK9CL55bKt+/sn57p2p
gKgGhPSXjOAACiR8sCY32yq0XtxGYvSka0YVA1e652tQ5uZ5HiPlBLWMYTYonI70
x4VCStuIwvkPm95fDETLivq7q5OAocbUTg6iPEBH1I+bbYbVDXsjIW2jvNR04Yi4
1TZyVQHKQNFdX6KSHem5v0ajVg4ptaHlKq9Qg4FCPowFDRkV8E4GmkjY8XhHx/DM
IzA9mue5xjvbuSR7OXSh5JlhUI8IA2H2xVyrNE5XVdkRPdWZ8G4xHEqb0w4pwOpF
evNbWoK6hROaWoAMIBDlJe9Ek+A9n/+1ftCvA4L52B3uzgCzKEavt2FCcL4c/992
jGLuPocP3UPEetAMhFa0x9bNKgWpJ0tqxm9BG2JcJaPLFZvX3luTFu8M06r9TfXH
Sx36CDv6GufHaF+BxRW4Yo3htV5nu+S7EtAl7qb/y2OOLtbagisVwSishXLOz879
NoYzVjZ7S2TzwWMqSIQnupYTJZYCOAzHZIbjhfVaE2+YBpzOddyJDqkPYgfzzoyL
6H99uEABSlv9nz7zfUQI9W56DOXrhg5+13mjYRrOUYM7XvggclRCdsaa4ZLbk16M
fi8dhL0NGw0xmrpOez1GFHeFekIbCyIksd6mAfPiDqGKKzDB/lIp1U95dh+OaCwN
P6NmSRFf1+r9w5Mz/2qd2LktItxJtvZLw8jAhUq/1sVqSzUkQWQeksLhYkmGOYBx
oZoawC5RiVdctqIWh1GHJxYisAO0N05mIRxa0sPafrxEEjtrGOinpU1Y7r9Kifyv
WY4uBYkqqnRcQVjE+BKQ+/uH2hONQ/jk0Uci8YaO5H0EcNGY84PdeKOEW4uNmphe
PTjTYEboeGAvkPP/5k83eK9arwqqKF0vmJljBxAO77f8sw+EII0aSfN0aoLfORBP
ZpiudxmBRqIyW/L1iBEQvN9+yvN8UbsOGdYWYFI3HsUI4DSCR0LUUw7hpTuBmEZM
rCXHsxx9CLfbYXqmzzKpCR7FEdnIb0w9g3yYix/i/4kqehKMgcI7klMePyjSV32Z
viHLe4uBbBAqH2XmBQYVpxnqgW7vOhdbXu7TWuIuhokXU8T+MW0dreBiON177EsK
bBedwHH3csTyH3tyi3Mk795ukhIbnqmwa8h38G26LF91+Ig1wjERQKsMNqpBYsAq
Uyn4QuNwz3ivIIQzHk2+LZEqNHlw38rwWS4d3hA8P0r1q9HfKiMdWcL/bs3FVpwF
a0W/sDgnRJIp9q/rTSmXFr36juap3HcMpYd4vAfhbWYyH2hMP2Eo+maGe3DY9k9/
oWiL8sNNbDeJJ0OgApCcnifCcD19uFutHLWMsug/AYIgdWW+JdtIBPJVuWW9T2Lb
bfTdKsfKL6oS88F4EZ0SmDTFIR36hzakzIofx+zvEcZ7pePVtBZ3WnTnbvaS3bGR
nyPRQF0pkjJCbeT1sL9L/y2ZQN4BtN6/HlZ/EXIJu2w81fpsx1a8YL3WsMzPZkeT
a0XBabFZS/tgyLc2rCWTVAve1epKVJJtdNIYuuJMhXlZNTuQ9swkikvj/etGZi3I
+zgLQ0ZkGm62iwn+nHane+uIS14ghPHckPys++zvWYoDV+SVVarEG1o/g3BJBbE2
BPWrQi1y8rp7yKjIL09DPx42BUICceUbzxO001l8NWwQpC5hF/pssQtaCSVkR6eD
ean2BKTn2DQermBdGhS9oJr4ZA1eFEyUiZO2JVkWIbfBzn9C69GYoJXGtqQllc2C
e4z8Q5hv1AdgQsJ8E7/L1nGWrAbkZ9iocEkNBu7LtXvBXtb20YbinJXtR9Uwd09m
sAfueHi7qKJCDbcjVBko2pgN1zMgSj82EUgQV0BZSWfrrwVY/GGOtyYlz5IcGpMn
xYFteP+EDpBULFx+y3UJ5QO4Zk2cVZTnRD27LEccn4ozNXjtgk4IiR0uTi/GjegG
aCUd/AU7/R7cSONYvxLVapx9zhE4hcc//5SN5zgyrzd2IAdRM/U+3nWRweIWVyJ1
gi/hNSN6t0JFfBABjkBTr145lrznIcW0ZYShDEQbeZlvmrCiB22K1n2sBPEDQr+L
El4NjyFKMOLdtgSO/htqqB2ZdapAc9rQ8HY1PymRY/AHzKYQ4/fDt/5qgG/CwpX6
Ihzl78K5RpLf/NBF919oZLQiNgenk/UwG3QmeUbYI0UKSeQMGjUiyuRT0C//lMsI
Or3QZJqQg1ndA5PxTWeomVnw/u4bJ8jINK7GU8buybRwUZVKHv+DT9NgkRl9ovbm
rP0CtA0AcNO8JoxQ4znI+rj5QfZWbbtwq0IWfoVSNT9mwXyCAAXAq4ZvJnv+54QV
hoFGwSuyvVo5iegGtaIdyR3mW3JzNwEL3OHiTVpE3YAubsIaaSjbsPpJAmD9b91g
NYNJMfg6XWHeiSXkDQCaEmvnSQFNvNJqMJSlto2MIGZefRGb46r2MlOvvwIp7guM
jX4/aiSD4/1Cm0C55Ip+xmevROBJ8/fWNZxjQKFClVvz3sKVwx3ppyvHDBZXbzbF
z1wUqDuDE+UMn7kaJXT0XEN4VLh0xGh4etXnMpj33M3dwa+p9IP0I3lXNkeOFiWK
zG2kurBAhq3tO/tmzmUTHXvtVlbAhZWeNmKtWBFH6xIxkYKARN0f89dTM+z6W+SP
nAcN76jOFpzb/UV7II8805WVMQxRy2dik2FZknpJzpjJfzsyTZCkhZIgg3XtFtHw
4fIJNp4JbBE6Ox7KhpcUEfJXSo+FEuj2GrC991BBAwV55+MaYEu/zFENEA+Hwy2C
L/nqOxgUHndI0/JQldAJrNa2DGC1GYcehXGcgJu38cU+AW9OEMv/XqxEsymY+xkI
a8qCNXsU+VCKd8Mi6roejkMZMkQYMIfoTrwynI7CtziF6MRTjur9mlKcLatjj7dY
TWvRxnUGknzV7CIjN9+pcOF7iFK5f6PKrSG4d5N1nPGrvUg2V/FyIfPrW/kUgKv9
rzi5AAUedtZudH4iNNteNdQCmCn0W+ZT/fsu6B1XnO1CbLrgBA+hk4kHkJduB2TC
1p9vA4r3yyZnzZpm6+ukAhThnUVeHAh9fn9UOkOSx2BDebnWkZdNl+U5gi6pYNM9
XeVM9xcd6kVV/k4GcaXtUMrvxQYg1e0IhvgjaCfofFoMTNJvox5vH8GDo6GWHPzg
5I4Lr8dTf/yY2YL8wekl5MaKqxU6NspcXzKYoUc6HB96rID/n+W2NtjUryfdPNHB
FbQt0rXfqLtfez+6TmpVjf2lLdKvDzbCJGTDBNAKpPukEgFZLVtiX7Y10rTckg4j
JrNK4GK6EHpCS/DlSQVISjwLoPX9NDQvPi395lbvUpDuB1mAN/a+smSkXo5ufr8W
54NK3tQ2llqdqM4b5FM0Ths6hbSAI5oHsUR/b9LiIshTyjI7uCPh4s3tdi/OAXsp
W1aM2HlwmrlwoykYHwVOISHK4Z4c7XZzOPuGx43Ner1KouWLK8RazjBiWKxCiHXp
czn2cFSxmsgNhdGLVrp18zSKwidt4NXC5SAhpXLA2QpOu7VsM1P5lompPJh79jKi
TNQ2M4/4UBZgLlWE9kCuMFLkRnbYQDejWkwZf3nj+OGISjXP7Cde7FjSM7VTms+G
gG9gJ9SySiOczd2zC4OrIuukPsjTHzX3y1m/INIHreBUlJAijNEWFZ6YQbrZo7cT
pKBroC2gVdz1yICmQVTnv+SmlzdTIQfi56WT4n2Mor21bexuFYdXWQ/pZGOpBIRT
dnroz44TsazSPFS6wx7Rw18AEpBg3+rSm9FejLcHbI3MXnCfXvIxm+j7WTC4qnni
23Rd17h6NGaVTQtrNwUV3O15cnNh/KRqZg/eSb6NCFse5tnbuGHk/mYugAtE7GKA
wRmJ9uhaHZfMZl+Ui0FD42ffRfGIKY799VTPbScaIp/5vxwXbb6wkgXAPzz/A0wb
TF2asxiG7hICZRjRFhZdARpp0MvugywJBWVGGYLk2jy//I21vSRNseVydkRMwr6D
MI0uaZyomoMkHzRXDPcoTcudaZ4Nl+RY9AeKyaPvL+CRh3DthwqDecto7HR/3TAc
1MWnXk6zqu3/xKNnli26Cm7vbhMY4N5LqBsyLsPv9iXEcnLcjNLbbPEdugxN7kTH
IlVhlec9Evv9wIPsDaxsX5yGiwF37fOZ5QDAoL2iLAUwHeENNl+uTqdRuBYoGDpm
XfA64tW13yuP1PuYzy8vWySQ0YXP7R3+/mLxk7+QSVDtu5ckAP2mGJQDXy+lT01d
W49wzfoqKO9RHnDbcVFrg3/er1B7BdmY9TdsFm4FWatvlz3hK07WS9Kx5Q5kYs5O
BLRRRbao6YfzLikpJIU8FB72Be29IL01K87wau1EGTcOpse/eibaveRe3WToUUjn
ikrZ71XN+vV1yXsc2UtvK9RqLGZP+T12RxwVIr2ot1LS2mhMl286Znvrbd0tVQkE
WzdisbRniG5JmqRG21y9wI9P3Ijk/aT4J1JSgyqmNZXJuhTwZPmOzGtJaQy31qqb
vXMqsTsLAEypQJZJdhP6HxfQ2ZjBef71JlVysMrTq2/pauTSVD7ymK3Q0bDm4V1Y
npDcMTynwbTOfFXYwzsc/mK31LScYPzR4b2CDk5E+yKa2o9/2oqZMCMJbQUXx89Z
sAhVIjYEE1v+RVnLdWDyy5evKpLYzMZfmBTmKJayOdksPbAr18i4/KgFZF12Pl3T
SVoT5A+HxpW6FkynILLMvl+5WvEfQvLnndUmhttl5BwApYBBRK7TSGsEHsF+ye34
y+bkw19k8zko3PXMBbAHSZiEX6KYgWktcE1bGCmax/yWNSDNdW3xmQCcZ3en+UwT
7pGfvnLkuuT6LhOl/B6VeEBdEA+AuBa6IMtf01p0m/AX/PLB3M6p0XaucQIALkCq
7SCM5PCaPp2Rgp4Y1rFKfX3HXPgZkrUK7iEfrsUBaJd4w2NOFuZZY8rBjLGBnXmy
j/NG2btRhlM6JshJamYcTMAMnU43vPJ2gBPKuGMHi9TqQGryFLEifsgF/Cn49xs7
wXfZnW5wV3FLpXqfwwha7/TFV067wlefcAvPes7AosFHsJSK8RTtgsznOjGf1uYu
1U7J1yUnvaormrlXCChq4JDUsYlZeszoZGjjsikw6tZk1ad+aYbvDV7sUKI/4c6b
AyY0Ckb8XjPWcWmFWNp1KgXrr2aVuhxwmpu4XGhOTE6Bzdtq8xZaoIW2+NHwXT9Z
C4Hl3tHuWmXN7p/VUqRddnxewUajyOS65n8rngoW08nORDayuvx25wEcL+PSnpVk
fiBktjllX0SpRVjdOwOWf38cNSUZnL2xn+kn9laP9++bVHLAeVmTp6zUSwGVKz5e
z3BpSMdxeEXxZo2cxLbhVn202BXo9CNOsh5/+4+ysQiK/jP5NfaJQbD/2Kbbh1r/
R6YTiqOavDpTaWSYuB4uWNs40PcLeiy9NkSmNj0ED2dB6FuKi9vYkrnQXywOCaCK
iepiOJ1z2x63D00Gen0CIMqnlaskJpQLVDSTGc8desmE6ERMAQm436ldWMtl1dC0
5UYgF+f1l2Q1qcInUjVB3prFWWUDsAwpYG1Mc6zP3ml2i77qbICaTsEpNZVtDMS8
YhGUyKWWIqRzCXp/nP373ekJboG/mC+p7KI3NeWL4/GpwD8rsc3ZVal9Ocud98oF
hcC6d2PcU4Itxx83pseVargZVZYewJkLrnwGsiQJC7ZBiGqfQWEynaeLj0/nFBhB
vH8BuFfBTLrmPMVNUeih8ICeWggvPfl00K4P9QratZo6vKSeuC0p6OEcRBZHakQZ
lm30Qm/NpcejtnrYg8E06DfF/PQFPnwau1uoMf3m3LxaafU8BMbVEaeMnu3Xz2Ur
6qX1yK567JIJMrRTTy2omvNmy1sdRBxUbde3/SbUOI5PT0iuFxcnHKoIm7D//D/d
+hQ8oEHVg9pvLEEbQUEUvNaQUaYaivlQM6QnVu2XbxinAR2RO9bUBVtYdfLcEnY0
/gTDsa9vDzw+1kS58dhfILAtjVNNkyCw7S7tIjjCmBO2UuUmgnILrNc4HHGa0tpq
9PlveM5CCh45Xqw9ZQNMbJJRh/NMVzuCwYHmClzF/vkMx4RmPLX9xGbs6LYZoQhR
0tjwE5ToJ9zWVKzSC02i/2WMHxGaK4oHzAnF/fWk50aLT/yCFMS1UhOpKlGhUdtK
/RXLzH0GERlbaq+aXgs5+WXUkyMUVdZKz9xAcXpumkXcG6ekPTZMNNCQZMWyOpxK
Y6ez5llsyBLdq26uQCs7926d+vJN88RjITII5XOmVNDenCk8nqAaWtDz5GgC+SBg
NP1qLfDE666HobBHBklvBsJWT0b49pFpLn3lk4Io8gSyQSj0m0X1/PKHHrI/R1XF
AJLVQBxfVQvNwakAth3Lkamg1p5NQVl/yePUi+PsQ6y72J1yNRNuCiSlesYsOeOU
V7YM2fnPeOMmRz7vzYjC4uv+WG7J5/xz6aY52HxunqM5tCnAwknBfOXBUd1efsbb
hMz1sgjsKkZkUY1iBC344rlGyzsUhsF7VtXSgfuLImNcV8qJuAXDXy0PCY2tPQ+F
wlImT27aZCBlaDbJjjz7JyOfbNw/KPKeccBF5NBY4DNAdPmUx4vqYSD/PDn4FTZ+
7uXw8KW4B4EU0ynVRRHMvytHF14Z1iqJXbRFcdItunqRXY4tcQg0kbFJoTldc0H0
51GtnMe6RmAvAfZcC5fvBWn++aaoURJ9Imak7ibquIDyhMn0k+WXGp+ngdWH0ClM
UFxBmpVa9l0Bg/Vt0PeYvg4EVkf+7bm7UEVP9wybJewWpCO4UpLxzFtYJs/oKiOT
GDHYcqKbirngm8GhXXkz6c/oNh9Yvcmx/LUVfpAoyxfcNnvUufPBijYcSXOSrQ6p
4eHnF080GUtxY10ngEswn3LUUnkGGdmAjOM5lcw/BT9KlHvZBRon2Kmo7XOoi3Os
BkbhuBMOoJelvegQbrhzwq0Jx/o2Ge58R1PDofkhwG3m2WCQ7taCjgNuA6TCqx/V
yyJYx3Z1rVrzSt/Lr0n9O+20gKD043y50u2VR1LdYDpOurxQzKIH1++ovwalxydd
6X3tzWshvARkadDSHWGemgJnQsf8Cyf2X2jC3d4jYOB5yEFKc87llwd+PwEA4Srl
vZM8vYAZwRlFTdheE5D60AcnyCgfyGCfG9g6hHLl+AEUsw8tpuV089dXsGQw9+5X
j2Hz+4f/n21oPT12xblLLnS96dVg1qDQn2T5SwEWDD4oAa+fvRdmuQZ+C2mVQcHu
g3Pc3DbgB0PQ3McuiqjRwyNLyjw8DJEDbWznFzxC74KHv5AiIsfjJ/sxeOaU3mxe
5rBLSxvM2HC/VxsZgvaKS517m9Nbvxnpx2aUQXzFSO3Ti+UGF9YyrBOUqJn+nZ6f
/E1Kkram+58Q4v4BepEvzF7eqozMes6ZtdAew2xwdlY42qY2xHVtK1r95obVpZWh
DV+sWsEmpTEFJkWY0CIIWCgxTUxQR7bHSpuwMulJZG26ASEiqIsA911/3YAcifbU
WkFjvjeN44fT3GAVkFFEmKeixXE+0aubHjTdwJTkCMETaf2DiOFrCgz0bllkQ8qZ
Z9CBXiW70rEK6MfmEhkP7qjwRlaob+m2ZmZ5S0cUH5N32kkZnMUQsp5aM7DuKwBm
3UBqAKzBQmLTWuBqSAY4TeKXoLTAZcfjKHcjJt8Hj6DAQ1fjm0JVO3PdHL1pELO2
iY9R/2RKOTqeHaHeKnovGSYpU2ByrJCxcjaWHzfNiVYJnOblsnkVKKA/EpHPLHYy
AzpqC1Pq1X5+HdOsrccd3bvrRWC8v/IhqOF9OSwK8TWiTx3xI66mEfrNloBao9cr
ZjcX2Fhk5IkzQPcvJ/5zGcXqPDEYYesc2iQgCxFulhafBqlYsl3dPsDf/ieOILqL
p+3INIKfJUn5wmlusLp3gvp92P6oLcMd52QT5K0FU6R1bNQFP8aiy4WdFQl44Tx9
NaPsUn9pM21ywfb39sRd96NbA3FnP1lIyXi/nn1NrvaojvuyiQcYdI5gELU1CuTA
L9W0vYoz3PijyrECI5reSs6xyWycYdeb0gu60gQyHQ20l5cvf0nfbAc9ruvxmRWG
h6jcId8Z1BEjUV/3ZVzJ2BHdj3UPmW3K94dGGJs38OGbkPVv9GBNyQ+EGmpJzkiv
ECCh28ufpmnLUOC2FBkuOD7AQEwQ1rCB5IDuHniMUyDH6Vsmbs7gl71j9VcysuFZ
m/QrsDFf+onwfuUbxzZCqaZyK4+7Kg+s2oCca4n7RELHldoAmnST0mnZZIQ4QSLh
FzZs5O+A673av8/MDuyx+/UtY776UvhkBGi1XzIux1W0jggy0HyQiHP91wwhoAuY
s/WLES/KxvEvfZbtqdbt7hjbme3yu6N57cJRfANVwBUWZ3kovWbR0Bu8B1xwT6Pi
OzvLHRdZted3JGt5UDZi0e0lEZn0/DKofoXgDfbLReaMSu+fDznS24qtDYnDouXN
98wjDpgbUpAD7sr6HOwAc8gsoshSOJD4HVufmxmI6/5alRK/mhvFYIN/U+Y2jUL9
emsyok12sFqDuiCuabp1Z2tJYYohjl+dS9vifvP2+2sVzSv9k90agbsbTd6uXPtS
U3LzneYgnGn23qwul+66BZkUaJm65ju+AdgVLps2MIY8lPQdtBd56dR6vPPCvy3I
secaOa+CgwECdjFIKbMdghdPrcUiqYBocy4DdvsgZXgKS98bwgUZQUPELHqAJA1o
VWWtpIUmoUU0i5retIfzZ+iGasQRUWU2qp8ByjPuIFULgNtuH6eZRel+yIc7DdEh
67F6SLIhMZfkL7QVdjrGBQLkaCxEYBwPqCzOtGAS7sgZjnnM+p5Aqp8yATMPKbBg
nUT9fRUW+RGGJGFMhHviTYrkBrWaBaxrtrBhE1YbSKXS0MeELO0wSfvKdnmojGU+
l9Gtsbr3YR2CAvgVYdVrVWszmB1mSThLLJUQApLjDyA6XbKocMXrgj16RFTDeHwK
Zx5Vmbk4uK4xQwmdlt5y5LA4GaTYOIhr0GFIH85vJpu5T2x+yGnTQjc5tsGluKfx
21DZFUyIX3FulIZrdeIJ+SnJueqTURac00kdvspWrmQFj3oRiC5gxtpNvr2vV/Q+
hxcRsANr5BAkovnK/9cuIm877E9dJiRJ53Hp30dXQ5qRZS7qD1hWtov4ir0y6SAK
IVgTIXdYdbHV+t7bWU18iLQVq3vDpqT9f1Sjv93qsbu0mQTDg1jBDhzx91OIAu35
DItI1mEpJulK67IRH1GApw/a9WdHrM6SZZmCbIbZIYsR32yMXXp8OAgES2FYXG//
a8OrQpVWwcGtbe4E1JzcMqfgX8XtCQon3yWH1sSCDycvNC0jajJQ0L+ZpURI5Cy1
p3E41Y8VtzCVOM0s+vctIkYHGfRY4vclN/wk38fOO2w1+eEtGPUf+BCUIGwqCN1k
L3bu066u7IF4uWNadoQUf/jzKqqpRpJZ24soweMgzGDgK+/IFe9PBtfT5ijIkEiE
bzP5zxvnEcoUrL8ELFrKENATM8RgLECy8Q9BWCt9YdQnC1ZKO2u5uQMNRrlNpkF3
FB9QlZxrwFArEEX+tnURLKsFo1fz5HptpeTqro/aZMgexeyggtGVw0eJ/WaHBL+b
bwo3qOWZvI5fdwpl+rumrsdgR0GXIZBoIySSobvf+22P8EnF3vowEtqtxnAaKP27
2qxKbT7zBLvUQqHv/R86f64slL39txGcPGxgSKV66U9VT19dP2tI4DtLZxhluogW
KKVgEOcJeb64qFAaBpZqWdr2B0+OtbNhpMHtJ7j7xNT1AFvq7leRvZZaVcqT+69Q
bno3xkfKm0LC4CosryKw7SXpu++UTCVjfvWRjnvOXOTMuCHLwuDc5zbwhCUt25L7
8imzCg0RsWqwUyNtHPMb2BDNpP1Z8oJdNJFvS55/Z9Ll5iIV/LbGJNo7xzFoT9tQ
M3ZDNU+ndojMqpNuqVppap4jahQmB/VRWh1fejVbm4MvFIvX5xD1LJwI8oBD1d6N
xK/9OjATSWfcAVUcGfZn+74liqfRrHvfw4Js6EUnIBLQskaHNVq39pqyU9ILy+7S
8Aj2BxY9y3YWwSyV9TvNiBJTREr1DIv8hGSM0SopaSARKKxY/8wKlKZshwqlVdM5
CBGDjei3irX2PUSYRC82VrnJruyS9WMt+ay9jqayxpbnMWw30WYjCIRgcbEBE2TA
KPQJS5/LDAZWIkWmb3zCO1qMwbHiXOsZA3Opr9pOpnFfMiF9iX3vtwMLUM908f5R
zKhFQ3JJd+4hYFrkrw9DToHpHHxIbkwUWxxhTM2otDYAod89/NfIGc5m5sQx5aUi
xonI5qpWEHUjyo+Dy3aam/P6PJErRmixiKL06+Kr4mlTx5ZtLrwfAuZjL8k0TtN4
0w5baSV1dV8OOM46GWhzTVeIAPGAaV+jcriI1Yr95pwbReVP9OmPGsCJrkHqttFp
Thml+OZhlKak/aCPkUhOFbpp0Dpc/jps0qBujTvPrNeLVUgqSHUY3eCzdzThIYwk
RIhE8yKU4NbUas1Er7GQqm+vAoA8SBqReDTph38uY9IPEDpIik2VCjh+rGjVL6+E
TYNIL4aTy3tldfMLWYtTBJx581cGAgTR9W/Tha7GGc06+DWS6Z7MbD9jccoiwzMD
h3h2ls37UZEHbIslTpvpGis0YxZ3UADy3smPRKVuRgi2zUnYUdz7Jgmjs6t9pwl4
+iObVuyiSyL9Q+npxtEr8CaUkIVRTxQ7f3muNX6xLvnuTTKJ5LoDapzUdXs85WyC
3GcXJTF3J+K2EVg7MF7vWcNKj4KMm6Mal4ySDpXkENCOWBTRLps8ftZXey9wOsTV
dIFNfY+VubTO4rF/YVBoDI+9kpNxzxwel+UdeMMr5DFRQLl8xSelf2VIJ3QCUoR/
a1r4bXOPXZXONtw/J+7NE+F5Utm0Ihslg9fGGvegQ4Yd/2fR76+9dNJKULQBDgfU
6cNTRlPI1VhkuAAIPAVwaIoCdxJZD/gcIysEZnfHFqHi1ZJx14WtbBtgvMeK9pRq
02hcV5BOLB6YjB4DwfonrGdjGAgfnek9QFGgo71H+1PGm36SjdsOucNbF9HhQAJW
t5r6UsvAu878VpzH7wuT1aMwQXVKJ3cLv5+1T56M/iAoEGbfcMMbVCPiAy2dBPh7
C+JFvmBETWosGyCm+u2wJ/yEjHISUcKD60p98c6Qi3YbJhyAT/UmS9zRy+TLzd/6
954lvnvj7BuJgQk0U0Montblb5JPwI4leMjlMOlL3TMKFfYi5zxlOQnT2cftxytx
VTJA7t0Hn4tYhlqd4qx7OVJ6IXdZuaq3aybDhTaXeKlCEFI4ifHkOszY4EEK9fMS
8Kjh6Dqgut0rZy6RVzbnW0jK2UlbgXWCKlO6JDw7RTESRbaVKqV4Qepv+KJRkB9U
PjAO9t4zX4HbH87XvtUpWhMdUroy2xDgE2whMb1a8zczAeNBoUi+CAIhky7SxjCg
RcJ3M0qkhji8Dq6iaE5/jq5M54r7FuPs9BRQdKV33e53yh4NJMBXfKwgv6ZXgm9G
MrwiDZgJe0BkW2baK2dActN5Yk0wgXjetVFAhKsv6VE+QbKY1t66WiX1QLra9lon
3AzByd3uSaRLGcCcGWZNPz1+i0yN8XRuZsE3VdRbb/af2augvyfSPmNofN3Q8/LJ
yHRgOHDgD06rxnINiS26hnE5p+JYrUf0k/7zA3gd3BGi389IhuuuVMhCf+4vz5bf
9CqvNC6X1TqRytumTgqPtak1UZvu2sZrtCdaDpLhcRp04hchO8JnyTRnPya5S8BY
LbbckkJvxwwfLHKUokr+yXaBro77UdAqalkdZmsQcIVLpn/FU18QqpDBqMERSQfQ
JvoL5NSiVmNJoUplIkefikVJL7rJsxJ/opVYhYErc/cCRQUwbpGVZg8i43oZ+OJX
tyegJofEMDTXCDa6q3cnJJ0ZkkaMDLew8mJEu8znQs7vn+r5csoWT9DsoZB8Y13r
W3oXJsfmf/VKPCDk4vb8nSTdDh8ha79KRE31LyUejgZWa2xcD7nCKyMSD2ZdNIlT
0OfR3TSm1zKgJ98oi0p5kMVXrC7tBRE73FoJDleStcuTSCQxZEvO8upijAn1npGl
7epFdeHRDUdHllnCKgbhc3RYPGr26j3FPTcHxphHT87VDz/PU8zaiifHFBsoQPI8
xxq3pIWITxGTMxvAMtROvf/gkLw6TK8WrcieuVzEt7mxuAgayzgfzioRiKeyLU7b
RE6vbz83IHFSgj0sI3f0zxR3OiILFP1ftVjZrIN8KwElHu6Fa15yahuWgCt9AwrH
6kwns9aDRocPHbfx3T3PLpBUXdjw+tuB6mgb3X59I2hSMLt7Fi633V94EmDG2IQt
8MgeKswocAb7V4kkWYuzfAa59TA7Sy01zweTgddDDKLeuHy/hTZ/WY6h/F2LmTbr
cECpCOvxrWWL1g+dsRyepJGyrIPR0i1HWVPxVXd5+U5IcLLcsA9DW1gNG3pi830P
r0EEl7eVKq43O00vCO7/7vMcFlFIep3bP7mMuVQzssw27J0w0LrdAc1BpKzrauSH
mt9RWNv5skiILZ8Otva1lruRQJeos+7xLrnzmv6fIH9sSgJS12ybhfWH0EyiiHkd
koZI/6kQtW/lsDM8VwQZqVPZcesBBN8CdpHzhRcIHyp9Jf/DaigNi+agxLx/cVxg
FTZd8kitv1SW/FiD5ULoqZb0djlZwcaQdK+WXuJpwQ62VOkHwVvwklhXGrtC81rX
mybLddpVYTLQMddVE83eq6CWnS1i7OmhnbwbX/k1GYd04hgpvKtDWK4ISh8Vn1XF
DkuGQgUkbnsDI7xqq++fgiv/qrUhu88R+6gbdr6jtdaYPl8HMFYkbgR2mMs7Bl+U
biPeoYCfjiUaEz/QlCgjXRdKGCwTbzp/U68yPpAoEqnkXZEs/RI7wvvCKbJQqAgX
w3ZqitLvhfQdumr9M/EKx8O3xC6l1yrw/E7AZ1Pxjlxa/XdnXluUfR2jgRcTR/J4
a1Opr7yreO+/nRsyJTTMDGMS8fsMjMfuekOSRKx6xilzfTmxAIZJsBlnyJr2NZlk
p14bCZEJQi9qq+XxWAyWFKFSDeu8gwUSNE+EclEQq6Twwxn+Ef8EFJzF2ppMxZSK
0xHCPVUZUwdZja5ZVtcq81cxfxPIzaB76pN5jQaEC8UK5aU/yu8y3LTpgtIXK/Zo
YJQPanmkJF0YVIszC1Rrxkk9aIKDPDSzDOtX92CP47OBkdLsbKhU94XqbZnz2pDm
uC7krLWeAwOuBh6SfBJcoDtrtf8pv7oXHEWW281ttSXhuPhe84ofPlcRMpbujkOc
QWnbbVttvbn1QkuU5CuRgouGNnc2kRD9C1TmL6/p1P7WIy2C33mEw3Iis5JJlmWB
gd06PWmT8iTp5s1joG2GTLS9bCfo+3t3hCTa1wFDo2NQQDk1YuUkQTjmIJ3BSbQO
yWFhH86H/fjh4chi1FQdLf4m8h8Kwz8AclrnxWfdykt/n9gwDYikS1gUQ59Y6Wuo
0wC+24gLhyifgKkugavoy2Py0n3/KBvxm+f+GyqA5OaRPcbRL7Wgjx+T2wJSSWLB
zuwx8e6cFmSEvWos6M3dd3n5iHva157uH/es+SldfoFjM1pZyJHkxh3EcYCE/SkE
focs+BXRqrk48F1kII1DgHGP16hxLhA9ca60u5QjAzZxio3ftD7cheWLsh05kQI0
UeddjGF91L+DJCdGtPQiVqlf6qJGTjt1vRD86DKttNUrrwhpBf4Vy1HSRDCJ6q1j
oP2EYrRkDZSj9AhE50CvsrLPjn5nUTQ7de6YWuMbb2qlYrL4lrb7H8TZ9ddeEJlJ
wvjqT/PCMf5/367AlaWCMullY+/U34oCcTxBbC8wOxhQH1W2oiWjO+KGef+NZutF
hDug6VJr+M+DqH+Mdwa1IJwoHpGlXNWh0/j/kjuJOLB6XPb5VhvwQH/BzuGQZ+AI
0CvcYfO4LtMCyLfXXUiR59PFEDpzVZXED7nj2u6ZR3zf1Pd6NyQp9om4te//EE5c
DEptJJGBxDuzPUIDLaFmlkWG815zVnX042hHRN9v7Nsb0HmcVhn9Z3uzA6edv0CX
9mEjRvyN98oq2Nv3jJOwowk06nzj4iMo9MTDnFb5lwTzA1uNLR2qE2Gbd66QcTYA
i/kN6s88LiPLE96NsjnT928DUvJ54XOtpwpgA8JwmXyhN5puxTELgwVfpocZT/r5
rmKpukAIgdBPG0/tYBsgDHcHS/U86rymErzGhCFeiDAs2WhmEKZNYzR2qYfEAmaD
ossLcyFZa54D2J/5DUAgPwX+7MPRKvtnaN27NO/FnjQ7cjMt+OIXkTHJ0DRAKpSW
ovCviBTk9rCK9qePoDYvyLp3GOj4UbjCX3zFtc6OKbFLPY0TKgS47eUXEVPWqI1z
vRlDzQDhSubDAJOGgf4FJJcsRL7lG94pVHk0EoVeFA5I1khrBak5v5FlhPU4MJEM
sGS3oBAwvX3G5D+MeOZfiGatl8WJh1rq46j4WKu/D517xY9UJRF065+shz8Jf6nG
Ps+s6PQ4WCr1vMUymwlpyo0/LOsulb3f8R5Vp72ua39vQa1pRy6MbA9b4D7pqVMc
AB0PHRJkpn/UUw6JjnAoIXFG4K7atqPM6hHp4ptvcYRqDI093gdJaa8Jy9G8xBQx
/iGIeDliBnPkkZByZq3MJVbFwqFVhnNorTc92rfQdXUgKawcmnwtW1zSr7AfcHnX
3FiGKfUZUGn+39pUNWdAjMbn5pgD7X//MlYywvTgYG4qa+HneiCmEmCNBzAN4pcj
TIEV97QSoSBdAK3FLT42iJx3xvY6IANOe8ArCaacQnYp1EbGLBtw+bco36VKXC6J
oTjyGDVldHTwugDPqJUsJDWDi9qf0kUsqIYgJKBMIOdBnqa8S/lUrlVzRMNBoGkt
I7TLZsa/NZYdB4c5m4EhlUzW6ocsLZWXpT6kx94wyvaBA0j8k9b4AThV4rKBfYdV
XYYht5TlHMqBL6SyRnfXitdVjQmw188x6vZLw/+z1eYvuIiIZwIvJ+KGiY86BDYt
Swcvb1i55W8UWP/ozUhzvBuEN/niKsNpAk4TlmIvU/B1lai94Bw1vD0Iejb8OEIQ
PaIbf9UklLg4Ao/FZ9JqUmJBbIClSYtJ6MDjweLnfbStqD9Ppxc2ckolkVJtA4re
yc/IjTujY4f+08GFZhf7q40Z6W6oV59kMAmkQXiGUkMRLvm6b9+LjkCn7ylgbXNh
8sSxum+jVVWu/vXiLudBoMmEp0NxyOqb0E0l98unljPhgCICKuZR3Xn9xNXneta1
W4iIOkMWBahmr7v/kRlmaOC1W5ETZA6Yk+rrb/M+UnStLy4kXu+icV6QcmlBsSyV
T/VS7oIbJwM40Ozqua/+ud/SaAD6B9kwUu/Kskhe8nO0xOQNYIDJlJQ+MEz3ucbg
JJSLAoduAU2VLN2menYyK+eyjE9D099HJN9RipSCz0IWUohSRVWk7W0yXLdkSin5
yllBjcZjU5m/+QqnCRBLUqeM9ftK1DHBWUVoTNTc86MCcP45SkUw4bVolW28Kj3U
ZmoyDAdWzzIPO0P6V64cGfeb1l7GyrC9ehHPdZYSjRtFuu0CuGPHRwvt2tX3JgVA
zEKMFL2v/dVwhG0vLIWTU9JbLyV+NgwEw52LTzkH7Rcud7EGrpybypeDkVWrf4MK
Q7ALEigriaEpT/2WjN2B46FMb1l/+ut1aG5Q/lCn1lRVYl//ofJjslM/+KjtOTY0
pS3eSLI3T1o6yKU8RnvlNgWXeW/xUGISvIg1wxw8zelCFSdZCShoVp0hHVYel8pP
fNkogGiogjYWr+nOeGeJOClxO2z9hHT+WaU0FeA4IdoVNxlaUhC7+i1uGwHZyjo6
z+E/+1GrfRUs8Clwco4GWNy1afEh/EinB2IWUXQeAfp+HhfT8nm97PSoR2pbIZio
+RZErKyyt/3T1+gGTNLsezWLObNrgc63VjnpykMXr8GvbGVFRm0du+rGxPr8nZ46
AFmP4UPNdTt9URy6dvf5YS01m4CCvK2ETWanfw0aIKlbwgv7z7Wv18Bu2KEmfm2+
P56iPhZflHz7+YGJ+4zyk7sGGVYoKaDE7wgTzhe2UR5eXbLrG2iskSfuk4dFFJOS
XFjiusXG745RIdovk8Rc3DVC7E2SsFHVPRIUSdISzFd84h/aVGrEbrY9XvT1IaBd
xTjO/oufsgpYlyf1xMVmghrGn23GmExrmixo0wrcgLQMv4w/1gOGY20XqcHHVBXz
yHOVX0JmuOyg+ul93kbnpwW1Z2ANlCBw8smm0O8qcWxl5QX96nPu97ktnNvy9EhA
LFdMQ4VEPnvquhsNblZXjx5cNe1RaPOCGRfopcLetyifLsIVVPIzAOVa4HG8WKAy
jRO3EKdLnEBEsEQ40ZpiOMdD5L4cSJ0XywQUfOl78pU/geXhyE+N+ep0clVHvGOI
iXsHuE7UIg74rv+oba0BPeZ6xriKJDDFjk2EmcxNLlUnlB1SQyk1/dUF2lel7YCM
fSG8nZssPXRBETVYqxuSnC6wF+u+tdUI6L3cY5t/mePh0X8f0D30ra1DxStz4YEh
+hkfrKV47qkJUFvIaIxLoPkIUl2fibdx90flYLFf9AA6zrP+69R2WCP0iGVlDpte
5TL9nJwr069dTNG0TMB2Saeea65co9IZz3P2B6waPrXqcMtKNc1VXHq/04v5Vkz+
XTI4yIN5DWnKGfBJFm0YUwwWaoDOrn0l6zCO+NBAPgLxkPdio3sUKJsRznAGvcEJ
Mb4MIzKUDK4MzFbohdS4PCuk6UoV43ql/vKP26bLctsc5X09o2GX3hxezLoiZtWG
dVc04aSGI+4OQ761Coswp1ltrWA+lZjPylbasaeljcrISBTjfkUbum66lLznDdIQ
9VxbiW81fCBnnd9l+u29nQrvOB+x99TXKlAl8yOeXX6mAe3erxZ7RN/+frsZ+9Za
3Buau3Dp2szoGFAn+KaBctvF71VqtrYhZGFWtxwRLx2nmVB0c2eNDcaO7ozIzZX7
upkHnBc9Zhgetr5keBXNiMgjpAzcRQckmRENRd45PXTW3oh6TMqyf66wL77VneBv
Fsi/+Ka3mKY4d3EI0ud9c52u6DXaIV7/KwVyxinu/IufXxvmI2k9lOeigrueLO4I
60/jTbfDfe5fTJhAflusEJW7azlF+r5Dr+k78V6GS9K1p6zzWzY5ZC0g9kUXi+DM
TfhU9CacxcWWPT+nIyULOmJi3uH+Q+rFMJTtYMtX+7gPpDT91Wi4bG7pcbdJC1/Y
DHqnaQ5F7ToGdSM3W1720DYc1mt/vSVXAAnwKFECN2PLCsBH3XKJJdYgGX6V/nos
qzsk3PklVjznxZC9OijxEATO3QRe4PzpVqIP0NB8KSCcr2R/x8Dz5w8dBm4iB02q
OgSWoS8k1wkeYPJlYsFGno1/004hmV6zKb6gF3WBpr2DaZSudVEowuFwI4td/WsI
0w4qpMv/CiV6bxdJgU1SHe/whn9JA9LorFjHHhCIZUnxqnc6PsM4MgiBcEmsSOIg
xfsPRKOyMHrMVjvK/SZqQ21dXMPvuVRN9WZnf5qnQjiGk7dPQqUzwQ/bjmRCIJYv
W8Y+yho0O73Q5BAT70dRqet5DOKmxCE97rMjXxxCAaocvn9wGONEc7rETSxLq0fA
qdPAEP1PmEKzTfzMdqRZrrlBdtCSmHgo+o70n28REzdmlAMM2mwguHWVK2rU04xA
RDF6maDqMWbcQi15dLaJcPjr6xqnpgKkd403/JzH2pMfMeudJUnu5r1eOS5RUjDs
uwQzFn+2wEXcTZ1Yu28BPEZtMlQFx4DdS7qcECNhPiC/ztozxQHo+QxCMjXks9sr
k0+8/tjBhQNglngDQ8aJFuH0crnP7q8fBWWBiOjjDva2ZafEBpulVnc46mLovGik
wTmlrz0tREZgKE58j6Is4MBf94JBzRaZ00kr3SGQCtSMzh8EZlfw8RSnUs0Cb/fN
QYYyXe1IZry7wIvr6C/skj/BMEA/LGPDjvN5JMX/zVUibuFqN0Ivhsq7vDPhBXhi
4kat3y6lUf31SJz/bpS3C+jGoRkh/b2EOqM7wuq13RVJEh6HhslCM18z/VbticYz
XhWyHcjq84EZT1UbFS6rzTtXtSzwVxHM137Lkul0YrVnCuFhc2eabymqWFACe1x0
nERXPrAd/SEHW8xkhGMK+eY/ZsgIWlsZnbOYpl60vd2riZ8mTuB8aNvVr5lABdZT
VUSABEwOxbV9c2FH7Jps8w5LL4hH6MFEpXBR+ZmP94Ua4RJft/0lNI7oO/Oke5F5
7PRBI5QZxzEwR1I3HkkCFP3nl7ITLQbB6gKXUCZRI/pdSSTv9+ewnqco1Y6ToE/p
ps3BTCiTjRotAkk9GOlprdYu4i1lwnNHyg+0Q7NgrpmtOuflGWDG50PXHqz4P08g
qbvbivAOh2WLy/99LmXpRjReInUjSIZ6rkMxXnSUp/H0qNDIsuNikFOUxQeXksOF
Z0VwhDzml8O70TBxF+iDsgwrUVeGAhi4og/v+KZjnCdePvetad7LtvxrefP+MKY6
uU8bYmFQds1d4DWIHMvDC0fA0AL+v9rKAtD4vbU8v8Y5BOdhtPmwgJ1AzeX+ErwE
VMsDweu34myi59CDaRNlPg+bF8mz5kZWLxsh7u/QNzsgVL0eZZw5j1s72IaEH28r
wFwCA2DcK0I6R9IRnYd7We6zr94dQH5a4z3LaTShM1qOHjlNtgsgc+zeOAHXlLco
jduD4c9y+84QOMV6feOqDdf/qeYLONpu14iPib2vLQ60opeV/xIC1qI/PzYEJTnE
71hsj5qsdtNh/rxg3E/f2bt4G9ruTMib13yqx+c2RziBOAVKqLEtHlrCd5Jy+HrH
tZpzVkLwPTEgHjwj6HSSO9Px+FGkN0VZq8cpvev2p95BXJbmEDUfrnOLuX/UJZbR
GhQR8UfnXvGmv1UuzLJTW73WFnHQA8m/o+i4eYPz9Hi1o6EzSmh8Hi3ksrKjwLES
2gXuNM27unsWKQYQQ4zSAG6DMXEl3FKi301PzYtmsBCwCYylEGdGzkPRqyMQymAk
/A6H0bUyeBKGGaFDdbC6c/HDPrLEPQtdcVlLqWmSSF+lTpQs1RLsCqm3V4WsRICi
xRa8NNUVLOUwdpEAJ3CWHJ+70nU6lDOVTn83XB8jTpU3GH+0LDh0MEUU1K30lMi3
jQnHIfYs4iO+G91J1YZyLofSEKywAx8rJI2xsCQRiTu+JGY5Xw3G8CDs0DrZE5Sp
V/z7d6gOL0zDpiW6FiiA911JpD340HOPgxig9dZ6f0kUAJj8o1SsucDMr8/b/jpX
OJjk7dklOYdSD0Pm4MJbTfH17tEyk9F8kuB/OXdgHouXyT4Emof5vJV/wVfv0PfY
Wihu9ojZRam6ldGNd7cNwRmlzYlbVHz0HqcCo5187k18+2Qmi0QKq9gfKjCxD5dK
5w8PeVBRx3OKkQnYoGMxMFcVNu8aCFsRkZPy0h9dnYk7m0b6fNVL9dk0GiCRfFux
0ULpcaw6k2ziK/EiZmHBp7GOM/4qZYVvrajz1pcNZ4W6BByBuE3mAgA8futEBE63
7gYuHzRY/8dZBJ8T8bMUti1mYzMrYPiWYmP8Eg0SCnUTpJ6snjsghDv+3k7Z6wb+
4hyVmpdOvnreQBkS3D8mxEldehMAi/bD9HAwuvFuLEHAVOELSuN44oxHi2Xe/mMp
/TBv0ntM/ZBIohAMa2kDUFKxNM8khB8v5amw330u/syrjhQoTUpzrZdXEv2w1gXz
ffTZ2GiVUS5HYCWS7auWjdsn3QZeBISCSZfUaF3W5a3ezM2G7GTaFcTIR6yNGfBF
m/zBXZ3gGy2v5NNpYnjwEahC7pQDFjcwW+9ZDkgVYVAaPV+vQOIZAnnLbCC7WzNP
GYxauJLjTBuVQ9JScRysfTuwuEKn24zSjTbl/Xq4Z77hDP80yahZ26biGYP4J+rr
VliM2yIIM2b879NU4EVvEslv3T/NPPqmAclEgAZ+5hpPMsdbEJAH16e5hZRlajYy
6EuwTa8HRgYYxDZ6pAsTHvLSbcAQ7gk+seaw2Oztkf/940Bhiq5hsF0MPQzsnxF5
mo6FwIxAJ/+nFnVHEGY6NdifKj8SqgSMTEQXQNczj8M6oAL+69kLcM81bken3CgR
XQ39Gaw7ty5RaF4SGz9oPPRxDmqk8U0xKJCNIdJlNTiLB5F6Fv4cIZ5Njiat5kzd
c/E0DFni1O54AmCZ9QfXAeIF73RnJMao3JWs0dxGda0iueR0dwhMI01ss5++WDAQ
8WfibXiOI0YMWuS/xPzKUdvCeDK4+cU8fv4yUPpeFEZ4qvF+LSSc1NK2a9F5pBiE
N38fKtSmbeqyLRECesR3qoio7Uk7gjpS/buG589DCUSeU5y/p6eLpQeIwhRa1HOZ
Ka801UDcrDHOtKHUf/MhhOW59VQcQAKL8Sb9gPPcboioWphBXBSFM512S/SrZY9G
jUOhdqvyo90YuJKxRL2QxM4uQBDjC1V7SsfYtiPsmEDkVVMgX2yifz6osi0imO/Q
/JgPUIDgubwWxlQ8Mwqekh8nxQyqD1FGSHALPqai1nHExd0UlGxTt467IJ9v2Adl
BVfP1VQ5g1aHGKGU3joXGocrwfrnyWW5pIOK+iyO7VxVPle+Ew/ieTvOtHR3cuWL
ytl2f7KXgd1EvPqBQin7PbV7nSVKS3wB6KSRjZa3xbTX4SdKKzrzyhqBPco3QlPM
F+MW9OEjb0IahMX5AFlnSz9q6Q9fOgh3SAtbhbqtCfeKCZqTKn7dur1EGWsr52Xu
ywb7YYpmFlroIk8zhrB3z479sVd8qjdcGjQcxCrefdeeNs7hzdyaH1OMFdd3iKGI
eQrerB/j2QgFC1GRVDfvyLyRZJebtLm7fGUBMK69DJDdHfm2AopZNwdYvOl2juOR
SjH/fctiNZnoCz7o/LQPlcuYTF9vJXhWgglngCP+QRTBvAQQYD+9gbK59cuoEeOp
mWxkRbn7PzXXvBHhq4CIJOSwIpfe2d50KVFP7aEV6kNcM2gBciOw7SGtrzpjA1uD
ym5tUmeV82lJ9XB++X1KgcCrwb9cRb+n3dlc42HuAP5vRj2uRQpeCMKtTGZc7xXr
T20OAyc4FuyGnwbQlx/6NfJ48GKHp5czRwnqs8UjCh41SFu+ev7uAmW1FM1y4FKA
SjE84E8isgIAY2O5wLvWhNKwVaN3PfihCqeHWo2gtEOtaMVyONwMdorXihOx4ATi
BrEcGd1j7SC9zJWfbbH/0yHzOjIwWEQNI3bdRGBqGPpTtav6szin3jZEoS156l07
6Eb2Zqiz6FrJEX0Q+KVueDtW2SS9y976i+H/CSH/Qelf/6ZFSDWvpna/Ey+cF+Xq
TJ7x2x+/YPMrFirPxw37kzpYgxE1XELcQtSgvzFzmXhvrW3SsGfCFJpQHIkzA5s5
GmBfpJg3aecArUT3UPYkJ2D6+i436pK3FmSI4Wrn3qkUSk1LD8UbJ3DCm0zNBsTb
QPH/Hv6bSG8IGNOYx43hFKmq4U5BzUhzf/LsW8JIABW8Rfg2T94GpOgdxDjC8iGe
eTZseXgOD4MY9aH7p5cj1Ab1cbn2/ZvheFYc6jTJV3G7VXnzt7Vrbi5QjNhkoUB9
Bwlo+D5Q25dlP3lqQDNu+1qk7kci6VWETycVIn7YrNPtJSRPMuuPIZSXpYFs3TlT
gd3Ddt7Nd5IFlWBHCIZUO/1UeGVS2LLptyVbOlkhVSXvZj6qB62QozO0WTxd1LPl
OkUbH4V0B9g85V/jx72SAqpFcsO0wRIsghPV7LQoJc6FXRui7GTYtu0Wy6rmlfwG
nnmvbRapSLKtDGVZzZRShqhL44yRKOt8Pdf4Fn37qRayoysTixuzaapg1lwQCvUU
SdDVbzJJbObvgemTYqSqIUSIgdigOIEKbZWVkM0sv1t7mQdPgwQddD5jg9mkN4MC
HI0OHTerOGa5REPYO64Nrr+P712hrZyapA4ztAjeeUty4oWcmtQr0odOctcxG/Fy
AI3sTChLQRlEW/7dwMFkmrUxjtJjKZOv2b7l6UcqBMDDuukl3eIEcOqqtavIQh8G
ef5qlW/UkZU9vkfwH6JQLq7wa2e317R++0MY+OvTT8Pdz2TudDUBPp9Sa9HeOFe7
+22SvpKMz2sFzzQzH91QyB58r78PKMoqHsoBLH497qmuSDKqu2pnCk1DbtYrYM88
4KAA7ndrIojw0u3YyQwITXfMkGAORMucniB54lPxLsiI9zfCaDSauQqPUclzMg2w
l5gvpOpfiFLInlx97i6pFjWlGGDskhYM1eGOrKt9WZ38x/i9Ixi1aTSsoEqamO/l
2np5m+Bq1gAyHNcaTgDW169/TyZK9QiFdjoq3Q2Ee1L+MWwPKoWbH9hZz325+LsC
Uuof2hfxT/iBsNaI9Q4oiL4r/J2Na4Ds7JUHQbr1wS2OP2GvjK4OKadQTn9yxiJq
QYaRRNCzIrcro5TNQjDVFjXEimThUQcJBp2OgyMIVB+0nMgnA/yKTgSX5trLGG3T
4Ril0TTUFZPW9OYCNqg000BrFMraNbdEgYqSs9kxzOi6Z32+I1EIJYa1CkjunwtK
1vxhfDnQ1vMNQddy27EHI85FcMyHkE5DfEZeAqMrssyZse1S3e8azL6v1QlPElBU
Rmr18vabtTQxEOdBWl1MhzpFk54oVVsdWgfuq/2k/33EWVHcSX3eCWNCAf9WKkq2
LJKMdg8deqH+uFW7rqPMbHcQULSfbAZ4JSMOVho28UqIaZudgpOF3/pJXQ7Ge1zS
6Ah/aVt2ineGmOHwIFM6v1pvmCzN+AiAoTAp4Dn1EAAvuvkdbozmryvWmxoNm04y
Bwhxr2SXHtoOc4Jtkho9LG16NydCGp/rk8wz9niQX8l33g5ImcMCM8S9umaN1e/p
hz5tvANxWfYzecNIA+TSTTgR/kp34Tt/Q1KOYuCVv1w9UsjhsCcJl74aL+L7dcx3
A77xu15PU3tTaCWHb3hJ/fjWJqlf2DVjdIJzOXGFjd6HETJO63dXArv/JUdIrBni
KEwEkgeOn2IPDNg5B6Zgt8vf0wLFko2RHfMVitsdik+LYkl8HJR/RRy9vgg2NBVM
p39hXRaQll3e6c2hF+na3e6+u7VHp7MSMgXIeND5NCMIZYHMLfgZAU/ZqEAB0aVn
UwySR5pa03fMWQp3TbbNQrPZdmLq+30bXLTGYWO3O21/halYgByghZL3W4ssvg1l
kNoKFBqsaH6iYoJEF7uTFj/TtGNoq4/LBG4rwKlRKxKh+rC0KukMfBmfllr/dkJD
C08OG7Hu0COIuMldCqNLufiChBw7r5Mt9hBkezg3AR/1Y6gzVi+EFoyNhXYhAa6P
k92mJ83QtQ9pdQo+J8bunxbmDM05j9gv4R5s/x3cpLHqZ5KcpaRfvRI4RGVrnsa8
29/dkH3gZN1OhyO7xgZKwQUufBYZUl+87rD4dyMDnhTd+12EqAQE895MIUmksPjx
NQVhjXw6hUv/s7Noyhd4hhJbHkwPEFgQVjdrh7FzIbstjq5Z8DcBaeasHd3hE3qL
QBD7zVvIvgGlTP3996wd37QP6Usc6VQ5hIsXUEyIbM2p/H7+IGtXfzHEAAArGVKX
A7jkl99DM/gx/zkIBsZnqLhKUkfRX1nzxZZjvMYmqEVqS7KqwgK/2r0wc65v5Idh
eOGOMQZ665gjlmqW2zAOq0e3RgPn6VR/5uuFMPVzA89/QLAZVLtSuBShBVNqLQJ3
FKQgxe0WzOMFuZLRM4yhXGuh2sH9TeXuO5UPrl6viFvUbhuwrqOtoYx/C76eh0qh
p0oNUBSLc/VEq4UO2oLflLmu60lpG3eRKE53E1dkTgGCrGC/pqW+DA2U1BzXVjQj
I7I8W8aJotLbGNjTcz8iAx/AGG02kdTPZZq1Mf8QgDg36nHSjugmui2n2XF8kDJm
jrS9Erko8FErF7CUxmPu9C9uZBR1w2kg/6srax6f58uK5/WfykafMm/O7tjWLioj
38F3LhG0PF1/YWdNlvSta/JOjJeBUloS7LSx9xoreFpfN+c4qPS5wYipGHf+Okcm
bjyjaKia6nDJ7VZkUKW4HfS1e3DqWoRjDffZUmY1BiMxXvIedQAyndUEaUu8ai3x
qrBEHVmt8uf0Qk+Ukz6nBdtmN67XpvbiqkjiR7q9lDumlKUjgXGpnolnqFfq5+ZR
I9NaWSLW36ZW7wqKrHNVmy5CXyh5AyJRwyAQj2kwyHYy2gydsuG3bSxsP57PsZIk
VPGytd8WyZ2zzf2AOhHGToja4dEoDeojaV4u/K1nv4lAQv9QByz/pmD8p5SevJ8Z
yxlJ7NCyFSMTef28nP+43EIncjfINQNrE/D/bm8r5Ji0x2/m7J1aD91NdWCwpDpn
Wy6mzv4sUUtfEqtg8sBXxLrWpoUXWSLHRmM3PZRlzjRwAmmHTdhyIzD1wD/AEDAm
CKqmD9rNPOHM/4y5+TVpmXZXtOJEPg4pqy5yLA9ofM98loaiyx1VaAx2B85nEL2A
kD8HzmzXFUY4iHk0v4SocjkkeC5tSVH4B3Hz01rY9zc3eaecDX6+DmIndAXCvnUs
t8fI8xn5164nk7LCez6Ax2LXG2zBveWthYu3yKIbP34cBa2qz4ZPF57BPWdYQzfR
okIfnGEmDUjZbwKANluRPvvF7nPTh1vO21OZIrYdhNZ+7gsP+VJPM/r78tyocXWk
NknGJockVGefRiHBYFIxMF9dMnsE0zpWesMM5p+Ce+OjsMwC8vSeGS1APN7oXz0X
cIK10dGLXCrvaUCBDYhfTNhxaojqMg3LKtbbAto3xoe/Au+SGPe2MYMMBnOSOhST
lcPCTQcsEuoH27sO8/cADT68Dd/q57ISc37vHvd/r6JisOy0u8uy4X17PZd2RQxj
VlbDnRamIHd/e4J1BjHk8o1INifYs3XyqEyghDsO20IVTCfIkh7Ci387IPmLSZuo
vXuCjiHqrQeXzFJkeFh5dmSJb7ptc+I4F1JOwaS2/Dg1Kl6RrMl2gXMkfbPfjV7E
yaX26OA4XRt2RHHdFIOCfneprTeJebFpEPuqc+a4x97scHcaa4H8h9BY1GZ3+fUP
fQFnsi0pZfBQeK9UeHw7mD5gRnqGsMipVytIPcutqV8L8MNl8HeyqLcUIVAI4qRA
+8bxp8VxPrC10v4Q4njiwbm+blD3T9GyYoLznVdCbUvbqVLsYMMUS2NZDG0MFgpf
n1YyLdRwRisevwiHTCZMvK55HPeORxG/yhkFKjrYKfvTNi/Uvbmqdkoqecwb/GSD
tVRnGNuOH/kPpq2rxe25KBh385DRZCxbYJkkqa86oG394/3OsnjDyHRgQ0IvujA2
MkiSyfy1YgVDk56ShrTEWaekTYMtRmmYWijNssDI4h+EbJOsmW1ibSHU/jYTDu81
UVDO2yUmqcu1dGW8EOpqD97a4oFcVD8OrVMtXJGJol5RZDK3J04yGRrLHh7EC4Z2
Eb5TJMF8xwVw8mcJ1Z8LbYoWN3lVHC2/Jsnoy9OiABIYXK8nwJFzZWdrQvhIdnwO
K2tWtBis3BqDmmWZ3IZ2SeRjBdR4LfZMZl2uAzwNk2zyntIdOkHjG1iLIEcp3ZzW
Ev3J3xiGxn868EpU5zinXTvxcFALyTs72ozPS+4P8P4AIxMYzSSve9rWlX/d2QKU
DUqB9SHddPdsM7QfPerI4O4NQPX72AoxPEOVLfL2+uFVofhykCjvpYWmMFwlqeiF
4C8CaVFVlob7BXgtRDwQAY5HA2zc6LHv/c8gm+0qfhw6r2pfTWwAPHQpSSyFRRlZ
lF4zQDrt/DYYtpPLCrkei5Io9o9Gdel/FU/p8TjnvlFeGczt3J/yHABJWW3fPd65
VkofAly71iLQnD0NXpZTd/xBlnGQDqhW9qEbnWH23XsjLmSUSDMiUpglh/iw5VmV
6N64vZ5egA222XL6cvFANK73J1gvbxnhbjBwZOxGeQX0qjHzlvO+1+ZPF9Mlj++M
YVRYOqsEgOeMOWI4CfsYBr4JpOd83AviTwMhsL6Aa9h3ym/IhIWMlQqyuAM4Jq+X
dE40NR0gd0HqtNZaZSfK0pR8Q18CATrELJvArSdL6K1Cwl4HrUErW2E2cN2HQml5
AFD2uowXjBqIRIrsexbNOEYNb7nhDYSbJtOvg6BvqWB7BfpuLRdjeV/HzjGvzoPf
Hzzaq8THsm2FF5F2PMWyT9jdEoR9WmYmY9giV2rE6wRLGeb4NeFwfJvg4XmbDABt
YDSX4XgVJsvoPO+WSMDNR49jiaOeKK6/lpUnYTDNRFlmwLPyRSK+wvxTiEDDtB7c
WxDqK1ogZ9NiPVDJTgOFqWlaeuyL3cvGC3ishGQm9I05rgoMpz7TjTgyfpbubveA
j/Wu3R4gnLDQfWTSj5hyLO/cHq6aIq+I8rNspe8/7HQa4Lzol2CUSdHn+zfZcLCj
upOcFyZWBR12XrMGnE4ISFTiW37vLeFcJsy7AdbGHBCF6jMwgL9DwTPkDPFKi8zj
V4YzpW9MieDpjO0O1IzDdsM5wTmXMH9rlqHs4obQe0O9Mde5K4FztVW99dvfC0bX
VMrpNtr8SEl5leK7zaEp46RwhMg9dPKSn2YOk+NlnxR0K459+djbEgQQL9M2Afqu
QWmBSwI6OsDJwxLPkNG5eZGFzI1dj27N3i6x1EMevjwFzXUoF87zja5yiVrZ7XA4
m6fNliKfB8xVMU6iYl1reYD5DI2mOHyT2jmhOHi/7lU4cgFxhgC+3H+UiGnndG+e
RxTRz0TSx25puLWijOTRYl20D4hBbYXWLmT7BQ3BISHSl2oxLGaB2AgmYtTKfKlP
FQkjNpX7LxqS1bD/avqJtAcUr0YJsxE33AxIcxROFTXnKZUnsULAQ+dXj9GiSCjH
+crge1Xb6NICqGKpUVjsWEWBkG3b+pTK7QgXjecdDXk4p+gsXnV6ud8irUEdQ45A
qoUHUj6gI6IW2FDTtBNcuoSXwJ/3tSKOKLUR3VXd/BZ9U+a6MfeC26V+5VW0twR3
0/7y9EtU6LMl/OaLWQptUBXtuDFak7QTX01+BVbHSXbB+RGUbVipGeocBgmE/d6s
Z7xz2umk7UcrmLIKmWU/GIsCOe3vyzda713sfUpW9i0yYlQWAUVaeRkpSscrrgYk
61vsPe4T6eRyiXXf9z1oVrvK8o5j6JPurht2DbQpQSekd0sYzu3RZNLd9Gb2lW2S
C9m67dQe+AgMJ+GREQMzca+xbhCASH/BCpkZ0CgiFgVq98/xsc3gMTIY8xqIRvts
8GLLjZT+1Qq8ebQjol2GVQ5bZVnxmbyWOMEhdCZAW8zPnhQdU8HtHzOXEyD2Y8im
fX/CMnzg5r2qT77r7pZKBQbrP8zArxRfFWmS9Up4G3rHANp+4IEem0b7VO9qxauu
XWBPR85D5VhkGYNqQKid+y+I6AZdl5xDIrnfR7nh9fK/FJ3dm8iITHQSqMnp5GYG
2KZ+oBkCfQ9AKXuKzwTI/PHvkbhBrUY7UNwjW8EovRGwhegBojBw1lGhPtQajyLL
E2ofDQSgJU1/X2w/tOfqigGTA4Q/Mbg6E2iWjgG0SYmMynqTYYdmJK85LUiQwHqG
+XRIWGEFzkKDikut36gkV9vZDXiVezeJ1N5FYF4K4vBkulsiGgyrfIcpY+J2efJ5
gKgdiqRcFLqB/Fak1XiIXwZBCUfAtMjx4To+6cStyYsd1bilLLnTLZ9glXhHAoRL
snGYP8azGOpbJDjyzGK6uUaC1aFMGc1b1zeQyBp41RvaL08BbTP9nI6cAISvTytR
IUW6gvd8cEQQ+J1obGeZx7GJizST4Ss5sqa0Io5GpQFWQazP1gpuQZq/OmchvnMF
SoftCQJ43UhLoYNF5tsZKAuh9A+v0GpsljTTRyEB7zCaQGC5XogR7Z2kjHJrj1ij
QyRXFQRnrg+vOqqx84OG3xE1VZouAhnwD6gco8LkddL+8SFbpjiskhKWKgCBVyCG
GqBJMXkl9lfKJzGBUVq5tOUtwcrELsTyhrxWZHmpccbysmFdpMH9ibqewy75uQVb
YXBgjLtZmDTs7XqWDSVJ0UeTYeZrAd5BFZ3dx9HMY2kWeBibUMcPX+hX056bqgGC
T3P9rAJ767bKwimPcNLyjZmfGbNr/c3zkk6X6xo+teq5p/BLOXKx3Y2cL1F1mc7U
UTpKtXpZzFx3eW3jbfRl5XXWAG0XIcZqXvdtbDVUGAgD1G/cVgJ798D2PQS7zaH2
Xe+Od4rEL5od0fmnq8qMwKUIDnPXwQrL4hu890HuhOH5SZWRHwl3HS2ORRxiV+G2
r0neU2olYtPctkAIGdpRxOeT9SvZaxi34OQxrYkcBLSBVcZKDhheR33ImB5MtRP2
V9+FUF3g6U41XYowroGYxBuBt0tYhmUJFKVyYOO+2+LI0sJexkCdyta8qTcUoILQ
ETgvsQaDREfcidLlc1wrGhTysR9G4+w+ftLBaRExXaqVjSemEcxMrbQj2mrFEcT8
7/Lvv6BQbOUfN80S0erLhekrZ9fYRC1+M1R/nNCsZ8xqk8zhGeMusxkgJDWmF4pr
CqC99IUdDEbrbtTt1nUApZUALAL3RbkRUQPfc0HRwsJ9La28pit8ovKebnl32FLn
o8ZC6qbzYqLhvgOCuweIn+NLXVduUPNV6+uzVYl/lQDDEir+pjGEKfk3jhnGvgpQ
bf9D8i7hyVsOS1LN21qqMPxEGQ+LfAhVKWinTujyoECyvtadMjphBCC2+aHtXKsk
5Ndyo3fCJhk5NcWchwb0MLHFIbpqcSUPA2FKT6YbLC2lnfjXHcfBQY387YqgmkJC
i5g6dR4YHbfUbHVWNpclFy/rswtbY3Ko4rDVDirNF4KPAGhttN2GrMj3YuXwWV+v
sKV02oYGDQmA4BbBK6iJ64MRVBX1m6SnWlWh76dAde/WU7UWloAyUorpr9REnK0M
acaphknCorY2iJuwyjs7jU3S2uEhqdRjnHLPZqAuprmGqIg4AUh+ZdFKLLUc3N0j
ARJipwDdK7UQKLJWrbdeiW6XAEKE9LhYgGWb6hdF1duJBLuba0Ac2rwDquOMthQx
YwWuwNyYD+GhzVz+FNO8bMPS5eLjxk/+zRxeHJAJ9/ge578FWIZg57D1J4Tj2Sy7
gvsnlfml+GZjiClIR+76AzmUQxebuij3RUlUAMHctE78XXZ/BBFe7EoDdSRapvAt
VhqgyD+Ly2iETExU/4XwkSelFhbAGlQAHOvqfVtFYtmZpNSAJeTJzUTozfoWTLQ+
/FDRwMnZbMD1u2IrY253Kz10VWWGAh06uTdWtvfV5Sf8WMfZNqHyR+pmTtfZBhSU
cSBTFOt0jmZSsLotrHvsYP7srUD3V3k/vV+N1gs9yz5QJrr/g4H0GwhLYrr/jfFK
kG83URipsXsYvAAqXttNtAzv60SfNNCpkHAeC6Xh6qDtoWZd++4H6ex5eY4lKlhX
4zAviBAF+Br5I3alR/QOFSyUV9zwJ+CaKDhEnGABEAPYOA/Q4BEvFABotMAhhEDX
QydXDjXsDQN2BOiiAA+H5g7DGnfekvQtf+YO0FMscoe+7JRMq5v1EnmnNxEU5HNn
+DuYCqNG9usMXy5X7hydOQJ4ogJalE4yPwD5uPavYDFL5faDwdFeq7LZSGF/9ZYc
as7VtpEBuHvs6Ha1vhrLAglmkNEIPBGuEhyOxph8upVaq3pgDzKhbdSVJj7lScqh
EEU2eSDCwCm8YAlhgqwI4OsWs/tPTSxoBfcEQ6bwpHYiN91SHRo4WVuqT5Wb1jrV
nqvt3Qa84sc9C29y1IjpVozm3Noy/i0GRc3lmaDMubEGYXiI+gI8ub/C39dbYey4
yxZ4hNVYBrzjZPZSjT1AavujA5ZpSbwZV84n39VUR5z1jzzRMaT044irpZMrbpSv
QwFUeVHjlo2PJF20TVDvCs+PZzWgJqkP2Yo9ifHsC4d7UWPw0ThDL330axeRcSaA
JNXW4BLy0sHVX4Fj7tpMdWNiewJuoqNVG/J2OLItX0C8xxyikgPRRh9YMeOIQxoQ
6W/u3Skw23rC9Jf15qN9x8hJDOOU2EefsSqZAEaTFYYqsiiE/F7xSN+PlDV1CMkY
7yALpdRgqTlPgi72zCPHg8x6yw9cXDunB3lAa2dq5luGY+HwOJGBekMX5UVi9d+T
pUWQtwilvulXFm7j+GtlDXteMJgOb/xYrn6IAS0ENuNxgBZCh0L5Xih+m5TJNfFN
IxBEgdgOqbFPCjcC8LikRU0xoHGJniYopOTZ5Z5lW1UVlCmhjfRDcWGz2ivkFiKh
FlEXre9rMnjA4dbu6X3KSNLE3yVOP805KlvS4j2md1z12ex8/h9qu9hvFs/NBJ13
M1l7gdmVq3qy4FTy5LIpGqOueorU6GQpctYXWg+qqIE9hUD61BQSjdrrxXhETX/L
E0MGDPNcPOeUeAW59elGTDCJUz4K6HRQX66VqtoI6Jp8K8hdnajZZ8i4LVv7FOVh
FHV4NaN3l90eFaFo9nF+mnrw4g9MmsDt2xVZq4FAcx6GWMzbERNLx1LCPKy3FPVf
Z8amWs7907PY/U4Ms8hzqW5TOjy8Ys2QnPVWBHdYyIcvWiwXAVbqT4o9XSSjFBcD
mZsoBNLEj0VdRobxT1BBksHjsQElG/LLj8LFGerbAvCU31uU3gZd4wws7rVow2BA
qUHTukhvg0GpsvAIyZIaZzSROnsL07bwO4bBll6KPP8UDLhuo/pwkO1987k2/L4T
hVuJLoDKeR6CDAKZv3iWxs6bkVhjdY8y+MVGN/BKiK8v9OOuxhUhHMXu6mCy711f
IdCfqvIJ0nhkpKKZI6sK1UrWg0Uw5ERg1uvoA1xsFv6Ma6CknrMyDy3JfWrsC1e7
jjIXX/QQSD2AAMb6ipVnj5V/kpvhBORbRcD9G0T9OCQYr8txEOY5T8oGXxS/p0Br
aOCsIh//a0ajkL037wrT84ebluwi0pE3vacM1xYT70YxbencA9e1tCnQnSQeInCu
+FttbUiEeNJKgX41ckZfIR7yqvEkIuAHdBqRKcboMmdWt3jJaQjehgDxeJGZQXVc
u7+clFnH2SxvsfsIlZRO4AHfSXmv77cfKrTWycpUdeD/kxJ0aPyuJjbC07AOEYkW
fDPCvXuv7WYersmURhNuu2KrkWcDYNzRDUuOONIcz6ayIh2VtoVXtURPnf6vppxV
odBWgXYDRPFXtp5G+2T1IJ2OCf2Qm7sz9qVEQw7/Ctnc82IemI9sc91QjKdN5vxh
Rf21IFrKv1jd0+MixvzHDwE+ZgUFNnQIrDzCuE9GjFY5G43aleztRcjDMR/bI9O2
qDkoTadJqGIGCIAjAP88lAoEtDyummph/mliBDjeQ4XMlRHyxxOEgLvPApkNPVrl
hun2jW0OySdzKZRTxerFSuNhT76ZFoZd32ccgAvl/xXXP02V4E74ijeBuxSOnZ3y
NHKJblBrmb9wAfQh+UNCkjXqcftB0G5yMltSVhEmDFgcM70tsp29EBLknJyW3oZg
SBk5DO7AdfjTt85Vt8SBJkwFeK4ZzTo3bNoKDiTxjYiKGYOcasFT4CTw3DdxcU6T
wR7sJNiA0fp3a2YWeAeU1EAkj6ZmvQXypHGdcsfr5rNzK8mcfgkbMpmHnGnEs/Jj
F+IanaThWSsS+JmxTIZSMuv8MG4tu/O8gOJMGYUGLiqmiVNItS5eGs5vuwH7ixRz
bFZ6g1F5pLmMQb7ssE2EomJO5vezWfqyIriVx7z1xvyseSzv9eYXX/mAjOKdZMyN
kFblS9kdGajXjAF10L6BNSKEv+1t2K+mz415Sax5US3mrNaKWLlx9i8K1CJVB0xU
Jo53ig9eYwr9povtT6XhEfiFPS3CViV2cpt/TAnZuI2m89qfAgdcg3hkdsnlgRmX
FMEdLoTi5OZb1WX1/DWHkeO0vVRFph4AjYfE6QDifG8xoD8p0wsz1o7R7u8w4/UV
mkOgL0/l/vpqoPQ6rvNrVsLiyKdTO4/xxFBxhHG8V6GYbJCQZHRs8O1p5PSlpDKg
UjSKx1aWp2HibKvpc5Or7+dqI0ayCe5qOjp3LRLXfqwD9n2n+M+zlRWF0g62HHsN
GpOcqO7PCC7oUBkehcsfOnjK03TFoREcXxB2/t0ION0wyYImjdLbI+Kw3Cv4Q992
A8H/pbKlXGjgwpDxGcSBntI9mj2JQd9Kefg1v25qdkqjuHOR95fSs7I3LLbi3JYC
BsHwgWezUSbkS7a0T2n163D4yakHOgkud5774IcQ2WFcpzBonOTDHxBbnJ6zgwXP
pJscsI+rldo7hhrQfWCoLnGy3s45Bqv79J7UsEV1xBzAMC0dpN5fa9vjtXJ6TdQ3
QI1fFG6CgKtmbYtFAJEXTS3w0b/UnkCpBqn9Wns7oMBraNP1UUe/vM3PXhfEzfgZ
Q8AhraKL7jBVxWP48JqE5KjNUVPEkRBjosFTb3dlYeEJoQOaMmHDXsgTXqyrPSHb
wcnyyyav/VS1m95c25obtmJpnKoxJskgJzWNV2jN4ITObscLiu+RBE5KnmZrHQVR
C8WWFxlaCqY+1x+ZAQZAfGVX3UJv0SN/zHvB66neSmwtswhmGO1cwBvcZ+qliSIJ
JQipx/T2cLveTjiudveANOfu1fS+mbrrgY20ZlaeCt9syukcL8TWxelOFFFsiR9p
FvpTh0Mxo+mN1Ql7X4XmpO3Br7IlHN7/G7OlmETf/SqXRf/fFqX04h2+mhgazmV0
bXHR4Gk0MdweiYK8fVaDYTnbqhXeJlWfx+katUv657UOa5QQHUk/U5qY+DXKC6fI
i+NzysVfmsRxGFUAHa1FpuTf9NlWnw0KeYUU92BHfhBio4L+yDne3N1rDTNaZjbK
hPeX3l8VIu07Kidjwq1Zh6W0GkqXkFGH7i4RljepgWkGIQrkpsDQQzRaxG8pKVrE
BvIpJVMkT4PYJ9kJ8b6rbSDoRH0BsOCYOoV2M4o+vYxmjF7kqkiJUtT1XvQW7L8q
JQKS9S3d09V1p4hIfSA62MxV7bpSLX7Xb2edaADJ96JVKJmFwwYIELqMs73MT5Xu
OsvZHD7YophInHy1JPN+1aKvCPUJaaFtYxarg31+aBitR2SC1kR0I9/aDA1zzjdN
4+zD9oDkxVD8JoRnzfqxxhS8s+SAN0wvqed+C92lhaa61f54PI/Md92vLQnxjJzw
GsIcKvBEpLqGGA64YG8fhtla9qNxfJskBfS8maxo6TK31Rerrfjepm+aPHlcJWKy
S5EXPPoef32miIBjfbWvXLETsc7C1IVD+8XVXVPCMllIhMjOkInwlIFs/AI5IuEm
bCkukg6+dKyyqsok8Acw804j0MwnqEvwIPGE8qlMbAOzJkvUudF11wZJ1rx3efBB
GEQFmo1XS4p9ADx310S4FdRAeIUHwmH+XUbUdjYFVy+iwiIfx/3A7UNj17ZZDm1+
n7Fcht1Krk5KClSd2twrRfqSdBqv3UAvO/3mPhxnYX+edIpirYAJ/XXfvj6EbQoL
wWsHiZq9SgqQ/cQbFJomWrlkSqhnMRAqUi+nvHYm3fkkiWc8GdyD+8HIAaP3U2Zr
ZHjojgCVZzJ5kLNkI0VPYLe/gWpf5F3kttUqP7STD5a+ANiClEaSbrcGH8BBETqQ
/4liygMxTi0147+KV8zGd9hCb1ZcLl+5qnz4Xws5HNsETytCNbdfIwiwRWWpxutJ
zzdWhrp0wXaqEcV8NDDBxz7ZTrr8c7uneJUU10h7dt7rO/dFh1yVL+HQLCIxBCA+
B8c0DHDVKUmi2+3vgFS7+n6Lm+eAOIb+ZX2vXqzPfaSxCKjtFB7tP6eksq7d1sHg
JsKl+VhlEX5f/3Q6qKdDXyyMMlMaYoiLLERR5eQwUrJVM2IBLJt7Y7QDuj5Et8/2
ynRvMk3gmCsQR7pZVYboKZS+5Bb4JuNBTs9wDbggTcDQ1w62tQDVOeRjRSKUWxkB
aAo0NqglQEWlcZVpfe8nUy5tQduP1H3NOuqeA5z5PGpf11sVfstcwPb3Eg0LNute
7hQAuJeIFcmhg6oXiG6D+3mjSQKW0zWHk+kWeDZw76QuiXO7ip7pAI7wv7JAfK9q
UHqiRdRV+sXmfXV+FOIcNkdU20orw7D0aB1DLr9oFA9JeuMhMyzUwYjtD2SspdNf
Cybi3Dc4tpOo8LRo99i+3HMTf5QL4AQZ/PrRFTfKuqBjnRvuIp/fA6i4DEWN6TIK
8yXOaZfYUX6ykSbiaebp4tJLf4KppuVO+3h3qBGrWAnzZUPfQHm/9Q6Hlu6zzTNg
WgMPrkmrPbzYRcj0WRp+qdZUUr6mxevPALNC41nBbHwN6DKSOqZ2pVvEPLfbHoDR
658AhQurX8EUV8nP2uqg1Na0BjOAiwFJ5ltietNmZd9bQrsj/MIBIy3uWtjIPs91
PVpRTDkZT2ItymRxSEQcbynCdzx1pcJFCz3D/PNvIFTvPW3Amcs+2tQDdP6YklVu
IreRnj8OJmPCsahg4Ab4txXQjF11b/NkIke6YTeeilvdSwE+z83g7YbaszNxCinY
URR+4O9ExIHpkaiprddAHs42zX2RInArb5bA2EPLeOEdMzf2oQ6ckU8lUgEgZGhw
B3a83+6rwU1zp3GoSTAjX+oLZ5xBXoH4OypUB62hYBKAJu7Sgcs+fTz1AcqLYTTz
gg6kdKLtUZH8CK5lss2oMZc4n62buinydA7o2omz6YeLM9Wl/ki1SjmKv+7CejcY
aTN/rbXNICDIdSntgG7+XHOPa7c3UDyuAZMam/QBC4rJNwmQI9Hy3pjFU4DQ5xSG
IRg6mdvojftJtHlT3odC0JKhlOOdxBjlZMujj5/S9X4lxKnPT+TwnW9wFEi2Xk0f
KXdHTfczKX2pM2OxawiuRfhmM92OJCCHQfUuaeMMjXKgn0/jG9LCOQvLExU0ad/q
jVhh5uAII4ELYfRLU4T5JolPmhToXbcq3CyrYhiAyMvKhYwvk8WjHTgZ9sYVQQyY
Lh3DZObnJI6alxAAJUohCTJPdl96wWazNJ8+mfAANTTOSwotuY0gJDl5SteOmEq5
JPN7Gm1ipbZVplQm52Y9hgRfgrj3ey0wFqRT5yo4TIKMFadTa9UMklitm2tjkaY8
P0Jw19+P3IK0bN8pkhfIutNEJL+XauGqqsHm3t7FygOcmSMvnZFs2Tqbx229SwM5
Uald3yjd7SrIo+8nhrcDOd4bqmrISPZnYlcJGOZnZatLzzhLlo5pf6VmLMobOsMR
fC/pPrdHIL/NCZCBzcxrjCmLBSpr89bsQLh8K8+NotvawhBu++khVeQ/5hWN/y0t
ZJ5++QELr6SUd9Qp1ZbueYgxWCP4T9ScPMBFsmHveHaKbCsXFNYXJrDiM/biUqAx
/MmIHjr5GrClbQz+kUuOZmAEVAab22jkqn4OOpZ3Fs4nkZMFzOA7LZNO8slanavp
euc5OTVJVu7hrzHnmw1FMbhx7P3JVcaQBkfmLWPZSmbJ8eodlgLoVSkDGeVwJcOP
/zQzqpkrSd4DJENxX5n2RWAyLuotGTZIGhG+uJMrB3wAm/YpZ174PfveNzDNH6uW
K/nczq8o9KIbrhJYt3kEGBAsqPkNJAgeNAzeL9FCOszA0IpouSONIn+nWZuuKL3M
PNzeOZg59W83hb5dEkmZptYTrgF+72OH7JIK0iCyNFXXv8zx8Pv7ZmA4p8j3QUme
MJMubTuGQHoPO8MBWhWYMpZuKM4HWpNnjYXHzoY2w6DOJzFoXDITySE6/P8kWpH3
Q6h3bgeXLwZxQdtxzJWu/JuLXZ2lcEdBkpV3znPDplpRMCJqBJ9/h/inwks/IKXF
QkguAkLjakQsw1RpH8+5nNb16zr1yyVNm4yaYRY1ka0yKymjAxx9LQ9FGQfvY0Fx
Hf4G0qgUk/W+4d7rw8QDwvQBQLhW48KD5zjoJbW0SCDHZRLaipaqA4hhkQa7GUIG
Q924DjZxnYXXAjGav/Bq0IEbxDG20Sg/Uad+dEoYAzVsYgW47VXkwuggsqIlv8ax
0eqevSg3UP81P3SFO7aU+/8SHTTr8LncT7NlykD9l6vl5US45ZPKMLNfOH99ce50
uAY/jc2MsxBybnS8KsVoVPUoXbsYr77QUCmIK6NV1wTGPoIvVVTR7CHbDYxAXktw
0ziU4j+o+jKp0cptybDRF6Md6PC3OCiNG396OMVMYxDF8d6UIHIGTs/RlfTmJxfK
AzOeOwzFBpmOoYqRM8/eVpIm+RScLUf+8YRim4C1jrwPTINE8n3jHitFTCaeQEt1
+9Sxcqp53MHX23m6QtLXMAR7wDU4kuSFj0kPvv88p73FUlhOUXKY2c8KFXnlFLV8
Xhse8wEBfiGA4dAoJynsbGCUB5zJCy74t0RKyxa9Us9K2nUkVJmPqBv/WuERCElu
tzlG3SBdR5KLiuWzPn5hlSQNIMzs5mI3MATkUIW8qI8/DWIGE1820A4/V06/PIY4
4Zsxumou45CgNGZuSiahs05laSoMsjbUIzMDe7To4KgU+olx42QSNwhQoP+VU/Er
5kAlQ4BmXmyGhpXRcixKJjp2MHv/ihMHWHibaSf9+ypYQ8CZom4GZBGmAt7AOGYh
AS1fOCDdJSasFeU6c0KAnxb6bWiJ421kknE6q8cX2m2v6OBRYdEZBQTgX1JGMdi0
n7hww/QDG++TLFtbjPNg41Z3iwQGyr125WlSMvr7GzuKnmpuH3MtZh/6eV9lbxwd
FS/STHUhVOZmM15cEP6h6WWp6y1LrkoB73N+Jw2ZIZWn2Lqxi6SB0kj1gyLZ0QvL
p+J3tVNOgjQPMfod2XhILTyYrjxe/htM+C8tDNj8bkS5qmSWwgY+4uzawBzGXzrO
daR736unv6z6YdsfX/7OwE0Vrgbf3D7hPHQEN5FQemJOj4c7C/4hfCUgcpSvWiut
9EwbFcmTTP2mkHuNvZqs/7ty1UQVNIe154blytrpoziJceO4+NOUwVMvdDaVXZpT
IMl1+d7M99+x2uS9OGh9Z+DEkQn5faDY8l4FlXr1fH1RF8iuPfLj/X71taZcor7c
MYbel+yq0kekvX6FXfzCNb9QCZFHVhXMKqj0IJltRSoYVf7iq2+nAbxetCf81hvh
hOOkDZgxi47rxNSlR14eJ0ZbF113pkNHIlo4bfqCG0kHu1qZ0YEbH/erXvnpXViu
X+fz9FPQlzMS6y5YDEfvOTKWk9JAdmcWtXgvCRegSJOdmYjbvysaOTKX/4jhH/7w
U+S/PnV/P31m+bbPS6WJSUoblX9KgBxSPWPzEuaMlXXzH1BmKDx7hTjLjFEHdlPd
WhjCVxHIQRW41/nz+l+vLkSGUirthr/KMy1GgUC5MRATn8xsseYejI5tKKdZWlA8
w5bzvs9Tss9JjLdaWHPJ/AfxIx5IR60LAvN501B8FzHxZxmfiqwWiquw6Xx6ajV9
1g9llIdeL6FzOn2fGt7z3YD/ILSMWrfzkhTN7sxv+WAmS5DxeTHmrLwlowfVx7S8
Orw7rdQCyPYb4OdAh+TG0UUZ02rNmL6fg70BDpBqMPVHmmXqtTpxhqwNvjamT8i6
AmoFTl26IdgKYJWWXb6sz/bG5wBdB2caz8t4NHfShLJ8N6hof+Cjm4L+lOrQCoJP
NsDtJIXZiBE8CYf2fTNWOYe/3afu60FdwzTWDPXsMqSqCt3omsYGEtw2Sipkwzd9
Yu6J4OXB7BqY5qB9Rpb5Zy9/SPK6pW8NPj+gkkb0Bls9cpkWBuzq9TFyxsl1rMDl
TeyXNejrxGhDsMVx+57suVa3eLxtz3LaAE7WnGeclMktQLpRJ2GvlInY8R9XgGfF
P/fsVflWQUslPqIjSEykREp5C9/2TTL9laTJD33TmOJiIj0GjQ/TN9LlvHJ8J8sM
DWF4RfjVBJezKLplr1SRcPJDgV4eBACwz69B+PrTX+MirZ7VBNX9tPqWbPpCavu6
78XjLOVeeGARuTzsJsMqbnU6WsuUBrBiZkktVWKSAtn1x5myNO5XoI5qDBKjbuBa
pL2d4oDJB3sd35LKuOUZuhZP8J2brLuCMN8pJtpweXSqSclu05ohZKxLNNMHVLqk
gufh/JcztzXHnP41m8TwANRhQb90sXXQiqvMvnF+tXr77YhfV9InN2CJYAiBZkh4
RBCBOIhIs09J92eETY3eBXp7FxHpzef2ddLMaxxb3cUkStb74B1Ri8tOCWz51ZGK
IELTGHykDvJAsbSNASdM6/SJA5KPW6j6PldyPSranKsnOzdFSjg/HiMsE2pFN698
GA2Sq0sKGSjt3B5NsI1XoSUhMWvUq7BHaJ+/NK/ai8aOF5z+KsMTgl7nzS0HVJAB
L1LHG0UjmVs71C7BVa3o44GThazFlw1y8gMQ+ZXFS0agZz9CeKg7zo8Isil8QBzz
NSocfZLL8tHfse7kxT80zqsEroYjMt37c0Rb/eC4TEO3aBWUTz/GBaC7wagwfFov
NEtev23Ipj1cSENi6Lr9rM98m8jmB7hn4l2yLIqtXyFp/0lCU+lkvCO3mEfKf9/X
30nv6yoW1r3LFoIzFGxyf+O3Z6Ld56wFqbdrr2lYUVVg79ObqaXlOg8NDjH1T+S2
6gKpSZsRZXyTCYJ9/4FOca4HjVcH6fNPg9AWpvSG8rjDuzt8GACG0JjQT5A9A+HI
6RkwUxxsLAuH5It8zu1ncM5MQhnA4O+ymCpdKSvTPJEbiEsWbDG1NhH+vcRJTH5f
sUn9Jy8zgzIzRfAm/sc9g6c5bQ5Z0cvRq6pA4KUYPQq41G23dsuBP6Hw4y00PLKy
CdqzOeqzWhXGo0qxJ2sTB+q6L4pcZdz8wqH4fzmwC8W3jbtBVPsK+MK73JzzN/NY
4vY5lDvDtSiybV4+n4PGAfrJ9Vf8QmdojxOjQ45jGF2QlecEQrxnbHGRotHbG1+O
4np1rgDuG+rGiYQoEfp2P50riKt0vJE4348GNx7JIfUjUY5huuAujy43kuCMy7Fl
ji1+vwNgxDc0wsBFcixgbUVtLZC6MXJ2QhPmSHeu8p65U4dfUQln0RpOaSwAQOCB
gA51KlmswW+at/1RZWUDslH/McvJO5SnT12pIrKSzNmA2lmolelA13YdCUxD6Be8
PA4AyHMvksu1WxMyBUH5S9R30n9/U5oz2X6akJPxIvhaviSY+xK6HjfDFTZvvR9+
sVS5eKEAktQwRnH1f0tOySvYXU8xRFQcuxUxA2pRQbDlft8Wl5J+8JXpqcpiH6wl
+2WpNDomyTC4Ho+SfmBgE4RHk84LC3QFZ2AXCAmo+9kkdBlzBQkfF6iZdcMN66Yo
rfkjsW+owteimz3glmWb9cPXd0603esYS5qxnzLBHdY/eMRKZBFhv5HcPWY9E7Md
6rQnMRWtn35dswRLaPumOjMf4iBjzTZv4QBskHFpcdCePNqt1wxy96/BQXegLFMB
tsxJteUZNhf40bVt3kcc2s2SjaJoU83wjJIGywr1H8UQx5IelVEbNWqH0+Rgt5Z7
npEqHxHRuIQxUDSz3Oss1IXPjapwdB7HZDrcJhkbHyb2GiRz/GyNjb8/ADWRa5YP
e0m3BtdYxxSto+jXSaiGDfA3lK7D5iDozq0DQFKRx2w3u+eDvOnOjFMEq5jKaWDm
WAMtahBxX/D8HPUxtFbm6Vcm6ZJMAKHWwN2Ree3lQY8UZ16AYrXQLM+8y1NBEbmX
pKWR+zMJ/7noDO9uiDIjyrYUmnINXPda3rG8ZJehURWjur4o+rua5+aa9Wa355Vb
vn8vUNoeWUDtV0gi1woJzJw546fmav2PbmgXDwtjqDolI4NnBTQe1cbWoR1HwLHt
aLdpFwyxJJ8AT22bD4p1gDmHXaV9Vr+1Sm8r1dIoF7W4OUm870U83J79DPnkhCaT
M3LVCAwy3GIbaDv/x54u7EhAc+p8n1jo8ea+FelCD5/hkWNop4Pm0C1K2LPc/a65
tvgJuo7gLlvSs6Doebnucctqu/pdxLBYi/H54YaYoDioi6L2om4jV6nOibYr98Ty
myuWtSGwxSLqYy0Gr6kvwFyySQoFBH96jlCgPLwrV8Rq5YUdp3/77CIGsw0D+64L
O5RJB1dQ/pcH628kyXj6vvGO/BDGy2jpFf37RB4nFJgYqt9BssVPDXvz9G0YKqDL
xkkWKm+r/pblp+4L3VU5v9tq9nltQRNXPBlshHkochso8afSPlwvKh1DqLB/efxV
PRQF1hVx9cjugpILbmq9KRbYzGbanlO8dBdAJDbTBeYve2AHZMGY85h0AsnC+MN4
s+6Vqmyyl1vLosgnD5mWNp4xkTNnaeLycgCbk0q+9MfaDgeUTGeHmduSUZoelO1X
qFHbQWpd2FJKhDXgCUMTcJqAwpIqvrkwG5wmFqWJmHwkGI2LLvRutd1TvYfJ+7C1
Gj5huGGw2c+mJmzZjlERSPenuQc6aCr/rWHI1o5vucabVCYZwtsD2uZSl8n7++Tg
8zfahd/uajCncW6avah3WNf82g5yUngOmVtHcmB/gLFQhdlCAHhwjt3wlUrbYHXR
TaR2n53L7suU57CjG6OpAUD1acvKXJVk9M1HhVft0SvrEgfVxADioDEo7JwDNr+L
F3jdMZWQyUw+CCxmB+ufZqbyc6fR+YDD+2vFckuqH+msHndFMH6aKuo/EJVq2e1J
NxTLMoW4FmH2NM9vPTGg4I04hSCodzi8CfPem0H8gTq1Fhnm2L9OWwInTxsh6pwN
H41lFr5KUgwyWGRXuv/Jd2STZTG7heqt+3TflbhITtH8bhM4d2Xji3hy4o1lJZin
z5dWnz5xg2t5HDVA49p8jfh6Fj3MbAb2fuApt7tbUuPBSHfzPYzRie+6mM09VJIq
3uFQ5ztCBpxWRduA52Sf69IcK+pSOPQdqX01mzlSvSl38GxurCgQ+UOvsUQGz3IG
P4t6LJGfDoelxSpAuEHclkkCq4NpFuvqjtwX/yEf1zmBmTlMHife9MZnDryZpLLM
IRxFBvtdEkd6OYa1zf5xaQhUm3jeFz1s31guhH1LYF11kbods+IO44lgbroaDfoh
RgzF7+wZduQ6TspqjNSeDNkREGpqRBBPuCDlff7FVvyqHw24bd8rlvS1d1Pcb4xD
XtLcgjGG1LOaLGGIQXgINSzw5tWM0aeLVpukvkRbm3Z02F/3+BmNJfuFgoagmsN2
S9tahA/DU9d3avhMl3Q82y6Fd8IOP7ADTmnLoh2/X1Hwhdv0weEOP/M2E6laG+zz
Vi0PO7ibXWDz5sF26DAIXyPqRlTwrk7N/LbzdVi/sgwSOYkeq714nVJKKpFRDM1M
aAP4Or7tUVo6ElSaB58gE+Ta2ujqhTA4IaROuo/DkDdDECLbT5Ng+7EXWmNs1RMb
xV90c7jSLH+RLZcee87lT/9prGPnFfSofzilJakb/9j7GIkzRfm2DzQOJyfRL41E
8g63QP9pUsn6KpRN3Na+TxEmn63biu8KBUZ7tlL5WMIL6mA7wIbQDNxpAts3r10X
XOazANPxKSwjRy75OZSbD10BULv1FU1r8mg67JUNcOjp9dMcyhU+adfH3NQhO79V
RnoJosybboGAoGsIz7EABFF76zR46Jq6W0L3ZQv/I7VtL4UrQdL2al8bt78H0O3Y
/anJnviswtke0DrMXtvHn/lMLNmfxbVkvFMkndcNq2johkftVtZdZ1kuKhV6UYrj
qJdoo8nDKACakQnNzjKwZ6Tltz6D+G6Tlz0QiVd5JwexFxWYroIebX8Pkued48QK
66XbOsE7tvCasZ8YLi4tdAI59ZlVUO12d3ikQRBAx61W/VDR3WvhfH4G5Bs9543w
I4EMzNIumifkRhqLrWTnWAlqtkRvNwSjYWYhT0kpXqlsTE2Qg556oY03ziRYMTM7
4JCNeTxnd+YOd66mk1RHyRb96O3l9YufBxtbTmKjShtVTqpi6iJTl7haYoaRAefC
/iQOGWkd7IHzhATrNVxyxpiBE3qDSSAffZg3S3cwlqZCgEBrAhN2Yodg3oFRTR7y
rSw4L5qto2lTsKPriRlUbYfnlb1Ew9wOIQWO2951hcjTT1Y3FTaR7oMIiuJgSc3i
MI0kGNpdD8sLniuGZ3rGMv+VjMSE6bEsMlK9fQfQXvA1IORbePnmEEXO6XFsEcr0
lqbFFAnLAtxikXqwuZ1yoNkCDFWhjbTQ0MwFtJRlW0uV6ZN1vE92gCEsFSeEXQXL
08LKWgQjUUQC1xB9DFY3JtrmDx9ePSOaygd+NlzImqy0T4kVrXVtm+fewsRpAxof
afUBQQpB9GXflvU6UGrNCsNYsK1zr+483TfBZN5j4ExNFwZhJf6UL5mh5p0JR/8Q
kKmLEFa1dSsI8I3TPvts+Ma0xS9X76MVjzHdHkYmLlDtUOVELViOB17ji+4W0R72
F1dyUXQYyuvAaoc2Xi7S2jNLdCcL3qV953C18CKZlkzSovREX4Sx2FGM3djlAEbg
gQDPVHKosQpWD7Q4zVzuYxuwK6UYQm4FV4anW/cVOin+yaxBGVdX6PqCvZ3S5BS4
S4yonv9s5n72LUru+syPjC0cbN24qe9qiMi5XEYkqCF1NR7rZN21pNQ0jeSHW8Fe
6MgWMapxmdlQ65Mis7zEvMJzMqxwbXZOdFecDa1QVDMOgmw7+lYMEL3dqK4ivl/v
I+tTnNYHaPy4McEYH0PccLLc1pSklsrzxBrsTiWdevZhdGnBSxffBB3SDN4jBjJn
/uSjj0+qzy5IWSsx2ZK5GLAhA2kffhuSNXk82+MHVanXGRatRjcXb5vnxbRs/Ue2
RnyRSQZ2Jr2y0HxyLhqQNlpT6HCySt6hdB8ziFAIbLqS2Naz8po3rOreg+AjXig8
aRP/BSk3LSImz0Pac1CNS8nrfOgd5Dn67fu7hP+m4MNakkC/qk0d7CnaZhbR4FwL
STqyKS/K0jmlgFTFR0dCIIT/POo/SqksEJBwsQfeCuiIFtNF8Lr3W+DgudU6cYLI
2isuXl0x3sOba6eQD9kBVUCtoIFmvcTfRoZr/iZ3HlRTNRuvb6CZ5C3Q1n80OCE+
JRiUQ2VAUq9ut1TZkIORh/YKlYxQqpxEGw793DZRce+/GshTa4yuD7B4zuLJFV19
okpuwqj613eMIAfCT1eBwb/M/RmyBIMSebt/gcp/VC0GENxCPJFbcY7eocWdE6xT
mjBOW2fWkXV2GKBPPUdn+GWjJZVP1flPmUQWHgpbsyy5wM2N8Vhm2flNwOrzvrc0
znuucS3QduADn2vqGZJ2C/pTolGPFZV0oiLO/8/YNFgcNmJ8sx9dO5R/Dn7OyiY1
feBeRaD0jc77h82RNCgKk6ggn1xo5dIM5Xe1VcjqJ6iwXOPeokBOYHpFSp8ppL0l
p6wlY0eMaIRYb0r1I1Ldj6EuoQa1CEu9mSRSujdXRVk6g8eXuW37dqX009O7e7n/
8wxNTvRmpD5ZAt7P0ogNUTHqck2hb30T3NIhm+uUTkhL/nEWr373P/EvrR0MyDXj
MfAdyHRCotR7r+NHY+meHDaIKTz8uEs5OkGDs59jPUGk3lvQhAbVESYZQFPKz3wA
L/83feqO+BxGD8/+RsyoZxn6DUdyAsZ/j34TUzDNwWvcM91HLE2nGkw03kIDkLQs
7aNBUTQlV9LFxjal47d1vRUzZsnf/KZCaZrz5ok3/fs6RsNfdBBulNCrzFd0ZDcY
NZIa0UwTXBq2zbDmoNzwG6C0cTxAvGGj/U4U4gfN2PKPq6MQQXh/NYsnffsgmXoJ
aJrh4Ij/+iwiQTj3lCWHmeGLrhIi55u89Vvy9bwv5KdyOP4UxKZbBWDVIk+DZBY8
F2yP1T5GB6bF/zGe3+96Rwn2dxTsP8JCxjnAmEvl84vKfDMoSqSILP9U4BqYTKa6
Af8OagYdHWftBRxLbmhrcXYl4+HczBwb6bJSGq8XLc1HUFwuX1JtYk/gq1GFqq6k
ZFH5g3gu4NuBWWRMskQJJ6/74pUFMD+0RHmXOPnGuYWTAiwgr9YJ0u6r1dS9+Zkl
gq+QeRuT5EkrL2EnmgTl9xllvBWKkgy6XsY7qzNMPBKdZvx6SrsxYoB27JxGY2Zy
a3jD9vJkZCt4MBgaowOBWOQVUnpxovtEY5hr5DGLfhpSjiQ5BSQh+RtYb3FyoN++
AgdCMezlgxrucDSCRQ6NIxr9M/i2gaTFJB560cAth/sVO6RSuk5mtkAq13Abx5Id
TS2WoQnuORwnYKfnnnpnSkPA/FxUO606dUaI+hX4L2HPKVUilJ/75Uyi4dsYfSwU
0fnJXZKFOTvwk3nWnWjf0Q+qFmkZ7/PURsyvwuBHHqWaVFCE1drxQdW0HXoNwcU1
7VmjV0l0lLolCTx0wATzbA1+JwSlrlPvLdM2o+kkD4ll92uovoumByk/a+ia+vCp
qiYjwzeV612Ub0aDdI67X0Bm3z788RTr5QxCHAEzKilZyJK8CncZJXmK19MVmoIE
FRnXMakNw6vVmeW+bZdKhytP5E0eIV6m9j8vC3K6DKR3ufJSkukBenZoi/9MiJUH
lYTUDE8aA0Sdf+ZEawcUmZkuxesJHsUoWtwFhoZT5PVoNrmYXvkIsefQGSHOILv8
lbxCMk25f6ST8Wy8Vl7s4QDfyWeKMTpfmvC57xbkDueSgKA9D7SI0YNeAEnZOnDu
ydkleFJOobi8mRQa1eCmHpeUZ8wRrnBhHXJFy8+jvKqBVz4wbgN5h/sEcLk4lWv/
TMRgZ6+LTAlBURi+Uour8f0Mw5cL+fTsUx+AEjhq1Qpdcim5gefKMHjIZaMBc/bz
nDrWOGIF0nMlrv74PehkNIwGflvrLaLvQzNvZSqgJsVA0guquFXUAXGQIlE0NaSs
A+s4yn9PMddg9GrHm99YyDRZrrsKmHq/8ZzlR9Xwo/7dcOgmuBByKEcthv+VwJAL
Uqth2Kb+Xs/DR01uVsT0wf/FY4y1uTC261QDjKqatqfYeKZGqnVic3l9G5UjDZRC
YQxsEAY7HcgKEuuUj0/szh6biQgBmZTUM0FEbg6pNmGhk/r5AEKs5TKabIIrreMS
v5P1gfd0pcvqcGpwlAvnN/K+HjPD1XfxVAaqE9Wzwy5PtkERigrM4NoXjy2iXiYB
fk4pcO8wY6G0jS7rwdHPEuxTDwnYfDbN0PSyCzkAQVIJVcwxNYZfpJSSTGXpjtDB
2y6pFsDonSx41YenTDML3UgbtIotrYrlHqog/NZDu0LSOKCC6M0s8bhilbZqMPKc
/hWapofyntmlmYJzDZkdPgPCPwmvayyW2UxV322/B6lkzwkGd0Sw9ZsqPHrhN6FS
hLlYYw7IXVsPA50QGe+ZNt11W7HRoZkl39sMfgvi/JCbHduSPJ3D3bkqTCfY8v7F
PMufPpcxdDSnkqi//7fdsIg8URslfaPtGydoKd0ytMMQIVx6rBhiv7+w9wkNTvh7
6Id7Bq+H299OIuhfx1oaxS+qqG6xOFnPpWPmqXEoOSKJ1W5tZWL74qvChxezlS7p
dJERqzKOYZh19Qp1MOgugw24gbfPwEu9vz1Z2gLx6iRxsfrHKjPhH0MVjfczF1qd
XT0LCbdDNKaY8UxUE9DwPoOGDfcslqtUDHZGmoDqD1WmX6ogKICSRsJOpoyBR/Qw
J3rb+bboo4OIPPEzMgyIfMuPaFy1Y5XkG4OM6FWLC9yMbGwUHGooEBkKbiKf/RS9
0cPe4DcpLgcWuhRP6UybLwuK73zMeriFXdFYfl8g0EPjvgDA/H1QuqZnFyZSf6Kk
Ztxgx45jgpX7eUnF2ZlIYPWYgeVDGgtr0gPyohz/b2WLGm7Yt+SKzDCR8UkI9uY+
KYDQCbzaTnlD5Sayaygrqk9S5wVazoj/gzEcAW3O7ZUaPQ9Fk9rkCZ7oJ8DPawlB
tQRjTFCiMf54a5Fcjui85YuuiHpoYfM4U01+Tr/9qqtGd83k8R/+izWhiSU52xjX
+0w5q0cs69A1AQOBzugHXx6Rhe5EPGjYLhXdKJvjMWaCL88f7VhAT8qBzqRtztDY
WvLKHXI3PU6bnYTKXWZzdSIC8eqbUjpAv6hicscHr5GM9CvbYxcaKK475P9ys7Ub
KOHvwd/lE0jOV9GmpWixmtzOYV0dZGiqW/yc+3BJuYzbngL2D2ZwkCFBOAFHpdLv
4JEl4V+ASd8Bf6kp/53flzaI/zZPd0KsAc/7ngQLYZ4hPOhwMEOTelSm4Y4rJp6b
d1jFprV+0lE+EDNcTdZaFbn0Qj3418ADfMJ8Vn9cLKOi1gCtdSzVGlPXaqwJirYG
JCXF5BaEUeSAs1sYm78R4fpK8wBumxUZfCZit8qkF6h4U5hnnUVElKx/GdhZZ8R+
MpB7Yk5203I7snAuFWVcYhp+z9SLSuxBw2DpuKpgSAxf5+n25NP9wmhktkRr8Xha
MacrpHrCKHk56XsVTGtMWfT+mPgwDDwOB9g/LwotgPLLSEQALo3qr0phuk+yWzjt
wqg74TXHICUiEe9XhGQevdIf9VcDnaH3i7SyxHwVY8g0DjBMCZefoBA53GIF7w8S
AxBO2PkXegURmKSV4HEkIDsw0RExXWdwATHG7emupMsnQvEj0HBm7ne/0o4t7PX0
UB6x0KN2xqkfz9jk6mW5pvUcawqXSeP55QvnP1Y22J/Dduhs/nPhKSg/+2dAC5mK
kxevzRI2xAXpAd9yut5oYmfvcO8JK9g4W77GEKia8JtDlSOQ0r92kFCOrvhN/TZU
hA9FpIeM+iD3RIE5UbTijoFFXhejKqP29O34/b21b19CAyW4MXKO0n+j5WRvEPDu
HcTI1YlMJrc8OqRBD6n7ZSKa/IYg+FGatSlM5VmvV0TtOI4xwE6rSs4qIJgNWpiH
xa2IlcOM4sQfEHV2F1KIoaaVtO5SsVfZa5AfpV2z+GTlhoOJ4XFJVUibMCSsWUO0
WxQ6dtjooIhCA6fm0S9KVirMcJ96Ec1/bCJ5mf9pgJ7j6qsWNY6oEOfpj/rvYXxS
vRgODWXyP3di9eVd9HYoJj5aLoFmLW77RcCV/Vk+87/96l9XHcdszchAzjisleba
2JWo8nOuquIYL6Dm9FIDm0qy1bler1KOXEKRXi4AooJvHNPeNxJgwlBas5Q82bcv
bJUoTpBFpCtfiMwkBdqsFpi+Z041kqSPEsTPdid9GMVqpntOFVUGMnvWq8Z1JZ92
HZnP9O1lvz96cPfhJ/KUzKH9mejEhbDw/jOWMYcCmF5i2+xqs/jzOSdZ4UOVbBCo
xguVQa49vTjs0h8UDfBsN4FYt8DBniV6gXUDDRcbLoDeGtAiXEQdDsCp/LZpfUwN
WRRWlCF0eH7/Rc4KYs2qt9f8P9b6sHm3X1RWe46PecBv3G/MbZNW1zID3mX6R6xs
KxWaUW71bg+jxsTGXzGZ/m0K2AnaIsHkh5sLVKlkADoxnzZk5YVuIPb95rgmUK6i
slzZXlt+g7gq1ZftxgWIAQCpiB8pQNZ1qkTUmfRBBg1SfLnpZCPB0rxNxGVtNq1c
j4kfKQKNhMLGs0WhobGClg5avtUrTngoramYXL+UA1urA0rlzgMjtzjKjxI6OPYX
+kmpWoxhmbTvBkJzQvLYq3UO9se9nyL2R7HSV1BSyykbNLerH3PWnZMkuU2D94iD
nGEjwGOr/VeJuYXcxR9spFlDJe/DfUmdllyOCY1JL/8Pb4lx/VolZZjrr9I38nK3
/s86kmLgZYNqOQYEGA0i/4Z3VR3rp3AUBEBqU8z/0t0j1afAkm+bV2TjeG/GYjrG
1kGtXKm3PV/a7xEgiFkh8uSbLKunT3c/En51eqBl3ZhWuF3jPCAuLfHFtIhFnbNo
ch+1WifKIXpOh1XY7j5q8WFiiFMry8FHV6AlAwVc/eL5V0Ntho9yi+2QczzCpUI9
lEvzNKGrbKHAPGy4wVoJpUVe+JwxsU/Qppo0phh/I873deQrb+YjHw6c3zXLvEmp
vkxc1SGuBaiFR2YSN0a7Ov4I1mGueSUj4iG9RnB5W9QTsa+j/gxI3yCIe19e+vyc
VRVHx3rr+NgwT4SqJdEV8P9oo50Uz7mLRNfcu4TlFnQYt02kCMA1F9y32dUvF6wr
YUdWGAaNYCybEhyPgF5lXrx7zmtAnrMzOYPc25Y6eMGOLISImqwTXBMbyimQn3jD
GvnEARuVDafEDOy/GTL3D5/57PCC0OEJkGgFSVCFBle8JBHJvqh76kuTfDiu5QkF
vZVH2hpDEyFQV707NEVOrPdZw0DvJzsuWsHN8TG0fTcLk0Z9GwBJpj2hKQdrdxZi
Dgud8LhfM+DKAOmyy2eWXBghK0eufT8LaLGlTHbNb7Bzt+/pKmSa5jJu+IYdg9CA
uxXn7ObwjuJsWfoMjz2mNCSY0UDbGq1X/BJ/Mwfha3VtGEr//T2fCtA98WoX6kkV
tko3gEDrHKNj9gQ3MHYxcCOAUAXVIulgaYBe/1cic9cJXGxbjYLu+sJPvAIUcvvB
PgnqCARDYlKz/+5Jqw70pLqCD0hzWx/oADRF66Z4MhhtOuoTOn15Egiq2A+vkrGp
TQljb+nMkrRMwDF9iqgSC1K5yO17CbbXSdzal9SW24sSoVddBcGnWYSTJ9aq0ObQ
HBtmq16fa+6GnfR4B5ZTlo3ujuM5Rh9cMtKV2LbDiqvfq1CD/LR0GfT43aPYv5QL
LOX2AbDvbF3hgw7wptFAAqusrZjmhQauKN4ddqJsgm2wfK5qaBeOFIiEhI2D6XiM
x8qu0tUF1nVUYKrXX6KMPOOnJFlw6uc0798VYe95RHPy9R4KFGBijoSvRxYFfOwj
6IXz6Rw5JtdPTweIjJeZvMaLjDC0DxMi8GIxG/22dGpQSq1KyQCS2qHSRTN9G2ak
Jvrncn/0ABbDxN8jWXZccBnZmpkktC2Suvy45ZTwz6oQNkAlwalXwCVdeToUNC59
x/TkmJ33IqBF4/61udDY+YOSB6CUxroN8DzkizR+108n2nPAjV2d3ihRYoYBR5t1
YfCroTAXhBUd0ls+dOz7O8xVQlCkozjTo5XRhzMdzdoZMB59BrwhdduZ+BaMEKQj
dvMfyD9A8cfLyMXvNcVYjKYqgKOr+ucI4F0kyBoxPkg3K1NfXLSe1IQ1VePmrbBJ
QfMFaQPhFm6UakHbsZYGIiiWIlWsNEh7TsS/h1Gip0wdHUWnlStJ2pE19ebMVedI
Tc66luQ37RXJ5Y9MQQHAE+wZbDZG/zhziEM6clA5aSYFEDUK9EzGXie2lCMYClSw
zT6oJfzPpCxZDknuSSWPEZOJX11fhQFLmibUySWogPm4JGAIL8Bl6CVZ2jklvyQr
zNbFMe3/jZrYfKsWfWgW0SBcbKlgnSRcwaFbrAFnCXd3H9dmMcR1MiCSf3/PprAU
MHC58hn7VOV7pHqijh3TrjgMRFZ9tT1vN0hr6RbmBZZAKwY8o/bNMs8+cJagF8hb
6/MehauCLMTfcUpSsHvj1EPTKB+GYLaFWvNI8dIJFKq8+vpKchCZa4wElKsD1Jzv
4Anu0r5m12g9SjBCmtki0b+SW9hXeIJuo7gc0gqP54clmggUhrLj1gGVIgLVxzQO
lbV6Yhl+0qbqBEDKaLLKwLbDkstcmyg2LOhOwXd/ZHU5HN6mhqj5OeuVxv/BpFT+
FERTbSdmCvUlDtciXX2F1uToOW6JmLhnsslLyc77icqp9qqgvRBN3nUTcCJP28Yk
9977nRTPxdp14lefGLTT1w==
`protect END_PROTECTED
