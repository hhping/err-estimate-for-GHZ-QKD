`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYTGwUXxYyVS9j77PDeTwtg0SS+ihCEZ4N5Pghw3hHKvy0k0fnYdmwbAkhtPOJ3p
TblJ+CKoDNOWOfGdlglymKg3mIreYVvPVNR7YPk5/5BrNz/9v1UlbK3axbpBCLlW
KE2CNEkUn7j3jPaR1HqXIaemuAAG21ShhzYtwdH7mE9guGbbOdP9iZAOy3FnGBqy
pEQaOHPwd3PgIuCjlKpRVW8bkNjPAB8Jp8e+Qzpd8aVg3vTWEUFrtFzHTBDnSiQy
svNsF6R1PtvQBB5sEkK2Ven5aRb6CjVXXca9WsYpZUSYxvbBPfrVkIBvSsLFqiyK
cQnUDnGbBbYizq6GMPpAeMEJZae2vNXARHw9k4gtBAeySMX5kAb5i4zen/c2rncH
76KTuytUPPHs9QhZtOj+UR19cV/hhyTpVZeqK697luVzQXBhpbSf4N2YjbntKuG8
geVgaatEF/JlNrxhngYr2f3higaCIcTsjGhmRXmMtEzPfVHzha6BdX76vZzDsfFn
rSzWMMn72MeIKnyfxul/+VJeHPtL96ATsUvi3Y2gX2b+loIwLRu4DWw1M8z5PlJr
thCJSNtHEFT7ylegr4DzWHOlqwzy4uxHcTurnCk5PFcFDN3FlwNL0xg8YdMhWx7C
tkk2EEF9rcc9jOfOioUsPH1kZSHJOXNYLAptVEC9JLV/QbRWZ1p09WjAvPgCRmOt
vT9Jp0p/yMT5oZCpYrpwmssFA42OeLuiVoG3iJiKzTeJLo/VKi37fdVlu9pMAEZt
trPw8hz1LrRMUmnvfmmTLj7aydsucauLwjTOjtX+70751ertlFIWt/eLdKUebBMe
MSwCsuSTRphcjuYmuQHn8ix7aFMKDH9yYwuZGRZhIP6xX5776innmvxcafSAotDa
UOhpgj3DuQv7fz1Gy+dKKAWJISWIh4VtWDKAssD38IyMy3np5A19KCsSMS36+QUs
cjIa2AkMg7yrTnUeecK9g834WyMhxkuCqv1Ma+rwLPQF3I0AWXXWQTZoYQimSLor
K3c2QUPYHBnqedEiBCnuy7lC8IP3xJSXGXlQTqWGIPtBigq3pfHH0Yx1CKzrOaqH
CWebP2oH6bKnqjaRzgVVnDF3C8IM3e1VFI+Jg/6Fj9sCoFyZROHK18OrFKUUMXVA
1DT70pmCCd3dvQUk2c4o0g6C9IX8shM3Rvu7NbUCCwmZBaQycF0iz/AMArtxV7VL
QODd6P/RReOt77UV4TgtBqQLwYti8jW/z/WpKgmP/mdmbW/WBobx8pmEb0GOND/x
OMBeMdBuM/cbESkSY6iklI4sXiRToBBEnqUoe6u7ep9pgmAu/Racs8p5QXWiGP7B
FS/6PiRVc/QMhQJrPZqBiWkfGMVW76G12JyvYPuvTgNwXmIM/KqoarJtGwesIWcg
kfHbvNJCYoGoJa+xgQiPExs6a2TpDri5fIKSVXxLO8vPrmXBHGsURmJjt+1Cw+6r
V24T0KcdN+RUqT8YeW145MYiWU68l/qUlmUiirHviYRg+KgFzLFoi3KA2pscja9J
c1crfgJHGAjzaVOQo8d5biGfa49N+40F5JgakgC+Jt9H7wIr/+lrNOLxBj2HDZQ1
/R8+gdQlHR+fmniFVjmybPX8OLW+DlmiTZmTecQpFguTPFnIFMV1G2PcZPFuP03f
8PxvmyPL7movrEQPBko9lEG3e0ky7obZgCwxjSl/la7gJn3EkFbWl9TgV6u6jC+Y
odCY49v6+/jb2ruikRScd5LAHavHT/FN2yD1ZV2R4qoPDlE6Gi96UBwjDtxYJVvz
`protect END_PROTECTED
