`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HVvtAHywzLz837/bAmyG7pQ7b4KuCxf/FX6Z98h7/tL9vSqGWuEJsTVmXA88QuIr
rkeZWLoV2nMXbXWD9c9QjNp3Y35E2y6vw/syPD6BISB4wLqo24NJclQ9i/+tazYv
jGyx8P9Y4SkoSvovJKsCC4yMlelPvUbDsg+uXVWOJsMCvHz8ZracLFipSCEE/xpJ
XZq2NBsNr4yhx7UGb4LVr4YvfbOsdJKiBJ9GVsEVJ3eXS6SE5Z5K+mhrpXLiGvdD
IwDvBk30vUOrzSH0CFvVLrVLesdtsKk/mzDmkFj96oOP6xabDTOd9unSnbK543fK
7hlUS52OuUwu061+/OTe1J9Qf8+PtR6e2+i9j7AVDakC6kwVl8XH9ohEXdfwhR0b
2wopgl3x7hjaeDK3wu6ipw==
`protect END_PROTECTED
