`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rD9/8XbW2LHX9vFSYxOor64AbWr0h/USfGwjc1iJnMlqYvx05OTOoCKTly34HAbl
1f52FEya2UyJTgTJ1AzWl4B+qqYBwzxi2YQ+eQ/YYYIa0FkkEdSAHWyLdGd+ntMP
s3vH/sruI64F+ebz7m/vRo8K7B3BZYTYI2WlzQJgwhRKPO98tywYb4VrVAEXyDT8
6BIqvHbnWL1exLEQo1lFnW89NghKlnthDNDMxvDaKVpu2RsxtivQuCcM3GF89cz6
s+kWMP7SyjKW9th1GIG3QgO8qDUUaRHAnzD974FAY7RQsvL9kkqoO5wLKM4nT4uk
0oQVTv/fHujdrcv87ZOFKzxjox/W7w+lB8mhOlAsDQMUiIvKKWAr4P/0/ITXyWu4
PyTVZkntDIVoPGdrtimUDdbfuPOb6F5U4ByezifavI6HNKhPLLfFpCPiVKBuVmPO
44fViLnjmD3GJuuUOGn36Hz8gAvF/garyEnTwWZbo8QKJMBuGTfHNKm4zaHqnhMy
+ixvrg7wBz0dsVu/+CEBxGk+Xj3nHmEU6ifTDjvFtZIj7RjQipovHec8FQag0vX7
`protect END_PROTECTED
