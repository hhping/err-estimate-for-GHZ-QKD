`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a7/Kp1Z+FeZj1RPv0gxtIT9XBCuFTjVTUDDc+dPygi0w/IEeC6h7X0dOzmaDGIMY
TqEXO5W2WIdTkhgfQe4hWIc/pVDVZfGyGvFlPZeAJhQMs23udVinzZLOE0vdY9B7
68I4oESmtm+L6Klsb9q9u7JnzOR4J1Ua1KV3oO2zuShGbp3No1lMIiYVVVo3vPK3
4R0wNlypfRmpsSoKEp/uGnFVYUfgbi0/81ANyvcggp+aZkhjdzj4JXrUPi5CLcpI
xyUKBuNPkF6W68WlaXTlEK0Cm/jdsSVtVV1Fyn0PBfTqpAr0PjVI5/vDl6AXPv2j
1MahT2Eg+ovyXQlHe9UBXgK8ovUvdAmtHBOzs/WgIX2ULk/48Uas2APi8cgTTQvQ
870QdGLx+2ctobG7QO1QZyFqHS1ye3fc/nLO3OYG/13cer/qRYXa/4jFx0CRCb51
rQeBJwTRJZHTiPfJVttnuGxFGEIr6HhR8oulKT0Q07HxXzTxZOw3U5P9JlFL7szt
PkXp+i9BwnHI4H+aYjGYAgqvQiJ/26lCcyYVFUQ6yn7t2UqyU5lOvT8vurqIYvoh
ocubJA4CmKYpTnDOBwus4+OTqVwBAnSe4tXBqH/SQnUOgm4VvlMSvNN0+azo+YUO
fQ/ap2ZtUZxE//48kzXmP3+r9Q2zDUyjKvv9BjR7hx/FHRpFb0Sd+5RPngTbpXCz
XD1Wx3UxCb4nedO46v21WgHYzpg318pBKKcsBEVEwIIHSIatWylEgOyysIVQuJ9V
sE43LNZKD/cRJsUd0WgfP2xfsBEdpgYlEkplM2j+EZFITl725jUWIEjy66o5LRWU
3g6OB2ePeKqHHv9ZsPtJvxiJ30whYLX3TYr2jBmr2/zAiin7YsltLR9gWRCFQOck
Wr7QvRsRAZMP/LXHempIYYmQK3M9/P/a4VSThTelIrER/TCbzAUdd7/0+GD1Kx72
JGrCwq3yppT3LVC7Ly7Cm/a4mosZfeRZyudWp79ubDk9pv00ski2ApH74iPf/Np1
yWQDR/tuGm4UlKr0WPu5q0KpJlfd9n4Pnznp0S50Pwui55RYuiJhoilOqgdqkfG6
AlQLIeeF+sGCzjGGLWCjLTCknsGTLfHYRM/U3MQTUO4ny56SV8iYdvk56BW/aUTP
3Q+ydAjf29jHeahJRguuyY0QjYPMuHSSjShbstuZ0OlQlejOdZfYhXcqAiJKXvDo
9S1p7HIdm+iAIpEdo1bZ0IXMKo8mZ5LhIEMUwIuVVZUNfQpZuDBr/CMELEJ7KzZ8
Y4GO4kWyL6uthpx6fE/L4R3Z4Ih1wr86PZY9Pd9O4bcNSDcGxIIkXG0a/toP+OwL
ShNEft3fZJAOAnBhFPlphdH53sxfMutRA+rdafi8PuKa41xGxkNsLXl7K31UO8TO
FFbzNYwwpk10kTA4ArghE/VwgdBuVLEU2QNZarGQ3DnqNR7+Gig2DJ1zK+6AkrRA
G1xEE0sQAT6EqXYM4Yr1V1jhViWCK3bMQEYO0yB5Zs5ncM1/DGnFF1u4+57sEx2E
wLy43x5LAYZ9LQ6Jsf3mP+243mTWtv3upStTohBoMUScf9/jFcKcG9ck6jT011LC
H9hpzeptGdv161UsJQPPotJxCZLXB6JfwUDw7Owf0ajBlu8RUhEhOmPwuP8N/KvP
7x6PIQ3LcYnge2i5Cbq2mcrjkvrUeO77kUinRh9Ep0A4pmosVre8wzWXIZczHtkP
SIrwJBiQee9bdtORkPQax9VqnMqmd4J2HIUvEFhBYM3FnoYVJbLXn4NBDpPKAQI7
vnB12A/wDe3xJAEHpgGyLVsvISdcUWUcX5FkWqAjsN45tdvU8QU8h2PNM2zK7AeD
gvcTxxCRGlE2OhGswjN9NqM1WtT4AYydtVlCsvYqA4adcP0p8wgblO7tsJPtoVT0
TTeZRgmVfv/2v8qA2qSvEusDq8GbDH1NRFyiVapFKLHGT50SpLWmSA+ybVCUkSYi
ysYvZQ6j5XgG7gJte3JnMHZr1gnm+659H/vcTphEab4sAjv1GwbY5dm4kqwJd56C
gwvjZdXUDtuaLXYorudGh8xl4mhhREt55xgNMWxNx1YM0u4VLUmEPfuRYIv52fpv
wE/Di76AUWUOik4vOBPbfpPQuled8l700pJPWHrwnAKB7HIMDGwANroGEnGuQDMQ
BBVEp36lQcWrvoGD7wAD5H1Q+HqiHH0w96dEcLAF15Z/Ux4th6+o7NRgdjMDlMVh
sH7uwysrBLuRH7zlMMUNzBPcuCD0NuaTpU58l1XHoMLJk8zwQATNv6CdF+Fy4D3S
XJyPYewJLJZNR59pQDTOCOW5h2yG0Q5IotnV5ZEtESgaaE/N8vr1KTmp82fz2xda
+hHWfNrH0sGKxgWL5RsnnpATuE8EsmbsN8Cm+nOzM5l92u4NDcMQ1guQnh97noYs
WCQTCRWTe6Te8La8BD0CAzPgNvXlUbyBojXdCTzAXhEpGATaAu44ZixoakpqjnVq
s+eQmqDDL6oIeSccbfmRRWsW8QHFgiqxwozAqDu6XQR+vhLNRH+W9Ow/FfDbKHKg
cV0OUI+SERF3PsRhFSwLH8Z2EA0zetcmJwiAh37V3DVzXUfFbseTxdKQrWxvU8zV
szUuQp3aviJYK0zRemXgrZmILZyzLbTEFRyUMXXtD1Pskt4dhAtYS5zPxuS4PKPd
vSVwqBvFG6g6bmYwjASklZwZQvIVqc4XiXwbMpk6X4xafGXgSlZtZWiZgPtKo8Y4
MWAX/jUO0NjJ7R2G/YKgp33ygLsLW7U0VhHuXpDIfffFHxvtm6hAhLPiKQrdo9kJ
4Y1aU3ESylTR6iNaHo/8vhXsmnCaTLHLc54ueBVvzC98fGar/MvhDebRDXSeVkw4
lhtL1dGOFt524ICpDerO/4iPYTBh0MshodqnAnSt2zR3/lXMgJwSvhcDhCcJte5d
syvwGaKnzQlqn684w6r296GYkK2PCXnVPep9ZozcbrwheiB0R31rJ6MgvoF1j7/9
6HKaPOnSjNVEcDf1viOQzzZmZdccaAlJSwRd9d4lUvhf3PLzIz4RDUW/cR9YU/Sp
sXmqIG1EwHAeBFUO5bc/MzYTcEd0g2s2NjxOJJ/YXUHwDVstUcaXlZ8qHUcn3fGs
6R2H0WPdWwn6P8rIaT7fUWgNj9NEWOkZuSGe0pJfenF4sBJyahimAMWcGeyvjla7
vtsLU4PgfeNn5H6kBtcoWx24EMOuRBflowiBoF6LsLXTxpNdXd/q6OaNO8R8R5YU
r5tZh6s4df2DUYOZwO1YHSPzoC7c5/nzj0B/4nojvRvtfl+46qWf3L3fbW4mLOyc
EFdz0YrPBKkhrfhhnx7GCN1FIDscLPn35CEY/rNWqcd97zcpnku3qCLruee1bR+U
i2kEsDunQdexBiFkAfeNsexTGuMUJ3U16JlugY0pP2veCi1U+2NNNZz8FbLNFZ6d
7E0O5Iv8/4g7E+nPGBpNfL8XdYVVdYTZ8IbKqbPFaHP67KkjAPILIjed8lp2dIbX
enAl3I1FWpluV0sWWMfVHgfAwuYjODKn48ZBcyhAVvF8m8wxyCaHHbwsZW3xaHCB
pbYlal1cHOO9Bo8lke46UkHz8mXJj0Fuuk2ItslPm2yY+KJeb//SQSHE/BiiSCje
wqq9V8dXBHZoMy5mPI6osyeuK27u0LXYcHkoeMBTMfrbSkaSBkdNv0BxqAzOJ6Wa
sJb/cD9Ct0KSOobEAJ9/jd7eCsz1MRwtRA2Gfvapm77cYsLIrrpE2oSWfiq4IHPB
SX8NIpHjWBy3kOlH5rDgWdbdoyq3/aj9g35jUw5zu9KVq+dXWYyqTpHMyUd3uV8G
liAuvlE6+ABYPvC85WLnBuIzljC4G7yYyeQwpNPZzJ+ADCzq4I7GeEE6n7grD+AY
T1qEwkVgXM+OnBsYszQ1fuxf6mlYyUBg/tVHRZw44FjsyazOtDc7UDBfaTaE6xZ8
4qJd1cM6blffCx4QExpUHopkDnM5d4/HOfr+9YkeSoqc9zwO+cIhZWy3rznU1k8o
V58VW7e9CsNZR0rDaNfCe5JsVz4siHXmTJanyoHruanvX+joNu6YbJHqu4HPF08j
piBGWmyXo+OFq/yDCrthugDXAgOQM+Dr4R0bMGa5tEabsqhTw+A1e4ynQYLZrH1h
hXFFNC4a2/LKLsvpMD9/ic1/QfGw9x5VeJXoIKjfVxIdgHgJ/w2RNNWrWByhEid8
ts50LXpmB1fTIjd6x5jjB36za4UNHpVwwAIRg+Lwx1p0v91WVyWRt/4kEj/+MdLU
ecf0iTZk/dRN7HmyxPgO3tA4aKk1apWjrXs+AQ5Cce6guuG21bqXKdpHS1uYFXV8
7K9soKovH5Y9zI2ENrXbM0p0YGf6Mv7ZENfCA6vkbtYqxMs9xLNl9bTprtic+bCd
o9lZXXeqDiN6BIg7+RqtRTxU1l8WvSDaG1bP1Tp4Bhgk2SgQFBivjGM0MsLCOmV1
kTe8vOMTrGV2K+66chve+TeAa5R/aK0GdWBm378hARHSn2YZCB5NmlK/oLL4LcnH
UQfZNtmDOij9Y8TmZPp4Tz2VgPteio6Q0mDDFdzraqb9qfSS3LfYfH0Wo2ICBcYh
O0wettJlQVw756lEqfMiCotAl5fAY9Shy7qMHP1YTirLvV3HBN4uImAgxiC4Owa7
+98dnK6NNnrSk8nY+mQaTIwycQconnen8T7fCfDIMh000mbTZm+MZ4BqBfgC7v4N
5SPXgqJqshtN0CEVS/eqg2eNxjtdHNfPS9b/phs0XoT7OpWs27Aj2ED7xlzzac98
/b+B/o7SnLeJsrIsts6KWFxG8aEOn2VTdp1vXniTxxEJEKY5Znk1ltx04edass9O
eQlFF+JXGHnWEv0N5Rn/evROUfRqP0G9/2yWU99Meg+NnfhboB8BIVUDGX51hK74
NKKdLgdjHdi//WhNo2uFz/gfn2wfPgvMUKZTvjephNQHLUq3WPALTRNiGWc6YwCQ
+DP4GO6re7kHIcG3zHpOVugoE4QkOgfrYvmy9EpAIM9Qx4t9Z9psyXKaDlZJIO9G
68P591XDq4nle4DaBgt+wiA9LMYFSkKKNmVdRXVXkVssxnKEHj/z7vqOqZaH28qR
eypksNr41hjqNHRblMgEGTz3RrJ/1qh/giT+AhN+3kMSSVWQPa8BnPZvbPbMGkUT
fhVJfLBvBeL+LGdOvb3sXgFxezyc8y6+BM00NjjPQ+Ds8N3Bj5/063zomwMfEdyv
pUBNgZdbl3gu9h9YEdc/toBklaeE+0oAniCLNhu2LCcbjWH91HVu63Yq3+xmlL3K
axhpOUq76PhTpKSfehGhcFa9FQCO+WXuJXvkcHyMUl4H/0N3F9igBNVVRz01p3nQ
Wbam9ANXY8tpMe6/CA+nhPPC0LT3gMr5mY9RGq1/B5+j6fxL+QDQFy48CiQxpg8v
hFSX86Ubo+6xxbr+ReEeMKfKc6/shSN3o9aC5AokZJvoJl9rLjHihfb5ygZR2jWI
1I+Z5klyp19ZswwtMS5wfVMmcnDB/QyggF9UUTeTosmasAeAihrVTqoGTPC0gss4
JL21IUnk9nRB+O91ykmSKb/CvfDIam/7/mAhIl3sC6ItA2XJOGTdrY/WqG7viMCr
VSqYZ9ZJf0lxXSG7Ex0hcPuEcE7nxDNkz08En0ODOicYJD8wtQws8V7Ao3JTl8+C
nbgozOumA1OzuE6700CJLWxL+hDfGdo1s7prdvMzk3Kql+w+RJTMYBzRYNSA16Tp
UZhzLyZPpI8/t68fKxva7IPbtD85xz8dth2d96LB3+68BGFi4lGkN+1ZMUIgOAAU
uNUdkjyI6ClJOHpSS0Gwlx7HBK9ftv/4rud0rGUcgPBS8e55Vl3vHJIULmih6Tsz
bN4yuKcQhrFx8GLXIBH4E5sHiWKlu+T/MZZKtQ0AzmcE+e60ucc0HDCBwQptrSkp
OaUNmMLWrzJyXT8kvUo4iYXP+GDDK2/WaFdRvkzxEGYz7kXZL5gdjNHlbDm/Jxcq
71Orregvbr9myqX9hh1tmjC1Bn+aYrDUREe16r0aWEAWCoLOMeaZ3qaQo+7TiKeL
wwdtFTm7YTh9j2abLuOrAIps8nex9A0Ws26qPZDYIJ5vfbGCpA7Zi44CR1WOEiLB
Lznno2I75k8Hify1KiD4TsJFpg+LyWvnx6HzA0gf8dZQQY1as2ZwpEbZtEehBjgD
TUGumlBAaDqCxn4L6ezabNoBkf+0WDNL4HW1OU7T1oDbDhsFEn84z5cXNIFU51zK
rQKOZOngmU9xpSsye/yeXK0l7do9oTXD7CNa4ljmiKNGV+Jol2OOGuDnLP/PgQir
13L1jfeUY3KZpZ2PApGrftUiwhAcNMuUjwehBaXNWTAGYmgz8EMZ8q9+hZVOF7Q+
fhvNb9UCKg739ArE8sLVuj4mk10u+1AjsLsNY2R0YOe+gUFZnA4CDLsCCuORKaix
0bl7nfNC3E2P+3RNol08PdwX30CHAH+GObKtnk4VE/AINTzyEPG5my7wrUZfEncD
BbUQZgdliiydeEwbph7cR4q8ItRbhrPPcMcmjzLnckyPTC54B44f+mThrajF+7nH
fhf+O7ud7V07VDxDvARtZ0OtFGD+ApbNlxINSy4Qs7I5CP29Plr1sjd+tYqJpYAN
hsF4szf8mEh/RF1ERL6gViR7/58SDw6p+/0ubEaQ58gVcKz8v57jT77UCajXQYmp
ntpI6ouya6gjOAgzr2wB8Dfr+NDEuhWgy60ttG6fDlXh6oLngIEXKX7Cz1yBPQVa
AU9lYTUwQEoyghiKaD4xk1TzQBYdqMQz/t2tkMnVAztaYfaQAGSJt1fQQEvPo3qP
+F1Xilf4HbuDr1FHxUVrAiZ+cQxIg5gr6SZfqEI0LHW/eyVyng8Bz167J2GboIhY
sEtrxRSHHNpnSH9S/f6gOjq/BCPckf4y9tlgECXyHHfSrkNeSQ3mU9aZwkGpeD2G
NPxvrHEY411g3FZrOMFzjB7ljymO0YASwr58iNITIc5pV/nfXsnQoimpbRbcbbu6
d/mBdsJ9ZvJ7SKPsON8yIQiqF/vl2W5vuhkB42pKvzNDQiHMvTh/KK3lWd2AEAQu
EhI0NsqKUpynd0AcZFa13hzSoKVakg876fH1RcW11OVen14XSQQ5F/9Y16AM0xnJ
VBiSLKcBSji89FegQ1PWw1f6X4orUrPdK/UHgqUE21UilOIfoP7177Tr4Q4DI90V
4gkNQzNYbXPf27sMKUexWL3cDy/ul+ydjqyaTEIhFtKw/s0L4hJsVNzO1UVr9V6N
m5UMFBeuEYD2E4xmZe0dOwJ7/bIRGANNmXrVBGfyw6YDLUZf9hOu2IkpP3Mw428U
LBxWiSjUABPOUdFFcsz0dfY1xVzCimEplkpKjC3nZADRinv67gxPeNbVx8A/iXBY
hwH9VrIp335vVDGmFLE72Wp58iq2VINOPEGVDACDM7b/5epKRriiRkccFSHwTFXK
XqM6XO+SqsSUUOZ9m+o/hlEQ4b96X75dlYf2SScveq0bqnLk1YylHQ88Nq+342Qo
8gbyKpZX+lGuqXzo3ubGX4dEIwUSCBwT/dKa5KOoKdfUrdw3YBoLe1T7snOFFSsV
GPTacUDsw9zjV8ICaw1K8VtZhAXWTC3VSOBkCxGkGBt3d0MD3fK3fStw0yoNiFWp
OtE732tNJo68XdHeVknskjxhFlNFYLBDoxf4MvlvJlqawTgz7wEUHSCFoFHaBmm9
v2PjHbNOKgc6lwgEgcMKmgpVCcGKQPKdlNf09zdcw5htEYlIB4BB6DDPdTKzeb1x
XnRjgiA8E9VbRySZpJ7K3AfsMTwLKumhUtmgd6sG01B5hUmrz3Q7bNMcvHyDDmFp
q8ocYWShOtM76kJoJZv4P/Iaxq4jgVqpwL9EkiAU484c8R3oTrEi58JnMhUEK88/
xPxFdA4pTfqogdBaFK/mLKwkZI+1CWb02uI0N9uOyURn+YHthAgT25Pr+PQSKcnK
eBumoCTsqiQq7bYMZt+b6RrNYoTcxkW2+HYebEU1uCXN1GQZZVV8I4kiMwTkNJsy
HKcdVHdyV10pqvvNGDTU3fKushnnh3O7tJCevi+D+PiFiUepqj66y5JPBjigTMXj
/uAcQyxslnmfYDxlR6ee3Q4Vrg7bx5nriqhRT1G4N0XMD85J3ewGfCemzazji6Xd
XdVcaKm3Fv9y+fITqZiBlWboghiBhf/DAiNA+47Pswgp9NRzxJW3Ss74af4T6siK
V8csrwmP8zvzn8F8l6OSlSX5lq5+m+jsnM+ZMJapZ71MYjGSt6+UTqkz73vAGj+v
3Y5n+/j6Q92BnHrWlvBO3NMfS7C07RKqqbFu1wcNqIZNFgDAEWOBJ9jzlsgx1eCy
fP69wPhuQZppmnj/3Fz9cHvmzZMZ6E18U7JpXoMmfgyh4A5m13xS5oRIQZRO6fuf
+iKOuMjYtbLdqE9Hzzbt+J6TZ+q6zzPg0bnyeUG0rVKPTS9+Cxx0khCeRMp+vJW1
7xVx53Tf++gQHiKNxdOMGP4/l8K544H9i0uNFZzHs1bexhslBBVtoiqQiyz+HgWh
SuMnk8AMzy1oXoyjKY1xivBPZFWsX5MvSf8MHFo2QvMjJMZ0a0p8s4bbKXng2xfg
tQVNh2dfH+DxlzLHhP7OFLiud32MqdE0prt3ydTi5Re6cC9ULkwn0Z08RSKChCvh
JtTzXi4u9eEgA12c5df2frS/kdiVvDeyRap4cDHT1iUOHLC7bw/HHU/yi1C1eyta
tiDGD6nXtGUFlSicUmo66iLyHK7ywg4kjUCZR3gOzeYKEE9TKTVMMAQCs94gdzfU
mAgYI50Fb7LnBoGrg22TtvtyPg1jEmT+lk+gnLfyIHCGxQjPvZcYRSIKdfq0dkJO
xrM2p5zWL6d6C427nqNGcDof7h4T1aWu3ncN3/OOFEEj9pCtu2umoEy5QrNsiW7R
70/D+UI0UknshJJUAmq9r4wCzPo2/e3ZBqUzY3R9RnGcP+ZBn9Cv70NEnY8QLWBn
RU1s8ntJdL2g63EASozfuJMZb0dSgk1vLK08R7tfWFJtXYaSF9FJ4jNREFK4ENm5
GpL2v/1JC5QVGshOmL2sCYgo3bRZEKgVDOI9WT17kp11ZhXCKisQOPVQ7ifAfGy+
5v3jezcaGnOAFLW/uQMgWTDf84nmU7kHp0+AKskazQH9FQNsEU/ctBNBEu7IYySH
GnIYWxS1b8PQ4ODgLwe2YCPag041PWB3esUx/RQ2ALXSSIFzYkS6U6A5tNEwHNU3
2JBWkaayL1okHbwGLysBirdTyeAiFOeQwlxpzy3xfrfk3j5Qp2rh+Tn5r+QxIwCZ
NIuggy2iyNsRR0459hB6HCr2Eq+wI09fZxn65b0g1mEOAHAzqRFlIkZ9fWEVRFI/
Esuq7V652Miro7j93lw7oJVfXMjc+Cfc/30iRxyObK0Wy8GJ1OeeO8TA8GsTbTxo
MlSd66/Tr/MkWoSZQQEZiuMgpCzSSNLueS+fkI45xNvqs1D9SyBX4AsrosrWncDK
1Fh9T2ejTmPcZTgvtHvmxR+b2zDURvukrklbljTKLPrlfoL0ixWMwiMVgJ2YrEXA
oau2kyjIl1a5WJk5KkpMC1CcS1N09W2/SI+XyHAU9L3HEcoHZUBtmE+AZ+E1BlIv
M1Ng6GRTMmDClESFGEFHnMxJLjYZEO84psbCaqQ8zr5vCaB2FESteJt3oK7aWtRh
9PXsYVLqPg049MO/seJ1+AwxZwmerB4+Fr4UOFmTiK2jg+KJWoCEs3dInZuAZ24e
yDTmeLDnp9HTIs66OQm9gmAJmO8rMYxrXzX4le0IkeIn8RaT/MiNNEQ8tZBhXrPv
2vPIFyqSxo7AdELoT1CTHZ1WiGFWH6WyOBpkUUjf5yklw6/tfr7gOWWx+B4L0OFx
NtrQviCjlYaL0R87JLuyR16PP27pCBYxbtoZmIL1nKkaQB2m7EGd59UMTqEqsOZH
WXR9wpTEdqWib3nrH7f3PYjp5R+z3/PEcOc/+vZDQaqhWTrupCMSkCJtvYXocKVN
pNnVL7LK7MRyQ8Dm9PqWZPK0Rlepuaq3AdXRjW1yn/b3t/zP1nQv4Q804We7n0GI
cV1xOP3gA1vIismQ+Mh+B6ZuUoOxnFCU0RcV+EutY6R9urtbqFGcyXttirXREwa9
cmyazyHx1Ik0X+llDChnVRCeEMXGSb6raj8LogBS1nHW1DNiuwYqOmciu1e3LszN
Hg+5zisBIBMh3HEK/Ur6lyNTEUjTbW0C1BCNZMe/TWEjxjInSEqFwBr8Ho1u2WiV
8KluhXbPoZ1KT5fIKjfETKGuueZeAOwUf1A+nYD1RPV90amdbOOnx5K2NKGucPqj
pNiGX1dSASEY7fstrLfNrZqkiuhoYngyDKSFO/D3mSeNTJUGsZCqE2SwBLBHnLvr
/tTWVj3ajARBJXupTRjNyQqolTQLLl9dTSzDhSpNzvpr1zxLXAQv11a8R32ZGNqb
eB/9QPRIRXkeU5aKXIPxjz0M7wIV+O4r7VNfzi7p4EzX+b/+GPOEW51F5tgJpobo
fCcpKpT1umN7aIvzx1q73fNXi3Wet6du1dz6hY9/WlrwT1BZ27wjxx/rB/H8huOk
lcHlGsBfNF/NCqybpJKXcuMKtEWGcrUSs6Wf2l3UjDbLjoqVya06urVLg9ZpRMdm
njEYVjJOvNU5gLBnNL/m6krTYX8szx1RD/PY7MqG7YZSXxzWyZJ4IvrVi2uuhlJt
rvIYS3k6ybdVEmsxLTHrQZlYTXoEXJ6k+T4oaAHdG7hsG5RyG7UAkH/+YgEhhUNs
ICrijE3HlRd97swLpZPLdz4aHOh353aMwnX00u0/wHmFu1hig7JVEPCk8UkdYV3u
0uaaVqKtEMFk0NsHKacUtT1y5ZYnEhPA463LUwvdb5P9ksuhxec8J9BLzo62YQaK
86AavRHvpG+sIEWAwbUIc7KaJPcWS+DgHwVCpPf9C+djrae3oCjq+40XjkpsyEJS
Vi3RL+JwiRx9yrA0+WFiogz7CM/dBkA8u4jBO2AyL2dS0yHUBwXLuc9f/QeX6zEL
leuaCIwuvRyqJ1F9N64Khhnvu1vIMGVmW3vxAyjCSnKA4uuKhs7CRMBT9CqS04/c
MWWAabGbEOVbMjY3j7Z9aC8Zixsu3BYPTBOFpIrQS9pUbsPipNhZcLZ3Gtej2Bd1
WH0s4Tr34uaio7LdcoU4eosEhN5iIC/BLOelVM4sS4xfv1rJ+1HDdLEzETfCo5NZ
eRy46+FQy248/TduOqhEFzh+Jy+BihXxrOdmF1eIQQOpX7pImQjnXvTwnk44iTO9
ml/KDpAu5xS6LAD/TCe+PvqThArKo3aQvsd4Yb0yqEDi2l3b73UfeVeQZfTVGhL/
GvWpIdCvRQRLYtCy3yhEnt+huhvuduGKiERiG5Nq6pslEaZ1hDgq0LLwR+key1cO
Y3rYAKHBdx5MAw8F9SWY3agzIJRlLcZ+mGE7gI/cXXa1pU/uc9LdfWSBab3ztJoy
ow69+VZIRHQIJjNleGmJ07IV++Art7ZfpkbFlFgkHTVWUwREMZbHxuQMWuIZ0PGs
MZTRMOMUOMciwPdf61SRQYZ6kYJ8pAbSonZ35cqIxlA3HpLG66hJ1122qEcmAR87
IFmSCxiNy+vjS8VAUp2T7jVs1TQSnGsufoxF2wbdjXIQ5B1uK1vmyVZqJpbIm/3j
OYQDdia+Q+/9ZR+3opms+e1wvHADLntW/D9EAhgIe/ZbSMmgE+uhmMUSQlxq1/Pl
FLHOIBCbXwqXEuxIL0y80OTNJcTYK6TUoQpZdLDVi1RDxxILXT50QooEINqWIK4S
5v5MHqJ/bFPn8tr1BF6JgB3uijfx3a6QRSs0IqJ60bK0xM0WfQCpnf7iOyxyeDBO
VBjls4lHaZYpG3jYQDPWmANs1ywveT3rsXJBV6tUtGQ+I/TvpJ/uz9Pdf72alNv4
IA89TVA5ENhH0/vU8+vOLQjdUMRT52Tkvslk/QMZaUZBRYWg0lbIld7cA8/ShXfx
6gdPSROBqV2WQZuc11ULlFx3yz1BEZA+jmI/Mc5eFZ9LiQhphx55X5kUj/bNb4Ux
nrUS2b7aHrPM4EKNDhI49tjbegETwIQ9FNYkwrAAj6s41OQQ+gvHwdU/Yxj3KTfn
amuhO/tYAlg6U7wRLo3H4yAArSduVkrLqtvCTpm6GJGwzKjiOqGHWB9RxIUNLgU7
3JYM4rnrkfKX5XInCb6gMoosyVKYtzKq66kTn495JFnEptsfl3eqSrsMdEWJvblO
G+m7Ka5FwW+dM5ZwNls/SiP1Qn6ttTLm1jCEYXNZNUDqFfxqra0LyKzJX/VY629f
j7L1y6GaKsqI/A/F/jFlfisa2dW7aJMKKdLxh0lpRTdy6MsElPTU0LGJPwIR02aT
pF8b08DkaWAj09o94JBXNU5eYgs0kjkMHXtBtDhyRoTbjjrHX7518hEek01+IGE+
nvochaHWfp+NUJKmhJeHXBUNOPjFoc7jZJT0PgLSn2BVCcjSzyDRsbYGWTHwrQsc
sZhsT/8CF5fB+Gpxm6MLBZpDYPm6gqai7G/w9NqRdgm6FvVBT5uRlDKoN6rfCVey
vW366Zz6+I//ebh1iS3eJyd9Wa4zA7ohngKH5BqfSPdT36Uhwu3mhcqpSu4M5fEI
D92mFTAhFBAgFvs0suXy2SIuWRUZvunrKu2+U9yHqRqYMfa6Ltr/I84hZA1ARfVC
5XBv0klC7WQebQHxoSRpRanwW/Gx0ReaVVxxkMhkdrfJ2OKPHXaVYAF6FsNWC7FS
BV0sGA+pL0x8cKhNt1+yAoJdopXx8fbD94ovaQ4q0Jo92WTlkhmxdgCT1UrHzluL
PBqFcUlDOZEGSGtnvt2TBqkJh3h0U5vXdtPUHJgeEG0bOTN9OzC/IGgnrOUovXqn
3AnbGz+/KLGT6FQ31mNXry6DW6VCSB0Zn8tlpwiHQBHd1Us6d2Ukm/0bomwzZwkr
ITT9xlH1Qn0XUO3T1E4GJ4ye2XgjMedxxv9iQlG5bHBsh19ZR6NkRl93cO25eIyC
7KmbbKUBwGkIAm6NDbErhJXpdQ3lMIM2xzNQ6iS2bYU40cGSFqp8KaTZeVCfYr5I
S1V+loZstUADdnHa7DzWqMyXgcykcRiB9xw7VDB+tdwM9tDu6Y/CExCAKP7b9Wcz
mdeo+UtWhxYxs5PYeB5Uac1zB0OAeXIqRS98Vo4DCF2EUJCbp0x7r4sfbbZj/fMV
xYBlCJTDUH9mP5TFFHzDFaXj48YURL0ItYMgEwq93DFZPDmfy4rcQZNaK392SzcU
hKMFgCRdUepgQET2FCiWI8VtWKypQf1sqfAMTprsvrvJu2m3KwuWBECyrQodoZDw
Irq1ktOib+gHd6F0ncHOSU0bv8ZWMVsDfX0+FpLVCJxozDI523AYslKjvPKKNwJv
oc6c2fhHYIhdrxwruw/xuE3wSvy25/BVwiPvKX5O5D+DQzr98Cf3IrYiWyXSoMCh
OFfQH22wVpHGW15aSkiost23v+LwUGKmuYdj5MpEvTYVawDwSaIiyGHNAs3f0So4
f6s0IszxMitx39Ms5Q19p542C3dU5yxlreDDkE5E9ZKoOa0gAr1oDpF8/dsqNMF9
XtakUKLaz712chUF/uCHo3AFEIb8rXydJnZFXu0p/kUQJfAU74F1KWFSus2tprQg
3bJMlI7HtAULPyLfCGMrT9QUCX/rl4mhgncUyEbDqFoirzP8M6OF0ZZynqdJqrFC
9WU/1s9ym9nO7yw53uXIfUb9f217fUYIG9xoJUycrslVUawlc+Sxlhyux7iyisaV
L21Y4FOrLZAa+r4Cpii8DDsFqhauI06md/j54PcNWgHmbZ3/XqQhwEtaVmGBhRB2
wWjjEe97g6G7J00DIINNe1O+mJ9WhbHuoNDVgAMcsmPFGKBUGGtcHFigW49MKhIl
d7sd2AG0mkVQPFG7RmUkY+hDQ6yO+ShdEA0yuMeakssRfP9H0NhFmqXYPP0eMVWZ
nKoFTkOHUwuyHVgZFMVexYvNBCVXOFZG+gVUSWNQPu72IDrvwJ2z/Vs3L2+bf8Em
c3WQp9zOoelZNOu3OUFZ7Bh0fNhrBoP6MTOTTT4puPVKZemsMNMjPeCyXh6sqBrc
QPYQODU5F5MfmMi7MZdGH/UQBRqYElmn/pwFSqinj8wAT0JIDSC/9h1F4pmUWs0e
JGtN6BPI++gIe/ZH8sjkVj0bkrEb/vHnhAGe5jmJhCuk8vpntFq1MB8n7Fj+64dh
a4Jxq5BOB0GmqWvW2KvIRGAwrPsEd49263ZnOxEYwUnwO0kXN05/gcenmftk2MMd
9OTMlSW2lkn5iEtLFYDJ1TvAlXk2a5NAAtRwwSmluJa8bJusnRstI2hBA7IXUzU2
EIi1/cKPSJ0TDZp8RomltMuF/ejCeS/v2CEXBbj0g9zfDTI27Icy+ZpX0QpwryYV
7HCD6jVf51A1Bv7ziXt6aStIMUblMKyYKxZKA11JrqrPj/2WRd2yqzHhKz4z0Tll
CUvFrNw5xT1YZNA83FeVJne2xT9bwNnvP3HrUX3tHoIQ8gXTEQTL+hZe36DRrFvj
wIpUUwU6e5z7NH8NZetB0xmaEk/JUurCDx+d6JGGmkeQ2hQE4jvyN2AEP9g3Y7ff
iwr8k1Cj9mUEw8j1H4jJZkM65HblaSjXxMnSKyBCWxKNRFrIMA2E1yX1CIyXt7Jc
MkH2lIYMJKTlim7etNfMD6ewccpp3BOxw3pt9BNtA5rY/iJa37cL+lsLmtF4pOUd
LyfKmGFh3iuHEACUL101jnAV0fcGxsH5WPgYRO8fw3Elbkr79IzmCm7JOhyib/je
DPb1cJOVK4OuGFZkIXoDtRLKemkE2sJeu4YdUbipDXtEPiL7eHggmjcn8knsPgWg
2DecMdmfToLNnysBgdOFdsD9mN55+UACvCYCuOdp0J6txVHandrmSEn+N2P+ti+N
XRZdwN3kOQsOn9Qh92sj7vxHlW0WOM6MDBkHZQ1YCx+mcdGX3F012zZgfA1bMCko
8XXWnrmHYirnkG6dCLgrX++5To84N+GuGpnwiZKDhxbQdKp/hPHcfmn6wTRfaAL6
MbVR94UP15J44k/NPLA8Qsnh9A2R0jdiwM9hdUe8+F7fAeyW1n59lEepJ0qGax7D
0R3UaqrfJupaodUZSYMTJsvxLKwO/XKohxEQwROA9OPPvRp8cL5hmTdxy5lOO/ZJ
sqWdbn/RDuaIcI5ahBJwQP6j2Xbif552X9fpyOF35WmefLVUFapTJJtVnN+nGvnv
rM+cTXWafWdCqpKiibc5VcOBSjvcEUmeaJN4mjpzKWYvrXGcUgmc0TEnb6Kl1iD8
z+kqJcZiAw15V9T30iEyE8C3/uU1cUPyaqe1CYeFXzxkw1UHgrgXPkYyLHo/MIkN
g3RaZTXu2kjLPyuiYGAAw1q0RgBrLSUG3vYHIhE8XfZs2zqC6GoMxntYKiNzFVBW
gum9q1eprx35noSke0fIWEw296F0PMNE+xJ4gIpCElbKmT/vQ8uv8ZPjx8jmpQxu
CiOl/hJPKx6E+gyELWIHSe/Zv6S4yCgR6ic3gM9YXE0fhCmVvGjPluSAy+adfvUO
LOLaT9KystJqZhGOvlTLN1qvYZo1VBO9156CiaNtwVaNo1XfKSQVEWYE5xfXHLNQ
DmQT5AGslPBsUZNESCoG8HopTmzrdokFRJeYm6HVZyhzagG3OlpwwypbFhBd0DWK
JQQuDMClPka1AYOhRyek7EZNAoKb27FmmL6LMdm8UJgUQj3kqeL2a06cmqz7kUWc
D1wKiGPY7dCJO1a9L2lDmlrAklcC/Dw3CrxCJlmTSpEcoxe9WFU/bnM9bwJFT/gL
p5dt7arj21iURYYdMV+A4PJIUD6LiQxgGPtLvjGkwzS4tuYNcUQ9ovP6Rqj0ffon
2qNUdhy8JI8AdnNeldol7exOoW0XOFjP1P9ujKyl2s83YEcirDcDcSHTEP3kPHv6
5mD2UCzvY1a72i4V7ayHVDotRMxy3E0bMGVASfJY5f+nXiS87M2xhE8gcwQnFZbz
uhg/gc+OfzXORaAx7FUctMOyJqstAXl7cu8Wkt2J47e2+dR6raFIbD1yIsP4zmYE
1Nink8qiVemjlpUhEHuBT3DVOvrGXC+izz/08wKzP9BRFKOr990xmWm0DFm8/rZh
DJodUygPLVopHG+CQ0Xb7GpVJx7TUnKb3SstnQguVvMs+MEvz07TRK1y4epbmMAw
ISaz2v+bR/J/B9pGshfdHKSeRtHXAuxMFLPmt6ZyUxdVjWETvE+b6+X1QRuKeqh7
sdCzsPbqUGaCIsK+S7z6vI5Urgwua5S06wuiJySopoMAvqQ0TvAtUePIQG78id5Z
Mj6mRfoJP4T+trE1MX3Aq2Lns6Vvrsmpj39whRygl7kcJR2UhnaAhN/MurZL6vG2
oM6xIDMxgkormDQnKieaDso86wFu59gFUlQyhwNokZjYmOE5b3XrgLw7jscpT/bd
XKDkBRbgM54m0G/n8xA/AouszFrM0N4v7zB3QkklSdkKOAfJ6KiNsO1kq6vhZwmx
sS7p60rlayKUOke1Uwq6QNFWeyBGEvmkRnKySJVEB09pQrPiz8IQGl6ilPf2rb/d
/r9JKSlmfHQSiJnDGFl/9VtGCF1LLgRNuYsj9l3hf1MYhiZbbhXTuzkj+V4wwRW5
FYKPBys9WX7sqQBGaVdjWg+SZV9T0tBPJ/pKMHIOP6GwP09FBQUvHqJF3KaLNJ7s
GMB0NigvNI7Sq5Knen3+Q+BMSDt0HMz02fRGjFCHEPrb8yltweAaE5KfpG1R9EX6
0HIFG3a62HqEWVug6qlZF7lR2bF3tFyDBMV+j//L6vDduyDE2gJYvupEyox3Lq/2
LR71KJgtLpRrfaBV+soyKItfHX9+HmGLAzt3nZMF/7JAqbdov6xWWDH+KE9fYCt9
v03UbefSo7yrLObuu15jAMixBSmB/5RmimB43MoENWrKQlN2GZo+AfSWOkTBSYL4
8HN/qqa6JnVwRF7c7GJ6SljSKZeLnmYJOeyqYupwgpbcgz3hXW5JSSY6HOPHMvFM
ObkjEFEYDciVZ1qMQmD3yFQc/oaQ7T+IlaJUfhJFUp13eUTTi2Ejwd1S88p0bJE6
zJTmEP9S1QZLFbn1CLPNd8uSjMpjUoJ5uCNmKBmUzKKr4ZoLMyNPRMarPhvPgy/X
fNDXFqHerH9svjVER2ZxoiN+U1NUJpyvinAHZ1xtNvbwYfQo3CvgEiElYsjLOzZJ
VxgUlavtJr8eOw9i3TEujEofoZRd2hfdAxyOj8WX7+g6ZlkAtrAyjgrNCb0vIgv0
tTCdphhwyOBXnIuByTDRJnGY4GBQrxzDUEcu1TyvDF5pDPi4vDvrBjNW/iiCD4ZK
hjVbT6Db4gK8j49sn5eZZqg2RA5opxxtJexUt3PrRnATmNyq5FQgKa402TFrs/o2
yH8M9NAlrgoqT/66yfontqYlpuqlVz/s5KxXgUMgaJfXwbxoYIMMCJzqyd+gN5ev
0uOLsZCiXnVftpsCTeAuL1xwFLi+gbGBxOMybkOHLo8gk1wFNfSQl7b2X6WKCfSs
iQ5FUMgC7xexMPnRlA0oZsI55r8FsB4SIe56RT8ZQC3UjAqd/znwLUhhyViEY0MJ
b+uAST9aSf31AyAWD20/El5rmmFdNKyn5IR4iys+osZ84kaQsiFV8tCYh/vSqhTq
sTN6haXS0+EO1IKJZfkm6XmklbMHOC1R1VyzrhkipsPRkL6fhYDoveTa0t8nDPpa
aBy2eZ9ygKJnkmh4nshUd6X5DZLvnlujVAuKtxuFi0mLT2rIZU6F65XYeCNggul8
6Fu2hMM5R8Fd3Zt3YaCIiU+tUuWhWPAF5HmpMOa6mMcb3BjHjBRQac/8tEFKkK5R
NI3SvX8CBWOrw6QAxHsspZX53AQ6TpQ63JrUtBzNRemH7OuBaoUpsE8Mjvf41rZf
03XlnQxPUjUWHcQ803QSzg3eDLHWureP1lE3aEMpj9O31JZQpFuzBs6AVwVTTZzO
+15ASv3mZq29mRVykYDB8qRCIzce22+Bw4nD0Cg9b7sNpUkSWvLFFcQOgbZI4zjv
HVKAsWXufLjlMc/DPr5xmjcpf5YTqzLt2cCMUsukUxjxqBWGxnEm/7VA9XWPfWgI
PqsSafa25QWYVMQP9U0oHHxLr2dEdV4vtBQVhvoeMKjwkXPHVtcCjYsSG9LIHurB
LL2FkdWzNdHCknUPX1a4xloiXeJau8Vow8wIC70YvEMPqLBJAjYMrEEV/BbLu3ss
6hzjHd+r5TRgdDtj5aCsa5OqOENBFZ/tRu82hKQk8GAhe3xNZZP1XxJeixFddESA
b6Iq9KzPyaqMis6TzIa+VTCBUppYigyn9Ynm9EubAUAfrrq9OjTYdrw8pu2XFwvB
TnV6A7SN6IKorfx2TAnY0cNCxEet0owQdksohu6KG8Dea2pLwvZaTqs+jTDAqUDw
houhrAHdryawZ+EqLkQ7kNsZvh26KPE72YUVKwBz7Sz2UyK2ExJZ86eQhPhjztSV
dNvP0rBRJrxz1G2Ca/uowaoGdd8Wu8J8PTCi/V+K5E7wAAN+W7K9Mee9vBqzyiLj
dZSfQtq6RDTXBw50hnI+1GSXsUTbsM6I5EjOlbedCnlCyxZ7DHUVty2Oism6yj9l
a8VjqPZredx7tILBrLjL8hKGYIcAipNNVzcooXM/7Yk7Hm3Y9ZT87I2THfg3bSIH
FcFGmPiF7pWJPwtc7TjS9vzRnGZzMrogmamOMVv4SYsYS7V28CEhAAYnhPGwU4p+
vL6TdYIgfNoZnhfKkgEoAw9JnV52GwhR0EQAJAr8ktkkNyIRIk+Iq4ZqQMKIRUAl
H5Ad3se4YG4x4BNFltCGR6TnF9Uy/1uEq5ZR4hO1Dn2K9lpjBzjhun1VuleTpZN9
KffCIW1UtCAsbh//2PI/oawn7gkVd9/VS7hJ1iBV+MU8WDBPXNp51vM26b8JAE+G
xC7l7+saWOWzZLJzY/5xtSE+z2VqHWOGAtjz1GAS72yj5hHjuzGw0vmuAopL36Zm
gaOmCz7xwlQZLNCtB0Xg3JV3LLzhFfa1QAIIg2GJdjR34eFtRT2EP3sckExXhqS9
8Ii5GqLo+lYcwT2tYXK9bEBnunGnjBq91ZrhsAHzKNq9gtNZWA0d/84a7my0BhQL
7qxHRu0Z+xdZVG3eo6caB27MttzO3Dp0vCH+uD0v6DrpMqhs2DfCgKjNqG+PuQVJ
1K+B9M27b3Jc/bDv3wsbt1h0YGyQMyhyOpNiXpdk6Y3uhwgZgy7Fe62dWdySndjg
TVhBw83R0CaQ/Ac2udZYd7eJQwlxAvYrj5hoGOMd4GnADg8aOdKVx3Fn3DBwxqJs
3KqmZRJQx6AAvydLoIz/n+bHVsYM+9rYup9WNcuQzPR6RGYlScldGNdgg61rwI/P
Z58k+NzRTGKPfX4iRsicxKLY2S9xxhdIJECFmZf7sCRB3tznHnRCz0vbiHtbfeRf
2NS31EFeW1EBY8CCsjpR5g+gvMsR5FQHHwwC/jv8y+Vta5OXFUzkEyoxj8YWN4tD
g90oqqIeixYfH/ctwtA9l1I3jpNVAfvnlZJ1t/y3ySK/E+r/5UX+GsmR9I7WYEfC
mewyI2hRD5l6IXeWTqtGMx/EygX9Q4LDhUv99RL0ZdW9blrVKKuS4wNKEbfpJyvH
EqZIaCniNyzNu75Co8HkKwgV96AeXcfcxSjpJiw9rqXnmJfTofOu2b93hyrrmL38
B1D/JOokplDeKtJw5NopTxA8c4+kjnhMK5Wnl4yNE8H5s00GaQB+heO5Th1e+VHM
Ov1GQL/eALyyqbuR710QP5NFyhezGjPe4Kd7redvmmDnQct0cbW6yLHucQuz6N20
5Kg+k9nGugzV3S/orEx+/VowJoawpNmNGnpimoZZ+xvl5kii1Fhr625yIst1ltxx
EIaiVaShyep0PfbZPwzRrJF5185Dn6ILB5Llocb0INhGCQaCRJNEjQixkWshjw44
rOnQruHmUSGUm/zBY202f/qxPcuOqDlePyburNy898SjV+J2VhY5nhlfLzrsURWi
oV7IgZJk5+PtJ4T6cyUg8nuTX1gfUlmrhnU2C5Gl3smsPjjFRN2fvnx/VekQSWwr
wVEVXFUFVC9J0TFRqNsn8UQ7fTBIth7kmCfb3VRWxKr2BhQa6qnwHJorB7b9me8J
ybLFNozrO5bcCVclnq9lp/KFdPGRN++v5ttkfb+54LU97zyKFnneLlygtN6BfFCP
L4om/XyH40TFnopqdUz4GQv9gOQ4fsgGiv2+8/0hqNMT9EpuTxxGkOnbNPtsXbrm
5sRky5PsJweoMwzw7goTP0lbZ+Ydi563Atm1/IPqaFOyBCP3hjXytvsweDPw4NgO
DA7w2eAEITZoKFtLZGOTQnRk6iW8rRfWrnJvaiL8v7FZxsCAX6edf4dvdsZRp60N
j+gnWMCa3kLqGQht8Key3Bq0ZQMsrNEen47PtJpx6ngdUkRPd0uaHvuyl2ez/azu
HQZ9qR8YQaWjLBn7YA2qUbszL6Kj00yKBPB6u4sZph5f8pVgAFg9IGUQ2K7A9tpz
PtLbYw/OgPwvbBvuO3AF89QHurv64nDMWblUfV/iIqRluG1X04UwMQu3jCuYfSBq
uQAb5oZPKP4QAYNKHqO4HCgDmP5+u7Rc8mWQUgnuKhMyRYD7q72RM9Tn5QXGbU8T
iEDkKJ6c+1icCZLNUSVBvRs8q2CplqqFJk1zgL65Mrwvtt7VC3/VzQMvozueVJqQ
CfCwmAM/+61ZL1qwwNHuafpKTvxXjXLfNpDtLj3pHrYKnWzkVskMCRe1UeUJOvpi
wLUT0P5TMpKRbJA0AmrlI7M1thb1pKuWU7FOLNLnvQls7gpr30JRA/lFx1etmlCb
VDqC6DsAAVplGmU78z+J7LkUF/mPG4y59/bYFusJNcRFjtkzaJB5+ZDQZUV3Stw5
/R3pUQxwFUgpmZpWZZjzCFuEIyxkeYdyXGiFEkR1Rjz+/FczQwFvJQzQIFjW7VgO
qvBiAJWcJHOP252PM0DCFilY/W+UGdtJmWetmeWf79fbGdQI/DhuqgfiUF7K2AxI
Zcdd71M3qFeiDWgZod3y8tqJJANFe0lz5SW4hwScREacmdprsmHvIL15e7Ddu5i3
AH7UOpmV1Fv0knn/YrC1IXe9GYWhqgcAciTU4MeDV+jT/KkYCwyMubEINfhNfzLF
k+y00OfVSI5xTRots4Xkv4ZgO8Ce4FwfbDUW06tioWnKjYMm3DiTls/ImDWLrAv0
ac6K3Kc+EuJxrgG/rQnCUAigW+8cdatMCkEWF+AYeX4SJsoHjpdIdYUc5WNJSMiC
Te8sPMF8S8WtK3uqDHXgjbTiLujHc85JRwOHVGL0wf0dWAv94G7bKHCaeFuOoNfC
B6ToyLBZKc1yS5mtqMQ4P41VRnloqXi4AECKagSWgB1/LuAMhk818+z7dlt/6RHZ
XoL+NAgqYscFyA94F7sp9ey0jL32WWPwpXVZJ0KUe8Sr9ebdRkIfOdEgqobOKxMT
n4dgohbb0/5ZVCvWuTcETYKxIbjtR42VqXICJhdosNzQNxC7jgNyYmfM6hWtBnwG
dkthvaN+GThC4QmGBv7T7Elqxg2hk6HuKx9+QHnK4bfUg7YCp3T4lJEW1GOtksU9
BVj7v9oZtJ1EHjUWZrWib3Z3McEZ3esUjMzBgC8wk2TaciyHeDk+G5PK80bfFvOu
isHb9pt7kphKbtFG47HJalDj3lyyxydypIQuGKOAmNT6ZsrzkK5hWa7ernPi6nI/
16vZ/69SO9Me56qIVXhOn2iPARCVa0WthwXceelUOM3KIvufJO+5eeQWMNX1hu4K
VZfQaqlG+TQxzdHxtWbw4k64L0QxgI9oj0ZS4pERSTEAlaxnv7CWHIOA+XKjeZLh
l0PHtrxJkbxBj6i9LFtXhSIZ5WX87VoQkhvWz4hENJPvRJPz8VwtmQXFvjg2PeYe
OejtjNKDwVAxhIpAJTH/bHgk0itEExGXK5ntmVeAamtHLKbuh3nVpmrripoVr62N
FnU29BnW/n+oVtezQfiT5SAiW2KK7xVXIi5K5b85/LVvzVv6renaGr11Z5C1dp6c
4ia5aSXTCE1wWYLggwhuXpMhVhGxlZm60lSxzZGZuu8INUjji9RfyBrxepTuM4Cn
GDmIlmg+ljHxRt6kuew6TAldCdM6wKoU4flcdmg0y0K1DBpo1C+wSKh0wqJTgDLk
1QQdGtRKmVwpu+sQ4syhZtNH0FhpzOkgSe/s8W0etXrtUQ6kK7CF7EYVLFREYFEt
o2nLfViX/vQG8dxB+v230VAHyIPPKINUb17+ZsufEPp+C1roBXCQbOzcPgkGL5rB
/fm0P8AIsF6nDyxz9eCLSRy/Z7YQpXwtSgESiMLW/X4s6BK3NZWsRliWcjtRV5N8
5GXpS7/Z25e7NXvGAx5Ublv+R6tCStlT9TdjiiVpUHar77O0LV/zScJAO0EJIv2V
eECENtyzlbLX7m5VzyVDmtJeYT7yNSd6dJtsYCRUtlr/Cojff6S3hvh+yHaBuF9n
s5kdaJ5+D/99A/LU5eXWgF3APX/otztZ2BQ1lnxPguTSMXBAn9m504Dxl8wP5Cy+
xALoyEafhL74wWuzFCGkGiH0d9aOtO2x1gpFsgpxVWqIY87SkKCu52NPt1x71RKh
BRsh/f48jGj6Sokx2UrcvH028k/A9Vmfi+4b2Bobaln2eJnhHNrgCc9LK8cNJwFj
ahTjFs6D+rtzuq9hz42WxTTn1GYdSajnovH/yVXZmBr/9jN1qRGg7+CU98MZajKG
eSrTOh/ryMZ83xuo6yalBwPkPJSbo7capoFdDySeHo+bD3+JqdP6e+G2j+k/eIpf
rRZ0sf8Ny5I6fD7i3HgdRu2Whtpne8vDo0RVlD53+JBf1m69wM0Sn1peicopDK3b
18pGTbvaop2vIwtZNr6K3a9Fdpf1uqpYK7o5ky9liKWRZEb5SlfHfgVPkx0sUqpb
N6a/zq3TcXpiqHv4Kr18IHRO764xUsZRC8wZIXwHxePAuJ5hzzFWXfwDEwMPWEUp
xN5wi/aU10TqJyvQydTPINV6PUqRVFyK3MM6gmFmDl19xoGxJhCNm1bRSZ9BHB7G
lnuBQcmKgk72cvKiLC6mdLu1J7ams2ySahpayRtS+NthErILBU9u136g/vxj8lMJ
TJbFKlO+/Mzp+gBEqTGk0CUhlHHhGrUeqWJ2hjHuXxKmpuPzNv5nysJd77f1ke38
jWhJHodQL71nPDKkpciKfVLviBEvZGR6cnpuQArL6yoI2C+LBRGo0e19sYdEmkAr
gPhEsJB4nzHxAquBHDahGZx11J8z5ups40HLqhaB7UXYdOxCrd5qGhWWJX6NI5U+
9utBdKMvCaGS2CaWaQMEMx4DXg2e1397TzxqbGiAbF4+YxLOfH8FXDRFGJ/DHehC
ops0vpF4Ra2K0bVMVKJk7QmFuGUC5c6yFR8ligLts8wEfIK62qIe2mO2aAvyqiYI
ZktnJUJ3mm3HOkwQePNt/V5cgPPJLHvM+CPadF6ZUtJW8dtMHy6xzCS5AY13fCf8
jBGHL6D873ZNu/3PYEoKQH/HaBZ5SO5/odVNbBJ6ohO635Ch20/Wd/JrVpKQsliw
RATWIfsE5jk8TOYJEpP467xrZBMoQjsWUsEhDMNyq8Pyy3sPNzm/q1cAnmY8/TL+
jVgU72wCe/f0yR0Xlpk4jojNYEyXg9+llEeqiULwyEMvqLQp9VB1glA6rojsjw+T
gHz1cdjIaIxGmqk0FyePhjevME6ekO1NKbDy0FEEogITxuHojkpiMTeV104GlVFi
so+LBjvsKGSG743TrlKegOiZv03rKEY/S1d0x18SxH2ChZ+bF7gLqTf7HseeH8SA
rFE4cHX+tMAyO1qTRmBu2pGT1hhRORYxqiFOpbwc7l+3Wkwx8PGiUAJhpKaQmbAQ
gpKq6TLhbQFpUKBQgVX3LVRrFrEzaK/7h9lXeiuggsobcIWoxkvUychlVbJJRmt4
g8aoWlXhPzCMfflhEZJK0ZKS9z1l5u85tZynM4TY5TF8JVJvBzre2OypJTuKq8lC
8EUumOzoUQd/HaCme7BPsutNmE/N/bZ8MPO0EGEIFYACuP2myDinyfN4B9nhSKrL
LPP7rTkQ8qwtlzievPLvgCG8TniXs+LekV4HrAVVWfFTM5IxsM/36oIJNyXCDAVl
9SHqrd/apGNpEp6l/t5P2bPxE8fl3vkO1/xyu2hfuK2m9r2Og9S/TlBh4dNMNjwk
VX8PVyU2GqSyHNGJ835F3lIMQccXLnvHeABdJQ15G20lu9FayffJ5IsdyPQGum3q
QDafJ/98pnT4njN1lHPIu9AhvzeYANnGaVrRVMYt0wO8MfJSMxLK0Z4nr65vb8aA
KjDhO+aWE4Yh2+JifGSDsupYx95Xq7COXeuXuYCHjT1+q54WdMygxA+kRbqj/8oJ
SkxbozKGAklptLhbFSwla4VtI8nshs4vYQxbdjDxSMkf6XJLp/T53M4i6XYQ54vd
oPEM1dB7nXWaZccjylg/AOZlgQt1YjxV1x/UodthlvFBhFdFNDnqIMHoa5Wt9Btk
e264TSa8vBUmu9a5kt1JKS/JaqOLJXOE+Furm2FGWEyaBF8+QZBa4iS8r5bJO+gu
outFENvvZKrmACndRXzHkLvR4Hb6JxKQP/66F1SpAOYRHWRCwjMZKySzuhz3hMdS
Iwh3O+gQ0btsobs8bN1dBOVoaHvUfw1JrokrfRWlItSgYeUU9j/4BOoKsbCx9o2a
sQ2kVlCr6po6KOZK1EFpTbeW65wSP2bPY1WlgoVuIOFX4teJ1Epit7oO+0pF7pZL
uq8L+yBqXOec5jfrwwmeTQ5PoGOa9Mv+GgWDvpvD9cICapRj1tmnD9+H3g0iLUsK
EU4wInKAC8T+Fh9RViYIHK/LT0lH2jjilsMXeToFQUlbQFmw23bV9DmWGUEO5VzT
wjvdmW8Plxo2204PaHbVujCevyoTMMCAT3ktHNQ2zNSTJJ9c2PqwXHH13PwvWQ46
v0HBzF0btnyvJH+muSs/78uUH3wo6t8nZeRllZF9ry7TXwn9Cj8YEWw8FZE+mBAf
hwoa9smiGHFFdAbHiZoDTF7+C05qZX9o1mEE+Fh+GMYNX7FtOd8l0oMxwNtG3Jed
tF+vt6teRNGwkJDGU5XyL+QuDOzSiyF0HOmn0QTdeWMNOV/Prc0fZ+3Q5ublpsIw
zm00TedDCQTIcMyvcP6UKwDvP9gy9bkHR8miONg5pKwDtL4eRWx9VkmGsz11xX/c
q7GTX5NwIuNLQQbMLa14tx2OLWFBYolpZp+pVb8mEghFgGMO39CH3cBdTtzko34I
HoSjyoq5hxs2Rz7ovROLDWxVlI+Z+iZlzkoOicJE04rKKU8usk1yc3AuEJu7P8m7
nvOjFRqHA55zMiy2V0x8Ek+uCxfqsYRos7c6lbggAiF9XM0r71ALnS6gCO2CDtzu
nRCjyE9fFt5qw6sgC2Aa5VXJkcNrdNcvSaw9XzCEtbYsNg2DTv+oItcDX5eahLEr
CyeR0KZdV087eUMXU1HFbNOlHxoWCb8XHOVsHfEu23oxa1PNMHFHza/UXTAfaRVa
hKI/tcJGbRDBRyIUU7APzeJV18R5qbwdcBDSbyK95Pf/RjLyTUErCgWtRS4D+4qK
39/cO76SllHToaYkcc8sEkn5uN2unuEUgol9BcaFVh4Jy/z+UkV6nAdKrw4gcOR2
Do1ZV+XPSzyEiHFq6B6zdlpgb+VjjfK/4fc2A7lx2jwW9bCt5y0nJfdZ/2HW2jx5
gdHMfG8wNViPUAF55RFaF8ogqzavDyN6KM0ZkLt7O0oJ3mQD3sx8EommWfQVSO5t
Vaxgc3bpqwiUVolPlQ798y+ofJM5gTL5eb+U89MhRd+OT/niWmn/Tdbvaa7T01MO
IY5iFji9HrWT2dixFqtb1FpMu1UXaIsEyCCdh/5TTAITW4JzpY9iUxhq5s6wwoCF
bkaifEVaMvjd6x6y+5OGES47cMLrOybrDmbzd+1lftVrUSz4EMhcK2eJ/lZ48Pg4
EVb6KC26kk6oMzWhJD5RbuOCZblV1h2v2qjRUlS0FSkyt2krj6WqRWgzFiAK0u+g
rYy0LV0lGLrxiA0HQNBLApnf1ShM6GBblTUrWxYrwPKjI7gh/aoG1Dg6YUOrij9g
4CH+/VfN5DhyFqZGQ9daQQvvEVYO5bc+LaB1AlbUjOf/byONYM6OucV97r4N7QYW
VY0j0naEwcJSdqLjBOlbTUoYK+MERQ27aZJyiC9yX8m7p1l3jwZbDmxnpfMvKpKv
hxV6UA8lqb2H0NCpJxEXAKBsTK9c7OCsrfsQBu0UveokRydd8pbWjrbF/Kora/qi
Al1JrKIGvjWABrjbbC29V+eUCQ0h7vGUWoplhN4j5Vo/fCk6FXZFCgqLNaRjP1y4
Rg/A7WA6pbTj9R0xFdqskWhjouqxl6mXa7lAlFU8JPXtCgVb0gKKoaWeszmO5FBQ
DCon/huQ16uiFdA4l9gciPilst2ZDz3hGq6oGIo8HltwL+N/+rYiMT+dYLyqkmJ9
nXfMsCaH1I7VOnsbOCF17gdXXPg22FVuAt1jeM/Qk8cC4IbOfYfRsz62zQTaLAkW
IXbK8EvZvPrkZCwoyuTtzUn1cnGCQJJWDiDno2PUgeDnxWKgWkNPkFVrIeY/xr+w
02UY7laeqyUHdnApId8JuvwpLwOVQ+kWvnhKyCcgNl+RytyN72mN5AHKrqfyEYiI
gbzdNKRnGjwrQCK++jv6xL1GTNNeexA/KSkPZxOPqmeDyAduWxAGc6YVSIUTo3pW
FIfXy/zmh0/vtznYWDt2mvjEQdXCJS0qb9Co8mssjUzF2ukaDcwEGaUfXc2UE4HL
sN80o6ajSg1FvwXMUPI4EYrkbFkCVDyHw4a0Yi9dBg8A8fRjMfBu87OvgAYfwFOV
NYYX2hbS/WVIQgTqyETpRUSAF1HwRnVqYc7QRvKkxM9rcWM4P5m39tL0lcLZB/Q5
j9TZJCroSBe0aMIdi7tSC2zsnNQUDw5ngz56sr2u19JcQ5Pw0J1prQ+QKeAiHHp1
XSEh+v9NiuuA1tIlP06oYR6+t24s4qXOhJ0Fk0YjFMtnLP7tf+EzAS1JlYtUK2vl
2Llcatw4kYezfMQ4nThA4L4BYgiO2qbnlk4g/IyIM8+1TUq548xeCtziMdoRsCA0
B3dHAxhd41kTQ/7kvMBubkJAylNquwc6a0ALD+R9aSxAHMFMzXDwJn40LPkMIrf3
GJwaZkhNVePRvQ4IBb+tkRGYlbvG/OMAZU6tXWPedmBfJB0Fk3CnXhiacGrF+8Bn
3PU8LmZpyLlv2Ptp1c+7LjjinDFqz/q97qga93Ax6dd4ppqjbuBB2FaXOVSC3M53
ATrDLbKQtC3j+sC0geY3YDeRHOaBQ92Sll71jX2n+DEUidGvhnaXhf5jqDL5p1wt
Y3NVLHvwMECxr/4LbSlaoYmKti566W//zVcviR5e9MJVuthel2BvSe1EGiRtt0/z
twB04HdFm6PEHYBGF6kJnMN/X4rX2o8tO9KiwQNz+0M2fHffku4SsbQznNmXJopZ
A/aJC3720erY5k2PxfUogktBao2dQuyUMUApjcHsUv2EV6uBgorMsf4b/FX8/BUu
AubTNJFH2V0tM0Vol5x3SDKy6cS2HGAFxYuFotutCBmCehyUy7cRd0RJb/VNI+/l
XQccVRZG6DG4TpZ1gqAZVnRUsNk5xDX4Gv18mgWzEFkXWSSo85+LZGKniHzM6MFC
uTdIIRdxBgkQtZhgtwOEfdjx12B7QOGFB2MFLGCLbCkt5zaJHmT6+g/mC1bBjptU
2k1bci11bfqx7QIOqVHk1Oa9/yofW4hjRznDb07N8BxxJUAVe7Y5uBCekXHYQdM8
8FJFE4C8bVvdciq2ak1xeWFbcu0jGLhT0TenabXBNPwN72a6/8xb0aJE65Yk9KgP
i/nrttEUhS0t8Sn7qY264+Gip4zAzT5R3hMvlS2Lq1IPVTSMej5VhGP6c+RwDOzw
/4L8Sx7QNxj1Ci87xM7wR4dxFMRjFSmbHaWuXe4XApilPhrejW1YuAnBkWuFBOjs
neizPHMqlqDjfls8PYL7zu0q4QMIMMP0AYv6eYeZ3kkQIGgQNfsv4hagbQneShPi
uYy/kP4DWZKvdLEJP7NqoFq8EahHYI+AURgzTV2IFfbtMLV4bxZ7bXqkfLz8lD61
JfJgxaeEZ8+8T7EdzK7QdA0LzCGWhxh94MH5N+TP/dMbzfeE6zzTU0VKaqEcma3A
3H0qLA2GvMWv3PbaOFVE8sXX41CfIsOWqcgPJvCYlgDFl2j/Vj1sRLQUnNk91Kg4
rZ+Wh8DlJS7z0U9IdgGgMCcu3v7tEI5ODiLMTpH8ZDqa1KNf5HAvkXlNCoC9yCl8
At+anksTCdGw1UT1Y0H4hu/lk+WSaixtrsFrA7QHVxgFid3Y2yNmQciefsIW3LUn
SiUwpoihnbGi1Npj1M9lMlhiCdig/pUoTGOWAjXfKM77C8jvryqzWX8P/WjBXc0U
X3QlHPCefLPUxDxYgThBVbBU/dwHr79z2BelfbxoAjUHbDMDg+ZC/y7SRK4hZ+Pv
YDZX8QK3NrWeybPtKJyHbV6CL1plHVO3q/LQuaBZDSyaKGZeWdZaPizkO1qpwoD8
1ZbaWcbUOz9KlCv/UNmMoi98ZR4iUFa5LZaejocwVtllvy5IUa22u5QwwIwiuYTp
ZOIkgSlSv2p7n2y9AvjRbCYBO88oL5R7WYbu6X3EkZVY+1o1imdMrLZajrTstNwi
zDaMs5dKf2JTbCAXVuICBbHlkj6IySZr13NJNBeEYMT5fmB4NULR/BpgETleURPC
iNn59uRcZMTDeHgmty9ReYCgpcak+NHXPtzkO2h7dYNJfuh56fvUvy9WfJbSMSpL
CFbkVvuYLGS0LJ4fnORfollzby0UeDkHc8Yk7BLD0Knvtv6L5SChYzB9H1uQzamo
9KJwU4+1tInRB31Kmvo3+7+YkxDpYpphpUzWRu4ixGDKUbvbnbHOzP0dqqG/4em1
SmeyaMD/RhbZPNk2J6Ob+N1jJwUthETwU90rvFDaFCP4kt8n72t5mXtMPTGx37+n
2a0MxqWd4zYQ+dk0bQLvwBpEA19ipl2KRrQh4EbDTdhG8vlTYuPEiyexcLochRLw
bsGH077ab8LBX4gnOCU71jx5uA9/pLykGsNwzSahjqTwgKYh+kZI49K3jetWfAuz
Vznxlw4pijTHkb2Z+113xLx1vVVMYF4TtTCoP8VZnRRM2sLEoabVZ8+xyBKh4FdL
NF0GvFWwi4OPCvZr9rVdHSNF9ULcMgbNPt6dysPSdn8iDQcpOJEgbcwli+bw/w2v
uZvky9cdM8WJTsUgeymeaKJ4UrXxtUhx7p2H8K9qLHt+4qKquc9QJ1w9cHgFNfQH
zdsdGjej342SGeuwNoVmDjD1T4+yVLm+KUL4PVT9eg0CzraIq6/+T4lBtJq04tQv
AS6jaV1PspigE/NLmDTBnSUR/y76VwQvCP3UPF1Mf74a9v5EbkiwbmTt0RbtfCSl
cYp1Qb7b6yisqVyGtqP2GyvGLZtq7M8gl2emCNN0pZsatHTQUYObAXlWDkBfH8A2
UvDHIBvMxuEMcbnjbNFKxjM7GECGgzXXQHu/IVa71rjZVtWFDhtdjnnZIXx7vWP3
R4GwkYCDz9I99fO5U7eEWXOT0EKwlHiMP2aoeYLvx9Btl/3BWT3B65gNXOoXIBQ3
PxfCg0jz7GbxDk883QHVva0rlmMYqxf8dhCqe/T0ydTYbHDmC7T1DY3iFhA83sad
yK/3OT1dMSYLa30obdFjOLJtA31+583Ou7eS0wIixe4xeurDoRsBr/YRgPKAByFT
1rnJ6OxA/OOPv3V4U6eCg0LUb7JZ7egU1fmoVKrJGv8WltSetKD8uUeWjQRBgKbY
T/+LNOaO1cIk/mWH/2834cJucmIwG7oTIiruJ9ig0C1HF9SLb9JSTAaOoPFVd6Jx
yHU0+FiAoIyP9T+WNqg70+jYongdtLoIeITGjzjKvyV9uFSaWATZlgzH/5dG1kF6
WoIieB9tWM9M1RJHFOPJYrPeoZJADMjQ36eNc7XcREL7dkCh60l5rOxEsvKwfaGj
Cr9pr5jmpCuitu9UdBG5piiGcz4BTAcwnc6XvfnO3ne6kVe+NNKj7o71YNwYzkrr
GjrwTHHH6d+THGdY3uqZI07OEIFlQ5aQLmzeLBpQoTvN2SVFVlJcFRcFLrpEwVc+
7drIgMQI9RTIYQK23TOKcMcClxLpATWsX7fE2+OATddUC2UNwX5kYnUe/TfQkwiW
1+oDh1bwyiZrTqABgC+pdss2vddOo89/EP/+SEtzREnNS8ryDs4SEBFhPKFFbEBd
5U8xw3JAAbZNGRc2RJm1add4VOkbRzK3DBs16woHQ/6jLplblr36bH9sm+fgKOoq
zx9Eb50UYjNnzZfmFGEv7qDnWfz7rnJIshPFGp6S3IHYvdsiZMU7HGzVYbFACBoo
Xlc67qiVKt3giAZFZxQjISEOostD3QNN7tHxkmnX5HvRkpgYzwZqDknwhW10KJWM
d4rfYVrbzpKu/PNaJr8rKWvLbe2BTZrkYV9M2X5R7QZXES9kCL29VDhmROTiRlaG
iKpKw6albLqUyHkEM2pzZp+3O0Uj9ne7kdr6mfYmuw/nwVBPlPTFUNkyHQbst7Rj
fmGiYmTOCK1QF+s7xOdQjT5sRYrhLzHo7/jlyQvqjCfnMULqA+QjGf9evFYThcs1
fsg06u0bofehu/Euvb+oyq4iefkCNivhi6GHsAgCBmtnwEucZUvK+J1I9nODTOOd
DAejk7aGGIy/BarqEBIesCFASa77xgy4Y8W2HDWLnrX/awIVr+bOC5QQ4oJWQgdt
hjxkmam2N2QlyLfMUTxdcsYcAc1KhEUrASDxWK2Xe87a3B2hw8/3TA+8Eh4erwvO
4vbcLA21Q+5T9WlN7UVdbUGPnH4NMcIRQRjwVzE37vudW4hY+K7t7odnYkEse2GM
AT/WTqL0A6SsP4bK3W38dY84Pbw8kPInBJaEHl/5tQ3Rrwo2ZgoWaQX4iyZ4IGlF
xjuK7sdVCXymvliXaVUqFz0adTE6QuDhSWVPaYz90Z/ipc5fC8/YcnqS1zcS26jO
zvVbHGh66Oy9qv2DEUKyDpJ5RHaWIiFPqB+6X+zCOrUP0TS/g7Mufzgg1hfUHM3s
0VLnBtWEACDNRtZUqzRby8V+EbP4QfxR8l6VoMrMDFujVQ5GYAitHt7AQD4bLBDc
kOe7HDF0yucgXKj6syMCl+mrbc7LD7O9qMIPZXyfTjsArfKxJqgXMdGZP8tfo59N
Z8BQOIWdgVjGNvuIZaN/0uvPyeZYzfS7GMjUclCQvrr5wpwvhFr8noNQBDb4nKNJ
mrMqhifxC1TdGQWLWyP7lqOSysXxoyAhycATtsyUTYUyl10FF3QJuBD8Kyubv7Us
A6dhpWEQMzEQDdeGmd5MmXIee5s33hmPdwu0W4BYD6LS2V5MsavAiXeDkfGufYge
Yn/d8NoUnl25Gd0ArQDLKToyofW3ZNr7yyXpLpHmsy4SFQJOEEaUw0ahEK/k5f8X
/8oswHZNpUGP8sLQr8PtPZa6IgZOhhdTKsevrok3Qoy1558N5WAESOSDIl9vYtry
fFfmrxH0IBNfPVpyqTw6dhXj4B5aQFgelU2FI0Ee/9OkKB+HF2scDe0HCZ+B2Ts8
uC5B6P/f5VesicYzyrjJJPto9wN3eZi/389igSVDYW2O9MWlLC8i6P5plagjszCF
fkUUkb0AUjL0hWzVp4XjCwFVP/G7ZX4Goxs871fblO/G/LcMUfA0MX9R3tKnw2p4
xk6fjdvnHoh3oaYjZPDvf+B+Ap30UZFUZRK5xmYglftG6ORBl3YxspUQVHUY/oae
Y4JLoe46SsAKVVOPr1KpGGE+3wBBQ1xm2ltDOOdSf3RQkYEY5PEU354Azt60QUXC
U97DOs0CLve9cC2u8DMQia5IIC0mo4Hr9zMYKpEhpPEeGS/TLsWfhtdtJLKzlcaT
xN7wji4qbWJuaxXGulez74RFQdY1dhUUfFwPwt/94okSJWyaH3/55ZTy7RhcVp/m
H4GAK3VLbMq22/ywIZY0OXiqzfY4UOnsg4rATJF4EVc5XgBAUfQha7RmQZNQcw3y
g+xs9jC1zg0UbGdh64lY7PxpFpJQoP4zNTsRbexZlCH4O4T/cOpopLmk8R+zL8KZ
TZ0pUBzWhtYeDGUvhlexTiRfwdbGlC1KDMTW7xRwp86AQMJpxT4oI7wlNsHHnZRI
BAQVnDk2+TACA8ZlOvr2BAiL8AravnhLJOOH9L+u1xsdauXE5MGZmjlUqgv+WrdC
FoBLno1ZZ1hw2tP/rbeLhdLmIAKfoBMjfG1igA1bZJbrXRAJK0JSSYG+xifnIUz0
8yK28Hp+ovHd6bHRKlGISHzh7KP4ABaiPDTn54N7RyVcF/81oOz9Fg+/ZKyx2Dov
SKblRkbacfVRy3syBkmABjnKa4Ic8AfghcYXWtSW+qVZOM+43GGn32QqOI0j+TZn
rjOyym4ung6jG7OyNDsZt9GWk4mfFt/AFMFzpX6zXrqp8I1soGw8NmXfaTd8LOtW
A41XwbYPc4r1lcS6ocULPbN3/oPjhTsji2VW7XJ+Z4acmqzq/dNmV+KywMUPYIvS
enGuDBxA2ikXRMAU2RJH8p94vWWb5kG/Y2PVgvif92/3yIsDnwhBUApR2YT/cQAL
6XZ7UwhsEaPajkU/Qk/drA04DDSxIKVTUJ+pCaYNPL8uh/A8vIFL+hvGevoQg4NV
Sm5tEKx8ZLFp/8i5lmCu0gBrfCDYT0xbM8zNIZNE0xMDwI5RSHTjavLQJi6KSApd
CsWQxlV8C1UeJSXRw0Rbf6nFLaJdGPLIOusRYwD11/tWR007AAZr4+YAt+qg7WzZ
O7tp0Qgxi3OW0SU4iOrfNgx+yoQ23GKqUjzP8cF9wVlFbTu3PyaNXZxXobvGTg7F
w8MSukzJT81c9HoTAhE6V5E40WHohPghiVgvOyj9fXlNFkOVaC0aO40i/ogLvH4K
/dHUIBxitUhjXJnfPpClD95mlorYbBNURv1PR0xhxM3sH9TC46YVA294NHdCZhQw
hsaDt+yJbzejS7UssVyEfhpLCK+HHnvIVEWTLN+5rIYgf2Yim0tIjPL81XcFDFv/
KykXW1fyCYK4DCz60X5myu+rXMbLCdpu5vrli2H+6N/YVSg8Xr9B9j8SWjkrac0w
B0D9es1ATlrK70Oo4/svFGUKlZrKb+gCrDrUSV/5s5RZdEu6oJ+LCcLfvoU1iqe9
B65lPLP2Y2aPnvZYOanBxm1c1T6IX6kWpiS2PGVx4qMWR95xWrF4WQiinDfIv3sx
m7xnI4XIQyhi/2e1Sxpc2RPRAcu4vCQf/MGfCfzsZayVM4f+QFdUQju9rezrlkOV
mgaXKtZxWEwC2bgNUyFx4Y8mJpD/I28Dvq0iNyXpE+ly1jMI0rnIxYOPTlkoJd98
wkkwkQcZ3CLc3VNo8hv+JJ4mvZX0dCISk9Hok2AwRSr4E5IQv7xwDYOSjR98bVik
/8D7eBlXOFBCubKA1dih0l35eepHNvkmc85ye5di5/fdzrYX1oUYl5ytRWWPX8qS
W6+LNeHBpoc5x92qTc69YBs6E8sckTT6S4h0wDO50PKZYOn0nUvGYRUybOpKl4P2
VY3afEN5H6FUi0uUgKWH9zVsGIrpcQDsrq5RNOUYmVQuAXUtJom1Xzj4WfhUj7OM
JMWagbtEfykutKqjdW0nHYoKsRBDgVIjgYQmURyYMYcVe+OnYuq8eIHKBURQVGWZ
ZdWYGxXDGO8eOjiK5943qax+IpxTVKn7w3JBz9FPd3xMJxkcj43IlOBDaqp331jo
PQ0Zk7HW/paNGqQk5ozjbkNIgnKVbYamc9ojl7YQi7ZK+rx/BVPm183dQfIdqjbs
kU5O6Cuo6QBN6UNJW+l5bbdvk6TTsb2mv/h7/vPi2JeAGnyxFbDvgvuHJa9rt4IN
B7BbjJ+xht9kPTge0XqDWoNmXvaPLbWX7jen+qTtqTa5oecJ+J6LM+ov4S5ukPKw
VgkAb+2ZvzLu5yTmjYW2aUvH19QxsbDYFV8y1nYNWeCnd4MefgRoa3xDwzR99ToD
cKa6nV0HEXB4WJaEtM5AtAeYgGBZZfQSqkBmgFAevwgE1E0vQx6XV/7ppUzVQJwS
qNYS3kKHh++WIY9Coli8xYQf06z8fqGplA/ODXrno7ksHJDcJO8jfhakyNKFFAce
R+u6+AkPqfVTFqoTyrrBe2xAQgT728FmbChUNiRRYpq9SaWUFcJE5HyxAiWZbzzE
ND59AfDvQvjuzQdXpetWOabvWQLJnsEy9ja/Tu5cOuNj3EQompIRvg+YkNx/ITck
KjvdZ7yjeR48b6SeospDRgpiOJWAzn5L9yjvYiCXFx752HHqEWTAFGmy27PKaSWb
Jen0pnrHQ+bB/+SfV9k6b9WDZCondk0rpF2bS7Y2lhp37nWqaxDHc0lNfadkDt8x
5ahbaGH+bVy3dzezTneEWj1KSRfsR2OVoK5iuaotDCpMfGjyj8iCewvLL/uP/bOm
f1F4VclBKCGo2V0KUoG1JDhd1+AyapHVbq6mJb8AeishGoML/ZsQIM1P4SPyBvAP
2mH8sI/XoMo1PylyMj1MIDBKGg/DB7l1NFePkzdpLY/TQP2gm91D8l5PWDz261OK
7cVF+E+9dv2Qatr2cZnEj4Jtk/+t/G1L9/0gPEYOV7clQbXtwX/htaAJROEGRVev
Y+i7etPa3MDK524abeLI+MJwTU7lSxnU7YMtXuMwEP+6IqVInZp/e2HsInbi2F9l
nSV8QYw3Qhq6bj97lJd42zmgZOBSxi4GWT04FsVonJQDls6dwDwS5YMVtCk5tAGs
QG4XpJKAREkXA8kMNCfFJSwTe9iJ9yUWIsKZWa/AsFH5bAD5aIrZZhdsk87jMQGz
kjVUakEyuk+qr9bM0vCxtj32PUyzQMb2uJgHTGAUYakwfHkH34flXylrS8KAlGsH
7KLzwoMF49hHsK6dJmaYDgVtSzxcN4xabs7lV8qS8iM+gw02+Zx0cm6f8GTlmhQ3
NPl+sJ9/qK99JiL9pjAjkrkVKNFx2QtEwSPG504N7TXucwiRDecBbILXcdtCERNs
l1S38CtF6IahOfAwgZuG0puSVXx90BKwnirQrxeWsxD3USVX8xIjgyVTSjDrcSSD
4cqtHa+47Y6oXmDTEwZ3BAOQbL3FcfWKdQnr046gpPDciVBedDZcUQEKXqeOIiIM
UcGwqehPAE4DPPGigyMb1UOM0alU4WO5vQRgWWD1saIubsXGW4L7PzaB246koYG1
6Ctk7ghMmUAsp91KgFR0mAVkLJOc2/5e208G+MDQbrGBEJI4iNoxa/vpDjI/z470
YyggbyqwdvozSLVFQ9lI8MXyAdtF+QR7v/2qQlwDdDa6PKAVlNo26g1hJaCmCeQF
pkLb/y6JCCZOgEmq1Ywf29roF1IndcpyMwa1YP1j6wD8MMEd+nnBQVaGr8s3PqUi
FUHLBHiMX5mtPcnfb1WbpdwjUdrumkdwriLfI3rmq2VT5IxHpbxGuIDfJ3lIwn4h
GNy1nPcDSutpE+vAc62AWH3HnghEsw4PIEAR32gcY1IwfzTEOmoqe+58AK+OjAfv
GIqmAiYR1yqWgoIOIuaPxhjyAumvuauWRYUoPZpQ23Fx/sTPK+IuzyeEyX0CL7k7
cNhxMPm70yFvhnDFObrRX5vL/C8tOCmHzHEwhMaTLIb7pRIxhhi/Qhgy/usfdBNR
dUo0Y1+P4bFh0k/jt0Dabt6LLkOsdntuNOWnhf3cUzveyp8i2eboiwuPY+DZzpLw
g4/OeopTt2rJIyU/EonBNPSvVl5TzJIpQNwz3gF09Ic3lQ2wOTv55vI+GCLl10Uh
nFoynUotirC+T5sl0KKL9epTV2IuF/UZBpr6v1XiuCH08fh7vhQwRkbP+ING4mRU
Fik+fxvrOX+TdelIEXU3SKE/d3dZIWjK50rDKLTeG7IUJjchdf//dEwAGH9Yapf6
ucM+Ube1JYFum4RfW3ALezwTISkgMXKs9yCYJA5qaowbm2nyt18bZzErW7DAz6ZQ
9bYzZETtTCJaHqCJdGTh/bWkrUScp9/px/rmUYxKPlo0lm3tsDdjMPFGTOM3Gglh
K7OqyUEcw6mGqAGEszXBPAU8kOhPmICOFc5YzmP6cAr+NFCEELaSe7OfvEBtaDZF
gMSY/iENVsP+ocvdg1KU7qotNZ4fQtS/lltu6zZGmsGQjQQGlg7pbdc/OBYxDnS2
LcrBlxZeO3gIYkCy2T5rVxND9EnqqOJzlpiIILCUO6sEit32vAsvzwimGXJVGdUA
7pfayKxBOJN0Y5QfT288YuKh/UeNMB6gJNSucHNOUTlYfZ3k+J/ca7qhNuluVlqQ
m05U+DR3SfUXv4hVDenwyx0KrctU1pONRfsLcWmVm4lYhbaz1X+gySZ5tskQOQd4
b+u+zR87lGDrKda2mUL0/uIB9fm95ggCxb3SIfxYBXpZ/Sq6Yi6ig01xcweWMUo1
px5jteVsRzoYPtx7erfDFFR613DvLrYEXzLy4IylfaohL0v58xvfZhrfFExKWhBh
3Pa0tu4syjQy+lip0b9qTAd5BGw07ocqTPwsSBuo90sRTJKTM8R3zioXy+5BWLGA
OB9sW9wX7jD6X2/Pm1XYD6EQ68Bv0nNH81Q14yOJuaiZjgtOG/zCeXzQTRZ38LKY
wA5mhf6QBe5RVKyXSvEqQFDVqTFy6D3HGm3EOJYEo8TZqY1aAeLpGk0GzMhOia9m
bz7tSaR7mu3EzmglHPPh4U5LFbrXFis2xSV6dgsGfG0JDnVRnLPmHt/6AIWANV41
20fc2vQ+cW48jue6HC7kbuT1xYzn/NNE/+UOhUUQ3BNvNaX5Ko+dewrHlhdAX3TV
+AOYiCBmF0NnbXXJe0sf1v6U1w4aG87/XOVnKKMHBgkukLvDUODoX/Qa7yP8apjI
UA2bGlAxw0iX7Ci8WSUpc3ANImfu4p/1+TZFGAaYJXMwn0Qx3qaiUwK+QxSqCCya
xu0By+Tj5RvWBi1I7Rl6Bx8A7q3duvEMEhCSpk9cJ/SpD36TIZ9xZRiePfu562bO
u7Vgp1iFJToG1wsgQHLED4PTFothAfhzm7mqhohSDxSH0p9h37RR8LglEDjG4RzC
FvduKiRHw7k1M4xjbd/S8AXLkzaME966puoT1zeZjhyQs6VgGAGrZv6ewxls7zoU
D8I+4zwAR/ue9XbXwPGI6RfUL6JFzdpbRSd1r/0fJE0/WEkUkjValM/MKqqT1iib
hclipCkExvVQ+zPInMMda8m0u7+tnMJhzX0L/AnfP45np91izR95Bg7axpS9PcdO
VpSKFR3bxRY/WXUmhs+w5kH3xe92phyGRyiNSjToBi4+MPCxn/ZgQlP2Ez1d620v
c8/nOl1a4xVm8ipl7v0OpzZpt+EQgG8OWwC1juKz3+tM2sIrOknnAitVD5r+5h1d
3JRy6LVqPNHz1WxS8LxfW91Jxiir2tmwR8hR17HERT5Y4fd7YZXDbeuBZvlxvl91
j9iA6W1heu+15qODJ8raOUxrv2eltW8xuxDsbyaMP8SQet3wbmsb0olyj10QQ5T6
Tr20Wia8MRuJZmJ/KoNKKs4LWRfnqSmQAjj7O8yo3zWUquePUktOnalG8Lao724k
NBepgAk3bUqQNS94WH68DVcC4yQDFdTqPykUujvjhbC0U8PptmqQsXjty3JQGwW0
UAGJhLz2AhTj24ngHhggNELLV8eifCAanNRdW5CXKQXCXM0kRtFObfL/PnliMot7
Oft+52A7zz0sZvZQCqEKsU6zfCtR43rnfWZxyeozm45bqrfXOVgsp37oVie+2YZZ
5cHjy8VpkuGrMSlMXyh6dAuqnk+05psiB0gz36mDcJHAg+NDV+MrKG82ymO0bBXt
N3Fy2FxCJ/fdBvhjttdKsgpnGbyv0snO+zAjO3O3rxynFf0UiN9KScUY8gLXFrcN
t8FDXE60soVQmWC71irAxU1giofgXMmMgnj6VnbT4qWjH4oVJhRbOxDUA2yav+vv
ZAl0T8IsMmqTpOTMQYnB0sUpxR9sLw/NkcJK3tMMxi7JF+aZ1Aa0YUswO2qR9dpy
knCS2go89j2d8B1Q+jB2qP10iF4L3CdPP6ZZDEjrSuf/pfPRK9ixB51YHaj2lqEO
lgvp253mJlBakcRrwx0T0IQPJFgGdYLm1g9eRN9T8zawCACgiw02nXmA948V9+0l
rI2IBL5jshw8ZbkBO2bSUzutJDTMe3T4oRCAIsQHIZdkTxccvgcWYO0CfXp5UkY0
8Wiwpv/vcMRjSMsMXOUQGT6nzyieRasS5+0Wtkjgi4t21c5HKKxJ4Gg5EoULWFSc
9f18XjCly/ItU8021AEK6O0lsgmOqSV9OLgZ0EHs5aTNp5lhJZSucHzzRGiJ06lo
u05nU3LddswjaWLac5RlJ7UCHVXC/NRAzmuetMZrihY0Bo2o+DmIGRpylTylQLj9
w0rp9X388S4eh5FZBfcWVvDFY56liueJ20KyTIgvVGmcWr9V/EnrMmQm3gCCd1kB
ErIyHYhpwDt7lqhSMjDo0GPv9WZqLso73x9uDW/yYc6hFnEuc+ITPzefr94q9avr
+OyPrNumrMhQicLkDjqIdAs48lmxNyu9jXCHv9UxriXv109ieq2KO/DMdEd/Pmk0
rhJimVxpGGIW52un6B0dn9apNJOPiYmjiP5y/3yrZjcochKLomOoTdBmUh8Y1cXP
fZWag/SZE1gGs1RiFQMTYvLiA19CkhoLSAKyH1kz5XUaXdqb0f6QnI4bU8Vt2vSa
Grk5djsLOivlzyowhCTIas1X27Mmey2ztVKMkQcUqGYpr8qFUWYW1101PDP+I3Mj
rURQzwqvXVmhjjWo7NQ5aP6PS6F2UH4VYZQBlY+KcsVfzE6NrCWUW6UtXmwj8vSn
SKjXWzg/13u90s+R7EjzRBisboJgmAnZxrrk5bHVnMo1XPNMyhIdhWX/O9jsyAd6
zzKYqaWE1i/xEkxVf4EO4E5QzXlpOP6ogekyHzgwPDUjbiCcQifboWsRCh4/RPfS
XU+2WFbMiu60Vu5i1sjMRGnwxWgs+ydPk5QXsfT+IcCyp3d/1ElJN2HLCD4GRXYk
yLwIgimS/LlXFBdQ58zGehWtoBOeOBLrWROL93HEFDy5+pzH95XxVFDzijpNf9aS
5o30Drow+OIc6q/cAR008JU3K3Ugp5wobAyS1EJCR2L0wJnhy6725pxF52nVKygt
lk2TmtzLaNJj8f/pyHTq6wcXVSFVC/djrirXOQY3K6fU0GNJ+qe9acRhrIkZ5oAF
/lw1m4ny53F1IUJWRnl54kbPMyj+T78lp+XYLZQgnzqcSvam9Ws5FeQLFp+OuQD2
3QeYdl//A31hBhv3B/fIr13IlUEadzdOg9EVGi0I4kW7Bj01fP4NR6Nje3dtT+/M
D+i5gpZx7inZpQJ2VmmjAZcyeuwu+dVWHm57qtq2yy/sXvmDmrmBqT82x9idigVF
nz+8Y75phmMsXgM35LTZnemzYlYBDGJoTUp3CRTfj3g/MTcGJyOOLQSvkyxqAtZJ
GtXQSax8pkMQNrT022m0sAt+Wd0wXXQeREDAszhSKJF0vsslwbV7dGqSxqcNdor4
LE67XQdd02iMLnZJkkS0xRpdcd4ucnmy+OCsd8DNyo2g6vqwULYpPOYEkY8BK1YZ
AqCZKP8X5yAAeKIUWrCLxXI471iLWXjqpesnKYbPBjBYheIBOS7/DKwimnj7NkAC
Evi5sOM+DZTKQtlqqneVxyZJ1xS9u4DFeEYoQAdzoe336etsLote0MCzb4iTKA5+
MBp9/gxKpUSPRARpcChmovzLirxqDEjCqkpwuTSZlwTcUH2S20K80YGHoNLOK+Rj
WYEA/m9B7rIeON8NuyxNWn76k3Ui5Nj3T21jbwAsWQG1yMRwemOa0RxSIHn91/3l
VeVwrl9zKhIEAcFiFkqgxhrp5P4VIau87leVYFGDtNRef6F+AFXkwulDu4q2Ebhk
p8GaChcXehsANmZuJvrdrDLpK3m1KcMSC9Cpqwb0TozPmLICO3qA6TmGPK4UEhtr
cnJSXIwMRZ2PnxCMFA9xdhGgEaTGB5ikrSex5fGGivQ28CzhwGmGCz+c5MX/AVI5
e8Xl5LirYfTownje/AXJOKD4M0pH4g9n/BAxssOzX8IGStiXmFTgkJKMZ1ZF3CK7
3IwQEd6KE4RJ9duCGe4bCQyogzmUAiOk1x/NiM9AciufFehymKxWjEznGGUwIPXG
or0DtgY/kukm1K7Y0nIQY2VkvYYywUfhgwaVvWo0LyHHTqW1OlrdFDUK6MRab1R3
A0U2vj5ZKfkGtwwRSSZ4++2PzUOug/76KP0l/qqJAG++Cu2FxadxqDNfz2KYjoD9
nOWkxnDks+jh5/0h38tKRb5Yfxd2GyQe/aW4DgZ5zh9SzYfHqhauFxE8R2QX1b68
8tYdorA78WnT2QX/F9DfnoDyYMME7+ErfvznsafbQGMABX30a9bbqk73yl2zIYDX
npbScWh39ubvNejI2TwKikqZvLmMQPs5p8dwkHriaF+yEpGKqaE5HdJt0kcvMkxz
OuaX1e8gT9sXNnLzJA/pFPHTMJu0Yn9axKoZjdvpO7g/VM+SyI4yfW9liI32EFIf
F3boqyII2Nm7lt5w56AMftAP7tK/zW75+Kqxm9ufcnGZePSTVNV2lEUZ7Im8Tz+n
4w158o9p23smp6znwE4aIvt8aN/sZjmWwKDFFvysN3/JNtO4hGc5mZGfTLuXczfi
C4TXxF2GpSH7mBQQrc7TPRhARp/9S37lpVXM1fmoRo9W3bGI14rwFgGpqKDrcV6o
3Ay75sIBlZjQ9AHgHVQ4c3oPHG9uxnSINYVv+BWH/aeU/KJr3tAkS4xizl2KiOo8
UjUPpbXNaFp5jlXIxAt6ppbxEPHfxiGVUx42rygqI32amKhKJkYd+ZvUQ2K6GFc8
uF7qszHq4dVFQrSM4cO7qf3vN2F+PbHCXWpHzFYq04oF5zLolAoxkexgjhWdTAL+
rS+5HY9pzp+dNy/RbeFyJvUQA+hnsXJBAjzbGKWcwPOhJ3cKn7gFm0w8sWfqGXh2
a19XEJU5XuwQwKIMr7tIJP1yKN1CpyyedLlUDFdaOU7787W86zrnTldc/iJh2+dG
P5xoTAN6x0K/7KolGrTSJUn8lvO6HvfIUx2sCCbcmiQFy+AiYd4YswhH2rPSQ1LW
wIBd6NNB5lZD4nrsGbPjBK51BQ64LHcx06zHkgI+KJwg/3cRx31FKpac9Zcij2nX
NW/+u79T20n6dYIf+Z8KA1q4C55T8qPW1lxIdom6FejoRCGALOtpTUB8AZHZ2FfZ
nUu9WCTRPxMY7ta4nJsco5KwHxaP6DZlSZ38c1cI3YZHzpLbvocw8x6RyCOyb7K+
6fo72qBbXj/gcuazlwPCX/dihE7562Km+jXQ5mLa8/WSh8ZgIUhPFed5WWlWDt//
hA4pVr5UC/wsVkKwBpLaICgcO28k3GHl9qLHY9wtdERVKYVP1XwSgSM+6J1tXyxu
nDr4lmQ63fTEOfcUq00n5Tr1tZB6H5Q9Q6NbVAy6sHXtsGDYaU3sVu7FYK64IfqQ
+lbIq17L4GYF7Nqaiv2jiPl/UnrTE6km5x06VYv/ESoUDork16Okm0putKFs12/2
skVt7Lz5v7uZgPeV5AuYuS20aoS2tnoPgOYW7iGa+nMKYQApnHaMBk67ItSKBIV8
rtIE54nq2DPiYGs0YdxV57xntqF1pTmQwgqaRPxF9wQYE31K/Bn23dzm1RnpEX+3
fwFSjtRknd0QxlSvb2w5tX3mRKWv1cBUjGEEQs86AUJXQmmt6jiK8S+KsOH99Ilx
Uj1IJ4Z9m95Dl9UveEmsAbkMF1Jly3FUodbzXgIN3ViaddrJXBdqf+VAMLN8c/Zr
kpHOstfscrIEjcARqriavs3DDTeUY6HCXw7zfi9Hc8gsrsFCmB5L3KCwUe5IHPRB
f6/k9JmJK4+EgXpttbdjMhUwxJEdjdTEk4WfoI9eKjZ7PpMNqF/oz8XUTtPlK3PS
g5IbPEkMRtZcpW0GvJlN79PquR94t4O8nONpopJ+2Nh0VUBksnbBaFmGiQEAyiev
HQnXzxC6W1hW2SUOZXl/ZhjwxyEeLgc1iI+h8WBk6rgWXw+6OQzHuxFYSz1Um+Ak
k/+RgUqvrpEBiWhTqsKF6j8Gb6/naouxRtv4V4kpxWk1B+jaTiGxbbRja38+OuKe
za0TOLmofqHRmJzIf48a7c/S7eDvl1HGT4t0kRlhxufbHJGcJ91QTibxOykGaqwR
b81NMxXTUbEvg3WVMKTVjTNLa3GcuthGtKyaeoWkjCPKLtLXnddjl8LYbH3vvA2N
k5lPyi7oSB6CL8yUPsrqWJc/5o9LgykhxD8gaexwbDaMJCaUNQjMFuHbdCLVMDKS
la6uzuPDRBW3bW5vxeUZPTxKIUM+lV/q1WnWfT7+ITRP9apRhF03CeTmjXAlEtiH
Ft9XlV26FAdKriidTVOCt7Yw/IQHUAQV9r0STTEpGtst/W9/GjtbX5D8JxRwCTun
7/3c+q550nqgcxz+w2ydizbCBk6GfvlXgHvCCps1hWFrA4j/5ZV1fV+uWZ3XuX89
lolhQYJ+GlWWguPHZPAgNkNnhPJqtUK74bZpxrEt2eSG5ek2xdbALZTi6uXWlH/7
vf0pmGG0hs8nf7esiUIN/ZPGZ9E4Rqq9ZkD7dbWXf4RhIitWIIyPOSLHGs5EAL2t
8s6MdFP8CpzPmcKQ0JFjEfli/m08uEQaOv9sTeLmumjGO8GmXHJIJ4gX5ASYuzz5
sC5yzKhOZ8qPJ9+tRQnMNLuzBfxe936VMre5Kh4T5D+83QudmwIIkZhEdMwE7Uf3
8zJjsvGHWCZPsqynn45sVRKne7sK5xjF5LvMcme+0UfpGgZT1TUSvl9zJ1ejgT3d
0eg76IG+WZemEpNpmBDm3ILAzwkpRlq3CCbva1B3BGVRAHtW6l5oKZrCBhF5krux
TbQFVlGbH0mVHdPrmdqIWZ4dSA+cjNuc8ekiZvro5BmRpOM/7Kk4YCf5KWPqpoFB
BCeWEzmIxb9pPL3kkgrXDBciqxxYyTBLBUKVZM2cpISYlXcTIRU4BrFIqIapFetn
jgtrIrdZPlbwLrVnDETHO9Hf/OyOeGLn1eaYaSXkoNbBrHyXaK8RmoyO/PYNluCh
NzfMqPulHRwTU/WmOOtQhJTh8qYbMQW5OfjqH2cJKl5O/8YcminwUXYbJV1MNXU9
F1wBUn6+XNuxlCI3tU4fv4y0kIeBEU6EVMJkFTxh0JRcZItVdkgVliyF6nEoFVSN
/h2HDYfwQeUNxY/NenYRVqkVPOKUEvqwrV/Q0eZtpV2oY4kqUcw1pN6JAXWL8HF4
BB5YlnhJhIbtgT0+dtAs/5tkNOi9X7C8KclJxqdyI52uHctDNltUQ3a5A84Kvgua
KlfZqzOiiXY4JBgSi/qYIaYYEuMrsSr09jRoXiajqitYuK8knumAQvl4rTRShAiE
M/5+L+P0vMbfzalXtS2T9IbprjbsCQnzXTR5cF7Lvokqx3JDREn2AjWK6WC17ho6
0XpJkJtTabopteir7YXfTSwP6fX67cXS6WSvJpr+QUO5WwJISPDQJ2ZTEE5fUHMD
9auGfTB1GqWaDNCNxrl6vEeuTEdxerVCBvvZaBvNEQivxpz7z0Gx1R3w97/MYJcB
5BLY5zO7cX9I2ZOXfz59iDIbe3WQcBR5mhdTrN0P5B04X6hQgmDQqGp8n1+KZYsU
bhHy/Ar5aKXK+gmMUaa3f/b/LsDT8WmxzleYOLcynDske1vobTyeRNMe3AQ3U4kO
Bzw7vD168IlTe1x/RlPvgPoIi8TMIJoPPCDLSmNK/phWIqBxzaWA7Ks/c+fRDjNV
0RbiE9L1V++DyY/AfRT/dtY1K15yCth0O7VDF5XlD9Jk6euRMM7XVFm42HYnvX8X
tzwqpCitzMeZsSzwrDrAuadzybEaYsMtE7kdsy9x/qhfS46Ns63Z937Hg5uj+cIy
may7Nl/jpByDBkfQdnm7abKjqPchK59hFOG4FgQxNyL/gMSgD9MNai7nTYGgycYg
bu06zAvzkhXJEUOdzW8AQIm/bWTHTElKyM8gr3nNI09tzOqAI7ddkImrA7fkZjA2
QWkaZbrNBNAKvdx6qni84AxGj0NYnpTN7/Ssus6IhrcMGRgrWpjOT7JBzt2An3Wo
9lQr21FrAkzKsQ6CbTeHtRja/gyDf1VetEhbwJCoMFkUn6rRat/cuoRDfiIqb9qT
V+p5CdDfi7zf97mzpUzaJ5o7DShMBGGDnWvlG9z722vc1xCA3M5rfKcNljxfOavS
mllFulsT3ZGL08ftW8i1SvWpYw7Q31hxylsxVga29L6fMJHolSu/m77IVsGLbznj
eK8Os6V16t7cXQfZtjo40lgoCq/2OyyJDUBMbq3V9EZljIasb6vTPmcNQ7PGq/A7
6DCmM7LWoLB6U93bAG4EvT7IU98gquyq29aYNpCYYQ/JLtBrACHq4Q/zvPr3POJZ
xv+kLYDC/OOdSTsSAbIdWSSpQX4ihcI23+pCMBTnYTqirtsNcjuqGqKI96q2w0c4
atpeOent0dUM8bfBKq6K/YZjRYa0iMrTGIL6p4NPcfML289N32GzWyemxZU1HLKh
54S4R3VP+50XoCqtLtqXi8AHuOskztuGwT2gLKWuAp8n0R6nTq9HiTE6bTMf/JKO
i24DGu3/QevZ/rrpYfop93vxlG7a4zocVeNYE/bJMXNYQsugWUWpByW8OnjCMvYm
sTE4u4rnvbwKGgN9MoJ764H/NKdrG62TJIw07aM258cTcaFaWEKzg0OxPySxYNlu
Qio6/uKLr80lLCraQrdXZg78iWN6b6h3cycvi/Co+eUwKcN7RAz+uPh1N96dtGGU
8cOg/i4Dkqdv6AFEj+DYCFI3cyMPmLO9BifAEqCZVENosKDV652Tj+KUn1jSfr9T
wXjHFl9FaHv/0aQOgfRNkq3bHbEIAXDdwOp2taz8XZ3GjmbL5H3OBT1lk9y57eSw
7mv1d5bIatPrxo2niiCZckTEQChP5ZQQTr/o65wc4pguu7+cxi/aLjL8pnFrA9Q2
k1uqv+NV4O+s+n/qCOBzSN2WPRUg6vKZABPhlL5gWys3KllSIYV9ND8RHXIe621D
m3kbZKguiOz1cMZXcK5mBqx+aVXgU/JXY+OFo+jnmZ8zexVbsOxSAHe8h7uS2TsU
Uao39WPQgewg0hOgKblzData75skpvOamiL9GzRNYSRbcvjhCYXRGlZsvPjsN8x3
iQAi0r4QxFBglDBHfSLwCgIiiHCxPTabMliuFt0zZ0wXSBbTPsSm3299iFcvD7Ur
hWeo7whumVb1y/kWuetcEK5HlEi6LZzIZ2cfmNlYVsbQDLz1deCigAjqhLbms4rq
iXVmf+NdmM1MfNFx4gZVOvW5AmG0qmYEL2FpPqTzgEDPRW2JS1ovcwdGHRt/Va8Y
ud7dZ+yV20yMY6dscGL3Owii8bY92u+Ib8+mYAiU5R+tyEWkBGfX7J6605oXgK9N
RQmOYKbgt/wtLxhceZfko5zuWYrHLLjvL/rCYmq9vgGhReGqAtwYD3F6kuq7i01C
CMauJNra+H7fw3Y/zXODLCb8QcsWIH99ARc2fnTwSr6uthOgepcEZMbvQsW3wR82
Qqw15xjgcuHH4HtigK4yvL8pBRPEiWFqhoBZF4y+QQlyommb5EWcBTyq05d6hBqT
ULLJKqI6dy9FVtsyFcg73tI9l06x2S3+U2wa2aJJqtJRh0coYO2lM7oWfcsS36Wk
//pnTO5Kch29Vpfivj9VsW7fkEdYM6iptQ/lHYzm8eZkPs+YcCVZKzKp+l82LO7O
qAX9EHztRIITFDIsFpz0EfsiBZ7g/N/jfn4dDwrfQZ70Ct/4yZoJyZVWD4/gsuB4
hBr0XgDU4iPYBCq8oSf0vkfi7SBIfAT+z9SfuCONqngNWLarpj6O24rtWtWgmzGJ
NJgk+CjeOPEna0axgngI2kwZKFbHulJpDMIx6nVJCjfDzksBw6P34rBroJhxBh7r
5NYbh/rw0fRCYQ5Vy+9EFdmMVTALiordd3MpK4TvoCwDFtISrMbXoGOgO6ROZbe8
vrFj11g+BvKqiLBjohZ4/WMMlpO5UcfHUI56nObAUKta3Rn2Pyf2nT3EmGnYov2D
czX/XaBB5JVa6rK985XeEdeB76mgOdFq/tNgN6uDXoHgQKleg4LDiM/4I+YUZChO
kyiZrYj7YSrhYlYmGpJBeba10mFBkEE5uC5AnmJPG3khD0cwd+zCA/g7IHljYIYr
DasWqzy1WWHC8ZbCCOM7YCzN7dhl3/601+W+LrZxw5t1EFqp5GYCtuQYOsKfy8EN
ovrrzOxaBgmAAudJ+hac8BME36xhgludHqZ1SaIV/xnSCY9ExbObosJZKMyoZS8t
hQl5sI3+KcWHTSb8UUrSQADXNeJTNTCTKlpQkDgmmmK5kFYr6qv1IGWNNJGuSgd/
XmSerF4IeRF+vX2h14lFKjKYhojkzPSBdBECRN/enVhn/Ix3UxkePipfUyIUmpwQ
GiSS5QCtRVfht8uN5N/T491K08orPMkr9qcYAon4SxIso4YlJu8vLSN23SfVwDKO
0cnxntTAoGSxb5q0ZKHjBVevfaB9ZusgKI10x5QYDW7a1qj6vow2vUJKdQ0bplNy
KdqDyVh5AsEl2zmVNjvVxd9dOKUm8SqzSC+8sZnZxZp3LQdkwXHpouB1XvtOWYTd
rxCP8PnrM2n18BwxNFPhGsVTZ8yIL/Qo6ea8Iv2+8m1kK06FIUGi8NpOXCGj88lj
2QiWo3eORfWgHMGI3iUtt6kVQZmr4kugP7Ie2eD9/41csClJYGmFdIubH148hW24
hjKa5IS1GB9KdF+LcR/d3EXO5RMdDxRXJdP4O7hFys/j5bSsbgxb711KkdTIOcif
TIXUvJP8jvWM20LAkAylLTphzsf3J+4saw63uDxx5MrcQdvctaS/hEZf72jmKPL7
/f1ANk5JXLv06zHqpyml7FCrpMDgBfCwX1rngti72LDgmoAzUAAUJ5aSJh0xqK8P
kBDSiGt98PE2CBYDyzCTtCp2sePkQgJpuwzHADQ0PCDxUiQdIWgm6RUO6TRIQHYG
Ew8F9tGAMh9hf2+toqxIgBH16bqYMfaS9/AtWtmrmUgYvElkZaM3XVBxB2/q8Kj0
6PywjKrJC9ILTwAPRkqQOL/1d1mEYir5FqlBl9jcnCCqxDLj0IrW/3qDgccfHoBI
R3T6syDwAd/vuPYw5oWGXMhiaQv5rPdpPNXkug8b7Zp6fDbMCj9f5jeKD5SUPgqy
gJRCwryTmOHP6FQWdcHo5zUyFifWdZmD398DitkcihQfguybit7n0WT3va8zqe4S
Y0rf2EkoVmf6v7PKqTcj8VRG1+ZFuNAeNyOQOsZndsp1tKbV/Cc1Kx0/R2/tZDP+
Sk9uZM+wt1N15vVMWqYR3GPZlXUYcTKIrtmYUXyKvSaa3eY/t/JAn/+3xW8UWP/V
rUJ864irFqxBBA/EOyv0YnGPrpHVFrMaIh6HHbiDqu2ncmQABecBpXUU+NR/D4Lo
5eyDIITT7AiA9GW49edDngJ77/R7jp2xHKJcTYI8RBB9Y2iuAkKOKZE6Yu+VdFRz
Zlc58dPvj06/wZASI5K0OOrEVaPcRNkWXT7ruMXSqSefme+zwKTzO5Xs8YNEVwN1
h0tvUanjdsVIxTYtvnSymAwbqEWGq800egE1vVAwpIzW4gWtFebQKrGQ3ylKLJg3
BUF29sHoS5lGK52F1nW1wy7/QbF254w38vg4rzV/nofHFYnP3G6Al4dGFbmFOxcL
xao5PspETWtN8a4akhvXqus+T1DjF4TJJm+6Byt62BViOy7rjXdr6tdZEa14Wge8
+Rtq/ykVEFPMnzhWgb26669pn901R9JFw+RpeTiBi2xVrZogIO6N/GpunCyhv6HW
e4kBxnUyMcD04UKtYtIC+mhywCG7LoK37dPUm6dq+Oc4xwb1PFU0rNveWyaX4zzg
zJyRxvYR8Rj+N0/4WO7wfAbUhia2SHgvIw9Ut5YVx24eXRm98c94rJ3IybJ3JhcL
ukuGcgPxmpaIkOmTM7iHrG2Ww2v7X0085btVAJtcZSe+6ovqtOnC/rkU8NDCBrf5
qvct4QOWS6KabyeaeM+wLt71RHT3Nrq/s1ZuIg2MelkWP9zZcsFH3+XIRd6C4Pgh
J+koGDDzdVdBoM0BFY5eeDsCNZ6/1azGKRcbQImSYQBqhY4Ur69ZVrv1xAFUnccK
/7+khPxUBnIomlPDWORBbO/TW2fMgyLZZLQ7QgVLHuMm+jW8C9VOrX2NQA60V/kA
Rom547sAkGO0OKjYXkJ7IrTrpy6ln7ePe4OwJw9KjeQ4BkHzdtdkq9H/BsfusLQH
h6IY6PCE98SaWZPtOogaFiCFMJje1jQkHIJNmbRWtc2WYKgUIHEQS+pgNr8SjdM4
rhvVahtEOmySxThnzN7L5Ku8U8AnmABww9mymWbpUk35OCXRaq+c7E0rO4kq2tzO
ZRRhg+bp44hGYO6FNumBbJR2M9RCEYYRhc/kXuXbPL8gJgU3FuloNjuMM+w/BMTC
nCLoR9MkKCNeCboD5tb2fCORcFG01IEYimljuFGsIs6TWyeAeybvdCe8H4lETAqv
TpkicuDtus4OhilzR6yu5wFiYgoqvGc7+A2TtdExQ9bciBTziYYW+Fm/2kTUOXwA
Hbvipqz54e439YNMPNwLRPW8zFsDsvf4fjDM6e2CXEcigG29FYTJwUgSVJF42vSQ
Trw76uC2dBhSe4XeS7IIjPX60/1b/e4En9wgWh7S3+TZ/0jUE8c+OYw3y1vz/+wW
UQY3sUlQa1v6VB/iE4TPBY81UYCHi3NZ7BwAkWeMTjG/ZCMzid8SiEfkUYfSlmlg
eNmxhBKVfU7rjYwek5TvAlQ+8o5im/hm0dL0c0B+wL5h8+ldLuyk3IG4ndZv3adb
IAh14gDn2WFJtx++O7Za1kqMwnmSW71kWfuuD8/f5e8iaGLT+jgm/j9TsgBIVYmk
l5aEUxzVy6t4Ou/vlAwSUVNBM+jPplyViHUtgC3I+zb/Gpu0OLrETkKywNvmNYxY
Gxj0ZK33ZEi1Gr3wszXRb7iqaL1naB1QYNSmGaFktXwPsu7/SyH7D5PSleNmhX0W
NQ/ff7iOvfvzgoeQpCL3GLfG6S+w/vqC6IHw8d3hoa2GYiekXlsmTg1jy5bMTjCp
75iCoWcxw4WTS5wo87Gqkw7QfpbAE7BkVSfefWSaCoJ7R6HcZPpfpQika3Cd5907
FPpRmA+6a9uLBCpzFNuZshrBXk+oUviLtRMI9MFNmESMYClgbSWOXODJPcVu2E4j
9eO9UufyTOUIzXCCO3LsCQ60zZjFPSLHJBWQzP1OKjv3eQWflFAKx2Jnl3kB8IgA
bdMaDCqzZumWaloYe/gvyprx02+udlp+3+A0UaLLcseuxT+rFDwGby9VuE2+1a8Z
X3ztx+vPJ4J/XOVt4iarZXqO2U6JJGE3Qzi8iY0G4qGiQd8/kydJ/b/MQc8e6LxW
Fr+TBUcdmmo9h+JnC4Mqtw8kSMUXHEo4C6cQKK5sF6fzjD18otACjPFdexE1CtAM
ZZErO6A7i2vhb3nSZIY738HCctP2MsyVJZNEvBc5aOHXYZ0QDcEg4j44hHtMwl8I
TQq1rDoSt3pQvr3pKBIGmQx4C1MT33AIgUzcSYTeBItYnPeEkvmwdz/lqBykWCBq
0GAcqRt5I+G/syO9EvriaR++Kcv30y+P2ivQFjpMN1gPNRP5DzSobYUQIwqeQNBb
/fyFurbhz30NYLuXOHlUiQtkDWIqKWVFGEZJ3gXivYsU084mFxvjfsVNFrAyqHrx
Ij/kznYt5s5mUzi1Vto5EnuCrBYFFleD/fMaaMRNhs4BPwCxCMxijtDkE8OWxuTD
x6+lrzDK61JGn6xktaDWjKKHEM0xqdBvSUxVFtmAcHixu54rE13NC3h/u1ypLWxl
U8tMomFSuEcAFLDoRNcJjGFLlL8Ef8q4seAmfMt5s8CK7VbVCCo+B/BSfC1hrp9u
mlYTcgp9hJ6xwHgLuuubay5QKi5nSLeA4TKu4Ncq406l4Y9N7acVTq8nNHcPIdQ1
HykCFPbLXJMG7Hh4gTz2d3uCJVwvfFG1KJDgYZawNHy2nid56nA8LwgU5OsOxs+K
T04lnMycMIjzW4uLa/wBMRXXe47/6QYAR82SjeoZNRLv6AUq8jvgmytLikbTepHT
A6NqNx6UHIbgZHDfn7riHRCa0H9XSxoO7HK+V6q1s+JV7XW4oZqfS07vjIBl+AxF
3/L2iCtm2uiQNEq99dp9t+1rFq3qQX5Lz0AijYnkz2ZjLkCarOS4CCeIhTFYUHYM
n1+pqG+vydy0JkiyGr/X8NVGNfvaFylVPCU/nalLpevE4bupQCCa7S6ZO67rv7nB
ndTiGHpKLpEwfIAePq4MiBrc9aVYS1JuOvEYw8Wht8HULe6pfnAFjImrb1m1PQPh
H7tJzBhAGmJacAxUkfpJPvNyhIgWlsQIQsQ0hw6bNXvt9JsGfTiZFXU1va5Lp6qR
Ev1snWLxv10BPR7IgBaHTox11zGtpteHMFal2zMjmcfwnDspxFFDRvFKwI5EIh90
wMqgIvimvB1Zx3VbFmLtZ673dCq52sbkCSKd4Nr9tn4yierQuvp9eUjueIr9nAnK
M1xeiyeH8cpihOhCPRszatVrwPqPtne3tWd7JYxmkyYyBSsFhWaEdf2hKjxcRurw
l4EUNDPV05VR7kQDpMBiggA0J1INjrsiCxUl9VMWCDHoSCPVk+To0XvgXNo49lTO
0X8MtZtMCFR89+MZoOtNM4mhrNS177ur44Gmv6qMDmSUU6KskurM3KwqH7Mt4PPO
0ASVtJxeOPmDPT3Kn2p2QEd0iS//rktZGhnhbkEjSmbK3CoetcjsqpqUHrHD3MJT
c6290/TMKMHypFWXlScuniYI+3hHxErfMF4Sl4KpMO/S5zujqH+6PILU34gD9JD9
wG11o2N5flxOrZp/jSEh73xf1jqCbDud+tGjVbkUhKuMAYMECgQX3fK8V7l7Tj/2
fVNB/AQJzBFI9Axo8jrFF6GjmcyWj/NVShC5erCXwgvYhbxKc0Z2NpTDYKgvrjrd
BPKOVD7P9cu4NG4sw8qOKAbE6mT9TWCC4Vn+Gtzw6lg+g2+z0Ayz4f5qr6qSBhTQ
P/dNczEC0AP9cbrciUho/hy4eBv0xAtFbwDWmSOsOK019pVTLp/CPMa7/73n5Ece
eLq55If4TOD8WBKvXpObFzNBAzSb/T72YNTDSsnYh8mymnTeEtms82ysQuV/JxIX
Ubnb/cAjtXLzdhAX6ZhTPpTwjtPOukw1vwcWgUQZHmAEaEOb/WlWWzcTPAaJNQy4
vIEDzd3Ieih14Gzm/3GftxSpM+MylDoCYn4MTd5Nrj/OhbbS3G7x0CpZ1DCpZZ1i
T9Zf0V71Zbh12pM1aVo0dtQYcZCcF+bvqQuEZrUqhD1meej/TTmnVlHItrhigEkW
BWoflXFZ+pJ9fO402npvWvjCa+iNTdpCujrrYyn5ieIW3Rk+81tVtwi1fdsXQqxH
bfgWrBrfXbQdwTfALPigdBrXCTi8k4vsJmtX690LnfTGC4XV31RUwEIu/8nVNgtC
HO+4KbWDgZr3OFcl2GDIz3A5elEfDvTgMl+EtEr/Ifp1j0ifCWIFy1caZ5Xcpk+0
WieWBOhdnb4WgCcs1qDX9Gs26VafsA90yGfJm7/wM4Tc6tJi/9/xW1FaH9E2ZLJv
dvYomrABVw6EJzKLrTlv3TINxbhA5+TTPP7DNgwid19spDwwohmbRSywmho0PF0I
zrMTnHHcNrH9Kh7dF/6CgUz0rH7MO/hhVWVgHOmiZEdrW1Pt8NMeiiizI4MrpJ21
Eayl72EhBN5slP3iE0Sm7Cb4EBemuQZ9mMA19cArvrR8t9AxemQSE4dpkLFCShm2
XIy4ZBpVDTvQMrALZTbhiMHqhEkKr5BAH78WtxBphEsTxmp1XxK8dseLWLko1T4i
/Y+BlUavd+h1Ljx4wpNo8S0iOhr9joSzd2/EdFEzcpDn/8gzClELjJhZsi+KqaTc
HSWxWHOLgDD6tHHr8hJr4G0ATE8xzXXIZ0L/t1yTyDQ2kW9D2+lGk5gBs6SgjX62
NLukHuo24+NXWRVRsFhSW/NgoNicTSnRCksQ4ZdBWozVMZnnTCMMpIk8ZCb22R6M
sfduWeZw6d7BOB3nr7/ofjtarAx5gCYFEIqwhRkxf0cMNC/fLRJ/BFcoCAs/u6yu
e6QiJ59sDMxmUAehfJn1kqLjW5z4xwu5ZhRqCXmyLGd9dk2fSNU285+mKk3zXnb0
EGd87N/FCfa1OV/N5D9qnroOd1/CSUc9TJzamIQT0QsJEhwur5JADYq8YoK/xDhk
v8VhUVfxr4W/tb2LsMOWqhbp7VpL53HkliXo+6v424VyYHFVjtOi3q2DEU6tZEgm
AHtzibHUxeh8hEsK8PwDO62O19HNVSKvzURf6BFeIeNPXfezuc2gfLlEv8GF/rcU
Sdej3uzOX4tvnLo28/L4rP29Qv91U4YeS2fn3JbXOEL+6D5G9UwW2kJKDZNellG3
VocjEL0nZlzs6ThEkPcNRdRGLgXwnyCL7Frl0YpURisTsMhBsyaFeaBBCFmJs7v2
oiciQ52sLkpSjZQlNpQwWstXsB01AHMGtHnFCDmnFsbWVM6/KyGIkxq4IfYEJB2m
mGvgN/rpem2DSbLFim4A4ApyJINCZPYVh8aYqBxNPC+/MAVhq3B9Ohf+aXLcarkN
5MS/L+svzEuFUY+MOA7IFJe+BGuhepA5njqYA9XzlRxKAtDN30KdzCIe0jGZr0da
ba0HL1mNVkU8kFNcLUmsXFOIs7Xypi+68wc2Ehhe2w7fgBhwEPTCXdCqSUad7upP
xkX5/XtLVt4d618koxMXs37K3n7nXRtVQ4LaX8ZFObz5ND17aZkM9aD5+38w6aHA
NpE8o1ZDsaJ4CeimFg/U/RtUFtItAH1Ap3ePYVIKgSaLLJzOmwZMj/VC/3fWid1s
dj7BKbyKESj3x1oGUef7R8+pTQTlDEFLJuHLlZSwEO+qqIKXI0lynlUU88bOUc/b
tSk0WPGS+5H4bBHNMIWkO14gE4lDw2PrSoO/4a8/MViYHlXvm78tCqB9G97WqyGb
PPCeyQw9mr4jhtiMt0VZu9TBwFPEmACRK+Yo/A7CPP0jjxOhTDEim08SO/VXKJPx
hHZ/QgM9CC1/9VQOFKIAOzl8kBjzYVNjKVO19do79dJj7aB4CU4ycTlAUrjoamLi
i1ywKk9l6gNX85LwNruxOM0z9NgF0zDAHLHkfEvdvYyotLQTCOaJ20h6ub6f7UtZ
PLPcl/yOWrNthy6X2xDrTT0nclc+S+Kn1rnMjxghCqgGZARuDpUhO9hkxhJbOHsP
+CBGMkgwCvAhQWoK/gZFOm1UKJG+C69uvG/AUUssPqva0IqxFQuQ0NlpGeL+yjhv
sKCWDG1VaYGVjhGIwJlVPPYDBjvIOwB4FyqEHR2kS7RqhpWpUCTxfGNkJ03sU2oz
I4DMBCvbYksidTLiHSfCVKbE72qAu9qXpvlC+z9JdYQju2EQ293bNvm8Bvte12wF
8snFhpyxqVdowq2XYWtNHoxL5qBXXlZBqkqEum6pKuYlXIs3MGc5HZiQDcaP4aQU
z6EPbbBe+R/BStXCi5M6FSi1OglYulwTTrenlzByDTDRf4hP/WiZFjCJR6gv06sw
UqLH4Jqs8U7lCj3OxsnpDoYJM2w3Jg9WZ+QPMzGz3D+iKBay5k0+47Yd93VEc551
buUHBiXpCTDpQCEvCbX5VRI/A8+YOPR1TdHaaC/kD73sYgm90Vh8aeeZSlfzhgAz
Dg9msTn+H6zmiJYwrcSsPwHAX2nEIRDcdo8T8YKqQlbqlzkEEfJlHFmC+5l1NwLS
v5zZkGgl/8lvqttvHAR1jPvFFNT2fSTkXXF/AGxdkUuIm00rFdIZfOmAQECvRUDW
xOsPiRVI0fWvf6/EIfjYoSdYg7q9gvCZ2SfEZwUQcj1yHTYUbAt/7y01qU4/RjXG
4AneX5zweCEpI8eGLQ+HkIN9SAOi06cru3o1F2oyYjCXUViw9thFDdtf75RxDuZy
2/kLJAPRQL0cs6eSJG5sTxYdc9axE3WBclNEF/Ri5elfMTj7mSh1jne+WC1lYM+P
dDA+ZtDsrW740PYNya0APt1A4pJ+LTzMoEG3GaGa+s3L/Xl3gGfCYcLh7n+AZCky
+Vp+Uf5JGRrOoJ70q8YbiQJA0PJhVZV6DZifPXYmyJzMZglJf7CICaFYKqVMA+u3
bL891J6RpAKK4g4ugRo/SmJpNnxs+vD2r7WGO8p9GnmW+Ue7vD/pqfGiKsy6Ik6T
59XXiGBxWRyTKnf/JQ/Y5UJLc8yU8MN6Rufdo10a6WkOm6FP6KHHzrGkbhmRascD
qtcKZVVXqok24UXS6hl8ClJYy3cZ0ciLhcd/t4jm0cg2drPZ4y10TfLPwd3ZqMD5
LqKoxhcv2BH9Jym9EDCCK2zfYiTMPo8/fH2Nt5LAdhsiIbzN7nqglU8BO+7t2yLm
kE5YfT3EMwX1xaTgrDZ9XGJBVePBH+iBayoNUxliKeOO0Pyrk/6b31M1O3zCOLZA
S5ibyfVN+f7bThHHM153wXbbZjKicZHeNSTR8btRDz3P9vEUMrV+aaYwTsvlIWop
aGpjTJhrKC46d+NHFl3tehxlfgHjTlVNMEaesoIdkngBF9Dwlav9pj+gJZQgn5Fg
c9siwgeb2C8hZAjfMuzt6PHdbseo+xm8wWnahPpzyBl2SidreBaKovjtUsiN78sN
aMKUFYDaMgHUbut2WYUXxgPSHzkPp3UMFhujvEddecEsSthc3y8cAua7hua9Nr6/
iQBxQaSL7ZQmhP595htYRlFE9mcHPdE6ng+3SEuNQVjq71BWnsjdQaaZGF6b1an0
CXFTFoDPfB07jo4YhUtSNrPTHoBi37LtNSTn3lv2tUr/hf++tTBx/o+IC8+Bac51
ZJcS2ADSX6wsOUZPxtzA5ni7j9OCsdLEReKeyLf424Z90SCKmN5ruw7nkso9nnYj
nuHMyEWVttZ98qSsPJR9HglksXLnX8Y0QUpHlCuZggsNlyxsf5w7m2Ar8Je/z844
xD7J2ugRF32Jo7ac7VRp6HCamxZBqTKWVLLuVfOwQo20G8IYU8cotPeneGO9EvI1
p2zLRVFlGI8+sTQLiZF4lvUvYtYmPhAR2G73O0DXMso+Xs9AbB4qpZlD2zDsYOTk
R9KfRCChbih3J3wXqU1oHQT+R36LdEng2gIhGlxGrQq1jNLgLeu9Z9320v7sWaDd
BTQembIeSylxfIebQzNcuvl20uF/AFRtbrEdLEG48Y0GeVj8tD47z3+M/jameKZ9
eWUe7mJcWxEt5IwkFXBfijmXqnO3mQrcJYsRm4rRKyK8Om9b14WY5oHNsJ6ZoY+z
DGalhuNIrKkCMNFWzUNGu41eXBJr2hPfBB/FA6i657z8X2k6vX87hvmjBeIt3d7o
7JTR8wI10YatzIHCPbvuOOup0xeZRj0MsTvZ4/K0E3GVmSpylqcAaW2ELEHb7Udf
AYFjbtjmrxW2k9lfXl8o+gDmTmMWNtJaj65FV1pXgt4XxUWEHgsnKBFqtwtdIxEg
Sca9ZXScgPMsEayzemHNsxBZRKs0qg9CsXu60mi38Gd7El6mxP9C55/sfDx9QzaP
PCNf5NU+ydRoDDWFWTl4G6Z03WBbpiTf+DsE5ZMbjB+K5FppJgfKL/BSHAaldyrR
Ya37o4lsv7Oyj3leIvuV6GXd5Qw657oPIwCnZUAyRB86w60WoP5YVLk9WmB0mt2+
kB5exIGgRS2DrBYd6vAwOOhH65Kcg4zUtAeJ4/5fWPUEyL8vTTur3Ip8KDF1av/1
uaLbiN3D1mdevmMI6Smst6GI0/IQnMmE0/BopmzjDBOAq2wol1reMWgk8OVehN3P
Pr7kih9hpMOul9NfN//PJaqTuvW4eekLcRLYyrgEr+nkqmo3yHZjzSczI/ZNG0oR
f8YE5/vUVH77YvNWLcSQYhJ41+GNlVnIMF3RQk+cdNov7q/BG4Jpcdh4QR+OVb36
Nnp03vsc0tp59JVc4p+bQK9ar6Ztmft1eSA0XVgt5KhHzcoprWdwm/R9YvZXe0Kd
O/dyBtvz7utbBfBtBvwVhkX9jKpATcJyuU3dMz7xy6rD7Ul6Jcykr2KKuo7kqcGK
WQWJPQvxIw3PDf9XWDgaW+7HHtPWuI/XBRj2ESJkCr/g65qDdmXmbBDzjEBI/SgR
LQN6AeMqZ1LDfCkp/khgEcL92SCbwuqBSziVTzE8pMC5betYYIAwqMpG7GBlnsku
MDCn2DyIpR9AXkw+WnD9gIGiO3Bba8nr8VVnWqlL0dSOzcdMFvtARx2CQq4bVRIc
CKVihHdVIs63XsAPOel/fcRwmOUOKFAuji2YCnho+3JOKtsvMUiT8dpgLT38QTA3
FGmsKQ7wQSnSjf1u5hjqn0zbu9ncMrKIYCxAdn0CnB2rvsLpCqzvbJNBJn9EcK8a
EfLgVrPQp/+eMPJsPC3AWgVKun14G3LOkGvUI2KxLjC6ZGUjkXLt8LrPSpxJQeA5
TrXKaPhm2mjrZPggnxhrwfw9najVfCCGIff6K0ayfw0=
`protect END_PROTECTED
