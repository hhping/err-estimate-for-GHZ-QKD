`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vhyf/mg0w2oRWUR9A+Qo/O6W7o4BaPkopscdgpXzssDdDVbAZ0HPDhwPj/Z5jIjP
SZSgsokG7YhZ5U5gVWWKRLfKGzxRLvFJCAxvIOIRbBCTVFTMjydCNn7Zz0sjmois
xQtgWCjqainyLh0ARqJQW5SMMzDU4O6zbH8kz+i3fuT/QAT27KR/J2+sNDjK2ACk
pEZgNyq+obeEfghdBXx5LKazRX7gVXWCRIq4jUqGIY7r6Xt65Bla2V3x01maNW0C
qDDRV3xy6x3Wq5DBtWYcG5IlYiOBuAL3SkV2Tl3GiPshB9m+M1hw76+2oL3NARjS
4VLcls1vPBxczGduwAchH5i/XXYkbOfgLc7UQpODwbNeG1EPo0GvP+lVsRFoM57B
RQqam4fp+4f/Hxg32xF4PofU9YMGxnpej1kS1HvJ53uMEtTmI1IGWlhH+ykHUBl9
/aQqn/3pzZOVhJBVsA+PF8eBNxJ8zqgHmcvsAzv4AIPYaP0qZJLjrk880KwvyFTs
QCycE8T/DnGj/AB15fUV5kqWIWlu0MoJr+7gQF/HXvMdYj/l97N/6o9Ls7m4nW7Y
m2BwSfwHfqVGVLx4mWoETrB7kyxA1/KEkXBRrW7mLvFBgweSXVN4/1HKYD7tlB6O
qyHahYqNrdCzXIjgbwvX94nCRa/MXrINLB9l73f1JQfPB/YDuEei0anm0KzLAb52
oVMeqYyrWLJS2+L71Ebo/WbquEsmmWtey+Dzvdc+hE7vlqL5XOn1/lTa28hXlxug
pLlUOMYF3GbVfuhHSG7FXcC7ESpERjl7gdhc/uXzgL0yL1R6Vygw4E4yYwIiyWHg
gOLxxuTM5xYiVBitsVEBRV432FCtlvTtEWcON5/du61VTRXi6Gt9Bs5EPLewounj
sWTFoPGfWC5zy2IIcrpPYK/8V31bPZ+JKFVoDlmY5Tg1NBhRTOX5Z9Uh+oOL//bk
IH9o3Ov01P3T0h9W1h2XyH6fGOPb9xma8RKSjxWss9Po2mcZx32MNDMfbycVBvaL
/XSA01SrK5lc4iL+RFTq5HjmR0qVPso1jzLbOQUMmPXohLCEwnvIESt3cux+Kfrv
u22mTBdxocJJRztQAtT4WlXCNtn4O7IKDm9vt0Cav+gX+uEqzS+0OZLA73WqXgHM
qKLtxAmEMgADVjOL+sbVdBWzkjpxKV9Wf1pmGuh9gNE666LwrrdJ5tSNL7kDsZuy
cD7rUE9ZpftvsfpC3Se3vF71es7Xqku3M4NcC01B/iKMprhg1DaIiV84h4k3QDJJ
cBuM7nBAVVuGq9Cx9R78owvZEMiDS3jcsPaLup0b+x5zY7ZFtLQjFLWOLEohbNG3
3cihQe2fOdBc8qomU5MyDjp/QLdQcL0FvzD164EJjZ8kbUtcF/UDAJRCUO2scZ+B
R647M6I/G598itYf3N5DHWaOdvlRFyi/acZUOn56oIpFrMRfRqDXUADR3FQdyWj+
ObJOzGoOEJPKhZE4e9SAwLfLyuxgU6VIeun0Jvbe6QO4W0+Xt+eSUcXK4hiu5rEZ
U0bUHSPXfVO8XMI/W+Y8CuIaf5umF5547HXXZ93NKzqDBd9dLISEy8bx9oCedR1h
BBf+ShPQCElQ/CvfZJkqTtxkc5wWDFh3B00wZnj2iBSVEwdRehjKZqiTA3r1DbTn
Ixhv0CdpRRblJHdixyKkNLjIrSF7zyJTmv1ZIiB5WbmIUKt160hcXAd4pipSNP2W
/Bro+kcAPddVFH6An/MPd4FKMgqwWjV1RxX/UhsBWqa9w08jkNM6U95+wiqlbIZG
Y8JuyfQhj/GgtHRgIPzioa/avKA1pcP6wrZomKgxxIF+sBfY079zq6vdL49tvwW6
ix7hgQ+PkBq/7y4cC+yQq6vF/AOzNY13/f0/7R8mClihpMM6p/F1EgwDS/JbS3bL
5APv7VNw3cJ1dCiQtFSywtaHwIupAGnHVgA3HRyZGzQmVfXBN0RP3zmhbI3zBrU+
klrmI1lLi0JHBTFN42Arwx/3Ozi4ektDGCty4jegJwCDC9wgcJlQGy0xrXmMUVlj
Aa7cKGZvZ9ThQcSFRsO3IsQSP7xwzRzOrPImmjYwbnbqix/hrW01QWOZ82iG0aAY
zD8JaUQuLjHX0RFLLxNDJ/9uV1dLp6fSPyP2yEjK2UOc7f7NPabfkzVX4kHcUjgz
`protect END_PROTECTED
