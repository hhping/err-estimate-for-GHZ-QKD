`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+RPsmbpTSy7CeODTO3zmG1UzCHaLe6J8g2xOmugnMQ/kZTNQzvQuPF/gaGwK7gIk
TsAYrxFcufRxGli4TB2R34eAMrKi6dny8AXEt9UWgNiotI8mspNgwum8xEXmW+Wb
PEOoJTzoVcYofLoQSnO2Ka3IVU9muDVjh4pcycxuZnx5lO7OZKGCDMhNJNt+odlV
8vDX6OPNsjFOTNrJiVmX1QspyPF5Gr3Gdc47DKy1r7i8PnQB7DhgTy719O6Im8v8
xaep5e+AvXzGDnlOotWsZDJj3742dVDXDsNtHY3hqoo7cy4q//hmrLg50sUefc0U
bwfc/lZh3fCreKaYKeTYwrCOgoYbrX5jPY+QEgeLIMFXcR3eHHBduKifIMyv/UF/
p4BHYsbBwEk71ahSmJH3/RVe+MarjXlvAISF26YSXHwPgJQlAvIi6gLdmBVjUqFU
4jeKCWh2D2agJiqOEbti+HQVWohxfjq1aCJ0NCmWVgkjUMI9Lt7nUNx0G9azFRc/
FB6oHuby13J5ICHsO99FMYvLyuzMaqkoUZxLSkx8SwlUeR8SWtnV7COxWQ3jz7aw
6wf/i8Xecx8SK93gUAX4Nh2eVcRBKuFmnWMqZZJuW/yNFNvEdS9JsEuNzLax6MQF
YdcX/qvlqR3h7xicuEJi0JD4aC1zw4ykoweJfXfi+NBPfEROtxhsneMFBwf50aFS
pS2HzKW+2SGMpBKsZd+nwS2y30gKoBOweNsGSv2hAoMfjbMT8dBEYSiWBLVcs9A1
yVZSKuBHZU4DFOjqNPJeiSPxdpWlBKguQBSpQeXKWgBodNW8dt4MFDh0OIW5Wl0w
NA/qn6hdr4MC9sL1blgC7IswB+1Y0bPP1M15bMqfYGxmaqbCWaRGPwyOdkfEtsUK
mVrXn54R5Pv/g+wxOVtTur019/E0Dbt+HQgbKdMefSnKE0Yi4rbKDGQKIDDb2MH5
7FZrzQ8+atxpZ9LAfKm9CmSN0o5TuUnXhKhoyBq2EmMUb9NOrQrp5ZisQnmldYxX
U+kPknOu7J06y2OqxT382bej3OF1t1zcGO7G6IRno3MnYL7XRD2Vmrae5Iz43GvJ
9muDmT0G7xV+Z7FglvobC09SqYOnm9h3BIO5nofE95OD4PV4/8hAE0fLT7xmZIUV
vBS6yAaRry9eP+RqUTKa1xRZ/r1aiIoxAAwbTep2tXe8wKgB6R4o4ssLg9WiPbxM
ek2e1PGRJEYdiv50UOtVjla/cNOFoDx/TNWVVo83gLCgvmC2wed2pTyDcaYM56dL
0ozGJ2Ksa1Kvcljp+dM3NVM7T2Rsqvt5RvQtB9eyI3j6DDmTPWn2JIXjqqDw/sZJ
kTQA9udHvv4oSNbFOyVMRI+6UYUo4WcbKLzhi7KisAGF+jnLhqWE3G0ImUoF+W8G
6a8vN59wkSnIbWWX/TxoZfbX7NfSOXaaJY+Fo7hEqMASxnaD7FuNCvE/QlQD7U+g
4EGRQoyM+i9XJxmRAv4yo1wZ3FmOxi6dHOgblL0KYeQ=
`protect END_PROTECTED
