`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fna+UuDs2ib+ftL7/+eqAa846fy0P5hWMUwZjcT2sH+MWpMq362QkzB/FZWuqDa8
FPEKx9JI8hQ9/2wNQiqLWC6VYtZMNLNIaAfGIJHNGubLbK0CpeRtA5Wrol2zA1+a
sMht0SbVyLcpQ9DGJ1s4TlbF+Et61sUR8vMUwe1jJZqKCEHa6atjYyd0bAKOMgmy
ieOv6aZrSGrUXBmQewdejXbeEGLkuRKf43g7FE1jnV2SbyA8ckmsFiL5jhfVOLTz
e+M0VINGbExH/JYRwTAS/e9VRjJ+u+0AdRfk+wHmWK9L0Nqe5W1cskNptgxbzo3Z
feBzdK6aoQjLwFpjY3tAOBCd0pMx4xXlwNwwtk6x1B1NB9YLMyQc2VJkJKwoxJRL
xE//M3s9ijFBxkNWyNe+xIAOW6HXFNPnrDQnqCg9265WQ+mqJ0qpYwLG6wDkI4sW
HdORJ8vDDksb5Zip6QURGw==
`protect END_PROTECTED
