`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/tb30KxvZXMz5zR47SRmt1aIK2Eq3Txh9/A7l6E08B66EyTHsReHAdaU20V0qkv
e2JeSKh+vn/DbYlS6AZ6gZFNOy513QRG6zQwYB9VQ+fnJHtud0ySZ6i52rEIUpZ+
mX4zT1KaqZHhpCRkcbtTTwezvgfEdSWgodl15eY1cHxZemXiKCPTHpYFxAL8j08K
RXHUWCJ990oC3mb+WHxLJl4fuKYeIyRKrw5V/iuAKbYECc6d3GEwTUKXA9m459Xt
jo/Tr7QQvk8ldN6cwxvYw+hrdzeyG/V88ns6wc8Xn+iI/nw/5KV/ZkHHs/v2Y57f
BiNGdNJOJdDQm9mVbQlkp5TTbzpyp6Ch2lnoBY5AdRbt5U6/bbHAEVtHvVLM+iMS
r0mVb62l6itGsHidVLi/bY5ikAQAJH1CQ6j0U5Rsqnr8QIC+BoNMJ2hqftGGFssO
`protect END_PROTECTED
