`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adRTF5zQfw/eCVdWNg5yHFPdZAgRT39sUPVuP5rv7qdZOKmJs+l/NOv4MQ0YilXa
dioZDXg5+ZnjDmJ8fHV82qfi3x3NuF4e2iCNr888m6kxnvbK+Dhyx1EfXCEfsYoo
cQHx4tKOgzeFFUfpFkvo+dq8rz7JdTtBmvl4NYhgtxygd4MggvN4R5KHZn5sFnXo
KS5dqA6AiLKcPY9ztF7ATDAuteOHT5ljamZ4L8eDPJWbiTvczzEt3rt2JWkQO9wt
/adNYksUG7RS0HK5VUY8JYr3cAJz5Dp/u7EkI9Mkm15Yeq32wVagvBr34qL9MfRn
eN8zqMPz14gTXCMsAPmKpvL3E5R5rCb3cPorpLmiDSu5IHuop8jUIdeX4UUWZpPr
Yw03eI7ORcSq3MINXKwltOwEQFNcCaKHD9IFgQhMpYOD8LOwW3INH+lhNCdJ54jE
XdmUEbQ0kd55WkNzOpoKGihfqutpsJ+I84Y5VXtbXM2o5UgyfDdFZG5VLoKXQwan
`protect END_PROTECTED
