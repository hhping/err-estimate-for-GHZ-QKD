`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dy4Gqm2anqvCy6sHKXnJ7t8V9SRDJx2zakJ+PjZrM/sgfvOpQnIMiqF3A+NmnA1r
rGzuwnlf/IrtOIjQWjA4Ps2LiiOA7BOkeYMzcLic+5UbWXRZjtiJO/eB9Ie49mRE
uzLvC00YcEczwUGeYm/rXDFe4IJ1iJ/dqFUiYWnkx//jQ3TnAp/X2iRQryB7yJke
T5SBH7jD9teKzTNfIXnxxYB7HHqdd98TNAoLq5RsspPN+DeXfa2hcdCuIjvuzLiF
y5wdfb+4sj5Jz7uMkQ9V4vXo3yGHTboUXKnhXGPZt3BXxui8HJkDQJAt5VMo53lv
kB1MMFS/4t1qz0+XnZuBHL5ERjBbiPzEfBsLocWB17f6obveCuKQrYlIHtP8S7W3
We9OCKAz14RF/SLZG5nZxdV7S+8LFHfhTUBoZ5WGVg9BBKHMXxzoRmJcTiVxCBg1
2Nz6BUxekCXJ89gdjRLoITSrRpCLlopDhK6hGl2iL5+uZ/WEZ3uzbezGEtiSypJr
/DiB+LpxvR9iEPEunClnVY5mxKYEItDfwTJqzgF3y8rGE+vsL0v3ugcWLGXDBDJi
yob6UGo14Lf0GcreDsyLMjgZZLIM49YbtvUIk6+4Ua5GMVz+1/epEaWH+ct1DUi2
KT30FrH4l0VTpgEoAIMTtpVyvCHsB/nnQcyODWEKamDX+34fUciuurBS9ybJbwD/
P3CcpTAWLhF0ux3WDEqfb9Xh7+Kdxq0IJOwwfS5z8P3OI+ALuqW02VsbOn74kPUN
I3lPthyowUfrRdDERwJ+egnNsey5iJ+MlqZDinxRIY4A090hHWamfXCVRI++R0GP
VAI6eLmHQ6fAlXkLU5VK9v6kvzW2ZJOhSs8lxLIiuq+VDj0+MlyfL8/2hgoKGu77
m50gbA23LLXmBmgiXWz2XHQX0pHwEUAPXFXLS444iiHzRDXHsHYQRhuPG46JynvK
XdoZuYBn0wWKTLJPIs5gYTxe+xV3Ymeu0/Hgp39vp10=
`protect END_PROTECTED
