`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fx/LTqXfjnKke3oA+TVv0F7qOGoRMSm/QzBD9YWh47u4uGttw7jehsM2rJX1tlF1
pz3z+YHpUZBaZbllhURyTlC9WKYLnmA0/sQs6A/gaxGg0zCROilS0tiYxu7GMGpy
uLmiKBUOVv5JlTZur16TlBxjR9UrAb4KFe/abHJtFCQkuISC3s1UvuClQY8t/44n
BpIEruMtDWxqdxMNZGhn8gSODcTUtmvzd3Nzy4L/8LQq3k6XOr3541RfLTWPeTg9
sReJ8w6PxzrAYRppDI4mvMuBtW8ZEh16XSzC6C8MABPWd2XJzG4hI9ATEV5Bj9YR
9jlT1XpzSgQw8PN4gW2U3p4DFNXdZY7CVSVboqq+G/Ydq9x462l4aUAkOoiwjxt7
7bRXrA76KvkMC0VTA6v2sYkrDmEFAcu2tPSWvTLJTh4t8TV5qOjAr6oOi6B4VqGI
bRg5i0EjL1gk5kdxre0WRM5MwLced/0NCqJ62ivT3CSHrYirfNEOne3IN0Df0eog
lkowdnA8Pp0pXUlm190zKnNHMhdHeN5mwiBbQsoQ3xgwF1G1cj4Hv8pJYZ2Mj7OZ
En4PoZ5+ktb9HjEqTYkRkPkUbJ3bRnXfbN9S1jI78vyPWuU7j3o+Ij/cLXykuNze
6+p9j8csUKMFXJGpraucnZCfe3ivLQeK++hVTFllmwLlRzb1UZkk9rlU2wRrXC9r
ipI/ttKioMwULuKrPi6aLRG4ZZevEa58/Q2atCekVr1UExCWV/7hpE0/8feRc1XA
85zH4YvAnie8bzGEXmiQqybwETqH1crti+g5gtpEoT+mBlqQZqrWs4HZrC3QhBJz
2N3THWNnjqLUcfYVGb5aJxUNubb6uG77X75ulT4WRo6W+XdmOv7N+L60kv+Uml0A
VKZc0uEWbNYYt9uAapijCmkW1SdfdSqGxKKYzgMKnGdKUp3eSlB1gmmAxXzxQhR4
n2X0aQODXg5fwCF4M5SqsPZ/wnKfTkUr9NXttujDDTfj9EdOocTLykkFMAYgFwZ+
WpgIc7/65XKgoG+ktXlDLS3ijrovqFGfREH9zTAtKzix484aN6RmgAWthMBqy1Uy
aEtnZF3SI8W61p/LwxTECiGC/fwYjwt6toUug7hip3fb7gpIyFWRVRdmZ9n79u4E
1FhDHr3lIAS3SURReCHhZE8p6MrPiorxtFDgkOLwisF1Yc6/8TykO+YlRnvrxsI3
z6qkaBmYzbpZf4/IyFnhxD2+lR8T4z/awWpNaNDhQ+O82lS9NARv0pfnNNf2aG5l
rFrCYupOMldFQlPsE6jYyWYJvukjF2sFlKyDVkUZbV86LjwPllb8Q5yXLkizfLRn
Z1Jl0BzvkAxcf7fw63UihlVWki57vMwblI0jVjT/btdUPooYchAWsyi+D9WRC43a
PUrGamgG7FoVxb+Kr4YRaZak0rRoEw2FEAzogxMAAfqx8nCtFXEfMYaP2ozs25Hm
AhNvpoamYIQzghGiVMTKbIicDeEuppPrPUYtzLL6jnhqB6nwwjK9BFtc33HTekpw
vY2R0lZy80/W/2vqFPO1Hoq7Nb+skxyfMuSS9JiyoXg=
`protect END_PROTECTED
