`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c96BuzI3fKnzLysjb9T3btfYk8o8AKb/xTR+5gvH7ytnw6jIm3nrhbQHbdCIttPp
u+eXAXHuvWb8g+9mjQPWLCtGwKPbn13wWwGwjZO1/GOGqDOUCF/RS2ObLqQQPB9H
FxCE1y1Yfv3c9w+zCwAfp3CEcVus/8/RFrrr6S8ecy1mw69mfMrD/EqLkcLVgpyp
Gn12kiaO0FDnaow8LLHQfxBTWtrBsizxqctwGj6iH/gwMYUI8TvVAhOAb9KR6Q1u
zjOZYzxIGepp/5PScAiBodHnoiXJrhiESET0GCow2FO0uE22Hk1E+m7Q+v/QljCD
A/p2uCAcoO90BJ1i6gjHsTZdNyjx20S3Nhk8RuMni47TgTmMbhGKDpP4Lti91clR
gtMU+c7TZGIucydUB1/sXQe2cbTzH1kswCqLApcLQivisS8+UgZJizmm9lBE+E97
tp4O4M44/XMqZ37e9g51RNA6Ej7iMyu83nHhHArT8U8MHdVIfCmZQa2N0/V84G9Z
`protect END_PROTECTED
