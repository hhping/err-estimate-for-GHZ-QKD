`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZJsT9rNSpEAsDlRYHKzY2siUPketNZX9i4Q5HxNdmQy+AyTE0YkQSmpzpb8PA5U
J5Ndk+huJPk5ZTkA5V4S95wAp9oGdtvGsYJAhjYNJRTEXZ9zQXuhHoiyRjByKyy1
wHZmE6mntLuWcsCLze2jgU89htL7mi5GFr7huXLnGs4sLDfxI5d3ODa59uFtHVD9
xUo4WkCqPnJ3fIG03UOyH//PUjBDzEBPUvm7lzAhQuoAnMjoSFltV+4z1kWoE18X
QXTiC+HTa5e/sLIcRDWgDfH8qoOb2XbcHNKqQvfr0GNn3Jhpmcik+3O1nMgz8y4N
fwPy3pv3MH3fJzTDmyIQ26G2u395nPY+M8n8erPhG2vxR4o32M3Yq6OsANqUDi7j
zmCtJt5bTrMIKY0vHnI18Dix0rUAjKaoryMfkieOp4t/8rFC0qjLh+fYd47fjT9h
mQJAvV4aZ7WTU8YeuCyr1scEl7VKC5GqY1EzrqD5ZF9CAO8qBx5EEw0kdtd88+rg
+opKQc/xR0sb7RGQ/495jWh20rm3QzcQTTg7HsuzmUaekA/jLHC9ODyXUYYnYGsK
sxlDSH6W2pRE5aihSx/ti/YdkUBtHqJxebxFQGFvAH2dRuTMmOr2W+uGx9+mwA30
L6q/dTV4WEhswtlrbCbYVSHEYKs/1O7oi0yjjUzgk5HpHO7K9lOn08D+3b+n4IHN
GSsxzWFbFIMOmVknOIZ1ApI4kH1MuMLFyKXjwBF1E/U=
`protect END_PROTECTED
