`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WL6wuJmzU8VUSA/0of/zMj5gwxCgsx5eF3nmdvR2DyxHkfHHyWJ5A9l9011FB1zw
2gVaTpHYRi/ixvFH56pfH9uBCl6j158cpMBjrD7SnKmpjHTvlVgYLACcIc/4r56M
FaEFSmiN06JHCycfVcdZkQIw9/6Oxniy/5aL5PqRz9iWkwMlda8+YoP8BZX3LhPt
4MuK0jiYDU/6hD0NyexDOuITH5fqrjTb+yyAGy4CxvaVh/0j/7EbVdGTz+vtSJV3
uVpAf35VnUtysE8V3SDhzHcdE0IRCVYLUzQ1EMVrkp60pBA/Zf/Ej8kcHX89Im7V
zXb7ONMH1/IpyrlDGoDo7kMtU/hmpZA9AVaLCJCfdimHb6WzuPvaROQg289KvbWT
2RfZSPkS6k5RHRCnMDoyVxBqMYddxv6QTx/txlDrJmml2acnA7jSPWFnrvn4v3a9
07bNoEd9HMeiaEdIr6h83MazjaYHCfRwpI1IlvUehMxuf0AYggeIY4Zp8B1tMpTN
7quhjfuqH8Z+8zKM5oMp2982pCY1neu7k2TdkFvUw5P+gy3xNYPzoy3Jg59ostQK
3Hc48F843h8nq5x1JGWiOAe/mzmeKPu7IUMpTwwtvS4P1+YYV6JgOrzxyugIzs5O
Xepp6dwXT4qV3oiB9tFw3q+TxipzKgGeye+0v6JJsNc5ILyuBVca45WAqULgbrAc
Qqg6+0OLHzGMU8q4z+Rl3OjfS9GiuQMDaqhQhTZUiZJjF2gpOMJ5lGlOIZkx2IWG
WGnTQxoYSG69uwaFsHAwoGfQNX5ty3A3s9ogFkLkKvEJz2fr9yILFeldVz30wg6s
hhxcGXz7JtqWf+pIhAe2GqUr9TLrLBvuQ4GcYS0/nOYBqJIqKuLzZEydrTheMNmZ
tbBjHM2kDHhHqsQ6txGi0H1GHBRZQ28izG7wI5fHMcso2e5tfOkdfrYNgHeYq4HN
ugNZjfunkjVIg/1QswTCHGBg/B8ls66UbNQXQH5AVSMgjEJw9OSBHr7/tXeoj+3u
8rAbbAjt1q/i312+L5H7DoPd/f3B+mK3/RXXCIp5RkcVjpAlZbqN/K6uFf/SqV3o
H6suVJ3BFhxuFElrdLuSohhl9VM+ss6Q45VzXoCrByXRvUjVt/NFm45R2TUT95th
44HA6ThvXzzMj6cttQGysKy2kVdmdSeFB6agyNudCxbQFZXoIi3xE4k6DHkggqAH
qn7Vuit+/NVjFP+gLFZntFikwdNb0oYhdLQJFSxBUzfiVCvNTbM9hyQLwOC/qFJX
me5ONwn2Sn/LMFOiz9OFtWm9RbuixDOmY7koMSO3EgYwOeNtwbfbYglaEJUzLEez
3E+YrymUcjE3xzwanHg4Ybnm20VfLkILM9psGszJKPmqxXAwAjfdE59Sn0Xw8RAf
I4DXBQzc6BM/kK4e34zE19aTnMFQs/EicyvaPRvtxkcYZc2hsieqQILPevckvNQN
onuZUwxwXWLRXqFizatm0YskgPS0w49FKyj7AjacfeDxM1/dmBmzjX4XqiDiNTsx
Qt03BBDI0jhQBidgmP16Sb1LG/WDti+sC1Nc9SK4Jg86CayYzUMSXLM/Vw4ZHFBq
WEVO6546nhkJuWWWz0LHQjEWmCOI/oY/9qyr4eWEiNzQ9kPqCjzQzzPRYInmX1nw
CygPGz27yEw5YDuNvILSZAPBw1WNXPAhLaqRT6412tY+b+7SXCEcQxeaXVvA7rbZ
NVLJbiEru9dwMZs8CbhaZg/OXmB1yFQKiDDiPK/BszZWOq/QLt2g0bs6n4DU6Asy
l0nhaShZPt/snu++YNHJcqgngoQEWAXRa6qf+QkKpCT/SNXW3dfAje5oxEinFHBN
9zxLB0a3wDKNyp7JIAjks4m+6JrgJJ4f9STW7u81yE/wRj/xFzmb6N1quZ4E7sVM
8x3BewK+Tnu2ElKmFBW/qiiQRSQ9Gm4PzDt1EhuZjvEfIua/Lq2B8feH0g7+WAtq
wrftvmhQE86dcRAFWl2gJTsIetz+5C61ksvHGr9fKUE0gBQrY6jqpnXIXMrUZQmw
ccJuapD+2BZ0agg1EHB1hDFiHL4A6UVUI3P/gox/ayt6+DmBBRZvzelAyxjbgSU4
swmw05GTNsQQHbAbcswU3vPLgMxb9Gh2ASpywF+zXOgeGvtd19pukXhC7JFfQcxC
a/uWYQ1FARERTGdlrn8PbhyNCjGsqjNGIuaYolbhCS9khZKXUY1Eu6cy60Ru1ieC
7OZ3jxdWhoTwDTiACkDutx0rSHK4p8ifsp626c5qsvOZ0BA0EAVEwdve8iwsDYk4
igAIDv+fy2n7Cj2uIi8RRe/EHlJ+ym02bbRN28aOEzs=
`protect END_PROTECTED
