`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuybwMlmI52Yvy6lx4YQz8t2PRbejtx3cbIgcx5yNenvs0ccZXnaqWGhzk2q6/Cm
bJ231Aj8dgv6OlwMRoMUFy7omCy5NyN59421M6TlApGjVtIoltlBz8yflvOf55hB
Fd2GjkROECJKAAetNHqx2anHw2tG6THs1LpyPfNrvW0XefW3jvaLUXw12nSofTr2
d4/ZRuf700oLghLywl7RkD9kP2uiwQhOhnRcu6sZMM90KerlfgKg3qa6LtTM0JDG
dWdcA8AAtUlBn5ZKhNWICz1EPe0LJm6KNWUjhjwbVgk=
`protect END_PROTECTED
