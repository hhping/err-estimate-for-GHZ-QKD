`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZA628SKekN9ZRamqxBrpxGsUtaWp1UX64i8OpWn/AYib7VI+baSH2jWoCDOxFAl
eF5/ire65TE3vI3gkrAGMfyE+yYSrVudE0hKToGG2hVJwy8ZOpWewjRar58cN5Xs
1tnIrXZ9rOJlQvuZh7a0UaB4y2P17cEOriqhVQ+GHrWM021C0XWFFYak4W/X0xqz
7P5nGwmV6bECW+0eT0JzwZxa68NKSgYu7vtqUdZIMmrn042Cys5gnJa7moeHyzwK
2s+T7KeD5TLJxbz6TJuE06mJz81VMDsD+QECuSGRy7C81g0a+ckOZMaDgVl0aRDX
KldDDtW636ZBG5ZMKO34N6jmlgoKn9LiCnVir5gD5+MTqG2vqpkv5KGt3ob5T9os
DV0ZKD6i97Gn5187u7ZYd/y6d5UgSzRnGR0JWGPKrLwZ5b1bjemYrejOojQchy1p
ToVTuGIc/nI+TJYsKSQxrJ0ZKjjpCYJ9UMt1kK6YogdUKU4C7ZcGKocEw2IkswiF
h1aOcG1e7+FY+8nY9Qbwn9SHZfCaC2bdDAdkkokgzDnc+6q08IOyPXXjqwzvBGRH
fmehB2wjLW2/Z1192r6dA3wT+39ldnkYVXR5DsnBBWpBw6E7NKJOyn0Vv5Y5dyZc
SNFkoYwXY9wbuRVfOPMyKxZQGbBjanEWIfzC6BjSeO5JA8vt+XKDlqpoLy+c0I2x
9GbjxfJrtFZqo0lDkWs6AvKRjBpn1QNMl8hcf5ke+tcwbNytTGudQ7z15Of1VQtP
hyjsF4Jo18yeVdHMWQfDf4yDGliJFWudtLjoAlqcYgsF6XQbNBKTV6h68B7s1XyG
LVkjFPw8h2IO7vV9mTm3ziwPDFsIFTJCkq1Gpi9u+qHNaLqRT2Dga2rBKKLHot27
HPtVbb122Su3z3Jb/hPTLcwMMcD+/IEsSlvmJ0fGI1+6a0pXv87bIna97ZRiYM6l
XDxEL00W19zHf3T4qseG0AsOIjLSW0xnU43obXz7h/i1bIMfdEJHjh47SRrmrvBy
WJgh5Es166n734yatZj9hJcaezSBY9CJv/panpEqa7vLFNLS7UUHS/miukXG5ig6
`protect END_PROTECTED
