`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zacwF+VmgI/9sRxawztK6SHCWldi2Zmhd+IayP8W1iaSdnYj/vFlrYPoJWLNOmO
u4fQaZCJ8hdKy/EdEXNAQgycJhdcsslzp/RnOlDOoY1rGsQnsSSlxrtViE25JvAh
bVkL0X+vCUtIG9Cwq5jvmJF26ar0MFrSNjvuv1SNG7DLgHyEYTH8C1CF5YfxGgTR
iKbjAr23NtTnaVZyEaOrHNsiYXWzbOF9KjoSuVNVE/V0UM08iCDIiSfzCZrxTqXx
EGhwRXBzAchtP+pr52+MO7RSt3nEDezk8aGm/pXRVLdU95zAo3zOWbCFcV/wi1s+
GZBpHw5M/swScr1uMEcuIgsF0jGpuNuFsyk0o92MtcDlsewF9hDa1KBjFQT8q0QL
fBFiTN8creGZ7X1LG4uXZahk+GlVzk4bHPoOihuqxXTdl2nVUZ6O6+ZNrPfenJDy
U1M3uoFEZUBzCV7WUWRU5Qh1HcCbKEKzeha22vLGao0jBIQ/A6x/Ls81UI8j4caj
a0VCaIJ9+Tol+kFXP7IIr1WmDiMkwQUzvxFmqFvXqBlYqH7l2abLi9G4/27k7Ot/
X2sVJRfwEmv0U30yoMT9z5mkgtfNMeiKK/pPBtvvIoBKlC1lLhBDGddtKvwEykIC
uRQqXsdotXCiZb8Py3vovFtTuCXFblVoWBneOoiCmdtzOihAk2IdJbxodhKlTwcq
89kMPytFvQ9kgf7MeuZ+VIV5oNiAjKxfJ5Vb9YqWVy9UJ6Db97xyCXgQwMPHO26W
5//Gq+ppXAZFqIv3Vo1FDWzWsmKOyeWHwqEWPltfsOwwg8cPXe44QE30vGJos48W
7rKIcgZVGRK3SERqS0elNfLFYb265wq6cvrhZ3G3g8y3ef3E5tHqX3jYWmqA8Yca
0rDsQkfuu3bhmBxUSR+e+dIgbc98jzKLlfqpdwBUgPDP3TXB5zJhlHHN45ssCPCZ
Q19KTrGR9RILqYEq1Vt3t4xRPtyOKSuY8VxGgt4GhAc4hEFefqH4w8u8mmIIzxEy
JaxNLZA3tgD5hC+H8csFldYcv5aEzNHmVgHKl/UDaZKzqOYxijWs4HkjcewehNSj
x/4DQAYAjMn1qPFA5w+jaQLBILVGObLy0X8ZRwIE6qxbqoBWrUmDx0OK/MshzZfZ
M9D1OF653oeAfMvYWlEVU7a67kFU2QsY6Q6D6UsTLjCUlWwlkeux6a3l5cgihiBA
bxZnxJARltVF/Tsed88Lwp5ZqlmLISLBEX8R7yKDNJ9f0m4P8kHAz3y/h6QR6NK2
Rh7gZmDbTuZ6dqnk+IWOCzZQk6m+mI4SJUoh/aCaQlflcysGYm4tReu+0wPT55XK
JiTbE/BoxXw5VdeKI513X4DtaylnUk0CHx0qMNCSZ1dMBklKsQBa9q9Eepy6otPs
88CyD6OtV/5SBHBF3Eryf+alp32933ZKQpzd9atwWVkV5Xiv8XmdTsryTj6Ylsg9
4xEjDVsbM1mY/+owT34JGmjkiQGG9skkpTOfAJLk20l1dlZGfF8yhHoITaKg0BmN
ja8lvgoKPZ+MijeO/F9I9FuHXtW8AcR20FLmhObdu+ZJnNRLalwCno1Ifizw7GE0
ZbY9bJM3goD2dRmgfTGKREhNMlRuWeVdFnk30pzfOwhY/dcGraHIQlGKM9tuQ73D
pey08xnntLQSBSLVqaUPyp65bqwD4GxavzRI2y4GdMaw5vs6qq7V6fFEZUVhRt1m
LSCNT33nrNuPBITtK9wUDGUuiWlys26NrF00Pv3NKnQ87Bu1Bhy5eMnAu4Jx6+Rj
Bf248G5IwFGbRa40RrIZjcI2uxvpiOYSuN6IgL7VB4jjbfglIlyf9w3v/NEkc6Gv
G2p66EkUhyvAMlKRXIwR8I/HjhuoRl19PXpZL4bbVI+YLgeA3cWdrS94txNv5Q21
WeeoKnh/5OGDnxRBHg75MEl+2GoavWUdeYAJ05viu4pWrFkooiAA3doFjYsRlVYd
sGIreKsX7ZF6uwFn1b3nB8pv4XQPSgwRZJnz06OoAEtzhPR19pM+PBi+qKz3YOso
uLm4QdZ+gHA1QgzWX4V1FrA7TOhD8ps1feD6NiT4pKaUwiHL4TBqnSrlfpI6yMfv
Py7PLWNOm8pooxil5jscKYojMI+L1qkTjqc2JCQ3901vqAthMxLIbrmh5+5ZfERK
lJwyr2XQI3l6AQnoEGG1hopsjyGXiJshduVoPucQWZqek4PT+D0l5TWfx8A9GPPU
M/DDPH9s7rBgE8kwNaUteMyZgz9hns/p0nOEBgj25rTj1lQWHynZtKv/2YnZ1Lkr
A9xt8HQrGliLnD6diFk0JgqKBeTyDs/jG7xLMBU4GddmJ1GPsP47P5n2NIFuFeDw
FiLMcmmQTJ1smvVJAGwNibOZTblK1FwkFeVTK05CcC6SIzWaX6bdCkqfjVTB6mnG
uQv7m6pJKCFidTdDYVm2LWjNTDcDBvP9TFjhJbU8BK9JBqbm3py9sgdrWL06PV/t
yZvG1RGq1LJK0JkYaj8DRAnWr7emM+ldXWB0STcFZkm3np3ZRGEu7yAHGSz4OuPD
dVmSWr+/0C+Y9gVA97uPN0tvxPa5S9n798GViZ+u2/SDvS4eI7awa2nHZ3gQaN/x
jBBxtPHkJM4RC5G/sot+U8smV9XbWXes5eWeUSAqlEXyehtONE8wFBewW3Mf3Luh
s9JNIanJQhjNc1u6PG9vXTZ1PqxztxOdDYNod4sRSnbAEGSmRGxCaFtiP7QYobcD
Qur44UTM7O01g5dP3vgurM/OX1m/G8msvD6zGBC9Ki4Gd9loz8Ldyc67OPQ0tWjh
+/I+up6XKQS2B23M70xIdYN9Lc47b4NaWOzkNtLUHixxWQI7Xzgl79FD14G9sRTk
absA+GHuCDbDWxInSdGUzyIcUT6pwfDv9CodMOy4XsvHohjjYS/CNd1mMr8VDfYP
LpKkwoqO4cppylzEZ8NDgiKUaZjxS5AUae4IfAVNjZIYPeQJUwUNTSuqLywvR6Ox
Il02P5fa7dMlyWJV+apXuUpLIkLRfv2YiuCSr+J7aUxE21/N5hgTRCzyVAueuJtb
khdXsywgPkhDxzeZy7jyX+xEE/caz6umO07xNvzsnPPDP5hP3GAjHG4HiPW5xz3A
o1875Qm0qgtVdDa/nhJ8vej3wBmH/1pD2vhHvYN+w92fujMyGUQyIMHbNAHAQsvx
RDFTE4Y8+TCuksMf0JSRvhWQi/df+8V36lzGmpEg/k1Q1Srb3kBD/XEzrMgxY9zh
TG++phQcyjE/g+472BHX7QKtUc2JwhA14ku7Y0gtjgJ0yJQ4h1Dzz+sGmnINi39L
A33dHrMXQHze+Ibpu7Kjk8l1+mLaxqBB9q+zC8jS1I7CI8ERXpR4BqHCdCHdr1mv
oYCQRMN2xJ9ZnQf9CvPjFNOamTjPhKL70OEAf1gX4gDW18aGBSXAf2f/pedyw4We
ncHNTe+nEkOsl/dxl5ZNHskom03e8DVbxlijk0UGPPd6wRIL5SpTeYiWyzTXOish
AWIDD1y4TFppTZwNRkwavy3wRqE7t8oTtjA/i1ubLYEWQ5Mmk6Vxig7uzfx42CAw
oanCq1kKNbNHl3yOBjNB7BkRCrrHVTELqwd948gHV72LQXJ1k8zJqNvW7cmn35C+
L8gjEi+lbx4FzEdHotkHBP0QOnc8rAw2Pd7bAXxWe47syGG0I8Xg+dqtDzCP04e+
uhLTwdZXXnEAyDq5e0muo0y2yAP2MzITaxONILKzVSlGbq4cBpNFcDBj9Iwzb2Vq
IxIXNSnBA+fEMXzIYLpPp+uuY6BHnSIfe8IkZKWcrsQBTVdcQ9rilyFPUBe9+bPq
Cv/bm+Onw9pBRkkCAr4b2B7qhkwgPs4oWo5hqm/x1a0eksXRBpSj/FaszfX1FzOl
usIHpxZejYdlNpn+gyp4pMD1WwepNvSDaPK+3esjWzb0ch6+tOAwxdCOYN36eFNh
3Y/haz+bVjMGMjIkO+5W6CzS4gc7IN7ESkxQ/Rq1n0Be+L/707909LL2FZb3LDFJ
S7939jtsPKlxcDZY2KUhDIr1ZnueHKmxogIOUXQq4TeS4NGE4dlOPctjUA1gnvsC
CX7k6mvJG1Dsrup7nTTMzJOT6f62Uj9+17X8PbSkvYAqYKuvsJx4JizkeleZa7QJ
sukDUp4HMjFt4C4mJTcCJ83n2lx+Qt6TzYyzpIzL7I87oVQmzXjnKLb0JlHHUne6
lHTrj0gDXm0MJHBXe5PsD629Fl2T26Hwc97lnfPK4H+eHiz2IHJ+wEKEDalLZ3Pj
0a5IHP588e/PkJ2mxeCG+9lNcUBXI5klRE3MO7FRrdKHM/pwSYPxmjFU624CioDO
vOIONpj3h4pQjTa6WNsPD2H9JnMiTLLhKIWMiyYlYZtiuMhWSWmy4sPpybsjs+94
3eBItQlIia58D2Gho9KgTijQZPWrwz1GC0QUyEmrT69eUFbaNUMiwRluluThj+Ok
rXefxAE72gPzQkoohk0q+UGShNRINW7+F84cRGH6Q/a19ZidWS14KTf6RhEo+tWk
vc3GjcRduhwM+tfLZZRg0pQ29xIYuNPa1TLH5gjt6kDJ34IGeB5NEJzV81L4WGw0
GEfd5yBRd2ggI16A1c/4eTCBsz1ZgnjEwRbNtUzt36EE5z8Xbg+OjtbgdjoFU5Jl
+VTCX66hagx1TD0C11HYOkMi4AGwNjE615ptmQiLFkl3TsR2NF3dkbTvtSgPNLUQ
39JclPrV/nsdoH6oHnrTegEMa5vP+ux7HoIE73JOnTxXhGL+UwTvQCPyxVWKr9oZ
1/0R93EgtMn3HnrgoFt3d7iSRwQynQ4t96+qGYw9VJCo/f6UGAl2BoxvqX2iYUNg
GbcicK60utQWvDvxuQJAWL8PypyUFnI5FZfCIN7ddLtbxAl/nB+o6SzqBxRUXfHE
DUAdfekvb8hcJzEDGmH2XVnaWZvjF44uxyYP9KIzJ2iEYF20fllizrb/2QYTa0GA
8c+syyiMpCTGagTOj8Sk+a3VuPGvJo2Kl/KjZ+llVpjx9EXmfzn3LqiiSadslrck
sjxaXcmfTPoYqOb3qxGSszCGBvyNPm6Mq57m1eiz1acwHIluesFbh3N7VXL2Pkpt
I1rOaQ9bvKIKuxnN3aMwDL8GjlDNfgqiWy9i5cfCLGV0Qm2YLyG/9mOT4jhgZEYr
VhVwik8ofVcxdbwaYF7OkrFGDo4VtU0wXXXwpAurqaAU2j3vF1r5n9HKp3tkdm0A
1s+fLeCtsBswFc2pcFRpl97qM1b6uBQn287OF9pIL4NYY5sRMVPDX24RWLDYliDT
yxVT6SOq0nryLTweAJBsQXle4snu3jROSxHLJoPn21O5UM5KkabB0+446nZswgYh
8ktsbPHaiy5DlodC+IXemXr5UgAhdT6ISGpG+qRTIoP7mrjgPKR9T2Ub8+Shqo1p
UPKDEErDkzDd0M1sR0dOZswzuTi1xN+iS7qyLlgC0eVk6Un/4W0XJnu93YuCK8kR
8fwHrLv9Mwjm0zfODSw1qDNUKsMroWpylKO5LZgTjqBobxP24qOAjX5ZnUKbb9bZ
fqSRvSkI9hrrV3goOG4SU0IY+RNIzsRYcRzKXIaP+xB51ngfCenloGQk+Ks2TeG4
znqYeMcMLTzrX2/lDBdUIXm8efoeOzw2nboeY+eeRBuVPcOsHQ5fneUr8txm5xV5
81sWYryEH7Xtn9XnyoELYljwFr0NYkSghwUGtE3gpKkjqw51uwD6pUPaok5AHaXt
2v41paZowyc6Ql82SMKg+fGnvn8atlV1nK+BLtmssLVp1jZrSR1c7b8u/ZZAH/IR
cBMpKdKZ0TAdg8piAN/Vx/tiAL38GebCPixwo170K5+CvymqxMaRlfuYOKCJSWTO
Q44Xs6k6VYomRYYCO6RUtiv2DDGOqfKPEjxvnrYSXvL+6ktDmhHA96nM0IEGcNma
9bYG/TrebKiUzoqKljiLL5IEM6Suc8gt7OPpCrlWu07XNWcyOrMYnkabWZlJB6NT
3pxN8q+Q1sRQX2qYG5jAwkrB/JF8eQd6C/9zYddrL5a6fgte1iWAGix4ST9CJnrO
Ai9L1m2iMb/qYfoJylNc/Ibfx/JnrOI5Pe5IxcYOs+G9ToijZ8QsbTKlFqqOk2R4
O0wHPxNDhx8cJXB4sU3FljJgkpAVhlekqIaqo0Cip8TaXf8YKfk34yDYk37OhSZh
3xhvN+edFn7q1tcKhw9SFjFBMYEAyUFhf4FINPVGVe4DsaLTt+1xXZsnBG5AYRoS
UtCeLVUvpHSO6oOsJT4qi/nE5opKBY2CUWeoJl/dVHmuDj/NoKpnAdyEroAIXzx2
OF4NLtFmCYzXsBn1wqB/dsVC5BhpOxfvyMLAIkNfP5gLAHDOMpxAXqrcBFo9siMt
j64obi5EfE7YI6S855IhVtZa2WQnj1cBzNmATA2Jk/UB/0ntpXv7beoD4rcrs4aS
8Q8S3KuqCeNjyPVRlvR+FzRqYy/SdWWswJFmR8iB+T12Nk6I3euPJwlVAt6SG6Ic
jCYRb9OODQ6QdZ/xXVtIklIeR8hsWC6w2RSfL/itvsyPUssKW6gNB4Yatfem6BUA
9+LJj2l3y+OiYlgPn+SjVDUT+VV9WjYShvoZf+cvgKHgF8D5JrecDTpZOFSMBdna
0q1/mxt/ELRtyR2g3uLE9StjsUjL8f5QMSHTNHrsh87lCSpk+Im3yd9nVf90XNhx
Hqsowm24FoG9JpMRmrVeoRRA7AC2+gvhOEFXJM0FrEZ8YGZMk+Jor8/3FBmXWzdB
zbDyXx5e0elcBeZpBOekfQDeew2IBkQMrs7r+8sl3IfwK/nOHLiuVZkaPuTxvQSA
bZBl8Yth0wdH3T05d1UQqUehKEg0nNB2hPMY3mfUBJxawUP7H4M4e3GtcWfqvOa7
sYx5KmWAQNObbXZL8skmgfNfM0usiHKl/DsymkCBbukN4xa/c2NQWNnjvQzCJ1/9
3eLciOLwGY77F10c6uSgpO1eIWMmE0nAKh4h2KNFKTFLU/lycVIdWH0Pg9Uw7rr9
/lrwkFYhKbU3k2BFpp42xf4gVddCeUow/w4UBZdkrNL6gfpf22qVYJa26uSb9GbI
JGH7mgZobO7rDsojb97M0uQgnme7pj0hEPCb6TiH6Kp7TCdAQLDe4lhclY76wH/B
KADXN1N24wePBxAUEwTLgnn38/GHQKbO0Xop5xgcvmCiASiOw8AFt+zDxdT864n1
N3pQSt+rEWbOQw4wafrRD2vAM1xPbp6LdzmHHBhqRmW5k393JGpE4CtZeWtG6rs8
Jyk4UKA2Ad3zLQ8jGILlgcHlJVn4vVR5DE5PunV3VueOzXIZTExHrEUnoN4BDLxg
KqhQ/v3TQfF43/8vCT3L+TjtSE2A3LVvI+LcT6JPqsCVJ1CjsTvzq6b2Xu+jqNDW
QwhedbKIN9R82gj+nUiF40K/7iegX4VY67uVMylzJhzplKtqvWa/b7dJ1w30qZTC
ve/Ggr0amYZ6cCet7AhMGirqih4WzVCX/PxkUQTzU+Cjnjy3bOkNYDCH2vYrWfJv
VOXLN8iZjtKCJQykGSEXdlx1Qluc6Mj8IL18sz+YAvwffBVplXOg8/Y51rE2HW89
o7ihgRBG6T23WIemZSzfSDByrXM7ugEP0g1vRykhesO6xeJ6wvDK9KpJjIwru1qg
k8NF9kQUd8zCx0vqdAvzIbVhI/RJup60nKS7oM3llsuXvymgXOPRUOHLze+DouMq
kTwh77ioLthw2wr7sJJJ1B/0+TSiiCJBncAUXKiP44rujVAaKOHBYxPkmavhV+Cq
c5shsWXSjd+R/QPny9UjwGbEYqeL5fGP3nTVuXXRXSFboYUhU+hdGVy//Y1jQF2x
IaHs92dnneuX0ODQtI80QhLlB9lB/09iIs0vKWNJz8Edm2zhCwJmm3xTCJ0e8ZV2
6+OuL5ud1gpxtiqQFgBNJzKZDUugPwpl4SqkaXNrkRicPMhDJYPdZTLZU9USOive
lvZ/GJsQoeLaRwn9qUBKIEmgumgpOC0xbb8Wq7Bp7w1FjnXWrHLYWo0OgtFQdYXA
+8OcVTyKg3MEhkW3enYm0q5lZRSOrYaRl3zMJzsHd5TJ30rG1pAbhXiS1Zt4FKoV
IqUNYfPofHCQuE0Sgqc7WmzEwhCmNgjlYYPQs1/uLG0XfrIhJ1uFaLV/Z7Z2f7dN
J4Zp0A/Szy/LN7I30oij+CHSe8GgfPmeChI5Et+vyCccW1ZbgoEcStVk8aZRbneU
5PbEeGgh6YxKJ9TIbqgrezNDRdxAMlXW5EuKORCtwmHqUhkrYW170nzgEfDNek+l
b273wdX7nT2CnguBEBojxMfyYXhq7gmrWsiyjK1BEzys2ICxbNfMuIZcS2I0oEci
VJel+fqZBwSZnzQDLiBE7+XSr7Tq//SisThTsJeJAD+ZkbHUK6qtaKhkTJ0ZMMja
ovkfh6fyp5O2KxCqrvrq5sXT5X+qbyXZWb6TRaRFCSB+AHv8bSa6R7ZySFHBeLYE
IIjUN3bGZb7O0L36b3vmcYRDc39yCMGIN9e3o1zRHYfYpQpjSb/AUWG2QsDLwKk3
/Hj1G0TH6GiMLKf1zUWsMXUlP6a8IWFHkVd4oi5THbF8yEihYPwf7bYNlIh45p6o
IZzDaI72DuZ/+2TYZduQgcyhp/+lV+CTNpkEe07YFrAl5KYGQYgeNGa7PXl6kvcV
qB5gMPINGYGRpVdJwajU7QXy6azDF4svsJZnz6327EF4I0SfrEKOOvT1R+23Irlc
VtwstKW9SPu5VORPxwbf+LDK6j/YlCjd0zhMwJ8P43LqihDyxnnPK5BloqtyAJT9
/g/zP1cFM0iVBFpg/qPuFJuwXFMOG5vbgdL6cTOAiFVt/kkbZtsFtqPy7DCsC4s5
O3ymUpvIDUztxiLXCY/2gNBP2I4mZzDyTl/2g/U8T7zRx92GhaPoDkmmWxXy+v2n
APqSM2jXNZGLH/1P1FE71E2lQUTq1DJyBc0kF+orMY24SoaKtc+tq1cwyBoJb8p0
UQzaYhwCDiYQKoT7jZT8OQNLW1XIe8g2bTggpCmciQL735R6GWObSSipYoE2K7/y
GjGrGXpxdQ2DJ9xGi4yhutQjWwnLFzeMbLP8tshEhhmhbXRAGRBT/RDqI7QXqnFQ
ygYQ5R/UEs8rYDY4HF04nIvcI5fyZFdbKZ0ZmLprdBa00aFuHhBrEgxCPGCzUw1d
NUCgel3vANqORaQDH0l+iXDARsTRVI9jL0VFHyMJdCoZbTMi5p3FBowUVll/KPo6
WVzmk+gSz6LDt47kAzJQUHoPcWseUuQKb+lGzr1qPRPS6vZf/thAt6A9af2Oa4qe
TWpr6ShSCwJYnXFvjKr/a94ZNgVAzVVnIbGfefVgzP5xFUITQ3bLwI0hnvNAe2Mw
ptTy7BFcgqKNuAzZEQ5Qoeg1fJofrSKpKYW1c7oYJQPjNxctYXj7vAxRYvlQCB0Z
g01L6A1r0eSCxtbIBAbxWmu5rtf1GWwKyt/tQC5L9EbEBNHYcaVEl6xxU9hxGs/X
mj+uLymcwNlQ4s8m0mfiNpDqnN+JPt2ow4IS9tJ+CW7I5VJL6SKk/1EeWUw5Eetf
RkOgaXO+QsYAeo+TfP5evFQvYG5vi54wiHYG/XDdc/VzCKXtHMoRE4jItV5OxQlN
K6QWhycGF2Hchxv5KqxL6kJB7xEQZJvWP3/KASAg5sXSdAuQHOfBJXNvXFTsyigC
ECzWHxFU7c9lkuWNAnPuKymuBxiMfLs3ckhgJGCSs2+f+khDXNFHPPpeak6olXEJ
omW8ha8EKRYXDFAvzVo04opoKsUow8TqyC11iIvlcqh+AFBLPebbyAdXILISYieL
kEAVXfTxRw3PmAJa3lhmm5RDQBINXyN7+7xkL6QY8rEq9UZBClaKA7P2veeElSG3
bQm+9yPve6As601NOPyVoqZw8AzFdUegHu1VQkV/szz47jPDkdq4JRyHOJVMSgRP
Zcw21fNW656WxBjHHZPMQP/mCYQYhR2ZznFcTo4ZgtsAGoFhESkJBq2z6FIWo2uD
BaPNdkCEJbSx8RFIrn5nvz2tpsnj0kjmbHvRilNksJI9MIFznDE9WRZTVvmmJyyT
BIseSnZKYfp5+4ocEE2je4VcCeFh7p9vBDroXgUsP+R3Rp7i+3/QSQkwWxVQ0U7b
q6RDoYPXaaLXgB7g/q1y/9bzRYKUOaD24eazK7okzFu8f9Q2A5M4jaJVZQr7etBz
BpJ3OX85XSvnt80fMWla3Ah+iPwkUHOckLof407Kkr6xLCczvt/2f9aAlCLyeNq2
9611B51yppMl6EKt/Erah8IK1xHmCK9pb1UOr1Pp+FuM9Q37LIr7cYJQ7VLjA4se
HW2pQ6wHq0lQw0gSXTnvFw60qrbAxRffRoSvBivQ0qbbxiz8WttSLcHKwT5puGYT
q21ANoSTCvW6m7EueFQnpYDKWEUqyfgyRSZ76q3xjD/bKhpOPpf919B6YuMTzKDj
acFLTCMT0QF/7/T7kScxxUkCvzntlIMcL+jmgZ7mE50GPGsVQLLAY13pJ1ynTJPj
yuukL+OUT7l8fHfvuNZXl2c0ozeYe+S0HBfEeNEzisEZ1Dz2vjoamOiRRwVtenD0
NZSUlY1ONpiBRoyzgLuOihBxzUGgAaPITS3N2KEs/3Vp/pd4IOX8/frN7g4VQyun
TCqYO5tNnINOGDLGdr88d9nvfoFsUQl4o213yBOtQD16YGnZeqVI02Vi+FWBt6ca
b7ao3SVMHhh4wxVzywcEuoL1uBsRY+RCtB3f4ODtwu215UxQJdN8HqCfg3KXlOAq
vJJeeabTj8pX0TYXDWpfuiiaDQ5v1tV4HK3GAXJNHNhsqsYDoyWQMqHpHDwH0VYS
eIUATs7pYcpEDT2KawKV0eDHb5clblBvqCG3Hwe3/4j49nC8LUQvToD9Cr/0sYiI
noKMSE7oo+LgN/eHh8R8R1wJgGKx57Yt8pomnrZNqtUXVpXpAK9LPpyWGhtM+xNC
Hzwx2JIecMOSTvVkSkdjR8/2WdPUucl6kIGCvNFCcMblFflGs5CIQ7gin2OI/wKw
QEhohvFSsSKbnHGUUnO0Hsco3lx1YeKAxjJU8EceIRPuog5jJnC484e/2xADqGi6
PFSAkNSc7qQLd7QaBBppx8sy+qWdgeUKtE2yvHKWuJJ/2nzSZBn/StxBVujYtzZx
Ro723oBxeoutVpkHU5ib+z1ZpNmMr9eurTadjKfgd6DwcVbJvxeWg+pFwwgmHmlx
Q62ADXs78zr0HLMAFsVvAI17IqAwqQ6ZK5vxPFiw/vhbwxoTh9AKwjXQLfVOxAQQ
+8ANCiGc5CNHpTZI5M6RbGMkd+YWEZ//h1iQdjEWFdzZNYE4mugkVIpdz2W+GWRC
YaJAxxKA0BSfODUgXPcbDzrfQTtLPL2UKgG491Vq3sJVNl5kuD3kedwvpJNXhKwe
Rijg9dv11WAqovI5IzPP9lqN+eKnSJiygpuoSmxre+zaaVX6H/hefKibPJy8Feic
0pJsSBTczAFkbBIS9jeZ8zNsLmCOCjNFvLJrfBwZEHrqArwd/stplOjEqXvBam8f
tPouNfUhoAHFAIYmIEPwJb+WnNw2+XGrQS2Aq/t842shSytFycQDm0sjPBJuBKIF
FtlAvl/tJCAgZNjZI/jX209kk2hy7Y/jZAzi6QLMxTcbowdZyBjjdZT4uA2/xPgB
07XjV9vbUizwNKewS821DVN9BRmCZTBrtpIG+DkUxyV0iNh+VYTdnh2Dd0yuHlNX
pV6eCIedhyMq1yvtt3QGHV7VX15/E68UVY0TgtO20u/iFEiQMh4UBlhkP1fpGZtW
zxrZR/B+aObWfJHpxqb7+ROp1o1gWJ2NSA1e9bOuobsygUGqIIstFJaCwpnpdVhO
y94vgLiWpGKtrGfBufpptqMAJeZMh7sLpiIkTs1iEl/Ij+O/r3xKPvKM/55WnjEJ
wwTe4siPh8YoUXjAC0VLHbm/tNCVXxDccSbvXyxvnwsf3z1DMI5OPlhb7i2ZcyFm
jr11j8tu6CnLXY0L++Bd6ADFhCKQdOTSjGlWtkarZsE6+EL4NJ6dqTmFW+HY3/mf
UXPxBLGqhFtM/fsqF2bpLhv7CvH4/1WfnjXqPkTB3qqemNf+dMSzUU8vD3u7Ak2I
Rs+luxpt0W/uqneFnpQudsHBg1nKs6sFUw/yjX0P/JLwkVaemyNjONbdu2p1XDQD
5xlCNjlMt7GfRJx8gOMMadwgPwXMU9SXdrtB3H2kx9WHPDKYDO+9lEMgHV5YelNg
ujYqFx3vKirDsNRcusUSuxvtHpxsLW90qC6fb2gN/mWvzmA3XxFkasJz7O9c+qB+
h8fEhZL6fYbl1CtQ5wYyg51uz2B4JXsH65cnuUnANt6jBqmgPIK96bpp1EY4zTLd
+aPS5skm9Ex6pyXFJtb9++tOT79vknDodKSnHS8T8PQXEk5J00jMF9+xsy4/UXt3
e40nuDUEiyLJSfraa+8EnSPflTdOvIm2TkjvrbQp5O06PjVTMYxIoMaclpOaCuzf
9w60O2EdFRTLdhnt3JGsjLL/negkXbrCyynSB3iE/qQxHVtlUZ97GdWdrzGgomie
R+rCjcee/k1j2fsjGqa6RKSxDdvt+iByPQyxTm7dUxrgDds+6G2Vv7b1jhNYscLi
tEEm+4i2aGtjqxfcMfaOei7FQ95VxmYphvpxulKiBhVEzLpjGKm2JR/kfjVYDwDe
cXw4RWLytz/uaIxN++bBLBmpmHzLJJCDWvas4znQCioku9qBNq2LP4LceOiUf6wM
akijtenXDCSUSsREXRtnDdtMU0vET/3W5hVkDUMrzC35A55midAwq9Yf5JyzKs97
jHJLyrHe0I+RMZooB3biZoX3OwGBY0X7kQrCLZoYBeMKu01Ze/u3F2zLS+t+zJpG
8sf19kRtgmcBAWj7PEytqZw7MFRi5BpHrK3dVX8/RnbTZyI8fGE+pK41Gs4sDDYu
jCEhmGyBOjBOpDedQyrsme0SvudtZr1qr/RogRw/zMC88OU2TarA8UE1aMduM5f1
H0vDiTVQIHVimTp+xdwp1TRMpBIre5jFXFgxWFnfGo0xJ6gnrtGZgx5BJwJZn62v
wwcmF9HE16xQs7anQxCwK4CGe6cHOg84Rp9JULJHKhFs5Yq5dYTrko7UfSnONcv4
910XP2hLsA0dhy80N2mNFy4CR1dplQskuGje8S1mvri1teqc/qynhl3TiiUhY3cD
6QVHpX+ipEfHepe+cYTj4gLNwojlZoYF2wAz214pasue/h5L0XasWh9C8I9mrapb
ZJeKaHbgSvjnwGqCeKfRIiJHB7eKZFlWZRB6M+DxC6CfvQ3mOYjTDW+k5uCVopzD
cnp/WIVMHc78ga1yx0B4I6rJVipneacl4+NSN6b+vq9W4zVbSP6HwfP9FwjnOl6M
/qbad2sqwD5D46SBYiJn2NWd2SmirsbG69dll1Spx8DUt1ze4w9MvIrv10iD9WBT
ylR6k0wF6P9DF47dNVK/G6l5gTOdcopV89aBrjsx7+tXYGqzP3f1EwsB48xpG6eZ
sgNqBvHhVpBr680mqVQR7COhdPeY92LtvHKKpjVH0w7sw9q55FzqGfBwFrYzxveW
5CuAsYvpPkY7M7bY9Qf4mfN0jcRflMOilHnbCQpC4GcNvV+Z8BqKgvcHdIuHkgTI
y8eijkvjSc+hEh2Nv+wHgRfzafxYotkxVYCgGAc+NuFFfu/pI6n0GBsTLK8uIK39
h40NrzOhl/vs8/c76AcCeNayEbvCBUDLUhT7ixSbbgsFs3fS5cWwo4goxAHppah/
6nD1cGYdkLW9/Md8GoNniYfm5ItAV7Jz1VceYW/u5jaoVCGaCYKQIcAIxNccjqkD
2mMPKnO0utfCBy9IsH2ougVSrjElMGtx/dIlBjzv6R0LK1zpSJHnV3v2fdU4m4YD
epApEd0UqwtKeIlmFm71OdKjzq3ijdeZGkmMPT8jLOm3JiUyKD6Eq2z65CtBhG3X
pQI5v6DwvdP/jjKELXddQ6mPJV52a03atJk9DdPXnuSqDOf/m5hFnH6FDkrFJBYW
1adezdp2AGjo2CTYX9/+eYkHnAoISlvoIZVRk8rN/9BeiVGcHIV8d2cKTSZxYvWJ
J//HSiAReFlbK0yyIR208xiJce7mi62JtOSRX/YrWeDixvaARBtAhbAsDXg+VPW2
btEs3Ic/zRtIQotl6dbMVb7O1zFG3An+2sgc2vzkOz9gkzfHBEG1cadu/1UitrIZ
8IwdMjgMOdv1YT7YfYGnEztJh1CCf14eVx64MrRxD2+NvnrDQsSvmhBbD2GnAq64
n+CidxZSQcYz/JlxIV2/Wo3uioPcL3C9BLgMMtxRJmDSabakf6rq7vKgirtaVGC3
Fwy46ZFUoGE/iuRDUsudOiXQOx6DO/WWxXucq0iWuOfANkD+gWs+V7NNDgNJgqq7
k9aXxKswQkV4/758wk8HjFwhB2rphuIlQ0SwzdjJZKdJasu0w1GavNAksNyYDbIR
JO+87FxcAcyCCC7xT7O2mQWkTcU+BA7NR5BgfQgEn+U/cS2W/nDJpRYny6NWShUT
RIBK+2OwoJsoyPrps7lbPVwY5/+59HNNz97j40yi9oOEdGGROHFK9q54p6TcHtSb
+DtfipQ4o8OOSmKADtzCFXq1sjQ3JaXzf6vZLHYaXovuI+VYwWj1B7S3iqlsxu7a
9bDxmjwwi8kKpY9HEIo3u68rNq7j5oljvrh5+a/fpLekSlEkwv5BvSNylLgyXMRa
DDLHTom8Cf8RoVuRgN9ZG6ij7ody3L5tUGxV//jDTbQ1P/jaH7yl35qvNYp6fGM3
vM/MXaT9Y+plB3LjVJZIGikqvNmTx20gxafqyQHVvNL3py+YkEHgz1YGBqr9H0Tl
beX1OJ5pvVYECeJxNA4q9aJvXh65lXsjtgP/1m5gKza0gcaNKzx7n9Onnb87gizB
YD8oY674an4SEIzaFCDeY86Q4TTxXJIViWqTF1LwkZAbkeSmsdQMEJABa4CCzMWl
mWyF/wer11IY2H3XRK5VETOneWbDNIr05Jtwlhp++YEiovc+jZDPkGmY57DDjLG2
vBoTjVPu07BTL9GCpZJ47raQGl4jmvA2Ut15RUC/ZsaYok5tnsY32IF9EgjR0/om
o732OwIFmc+VGQ1J2Sp6Ew/eldozQA/Qg8h1yK+SRyQ5JkQkQnPEExmG2hnE6SOW
jFKm1I8Ek+NvAaiCaPio0YjTFHlsTDpT+RRrwMmQ6yaHuZWaUx/N4Z2XGoLP8az5
bEDLhtVCCWrFIl1ZJ3wXeD2MI5r+/s49/KEwVO760vmUtRTQtJwRdUS1/yvBptsY
m46OGex/hvTfsJf8ghboO/jCtEs3A7/EaDp/7Y23sDuZlYhqZjVGq6LQQRBjlG3y
ow4oSd53+Ojz9SoU6dKL5X58K5ysazJGq7rss4FSDiWA8YkvJGT2KxejWY0h+wYl
6w4RiyLK2pJPO8CT9nu95JZjJgHxcnbMa+0dxon2ei8U5Lc274rQYH4AZvb19if6
d+GCoOoLYhAOFRYbsl0AuzqYieyMFKzp6+hba/f2X92z5drNG28CW7basPOqxXYP
e9CN8fS+GVmGOuxmlTuDruW8RZHndlaylP0vhyKfIOqi4L0LgoJGD3nk9g3LveGZ
ToZNIM0UY65zn8Q+zX40WXiIstKYhgu6Rz5AML/JlUkx+V+0aQQCSPA8JgZvTKcJ
8wFo7Kl66EIKyCy2qyhx7NjBH/+f1VPXDxOChOkeh80l2FEh13AR88ddCLFiLs1h
jq7mfKNJWjvamKuCYl2RLTgftQ+/XYcxKCl4xx0nPFSvM7fpfQfhPBlBZesDd81C
tqLVDCfHPdxQs1VTEZKI0/zNyy7CjtmZTurBA/cXpw3NqQwt+32jBtD1OI16EaOF
ZLeUabwtwSIuYKuQWsG+NHCtzBmqQvVeNAKwwpne8JfsTKZNu0ue0VYjX5Ujp5JU
IvCT8punktwwJhxag06Q7ui59eWpTwrvzhY+1Ro9Gz4Qwn1cfu2x2u6EmIziUeoh
oWbpVopqtcDDx1Qc2qdbYWJ6zgOXuep83Wf6OsdOKAhSnTz2Mncsl8keH/u3/ukF
4ryCHLHfbzT9vY8m94obu1Ddpl2Lo4Fa9HHm8NwlOh+JwB7XUsN3Jxoll8wHTxhY
d9bn3CxA+SsSN4EXkVXy5WxHtCYOad8D5Z9Jsbtmr8BkRIgfxEyKS/eTLYWt0UWy
P23gX7BcIvU7mSEn1mPfYsFaZakcSxcXVl3gkIcmD347F+rh35G3rdPYbfErvGxs
qjQHvKC82FgLUBK+PwcsBncf2COOABkttw9a8Z6W+up8yc5LXzBacW3sjYYAkEgW
IkJCTMZZ1qDQLRmKMT2EEdX6owlEiAxZLYGpQvHyBOSeBKeyDJAXj8v3O3TsH6ma
FDznVm5j2EL4gAWB+QjStRC7R/9/6ZhZVwcKDjo7cvIdSz7m/TR0HSn5VrXIYqlc
7Ora1K1Zco6AbDGJcQ47TeVQt8CIQ7pfa5k3hwE6sec+L8g7Veuug2SqKfnP5kvE
OCufBWZ1aRm4viW+4pT7TpDMSlrynrQqP7m7tahQrlQ/0qaXHTVQERvCTCHA0e+h
oKDB53YPNmPVHKQeYMsqK3v93qNHw4zcfIYGuEnfy3OcKq/+uEF7FyVfrOTSDsZR
FdhmJPdG7yzI2xzDZrsmrjpxZhYs8thU28uFNMsIRVOvg3IzQAGBqrygnFB/U1J1
yzfyQ/BFmWg53rFEOaRkyik0lNpLAvLxVSc6TSfp0FaV6cplw0o44TcQTThw4XLL
kRTarQHyx7+9YQKitBw8dNoq8sOqrMwfaCZTSVIzHSA4qxTKrv+O4rMRwzN9Ydec
qJUFEe+uCRnut1PAkfued0j+jxMYkj1/OW1Ee9Df4gBQdOatvHNuCt3/jeE8bz9Q
n0EsiDFTuBA1COnC1yJhvgBrZl/RFtGqBc1Vq+nrc5HmkMBmKKvFTiH3Exa0OemX
b+b4zCs2pga/AQmSwwa5Mhk8f9+zhZr9sr0qSP5ITMVP9HFPWa0kWiLJr5Nuwyii
kP0xs/hfpsfD37uzXbG7jFcqEPZwnorZJooFcNl+WW6EgCN1FfWiLKaj00ue/YUW
3B1cQCcaaoAXdluxdxSwYwWdwwBmY5q07R7fYU1BZfaRWXuWgNepzSkTir1Ikv7G
W7nudICMrxMaqiftYgY5QnnIgrsKKu1PmPyoFM5NWcaXstPfdMMMzKgMPO77C6uH
QEMZ/q5xocLfB/+UklTwjKFiLiQpQOYhUSpDPouasv4JqLm0FZfV8hGKYkS/HYOz
+IcbSEoUrdLHcviQi+skux8thtJ/AD6fs84v+Thm4Cow49B9hSoGP28RsPaMMvi4
TvexNOjnCUd3WCbDuT6tRerpvokN8xapPi+DWnbEjlOFxjzpV+AAkizmNmtJmQj8
FMnL1NOkPjq1XKPw8GVPqI8aOVGP9nxGsYWpi1UoTK+r0OdWYJSCPtzKu/eRTZFD
yPDdDxrP/V+X3cBDB2UgqXRYplPvr8c9HTC+fvAbN36ibVqNVs4+1A/DTZKf+ojO
Kdio+b3SJ2ceLt/GUebuabcGRIicxmZcXXRU3Vci2xCQcYlgjYPm+00hQZjcGzxj
BWm0En0x28jnicpHbHqhHL2cEIt/rern+DGK9tbqQEDRVrqs4S487C1FNvSszYCg
uOwFOTsU7fABXovXGRcVkAYhiB+O9gt9S8cPzkv4jqM8tRiJGgkZKcCUurZW7jN3
Wqxsa7ldD4yWeZlMw2+YSBs1j+3+Kb0/jpuE9LtEVleWrQhdZFRZ6rKtol149lxn
m8XRtInOZhgBEAlClgmXCoYcmNV6XPJJkRa/59OwXZ5quigmKFRV65nl6+5GPnqT
mfzSWIFPJCYwVmeRSm6pAQNBtB4EBI/ON4GgelpqVuwH7nsdhfA1/58GnR5aGpST
ChKtRtMEFPfb7FV/NhE0eMHGPsAjouvBeDIKf8j0nPD1l/huV4ChM8rGmFaoFWHs
fzpTi9JYEjCyPe83oq54JWmlRYUuz7pFmAQAcMzZ4Cp5dDMtWREDiJ4a1Ewc95wX
/aXIPqtnBFzfgjfEGks4Nbc0k1C2N0+HCOjS0eqPScqTZyNMvln2UBLUhy1tb4j0
qdVFCmN7wdbaYZw834IZXg+aibSDht1E0yXsv0SuggcvocqHY2UGNtd9wl/kc+/0
l363QgwCRPLkBLzT+p0QQ450uRziGvE5JgKbpVmDmZBJ9hlbgzQJpFXEsGPUTP5a
yeGWC4NZghpwkr9qMabUZBOHp4Fz6zXxcfod6brVGnqFhP0S1H8uIBb+mofwf+L5
E4KwzG5/WlaWGP/xgNsXgAl6+qO49joA8TKahwosQGy6LPRcrWurU7T3HZpZ+qwZ
r17HMADON/oFz4xNSxdPH8lAlR0dddvhuc7dLLs8/3XK28d1y2x47d2JUmWOVkBy
UoeW0xAcaxLodfNBrGqyZVK1nxcoamBaftkCBNwoHw/IXsTW7wgnCCCeqW7DSR6w
3qKFE37edMDhM5ps8Hc5Uh7nhuHTNscB8Ibw59zp29EsTEt+OAYS2kHPPGUdFg02
m747HJKVBbSJDI+cg0p3fYwpdPGJA5qX3NNQM/PhYG3yHvpEFnmpBXCBuaZT49Pd
AKHweKcqAJ2fS2V10w3lgcJeLegYylomI3Q+955mL3x6rvTjCW1cT6Rb+kveInPq
yo2w06S9DtumgnQs7+XIHUX2w9w5rrUdya4flPcimAcui/y0AvH2t6l7TeMRxFMQ
PXf7dTq3kLSZqLa9Dv+TehwdJhuvxntORg59vKPAJZvbc3tfyffEOQNds6l8V6mP
Im/eT8yILKaT9CTISTMO8gQKaStoz3CTrAqFCHjyidxjSTXfI7Vy9YCBI2tnj4bi
sbMQrZcyWjGbZ5Q20XdalaD7r7K1lrcRshzq2iif/aqITOKYUVYenX+SMOieI6J/
fWOs+evbc5B0UaDnRU3Suz+57yadMBohNpVUNj5LwLBQdd/LPs0OQwj3QL2Xfxal
SjfRwCiqago1X742Ze9n+pcdSxsib/f9c1iZhYUeGc1bE50VlByEp8lzbRb5h9Od
ac3REu8aqKqQWONkyb2MHXjbxDX9JuzqMqGkaGYzuEGkZfLxc7muhZ4u30HGqtNV
NqlJuQplvorbyeoCFGDLLVrCgoKB78azwLlA51p5A5j6vANfkq8Bh6tYkQq9G+Mq
4pDN8MXtOn9z3cDLhYNn3+P/tEGiAvT506el5HF+OW9ue4G29zbuidn+OsnwCat9
BxPH25617qwqF9FI9CqitoFWFZ1+3oEl4y5tEXUKuyIXnvy6+S1/nOnkzRbZaiiW
OK5q8qF06/tEysVap6bEYS6u9i6HRSuTBWAc6D3Dri63MTtV7thu9I7YP9a4tGm3
Sev/3XI3H+i+ksZwUDlFREiZ8C4fKsqQGm6U6KWnZvK17MIaSrQiPb+X+oggYer4
ER6rWqDfWnYfzntw5p0mR7flcorDxZbuYiJo44aPtp7bVLSwHeydp5tIqMdeyQVz
xTy59r+q5FUiGuE/m44Ha5e/FVZVvMDZvsWh3JZRDYdeMx/7WI7W8vZWJxQJ2tra
EcOMS0smhJBd1WQ7atfJQdXAQXr8qyGCcj22PNuNtHPVRvNzVD4o6cZ6ujaq4rXp
jhSVaYDbPAA31ewrU3laNpKQKg91aPREvDZS22MinamZtLJk6EYLM/npdqH78efi
zqDBZiUw5cn7zZ6La43BWZj0xYgjpwVnXaXUdlnAWq+ghM9C2SpX3GYpC8gnLAOi
OMN/b33ekXaiGl6A5gO0hSkHqF/9qImjbB5R5GqRgFwjaOVhNi9eQvZfsqlFVvpG
/+YPqyOTePDP8q3JKs/36TyVoxsxmILwtzrd/MABEM3B+oHGTwmnDngKt2wuYjKy
uXozrALYrHwjAXXP2pNdckgsnTOFPs8m4/RVuTFrECTrZctxHb9JPeeKYMrL7rbA
mdxU+Wl8k3tW3R+luG2vZc5QSFFbin+M9i6ASZqN2d2U+NUsOZTaqebbhSbzE6nL
hgzeYxZo7GnF7LqZitmEDJZF6a8kSUvdDAfFpX+dqbWFnAe1LrIO/6LPIe8qoBYy
Ut2x84bxN6dF2WmrW//zx0B42vlnS+6FnUhOhgSc6Z/toCHAAzUm/E0zqZxdSExg
rIVYuxQQAGP4zIZbDGXoltEPYdPSUE1DPoioO/kVcJUi0BbWw4i0Iryv45e0//hj
lw3WtkrRVc4sVHlbmu1Lo6OEBJqypkE4i5+6af2CAO9WzEDAti3BHOZ9JSzfn+NH
n4CEqjZx5WZz09pTvPYFToWUTIVZzYsUE5CJIgbtmjg/cg7VFFmGpfXzgxLmF+n2
H9+NydQseoharaCBhhtv+zRZFeHbNe8srlFO3SDdB+ose98w9lZbX/zbhXIszUVI
PRyCxTrLXqmzU4p4irrChIxwalldvtYrpNTdh9KUkuvS/348/pTiRqsUg8g8firZ
uXaNGUiEcd0SMx1h4ypQ/dvJdpFOm0IwuiKXbMGVBvY04YmtVPfscQqPs95dYPRA
B1zMoi8b4B/M5SRwawl+/I+ArE1ncS4OrkIGNE3dKNfrkBENLnF8Y1WBhEPeQi20
dui0sgMPsxgl+hSNdm0vpvDqPBNWBCXGiMkGSTEXQcfEZRhUPIEe5bHuY9jX8Y/T
nnIOOLhiF7iz/0MnUAirrex8mSLdcNB8xfSO8D/NUKrO+48mBu6E7rM3nJ+Z9bKj
S0Ju/72K7kd0GzSYYuHREV3Wt5SU/1NBhlpaYFAuJ4HzpYgR2rMPiPkoIZScfEPn
BK81LzVliq5KoZFylCyvtloMmvzZiY668g39e2DpWdj8PrawjMQ5zn4nuxxveSEb
w8BHZqS+7eapl9QY0AHNVzJpTMEgs2EzcflEuzX9X0YGpM6ppU7MMQqn1EywRrYL
Irar+cwNSSs3ql7CJ88TmYF3eU4GA3gMcvAD53osh8kix7I+R2v+BOQq7t3zFcTL
KdsH+sJt2/Q5bQV7tLUqxws7ExftxkDPUE6Rs7p5gpnvAAnpm2uaRI0HANQPyQvF
BYCF/DpHEbeQRzjAoR5X63CSCCKNcIe7jX2Ifra5IuYpSzXnvzKQXQJ1+i7sBzBR
R+sClEmlM8gmpxuyCR5rb+JNkcpJiNWL714PO7PVcRNTSNqYNJxMoGO0DVSRLnHV
+mNr6p5BgFD37yWTDxEYIpP6mFRqv0G1tZx7Db0vxBVE7QfOZk6lLo5Rn317+u4K
dkjrt51riLWepdxKCyddeGZUICLmKlQm+TNSGKZfliMbt7K47ZMjtn+U9l2WTrMH
vOQuNu77+9oyW0V1FR5wEaxmI28R091MeSqNpgfGEVLWrveURztQce+8sHqLTKeO
+OefEIR7QR0J5KqAT7OpwnaEh60J9EdS6hoxi378tfkUcIDpcwrZcGlsh0otBeLN
0Ga6DMNYG2zgU8AuGtS8RZ3WWi/JIZ33ibmUh4RtGRzd2iKWIVC8fn2k4wo5iw79
ocXgUj4vh+8UK3qM/hPtE7d3ciwmMYIJ/3TVbSeglMRZa44gnPo8v6KAKIReRBS6
hfaNiEWcA6Z2+xQUlFMDpJlKFIIB3F8ApcyGPmAtYFqgL6Uw/va7SxAvDVsG31Vk
sxCoW1sbQjxFYbKom3Z0IiNWzicMqGDljBh9OIADCHYSoklJ4kacXSEm6wmpCJ8Z
rUf4OvkMsdgwj6Zt6SqavzLDmZaorYj9jnH2gjdDtITKgJvwPoPCScSkdlk5NFL7
4i+5WWUv/cY4oYviHubLXo1Imsx4NooIQTLBldgO4uS33mSFq25Qfi99mFp6Ji/t
1f9iL+pL7/UJRTR5Y5vfl8FFaTjbiojFDIJ7SeSeO1orevRrWm9sLDnABgXcRXq8
eAUoRJlSJF9ysRnzOkCv8Oiy0iSM6OCfEmf5u0sg1GGDgDj2tzHvklk6I8AlvY+H
5mnHNUaHprecnDggsmzTIY908YiVivdp9Hrk4NA+4CXtrF11uqy3u6/mzsNLQe/B
yGFiXvX42UH44GwO8B6wIvxgKg7NhN0jn/U/KiQYbkGMCOKc3ySIWBI4sLvjgR0P
DzfHKjuwYuKd5BWzm1x3vNkNYxkYQOX4uo3Xt9k1CbrP/VSSS38vhhdcJpLPqPxI
cF6XwFK95NzhmU9wQg8o4vKsgYgAMq/J813mu7AGawM1c/ipCwZMXucCEHWSTr8e
Ej0TKPuUy5qWzG5QZGwPhYBSjOfjZ/JXff8oU+O/tu5FGFiraiWUVN+g9NIYFci3
DMyUarhNw14kkqmkIiNeVAP0LhCwv+ReawUhx0h59KHrjVojEsz334Ul8DDkNT10
NE2lxdXG4Zw27JSzXkBxLp2uk9RKTenqgLnipMruNsjl9fuwR5ydcvI0kjaee91h
pOsmq+u2HmVXK/DmIZFWUlrjzQodDRhNwhY5vR+cSWJ4ORYVYyKior1BXh4d2g4w
atK7sJSH3YH75mp5skYH4RBoaiukmbGpq9Bvz6QYQWEOpwb0+5bBkyHP8pH5jTjO
WYOdYD1Gu8V/FNeT3B59KQPiHBBsgs/RYrNQ/qDkTFpYzhQuTq64DQmlqokfiJE9
ztSFNBDVjrfApzK52/vXZvNsZix9I5+Y+CWjC18HJT+zWMofWsehWPiVbwGAZFQX
0lMF04WCxyrNmeWybsjSTuruGRWa0tIZEEaL8Fw9/MvTMM9Z28M2Y87Ir+QkVjHO
ZlMubtJjqeBbSv60OZUgKQxpOENaeeo4ZnixqKUTZ1ZI1UpYF8Yyb82W82cL+9dI
krgmepnhkh9GxzFB6olH6kdTArs+A6zaYZCMAzJ70fXdng6AdMUximevp42CPbW4
SPl8d6Vet3I0BezHZbiuhQ5HWLyH5xM88HphYnJkF8aMebW+bHoI2RCsdggKpzS3
eBVtB3BM9075NQl8uYhbq2NSs6vtrvQIQ4YqtLCFdC/qmjmO9b4RUcwiLrUXzXvW
LR7Sbkbq1dpgu33L4aHYqEZPtOGLZ+VzjAc0TQchT5kLqQWZSFJQmIsOqU4mm466
pdxh85UdROlFzFDdjdo1I6N0AV83j1KDGd+ajs5qkpLdQtcdrAUTpzpiFJfEapb9
MjJV/9bD206+gulpeeQZo52qxpAUxlUFJiabWfseGq8loodWoFZkGVIAq/jcK8F4
zD+O0allGkQLJtLRjfQDe4KDjyO0Io6BghwvvEXeOBlNkkN3rCDPZH6JtY0KVHNC
vltSx4VsLAHvXkFh4ZRO+JzKCUlYVjvGLFdnmj4062XUVOwjsLa73z1Y09orXI0t
SO7o3w9PgtH4vB1Vfe7oB3j6zbvV4vKp0QPJHfznF88snWtO1xUec0CY8RtiHny5
kdGkiOlxETB1P0V0OosOKQm9P4Agu+UMPm2FAhrumFkizKFGkc8oQanP1cpSGBHw
MTCLJtw7+QuYYGU8XyQGQssl7eSSHZNBfvO86LjZbteksVdEGNL/0hluHk4uJwxl
xBhjXNMFgWGB/X6+Pz5eO5xkb+1mSNstpJ8pVMoc1+jy2ycsqDJ25nKCzCpYOpzo
xGEqrKfJx8ekuCv3drJtqNv4i+Hcmc9iU6MbA+EmICjjOv4dsLGRaoFIeLCSB1pf
GcZfTilH3+Cu9BK6CZbdEQ8Fd3uGc6XY4JpUb808WDzksGBH6nzr4RaPXZx9mdBX
EEi0CApU18UO99KL9mc5Pf407TjtN+9FpOTYRpTj1EZ0E9r0UoSAR26KDfyieqv4
uO1HmTTzbaB4uRFHNYZxKyKvFLo/KUmdSGIE1mp8HCbUZseD4UQii8tWOWoDca47
tNSyBt8rXyzwHEpalBXk9dilOxk5C4CPOvXC02Zf3OjvRIUT/vMFTp6d15TRUpCi
TfOvhPHAumeA57xKX8i2gr4IGcCYOlIPruCi3cS7rviGb3Yefl/tBvdYFoo+mAwL
DogFgpxlf1HDSFgyfXTBq9LiB2LabB4Q58qkX5Ky/0TENbGU1ozi1xzW9UIRrMA7
ecstgiJVEdVZTbDfDRBqiPIWhDXgh068rrxbgz46ULDlMkLeTva+Jq32ttf+gLIY
LbwoBBMhnfZ6el/anEXa06bQJP+xbKX9PJwgFShZOFnkLkk+UVUaD+1HVjmU5yg6
mE5gtA1Sx3hWbRP9QtI9oQEc489etct6Lof5HU7Vr5GkgeJGg35UaDILNnQ1r88X
3cLmBaBrXj5h/ZfrIrrkOf+3DSPSjZDg58amUsa8HOD0LBxfeu/m2Y6tqe51aBwf
vQEL4WSXzgpU3782XRgIGM6ZTz3MqvoALkbrA12h7WIVR3p9ohUhpMNl383wG1D3
hyoHLkyYC2yYNEBFChOAhAgnc2l0gtU5HZFf8HCIucBSdqWxJ617oX4SEHKbDV3p
L24BeLtlwdV7yLe1mv93TdyU98SSdVU6zmXwkhHDa8l4uqyQ77c27Zt1SFm4S/qs
g3u+AutlZgkDKxCn8fJlDU69uWNl0WL6Fcf4VNTAdXEK9IKX1M3y4KodQIux5R9z
5SKslFY6fW9ZeLpPaHagKqO+QKSMEvF0s91kh/czn7lLLJ9ZyzCRGhOB3I9TsGuo
LlSgUSBiYV1BPYC3oz5/xtY09rkbUednVCm91LDZ/VjfSKlbesurIu2i5wBlptmt
2E3TD8sTgqTLShUvcyFdrs0snWF+KA456j97Tvvm6HdIKEg32rnrU/wWmLKE3u6H
QyTf4/AJ3Asz9HcrX8/ToAVBxGF40AYdpn669lD5bMEzdLetH5jglR+UTaht/mL3
kM53R6bqFG+eXQ9RnsZpclVEcLsCsRlpKihfsV/+L+S8lpbmPMn4gAb34w8SiPIA
aOX1OUbjHgBoR/TjE33R+yqxWSB8EZswYZFwXHjYpUO1m6TBZv4vHVhaIxVITCA1
x6jend+apVRx3pyWsO5TCImctBrA24nvGdOY20dkRKxsMJo2kO95jAedsSfTQQP8
47jFyoIq7HXHLH/aEIDWnD0TVY+kc9J9EJpxKYTNbQgQNrva/hxsost7dk2P5mB4
74YAgatxdlZhRjsvjXkov/BOPMIM5AylFXv73ORa6Mr8blHS7M5yMHmDTz27Jh3R
reewNCz8C6LdnTcpnwYZXoWCjTFUACv9j1qxXGR5p0+1NIYXM0mgO0PRKGgvla/P
FcD4k+3YeO5Wp7kIYwro6AtWVLnmUSZFzqxYM2kTMKaG3TmeTtBaBycrCWtjujLi
yscRcOjdnylVSgTVZwDforM+hNR/YSjUtML/lAquYpY0x/DiyJzB+iUNUzDvGfRr
gep9FEtgaIEAQ/TBBoDjB7lv+IDHmQevKG9jklfcFgp6E9H1k0MCplJSL6KmeW3h
lST0sF+LY3PquxjP+Eanao3b9b0ZdzuvyZ0bGtHZTYsf3xsJhesx9TL7F8GWzd5J
FuuYYaAQqh+b02KKE2MtM7l3wRrYiQpvvN1XOdrMAsqBO/iiyA4S0r0lokzhDXRQ
aPtKxOufMOvDS7Z2iXCBogEJlSJbD4ifDI4yR2YWTBFYiKKG7o5kx84b0dCfh25V
sP9ihSgU94GT2fGkW3jqFKaBEHXXrV813LLRok/gKns72EvYYkQ/Tdy5pNjaKwtL
NhtBYXjstcp2mPU4iiDz7XEsYhJAPRY3Q+obVG4LA6FxlDmJY4lRdT9bNYqtRx4R
dXvR8kxRGiQGVwWZ33p07+ZKg3AqdRKESRvYW1US8mh52u1jefkR/ZjGo8V3tnAj
4wLAxlRd/XplIy53vlJu6+C/8dcuHbbDWknJrf6liinfTrONRT9fcZP/0yWuqwrI
1NGAHKXSRvfXMeO/E34N6iFMBBroq9l7oSmFBr053xwyb65IHr/syTnXRHeIQBfN
Nrzpaa2URSEoDqvDDjpQgB9t2/gNoA/34hgXitHqtMyGnHIs1chEJDhn+g68DX6i
tGZTFqkxDOV7x6Inx/aJS6a0L1kntXjnJglw3Bc4pNln8NJqTFEvU2xFh547pGOb
EqBkVR4DllzmsBd1MMDrj8CjpMvg7+ZuYXa0ukqRj++evIxo4+wYvJw4GBfsizPs
t/8yT/MhYe78tOLGNnOEG4JobRHZbToFbDIfPgn5Ba+YMxXj4IDWHS8Q1tSja57h
5YVtKeL66XXANH51NqTvoQ9wGf+O5fjeUKpfF0FGKDFoTD9coAvFCfHbbY1ygpWM
V2kRXRk2JjACtyP39xE/LKS2U4LRIB9UBFJp804iOeZXIQATcYPAsKeg0vR9z+rt
G4ccqBjg5eMuZBCo2isos6mQqbF7ClQ+hcL33qnDeypEk9suBvckN5Zt6VTSP16f
CO8KcaDDs1t+P/dw/fVpWrNoZ0qKRrFWIS5VC3dRluKZFFTgKTSdQURXZuSKzHYP
TPILtCZRz0BAfp2mcRjtRDBMPS3NkKrzkDfqQ/70GpiQkVdDl7IQqn6HyYc0NUdB
WvTwI+kgzFeLjsV+jFm4R3AIm1ri2dkTTrMx+khCU4TYZLhMLS6zrwo75MzMqIA+
AD75JqLUU6HF8tPjiL9NFhKnfw/lQgJ0AiLPPvUZAgpUFqxAbt1P9sJDOdyUVLEf
mipndg2E3BsUYzDEPPCySVnPdFX+rqbSplduh3YZZHEqtQWqE5Nd/O+O1mi4+tEB
DfRFA4UZnpaYNfaknX8r6Jvk3lsH8lJ2MPY198knyZZY0yUhUkT4yP377mq4HTVJ
3uVqoQi1T6KMjmgJextjzLY+ulaiaHmVoU2kGLk4y9grXkh8f98WT0q8Lr/1VU13
RCgA5BJpcZQfCOT2UwpBXDm7WAsqpHFIsrAaRJ9Ol87UoUl/DG60x/64NHljdWbz
Vy6rHueysh1h3i8HsliF2x4yk48kBIq5HTYb6CyBM7XLHy8VXOmk2rHP7KOGvvfU
2FTUPglUBBH9FFIcx6Zc6G0USGFgXAc4Wc1eSkbofZBhR7Oyo1NM7+Udlz8nNil2
7HMdebIXzc+OPbW1uq1M0stHvtZXgQ5+y5EYOmOXVXK4HsUtK7ZhmTQOru2Yp2m4
NjHDb5YuCWUfvDFkEqEaUbJI+0Ey4b1OXYgUk4l/HKOaydz0Sw6Q7qvoJCEl/LSq
Mi4dUIIqk8XmGX1BTW/yagm3DmbcME7vVebuplTilMxjE5JPZzgncHAZCf4qIUcC
pzOP5DOF61yu923w9SbxuL+7btl1LNXN95u3wmp6bEWtvqa4UWmmFAL/q6Ihga2N
Phkm1fp+H515MaAmmRxTnyDNCNSFzsuzSARUCa47x2X8p4X2B7pwTN33q9kazSUT
Mn2DG/VG2nVvBbcRkuZ9d3XcKMlrYhc0RG316nbkDNgSTpmJ3foIqO1gBot3cRAc
FVGP/rbwhUalD3FzR73PhZ6YRruegbIEne+kM9V6LEDQElRIZq82KSOzYhvioLZD
4R9PAqYsathAA1HurUBxXrnP7EjIdfU46jjdLRpyttGHJlR4aKZeQLkD9rHuwgbI
KN5O+x6cwV/6R+2GVS8XW2+1+IX6XQud0LIt7HHXKi2ACdXnAU9XJ9//lkXdz8Gu
BdrQ6kauX9ZEIBC6yQ6eX6kIMQaYR9s55UwvyKm7elxrB06lzZnKocvL9CKmOKoJ
8huS+FLdcTMiIhWD2LXAqs658OzGnBj7B9lmrsl7KMjRMRBe7OB2VAAgRdxwxqik
Zrj56p5tdHqaE40hn4W1F4/5brgJNvLWbFG2Ye+yF+qTJo2urgas1bEag6qNn4UD
sKpemb/luWzZrDfJR6wxFdZW+kTV4fRYGynIJw3QIsjgPWXi/IiFydMXuamz83Km
buvagYoFSP0DiyK9KK2xlCXYCtmtWwtw7v8kDck/4PZgvQfSakrgp7S8Eva0Fsg2
tJsYOM+IDXM00hI2vMXsIgKayx34QFSwAZlk4aFl49YqSwXjgtCwtyI4SV13MyRH
k7nnwNsrsa+wB11NHwehN7f0x8XIT2k26e8m6EaF/cwOfy9tTe5HlMNgPy9AP40N
3B4PZ350LRRdNI2g3BICoM28vuPmztYN4y0j/SyueEmTzsSwBb0k2SNWwWIQkBkJ
cKWh5XtYvqgob0Qi5FOGy7yTI0j5bpCgP98TEO0u6Kop2I7ONWaH2BoofMfM8QU7
7Vc7Abg06dBye83Ve9MBWxgTc49Tld68WNql7eplyoOnKzSNj/p9zaesXttxBuGz
KegqM9F/eeTkAo6RKlRo4n3Y8I18uM6AJweWkWMkSrR22zeWwtfxMEVbMOqsI2Nd
PVZJc8XSxPvViq4tIGi9d0yJKjlU72bX8s4IQMs8qFlDXzvVhaSeQOZx1OcFkFcF
SwND9g+pS6PuRU18aOf/DbM7pe29B3/XE6x/UnrjDIAYRNyQkz5R+TvwsE7qc/iK
+uZCow0uhGZVs2nTl0CJi2qc3f1y7aeQBhB1Q++LG8zbaqDaKdz0t4GTDzS6uVzw
JD4qxFvYEif52qMRTY78G0gmDfC+oXoCizvRZMvZkwny03XufQR/KAiuxU3fFkOl
BmWqiz12/MfzLYq/keudeeBHRvuR/fNZ55j9Ud403wvS3GSUXwt2DsRGaxVeb1Eg
YOKOSPIOt3YVSgeSEQFREVLzXDK2nyYI6AGWS8OAx6l0n7TuEky+YflvdMiWkRfH
SBY9mss5272quZmmIVFS2sWIiJyAgNy81AZhZTo5bTJRwU5GqhPDYd/4utAQQC+I
qFBV1hEULOpF1i0gu5aCI3530ZkJd2iY7kkH07r2XIFVzUPCoZnNzcurpHNtaN7l
R1SRokkSDCkRm92jE+UyJ8feDf5NLvtDLc7ApEU61ysZxePbLWikWsEIlaYtp3Et
fNicumpOV/yS+qtxjgFK8KZJtoeNFsvOhZHmB0ha1KxM7PfBWESm8k7D8tPjfHId
vwzk3nwyDB2mJPIxnwKNzxkVsgSvWWXee84mtr4HpsaqNhY3hleR1rs0ulte1Muc
OB0kuqVUGoyaLh9dp+tvhQOU3pMjo9fqHKr+3nVq0xgH5yRQFv1GxMcUJLG15HRO
jhCTVjsNHtZrXCzu04HDNdJh9w/ISN+dA6I6//dt9koHNwOoN6lEAWREYuFacULY
P48n2raQkh6DLxi2XD8qWVdPB0lby/3Ne/nBB/9LilGIX1U1ViHZXcr9zOutqDy+
Egzgdfu1sos2MkOXIyCYG0oGcjBo/8tHOn4saoK7oYTL0AEoWnDjJ5ude/g3OKSW
L+ymByaP+okGLrvW8L7MDLhjdYSmLnLlsFyIWY/8kCtZOJGNJph9kbqhA+cNfiSm
vH26/z+MpFeOwmolHsw/z5ZZBiSCLHrzqQcu/x9BqsR5W5ziO7dEkQ6JvsxOjldx
QkYMpWgMefAQeqSV6eIFqSBd3ctYMzCiJfoyKh2pSSz1q6GDqvV4ZkZmxubTYRUt
w95prJrIa+V3xvItJ/QDv3H3jRwKya9LzysAk5lvTtvdVjUYpIZwlcrAaDIka6H3
UYiGcX9IwG1n3fU/75K/F+XpCeoYIsPTa3bc85RMP3/MyVBqaxqitlRJzNYU6lOm
ajB6tqUJyeKTslfdUphxEXCH48d4mLCNaqgBGphaabiIgPqCwYKUYbqcYhlrtz9s
ldwUH4n/x0iqey/XEjGd+c6eMMD2Ie027ZeHloUXBjcJM0ZEEUXdzQMxazRQulDs
0r1udiWSCEGgB6E0sMzrebdG2ASpSYpb1rrGXxCbTqkkSYGudbbb+dHZ63UY/Wpr
tSkfkp9Jd5X9s7oXqYBCu+cIOx/blzqPckunPmJURYHF+rRYzfv3MaeEeNKlVd4v
S7mYmFCpOSleOZGeFbDXRQR7iEPh+5ibmCHQ3xRNj40SzBK47YedGMP8Y+0sHsDD
nf8CZ9Ww87EjeKlgZUWdstAWIt7yMtgkXQRuT/T8gx6BP3k8N8KPpS/Kifr0nP19
2/+C8Fg4+CXfB77yZxd8dAWS6d4aNXK6I/1my0oz+xM0GQpRleYDeCbDM33N6h9t
C3VBng9Yiacs8NCJr9Ke7WjaEYrlBgSRlERs71NZI/I3sCJCJ8wHN/GT9nu2p1zR
XpkluaTNohwF1vIXUT2iz7bHz5DM7oLuHAnwjw4smJhjILN+s97/BsHo4fb5cnTU
qD8K43d4ofgz6PG292stN3CLO2oSzlAc+Wfdr9HUU6gjyAUB8C501/1H48Iq71yd
Mw7A+ivepXul22qVI/wK+7R+adpGY9n9rXRYykFELCR7qXhMoy8q5+OEUAepnsIW
0UpcX7a5WKZAX2PYseXjfypMDG1G9LEDNhGIDDQ/IfrO+Ov+7WwwHhMm+Jy+Cnmh
DdgfpR1+Bz5KyZxwuaeH7XMsLNwrF+PTepPpIuMvFI/9eoTpNQl6bwYUM3Hr/F/X
P219fvcuXNzN60vP0EScrn3pUUiG0F9DjrRLNxzyKdm6KI7VIhzHS2hWeXdd5dgk
4AW9cvhg01vRJ87mR7sqwp7wJfX16Emkbp1Y62IbJKtBn4KS6f6IqXGHQNGimhr9
3dcaFrP7ZRsBpKddiGv7McntdNh+tguDU4MVdS9zMyRcUm4ZnUMzOtn7MLojZoSP
G0YBjb/Gk0b+jz35JCyDgm4KYfrJju19xukd0Kq3woatAUG4NS9xS9zi2UpC36gz
U9wRRInUjhCOOCDfnbId4Q2oncENMtrLJluBedOLFcynUhOusrhmc89UTdDt+TKH
sV+NXB10uz2JmnNDCN1cbVBo4fukGrZPVDF57ynjjRVEXBVe04rrHM+e0rTMhv1Z
aUmJoQzAyI8IzO+uJv5ywycIjx+t+ZG5WzzoApVtyxP/OJApng1YEuRm2N4E8ggU
kJ4VNMLzMfb4ZApUtDhn/7XFjnpWBlctigb3vqgt932zrS8dr0Qg5Gl5qzunm2FZ
PtvQDfPJHxoIn0DzqSkDyFyQgSRPMUWHMfuUgc5BrJ74Pv9T9/n2MxqLxWewrEPx
fxtm5+eVtAwsYvf//IDRW65TWHwZcDQQgKE3g2kMWiZSvEHI3xsNMQcXNZQbsHZI
xgRMF15Z3JEpxNmqLmnRNrnRGCh5nFxc8uHH3J0vlv2JJFn6gesvsN4+QdXWvWch
4PGvLfhraBeRgGzoV7UEF/Pbz3Qzcu0CIkQ6lYoWt81RWek7gP9nLeAQTQTePRkd
YRWz1lyf9MW6H0y9iUGBME6MmHvVhJRHgBeWTKxDtH9tBUGlpTX98YBnRC1BKBs3
oJxLcTFMpK8HMUDWXRJemmYQlBvYUtpbuR7F7bQk870M4CwnJnyMvAQFQsmyjn1A
6HtiVogR03GbGQSVRhs57Sn681YrSKqzS5MwzohB4Mqf4xnI6LrL29pcYrzJxhm5
OoDa2ThcKX4TgarsMpWw7VBWRp7HYpn9FGfw+buzEn2+zHAGrFNoKGSzJuBNICbN
7sT2+RE5i2OFaCEneTM5mTYuz+owCEO4hmecfUjLutMGVRvBKDCDA0jRZmsIU0C9
m5cnBgRN28PcYxI0glXYW242fpcgMLw3escBBdOcp6/QRTwKpYU/w05wHnGEe5Fw
ebNrQlFZ8h7SrbZBfGWygkhmM8uYKWpveomG4wdQAd8fEv7Y8avszp86uLNnevEh
/fcihryDSOqnk5WlGPOYI6OZnwUVvL/FaW99bsz+bie4tbYWm//gurGL+t9MU8Rl
4W2gIiHdLL7Qv7LUCxQ9+D0lj+A+1tHbOmrL5z8UFMTFdWkXhL+7smaZt4+ntUu2
ayuiZcrtehFLXl0YRakONSms8W4cNe7IAKhv5yHsXZ66MBn+2OYX3LC+GioyXguT
1GKbZJmXq5n5TCVcbtuf5q2ErWad/gVnraHY8Qm+uAfQUkJwy4ugXtf08JY+r69u
KmassMy/15AvSLTpFgFICGQNIal9bka+4NJk7dFqUxsVL5u5jufoPFwlUuddDR0V
5YHbIfq3ug5sx1I0Wrnwx/Hq5mHrJe/24aPLWsaZT7lv+6vyVMTU+aCY9tH13iFQ
vTLXLgKRV2u+Uwrt1WzdzWaaNNX4i1rdZdngbOm+vEbHZGzH4/cL3CtgDOVBw7WN
oCehwqKAGXcHJpwoZFTaNmsE5pziwWBOaoUvrmerhB15ugo8JZxdE++TD0X1sx7u
tIBNsJ9oezAEAWyqNHC8wqTCBop//+zn/8Iisir3iqgzug3cuzOnesToy+N84Mo7
9/61kpWzyX9LsFI0byw34fMDDqWsshNpo23JivLdtVyP9H+L26Xb79ZfstBlMZT/
BxRSV3sZaiJ7HT3XHRLD3jvEIZkxk2zp7Cmwy10gDENMtTpUaPPojHwGCXz2Hglq
hfkXg4lGSIyjeA4juyKeBsn03WWnYQRwCcgM05PVqvD30disaTAimQlkxEV2cNd/
1YSWyRdGzXrzNH5ZwSLMvEFt8Vql9Sgu7wrKrSmfWwroTvlmSAi1LoTONXzhZ2mX
Vv1hGpv95CayIoCtCdiw+cULM4efc90D3tqH9JMw13tfauqYnASQb1nLnelSBLGa
he4kuHq1Yt3VUqy7X2BrKH/5tuLEbWdnvL1UvrmPNGUtS9XWBTAoYrDKGv8H1lIE
G8aq+HXAzKkSqZSRuzyOHRgvop5UBGZku95ENLDzeF5ezMecrsLKvbvzHm2/W6Ks
evrQWOgNkxG5LSLbtxw+7iZaa7hW32MdBhLi2mjluzhGWJVnJkgUJZhxbN7NiUWt
mFAWsLIc13DQOzF8Y/i2pDItxnRW5GabZxeaatPuRJL43j+5BkpkjIbYsGpoQ5rx
FQSHoqQqc5ioN1YoiOkVxhNsc399I0RMpxrzX1zYvGRcYnNNWFIX6MN2Qgg1T8r7
C+LDUOWZ8gbr/sZ92lyNKKg1+98QDL1WIH9BxF3J3j72lKlMyFqUJGffrhexfA7L
3vE4YnuOdUClPridTjAyZUaLgDgKBTaSJPdeW2/neGLJTPzKJ2pbruzbXVLMaIjg
pvpd90QFrYu2184HtCze1BO7oa4UFS859YemosEawj+C0RN6yeSd2x+0d6f0x79U
U6JnRPMcDto2nZvb8/ZSJPas67Yk6+r5Ai9ePKQpoG6UIHCVVswX1lkIZbeIJzEq
J8g01dYujsxrraLvXq6NI/qUFQOUmW0ZnYxpXEgfuqqqDXvjsA0CVq+9fOrj9CEF
iJeCaWnmQeeMUhcCn4Eh/2jmzf6EjgB8a67ZRDZ1H2TnpEP8KqKSPS8ODfDWs/hq
qrawUerTh3P3gNMT3hp0EBVxgpIUrBHQDJ/n/LS+XS1FV5XqG+P/E1w14yUHmFlL
bZBTYgOPDuEidPn1B3bqoosERIrnCgosvdAK/3piy9gCeSQT9a7r4ugjg/FkraVY
HkTNetURgqG+0To0/ppPiPJuKWzYNEPvjCv21Tfh8H7ybKESzUpTaeiBjglzjNyI
u+pqBlH4xmv7oyRWV54YP3ALeWDgLGLSI/PNJEE0UaJtPv6gBHI6SRzAQ6a3LqHT
/2FkJa6dabNyG188g9zWDDgo2yXBOeUl3BO889krUGwcY0CuCQoFwYXh8LBrdQ5J
MoESAnmCvHyz9BCd9Ogwd2ZYPcJ8k2o2F/VfP05oAe1nX/vI66gdlg9+CC97V+vE
GCAuekNk9oGi/VSaWnE5ng+S7MXmgJbsa0dTGVyejT9AHyZEKOHUy7Sfw3jnTV+P
xJBu7+b5hMXS19RCl3dCYqzp7woJPpgbeQJHHWIbHAP6wPCHwwxF8jM4DJqWqf4E
QaFZR/GOFfnyuqf8udyZlnuCpczm1r9HSZhNJtk5CTFM5vG+jvc/gSrEwgxil4B1
2CbaisM3lMeuCjittPPevGG5fstJhcKU+9ItzcWVlb8VYiKFQECst6LuW4bCwhxf
k7LRqKGznhe3WKwpN20A2Na3WBTvV9ikNqg/QDoa1kVQLP41SMKCzGu7zlZLX1MC
pqvRz0GFXOg9n6lVKlwFx8znUT6JrF9GuRIZD00lCPtu+PRqymgRHTj/MmRIfjfw
pUjVLHCwYdpLTVIINrJCEyzAykJ4c+4LZ6QENSxig6kkLysfhSW1fZlUUwv1n5TG
bA53AOzHrRhoPGWJnC2xlRTkdnnDbHs0Erojn7QqQ7opygZhJYYO9jWmnwRuo3Dr
hFTP5QOn6IiW5LMfE291p1CDoDtW4JfisF3e9ROw50UQt4ya/VT+gludDCoL+64W
fb/aOBQGbxO1NWvKt3J43UdZmoT6EJ5ZE5GswI8xmi36GNTUDoPGsxmRfzuNxuI5
grrzxsGV9MUv1FT83D8bR0e+yc5BBuIbRX7FLVp8CbCTmPsjD8FiGaRgZROqNKk0
L8G0WE6LCoVmHOm08jav81/8yVyq9MUR0TqWdx8eww5UNpqNGBhuLbgPRC0i1XjL
XbVkSk4Dtzbpowoingx9NwzuckJYAP2ufPkviMPp5jYzTkbonkh1ODAtGbAFYjt0
nAr3Z0uULWnuOjTuB/8eGtBrYXJKxMJlIFTI6uO+KHLY4YT4IZ1EZKjNyVuqFrIp
QgpGPSmSG7+T5NwuV8y4b9kqpZvVeOpzpkl2AdFVbmj+szV4m1eNFmv88ulPq7wA
EQRGi7yNW+a/f3z1zIIWWPLXaEcR7jfeeqpj9WLXXNa+Yo8UbWzLO6jLLF+zuvD2
oo+j/7yUQBqZG3IUEWlD8rGR/AojVTUSwKhIO9J5pE3wc3DuvZJ06s9sav6hUdzK
wRwkhUjUKrVeWHYAfLkNhlUm7TF3s8x/2VPgS60MDwnibVqtHsEGKeTSmyDyj+Bn
4cVqYAhXeJneIY1v5JY2PFLmtcOsZNmvMMgLkiT6JHZRM7qsXtzAbUn8F4232VFs
UWKLmS2Sz/XqG5BPrTWAEyfqwfNOsVE8gWxrPf4DP0uOM5ihvIz0LFa3/b1oCK7H
NM0wJwDxX5JdhZvdhznq7B/d8ry4+6RZa5RyUeWZrLw8saCFMFj0/ie7i4LN1zpQ
sfI8A4C/eLnFZd38rvqghjQSKBm89JWe9bei/CkXnc9WDC/DqqMHdQUtCiNwRUjO
oT2DX1/5upDpNibCjy1Hqr6wjX8SEZ2UBybrPjSxuHNEo7i6g9Ut7SzXNX75+2hW
hzF02Li2H/kHBV0mk4xV1MDW0SKchV7j+LUpiH45e5KGOPTdLa5U9zdDq+wCjQha
YC/+pWXipYcRZrxMchyz2ZsDZ3wkXRlQfjijt6OtvzDU9Bd7/aBpxYOzaWkfxf+A
RM90U2jAU+j0JiJ0DjlxkxlIGhHy75jIDQNi2OAacQBHL0lKl2XJvsZlbBQCSF41
ILuqhFU+9KYxEossY3MuLfcfn1AlmMc2+dGJ8E4UVkIHvftDa/PyPAKXVNFO+dm1
P+IpwwbmTi3agoSynd51zRBaeUVU8S1rzM/nZ411uvBK9atGWy5xzy3+j5bql4CI
GV6NKrHjG2+FQNDwR/KoO+pDPOVct/mpAuEVW62j2EJh/6jiuLBHwVYvVpyir2dD
iymV3mqEhpsBMiE8308UhsxRp/9oqd1boFMPQNY6uurFA+bJbxlbYC2iCgmpqIpF
SvTb8Q5wZhFSJiZYeK8v1+Bh6/3/lhQJLazPmAF4tue1yduZ3LB8uKguf/NHLKfs
NFzYXc7TpWn3OA7uD+1LqoqdIjLHSPfeWQMw4OmMF+CkIG3NzflGMH69BhlJZ16Y
W63ORNXw6fghg+sylde2cHQgyksge2UbsLoyZzb1Wbb6prSs4xWm5Ca4NVCHPNSi
0xF8tqLinSLJGT22idFMpVMjE9VYxh9GrZKKuWy44C53FmOu3Q6SXALl9ts20RRy
bjyweP7O7beKSxN7LAx/rp3V4SmUCrgAHOczPWZXd+wBiqV/lZHxwg7unpBlexQM
dq2dQBdlc/Zz7+adSWxe84Yigf45B1cDE3RzWk60+a9k+PXRGGi7lspqIV33jbyn
omzR5N8mka/3YWLXZ9BgzwmH/K0A02pIZXRc29R9Ayb8sEp3rWsx2X4YyfwfSquT
Cb+bCFeiD9cFZ6cJ/qax5b0vCQkLwwyMWK9AI6gZPXgl+lU+4XJe6LcdafTYCpiF
F6I92IdT5RXyPgr0pV4oo8hqpJMtGQLDZ8tHaZBTqL5zQnu/BWm2Ql/krkLiDrXV
fcmYZ0eePyCQRYvhoSxVLpo638NhwvzSMKFVDVk6YR1JTda2hJRVRnAj1Qc19ABH
5sbNzBFFHR0AZbLC3FkuMeHsg+i0xzN9dKVWb7RNM9Osv5FsixEG8259oFUGyJMP
Vk7ZnItv9QgUK+EUL+o4/u9j25bJcqwo7GllFEeEYzHF6VHDIOPhg+vh9NyRC1U8
8PS86YaZI6YtaKt8RyV1LUj4k34e3HScfMSsqEalTjSQraKTkycu84NbIG6Yu5jt
9jHjdHMVu7COrHzqkUWJmGxKUu3jK9C8FId2Qf2U0WljC4TJclolNVDffh6qbAzO
APMQV6n724k93GVSfjwtpneEo8V1fr2KK09G2Q7O4+FC3v1AUgfgRhek597nZXRp
Bxg+q2tLMQGfF0FaJiWDH2U1s9UsWAsCcK/6V33tixHras/bTqoZLZY2tsC8naa8
ZMWBW6v4++zFqUKxeXxoNbvI8NmNPpTfX0igCofurw9C7MIiak+K1mJ6M5cn+uUf
TDgmWXcrnTCl0r52Spi/OCQ7vEd6CK3gSPw41M1FLhGtPHXTwWzktMe6NwVKZf6Q
EP0rBFGlNQGeAS04wrRti4bTJNJ68TFqbBc+2v6OmNB+OG27JbhZengT7ReL+JSq
4nRAEdlDowgHfpKJn2YFFT36lRNDU8l6aLeMFDbHAMLKDuFodiqVTknocbN6bZOc
xYDJDYOXnQLc44lpwCAfiJr3HueXTwXe/5J+LFlVqkMCrWtopAxz4+DOeDLJar8c
ZEGHSRVVn2S9oz26RbYwuYhK916L91Ee1OEsCIh5EijxjqNCSvWlKZ76RrMFvzFx
760At9UDN9fabwaPszEMLOinB/PoATggO6xj/Oq6BIRQA7Sf+Dg3cbKUwJm0Rm2y
ggSH1clFmEVwLVBxtmGQ436wFCzb+rXKarnoMiYL2QthG2uGEWv1a6ubAbmYbKoP
QK7O04WH0p/W9v49/C9ioX3n2YXiKG1tNbmPqUtUs7va5evKtNrOxxtQs9oasiE/
z2GRUoVjXg05cgLocdvRmXGZJByeLWhX8KPDhCfrxUgaWilhSKMj9/hbO1JxsGhO
FlAGVy4FKsjDID50Z9yP2M6Vto4dH9oWBn0cJQsD20SDQy9R6bVtybh9NAJD92Iv
79DNnMm3Od0TO9hRgEphk9R+ZxWp3Q88SZCCGqq3hPeYO35gccRueNm/JZ+6f+zG
FWNiCMf0vnJsAYNt5+UP96au7yRj9Ewm+l6Lc3/ZR9yGQlNCoq0dUlSk2e1GNgUO
9Qz30B7JzGNn6ufF9D7cQurp58uvoxSzhn4UnxbwUMcuqZYPhWIibUD9maxF9BvE
/j0G/i4wlRTadVBHU5qvrb4wEGfQeQNKYinuIwA6R3I088Ty0Az4cuNhDnPwPfA9
PKH9hHs7NPNi934zKoGsr60yp/TNncpGJLLmih1jCM24Ok0J1ZkUMo83GdZcDdHc
ACvwMs9DwKGArgJGfviYjWmf1k1mobDQY+WB0pnktd1RYFyU/cPZ0PslNHcF+WMo
1mdtpgUjkSJ39OxeJa3DAiPiOCv5rM8Xnq3zI8ffwvV3VHUdV8SOyyp3dFfWZDfr
qcmVt/0VDThjTbCtfzy4WfIYUC+QnE7zutUj7i+/SnWopS8zLR4CEih/Y5NMaPli
/SltUnxsIbC3bAeqqXI0uGrYr9TW9rxXK/Orp1xHxW0xiISmx+sGYzIBIbeNJDv8
b30tm/i3GXbqsXM7JUzB5yFz3NAejwSNEA32AgCVtlGjBwJTHQyxhz2sekyiybcq
IwnBqa1CDfRnecg5KjYUtUFTUxqFf9Q5nxD2B42s5HFkMYKly+Kc+e3C80VEjqxP
/pihMO5v5736rBrrVJo+3DSD4T6Pz3Jy9Lc++zHC6jyDDY/Bb+xMjqun58+t+dzL
z6Q0/0BRt20mLCrsF+MYcpscb+X3WoAfm7JF3bav6covCysV0RcaHXthgo2P/ctb
JwEQ+7n21Z/vzqj9842/fjIG7no/MvEPuxMrDHQBKcpEGyqY5A0Nonv0gP3gg7TN
Qb8NNn9L3nVXycFbUW2/ZmqMwI083X18SWqIBG9z2wboszN8fM9bilKsGMGlYEK8
ZfxbE++k8yw4b8BXe8pLxYHaELPjfeWz6rXoSU8AJQE+0yZk/CtVKyNJrGgh0Bht
joswo+PIgqCxbKGrz89km4Gn8s12KTUwZQWb3CY3dMHoZe8W/cRXGBYnhFF1deGV
qP/2iO2X8xYblq/uVMXDbscyvf9E4z65Bt0SpiJ3VaoJVRps/o0lEpBWJu8MCSPl
9hKFdlyz5PrqFMw+msa6X6qdJ95buWPmwP8/wYn5hinog5z4H3kixhnpRZ144EN1
kL7yYKLLnUrtvrR6U7tWy7Gq9ggfBaDi6az16yECdL4OH9hoeeYUJhk2QBbVnSHI
mI1GN6Rse8LEoJyHldT2L4NMrpI2o59mPJbb/uC4AGB02s/zFF79WDLJ1Uns1+MN
wgaees1lzsElFXYs3BpDpaNbycpjryaI7ZmtJOOIWYAtPngi8Um0nIS18XJx6yh0
aY+xzg+uRPAofho1vibqgU5P9xf0uc/2Tc8HNP9Df8tkWZcgjUBe9mL3+ArWZSZF
bXZ4G2AGdtxCFdcoWcEXFiZSJC+/zWbfnoayDSKq8zYw7FMFf4xTNjrV2WYvqlra
j1PlVUWzK1nHxeTApKPzBO8Hv9/8QFvWHFtxujSHMSqL+UrF9CE8IBsXuS5LEqk3
qwMIM/MGAaUVnKlT8rnJo0mK3sRu15b3We4fykplR7dMgCFIXfO7EyZuzmpmGvb9
YoA+QEuhcUI3fyWcxPsB+hCYo1OrM1s7kPaLyOTx81LxfF2BKX9vuPCTO22hMQl3
A2GhPOSroSidM+HMg8cqqeSWS0XDXwq6yk+sH9Um2TklXgRC/oKPqQKQiDD2IRWs
58DSjoVYf/g94Dqi0nijiuZYGKmhkifDoNOsVqrKEmMsIjp1Q/yMaoaxHXEXmDGG
tYZyxNj/v/H9TX95NDwCeLnSzrmvBNbAAO+5smwurPa9hbJCS4xERaCVHjvPXXf5
ZxqTLI1EpZPslehHLFT+8EgZkRq9xn5AqTOk1Yobh6wyWcMIy0PnYAFD1HYkV3bk
jD/KnVf+bhE4b7kgmgQo7m7jpWE8zltHxKI9uQYJ/qqbnUqyzCcugga4gvmhqxIE
YGTIlqsra8wnKWzeDJZeozJzq7rWtSKmI7x+dK6T6mCO7jEDAL4VUtkAbixsKtCb
2J/dW/Nw6SRrXUi7INV+Cqruc4SimNQV9Gv03YO3wC2ciU1eD7w8v/FEwNeB3aTk
5FfCzdn+cqsm40Czr4/l0sqLPJIKlmMVX9h04uoo3AxXUHq8Yrj+io7jNJXX2DWc
fwI8TOXkYDyPBK42c+/Hd73J1SBmSpJV6VJjV9YoAFYo2rawg8/mdYAweJUyraTC
2uHNB0pnFmH+hguLF0exZpS+n8eHUTfbpjBG5Q/xTnj00YKqmSg52iAnoqGHP+lt
l8ZJjbWu8UypIEqoG4CVNJchmqYnkJWpSbD2GDAAV66FJaUyt4M5QE/tIOfWR1ZR
Tw8ixYmIbAixhc+fWd7IHahCXIBS0YzqqsOnwny1CGshJftb3ohZF1bq/qvS5/Rf
BYIC/jyFCf1qbpIzU2VCzZwTrqSXqBVsImzLN/nD0B3hvtR83NqwjaBDDjT0nQn+
SkeehzmQd6L9+O9KyQ/4LmDux2mRzIV/DO62lW1Iz3hiZ3Vu8cd+t/6uQWVs1eWv
y61+7jfqM3ClUiOBMJjefO5GQTelckFXhCfjFoV+fjmUTYOdFsSHJDS2RqV6XzRD
nLqZNtcJY/gFUcyVflieaSrJPi2TrOmXS+1ehJog1MI6xaiQv99MPtT6u1iDsvSZ
o2Wa5BR35ERtm8lQFToOulEUUAKnoJYg45WnShNp3Sw7UkOpV28gsLYPkVMDmofm
oAq/8m1vafMCFf6q4ldVOmJVjPNLLnyj8eSMRqK3X1sV2NLVCH7wObILYn5Mz/er
Ckl2Bm03UvsUK52Mnuv8Sy/gyP0kF8qugCFLylZ1zF3I5t+j12VSu4/IG9sfgnF9
u/cXTpOTtg+NyZmrhUtby8xqdni1sCuWZ74Tv/rrWxcmSjKRIH91a7x7/OcnMzaz
OjUHrgixBIGZh5QoWXOnYrp6cusUheZpFXGsqR3j51fuR6uvECBUBL/QI+ZDvNAp
nUm5W3+ewY7JjKbp2MTKmJDeUB/LFep6q/LsQbYJgMFFXpJ/UFnRX3G1JmNjuV63
SVMLFwn7ULCJQPv/rrJUJKZ4qv7Oz33SzecWljoiyXOizK0GnS13azVkJWhV8iKG
jeELZuQ9/I1k9ACFKphT6/alajuxEYs7SS/9jLp7hEzaV073TPw4NEsdkd0uGg5N
aUWL+FtI4SSzrecEoEiiCGzqjIrpRdmhcu3LolDR3Wj4HffPjvHFbsSD6KUBa79y
wzCDyrcOz5RhEzI0ZZei7GsnYQz6ATQf3crBUDMH3XVRx/bqKrxy6pJqQQeIMLMj
k3g7gV5sgbuZIxAoVeWxG5j9T9zqq7Cw59SzOs9QEZcIxTM1nEejm3jIpuWwKJcm
D26sijj/IIJiB/NBgmdXWnma3Ss2HGFxbHtEUlrKEz1r4XoJENyIl5B5tqttwJ6q
xD5EPwePzt3fORiIMcGtogZC0bc9h5kmSbkGb/MD9D0A2NEAKAdTGdF2cl/5a/G+
l+UhydIsJXP4V6y0UTfWkfjAwHWIyLeHSROV7YpoXUuEP/0dWZJb3JusY2Q9dKlw
p67KZ3liML5Pea2Gb+v/ck9EduhZjnuciel3M5bZ9kPJTAQ+P0wCWpSKG18eGrlc
HZNYyRrSNjhfPGbrfzTpyaDGP5AuClhxz1O5YbNdYoSRGTi30Z27pxshNZ34J1wk
cWfd7aBWZFhDux1kAMskmIa3+cv/k+e2to3lDKukKcICI7A2XJJnxzHNHDaFffy0
uwEgmDeL9qKdnPM/vYVXPb5UYaNo0w/IxbsiTacaENhwTFs14vVnROk1OXHV0Vwb
y2Yy2usD3NkpkewUdhqZTZL26dD45JTeBDBiVBe8+/drrmXQIJGxCNYGFW7tlbgN
2ZalrLtUP2gCHT62EpUFYlacDHndABul9qF87b79VNum7ap2fZdI875AEblU9oMB
c62TzLf99Bdt6yB/lp7giUxxHMNoxpt31mBeBnioDc2Ujysy7cLHQnvIQXEXZOBQ
bUifQWJzKjPJjKMO3cK5Fb+SxRRHTfZVcIWotGZKYoldWI3xPVwmhjQb0yMznorS
Iw0nrnGT47zbWPQYnW7D/Bw7lDa2paLlunj6XhFZLMKZH4nYu5fz+nR13GnAdyjF
lW1Cm5l7BPHyBwr9oQVYxwDiYQ1PUkyqG+4cT0ISBrnN93oSwFt5yhQYC1QKILiJ
F+sn6ihtybupCCWgWQ6EoQ0v7o4Q14P9zI8xua3oIS+Op9t86vCSM3gb0X4fsrY7
rmWSNhPxyqZBDMXWRwfKBSSJtuOFfn/Wila4/4U8HoiCUViViPuz4cc1PB5ZFDii
UEiDDRvmvLAvmYqz0lP4NZVlYOY338gSRCn9x5zvDavJEdxjFLhIcm1SwNI6Cmc6
U8C67yY6Tm4ALc6bcT1nHZYyi2WEmhDvfZ5ZhHe7jXt/MpSYDcFpa/AXFAG+/r+j
Hpw6QB6baxJvQKHcwMelwzAr6frhE6epoYlnUReajNJ2aD94Tz5c05C744s1gpyA
RlJhbzJ07MoqFg/tA9EcvdqEkP6O4MfUOL9FVPa73oq0BC0K+Fz+9QaeBa4l2YE0
8qNwk/aqEU7cGkTcG+sn0rVx8BtACyASl4Vudc2lP8/Lr2Gl4fgK7qwFbazp/ifD
2XEcTUWv6YwM5Z/fbKbff2ixM631wqgbUdFt46fIjZaKSNefDiGe3S9VLLTpdvw+
DWSWwhq6WB08qX2iVHhHVoskp1c8zmvv/L641zAKDaEpqjxUULC6iQeM4lsDK4hM
B1dC08yffDgfl4xXq9y+BU6PlgIgEMFixowjjI2zbsy6cOAjIUrKwU2uWVgIgDGr
wNaqXOIJjxkBvX7kZe7OQSZLeDhpH4TFQSMs9RJXKG+iKHykF1QWZyDLaRpYlRKW
Sl/qePXUtABouLYQC39Ym0LwwesPMhTps6mpnoKP4p04ztYENhZRCPHvdfvTEOQ1
ZcePMkxfiw+AWl8Q5PB8ualicJQdThF1qyLKfOdC/zA/YrkkOrtdYhMklzuePh9C
wu+AQIG+ULN/ayhkxcHLYiJMKpB3Vx7w7dbitG/S3roM79DEGXTzqeGeCvgsVxgd
kdrhu/86F66GucqBA5ixSPx/xHUxys3qu+16g0VXXFlTdDX3J3B4PM+1YqLtWdO6
HT4xIth/ivbx4WDITtEHCBKrzh5HR76j7iC3ZE2NS/JoQqZs65+U8dquKWiyDKTn
Ct0mPn8pHoTPfisZqhkGWqjhJM/rEpHwLRl3nOA5hskwGCLCph21miGjxNM+VsRJ
xASZbh4eS6NZBWW2EUY0s/7NWBPCLdzrtllwClM70ucl8YFMdFhmXkuZa9jc3fek
VYmoBIGE8tK+1QYVEA0T2qon1PABhL6WaKi5d2yiNUnjpaQwVb54ccnVuLYS4R6W
FY8/23fB+ydy50jzi75JuxChtK0CGmSJ8CSkysJWECJS8qYKwlYbacjJOzKYvEbK
1fR+/mVzPhXB0ffRgcJ0fSUnods1o8xci2nwdlLlQdZMotVmEsWSmswEcOmIyZfJ
RFbsGH/I7FtVeRUExLPJoWyDL3c9bID1iVROzTmml/VmnmW8mG27diPY03M0wcTv
g0XkZSpwPAwS9NcKaSGYfcm1doV2rtF7R72JWaGeqv9H1yoaRFEe22iNpXL6bdg3
HA5dVbdLO3w2vvdICSnACzo8lMoka3w6rWRSZVw/m18fLVp4X9IHHNjlP4bAyuNP
JfDNrBGphLLensfz6G83zBP1Knv3y33ol2fZCC6oiSh7E2dNdd6AvxQ2wr1fRda0
/c2gaGSix8a3F2M16B2J+5kLFO1/qlJssA+BBpIejhhTxJWNpEIW/C48+R3mWG3j
kHgAMKE01+YZyJK1PYpCjdOV+KCHuXwukGL+xh7DHgMQNv/qoseG8Z9bhUoGHA+A
iFs6RpgV6+ju4Ky0R2eaCKpFaVP5bgzk2v/O55fZmgJhWzJHOzBvLfzHbSGhUGSG
7xTUKzHWwt78dU8Xa5mTL90sRWZfCuXtVvT5xRknWRuQ16QDaC051B9PEpLgM483
YwlYJCpi/AcmLctH50q4nt7lbZV1VGSxketyMMGHFxlPH7oHy8l+Ts/N7nqiGT1P
VWrizHWWtwMo14rlDTg9cesQsykGh/LZVPMbHVf0fPBwFrxdC5O2MxInRm0bckyr
F7yJ2wcYGMBSc1pTTNDSFOHFTaFGsefs6tcnHkKW7rb2dEDtG73p7dokaHqR+yIk
chbg9PXcrA6JYmKKdJRZT/2ZQWQ2jd9W9z9sEpMEuIVaYbGf9RdjztBWvcmq6D5a
/Cnd0N6uHT+PKEIifiSJV0D1JvyoksZtlDcKGmoxtmDsV4lfYnSpBUECgHC5cCZF
Af9o2CEEicQCE+/vU3Q2Bg6Gjr3IwbNPpdY6RAWCcCavVr1Qa4TTSAITHoOyy6FO
4KNffkK1v189EE7Cjsrtoqi/Qq12Rzx2TYEdYD7675/iTV4RZCgEgc7TnmZKWJlO
BHCwRsHtEPRVW5edQtT/67/QT59rAXZuq7KDEYUDOgFCr71455jP00yqGqmCBBGw
L/fPfdKqkV16lKxcI40P1HRNCLx0+T3ssaFNB0N0lkS0piYVYaZasS9HyOOaqsYJ
SmU4VaYrwGwyEnIkHic7iJzh1Fuijt1Du7oyISWklilUBr+X4cXcD2vX4VNi8qfR
GmYbyCJwwMvJCRrckN68PIL8vhikwqjBkY7xUmeOxoiko9QiRcFFuuO6cafY4I0A
HEu3Tta2W5jcFYi/w2fyno08uoVHcxCkYUMADu/E//yO7HGQ2ojAfQSJw/6Ol58h
CYQ6OvwQ2za1yvw0rsQHk+drqd2LMVOkbA5cC6AMjMBxrAuGyg8Pa62oNmUFTe6G
b1TksS2rBKNPbso5/hfI+hzEmYOVoaku86bbuSn+jz3hD+Q083zO7hUG623MyVDv
ZEfC+ai8SEcSg73kisBvADTgSrEqPQZMrB4LmzXwRrBPwXO5005EapDL2ixjdK0i
e9ssYmVss/8ZUYhBLkkcMSOMhTr4B0cFxjMtyin0c8ECAt4Oxd0D3UEJwQixOuHz
x3HigWOTKn/lZ/9lagKdETnfKztryzdtop6GUuSkV8LRXxcIcU17oq/VOTYuQ5gR
mCXcsX8MQk1jR1PpWNbFNY2xiyCs+2gQQRZq2rl/5vCFhDwQbASxf/jPFPNaYsLK
7uvJueldyMOFRSNuBhyEzjNDlMqKcN/+RkkxHsU/Zd8rKz/HK0kwgw3dxMfAeBKP
1eex52EqW2Dw8nwF0N70wRH488LdT1+q9d6yz9SAILAt65vV1KH9rehoBSyQUyP8
3hvPpdvONOW/zVdJsFCpkSsC2pezwbF/ffj013jkA7Ru753NzfdGdx57dq9h+Muc
FN9+D2UtsIHLKpnO8DoPo7mQEzCMS6TQuY+FvI60yYNpL6mCKIvZoqHAfVVbZR/P
kav7d6G06Hamfk8ik7ZFzXSlvNGnUgyU5EjysBNhxuSeOoItbshpXaGng3kqBZJv
TaoZh+PHwL/FRlDTpRx01XHbZEJiFk5/CzxaTxviXd0lKt5+yHAaIIy/uYwyAAGZ
BaHku8Y+C6bgYGOUsM5nw/FxPv7+Ka05WaUBTqUrOdj8N+WE6xIhOpIQ+JZ6M6jB
SsTbi8J9tLQg90+oM5owm3HoUMHe5GVMK2t566h1EYlyP+nj4c+eh4R912Q00qXk
aX3tmmIXnn9DOE55qjVBuxNaJ5GAEwmdNs1X6ZaI7DzrDmZnj63gl8inGupJdhkM
TXZHZnKGiQOwcDXU9V5WmZiiVFwd+F0ytjue2k4OulWiLgWhvIbh0CChqYxM8/lk
WDuUtOCAMRBwV0IpceyZUeer+kmdz3AgXb3gMW3co1Wk9oG29f7/bQ8MixDEd25w
4KDcWSkxYiU8WkBlipEccHbNuiKp3C2lmnugiRI9nyFBqQWY+HE+mwqSue1AVpU5
P8eEOV1Xxzs685xSAdsoAyWVENCHnmnY6t42X78OYO2BFn0lii7r8risfaBZGSdb
VYis0JAZ00y5pUOCYGGMlPA/jUxrs/EBOypW4KdA9dZz3awo7ZSWEG74vsYXnuJN
6DmCVVKYFdZcH5Qqf7aTTmzFDuNHt45QTn/5jMsQvDklOnr9dz6kI6gq1qWNbaX2
4bSPnc3MRwX9GgMBLLEtLyuWLt7YdfBxATaNkTmPokLpy5Ac1J6pfw6dCuUgJfra
Jw6RpMSYKlyuhRAl7lTtzGt2c967qfgqBUOMqvsvXmWJPW1Z2u305a9OTwQM1Q48
wZiFqRTwoIm8AkqcuqXQiuJgDv2tfz6gt/E07g8/FVGCi5RYM2G0nEwh+JzIfbT3
4lf9l+XqP3WilqK5x5lJMbuX+HlckIURg0hAF7qaZkiyykTfLvfXfa5z8z0ZSHO7
X7k2svnp5OmeiYj6axc94IzWsCMv3b+h/qHaNVSjaPssUyJxzb9eOkHpGtSvGICw
yeTgRq4OOiojX3IZvlYzCB+cHfQW//f7DVsh9ivVnrLop2l6RaRFPoBwCMUHPYAt
xX8ooNt6ecpNyyH0OjG2bMIfwuKBKw5RQHEhkDbPhYAYnED+6rUoU4AvgaIZPgHK
lfvCauHJi9z9f++rNWXwQQBPK4gcaurNyOCT8RN2cGHQ4np34FAdUTZkvOW7qjZS
Dz2dF+xuDvGi4IFJgU04R5BlEgA3fp46o6gyGtVOsvecR7NoRVmiMv7ZlaE0meCV
XKnQHUj3elhLDYQzQOjowYXDSEDoBzvwobMfpAWh9sivwsFclZNfp4Uw1NiXCSC+
DJDHS5HyGppckG/v6RrLM93DqZpU+SA2meQEIMIkOxeM23s9Y+lKE0eIGmkglPOO
cLo8yRaitdp2Kszrh47ZrPR+qpVdGUDzd4+Dy9ZUx2PrmpMlEPpbi1sH84ZkOSur
EeUaTejjDtT7SY8bXij8q6ZV9i71qxlPDa6eBco8Ux/N+cPs5X89W04beSHE1t37
9+W+s8nN4wxTihGjycBuoHs74PqPraG3FdOE5VlFkqJXKh82pCKkJ0IqbBof+lQy
pFB4CpKJvBq9f9RtaKeWc5iSGVtbIjK14YGg/AFHYr43gxfKlpDVLcVsYGMq8r54
vIy70rCZ7581iuol0EnCPyjc3ZeGxkDo+KwCRc1/x5eYzdrxGYbfM2sCi1kq79xD
bRQMn1B0ao4QIUghfGJkq8Xy8HDTtAT0nZL0D94zDVi0LtQIDyuRDjeSZpBauNVg
4eV3BGQT4RQckVX/dg2nfnoRa7Vvu6SRESXlNjGkbCGFkrkkUbvFY5HBMEsF4U+W
1xykNHfmsRAPJ0LmEfwwXBNQ1yrXwJuwSn213cedOGwtCecUowaQjSA9iGGUFGG/
bMYsH+mYw/WInr6MFVEbEtFisXwK5Q1MZxqPiXug2rxUHeBPyaX0zS4f/o7B46In
JYi73EL+oq7xlLp4MsZLRBBG6RvcYVv3l0gp2MQPVamW2ZZcZpRjvYoaSSu2OO9K
DzHsHgNNeUx2dek/RARjy7W2anlIxJ1X3DkEbFfnwhVN27+vM8rDw9gWxrBBm4IY
kMZMwAbdpXiDpcTecmEySNlC+icckBgH3CTRSAUlHok+3ynjgXrdH9pp82d9V6Hv
rhzbN6X0Edvoukdg2aLHc+Tqt1PHooUbRqroogxUxF/lJUwok4YkvExpx0dVVuSr
S1pXxluH+EOb1pHexylA+pRh7btwh60QLyizIB3d7MZqrZMi7jS6qRxuDqxPlr23
hms9fFnc3/+GefuV/2r3frCq2cO5XSbVh8hbpXvfhDFEYWs7UR0SMTGoY3FKoN1S
RI3QML7oofkG59xMPTFGgQM/weOuy2kVSQFdbavmUCRcSiHdL51chbawrRfrF8QC
QdfmwR3XAKf5Pg1bIB56qQDRyeSr31jlUyN5RsBZVUBkC8viWrRM4uWYzMOEjDE8
f9V02X/8085v0VoQ+wOc47FF6gEBMnSQlddVsfHHzIM04wI1zmdfK/vWXeGK/YhK
IXVTBP2PErTN6M/niuazN4t9QKr2C/WEc7dHRMrWLh6k6RyLJyb0SO7ZhHO7fvIr
9n7iszeHZxtrMzHIDaDyWaCr/YGck5iC1372aFWVqsSLn05t5eHep6+0za8H9FQ7
+5WK7bUjMMPUVXVvqJKWt5aTRuKeLb4oIQikrT7A40kIb+7ZP6iRlRHpyBj98gGY
XsqbIqGbMNBOczuofWcdUpQzqTzm5KRzNAfAb+1gPOdTQYdFDJMoWGRS9HlP/NZU
MpBqMwV0rm94hqLVhvbUCmXlonOBPX9A2shcIywhgWVQ5zy8KAmsZvtbah3OhVdQ
09O4y3/3bM32fmvDq019nsNdRczRk0lfj7JiOvBAn4KSlNz3S3GO6CcDS+QllPNd
a6WgO6olMw7SL5Qc9+4svFeV7gvO1m8fMUFhnHDOTVDixuQ2+oAPypqDWC0bd/G3
1X+mQVZju0fml8Cph+7cbvskz2jv34Rqw98biOSS48ju0cit5ythRESXzTBb29Bj
NZV/g0sQrvJZjHlilqKHpcuYYTquMmLjybswJxAVzbNjXKBl5+yLT8tZ5EBM3urk
wm9y0AGdouSeKeqq5+n8UC7VGtRbUaOfaHtaFepD4Hr6M0ck/u7AOccRRHa6iIYU
VSRKJa7DDe7z6gkoa1CeTvzP2v3HN6nVuq4ttRFzpX09lcjzXlUGUfwMzb9akb9C
JFOpUnEgX/ufBDZWEbfVVic5mwlMavsI6ki48YYrL8YXfb/gXsQJ6Nt2hAgx0ReJ
2lD5FgenTSx9ppFKLT58RvHxtV39YPZBvf7bcxjctA3xKz2h6FVtAGA/MtBuXJRH
ZmFXgQsGIG8yF2Wxh6sm3RYEquUbXRLwnLQv5aD72SpLJNdQZjpwrFyeWDgzogCl
VBmRyTSzTHO0tH6AEkik3JOisdg6Vf9yfb3lk3AOOxZDl9AxwlZu119zSvyQBHz7
8kWS9j7TkdfydX4+6TjUi4myq6GhAFDFIvVF56gSvzXKA+68DEhn/GYfQtnxtxdc
9w+jvWt9LnvYOBqJHo1gh4t6Jydr1Ziy0ICufQM0bRjD+CVnpyzXBE0bI3KT1nGo
NrcO/fYYg6TVCLjv+u+xwDYUPSc2ukPOlxOTmp0IpQgRSv8y04Cm5AolAJBAHzQ5
YRwUswQC9YNSdKGeJ7oXCgdmiloCDV6xEtMdTPVckEAmHtixqOdgcP6mBuTU+Z9w
i5xJd/77RRDJ1Zzy/gGUJcE/CLoghfZXMPAcDfgtYKKnglk0z8t1+5QR+fRTOQEC
Fn0ueTjOdSPYDnixQcwlXti0AX0lCWzCAl8n/sAgfzk512AdPeaH/qRMVBtxhWuA
cSeLYSH50Tq8btbT/IDVXP/28TLG0rgJFsFEugyigLWNH7vlyN0KxS1jUB4cl/kU
uEQD8okGTKG9d6F34fcNQXnBXB8D431T1g8a6QZ9iDCIAp3cOtMk15DfhDaYnBb/
6rsNW9+ubdevv+nyxj/Rbrk2yY0Vki9oeoBS1BiqWmpSY28lOg2meSRlo+BlvB++
hrsN/Pg6vMTJjcLywggsSlRAxoprE7K4sdAww0h6HnsaZAfZFrUn7M82siv54LyT
54LXvuz/Rfp4cKgsYPl4XuWSv2UXkZBMj9j9R0cB8wocGEL/pdD8xxUa2bS7WpVx
5uhT9Yftq8cS9yYFqZm1tB7duwVvIAxl4/6s6DEK4tUwQxKSZJ/C9C5ERjLUnLcN
KWq+8Z0pEVwR7PQtLX+jJU9OCj6rFCXyqZhy2Yr+1CaL9+HQIePJm7pu/XSnO4Xj
snv3tyMkIOPD9gQ8E/LREW9optP9tKhgveG3g6IbFj4vQULXi5mWBWqGKqk1I5PJ
DCiCmSWXEB1zXYR3cHrSw392zFg1RUH6G08OJX6nEDVtW1SCtB2bNjxKjknOyyJT
4dvbkW27AKmTkBkAn5wHp0OlGVdpdojUb4CeSfi0MSw6ASBG9HEsc4nYLrmRQG7E
9mRvB2/9hwaUD0sh99YgJL+q9oiZY5OrQWQyU4qN6Ix4B9N83svMHBy1GLs5hhVD
2rE/z3F48uIXmhSW6nTV54bl3/22xCRpSXbK4eGQOzLIFCDgtXPHenIXehUUMj1m
fvz8mHTAT0G/ywajN/urwnOPiiZJe2dTnA5eLlNjImrx6kJ8dQ0I2huM30CfrNis
4+yXcKdh8WZuuSLJfQsubyYX/vveSulGISOGWxt326ZOTezlUgCtCeeWH4V/TFl+
/fJgBdAD196Q6MeZcrQ/qHxuNjJu2AgzF2EYHzz2uaTj3fYYCkoWG2d23NbngHH2
A9tk6/qv3563L5KOdCTzQLaXIWJjC+ZYqnPbxirNTXk0d9UOIw8qDgx2c6AMBySq
quDpVRd0Ydj4IkoKAVc7vF7gP0QMR657/13er19UDHjHSTk7iVgBo1brQ4hDkgPI
iTOUs6FjGeizoH6Ba3mZLZ9J4voeGUg9XjVBsiAxLOnp3ux7z6qfIxzrpoqlspe5
zAOPN/PsmReAEzuFQDxvMkUnnp/aWGxdXIzI7XvQUtzuI1gE8V06HYzJR0sMYdX/
0/SxmiTGtvcT2XG1SZ3leZ/qg5HtedMzxOZ+7phlfwQpT6MMLVuEHoBQUdPx5MbQ
C84l6FvDaQdBzjAYF6Wd0djvT+gN2WmK7MB5+CIu06g9TR9Eo6FcELTUHs2SIJTx
zTzR+0Byd1zFZnlwyouU1j1q4PuHCQd8kiDfepPy8/zQhlTyItZCqJG1ALmxZyHl
vxW2tfMsUnFH8mF5YFfVBM84I4y70G6AjaGvC9wew0u1Pzn2vkfwxUzd0oHf+b0E
3Nga3BAK/kwn00uqkZOQa9Xnbk0tzeeor+8ys6GubN8+wsURvNSHKchuS6DwQPpD
uCxHoRC1LSxMOHCQJCI+JPEwC4fLcsVob/W7FnReLydz88IvnFdl4e5Ir9bOtVRz
2/1wzNR1bjyNOCdiyKHH/hObk3w4PAr9L3vp2JlYdHr4Hiy/qWF62pK2Adfw2r/8
m0w8rHQzwTWaGs1tINz1R89dELAVDAL0lhFQUkdhqj0cKrbZQHeK5cVgYpx+3tfw
eqIFyCi9DEpp2pitY1J0oSG/95wmRQcxyJZSsN6zdRjeZ/i7TQmTv4bIn22HcNmn
WUmhEDCl1egZPAaPkMNyRi3mPWvTPr+1dIIxGeW2gfmBzPl+dhOS7EUQ7EheGvB/
1Shd4F9ggzP+Htbib3ekA0dsEvLdFehie21oTHt7nhdv/ElB/zQGy07wAZJdmbaQ
KfzK1h5MLIPRzDyYVPJrGSNDvpmVwowNpoAhT27N4aCAgn2PIEgaJYLgv22yFX0R
846dNKCo6eEGqClkvlDOEoFrYwzczW61oqdGDP3g0tayTUDfpCatruHpjC5mXP3G
yN4O6Ms+1prTLCz2YNcm8fU05tLSmmjLbEjbodBko3ff3yil+OIdBM8mXWe613Fd
2TOGZXrDP8DD/2/tndY/w4mUAfVWh9/3sVVUEV3mJnZrsQW/TzanNQiOckU9TonM
oS1REZAEW+6AwgOZvfeXNVhfNMvz26A24serbyirI5AjGKKF6HGgeflf1gSap03Z
np7YKfhei6NWjixZOXmL6aQw5YRQZ3WEnJhAG4OFc6YYfqrPJlvAQLocxYpcPPME
q36VuNbQtze/X5jbWBYLIht4CpR0P3zfpmSVMK1h0u4g0OPJvLgYKzvKcc1GJ+2Q
sFJF+gHiQz/JJP7Yl50K8Yh6R+YHaLTBjK303hl6RVb94o2d3oSghRx1Fej7eW0x
WzCSocbTf+2UprLprqwCxssDl4bBURqrKGXgy34GJZ95Syuj2aszPAnuNckfqtzZ
lKkLfHbruvqwVmBfgjPaS1JRAu+9yYvKTTmf8z9m3IpMpkD1B9x2em+cjJMqCLR8
HM8TSDkpmAHv/WPBIGBUnKs5T4frtvJmH9o6xJAhaP+aeivQkj9xufQSt4oa8REG
k+fG+k2m2Ns73b7qRQV4/Qv65DZJwiqnPrLh1yJn5m65WNX66S3aNOwx3CWD2g2w
Gq6zRaDNQgZ1feL9R7gYv4BmBK1OPpt2oAGBGgPcK6PoEUGyrAsplrJGtJFZ2o76
QlucjhyiTPm85TMVxisZl+qYZP7zYWW2L4K+jUMRYN8prMH4ESCA1EjZyVP2MBpB
y3JOk53kOqfQbP1dJUbeqtGQlKAVW29kfxpSpd8A9+wKrXoDmsHg3dhXn0U3IgND
Z0D9vtfAeZSmaHzNBAQ/zhDvoHDBgUUdZI1czi/lUj3ney58IamW8e2OVe0P+2tD
UlgCgn7upgTkscYIvgNSC1OF9XfBWERU3zsEIC2b6CkCr34u/E5vJfNon4vigkvs
+VL0Z+xz3AjF21fbR4XkFfFLWoUtxV629lC3bkpBNdis27yzgPUVAX5hcNYGjMqo
g7Zs2As0QToIDIEKJxUA21+JSJD5FnsyBjYi6YomM7LnKBAqyh/hbnjBsKf/70Rv
/WgJw+Bp/WcCf6bmDZBMDVEVzaX/0J78Yansf/7Ez7ai/qxLZvYdCZnCVV0QFhJ2
6YCyasoFc/NqdXk44pEYUx8xQA5kVyQ7OMaWpMwD2305J8Jd4fwZsCglEMIYp1lJ
80Xv3v2WSI+aJid3G/YWb7TJKJE5b98BhcPgsKkTy9VYcp4rKTAZ0johsstjgUCE
zNhUxe+Oc/Nf6KEVaROM40W9edOiZabEC7kDkqvQerkqE7s926f0m6R+nsZTxB4Z
XRFHcV4o6UZTzwI2I4XGZwQ9N2xCfhQgD1U73nfyAGLv0ARBvhJBhk8+6VR4T0h5
dfxcT5kMxJ4JYRcqPUsgClqJhuwr3prbkUCCZR5HA1wusp+xGJmvY3DwfWVIJF/1
0RD1DapzcWRRtN+cNpRNY/8OlAKDIK994V9+El/J0+NwCi2B4XvJHzdvvOdlY77K
2Gxki0Suyw787sPPSw1kez7wyPvsa9gHXT7U/OczaI5bQBYykzQtf3cWH31TIEtH
LASi09IU3XP8Blef4kNWqNreDPCcoyd+0NCHkn5tRsXTggMumtw+Y26IC0oc4t3c
7dCxLH67LaZbekUtJcNLDYPIdme2yi6DE2q+FgQVlUnN5uRbZzr5samxEDnTEdDD
ZnFMvYSB0TFO2LolHUbaro3Ubc5VTYfF64kB2+6XR8HUsl1mNUF4IWtLm3vb41EI
th/Fwjwm/6xEWZojsNzvWH5GmxP/Ym2aUQoxPWcE8sqb+mpAcBFb4DIir4M45Woy
rPlHP/Lij5XdjcFMELXv353i6V/aMlJ6rz00YI+qzci2Zj7/Qr5dTl4+ZOuxGoeb
yvv/dJGUV5H2Rz56GLQomYdGdw3nM04tA2phQqnNfquX4423zB2lfTz6zLGenXnr
JnPTEBhJohFMATZWlfWCgb2lM1zetHErVs1fNWMkXZHwU145vL02accBTSlGU7pE
4AR34Ei3O0WuIyYSMlsarmqRKSdAO9LQWaCrrznn176VGFwHTBw6RBCTRl/fxtXU
HhxB4BSi5u6p+Zwmf5sjRljLH/QpuT7Iy69pN4tgSSzBHTn967uuig/mgdO/n6ct
nsxMWSR11CIlDK8zFJsSpMAz4w+hknXrPxnYa445buEQ7WS7oI0ndLOtQ0fPgXkg
RQEAV3ymt7/JKKIRXBr6oivj1hj6FzMskNgprt+JbIeol94C2nfOqd/bDseoR2HH
AcyeVba6UTppc87L8KmJHKJxUqy6n3iuyCo7PXBzgMPp029M+tse49Pf0w4BeEYP
4uSU1ZA4XIzKIGRFKKQv8CF08OnjycUqYXpmImYln1K09DNSckwzhXCSn+ZUOr2q
h5GrhI98a0ArijBhHP+7vqLsDzn4XcM0Z+j44XlT9cBgEKBrQMwchfhZKxtdxCe3
rBPGL2J34UWB2e7oCKv/DTl55qXsCJaK4p8EMSUnnA4Lf8TXyifKnbIO9XpkD2BP
ymY1d7rX86ykvs3Kip/gbSqV11B4KTwUznWRLB0EkBPmwNvVxMKMN0n9FSWiK+8b
ayE6B78ubIpVswwoyzCkKy90xJVEOEsPLVq6k5zm24RltrJgGiXY170K+JZVImDi
C2/kwtGsFeMpBtPYP4l7inU4D4T19jABK88z8MMkBTesZ/Jz8rWPTWA/SKjGvdxS
qkrcf6HkDR9oYJckQ7mCFRsEAnGkyxz6rDEJZiikKeQxxTpbJ3qO26sYETgBH9Ww
JxdoYUqSi+bztJ9KDuISzzQBzMzgZH3uLW+V5nlttXJzWtSldxtIUKfqIcaXEX0b
bAHQ8uzbTeaXI8v8M+YoGgAuLybQ3ByyksVPgDtkHJs8ywVNR1dwdcKNI4FysmP+
+9C23FUezEhPnC9gltaB1PvmCbpt/+iaZzYQOVTRBd167viqh9KPSHub8GgJxi3Z
wK6QsD05ieI/QowzoyU+0O2rNkwes4HDCcmIl5EGuqnN5p/O0AazRwwhTgDfspsI
NJ/+TdgeoN5GBNQJp4Bfglji/UyU/lGykqumfdSZZ9gvyUmQRB7r77KO3zpazYnh
yobcnibsBkaao+xF2vFhGh8fkIXQjzq6ppL5UFLzUOqZ13jcOWdeL1NSFuQvCfG1
uIKC5OHKofr8vBhkWAJMkdKPBI8p7RgUsRMi5ANX7okV8SYtqtNjgj9HvR/PxOJW
vV7+OJClFm9Qyx19b0+0t4FGJlGhBWyEAx44NF85MWBpxvHXYBJ/8CabaBokdG4f
cyezNdSXzsaeqbxdpo16aoU/UtLL6AZ562wLgyFuimL+IwWOc9C8wvqrRH5s9hpJ
MX8Tmb16Yt/DpRpR2A8EbcY+TXGIy4fGiDgCEpTe3j4WzoQa8rlAuAtl/Xlm4ixZ
WLqXFvd3i8abNETv70JTwkCVbe9nviq9lu7rU+p3z/jh2kwy75vS5fgFBglCYSy4
S9MTkhgAlehm99INd/Kd/RIcv08psML+2I9HNGmupfWmqDjZRepzZz8EDA6sQJpa
O8V2Nn5DhIwCFAjikgyewlkpe0IlQccvxNAT9iPZdelE027P5NdJ3w4rhQnkBKQ6
4hEVde3j6NbiIDS2jk9i9ciomLTatBcDgfTZJR1JPLjZyIwfgaqdW6jinReItpEO
HfRDvU91kDm5xDMQ3E0hZi8kVxb5T2dmTF6b08U5XQpIvqqiMZUv3doLSi9oZ74F
ki4F2Ie4swmTKezwkGLQutS56QTw7RVLU1QbrUCCC3mytSKmctKJXXUofvH+fMcT
EM6oBkEl9DO6Nw/xT/0iJTRX6TzKmDb4t36dhqV4QZnGZWAN5ynKpd56t/0WxhDn
AXxG4880so1Ig+TKmepBcADUajXDMTvHYjhFowKWw10zEp8PArDK4+F+7SKMaw4C
3pdj1vOdqLLtyxKjQiujbGP4qxtQXsTKXQ1Fo2km/i1slnbF5/iD05Nts1WyfDwX
OA5LjuiEGb7/wbskVIMrNRX8hLzTSOPPjFv8/hQNiWepFGoMboIQdywOvdtIfsqh
oLiP73BQH8pcGyEqnwrbN231AZ9fJCpGtJTXjoYLKrcyYDuuUv/ueQtPhRy3FNE4
4vLFGWjeaC48t67XqtxorlTLCqRvinA7QWdSvAHkm5SepEgF2H+5HHuFSrBzsVd0
PkBciuEtuQ0hTDioCBtT/UPfTRpKn759VFDkya0gy6qNMVQRGlmGifdiYZeToJI8
hL6567A8OfhgPqLC6J7IBXHslnuLbhRcPWLZvnyfjTafu091TWwsaLIRMjBUVgDq
ODJofGe4gF6OYbPRX763ae82hp72v1DKrf8CXBiCQi+XsfiGJ0L0MrdcRlLnkaCC
2gjgJyHO0k+X66G5ntXGzY2faRi+Cs+jmDi1SKr3B4B7giaqfvGO6S5rv2BffG9I
1RcaQxVNSV4MUPuM/UYCABNd4pwZGKdPM+6oN7r7r7En1aJ9us+4A7RWzfLIC7I/
0w/r8uyjxQ/5biszlLlH9d/yGvurbYIqfWRcklk+2kzKJcEUqwkkr+LbB1hkacNG
Rr/WYD/Phb+WKk5vk/9Hh+CLndJny87eoSJN3TLV+Enamd5vXuQPXOsKECXRyPXE
62HsCklmiZFXyOKzSWwRCW4KPhucL7u6BadkYnCNgdO1KzHqqUTvERoUlbYhjlHq
rVAd06wl15RQZ6lNk7sPL/6rN6ViJVB0Rx4QHZjl5EgtFxYwP0mcCK0P1TD+slFU
UsEILpQnmWkIOLOvZy5lvCttIQAiMERKhnkk1mzE2WLpJifsIRRw1JE07uMMSkCa
H7ZevSPf5KECMrkvgHir0tLZximyiR7u/L2Lg4jv+QOpFVZooDoeu7zkvOJjsHTO
vF+Eezk1Tw8YC24xZtloelNw98Tr0QRmrE1bbzjrC6g204MQ81bew6cY0gc7BZaB
tJah3k530IyJgXmxRv5LJpL5vQb0FTruFg2rE5hivYE5vhEKZXWkwcpmFujU4fnV
oXFtJa3nE5l+cGMYXVYsoR836IcQa+XePmqnyxYi9/UG/5RPDj4mFI6kO8Jo7n0/
+q71ms8JXa2ziCADfPCkC/j6GRAhvaT8QNKVZfbIPPLH8mG/VEWhNVtoq1QwF17H
j+/tTPjx5XmPdPFO1PAbL7VAE8XGj4+5DwkFMbB/asYLuwvWTsroQagsR3tszfcf
WjDArVegHd6vOk8Tsz4xx07jNVUDVQa/fCSaqyBdNaiu6kw00VRTDjkIKJ+4pS8H
993R9PAOLQ6j1oQlqVaOQE4rmFNWnmMoAqwcB2ZxCxlQn4H9ewDriFcd1Fhnjauk
UsKdFNvj3ZJnAE5q7H/rI0DcO3O53NFH/7Go+zVTWcvgcNkC6qTqE0CdMC0Se/x2
hMJ/t2D5SHXGowGhSAMZelyfRGefNH1zlub+43GAh/GLeIbOwlNPzeU+JH9gcmqf
dSG2jpClAgHUSjkYNr3KtSVPSCZd9JW8QvKNcNVYtpcprAvUiOyVnXNggV8oADS5
9QIow+/eh4OB0sWbYFFwrOztCpYJyiFPY0LFFdptE21qNNyMmb7wsAglt3e5yMFf
0RMsFPIeosh4BIEu3QebJwEtt6J/5d9Hj1HsSPa3lhM0kQALEs+4YLRr0salcvNW
fUiXsc0EZFGylnFX15zYpqYhSm4wc5ZruG9KrqxbD7DHQZw+isTgOsUPoz6zOJH9
RcT+Jz1rsAQ1mK8bjOaYjiJ1DDtdnqvsFqCNfsWjI1MSuGuoLDsm6LYk2fRz2lmY
f6UvrVVM6JhVLYyqYtQYaQ/vgGZGn1Ep2jZj/mSPP0dFHHjVKbSo6BEGRcZ7p4X/
8OoZhPzqMtOyFxVhzfTsyJw5VbyoFvfyccs1RHKdYb0JnrQ+IVzCt2Fx236Qp7gU
0GA2zsESyemTif+0XZHLPSFuL0BwEGIEZiNGZPZ1fCexFKeN5nKYo0u0wMWfFP4L
M8GO70k+cU85P6AWF1r9z3ytSS5KK5pPaPPFSuTRV+PoSsmYbx6Gaj82hCsfKJjU
UJtA2RFGSetXjDkVCv6w3G7mcRulyr7Zp+w+Tp6QGW2EJEcWOn4bGWL/8LgjegYT
08kUTDx6yvw/jVLsklX+KpMJN9Puwa6v0Xb/+9MBEXc26Rfwyn3E/TOCSgppyI4W
pvCI9vqYkXjoW9LwDDopGkA05+f4Qjz7DnhM6FpAFJp8jo9+MlpCtrV9Bn94QroA
i2WopIFs6WwDSMNXbcXcDB6Wua2ag9UvZuu32sOE4urkzEk4xbJzBzFXIM+HkJ1b
xvjOBV+0QNBxtKf/Q+oeEMW3g8PRgky9qJ7yz51SgLYO11ruO/z0sNO89X1C+Deu
ahhqrZ6HDdNU7TkicC2JTsKHFI4X/Jmo7Qfe8A3RQfhkcGbjn4kitimcnXKsXeZO
92b0c4pPJTlHAeMMS4rEYH1WO8P5JCaM1BygMC47AFLBl/VfYZuRT9L022UqfPGC
DoY2ZvkD5AMA8eBnqpmdS1MFhTYhztdvVP8fAvjJ0bXogJ7TmxuWNJNX/3Uqzk/p
WrYreJ0bwaiZ/9nGNvQqYda6Le13Ah9UdwRGgyOwf+hNVUuhog4QR8W9HqgWGhrM
m1U0dc/wnA9hKIOd9QWqvtwr4TqVokDrXDuRnBfykTc16Xv9PttiQ2M+r+hpIj5z
wxZUGAXouUUjZDbyiE1df+zPYynwyJDLg7P5yaGGuOu5PjuuPAXV6lMOdFhteU+O
T8Aay/ouwGzRsuijZL7WLsB0zLiTj8VO7uuV32NSw8dSzOO5ua42iA0AWwXFgs5H
Ik6B4olvGytWnawIN7edKBlsRHe2iKI05NJSJNArFsZupQofgTw9LoXl+Dfm0Bfe
4FclxqarOQWM0u7nRYV1OAoWF4gCyC5LGFFmExrcncYXlIr1Arwwy9y6Cw+TA80Q
p8DKsvJnd/SneLSpVPY5f/yztqrfqyuG3TMl4JjFnZrjX05Jm880wNNSInWN3/zA
srjrSgp6WfHZtE8+ALZfgJ7FQK5JyKvIkDsPq4s4w6epOIcerkI9cOSVFvv+JTIY
EC3UGzlSAWcYWphhv0WLIIE6ROoA/Q5BakrDmwgYXMUcJO09sV+DyCog5HhMsLKT
iHopNJo3mWSi0UTTiNEHuCxOS8wdBijWwUvMUyoxnr3pO0PQTY3gXFb0a5IXgKR0
Mg09UVGxDit1CGegyUmj1CsgDP8F9RQXGVqBTq1u44xxCFlX9Reyp+OwH5FMwV4x
Gk4PQ12+pFlgOElb4l05JeMqH9Pdu4nHJDgugG6iYUJyqTQUER7kIdbhhps/Ntr8
tu0jfFX6FPAxfMUcGQA2j8CXgtuofVz5Vjmbrj3hSItk9uLSlDDNF3sAVMRMMrFH
Dh6cc0cLT0pLP/COKsIP6FNXwpSlTbMysTcuZxiKNqU3aoil5gQXmz1tFSTicF/a
E17sIKV88GDHkTdVLKU1bpL1raxl+LDNdfPvyxvekBCV9+IRqVorR5LzmfwQ/2WS
1BMAUcYjIVN+2kw8rIuVC9gVkz7MZvZ/v82D6AMCV94SkU718MprRiuL1SWX53Z7
wcGLapQz8gp7jD0OFC1y2MsczC6gqrMe85Z7BIrDJ6uczsE1BuTUc7HxSG+H/J13
X0PX8qc9XD+VgHNO5FVShbYhYc5SrfKHXuwlE/Evl/EqEhj5aCMFo3KIjdov56g4
9tsOzPVRTjDN70lt1Hvq8fduL4pUPpbKaiyIOB2KSpqJZUhyJmww00peiYGQacGU
OsAVpXat8X3u9xW/fZ/MHwydw9a8eT2yyGmwtdb4S6AppLoGnjUY3mQNbmM8ltrR
FRQwxXvWqNL+g1ff8SHumO8ICihHvH3XwNkN3EkEsThuzvlMJFk6s8IaKt3pxfSf
+jonfe/QqzrfCwpr9IZQJHGzqDHweDOrcOkRAkbWOZwS/MFlmD70hKoRWi4zzzhL
xvSzvnFMqnCtKi6TK1j9YPaMF4Ll1gbhlPySxtnFXxLxW4Y/n0HOiaie/kDBZVRg
Hyv/6b44x9RRq6O33GYPU7sV/fyNSsP/XzQCmTcI9fgOVUoaqCuG2GvfqclySPeX
vXgiCae6G8KqBFdwh0ogLRtEnG+CRYvY7ruAILcwB9ZHTWPA1N2Utsga0zP4Q9LT
G/hkBj/HLmx/zfvP/UhAxaopieFXQLwzansDNIXtnN0unAyyRDGnh5BunWYH5Mv2
/Aczzed5/+6RANTgYw+kgdi2id0aOtoddmQ+CYp06hiwJtY1gYu3yHVWMk04/nfR
TsZnbrSYVT9g6tT3RxxmqTOG4kyS0J8vuEattYZ6QaqTSC1RXtUHhITHKx+e+/uE
cmJRKTbhTOqD4FRECk//RBQQ58EyZEzbHfEDonXiGHNd7dWLjMbOn//zMYdkfipD
KmoLyvwn5eu2EqRF2QGaxCeQNZDeXUUzqg2MDjlXpvikQlVK3PKcGxJsQ3Me5IxJ
PLkxxFycB7h9LeYeGNasTz3dY/3YonBg64oLfA94lU3Icpr+W+5jyaz+IV7lpcVG
LzYRXvLclB/P0Tn6lu1wVCC3GEJ1xhn0tOomgVxLCKf9h5UAgRFprm8gViGMNYG7
4u0/AZ8dwvsZlBWJCq0YWZQi4xEL4cg5HYf9qeimAqI0+60oTbN4LNYTL2cvcSCj
YrGdpHMshUUe7AbsuOAFkp7+rf3xg8OC5wairN2tTLpWq9AWGetwWD1owBggSFkZ
koL5jrhDvO0PLMOlhbrrNE96LyKwXxV5zIqJk7b7tSFRmQRZeZUoflywp0EEDzji
LcQXX2mqL63yClKxRNEkaS7xAuocISkX8Huhi6QSQ3hzmhKziTx7vru0ewv28bRE
UZi63LmkIJSu5i7rzZVYNpJp77/hG50yheUpbv7K+liUinJY6ZaO7pOulBDUZouk
tRgqngx0PpBSIFqYtZD7jkrH5JF/Ep2UEA1xpt74i9XULuPDsKO29goAHw7oKQvI
iqdrpmGBj2aDjwBZ5RWsTBi+05F9tDe6QTQUfqYRYYdxv3BtGHcmVZAjKn5SlabF
ersiJQswXbhP7uucBKuXKxqhqpmgh5FLlqM69UZcdK+EnhS8CVxDdOMFAO2PhW6s
TTET002KRIOWgTT6/n1W/MNEHSWXvKdTQP9s4zIJlxQ+xWZaLgiR+dEICOkikBg0
pe4x50Fa6omAVLnVRZ8bjQ2Boo29JvpVBPhIRJdUIEnhTPQ5KR1ztw6X3ZCFt6AX
0qQG77Mw5wMpTdK9KUTXMgwU+hUQPRgzCQ09kg9CfLFaFub///T7RR+Dc/91I7Lw
KsySRHb/bFBYEebCdrjE5qp4cj9d1b9zwuYhUgFI/8aQdSTXVIj/drWS9bNt+emc
gVgsnTdS5oGuDy3l5WT8dYZi8wZvUcQXWA634yz/kbLN/ebDiDJ21HkeKS5UCv0S
4eXF9UnZPK31IdipnNfPiSxQi4jG3B+HPYDNmaH9STYAqltOX6aKZgRAFEP77I8E
Wc7EVUZWNcL9KEUOd/IKyZo8qx1jISDomdzsMKkmN4T9DAJnh4l5rtZHpbRQDRD4
0IhjgCe41v5gGC21NBIxAenD1trkbwU5xwj6+75roHqq7DfDOhpvP/zft0qYa5g7
q9wmJ4Q/wPqa8vXJjvZvbHm88BfgF1YXxc9o8rXlblG6+5AMoz3Zk6+7GGbVTPVW
tKHraqKEhAy2pNMd4dMVrYTKxEN4ZaycGvE3vzHGF8XJMcG0AQxR4LxEi+Mkpjj5
5xWZ9Pkkf6FZpq99w072LQDviXn8R70KO7PO45tHnnPr1F4rbbjJYoO/nHyJkXac
+CObZcTT7Sukq3NjN9N7PDjT2gBmu2++Uti033wlvXT9UW57LUXBeBVfOQGL2lq5
1YUeV75SGvzccO6h98KtXbpHdUpS4mzCrM3UqABqHbSfdkypaF+OmzryM0jVmcev
ZMqFHDj4UQFb+2VtQa0WRhF1jABS56ujHeCTTGPnVqknvUqgeBtLmc5yV83n8hQ8
pEszj+KMzY8CiXbKE/4Hw3v8pomkbWIzAFswY31YUaYoJNgsVDJO3TNNWHEPmszT
sTMVI+ML9A4Urrv3uH4J1Aw1571Kt2TFZaxHAMALIwQJpZ2W8inwSj0aC5CpoIi/
okcJG8taRUpJ/BlnkkfOmQ7a+CjQ9LHYx71LB0tzzE47jKNQ7wJDeZSnVcrRmcSF
PmwP6rc7Fal1NouJlE9imTQ393+VtwtkwKDwBAUCNJqwoCGR676x3H/LSU3O6TZw
i8ze/bLrcmYzd7oc59f7F/g9JeJY60Q2VvHCc7BTeGwpw0RgSdQ7CB5vxsbLdQiZ
+WsiMBkugiQfhVmRMtOP/cCAprZZ/y71gvkuEa1748pd3o3IJTr/+beSweOkaoJb
et7dy6AiEfSqMKGz1HM93ej0M2UpsE84SrLLZmoDlIF38dOUO4V4HPzNSBKCQIZU
XrgvCR++7QcuPx6kri9pPKOzyMtis3grrWdVvXcIiWoLt7LXOPXZA+kr/XxG+m61
24PYeTG2xnAGX4WhsyTb22o1VIah5eG5wiIVM3Pyx6LhnJyZWTfu/Ex6E6iKGBBq
cW1MoFWFiN0QyqCfl5DUlkFmDLO83YsRVSQoM8c1szpv9MSjpEsnzEsH1LWzXYbt
PZIgdY0tLx/IE6IOKxGJOOTNb9UxcxRkMP/QzhMk7kaMKw10wH254JKj/EzrgJ/Q
0w2Z313MPb7U4gVQ8vwgWfqWtduCQ6PIQ1KsbbfBYOJi59u8rRPJu1Y/L6QudDjq
ZWDEnxbRpTmsZC4xdlYrMm+eSwD0iiRcFqYpDosewzwxA7uUZ0Tdu80dIa+JlErq
pyvZQuF88uTV0yKH5nIjGr0lZSHY9e3ZeZRkAwpeXY0h+7bQ0HJGh3vw0garWnX0
wo/ri8qWsiIO2SdljrnFONUwS6hIaQ5y598BI5fR2/mW/MJyj47eGdb7zrg2UlkZ
x/OEOxHt+MUFdaC6umxyAji0QsVhKpcW2ZEiAot7RNokIMgxruDM5yPn4xT7UdzQ
UShQFRzLq1ngDSRwqxDKYiVfHikj7tqBzXq1tG3xMomVlqJdI/fRHleEVR97KsOU
lzBokJ02GJYCKoK6sWJd4BKd4dhss8G59AFxx8ptl7VgTE38FyVZVh65wOhZxcCv
1jjerlIrzjRh1zADxy5TyuFoqFF3Uz5lno3TBEazqqRiKTtKYIhVW1Bz2gpje0DR
fvUoGXGuGqXu9CMOcgmhpw207e1saJoROrrQmOAUPwuVuVOc6q4nPbD34l8sJYu6
7nMOc39vigK/Mqa68YWkWKygYGUqFPBUjCVYEC7Wmsen3jdBxpb0Sw6sZI3ZdyRN
T6rK1cUi9MBtA2ZBOTD2PrTtUuarhVqfHbaa791DFanWzL999/HQytkdgqQOQiWD
JooMU6VxX+0K6iiJZ/2lCyC6txikZYXWNqpvN+ZZ2KqlRhUmKOTZJJGRyD7Tu25+
cdj0LK9HFWr2qNJ7yWmu5g==
`protect END_PROTECTED
