`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYIxMsxSgOhZf0kMQPTg87BwTxEgXGy0TqrRp7C0hNi9xKdn+zeI/wL5UPSk+n6F
Ja7Q9VUNjW7wzzstO+H5LN267p+PSXQOo9IZXxBoQSFM8Wy0kv6Fl2TEgpsuWxa/
/oebYjP3Ux+r1U5ugqSZgd1xbtrD3Cxotqzm9Gq4ThB1za3gfjZ7PxmdgSpRWR6H
nKya5rQgiQAyivVIKLaseDNoBknLVHLBZYnF4UuLBjSlv6zRUwW3a4APHk/exfto
1P0N0jqd1mYPYiSlDvE+jW0D3iGVZX3FuSD1Jx0KKVaOHBUrY5SuzybaEYfh92sK
lUxZMzT6dIFGhv22Y9ANC/42OMLm1e8A6E6ocWX8DnElLm65SbBqluqTS8nk07f4
beeAw+Ra9haA4IanFkFg3g==
`protect END_PROTECTED
