`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YvSdEBsfGXIG0GSUrQhOIHuUhwl1dxqdUT6ZnsagOMCD+Yxd2bR2bv1bp+NdqdRj
bvVqxRMfIM6uvv4ifO8V5Ynjo828Gp20zhKG/UTU2E5GldfC1mFwMWEV+UYDtZGn
GBmEI65NrsOqzktzlm2imyMVHi0DiKGKM+TeZqjX50bgeTcG0x0UQf9QC723QDh9
Py7hAfVsboIexRU8O5X93DIydoA5aidhOJw0mUuilCABVWW66bBHYt2NQBc7sur9
7W5Dgu7iFzPtC5UZfwBKwzhUGfFgQLtMscEO3i+p7URa37akynKeXdg35rPZkbgw
DQoHOBruAcU7JBTIb6CyA7X0IWhjrD+4dl5Lj8M5BVAhmq2yqluD1mk68ItbkA0i
Jf54toEUNM8/J/ozvX0ziQgA/AGZXecbgO/lEOY0wXofajZGu4V+yzJHuQOjxhot
0l9q/kBnUQuhDCVr1aT3fJ++xgqZ5g69stzB7Uv/XTmfJzttHHqeJ3EYQ2NyQB29
IMzDZh2t/p/CVV4+ld0rPD9DWL0s/7SGusOlTc+5XybowbA4HrhqniB7HNkkr+G/
pOkfhEP2IW508zyKmk/+AEUVMmtmefoEU5gBQ9lMMeV2cl54B7VNfZqv03AQnTZS
WPdnRAWIEKmNlsqr3oSquWpET5QEyKL3pvfUtOoFuzSTpFEd9L3xvjx+eTabNXeB
YtGBrHjUVEeRf0XYA/QViLWGbClTxPlTgUBT6dYNptYOstaGbRipUXI2ukcbIKgX
ssK2MKqPH24sbB6AFr+T9Jb14Dz75/wrIcfAo50c2uDh7+GZisLeL0vT4d2k8PfY
4SvRtOLy9tAyaDpHXCqe+MQ6kIkzdy34Pz4WTSXNGmLn+t91L5d8gHS4oWZTb2Jm
+DLPBvGrIw/zOVzgpRbuaSsDErnA5KBnsMpcyL7gHR4=
`protect END_PROTECTED
