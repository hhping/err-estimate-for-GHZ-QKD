`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/gHTgW2N+sWL4C1CuCkod5dZHy1Cn0XgutHXrzgACjehUGPtr2Znud2LFMQ1o1W
aPc4GcweOENVO+UalL4OTmcPleQ+bNf+hAad1ABQyUrk5Pn6iY547Hn2BrCm/eq4
zwItJOxs9RoqND4toL7OXwRBq6XpNIpChX0iXi0KcdNHM50xuh9V7PNnpDvMx9TI
cOkLSYtrbbPA+Ci9YMN27RDWoE/2vF+39dKwCSgJKuR4MvhZ1I5F8ljIdrarQopT
uJ9fY1uCMAB9ibJO7q8d5SYC/0EBKis+nH7/9m42qh/RzI4n2ys6VEhY4Eg3g+uy
JMA8DulB7o+zL3Mx3gsCL/B8QOUprB7AfZX2KyAoecjAdvqtnyF3cgr7TGFiYNxa
D9gdxMaXEp9F6kYJg86pf3IQD3bK93Mfkf/LvvmXTBA/TBfkXxseUGNRXYWSXvyR
DMWfH1WrF1ROBcLo+28ptSI/ETOIq4xO5r2wysRIQ7y2nwdPrfyW/AQgMF8irhQ7
vnbj5dVk5pcGxrnJpsbXmFRESkz8O84O+SR43hRH/aGg2wA5Oxv3atXoxKAkRHSi
IBjkBBBD1kKIIV2J9hsWjhDSPJLoGe63ru1us3uN2a+xksejRdtIHIHQh7zUfnbU
RtTsF7QyiJe060nUeMF94Zj63Am3a7ggANMukAhsgC+ojCoODIbO8WslltdCY9aC
MEZgbBFwNOf4NywlGyb3zKH3XnHISZCFfyF5VU65ht8=
`protect END_PROTECTED
