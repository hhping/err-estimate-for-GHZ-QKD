`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XYS1so/QF/0jCCWQQ9nyrH1l36CLb/ReEpEPrMrExdhUssduGaiY2xF91d04geB
7wO3NWaIe2Iq3UiQcJe6a71MARACA7yD1GX8CgidIgRA/iyxACK7TvCcDL4rgcdh
3SxDUPICJrD9A31yxYGJvl+Cw8FJKQlFFE/Eg92XqL8I1IkbSdbqXa9pdZhvEoZ6
9XkpIp9I8My9O/ciPY6qpNMlbiPQOMpLtVSK/X7ercQe79lNO947walqzHGhGnhU
oGFRmiHKxVWXuyzsRn6mwPH6q2P0tKR2o0KB52t9+1DBkodEvEmJkbAJ6lBQCXMG
YRuTLTWXmHZ2uOjLEPOBsYgrOV07erIOAiWOkpnTtHt+a/n/6s/hrDJRT/GxxRyX
uR2nWreLBwWvpNu54bH1TYvMAzqYgSBkRFe0Ypx58Xzx4JFDQKftwxei4BL7+WD7
BHSSFuk1MqD8eW9fhFrA3RxvRFqIjuQbzJeFeoG67UAA62lhA9cPHOcVLKY6kY+b
rcVrppXHkd2GceaKsu9Z0NjfjXm+qAOHdcYHZgGwexmnDW/M7GbhCIVsI3luRKHj
MYPjq6creg8/2BZOulalNWh1AEiiOi38iiUPDWjWng1QTmIOhwbxHbI6cldfBHbh
69Jj1SkY9Z7Hns5i4noOmQPWEmaCFD1/jKBCaLWp3nzAHWQb+6XNLbNU1L5JL3UP
j1MSul62VkVWyLclv2Ax2NbCyxt88Q1xv+fSJVSXtJLZFq662r2p61Oe88ql6RRe
rJKCtE/j5ECg65tuAmtS2HHvjseSWGaScFCQCdFxDUaj4iyM9W8kZSNXhqLvMEmD
rlKzTab6p8YXApOi5t+MWKHWr4AS6c4H4gOP333Ybr6+U35P7Q9a212qOsytbIwN
0Iq8QjD5SR+VsvTQSYj91LmxQdCm1HKz+yLwnUAICNCzWkVZVnjxuvYW/oVZLxXO
3iefjHLDP3zPOuHILO/ddUh6baghgtH8XyK9bV9E/a2m0vk3TdgVSK2KCsDeUhQr
`protect END_PROTECTED
