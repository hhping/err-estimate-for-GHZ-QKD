`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K80Xn4Ps27PdMoJxpvxtKvE7gvNuxD6LONVPAyAH0goCiB7Xajw1MSmwoQdriIvF
vA7UBSaEvZk9zGDpwJ1ZrK4QBwpennHThOfXv92lObm1Sm6rdHT6dG9Tk8E70Jvr
3TDNmgs1lP3cirwYf+/x8MHOT2krJRbm/cGhCmSa50MQWOR+adutLZcFhyqpXy7l
d+zSQKgodkh3eYwv2ZFuFdQQiOPBxJvrM4DJT/pXYd/HOUlnBykGA9YrmwdG3FeX
zwHdlttPkCaJOycLdxOpjw7CATYTWn9qMGCu7kTotNC6DrlxfYahVrVaHjb/HyIE
FDS7J/rr6HEEt7j7SdtQfhi7JcG/HvPttnKdmz6NtvsL2xq9sGpC1Q4EcOtTQrNp
og8mM1OqNumOR4nhA3qYtTA7yoLSSeQ8Cjo6T0tf4pNmyhgcCQ67Sa0KqDrlMH59
8+lDVyIqw4+zap2VaN/JSSlC/obaa0WA31r0hKxH9DaC7aTrTLXZ0A9XbWFETu8O
vHd9fkt5Gum4Yza3xhyn240SaruhQ57I0Yf8ho4pfw17yF1AxK+r52wonokvjscH
OeWVTCfusCscxOjbyfwXyxX6UW7uJ3Z7FQ756GHOPvJifYMxhjMmlXq+thVYwV6v
HrQcIDBg8I/01u+YC2cRcFTBfMZ2We32qColAd8JU8A=
`protect END_PROTECTED
