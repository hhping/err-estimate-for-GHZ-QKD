`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovpneAf8MJX4hMznyEF76IfW6N/sjCJYanbL34PhXGbJlqMW+zxs+G4j7kXg/qfq
y2g6atSXBye5f2w5RkI91JFXTjsvn+n00IS0wte5Skf7fEVGbSVn+ksHWC5pBvv1
XYDouXlh+beAv4Wlp+6LhP+bAyv/cCR/SMJ5ydgD1xn0dWTYkfn+y5LQLWyk1vCs
gS/3FWiKqthTVDqaOgBRTcAo19X3Cu+ZiFOzH3lNwI1nlg80HGnortPXGhp5hh16
vEbDQByzVdYehhf9dBa7w4JTlJSFyBkM5TufOV5KZPkPb6Q1oANdmrPBbr0JFzzW
Ndh0sPH7y09lJPEjUgA65YfYhTT+4AoEUtX1GyT3T8O6pjhMpBmHLsic9iqTwmTk
Ud9G6LHpbR0iBzSPeTeCe3gfOb81fYcs4MNXn/JKUBq1qBDH684mAicTa1GUw8x9
F62imPy3jx0Ua4eDlUCzn319SrmyGySyKV3ThnfHsL2JWyY1og0/DzIU83OxVJND
gVmJ88hKgEjoO6cpW1DDdTm4et0ik5NAdQSHEKBpOc57Zov1abjFN/vaem0fFSKg
z8Hv4Rlv4c9nr19vlMWilGgmVKU5BlYBtX64ZkNjUBKDpU43fjltgb9gq/ZtAzTg
nx95XaiH/EfpoB7smTAJ/T6wRrx6wNA2EQ3ZBFJicmkARhAGWpCLB7gGctfmfqH0
cb7MW5pJMJTJaElzXUoDj2Hk7U0gZpsD3ojWjHXqSq1QpCD/7aoVx2eJXbXJwBZH
HQ7QwJgWGtWfkxhv/Fc+fL17IACQO7zZ6DxHqxJf+/NEX3/hjLHIcPJ7u+Tz1jJ3
a1Q8Uc2fkA0bYxEapmZreF7JJywdU8S9NEj132QQglfkwTKBh2dw54QLGGLREoln
kfkNSVy+WrQIshgNia2pukr3RAUeoFOW8o4Vd7ttkb1Sg7YQb3IPAss4+5HoxWHv
yCSpodSykFvd/Y9JoI39Jhbq95BICYNx5qF3KKjQlzA2VBcdEsew2KZghnYZKSOV
V/eWIFoTvhYPDwoijMcqFa6hklBMxjPiJ1ILxoXl2bArnVZ8ZVlisdL6LyCzaK+U
`protect END_PROTECTED
