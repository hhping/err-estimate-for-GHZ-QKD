`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2d2HKvQiwoEBLjQJsNzNFQ8Ylr7nVdUQR8egL2m2zrQvTYqZ6vzqqRbCB0KDdfZS
iPSJkWMzH00bYF/FLRh+xoxmoKLtUiIRQnOvE8wVpUhtkECSNL1igGJ/dUrfn+5q
KLlv4BjxgmfSgTtOfMaatQH9TwZdQPjNsY1w8UMqxjQEM+o/w7Kamq24f9/jNM/g
rqfvqISGHKDNwFj7VR8sC+3cNJmOCqBajslQ2iHIniiUuMtImTjy/B3SBA1glFjV
YfI0XvrJ2iAL5szF3L9X9M03yEISVZ/1iIeLhjezsewUYYGnScDojjkIirh+4Z6n
ISCpyU8UqMd/bO+uHOMzIReNofO0aBiKGQQsyymMTohOt7Y5FeYFQCCii1L6PvE4
kJOMKZM5B1lZmMFrCsinujV9FGLlmu2j6N31VsjYp1XXrtch+m+7fjWVgD04HEnE
Z3xTniSQwyKvN6nfB1CQ5IbjjfyecB+OkpCGe+I4sJT+cMnQ4XXau5ZhF9npvqsM
z3CvZFNIaQmtRLcG6jfRQdF+ZGGYAcrJz2qqwsSWkQkUp26SC4j2EJt4VqfL20y+
LwMLsmmJtGUUTn7wP7sN0+MrjtlcyQvz6IbnoBNLuJQ2m94IrEDwlVCxRb9zXMrv
Axoo3y8sMj0jJa1mlMfHKG5HPDrtytA/MUd7WVpdDlWdOCT6eYWCIcPfvqhI8PyY
A8TMvUxT3kNMvpMrn8kz4njllpMwJ0mBylb+hc2zUNMOcm7QtYH2EakEQ+x8i79S
mjtDAd4KN6VibOVkUi8ceM+BqYUReoej25FLY//Q4Dmm0pjqUnjJkZjW3LNCEcNE
PtKMsu+j3E3wzGTTF4ASHAwsouHGM9qCurnkYnO6L0rhLyTyf4ksxBpI7Wo9pc30
8LLQf5t4BJXNvGLVdnIpNHvcJEX7S7RInRP1B3YS/niBHrMWflS9IcmUuMPPsyxk
VrasEtTg9N2vbR+l1/AFbVUUJ/l2zIRqJu/x33uyH+kA1GobB3L2GeU7ZJhLqTUU
Wbv1ILWYF4RuyZyar7S+lg==
`protect END_PROTECTED
