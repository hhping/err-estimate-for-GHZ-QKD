`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d0h++h/x+vnp/XysiER1pj4I+Jod3j7dPa6ISmjAxRaypi41+Fh+vhmcP8q3rtc+
zQjfpBCy65IB0D2bUM8H4Ssa3+hH3oMaS6VcS4DjHx6iX+PFk7C3JePsB/s1gK19
tJzFpRzlBSnUktdtuotjHf0rbPDJHd8yCgPTQB/4ME/znvK3lQGVNG/23TpZKxRc
+ZAOXDia7nUjNRnv/DGDH8V28aJDiapULNwLwSaTiU6xQM2qsXIl7rYanqXoRpHo
A5ipKPSf664y/4g1Ke0aPa3Wj+DLsu4Gp7uB5fldCZd5bkmOA1wKWcpECgJvELHV
t0lN0P2Et7gYKdkd/PRHOJfcx+B3baSC2YWCWo8a5FQ6SD+wun3VS5H3Hiy/IRUb
Ekrxh19w/U6vbNnnt3mm42dvFyhx29MrD4qUfn7aMVJphYHaB1LNc7CFHNy11Hc2
GAsgZVPRpiGVbYGAIhyCkUwDhueUlL9CPZfMfstFoSyG8tNcLxYB3BCEk3Z+6itO
vSxyYkaoAiA3BHgBs/dIp/tWSvxLfjxvLTvv3g/vDstLcuy6oIXfp2+yI+ayIYG4
CogrCDW94v7M4hFsUwqyMmuxWT0HncCatYZoPUC5NWn9iOi7P6/6AZiddqopmcwI
C2DdkRHl2oVcIHhh+4dXv0QzXeQG0+DEYJ3bkR7I0bkNsTHXcEtBOG68ZSyQ1Tpn
LNu56AIU7myRj247qx10IX8ZvtaCST+0sInFZOH79hFTUsxivCx8Fhn8DtMJCB0F
xRn6G7s1m1oFTMTK3sY/GTPOlZHNN8aWOsVYrM2z8NcQLrwCb8dR0C3BAZ7VPS+Q
d/5A0MuqbJ2dhy814kXjVgHQ5NecQRNwefsexC7otbu5RSInc83FUt3m9Lm7azYJ
rs4kBQ0A5akLYkUABAwZLXtXfIq+CudP6R8GrFBRihIbdg+b3+DANGMHiNUzajBd
vB0MWUBxvyuguV3MqfvKWFCDZ6UC5a/EP8Jcy6gAx9ulH4kxaezRZHAN3517LQxA
sfNsJuwa54S60f/KQmj1BT+Q8scfh8xmhv81xM9frkQ=
`protect END_PROTECTED
