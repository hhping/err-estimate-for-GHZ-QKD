`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ao4Cl3KUk6kgVm9VSxL+DzAZBTtMG2JcWL5L9YwMxH4POIZ9lMCp5riLXao63K+M
cARtUeN7tuVrKe+44bPx4QIqFPNXIevl9QckV2fntP4VHaRALgQpGcq7tXA+vW5p
kDjAZ8gqM6PoAf9eoqtIJv04PUlycfNZb3Kz5WDckhO8jVQ/zkH3nbinjksVhtaL
xPlneOw03t17QyJhXUc/w7wMuBnnLM77x3NB50CCmwjYVii1owXHqB0WsY6G5fbC
Icx7OdPXmN3h1ER8vCuw942h4YPCzpA7PTu3/gltPC1YymVJQbi9e0exd+FLEdOP
9HV4NKhWU0v/bSTZv9nNtZ4fhCUnokPzkiI8apDqSM5l9Xvnny9xpOZpUREoYZhS
wZ4rVzGEEYhzD3MmFCcJLLps/0P71bVynpwhZ7c5BDnbSiFghdOup69Pjsa2Bykr
M/Y3MsWreRls2KOhH/tQNns6ZOjVLAGbMZMrLyOqCfxMu5uXbUM0sZQ+opO3DNoJ
ZxblzRhK5VUOHsVOIRsAJ+lJWr5w42RJx5ZeXVzT/6x/inLC/LS/kQmG4ep4F4tO
5CFIn+xopOxh8TcF4Wjl724sJBq79oijI/wzEVe2mfOf0CVk0Q0hXOoHz3cVIOCY
J0XwrkfrylEzAq6Mo6SrHpkH2p1YN2Z/zAsU6UVeVRVR9/Gl11DllDEx0GOlr7ot
M6wLQ1/nLFOq9H9RvzDmsCvnGr1/10NEvcHV8D6U02g=
`protect END_PROTECTED
