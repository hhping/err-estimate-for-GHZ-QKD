`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YPF/R8gkt1vrMi0Ayt79T1X4DLYd3IZizsy3rNQc3hy7vAc7C/Sa75ZEe983EtKE
0UCVnTXWBK2HM00skMHNsHrIXN0foFtInoKcFZobJ43r7HdLeXKYaGRG3E2YeHLu
LHV83jCD9+qr6CZ5tu2QgobB0OTY3So2jMjH21hy70TF9IAKbUPdBNvyE8pTHoa3
ZdlUzwZQBZ8ExPUHPZtBq88YjdY+voe5G77XazkWJLkGbvRGKeNerdZoZalt0Qhk
cJCmnVy4jT3AugYoIaU8uc+RctG3dfV1WTH1x3t7tV4=
`protect END_PROTECTED
