`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTJzGUWzY8JtgUIZpP/eWZgBOmdG7M1CaUPclALp4AdVdB3umh+wb27ZkbvIAeEJ
m/Oj2dz0qGGGaScoK/Th2ibiIY5mUv69ekgp+LpU7alkbyZmAgl9gs+URI74Yeyg
tx6cpvcD96PhhoDW0GAxkkImdLSVlGmDXL2Sgn/k0tWfBRlUBf2PzFvdlp6Dqysr
dwIPUFQ+oJnmG1TcLDsEmYi//5YSJagS9ZGVYdvPHEk5myLuL0VjuHOy2pe18xNC
3t+LaDAZrUTfKICXn2OK43tyBZt6HWWhWdMbS4LHMpTYjgmkg+leIhNoA9RQmCP9
WODvnyOlZ+CWzBUVv2UpiNPPzL8CmqjhfCCFUlYwgImZ2rEzyAAtv6+eDzziqk7R
5Mn4Uxn37pG/ZXdhs9U7Ze+1KzQPi5iCJZb913XeaC5tsAOy/4N4o706q+hyHq+/
fLSEI6KoumTL0IevqknjLzE5f7NWBfOfqgxwoJXX7NSj/TUErzDeK369pczDAUk2
vN580/2jI9gEFzMcNv5O7e3cpzqmQ7ho5wsuwTzuKHyafHPzGs1f5EpZGeu1IqGI
EZ6udC8qp/AzJuFS16Y/tyjn7uD1XhUbndMhCBYotbpmeucSDo95i8XYzu6vyt9D
YFfyWUTlx1wM/L6JBIJbt0x0kI++LC2rkPVdY2Auo/jpaCiydQWVvr59Nep0RTKB
MOnJxN22JvYn8Obeks9PEV9V5NkEUyApGFztM8iKJY3TNQNmq6kya1yoaiAhYctb
qlk08m6heBHpXUHeIKmKPhsyUl1GVmRpwuULgsEPHX5fmYXhsLXs0CcJDuu9v9Xv
uqgfvu0yEkZNK7++TUWoEAjFxKRvwmevqrsqMc1IsACbQUiAYqAPoc3Ps09mT6e7
1NYsziqAbKH9lHOVDr2X7nw8XrH7Fdmn/YlhBV8yfEgDmtP9yHy/0XblWsOXZsZN
yvoXpcanPJnaSxkbyrycige+Ig4X84twUSwbf2xCq68iY6VvtPL4+H0ujXkWmcCg
EaIH9pniMBw1P0QKwXDoyx8HFpIvo5i+EVA+3zVh5nHluyIhmJ344emyQB6wNJxo
UGw7h+a3eCwpXicjyCnPGe0gkxscQ1EDKTonjL1hgkqf3wvls5uUFv+je4yHPuLv
vVlNp480EVJikOs8i4zj6CbzK99Bc+5AP9nGqiru9K6DtF4AqmYy6RA8Ss3X3jXG
wchWr6kepVIPreAn3jc5b28O1tfHAtEqS1GRRb5/1uQps3JMppzALneyWGzWI1MQ
y9ke6YiOWK4vROupMvckSaUfhDrlIi6cCzpkbKbzDbp6NsLfFJZWeJrN0q1Y1z0p
Wt3QU8zjMfTtGVDL/VOhe+39+kUcZYXqSSKQRkpCVrl0lzo0UAnIlb46IofgwBRk
IXIEC6cFua7IQuQHQ1RxSDemJpWtcAepIDPmwlgSvNt74yOKqZ+N45LPalbuLwxw
8nEirYMwxHmBSXcSUTBuH3ggdeP2O8DZCVqVxBAacSQcf9Pv4hLu+JE/bcybDpln
g7Tb0UEjBKnGH/qd2y2TNC6iW+QpkYn6JDqR9Hr/qnJh54roVITT13W4RY/XdmcR
gm+eE51YPfVVVkcqu7Zp76ArV3Bp33B/vTgZ3HSzrY9961P6afMDj812/rGcYx3o
bcU5LgAB9jRC26S9RmqSj8Wp0PrplXfPZiQk/j2RovHk4uKiw3uvSLN/jRyjg30T
N8gpneHFpKObyXJJeNsjg0YnmJ/MSv2q1qGhID5/dnCq02mjES+imwex/iZQvEg9
Um1HPFCujDIjcgMzlx7hoArJXz8ayuWtau5SbJ9vPI+86RnjVWs7cG6vfEN+kfRY
be6VmLIm4tAC2ZFgBYkBPnDnzBad9hP5JqFVnRY8fqn//QJhIc3eriOu81zi3K3T
wcAk6k26Q2vciZZb79Y4CqYpcV6eh9tGuX9z9keCwD2mZFHIwsAgLyPrULJ89jyT
vax0AT4uPNQvj4ZnbOntbAVoLNvrGthXbokTBaA35N/X/TOw2an0zyDTnWZEA9WK
pxntOUBXerN8A97SgJrW3aXdt2PytM+ZY6X5g1nQ/f6MjmxUx4fEGyRpqBOkQEUQ
az0ksGrdOHed0vMOh8WdchweKVIZbRVFfPFsWzFsilIyiUddnZH1RZ7X1TBMMFr9
fQjN+iJidDDvCI90oVnRmlZyDJbz9DCn/Zo4If9JZYEhBd5YZSrvM0CtMnPkPq4i
yHzzjeB6a1pYQOOOkruZ3iZ1KzD5IwX7cMH0icEfjICvoWnxyMAGVm1oB+8LrxhA
hX1axDETlqdAEdSrPphemFu8nM4i1fVVaMmm56/anZPmtACd3EEgs67SS0uIUfnv
9WxnYuKS6H/Oyy1PDF4Np4AphGlyHWj7jdmR2S1Xu0DC5N9bESTJqzccyPiGw1qd
RE3349Prdxx1wmsHQrTVOJrG3waujFq8BzhlAXHZGa4ive028d9uZtR/6U3Keapv
eON7voEj9Y8TzcMGmXXgGPn78o7rG9s0gL57kGy/OyE8A1ohgfGlHX5TcIZGkCOR
8Prez8/UaHIQGbIyzBmJEoUNCLeDhAYKkxEeC4KKMSYwi5Mw8Ac+rXsaaRxIzzrc
6khubgg7ePHv9tq8JD7FQFJ1WrHZneJQIEiuiapMl4oo86IF8zDDiKxh8BEw2CPh
413x1qQR/0A8msa4XyRcmUOJqMcHgic4v3Yt+t/zzgXXZ/LwfmzAy3t9NganJw9u
Xpa0h7lq6KntYD2EMXG3g7wzFGeXVk2DKcLTzkE0bIM=
`protect END_PROTECTED
