`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XYFjr1dEuRdJvS1tJDfVAavHCAONI+JYVPQML2l2nFBMlycn3C1yIhN8j1Z+0RwS
VTAsBoJ42QnuysrTaHRm19hNJr2I2EJ+RwlXk2I4C4LHY07UwglWy7ncEeCM5Jnq
d7bj94IPEyktih80MgCIiZsBeCCaCY+DCxSE8h59aKCVLuomzcgd7D6iLSz7bEQU
Vi8YYZB24Y4fDRyFfRA7PYPAOpMZ1b59Tclt/m/LAAw=
`protect END_PROTECTED
