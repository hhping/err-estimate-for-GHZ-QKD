`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zaeAByPLTTT00y38ynWGOM7xxWSMGIEHqKRLefFtTUXF5qgCDICu5agjcsRjlj7
hLSHoVuKMSp6qF8bjOitCIiBQ7L79nPcroGA31vEriVD/bRHhDGDFwS+5C/AZ6N+
mJLxbSudBNB4qi0RXFP2fez4yfL0NAJUeO67Vpcx3kN16cBIwo380wX/tobgNO//
8O6/H6ZIISucu+zFOvnvQ6Y9Ex/fYCFqm8t6hXNpM7JyN4fHKHXaqAngoFmAny3m
yG1WH3MHDMCCU1tNCGBhidlvMOe+EbDdVrp8UzgNh6bNetwGQufhWrRAtsnNmzdQ
JkWTi4dd+dHowkgtV06FmJH1pYhN0Zt/OwAzkNQaKR0=
`protect END_PROTECTED
