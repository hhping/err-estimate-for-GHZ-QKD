`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cHPg3re/IHVUCWIlqEzyxSZGcprSK7QOymF/JZST/t66nHVN0gxJNMezE4ZfgfZ
3xYYghPyxbXzXCYNV7Y0EjuoIGyU3+Xd72TQf8eCqFYTcw6Xy2XFciQi77P4gnho
08wjipHDNpBfsIFCfb51XyDnRfF9Npm5TUgqr4actj71iIEUP5YCw2MNrJUeQVXg
uEKsH2eH2ejRy00XPhFHMp8x+S1pXUtkRKs+9dJd/z2XKhtSQzwdQoeu6eL5S/4F
kKcJYNQIYNqufPhuYqR9u14nnRFHg0j2vskXkFmV/Bk0gwNU6mCdamNf4ZTwjZjq
RF28KcunFEdQbjfm/iGbpo6zxvJPXNL7ES8wzf3+qVDW2NsF7a90JrsYTOUAxeer
+us9S19SWWDKmYMBZgebCIg/GTHTVKe/hAH3HDWuzuXW58mPtkAPLChcJsjjrRvJ
aczsoeHueyRjh455lBgpT3CjClwGm1XAJUFWz7eRbtpaZZN8dVvNpTleDOi6dRmQ
6IA9KHkUobfYTcLJ8BphraHIhJgAnywBAVqrwvoyEJQiyvsvmLIHmOH+y+nWnGJr
ZPHWvK5+9T+9aKjO0K/0NGrbiugfVonUd9xjx6yjBx/A8XXF615VUPwRBChx9L4T
rRCCDpUYJ/QqlUfFjNIM4UGQYtID7uzzWKqTlrF9YhwBrChD7sF5VkDkBjH+dDDm
1Tb7DYvx+UFNEQdQQ1sVw6qWB5wmT6NqrzPHznVamqrVqZY1lLxTlIh4tnwf/P94
dIYxwXB97rUSecox02XaJOFZ2psBpZPz8Y0fxniFlhjuqyxSusbZMRXGgdyDXpvh
s+9hwkk2esPX9b9UcoRdUA4w0dFL1NX7wP5j/JegnGQJCRV6aQoa9gU2YM1pcEk7
4/D5qd78TzK0mB6p3MNY6+0ykiJ39z/mLFwC6maR/u3q7saLhVIGMJpoDDt0+/k1
2WPneUNiE4p8QDdsHV0BTIX/aKuOwWAnwpJengNdgamm3v5j00I3y2gxjLcmg9PO
Tacb1FIqCtyHy78uwVw9mN4Y0bpjKBa8TGHC5MXYCksGIvQVsUiWaQfWtBwfOPgB
RXZ1qg5uYx4oQwMFN3WVXcsOV4t72frI1SL6VOv8SBoaufJxS14qUOanlDHZWJC4
osAjkauh3V1Nd2VmzyYnkN4vvE6WFzXGaTSon9vCMRDiW3VUtUUol6dLjfv3p2n5
cpvPSy9+CGrrliCutrGyV2EPvCN+CeBk45pjfqcnJYezsEh2re99IrJS/6tGxKnc
oBa8pt6X+yPMgzMNyxGkLZ6L5kN/BwdgBw7bjZpRkPcsc5X5Qc7VHLPqdrwFGbl4
ZX2rOnKyD5SU+r4mHpARKZ2AQaWzRYEpfQh0oZGcGEyF9CvytoqYI7AU1e10uGcO
XoJU0c3ePQTMES8rMcD3M89PeDmwhQyYuq2GeYl434qedE9x+6KLUlvMMhcoV7Jo
5j8iF2WRVqNnKeWa/bOz4sggbTlnQuoxnmfC1URk/R9QtB2tS95KiSSo+VEiChkZ
y8n5qw7jlTutWS6XFRUjxzta/YHXKId2B40loAH9ovyzD0EkHVypF1O+f1kF1V37
6+cOivcOgl+wpVzLQ93Ftl95XXAlmqXIR9CMrz/94RFm5Q5Zk9h1NvZROXl7sI3Q
oqhwuHW2OiGrHYh1TdRlh2CdAMJOH8dt9a+Pm0NmIFWFYLlvzW2mFE4uVICr8tzg
SGuVS1rBgcV/sS+X5qP+nO7BEofMnk3IhnfBvVY1xAVRADFzAtGxExXWsrY2ki3G
xH9FNduC5Rd3dn/ICqSEee4xGTgiUg0Su3f/haJQheMX4EJjfv5CFgvzzye9iOPP
WBVuWNK3COeunp9HFvEQ41K8vL0/nGl6GaCkk7C5/UbJQxtFl1ijjaj6HT8ozWuT
0cTqpLY6xyRhyIzdvbc5SWPnSADzadURvo1gRygAWVMXd9utLxisJ6025vJNurYX
VLlT1eaqCr/BmIVgGSzqdPRXmZI/+sdpFcYtA9XJ2FDQ0wXbuOFiBTiumqjGwyLP
992uVSXsr61b60iPw35D6nNbUkpUbUkcjE5dM9OS+FpfTqgI2veGEKseYIcPNpcD
i+ZpbCXvHcMA19p62o9TVl953AUp9XvzNbnSvDYkntBG54aal9d2T4B/J2XXOB+I
1XkcdonpJtG6Hgl9lK4aEL16L3OEDEHJvaLb3kwrhLAv+xSwBiBdjjUT95LcwvV6
EyNWm2s5LIX0hU6jWDiRsPZxwjqjsbGBsAauoZiAYsxMvGJeMNO+v/2PIWjrl4Ox
g4FLHUYtnp60LZfl8YgOrzm+okuwN+nRg1oyWjLVVWbMpS9Gdw8/DNSGcFRagWgQ
BvelhLI7J3IB8+hBs6wufQRwzrmpsI6qUvq0my9KJZxNM7KxmAOi1DqlvfZQpU0D
IG26Pbh7uzBGVCHZt7+Bwl6rHyWvn1gBDTJjCepOEe2Wh6YzPgHwolzX9tv/lxgS
JMjfKhxSFKD6ahMLvukh6+99svqJBGVS6BYreRZv/lLxUVKgB9yp9C7ELKLUe5Dh
vW+GIkqH8zDZtmLRL7PtfR+y+oXes6WQ68xoeeGGUC82jKhTzAXNZVeuVNkMbqx+
oBbV+E1wyjwtnGBDxBOOfH6RTC5J7wNSR7DTHbiUydkA1U9c1+H+nY6EUxHiEbdx
aAV6rBAfbowqgCA/71tWbO9x8IoowO4jCc1V+4iTq6ZeHpNepbgSJ+ZUVtpF5P9s
QD6lt4d50nmWhOhxJpgGlZ3R6pyn13BrCx3xc0zenW64afdziyS1V0EawFddIrxa
y2AEYB2cC4Rc8LBeAKf1/xlA/ogFaKZ0YXn5gHh6qQtWnbOYfMFmAsF+VfLr+DH+
3jkHld6CpTQ9najV9sP5yqtqHjIoPMoPDhIb4uqEYHn5ovV4WtlXjePJkMQrPrrK
FBSSxn6NFQtR7qEJKVBt1HbpC3lSE3OtbsqC5E2OIE01Qq5sV9aET3OwzctCbVRO
jRxJGdDFTFPMwYpERNPXEi7P/8xRIgoqsx5aZVgYXxAtYJKb8zzrPLnn3lx/u9Qp
gqaYkGGGrQocqunTg+t663hpeU2ttlYebh7PK0KW/91tn/DGtnVtnJECu5I+dkb1
gB0Yf9ZGQF8Rb/o+jwkp20SxztLd/nhNcIUm9clVF858yvhXP/tqvP8ES9+8JsQL
pycyELD4PGHUr/+Az7AxUtpgOI2G+xqXE2SaDPbfIJEKh2zkoAuVF6rBg/PWB5qc
bV6Otk5iFp9ZehS8lBY40ZQI07Swpods8q66213vvVN4fvzZLRaMuzaq3FX/r7Ty
P9felEvFc9acm4qWHizQNMgdvgNyrpCoXM4wvdsRfa8vBdkYju5yZ2YhF6jKXgNl
1ihwBbbt6ubLmsPf5HMECJnh0Deo650EH5wtodqUixitA56dN4mMa0yIzUN0vnCi
FJ97QHk86hLVZMU2+G78IwjojDBN9+qt1gbJWLYUqCehvKFbsPlHFhaVDTrj9psN
P9MMT1LIZOM5LEa28WB5LGj0PT6Q6Gb+s2uBK3eQhXbtMavk7WwQq69p3kod5sWv
7S83c/cHs06b+HlMBKHfdcxAxstm3aZ8CaoiecVOR+KwgKfk1x3t3AObumyCBIRH
Ks60tzGo96PwNHif2IMIrK7mvwYRGoz0TbKhu4tO1SdLhifJWyvhmbCmoAI+JQUk
DNqlOMVv64QzKRaCb0nJCXrATMpOEY0zNB7oRwxEpxWULpPxOBj6AtuxOtjin5+k
4TTRh1bQPM7S4NXlpSRmj6VTP5O3OhfRRQSRGIAbUkQ2ZuqYyFaK+3f0gucL5K0P
QR2q6ocBJAg7d+vheuMRm1Up+ZgQwfjXFAqyfLCwWCDGorNDCezWYq3io1DYYNu3
K5jZR7HReUK273gekuheXi9k3hwmF7iIY3OJWdkUj8x4tSy+xnDVqLbo/aAKzdTz
4oCxEfd04S7+bSPkvrAWRlr6wG5C8pPDxQZKx19lw2OUk3T/skIkNLLOJKo/8+45
YHA1ZHnSJ82doDrUzAHsJO0x6uPyKWpjv+qs8Idf9QGAKAzclTyK70P8PHBS4T53
mcW+vLLfIRQYqGwhnO4cSgHyUCM65GsfFtiVkPPmSls29V/FOSkVvyqJ+5S2wCC1
gAO1/mlquSybzJ/I3fTyFx/8BLHEMdC+FrUBzT9L72yxVf9J4+hhlrOOqPfX43Ni
o212MYEYgTr9fbxk80bpi2JFWyrZ1zzAr6PESx6dSpEf3hrxKjP/S583PWcZlpjG
B4b96jIIJWiQamfjNpgilcY3lLB+dp+b131uMVXJWiisdoRt6K0bqgtqXyfeys2d
tBa2VRiLpXlqk3E03uxQWnsC+ymtxDPp9vZ6Hg9IaSpNukClx9nvpgN0rG4EEzCX
YOdhiv88qymo2jY/3XtIIDaTdt6/WhBDKuNuUVi4pRRJn3VCtIuK23uSVd1yJGVw
75pAwDt+Aekv5JEH+3py3KIczNnclhkZ4LpJi1XhfgnyIj/ECs8q5iWDm99iJCW3
jfrEdTnRVfOYzCajBJ4mqTmPUsMB+TImF7JNZMfZAXc6tIDojZKtnIpBux3tpdz5
IVhnbX5h7UTVtxfkDAZOnL0yE53a6juXTeEJ8ifkE/sI7knVwP19W8YpgseK28GW
R3n1VloADnJATUvwp7/vw/t1IS5u7tFDuhqPPzYICFzZmvidVk/W+GWUmE0oSUBk
lirXbqxjKclMhxaGByCFugotlKQYyRrlWi7x6FiAz89i4zYQYG1jK/RdY+CVCduC
BI7k9fU82ct+naGfTNIpLslopth64Uc5xlqi6rL+oGnqI1Sh76Au3HGzGbX0v/pe
g776A8uTlXgDpIJpldvr/bf5/MaFMelpBxe+7UvLs8bHy0wDgyNE+wLN4r/b44cz
8aCCcAZCOmsBgTeAGNI2tG3G7E+mixSFbE0ImCEveRDCRTyRHTuFwSKIOqugOGEg
o1Q8bTMMTCi9MKpF5GgZURyUgbRo48FpZaXqN8JO1IxXCCJSwUkdEXOoEgamIm4V
bNCAqNFs4EERSBPlRw1hoWIHk2ugs3TsssTjGMUTaBSCeMc/F2bkaU2osAj5NC0g
TOWZgLyXhe0w18udnXN2KRC9BzwNGmxujKW7an1B0CSga3uyvo8fQ5NhXSZ+58S7
0RyDtJT/WTDw3/C13UJgYOCOExZ4T+EnZLtfvVLwYNKCsIavqFCDN8rv+vUjSaA8
nNzS+VUyJtJWHIuSGfSQHgecmwRDirhknGA/tZuge0YIrb+Rckz2/j3UFGGEumm1
v/W8Szeukd4V1283Q7Aii1wU0cZDYCf6/XpLRMkatUyV2ZSY6cVUhCwuUE4zUQMj
xW059sJD08zi05kM4gPY8W9MHYHO7YKAErnoTwsc4tIkGoz7kUE71YudP6G8vhYm
7ZhcQfNwRWlgBgH6QMBF1b1ep5EG3DJPRzSvcn9ThbNIGSdT96w6iavsnn6Zu4Rc
nbbKTAHfyz6eUDWZF23PzsZUvxhHG607OUelnyKukAszJ3mzNrTDNiXhu+1WR+AH
AeDTM4yaNhRz0bvvzKS71DS4nszm1GPn20/6+3DoFp7d5dhPd7ZtLbvryMb/AqHr
my+J0iMf7/QJpQls4nNLVhIltXHW+/DkwYgDJRXs3zrO9sgGEGTrSHnSyDIcbS1I
nkUlSXCkRqozBUcj+9yigt0Jq9+eOr3F1frHfyzy2/SAKQV+kQmFlq5Cg8Z0LAzq
GkHm0ND9AbKdSCQ5Wn2JVvbKDJRVr9MT/rurORhKDsBpN2dtJMRtF1cu4f+Es9HQ
+x2MupkYqWYEnXh6lxMLGoQlsI77DOHA7/O583nXxUZofhKL9kaH4B2QopCJn3O1
KxwAlBj7pFn2jwYQ02Um+gLDEXbYSQ2ivZ7M2GK+D1js1393KFBT3/qXELDatH7U
rxTG8RklGIdT9g9Ts86Ci+wW7qdCs8W44eHhUF3+vjN42KIrPBxxWxupAFj4+fgM
iCRV6qVpdMahabiVezkn2exTA6vY7WYMx0WbvsGDPqkDZ/DswCouiDmZPCOHxdWe
AtNDh2sHYKqSd4YZUj+O3oSXnaJmXWkYdJwnBLOZIoTP90LTVBlWjSyfQUyoPnT6
3PRVJPt02fMg2Hpwatfi1KQkgyr6H6NEjU0H2rI120CVBoZUAq93XtRO1zrFE/zr
aQK3ZyglWrBxaL0Xzj1pBj3jg5MU0jnDSEsXwerdGFRy1YQLigpqYLWnp1UZ9K6f
7Hm8c9AMn5VNFyPEYf78Or+R9VEcJfslD495U2I5LfDrp9aDjMTan0L0tjPnOCX2
fI5VPG6TRaGl33ewzo3Z+tOOpkcH/nqOu1A5Gj7Y61HOWNPH/keaWkkDtx1eimf9
3GFtOXyQDcJqeWFECsRTJKpnT6rGuPbJBsIR9bZxjL+Bh2AfaQMumOm36VqCXcf3
H8ofj+Cpa+gop3KMvyBbQ7kil84QTKUyQcld7wlnmMHToKb2G6A1vVPN0EfwEcHN
ko6wWjLy7IDjkh5LCDWU4TLB149IRE75lOfbAfOVNy9tLUa+5o2dkUsS0WZlNRhs
XOQCWn37wUo9qpteBH1TaNLSsglpuzFd9eWxHUqTVtaS6QnV7cHlNAY6hJwobg6M
tS281s/FnZ6VwmOGs6EnHrbqy6KwM1tplXX+3uJsL8r+jj5yiuqdbeYM3HUmNSZP
sC7XvSyfnjbWjPyjjvVrf3r0XKh8iO8n8G/UZ+45vvDpZ0MKreHUbEjkJvgmQTDm
aDazimARn5H1AsuTrzlTfB259+TKCLoAJFCy7GiZBV//Zu12AxNwpdS5YBCfr2Pl
bfU43KDSI4QK5TTLa12wTqed8K69XfFgmaWmAEGBNUexLwxlnROnHrYweb40Z88S
tFy9vRiTmtuzeIjFkG8YIpfviotoGMhWw51xyYsZRpXtYXYGqd2y5MKZCXYo9LDn
fvZUxnqcBZOuytkzLwWZKds5TNrxK+4el6qwrHQ+fANtExEF0UsOPHIge5eJ3C64
DOvJkXXKpoubDQw0b62QaM7BEihyq0//uSLR+hFczv6yVTU6i3GLx47NAMK4ToQ2
GO08Xj8+kWS+Vk1u417rZ1u8Qui51/qawTqcsdm2dBGZxpzIe11pyFqbDZ2Q/M0U
QARiM9g8PyJTOQBlHZDJ4kaufF8Vn33/Ucbgg0qSXsaYtPIZHQ+A7NYTpz/Ln8Z3
VIKn6FV1OMbMy8EvtMra0FpWZPQxa/5jYxVrbEqKvFDntnm5slep6QbZ7mgw7dYR
gPAYu7aSDVPUGGt7EzblzjCc8xdXI4ENyYtmche5nV9bsfUK/DrjkaJWvMWR/2uI
4ZVlNfyhcmZykZQIXG4/0+nE4oLmmGfFVz36/RhlV6JOUSa+rwUdRNeSjwbhDLHB
uSzapP1gpYmoEGS7svbrv3yWAp3xUMMoq0pxcMcmo8IoAYcLVlj81NTMVIdG4ZNF
I9ljUTKNilAaU9Ma37JQF2VcCUrCIqMaUITgEa3E0zSHNdfh+dbYQC6hZh+m7D64
PNyru0tCwdzCOFHyZkytUjHcdznugSD+mfJm6krc1fRvsfyOB5Qc0NrBPd5zSwtu
s2dnb9LmgehT3esP0LpyWpU0aQ5Noil1I34tlwPW6aIh6JLQdZVQ06i3c8Mt/gAj
Y/yPJ0ljFaqfETyVr/GykMUN9vZyJbDOQo01TdcDUN4doEIfi9D7DN8Th7JxJ+FL
7jTtVs6phhyPJGc4Hzjf+LulACIbptRkG8Fv9XGK8z1HktgWe2lLoV7WEOscvEu0
xJZJXRgndiTqpNp0eEXVpIdsfR1pXH2b30HUGd78Ph+Ld6yzvO6/tYfsYg+j9TI5
hd+huKqombY7IVGvsYt2wBok4EUJgr7VZh18QzCzN1F+Stn1QL7FVQ+07qVUY7kk
vCKRFA6LxAsvKoOsu1PrVN2x5m4Tb34ZOnU/l6Ct2YESx2P56BX4exioMHqjSll/
jykb6//l2ZqzbziWTcEH+LJNH0Xp8pMJ8kbVsDQEoiyt+Np4f9RljKgKHRiM+3uM
wg46XP0pUCSStnzp/EXr/fLgi3oNfTb/vtyC+yuFp0XxSbTs8z2XrsHo8UZ/KUcy
dqmtFuAzpr9lTQuWetWWNNoM4hDLplxAgxx9noDW2Daeg8S3NVlm/Lh+gauuOCzm
XL/YRpKZ2UXgxQipwHjfoweF/sWM/ObdNBDFiP6bRIYpfxeICSNR0s+gynS4M+7W
NPrZ0Zvo7Z1erQDbx24DUYpf1I0mMRkrudb6k4kVvub7MvOuDOYUbFuuTwUDU+PR
cD2vEhszUGCQKq5tVvGQc8L235EyK/BNqxo91Zyrpqy+zB+DJxi0D1KmoOScp4Vy
Wp0AAH9h+sLKc1baIm5YfYegUpPg2b2Hr2dxwr9rAlGhiXKHYy3R/IdV0OSrcdY8
zB2z4K0bZWPntpaEwv0277CjcrlulLV17MAb+2X3wDI+tJr62LO97CRBjZKCNkFi
7tbNSYU3flv0pnS1xC0qVtCREw/8J9q7VhCq8O03TXRX1bOIIZshQcubCKZqeo1V
XkPAN4po4J0gvFlYyBCKcsFRDq0ggy+ISQO9vDdx9wjh83vnq3fPnu70j2P+WUaQ
2+rLtuwNwl6SrO+hPp9R9aQiQ7EgPlbHy+rayBVCqDiskckEK1TzaarCRYHw0mF+
NW2anDZV4ypcjLsgWhhQD2DWfKgY1nQ9uBE1gjH3DqqgNFjYPNQ4R7iQT0o5+ppK
8Q0KtNNexP3AL3Mua6ls8nGHJ264zbo+0BO95rXHK0uti6fjYn8fpcaEC6x1OoKR
WJggINpaxPYJNotfx4dAc4+MUbQA+AnwJTBseVp6K/PgjHFAL7Ql5eCn2JWtyBtc
KcpsO4ktSBqizGECKe9eCOybz/CkQjNKJo6WBx6CS+po24jyNOK1CmT+PtQ0ubMO
+okHlXd9dmo5OeHdGKDZ4WalPL5EyxK80kM9G8TAw20ipPJAn10aDDH2nhq2sVnR
8nTnWGEIP6ExVDxwaHAH054p9IRd1bWCZtvqD0FZ+CmFtYWLZUH5wwkgUgK0cR1W
E9Dd87Qly2z6spGZPM8gfSuIvb96D3qxK/w1baQf9rmXKIBLW5PsblVKSufbjKlV
6493AIXR9XPpYJQuj70uir45DWHG5U75ysgQnW1YIlrqzBCYGNzYdzECtUkhhb2k
auAYGFhvHaHscwmkkwsqJLiti7yKmdoBj8nEVP94LQz03s1oeQvzN/p3fSfuaYUN
OjCIa4bflSgYL/PrPO/MLOrp3SZEc7ycvO+RnbMFoikLdFBWLd0KQhyyixbm8UAf
3keqHR7M6qCswiH0+BKOWhEz06mPSTRB6hvy6O8P1CqyCFc9TO8LdNGvpelSkMOE
BFQlRBATepsWfIns0v44wVxltsJVZVsvbTn7T2F6AkZXbNFrGdehmSV6xlqC2pJa
sXES+H6iUzuMhHEj5VkPbWICU2a+w3Xr+A4gR1CqgIs/ralO5Kw3D4kUdgaVt9R5
SuMnyHARNrwM0joVuAE2cfI4f1RJR45RvVo5jSroLnFAOcN2MkR5QkLuN+WMfl9b
p5jyoKdUHczDcQcVSfd4jY+cjF1xtU3BqPSq9OU3v1uMDeK9O54GxJj8zxPRiiKv
7kdslj1sfdj4Cai7/DPY7kSATy5XzVcL5yCzHsyU6iVKwOVni+5BUzSx0FPPIccy
NMsRVlyL9plfUPXWDoGUv2wg6XjqQqmo3//pLjy2FCsaV5c0gan7QoZscf8Fen63
hNmY2BISEKqRoA44LiC0TrdnACSLuimge4j2SNNc940b2tZCoiAy7lSl9Wvf4TGF
EIh1SHlZ9dMHdlRDpdDpjX+iGac1kg4U/FSA/Rz9DBkxrD7MBp/s61i5NiMvdGbS
bvxgF/oCGNqr8fOT1jFHuwz5FFlhgNqYV3whYcEDutGZUBXwQjSN3N3Df7HQcOn4
2BACtxNIGaz5YYjnwmrAXW77j86zCAjiY9EnDMYV5oDzR2MC4LgG8Gxq70JrNcYU
K2LDSBmj4bkj5Tf17Bfe1qUMS6CB8nffrvUNwty5jy8ptVokS1yfLsxquOucjwxY
95mjys9TjWlpROhrij+7vtK+MynlU18hNQ1Fcje/fpj/KZ6fuM7og91W/QAnEcjR
noTOImozalVoBfPljgEA2CFf3M9C18sRkbwVTh6WsH2YCsVmd6AxnjQVsYRfNkAu
FHA/SBPQqQMgXu0dPsUAn/Sqq4Nmi4GX/SrauG6t4OZPQ81hfUb79CFY8fqsVRqM
WPZ0z54+hf2us967+B9R25BCaE/0pvkUiTzMvtM+m++FYuh2xOIgX9UdqQrRnOW6
QzvCu2lcZZU3DtSM3UO7IOBCgotf4HcjCrXE1MW42j960Ap5bW8sta6bb6085AV6
soYzcO2NlvJUj3a/uEIu0LEGRiYIeXJlgAKZDM4qzLa9UEvEPaibb8klzxtfp/1i
dn9w1RMF7Z3oYtflFUWLag8cbCJK3fvme7Nzq55ol74BfSUOhxJ/ILz2N1JF9HQv
liVLPWy3IHL4Id29SsNkiLbwLYClLPCLF+ezL+/MnnhXFQwRkxl9hKy+uVwcixfJ
ek59cHSZoANiY8ZWzOEv41Ktanpx5dj+hEQTJbz2NcB4lOVMvV8aElfo3IqhQ2pH
r8t9eIm/P7Q1XzxDXFHgXNDjUVkDfC2t102d8wRr3dQjJvBKvQeUP+wruBWlSKx6
rRbfCH54rnutnlSnlFQNvRQQcQ/zhySMzTUdvQNECZH/zA1oIX4SGKp5CmxSSMUF
J4NES2eSL0o7O/4rHaPR+H9VsjxeTpSxPS8xPuZm3Iy3xzF8mdBVPZtaU6ymTW9y
qO0oII1y3ams+96ed4ddkGYJ3sA+dJqIXMXVjr2pXzfouhIHhCDjrY6m92zRQBL4
EhlbywgTUUxfHvgq5xSoY7/8UeHjTDCqnEuHDEtQf/wC1HVS2qcC8dBwJk/lnWG5
yrKAMpQe6CyU7MOUO1YV0dfcEgz0hzyXfBIhZSNrch6EJvKdGqX0pDcDqbeslS1W
tNtpDaau+butHqvSzFavoKluWW8youXpHqnLLgAyrLATtqp1B+9mob80ipULmwhg
N02ISo7AkmJq4OJHDNvB7Bhv2JAPTERBN/c7R4NMOT/EZALH/fTP54WFgKEPypVm
mrP4RjPXiKsZdGLsiux+vMa4SEnELamzqEhLcPPxluIh8BhegOgo6pWQwP/+QdEF
XfMvGim1LTKyclQYUbtO3HbzAV5Hrym2Dn3d+W6z5pLTsjzhAAQU/hsPY2lCwIPg
s2wje0bU7wZhZG/OA98N56SLUQxueObyY6EIutQZ59hEQ0jBfd1zcG6wzSlmgQKj
gkVPOSz6syEdvyjgFeVYHlV6ouE+gtf7UrseZdyHyiYdEaotP9VvLlTaxMprlqcn
knbrvumcMzCtQ9OcGiXeO8giMgzfwyG79NpXtRvmYYINerUnr/6j7lC0NhOIHnqm
wNHVMixeVkHPNARdRyftB0flNnPJebzT4hTtTq03ivojUC8kkNWJONsdg5DOQIwA
pZIwlkkyJqZhJMts1CkR+Pmy3mqsjXeLBXwHv0lanFk+YDpAK1VTa2b4MPXxewRe
OzSeDr/aoWzoAypMsAwLI+dQf+HT8Dnbjo3/2F8kDFvesHUAjKcvCTJ7Lb33YBCT
HKv+xnjFXGlKVFpS/yvjSc/CRV8tbOQCxLBQEvP7dqDN0aP7W06S6nJcBVeezTlU
IUHrRZA1fB36fmi1JZW3GVKSiRo4ZXklNM9hoo7YhAwPy6NbmgkhMGdUjP87Q622
1b5LjH0OIZfuoOx2QN1lspxL91m3C5/UFe2+aLbZq7DLvtW/XVmfvGSIPA631Tbm
T3N4aVhCr7agec7W9qEnMfsDucuIVkX2C4EOvg0ALx8mTKGa6m30SYSHYlEbyF75
2EMhoj6YSnaH+OPEKPoPmmIGOyunxkfey2kRs5Cd1weMsr7XRsH2b7iyzaN5Ftc5
EwToyu/Xsgxobt7rNUdxUyJ4x6vV+N8qKKZ8z96zaBPc4LsE02OXS4VGFStKnWDR
ZwqznXewoFCxN9cyqci+jEIMBHjhpYia1W/UyyXZt5Px9/lIMN2x34iuemZ6CeP/
GS1hroE+VVEkwqFBXsgEqBxWLS9QjSHnw3o/Dio//e90ApV094CcYLHx3HyGsIAC
fs5uYvp8YObFZmxRY6A4hHumQbX+AbH7jq8pZdigl41f3NNOUNE29rG4Dqlzfnec
s7u3jcuu8kz/PIyFuljOkSSrM3obA0Atgbkz703bzPoIoHPYMy8ifAomu8MQZUDt
I5ZKl1QDer8Fi74mInGrbt6KgTCpVD2lnsGJ69UfhKLTLF/ijPtmLoUrD/jn9vjr
IB6FoRlLH5uqbBVk/4Adj8yivd4uwBEO6m/SKXTWtC7/Kb6NmZchwRuW7zNlQdM8
IyEvXtfLeIjClpcErHil628Va9iBDDgfPbKyjSQMcGhENhnj/ChnUpJCkVqxBL7M
A7jy803T+FiZNY0BHvBtHPO3H0IfKEJ1oRUxe35iNitQHpozx28cx0o4mPU2TEkV
Y1MMjs1JpvKga5oBZZbC5IbTmG8QO4xr0/lxuT7Fd+QkQL8SqdaifaCH0yVvyw81
VxpkE4Qe1I04U7j+L2AAvG9ukZO+L7vzDYB3Ptw59jhueBRS93luv/Lh6WkMQknG
VhFKRC7/AZDj4+bUT2xUJ4H3D2vhCDhAVhbTcdzWyHFNWSXXaPCjyf90nWnMqVVE
nGETkvMYhZZ+q6ayn0lfKTesMFgn4G81GHlk49G5Zmsx6WPfBPWZ7UDwJQ39Kvi5
c7Z01G64pZTCiTXmHxv5ITMqTC1wTnn8kTd3mwP/+mrvLfMv+EQhozQsrWqPbSo9
W/AGPmoHKq5/VKTAF3Bqyxo5yY38boM7kV6l+YGnO9HMjxlBzIVbpRWvAhkWrCLZ
gQS3ZFC1i8myFm+rHCjAB4FfKjpgwjQc0H/GkwMT85Zj98C1eq2z93ihQEKVJ7vC
Ydeq6rzjjOdzmsVDoZGGvduH3iHixuGVKLEk/G+ODjLX/Z9PC95Y/D1ryltdsXTQ
lymNeooSp/n8wMyk9l2/qG+xPVLLIrhznnqmzIuFBZ32ge5fSXVcHPpkRq1tSKjY
nUQNQlpAVuPPxr+j7JU6zFPEWTxNlcbCgwercKNHdrCJOwJRqXR/XAiOJfyIMCKc
PRda/HoQWUXzD/5n9PUQs+UvoLHPotTV0bTHt4tE7h2lkpkA/jU5Uih7HzgzKfk1
7pVR/SB+B7+zdBM293witRAkXlHOPCokn/PQYmoXsXzk4ntJ9I4NjbzV3PWNKTnV
e+AQb1wGi2dJxC3fUS26Fh3njCoc/G9++c3UpXo1nljeWc4y8spLvNJG3CVXgTAG
xFzxYkBHi+wtGxvObFJvj+SAC4g0bY/g9MVgYWv3EvBiDjCqOjY76cAWS0M7TQoo
3bDO4hs5Ip4We2C4cNvwtrVLCBjKGm+/xzYspo0F32oonilwFwLYt99VU0CQ6eK2
Kf5jys4ooemQ/S2wvZ3ARHvLFz4l6IgA+Rhxo0tXS6kSBuYHWwF5DeVammh43Q16
555rf/udh0jE1B/TIfqvitSY3TZE4mNhCLtig6iEtH75Pv1H1dHu2FSd92MLCRvt
PdPMv4IRnmaAOzl/4ILueobBJQ5jHW+kwyCVM1Le4brU+/a52qCQt2ymiC5QVuGM
tEo1RHu2ZHd/XLGFFwiUg4iVSCHy+p3TvYxva13W3Ja8MM+qkdagKmePdkaLhSqx
R0fPWIRVBse5suIxAMjSHEnn0Xu4YHAuUdmtYVjO2KN8YmCO9i5dJgtPs8EySO2Y
7ILj09ZuFg4+KEviK1whsukAq1uQP+u5rn+MlJyMgmxBCRb8dDQQAptz+zpLeAcs
9LPusxTdwhDx8HgWFh7xXu8Pq2BLMn4leaAd/pphcKuVCKtxE3qHVyUS00zm/kxM
humHnv0tiXxLnjznIRXC6nVzhuZkgZA+SZ4WCJVb7ciXSyRJusEpya0W9k+83qg5
vaw8xomWbVQA++ByYKJ3S2U8fNxZUe96Q8w3rQ5yn09BkAbQxiPPhLLFUKlsxR92
Y/XlB/9DLiCopqGjn32KUMkRWqynZ3an7jTiE0BGP/nBTK3wd+NWAwtZeM7+OXAa
Hk7X1Z3Y9g+z644j+DekJpxODnkJhY9pgkZfXqHCfgfRdlMAs3mE7Pvs7Q0WYRM/
0uUMf/Otupo8FfZTMmIyRfymNiUCOexFmQD/K3fB9xg0X2c5owtRrZTCs+fvCczc
9FH8agXewWAT+GoRbgk/kpTKkiG212jJVgxlSzNdKQ6Xd/lARM3KgCoErvtjFC6a
Ip5GsjPEl3zUlDFYaURr5DsLTGfJILHdNlZDeVMPGJERf9Hvlxd4kT6ZBuYLNnwI
s7xXdzRE5RxBj110W3fbCB+OUI51d1eVlVLekrW5yk84twyADSVdMl8oq7Wi0e3/
pk3+xtuomhVr0EnbIa0U45fQAWzAmDHhkOChjoD2Fnl4VroJzLO3Zo/Z4/GubmO9
rO/q+IfkihtQdrr64tGtZxUpLy04dzq35R2PMee74I+aujQCu19N/E7KNEqQhbZv
6QzzGWBijd44v8JiRobuIr4jCHQeLxFfzjIyOd9s6OFyFA+Z/ONFcss/JxS74A+o
F8xQOoBRp4EUPCgvz7cmXQRqXCN1b1TcsdHiFnpKbS4iwHZYE418DfPYtiN9gmiD
LfZjeK3ofOtgSy81BbivzaHgDrugGUU5bBqs7k2PiNLSvpSbrjk7HfammwaSwtyP
/qrLidluHNJe/8fjJjaTbmz1dIMJ22AIRrLwheN6VUfa7rUNxAPjif/aE/E5e7Uc
Kg7E8JwoDVL03HYqP2nTZyoiqPbo24PDaoyxfZTfS3d6yF9jnSqTDtuGpELkZnz3
sTZv+YZLgC8pwH5+zbbKSzfQSXK14UrCfJ6q+UQMfC7w7GpSrGSTXG1SXjWkU7SB
7JKE0SBd/2639hd+YerTTVB8g9RF5hvyVYfHZJpeeEWfFfV1DL/A2Xx7/NZQGTz5
DtVa0ivwWfKY1ppOaHWzJRqNKivFERz7981Wba0+EGMWOwXXFPUIPPfHsSpCGRdZ
6zvalB55JqDTNkaMNDSbZ4h2G4PnSx984w/mLHD6UNg5UCy+gpDlZFh5FZjaaTBI
SbEZMMbLOJ+i/qfJhg/twpCPQvqbHRYzB8ey6GRc8M3U/RRrW0UaOj8FaESPtrbx
p32XFQo6jwmbao0qN1avPET1jTdMRRFNBr8i2cnBAlgtibgM9jbUhl7sq69/vmhJ
nXtUytfU32305i3v8AoIEmuK6PItat/Nb+y6X16zcAakFkqLMwtNfiyly/26pm0y
+07Om+HwStTFJieeY/Xt1bQ0AcpQlzlcKar0rQBGJvOb9s32qXUiNg+RO1EZAxTJ
F3CQgGigkOS0zni8vxDKA1bug9Ldrn7vuUqEzFU6J6ztIZXahfUKAEfiu+tLHF3j
eL4th8WkxAW953qmylAQtzfEs4KLz9J8FxJ22LEVCIFmG3YPejc/UPmkNDCBwSw0
vMHZ9gT5dwfYRoky4zsb0iHgGlw0CyxO6qDoa9CqOOQiVBvFWFzV2rhlG9tqKSHU
bHSJpcx/WOE113zvX7x43z9EAoGxSTY3Kg61tRF80S5NENS5LvKY8G/AwyNv/U5+
MFHF4FlTeyQE5XEd4R6bEGcL408vZSwWNxRLE7iDgo5yTC/agZzrwXJJmfO4lf6+
1Z9UkE35pA6YJ6lyPcJj0x0MHEpBZx3LaKVXmoQU667rPCsdfKWfo/ZNUObXHuSp
upaTUAtJVRziYg9Qo7ifAQQ02kxemf9Zp+WUEFaG4FszsOmTs5KnEFp7TpC6OTX+
2XLVNbjFfyPJwGyqarGpLC3b0GvZl7a/YNycI/XZdH7nuzDWQ8o8DLHJigTfhIEV
HbAX6ykyeqi+zts02tInWT6MCq8rYPnWO9OVlXg/nCHcsQodko/sX2Kn3q00EbCs
kKpZQbQA/gtiiwA1A20KcbuRmuAoWf4bxfqhKSohTdKjnyftBxNyv6grqkLa9l3R
sNzDHdLUrtTLn1PXXH+pXkJskMVytJ/2jdPQ7ZlIZWhJ+Vw43L3ylmQwW1LhWSso
xyi8WKoV7MOL6aN31zojF4B2rDOP/Fz9tCutdAJmYj0BPx70HKlNcJpH2kt42nlG
lgYTo7Gb2WO4hARswrQvAyOknjor5XThLH+Jz88Cx6OMfBF6KxOs1epjyfWocwl1
S0tokehws7KcM3WtMFOiZNO9YIZ5DnXIWj6oRoePaCLKjLsf+G2XE4FYE6ujJlBG
o5x8iWuNdR2VvsOXdM4rVGF05H1rWUmGl2j0UFIqazZEaRxxrCa9UZhd4mt3aabz
RRqd6e+wx7ahf8zUArbLBWpobYsc2vUNzLGE6+XIle3Zlxp/49Ny4/Hl7hJmvuCc
qUKfa5WahojgnZuTqFFpXrKm/i7J3LnjfYDOQGXmwmdD0Eim/txuabvm2S2LJPD2
eSsrPtqiGInKapqMQjn78azmZ4ptj+GnrGGJI8QdVb9XJHUasEu2/EYpRVx8FgTr
7kcMBcGk2of9ffCfb7h4dfGfMuU+5wzFybmhCyKuLIqocaQmdWKB1H9OvETmcinZ
qlS1h1IUWpagpCZw34kgOuYi+v28JAkUrq6LfwAPAyrFRbI15quwE2z1HZoAH14F
3KsGzWvCgzYM15C+jSvwDlMNmWgGtuxs8nk9EQoEyQTzh+ZmtkqsxkF+rpIl6101
gzXOefcj0yZ6+30gfe5BDL5ks+bp9Ca2/b5+8/CGvsGHWJlrtdlofq+WClWVb/I+
6CTvg88cTrlduq3EdH5JtL1Yyttfv9OhPbQcFczFnEYhR12SVsRNzWk4srKNSStA
Aoe+jX45hNmzPohEd74V2nuj7wgEl2cvHCVxVZF1bPIrucl7O6jJGr9SiNqSY0/e
iaKS2wvKBsxL+JzD2C6gTzXKL0/J02lXaluClNm5MZoQZQvnhaGgmsfkVQn1dhbv
DN7GiQqhBeTIg029mtJIyGA62hTZedO/w9wcLnPrvBb6a+A7EWrraMMCbu97yQz5
ONgdpoRrn0ka9b4e38H3fGpYoQ2CwSlqttOfXVuZE5vGeaJqfIAeWLe7ThVM96zO
FQ3iODywsC23T+lV07ty/g==
`protect END_PROTECTED
