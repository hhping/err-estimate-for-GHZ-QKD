`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G+lqOjA6yFLPPf6QLS9ZcLuvUSfSeoB3QRG56WnFEq0yBcXmBRifDFQeoMJefJUB
M1PHR8JVLlWt/f0Me1Gwj24rsPq/k3fP0pcx6UcBCktSc8DzoYHty5v9Kdz+hTjq
4ZX8m6+5gK6uzRwHgUDj+4Rr/D/2ELOiION8Fzo/Fmnla78zQscrow9M9bMOWT60
kXS9D80I4Fvs1NBCxKjcTouaqQ+RomUKfrqKSY5VxBjbkQjCcv/oLbFlQHc3IoY0
hKYBbk1UkEPrrfeGlGizh91jD9RxEbm9NcMM3xmTfI3r8YDJe3tOfU5afalukGvk
njQSKkaisbcMD+5qbk1wosQH+q3QV31MKsCgEAgB/MEOvpY+Ro2wNJYsKWY3yGVL
4DZrmGCitdku+G9Wd3N0VCVLdmh7fkuXVAt2eK0Jq6RdLUo/NZ++R0pjcIuqnVvn
4khi4sVfbsk7XkdDWFDwQ2o671Y64xWOtiu8ItBDPr+enNKzhz/2TOTNXhO4mw43
Zijqcy1qrzNvJPAIOHM6674Nz8gQRo49sLJTdFXo/uI92nOQV2AeEjIXPjTTY6kr
gbA044sdFChqzZqSnIT2lJIyuM0n2dEv2hG+mCeouECDwhRlDY6euEfgIbP7Chyp
lL5vJjqT0pkEo7cWn2IQkIlqTGF6I+t+Pl38mYjVfY9UUruN29YkTTxGySwD0e1i
aP9oW9EGhTns+FZtxfM0HGIqFin36GXLHb5idLuQ4Y9NaaCcIRbuT52u/KMSgRJn
0WaPnhq6M90TC+EOEPAZOaSXhYR4nvXliXxhUqVVOAop0fLOsZFCbM3c/y/pX06y
+EnWZuD+xK8Oaf3isAiOGw==
`protect END_PROTECTED
