`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/PwnlsyQY4mry8PJCBcLm81fUBT9wYNldt2UTz5+qKAnlHtqUeXflUhapZs77gt
IClCF93jve/9/0e35VZ0emLqERKuDiOed9pRCWHA/tm2hSrnimAmkDsDwYEvOHC+
w9nGWvAj4aqTitkgLlvCeWH3/bKkQ8RhNQXRZOgsEBAS6MdmSN48CyysfQA76BsA
KJn90VAyfMBzYT28tgs6EfCZywSONtpVRDqp2YUdFhzQkQg2SlS1PWtd15jzy77g
gDX7AUuh7Evqe/HPFFuufZeJ90buGoXykWuoYbfNqwmpbIs3SsJRfLxLqqwBH0hT
MTWTyiMYQ7wHYkWOYwfun6ns+sK6TsuuJ0XUdhF3YGGbM1qENRAyYK1JIrQ+3+te
Qtp/Z1ebTUku0bEqIrzEF8vsXPN2QQGTls6icsid9/gDuswl1oXeI4/FVTM3SG3F
BY5yH+tSR0WlI/FpYrry9GgNn4omrYWaGyxq9JmnwTsKQtTgfiOID5Lri/ocBwec
gzZB+QjqU8jH8rqy+568VR8+esQDoMu+Of0Y4PBsVy3deu71OdLodJTXnRysbGGC
hvdZa3ibf3IU6xeO0VzWOxrCrmggrpIDL7XWwO408orShgGZwP2JAiYNYBBigaPG
u/diqrRbcJFslAZzEG7s5zEO8CnN/Da5wzzMlPDx/mkPPtJGxqyJ5pg14+6s53Vv
wEVgr8QmbhO23nrYtsLPVdfbXxfyQ/dyC5GdIA2jHBZMpYuHtvZv0SCp/jgx6bA9
sn6UMrQjrSRiH0VHkJBBgfPZqIuIuttsGUQVa9tFWP4/3nO6muBZ6o5t+DZ1BOnP
OsNyowqYRKQF82VT/X2VFtQdwY8robE2SKApTdZnTrcpOVh8WTuI9p64+Dr7Pd27
O/qwz46fKTNadWsEoF/eaKAJqns8OEkR75m/GHH08FmF8LaDWtzyT+/oIOPUx4nJ
LriOdAZbs29sXmlr8W1rSw9GQWClSHEahQOhrwEyRQlE1jGdRAHFcsyllHF5GAQF
cTQZBUDX1t2zKFXodBmv0NSR3AkCDVUhwzLSC6oBnhE6QeYOYaEJXq8ip9D6jNrz
VSXtjCUZ5fpu629/yqHXlnMdz8RqWVFaXWUN2VM+wEcP1RUAYEktAcv1D/eMho73
961FfFG8hfHh4FnyeZKTbPNKO8djHCrKj39nWYuQGf7pRQVBOmUVhgJlcCf5LQfE
/4NRUWP04osLAajfmGqGhXlATYMjyqAecYMF2kcA8f3RaIKTEdQhwCD3aZEd+egj
gepx4iDkZfbQ5T4n+vC7WsGvgNWERNH81hhhqGOJLSNCnHOiCRWujQNI0PvbJoB8
sFvnqcApWqEJhQb/YawESrRHYRN6eQa3qsZJ8ybf6NMYmHEhXCPdNC6abYhEiJSL
0N0ob90M2HkS5L7P2VC+dnBDcj6evFfM8UdT+46uSH6CDjixAHOAa1P8QKSnYSet
H8soj8XrljM82kf8CfDQAjrQXpikpcLeTm1aIzY54ZE=
`protect END_PROTECTED
