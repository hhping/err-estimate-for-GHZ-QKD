`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1N9U85Jg5UGaDK1B9bCsKK0KUqgpg6cJ2ocT02WGCAaM5AqKpjYFtKvaaT2//cA
WFJ/kMWQPP5EEuqqCR1C4WbCCqg3YALGRHXCOYhZSLeBuWjBmyuTAjTf4qLEQg+N
KURUQKY3Rp2cVlLhhXxohaBgTyxawgyTcw8c4WFq1z9jpEmb5uhHPavHo4yj7tzn
VLpBRbfLLTg4CP9xYOq5FQbjYR2YfrBcdc7J+QQ5pnFeE4/QDp5eHSJf5KGHAg6Y
Y8uAXNSapE5xczyKTMD88+r9w1cYoV5OCcNZ1zb3F9f+4W+4kizfFiV06T2zZYbX
5KImreJy2RbnwRiZD5xedeXfbC2oTWBiNyiWNfJHp43QmP0DtnMQFV6UpRSuZsdg
qYJzlGVIbKCF0/GpN9noD7vyk1UfbG9bV9djWPY1zcnfheVdDcsDwCeHh+pMf46e
0k9VnmUQamxc407IJ0jIyRNvI+8A6JjZH24cH4UrJKrVyakyBDQTPckoBWewwp6n
I1bfyX2G1VNkEG89qASbGPkCMZ5aPW51ws7kgOdOwvHWyQalHu7mq5AGAvYMWazN
vpgIMsrCz/E2u65/+lx6yOIRANKAIGa2x5M+DA1fh5mbqMpwCAAzmiSM/l1FpkhJ
x6MqaVBskfjK3wUdZfm5rpCxFs7YBhsFJvNo0pZl/ZltxNabHEWvzDHjVZGnTmCW
BRLSsND/WrvHnUyOz0xOmpryizkoskqgImPcO9PF2hbKaZ5rOAxdwGbjDuOWvJog
Amgn2RGfkEAaoX7N3n8mEbOeNVKYc7icbP9OoJWhRW0fpUR+Y2ZfRbWRQeiu9imD
hWJI6exTqnlgFNt2ImVTJccwqGpDcfpRAq2+PLeq9mxNXlvSy7cy9lTTZUXjRr8Y
A6ITVCdna3V3IP5v9Z+jJxOeMjcJdG57t9AFLkNY0+itcys3QUo9C0bHjK4JzUwd
gutH+ZDvQJPQhMSoO4l0PBOfcIzK1AjJuMByK3MAQo8oJP2yP/SB4QjX1zWoUZgC
BljmIGLPbrVCbkAvMRyPL0+Idcwp34f8H2K0Mr3kHpVk9Xm93D8Zp+aJ8API2mOw
+/gLet/tM7o8+FPTq2UTib+PzJ8QeXPv2utkGZxib24SMZ9pXydpAF+vDJYi0xfz
2dU+7bZ3xZJ9syodNZvQ0meAstqaMPUaZnoMen3EMwnj7YdHrem0KfuftyRlJahe
NtjrGfrIcxwtZBkUo448HXzJdZl8ZbStmNXz/+pH6krcJjBZbW+CNsuZ+QMpK3Ow
K0uYsBPZw257JVpGJCSLc5d3lmZCnsPvPu8S5oKzuyhmYhIMzDkF47aV1Jp474bE
LvJgR3hywjzainkZoMNc0N1mZQgja4vnnkIthAHV5cpj3rUujrBDbW3XfYp5VyKH
95pai1JWrOTCer6IyPS3MPl24O8uRDTK10MuyJsXfl+sgwcUhRwQ9KPTX830Q6WP
`protect END_PROTECTED
