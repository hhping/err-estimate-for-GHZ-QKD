`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXiXEUJhIBK2RZKPEvkC2zlJ10lUkdkXLyZCKFhxARzq18sC/ixNiP+LHJCWLg+x
poHAnyakT0FB6vZ7Dei0V7kwV6ZSKb61ONr67NVLkev3WU5YQNcgl3KwnVj3ptsP
43NEsiXPXqT9LnI/L1trA/qtqeN6PfjdC2znwOlzqPho81RzHsEoUtw9ZQIZzOTs
PqWWdhdUryYCJpC267YW8hyGkA5noM1lMQ/swEHBFGE875q43VEJPELh6RVwd+1N
KjOM8wSOCM3xRN+ZyuHQgnKCWSGMtoloGB9SVReUGgEnggLRgZASYf05+bQVOOdE
KndGnIMR15dS0nQPk8MqNSBC5YkstcbAv5WWNpm0hNHX8tkAAABhHP865byRf+wf
XfnohZst0a/9TkhQiqG3a/QlE1GbWeUDe/8DQX+PUaJvYNkLzrZGBhb1abu+ERmw
sRVBNnPuSgyRL71QTrC/PpeLHHMPuAbhJjjG+uHZtk5uzO2Z0icfCZejmtssaQvO
rr7hbkDe4VSidU5XGj+fBPzQBTzJRqq25dXXpQpg1W/rIMUyTwUvfx40JurECPfL
F8nDcNUywIRjGyMF2hvmSBw6/2/Oa7LoxDoQ1TZ/stRNl8dJStlLDJ0e5iN5hdCD
AGS3yqcGvA/8ELGwcv+Pdqt21jIG3OKFYc5VNoY7NdQY0rAc93MK6rgnWGyL5AAQ
IduDXzzlN79cV2zklDTurQ0FLOUz5dIgSUm5N4/vTmjD+4XnZwci3wcOV7/1cKEa
/aRjhxlkuiEo+bI2c1a9sGpSMaMAcWSC1xmN8LHXm76wU0nrR4zADoe4Yb4Ngstc
u6rq+j3TerpvmraNr6D3Gu91oNtKkbYYUxyTrQLRqW1wbswMQovuRSAPOioPLRrl
47n+6e6imcRYksi9J2jim2w7gGboUl+0A81m9RR8lpLxXgd8gd4UP3/xbD4zSVOC
27+6HwhqRLqpDwnrm1j6ty8CetHA8KiOvSwGxaSp1kU=
`protect END_PROTECTED
