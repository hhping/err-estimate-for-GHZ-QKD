`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cMM4/eEfLNjMVPBdPBb5ZF+qB2QK4h02rKp15Fs2WVAv8hylEWcxmRBDClimM4q/
X2md8xDt613wAzFDu2r9t4CS+Mm/h+zeC5gebtbMsAJMSPsOJ/nX8bkwmpLmwiW+
FmLZXF45oh63sTKqzMnl4K5Gzw6+VkuM052XtmqOuHsDFf0IfQhcEqP8NwOg/5Lu
DAc7hZarrJXHxhPSO/fQpe+6RJ53E+lk1H3MA2xnmCtdzruCJXmeaDU5ygeV80XA
2rgn1uKc3EYZ56mH1w3mutWSZpeUnM7xek9ox4nhI0OjceU1iofRW4+CBbEmFe2i
bA8+ViK3kJ1bf0kky2kVdlTfMDj9UszGyKrIltmDiIF6yW5b7yki+7X7t8BH/1+x
8b6dR/kOZnwjSeqy4sC9kA==
`protect END_PROTECTED
