`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RE5p/PH3rZDfB00lW8pfe0WzhzvRIl8tEsW4TBLh0RkUaCrax/Mn4lDCe12LLz9j
D+UHnVpafcoCOhWnlS1TSiJqu5oJNL9yE5Z+9dZNuWQ67tdfnCU3/U03WmLTDZ1a
GDFUzi4MB3SqJh07SvyU4K/CH0re8FxOuAgVDnniHjlx1fdGGnUT5CXUJIrp4q61
qEqhQvGd8MIy+lSvhGy1cnPyBKSshdi9xKMhFm3Op3vO7BZ+E8MR6A0ldY3kOaao
MfSFPZqg+i1VjbTm+LGr6IYJ0WiprOqBemxtGYdCOIbfas6CUwpNNA1TfwnlEGtY
/Ge799xm8gm1XIObOpo6lgO+mBymNdpPpYMs8PRzgZv/SneGTovFwJltAlnfqYg2
klfffmwCZ1YFJK4Jas95xSfTVzDQCDtsEG8Q5nm3oTJktAT/0xs4HcHf1Qp0Cvy/
qy/jXw68e9i1QV/JOROAi71pTBm5GNcHZtDRMagokDirX0U6/kXaw3lgdpfDeQ6l
1jkVuQXx8+Y7RUrLKtqqiq0Dpob1DTEET3IT5NJxb4/bD7+22JgwKX/yxa9dO9vO
jYE56+IdkzX6iliv4zb0tuYj9IyUHBXPsetFDhiMNid5JaSITTtl3Iko9geAQt1C
8wN2yhb6btgZFYYnptKUKYSbC+qlZ9J2MAsrf1zgfqr422IBsNTWrFTK8xCBLqB/
Q+oEQDLHsM7TqfsCNTLqK9TNmbC1y7A+5HJ86Zz7Uw6hdfXir6VKzsDc9XKpo1sA
W2MtCTy12Y7tt07V9e/saDi3CQBdba6vrUUuULc7FqB2cYjvYAtF3Eaqd3ptvsYH
+MaNlQvVXFT2N1MceZAkEwSzDOkR2Acwnf+BQ5018ZSpc0IxTmSfanwMEItufE32
9mGaRiS90udOF/MGxXzLfRF6rfnaVplfK0ePypUBHMGpox7jjZlJiKb976qLl6NW
duLEZsJGEWeY7cwr0u3YApc+HvbrnFyo6m9ScmjK1zDxSm11N1z5Xej18m4bXxn9
WtxN/1bWKpq50bDEguMsOzfXk1JeSXQ6LJzqSD5BT9qvIzRWFxGHE4Tq4fyVamaD
1/YHgM8MtYp6XFfHZE0rOxDqXgzUwfv6rm7swogaVmwX6Z/RqcjS4iiajKuoDb+M
J1QZ3djMpR77ctKnBK/IlR8uceuIDLe85LHym6PtgziuaIvQQGDpfeAulTUa50N4
nXorqxQDS3zUfP0yukOpHwUoEVdP003X4zsOC7E6TyaEA39o8uBSB5iBUB8bdHZL
W6FO6CRUKi5n9w2IX+BQz8IbtZEgBCpvNmFnNh+N4g9+rjvEa4gGgnIta2R+QEdV
bKJE9gjnuov4hv6B2YHZi4aNt/udc17IqI363N3ms0tsR3y1LdrMhbfcUXYusPSh
RVzGpmXFLbvpuvSKAtsXwRXikQvdMlYlGubfV2moGInmiFi2B5AoWaBML471IYr0
NvMwf0DLZEc0jmVDP+Qo3kUMyBYPSYxBY4PgmrAKImCcb8csKN0m/LJjCBf1Mxmf
BQh9+zhbLNrWAvf773RYtDoVVz3hPnPbO9uutRIz37A=
`protect END_PROTECTED
