`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xc3FFQcI0q/C0LH51lGrwkg+CV/8aNNDjHA2hgciAZb0pr0HckbZFIBW5txWWU6p
oOXj7cn7OWA9tlWUvP8AsvEueLBGMRVLzSRwVbLtxaDjVmOV4gUSUSQi59hro5oU
TQwbrjJv4FBBolyAjQmIec3WMEj47lxr3Jdp6E237jRBL9G3g0gcN65l7LES5x6P
gbVhS9A2TTi+JTaH2rbwqfME3VHNZJ+bky4zgDsdLpftMfCokQ0iIi2E4ZbJ++hM
RDHV65xbMKbUIhnXVEr+6h7bgMNnSwMQlVb5xyN9AAVk/fNUDcSL9WUaYAUT9Rwn
Ju1MAcWF2WNzIaWePuCzXwop1E0EsRFloDACeqkzDQOKg2aUm1GQnVLV+jeLtrF4
8sf+vuegoppP9R0QfMc+SqcjLlpH6YzGnAN4mxAG+lTu9tKdRoD1+f5QnU/7PR4Z
B4ei4ZGl/JTT3r+U0LivChQCc9Kd3R0Pdiy2vCH44Gfakbydl0HSOnPb0Z/4pDUu
0dh9n02EZOTU+sf/dZ0YbpknFQqQV6FaVHJtFLT8eUpwvhekEh6i7Gic5hmr3Gax
IZlxZO+DPjMhb/0hl7ScGRTAWeadsyXPsPsWIGDMgbvo2ErYlCVmmvIce9HwdEeT
Bj6MT2UkN9/w3eR/iaKQviO6uGJVkC5kGv9TJ0zMf9RKg0kdpmEaIhymO1Jxzhwz
YK8HMAO7lHEpMgoft+beYodHws+Fr7+IdxM9hxGMJl/s6qTWr/CLw0PivSuLRz7c
ZUCYIm2F68wogrGq/Yq1nTOCY314ZjicEeSEOH9nlD4EsZhKJnG904puOV0F81ka
stTmdA3JurzsRUR07t5UaoV++LeliZJQl/7rC1yEDJdX/umFuzjWJA7fZj8eRYYg
i7cSdWQDq5VouR9esXtbTunSkI8bjJ/YiDDiOwt7U48WsLA6vi/HFs4rvRdipCNN
tfRNC9lDxKnG/dVoIrVTApxqNM4IYAB2Kak6Kh/03pP15KR1IQDB51QVF+L/CySg
MjhhPe7z7h56AmvNNCDlcV58ei7uOCMez9hgiQ4VxKAn4x1M4jFtlTwpcMxnkmXK
rUPQN0IJv1e28hOPN+YQs6rEx8UKtBKawtKw5IVkHdY8QCBRJrYEBeQ76JrL19eg
010tBe8Kb6zbSy+iqUJ4sOPhphAXJV21+5txupJY3Z4aXH76r0XMR7aUdOyygS1U
i081RtbEsmM5eaFPhcG5F/gaZyQri8/c18HCRGABSpifJkbuSR0mYLNm8ALECsVD
Tubhs1HDvicp4z9pC4iQw9yYoj9GPUREPvOSY0KGuOQgRtSt5MLeCWJtVgI692L7
STIQJ+p4O7s9yKJxcR3fH8Cl0bdSAwNFEe4e4cuEx+C37tHqEatEDQgx5yiTJSoX
L7L/Z06p+3edXnlg4ecVYggbujsVtLMSGwnwcDh916xZYZfqGUgw8Wl4zUNTA6Z3
VZ4lhAn+8q8m/Ipggj+AQ8LaG/kJupMKIM7ZlvC/qwh5hzutglduPwShmJSgI6t9
wdpPhv00A/r9OA+nlFHSwADvmTU2ilw1MvBmQXhOn2VyuAoCLIigJUsATLYZbSy7
Hzyr3UEDSb4JGO42eaOxN0njUsOWW6nbn1DHqaIy+2o1dqby5uvMPSJnSD1spOhi
NaSAEELKTkHcAQ5q9pkiqpRVubBkJrajpCQqF10qexp70uaT6ZGnlcYSnMXWwbZV
67bQiodii2kW2F4dBzWyTkW27aQunYv68ys3WZUnKX9ZXxb1O+aWjytlBaAeMHmg
E6DXry2Rg6l29t6Zpw4w1ze94QqY2CHE151BwHrw6o4fzSXmzOI34u8qU63+ce/l
ahcbc7EtNNA5A2cok/r6dA5F8SNWDXjbf/MOvyYUqIQaeirdUAu2v4FcxwXGvuj1
z+ffujWvtZWa0nPYSVSruKRdtGG8WTtffR7CqLuaVTFV2C6P7C7yormYRcl5UcV6
hq5lewomEqdkMbJ57jyAXozuIIwKgFfiUxRdU5ISLtxpi/pf03yGBBFQya6ns2G4
liQRtpk3mIftcHKeRd5/d608U2lIooavoBwGM1i2johQvWdMkv5q66aZuWNXIiyq
4cov0wgD/V7DlxxGV30BcyFbJlN5+8Cv8SeebwwqCoek/oEJp2iES05kvx1jEUhs
UEprJJ1F7pQSJFEugBXdXcsJ+65ZY+4+McuSqZc+DXoBWmo0FC72omnIeksx+0zZ
HTLXkk92yXKykgL0qV3u2fLI73Hu3gnFzXKxE1SHkkD48BBc0ra7msTcSmD+gKiP
yjlosK+R1pUGZBlQDDZR0Z/oWMNWVQDOHKXZ80TRjOGa6Ea1Zo0fxAhEl96uUCHk
9KZa6P8f5mKnuJtWGhqUVk+QTDichyBsnEFMFPXUFxn+k4UZWUOj1fDRjFRXD/Ew
`protect END_PROTECTED
