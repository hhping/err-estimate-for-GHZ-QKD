`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0s9qUgO253sNpK2gV95h6AJRM4FLDCsbMllcqkc7aIgdE/6PdT3AxDV+tL+23SoW
xVPBecyluqrughmp1gxgK5ezMdyr2WACDUoIgY+9iL8PtF4s+P3hNrludk2ufd8d
zx3rCy2rUTQEK1qgzAeGwedZtPRbplwbeJQCoDJuzMyQtPInLsl2MYnzR21Y4d/B
kZqYTYNyNW6VM3oIeoLH/vtsQVp3gfPyo4Th0Q1Wgqvx8cBypBC/eiSoKMKxOudp
pkfR+verN2wLOOFMG8APMCkPsnHVrCfzVlMprLbqM3QtY3QzN3zHRlMdwIDmbzuE
PXyoHH9ofUhSwRbX7/GZ1HxQHXQrq36i6tcl9hSH5n4VsfH/hxcfdDOMMlm9nzF6
H8xL+dYAlAaCjakwSINJzi712RHZabuCOqQz8yPDVVzNPGIYBDhM2wUy78gUgOiZ
gVU1H8U0rbch1rFuG12N8sPAREz+CNZcl/o2aKi2pXDvb3vbd/bvkl2ApA+hXR3F
GUT5ilM2m1Z4kq+kCXw2QWVb0VRNy+SWGYXw7CvZojEMXm3Piq7Mz0Rv81cN7n6h
ZSI6i9XZ4oRVzg3JwgjQ/0MoihCAZymxqXuXxbZjuovjOHwsADLwbtc5eSU6uaDN
ALdDA4MuOkEjFrpAcuqPO8nHZWY+rhVmJ9hMZP6LQ+U=
`protect END_PROTECTED
