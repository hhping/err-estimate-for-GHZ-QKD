library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_10g_tx_pcs is
    generic(
        enable_debug_info: string  := "true";
        advanced_user_mode: string  := "disable";
        bitslip_en      : string  := "bitslip_dis";
        bonding_dft_en  : string  := "dft_dis";
        bonding_dft_val : string  := "dft_0";
        comp_cnt        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        compin_sel      : string  := "compin_master";
        crcgen_bypass   : string  := "crcgen_bypass_dis";
        crcgen_clken    : string  := "crcgen_clk_dis";
        crcgen_err      : string  := "crcgen_err_dis";
        crcgen_inv      : string  := "crcgen_inv_dis";
        ctrl_bit_reverse: string  := "ctrl_bit_reverse_dis";
        ctrl_plane_bonding: string  := "individual";
        data_bit_reverse: string  := "data_bit_reverse_dis";
        dft_clk_out_sel : string  := "tx_master_clk";
        dispgen_bypass  : string  := "dispgen_bypass_dis";
        dispgen_clken   : string  := "dispgen_clk_dis";
        dispgen_err     : string  := "dispgen_err_dis";
        dispgen_pipeln  : string  := "dispgen_pipeln_dis";
        distdwn_bypass_pipeln: string  := "distdwn_bypass_pipeln_dis";
        distdwn_master  : string  := "distdwn_master_en";
        distup_bypass_pipeln: string  := "distup_bypass_pipeln_dis";
        distup_master   : string  := "distup_master_en";
        dv_bond         : string  := "dv_bond_dis";
        empty_flag_type : string  := "empty_rd_side";
        enc64b66b_txsm_clken: string  := "enc64b66b_txsm_clk_dis";
        enc_64b66b_txsm_bypass: string  := "enc_64b66b_txsm_bypass_dis";
        fastpath        : string  := "fastpath_dis";
        fec_clken       : string  := "fec_clk_dis";
        fec_enable      : string  := "fec_dis";
        fifo_double_write: string  := "fifo_double_write_dis";
        fifo_reg_fast   : string  := "fifo_reg_fast_dis";
        fifo_stop_rd    : string  := "n_rd_empty";
        fifo_stop_wr    : string  := "n_wr_full";
        frmgen_burst    : string  := "frmgen_burst_dis";
        frmgen_bypass   : string  := "frmgen_bypass_dis";
        frmgen_clken    : string  := "frmgen_clk_dis";
        frmgen_mfrm_length: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        frmgen_pipeln   : string  := "frmgen_pipeln_dis";
        frmgen_pyld_ins : string  := "frmgen_pyld_ins_dis";
        frmgen_wordslip : string  := "frmgen_wordslip_dis";
        full_flag_type  : string  := "full_wr_side";
        gb_pipeln_bypass: string  := "enable";
        gb_tx_idwidth   : string  := "width_50";
        gb_tx_odwidth   : string  := "width_32";
        gbred_clken     : string  := "gbred_clk_dis";
        indv            : string  := "indv_en";
        low_latency_en  : string  := "enable";
        master_clk_sel  : string  := "master_tx_pma_clk";
        pempty_flag_type: string  := "pempty_rd_side";
        pfull_flag_type : string  := "pfull_wr_side";
        phcomp_rd_del   : string  := "phcomp_rd_del2";
        pld_if_type     : string  := "fifo";
        prot_mode       : string  := "disable_mode";
        pseudo_random   : string  := "all_0";
        pseudo_seed_a   : vl_logic_vector(0 to 57) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        pseudo_seed_b   : vl_logic_vector(0 to 57) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        random_disp     : string  := "disable";
        rdfifo_clken    : string  := "rdfifo_clk_dis";
        reconfig_settings: string  := "{}";
        scrm_bypass     : string  := "scrm_bypass_dis";
        scrm_clken      : string  := "scrm_clk_dis";
        scrm_mode       : string  := "async";
        scrm_pipeln     : string  := "enable";
        sh_err          : string  := "sh_err_dis";
        silicon_rev     : string  := "20nm5es";
        sop_mark        : string  := "sop_mark_dis";
        stretch_num_stages: string  := "zero_stage";
        sup_mode        : string  := "user_mode";
        test_mode       : string  := "test_off";
        tx_scrm_err     : string  := "scrm_err_dis";
        tx_scrm_width   : string  := "bit64";
        tx_sh_location  : string  := "lsb";
        tx_sm_bypass    : string  := "tx_sm_bypass_dis";
        tx_sm_pipeln    : string  := "tx_sm_pipeln_dis";
        tx_testbus_sel  : string  := "crc32_gen_testbus1";
        txfifo_empty    : string  := "empty_default";
        txfifo_full     : string  := "full_default";
        txfifo_mode     : string  := "phase_comp";
        txfifo_pempty   : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        txfifo_pfull    : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        wr_clk_sel      : string  := "wr_tx_pma_clk";
        wrfifo_clken    : string  := "wrfifo_clk_dis"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        distdwn_in_dv   : in     vl_logic;
        distdwn_in_rden : in     vl_logic;
        distdwn_in_wren : in     vl_logic;
        distup_in_dv    : in     vl_logic;
        distup_in_rden  : in     vl_logic;
        distup_in_wren  : in     vl_logic;
        krfec_refclk_dig: in     vl_logic;
        r_tx_diag_word  : in     vl_logic_vector(63 downto 0);
        r_tx_scrm_word  : in     vl_logic_vector(63 downto 0);
        r_tx_skip_word  : in     vl_logic_vector(63 downto 0);
        r_tx_sync_word  : in     vl_logic_vector(63 downto 0);
        refclk_dig      : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        tx_bitslip      : in     vl_logic_vector(6 downto 0);
        tx_burst_en     : in     vl_logic;
        tx_control      : in     vl_logic_vector(17 downto 0);
        tx_control_reg  : in     vl_logic_vector(8 downto 0);
        tx_data         : in     vl_logic_vector(127 downto 0);
        tx_data_in_krfec: in     vl_logic_vector(63 downto 0);
        tx_data_reg     : in     vl_logic_vector(63 downto 0);
        tx_data_valid   : in     vl_logic;
        tx_data_valid_reg: in     vl_logic;
        tx_diag_status  : in     vl_logic_vector(1 downto 0);
        tx_fifo_rd_data : in     vl_logic_vector(72 downto 0);
        tx_pld_clk      : in     vl_logic;
        tx_pld_rst_n    : in     vl_logic;
        tx_pma_clk      : in     vl_logic;
        tx_wordslip     : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        pld_10g_krfec_tx_frame_10g_reg: out    vl_logic;
        pld_10g_krfec_tx_pld_rst_n_fifo: out    vl_logic;
        pld_10g_krfec_tx_pld_rst_n_reg: out    vl_logic;
        pld_10g_tx_bitslip_reg: out    vl_logic;
        pld_10g_tx_burst_en_exe_reg: out    vl_logic;
        pld_10g_tx_data_valid_10g_reg: out    vl_logic;
        pld_10g_tx_data_valid_fifo: out    vl_logic;
        pld_10g_tx_data_valid_reg: out    vl_logic;
        pld_10g_tx_diag_status_reg: out    vl_logic;
        pld_10g_tx_empty_reg: out    vl_logic;
        pld_10g_tx_fifo_num_reg: out    vl_logic;
        pld_10g_tx_full_fifo: out    vl_logic;
        pld_10g_tx_full_reg: out    vl_logic;
        pld_10g_tx_pempty_reg: out    vl_logic;
        pld_10g_tx_pfull_fifo: out    vl_logic;
        pld_10g_tx_wordslip_exe_reg: out    vl_logic;
        pld_10g_tx_wordslip_reg: out    vl_logic;
        pld_pcs_tx_clk_out_10g_wire: out    vl_logic;
        pld_tx_burst_en_reg: out    vl_logic;
        pld_tx_control_lo_10g_reg: out    vl_logic;
        pld_tx_data_10g_fifo: out    vl_logic;
        pld_tx_data_lo_10g_reg: out    vl_logic;
        distdwn_out_dv  : out    vl_logic;
        distdwn_out_rden: out    vl_logic;
        distdwn_out_wren: out    vl_logic;
        distup_out_dv   : out    vl_logic;
        distup_out_rden : out    vl_logic;
        distup_out_wren : out    vl_logic;
        tx_burst_en_exe : out    vl_logic;
        tx_clk_out      : out    vl_logic;
        tx_clk_out_pld_if: out    vl_logic;
        tx_clk_out_pma_if: out    vl_logic;
        tx_control_out_krfec: out    vl_logic_vector(8 downto 0);
        tx_data_out_krfec: out    vl_logic_vector(63 downto 0);
        tx_data_valid_out_krfec: out    vl_logic;
        tx_dft_clk_out  : out    vl_logic;
        tx_empty        : out    vl_logic;
        tx_fec_clk      : out    vl_logic;
        tx_fifo_num     : out    vl_logic_vector(3 downto 0);
        tx_fifo_rd_ptr  : out    vl_logic_vector(15 downto 0);
        tx_fifo_wr_clk  : out    vl_logic;
        tx_fifo_wr_data : out    vl_logic_vector(72 downto 0);
        tx_fifo_wr_data_dw: out    vl_logic_vector(72 downto 0);
        tx_fifo_wr_en   : out    vl_logic;
        tx_fifo_wr_ptr  : out    vl_logic_vector(15 downto 0);
        tx_fifo_wr_rst_n: out    vl_logic;
        tx_frame        : out    vl_logic;
        tx_full         : out    vl_logic;
        tx_master_clk   : out    vl_logic;
        tx_master_clk_rst_n: out    vl_logic;
        tx_pempty       : out    vl_logic;
        tx_pfull        : out    vl_logic;
        tx_pma_data     : out    vl_logic_vector(63 downto 0);
        tx_pma_gating_val: out    vl_logic_vector(63 downto 0);
        tx_test_data    : out    vl_logic_vector(19 downto 0);
        tx_wordslip_exe : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of advanced_user_mode : constant is 1;
    attribute mti_svvh_generic_type of bitslip_en : constant is 1;
    attribute mti_svvh_generic_type of bonding_dft_en : constant is 1;
    attribute mti_svvh_generic_type of bonding_dft_val : constant is 1;
    attribute mti_svvh_generic_type of comp_cnt : constant is 1;
    attribute mti_svvh_generic_type of compin_sel : constant is 1;
    attribute mti_svvh_generic_type of crcgen_bypass : constant is 1;
    attribute mti_svvh_generic_type of crcgen_clken : constant is 1;
    attribute mti_svvh_generic_type of crcgen_err : constant is 1;
    attribute mti_svvh_generic_type of crcgen_inv : constant is 1;
    attribute mti_svvh_generic_type of ctrl_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding : constant is 1;
    attribute mti_svvh_generic_type of data_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of dft_clk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of dispgen_bypass : constant is 1;
    attribute mti_svvh_generic_type of dispgen_clken : constant is 1;
    attribute mti_svvh_generic_type of dispgen_err : constant is 1;
    attribute mti_svvh_generic_type of dispgen_pipeln : constant is 1;
    attribute mti_svvh_generic_type of distdwn_bypass_pipeln : constant is 1;
    attribute mti_svvh_generic_type of distdwn_master : constant is 1;
    attribute mti_svvh_generic_type of distup_bypass_pipeln : constant is 1;
    attribute mti_svvh_generic_type of distup_master : constant is 1;
    attribute mti_svvh_generic_type of dv_bond : constant is 1;
    attribute mti_svvh_generic_type of empty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of enc64b66b_txsm_clken : constant is 1;
    attribute mti_svvh_generic_type of enc_64b66b_txsm_bypass : constant is 1;
    attribute mti_svvh_generic_type of fastpath : constant is 1;
    attribute mti_svvh_generic_type of fec_clken : constant is 1;
    attribute mti_svvh_generic_type of fec_enable : constant is 1;
    attribute mti_svvh_generic_type of fifo_double_write : constant is 1;
    attribute mti_svvh_generic_type of fifo_reg_fast : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_rd : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_wr : constant is 1;
    attribute mti_svvh_generic_type of frmgen_burst : constant is 1;
    attribute mti_svvh_generic_type of frmgen_bypass : constant is 1;
    attribute mti_svvh_generic_type of frmgen_clken : constant is 1;
    attribute mti_svvh_generic_type of frmgen_mfrm_length : constant is 1;
    attribute mti_svvh_generic_type of frmgen_pipeln : constant is 1;
    attribute mti_svvh_generic_type of frmgen_pyld_ins : constant is 1;
    attribute mti_svvh_generic_type of frmgen_wordslip : constant is 1;
    attribute mti_svvh_generic_type of full_flag_type : constant is 1;
    attribute mti_svvh_generic_type of gb_pipeln_bypass : constant is 1;
    attribute mti_svvh_generic_type of gb_tx_idwidth : constant is 1;
    attribute mti_svvh_generic_type of gb_tx_odwidth : constant is 1;
    attribute mti_svvh_generic_type of gbred_clken : constant is 1;
    attribute mti_svvh_generic_type of indv : constant is 1;
    attribute mti_svvh_generic_type of low_latency_en : constant is 1;
    attribute mti_svvh_generic_type of master_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pempty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of pfull_flag_type : constant is 1;
    attribute mti_svvh_generic_type of phcomp_rd_del : constant is 1;
    attribute mti_svvh_generic_type of pld_if_type : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of pseudo_random : constant is 1;
    attribute mti_svvh_generic_type of pseudo_seed_a : constant is 1;
    attribute mti_svvh_generic_type of pseudo_seed_b : constant is 1;
    attribute mti_svvh_generic_type of random_disp : constant is 1;
    attribute mti_svvh_generic_type of rdfifo_clken : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of scrm_bypass : constant is 1;
    attribute mti_svvh_generic_type of scrm_clken : constant is 1;
    attribute mti_svvh_generic_type of scrm_mode : constant is 1;
    attribute mti_svvh_generic_type of scrm_pipeln : constant is 1;
    attribute mti_svvh_generic_type of sh_err : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sop_mark : constant is 1;
    attribute mti_svvh_generic_type of stretch_num_stages : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of test_mode : constant is 1;
    attribute mti_svvh_generic_type of tx_scrm_err : constant is 1;
    attribute mti_svvh_generic_type of tx_scrm_width : constant is 1;
    attribute mti_svvh_generic_type of tx_sh_location : constant is 1;
    attribute mti_svvh_generic_type of tx_sm_bypass : constant is 1;
    attribute mti_svvh_generic_type of tx_sm_pipeln : constant is 1;
    attribute mti_svvh_generic_type of tx_testbus_sel : constant is 1;
    attribute mti_svvh_generic_type of txfifo_empty : constant is 1;
    attribute mti_svvh_generic_type of txfifo_full : constant is 1;
    attribute mti_svvh_generic_type of txfifo_mode : constant is 1;
    attribute mti_svvh_generic_type of txfifo_pempty : constant is 1;
    attribute mti_svvh_generic_type of txfifo_pfull : constant is 1;
    attribute mti_svvh_generic_type of wr_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of wrfifo_clken : constant is 1;
end twentynm_hssi_10g_tx_pcs;
