`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qoEhcToMwt2wDQXPSbxwp53FlmQmyi50tzHHq2A+DaJaOhHqlAuAvv18v/pghSDv
BBPi+lUD46fXO9Ku0W6DflEoByOqyc2ohMN86PsJdSbdQl2Z3teMrte4loLDk+Iv
IwAUlpmEX1MjM57b6n5l0z3iwfA7R+wSzrvDe1EwZhUy8RtmtBnt5MDzEQy3PXTo
FXr08hgpuYR97sHi7JbWB5GHwWZE4A7fhwuwAE/tyOof6wxcx04pkTlyx0qV7eh1
6HXCOBoTDopDicHrgtUnGKDiT/sz5KE6jNxUrKLEqlCjpDJY/Ry+jhK12Acug5X7
Jr0FILQGJhrthA/37J/jp66Gw+mwEOasTUdVHceE1Va7uQ2hgoTbvEj3jTMQzbKb
g/LunRzIlTHFY46sDjowD0vLWLeWHKkheXAYqEqfxMwnNFem5ezSt80hLyOT4iQQ
6nxJUhAY+io/mMzdTBIx3h/5kFxTDyC6lsZWSHHzJ04tve2XpoK7xcNCjps+Wf1U
ZeByzrbsrFvv/moSjm9V118BGhelBNQxmyErpHQztvwb1lm+8lOQXY8luiQjDucJ
dMx2T4kYzkCwqKaSEfsvh78PSy9g0PHdtnBowN3el0JvUSys6cx+XG+GE76D4nmc
dO9tRAtIOrW8NFB1bTiNxgDURDjUy8oo20enu4/T9/FgPOT/tm4ofqSGszamti7s
1u6+83GJ84EW5zxx9sy+x3CXVNGw5GOy90Xg+X/zD11xbGPw/18e2B9KXDuViFTP
W8Ug4Hh6a/YFmXd3iAhtNCavYqSCED45tOobXOGO1RyNc2OBBcKCCfRt/8zFcp5E
YxS3XSpi5JNOvvP3KXPspWLB7qIHt4A94E0WGSK5lBB2sFyu55pkp+V6Ndw2yu5X
VL43k2r/wWpJEsUoFdFkvw4FMOp3qZzbMLzxe863I29aMa9P2WE7gr2uBULeDO0h
9Q2M1+WaSxqP2oWUKdMsg+heEzqqoJdUB+4ALg93weDzYrcPgsMWABEWjGtdl3bg
aQRYfoRegl7YsE83jY+Q/Oqcf02AElNPMsfr4Ce5GcR/NoSR4THOKvT0ahsanil8
yP9g0CuuRNF4AyTRrCun/0IUB96C57BFvoqnicAJ/4nkkA0nykWZJeK7aLORzT/F
YOIup4C40aN1YtsAXlqY7yShTiahZacfpFMzZgkWVLQwQq2xDh4ho8nAi/3OLw9n
2P+LMeBPNdoztAjhCK7WqHrnSCvhFNtsa3j76xEc+hBH21xuokVeCRKxMA+PPqNA
NfQgmXmnqgVjq6O0ff7atn3egwTdG8ISYAcLvErnceSupcwQ73wEJ6gS7ITmntII
n4BW1DBw6/3MTZDWMLZdx5koKoWvHR9w1JnqBOp6IDsTkFaWxsTc3HKWw631AjwD
Qj3C4UpMMqTdapzGBcDjyBSxt4rblIa1b1u7qurj++AS4Xtcz7obzLYFVBU4GX5x
6MjI84noNwOueYXF9EgGXRCVdUinaSo54JFrhq6jgP0ELFv86Z5VfY2xSPM2WTKR
+R+4N7SdKHmyIwVLWmkXxw==
`protect END_PROTECTED
