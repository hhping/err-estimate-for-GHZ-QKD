`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bysXPo/PFLN9o/dTWw1oRH0SP3gaTDONl3wTkpKPDRy63bWzwPjEoE60v+eCZ0Zu
XVq6foVd53LVd+5h4ALOrbWSxIo34uFBWX9IwW4Dk2U1DGOTXW1Yxu12H0JS4mH/
cpHvyqEKozxkOos5giEUq/buOJKZ2vd/RQNK38fKCLsNJDZi+scCUGCEaT4OU9R/
4dApo3U9/KuDO1I5MJxNqTRCnGa+HZdcaK1crFPwKIooUJZHknqc+ueU7NBagWnT
a8fIimP/BPpaxqqdRNrWoGAsYlXuKObNbFqKymtbU7PkCfeWtmMn/v+iJshLUzRQ
aUEzD8+bXM6HV9HjZBADXeh8wVp54ekCmSoybT9LKr4mEwk7WuMHX3Ym3VFal0cU
ydHKuhY5pvmlt+X4OEdFAPu565lxTJXByuvAU73fFpsxiH1VCHgDH6WRAUds2rjV
iYLkv0+VaY2UD4N8he8cgv3bHiF1ljr4VixQFKgubfny/3YzJBHCrX6nTEoVuXav
+4mvth9ykyH+BhwlpQSfMltNK8iQezThgJyHH1TD3LsHcAa9KSZi8XljJm44U6Tv
NW3r1I53Y3NkUqBNlzUUj90hkAPPQ8uB1EIIxQIBIqexf8jYPPB7Hjz/Xfpw53bJ
gYcucLflwhzSFWBQAe/Vglt3KXEiYu87q7eG1S0wFBOk7FRunsI8xj6m9MEw7n+u
mkmHukkPnb/sL7Tcu2dxZrvIdbAb3LtXq6UDa/eG5ulKEGOUXAfYx7dknIGy4SYm
NauQyrJZFLXgkDOpoTyMDiCg8iPXQlN4VPGSir1U4Ipiou7nmEfUmjL6Z8bn/vzG
poW3pJdDhrgLE2GPwVFVCKTQQPGMIZd1654e6qePQtBl5lVw1hs80XHhYNoxie/a
AioH3lrIwO4cpbAA66CX//SEffNPItkuEnvICCaQUbw5OWgtQLZXKKABWYWo1LMd
VlJguVbJBrnSaByDqRPlR/OZPEOCGXOzy6FqEsT9t/I4NfAMXBlYLQvHCaX993U/
hEpQ+ZykVaCz9PVgYg2en6YDn5zUNmMCUAmLDqbnqFo+WPxP0H2ww8dlCjNgI1LK
00k/Z1kcs7A9GM1x+TMqdTYeOh0gcindLNE67V+y8lfRucmLUXMYVSfOV0zjLPrO
A083VuQ1BnQtr/KnV9vcNThaOwze+EpgxbfbfwjXpkDDMbyc7M3rArWzsc0vhjKP
mBzpThcXYlpP3zLItG/nMqseu07hra2337Pd9j5NvMFFEiF8eCVUWR7A6+4RXhaU
`protect END_PROTECTED
