`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hB7jZzQfgGK+wRURtt39ZiN057/3npG9Z0Cm+67tQx7VnRPn3X0uWp7ay38wP7Zt
R6ueLJQP4orcIvk07fuATdzmba4KEhABzd5dyowz62gXJaT6+EKJlbHllnaSRkpp
u1F+sWaIX/C0eDmrxmVm+JnKvRKJWTMnr1VZvfrlyo6ersz+y3F3ZX6jOutakDHy
y3C6xDc0lclE//wDtehO1vgVnLx97biGqHfFIMh+XwIUuuzDy1dQ2P0U530xNV2A
n9AcvgiZ0HdX1Sq9ORccpbCzT0A9m9pOLdgwSuf6cBIz2HAnqUq0PEQxULzj6eUc
wv2hk8KEgPX42JBduBNxAcIn9dPn7+WhPA2uWK9eV373gsG0NAWmu0wp8cTsEyoW
oYXe6M5Rtn7rdIuyPMb/S5RXjNQ8K9yAP2y8vFmCqiaCVwRXr1kwtRtCNQQypjwU
Cl8y718M3RAjniHGIAmEXnEqXsUrvULTql/szRngblo5NJk6qTEO86iaPZhkgyA9
279E1pjaHhDIdqBpz937xQgfsn+K614PceXOzD3or7NsU/KifmXLB3Tcr0bFdSqk
yBIe0QBuqyDCMvniHr5O1VB7s3ekNLGwJs6mk8MPNYtFGSSVpKXV1z7sruy9CILU
PjNnXBmMjEESNylyfTBrsfC+2hv6njcwmAQbEzV4okg=
`protect END_PROTECTED
