`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wk8CuPwrPz6wUBUXDqeKIHY1t+MmoJnmkkhnGyISGRTEfboAPZduGbwDy/uh+BXu
MLkkPUwkwsEujYAOCAxzUnRZeMK6BmwwTc0PyuLAEUo+AMUG+nBXAsa4uTZulitv
7v8NAaeNYnaiPP2gnEVLUjUk97g4C0fTEqn0c/0yjsI/4t3dYAvh8eOxGGAHPclx
wkVYFyI/yXYKjG7p1TlBxJ5166UCrADPZudBL0P3XZIr+Ww/LRmOEbjqvi6pPOXO
hyzmwx97IX5VsdG86j+tjNZ6+1ipvadgIwBluV51n4ViZQWKJn3t1M5VnOO72AgG
YvN8rk//b7Dsyq/N4ktGZlBJI36IwuFg/VvVAhfSY81CH4qmmUaw++A3g0QtY4im
a/YsgTUseuZM8Mfq9b34F/FtfxzTiwMslz53jdYqqSRlqUD+OrcAVQhnMRTSqazT
emsUiSXh6n5felKbGr49EsfSLxPiyABxfI20nvjQPrHSwtENUtCAzGRXPrRfuwcC
Dt+86XWg4/0BtSw8Id8PsbH1escPnQrSFv0WSNUA7HG81zfkFAhV1a/FuCuuwmBJ
7X/kvhDbbwewxlB5jO5iASK8hw89b4cOo84be5sieHlOR0trrMJofdfG68EAX3Wb
`protect END_PROTECTED
