`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aiAEwb3XLe8ogsp7LMYKHuHRkD/oJTYIDwGLqgkfuB6mg1eKraa2Mw+RnyJKEsR
MEbnlJoQorZEErfDuIwwEceOIiNp1tPe3lFE800CivZsvyVWCTDEzwFy+qvxrVi8
t6Jrp3qNIsb0+X49cFvdr+rdV9HFrn5k92mES5LSp7EvdewAMiaAjPb/Phgs0dRw
CpiOiwz8ZjKaItq2+Qq+ezWXD++bongTzqWRyBJ7fvIw/gVHNBsfgA0+7PiSvDur
zgUajOxy30XTSiFoOOGUQYhJlrewaWLDPK+JR85N3mmLtl8Y4clE5LYmj+cG70H/
vkq76Ye/74folsWoMTNzJRefFQ3Ysqwlz1flZVAktfrp71XiSD/4jpTuUiQ9SPcH
KQgIZdoCd26YaP6ubP7B755pxCK8S6ApnAll+gAriQlF2QGG8fAf4EzChW4yGqvZ
GxlI4NivJAQlzhEu8vOEGcZ7JP4S0YIwgWx/f4N5M7OsxZpSVmZid1lCriM/hZTI
ku3L0JCZKwzFNm0Lx+E82fFvjnbNjkTMN48tUjtV3cjM8s8rqssZ9aJwwiVQ4k9M
43unBrQu6kjWBM8C1VKf8/KFptXUC5x2iOqQ+qkEjktLK/7tFwVFQVmlRw7RykIU
ZN27IztoJfG/3HSKzomB5Kth9uRf0FgvAmbfXe40ZNuaSRDf/BkyIhxTRnRyiDYS
J/FZXS7lgsV7xbMIiPkjffJihypgkonwl2gMuRnRDw51C8bXvAUGNkeQ6tbNrRQR
AcHZEgLHNkmcYHV80QEdOlbzKkXhFPDYY7M6F3LS/qYTm+gMUKps4KnaePR2bX7V
Gg7n8KfC4DiNgPizvQpAZc/cty9ck9nLEnQyubnHAm4jBrKOpDPztF+SH42S9SnL
3QDE24hKibpftmfOQRTE6sNikci1A131rWss/lUQRPnrOSVzMq0UvnBv85vYjDE7
HQbXclkBL2P3MZzjNQOV1gTn+wyiZKne94XwndDpsl7Vm63GzxLCE4BObMlT/1iC
+dIiHRLz9wZWXFZSgIagHE6Dddcd3CupinnIipJd7GYEK4JhnHKXLsv+m9TIASP2
NhIMKt3hjAGqAA1ZlDR68/ZdD8EqNAdWeB4LIusRfNs5qnsIEI7xheg13Md+wMK4
J1N6MrFqBgy5GV9dUyDZglJkHTdB0YmT6YHqOgcZePQoDH3cIfjBVImZnzJfat9R
gDxvp1+lbjNoXCc4HYgdhvvfhlIU4vbqCh6AxozLZALSlfo4D8reiC5EVPza5SF+
80e0XwpfDjgfQkVks58TW6kSpYKnBp7zRVtDJ6ydYuYtgeAtX2+Sp9aO9fSXKTO9
jhqb8oum7ZN6j3IIRwMFdj38GS1I5MqnhLDaPOK8pzYgarU1Q9oBGnX3WOwsNIvZ
a8Xhr31OdGiGoNt9tV6CCZk234oIsjC+e63E04Ef57WQRiSFQ1mAYROw4YSCxQ3h
YQjBUs0KpSEoJ3IkahrSqeNViSeSFNSdHMg+sCGqWTZX+QTV+1xcGMIdszbReNNE
sSKyWr19aCtOUGlLOVeESuKmczA38Bc9vLmgIcaFev8mZTuyVZy16JeCAoxDY+8b
AHOG46YKy07UGt6lNt4pVsCNMrsQcwG3yTA7lPa+9U9zi1svRXD6N7sL/R+HJ0SZ
7CSH5FNKCQUR/ksTO6US6gKybgS78zxcMTYlvSCI2KcvUeIw8f9tWkX5VLs/Ct5i
iwzIXCoTyZETaWu7xRf8rsQQRhFKT3B6R6sooUm5Cgu9mg3beSinWVu5rsfQsMvg
tjVALMl2wTS4+2gQBdGUXzix6m/MHCxBaJdCUA90xdxL/hvQoyT6LJIEZuq9MsAt
aTqxNJRUjpkqSDtKxf25aHTaBRN0h7B/U2R3RiZLpZZKZOgU4F8rEiOP2fz5ToL5
u2P4MZhwaiCqzFRgJhhyBuP2TSU9MIr8ooZsdnFFdxevKpUxfEIioYXDjN1sUG3d
MGmN6jmTbCbDaebxV5TjL8UtSs2+sJ+arPSUmfSji/k7nE4uPzaDhGW6LvTdcYAm
BKiqGh1BJ4ABn3tCGTDAzSp6L4VcH/7PV/PfKfspgm+aOBQotG17WeCQL9lqiyh/
A0Ewgh0u3lCAGUNW8dMD/4DVKyul5K7N3TrW3Bb3pfz4vIqdnOksLq0hD6QjDMG3
crzVFhsmvgiEhtNAQebpABEgGUSRGArQjSiPqPyGpS0ZA0L0UOH+0CH5XGVuC1wa
rzkDTVcOnpmWBAuiI1XvtLf7FPMxrYRo/Dxa0uh3Pdw2440SFBZFxJsfoE83xio9
hIaKeJmwB38f3myFC0bUuyApijL1+JgFMgZv64yZNpLqDz6nL50CxBSMZQ/buRbG
n3YRqeSMA0WC6Qxp9+CDW2rCT7Zr9UvJ8dBAMVdakHnqSTVh862mhrwheaQUZsHz
zR+ed2MGWF6f8owgRUrp9jWB5rRfqgwQhZZcfzoOlGEJzxq0MxRdO1SR/sZDuAt7
sX0KWhEEfX+tynadmuvZauSd25kvmUJr8mHfd5BulSpAAgVmedVVbnnhwD58aqy5
inyE/yo3CqV04RFiDGHmJjcMkD6NaPy9wB/Y0ohxDK4=
`protect END_PROTECTED
