`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lV8hDb3Qo8b3wC6OHBoI6V9ZYbm7F4ft8qjChLD4EmxM8ZCqvJzaNQPT2gCyxIwb
X9KX1oZNKQfrjNh8k6o+83t31yXvQ1VkmpKj6Ji7uefEQs9F6MgrXMYfTzXUk/9d
xGehMlOWcTG6iqupdRlVZRLMmMB56CtiE7BgmPJWb4vLd7cm4+w0RQPs2G14ObYJ
39gcN9PJvqyo7fvxUKfhvmKqJy4EoaPCNwfLHOVgXH0GKytYd0t/f3erPzqqDWjt
aBcPiVdcpZ71wxO0Ebx9nph6ISaUbEBRWz9i6PQzwos9plM6+5xKPxVOcKLoi8pD
k+9HovQ60dQG5lgXxWkYb7EkIvpio9sc43XpHtBVBrnlBKniH1pcfk/pm3L4jTS8
GjWAABE7R9PhdIt5XdzzZ8qI+BjRvfpsYzKlLB5Vy3uQwQLfNbOEdYheA9ng9aRS
vuZo1Q/E1a9B0IIPAHtvYnnCNN3O6ksenmsCSalICn/4balMDHvpycGUZBpK5OdS
vZqCRGEu7g8EI2FC1zcwHKqPwHsBeRgJ+T5269gh2O27ljxlK3Tgn6UY8aEEKAqv
+y36KZFcDbAgngWOv725l7CbCn7oRmN2W+cW6ABIuxEGujMLqO3vqKExdQThn/CT
URas68DVdEN2cHxv1L4Y4yQUZ0fs0Vv9H62quihVgrFBu2bf55WCHigd+WdQUlvB
XBUL7pcSUxsKZ/v2ph/LL/e1VgsSnSVbsaZ4J6e8pDt890NOeckcxSNqtwjxarhG
CyLEvpbg6mQCYSu7Pw9zT8FvJlrlN1ksmxCSgsp9qSkGCyeAi+makipPOkRAh6AU
kxjMElyrLk1NCMwpeATNCaGhJKNNCH3xYt+ItO4I6ig23RrAG4fzGaIX/6RxmYl3
fa5jJ9AcjX/rO6obFeNuSfxfl+gYnZGseD/fujOgbGLvUgctVDhNEFiuMYpzmYCb
QAt3Vj+QoSqD7xTe0mG2H9f86G4M06yfyReQMlluiOxkdR9OfO35hBRGINZ9x7nj
0eLv77VMhHduKnlrXyNfO56QJO4CEZ9UBVUH+dG43yYmghrxKLNme+CRriwHL9NK
u8ycZSxqR9e0jaVXj3HRVh9d4N+JXGUV340H3ovh/3RlKlKiH9Apg3QRMOiMCIqH
XDg8xKxsxOVc/3Rf1cvyOAaPcII5Y4LOBL9BS1Ltq6IF7eUpSaZ3uEjH2MNCjQZE
ivzMyIdPkKusxQYAZg9+2bfX0796Gl5GfuPDx0ThE5b4shYUIF9ilVIQR3RiF0EE
C4Sg3eJot/iaF6ToyHSyAFjRmRUflLK1pJOAMqimOf6Qt/F74+uL4JiV/e38EuHl
E+LKEwvShcv6O4YoynLMfYh4BXMZeRHH0q+qS9Io3/88+ahdOWrGtRuQcHg21p+W
7yiBaqv2sh8+OlLoL5hWvNhYu5FU3NXC/DYj7QgEBA/HR/Kc91VT13FdhMiR+FGs
/TbMu14zYnx54tjSdFz7ZdX5mQT2p4P8jMRu51zu+WY=
`protect END_PROTECTED
