`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mqkMWqR4tWybMsUfTnN97UqrGM910Kw9ycGU9aNhc9+UJvxa2ch/CJdARrO6C7Ct
DpV3vPCi8NmKj5NzACSqJYkf0zS4AcxxY8dLjUxV2gdKpLuJnbk79YybP/ZTqp7O
IAa2z4rP2ErPaM+NNdydl0JQRFB0dCWj6fBveQcenEe/FnZRoeAWmEYIcwf7kNCL
dNJc/M+Mp8cgR1GPkORsUTYooXZjPzOamgfnZ+KNe/GqA4JVC0ln+8RDHaMsFJlt
4XcFbui2jTupcCa9g+Y1pdLMcEp/7JqWBUoOvCLbc9Oa0mb+wVe7UH2ZyJrKLeNT
fPRY0N5cEYXXEub0vUSLSfSWjPO400YPqQ2bwUKiFqFNZfMxb0IIju/JycMAZkSa
5x0YWWrnf3c/FlHGTML9IvQmP98gYvTw/MsorsyAhrdE+BNaYK4j/o4UE7GslGRE
hZOmOXcES8r7t2tzfTyQamNati/G+l2CEN34H+2YJUc8S3OWjMwOJ1vOmmLDdd7r
iweCtVa6c7nrifBH6F2iZsFXlsWArvcdr9KC3I/U6MaBEkv5242U/6wrvFo4SO0I
/rOtksiPW2sa+q8+qMPWaAWGKP5KvTj0c6eusklzt3oap7g0rSL1OMsmvdSQ1ano
ZNfXs0LxhI6VvTNqsG2f4zKEQkb/hgfOTPUyAeQN/MqCr3r5H5aiOuW+gzRl5rhx
v26O47UzpWoZiagO5UfpNftwDpV2ec1xRMfZ65J7juU7eVUrkgfwVjl7erhBq6fu
bOefJWrznVaqaZ37mV/nXMMJPGfVaUw3Axj/0N8lgu+aYrxpa/BsgTM+R46qp6wx
epK9np1a9pwPi7qLXc8L2LV7ydBBUc9+ugJdmml4lYC5M3BidI8z82VN1BPJ3nyR
kBBUo8hEtE2WMEwpKjFNBkwX0AjJa5pLeM9HQix7tHt+RLHYlpnX/DYHCLjJ9R+o
KwYtl+uAh7g1yO2rwgPpL5hSrLFqfpcH/1wR3PMrtRyO/fpsyzM5rIjQNJH+mAra
ALBLSTXHVAWKKNP5WsFaKp17k9yhTYkTKad0aRL7UoM46Doi8867O97949uOPyUM
JGMjKaG+ZyoAnEkjBTN87uCDsq6/VD73Xkg6Y71mW2efLhx6Nwl5H4HLPDQQstQP
jha2j+2/BUihsD+Zu9fOOaP8few9sEZYK9V98yNqqY2uCuG05Zkhz9i5EHSAF1Gl
zQ2l+nyJzWnhtPnN6SJ9zyVbAwA8YpJvoiX0bO8Ov0crGNbOLXWBA3AQNS7vBbaL
BDBwIQHdWrAjE5pSiaWbUNCaDrPk3JRT3N8gBWIpa7CR8t6mRbtb2EKIRpu9SpZY
`protect END_PROTECTED
