`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGJ8ue+L3lSpJ4Ey75kcAmlp6CjBAkO97gCby+OJ8A1B8RoPq8NRn8XdpjcXbSJG
5C5SXrmaKmTPD/UsPpGVA0YtpN4ea7A9PL9tE223c0h1nvfTxmvG7MSN07PRK73S
wLkNkwaajWi86WpwatoUR7jUT4xCoIRt1xk5tsQyRdmOR15MsOrle9yvkYiWWw1F
CYWuJFTf7Qm3UM/i9ZnpYftXLVzXNLo5gbkj50pzAW8hu7S6t9eFCFm9FqFpgTH8
bwKkBj9L1oBEe6wqdw/BAUYijMzxYnS475sVAN1PNVgbbvQx5aZMO0X0Mtxz+3Yb
zVk43m2P3ddtSBkm8h0hfr1Zf35EnsWVXrQKhNPYw/v/HALvtzpJwlO+CPkXcZCN
2ENXXmZbdhxFi0+MDAPBK0c+XhMIFyRptlIJpNSXE892hVuatOk+8sNGtAou8kTL
zOfNdbpM/kZyyH0spzgrTWYSyinWIFaDxNKN7/f07a74GsBhJ1hG7+ALKzHoQhX0
XCg/HGjlyJFhCu7Bhl215sZWlUAFyvg3w4fKuKDSFG2N0mIm1cbFsRFFAT9Dx93B
UFCbfycjId/15oYCKhChdTx5j/fD2MkLAb9dmtcXohj83Tnthv+18qpjz8THRClf
IxVmNsrMPTL4n+Vfn2KtBqGVZW6+gU2699b3EW8eNbg7aTVmOnbgWlR2mLi0hDV9
I+hZ8/94E3sEq1HgwGXj0GHycuE+LiLmjCmYAOgNnanQhwgsQ6Lj64I1AtY4YVH0
4f8cfofDLHWfmhqhlArhIHipCZ8nUkgsha2uG/HydH4fF1h6EHV8Khw3IqwzJGxD
IYhHpBXxTNIC/XjPwdGGewlXfLqKl7GDDLWLnDSrZCKT7x7xDuRaIDvhV4hUN0GH
u90d5ySiJol3Qvw+/sRA5g==
`protect END_PROTECTED
