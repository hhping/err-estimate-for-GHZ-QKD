`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/m2vWFdfH5u160KLjG8Qp++7ClM/QFhgNjhKhDAKV9tN0IFyyThZyvVgSxnX14J/
U6p/CvksgTcpB0qeg+gvwpYyY+sYJw+iOhArYdMU6WHYbImRbEM2n+cnNLqwU9hM
qoPc0nN0YcCQW5tylnB3XAPfCiCCcmMdpOwJKSMULRKBHTqEGxtqZok5nx28YJVm
q0TcFyQSCms45wU8NKIzq7Zom2y3RTO1Cim2MQE35zrECnCI/iL8s6Ri0wBn6iXI
DGGRw7y7h8L3fX9dFHzstgt/xc2YyjQTXerfjcoEpkShEnJ7fIv6IzpSro1FYdUX
uxGwa3Psga9kfrkBlsQbhicaKunhy1IGs1YKh6C0GMF3YSyb1ecRXTLIia0FN7TU
HsueZDvPjP2R1mM1p7nQ0kK8DlOabe9tkU+UzOV/334CmDQ82mDoJYZk6GaQd4jx
BZwaonKTW2OaSNQZYYCxgWCemy9sj0uQarvm2bg0iL0F0v5nghTLWYW+qb3qOyzc
stjf0je8IJAwkioCOdGjRVi08jbbSnP5lsg47BQXVYD53SI/xe/H3gv1MaB9czVc
doFDSZxaqFce12RDAOuveG8riF20mZlWzTMm2kAqVZKRkm2bjKVkDkcpovBUuBw1
+tZtLctThaBr15nMxDBwtw==
`protect END_PROTECTED
