`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVHQaFUvsRsdbGSfW1JTq4Spuc1n3LPGLFmm3LCV0K1ibD3H2KnUQ4KbmNwO4EID
LrSCew6pQv1qOvIo9UU1PrbpJ/YLkLKStUlqX/4EKoe/ru9Hj1Nhb8dKRuWODw/U
DOmbRLLsOWv5J5uUVRY3XrV6zXkbDgc7cZ6lT95fbBrTQ+s/WjJOoNlzQz47KXqz
K9ztrUxsNmHEFSnfR4SZpO4poJUcF/H4qJtKjLGhfamIaNVb5f3O+pmGqL469C3i
enEkaQGK56f2Epp3bFv/xYjxo48Y8r/sBXa9p0QoPQAqL8eny6XeLZG/KfLFa3nx
dlRdi53U3LZTg8MK3NK9j+3vnOtkI7WjHHrJCSDU19IYEZHVDrG1EisFJAcQ6jaI
6NCGbrZqRJFGHfEsSGcBWwnYcpu3BYC1bl1YBHYsX3YEdJ/HNnn+bGnJsev3v7yU
rguLDyZGueGMlXfDgk/AaQ==
`protect END_PROTECTED
