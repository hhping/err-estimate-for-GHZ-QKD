`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYBKgWxcmt9oe+PysrYryZ31YEv5KA41fVOZuZnp8YIS+YFvbF/GZXjHQc4oqDxR
K6rmhZcykG/XxUiI5hHfRPbqRnPKxNhTc+XhpWh4ZGubWGJzdPS7Aql/td5tvGu9
ejiR78dmRympMlzfx3HnYgEWmNVrYfbT2XKBccSrAfm+178hp2VeXyQBppgmAm2P
BJA9NaYGdEPuSmDOsm3DlMyMhCTgmF5sMV4Q27mIkdxD6aExlmgtpfpGJIIykN7f
q1tDc72rlT4mhbjPD6la1KQUhjd4x9UP5bPiVPYY8W8AUXRlOMOQRQEeUXrzZYY2
bpb7P9aW/5qWHnE1gCVgOafD5om97lZB7+cUYKSGep9hf57a6RxA9c3ZJPy2CzlS
3LVTYa9h0Z/vcMI5HRAh8jkz3N4WAOB6CD8Bww5Z2jaZmm1dsH7c/GSCN+tN4Hzc
N2C9aCnllKnyAkE7yvBhZeZa/x0cAN4JJfZIgPsuzsCLhcS1gVtSv/7nCt2YGX3b
gtarh/5nThbllFG2PfhIvFyxXMY0RETM0lMZE3fl8DSwq+iSVnydYgfyLg3/gPUf
nX90Sz7s0n1luotfnrn9WIpPVWi9mbgmbzVAGcLKVrGHbgwMvJ8ByXVa3Qs50dPv
aSm2oTB0deKqGyb5bLd16yaP5Pa2LNs5WWT4C52k7OoZb7iIW1CcMdcsHt2Q4yxv
urzU0JwS5+UfDRX+9X5WI+dfukf7YdvjjrNt8GHaNPf43AzZiZ0QZWNyJ3v4XU6s
gROsIjI+UYnYPvdZwW2qIeqiXEhEbz+NhuxDyAklALb5io25uoDlYpzXTAXuFyD/
KBUJEXyppBu7/mzHbcpScdwLue4rpNq0EldbjHm87dklH/tmkadrvyB8Mp5EGI5E
i4LsOv5OcKhnqeH40Jid6P2Yy+XgskdwXZYq2kchQeaM3M//dJBgQ3ZBBSk+DdK0
/Z27iJORglYRg+dyE6FxIdfu22/TQYUTMMiuZakhp99/ygfwOBsfkT08vJ+E8W1W
Cs0qRtoyb8cLoAtkPOo1CKRW2uLCONqf2+e8uqDE8/OYiZsdkdMesnmG95vvHpgb
txudy8d2uq+oZgfj5Jd+LMyKRgWHzEyLIomAN9odCFWscrwwaF5eCOge+K6eGpxX
U2hYc/L8X+NVpLWVGfZK+5pSvRIZK2B7DiHpk3X6FfQcw0HVt/rx8WK/N/ErzcB/
i2eAYwZOQ2KVZwkrWCu/O4GHbV3Ux2Vtt2qmOFeGYz+mF53Afn+UJpQvJ1OQJ+BM
A3vcXfo58uv2JOsKGPkzgePTnTdyahKBhBz5ndSMJ4rebHW5OdH7uPk0D5mDSZwH
rMBvA8+ZQhZk46VlgmWw9+GJT3A4JCKI+Tbd9N6NpmpzrzT7LzjW9qC+mG5KGItH
KIKAxAc41FptJKaHMTEXbUnGcI33HkF1keaPJ6uB9MDqIJfDEPKw6TUnt4ds8jFf
iOOciHo6nCStbw4yt+9PW1uMGw9m0i/0TYw41LAe5T2oKHCaFhGvzLeN+vIkE2KJ
hI2gBeI2AR78ItyAOVdCo3nppQiOIEjZz72N3omofJkUlgaNcE9bBifT/sZYCnhJ
Yxrw4i9V71UjMOqB/enzew==
`protect END_PROTECTED
