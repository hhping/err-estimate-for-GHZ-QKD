`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2B1Aqm9IheN3I2Z7qEYbTFKRt75huv0wA+mkaPPE6YcbAUpAJmlB8l7uPqCaS8j
Izs2igX5K3PNO52RSyEKPOQqBNOLQrA2rBNBech5E31MDHnCaIyos68QggjDrElk
iiWsN8iFO0S3h1Q8mKJ3o34poRE+AAqEpsurOP+MqNksFS0Es6L7kNhE1tVt8zfg
jX0E/+gZ4+JvWHJsXcbxykNA/+j+PP/tRA/wx+0mttw1SqgcT44+PHAXgGWE+DyR
YZriPkUAfcLebNxlqnWJctWMc7KqotHDRUvyJnuVCOUx/UE1fQm6DOOMFLPuZ4K+
3/zvpTzmzLWiMQ266x6wGDG/row00Bkg2Y7FGu5/WEbCo9lV2MqseZi4HPVtMFbb
pyDaGwkkgEScc3ww65VBeF8Nk2B9/H3R/8AYO5ki7qM+gbfTw/Lo4XKs0DT6rFEu
6V6AxOgRPGAwgVgZL7vuwh1vHVpt3wWd7vKeEnUCYY5TANJzoz3W1b94YjZ6DzKx
vPbD6vjfMN2aRVelMBQ6PYbCykgInVYEwQwqaVx9P3SoqQRJWuppNuPuTA9Xuzzj
FkfOGtPFzl6MsLaUCA6jdUjh+o6RLK6c8idL5H8foBtURTjlnjmxyhLH3M8sCJAP
zF8R7NeXeJxY3xbe4M6+JXFEFbibvsfXuTdnsbB0396SXIzFZXY+LyCEOLUfRtVn
zek1tWlvuBkneXNKypDkAwQ+8t8I3xZt06O/m7iikqCJKYU8rBeIWgvQR8tYlXsI
5YkWyCHMbCz08HTcVhY4Dpc/7e5xdcFNk/dETYWfAYYJZyHxTqwzb4tPblwPo394
VIQ1j5G/Y2P29+yECIAwlzJgqsTkTZsM4RWNMBnmqJIJo2xpd/gEZYMAxZpNkDXF
N7BL6RpuypKuE+31mRt9oMSH0y6/iqwO44nIHmLmX2eRHdEAoYxSy76IlXDd9i7E
B79gVF9ag6uv3qL40JBKLE84pQrgqj9iWZ25W06OR1N7P+7tp1rUzz69RgQ3fkOS
Be2G2pwXE7WWGCRaObDw+8PNaKcKwGB2VdLPTUptE/CvQYSOFeHf47xLv8sbnQOt
bXjArsXF8vhyNstpZ4lGfUAO2hDX0lzy+f7l2eaT+mboAifvj+ox9N9bzaI33HXs
ODQ2WxWt/krPt2a8trC/Pr0ISjRN+AKpFlwsL5EBqAksMDfla6golXd5YLJDEvvS
DOa+mF76zHI3K1owXlpzulG8q/WA+y8RVy9rUkngoGGbwbU511TrcZBVx3wREm7E
i2cf/e5UwEJSNJwcpB0NELFBqBfUtM+PkOLFxU6TDSqdz7l+/2xpGH6R2xZ1mVVz
cOT9cXdzL0tIInqzmfSOAzIrwOfqvAV17yTi4Ue/VUQaIEPnBe8s4jquudVKJN2V
XTFcMPgpEzXrU/oKBPivScdS/bbps1LwYbRE7SrC/ql1dvrGvmHZSQNMYcbxE9Kj
/9J8jZWHFAh2HvNZ/g8A4KQAND2VFkuA+UXsK8ef0r+NtBQA3KjB+43ANWGvsqfd
QBhIASb1Ahc89/2NLtEF4RyjAn3NoXZgzy8udpRXpbuXhlhC43jTFpMcyT0uhNdz
8d+0NZMuRJvoo3oxPv7rFHKDSQG9lMCvSEFBxALEcUrWFR6P6v3lY4ENTPA6GfiG
6D2TLuLMx0PyIPuEuN36dDphkjBx0w9xDlQcXyV/7oC5ou5tMWV8LyGwNP/vXe8K
SsEs3HR1jiDSQLQB01bOMImdRbMHfE+f/rBYc4g+LYhTFbtzfRhfeY7a1jooES5/
EPMDClHIn+VgAm4n8k23fzScBTrvMdDqklSiu6fL4ekvqV/jjYopLocISyLAmLaL
Um1IXSwbEVPoHHzRfJ48ir7G7RwpEyg4bKZgNb1NafxQndZrGdHfk6fLcijl+7iv
67nCJPkxISlEyE4fGrY0YjZfjmw0oATzTkg8Hp8csdW+xJowyEexgmwYvo5XyoQo
e2dqYTkQuoLDOuR8Dhqh5Z/zpBN1RyTDVBhkh7zolvi1Rg1n4jLh5nYIFJFtPtuw
aJqdUcHAlJ3QlTxH6nqI1smcN21tmiEd5+hpE0L3z3X4SG8huFfkgXc3mnRuVbnw
d9NFZWbR4GaV4XtdxocAl8455Gntdi4bEmoaodosGB96e7nGOUZpICVPQkxisHWQ
TDqUZ2VPEynUgU+7MaItIQRrvLTyGmdcJHRmFDevll9LgileN8cYVk2WjOKmTStT
pW/4NOZK7gY94BuYyRBBMSqAz5GdMGgbdwhdapfaGeVyEEQNlBT/oq+HkTylQKjn
t0flV6v5eBrTIADYQAkh6vwwtx1169ozOliYbqpIMcx1ii9AWI/H3nM8En8DkhpF
9MHu7Bw79r5dSpjzBB/kFeQhk+N4PPjrRwe84sd9sp7M/GsoUZcWqAGGfo4e7TA/
56vfW2nOmLfEszmLwQ+YiLYbLe9F80innNjivbqNjVSP/ixHgkcUsZmnjOuNvwpL
EO3kqebqzwOIzevRta0AFEqbsdyxxPPwwaBemAOARayoRFSCo8cbvdB064XBGZi7
Vc5HPIviY+UbhIqTSw44juoErLMJFijrPVXZ717e5fr9XAbJeEtnU+Yb3khUhR9X
+q1YG7o+fk5fE7t02t1awcLBXGNVEf33vwRz7cIRvCPKQ741rL4VYIj2NHuraoK1
naaAsGYSIpkZE3raTeLY97q4Mjp7Mguk3ZopTyTtkrxr+rXqz8cgC0uCp70OZvJp
ww8Ni5OZzkn/0Z0OHQ5gdF/vivPWFp7EnWJj9205aFD9ksBCLRYkS8aoi5lwNkWo
7HYkgYDSvmjaymrHVl7dLcjyDpzYoI9jmpkSNW35xxjG+/+z3TsFEzvMUVL0S15Z
4HnvrSIMYB0IXPBCxP3IzCPw9QUofwsmeSdmFKsR6o3dQo72ZItgox9FDKdH7ZeS
aKHvHyL+58GOzsbZe6OK7cnT4h+GxY3W9CuaByxIGNOo3+0FQ9tPdUcehL034Udb
D1dNOkROFiFIREgLVCvHyVXtJybPFOCwhnbJcGN8aydleG7u/UmZ88l8ZaF4MmVp
QVnQPi9f0V3xK/Lcw9moxXVTBQ9EHTSBkIlV80Qg0Vwnut5PaCq8mf/MH80eF1ed
fAUpYPauCDwNrYrqw3/grxY+EHZ2HJpslk/THPbkORBsKhiq5vhJVDMqSX0riMpK
P2IVq5bA1imoESjH481GzOvZQHbb4rGY2SD6uNjch+lUXEPLZNtQyBnIDICCXB7G
xBumlJgBGNngbYZ+ikGr16ORoUhODbufGpI61BJ21dtArT9Dbtw6+gz5VEIKNDXs
Lqd2tudaWBZteQuepRI3h67WkoYxmhb9o45WKhNpVXTMeF7kwheVR8QKjOtoOJjn
unAbRCfjJykDZ8TRrXQASb8TtK5uGoxB7dgUovurUfEeem5kqZGlTd7cqyM8dTt/
ejj/Rn2dWkNm1lht63DXEa5ZHlxKeNyeaNmbKjPL+N5LKLvlVrIT16rZ6cLcfcLk
+fH8BXQPWe5FhwwKOf05fqgftLs0f9Vw+p+TofB5+WmXicrBhAI5kSIpyO61yqry
YKXcc6lbN/81mOY5X+FfIzJa8Bd5MBbogvT12C0BHgi7eOHBnAZxYw4ye8LkWgop
WvrP4ldBYeo5Hlw9HOFkm6zo6Yma7H/IYTY8gujcmlwpr5MmEyXhqa/Wsw2PPNxG
l52gXUPHNjcjMVGkhcG+locm/vMlCQQQvCPg8yzpxCkf9Om5i0rR/faWuSSthhsO
tAke7G2eGvpreZBlMFF/kwpkGzECWOhlF7dBKDbhPdA5jff5t/TzHDrJys423LbF
fJ18vkwseWTepUPD5T8iW+Ouh0FuoX0g1+tY/tP3kgPtVaMIPeo8rvqtX4z+mi3u
3TGhgcrOr66jR55pGpuR1Mfjmk/Ap4k9M5UbP+3zEMQUML7TXSd5HxOpESg8zkwx
NlFPJ1+lW8wT5pGsWUu5Mcl5y5jsNU5NKxAelpJ/rniSOFHDvUgPacv64GvbBoIN
1KGVw3FPyaXern/9H0KrgBePOTMSjN5s99Gr9Em50/0Rrk51W/FfcjHgSp9nz0p3
gnLrEr4QoUFyJt2d5OTMZq13zZgLVNxna5WSXZE9Ggyqc2dUz7UXJvrV9W7RrW2N
TS+piRYNPkUUFZKdceVojMo4VvdQehRKmv1K/sGQ+CAIxXLYcN4j8EV+3j1VOF/Q
2vfznWgp6mXLjBb0PGd5tnm+DTwlOfQYsq+ROO2juaaQEYW3uTFYin0sSz6ip1j2
3KVEvnJ+jGxFkGXpi0nmMJE69dJsthLzyNvpPG2bDQg1GS9z2V1EOkC75kwsLZiT
T77krAFchHAU6lVLDHOOLZGHBlntisMk0II9Oazaw0tX9/ObQBVElfkh3dr79F2O
Ig+MBjk6w0nXNxL2ivBvppB1a5PHelmM/cT+PAaTKrsxsK7cZ3qkrhv7XbaNq3hE
uFNBW+ucUoBSaqypnfxCE43d2msMhxW462LCL80usgpWACFSdiloS4eeDICSNcMq
Tt0m+PcmclplAvohe/kBQDAdHrhIzchLGflqUqDC7j1QiaMnfqPYZFb6skZIE5xI
0akfJH1qKE6Ucs2VIn16sRSQMDbYrDU5q+2DlVG+y7Y2bV73CYh+EuXj6BkofqDE
7qxdXRhejN4qyiZlDlLnXZwQvkTvQFrEpbZdKWRMCFSpaTNBTttYtXfb/FsIK6eJ
+HHxGOe5dHt2YoK51znCFY/ANBCo03ndO7hU0Ob0IDHuefY6e0M0IbMlLYfv5haQ
1dD/az8kvfzJpowF49HxLNHmUBnvg4AQnR6c57CR8CdiHyryo9ATotJd6mRr90zt
fCrclYWM+8dPBX1uVAfMhq4KsBcX0gJjXkDLl7XzX8dZw5FVaRoNB2jOxlfh/A2m
cu9fHvDuc2LH51WeywbYJWKciDld8YvyiTBAyEwx36gI3YbEb1Iif5IrHPzTrVCd
0I4cYWBORY6fyj4E0GE7I9UTP+XTO5hxsZoBZpIqiUPM4jOsRNOeEFf9ZN6uESOy
RftPq1TwsJnZHOxCkMc+BL53cRW969HCMlMvEAtkFCSzM9ATHQWwH33EkMbtJmq9
990qrgJ8olDmPNznbKOIC+zKRw4U+he5Y59cV9FTcjMPetYimHZj4Fx+hngBPYJF
r/YZ06A4diB2QXmmFd0x4f9VwAQXa6ksE2Ij7mx5VzQsyz9RWsDjnODtl7sDQNQW
tLlubYucTIuK3W03MpLauXqRgw57TZyJsNmKpSEL+nZbmnMTezebfl0Fp6P1FeGy
PUdiVhBCSefoyflc8sjGKrrtiIPoTBe0U9MqJfWO4NloDnl5N6W4ZMEFc7pAubF5
JhQ2PNXvyoA1pJWpUtq2FiNk9tChaYvI1DO0ScvOX1QRryaNGNTl1TsqVA343HyF
Eh2bHXyY51EXs2L5mJ9hRG7PlOVyN9tnlYvKKBp1EBSSujIRNq3wmi1CGcEQXKlF
6V3TPSam+J+3aLdVGBplTrTV7+L3JEtZVpre0sCUWT9g2GuDrVwBluz8i05FIXMl
oaNkEKLlVApygq1Al0hFpELVo7P3VJ9/omwltS9z2+QMaVksDTWmQ9ByVKZZs9k0
jnjcltFRLtlnNucKjjBpteV/LmnbjSqY8nSAC8Mv2dNOnvKGBtPxWFbLHuyG62/y
DqYKS5rtNp7qVfhIzUyaXYF4qkCTqpKo8rN8RjsUfYZkdKqqQ7ju8aJDcSGf2VZz
oGgDpCISvgMw/eXvkuobIk8wP0SMeiuUUyq0pmwfeLlMieo8VrIgxmhlfyh5qW9g
zuwhQk2PlUJ5Cw22hpUohgi3Bs1cdgupNLVkd0qLnyeqVpwo9Bry86gyf1pQeOWh
HMBy8pV7kpLpSI7duof3qamVm3Hf22QNM5wqq31+MIihZHG5CoNKE9pPF79raObr
5e0FEg2jR/hDYdQ9Ao4Aekzpx8/v911/UWe8vCTO6MDTHu2tle2hXAMZA+F0ip6w
Qf0dv7vCnQK0UA0Ww0a5jgHvtxI7syFejqfpWYV84b2yqGvhEf73KybuT89yMHQQ
QINxIpN8WRd8HZFYeTDG6Z729WCFIju/ep8vOxUxCDYwzM2tL/3dzUz1AU9bD6rZ
smlWsMRY0KfoM8ptadeyyhEQ0KVHrPMd23NLSnlD8GfqBMhIZqvI8RFQFVqUVJnH
xn+VzV3Ov5ZzUotxwqMi1X6rN5gYwk7nC13VZPA4oKeSQvoMmhcgnDpEyRNMg9Wk
AwAOXAiOf0X7XMr7hFF0cx2HhcloFA73v05tFiE58uqUXRfGv3UsYN04lhJ0Jour
8N63uR5F5+CXzQ2aHfR6xNKvHusFHstN5j6gWQTY6utq+/2E3v8l9c0kTiFAnjQI
BJ1U++vEVvMCRVqo57F3f3pAZofG38xQE6gv5xxQ9znJjHGKqdQ9GwL9nhSwseMd
G6j4bLg4DHEJWd7d5YRTVnaa9uaPmS6zr9znpdMOqjJw/flAY3Swk0dwbrvR7u04
DQmBCxxenejB8pALnz8hclqLrHoX/9D3qv2pX3oBo3xkPi1eLU/9yFEDbBy97FD7
Dj7gntvo4L+OEjenYMlrciKiAROUlIdOmY9smBP6NP1DWtmI4+gso7rTAWhET6wS
jgx2u7UjAv+XXJJ3KIiezUCtnACHtNBEx4AqM73EBjTNqNATICU7xsnA4hG2M4Q0
Set42PFFpbGNHiHRDJvtaQ==
`protect END_PROTECTED
