`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRIFCBCsFaLe2jLSg+RYOrNC+T1XfyeJT5ElkY4/eV6uWH8M1sMHa1SDt2aKoXKV
N/uywwqGmLaRn9ZCNBL7LUu5OkjbO1Cycdpr2NuJu1tOXeqjKwDW2/rNScJiOzdB
ynnx+CeWEKofshLpEAuiqjmOwrqHXraRpskUgzbtehKt51UK+58zOFBWqK2MKjCy
x84+0I7iJrQNlb+UNEJMtPec+jRvR+DsnqJcgxkiLuWdxBJojf+OLvkOp6NJkjvm
qOSuao3Z5nPTNMEDM/X5ZmKOoWE43LGsfd5cJf+yRa1T55hAsK30gVESMGEUq/fe
7a3GfJ2w3FqUBZzqesbo4Z5Hu0lpJdORRTG5A4TsG0a8UikiBEagwW8zH2sxXJAo
J7AJhkGvyI3MsRBnQe5rDJoQKaGSsVF6oL9Q5R8+rjoj9dj2NfQYNUAsAvtymMU1
uBF/iIyO8V/n9SqeWmfS0+QL+nYGhk7KbDKnPSMZ6sjsXvRTJnScMMoJXqJhWwy1
9dyZseEOc6G36iY67qFdSr/PFeIdsbd834akGBuD/o1nI7oAkq+GlsAy7WdDgfcQ
edZo43NSg3bFMC41ZE0YYnR5k3rbGIOngavyhVC3PVjrhwUTn/SSkecrFMR2ZUXU
nzEygLPrlscB4PTi7RpySMiprA4WnZDSrHowtc9Nk8VF0NvviEwDkX1wkkaqVu86
RODfeSvatWuIw7wBPCzWByjW4KfyaBTQ4mPmw9ACOdJOvP25O6MXg41WdzB4zDSs
a4F99odikkj6jBOQV7vocxjFqGN1QYs7or2kIvBszJAoidCREsTAQ3IZpNBn6bpP
iKEY3Moqf3kXRIXZc4R8nxyfJrvMklJT4ZAwuWsVNZ/x8VSFMMWVew+/4q2gsMfn
i2Pv0HKTu39+7v+qwZfNHRs8ZEPYEoGyWgwi1OkC4yCsLRhOG1zl7M1g7gkmsPuj
TURjNMGy59u9W8a9mqu3X6S7nBtl7NO63diV6104VHap0vXlmd6XbT+fB/E53xSY
g8CApWS5ZCnAx/gC06MCc+u+alM1Q1ebDa9KsBYd96NunJvXvLWdqcg+Z/9JnI0r
+GIXBQLdERzXpChm9zRoprh07NCagA3A6fE5RazR+vhmZgYuPfllccPKGf9J7coe
++lnOx8OukdZw1JmhPEZG08HCgmwleZZp0Y0P/VlGuU+OyjDj9jIOXGh47nhqbqx
YbRmA6WqaHXTLm9hUHdEjc5WcOJH6v6gYj3M7WzE34DCc8l1oIKVNeBMnl9gMUWu
N8Tbl08Dri0dWZ5jLCuZ+zRSZuduyImAolSMKOXfEJySaoeyOoC8jp3BVcZ4/fbP
bm0Q1nSQqiKMI9lBrI0NWeFG245tHpurG7Z0ua/s41VWYQxGOe2a9couy5MHm0Gq
GX7C/KO3JlALZw17KqZowei8o5mVULDvNx+pKWQx61+acwA8zA/lJjbV/TQykv8i
YXimOg8V2YuRXY7L+Sdljl8+uOrk/rRJA5tgV9IazEb7upF0ZTbWST2Rcfqs7Yz3
HwmFGLO72/lnzhDYVpp/d8e18MEVk9n+t3z8FR2rmqdB7HnD3lM3XvPnnCuNSlhw
aAORDLQxd2XJWIsfHtx8FP/TC0U1Gkv8RhfVGB7jMuWEUdcEqPdLmADm/0wI5ySF
2UkCS6RZCeiHlE6WEjxhPAg9VhnZlsodsLC2yFqYMFz46HusPcIMGN7Bfj37XyYq
Xnt3Y1/y1g5kR5PiNVE9VhMnBvLWBQ6cdshUZLs4EQumFuKTFsqtukOqbJ+mzlUN
4UfZhtDbi4N6LLpcfHTUgsT3tY7lnEz6PQa70XcD8Xf24nf012BgT2Pm6wmwEVCk
rusyeFk+gQmVXZI9NRx2c9ZKC+oJavw48P556dIa+0lmps8R+EIFCV8ubGg+GdsY
R/BdAl7PtUdwt1Cr+xd5+6J9Tw3VbfdtVsgmigmEuvFqXGXcauwPY7+4Qk9ALY3T
yubshOM/pTSplAnIbE+dpdfJVLkr/9d4FuQC5U81r6HV15GBatvHd9wSwQ8LVdrx
fNd9u0eu3Uy7yGJYagQCxyZd+XV41pa5PMgLbUfl4NvKxAKJYAbkOSMICZsBgkye
CZnZucy9zKf9bWv8TxnosnFkzfGSgs0GMpIwkfjKEpmf5fvScE3unQM90tbUw9cv
9IyPJP3HV2ZFf2jSktEfBnfvVXCvIO58+bsjyYtYIKm7yUSQ14Wjd1+tyH780czy
nZP1MKrhXZRpX6NJ2rfhZ8MKh5wKq4WzrCIaHm9pNzNcPT8woQWA7qjTeeJ6YyX6
Ep2kMj7QTgCj8PJlhckbjt+3xe69B6PEJiuhLVsZjVyb8xE0IxOwQBfG2JeqsA7T
qIXcbXKS6vtpM0bzifcEssFLFmtJlwyS8QrCuQ+Ofxv+BYVulRu6izdadSiwyLFl
O+2ruqBvkoHUHAWQJle2cuMZaUQcFYSM+dakUARLVUbFxY+R3Rfn4CwJedmdX/Yy
d/LQTdbh1GRZMNBIQBYwmPAFJURpEiTXnUhuMKunv5u+/NwbEkbz1oV3EtQCNf5c
cdZBrWKLCC20MX3qLIG2CeBFNeDYGPP7PC9g0ilz9jXUZLEpDmVC7q3vS5h6UywO
bMoazClYR1Nql+hwFOPuEeELrOgjge7Ihh0QERgvjJVbxLEpXwfFg6lyxZJPGE0R
Rc9kaGhmOT3zLFR1jhgDhwI1/dL1Cm34/XqbsirKuNOMyxDA4gH5fOfsmD56Suji
LftLxGIpdmBv5LmM+hIxjM94Job5R7uU/OEGezSK5D+i1qP0RsSTf0VBbeZOeZ2d
W9HmFYVNEkdnmIU/S3wb+EmSI8y5RueBfU/6yTqKhUHCIHuS1nRF6eTCz4FvyXS0
6xrxg8Rrs9VFwl0iUVeyFkcskUQwAGad1zhff2qzIBQWa2aqQWUvgd96Y40n6C8+
1ODICfI0oiWUpegx1a9oMH+kLIb0QLZdezyDgMxA4JpfHWxZtzx4/v+aLoT46Sjc
Kkf0ihbO7ZmlIMqIZSSP0/0DbiQFdAOB6FCwW+UbnirIbCa3rYdsBv4nboXFdMBu
oAS1yvTk3k/ig8k1utdxyXE25aWNlfGB+tiVM6FxJE6Fa+mjSKuXTv9ZLTC9+CcS
f514JAHBs0xvcjtNKa2TdioXZTSpCU4ZNNiRlR21xMKSr7CdrRYaVSR+bmM4+0jU
ksu4cm1RPWcutOHQYsmIY9cePJd9WcLlJzGn9Lkzru4DHcQbcgIPfk1og9GhBY28
8RO6Gox0SjO8ANUvGZ+MeHLj3M2Y709EcPQSfeAK1XJCFDD+0lZxXeBznHiyT8/i
9VPxOZkpZ1uMdDLp402ZslRXhRMN1mGvt+8RaARRtW6kJirPjIBsxj818DejNPRS
Up91U28Tnf2i7SCAYja7qtb9HixexPIet4t7bgttpmRX72hNY9g1xR1DSaxUo5CH
Di5LVr3tdcnpQ5+I5dncDkEU/NeMvEWJvVXBBNc5NjOcE9G4nK2n5oyJrU7SvAjm
MPrSm4MKuT4UrWmkVq+WTsTCSyf2yGkaCWqqjDFqxlTBBeSVjlNt33qMBywEN/bc
B47CVjQL3B5KuFRCpAK0QzNJm/vrsj6SDlfAXFsKpQ0T6fFEpJG2AmnrUG0YaKdR
F6/dPVobv2FSoRoB/g5YDU+P4g9eEFlMlATJHac7HcHF64HxXNUEHsTKEweQPOGd
hBgxU+qSUrPLTOCSN507uO9+OYhZTjptc0EvZWKKKfbwBE/inKr3uD6ZL2thOFfo
HI6kgUginA8dUcyO/kFWa+ifK9RgTdnEzIsOOmJtkk/1JEO7GOcMKyURM9X2oGnF
XFOpOR7kecQ0DBNJ+kLXe619l4leQVVxOFFl1mHgonYAXCksw4ZL/uJXSBOF89e3
tejEQStHyW8Rrkz92osazjDTaSCsjEQyvi50M8jBHQtE1XF5+rSWpKrLOM0Bsd66
WXyrkzrqiJQgM5tytY7/R2csa4qQzZ8/AWTm+1/Ld/F2TzgBFbwft7uFoRrNLEoS
gNGadaGuBsHPkHoiwwFNH6hsC9fayR0UnYjV+ZOsWx8wLPeryC2TrQI7wgeMq42k
ks6duswIqSAe0CJm1Ys5dczRQH/mtejlB56rk78OJ6ysQrYzChS8nZIZpLxMmqcw
a142/jU4f5bLv4mXTB5A2KiTnbKy0FXqJUqvZtSBuePs0zFPSpiamawTgqxYzcO1
Y1H7Yai9pByq7XaH93Y3iJQxDXTkDHv3H5GQbL1MDjWER2QWHXoAwDW30LpEnnso
fSwHbza0RnbJvsQnHBhra3ERNEtGEE1+I3vLREBtkahM9y6+awBrqRcG/8/3Z4XT
hXavMKQ050+Ygl58cB2JV27sQG/jDscSySO11fybXFoy9a8lWBRCMNxgx8/7gIf8
k8u+ejEnY+WLuaMw6X0zvA2Ro/Xslleyo8Thl83YACabrn4JucIdcUVesdBW5iaA
KYEsrlm4J4CXA11u9M4IQXyAOv1b+onf+FZVWEXf4EJjMfbuk8qzhmcmHcTjIR7S
9iWbcUbMX9EROW4ped1NEmkqeITyGYBtgeM29Sg1ZkKyHi4KTRlEMjphIT83KzWq
ASqRz7kDnzvYjoL3dgCXhdrAAHMBKf7VvXo1nMvOn61LN9pES0ysC5tlW9SQv1Nv
NApvhF0KAGLK7hGGsgnhdDfkpyJlSAVWu/mO93sN7oyrypQulcS6WgLnidKimyVd
7VbXMnHmWhfftRCIR+80BmWV/oyrJCf3ZtSIS02gpHfLv65Q8mg/969KXZ6+gOHm
zvUT0ByNmuGMUvT/y5mwSn5h5uDzAMjKcPw/jV+lpn6NB1JuhG0iwiHKjRmBytPH
5PpOkQM8l5inQG1xNbYSnT5HggFv3qNeKYDRK6bYm31CGL7ywrngvP3aBbX6XOPI
+vCl0ZLLkNAbcAARhSa1pg/33EpRkY56dZgx30X6fv68tSBfBEX2G74vAxX9ag9z
Yo/TamwuOsdwn2WfGVvDiJxBd9+pUlhLLbRL+T98n9oddeT51TV9C0e4YwixsLA5
WP71maJttfKwdWPO7OiifKmL1I4sCf+u95HSB6JBGFcdN8/kVMOuTtp7DBN94vJN
P8K8pzWPYbFzvrJUw9DawRHlxj4NiifmhGDIj79uyyl3DH4Ivf153swT2SXzcE8h
kWnltcyF/0V76IsmIgrHjRlJG2ZkUkYLa0tcPs27lOs=
`protect END_PROTECTED
