`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
keEgkR5M44E8mZ8H0mHQJTNmwnjdyBavW9Kw7KSpiT1+35SmeOMgbcXAWTmunw0q
n1fCBZj1k04KO2/qI5q4Qe/p+DzguOa2gQL+842D0y/F5f3PPII9NeC1a/lNgu5v
z9IzrZxWTElsHAV3+hBqidFQ4zKFdv//YyserhpXZVN4PLV2FwzGRH2ICgHDoS+c
O2wiEjmqo++2650gc05jRSb0npPupdHF0/RbgL9PTgnZr0mHlZHkiM044POZ/6WR
tJ4PR7LpbDblje3jbisCyAYu/FT6i6ixUUNzg3smSGBQswl3KQG9erfc7d5Y98AL
mnrGD4tNvLkK3AOeJHg7AeqYjgTHLf7fXTuApwVKPrIxke6VZJd1xD7I5I+49bGo
FbThdaOud5CYR/hNKiptZXOQuSQbbwDkNAT1ggxSt2IEqMEfosGCSfkciJgcZHLA
ajVk/UrX5V/oAI7xICQ/bG42itIW/quqeSk0bI3q4F9CIAwgJ6NOUypnPJWwZr61
QlsB1kR5ZMu2rFSuhrZVpiHPtC0Zn8FNC/cHiwTF+RPNzrWUzjNErf/Dt6pRg2cg
gbGGtZfd/HQYYaAPJHZlCqrj8+Lgu34VGXsL7GjAqib8e24+WP2nPgrXRhtusx89
LPKbKL4+1Zn3EYtQuf9Ml5HjHhAqyIgnUM4IKRGDmbs=
`protect END_PROTECTED
