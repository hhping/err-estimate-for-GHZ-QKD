`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f7a+6wSh7JgjnTl7qD1bM+LxuTZTAG7SQnzbE66cnExkDF1b0ZKTzLWiE32gLXQQ
d9dV5IeT3kVwUVV/EXGgP+JxMbxysytqk1k3D2aAp60ftm1Lh51xRX7evJ2gdxOs
mXyfCNgrSvpWJJQuoi0aZ6FYV6YhVPoZuzUjrGz+lXGTu1AzOkfCQrm+zaZt+AU9
3aPG+7P9bTwm7bcEwEiPBZzEHyWFMcmNW7HAPuqScRVgsA/KhGEi070RfzlbMM2M
0Ld0XbFfJ2+E0UxM+0oBpQHm9rsJjnpFPWNw4ktpUfr9sDRHy40d2tEE7MFF/hSJ
Zq1bpxCpBS6BfYjoZFlwjhkixpgkG0b2LbHPz9d71jnJhbkcG9J0a0bo/HN9v8sN
9JK+ArrWhM97Q/NqXtBDVPVCoNCjBZ8Vl1++POCz41Iz+bDthLT3MpYrNhWD6wcX
aitYUWM8lNfXpd8nS7xWYiYLfqI+YFCm1WxtDDJe6oF0iGUwhfs8ZmNsVT4LQzRo
+Kmet/lV8v6cI0oZ/QiDHjm8++qBV/c+GrY/VLTHi9cNMnw0PSpZoiODBTRmrDdJ
SoqUhfNohSaDVY3GhXf6WXAI3trqqQ0sGBWqJ0wx2U4cdjI6cYfhxk+YhKKxic8N
qLD6ry9eMZz/S5Tj49jPGT/8AZv9U6wUm5Tt95F9WpNMpO9IDHEerJTjEWnm0uLh
hT30YJv+5VmktdhIOeVHSIqlIxmXvSpi08WqfTUqz2beKwrE2OSyQx6kmUGv2utZ
oZe5ZXJWRBD07IrLf9titG375nmz9lCzjBLcEl+PmOR+/L502cpg6vnk4bw6uhbk
grPPGLkKFJ9XEDfb3tvzwhTL9otlnwFo4yWJP+lKxDNahTf8Fdd8mnbfHO0UohYC
hpgxJTZLkxzzYIhu8YLFUHgHITNH0C2AoMZhn8lOLFzyvpkY2MZm3TNEnxcoxhMP
X4mXVRNaNuAy50SF9+daPiG1jMdUZLuup+kUYcO6pcKPo3YpHXHVpfdfHQVXzxTT
abq1uUC2wStb8QDwCg3BRC0L/Hj2Gj1Lo0+e9LVXBfD/5XryRKOjE1BmYiotH8eQ
4M6jwSqoXfRtK2MtNosjsBoFREevrqRgGqEj0ONEsx2eluBwbBmrkCGq23ObCyzI
4sAGaysqCJpTiKTrJICkwRCepGQ2CK3GgTHImNmk0fRSYi20PpUEJ8W3C1egPg0N
my+b/lJtccrnwzxyrHm2SGAm2nc+LnSbGPyUF6lnWrXZ3jruUhxXQhgGL1jiLpFE
Rwd2nxqYGAbWTYfSZidFX+XJ2HQW31VLzAtfBRUe5GrCZD8g7ZcGixieVnx6AQuU
k46qFAJ7Pl4c5lEdMHdcArOjiucEXPr0LB/4xZhscnRHmIbNB0sCMeoB+EfzKfve
+LsOUguwKPBxr/eaUvVWmK1JI2+TGixgg9hr7bwQt5kEX7Mhw/oamEKNqCBHKSp7
Tcx7ljYIjERpnlKJY++/agET1ccE2I8WNASF2DqkWfwiBGqjwzmAqREasXji2ang
8aSPpB2Wi10K4zxEq+uFGEeS82De5vKOoIiYu7y8x+tZrEWzG86ykrpElUYH5hjV
r8ffh5oD9XjBzr0BTlFewUe4CiXWXxXznkFJXTTGHjkuJT/EgmX4PQmeuINpPgwJ
c6zTsemN9gHpEMrpeSOk/CqjXyQqB5FoeNhC7PLuEv33iHgIXNfzMo2EL9NTjv+L
RJujMSMEkvwdxeB16hRNSfS3JGUR5pJx1RJtiY4eP1+TsYeUzSiGc8EbCID2JBkS
SCEFfv6mEeY/fpR+bxttZRAfVjpXT93boWge6G5RMvMGK6JqLvLlLZCtttRaJkhm
Bt87Bmgy3HRkrSSkFnHJWzDYYWOVoTS96LvJJvdC/ALn3F0pmrSALdB6agsEFe/v
ADZMNNDtcGZgf/AAsOHKuJ5x8ZHfG45d+Jgiz4GpNWVIV3hhW5rdSkpwiEFJtnrb
fJTyVbo/vgZyLUpkUmF3BCNgNG698bux/o9tdDT1cE0wVauy6SgB3AoaoiZyp0SJ
8pFzY/6x+w1Aa7/lyA9teZuXFs45ULm3IQx9Pej0UIQ10Pk1ezVuekfEIPvLWCqo
nelGFooL4pSlsX+go1YTBfQfTyXkGfZUbdQqwkc0VS6fez45hDSGCmwTKxi5AH6Q
O1tXpTy0f+R8cZfBsRP5JYJqk5MnQIPky/RhX4kvb714hG4N114mWGu5mxijnrqE
`protect END_PROTECTED
