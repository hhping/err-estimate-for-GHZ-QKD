`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+TxYRwFQWhZ40C+91VPqZeHLINarHXuLEizoKaNIdLNsb6rIx+STOfwujtYUNnb
SvtbGBd8a0HzJlKcZZY+5ZDAvEanqDFKjaI+Sa3O0G/ra28KP20qHDjCQ/gMwrKm
HpsgGJVl/0eTEelNIq5eMtvaE0dEg3su1X9MyjRgKCLSDJIkdKAJxlAUOzcSR7JZ
0EYWzg4OLT2tBzHPwzEsFI+X8EX2HuiP8WA+fr/eH5zYf/teYMma2jKRMTUb6qG4
V4veGrMEFjAAzwn1q86lNYodnKA3dxSFAgeSmurKuvTy7GwwLkNOenGPYauFxmsc
UWmwGi5gfoLJvdVz4Yl8N6m16aIUCqzZm5EXTEWhoHSE5xEsd9F7V4etnu+GUFot
1myvdXOvY0Qeeu9CspencMj78n8Nli8eEUrdPEwLlfKGaghkdMigv651PNpbLP/F
v206ReyvNDaCSBoGADhZ6OXsEE0kJPXiQlDph/8XnEnVzv6mEKqBMt8liRwpaNJR
AKJmKQ0KrYW0pasVJ3VdWIRAKmOZayTQ8x41kLWC23jwm0zCCC/Rshe8Pfao3rK7
TZwD4jtfQN+/OWBNqazT6I0jJFc/lbHZontZTDdKFde7GcZW9z/VjGzHJ0VxS6Un
e2UntXqlwUBGMC7XwVTTW50Lxha3QLqTFIL2VpmYzmxdzsYowfHxfLW5yAUBWbeC
jP8bFp629aR+0VhD8mWMCTdFnC6/bqB7ef04Fm4+oBjbAZ/iZi7a0cyBe0+mB7VQ
KrtnDiKlZMPkeZPrWN7UX3L8DudfVKF0IyC4i2yY4KUPz9WZ3UoJP9jsrqrlsmXc
hOWLCMUZ8HYGdz3Du0Qw/VdHDYCoByxnbsHLP1wS0DwJQFu/V7oxqhCMpgxPop31
jzpmPKLPYs5pLerKG08JEF+qHAjgyoUilCXHxAXtBl1JePRYTNneVQJViCRyH4jW
TQ1ZIbQJNE34xH2DDagW6yv31jyQqby/0pO6K+gO/EhZWrivAU7bcVA4NnUfRpWN
NcIgEx+eatJFFQ6L0xTdn/yB43u/q8ioKJEcc2XYwQblrLS95jGWkCWkT4AW0aT6
TOPRhOMgICmPuZDObbu5BPnGJ964ltueeHrEZr9/TT8IjMJvbT7dsoudLrg0xF7e
UZGvnT77SLWSaXKtZxWpDGm1ps8L9taF/3XzLab6JpRgLpEn+3jSlKKwPwLnIaMg
c6TOG1w+C/Rq65VruTUQ3HhHtZd4A6pn/E0POiajOVWpsnmSvjwgGPgXnecmKKLt
ZZhQxxmQ0t+oa5eWonQioZI/vrvE2TLgsfBsZlLnpVEIY7pgwZjusKhYPe79Idw+
6hUrK1BM0KnOi0sGBUPVUGgkWJhsI8j5YQ42ebJGob2LaWlJau4aJd9bhSyt+3kL
PMso3yyWejntL5iHufMs0BCij2vzd5Gjl6Uwk2bPIzgiv/TvebB2YbIWKX+lu1Q9
VnJUSdOMOzFOdSPVbYJ6GSksgR+GqDnDm59LLHkESImm4ZCzCIbSET4U7HYi4P/6
4rtFCIs4OQoo3ec997ZYukm+2PhSlHL6+YDIzvDxIlTBxUIR1Jz/eZ676vRP37k0
dgk/SpGuDAj31Q6pgldaMlh155wDy0J+0k017smieIvLd6ekqqDCuFnw+KHUQRDA
CZRXy1TMMVr+Lld+ZjBtEvM8vvV6CY4UwyYZ7toI0P0BxB0zUxoK88lYxNIhcqoi
V6/R5R20+o7cM/hYebCdfKuLoFEoSm3kiMUCxQu6OLLwCd2TVB1LIMG6o6wU1caM
Etwi+EF4yFfAajzUEXzp07Txg5N/TElBcZbJsb26MoLrKqd+8dqPqmIL3GlfgKtS
9nbUs38POZAfOiJCudEa7Kjr+a+DXKznGWcTeLPMKXOX8/EFmUun6gVwZTHM8Q+0
UXWmVxcbPL7jyY0UlnDBghQKr0Zq6jTosub7ypE8gQmDSLuycDtvz2hTAbbpe8+o
V0sQjumEZeWo06/iqWqNIL32PFsoIvcS+iX56Jxxi+sAzqAzJgk2x3LW0UOyMRtv
hgmIc+6HNZF6577Gd8NUFQ==
`protect END_PROTECTED
