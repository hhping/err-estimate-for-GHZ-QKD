`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqvX5G1i/JrPTW6FSvZyRJQzjXchIFd8ajNA9LCWOXh3oL5nSd3X9P0Gf99KNdGr
I5WWGB6dsS6451jB+xzqHLTeHKOCMVLK1eA5wE/62iZzqkfnRk58hGxGnLyQe/cn
4p1jhm1cFYAQz1OFKz0DLemYAA0bKBX61HEIzCQfXU3mvYmc6/C+UqECLgjrGgsA
gwY6nBT/7W3TLOsvNrCRjRuZxMtIEsva1KBIidVEhP/xaGjQI03eelX6qjMod3JS
i2OSo8o6txka0XOkDHM/eqeNWw3NnLF4hxnEGxxWoCY/ojQKfiKpWwVaKdEeYAR9
R/nCJGyw4k/dACYRrV6v0Y2ZQhMRGk5dGeWy8TwPyJ3rdWIx8TCNbERn4KIDcvIf
ysJ+Olocye1lhZRVBl90oV34O9gmW3m7BtRPPqTLbs+ZxdB8opA4dwqCr86/T7ek
sfU4OPfuACBiGQ9xko7cGAEKNE5F+cz5Y+gmIBT90RhLF/tABuGlh/+N7pAIpcz0
HQq97P5fCj6jtvXVmADGI30r/dy8x16Zq1ymvrx8yeYFe6tJwXRjaJ8JPuPPhCH1
FqS6rNg/I+fhqoTg53rREkvGO+Dc59x/Ym0BqYwrF8ZEFhBwLdJYWSePnwSzeRA1
`protect END_PROTECTED
