`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIxC07r0LBBkI+KbpoY8NgzV/fG89kF/oBxvPS0qXDQTcfwXfOMN20sagoEEXpF0
8gEFE/1yrbdZu7uyqMbzLlMkEWCCKk5KZfQJ2Udot7PHCaFH/fPcSYoRVmCpCGJs
AN/veCIlaO4wmpRG2XZrt3cKkS7xsoxFhsnnhSEmlNo5V6Lc4nxL1LS9iuslC+Qd
yVXcRhzMhdT7ILwn+FHi0b5vg+JPgkUoV/anVggriUXHeD5QMO5VystSfEnzgGvt
SxUfT/0UAwTe37E4zwjoTypmArBkTWD1NMo2J8hsoRBOtl3JGJzzPs9UJX+xL3Dc
sOpJ6V/6o3UXYxxMKADLkLo8Za+/a9LiSuz6Pk/qu/gKT6GuL3SQGukDuK21erv7
j1nMN3zCV3f1waUxSuvRjuXTP9n9Y/4M/0JMatstIRCuSkl6dGA6Siky7988Q7xS
zNOhfK/gZf7ur0RWv6MWioGMfIK6jY05DcxF3r0VUfTF41nsUDZKnMM3ef6NaxQL
YiPidIVELS1Ii45mlX7a+Fx8iO7I0LJPwjraM1A711kR7OrYgTcdLN4qvWth4nk5
7jpYWPL6lquX+RgPu4QUp+7hSFNzvg9a31FI0JC60/VpNSht0z/mdL3bzOcVyJmW
hNWjUTyYgWXSo0yEUp0qO0Msbqf6O089Ig2G7aVUcDtIQcLV81DRe/ljLwWgozgq
zy8bauShHaBTT/XtJ4+/9WaKmZX0plx4YOtWkGDB4bLTL1opeTj/SuegLuzwCg+u
x97EdNIfK8L3Kb3A+8EfdwsX603r9rpWKnB2k3IqGoBNprTNBmNbpTaJ5iP4eVUB
SeO50wKyxva+euhpphF6V20y22AaSdvqIYSXxlWtghR7oI0GCh0H4Mb64sMB/Vvr
hsfvQChLYCB2/iqLZVih2zCY8ZGtP5M/I//7yoWwoAkMBPcqsUy1FWDz0rW2+mK3
yWWdZ7B79WJqm3nFs9yOTYnRrIv55lGHKI4LghY5E22sgyTZVE03GxUNTxANlmv4
aEnz5Uucaehgmy1q5k/A+i4Ifvdrt9GO6VtOS/CELvkRPia/JDfxg/KNE6gLK7xk
+t2HYlrRFdIwTsJPaL2PK69xjgAiHlzjlP4kthyYTd580Iro0rBqQjiOl2RdgDeK
HOuM61/eHM1YyfexEACUYTnXB3wUH7b2oxl3zZk+g7/OEUNCve4WCxDSM8zcmLTa
k16uDxOhQGv4ndvPPeNDUKTqhgRDJWGkORELpD0iFB3Zaem7W4ykxygX7Si6v/eA
T2dHx+YEVVB7fXAs9WKPgdtvYNt31s/fE4Ad4qAQKLBhFxuojSZzuF+tByvDofPB
ktwgv4UUZqgLrNMrDGCmdQ==
`protect END_PROTECTED
