`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vmXjqAUi3LgseKErooAOKS2rWYTgEn/g2Y0jbkBr+0p/1D+V9vk1OMQL9lcc3VJ
hsv2y3CSRkGR/zssWZaSRv8Bv14+Ilwz6qcpIf5sF/UPA6o0n046Gi8JvIvG6fm/
8TN7OiHliFoYEF6I83KRR5YLVNMvUzXDkF9vsCSQ0deqAlmMj7SFNLJRiDXmojGS
Ne97S/Nf7IrM7VIwf+saZyOeB8Dk/h57zA7HXuGTv47iSFpOAEjDtasY9VVsftpE
drHWwtHyFeXHuiUmCMitf9Xn5hA5TLkDpCPF4nhwGF4/cTo8jAJGLQVN/ggmBvKR
8k7zO1H77mCRjo5ANUCPjxRpAb33j9F+KBrdGW64mSq1a5WwhXL+UlJ+BDX+bcQn
DwqFmxrLldPgCFjSrX+zMnodV35rH0aXkUv854ZI89AUReybFZBBGSej+0Gf85jW
ovEvmlGnjCEp9sYHezQD45X/mIEmucSB4cpwfCuNiXtxLmOi5JG1qk6hBjhZvozN
1ZScyZt54sfLj24WVFZ8a3hTszRXL2oKGts+BJABGxprS/I9Ah/y47hTBYe7hcZf
/ljEzpoK+2qVDeqH5gddHyb/PGbfFAbQ5F4Ek4FBvMWxX5nwtTnUuMO8+mk7ezUC
57PuHFGaTiyF1IGSA4iV4tbG0h7F57UOSJ5tdFN4jU3LvJL0fVTb7ykUtBXCuuzs
NUUovbrbLufKVuYkxpA3p3tpYCjqmp6vJGMZAvWS5T+Y/DdRUqX7FkwaFkUSxrh+
eZOF9Y4jN0vFigt4sjq+DBs41x2yr+QbxJKpgKOdTiq+jToHjxuxOAj5xl2Ao9E5
3LZVBgITQCTMCvfOWtADhSOcKr5dkhdwSNproDjKpJ2xSZ2lRkmKGpJ5dCkiOWYf
Ok/00Gjd5EF2rdugiN0WRa0C6FKfLdytFZH+Kz8hlbRvSgctVMI+TKmztsuYkDVF
lJSHxUIkUzv3IRwdW+spz5OCUqt8+Ui+uKEz1wAzjxIj18vfmvUFtwlWr/9BbUoA
1LSwXXVERVRLBK2yvgG/vXUYA3bfwZogDbfxXGi30D5XiNfY/AZ7bTGEx7DRV+rL
d/kZiOksTki7Vssw0Fq/uXQ0gGRrfLuIEmMa6iv02wkyX4EH6l6ROznZr83hWl+I
CF83qv/4vHDa72y2sGU/VZ6GddBQ0qrefQ+i8fmo01kVJuIXEkDfViVbM86hc+ku
QtEN28e2nC44sEdBZaUDxVHExJbI4o7VukHTZmi5kVCkfhyU1LK46LB5tYdAqT6l
wzWQv1ptudjpIb81O2dOKJg5fJaNrZwbCLmTobKEAwNCKnGeTDNkNCK0BoTekpAw
20m1YS62VrcfMnAmsMaP8bTZM/sCS6a6Nl3yBzDSrITXjBQ7UauX0NP4qLfUFgux
wQWK0KEu98QRFHdrshM2D0t8UxMbxXaeYJgi3LRZ2hvg1EZSDPi7GlmzunTm3lWX
L/ZLrsz0fsyxAHoRGKAeiVIh20aXi7afFV65aiQnzsttL1SLZ7wkIZULRC064J2f
d2lDe1sxygFpvtXNSUWrBJCeDGV1r9JX4zB1/JuzxRNr/5VLTn7+XcVr+Izj9Nkr
D0Ne28GtR5fQI/zctOO8XaDUkhIGTt4UshE6K74WIJnnSOvCE5yZlrgEzYuEPUup
JfOuT4GN+v3MISrNt03wWp5xup00pNg5+BF6vrT0QuLAcFvPU4acUNtDczJHEkIP
nskVg2j3Wi6i4bh4mn8JepnckMjTqAT3yyt4HyrgCXKZwo5gNezSim2YMyTlJKVB
WwCaT7zFNlcUHOnwEIandnRsVptPgAfhuAOWKT/r+EtzSZrJHC2DzKMkvi2FTago
NDds3hAqhBjo5Bk7DwDzPQsfEAIBriDvzImCxJrz0UE8/yNN8s7/4V9aky/mS9su
WwmymcAEmwYmXebOLxle+TVytEhMzJ+OFPVJuI/49s6gT6/tvoev3OCKa2lw9Kwk
HV3ahlZbBa8szQ2c7QFpurhKN89ZwXjLwZCNHERzKUnwLHnpvJ6h4LcZREBZWu5q
ifgMIayv+PXmxnRvzIyIBHnlQpCYDpLCdXy3wJ0t0DRmdoN6z0u2j1lZYIITsYM7
mTc670dZUgEsKIuCh0KJ6N5Yb/p898dLTTRsItp1sS0oeF47+Dyv0olgkukj02ua
8dog1rMSJ++BsOBWPM9xNDQ1nHEMdmDxceuEDbQtqCBHa14TF7MaZkKPm57U8y60
SXYr2v+Pl8tKUjaYyttPGbyI5PPL4OOtLQ8rw0jqjyU8EZhMqsiUty1z/87qm37n
lxEhmOYpkFvOqW/u1hOfUUuvO6KQh8l9Zciz1VEQFXHBhkD8vjiBZIzmZ+EirbCF
nP/BsvrBS3vgQm6PGI2fWA+oiZvR6AlkWKgE8CJIXWak7VNlA2AFXneZ/8UkgaD6
/qyhsm2ABU5aeoJ2DNzwI8Xl7mxX6W2RchKsEFWwlmvifNJcO+WuTT+1VtO9b/Nl
gXsjSEBEPNiAA5fkdV5tsKQfvAKkyuPgfro/xYeuMWAI0JzLBed0TyjzRn9wjfj2
0MnkIzsjJbFpYT/M/EpYT7kvr+4Hgc3d2BfA1UElxqnMbunE/pJzvUVU7UWRRxTj
2GeIU7nZ4RLIi7XwgjZ8xdEtvtQOnU1BGDHoHKP9FYOjlEDzNKlQh46b9QPrpPYl
CotfZYdukgIqiL6v/FJvuB14AAWRTpzNHifAOBZN+iXNu5ou4T+e+3chu4zBfKzK
2RUIJQxK2QZ0a/A8/j1uzAZporwd7mPQP29zLZeO5qypmanp+hz2qMwixAJtb+ft
2tz7jbpxiiaqxpHvO8Erb7jDpAxEy3hYo7e5sKcwzy/0z0pkxrRXv3KGRRMVxIys
BEdSCFJ6iYqeId2FsHkiCF3igk6tcLwLTyfFi5YaJKJPFC0O+YyCwHfn8D9e4eyB
qyErpudZyZGOqFus3/cTQChtmRm0cAIg1QDTjm4U02EW6EChVPX4vXpZxDYQSVVL
fPjDoEl/OrSW6X14ChQT2Tkgy8+MnSZH/cKRjqlv4cCNV7zIc6W8lhLHqfxj1SXS
sAgG8rKhvMerhZsSjL/M8OzX8D7oMPGmjyuksVOcjxA1UkUODeuxe2dwRfrdxozO
9cVSKizWpbu5xsvuMRdZtbDwL+8JxI/iUJSYNjc/YzK2wuwDhUSXP1rfWi1znH3p
olt4Xn6rHavTJG2VuNnpzKQOrnDlyUBzsy7wpdtKoq+LT/LbkZilLmTArwK8Gq9R
swrthdR5CEn6KnLXbgdztPUIcZ3YoH3Xpk4LGKvkn1t/GzDdbACl7/JW/DaFAMth
RoUQAyy4cPWr/Wdq9OHWY7tKcEUerBExeC2nHM3fR0ofNfUdqEkJ9k79K2v7aaN3
3hD0XADPF8fZncbTlIEyG02q397SzMHN4co7NyE6c4Strjc1hxusIz4TbAOxBbJH
uhvJYqBveRaikOiMrfszWgC1xosEu1tluitvwHJjj/gwl9pvOONkJ5fdGyOMnl46
vnVGZTzi56QGsMxy/vtKX88ZYpklHM/Yx66EIQrCnGqENd9zstJ03wOjwfW78Jyy
CCLkDt8HYR/U/OxS8YGmtbeEWsDuQTPtu/jzl30NBItY2w3CKatsRTjGy5kfyyxS
oFuJVRFaxcJ9EZNXkKndQEkb47YwTgdURAGWQ4jZCx/mhh0XP/j4bIl+TfATeSav
ddPihURH5Z8xQN/V704N3FNC7HeFaYyG92mgRfNhPVapSaHPMm1gl2/Le7NlWRwg
z5KdV88P6fb5trCPrcoCjeZYeyEu9vgnRbMZA1C4Vt1qGcRz1K9Db6V1a6Fhje6n
KPZvjQ88WIjELIz1A9ORV1Uur4xo3sMldyS1aKI/TGv3YNxVK518RfyLwIA9FbCH
Of2P50eWGpUdbV2TPltEZ6XBw2uUyR18dfxgT/EDMDLdv2OPwRlS5Xsv2OKJ7oyv
qYB92LdH2EcHA+axOCI4cRL3J2lIZKlePLKX9sBAe298WE4KaKe2CeLPJlCtUxtz
2cVTV22DEifuJ+ZzL3A/4R1c3WMF6dORiqrRx2Q0JOBbCV4rVsK/pZqEwdbjyBxj
GP/2o/YVyWjCs94c3fzsCJrja57ozwrtnz5HuCrrZM+Weid+n4wNrf4w9eD2dIDN
SZB6+tPmPQqnbqchMvdBbCMdUb9FOicBBTsfc6hTFP7OrNumvlpF8wAs5amiZa+m
iTLTi6kdJudIbfwgFW9n9lZQSbygzAuv+kPtW9iCNjOsAOF1Z4kA5HryKcra054y
4zkV8ZMyCZtBx50UU0L7obFCaVRjE80ZYvywGN5V9mlPqrtr92tbb7wi3TAD3P1e
DEi0re0Pg3WHv+OjL6W4nFg8MZdgsaHrwZNX/Aw40eQgMQGsYa45//wq2x6Bo2Qc
QhzCmojRHjzCnYtBRZNyHkkkl/1Z4T4cQmVTuDMoea3sMyZvWKhwWsdWgVWDjDan
dnip1kIwsFc+tU1Z3Z6dYW2zwwVN4giSmWMMYFYFYi0A14+xnYvSzlSu7INNmKYt
K5qcqhBr76xWFGqZmbZwj4CAyL+Hu56NY4qKu/2GCnhGHlIlAbLXhASqbRKNp0s3
zRIXk1KVB3rLFsnZKbRaOjuQWAd6UlZ5c4rIemNBJcrzaqBAYBdLQIHmxOG8m01/
wbaOzE5ykHpngGqWpM+9rF8gxcHQ59n1bVzNNe1tle3TSkLVik//A5VHHdCWK9Hk
VR/LQ7LWid+Hp3R+QT52l8ug6rCiRviViS+KSiJJAxXZM7Bv0jlAtU4HgCmez7WS
tvzck6yGs6wIbfQEo6XjYz8mu5D6Ll4hl5vWncsKvR4Quhojnk1bWqOaAOQtvcIF
paCEbJBnFYMXjOW3QFUHPdhW9CsJRNY+OZ9Qxy3zM1bbqPb2L8agCWk+30Fz7RyR
zoLtJETz0ieH8J3qvS32RdsY13SVlUgpZn5Ylj8r3Zx9RvDDvVJwURibm5XGM/vQ
Pc6RiZDdn4pPnc6BGoT3BYh6nvagtkZI3yuBx2EE0neCUEfGcQ+PyME5zF2Z9lLx
PxYokw+bg+jqnfvQIZwTTwhP6VMG+UDHRYn/r5oU0NmbSW3tX1Gx4joXJ36ouF1B
JKnpWLBTRo3TXkfrLe+ugwgen//0bVjqhqapIN93pUJQich0UWoOGHmqWQyxkLNx
yo+rC0sipvJbTFCvykPqQrXaQPNISnqSB39vEwXUg5nlfCKYtkRl3iHiGXXx1ye9
2hEdJ3nrAItK9Cfcjubi10nSr2gXUMzchG7QOMbkyaIZSpfnqH1CUkMmA7KC9V8M
fAUVbuFzfJhaXlWwMd9kmnDZAzycbVqWdIQ9GOsdSRHp1TeqoGE+UnhBK5wPGzuQ
r6Ahk9vUz0BpmeCetkDQ+4K1Jo9nTBdow4hc7AoSu/F17xa3+YZ2j4hO2cu/WaRt
UEKf8l8/dQ7nokC5wHFIxBlcBc4bNjTcpVny8RjU5sETvzCjpot2EaOWTBWnAWGY
y7JFNYYTWZncsnvXzez2glQz2qPfp+zTw1bE/7jPu4/sPaF0b/BwRPP710VgqX2x
p6FEJ2n+E8T9ccCcRO+5kANA34cvjgaLeLAHzxhkts2228O8sWyaTi7c+S7RDLcQ
/Ryawz8tCogKswPU1BfgoVztdfsQ7ies1QZfkSb6NAhqNm7US9n8qvPjapkWRzMT
GxqgiaIDdE8Q/voLkKYAg6ljqx31KoMxw69vooHxmERoZzW0FSzCETfgbvAnrIyb
CK1Ix4J+O0RsYZRRWLQlUUkd89yECAL3o+fSe4ERCBJLOtJAOpGxCvr+f09cyyT3
u+glvUraU6cvBacia/XfNEY3JqxE8dPDU9jWbbHZafJotbUXoA7W2gzGAZjyhyUV
5DuMp9gLFrP06AAgNB5ZLTz4G/lVvbFdyoNXRufwJCYTOQymvQVcjMJ1QTSCY7vB
5zi05L9PdHAexgVg1vGV2YcShQBqKBaWWDb8lO81U4P3CmIgzTPP2YQdVjZ6D2xL
osl1pJPpdxvVHtws6U9GntWKPckfZw9xoAqNK5tqnY3BgUtn4wV3B6kJm7JiBTlY
UQK43js4zlYvFcEdxvAHJuxJrWNKgkxiLrwCC5Gs8j99Dp/DUslyU3ni9Z0wbt/J
FLk6u+Vq5wOKP/gt7PVf0k0q5rc+yurNNnuuXc91YwQNftGziL98935igNDuhBez
5iwf+juGPrIsGpubMlEyf8+eacQG1A+Wu9ghdarNRK3QGIhrDx1U5SYrYgX3S4RP
yoLKvpYjG9h+o/NoXeEjE6e7J4VOq9/luVoT67laBL9i+brpwIxzBs3IXkj0Ay4Q
ciXK+BMYAZ9ogo/ZE+tFnPgn0sbJB0OMxXSzePlFRvElukkOqL3l2gYcxmz9cvtf
q83wluEiiZJSHNkvNBGADeG0p82iv0cMOkX7VrwwnOT1UKroRUYP/m0tXmgprYoH
htc6RTEuNdujZVuUIBjo4k1liT3fw7cJBJyV7GQz9pQJDGZpooJwYX/c/wkiKG1E
AV+6yHnKJeJPElCnn3AyOV05yoTMS5Z/YhjaaqpFw+M4enbolnGb8H+QtpJFapUK
8RsQItdwo2AVb+E6bb6r7lRulIFHftpEWTLME/7LKMOqkJnfKLJgnRIa0VTe3Jgp
aZ56YvVkolAW31bJBJ6SItsgnCnzgi1snANtWO68L1jMnAlShi680sG6tPSXFPUn
BwzJb+i0gEx2Jk61qqfaxvvG6t3c6YU8qnj1Xgl17r3LVQnd9UjgFgH0yFxj9lfb
g6HbuCiJ48GxWeqZJjEF7d6SnRcuPxv65pSGlQL3T/s9PChlNDSumoETaVr7kGmw
f4U0BLczuvFgxLmUv60CGc9A8nu50oFRkeberEznmusITchxd88bg3caYl6w9XAB
5F49VXr6R4C102Q6inhggzqkwcBWeNM7k2ZF+nk1wE1urNJH1HQEq1/HcEhjjKIf
CkekflAgX9A6PusBbgXJFkk+90q4BJjKHxW3EkhdXRqtVWvvuGJ1R7B5A0/IHnty
ag9rv3grE5FiRyDp+Rm90mQoNAEjsXAoYhxEFfYcynbHClKKWsRPEfaqqzUyn4m2
ZEAW2dBmYjIz5IE0ulftEosu8rivt0oums9D2pRwDWKAm0yiiW+kFiAqKzzvCzYO
a+vr3O7RLVxzgR6OvIaZExBPrMLTaxkwe6zJdqLNHXyUpMZMP160r0aKKqC8mofN
5+ZNG+xn+SbgdovV+pNsxeNXXor4GcIow4g2Q3J24Ozw3HrZKpujsiKqj3AJ8RKA
WBF0xEYxd0vcsi6O0jaPBEfW89qzpFv4n3U4W9LyxqvxgbpJyH6wU9kXq+YJZRCz
0629lq7VPlpfqlzEag9zYdSs//8r11Sp+zXWkJhRIdhnMQSIOqp6GKDtD4sbcsPs
ddYB/SRFBnV+jfb4LridFChv/k3PDZXDQHOUb+kD65JPh/7h9LByExl2hLcXFz7C
QnbDOKj/vJJFsIg95OROjUP+JLSKbsvWi1UmwAXoe4jiRaRlE3jUUQ7Z9HPPwA0z
zuTQrWjkvzF1F2A4+GxgN97h+ePl1KfQIyBpKvvXwq41M6T33uGBYMcwzH0fU4Yx
KJUY8flBsUutdIJ6gm3MVGOu3hPHXg6FMqtUovY1rI6Se6nsezC9JyYSxmlgbw/M
cgheHh4ZwVaV9dJv4ZKaTNctJtqAVKPvvOU6CDMc9GiUeer4EARdrXRmagAAsUgu
1npf2VsNyZ7IFD7QU2Xp3uq1d17Tz/JWuhTK6USWYcvw66XL7C01iz9mgi25/xEN
EQZpq43zlAm8/xOiX2c+OVEAJev8pvNrq5kBxkh0b9+xjSYSUFT1ulbPZWJYdtKc
ux3SOYcGEDr8LrGMKKD6xl90t6PWM3U8/sN005kn2zKS3vwg9qEQ5WSGMdBUKojc
g44zPCh8jdQbz/W39+ENqCS7mJSrrJWbhG15FP7PDKDFTTELzKRD7xreyddQP+Yf
CmgS4QiRvlJtNfnaxWn4mMVmJe9SJOvVk0XVhoIHFe5zMYZMqQxq0HEzEUbFVkG1
ugavyk/gF250b9aM/xxujHdre02IE6gxSUadTMzYVXfnoFQDcn/H5V0wzdgQc4wA
6rZ4hTWgZ1dY67gKEhIWpSAGlSMVXcrGs2CEjnb23RubbjZg9VEmUCQl4Q+FqTf+
+wJTFZnNkHj0Wnyy4KwOvDoc2KcWRdX4duDDMpssMM6VX9feaszwfQzq+zroljS1
YynF4meenyDvLzm/4wA+6dNrSsu4bu530WKdhPYUKYu3gYyiKHYv/pggrx/7c36s
PPp5gKp2BfJqB2ht/xANrexKm6qYZGFwvpDgYjhFWBjsqi1Fku0WqwN+zSO2gOoM
VNjSTtRMP25jNkzAftrU74IM+517A9J43YxzsqnM8sjwdMXByNYRVsH2xbzoEztG
SwVX/KrRXMqoQlbVtyz4GvpXtZTBreJE9Gh7jWxLqvQtISuSkOhPC+ZV0WhPGdwd
CUzHWzN3+KCjxFgUfbDShy4JGkRWU2ZIeNlhQ5z80MFDEXh7wbXCa1wTDPaT8uM6
6pk/8ss1p2QoUmusdWKAwfZSzPTLIDKmUz0135c+/b0/IBc5PJRPtbU38k5n6E+8
PGNc4zrszF++SyJEkKGIBf0Qp4XwoqnDL8jyekgwM6ispOL0gO7o0T5YO79xJ9Ms
MSaNqWXkzP9eXrCCslTNEkruKuyx8Kt2/XmCuy0JlgZYElZLmPkk3jaulwsFHP2+
fG+CrPlA0wlbcPpzXXP9DoTgMTlDaliJ436tDesv6YGr6/eU7TSZTictYtmdb8+A
qd4ErvsbqYDc042TV34wbwIh1/B1IlQBKWy/v0I37GVuDaab2oeCL482eLW1Lv5J
Ky6cggdbzWC+l6AWvReHARMPSiZ5LNywyMNFRBjVQXvOxXrZa2PNnQKpWfi6KB82
MLc5V0w+IWTycsRse6v3KDCu3++3Y6ZUVh7SDikAsy8IrCAdeo6MsVWGoJ4LNXKP
2vSga/UonlQjhfAaqNAqyndNA+ApoNwSSbeAa52aoTIbiUO6viNxPAsVqYGGIKfO
mMcI3CAlI3UlJnCUF+ThXOa/IqtEJD6OrsbzknFxXN+lH07me7o5ZXy/b2otJtGK
uTjB7Sw3OiZOZ/OTVaB3ExOUN9uL2+Ct7XdH29RIJ0Bj3T18cbh9wZp1Wdupszlh
g8gksmCc6h8Esjwc9PW0nq3MeyuXzZp3IbcsTgSnuCFS6eFZ9EwDOHXmXX/P46KY
KC81LZsAdPJfsD8A4QNTFKYzPHYmLpjz/WeIkN1hIRzJz8OQmnnt9nXazFmTkedP
d0q2xWMuklhkx2hKusnctekxKpua4jDT+hoT4gviDUphOA3rdzbluWZHQvvcg+E1
mJgD4aceIMEjqSkcHX4E7vyZpg0o0hnfNp7uCf6uKYEIWW5z38rr65CAQ/GAUGJs
g4cWfEWHuZpCb4QD2wFX2AV9Po6mmo+Q8Odg+tappyYHpRnnMoZawOiQml/wWXQL
CFZRjHjTqyCZGYl8e63L8GhDgI6UFE0MnhlddZrg1dVRGiIMO8uE3la46L5VZopf
CCo9J/uDlrAI80POYe5TYmrmxLeJYAPF6ktE/O67lVNHDabTkw4QzC1oFtjLlga8
cGGVwtD4F8TbpH/+mn8CkzqshDyexfPrXn23u7Q7me+xJrxWfNyIxGxehzHT+2uD
SWmyIeoYW5XE+NlKvQvqo8ov7X1VrpyvRZI5jJQvtXAt+SXYmgkiVjpnho9cTur3
POVt6kutajzyfwo5SiNDu0qvpjU0UKPre/A4wNSY3t93m4KPG1aIEgbR89RIrgkM
PBFXizFahW9RrssVHJUQqTbjXYxtOylMGy9ryJFHlqbpdCDowWL3PSuksoaocSvt
NV69jagG9daw79kNKUzOSxZDozq8Ua+K4M5aFwfCnC37JEENC9ELLqnCe5F4NpoH
RNFSGYXEt8jaLmjnOSskok8fgna7CE+WKIiGzBLwZhd8yHK/8mXPGpBUROH6wNVW
JWEHKK7ECsK5PMrNYOnZ0fFlb8Ne+M8JTKbmLL/FZdaJjGabcyMFMWJ6VUmOUkzO
EOyVp0LOIurz3q5YrY1Z2p/mCWCFQ/9KU9xrwvsi+2n41s6s2qn6V9Ot6QB76y/c
sZic6XTaPOuq3pyWFVLN74g/HvvyxfWNFysgRijBU63zSiim4YdhgHOyWwSWM6Ik
3iVIhNNkzHFSfSyjrIbYwCiRsqoYhaC5Ffw4R9x6FqFnCJbt+DIdtkJxFfcnBDLM
iwzvQMGKv++GBcX8Vraypo1ms3eFoex2f2rOMCupGzfuKHQRwVZSM7xkUnVWVGcu
mj4HlGwwvp3GLRbwvaiwUm/vJ/F13w+jMKQTvaXcYNhc/kmaRqwW74jVtos4Yi4I
70TpdexZhzcBxhodLzRHwwGPjISXswbpP4tCQ6hFHhw0/ZLDfjwgw8lNglGowBr1
xVDZyHEJzBDzOAvooVLlndwPeIiK3Os25wyzwBRiVz36P1e3QqQK0w9spGhws2vc
kgJlfgESCqqEfBCjwSQWwykcssnqWIifFbGayCv995ZZsZHKmmgdbgeL64YZjAcZ
QYG35Y0+Cy4vlnQQzzEj3gdnmBhuTxjLHDspCm53ZvsL38dwWK35hrM1OVyd7zcT
vNtXV2DRnyNVEAxWLDkoWTZ+QD/VwIvM6MkDWOKF8E3itMXrO+HeIFR/sU4ILdTd
+i1I9zkc9OZd2SXqZiT6BBIO0jMUB73A6sLMHf+L2q3ohNw/5t1kOjf/u3kIZiy+
qYU/JmvTOK+8/I1bliDVhIyQ5kbBjlWEzWbhymcJqnWPL+W8GogxnJADMvLKfjNP
17yVC65RUQ5qALBnpBPcPg2ogAcwVOEOYdggY8i9azdWrYs///YJCvMtooHY47Bj
hoZAmOno+i6tXtzkMon7V6tC7Z3WYuin+PLQWkOwEJJY1dMOab/t/rPIC+NQbxbW
6g8pCN+LVgTdzfc29KNILMaSpEGrOoGmIE3eBPVRC/2mC8wh/hfCsY7rPGAcHdLO
rIP4M9rVr5ZzTQ9yF8euOCz8hSFhVdMesfvw+zS7zYjxMLSroOQy2iivVEdmPuJp
jhAk6YgGpS3HmJrJO+ONYR1eeyDxaRT9OPX0aNMzvnzsOoFSNI/hPhf4loX2tkwg
7KzX0j63X923wYLU2qtqJ8XoDgfqnByChLV2BdiEPwG6MhoGieTLPU2hBggMmhj6
OV62p9oY2ByaSUfsXYR67ov2BtDThX36bvgtXH0IZOgyuss/q/FJ7+5nYyVFNEfE
q567jlzy4Dvs5NtAfoTjkHU8464srGHelWbT9Y/dqPycc+XAG/tp0nF88BrsJM8i
4vo/WzDM5NKnzLZ6TnInlMWCGtAHLLogfNS2bOBiqd6OZu2fyfi8xPE5MEeT9gvV
D0bSrOz5dPI4YxY7HnxI95KUCEHrSyEVU8FvYj7i9+5PfN4m4FfTNCMC/1POb3zj
+lwIfW5KbTkW20pXjHfrml7cVVTkyNTffO4doVVkiXbkjnkRoIbdsXV/4Pjvb4Kz
`protect END_PROTECTED
