`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99O/Nm0YtdgmHTAMt4FpHU09uSej80UUACxSXmSxDqeyvAWsRP6Kgji2mQL78dyy
eVH2a+O7FYAYn67ujqAHBNmNuXglHUFOx/k94sribngdGN70aHG6R7Xg3VoHjP6Z
cvIaRFQaCKlO87v4hD8iRv1t6TdKKIzd1qjQCV8Mq66uEIowXre95tWZhbb7rnfV
htxhJepcjR5UTeW4FnXK0RKMvJXV2wNHbQy9jHOAOK6xwG19JgCTKQPLhTzHFuFn
7VGuHh68G9nXg3Dj5HJxAtF1HgUk7WkTNwJVak9G3ZczTc0+WQfFuQgnRxFRuOxV
bUwtSN7cEDAnu27isB9a3y1nWMWjy3fi8q4iGjTssjxdM5zcrlkQn4i8hKaxDhap
T9mm0iAyEQAqcYl0G4Y/wRbs/IYUTo6NUx2awXzAhvHcChKuYg2CoH4OaoHTGG6J
oQAUMyX9JIiWGDZsgZu+xb5pAZAutTp3WOGEfyW64JJxHV3EzOAGMTMu8frjgzfm
w4+9rjNGc26qH0EHj4uwukQgiZMN7fPaDAeNFTr+XrEC6xTp77pkI5R78Z4KKR6Y
z8QshbuBRttj6qP62uZqPCZNw0Nju+o/iMKe0gGfB4kb8r4m+6kSqHNKbs66ZRXc
`protect END_PROTECTED
