library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_aux is
    generic(
        enable_debug_info: string  := "true";
        dprio_base_addr : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dprio_broadcast_en: string  := "dprio_broadcast_en_csr_ctrl_en";
        dprio_cvp_mdio_dis: string  := "dprio_cvp_mdio_dis_csr_ctrl_en";
        dprio_force_mdio_dis: string  := "dprio_force_mdio_dis_csr_ctrl_en";
        dprio_power_iso_en: string  := "dprio_power_iso_en_csr_ctrl_en";
        initial_settings: string  := "true";
        pm_aux_adc_vref_trim: string  := "adc_vref_trim_4";
        pm_aux_atb_bgbyp: string  := "atb_bg_ref";
        pm_aux_atb_en   : string  := "atb_global_disable";
        pm_aux_atb_mode : string  := "atb_default";
        pm_aux_atbcmp_pdb: string  := "atb_comp_power_down";
        pm_aux_atben0   : string  := "atben0_disable";
        pm_aux_atben0_hssi: string  := "atb0_hssi_precomp_open";
        pm_aux_atben0_io: string  := "atb0_io_precomp_open";
        pm_aux_atben0_swap: string  := "atben0_swap_disable";
        pm_aux_atben1   : string  := "atben1_disable";
        pm_aux_atben1_hssi: string  := "atb1_hssi_precomp_open";
        pm_aux_atben1_io: string  := "atb1_io_precomp_open";
        pm_aux_atben1_swap: string  := "atben1_swap_disable";
        pm_aux_bg_powerdown: string  := "pm_aux_bg_power_up";
        pm_aux_bypass_bg_voltage_to_iconstant: string  := "pm_aux_normal_operation_for_iconstant";
        pm_aux_bypass_bg_voltage_to_itrack: string  := "pm_aux_normal_operation_for_itrack";
        pm_aux_comp_minus: string  := "atb_comp_minus_disconnect";
        pm_aux_comp_plus: string  := "atb_comp_plus_disconnect";
        pm_aux_dac_atb_outsel: string  := "dac_atb_out_off";
        pm_aux_dac_data : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_aux_dac_data_sel: string  := "dac_data_dprio";
        pm_aux_dac_dmcn : vl_logic_vector(0 to 13) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        pm_aux_dac_dmcp : vl_logic_vector(0 to 13) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        pm_aux_dac_lst  : string  := "dac_atb1_disable";
        pm_aux_dac_neg_trigger: string  := "dac_pos_edge_trigger";
        pm_aux_dac_pdb  : string  := "dac_power_down";
        pm_aux_dac_resetb: string  := "dac_reset_off";
        pm_aux_dac_tstbus_sel: string  := "dac_tst_0";
        pm_aux_dac_vouten: string  := "dac_vout_dis";
        pm_aux_dac_vref_sel: string  := "dac_fs_full";
        pm_aux_dac_vref_trim: string  := "dac_vref_trim_4";
        pm_aux_dftcmp_pdb: string  := "dft_comp_power_down";
        pm_aux_iconstant_opt: string  := "iconstant_opt_50u";
        pm_aux_impctrl_tstbus: string  := "pm_aux_impctrl_tstbus_sel0";
        pm_aux_itracking_opt: string  := "itracking_opt_50u";
        pm_aux_lower_limit: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_aux_refclk_div: string  := "refclk_div_bypass";
        pm_aux_rx_cal_override_value: string  := "pm_aux_rx_cal_override_value0";
        pm_aux_rx_cal_override_value_enable: string  := "pm_aux_rx_cal_override_value_disable";
        pm_aux_rx_imp   : string  := "pm_aux_rx_imp_48";
        pm_aux_sar_atb_insel: string  := "sar_atb_in_off";
        pm_aux_sar_cal_b10: string  := "sar_b10_cap_off";
        pm_aux_sar_cal_b11: string  := "sar_b11_cap_off";
        pm_aux_sar_cal_b5: string  := "sar_b5_cap_off";
        pm_aux_sar_cal_b6: string  := "sar_b6_cap_off";
        pm_aux_sar_cal_b7: string  := "sar_b7_cap_off";
        pm_aux_sar_cal_b8: string  := "sar_b8_cap_off";
        pm_aux_sar_cal_b9: string  := "sar_b9_cap_off";
        pm_aux_sar_cal_ctrl: string  := "sar_rambit_cal";
        pm_aux_sar_cal_mode: string  := "sar_normal_mode";
        pm_aux_sar_cal_refn: string  := "sar_refn_sw_off";
        pm_aux_sar_cal_refp: string  := "sar_refp_sw_off";
        pm_aux_sar_cal_top: string  := "sar_top_sw_off";
        pm_aux_sar_ckskew: string  := "sar_skew1";
        pm_aux_sar_cmp_curr: string  := "sar_cmp_curr11";
        pm_aux_sar_dmcn : vl_logic_vector(0 to 13) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        pm_aux_sar_dmcp : vl_logic_vector(0 to 13) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        pm_aux_sar_inbuf_byp: string  := "sar_inbuf_en";
        pm_aux_sar_insel: string  := "sar_input_off";
        pm_aux_sar_lowrate: string  := "sar_normal_rate";
        pm_aux_sar_lst  : string  := "sar_atb1_disable";
        pm_aux_sar_pdb  : string  := "sar_power_down";
        pm_aux_sar_resetb: string  := "sar_reset_off";
        pm_aux_sar_tstbus_sel: string  := "sar_tst_0";
        pm_aux_sar_vcm_ctrl: string  := "sar_vcm_900mv";
        pm_aux_sar_vcm_en: string  := "sar_vcm_on";
        pm_aux_sel_fusetrim_cramtrim_adc_dac: string  := "sel_cramtrim_to_adc_dac";
        pm_aux_termination_cal_ctrl: string  := "pm_aux_termination_cal_ctrl_0";
        pm_aux_test_counter: string  := "pm_aux_test_counter_disable";
        pm_aux_tstmux_statreg: string  := "pm_aux_tstmux_statreg_0";
        pm_aux_tx_cal_override_value: string  := "pm_aux_tx_cal_override_value0";
        pm_aux_tx_cal_override_value_enable: string  := "pm_aux_tx_cal_override_value_disable";
        pm_aux_tx_imp   : string  := "pm_aux_tx_imp_48";
        pm_aux_upper_limit: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_aux_vgen_pdb : string  := "vref_power_down";
        pm_aux_vgen_sel : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_aux_vrefen_minus: string  := "vref_comp_minus_disconnect";
        pm_aux_vrefen_plus: string  := "vref_comp_plus_disconnect";
        pma_aux_clock_select: string  := "pma_aux_clock_select_clkusr";
        powerdown_mode  : string  := "powerdown";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        xdprio_aux_wrap_xdprio_aux_cfg_dprio_sel_core: string  := "avalon_access_from_uc";
        xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ximpctrl_pm_aux_impctrl_sel_high_code: string  := "pm_aux_impctrl_tx_sel_high";
        ximpctrl_pm_aux_impctrl_tx_enable_eos_det: string  := "pm_aux_impctrl_tx_disable_eos_det";
        ximpctrl_pm_aux_impctrl_tx_ovwr_ncal: string  := "pm_aux_impctrl_tx_ovwr_pcal";
        ximpctrl_pm_aux_impctrl_tx_ovwr_state: string  := "pm_aux_impctrl_tx_ovwr_state_disable";
        ximpctrl_pm_aux_impctrl_tx_ovwr_state50: string  := "pm_aux_impctrl_tx_ovwr_state50";
        ximpctrl_pm_aux_impctrl_txcode_sel: string  := "pm_aux_impctrl_txcode_sel0"
    );
    port(
        dprio_addr      : in     vl_logic_vector(8 downto 0);
        dprio_clk       : in     vl_logic;
        dprio_read      : in     vl_logic;
        dprio_rst_n     : in     vl_logic;
        dprio_write     : in     vl_logic;
        dprio_writedata : in     vl_logic_vector(7 downto 0);
        pld_scan_mode_n : in     vl_logic;
        pld_scan_shift_n: in     vl_logic;
        scan_clk_in_impctrl: in     vl_logic;
        scan_in_impctrl : in     vl_logic;
        dft_flag_down   : out    vl_logic;
        dft_flag_up     : out    vl_logic;
        scan_out_impctrl: out    vl_logic;
        tstmux_out      : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of dprio_base_addr : constant is 1;
    attribute mti_svvh_generic_type of dprio_broadcast_en : constant is 1;
    attribute mti_svvh_generic_type of dprio_cvp_mdio_dis : constant is 1;
    attribute mti_svvh_generic_type of dprio_force_mdio_dis : constant is 1;
    attribute mti_svvh_generic_type of dprio_power_iso_en : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_adc_vref_trim : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atb_bgbyp : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atb_en : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atb_mode : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atbcmp_pdb : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben0 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben0_hssi : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben0_io : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben0_swap : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben1 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben1_hssi : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben1_io : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_atben1_swap : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_bg_powerdown : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_bypass_bg_voltage_to_iconstant : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_bypass_bg_voltage_to_itrack : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_comp_minus : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_comp_plus : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_atb_outsel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_data : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_data_sel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_dmcn : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_dmcp : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_lst : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_neg_trigger : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_pdb : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_resetb : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_tstbus_sel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_vouten : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_vref_sel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dac_vref_trim : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_dftcmp_pdb : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_iconstant_opt : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_impctrl_tstbus : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_itracking_opt : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_lower_limit : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_refclk_div : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_rx_cal_override_value : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_rx_cal_override_value_enable : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_rx_imp : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_atb_insel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_b10 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_b11 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_b5 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_b6 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_b7 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_b8 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_b9 : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_ctrl : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_mode : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_refn : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_refp : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cal_top : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_ckskew : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_cmp_curr : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_dmcn : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_dmcp : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_inbuf_byp : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_insel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_lowrate : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_lst : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_pdb : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_resetb : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_tstbus_sel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_vcm_ctrl : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sar_vcm_en : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_sel_fusetrim_cramtrim_adc_dac : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_termination_cal_ctrl : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_test_counter : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_tstmux_statreg : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_tx_cal_override_value : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_tx_cal_override_value_enable : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_tx_imp : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_upper_limit : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_vgen_pdb : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_vgen_sel : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_vrefen_minus : constant is 1;
    attribute mti_svvh_generic_type of pm_aux_vrefen_plus : constant is 1;
    attribute mti_svvh_generic_type of pma_aux_clock_select : constant is 1;
    attribute mti_svvh_generic_type of powerdown_mode : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of xdprio_aux_wrap_xdprio_aux_cfg_dprio_sel_core : constant is 1;
    attribute mti_svvh_generic_type of xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr : constant is 1;
    attribute mti_svvh_generic_type of ximpctrl_pm_aux_impctrl_sel_high_code : constant is 1;
    attribute mti_svvh_generic_type of ximpctrl_pm_aux_impctrl_tx_enable_eos_det : constant is 1;
    attribute mti_svvh_generic_type of ximpctrl_pm_aux_impctrl_tx_ovwr_ncal : constant is 1;
    attribute mti_svvh_generic_type of ximpctrl_pm_aux_impctrl_tx_ovwr_state : constant is 1;
    attribute mti_svvh_generic_type of ximpctrl_pm_aux_impctrl_tx_ovwr_state50 : constant is 1;
    attribute mti_svvh_generic_type of ximpctrl_pm_aux_impctrl_txcode_sel : constant is 1;
end twentynm_hssi_pma_aux;
