`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yf+HjlwEVIRI49pqUgbTXbX8INUaaONWKuPjRhguKIOeiVbCrCtMbl9Wgefw4HME
/WW2sVnsqJI4Aum7Se82J7EtsXg3vUadSH13/Qrdh6hsAgQMl3InQKE0ESCqpcJe
zCyxJx16OTODNND5tx4150nLBu5yc4JPj2UGJX2gUaOpeXko7E7eXrSYrBh4h83R
OEymXJi7txyAnYdLt3d5tU4fxwEzSS3RMsf5OlCKCLpEqB72McWg70drufeLoyN0
bYP1V+RVDfpH1eoVsSSNQcK6/rGgIDoxpLDmpSD0LUUqJ/XwzOleEF0jFD/8Cbrq
0jRYvmnY198+eYbeUBDp58UB8HRkmhmSEWGwOcOAa/epjCgM5BYb3IFzjR+Bx4+u
7h4ji1enm10QYDm2yWORo3KJqlA5lyJafT4A8DARf65sVVqLROs8ZhjeWKqxEjzz
OSU5K8ITvgzJ8gZ9Hf6E/Aopq3v6mr6xEPeGHkKWjy+JyrS36D0G5fiL+jB5eC09
M8NM5mX0MUPd3zA+j1UrMrgVrlHlJhnIZrfz7LcBC+kbeZH+aSTS+5YKh/cxeAJa
qyxu3Iqcv5AE80zwVdL7fjdrvaFhjlZlwKY0BDf5JfzvlzH0BZi5XJoWDQkgkGES
CRLSLIZzkZ7CVbf4j/fd0eXmKZW3RtaGLDZh0VfpIqIuPsIBQHibRAwJil+SQGaq
NPFWt8KJr78yjh18NERGORnwO2V8VJbeiG6/DIoEDo5izg60EEZVrL1NAwGaKHJc
a2BXiSVzEoIxlaYfBktEcNvfrLvz5OdJCJzT417QBNMKVGk4B7bG8WgUqOGDypYc
sXDpHcEYAIxsuMMciaktZQ==
`protect END_PROTECTED
