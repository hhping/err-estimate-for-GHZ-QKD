`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2Bt/r999Wg7mMY/Y6D2Vqc5hhAP8PRaABpN5A16+3IV5C44k9+x3W/iRzoNfD0f
0Ve9wh4z34dovN67eFL/hHTXl04PONKso6ifXgyXunFEoQMMAzZrgvuG4/rYvaD3
D7fXFLucqgYi+3MDihqpLp0KBAXhtyKiw1I/YdaC2H/7lr7Mkshdpj57nD8ErvSu
fues6MuiCI94pNPoQ/w2BMkOumInuLdgJz5Z6sbUVX6BoGEoSlhfp7xz10flBy5n
nUCL4b1ybAWQeB1gFyKnidJgVlQ/CdeYszxLKC2bReyldgazCGPUD0MQOW6KewHy
M9yRfnHk7U3hN3kkq6VhEaynjn62ZPFAA3QLc1WCAZE0djyfsvVCLAJ0bPC09QkQ
6lXi9T0ilFiVtSxp1FjoZ3K7Jxlgbboj9WYYH2cZn4bFFH/01LRYYTlBH66tr3ES
ETwqr8AQR51mcPTo/q+F90MBpVTdVKpGstn86kGpjgJu52V4wXx6PlMEnqoMFCtS
GMv1j7HvcO3nhyXIMM87bZReQQ1JZbdRoA4Qgup1Leuy/aDP5iPLzBmhFCDv3OcR
M3W1kDk+KBd9M524XpBkpR56+z57CMRmeCS81EqYNxxRB1/VSFad5paI0oJBMgo4
IK2WknsV38V3d/5/W70WY+LV3Kzwj3O+IYUKgGkHqoZNj91ExjDGoqS5pXkuhoFp
azcfehvGZJR6LOe1WpBHJnPV9WT+o2ZEldXXkJ+Wy+gYmjUKMPyhTt079okQ/k8i
L9bYbH8fFJCWFkHY8esCy8GhS4r+M8h8kKZIXmNwRNv1copsh3g45CA/t622w9em
cdwiLduSfIcdW8vf0TOM6ye7D+gjmPPUj5+G99jSLxPxXW1SCS/MwLU5b3OJOV9F
M0Lym9mjY4JSHjk9bsq/AWup1DfQsrSt1QVvYgw1iQbCijJejOpBLVG1P1X3lQiP
ANQN58ACN75OS1c7Ocx6WVS+jkdMP/xAWRdW3P6ZmuJ9rwcgDFfVJNQe/P2TkVlT
q2rEdoalcpajHgtRYTrk3oYIxlFmutl1HijgcdI1y6nlMMdd/XEfX2HD/UDLRrUU
+oA/yzbyQ8Rhn34QIk1WsIAWvTpCI9rv28j//4p8pmjqgzMz/wPLQuTOQhQ8yzPZ
ixBJS+tMQvQYQndvLM982u74H0FnL9mdL37zwobJNnuFWxjAzPBR03OXoynecNMv
W9dhbED/TXGP+yyqWQyCvr581rqjoqTeXDgK6Xoq97yDtVFLpxPJBmWcqztDNqFa
I2mFrsHk8H0fiWKkWgCNWSQKiLg1frVoYAV3fi661qGB3oCfPW96DmzyCw6k37rw
//cqFgg8eQzRQs1CcUw/hx0gYm9qBhBmbJJL1nS+DPZsffHXsyHOJMlnySWoyBde
xrw3nU5D7C6fyIjhkjzwPVyP8vA2V29rfiSi5NSLjFaZh1Img0Xi7eqEb1T5Q+F9
k0qt38ETxp+HiTprh5sip/HWyrBHa+74TAoKR0/9q70pzjNDVtrrJwua2OuItBfO
hEhwE7tM8pm7SVSmlhlc4ffvsNQhwvQwjW3RFXeyZ3kfFhoF5niFl5vaT+UZj5JT
Gm1xG/jfUOPmXCbeYhDGkh0l3N5bc/HXuPkRus2w+YwVirZIOmlaGJYXMmbB9Mbd
FjIizk1TminR788ELH/ZCa+IXPjsuy7ADzU8C5K0eBC4Rjri806FWCw9zqpnCXPB
g13u18fiFBmHjAS2Iqt9JpOamrg3wzGXnDE2nj7Jf86jCsc8VlkDAuO/qvHSfeJR
rVAPA8qZqC+Fca37pKA2cdNQX283/TQ/YjsGsWoFO7HeqV7TPcgctf51wYuRAxEU
W3fkKVvzZWny4WCTJc22Gl9K2Uri/VcCi2gzXjCHEUaf98OQTBnmkGwU9Mo50f0a
NRiECibLwewrQGvWlBPJ8FGvNCo8/WQ/295mFsgkZoo=
`protect END_PROTECTED
