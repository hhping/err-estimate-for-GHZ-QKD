`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yjKGH2wbjtR/EmQf5ZvggKDnRyzzflwpvK/G4DhKCFJLNMzlORjjMH0A3FulraY
8PugbgwuabbO7aM/BvhKpxkkxVTuaFcORXM7Vd8iMy9fsm2f+FvhEdU8xerwR7BC
M9vFXv1Ln0Mz+M+W/VK32xH8rqPRq7A1uwNjlFs7xgaKnxVoGoENv+xoy+DpyOmE
zfdgzi0EuwNVhJOSjP/Zdsdj66FFtpy+rygcfjF6mIcZUNeq/2uRB/e7aMz2ey6/
13+HhWgxwko2Px1E/L56rx720DNas8Rs36IM72THqhNGkkTH1lYMyvRt6xr1zqro
tm+fu8FC5Ak1+VdBuZ3VrGRm7b3a9TJgO49c1DB5LpESLmmm2aYZvhXrrt5fIj19
mNXFXjk2mT4hEQYha54eocDmyD9sJiZk3iSkHz/TM9rcAtul7R5J4gQY/5pXxyU5
HUq6f4eOOTeeQdNKwt9PPCY/ZkQjA0oNOlPM2G+JhAHwpUsFej/545k4HCo0ASob
rMSfB1J4F7Enh5D41EWVZa9IWs6+Vo/q0KkLjbIRNhhvJjuCcQBuIPkyg2n+/R7c
k/yHWjja/EEnd2d2HyeU9L666fr6xkKoVjq6Fy3V3f/m1rCrVQ68s85k7LHz9qmr
YROA6zxO1G9Fk4OmCSanAW66HpjVmbgMuMKlwoexiPUlhFyUJpdUiNsISAVc+F7r
QoMwQwp2lUYl3BV85txXJoLS0u8pKWh58RKuFx7Ymi8i3HwjqP9oiXk52tDqerbY
IGNcyN2a2Gqd+Du/0uGg9ETesnTKILGwfsn8gfRYAYuhn0nRVkPxGrmDbodkJn3n
Y5+iVILWsOM7M5eQZcG32BGSSdD7V3AGHWuHf1I5qWdg8VN8o5HPkWzgr6ILYys9
Sej/3kr3eQ0oA/y2NF2RbFcrIXWSo9fHZOhxx6moHySXNW9SQZraebQP68SSU3gP
jw6l3ARmugFeX9y5jHR52NSbPTSMORVoVYGIINWlMCK+5w1gXekbIe32nUXmsCgK
akyICy4ysEkt2XyNgsSZFKR+IYg+XuYdJYNQZU07oMd1i48i5sBD1CQ26FGo/m6S
`protect END_PROTECTED
