`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6fvMHS8lSkYbUZ+eH8MIJblIggbgfsKr7256DiMGd453k1/JzNi3gPPtgBopETi
dYoDeBob4Z1pJNQ2c/ndqXJqN4aq6hLDt/NJJkN5mHnMBTW3gb2+48LMM0s4RWFI
6BgGyAknEHFaay6M+7KlS1zJuBWvXthUiAXNGnGVM4zSK1rNcpEka/KnVIx+MT8Z
r7+R/jO8cp94EFshk+ySQjOxPABmJg887klbxcXH/obnaMOjotffTA3O3PCXgXfW
R5fZTrLs4bnPea9FKDB1GYNKj9C7wUW0G5H4sOoheykAa3ziXvzbiSZiLjTQkM/l
jk1Ba/f3xi/rRT1Tv2LjCJhQjnOGUsgCOPqUL5h9juSIK4HpS/HUW9ZavvL+p+xl
jv8/89Y3icgRptyDSigLSxrGg+Nj+/ogWNTmgfVJww1GH/Z9CDwDvC8KLnmebl4s
QW+Yni83+mCZrHrcw4+r4iIbiiBZls/7CxNp8wWepWAai4s309zmnUgIpDIUDvVF
mGZ5YjPcioThAZ3lljWChg==
`protect END_PROTECTED
