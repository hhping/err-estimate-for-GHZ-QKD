`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQfCjmD51WoudH4rTh85j53OIm5d8WUEqvXxLDQ5AF7QJ6s8PIl+PL2Gsf4fyzTV
uS6NswxcbYIF/GlE+2YwFvDk8iZgpMCXi0+LJZH3WSubOjgqOdCBcQQcmJ4xkHSb
K/Q0IVLaFFLA+7kRgKBw1J6o0CLO0NGYMr/Xe4rSUJJ1TEgNRu4JKcrSv54tV109
NN09xZZKmyWFme7HDXNzBQ==
`protect END_PROTECTED
