`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CoVbRzUn+XBT9lfdE07EFLxsECjJLa7DMeSnJQ85V0PPjZLIBgrPpDXIgXxQfCCt
XsjXXkV5Q7Ua35uuobqDb+VprfuvC/Yivqo71BJFXPr/X1336CXI+MxwlPHhxU1s
c5B24siBRp0MsJ5THUJgsbov71RbkdIHVGmpWxTgGfqVuroQ1O5nrmxyu677p6we
mNOHuYQ6vexmNXn7+/Ao3A1OL43XhAR1CjISrEDXPAClDgdIBKYZEBZj/4ebeuml
UuxmOREBQJ52n6+S4Xnv2FYgvZADcaHa++WXBb4JSOjCtkaw38saktdk3RiXMN3y
PC8pBBK0/BX/80eB0NFb2seYTQllO4RlDkuSZF5DegcgiFbnspkcQl7W7r9PxrTE
3nkCRf+wQtPz2/x7BaPQdtZAPUcE+dckDzK6UCPRyz0evwE2QY5cmEde4UXZFly1
6777DZlaAffIAO5xlclX0TrKg8LJgqiBd6uQJXFMo5qkVc4mmVZbI+8aPkhwM+El
Amm2qnWm+SLM9eZjb2jQzIXoGoqML0rMnem6XNaI8ZTjqPjUeka/sLWn4cHpJU4U
ja0zQLwnSYY45MbNc4zcIYcNnHnqll66WZn/EUeI8l9zVZUMMV02mEAmtKPOMq0T
5yyW7JnXSbJ71YTs53FWGWI5K69UTFBZCTiad+6A3j488/5fE50LFIHw7C55gGjL
yyrHOZXwDVjAm6uKEnrWXXrdg8CGeVq862eJSMtRr5m1xnD15vZc5qZWiRFD46Jf
8ejOAAgR++aZgUk7RLbJQOZgn9Zbxp/lC9AYuJML0GsnSrGpZP2hi2TOJZ/FOfAg
3r0OgoMujOhimL9T58t8ncG10eGzEsYfj57H6xNMQaBBoFC3OwmOZgsWVgL6pR52
mv6o9GfQUfioeWZ6DI12fU8TotvFc+ya5NVPh+huwvWRALPMcvNW76rNgEIG1xmX
R0A7c0y8KfjuJY0iLwysUxJOBmcYonfBG/4O1A6POc7igV42A+HivLbk8CxoRvVL
VbUmUjC1Xl1r5Zs8seORyIIHbg2B+yBNp6lQNruPRJsJBmQE06u6V/UuBsT4AeTr
e/Cb8b4uKjdsPFCM4wI0HCDxmWAcgaPvHqroJwkZvKkMqKsETZkw/+DcbkCVPv8r
Zi27+G51vGedQa9cbk3Pz1krHcjCyBgZx4EpwChK0Pw=
`protect END_PROTECTED
