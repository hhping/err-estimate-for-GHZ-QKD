`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wALIUWHHLrNp5KHlFxtHofKeILWh2yPYqx3r+q+uAcGTH2tuQD1bkZ7AeeNDRkpV
HxT+EGs7ISlazG0aYf9EeXWeCrHGICdcXHCcBJE8IoqOej/DhHV920HJCvpzHGS0
AEZQGfAhHKC8UBoKA8aPrp6phQ54HrvcfWvmxFez2hcYmwPcgzZDeVTno3YWbLtk
yil1RhqRcWVoa+Tcias3kd1+lLszkilTTV9Qt+DxrymwKBB2yktZWz8LmTG7aNW/
rbNO3ZXadK0S7fyz9W13O8yTOrJZKCBiHZK+keFY21UmPR5azBK96AU8Cv8d68S3
9+nw9YjQdx5xLOiHpYCgCq/UHrgorPP47k8FlJZLBg5gdN9vZgLFh15miJQRd1Xv
pTX63jWuGotXlBaIV4O6Rj4EZ32fmUNmLeA1vlT/liNC8WmQWtrSxr8kboShccyI
zdLdzZYjJlZN6rUjLpq2zFrXstIzh4qY3iQfAcVKHxSSDE6z8cEJSqBtxDgUn3Vd
IwdRMmg0XknQQQx6XotAdK2igka2rZ7iJ9gzTKNfFI0T+XeCq6ezZ/1KoryeZBfn
ebeSxN86moLP+4zFKwJ7Jf0vomM/jGKe+B2vM7UXI7Mo5ulfrFilAk0PwrbhIyR1
MQyhbkDYp5uH2D0J1Kf0jd2J98mVNlrV5U3WrpegGKZmRSaIbwdW0f1Dj0MAlXop
EBQpGq2VrKAUawafzAdwhZ6Sn8VGQjDHZj1HqxkYBG6nmyV1r49Ne9F4WuYA5XzN
tdI1zS0/BVUrmV0NUURO0j3ixC3LomncF0iUIwEavu90/y9qVUsz6/2fTDUSHZMt
NMm+vu9RYZzzxCUC9sxA4iUBA4honhaMt6zji1uooCDBoKEauN2+5+JXi5R66tqb
5sj7QadGzUrLa+yK8OA7r1Autjcm+lK52dOUYveG/RxQFmo9yDcKFoh1gEQNQ0J2
xF2oYZBKkHZwWaveL0mTLxEt3h6GLuyaKdwIwuZZU6jDu/TnnxsOED5cX7duGwUg
kb0/oBF1WkBBmjxD1mIAi01iAokii1sUpTL982t+QcgpUjuGpYU6dzK002m5USLp
vs89nmm0Atq1cZFVmQMpdKsDcG51s9T6ALaaerPIOxHoml6xUFTId7AthE+7WysV
CSI4eG8rIzd51UowEPg5hg8oMCEaDprFIR90yLBmuilqae/0SdQ0H7WEXtrZpVeX
vRidW9Z0Y1+r2uMwQATwI87hcK7lUsnCe5z0IRkok8EmvJHZdZz6f5sPK1LqxsfE
enu2aSKXAUDlm129KmT6j2Z29iR6VaSPWkGKgKb9ZSFJn6aaQguQHSLpyjMalSCM
l0tbOpyEwjlWI0qA5hFeQmEuP1ao76Tzwoqp8AcHOfdR56xNhlVm24SNRENN7Gam
/dVxrnxAambGKYfALPfOG7ULFrSdDL7+XpOKQ7bxHTHsPe1ilOOncnGPjq7vWr+v
gKLYEpLFToW6Vaxj8qvi2Nv/2s6qQuC8lwgOSzcO/aZ4gYh8miL35cl/thYCc2lt
pOsl6DsPLPJlTIK/8QGOfROBFudxpI/9n8le54VNdr4=
`protect END_PROTECTED
