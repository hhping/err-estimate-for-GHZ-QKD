`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GX6fiPlKc8TuNuxZx8x0iNu5xdIw9NHLHEbgJOQzjXTvBsb1dxGh4feXvnVkRGyI
BoNxx5fNiyXUk2KDFRlajaTKWGxuDLVqX8C1jrr2bnPqKQL3ppszl45SEpiOOwXk
+ttQMlcBGKihZ1GidQemULH9Ktvz/rj2rL7mgBbPHCa8whtBWwjxR3qRIcrAgGbQ
0KUaYKRWjsk+yChKbXC0dI4wGksodEKQBZ3qioYNandnajXh3pOIHU2p3oBsIA2L
Z/6UqqDBWzvUJLRN2KeVGy+FWONk10hibKWAQMy/KSHASDxBydvCxOduV0HZ4n+W
GzRrL3IcvCx71vJ2H1JFhtY/nTtk0SbxrQKUfW1xR3S6iwPvAwidFhEggF/AmVBl
30T/dFowKlHQEMZEVkOvE2QDmWfxzhrP0+cp1b90IzINVOPQud/BtRb1/FQNdRA/
ttqBAcFL7EGKBBiRTiIkFQf6s2cvXZomYRci084xrwWFozcCH0tqC+ngmv5Q6qaM
D9Y6UiR+mJsc0/HYz7mqmuggDcLJFUyrqp/RVxJLBWNR3ar7mPKJCEE5H4Eb6JKm
3nHf2S0BHVUict/DLqXJ/uo0bBFEwPt7hRFHsA5R5R3OuwTLxeZNdUFpssclbZhE
3+M72DagOrl3QNlIQUf+hG1cM5xxOOnvs0T47WTjK6x/nTmllYHGxn8Iw73njQUU
sXODwmsZAiZL5aZidYrOpgpnIXt2x4eV1Mqsje0782FMa2V24+hPLZ2AiY+Loc+B
X7GyQ5c5ZaQ9FpfLX5sHXbXPWaRvhkJ7C9PzaOkhF2ZPyulJF6iAo+u3u70YVibT
KTMbDj+EpRR2ta5LinFzSaVb3FAD72+rwviVyLAB/pyd/nw0Z7GTCIF/fCHrke+H
G3eMZ4dUU/uN14vw24yDbct1BXWh91SvazDXvj8LuNr3xOQDJnkxuaG3uwoQUoUe
FCa0juD8TxJ4cJ6U2IAsyaIEmoVRs5vCNIgHDCZSEP9yNjimizsiMII1Mjj2Jv0C
ByaNJ191Ih/h7fEkfFGqAy6XAr92yGgmlUjCKLJFA/ronCF+nmqyinXpioeSdnC5
SuANMvzoA9IskqhMyRYQ3k0ye2Sor/OTjzvKmbWa8A9JjnJdl/6MiDUhudHA2Yp2
a7oI0U+tzuN71yPOiG1KPHwspF9Vfnq28OYySujAQBbgXQDPrASHboM+YtDQBRa9
KXDJhfohFugqWlIVqYL6vzP1rTpZhHDIlfdE8HvCyOsCMSrUq7ZD39vkJVrVpjdi
78Jo/y/RISWCX2ATwk2koeHv87Bnm7yIYMQ3SrtHoDuaS7nfJdAicuoPSKO3/nfv
myt3K6n2hiuguL+EIscH7tqPr5Gkqxd2vgvAOd4iPlybY6i+XpRhyt9qB89Uhp7D
PlgosI6MPLj272CV6CV7lw5t7H/i4MpMCvOc1vu9pGz72ESVXGHzqYTbkvRN8/19
ncpP116j8RR4YEbwmD2Wnt3yxqJeG4Vvk8wKbmSJ+sgsSy2M0bgyzBYtcAebT3Ln
rBXBomHwT3zMKytVqcyu0VAsKB6iiwl429uTwQx+DeUX1yuxqbz1owisLNvSGQG7
I/Kc2nwcTHnVzVqZLn9KyLXcAXlq/1ld+h3eKkaHfMFaOulVaUjsCuT1EjH2Zp3v
KPCtlZAmOxkfNdVBKK92pOXCVb6MycXeI0jYlMZMuOflIBQYoZh73bQLAKocfaWY
`protect END_PROTECTED
