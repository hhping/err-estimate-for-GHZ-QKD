`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xROUBiF6IMKDK/IM58VdmbXMwJUzrD11p7J6II5Q+sxH7DjlkaVg4a5KNIikKCPR
FeutLsyLtLhHi2Yt1MXMdJq1g4AaLNL4w4M4DGKsVMiUIoZ+IXklX+bi/bhou7gJ
64UxuPMyrA/lofi6NJUPoL4MoYjjSUoksuJmOE6cJa/XhNqVsKO6IXfd8rStKPKZ
8WFLcVdhaHNQEdk3I+ak0LSibNWC1cMdyIxjuDB1i1TdaIO2PNwIZ9PmmxgDowP8
CwwkrrxFfLrDwUnC+7bcEORoda6QjkoZHgSUmp66v3fOnziFdgLln3wnNTvZs+B+
MYiTVdUsjWpPTw/yBPtauq9cw/aQJs0kx/8A+d44r3Erd/VaBsX9GzYXb2WqALzJ
T3mHLLsdm862rSHCPXXue4CJS/EIUNw08fhUh4iUw8Ra4ou8gtcSIXu3mFLEfurO
jrVoBkbUuhChruv3Aa5LqnONEEAii4jwpWS8AJk6QVXHSxLtWYrv3MR4SUD7h/VY
67tZb2X6lO8XcTTfW7qZmEUAgcCjuxUf9oYeuk1rB1c5XJkuMO16ZtTUnZFgag/y
hhYPd0/KnT62jEhtvK01UAjygMGbnKd3xQJSpYDZxmRavHHqKCd7O5qbiQdL57JJ
z0hAgrrv1vMpuo/k35dEApEtZTB0BSbdGLhUHJ04jMRJDIVqZkP98WGWW5oMcF+K
cFDqL9qXG4iVkMWFfUsQDJB3TnMAyTD6OXfFoD8xPmdak69nf+foAw+5ffM5ubea
tO0abzkjYcZFAyAfNmprsrOe4AbN98KBvOddh6RimOc=
`protect END_PROTECTED
