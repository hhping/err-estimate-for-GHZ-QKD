`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7Gl47yXFueCBZjr0H6bEr/YY5ZcOdVI3wlDGrTaaPJtaFJ7vKwgbDeXO6sBEZ/v
mWfdi17EU85wFOWQixkfjtEDnfa84AyGFIfSz9a1g0Xoi8G7A0rYjEsO0emTZtxK
nlHt9duKFGeRl0OrgW4D8MbIw73yUnXYdhH/sVFBdbILD1EL1dU+EZoKvn1gtItd
HR9aZU9q5Omg22ZTupyFFcvErHtEGLlXIZsXJ/EQb84xKXvv8lsrIfxARi82hBaG
Q4jMKS9fXuCIcUcz9Vsau312jBy9MITnKgSVS0A/9qSahbWdIh0q7CLF3Qj3GRLW
ViEe7114zGa9HCTLRfK+Fkl3SttNqUs/jhX66FE8LQTZ3aihkrasdKOdEVDxLhMb
xOxq2WX0CNrcdh6r8WxVl4Fcf0pPU/4EyBJ34TaawBpBpIKqZVmks0c00ZUWw2tm
mA0Z5beUvBpgX3VlJStqsU+i+WbviHyTIMnLatc/xy1YZjzZIlNNmpyQEDzeatw5
Kua+0LNfD9gyh04Kap4aE8wu/eu1DFoTDQ9m0uH52h11qAFa6hKIaLhQVvh6XUaY
8uBZR2/e7vrjIB7MFsaJaMBpDleplcrMhIOW8USk5HLiw8Pnx631HCRmue0bOwgJ
Yjvxa3OUQ5zslIrsBY7WdBimPxTzGPRTOgSM8y/tDeL/DlJL4uBSnNjX/vnUa3rw
mJ/OcrVNGVaqc7fe5myWMB9FkZRg3q+W2UT4RftX31tYETeIOB7Tl6QsPWRCsWer
66CNWyiOkJIHppuT8pSrwA==
`protect END_PROTECTED
