`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aa5v5iLr6IW4S0f7xfspM3ePMOWZDdmRl90Ljgvjp2Ai/tJqoD+P98vx7DSIb58q
ntUE8f2T7BUQafWeDUtrMxP2hedY1G7ItMgydbHrnksb/If9B8AfCiMn+7Y2SY7Z
dzKzklWhmXlmwvqHODr/NFAJ4zVN4uH+X4ZlWtKPFmoDRLvI8ZDrPWGuggTqjJrc
VwkqjS0WI1L+OGPW2xB913Isp2lFs5rIyOkBWtAMsTpbQAKTUQhb3HokPWT0gdXM
3nrLWDBU5eDczrvTf7apEKJxhipM6a41xOphXrWJb2GRJQEbXMDWXWiqBcjIZ0V+
GTaaZCfjd0SkCdZTebWNRm7QeSGyhOFpgs8347GYa9a++xK6Y9DGl/3aXv6/KxUm
VvdmRA0k2kou8V/x6aQy2IoVMBNs58KJoiKgPbAG2eCIhCClU+v6SQyurR6PB1Ou
gWLE7CDw1Hvge+iqnq9JHA==
`protect END_PROTECTED
