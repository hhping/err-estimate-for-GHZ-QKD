`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xwLLThUCD7HNpY80H4dRJtK/ka9fj/zoBEXDYqg3t63nRMfVfuoFp8Gu8L6UBtx
1zLKfdZEN9cbV4vOJOEN6MzEAKlRCzqiy02G7yNorgrkHx3cHpmZkNv7IUIYQS1r
KlCuz5vJ8RqQRWtFYdYi8/5/1OTkHZUAD3YmHHQAx2cw2zZRRDkxfyGiHzDqVm/F
SNH71R0agFl1VSz+bfLNdZa1bw52UyHCaoTcV8FRsLBDUCbmgsLQZBXVeoFeK7TW
+5gyQualMRYsv7GyyzckaTQnhNqmo9tweZyXzUMPuagdwLFxIwmnNdUvwFwKAc6w
8kIKa7Q3v9hAvoYQ9BdcoB204r2uqrAE5g5rj2VawmhkeCU5iquA3I4UXLvKBpja
kesY/tJhgL4JwyFQNhkshEOUrY2y3LV1CFE+wx9lHcgCQqVqDGYvtp40xR2OCOQC
wB3Z2BHfjo1rysAv2Ku1VeJ0tyPa1Iz/97jkhWcNwiVawHIDMo44y4oddwvw6SYT
Si4fzNkveC9D/gSIovtt+2HWpBUeU96fuvpc2IyL1z1htbRvNItiuc0Kb0GauptF
FajpAv6QmD+afMHdewHuDM55svNDku1Iv4vkfuAG3JJnJYA26Ck3zHaovMbktoCP
kv5uN4gBsuS4LgKkgY/FB6xf9ewnLORhb8XN07vKHUQMm6XV7esH6usmlkQYKGXN
oPDchV5ds+9ifWIf65UhD6qmtSOPCtK5h7vIZ2wlKIxUhyF+KfjfKXa8hu1OV4ne
Z7Rs+noVdri3RCdGabe1pfWt58oIHI4+nXuvW7o90w3iUnYX6ATWs//DYP92vYwa
C4vwW1p9vQJO5th6JQtOGVChbWfDmWXAmiozDmbDy/ciBUeeL9SXnCYD+89XBPNt
Hg9nwqWZsR4o5rCuRxWl9QQuqTg137kJUUUZCHadEfP5p6pgPW1dDiQWd3BtSe5g
+PvNbjI0k7PliaoBo5FceE8sFSR3HMnBe48aNTfzSX7LNKaX88Bclmgkk0vciFmR
x978TRU6zVJg0G6EeuLm4N9gCQgVpQ4POsOgrrcBObuYZ1a5qKQcGlM0lEqQ6aGy
vup0EZLXXor0w0fPg6GlmVklkwnEHYNPO3a7uD7iRpzNtNeqlLV/PAt1XsfnZ0ws
O6yBf03ZGo1gMsJ3SesP57Nuj0gNBfadOHiIYgJc1jQMFATa9bf8Z93nhLQVeoDE
Zoym//yBpdoc2QZQSltgcLgFapYdcXIhKFCZTtfL50hrYYbAyV9vnFbrM0GbwKkA
JSWMy4/R6IFozSrpvnrh1mwgTR/Lw6wg4QpXuLLGZSu+UIRoiB6BpfMGUYwKLYh3
UrD+qcqKE3p0tQRIe4APKW6FiJXNCWGetexxJ9JnVC//IQlqZhcVhNCIgBIAbb+u
Cfj7/ysQFTU+IrbRGZIkGHmP8/o3yMcOIvVbI0ClR5yxcZcu/voswiEZ3CqSNI1C
AiNhnG5iuXfSqYIlWxDf+LB9449m0T1X74IlCVfW/eBJv/p0Px8NoR1i9Bw97JUz
dtjvfxcdLNsPczLADBNaEKtPzu7FjJGPcr1DxwSbOT3bBrwXgNunNTxittW61Ddq
+uz6+txSzm+LbteNzmX7yf+kN1QScFG9rtgEHupTs4DMlWemYmTx8/J8v0dIJvtE
qZsA8NBVVdmZbqhBg6E16Xphy4SPfZElrO8R/5Tt0c7jmfbXuUw/7NWW/wMhl2LE
+IzwaoFabJ9tjF8D0KvvcpwDrVGbhEKPWOWBdyPla2xbqU9UdCN8K4QLoaCBp7ib
7tP/zbFde7/jZf0Xjjq4z88Lhh3pMHevLYCHGVlATFxqk7UQrirtSSOy52KjqlDl
TQP4qLuBeYodd4lkz5QDu6NH+qG6fVVwzFOWqvmPtF+jUWt2ALquOhFSRt53ajgl
H8/F1Dt8WUoZ81lyjuwxYChIk/GhJQwVbyuXrHn5Ua2BejEg9Bic5XE6HX8eCNoF
Nz059X7SBksFNyEp/lVaBdrSsPFfjtAQ37o3DhhWD+fY4UGdoyhEtVZ1BAZgge5/
LKLscrpVjZiAkONV5qmcedHpOBmf0ADZGqDLMDUeearZ5MpKvuyYGin8dVes1ETo
jwSm7gPOSBu15ezcKRRDKgInYOskJLup1VE/5XQlJ35LhCZ/cFmRn0GlY3Jac+QD
+Qu5mMTMs9nB+jDZmD5OcZdsaQ6nSAioA8Q1gokEJBk22LXERpFCUFfymPQIfH5E
mPJgGz1OAZUq+rx00h41zzbnIMjhrkBPVIbh7D8/P5Qr3SwxnAiRaNhKkQaN/zxL
hEfopAbY7VrZrQ2TLhDlN7ia5ChjfgW+N5K4H7FaJ59ktnKM24xQsosB35Ram3XU
atL9oHjxm+77NSKH+5bExoZ9sOVd2ZTWgDUL4Ulvs4uSYacT1hWUpEv/4A98REzM
Jrfk9CiItxL8U/1hoCj9SyqD0j1nQg1oMKTunB1l4UFxX3sjFHUwgQkto92h/VS8
UZwj2c0UO5Qteqx1SIXmZj4YxE50VVVpwiswXLK3ZTz9o8bxa+runxX+/VdeeBF1
SsQimxxH5PEJGb1miLDi/zcH02cgWrNnSHz7wxxbtZ6ZVNHT2mqQA8mm5idaol/2
su0Ncja5zfZvf6sui+21J87EmeNH9xwAXSBU1z/2Vy4Fufr7ee6prtLrzq5mdEDo
jzqy+hmWsrpL91ZmLyblolBiQ8J32lZJd/RlxkcnpqTIBioPGIlnQx9n1jxRed/J
SUt4tL7hdnvvuBygLcYdCDklQtHhV3DgMl4FpOHOq4ErR20+8KkUx0qky+QgmzJN
rmdMNDpIpVDElwT2NR7Pm3Bx+riuyY0SUz1niixKFdKw/yubNQGz5jgJPjTDa72n
TtJJBGzVZrws1t9jbI162vxW+BcHg1AdsScwwDFGDaEYeXEAc6u8vMEuoj23O68F
IsQ+AWCCzZ321ZRRS7BLLDbC0cOwOpC1SkomE9oLii5OkFDYKq9j9SkarimOUkWM
qvCsqgKoZidW5WIyLVfuFBb1srUeZRUxpX1MMGVxf1Zp6tyh+2OoKqM959qygOdv
wLUu0h8atrdUJCY73T1N6OyYQwUfXVRa3yp5miZeN+JExqKSzZ4SkDdiO/Cnrhoq
fnpybdbGNxL2Q4Ih4nhcMduuyj21kFvWFBLX65eNNqrQ1wHyq/ZuJXokmRSFlmTO
t9S/E7aPPfEIL6w5XBdDSxiGvxRV0c1LAT0h16I/KyUrkN8Tie74IwFYbWMRx64p
ek7uQpJwNCJIZq24wubXpsHibkH6+oUGEckaIfiT8FlAt6paUFD/x74x0+1MdLJW
aLcIc8QRDvYZSD2buJHUEtfNdJuKU1/EXFhV+d6anwRg05fX72FMGSr5DQlfOwAX
sg7X9XkLXuklsXahDISGtCUms6v8WMkMPmirKnCgrnOAjYeS4d53AbrXNRuzEJR+
azFyAwQeq1w5DopyqYhaKXMSNl8t7SWC+54Ps6AYGlzn5nOvubzs12KKHTYXegtT
BK4xCAH3vlYFcZQ0OTMaKVoyRpOlds6jefC8tpptrdC6X5Tg0qmh6FkD2wVneJGz
+Mbubngd0xqtE3LJlhjyfLmsUEwySPFrb8N9ulcXQ3Z5gGqHF7tLujiu/l4/sb/D
Vv8fBw2RRTAMvo3Itu0/x/lLBdU5PPIFn0iFAQfMQWWPtHZn+ZmW6MzbSU3738FU
H04pB4IDWRYaLc79eek9zhMKeNCdRYLhced9kproBivkWci14HFnYh46qxhTytfI
YvbjvL5HBOtZCl/n7Au8hnfWxNucNquWHVydVorNCtQKmBZFjmp8JrpBlRQK0Ur1
3vLuTDu86YyCcV7gmTOC4DsJTD2sMXLhN9773wK1b+rXfkqdLQ2XMaPT0Jht2JTE
iOQTRxDaPYInZRS9ajLRHcZqqJdEt1zeRZNDG6R9f6rEaaUe2fKZiJfWObmub7Ma
DUnGfoepRJkv8QkZ8mx0I5ad0FzXajIOhLOOPgYBd9IBIDjDRbI6eX8WQ1HqqAjH
Ywn3KI4lrWE9L0IOtyv3VmHPeMp8guXQTbvQVqlKSakpTJ98D398bqc+0yPf25iz
CT57O0LeOPlhWhnxec/0FKyQEwfvzqbaK3NYXufoicx9sKMgfpVZ2plfOcuj/Vxw
DkMHk18D712RJRs+80NUYWXDvo+yZ6Pf5wYm7U0zqAx6r9qDu02ojFw6jyZ+/o6c
ulDvjEewUbj18BeEexoMw/jew1DAmvajmHuzpXYOij9rwQzTUuDRNQX7ox67yMfi
6FHwHlUSpzmyeMHlqICnDzyE2a3dmG6L+7HTqsOufAg6RORPMNuY0/NQKKVo4s+Y
drPWMdtU79ARu9RNL2PZw1uedCDqCMIQJN4gvH7ezIzvU8pUOMLTpiEPdxc75ipg
VdHsNVvZ1TujEj/38SgU1yVGiGOwqmeyO827fNPHrfO2WAhKBQSLSZGq4zK4+LTD
I6XZDoCz/tssWvWeUV9Lb2xpfqYCVbmg+tsLBq0X1SK1IEFPK8UqcjTCZOsytAjE
Xsy90eb8o3DiYh20AgmSLuzan48cS8hhawGWbrgjUH0yMi1twYD2LJ0Tstlhal1r
JdcKO/Jc1gA350/xuRdEQQqfqhJeAyHqB9stYv863msySacqBRK3FDN5A0unUlvq
/Ky+eQK06j/0uYQnZkamDBVVNmHxL7x+j49GiwbFgJaSv4VbdtYuXG25YsGMlQVq
wc6nLRMDnBxd1WUVdL7pez0pareOaUN7WMYvMfraIw/7F7aWrelCY58T6t5jGp8J
PMT8Wi4oP+UR0h+AR5hTsvZG/cS/AutRN9knO7PBdgPyPoKLZ2ef8xKwOe0wDf8m
hgNeC6/fdA1zbHUtlu3/h71qj74glz3N4z0tlATGuLHY2T5YTtR1TrrR2asR3nIz
fINwTtMzFq5wLY7FcrThkKUqxilbzKS5CgPGvqVd7LgKDdZEkOAeATV3gtb8DMqm
UlRpAaNqEKBk8M2Ce96Stp2YEHZyDV501GOEi5EbrU7XWi3EQulDkMqrJqOIK6x6
HK4eBt+W0xOngM9iwO651oIYfUVnUPNbTe/i9JkM7TI9PqCLMtbXeoOyECqtXJT/
+KATqcsYuZy3yZdoZUYQ7A+zWKhOt2Cm9T/mw/JZQ+3retEFdi8fHWym12Up0BNB
39Tf5soJzldIdy3iIvIa/TBkOLS3VBEWfKFLXDJb0687zlCeoWtP5dn+mktzXzkn
G18fuJPV/tlVaN1ASdiWddLb4jHtEjGQIg/FWH2rYM6ac231IQ/ENvypCbxMKvFI
qB2ahHJkRggRm2Z5wy5UgCuiM/JJ7jRbuI+3gmzldqftrA/w+StkaMFvthH722jh
zt2L/ksnu1hC1X+1rOV2p8XZhgPwIAQnWUev4t2PMIFSZ2lyrb/+NuYWF0Gu9kQB
fwT0bwvUQHVlytv1OogumwAMfsHlCK8jxE/z7QiFvEIfs+o+M9WNXN1M8u6MMpm9
cFIYeAqDLW75Epy0AK1qqCackKCQGwlfbLe7Mln4aTXAxl92NtGGVnMec2kRkcT6
MKGpnMKtC+c8kIfV8F91PvIqiA2EVc+mHI0jUk4NzTg2eYbuolVqX6ZNM8ZTa7w/
OoPfWz05oj837TP076ZPamQsm9npW49SeIsONZ/MDKpzX10pI4TDZTf0QqdQ+5V7
DVUwQ8Vam/m+f/qHLhdLwzw2bL2O6rUDHmsGDzOG48EYlz4d/1R4uq53ebQuz2c1
txji0Yg4cDI8Bh/vtOM8yy1KXGxKSETEH8QIJOZplrADIk+h0nFBreZPyZOugHN3
InXtcZbKLdQubywC3bn3mX3QdXq7U7wXRVAZ/pVpTOOhs0lCKNeqYF7WKnvrRhWC
d740W52n/l/4J5vpDOI/tU8qOYOyc05Y3qcwOevlSYyTNxTIXrs3DyAYVD/1lXgG
KBZ1FpsYCaVmWbVzlgrVTf4V8VN3O74VycFG3zY3UW/KexHDSxaA6ajKMusCsl/4
p6/Zunz7LMdGsG4ApNrFMmVrLOugmOX6qfvjh1vgfSl55rou9fwhmVWQ4ZIOWid7
gtBSWPgMIBVYN7SXKFo9XLIADi6gsxclaa3TTPz93OaWMhFpLmHVC8OAFsWGdBAm
1O7CT4jPSLkfCG810h2hXJaTCvYdBVPYfkMpD6fdbG6DYthycFiR2VzUKcp4X2Qm
qlnHT32LVWrB5eLOZxG+xJNvXULCflxqJRc92yz2gjSICck1Lyfpa0ThcVv6qSQM
xOQEuUP8zvGTgTivIsMfFpSTotRXitzJ00J7XHFXyVermEe0ltrqec0TWWlGTVKl
gtHKtdRbUWfo20yCYj7Zzitv97EWgpQqZz8Mbz/zbGcqdeXs1jMWT2WuG3DVXNl6
3LiPB9pW9bVDAj/VV53XhVUp+Rkl3Xh87MqUhVWyCQwfpkNKzm7ik5k4yuOeSZCb
Wv9QgcXfaVvGEuBr03x3WGOsArj3z/GNOS5Kp8+ytWxvRioqwihvhN45bioey2WB
lRkB3a2jxDmvF+Y2ePEyVkk4umXfadXNHIgaT62/B6wQ1gQr912k7I0V4Sj+V6QP
JKGny1PUcD1++7xomulCeS+F3wTxGhxxsZA9wniS6GMwW6DOkV5Fo//TeOS1WnCr
68oDE2vu6okNxgwPfDg70/e73bDlDAYxy3sXeUDWjYHxByFeGpVYryqpmkb8Sy29
6PruUX1j7qymWg5z2+LLnwG9dUZglu5rwxiAGDA8dF2YwgJpFcouG/H/qJg0+Cx/
jki3v0zaWtolssl7O1HW1Ky8GosUgJIWfSLl/pTAMIU5ilQAuxYlkSoOEfEqzFBx
1apBXxITMVR4dmfijXzR2E+GEp2dKEu2bnWyWCN2ZkP6e9GrbpTfab89O4ZQ1P3I
Yudtwpt91ZSvk7I0Dz+fHDmXhVwV0PglO7qtpgJJdKuREphPk60colP1Zb+D2Eoy
mZQwUzW05AUDddszdUJgGqiptqv6jRunfypVw2ojh4Ic1eHty0blp8nju6thQScG
2KGL7THMHbIJGP6DeqyH4uisMqLXLur8hJGZQEZGdaEVr5MYP9uavDlyEMjMCeu0
geBrHRT/FT0VrcT94qeeZ+n/7uD9jVBypbvW2gW8W2dbCa/LAtpMN1/77utgEBhJ
66YbUcHsIllCzCTq8Yy77UZ/QYbksq86rYawteLsBJSzw8xktj8yoHNZYHRClr+1
t4TuUYnGirLdaPbO5yUwHnZ4kUThbNpaAvd6dwmeyKrijc5JtbblFzx1gW9dKbnM
2I0Fd35qVC5U+dJXu5o3gZAJe3Q6Uixq726h4iJ/Sh2BHa2r8XYFZL3ttZWmdune
JewnF4zCtTqJvFFXWB6gayxSe9+GFOuspIBy5qkpNHkZ7N7FzRaoK3PTvkKXV+aj
nLtOvG+GLCReageUywfi9wESj27LhA4+CvRPLQLVGzif72Ubtl6OnAhJjRPDHpXS
ZtbGdipvOeDRLErgqrlFMXAioBxjCU53KLZNmPjJYqkqbecJse1cMp6xHOL44wIw
1m5pNcHNjd9ertjoPOx41ZXzXjXn+DkSX/DHYNUkznhTHh1KcmlQHdW0eMOhnlrh
d3aUt3HHx/V32+9QF2xI9GoXTsv8yS2gTWAo66xqbA2D/nPLZwuyah1wp4ap6xjW
0vocqMKusL5wrJiHqo2t5WgDAzrDB4VtMZPa/ANnqvEBt6eoqvJxw6dmwnaF0SGG
wxzJ5OMxOnC5m9+3c56SaUDgxjNmDvKbZI9op9BHiFSK5rUeehDe+MnMMpzEOX19
eE9Zztcz1zTqXU6iH/QJszC1eWeO6LTKkOmbSJBJGjnfaAJ1J1eN/tYAc9Ue/2d7
nPfD87/HUSWUUrz0rOsKTj9j1/ZmU5KJmRidEhzChIAdoGy7qRaS/9mh+JCO6j+q
EUpA4s6AL+EVgMf9C8ZzWktTsh5gelHFERT7gmh2YmgKn2c89BrwSAWIszt4anxf
7w/R/p03boQ95EpcxPzOdv6EoYE0Rb27G+RoRcqbxVbTTLjPhB+ErXNcikA8Zd/9
oWBiAXu3+9GbsqPV6Sl/TzTMO96EevSlFr3LCFd6tYsL7ovwyKnPCavYZskG9Kzk
MIR1VGvwzkM1UqE6DqBuKAlfgihLOfCgvrzrcm13GeTWk7PpEaHCOaSgXlMeC1nf
xGTs/wJH5c9OMY52MsSlcIzdFw9msXslQyH1irsSyXE5PjiMQJFBEbgvjAug9rRB
M3gjEDq6gZa2JUPw7W+z02G2/LK4szW4gSPaZwAlucdqEvk6Fqvw2e62Ut7KvORB
ZxmtpuwWi+G55a4TZZ1eIOYREM3AA0XCCbCWuzP5vUIf/m541+TC8Sb7VJqUTOTI
D1NsU/Qhoq89RqDgpkY7HFAIBbbbdBNvuuBh2zIkfnG4+pxKBVHndN6i2CmFYGaD
5/n++a43RAHCC2reMyFxv/xROI/1UOMUWc1Z4TWjhV443nTNdeu9JU9TJ1AlSlEX
FQeO9nhPXbpv/ZShE4tYnggeXJbR1Au0b1Nk5hg9tI8qLLwZPgWLWcQBNi5XAPRx
yPytwmSd9zGSSPmMj27ytArhuz5Q63kL5ugwrMikoca9maEYZ0zeU7AUhRzeTo9c
y80bMHtFYnh9VwGYGeU2xUWwbD/3eVBtAzDTt+JnCo31i7DAyM4vvJ9tc+y+8N0d
8vpRGEWFRISZ4ZCLqeE4n8zUQY/fT4rPk33QoVxO38AYsHZEhkNB9RTDw8nZlSP6
EDY4WW8Wr0qlCC9ehDH4F8VaMijJFdIInARTVEQpp1Hd71J6yCd59elokTpUPhNz
icP6qyM1/78suoePqoaWcy/CYF8sSZZ7KOqIXYc9FlsE2J4NdRmhwj/thG+5fqya
1wu6DW5BhY6IoCkeKXaGGgnX7I8EP9hvmDQcWM5lbNX45DT4lSCXuCJkmXHHId6S
bUXG41AL5djkbf36dBCvUdgnUGYDVNh3JpXFDTwH/6y7YxJnOSX9eQPsIpHZpak9
IOgI6S5AXSY/VAAp2wQ66x0sYqJqLAT+CZZJiezb1SDIRXAo7/DtNRRYIv3/okFc
dL6x8nWt9cNuXO03wkP0FPS4gkQ9a2aK0Z86izJspIsx3YlgxhBsAcVBXVnVMgql
SY0ey4VLVrM4EvXgMdawkK5aS97YKJsWE8rTV7V8KC8y93ozkvnmuuJIqP0TM+ZK
dItE5Wwz3v4yedK/BiHz+QWnaFeLBoFsGONwip6KuxxSFM7cYE/yTlkoQ3oZ9fUL
fcOaiZW4fB3l/M+2qZq2m80byWGojssRv5Siz5pjHNjQG3VPJrTK9pg0x2ge+vv5
oBQCU1/bQ+g2RYFm4ZX7/SwXNvzaMfCskhqsQSRXY7aCf2DyQg6N0+oMm3WcXeQm
m2aSQr6PBMnFf4WcSYJyYPXqdo5vdiTij61Yl9SL98978zCNs/evoo5g5d1U8UZV
RyDsUKgqAVCpPZZvJW4nxKtQy4FOVVmnirPYcG/BW6SAtFch6L3tUbCkl80+rfIB
pwqAr0SDm8xN3DbhPA9B/CZs1O2Ul/AXDml0tUkx4xhxTmUv32aOiFMCiZoeGTe+
Jplnr47OCu8vN7M2ZJZa/vChlQ3p2u07lwZcxvSCZr/jG6YMOVU5i4ZddQEuge6e
mzcvkAj6+52hRXakNF0oB/v+JH8DLJX1sKRD5MVhk02wPHgKTeO8sZ/wV6Ol+B/W
XaGedmNFHbeGsIa86eojWdWi6Wq99ay3mFfryjRKf+vYVM82JExveLDKGFEhqt6s
PI63qoiu3pQQbcHqfLxMfI4lkDe4r1eyjLqBilzKUl2TbO/bBDAXcvHMi197PUso
Ic8QAub/iv7CCi0wCba+wZCnfDLenyRihXy/qodbmvu1+FYOr36/RDl/iQ65T4wJ
7GNCdh8GP7QmbuP97ZsGjz6JkTbum4ZqtZ+461YFNMS5aAOrEEa42GEgG25VjVVB
AuGN6vjKw+stCEYuMK5DaKx2F6vcuMEBhAeodR4SxxQO1xo9w1VhKGEs6e8KffIy
g0qDUvnJnDG+WXbd7PTaCoVbSFAs0HNmRSLnXKMa8zKKpukA2dQGMPT9CpDzgKIg
HQFeKwGNtM/39EVaNn40q1RrGLwCgWsqS8jWg3ajPG+xbOLITgsM18qyCpv8kU9w
8/RK+WAjPngR69CoiXvAD3SDR5iBjtGnb1JLzR1YiQWG7EzC8tXVjZmAgqJYaHEu
fBqegkvSjFJOSX78dx5DvattRY/9g61Q4V15eXEObQ8fG0VOu+PArHBpY+E9PnMb
wrTgoByELUTvHq3vJ3kTsH4yvVYWz+v/ckpQjX3oVbpwz2d8tudU8TVOAuutTzrn
ooB1Ohu3oKOH0ttG1/cG/yTdZQeOgwdHm0euaYK2hnIeOVldXBxMGxV7IjSa1yHm
RPZMscvKeTFCc0Eq+983NrLwhkU13dEXLv1yoS6not6AqgibyvGOdYiIUKWFs3EN
0/Cae5qsW5UQkiszFK+vLoDZri79PoRsTqq93RtoD3wlyQDgV8ZkeIOV09jLvtzH
Ov+zSuXArNTun5iHDtdK4U/sMO7dtCbu4UN4+5m7Ut0jLsakAw7wvlnkmB6SSMhe
c2gxmS0yz3Unt6nLa6QqZRfKiu9wK1uDhb7UlW1Utl5zSV04/X6zMHAeNBFs3o/L
niURjuBR4GnVEO1Ihock9M5sgtZ1/fA2FQ/Cuamkeidb4iU+WdTobVnjk87Rm9Rx
Sh6KEji6au6+1zAHlYsF1bv/bXIlMAiAXpQ3LCkYCe4np39j2lTZ+sTW10E9rCgL
nOgY5IxSbEfhaNP+AD7xZIJ8n1f/aaLSwJzn5KYgspGUD6ndB1iFHMSfmGPDzYEy
f1B0N3GMy9+LHLOztP2kfBf+E1QWoeFnCNSDU5Llic+b1MIPX4qL9MI241jUmSXa
Z4NimSjDR7T4b/35PQsAtQR3ln/D1HiN6tqJhX0V73IeMK9xHjoxtobJMy6LKKPP
VEPnUDH3JGMxKoAtsyVi9y3xtt54aB5Katr/8DCrHJvsea8HZ8YvNxNOhzlel2+3
etn3tVfGzA5TyycutEYkPGSGF8x3OI2s10B1k8utdALHRGhrQ586ED7PbbfiVR6u
Rx4I5LS+3tmrBjIuiDd7k35ohV2g1DJf+PrtSJlmlseEy/Zrqax10ctOfd82csCa
oFP6kfOXDYq3ISY8dRlQlKxVayDl9lV1D5NqxLwitk/gTq/YFfwgmqxvm0Z5n8UY
edi/dQYPyEbwBK2mvVDqmMd3TKrAofFrCSzrV0IltkaKcJ5ku2dQJXGFULcw9TOW
c6h3GriDGNZsDEyTQZ8gqap62MGcGb8TfRDf0x4/jt5up7HB+658/Oyo9NwbGLLG
4aLvAZCbCv2NTvMJlKZ86Mn8AMhniDpMBnYpfNwL/mWPM+K1C3DleUFlHN7Z4eVL
iz0PTaANrUQml8gFRshYLlbuaSQ87sJ/s8lYgtQfeOx8JTzt3zLy17C4lIGxIo0L
+plrGc5HmSrbJRJKSsjK5ujvwWe+YlZFGULCv9ja2pECLk0pU4v9KkvE+gekRCk6
oyL292AM/3MIPyz+1ZWZgdam0FQc2IFmcl51YOGzasjYtsEXosHEg85Rh8RO7KZk
TTAmzddZBuYbGIdmI3wbHG5nNH6fG2P0ZH3MxgJZEQuR5vyT4DhYFfvkIlxYkovC
RS3MvZCmjzzSW5YGrcdZ+9tJZI01/MGxSBaMQbbcjNrBBPxk02hJMWh39xZ1TrWC
/jJ//ua+uX1CPJnT5bV6K2IzDo9yK4w3gyNwb9afp6IKbyfpNpumOUmFWGDUj4zw
laMOjrcJRboJxwq/N1cJ+wErRj0O3gGm2JgQ4g5eARtVNdmEfqCH+ZqEByiaMBKG
0+85BHWoKI9Gr8DwbkUF1v4KC+tkhejpk2ado5q60D3F/GhrJ/JWWgnRp32smFq5
POI1KWDmXsUAJAaYkCR5yf9/UpVt2azfnYn92FoNB1hDoPig6guti8uV9/EK7GuJ
aBnzqyb349WDY3NL5JsbQuA3PhcXoXUbu1ee6zXaJno6fWKHHVLJc0klhtquSuCL
ZTMMhrBxYneW4ZCk8uTuZL7Answ1Iobtbv3brbO0bb/5y7LvzOvDruRZngJzosXM
DRwnxC1OPu+DZ7KQ2MivXqEMMpg95aPbP2LMYR/aR0AL5JLTS3tdfR3DmganAsrw
BlMFPijmJvjPyGL3tCmqd+IkvQgyVIpsRFMatMGs+db4/r5cHO3vT85Nc1GkDP0D
y/i8qApPHPyfUQFAuVjVOoVEn2ZEsHhwSbz/yO4mCKcYs0H5qHgPZ0CUtr48qLnS
8y6AX6iMMJUrlsPp351C2PgINWXFItiL+yF1ic6JR9T+gqAFeWVHjew1upfVl3rU
5nRDp97Nh+8uI7yM3DC0DzmXiGzUZzbCNZGfE4/JWdLfGJPwKXTXUI3oqz0OgHSF
XugZX3reMcvhqhTSOv81ZQpIWXWSvI02xHgfL0DAy2DIDLXLVQ+bCEC8/RQeN0L0
CFQpPv0xDubx4vONB8/qafJjA/H2NYbFR41yFUwyQLQeoJJl9lI+Fu/BALCgk0Do
Wmb2Ao5oNjr4oeawLWG5RHhfxPMBuNpnL6Ck/SssodsGQuOBchvo/6dWHXkJ5f6x
kkotj2aW5T3aIRb2EIGWurCJyfCirYW0bRcSNXyLRcTHUgzHFnpJEsLkrncPjcXQ
SPeMKuVRBffr4ubcPj7LHTwnFGzsLQVJEN6DXrY0hFqUY/j45SFwCXWlU1Q5+UaR
ik9bOYpaSEP+Sk4SMn9DSnnA+1DzMbw0LPkLfoiYEq3zu1oERG3SbUw+Z9SABwV4
uIOW+AggZapsZqpiLBJmPNARTzBV3RB6mPkTq/mnZrREHWdevlC67VTrbVm6jII3
F1t8qOGnUsalU/ZEnwu6Cafc8EEvBglRmpS6Tn9gd8tzv22RdTDnlUsDntCIdB8I
Pyjo6qEP4os1gY+xCvOptoxN/YfzZAEM0WAJomCoSpvCa/2sYHJJ3xmVgzWp9jv+
zOU3K0BAUhmvVHvqCEFrvuvp07y83yoaOcsAXQbU7vunABJiuFfJWcsJ4glpk+Ue
+XS4flaUUYkEWVCsuOKdaFiSWlaQcZUORwkzZoOkJ9Ec4B4HGk1bFA436VQXhnRe
jEHRdZRRqu5nmoDU5ouj0F9RVHMqBzGf4WWrTKmfOMe05rY2cWtMlKLTXaBg8bBC
ea+QShhTKsfcy4HZMoMS3YoWxJNNinB6n8h8bMRKpzNzmPTLuWduM0Z+CjzvSdAK
5+NRcmwWpViijUwz0rc7j7C4iW9wXdm3lm2IpR/fLZQ1dCG1DcsjX3yTu4LSndUw
QN+GEbGUaI6vOkEBx19Sy7uIKx/anf6gPgU4NLI10ut5tDYpa/mp4wY8LixNIXi1
7PUejgDbVPui+N764NlU36z1CgyuTOrY/HXU/GmX9l2cmVQcm7E7lhYyZAJgjlIT
4sDGeWpzYqJiHKO4cqEM0lULrqDWzVImRUZSQ4/YtrXmo33DtidBwRUPpmxHnh6t
7IPqGqhUAqu6iOaG9/xwN0LidxtNRJ2KdkEboiybMpoRlLxajw5c+i2LgYeyhooR
uJFE4MNall6iQJBMSLXilI7G8XxazaxML0KYAwFVmoVeRyBvssGCzPGdzOYbO6yc
nWlbFwIjGpHr1TtYFtUpIHZ0ujybmlucuqpDwWU7lQVgN/9krqMRPU7YVjALtlS5
F1bO2iLFU0CL5VAsW9Kd3wJFvECFRIvhsLFP1iDyJDHM1fAbqFVEPDx91FDy+3wJ
rJ+ZA5ZPVD16VqqQREkVbFyBmADXxO1OAXJMoOHTG3cXpl3W9QY3CkqUtJtAdmOv
joupGXLhBIg2HIUUEOpZyl7QCewc/cBo7muN1YWzQJzsSFU2ZE7BL+OuSkPSfTeH
C1Rv6f27rf4gGFGhQipQOsIaHUqikhxivl3dBBcb3r2TnijRNe1mx05drobAvxhq
a56UMEUDSyAYlVqjaL6rkRsRqRGgkppo3HSvFuDiOTWbt1W2YY+BRnGcKcELTbka
1oD3imFt5wY1R215jo8eKRC9r9xj110nEZSKPsZJHtUvm+LieKjQKEfIEhJDHvmX
yMG7HAirIVU3ix57TrOEWZ13kwPYxzIH7OkmQqTs8BuO0AB/KCltX4oS7G80ECpo
snTyt+HT9XlidAsgXK5IP2ol3U2QZYbYl/gW53LPi/e73fS/KEEvlPTiqraGmhFw
iOnUZdmrpaw412dd3ziy0qVCc1QdWYLAAdCuSlJiB59mgXkHd8o097ecK6cOncJ9
ntKmr/hEY9wVNNu6QbvWKWjxE69FTL3NMfgK0e169gT5KFSSOhH6+YQEQmupFrkS
dhJ/g5ezkKQTrAnsTk1z6At9zrLFA3B6uqBuX0dGpiSyhLfczSK9YOdW295y2rZn
QbDuUBnWHccPu+wGBFzPILmIAotql9yRZK41++cqpEZmU75vFKnF3QoeDks5KZn+
WUdE2RUKsSGuvlzXEtkzbudeJdb7rrNvTj+OdFM4ikPije449Az8EUA3Slwsj+aO
zihqcQAOg7k8h7afxaQ1A05z1reAra3fauo2dUwxa1qi9WEsG6V6TRD+aMXAFR0J
ugcuhVY7BiyzhtNSC0fm32XrjwrNj/x04QI9oEdG7+JKLQWdvphq6PFZTHv7z5GX
PhEVYXoh7+mpz9yPBfLUz+DVW6fwwTLYB1tFHBjge0gqOHD/G56oSmSR6YtjSkB8
+Di5O0qOKB0aQiHQV5748Er8FNz9m6/+MZJiPvBhAm1IayxcfDFsNHJzr8b7EZPR
qBQ06hWlsEMQ2T4SKNPr48VhWUAnB0SIf1u3cIpYBu5ObnZOAjK32T+GI2RlU8x5
JdiBswu48ukeCZqKFXSJIvDcBdCt/91KQtx4d1m+/mXbpcf9NnR1HDgW5iwTDd49
F2miAT7XnWb2RrHAJ84HbfjVa+ZoEVLgE7yJgoljDr/KQQx6f3io59PqLOtFM9RT
h9FLGyDKJ9VRyMFEMbDO9bRp2CEI2ghldv0GCEvciE/SYJypuyRTv0O/2aTTxe07
nzR6BvL3AwxmNLf4ZOwls3DtCcb54yTRIe1rW+KEoGrwCsqoggU1be9fZA+PiSsm
tJ3z57Rcet5KK1U8Sc3aWGZEm2L0ckaVH4uCUu5uj5v8wWNaif3Po46MvdNO6Zna
c0Oo0uhtUKZSobW/LFHGK317R9+QFFnMJ295pWRClZB+2bRM50AKR5OE3KYGVnm0
rObXmuSySodurj61Z7H1SoZmCGjgy/pM+6YWRZ1IGWawPFg6N+yy9yjAapAdDoff
4yY8l60NADVzUDvIrVdt770Autue3CwSqk2af0eaPogkzf+/3GA5PCuXVqkuITse
VvolvStb7S52VWQKHRPAZ5yNtUSPtL0YFAMjO+6ys8oKFLUWM0vyfTky+IKAQsOy
+ggzI33eCpYHBoatGQ6nsPFtTsYm9twbtVY21bjQ+7EssP/gpiCxh6ZRf7nE4srZ
vO1jdnBOHl1iCncU0qXDM9XAKfsisHay0l24TbHig+RRdkryFn8jCEaVpxQd40I2
JDUlxdRfuaRQdwWK+rnf4BNr9eP4ff36D63KLix5fsGcuovyM4HbzIzY7wH+mcT1
+pFSsQi+LOA/bELBRqK9kI3dQKu6BJ9+3YRqkK8n5xtwVp+AtYPToj9j2zRwvr3I
ftxwI2kj7xugovjX7k/oStDfZPVONHHeCpi/Btx5JioDd1qx4iHeY1ALsyhdUJOi
3x9Dt8X/iYo4GqQVTYQ13Ezj7JZzkopiaLrLmzinVsz77V/DEwSi2E/YZkkkhmUF
MkgUjv3z/0jCc7rRVckLp6rAke3yULvNd8/T7hFaMBHBPLrWVQFehzMw/p/d6fgh
PLrTHYEdW0vR9k7Q0nWmjPbX8AOcKWEvC/7e0t7aJn9h9B0inFyMUQGWZX5JPrvh
v2dhKpoMN2kSseLfgeTMBZwmHzdOSb1edt4W4rshLt4wDvx5sc1fGd3VzDD7uAIl
DyXx4ta+UTOV0OIW0cjXrLC8zHh7meLOVdWFKhnabOOyt/+4YRN7sGyov+qTVmXi
5Xv9DlK53ilysBBSDJP6rt3SLPoN173JhaEEh5DOCK7HmsBXuc02K5WZcVF4ues4
lhVkDL+spdh6Ob53FJhMXPq4nWtIjSSVnTyTg+Im4QEmXzQlju5z633lAbfWBCQ2
6AduwJapWYKkChbkQwk2QDXUSykEDaDZqB8s9axSOfjbIOHLQF939gfrDu9ixvF+
IlSOLNHRsegxTiM7ROoAmkiVKof65kFIkisUSjOHfjcDcq/KBq25og6aY+iHBAYX
vPLBvxcGDxqZ7f6CvG+3r8K3SY/9+sxN5D1yG2Hys47pwxErduXXHAv435CrcrWw
BB4r2caNzRJBqyEpHtsZWE4w0EJa+eM+NfLBvBr1FKrf1ShMlwCyB176hAaLfjnZ
KqwvZo1jwbx6C67pyNL0MUoIqwvPAFUeXsLUGZeN6+d4uFMxxX8wyP25WIz9AOvc
XqmtwjCatKAFPOR5hn71JgJI0y9wlcMe9CdzAzJRdBBlay3ijCuwktgnCkwOznB2
68ikL9UxPDmBswhclysucw1g7RYvIhSAS1p/08S3mEdSebKBIU690VvGDwg5vSbM
PlLnTPVGW1zAfAaVu+Efruegh8qt9LV7qCuh9aJRtWP+fOhvE7ZWMd8PubItNgF3
E4MNkCW8y3Hd5QrCDiWK7GNjvHUfVXmIjhnvjMAqqgu+Jb6PjvbEKLZTFHQiZsI/
iyxBJKUB8/q5x5G6ydAEGGdk4dUFkFp5sxhZKXRc4dEKZhWnlwTLJYDseY6o0FZh
JMI33HiQ1uifn3lwhGI6Bv9SIuBjY//uV//8YBI+FEEQhsVGUHsgJ31cauWYVskq
k6UlQRpk8S/Ql18bS6wNSahyTkF0h+5WYI2qin6KeKWVwJwOEEcSvGq8VcYHcj1J
C+2oQ2fVyC7EENxguD/VQBfmJSUFVU4l8XHR30MxJ+adn8EtFo31toYCi0JQMirt
JSaq8wxUE41Gl+87Ehx+VWNS4caMnxxC1Uu7ZIpCsaexjrDhJbrKvrfPGA7wAyMD
QdmTvHoHZqdAE/Jc2QIwt0UJS9GRnFvIX66w9uS921biO3NIdAOQpRzOD0w0GK2V
6jzfNlgchbQFIJttWrhOLZ6a9E8+MDUtsU1T7Urj//vUEQJsoWvfU2gmhZin+hsk
8IcuzPO3mL5nBqK64lYdHXPSCC/sS8A7Yp2DqgKZTYtywen5K0PBUuae44Zf2GXE
JDHF+I5zHBTrrHOuuaXmlNDtm7oy7/XwHUtejl3cL7U2nCZ4YG2ygJLntlbFUMCj
oyfOHfycNdShmJch9aywyXLV+b3wbxvYK9nhixVOBBYw1rn4kB5amsbQqZ2FfiZZ
2fvCkm5nImWQp59vXcMa+iCSAP7USoq2LfyHfX/MM00Qf559q7PFp9anzPwy/na8
5PN8L9YrfzOjdNQpPXOc8z3FcHEhCmKDDeH00ipYc8TRG37kZO+rfsRyXIxO9jNU
xvQE0Ud22lRzDwM5CR/VnsPUn8qJ47xgZ+4pfw4UGoXIe2vJHoh5nrO31Ahsn279
rKLPseC9iLwxBFzXizu3yFH38EGCrADW07Y1d9I5Jb8Xcsvm1RGRJsnhLsLRXVMb
5GnAjnKqwh49p2x9ZRJqpFjBkgBCahw4nFTO6ej4P9+NiUZeep1DI8FKlPnNE/wr
vXBqwCAAB8vMgWtwfq+Dk/W1RWP93+dVW0zYcEbD6C7NecCvylQO4KZmayXamyxP
dfJD1OZwPk8Qwd3EolB4nqHYw1NqgSZI4Ui9/mXwGOyUWcbSRw/Xa/Cbvrdf7i5T
1CVTk4NoFnulWB/LU89CF97TteThxcGWMMvSUkYYRvtuQuhIC2MG4y6dUOYu3JPQ
3dqmO3Lv67KIZVwMEnCon/QpzXKqR6u8aMie/AUCH9mbdNHsSgjMigWry9RNYfGB
56XYnyJAR26Kccrkt3OeHDdcv9adWHsOyDql0t7Lwb7RNnnwjH/3VdpF5cCnShPF
CkMrTlQTwfYu41AFuE7OfPKAgKoEkUi7KgHORySSoevG8PASPpJ2tGrizuEY07NV
YzztrThE3yau8fPpz3D6v/szMEplRzJKEfXYUBt3iA+bFbO+6ZytW6yTRpikhGlf
pJCs/X/7RmIr1o0zOcRuI42KxM4iGAfbiF9suVMsNZl57AstScBMp3uB1eM/7W7L
OS1rycUsNeupJX5I4R/dQISz8HNjkGw1ICvveq37FVB25pgzOfvtV3Nz2SGABnUl
Q2u7fKOqnTK1Vap2cNjWvXFQ1m3FK5YYEpRtkXfWiMx8fF/wmH9lOAnznJj0PKXa
DuGnZ1LzZonmAENuIe4MUdXpnw8BebbfySMMEZrnkXqOXGrp7hMydH8ZwMNad8Q1
0+od+oRp+5JQYkNrB4rCxItBGqIPVy0rMGin970Uyp7vKAZfeKt+1w2opyedhIYy
1E6HaZM9PKwVlAYY9kj3vKRWZx/LNfisdmAO1yHuTz1y9jBFtM3B9/TI0y9CouJI
ePNGtcU1r7VbEZJj/QehH4DxOhjetAe1vWFjvJ8t6haNxwlvQ9CLiSjXDGBiFF0i
q44Zz1TU/iFHQvAYyY0vAGTxfMy+xHE7qHBckJoOs6sYBp7HEALuWSDt1UVVrCv4
072u3uRPUMHMLsgqrZTntTpICs7WwXAAsYtiFuC2Lwn7CRiYCxJrUKFCBs90V7oC
hGSi0P7Fqoy28YPeeV/+aT0NS9cFvc9QNMCYovqKu+Rbl/lNS/I5uFsiso3GTNt/
2pTPMWJnbtuO/xN55kLBD9qE5Cnm8O7RbReh6FAeoVvaktrIYT0gebnjSaa3qP+e
DM4tKQYE6BOXklRNnvEDsOW87HBEQMlKX3rWwM7p3iP43DjMsPQhca9doxQA5FvZ
S3Neybf41IEe+YNqJO9UUbd+Dftk22WCI8F0OJnV8osHfaqCzRTHxIFdslZ9xNab
w+rPswcqh9uFQ+DPeiztncwJ9uGtKt9JN28IXAttsp/xRZjAD07NvV2Vz4lZyp//
AVu1IQqRQ4IxM4sqUGiXaJa18/tbaE432gfidM1i4RuH7N5aNupSQ+zHZ70A5FGh
kxy4DDD0ePVwJZy7/t8J6XxrS/jEChilWbkJa8uyuhtVmPrg4QDd6HJQw84VH2Ah
czi7wkiGuP64IVKhEh/c/oEiZt9oqQBNMQc07yUdQ/7Gd4ufCH1h87nX1pZOFjPD
Rna0d0XLPToYd10kDyxCoEjmA7jUsH4mMf4eEuLpN2XNcUvcgZc02igXE5v0bK1m
PmabyLgrl1OhEo+tjgpagqb3ur4r0de+zNb8f+fDlsovjwHsth1vxQAtDrjc2bAB
XGb2W9lQVfXC/R5Wz24SloEadZwkDj5aVIUp/q4zXRy1rjV8WcsOjR/m62qehmX7
6vu+swdAjXi/mEMHSDcgB3nCLOtZKytQCmX+fTIWWGbjFvupi+hNTUNIdKgt1OBu
q6rG/urXa1xxia3CIlrGG/vP11K2kg1mh+eQIX9vDxzYe/S+zc5AHW1ueLKpflEq
3UqCP81fyKIvVr5zI0LQQyqpN6OxFG4hFxd9rHdTrWypKmcCTAqkyyRQSmmbLBHd
/g5K7EgCb2lkTVYtDsuXciozKefhg4L8M1tOvjVkWgU+U5RuitAm4lLUPICJjpsF
Blw0ImYLx0/Epedj+IH2hp2NtRuU127MO5zSwBvBJgk8iFmzphC6NFmfOXpPGC7y
7nisPHAxjJ86cRvRMCtSliKSTlctSZp08GT9UnOYUZJcxRALs85DZA7jImHYjG+h
CDGkh5Mpkvj3/hpjHVRkF2vGLvv8LSi/1qDxQKtJ3LDtW+iVVZ0d1x1mrRbkEIXG
MUPSNBT7VZg7LpQXZqbGhv2qIaaBiB0u2ZkcU2bEXsfYKq3jKFWu3n+sxd0sP5K4
cnMKHKv5IpeBkWrTZqDqPReGH6qV5gNXFl/1Gfb85ypNHikkkxMQCsTdWEZRPmWC
nTuHNnn7IPb/rRs0BxGIlbMTMLZfdRs3QtKNv/6ujANk9JS3hovCxAi7aEKyoWI+
dcbWBXtWKtMq7g9AuDdHZI3ayfr+5g87Gsd9ZvoN0YngOg5n+Vza1WqGqi7BpoxM
3d2BuuOJVXxhbtVcRq3OyHbo88HtOlAA2tXjU3pAHG80SRZqsjOimAOT0Y9eyS46
iPl8jN2mIDA7r901P52sTpIanXB943Wb6s5aWEPgfJ/5xCxriWPMBd4vtFOW7IVL
IyWCOTsOLVGdejTucoLpkq9GNwcF/Gv8F5zUS/kIwyCsY6/NJ5EbS74GDNSUAq0v
NErISdHle18kwIDDwvvUVnDYAtUl/g0kjIeTeFpM7hdcqARyvaHKl7sK18b+PmCG
bUX5tuDl6QrKkxjqA9yQBOlkFjrrx9XmXowsfCYIJLPvdM9RcxJ24m4XOdBw6dsA
ozrkbp2vkjigAXYhz19VL9wcsYyKM5mUi71WPgMkBVLz1tdxHSttkCnz45fSUyBs
2PQ8L46fSRjnK9LCm0rgidLLwliDxT1c1pgiD8U2Y6jAOKrXuqBccUnF04dtS62V
bXE130tnSk/DOc/pugz4dq35kUT8rM6uUzTUYJlHTreZvISzMq0Oxi552zLwKueG
mO3FYdwr/aG9CkuMUf7qo0rVZo1vlPH5GBMKFSyD2YEaiMx6XgwBs95LFSr+BCmF
BzcsI2Qz5CrD+Op5StzLiYRGLz/KFGH9KvwpFy3U7g3ciS5Qe0owUiWJWGJ7xX+k
2WqXsrUpGIcd6UuRkWHXuBrxrEyUdYyq4flh/KD0g/X3xFVlTp8LUtHEsUwZQfV/
c97DAlsLp1nFzVacUqRoUlY3PoUqDL3atkrYqqp17w1Vlabs3G2F02t7/bZ9fWcm
9ioDPrlGAq1scUHfs4K/xcp6l9ba7XovYTbGjdRv1kFWzDAbPu6PSQLn8/GbtsqI
htlC93JQ9BZSNHbYoorepJ02wMphrT+iMV6JT+R8dm5Ck2CZSx0Ofv9qKnv8B9fD
Us5IZleafvkR0GlA0kkdXH/v3k26YFmy65MpCWsp2/Xnbc0B6+iXkEpmjag3+GMc
L1ItYEkddlzFCVeZYYjJIkAlaKskZbWPb53zqqiBZvl5YF5wGMxd3CODN1kwpxP7
kcCGxFYvd3LJXazZmt4Ne65tw1pxwkWaz9h+1IfWfiXMQPoJpgnfJ5pbgsZGUQvK
vhD/N1wG2V6z5/R52QKFhCNM92X52tfQ7ihFeL2SHMqKatnv51sk+OPlHGS11vkV
wPgX7dkfSQQzwFGDp9wbqlbuCF0eAPtQaUo5s+j4lRPbnv7mXt9OL1mfADaxgXH/
mSsyVtvg1W20AeTK7RrlYbvZGZubXp77SIPSo46eBw4Hle9726Jr2uGJpmvXQpu3
uXuzCCLa4GBVmJ5zQqY0f8kcnxHUgdLBI0Hp6aNs0DWQLsSoJ7eMG5E+zaUYLh9V
WWbSKlm3kG/6tMZrRYNee4A7qFLZCrdJ3YBRbNc5DwV56AK4Mmn2DKxS8t6OvgeG
d4zNXe9nNvo6YF7iuQNe903WyFCqC7IrPFRDy1wd0g2116nc0fO40izSaB6q3+c7
OkZaXpTPBP9q9WfnLWdNkF3JHP2C0W37PzeANzNdE8RIdMjZKNuIF7aWgCDmG8vC
x3ZB+s2Lz39o+oyu6KF79PAEyZs4bKDHqXzU2i4o9r+03lI6Q3GpBP+lv7MngrLC
nVoJeVg8HFnbWMxcOWge0jjt94JEuFqn++oSY5WgZRXvv5499zmgROcjuGEivgdl
VBAgi9+whxCmNvSYaocjILhBuvZCALTcsP3NhgZpE7BKU04hzyH19WIa8nFIFKiK
68h04KOhM8jQsQpAXFuhswT+RNuRXORnPUbDnGXVwDj4mMiaHj3ZulO1jKUt1qoi
s4KZiN0kLjjvJKqO9Tnk5EtRuryTq18FeSn06vzr6lDp8c1OKZMaRvQZV83Z2DQ4
EuuUlTtT/aFDND/BlvZNcaBwyr08YLNmvYpy5+wEhTnU805mIryfJszTtIjtkC62
qbpdGtx9tEPhLf0B806dlfRX89g+NDn6nJNv68BwOLyODKpc7o7Skj87eB+BSIw+
c46ySUMuVq7FEwrJ0u2LE0oBYRmv7rFZn2SQwG6fG/NZOlUFdVyj53nRaUvAqzPi
k/0e5FgU9dXNhC7wDuH1AuKQ+dzePT3JNfOzQ4l8PDbGO+dTDhhbYBbDFdMsugcV
Q5ZVMmX7aX0+nklAQTr77YPfGbD+vNT7a2KASsbFIYhEco/+mMGhp/qGBZtpA/ts
urF1FcG/gJ1MAMqnAz/SQKj1sFGPqDvS8ENu/00VtyYuN20tfR6cb4ZgVs4syTby
CxLSkJ4H32eDYw629vDTUzBqIFzq0NSuKLHneu3KFR+14PJN966j/FSlrJ7PmfCV
kqpsqeos11Zhjs4w0G/+2Ui+pXUnC7xPCYRnX6mK53M9D8rly1P8ByONKpnFq3hM
w5h1gYByMnWJcmjijwy3nh2747zO54f9fYHpW1zyqQv3TKr1xr3X6y12y4jD4BBK
jYnR3fMkbhQU3g0Li0bQfjmc9hLLDFJkiowezgKz1rCW7ptQtP4Gs8v8c3wuHI7C
gcWswoXJWQ2mzp7+3KWMQod7LlVkJpEiuzVqKNx/f24OttuhOWHIR5kY0zpj+LDM
bSxVin+8FF6zFkrBLapTCmWh544Ujoa5dtTrFyQjHcOTCu+bTDHhRDuy95tPx7cf
0bH8PGADLt5W0+eepIW8x/hWT7uXoEjEDJMQy/PZs3GlzP0TlGFdQ7hqgasfmqWV
TNRomfHV0Iymi/JZqPRZZiGYPEKAp96RwlvLcvyuzs6WbWsD5fFS4HmVvWneGdYe
u+RPCpfzWxZb8IfipN1zqeUv00muHnMJlJeviCetvKVBvOfmlU0LQCVYPODBLMCn
me25jXdjEVILdOMQP6zlFhjfR3tJ8DzVQwKE0mKM4j/xLABW6GhmT6+JJapF3KLl
GQk1usmQnMxc1gl998EGSKmycDEC8lSn9m8vlyGKhuxNdQiFNmKAIeF1wzjTYCXM
O8JI0mHQZAfgEPtnTO+TwlQYl5SCxZVKdD6+aMCS0m8W/IY2fDdXzLZRqnfNh+G2
u3S5DmwkPW/+S66tHqQZBOti5iACfwLU0H1H685lx29qJbbSBmAPWRdNn2wuz8ED
JzCXKsG/YqvdGIfKNhFpGGbgNHY0C7DE8u/2sxpDV/9T9IGOdWTvrIaB5CAPCW5C
wyTxoZrtVRLldH1MDM/FwpbWMtulW/+dGr3ndrF/QS9wiPtOEAVCiW6cXKTkb2cD
w/kyMHOS2EmUrrZSJFnBebPD+PTuk0zi8du8l89ep9DU2hLDCjvWFNK5OfgMaPEF
+LQG2bBZTBbLU9yVWlQfTFubdni/MbJSNj6fbQfqXl2OFhd8vLQqL7WSX6A3UXSy
9LTJg4TizNKS2Vrby3sMmYaGRT22UiILZyabAnIj8bR1xdvlARiyaIe8qQWgC9y8
u81ludXRJilax9YowSKltuNNNmpJKmd2koApzQQA5AMYlxsdrkCCe+1oWLemBgEt
E9RMFCb8ZwurULx0SqonVHvEzLUc/TdixUBup+Jj8lPE01PcjOopv8dmQmQNPrkC
anEOywOFaCm2I59bmfSKtcYiVhJVKxEdDyk9nmMwcznHR44p2+KbgHepKne6av55
5xd+XscRRof8Yq0an0rwr+skupKj7bJ5NIlNdadHDOdfb9AkMQgT129ho5jRvUx8
TCzHVou4Knu4yxVcs/sjiBN/YidCcTFo7FTuHALPtiU8i/0SSoT4hEIB2FshKEjD
0ckD7eK4au/HmyeKMCHH2AyGqDEdabkgdDWN5DZpKjxwb9vjeS2dILfICplB/pet
q+GkE0FFqYc86adjE206sI+yk3GWtmfmylTQQJfki9l16BMxI0qp661ToPC8c5Fw
V6NuIcFDzvCD9w+1pdhFZOb7M9q4j1LSoh2c9xJICtmVaDFfkhv1+OGFglgvSlaX
v9NbFzRNB1I2uehcmA8K2cW4bpWAjEgsM2gokT4VRtofJJgscpR44+eK7+Td2akE
a/l90DCh5yqpWgen1/92frkTn/F9oDOvUaliMdFsEZbfWBr3RbWZ81vuYBn9kv8e
rU9+hevQCkJFaBfQihbRYeWiByXWP+PDNiEJtyOcb30BPBf9ydCgReJ6RN4wDlYB
ZYJylOZiF9i9wQp9C+pd9wPn+8tKPHZgOPp9p3PwSZXGpYMuHCXHxJ8vnUpPR2IY
c0oiSvATVkYmJjIL9nidY6fjQCbHt9fwMTDWJS4Gv5qP5KCKn1tcL8jN2WJBooUu
w5qu2rlR7eXm+xZxJyacVn+m6YT5YCTGLhfdnvp7ljJTojMu8PYfinQsVO26oaUi
1TnRMXyheJFxvLWCeQ2sFNG+RdnQoVE7Xyn0mYIYHvpVehuFUaDgIVf15e8shfdN
GNqw4VW5bvp4ymvig0vdI4Ljj31EzmUifHJF+R7sI+lIJFNwDcD/lMXuYwvf1ipo
3+FpR8VUSAZcykjIb2vePmsRgX+cfaaK0dHpqEvi5BOccx5px0GKgxKbmD88d9l4
bsWY9YNO9o1KXiGbGJLnbegMyaxTiEyraw8nJ7pu7J5oFI7gK2YSFluNXkpc3CV9
UqAUD6tUWu85ztlP0JTfUIJ1U2zddllL23WZ8pouKDzPMq7qucOjwb01F3sXN0ic
wvXzqyPmNfZaReyTEE61ybAGicRDpdXlhsP/s/RnR6j8lNL6Po7ftXQ2nGg5pPaF
EdmZqIXu++UloGy3PC9eKAh9v5gdfYTl0Lkzu4vKaWI0VCcWZmgh0ko6GVfn7YEA
GdMDo0BNeuPqM/nnG5zSEYCKda9FVHcOJcfOFCtmxnWK2W3dbEuqet55hBky0kEA
729poDxKOYiy1bF1+UA7hGLanQIA+/uqw43ZeggHtifjLYlrPsyFKRc2FngVZmt1
evrq9K4wBOfHRgIyQ8n59Pi9r966gqZW8YEGhL0WHJ+xSUClurS4ae+xTLyB+0Z1
kGLNCh9vI0JkqCpobKR6eszF6cro1IzUpL1qEgpCKC7VH1avU845MEYHdj3qRMXm
tCw1a/f1TqK04HycdrKGckiidPc9sXr5S/dLgAHAxgsooFy/kmKyCOJso+MVHt+E
oAU9Je0jHRYLZKLZSGgTgaS86HJoMAXsuw1E4tLIjD5Fut+uOajOmdu0H067/csf
LYvClpOx97RMqyCvrmqP3481HgMTtgLxBXydyIMKlwEYv3Sx4Ml/T1PN+flSRZk4
jCvm4TU1vxaUh3kxAEaV/owZM9LKlzb6EycOak/qUTDL5FMf2QKXCPO1UptWle1g
zOCuq5eQuzLN65SK9IvruOC+u2YA045SFj35GRFDjH1xokgl6FwtCS2FUxusodNy
qlDX1aXFqinC8V+BaeRUemHXsbAa6XjsUqBK02BCU8kPESqpfAcm/u0patGFxAqZ
xYO3/nxozKiviphgT+hT70xWKahBJK8w51jdC833bV7PMSmxJgP0vhwUNL5zyoto
4Jl8Cllcsxk/G7qzQbuoll6Esmf72MEIuOggou8x8yT5k9fplNN/mwv8m6iR9ClO
CG7LFK1wMCa2Eq8DkxbVfhQvwu449K9VPBKBpt0+PL7fwGngO5BcQnKzTNZOq2fu
RFHCBBlZC/JEHDzzAwzff27plC/HE+lRu9wigvJXjvTQ2SVOMd7PW+HeFT5edrjC
KeUfegESFENLfaiJo2TBPZgnAnwmDYDWb+bkaNqH/oUqiv4yMBhY/+97EsvqMoME
oVFMYQOD/1Cu6voGIRAMWgdjN8/7z5sl6re8YReB4CZAk3Wh7HbBYuCWGx8VDkT9
GMW93tOj2B9ISjcmDR2cYJ7UTHBTrCIeqdej9is3MgDq0X8JebzGq0+I03EwUTmo
v3i2PPNVaGMNXUcRXjUEvld/KRsPIRlRh0eldOZ1NetLaEsZ4JuaVEtS7n5WW67y
C1z9SqBTcRFNZALLVoyt2v9m285/rIPcP6Ya3RE44cbDNlV3ysKTHkigO0itzT/K
C6dRMUQy44QO2sSULV4hH+yhtzepqmMMhGRzovq/8dzpxD4LTYZHDZC3RYQe8FIX
N3iNZQZPjQGrPZVcayd9N0b6PFv2fOWQsxe8QSDIDOOaIFP9T2LwFpyj94fkU1f4
lYwwpEB/MSMxcbOURBwy1B9fhGiQgaW0tKWApo8a7mIrjLVEMhC7/528vVP4F8g/
Heibt2Dn3Tt+eQTp8fjLpb54AZfjKuG9cWvgQtiusK/z9SUAzslPG84t3P4kGPsb
bLAAJME8/CfvCDtTck8Uubso/gA3KiYcqXvGnVqU8XlljV0MslLCrFwBAVTqoiXc
B0g8xM3vbqkxut2P6dpXxs15SlCF0bGesJbaiNTmUt5gkCU6mqPp6YFW4SvD2mg/
W0lNYNYGgSAqN+gvwNZK3AfgF4+95GmpZc80GowU2RKI9/g1/B2bJuznHuqoKUX9
BlMWoQjoPVg2vdUl8xgr6GpGiT2RfinUMsSUuPVAj5RNGriBwKVWoHdTkb0XsNeu
sfw5d53lLIvvNWc40MRwbD7O0UGz3tFbD9rjsCXxFJvOh4mtZzI646tY+oESgW5I
gjNxHs7hQ38d+qnlM62uoBsMvY9IsJtt/vvZQtv7AaRd8ibXOg3AP95SSgGCrnku
rx6DdgDrx3sc20+wLjN5AykLbSa6TzZyPY0ykqLLIn0aCspKtVSn1gxQm5vqC5hH
unOow8b0VBEIcp1cchiowMv2Ld+8tQSpR4OIR75OVtLoVR8Bhvj5eyHysRlOm8FV
bO5VqUqV4OqBw6lEAs30hHTz2+U6znCmSDGGil3Es9a4YJ6fWEU/Eoz83malLTUo
TyP9DXL5gXad70zSPDHvI5S1w7nTfLh3eq3v85MInXWwxRLPfBwWhnZA0+Lm5v6i
ykzViGXkUbTmRDFDVRIPUPOgyxSky6uuBmNnfr2CdZpoekQc1UdYLG7eFzW/pUF6
hBYgzHBqV8YtXM2mNzTx+89+SNazTT4ChJ6owJD0uJaRajbOMDsgTMCOYlTMf+jY
16rOPyi4ckh7f0tbbsDfKA6Fur3xcJiZyITziYpN498vKVAZidycNfu7qPZQOQGt
OEfBPgewM0GmxIG8il0BfoJVRkzdt1Nxyr/CO+YvyiAdZbEHvHZXI/oFJVO7TP4f
iMNqmIFpNek7wMa9MxPCTu/t6NO/zwQnNjATPxD/VXxEkabtRAFWS+wlfgGiQz59
G8tvZ22x0qjxVrT5x8rA2aq1PmH0wFpltsQHNodMDMrZ8KlWXbb9kDaMYxED/SdR
wKFFKuJeNumfn2TeMP8lCgxzv4BlhqAcOJZ0m+4avtNFusq/tmBE5FXi+dm30ukR
rcLz7xknEQYu1BVPluATqgPeZ/4kdeWPjWCbA05IIcFCYsDESxOl0MZusnU4QX6x
rKaIFBDSUwpBknR/S+2d2rTZcO/X/aOXCUQ+1fO0kzHdEN/GZvjdFdFM51g8iRDx
/I+1E89fvOne3C69JDYgs62sr1hozkhyeQSaVlpj5mmciYK+I+9lwzgnTMuZULgG
Pjn25h4xUsBb7x06aBLlZtGrXvRU303ukLATU7ec6sld5kFTURjfypxZecNCaWcv
Lqj/H+kq8dvcN6uclrrlODn+KjR8CWV855xgH27u2joMh82GOohdI501YtuhSed9
sS9vwcbqq6wO99izhbXDgDPzcAISjNQed5HwpGF5BJMwjKenrjWWhHKSWwL9h91F
Igw3sO7wNf1ra2KlzF6nAZgcPs4MUm8O8vCb38BV3YZfupzdITh8eyOiW3bHQDp4
EF7DCqqVafBHvFlSvbjs+n1cKmakcALY7r5MZQ2jkFiX8pn+pNpv+NoOx5jyPU+Q
4yC2Uwes5mb4mQF9bhtxhzo+JrvSsVHrAWPhY88/jYk6rQKg7fF9bb/7b5CTwmHE
m6lahUYckvtheb9ks0mE4S96bHQcwdW54XeXr/bcKAmTRYY9/mg1eWn56gI196WL
N5Y/YwFCGJNdsO3q6inz8MbefKfN2B8SMZengTvPXcxRgOT5F+Hq+emt0zUcE211
j6Ix9npE3+Prt0HfdPNSpRzYmRjaQOb9lplZl78kc1S0+nUu5d4jjvMjGSSWvAfh
EBD8qo5OhzMhfiSk1hfMmIpI8qBKLcFKbkxNwVue6dJNENp50A0LkuSIgudMZ2OH
3Nu08pyzThViEdgE/svy8L4abGud1f6c1gfW1ab6h3N45rTsj/A5bKdJTRsz9SJ5
xprcM9UboMA453K36QiZBkmHQyX3yGwZgj2WMnRA1oTOZqWo55M5PyqvinBmRSYN
YSQRPSsTifMGbAJq8STFEy4VVCDetIQ4IJHiTxUzEC4Z7tioVVZiKgVDaXbJdSyY
M53cCAZeLpDenkcbS+mSKdbvMf6lZPP8YwDUyMNqZhnAB1213yo3JObT4oy9OKV5
QT0GrmXfa8bkMIEy6rZRLvLqIy8oonF1ulP5erDB6I9jLkVxqZ+wWCrAH+KKkCQf
ciw4JIxEEQee8sNAbMF//HepddKeTKQDsWWbrEFRue3lOnTnzDg2CNXJ3YvVhhod
9YPboRqJnJ5vHOHbPOMiSm02V6zOXNUGd6IdvW3aBMU1rGhYAs+wog7EvUEJXjsy
XtVHi9tvtzQMHal2xv/FxA74se4dWOH9DNxvHc9BkjJe8t6ksxZFMAVliIXDeAOw
Z2lFQJnwPfsyYejiLgBw6/cIR0liMm0YfKZ2g4od69iKdmRRVk4w4/+8fiXlW67g
0zW9bD4ff53C7vWs05oLXFY3tq3sT1k+YJ+jYRUL/LUapHADSbqDr0d8HqQ5p/7+
ZUzMPcK8r+RW47L43EGgvfmBX6RfDr/BF+tXwyqnCXcUIXlaxLMfS27Dr/rJo1/C
U9s2ajyU0+o2Um0jn+n8vA6fdLDh8ENLdV9d+FTjd6R7xpDDYguGtNKSOJsjZCsC
VkDhcZd8e+Y3Ci77SlyfmFKA4gcemoHxZGTNzvFIQg3gXPeGxHrIRt/P+KKDKVPp
bWgEm5YVErhh7GIeYxaRnfrroA/SkjJGBEzy/kslAvZIRqSBQC93dctn2TMkkvnx
Dk2g9kaCbXhXmrjwcqhbrzgubO0rvpFaelwdJ/K498rh97Nk/CZUaDevjvP1QPlf
u9V+qMVE/InYONxBE3z+yINAyhI6+/ZLJURuNpl9UQt9Eaz9kw75ZZAhgOWbEBuj
V/x+44hznU5zEjcz5TUjEhPBTtbo376iGkjUWjgjAlsXOr+rAQ17F6/n5SeywiGK
nb7ZJBM+dlRsAAjWjy02ETAFTvnEDduarq4GwmtK1BYA5oCkFENc4SAf2J74xUTf
KLyfYAbBO8TSNf564vTEPkQpuX+YzDXBzxsscB/H9dKsTge/Ue2IQSFQ8XcnCywk
x2RjJ6Q0r2QxYuAoZi6ETcsFuLzPGvbgjUhK6SqDVjRU+4kE9HkihxxEH/fGmya0
SMbA9yObNfJFCTWwEsFwEkt68/RVNcb3vCaC+7cW/YNrlMQFQh8jdcdaMPZUbTZm
fpM3KF9hIxG6PS5St7aitAvyFYmAlp1xDusxw+0m+rRKSswc6NCtYtBzg0GnS0In
SeajP1ngLE9DSzvZf03jZrHqM4bQXoro9V5gsPtUPWl5oIr0Q5bnSfpo1nlFelUy
yqkYn3B6/2AZCG0HQJ/16JnkuKiwvF8+qchXL4Ign7DGQ6s6MtR158uAMeGAd94t
DlpxG0mBgsRWDDXllW4E1Dj8vKcKKxnzKzNo/vqiDnH1q3+odl/GRGaazBaPeizI
ZfWGMUTuyLHrlulhyJr/aKYYyXMhP2tjC4jNg6afKnTmYnDol4sF7q3nSp0UeG6H
9CwQkHT1TrlJA/XgjfAnnX9goWR3MXQUUCozIZjrXxGAMZUDwLIAOKh+c0s4DyQo
Yeo9Kaq/2OeummOklLzor7rMESNNcpHkB07DAXnf0KJlacmBQx/zM4riMTMAjD3H
hfQzCtl0O57TSMpp82to/SEMQzAEjVZH2+a4KFJlJfsOJmUB55CJT4LpqNaBEz2I
7DRMw+Ba77VhNXJR9BB5irrt2MG+BJlluaozpNK07hCqgeYIHf+YcxQsyPpecIHY
0O0TjqVfBLIMh+2B+s3mOX977fd1JrwQzSi7AAFYzAeDQO3tflvlQTl9O0XHc7va
xRLd+hGeDoKRwkyW3axdm/QhVWNgYaTdhTC3ZCxCKSrF/1M41p8zBBSj2DdBQshj
BBspPac+NtkrtwLfyNmXasPDukbulP5EDKBBTBUg4z0OieTIsSEaP89BJq1V4NHO
fmGAV1F9k3CqTaJ+pEjL+lcakpPCAO/tiazSMDChRUrxAd7ICzu2vp6X8O+BWCcv
dlNLAgisdjAXhItaLg/AltEFpUNDcAWu+lsLTcvf2CJabl2nwpNnzgsZNlTF9LCs
p7kr/Na4CbJ1ohbVuTIVVk3zXkO/EcJuvx1waJvOjj6+l2Ty8QGkTZULRGg8Cuvm
/GJZijwkCB+3UYw+qKq+CdmGaGpWKpiIteKg2LemzfzakFk21a8JVct2HUjg/9Ee
qX4rILMaFYpd8uYMF2/zWKaDQMwiwIpxlqYaMDBUjCnW23K5pJAaIwjqVWUJRvYo
XsK+ePF+bc5Qb/SYmwNgOF7oLYwbtgaRM/K4JQespbvzmDgyedLJ/1avPBbwVgKZ
jbdtoJ1qCpLsym19mF1XiTjUhT2t+heHTuoTwZhCSq7rT0RuCm7bn7Wm8gIWAUfU
g6lMXT0i7upSN0OsJ8cQtEu2eL2+5Ujt0vUUj81sN8sMUubyqiK6BLVPkc82q/X6
OZ04zo7Jv10ZOcl4sAccdJKaamU+baVNw6Bjz457VYCa61twpHZzV3lh264554iv
2x4N33Ts3MylaArVzxCM8/EkSV0yYupvmGqyIXBVjbKrArp0hW+DCL4aNfsWLTw3
BdTqUycQqdnO2sXIIfJYesZpssKt9cRGsr2HoLiySDpQNX5wuWV6oCL2pV8oFgr3
LIq3YKUOypU9e3WG0aDeesapPHbKmiEJYtrudZvmlWjLC84GQihk90wxqcvcX9b0
1WpIfRVNwjOPcDm242tIXK3uLO9kLJem0BU/vxfRtG+aWmyL9SmGROgF/8PWhpM+
cfuKrouybJ9dcEdg8dI35fhsCqmE1Cv5YOXgXGaBrYAVQUSmHfayEYXcOJLeEJ4M
mlpqphEwNmVflFgDLO6eNCsMTW0cXB2V6K/ZkvgtX9pGXwLWxRKsxBS0BPLgsmNI
PpsRBXptHESSdK285nZzkvGoD5e7te6IKynamUVU8s5ReMmclImz/2/aYaF/ccrQ
414qOW9VvnlPXcknH0HmG+IGq/S8NBKbICiiGpLN5K4CTKovpkyx7jMGAsfRaQJv
W+FfHNJi19/WtzS/aPNMvQP/HEAtbG/jr5fDd3O1sqWCQPyOwe5w+lC7cXu8Swvg
QwVV6rAR5n5+DaiKKTETOOGefCerUTV7dPOanPC9x7+On1zWaPKu3fYbGqmVeJQw
sJsL7YG+tLTooqwlhj5ux4meGe8aPY8goJjW6OMhjsgXJwfemiUmD1XlNin16Goh
YjlZ8PlK0PKhGe3OoMheMAMHHdyffDCryxP+BoKfCwbKPLmvT6AjUPL6uLnVioS/
myXGi8W3FX2CmMKnNKml181MoTW2xNXM2tP71UDkrnlgkYMTlQPB4RRdYjRDh41K
zotZL4uq5PB8AhMzpoXHHVhMmsVW+GBSiTzaXvng7qu8BEqPm70UOvvf8/w4rbsn
mn1D2gdO3xL6eFvgRMn2ocnMouMC9WoTFLq2/Qy9D/wQZIMu10WN6uex8q/m/86v
olMkqGG/SS9S6TpB7tSl3ttB+lSkZn8ngW+TZQdW+v1x7O9PGrivm5kZta6W+B3y
sVdU2ZIW7ZJ+syqdd3OCUVO2j1Bmi7AgiprwRLIoybcvzAzPx3uWsYMVl5roLFkX
MGhGBPjxCY3+RbneMiHUgs4dLkdCt8atvsT4s0WsI6VtAfCFMfvzEOMGRT37N7eU
CYwdbqFCvH1t+lOM6bOMKI400pgDrjcyNug9nmUTulGM3PNsOVv7MpO/GzD8twbT
mXk+wA0c6rFa29XClN9VOXgeZuGJnSKQafBbwlsAu/MqpN7BzDXwd40RankucnO7
Ql9JQdD7Pu++7PF1LVs+aY0gsbsQYYfrPdsnkWxD7AHKbQoVjg0UCRhsGtf4g0CE
6l0vS3IkTgD0Q4fYzknqVf+kTOLyPkpOZIIOzfHiwiJmUVrOtFSfV3IqjoA1VOwR
Q1F3wBYVaKtSKvVfRwdrOplyZPoBumr8WHIkyM6/znp/OeZc33t9s+O01guEtdUd
N9ccLZsuMf5qGN+1WtSlq4ZkP41pZWugHWDXlmGFxArWhHLjjwujiKgWe7hTZYft
qpdB5T/sSIBeqk7SgTWPDvnPvOYNiuSkiMDjhVCDaMBHihF0d8JFmsV0kQZbqIYv
hMzJM7YASQeIEi31FmDIeyPDPqpMsdrZUpZAVaxi6bWiIqk6+MCB9NPEkpjSJzHj
hsAN2WHPwA+gfVphD8G67/ZQOoc5E8SpLxV7LisGQVoomOp8/1TUGfQhP7NgB2kj
Nj7vy8qqaByig59T/taLfc1QjU2QStsoB0xHOpKFsEZewlbtF91MU2nHQgdm0kVI
B3aN198CPvNpcxPByMiIRKwotVYam5OZ8oc2o6+4FHwa45FxcFWVcGmf+bdIbsY8
lp9etCDoJdtMLcXrT/5ksuJil93CPE7fJoqmeuEY0fVFHQgmZSMFx2/mZkKA5YYt
NdfnzwGDn5f16b1y9SHyOlcEmt5RGe18lXUaZr7XHhBu6C4Pfi8Lhn/qotoRgNXm
DgBxdklEXCUw7Ze6GWWV18tQ8cHkGJHltWXx5oU9ckuMHAGerrrYRi3+rySvhieP
lYgTEcCE+8YfQMqJBLYGqEzzXSvTRstWZuWV2eLWN4VY/qKABZcEf63YerHbRr2R
5oeWgg9TpdOFCgd1uaAZ5pWbFXAsbzcvd9eQrsLx7rBiafeFisP3egxRtiINrhFw
L25Igq4ZTeY6lEi6JWnAdkr0gZACc4fwLROlQaVYcC4XIqr4ggwP3LjfjoeUyxy5
ZTWlVxb9HojJAvEx5yb8uSIIgh7A2rcETpnVMBTCDWy6/dFU5PLJ7DZcDjcy9Rlx
KOxnIsXXlg7AfRePaV9lUW9EubX8XFK6XxvKKze/MnYo9N7A3lYYjkcoDRTL3kAi
2e8YX89bKYb/xB07olj1GHiOsyCJr5E0RlR5YHuStG5AMtgVwMvqlgTP2RiMPhAr
xb7oBSF9CMxpPFcbjztrbBIXwC5dwIoGy+/Cz4y4LdGOLcGcPU2+85yMT8g0GPrt
mStZP8Gx50GosOF87oa+o1p/XUY1RIpYPp3eW4PTxTpMf5hH+zhX9+9VSx2RHXpI
trMrhw/V7VWxwteFN5pbVek098bJZ3BQ/1tejcSicqMVGvbTGf8avdhyaf0exN88
PFETI95jZyYEd+Mc3x3ND9zQFcJE1MLvCZYYlVHZwqCxpzyaotiDJZ0yogw3x79d
RKkGLz6uIuj69dOkCytTYMb8vtAnZ67XNB7BoAKGW1qC0I4KRz7G7lm8PLknBoDD
2Fb3LsW4G6AZk4DPwwHDrCJazu9clBWk31s+FN0CoG+1QkmDyPtFL8BlOUJsfU3v
4FQ1EvLgvZKVw9J2xslUTEBSXw6VmYv8G/urY5EjNxlirvpsF3v9TXUTYZ3Gg7zx
r0B0Ssb7KSeNyXz4xqgWYPul9o4w3KHcGnCCr21BETfCSgs042S0V5XDf83/QThg
0oKJJW2OT4GDVk0vnHCQ3TcjyMtSTh7OBui6lvf3S1MJULZeK+PxddpIZVMSG9KS
3rQ8yAw3+xMzJLPUHBiY21jtAT/jseZT+entsilZ91EgKK+rZXYLOo9onbPPJslY
qdQlHPOLjYVaV2X7adQR8n16cBsF2Zjk10Ox5c18st4409Cu9FnuwlLuTd97Pcg1
kWndAROJScL3LacVjrLmoXddGGvf/qNkByxb4a2J6O8AGy+HY/Omsx8VfI1d1bMB
P6z07fyEYQa2nnfCmImsxfeE1HcC4ax+tDm0t3EQYA/nSVaOwPVNNYGewTNKYf1V
Qgg+v/vcrboVX+PcC/vBeJQR8emLNIRMCSHyhrDFJtAZecCYEM0IwcRC1mVX63Ix
t8uC47peQoto9rUWR7W3b6St6VS/VatVDVEpCP+VQa9vuPC+iSrHbIiSABn2urJ9
N0xZh7YZvK+7IdyX5HE8DKAdpsWXH2d5F8zfLHar4eEnHrBKdhDXccDRtuRkW0yA
q0L7nppaZhrvPZ9Glb0/j2y8ju9pnuEBlRiNaczyFSR8Y4WIRNwGnCrwkQT8oTOA
BGEkFNCigHitpdejrHu6Qf4aR412Kr5HD0Blu6LhxPUhdfkEvTKhtc8wn+aT2CH5
r0S3aSzEl3WbGyzHOrGC1GTaWHU9xQjIRHp5VB1zXUlhLTeNLaEDlaoZ4aeTtM40
JRbUiQiUgrypn9OTyEzghmtAwjfyoeaQ+daQy6pHcZi8BDuOkj32LcEEDRJLk6e8
aam40STyTfIhRR2AhWCR7WWbfyUV3SB/KMLRbtJALJejzzF6o/9qvxnxLv0Yi9cp
Y8Aj3DQpyFz0zX16Qw/unkz511ZKm9u3bXIIHOfADCg5FoYUlaXfEbZrpA8HUTWA
eapjz6AQMH12j4cEnZ3o578P9gtzvSkRhA+jfsIZ29A6ht2xCL1dghQF0saJAvGK
6IgJXAttzqGh12xbvHN6e8W218wBLGAPxpKvf2OGavVOumOUy3dDYtewBr+WJdZI
aR5vVtDgtrPFBogfQ4LMinnIUkfsvYIRZwJ7HRNy3ISjk2h1FMIwV15giyzx3ByI
lcZt3wI9Jy6gEVwTNP4A2oHCsj6v9D7FWgOa3FM3nXiQbWRpXRIzyEppLlntjK22
vAwN4adcO6jctBbgpVkPAELwQrKT3MlxbVo83K+pULJwzkeKLnY+tq3CO/O9tX5W
1l+0qq7lTWXw2qk3GpAMmiFZnZiCmq/SWphzWztngILDZQ7buTXdK/3JfTFUuC80
RQM6ueGfrRZWsgaWEFE5qalZXfDbnJwMDuxDFEqOzOjn2UeCHOYaj0OWHmLLFm1I
SAr+8M5fMeoVWVAQrqo3D9JGJjlUz11YSzwQZgQtjzbTr0QaMfmUECYD2ZeD+YIM
y2cPesZzYPIL4STsPzCMIVvEEycxI7Rk351YGtKUYM2oUyIz1y2wY1JHqYVlGMGH
+JYVqHta6PfXQuzzCZHPhFhOk5NO2zYEwQUMn4RWxdqrOmUaEOOxA3/VHrjLVIer
TwlcdfFUVWPuVD2n76myVYqv4eNx6SUDzLZBWWZ+KwxuPDxbdKPIla5cODYdsrS0
gVjKljz3CEUB+2QFc7mSTh+uezdZJy0dVep7bXOzb6F/GQrR8lYZiChsQjk68qc1
zI40KML5QMmgQFm4XApHigGvz8R9hhAH5CRHvywXFXgBUa4tVC/c7/XFUMw06aiD
9Jrk+XrUH3TYXTa5AwoFl2F3GRH37yslVjbP0eTzqwFgup9TKnEmKttelTEOicxp
7xJnsd2X/b3y3wAW5U8Vb8R5AVX8gNVQRb1FZPgtA8b4/eHK0V3gTCPygsS248XR
PlBsgsfBhFfv+8RX7dFku+77EK1+PkaCxHldjKdtgrHuv5TqFjBM7dz59OgYnUlX
/EiNnceaEzjwhqMltAjWCKRPwO0EP6RsTYUxncj1qcrGMSmbNNGO2+pPg/TOQFBX
WsoP97lgYXQXXyiKh7xTU08Pw7EOlRVi1VU/4F64YMYlly6GRfZAnpwkKPjMQigD
MApmwLSpd6yQ1NSlLHK+5JxOXVupM8YgjhdISCeabJo8qI+MFHiIRocZWjEnHNOr
jKgAflGGmoOhe++M1z2IGZRd+TlsS7we3j8iuPAqPk7ORD04wozKRM1KeGp58yHt
WsEA+EJH6BwclkhfZNhfu7CvZYKYg7berdHXvWh8VNpVkr/gRuTXr8UuFYBmNyNm
AL91J6er209kuS5ascQ9j0lIVyjnoCHzlz5vyG2GTb3jV6U6jtq0U2Rn1a35ao1L
Pox86NqFOIn8fmVJYlowzp+XkpAFAQGGmUz4BuPUCx0Max/e1B4IW6tFqIqEUJ0U
rbe+ZdwiMaWC44MQZlBSDKZTgmNKJYWBaIcjWZ257sYDNWJrwCN7sf/rv3a5SrPh
WrD+FqnrThnCnIhzG1jHnJXaWEZ+b0mSz5vRsFoeXS/IWYLpd30U2v/qOH/YwBfn
iDmAEfiq/uhYwQMhEJvVH/V8B7vvKZaDSM3zKKjNayy99wZ/lUQwCzXALxEbLrXm
UcZ7Q2xY8PN4tO9wMAD9GdTCtu4MfpevvXir7KYWUv1WICVBUeCmcVDsrImkJMTK
kUacSJ3QnMmu+atez8K7rGiTGNm9k24+rc2UReXiHN5jRgGxWEhjFA8cSp7j7thT
/ZfYtMKDVHBVpmmmgP/2N3pXbzQFcclEkor+ixnqKsNBj78wZJ0ue8iPjbP8J4oA
jmHocjc6DtYyJqeV7wyyARnmus7eedMJx8qps+sDgHCGYwPPYBapACNdUA5llX3o
Id8zB9Kz8QDriIa0KXsipZvBVXs5o6zChMkQ91TQdteDDBtnCfZ5s71C5u2AzM57
h50vkGDMzgF+vogxP8Onx0nb5LtyPmJUmQIw31qjWGmiVbN3F2b9qELuYt9jOfyH
tKtWa/X/woWZ4c3amyIF1WCBN4adGU3zaHee52iKdF4e/WIdI5Oz+ht7tGWxxRlg
H9lELEdkIpcWfTngaNcI3WjUlhQVcvkohcJy/O5Mhj57+azZ+3ywlosST5JRaYq7
qmh7EMvDG1kLzWo3Ih+fkglOM4GAvIN6lBmHxfSpCOjqc4ZMw/HKTTcWyvUEt0jI
h61uybmGsNS4Ps5UvyvV2IYo3si6gmCxx3trI+XilolbTXZJgfzSyZCCVt+AlMj4
jh3vwRuCI+/edoWOSh6+rdbbJA2/V9Yfscn9jh+vd2LGf2DUPCECeZZTlJFQTa9C
3r8dzSeS/Ga0lB2b0JBbfTROLMh6QmuyhWSpxnOnM5uFnFfb4XzessknG030JXF1
A+BO5rrEYSrIlU1hmNoOEfBP+UpWA5jhhfyspL12N5aRYwJ4FI+9ZMIz0AGSskWj
Q1KmdZLt7JmiDCv+5Ia8XG6X/pCAV0CNEHifrvLqkMKi+XsmrIbplww7dBa/VoYm
BJgdwGfKG6Ag2VWzNu8znMOk5XnaXsuh9Iy6fxIq8nuyWcjBqgQzgQntgW3PF3To
D2B7nusfnUI+X/KqTpyKpbxw1mgnnd69M7Fgd1JFsYHAAVT5Sugsq7pVW9Hf/sMv
V9nEOLqOKlEW8RLwe6/iCcRvb2Dwi/T6aq+AuMlY8V1+uktqbkkllbVxvb5oWL9Y
AEvBjbG8rRmXKosu+S36wuOxtpONkQjYydSkclvxyIqapvkh3G6tMbhJpG6NMnZJ
F2sPy4qJe0g4PgNbGnKDYhpn0xfxIyVROyx+NFL2nFFKixBXQgvEs0qE2lFayzkq
MVxF6n24dCr6ttGBvIyQQwu7b9MMlSnu7DB4fWr6rIq99Ns/P3hm3CqFb6ZqrOyt
+ys9LijIbBiOwdzm4S5U3Tu23Lv53FhM3t3YjPCOgm2m4O7rOmQWa/5bAy5FpNWG
L6+WqQQ74Q5sb3YBv+OW1Lq2wU6eq/Mi8t8YW1A685JPfnesHi+P//DE4lex1pIR
TEYZiHK6Qw2BAto7utQDsXgzzxXrl3GyRZZ9GDIGyi7wxEhVF8n4m5WYWKf9NZ6/
XoB0woW5ok/PFtBzf5N+voWGoGFLQeYvWe9v76s3m3GqtKpuhcH18BBM9Fy9aSMP
Yu3xd+2URKMWkqcpojtA/jBbYYXdgzVmGvxAJI5chW+ruOHgJilr0PontPG6XqZ+
DBX7ld4V/Rt4hVIawBiXOpkLaobxUl2e3ONk4ywVgntDyx2yUmn6ECVa0L/C+Uwz
nGXg18zZwqS1ssXWL5esKcKm/FNv4v8L4fDX8NB2l8nlXFLSreB1L7YaUWYeDLsT
icOXFknfKK8oAW3WKtgqafCJVdqTHNUFBJV5rT4vSWI5q5yE9FyrDOVbBKGw348F
rWDplDgqFHFe53Mi7gH/81+pWAi4D1dqvAJ6STbVOmCefFVKw2kozyZIOtYNNc6u
CoTkGGtys8JFu0cq0SZ45BD851fHxrejZ6F26tE+dSKBRrmRndSSeudUMFM3xOE4
d0prPLUq1e07Do3Q8dFxBovKj3M73bbDOMl0XxR1m1meHRH6PV8BKGehDRJoijbV
To0XRqKTqPFo6iW+JQW3DEYOyxdrgCyxi+mFPEMFv/zl+SFMvpeLciPr1NVn4vns
mhBkMYvvOCrxn/Zo2NgoMM3grmYu/wPvgcn3Vunn30XahF06hJHtp1XR0xOF8to7
TvvDYMwfZfeAqQMNbRnha21kwEaxisLjRMEpfOaH1izVb1PiZfDwwYG4oQr3Afzl
E3jE4CiNgFoyGNA41E626T0UlKuh1nbrXi5lljqS7MR49xZabzqMhEdpYr2Y4w3F
AgQRNvUZeGZJ9rPdYU2hYvaRLNGFjl26QeNGOhBhvAMFaKb+AFScoGV1bP83UcLb
ooGFNpVp9FomYmFnRtD6rmPK6yHtrbT8C5nIlr0kUGkygP0JRE6jxCCkkknK4zmD
NPgKQ5vqDcqEpxsxpxB22d0jtOg2UJliNzSOctrclz67nsFYpmwIBovCndxdtwLd
4mocCibp+/txRGlH0enpAJ44balJl1xBKl7wnhHi2yLtqmFyf4qdugn4kui5JK2q
UaF+hcd+p2AjNIryAXjt0HvCPaa6RlF2TRtQI12AD1xomZ+2ZuAnTs1/jJGCt8a3
jenT4NWKkZEuSqkG4YLKYbu/objmRu6dWt1HZkC9ZszNNxufN+DmRFpayqNfNtR8
QA7OxOZLC9DIGeD7kaTlTxKaiBemwPKSsNe0KWYRzFqGRtLOkAfEhI5CgFzLOotr
65OImVLiX9i7flviafOwPQmCBGSsGov2zX2axXZGEeFfpkh8RmmDHRcKXayk+KKR
ywhZANa7qyoJ6U45OY1Gigsty/dEwkYBOohCnLQlmFchni99vbUO4+Y3992mMXR8
TtaavOMf2Riq75C5A3B7VD+4kie8u0hNGdAibO0Lg4MxqjZE1VZVAD5TgQIWvsKx
YtUKkSF/ljXlwB2CwuO2w8c4ZTCNIGJoAhHqFbHt7C2TjmXuvsd+wQh1CYUDiA4a
dWPdLWDEzweg6wi+4ltCLFlh5twSuDkH/U4YtdieAlbfFpcyJ2BKAA/a+3nXDwRn
suc23Qwm10VoVmK9idTkcbAhv+AFTaw/qLgIjJm0wZb/V37sgg1f/3r7JNRRswcz
xiMZGAqwD4waDsLIPSiFLSSs8LW6QPALuFrC6XW5ScuYgMkajtXRM52nejbFPF9d
xTtAldl6JtrFNjJ02vHoQ7BVQvM0XZmrrZWja/SNQ6A/FJ3l3ywfEkN7Qdg/yYho
+RWvEoGppcgMPpt3to2mcIAOiB6DXwxKWE5NPs7COK4joxU6WNquyJtzaZuugFVl
WZ5eDawYyOrtq9Jurt0yWz1/NHVV5f7dgKIPVQIWl+dP7VuR3B6Xa+vbv3coiG+e
4oiCR8iXiz8BcHtucuQG+G2xj4Bl2hk9VV41DXAKd/qdfM1ftme5/Gh13F+GzwNr
dY0ekqxlyCgsjgSQLiXhpYagcS/rplN1XN7DoJ5fig3RD8zKR9snw6m7nB8s35sF
eyiTMkUD7IZ08AOPUcYc50wldjM/mISzLeesNS7TnwHEWnfM7eGMo6mIt3ZUlwca
6oWIrhoW5/hofkRODaYFONN/OzL3qcyYK31S1Q383+t98y9gnQWvXndD2bJ2ApMG
I+/TmrsHFzee2i3/cHjknl4qnwhRJOr0QsHyrVHLtcdYt+RjtWV+Kpvcq2PNRyaN
kZt00+6/mi+FvUmfTnh6MYmiqf5Eu9rjPT4gAoO7V/dySmdbweUp4VNClGrXeopD
DVCYCrwUBa1TPn2nHMFWiw32VoVNTHnTb/eFESwJ13hUdOgwu+IpYGqSeNfnigNc
DedZs2UHHb5XeUS+gbs6A2OZN1mQXz5rCFI13vFIJk1QARvA/tBRElQan90sP5AJ
mzwXyqv+krDa1Xgw+LNk7cuI4b6Dkp8i9OBuafVOy5m1oYKTZKsooff46/1WQMo3
POEMZusRiM81FjM7pU2f4ERoiCvxhgu8buNAgEHc8AzYlxcaSgyAPrfx0ODry3cW
srN/tykFu9O2Scrv5hSQymwS+m6xYTf44x9jCyx4bgtlVZzDp981V0a9CWogB1wY
bLYGujXbNzbVg6sI909JXMggB+P49m+SiS09Awt6tbkkXn8PUrLwv3TswtViCuMk
6FZaTIJ259KgQr0PbkKpm0pycObIFqk+mmkFyyLReWlBqpu/d6pDDy9jHM3UPjal
Ok1HjIxJPI9wFRHPVPv70lzBdht4ePaPsZ6+BO+ZFnasBrHIoqJixMzGC7Wx6bBI
G1d+qqXr0fpFsImVW6NbJUCcCdP7iuguJlXqa2vi2fth37YgZzNruYszI9jxu+0G
mluJyYCZECkmgsr/E8cCjYuoryRP5+liRLcoUsisXayQPhJ+jOy/l6NotUQ1QJ6o
qQ16OfaCfGU+ZGFM6BTJdxinUKJ88twX9qgsEOHDi1R73e/vk/96Me4Qnc8LwNzV
FYgYnWekFwz+vB84omDILkMcDN+pqS/GYEYJPbhkIEs9XbmlfgVZR1hc8QwcEKbH
h8UAmLFc/0KmXbmyDNONNOU0KaSzvvcy+Aevs2++QwjSprrZbxTC0jYz0AeiOLGV
nNWrp8qFDARsnC0Qx//TdqdrBkTQsljlOaxaY3d9j8jIjSl/LWPEqAGlbC+ePis3
FV34ams5jqYBkz19iCQejgEewHWirA3KCE1BN8ZTz1KqB7I27DKvBCjn91YNhoNC
6Rc9pqupJfg3URF5V5bBqKLoUuCTesvREyKZjrkr6uk03/714+xeeVYeJ2NTpxzG
qaCtoDYu536spUin13I0M6FwxuzHbbT24D2FsulaKq1aWdfwO9TSwOidMI+3nLYG
XdM2FY5kfNTggzFiH2dkjH1BVwwPQY3rjxv7/qo5Tr80TZ9j8E3lF+0dPjcrPYew
WydZ/aaSisGbvbJmrFStC9yJDYxTWA5ogi+Ky33xk9oLejIBjBMd+HiHrTHdcgAO
63bnBobOqefmance04oalUQi6bT1wlbj+QUHIWP/XNjMN8JpHQi7AogYVZP88qHG
f68UqjKEBgzccdCLL6nf6D2I+vqOVFJWheggJbZ11UVWSHaCJy78IIrfC6acUFFV
zuRvTPneqLfh9VGxe9NfOzUQfimK3O5+8ZZmAWlM5uRbXVw35ugB/51sG3rmNxND
P83+SLin9kfgiJZR8QsTTMSTPuzIPFNruUiUKBr1RT+EmDijvGTZg0jjsHDIjF8y
rUwAUW/hfrqgDDwDjpN22xFZpvX2IV5VvSAYT1pOiqKwjOPB4kghxTotOUCEbJ6R
dq0hgBwXMjG+u96iZWpioEjYv/cjwu+2gX7vAXhvR9SwUm4BYJglz/eTMqKMBjnc
m6ohe2kiBD3zTbiKj088+HewYchTaVFQHpPWpFUkwxSqzvGmG9bE/6RI/ZzBwy4T
uaW7vmxPHalDsYRTcxpjPaZ2PCizHcVBU68tqp5A5fbB6Igla35tOXYVeqK2lZ/a
J9rfkgWbD7UrOaadlSFKJxe7N4xfflfzrrCRY++F8+ndoRHf64h6gX3shAZb0rxO
hYwhXRvjNpayxPxE/OTnT0AlZnzmAzNF+qzZrtuo4EwKSTplb0b9Expp0rNvDhwf
mpgp1sqW7ZoZ3GhmgpUNMt+5aORf4oH1/UlumjdyPh6rMiinj9qIMt7dDSh5G1JW
U619bvLnDjIItdFlxkNBp8J4o0Apj6TI77XpLtZw8pKkJufuKLcIKPvuxyCfPinF
uC8ySCVfkdbHQgS+lQWXZDE161+0Z5Th998IhBjjat/zUo7RR6MwLzC9nQWC44LW
lRTvtS130qcrhTIkc0J829/HSgC6lBVU7Oe5dT0YUYDQoUJF9g4ZTwHpVN2akYqN
yAoIR4qhYEClL6ali6Eykd8Pb3Z4RjlAuUUq+INQDQozm4hY8qeN/c1yMl1BZf9J
3uT2CkXNsyp91NJvw43bFvb6p5aBXyFMnQTxEVKkU+9OpQk96lXyelW5J8hkLbGh
RZOB5M89sfcpFOsJAS8/iQJ9lR3m0AMM78WJLqrJE0SMcQ2R1u2gf//u+yeVfA2T
ovGlLc0b3hU691lJdyeJdFs81Re8xo1ShW4DxCspf6Db8lNqCLaFvgBRrSLyWmwG
7fP0q+CfyJby9a8l+77NcgtFE49TRmD7RT68adyY5by2/QBTrNsluBHSiQP4eQRy
sATAY8OjDAZEfNGJ+YuDkVLwE/lqzWEJg2Rn6QQv1CY8Sd0vstJZ6KIAgvuxbPHH
UCAAMUqj2+VtRy8gnGdE5CAV15RM8h1cCzYxB9aZosQM+dnya18t4lPNw0kWGmKK
j2gtHpSrTZBpi+tBRIeffuO00uzXTrEA87dPoV7ntWZ/8A5l6nMojLpUrTZtN7y8
uk8cLlqMK5LMUVCI9981GQ/zcJj9Ra4uBsKAQBvR8Ge5LhHSi+ci5sMOK8rr15bY
he3DSlw0ckft6PMQ//Qqe20dgKpEEGFaOvrD2Of6/KgI/KNGGji5McmKtqgInRw0
CumFsRFxNSkx1V4s17cXxFmiFBFySRMpkw40UrMgBhwz1L8FE3NHr0wqyEmnzyCu
SOpjsEgE4kO0QEpGfVFOW4ZvFSXXSAXDXTb+rPCKoiA6f3e1p6d2gNOpJQL7AZmg
kCTzLGgJHCVdg3gX1lXNkg6DcOJ5TgGCj6A7jNZkkRMnzpnjFliVEtx2UspuXhRD
yV8As1JCcCjMygmGfFb7tYh1UMGx5WQUis8D2U0koQeL8Mu03kl72pDd7qpTo4t3
hqyolyxTw/VPovAhWxSEtTpsj1HIciVADnKEmPUReHNtnrcU0U8tfJJKxOWkH8+8
Ig9iD+5YA54bjAnrGbuj4enBPIrCKvKT+KTJpOqBWklq2lWyRtR2UOa3KBl5MPlG
6ECPOJUpOzzNuyPxVqgCo4L/xgO2346XbUFFCC7lGYOQxVavlBcRjOKfUcVQCR+I
DxRT6ZloTQvmgl58z9fXkZx0zeatgDp1qB2DskVUw3GcX7SsXw9w/4wEwjMr+Rwa
qCI6QPz6tEaTOn9poBQkr1oKNzOnuxzxNlR+wPNihYLOvnLLUCab82vnzz0ksIfD
72GrUe9y4ZZGDWLjJoJZpgdrApVTEq+AAr4NITcTwYsS7QbTwSgea5QsLd+2M501
I5RkjxqUWM0+8GHzXeSpOGNEabFsI3H0olWsRRyAJwCxQ/xczb9y9S68BSyHspG1
AHm8ah5i86yFOOKBnFh2KFDdmsnb7PuGLUzILl9DLlGd5xTaU+VElhZfkp0Lfc6u
h0VlInr2isndrxkMwvdDv0ESh7wKLUzmjx/tSBbzofx/cp5Q+QcKHer25x6qMeBQ
L8KqfANjifhZyp6U0xHLgeSceb9YwLnUuG2KdXD4Kz6zPyPtDOS/k34Z3Ptzv7Eg
U6hHxJB4ZzI40McBl0COqawpjWkZNj01+QC+ZJgmltRVEgPHONQxVs8HUoEvQ8aw
hhH4EeXZoCGbKSVbvgarjM0Stqn5o9A+5aDFUF9wGh/vikDgt0+9JNlBpmijpUAg
YsVL7VcgKRwcMV5Xjfrpqq/ZNMRaUjR/xbmFxBkQFv7FNc6S5Ot4X4h/a0oUrTPT
pbsmhIBFaY2wzAa1pork1O9XwMxEWjON6Fx2m1XSQo8CefhA5BLXhTT+RcFx+lE1
oh4Q641b7djZvtW7tQ7KnYkqPfUHAwvllQ6PQ6Mm+GstQUGMW91b0llMcxhHLHzn
jHJXMDBTK0haHT8BU7qcFp4HL3vaucHQLH40Gy5edpe7hbWH49J1D2+rbwiOjk/Q
hbzlUmXFvRyK8rsNiWjue4xIfs/IO2sxjgGuRsJKRXEX72+pbNmWjDvPfac2WvSc
I9Xrqu3jEBAlRT3Bahey6EvJ4yVBKsijiZZExYbj7pk/xfRXMdDGbVssoFwcLd4s
KwV7wMVTs+vmOvwoMlGLMDEZTokn5ie7GeFs1qHsiy6ZZN3u/FenNSzyjFHx086/
/dcVr7F1u5U4gBvo4YTKmj8et4xx1UA2+Qd0rotwdlC/kqQLEFiGUHKnFU1QMl8H
m/Q/6NITb08P4I3/66jdGBj5ViesdNgFTBjnIQEUBO5cTOpk89+cOEcsybfMHR+0
SOpdkyTBsWj5QibtaI3FFJfQovPDp7/p4rBsMbs1DPMJ2wpQq2ZQUQ2/zgb9bFqI
97wy0lbQEeuVnHi/oihDn9hdxXZAlQi7TpTJEuUJPWD3IfithdafiitW2lf0hZQc
lnTuvNOLs26ATurzOt/PAPJ//JMo817Gzp6Fime0+c+SGowUt9QnCxRJWIApR5tF
c5EyUxROtHr/dGZDKReKb9GTRfHZ9ze7xOMj14L2PSLon9i3oP1fsh42XCwreFrZ
3+sHxmdqpV8Z0M0onBrnx1QPcJ8y50m3uhCdqeywIey/NI+q58Lu8+QlM/xJ/Oh1
olK5nWiN1XnhRT+GunVzqDspvhmW5subGDRpQtmmey7PScvXY4T2FlU2ZB9abpHb
NvltNkUclMHDMLjnxvmbofwHL3OlDp2ISYBHZs/s9XMf797siPcfLqhPrgJjAecN
Rz9T3UbBAtYfIG7RRyCwXF375JBb8dIQm6r2IQxNphTU7QoqSB32Wfhvzsnj+rp8
3K+XTLOivwbBLmzyc3CQzOQxTPYFZ5W4Vhs4fHElTeXuJTgFNPeP4CtiGkFV+Qjt
EtF/ydr744Oivr+7KZkZVwX2QPzzIlCQa9zjJI9AueucXQAXe2xdSj2hsQ11JhdJ
tU2fUe9qTbyrbX2ZUhyfiLmza9QEW9wekDAHLy9mILKVovON4ymUxz6NGPJC/BCw
fgI3S2jNO28VNu+q616uWreQlHeCUM+jZy4bPVdHy1mtMnTMHtgl9R8ZAy5KHwX5
pA2EHnrWgkBSv7ccnNKeEzS7HzmGcuywS9qZ0pVT6Qhzfb0gCsyqC6R5k0h8+QKO
D8Ubd3h9q0DtSyk1Jv4zQOvFDNKvr1qHgnS+vNFc2H2PgpH1LEQR4DwBTmoTaltY
/C5u0oCdaHLzg5o1tXXOHPuianFxRYgu+ojcuSZ35+mCjIeYQBlkqfCMeC9NMHfA
euCjRDjzHgk/2HmZkgH2hO/XQUw4eyMTFyPNDZz27E3256iqRiN8I3Hw7VRR1TuU
/A14HvZLLnN6LgT0Kylc4sgDc9OvD69OkkED8a2IQjnTMuVcUXaymUxyWCAv+qHl
liXfASv+fobtxYK9yp4NdlcyK1anI6NvyQG+uYiyjvOz/OayoNQZ1FlsJRM8QYF6
VvTxn2NXmFcNV2hKXPmdr2Ovbu6ITxEBhhfpw7A1BqXsE1uaqoI75zrkJqnCQxz4
s+2MM8EpRLm2hf97vRy717EJ6wSkWiQLOzdbcy0XbInTBBYv/DTslGcdiL0WUQeA
WGAIRpAHlwVDtGb0QSKIX2J9u+nl8Gj+d3N65YBb/7TUUUvstGpdTPPy+nahfdHh
row6rzMZ0pti6pcYH9oDJkt8E29aFJJvyG6/vmmJsainoqehRdHvCOw5bq1AskTT
+fA+L5ZU8LaOAQiVqCAmUdwMAyStSvEpi6Ch29eEgB9CjLN+rftPfAzwI3mS1GNC
ePe+hO/dE2Yr3NiypBKR+iyI9fjeqD8PlbE/gWt0CyvKG09zSytoz1aQsCAZ8sf5
8/KRDtc0NeScFavH3JGQ6gdgGvGMD1IH5vm2fN5jtFmPaPxxH238FZUMtBiyPT0H
TfRai6WJBUcRNJ2ojV1UJ8kwDNGGJ4PQjrQXuRqFYPK2ABm3Jf3J5em89+bYWk0N
0xTrZ2N+aFtCDftzmig055mMC2IYKhFkPx/1JdfUqKTdGGIPXW/dmSQue67ubrcZ
/nnGqqb4gNxV/WOTRESVO/feUou9PAOGwkBMuWYhPBcRAQXNoM5DjvyFi3fD7FHS
WuiacIWnbc+lWxTeIdSU7ioNXQ2iZIqffvyft4UtwD2clnPTiD+iC/MKTRvmULUY
yjv+UM3t7XoCUBq52P1GHl+edRuhuGFbdTZmc9F0zjwVGNGJB23qr4E+I/eJINwi
f6KKUJHPX5l/nZ0e2iqHf88ea/XnzsaDHKXQXJli0HFrmgAFfC93NzvTkgRqxANP
dprU42AdlCE5bNEee3Xl52Y7wAtif+XCrQk58s+1QSbc8dhlnFSgVsQaQNU8g/LO
b9i4VHkR/YymQaXdIQGOtvtBCPbAT73jIf6xn6bmifu2C99mSWkNPjwi/BrEWrV7
XBj36J1si7Z4EPn/Fofc8B5WPKtawJr3awRg2JFWiL/KYzDn9C0AS5lPpHe1euVn
3ehFyTVU37e6Puxx4vl3ibXsAPVoF8vhj7/f4t/p8odUKlChVhEF1PTc2IiDfmBg
+D+bZzi8w/+IDQgZ+nkkn9uHWdih+R3k5ZLgBNMnOBv2w7DT6Fq+CL5yOIH6Rm5Y
iKEG7Kz/drd/oAne6qtiLpmGRodkBmP55aTpq3Scj4RKlsNjgfBmy/1Rf7/H7Pzw
S88KjkASlGYcvIqxEeF6vfk97LTaBpC4NK6smyDet2VFNaJ6ycC0Q97BIE3/2B6k
jsL0K6bNbvkgo9OCxBPqID55WrxQbvWehLfWWjLfVYyXEUTxscCvp9wCgrXw1I2u
jxUKlQwW2KvB4TIgjUJO4IN9O4d23GXvmnM/k3GJCjWIEYmvhHm8PqyJ6i5azQ/s
+auiSvpyxZQs5eO9XyFHbHzSLjz0d9MPWAECG8r/os+8rUG7mhMBwLHuKJwY5hkj
yh7Gn/V0+tODyUArNgoRTgte8kNhh/KACCSqBWzyw2ILWnqSVW/u9oz4S3fizwrQ
ZkeEt/16vWcdfNJHwX574R9fAj2CTEnX1VEkLV+nVh81c9A/MeDsDO5mqSZVvfyr
lbvtMHA1gQPaNmAbxlUVJOYz3DdeFjJ2X6CmoeKhped/7iqWGWM2FR9HARUaxqPk
KTjOX0FXW2jfKNVzWcHabOq6Qz+TgGetCE1nVpvCDtbO2oB2Mq1Qwzm8B7/tfnMr
FjoGZziOH74IBqJaZrs9Nx2JPovfCVCN9daV/COSzXd/DsPoODX4X7Zx+7gVEjr8
FIUqtGkZiCw9i2UXCAQt77XBYAz6kciG8z1AutUfKHtyyPhkJSMOT07mcSHeQy6j
ZnHULwd4zLDMkxLWd/+3ifEkVc2HqCNA4laTNMq/4XMvc6xu2sEqaHM3daGLwmuk
GdUPiczTlLYkLk+i7MJ3dk4ELVNQ8oc0dwusTBsCpKskLhBkReTy4IfEgYqxDiSs
1fBNNhTmcIdrKB6fz8F8PTQ/bgCmgdU5RniRhLYZYbLl2mCdRzoEHsgusLzIJGfN
yAjpEM3YaLv85pM513RxsgbDxuXM1JzSbioLEr4YBbCUC2BtkLcwLr1uOCgisw1R
XkaVSZ/RD1nE3IqyQZ7Sc+7SnsouPdV4Of3nXj71Yf9obVA9JeOjx9PaFNQQ568U
s3z+VVxHxzOd7XD9qko9VPiZ2vo9aYg5NGRt5y6D+6SicsBqQTtXsjE+0/nYyeJS
Wd2mfmX3xm3rh5NJMl15gNojwilQtdD+Q7w76Q7WtFSpBRVkPh+wsBp2FW67IlFr
UfZhOnO8f52f1WXt22FW07/KijDGhRnLdgQNXGZYCvNghFnfmtVx1q6eO1Ih2LRC
f6XfJxal5XeXRdh7z0HJEFJV0ps6IxOMUW5qNwD14QgViiw/j3Utk4XZIEyiLrkQ
LezCk8yy1zI8+LQo/xj/kBWPW0qJ5kA/NLzy+ibd04dMcdsAweg0Lt7AYFj7fZBo
aq102n3S+i9p9gm+8oE4+4QRCIlc74cwAUJr7aLF3qjgSD4fmF3K0HieS8Swg+wu
SF7Ueke2gjMXgb7JJT7KdRzqC5FyafLO7CKb+7mJQ/Nd+YS+IZX8iWFMK0pxlHKM
7d0wOmvzrGpZQuG5WPehBCHCWdepshJuNYqZisns44Cqq+4DzSeBNx183YSZcLew
BzuenlKlRhzInb0hQNdqCtnUCZ1jk49J2VrZlz6plEkQfmIHrD3Qksi69Oqey0Ec
gk9VJMWPRi8VDxwWFCGqbvjkXzxwljdVF40M58IngfyHgrWhL/JlhJ7XC/AShzQF
U49YAbMDhMYa9v4ngSRiqbKbHdk1tr4eQwZj/tMjNB8FmumyIeTegdPjWDRAS9AR
xzbRcfo8X32btkFwOFM0iGtrdRVyNRChfJEOcx6YNgTwZV1NGeCydoMVqm+sGAgw
XPfCihUih3KPL5szoiDkjNRqQig1goheULh0atgNYapBBn40Dczln4NLWaUzOxJI
mB4VN7MTP4wWIquiUsPfBzi9s0HICy0SJ6DBbWcyTg2j7Mh4UCPgeWJKqrrKs/ye
XvT9Fq/HpYk/emY/86jod0qoekvwo91FofS9GbcgOKu4kOzCfQYVQglvhbYEhqj/
8ChdCrFEu7nbLm2B0e9uNuwWHMLhB9pxVqfKFXNMWtfxHwL2rbDNE6KkB64PUILN
d1kwzLFpSdJSCxk8IMVQHICkVKscDIS5+qOAE5UPJhnqw1EdoY9ICnP7TWTaAB9W
b2eRpHFx7nJCdqEnT/42JXV8imXC0GUyV8lC6ozE5FpMUVz8GUWe2GHxWpVzSDIU
1bHKFoU9mZaRqO5WmpvIODMiMnTAOni22ULakIUlDbyA0Mmq38si0ww67jg8u71g
FoGouoL67OkpZ0lwDNoE0CSPorvZzNQ/Olg2MiPZXaLUjbrvXKAqHjn3M1Pcc1GU
K6Gie0wx0xa9ehu+V3efXsBRjnaKQIpG7JJoAX52pIfYHpXlcLvov6+kawpI74G1
0FusBqNdaUH/ix3pdAtWZTgC0pAhcePhKT2WPMHHpwnV6kv9/8VvW9/mDKKQ4FHo
xkCB84N7+384Y9nwgkQ0+vdqDCIidoBxdTs4shm3N+MS7OhpUqxg7g5141nVED22
W74vTER3oB4wTg+XZeWyaRJC06nJrNhKKzFUGt+sfP1wu0YsdKy8/54C10xV1hDt
x7g28nR1vX0lsY7hLInux50mcvlJw6w89EFtKWQT/9ZTlQ6Vle5IYUdqCwtDhOhg
UqwA6gsD4OtFvKG0nwUJHu0ccBFGSEe7LBjdnOi6NTwaR3Kh5DyUlmVDnlDGGbn5
B5s4D8BuT2ydaA5LMoVffCwngA7SrnxPDUBfcj4VxEttPb9wzhmCUnKQrbAKFj+Q
nJ4yiyBhsh9qt9jFn3ReOb3LMS1spua3i+XWLn87rvntwso2YHrEwsCFqiDtS1MU
K7GduONiXtuPkXO72aQe4Dr4yW78ztVKE33R6u3mIC426/LQm3CFFbaCy/ePnkJM
z3RmobLoSnwflT/uScmN1+V8Od0+O2pn9QaPdnXzRAfxSLAxi3DUBA4xgoV+Utmx
yJowDjVoBfZxJJuUiG8QOewusSoFFVct2errzbDf4JxNKtjLHu8ee7WZnKYx0pk6
Cbc9OtXPrPX39ySg1Dq5SLxviIxIBLUl2cizm6cuNOFQYbKP2OXE8RcgG/5iu56Q
1J44BBeI2w75VIbPPERGaPqb93ZwcWelIRm+6bsAh52Ypga7vFV/0fUGP0wv/ubk
NHZYtHKNr2fuByY/RFhjMwzhjlUYcUlirVgYZyCrpCz4GtnP7BEHhS7Ion3p7IDd
OUHi/J98UC/IVahPzRp2OTIBwzeUfZeRkkwHIySpP6L4VkLEkJkI53hkNtj6O5rY
CvqvXcpigkC4WZxmhQGwaD+L0RVUbkIBWBW2pa39pFciuqx3H3futZ0X+rHMAIbU
R5W19a+EH7IMncdpWGnWRidEWSv/C1DnN/mvKWX26gQphurmNiJLHbN5dLJzd+Kc
dpAx/uNv9uSiFpsQMBIN1//vUv9CWFy4Z7ND3003S+kJEuYQGK0tZ97PzgL2xheX
rm890JuaUg7vF0MKX/2h6md3QistUYqHtxrMzC7WuMxVi9juZjGXagY52VOIz4JO
p5e7CLOfEjtqmKV5p7NoaRV01Gk2GiFSee+zhg08lKMt9Lu4pV96XL45ffGqLfb4
CvKtUp6x3Kb0C6hfu//jANG41IzI/B0Cy8Ti2U0cD5Np2VTYphYZcngyeoTr3Iij
q7yZx9QKQ83hBTODQygM4h4UCFEQ/1Xln8Cu50s1fU/kVNMlbUQ3Al0oRfxgGfpf
FMgOEfUg0elx3+vE6atY0RUZDRu5m0GTUHvSohE9Kf4/4cagm5F4U8gRj+Ee5ez9
4JM9llAfNP2wduu4yJeVzcqs2mQu1Lv1JzV+hd80nLymEBMPynzFMaGQaf0ChHs3
r6tKuJFvdtb52tZJgGS5j5KJcezQhDEgL+6k2niWtLIrd+QtkBysD/ulw/Gg2zqy
KLMTaX4dXzSPy+Rhhjrx4y/OfdFz7r0veyCzECvKDEzi6TVoCnP5RNUNBVF8YmzP
l5qATOdxF5XG6T1NM+MjpphOlY6Bug8R1LU6pwyQA7mSATk/G6nDxYvane/cJk+5
J88UNWqOEEwab/M8hdX2pLfhIx3iwa96jcj1sUKDulHJG+lGdsUeeVKabElt3PMl
BN10qkzbIVuqmkPwyROvWr1WdhSEypWMmkaWjyNt00ud8gcC+wIaeYrPhpC2EPJ8
dBLzhugOHR5Vx228nAWV+rPEQCjGLuDfAVCvOVBjblAGJkBHCUwh2HdQzPR02X2Y
S67/QZAPJ0KKa/F9ZZ0jTiIZ89iih0LtJ8Z8B95MdPYjt1zwU+7Cd9Wp/5MVxjP8
VN/d6C497M4bgz2vqjFrmcdjnZUwPWy2rP7WtoWEU9mVgzk+iUcuBYpL8hjEsf1N
FEtO8pqxPr3PI6yKF2AEFgWBlX3W70wAHoCX8NEDvRljTvY6MuhduPESw+qrEjdx
HAQJx/2+LifO+tL7eoY7+xlQFTrSt8JryV54pGPisUfAmVtf43lXGrs+fcf8hQWE
zIoNkNAdQTWiwvx/MylJPnzbQgV+C7ACqRz56jJ3JRuGb6sZkOA3YobNgVBlXiT6
rfUf2cU8gi5fSnFIP4q02H1d9jDtpWHyZV37Vcm9/IYdRYytDtHqlG9AO/NTOqcq
FepxC0TfsD7uFiD+wBAvD9gtXdBL5or8wabTVYgrvs30oYQrTb0t0gE8R6tQM1J6
zbmwcs6S8xYKemNz88HXHGPDuBYjAS3+J2x8GdHSmwxwxJagLUoy2na/HzQb5jPs
gTCFdXPyU9Exmq1gIq/NEABE3Nz8sLA8oRhRJx6suyjSVjm5AbO923ELZ2fKIlSX
4O2yO790xO7Aehk21YrR4TvNFI/aENDbEr9yghqe4lzLiXHed0xbP2ZmrZZzOH7p
HS0jz5G9y3bz6olItCE00QCjQmRq5vzHuXDlbLy2j8W8bgDLsRV+Ci2GoQGPiKcT
FH7oWnUIt61DEs1OrgOaxidxVC68mmF+hH+UQHrI8V97+Gc+OO7d1iNzRGx2PT1X
hpxAHyPljwK/IhVsNx1c9vSVb1/jmCb+3X7JDZIVauvk/i5DM9r9ZOtKpXHqBRwn
yI27icSk9Jfpr19dSbSnIzeGtw7qkfKZd5jZ+mJspG5NQZrQCl1ZqEfz7WYsq7Ml
j7zzqCSCZtUMSFno9vHQLfaoSd+GxUdW9m8777z0zo6DLaPPCw2VDyW1dIzxw+4M
3j1Mo5BC2Gl2hfAwjje7cQmCeh759Sm40klXNoz+Uilo3fOnDZhP/vkgCS6+byQB
GOH6firTi24TA66GfqWhKyWBqKgcDl959WRR4EMfCjeXlyYfLK8uWiTRePiRCt96
EyXvW+IclGbmhu4/zf1IDPMqUBPN9AYEQzx687x5FggKcy1NxFUT2Jcz0OLTzOud
4oXZ/DYib+XQq+xOqUtSHQb2l7q9gGT0h/nh9qBl+XIRFbJ6CiJIGdpbUhE+AvoV
zx28KuOIijBcdbv7cH4HByV+SoCsb1zjPIvIfOTfsOJhM09s/OjXpHbv+8mKV2QV
iQB8WUy5Yo/MsGJ5SREhzu1FnLI+zh3XGhdVbgQAJyKuy/o+kjm5Jb9re+PfGr+9
GiaGob+MODcT1CId/TlwhkmN/hiNLQ61BNgBEv8fLjbFymaVYS/Czo0vu3/ZjjUP
PSoQqEG947esiO6rWR/YkwRG8nPN25ItXMM2DtBHv31DuDEoU7s/T+FPB3lwg09x
Rt10E6frkL+iBpsC3MMRJq16//+zfMFZWMhIPsK0dk0S1kF2WmaQTfjG2q37orXk
TooIyUFdYEq17XiO5wAWvep52YXLu77TybzYFH1fkTPEQ36TaFiXo6S+HvSytwVn
NYPU1IDjuIqJ23w8ydOAKloGUqgFINI75rbqsrPEG1sWm/UmzsoeTjz5oQClGxF2
sHKi20IH+Rz0FRtob/2XP0QlGjpF97Y+1qanmQXD8jAQ6B/bWKrKqN1BY6jzR0Yf
+OgdouDEmRntaojBMoHb00qfyOPo3Qw0HTaBmMTxdSj5OJmO+zcxKzEwP9AVnxZQ
d7psAQWumXrp0w52RbFeAACEFzv+3yeH2EhTTdT50a8COUR0A8uDcGyIBrBNj8zw
hIZ/LX2n3cbleHw39IKaZidU+UOaBId9JkclgTYwVSAcwnuiqsBbv5b8McSl8gJ0
G0Ier8ittsRjCfScYbZhc6EC+wsHkXxj2SbXwy/kpu9OhY+aJ1Gyjg7QawOP9PnP
FS0nCZdh0AMRvgIVVXWF2CKa2Pwe8YNeI2j1sa4ZxD5HuaID8w6YYdt3UPQMgaNE
L1hS4rur+7I+VU6GWHGIBZyLHgLb1rI9qjXwILYqUDimsyaLiw1uCuVYj/MahG7C
2H8diiFQ3HduKy8DTIQ/xvL98KvFdBfSV2FNe5wU1uZE+GPPq4mMe5tV0rFmuVZR
Ex4YtRc2EHxEK6GZyTI124LJxet5q7n3tIVn9oIY59rZW+RbBgex/PFa/y17A2Lt
S2jSM1PuNkUSq53Xzc5ZdrVTELTKIYq0RVVWUZki2F9NAxgIMm86GkQ/g9qz63jQ
9OBJUYMC3HN8HY+hkNf4eGWpOUqBs/58DwjhhW3MYxpepBiyDtA/9um/i3NqKPZv
KwWe2dBtuFimD3VjIa2DBqh0NcjXvhFZnqeuBqQv3yOV7C884OtQZUP+fj4ktDnF
WK+PYitUtKjemB2fhV5xx34nwrqm/zmArS86gZT9Nn7cLizl+CGKq1fIeRIJkUIN
e2BKWutVgK0vIgj4v6CsxgLAXKP+cZVoQNrIiZ8PALTst4Yhj2Y3S6QhA+3koAWd
ay/hppZW5WxE1OsC+E1G4nt24egrlhKCxvFgfPScVGRK3pLLd8LfoLzqBz07sg9f
rQ6OfvSAvutpZQhO0uOkLm+iyxC+PsvsIbEwYbh0ghVnSTFMaeUKFWG5oUF4Yk92
rauxPeFBVW5BPb4VSuywbbTvl4x9eAlREQG1MbadtZADtCYE8T1qiH4mm5R9Y61Q
tiUwiPIdqNaxzIhajRXLyD8RjC1p00uoFcWNJ7+b96AbFg92x4dtmrixzu49fYsB
RyIzXxEIXLtyppdZWmy7lOEqIDDZ54gRj43so/jdgxJBy+X6NLSXxUD2x0VfGwPj
GEo/N/uMX0MVD8JUUHb7lHsnjGZ2a4eQezPmDA4h+WUNflotc18EREi2gVJ4Xbkh
cXLomZCg1QwOgbTt3mGvt2FxeEOxVMrIVyesBTYeYeNIocVQiIUUO2ZPtVFEpqf/
WVi5f7AHP1tg+LDDJVBADAwgSTYG0ywy/3mSdyhRBMOsIsbPIY7gNGALWyz1k2e5
+qbJNwMeQFTZoCEVWonL5QhGsARHepPfqSRr/LOzX/zVVSICb0FzkK8uUq1o+BUl
3JV7nRJeXoMJtOCo2pZrKKNHmReVrdI7tlTa1ODNYEV8pPLunA92J2G6u29Yn7CZ
E1ArHttSF88i3e08EQs95RbSv8hJCngtG8q9qraa9BzXNqBkHoxD1JVrZrWESjwi
4lCrl7hrW5cqsO46eR7T6UcRVzRLaLmvdDY32AK9tTgr+bnmVLhHEN/PYO9FShzB
JYRQBlkGI9ms0nPv6Vhcy5wWamGfGUpg3n/L2EuTeva+sXInkjyO74YjccfruaWe
ATBboS7tnfOEctUC/EhGyRMGL/CKtA7xUBFBqbS3qXs9yxhWjmPgKWf8tFMswhhw
x6WO5+W/aBi2ui4uq8OCSPHfuFLjH7dEb4KCe/TczDMOXtsHAsIYLz1R0eKJG71U
g2gmQafnzviWWLHJ9U35UdX5m3X4n+uRCCBEJZkG6sxoWpIDqLNg8KoNr0MWpeK8
KlY10jB2/y/i8veW4ykBimXlJRsuH8CjW7/qYD37opjbpBYk1zrN+/Z6dYzIZzxa
ryGpnJoKpglfTnWSEhnUC8Wyfh4In2VnhsppiJrBjpNOGCnj7v58l7EnTEteht31
NTezw837ceQj+o+ggOvG8OilajyNtSu1EU+CS5seBsU/4svlzbaBPeoCBoZsztgP
WtmSnCkDDr+jwKe0TAQIrAJvyulvZE4etmMlnoMVdk4ll8OreOvJKAhezBFW4o5g
4a/gXXPJN/FpCV6caMjP0wSpC7QPi5fFwvOL5PmsOL1WhCroT+zmbbWU/VRSHsgx
9YTSLGB2AvJL9xZnf+wy/vxIFZKLFUFUGig1L4zBLgXYqthcmTs+FTfjH3h5iBYm
RN0Xn/ir9GRJoR+iI9S8lCLfTEE9o/kCaJy55c/aiHjCmtbvovRXVqeVUFpOHcYT
8Ynv2rbIMz39fdcXsJAK/UOv4nmWxbHT+Wq8+BVi7thaOQq2ws+sI8SNR+dT12Wg
Ug8ny2pQPOsrDmRUsFj+DNuqf6LeU0uOy+nu1//1a3AoekHGCZRCK3glgz5YOiWW
cSB1gNt8Wv+f9kaVKQqFP5SDTGYv+1JwCy143p/geNAE4fof4ltdxrCXeV3zqMXh
l67Td/80nQl5sF4JvItR2cijctfQ+6FIB8iNHRXHdFsBDert40Qk1pE4dKhkwscV
DZgHmWWiFE8ZOty8XIgeYTS5z/lhwWtz0nSQFch+PtpI9xMTqSapm4UEjRcWFCvI
HKUWkbpZuG/6pezHvjMSDMdcaQ5ebDNK3aV5dOkYPRyfyv57cQzfUq8APqWwiwNx
Jjp2eOGFqVrnxDF3+y0WYltEVI4QDB7x7OMKwjDRucslUQaTN7bLoJ1ewPYRAlYk
tUXeaX2vMvgpbXFXUYR2PxG53UHuAL7p1ImxjWRLyuClUr8/VuXNU0diETfk4CYR
3A/nCfu+ZXtxfhOJdhqMKEj1oYjhfANxrxXeRYUGqDr07hJC0JxO6/NN4TYOIenb
elkRSV/KuIj/YAfTboPHDUGp8Z3igQsxZVKaAE34/pCnCF/wEEaVL7LARB7Hw7bt
6fzPMB39V1kQCadb5JNZYJQfnLfve13Dk8lOT4B0Pu+i2mvuwRLcTnpmejTTMjCi
UntG5Gi83Xz0SWQVjHQvAvKpB1ETVbS2qUbyP0qV41oeSTGVtmqUZHUzhAylfGOT
W9Fkj0zCHMR0AgKm1vMh5VgB92RV7CbLaau3c6iWQV2lejgHS6zysAp2tlRzPGCR
TGkU/IYBt3ZFUV3Ra3w4UPv7iBlXRgE5aEO75e7HAffKwSkQv9qcnFtX/Vc1hgsn
OCrPjAGBUd9a4zPk0oO6kzibgGUj63kk3b8KW0zVGvFGGFIphoNjJI2toAVEo8DV
pYta+xR5EkY/vhDV5c6vLhRpKljPKoPryPqx3lP0i2133FeBJ06y8lJWqctJYakk
ZcBrtehm6FpJyPXKidB7xDhYVoV4IzZbpfOO0kZz62xVRdRRxFqmKU7Q8gAcrg4k
NXiW3B08SuUOwAEbhSc3cvhK+7/l10jKNsKbwKac6lqGkuL8YUVIIZZU6tw0xsZ+
mzMwtxA4pm91RgZnCb/GjoWeAaV6vqNAR5+BeRO327qw6+q0VzEbK3Tt/7hjTcye
ovhMonreNew+q7KdbBSalSi9yFN4UzOFvNzBA0aVivNEGPEsPTLBecWbs7CN5GtT
4acwD4vkw9fHvzVYROrMiFfDGeNvMk/o8bWGDJhI8XouZc/wHtXq5Xjgdu54qxzB
sTLSyg58JHLzd0jC6p/zHpt6hqgYIk0Mjc+szrmWP6HI9nLMGYizr66Z6Q5cPzC2
/2jV7k0uYIbeKKv9emSYCYZ58cUKhfsuiIm8Aj5wv9CrF9s7bEUblsgYpYCMFi+p
xE5HX23AmLzSaO0v/Lxnutu8FNjzknLMF1hboQ6/UKY0tPfEyB2N9c0gKt/QdSHz
I2toDb+t0RdI/CU4Qrx+wELyRvrUI/PPvZPu2RCC4idAm+Pk42W0pIEGtNNaj0fZ
7lt89U9YoYmc8+E3k22jUXRmX7MYgXJm74XmpBRcPiVgQbKwAckRhhrQMqNyS9s3
Q7TFXdHmED2gltXevSK0WZcirhplCXwUvnD7ak3Hu9kyHCfSdPfiD3EAw5+004j3
tzKqEE9+fXkhroGuiW4ss9g5SCe2SnXJFiLXMdKjzW6Ne/NqNT2NBh+VNYJtwMnE
2c97PHThJaEg9LQYptkILzGPsKpPiI7va8/4nxs4hQP6kXGIhr3QtD46AbP65Dz3
QxNGOZjfIcF4h4N51QABU51K5cNTTQLTSZU7wiMWucMkrn7cSPp+zpUR/WRiGOdf
4xgLV+YvtkjxfmgxoRWkJvAwPPNI0BNtiCP8gIXRNuNzdeHhY5N0vp4H2JCxmpRR
Go9hPWRhMI6US5OGVPriLvchHSBFIiROljpbGcr5JuVAilpRu09lNNv/zE7aE3wz
XCJCaAo+Iy/ZdtRn2smHoENa2Rg+AyHPphdFMuriS8a0a4TVx8SvnWVqy//QBGT+
TgIFJ3tdgtOk7FR260c7jsm9xmLrD3yjVmh3Y05h2ZTtxFNunZDmmcksm5kU0TT5
2jCgylU3Btfd9h6Ba4j6J42A04iSSXVvzR+u+izK5soWlqDPMOFMC5V/Cj1Q0+2I
UusJkwRzaePhF5/xRKScOsxtnIeRtroSx5JDm/ZKYIbpu4Ix3Jyti0RP6jP+D5Z2
VgAQlkxNG77YUFBHG9zoaIhNcC85Hd8qAosrbXlO5/N51YubG2jbvbZSs6uSH8o9
RMwLE8AmLn+LQLCdVpnEn1wq8csfJOMPCMvPL2q1r8mTWsn6G6mXS5PwPcpU4Vxn
/mFXV3KVvJQcpvRr8JfvJa5+3p7qovCDMHIl5uBC3FAWOYTvHAc5y8jGxeotblZA
QjEas6V5XF6LtK7/Vitn/XkoZGvXp4bVXSwxgSyUioMI63Fy+4NmLqmxbuE+m3Js
Suxb3pY5dzkzKMgkt/fbXHO/9vsmGZ7SIWXMA+BMr03NWLHwQkIt3hcRs1wU5Q9o
+8o544ZFQS955CUEQ6JvqoVVR0chrkehn+8a1vcsGmD4d6U8Ejcy3gM+VBX8SGCy
uW8qPxLXzFdGthqFHzlKQ8HAODmLQbC4G5acMRf30wo+5qW+wAbVlA74V+lZdEew
oZkFLL3aH4SaCGDJb0PKpwly+NRsz0MWB+lKKUwPSLXanjfkRKWCHD7rG0LJaZwX
/LMjJDm+j2HzjYJ5mSPeUkVLJ3cOwWNmvgQK45tWprCJD0HWpco2k5P0lCm0PDka
YKooOXmmtyLqrH1wuey5cm/UQPdqqRKajrqo74gG84omlABWrocs61FErPfuEmJW
rHypC6ND059tQ2Vp/7DSV1LEo2RZ+x1+XAaXNS88U6I91711YpEWFpCGdJX6Wm8L
5AQHmSE2zrG9K0+1d3NhDZj7OBQlCD2LR6ImDe5Lec9DucKcT5lnr89WhomzT0YS
QshbYI8agYQrVlaKAoKY+qAabcblm3JISVrb15vbb/ibtknmAVCn+UkJLbwVLpqq
mqdnM++fe1xDm5ddzpwwjjARW07DKjT4XkJaWcKf3YDsOG3B/lvfr5AgU6o/ieXB
l4cM6q6VHYO9LPE2d74M6+Y2qKRGtPFJAaoUP9WNiWe6oRoIbHq+I5EpNDKtikFX
qavQGeeJawf+NcWp8UbL4crNT/unDkOiRmLXchMInjm5v+O4vKA8PkuQ275aNBx3
7a9kie1YGu02rfeyUYRPJc/D/afGjIsVxE0M+5yXz/8yxyXtNvP54fVPo4QXQoAY
1sKI78o3MzemEtgD1rk0AqKcqbgE7bssN3HhkWBTaKfPgEl6oKEcQpF8mFgp9mDk
TzZdP17eZCPczFim3/Y0rVCO7g5GXJq2OMTHrYCz6+C+B+M9AN4WzxAjonkendcT
UQXlUFKGsEHLNP1CPo7eJgCXRjvuiZIb/UOyASR7JnMHDsKIcST2kvSm/EkgJlpO
aQuLC54igWNFdLrJsRs5vv+TNWefaUZSJHOtMuO+PDgels7+x/uEbXCM8eO+CwXj
Phl2+3e9sidX+VsjI282lmEkuC50V9RQPBHoJLg6Nc4yN6odAIE3UgWIP0qVcqgk
vd2vbjU/pS13bF5VP0j2ba11eVXP8XVPWWcezMUk8s0ppkNFbOsM4bklRTD0Lp+g
lLU2jA7QLnngoTjgKdcAyN4xBlBTobLdLtsWM65vsSUwAvYv+fEL73bXQB9rYVWI
MHETeu9P6vJ0d9aqVhFeFCFKw0QRSsdCAbWiBRRxPEmLktOvzIsEBQzH8uvYDtIS
`protect END_PROTECTED
