`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqdCB8C1G9K6j6vhYht3eJj2aUOYwAzAK+BZTB3Oa8LIoltbaWwLalxpCldwTMG+
5CgEqcs+8E9Oo7Q4KA1VyyJQ7wXSPmzF7k9blMUgiUBDqq041Avw76TTjrBg0VvM
POhzhlzL2bODRNhVnC/NNM4PoiOqTUxKdUUEKAQrnjcHWPVH1wcc0/LnBfw9sd5/
WLC5wWDDKZCtCxER4ZRdM8mewqpE390VW25RrhRdL32ZQTFYgxmuuDb3jBBKwiqg
Axf88s+T7q7Fro2gurFK4k+9B8rTkpL2WaYEFGrSimg6U7PraagBVvVqBkv8U0aH
fHEIrV9f21tujcucxQGn9IDXBdxM2tmFeEtfzBFso1wNbM62ylcIrCEsuaEE4Ggt
kr1bkp9iK1nQi/pVmxVgvqEg76Wid6O48AnwXzZokqGKaMQnXvS9p3kA3p1nc4Nw
Hrl5EHQ1JUpdTBMrhD7DG8TsK+M9D1sa2ZGWko25ZHDXbmiAhni3h+FRu+DP8FPi
NLp+qKK9FCzoCCsLUvxVC8rIuS/IH33peNam4uqjQesDaC6R9YYi1xjFhf61kCEt
fx4NWq5o8yABLJvy4xRY+VZrFZcLgl8uBX1bC8eiFfPvhT2ccD1I0qD82T+48PHH
3sHJCgARVRiuZ1gn7gNwpCL2kxXETap3Gkrb6W/rM3+hqK966b0c4JN42vHgqOwM
ZKbhUOTueM9I+FTEhIPrBKdtV4/AIas1ZNABGR1bWUJ6/BK9/r8bjoK/evSJEPjn
EUiouOGHz+vnDF0v2eLZN3pGth9PxdYQP8wtZSE2RUK3R8+9H1IHzzmjMuDESvFl
RxAALUnS8QN4eXOpyGZ20DVL3D73I33yYlhqHfgndB+CXx9+cYjYZyxxR2KOjB57
mU3qguuFFOXk/zuVZVxJaaqd993+4QdVS7adr9QeT3KGkQyOVZEjZ5WdSPj39hjM
+4A7MhNVPbqhM4ntuw59UIGMR6LAp6RdDAfvNuOFbHnOqmM0pbWr907Egt6EcQ2w
XUw9edmTEn728dq8p64U1MVqkwkDPkQscBj8M1HIf0o=
`protect END_PROTECTED
