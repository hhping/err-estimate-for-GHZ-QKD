`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KT+OMtItePerftDYoiE+TsLB7OaDHFi3Eh7xrEkLRGtN4Q4Z9EC0I6jlKJxqpdTc
beqMSqNENKIWc0jRI+qeJmO3FeWUf0+LgDQc4S3U0FhVGUIdceW27MF0b3xfRy8P
aJcflWBpqJfLl6Wf2FHFEfGo/FezgGoOp10u494FW6x0c7ti7FxuhUKXRv+ipzUR
LvfJstcQJ/uRGBDGc+bSqNLD1RFCDx+hF6uCwakT7UnWUvMDL7Pag1ry3DGKKq0t
oe/IW2FwicrSuOdjBsHD5w4mNMZ4JQVVJPn4y4US1ODWTPKIh92i1ijlLzTYg+jR
vi6xFvsJFrbeL7+tbZ5S0ALhLZ5FfRgZQj1DY17s6m/zQZPDmqBDycNv5EMTRN7r
R5NZGorDbuvLRJpvhk8J+mNNa7xBBAaOjUQVmqCM8xRin7kMlmf1ee4FtdifDf1M
S4yCMxSbD04Q4chkjyZMQOyrXVjUt8WVUFG/kO2clwRvk1RB02ndyVPnKRkZ1J7K
mtB2fwFOBHmX0r7QJWCASbdCi8j1hrvhTsKN7UP7OlekNQNuYBp2R5COBNruoemN
gUNCqiGiyhJLPe0ncyqe/Mm7isI41lTYa3lBTbLsy81wLtMHc7CfZJQx7845d8jZ
Oqz8vMaCTyNK95KuN+A2jLQ4kdRyqYLBXxAYTNyOB5yuSzuFAGVv4jaCyzbXvJjC
6AuL4p971H4qjuupC1tIDvZOQTb7jUrqPvfkCKqTKjQ3vDSko45vQdN9PhUJIdBw
ZCofmmKcXIJIhLAs+Zq7AX7HsCUaMDeAI4XZSh90RUglA9qjgm/DnmRVI8XNs7Px
xLtunuA3Iw2+uny4oTD5G//m2t2wJIglwSLqIUsShCmfm4MK1RgpRSKsjjNeZwLu
vHN7I6yWXU7oCovXFUzA2HwgixnivoeJ6AGRZixw9gNR+pe3w/NHXjxsahXiCOhE
Wsh0x2YKAEsDNW1zVphOQXy0FesNAA1i0al1V069R3+Aaf+cd1g49IiS3BIbH8bA
p/7lzP2IRam+75BHcsiBe3iC9d1rFTHft8dbBsXm5RaNnyvmo9utbfIFuRT+bBMd
9VIZH1b4E7NrZlf93ZPWsfPiwImI6AUrNNo35X9VC/NyE6yh5CoSW7cOKNhRengo
mqbnfXJGsUyNxxuMLRsurDlEQHHQFX3VIBRl16GNi43ggXbfFjYKGD+paJDT/v2r
icVLNmyMSe5ey64oM7PX7IDAu6r/DrM1KXDgRV9JzNy6nJSyjvJ/ZdJGYL/Zlru9
nKQHmKGQ4KiL5ld/9JKTYrF2hY8usSX2m7cJZbVjNyBh04MOd+X6lbtVNFS2rL0N
Dcv2vE58Xm3UtEirepenPjWVeHxjEnLYifM6Upok8xNMM4kzAxsQGZ3AX9hf6qFH
f/5T6//7BKIDSm7STRAb23EVQxebmirJ52otrhYbF0LYeoFwO2C6V0kNKbfzP383
Otf+qwNdkRjxeRxKQGUE5KMw4pXKc4FkXRE69fTt4PAMMgxnb9aG2oudeRnDhWyy
gXedjO+e+XTBCSUCSQkbcI/AerbF9qO/+mJeXWVvik9FYu3Vyeu6VjbINuq2LUZF
gWXpJzlXH05IDpM7wui3rKBeS2j2CRNN/yAWmgjG7DPR87TZodb5JJNnWf7B56qU
atK0b6eidgpfrFmo2I6X4ioNohRDMBWb/isBGE02G9W9l+n6+X9HGP6vOq8y1baL
HM+YstVoIl0XFboz0rFwYQwOPagU+f8lu2a1KWYLwgFxw9T0yLnuRnTM/59RjagI
QBOlrW9KHXI20p/H3CWR9MuS7tDdP/1MT8AJ5enFQE4iU8GFaGGYhGhlNLzvQbSq
IzMgA+A3ZUPGUTHUX8Hf1DIAPZKj2Bx1a+CluIF+Ovn7iZ+Fk3D883W5YE4aHhcx
BwAmWLnYgW457fZXhraCuaoVSZzyJ9xt5rwDd7x8/3rDiM4TIIgJQ4ELgPrBPBrK
9rbxUxOxuv5X/qPgdbiE0N6GxoUBNc0knNk1C7dH3V6WfwZYFH98zdIZpdHyCGwg
jr8oVpk/5nt81yj8ij9S5F5IPbcCTGkLY8C06mL8AB6K3oPtEf/W+UhErGx/qDrE
lufRvAQCVEDkmnPOn79VQ7rnm6LrTspVk6t5mmKKBHRlNRowa3rekuBOjhFjneE6
VU2O7fNdl+wUmKwM3yYzBGjPdPc9I2narYjWOuiAsfY2REkK+jP3l0PZMjOzYYRV
fHGRyfQWr5lxsVQya30oiM+KB/3f5TPuaHuCAFxViLR1CVjI1SfxKWHAAMbv/FUs
ouk79N1UU3RAKKFmlagf0ftQkwut4h3L3JyCubHkxmnfSbC412vHWwYl9h2Z1Zqa
m2bWSrlSQ9qGBMFokK+JjJMZhwS2w45khCknRu+axpm/HCMifxgAJ4et9Su41yJA
/SOH/n62BJAitXQAKGmj1GirnXVMk3q5NhAUDTe5K3zYqXszEPkBK6GBEZJW+Bzo
vGx2HyIpPsDqLGZuCm5IcEPHFABTPSG82rZBEuxtdbeoA8C77JHKBzKbVo5hFAP4
EdwNkzOfH1b7xs4H9Ugdq63M//mFY8yQO8THlX+FGAbn8tGcNAj3FxI+B938HD3h
bs3flZtidRHrghB3CZQa0nMXvlSg70HpgMlm0+otNi2zFL5tAuja6Of013Xpx8Vu
Guf/9eBD6aY+qiEvwhW/G6Dtqe1eUOS8YzkfRuhkgFroHxtvi+Qme6xyUatfBfzw
UMp13BZks6sMRd4m5S/4P30wJggiKkaBmLds1cH2D/FWL7FdsuaLD6v8mrSDuRoh
/1vk1bMl8nxaQ9PlXlV0RjtZ32cr0qZfs+8PSqHuz+CHyHIT2AjsOz0VHujGw0TH
tZoOOHlWg31OL1B3FCRMS6BncKy5WgQfwUidOiQJo/Svakrwl7OTIc5nggQ6wkng
ja1maMce2qcnOjfMcaoAZ/aVB4rcs2S2k8JtNhfRj5JNh+B5KcjzrQq8hv92oWZM
iAtcQbTHbCWIPuLVjxblR04lXa1Ys0LY+Fuo/kwZ9LZNmwZQXmjip6ukHO+e0Wqd
8Yplb7ynh5Hm1pYoD6yvPMplRBlcrqjopE4mZSDAswnUa1PLtCV8ktdlcqC6tQ8g
xeFdXgpOyHOWiVg1tPIyDvf+db0BFO2YrOUrhSBcc9x3FxWr0ImnRwEgMixkrcfu
A6mmEOF1QnHria9p0pX2viGzJ6S9wgyy7HY5PysmLneT5m63z82FNv0nkz8I2R3c
TOmtgJXKoOR2xpZceOeL1wsxY43sHNwWrRc4DSZg5TJQvoKqiMBuEFYSW2Ndo54v
MQH7JXk+ypPvUW63S8JMj/PDVT2qXALMvvYW0CQdEIc7dWU8qy1T8uVkyae4zQeO
8zG0GHsDC+b/gRAsUgS/Eq4f+lcY/OMotpqcTjZbpTCFOSfqz0GOtlqM2Wc8n43A
cWhXrMAkho/qp0SfTul5UyAic1r3WEAd68WMksu8CxvFOc9VmR+8WOsU9PnkESm8
x1emObKRvE5zp8wN88AEmWl3BKwQvWcma2oIMQwfaKDgjey87JlNYCrCk5eghP7P
ppW1Acj4c0p6yHvOhsKopIn5quvq4bV/Ni3/EmsYYRXZCNTCb4tkOWAuF+EnHeeE
+9BFJxJfHqKTbj1nmkbb+EwJPs7jKB0cBaiRx2+74ioYSUDy2pymkLbkHFqW+CYe
AuQTHEet88cZhZyyuvvfNewHeAo4SunN+11RBXRawFaOkMWkjRRy/X8slFdNWRPo
ly3+G5ijECufq1FNwX1bEeyJ7EUUjjKojCpr7tjw5zgAfXsCpYqaGdldpMp83pZA
pSEflGnKzqRwXYBNCHwPB949U6qkPxAoEtEtd2ykMhNRv2Iff7I7RWguu5UlfJCG
f7lxNZ8/iKfl1w3tmtkIex1fhJ0pKMEW89GYpxyY1woG1K1n/y4Dyo9NDeMXuvgY
XNwtdT2gw3ZaLsSIMDBndcEo3OlHXg+pOa1/88gd+CRJfIuG8qF+LPShb45vRJzo
0QXcXo+lrZqWR432dJ3/hGSGnZhJOOzQuTjywgSZNRe6RHRYFvr1/CSCX5kQX84x
zXFphZo08BlI0GiYTbGas5c/5xvNdb90OCn5IGqXVu47lLLoFNUyLwDNSDUHwa6S
VKv/rRI6qApI6y8e4CK+8x7jAsNzW7xjSZSbYwVfzj4=
`protect END_PROTECTED
