`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3ubddAP5j34UKLWyJrCh5qW3MZUFCyAwrPLWI4u0y8zNn/5veY+rMXvtzbsA2hH
ayplw2jgauo/UcdVqmcw5OF3SBr8aDaad29PQx3WbY/MHbWDOqLlVzfu0+tIFkki
gtrK6A8wntDWcwSAb7Q3Q89Mkhaea4DiySlQuCD27wEAp2LkRRWIF5lwl0z3vmBk
kUEnlVlfGOMYSyQz+kNUh/AzfFHiqf9Et6g5JVYVHRh1Kd5+sTIjunNm66K7dK2o
kCAr/1n22aCLPHN7/ixWGCRqTfxdVo2jGpbAGGMcz8il/h06iP4bWFER6YzYe9mh
F1P3PlJuED4y30QkXNho5I/9Pnd5Kn5iDPwySZb+YFrwgNkt4X7P89hz/ebtzYun
dImXk7LTDYnrBMBpc5bQVuwe/8Tu3VokyUN1kaXxb1UjeQ6CdxWvqgEtClnvTkk0
9dstPiAE6TZU2D16YZmK6oLJZVWF9tBaSO1KlT5SIhP+XvOsRTnrQzC/uS4hTxUJ
0RbMhTZIMh9XUKOBkAGDoG3VeU5LNayX5U2WMrKFx3b5iB0KFm+3n2kvDqMERWdW
9jNEYhh2xqp8F7Xufx7PE1swDG4OCEwBb4HOxZSZr+1TLhAaeqQEOzYBdPeaJFAw
GfZ41N1qrppmXkplAQkbcaO2ta/crYEJvJiHCFfu0Fx9mhglHTaPz42P6oYI+ZDe
HpLJAWlTUFxbhHXhpw0DdQp9nd8TZARpjtD8y4K8OJlr8KJEENSeUjompSsIxBu2
9S+wV4uAfey603yr/WlyQaID7cfmYYJvuc5h95kksvUbRdhqvlWAAW2X7ZrhT1Sw
OMFgZ2Vdz1WhJC090fNLBbsE69iVivkeF5zKZ3fELSBiZemaYItQsTuRrhr3kOu7
l7AOiQajN+xk27yuaZpv169WYw234ISbKuHLw2OzomSF837bgF1Ib2U6Cy2s0SIS
X1HXbYKwQtrxVXUGnlQ3aBXmByLhO5zj9AL5gb2yArp1dfdY1Nq13bV4HxoD2Q9K
CNASiZRZK+sxPeA6E5L6puG2DYcntprmT64H41h0O4y5gdT2Gpvc2Ifptbf4G+Mc
yLS94gZS3Itp2Jnu6P9puTnZYVAgsUe/Y0pQkIj9RyBqfJMOKegr92sdvbKBmEDX
9msQKRthQ0HDBfH75MbN94iP4NUcpIYj9vX24FRgsIhESrXKUf9AJkgAxd10QgPW
dRhmd3FVFdAzSPBVhEDuCHCh1JjxHU9OiefL8RaZ6dPcureblKWOLM0kaLylP4Cn
zmxCyLfIO84aQunX7yEI1XOuS8Hb4erm0/EN/sibh6t7iIKmfLIjmrp3uR/bPR2J
lKtCtff2tKAgChyNyGqoU/pDcm3VeUjd1yRJaRR58JLGSQ6VISLXxRcotBe2VL9M
j6Z8qyyshg2jXjf/Lte+xLW1l1YQx/JAVY3uc8tGJ5+leNvkvXNDYAQmXxv+Y7PI
1BjJrI9nxqcFrSedzAjRkx0A+02ZKlmM/xBwG3xXhWVJiwMfb4mXUq4aIfikHunJ
lagmwWs1r0ZJkk7rDlNPtWvnAU48LcnG0DZ43Sg0Gpn/GM0oI9w6v3HJslSWo+tw
jWIIIjO4uoDbkNq8Vmw/QKBZ9MbnUVpLPpq/+JUJ1uyAQnOAsMCx2Ppvx8dodeOS
YIg9pHAgGclRAwj+L+h4Z7wnAvI50qJHr2OfckhWH18J3JpxYGwTHbfCZpeV8CS2
Me9P7TYoRAK99eVm1l2Jt4HLquWkYefM8j/gQZgxIfMVZcUa+vAPN73kzpG0i0Sr
LBTRZdEh5LGvAddvlFYXVM5UMXqmNH1UOiiRXtlzBXgASwBCfwQ38QpOKBZlY9+j
1yrropOumTvYpt0lBoofk2Tru5HCMt5+MgUBOCmz5+HOHlOQCdDxtnIPP8qi/uWI
VCCpgyzYfBa/wzFv1rHFU1EvojgJdA8/kuyK2M/JAwEejXVHOdHTSsEqbKWBqJb7
keLE+5f3foRX3vIzaO0Jo4Dvf9nCFGieGxq/ePl38Xub1YG1QgNW/NeDtNATpogi
nlRtnF47iqdafrRR7j7AV733v+dO9TUuebYjcIY/Bwy12kQ+fPxYzkw65P84jLwz
352MwghC8aDi8aElNJuyP8VB1oBpt2K0fCUqnOO/QUg87GYwEplqql4bGvJy5W9c
i//fAr3sn5tY71X63awJ5ZWbnTuOitsO8+pLd5380efPiByaVhDWb6E0yHs54DPW
`protect END_PROTECTED
