`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xCEV4/HfEoOSVnudXK/01drrEzciZiOmJO2Argio5ek2dbDUSv87rY9rfIHqsagJ
PKFHDIEK3PYCbARRUskkRh3rnsuq2DFSSCAzG3kk1LS7EkuebsRRrJSSTO5OCQrM
ZWgOhHfwZ8VGbw7wCVkAe5CBMcnq50qoo8xXhF5kj0XuqoHjhgyQtASaExRBR5Jl
BTAH3EAQeOYK3McqH086YCqKW2V0S+KRGh8rNSDFKZEoH7yk3Byqf1/zofDtdKEA
s9ujcYrLU4tYginb5DUBTPduaG2gjF4D05iRt27WIDXtIohc4B2S0qnE8NgorNPK
1bLIgr+BcdGfTUm9zomFvr8rLfMLtJJXenKRQGUsS/+n8SgZBKfZPETp9LcBmgQa
1OECYL1dY93vYtCCFRTnf5MSIOfAV0z3Vm0jOs3Y1riR6SFp1QCUk93NnYJhOGWj
AIxsAaImW+Sg+FksRizFZ54a95HOi2HvU6M0cw4rnuh8WDq9F4uPtJiOUZlbyfFF
2kOX/klV+TzM91CXqw4Sgp+j3Mcyd+xLI8UIQvr0tRwwcEHk0x6myD3kXE1J1sd3
Fy4OUiVHeYNaCVZ59f/BTAOz4GrNznV6ZYG/XW/0iS6MNtOzj/ssTgREqJH2F8TJ
tzJvNZO3tWn++Lc01Y1iSNcXvpaEcHjreGbOHcnk2ldVLvn2vCPBsRm8kToSNrQ0
HwJUuuscLdXBhtpm4UJ3tP8FfPO8SBnZHbjApzUfsKvLF5+pCas6HLe6XUpUPkdg
ODmRm7/NUtiFZpEmNUIyFGsOTd77/ESXg0u1m3A+eEKaOKsosDWBFTtAMnKIFMmM
0yVTvNqvQ2uhfspAwiwBgiyUDq6xcOoZkbZnOAAnkn5NMGRV6W9bGV1yjheBZhDg
rRlGJAwMWOo4zvEuY/bOB9dujtH9+O+Tl9upOlqBrtB3xkVGnpAsbvD66ae8ExhB
mFT+KvJKhOHoZzfsRaF/7WgKl0IdCdIlVwevYiaTUlNbtREKgB0RLvwzSkELSdtB
py0q4znSaAp7M5h2uwZzyhHvKljZTYn1ZKusLRA1IuW+L8gSwmWGsecKyOsIBV+s
B2s912bThzBRzt6/mDQc+jFMZ58iHTzJJ5ZUgvgG7jbzY021d5ZzkCEV7FTqshzt
B5m1Hn+4yMZAyqeO11uzaf+ueqAgJMEHXqrryNn4yrmXlZHndzMHnX/l71IKnGVu
h2d00wCAOHEXi9Pcb2gU7Eiew2loeZ5DGgHHvVFl+QKy3wI3jX1wOcUSzWGt7qAz
O2xwtwlBfcLtrFUftwd/h5PmYoEk4qsC2WdSaPts+juTIonYS6dVOyJ2ajm/Fszw
jS5pMM3Vk9aZgrPsxX53xJMzvMU2CL7j6yV+BtzpdssSFqL4XOyq1NSSJrEk3mVo
g5iJqm8T/Aa6bhW4QkSj/c/hpVlL2dR9Vu1n7rnVwrjI93jikVdCE47QgZGN1cbx
7OvJZDMytMNndofPH/Qxs0Xlzmi0wUhai78MLtGMFPhupNaAdQRRsKIF8RzQ8bN2
eSHMUWAF56grv5GR29BX2g9exCQMlYIcdV1ruSe4CLq7DFn/uDg+HiYt7o8/7KM9
AfCDsvM/dgQG6Lc9GD/8DqopKxF/R3NO72omplzryLrk8nnjGEo/3pO/CVpRoDDa
59uI/IoQe/INEamB+M5XoqzlDAR8mmi8t92kLnz60ysRv2OhPoSSKDwQPOqI8BR6
GTZRuDFLuw4HjHSZ3oTwYcDiSB/QZPPdesn45glevI4Ca32FLT41x3s7/djIAFdY
P/unLkBJMuRU79In39IgugZ6OA7maai1SgzlUjptJE3AnbZE9+cHxiOLCJ9b4Jsu
fxaxk/X661orORIUOs4Uu20cC/F8QyqlY96f+SvJH2XEZvuhqDZwJaAfvOAe62Ez
DQgIjGRs0LmLWxSjE0PXIJ0rEv5fUmxVVa7aY6JxRyz1rayVdDFFG30V8cK3/3nr
cApj2AUxCbCiaxN4yljyT6jCJGLtPZXRJ4BTNtkwcJV9m1jC9H0LUDdNqjjSFIuP
CyOyLv+oZcpvcFg2NJ4AnFlH5Oe6DeZ971SDQ0YBglr5AmZ2olcARGg9vOiCpW0F
N6ieSWMGoQi7pMEvGI3/RLGykDMqzi2cg3NgdTcmivyrNmdK8SQM2XbVXEbXpIcw
lTHCz6jqu1vnwkxqLsLhehY3M6+SNfA1Z96TlHOk8f85+fwhFVHuuHnfeOBvuzEf
CBI5WdO8SE6ReB62qzumzJAKvKmbhJ18CwkQBohA8W/frvXzC72UuV0ugZZ6icLl
jgfghmgPasiRx4Rw7LHPhJrF37s/yt7/CBeKv3sGmeOVPsunInxRgcd797Azap0M
AwEU2X02lCoqACbNcg9uKL757d+LLkyCcFUhn6zq/e6BROgI9ap2hUIc5M7wtJyu
JB94Y1rYC6kink866052JuirCAi9n0PQg2co+xAye/1nwnQ1OJ76LfuGgMPem9bN
1buHs1RTgR0PrZgW5LbV+govPcNLQPm+cqCYIsm/fkf5/fUyNG7notbuyuamtzXs
BsiuCJlq+w9FJcrlo6/ThGpbD/SxDrxiArg496h1wIWkjqMrBUi/ImWhM8oCwxtC
BIqlUUqCwnNQvwPiZNiPQrpFeoPMbxeN3fKNCRQsxl1xBFijlKUn12P5fiQDB++s
fSVP8Q5HYVjBMeSpEpCOsbOmrFJ5C2N7xBa4hHyG/UkCozqUIdUxzezY+RP3Xw7Q
+Z6MaMqC09gpmD7bBjYkKrYuHz4XGXYafIJUsdD6QA86nCHLQqYteqBjRD/opo39
OcDhyOSV3J0kMavc31wD+mfReFshBAvUn/aQ1A6ydXO7GMvj9iOJmnvpfblq9jpH
8pK9mWV2oMm1XaY85spQU2jyBUo9EauTbp59bSpzgM+ObEejAxCINMULKEqnppHC
I2FhGQ3nx7PwNAzuMgzyGA==
`protect END_PROTECTED
