`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKBXuonF8UrAUtmhUyG2NRRHRzAR7bIQ42xq0NsyW9wULsCJ7eNqe3iQO2wL/L58
8vAJnNYz/RvC4leErYpiqYi1jHav2jGq9zjU+VXFQDQtSfXQAi8+L5bdLU4Mc1wM
6iSGqPvnaF2sll1B4wEjM8F9YE3+a/T+MGOpZNtGD7R9qwOuuuNv5XQyEBo0PV9P
kE0nXrPHwMuo83Ym/eQHWZI8rJPFiEAOkzT5u+tPDpQIZfcxU1VMFxWSjMDaRCSO
hgsBp3V1Zl77V7g7BllRgYuZrZCqWNQyFa16MT7GV2zSotXQ4ihQAhnTrTGLXvP+
dPi/i68GAsHss21iDVD1ZFlT++jJE2OwacAlHS2ylytFCZiqmVaXz7dOq6Adun93
ACGLeY2dJ/tsfynmqtd/CN4TA8CecmR1CKPAMNQHlclS/ZYlBMjFJpMpeBJp7Nja
AIN37sTh5+JVKJsIkMfcLnsksI8Tcq2977m0s4nJEDiADXrfaA8eOz8o/lmqbMFB
2ubIk2uirc45FOlhMl3XUjHg0Fvcpknixo0RFANJJjEg6noYuv8n7hZtQF8Bk3We
D2V8tNV7yVNM4jQ1YFIzuUddfszZV1InMqlWg/hk8HKdckCGL95RKHUsuscHyNyw
Np4M0ieeiquKlfMKJLRsCGb0XtFFEv+/4jv4iRXqt8twUOostHBmCeec0ydaydTX
qPzlRC1zThG8PBIR7WdTmMtrF2RjLlvMoOCwsGczS7ukSEKQczEC4t8dGRm2e1nE
UyujJRQbtFdCRy/z+8tbVqrGKslhnjiilMOlAMTaA/zlML+j4Py66qlA/0kkkqV8
PkdnnJNSA9HB3NMXxkUtAclFh71Uj0x3oj2wedKLKFPA+OEaGKA/QZP3QQ+dY5s6
rkvzVk7ufDdT3E+/uVEILSylmPP4zWdIV14/qQHuPwBXfxEfMGjzL0iSunv4OXpq
Ff+jjOKFyQx7+0LHgIuHtxbGbSkZ5FMXFKUDv9G0Ig4Qud7V9s8cU5bzfxI+OFh6
YWklezNzZEW5NBcvYCdQCmZWzUKW1OIF4SSrgWhKhy4KumtaNmxyWzshBK/NFDV5
TjH1fjwVQlfRoHWAVqbjV2LOphbZIWM0ym4ubcFPG4Fc+zVhkbpWtP+asT2xceK2
dsBuNQHIFTTMJMx6Z1rc7E1VDtfeRH4woJXqtlOFDN3DlfVEsl7jR4XuhU9MpfTE
dTeUK6R2pDFs/qKAhFMIFvQmBhI2Se7HpfymYhvahT29qGN68RZEbex1jEgFypyx
yG9wQhZD8PVskSJEoRGEqESShpWNYqSCpZsDdufqgtmOfP4vkMSu8kXmxPx8yl+i
m/a0b63TJ57y3V8W8qbqSBsUEXPCgcalkDqD+Xc6qEaFBxEEC9KJsOuxvjNI5RyK
fNaT5MviDqXq/HjASjDhTmookP4jrOQvIA9Ih2c+LfDKFyr3yWJ7xkufvUtZ/UB+
QDwobr5isiWedjLYtzBe8RPAR50aR/OOadoS9fTH9dEQk9KnS7n8TCAPclVaXkfu
i4SqiUYPxXnXJ6Zln9oIp1mgv3aeMXqtgzb30ioA5OHtjeeuM0mc2xSKypJESfPu
IAojtIOhzPyPIUiF7yeFRzHKRIy2rkksXDKSasNlj/j6373lANZha1sVUGIsBy1r
x95a1X2jUaQ30uxduCxLz+QQeyCjowH22zPFS9jSEgAYzCekBhtfx547bixpEO//
VpUjTIKJgiqaFDPs29cX73HTQcKlayUEgsKDulg69L9VMIEO7DlxLepeE4Ry5PAI
97auZdB1+CmaHq1F/Mu/eEpeme5bwr7w7CTWg0txlCdh1xTFm0w6bZWDADqnBq5H
qN959MoACmHBOot7rxIj+L1dc470IFkySRLRO4YFW4abnSn5nJws9PtpCX6jhZyu
UXCgcxSQ22OrJbpuEcIFK4o20PG8cJurydi2dLSH8x8muvH5mFRK1VSLZLXvBMjJ
ZXzJ6i7MHrRpDf2yKO/SSiDjScu9wtkdUUPnFRVRo7PK9IPnteBUYIXfVSrCF7NS
B2WR74XbdhJeKxN2B5vdx2tUVpoHQRHv9asHRaOulCyNE6As2FUbNbUIzU5m7PeY
1waSa0AHn6GNXSKFVuk/Dy1dHA1TD7hTIWQfhvjNRiHrIOHfNyEQM2znPnDWhuZF
5Qnb7q5vO0emyeGPjyOlE77rHh20yO5RDkyDgZYvorf7qQ2XszeJDvMGPSt6f2ZO
N9zpGdyX5De6Pm1g9K/xL2watolAz39J/covA5AhrCeB5bfvulgFnLte/oATVCkX
cZzya7o5aQSix31+V3R8toLALF0cpdrCtU5/K1CG2TAgvaiu/95EdbBcM567YcrJ
OjBYsi6C+BgSxQJf5S/wNtFMIVDQf/R3sR9IPdaCCQEezpuwMB3OWJTSuJTY03j3
gMPo5fozRlEjdLaBvwkSwgh67MZ+G8dHlQvR6R2qw9A4FxGWgPvxoDQ72YOTICpC
wCVadtkLrBijIr+MHVoUstrH8M33IDT+jvOxezZdazb4kVlDfYQLHZOU4eGdUiOq
ytcID9XOkpQqmurNppVPlaVuPrhd++pzsmi3gs2bqMSRNGECTy9bG9cwGdrb4GQf
9HMoeSFN0PWz3+/IdBdKT1uhRoxdggYfcvp0i05SGaKn08VGTcSvdBeAsxbXd4o0
UGDExDbU1h25RLwk/jApMfmkepWTpE0Tv8cUIbCAaX0UNdxNEtd1KWeVHGZKi1p9
Ko+mtwd0Ie3TBrRhS6ZDk1a5STlJpcp307GNZ3ICbj+pQ2udFmLeWM7UK+R/84vK
8tXwkqTrttQFZ/kF9Z5Hd1TgOJMhUGaD8/vki9UHGWZeKBq/daDsFTv/9gmDLh/7
a/diH5ee68CNF4OjkXlVfp7cmQFpR1LoH1q8F0SWSShAhIY7M7k9nSbopjxnzdS2
k1oiFeXPSI51FONtWwRuwPdGsFEvCNA70/2QTqjPYMiPrxQWRcf8foLjfFxQFI6H
wn8OoVnyoRu3TrUVe+zTJxr5WIeENgqhSUV68n7RkUx/gud/g9hWtaHJjcLbtLlt
z1YPJQkSICekycfIwPhowSy26lCJ6CqvLFzBQy0AcWiobNmeZC6PjxuVpNOE5VN/
63mtwWC2/mZ6yjcx7XYULGKd9Yt9jhYIqaQq4nu7t9bN/2/ct1vclBlmIAmJizrH
`protect END_PROTECTED
