`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7EyIO3/Kb8LSTyQpGPLPqNJeXMnDd8U/EjwEtMHX36RKqTmtUVH4s3uhAL/pCbrS
5Fc/WU6j+R9tTukSRIWAflc+rjYs0LTkIMTP0mrRhLB8EGvuDEBuIVALIHq8BS4C
Jm16c1KXA5fEi7u5aLDRhy/0Nj2U2dtIE3EXI4NsA7+bzVzUTrUiysYmxmHUJuio
uICoCTI/OEIQiyV94oUAZ/pbZpR82SM6guywB/NNwN+ZnQKc0y+spCYgIQuRk9BR
jYRA65mL7RCQoMgJavRLi1e+dD/erJlGq3UEqwOeJE1fFbPUQmZUHYjQUXUf1400
uzxr82v2v/xohYrQVkwX05SfEUueteGy/i0vZ6oRoFuIB+QinckkrZWTdtpqWI98
U6ZsVjzyaO4YCcPZ2rf3brqdVYdXeXsCR1yPl9PdSS+xHbf8KMqWUvYLadAmAc9g
X3eu+0T04ncPI3dEwneUhTHAJKEyoCzEkrStmX/HeP/zAt4U1Ml/4ZFdnBFeja8V
XdFRxZqBsxXpNnjeTTfwLskXPmOMl8LloD1lY8XKhWPE6sc+A1XicGFr4ZaNkB4k
uEAfQCG3J/9m0iJVpMHmcqRurmvI39JJGjgxR03gwxANrrFvIuV4Fa33D763pzzd
CZlIlD5S7tjgouSEuHOxj4VL1fVNKYGC+/HAn4zVjYs9bsiiQ5046h82HZiogTwv
lro81ZXMvJ4UBXjtZCO1W70DM8/h5BppJeLdhXy4dEtYYEzDz/piS6f9Yf+NbxYu
sCT+KKaEGJBLJSiVgaUFUQn86na9gN+zQdlXOt/p/N7NuLXZzGGVJJCd3Z9xDexM
+4+MOhyW7Q0AQOqgjTwz8qinM7mTbGWhHJXTnQOw17N+D72dV3kB4r+i52zWySH6
wFfiC+ZaIzZ9wF2oVibwR4KRhOZa0f/io+DweT83FeQz6sx8LnVeKMN8GaXx2SOc
Ygig4bIWk+CpEd+aYazTq0ynGi3cQKHBI1rIeNmjOmiXp7cRVPK8XyYGx7WRjmqK
dPTGXU844rH7zp1u/jhfD37XbOTHAIwmgkt3HvGneo52EL8vNrRTZ8sw5g3i8JM/
xZj21TmkMp9Vt0BiWEMqDOcqg2/0axnGz8dQeaazkTWalmuLToERfPc/EHLsElOz
upQAIMjuR7C9SZViu1x+2J7droahsNvwRLfl/FAPNEdbmlzfmQxqefkf2KDEJucJ
UfaoIneBpb0yOHexYlISAUusvISZHFYRqzDtRbVryAaOpRgerfU7OnxxiuEJHg72
JezZxJd8a8rjpyVFGAcApGkmpSSNr6/IcOH+pPnIP5QbZ/DEt1uAojrhRZwWdNO6
PR8aoWk6SARYvyAh2Rz9Bqcij8sOXwNVVbp1G71d7fQOXqWA8Zl1y+eYwoglCI+y
58aw+xT2t87Xz+RPVmECVEevKxegTxDq7RPy7u1Yzui7DPC4zaL4Ng9glLxGVF5A
Dn8obLpyAyvaqe8c9j0oY0vqnGmIcOUGR3zdojiJW1HgJdEbLD7e3L6uVUvc6jIT
b5XpvSBIjLZQljw+soLmx1WImIw8SdsNgPJ4iRsGeu+pY9o3QTyApKn3B9XI9oqZ
IXBCmM4xuW6lBr60tDyI/Yllq8G8JlU+IyDgC0nf8LkN3CpsTPacMi31VaK/kEhJ
qK8bGScOvjwnMqR1XmPmSMN0teVa8fC5R1XsSWyFN3oT4cSh/QtzKGR/q5wuGIMY
7loSvY9+wtaPfjTowUiUZvrvT4GDFNzL8k5qQxy2aj/q4j3HH/F9lOZiH4cxhv0F
GEq3CYbqS0C+BpK0IQA86cHwoIKbxEZUadZmNz9hC3jdxE9RYgNjwmR68wpH6Kzr
ChCbPLVhgDnnN9UVx3/8lv53KihE5xTinLtM/MpyR1AIJkLD4lFn/8C9bBnhwxhU
MMhV72ets8yuHhpVNhhOCxSa60QIRoNDVO08nLUcN79Ko9DGKBMkP4IfrFFvbfPe
soBdRtc7FwVrtsgf5QwFS2l2P/zx/wWBZJXc2xtifcewEel205qPMwy709AGsJZ4
Fc0zFEBpm9Al5Qew8al1G1J94YADjg+DvKL99cd2LACnhSgoQ5Zt/DNRPzQ0QfsP
Qf7/Rh3vEtczYQTXaQSEbmcwtI1sPEpdqP2dOpuQpVcTag8ON/Mj0VVlkun83UhO
IWaOyqL8hi3NE0NMosiSISVernFSEDO2g13KC4ByjXcTV79oRUrCVHsTjm4+2kVC
ArmgAI+CMupmuW7+GULoLXfHx0VLu3URBnpLSkHZj8xt4IjxcxDUvzDJT8HUGulP
42qZt4BmLXEPgk+GgDWfply4h+Gh3y7D67o9knzLq3XLm8bwfPtdN9OImqvT90qq
fjq4eeVAWvzMHm666BhlMKIOflO308g5jylzw8gF73GAUdEwr9kdyZ8y6diTWZcs
wv3oqP/lOF0Cj3jO+vOrNJ+F89N5vtxNNLDnm7SWl6VQfxojc5ct1KymB1uRO5OA
R12BZodCLlydMc0chLGkrVXIPGOti8SQXb/cq9t7dWR8j0jWaymIpWIxisafSESR
rLZb3Ufa73zNJw7ofkOC11edtPxerUJhrW0B3Hplp6CEdmKB0wPnfOPj83U6W9o9
ljJNnp5rQ4ZWM7vzsCU1uvKaxQISPc7L8CzkygGxfcXb+yqnYr+q5KzF5jwxFgbW
p7TGxCsiMtZiuXBc6HN+UsvZRGZKV3IQWgBg17gbqNBnUD58kBD0B98MPjOc7zOd
mkFIYcrtHHKpK5vQNFBUAmUJ006+dACk8uH9g2k3OIDBO8fQSygE7i4YAANbkR6H
uICMf5me+YHHepqtT170zC68m8GvMUU26cCt6NggPTpVVYgRHqSyeoUjSbKH9GoP
H7daiYV9ff0Xz48fXgDj8lccQQA5wdu3Axf61xn8RzjH8lT9KfK4YEO5tNGakYe8
ZL9oxdQyHgrVNy74dxyaQZXapi898ZKzdtNYPxra8YuVJ3f7iIWJE7UM5YnmA7Df
VlX3boMYiE9YzHKR6Jc9zyR7Ya5X+/V5HS/DMXJCzLTK5Egnp7/h2sbeY7iFRoyX
lZVgO5MR4ioQF4lcVXEQ5A3HQW5jlGJVO7Ktc9gYUCjO9vIdMBhtDJhlGSwsRd4a
UuXTgaT+er+5VScZZu+MPdaSgBxyyslrwO+ddHjKKpaSRWyoUAJvf8MW7+ceaYJC
Y8lFALOdPuijNxoLbUZMrLUXZmM6E/7VZgYqFUrysfrecP0Q1tloCTdbrumF6vv3
T5+DGXyM8F/vB8bkLP+W6bA2smU/CcPCTxjrskDnI2Vq70lp5+REMoIw383kUKxv
U/aBOj+2nl2SU3oQUxrdRk7Zy7059iq3yO4pMxhieBLHuokgvGm56IzcUfAjKYes
7W/fuF1iKn4Qdl8fxcWS9bsCG2XtsujJmhJSFEEawZGsMvnuriLWIz4GgqoJMLoS
UdulWrQm9N/M0I65RNoc4AmYJ4hUX0fSN7/vbPOKK+9F9udsuXkA1/3YGGj9t/Fa
DECZ6JBwdf/VH4NKQufItq/FNMpZlJzoXcY2hAc7crSef4W4P3643w0kDhHFx0Vh
Hr84zMrmnBs5xNqSxsDbFo3nrdLEZtjh6mGJYVMbTjZqmnzkmUPqa1L+O1G2PF9J
QcDFbUbdU4kWnDOPdigF324zzDsML76Z8r7KP3Mae+GJ+Z8TLMABnnulxk3PufQ3
myknPmaj8DnxwpoDmfNPFFZPDOTb4/wgUxMviWeYQn/f+pUFj4tvCSV+cSAj18QG
TzJeWT6ddGkxWq8eNeRXiIedCHZW2mLMPflltpPJuMp24TTHMHUnHgMQHrjpOz33
b6A01+to1c39FbolF8J+TlVIBYoPtzQjvw2I+TcqPMNjThXBTYJq13Wy/+PJnpY2
jQJ5xVEfv0ngufy0BajkcenS54nBu1UrVcPcuhsGriPaexLQhxv87CohS/8khZX7
gHsWkwHs5QpG0PljQ25XAd+Decp4PiUkUhXmBFDLYKCfQfzh61LzZgLjebEeotsM
yMZoeaXRKXJ9Y4CQdidvGhSMepRfBPNrXgEynMsIh/TQjbMjRWwdawCn/Tx3wAr+
9qfQ1PELfGPpdVtavQHECkJ1oVKY8k4smju9FhhCs46jVODWHsi0dYnRA3wZcNEX
wP1PREO6oVTnGzUSekGjUBAj0k+A7VmvKt7k1veM0/CMWgohm5mf9YnJUGK2HYcj
uJEcudWBZmLZPUshXCaedfUa6YoSU8HR5K0xlc22snAfIsgruCoxe5r57sYW01dQ
jgRsPRD7dzr22yfxpHsY5hXs4e0ZYeU97syz2gz91zEsZgtybH7zmUSUPHz+KRiG
XUNOSrPNoXW1U5pCmDiNnCiYYCy50mu4OgrhEF0t6mPB81lJex/BnlOsEcSmnT5V
UdLNYuFWJjAB+qVwhe5AjY2wKqFFyLFDM223WBHgVU8xRb2vm1Xb1ztCvPD6fupn
tSo4UpccILqVB6zj09O2VxpOxN/+cedtc+zDZj6EYCSsXhaBLCnXEAO2ULHgTywh
iu1lJlqaHnlDwwMEUZa8MpkO0cuEFddrMJXfXmy4N4J6Brs32p2r1FNSxtcNAvt/
ndVBWgWNYUm1wZB866fdbqraPmCkotCUh5aHTidqNFwpOCzwpLoED8kPfSCjsCkR
xYOXMTKkc8RQ70nlBQp2TZ0T+tIm5YQ7FqkGrK8wA9OBXlTiQeHYrcP0P2VGF77L
cKIEQIcdE20GKmA0es1rW6xb3/2gj3y+/ql5uxh2HxoI84vDZX0i+IxaFpQEEKVZ
PNAKPD3c28q7h8/xCUjNpCUQpiMqqbv+aT64+rzmXNG4jGtig3faQSDnU9g8geUt
HVCLH3RrxHyk3WtVyATwvGFZFUHtBbMWPw/5x9PuiHjdKTXt2Q1ZCd3y0W6WdcUh
D/UV7BfQnw7/9dCL9YbAIw==
`protect END_PROTECTED
