`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFfDtyzdINCrM1uggcBtJCeZM8i3HVGovXdPse1GZRZJMITvCME5zCDtn5JX1HB3
7xo9cwtQS+hupfdwPsZPWAcgWPhgnaIjvDjevL+WR4V5I7npU9Fm6Yc8ONA7F2VY
XDmVcDOKo1WtRQCMD83LD+Ls9WEIGWttd7zJB5sMDCUmNf3w+3hx3xGkkoplVBnt
AGVixE72coexCbOmBD9T3LLsvdqsu2drTSKaxfqt+BzCRZ2AxHOPQuYadJVG+rGK
QR54/VVDElbxAkJaWR9op73o3e2e+Z/Aab4H8vm7KFMmxioLqcfbuxS4e5JgCOAL
FspKfAOup4I6DDOo0KcAHnGe6zXXR2yuFoxz61n+hdB1ShtrGTA9NXTiUYE/Opcf
I6vbvh5hAjw2ZQetO3JvMxsHXR6Q3ii+APwIQ6ZIgFF26WJLSgJXHQVYHvYQuJvO
ZQ7KsNtEWdZylrEMbKrtsKu3TgrCg9rQcDmZxqKr4B802l0HvT7Lh33aiWc2P0BX
bWgn4Iv7xsqTSP75YrTY9wyUo7xUPpJso3puTQt1QX0P5BuLI0M5vJNMomSDnRYR
G/19rnsRSZQMa6oNyyfpwiKi6LyaAx0B2AfhxeUA6Sblf9knkP1hbXne6NLZmEUR
UYjN8dhbQ79/YlEQWnmydF0J43GhN1dHgx6OGO1V0hHYWQFO3yBvfhO5EV47/xDY
lTnHyxN/et9Eu1g7fxB5xFsaJu2cah1p9rwn58ln4wWQemmY3kt0c6XykK1Ff+VT
AmnEVwZHZNFywaigwBOveUUbRUux6frwQ3c50CwuP2bCjdhzixYsUXincCzr3LEd
wS/GElyXvefe4elf36ciH3SgYvjdkEXAtahQ8DegNohZl9MiSCJ85x53/yf36If7
KXCqqmgOoqgkEsItRNNyMV1iFTaBTjtt2Q8BGnVoGlpI2Bhbx84jeHXxby5v7vKU
x5Gi5nlbtPVsF0k0Zr4BFvkhNLAHTdIxTT+eR0XFjNEcMOA2rZKaZEFqmsBUFIov
zUjaYAgyJ1H0+ecvlAO4UEBIyvoGUAwzIW9JAkz8IxvAiiJ5Cc2e7eddoTQ6OPOz
AkQtMSaBmybAMoVLDcA5tBaW5L+c8CTO/3rWJ/QAoiAOqF5fVdMxPrlODDuVN0KZ
prxEdveYtM/PPAx0sPiZxg==
`protect END_PROTECTED
