`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SwOerGu7Yl907txJVUFU0rRIbA59UmGaR2ULtGVPclTww7iShiNqcKLhszIAs/6U
HEt+hCmbmtk+os6VRG3XDjdA5jvE/l+iqT0mDKbYuk9L8VtardJzNxAWQuU2pXvr
nulSMG9O17wSeCIgEvqGA1O5wH20crkiGNKgXFs2Rrt7QalCvSvCy5A7wpyEX40Q
YJrPSOYJidkvyjMXZ2DkYDjpti0vPufDSBp6vB4nGdkIlkVyGmsXZirJj2ZkjymV
1Rp9Ne2M08kCzP6uTeIpSR/z8d7CncaDfrRD/1zED6Jh8EEktb9++O9unBgpOgfm
FDnaG1u6vdi9+OPwUiBVvFGmuVhGdbyhfjO+dzFEb0eJxXy4eceHI/qTB4gnCDy6
y7W50Eiov4Fu/jzIEcOFwHl2UvXvpdlyPN/HXjBIk4cIle8cQLvi/4xpl2uz+tCM
VAx//cOyEGiiBY6zPgJpPU65E69K54D0FjCy22UXZ3csPHPRRs1X2g1819Q9t2Il
SO1ciHch6EwmB1FjeFzByjwyxdr0psPHNwxXbpJ9eGEmxrSv6dwagVH6ozjzxJ7s
NRn5ulmrkK0CKlO4n5QCd9IEK+X/WzGfyHvQmJ2BLpNtS62KJUfRTDDMvVi2hjog
`protect END_PROTECTED
