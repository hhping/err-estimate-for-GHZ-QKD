`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lBRFUoGdQ1eHnRELhvxVan7FfjNGoTNVq4WrE7or0vPn16otwIlj7+iCB1P/EX9n
Ce7HjxoNKFTpQX2ggNQxOfndbEO0cZ3vejI+2QQIKobW3MmcPaXlAr3Hon0JTf0S
Of5fODP/xt6yzwBtI+w0WRhP7WfUzUrKMMIzXjSOI0ecoy6bxEfJ/iCwRexpV4kH
IrmeXnPYLSNqiE/5FnESIH2jDnC/ljIz0tqAHuVBAvZvE7Mk++DW0jO9Pfi7ShZu
kAyR8Vaew3IR2ram1576WLAFAymIegQgOSUo5CF0dSNBs7C6Yo1Je1ZA/oF7MOlK
2+jmZln1diEDc7Dibuokln9Pu1aU+6L+lAlYPY/9C1aBP2545K+RxjO2BxCq8j3b
9iMrpHhgAg4Vpo7w4QHO0jOBh6HyATcMLizCpTb8sqDEMpuPzZkFWKaiouOEfLXe
sPWqhCH9H6WDLOJ6TZ59T874n2SI/2euvWYlAdR/c/dX3QNZzm2svzVg2DFvaUkU
SezZWtC3XwVuyQdVPNCcI9qFeAfZ21lrDrGTh0znGg3wTtW/7zlktKsMS3W/lE1G
XLXHzr4lMlI3seQqwjAmRKCgz4unlI6HRVhSVub8TiYnpy/XAmcU4VOC/lEchcs2
GQmgoZPeliWv7bCegm6yRwhkt+0dwvEcaj1uTlhkIe2MWCfgPqyyl2N2XRJ6e1kh
`protect END_PROTECTED
