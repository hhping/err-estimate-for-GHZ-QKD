`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcfdN+NALUr79nCoS0HKlyuqXLdsY0I2YpwQM6SW/Z5xffY/4LphBlwp+zY4+hvJ
8cl8x527CAFS6QaUsC8o8BVS95516shmJ8nkpRoltoms5VLiWMy8LsVAr5WqECOF
JgdP8YOn0Ht3F9LLavQlGcWVuXlLSCnphqNZid695xk6FP80gb0bBEhLtEDXBAPg
dJBWP5cnPPLEhGWZBVC6SBlsodnu+RGlKW0p5i1chefitb0sGh+KFD3Rg0zVrwCC
6YYczswu09CvFXI6cCGFbwWhSxrmuhTgyAgo0t/sHgFbnxqeGXTH+XGtYcExQH+z
uwJ/zo8Dfa9YHuQYLzqOQdXrROlS0qvf9U14+U7l6hL6yaSxzPryjrfypHphkFQU
D+1YkAWyVv6CsLcWpQ9FBarAKhMgrC3RG9+9PdDHZ5+nqH3PVq5Iy/sUlAHFh3Vg
Rz43CIgXqlcIQqnOOpPp5m/w/s9KdV5nXsh4X1Ln/kduy+IX2kPz9Rp3Vple3tJZ
gCsaa/wQ1DAAeX5sztGZi6Ozha2vgcJjVUf1MBxOuH/rAgOlpCBXVLHXuauRe4qW
5ZrwFGw4On+B9qFHp9Jze13y0LXFHUk46vMJo9Qvl5zokws7izzeKw1sKjhG6E4P
8cgJVJ0Cj5YZ4zkJP2nqGUC4PJyt+FfBwMeqEtcb32o=
`protect END_PROTECTED
