`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pY4kerb8bn7Jdkenjtdf7NRZp52v6TlRd/PR16kPGKOad0cUDy7D7soYv9zN+GiY
UZ3dOVKxGpt1ZRaq3FYCGzNMR3Ip/uTBIRnFD8FWYGNukQ6Sdjq1QStF++kn4WM9
hEl5HyCoFw9BHjCAlSqbdPucimW0HHeHwwegejRi+8EnX5AGPVHBpPAY7IRWNKZe
NXMdrO0hppNLCr22FAIH4xw7g0kfYZHJjmy9P9rNkFXPLkfpBc0b9WGo54myC+dq
PNI92Tg+GYxEilZOY76A7FejGU0Hv5KuVlTbMscyxGfAeKLuf5TstZf7PO84d7LS
MGEeADf6MlSefXI63mz2D/UeugQl5kNf0TqzsupMOqd0l+Sw39CQDnBTRz74YTIs
09c0+a6gHbA3W4dmQXJgvhTIhHP5Lo09PnRI6eDMj3opsfdMIFqTlxmx9UXtazlj
hx5ifrt09iTUsRhnikZzGvZRPOyh0Ub5RfDctsWBhcbEuT7Lqwwh8XhfZb3JraOm
SEOngbM1UYbfI8/H9vxglaDdjVZoKgukuONtxSVcG8wsJd7woeO8YFTPkwov3Djp
iq8tn0+ByZMjeHj/Uj5SAWbaae5NluS7sGVDz6B3W2Jm1r3yddGfC8LdLcI37gn8
WiqXSkv+vATnl+K9j8Iigdypa87K7kvWNULknp94uWHoZYm0/Ok+zg+Xg6EEOU04
wSkHT4rcyCTVsbh+ac7Eoh6OvLD70MyB3SqE2rgrvWdfXPdGOmbXg+XOBLMoUzeX
znhBG7oYwP09QOT39nKQRK1NoI2Sat/VSLxlLYuqdsItUtblAG7aWLbbvXCq6oL6
aAy/dcG5EW0KRJA7ElnRtEPy0pYiOxVKAcinG02B5o07Edi2bboEicgBjEsuuoNL
lkFjw1DBRR/sFPPzrZ7aygxWlba1vlP2mbv/l5WGE6T6GjgaKj9O3QuCryBKeM2t
QQ1NvGpi9ih92F9J3yN+0ciYtut1Z9zMVvfFZFt6rrFzRJWtaNaBJHzhUnIk90Fr
oVa6Thw1SRUBB0dHKy/Yz/WA1oCPRi+0j4MQRrKBXYW9BayElZT2WB++1IIcnx7F
hxOtvbAUe6x1Thn52Ri+V7V3aaJv+2xYhwuN5KjDNYMl+X7IgQQY3MKpcGHX6739
lipF4KeNmgDHI0wE4vAzyTYSyasd9iwyHt4trwXI6v2foMLZdNr0gXGyu2+OUXZm
noRHh72lQVS9kIW5smQloJKtgfkvuBdcvFaArQpcfs/vWG7RsGKTh7PwaDN8da0Q
z9Piw7ajf2QWtElN3JIv+3+wsJ66w9+atjiFliODbxyiUoMN0M0VFQcxNTTaaTrD
O0eVdW7o1XFuIn5u+sEh6y3Uil4TKy6plZuShPMi6KT/lYrkRHrtEilldL4fnKOz
nGcQmDSke3qDm64Jkscw1YHPO7kkUvogJi/tdE0Ad6UdGFS7cwKqItIkwQ7g07Xa
Wh6Ta74tbqr2xR2Bpl0rJQOfD0ivItteFSJ0iuN6FD/7CIQ7X86fN99/IY6stXgL
pksdHXpOj0BilVG2TodJMb9Jk8YbfzITbsMTKufFDWaSQiDijXCWhpEUa5VgTqEj
vT4SjaEiGSIfz30pKnQ7ddJs0+lQrrkgJi0XYpBrwDVavOe+NvwWmBBZ6DytHiqa
0mc2+u5af0ctEqR1llNUEmACPCPtDbOL/6MFJUoDhlTcvAp+++2ITTFo/K/Qrv+P
0lZy5MZrrwL7YEjlctopQ7c3WztYjOtUBZWG/hAgEh0o2FcZe4J6cT8p3jp1YvJ9
gJgsLAEcdH1OOPgwzMCedCFFfy7F3tSQyiV7q0dkoBEcVv+v5e0JoIVnBl4ZQl09
3rQpa4hhrzK1xoPriDrtHK8TBCRUGX4Pt6Q0VYO8/6znKW8pBXdB/o17SL2bwUDP
kel05BLekkKpUqrpwdbChMvYdA2RGUvVv81wTDONJY0Wxr+zekAnEgaMtYwpeQJv
uh3iycZ3ivSKGEEzhrtOHWk2ONOxnNPq2m/xbJY1xgWkWgKC+mUJxL+4XYBGHGUj
bJcqgvQ9D1dILKRJam81ITjXvpLULnC9BKo/qO/To54qAfXKbVlosKahKFWqwAek
AGq4dwOUl+vQYAX0cXhB3vlx6zeVN0QGMm0J9QyofrwusTIsO25i2eWJxt25ikyj
Zhul3XanEBbGHFtaNLL5iYIP76HVMROtUCab9ggYqUceG296sd1R1GVvpAHYQw3G
FS6+VjHEd9T46+SHkW2iqzKu+Fvc9XSVFNyG0GLIkKv86JLealBnqeZDszPqTJGe
dQyoGPJ7i1Cwpjd2JXGQt2zexXuWZjALfJ+R2bML20h7HE9hoOPKenpvgOa3AS7E
nEbnQWcRxiO7r7h9/tQZdRuhcWPISqHKI5wStABVSKBUcQZ+YjZXRZf6sIGc7d4F
2NF+tL+LPHNbLpvomVZi9NbN3e53TQElaKRJnoO1Z8YrcrYxcUKMYcNRzl4uukJX
MHunt/oKK0hHVTshP40GYoX3t/wgUe677ML4mBx8gDbd1v/kJ3ZG10cVmr8zZihr
S7dWm0/lnJ87JX0jwCr6tYOU6aPBzgenifTBAPblLR2CST+ZHlUGcq97CC0VJdMF
s5wlO7beIZ+jbIY8C8PdLiTjGyGhHgHirgsvZ0OWTQxbQUBzonN7CkyJg702EXkH
hk6lTTER00aj0nhwCkF6XzXOO5Ss6/ZsG/ktCbWLCsAmpGFERwEoBgPGCCs9Kdwj
z5biEY4vwZg87t0ETo4pyo/yeUzmmrVFW7qxKiGwEuSb9FQi8HvEXwxfHyITt9e8
cXW2ODrkWNQQneFtBKMGPIt0vqAvn6D/JdnyKcY3t6PqLHlOb9116bH6KN+lznfP
AbZoBcknnwhp7F75vwl2qj8FmN33b0K1pS8auemGHLClVMr7/sAuYbmpPdXxQDXx
i7snCJSc82/4sbiaIKEvkAw+iychwJbCRTqNJBm4IxIbV8jPHBzto7HNVuirFalC
ioIa83ZwmcYFLvuij4C7ec5dAvIpjDQjLfKzooTdOVuFGM4xzO6VeOdXGe4UYHw5
AON0karGacO8/mgMH8/xL8uflaKSh60uGYiisSwRxcgu84CxaVRZWdcfdvtujozK
B8TI69OSid/oF3WgcO5WKq9iaDEwt4Xe3LdxN3tO4uVaHwlz6Y9osEpyO2OH/9Hz
QxCFwc6yrYcggNdjDfwYopWJzazxAOGnWZhMFc6bpyvZijWfDPxYkQ/rAdkRou7I
bFSR3UZyqKfRW6PMTnxgdCNBhnmAsi+uUQ3Mt7yyweVFoVurq967OqM5wkNLQsqP
RlNOYLC32PCp5olLEYEkzPSVD6rw2kUC6gcpUsqiefYwaiHr1bYnLNRNJhMewCg1
INW3KPGu+vyIDS1eGQNFRDXISL13tdU26cRmW4phSX94bBLJEdwQR1BmMtbU3pqO
m6lplLipSZf1gH3kJsKJ53/CgG/yIYkDIvWiySbtd+64gj/7oRsuOomHREWSN7l9
WUNp3shs4sXAtTPx9Kk+kGV0YvmGp2b85Vq8wnC8ifI8lhYd07DXTAGmclD7D6/n
aarc+/UpYIn4qoTivc6wV5ZJzwhh/b9328+8v47ky114/J/9Hou0L8qtSOd7QvKk
B3eDiZ+5+A6kr37jjA2XLWfDpx5DnMGSMWrOMjQBt3xBrt4z7Bhs8tPKQ2eLhU/6
bUMegGj/1piB5Y5AgF+UcxrMkQkVFThUsS4wZCKM6ZtTCIEQO8f9V+aN+IVuH2sG
X0kt/cmtmcWTvmGAD5ZtvisMycD/v8bsT1qgWlFM60qpxHdT3nTTK4nNcnHEKtIR
B471RM05NBB/JrCw5AynpcWtrDFwt6xJoWRKYxRztgXh7S/JupJKtd0y4/GLdwhS
S7jTsQUERONPi0j3f29PP1DSMeU+1dz4kdujfAX/sAmR3dydaad6zHmTNczujzzK
ESfHk9/imcOX0vj2fCehhpFwtXTRQIU7EgUA9yDxkiEy4AFrktUYix0kPuqWJPIB
HAUj8DYvxgYTUZF0b7kaBR7efu7FAeMcfVE1tOGkrQ8QAngQF+m83cJ/jT+R+Be7
Fl+xjgDi7f3NCu6hS9DTlHs7fTfMYnHZuEFCw8tVc7AMqbBr1fSmUZ90j00DhXq4
H9XbIX1FzlQ/sfBSptH9r/a8PdEDFNMs9lepq4su252bM5UTv4plsKtVr3ZAbk/5
VRUJ4mk/yvoSnHvr7qltaSd4KuC4lGnpR05yl3x7f8RhD9xOM6n5HaB0UfNhgR6w
EV9oztAt40Ds4Ix9y4cQbKMNYC1I4g7kbSjZ8B/PsEl+KtZoprBAfnYHWcgzPkan
L6HpvHEoN/6wQBIMFoOayqTf0Ca3WUjWrGrOqt7se/fHcMwzXtkJ9PlACthmf8o2
u6zd0o3MVuuavwMLx9mDeHwfDK9yJW94nrZkohgE3EDkapDZ0AA4/H3D34yJuTA+
y5/BHVroEecWuw6YidZpU9Yaoa1pf1eMdaPYVgokBuMDkhMzXG20vdYivz6q1rU2
izIpBMKS9VqmBysVsdC0Ds77rIkSjTNS0JkFyX/DbYA7Qw6fwZDPv+2GhWC4fYa7
lctAi974N0ONvkJFbJAxA5qD8LLDaRuwkcxyhbfCnSXyEFlIzGbn2u5/JfHjQvNS
Cui1lqSdOCzBrguA7li1P3z8KxlHurlaOKUd7Mv7vefNkLlBzXHGihF2lBVvnviH
i95O51liZtokzfemCGRS98sw0frFg6lCCZ0K+gG81sUevftjMtj1+p5Gu/m1mHCG
vDR4DM3X3wqR9uF3SV6jzkL/+2Nszza3kSAcZXx+29MymtyhnhCL0hpmmGtZKU1m
Tj4mS2PfpDY5NVTYp8W04b0TLrM5YDnh00gdfUQtXxzdbWsVPxL8j5EKHhU7xnpC
aa07CXJvOLu6blxpOltsKuOMPPmFTbfmzapoteai0CHjaRcX5E8W7fMEeyZhbX1H
uKaM+OZnrhQMNxWA5iYj4cus8SDaZsgTVqa8Ttu5MQUGZXeTXi5etvgRYVLdDzdj
ql68hY4idynUhjg6dpJnNfzO1vtRiswI8nvQqTuX8GBYFk3qFMuNM9mVyka2P9Oo
4eA4yrc1CBTXngPUpj1zgvUGU4iC+98zTHQ13pgGJUwB3FwD3dsa2RUvERvksJBJ
Yw5rHZGzB6rpMT9QfomrtrfhqFo48tAZypCN2vjTzc2BC4FC7JNZdVBRiITYJEvH
FKewZkDrb+88DN3rzQ2hIT+ql/L3zD25nDkFf/c07xOJjheh6yJ9lktixVHyVnyz
T/qlBHw42jApzK/UgDeXn6/pBFedgraUfXbgBy6ZbQjvKPsakR0iUF1aeJWWT0M+
josSwHW/soN4RIZ2eHy++E3QJEGb6pNrfyU9WZQ845BcA30ZDq8SboOvSa8ZIRmf
`protect END_PROTECTED
