`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxzh7jL2gtYOwqmuWRLivs9RtnqCM/3X8TYPMu5Dw+jdFpY7uftsyU+30TNttmfP
dtNnyh3OPxedKLZa8ah7qgoPA2oOIDCFAHldyYsnZ/AgDWW0eOALmuXx1wFNZ01E
RwwB/mHvJEE08pPnpZwYRS3IA3RHWq0FDMdmOIqedMbGr1dEhj8YMT8phqMwpQYl
Gzjhi7QkiLZ8x1jGxHgpbhUMb3XtufcH3CFPwsF68oql7j8Lk7u31Psk48zu6Jn/
kbaAepVkhwP9QFnECXsS4+jx34AyXvdfK1Zq/3X+JDktxAOteFuFVEjUWSq2HLGe
vNb78t91RnF2BqVGrkMZEvDuxMARSnXMp8A0L5YBxlhrKTM0J95rjwUWc/+I2lAF
izf7QKaTKD/orvOkiUgkq8M/nfGI/aSjGA5J00mOewk70AT3NPGJ9mvgVm/bGOK1
brbqGw94759cHisQoxXVE5Mg/7vTTWqgYP0+B3A9nsIMUIEQNnY2wExoOTBxHprM
/3DhnsY0P8L0MibmODi5RX/i/EORatLRmfrKTyvRcQdvQjpOdiftH2sX8DUDTHtQ
3lq8fJEuuUSbrHCxAyJAryshY3RKu31viM9g5JWhNjqNYEfnWUo9RxvyNmw4quvM
3iqIczm7Cu2N6BhgBmNWZdJZMawbohHQdFQuih+FrADbarNm2VYRiICf0j03TNB3
TAhHRo2mGAyTjxbNIkFDdKxu5mGJNpspJDvd1k16yeoJ6sRy6ec93EprVRrqGqDH
e1X0Tlo05pUJ8QPzsuTcOiaDwlFkGIfKCG9iLeq7aC3V/UfzXnrHL0CZhNUHs337
a2aZbWNMeMYGoZn9YRtOnhz2/NjUEZkl+wgebpQxyLAReKJsFdbagku5u0Zh+ohl
YmuCPzq9QNvyv7w1J6OauiRDhUlA5Xrc63X6fJFzXWxQ8nzMcQnDkE550hwRCIIW
wqD3i8lzAQZ/N48xc9TlDcSmiKIGihwIVf+L++F2tRZ6sIN97WwAiLyvLhxCp+lU
jP1NpijJa4X8dTJncTsrnqJJmWT+HBtMS6xvBHs6yNUKUKg2pKjZ25wE2xEMDi2b
sobXHJEsdzqHRswKN2wGq395InYXFimGwmMjahfFu4uHazAqTSDueRDzmCOFyaPB
oiup9b8wPNIaZKG/LrIhZJOZMFK+oaM2bBlBXoxgEboAzawxysIbkqBop0deBlZy
tt0nCJtTeyCCvt6jIIOccROR0c9skCjrjitm/LVO+PJ7sfsZ7GdY0qDPlZLKROy5
`protect END_PROTECTED
