`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLAVPOwwTOLvpA+hyHHcsHCI+oCr5jghD7YRt94cBX1r7/4VfyA7FoHCKf3l3bKD
gOvW1jGWjjE1aOu+ssKtQTRstZQ48VM2swwd8ho9ZPIWoy+wDJ0npyHMoseiBYJx
2qavsHvFh7g0Rfl7nmMCakTvSgeMUNzhvG/IUluR1WMjxO2M8JOwGwi0H4GPvn2d
67veYCP0W5oBiOKzJl15Kw9+j92tHIAMwmAslMfR6tqbIOgeNRUB/cd3hOZMFErh
+sFd1ooWZ+z88bV5NVIgPZblayI6UxNRFWdkyq1pqBsdqBjcTqF61aJZToDU8GJS
7W4wHGTfONpcJTCcYApVr0CZNsHANTGst3QoOKKDzakOR5B/MgWgifqSa2iGRrv4
vSavfupLLoDuumRitRm21pXBf3Rf+3L8EjzhSYcWM5SJlExYbLmVnol3eB0sr4t3
I+P/T+zT0sk6IDXihUd3evX3mzIHnKCsZXCVCuCxI67MI0YojXPkhcho433AP03u
mp6/+iH7lYUTl6lCtgMjHUV3DlnUKCJJPVC7+xGBkaOe6LiRi4QBWd3ng8Nsn1ym
QepusWq6ONORKuWC2Hnl+lqKi6bTwS/amFGpOhHEB+0GYcUeooT9C5TaGE/Oce50
OqvCCKglK8FVLa2b/dGHyIZCXaKju5/NeLncLx2xoiNg5SmmuV6KMtFdf9F2J+CZ
SI9Q5vvWZbbqAz+CGFD+UIQpI2Or6AqxocG+pIi3OQgSKdhLGhw9/0rWR9xyjjBO
`protect END_PROTECTED
