`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XZN2j4gL+tSTkZe2sgfWAdKHVuM5wZhCw8kR/LW+IbsUy5Ku4bamaOgVwWe53z+p
ObJ10hbILIJbGO3wjxC72mJJnK+5ysd57CKwUHsorONR2NBjpxK3bcBD69Ddyjr4
Cny+ZAxyHPte301RkbeU5eHGzCVR19nJAM+/bxT8/1MvdEEJW5rB0ngRiZqboSxK
tlHtiHLOLnOMZT83k3riRKnYLkPoZfhKcGfN84YpnH1gi9A5X49D/tcEThLtKL8X
i3rfzNxQBTS8qAL8rjKPPBY4rw9dKqD6XoZP791BE3f2hVPbb8huMb2ArxbHa9bV
Y44NkN3lTK0fgTYDCKjzcmNEdlj4oqrCHiknFdjNDoxdnXWvErtztseh7wGlV++F
Q5QMVFNcf4ExhDJTzqGQF7TADEkig1V1xD0DOks8QCYvrc6J4XNtZvj+uqvfRe7Z
ZDI6OzXJkoi+BMjtzE4SzrB8qJwYPhotuf3BlXXJ5EcSGTbkFn/o6Nl+jAnk0plz
K9OII0NNYjXFYw44d7qpJZOi3rJB8UXGbm/ZXMYRj7kTYkRXVHBeOos0zDqgicTt
0vxqqni3qM0YR3zmHX0bMw+0Urvb3wiLlRKjMiVqHpxrPF4e9tVjSEXVefZN5CrZ
b2fo9WBOFfr+s1JcmEI/Z/ppthLg1XUFr8rRS3rIRcbuzQDDPFkI1WH96xgmdFgT
xb08z/M8jJZj6WX3kyUvN0V5pHlAlRnzZIq6hGfddeXyBVLOi6+9Xw0ULPShVWla
kNQsDhm21Ot2EBvDK3EiheuuuxZadFzXaEj5RBE2qgE=
`protect END_PROTECTED
