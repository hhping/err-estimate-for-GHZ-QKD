`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mnFLxDphWJMvKiRscVDlC58X+sbQHHHK8Ykjk0S+zNKALoZbB8H52glb0UTHHk9G
U0KPpLk32aDzx++SleH1EU9me570gn0/MLIWsPz5lzE91k8nsoYi6hE5HMtOMAuq
Jv8T4uACepNhx+5fwGfY1NIKrALh6eNTV7f9GCNi2Nc1L3Yqaowhd75Az+NuusPU
K3GKRg+V88l0hkMrqSgZ92XCTLx8RstuBntyDXJ6+Wrg1EOmq8ldDZiPqvHKjTfn
i6cNhIjNqYWz1rOGB9bhurvkbBEK8//Mg0a0782ehJOCE+DLz/7kt7cl4kYSMXyn
THLKY5pWTJBjsGQ0YjtwzELyIoOl+AMauSE7qXPmNASUFU90nzqzCBAEeOT2dV+m
EHDN876J+raOvrg8v4Q/IBTmby9fIFJgI9km8OkoNF4YDT7bYny7vIKBHtalPc39
kjr8baGO6tLwsEteTNsSB+pSCMGtFsiRmz+WjJX8OAM/fJ8czTYQhukoG/Q4l8CC
S/uTU3Nk5GHqc/5A9EhiUmUZZHfI98F5QpniiRjvb/KHNXXc15N7jaBjHgD1+g8D
Q2gXqBECxY+Y8FsTQBoNk5R591NDGjUl9I42xR1cy5TEjcpPLEuytaagiCnL4Mh8
LZT6mwN7zi6Jv5tUrGj2PM4KJZ9g5k0Mzu5zo3bDlRmQ+do+CIidbOnV44LrM/23
Qn6/qlLHq3L9TatyBqSaAR9Jw4I9Zwb1ypwuHqhkuRT2NpvpPv1dtnZc7KaZAxSw
q1cLMOrTy1ItHZBf36tbYb6cH5CqVS+rcGJIabB5NSXN2sjHTjUW2OVzUsPPgsGB
w351YlCiSt13M+qeqMSESaSzFfGg39Pu9bLmFzb8/Opq48j5DRtOBzQb6i6ldVBS
VCuZUDMP/9nNJa4z/cvvj86d1LPkKZSGRaeUZeFgLzEEJoXZ3werdQ5Qh7IfKEMv
V/DyM/stK0kkGz9O3gMWizfaWfNehNyKEBBhDUCo24mWnuHOZ9Cc7YK3K5V9C6/q
8DADP+SjD1BzWp7mnvPnve03+jHrVTCb543ZC2bxjnSy+pAj885GC74FCjNt/9z3
tEZinVQyU/TSC1WfWeiS5rCyRy6bv8lCL6JD+uRuAimFa6zzz3/frBR7ELkmuSH8
8E5dLVEy/0ROCIGnCaijosPFfAb8QGABP2HJV7HdWHkcHvE7EWRZ+H0Nj9IEoFBi
CVAj71JP0lhuiTt3qLMqYgrThQZEnL+V474Oo4r2jVq96EkVVPM18Tiaesw+EOPi
DuWIlbuDmIpCJIO0WZykDwCDlKbSzbXpCLnpVnMfsziiY3jvsro+MDMsFXJmTI/k
UiK5isNj/VZL/djj9M5q2lD5NN3ytyL+BsrlWqRkLPLrVVLPo3ghFpa6fuLKxWbO
h5F4CZKLu9V/23HX9nWqUMBJxIGnlSZNfxouuOqatiLw9Qo0VZp6+qczdn3+aAis
Gex14t3ouw9pY0X5RWbSl09VvxNGf4fUxwnTk8Rchi2Ug9bYO+NyWvQpeZ1uSnQc
sI8TDBRM5G2SMYMxG5JIw34psaA3r7V5r6iACzuJ0sTDigXvU3cY1BTvHhJMKaDm
RyyV5MZsMegrNWIi8Bm+NIgpBWXIIXqUwPfG3D36lNyY5+NfdjUJ8CiwgGDmaP+S
oZBCGfp6L0qdrC7gDgWt68ZIDybDGhBrFvgrIZCPHuo=
`protect END_PROTECTED
