`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9Hb50bZn397hbZNObXvyJHLUONYsKXpB5PROtT8IKXWvwQdvc00mPDyOCgtvYUv
TtjQWAI5u/vt+bYw5R2I7py1KZmxAliexAqEVwNP6Bmn+BIy6fWB8TDiXT3c9LbA
CB0kPktB9Rl4SWZbgoFBfZakUdZkNw1fA91OQKE1HkBxgQ5NbSuLU7T4fFm03hiN
VIlEanSuPed/IJzBdWmB2MXybjKaMr7OOg37ydbHqzC89BPode+OUqMvh2cSvFA2
2bHeKWI2dMZt+0siUFklklEVgwxU5x/VqJgrfZiDvEt0+Fcj2xUUBA0f0EvckMNR
Z3RYEDbRtasSlgnPYLSKFzRcFE5ixejdW+++swdRYH7t2SrXheetDUdNJHkhItND
L9hnQx25cAVxlJ2Gdjpx4cBKV1ih0SYd8l8Dm6xA/ENof2jProdqMIXuaNe0wpPH
d4EZHd8LMto6whsTFOYpK4qlvPctmTh+y6aqmXySwRLLC7Z2sd38HkF66VLlmpaU
KGNobI9dzMdBnLCmbqq4AJCEhurggH16Hc7xYsKTJBgq8V1vcdJC7LnjZKIAI4mk
89oszMm0Q3hbMYq6rge7U94SxqBUZXprSvg52y3hc/RDb1IEEi26mi+/u0JydPja
gMhyrmt8V/kxDpFMEEG2K1AVrbjzM1mm/oJQW1Tet1iumQ/SDEB0zaLydBE3ghWj
+D+PXPwmBKptEshxumRPlByBAoBlxbTbmlAzYy0J9AN+PQpQY7JlX2eylMI16dUN
he49HhqFdMGNUq4sdNBfwADvhVrA5V1G7O7F3EAIP5AyJSHzH3GCO9jIUBBdB54W
mnEqD5zVPge/1cqVjjyQVIROtLw+kCYgEa4Av+rdS+C8S4ngkb6fXRn/Cmaxb91z
RIz61t4nRAx5h82mUrO7/gQ6pDJBnx6Uwkt7is/Jz01/U7AP12rD+ltEQHGh9ZHb
ZB56g5+0G/S36fmFntatOjyR8BsY+EJldKFPHhM3RwhVbZg/prXeT8oOSo3fLSI8
+/7awy4/UN6qckp1MZQFOjYpanyY3oWp+Z/HXMfDlipdAykQ9BX6g9IuaPe1ANCJ
CUGQCcBmr+y2CXMLJF72mpPuH+iFtFClvpU+7PPLH3H0h71ltfK1gTS6+sJ1yLEu
knDdwjNmp+OEZEhFK5WHDumPsehDJGWr3YkQ4FHFOf78x16KjMSRaM/zj3Ku/PKY
zMWQUDT9/UFYTNuTrE4LuX6JHUtraf8riJwDfVZTGcC7Vxj0ixZq8nZ0E0pzmEUc
SodeD7PDG0pGqLNeWCCedCdzQ96qi8z3Ms5B3oeQtvdz2cCT7XYf7ODXigMxOskg
s6u/mkk5MEQng/n1z4GGWfAdEycgUgRdm7IH3XUSnejRYlPilVEEkWS5JifPcY8I
jroGsJ5veCHliYv4g82Lecn1BsE9ECV8TLxAKmOSRH5ql37QFFghE//NWT5xc1f1
UtdyGviGdntFXA6V5GcBBPShmBmnSpetWNMii42UTWJTQNjY+fmXX/ls5th0E/tk
UHCbBamNDJxYhsGYL/2+UuDSK2yCLXvT5DpDtxHBFb1ISFQLHR/xX478XMwTwNWP
uE4gEaQwLqM2uEmMoRJ73Qfb1529eqBY0iiaUoRZwVbZSNNEsOWasEcFWjEZaU4b
tRKMH/UQA3rnfTwPfWG5ZTmGrRZ/b0MfK1g1BlBKcg0ZO+yakoD1Cg84J68Z+/DI
cVSZli+RtC2d9XlMa5tggFOqFpQxcMHunR7tZyyCXPGv28B8tJg3v0068+YYfjHi
06yiO+T5pik4b7b3HvLislcHXNAf217ddwUFKGA8eF9PXzkI/TFwPcxmERA/sgVJ
3BwBjJ4lTHElbuuVcx6uaGJhpAKyAcjFR9EgR1+Fyg3Y5t1R0ynhhehFrVQ0nDgO
Za1LsQSRzZjAtmQWdcUjWV5Du/IqgnGUXoN9M2lb1tS2Minlsj1rrTFd63/jd1wz
n3OxwdKq83KncwJACDR6r66o3wk6E6gRskmUbPmb3NbJNmx/uUiq1TnWnKjHJZdq
X4j4PNHwvHmHK/fSbJKLEL8Uu5gNzOHjVp4dTkjydJUpQApyOxPrZ2smr/1ZPrQK
ZG40/XTzFikdfXKOWJJ1Z+aUURXyw37lf+5bdezPmLZ3XtY1lEbyY4C7J4qVV7jf
KLqms0uaDZTbDi+hU/3yS0VTnLkqXRhMPpzIy2T7CaEHLgYouRLhI+xfEpB/diOP
QKaAiGQ8Dks3RxjtcGX/0g==
`protect END_PROTECTED
