`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4o7fq6fM4lAYxU++X52mkip9MYakJlshMjm9vPjtN7QA42SJq45jtZcAam08apR
mSbgEDwb81PQzxFF6BtBWQpa5HnmXNDQWLtacCUULuuYo6/pWc5BvM/iFL3f+Zbc
9Hx7Wt30GmwzTJVOum1/VzeKj8PPxt2Zgn0ShKu+aZYU31dLDfvL0CIHyVySs63Y
tUyW+IcEZHVgmzsT4rK0EeqaAXbUUsxfKEotdajyxnDR9OZq5dHb5BvpAX6uEQYu
fkXPyHD1SCLUO5PwbCrWN2EvNC1y0kf7n4ooWTzi/97c8GZL12jo3P9qzLRNCZqF
fFlDVXaVbsaom14DPvqKsmPupOUr30m9EqDYADeAKY2VVFa5/vPCS6iCGGmKKOcV
P+f+U3F60BVj3BSQ1uFuAwGvFWLAxE+1djBlbjlRMeajTraMGGxiRyfw218/SWBe
YRpa23Raf8GEhPXOOfePUF1HtWCi68U7DH2rxgrVMeEWO7t+U0I+ck5+mrAtWvuI
25cZl3y3sIPIRctG5x2haGNHaWLk4PQ+agOobj7aVgmkf0w02PStFw1+35VdEvYI
Thdp7DULG7erVrU8aug75BQPiUL+zYiwGAcqAhgrjIJ0WgPsTEHo3+e/16hmGsZV
tuOHqHtR2bRAfd/ctFP2UX32cu4fk7Bq0m5d4i8RKKM5V1Vs100nnNKj3VaCx3gT
oF8WU3fVJBwXmANVTU6c94IMtIDaCz08RTIW1zBB9vaiESh1gpxBpnbbMB/R0Nkn
`protect END_PROTECTED
