`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZLjEqTIti5yu3CgKP0TEbTVCf3jMUkJd9G/2SNjAuD4QOBnBS4ObJcC55bolujb
4E2iQz31YsDcClcZUzvRh0KCwhwiIUGRFo4YbMDd/nx9PBeHrPyzjs2losM1tweV
nRPy5lCNCLVpOhWW49rhN1ZVuZaOfBnSa3KS9Ld5xHyPCR26oYyz2401WayUOHpc
dLCslV0yWQAjdcgURDCM9qTFU/jvcnXOG2CVIs6CrapJNT2Xda11OP9GU+/ZbaFR
tDLZnAInJryyH5dSUvIe65q12PIwI2x07agIYO9nvxtj69Yn2OSvFNbO0UTIpKL0
zx2onzP4qvWU9Iv0YMDXqhYbYAhpACndvZLLmQcjvTaaftYCmMJtEgJCv3mlbLn9
xVouIR0LxqCNO0IlqLfGd1ki6pNLpV6NcDRjO6ap2jtv12ckXi1MY3USv8jJUEwm
w5WEi6wo4jWwWYvIw/EWUNkrKzEvAPLUsZ0v6ycnHYZTYFGWPgptPV/CHX6no+IY
FecSfBWS8gQt/HhrnQvDr7JijlubEwjgccxvvlAAGMb0YUEGyfKKvZx9b6oH6Sno
LSzcV0ai+sTu3lpDGyEHc7HvUvSvqr44GMg5Ov66y23MuFKCzBKQl6GIXpAbgW2Q
cHJBmLDNzDiSworRmKlS0fXPgwhPwUOenaR+31ftj6M2hiVjdRoTh7UJT7LEBHMW
2iOfHCIjto/zqNfn1qVv7w==
`protect END_PROTECTED
