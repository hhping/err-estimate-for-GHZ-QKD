`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8anXiF7/C4wJvsQoK+Z60yxcNyU87dqPDdBG3Kz97Y7+f/n3nCN0mY/n6iAaDLSc
AUU7Se+PWooh3xXgb7vYdUm+oQw89c7Fg42M+UyFbPi8ZhrzZ2ryVfLdWNxt5lF4
ix4oVrQqugY5aGf6WJ4/E6xm7MLB9EUd7fYmNK01WiysynaA678un3PodvpHkID7
KZikxBywB+f1jYfjzl47CZB7gpc+DkhI5MEqL3ihByFKaxLQSuxGiQYYlrTRKW+s
8uPau1uLdTOVorFXMzn23TO/JyoYXks+bViyJyRTXBLRDGvDXV1M/zB58tsjHa3+
1IHmdRXqSp5Py9oWPrAlz6WwEIoRbtI8AONUfHy6wKIPHDBeiLk26+hMlIZl+kb9
Srti21mhbfiDszT/VfJp6+X2nedmB/RP9VmGEO4x7acjC8BySEESq50vo/YWX6gb
Kkmbqp0lSZaMlTgK6nVtSl11tMknHR1wAk1AIK+Q7EHL+EDTZMzC/21ydfOntqWa
r+uW4tiu5oO+e8Ql8RdIe4h1zoIu9Aw9k7jsu0Mw01G3pAsHvW80fQnJfT9HPjZ4
zpBbkVfmWNIAP1gHLNSLDBuR7/84tj6qOGfRWovaxLD4/AnJATHYQ6V3DggxRXuM
v6wn8XhQS3IOTvvsIwzEUPZQHr/PAaCFB9L8FraC+b3oiOF9VHWePcQ1JSP88Pq6
6VFpOy+sqxuFvkglgEsnAZwVSc9gjVB3eK0kfgaM96XrzQd+iVyC8JFKFT5MJXCc
cxMoshHqKQNUtmpnmJ7yruM2oMKMToCuzBJTDJWCDFl+iZkxWoodvEJyoUVE8B+x
EpPt+A5rSGNiR5zhwmq65EafQWEqAHODL3BSyx+aooayxsOQxECtrVJZ4i6SFGiS
9SyYtQ+SnTPRg7SycZitb1hkQlS+sGEJ3J7qyRywo9SVdCuPNQVle5WPjb+r7QOT
yCojhQm6Ua9U4nvtQQeMrkc/RDtiVeKQlUglVEdG2Pbotnez66j2QgIFXHulMM4S
CneDSkiLho9HXXccB+CiDYdNByUHZjMAyLjcVfyM/pIds5fMhMGbgl+RlmJZI6i7
sMUI5nDphmp4b6YnMPmMVoJZ3H8/QQCQR7h1o709Vw86IIFdeBMIYW0LWsTuFMhB
1zIk4OXu3zj6qrjN5IKcpODTsi0YSwBTYAznJfUwZqLx0ecLm2rDzcvunPLjG7jP
A0tdZQNePtVFZN7DrkqDb4QXVaVjxVCEsmbxwKC0XzcAXYX1t9C4cinbTLN6jKub
+f/P7Q3c2QFI6Iy9J2KxpAvmey5oyuqerrPSOEBYJbRvelarH5VspEMA9WAuicKF
QkQNThUHuOiG2LsiJxsc6yVhKwH17sfDbjv3L9SPioZDKa9XEP1uw72H4UnzmoWn
OcHBCPJB32L6VBgwpZFD7wMMvklDYVAQLyrx4YQPmzwlwNDLF5aMLQ1sbakpjKN+
06Da4zKCv12Qbuy/hoGKBvMCycpNAnu8befPS+bZKvwsxK8UMEr5n2tHKpPJrbPQ
h8+N+xr9wa98q0cqraurH4/Yeri4CB2fMG6yXvT2XzjpGjokyLx8DLjvny0b3GLa
ZFlnypwSnWEvsoHq259iNIJ0hqC/ZUSIS2S1sqfgdIqwcuYQMi1dBuxGxvaQ003d
ohRzhMA+PhwaK0uAadwzVA==
`protect END_PROTECTED
