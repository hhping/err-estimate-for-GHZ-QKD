`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FED/LtPTVMASXg4uf0uS7PErzw0/fcMcOx62s3JFZBfwVowUaBcp1u37vrk8WBh+
zmQBg2mAvoxV6jB/hBCarR0S+bqw3EOHT/uveroQOyfNfgXiRunDGtsmeQC6P5qQ
+fgx7lbhiFeChKfhAG56Judh5HF+pDPhb8CNdCX2Az/t21JN04fPfaQCXmDhz4e5
hz9kM1RHUnSH4yPBP8f28Wu51Tw9cZHSOVKhdE9mLOH55/1WQgIByRoQbRP7YmC0
8gutyfYTBXXo+0cNZYljIZqncdPKe1gOMv9BFyKyhEHwjS+mdV6NUbJ+KSmOyzl7
BD/yG0QrVAi6/yWVcFyv7n/oYVM4Ox24xnYjZ3f7M1ooiW2+wKAscQi6HCpewMo7
Dg4+tVy7zV73MsuzmMqVzv7Q0cmIvhSMDKupUreHY24=
`protect END_PROTECTED
