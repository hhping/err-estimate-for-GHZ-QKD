`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jXfKdnwvZeOaRXN1ACkrbCk+5KazjnroF9rQFtD5YZDgQtn23LXe5nZwIZhk1p4l
QQmV07sPHf5+zWyeXEvUl4wbqMqyjxvYdu3C0I8i09C/gWY1Z2UJZGNB0d5mIhqj
1kH4ltNhDNQ/Fl2s8kpgLNvJdHM4Z5YbdhwixWqenTMcLlNwuLvoDwkeQ0UUzd4E
oAnDCROqcYugfow2XFKDRkjjlwWOYIr22ZnvXKcSoj2pMtPwBREyKArvEVyMUD0I
iANNILt1nuxXnDTIeRYjDfwut8Rm1ARVJLoBOdz5IaiaqV+xrxY+RwwuxWusVHe2
h+WQeOFx5vX/RspIs8YAXgbPmo7oe7syPDTRQmqXBs7GDRzLnBBCuT4syxZ5GEzU
QQU1Z3mTV75ZLLDLLjMKwE4zXEYrKrwWWtNPxu2hX5pEETqTZIxilgMcM3KEFgUw
NAqF5ms1G8+0GsglVkZdenLgTi8HHkCRrWsEclfG8MvecAWQqgn1IvjpDd1ZQOvh
2PXjTuxFaZrNCM6NVAUbw3bO1hO4dcRJPGcIH5+Cf2RdxkdlyW6FSIAo2zCqMbRm
Ld+0k3wgbATiEeYp5167W3NAXVjWg1jSqHcfEJis4vSgVPBRg0FVKSeIEOFhgl5P
HJkfW2t9jAjdwER4lDY9P2ORip/1FfCnsv/Kkn16i1I7/t2IieNGO2ZegADkXczl
xkyfhYVI6iXxUQLqNc8JD+8UHPt2hw7uKe53NCl0bc/W/WXGZ+z+eQrJjYLocobs
OBKhR0oVZDhj+XqlgM9r2ge/jf3BSOWPU4vinSMxC7DV+Jd2uJBiJ1QaRMiuxI1s
3s99P7Se56b7TkoaOYA2q5BO0hSTQDnAoy5vptsp6LRMKJnUxgxLhtdHxYUQDe+p
XQjqUxXrUAXL5VQyk1h98A87Izy2ghbOONYTTmB3hHyHP+bJq4/AqpeGyJgcVuZy
EJKmMkNU52qGRCrBEiXILXHs6sAq+XTC7uw7DboC5VPLzrG0aSApWnRwBYYYYfDG
m4WZYrpXjk78KOmf5j8ImeDlhQaJGWbKNGZx5IipT1W2m5STBlOR5+HRSvAzbNhs
KadK/dJDqirw6BmPUKrHuQ8965d7RAIFOG626mN9cIWd91Hoz8dtIJiHC+6xqRs0
J6/K5+rO2Yj/BxBCtUxg8tkuw3SSWM6MqhJMEKrQ6hYEiE1UIRdvcl/Zk+gJZvEl
T9J3RJT4KUzEXo8Gdk1zTkTGXuYeV1Y75bxi2FgGs5xpjuX8QLbnUMRtGjc9y5ej
XJuNGSSkMqx7hdlBY+YUsCwT/AyomucPu4VeodF2s+P2QX+QZGeaaG8Idh4WljY+
Bf2GvH+0i/OmHtCNfGgk9sobi0fNr0UzLZyzcEpwYm52ACU0UWGnZLMCN2eTCCxg
Hk0pWHbtT4hK4fJbw+xUwD/88PFRYYPsnsXU8lkWP+NaZlI/NEgsOOC8JRmEU1Tx
oGYkYBz7szbOqrtutB2WPG/RaU+L4QB2nlPsAMg3E21b3VxZJPXdqkYx6XG56VxX
Hs45Y4onV0u4c+fcVvv3PB78+t5vt7BbmpfOeZycb57hfmZxA9k4E+KI1YG8RctI
dPnkN1scKT3mR4kNel63AT7/gT4qdTksalkD8HItrfpjA5F8/dwOGLOaSEDu5HHo
yW6gx079GyNSX/QG4a7CuxJCIRkQYh40Ye01LpJ3Op8XRfTHNuL+1bDYXqk0Kez4
3qkaZtr7PRr2sCMUNd5L+sKZrstAqjZrFpg30sEoHmAlTdCqpOkjHSDyHULjeQfo
0B4JFsEq5KmBoxs2D2PBC3tDlhk3MrCXMAE2GatTaEkWvA7QV43RPR7QxpG92Qmu
xZE9BXOcaJ8G3s4qTpib6IH9WHu6B5I5H0cF0AVnfc2EL0eHTCw9FxZo0MLGDXG+
wNAHaFIMtkVyTZ+a/vWlXlNeBJhoIBcIBF5sT6Qb4Ls8KyYFVxKmNJjCLwHNtO5k
/dV/2GX2b1V1kbgP2HPAlv1BREmrI3wjT/XOSEIYiShc3LdBVwm3JmijlVezDDt8
oeJBtTqn4riDdrzPi85ebA5cXI8auyHTCkIFVk2+83XfJfZIFBbZtMRe8jCcCVho
PJRgtvoQA7VMN5iSc999a5gi/t8ORbGfoPubtZ7MNnoLAH6wqDtPyOZaCvdazIwJ
zi39INZRZfiMqhG1p7sO08GLAQCdyyG+b5ty5ni+W6vp+quYFOfJKXrQGRQ3REkc
33SlmYAfKEsJIgLXYSmK2Y+9xwLUE26ElTAp4ZMLi2K5t/o57NyRf9nW/5xIqwgw
m1H7KFkTH/wDBDkYYHvH08tH4Ui2qsFfyBx8U5bIyCGV0NeX20HwhGViCw8mfUfq
cfpaZgNzpjt65Iwy2HsJJgJiRkaJe5ScSeZuDpDa+s8FneTMqNrGxlmjAUHW5JRE
1X7SnunGWkvRdBVAeIdMahTnLP7QthkvOux7yMrG2BfeYf3InsbRnpzWkEmIqE5O
POfBgtGdpNOwtv2ghRRN+K5V1JB2oeRzsx74ys3zpsxzdWn8w4bSC2kvKdEujwui
SgCcaW/ZholAUL65xMnPRSPm2H/WjsUGuflhhwL7WZrWgFL1kraMJHzghri83yQN
1u9Bk288Eam0olHQJbcX3Q1+/Zv+YCSoRlEe6vX5Ib8hjP6I3a6Qz8ebZY/LnZot
RjjnhwYWRUa86nJhvFVg4Q+nUjj8m3wgnQb62qsIUZA4f9GdrB+Jet6z44zu/VjF
0KXVDt3sdLqxnyWmPXPriv/izFX5/yb34Y4mDlHSSYRZNOD349EwfzYq/adYIfPV
GzMAdY3PX3s/s58bHpWWavcmj8rpJ/oKXw4FHCyz5vQe2SCROvCZFWc6+AFENs9b
oq4KO2/89y3z26uV+R1yAc281DJvfvmWLoRH4OgBefmIGcZ44bmr2hcc2VECVuze
j0cuD/PnS1EoolDtC9+yAwFIYyjOpg7soiZ5A9R6/3d8rGac56JAAaFT1cuVgT0X
8PoQiW5F/WZaWwv+LAlrWMAswWultpRiLRF7Dp85NsDfjYftJd9npOOLZkV/lbGn
Q39+xvPDHTbyo24OFCcQyR+RK4n74ChwtU4MSnFERnh2JBclgFw/gHWcp0+U1Sil
x/7+7mnxAHSIosY/jVIH5Q8czSWlI87GGt28TzHbvaqUTotZzNin5mdSyOPGd4xf
84ydCvk925H2ifq6RIVRaBLCWEgyNfsjIY9XAaeW8Xho1VGsIVOv3PnWrZzCOXOO
u2RKy2AapECdZtiAnaCxBnVtDnzTX+DWH2jqUU5jCNwtupRxFTTmYKBAnb1Nna10
tBdx14jen2lJ5XK8lecv2TYmBXAdUQ4MrLFLXE+6odzGIkn5bgErNzUFQhN5JZ5s
QiV42dhzlA2k1uu/u07qNxn+rezgxsrMkwnCHNETECw0SwHXrVsdOvRefjc4ubKF
qo3npD/f8WmGwXxn0TVIuThrt9wUtNaMQeBLFbfRnQYJaFSLBYyFtoUSOov36Kh7
PvTJswYpv7Z50wpFNj/Hl8WsZ3uQz+wcpEemz8cP6T6S7NiNnRfT+vgYa6S3tLUC
4aNxGfKHTkYquO7nRpLLNbE8TDoQF9qsfzI71HVpiIXG0W7SvZ+4LL/dDVSXM7yE
9kCBTAC4BBdGCy8tBSytdGXOB2a307YoCdWedEPgmk9xsQk4Me0bgGgpOv4fRgoZ
Do9RhGJpCmbNo3UYaItclPmRlsnDgil9iTcq6nvQuN6cKjcYxlyv8QHYj15gqYZo
HLrBH/YoEU+ym39qU+PHVkxutKOe6m9zz/TU1djC4z6hl8BSohlZGI9ybAr2ZaMw
bvlxKO9CB+bK+9i7r+MPDrGFvguZUitxcOdOACVGY+8XQbInYgFPNIC3wUcCKhrj
GUU5DZNwkNXXKOJlG/CHNxONE3QtVTQrGlBPLcOwei+aZ4G0qOh+zKi3pDTr7UaN
mQu6NQMRaQpJQgb9gpKjUzgLeErNiid6Qm8UPLkoIU0ldXvxL9soAgmZMWQUQPWJ
Y2fdvW38WgVpGlU8mZTuGCCw7VWkmznB7i7pxXnZxvSYyNS0B72l2pVmFMiCoz/2
1QuwX79AhoxrsQHsQXKnFNgY12dwPHSAzfXQaRhU8OrVf78kTTJNOElLIwjF33Lv
HbAM0p/93CEDwb0kw5/E2hpL00AGLFFF91BV7B/Ge0Eqp43DpcpxsiVPfjjxIt5P
VaLJ3RLUqt4CARt/OPmVuIO5vTP+S90LKPPWDyxZuZ2BTol0WfqpP29NyoOF5Ep9
KbEt4+WeM+4g2+z6xDFzL/6pZur8Rb7Y9LjgFz93k6Ns63PIoibOc8JurPLCkzMQ
`protect END_PROTECTED
