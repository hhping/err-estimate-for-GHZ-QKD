`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AW9sHIF+u6J3QI7+U+KHNjy+HYNUzYg3iJ/5t/TgURrWV9tA9LXVj7zZDGAAB9/W
/JQWxngGWLeV9DpyyPnW1fMxK6QYC1h/THXGYQ3paIvlmCByIo2dCMPTpYt9CgK3
qHQ6iciJJpsj8TaF4Z3JtpXkBmJF9pvgPYwAZMue8M1CyWqUbyuschy4NShtsvF7
sID3xvCIPPwLU3rHW+wPjPJ4u2+fEMLUlFYcSQwd+5YP79HW/lw8NcHuT491dFeB
MEgwqo8ze/LYH7XlAOQ98n82eyPRktYB7TLkTbvLWbWxX7MdGDyX+xWQvES3Epru
LZtV6CTBn3ULlq++gjsIpS4rlztgJNQ/MVdDNRXUMoh5PdGIeR4WaMYDE4YNBgaC
PmeAUsWNiEt97v4T18OvrKehqML2CPACsoak6Nz/X35d2PQ4YP1F50ud523pk/Ih
CealN5r0IY1b7tUGG3t3K5UPvEtfrJIi92eY7THHRNyT84LUL9mwqgFBakpmGA3Z
6aP3Jj75gXgpdXbeDhCSV6UNxjRB5DF+/cQIhMtZ7msLY5O+r1yXEC5BGsy9d6Lm
1j1rBJrxBsYDCO0tRKUgwUwAiyx8UlY/qQ4NpvsSxSM7Zk94+WoWXXx8/4r6nOq1
JlzlKQXfB5MqHM7w70hxC6RH1BG/mAcKaGsFkRLR13V5flbowqPUpDCTm57MtRni
blc7y2tG9gKzPghe6leQryOyf/6Il2ZQFdkTpen0Qxkr/A5zFhgPvGXZ5a9YFf5r
Fd8EZB/1EpVhhi+BZbs8QME4B2NjfkGd6RJEnj8B8dc5ATixMppuVKqjZsjYWx1Y
qTiyyt4Ps7qfsz1hhjEotAYSEKoZpsCZRUyIVq/P1RzgdDByOLzGHcYVqP8VPLN1
iDS/q8EQ53Dg3+Glt6KWbze869yW+9A6bQjmdwKITgZ02QMpJuA+a+Qq7Jgy+IxK
LpBN6jijxwTEJ7QA6Jf9ZxmTkZgHVTTw6QBSrVhWM38yzOQuWUrdhFmkFMiUTfiC
MpdYPzfxTyJd1aWbRPZPlZnnWTijpHA8y7fB7ETvWk9mr8lCQfvHRx5qmuWSRtJA
vbLLUaoFmACljDVTpfOvaJHadfOU2dr5z7A1hZ/BkXOLW3/0hFTouwpC6Ul89r40
FYxPWk+13h4uED8Bn7wGHTVTTUfHPqY+1GK2a+D4IMC3r+SWRfqJ1kRfsOwuTtuN
TM9W8rTKMMhYrKHTA33+kw==
`protect END_PROTECTED
