`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PvHP8TcyWKk/jqzSaKUovOHiU5Vs2mphSgvXFtZkqgqVO4IYCR85hWOKrkqX5x5H
7PV6lNYZXSFoIUcpO9wSobedgAHVgmIZ/tVMdo63btuv9TzeqLS1aHsb0OwYWmNw
dojNt9t6rkEVl/IH/XkUQrd19oEw/9sobP+DELYzy5aFdoPOg5InDJ0LersLTh8T
AkxMNvv9+iTQtmhZMizr55oyNBybWmSP2LBqfuU2JfCv3BG7S3PWKH/aj0DpV96J
EE0BPFPWsNfYwJvchTpBcLShsfCG5XnWf8JTSx60YFbBer38zflyvu34j0c8UqF1
ExCOHcy+gcd28etVbUYWYwC29bXkUTrLIel3lvNKzRQ=
`protect END_PROTECTED
