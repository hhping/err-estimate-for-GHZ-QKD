`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWtvNByu1LBtmZ7mI+ak/JZMhtOsbex8+9z40rMq1y3CSWnMByy9EvRIIz1AyXut
aTnGSoW88++uatdhLHcWlkQB41dd60gZfAWyY77HnhA5DE0RaTB1Qtq5kvpTJGRG
NKmStgx9uBCslraaKMAShwRMhLO9m9Fse1vNIeBabuJXXGANshlmLWUOhJztAEcg
RQS5bNugK1XZ8cOJe39PuzHP0x4VgBnlJO+BjyuzlHkgx3gGdMvTYmGnabUku3mU
/GgCBDC9CyO+ngmha6nii8jWwNoRklh/hLb2BhhnnJb92WkUUrohkXMJ4AiqWKiK
vqx2awqgAhU3SDx5FNCFVtvipm7lbzydfHCR4/KQ8rA6+HCluZZ21OY9XeUZeR2L
xnRiTbEfPCRet5TB7zm/2kcvI/WTcjSno+F2F56YrMVHQ6A4zN3QD2G2BwK8hmz8
`protect END_PROTECTED
