`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xu7W2gBLbiFxzVSoe99GmePNEooarB/ZZxcM7i6TuNCNcRPWuAyGf75EOD/wbSmi
QpILckZ+MUtsOcNzlAwf0LviVSdmZu/aO+ZW+xmooFkFWsT6NS5RVfU6jXEFZK+P
fSDesRCbBATq8q86cvj4kn2gVwTbtSo6Ce7dYSMueSBjCH05/RHVRcljaLFmyu9z
e+02e8Q+Rso1AqA3gGq7M7L0kMQtX+9gENFmYhpQHQV30EA5x3t8o1T9sYbBYdgg
PIUqzNQlGVPUURroCB7oDRklhrlgyKmDRgeBUrNwAOKUA0U9XD3c7li5ukDupqz3
c5Cin50ejYhKo1KEoAeEDoGbWEnDKOoMLkJq5D0een06d6QN0qKn4CGY5iE//gAz
VFWHum7tFGqYlpuQr1OhSI/kRRvoeE5n0OJVs/hBhkbd49DBIM4UScjCpEFJa/m1
faQchMaKg2U4/rWi1vnPMFI0FeAvVsckBe7WorOqZKF8yghtbcVVZo8vsPrgTRtr
4xUDkOJ+mcD5wFMa7t5N2RLGMvNRHjGpSMx7n/jxzhOhM5TLAiEup6fGI2Hz/Kh4
V0OkfgmWOU1T3QnrmX0i9eQX19yUDSqQbKvXpdpFRiDBLOjSkSXaAcjc23AC9QFy
iLLMw03PAYqU9uGGzy8jLXoi3BnlbwQjtvFr0PkEPAz7RFgy7gYQM28vGDASRIX6
ZTKe1OU4LPzQYCWtIQUy0p15DeMio4/QJ6X26MABHpj27lGy1OLF4sta2mMGEo+k
jHhMxc/DK/42BwiQsbry+kqsMGpugZVYOaEgbWVG4RrDIdc77Tutd7HQ9t3E54Kp
hxSdA8amrXhSjwECv8hwUOd8k6X97hZqUz+T6x/Iy6VrN01SEq98b4FXQUA79X8o
/H297NqTvfjWt9RUktn6X0V3coZ9pxe7nWFVy2TkG4uGNZBG/qE1GYvhPQgiIG39
kI61lwf7/JnMhaP+lOq6SQW1rwWY1hEAhYnibVmMo6lMuwMDKzB6rYP5w4yqpy27
ihKVx15eiGSrU2v7bqxrDp1cD7BdhSxoxEogwj8FPZnVyKCONmkmRT8UaehNN9jT
VJzHY1PgiIWBqfrWx5+x/kn1Z2kGxXXsiaM6IuwS67h6VufJdh4DzGRaMufc5cJ9
zaf2z9qT7eJ40/PsAqoMrlgWbF1YFluM1xTDDIHgE7ODvAhzxlspbBFO31sXheSC
NWHEn38QIyFS6IfzVGPrEk1iF8cJg74K8ITxn6htrBpwKiN3IDUckp5MbUzxy94Q
Vy+ACfxPSmcN56TQDA5nvX9u6E9yUlRHP/5yzNU+NgXPrNiuEl8nfh8h55qvb4I6
DYFhXvBCxHENWG51bbm6zQ+Wi8Gxjp0QeQjs3g0arV4mWmOW1yyPumJg+LmEq6u4
81rJbgwlFMlXLxDlkXLqk/gxHk0zmGTbUVXZo69kgU4Lu+6cOrU1MUrxCkCEbtx/
zcJswlVA0vASsqAXosAj6frL3BHstTLGELITIpnpC46j5eIq6NG1jOF9kqbp35q8
idXpSNyzU+7u8ovwW8PakvjlGJ78TMhwMMEVQA7E1IXdimiyh7mpkiRi3FYh1w/X
fu+g9yyzu3MMbakRf+ySQaBOAKs/GH0hZ1lcnjXWG3LOGSDmIsVzq0xGm6NS4UxK
WIj7SnfbZMlWHs6iWSiFXlMhtiBL2i1hqmMZbgL9qyFHAZ5sfRsL2s/pZsCZgfjs
eEXt2MZJRDZMZETfDeWR9Vm5USeZnf4FVP+YwEdlgY3nxG957m4ulAG7dcVW58gv
m7q01eXmBaPC68zee+WmDeoBe4aecWM/hSPCW+qbmvR6mDOklKxQKw1gQIq/aYNv
5VbCXX2NxVfVB+OQ59MdnmTXao3L4fp3ZxAQvXsUf+4imWkq7XpDpjIQTzpVSz5V
t3ppMju5WO2OSC2u7C+8hki4+KnMeUQI5larm1kRGHpBrLnLs3mtC0FKC3yDug5t
6XRcKv4pNFXrKinWhDTL1AqSmTIAQFdYcJmH8pdEEr3KjwuQznIl/cHmaaYrejpu
oZTPi+15TVbS+T/OirE9TSBo1kOwc/j6ipCsZBh9CsARU2k1cleo4ujvQo/rgoDo
yO5CnkKoK9pL+nVKk9fSinhl4iW44fPnQDLXCXKXhiHV15q9Eec3nTITOBKcUKV0
XTqVcUtJmwX5hIz9OrMHgCu2DnFQrMGd3kbMThoPXgvUK7aS+rTh2X+CeM9CCKhg
iHOcBCpZ/FRyWLXWaGAw2sC17OTaRqkffKOUMI5xpHzinBfZsyc0JW4WJItniX9O
pJgFCtTGUja4NTpHu8EgKeVfnWFfB0j32zDNDTuHm4vNIFMTF4uhxRcdv1d9oBpJ
hvFi3952WQkozNjeEsgQy0AGKFKy2GVSRlq5mgTM30meE8tADKK8r32LxPXnut4+
xpRuFlAabmEmqj1DCESB5pYmtt93II+Y9l4DweVzNIrrYZIXDkPtMHWBzatkRo8H
EUh46BHPQa0u51o7dKaHNJNw0ceo0EbPNmqOth62Totul2E2FVfzN8q7/aAg/FD8
Aifzkgtaq+/8c0MuuRPCj25w1wN4jOIsdqxO0CrgMo44vGh2c9aSTUQYvndPiWWC
`protect END_PROTECTED
