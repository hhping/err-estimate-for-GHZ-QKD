`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAGqih4+G4Ir8/PRSKfpvm9oJR5/pVWHCCYWPio3tLo8bkHwAdKEO0eZX5hgYcJK
lnG+JvJGyvacSlHxVeGOdjtWvN1ieHdfmlTd9uLwQyfB1Gd5u8F1yOXRECzfVBPY
9nI4WRyV7OCIKA6A9ImrvsRACOvHC+AoWZIeFUSqZy2aJ7B8NmYxvsLl/dDh2PUj
zALROsniD6YTTfpBs1LlWUsoVXDVmN33n3PY6W7m1f9hPTG3f+Qjy75oTGhhwPQN
7xGsJ5s3Rw/+5HeCymFW/9+OndEllERqXyEkIAeZ0SmLsgjiWMkOLKeUjJyps2Rg
m31ElG76N6kM/NlCM47kbBfp8H9hxhKQu7WODD7Zx3i1wK+tzUAjyqaVeb15lo2g
cxB6Gw060idASuqlcxn7xZgelt+ET3s3aufh/jHMZDWyzu/uizHDFTz0fPGsmU8H
LzkEA4DEjTvvqpLr70shXs10JZMgboFHMyl7VKEjhG79Xwx6HTdzmmOoX2Fsus64
XjSHM0U5yHMLHPCVLQKjEAbxAg4tQs/MY9XOvj1Uz2R6/oYk6YlZEX9Gkj5ArIV2
rwm6HTz8lVsCW+mupONENiQuEPCOto151ekl8JEXoNyFORFgzXP/nP+wadqisQA/
UylHKtDNKY1PCPwQRSRxUK9tFflTnDPe6XBJCN5ryGTOQlFkUI9uHiLDvMch/Osk
AVPGYmsuchaqjlPZ/d+o83aOzGtMIJ4msIQhThbmr4F09kiu6TImq32x79DVenjW
0mF1N+lC2RdErzLFOOYRWwVJr4cchUBe1ErBGzhOqFdvHILcnXf7kSOyY8sAuewj
AZciEqvhp4dPJF92/H9XLME9qL5Afb/Ff/hrK6e1J8OnrxswcN1isXZRey1bchZC
ubpp2vp+PajWgsmjuvYmiroCDZmS1DoGbuIs/0rtgZZRzVBhGLn4dRLE9uluDtTa
uWAVHwt5o5MCl7vRSVLCHUWFCn28BBcI+k6nWc/tE03m/siJqNjBGYXbRythPJMl
i6H3hcZQh2g0Jp4LmcCEXULVZZT3XSJdRUdur4PwVYjNpepHEPKn3FIyvksgE2cU
l8TKILxURo4XiJAHgyrZZ7XrRYRHEJ/R25QQGOdqqpsKH/SJ0Y+H1R16uDxI3JTJ
gsskgNsAZ99NZ/KjLf1ozmqRkU+QQjHZoZ4FRPKGzCvPmvpBsz7w2oF6XFPE3xFV
7SoOhRu8HMJ7nCHwJ6mN15He2hSv/ByAU88sBbgxuxjDsbilVEtDG7RH/z8CsGRw
`protect END_PROTECTED
