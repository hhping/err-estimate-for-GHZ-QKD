`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PlKkv/PcrU0W+0PCdWBwLNXMJxrBV8H7LwpSlJcLC+fPyiYd8Y/DUTO99UgTB626
mOP0bjxLEfNgk8vp+e2ZnMJ7KEXiMlTmvfUAswPQ5gzz5+1XVQZsJWWf8zE6v036
9UvJkHLTHE0UiyVRrSRmv4LD9VnEXKBlgoz4P/n7t6NIb/hpC5VgXTV3cpRT6kdH
2oeNJmE326/kv9TpuMsezQ/mRigrBVHIsnCTyY//+nH4bkoAX4TSuT+WebRufwki
rtcqFwTDKJ7jfz3UPrV4cAxO4Esxc4ghPg3RYOvPAsYSISbxUSRMxa6pM5PomUgy
zR6LRElpfx7197VidyB/xKgZKpF4sMG8mW65QjeJwT51OLmnM+3e87ipA/2zghqG
ScbSUiGFz2TyySEliYgjl0wzZDpYo73wmYozjNOpm2F6fXSn4LAzfw46sDDXR1uj
++XhFoV1n1d0fpXFFSZ74zlp2/87n2kPAOKPJA87p3IQ+wh+7YjAjU6hrSrZ/udG
fS/OO7rjIuKuRB4Tj/YLnA4KixEwME3y30NEDCCCMfX/FLBvoEKuW9HTMIJsVmsW
7tdespNVrXrlPawUZvuDm5lJtmQiaETbtQfdYBzQv5LZNd9oNcK6xxcBDkNM7oGt
hNC/9zxJJGLHIMt0ADZL9kDbn44LeHiApGNTeA1M95AayV4vfpmuBCWR3DYncuZ/
wzKdkaouYJSSrDgPX5di2EUkTokxoHpMJvdaIVPxL5ug6B5dGuSDmtJXKXmFRo4c
M+Fn5NrrnwpXngFqveQFHaN9sywwx/6Ju3GKSJs49u/Nu/4SclCKQFS8/p3a3ASm
`protect END_PROTECTED
