`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+03ZgiRGZpK7lgPscl7LpVpa2o81o4Ba2M9sFej7JSi4a3cHyhYOUZUozm0Op5R7
VTqtuWu9mN2f+fH3hn1/lQlhE21GYW16+jAoW4IPj5qvnnOh3xJbhADVmTEBkAeo
D4/zf2yRT7joROZXWU7ka4Qpu51m2p9aN3+CXH6EkbdZvbJlt+xeCdH+rBjSc3/8
na+W1F9ujR+CEJL3mAFSBhOPAF+PNkXEhOpOsbW9RSsz1pcCWBw2fx/YEQ7+ojEH
3sjoy0YnFmP/CT6tfmqTqIAbW0K32a1bpcNEJDoqrm6je48ML60ji5WOoNFEB541
JKove0BiQvMYnozAWMfmYSw4Trg4suyStP7mXQpP9qIq2CF3EzLFn34k6Nk+3Uxq
7eALHFuqTT0aTbw6536PSUsyzUHfNlgpnElit6ERR+xE+Vq8611gADyxPYe6NtuW
SyCopuGS8SM+abV3B4PJOrqOqfAHJaA3D2KwJngEUK8rSM7os1q243q0gzdHsymA
RwG9A8QtMPXUQe0GrXAt/s2/nMAgzuW9sLdxk60rXysKK+zS4F6mZuXVL+V6OmIN
mc3tV34geBBia1zTnxWRSbxDijez3qwVi3Bx7n/ihA5mlpnv7otaW5BHYPMSj5xg
71YU7g+fvWZjrMLtyxdAZ852ZZJUl8cgVmxEx/VGovInq90Nycw0JSipLkHa7RGF
T9dJl8NuK/IMDKey2yl2Y8zn/4kHAV3pXHroX2Lk53MxQRpas7MA2sRgw+XG3rlk
3KBmxfAgx7w2wiNKN/gOtlqhxdQrKBsqXxfoA7Urcq2ultT5AdKk0ggHUw53pMW0
XJwealgjRZpcSht04c8GbghZWULOb2oMKNwGR+xPleBIFi5Iwlpzqn1K8qf3QQVZ
RkZz82HCamOM67CprXNXaYNCEPhKy1GscFrhfXybAKr1plbFJx8WmtN25Aucc/q+
NNLZX2OKbciOFI2Wus/de0KQNu/K3bUIrWCILNVlDi4y41s27Aj+rLKCgmm2IyoB
//H/a7KAWol/W7YaVmTtOvcNnhvW9tf3OTTZoNHeslC8PT61HFzJVa3ODr1AXOR+
IvBuRuAaHzgi3BAfQqDdPCDgXw+bl4Rv0wmslqVlov2xooo6UYzIwUeME/4a4F5/
GXw8OheOUE1Y3AQh0Kexx5Yq+x7W7Pt99ue4SScRglU=
`protect END_PROTECTED
