`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWhgvMAgRy6VJMKhM3qcIYCvj/GYBL9Ra+xAvTk0y/C3NMHdSWKrM+VDGotLVxV1
+opdQ8TNsA4aS5R1ion9hPNpS2ybGc6/MSdd9PTT2WZQiSvJsa9zmtTYsw21Ha9E
5/sHcuGzWi/mjZK34RAdSGG6jyeCsEvIPMTByujgkMgdprv+HAAJvPegAISSpm77
WvHnMwWD1grTgMVPEsoJZ0oBUUwOOwYBUUuxMufz3rR030G8SJCNrOe3Ox5rsF1c
PhevBdv5OkMcIQVfDry9Y9Hk65xqg6Q2TleOqJmibJAfeCQhOuntE5RHajisLExA
JD4lrD6Hsi26Uae7LNlAMpC1aeHsO3QbExx9U5XQnwc8Nwp19/3dxp5tVlulMdqp
T7daRa8kCZGKF+SF87NmhJdkQMGZgRpxQAwh4neTSgfQ5Mcn4mndbDyH6Npakp9Y
UMgXdUNJhjxVvrold0T5i3HfgkWjUrfcZCwtHqVpIAMbisXPW+m+loWXdGZFSbs1
yaLGuG9VDidd2xInhpcucVrtUuUiwoo6/8XjibHIdAXaH+N5utIfP3mJFUsdaHrQ
cwYucKO7MKq4LKXn3rjGXn4xVRwpl6Vjufv6WV2EQsIrvkYwb0P+TRowmISxsFci
7SrlTfjVrO2I7hHk6IfiLCxq+RJ/d6TqQ5swXO4bO8phx7nI7x3gJWtkFdXKTV22
sGjl9PPLbUTyEjnwM2wYlxoqmKReJsf2NE1qJsBx2zia+1ahExZKmgDaxQS9+eYs
iFS7gmKh7h/XJUh8rNE8GWFJ0NbJJiFN46ywplI/sWzZY8u20QtDtlpH4p3our0B
JyMx9ymg0zRgOjEYkAOxF9RGH+vTXCFsb7niaGqhtu0pjcU4mcxMku7sbngtQfeP
D4IQJsnvoOc145049szq5uugo5HIs4NsJIiBlwoIvY3j/Fh2AzixrUbbCO6q2M02
4i/BB5JD0ZFoG+8bvgoHeDRFLAv5w4ufpQDRMuhhZ6GPDvkiGpEw2eg/3h6FAiJf
3z5jGv4FsxN7j3Vj7Hh0L2QBErKx7tBt5Wi6MeDu34rT2X4/teMl0qGmylK4Puvj
X4l0TUCsSZqmCz1Tk4LCxIyRgQsir1mSmtlngYFylZreJCppNNDaJ6kG74eNklfB
56QpsJpx+LYpJrNNW55M7d3ppctWUXroMIr+88A0SGHBYhyRYg/0oIDAYx5+Vohi
ph19LcDI4/zNcaOjKuUfhIRyTC+vJefDUiOGqdTlmu/zQ4Ftufa627RYssBfRzYg
`protect END_PROTECTED
