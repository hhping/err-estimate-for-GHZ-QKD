`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hE04xW/XN71xHW7dOvCyxtNba61AmbpO74SLTDU/0BLxfbDjPNI44XHpAD7MDSq3
C1IQDgM4YPveRZ4cDx1Yl52kPEgFQ/G8SoHkWMTx6EocIx/er3duLzfgEnJfdM0+
VAMvJ9s3x81Vui8/dz+WPysIlYc1ZZBNr0msyiQiUTw5mIbHbakZTara8ETHFtch
ZRuKsMduQMfHKWhk/HoGZSJLWbwz3DXC8YSHIKrgK2nhPZPf7jPN7uWJDWPIFrRy
3UqB9cZ65SQCMuJyxcCkwRQILxbUsZQIHn0ZXNf2zrXZypicELfrNG7utbARmes8
gjhFSjTxnOZIe+kYxPoJIXjQ/rioobQjR5hXPGyA+Iuc03w9RLhMpX4Bh4OP7LN2
f5EVaS0KDlGyJuOmqxsfub237OJSe4IBHhMUhPnEz+pyocbaZK8NGGwXo9aG+krK
OzmcjhGEUh6Tebh3uB7TEWJ8M+7+0U+FtirEes8Y+Yon3J4vUXKRbOmUMsWA3eIw
ikqtkrDreWIYkTepSCRTlZJMpCl6WH0KFXI0HzvX+z1M5kCYfP85c0iFunWMFhyt
UMu1YQi6HFxSosLAxE8jA74Fm/QeJHuqj9o7VlhRoX6y+yTc8l8/v1A8g2Gnk7lx
XEZ47N1G3TF44by/FaLrGairqe7FwIq+dle1vO2F9dzMRgCOcvsSxfYcGaoRbGwP
04tXR4zDTXRFNPwzijeH7pd6tmyapEgaxBg49goD51w3R9rz8sYVptymocqErkWr
nC1otSlzVnFQa+It8zQzp5D+RRTADKQeyW5CUvGF7I2pgCZRVvUyb8KtdVeIY1Pb
u1GonkvRZIxg1w0i8zEPt5XVB4qEb/heZyGdN7ZE7PubwhL0zHzjXLETqVE4DGpF
IfZxHA45IDbNAkK2yb+HwazxpoHzyUmYAYqPplDS08Kvma5/d5LZCHDRuyHL/l2E
WsHVBrgWptpkRF5o7vAjIB13NIZ0//GCkKET8tqn+ho=
`protect END_PROTECTED
