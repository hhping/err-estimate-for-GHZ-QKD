`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhBSjFwb5shGumPw1KeiMlRFDN4zpzMZ8/9weAPYAqRXZzboD365IL3xjBKXn1rO
Q65X/f9LVTFSP+8EOnk4wTu95i8Si/zyfKW/o8PlCBq6rWazy/HM2KM/1CSVs6ut
Mp+Z9kImNSgHzW93WExu5Hj6Tw6O9oT5ywhZhr9BE3EpGHC793YbV+X0w58fc4jS
+kHtYALzKROuNosCW7aDEKugQ2HRLgk9ModZF30Ksm7MOaquWiuuev/f42RBwf/o
eqZkR0Q87RLD0yX6sw1+R86mdm1Tyq3lAMWb1+vPttcfZjB0QrHabCqx6fcFv/Vx
JjjmZhPjvzuhUam8GCYvsl8zuHBHFLG5nt0FcI9cHGM1QRG0NPBn0zmk/cHplto7
sIDZ7a6QqCL4hS8uL/Vi9EjJztitT2UOou68JNMBg0Pq/Z2uWMIKHiJ8ObiLVctl
pQvi120d2s4BSlFBePNU29d+mIalxBL6cz/NAX59Jh2TST6glc4tm7J48IG2foQs
yZM2ePw70lND+RoRzE7fGsJa2dK/0pfWNRnMPcXufOF1M7+OJeKVzQeSvhoyVUqM
/v3klii6d6SJrlBANak8IA7goHiurVMcxmg3Mb0frzl8G0Hz7RwPglS0N/4fMmhG
wD9rZa+onQ9mBGzRQscNH46oejC0rfXhJ6iN3YNHbKodDkOEPpI7m4gqV5Vs+jRT
LH4eh/WrNy6Am+Bghpf4jZ1+UmZXFQACHLxX6TYswJdBw/VZL1yMId+Cd+rgvCh8
356NKn1L3FE0n5FAxSsub51X4Rph2Rk2nmzqgzrHO6bcd88fzjwlum+wjhj+3GTU
mv0VzT1G3Z1w+CAp3vHGOcZ98fh4Z4Vey8lxlCoU3b21SM0N4r7q2b1ORLqZN4aD
L5d8Cm8/UnO25AepWLhL4+rfXH6G5UbI59nMALN/I/06KShTcFxN6reFFK/l88ht
ePOnwA4EA03Ei97qoBtGV2WblmjWcGenlyXedpsTN6D4iqUwtsw5MbXDL4Qk6CNg
yrXMyHUiZbm+g/eQp/HDjFQiqRdQgQMNhAlBwgfygS2H/dJsQ3/BjzQ+IP1Cjan2
EfWhOLJ7Iz0wo/cu4SMYdEIR/bWrQuMfgMgCZdcKBPDArOir4RBk0f2FPLoHmfHD
i3c3fvel/ujT8VP9n+nqxRRaDg26hIHJ49OgzI8Ulh2z7XrFh1x3ZyhXcHygdI7L
x0z2THfV7QkIIQQiKIoBH+CRhHkUmlrK3+SdPqtYRwktYeAHCOUtSUsHn/a2G06x
G/1m5e0QJUmclU2T5kgcQ+SDcn29b0K916nOjZ/QctK1u4UrCz0IZEeKH/6LqS3H
pXYgGx6k9wydEiRVpI5dqAvqeTb0nAVz4EcOI2XZ13ZEZIpKvPkk+UkQ7bfnVKOZ
yA0s2xjIh9kbOTh3Npnr+rOz4hJD+G23BR5vfoVDnzXnjOAx1m9nqYY/YyFaenIs
WKFTQcxbsX+NSRQ0ez3PRul7yyNDhdsY69TU1DG5Kc4MMH+qfBJkDPAYaW35Pf+t
m950VCZ7XDUJIwnEuLZDoivnTbvytvosK7y07JWN/F/W/580l/VFl3rGOH3s8Lhw
MrLzxLUr+JxrH3qovPs5sCNMYOTSwE3bVB7fH8AfQQQolMFG0QFAuAPvRFE6wDI9
edttqF7pP7lQK++rDyJrPz6HrEyyDvf0JPd94eAIpQ1CZKDt5XjKuR0ah8g9Ml9y
KF7rMju/n94U0Sp7cKzoymt1deVKUc8Pn97zLr5aNo7QtMrk3NQ1DhOq9ixQ9/sa
a4XGWD6lEelYd0QM/TNw2Bl9crmZ6GpU2nNfX4oOvAr9gxn1A8CoZ4se7W+GCoMc
0qFdyGP8r9wIw1Xzkn0UTy66V2LqW80vk90D3ShFCXV2Q6cg/KtOqX6ccG2ZubR2
z4sJsbz4J/dTkHd6lu1TdqswQwBbtCS+bAt1Nm2SCGRGELU7rN6mnrIPM3nXZ41r
xVjC/WX1+YcU22iishkkAWCXpkLtB7gGp28gpXNQFmGTFtph3Gl44HtqfSBIvcSC
qNGn4M8fBlnJru5/MJCkkz3LkxIWNe/mqoQy5Qbna445u70zIz7owT6becTa6/i5
Pzj/8sh0APuprA72C982iQDYEkBRciAKhM/sYMk6Ocy0rcqCyLODa5ljob0XzljA
cZBciwgRUxYWkZWJTjAXYxj4UhRkwFsnqHXfZGGO8L5bzgNL+QHufl/Jx4ZaOGG+
Q9dXwxxnhS66nETOZ7VjOg4RCv2EgI81LV4Ox5dfTV3gnjhcY54o36waph1w3M0D
u9W0llIkWS9e/bddHkoppgyaJcJvHiiw45tLgSBX/sribKdCD6hLsmSvnxaMA8NF
vcuRr1BVO+Yv9hQS0XXbPlePaGJWrvt1+BHvKmx6gs1NFrdM1qO1c4Gp+YiJoBW8
ocxhcGcVSkfRhfmRWODw1DuLmZVO6Ex/ubPLjoLw49K23e2oHQ6xj55PWIJVRa77
6BQ/YhOk0CBtF4XIfaS/YVyGA3G+3f9YLvCoe0K1G8YAhme5LNJvwi3Vr/nQewx8
Bka5VLI4B02pC/6DaBC4VYkG4H+1DO/8/nUVymZc1G18rYDpQT+4PKhD1ngLb0U/
FEgYAHOaAxzhJTPUdSz4DT7Jx/gDsdWQ8TghgUXvZdPvLzuXcyXkW7rZR3DQsXAg
wO7pjybYLnEdY3C7r5UJZJDeOQsdFyrSEGr8Al2ziHrcc0RYKcNbhbL55xklg1Pz
e91y7xN2u3NRAWANLpG6YxMgp0mx3vsVyLi3k3IZHgumgWnqa8y2hCPNbQWc6w7Y
1jTuxulR5eFRupUL3yns7tx2qyyCMMb8re0sQs9ev8b1D8i+f0s8/BNdSuHSTekx
BqGwqdnJKA7rCafzhAFBmrsFWy/7A7N1ShlDGwdGWOjyAsNFXYH/1nZ1AaCuUv13
/jKWF+l0ZmVBqKp0UqhuplXKdAaKefnhIPfTi6oDanOWuEPI00kTp0f7XatSNDwB
yOuROZvTvciHleUFkhWEN7GHjp9HT81xDjr6uNPqCfMBMZDPn/V3dsl5MnO+XnVq
ffNpYU151XHYn9m+FGcqqKwSIoQJ0hlW5ElBl+G2UKW4tVLintim2SL6yzegghe8
BJM2lt42SW0mWNrfCFev62qgAhJPxlhDboehvm3EKbh3aEshVSnlof780Oje8uB4
bEj865kw8foxdNsuBf4UeDwZGsOekia0bjjvjh6rnUF5UAC5oRZ8ZXwZk7ZRmbQl
/sMt2FkaDBAUY6lcfWB6+kD5q5MR+Y4QDsgNlwyCD54yb+G86OtrSTppX22sIEuC
5f9xPpoglnMVq3GlHu6EXdPs36Gy40Rp7bvbh6zkjLLWHdjmge5wJVAHUNPqc7JD
m2bogSkaNdPC5Ynex5bgig16OqBhU07VKvEbl6Zw6jGlwM8MhdZZyybLZ3bNMza8
+k3G4tRn3dMCpbSdwazO9czJiof+/jGoujHiQeSS5EjLoD4pd8AZtqW6uCPRlbcf
HoqNHFmgIaVGyRibzj8icEkK1XlCnUp2/CegVMsdjnnKXhwJCDSNwExsDrO1LR8F
PShMSISxT5xO8lI4elh5XeTWr9K1uD+qFPXu1A0rq9lggRAtaE2O2QNYI2SR+ojp
6V9LEoC+XZN9Pb6viII/P5xUhycCGE1tTl1Mo+yHFJPkssyOx3mGfoW3sf+g2aV2
v92JLbhzp0hMqqL6zdrI5qH2XDhrPYITAlMtzLtKjiTUxv6K/g3IDLc2QeGtO7Fy
5N3HDaUslaRECw6N7gYrL19nO9vPoS7aE4DubXhSt/fInxH0M1ucNh5c9NMnNjc/
kHY8c0buzblzXG9LpfscXEUjTZ7Nms0yoODstIWd3ClGkIZawqCm5U/SHzs/yoDp
xq1vKc2SFmF6SIwZH/kZsqIGZnvAR3PwB2SWDJmwxjk=
`protect END_PROTECTED
