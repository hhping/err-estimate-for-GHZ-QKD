`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1WOoMCltyTvhx+HeXJvNg/dr4AzlP+Uwbiq0LDYhCxYzfWMi+6RLzLBhMHr+Ures
+kojcfFp8fnR1BNHSNyLvZjJGI5gq7ITcquVfOfe1u7fmhujtzGp00LJs7rmU0EN
USAcX8sFr0RnHyKtN9M/+XP54GkEyM3wKZdlI0CSJ/Tq9EU+MVOtELEBytJAu/UC
EhzGvd0Ugrq+mAbbeyMwzii7U+5NccSpduQL9LtXk+TcCN0KlJr4XwE7qZ1PrEgq
7kpODoIjE5vuMEugBBat43afBXVINiYIF7Ay2Bk9HrDmSXJ/8NL7H0zfoPWRmL/V
ON8mSddAttIXoA63kcxg+2xffIWNTQ9fEEu4vzsIsc4=
`protect END_PROTECTED
