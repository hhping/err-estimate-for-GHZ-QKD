`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LsbzHrnpTgP1S32brvL9yssOMMX7CIPHwAMBlmTZsCIRK3h+Py+kCMSjMQhbv32D
f0no5oI5jj61FRUhbxYpDrG1bzOB7mgDaGtU+LHGTHgUGtA+ltpxYTiceT8+c6WJ
womTPaL/FaKXz7Ltw4nMHIA0fXxkmBz3m0WV+I+k3oJ3D6rYJS/9lUGm+psjSBfj
XiwdWdv84WdRZwkuT2WU29kH/y09qJVxXVG9PV+/RL82ihoaNJpc4H5JX7kGwSM5
rJZq3isg7c40c+39tDDxXB8Wg69R/5+3xXRJNjIGKxyqn5biH1c1jjbtktjCizYa
acZ7pCmzWoP21NVM4j15KzRy8C+QJJuvZN5GaXrXwmHbA2uVmkyKH9rHhsM8VgVC
uUSOkTfRNFAe4Ryt3tSDDLP3YQcAnWH7wYY6cW6ikeNC93arJ5fYstvV9Y5O3EaA
pP3fOtdF7sWDxNwsIf9kwoISOXipdGzZOqjmMWWXpcinHwJWI8MpWxV+Hgkg48Ln
IoERZg+ltac36VHawGdweSbssXcXsLGojYy+bG2MtpDWE+tyCrUFsCQdGTLRJyJL
Vr6VKqswwmMuvmnsw/GpwoFL5kiMV9TJDlq/VOY7oFAt57zsnpQg52oQ2ahC9SJi
zo02akRUZjQCMfH1LbkeqBo9jwbfXgdGJnNaMsiBOR3nvdva6ywe4lTGI51YV44e
oOhBG/OSvrmRZ3CjVp9d2Lbb4LZj/+ir0yNpVHw+kCwWg6Nsm1lJZ8h3a0lRJ54O
yuOEPVeOSZg18nKz/syiDu2Yl/6DrgHsHynz9yu1smZnfO/wTZ5JBEnEO0AUfXkd
GzbTRmij4ngmN1ZQJZ6LqNuv6u0B3KAH/bRnZ1AYvIFfGkyKPkns7epNffwnDHtX
7j/ClQ5ujGz7T1/DKPyanYHYhI+gx5FQnwB57+4DGi8A7cBv+25pXMgoB/iDbfcb
i5LdeoBQuTqcOwQfrROES+xwQ2omSFLRFFpCrDIf0I1atpPG+oC33KAVdOGldElW
XLQ4YHYbvxF9RrieaTMJARqunzcvM5m7c0kOEEPFXy+0oTa6KsFJTZ2/yU3rwC0X
7AwbMAKPN+7yQCJImY5VFRMKmw20P/brEGZFhZ3TlwSdvr6oOUISTS1ByTI8ECTs
grEJ3NG17F9Qk7eeEbeO/okGceVHTK5CWmMdxo6JO0WfPk/+9UOMtq+QmNOYgETa
A1uulTJpgyOSQ+VOgaTttk38xzKwlEgDED72eCHWnviSsXptdsTRc9BV79R985FA
vFNG9GHxhx8jV2QGlbpASEHA5X5HxYbx5Pn0d3P0JXtYVoxR83hXaF+RJUuSoPwC
qfQSGAi0FLOZVpjK+yeyUktLgLeTLnM6FPVXDVRhQfZHfU1nTBxgcSi2LX+MFx7x
wpIwdTggMJ61mAc6pUuxbCehiHNSjhL9qhR4NMFAVCWaGDD4HwqncvPVY9HH8d2x
YdBvxXndtPUqHHzdbROhY9ozP+CX6ZEnv7NCJLK5Btx/QHAZsSRT9nBx7CIaBtdU
qFuMtv2BsKQrRerh17Ss9pGftFjNI4OZXEXLc3JNS7ku9oh8U9JQA73Qw5daUg2y
ZVq4NJ4l7K2Fytj98u9Pw/qJcszFRIg+/foYpEfBIc5/Xw80DUlWd7g9Gt4LuNpY
`protect END_PROTECTED
