`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+DB1mlUxKDUjivZEq+f7ypY/iwCq7qoggeoISUmaybpPGwDIbFlFXQ+uahl23Lx
7PZccFj2BV6yA6SL7mrC5Ax3FMG3mqRdDDQABwVmEn3pCKtkns79a9ZyYFKzAvEL
A4c5BCJiL1BaeZEIvkE6bU09OYwPcBrqS2wu/bu2g4LWN6n+i7z2+09xWrtzcY7h
FmKCL2eXyhyzbbaWuopmtuLhp9Ao6Dgue75ddLWUHhSRKY+itNg2ZuSMbEV8H2nk
KCrNujkgguLbs8RHHO+ZDeQmiLtsCeP+0MhazuZc4zKFJezroF5Jl719LC91Cyz+
7AuvDz3IPSYRxbpdRv7GH7wCZUql67H9WU9TbrJOTqDvh5D33HI1Qps/YsAG/ba+
KeODV045sPAE5fhbH4SUDaz8sN4pYnn76hDICnOgvMso6bIPugkwKk0bEUR86aRR
Fg4fKFEs8ydVAoUylyY6jiMyJN9Ok4iyzEcGZBPiDwKkOE9HCEXzfGAZRYiB00Z8
T01EeyOgHjVrw9DCPBsrF/ao4D3cLHbbJYiIa/bnhvezrP8QdHxeqrvLu3cbCFaH
KWuuI1CklGHIRjQV8ai6TIqesZx3J+sxD+sOIJVxVjoU6Qsi8pU9y92JjYlzJmXQ
QhvgKvVSy1E9JXm+37QpkCE/xNBVTqg0ix7/jUZM7JtQbekV5c8cfdwI8O1kOxGi
4s0yLh1wZSVyYBCwjtEkvl5Y1yucwuyk5RBH33SVRS1dQ3KheUS+1NEu+GZbDwZG
tIwuVCDhdQ3SkG/aJSlynGZRe5ulBQ+0hWX6xE0qMNva+J4eoo7TPoHZ6/BvypBO
ke2ti6JHwqcDx1+BP/gulT27nugYaX84ay31aVoJhWy8RYnNkhj29BgDeL3TqKIy
Xlz/E9+TAuFSqCff50VXaDuETi/jrmn1ShYe1NEm27cQZdjd7vnQCDdLDU8ef6F7
xbM3CauIGNLozOxut8n9sBSVBXGPj6ESH3Bybxg7Ajp6EbV7aYFVA9sRfgj36qqf
L5N8/pFH/Mpd2uO0JpyCdBThPaRe2+/uud/sL7GZ8AWj+8MN2hcslMdIbRFR4PZ4
ETuC/npNyeBApnGY6RNQO5gveLYdNkBmTIG/PXj8noBGYhHKyEUBvJ6cUsdwt+v+
qIKYAD8R9gznH6ZvT1guAGYiDKomQCbnCyv5H6d84RvoShSqks/zCtINTitgqxRZ
SollUVBGbkifMA09VgaRXDWbOcIhCK2+pU1d47AjQOaf7YC1p+P4t63ck7APhPeb
y4hjJAZbIqdWUKV6M+A9M2DLANJhJKyCdxS59SZQlpeQRvCwASOj2pfnCFiNwJPG
`protect END_PROTECTED
