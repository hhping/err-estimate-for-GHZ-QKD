`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mgvXpopcSxuM2d/ZzG58ALjwte3YWKYU22nitXFcYUeI6/Y5VnqhWiazkgOiY1iN
jlM6+85Apcmmy0HiS1TNH/bMEoD4uBKSfVIxuQmhPUVh9reOikfq7TtsniBSxX9w
Ylae5L85ZZpic/bte9jdB2RGbLn+yfSEk/s00lsKE+QykG80ISKYG4mc8zXOdNSU
3faH3182OWh19S1cfOf9MT6YY16gcErAwwsdXBxCmyDsV2kbxmSqm6RXXGuX97Sn
sdsj1SXrFwH7VPFdkiFHco215Dzvj9Kv+gRHeooBvZbP+Za4faR3+Jvp5JfHtOi5
DGqkpOWxvi3bxoc5naozabC0hbEUNXQVuaWuUCXfMvN2qtxLVcQOOsufoifvvm9Y
g5WfhT7Z8lZEhAwAAVEXywGbLSp9t9jKQ1pv0pnxuKHqzwsO74DCRXk2ebN7K6b8
kyybbhxWQ8PNEYGDKc8Xo2DTZZ1m/xZeqTOOS05KxqhWDz4g7RJvSd4HoWQ+QOhi
/YNuYhG+t4SEWgUoiwFrrQEoi9GHEcfC6Xt5Q4vS+9ch3RLvj1GT1LyzOjait8zk
4D+5DtjbE++xlFH9ghvTFW13HUqSwJ9yFapyrSJDXzCB3AJnCys2sIe1oCEGAJX7
z9Y3+nlKVhhGKR1ZUujrf3HH5QBpAOKol62i3zXIRadQFJNxSyL14cAlcZLz2iVk
XgaHjTszVa59oBfFh7Iv/6GFEnEVJpx3xYLU6TVoHy101BdT0E86Yoxocchj+jpg
3R2UWT9bIx7mVBRWP0+cfevgju3pCTEuNhQZLfA8KVSbjjrqlQPCTp4LfjvmwpQs
ePQPeBYLYzfqOM3ALGpWV0f67b7mCJ96wBpzSgh2C2FJRaBcG52JgI4brKcU3VyG
eLs5CicEHwmRCBQTN1smhiSqicXyHKRN2Wmkpx8cBkQ7ZshgESIsaqq8qw0tsB/U
h6L/FYhe0L0mEuc8dvwgsiYwvnZz96r/JPMncep/RtBJ5mPtJedpC0w+WEIiynWW
0WCKTFcjNKVFe7ibJxXrC19WM4k828caQOl4xKc4tofQYu+RM9IkEV10sRHjg9pY
I2lXYSID1rS18g9Uo6+nppzukXzCRt2DYq3ir71ypmk93wW9eQxeTBiE/mMOCX5J
GUFs0dg5CBjnINpQGcPbK7ZQPmqVGXMMuCnwSt7M33GGx5E4JEWnUpuGrVR6AN+i
pfs5Gz2WXj+VTuJt43yElERBesMoL3ImiraM3foh9ismburJY+4NH0LZrBSkEdfo
kdpGoWSxLq/OyzPgAsc4YYaoHRUHtskw/MQxXcPuqhWfwMHEaHR3L5r28ZZ44Sx8
4WrLD1PSUR6V7lO4SrNMpTAc7Dzr36UgW2/KqZ4OROJR9iHj6QuZOhYdY10ugTly
PSoLN1hF24+vG0tpBY2LWmdZA3VsosSc5a2EUs6PA6KYCcbujzJjtOCPhjZOcGoc
TG6RjYCZlhS7hUb5aKEq/KrDU4pVXDxeRqIPs7CApWF3kLa9iRpWj1+PjXM7wAja
YiWJAtXpxPo2ow+AIPPKWJqSz3H1vSN51PHJ+uBhvSbdFqtdDGiRKaS7h+VXA/TM
ufLQMHS9YglFlK1w2K0KNhV7MX2BDa3z95JdSgB6yLPMyVmkLtVsr4RE5Gs53+6A
JP0AB1jAsGUV+8W/S1+fanPR3Sqew9G7SDgpVqnM4DjPRkX3HLzBmCXKSCIB0Q07
X3orafDO76Q2ph5UdHR8ytLsn3NWZYDHAac5MFMAGYDxq8GCuazN7GJdxzp7sX8U
QedNpR5ro+nMZiAQJHCVTqUHSKGQov52QOrPxezgpgF9S2FzfsMscVWagsZmmPZ0
mxqWmM7vLV7mq5N/rode6dAs3sJI2v1gEAgNVLfYAXNwfrJN7VHjw5u8MWpxgQLA
0tjtTbTfKns8k0k+0m7KxigUaWN+DDOw1cV6T/iByrJmswUmfBJkjqBdpL0/L3MI
AEi3I3Qm8PGkgiVFk17f4PYpvxX7QU+LO9ffSgDzMq/yq9CZ1CBrk/fBHILT9QEC
h567mzkgPGU7yQqkIF1ynWgohK5T6y1uP60siudHsiS55QXHaq8HDt2CQQgB+6OV
HdYrJUbS9UDATA/vlgcOdQ66wUtQj+JMyJQgnD6II9oGEZgOfPzbYXltTlcT/Bwc
TG3M4NArpce8o5X9gwt9v1TsGDQ0W9T2CTh9HYZ03zDmHiUqE5QQSF4WkqV7oP8e
hLNd+oCJ9Jq6+dUN8sDhxlqZ6D9QME9cTBjVO4lw/ebCqyWwNzsU2fcCjDNmznti
h8teUI98i2l6yTIqPP0rUlcLMqVSYyz54x7+aDhosWapBGUtwYoTd+fHDcrAa17p
PmQn9Nhu2Uuy/BiYB053vrj28yIolG4gOUi1TwROCXyRTwmyLEJfLkl0i72zAl/k
NBFxh3fQU/Prai1cjHuE1Ng0mEXvmiNLPca+3uHzQi7Bk5+0e+mWWxc10tw+X6na
kWuXFZq0+A/c7QPdCtjj0HPZJ5Jc8OB+3cTr3Wg0zzuvE4dpgpbnSPxZWoMyz2SV
Rot/QO5m59IWQPx59xJHVQuhUL4ltS1ILZxUHdBSOwZ9zEjqHDCs5k2NovxACU5a
/tQovZarrE5g+wc3z9ApGL32UuOABK/bF7RxwRqWbJrDwaq5xXGMHlx49w81emqU
WK5Rjpe6jXDw5/pG4VpuKp2xtMttLQI3/Ir0gbP/3laILRrHIQLkH8MtlUMu/omH
+dNziSymi85wczxY1YmrJA2zep6i2GWQV/sbUL3sgJJ6PUVgVpbn0awFmCtNwBcR
ULToQrhNDfQ7hyDpzf6kJQrURWsjKi0+FEoEiDYCF9B0udjes/P/z7uHFLkuEptS
r+38dAwL9tPKdtpDZpLr9a4UsBVl0uL61RG/1PJY+blaKSCUWCmSHR6vRCFADPog
LWjc/PVrDX7aNoWZPPDvui2kduy626A07AV8VqQOYRH8v7WGUQWzx3PibLYNr8Rr
VUju2XIlDMTrH5unw6NYkoYFSeF58vOk3NzjbAmCZsEZPS3TL/++hjbgj1B1LcMd
bp/Leo6baZ101TLpmMZsu8NrvuYjzE5MNwTTmBWUvHEd/BhkngcPo+JsdY2u8yr4
JPOjWITeNzglSnXDl5m9cKdkviBVk9L0DETTighrlkL/lBqmrFMZOOBr3wWNdi5y
Tuad3fxMI9FSGzWg872XBywjVjAwtgWrqFnuT+CdxiUpll0XA2/bNvKGbVvFc2Bh
uol1hM4rRgzFhvUxwT2CV6euYzY2qnTEyehT5bep7uuo5RScoMATXNQN7fu7Mx/I
6StxNvYu56Yd67WOyAgw0TG+3LjLbMkDwBIxX4OIzX1I6Fu0u+0cvsPvRGGidSNI
y3qgZBwptpJuWf2gA3IfjGgCJaZjPAmBWRrRjwB8PYk9mbMt05linxIwdTkJdFwt
YjjcxCCzfa/XjrRhyUD6naLT2Pwm/LJ00defbWsh3eYL125Kh5khvh85hu1pvCki
ltTSbsRcu4ttdhMoplbTWmT8ibR5BG9XAvae0I11/VHqcCxR4EeCOxLQ9zENiZ7L
Ka8wowUEy7pINy3gxEEqxqjZLSfvD2MQ4k9/i7PsGeebj67QktI3TycYhiKNEoVA
CwNedOUY3iMBf07U8Yg/yQHmZiJpSP57y0Ae3WdfxHWiMdh9+iDz7O7qmiw8F5eW
1mrtjwWMGb20tkhWj71zOONlaWbUzeqtadDjhng5CfWEtCZ70BW4+uoZB3oZ7ngt
ZGKf2Z/aEsxOs7Rq3pbnzwzXmpFYnYW/wDTwSnRf1F38AFDE4D70TH+1MuRtij3j
rlScMQHMiUAmZ8bbFzM2e6DxhLXhGNsZwpsAo+ePESXCXIcuAnXxKaqsg3ZhVp9h
GvBkVFLGpJYk03xrjLjfW6ETzNen2OBbCoNfHMGX1B7aQ60voPo+0BekZDmiJL+N
gGmdAQ6DrF+6Am7z0b9kQNGTZ+YtrXNf1MJfMaam8RBmUJ7FquHt9ayXD2lVeoYF
9083S8KAQs9xHnPGj+AtYSJczlaeYXA56eLK24Qvy0+hX1i64Cnh1WgV4yUl3BCs
huCBy8ueDPP9MOvI95bLY2KF3cOst6VMJrW164DgOiGcE9ujR/RzJd/+HX2CDYvy
Xxt0ZCse2XpwZp9SHmeQo1qnO5mWrt6zfNGLTuvLiWNQZCowJ22+VjviJ4ammTRt
cdPHaikQEpW9CFzMlnyTgclRJQT1HT8Cbc7HzI0ABBK1qOZ+dvmzBqa4P4XXEv1u
+WapQOM1+Q/0RCEkfAS9jSZpEONY1hOT2dRPaLQ6/DSO9kjYK1f4ExHYsk3g5/kQ
GPUQ74pXLNqHwQCjgkI3jfsWPDudQ+0hRZK9CdNhl8LTXuIWn5eGLBq1URi5vdNi
+3Ptb4atx56qXagGh6lrHKc/a5ounJWh8B/kTpuyo+V7MdU127rkmYAtPkIu/ASr
CmgCpO0lO6ntvCvTK1hjHyvKtGA1hr4ObzMBdp9HFKV91qRmz4UjjpRvgQOhnxkv
o/LNAtk0pGlG9okkdJtCE/1EuNxeJlyZQXc9ZNv5gC8FELRAGevZe8t9DMWlYrsZ
AZaINzIBGTn1/3AyNAitcw3MzKKMH9sygyGj5POc0LA4u/CNqZRWijrszhJYbWm8
skpGuWXIGqBgj89Y3CF6clKdQR5jb1W73kNaIkdZc3JmegaA8gKqzuA2wHHLZVGp
pkw+v4/Na+UsNxpaO/VvGzX1TncEl7lLPk3UZ0RQhKsARSJK6eScySqChoZY2ZPP
hOt3Ch/ykzKYcB7YsTmPx9QTfieCnJbtZIS1H70+CrPumvbCuXYe0lWoOlrFcbBN
3RsoUXVlHGobM2f++e5Rn8BoiQ2R9vSLSOBb19ZpUwOW47dF2KOBeC03BRLxpAi5
4/oC2msazChZB6mB5LVzrZbb0bG5gR/l4ZzHFGHrkdrptCEupZX/O3vl7j1b8HeR
BvyfzLo2oR//XiwNLif+p/jGzfvJftiHU632HGqjQ18RaHiF8H+NWlvoWzOeWS4Y
AagTD2/Ty2/Deo0ZkBcpnzi5CZty+Hmx98L+1LfL1sermWsAYtKGAKM7T8lsFEKD
bA/3pmdVaiFgA2WCVZQgRlByE04jt71mxV6JyM954msUDZ4qNPOKQg6yAKzcUW2Q
tsioV/47PF1oyOceW2W966TRRN0aoADtKLEMMKaCXSzZ3br45DMYI1Fyo1p+P1YX
tTlvFhKSG4O3UKKUlTx87UfDRg/KZJ9Y/BOZcYN7KBsF6a0NiweOYv00yKQMlnv6
ywp5BqDiC6obnXKpor6CUYt1QM7p+3FRT31v42+ZAZVVfWQjGbQrFGlOx6se3PZx
YZWACh8fpBaQsyLQ3SViRnKum3N0jq5HMXtRoOeH5MOyXyLnxb90qDuLLQUVehgu
4ZdPcJeJZEGfTfo0ad3Agj6y981dZbksJLJWK70MaMOqmT4gWlmhCKXmWaNgEPHA
LtsulFoZV1nt3hxvfe37oVOzZMc+gfnyV3o/7HMBDioA9YQSE5eplXUXuEmbIdNp
SYENgWAweL7oTFBX1XJYI9qtFRAHPhVpYi34JpZabP6ZXAcFRrW2JFk5jcOEhJKn
qbe7TIFZ7Aoq0CurbE8bUFfpYldqrkYeM7okg4GW+211RjL4TDkdpRIaKx0ZOX02
V9KT34HGN/BGKbLyf9tWB30bG+69QPc3gLCo9VkXrVsT53LjL9Um1XPcjT+5c6nR
EZQ5OIAwE3I0iNaJoJ5yl+6DLEg/DN22Go0nfjOXUlr/bbAkqjwxGpSOWvnnfBUA
ndYvrSsNWnKnfKlGSLtVoRt42NNPJLxThl7S0AoCc0RwA73C3m+N6FIkZ2+xF75P
sRQTpHCQL/k8L0Oon0OVkt7huO/7TNfVPZyVNm6HgtI31eFg8aB4Dij1exQwuIar
c2UaMnvyLLzrVpf7oGSxQHyBMTN+aJqvUryb+LV3458A48uEd97BOd3khP6ro2IT
oB4JSChGGAiYu7uADzyAEArENbFA4/QiFWoEaI6xdB73ErX4xAGjJJKTt1/yQUmn
DiLfSK2h+6CWmh2Osyt3SyomUNpKwW3/nU9O9uwcIqKqdNvWfElajW+83XaSw3EJ
1czXHJiXsfmrsHhLLZ8O9fO0T4S1TGmtsKDvZXKTyi+H+sY9NB/lW6IPpPNyOSmt
U0g5NoBYv7EMzNVWuuceFDBfabu871nIJ4EdnRlzk5Nq/y1I33qdDlZw3Ld77YvW
pEXzZy6WgOVfMh0BgiWj4m80J3QttlFUl7TLOG9qbt153CaR3MK7EoBzVQE9BSOa
oSE7S7LH40Gmdur4OJ60MVdDOFJMxl4vhToFuvLFGtL65+E4cH0L5dljnxF4nHt4
BH0VSiw5+K+HvfXs3j3qFAmEnLCfvItX8vLr80XG8FHxYsN+m1SJwsK4FloCZbHX
scAuAdJsrtyWDkObqLJBQdvtwyDYb1eSM/YV6LWNSpXjY/N06vipfLqGMt1/n068
4LGAAPjSemklfYVJVCJIgmLdo+WWGBsgIfbsJ2lQbu1Ob/V/i8SsQKaSmLdhnwrJ
s2ugdDlMesxixs6BTbZkjpLFr1NABB6/47mO6JoYbnEC7P7rEWp7vRslBkiAHgS0
FJkevCX4JDoHT1aWwsrmY+Dwr0xzYTv9FRUko6b8fBlttwJyr+DK4K4niIHCNVSH
jz5Q+7BpY8k1kyK76q1BSYlZKwC7wHbAvUtUi6laPc3zdKm71VkxWQr6iGIAVtgU
qsTixkNiIVuiiIros41FDMAR9xaNgi3DegT9rJLQuQ1x9FbJach+FV8dGarx/FIl
TXLYZ1oglejwODngqOTk8axPY4fy2zHQih1/YNUAN4JAx9y5dpnfhoRNTpnwo0CJ
CGRks9kAH+a1N7+AIzRHe/VMlK4OxpCnWeWlPfWzw601LyQKNpXRU9Mtq9qL57hH
VdU0I43ui/y9DoJS2R5HNAIx3L/I8qvdnkQT4io2S4hgL3+rT/gDbx6CctlPZHQ0
9WIeKYKFgg7j5i5vQrqz77Fu3SNQIE72SFNo2xcKZ6/YvKgXtftFFq6fvwfxjGF2
XvbEr6NuayXiOqFw/QFtYdXyF8MG94mSkzEpBEEE6hrTMHhzBtur5MUWAR7tRiZ8
InN1YGECY+9Sh7kEWsg4t0oogkmestqubHcfVloDj/3zXxzIT0vWYFPiY4X6sIGh
Mi6PK5xH9PMXaX4zeyPmSuVG3RyOdj1h0AuEB3hRdxgPMg7qGm3Xop39mzPj+7KW
WoDEAWKuhxLVCPpM2xpWmqgyvA6jZ3QtoQuuoKT6Vv46SxJ/jfPBCxZez4n9Bb+9
UKgrBJEcuy6uhtt5bOheeydG6B2L4DgbELpjZcyuIlOS35bMQ7LNCxycldWbaDUL
AP3i7EIuZHex9YBcUKXByFa9lyfIvdBP2xiw8m5JhlzMK5tACEoz+Qu4kf3GeH/H
FbHoSIOeBEeVDB4npY5VGJkvnD/LlQguFzvEkTZdkQSRGHQhxCl1FZZ+w9NCyMR0
0eFazuYABJfHEoG+Noqe5AfcE6I7EbN3nsMjFCOTjGmQpwU1J+/g6pIdyPJhCGdW
uwYk03u5qvOIVmJoRH9VJnyzLBn1M7gG4vYSnVUcY65mANeCmBC4qy+fL3JTgv6D
X+rragsY3nirQy0AHpFyiAH2DCj4Vu7FntjS48s7AHK1EYf3Q8ZDAtXwjU0Wx7wD
RGsrojFN8r7kjiSE1KEVDr2E4FKPL9Jx7oJKO6BVeIiSLq4cX037HmCaKVZbsoVd
dt1ZffHV2QbFGSLPR60aHhuHP8KTBh2JINaRaeSmcdDpUjQk9RrFqQoYIBwhjAyg
fzl32ptrMFzdR7ODxuI6b7Qgcg7hhVOQBQzx7hoqTwRTAAv1ovs+mUmVHfxXW+I7
Y213LDLd8XjK8XpYMSZ1mKmTec9IJcF9gpWPYRf/TUoex0Gha96qYz4iwYlqhTcl
V5mvuAJwGehD4/7EUZKCKmGf9/Pm0nuU9ZYI1s94f/MohrYOro+u65ysVGcnaQiV
kxJzvX7Ucrx38MUm1VdAwI6d13ylr5i4NDw/+fR3UsPTDFj6GAoD6S1kJ2qm3C5R
EACsfEbOuVWgofxyfW6kHnO0YndKDAJ3uMKXedoXBk/ovOShJ7ibS8pg82TzKJvc
nc58CB+x40ayEKWdtq+fRKBf2qwfYjnd3gMvBTSxv5ztGKCFjNeCKxChY6SVd7No
il4gxYkiuShNg5/87uACX8j5EuSHfgxV+4BhkE5IY1YfLKQ9XPKB6boanf8xOuGY
bVYy1hZeKZdj5FjXbIrHd5zsuB8X1VnvIn/phvwaW1TKfK18yxGUOQBxC/PyNJUd
jF3AmrKCnA8RfwaogfnlUAQBR3Ckmd2NZ/80kuDuQESn9LiX+Roua+O0ja4YJZdS
wEwYMtwGcjwOKgVeB2wpsuuoWcjNIgLtRH5auXB+4rd6yFbpHCzzUHBTmJxWUSO8
GhzxqJt2ysNmJFNuwlxAnh7M/gHWZHI/6StTXVhJYkYCQGEOiH6qRy6WVpTJcsky
DIdtBRHol1MEgubH6jIrSYBre9Hv9uervwJiKUWjGko/DMoIJw82YlDzMzLNmjst
Y1D2t9yztZbiNlP9Zn/Y7G9eIWBwOB867ef2zIPmKpc8XnzWl28clhH7Qqb8FXiU
4trV/zmJiraCRg6FaujXeT04yqw6iR8RuinC7QKDxC+I0IbIF6ddUGb0WpSPsz1n
3rE/UhXGh1zg4TMsvZYAmi5oUexVnv3V5NYnPheKiKhHuAL7U9a42KPTNvuJBtlT
IOHDcFXlxa3u2DFwXHFcUuKAtWKLtRtwoIXokwDpbdTa2HYyYUn7sbAsjVDZSyb0
9ibTeRAW+gU/Uk7PHRjUr8MWLzJjgA5sgGmpEn+51CrOT+ioGBUlr5q8GdYXm5eu
eAyCwqluA4hd8hoOs3u3bVS3eT4lCvIpoyFb4Ybd7upSF1E1SCrvx0TMmJENTAhm
BzOxAq7ex8e0pYqJCZb7uIRkZAwd2kMktYlPiexyrgIssS7VX2EHl8MFB2HdxdWC
vJ0KLzZhFVUhz0JQrriARkvmUn90orW7JZTAPk2eBuYpPn/wIoziF7vKoilzkE0A
A93TAFuwapLiEDypEcIwXIERJSuYhP4pPGPHQhFtDKa176h9B5Jf6GIPlxPwJAM8
eyF3vLo5qizh0H65l+p3g5XtQif8QksWrUePy//FXEDTGZBCSYwfpl7GmXXI5zVk
ijk5DHloVCbzhX+pyslfLt8f/gvqQBD2LJrHoYL2lHYlI78c538eTZWPeyQmaBXa
8mI7c5zFYoGknF7xX8cvXMqF/2cVSC5GlyT6BgNy9SyJ/EnqzOeZvLQVUYaxSY4s
EfPhFxp+18ElmYvziIB+T10ISh7Sa5QoZehabSKz6BSruLV99cqpKePckRiAUKvm
FM9pXUwYVHDALRnDix3sARtT+73epo1YF7PkGGoJA9NB8INCpuhA59834PMvzihg
nW8n5yhmS2kjtIpgyoOZxi/gqCOYWJc3pw1hzfEWVt4XZkq1SMdDWO5FlTMPkPlS
AgesPZPZ+TWj4aJy601IvD3uF9ooZDvOViQqAkTS85Mt38Rbl9GJFSMDsO765XXQ
LzGkEX9ojJHV+ji99XYECGI1EjqEqOgajMoZNmljz3xCyUM+j8FWdpMXgfjBz9yS
cHcYaCBfeq3hwbr4vPFONeYPVxmmHApT0wZySELaY6QwCJUynU2zt8hxoyelBVTO
yllzK0RtboborkzYNqECL51KhRh21WWLXrtd3xLqYjEL+IcQlyyDgkn03jfft3e5
cP2Y/V9jVB87+wggAliuCqvgZ1zuNg0/p4wWUhE9MYSGPs0GhWx4qgx16fM/fmd2
PkpZeK6R/qk8PPuSzcdVB5YiI6BX3fwaYiNycJ3Q+boDC+jNXJ2z83XwSyip9tvJ
U2WV8MxyiBkhA7eFN5zSzspekEIOVN8xgRChZ/OVDcX8fACtuwiiCpw3mFKLf0AE
UmeqixzaLpZ8QmPbm/5TLN1mblW9Yth0AvpBz0exN9/CUh4WQS3PfQwENff9WLJK
Uh8sihEzx1I/D9oJ4p1oEJPPvt9r8XTZTk+C1zExiX/wS76eldkRG9YcQSZ9u4TT
A8rP9HHWvzA5jqeBrZCArp+vrsDzxc3Tx5Fq3Rk3Aj+ONmCLfX6AvxDRDsAtqwBK
Lztp2wnnMrJs8RLEhajrAclOoYXOZ/rLdMEeCv1j1oFGXA10u5DZTQl9/DPZR70T
iu0uSaG91pAJnPuCXHoW+6DTsjiy1P845lBbN06IGvAlk5sGPmXay/yfjmoMCFYB
x0OtrCjNOiRB6lDWOzqTd1MOKxy4L/awZauTRM7x8HNy+hHJPHhYwSVOpNUAq4ti
VqNtl28DNM8v+jZQNiKqLhUkR3vZO/x6ayYLOP8BNWViOCD5sSrBgvI/ArwfOfYu
bHr2FZDlpHnHLHhmcavzrc9vnMp1BkMvH+TAOYHqUeJRzbvd2RbhslcntGx46H+0
qqrY/UUh9wQZ9OBQlHjG+bJ/E0d+2awHcjioPGMTe2ewlaN1Gh3ti8JomjeHzlOS
Ve70JhC7ZlftFBXO0S/+TIBgSOgYmc3wIdw4b3mUTvXIzRXrLfb2i8P4WHlJBUUY
1/c3g/uwzv+6mgiNNoM0EE/v28Mv71/3J+pki8akVSaC5n2gNy8DtE96ZA1gP8X6
DnprEuVLY+kU79rIu/gljh7wNtalwS8RwYPF0nDmDWYIUKw9WSAtUEi7L7jsjT43
Fq0LNO3vP6FKUSjTJCkAxYHfQu+sGJM/ykyOXy+xlqmEFCL4vnCGRvR6Na+ppfkK
lSnH4K2V9efWGZTqNpNpb9yq3mp7R9wHrJlFvW6zpZ8g2Ku3WvN2z2x8JhdFGFnn
6OaYZ5CURK7DHStqJuxuCgYe0zOyrZK6RXNya17xQJpTCcah4jwLgsn4Pm3IKzim
kHgY2rx5eR7bvsrQsL9PKCqWp4htVtNMv4gvJL7EjilCeqs/8MaLdjb6l4Zv0eEy
HPW84SL1tzTuYU5r9Y51ju9Ckk8sirzVJw//hohuM573SCRAcFIksdTI03LXgEe4
ADzzR6GAiD1QPTWfJSlz0LiEG5HIBuF28j+YQId3o0NRqa6PzfY2XnUPA/kqIy2z
qx3Y0lK6ulUAXsJJQ6UBc7lend5lvLbdU71CvwggSELrtWiFcrrnErjtvlBmbUEe
5erZYUilnyfZRUPDv4hjcFCKrGpKHQcEdLDi+carm6258Qhh679DhyUD6y0GlnnI
j/MSnZgFKxjWQw58f0V3OwVYpbKIK+T7lmOP9pIQbiYos0aF+82RwZnZGjjI/lnz
teJc/p9JxkvcsbTmYOXi7d3W+3+NofFgZwezuRGVBqizR59BmULJiW1LgmhgwIDA
sSDNo4zDMgypcfO0Bn84gg1/y7t+PfWmlpLa9eyCvT+PEE9c1eODh9Kg48MO0BRD
4P7nShVjj7ca3O+VLsXssvY0KA62a9bZNixH/qaAWXCLtqzwMgW7850rhmfepyHF
lGu7o3mjHLdE8nlm10trOu+1BBSR42mY9MGKDr0aY4+rfxwVcyJ5zTK5iY/bedui
4i6sIvFG9HIz/krKgD2ZjXmlS1V6mVYzuOA9JVNp8ZPB1sWlVkd7IYdPguP20YdZ
QgMc8vQzAZXslSlIFyVEn2w6RxZlAQVSCo+pH8icwgEVnkvILu86Q7lIX+SzNOjv
zL2wX7LwemV7aDB/aQbMW+do0Yp3ngjtJ+9ZgDUT0+nrYO9Y/hVDLPG78G+Yslvf
/sT3+PP62gLU5JvIIAXv6vS9mjOmBEgaHO72mcTbz7xsJP1NZezGSFeFrY52ui6D
QUD3CnigssFeGkgWx+yVr0l+E0V2chwz9NhxOi55B07DChYmxI3uWDYmffUnsir3
KEwRUHb5JC1jRqwyUsgDUW2D7mUrQCtdqAUq4p/n8vphHGQbV3elxSRYc1Fi//t7
bsD3hhl15Kuukjzsg+ArC/Zt6NqcIb8jNRVeS3TKZ4xO7OivGSNF5d6aL7a2D7EZ
wubsy1klIjqWyj24jZtILJyYNOebezXeFRKJ1iMS1jHC1ryMGOkQ1Cgjov4oWE2S
HiJxI6aZMOFWcSJNBa0jhukwEloVZ2tuU5TTLI8LB9KiTKXIqSiHQDdPwJAcZaQG
vTsIrOx6EtDp3XcfPWNOnO2gOGCGMNYLe5UZwkrUWbBncbEJz+16PANENtLmQOiR
/RZ3rvlTnlpOUTztPXOEEnFSRKnNCZtqE81T8SPR6oFmjizirYgNCAB+1RZwO3Mm
FDh2dU6ZXqa3kS7dCGAxrpq24mZBvWrLZfKd7tlaX7xqFKUn5KAN41TbN0sYQ6Fw
xg/MbVvM06WCNKSefpUOVFQ475yucXV5Y437zDqL8dVTy2i/OPaScqGJGfzlf9GS
82CjfapLXXVfyxhVGfV1Tt0AYgAMPxJLVJTFsSyjdEE1s9hzKaJZjAnAbZy3OdQ6
IPKOIFSc4UsLow5XCV6a/CfyGProaK7zSuQGNxjvbR9hqD7vhQ4xRXOz25x8BfGu
quIq5i1qhiWKpCYL868aFOOOCpqfNlT4hP19vkXMsjNFLAWks7M5MYm+69NZcHt9
THXQqxh0vWnQzyjUxT5r961Kiij0EU93bRlIdkneqPx0go7qEwcrOuj1oTMY1o1N
sI5sqTA0VnlXNaWQKvu4d7wSsS8f5bpbiIUa6hMZuzBXJFNkncMO/2aXfJkqeuAN
AAXM3LbJJzm1QKnId731zlZHEhtjkf87Bc6AaliQYEVpmBmY4l+9wVC4ETxQYalX
JEcCQLIAwG+OCx/yVDkLPR6yhPNd5/ZWOlGIQLHeGFyrZKLwOXgAhpzahs/WZPzU
Q4BbW24OQEZzrWtPiw7l+FyFjaM78AbbEA4ZnHqIgORXBY7TFZUXkbeDp8cUwE8K
ohp2xYTFO655WN+O+vIJzWDkfnxRdHqsdTjIuEzbQ5lKWJ7VeYDEXuXhh/yHFILd
F1fAmkai2CD8pzkwKjFVd0N6p/gqty1nmHDzmavgUlWKmjQb92EMUNayC2QnNqcU
8ZcnKIuV/NrLLdYy+FtPT7BBZPL7W4E87n4D/accWV+KWcVBYP+WIn47VEVwNzRg
SPFFG0vO8kPQ/pFzEA3x6XPHXGnVYpJrGVUVOe6mM2OHh03PPmfJoLQEnnJp5aCI
M/bv7bCTkx8/gv2hIR4L78Bj5rGa1Clbr9Hdzw1R0EkiK8A2vR/HdivfFhqpx166
3pMWmNeZvcLW+yn5PkY4hhF+pWnNkIRC//TUvgDF8MVIpLUk60MZS/DNEeLmxIa1
cnH+jv56Y6slcHniNx5NlV6jIkCsKKirD6GMs+rRiVo5Y0OFSGYpkCodNVoUL5lK
tXe7X/FWzEs980RDd+xtJMd7CPtaL+6RPiSIpL5m+9HNj7p+2EhfIFft+IiWNXkc
WHiU4og3WbRwjqMogUYUAek1F0tW/4eUZF73nJESsYgdav8MJ5CXybWT33z6mF0U
npU8KTBsAo6tMwTgMsB2wKEorn/7BsSh9TitZo3JtVE7Kp8VTytC3sjjyPzMQfF9
bYALpCyd12B2vZ76HnnbSS9XMO37znWF9icizDQtOrT4fJrq9nK2a0FRoWwwnQXk
FJuBZ9s7RHfuv5gUSGQDcIOGkd6Kr+Lch+JQazxh6fnULK1EUOM4Rlh7dLCqbGtM
ludJafjriKejVEl7du4NSrLEGTZogSuyiZpINosyxREqAYbQNbU1pMbjIIewQZIb
K+bNbPwWK/DzDoERVAeyOZ83wWuT3lftxRKXl+47BLMm0R62+bj8p3UoxKe6Ozfi
Q9nLJBtap2jhpGbUnTPIEOqSAWXI03DbiK4ubDGCjwIE6RJCa7P9R1KB2T2hfa74
w6PGuGC/Iy3/jU/JDh71yorKkRK41NI2NNVgg7Lb1EOvv9StQV7gQFcF6z/br98c
HlQx0Qg03CpPoUep14ODp4heyTy0PCOEsgqQ8mE5Bv5yD8UjYwRMr4tz2sMuIRBs
Yd9LlYnXiwurWMhkMZhP3e/Awc1Achl4OEkTiCDrPUWkGL6q3Uoh2AM7ZaSEUWjv
ujKwFFgFe8Z9UJIqoxcwyyxobJL6BRTZUGmtrORid3jEGNjplKK31uukj/kT12n7
nkuoqMSx2Cr0Apuv1WYMs2tTD1ThCg8DNQ6dAfdyESgnroplNaMSm5bliFAOLBIP
SI2lI2HDEoMUvyorP8wGN6N6DZ8Tdo8rqjeSqPltNbOG0Hb5Vl2cQsGdn+WXNOr0
1BT79X1VnQs76FwqYHNYDOoenTs7goKjfD00v1k4/8EuYepT4RwCyFWE+zDhe3u8
r/82NXkbt2s7RsPocTzF7Th504380B5XGObeDf+aDb9lZE1/ec9nvDUOArsUFQo2
53DeTWoKCK6sptokv1ZO2LfYjN5Hd/a2MTdAPlRZ0deaPgtOA4JPK8FWcdYQZC+u
C73WtQqiLaJOU6BdmesKPoHfb8XwSHCP0Dyv/2cZPyuxLNJ7txN0/ST7GYgKIdEL
38EfydMe7xTcQBatNG350Lbiojw2pukzmDXHMDSXQE1/M8YBJsKVR/8N3mfo3r4O
rm3LRwFvP6YJVyHUt0NxJRqEaOhNSdRUjvUJ4f+RmNL2dJEmC1PeJL//D/xifHkc
6wbrqO9lTXc8/d/rgWky/EeMp3S+mgQXiaUc2ka4lDGgavVC3gBeNMPG3IlHjy5/
DZkxeFuWuMklfa+TrSm5IwqhurO5mgRCNFvSHdERpFw+uwI/Is+l2qdUU5larrbG
VO/kIzWNvoe8xXlRDiMj2kvnqYcyowYbAFjcKNt9gMrYgFxB0ptfyVBokQrNRWx8
kP9isN+eAseFbttXHv8KV1OOKU6/gWjUOVXg3EZ7BBhzwFWio4UJ9GkWHtxg+TIk
+qs987mtW1kPpWpfbJ5IX2t4yKniHe3bBI4EepGnx9YfDZfYhqb6vw3FZ4dqSjmF
BhpT3i86t7KwsH3I/rZB7ysXM/6Lk+osZsuCT2jsVyy0v0KwUJehXsbR5v7DzSqE
NINrn50vRafR7sh2b5OSSbN7oeEIJDvp/DOE0UzYMz1kYydcVXeR0JmgbWuFdJG/
MAOYxMHHhpJvtSt8RTtYYEbq8liQxJ0/Hv0IkskITFyMbv87jjzUf8IotMQ/MD8E
j0ifbkgh22vH85+S+vSKukDBJTx7qmzOYSB+Rvs38FrCby2xGfkUF6pgmjVMBfkl
ubkBos+TI6fpFIYChvG/b0+8OxTpOjAqf3y2wUmLimwQp4kfa938AcPKXW6N+KEw
4TN3aZoxeJKnmUTMwhR5ihqO7/7zvQ2wgZhC6RY3+xE9yAWsXwGVt7Dy2ycdkSIF
jdX2gV858uvorF/ixuXbmqKZ+iNcHci6mCmj+MGB9RNQHG2MhOaAiwQUd+boAaqs
pX4Z6n5LXCrcFyMx1yj+vfuPRuO1QcexloRGnjq8bBxFiBugOjiofWTpWmWv+YQl
UVnU/Q+YQtxoU8CfcyypbA8Rxyb0EOxyYsX/7GE806v3PnvnKJFO002Y5BhLGijn
NeCWTTznbEVbATk/NcsHNbwUbRRl8YHVyXpADQj9Y5DUPcolHxq7qjbkiaadegmR
vRDCoSYrx/va+Sgm6pdrKtTiigYwvgP4B6eJjZ0vYR41ErP3+b54btPAG4c8jc9j
YYpT5s4zplEzHH/dvXUH64AcE+vyscVmv7MWbc+8l9h+UdCiLtGzFDgsnkOkBWrz
YwvxpFXk8mI8aqYL9ZBVi+S1xxZqYxjieuOZGEcR+HHGvcg78RWegPQuCKaGn4qz
qTPEMa5XciBjlj/fANiTmPMxANn1S37QlhXwvD0Wut8WrhkoE1dmCXvOTgdaAyMb
mXNaceblw0At7ouHIAAQr1cDqXf0XZRhYU06a8tOIRHhtmG577cb7Siz5FntEDsA
TtKayS9BRnWvqA1KWhCU9lVQakOjIAr1nV3BFGODOvtroRnoovzK+IYfoInKnjZl
2934vmqnkDS3Jy4Wtyw6VPQSZtNh55fMVVPJEDGVbhT5lqv48dm5PV3lVBwi26Qk
wVu4GdRkX2em1zwZ2mZejfcepiHAco3WNw0xp8J5ucwy1Rf8GPIAKtcdCI8PcQVi
RyknYZ6+MewpqxwPIofrLT5cRmQQHdS3tOb41JyUXrCirwEqZt25uRaVgQ7Z3hHn
p5XW/dQwL8QJMaFkuwH5jnCwKxrRZettrdR8q3/D21bkl6tCtHyLAKMbHHO+svrp
dEqJOwmggv+r4UCpxd5QzbBS2e8KbRTdiEzl0m6QKFkqtQBR4D87ENoe8VYI6Dez
SfY5j2MN6r+GpDKcP4cYjIcdKwW9kGiNB2b8v+e54vmtklUfAae9UAG29CChLeYh
9EZqDqp7l0MYoKZHjnuzCRmOAKSA69V9n5e1/J2RG5MEBHyL5r1OCv2iHTtgrD3v
lcIsdEDZ6gH5nj+ZGqESz+Rk/vaaEYnIpBdYHxeIi3Vo+J1eJ29EVqTaWC9kz3Df
u1ij+pTmu+ZxsKX9Avz1lKFWH5Q64oWKyrynNI6y1yFXX+Gg1/9A872MgWAHZlB8
vN93xykYTuynv7xGblS/cKou21zeYbmTrwEDnQie8ackk2X4rZvpBGnIQEP+Kdpa
rLSKtLQe2UE63elKNd1M1R8zknpDach5GHY8z/ELWB9E46gdncYNJ2JNOreoYeMs
OTl95ZvOYvQbQU4Uqk62gsAOhB0n0hiH90qWW9KNS+eu+76eaKR5ggJwrKZsTnhD
vOtl0/s+MA9wy7k38DR85qycgqYK8H4M2dL0U/qk3Wxj6L4q2aASLcym5RFRxypI
XvBOeSlpic178wpfU08jLJjrJQjBiANDK1K/EWlohSgcEyK8Gx6NSPfSPwC5a7wF
jh43BxeIsmaCfNvPXv5sEpsuTAQDC2tu0H9TJ5bKLuwXN9/hlBamKMCaMeiD7PF7
aNzO7z2dnYjuPC3wPolG5DUbWw21h2dpv/+K8//phjiwFckugCIOt3TuLgzJtZ2Y
I5FfAM1ifHJhj3TrEUT6n5ykNNc4lvEWA1tLO840tW2SJSsTnvHYoZ/G/OcyVJ1e
NpznVYZlAnLQ0QQP9OHW7jKOhsK4ZkJ9u6GK66WAhmO65N6UGZ5uGJg7bZN5Mx/R
lpPDNcmRv20lZXQc5Fpk9FbTahqqS3yiT22SJAb2BIvTdD4TbMQUUjPQp1vuNpuI
40OTm7AHCJ2ebytOwhuiPK3RpJg5KeEOGUnAKTmZvS8x6LLB/dF7CNrogNhjWfRm
BulBRjShFsI/rChuoLagNOwFU5jn2U0ECqNrgljk7bfJKWIDn14NmOd61N8FFcgY
Kk0a8zvcUdXEfBW2RUG813GHQVYFKEGpphBwnqgUFkv3L7Ld5Zr0yUt81iD3RY8L
Ke27UYhl3ZlAxfw1mYDURO2InXwk6qRZMLxkLX5HqSOppLYbOSjyqAUf87SZw5ck
/DNaJfXyhfav2CwwfquS9NLNK9+3GA0SPZ3ZS8jYvwmnP9/yfc2606AFq2dg7waz
u9LIPtTsnssJbeLdl2lFf6XXbfnPY/1/tYir7A27xXgV68DIM9gDPMdoH1IIIYFI
cKZ9VDKpp6/hdxAfeydBczLyQQIF+r+YKLhZkZ+tyjVhd6BQIHrvo16R5wgdJtrW
vvKLOY9MGtOxwfBDz9rBAgwUIlXHfXiffBUfenP7dqteO/fShEBoueNQQZa8nznr
8MadAXdI8AWh07XsZaRvYq0y1RCYYPHGEAWc1XhIHUIut1nofXc9SH9bFFK4ABrj
EcTIomMA/r2Sv/IJwRebCjpJycWL6SZ2Yc3hSdc8lToGJW4DDBK3QDRgg5id0Uyi
yKrN7PCFUSwG4EU0hvOcsNr10oKnajDCUdQwSPHOqT0zQEDs8yq1zP7HTJ5Z53zG
9XOnW8AFsHtska82e6pfsp6wHFd2hedGCC+raJbi6+CsKxAFmShFbr/xwLmvccLN
bCaDK/FjM+oB+nre4mkeOIVvzLwwy7KD/GHi+f70xGYyUCTiuIFZ0EyU4sgNivoP
EfmFqBZWLgata0OFgARXxkSr7rsmQdKfwrV7PQrL05kBD6HoNc2cFTnG0FDNz+y9
HFcn60luS69LkwwUwpW4t6rGTsihieOkCr1MFSpv3+5usog5JRsLVUnh57KyqC9n
qAOifzSYhV9UkYvFBSMRq8bKCGhV5dwlC13np8qFnMH6hhBHRIMYLsSeNM383Iz6
xnKTlS5N2PbyQShE/Bz7InZBvkM2K/vJCh4l084pyrlISSqC6/XfRodcFgfX3p11
t6y0Fg9m4azd5X7GFqfdBvT9ela8KDhrnvN/AYjBRm72molNsZGAJI/shKVHrHdU
Na1583306F8rXUCOxi0jqS+AdvP/adI2roamzb2AztqpxWKI1dtVLHJqSgpcRfbB
Fi4yQkgAYJgLDSGBiIl5VpTuyWfORgvvMqs1K/hycj8QMsBHL85VyeJMX7C4lzlr
tODDpQeBWOuPNJDQ0Ug9yLqNwKt0MCd3o43CgxjIbsowQvAby+SuPsCIvjN0Cc63
ET65WCh4LPsOel7ZWSjAH4ubPuaCNryefxjDF2+USIzCOMICYTm/mv0kkS6t7byr
SE7TnuCKBhWqoxCNtSRw9pxdCvrVtnm5KBHJP9vfFoajKrkS5bivbUmseV6b4QLV
YDKWeBJBXAnFBVBHgnHX08Z73bmEO4UP1plDf3oveBJa6zTftHT88SKd2hQJBeBr
Szbg/ZX1stOQzB4pV5Zd93Tb2yN6gZmhQVPDi5SPmg8byreEvoVShGaJKOCyMBAi
pcYsVTwa6mEPZGIMhmBht2cqgpLFxYGgDJmWgLQQWNUA0TUaG3Vol59t6hiMwDOJ
g5oey0lAvFK9hveTf4ASQUBUbrepDygnwJZL+AaNmZDIBE1b0OMZLyFSqPRmKWkw
cEuMo26oUo2HNFjYi/KYsOcwkXxi+OZJKi11tkY54YrUa788HwGLJlLPD2CGuBtN
/mgtWCLE4RxkEjjBob8WH2njuxvjRJDUOf3zQUc0MlwveitCDg73YBEzfQCK3V6T
dE0LWiNsx4LQ0luGGZoYLNV0Bg3QvNwxyuKO5Wu4UjZ9N12CT6Eud9rLYH4T1wR+
9nhdP6oq7K2bbpcAwYaU4ezMeXRex9Q0JzjmOZ0ugd+KK0hetu5qu2L6Rh7JfWAb
SLDOP15CZf0YdKboSkMV+LomSClh1Rw8YtiuXa/h9OKAtj6IOiTi/wGsKPceYE8h
C9b/Elqi/3F6bBgj+GEAXBQzrNufRx5GrAGLwUW9kuL4/weuQ72QpWgrHwy04K2o
5LOQKVFWI9tMZy/RKPoYXByDRu/uYXdUNcmvf6mLAskQ2X7sBu5xFLVNnXuy0dIz
YLTm82/d29iWnOS3pYYgq07Ni+mgDDG6gScKFHqU6PTLyDacrjtG0pc+tyX84pJM
6oKSCM7vHUn6hdzjst9PoP4WyAa/luHs4c6gTxaz1MDrZ07qDPU4kR3g9VzBDRlT
EUmmMBIy5fkyDJonioFONg3uCHqrLnmCQfbg/AIDP8um7Y6PYvb3lpnS3jMBNnuy
2/8cKkIyrVafYukJfTpsy8k642hC0uEW45sLMcBruEUlZ/N54cwghrUW3JA1P4In
u1NVp5H0g0w6Yqw4bxGMiOQhICLoDrQ91ltXY0+Edr7ew4iggM3FSsPqGqPZ/qn+
n7Pdvvv8YGOHLfMtkAvpmesh/6RZbZaBORkzi6EeDJdp73c09kTEjaaR6yVY47DQ
l8dms1XrPm8jzVh81AnqEC2Mj6GgqNFDdWqQWfTTghaijbNIRWAKU0THQ6ve3eba
QsYZALIH5p0Yx9MFbeophrW1h/E2SreeFKQH9PPpz2xxCIzaoF6thcs719nFvdTJ
G9FChldOmMSiDaGDwuuDE87v91A4XWUoIYl2gT99W9A7EOfTln9g6R1ji5m7mWLR
mubvkxTUkWze+4+uezetcORJsznidZUMFN41hzN/PuTrKWm0jOdXGqhxKCz1qxlD
qJEUol/BpYhlmRxv66v54MUuu3CeFUomjegz5J8PPJufZGsAYbCIza/+HmokRsHs
kzR8g4zT9iYAN4k7HP9G1tuEHgYhNtY4jtYYmlFwl5nHUf3632gB0PeW7CQ0+6MR
2GqnAO2wM3JRrvJvRsRiYcOkcJvTPfQ2vRlmiZ4w8TwvqbJjODeUm2xR4WdN6EfT
R/WIS+fakTUQeorUlJsoI+Xi2FU/DdqOczCZxoY6NuK+wcjj7Cs+tp7ky3NMvngb
sCszM3dLmqog/SS+5uJWD6tHZ1mU0kcCWXaSBjcddJnk6YCXCg+lLnV1BeJlKD0M
g61eKhBHOOeefAVoSbMefzxHh71B+QQ9aWDNyPJISGAX41IxrRbR6fTjWbZHdv0F
486yOV99CZ0ruEbJK3ddQH0J5ji4gS5qXOHMqFXr6w2LkCUFnlbT/0yAykM1uzc1
07zK6YCL4gZftF0oIrN1bOcZq8+KDuMD5uMNk4tPxcwOZRMa07vjFrhwcu/QAQJv
OhOYojopVP0HcQne5kU7pwvdvg2e5z+Ve36CDaYirBJC0IYQ4aC1sl6/T6pRSSMQ
cAczSBqxHg9KV77nMhs0lnjrhR0pKs8vd3s6A5ufdP61q1Zp7SNv35uJEnsbJBFs
DuUXYRo/tC31JAaqzKxl+dCHXsMOe523QbdnlUwN2+5eBkmUTQaV9WLqHlSgkwo9
a8YAEIw36rZm210lM48f582PMHfUAR4Av9MvKORiZPWKQFAmDiRd3GQ75WDUxl09
ZyEnnu8doIDNAkfg5ZLm77U8gK8CnnxeyqOXaHOIVYUC3aG+2tjRYFRC2NYHtJ7f
OFsU/6mbJ8iFtKUF+dYWo+gFm7OFdZH2i2jkm+Rb5AMoxUlYjKa96UEetz7h9LYI
aRJ1irx8c8W8K+lVLcJZbx7tXft+jQoNT+mhiB0fF7VAasH9ejdjusoQnXp5rTJM
k248EZrB3u1nz5Pfi6bL84zC4HwEboThSOkFu0Q+jQh/j0sgUWZl7j3kojkCXB/d
vwfx4rAQl7UdHchnJ2J7ubGgermGZawQvlSomxCGAoapvxA44t4S7ZEm6cZZUbjQ
2mN0dtDBJTo+cyfYA238pby5gS3Bjf9GkEz8pKSpFwGTfJcEKU+DC34oHVR6JgE5
qlbYNk1CO/h8x1UaIrPcXoCAH8+Gs7+ugYG3X53y8W+GRthuayGyUA7v/NSOheg2
rToEHhb1G9bmFayyztOYsUis+sWtrJbnOGIX8q/tOPqmA8dqSqSAQPubZvq62TeZ
16BaRpc+IKVCK7Gb5qP5EOP3yPwR/SBsZMUPJevZklQBq2v9bvZivJnUeJj54SqO
2bwKfbvvklFyK9tiZ5D9o0KOAytebckgr7yEIdmG3h7cz20e2W+DsFQfJbP09HEJ
Rz8JeNcmDecGCV1xFzdWkpyyGeDd4TL3+Hlrfk1N1CofRZxskACGP14QeVe36o6g
ZKfJRLEWGJEgMPTm4tJqjGFTnRlbj+jKRP6SbrG02eEgC89tqpn+pu8EJaF3QgSe
/nAMSejHSn6UtR53NDwkjBZklIySXFYNdwcToNHwbhoQHR+ai35rFd/Ks/U1r12+
jkGSrFTiV4o5QJn4VZxgYgQ9WSvC34lXgoPGdnNMCeg5imkXmrlxJoE0v6uEoVAT
0rufWe6Df0wvj2HC60a1nAKobEiZigr2h6usiScUrbiSSRQQfRCL2mGMX7oZWQWW
+KPuzJ17M1R73DagxJClzB1U4IArRweJCZbhDUvqKZefzzxwBvYjI8rooSRB+w3h
XZvG/3xiRob61tK4EhVAFn34M11b4ZBNxbAHZ98jilsCCTATEWFSsVLFI3LP/mgD
NOFvgpsfdaKW4DNYOqaZ24KiHMDtWjAVOebhIUnX9ip7eQYnwprS+vDCQU+001W2
IP+W79fy9Ma2hcn46Vak3ZDC8HfuL8Hb+uQAJDVyxV2Rv86c+FqPQuLqDpeMi/b4
9qdw42j8uTapqDJv2GoiQ9/cRV4fAqrFGEuxl+x11GX7BXckMgfwpLbpn5dLCWnn
GHkB9Re0I4ZU7balupzRax5zOA5JE+FRAvmlHGwhjnMIEt6OPOshLRgXGwUFzw39
5FE7m/7d4+lHNicUvnUf3n63trkW/jUjIokrf7RyRlutSmF5hPhrt7LGKN5AeQj9
w/Hck7pKexoe/RgafGCKEvILRqfSwpSLQ45vDqaLb/eAYqOJNajKKeiP7+l4Q1ke
gcj2OJq5KpMiBv/SV6VRMzYG9MJld86UrP/bJj/2hzqiX92nq+j9uwiE0k9HZWiI
/MCJTh4FiMLs3vD8fJMpkYAdRwUdff7Nta0BLk04PHwHtgZIbXRePmbIAt5Zkgrg
96A8/+JQwAdBviv09HbkZm3SPKfFSdOrUOJieoNt3rrkW1454x6kfT1wZvDM9mL9
KhGXWQCeuHTItBkavVvCuJXaqjScFM6jYeqthiCQ7M/gr7kym3SaAnP3Kk0WYDRF
VRMpEtpB94QeFP/gqBEf3ovteYqwI2/xaE0MyrL4yNYmaecSF4SVNNS2XbUvf9X3
UOmu0p5cSCsR9y7pdRYNFT6iRcGENyCcxTal9t84XH/sn9z6Mugd+c1IzORj9KmL
BkVfaF+8WYlM+qTXo5pLzi2DJAGhJQqphIoTQBDzMNTwfLzUBUErKk1Te6yyPHVr
/ZzI9Edc98VQ4pV+z6nQh+4nfACKEH9jAZSjQj9PBxf8+RTM5SDpKuy3skDMXTNm
WL36NoV42sD04hLMfvxxgK8qBFqb1MRjxjB2bMAlyQ2ptsJDCgqHGlT4WkxTPwVv
2daS0OpBU7cEQQEgWQJ5T/C2EY8nDAeal5hFONgLutwoA5PX/NJp506XuYZ5ZRim
1CUvR9eq2U4oIMl1/c3mH33YyPV3AcMOEJAY+s2ysAwR61trBY0mRynB2DYjqCYg
o1GMDuu15kXSi2fQf/ByBtJyZyVgbSLzAtA6VE8Q4NZWc1c4eStCClT7HkoR2Ync
z86MS1/QoFAmePjb/euMPo4JBVEN3i5HLGsHinp5H0U71+hyWJmwaGjIqZlEOl8O
a3KfWZI8yYKKQP1TjPaIjGhRxXcl5SmsHUZnDjGzkTKskQruyHh2DsMbf5gNxvW5
poIq4II44fqNjo0/Y4wn5+bm0HjbTj57mh22vm5pZClbXYcKRZ6NnndSqMkxo4ln
nmSnQ/xnAXOfc/A0jo1u0kz9tKWHaDGKY8CsG4RduUi7Q7UZmPOqzbFmbPcTihO1
8TMQupY8CoBFu6gFUj9ljUNoS8CTPZuszcKjvc1SKLX7wwNsTlFXh14qTbTyx/b8
oVIeBO4y3swgEFqwrc9reS+CwYtfTrU+vKCJvxHtJTGKKB3AsrxZ+yBVIt+WhCJv
/tVzpX6Bf7MDplG+/RxSc+Kdc82PM05in8LIrPswtY4Qkly/IzvdfTZK1MGL7zvn
Lku0DWE+JO50IWRnVoNE8q21hb7BnlI4Bh0KCCM2vfvGG/Dq4HzwCd0wAYMic/BH
FdFt01G+eFNgS+++W4vISlqCXPdsDsGYI5xCwjngDqidcjt+RGIK5q6xVBEcE9sJ
nz1K0hB/w33inMrFSb9Y7kRAWLqaPnQScavIoxfF1mccL+qbbswXueJ7CjMa9i3/
nCimJrzVSQiwXikor+0wTMte59mBerUqlTvOjgdIUM9sPYNXljtx9sZeNWYgkfK6
PjQT4AWn39A7paUqtfA3N+stpuiiAr+5sWL9SmB4ZJuoAYbThy6mJ9yLV/t0YrVS
KDMIWDgnYOk5zN3vs/x4HvEoN40E0k6hCp4cmirEZXd2qQYM5nlszQeb+SZEQ3eJ
G0CLxLHn+Brx78jTZT5rQrx0cBtPjlEEXa8pgx5Ep3ovF6gDt3knmLQ29xGKK1AG
n0ovjLH6trHNK1c6+XrN+j63h8F7XmKRKgmsTQJgAD5rd7vtvq+MNJ2JddXGpwYZ
hnnPw7vgI3Oblwzku0/kV19ahpSHZqg/s4vKEUjP7+AUv10/md3Rh7HoKTp3SBMk
glplyH/eDQMdw7px41n71d+KqI6s5xJntSIgxhBtQmsuIo3u3bYQs5wMqR8OlQFx
XVGkxSrJcylcOUJwKvfTv9k+xYi1kr94SwRASZwssaPTeMRhxECiXQpGwre75k1m
bNZU/h1Fm8d8zBoMGb1JXCv+tVTZLRDUz/VBS05A4hS5idPgA42j+bRKRYmbEKyT
Cnrb/9P/Vvx4/Icbeof1ct0gYVOh/WMi0B1TtefKxh7WgoxYIFgmmh1OJBRCBnq4
q5XzS6c+6igeyjsW+g4eavTFHi916rEdPzCdIDuQxaecMBTWg9P7NFvdNNpSh4n1
qPD5A0kEIGN/JFty3axF5r9Zsp1VqHx5J27Q4Z4ToQ1JUqr4xoailKDPSLdpzeeh
8J/qvOrJHyQujaOtR/7g4Jvf/GJkzPXcGXqm9wlZiVyXPQePimT87QNN/gBveWvC
FtV5Jbr0nKo0+/sf+1ov4Z9YroXhOyYa1WpmanPfb1NT5j4Y2cHkHjsKlQV0VFTd
cQLFAiGKN+fvGhjzDPolk3tgD49riJOyMcLDgx9+dMLD8VypHOcOdKglHPsoXboO
stHyRtU8Lk9Pa3WmllQpiid9oklEb//L1WRjCsGX2cn/V4XqLWezh3UpJVVlurF2
PK55xr2yxcDEDCK59cO1cc9lsUe8L+lgx2A8ltXegPOawGFXBuGY66iaTqmkotBi
dPDWQ0zSWZRNovtOPqa3ymmiAHclotjkQxvG1NAGImInb2VJUZewWOj+I86Acqff
DdMJkF8oZyu0D+H3g6tN4E+zCaCAQcST++q6lCCp9SfmycSUHvGDcuTXCruH187m
RvEkUl/VLj7lOyMCiF8xt9zOYhiDP9rHw7c6gah5kn8XBXX6GM8vR7LLZD4yWQad
nwujRqOQCcARi0NBPKyqhHh3d8i8aRqVpTGjUQULqv6yhW7PqJZoZchSznrIRCP5
apVwNFkgLOEXih8bi1J5gm0dZ4rjnsshRZA/TX4uBRysyiJQWO0eQcozEaEHU1g0
ZTQ8TrW7cyAprNYQI1IGJ6mpl87wp3WHgKs5g72jX0TkIxwIAMuKZ1ie5vvnsj8l
MQIn1T9sB+uOe2C6ee933yKhAK8VBFMO/yisRD7OjPcGmrPUzd2Yw9NpGSOKdbTg
gtkKkPXdb8kS9Vy20BheORZ7En7pGTyRJYEP4/xSc+X3NoJFePB6W9yXj6i/TNVL
qndYISv/bJV/yYGZQn8bPzzO7H9CtsdA8bBETDIGCtt68ZQyQIF2Mim8bqSwqGtd
WtpCRhI1YX9LAQ3nojNuqXiZ74SXIqjTb8k+6RxiVr6bUOCmnUT4r40GHmEJd1rg
R5UXiSPEuUV19N7Z2Zv9z5LwAG+mj2zEj/ID7K6ACtN0B0XLQ8XOX9mcIRj3J/Cf
ZT49gEYbRlnFgCu7jLI5P09S1uoSeZjFhQ0kxuREFBJ7UcRHeoOpsLEt5pBZaqAY
Afn12HNpScrcAhv2P/670XnlVs6t7pKg0vnnNcHjlvIQqoM3/uOEVArPJ70NRc0x
3KB52qLQNr49mc+WfHTLgmEgl3qKHdVM1Sm5heuYn6Y/klIYcPN4xm2gRtaSuXsV
Jp725qxhUX0AdEoCiKBOtcEH3HuA4XyVs2SpR84mm6KN0EVWRfh8lAweDVPKiZcu
wLimzPlvemHNaqV9gEqQ9qN7/Jc9MUV+VCjdtNv/mdveeyUyMD5FdRBb6KH9MvR8
DbIUfjqB26oGGaDKMzCBVP1pBcOrWY3/JVN/bZq9SyLbC4pUhrpdawHv2xujQPa9
DOyG6RR5lNMU7lizRKYDLtQ0cEVB0vUiOzdV1Tvex3Tn0N66CgZkgQHfASUaUZON
BTESClm0jYiJW8CzejpIbUHkdwd+V/GXMguR/CF3HP0VpaVoCRe3PCeosGrAlDQl
w9voPeNoWHxcW+sV5qsMsLDGlU2m6/9/AufUgWYdFg4wNtI2j55In6uobifZlrPe
GtVswxMBsAvhnlqP/twk42Ib4wVv8RCAPSE4IGuwgrupBZqMVSOLjj2HFiSq73y2
ikF8TKECCd54+Mv1O6sX0sx0yaSLdFOWPSwWlirfJnwjUByAAV5o3X9WU7+aa9UL
gDDcDLJ0I8FLiNxaR95R25rF3run66U/vRVO88yr6tsiSRKHUWCdtdwsUs6Vr3pA
5AzKm8Ds0FB2kFycagkkBb48PRjQPlzw+X+haiiFX2kHQUdA176w7MZXECFohILY
pRI2KDXhgSUp4njecl4CVMmJ0s0loalVViOmyKN16yetLKzKAAy8wbJXSAzET8lc
2p2a6JXClBwrUEf/NpLFt+X7vcFrJm9xbvc0JaNB9yEwQv/br/1wh4Rwee26PaA5
dIDOupZfJpz17DGbh5tuti/JNZffCmeBqyi6NNXWt/KRWy9dnnBDc4g55bJByiKn
ISCsZeJN0yPC2RsJ7ykJAI8ww6lLNBTLR1+G3TVjgNR6n0sYr80aI1ng1CD68fEN
GICTDzRgG60oWZuJGJB3f/fIMt5dyUnbqE+eC1E92bMg9X0tzv3ROidpWA7S8Z5x
JYKaJMq++pwaGBk52RxupZkN0KRV8N1WUHwFupkuJu3TsdGVtCMXe3zj2UauwNSV
OA2pKb8pAjS4tIqZBZZ7emiok43VBpk1AVTvohg6HrvyqzXv2twTMAdo5KkGf+9l
PNXZ9inxCHlabbx4sGZQgYrYmtJcIT3KfOlRndeC+dc1qO/JjHOFw7Zio4ex2LID
CqRVKROxLr6iO13M4XdE8jSpgBPQZw0Wyx2g7QMoznvVw1PFFXHIFgB1WXw1ha0H
pz7pInMzaagRguhvnUY8g3J7DQT76EUMKJopKDrXwCtnwzjtyo8nIlhLdfs3O6/j
8C3ISuub4NFCKo2T1M0fYuTDWYTpMCpr7rPZKSq2ikASWEYpRbGJ3EkFY1Fuecb0
J4D7bVf/IWee4dPzK7NhOD65moJXpopGhycPzPC1H8sK6M+eIpZGkP/X1s4t4PvB
CxShLND1xwY1SP1kgydlpljy2jUYfmC/uNR6VTgyKec+QVAQmHGF5zqoxlebtKFu
h0ojm88DUb8I0RWDQViifFQYjbOdCqOOg8kW1SbvhaQUazbhde7I/J8chLzE0hD0
LGhYv9+y6PZDPvj+xCFrEbE2ohI9u7kBYe/Sw9dgYne/jkp+lHRF1GZRsOR1Rt0A
dZ1x8uXu3LLWWNmL/GlI8qPkzD/nCxOxnh+QmAgcF2b53bske6j6eAtrpl4jXEtO
WQ5WL3K6dTJxOZNEO8hgfevI4zbONXzROkVfmiZ2x1QNbUFOtjHxh1SWZCAi7zf2
Szr/PH1UEu3mUzwFZTva7JhO+oPqao9XwW0rOn6AL5uYDPGC+6HTHKBrZyXAxwwB
bBOcnTvEdN2n9FXUTI8xi2DKcRYKByg8J0hcQhaZ/CmWUK8MwBV7dshV6ezjMh3U
DxTciuZzpNNx8wLjukGVvD0IG4Nsg0FinvJIK7Hu3YbHgqWfzSR28PhowSLITjo4
/aensTUTvC/12FS3foEB6v/KycDSTvNy3aI7KIYK1NccvjnfIgNJHMcZh9Vn28N0
y3Z4d7G3wSgGqJ9knn5FSqcnlGosHAfkgOypppZzoy2ZVuhJqs+bn7gmlrlJ8A+u
Sr570nGFZbFLLCcoASl8YQ4/qH9YXqQO2/46BUwRfGLYON9Us2LwF437+hvFApGG
3vruyn759eLcbp/CPLFjcR8rIemR4U/JQvdeh2g9hEN9nrz3cMl8NB/xQXK7mwKd
hRqlmpJOQC1cFfAVQaJt+sHs6il3srP5PQvXg2xXmUaU9KL+rYvGtL/jQ/vGXKw6
XNKxkwJUPcZZcJ/ZeVJw+/YwlWqRLJQcGFpw+hR0xCNnLJmyIfO0OPAVgFzzAgPu
T2Mc2Fk77E7p54VU21Q/Q6YX+8lbgpUHcOhXgRUUUxxSdjan38+HcytjUQpGpknk
hS59k9p66pw73HM9OhU43fJQt9QACdVvLwmy0JK4FEN21R+jduAAw/HmrVVpEdKA
Nu1KmgFQoOF8WNvsL9exKArQGEaQPM3JJmKAD24NTzTotIue3py82UzPmHAmDYBI
Jq7CGPltV84ZD0iwQt2cd5xXh3OnjQimX3HZ8Zq93iUVEO9M8hEYUHXGeoHhyPG2
22dIHr0qGPUzoK6Sv8vLn/aJ6HNs0YIfOS3UXErSWlinV9+3OyxPxriPvpbIdbAa
QZOAUAL81z7oB5rnfntPgVhQMktRqtTscRsHX1Pkl8cRR+vxA81N9NVlbKvFkW/4
fi9ok3KBSCeLZOCRiaNrUmuhW6g+oxjjsHtLiD+QMEdLPgk1eLnX/ajIQGidxWYx
JpUwNAS3++/0daehYtyEN8yVsSto2aRy4wc+MoguInIQKsIdl1xs31Q2k/FCJ1uk
A2KowLSCQlgx0oIFn2vlzr55cWL0iI8zGDg0cJXhGyLGzLC1X1PLvf8X6TXBCCN+
2xsBM10pkVV/rl91tYXsn+g7vVBanqOuVYwsa8OepfF5oOZkkQZeXv10gTr03WpX
8QfrZnF/HOSmhdxfNGTfxkAQr6dQsZAs1so8jJUgo6b1Ub+MbWG7Bdlht32hyzii
8qEXBVV/dX021umtN+IlNZ1XXQgOvQPJvxzgOvHhvZD0ARhPbhLXokLFx6q3vC/a
ZFBE/+/CO/bg0AjuwZFdkDsE7H+pvaTfcBqwHkmRPyHotjNZ0zpEL87dmMs7bYH8
IkrniwwKF1pe0jMYxLpAP2wCCAE1GIekXcym+ZRy9Ja0hXbtCn5vtfXyw7b908WI
4nsRiezwcv5WLr2SvTQXF9RzNIUU+V++ycWNi764ymgBUCwsChuCA8SQLNjGH/W4
0SFz7YXax1fMt9dU5NfPIbLxoRA0xTvFr+FTeD15FAxha3eXCihqEoT+KzNInIVn
kjwr0YDvri3Ab/rZ8Mzj+vnYOeDtiIUCmtZuqck6y1wFGZTh+cVp8iduWi6BpGnt
24EFfg9WZfLV6HcKhjCY2tcLsHlvYfSN/dVCNtxv0uLagHuYBijPp/brGg2ymc3G
E3kltm4zcJ9HTCZA2p6vndAraTMiaBFo9TLj+6w06OeC6Om9e21FpuGwHzT9tujs
eakf9sjTyTAFxq9IsPo/Ib13c5LfEKD/9hohP/+mUusfKRiFd2HcDljTlE2ri3/i
UCY7xoDA+0BLvsF/ttBzfvuUm9aQN7UJY9bEb06YrWdPaiA2t/f3AkUFcJeCiAYF
/eT9ss7JcIWF9u3awTHTEbESz/6o0g5zXBFruqb3j2w31NkKBpQHky1c6r3d9u/S
pcX200U0WmmYjrIbm8Bcb2bAGF7l++bfG1ljtqFx20irQ2DY/OL7jFAeEOXjjCgS
ahW0/smBedrdFSPxTdFbdYeWfHSmZQfHo5jKSHsoK3pNrPt++6f6hv0HelYe1bsH
oiKk7m1eRQOKh83L9T1VYcfSyL4z82Pn2QbNWCPapRISyPb/6ma9sFeMZBcQVCNM
Q95E6QXjwpFr3l/lTDJRZKNJSUv16e9qRsSEFWLsSb37EV++5AIICE/k5lpsiTec
MJN3ZHHojfw6HIaf6yJ2gHqdoT+JGtzDOHvIW71mOYDYJvIPBdJmHuOmg+Xtln6c
pJriR0Fey0lXOKOeg97s2VMRu2v7BgVfZGInnBQI0Ll0xABZ5hOXl5btX3oBBf1y
A3cs/cpqBx6rYnC6mYluT0QTGmEfe4ix5KGDPP7FEmXNRBPYGT9u3pBAhGSwuwlu
Bqwtz6kN+j4DtkEXDDxTe2OPXYFNCuyoXm36ih7wEwFWAax5jjvM15eKkBlLnnEE
4i4ANomNThcT7WEdlF1u5LaEdXXeh5BjXZGWpgQKO+JTvgZ0QZk/vxPIPlSV+LSi
kVqJBvc4427YgiU8SUAy3P7No8p3QTNU75OAvPVGMXC6d6uvEo+u4ulqa1JDNoN1
/G5o7VEJWLis6KGh2gCBuz7EUOgN33EUadA5jtzvLd//8z1Z8NZTZeJu6YZrW3zu
edXrWBW7BTT6ISPCjLSXHtxD0x6BGcopAV175++8NVR9JECzXA+s8P9RP/Y55kjM
uoPPgHjWgFEmAzJozJrkP2AcQFHJtomrGM5YS7ajGDqaUgFVhhS3VOh1nSgsi1XB
fhAyPimX2T33d0OglVElOFAJOvvCgs5RaMwxggGeBeFAiUYFLgr7nXjPSASCyH+C
dvYWa8gzi8hTDmoHoxGROfpb/R7N/ukAlRPf/2U/CTS3QZ+BNQ26txe9CfiMsXkS
sUNFl9hUMMXnb+DiAFSD0RB8lCfOVXKBJOe9vcpYuSvSI4y/aa7eHfoUBzgSpzyg
1fIH+nK6gzBYK/NyTKkHWrvEh2N1AT8412poOb1si0SutmqwI2dqs4GqA/bF6vje
5XEa2ISl6DgoZjFnCOImQCjCWhKdqHdyFLa/4J45wVEdl18niQiJvd+dGTCHgiCa
4Uuw+TEDrnIKrTeqL25qzQhfO+HMto9XGQdTq1eYoWNRqGqNtoSFxEEekHQttySU
uX3rHmuDkwcZUiU8hs4bG4170GXIPt92XbeAFCGNsld3AGoNg7ovAaX7YLu4N2VP
vAxU2dPMQuaqew0nPkLzqtS7Uz7N9vEEJ5tcQpAHiByXKP6lutXsOLBzOjWq5B5x
nFoif7XcUTgFXdI+wjBHlN0YnJzpNaNwIKp9yCsRsIE3pHa00enZY2pWQRIWUpMg
FONgUUK3jHKSp7sjta5bSorzL2jpaOKFQDwSqftgQLY+7VOifi2m/0Zt3DJOVo7J
yo06bHX8XzjUZ/95Fv1EfXjE6jnfJSTYEpE3ThGP76PPZ2RnILGNo8xzVpaYr5ig
jgBYHmeiiD1A7HDn8qAnfLA7FY0FsZMU3lac1pTgAiQIy9VwsowzIWpaYjXGGcgf
7T6rjW2tudAAqdZhZCOXMgOUrHru1MuyqpLS3W+HQq/4rYKEweTiI7upqNqP36un
3mkApeDGwkkWleqEUC9gOgoNWZ7gcXBkIedzLbKrBCLddeemtafRTaqPAbWZp3zY
uPQWwShr8tKdq9Q9PgMR1km7CqYqr4is7Ie6mKX2SWIReUKn67HXUo8zv8Dt0EHs
RLBMU6Ey8h+w45WNm8vpd/rhUZb2Usqq8yu33vVEyytQmVNKTrfTOvIJgypZf8h1
v7ZnAMqbpEpyzLBN0qoNTfm+tL7Pi3+KFriT1/1PoMb0F0c11zQP2d9uVpXjRN2O
TMjbcwXLad5/9W9eD+vr6IOmG3uuEZ65JSCteSwXl5e/yGyLFeZvGlnWrWyJ9tlb
Ptp5ZZsPd9KdWg/wf+9hpiL1/BA6lPCoC82iPcCZ+njm59EKv8fwbdpbjfMyrsWH
gv0wHSQdY8u4JXYSv6Kp+HwZbFmUoxN7wQHU7LcvgNDqEAj8Ie1XWEMUY3Mh4ZCt
+9z+2Hu7SuwhAJ9y+uPe4Ss1Eut/swfz9u5b9VXiX+g0RVsOtog8oHwpcOCW3RxS
VXd3eYRIyGIUfc5Ny6P0vSNeQfI/UCEGiVjgsHjZKYj4sJd2AO6txitP7OzmNljm
zL7WPzjHs2p7jxVsNUAMVNMieMQB54Puh4BkmZBMDfKyQIHIlwHyuxFNwxnjK5UT
x76WwIr8RE3z99aS1Ezm6m+NgWcCXhGhGUeFrn4Vlf4OE4JH2A5yMogRWlooKUdf
pbAG4GA9w2FO8zzwjKQck3T56wt+m2NmyRGauIZ+YefG0Ck8mHxZAn0tyAjkt5Zo
VMctWLO3AikC/NuO6h+LpU5CIc8FBgryMrs8+WE007ieFBJ5YFdjRq4bD7hWfD7j
94cY0+LgYDcG5rVIndV2w490Ygj60wePwsZS8AWWzJJ254+V2I3HxuUmydHfyzPO
0ayD80vHXbklDTMPBpJdo9dmfv3AZQhS7S+EsYJPSYk3Rq2551QPWIHw9yU3ZKAc
k1QqLtkIHwkKD214Bfa78jMp7ElJGp0EefZFv+tNxgdjtkaTPOeapTSGSCdyeG3Y
Ohc+K4ySppDXX8imvTjaA5/8Qs3Pc84yLBo8U2vupaKzAbo1IDR3mgINdcFnaLSN
oZ4ML1wIEAFp70ePc4Qn9Z4vABJU+wxa2s2queK1WU0RhYL7PRmbrXbHyrGpX2hP
Tn1zaLwLzS4q+K67EquhWP8qPtFQQTIcPnku2JuHteL/tmePrC6ZAj1NJ/1e9tGI
RT2et96lZELjIa2Jn0h9Mu44LBOQ/fGoRRXP+1mKvd/WpC3l8mwREmUsKi22Gala
ZbAjdh3FPS9l4JHsR5Pg9tUfDyPdZmJrnTh3yQtohBKpvHsO5wf6IHcquwJxSxqR
Npltb1qjAxX8nLlWIbp/7z/EOJSVgJ4OWUXHita6uoZkO31r2Gr+QV6LoS2ofHkl
mf6390gJHsvkkIKOnXnu8z4AhGtHeRI3/nbO+Etj+AVkD1HNDIPDzUUYXSuTXmZA
8gcJNKdDA6zhV6zNHh/yX1Y/Ri1l7Kid4dETAdU6UVV9TNXBCMN17EAkG/5Gw05d
1NwSVuo1C/1jrMBStbjwpSl9K1yP0RxhQS7TeAgxc4m0R43eTd6zneFYqe08CgIz
R51uUlC8Nva9JBb6U6nzY4Y/v+OHl6O8tr5Z20tmSDfpMjhhz7RehFrw+F4ricQG
6Kxlb9XNuPaUpUHNZ/u73bMdzbLJqn/wF0GHMV7kPdREEVjXN1nG+5ehCUI2dw+H
ELyFcvCc/uykeqfrE+TPbytRkNdeHPqQij1OcHR2Ht0NB8M5KbOIbF7fMO0yu2ky
X9yBr+3OgHqlf8Ua8uNJnLXrzcOeEOyM7tzyfiin+qalcwt/OFrFX/A0aMiyIRS0
66lh+HKpQ+fUp/5KRw1glmKIMc7iV0R0JXvszCevRODuS39YEdBJaMXPVHYFV6tt
JeeNNx8oL306QO5JUHxUJMX30SCVn3Td/PEWi7L0SPx19XpyuII8K0uRYbS8kW5W
N+mLv72hZAB+k7w51sU1YW7LrrgTzSwCtxbDw+I7y5KJWeE5lbhAEPtzcgf8xnPo
Rlo29JnaJcbi4Gi4NVCiFZCDMrH3SMVRymSofcw729sedvgdycWnqL7fWcxwsI4a
yQHMYkx2P2hK+fgrflHmK7Vv6jwOGM09Nq4bB8oyB5kokRNWYMrcunyxWJF8a57e
k0atkWBZzPtvInkof07+2YxuxGmG4XiwnvXzirzdTpIt/d/w0EBkOQvV3cjTYs1m
h87+nCvomBUPjwGYvtIH9JppQPR8d1WbBehtRnkd91xEU5LDVo/3F01n1BVqej2C
zkmOkOPODJZQSG1luSprbKZIJr/s3rBKQ4D1b3vr0mzDCcfhiS75p8mjRJZTnn+/
G3La2ezN5KxkFjOvm5PxNotdTeTlMNfPfcDrju7U1+mLOjHLq2Rmr73CtTZrMOdJ
o2bssKjZPZ34PjHKX8hW83AOLymotMw5RZd9x4YCsnaVrY+rB9WzLTEpIamLpn/S
kUXgyOeOyN0mR2AN9PBuTnaqMLOJAP25OZbBUPgICzIw8+6uzNIzWAT2YsNs/Mk4
8KxuHThwkrGKTH+K5chuhKLTu2aG9iZIO9EECimL4F1lr+ZrrIgRmYKVfnYmu2F7
jn+W5PrXBiBdWp3T6lL+nYxoIv5XKPLnDQ+KJ/snj03fFG5QTN/POM+G2fKwcMIl
mUsLqJftvd/gpGAVyJIrC/umSVTi3NzFtwyGnTKjf26G+i+cqqiavBVDPlnHCIef
3kKauSat/3Wk4wctOBf+RoNja1SzwLwiBjjIyJzzdx1IKJKZmmIUENn6w1xmoAOQ
gHmjPvLDTmP1OTWiMYxYRKCecF7FYTtwxwCNQfuKSwLxtdtoO9QU6r8d0/bCms4q
CqJam4n7Uhz6Jit5ryVclqXtFFK1uhi70CjoQXTrmPlJcDFYi435phRgCYA+k3nd
0lecdnUoEdyMGKUVGqns2C3LxMuM0gMDCLBntq38Ccw2I3pvYqakHJQFi8aGNGmy
9gZ16cIjXgL1G0e4+A3lUcRJARVlpE/Nna5ndZnoF14FNt3jB+zUhpBSqJPNIzMu
03WiBz4H8etlcNi49a3rNsWi63uibTEcFurm2GI5fuzzJEdiYgr08Tth1wLH14tL
O+wVJNm8w1C6cEsdoj76QR0mjiYXPnFYHmDs/ysSeR08KGpKQ8K2wAsxMQ+XsaQi
Vl+pKG/TBM6NhAXayDkl5jRbcRzPmKMWqMCI7l4Q62r+eWwyrj4J1dIqvPVQEGNC
w3dvBeUTgKrgHvQ27zeU8PWWeBYnh1fh/Y5WSBBelzAcbWdqRlWEE/GDLejEdQbH
5VwNV0WNrjhjHmnwnP/SeLP0AxfKTJrYgX5dIuag0H+KHXwXwMVuWeD18N6eXaK+
r5MK12qc9Lo+1/RZECQWSrHgkWPOJB25cuCRBOy158YdjrltNb6hfYlETMaFMZ2Z
HTghnicbL2Q+ULrKvRICHKZHbzM6T623pGauRZY26wr5cbfSe/v8kKf446wEz8Oh
X6nIvTqysvnuBtNNR2EBztcI0Y0DEblCDTyKO7QpDPYzpzZU/X/nhxSz7ZSjhSua
IEBTlAf0hUKVxFIhRepeak6ajMqtijhmBqOIs1LA4G+lZjK44L5hdW5o+6xrPn/t
5Y5FS9aaRdPxrHRnHMZ3Bb3+S9P0BIGU32ihfOkeX4W5FYh4/CaFPvvdxIG5pHlN
obe0iXdHeATpNVFFwEEBzcCtichrkvSU1Roq5BnSRp/wucV4zKxY6nD5DGm7R4K5
x57PMZowfQtxc8vvMjPa30lI4du0uTqPsvtmIplXQR12nIW4vZasDKYZQrB9oGi6
YD3jIt9O7uGeZ5RrFOSPywIps4TrKPadO8FRlyfGNwrvbhXjkwO+D84CjfvpQQwO
voL03DfFP/FnwJh//qMXby6/khJbUJroFB0iPAmU30REK9alajqJW8YIO645l9Lm
723xcOmjqKvv7FYvHB/LwyszkWhgO+4O0xnEsEFr1PsfV/TVc2lnOrKbvqWNx2b7
g016OQvKBktLDTu9b9wXkgpX2j2GW3+dZVaCu+N1j/NPsNKeoWLNTtZSCWqoEJzQ
8aM4U0aKrgxwzU+PR9vjdeZGlwMYFlOEBYKur9zrXE9ZEvPl4kXHLMa5Eo7Njhgk
4injTlayf3bTmLt8tNKw+CZaH79ei34+smwGy9WUt/P5/bpQEz/p2afFBYOuXx5D
VL/Aa3U7eXi042RtbT+N0LY50HsgYajRtmoq9EVfUNPKL5FpuBnCUJXak3U5oser
FpSvyddCtpGaXAZvdVSOzcL2ukWP3WO12SCbSJ4P4XFEco+G0nLBV74oWYPlulus
UPcEx3L82SHE2p9VwYHmSA6gayZXMzQdWbDbbE2pPx43/uBKMiJOgYXmosdUFZTA
gacITKQpGIJ3708/G7p/kZbsEqq0wQxULdIe9cWhuZVhH8vFJNwSobOO13PJmcmJ
Mw37dX9OkmrMO9soltDNokcF2CAFucYcAY75RPSZPFbH2PGB6UnGcD2tfoZb40pk
UsON0v/bfVvWJpfi+DpdCg5CUMciY9Pknf/1kezS7rNVp2FfTBQyhdF38lyYkKdw
ddOb/TnPN0zwLqp8Iv1sKMEkPd2ICfNCie6gZMn6D5zSXKlJCUTHOGEymxzup4GE
FjL/uxNn6T3e8KXXrk5zjmO+c6ayqVL+l0zKM2C6bb9j5vsiq4zZ77mfsab2SKSg
NZruZ7Pv66gkJe/eHs4ONcZzysL5yTQoXa3hPGoLYY36UxNwSoFFpn564WS+lj50
BxmuJFZHjsa4M907FDIlE3MoTz204/2Q3tPl0J6rPs/aXcwVvZltuIwJkytbCLKb
l9T+e/QM0xwfFPyc6gDK1YD56XvLRh0Dfua2oNyLihICJtbZnEhql+xIBYIPvt2x
E9QeBSP+YyzrwaYU70sZw92z1w+SATVHKNrkxaeRBp+mDbVJ2TuWwLa5oTgc0/fX
863LnDkVBFPiM2t0t5G/ofVnM6IBb4a0V1R1jeai3l9jCetYbe3uq8VEk3wSwDwU
4/2ZtlIPw+FGiVOVdvVFAVI87F7cPaETEhiEYlIn+bpcoABkIzK7UrONNkgUzJMW
XqJ3Z5PEMvvWG7crNrFU9MDju5DI2bWsJMlq07SalQodrSN45yP3h2I5jGAtXDAN
XfXK3jw4NOSvoRLcDL5wHYu2a72hTl098ykL5gwo0XokhFdmBU2qgK4ITS1J6IR5
2c7fa+0nJCBZ3EIbWu3vac9HSplLcLbEYyR/8mLX26EWpE7bpb37Qqfe54Wd3bsD
IQWsg5Lh4t4VN9ZLuNkUD38FuKtTtcEhctIebvDpPeu9/G+8+sR3qhX240mx9ITF
5xWJuwS/n4DKpm3kVx5Jdb1ca8+FgZvOsLiJb7zde+jkeSkl/RT+tpABWxhXkMuN
s10xyj4gZVm+aa2RD9aYVI1DpULKoQFc9YfVIqsb4kW3C7B856QAL7tHUbXprVFd
Kx256cKd2FlX0Gmpk4+4yHGlaWz2+xaq5CKPYNUDZemq0TNcsCzjJlB2PNDT9eW0
JdIHJi8odh/35YfzxZjQAhdJ9Z8Sp1gwwsDBK8d9o4Iafel+ZRZoK1594NFFimq7
lehXLmF1Nf+HA1NlglMROxcldnM0/nNHDcGabYnONsylEClwtdmkDIxGUA3OYzL7
YIzfK0BcSV7s6PNullftyP0gPu3teCLH5EOBt1HEoV2uJCGLd1tyS+nyAHQR0jG2
X4qq8y6aFlXWw5tY1A9/QLI+xy2YSXBGVrmlhlMRAWP2KHYs+DCv1GjsUjew1V7N
RR28u0bFARrTD9irTdSHKe+d0rwnf34aBavzpyk1Dym6mNQGKnnGUCGTVWoJmx0l
9jIGWAoUIRfr2wQG4kqHxm+T3XRpZQn93d61a64zJ6R3gwov+0MZIbI5o76x2KZV
ozseQaoQJUgqqNZ/edFPelAflQtwYuFCyFTe1sxIF7ZUgHQDD2bVW/vfoZidPgoj
wvUTDbMxIupJVMMH+B/Q6mbcr8LFnTvGZQXJqAZzI30QiOAzN9/tUEYBYOzgsAxB
0QIVXYvVOO4/csUqmk5rH0YtUUQyUdgDraZX/LI1XP2fgsla08tMe+HMYZ5gQLHf
Z9SnYXUA/fw4Ssq4q/PXQWMnpmjcqjOydLDXfmWgeqGE68cPY0yj28JEs5m4J5Kn
map1KxkafEbvWF3NcCCmWbUiEwe6sWtQ0wfSg/M5wtIAMzLg8IGt+f1HsQslByHI
qLYv4KvJVfjfE74ISV+3HwWGp9Odt+WDIOLeMwHeLqfhMzaq5gkdc//V6RYeLbu5
KXZI8EtJPxNwCvoFPb0bihjHd/ZljcDFqxGn5OiY0CipMGFO+Nu5gUOR8COPsW8+
FI6pPNODDiyck5bDpuH/I92s/mwQfdqCXd3BNgH1EU/LO/yEtC/Xk9IktsifEiIk
DFyEIExGthGdO0ASMFYzI9as0OEak6azlgie7uXo9JHsQNXITbMX7PwKF/J+sPjS
JJJI8C12JRzXFeE+lRMNeQcfR4OyupA0ZQAQNue8gKG8eVjJs0yOkYLcZzpRZMqp
BciujGg2qqWsbKOGF+vxwD7wE2opnR+dl8DlrifBw+pVFkk9005YXLQ3hUywUsUX
jN59nCZ7iN7HLSH07hBsPq5vgWAknh/dp1HoLgUv3wM32+XFTwweTAuCAJhzh11j
Fs+ZFfvDGuzYdp3SD5qmqA8W/RzTSQSJNPAcye++eFfZBqyTjebRNM7qBdpTHhaF
1VDyJmcP2M9ix0B4BgE5qT1DSOvQ1DUOsePwMuFH1L6TyXHrQFsUcJ9NbUUEPZA+
QUHVstx7DMdUbeHts3OFi3di/Opwkt1wFRGWA85nYCS7k6yufQYs+SclA5YLd48p
dTMVTCZh3d5HTrasGyuHC4i0uOWy6M16IMBWAUmudzvbsSCBRgiNF6tIL5f75yX/
k4EwxRL7Bm+wuJRuGdVo7di+LSweILDplWevzTRKOpVG4uq5YfN7/u7d1GTH3ge8
5AonmUvZEPrKTiTy/8IEx1CpqjEG7q8iPWmcDqQEOKJcwATkAyLaPIG7Tl+01LIX
uCgblhWv4KELiKesWH7d023AR4GDPDC9ga7JtaN8zcodk279TPxbgiVmBrZhWiw5
jdsLkJwiEg/d0kbpjJrwTTADeZSawkDJCbLuWIP2atHOADNbs+vMyGD0H7lyakm6
NRakg5dBZULa4o5t0pghP9Qwo+6ovi++BJPXScw6c8BDNPHnOj6JngqfUe/7Vakp
kjviXpMoVYIejs4RxebrAGkR/jiHgc+ZM6N845VVDvHpGcpAZJtehqaofRdOS1H2
o2WF8ga42qYbTN+YKi6F+kaZ26dS/C4804kxW9FoegLixLrQYzV+mLFFaVL9nshd
2wKdHRME1PuziF0nprgJ0ZKJjnPPKM0qOcTPb1x2fXuuziyvRmQKbK1a44YLkPTh
S89TmzedUG/qlja67iUXLKNbWKgJaPDTKk/1YuZibr188demW5b54jCA9O5VDVmk
hZfoSwpXMNJnHvZMO26erMEyKA+g15y0uFFBgRH9MKmMWuQM3f8ykga/VvBTuIad
Uidmle2EY4QsBDW7Qx/yMeH8uX4h7MpKsVFFqPiF0CQC5zC1t74z/qiYgiV4cwUN
1d4vCiVsRgooccDC6OKLnGT5Povy/9uEIe0K9mzCwBNTn+Zjl2WvxUjWL59PyoG7
aw/GuJ3acLNqTAAWasf1556A0w0XJRgYY/AfNbdOgn2AIiSp4xV7yHC8kA2mftUK
qN/FHTcAyY4ZzhcL48KnSxu/uC0QQ52J8crvQhjHq15uOOcrgnei5hxrKToiZZvI
cYMbV93ONEWJnc9gEP96BUJzrWOpCzCmYmRy28aMsBKuO178I4LIs1qGI1t4bXms
X1pLZBVYhEqDAC9GBBtixOlM8eXI5CVp93w6bTJnCvtl0KsKewZNEfDp69FHgx7e
2wcV4cckfb3+pgMYd8/38ZTIoEMe2MLc36cAlIfMbAdjYGWkniuOCdx6RR8mK7aQ
ufc9P8rNBv+v6GnfDqwsAfQSWUXG4h4uS2CTqn78jki2dQcg7ms1TAtGg44M9+YW
+lQc2NuOH+8xvoloJbk3DgLRS9OyNV4wTyuY5D6E6Eh/Px4EW/9bW9+1hBgn2z4v
/cx3A47oNAViWj+lETo0ybSFpffTP07IsYfdajzeJ6UQzkdYa1stxsk6jj+vU6/C
tOntgtPb34HXn4OVPU656iBrlLKa07b4bG8cU4OJKDzkOR+ZA1WoN76yH1OGpa/f
fiPyTJ0nBzM3G1qBTBIb54CdCqpO4IBd50bzW5aH5M9FzxGeb/Pwfa7x91ui79b2
NoglfBEEADAm6G6mVnsN9D/ghI8sy1tyac6jxAOcSsgfYqWbLiEeZs5M+QO3kGe9
qpL/hQee0I7Snyq1PA2l2gd1lJ3KstFivFBVRBEoYoX1ULJm63utaGPhHASboq72
WcgQ12I6c8TE+VJBPO0zQZBJuHs+SIJPsi8H5Otvho4BDvb9J8BY83jqxwe42L70
kmHmAhYZCJmDeh2vpcm1A0nPc7swpdUXSwV7Csx9+9hSEE+yE+Nh7MD4g0EFHLSQ
KZZEcZEFP3GXNCQTCYUDkvdmqRTmzK35IjY2nnLeb6hNPrvAGPX2zh0J0c20F828
pFbZ4QWzhPnY+7+vxntq583b8eDmOQZ7NFz7OCjaXyyDNs1f+WhQ4EmUQb7CexX8
OPEqbJX6NOZn1rHWWQL7S1DvWQ/KeZMNXIcrEJMoKsVFVcYc6F/fw0o/GsO0ebRH
2SskEDl5zVHBkZbGLfEUY38cE2kIJ6R2LOwTEsOAphV+NWeCL0zRLYMVKSfNDHt6
EcdssgZpTKxbzGU4Mvto4s/q461Hj1iP+8wXhUi3uaV3dJ7Kxl6kbqTOYTjmUI+3
Kmo21ZnhUHvvR7UUkkjq2nzYvxeH1fXSF/33H9HCwhyDzutRkx01yCGBxI3IYiNk
QHNiXdRHySz/VgL24/ZOa5IKilFqg78SbyuKqoLqC8S3JUfs1+k5EXecTTEZ/YdF
zMXHP7XHck0f3FjMHNktUxFO4NENcox7zkL2lTDBYp5Z9oZ/i8Ylpf1y3GIE19Gb
Q8OFx1NBqOlFiehO7SEANTtl5Nt0PtZuV+QLFuy8vXxQVkyWAE6G5E8qLCJULdrA
U0GVSo6q1taakN6qgsy0ZKWbZXcGA2wEV9A0QnXPEOg1fsbnVBQoY2163jh32ZDM
sY0MVNecXQWskPNP5VOCj9UCXQsvorEcvekx0abUcOt0APPb2sVMduNNo/QNQXX3
bldQIruMkykVCNBgUYF+tqBLru1P/hypC3ht+dYu0PUToL0flNHEOWwcE/OcnWFZ
+7pJXCFpOh6qBYIrvX7l9R8Ga4ArgaVmht5Lad4ML9zbdnIjMCl/mYF1BM3ADOlz
VDxp1zYNO9J5hfV9gprGj0450DBwxpMpey00wUZF1948YiLTe1xqyuFtvyvbVpho
RSsCkM/WsQos1dYuK5o8JeBv/VlsL42MNa7+tKmTNqwgb4o5TiKGoZTjl51P/2iv
e7cizwx+Nw/UczpGS55B6+lZwwp5DH+ccBgHUeWL5hoAS3nuxXag1vALqLhaG9cg
a2yMPvLf6ic89DG2S8jfjS3Eec+3CLdkHKLbPXw40hhOdWY6X9NrcOGSdNBWU9fQ
E3VuAHBxLAOV/XojalqyR22PUDNEcfwemGfLM6jP7JFrVg8HNr7tEhdBg6D+awEA
XdFTLfB6Ob5JYdVITe7NV5eG1Nsl83eUYYnO1DMF84vGecGJMBP/DeXS50Nb/coB
EVFrE3E2AgFWT7nZh5IWiRZB+IIlc93mo7tWphARuHbHwK1wCXSdjuUkOJBMzQeZ
KkVQfd3TqysyTwqi1ngnFbJ6LqOzaMclFiV1I7VflMrB6Kfley0a4UwmwNfXx1I0
XkmBhIo6nUPew7QPhCsnFvVbmZUTW2558t278cMYSRnlv1EM5xMDiyfu3/t7tp2o
oFDEbunJV8syuOlQv/2KtSES+W3SZWIPUmw6qq44A1kGzDywKjV0dbpxgsk+5v+J
J1Wid/RiGRxKZyUa88vTXSD2KSDBliec40DQM+tcOkuCzFnkHbzS180VhxhOdTPn
opvMtBDpNmUQNMUrGorA9LmZZD6eCLniaMrt1CcaBOvVDBtPVIyT+QBak7Vuw1xf
GAluEJp+5JyjR8ZoxPZXnUm0Tt/mm/ujnjaDQLutMyUhaYTs7vmDGH5XCNtd0Tj/
pf7uaqCgKqMe+t/U4MzAGyIUJ8MAdlOBS5Z+sqmHsju3Q11piXm6/QzjIOq5ZAqm
eQjR651cvID2jfXmtNS+atduckgpj+48V212H6xyu8ZB0iE5iZcV0R96t426J58O
AD5cfVZKSk8HemXyE35PKPyyOXbnt3XO3XMc4cVksldTrhQXJX7Xf1MQ3G0U/FN8
gLi3FTRhGxebCrM2w+b2M4G4dijzKnsRdW67VhebCkwmmlF676VsY4geMYLzvGEF
0BGjdlyTxCyrA+vBnSh4D5h36Q93pVp2IOMaQu+fFLZ28fEfnx44ovxCOY0C+7EY
D84JOASrYVOuNTpqdaMy2bdUQ0XopfEKy5YPw3CnTsR8kIxqAB06oE81cdYga56a
+cxaJlJsamvOWO+xbTRpHFhbd6Ba8oH7dG27anNsMUPCwRRHR4Oa15gBrNLxmDny
j/+Sow+gjH+lhA34cBqw4s182fCE3yKp+XAQcXqWY92dT3M8ufS9meHkXdCG4Qp7
MVLgX3cCBT5zNE6Pv9zgzpwyQV6uslBIpKP9/dcCg6zQYeXcmkvqWScTw+aggmW/
YBqsVLcoOWSuBa/5kR5H/GkrxkmFIVv3PkexqHTbxbv2rg1hi3oc3FC/sviCOirm
prIpaqngnZNSmO/J3n9rF4mCievVeI7fJmDUohBGoaPdtLQAwTIpge7FDs1V42HZ
zL04LMIASNhdpaFZ7Y94Du0XKYyuOhmrJ1sVYSQVaxfIy/0Pwj9MCl3e+XEWnkMt
wW9pytfx6EX9aQHiWpbb4O7v5hb5SwlMLgcXkRbsfB4JL9G3hCQLW7nF6jl44Aza
8Xv2XivGHLvM9Stpy7jeB2kQst0PlWRa4pTTzqoxMjH3hYBXeHpMXbP0Wurq9LBW
Af4veSS8C+VUPiaUNE+PyfsbfDHaze7AdHDQYnFljNB1nPURMnIiuqpsSCrPrzGX
eOsNqHhz6VuazJ6faF0idt0i6a2eMRb+5Dc0cGKHnK8AZmxi+vfsqzNvFQK5ILGY
pfibscgNN8/oWM/jvZdNErcnzVBXRbVPS87NBGbFthFMVIIgP7mFaC/hg5dMz4Q5
uwdB6VtaSuTB93k+KBF59EjYV+9dcnk65713md004c1pa+2JUGYYC7XkXvbdIWtF
5KU1FTdTyG4G+BrrTOu4ASSob9lTNa+mGcmhp3g0gnTF8D55H/Hj0IQy8n6nmmLo
q/PJfEm6XGMWeIdrs5By13YBBBEJhgky/NnY9ZD8Nb71iI3AEdMMT2/qWjPvsKsp
3eBLqHg78IeADfpTmLpF+8Rx6BHgVjqz1KG67Bl7ZrMbyRMyfGAGeXW0OavqFpM+
AWX8nDtG3A1D2gKwOiHg4k+i9Ta82Vsq6mRSLfLWccglKbwI9mcODsbTwW1CpIHK
6BcUDuSYpurdQIIhOL7LXgvV5s7eal5zQGccoGerpvlY4vWgguhqMlz8qeU4gee0
/TTmYkdtnDtjqlXVF6z9Q+sxPFSSnII6JZK16yY5JWIsTB383zAZz9mpJgoOSfSn
4i9u2LmTFICFNVzBKxLUaEg/s9D16tL/q0ja7uNWnrb3KXE/5lbGBEMjvEvVoayK
Nkprp3y2Jm6AMg1OzaVIpeLQ7f/H07M62TJ7zLD7mlskDUPvxvyI9oDsmadb6ROb
5qVBlQ+9QXPg53ILJZfJH+xPmkRp48YFT9mb1gVPKz0MtNhn+MmvIzUjpXNQs8km
Hm/HK3HPrtyrb6+lsq30K0KMvLcn1uehAKAd/Sk07OGCMdt2TTsqsG1OjSCPkyRZ
Q3x/iWI0fhtv74EKqfLAbbtDtyejYMcahTUPSSb03TmQljxWOs5DNsfeQZ4F9Bx7
ep/8f+mZD+fz1DX+/iAsnjAUZwwkvv/jjD2unGWX3gSVx2rpvk9UadQ2AnGgVesN
l/Wj8G4zaCgztrSbCfYoCk2UK+lgIC/rj1wSRyMlpTAyqNdG73IkmE4UGNL3R653
uU+83oiUJr8gSfe2xvLBNrqeP47hqLwEMCecKQbxMYmLzTFbQyePLOD9DawLj0En
bNkUoVpdxSiQBKRglM75Id50cdSt4MRMjqNnc/O4nwpD+EmVUbnte0t3qHNoqcvM
qocAYGOEybRXAkbOTdlk9IHPlezzsrxBE+k2h6MbsLKD/0Yvae0ilTifzO125sDC
ABuxFHbwTgXNr+iaJ5FdGe3IXXCq3TE4oRoCo2D1P5VLtie3hGY0ZTNFFXrh10bT
bQ1l5Jn3ZCje2Kq71sHTlymg9bVzv+cW6rvUyykSpOll8YRV7zRKeCQUOQ2J963K
nSsEUyJ5Siw+KUCWPtH6AYa7EOLz7L3xMIwZDV0ZlH0mHBd2OAFQo3eOw3sbY2Ai
iFA2bDu5py1ciamJwum0TOAmpcEtkPAstrGNU86HDcbPR6L6PLNigOMSM/003WBU
vbEtPdMtt35TQAMVSDLhDBp6oLSje7LE3DyxYyV9F/7G4dJI6VNMAjZQjixplnjY
BTiHo6nDcWDUehabR6Lflfo/uUqGL9t7gM+hwhv8d0nPAr/Y15PHI/kmjLxwn8as
Z3jfWNK70UJIGOwxM3/i5OhSXuTBld3l9vEjt8qpwCKETIQIyPFkHJXe61+LG0XL
w0/uiflj1pdIWRvc/uyfiEtUCnuryNeyrW0RkzY6opTwGiyaIk0fRbcB35dJsTYI
YO6l4W4/YQZbUy1qdQeBG63oR1tS6jd/Rn8Ie5dju+i2Df2TEimBumq2yNWiJtTb
oXhMJZWxcaotSK/DKPbQXNSYVlP/oO/6XfWZdDeNSIyoMRVJ2NXm8cjp/9htj2Tz
eEC0c4gBaZQP2bQCm0lRic/JJjkevmvDWXWST2/k9JfhxsyNhUQ3ZLSHI8D6O7hv
2xfZvVNxwgTQDtN0O8TF0pqOBYNvo6QnaLFIKuCDRikJwuBbFnXGXWXm0y/SU6/D
J8/+nBBE5CqK9NoyfZUMJ9+Z7Lv+oCUPlZA7pXFfjLKjW4n+6l5RoEHYff8p6cNR
25Kt9P7g4pS2gqUlSdb7v8xAQLwzbTQDcRPHrDEZt4c0xp/ck7ovXqY+gjYfKcnM
mwUoL4Zn8Eokx+x8gjDxEfNUSqTNTZx7Ptv1IsJRYm90uUM2C8+wc4pZzASpTEDO
IWCGRipBcZfc8XeHIGSQAvkWrKtfOSy6Pyw10TtW5i/mPNxazYywSKBmsM4Wo5wS
3GYMvVJlhHucPaWXIlRRB5R9V9/WInXfaihAdBN1DDqA6evGfdkAMIWCk8BcsQiy
HHRpeWLDGanGFMVfCERc6qm8G30uTd9Itege7ObucfM1HEWXLTCLJyYBxZLOZbF4
FyivEx8FZSwHQY76X+1+mXh7hOjSpf2FNkjdgBLDYOdP0gktc8vZX3BTLpEgEfIU
SkG0xQknaYPkiXFetnDhprr64l27sBa2bbqcQzfkDVIyznU8UTVGIjs4cgVWEmmD
LiYNU1UwaQfdEIgbyNUYrxUjaecu8ubxbRFSeTHqjku6JH7BFII0rzbNTwXXX80Y
LULpgDnU4cesVoC2ZNJuiIAnRryczuwpExR0lkwFQP2iv63U/p0AxALfd23EdMo7
+ZZ50QZh4U6TUjFzOhmhHdJByp/LBdCTA8ZZaYw0irrow7hC4cwGSRit+4WOenkz
xT9XCofBHlJraDEyhmhijPE/L3BoBLRamd/0wIP4kYvbGhIrFbMqrH/xVYzYKndh
COXsRTqex2NjeLclE236U2HiiB4ddsiuNwNhoyAI03gfb8YPWKbnYPuSAUYzRz8u
tedQ315mpuUlVoPX17tv+ngSfaxw3tev7JbeijZwNcDqvmI5I1FxKJ7Regu8jcr2
luZ6SPSOEUrR/yRXw3ais9b5ZdMicbpWek0Cg4pZZRChFh2NgqJxDJq6usu2c/bw
6Ib/NM0y0Z/kLkXnYYj2X/CFh04WGDbCdUGKSvOSrO2z2mBXceNugCMwpkUfWlU3
RUXm4DHbqFelmw6ofHngh/scrJZ+4MPRC7aFi58ahIZvY2Gcw7JZh4t7T8kurIFr
ik6YcKDjEgIP22+VmFxtALcG195cMUIru34L/yo1ZgWOB2HTHwz2WcDUpHLPhRvF
EluZWH9Yuc48DXNm3jG23Q7+FrdYX6LEnLgxShJqEOe3i0UbTfB5ZI6vMN/hdg0L
Q3U2O6OSpUX/EIAzjr9T4F3I/iH4A0jx/pAnZqxP0ORabGgiWdd7oXOrp7d5snMY
w9et10Ps1V1GGyKaQpgFgmMZ5IlSrDHsItUVx2eQDiojoBBvIQQwEInTDHOUtyM8
PnfMSEW8uL3q5B9RLPXOWrVcn4KsIjCRNJmZfaCZ41wBm+JYtwg0Yn43I8cuGSNv
u4Wm2STvdYPHn/Lm086Sh/V8BxIr7LaipcIWNrAzSUDoklmIjNH2y3eTSFIJkVlJ
L7QtCEeBeXiubTRPUNzrlvYpWkWat8mhAsp6XuwtSmORxYxTYqviNkq0ZxQGu40l
jpRHJMSks3jKglcvYDU4GIZcC5rXhJx1Vg+nFJR3k746By6WAnovChyRzQrkMhP+
1X+t0xxtCbMdjPWSJ+5l3WIVrvMYum0cqYPZr6gG5q0rDbKTbvol8CGvbU6YmbVr
l7bImDpe/jmXAmMBEJsaOAfj7k3wsEFeVRwu3ILydoiwDu7uiAwUVDpmAOoRN6T7
YSO0xp5vbJoJA6P0DUza1xCr5ho8byk5/Hm7MnbV1UUn0sv6olPj78vdb3BPR1gT
k1NHR/1nSiBRHkZZ7+h/HsznV8viaLzYsJRmBaMdbOhqdDkBcvHhUkHSPuumGt/x
tY/JXTFHNBIQZ9BrY5ll7VVosM54nt1KMgKHHw5zmMzAG3dOIQpgjvKqA3Ce6M0U
diiSkwa34QZMx9TDrxQHojIujLcWRacmgW9WjuZl4P52Fuyr9luadWBlUh2RET3S
fDUSb5fNZrCnsp5kYlRRXAjdP0vN6B3RmfrrfJTor7l+8wj9dElz4eu/gIkTXnDo
J8uHnBWRGSE4kjHrLlZh0fsWLsTf60yTotBXcWeQW9njvMEBs4C/9KBmnhgiM6qv
sIOB6y1jVjMfmpC2nBoImFI9GDofqLkOxUmjbZQ6jjG1SPKca/5PJlv12ilvPLGX
5PeYRfHFpC2JVTKLovA3aKli3Sg5RhlgSIqH8P4sKu2E5ILJP2kg9veOm8CpgGVq
cB9H+IVs0gGDffN+0AFCNJ8v+jf548m0Plx7kz83zckoydRxlY+ZbGykijzyu+ur
viD80q7lVf875tg3xIOeUd/XAX95mVUayDENmp+6CQhwx6Ask1GPnNjmGPvOd2Lr
QlwxNZljhuAjitct1up6OsB2L4qf8BJ0OFxrPOLUz3TFGW7idGamPXBvff4px8uh
VwrU4S6EbR0ESzrUQr08NYxjajEdAUjTfKEDWZTg0eKihTQHsLvh0ajpTmj4YJYF
GqCLKrcArxVQbTrwmJDmRuTxyVnIYkhexPI+v/kLsWCgKHVVKAc15Vr73I6XjFc0
3/HCCMrKB+InN0WYa9vL4+6LIXkFRqQmaPxUC7ItjjYeTkdVC3q3n3qffcC3iiON
xDE+/qY5dZiHs8eCr7te1HtjcQr6ZX8h7yOy83FgFbbpd2glRf6Zpywl/N2yLWa+
JpZzCUvHM+KmUR2W4rjYwWj4O+RUpS8JdWP62+Mz+K0sCnmAobOLdy4iJhlhGV4V
CgprArV84ofSUk7ZW84wRISsBRQvlMIwCKxLVprvpcZjQZe5cOfrYH+J6avslIep
OM4FRRDuz88J9ebb/G7shf5YPDNLsSjnP60jVR6GzmYbSxnW3zTdJ1IAmsTsUNuQ
GHUKPXYml+vYtvv24VPDeE3BGqL6moZ+qk8UtV3efpVP8ehPAUAbDzQJiyfdeUpv
z8Dlvpr+yqfAikQUGsO1YXwPfPHZcNaunKhakD09nuCQPbXweuLhvNNpJPN4cEot
Zhpw+JosVokT4tCUA4G5QmfHzKwakCwJ6FNfK0LqGE6Y1Z4HV+NcvdCALsT905qe
hQ21QjVyZ1JBznmvlGbGO3wXn8GJry2NoVyCL9je+yAMWMtVUF0AsICanclKI5yu
SijnVYBFc06grVdHU3OPMSd8Su3lIcyzKlln6kA3r84q6Mi32Cog9BHdCFtROG2g
mka746EqBaH1RFjgYzd4S7J7FMPmIoSZGaPIFaF3t9eUvfu+zGiSYA45/Xf+sg4n
+2MnePiv5VDyqsi1a+JGYET3/xdq5gcZL9iUpCiV4Rimypjeyw5Z5vAPcdx99lBW
yMD05+BugTUZn0Bo6zkhkDs4Fk0Ki5bqyIYsPWHZD4zcf1EGb2vhQt0yQ+s7AsOZ
YlR6P1zOeaiTe5LRe046OyUHYycAl2rWVf0Y/06nufrG0tiwJByXY+HpscvnBdFl
AGwldUeXO8Ud9lVXRnVuJ4sgNbooo6j3lFvK4e6tNSkRRAUOvegKRyY4C9P1GA9o
zqR52mXEHFiDeFtDfGu29b6cdNxp8q1SWhVZ4hf5hNr5OA+tXw62aZ7/eeUPg4fn
1jU5MsD2zuVdYrfwT1QUivcXbjpJD0tiHZO5s7W6j5xRiapLkE819WlpWHFOMqJh
eEjz3gvvuFfEhDtkKXBVBctZWMZ+cgLMMQjguEc049Z2kCTAh3pXgoZpTS6U+1W4
e9cbkG1QUS1BIbEHfmDcUTRAZbcxqe9fOQETYlcatu5kOMPOvi3bedZAa1pPU/yE
jb1A0NUcKYiQdDf8It3yl7aBr20+KjddO3/wSXLWo/ATCMbp9hVLYl/t5aQBJo+E
4m+y4BSh79beA8Z72JmJ9w/jYnmnSj+sVbbLfmhjRVlKg+0Y9CF0LMYVPPGlsCRO
J1b5Ek3M0P3+gK1PKVg0uDkpkpH1GoeiAmBgU+vLFP5BzJ8o5C8cRTP5FUhh7wDu
39/tEx96auCw8pu9c/jt0Lr5O09Og66DoU8Rb1AfuctfgR50F5g7i7GNlJP6PR9E
PPZtgSVKitwuEjQxvmrzkS33ZND/QWbckUFGuJQXepAuH3IAmeFrr6fZ73TEP2sC
pypoxq25LRepE+t7kgFVOkpOyZTU+NaDVSAbi5hRSRh6hb2IOgFp08MzVKNV6d25
4cfbn4kfAgiTuM81KUbdlypNBYCdwXfJp4giu87R+V6V99JU0vS8Nc++dAXnvcVR
taXAPLqQo0/IOD74fozecWdseJ/S/XZqxkzJ7iE+i1AWi5QR/4Dswdsg72nBKoa6
Lnc++MCjgyGEK0fU+nTr3pY+iVdOTjqNKa94s1sakGx98nSj5K2NHwnntsjPJd3K
XkQ063/s4zN9ZPGzruOF0as+X91UcfDBMpCccFNYiS6sEJ/ddcmqBtYQ6oYjDXH0
ZcvbwgRoWmVIugbRjxyMKN3obwxgm5Xuf2Aa8CJM3lkoU6OSoCy7h6G7hEdT/S3r
KtD2uo90E79FQUXw6SHm0XOg6WgiXZghuVAVv8JPiqB+Tk5zQtN4N17GF7NefiVi
3Sfol1vz4PJ1/Su8iBuI4UWiJKpIFFgzWvmnPgEJKCOI6gWKLkn9zrnIDKjdfF99
wlygsiF3fOz5Z36cR4XncST/gfQXfXkpln9HlWGT+WS45k9BtpXAHjrtkFeEncrU
AY+QNgqtgWnYmycLD5dGHUdQhkjcKc/qt0KDMUmSa+EiwCdoyFtrjcLOycyDshmY
NGyDminx5UAUQNGTGIDUvp87s1yaRmywIWERnXd9b3i1jUC/rNfUnWmcpGjE/GV0
lmtW0LKNRpvJNVSzzLJ/9IiHIuh6YtiTp5kQu9ahUTBFmWSDuQJc4SJowj/UJjZP
hIbS92rgCk3LoOF89vux6T2fBvrMVEtXRUsXj1nDrE4/NOwcjKwIsSJyZMQgqWB1
kl+GZHolXj40VneduE3NglMsClP7Kmwi3NBTZ62V8uPkxTLams9eDDMKxVWjf5oR
AVPU9b+QYmiYhbDn0IxcQkhVVGlpExVA/UkId/+Cb5Jp1PCQCmHDPd2cVWO2vDEp
kQWd7Wru9ZfumhwooDMbpuV08vUbi3Girwq4+JkxN//lTupFCaxidAf5yLbPljmm
HOkhxbeSNrVeyfkjP+euvYzrw6JeIFP6tHEQv5L//RqzcDUkQj/bA4BI7FeKEK6n
qWyW6GmUrePA+aemuJ5I7pfjbx8mAeVtRkkRN5MeOb8TuZ+Mrbg2cok08ghkybvh
gy25r51eZUS6/mRn8EVOYVpPhMtD2hW26sstRd0Sg+fr5urCtiXkOP+TaerShC8H
OAfxXqaDUaHSGpdImqPX6Huz0ZcyqwbxTYTBd6YWjW0c68Txc0KS+XjwJblntEc7
H3i9/2RykXNCsfw53Jp827PsWA8WsRDvbpcyjahxwsXYgqBqstY8YXf+lPsfNhGs
7wYvwW+hfVANBIFg4k8hpcSZkYQxeNWxdTj3EA1wuw2/8/ZHgz3OZf1W8MVqYPiW
NfJs7uP66gmXUxfuNXRTPa7tc/+uYr37hh1vd4sNGjTPaZDpQIhob9YVmFLIiPZF
hPtW8qqDT9JtJzQUSButND25fVBTuC8PasgQIkfHZTi9lAJJsBj04lfkr1Ln/xSH
FT+VNlPREax5tEOfNeI9p2KtIAX9JR9Y5bbEbd+0WsBrVQ7Ppi9jifWIcQdBkewb
vQKwJCIMZHCp379zbtyTf6EZEwUJ7SwS82sNPeUQ+2Ts5f2JshSKlyd/fIRAgi4v
OqXH2z9MdMkU5086BRgd1KD6MwAeaLIYmhIUSvAGWhEaSJV/v5F1wclSoLGR+mgN
tWjIZSQEJTGvRDhT012BZ1Z+3Hd2tfbcl/cle6eyMWlitUL2cdDUr+tkDu1FBaTs
7nySS0OIuoCRGzi2Eta6xCA4u+LPMO0Q3vEpUaObmse7sT0kYZ5aOcJQFPgYvpTk
n2oq6MtIiiFCAZYgjU4GxJqHMWHDXxodS9iadw1elr3hSAxwIJu2jc97+/NGirxP
vnYHjrHCcqZWgnlPzIKQOsFHcQ7uaYcG7l7ZOWnbugt6XdWdFAkA4jwE9fVME2UL
lpHSOhfU7XX5ZCTQ5EK4QCMuesC85wUFWNgecp9bgnM/vLIwmF+CV/BFiTyAmteD
crtshxNTGyVS4bnX+hoZSNUag6X0sGDovdHavR+/eeyxWkYDaJ6x8eAJuO6ydanT
IAiyRTwFV0hOlqoQzYgzO6qnlSjmc+msZTed7zJoT4Dc78LrmDK6t7DPLhGZ3xGB
IGHmM4qftjHqMVjG7wWgI1a3mCwXDWSUtcmtjNRC/DnVRk4ZEk6nBoBicjJoqR4e
YAwymLby1/+QggKb2nlqQMIdvgN7RLFcjXfQj0tCedJgZ8MBZKWHsK4hxvGrQ4uZ
tf7xQq3KUHcir/hYj2ZGDAicXnY9N4w4CEmvVOcjwHBiJP7FU8KuPI11KtviSQOv
yaXDq+kf4M4040HyRDbhPywua7WP9AOygxmVO6dc9BzamZjpOjrOW2jrRKQmZHjX
OYUfFCyPA2ZTLBd3jJl+2FYXiw4TjN+DBV5Yaz/cURBgNxHbZ5Ta2Q+BjdwgzklR
Qjf1hy5IPVP7UH9YqjbUVkrmIn81JDH24Vjv6bi9WNSfkhfEKMOg4fA3jLUJihnf
Vf9ejiUMaOykFC7lS7PRP51cJU59zpiqOtArLXsvwzXNUzWv2HtVHStOWly4xOq8
X7498EYaTICPsltCk3voPdbpa3EMZ2ccetC2/rSDs7sCuwJmvjOh2UrzOufw/qhm
Y7MjcsPcOQjld0FhHesB80nYOZ5BUIqmfgqlYPpGApYfwFicIDmla7a/sW2eDpj+
fN2QuLv1hnkDbY5bb66RPFyFVMXcJRy+W4p7HPJcHEra07fPfRmsGo8uV8D4ATxC
ALakWc/Lv3K/meyeTw3M6TK8saqOUArmMTx5B6wDEysPYFi5WsqUTt+ekNrjb1Ne
BT96JCTT3AI4lTcOFGz+2zqs8LHsr+elrjpyT5wEh76dLW/xQDoww9ks7DIQXCGl
3/2EE/eZDUqbWITTbDfw1bWrMH5+Au+6LRiKmqcwD+PxwqhWkr+HuTYw+5dWmR9S
LBohxCLG0OkGDKsiRUy1zxCOkWT8nHq+Lu80cZqGgwy9K/tZMwQ3J87ZtftRzBhd
JIUbsxF7CcnrIFF+m11J36Mvbp3nTkJphOjUldS5RjV1LZNU0eX/sYZaIRdPsxlJ
7us6I+vELeaORsBM9Ex0/DSIvWPyxnocJ055HC74GUaRYIDz5xYV/3FKW7m4aUaH
iNsW0yQdU97Fl8bt6HYqWLDTGZjNsqiDMoMdVrsguIw0P846kQhIUD4l4MUtTjTa
0MM/Z+rKy/elcix/yS0lQOuXJJL7WyxrUNUY7NE84jm3cUimSNF/iQEJYQWjPMXa
/+30kISaOCZsqGV9k0rcU16vDIo2Va5OVPDLPdcSMun43w+r+pyExYLtTUCtvZ+G
uW1I7Y6Blwc8YQSZ33qDWKUbCCzbcpqga845iPzyCXBGVTjPF3TAsNTripGGOh2h
0sHY1iK9Du2I7ftsO5TeaXcs7m+2UTf2xirJQEvnuEzRj8sTCmo56hvNtH8rADs7
YyY50amPELAy4B6MLmSMOf3nEOaqeNdueGtnt+B+G1cTFkly5Rh7U9us0s1bB576
fnacuAGXzYKeiG+0/qJJnKR415yxaH/P9f7FLp18iZ66gO6LvqZxaiOEaFq/6xjo
qnO7gdVtIXc2sRfWiUBJh5sjBw8hlkzkPVAQNm1KaIz37M0Tw+b/kTFAHmLxTaT4
luBtE5ZkP2MV3cga7gwArb/6xxMusvvlvU+8xEuNcEz+GlBap9c56ScTo11OA5ET
b9ECVEXDAMja3JrByMHEOqbKlniQ+2/sid6P2MAFO7HBKVVF0lKfnrvQfCcOWDu9
bp17Fl83Ljinebhl//vJVTk8pOHBxEBakHJabp+rpPvsvCuKkQ6Kmkn1WkbI9zs1
xzOfsXl3YddbsuFPREA7T06MQLndo1GJmQLNWXKuIQ1d9EyGzoY97I0QdvyZKBSm
8UZXxIX9yvfR4mGLsrPjcc0eMblwcHq9FKIGijNIFqb1noxXm000yOADXP/aqaCW
GiEeSLW7slJbDJjskSCX0wVP88ztJLa6wOPGTOCrmeJm0DB15TlpsnE/xXzvPTN+
0bCrLZPD6tkqN+3hkxXjTmbFsVhBZX4ndSA0oNxown0ThGgBbpO6RDMbCzehMpk3
tAXx8h7ILePfYfFAW12FL3Tm2vmui9TjY9P76eFuwPr6oDjjQU3YYwkhOK1maAMz
94cq8xr+Jm6ASSRQo6uWj9AwwYMb1x7wddaAQkreeVmru9zkK7aSZRU/k3CXNp2t
3vyJppZQJTN8fdKocsVeCJLDYwaNvRNQe45fGCyoWCkZLZYw1C42B/0IIJx6620E
yJHrICtwRx3XS3AeAavbtcw6zQNwJCC0WCaVFLY+519MMF0PXZWxcNKTSqWA/IXo
V7IVgshruGYPRqgLPvkSFIXKQgJB7lBLod8TWZYIn1H7ELdviRDK8R8P/sB3BvlP
+ZFVUDXc7AlZRFw8fD5mTIIFRYzoZ26UQ9qRTlk0HDnegEbDECAplcf4w2z76hbb
F5zhdZeXvODA6FdHwW6oxBFlcKI5MKTLKwCIlTk7jMyUjRKBk5X2kG32Cm6IEWUq
HLb6EtnNVWa6dI2ZD8OOy0XdEWBmJz9A2FzIknYE1M4HWG195gASZFVEWx5lo0nA
xn5NzFLKBPIkVJzh87jlU+NjwXQ280hRiio1eysrWP9zLBEhm8mOLo3du6CVoMF9
pEHgeHkZtmkM15eMVTh86wQkFR4VJQgOEbs1QQ0z6AHAfEB7Vz/5/Zi9/eYrSY5j
EN9NNPlWnV6Xh74/7qI+CXW/fGJraKrJXMlv71XneOG8YD/H8fRkpDCKpHLHKowb
GRZR8M+KKymJOgKa2MdUQgRhhtFOACwllwiaHYUKf9L4jWw3x6dQegY21fJXQqMV
p4eQvT+tS+iXIO5Mmge3+g5Iw76JEJJplN0MJ2E5jW9Qn/CNNrS0maMPLqOZMGDG
uNx6FqirY2Iwmj+Ct5FDR9lQ++FghiuoRFwK2IXq1+3Ti1iCKnYZ8JgY+WIpFhlI
yE13qlWdXVRpNDZCc1J7YmO8FABk14Z9PyZrWOYGti3Vs7UrZaFxdAQiux7+405T
q8w6v1ZciYN7+tx0gFibs9yWgFF11i0ykZphnBKvIHKuM8vFflMrrTk8qXkFLG36
KA7lZS6Ctfd5ilOqu9VSYZOzVq/6MKdsWDkOEnq0BC53FkOttrVMqLC01DZaIAsm
oQ6uChb6zNY259kL+mcy2IV+n9TS5IS10oXZUyXWKHweQ82SyFg5LVOUq9Vybr82
k4obuUknP6RLQMdeZ/rdK4BFHxM8Y7pq0N2HW8T7719YUCPFyvd6pNQEsF8V4TFe
iV9Ib81keITPzj5xoDpFNeIdzsHifw88u41H870pEXOZNlH4zjGkRwKPJpqbJfVV
pHOMTx+GJjCmFf/DhHmrSRdO0DpaUoqE23wUnwLsgH+bpS1C+pALNJjjD64SfNpp
CTFnHZWvlr7ldKhfoA75MCktvZsJtCmT4ugyAuzZYf1xwGbffgRrnx4Wja1euXQQ
LgI5OpXbeToWDNNQ/QofZHlO6xtEFQMfRvQKyHH9mJdQPuGuWX2Z6ZE4xX3ndriO
a8YFdo/56TzVwiZJsbvqkSwDU5oBGqbfxP5pCznVvH9Ms8iFvWgS67nxSeF2lgac
JG6w4UIOo449KG0DJFXNdkDxSDGI70aZ+dKHVExZc3WUnR0DXjb2Rq4WLlHJPNQR
TZzVvyDy9y2ATS427/gJKHMfRjFddSZghSKfslUrO+lI5NqWvicnC5qVW1gnvktX
CQLpImCtRKF4IHJKH0hypdwWxnzN88T8+ahm2/IqLq6hKGXVYF3Mo3soqJg3kC9b
tzHb04pbVsnbdMYXtIYadtHXEkSFah4S1sSVeaq0mAoy51YkeB7yjVy3SuYYfD8m
7nHDz3GXqsmqCUxd1LsY3nWEmsZd6ato6Mc5Qp5pV2zNwpNqtdltwesAs5wPew9Y
ypB89+Nb9CjwFoD/bYvde+c0Bs3CdSMnOUku56J4uqEeUl6vfi5F63J1gA+aGbJN
4FIBCGYassT+OqFKAmoD1vgBh7yChsDz0o1rsa6iGxTQNJRi0Be6nkRcJZAoakrV
2kxk261hojJLXOFRlwnetqT7r1TpGetV4G7dgBLglzI8XVm2I2YrM+vFptO6bugR
AEeHbFNCVGi9jFK3addQbhVAzeI7mwjMAP1tzvIMEtVvQzQP/kLoIcwdhRwJGsvK
DKKKITw2w4KAuHxoonqrZNE2ccrEc0iPMpnoWAQhajuOukTSw+reqa747Wk9riWY
NAfpnhdDRivv3FdhunVeYX8mcJIO2czAqzAhV3ZhjZmkX84zk1voGwIjLBwliD1Z
OzuNguNKeJtFt9CLT/sz23OXIRk/uYw2JBYV7MRLEn7TYYfHRZ4q6325YgD5LP51
3uNCI0ZZC2tKKKlN1kXh3Qs3bDEerpyuuuQDo2atypOO3ckaSxJcBz5cuQ6jxdCW
QmYkPpOdNpnc9lcdUKJzyVtvfiDCaoIYtYT51E41So14Jf7JlhGNr6yE+Jlx2QCc
A8zwgzkhfDmiU9rKp6KVKD/GVPK1JC92Q//5HH+GqZQRqtl1aLx0jv+6kufmnASc
oTAJQ8M09QSsZ4unmzrLIBTZ/Tfn5/NWNX8hZ7S9fltiklqdMpFvojrc8lZvYO4z
my5gsEWJKY/kyknES25VVPsTHBGTbGiKPNv9Mn4JIP9zL3ajRPpGuw3CYmPTXqxg
f58QIne6zrC0IPqK7wFZW8dWzLshHwCDfrtBaL5Y1BOkffB7mQmLHsWqkiS9hvRN
Y7z6F8M87EHnAQbhGfkSzFsa3CIGhmS96iIu44fgn2AXdFUxf1mwDWzkFoaw5f1K
nN0HurRWfQ+m/IOioQySTJY6yL8aAsUQQ3Ur0azJhLAQ5J1kLLPhr8sso5OLT7Yi
XWxACOggChDVB4TVzx6uDGTrcsZUjnLNk5/GNNVrxmQUMLfvNW3f+hdoKbWbyRfb
BgJNiA+mP9eZAnP1iz1fZ7ZlUQkKOv3PWc4UaF0yZpo45HKqKsweWlAakqwyhoCY
fvIW6cD9OhjjnqKV6E/G2qVOJKp7SuURwvcP58IK8m2FlDQVnct+NUokRuP90RWx
zO/y8Gtxfa45yQdc/XtBiI+07URtR22I8coCH0jL6i0TNQW1qzdTcehlANWx3yrH
BhhVhu1R937iKu1z/x6mhhfgzlka87KR3mNrDMQoA0TX4vxubF0EFhNR74S61XzD
tIwuxs73se1dddEN7yuWpo4IhQyOrUyTLPTurL2xzC3ClVUs25bU1CKAAm/CD2wW
VFATTIwx5OLIoQI1MePC3GQdlbWm/keBZzWM9+QlboCIiRESsExzXMuLClkoTWB/
ElhTnBXMZJkvkGllmPphJFpc6zkY0zPxqNLL3otsqu0MoycOi0l5gClX5DlcEo7V
H9CwiBjaVef0CBentNHRU/iRdpuDMzxkRLRO1a7RRYO8aYyuyrEudspNHS/tKLRF
gMuFxRjJaGBtgYfLSx9ptFgpm9LhngSnrmrdJ9rkk+kmAHkH1nqVthijn0hTen/H
mcDitClZmb7osXEoGrtegK6dCSCHCWmQmFkAbIhoCV5WsMdeaf5ofBufRaFuZ2wX
SsAsn9pmepOHv6TcBan9mO5KpbDEbQmT+/3VTGZ9bXTSSSlVMpTTnX6MO0ZdmzpS
1IwD5vhuxF0KRgTD8P6AdJ/dBI3xVJIVNb6+9tdXfB62+sZKrZYSc1Rg0gozI1AI
6+0iq1dtxekZCgM44P5/1bO5WtlY35Zrmbz+g0+TEGzXMtWYOXfDWHhufpS+qVYL
RbK8aYBbPQ0ERRCvOm9TOr/Wh2OUk8xMlhszMO3cMCkatuvt557fXoqVkiM0q4dA
4DGMdJSbNrbJ4Rq6RXqEgNwoIOPJLBfKj2JugxcPcerFuTBDtts7QXgw17jReEmJ
wsj6TA0O1LiwcaldiCvdf+xNSukLFfky490VCklb69P/Hyr3G6HwJJUs15ktRcat
i9YvaGBbBG2sz4knmcnTxofTqC5Icrv465hjBT7dZtZk4VaGDS0l8iNveYN3+Ihe
QsKtEShQE510rA9qKA+MjstZimu/weFwKa1a6Awm4TtG6nJ+yOYP0lJxFr3p7NrD
dWj7KkLyv5DGLoOLqpHh/59PPOQn+3Aw2ZcIfq3HL/MCp7iD2X4UoIaXGGi14U9E
ie4XEBP/8MJEj8pCaHT/J/vII7pFPG1adFpid6MwYWgKd/ZUZMscoK8s4pPh4329
J7nDh5BvGSdF0LJ+QOKXkmC6uPxizqddglG/50Mu4xknBx1IlpcXWCdCJ67j03ll
33sRalI5WD8nsPyOz/NwEcieUM6hZ7pjJiu9P/0xxuzO2oxQ9BFLE6JGV/J9Xshm
/dTNbJVpkH1Jc+kaftOlxXIE6BCQpZfj+yaonneorYcaeiP8XCRMkba7ka695roQ
MLtbteVW9xwnNDqKoOtsiqRyK8V4BgXyputuDgN5tMHqIj/5yfdg1iZ7TV6FoCsd
/XC1jBuGbvPlWzIIXlVjHNSAadkjuc/zoYkFMGrGEBqp82lLmcARj0KQw7RdzzXd
AH3lI1Uy0CErIuPvrdZyoWcceVhyF8RdDkuNOc13n5AB3fybI/6JgJwl13nSc7XM
JZ+J1t8XsbcjRzETnYcxVQCVelJlWP1WBMcwNRbSjc0F4AVTE6kUPJonLv2YeOv4
NHss9M80YWEBQ3NTWsVlvLEjifcxy5bRsT4MRHE/xTBwDHrzeOlgV4O5ctHnuFoT
j5HXiLeXaqcHkLKngfsMOVcp3Z89rP3ma8aJr1qlBx18TUVi6YHt2PqtegNjIkBh
mEx2ICePazd4iRnReZVe9RHLlNZmdUOusnW5s4zE5Z22Owo2UICk4WuadlldMPee
OjG4M678KR5DU5yOA9tNwF6IXYlnZRgiyiDnJplRdb73PHM/5crG9hJ4v6gSEbjb
9KCEc945r6kY2ylZCtz1Bopx1aB129s3ZFKxHgt4zIyqYWaZYUGtA1RO+MVr0Cyg
dxtFn9h+ISQI5mnJW3Mnovs6PiVyRvR4Kdx89xTE9R5eWzQTQLv7RzuPPSURzSd9
IYJGA2jbqupe3rstYKHUKxi6FLkkKzfR4PIO7Kgx5RzkfZ4fcaPE/5u1XeFs9fKa
do/hOxOcqXAxmL3Wii3UmFgdya8dNNEE8I9tSvqgMTONesQF+b2VTmY3PDltA+RT
QkpwHXxWjpniDC2EXtjWFif/ijLsfRLU5XMS38TjaY6jaQiPsG6cARv02PQUB6zo
5XCBm8sqZPo9C9zKGyzmmHNEjsusqcjcyMPFNjFO2GNZ0biazHPLUE/ii4xitn9D
4+Aoy4oHtY2Qwequ8kiOP6MgbR0Az19W+9eSBjtx8TqrqImKnAm03+DproZ3KA+l
3+YDJdtetStXHD2jvUdcs/wOE7UJWOBtoGpl6K4wnPv4IZYz1QX+tAzjTSuQAyge
PsYryDYLuXyNMK1cOs9FhquvMWBR9d80+mFF3XrviuVr7eaKCtdT0wvM4VMt6bpi
8Pj20B/Ed7qWeBVVwroOliEk9Q9NIcvjynNi716j5x9n1j2LrksvGgEsUmSRasSy
zHexphdJF00WnjIuxBlLB50qhZHR4nh6Z6v88t69xKBNSBuJO6oYwYpLHMxDBsCz
+rDKlOm/AVuZjgPO88dY7Q==
`protect END_PROTECTED
