`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CauBsQmo82yvaoo4ONXMA5JqjvUoAUMfCePc32ic/B0ln3AjV/eesk95FADCBNc
M/KFTZUxFivAtFeNbeg3Tph42m9TRDcifuCGElHpDbZ/MopCTNwVNsDQ3mo7kTIc
lkUyCalDc+X7ypnqRwD2kIsfSU7CcZl+ZIBwoB9ImYv4UIbow9uJ7fc68jp5btLF
38r3UMUGW788Kdbz6cyk1oB0C+BG+g3zqJ8q1ZIONDys1G0qTyWJkCZQIdcg12py
j1P9UkGYAtT90kJvw+QVRb2vqF8mpYVkg6FKKAbO5gZ8vt9/PI/2dQGBXqRVdfr2
r8BgK7L1t26227ZaOmy37cJeUozfglH5W3MyQMfGOzaU2fveIeiWdundqvbhRv6v
ovgwGbVB7WnE9bKLGnvjVOyHetDgfLmrN17l/AEJICLDYNUIIW+F065i2adOHWn7
HDliBvLLW5unhAVuNKXcsop0irGD+6eNgtmwXNc2Fv7uYK/f7jwEY1sxslyQgH0u
RHBvJYc8lwOY31NyK6gZvEivUj+xhaKtgVgQEUCc8xDqluT1Z/22QWVhPU1O/V7h
xdqt9E72GSUFsc60BxHlhsqI0OdXB1VBSZi+lh6IL3rWeToyLThNnjFoNnqCMiRD
B38Xxb/L3w6bkWLgjMmPZgSOb0AsXF1acuARyRuTqCd7RCAixZcMaJbxB+/T0IH1
1wYiZAwHgu/0lsATJlo8ryq8sUK7und+YsZlVOEmPn0pJIOTj4NFIXY0pV7h2u5/
`protect END_PROTECTED
