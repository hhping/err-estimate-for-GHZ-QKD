`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ewr+ceEWk9dn8iplC6w/+1xPrHk9o6ddgTxnTfn6ynpGMozz/izfBzd8PJvD3pN1
G34gNLT8H4VPPBRomChTkJ8TZuakwXV0N6GDRFmBxePS6/onak5D3zpQcBurxuaj
tGdQYVSqjZkXtUs5uBEVGsa54zCpwHsPZElAXi1FBl2EDQQCeii0SFkD0ZrRQeYS
re+1xOzJu0OVP3GRaEeuzw0pGdt2loynhaWoWr/VNeKSk3yS1kF0Pd5gx5pmYqTf
Qs/N2Fmnspyzcc+f3TSBTgsx1Ntbpif8H5wJJ8GH1XH3uPlbv3g2THRVb121YSqi
mCtbRAGGVoCVEnE30xIhY+rTi2KFy3wQqYXM1CvLSARABrLr8IS+5hxk3+vzc6+B
/6gVDOyjUkVpNZ7nNHl8wm3WrKspng8VuM7SW+/K5dF6gOWklsT5jBe/rRHg4cCk
wJbz1Lf2PsetOV8E461F4x6yKA7N12kkUo5zN7CpHZW9h6gSFwi4WoiJskAqDQog
eyd+WyqaOEs/NlWVdFsdz2Dvf27P4LC1ApWzutLajtmA+dvmDs8LzMATlbAm36s9
rB4+U4c9S9uEKSroSIgKeJn/4rf7R2gInJprIkDcpGQWxnLinPPjr0HKuScMSaRa
bWzJcLBwC0TMsnYYek7G7hzWzV0UJlihC6rzJex9zb4PAXWHtg6pbD6+TC/G6Fn+
oLDisnCX3UTABbrNqCSaAaiftffJ4KWgzIMilc99KXfuMKf6YJ5/LB31BYiD5gXg
RRgcRQCe+KrG53Lc/xRJ5hlhAD7kS8Cp4to2ydAY/30YNUZLmK9gtYpilZ4fXcls
`protect END_PROTECTED
