`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNvu0ClDfQmgrKdhOdAwZF0iEHH0T/Df6Rm6vPgKoM9FAVjX6mmfPJ/WXc1s/dT1
ilPDrbeyruJ9n2LtdiqQF00RQ8biaewworU94XYbtTRMw8eTUIx88Xf+PqBAA2U6
LdQ/9yF8j82/wMHY5ALFs0yoC8nyyqphwAeWtTw3xGClZuXp95/HcmGJQbeGob/+
6j2Yw1T316qIfhY2lqnXyE71qtHS7J393z9xtD1jFR53cihCDWn/1QJUAaPYRD9q
uPyMBpk1brxOREPtFCXmvLJQs1fIpYxYQVPSNELtp2FwGf81TLpvqiFLbE4vUFTH
5ls4FojyV4nN2RjDfjxhYf4T9ltrrOpGmSx/dwXnll+EzZkYYQqEFwO4x3RrnBgh
iabcd3hmeZp8LexUUoB8+7XzaufOgEgelJmJoeJ10F0oHFEhNwc83KCkk3RuUT4T
FgFgZoC20nVhZIRhm/Fss0yk+HKEyRlVH1zy8Rgp50O/FaWNkKKze7mmRjd23Voi
cHgzllIr6989ZyBte7sAmBS8M4jxmAaEdktGmvlS7dmgiyWuD6AhicMiTQLjDo6m
UTQYrrfjHTaCvVMIOBlqQcpv4c70PPusM7+ajxVo979d1YrWZBDnfsU2zi6/H8s/
8QnWgHbkLcdVUdVT7FfKvB8NtPVxz2RcVns3Ln58ktdDaYuUHPuAHahcmmTyGuVl
G63N8OFrJzUU9zJ+wwHOqK5laHQm9X+iD5Y7GydAn6BFC0/tdBKWn5FFFzOF/cJY
4RNJHz6xdz3otFPg9onER0BXH6pCouhcn2kLhdVoPFIfXbAJ01D2426JhZ/n7PO1
tU9jUGjoLKD0rkBIfr+GASMvlsAANf/sIpVgFsyBOvKNTSYgrmkZhnBGXwu1bCCi
lYBU1IAxkDpX5IWJUyACXVrFcU04Kh4sokWOUtV1l7QQTO5jJnd+1fQyK6PtvdTz
BcCYSy3JoUgYkU+YOrWOoK5Qh31m0z4+USRVPruGhICncQL0aVnod4OT5C/ZCqk/
pshctVP2issUGU0x/WTxYqrCi9PwZE56CT/668zAQ7cfyNRr0mXu7odyK7lQ+t5z
PLtoOHOJO95qS0evtf8zWTz3DcPcM0eARIjh9HFiquZOyrLFMI6x+sB3OzRuLswC
FDG6jbq0iOx8SAG8ikTQPYdL3zvUj/Pl2rU4nZRTndUktpyDCj+KIbJejXs2cV0c
jgq8GeIl1MKnGms73CVRKWKcExDC5bsSrqzkRP/LqNnGylGOiIblkNjzYEc9BmWG
R5xYgKX8YIh6vtMtSIZ0yA/gzgZ3eXuFmDmRiMSA+x8twPzcBgY2shQCoF6DAVe/
+jv7w0h4Sa4M/FXyhGO/slAjqd5F0719VowSZxIi9qHW/HUVjptSSc6w70m7viVZ
+/NFn87LJMaXTpnhoheKCq9v+a9qdb2TYZCgjIJivpMeva+nOQC31ZPQYCCUvRcB
RGVIo9SjnYS24mjCbRjDwqMmTE+NkMfoUk127pq1quy7m5Jkjin7TLKZyfxCAQ/R
iNOb3hq6dIKLgHomVRWmldXQuTqURdQlgVZcB1jMqTM/Z9rfsM6qr9A5V6wyrVtn
rjHMJ/HeCfZHFnyv1Q4sa353FDnll2dzWGlMkKduAKVlXFiFhvpbObOPXiG7azUO
9nYXTl94E8y4KEV7z/87tRwatlrm2UniYZRgwYzvxeEef8dFiT30v/t7EMlwc0cC
B5FrNf19/5N0qmojlZ3xC9Vqlx2TL4+VNvcbwrjx5qNXEZ9cgE4uMI0Pprtx/0RG
i8V1/aJJF0D3qS4YnW3BN67P8M2TY8hkL0xFCNSTmht0qAEjtoaHOkvDJSMtHYq7
859aSYCQipEZG7l36e0WwNfxBYpKpiev3eyl0tzWtGUttVUoOheQP6MfsVI8RqX5
rDpHGP5ZIMIXDvj0FdGWuN0a4a8dwwA1WA+fAnscynHrbc0kVXP7oKoi4GBrp0u9
ldbx9BSEWsyftNkK/COxGDuxhlApo1DCIKlz+qa+5q9sWx6qZBaxy5TXP5Nfa9za
hc6GgYm2xHFrPqWlS0jg4L6oWch1Gl+VrGDJnsxIe0cTE48Ue/D3a4TxA/qA9tQR
yvkGvdHWZYAlPdmb0VDgbMVLtozqHXF0FO9TgMm+4jP2Js/XbyeW//Ch7U55UBtX
TdMX9r2KPObmxD4AveVVQLq4AWCTv8WQtxNToW4Ce64=
`protect END_PROTECTED
