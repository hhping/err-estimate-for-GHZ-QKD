`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3xenOKIU35pmwPjTKEYvu2iRxGB3oxPjwJHFKOfMsIMt9qVb8wlcthyLKnb2UjY
UNHL3YOf6qWm7nE9dlXxMH1Ezf03HJKMVdx+MRH+LPw2AuyS4NJliXzwkU/pyNhp
O1xsm/HQWpS1fTb9ypFEKRK72DgAJfX3ntWiqiq2JhacteX5Dy8mr33ytVYx6Bdc
lUpShMAJDJzFWoYA+hGeOnaj7cg9E8+8YmNCMK/eF/8wUI2vPqO6ctYE+RLZvk+s
MwTsiJHYWKMlJJURleU9wqPML5vu8zqz7aLGk5koVMcZLEOEdtAyE0ev2cjAe2Yy
awt5PVdivQWCi9H8Uk1097GkbASNGf3me5vpOU1hXYJ1joykwV8VX8Kwypi81Jpp
Ma9TE8o71PbuW7iD2hNhJLZr8BPHMVNcDa8Yv3aeS2PWoXplmlodqUTVBkqLQ5Qr
5pFahpyTHcBSZaOSbBw9bOLSL/N7vQJLd9fG9BoWkZf9gCaTEqiTg2/GFDFw/G7A
MhVwKLRzNVXBJ/Nv7g6BqM2bxwngsb65r38OPxtrm8bsE2NON/ADb3Lm99gLjESS
z4QFWCffV/4077/BazMkS/2zWpZi35IDd/LwJRVlLYiv8G10P9/+0mE835rEyF9t
msLS1lC6KLomFc0fYS2tl44xQW0qAdGPfhkrXzPS7sGA9cDN+AvrFdV9Lg2QnKBC
KAccLlPiVuj7wYZxCKSDj9b7AxwfBlQeS0RiAkF+inR0ypw/pYCIYeUfxsKaAAvp
Sh0iSKgq/q6pvYabEObEWMYhQKaYrCrRO9c6Z4Wvo0dUXzuigwcwABcF+zfkegJr
bs+KePqYoNL+fpSvj9ZfS8b74S+iQxFA0Y5M4Yzpx9plb8lcpQBoyqEpk8B9IfxZ
8QgrHfZ1rcmYq3d16CezKolauKY3DjZGRj3yIO6AgOcrDpz4DLGYqNOOEsDpgOc0
H9aHbSJxzq6+wCsB/eglRkYjFLj8Z8oUsC/Xzh0vNTbN+nNpG4x26mW2cVpK5+oZ
tw7kg4QS4XVssSlyGzbt/fBIGMdigA1Ar33Ja5v9Ec/df1bfnvf+FI0pEW7AF+GV
YcnTrl+C1dWQoQAbf7Wj48v65bBO4DdOz2/rVJfg4P34Sd2YiIukS9dKlA6Uhzt1
iGj+jxtfrVxUbfgZMT6C/LzZv2IRAfqdjWBZnKvTWe+Rzem5ImcsRzwuvu1zIsJY
yCsd5qcDzSoJzeiLayy5IUTCfK2B8wSCpDqkRUNggHWu3sOCz2cIM/so13iqkvXW
ekn2GLaO25km7VvcbOYSvJiCliwds+d/Zl5mpNjwLbPHzjKeO9Zp2TrTbXQjLOIq
i8UmWjwRJlzNFl488SmqEUfPExsLWjRffPk+yCtm/EJVqTDpotkhPfNDq3UhfNcL
Jzq22sHrY8s99aAOn9hEIW1lWC4fmAZEuTV08SO+GKjs4A6aSxsZz2gcCV0iFdcp
afd3DuBwtSDtLNU6xJ3ro0CeY8uAXuB4oo3FZmdg+QKqvSV8/ApRqDistr3uu7zs
RcuNyAzzqKG1xl8nkuZ4xOjYWWQt6rog0BQ/3CaWvh4nHpp+kD/0uhBU4Zwk1tS1
ou/Yo/k1S1WVewJCBhhZZI2izGuqMv/TyReqGxVU9TSEd5yEbmOi1knZU0wMrAH4
QB1aSD6f6tEnUiT542bDLt826/CWJlvSdSCfT0I4PzJzTVOcLv3j6BnogrY0WMli
9HtKheCkktQI4GKm8qyEX5u03M2i7Imqm5s/uLAr4VAyFtvftv4icWLr7bX/YrLJ
ISAExBzePbax5GFI08HDtg==
`protect END_PROTECTED
