`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PISlbRWu+TwhilHQEZ8XbWynHZRfOYlMLZC6BVO8Rpo7TANhD9wMG/cKuSOGJcUV
2piJ48JvbuGl3ETHouWQvto5V7MBIIFQ76ipbHGp6+dW2CP/uhMVKDASpNDpRrmM
768JgACRa2Nzg8lt6d7YwYNlRQVSi8ihhwlo/IkERnAs7FMuY50dkeztZSB1HeIe
v6mT4UcIaeY6GBw4Pp8xQCZyUNaWX+ENT1l7T23vqxflV1hP9RkfwK/Toa96L/sM
t7lpGjTKheRrwum6JKgPDFm+1dLTqRt6zldZTjnEQ6lfHO/FZL0hlV27l+Sso+L4
5Qly/IklUoOIHMD/DJJj+F6xd92eyoX1/g1pfUg4Nlo6PFaf0HOcxypVZtizPdHA
WGpodtLfHsQJjGl93p6zUqbu+4wANImgKIvBn5ZTQ6KXViQ+lQ+tbGeslsXO4bG9
oC9hVLF/E7/7h6/fEoA3FvI2YPUK2sivWv+CABi5PzURAnvrbzELSg64JxBkMMpz
nhPN5mLjruNFS60cjKx5b4oMtiEOtUC8/kns+t+r2WO+llOq9yPaj201dtjafqiw
9LnUu6u2ABofFctZQETZHxBt39bDeVlwsyVORUaXZTpEUOq8OotWkndck75jZGCQ
lZGVnKYfPKhOa9TvVB4G6Xc34pBJqrKz9ukJPAtD6i3sCOjBFKghqqTKduwfo0ET
6K/L2v5W4e7GUX+7qiNWeE8XuM0ChcNefiEqfKcstA+mKHzlL8gsUYRdBwPOxj+7
7ICYJQghs5N0XTiCts/s/pSpsyqHG5yrOKcdrEWT6rPAyyxBqm+pTDt6ORlek9Md
i0nqMV0Jo/kWpJUsqY0ctkTCQg/mf8bfwq7j/lV2f+CDUyBohju5wS5pM76H4TK8
ac2eE3SLpnQ3zFqqrPysteNaLJDZazf3sEusQ+fWZGpeovsHWT8AhOBPpiFSegga
w8bTu7SU22i6XNmj4JB1upaj4X7qmBHjlR97jQgIuQscjITVEe/JnEVmMJTZ7etk
U4FtIjUyhJ2Y1frWXEhmKkkdJUMPaAzPrMI0qnVKtd5eDdEv2BKTPzvfyao7p/cl
zJETjZAav47m7OXCWw9RnRpzJkUlCVJWnkhetlzpmGDnVyL6KRQ5B6YN/2Dk+z4j
V3mYERyUcZWoUdBkwRg1HGrH40EqzE9bYfBCGrQ4VqqbufvtZUPxpeLpV9bx0QHR
zSFHajNWmW2F0t8476f1ErMVHHAtNRpjzNuaK6L9PJZTMY+CTe4IZPnnscBivTis
dzfrKXCvdC6EtYRrZ0cdITYPK29psU/wVv2A6G0Gu42yzWeD+lIsen95B7v+/18w
ybdkd28trBNuUtrVOjjTDTcVxHMK1/WqsctpB6k9ExPTvd5cGa+lH08f6WfWPGAh
paY7JuLHmuKROawrq0YVs/sQuYovHGZaGg7rawsT93B03ZiZ9cj3ynM2shQdBgJ/
YXj1Ggn8lWeJaRUEiathUuEc5Zf8L9GfptNSd0P1oWvs/n/+gOurDhKt2WhncRSj
5liitN2ls5iHJH/HcmQt01j9hIsfpqInow44GM9+FvE2VnIn0duCi0yYwAcN+Z9d
05vTDSEwihzr9FBh766gcrryqaoxc+21L1lfoDbqDy8+LXFPNJSx9cdjzTdAOFlC
N4k/cme3Cj+zdynrgVut0UucafCLEOkwIbN9+yGviTVlFEiN5CYMivmt+SnKDmQ/
JiPj8f3050Ii5elafTPSBzQJA6YgcxtCnHLfeS0NMkcLqQETo1XUmTe9+xiSjkiv
P//Ze56BDs3gK1Eppjg5pEf5g+Stg2qrxEkCfpDAu/xQqQxUy4At45LGRg57v99Q
bK1XGQrybOKEHwI9/nW1CLGoHbAUtYmpaD933SByytqMlE7kJJCj32Z4hB7iDRzR
9l+ny4UN6lFx5kF9DE/sBh9OvbkFtue268q1kdRr/b5NYcnczP2Id+b9tXfz2Sis
yhDkcpNHyDWd/FvJqmNzjrY459cPfWMo/efanMwVdXd1T1xTzWKJSN40iiWptegA
2F23S59P0fJ900Jv/0YwlPveW6hdnDRf+om2++93jcTOykYcxYA9AfEc2Chq88LK
tRWSKXvVPzZZAq1+wmupy3xw7rlQow0aDFOvWNn7PSF+BxETCD7Dv5HHV/kY1uIZ
o5Sf9xkbeP1csu85sSwF51A4g4tUQjoBQsxJuc6UlLsU9B4esmvkB0ELalQ8mo3Z
+ztFlk86y/j+EAPDlZiqn6DsVEycYEmuud9wTza35F6y0yR+cnICmuymjqW16S9p
I25Kyav9bSR/IYLVkc6SewCGrwKPVpWL2zdadRX0eS9RKiIaEZbTkwg9DOCzfvN6
QoG2lzrcBzg7obURkvNmbgs0yBaNkCeS527mfa0phTG/SHlg/6wjJh7aIoiWi39N
s7v3YHBvMYZgWii2PJY6UoewVY/oz29RLVtCGmfIj+CyfTpco0O++ws2sDllfiiw
sgWW0wFTWDu/iD2sIq5nHqabZwfqGU0ERN5bf8U36ewIkuv3pP+NZxoipbxjT2fe
ITNU3U1NQU559GeBiUyCeMB5VCg91G+ih3oPoC3J4nWZ8V0XRGlg1A0iqJWAE6hd
XeH2KxLS8t5fYDQTt/oeByfEbJae1XgPmSZAIgRVkj7gaoIAKq232KN71pL7azTW
dK6A3OmsN4VeJLnoSFU4+yGSSC8s+BXSw/nwxLvGmTOqXIp5d/kKCA03g67McdVe
Wi50LLZHYvPEhyc+z/VbHlFiz+PKTbmGqKYwCEUP4kEfI5OEDZdvUMTiX6USVitq
ctK1Chk5oqZhaAYiW5uer9kCGWTk6tuvOHeTNKhUtLdZnq6v08/wErPVwnAd8318
zsEudFcKQY3qk2qZ5uwE3eLKZlSNUA9hh90S58gdA4sm65tCdqxV5elK1FAyqY/S
O94NQFh0OG1MeTNkDqEkxK8dl6byCMKi/yXoCAbI/VsDZTLDWf1TbOpUOAMnJX6X
xu26pCtgQ3SuIKXKqUd6ZzzKQOIi8pZ1lNn4aXOwXTXi7kPziJ4iBKJOmNoUUqkN
pnFQnq99ZraLfo2z8sZHb7bdNwokmSwOSlEdvQhK0Qt7UyaOzrBieG3mnL24WyUO
BgXaYOV49XGmAw+d5cGeWCLtqmosYDC1ThMOn04RpiJKQ+GTTESB304in5/sp44Y
i1TmhVSUbJzi+878141CCnJH9U6ON8erzgZGYgCjMgXzdjKYrztxg8w1Df4vQ5VI
YL3NqzwIsmaX98uZIhzJc0VorTXWzz3MhbFvFruCumOqgha/HaT4AZOC6+JTP4Ro
86Iqec2SRjClqqio9Nh92CMxwAMMP04g4/1tgyXShHVhyZEM2ow61+hzk+DlO86u
x3SiyOcuNPg28J+Qz2RY2tp4NfMvtpbhUP6qq/1nwdwvErXJmTKbIqsqYvMoSeyf
zsD+EakFNvxza9l443mTEDJ47upTPH+RBcUOjQ4YxkEf89kh2bTb2ZPu91DVfJiy
3y5Ycajs4IWVVFeaTEXyd5ffS2M7zEZ3Pos2voCFxbD5bedxPF0SS95FTHkSGugt
TynjidOhOIgJNunuflRGQpPJXjVvq+SIb72uHLgwVUaBcFXgLB8O8YtEAyWD0WDn
U+QhNA42Eb435rmDDbjcMZyMX3KLJCy4D3Ejbin3Kgl/SybwkMZ4I3Rh9obAVSIa
MvA1scxDBNZCK5HJklR7MAGV1blvZxQKzO+L5eunQbYkcNVTdZVIEcWuFhUnpqWX
Kb4nWWXgDTtgUgyOWleRnZXk0qzAwm99VgYkNa3XUcQkktvbrAahRhugljSwCucO
lubYRVcKSKaH2hpZAOPH0v/QZCu0GOD5jSrj3UJrlJnM88MUsVLPf3SqYu7ZZlMZ
SCM7bY0j6O8RoGJzgeQEPzxecZP4fr1SENovzZrcM8Sq1bOW7D5iZaZDVL2gxiJu
gmiiAQWpsG1p+gTduvJnQQhqwcz47Ph2v32peHCH3izv3q9eeypgy2WV2K136b76
`protect END_PROTECTED
