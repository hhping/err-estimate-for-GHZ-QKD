`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sg3SW1a4K/4pRET5k4I29YAe/OFE01dyRge+RyRmsXkctdRI9pVO9/vYd+VB+LfD
MTQ34TCxl8fnB62uasccMLmt5O1h/b/M3yHC4+BlSqNL+j/KM5g7UmXWfF68to48
8fLllTTI41dwj6GIpcLu4eir0GBL09RApt2U7QQAEkDDCQNR5OXtQdAP5zJ4dAhr
vpf+vpOHnPoIrjV346/zZ2UxODPEWMbwSNwCigEDuXI2gwhglPfkvxk1mVhPTzYw
/Wcd8EcMW24OIUnYC15TUILEk52x3H1p0R0MBy6QCdMkI8b/a/PmCZW0c8UNKjA5
SM3MBlkewjaaTBhwnh7rrnwEMTqBB08ZEoIbrph9EYDxuR7ab13iH1Rc1zjgQ/Hu
5U1sxnW/4tw8q2riqaDpPt+4Mx2DwD48cysUwGJGKoueHeySs01uDNG83+PlZqfT
Q3AtzXK82HWkLjM7aEntrUovf4zHCwBzf5xMG5nNiIIo94f1+hochYmy/l5hrOuq
4jmjMRsSb8e4uNxQbwhmlmCpUQp6lvAC5xJQPLzqs/Bo+gpFiD3HGfU3kLM0Kkij
3jy8gLCeezruKMgnHJp3905AMCxB1cNO2XT002Tan+R5TWNXXs4To4I39kDrgKbI
kdnNrlEn6TP4nF4Sff8CSkmpdZucU7nZgGmdu4HV0T2AzjYWWDKwf7mCA44MgxFi
fIF46j51pVDNIgT2ICC4/PknkfgAyqvBk6r7j2+GFXWXuDz1eokFRYN5g5oEzbW0
0LAsi7dTGgbFQtS1ekgSjzxt6zeEDg5xjWXHQSvO0JfzyiFJQB1U8tqNkYoXtHgt
Ku57cBdFI+wBQ9xo7FRAwBJ9YRIX+Yw53gqOYsMyfsNxqPYoJk8vM/8x0L1AlSQn
OS/yZmRsczoemERtXNAo1qU5f1Bts/mMBrDagZYUtHk5zOPKVxagqSlKKF76pk0F
WA9TpTReuqJhRUwjHdSGEOUTVjuT4ogUsjXeKrPck5Lv50dImsR4K0e7wsTSrMy0
5/O7PleN3h67emYP8KnkrPeujYgdpxWnkpHf6yJ0wS+rAVOCuqEo/RHT7xT0sMHr
LrbHHgBsNaRpnBUyFiYTDfBtpo18WIlz4pwjQFI16cQf5fYAoj6cODBk2PCsAJq+
II/MBETKSMBqb1Ky2VCf1R9vBzDKPe1qSaQdVQ0asHh2/XkPqDsyI2s75KsoTvMt
EaeGTJ7KIsY0AGAH2Z8GBOyMy5ZYZYDVbFUxjvk0pAEAdCJsjgxr3Xghj+8kSxKd
qSrHb7Qe7LPgWV22aR1uJn7ba7iDof80kdH8N0WSD5efxjePE60w45eD2Xh0d3NR
yPSccQJURk3n1hAY4EJ3bAxlatwQv8ib5i9FWb9B0ioGWqKbShWC6neZUBHyQ/pz
0ckDUYSJz50fdet/Zx/GbPYXOAyLA0oC2JsN8KaoY40vJ2+a6yAEp+ktMwdJiX3N
WU5Jm2J2jUCkVNZdOJFGiIVhE5Bs8nW+5B1WqJqFTiTaZBOuQraKWbT++Bn7M12P
BnA8oSDxBfWkuOPKLDwBnA/xzWZPLXa0B5o9rcnwByzaRAKv/87F6ILpEcsb9nGw
uysYsRWxNRVV6XATjeTDGP1I/zwG39J4eDymwx4/7gROKe4YHnjYbkr975aiPsms
3KH00z41QVeq7JSQCjz/Y9ZClGItCjLGvQGMrQls3Vm3dalggMoBhTk/K7CVTE+D
hEtwe+EmW5bRCSS/cWAAms9fvxp3nf+R7OSGTKxtJRbMcqH7WhGWwBsCUudoLXmK
XDj/o1eHOIZacoCX3AK6CWINMSbyDt9jsiseEcclsjawMrNiP5mjTHNdsvLtaTQk
KBJgrhQY1CK2W5EHQrm4asuAeL0Yz+0vfnsNrYuQiJroXM90m8adpI8aiQuzuHSN
hg4418Z+SQtXpXJYxGmyTw==
`protect END_PROTECTED
