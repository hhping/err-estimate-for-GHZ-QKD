`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cMI37rhk+pqoVD3mUmiycMyZnKIhxXiCbMuywT183H7RbHUGxUC75R7wIM+OnBtq
fH+pyOyLgdIf0v0TEQiYDhSOqUqjlZiJ9ng9G9aSOSB8PnZVm231GBMIDH7qgAU9
5q0rB5RrEHLEzQThkHAlnK0VTQNrg4QIbfASTViYN4kDHUQtNavb2vvfW/xiX+xh
Ya3yNrpQZp2cOt2OnOQvWId6fAmiqwgI77wlfUAqU+PfF9UL3sECFKS/jSdw3qDF
IcwD5dQJiqpM/EKW4YFkpC4AbEOXq4aXVDpEB5leOkoQmkXHk0W2aOnhEyqS1ywX
MzcVIKxJD7Q+3iXzaVupZIot+WmDfC32GgYkIjZdrcB8XuUJ9OQyZN1lxiyjf8G2
WnnS+fsZuHI2PxhLGmjUBdZZKIPXYODoSzGkD91PhKjH3LLrVzdUYR95GDv5WIBp
1zUnOanpiFZUx7wn+9OCNkOtvRC5PjDQXnxD4IGi2as=
`protect END_PROTECTED
