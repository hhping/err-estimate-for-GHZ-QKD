`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lPpXgrK+X1BHKiEVN+bW1IIdR6qHDRizCtZSCgA2agPxaQt/uCmb8M7I+QYQcKyv
0sPfXIjEVFmSaixLrb6xTN31Xy9x1D8YT9fh8v1bm3jmjalOec4b+FP1MYCMcTIp
GtTiqHvhFwlhWG/NfStcCCPP/a9TFyhUG9uzjHl1dSpGJnkCPYBgaANGQPo/3o4a
EquTWIfwr8sLHAJYKPV0stpshPgrKH3KTZJBuoKAuy6p78i6gu0qhuV52+0j0iXX
e1zm4SDRy2Zt68y8I+UQoxUFOhCtR4shCk9Strpzyy/HmEQtZCn0t9/29lbKd3iN
bvbKDr2kxScd336BfYYqNWrxlyrliOaGFbD7VuQqwX6vANo+rKZiye9a1bRYO7b0
+yq3reuvBNFLFBP8P4V8jCZ1uEpeIkgvl/ssdU+5JlCSPHB65N2QLbQNS+8Qy0Km
hF3Ta/7TTTM7a+sVbxRURKMPU7wkRJaqviUd+wTq80OzWXIUa+f1L9lNictUB6BS
va7q1csPnbUsAi5GD5wVCM9P3SxfMt3jcayHcpq1nSafImdLO6OQU5JSd1tnXqOC
uoMa80W0LAFFAVi3udZTWHPvMkBHxCv6nV6HDbguOiOvysTN4G4dCM9wZDfgYsRz
HIq5uAyjwtwq9zGQ3FPbpjS4rjJs+f471xQ8+npVUJBTeMNT7b67Og/xdguPV5ZD
mLjINLMLmyywNcaJO++iS23Jor3XOBZnqbM0IOiLu1vgxdibBg6areuIip0n8PN8
bWXS3DgTWWR1QTf6uv04Yq32HTc4H39fG5ih6+Mr7Nhn2srEelV1xfsxcVOx8/AE
EomfaYDjMfI/msrzzKh1BMU+9JzufQVxIzwGXQuE5zttwq5T4AuyY6kTDmxn0y49
jqBjKxRYRJPX8TNyasyDLHiBD/d5LvVV3cc5xvoa4fTmo3lp+DEHUKidBEc6gvxJ
LxBa8crDNEffLc/32qnyOkKT+gh7KMSXkTNFdyN+xnZPhvl9fPA6nJ24qCeutXz/
7zZvJV3TwpLl5dTF07ql9BeNb28FIrOa+p0KtwMhnzkLBZG1pKRQQAOJBh52MhUV
hs2zo9sAHJgR4zXXzqzkd9rM8DrIWBhYHeoLj35a3lY5aIxFKpqxh5TqQiJDPPhl
KplaPnwrvkXfaZGz1za+Fxw/9MIhgy9U/6B0T2pxMXn/dVfjvWNKFXdvnoVcZ0m+
cYHpISjSCZ0pgJt5vEPNdT9QGk4f+OMfd0RfjiDTrSn7GZmmejiPY1nu8BmkTmGz
p1TF6B/2NvIz3/pzQD6t5FV9DPwpM9uB4Saa6ySLRCfN/tYQkpYwZiJsLR6DFt0k
zltF/pDPxrxKjdxeJjpp0FQ4ZbBMLkDxLZH7foN1Zel/ojjAF3QaKYMVqkCJAiGe
uotjmG6iF40p/UE01o5zcJTxIR/i5QuAGW0hgf+/HnOP49V54oNj5reFr6sRuj5l
7npSfwN3cE8leW/9Wtsamwe+xgxVZLNqK/83TiFoT4T3IeijG9iUy24EjPi/EqZY
xXoxzuv3qgeCsz/MgUV4LXvsEpQCEqWY5gNMFsvyZAEJcvNGks3m5wFB0+AtXnIH
NhBxH+2UfTznyNVFvZEUaS7AsRspkrkecCw3p3riUE/SHZAr8MfFcD0Hras0PjoK
IaPNj7FSy2RIZaoUBw/xuVaEieiNOyVBZJ02t16Fhe3Ukkw5+tLxqbv/oURG7NNG
XvxRz6V6+y9U9bHuIlxbWkDKiLDJizQPWFbpd7qMFdtwJIaWrWtVAlRzFxX9l6Nj
SOXLxrWStdHPxu2/BbWuPllda014tX1H6MVHGU/126Z3Cl3cajc+EJDoK5/oMKLp
bChQanq2VAttaKrFrRe6MY2gbh6yTitwWa9tFJbqo/SP75WaIa9lhz8LjiVrFdVN
5uIgr5oA+jVW04FCm7xONgYD6uLEnWqmGBTQcl0w8hThun3BKun8DgLme/y2VcgN
aEwMN3VsOt7W4z8RAC7QKH9QMY5D6WOEG+gnpHnxUOiwTbt/abI/StIdDmOFLqxg
d3uIyapqPmnp6aasdaN/WViXy+rgBSYptpbOIsH38JdFAsygnQO0ZBUoV3eMmq2L
lZ28b98hWONbq2VAXkDmRtnTRClgvJ2I/KqrE0hYkdyucJBV+Ny5ioc+lgpHJLD3
tyeSH0UDAgP3XL7QNXNh5lmdugbarniGO2T1/xGCtfhPHWmuIzman6bsRMkXnMCJ
sss4VOcZFjbGw6oHuPf6bMjmXVEQBmobmqEz4CTfQ61h1pHFPUCBzMHGkpYp7Yrj
Ej/v2TGDTg/kj9VPdJPNZj1EDij5zuMggGsfaQbt2SuEFrFRUlWJTWnedA/IS32f
C+oNaKtXisGIbz7m1BQBbaAC9YYnTvJEhes3Fe2XDhjvzxKIXgaxJUEFoBflgATD
yOU5fFK4eqfXZbdzirisTf+AyoKpwCnofszVQ9k5G092Rnyk24+1aR6p4wiXyrHe
eqibj3RwAu7h4BhJl2WjhcA2acgaBDmmKFA1IcXBFpVHwWf2pkabWKaMTTktWA6E
`protect END_PROTECTED
