`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UIsezV0WZgyLZOlGtyui7ufcc1ktovr6XX2el7T4nDqadv+olfHEuP5cJIpm/QO8
tqaD06/eeLDxiPPK3ZhWmoq/0pFg8TrPQGxcmRbiYSQIca+QXbpxSNHMnl1DWA2m
Y6mzC3Hgzxr8H3BqII3vp+nJ7IT4bsS/a8f+YTWq0uh93AKJt+bMdbmNgg4IfBht
lGs4NbiaOVT0eRoUXBxFkpkrNWqYfKAo31vs5rakoRgBzLw+T4DP4o3UUTWjh61A
T0xWo5kFdobe35e+WKqDVCopf/+1KiKP4iUGRHnEl1lfh9gxwjrzYCVONNn0ebDf
Ejf96S+k6+DRQ7O42zs9RsuLnAKd9CkNWaKeqHIjGuAhXnUst4gzHMwQVCLjPc/9
t6Jg8Yk5R6dvv7mmhx7h1Rl2K2RbJMwI7ttkL4GXPm07FYCbOAlSv+Hzso9rK7xD
JQPntPZXqQKPW0tI8zfI05b0T2ZhORGwzS7drwHDUdhsGya1qK1tFgrW4Be2KBGF
MAxdavLB58JVTINBQIcx+MiEGyvXVKt/pBVLPjArAv8fPZy2jc1iGJYSmWWOFDUl
xEAJ7DVx6scmaJwdM+qURpkLpNPD+RQk/8kd2hol+ByTWsA0Deapab/LXE0FmOUk
BpQzH1JmJcUoXjmUvBtUjzNkH9oNAqqaOrcfqwIR9jCY3qrbjXf+j+754qKHeyfb
/R8iyOCmmBWaPgSYdQH+mCJiFsQ6L/wmLW4cD87bKh7Fu4xhLKlrKWV8yIScJGr2
fRV/cRE6vvNHI/5C9GID43a7e3tRroWi+DpOxqIpC/JU7Nx1CPMPC/UXgJtS9fqR
`protect END_PROTECTED
