`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yC2yeiIobssnkvY6/wDiRQDxOpwxqlgwwcvQmOJhiSgjNFnY2RE38xeKGEchkl1n
Wy3bXH2XXeDKEPHhasVGD5VcllQnTZi3GMnwmltZN9cZNdLlNmpMdrHEdN6dzgSS
N2shb5BNweIh6JADSi1xmgyZ+9TEZmX9rB/MgCQqDQ+ntEjlAUNTBSLo/csWDpAd
XRBL/dB2vIkqvQ70WEww7fqZwmRNbmv5tuiDFwljFYCtag4aSZCMR+FHRbwz3xDR
bZOnKIimLb0/eBaCS6AWOoOT/G7TUFYQ28wixgSU4PuBMEM/oORVHN/aMYLOVCXv
wofY0Ka0FU/u4xPQjGZB5TUIfUtwOuz/PTM68zn7VWx5mEB3jdXbApl26sRBAQqO
R15BYG6SsBAxGnFv10izSj0sYd4PAEAsKCaUI0xlOBOl+NoSKHRrRVCoecy9Arym
D/5yCYE5c7H39yLzbiHbhUcS3wxhrHQKjvb52HT/Vn8ou4dkKHb4YE/EIBXWk/0i
1TNc8qG4HSQeXdxkGo64dLs7J9NnJgoXqdGHvOr/3L8UByp7o0d91SLgO/kF9I1t
cEiSfWIwiwFX3QMt9vuS7NDLVsyCcQKtaAz/DMMcQoqe8HTARZMkO/bepnNn/U4i
exKnzO7yru1ohM+vzgAk7FuMfKzTutfKC8CoUwnMSEvtU6eEmlyVykcCcVx6gDP5
71j9kQ9rS639HjGyQG1B8JBt8gbYvNMkkdkvkN/xGCg=
`protect END_PROTECTED
