`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5/Wwr/Z4othcKC0NzV9M57s8phorjvvaj5ZYrGHq3Nu5hS7sDItT6o4goojXxf4
pPxNRxv+UDjRZVS8wb/zToD7A8n5XqlEzqxIwS1mS2ThUWdnBNsFtE0S8vyDVaCl
CN6OqPXnvAcmtXC3B3p+2+s3F3++bFpjSonM2wFLHBzy0ZmMIw8Pe68kXjnAvmQb
xQVTicUtIa1EPlxbaUZ/tmFu7cznfccB6+P4rSL7Z4pMdMeyca9wOyI0bgmJkGiq
1abs5jqUbfnCwk664Rsq5zyAz6uC/vgOEonNMpZ7dRpc6mVCzQkP+gqPd+aWFjoB
SI9XfVeTtZnSV2kg5Q6jU68wEjBFO+kINMdkJfWMPMmdwtcgvXxt0xyeMK3aUJv/
nVYWi3ISPpSptkiaZXoq8NT7HUA0eUCihL/ve3imh4CwVfmX7nM/PLID3eptqGVd
9hOUSMPFkTjhxnAapXj7ZvamRtaonsllBKTPtB+IyH+ePH3iG8i/WfdGcArsbFjt
WWo+nuciS1I6QH7wNKTPzTIo1rX2XNjuwiBWKdRMQnV9SDrAEklRtEuqgfztGGIS
4oVgzdGzRclsmDw6MYbpSgleENltTcvVVmgxFiBMeisrNmmnzRXqG6duPqfb5CpB
26q1Wd+I1gciTo/n5IZsD6MjRW/zqWmTZ5F3WejIRyJuHE2OJyN0iNdcyn16For5
eOZr3MLxw7nGCD3PB9015X67gcfoDJqvwZnonwjUvHXK+wsuEhP43LsHN6AW++Hh
RuJUcWXfgevFmAyvlkR6/cJLWDcx5ZPEM+mGdI6rooJV7dBC7nvoDxo91G5ItV+F
`protect END_PROTECTED
