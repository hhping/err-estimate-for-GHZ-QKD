`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ylzidpdv5c/eJUoRHOZ+a/JHUipnlDNWnIJP5aTk693/12PJhEegOWuZAE9lGKD0
0wv+PsOXZ/D9Ub0SaAKyh7rjY26zXPNXdo0nZobfzWXbahJ/P/2RzysbpbJIkMsc
IjuV560otfbSJg8mMCYgiwaIHmJalcwflKBJwFNfj+Glq5CkONYKZD9ds//aVrfB
Yizcji0zy2rTo0dArKN57lfeC2tRwe3WnFPoe7CAJf7SA/txcACi2sd62R+aeLoV
1YFE5Wrr/pzsDvwUZLPWt+shJcZgxcsepT606PgfMfnUBJI8M0Crv8szRDNd8/5s
dA/q1UP+Rqs9dukAEXwyrWk5wXIUgToy1WwXOPivGe/S0v/JUbOkroEqIapXgkhv
tCKEHO2hZfiItMJBdJfiGqsUBUatbSZeX9s6mMqX8tjxQMGw3oeHBnXnrV/1zG0m
gEZhX6JcAEYKu7rbeDJk4OqmiNTqfyC/cbtB40IJjIik3Q8PGnTDizWHSOhSqV5n
UHCfeflXk04ueFMBK9QVrfOjzpoqVh7eo/SLAvxLVknkjFUJOzTZqwgfeoQ7j3id
YklkBRvKxsXwksKvXEq7qiLOor82aZUpMzswkue05pntQRW7Ax8DIqh/MSx6ncGG
cMeE3utCg+R//7OyIbUK/6j9pXS83kiOsVOfxBQNIk9yrvzYrojj4xN5JjyKAwYp
PCfcroOmN1YQ03uvOQalkRRGpLBbrLvOFMbH0mYioUFS8oskej0swOabNJNWh/dQ
joTyz2L6xJapiiznk1wlQKwuVdSldp0CCGymEQ+dLkpofDndQZyLVTfeLIuQgRhi
50Ty2EYupwhHMkgtUOoGreBxo009GCeMZZ2FUd3SuqWofjVNzxH86SUV9vMQcM79
4ug1SFLIaku6SIu0xw/4riN7CJr8H03kgrYRpDzOPrTTut0bXIg/lwGQyXTKCaPR
BFXA+IwR/lH6YDL1D+s1veKwrEAImy+zKL9SVFubcKEAZSrGLdqez5YFEwODofkD
5SE4iS6odj4xa1S9STANguUzZNBAwdj9SsQkRkmg/ABHAJCkG1aQkw8ejw2/6u9U
DABKke/Wmu8GbWqZyRH1EQejv8pfQiolLDWzHuRPR1a3ZwQqvG3Xqu+dym9nwil/
SRoV2TwKjIfW9DdnYXCc/Yf9e6wF7+cYE+fN76NktL50mh1kyoiVq23/jW+Lx8QU
D+xftso8p+VZw6SoFbRKYAdQ3zFjU0fKI8rs2wlMAWY9IuT4nvL9rPxgUMPoIIYY
cHr0whV+yM3vcbSDhHpgdXWGf5PvgKj9jbZsCpNVpuLKXVWLnpb+/7Mh3s5IgN55
0hfHUXnSJ7dX4cE73xK3chAjS3W8kOjsmrgRWHXzylT1/+1lDzrGIuc03599MSxw
keIIg0+v7xWtPxOUx/2YJEqk2blck16xnCjD5jLvVzW7xZpPJ5uWMMfGEkvGyBA6
51YOnqaC85lBI5wwMM3OAPvlWnfPNLhEOkscQiNspPPZc5MNQT9771x25N10CQdQ
qv/JER5XyT/nic1QiBYxFD9X88/FWIzCPZ1YkpgPJcSqc0yuHK1vwwebeTB3AMrL
tlnVzSOrD7OPyZ8uYoUgJQUILLUZKdX3zkKk0T66ONKOKtUXUW0soc/Yvsy4aEHd
c9A9M+uDYBBX1+Dv4FRDeiFLrpQckOi1r+mH3nnnFRTtLHwQAfKLBz6bsgVnmx9P
D1NGbrJtQmgFSMmWW0k2v0Yq90R4gB+Wp31jtl4d/u/ECc/8ukmVhD0uivDQRZLY
12FZC9Yo0gvsS3di/kI4A/CZqlKzCV0yjd6q0toBTgB+rv7vvs92k6d/exmMtaRf
4rBNoxeTOSrenxM1d9RRE1ljpBvnSIz84MPBXbp6KVhpFOLPWs8e/9i/C0lGqEoU
9DADp3drSzEptqo63O/P8CttszQ5SUriTaDi0wJGDr7MNhDasLIB3GOvKWfMZTDT
XoRWI+bYLoU2GDORLr7oc+wU0HwYinyp4CXUWZCHGZk5NED7YloJ15YT27FpQuN2
o9W91U+2V7KeYFtS/YP34DS2mKtf7GXFFoRpd+mxfnhg5ibDjOsNTlphMRADMdHr
hv20M/FdZQUACt1bsxNA+Xaz2AM2pTCuRMls4JJoMXU1kSqDwlaWDG+2D6PpNnTH
JzTMG9UT06Db+dcdwRY4iGeBMoJhddi7GyXnePXGQFdHQP6KfdKiNsU5YvXv3Wsj
jldMsybOuK5LR9oI7R8oRRaR3wnhHHM+KpFjDW2/2k+LU8jmBcYjJAr27oeJc+eq
U0IJn9wQO0UrvQIhvcYVO1OgyLxKfrjywEzd/iWROtu+NbHmMSrMud1FBPRfVleD
/KfLWf4LFRPBPlnyX0F8y1aFuCWpoCRE+3zg9GUTWcurwLdiMkxjPXZPllY6oJCl
m67nnTDel8hKEkTEcoaFb+Y5R1nkevjffOzri0xgE3M5yuaZYxTlvqalfbUANBC7
hTkgqnm1F+KmLy0WTQ6UJ3mrg4bcc3mvE0jvgVGeZTvOOWyDpdxY0CbmD+1Zmzfh
MeZ5L+fHBzeQ/ldQmBnDKnxxzATMLvD7miE7I7JvWwotp8fcBCaew38GtRQ9lmuk
PTvVZKhTvxH03pGk+oIajofK31NEsBpxVmJEjsYmeBj+KVSXJpVgl3JcMcT6N+iU
/s8pz9V+fTskn66oRycUco0b1T0YKC0umF+gty2EBfyUdx3YDRHvbvs6KotJHy2y
f+XybwwkIfdPHcLq0TU0gi6V1vpJRDOXUhOFcGDQfGaZHXihiKP/ZAvWwtJyqHm9
v7CQuw3ecC36zv3Pj3sLdFy0t3WgRR4oJMicsJ1s9JMZgxnd+ixI4m2cd/HZaVli
rUcN4jrHv1r4WCQVYnywXeKZQn+AfA1n56XGJ1JjIXxx9wXB4P2LclFbjdqVSzCB
OshHM7bKTORwhFk/uKDt93WU8FfA87E3Jdx3UuVLCWKuHj1oyFZhOcgft+9ztRpm
GY5T2bYG8L956ALbvvkduxkSA/Oq5t3tQuy8zKPIKgZYcJinl508d/KHXdLZ5Hku
V2X9sDg9ePmWPpCIUr9xUYBNxlfBpZinGU0mcN41hOOW3c6mEzeinTd8YfwPwjbj
XJofi15MvoSMES8OCu8YxRLhrESmcn20gie3dyCWVeYjMyJs5SYXx0V6ppe7rQoI
JrnN2G1XcE/97OSWB0pSYMvrgJr8DOCJzuQXadWlIIFuKtcKrKqT3ic/1ZoITmf9
vt0bRz9n43dURpmYEbAOAv1UdI8e/WFumfyapRzigmpBWnhK7Vk0eCZXQ4jAJFid
TTBcH1cSKjL+14jB83aeWTb79gmW8ZvTv/2WJ2Mj1XRuTtdodJzoZ0euz97Ixnxy
0VV1d7XT//+U2yj8zjGTBwffJDu+chglvhexSZszC9dshrzVpDSU6l9slmUcumTB
H2efMe7JMXHxpxt1/n3ZQyzsKL/PeOvrDWaRYsjMo0xaLC7SHfIpMsPngen9fJwQ
OEoe2hYVlQR1UmIIlsDiHAk0sl4lGhgdl23N3yb4jnw+8siLvrcWGm+mLwAs94Rd
Ghxap2NtFwf7sBT2Vw3Gz+uzDCnN3mGGBz9PlCJZnVCxbMP9EVG5xstKLK2j7dWS
SuDj96YyNwXUgL1A2fsrfv8dETtwwdMgdQpvhPeQKZZHcDYubqUUJjNk53HpWXlw
UN5oPbD+iHAost/8nAnOPsqWr1csIho8JFiN75P4KNmAdhGTK0N2hszGdeEnQPRG
EydtteGRcuBNUpuyFIFDHazccRuwgATtxpME871Mp9ufezZtds9qlq4BCNj9xUF/
sxjkdx+lXJeytYzmeUsKQWFxVNqkurURTkh3kglHXZSX4GHcfMA/HAW/z+eqluEk
sYSxU+0W3O7xYxM9evBnjvgQkhTn/VybtSt1mHINLx1uf6p6AIFX8cKg8dfkJ4dQ
U0mxythTwTKMY0WaK1sfzX34IDLc7sQZ3eIJxiWiwy0f8N3oVExAOASuTdszwQYq
cqOjcZoFrql9/hKo8RnhQPIlUNEcQvi63UKfBb/F9G4fcmdYVJiczdFNk5EmllE+
F3ByBc6Vvkog6EH3M0hteJ2B16Limm3qXop+EEeYKN9OYOvj5yE+BIy6hR5PnqfM
Ajnf0o9Vmcy39aXvrbGcXgfZXrdVrmSInWq+PEf13M1wCSjyIzjUxlDR/bTaoBq9
7fHvuFOj2wClDl1wdbSCkRzJXHbE9Mp4NHATYzSc6WRFkVtcNrVJnrVgczRkYFHa
QRJeFbJTg84AP58rsuz+fsdQmnVZT8FQrKAkTdEyLnUCIyWOiwUwbK99Re3qcrIL
/SxvNJga4J4TXEC9xvtZg3i6Z2Zutl4Yod9Pe9WgNyYmtgGrP/+ss5obd12dFeqG
egQiKWOMh/kVC+73glFIMIwBFYs38H8eFK789ABMVQZ2AFITLLZBaQlfJBVjCUi2
a5rwxShZTsDS4CwDr31V6rYJARTIGjoa0od0JU3fVpFzFLfUvPQ462uMrO0ibIFw
dIQr6wUG2e4pDNq1L7A4h0q45g/fmBY+xWkeIVGWdaaiU6KFXhmrJGesWgraHjWS
gtkTH+Gxq2rwhgJAFiEx0ky5HiooLe1KOpSHvJmeruzg9Lf4M6n2W+/PgEC0s3JX
4LhE0aML0cTDMWkkoxVWt42y6148yePRJ76Lb7wsRbC/Vtgy7F9UbTmj/3ePoKVD
kdCqACEqBH8nBXK+SM/0QAMFuGoIBeXQGj9ThUzxKC0BFlX3WRWUgJDW0jx8pWSQ
nPrWXZhNCRpMkk3GdkNxmEm6aRXacRHq+q+BAOGv+LvXfm2Uhed2af4XV9Bsjaw5
/sZeaFl6eGXMdq+LLCiKxwX+RjRZd2RNQKW6ViyUNt6i1v1aU0L4TgifetRAQoHx
BvXKp3Se9KXeVc5EcL8GrzI3w6mASMyhdShhON3BZmbZbLacmzulM2J8gaql2zpv
DvD02U6NNhZbdlgPVy5CikmtZilxaooz7vGa0ebuS/GAwaHoK1ak2huUHCcFS18S
Kr3VnFcSmMUUZplEPvOrhTikScxZkzoL/WJMrmWqAA7CapJH/dksV8zq7yccGVHa
xfxeG4ImPNrvlr6iOtJfJ4a7SJvlpVjI42YJzFZrgbaVfcm1GFw3lOoLtMGEgDwv
ii2l0CAJKgqLheVf2QmJpYRRmN8MN/mglrn8yUFimImWZrDLbCL2SCHkvbFvIM9i
gglbQJjGrZzoOtMc5OjGH6X6jE1ZYG+K+t6My7axRDTlsraYxuKfblMHO+9sU5Fo
1bl5ML5q2rvL24Ob3UDWatEGvPFprefE3zI0H3+/uxlJMTPPeDDJyk1cStBAub+f
IcMC3S7xpTXUZLzaS2NoQNE3HqIyz1568AldKCndPHJuQof82wHHjCL350W6N/BE
gA6EHaZFtkVQcMm484VajN4Lmbd40IzWnIl6USDVxPWHXwCf/kyWsBadLyK1WwOB
GS/piKCkIykhn2OaxbwL0j1ptkGL/WscY+tAAylOtjM5PE5BbezpoOpHjGdh9iwn
/3oVz9TdnP9tAPXy4d07wH6bJpdH0lLqGe3ToE2jcD45X6J8IRP3N9EEbhkug8G9
Bb1dzuggCLXAiyLK+f2P2trCgODjOoXTISdBbZjdzbEOacYpRBwH0nsHtD/AtnQk
3FAZO9MTYZp9S8Ujal4LM+P8PpDVL2h9jLYQoWwy+xhm5sc/R7w9UrkgG8i3vGoW
Azdt7l8HJeKU6ofcBV95lxcD5AziMasdW9QJQFrBfZMnKCGKl87A4AkvZt7vbRBu
x65uI1IoM8aCcozvb8E4px8iywsA7BypTf8YWwJbknWCJp1tRsyR6sAS3Ev7K16I
FPuX+MGTP9BXAl100d+rEb5SReS7VM1I0DV8Sy2J04iMdzehsr7qCBvkv5Y9rb1E
JRBeDVhQVYkkangESiJgcILOcgM/eBzeyBIebtzwUIti+56eK7cqrhPAr64OIzTU
E6Y550aOc1BwRkXIg61z3iHtDeYzxGghcoPp2qE7vlFfez8QS5rRCWcsNGcJSWFj
Klrl4e3RaA4oQd2bvvgd+QfzQiRMziUxS2WKZmMGMYsKgtGr5nYNYfUMfvIniAlZ
Xp6qKK0pNYmfziJn+hI73kwyu/dwBUrQSbXyRKB+ugBvVwvPRwFoh+ayjtM9TYDW
nm45MlZZeC1+Zys64ULa9mxjjb7snwZ2MlTrZ9iZUCq0LzydMHpJV9WaXH301tYQ
P/P5u7MuzRNciP1QCylfc7uuQnq6DfHK/TxbPARGkTsjjwZ2m0YvlibkiJkBfGuK
KJELYUazUXiOvnWzDd6CGPwe51lR2PZm2yEGuVv7yKHyE8d02MWBzXxsJop0wQkB
n/OXHVI3c4tCWJrKQXs9N5u7/fluOsRxkCQn4Zb0D5HlNvQjTzZ0v0Cb1UhY29ng
XMvL7XKNCPJRv6MyI92eHebdD4lIBvtVOzjD1JzXZ74lZ3Ug4FEiLFm9qca6Jc0n
mt24aXp3K8Mczyf2zWdqCepjKJer+fm+6RAMUF5aNJuXDawUGrQbDb4Gnm5RVPnh
/LE+vegsKy0WDNt/AyJoiY+3WHmJgMfieqzygTCEP5zrjN4mZJDIfw7I85c8XiVs
eNAp8wCVHSSb6AzgIVwyu3CwyPcxnP40qYGol/mk/szGVAmOlQpXd7gtUyiR1LzE
cHwdiKNI1wJ4LUU5fHbAF7pJbQj2lFJ4rFUp1FArkXDQjZ7LpN8i+IZF2PPo4HUJ
hFELE1n8YMPimHMS0D5psOIWHs9+ryNB3z70elIfPNsYeMtKJr0EjQ6JyyR3s4Wm
xD+gXgkvUEk7Epx56leZh5lO8nxQXQqivKzeezf/8p6JxZdjMEsJa8IW2UUPO+5l
8cX2u2905MdneLy1lb9xjp0zG0pE5zAvPZBdi/u8gVSVr+T6BNpmy/KnztmMjlaW
ZMEmcYajxx0rlKa9BVphGpBDJ+NpHsPML/oV5YEkixpoNvsT+xfUOWvAR4xjXUwK
9NySic2Ct/81xW9e6QpUBj9EdsNSQhaZAsEcfHhT+uli5XZ8H9Qb9vP9Ycq2xs+C
mBHhtd1Yr7DdkS+QbSvJALG8smeO/byXOiSYUXlT72OOx9sYYx07pibx4RxrHIpv
hP+pMXyM5nNGJGCaYxgJq7mTxMUGFXgHymU0rIezu+MLNEJvIZkUJeLEePpfi5hP
vYF3KRiLIeljxDDOT5nPU3gnRcwyD2Z58eoUUcF0JK03emopH6LpfbTPCo2S2iBX
FrTcz5phGKauXnMyB0Xee8tG24jT7M7h4O9V0zDAx7RQ6o42OdumY08uz0ayjGSC
lXrZBP5xDiFAX7qaLwEv5iu7xjUeyQB6YpUEmBsQLBSwWIxSkfDZkQcroEgyx/bQ
lKrxpE5RVsu4k5My/BHy5yi6XVxclkmaOvqPp1ZBDBYlTOG2qpF7LVffuQooaL5I
7PqF79ExO0ayCsmD2bXyexTv8xfmAkIOkPT/h6sVctqswz5cKMyE7HMGV0mtXFLs
YvuK/ZEjIHNtm8QhQmk02zgceUlSIuZ1LDp8ygZosYC1bTTP/Lsh7kFMj7sS22Ec
xeZYUXTBNDIlUJ4+YjIHKZSY0wC0SaSJoittpk6e0tSOJ133l6Rln56IHOUMdTUj
mzUE9nrTZ67Z/5PEQV+LpYS0KXQP96yB137mLtLNhtSlAxHq3yKRvNm2fecefTHK
dHXalu7owA6JF0UeYYdf1RqBAsSDQWDFB1Zb5KHb4g8nz8UUp1VsgJCkWUEFkRsP
0Y3KonbRKP5DosZg0WuxmYnW4qdyJXzPOrw6gq3YkMrYtHUuoAcSjL1KhO5df0Wk
VXjEGUOQ157bPsAVQpK69/hfXEoscUXj/k1RkHzbZFrq4wzalqcp0bvjYXWdDMgk
fayNyfp2oSPjs3dqHlJMKz1kygW0ILTTmU4xxfGzzUOuk+TOLsWDYz6Pyr+nCxNO
EUE7GD16exFCW+LxP2yFWipPveDibkODlhgng4GrAvp2PSKlZYCmsArhS9pkW5an
jVZEyEK4Rk7lwRKYyv34XASFbvsSttbiwEEWve7H2nU1VFtPiZ+w7doHrxmGGb+H
L9nI3sPbE03B8+4Hu53xFQ7wxZOiq27NJFad+cjzwrjK45366PfzfoXx/M01G45z
LwT5EttevHRAtonYEIqSAF/2cikK1dmEI5gU2m3r2wWcNXrZHmBiy8cnEn1dJ4FS
k9cQcdQDOy1xM/f7wIEsom8JujJyOg5QPGAejJ/H6An7b/97OCJSwE3KZtbdnRJi
bKzCRcoQDSqa8OtggVTxmQX9Qj8iZjE6f8wC6GOTihoOTHErK/e+dVByrXhP56DM
flUlCRitdxIqprk6UWB1UH6i8DuxH6tkxZTi18/h+iO1BIRevTuwF/gYS4kNF03y
lsuyq55cOblSTkyc3Pb4+Q2cF9fp3hDG61BoOO9qOwu9xTw0ZaGLz11aqtdnNalA
PnLCu+vaUce5fo7/5vVO0WSE/mo3l2zjhWVWU0Ib/zkcIuuJ38EinBnRG4IkkBFm
Pqx+nDHTbW2pwuSiYxeqAdyj1CMD1PKR82LZNRtqeQnTPS6brtomny+6bK/ZFihX
qBj/4wWAVFEvTvq/rifgzzVrCqy9w7nybe8jGl1vYxDEMJI+U6NBw661aOxhxH8y
ZKMp0dAH01duvjFRXx2kTXeSeCKQ6suOpIFhFGj4uL14dR5oHz558QrN3mWbs2Qa
1JAUC33QPtmd1a+nllTH10MkgmCa/stAlUS+7zMGofZGqCzy6CS/E+XAtJjEAqsM
FZcT61zPxOaq4IxhcXoN7mUPo46j3txGj9xNK88L/jFExnBQ3FIt2IoU95E02IOo
+GV4rcO9+rd/uEdtwNbAsXVwoDKog2T7814GofVkDBeVaPJguXZEi4kynxsUzt17
QJsTXHIH+41ViIxL9wNRsXFWxMCo8TZICamiydbRNJRFz7E6YTufSWJ53uLjo6ES
YjABXwouo8M1k15ijcwKkF2f/phHsDQrxPCGC//U3KzpqJLeyMgyt8Uw01TgY9tx
ukuoi15EqZocw4yB0tC3GkmFlAxGgB4UiXxHsVG3Onp7/pjAv/WZHUANzvC7AW8w
21yYQaH/w0gtgJtlZmx1vhEPJDChP7iiOe1H8Ym8db49faR0mf8MHAqJk0JJ5a/c
qWqM6C39cBmqN7MzsHgUZ2+bTSpdSLw8o7sMBCN1Lh8MEFd6/gOynvg0NX1rIugC
Y0AJW0ybS9/nuCdnsV5TOZgLfWw6ji0IG7bg17owKmKLcv/LCrLMyoicAUSI07DL
SLOausgigmuQfdiifWpaQ+KO44JUNGHpWVDgGBrlvzNOBgPClBrMenPIwPaJixF4
A7ycRnx6RQb20N59K4HYgtJqNOaNf+WAraRa7DT4/sgUa7DKKxP7/2tx/nhgV2B9
sjabHK0t2VwSPq+LgzZP9ipKbAA+euRPgiRXiiCLIwDASijskoVX+kC4u2x/8+1E
yF97uGvXPdyX8fU4l4b1tZYTpjY5OrG9944IQs1P3c1xS4CUI5RA00jqcu1rFOcN
gi3sqFU7Ka26mML+dz5rAI5hQolBO5Ya84uA82OiAA1bYlEei5FNKqaU7ktRSpBI
AFBT6TFUG/MUo2j+gQ3mSh4YPy2mXjYiSJ7yrlkPCjzORHtAIxyDhS8TfEroLpB0
cvioptv5wKyPMqfkCOguqL77ndiEEAjj8jPKL+xMRhyQKa/qN3fkWASWxS44gh3F
TjLaeR92+rNYjz/3Oq1iRpg2zGLFmjIqf5B1JJApSkSOfQxuCWfUlng1XnBEOjN2
KRiDLb4VYk0UZEXn7u2ckpZ3FjvU4ZGXZ49WeY0oy4d+d7NJ5TInMoWymnDq8c7b
8bhu+s8FgBNgG51XjQiLku/CYSXql9CBrIALKSP5qEXXmPQmjN3FS3QWV9yOF3qY
kInaSMTyszNBj8yQ/ZBOUHM/Ii3rttV8zXXFIJCVKXgr+74khh25Gz/4Ll+gy4Js
9kriWORp5eGW+rKUzQnOUJ292qPpoNgofSm2bKWvA+ZdrjA1teDM8N3xEmpRSZgs
kwgFBsQ9RUvqc8iJpcvMe04qwrmP3M2M3tGOpl8V+jk7d0WokIUzzqg2nTsp/M5K
dc7N+zwsIcCf6CsaaQE+gxWLM5IeGxy+76vr6liUGaUx1PaYoqJS7dPo6aHYNBVu
w8tVoXlt/07bcpv4b+UbhxKsQCkNtNmnTATR7r0lqFI9D0focecJ7qlalBXxeFOu
gSAoiIz6MQFJSaAzSdyO67lKPvm4RETM3Ij0arMEJqvTI92CYauiSQyXslW8vQAo
WbuGl/XgyTCGJRYKNA9nen7TdTMk6k9kiF4EcNdymK9qAlU6lr7vTutQx6M2y3BV
S3Izr30dOstfrhwPgNuVDzA3iuZAwEVz+zNlSW6GCW2j+0dWxmBtg/ePOPF9vIJP
DD1fJ8EpCcwZaln1MEmtpnldny6Oz9pfsuyfGtA8yhZ2ffPr4BUQysm7ZWz0F7b1
aMaM09OBmUkTacnO0r0kixVnkg3PwbGJdIkEGTPfu5R0m+IJ8OCQTIfe7yp0Ko94
sOZUlIOQmK536OWrxij92qzCaGs2Nnlzt2xkn9cuWYQ94ezEyXENbwV1nP3bU9TU
MhQmFehuLk91zhBIQqvJSQ3qxn3vlNGDxAfdSZSttrIRy3JsmJzU/T/A40PNYkjk
Th9AtauVuZMSiuJRFJR1kD9dmIt15mCRVRazLhDJSRmlwSzYAUNIIMAisiVhAH7F
UbQUx3Ewx1XaWiTaZJjeUQoP9zCauB1xP72zfwcBgU2geZLnORJrTFY81yAIy7CI
NwmmD+dUZqKwbpt75JRh+GXc5Ff0YaYUcam1Cq3iFj0lg6bUChePXx5Qjfp7I1w4
4YD5nvhpD7gC3SF+PZpUb6cnEjB3Hif1AJbf71eJOPjgPfTkoTLZnPWNWetrubsm
IUN3LibQ2TmlCNCT1K5Hn9RuYr4zy3p0Y7VNhRWZfT3H6BH8pDxwMDXXxK32bsGA
rHYV17aVikK9HmXh7y1JbT+f64o487tVKqBXD3FCyuziau9wsxKK33OHSRADcVdd
meCHeDYL2IZlrahmf80xHmBENjX+H680NjGUUoO6KLR+CNTqhWSKm0PeqmYXx4A+
0kfSFMK8qyfqEY894xxMnjf8Na8FDb9OihQlCd3vmKTIi6EZJzGnJYSKiBI3vMR1
EfIbo2cCS7/J5HN+wU3Bz0WwWK9CvePIA6oF3Jv9M8tmC5N5zKsbYoJR/2U3Ecle
u7MojLDq2aAE45ns/ZdcIVLn8NWY9vcDt/XuwzUBlq/DKGCwmkoSn3ZalOFuFJt9
rSKSH9HrescrZ67JskDKC2kG++gO/1H0QlUFvieAWhW9aTQFh4NnvrlVTkb5caqa
FE3RZHQ4D1Nrrap3oVQXa00w3h/TR2GcYyAtsPgtiqsVU4EX8T4UCyFe9k4DPvH8
6XEeJegpzRP4qgdTtP3GH9PgoBRPkNG1O/LX58QiwPuGm3+8d8RBqoO15yYbkoxR
1YgTtWQhZ7ulQMR5SePE+BxbDfPyzRrbukzQHiI7pyQGmaYpSKeUO+pBOSD1yVzY
U547SFyMKSKKowqz0oLbWLLBJM1Jnu7Xt9lGaEvLNl4hiYwHOVvib6RVL3KDKNsd
3X5QfVSiB/IUITY/mEwD0FurSnLiKiXRKke8WD5EFp1NRKqrKRBv85kimOEf6LZV
1v2m5yZXTpV3OT1PAId/nEmKHMT6IgV/WkCN5879TQhwh5W/qhWb643sdyRlpXL9
HpLyVzGub83H4CkqPdwa0bDLXvofbRQ6rltoYVzlzCdC/ftl0OMappL0wKTnUxMt
LuPYGhb6I68FBptDy7F7n2dG90olZJ9vRDFqvtBhT+z1YS+bfihuLPFF2nRy80/X
FTR+T3K7Uw0Z0XVqPUklJp0zlbPYAjJizpKluqGmy70CPQ9Meh9hdS72iby/cddC
I+HBgM2kgzaoBpIpEZ7IiIf+V8/sNwzRYZTVBbyMZAmo7kPwX7LnxsU/x+rCbFym
9HxNbIXJ8dgCXc0+nKK+jWtDvbyM7IFzhSm5lfN03vKu6Xp6N5wMErmcyP2AOmKE
9gNaZuKm52TXvVXnW3UyqxvxAEVRF8CO21DMtSz19uI/Qxn+YUzlM0r6ESFN/3VO
+AiLfFTLMaoemR2/XEvYiRLYWp+glkcgU0MOUKIqrVbCU9TB3tVOQeVxOv+s5dNu
33GCtZvk7w8nvonxmsbdP9uSZU8atYdz2DJuGXOd6TIxn7UNUuYfox6B9N92Dzwn
78x7nSV4sal6rr5kmJJFIzXfvFDGjyhrWnR2QGkK1aDXbSP+EVxWT8wJoLaU7QD/
DK0JHFlXqAIv3C5ym5mqcBXeqDZBtdYheeUEmIe8ko5w9qplntx3bgvdlJrsF6dy
kxHXrwLfzM2qk6lbA57VPvQX+C4YSEyv/N3OA+7Qfua+W2bM3qiE6ao7dDXvHxsC
BR1f6QvNTITQNnrJlSm3D283Hv5t3O8R3v5BtTqKdUu1Xvj16xSCNi4o5muykYlk
Q8IQtpu3R5Qene9dg7g44HkDElOhqaDelcw3QB6Rm5olDqnx0+wNrDdJ3uvU+xdy
rO8ivUkQc8lSbB+pt7nQn/w90Y0wdqyYdAal3ALDBQ/84V20EEvzT7GRJ+W9AGlk
N3bpLqC1iwbPRryz2vyNziOHPmXOwJzRWy43RMxIOJy4ydXpDAxMuXpv8FnrH9pY
pVsGvuP1aSiRaRz6n1nugdfkH5khf3leAqWiZCemFz+KlQyVY+Dj2BeeZtgSoUTr
enjNLRrbExWrLB8GWp4qfoilvDpRxOz9AiqNqwpTXCcMMKQPZgNIDNZrLoMFmKrb
Mjpbt1H98aHpgYWMxIUBnqCYyTHk4+3ePrpnjokCOs4SXmV38E20Jxcvhi/UyVI3
Qj5Z8JGt6oZQeNxop5iZSH+mfeHay616/aY3jXvnGYJgea5ZQQGQxFfxSifeZ5Yq
ZksUhJl9alRPpbV/VhqWqWRg4y19lNLL1WQxTJM8KakWo3VEcgwB7kT5EVMCt4ph
4iWDlvE/YC4puvqy8iUwCvD8hphJBof2/GJ7iWyHiz5WGY06QtB57IubYv6xv9Z4
S6OiA9GPrRC2yRLxN5mdv2/iFEi3LKg5GvDQsmoxHWkz68rSlwAFJSgI+e8nH4FS
I/EjnmF60PyQVzVygW/Zgx9Y6xu/Y6TH2nhzy5j1HAUxEyAdHF0Jl3jiM/XPb58o
JyfEbakD8w/REhluwrvTrEpoIrDRzYUBNh1WNKY2R1HshTTJbkrcvrr8fGweQfMW
hxR7LYTdxucERDlS8bqoBJXZG9+UoBqeT85HqMcLNV2E913s76ofQeVYwwqbl91b
tjdAIzVVu4zDYLjTM1AkfjnyjqHovy0aLK2wgy7NAicaZWgEWR3VhafLQRuHD3ej
7YVNPbkMbpnHRQmONm3wosqzZFsj7Mo5SHTozcRnAC/UbQe0l03ZG24R2hP9dxXZ
rPpU/0zaSXw3t4Mfa6UzklJ4lmDecQFfIsFS0QQ6kRGh+nsAZVT89Q2IfYYTLbTL
bvibHNIrKkmwy+pMp9atULEsGmko3Rox5U95sGLjcsMvDNknoy9DiImRh83ude1Q
+YsqNs0vtP73CqD3zeO/zH41zVAHwvIhsi54+lVq8+Fi2hYERZuFfp79Fbs5hdJR
xXzT4MIoSTBYnm2JkehQIoHTzJtFndO/t32CKBvKomo37KOO0U6XGdSIO7zTLdU2
i33z+9aSSdxJt624T0zhjxnaEWoF3HgtcCyYO/UwN0WOKj66ljq77QYTDblQsP/1
UVEdbWr0mvZjTii85W1SppkhnPm9ILVF35Qwrzq5RkjR9xkUyy6PZTHNCVPytyKa
a3vJBulh4D/whAGvZX4DM6zvzjvyb0505MYqVCgm+XDIh1p6ewVaTPwz63dC4+Bu
nJrXOA74gQPqYtJuVW8BYvdPMgGvfdxrSDEuizw54ejTDS4343qoD8MiWdEdDjhv
ngkKWGtRbEIkFypp6EE7M9HUdB5Uan+6wnOdzLKoXVI96uCL/4Iy2eu1oKDjDH7Z
cKHtHlHcK4IjXrjldW65FPl392jopLAu96WBG58h3STr2pLTXrY/MZWDNHYtDPsg
kL6AqI+/W0EzrzXFq0QEdIBfw1iIEhAA6EWza93Ev0Ek39Nfqg2u0axOsFdLVGX9
q7EdJMmhst1UNFiklQC2GU3Bceavr4UiPiOV/CDf72uVO/PpENdPSppO0LGetWrA
6RvuP2szqgZldHJU9t9TjI1AbJ1vuwlq1VIW5Tl2rsZRjpEqGlht1/9iN2Lsm12X
3p8YoF6a9swOY72Le1ehNKQHm2bZdGzFgV1V6XQBxg1qzUJbSI2Em3gEfqyWakqj
dZTpu2yIvPDH/J/fP4r9Qw7cCJZWvtZcK66k+CyACbWp6KfX2QfP/jU37hXZ6kdd
vuFNw3SDfwiLtCTSHPEmjPBM9trOQkyczJptdjLiZHqymRh/44OBVYLSCLdO0jt1
znmqkd+fcLAMaFzT/wRmLmV+WDrg03shhpnPGlbbiLsW8mCCP+jGAQ5qPJujij/t
pgNWG2uIchXWySjshAyjtWvM6e3suA3IF9WQNPCK4euPf61ZWu178mb9ddaUXNb4
S2M9+ApCmYQH/qP/dLnfxTeyuer5c9kHeq5v5Oma4e8xVt5SLbRbyRBl0/UrVIH2
DYfEOv5ejYz1vQ4zT6ZRiCwCYh3jClgrkpHbgq9My6RHwWmYINQ5UW8HFhoyc4Js
ZiIBJsATgukxOs8VoNYxR+9OPgs7eZP3bonSAq6qxHCExH87hrI0KycSLL8QlgIu
owAXYFul9VeRt6MR2XjnTt8htjhDyDfDM46BmDHD9t/lLZv9KpOGx2B+YDs6V43g
U1RrsQVGYe19tgeyojMUHg7/ivXD2lvWh85yJTk4YwGc1c4nOtgC0pSg1XAA6CtT
fKhVZYKVjGT5dDYvH248HZaoIEKUVDSB9aIXFUt+1a5CwjPj8rg0LU9L/6iGRIYm
/TvtbrrtJlJ2R2HqMP9ydcc28O6SlR8Rp93m/5QiYv3icT2iwEBG+m22je9lz5rN
zQc01y0GdeOLQ+RIiTe4kTrPiTLIQuvL8l/d743sza9pswL2zhzvF5GOLw3r47y8
2J8CahNBeZfNc5cNQyGf9jmdVUKSqAGVaSyh31opun5yt1/yZOjX/gc7RtNazW1y
VKol0psFNjEDZBoDSP6gQ1HXVRFEco4rPY+4lTcoYvYIA26H4vsMiGyXsGXjif9i
x72oWJbP5LBUxs5Ax0lF+TS/rBNP1Vq+B2EbwrPuGNBxDGk6it7Hpxd52wFpn/Ub
ltGDCAJ5ztR5uVzHwSIsD8KX3NWeZjspQ3F3vaXp51+FYbbQQ7HQFnXQcgEg1+s3
8Xq7p5xyA3WI/QzMnIk4oMvK7Jdu1PUMfVkSimpQLYw2uJXIBGvIZOguCH3EbQ9x
xqN7qXoA31/Hl3TtXddy14jiCLm9vpLEnhGfO5awiIln2Vj0zZhotRocOpi2Cb3G
wUT6FO0WahKPVBPiBl8VlRSsnWPfq96V2Ne8lH6TLAht2wZYNgY4x/15+yfmNMJ6
y/1DFlyBByrvfT0kD7KA0zLaPqup57by5FlNM05RdusVpEPKfywp/Gli0fgLRxRQ
qrcjgwCCimEXYWCRLj4rH2rVKfb7laxxUk8gojMFqXQHH9L/w2dDu8EoNHPPiyv0
zNiI93oUMxszTGaBSoa3kSfDtuxbVI01OamVXMsXeOflxlgMLNlMp+BxAq82GiJk
o9EOD0jqdJgcICX31VmQREiRuymMEVQAu3etZt7RoVP7ZUkTT+DOcH5nh/D0kFb6
1h4nNYKlZb7Odq3huE+osghUwsvjsZSufpKMzvNQXYXQuIqn2KScoaJ+TKfDVQ3e
2BL2bkwqg1+K48MOzQths0qP9RIHIk5dLWPhegFiMt0fKROqQciZ4E0BZ/Xo9l92
W0KKoTjZCN2ZFWjOvDvRDtSFDf2EkOdDXmwqHRxS1DeBYzFy0/iATFBr16mRF/Vk
ZsiATX/J98SU5fNlcJXV0Rvl5a2oCglERmNPeAyGPjHyVQA72sZnVZJ3isogHewk
KRDivdy9+QQV51PXsac+GO9coek26fjfYK40QakRy3sGH1yXBwzTa5Kl2Mdzf2TT
pJRyuuH9Tq05lvfXtEg4bQj5mmFU/tca1RzjEdFeP/IKqm17O1fkowHlmSn+Eocp
hszE0C2q9g+hdC7+yu2LiDtmKQQDB/2lNRufNi0twc5ScSJedxOHjbr6Av0vNTPT
UnJoNKDMFfUDY+eUMmvPQgpRlsr+MbExvPE0UqkN3LHa0mmiNG9BKWiq9Hq+2b+d
EpLlg+vGafUEOlrn/cAuUmdv5yAcYCAL8kt5MP6GBE2H7A9jmU3r9RZM5NG5/dlQ
5FyBE5PUL7En3b97etLxhmLWzaiDnUgwjwG/PJCy8CHyFJxGuxPqCaz0pwK3zOrO
6I73ZWmnMZkAqTXVE6dPbQ==
`protect END_PROTECTED
