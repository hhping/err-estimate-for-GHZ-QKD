`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HG3J8xgTBFS5HTaDDct5tPpXexlvfBRmwvTVXv3/0Korz+ei5qDUbExioJ8kqw8F
zYcQQtHwDhDFyCa9rKZUQMBP0R0KwbsdYyv+1JPuYQTBs5gNiGUt9wwH6cH3IR9c
e99Ax7VZwaozPnF5zLzlcMKf5zIYhz+tUvwMrxEoT6jNQaNtSBoyo7OH174W7Hwl
RUZwvR9PJdjO31NlMF1ywf/OHCOc8UgS+ueIWlUvl/5ROKDXMhAxMGKK5jHFRxQG
ypdQEvIkTsbwdFagpbKQrzXcZqDUadOFhcKUYorpZArodZcHAiObHgwzuz8s1AmK
gIC/xTfKQ0XwnTYZ+o4iTbcNktqOFZXZYAxEOt39hJmm+39tyWSCC+htTb6hrvCo
qL+5nJSwJ0cqph4clj5G4b141F6KeUDEwFlTMgeLprswtYWooOR09lm8DJtUJ0Lx
bAhID5UZpKqGgwZFEXLooP5S8Ebj/NztBJ6TYHpaelxHgP5zLEQUmOeEt+RPulWQ
HMhGa2Nz7V5PuJbYIRElOqddI6+vuklZ+CLbVGkZhjOUYKAgzNxbD4TYVQd7G/PC
546UKKiqgQ/J1USVly0jRWu4bFChD+/fd+DkkE2CLaZgv/3FR0/XcUQ63KoU8H90
3tivtrsINQcnDg3E46veg3d4YI8p7Z8f66cw7UuKr+BHlZ5iVfs0tK62H7uWrjZW
+IgJrrIlXfsMjX2kvhWWeMsJBxy4acfiL27RcEwr/AvoTXCcHNt71sJ9QS/4gXC1
v7Vc4y9BzShDCE76MdI0W97mizPtGcfssp1/JgnJAhIzzfKKPPgGPjnVPxsemIb2
QndNzzNP4jMtgzU3XvfXJygxoCvz/UKx0mv0/LyXxH9crAzKX8+ZqbJld2/zkJXm
y8I3XHKNpSsjjtlQpt/OdGqQ+Ov6qDwMjSrAt0yF48Rso3dpjnGgkT9jmH3K04YP
Rk4gQ9h51xmDYFrKrPlDBZZIMp0lpjjTDiK3WnSz41SjAzPO/3z/ByK6I7sl52JQ
diiIfveBdRJtCH/iLryvO5fN7ByWQG+mRWikgaR9ORMrL/Bg3Kfpqn6hcVT3FjdI
DD5Gmnrc0PeFZav4luc8pu1ROdaYssB9n384w6+1fxkUZRnRVGTdhXsqc5X53XMx
/kp5/JW3SNXa3K8J7w3HxIAEA//vECfvDvnk/HrTd5QwFL8xfOBK+NOm+p/vfP0v
USuFDfxXEnrpicWzc4LszUzQ0m793DlCLYAurtppO7TtTfuqcRO7LK0Evc5xZyN5
UdsaxySMt+MNuGnT07Gy1CMah/sf2YWql6ms8QqfS8y9MZqYB5LS/4WvhiNwuxCX
GhEVYlrvfF7360Bgxo2EFnN+lGX6d2jRRTlzgykIFIVIni0dXk51+MIouyx84fl1
DCL4l2+aVWsenCQ3ZPIA0uHI/v1myIpboMJgE2ACOXr+Ftnyc6OQQPXH9udT4XAC
3aaF7QybhWR0uBu9hJoiopwlehQXHXRmqiFlEaYs54+54jIBpCkGkoa28tFXQ6hW
lGPLHNVCmcSZOx55s96A+bk3iNeZqW3cRnyu+9l/jzPp9haF8v9o7F3jrSiTbuo0
RJQbIHZamk8wqGpPq9xx/otL/53JHuGQekXoi0iZdBQnr3xLug/F6HqEZupy4rEQ
0EhQuZzuGBHwswiYwW3QOJTBYdoNw4Ag/x5frKvYrlaZNkGc93sxWopAwWYofrUE
GI5+uKAi1/vG9ZLGUvdMqVD/yVeoslWlhW/GLXyqBXu89OTF9ASUILr4bnkqSdaQ
lJLVxXCqR69ZyTIxZGlj7l7fBtB5zqDyfAThz4pHFq2gNijXYhJO0bIMr31QlGXj
7rbZ6muuy4UM7wQwaU84VY/iVDlYmCccvQUGz+p5wnnHIUPG9ZHWKDWuqbc5/3gj
AYlWmjD3ZIfX/Rwn+s8An1sXKRBeuOEoo9FuV+SAtg0juzc+QLb4J2y1VPATLP/x
pXNp6itxPxu2AKDzrf4wb7N3XlekMHINQ+2HrDByBez4PKCYysDWM/hUnb1Nz2DM
vVXHfNyhLe4ggNABH0p6LeVFcnNb2FuvhPnYc8ySDmmrDCWIhXyf1TbKMxDNwNs5
`protect END_PROTECTED
