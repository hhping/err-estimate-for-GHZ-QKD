`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xpkoez+p23UzrjCX4ox+E1E9Q48emO8N8U688Hgh61CW/PKZsDckXPRkHDjqnbXn
fKgXE4APmeQxWNd0bz424M+YRxeruNBiGC/QovnwuWQmCOyS9SNmxGYSanJttlyr
szpKEnQNpunDEB8hn4FlT9X/M+9KOhi0cQUESf7nEybwV3OJGf+G3YoizhqvMH6K
i2doz0ZHGc6nyZlWbsNfF9YTJbPZPCB3tY1zP/RX4kbMLedsmZLOvQk3gbFxMEly
EKk7t/TpM0EabLEiLdRuD3Fa+k70KIA/JpLte+t7ojiuiOTRX8oo6IPU/S7DArfl
1QbDHamtGFR4CRuEGUEJXaWiV3XkkmPkqlJLWRMwBR9ZLVZO7FaqoGkQ3rl826tW
nx/l+wi7Jyh9ON9xW2aMdj0saJKKqcmXLxd6ITsZhWhxE8P2LKkv4K0betBsEteV
ORwfOZ2xWnZ97+YrlVRcnuMAsYBlN1MG/UNlbq4HdAgBdVX/PIc9rvrvQmEuJS/I
XTny/J+I69M05kqUFN4G5hS6jX5cfsIFM13+3wjfFW+Q5EXKxPO7ZN9IsNWHpTrW
PJRe1S5RJz5sJg6TiYy4oaPrTGi0uJ8/UAp2FHmy0hYnE702j/6qs5F/3kHCcQ0G
h2Wn+BmL1/z9q9azjrYYiI/KwuHG4XDu8THLY1m7KzE=
`protect END_PROTECTED
