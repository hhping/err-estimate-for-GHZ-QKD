`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x8vj6rjpDzeo5wkBPerWRxl9Oj6o2womK9EcoOdwE2LYvFeIt9TudXuRBQWMugI3
dpjKTMawplcWEM9N3GJk2Fv3rCXmx1PaZtbuI91LTAuDKO/xdaz9pKGsK9Vz8qqi
yAPzxfJLBc5cdpHmlgE5cO6sClhjGhpIN/jtGEtFMkGCF7Y1rsPMNNSviY6wY4on
0PYajeEDjLTfJwVK9vQ+ospEXRaPNTn6p3A7zAPZbkeUyOHADWPl3aXdj7LmRLcl
/b5Uj/JqOXTRIMXTobr03eeWMjn1XivFiKUksvwm4V+dVbggCYTLNh1OTuFPMXmB
wnJKwgHodGhOwWHvuVlDTsSop/5KUzv+WiErHMkSBcZSdVa2X8Z0mbDSO+ScRJaz
gA9lyDRGtuN5FICz5Jpyu7K5q1jqd4qI/foriVVdUEQ4h4yoIDDmjRXPW8LNfmJv
ksWd9HV/Eke2KP/zQHuaUq6kyYBrmAU7xGKobS2n6c0P0z1c4s6IXwzOH1A5yjRu
4EDjDSd+uI1vTh2R96OeglBf+RU+VlCAyeOn0UMPyNf7PM7gd+53CeopeCZ7+8LR
mu2kSdAp9S0l5+LnIMw6N3cfvUylE2kNlR4TYloTlbxzj6ga0buMub2C2+UEx+w5
Vf2rRkdGH+HcgP0tBy4qUqVz/PmcRFYVh0yBnZ6KuNBRpMcCso960UmfgLLOZ00I
8s9B9s3RAdQGWOHzYEKyyJ0smWrrVFO/IbZuMlHWhFSm+vXS2UZaUwyL7PLVKia+
ysz/v0oGgxNcUhLd/GylN+4m7P3Ut1EQ2mMcdGwPKXgtD8Rwt9wx0k/wvB5GRroC
Mzt8KL7Oe5nP1CIECXkgFoIq66uaYmtNeTbdlsCsuUK29uiAU57/vOhNmBzJGNn7
gxDyx5k+JaCv18OnALUlfNLiyFiso76YDg424BjPRzVnMx68+l5rGXgqFWOXwu9J
jfDbnC/73wxsNoVdJ5cgFH6pgd959Rdcbwgue1I4Ga6gfT56moCFlQ0MOiJEJkfT
PCr+0J+nH9Iz1rm4dTQwybvoam06sCv5wfQWEPdJwPZ3HutdaoylSoI6cJXwKoRU
wFz4Y07l7T9imDRQL56YRhecrRM/OvPeoKFGYqEVxD4Xwk2CH1LTSYcKQJEusZX+
BrnSe5R8RlSBrr8xwWKMwW31jexnq0coSCoaNvHvWmMl1tUK+x0HwK7rSMvvIsyn
Dfexen86PP3G8S+EfYcCvP78UhrcrnfrGSQzRFxJflLt31gB5gURtNzZ9yNdp6Kc
x/E2iOIpvQJT8rKTsVy1hInUvvpalxJ3yGPzHZVBQ+H+B3tMPpWdHW3Nur7qdxn7
fbjJECVRBX/k3OiEvK1JKnAYbH+ZMnnFRPtvHiLzR8T6M7JlSRMvnSqXiPAM1R01
sphS/Wan52huVVHthPLZhqrNjWqWCTL8cpXZehqsSeN6FJp/1rM0UXncKS6nEgvq
SyZjxYW08H6NjtcJljqaDl+oAv0SMj/QWWlIgp2L3u6y0/cnUz9+sSuk6mnREBh3
EAQMgAFaOLXfF/jXv1GnDxqTaPGl9Rk26weK1nqUqKmLtCSfEUmjZa3DOG+A/9rs
faHxgispbFLzuuPhHzzSftipOHkrJcJwtK/X6YL2wI8bQfM/s9szbzWNpq2iDhkD
lQG8fdFqaYMR7E2YaHhqOC09F3kvGBebODF5d0/o8lm9eLnsVE0QMbCDt6efW47E
wnD/vlEBjP1p3cWSCg7cQewMf1mWkukVNGVh9vye8wV2lPt5BngfoFhIRs+fGMMG
4U+myj1Kp6s13YlNhmbxmOFlI+NSaY3V/fvI69O/iNqc4TheZWagWPqttqN/yXnv
yJuJvvW94It2tQlLI3dEDTaj/g1mCzVTxLqmwkHYJ7RbZdAAcS8D551def7nneVn
5Qrerrkh23qnf6GR+v872YulMH3YrkjWy+s0ciB8/g+e/6cLGFOnyoRwDVT88P9Z
6b6T9hg0865wQS432cpRUNolZBo9frD2epS4lF/K9RKVmcE+vfk4ZyvxzHKizte5
f1klHRD0lyaeo66PRLjUhty8NpPWJq1qHZs9pyftXF9ERvMtsVw5dTdoicBMxoRH
8rQEqmMHrupEqVdpRuGzWKO3K0X6AE+mb7nmQJ8uZqu78Bc8v6T/KSkF3tv0XNWs
SUBn02IhEpz5MKDInjzWkFBrFj91nUuoenQDipgRKscP6mjJ3O15CPzvl8PmUIaM
eAIHxXKUjYBPkZKj0XyaADGRiKQLD9WKRY/YTv5AROvnUeg/8eCzB1rHZPV5Mm68
Ohcg5qtjmuCtnR/bbJB6Su5xKy65desmUk6+uVIjDuNvKC0Dfv/jNpQI/EY/aFE1
bFBHJeYmSy4seyhYJD/WFBLVn8pPME40+GVeF8K+I/Tt3Cq0VKV6F+joH+HahzDU
/5Lz0GU0upH+SrU8uSTK5gSZO+ppKNfyz8OsuVeWTvkgRovuU9xIG/pKkxw2Fp+H
+6KmoKxkzrcaK2oBTd1jgBrmERxdzrTGq83z0QofQBbH69f5qRQxzYVRaKEt5IcB
qUy9uOwkDqOCnXFm2hbd9Z/n3tDnbdIZmX1Nuz7g+sS02CBVB/ko1FVdFIzM0B5y
9rZg3N2eWLlvFzp1WcWOQXsMLAVxHz89EGb9RhFipXiCJfL0YwOh6695KrejQ+Ju
8Po/FO6fw7VQ5/7BcDoOBVSpYIjqwgCZ7020p67py8I7CKGkbT+ykH2Nhpx1NXTc
IG4bK6VqwZZYkSms37SA+s7TAHdudEKQvGvW+zQmqP8k8+t++2zqxaXPx6NQmZiR
+FxhaZVrXhjcdyibxxZ6Jg0B4xrDiKTxd4faJ5QRp52ofYAPZ1p+DKai1/Q3Y8NT
NpfwoBq9HtLUPyFcDu0EsoUVasplyLnOau8mhVX6iJIfM5VbgT1S6BRqIImn9gv9
oRkLT3YRDQehhWdNRQGse++768iEi5++2nVgzknT4HWeYMCHGqOlhY+BRX7gCfzZ
CT4flM8Tuiw3dtMkBr4mKKHpymIpcFSwZxTrwfBUvRkvZUkzZQNLpDb7suxa1J/W
+U1Laqj1M218JxEWsKCn5AgJIMenKQkt3jqTuvcKi/C3DFMwMHXrExLfiuTp3Ie9
gbPB1DjGmEGRHUewLN8e8yybLkMSWk6BV+fWLomGWR5W6TXbSo54vJL4aJVqNvYP
CP5UDTtn5nbvIXF4iRbvn2QaUPgoQMlXGnled3/lAl3Ckt3U3V4rclM6QK4GYFZQ
CP4YMZGCpygL/A99QSesDZY3ucG0wQtNXYo4kp4M4NbzFdXBwcAawJRtUAl/MF37
NEmhqLSCuGGj6HJs7JRFyNxL+ogseDtE3HnKUcnqa81H6okQZ9QSuELkrlkfzXer
kOVRcYSkkIFV/kyKGDni7mNwJI00x5jqr6EHkeMYyJTgUygi73c1EdW4eUcc/4Di
aW2a292O5pKKkfB5kT1yUW8ynbr/n/ObDCSlLfcEdIBRHEftjWimt97dG53p/p75
FSyyV99OmSw2mMXmWyQhq0syvtnobGiEFX2/uEcEYuh3/iWxQybPStPuKOy1JsOJ
My9ncTZnmCtsnuTxj6x2WRTMV7Kg6NaouLvo+xhE0NpIJEhTSeOpsN9BZJ4ErshG
kVj3/ekwyNKGPqtFw2PGGo1MfG6p98b6qyT/NwWnJtF4W0tZHAxS6rzwPRNXqjGx
sne/PLUnFcDcpqT4jB5Yy0gQNOxXAHBU7yUQAAjNzIzdJtcV3u8nvpiGWwBXLRRh
0NOPDSjHryuSRgl/FOTyb2rOzhQoba/bF1uqWviKPq55bVO3AW9iGiHnfQQdaTHO
XTczrzg8t0+nehN9pIraehQZWl8f5auDLL1ZXayjR08B/0JMw1rWw2z6/ydFuXad
Tkk9k8GXPJVH5YL/htB5OnIo0HbEYbrKHgm4gDPeS9tVyaUH5I9bmo4HhuYuty8+
RyIuLyMzVJwy5tff5EALhCctdVuhTLu8z2xJdKamHzsNe4+2ljFZMtBdHFZjvWra
wZxDxOOB2q7sn3k9gAw2+ZcfcKVQAjgvAyixYhPz9xpGGQh59J0TdWNwZ/vcWVQ8
LfJRzi1fzl1rdJg7szmJ9hDrltHu9CRV8i5eHpD2ZHufe6tpQQC9OHqUhplgcUnN
P8Ea4OXiNh13A2pkqshH4EGgA6Ej2qLCuyIw5BNuvdox5gJLSemSh/zYjhsxlNqU
YIPWOZfBgxOhXo/BG4MS+G4+ibDnX5KomMIzo90SBPsQvNCMFMHAyolRFjzn8ffa
XMLxdiQVH3G4+eX4uL4YrkO1e2xmmtnZ2Clflb/kONB4Kit5vzHAvC7LpDtMEqM4
CNPft3NbVBjHUiUmgNtvTjbHJ5siNUXgHbJlK+nR7VtyxawQYFZMgfsiVuglzRMO
wNtqr3Gy9CQZs48Ww/8Lw9D+MGU/uG/Qvk7dbiP6VqvyAvV3G70BKcqocYPHScqV
JHAT/9um+54z/7YbvzRwmwynu0GSy3I/lFlC2S1ZSdhvwmeCAYOsSv1zyRXJ9blR
nWqhMD7bTd3hkELp5Kc+/C4fAahE8D0TCNlTUbOTKyywPFM3TchPkpgpCNy3WDFf
Fvt5Hw8JwVZJlwNOYbDwBtvMoeT5Zb51Zm4qf9O1D7qt7P4nEQ3nagJfEMbajvLa
WxmpcSTkYvy+SriovNi8EMk+2bn2VQPs0065/5HjOJyory26yTafzgBEsy1XHxX5
M+6degWHhVLRDOMmF1E7Vh330UTqXwnRwXafO+BVZ9TAkdWBmtdfXN5qfi6MLzaK
pzZWix5rWMD/yxkGvHVDoXs+r8jFYtz86VEw1PxDpJuL3qX24joeSpgm4s0LtSWK
dPE1YwbgCbmLuU0T/MA6KCt3uaSol6RoZEOiBKVRswyKtqChDgQCuetNFyHiM46j
/hrp0YrDHbM1YHxOyn/b2N8v0YJPt3glfM0ceKcELjra7A2BXwikIPRmeJZSG1yi
fCj4CRGut0VgEtfJwCvCPDwCu2ck4yxcrjaAomplOq4GDLJy/9rJWY8UT2IEVznF
MNYXhfEeeNITksSYiYvgiPH3ChpYHsrU1+Tbk3DoeHAilPKK6ZKbQGhiWJAx2rA5
xVhsyUsb3MiKrFCNUszfTJWH5lDlUCfTWwzxUtghMqepMZZjti3ZCM1pmISGKJ+k
f0GUqmoB2LcrdFelP4CvVTOjVSEMlGKmY95s75fIp3e51TF9LzaydsZciw1Xh3US
cwh3KEm1CalrKkOEL/9TW0SRnzkHYsoYEUHJKOtc27vYDCfGQ3R17IvXkhXce+rM
zNkBo+bl37MRNBLWno6el91YkObLuEjUfsL1Z05P4ILbeRDK+S0upzxE4QPKDPDP
7TO8J3rbMI36PBUunNWNN4ucYHJUVzO6MXqym9sbBTVvFPHb/aYqDWRlAHBu/goO
a1GwWN787xy8cg1J94w0/zQywG3OqcolQTxkIzXP6Nn0JIptlF0C2tzYc5/zT6Ur
Lg/ZNkSLoAcQIveOip0dlgRC277CWrUZSRh910lt+I6c5q29AuY7HW/AUyWMU4ww
VS7F33BzkvsfXFmv9OTkQ241Y5Fk91ppftOyqtxoPeAFNiLjUQPZNv/gIrFqkv2x
+8uADTy3agHieo6L6wdt8Wh3SAsgiUGCPMWLLyNuUTDq5kf+DBIJXQhDHkzjWDMt
O+7YEFbaBRZ14khjTDuKGUafKjdhcmRuJFVaxZNnz/OWDfgU/EcOw+jx+vVOiLqG
6ZY/lxf5WUkh67QCB+/aXS011H4rhyaYlxbsmsRTyRCraHLm8LGRwz4pD9FfJNjm
pp5mXeq6xIjQ8aXPRan5q2Y+sEFedjP/8huNTVsSu57A6QAPKSzJVH2of15BykHG
oWCiZz8aBiamLWBzFw/0qp/+Ip2EK+TFvjy+jYyaIvk2mmJnmYRlZPr000WeIwL2
FwIwmKsEH0lSYyQUwvJDxNnmmztk2CJPYZeyG624djv/pFpOy0Fag7hptrDV00dF
T5GQ5ckkscakiHN4mvnAJ3Bb2sk1TArjDPUiB6jNicS2FGGsmP75TU4+cR5jeVLI
HqYLyHY76erkjwIC7YBzNfAFWzaWRW+tvp3r4zH2JQ2ObQRZm1YSyiocQihetHaE
wlJQPNNDW1CcT3JFXCOi5qV6XWB2NNUxg6hk/UgS0SkGeGZaZq/CquZiEWLPWQHh
iQ9kgNGCj1++F7kLMVIh/svdsv1Nz3rwdcxe3UuIGIMgyMHhEm1JOfrOg0KCfVDa
CIb0zMzSRLQ0rNtnq729AqEdKTovpGJxnG/vMP9ElPCtOYfT25apzn/erC2JztiP
CqFOBNKugXPMAm0fSdpEYMgGAdYx/3eeiHsrBhNVqNh09ji8KL3i+w8AOSxqRV35
zTCjX38QAn7Z+ECC18BRCWDaQvqiN6+pxj1JeC0GNN0GU3XTVKB7GqRUnwQwBLSC
9b/5J5ZJn1w36TOBcOX13sDiNPmpF7bevAvaSd3CYS1fgcD0+LG7Hsoatra3KhfL
uWvZIsoMfRGxc1DWd9SFnNrtlB9x62SXd3mho5+KBJkVDroqXIbEkBQKzch+gc/3
73oC0fk5289Re7/Vj5A6+U3OM6lGdnirFmXfuH8XH12NoIqgffDk0Bd8e30W0US7
sIrJJobpTOlQg2n0/swgd+s7MRl98UxeOZafLYKQR+Ny1awAkYUztpxtESFIYc6r
sqgCMX4MSsyjyTs+DxipO9UOvJ/lKQTBQr0taq6ZF1wuyrnHSteOD1Ys+5zPJhuk
KSbGlqDNtcBQMKRnvdK4iV2196DhRJ5wpD1Ux8IBPYG95m4FlskLfg4PpF5RW0aD
ysMks5cYnwo0gDOBncGWWrcLW1Tip0ykYBGPVm4+az2/iQYu4U137aaUVna6NI5h
hOK+S8aMtYUfyDYTLptu45jstqDRdb5q/irEN1/jSMdPmfMcneEjvTbUUJUPfhF1
FelC1xeW4Vny2uFtcBP0e7J29lKbnG1RLf1uDeoksDS/KMWMUll04cj0t1Uood5v
ENhC1YimazlsAssfQ51cbnGjRdETGF91bKeJsvctiuv1NgUQo1fGWGdMU+iUWE3G
2Z2B1Y5RfH5S4ZS5xZYDQXhOreNXLJq0Vhs8CbHiAhSxJtrAp5WHZjVts0v+Rtun
YBJzYV63RKOwbILteKQMVvd+Xrtr1FvpC2+YxPqFsw8pYP95b9oklLSMg1XEeZEX
/TSaJ4aupa0IUiAUE66mhLSX6ql26ylBAx/Lpdt3Nirp8X7NjW5bAGsz8n/RX8/V
IP/FZIG8uWrXJhyBmhQo8Sn7D6etJZz7aXNRIkELB1QDcO5u3IRspDdCj6LPL5rL
KC57Yq2WVXJrbi7jkY9LzaQg47VPaTvksOxtNWS7HgzUZdnxqE+GCHx6hqv+S7ad
DOC8WFUDwAzwpFiOt0EBQMKZ5msA8DsUEJlnoEctyoqssn983ryYyfL+lVbsNDEd
fhGEDgrvM3JcYwgZ8RmscX9FUNR6ecPoh8jpLmybOBReTYI3ZvJdNhVvQe/6H94s
PdmZWXmU6CuxJ0XrqrW4/luWKxkVK5Lh2GXbn2fnCm0v/hNSmDblTZncA6rbKTgj
7d1OxxzGWAiWpUXXiVY7oLxIgr/PwxEU7Ys/StpvID8KVBLXee8ZwVXfu4aR0qiJ
Noth+zeFdbGnyTlVEjNazgP/038Y46lJ7aQzductuUm4gZ8GHfzLWL0gx1zMZOi+
LXAMCU74YBETqFcXSHP+aVnblrsuKYmcv/tJu6Z31gGgEfoC5dsMJhbJJ5GmNqWJ
6mN8KnmH6YHAQGZCDvZx9lM0PJpAjdNKYNuxDHMRqfOVChIyTGmRKDg0vEenFTAW
QB12zh+vLIsbk0zvS7nYlVL6ItH6ofMyhJjyflmPiM3dbJ6mU8N4kXcNWnkYpS3i
qs+n9ZC6gpyQ/Ki2Cfw/rRGuhR9lNyd1AKZZYMKdMtDA4LZK7Uf2lBq5IYCZZ/69
3Z+0XGcebiaUoVAgP08PInZbjk/5fTQmdnnJX44EC1CztCtNCRRe3nmbnlvZ84jZ
MGVaYQRkadt9BAh0dbxTVG8LYYRtS6uDWj5OkeLA50Ro1WLM+Y/DFH178yXnJk/W
PrTbFVH1KIEhqMqSYNk2RAWwINaxKRQ8Mtn13vurgUY4DPsUx1SSroQsuMgiM5JK
ebPSZpZIcmP8+5Ha4ua4hMTqg2w5CmQ4Ou+WXJF8O9Hvb44pR5X6n/ivo2+rjAXg
51aatu8rUrtaUopF7Lkc6L4BDH+TuVmN7+s992Op7fZsJfdzN6ybNtwZcqdkef6I
GEV0dssVK8AlPoCUzsp7HjvdDxH6MN4RHPMW9IHw8fpb8ClhOFkwKZ72FAY3Pop7
Jk6yknkIwaUhgYvA3CqNcisfRd/xkrPjjjGAXANcNNV+Aa1Iu//Fc+vh89duUY3+
s+hTYgBWYufFEcOLI26Y95ZJzf0K30j4yqPafO7P0XuadcluTTA8jeZ3hjIdA4ZQ
U9Vv+UjN8RnQDiarJ9R4x1L5C1QrGOLJ5bqHVR7aKMMmw2uU5tlVmJVI2kDDpY8d
mIObu8HSPxpMXnLriYUkRUf25lR1pMYh1W4ROzQ/if+jedJTa7I7HHblkRtKnzWe
DNOs8tlWYTc8m89y0+Z09F+qdPWsT43z2MBetRNMqYBFmK5Q80Shiws9Jc3qflaO
euPstEhYYvcxEPkGySbZuPmG068pyfuSoFJzC4KH6/2+yyElPt632zeNKMHACZjH
EGg2BkV4OjJ3eYk4sNJ1kmCrJcp2bXFJo74zyT1jvLP0ckxAixAwGvkJFuSu4mZs
fiXMWsLPtF2H5r0rUKnPpKedoonuwQzImRgmHQLON3KkpQ6EWo/xV+gZdEz+BsqJ
DQ4+mVeFmOv5Bad2EMCUGM/LS7pIr2nelBCTLR3u+HcXGzdb6JJ4V+2xy0LdDoUI
phZsAWxlfAwVR7UPQC8/+rYmbWL6iezYfZbSe4PVuxT1vm4Rc4K4OXm28BnYQA+p
8Lxr44w+zbuNrq/b1PNN0NVhn+RMR80wVX6tCDtnBUQGZf9+LPPcpF1xpouvxSkJ
4wrijxcyGnv8ETZXaYnHQDX9066jmze77iXg7A5w32s68FCSbHQopgREYIjD7kgK
N2wqhylcnOVnNJSIGuYy8tcJwBUlZVdxTgolV4fpfemRVRk8na68ypVsMiHkOX8h
+pZyisjUzWB8eNbG9AJoCvLvoiahsG1kC0Wveb9ZC/MlRhMG5G7+9Bycu15s05cw
Z2ejfH1pPhHLjQEnbKsHzaMagAXz1WvRtHp1iPSRGTwEDuGfmev1IqPojSp1zbi4
VgdVBh+0c6sFowcbbGNUPS52+f2KJJSCQ/M6lX3B+ZtF9VUfapJY+D+dd3XgRgAt
MczOMud+pC0GujB18JjivpXes5z2bqj3j9LaY7zVEQMvK+3s1dcTr9HarbPDkfLd
x5RblPKuJF2sKYG+HUmNvB5IDW/6MnsyaKGsN4yrAmLkeXE4YZX2zo9Dob6lQEnm
SD3Sk9kFWNSmFB6h1CigIhoHE1cecj2LqymaJzSIqVcswslKIr60cxNAIk6pRUsJ
a5iEfQ3yItBjiIEzFE4t2dHrYuMZb6YZtPDQ3waXoTe5suUhijJA1uCBKaGpZ2Mq
QdOjtU+iU34q4wpfKfU81/5l93HWPKuzlcP9Otrz8cZmrUjZdBJidcWeCaS7+HIi
YujMiluuZ6+ARkTAmKXQs/zhTqFsfiQuRhczruiPOMvsjD+lSfcpGItS2ZQmOz1S
FCECgkhmjX4v+ZoIJDx06fwsvxiPyfopw7a9FF4bK8+2syoX3x1ta2iPCsaRolW2
3gsRz0EN7LBB60ytVVhdulpRmwPrMLBZmNxp292VFBrP69U+o3gTgffv0j4Qamuw
d0Z1HUvhFmnk/Mk+WhC1EodpMmoA6EWQqF2wJL/y8pBhXC7+aAHJOy5bAosORKNl
C20O3ffXaRMPA7NzLonbSVZ4zXQ8t/AjiEBOMNxwZ8wvDCyIbkkTG3c6RsnFxuA+
/wSUpQBtzZaTVEtLJm8t1moPmtUPAY6ThOFmxjojUvThZOv1o+MMZtrKTnlU7qSr
4y2MnoLWdVTMvkL+pHLbsskn7EuqSA5eAJR+aqYiTfQf4lt+o25q07Dhr83K847e
wFMjO40QT5olW3gHKfInCQWZmDQjNB+zZ6JIXCR8BEG+Yin/NOXX/Jvv3Dyp8klk
lKnqQKiZIIqoH9LpNxc4QIvj4Tss3TdnGO/6pLlZdrceFOEeF+spapclD1kmXQOl
E5QT4BRtDWpwTJfaluFIDEd+cI92cV4SoJEpdTj1DnrlVESUiooPn7QcYPtHk03q
VbN2EuSdibI6y7YCJX56KrHhcUjpR34riGDHzLbU0VipczGTxuswVTQlst4b5EUs
BPgBC0rVKiohVMQoPk6CfyN/4dOTLy3yBc+riN8T2KRUbl35Cw2dPIIKJTzVMWi6
WsuzvI7hxGrr2Z+HHEv74apK6JOV7q7+z5I3GXRNH4HYfRe4r1alXap9oWxawOxZ
nnGNVN+T3vvhN8zvcavZ9EtpEhVzS2RbLO/wuqSofgPpzmliG7/YFs9eJQNHWlg8
HGWnZ8hCck+TgprBDg86fPSLPhYPwAGRY5goO7DDPaVagFk+DyKPrejTQyeU36uz
rujL6mzVxDVLWoX1MzK+4JZuNgIHdWmxWwBhivSorCYuiIEOK1oTqE2TidSUEYtc
KdW1PrYX5QSJgCSqDRubBusikCCb+2/ppDk2xa1r+jtMWMGuuYskg4wRgrhZtdZX
+KufhVdFVabwQHhAGU2zwPBxPxPh8WmOBl8LnqUiNA9vJSjxdXdlfxzT+DjuuG/c
P8UpjbaA/PTvDaMIerg3Stk7ObEt1hFpM2OhtoWNAhjxEDY8KJBdgzItDP7yMy56
yobxyOx7BW2r4TyZEsT6QyZkpLvjTzwgEVojmQ7bZu0AFAA/wS7+d85c3//seqYK
nDCXIJSuiLC5uS6Ietvp3tHwbe9blnj8TROOOVi3bz0D2v6afTgzRE8/Tt8Bx0WQ
xeBtWB7uXBanRjnec5ZwaOxq/nBcmRl0FWR4qWJkr0y9ekG06f59Zrf4ERH8V9/a
tAbSctRx+9pXYUm1QpnMLP2Ozmk4+PLgOz4etn/AZRqhEUSTDuSXB/bQAkqPnbNE
JDfDvR/wBcC8o5ou8zmmKFPe8LOf0KJlkX7j9ETwIW3iTzQ24wxRgtOLNqvBhSgo
G1SYKs9zniqEdN8PFQzinGxCa7Xv8Id54H6E+AioJBiEz8LJmCKrwPur82krR/pC
T7AUrE5b47ch3WX+aCS/HNewX7snu2JydmXHrS7D7JKCIP2TtMTBmjJoPaU+z29K
QVsanGTPLZfGcAJ1oq0ZGpkofO/YCyBhdU1I3tvGlGXneofPkgv6LtlW36HQ9O6g
M5UhMdyEjKYJuSWqRVCv7F072hJlBSW9L69q1jRyLVRFIAsWr+lzsJlvGigYfrRW
FsYFbluDYQ+hDqo6hrz72R1WO1mpWsmLfmWkRl3IpDVlcz0an3mjxFdRSZ25mWhk
jzCPnf4SML2C0Qlwd6iirBexrbInc/cW45GSdlRBAMcdRIu2z+Qnv+g4uUmRcTem
2erXqjFhTYG3BxjO8LFQc6Er0S3WLTkxiU5dQvYNymJoCJcYS2wiqGORbGnDVPzv
r6CDn1fSbuzJz4HkWvRQa5absJrpiLzg9UfFOFCLWQ7R0SylRpzJiMe2bSTBCHQq
Yj+aXpPjMkw3bjo/9/rV5RefodARKydJpEplwwNsm/2RtPpWsz5shnoE2qb/L+t0
uVHOkZaphZxkOESk46FYF9f3HtNjQN5uC2i2H+6dPIwIddt4k3r3qx6LxFdCm8jy
Cp78QP1MXzaLyEYu3xtNUnVXbkzmHTPLRufczM5AP61FkWFFnqN9jz6RVyFsd46w
rBJNwyNDycHBQ5KuaMscSiHdFirPhlvtEjIranEj9p7zmAC5pbtzj9dm2S7Rbr9B
Qm4/HSfLky0ZUSLRjUu4ty8oL+fJmBxSgf9ijawJ1sv+uTefshqGixA6p5sV+JT5
TpFGidZDvkvmvtDMy1BeVQZv8cDZY94P8xVjEJKKxYqKjd3qpm1ux07dxTB86qe/
HHAd7RGVDXXLRdVNyjfx4qLtmNxcP7omFNcU6CEqYPU8im579y+2ediwYKk8YGWQ
Z4Kk4Z8vHebCHMgxbLfUL0/sDWrFMc/J5t2kp3s315rlnkXoWkqPeTEQp0xhFD3+
5Fwp0yKGmzWPRnM1kEIJRmbDp9NdviztRbjI7/IvFoAL7tyDzQzq3k3prQIB8uaK
HOAf+Hek4v5HvIxJJIuXc2MFBu0syvUlCqQi5J/oBvC1dQawR+eZHumgmyvxB507
xFd3z7KJvuYd+Jy1vymZlfQ2X8Q7vr1LlO9SGtffKXHOZURuz1mW2CRyTLUeTHdL
SsxX22NZ55UtQjEWMHS7PXBMwAFiAycPFRiu7MB1Vw76fOpCbS6mCua7C302SFXp
8LjFJBc19R8qQJ0k0JqoVbEBUgwrsVaoy53LySihN38N8vZtdxdym545lGJD8rOE
PTmiglxZdeIuSoORKXKwaA4wTD66+UG7FR0/vyvl/6o4WJ44UX5kmqdGV3xupfdK
PbZWqp7z1E359xzJAAKdK9HX5R5ON57/X8ZfXXBb6TxINjFmAC/2fiQLlrVojt5y
8550PzT7rBRKwFn7JmU7Y03Dp9Cnxadz85qJ8xMuknM+42EsTEFsCx+1JIScodKO
9M2B8ffn6ggwJzWA4ETiFKppvz0yDRm8V6ADQpS/628H7BjqqguIp1l3oVTfDmyd
YT2RgujCxnF1oOZJ2Or/orCbG7y929NTegs1slMuF5Fss2WV4yW+4wx8zb5QCYvs
JL69D939N2ibrDojBdnkTlX9NWtCfk1AB6phrxjrmlwJZlSBzKJ/rQduXKhlf4V6
PsWPxR0ZLGbp/31WiFe482N40bpJj38LVhk0VPlnW9m+COEDWBF5xOI7O5UcIUD5
ADuHWpk2EtEr6zjhiA+RUABKe9gHxfQUMsqs2zwdPpnJY9EcVtyWT5ZX/ivZkNWn
i5v2hz7ArE2Ti6R9s0T1uW3juZix0yQqzzGg7Ie5Xd80UcVyI3qm1YlfezSw8Hu5
3PhucM97QqrrK2VjEJQgY3i8EF4L/92K/7MfnK5/2l/xY9occPKdAC38U172alHW
kossi3gAwdJwyoJfxLewpPnNa03A7amQDMeP8QnnGEehstqgpJbsWv0KrUNlhnDs
KwXmrBzC8AX0uaPsCqN+0oGtg57/qXL8cM1wuIFUfHOVoXux+4zsZDU58uV83gL+
U/EEE88SlVwGv4LBNMEdLK0hbWxY/AFo8ZO6NIp23D3ZWSXuBUov2qbRHwLlIVgF
3z2FPFgrzXJYVsG4oX+fRgeVtMhaeZaS9YfmaV03ho9+BnX5AlyoWpSW2McfoKiB
CAFaj2AJdKbneXgvCIR0/Ej1DhuccyfTSU3T/+lLMc0ZO8rCicoCvisbvwdFRJBT
X8FyIosNJB4FcPT5Of/KPWPS3pzTdb7gQhupb/94MoQpx6kqFXqZOw/ajuFSO3Xi
DNameRKbAx6GFiwm3wBdUh/Hjg/TQuHHwOu8kqSgV2yiVaAp1ibq5usIq4nZqlQA
kHcqzSu5FGk9ePuiOz6EqWk7UuP0gxewBuA13Bu3hq957t0lnN3//bc/0L+Vlkfw
/E9ClHRofPsCx8Jz/vT31AMkLJaFOCb3scu8xhN+IcWsYJSoerF4Y9y4v3tnddh5
Nhe/BSLgDEeGkr6NV6oRtPzdPMHQbWYfq0B4VLx9hX1Jj6wb1bj3tSYr86foJTwu
xccqRt1HNH0oEQMgviNbWKAmG73wKSogNvYbuqCI+qlv/74uSeK8JVBqcaUdbeNP
mAa5Qoo7p+LfL/Se25SgcuyLhrmQPDtsf6KfgpB+LIVxITR8DZGS0KvHlI3x4fam
2oxJEt2isStx0OBKGEkb2OCmfMgbDdgqVzYMg9k6c3tDHJC5xb02vl8CLsVvDW+l
l2VCVNUeMO/nf3C41URE/+a5Og5GNK/T8pZQ8zrh4SjGpv4W4frHdgnuKd6GRQyt
z9ycK6kFmgouycCrzeGqRhZGEjOyus8Y0DuKG7Dp0TZBtuTje2cONB+OBgnJiyAG
KrtnmefYVeyf/avvDgV7MRe4Ze0ENNUj4RpZANz0nj00jQGtsBztbchsPUHQFaBH
S01fn82nZkDASP8ZXHmbhmpl3E7AU4ucqLqQbiaJiBF5J/BcYbsm1RH56/HLzZr2
DvTnrBh+7g68hZzBd3gFEvhUgruAYSF1F5rgIgbXLQS2wQCJrhmprJaKZTOr6pTR
PNjZRqykrBaz97U3IEPWbR54lmzq+FSXK3jnARLyz8Xc3xg3JLKR+CjgtY99X/vl
mbX8cnmiLE8oc1iRYUiwdWZIq0pQcMzmlJv2vLfRdfQuamaIuNyeTJql43+bPnQt
FhKJXNI92ryKD08LOXQ8Rh835BGa5JpcBzSsbEVg4Ui3+FKSDM1iUBFqauW0sja1
/odt4fBGXAu2mTEGCyIgnW2ijArbJ7PxWbvFeU7NEl3lJkZMefFGw8482TQl1wAH
mvHmLuOThBbDPrcA4UgQB8ZHEXV/ZXTil2ZLuAFhLSrh74fCXP3h+e6EB4J/hBBy
zCSCe9kJen5votqIu0LOjsCIkrJSxoXAWaLGzLYDD8y9rVXLOJ5TAoiyn7Ik4fRw
8vXixwH4KIlv9XCbi2/WpKkqzmsLStkcqujlTE0M/5z137JRHR9O1xWk0OdGNZat
n3TXUkO+xQH6d6UcGRUjBsnWm1rVGrjato1Ygw/KbLsNh0QRwlgM8Tyaz/DcGRq9
AdAoQI29YMGUdLGY1W3JQWHrLLwc3BHgevZaQ9DTdMDwJlYOYfJk2HC/Gz/U1st6
OyiimmkOt4QN3Ru52Xk3jK0Z/H1A6z+ivX2I58KwLphWzij3MBhxhOVwHCMq4epW
PM4k8bmNvi6H4PJ1DyTBPN/auAQFsXzrfK/Zz5ZZMQrRqVv44Xwc1RZsy0ndM+tv
0gS3d1kCSePQMIQoKeWVGqWERv+urpD67zg70cfp3RjdW9IfPrbajw/ZkwD52+ql
Md4wZ2W+t+zxTQrsombbx9ddg3F7r2Re6zLAnkb8xMcZDA2/26Qk+5eu5tS9yXe1
yvAmtgL2UBmGfLvZvK4VpNp6EzXSRo+1/vdwYcWzIlsSnP4YTbPGLd3sq8FC/2qd
kHneQEA42wH4tjFZihe8U0vL1rJdNKq52eJkkvyn66eozwL5MGGGJFrTDwFykEEA
yA+xI2YVZ6lzY4ioOXpXi2bRuMAiiDaE3CTOnpVHhTZhTN8mPCkiEsA+W8wEVnz+
PZwQ2Li0BLgFjBsvjeEY3vCWIR2tWofUB33TQEHwlvFR1b1r+COqJh8lFUSpvq85
JL4O4YfBnQKSAmnBcdM7UcA32nUjZkEk7atcbjF3RCHwueStT/jUvHdLTux9Z2qt
BSMBCyh+twIYWzoaPUf3uxm4Mr6Mn9Ls43+U6sLT3Tx6mBxkh3Ot46ayU8vUD3Py
bXyexKpKlY9ZvfuxKnPJBzDzsJfYvw7T2PccTfxH3tSDAvCZqt/V9vInhWXEmzMW
3lXhvIHOQM6zKDbD2HXWqCp83c2HswI5SAmQa9Ukt/nLvWfdxVjFIvO52tBvSkzU
hhlViQdMi/vd0NlAnMGPvk8LuFWI4msXnKMnjtAnpNBegrEfJ1JfYUKwDktQEJjB
pNTO2/d2MTO9YBd4Ry6QYSc/VnpLF8k+Tc/p7DHltrtsJGhaA/MudulY+W7yNVPF
5OnfkeY4g3zMhdUijcyA8ogZNI8Mapf3JvkXNwckJTlNskSDW328NmRTsYQiNWMd
hZUF50hvFGureq80b7e26tThyK2z98NekXn1cYhruVoIpYJgFTmbs/nldEM2LemZ
DM1AIF8UOBxj5Xd8NY9xpRtP9ZLVJ/JmFewjg3Rwi5fssHbQUFDaPhiVKt7vWkhO
5UrR2aiRzywgR3hPAmF0vxqhSz4PaiE+b9GEtjWCOyvL2nouX0Ei1KtL1R2UZ7Mn
6UI3ssSKTC5v0HmP6Fklutz9X96BCKRToGUpXjElMuiy1Jdi1/Jdepy7r2zylSrw
Q23yPji94aiXHTRurY2REA1SthUU9rrupv9hOgWjwgJTd1sQpgb5Kt/MPSkcTuaO
T0cPjNmCoks2oSPBaYE8rpLRETA83o4wc0nY5pj6CUrrUo6yERQOIj6yH0w9xnLJ
cU01cFHfoP49cy7ReQ8auMi1Wj8Ry48ITb9Xt3tBpwrMgGR5pZQxscWHHPLdGTnF
/Osak5N8n6/N8ua/NjGsg7tvuiw9gQ7sPRaq+3Ms0VPh3NrOXNKW0+CoP2dwsaIt
8/us3h0wueoBljo9sv5CL87QCOSdDfluc9se2rqLCrEhrIv3/MmpZ7ykcstsvZKc
Bncyk5WED0ah/3ZlSzHBTZ0lFLpkjvUD9qfRtZa5Axu1+U+kKmk+yQiKgycPgKPB
Otr/rLN7IfXiWjDMjGDoyHK+uJXArjHs+bm3KJLPE7IGo0CgPkqyWP0wdcQruw6+
XWnUSm50a4+P8gsPQ3nlwhcDByQFFfjhddGHoyvz64gxOX7VonbiANGT60zTniF7
CmYu136tp6abtND58QFP2iKER9ANt2my3f/S9vlUmsh6qsGSx+O9mQ6ETGTR72ZR
li/+oEmSIHu2wKpMRIcirkjKrXh0Oyca2uWq+CiL4yO8Kt/IEobu5p2dw8/s2uNm
jCBWq4VxGj04AFk1Qbb/FC1298o9oBAUrvAf8So5NP9spTTCtGvXeB9JkXgFNDgy
hhZSe2gx24unGdsYn7AHlo2MeYHskULrcuRODcUKS5wL87ikMDC/a8bKMFcdy69H
ushLUz8TTz8O1Dr2/N9fUeEdIzuHxvcdsrI3d1yaxX2zewu7j/S1HAVT63wmp7Gp
OaPEtVqJy7LKLSNk5r6Hkqz2B0PVUCUmJvm7dn2/PdEvCW4jD2XlqVYVB6MowC0t
Tz+W7xUsxYWshAShdHZWBLRHex2M00nddXE8ap+nGj3SnSQNpzqVXSgglDf3R3//
cJ2ed0OUdb0oUjxqLn+SeHAAekjbq2S0Qlzs96UQ3AMBVvd0bePsvr1PTOaNwMXG
8HFx+WJlcU8ZaKmbWkr+GVGBxDPEuo2zsq41ovhnwZo/4+mNOl5oCZZpQ6HQ7SHb
0R2y7AGUAP/L+lAjMPdsGpUtiASkjalvbWTyal2GHD8kE724Gd3rBEKATEnbdoEA
zjQgGs6x6YSUFidPDdCCzHNlHJ1CO7t7rVkUNQVndEaEG8ornlZI3mhXd2o5QnaF
QmS2EEJFypvlQDoX3vEUOD2Bj9RjheiswyiehfBar8Ate157/tKJr6UUjK5SVfU6
lgoUm5ono9nH4SQMsxqpgQ+8TqnD76i11Im+TuE/sXBKk6vvIplG66N1kEWBLqLo
xVt3DfgBmLcwu25UV62V+rbPVfS7FHeFavebr/LCpI2VtQbQF+6I8dltns3BpdNW
S1O16qZfbSV1jXHYgGCPwlzUTxF2W80gXbVlpZ73/rWJi2Gc9P7U1zapwH9lmyxE
RfFmDP/eM1cO/8pAt/8dhipj3v4EiWrAv926RjeW2XSgCGMu3y6RS2jAQNmM79hV
sleGD2jhFC8vAvbvNYfoZACl8aLdvBDn0UqwCxKkOhg1K25B3bJJ4GXuxS5vx6Cn
l6BFAUFE06CPL/y2AevV6fo2XShTgtcEuK7rk6YmkioTmftDLTMclaf+IXlTuWVi
ZKK8fErSot7FOrmf7D3k2jNZY0MJmB7821pjpTQY6+jyVJ4KjigbgUEdLrwqMbn2
1nIpbJX8tUO1oo2kpUeMMbjdXpkPkJqR+1fPQ2dgU7cv+9VqpC2t0447S8KATrLs
uKrLaOcGZnli1U/dF703AcPrWYLXkC4r/KBuDosrTUfJaAEqK2J4ZLG1nHlyrS+i
pQDeiA3IBQQ3TAKYe/sFQUub7sKJIlmoWFtMNRUy/hZxBdINMDb/C9iXekzN5rpQ
vO5xmMjuTa+z0ija7RFL5ldvK+gHrUWqfujzc6k69rgWSF8BzVu87VATwtyAMYPh
eUpyS4ItwL15EzxxlxARdG1/i1Fpk/T+puUMEDOHcOLyR+r8UEzgrtk3lEgyl/fx
Qc41sZHmUk6YEhIybU7beXwDIs/DSES69SToUrM+hme/uOimYCC7eyPH2RWKapHs
zVCYhaa3vxjc6lm8lheFgsESx1d3QLl8V35UC5WWbc4KoVhkJxVJK1gQp79iBYzZ
mWjOSp/NpTBlIJfOeila+JoQZg11pfGFyHHONUDRR/Bl46GCUsoX7ahFFYYVS3K9
8e99H5807TofqzsAeE7mK0UbkHQmNvzxXYd/QJlfaRnsleE5qj5/2Gv7fQiKeRDS
61dgh6jnh0tgETH8Fz+MlqbfkVZSoFT2AE2yN8wUyErFhYG8HZr5p+GZBQ8cndDL
Voc5S/zSYHTrDWJABYkcoyuPgjNUIPHIvBbAsGLPbT4Tgfmz0ntrsYTdMHOklauV
qoCl+3NSiMxPfzeHjOjCPY+DXqD5/JLXu2Ct6srBeZDKCROkc7GL85kWoz25tno/
xK81iB5u/d6Vh1RMvTtErtEsJNakAMu3BOQplCQwV6K5tJ0Q5sx9A64IgnxYy7SC
ukqLdGH+Rtbhy4mht9vWJaXbHaTXgFtazevdg4x+kZPgOIcJHZsVCcFFbsoOY1KC
u/2RsMliLvbxqQZtCIp6FbQHJfZDrA3/A3rUNPJKb85UP0xQLJ+Flzw7khvM5Zmm
XxW/tPqO/gqKVu6LG8en2NMppJLHIE22//UUw1CgDnYm8Ef0cvP3+YhQalVfxF7H
jytp+/LkrvIuhOdLeb0OCLVHVOamFSM1vwGOfdRG6MjwEWZmhg7RNNRvYMGMAuO9
/DhwhkSbi/VD+NzQIPXN3z3/oC0LHQ/WxdoycPOm3iUSvBUOb3Dn5a9Yyswh9NFK
6jpZrLBll0VpfWrnQdVU7mOp34UxrQGTGaLPglPMx9liGCeC31NZJq+bfDMmSRlW
opUne52yXdKq04H/PGPTcHUx9E70ktSlWjMLnjKVdtdBtdQQllzHac1sHp0XKhZ7
AL0IZu6x/DJrZ7P5EhfczcCYwsXxHpQyMrx5GJLEkOqpThrhGHhOLkkycMGxLnre
hZjeIqe5tOiVT1GcYTVzrjWuJ/ISLSvSVk8MWARXKTBoTcV0SaPP3f9ip2HVsslm
9tzb6gUF4RtcOjT9GJydHip8mUUS1ZTV5L5VRKLw49oip4XRCtrFqVl5M46jAfWz
cOYyGXQGkkuCMj28IIV/ubsSQea4AkYTf6dDzZ8ouNbswpPmIk32KjHBR77Zrcgt
Hk3RcaTyhm0teb7JtZpeY7uTYZp7Sia+K+duifSspk+xQPgc5g0KKd9SZDTd5Gz6
dSvkjugXWNUy18ItmsuJE+j268KAjzU9ih5S2j2BEwv2PAK+toKYsFzQxqo9xgQF
klL3ATVKSdZi3TuajkMkLPn3XJxu9hZ8F5izvFIWIS6wb5jX6Klhzu2jjceiV0gS
sLwC7AERARjJ5CABt+uSCsu84Iw7Qe8SvIb9oazcWl7Ne7A1SU8lJCT4mY+RxeyB
vn9JB5MkEV/eHscO4kis8OnqZvir4tUH4LfVOXMeeUtB+mvle1PP+ZILNHdfXEIX
s+sp2JVXRayBUGxde+rR8ZdaQmVRTAmNeB0oIzkxr9/YvbPXRsfOSzDJEKsGXkuF
qEqxTvM10IUsOTgzl4AwBwNeav/SrbFpGsHcXnPgcRQXf/np9vTSYNzLxue5CGiw
ILcAwY3aIN9IALxoKMbEGBO5l9bGqrjo+JPwaY8b78kG8ij0iIS+je1LxA9/u3rE
kxSuFTqtKKqkOzEtRZxRs/FiC6s1x+dkcleBgtv0mhpOgKadEceyT92vO6OaYImR
HJuwqt3hSG9IJCf20I4n+uw4rLY/+LaKH6n65sDboG2EpJSYdgzTTm1+aOAcmeYJ
XIOniQTE8XOqjR6gK9tvAS/i+MJMF0gzMxfuTTKnQLr3CJEB2Aty9jeicHZOUTPw
/7vP8cN8pAu8ehR6LJCJ3CqCQBY1+1IC2088mTt72QWPzWZ4RMebzxBPNTypu/S+
NkxYkWL4ND/HKEsehzyDZgTzlAbvZQuarrSiXJwp2oCi8iXGYKPoOUhb/ddVGKFf
RACVJ++JDmV6eltsGkzr/ZA063rLI51bV3sONumW0QjLwBAv8PG5XobGWQPFHpX3
enVnMiykrXv2dmjTRrBbwKZ666gX05+FF92bH5SUddxzf3KInRoeXs/lT6Wsekve
m8etbPJdF/P/myiKf3rIQCHWyLUHz8VVynBSbzfjxeO/bsQovD10J6kfakdg+Ugh
k/yI1lILjqb8PZpkoT773jGvbGsxJ2Jw6OTSfdyTlSW+StrWDL9xednbtA8eFMDa
S+HT/9tYLY64gogXmn9rwWpwe4TNWm2SjciI181wA7uFmQvp8X7qGJd4ScKuF+GG
/P3izW1N0TbAHPwJxKw/KAOp7S2xhcQsEpxasD8gUplJ1iHfzpW8R6pCWxt8lvk6
PIoUF/z5xyQ+qHaMpihJSbM5yA7eNqHWBhWmkqHxuHqGRWNbNqqN0kPrzgdAOyJ/
wjSPBi2eXyBd0zbn1ZXnxUQSlwB0e5dX3FtTfQrQTbj2DSLWHmptc/7Jk7qTrMSy
FHkz7gLJwEX8d0adnofdxBcDaji7msBSEzn4/hrhPb3zAcD+/+TIJ5x097WpgLCv
D8fq+G7hw7g+rkCRnC/DghJK3mPCGnbuHGiViQcvJykKTuwpggEqahn8Yrpt/CH1
BQofK+n4wEjBWeK3drdpoU4umius0TGSdLp7PHpJvjp6Pob75RSPCQMxvzjixJdp
PbdkRdrCJoRvkbtwr20MRzjXw48o00uH/xKVVyO7zLgmYkNqL2v5in7beZ7i5mk0
+2YBDh+Ne/s+8HBl+dJ2d1DO7DN+J5wdIhJsxaZHQ1mXGeEB1oodGvxBw6SeJyRG
2AExQL9Lm42iozY0DN57Owkuq5aAztnaZYrcGs121WwWQhHEO5t6EMZ14Lv6Dvrb
u7RaVn3YzmcVXUBxxbLiYrXZ0T0ag90fa+vfc2gOhYhipZr2aNqqjcrD6atQPaUW
K5sqB/agOw07dJr6anpdlrWrm+E+q9/8e85LZN3u91ay8mQ20nVfEqVfVptzaOul
SLf8dGKsd5RJiCxUrUKostCM1VJ6hX2TM+H6us4beTilcioMkfx4+ok8VLJPUdk5
X6KzplIsfWTiXAgh/ypy+hOWfEhky9Q2KWQJKUKNed/DsocU67yRSSqoX1TJ74dd
0Q0ZQEnVp/A+Yf3H5m9EBBs64Fq4MD2hlb3B5aKe6pOSVhXtCTMQ/SGWRTMbDWDH
jbDTaJhQifw0LlncRpSZCyM5SqwlqnsidzQsc3E0y8eCo4rAEEZpCb+sDUHKnnu8
CLCqFQnwaCLy70wKGW5cS0FEz5S1+eYn7+m405jRsvs3QAT4k/NSnh1rDmAWGwmN
SjkZ9ROzN0mRDTRQdI9m3oipoDLWmodPaZIFFNp+yccrH4qr81Hrkj/RfAsTjNK7
2hIrIFTskwim0nP0vuazogqaaLGOXplasWm+ZuBkO2z6+uzJ9/wZiVaNVURA4HLW
7SR3P4uK9b+L6qvCB/aspEubf1KXPNuW3kZ9d1l+RoDOxNAfG6fRULC5dDXH2DUU
ZigzViSBxUaakjzJ8qGPP6sEsDb08Tjwp2yaV8tcEotFf4MtWI95KoKiYK6uxPla
lv9iXnNHYMlhGsfER3fkCXkIzV8dZOg8GxUXsoSteiHJD+TDIm7YHYEenTUmZelf
Zm8NLr77ImztzhSsw6a7Xxl4FuwqYBd38+89Q1vg/VpZm8RtKhp/xP0rzcedR295
f2wfGn7BuQEHi+zf/cj+bDSuSbCeZGaSpXDiKpUdEG8ooMWErXPXZO714qiOz6NA
HbIfVQMsHj1XyEcIg28AyHNfu1Q3UaB9t3sB6vBrdh8B9TNWRbPD3yE6IjVd8QaP
mtttRi4yuZRF3JzPaDC7YZ3UTA2YcnQRgLsZROm75t4PWMAG6UopCS7VPES+NjbD
ifJuFxnjxs+eXOY+8mEU+XYyfEQ4comkYm+HBuT4wEpLmMnLl0XO0Cq/bxODMWEB
mhaCYn8o1DPfZnX5IUAzjN9e3CDHmlh406BykxhQnb38AWa5cmBUvmjQs1H8Pz0E
soJIlzzIprcMpgX5jbMt7oDA1DmjE7UDuxVd/V9QUjQyfCjiQU/S7Oak14agF80t
ZlS2crxkZfIjcMdYEmr/NK9cekc35At5sX5RhUcT45sUBzQbQQF4GcRkUw1bFDyA
qGs8QEPSFBWzhVcjQqla/2ud4GnnAsuu2B10fbEwqH58faDwJXe4Bj9umGWROQvT
vfhKXBqMrZ5DqYRfotwzlS/Z74n8Cl05bmS2tzSGGmjbNHE7JTF0TF3IYglHykyT
BU38JHE/v8Vxr/pw66ZeXnUhbXZf6EuR3j5m0YPDdgNP5KLmxrpIhd04IIYw08Nr
LQkTb+48zGCgNSsdSua1pzA96JLwi5c3FcuyTNEbwgRqciFwngrTxAuu8WMrKDop
qwLbShTCbadiotcXB0CRdoPzqimI1fYScGOnQWncz/A4k5EUKOKO1HXcvorHzuYi
ert/tbGzZNfEuZ9ZWfDXB0NIqtz5XaU9eETPDo8u+/d/NAuvQsP3FDrk2LeN+p9L
NlI0SqpOwu/iq+CCbx3jdJDEUYFHHfbkC0wDVLVsbe80lryl/PxItwKV1At40SNc
jQ1lgEWeDt7StN72M+qa+jq1+Pu4bZTB3aCK8kJHuFIELcM2FMpAYhTGmf/T1IB3
gSySHCOfRtFH4TodxmwlPknb/kwpt9CXEArHcXlMdVCA4zDQFmvseoO2Aa/n4S/3
2wDCei5Y1y7eP3Fmo6upxX/kzcSVzEO7TlUTigS6WPkE2VrIUHYVFSFqm0UoxTsP
A1TDwHOYIexome0MpRmampVyrLK2/jcOpY0C6gf9oH4hps1unE+QadIDSRNg4NGk
bal9K2ntp1qjCh3dpjfZJcxLNsxRf231O1Dc6/4435RJ1JW4HuvlMAip9x/3lFH8
8Gb/VLhz2ATVrzucw9twc9olf0aB862/NkILi4ULmz3YBBvA/vfdYrsQZeu09dMk
egw7VXR0REtvHUSBBHyjwDQMABZMBrWmZbMxJY9jHoZN79vsjuNw5uT63IzeN0Vy
PU4f2JdXFeA+myCIc4spQHj6xXuAyySlDAow8gMQo8qgPaSd2P6ZfOEWe78czal7
hUaVftYqqgpIwGXYxL85at3VzwEUeftuA4OrBDLgel+nLpJGSnDTDTqR8UOkL3fV
6uTVRe0La90GV4YXAqnJ5B3FQsTwuPsVusJArhu1gHq7S2jBujhy3f6UEF6RyUnO
GgRS9tsCBYWIrTRoOmxS+D+K1qCkavq70R8K48qZ/hf4a+flsxFLL8od5aN5CQLb
VrrDCd5mK2gvGzUWZiLiYxsalkdf294dvCnN3pHdV2kdD9Grh/LW8RzS2IlZn7Jp
LcD6B9Suq8spmvuQU2ypfkZJIj+FZCaS828EtXuogwldDl11yyWvLCg2FSBa2/lx
IFzoskkdLsSlTvl8hLggHlJuzuc3qPrbXReLoBg9401zv9E315mKm3rxG+HY7C0b
3j9lmz8YsU1laCo7QzvoV7sOoxSPVDy8o78Orps0FnN5OPpRI3TiqZjwdBzdrBPA
QsEtB8AaQ55fCfnAAw+kT0dDVlJPTOsUpXiQ2d37/XyRDfZs3EDH4+mTTE0fWpbp
Xe87ivo4VDHcuexg5u74x6N0waoWdrrMEwXVXVYb78kBwF7P0t1r4IOsaszq58VL
Xnx7y6kKw6Qkv4JbRtZ599/vwaiUovu4lPBCTgsas30hQxZ4OT6y4322/L+eyoDp
hnDN0Yjmm9lf/NbxmiihkUTh4y28mFc0kvXkro5p0Q0jXOB3VSlQ8gtSl511PIk+
g7PF+ZGw8kpSP+PeFoiLkoTl64DdoPNgpHjC0rBF5fguqJBXo2DiACwrudcrWuas
knLFYRZcQfpIu1EIQShOkfz3gKXtVYH5R/fjHwzj5biRohSH5foJjDUZQgY+NIGE
mSGvggxvulcOwRyMYDz8zIZ9igLzsi4+ti8fwU4PEI+EqxRvK/n1dq4FUumBpMMP
4yCTrmo9XVM1jzKRxd2IX3Rx9506HfqerWliP1lx72U0/DW5106zBh07pOoxbsX6
zM3d8b0RLfmymLhocuVl3tHycZjXGmkNjNx/FUjG/UEXcp5Ssj8fRM6Ws62dAHpN
oe2bKFz8h3DM/TckKL5Ak+4G4TuhYrdb5nEZZRE/mf8E7fzwvYMiibh+6ThUtaye
vyxpI448xZlw8w+lKmf9fL7ImvgSNmWArAoDhZYCFSp9CYiuCq2XhsOpgP06Qf3/
UndXlZ5GDMd6Bfg8Sd52b7iWxx+Xl9KQlDZrZe13h+lWYSnv6QHWbrdhCIebSG08
hI7jtKorRH/EoLtonXIAmKz86pmWqKJiRRhMhphkST78jBGeybOJmB/ZtmyqoBmb
voBqGaNAjUmIdx7VMu9zWDtQhMmeGfI6R1AQYXHcTqo59WeOLZJPSfm73MSifGzR
wZ6jE0XF5uaMWuR+/u6uhIg7QWE9ALa83TDXh+1f7J/1dvmKO3DZe8nUHKlVYEOu
xwrZiWs6nq+e4jyN6l32wWd+y2iYfjvnLJw428oyBonacDwkJUlgsiUluWr2rrz8
Z6as52hlK7wO4tcE/7qSJ1iLPbbXGV0L77yM0VbzAq4avbSjHzrfMtFGavHsTPif
6VKq8Fw0+iQdUijKwWnxRnmzf+qgrH+A/dkqWhzK9ylX+Jt8ZppXmZomoJ6LG/Qy
LFDyGeYOgRM3Wc0Dt1dFa7k/puEFRNtIVKY2FxocS40NTa3a4IMpBvmMlsjH6qXE
Zdpsua4vP/48/KdiRM8EzLi6g2mnznC/J/cUiIszOlxBexjdKl+7CKTT8p6PBEUV
WwbqLC/lox/VQuPVOzRYBOHGN6mCWpU6EGn6C6hsUlQQGebMe1k9hs2HyagEBooq
uJS8ol8sFoB69bGSdpG+UcD8FAXhh84NqSuW754kcG2suL0N4gDvKgBBh2kttFJm
qmqZnhFgdiSLRmBxA4yBBKxa5+xBIb3fTVgroM613tOIMcm6GUJKjl6KZ80x4Szi
VhfT1ctYo0ojpBOB+lUHvnQnvn99k9z1mftUZZBsXpH9iPw7aMWZQGUigCuO+OsG
ujYrBBhB0dgO/abqy0eWRUrUYtODktiQ5ucy1TKDmLNMb2W4h0dj7a20/2jkuzji
IkByGPv/X4n3wk+2WpZxWmMP8LQXBsYGfzshXGVtkDXEVOwnxAvZuewQXnTuZaWo
VxEH+tRohXUNyalByQyNINYGdm1qDYbMPsl+GiEeZXZzqkZtAuo14n7CKxP9+4SY
NL7HRr+dlT06EWRYrTRKi2pUr75EPGJqXyuaDN1FvN7ntQhYQmScZv0PPOYLMgoQ
8orW07mojWo8gAAEJFaQl75oblzy9vFWs1vhlmFV+O3hDJH9j3XIt0oZLUI3029T
zinkfodd5fXFtYFqVxVtkqNiZ9N5tKIvT2IcLBJ1VR4lF9OAGpyEXrE047Yj7CCq
7NfKSzWpE2bhOtW1wr8NQmJvZ2W5aek7ejh6o6qOylOL9TOO0iSM96BYDpbMGNJ9
E16Z99gRQ3Gh8BTD6urV4NJvAXdBzUFJOnROBLhk5xFzpALhXHsm9Q0oYxa/8xZ+
Q4JHh2s8cA9xVfVtEVQLjalbLdVqf9HZhAdI3QOZU4wqlmB5tICTdrvmV25TXhrj
Z0Rb+zP+7rfDP16Q+VqBCzPqK6/t1kHz6shUR7NoHFdFCpF5OLldywEICLfC2Pgm
imXeo7ZPCBvmgSMhRJqBdtE8j1Eo9pbcMrawvvl/kwOiCZDBYheYT6YHldObjGRl
0HNtxvElPnRMdCv/9P25CFqA/bO1tR64HBBJEgyp5/+9M+w11yY/ZvnWCzkOZf8D
CJn9QcLPf0U2yhjtn31zWyQ12ODzrgm8aZJYbTKZ+Xx4g1i7csP3q1Nl40Tb7me/
yiQ78BaWN0p0I3RfnWbgZ+oNFjBMIiSZBVsaA4/BY+FdkREhiNDQ0JNMTkRRktmm
3RQAdQsbPeTif1/7CbhPiPioC/C0lmUj7/+bmYnQ8CSvoVoZ6wWNQ3HMp5cQS6lp
uKtWSmbgGFDqv1roniPpa+MkF5QtB+BZQqD945HOQ6F42fcLEBl7eMRoO80TwalI
/O9Y+K26NqGIpBTeWo8CCgdaFxwWQATkmyACUKdQXfPeKQXeAr+JO75thnrI7ll+
8h5Y0XXwB12kn90yyRbGDYcY0pIBFr1F1Hg1l+LfB3WcLpO6JcHFQ8jJ+iwSc9ka
lzdNRTHd/6cESfLTEDpx6ZKVg48ZkzecnQcDVUyPbmUboarT+/irXwZtj61r2Lsr
cm7VcMp0pLnFOpLwlMIu4BCWTfXzQ+lInB3at39tml+fLU3hdx1sfjZkuURTr+hr
mCivyEvYCHyFyMSFEpoVHhffVAZrRzKE0eLEPGz49S1uVw3X56ff2lUpy2DZBA3r
K2p8pusEMc7/E8tDb6ibvte9k/3M1hbaPVFTwNjXF58OxysM9xDinx2/32OCVCZP
YPtbJyjukGvhz4Ke6g0c3Dcjeou/ZfHwW3S0ffX7lo+z8zVzXQdt2Ppd9d2Q5oUd
MIcxPFhaFcP0hHAjXLdEab31rmZ6HJaV+ZZd/unPPDE2Ibd2Dq6iLKmMCn7pvRFd
niFcATa/vlSOo3UDvA5vJm0Q2ttCfrJcduArUiH8KJ2XVIFaY6EKZllJ4X0jR0Zq
St+BZBEHKXPa7U7DaqStY7uj7Ow13yMzYtUYm20kjKeXDlWVpMEu0G7UZ4tfao8V
94wODj1cocMZNDf0QRmsdMOPAwzcXvz2Yc3a1iLMTz1E2VMUtRupcO/HXmcPJYox
e2iWcXluuCclmo6vM2Wxbg+WsR1d1l4O2qZgMGE/lijX0wKjKVphcDI3e7+kRQKl
BFe5A1RaPmQ8a+KhtZflfuPGcOWEWMX6cXpeY2P6tKd/z6jJn9mQ9F8125zaoy9Y
KHx7h2h5BZxz9KUQx5W/LNtGxnHqS3KT308VeaF8vz0dgTvWuuppbTqW24jHBg/D
zHounha0WwQxU4BoOqLiCdKH68glNdcqBc703SJMaNEUEX81yEmOgLin/pqxj3tc
Hc1EgkHfAVgwBl/rtsFBI7mK+QAqCKHFEMyRO7jmFjQzr7TkcvebnZ99LBUDjb0k
i1MwSp3l/1GP1lzKwV7zEng+qbWOGSVc8a2FTjn1tyIEfboy3oj5LbKlN64Vj/Ps
rkWpCDSjRAf6ogiP4JusLo5QhoxLkDmMAXAUn+StblGxCLLi0uuqkS09yeWOBjcb
VhmSR9WIDSYspxPpyzSnSajGoqgZ+NdNdeRTL74AN29Hd3InDzJm0yq7Gor9CTe+
7U7B9AQkbVcauivdf4FHfy5hnFEi3o78V71y1B0w9g9+UIr2mCEJ+edWXazLrPOW
Iq3DE1WFGRrK4AliJJiwFu/Rzfji0OyfZ5xW98Eo5kgZTMWYgFBF41TOXdlQ84bx
OooJ+gieVMaJNMmheozw+VRfmazYt4DduUwvqt9kD+Jeeq1s6yKr0XDzgmCfb5Uj
FtcmfDEdpRYuL8nXBMbX7d1/BfamVCzdt0XOJwPAhaUBn70UbKANOc6P46thugOP
KuBBP/s2TaLUX0vGPxiUlz2hWercmBjPvL8VlHZzA++BePFiCfbuD2TbOHP5j9sd
tkxyXe4ekiZyD5sC0ypGnHSCmPKbPUiB5MYtITwm01C4hmpEq2vrSkiTYTYlgMdp
HsPcrl+tvcWwwRUZxg6tMf9RTqD1UHcp47B9EzBYPOYv0XuzduwAJ9oOQS4BiuJa
IQL6JV/FDtBIKbFJPHGxKMauBt8/RHpL6y4e+2JeMpfe9ucmlbY7Qb3PBkKjwkqh
tJx08pCLTZDZnzWzodyVSjVDou4hWqbmi+IxmW7hw5rJFrB3FFBNudsVZzE3Eez8
BGzP/EdzykaWNFUo4TVQERmcJi3YI39sB8cnBqe0Ri2s9htG8auQK6Jj/uoeS+qX
c2PKOPNpI4snv+KaaYT7lAFsMUB4H78KxN3KK3IINeP9agD1HjhqxhlO7Kr+ysb/
R8+9/90wdZ132gW1C2ptjny/PJQm/exG9gcXgrGPmQUXiav/vL16bHPxetKE2DH2
rdu54uAw/PZuXKTuGeyYThYrhSAyTiHz5woTt/JDkX8n/ZlTd8cydxaPBbVEhyA+
Sel2Vc1ob5BNO3mgFhYtukJK24cRb3jWt8DVayysrVKaMq6ds5DDheZTj0OtDJwa
oRSQYFJqpE00n/Bl7c/Rd/ZOS6DOyy0Msz3Up7Hno1N9nblruyf1J1Bsdkk2Fyqu
rA8E2ts30PdNdFCFC6L/GRBoPI6269bh4NzsXxRqNStZAjkiHinQZNS66rf1c5Ab
+vdiSuRR3FR34CFr1n3eEsxuxAGine/0HOly5cWuEGeZ6zyz5gX15AKnq4Emxtnr
zh/p7pE2QORh7HT27CQJcXWKgYCkF3CqLsTwhr/WD79EiFA0U3nXO+TF2o2hdrW3
pcLo3Ca7I9TNciEdTlCZu/37D7lfBEPPMk9QpFkCOpxEf40moHLHSoN0WubMUDfR
dtZ2slsdhej4dXAb6FmTrV8O5wB/AFf9H9tSxz8F9x2yEJewlZs6Fi6YhBwXPedY
CFtY0mDl5hEncB4DuzuhaXoHANJDPNZoooOPldvI66WolS4JbDAnLdLCXapXaNY0
Eywtm4Fi1yiO+a5RB/T7dcYdaEDoW/xOUHqRPjVlTnh3+2QM6XQwfmnT7l92wgdO
tEgrC+IBlnppk4ZRK1Pj/H2aJy4WTgsvEp5HI6YRfyWC74XWKdhEb1ILGSvpKVQw
0D/z6iE6P+7tyt9u9NHq+oLO9BFa86bhYoskPjbsIdsErDPFThkcsp7Syi64DNwl
OcYww8YV9yFDPiZFeMYMp24zipqAqVmTJrBA9KiIfEbOAFBTjrkRA4D1DsxOYOtk
XkCW0GhKs5lPjhW8fih68+SEhdJpBqMnhqWoY9BhJM2VXvcTcLSSS399U3mIujDb
je3+9gllRm6JsysEtf0PnT4lo44Y91Vnn2LFpO7b/1KWa4pKjaxMqd+oMYmKvxlQ
hCkkpx7qywZG0p32NRwmGzFeKJZVcUl6wSrCU6hqxyuvl5A4cpIVSou5Y5yqPEcr
tc/FoEKW+r7cdqkJsw3oTVX7ZDf8/uCSjgteCeQ3Wpeal7/gJD7ppDdqTRC0VjTQ
Yqs+aXD6EZLqRtgrd5fNTQhI5EpjaMs25lM3WS2lgZ7TgqtVTgNayYT14Gy22FiY
8bycVNcfP+wcfa2lr6B3Pwqv/zTD2kXRlp5HRy4DTW5egAK3ambN4LQG82lys3zX
Ab+6NfKCh3TMupjNr+01NcUocTA4TtPfHjkEVsEk6OS5uJMuOT+drTnBCBLMNfG8
OFPlEkKWSyC+9yUzH+56FgDfblduBU0rlpGYGXeEtfUle7aEVkkChI0YrbzBNuf6
JMKFsehJzpZL83l74NrfGn4OU3vQtxICfR/wa1WuQhj1NBKGY4NtyT/dg5LLD/WB
EnIzN7IxBM+WfBI8hZHMDZNLxRy6o7vzGIvKcio6fz6XMU1phBxYblbCi89FLIO6
JRBxg8Nw2cnJF/dOzWYdcOWXvSTvr83EWBjqcibG0fGX8BUlD5haQTl3eTYrNe6N
xtLmgIvtYzvH3w91UJNSPdGbGk+OkZvwq0rk7TLkXE38tDlYuwx+rHA+57ROZyuR
C/rAlFIiaow97X2q3IEwTU1lClg2FSjA5biCJMrpOa3XDWWek8b5v7xivDv+6+4P
tBgKKusZNm8wdnG3MClwBt0Le0J5oiI674zyX5pz2Q5vGcfGu+66Kgk/8JDkB126
s439W8gQmaOJqjuGfYXDT0kidhM0VfHhZH6T20v2kBqGLe117QWu+kNIU9kWaqVK
CqDXWsds0XUWaVN9aCPX3wfeOwIthDFGw1dBC8lTobujTfQhKn+4z0VFJxlli688
tCV7CMEJev+vKz3m/wNJQxtdaTvH3SXFecLEBGDJq/4tb9xtBf+EpHrV2Uwl9dT4
TUUyLkdLWp+Vw/X02zzjRUWNhFrPl2G4EzL+e4qh4cW5Fn2cvi9RqT/TkNbYTbsz
KGBanW4CeYLe0QmsmiaJYWwlh4BVqaOUdDzpxhMMJbg0DH9/+Gh0oaKbUIOFHw53
THZgDZ3pR3jHRZ+UjjSNbov02YD1kbmqoESJR+Hv3SQsvws+4nHV59FQkhKhX1dI
6eooOmb2OI5OjjKbp91dtCZ51rEO0QhVi+hrh2EOxPrxuXyDdoqk0+b4WIAhk6JW
rOoO1uZoC9oL8zorvz37DSGwxQNZAifyQ7kLqhRm/WgH6b+0GBj6ICtIJnlJDibM
mDXaQhOVI2C3D5TuemfWbT336DBbm0vvHLd4bHT4FRpP6OOOe0elQpcflEYQ5CvR
fCwz3NHXvC7l4fKuna0E2eajQ+1QAmhfaASFhykeE1cADpjdkRs794Po9MSLBmqx
Y7A2b04v22LWLyKg2qw73DGobxvlCJfagt2sFEuG1lFp8Vow1sHMTRUjR+r4sm+F
Oy4hGqMOZ5Q3b15oLvP4o5/hfO2jz89do7IyVrIAvMOKD96sBz9BsVna0oE0Nm3i
DY5jR3ftJdRhGMk2KYyeB+vDB4o9xShKIhuerDCOO23Dxy1zphkOJE7obCHmYP6Q
0rQcQq3gMtZFUhEpTVoT6H7xAT0uDHJUVgXW9MxFp1WlT9Ags0sEQqnKALDeICt0
SFyfl3v2kfG9G61vqFbRg75tGOoPXGVi6Iw7mWG9M8BHPkxuPKNCR/ifOsVuxPFq
Nsj6JkPG9B0R2eKkWICKqgMDA08mA9ZxkAwQvqE7uv2vOqzx+hqE2fHSSXWRWvbp
Cr0S/6fCMB1ZAH53Zsy4lvNU91TMGZiRXfSEVZIaG/SLjG1ea+KiJNl+IobNX5YS
v5vsoHKxH0sq+kWghQQcjLVBsvXHJZWzsuUVlVFYmCv4o+aNVCM6O6buzvi/ALIu
ODGT46bhKxjfzmZfH/6jMhYcNJBx2j6IeqACflCObTqX6DlkY/dvHy+yu0y1Okxp
EXVZI5W1U0CjtpBliLeWaL2wiq1HlqBf7c/7mLuYW23T8jz7sD0pSMlwPYPqvZD+
wmcAh66lRU2kmMMheGeXjgEkpJ1UajLLv4Ut6/CAHdfwFyn7Y3jaFE7VA5yNxE/M
Pxa1O29SYbNyoGHTGdf1pd40uBVwlL0uxVNhxxculfSFyQmQj2Rm2Vm4+oywCHaN
1ksVUrsiKR3qnfRLPnRKghFMATRqT85+FlUrLRllo7vhSCn+lvnyfsCrtF+gsodO
KQB3/LZcApj7GG5L3nhO7mteGy+RHN7NJPmgGuW4cr61vF/Uam5d18OKis96yNKC
BqD/xMkTofHcqNsCZIX2j/rVLQagWcsynAVuvx3p1vEAeaia+4mGKYqp62vrTyy5
GizLJCoZTXIxsSOO0fMfthYkSmCpgEKaD625/y2na0V7P0WT5g50C4klURCFqn2P
kRmVpz7dW+uU/ltu6PiaUFVjoCINPvQiuI1glgBEoy/703pUiuvPJxINCo+0E81r
5udYUsl0erSUUfp3HPQ81CrhgFlzzWSMZiTizSJBUmshFIC+HUugcOuXTbuUqq8b
0rBn6wRCYrjh1Kk5gQ7g7+Zhg6eVEQrTH6cGI9ws3zq7WpZdRAje7Ato2KpO1AwT
tXtJ5lswGqPPoXtGFDbGLy4I09BZdruUXbYo+Y9p47xUttQG3hxEQjNGOol/+kDx
bBQLtVv29lDJhk9EBjDrXOkEuUyFJPIMAFVnT65VcCHDNvASrWU6mIJZFLUIYZDt
mWDYkPwfPFLiZvly9EyweaWwSdVdU8vs7UVR5OcZBpQGnMl4Oz4WOP/PmQ0htSKT
1NIg6pGNV9G5kKYrMOdAyb5nA/zPdI2YbYo/dP0losmClyp6te/e7uocno1nKu2d
AUyLcP25n05jOShvlBu7VRO9AffRlOcNn9nULmrtaEv/TC2vGe8SYcsGiV9L7Ehl
TyxVDl1YrYYLg9XySo38Us5wRAXD/xc7LCpqbojk6LGAnMneqKjfiKR+YjXQHAAf
DqUWcdUMn0VpvQQCHRgXPWuTjBJ08CQ2v/63JzrLac1eD1RuM4BZAoetkLmiEGie
GZBa8KIpBmG48Vnmy1ZKqSPBAJsrN57DcgOXyy/QPff2ehXACrs0A0vix+Loaa/V
RUUHJo+yUSkVXB89rRHi7xUjtxdQjWG5iH7rkPlndwKkj0rfUQN/D+t0a0qan0lx
ibFXrLZ50imXzZ9knP5PPw2qTiXlS6k183k2MciawStxwvBp86BSwdjcba/oYQjN
IJyH5gRqlWb6WhFyOmM9xBioQaAPnJON/0TtmOiE3s7l08y/+33HfqNB/aASSoIV
+z8IEKpuxdMkjgMAomTBxMhgabeI0Td5kZjFpG/tVMjW0BpcRcTrguG8Lc/D881M
QPuDFEGqBdZC3BwOM8R86RGsuFRu3oOYHRot4U3hkc3ftT0inY660LWl1Aso3Kav
Ycx4+YBV++BDQMeGzduvqdE4+yYYmfpRtibGbB+i+usOsEjIELqqRv5F5Gs++PEv
yF/4dE/XZUWcf7hNZnmUSKqV1YyCZXN4SJYPi6zeLvNr0b1D1/fMMCg/ieg4oEDr
yLRsimaJFHf8YwyYcupoNHSl6ks9rt3hp9bDKsi5+jghDVr7rEJimH7yvnJ8jwvq
igG5IjPfdf5zWypBYTkmYJyYkU7UUd1sG+3MoxJtE4LBRtZvFVIA1pzd0tx6KQpA
4a8Uf3SiE9kxLIYE+/NwBM8FSe9+ezJq0tLALBriy7Aj9P9oITMw5IK+l1BBjORi
YZLz0nErUX5VVdRZDx11k5YeQdK6YuM+loL9n9JTWBagK25TZ2qIOxwnt4rSB5EQ
B+Mr7+PHSyJkF5NQ80Tlyz5Y2ianbPm7wUU3ehS+DNYxFC02RSYLf/GsDVeJfHvG
ysKU6cSdghTrQ+Eh48/KD2aITL09NTuNNnMANtAv3trLaGMFET9ac7IZiZdasbaS
4Ib70fuH78mk1AV6/mxcj5gN6cg6w1J7AGJGVz630JQLXuggQrJfRqMpC6cw1Vmy
1SvwMykF+Kjeun11+BTILp17hq0k/OOP5GKmPP0Nn+HbKNm1EEDOtZ7DGMRgFYXo
MR6RH98NL/okxSCVzzJz7zimtvtv4RsVv6tdqRs8m9NX2TphmYOMdII5J+5FKay1
82HR0Cw7hj9Qlto/fYONj6rZwHs4XVMS417rBVEvkRN681Lh/JruwRIl8GwlakzS
ezhVXEml+Lojware/HJJFMGFJ63ywqq1NYCL15PQtmCBIGjq57PhSfB60Cp3BTiE
dd6EamwkgK9cr0pQr0r2wzJ4DevLWGybRfscrRwKx+QZ6YvajOWhpOQbsp3DwcNF
vW9vJoQpQLpE3z86SaFH6mREBEJhGTJc4E8+2HKNk/D74JRUXocgrKqXKdbXrvxn
OV9GgqLRD/iPcFTZEV47RA/0k4p5JhxNb2Rj9sly2OiSzc6RdZ0PGQnCyu9sZExH
vmoMLHVtefro5i22nRQW6MPLPBDnCwX+SJs/IwOZpgcIaw1CJWZClL+JYcfeKH6C
hMkSq0hEl9sroPfkro5/Z3Zqody3gLo9hJvZ3Xnh/cNNXpTrfU5rtiaSvvtvK0rs
v5eXvxTem3e2tx6EwrzM95wDY4879+vGH7MaNE9S/5gZgvE6rTQJaPT69OmCd2LS
clXr5PmYI/DPxiQImhGNo51Ko6Rnb34yQDgnA2XxiZG7AsA3emzo+xc4Rd6PRgi+
iDMHgfVMlECSgBjuN60ETR3k3rdVQ8mrC0JW+3A0WG+vxPi9XrInJJIQbpDvKkD9
YO3256OVyurZ8Ob7PPo0QFZorayO0h32Y10GDkUjCymEGMrly4C1X5iKKnMRFPVO
72heDN2CoUhL23lO9yroxnut0kTlmdQcqtPlhK69pMJtTB0uT57RA/uW+Kbmu21m
W8wOhlmF7NKKsAhypgxVBo616SbijaN/ncYlMrAa0fZL2gBsgDe2oX0ovHI5oMzT
WjoOTXOVN0MXvE+Uy1l+SH1Utq2t2BSCFm/seDQY8Vtuc+em1KtfIAq6RhIilUqY
BZX5VuN3hQD7vyqS3qxHVOwXUJcLpvcT91utCOUB2OThlSCcacG6mi9RY2RIanLu
muKXEtlW+iBUEpjlGpYmL5+8/QV2K2g79TYQppY7bRjr0J74/GcV0pq0iwPKGxc3
3teUnzd/4NTtV/CMF3NAHyjECEzKoOBDdn6j7Z5qY9HUigGsgTAft/M+Sx1nMmio
OAY18PdZmDulCBixKE6yRGY41Pimn1EAhcJWjbKBkHs7St7xIvMaQ/CRaZS2d+6I
UrDe97maqtXBCDAXjjIDn0CEaLhGIiGAkZlI5aS1WescbSWz/nqWGjXsXUqb2pEr
7P2DmDLdRlS4EZ4bKQWKhkqfnbD4vfbe5d2IyMRay69c8OItulbRF4SYX10EGaDq
oKGXdiDkki3Db0VCPZO9et9D3fP7BHg1aUQZnAzGBz67RMNAt0Tf/x1XenVll2oj
XVbzpDAnRGDjy97tVeMnv1/RnPZpkwcdFl3qjQrw94ERyviQwJaC/3Nt6NXw7vq4
d4riY6cOpgDCrxAf/fU9c3Gl1tmQZ5Bo74OL4oXU5edEIS7b67AdYX0Zsge5pne/
eDhQrp5lp33STNgO9lVcB4u8gQ/kldShhVhW5d3npDJgP+a/pp2jciujjI0nlzKr
dbs/fjQIbyK6dRv7X7cRpsbOSkomRfNqbS/aqueKx81bl3Pg27jaHtopBwynNZLU
vSmO+UPMA6V28kr5oMq0VcN+xdIAImqsN5FnFe3aemu3umz6XnyS3W9rNig6YU5l
Shuu+gSq0AMRjpHlqOvo70++p+6eOJF5YM+Isric+2AV3anSZRMbRsZMf+u3zhCT
4I3dTLrJ0tAYq4lNWa5OTa1UP5eBv1cL3m8rbClRHbvsPOApTEKlaKlOrToKMoBB
zSKEayAG89s+Z2sXx8llogvIPx57baIvM5nwzY/RzS9t+YFxN9CartSLJ+p/G9jN
HYUCZ6QtTmALcliYBpLoSSOZ5jZJ1xhv4Ijpx0wfrae5b82TYkxD9kx1eDel0MsX
24FrbxE0XK09gryk4mieJYEGQ13qj420NdAI0TNQwp8/Sh92poBEhbFScZ8jlgQw
TJmQXPhYStA8iC+aKeHRmvcJYrTYGdQ73nHWUaIbMnPjHZjzSUFnofUjdc9oVStx
Vm+9B0OxVCYMHNZ/G6fGoYFFPiVbL09uwSrN5+8r83er+eA0prBBS+ITNZNapDJN
Hw0DVzLpVeKuBwvcvY0YoNOXN4SHpkEzRuBvaJ+46XeSn3dXfL2MDbZTEnK6s5rD
YxooQ1T1yhcClcWjgVDtZQK6HeCOwJzDPzJ5FiBRoKtT0SUH2NJuaDmBuTGXq+Ef
12PRBZCrP7VIraX/csycL2lT8jzSpvA25iFx2lOBESvEYqUTIl3CMNC43PlrCS77
LG1eBsUbXAOrFFloWsSLtrZ9mMTw+1i+IQJucMkfh2nFcqiMW4KH6xR/byJXMa+m
KnPSKGyyWcsgg5jnUu9zW1KSTUcLsu1OgfXFT2l0CUgbcP9pjYR+3hYqriQncfDA
aBVGbS1tUsFuTDcdoi5mbv6+rwHOuoW3bF8onE6vsird/y917GtkGS6cTiuPrQpC
SMaRPUVWTP4PI/x09z5SlVwiiDjD+iEGie4nvY+UQkw0IERIh0KspcAUoQMdbIIq
Yxrz/mqHCLITwK25q1wrQ1w42DCQzhZbt6FFCiabNe1EER/JjGARXQT1j7mtexhb
IZUdse0OOmQWa58VoFc51Hsp1Qb4zPI+OEFrNwaDF0whBZWCt15flihGszXJ0GkV
UUxCmZHbhqkY0FijnxXdJcOcEumxhnx7e8Yhc6ZDul3p61kbKnpV1IlDn10pqTMm
DNFtbGW7hJ7hqKWtpTHUwLAiLq/6osE8gD6TqDTi3gq7X4gnrwTvb9vCYsUusnOO
30SfriIFdRKO9h/djKurlRMFPCLMwxGKXtpER+HcGTBHkN3KbvPZqea5z9GyBUli
d8mmkxmNxdqeQHBSt5d4QKVo0W5sxbTBIE/ELPF8Kl9Fcc6WBioEtHyCG/63F1K3
hE6XNxZQxA24EoCzc95vAJ/5gylJy0erH6YsxKdmbbg6U9WjeDZR/K+I6VyW4JkN
Pvq11/zPsLU7SNj1LQpOGNXCVeZ9LHyumWIXPgh4IQxl77AUzeFyUh6dJyJuFdHj
W7B9Oq3Aptmz/fX5nHfjYio3uSysvrDLnD/EOGNYDYJgmqZTlQ/UO6Ijliu4m5ih
K3J2yCJW4mS+cWyOKqLcMZZc9f0r/DdallWKOe54AX3wj3KZIlMGPig90Z4OuhEb
VylLJXHAIehOZv0tnf6h5UPQVM0cHEnLa762veDsdkO+GKAMLS0az+61f3kP7ewv
RsmHUUepDMr/roxk8tcOU2PGToXuZS8l0q0jUrxIO2ItNKT94vTWY1kRPfEnSKjE
xjlRebUEXsOtg15MAJRJyvXvnCSHroVmgU6WiYkX6j16nAjuyiJSRWPPXndnDiZq
lBCP+SbP1608E6686wsUMpOS42kHKwud9r7k7cjeCmsZtAkh3WQxI6Equv4OzKTL
gwHEm9RQmuDTH5HQCpURWqPF2tgY+tJWGS2wqx3U1oZhCcrSu45Tg48yBlAZmLhz
Bu++nErtPMqOgrcMnxytp2KHmm6uEsWhvyi3Z4KC/SKfDdwvz1BfbIkoF7Dm8CEU
KOQhSeRwMmN5LDQDBPgCmyyfCQ9eIx3DXQqk7LmJlilt5YMUHTsMpTmr71WSHnPX
OaCYkneVUs4FkPkU2bGBq3Qsx9zB93nQ83C/+uDGlae59gMJuuOjh7Y3y5L/nXkC
2429x/+CH8leyS7qTVzZI9t541YOxouRU5f8xIUz3Y+fT1mv7Hzt5RWCI/V+nj/b
+tqsvNECuqnN+WtS1w33ODbuI+/uz56zWym1ZfKfbVbndg0GaAuHzU/cs/K/A6TT
w5CgOujZBj2t+Ur6h+ZciK6lQ3B5GSnHEtKY7B195uscQYBDvh6x8RVX/xjYGWzc
aR0ti2RN0XuNVomBHWxOrJ11sj+CUEnl2/NE2MdY4HHFFffnvE86Su91/ovKtUdb
C/DHKQnSFDNySTj5oF54E1W1+EmHNtlvZF/px9jwdpktcGzlOukKFJNJS4sSZOI1
2ELRhW+eDZEAqu2wqsjlYYJmrXiE4Bq9bB3JgWebKqzyPmdPPYP+QHRsHOr5BJ12
vEekqkchlT/HPTpODqcnOt48P79Sl9XGeUEy0l6Blj/2Y39u7OQ484AphRnypHsL
SaSHYVT7Mw+v2QjaY07V703AjlYf2pmpKDh6W483O6rGbLBIdjDO3nzl286LidVW
in0nLO6ZqQLYl8LzWIi5uEjij4ptr8oRVA89fisEw8n9uLAVavVnjBOx8JnTGA0Z
6DSDXRsG/P0ZZqfDOu8ik8YmrhA39DV+yYIzpuaHWxj3gFYpadFgi3UpaGhRR86U
4Ss177guHvaBMVWLVJd6u1TNdjwjbqKco1DnF36NK7nzv9Z3yLQngOyE86nA+iPy
It5eozRk7QffhwxCewedNnoOInIJkkYO4Tqw/dbspTgwAYT0I6OGhXmlD7EoVqEO
E2g6ThxbP+sr5RG/MvqUzM5ilTs9wgmecr6bafsRxOY7haPOSFxxc/sPQR3Q6G+j
v8SOi4KE4XCzldAw7RE0bslFcLM5r2DuYnIa0+LcVsm//HD8S0hFg8io7CIZMzT5
sMmy4kkxFlDnSWQQ+0vS4C6yfvawIWf+ZWdLKMxIsto86ou1o3cr34vqxou+nuoV
81QgI9J7Az3fCYWPTYMaAisg1ONAStsACK/II8L6tZMeTGx01hNGqR/niVm5Rz21
t8gipxiWLnWQcJ6HGpdZVya7yfZgI8bqPapcce6KiIo2++IhJejQuCpe28lRG4Ya
oOtIhGp4QWm6G1/Rl6hHTDb0AkB3lvYxakMIui1vrDenNbTcjTRPly9N2tewyHJv
Wyjv/wKGxhqu3hEQibfQYXht54TLPDnD/fwJcikVqr8x7sOeap90fV3pGNrvrxlS
SEMvPCgNeQFFnjZBXILqkBPGYWkPWKH4BwW1WNjIl1JexgGvoK9OXrgCwEjI6mAQ
GqtknJJIhP5TwG/4dsTHW6w9U9osGcCwvWiP8YNyHhyEtiZh2+q4tK3OCltny3c7
YXwKMnmRgLmhrzHfPVzHd2rkSMD7OTDS/saelcW9dOFnH1ETKtcUg0VEA8CMrOxX
HzqVh+UXVdO7V5RbgKzSkHN1651n9HpxShnkm9OpmL7NiN5IfSTdyohxKk7L3UPq
psEkXn4/lASMpjSmcj4CxxyyoSX4DqqZD+vpbwAcU5NBTBRVRDbmS6i8fspUgvDe
xVsU9ET6mSxnjCNDanTFaP68G9ODQTOUKcG/XrhurP4fgfn30B6dDoKSkEfWk4NK
Vx167d2FKqHZvM/0EFGGs6md/ToMHZQpEYeWH+jHEr1HMZmcRYZkeMx3yTWElEXJ
Qp3NHEeTX109bRNW7FAgDhqPZBDR6ahXB3v6KCwRh5l73u92sqYBXnUe+VTvlC0F
gL4szhNvPTMgmU0SurN9W6G46gU4lAhX01UUPplYktQgba6zM/ntur4sEnoLhIDb
1yVd22fQuCRha9NOOtnXmoyENJ1uuiVwFxEkXyu9O8GecjsRtdxlcNlhdEVAluOv
t+DbTkEH2W99kzZdGJ1vgsJQLWcrbUg6B6uelXVvwUUOXC1kcJsvVWyuGIvvamnJ
tq/UpNiLL8/S3hY8R/57MHujLe/16hRqtwN4Ad3p6bFKbFvJ92vVT2cqaqb8PaoS
xcnWql8cKiCyTpPwiMb3IzuIIXDN61nG/Rh+xkjzim9i9sXiCGzIfiVw8Y21AxSB
lfHKktRtRgscnmLSYO1Xc3m1Z/18HVS+41SyYf3OtpJK5TrVy7H8cOOW52CpgPMn
/JbnrXRR6MBA2zys/FkiAITLrzC1svu4O4SzKngoIjWkctmrZSnqO3eeDAf4mXki
8JYjpcV056gW+rxFjsJGkqtf0Q+myrDwzOfOFNIm67MmbnluLHB1AX5stUOz/nOL
LOHv1XhH1pS39bJRTlvXCzZUcz3NNsyneU9XvN4r4OjtBkg564wEtgFi0q7qPoXq
/2/JttPykfVqgQkpJ87ciPw6l3JKe+mejin9cgFvXVKOSRZigIhhdNpT7GIoNNRI
25eqdY0SqgnA6hnmBhNOGZw3pp0s/yRYLjsrdgYxt1mWqx7K5JGj4HbLbfjs0eA8
cUMVoEPWlcvRuWRI4CrrSZhPZgTzESiJ5O9p/NPk7I99V/3qeHH1jfdC+7SJals0
uXsJ5vjsjtFsr6xRFKVeSfBJEdakX3Q+ZdQzOXUEHULgD7dzUv7mL+vx5yZmecyG
uTWQOryFG/vW61wRQ7KSlp6r+lM/cYAcJHJSYKNlPE9G9I9aoR/VGFyPGT/Nsl9p
ydyveIq6zKoX0N5GRz603wzPnxVumC1k2PrDQva986eZcfby4IETN6KYi6+bo3iF
Potpjagrbv6zpY7dEkJuu1JSgMf3wU2Ew2Pzv6Fymy7TBR77evLTzsOloSXSZyPh
Uy4+DP0CiouLZZJEtE3XyUUMqlesbOqbIRFNENGNKp1Iy4DeRRaRZ/mdIfWe66LN
ciyl4Ktj0vHLwnftP1Iv6I1RZaZvRlcwzLDfmebpiVf+cYS+/MNZWeZxenaMfEva
AzkU/52HxO/xNDeDgi6xYDLzYCq48PRJvdgYIFRhdoSOQl4lLLMdj8/XpIn3Rl00
U1NSaNxqYWIIFMg6DR5Pn3RLXXQOC93V1AS5IJS2yeSC6/BiaaFsa/s0k/AQuz8n
fsAXH20phXoRxi1xJICgFyJyKYMD6TAxm1bUNWD8DP8jkKrgL0a3QSyJ1x1Wqjjk
iI98l40+QoYF2a+f5GdbwmfF+mKE8iguRPICr34odt3shgLgJ1pBfw0cun5SqDdT
WaT/E1dgGlGy86j6TuGxntg1NeuEuxYBPiLv85yPaSmBL0z4YZrphKe9wy0WwfhS
xJgr1AT4r3S5Qlx74KUKpD7YZ4tTLuJsPJbXqkSeIDFZ1pKyzMdLQq97yJTkdmN3
YK+9aK/kFzwWSXOzxKiDE0xEGs7yy/wZUF5EargB+LnhaS5MhHCYJHKDx9Dkvgvu
6Yux+MdnbVGUJYOWYZKLXNhQko+dJiAHwfGJv3bhJLKuYPHdWcAGRUvIoL1E1NPV
Mpb17xPn8DmGJgU68+u8hhhNpd0mtHzXP2A5+u0xayvfC+00Chi5dZFaiYGqXyM+
XZqJ1ttiyga+adE1prXwacQMTmJVktTggfhW2o1hXn/kMH96jo3WGCpY81oKy4hV
/h6vfuO6AkgwmF2T+9/5TKm6bipfT3H4hy86mCH567eecgM+g9VDtpMyiXy06ApN
4vB5RKRtcehlWqQg53Jo8bVFYE6IuPJOZ4TMw9i5X3AW4Gw5vR/FJDVXyaDnvdeO
0bcIyoHAba9lMhtUd9e4n4aZb1MjiTw/bT0iUHxR7r4OjtqCTAW9u366Mj26CIzB
LPb7zkWbaZUr+QKYT89sqefXr4gTjLJLcpbIXM7siejhKDnTDHVfPTPsSiQQXG5n
fOUIny4DNnCFgwKoK1/lQA7puD7NKqACaTfLm2yHv/L/9IxAQyFHY2xxmSIrjIsj
21wVfhfQjz65rAInR3bipsLzfUwzxMosg03WlHUOFyYoSRxFGEju+ZdN5z4gFSk7
U+qVPK4qnCPLUshnCxknpHHw3xlJxOC9CtP4hkEnvvTSG95i3lhV0Lcc5PB0Oy3o
6FfUyYCZ3QvG502+WmIjvlkrN7m756CYnYjuq0QlQlABUXz3TcsClpNHErZYlffv
xdTUo0qi+Ps1I+ZsSBlGK0HX1ZPGcVmhsriLvpIOr5SYH6YRrJOFpHqwZpHl3oyb
/6EfhteYVUBJyVt9eHmBooCUreFuwvhtZJlpBWN9PPNIWraOmmLw79n9LtAF/jHv
ct21N8mm4A/jSVaj16cm95u7MI7swpYQlWacoCQ44ZaQPcvyGThxakh8XNRPYX+M
tmjWGHJYiYjfFOilKAXFvgoq0RzEBkI0sRrQT80PH9++acBb1RPu5UalAZAlPvd0
HxSlviXfsWSBdRbhRzzjM5TbN7WT+SOEdy6awPB1i4sxz/UvSsiWAqrrOs1VB6Go
lBST+m6ZqugmJBLdpOqSdL2vqSVsFPOPX3f0XOP57TqLv75MuhKvXXgSrlsmFPJw
ObyeW5cI1le3BPEm2C6gLmbl3mdT8tkVP1rkPikzTdoiRGFt4bojd/vR/aOfZLT8
zuBPjZRLtwzuuIoCoPX0KNaD6ioDXm/8kRgEvm/J9J/aix7BU8s6L8Q5KsF1nNrb
vtY6t5E29p7Pv12RxxhzW2jExpzoJMH1kmHsIk0Y8MrHs5SbojzcSbdlUJgPrw89
1aYsTjULQk96rbnuAji2NhxY+xTDujIQi1bhzfr3ZYVl3SHSZmnlZLz6bBoqVjVA
LfULIQZi03ZccXUHMZLSqhfTKhs883tmlQfk7DX9/ZWXWGH0Qk8VvyJoHFslZ1Sj
Gf0Oh9+5/tjpr1jiaipEFTuU3xsQHQU/mJvIQfJKIguv81mu+7NJttF7jsQ8E3Yu
VFidT821u7/6htnV1i+zut/6ispt2KkeeUiy0Pn7gtFKn1VCqPWtLaAajHgmtIlF
azQuGJacrvKTufwEXnt2tlVcO3n3ZkLYAFsXxBoe6eEU/slSaWULFAsKyuPNrAfp
cOIYzASNSXPBGYV4clJTBstJmrbaCZBKK09eTyZUvIGGvQSWJhpME0cdC/aok0ph
xsLzpnVIfyZvO43JucJXmhtgeJRSA/8ZyVQbyrAMVdgZ0IWOtbMDCmmRQYJe3xtf
BjqYr7vQDWz308/SflJ4f5Xm98tqBODHC0PFTT8ywYsAxqp38t2iz9vWQ7XyphOH
W7COcaz61Qs+DfYF3W+AiEFp9zm/DGiQv/VMzFnuEidrHPySp/bM08VIYYjYebO0
zk2LgQ4gcI1Rpe3SIYuYLKyoul9FOSADJI6hWfDvPGO7YixPAtHRbaxnEWJeOVVk
IW+JfAOED0besXRJwZW9HNje9yriJLZJCfAhMHMCRrwKM0GunJHsjPcaBEayQIrn
MIvgRdnRNEfM3gS5qYRSgibsI0iw44tYa9DOtpn+wh/7SceEgpHJmHUbvOSH6ewb
0rXtDSeKI+kDjfhiGEtVTBuVEEAF1YSygQ3OsLsZ1c6bHHNZxODiR31r3WDlwX96
VRkcZCQVL3dagn50yDf+Be+VNnyOsT6Gv8Qg5F4xYyBb5LBJvUznO8TlWEUc3DSK
DjJTzCylU9s12jJNv0Qlf7TBQIThBH5DGuPqBgiPxCVw5xuYaBmdVEu8X/EPtlIE
/pA/eH8ht1ihZRLRXqPO5bzE4BuSaP0+Gg9VbY2Z3rqklrDV3BEyaq4/JZOjiSBB
pnHtQMP21euq4+EDSOr3BMzSKikYqeX2b4ld692r8fmaV2lI17gTTjIpDnhDJMQy
KBFHdTsuXoiQmXWTrxP8e5JfzGarCZ2NBP9CfVnch8M1SBCNlzs3sb9CduQAuhdC
mxErpVVAfre88kDl13BiI6oeQ3D83nlwM4n4zrQkN1xRPOC2R+4eI9o195JDHaVW
Arw+E8S1mvcOTDqKYIfdPIeNzTZIqfBBB3tDYnetDRmczWeCY4ngZDuIlgluIQcq
QIlHdfjVtHkbFKVM8Xk+eAIr7qz4MPfHsqU8eC17b3Lsx6jMn41WV0qobBosukKb
TPBzIFTBf3YBIOw0Oqg/Jb7FeffEsIJGY5/2leqtoFJE9i7t33DksuuJpzKizFM4
hSh6/5hxcEHjVaR2qgXXBzMmEn+hqRWOb3nzSGOKKgqgkhDIZb0TOj77UvXE9HqX
zumqUE1hpQnn9YHH9HR14D/Oeb9q0RUpoyU6RZjYNG5PAPE7rbdSKdZRj8koAFFP
Lo+4ekZAPhjkDv9InY22b4fdHHGm+M3lMHpzCs4LrDTn8YIB02LFqxjmH/2uZXBx
i69qeYN7igYjs9WhqcGtb3HgnH4oaivcunx2mQ1AQsm0ZGw0RR4UIiOuufMdBx5V
n7hnRFP8NMAxeOIG9HeGfbCKShMZoo8M1LXO4GvY/wiVHQQjq+a4o2Swz+Vj4/XB
gUB8wsHQrfgig4lnAqM8j6MOPbnJfyyOmQpvRDvWQReL0EBWBs0Vw766um2N0euX
cHTB4B84r1UXxYsIqjEoXkt0NNr3dIv6eSDQcsG1DggEAubsmHtQQahxNY+GuW+A
pARKklz1CvY358DrDffgNU02ciIrUEqv4M3XlFfH5w20RJ4+g/oa96szFhdmqAWA
9voTYi7ZiqMYyXHhJMeNucM6/ENIpi3WC1feSZNz5HPzjAOQCPKDGMhdAHy1T2Ys
Ohrr5kjFs+hGykLGrDPJ2Dkp0mtkzIPHJ2VAUfK0/fH5a3TvpF+oFf0M6cLPyVti
E3Q3+0IZYL47X/W6L1djQZWi3+md8SXcuhp5h5oGVGUq93c7H+HRSCxizJmNoXjW
M4ZCXXWVcrKioW66uYUmbiZn0LNR5IxHov3yodBmmPdqcQeCBfSa/CvtgWCU2aMh
LMGkyGfndp/qQScesohZR7t8zy+p0uZn2elRERlg+JrEBXi4e0FI88q7N0BhAhjM
Q1CSaUem7nFljNiORSjMfEsbzhQSD1rlsnbp9yCrlL8UeeB4xCl3onAg/tGQaeWc
VJTCJzi+pTya+Ab97+lb2C2sRNS9mr/zoesJZFpEUzzOrYgXFwQtcKwgBX8mUPCl
X+UvGjIS/qYrB3WLrQ0LN8SvaEjk5DNBOEY8xt0+CVtQyX0RlteEUEfE4uCgxEzf
/0ZcDP9U7PCHq4TnAeJ+zm4WLN4ws5NwnB40NNEFOQYFtjVXvgOr2IwLmcUdDdAA
2e+VJddZtRM/chvyRIk6r1pX8sbd5Bd+t1AlYLOZyZrMH5DVl58TbkUEpncBVKep
5r3tz1XYL9y/gGdYe2/htEjj8JIjY0RaXbyadQ+6yNFyqXToaGOSvNxILa6GI2nP
pnB8xvR9MSsNAAznCW74sCPYVvOXCdzlLSke9UbUxzvG8tn5Dgxapx72gTe/BZy7
a2IlaRwzuwOc1pVGjQglzF7Vd/1SPRQVSMUtOF/lKsZg+N1BA314uCF8hU761/i5
f38TV+WwYW2X7/VRn+lKnor5aJGwcmqqtzaaYQX/pL2NYqT+c2MJ3ktYmtpWlSpr
UFzMCPPlVqRnGSDib9VnMNUGaX44RVTUXSL2XfkYttLEasIyosSz41+IyxVCg1Dk
yF/i6OiwORNu5kvA6bF6fHvofNgcliXzt+++YpEIc0rToHD0muB2WDu7kDURAm3V
moM79Ww9tKAPxLGfJZIO9VYFDWvYhdp4aOsm19G0x8HqCkc2HLwCCN4cB2ZazXA6
PKATQOjXJ9Y/YvHR+ltLVJxxYJ5t4J5A/NMa1MY2tgX0O011ZKR4UOu7ncpoGvRx
OK6jWc5yT1FAYc3Zo7XvXOHcOXG3kj8AkEUYotJH2aU+meglvd3CmMEDjBTew1bG
apfsmtDhGdCEfizks7kmCfftCla/mq2Eln98WQZKBUYVwCh497uXE+VW52wSxMwA
1I3dBDUbwAmlZI8w4c9DxJLN2TuKIua8Q027JjEDCy1qfTe+gUZgLg4nx9k5C79b
Cybxka6GCo7FiTzevGHl1nI0PLtcuCfdDRWKd8B1MUTg3WQb6oVrLlD6hAUHcFkS
nI8wOI46YaVGy4qMv0LtBtj30BLI8rUAr7TC5iUs9Ild+dBZ97L55MnZfKKrmgH1
OBrzSzI3kpPduj/txJASLhv0MQH7jr/Vd9AmCBdIZvRr2J9/qCBMPAf4Qj33r7pV
Tr5GlJunH2rVllnfN06VPbDddOPoIzxs2czV4K3xf3NlH2ASKjOY6T6+F39ZFuTe
tcXSUID1NrGyM1Bv7zXwaZiU+nL9KYvIWy3BbcChhpwzOX6j4W5e4D48WyQg2BjG
nEzGTOY/r6xjijZCPUWyr7oTdVsVBjcAXmRWRviHqH3Q9kDB8HIjMcrAoXDStFxV
VK/w78qmAVZ2dQsHYyKXVVKOv4ndw4oMqPr+x/hx0PbXjDLzYP3xC3wklgJuLt2+
oV0o5ro31F1IB//pa9YbyKV+lOmTEIw4+2OSihSL9f+YnCbHwPKGOi/BQ4Ac6b3z
+jCcjHR8PytyiQESNINxB4zv7ObgHBvhOBGdWBNtnUbtJxnYqR3Sv9FoYbgUK8r9
+BNGoyQssrZQf4xc0aIzjZEz+LtmgTnxSEKvuS2+MQQv5w5CY39ZbXGtgeev4l4n
tVjq1fr5N0TobF29vIQICczgUJhQr+zrFQNSsRVFxOEQCQL60gWh78ay0QILqUQ9
y221Lez2qkRzmL9rt2W8oU153udvQ1KNGDFFwFHj5qFidFmCSe79Pl9mjqNxqnWB
dI+p1rCAr28nV1dycZt8pQVs1NFBGESpXGJLHi82Hv3AT9BlJ/jB2sp3aZNC4ivS
ck0diWWWVhWW5pMurAWozK1J87LrRNPdYMae6TXZFPTe+ffXjPRupiIXL7luK1Hl
/95yzLV54oIzKWDW684DDHN2l5ErU/T1ZDwjZlDzerlD/dNjfeJbNVKOVJqGIo1D
rURJ5q4Bq9edp2481Utc2DzFlRzB0O25//r5d2bTlb8+0Q0+PNkpeXGjDiEl6xpJ
KItq6Pccn0JI9BKi/JTVf3iyv/oKoO0n4boQBgBN7G3Tlzo3CH/CqPqUcuRNSteq
Fnw57vx+NolmgQMZxGVx4NPnUg22NvcEUWgXJ/RrWIqC/zAveNXB+g2l/DBHXXum
KLFtUlOapMYLYjtkJC+EGmAD0OWg8Fxo5zpKCFdjaeNWYhfNLfGzfuYWLdt5B+w0
3tsQ/n7qCj5nQMZ50JeJR8m40aksNEasZnoDPRQqNa2P5k8fmjdnPuQdfotI7pCh
26WcH+NbWFyo/PgmAAyJhDmFf0KYZ9awghLTrapeiP6fC/xbc6+nMvehqMrParr1
IMYCdXciF+MUtWFnR+lZIEY7rO/ZhDI3OnCKurwcaMJYwV9WVRGhBw7lkdjXRlB/
eF6iXrhN7rVromBtG/uq38LPb58WmuIVFaYx+T+1UAUcv69zMfOIAmOcoA9JSp1y
fzM1zrqGHMpwLeLcfKlNDc1MDPA41I9bXk0cwjHL+SW+1nMakG+owJH773f+XP+h
x3LYO2ybdy2nlCrLCh1Ry2b+PXsQtrSqrz3lBw840t9/malbFfqAauJNAG4pqN1R
Tv82p1esUfjtoTraCArp28jbbkpvUeXhYNOuIrqBGOyyqWDWCBNug5hrVFeYKAyO
rICM0AJeUAoeTxNnCJdSf51xjViP1PcHnCeY77tlujx7WZutvewXhW2ygH54saRf
LPbKcTYLp0RE8Jq5kjTjAz6ZyJWux5NLHhVNagEIrsY5E78ZDW0tEygPh2yrRGrI
yuUdoFczxZ6qG4vEj4G6LbM9CvWB7M9ZDrRXY6nvQnTUJ6EyQbSa4MTVSlYBaWRx
pC6d0uktKI0XLnSpO3KwSWsNS5rp/PwXe1j7zh3LAUajVGg87h56ZFPsfVVsYQSE
zrS5hAbb95ArRBLrW0zWdcNyoxVVk1OBk2PTrCPS4P8s/MGmSBPcMuYMXUbUvnUp
nkBJBmODcx4BgDVgfyqSAMerZSXVx5gZChfePEQXm8mTTBz+1YtETk8iIOwlYNcE
3NhNA7c0w11xcKCxY7SZe3vGVi/o1niwdGhWfm7DyKN9PpTpbh46L0+8OAOU+Bv8
Nugtk5q/3IZYn+J630QeiXHP8qKQoyO0F6fplsqhdK74vVUGq93HySa+7T+cCBUb
D9rmUUEerjPXRpux3RQTz6JK6PXarUhBRhXOPGxkhSCoy7JfqMgN4oPpvJf9sJwE
BN727HPPnCJDlAXVk1wooUBe9g+GzoTH3iNGCz3V5iuoA03n9Sk/BeTqeOrO8Gzj
lJqEFEUf81AWK6+2CbESv4TEjlGAPIzio2gaOk+25zZVvjusxz8q+ib7s5u3AJzd
7M0qy+lyZsXdEah223ZMo3DDWb+ySpEkoaKYbwbA4j7vPBQ8hSGQLvflztibRNTO
covVlBxuvSJkkVbhnedlXw6cEMYPwDBVaLq/SHdRSb+ARn+Qeryz7KxQPbVyeFVf
ACfBNHlOAwbIYlgVrxPEHQfxb5oAM8cL9GsT5eDqsY/hloIaYjBy/Tm0YRKl8R6V
TNbn8COV0U5sZoodxtuDiOlj1o9xvOhmKRwGKfNZbDXB+D92mhSaZCCvOlJprijU
NF1e2Q9+xbivro1di4xXSwjmB7Ejg+rVnjgUIVi3wctqsJkm9gC26yGKNLpRvMJ0
gvMLHTJ2sjmsAjdo/4QBjLP6WS9EqkFH9aKfE9eiK/zHbgENPaONEoK2BtGK2yqs
bRlwdaPLxc4DwsyxALWet5y8mZr4wgxF+LWRAHJnvge8miFWP4ArtDT3MhjLdFp7
IXj5uGzqPrBwKu/IBQng41ET5XhHNiFnyPxi7mz3Iel5RY60EWjZ8nstYbRwUR8i
oXfVNDt326Lay7y9BlQQdHWws4Fi9uKaMAvuqwxVXxoyf5hJqtGlUrHaWJnXmf98
pE+GDV5Y7zlmwvkXb96/LhMNdqnInBY4q8ttsiTvv8NzNLofmMZZpo25BJ82N7rH
1du0Fjj3+7fwvXNrsA9pG42jtyTfI/crYvzEtDZbOTpVuAiGlsGYErqD/OFWqHym
z+VNcRpLc0fiPlpiqVXohosWnZ+aU7r6HQ6J8vG/CK8Xoc9u4mhmrhLP3cu0jaPD
FHQabY+RUsFf7Tl+WtMwiqojW46oENC1ak067qg1UqltczOhZqW2q5QfzGiOMZUD
+f8Z2X0LxnUH7pfi0u34mdrdiGvGSr4vieXYqTu6isKF/8PrNqguKbfIMBsTeBNb
M1tcA1Qn5EkfkY9N/7CnjoLJDwQAyHwUqPLyzdj+viF755ZPx50PnfZFYUqAXiPb
hzkdaTTrBNWtRmM+IxA8J/AHyKBWfuuAgbWYjUwqrtm7k5bU4aOu4iJQstev81Rj
dYderM2qlPeXT8rvejis+ZXvZoLW1cYMPbXXUDhoPNlmFv8JrjguG37lr2IqxHm8
mzUE9inU632evXir3SeXfmaAwcOod9BxJepmf8XB437rWTm9uVV6YVHBNBNcX0eC
9cINHK2rpCwsO4gYj7QNYiSK0SoB6MT32Pkiwf7fAl77SwlIFFXXj43GHtk/lddc
MKdGg1YgzgaKuz7qzhkUh/UHEvWFe4IMxRRK6YdYmiTpRgfaJNXXRmn4o6EiHnTB
OUZTeojUYBdWb3rAKeKinNgm0xBkuEC2mrp3GxWh5hDQlNpLyZsVgQ0hMxGtwAdH
CIDKfP/78ErddRDvj1YtmznrrKet1DX4Jsg3wJSNWwDTNSRctgTfPCFunKcHN2+U
+fg3Grn2iDLU/+fN88+HCdi2uXaO+WMy8zhLxPyLU35mJfezFdb6tJzj11JEuTJc
S7aLp91yd8/Cbt1U2bToVjaUZ9XnRSKtFZQknePpPpLJNFrmGyr2WhVBan31ZoAZ
sZm/5Z+l1pzeIUiRI93tUb0f/dRrWU3t8ThdZQIPEcIrcKqOgN5xBVB8f4J7lj0+
BWl6o61p2MO1IO1RRTIHiloRN8r2+63vjAuOiF/vYFpPnrVS2EQuwFyBM8JJkT56
yMU37ZoWrSi35Xl6bQ9IAmUbeKdSnsyndc4kQ7IX2RBnkMkZlNGiXCIpigYIqzVB
mugPMSfVCukz442oZHWixxZrEo6jPjLlknfUXk/0OK4XDd/p1IgroZBbDbfOjloI
KgDEcyluituOmXAORX6aRi+8TXzEEoQwc2sRlIBhyDtNdWf82gDJFA+/g2mzTgDD
Kmjw/j94P4csyHD2F2/GY4yzEppQzsanEd96Jfu4Qr1aOlQKNXkk3yPcW7HhrAyP
EIs+lw5fpWsxhztU0LSXMwfusikL2s7GLYuISw+PztvpqYsjbAui/mleIBCR8x7R
djhlHKeOSPved03LkxPqSapPlTdI4riz2P+X7TI4L73vrCXBLTdSIWYCQ2HdDD9s
OcHT5ysJK35zv3CmELV0OgRy+i2BTEeKRmFwBbORnJZ0XH1IaeUjwBHID8r0a+NJ
C8CzDn53IDp9xwlzH7UtSraIheHYrH6fFVBGN534yqMPf+zvd+tON55joKWFBo3i
YwQE5yu8/N5trHVzcpm8WciuWuP+nraTYHYhvfVamhOUa3/rOaw8r5uayWBk+yvF
NB5DV5jDUBZuDBwlIqkOEQ6sYVjaLI0TmOC8vnpyzd+uKsdPaQtWcLnlFKA7egf0
iCGJSO7eGdS4ZwE6j9FQ5zx6ocqVLK+7WEtIY7hbp2bXw2fJHXy7h/V01JHJTBzN
Qdq2TJ7O6fDR549Rycb9McmunkY8lu4g0X6k1AzbTLDpSIQ529DTVAlxKGPQTrvH
RrX/SUoYzApcJrVK/lU78sRsyKcGVP+eUpr6X6+vISXt3xPKzD7PQPWS3PkkQy3n
y/kEvlCdCvnWr9BG08bFhoQiO48/7UvJ4qYpV4++b15+j1BrYsUV/MDD4Pv13IyU
u1DCaZ1w8TawotgROBQyTz6QZXu04a1cpOX5f/fKacJH2VmKPsEsQO++CIb3J3Yw
jcGL49MR2fySI+UmO7tzxiSnhUkurVoSbIJReTnwp+nRrrUwzMij9FxrHcpFQe5a
UrmcDsxCbCoktge0LtQSXrURW8p0JEqXvlY7ad/jh5J5/kN6nf352IZfKSUlfB+O
66s1tw8L87KQPp/Oj9fM66IZLnkR8FI16jE+7mTW81GQGNPbOPxoF6RRxumST4rB
9y2jMRtmqeV3Y7SMYymmlvwTA21cWZVn8MiCvOwssXCoctXCFzvQ3UdAif6gI7WP
Mq7+iHNiGSHU1tzI9Ql7Jrx64tzK5qJKTRrrzdG40fA3lolZUejr/IgG5jYcD3cg
ngcN3tlo+OaaHAOtWUbyQBTk0O2hsxUcMce+QWM1VHuhPxMAHKKsikobDg9Zq8r8
gcRbwyfv4xzEUyib8jyScphioTjdBZlA7KZNuDeTNHq5B0RI1Jow8pBA2VdUUfgv
KeJo78Frg9QM3O+bdYCCt1U87x876AklMfzCmiib6vBmDzST1FF8B4X3TY2Rkd/H
i5mNz6v1ttNAK8bMrg1LWhGukQtoNscpK8p2qJSlki5FGKK+8qqgYa8zfrO6iXqg
u1OS30D02cd9iEXmu/KqzwiqlwTnZIfelw/zGxvErHn/NXpY/1X8iCprfp/rU5Tr
fTzf4qJ+fTxwzVbEIgRU8c94gaEy/8zeNyxxbpPaXl5owjJ8qxW4e6sWHVtQ+Aoo
Qu39Fkper92jwb5YPk5dSbNHlUqy2g13gPLMKdOgw57xRzBqbFFGtzVDUKFETO11
0ncLVicNNQN05uPmf5CF6mMIZ5CbQmwOVQcSvZNrG6nZHk508Th0kwP5XZKeE/S0
zQFTRtFUsh8n/DrE2ty5K4xTsDjooH4QrbHN1rqfLz7y6p619DOY5f78p+NDuadv
11LVAc3SqU83OW72jO7DFrcxBgsSHbvbsODvieoxAmRPR/mdU3AAfsMEgpmGU+yw
ZHIjnmOVKX7y1pUgMkLBn072cul21V1ymhi6DMBnAIXWJozwNOmIvXmwKccwVHZu
iGJcS/0GpTo/EYQOoOip0QvorZQwi35opl3Jf2HlTRG7IbFcQRS4JNuygvRgjs19
LNobJxYHDP27238AsalLvJ15m97SqO/pwR6kHbtIeRI8/U2Xau1kILsLWR2g1+/Y
rSIhEI8agEIGGQ7baAphjPM6sRdUSm0pXLk5R/R4StIoa5BJTSsQT3m9P+KgKHG0
BEEfpDWZDkdP3USiGMQYdc940EdIqYVTAD5dnyQUt8EjtvAeTH5X9MQ6g0uY5ucX
flNvdhDOAe+mPsIMBgZvSADpMQaPMhNfUq4BDfSdxJoaEkXmrSKMh1hpyZgi2293
2+u4FRVZINKp/OwyPOQcfKPtgFecE/P6JAamV2Oyk/oUe/AQIT4cAEkAGtlAiuxy
72YllI5ZC1YXqk/XOLZ6AL+MDLBqmgjHRiofof6MNeX3MZ6q1OnXpI1b5BAZp1YC
uubejzaeJ0Gep3BuWZXf+TeeD6gg+gHquJ0Hkag7HaNxyVwFN2TVDkVH+WzsifsI
JPZigR5A3UYO2GOvdK8VHH1AC2A5ewgCGOiAm/mqNBzehHpzcAJxLXjY/B28BwZc
ClQTI+ly9xhfJn5+jg2CgWIEm3RgTPRuKn79itsqinM5pNszEd3DNJzwyG/w9oQU
ZZzDTbwEEoZfrT7SzIuhfwsB/+LMRHXgJu4bMYIdz5rG1J8j52EB12pw9e1NZa7Y
PKqeZ1p8LD0tX/Ehk3Vfct3fUXFhU4krO8xfCXuDRS2NDRUzcrH9RzHf1A0rMwSw
PXCX3bLYsltPp3Hvv1uglJ+KMeRa7ljdyuR9d9gKnl+IgCD8KTp2RqtIozeX8f/l
cw5KUD62NylCvmsMU7z/kDFVcHkEt4f3Y1uyV7Y0Jk+reVkwWQsWjeYVLbbL2qgQ
wwNnydnSAc7XXK7/oVBFAxfieJ3uVHt54qaUFKEXLSYlO+oXxxa8H4sYmvjEGfxy
5np05LPDqIF8JulRSG0simlxqzklP8kf9X/elFBuyd2yFf+Wzv/s0+S2IwThAbRW
NzXDWqJ0tg6ko1rV/mymy6/Lzfly/2SJnhBsEudZsptoVEam3D/SoPtMNkBSk61b
/3y5TY0c3zJu4zRqeSQ6kNN7cmj5gd6NVuxffTPFxZCFsVAa7AjYGvxeUn89QlkC
8EKxnTELrIIIqQNGq0r+9tlK8WWCbOfQF+gMLcJrdpbrrqwdUSY1PoB50bmr9v4O
JvOs451SCD2I9OXdtg1IX3LyB8VOFJULS9qcTwBFnlRnmYdQ02wkxagHnIYNviBC
9WFffRPRE/EXzSc8d7NGXRXTkRGQ4WuVVN3XzgNYjNW0veo3stIZUFezba/gFwIq
D6OJJ0SnyWWVVZFsYQITINE6nQ+3NvdilDwSbaWaKPMJnespR7VTXe3mL8igE+fU
0z1ytL1ypIF/lE7rjQT4uLhPKoeg+F9SI5OQaw4CopUX/KWwSzGoieRfM2sy/1BZ
E6NZ4FO5z+Xpg/XDNSDNt5Yxg5rEJp8Orw90c8lQiQeDH5F1jznIVFylIgRxcIrH
5Jfwp1m9qTLFK+Jnuqi2TZRv1UD9WDTxCwUujGcP97yIM42fs9cE1KYjhdbMTLmp
qiz8ezJCPC7CQluSeQkQcTSSAt6FX6G4XcEhayfT3XzlOpeAGHElvh8p+MxlBHRn
CZEiiNGw5d/X23VlcEdwm8vQO6FxltYCDF1hmljhmi6argpI46BZB3m4IL4Rk0Ti
rU2Td0LAC2rs63XZm/QHYhPGj7mt01sHFYQlSLqvL3XG4diLpGTJIt1aahT2W6fA
3xG5Cevg94f4WxrnnfdhZoRSus+vxobFIkO2nQfMK6oLB1m/LVkooGb+sguth8fz
PyxTOHYLzDbN3ToBILGRtY909NAbRQkxZ2JW+NFpvbuxA+DxI1L3k/Zs7O9t649e
B9MoPIFDy/4PteB3coVgEs7dqbygO++WwPzrgx55EXIWJbCmO8+wFqZhHFFiGtvf
CMl2cJsOdw4HhC63NUNJG4wOPqDap0buIfSgj2nwmizwxP8CeUQvQYyXcYGx4BTP
hw6WEwpQqPNQmvrHTiOc15Gx691qET8BsQT6vbfmA7Uifzz7jGWHMuCjKkdXh+1E
wz784XYnTy9gbXMaN+yh/IbttBxD7c0/JBfM4c8MYgmiNpPzfwAwlntQDYn9ET1R
yElsiaEnfhSBEbBNMjNo5SoyMUvXeYURmWXN0pqXaYHp2PT4twMLJPvVV3j+oG3h
Ktmaagm67ccW+CE0Bw4HIAsm99BigpfKVXBtEqHg2CqWXhsGUTLtKBx/zmQrwwCx
xq/YFlLdayJvmgS2Zs0t0wxgv74UMygwRvRZKXR7hwhQ6U6kkS0vlSU2uVSNkAj8
iuKOM4JceVXhtVdSov5YvhYHcIpEtO71Ho6w9E9PGWZY8DMflxnOEqV8/sOdk8gE
VZq7Wt0p8Hb3wmD/LpjnGJ+NihRlmK4amxtjgltDEvXnXm1Te/55yvCbV902uusk
hfnx6yZGUDZEjFrcw9lyaO8hqhUrFRy7YzDSsR5CpMWYmPBlG5E7VbgZQqjLTPvu
yO6vyNcPuzN5WrjgtzmMucRRKcTdvvTtIlDy82feS/6l0fmSbAqtJcubrLkV0BEn
yNejI5MyLSuZpCxxXGNy0tTIVY7csd4NgdGH43xiTTQycCnxaMqav0oIW6JCX0HT
d5cnLh6/q/l14N2Q5yCmrkk9zEZAdRtL2B00E2IwmVoGjlrQDI6ICPe4Oew+QUHL
9G4kCAmj/m9EjElJ5TVM89501k/IEO2qYDStOio4ZXba4orcZOwm5M6seU8tn+Xy
t9+LobFg9p0xvpuDcnDbCggE6r7nbgVgGPGK1o+BdpLQ1MEnhuMtuEnQkIBDwfFI
KdKfGSyXkMnLBTaAOhLZZf81NmodbU+d2LBYRhA9KYXYVoX+SIEKHqq8n3f3hErD
r7cg80S0TgRs6Mgb3QRHgVP4KwYxn24gSnshyfrZlJIk8Rui+SJLwTBy2afqp9al
98Ydg7m/aqlZP1/6KvQRKOPPW98rRRcaUFy5yJAN0O1k7gPOBZDPt8jF8JIW2bZd
QDLQ3VRRSMdeRWIiPCaS51o9+4jqTplvnsbTN9XAfJmyd8NlbUtBSEJ6BGk+0lX2
ajy+aiF9bW/5t7pzb6fHud7IlPntAuy7x4dJhH2MNVHmGR8NAshsdfp7FHGuVf19
hcOFZZayba7qsSPljcMZ9KBedfDaqC8sCVpHNowdnrsB3ieYG0pNzKapi/a5IEJh
pXOpxdD8lG2Rue5ksRjrHszHrFXjXw3rbaD0c+mQ9hnk3gZrNtPUKHdfttBMZKN7
gspSKGucskwmuwMkbLwuKRGvZAJPVEXIn/t29mGpcI3wpMJaKgRmrFB1xsRPzQm/
GKpS9RpexCLDzom2gx1Xw5XZBxdJ1dKGWat4Sgce2ckICN0aICDxF5MwX1J/V8X2
Wa/HLrhooY3CzOEKgzynuemPWFdoCykrSaeWtxkKQuQUaqKA9GAjDPoMdYYyIvDb
uYigiQWSYfij79sy0Xs3GsLs2DQWuuc/beaeU4zGjfvuVL0hFxZdPJ/9MkS8qIkK
U1XCn5RnQuiPNs3XO2nDK0RRxF/q230IVEoifxdChDHsWDE01GsdVk/p1+1sOGNu
Iin+LIq5RNxtLNi96y7M2jW5ZxBHrtsqmDkWgx9F3iM0HvTDgq/MRJO/qh0Cvlu+
lD9s+sDkoKF3oYQkjB1ERbMviwrDTXkgjLvwHEDglhII4Tbj+x/wK0v2Ge5JkVKr
Fg98a3sUW3SD40XLCvfhLM3LfAc9mhbNmqImOuyKq3heTtPS3Fuqmz3taqRTyUuh
M0/FtWOzruJOGgiZ+C+YB+o/5/JZv7lDHG9N9V8m7IYWUjBI75Hh++OYWh9qhilk
KIk3P6RGng8bILfbbO6mKr9z9iOMox1bli9Wx7ePibzhlIsAxCvLXgjzG5mQBC5J
ZGizMSFQUou2a40WSjdovdsVoqd86rFP/j4Oe3BnnnxGf/TIAWYQjZx1wkd4a+1j
r78ppUjg6/6mW1QhFMqN1kgYYSchiMiQaJcaCFmmgYJpZvplkkFywHIENsLr73Yx
caKesSd1ubpcKqDbN0ND7yjJQVdKjeLZz/QiG4ixaa+HCJA8gOKWsQgJ1NeI/9op
uBROo7/YC6x0HYgnXP6kui6x+DxFAQX5KRu4vPPVZN1fbdBTjZqh4mSo+h1reUTZ
7V0iql6t9e83tl9k/FNyo10j0AbRTqeCxvOd7HI/1j8Mcw0ny7GU8SLSkxO2rPDb
JAKLpBAQNMj6I/omyN0x0nlrh+8YONCLcFnh9hfFC+WLIWUL8MotPR1M8Y0vxwi9
gYnWSe0Li097HPcfgAkNrl5q36hBtOXaOFuT3JU+O6ayBFIJ+VO6573L64vBs2UD
FYWFvzLd1wmCvwliaQ/uFOLP5SWk4c7CZZO+IrzS43ZQzg3aPRfu7BTmn/gfA3Vl
7opL+D1QPm3nbfYRVOW8aLyM8wH8WVM436BA0LWali/uJunRnwcwzYxk6B6BHpNV
nRp8P7rB3MDMSb2RhxIEe4eccPjuEc61QqjA119Mw0HfFlkV1MAREBvkYqs3Yz+X
77YjiznmmhGbhnrpoRnBpQ278RQJDffFRbpiIGed1XWmJFPApdQrtIDiTlXsefB1
fNNTjncNeqasRVV8YFOE83QvRYQiu/75qJU/0LzfMQAaNqJryEKdW5Z6sY3kS2oO
E1DuvpJX7rtyYNtxnB/drdAi265JeHjCyMUznx+aXXwgPzcn7FAddQPufGneRyuB
43isO9bKemJHy3jFnN4UCp2LEPNnZFONRX3NmCpAnISUynKq5vDlRpP8bCNs+XGH
RKAzN0xyokxnoD0TYJcAmtFc3UTFGZUzZrFiVXNW3mdbp87GID/PDKwEdZdz0IFL
onUF5S0HtqkX/LXSb0lMeRJiFaPZlLGazeLR8FsfHBLu9/p3hkUNXZR30xOSlfFQ
go1Eagj4PI7+ydyd0gZeELBz/7tGZ1UV+Yv7Dnf6H/xZzVXYK5kOEZsKWHl59pPm
SD36fgnhuKNyKMQs51+QBLlglEcF8KVM00uhF0kIk7NG14hgv2gQbMkg0qOl6m+x
1oBkCmuNi9vC82cxEQ9d2Ple1Eo5wzTZg3zEY95J0Y3m1DkpYHOQVnFCzpx3Z2tZ
JPek4Nbt8iiHOjyYbGMsR3gI/Qs/3Lx574SZAmTZAIB0eRwbsRNqX5aGzM+BSBQx
pK6uXGnaqGIQKg2lcGmhwjIR9Qap6yCMW/LBTvGLcrZuawjmz5yekKgJpc92lzY8
+3W8iH8cevD1UET0h8NVBKkqS9wWEe+/yZREPuQMde7qmvHqfvcuEIHrbpfsbvxD
nLtHkCSPG43PaSlH+SD1AYIsCqq5n0FMGXor0sz9ZXFRfDno+1cgVoI3H65nu6MN
M8MTTPRAPAhIFK8IRjOqVzX5dg7Fa3sOyIOEkSPuuo7pC0N6e33bueMPRhMW9Fcl
p1C9KghCCbq9Ri7hMfF13yoQWGRfVEF4j1V4xL6trKEDka0I1hhRT4FBWuafvWP2
vMQ4Y043ZZ4SF9L0TXk9iRBvXJaQv+OSkiLD0BilttfBn+fuE98qUWIk5Knj+7n4
TjbSO9tl4fVmp+V3g4GolxE4eha382e0DYuLEo+mdIBk8sdZZJ0iCPveUFAcMD3m
RIV2XKeBJqousslVQaqOkiMTCJ4k3Hwship2SR7sqyKENRIuWjJaK3j3o8UV96YM
VjOO+XlrMdFn/J4kIzThHG2c5VXHFYr+BK/JtyhC13ZFsdJSiMtAHnZ/iueEMHoo
GJo42VX/qVA4gD0JexNvPzvnwLp6Xl06sD8SOvzfLBZ+orZuv+czNzp1bC9LfnW8
hlB/Cp2MKUtj6DQ7TKXK4ZBngxGX7J7ct9QOEi+Xl4jt80qOHUhftQhLkp8YU5FZ
CShhf6er2h5ZAo6cJG8wN4Td2sZW6/teqJ1w+gRFjikEFv7mQj9PmZ32l1K22B1G
hQVP+wc0nYu/HZh8A9ueLvkm6T98hyEoWJp4EUxaawmxJLm823zOitzcjWjcFB0l
JwmaRb5tT6YkyAl4qbGdwUljd2C+XnS1zXyJipTOETBP5PH0nEdvonoT6wmHcyB5
rFb67KsXvKGO7FpkG1YEec7YK6yNfupylEdcSLV5b4zcqtZQnpKsPA50kXTSD8qE
qIysLPvJRzqaW59hi9CrKMyvH0XwLro9keylovdWMoF4MkS6QmihL3JL31k5i7vI
qsGvrnsQKFYQP8094GgFi3uccinqy6EZ6qo1LmzkUj7KU7iTlnsYZdYrouI/EtMX
Bk7hi46rL4HV39UY8WdWCDlcRL2K6gsAC25SbUVWVPUyzG0kDlTPngCa3IS+5W5O
pzRQ3WehpHLBnsC5hg7n+1YVNcLEOVQn+YoyT0bMc0gn/1hK8C4hPL5IcqGrrQlj
+OPRYSkCKLK105mp3IVpAc7DJ3kbo/ZGP5ueIp778tfXKa04TnN1zROQadHjDbex
cC5hhMgERdtwbG7WiNOo4IQLFD2vzQon7lXIw4MIeihZ7iSHkKkhZgbTyu63CbQW
tpLj3fr5mdmVRtLX1+u0+OPVIUjBP2aWhXc+EkNQ+BQdbMTfd3Q53ZV95ztey8RF
X8LbO1OL8uTGhpDi2a9dBfEThjhh6mXc9m8QxBfmFqWFB66zq9CkOtszI/MTj4gx
RU5Nb/HiOFDVQ7nx70xIE0zGGTT7u0gyv5O3URlkbx7T1lsa5mp7GISlaeD14L/f
1ZGhvvzzlRIFctGfCt6rEQgY/lv9bBN3MSpZZmraqWlbvWN/EH8w45gdeL73k+Ow
9ii1Mxo649SMSIbe2hfjLeimajzLorQ6j0bzfGXVwloaLaKhoKP2Cei9yOVpS1Pq
hpg5Ap8j7vogSg7WQMZIp3CNo7EKyzAP1Qhb38kW7pkglJTJcdfabdJFnShmDoZD
uCbNKhgD54+1uMYyNCVkIt68mJF4NemIlWqm3Gi70FjzMLDrifW0pq+Dqs3iknSn
ci6ZvXG9opTiScZ10SGZX5YZrtbTli2nMIKHXLixMhd1yBYu+hlDEH8nq0M3k5EY
4RPZU8oRdKWTIdDZNQkUeK/Q7fVCSlnV1IA1pfj1udPul7vG3hSdtKeBxtOwiftZ
Q2z+74i12VHHWZDw+/541fu83/95ZLVH+aNdklvvnFZl9+RWLjX7dvD/vN6IAxkP
2a7SbFWzQ9aaQTlo56uzOLXlEEEQqQ1tqAGI+EdNl5ZOCfgBqsJrpP85EWcgk8PB
5O7Bq0aI01PKX/ceoencdYpv9mhuXl1MBL3J8EZ4YM/Rf0d97Hay7tR8dk1G8A4j
vDIawlvBaPO3lG/AFI4JVKQh2lcAbABieFuUi+M8m7Ma1ZzJEjSWPXywOasFABWT
Uv/V3Nh6hv4BpHdFXE6ZSjPe6fdvlxA4WTWMwxExUrqXwLcRruUb5+TWNA/h+4J6
EIozHPzga+GzRRkLevRKM4AFmght9iHXN8MPwRs57Z8DqlqZk00GZPMogBeQ7DIA
4pWbjxk90Ou20jRGyFE/cexzcGplTUNCJMJHUkesUqJf/rTZszqDiUM1TopmHGYA
unMWL8shsi9nRhhKWwUqvq2KyJYHJvkRy9KRjchm0/58zE55yB8mXdEN5bZPvv39
gfGXxoQ9U9U7iqJL/0/ymD1WLyckRLRhZuysaWsCLoQmh/VjOPYNsAlJ23G4JWC+
cmNBdr7ONbCrcgPgaAtdzje/abL/ttvNVZDnRSqmmcXRJ9Clnqae8Fm2dqfaL16d
ovVs9LWXpvBFuP/8W2P5TOpHM/bzZgt7/jYFyovpp77PLkKbfPCkIfZgjE8wDieN
/mR7vPeU7+uXHgSdkSqvQzPW4iDSND9Am2WTfq0U5XWXyG+Nt1YPPtiOnC4alePX
FGrfA8bAQ2gvhEcZu4JFOENW3V1luVCS3Dpj2owhFHBEtxIj2WPR7At8yPdyl/Jl
+T38Actlk8BRbLGndAKJCf/wkTtCiA2VLycZHHkBnDI39RKN+BlB/USEuD1Gqq1B
0ZEvpBapcH4C825XsKaHwqxqqtWheaz51BbHLRhKsqtvBTenhwA9+Wi3cYTwvy2i
hQ6l2yQfk4kb35+Umiu1GnS6rHSfsCiKBvIuFFkM7U23RIszda2dO2Ikn5TggjXs
eUfL9WpGcAiRjMcgRWvyE1mwn85/Tx+1N/puO2RlCEJ7a183p9x4S8YM4MtA7YKz
vM5v6xU2vsrOTR5mNo3dRC5ltx9spynr1L8Oio6VJKVfKL6HhS/2ZSzoWAVt0xdc
7toAx4UE2Rq/kAb3eFRVmjpNSdceKvFatJZOjlaFI0xL5ZkoE4usW7iHVUyqZ0I5
xh9DJSFGG7FcmLGr6eGxQTUpYMwFkBmxvLrZO5vz6+397uYKDXhGzODhwpCbnACn
IS3Yjwz9SrM7NeHHomQDIRPwemhrxGBwuweW+u4s02whA/3S4/TI8LGPRUmgnjP4
njzRKH02QpoXIYliv4cUTx4J+DlmjFKZs8w7xdxAYaMIcywsY66OW4sS0dQ82OVa
ZZCF4s3bhEIz/aDe7/wm4w5dePdRydhRDbgJ1emLZ3ieaJtdR0Ik5rg0Kj6WqtxP
6163Pyy3Gea+0ik3APq7yGIwIzIAVa13Sm0rsMWJmYTo/uNolO/dUDKPJurccXT5
vUIV7KwPDnq6frqMxmxsvEtjXMKTfVI8DuOIXoDvW/r37SWpV2kDU4f1niY2S8fw
YcOypy0kmaVJEqtnbjJKgZWgvX5pTL9tF5yYRblH0rRd89ebr7dxAuZmJQN6srfN
V9H73VTLFifIbfSo5vviB7DKV67JTK1zgRce+/5lMBq/p4cJU8y5hegdlgJe/F5x
XgasgE+yu+uk9LzfJ25O1i4LbsWOCvGloSLZDIiRfjpk/Wm/ytYbng5UkrjVsUhN
DHovDMozvebennEUnJWB4YCrsfKJbRXlILP3ATyzQOyEyocQo39wVi0AiAPUyRAc
pso1WpZNTw4gj69o8dJGJYvxuYuJmz7bKWxfbnLCRae4ZsPHwUyJQ+ioIVFKtJVp
fqZUcWGTLO+nwHY6di/dINwNJBbyXaUxrVmZdCsYDhnNXmsEOFZg40FJLEUtnREf
J1yLETljHqOkYLCnTaszrLOKmKMxst4XcEHAL/7Q7UuysZiDYaQ/0nu8lBhroUbj
ftulcXpNzmzTEdAz2c2WB5net3ZAE9LBTQOonN22RZDAGsO9UlRRehMY+tpKH2B2
2yYSFkLrfOoh+VN+6Hcd4vZpAq1jQr2u79MdkDt0uIexXifwAWJoynBftriugMza
DaCxGZbrpr2F2OuwdagH1VFYhzbdYmaU8XMAmCBJA/fWwFll9Gn6cTRhV3s6fDSf
k+Zk3UvAOfyGIQ1d2HGltJvmmhhaJtEOVE+AMBZFD34XueSrssgOLADM8SK/scBt
gMmB8CAw3JgcuqW/KT1yV28Gx6rMZAmt78lROteK7GPvJfJV4GO9TPD5x6alFP/T
FJi1VgfBhMKxZvtE9xm0AiDNYFA++Df1W1aXFddfWCBLS1loLIOWS4P90eJjAvMt
sJdeEwGJefkVLqna8uu21zWq3om6qml6tDlXDjwztAmlTlE5VbOupk9TtwVQpuPU
6gmm4ZkeZIDRmsOX9Luk2DhM4Dy8ZMvLtwwB0XRDAklATBj3YmZs83L+ZpNxklDt
3VvXncyxJaqCJPttL+TYnQq3cLAOBRq/ys3ZF6jzVBKWE4zbnGX+10IVe0S0YfhB
H1FF9HuF38H+OMn2Kr1L2iHa5GTu3a0q8vrQLoy+XngaoaJ8wTMQh/PSGd41+vF7
RZffP/XLRxZ9buA9dPGMNXvFnq5tjp2rUJILoCPSA09cmar7mR3qlV2URnP++F6I
VWoeyImjpy57Jv60sVU4dqoyxBNhK2CaOVzsrOlLBuV4JzTlbvpQSvXHge8VnM4f
gfbHLMDjhr5v4o5xhy9twrewGmlbM6WZ0gJ6TW3EbHGlDVnC1D6mrywkAoWCOPVr
2vdZAEAuLWAWizPzO7MeYbVuYYZY76C3JtlVHYB83eAQqEc+fWBUrUknDllJVFV/
BW5DWCCFwBn/yULNVlaBHIM75iHjx8Fy4YFVQTmy6TJ6A7Bae2KiUuGyfTvrfKAZ
buFEz/cnclIoB15cnk4iRXEhXoT3bXL+Kkj6auZ7ov6ksaUkUSWTxCJDiF61ceQi
qeKLjMVL/jIYoq/9ZK11DxvyvTqIY0OvI07gWRP2zF9sp8tvKoWX9sqLPoiMdCZL
1EuiBYhR24JofuZ2/UyTmSt0nun2yeYvYPqTG72Q++OirFJmKlwgcNT8nTuWjlkL
T+MguzuZCwaA0B+dotdxCuHumpc4OZN4zkNF1rhggmtJ+at65rrSiVHBVae3UCHm
u5/HhX+dVbneNoAtDOhAZGg1oVQ0NJo/JuoktdlFr6Kxx+aMkQnQD0XL2pXJpTlK
DdMpPp57CWr0Al92Vv2g4JwM5WPspwgpnCpr6BoCQ27ekkvamW+d0jhgYe/eqHhM
rWftCYBKwmDpHfAQI/RsBJyOZ9m/azr5mui2WxmVuvQD5zRFF/eY0VoarGFkAAVZ
ZDeQy10jghX6eNltFks5sKr7vkiTgb8OaoCGNo8Vx3ovDGm8iUBm5teGbPbQ9vEu
px63DRohFGlPUrIH40Twas0cdPg5Oj2Wm+WUWiBkgDI9kt0y1TegNKqwv8uTOrNE
S+FpTeAR5LiFR6enqC365WNckM62GJTfvs2L0CXWkyQ2rVwZcv3I9/tVQGAVNpF5
pOPAoFUTAYZ4Ct1/VbDzyGsVKq332XsTs+4SqZJ4Y6SZ4lWGCqgaXcgcBuLcd3/I
gBPROc6G5nr7HVsE5LdITgRnD9+vJcUAc8LOYHRfjGi46eGThlZhYTv5b7a+MtMf
G0UJfaWH67vhWAKeeuUF6gKBrOFwHLkNKFNeSzfS41ymxuiCCLr/XEjdfs/YtNLL
hT5i9Ch/Jl2gkYggUo6bXjN1ig64DTC4B/OV2r8BTJX2T53p0TSWZSIkDUrIWlN+
OWVwCIFxrLaXWxv3gZ6RcHP2M0m5IT4rJuj5j4RnaWU6ZReKmIZjNvcOcm1jeYGk
Om0bhiWymw9w9Tce89z4TJAPcrHBaNOPC+7CHGCXo+rT9a9okbz/OCuNCymvmjRl
WUf0VxxJWXp/5BBoU1TR4y3e94b5RKeRpkpTlG3VbaOV3JqXnm0/4Y3EfpzSKrF2
BnI+pHpQQ8A/GWZwDCIVfN5a0cpDaVA1xUGZMCRWzGH0Wpi8X6peOHhI8Zh91WsO
1bfEvPF5/OkZuce/Gj++AJJc0YYfnkwA41K1AbEn4ogOTzBH+oXgfowBxhTDLRZf
gtHf7SIbZ4/3Pct1QQoeRaa9P48oAYwB8XX0dkkp/P+TKVazTb0qpMrlcrmwvyzS
ObKS+ICiPaYcuA1n+oXd3uozY/NgSJNrR/Cz7VouvZ2XSNVzrZePJtHrTRJGE4do
fjGoTcY0PiidRyQOKUk33rE7Nq9hsZZdw1XIfuU2SPqZsaC538LZCHp/uXuUv/wC
sR0pzX6lWq5n1PncZjcqSeAmAAl0ft1DvfceyQ5SbxbcfO4rpcndMAfV5O3RGb1u
vQPb7CikjkPFz+Nn4rnCqqfT1C56SreTLnrg3o+Lcm38ctjK8JxF4cB2XmKx/jyC
IMOR8pcEjir0UEvqmBWgG73Yoc0alAsuM4/thx35KglOggPYJnTmuNTI/Mh8FKRD
UDPf+p7MA/9qRqnxAS/XpgWKGoZsl98yJWB4zfLkpPEbPL0w5tA9Ugl82P98wRGJ
DXCA7NiKlPwC/Ngfl7QksH61sUjQfHbDXf86xafnoaloewhoCESOOcJxoUo8TzRt
TtslcCz3p9Tj4kcYqsktJLITbSze3D3jQqeumGCr4HENOUVxa30T18CZv2YmaIbj
fMYiyplMagte57EA9dCUqIlLjsdCCy0h93jhRFxPyZpQ6ykHknQqIYTzeX2aV2ho
D2Ymj3f+h6oSB2e/phXIUPBv/37Ow9V5fVK/v2qfXtzPGDRbTirNSqY81z6mN/VA
nOcg3Qgv2FFL3EYyO49igHhJfrPBGBHFHf+xNKW+5NkCq83tfJUwN7cCuIdrTIHd
UG417yzEm11kRueXL3h+Wbb7/mRfFdliS5DVNvLR3ZmM5RhRw6B1J34K1aU3Ykuc
dcaXcFKB7x8wS5bds3hk4gZ+RWkds8b+Bnz4bMrgAaMrLpwGFWDh7aNNLKmZNWDN
n6K0hUxonSJ60Go2dODLEGu/G9rYDYPaSQ1dozpD6F/5ZHljcOk+/LV8Wg3NBoWt
wy8bN5VzhQI2hkvc0ej+mn8oahKPA2DGrkHsmNApXmPMTCpf/9XkofpItDP3kwZL
NPeJtlAkkTfMS1fpoJNcoHWIMOaJkgeMKRbJcoP8fGXsZL1gFvrWYeYC63er7/E8
P7QzNS1/zS7/zuv25KPoUn6fSUO42B6ALFSIGRTTRccPjCbCdjo2hgDIPFLHhw6p
ppqHLGqocC7AERh3FwXeQCjqtCLEktJ9r5I+CoyuNOaULJ3suduc803rnH3lTVUi
8IbzmS5ReQHh1nlJqcbdY06Q7qNjJ7djY+IdPr/NYEiV+cr7cyx2H9GG2RvsA+sY
igx2Gb3DIpK7HpevxJimEyexZVfeOSdViG0BwYrwCO1LbuEGLDpigXUol5+1RkRj
vchYE+CeK5hMhchCASb/jIQu49su6IF+GlGUUW3v5AQJ0RClOfEh9gcAam/b7xlH
Qjw6PDcxHRi9+Y/rRmdgSNOhRaj+zUD5iOMZEF0z1lnsu1yeH8Er7QttVFGH7Fl1
BNY5D480tXJE/4PHRIwrOWiouMnunGozByWcYm5/0kZjhFDVBY3QUcb64VvM+a2I
lD6uCCcqJ1PI6J0sDPhDnXwd0joMxFDHirguIZPEXVlyAuCi3myoKKMWelOTrkjn
WZt7GLIbsgYqcx5ZoRSQujP9YJMRtZAMPWpYARstiZkQxohhXgI+O6my3KzmZoEd
4YVrxhZ2fD7+kdmFxbu97y2ZaVhD4xttoiW+Hd/d/HGaLExjaCCkJWQfm/gD17gF
/Fidd0ZbFeJP42/Mq+4gYJh4StEshzdCqWevixB0zlO+oqoqi47f/bsuRgCqKEBZ
99Ka229cVdm2fAiYPqf/+14JaUPjU1+Bo3vaMItUvKt3sfG98udfKtCeOQ/d6xEq
o6MYzJ/88LFQq6923FWVA6wmbRd6iKUtWowVK6mX6oy+D/1JaYiTMoSqRglSbe5s
BYrBUrAmAAn3H8WAvEsm+F9nx1UVNWt8UC7VHWLGNthEb9lsGpM95bigixxKTE9H
D3kejl80P6x5Rehd+bGf1g86hIZLF46EsYjd4Ax1O/1upfTVMCAkKQB0g9gjzznD
BztHWumgWJmNtYfK4eNS/gzzwTdQDINmp9jCDh01q4mZo09MsJMKb1yRBEmbcj3l
KPoZDOxLPq5jLFZwaZtrIPySbmrM1hYBkcRyIC4W/NhnoTQBxIfcfawftX4GHTIz
G5S339kDhZ4VJSLBmFvNYl+eh9Mrdsqu7reGKE6Ot9vQwIccMc+HbL9Xu78Pe2/8
2ywyNZEJh1QmlXhc2M5u+qVXofsat+xflzd5gpqjPthrPp9SVY61thHU3cX5UPsM
a3H1m4LUcyUnvADQt1Oj8WotgruIO9GIKBWsHVWdm2obkJCvRrrAdX7OhwKvJQkD
EUcXDVcutsxqK32rP58rceVIEEB0CkD21OWV4iQneYTEhfAHtbNkRwAyHeClOfh0
FkJ7C7LMVAGmA3UVVKjdHyQZUF6hAOfXO8MBvHjscQM2S5yYDe4hK1fpbJ3vfhOV
KihJo+lQGBSOZc5U1tAhta3EcsOa3+aRcYhmpDcSHRKdJrHzKBRQVRl8JF0ASOZl
eYdcYNucRdjymP7wA2NCWoArq/c04QEfEq0/WAfaGHmCw59P22U+HnJiWN8/oHKN
zPaIPAygXu4kM/iWTZCSIpVMHfi7XT2mKQ7trnrdotYhUjnsuwACw3+N8++cfvAK
Jbb01RLTLIruJpznX5UveoUtQzRnp1/czfqVg9INirEYDMqiIdRwRhLkL7kIwb3j
W/5CkZpUDywOcy4Q14QBZxaSy/j+0zGEHZDOiiroEeUgZJBgk28dn71kpvdjdzqs
9fbyOUqTMGOrOMi9CEZjq9j0AvXz+q7cERPyrOVp/6t4qh492Zdhyog3SQ4pF3rD
qKjn6vxdFhVhYW8pzKlZwaUmCgZyVJK48Esae+IGHRlEQFoqJ870bYGjuwB2jQ6f
pTmidMqWVrz3ljg/HnXTyQYYRyiPbcNfjBTGWmd5i6Gj5RlZWwOmkaa8114Ufe1P
FPVGTcgdz+M9ADJxy5VMyw/RHm2nIhhG/mz/A7b7q7sULri123vhAMJi8ZEPOrCy
ir1NwhQ3sEOF44XK6a5Ay1WPcDtonxLc2A7I+rmRNFeQ/iGXB0Qjv+uh+GSeRGP+
qd5X95Bi7t/puYiveeBIyySDYkOwEbHnew0DlYpp4E99GCVTJJhSsNBPGs1bJXFm
QmrDxx8vJX+/f3ptRbGwRyZXWAMYkJaAXQqjFDh+fVWNFZ3Re5M8+lSr9O8ZnSuu
BNOzMZB32ncqt8NV4JnKaOMPhguFKLyBrTod6jc+FVuezM75kGBFmeVdpC2XZkS/
zmbGuDAwMFB+9rufDEY61wA5cRihg48UEkNnmVtv9IZjCjVLR7MnYc6h0D8jyEZS
zpr8/4PyM5ARSAQu6Vg93CVhfb8j+Pg9l7M8RiVgFekNapYfpgtig0vIG98+DFJZ
dFus8TE66a1aupHxNV/kCELApufaN7euvIDagWT00vjWw3uSe+hOWaKfyKxnq8M5
7cqxoB3G3MgZlVGLM7O8ixUZn0xvEFQsLWOXzrejkGsF7dqj13ICd2Hhp2/bN4wy
yzcV1pdkEGe7qOmyZhPd5fzgWVTYODhiLDU51HdakpuHypwlG1+MptesUJg/q6ie
4KKdtiy0xgNOuUggB+NdmfD9O5rAycQ/Yh597yf/snOGSWZ8SZWvBi8zK3IQ5Vnt
kHd5MJV/EeOoF2QfLJi/JlhtsTqEGdrmL9zhI2h5Ca2oJx3AoRa+KtSp/xId+EVq
QEzoidMEp1kLOfzUhfGoNErwiVhqul9Q3mNRPLbLZjpu+VDXv7fJmyhLjMpPkjoA
vKTn242683B9d6dzjeiSFFXLJk/yIFxj+ogiLVzAF4GKjd9tcU77Y0SjOABjRfIW
aSTXuAJxg8Fa71IKciW+0s4cj3Vqq9rdv2zyl1YVXW/dNb4Jmqh45NHFptmWBU2v
GLbDXBXzXMenw7Lr3J6HxacyeX8uHrF3HhMxjLO4aVhAxcdWD4J0hupkh1McA3KW
NQ7P8B/AtO9I6oTvIJhgEIXv9ehCkU4wMHkVVqUdkLESWUrJ2uWp9jggcvU/d7Wk
KffHLdh+CpVpTdDYYKJY7ti3qsBVL7lmibCGL/tnqby9lxlHCBcn3SZerNQwTQsO
l8urYh+saW7/pm1zxVofPszX8cQIWZuQqdQirZ82/oSjjboBW/TDcofRXaKfHbAE
sIeMWQHf6r4Wi9hcPBuAd+yXuHh9BhJ24VXeTZx+ozmed24CQDTVp45sZNimMUzo
w+LV+26F99VCnBB3byq82rDsOAg86hV1xS7mKCfpjGobBFCihaseN3CVS/JEzh5j
V3ccYRp7fzCXCQHzemolf4zMoo/k5aJ65Gv3Unffsl8ORSzRkPUXs9b0m/ORbsZf
4IOm5Iix1/B40JPpM8HYfTYIfWfDTz5/FySykq9jPK0IGzcojeomCjgcJOpkdqxa
GuIUFVzhjS0WQXvDdN4WxlU9/R93Y8wI5VDNYBVC4oENOvuQ0/Ly3ERnyrTpy7eL
sZcbN8V1lDo5jqjnO3ae/v3nX20R/XslE7H9rUy33hCEPfczeaN99j01yoSCV7bg
QpJ6mEDOa4EOJPZf6QLp2t3d7TC8TyLxu/+OmgmrOxK1Oxily2l3/ptvFvyROSsc
R5q4zzUOpCGRkF3eisdAm5l7jUr6k/Ufd5/mFEz+BU+ePDrkSJ0hExB3v6OJJZ0h
o7TAAQ0rmIMz61IZhk6vh/gGKwuHqzNWCeQEPL2kfWpo526TFCkb9i2a5LrVkZTl
GDylbshctzXmnckqrnH8BtRObyhcHlSQklkvmOhhyNhCPacBRD/X9QODl4lH4Zup
bXmGEqdq/l4SxN7h3zJbPyh6KSiOVHZn4ItrSbYp56c6CHTVxv8B2gxawyLSWY/I
`protect END_PROTECTED
