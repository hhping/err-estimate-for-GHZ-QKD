`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/Gw7HRq2UgjqjcURHea6BQ9+SXA5LS48ithuTRPoONCIS9GE6XkffUNaTKiliL2
VjOBFS6S0UoBSgyLqkNatwg7lFOsiszFq99/WcM2lq6MsDCtUZ6VCWhmX0MsNhj1
QX5qTHqiIofq2Zr8as2Jrm90w0wudegwbaxYlaGjF9QCayFOf5hH/9k2b4r21Li0
TbPvqBqK5YErMW0IYelKH9fzXM94JygxE/7oaj2fTqelj+YnLEuG6uIiN8oXWpf1
81tbAPu3+kyQ++Xau68874LIj1oOEerS1gyIIjyUyj8hBpW04SmE8cWTSSV4FlKl
TQLzOQo84UytiVIbEH35Ws3KGXXJkOGKnwv6qfeUwusFeasG2QyqPwfS8bi5nX3u
VU4lXl6VSCWXHZAZNWw4cBjGqW0+kmhDLUekgnB7lcVI4y8Q+LSY6ooKQ5wte713
CyU/644b0+UAuAhDvoM1nAjaiTHizuEefyfwVdX2358=
`protect END_PROTECTED
