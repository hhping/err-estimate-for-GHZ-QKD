`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hishkFR0IPxQmRzALGr7NvvurCpvhL8WaKrrie9v76xXH6WNzlUxXeSbeDjrjQ0e
RN1B2JpluQsIxWHkwTlqhuHDvYSu6vbWGNIsXj+m9BcH0sD/rykUC6YWo/bCx6KA
LRzqQ653Zp+HIh0jh9lJxhC6Eh6ItVM5clfeShR+CK2KIui706aoqzKr3OZRcfSG
8FfkmF0xnMg13dVBgyo4S8lu5NjFoLZBR2RFDi1DCmxvbhXLh+pVwn0M0UVimIDC
n4CcLXLTRZm8x0le9WUBYYKQ8QcVgX5I65dNQT+u1n8xwFVFRzXRAni3crfNi5W4
Q+FvWCsSpvMVovXti2yGnpgBNi01As0m3kFg+sFrxnFhM8jFNEFpOKzWYANfoPk+
O8QNuT1yM5CXJJHH7Sg8J4UVTGnUWYQgzN2vyFrRVgzVvl/WMtVBTFCcCycyC6WB
vYAGDXlUD1oGwFLz2SbQUCXjKVfiD5K7X29nI172Q4wBdA3aRD5suKDJJHkJjKhM
vn7GDYWTFDDh6CEkw32k3hr/2ywLTN+JxyDYH4eBVHL71ce0wqZgoIRbUdvuMk+U
fsObRRyKeVrWyaV8k8uUr3Gzqz0bWU0kmmu2i0vYJzUKoiUthUJ7Wva0Sk5QVzIj
GsgEOQ0AXei7OTOveRyiDOOrIJRKuYd7q9X63G5/Rl9bqP8omTgdN3W93Ctqu5bt
+K8oQa3mzytY2sYW75bW4Ams7XDWav4yVmQrk90skVeBup/vlafJyhhWGC2i8n7U
RA0Zd0hid99DrUyT/2EX1+rLWqQA3SHReS8jlVvn+eHeWF6Gt2Rf7zpxuOF+7/Hv
IBwTVB4zEAvPRVw42YX07tuz0XnB5NUxKO6qM5/bFGs1azmVIWBlhGyHYHpL0L8t
r9byebHQFN11raVVzxlCJTPfh6HCuEE6WHgwyf3r6vyiDXaprsrsdGRo6O/ARUPe
VIAAbWOCA4PPHJHFf8jJAmM2pz/bLFg1o8t57vn7/ycPs5quYyCagVUTbYusC0bx
XAJJXFE6wY9O0EYfb6jnr4VsnbmA+wLOft3Jn2f4+PY0kY2ZEtt8Xr7iFlrE9Yk5
K3lsKc8Hj/9iS/e81KjNPocCGVbguCvBUiPgh2M0q6yhI8JTxKtjOPWqrPjLD+A/
2DwveexLlZlTcuxk9uJL4bX+da6aEQXz/4kq49mefPEgKRwSoH6DWfZgRDjbmm/z
t2g9FBC8DOfjDfNv4AhwvLCpE7gz0lLYITv4SF6xYmufUeEUI8FrzIG8o8ViEe7S
49XvOM+cKMAxIsFPNdijlrcMxU3Ywvqi7papS9jOXYGyeGt+Tnl1xgt4O7GVCFEb
ZmFPPe63YUi6Z0tYxoePiqFc5QSBgteBeH/QXCPUNpS2lv23kQw2cIcpG7HytP28
37thQGGOUmUeytUFLO0DWxJdhzDj0OBIcSBTFtxHU2QezzuakFQm/4ORaKQZwaZL
7tRxNd7TjTnEM0mxIITKZ5tkdrvqWvX4KRGVBO9mp8dqlnZ3gYeM1khahegA7WHO
JZSL0gaBHjTCSgJRre/HLjLsBnp6GSwTs/lZug2hJuYtfqrd+Ipo22X+UGbYAC47
adguZYWofoSk6gQwO8ooFCwS8c/Gd0FezB9HwbICrbvMLHxjO5/0EidPfteb7lo3
83wU2DCpr5Z1RZVnO45RoFAFQYGJz47THAvtmvdbzxuhv+XWq1VpPESkBkibcFGT
2CafYJ8yVhghMeauUrsuLd8m9OpcCVL6/ssfY62mf8pMYIjWtjzzl7/qfw7IE3D/
tGZK+k2wbgm7pFqIk45S9WyE+OGKLfWGzEQbwvEC5Cng4yAHIQw/bRRSKP3EXwwO
QcxT7x5c4+7a7pzVRUcZ0NKXNR1IIjH33IOtZC3V69Hl9aiH5GU+g88amwiYqS3i
29a62r88tqVLdQTuZqueJjcnfxIvyKYcGcLYx+wFfVC5FW7rhUqyr2tvqs3/y1aC
FwGHbsn0GZmvJcx3E4OZ4a9RRXkaC6lUhdyiRly+RnbfeTN9LU/ywYC+C4Ose4sT
zxKpnjzY7KsuNSrSOWsrfDuvT/CG5vtyM4uDXsqvIaRP7WUOHHjVkFyFXgEdMRwF
eCO2ZA00mRSxNFShak8st505e1ALHTkOSXCs2FgMZKsFGu76g1Cs92v6Obw1oe2O
giyBvv19tC6i1Ly4bMgv07Nmu6G4gL+//3QrbwCtFtBWHBo7Qi4FOjBJdVYGJnTs
XSe7VpzF1YWAoKsVQEeeSL99cSj9xGDnItc7i5P5O7nIBkv8hqkUpkL2VhuaBYM3
838GhyE4CK+qt5eONCy8p5yljc+RpA2ZL3vKURsfs3fgOwON0a+AU1VmTvzhkXl2
CK8x0uv182dOvxqtKSJEPQS0rYvoP/K/2I+FFZxmqhpecEVPh1COKHW0Jhf0L75A
6bFX9Aa/ku94z17umW7i+mfftXPMF5fZrLDLzRBVPMOYDP9I7ilVuAIuG/L9JZFZ
5olvLBDEfazDoBCvEJzI7HT8vOpNAsEg2qFL/kAi0SD8sTo/CPZEOdAYJVGknfDg
2XeW0RtNXeGuRxndcSffnu9zZcasIsLQ6LjkPpX1EHxS+/ZwOOO6xxNMFdygmM2C
6vQM8/4iHPyjn7tUepkxTiExcxs1qglN6G3Xu9hAYJU=
`protect END_PROTECTED
