`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXh9anTizib7cjq2XGtA8VXleZiYLFThoJj41pstA1Ypzq88sLrUfrAtU1DUjP+d
Ho8wet4T2YzoSJ94ZJhEyKgyIdK31B0hqQuMRxaknGODHbmN9cxNaoogUOOfUT7B
O3P5FXRDPTHs/X+vE5JT6SD5YMi0lLg51TPm/6CONpGHRG2q6/H2R6HbeKlIoHUO
N1wJEFHP5cY0PO/diktW4RQrnXplvDazAGXPAGo3AgPxQsXq3MvQeep2yiJNhXMW
axxpFa3in8HyN79xQcoswxwJu5QSjiQA7yquUpIwVSy8F0tO09cJPWMg0sXh0kGS
hHVqCAOL8ak6pHIGGG6cIdANttJdH2z3gcVfcf/sT2qvq1O0oIMQQUNDN5Yca5ST
MMulemr9vRSf+OJhBbyQ1wq/vll7Tgh5RIO4isJSJentHDMxus3/+2zgg+9RQ07N
shGhZxTMmZmyxDFl8e85TR8QflO+tTqJyT9MSHa9rFzK53RpIOwBuqdraZ1mjvz3
y5YHqKSLBsXCwJPL4f/PrKpBVmn96QIuxg/O4+I2zik2oZ0tsrzWI3N6gOHk4hA8
3lCmIy/+ezxAzjKSzckYMchwkSOO3Rt71ilUfRcaJTyf+LBIMynTPli+x089DKoR
eV/0DCzBkW9DEN7rEg4Hn4KuGxrurb58U70tyBR4mnOM0ETa9TJU6V3havY2esCO
FLtdxyVWnZsPOC01GiBKmJ2KLVwMQ4JDU+/biTbT+IOZLmaCzBs6camI4epF/hmV
OW+QhCdy9XA3rwaZo90c9frSTgl6e9Nbw4war+D7xZcI3ySojAfCWZ9IL+rya6uz
GnU6wCp00Vt7DHE3F+6c+/Oo5bW+AHKBY6TRjaXALlDKTYxKGFGpGazBpzvimrRo
sEANHaS0W144ZevOmJDAl4jn9Th5kD/hEIbVhKX0/5TitNizyRrBq9detUzfPTHZ
EkCCKKAQOI7Q3NbRAkV3XGUyBNbKiILu1WxYZE4BgHnoVY7inti0qb0+J1A9bQhu
+MJ5XzdRRg7cePM1Uk/BQXhrRkV54xGBl0l5zKd6V46e/1Q4B6P667NVdgyn0syl
nVfFeAAMEb1SJ5zZ7YW3yVu5m7Y8uj8ZvZRAXfmtpNojwvEv03swXpJQ39KjS+K5
76oTDx3l0TZe46j6hmocbsXrbXcKDR/bc3lLMif+W4GxzqiKpGCFc185yp0HCpmj
65iSzZ55+5x6DAJaC5Bus+IzxFc1euXlhEFpXoiRiYqCa69IH9nhn7D21EPs1Spp
vSFkR7VyhHzTAIfwt9PfUl/uQTZ6ucRACbvmosE7Vshv4w6zuvRIsE5vT7EFZ0PU
ldAY9oLV21q/WKq3cA6IZ2oclJJ/LxHBACuV71hfX7t1TfCilbVG/ThHvpMV8Mdg
7a8FPFRYejgNr1uYNtdIKb28UAfx6lDh/9rCxxLtSJByiWmPcFRINoNZ+YtxipBi
Jz7e5HGQIUBzP25i/Lkra8WZmFaEPd534eGlubzVPbvkWz5JrI30ETXAmJ9eSyJ2
35UUtXDucvJeqyC/gU5n9b2pF/O6acX+FyN9vum1X8qFNLOA5nnGSJEs4+9A9Pjx
48dX/CnV5oykOlX5hxvPcbF6LJjia7GmzaZ6O+aleL4vtHPLhUpZTU6aulB7SRFb
ed38nVtNS2rrcTmpm1qHai3gy3srT5zzHbV9Nlla1Eme1DWJw5tK3rKskMwGQLsx
QUnt8Op7eAzG2e2bK0wTDldrHH7pcEfJoCsljNWoKVlWvlNQHS1WvWdjIEXi6b5U
SHCPXOrt+puMw9M7uYf+9iL8xyDbNTIZHtPryruyP9DqnAq+m+INdvRiRGFTMxNt
XNcQgJfJXFA0WNu1lTrL74yjoVpJWyPU3CbOOEgzxKyqqcYPELKE0vClF0LappP+
5yu9DA4p26IMtl7BqM7xzy41NFSWHYjv+BgZEO/q+aqPqG2K2GopXo7NZJ13fq/Y
uZgb3j5M3UKYuovaF2DXrSIKELCPeMaHbJDrzw7lfiPDAWKo4QpKRgRZzUfaL/ow
dZ87V2ywyry/+itOgW8QErTsH79DFtsW4NBOZWQveVyyfb0Lr0tGXj82trxgd0k/
S/N9KPAmLpSJzU6FVM/CCbe99hbfNZHuQpxSYKLVg5j6tC9YUEwx5FZu0Q0NlFSx
Xzf2HPVBE1vQFiFvgKOxOVCDIb/NZ8rmJIXrZ29N3+xiZIsIrDw4NOXKb99QEcVy
dqeFRZanOwisgxWtJmh1pHw2qaWJ6JjMtJmmhZxnPLZnIG8fyJrDJjRGx8UQzaoj
18O2rGoCcXLCMgUJ9vrjzH21TB5MyAYd1wP59dgxpQeVJt6PIoAWxeFuS17xIGeZ
5divjDjyad+FsXMJuEbDE39htKT99x2WfXvCY9akafOdxvCCzCaQBnBN5BMKgbtd
sqnB1fcvsf2S4/cn9rtLY8EpC2cW1YKvq1g6ky6Ph0s=
`protect END_PROTECTED
