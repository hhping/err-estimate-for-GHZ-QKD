`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uNlVgHr/ko4ZocYuD19bgGfmVH0Baxv+KjLudxEYFJ8GqS8v23QOiJVpr762VUP
DP6NsqITJ0J2+LAIpQgcKXXaHnxbwuwh2MuRODTI4S7I/tx+IwmMxw5VLg3C10rc
sO5FLo1irJIR04ujNBCNUPOMQYAKSezsXE6F6WycmaKTDQDBEnzd8Ko5/GayRjhn
A3r/qPEWmOzgDqtw7SdRVx0tW4XUeKPkPrq9t+EowlkOofNHHLwnIjRYqgUGyI4a
YydsQRArEqeqTFDQHaoyD/bmPiOfISoMIExd8j1JEuQUIxKdBHBdgzQQIhGxzZXO
h8WVLBvk0105hnTBWCTcy2ETUc+UamWMdwznIqNJuXYuYj+g2eXxmyjDD14C2jH1
Bbsr9GOXSThXfdT1dlP7e53+fBetqYx8QjfIoOZ6SXHmUAV8WKRnJrpVydvoFd7k
j9Hn7r7BwKJkAf2g2BmjVg==
`protect END_PROTECTED
