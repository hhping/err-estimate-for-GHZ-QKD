`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPdTXbXJCPUDqg0CqvVk5tJD5p+oWnNw2CAn3PyfdVBMZBMbCKmEOPNxq7pJGcfj
9CGsorE39z/RsWNN2t2pJbWxON1C4+udEplhAnbfWN2U3fjcl7yWzkDh5z7KEtv3
T1sbAAf71fzu5Zi9noxep5wHoY/4gQ0zCimEmoUfI3HscyD5HdEovH/B4iETIXvx
4vBVZ5ABxxBeQnWqzWqpRWSucmQXurd6J7u8Ph03dOJnuAJL2jHACz6AUv2Gyl8t
jRUiE0Zl4ay3ZYdC/yrQwSesPzWJVIHCd8FSQsLTT5Uxok0DOXtoPZYhcSU+BEf1
OQL3o4x170II6qzv8OVNPYhrvrPc9Yj7WaTxGzeDXG6f6xYFN7aKkgHjbz6EQt0q
OozzV2PQdsZw6TNXBWDf44ldsEsp1qOImOvHjVpNCclTljk9DzboW6uApv4uXM7v
nSoq3+jlAQ6GTDgklG4G9bdTdkyg8Sd95XCFEpNqIynD5JjnZxw8BsAMzAIMnEnG
L4/NzXR2XhJNZydrDsVtXnnjFKbY5bNtl9tW+On5gtd3DBopw3lI1oh/KAfble9s
oaELk2zfhgo/azvroujNteVIgFoVVG/ri7c+dVWg7h10wNYzX+0zm1v23BXjYBYt
Ju+XIhz68icL+iJ9FRS/uuoCZb4bVGlyP+SNmQqh8yqe1JlxB0NJI5XXmjoM3G01
4VnQ128AllINTpAkWqVBDeuNQtyv3XhQFnfOCDs5mZZWGKcD4bI3y1BFGFf8/J7H
70Lmmq2yujkRo4JlT8MEAcY3ymlZLKBLEGLo/32gHkgzRmv7hrABRiRag36PtK6E
aF8oRRpokBpHiQjgVFX556RrHSX/cykC9O4+e3hAkVWlrXoIBuEFjQ7oT8a4Wpsx
exTibX20J1CEhhuDf8PUbcehX9V3SKbxDddouIbEsOjXNhsYVtnWC9dtLAP/OuLG
l/+hZknZsWPbVbG8d1ImOLqbQUoKE785pg3Fc9QNWL5EzJBFGAYq+kyzn8UAsWY1
NrFk6uMn+dB7owROEP+UNk0SReZ1YW5IL2n9rMKzpQmFq9UDsArEbnxG4sE2AO1f
R40iwQnRBVYl1hwvTbsHPG2gr5OHyzVsWq4FUWKcwAwG6px7MYogBXXCy4YL4udT
MBN5aDS78fnYhyOZoGElvSu1hMF8JwItQbpM1teYYNBEQ23ijk4zNtDgkvB/qRyQ
ALGn8Gx0ilQeEqcFXgmfUVsfVeEtr20T3Sy149QcL6FsZ+goaYyzMg3Ok4ODBtje
wV2IWxra7kDisXtsmkxU0gvB5zeEPUtghCLbWjJ0YcMlyPjtNKdRdxuwlHL+ENvm
CUC1iItc2A2ga5fHvT1WAY1fLAkX90e2uO4ULKJsId2pA8vOka4aFzwBo/owax6y
X+pCQIqHmVzGH4Ab1+K4Q8mJDeKb8kV42MXzsC2o8SnvTWoPMTlbGJfuYd1XdPXA
cgJkjabnlPUjNYphmcMvdTxK2l/8UtqudpKiU3QEVsOnHJu2LStUivSfwvfJszAN
YXQgG5jf7m+CmShVfdkyfk52wrldq7pAKjZzfl59Oxxm3d20e8JF2j6I8jcGRvRi
JO/DVq1vrwXmD0NgnkHhUtrkePq4MV02VE96v3FJuSZ4e9aTuwnowxv+d+zzoQmb
azaii9HhFfI/3A2KP5dXGvziHk2v0cGy+lOl03cX2wzI+TpUnzVCmIx3Cc7yJ44j
PIFOXzIGNZMP/N40Qw+YY2o7LdR2uK2kbQYfc6V7b8QBBDm/ZspSxs9hHEyku7eX
ejmi+ttVsgMyQJHeswwkwvlpbpe7AdmyyNS9VpnLgFubqBNlsBVk1YllOomb36RV
NSNAzdIcb3bAZYNjmXUoEexC/kr7iYjfh1XuUsKVWW5F4FJHAH5SrZlhWohk5hGW
kZMV/QYl/KIiZTF77y34Ii9zBX3RtUrrPZHvzXJvuktSkT4waEVuXvgLJYDNmyYC
0Q+nkGnX9paQvn46AQRcuY67L6W8zUpaqpYl54MI3Co/paz66Rx9DniL3ar/cbJq
Zse3gtzRfW4Wmt8unBGc9gDdg6fqaZ/eKMV83mX2Z/m9xXStvgYwgKMASNMpRvi8
HIuxf+TWGnFQPNriDlQLn/Iwy+AAHw1HnhVJxThyomFd3tECHJIYQIo5Cli/u2GJ
LhGb9WHnodc1Jw4bZStDD7ysObZBHDsZyibUXm0T1LX84eF2Mb1+EYempn2/dlgq
j2kyhKSWfUSs2UrgTQk84duXyOoNZ7YztlZI1fup8aI2NzstwrRCRK2N5Sdz/Plh
8fu8RModAWP74wlzuHHk4hw+46gacJMWR1YAACY7d6CWpPKCZZMyDrJBSX0UdDzd
b8Y7oIGZqbBITOncFKzwTc9zb8OrRCy4XS7MoQvOhFCn24yeQlEWHRRM/FhGxmzk
NH5+di/Zn/DvgVjS1BrtMWoRNENqMo0JKX8pCN+16usRPe17cb5+Cf0lbSA/1qft
Gl+XvPpxlXANhK98yjJPN/umOskgrUnEHxBAjedZKxFo+emI2wG7a+vj1QxUn/V9
ehTEMaYm7ldYH6xdx+bzHhPNMR2Qc6JC6dx+MnqYq7oIL9jusbYZsYy0KFKbjRrW
fw01k8+ruOgh1qI84REUu0tsqhzexcbyMFvEaLOBOY5Wk2bjRvKb8ZQX89iind75
V1UOWOKvYN0aYF5Phcwc/NH8w5gwyGG4rLOVCwQIq6llQ3jxpehLtVBt/7rpeFWe
QGWXrimnFqGFS4r2WoyXLa2SBJJTf4lf7nItESvGZB0LSHjUuD6l+uiQgO2vrZbF
ei3lO/xrG61IvhKWwuH+By7wODF4KCa/JlZvyEFjWW3zsyxjvoyErBN3LwYQeRcL
77fcK+i8DJuLR/rhORGtpaMQUowdQHoEMfea6hkTgEGygkQsAi11MMZys/LM0Q7G
jykD4Q+CzUM59FuDwh0l1ziUZpBFzjdWSfrF8dvLTL1CP+Ifywq8O+Jdo3RLJ+y2
XusuN0MBSfccl1mCfvvRddG+ALzpWJgtEo35q16dKRDv3asFM220hI8l/phpHd/a
M92qPbM9a/ShrJ5FPuQORj3s2p7l3uG6QMMbicFuS2ZlVOYoWHIkU7/ePumG7IDw
sb+/lvLRGbTP7So0TSxk7ly2rq6xmgo7GkHuifc8YyNdK33FDMvxYjDbztZaOEDN
t2K6nb82BqBOGRUNfdKr6AwjANe5rQkPTStEexIJy79hMbQKSFrquZwt7Wb8q9Uj
f0SOLVh5w6DdoqUhMIkz6lDgMINIINQBnF5qcmG2i34V2CnzGMVhGlLlOSCR81Pb
ar4DCiOITSiB8etue9/Jm/zFoP3sM2/BTsBEvsZBQKECk3kzjGtYpvp9v5ajEBvo
9Hb3dvhaHy45UF2jX15weDloYUi8uHFvGaf/TKyujFbrQCS63RmibhjK0Vf37mpA
xweNHPiJMwdlm4J4YjDIyrJp/mr1jZ817RfUF3wLBynp96G0lwwKCW5iM2JAn9Dg
WeX66XoGoVKg4oVwUUGk9g38zF/36W0+0vBszu/8sfj8rXk/jGY7JUq/7HMDz8dO
e2pqX//y2PJHG4SzTsb/akVsZOBZyn7ixFtaCIuMSZ5TL+JBLa4aCtELOhQDz9rs
XR6F9R5wJs7f8Yal6UkRIlCm/gRQe91Mcshke5pRsyw0hTURXBcucaUKd6ZO/sFa
q3+cRs8zVyfUZegbi2ITgxECaZQ+SzeWkJOWc87FT10AO78qzz01r3EOulBoQm6Y
A+wHB07yRtCs4lPdlW/YWdlvnAeVlx1hHQ3K80rjPtb/4ZLz9kMxtjtU/A9AoC/0
gg742gOCAZhAsBUjbL0AYK2CwPPsd/pwdhPsyi489Vn/afX0lBkHP7XYUcv16z3W
OE+ORSy+F9nBJBeO49+YRsJwM59eQmQBbWn6hej1Grgf4GpWOLdtSzeiK/jtyrQT
Lky2RZ55b24rtru0fTUgNWzamL2YonLI+Vm+qyEYIrNUqABcdPKTSGcQ6a3WtH0Y
7k8vZB96RhRh8SbhOi6tUtNme0W9TD3xWekbXZm00J5i/GHvZXZKNE8anVmU1SMm
QTooRb/XGSu1vGepexqhqnLLbiU01AhH/NcWEVRVqr9mJluBozbT3m8wBePUbBgt
7oKMxs8F8dvhyKpTZg8PLe+kj/p61vbM7MGsg8x7EbbeIk71mT99gSjArHvQ/RNB
4POm8uV9PkuyjZsEe7nglnJBUvI+G3Z7dPVARZqE8mHAUpqtAj8tqtmBwwYCVlvb
zr5eoqqByurnO/WAzfBkqa9Wr9JyA/Ts7/ZbF4NMTpgP83m+y0dZaRc+iMq3s6KQ
RUv7dH8MP5Q+zU//KOuBl/b+VAGNa9/Pqqb9kkQgfXX7lPDs2SPqh4UoKwBeEHf4
j0N9plcCQOnRlHYqDQOloqmxr8tX+lEVTZAQLOMNIG7iRngVYvpJBXTZ6mEIhp8m
b0tQC/2bjgOP9VNQcdxnZ0qrFYOTIEA+HcXz/tHN7HmH/HEuEEKerlbtS4LmVSfF
KvNahB2+GVDgM9krcGxfxLNnS9hxj7212iSMuY1EyEcAJPYQzuq2zw4xT1PswDfy
0CsXIiPmT7VqALwK5q4Xr1TdaCjnk1RdwXb9IHIvzGelN5fW7TOkDnmzOcljazf9
brM4T5PWvTNFhkUiab8Vkj+LLsl+Fdn5P0VjsMqriUxlN/L3JS2PPTSEGGszOmnK
5JNALj70FjWx1qnTGYIQKgg7Bneho4DgZbi4enmnQyj3WPdusbn5NUfBVHrUsFCW
Ez237UwRf/MybfibfPdwwuhaJvxc1CrFKYNpia+ouQtq+6L3arKB5hsclZB48k9y
6RfCP/dzHJ9h06149W4yZDDc4AXX6iNPOaGXncg6qTScSd+ZrfAK7vLmX0iNl57w
SFBaMGgPOKnWWvfqU2ElejwgDDWO2+jIC+QIFPGF/9zogiVBeRw4AQZTeilsNaVA
yiOQnFUM45AWKj+fSx85A62EmOV7V8eJb4e7y+t+JhH6Ynmdva7hBELx1Cwe2Q50
UJv/CoRzbQtrxPDGabMsleHapc3tw/Rw3Pd9mcchRoo0OSJo+hB2f6gpiLNreVWH
GvfQkg+sw+BO1GUI7dJfECGL36L929nbLC6fQvPVtKbdpozyFA7G40FzuP+4wbDX
u1ajK7cUMu7/hqOIXEgMs4yzMJzixlWQXb2f8bFUvcbgWWson9ZXiq7HlGuQfF9z
DfLcYxitZxqWniEwe+YXSsFq4iw+YXoKCKNAZlrKZh7HDaUEbblsG7vWdh6xDgT7
UnGbRwq3lzSbijoyj6FTPiuxH9XPz+LswLLCbIiumtzckwWhi1aJOI2wT/CEy1bJ
LPh9FCZRu+ijkZxARDZja5V0I5VcJuQ/awX4kp2hWbBY6W5zlRYks/LZwRdvSHbO
yuWPMQGujWI0XrhDTE+ETNG7W4qPxZzQhTc+j5SFVdE3NZ95rkPAKSO5biwapQNv
RFppURFxFZR7de0ZFeIawq2r4YeJQUD7Hris72xz61jONcpZGk8jsvHSZVPuW0d/
O6K73V1Svt6QNAA0lE71jsUeZqMadl07Syn909ROcFRC0GP1/i3IQ+DOFeRGkQpC
+sDYbYvKy8kruGY/5yXWFG+6v7IcUp4cfeqg0qry1/FNJg0GTw2VDXBEoWSXVLRB
rmrKQlyk8BZLVzzQuv3JS3BplbT38Pva0FxW4az0Vs9ZxTpLuBcn/AiQjhufier3
Y86ofCmr0dyyblwyI44He7qW6lxSMtFGEZBU1ZOt6EsNNi2fqbyVoK+fARP3yHvM
uAR8pHATQn9YG8qGl59knZsz4so+xRFlucilDWuANJpQXeabmJHeCDsmLPlhZ42V
toWgQB7aN9jEFqadfvupIBkC7RTKS4LIIOjUqXly0q4avD5jCT7Y+hxITd0BQHtN
q7J/vT6JRWnbw+i1jcHYx/Q4ocdleKgP0PosjjA8WVYGlHdKoE2z1mUzy3OXfDqn
SXfyp9crHl1i1LFdxcfM183geerYnh5w2yalYZqBafegPPR8UELkk/1i48VuQ6id
alYsLZb9cxNGie6s6xGwhbAdscpme1tRBWsC6Ca7jF9jR67VTHUmMO/BqNwxuGAQ
pwsHk8GWs/bBlnQp722oIlh5yWiWaO4W8/nrLIo8ZJ/QCHhalToS+2TQ3v4XhYdv
m+5hHWRf9reg28KXqs22KHoSeJtl6UrqPtSwjyjzvYCJRwItHEXsgs1/7Iw64hn/
WrdPBIWGvz40nBxpIlM9NNosOoj6OiHO35eemjZ0ff0HHosxc466UPmMSBC7Rnm+
i9mZsu0eRyoynHc/GsWQtgOdF2BW3W2UR+7+8juVMahffc8Z6ioq0qgGuKM3cMzf
309XjiTibw1aGtT9+W6s8zLCUTornHOlvMEvW1Dv0rITp+wUx3Z61WDB9SnUgh3V
nSGOjhtItzZId1CzoDjDTFG3Wv6SBDMq2scMd8E8YcjfZY91Tex5Qp99x+7Qq6UX
t4CQroHaNOZFaMyq8rpRYYWyVr65RiSCEk7d1EtqrV30G+T73N9NF5/owXlu/0jw
PZjZO7QQpsEKJvHpoXo7AubXVInDfkBGo7pklOfSxeA+Rgmva0aZECFpJy33ZOm0
gOvODiM7UehIkMARrQQop4nryIJBPd7R5cmz2Ge9tWeMxlIWfxmHcBoNhvo1rlPW
dBfb4tl/kwUkrPTNZPpbXdPwiT/hAYBsUhxu+wNJ9cJmzKcy+eBYwneeIcE0Tl+b
DxBGyh+57WG8kTBVUWjPB3T0UIDWRk04oMY9htMfqwqIxxeN4Kr8seVKu+PtxTyl
O7xLFNmv0trzl8vEWwIXDoVRonsdtYG3qN0jPuBtxmG1xDjfbU9qhxKsBtT2Z7Sj
40YFxETLNReCu+/YBYMpuvhE3g5Fbj/qR/FgAwwruWfFjG3J1R6jOtw4xJDpERTo
sYHXHuWBFD1fQWSXg5ySoF0oO6RTbXay1I8jHZ5QWbbchrK+XzY2v+noFVRazH3p
5Bzzyca0d3akgZW0/aijdKlz7UXs+hia3z+PWOyAfO20+v7Ncok5jH/WpE1ofyZj
md/rAEfDZoxEZDmuQlgphthztr9YbXAa4WX9GwFg6eQEWTi6lRRhbjinBxs4V7le
QBxQqfp8Ig/wHEfoLji5JI0PXuh7ys6pkIBLHaNxHnvT1qGeBCHI2xKxCcAf0iIq
3VkV+eP8D4w7j2TuSaluDpeWT3XgmAGwW48EzmkNU+T7p7XylstN1LAg2KzapBDd
CPkr6tsprgrVQenTmb4XdyIUFvVK5YwT60zUzmmo8gcdefrwBKv5ZMvTpCjL54oh
NWzXKyh7dWunbSzeZI/6nGePeVpbqpFU9a3V3WSDHuB+0SiyNm3R1cdJ3b6ukiqX
tls+kjrCsigDss/HTvhx895/uExoMHDs5PkI919+OFnz8nnKC7VQ32gks751VrfS
qS81wpt+3s4ojUK9PNdHnPRDQW00RUSchp3Z7JuNE0Kq/aMKwhkBN13GJ8qMHy0U
trcnPepy26oXPahepk3d4wH3ujtkD6N/qOpp3IWLMZWAxWwLTMswmVp7h5Eti7Lk
6LnEYuanUoTfekgq8gZTMh7gOjld6ckrOjN0JLcBGNNU0eLMY77EQrq5KXk8i64U
W0ed+CoL1tcrbnCikc/mO51SQtIKdPVYSy3MwO058ipPeL+dt1AoRlBmb/Lrx4S7
TI9pkf17TBHyVULJK+wkzXJJkZLxJKfdUD5leue1QmQfqvX4jNZji57bx6LTvIR2
LMyRyJhSX1DQaDxZDQFVvgcicxqq9SFyi2bsKHi2Nl7Qg6NkiqgXnF8BP8kYDH9e
8aZJQpgOslUUxaCozUufqES54AexZUP2/ro6/AR5c+18nI/UQLy9MHWh11mivm2S
BnI5EKB5J0WZvoJJ63g31tZA5LcJfDdFcPQAVBeLvX02NtZdXRZcffu0oRMRPQZp
Rpiw7oKeqHMoVkhlpcxCkzJF/JrsWRX77RFNmG56y6WhsjQ7hohAPG6cr76tgLQt
GDHKyVL2iCS0xHR+17PfUep8vhTShhN+Bvflv18PZXIIJxbbe5513lPQroWCUkFY
XDZ70WmyOOrTLNA4+Ti6ECen9PpOhY8gZXrJGZhJ9xatcSHMsTSKAX/3Z5fjGrT3
oKsYaNhCw8KH8Cki3bZinF53VwC6z0d5F+YUrnCTPLeznFpHS1Z8UOUukrweb8Vo
Q+od+C7T0+4rF0ciZCfgE8bUQGGuZ7e+1ZEmLpnmwqGP7SdIqxe0bCxn1QyWeVpK
Prn4DO5o0CfG6x5hXNS1UzGdPMlqpHfyE0XwNrk2EAEDvXy4e0Lb/CVQw6j/Ezuz
DUa+Ok0QB8eQqMLwM8Z/LdkkhEl5+I1sWZk/1uYLK7ZzTXw2XPS6VODb7WnaFzfT
NKctYhgEr2kAPZ6pnA8kapE5P7RLx/AW+gvNTf3r+xKpX2IOEHU9bpgjY2rHtbPY
rEin7ESf9EGDgtlwP6A6Ot1WDWcP75OvFSzjVXi6/Kn4fgz8JmHsRaCMY2VsA6JM
e4fAIcfhVQo+zrekYl7ggs2AOzTR+hFfcyXImLfJw1AuuGuK7Ya9+sVxDHUw7G8n
mRDIPj3BjS4g91nk7vJw2CjCj8pIInkHjlGXA+OOm4XIFEislOI+SwAk1t1CQXOO
wRdvPVcantHy9zJFCRwibnY13sh/Fj8qClPiTsAxwW3CpHLlX7e87QFfXYhqZb0B
ijvbzvpWS3PiX1bnap6HVoApTs6mnRXfXyjFt00su8JJYpPmv1HpKcZcY3dp7Tsw
hUs8C4736UPBkqqUjOXSfmDIJ6jJW9Ut6YXBeDEChe9MrDYH1sFwVft1/2fHFBvC
MPemcVgV2242EEuFJC1aonGG/mrsdeIUBFiGU9ApWhOZzmBZsef6jcxiqvM61UBh
uSOxa6g/Fr9thNs1rEp61DKsjXTW/GfTrWXH0apnfvBw6bAKufYbe2u4ns3XGBT6
97QNMANpNR4/r4ix9dF80vzzn4XWbnx5Df/RxlYdGUAYPC2yjygCQgkVxz8p8B7+
kp2Aj8oedFLdJijKw+fM5y3jS3U+50frtHf8EYLc8VIGS8huK7bpbsxup8L+KNSC
9vhXDhH/RZv2QYO3pXNuv7tUh1Cm1HFYecInJ5NpqLweTJsvv/OUlgFyAfQtc2GH
b+L9qvgS1oyj9AwXR8WA5D7P+7Pps0W/QlNlFmat4XADWa2DQX266YSneSnJR18U
xTNWPfMr5rGVIx62rxDN8xap6WCgDULsihTMcu6mMHOtHRXsWlYVtfnY0RguKby4
oI4LbLfr+e0FwBLvvIJ2Vg3GG6oYfbWQ0wQrdoy+h77NQvcixkqyuLZofeZVoOBA
jE8sbGkZknO43BTsAfvRKGe/LOtefccamIzpIOhvAHIuxl4VuCivR0I1gKvzsJU9
2Z/VQKZ7KBQMoLVh/FarwfAguWel9ocCNURr/EzhoY3daDHJjhRTrLXWQWafeQYj
zEFk15IplbjW26ofk22cJoZG3Y2Nm3dSx6EP4XmfPj57GMOjd5h4Ts8sAZU+tRer
zLR/kxbLFI1wNb+HlZ8VctOaqZuF3xBjdXtEQ+6+6VmPXE1MtdEmxOjaRfV4kiZU
KTtcaE0svfyLd21pFEoP4gRL9tDVcz17PLRvNR0q3nbYp3uHp6r6GMWReDEYJ/1R
k37JFyKuTBpX2I454RY3udzehM9UjLnop2AN2OQ4ETNv3wC6ruFa3z3UpvlHVe/0
ZVyXLp8dADwt+R/Bt6Fz4Le/VAhvw/YikvC5OQNmowu9MIUfXmJnfWAU+ycHFqQD
0InKSV6aPIvjYekC3CmhAVBjG5T5uNJjNE8nuxTPGJw31GJgRPpuaBA0KHRavsiw
itAN5M72sMLy5EzzKxgkKy+q2RFMttD4xnEj8JOfDdC4tjBYzwAWZ3BFmUuqTenr
SVNawly9PleBP3hGfmVgsQAVDVyWjqUK5BBFiFRjgIzXK8DEZg9onla3ZKdkMw5k
ZWI1dWkrIZ1GSycidREY4lXabb6YGeD0lWE+P4aLajEMV2esHWgE7RvS2XvOEevR
kcLb4W2Mhz40lO/Fvx8OvLWGngF98syTIScQhHmSepDmdamc6/jZEWEbmqNkceQG
jgul0oH3zILW96EOBmtgIJG5W0M4iqpiKJXcjVJkReZqVpdeMB5OgY+IiftFSjCK
Rp0IDd0REzFo1Hhj7jYPQwkpY8A3fbTn5/x9oV5vIh0b7pEUFUyQY/4iYs1Q+4T8
7uuINqS1CkVuxWLe1YcOKSmVvzsoYDYoR7Mc02Qx5B4AYDQKQ+ow0ArVy3zYqqLZ
HrkKmiiMSc7tEa4qtbgwscoIO8kmfZeD8Gu24dkAV/3ps10wgCtX/FWUBKa62BsF
/s1saf2TlGfS1PT4tZIv2fNF+DLC3Ky3m9fAVyuGIwkqicS7heCzR/rXGry2eR0Z
ZY+VwYqm5Z3vAULL/b+piuq3iAPA3CCMg7ojFFV2RL1R8H5eQ+2ORfhqQF4G8kSM
Hv5U9CgRCcrjdUIQkfOfqgMWG1iIE9blEmnLtFJJ+PDGLrzyydVGQnJ9i0AuzGpS
n2SjiFS2OxqdgoJ+itgdRWWFozXlTpIyby7jfKkPayJv4N1H5cbR8kSQrWtXVKxS
GUAbNZSQXIiKGqAg7ol6UPpQYzsnxhem7eC39MSaD538sYGfdYM43Q8aSP4+32SQ
QG3QG8TLqzh05NcwWh3pdYn/byJyVctsE9Bq5XOAlvhQqEFG+kHfYerBEfrzONiC
Buw+FU+rScsuIOy7wIxsAlhDCb0P5D1MyQNZggptDiA2N72GwottWjuUPnO6v1rM
bwsVm9PDOR99y6UWJjn+pDZzQlQXCCwEAfJ3EJV24ZapozjgOHydFoMVguF6fHX9
ufDUmCbuXzjzSZsImJsVj2Vy6DlDx9cjd17XQUZxT7FXw6opWBqn2qZPHXwfSfDO
qjh/iUtYJtJosHk3g/DOJzRTRtU4yb3rrlxhV9lRh7HSZ9UvznBignTUXRsEpYhV
DsIDaqZj7x6vvTM9LtG9gF7NZL0xxRnCo4H2+wuQ9Y1FD/jZ30hStrD/CjFrMnE6
x3/5zKETAxBiuaz7KhA2SJXgG+k2LQ3aLzVppY4vs6hZl7MNx7h1Qqf3dsa1I8Ak
cdAtk6tBc9RIoBRRlMCSzrdx023NAnyaPkIcuSdpALoxBseZAMBAZbk53aC9coQb
A475uMbOzIXH5SBx/moM16aWoKfpfCrmjqV41XSoJi5kfpWaH9jm/vZYWbjrrLqi
P5IJFyCZRPqEb1gffwdO82dwcJ/7BqBnXHciyzMNGjl+biyGyTeABibg03pVC3BI
nm9RfVqDVURVnRdhJpjh2RCNFIj6NLl58R0WM/43YJGqo4ONAFk1J/m86Rt55Kk5
YuiCuBqR12ZaaqcGARv/CLASX1H5vFfd/61EIYyy+vjyvpUV+m8UZi1+eJM7VB/0
0yQjGCjmHKGJPfjNvobkebvjfRsx7ETIG2dZY4bdZyqymNuFVSd+ff6E2yzkoqke
Qr8cgGm4/wQr0mhcYh8y3Hw81wa6g+Eu/eWla8LJtrjlOQ+0QSAcK3vad2zF/yEZ
okGOj2vu55ERhe2Eot5T6F2pXZrSdhYEa/UD8JlkYt2nfKYyaNB9fGb7wqaThMsN
UAkDLkkNmWX9ZxJTxx2Ua9HGGzH92Qk3TXVpgceCCE+nnFs69bM0TGCE+oitJCWn
yG5SOpy/KIPoMMTOxP2SJL1A/PGHkhIqk8WzijoFsgTeRbev67URNJb4Pfi1IABi
wtulsCsf1lWWPQ45OEF2u3M1RBJUk8qFJY0qwlX/7BGt2AKFnYbi6US5q1v9mWWN
KqO33yOlx6+qtI397DxwKr5jhvuawMcdwRQPb6hvUyNKhleQ/vtxASS4lLcNP5hm
3d8gm1uoiv/sAqiMdDgocjShVEwET5CxIVtlbyInkn9+9vTIcuChsQjgRHLKyvEU
CHtYyaUFvgoG3x3DqV21BGAQ9ULJ+54DSph337/Yaf/0S4gnAkVVstGMXDGasKWc
lKesp4QWZ0zgirNP7nD1+9ycqOnL0R8eQu9vQgS4Q9E98kPO8WN2hMAO+PEVMAdP
Fop184wPqOYe4BoBCt6XyU0lbl7ZYdbbKndinHqe5rAH9SQTtWMeVMCYonISIpiJ
iqdDBOSzblsqZUpRv0iSSc/Bj280Djn5Vvvzq5pT+Z31OlNf063ZvKN+998iDe4f
bMQzWZXLETptp5sY00181nO678OSJZX2YTNQEZ1fVUJE/IDLg6BH4cQZWvQ0EkmQ
qND3RXtsBdG4FAlv9vGgUsXNMKh+uM038z0lUWcJncA/14cdt4XhMzKztQ4vzIet
/10lQr+wtJ1Jn6QPWWpGBX/SmZRw388gT8trlBhBeOn/WpH0Y6dXd+GIeBEE25lv
H1mXRtXmQKbzOZCC3O5Vv12wZJ89c8T0G2mH/Wwxb3JcviFw8yZ/uJ2t963iRGfA
W54y7HRCI47pdK/OcS0vgzB4PFL/XlY6f53dtgTDEfV/vO0ARUgFxIWnm05ERHQp
KuMVtQMHY5XWUslqw32VdadfnYESPvENh925DfIK/QgskBbHJ0jsBCTasld2DCUt
nj4Xm8hV/Hhrcr42rY9SysITdkr6YmRz6yEB5iYCpvCzyG6hgMu/XbNMLoJdoCOC
zWwAy3WDjmoYzBSMcVHtq2YkA2dDDBxnfeaVyb3BDQZP/RNJj4ovwaRnPT+c3rJM
gS566QuupSMqmQbeA/iZRn06kKmj6kOgYgtWAgrgTMxgWr/LeS+BpwkkC2amceam
V0p/0g9ByXc44CBFF3thgJHZO5PVqTPkDijt4RqKj9Cw3tcI2qa8hxTINntQOjt2
3Frh+C4dLynPsVskGqI2V2mS0K+z4jUqUejWf1uYlvhfP/XA0MJyjbv0a60Dg7Vc
zFotWnevru87NBbYkz0oZMNS9VXBbzHAvCCobJBBSi5R08XWVWWcDpbg0V2CGnva
AyyguZKbQx9nsKi9DQkydemRFcyMYOYR6le5yqDMCQoecyK+QPPoRzMAuOtJffye
Uogx6A5XAVBdcWwm6wsLzPjZyZiwDzsArJWoqPVvSIvqaF2M4+HLymQKBWBtU1FF
Y3Bv8ON6xXmerXXjFeA8JaL8RHV221VxpIDE15IPAjbd1wLAjf7UlGDWSmCqyXYR
BOJCmh2Mm+DiI7LezSGvhI8l7M3Jw1ANY9ZtaNj2ByFR5jaTB6VO7UA93QWOpEzJ
ESPnIwDDWbAC1za9ZK3QThp64W43760sgxhHk/yyfHcuUzseZ1+Z75kgqcM5ouzx
F0AowzwLLh4qkTO6sSWaw/p6gusS89BD5sW4gzFiJsT7KTjiXoRhYCMm3PmY/0t4
jipkTfqCz8FnJBulu7dcG+adJq/qzO00Yog0ztpHnHLZ9nOybJx8MLyINOcotjpG
rf/ArXQZDLsQJz8fZFkA+wGwJox9PaRb57iOSm5UWTJ4eYl7SIzZulxdHPO46UAZ
xgZ0SE8sOSanuWfjnEhTI5ZXBkGzq9xEqJP8eD25Dx4D0LtZcxQuEpo+OzQw2UIQ
QRUrF2TE3IFowiNaQkqglG7HQOPM/4+7Nyi02g7UrGpYr5/gRO2OuFWF+vUnP4pR
XlZK3w/DppL2sFzlzRB2fusKYm9pKhF6s6TR9xHCaf0tzf7FFDZUuGRwGTwiuUnL
TOV22kf7foge07H3KFEPZWRpqQYxA1SB/6y3wy81r4yvuHd+UWqSpBWo29a4+dWs
3FMWi7aWYFPJtOqXxn6V7M+lH3KsHJQw1Roza1v0BR0nUZpIVsxYjiDprLLcNhD9
QZdBjNmjmWuE1NLb3/UcKrvBd0OaUjQGsyfhEMPRVUvZKTSVIKxsJQlj38s2yHnv
JL6Q5qgP/IS+P489ZyPm/UttcDq4ZCyrnrJgAHFGerLHBzKrzXjSFsmAxkAw5i/z
AgseBGNAcU31va0qSxKZU8pfVsoGKfmepMAuNMGb0mZf0D7di3gaYlGPtLpfnRAi
WMwdR0fOwx+3Dm6bvm4hBgjssE8rM2+b07cWA8CrQEYpitXJEFuoiCVdGeAh6jjZ
EwBwnSkpyKV1b8n2oXnFst8ciTfkAxMJCPwUIYtvVHBobQ3MSl8Efip2Wgyami7a
PR9mEQzb3qqrs2iJCsQ3RXeQfbMwJ4ciJbwXpslD97vupVMuT513JZ5wHbbktfbI
E01OBjGUhHodLQYsA61QW1Fc3oVA1NvBGBLzO4eS+n94qOyN2BEFcHfenxl792Px
2LlVi7kGUmesMEYFEfY7iascwYBfs1lMRWStXdLskzV2VplhoduIP87fUXzpRvNA
ceruXrCjYPTYzX7FbX2iWN07H+e/6c3Zb91U+5BLBeroPFQfCj5wmIR0GIaoNRLB
GeSzy7Zg2/IQehfijwEG9MuU7UxYQgZfXO5Xf0R145j8lFyhKgUK5IiY0HDorYPZ
bXndVcdYOslA1jesBBPxhaOPrL4FsL4lOjYdrONjh8PQ7t2hdTJXYb9fGxAEKrxS
1OMR6IgZHOL2QDKqPdeEfSUO8fu+VeZAkb48bkkXxai10a1scKeDMsG91bf8EV2u
DsRUlFzmA1xdsZUaBSevmzonDZTUGCcnNXhYyvbSxV55r2ujP88h1+yvVWJ7g3ZD
0IJ0imLTDg05DqixxQcYJVGFhin3pfaGLN+tNcyeZzXMODqdL1mqIumc/pHn6aCC
ZJAfo7TmQ5ADdMJL36d4p6kxXDsEq/sBQds7g+Jzv5+8gUDv4dRA814yvuL8hhQh
K0bTuNPEcg42GVQlV3hBAv2CeYBf7DdwaMoAt6FfvQ6peZiknGt9CHF0gs+3Rp3i
XzNop/fV0jEvPoHykRHBm1HqCBeLIvhFRX8R45xJnqXRmoXwfHUq3pExb63+80ll
PiCN2+TaGLrb/AwsxbhT3qMl+bqYY3bOlgjDlnTO4wJHNX0YZNj9pkVBPPyyvDhj
6DzocGel1mJWZJ9CjEKF8yX4t+eX3lGv6ffzjTndUA8GoYNmL+p24FwTWSC3Fi6G
hUgJ4KZ7wZL0nd+OybsVziApUJ8ruj+SpC1D209qDv8aOymQavowC3rD+QJnwrA6
6ESVJbgPKxTc2U1meX5muqYIJjtCKp0f6+cX+OP81Iudw6MIE6BV87Vd/OmcecUR
aTuZokr8C+RsgddnA+dpKo7qe1k7ROViztqcgeFc6208aEPK8r6KRKWE+uu8fS76
g0QEGIOScTCgMRb4O2t75XcsuV3wbcmw9mwsXyseR62rl92Uv0/YMlrTRsNmBKvM
u/L/VjSz2GUJsr7gV9oGffTrLJC867JCdSIhVRFfN2s+kuFgGs/07W+LyVsjm9M7
voVKBjajylNnPvzHR8jFEJBBy04mKCUgJwxsTg9eMPHRLv32i7KJYZWGeKcCel6n
kZCnvzT3cOB0Xl3z7oiflpdJXNJbINVDi1XnT5mp+ycjwT2cEEA4dqt1cN7grqxi
J4xvg2GnZPAedF0ATM9i0PdMPoMDpByE7Q/D/c9WiuRpN67yhBxa8UQAqB5ymLFG
YItCy6QQggqgzSl01WvCvQm+1zi7FXyccZSu8PC23ys3s8JJcA/Jl35arKmWT2VC
r3U9EVIJDhm8rWjHWRrR+9O0LiBXL7Tg9W/Pmmncj7z4U/0hlrdVl8giVkn3PX+z
tWTQPoMGMctvjYKHBksyo2NiTLBNkyuTaC6A0HC6pbI=
`protect END_PROTECTED
