`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+QXeNYdlrD/+J7HBkT9Rh1vGMMtaBiQFSMHmsLA0kdmB7H2z1vDbiHKYcuuwg1E
zOjRMZ43oAIOlqqYqls2oo8m5lunCmgI17jshg8AbFh5GzFdrgKGZ/dQLkZoUWZv
FPM9TcZv2upQX/mHDx6CbmQCqrKAEZhLfi10w1gEfiggVkqIH9tcohshJIekGC7B
iyhOwi9V9E6CTYk+1JIFNgT2nlYBDkbetEOn5VwmKPQsCQ6D4dZ6hl/2p064P/Q7
gmtIWXXadSLgi2qRx+9xM87dApgQYg+BDT2UUXft7Rm+735JOdCCrtwiNe0VcSc1
QHcfQrIYtj/e2Gs7lndPaTvXi5/fpf+SNpZQboqUQ3P0VZds+dV32yeOQZr5n2lr
A9ZZebbxmjMGr/efpMfHezZreyg47/PMMNSrxtn/jsKfGOV1LeNv43kBOSq4cpC6
tOjyj29i1vYvhmHBYVzyh4LXzg91rhnjw8WyqvsUtJBR5KN/Q462txbexQsk2RvO
4++jd0+o1eJYX2OpJu+pkWPG0UpEkIG3s9a305nWDAkPp9AsD/sVRtXXwGNOwiyb
l/1mlM/nSGb+IOz+BBmAC16XEWG/qFJr8b+lrHop0eC/GJ5k9Goj8F2ONQ6bmLRC
NKqW1WoIwriy/F7nJ9/z2VMkpMWPyUmAjeTNoeMfnNjmTz8BkNhps/fRxjVqj3H2
v6Un46rUmtDZBMllC3TRUtrneR7SrzJH5t+1R4Ch0bBOS/WQfXdOC9abREL5M5lY
dvL2Q9j/xawhFitS/XFezQJQWQft7497KcxdhqsIrHRTG6IIdbN+RWTx9rSmzTmJ
RicF+vfNKTP7q/77i/f8t40vMzUwYiCarASJjdL67c1WItNfID+G45wUpjgUrw2H
l7cz/Xn9TmkCsllVebr6sPZaeFmTs0mZ2CtVkDpDVfi8G2z19QHLmO2w00jUkY/Q
ZYzmK+9pbwMA8fz0IrzhCSxCwsccRj060JI6QBkIGkk9o/82Z56lB703RHB3QNaR
TrFjQ5CrnGHvogtwKPGxDkjdEhCCN6iHpgwhZwhkc2T6NrHAnZ+YvkfXhOhT65gF
FZoQ+LfMfK4uMlCOmkgijPt2RE6Bd7mQT9fD8dRmqZ8Udql26uiI/8J9PiNNBDGQ
anH2ZhQFEKdX8LmIrxJ290m1/ty/lgDXplAVWNSbbrz34XdAs4t+vG5rpl1/Q1Za
nd9rE3bkLHurs1JhmmXBXKjBRR4GTpVYK27/V3hSn5BJijOk2AHMiDJtm96Ha48W
pOsLYuAw4EwBEXsMYzZwM409SfO5ffRJztOhzi6VlxxpryxFWO1yJz7gxTvHEhr8
7RAjLKXx+/aayhh/RueQLDHRsd0iJgmPtHiwKBZJPAxZzO0LPMFzzkKEKFYzmFyI
KICBYnk99hSpe91AG76V00Ps21M8Zp5dIPB4V5puXHA=
`protect END_PROTECTED
