`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMLyyWi0PBtCbdpD0sT7brLPYjBeU28MBRXWvJP6q/PjZWFw6MtPqsHgbi7nkF46
dw950shlzGZr5njE3R8oXPMDVJXSLa/YipCZFIJk9ZAuEWEwMvSwvtOiQHjNkuB4
fOoGOsC03mH0KZ0ZcMmTiNpEpM63Hssz+q7wVUQaFRsZ1Jb/72+78bZNoeB9Ld9U
iBNt131bphg9PAAnQqH+7/599fVa7hAqnakrQnNSflLCZ5969LhBIz1FpHGD6Cl0
5fuB5kdSO5es39iMHWlTW6DI1gQ711IXTvpGmpE68PlV9O4jt5RscOhPCqerItLD
I+wiIB4RwYBtLVU3S2cI6GFrevxo0MuF57jhFlKSaKnyfp+hir1FTWke+/qLTwxm
fxspcCR6y8drCn9mzNh31BquS9ooz+YQKM/pY9GWfAddok0tbCBk0uccVez+efC8
oz2iNMu8PEQfWOKhaWNUJJuE+mI85VbzTzdaxy57FPU+JQIALTEDlV2S/vBtvj8C
85u9P6GUUF0q4A7HnE2oNMNk/4XR/mJ7tJoAORdMjm9Wp2aIebQTSJeQ/VhVKsnm
bKy5giVAOPUYTiDo7dcIk0ce24x1I5D9rJRDd5GaGbLD9ijcw8X9sl3/JS6FuaCS
`protect END_PROTECTED
