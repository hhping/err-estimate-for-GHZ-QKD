`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y79TwblzK6108FDlb1d8/F0/wOD/mk6kGuULe6/0H18lOa8Wh5gDqA6E7orC2Z7w
oeGYSo6OrhFoRJEjZaBacO0r9VZlaTgIIbextuV+EKBLMcd25uNv4lXC4IEAWsU4
PZcU9Gyw2L8r2R6xEk++PC15eP1VB8Y+mXIZ8Zd8Ceq98yJRtJZ+rH4uVMOL5hE7
dPjOtN2PEBS6umqcmgUsKh7M5rLB0DdzGWsSZhDbMAnbNe1dENtedT8JzkZlhZGZ
UDMglxUkgdL9bOnX6dPO6spL2fPZucqVNqyfgUA+3xzyuQXr5Ee1Lt+NTq5MWlIN
kAGKCE9iWqhlDCgHj+frvOjZELgEgZIvUKnZRC35VlMssV5ZgZjUmqpOtTccU9iL
aZd8XMe8lesY0TK8Sz0hiJjOQeoBHlo2IajAAwuqdiSJTSZptmHOE2DFJ/Dcxa1L
77sD6Qp2tE/J3Pr58owZN2wiYIDgnn6p9sxnvkN7x9jtCpK/xksjWB5OctzTok2q
tAa+Xwosxc6JIGNXyFIycjKFyXzRWvWe9Cz1MSgTfG2BgQMZ/pF8LUR6B+6tNFox
2n7Z1k8Zm1IYxZPSfIRi3CLPy7hfkf091ILHbfg5JvEKTUc660th6Cae5qBjPszu
`protect END_PROTECTED
