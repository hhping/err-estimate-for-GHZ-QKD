`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vSGBLzn7mnnSGB9vdxi4omU6HJiZ0HW9TR0CIQhWXVUYDQkvubeXnPYln8VHBE6/
38VsI1tZlWYpwvZd/jG+x8zF69we2Zy3g3u9ARnMEfB6hAh80Q/5OKd2o9TA3pBt
y5JyjdfE/7KIXzQsQhteRxQITNvaCWV1eyR8thVKC+Dm+6PD5AwmEOXH/OeMu2ud
hO3BLyRq/Zx7z/HWqKeLKkG//V6toI2oqUG5VcXSmGgJy7+9PXVdkRQWH5/UugAN
GbrOt26Ps9ptc+eix+10Wa2BeR6fGYzZbZURbGkv5WCUkSdD7RLv9KK/6qDjeLOl
2bilacW760VOZ/Zp8gm9xlGLhFwbx5wjnTlSTM1qfnSV0lHd8KkfgY2FfxdCKUPC
vC4uUIyjoYSk5tSwsxQVA/2ZGa2Psdt7NeCann9ZdQLyA3cWVX3ruce5a3CMs3jy
NhXchXJcy8TVlKNdEjfaK7Ptfm8Gn5uX3yqyAxD+1IjYwHF1skRHShIA2DltypzX
g8kp+tNFTX26OiOL9DhxABVOH4N/3v/gxjy4yuPo64SpY1ZwjBvbyvuZJTaDTl9L
hR0AmekOrdfLFFM4oX2EHb+RcT7qIHKj4TKSHfal9hwLRkYPw2NnVWKEk1cldCB3
qauMq7cftWULZfl2gtmOlYLeRlaWUxmig70/Ixo2697L3DM2jX1YWobQtRdqaUB/
PaAA4iDMsOk6cQGJvwEieoKPjQJ/dpUeDlDFVVpeV5wJBh03yzP+i0QT36WpsRRZ
oBUErFmx1UJeXhUYtjwMDS+1uNP/ht3XWczro4WLqUjfgyJ0GwKRFy8Orn09z0CS
6ffzJSWTb6FMwjT+X5k4wc6Wz7exPQOyzxZXG32XKhl1kFoYQrmtxq70mGzPxO1x
jCeRnPOLmxkjizb1ZM/DTuThQAu62vwezIckW2D7CkrJeBxzBUgBD9aQQ1tsYWS/
XREJ4eqgX8ED4ngtkiHUl2waE3h/0ZvhibQdDfMFTzbncOEmq7E+uJndy5uqq3pd
th9xXXtM1N73s7w6cwNvFVgf/NozH/4TguIKnsF9Oz2Tog2NhtyBUAIrL4hPf9TE
zrqyLkeVyct14PHuBxdNqM2MgKhXAj6A30Xc2w2j2CQCudEm6clg04jmJyBdOkxX
oJ9Th4gGIl2FmD8hW/K0+QHzEpTePacaeL9i1uDeFraXcThIXzer73ifY50VoBnj
T8F6TWDm9I0A04ZdB1WNJpWnluONNuAlSOfZh5lPQNliXVASvcuFaLskD/eWNSpL
QtIyZLHXoRERpNr+iI599ugFd/csvZhz9DWC4kODPg+KI7U6+Qw0jgE7UEc5Oq3t
lVwch8yDMuvzQhw89McqH70ADKhYKeqvx1xOVMIMk6zJ6fJGElodIwqpIQeqgJUP
gpyPDnzh4PL570Bxxl+Od37DAYYUlcijXZ5hXcjorrDYTkOkN2TOnnbQcccAqsV9
rcD8sQMQ7GnSzFaF+4kLGIb+ZR8wpz7ZJKgX260U76MZFreaygtYjrZu9Zvt+vKs
aFD8dWYVXCvTL/gLYvrTor6jNlu5lglvt03fsOUlKeZBPPr6SYNrqPmHtyNNfLCJ
+NVFvgoRt16hq/HfdBuj2/1Ow8NXzGnt81eauXavM8EDaGuRc06F1NXyZoTP1K5e
zpilrxYXQO7mqHsz2FGCEOLRLiUrUjAhXHWMFaM9l1B8SgSLzGH+4xVAy5UolWm9
mjrGNWOT3pkfq+iVGF22cOftAOEIhzZM6o51r/YMRdc=
`protect END_PROTECTED
