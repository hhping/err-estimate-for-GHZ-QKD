`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fm/IGA7BBNFGEOdgT/6S/nBQgIiOoogNxhN+ykQolf8IsqnOHTxIn25laKXDC5/
K2zY//SvDULagAfe7HZoSrap1eHlZGJRs+0G7SK8dTJlky0NA94ed09OxokXT15C
QMmjrYcIUC28ZKCVlbBy2+PtcTErVFIVRY8hTLDfl0PV2XRE4uOG0PY0i0AgkBKP
up2PWIp9sEDNgZKipo8QofpeDZRhvEKnl/xOQiD69FZiSFqE9qv79AzP5xPYDYkd
LsG4D9UT/Y1M4Oa4W0nYV6OhamzU6MIxf6WRIbski1rRPwaT0/ExrhWK9x7919gI
26pvIf/OUtS+GgS5d0MbF8lZ/CY4Vdm6bQnzYuPJ1RRRgjD6m/lfLoRHkDVtl3mK
da3t4Ry+/V13Oe8Uzw5TcvDosZGRQYD7EgzfIynRKdZ+bDXI6yGBezfwj6ATweun
ic1KH6GUvj1P2xri+nZMj0SMwKczgvu6SToYSyigiutCVgiysmrYHkVnb/zjIPT4
QkOAfSGldXk3+lsftE1WyUlUhwy3W5reTDaw0z4C8Ll/EDWL7am+/3yYDM+R+jxX
MoRT+Hhlw3xcyC7YMesB5sCOXBwmMcrDWXZiph31jVrsk+I6cs5DI2cLFMtIrS/D
38XjbYsRWRZ8gNXyWjbTv75kCysYic0lrGIjHTbD/Ec9b1Yw0HnZvVHWb3Ha5mme
flgD5JWQ/XvvLNUJkeBIE5fTQKvtCHaGxiMfWHXx+5Y2WIKU3xrgwPtpWXf93jb+
xPCMV5E1b2kf58jRs/Gjplk60fbLGoWQSOiDhCP3KaFrHzTxZTufqB0fqQLkigPv
Xaj8diM5d41F/2MlSUZzxqd6TtvGR4HGVegm3b5zWDQGLhcv8uAB5r7NPMW9AqPt
9ZDgNDqpu7yxOidJm/mYcLEWnRgykuImIMKeYk88OwkGzZkbvC2vTfsMdjPr7urw
+lTjp+lOhJ4q1ZsDAo2zzamRBPo3lh2TG4IFGCtFlFOTLomzhLQpc1qZ/rhAk12+
yRZyJZuQotFNcwaecTGzkThTw1fqAN8VqR4S0xjetMTactXHMD0yAvr8jnKw0JGf
zDWO7WnRZK3YPMWUBfOjWjFpBCjTma4vXrt2+S+wlvgE4vq31su71hlQInt7DaFt
NeUNrXG8SlAG+t0qZXZGBdg8FT5WWZiLUAfP/6Ya6Qtpb49Gi51erjTfKzp41gCi
E8++DNG84v1L0ERBuyo49BPnmeftLP1sqYaBD2VyzxqOyWri7YSyDq+dwFxr3OJL
ztCE/2NccP4hAW6/SFlzmjXJf1xr3gEgty9Krmc3pmEnP87b8z6W1LblrDT+wnB+
twoQpQt4HzjwLR0gFYzmz6YvsEGPMkhN3Hu0cNt/Q5wnASdT2+C/cDWlkzSBejTq
FGJUaYMIiapmEZ6grycA6cLOU81mv/izuagnc+iL1QTzSMzrEwckG7XsGHwc7fkb
y6anzmo+ImLND43WBz0NkhLRjVL+q6hrUNUz5OwIPsPoTj1LaQsO6n3ce/EuA9pk
qrbzjX58EoLbA/JVNdfcM/M9gWpLJj09HhHDUG782wa/Pmhwo/F59Zj8EKLcWynC
eEkV2Zr0RBANkLH8afNeQC5tNuiwu8XbD36RVIpsU8VT+j7h3MKtLSnztXUVtB9B
baGbENhGQFtMaYRpy3a72zD9Ih/K6EzP+j+4Oif5ENUvM6uIVqE+/ZV8kic+IM5l
QhUtmqZg26qjaqlGVRlt4cFFk2RMhqVwdR/rvVid9yyvuMpdcnMmac5mnUo0B5oY
ByuvNOi1oh88KYySHAlU5RaFY0yg2wHjy/UfRpPd+sjSX2ZZgvQYkJP7IeCEFL/O
04XDeoaa5fPxSP6/VY0N9Sx71uePbmoRBaE+8I+AHkz4k75+bw4YXed2lc6x71jE
rHj54aFqFKGKfO9D2iQcvsGswkYNr4rTEgdKg5ZaCF4hZ4VzmH0V0Vq4S3LXlaTK
GhL7oc8vnduKfT0T5cvETyIWZBNKIoi60WVcV8fYlx6116MsKB7+P5fBgNzZCp6C
ALT6ErbvLkDLFrqawKglhxTacgxLUAel5r8K2QZHnFRMf37tYRpZ6k1wJOMykbcL
I5CEcmZE6LhtajePHDZHIRlM/QzLNcpUPHKO6TVGRa278NxfIw6gwFlNym0ynC/H
XqXBGGiDihmPsxVZvGu/6y0hWWkmiz/R/R4Ql8p5/RIzTKCyThgSh1sc+JY2bzG2
PGvoFGUEWRrlHFdz+3sJpz0HzGvmnRvOcs1R0odfFdS9Flssnsg2jB1JA7iCmPUM
tQanAihtrPSZe5+GoiZqFe4WLX6GHjRiGs8qgyzwjKugq6Hv6eKbbpgWhUmz9mOe
9zMdtiX7LofHd2A3MchTLyhs6KjXYW0O17yidFSCwngWDMmvg7o/yHRZKE3aVWYp
I/4zhHuB2ZgCArvQn1uI/kZl7coUhOJZ4chAMxzm6zQYYTZ+aIz+OnuX5dgQMiKC
IXjkg1cY33bLtHEPYT9FX6rovQcYSsTuVYxcIwBfjTZIdCKff3GUrlc02kid2RNc
uJOneh27cPbPr2hvbOxVMfXKWcYu7xTz866UaIb6MWnjAf48qJ42ZmGLxEHZQc4a
3yUmyBKouF2QuPNBPQkML4uTipXVUeFAYgHkV6i2KzMsJGtEn5LSrFrEJZRjhjvy
2WTuAx/9beVtFkXeTYqtXR5D/MrThF9Oq2dBira6HGJFgm+O6WaUT1JFPzv47cwQ
/izEAja3Arfufn0za/V3ELtB037WQVBrgf8W+ya/n7qx0IzapHt/cwtUaHAKJj9r
5Mgk3RMjIskqQCsbrYuewWdM0KAe/iin/uVqrBH0FRea6ZiR1kB1Um2SU1yV0lFG
1FCcVUGjGW0qXpcjbEUnjnILJ/0TfWzL+tqnZvB0oLSatmdtysxCpdXer6ppvS3s
xCdqpnDws/hXFquJLA588Czgwiv41MNyxwnCM8z0yrV+hdd10rJ6413TdDCtKuqB
U8QrdXMzUjDesIk6xDhjFCMKHF87PrLzBD3ww8R5eEQ7GP+8R9MN2gG98Ztl07lg
PCouJNCFVG2EeUBTbnn7jHClBoSu9fOf1vClRs9rHCNpb0RtISxBtlbOy7xOsPZ+
3UC/Bl6xwJrOEPcgUonciB8C9zl6COUFCD82hGkmEXysUsKHIocX1IVHpQmSahZH
L85zt8NfHfV3B9nYy62iPiDeu22Glg61ovyrqd1qzA+9gMZ9WHU+xsisJBfoS/gX
7s1OSI75RGUWAcc9y/aUMALxAOk5evHBoikqYGQM5SXS09cwxZoyVfU02Ephe+2r
9CXHAaz7Zd7L18lo45b06WVp7mHmMkHRTSxWCzqT8HdWXwr+cAz/ZxQ0UARTpwpd
yq133q+ONuX2cqH9ruckxCVh3iWOXFs7zMbGx/EUGdF0w0qkdyMl1x4RtEsuXF63
xKIhKJsosIqhWi6ylglKPZIwhejWB3PQCsZ8b2FVXvPs78ttb3kfbnQ2icoaj3m9
akeTceRdXqOshMtVTu1YqW6sV/ong082oE2wHwmPbuCnbyeIlYL5LCA9udOhXu0F
6KDWvv5znNnNYo/fPeLWriwIrUKw/y8pgDECR8IHNWS2QzZcfwqc15n0DMipmLkr
pljUXbOmOcAgCGUgD+7ciwJNuFlpPfpCJxUAbA6vgaTztfthrzsTSFTtp7ZpFhkP
CnuHqCNnXfAS57OxhX9oWdI54Pxr51p9Ykf4cMvlIDzh24lqy4SJfoNBqu10vcuX
3uPNqs4CvPssLBmVC85//63Bu9Ebjzr9G5szVg/e2IUQf9dNsK8AFTdReV3KdwRH
GSee1n17C4tqq12yTK11AGWo/5538rOvUsJvefEsoDXfSDEvAe2jzVnJslVZNcMZ
c1JLATMo6lctR1UKdNihcu1JuYQBQ+00TTAVHN3lLrJZ9PID1sAKpwag+XEBh5Nk
herD2pW1mcmjeclhiSNP4tw/bA4nzJt9XIvpfWXHt4/Ft/pQui94ifVxl/xxaTnw
c7pX6xArxwn9ECLYAsOa7IttqTK74nBFFQpi46Jb93DHF60ojjxIiJQmyqkMtS4d
o6eQPKYE+Qtp51aVZnYn/cwkvrPzKhv0MtgqDVbsi0a9MORNZ4XliX/jPVlbDHVz
IfvcRbhZKNRJy3oKTtO0mh+tg+UwZ/4yR6FMZgMK/GP8uYc87AYH//5UE9tT6JX1
AZvs/VnKR90914LgxbEmVZ5o7hL6JkJlUfKcshdrtYlH56DOAyje8pxBrGq3oQ0l
ddwVVVioovyog2YdOwv6cyBo60qCJM/yZN9dO/CpgwIJLYphgRwk36cCnLu1i5aH
UPMgiz+mIv7ncZ52FyeVtEGCJKNAPIidQPohG1W5rOWub923XpRxEmRLgcO14dXx
HgjdbUegCGHJRGC0g63KG2tnIZ/E3taDS3jECwbw5JKxbPLEEpNOM0B20SNZSENe
Sh+ltZR2ChsZ/cxGiNxBbXbxohIvuuJu427wkUVx1U4lDSql0NR/thFTd5w777hX
SqF+iYfVF7g36FMC3ZXkF/mXVw2Bxbw9MJzsQTdySk6GbYOTGWz1McVgW+/ib8uH
Qz2OtYCdGLsoAgPnd6mn6TYrdaj7xc+Jiq42xJLHlTTZ9y2tu8fDIvMgeWVxV/0x
iNyjBTGVNVFOVG2QvxN5hNKN/JaOKqcS1MkMbC8JlpH9fGs782cPZcJEubfoTQFc
RpjLdpR4/Y57qwaN+C9SFQKM6EwY39FCHOdLfzcZyUFARJpn2tnyibyYtr9Iy4Al
UTTnNgAnKagzXGpTKHAhvnuYdsJzGoSaJaeqin4jeSxO7Ls5BRJccxa5sMazWKxH
qcCvsCPcpQjXxiGiIfCu5d2Bbj07PToxvBlJQRADntdTp6IciShhRtsN+SAauBpA
IqpoGG9j1sYJpp+FrJNYI9aKOKv334+pr2eqLWZ7tkqC+I6uz+0YeiZEybJQY8UE
s0cvH1Vb/eJ0eM3/fgefvhX6sRpup6Ean1XI9yg3YFFDBkiEiDAzJpizrGGWQDfy
nHiQVHd7EVl++w1Xr0bYPVSsaXLEuo0n6qUhTp+mfM0tCCIRDpWgcsh8kko3mthk
HBzjosH6UmG0S2gSQxMB42ckyzWUfS1WU7zxjxHTiqH+9RzNvvECAIWrs9NQdIig
FIahHKHQ/8qGAJ0cq+qqxKhqRrMk57pA5l8e5r9Q2k4bcTBdb6gmKm5mZetU0cYg
zRaK7j8NoAszHCPazBucsQXwgE1eOuCMJlnaP6h41yCumh/om9Xt/c/6NTRf/qr6
ayogzFKOIfl3JjkP69t+sPQV+NxHlsO7XWqTjlnlQucT7Hh43Jt5RS8nwDoSwFnY
1Rtgcgr1X1TM0gNRtOslTFxRETVkHDQ55QCNWXHKwGKZiZh9CsctW5pJfRuZy9Wv
hBYmbUCr+oGnuTRsc2RrOilFvwdYnwOWuE/qXlhvXPlM9tbZKgoYxMnQZ4eJNZY3
NNlOdeUGz7R2+LJi+hPhhqq/pMirZfDIQP6/7iJFRaXmcjOCJyOuwsjHX2LNs6mO
feHoAsU6lTUl5GNrqxHNHSvUjXdrW0ZaZmccSPG763I3zG8unkv4LnX3gFYE4BJP
0vO6LExTDeFgx5ZRuUk744wfuhyf71HUVJP4915tLPRIK/27Oy7JHU46CoLYuRLN
L6rmtZAzCCAUwgCtEME4xK1pmo72VrnKtIiW85mbxelzpDG5klu0RBtBEQab4+vs
/8Z2cFKkCyzMb+BE0DMg2dbmtu0UQ98WQeNc6MhfUhuUn+PP2t0JRDtH2eq7KLkx
qJ/0vNFy/Xx6Zlo5CGSEdcMRzglEB7sLdspzSbO4dBKrLk44u+xqtYwJBS26UCbc
2jYLXzirVailo/jP/2LZ/POHouxBqdSM2pIyJ2U+kxoQFJUX/RIdmCUhS5WJ91Cv
58k4R8YXkldKryV33Wit97sBYnWzzjAydndQ6LBjNjliWtStPvbpSq68xV/KUriX
rK1aQPIN5c1qZuVAjcwapH0+f4v46tq2fzPNPHg5S9bGD+5JL8Z8Q86v4668Ma2s
POiJxA0cfSGHp9ailPb85MkVUpCKY4RCeKDOPTiPkYV3Ab0/rC+Src+bZjFqdGee
8cQA3ytUguvggimYYQGyad8gFnRjkrBfiGS9LElLaVqpyDpqc1wuxl+LZO9oE4WJ
Xai/wdEH8vyClvmf3cActQXpsIfHqtFIwRLX9+v3QxVh0cjvJWkPhM3GFH9vf0rR
H5t51zxxbc35yn5k4a4FjzWO49EONl9H4ifPEaWjNaU8TuMsKIoSduIqbI93q+6B
hdjX72p9fwwyVieae5xU4OYNbtDgasXBxE626mezBkaqbNZbBKzEbSaKleOAE6WC
MUTMOqL55jf95C0qUmU2YaAmXl7osNuIfHgn/JAoBUbcR8HRN8JqHa92Ihvk55fV
K7k6pwI/V/ZQ1omrgOta+pbCa1Ex8xZ8QduI3K4I7BsVONzdp5frA1DB0dnwEhKY
SBn5rcT3e2gj7CJOZWGPI8xoAi5kRuaxFrrRjhgi+6yd5z6S+YewRVSfK6dZgaQc
EtLFU+IC3E/xOOXpd8d3H4/7mKCsVpcLa3FTeEJF96cp7qcKoeHr3+R+Z8ifkakA
c6pO38kk5pHRhKwhWd9scQzfm0oMLjyL/U8nC+vEZwgHOYhpXw2pqQJfcv4G++N5
B9EEv3kfWfP7VTNl2D1hq+RP5L8Dm42lAC8WeccNJyZKEAuaTOOxig/nGfSd2QgO
1f/Kj7eRenjZHXj4PnCCKLiMLXMW2ZpamQPgTmbLSSwBBN1g83WlFDnXclLzZLfz
RVMw9nwePNdexZ5kIlBpcz064E64d33+loQms8/J8xnKm4mslJ3lZS/3S3+KDZAm
fokU77dOanWyeo/VHrr3qGcpWSnCf2quMgnaPlhsv0SJ1gpcMxCJetxrmj3OZIKt
rSQDOImpWRBvoYKfT129S48fakzStoNkDx2ehjE1cEkpj2SwqhMLxNcoFgH0+QF9
S5xvL4sFdpckYLez8PTz09XJtCsWcHjGLHMD7bjT0F3Out0Ek8kq/rtJ2fWkXBDA
1+nknKy2lhBFEbhDAYBdrRDvLX+Jz1HgVQJneWfkcKehV2KuPHeRui6IJARnKgBX
oj/0PNX7VfGI47y560VPqIc7OaW/lT6LDGETYxJ7BYT/ficP5tP3G5xsGyM5I99Q
AvZyBfBqxPoMKqh5WnUwtpx3+0r/tib912tvwp7fC+VAlbqJcBzaLQSiILcyNvIt
hk4F5IxtcPwMFrSMiZYU6zGIk6f9uyDM9Adn5uNB+pb2TaKkCiq9HHvO6cye6M0W
NTXcZYxmiXLDLYjdsWYmctT8l3AB/O3ZzEx7qTmE5rBnWTcd7kBEspT2GayMm3LQ
IoToGxTJtX/JQDGGrDnTd9B4/qunk+OwzlQnlFR99vY4ko2iCiSMe1OzwST2weG0
+VK1Wz4XsC6LQvltiJ1LFap8WM3PNZaWlzZsQT9FBx6OR9AT357ZXnyXu6YnLNHW
ZjGdEOgpejbPKK6ew63j0NiFLdEzDbq+DWlQFhZr/vw9/tRwKvgjQWAwk8io4BQw
9yso0UpKAjm9KQYm0zva6pl6xP3zpzccxD/2QMFgWrspsPJP5GFgp31Sh4bS5F3m
uS0LPU2IpVoksoyy99GWiSFu4rikC03e866+D+omCovD257equHVEj8S3bxyeM37
lGkCTTQS/GIkVCNxpEAxQJpT7z3OSzoZZ97+ICpxZKfWGewRvqUhMOXBrRfvlR3+
1XDRwOjzbmLKKAJFuC7jY9tbmyKjlUHwIIWpQiQ2uiRZFL0l1bpjowT57T03tQyl
7vPnbTI3+rR4HCL2DBXlvFnPvSu8l4PpImg91jJse3vS5TOsAjDTk9/XEh0Y69h9
+LsSeSVC4PD0wXWZ/p3jZf0y6bXaZvticir51+v1aq8674BUbutivWCAWKQIHd/s
ITSwyXSKLuGjr9Es4otER7/0tFsjonlJJXS8WiMU06sEOpoILY1EYwFzOIH1/IJ1
XJf6IDUpN82JesO8hcrTPuAOkgAUIpDzn+7u2nLaOzwaVzkU27IDnJ6CQh0hYe1/
7xGA7IiDZGJzPAuvSSNKszHCCBLf1ID+FgRkqyxdMvcHiSpEA7l+/8z0QVh/OB2H
rIN27tEV5AKucVoHggl6QQq32HmU6WcebZZnR/S0jYAWm4Ti3KcIOWnt7lHpKJTB
OOtjn6IcFNK0riKIv523hS9qYlKhnp7o10GqouD9AlY986pvTASjcWDFNdsvdNOs
uhBbeoVkZr4otXog8qTR408poymEmr6HtPESclwKvqK96OKaoOojt9w0EP4hQvdp
GrWlNHx1t2SOZHRlap95cituRVHqfv+6aV4n5yq11j2MRM0GDAplugGbOw4VHRTG
cxaF/aiHjA/km39EsvsUS83aK/TAsdpSMKdImiXyaPhkZL4vI0MxRY9/sD188h32
/qkK/HHEDnoztvwou4JbMZvhSuz/FgK4rbk587JoWhYFj62B2VdBh9uKGvQ+IFDf
R2dJmsPhbqJ7Pv2sWrpxL1zv8P3iZj/qMdpP10PpI/66L7hfDLRBcrmwORjwBI6e
NVj283Ikr+3ivOW980Kk77GiXcOWZioG8gVS09HVLJNDAPONjSWF6YJpUUkN8qed
snAh838ODBCvX4ljB4yHnA/NJxYQFpD2Sq2oesY8+L5KEzPlcZcWUVBBwk023h0J
GK66UuCFI+I44dkVr71jKUgcTQvC6odwKxv2Uv9y3dPJVA9ZgYc64TcL9YcOM++Z
Kp43sIKnyVASOq7kpaWefvzhAXQyXeRoMQIhJzUiG8yrw2p1tBY9MDgjW5pqZvrM
VTVLlmBQo/tfrtOqzKYYTAzIACHtOahbc/DCXGKQaqhox+T+WFjlLlqxSdJFT3UV
m6swONbZVQP3bVBmH1X9xZdjKKkdOqe+/bo0zEMLJryY5jvwFmvsTKRRQM5NPKhU
6TjMrodmiqne7o5QwyCQ3SLPALNyvO2yARROEH/5uHWH0MyZDqP2AOZW02xl+ZeC
vQ/cEZ7cSWZNRBpmIzNAIp2QlH6THcnlfvghGisAqpDU9g9EIx3gkW72m+LzCkwK
V3eGbLxpNDZE6i+M4XyVbkVmNoiIfywUWsHImbf4ZvsEpUX6Z3b7dKU1ixZPPWT8
bFStjLVHQYIY3k9qKAVer5G/SF98s7uWFx9zm7dNv6IsqdFpg85NqYvciBMoaxnn
B8f2oT+lo2VA2bfPcWkaOkHYdwG74FdDpuKilq1OnmuXVoedteMrN9KEMJEeb39i
ghju0j1BoKvjfBK4UW+zjvsxciWDQL1keTrNBXBtYUE7dj9jnoQ4pYOnKAmtn6zf
luGZscmrUBOMCP8HspeI1kygYXLfR79hPNhbEfIoKMyGS/v6NLY3AJpDJuBcBxK9
UoOM4Tyf6FP32LqWwTed7TmK7yK2vi9m5rSwXJ12BUB7iODc2FGuaUGhnQHFLZKm
4VYKeZuoMJo9CvPn2T5JME4+U4m/wmo7kDvHY5HgCx5ZDmHGUH6UeAL82VkfTV9M
0W8UO3857+n3gOhZDl7ReLc+eSNwpWJfg/xYObw92fCRDU66DuJRC5i1avTFV+DC
bcESs5hlC/+ErBRvmelKk9kFx0OB0v45QW0Hqkd34yWYFOCRwDgyr0quyjrdkCEB
m1Vm5YxAe1xVllgqqivsnYXN5RoQjDPmXqpKszSA7tv/lOt3FrXCcuqXAtbS1CjE
r7YgW+/hND2vVkGoDigU+ysHuweO3Bd0nehRSqe5AntpwuZh6zlJKunynj0hB5bt
wlUYAWs6J7/D5hS4fUYpmfANZZFH3QQ6amzGZHkmbHs4Am/nQPo0u5W8abxWDzS3
SsW+5npgXB+eN9aUaWrLkLD0lMEsKUqsTmMuU8Ja7pkHr8o7DT9K0D6BPB+63nSz
RpayZdb6CNjzSrVfmu6Ga573U48bfBRJgFJLDmLKqOlTtwwnJzygemqrawH2Lmmz
MbtC85zjCozfRamF8HWTU8TPjIx5EWC4XP4ME1M/iw43zsKg/F8vrChqFGolS+ok
oJ+p0OcmD3B97cQZVb0bkMfpEovz25K06k1SY9UZnvtDzB9UdZ5mIwqJMWn7X47w
/dwk7Cd1hbkqAQGn38sxQTlBrsg8Wqw1TzHjUZF/HlfF4Be5tYieMpnT6Zj+1qCf
XRtWJB2YhCPEYoa1Y/wotOXh4V71DX+PKZkLGUTQ7OfhCqVfp6GFHSPxD6Vrob34
Q82+ydHvMCGB3Jm9BhhX/JOU6QB27S1crefbdq4xlGvt8HINXKu6Pu9M4kpuL/NM
gsRm34gBjy3708OCzVboqhLMJe1mmKsdP6QO4Uyt5qB1MJyXz+ueSJS94f2gLLit
KYCtQA0sMqqa9uPKWGRG5b7pYv8guOSYw5CuWosUm3NTUz0gw7Oc0QrzHEyeBFwR
DZUVzCth4s3N3Cm6QJsYX+DN4/SlgaHpLAqXyk5EfAJiV/pTY0Njpu7bviZAp0/2
5grx2udpWKZcQVgKnRTVuMtxoZ1kF0drrt5r/l2pPP9RYlQ/zMD5DiJ+siPMWBvb
N8lsPCPq1OQEegOx0e7X+KVUGJH9z4RvWtMA8CWRiBpR8q48KZtZlpazABiclwRg
l8i4HiXKrt9EoB5gzFKSCa2X4PvdJfpHIlFtSkQVYN4cjbDcKA2isoarozoaZX8X
pU126ee4aLaDy1dQYu3djklzLeTDtfT/iY1uPMZxwBoeho0O0ymaPuY9U7ypoImg
oEds/VOwWdBJ7F74gV8XwLrjVEcTd1MSxqvU5Eu098SlU9Av7/2GSSobm8pr6nS+
hOil0mFzzS52GPvi1+2u82ZzeKhKtDCriOWbzFU5xtvnccCdq5VEQ8DEJNIgItB5
yeVI+gSgLxmTZZXEEuy7hundVEIRrsyNUWFkDgvKLvn5qoCLUw22kfHlZcxc3dPn
dIh3tdpoZRmtmsf0PDGqV6TqfifvLdFGCo+W8jGgoD7KWbL+TYZK11igDZ00svU9
YY7a9mFcEaKs6Hj0VtM99J69SzkSxH9Qzd1bP0ojhQOS7hKF0OhpMlKOOCpmpRry
9QhiPJLySi57XfuiUWgjXOy6z9Ej1Dwby+H7I69IUG2pycc8YIEbB16gJpsGKnRz
mISTY40Y+KsUBxJuLjzQpGOOPSMZPBCnWv7dEqr/Bi1YzI5DTFsf8uHHf7e2WNZD
vkp2u3rdCDXMhg7btuey/S1RIy95Ou8ii/eskNOlNkoCMv6vHIDnYRJELmGHchcI
wrjKw3qITqgNQx0OdvdGAGBZjKaUUfvJbqep8UVpus0sEJAY2OwXIODXn872o73G
fU/wEH/m94zcedNiiYPlclFy0Z9TN/BHtbUi3h3zdLnBqhyCnrZ9xPNmcF5vCwXC
8wr0AjvKotpFzzzwTHqrhJ6GhyhERkk3Mla84W4t3Aw8xb7MZp8+3IVPS2rLy5MW
k8rLVDinlaNdgZRqY+E2sUu6gYLEemAsBU03MWp+S9xzSmMWAI1WLZfkSyYbmW02
Ff3ydInaBluZUBmXtGT8XrWwrsQHBHogW2JfPWNIp4dPbvhLbhuxNujSEgdZsbDi
faCv51Y/LR6ExsqV5wf6GEUuCvh3koQFrMl5FfL1S++GaYw6MWoMQORIV/1KrcO9
VECUu9qQhPfC2npryMGX9T4ugv2fUIPInWTIPAbAZU+vi9iGjvJfy706esSOsB+7
Kc/OKmrIAz78xX5oOyOO984l68noVSRvsZyh/QbMeW4KbVELReSqb02R0pzs73xM
z30TEAOtqAFuqF/u9qdpX4E4zzzp31CG4fHyEtsSxe3Vf7vfKD5jtxErDFxxz/lj
cAcYVqKA8Mit0NxusZ42atVHigY8VXsnl+IaHQ6hTW0xjy0T3lMJ56FEsvNvHuk7
g4HyoSpsYdDvCSU9+5zRz/ruJa8oKmeL1Mc2T7tEP69hL9f7ieaBTiuZBQQvQKSs
f303ih1DxYvIOjEAu5+cSezQsRvwRSEJ9YYkEa4EDXwzViS6I9gN9MTkox/ghkyc
8qDX6UWZeWGt8AEnn7AXgdGh7b4MzrBeTpSD4QelyqtEbHoArtnBsRva3PsgmBEF
URxY8IhJFgZ+NE8MgM3agt6bByNIQqZZOkSjeyWalelXixQtStHW1BPUNh4Of7uw
s6wIRu6zHokUWX+8lDqhW1M1vdjT/gOzKIxqreZWvw9P4YGae/dNwERqa7gWkLKm
WCmLWCTTROuFG3MMFbwW0SqoMn9WStjun24t5NPQEZJusC2USRib25Xcj9JU8DXN
nTHvKw9/G7t72LIImipOuZMmNQKqVlRLQY5lU93L+P4n1KC0SgvI/UdIx1lugrTk
S9l35xJwfpfNJQRXhzJ2n8ccLGDSaewHwZuB7hU171bcxS14R1PKnsO3XFwiPuwg
ydsag3Os7zerZVQkA6H39s3Ud8CYZj/1NnHcb2k97v7OSkJHL6L5TjW1cro5Ym5D
ThTcv/1axRJkJikGVFQGyHZW0gH8Uzr9cFyq23JmIu9lnaPESCpq7GIN3mjDo9yX
FT24Y1+4UXfo4IgemzhlYbEn+GwsJ/50d+WzIsNicSFCCVFQV2N0PjbbNntRJdcq
8iQ2jDWElnVOLK6maUK3L8aiRqY/ErzvEvyh/XaSJqk4YZaU7v1rGjWtimqTl39v
4Ku3cbyT2aZF2FRWouWLSl5q4648cc1QNXcOZ6mCV71++y9N15lmtLfbIejj9tRh
8KN2WxKzqIaFazYAhCM/JT/cPUucWYKI+Y6QS10e0+IGpO4ZEb2Ztc5nH84ymVGr
J5QBjY5La0EI14ScYN6Ox6D6c4GljRKt8Yr4+F8dn9lXE2u3FwJUXFheQPtet7Ju
uxg6vcuHWC4DC6U2PjtxDnHeWaR7ujqUmOL7Rf927cV81EyYee69lI1wlBRKaEjt
RVPxLCOXwMCoHwHuG2CKBYyYiYYt68xkeb16t0EgJroCJuQseNwBmydJFMsU44os
9K/13SQ3g8yVmFZ30b4qZ9Cy4im4MKf7Deg2np+IeLc9EnmXpMzIbmrAFv8ihko9
Z0r9mJhwaE745PSq4vcy69S4VfR5WDOEockNKObdlTxNSZ1IqvE21SFyvvkceRkW
Ib8Kmq34QGpWDzVf4E9qJPqZy4q92SMxLpmQfFhwvGhGB+l4nX/v7o7lPJ0wwNkm
eAcFIthWOT12dNQb3vUipsfDenDDHTMvbYX8PBGBzRbkx8VPpeQw/QI7EtpniTWy
JmPO+QIyUJu+fP1lBPCWA0B/dZu8IcgrT6bGi06QR5XduiXTHT9l+Dh6S2IqWckC
MeqLwfd6vSUgbWxhUMF3QvCZCWJsVWGoaf+lvPYGxgyW+BTHoA6EcPvkm+ZSvtXl
25d1zXgnjF+G+VFkCqhHwIz0Fhxt6oYoYIwYZxBnXg7QCaizo5oNZkhEcgXyIrQy
6u/BUFiT6GF02uOoclIcErYDueY5BRQMNcA2ZURsDGNohYdb7eH03ANm7lHn0lhf
E0dJ48+IeTmV8D+cMObEF8DcUZ39kK+T3kkZWtFsc8VkjoEICFDRzxNRRMP8M3w4
vwjE083Mqd5/DI9WlsOP+nDXUaZeJ61+EruSor652V9WwrdsGv3Dg07wcjEJuV+1
3oNgJH8zOelVleXNNvp4nxvzUMJ6mZs8kA/DPxvqOSdTM+WRWlje31jjZeww8J27
JZSLiBhdy9fImM0hCAHYu9yuEIMuKOAghNjyOJ2s07XpqQOdfnD2Hc2GYr4nC/R+
KWRnRyfyi8ew3QVh9pUdr3/iteBANcQcSD7SeHVmqPd4IrFYm2Ssh3xqOAaeNysC
9hrCSKDOD9hah77BUTez86bYUWB/cSG5gubapovuUkLo+W/QEqh/ldosEgA9eoI5
VIANRwDe8kujojRc/k958lWv5ggmoOuUbJFx6jQS6E0YRrwrGLoA00llm98XGT6z
z1bAOEI+PzPz9mG9cmP/Fg1esiLpgVEBvF/ssLUmO8DGXKk9Q9mxpMfeJhqCHhOc
TzRpWQ5xFaNaT7NKYUBe2b4zEYbREV1MiPWgPKqHK06Ias7yNe644Z3RzQpuSEjD
567k24JMvEFuFimWn9mz93k/dHpLPDSoXteMCkMUUlWfr7vXEVWvsusAtqiFeEui
tXx6ldGhtM317x8mnCW16peA4JWN4aW0JZbKOmI0gIRtkc0/dLGVzwgGEljv65xp
6VDjwVkKes1NatdaBmNwFQ1A4zHS4tbV433gkGi04FAqJW9jPeG7ruKV5xjqWdnK
m2i//iOPRrxxaAj7f1h79KEc3vOoy6j1j3ISJ8Q0HRfkTkAHmjFx2he7IMQm7Cgy
q7thYwfflOIzzbCibCBz51nBeTOgGilb+UxebSgOsQeyinE1gycAseG1S/qLcJoO
+cAI1qf10wt3/98Q9Q1+z2FXWFlzuilprxqI8gia7PYZNAcLmbTXNgcZVzl4SdR/
JSv/zDFO7DyGp8Bjirl/R8KPZjbaW0URe8IqLp0wiz4XL4x5nKltrn4LLSAaO+x+
DCvSQuucDIjeZlvSqduGwsQ48q9Wrw+WqjtBI0xGbZtxJB3maIv3vFFLU+hFDSre
mBkRoFOv8Qb2O5IxYq54+Qu96OjYK8VIPhGq8JbGXH1XFK0kykKHjJxdTf4oK9/v
bTAqA7bHFtgvWboggRekv8OpL5pznscnunhFpJjQ8iWdYfvDo1Qzpk3VW8npzkMw
Qnr0voWKSuMjZAhpTO2oDcHZ41xlHu22Zoka2A+sZ0pATfQaPP7FHxG4AbsPK2Wm
gx1cXAw4mnztv+gaua9xdMpAbQL7pZfQpelKx3WGkW0j7k9YOwwLAuZmhtxSzMdS
xA1jqT2g/vioHNBBJsv3O3hwWAy82cz7wOqBo9dgXj0QIjKFuTqNjOxOg2qvKKsM
x6QkIxAmSQ1YLAWm9pCuBe+wAJ5HY3vwWd6UU3O4Yxk9J4QU/aTltRhraqX0c5Pd
QuaSGAdUjaamIduwLOBzzGLeQX6lGyLyzZvH/PvC1AqmZUsiJu2i4S8O7JaLHj63
U1Rd4zLIuHeD49wqnP7U9YXFG8VsyApv8pkVu9IoETxh2axFFP/fJC5UHPb/wIjR
Gf873qBgfTY2nOEugJWlbAAnpxIPg8SCXVDVBSOzgc/q9XefF8RT3OqRF+xOzQ5o
OR/vjY8IcER5R0pVw4QU6ZtBnz1Nuh1I0Ad7BVJi5CweFtruci3qRSRRfl25L+Nr
WU6cqAg7F7vwIRsH8RIKBkYLeY+cn2UVlhCZe5AhSYQGmGLE9ZeGECHWGxV2gYmZ
DsHjmZ/wc5lRQQnNLrpUr5HdCrhRbnsfS8Kxku0k2VFT977dGXRT+ROtzrtcW5Wb
NDxusw8NgpzhoYDtz2tnMYgr6P9UdSenvR9nSMLRA2i0v1t7E+5VWRQUkugr4iBQ
JVqGnDk/V1Rvj+L2486V+VhA9vza5W0dGWoGLCSNmydRLfVFBtMkAO7Zk4lf9W/N
8+fS7F/lCEH3ErEwtNeM9zJcB1khrvN/gbm99CPxZ+IVrDu0TBzDtY5dTrINTfKn
fwDW1Rcm6AlL99GFYdWpk+5Hc0h1qlIp6tORw/Yb0hWdXn+QWepSnaqIlIJRxuFs
7JGID1yD7pjL928OAbypEyRfjw2hTNarYPKlk/C8eb4iXDMlCnbiXdDJhzZGtdWo
O8mtbLaSBVVHhkCI3rX66RXPIclSx6aU3mhUK9VvSgQprLlA69tSdyoKOSo7InxM
oPKlXZbWKC5TL58yCaI5eXAPQcPTnsCKX8zDOZvJe4tYKoy1XZGfIvhU2JObGtHU
qM/xiX6c3obSHt88CSR16LKmEKMix7lhlrNcCtoTLQondlylg6etB18v/4maLzxu
AYO9fgrRlW1TqDQpTGjunZi0XQ3ZCh0wmWz5nSfvvrdUlUeZwzIYtHu2X2e+NtdH
KeVrpCyHLNJij3icVv8ey8jr0hp49ZSyvKmaGT2DsxTYfs/9ZECSNhusURTVHBWT
4z4mKwRHtW8x4bBy2+ZkW0QmiMHGf2PFGvORvFzjAsOv8GNt7X8JGyAeVGblu13M
SVqLAjIDHJg3ew3So3SyHS0ibH5nfE5dfQlLO52fl7pQUL7cKjf/debVlV0yOFpM
8waNbGqbtwVfxlu1hD+o9Kp6mti2HsBxi/CPxlYmvx+0qEXbA2AkLimWXnjpZwy4
1T0vrZkxRGQJvSo4cmBXsudMZPx/+jjKXm83JKUVEnin6dYN5jOWi4Xx/l8Q3MU/
YNUf3wnxRLK6tgbU2irHRUsXSPZ6Cmmu2msXK9mLC8+tqyxkjrr+0FZm3ybGpA/h
N2jo4N/qvlII/SDjfPuGjMgO3KpLQwKFc1qSUL3381qnDRbeXTKLFVYkpVMAttbR
4h7Die3UC/tzExYyiTxnCKNTiCeK7QYstkZS7f21AKi6UTS6PEhk1EsuoD5sBwhd
xSjRwmb1iCDUt9+pW5nuLyG1R0P/emQtSy0K7n2W3QlxOrDmwWjVueXX/B8FRowV
PGMcITDyuHFMkrDErSs8Z5xDxr5no4n8FILIe+WMBiIoh5d46f8N5BLR8F5TGiu0
J1uDxP4lf+zNtzkb/0vOGaBXP7krbcVb47++/unDtwa0yUQgoOjWW5IklFO+E/nq
n+o/RQUBPgCwL5fr2fbaJUeVGF0qPpGBMTuLP5MrkYCOphZkugYXdzsL3FKxUOzJ
W1C2hAYXk1m5WJU3MT6Q1IJsg3/0W5Aw1R9H3qEjFjDEwcugCyT0LDBaxWCFEpGt
Bz7in1xbTro1oaE2u5xXc19lDktohNawHQWkH/qzWQ4anJXo+T5wW00+crzQjzaT
yL6Rj69muWWSaWPQMsYa+fcje32M6B+RExk7SM5o0ePcy+bKipOwS9FYsyhUjqS1
mewyTCa+srup5pLn3DQsZEA6R4AAwZr6xw55/jVSSkI7dyS5WxvjMNR/25z3Lvb7
SWsrGyMTl19lh47q5cINvRrH3PvdpnT1OAG7pwbhMcdjN2C2WM7fjjnyYeIQ6Yvr
sibcDkcxslvsVmqUY6PDraG1kzkcP0pKneQPHkCZ+jiK8DkO0UVaOyZ92xY+2Iae
AD6k4d/dqcCG8TXe2cbY/7TA2xOOFcqu14eikpRY9MMv0YOsQjhre9TncpBEVoAP
U5OTh5XBc97Iev0O4QawDErv+l2omqwDn2eyBZg6fDlIksh5uHPRjNNDhIrDDXb/
sxMuCykaQx0gjauCdQKXDdghIKhGzB1GfjWSYF+4jfo6ZgC84KI6BF9HoOzRjWZO
8e5lhpXJLYACxxRZZqpQuew1wel2yRXVCK4WtZ6tnuZMvo0O4DwYXGdFzXzwxju1
NdbloFdn53o7lrhwB0YDSi04JmzcJYXKROrBEQSaJtXT5EYUDFYzQAR4UMHIFuhM
ffgkuLWilcV7+5XBpA6IrPf5ALDTDqa9DWXNATTcKG7qINc86TfUd5Yd7R23IZhf
gemQzzHsY6sP7RNTSl0iIxfh5aR7oAvPqMouLaKgZ+zj2W9IINvundcugGDaRm9e
TLkZ7EAn/kmKYzFJDOKpKuNnlowaC4YWPxETpxnZlSbzIMX54cJ39XdNBEOr/Eh+
ihkPjvccz7KKo+VQZch+Dp7tSObNdvHAtVojD0u0iGaVTFlmZBdp5yQ3vP+L7/U0
moAT9u+vuxrmIhUAmai/Dy61uT2YbyA5awWj5vX7hEOCxc8Qjzlti1t/Do0VsN4n
9aUs3n/drvHC/9jc0Zssia/pmMMJvRcaukhFZG/x+ygSy1CeKZ24Vu4MbR4Gfa2i
tawwdJwQG3NQdh4W45pJWuLUi9oEMQw75GnandWOact5SFGlOxd1ES4dnLydAzCC
IB5+dQbbMiCaPtO7bedDGNr9DPnZiQxTmI45Ej2+sBtlCe7WFoYbUwMTAJDzSt9K
g6xG/wV8sgWV1/X0oauacePu4g6knRl0hW/2bC8hTxocCOTiYAavVX7ZLSPS/T2T
3WOVZJrA2LMTVjTA7IGr20tDEo5uE6GW6F29OeP3wxYj5Ktrp+O5Gvi9nrgeHOOh
7NZSanNS3M+da+QbqPbUhfJlcSr2CKYpDuTgicraYzAGovsFWFpyUK6sF4+yyxzg
pDTV/N0fCEchd5tOndm4ZUCgVCBif5v/YsgDAjHwHlryT1LWha1+pIVOJS2HtpEq
QLd3/KHmW8Qg/0zpae6EXAm4lb1Qzqa0bdnCL++iZRMt+GNDMAqg06Y+GfMWGoRL
c+vn/sN0shjLhP+NczpiSkrRj3EKEgKuZGfy5VekxIme1tQGvf+FC5r+2trK5P7m
nviQo5I/FB1kfeW8WlpC/lcRT6wIr6jsHkvDVvfJzHAv9gvv+xH+E84XBzjKy6cd
7zYYJH/0/RwyqYQv3U1zYLbZEp+ZkUD61Xk7kWbiu6TY7epDzsftPdH0c5kQGbXy
I3HcXesoDR839/6MG22BXdI7I29uYrlfW3GEwrqKt38m9GLvhlbPDy8f1+uxTCuW
y9oLFBqIq7UfszaV947Mz1ZxXgsDInc1nwC6utrrIwhTL7sBMg8dGhNiKSwNwVCH
cgqjBZ7cOopb3/ieHp0T7w5U8GiPEZCUl78KWFuSDNnmK+hZl7QeRyljkZMqtuuI
L7EARf9ZQ2r/xk5F3R/wxlk7qvgWDlp6oW2Slk2ui96o4RZfHeqcWAETCrf6eedb
+TMdm9+2myMz9B/FIV9sQDQv1jlRbf3fUssbuDyOHjzdWR8w5x4e6uUCmEtuZkc2
dX6GEvGJBSQ0LWI0hDTY6Df0OvsOWIa+nuMDRBmwwX8nux5065Pp+TltlxYEr2UG
S/UqtVtQgX2nc8s20x9op7amL/f+1VfgoyWa/Tduvl3rrIhzGsZG6Yvgw/sVTQiJ
5p02PDUmv6p+ZzLRLbsEHfQvUdK94cyTnkAdgxTGvVbGHPciGGIKd1FWIVsHM7QE
78Vj8+IwmJb5QM1BVt4cHZM+/9vhLh5lXex/P6whErJAIU6r3Hj6Snw4KvyqqE9u
xCBlRuxLX+1W98zVsA3s7LS9Ipt88mksVZD2tsoiXm1p14e7sVeFFgDNYG/R+rKg
nhciEpprUv6f3JIHb0D4aE+GhmYH6T1z1VJfdTMRQLQDnBcbfuZhjRyv8f2gzQRb
5DFutcVWJiCtS9FjfN501zvlpUqD4gxG4fepqtp+5JUJA6Vn0L6+fZeBcVMK4xQj
SsHTp2BiUIkf9fOuMOuoNguIs7A7/k6ibb6zgdeaKXvAyoYFvoBAZnlosGDGVRVS
+YYUhZq5mU0feJ7fI6Z6gRaKKM5BEoXu4DZfkuMXRJOuOp6cMquQMib249XGguh6
bbOr/oQYEU1CbXqQO6LUVf/tcLwCBdQoTgQT/L2nY3pPszBkh1vqY1h75EViWRzU
adQZ8l4BwXqYAO932haI9LJ0q9pFnuECKK9fSsy5uyqXPabBTt1spZb2wJjRY8iz
zg5Xm99jhED8Od/VP6xERUbwOvfivdKFOdFQDqvH4RRWUZIMO3OPLmTea4u1aCBB
0ORXU0Ql7276vfRWHckhLn+/P8BI4IJClfoRYFhP/j7xscOnwhesP1KYCsslV58A
TjJsWaxT9j/4gbn0DBc+S3ZHBnET3B6mTMMGfv3zrNoc/ZDnqLy/Gv66oRMkBYm4
oJCnaQNQMIJV4Ghe+Dpv4+J7UKik/u3xUoQ15pivlon/2cUF4NSJn1RF+iv6URXg
UVkJ5GcOBVbPmSsv/eH40MGMrsvBuUL9Ap9ePn+qyzmLKP9fSrJF6hCI9lVbVfF2
CJvMff5bzGBgQFRVuuh7rlyerEc9bwezMv0zHktPICT0XuXTdetjmV+4IoULGNXf
ho7DYScpCky5cc4BcN7xY5J7bzvpaLkruWhiNzqrsVUC3oLpgxn7tDlSwiaqruLB
zhVlTcyf+SOtsToh5kyzQB8TIvXL9+wSdM/S4C1CRlHI/24dlt6HtFqRTchdR+eg
/8q9NURsgfB0/S6afzhBRroAexhdu8H3PyF8WCRdEhAs2Uqr3Led/Eh8r0wMucKd
K5iSkomrX+FpD8Q/x/v2UZrUUZC4iSNHhZt4gY7z5YGapGzj87CA8EqpcbaOMICM
v5fcPSNYNd7hC6UP7+1ihfrUgyo5pL7PefVVnDPFd7czcTq+mFz4ct5fIv28VMMF
XALcb0sw8wvwgQ8MJo7AJ/SNdW63HIUNcfVLVr8Zpi1V4X5mcMnHSFuoQNzN2XzT
vr/D1Efr4M4G5noS8NVmL/6RMo2NniUIeO8v4nk2Yx3Uvo67itm/1dgJC6KFi7d9
dKC1S5A2kS81M2GB0S//RGD0WIm/y/UgOqZHz27cKNX9D/flMCPpNMmI2p1HfoLG
IB53ihAYQpqw/JjkUoDCrASUFXQR6O9okZaHSxe7ELNBm0I62c8yJWEmncJetNaF
v6hfnbNvqXCDvFuKu4NPNdyCDz6B4NxvAeDBoROCAndmwPDNef5DBcFZMascviB1
mVnrV3av+IBofCN1D86BBJIauzxYMAiqp0Mitj1pTahgB95mgCq6EGwmCQgA1bMp
Y8kol4mzGE9y5fY5oSVYWG09YdmKgpjfWqogxo2GIRY8crboulsXVPiVLAZpyciY
cOMzZQrr8hFArG6aiYc2Lz8iEzW5KOMPm6hAaccfsw6TxKg1vc6QRYY23ibNzYYC
gmQ6VDlutiwfyGaaTCAA/sKoFy93V7Vbytk9fM0ikTxR/w2MWcEuwGmIytPoflRl
cDKRfAPhDPZsxsWnzUN5wUuX/GIyBwmppfhSUvUvWUmusa4+NGG0N43l4IMHMJ9W
4xLj1BSCxQ0jyJiimMQHmbBdmyAAN9q5O1bBBPO3+iPRWXi2d2RrhuxKTm66Ils+
8Mm29fR/VE34i0KFA9ssIwzGpwIGpo2/vaMSO61VU/vxF1x63bj9u3Pjq9C/XIRL
Yr8RB1vwoqKkbSJz0jPdpDqFZW8JJFkqEj2IDKkBqzxYdXvLq00qwCBZpxsb8lLJ
rVEd8en9aQQCd+GDvFQXeA32om0oANSSp9hUG9pcMqmMU3LwLa8cxWxo+CIRjg7e
TAQ3NBxn/aBtBBFdrNcQWD4hlpDX47LI0WvLST6upZD3btdbuYGRnJZJ9svtvExU
hKHDrpgKtAX3V7XwjFbz6VWU3OeCeT+vb0LzqXpaQkbJC44nCN5us7V6qZNeIG39
D3K/K2zzCiVu2Nn6JWfaVee7R5yGmqHkeBLsucRcMaofl04J1Ct5uWvhbb4BFT38
K0W6cT5QZcUh68JzUDD8XymfZ/NizAFX+TROoE/ISBDOUKVvr8gszdrI9pvh0Rn9
obtMw7vOw0kYhMK3vlx/ijK+0K1mt386ScFEk84S5zyxhj2UzITyZWZaQwtfcamB
urhF6xITJ8+QFxBrdGxwMcn9NRv3cwvFvuI4fXv6s5XB69GuKLJ9aWPp+srOH50A
Mw3GRhuEKkF3PWSs+MXyFqyGCNVIAeLyo6eWDvmxFX521cPFFxrx/9I0M5ENRSLU
sGeRcmyADK8p6qD0a/Mi2Oal+mjIDzgV4kSfOP+gVZskH1ATYD3YnN3Y36ZJiZ2Z
kCxAU736HfFnCWRsTvRApenF92LZpirKf9YoO1S4GnzmGJeAsvdPbb0/lxx+ThO4
s4Y25fV/MXXDHbmQrYg4dW8hOzHTT5mcPtivZeIIOZNPS2ONWacJJkMKZ7OAh6V2
VriRRLa40+TIpy2devhO6WQ56YhPeAhgcfJD4Th3BDYXHgkrTkOAkv2f7XTch8cH
t5bfqGSTORAaVyTDzYKSPEDeWoynbfYdc4+pqt5jGVorjU1/7Wp5r4FfZGZzQAIx
j45ibsbEXedsgSjvVbA/H3VFmH9ism1HfsKG3jxq7LpTTldBQrZsJIGgGdEFlhvR
gVb8f5WSH8qQPtOy6ECWK0Zu0q8HZ+GuP30o9Ffk57pGgD4fR79LX/lnEbdWv6Kf
+BugFecH02Gz2qzaMwHneLgjqAv0MMZsZbOsGsQ6y2vfFtnjEDapr+zNelnpqphC
XGc7+RDIICIiyvzOWjrlXNKkbeJdTMS+io/CFHs81oBV/RswY9lLaYwDREt9ssa5
JyAk4DO1NVISrCXa6haihM9XQtIeq53/md03p/8tsx5IBD0sdRfETv9tYuXptqWs
qtVSKQcuFLJog9fC+BAilQMlDAKoPsVai0cZ7bgqwEgzkRpLo/TlcnIdwJdUlGIN
H17F5pjFC9xMOhxIQbFjUaQupMawcxMMscAEBdMPU6rR7OXBHQ6hWfePbNd/I1rj
f6JV1PGRB0DvPPLIZPmDzffGNiobEhLjhzK2/SE5My+MrN/vcERoSPJfqppvCab+
PVIZ62NSA92YWpC4np67nPAaaLB1n9be43w8JqG8AQZ+YFv/A+tn7j/eFo5jyJdH
RmhqccFaQuiKzEmU4PPnxsEyJHYJHcn9Rs+7SBVCI7LGQqwnhHoma33T/kHnNsOd
6W+xwvwpUKcnnZyEtr8Y22Wi8iDiF2yP9ICjQe97DW+e2tmv/aYZFOV/T8wqD7P8
jzv1elxZrmAs6yQxXelrTWOC7iYb+0YIOHM2rrMw3yAHWvclXGsr0rwCLROsydXO
Do9P2PU+gyGxLRlVF3zMdBs9CXfTNVisBCoIgLew1/FE76Vbs3EH3NZjgRaF787a
A8NIynZjRfIbpctHejP3+R7r6yCt1k8QalBjH+aHJ8XdWGyy3Dl+fdyVgj85TXyV
veeTPYzaY+2cPKrvykSGnCJmde8AtlayDw+lTuN9nHNHHdjBHfasTz8PnTVHFFaw
R6I4XKsCd6Sedo8zLv0kz+1niRDv8XZ2c0Jd07vVzQn5ZJCp+BvWqPbzihudvnnz
snuKbvyaPrGVpUIqjRiqKlmzrPZjIy7LraHYRe5wNln2j2SfBjQEoJqrNqA0vQIc
uRhknPwhjbuGYbDJg1sbnEG7fs2dSn1f+RQ+vcquj4t+xDLvFSqAo/z7Kh3UTWBh
crQiosmPETmyQY0LYU8EdO5lYaLlZjomtG1uLveEb3jEUjn1ch7GHBN7ZLAIMizm
slCKFgvwbJHsqf2n0/1N/+rzGse+nv12tT72ldAlSVaILcCy/Fa/aWKrEyfduwx5
frm/1hxB2xohX5ufswHHVfVwFSzoGUjMsIlRTebo+HeRhMaJaNo+radJ5dDGTgJM
A653xjzA47I/4R2aoCJbpK0yj7sLxheKkXrRIBWyguNc/Q95W9eLKH2JVvbcWcyW
+y91BuMiqGlC3xgLuAK47eSp7T3ns1mCdT/D89lb79SOgeqk9CngDpzI0tfneIA0
kORJgsGqqpkbac3KfSNhpe9ALX39JFyJnW1NU/PiytPMxB689O+Cy1oIeq7zaq1h
mMaBNaitFBeruxmvGeuNlKlcbs0/1jIYg/UqhjM6Set2HQ6hOlyalL5CHmLbJ7hu
La39puM+ROAbXrjrk0B8J7yzBSy+FRgXaBaij9uKpB25C/FJbBE3oEEw+Ix/4zMG
e2t2T291xmM/2l+U4iM80vI1SA1Vlj1MNvm6XYO6syWCrzbn5o8QkHBa7MsEokVP
G/uJ3GOICanZdYHIFcnH2ErcveUVzjbIbTcEtbgdGgF9XCWYrboxhXwbkNKn+yCK
gB/vm8KquDGPeC2NYR2mvjs7E3dHkPD5H1IJKQ0gETh/S43iAU358zZ/x14LItcN
60evXXDT5yIn7iL/E5+dJyZRLkC/Ap2iWwU/wLnP5qyIIT2R4139CJo+S+94yz2X
UC10lvN3P7l86MNd+SZbn7j7Qp02DhVX7ESyqjY7MuaevpGmlpVcSbT5Lw3J0e2F
FIqIqn+WjozT904bpHrUrpz6BoCLbQ4VFG/CepvqSHb7pwRh+cT/x1JgPQk8Jkky
n78wWvNHn28D995+Db/kQhsFKTfDDjI6TQ+ANLscp76b9QOTXhsdPXOqSK3yMobt
zsG/V2mwoCYbLO73SBiTdyrY2TVIQlWcenY66ada6D45h/yRIqXITKVmU7HjxtzI
xjMlmGBX/Jl1jiapt+3EDqZw1492hAIqBIiOEyluyaAJVZmBQvpBGAduiEITlwme
cp9uAxxvHN+V2I6PSbofA/lD4CEVX0uX7H5Qe9JQwmoK8HZwfM6fmuWIJFQSEAOz
nz0ZUksyf5Lz8hHk4ihz93gJKd+kd7pj8I/3uD+vAZC4CsMt/SwtNj2LsXSreLtU
Ci7xVuz7K3u1MVdjPLK7em/Mvkz5QrJaNbaZFs8dnug5hBwvvlyhQMXK2JAeVq7D
/YV7i/ma3olztG+355G9pc4cKBHRt5yx4nk3oDG/V9Osj3vCmB3ocRJ9EFM8WbOE
j4E2QVnr6X9iCqu4sLCoiA4gn1Mfj2LFHns4utQWCylWd6tsHcWH3B45dL2ttmDs
cMvI+DFNVGSj0KKcZNDDovN1bD6OY02tnSL+yuey8vhfEHfGeizOz+cd8Ul1+Qul
nXv34GByly8LNNlb7Rfhfy4kujHMu8Nced6794g1k9SwqVnvzp/qmI7ZebqI/hL3
J2/JjWj4oko16qBs3JwgkzZRlpyhyZgrV3kZi01r1U1zWZHSwqPtQ8AhjFShq9rs
BZ4Lj0uM0Wb9Z+4om1sXqat53xLQF8GSmY9ZF+tIx5uCUVUu9YgaZE3Yo/pE88wB
p7SN11qIaWta8Crt1psJfG2J40sTEnX2eWhN+Mh0rzYTDTv7H3iU6NsBnE/NjwE0
ibgFmXcd7g8tCWLrgq1hwZyVChItQQFFVgzm0oaKFzoMSJPCnnHSybe3W4yN2zFm
VewKHGRg/P07Pek+K4nCntw5OmwGNa/e86lIyrgf8hN+5S8jIhwM7rBl+tl1+hVz
HSz6QjiZsM/sPgcgEcrsLYlCDuqgGUZALgcSCIRMCxAwMBee3pKtBDIZxa/Yy6bf
opSSIUCbfjw6oroz8EpGAtRHK/Kzv73TeMmORs3UcY42pgg8EL0rXLkn5MCEYs6G
GuczohdPEJ3FGUcwKU2P9yOa+B7eu5mlenI/Sy3ZJCrGqBz8VwZUP9e5WRXiuSEa
urPo1+3ImdA5qd1eZXzFYo+i/ESGtIVzBtPS+A7pCQ9k9xwqNDZig/4Zm09WXiE0
Gz+r7sQNQbot4sNFJqOH2p2gcuEobADdVLu3pTryQkMZYCz8fMS2PMo290IQkrtk
sX/stIiwLt9VwacHoAGUUaNsDltJazsbnyrYcQdxbeHbXhPI6zWYb3jO6ivs9DWw
SL974VhwIeB8PWIfMwvRBQTmXeTKQwLF3TtBKpB46mRDw7sPhlnSyH11+KnbxNnP
Jk3HcMVKHrbtrdtYV5ix8pWbd7yq9h3p5dig5gjk9Qs925wHeYkleC+tTk6gtlP2
C6INA0xG9ooKWQMB3Ce+avxo1gHLFsQd5E6Ja4dNQOE1UMalFQph6CGX4c8dJGeb
GzktkzS5Ubfie6vxPbD0tNg71enGl5cL7PzQb22p+m/DmDZ6YGBg2IEwEUPFtlZo
4M+OEvMEY7WOutB9n5sjWUWaWhw1OiQYDMuowCwn9bdNQFJiwolJLdeWEj3tEN2D
HHuaxaeP0B9Xs2eU5gQjsrDrpFx+ar50cePx43gE+tSXzaUJM7jXFeiDvpkAZLNd
haIYLWDwWwxUrF63hsmB6KAEJaa1LWrmCB+5p5uogixhAoguAKAwXezJc520f6+b
B/BV//8DXeVoQfmO4n7PHee1ivjAbz/4FKm9RJNk5gNL0sItsP6uCQAo79WsCmhe
vD+bqWqpT3+j5nGcIsp2g9MnAtiDz7wnliI6Nrj5vilyaAgwultaXbhHSCDPXM2h
0l1V+QITFXhKAAbcsmOtlKocAO3GF3li5GXlNpp+GgbFMfRP+QeIjmBORepdF98L
jCWq4BXzMEpHKFGkwt2EvAZ1ZAbBYHkvIROGdhFDqR3OSi7EHurtS4j2k4+UHEKp
8LPuwyd6FiJWU229SFaudsiGstRqy3Fd/q8Uh8zrAw4nLpmfK2fSSfNkD7k4l6ud
RtkJGDXP8iIZ//uiUo7p+0VJR6GckeKOrMI7Wz9NTOqrfObhb/rW/Dccuwe0QTSh
xSOA0YyLP3c+wBl7YhJT02Yk6uShMgCN8ufY3B0ZEt0Dq91KEtmYFda+NPgq/+L9
pTndgZZ5xnRyPG2iJ+dPUOHxYCknVPJnw4Tkb4oTI73LoJLBsSHjotEVnF7yrjCl
IMslsmQ2BDzX8W+oHYlm5TzZ1gQ5mDbHISQYPDIop/LUYVhRl8CQomcZXZhFFHul
ubjZDJ9ZEF+1fBN7gUEtqITBKNmwP79aYJrICnxUyA3qx/JKAbgodsfOTacZX3pq
3sLq+Km6Zzfr3SS1GhOp9c6XcaqBTmno2M/TtMwSihJChU+b2qY01Vv5yvFIbLje
h9/vhF9JYlgr4j+QrKXqOd5TPT6LTIHVOI6HZVmSXt/qLjPdU9141S+eEBV9iZ1M
A+m1STRDJJJvL5StH6vJgSi3TF6UCxagWdZur7HRKJON5tsf5jup9MHHJTPWtJPQ
QaSNvl3OERFxaHHF3uo5WS579FOcWnxnFD5JFHrBwo+RLbRY2rwySpu4D8XCovyT
1Y6UwM7mJiWnnLNd1skx8iNDUqRkQz2iFpl1U4qUsDgLC/XSMOvfTQh1hmVXtsc5
Vy3bkp5sp6H/h982VoM4It3IAl413nflbv55LNTmcI+PDn2X4KbG2uMR5CEk6ca0
tKyFYphQLSmVqNjXCJz5jMVuiYtPsCAc44I+P7PH0qVGoRZBVtJUFgDH5AcTpoKE
GBoUVfUQ4x5u2oteDCw+YB2He1TniWFO0HBufC756QSdjossJSmi0iPBybwMWY9g
MeYzp3Vv2o0lHHdN2hAdSXcXCREGEzobpKtoM4+KcztdCIIsg/7MDycWmu8To0RR
/aakpIbKLQNVTl0AsCsVl0Z0Z8Liv1om7LArL6iDvgamBGZHTZwC0tL/EWuiPLus
8ezPdWfa0W8A9cILdbXDAaCxUG4Rk0Bak+GIonSDRXC7Kb6f4RJbxmRYomlUqTad
rstVS/gLoNPv+lOHKKLsYaLolcV4cZZ2PG8W8OMZ8VgddPEvNEEsJrmxWcg76x5K
8SdljgDnrb4OPG4/PKcrYDVWuZ3CzQTuA4fZbmzUbP5CPPpp3tyhXjqhV0x/FKGv
NVI5m8c8LlI6WiJgC/fvLvpuWLGXRtO6GVhAAdLeXHuxO5c73JfJibmbbJ7DErxc
4eOtWHUGHuFByZppVFAl4Bt1s/w6x8T9P9E6SX01n6UVWtriyarUU2Anau87e0A3
Fh0hSdW6hHy9eypcrofmFwGEkFiTkn387r7Ef8rjIHQi+a5gDM0KgmzDl8OqufGs
tHKlH5ujoDGTBP/AiN4DVzXsOIOG1PKlKJ7h7eQyBp0qt3A/znL9G5ImH6QQYnvV
PTKIyPAClI5wACCRInNcW5u9yIPyo6h0bwoVSQOaXP5FVSdA3upAlpVufLCXOq2n
xLCMX8LIH3uBcD70YlBt7Gvp2fxfvJn/2Fi6ft4aCZyg/nmC8LwueLpYZzYbzJSb
RNv+vK5Wefqvi+9ZDB4ZcW9e6Eg8142r0lmgZqqCyH1ai870gC6bIHKszZTaHt4C
2YDJy+pGsrGGIifO93rmBG9CZq6qZaTNzOPXI9MB4sBMt/0c15FDxp4nYuKvCLv/
t99Ozge5h4BoLqyO3WmV2Nq0zLad2jZHwkoQkalMzBabHSTW3LgeXE6vRa8fK5qB
uQowKHG2SZAGIR0SohnHeuiIUCJ/ufoNt9oBU9L/zGGws/E8HUqWuGb62TokJYqt
Plkq6vbzdD5w9fv+Fts1heo0HcL+/ITr+umBS8+OTQbormiG42sZEZmRcLgAodUj
RXXQvDbs/lIIo58k+I10IsXDMTeV/4yDcZUGw1NWkco+qPpUnXjkSRov769NWBkK
1phn0Llb37trSDyDFw4YDjcju/KuhPRLvGli9sNSlmpjWayRYGGJ98kP1sELR0ts
Ze/ERlINheJr6xvguhuSwvIKOLxHCEcpGbsPBc3Piv7/rpYGrs+pWvkj5JfV9Y7m
w/TuQbQbe0ZSKw4b7cQWGnq1w0UbuG8fVqwbv13ZctNllW898JX27bSGnOugxzvw
9KNOcwRyUxvcz/Pb2lrQlRdFsND7we5v2CsXwGSaUNlNZY/RoS5LCDKk8aKRJqyN
VLWwewGDMSX1DyuZgAZCWV7gml++najwGfNtOtwB46yv3dfV9j8GlPCHw+r7MLgK
8E1d6Olz4ikEvvZr3iM02eEjk3CIRWCoTUZzpRIjBGIfYo0T2t3uzyOp7gpp4Ooq
4bzIbae8q5Ef2Ajvpk8yHS3WGih4kJxjysNkyztnpx0I8mcwfhlqPmznP0UfeJYC
ws1cA32YEyIts4xCn5xpYmDAiqSDVR3wzyAnDlEeWbWFO9PEc0Tagax2bmzTuOWX
osKXG9wKOqdcHbLhxQI91+0hCmpi44/dsqF5QlgwQM9PRmi3mvwEaUFZKXhfwkl6
KV4Hlr96vQpeVjdpZK307jPPv5ng2oRw6gb8Gi1nDvYbzz/w0BVuNX4OeCSuLaAK
NPV/ExH7hjnxivo8ZTTQWMPio3deKzRBjTuaGeWKXrI6gvHfNxe0awqGK5bVOfCp
pNtybtSGnUIxLtT5X8JZAqufAiHmzqCxxBoJo63v4yLpFCfmhilAPeV2POaXxpVH
jhMDQxb+Sp7zEvxh9QduV7NZSGJqGhXVqVa+x3eB3i70u8w0zRV5K7lBCiGI4qbF
EVFPhfPe8uPOsQcSLH925bZrG3P9KgL3svM7eEcyxrdM+EmZj6kanFggHrsEFfik
LkBKrAe6fgpTHBOgGQe/K97VgkeaEw/UGXIoShGBmG4qkBYbn2Dim51xpo/03feR
6QcnyqDRMTC6XCN2U+vUE2vGBVB+L5EgKCc5fgDrGXJVSNN6ViMDT/hh6DbSS1PL
zH86IMH0KT+MJXA/x9s2WrPjJG/Ex+P8nBjv2vGYapIZyGv383BQwbDjT5q6wLun
InBAuzfcxr1fw3IZT6tPi7qj4APkGhqX7uJ8h72hP82S99RmyVd0HntZSjlM05oi
ljf/th8rtWh4khHM+H8XWSmEVrNj7UU7XoT8Ptg/oaBEoqOznps5xAMeWljtLZDw
7hiERzIFkZ7Jole3TUHYsRyHwwCaCLk/zT+te/o0JQua8hu67Be7BCy5P+6QAybE
lDWKY5gb1zduQWEc3aSQlSH4/Y1m4UsjfV4eVWKI3dJlhHAce+wEZCdwU7Os0UGq
SjfIjbtXuq1IdUMcJ+tQSC2JKZAMYbBp/U0vpB4O6NFXUx14KDAlfjh3dVsaWQb1
+R8SLuK28ZAm/vFdHgjeIFja4PA+r1/su2gRqZsXHDKf/wL928kCOljp0X8yyoLb
ukTTs9VrNMs38Yo9zNiSwJvSixoJU0r18+c+WQtlpzE5B0mbXwGoCKr2o+QEGYOU
5gBAVhMc2/Ig1mfkzJnlqID+yBJiBV/ImWvpVsmxM5pWtGrFiFQZVWVPxJtmplBv
UkvdYKUtiYZSPKEYuCO96BjAJt3A9eJ3VrRItlyrzljdBjDl4j/3ho3X4SnfE+ck
A2+by8WMqXm+GYu57INP6jDbnricbfd59xb+Rcq6p9sFniqtzBoPiX4NThvnESbN
oc8eEmH7iD2vYjlMGfdiHHPomlsQbt6ULgquIVl2ggTtMHlL3ooI6njV3RkG6vBH
7oZaN4pJJIc5SRCfy9qV+tL+A0zkeQKhlW+GCxFVplD9pYI1r8gfJqopr46MnzmN
6SQRHIQxSWUXj9eLqtHKVrpsAVX01AWrE+LHnwuWrG9cZYKi8rZa8JJp1+6evaX0
SgUQR2vhmYSWJEF9p3NUfl08iDe1i6TgeAKIYvuZDngo/dYivvggDPMNOkcP3A0A
9cEG4a5MKugXbrYQFeRnQtSuNXj+qZCiKeCxcFU43aMwljTQd61YdtCvmKDKG82a
Qz9hnkq2lLzvw1Hr4+gCQghSR8HdhxyXF0r2Okh7FdlLMcvIc6uQD262VUX14nyL
zV1BgbFobshaAn9Dyrbam63Fq+YOgi79faiKREzy13mkZoNi5sFt5Auy/PIJumXx
Px20K6UYveHWYPsk0oMYzefFLXOz4yCQIu/bbgWOU9zZ4xFipHXsVYB1Y3RNxw0k
josy03+ndNG4edPUL51xquKUjtj2KNMcg3SKFzwnhaaUuQN7vIYvGNdmQkstrQYn
yzBMuun8dFO9TirNBgUt/ggdDZPoaD4uw64CLHMQhTL3i3Wh2mdov7ScffRF5sSa
J6mNkior0EN0doCRa/dnOt8LG4VhV/6r4EIkiAeTb6/dk2+GLU96vFj66/KtKjkz
xkGTI/b/DHcwE+vBmi/Y9b+7r+oNkECacKf18f92DoRTo9W+y4pJzqVd1HUX6UoX
RtGwsq5B0u5ojhZVBopZug04zzXTW2ybRhuVkljCjCiWNiUb0ChlYkA1GESk+mnT
Uyv9r9cO5ycK0nawzOLyVplTExVfvn2FEbbVkjc9Ihd5AC0v5u9ub57rUSUtbuzV
Jy8Gm96mdbU78TfQxnP84ILVpZIzN9mvYiqh7/rOSsLIli9y3xkzBw0KvjkON7na
cXX9l0Tf/EX/GSBx5u8s1zXScwreAnhaPrefNfLBJ47FqAzA46lxXHVREgYsaB96
fjEcfTiUyvGsnQjNOt/w3b4KCSoT9YVkzpWMSKB6dYlmd+nx50lnoMiKroN97H2z
oODKf1qn3MGjkSdXY/HGcFXjBz9p+J2dZFm1vR9/SR39AFGwJRDP73nla0q4fDDD
iz700mGBddRHsq+OHUfAHlDBkt+Uecs66WFEiH7SZInJsaauijW8kGBzLeNGslhU
+kvCkzwggpkyjF+UFHsDj5P0RxzXgM+DIcl0ZuFzYnPe85MEvi3+diIql2qYQ6QX
KTx5DHYhedfd4QB6JHVe3fQ+i543W2g5qPnGOCRKMjP1ueVjZ3t7XJ7934L1fmHM
jeRoaSvLC2yGx125wK27apV2YswVUnCPPOFd40x3XzzqQtETck0bKOVlqMxP8Cif
HO2LAPoRe2NXG1EJJLQQ7jUerQZkiYA+6fzooNCIirJhsnpE66ITbjf1smUMMeUw
vAcvGSr7rcqyDviI0Bof8RtSDs7GeBwHuRzAz6shuOgN3IY4O9/sFiZ2Afaj/LrX
e461JVkp+Ri1HFWAHOmayJliVln2agVtB3FGjcq52EgbJ06W41xWHRTj8qSde+hr
bA7mGAwth6WRBDZeeKuqVe4q1z/Q9rhe0wsJl+z4LFcu4a5WnpnWwxjhPk35cEBI
ePJbLTEb/x4EbPEOxD1RSF0UxF6KEQxOMn6u3AaAUV1JdDqPu/vgDoZcdEctEEUV
P4E/gFy1hELx1IDPZJZzml/LX5VpolHToWz7EJk4Vy/XZt53Nx1l3IG4kTIy0X2q
/FK6VWWbpOYn/iNDY2fPqBsMvuf5jEbJuBleGv6kn2t4uTjEKmUa29xWUOlVroZK
T8ClYH3RFD1BG4TYa7xO0SqPIqiIIFauLQvXCXQ56nYQIVegyX3BmsxoRYXAqeHb
6zEKTDXTMMXJpoLcqttFsBVq8czahf0Pg4fubH+ih1opEmaC258Lu8u+cHwPPaAv
suRT2OCx0og3AH8zEpc6axX+yN6/qx5+JCzLR7uA4AJ3ByAPhH40NZJAsMh0jaTZ
8iC1NqlOmtuRxxLQdGb9QL/29mjOlcS1QWhIWevhxXERYONDfZ0cD90D3VyCzl3s
mb0qep8rHqm3/yh2IwBDjs+N94Hl2FvxGRdd3ItzIBplx+zO4N5Lzewpnnm/ZFEH
N7nZk7CGL9WYq+R5HhWg5et8Op6SD7COylEat4XC2oW3KClbG9PJSBfe5PtAhCXe
FAoYQc2IXWkO2GyWpZj2H/3WadJdRA2r437ZWTdVJeSlzXIZbeQR0QZ+lo2PfkH5
ZT6zKBRZXT8BZUrZS6NLwzGVVSd2m/tRwvScalTp61JK9ALTn7iKTj8BSKe9YFD4
bNXMCCFOxmQQ/+POwfLYHMeYeCtv0f9k1PrFuiJ0JQOr4sKHXQWLrTVkPg8ReDG5
NaCuKOr4Bkl1citZVbA8Q8YlqIfKAAtHSr3LmhDuSAaqepCyLCHm/r7vW/a07EMx
ELouGbSYjohgZC3wi/fjF25POTH/3cbPu7kkLcMKRoPoUxzEg3I+9SYyZmU15516
mbk3haaDP9sDFQ51lNjVCf7AFClhfmgs9dOZYouziB5epEmXcrupoN38Fd03NZum
pvSvDRi+6tdnB3cMsAuJAaAOwFaxuai/z8e0Gas2VdMFvE3Y9yBl7T6qxUiJXQ1z
SW3UJNxGMLvA687NOdgAlRl17+7T/kUuhskIIGuPb9zJpbn8jVLfv/wsxKKPtOLs
UiNp7sl718CJhe22ym8PsWxMSqjmpUXphagKGLbNFsa0ZxAkOmOMeiWWmQk3vhd2
7SOqeSPTAOrfMkHxomdzR7femwG01yFMoFrgKUbBxepR8cfJBC1N32OYoKzzuNaf
jzolVKzyFT7TF2PHFrNbNoe12t2XeNUSrL/sRnQoWSpKrqms9WvV/Ppn97QmiDD8
HVP0XCBwYF1yYHillGIBXZ9N6vSkFMiMGxTTOjaymUltru7ufriffvG9nS0kPfEO
WZpAyVsZax3LJnnumtwR/DADs8wCs8R0cUX/q3Gw3bKORHgDCRHKstF1IT5cbvFz
zSzS0ybMsTeFqYi+bxtc/62anbm//HPezjAe7CoTcARL9ziJcyuw2uuH/QUztg4T
w7JcvGWXFV2lmcLxWo4/H6voE7fHjQw9kcr/hpAFkCL0bJfkUhmmmxjyWkCM63bf
LDFphsAKqTlClH5UDPWTyHEYB0N94QtyPJi8nPknRcxmz5L+Hku6gf74sRPbAu0l
wLZSLef1VcDpKWgtq/trm1MGKu0RwzMlBjSV/iQlPPUUoszDheS2dma5vin85o+h
gM78SAKLlrZYKHnIFCwMNIRA7zaUw40xf1ZgIGKMikPIj4LvDcEnf5Qp/i1u1k3U
bpfpXPltpDc06xf5CTwHO2wJ6242MeTIibvGZPZxbBddQS7dWr4KhKy+FzBquKgn
22SBIYQbMERMG6govKBwAVD4xqet0xNmCZLHWhpfBYzg0Ve87ur4xAen+w3Yt0bO
rKL7OAaOI+eVYy5V7RqxNGDhUfChaIp5GWfBmSIR/o1lmf5VxYEp4hIZ0BkZ6eAx
lZanvoFsz1GSl93k7HBjrcPuTXAi5UD5X1ipBMrbRZLJU1Ce05AqnziF5QFIMHp8
4YrhpLB8RhJmzrUPRvIxTdKoyThRlJHX9enVX4J5oO1jrcYSTsM2bjrSg+XNDt80
nAUxuSEZOICA/xxYcWaiygvVMo/Hw1j9zXHd6w8CcEcZyUGKal/i72GiWThKALRu
ftbrPvgiULD2mRaTuUzFS3OjJfTurVXwQxxiInhyhwljh4oHNkeFcGQot1gDWpNt
4a1s6LbKQm3gjQsq3HSIOQARKzM4TvgBAGq3chbdzMw6jOZbJCXhuWzLqEkTYM10
zA/uzESBjfl3eJikxmfTbKh+w/NMXI2J9s4snGiNO0bWoNW5AGCy1PwWXuURnNod
fUXGAlqqIoySq9hRvfDcPBUy2oetj5vzQnYDtkq2iIpH5SD7wECgMPIZI6qSegXT
6d7aP31uwieB496RFRwJVThtHCVEGVUwDv294Rkyd0de9/zWnv6oy7yJCASJxjeS
kmbgtUGBxQ2FLauRNGv43zSOXR3xVukQSdtSRMDf6nspqh3tex8KkbYP+Z24Izqs
NRho08sh+Sawa494jruQrjsjg7S6XJVyO3tX+sFU3TzRx9wPgkxOT6ij1GScDzXL
EcQjIxtRZr93BPGwbi+W6CSlh5Cu+PhjEYbN78LoehmeEbsrKf4WpTeLA8UQaLsi
67dFghIlQZbUSPMMgn7HKGNOUFmEdqcWJoePNqPQjc/4VmwwgaNbqzDS5O/cssT5
yJRVBQHQiD0CoW7AZ0r8YOFA2dUonh+Y88pMM7GcWsRaoJRVmV0f3GC3V26IG2kK
/k57iAl4roC45egi9KPCI9/aAacj0ncAshFs8BgeBaMRVFykVzWp0gBJ+vAKkUVw
zH7RWx/GslarT0KCLgq6GMwd0WFncedrnE4vqN5kYHIk09ESgYuFOR5doPdYmcvX
oAwU1W5dQhH9ip2znVSZUVXaZh8cJ2WIlVZ6ohTqRbt5OPZtX/cABH3j2FVDjX8n
y5SU3SNZkjjT5b0lvtxUnxlnX4ovdvKTDzR1ZhWoVUhVV+Piwe5dx2c8NdU5qXTp
+5qt4apmqrG4X8RUlsu+fyc1sSrATRHFaSzOX0+k9TiGJv0TCFOyVDjckQ9XmlsB
+390yh+TrCzNz8fhN1VMJX07eabZUq3dV35GZUfhqi1kr+Afg8pzBjmLljBEZHEt
RGFWeVpHEi7VTK1jDWl01G+ordQca/uqwIsHjvttFFbbBeu/hy+sGHN8eYgPTuqa
QQopeaDd92id+odpLk1wCY/fLXEO+bmioVf1TQ7Ql+bjD2AqnUQMJ9ae3GKK+Y2g
CVvtP2nbkxARVQB+3D/ilLwQB3H2pJOrhc6xpu2dTJyDrSit/sMylL49zvZ2lXA0
x+DvZNKeZlz0lBCMqwEgBavppFTc8bhUa/IZMae8BgsX4CoSFiRNqpAsqUVCMZ8x
fUNSx75UY4VFeXWCyYf7g4wcDeQcgblum9PJuo2OXvS8nCknzcGLuLjQRMvhDWY3
IdcspNJ4OQ3uC8MUJgB1SPNid/RPrfBnlSv0nIBXnKx9bJEZd+KEgax4W46RqghM
uDaPTX7Gf1XSzkN2gzmsMnffqHnETxBrk0ZduESX+f4V9AcllUDmWZV8lCsHKES9
KVRG2tQ1rOZ/2ZMOipjr3ggzmaBCaYxOVEs5lSrUQYpT4hZzJSN7Pevsp1HpWZgR
EClTAgtVQvuiSoWxy+4PdCY0QrQvzqJkvg7soDZRs9FXHry2WlbS6n/9CBZWE5JP
Cel76QdgKyeqxvyLNrnrTApnlkbIm9mT374jj1Ra/FWLv11jgWsErvC7TV6CwZ4M
sW4Pn1frr7pJheASAoJjHGGbHIia1p1fA1uvO729Buk8Z3GaHQjm4YpMQJlPDZzZ
+SknGzNUWQUTr0PUXocVGavM3YbNkhakHm1gEgoVYGey013x3OMzmLQOSZmUyQ/H
3u1fivutYiP+CQHLmViry4obQEXZPdFxtw9Xvr4ki9ELSvCg/HuPyBrj0fUkL8R9
8e+nJY3XF6fzD8DkAdeLwKw/BwBx/03Wc4tB2yNr+2aRZL42bYAvjDsK0libRRVi
eXgSdJM1oRG79c5yqfGAj01af8HEyXm+Z+dFCDAv3vG6NbDGwleo9U4X76jbQZoH
z1OMzITq5x1106ZDVhcPL9rfZEhC8xGe7rzwrpo8ptbjHLUQPmq530c+q+P8edHq
HGhP8TqllXYwmk058WEmkhY69mI4rpLc36MRPSnIeaCXtlhjAX580MOWMsCgGRaF
v0BZEvzMWct3IAud92tJihGZhndi25OXc18qPxirKTkd5MUPR16pYopN96h/88A/
/ia/+qYFCjMlflE4fjqIuATdHt/HXyAXZrQoYZp+PP3HmhT0M1xx//p2UJKLldI0
QO+XRLhfDBOZ780F/+mLrbDx30tg5qds/6wiDqDfJfctjPgQ+q8m1cR0EUSggNjT
JbS+7OtIRuo5BY7yUJsSxXbJAuegv9bdKoQOBxAawO49/Cc76+4isz1eVYkowmK6
ztBpwBckh/KJR83N7rm8qpGwvWqYY+nYA4t0UvOQHDQD/fZBNoeNv6rLf1dlVLXM
BF+tBfPNJscppdfxi3Qu2lNCdqZw56hm3rWFQ2X26wLeoYnfZ/NNeWSU+GlLdpot
1GIXF4DYoLx8oY/wfPWx/ws1Bz114O2yVKCPUKvfLr9n4oFHi8CyzdfL45Dkla3z
35PjketdRvULU5daodshMt+h6v2sePbgCvWxW3hnqwsPS8TjGZSd0wcUsHyUV7Q/
PkNfwTMarFoqRG7UJJJHh+wxz3wgMtcAXBlACBp2Y7nlvaGM3f1Yiiokn7DXWCRD
pXtr8uPkTWnj+DnjhyiF5vqNZA6bCNzPHfkFyBs3sgO8vrOkWWjyODPQDcCIXVNx
KES21G0/LoTkHtpstOakiNN2a8A9vztfiuED98MhH2/NA0AUmhGZ5PoQ3p5rRWZ0
ZRGUyIN6FE0JQSgEyj+oElq2H/0i1iLvulefoYYa1zUanSzXlHI3XXZUbdVPeQeL
agjkKFt4yC3zTvSYdAhym2ORgN4NYr4EXlTJJXeMfl/Zo5QKgOMqt1lX3lkc96lm
hUkz4U8PajmopQtPbYq+w+gpT1Vz5sNpt7z9qrwDmiOiLmrgWZCU77Q3rMzXuvVH
CaTyEtLmOYO7WOjg8zzXg/PG/xK+o+ofbSfA0zIxnF0GbvmjqpYNlNOtZnDcy8Hk
y1v55vPTF64KALW6o6c4BDn3SEbrAAxLvxuAltH6zhV+O+Bd2MYCpACaf+qur+QR
u0cAfRteK+Ga4UWE3FJeQZbht9pHRDKjO8Zi2PTeVTuwH2njFFOT/6iZvuSqpnPe
sVXcib5YQiKH+rB8peEyGFuqqEpnFRQXFV2kooQYMrA3UUEei5K+Izr12PDvhCEZ
Dk8ZNaE5Gowdsrqowxt+NRjo/lCG1yclYLsPWqbbA26xO2ggrnpmiNl9dD93xOqs
MLHmn8Urgrcv/YZRTvdCaxfUfvuWz6pgnSUvUSP4edQq45krmM5GyqODoKBmeFUM
C2mhcCuIkj5kngHiv8TAZI5LW/2n7OMnjgqMvaoQZFUJ3ODSQ/173Yd4WdQbC+uS
9cEJzDG+GkygoN4rvdXQLuPkLPI25EDY8xdX29D04px0n4Q19V1aPvOV1NPxw3yK
0+roFHjxTuypqBLlW2AoTw4vj0lrAthilU73nZNK06YBj1pryo+C2S78JvWwwTc/
B0FiiqPE9dWoNoFqJfqqMjGBwQmXfgGxI/JuVIX3GijPWjVhx57piF/GRNkRFB+E
X0hEjY+QrXUub8DzxHO1uzW8le2GwVlrsLDrRNWs/VPYA5dvRz4gIF2g/GwRd1nL
HxezOLe+54qXMeCEb3Et0gB8JjbRVuLaZrzsxnpZyFDb9FxFy11qq8SLihlych1N
vGyQKectSpOhVg9rrG/ErpbSTs8+cZkk5vwKqFYusps5FvGa+Wz/QBy++4KIrmc/
f+SOQPKTW6/2sSfdmxsC50kPddlV60EkK0AInUUWZ9jkmGx9uD3DWmVI7gW10rdv
+SbD6i6rJ06BqGAEp9tXuyJH1iilS20vdkM9nAzi8LDVtnqmHV87gxNQzbnErJ/U
1l0EiBpFr+yXPFzWs+S3EJzaGGG7Jd8UeuzAJhI5GgoXRbt8hAYafRXw+5VGE7Oj
b0HvTssXCPlqFcikKHlzJsmjPIBt4BscS2GWnzoStdK+IipmFsNmmkVZZvWUt5gY
yahmtO3xguy1EMZFhTu+hkHtxmJMmvdLbl5x66ELrThMKIBBRK8GhHCDyroRII40
1StRutYjzkDgYTwwj/dqG6JupUT1f4wT5Ng8rg/9Op2zYD5Pzq6S6RolJbB28WNm
UjCT1ffLRbK80krxSFBodQRwAKaDDTTgWvwrY4n6xKcnqGcI/A9CPHjthP7O8xA9
ByFQqoa8UpnN/KEPFbngU0NAshs2Z04e4y1G1f9iPJZAjH+oSAlyLmufHfu99d3X
54PdBK2KZ8Bc5aMqvNcgzRsj/51civKosAdhHfEldNmfgzgfnIJ9tSfOiVhRj+bN
cAdq3IXG3Ms15hz2kQ6tlKZ204FPJyFDsepadLVDY9KOlClTr5HYzkx71GJRj92r
+GTxSsaofzH2zyr5bMXnng24bn1MMmIAS3FxMfwWkV/Vz+o6E6Q5h6HijcexfTw6
QEPsp2flhWovAg8P4a4VFpJJguFhbbpfqerEDalwK6mPdQ9xyHBX5NAog/XOlFFT
5sfndjIKFuYu3p/xqgO3+zprZwDrx+/IP+2mvlRYz0Lxd+E71DSPNQ/cW0GAJSLm
FrONAmGwK+D6l6apBQoMs9JGdv9RFyJXvKZ/u+AIdVePGvkSkNSjELzJy5eLYJhf
Tjti2PBpHRvTb0I1xbSaEJsKqWIs2zr8ZYdIofS8ysEgTsndJIGTPfD3sN3j0fJC
3yPlprbzMLXwEfPxHGNQ1xkNic+WuEIMZ4FByvl/3HyRhkHxLDpRs2Adiq8v9AxH
ghkl7paOfv+IZApdUwkjG/KVPZq+NJEv5H7RQzeptgMu+IlHetdH1zrp1YyN9qtz
hlba+fIgOcygU0KEbpvFrZFQFW9dgiY64MpSUWA+/pHNLDPYOvbVox2bgso7Rh3D
yuexEu+Fj9YIp16kLLwdbsPc6rHcbrtV1TyObC/UnRt6UOMgrPblTtfXhslKmFtz
Dg8aFzDjR0ee9ishhzJi29EnwF4DUuur+pLwy801TzyQNQZ0Bm8wnfBSDYBg1T2U
Zpe8zAIOAvCTOJyEMwbT67tMoWOOQWlCnKNZ9rbSBmRF5wmdKF4/8axBeTYvWuIR
eF0fBwZlG4PXyl84ZG7gx388AR6bmIAIgboxtXkcCCNIrag9VTFJMwcWJpjguAHU
42bcWI9MV4R8H7bIUPc0Kl57+tDQpJqSPDZ5z1sU3nkE4f+JDQ4NxOqFq2QBVEOU
LtYcjx3gWxVHpbkeP0fdsZFFutu6K+BlP4KQr6CslwbOQfdWiuNut6GOPeZ0zh9C
TQacDmwAWjnazDAIxyR4QXHTTqFzyJt/RTQnoUE+07YoXvNwQ6tE+u4WOreZEhAa
LmDdmWPQn+e/FLzfI5ryt7px6754UfqeBClVK/ieudsnj5X8jsKgHg5kDihwJF/u
UxRtYmZ1pPl3TGpV1qYKtpXx0kUh7S8Wt7oiYyDDKF6ZzhP7BmU7ZG9k/HFgKmV8
8U71A34SDUgX2kCJLcDY4xfwmAq/BW8W1gakKtP0e/Eox2RGYuTB4l7HKBzOKYOU
da5eF+DCm05HrBRlbrwicyfq44U2wMwiqLHJ0pSkjWUOoqewSQzwxFqxbc8qzSOg
2hb2/d5dYJlfP2MREm52DXRQVUyHuFN2yq6j6O3APmTo4QWg6SvhPqhHMof32Erj
4jsE4sQUdE/ya3wc4EP4HOcOrmWwXjaEn7bfojOTI4v7IZ3sTjIH0dLFhr8VyuB1
EfPtfi6trtnmQUqB8qptdA/FKOro6Lc+F19YSpovDb3DMpF1FehBrfKFpBGzG43e
K3kObXneuSzgTluWwrswBx/ijYoQLdarFC6XvxVp/tP8HDyWMHxUNo4tSYKYBgto
lBXROZC8oYqGB2wFfdQyCWs1vowBku4a5VDpra+FFi8hfgWkEr9p3Oe9Znhs4aUc
PqsQpxA8AXArKhql1kc6VfoqRgeXn0FCq8j3sro1+pAx/v8ZeFiYAtVP0SILddDh
+nVB8bJA3lDCLkz1Vckwm6Yt5yDUrBTy6sPFqLkLNUUSK/Gfr7MdUaJfCsvcWNkw
IIYJt4Ea/fjvi0Cr7YWxdJldaC+AWIDvpMg5l+sKGN+hf7y0XcXCgd+7i7MM+rtq
rAGPdxoBHsSesdzv2yBsWHKr25vbbUox6izxVs/oflqFmnE0nU0N1W471ElQWgcB
3aVietWF+VXaTSsUul5I0wZcDxLEOXvNPqm/UpYbL11qhwDsKIBQRT7QY2fJy8Ur
PQmIpIn+hHQ16JSMMZqaEnX4XLJ02/XJ8us8YZzD1a2Pw/xzwu5bzEbsdtOwXfL2
uJPd+b7TcLiw5vAs5i/157GeFs3klglKY0QAwu+xHrlHauGkPpEK0YkqMcSdTfgF
7rGj8PzO+1K4JZyXeghIcwD0CSoFqILLjUriyF4pbnWU7y3knyJ0jOKdQkQ7YDPB
/1kJsta+1mAlqDCifiQsv99EhTmmsm2eDJbu0wrAz7eS6rfw/t70DP0SVLM0e9a9
RReWKJOM89QG1Y1Ct18uZYGoCOOv7/dAhs1eZGIcNUTJfkaGtqA4p70/HmrtHh2b
YMrdz7iPIxM44I7MTYuP5oSpX1ooRA6dbBz9yvLJmNTr/pcnyFSMzYq5RRDh/UZA
y95nRXJs13ByeSJTHQPxUcBHfDSQIoPWFqYMTDB9dACZbH3wd7e1BzteTN6YF+7/
Lebofste4fgDzQZm0fmIALSwVLZ6/gJo6rDa8Z6N/NpqzTI0gjNVBugWrpW6Ej65
vi9f2KdY8LNlUmUACg1NWz7wYvxov+xUvLiuKNjvOhMlMkxzAfxclwYmPgb9u/VW
V3/wp2ksN+7rwLX4RJiLWIycb5NBCe9F25hhVxVsd2adoJnMbOgSUKVqT4FiBaLm
24D2WmsBjE5Cvlyxqi9S7Bkeatyb5IDscmtjG31RVH4uJGDF7P5kw6NNN1pSj1mQ
bsTRuIIaQrgFk0aIanKD2ugbNSJhl3DdxgAcCwG8QjN7vNLWczcBYF3HhrBzMFgu
1xUMavHWzE+RTZy2I6HjqB0EplXQrA2VXzhC5rPeR50QRixO27VpQcU6jgM7MHfz
PBpZ1hyVlsufR5z16ujIBiBnYGXxTcw9cRfQhJJEHw0+ODfQQFgm7bKP+MfYcctm
gR18CO4sTY3UT4WS3bgAOqyb9YPrGr4yj1lnPC0F4mTriofnWhvAX8bURdslZvcm
i1ZXVH17+rroLUDBYem7ZEq+XLXk4cNgSIrH90DSh+EGgX8qECQK/Fio7BLjfLYQ
BDchIYgx3GM+sFE86POWTgonPC1kdTncV0WBsPFtvueJEYZSae13quHm7AmKPlX1
Ba2946iR8mTcjdTUKxBO+5oUrqbnn1ku5hbO2qeI0EHr1pLkiVhpF9b++zY4p0Gy
PZIrn1tro66eakGmx637lchY1YblqDUI4PdGL8FUITfD9sBs5t9phvDu56tTnNad
rsDBOEfPfQRNLA19dYbW77BTrilr3vQTqVzPdoDDrZKPL6IIVBrBenWEQEQOpzLq
kamteaPiOzuwTc4+qN2RWQub2pxoXp8CIgr1jWYH3ubEqd4GofbXLv+6Ey/qqVbY
fjqd4XEU92OMIIEiT5bPghb16AyXJamZYROpyDimSOMFVv2+lsdfLSNZWl7aWRRy
qbz16GP67zaPoBxh2iGKWUKnFY7es+aZrlUMKBRrYRLl1ueEWfkoMbC1MjRh9Q/U
1orDCxM18/DEgjVmSo0SaPIZKVy6Y95pUgOtcx8Z3DlmlJo+Mev0rWlkSLPDluoz
cqMjW49BGADaf5WhtShfX7MahQjw2L/SvCOjj9L3ocXIiwO4OCFRjZFHb7kzgcDE
2VelJm8WzQAt15SQt+Qyht0uLsZMt73TxknL25/uE02x/jnq/ARBs/oozAbyIca+
DCSNSKNexXj3KVzN1i4VTrwI5V3eIJRzdG3hmwjtMs/4oUVeX/uh/Ds8BIh9TW5d
j5ukyCzR361i/fLKW64w0IHJK2JAWnFpucsavVpOA6oVhJG/d3alsBWBgPk9T0yb
bPYMmCQLvmOmgbOPjJNPEoK5TnvjXIzssCV1AyULXZcb7K8pt5IhQQ47loeBKqt+
YTjkgEVmZtCrM7pKzIXryc32wBt9zrHmscA8HHEyiMwpfuODifUqsDURk2WW8efD
H93pdjCisnuwHwDInq+N/yUORDD92okPQ64YjpGdRrOAHtGEDhxDSYZuFF6dA1qc
swI98bH+UjJbUD45UHfrblIeJVY4qrd3NEJAmrKhu9pH5qOo0pNHGehcTsqtF9Gl
ZlOL+DWqSJJvoerNf3Gutom1dY67CKO33acWimvtiic0YJ/6Npu0QN3sC2Q0S2LQ
SIC4rrpGij28jCP8Zq07TD45Gz2xDo5HQ1mkQosDfTbrBZAlRI9Erwo4xi8YvBg/
o+678RS2irEeQlREJuBDcSQAtRLkCS1l/FXn9aqoXc2lIAJnugGeq7xoOAm/NIfx
FEKQ9Htt5h5elSLZ+6Z8VIm+hA9QV25GNtq8e5Ed1kmPftZJlzIZEdjEKNJSXF3t
5adHdnNQpI1Kib0hy6Mu85tSO/z0/AhS7Lb+uxVeSJfqcJohlvsuKOs737lQc7HC
J32JOjxPXR6t6v3xlm9XEJEAxNfM8+kuqK3P54wS5nqCqfq2/FWPOamwyb3TW3QC
H9OqOPpbsd5yMoEP1CO/OxPK4BCegIZs7DTHlWiobRuzRHqC+nhuVNQqdhhu5ZCh
dii3PI3EsDhwDpFlOdPWv4Xrnm1QuQ3UOhg5agLZxKimG5C/UWNShDEyGE6v5KRO
B3nxtGSd6KKyYsZpCBUZe+OcK8NCgoPXPa2ASHB3pVujBX93vThxSrXVzid7a1/H
eOwVCVgyGeadiP5Hhjwdvdrov8gnpkaUL15epXpioqKICZnoD0LRBwyk5W+vBbGf
Y5xD7OY6nWvHqhqn6YwrS3Jv8msuSna4Izm7L/Avgfomci4oTgwrF7r9L+6cA443
CikeSs9B9rza7fjjO5pgXG4QhcRbdRA7CyTTbnOup2FAJ5UU4WZOMIGyEiJ+AgOr
on9db2kR43hSEJgE0n/HpxkWvM8w/p3/2XwMb7rxgWzGMXfSJ0/9hUl+hz3mwp3O
wdv+z+PGvMRsKIWr0z0O+NRiKbPipqAf/i32K2SM9YtrK6eUWZzUdD2dXaDvy2P3
OBiAoe3DCavtDwjQLy4QZK4bd37v9wVcvy77KxLY71ibNnlBQiEuZkRWcK//cx+Q
fJf5WfYG/0+5rAANNrz2hs+68Wd0sV6ojpppcZcfu475GKcbXn9oVkzV5vZD/HrH
6EX/TCc6w4rs9RyEL5Jer/e3OlW3lizpypVnI5/fsnUm+6FA8IfakudJsvFNC/Nt
bSByMQZfhxXhPfYbjMjdaCMIpnYVl15JlXZrOv/nbFHSzvSUk04ABmKdPAgmcho0
u1i61KUh+6xkkPZSIY7b9xQqEf2NAEWrddSfX0RM2uNgHGeyHbHaZiHg1bQ+U2Tk
aVGfVXKjN0t7hekKIV7mi15R9MjggLrWODPPeZvF1gFKjUZY4l39GoW3+csVQAlG
pw6/4TYwx2kvE27nv0789aMZ+28/xuU3yiEQq7PGHsQlRpCXJWd9dWQCqwIhHxul
g4jCzwssgPYNWZTkEllupZhC5DP4Rt5cpeYwZnIE3D/BcXejBYS6zCgSuyxjd/PU
oSdQY1zF5+9Q7kRWVRL3HPflJ9Y/cU2SytRivQGWXRgBzy83y+n1kozDMwBIlFXx
+9hOhs8MB4QzndzsxpLTt3/s1ifH3DhnhJPgPkuDtukQBgKH0Y4K9mF+0U/8Kbso
WvRxocIwDtkjgI4IMxRQ4WhfkY6DkApsfSIOuDp2NU6sPNibwmLarjW0gy14HmnC
bdvpRqwyJe5wkPdOpfjv1gcfMMON68SyM7J9F/UUhqBZ6HlfxniVf+ntxi2dICM4
a+GvU/Hcvo26/fKFt6DJE5f411s6bdvhTg1g8vV1CN3jCE8GcEH8HC22JecJOZWO
KewQrGrVzIj5e2av85IHx+E6cNz+eJPKLX04SOOL53N3f68RHiauDII15Vu3lgDV
TiqyH2nF1CxqY8aqt+MQXQ0lGet0D+ZTN+vPyduiKHB1I8AO/w4fAR2aImCb3SJy
whAjHlGVhilxoHyUxJUhQT+YnXwnrJTz1vOyuzc5z3aQTRFj16rCAxWR6O2HtURc
Aqu4O66nB/+qO4i5Q526dNLQNvOJ7bpnB4UV8ZC57q1MmsCHXJ9UQPAVt5tSNh2/
zUFcUmYCinfH9h48Gl7fx8zDperj97K1OJdlF7hotHe45Wed67LvAjuHt70hnOmK
sOw7nE1+AXTOqvbFu8vgMv+MgX4UM5YJT1AqLf3NuQ5KHnPEHN5MqceZrjEF8PgQ
Yfoyq3700ZQBalngNfLYm2f7OI4RNQOGQkJHBxn12cB39oMcVIVeYvnVGw2wEtk0
9PvxZ7b4c5ZQKo/LN3YRVnp91d5qYOX5ZAGvkP7b4RopN1oJLWEGGYFo5UVNEeue
Kpa4RnQhDm44piYNhoWaUDYYsAlV0+lVnLgwX43qr0Vwg7L3HxI+PkYiCP0KMIgQ
7JtMSeMvkfl1W8TMqIrg27rtc8CO2nyFtAhpbHt+y3gExCtmk1OTJRaqK4XXL6f6
R3sGaVLHmPyyyQ0YyoFPiySI8m2tsvALgY0aXhrvecDXhpHV2u5WKoaAAcOXhrDJ
oZ4c9nWVWTEo8fsc462hzau+UDOPw+DZszOh6Deu1i1/vqrG9LgmjHnVpk0fYAbB
CEdiA6OzN1Mzr8KY/xV4XFxhtQezDzbsQ3eiLgnfzcVvFi4M3+yeu/U4POUo9hpp
kxmM0mMMIJRgIuc+MA3rYT4S+eGudUKx20+rSN0nXwA1NRQbhwRjCy6hU9dM3KaN
ngMH6Aj+VBBNdUrL8ddvaVHKs2O1ckgPb7gVCVitBNRfm/fj9jxRb9bc1nxBNk2C
qFIpEc7i7ctIAaaIzZY+eBhQQnrWq2O7ndtlOslEcBV3QsuQnSOjxyI0zK/nOZ4J
a2HXoH1XgswgPg/NjISy6JBerfGRIsM8NTas8+tIPpsypO8oqBEVK5avDSyIVLOu
naWgE1xAcv1jHsIhy/d8PuqHIV/nh9VlE6c6C5Q/u88p7KULdwAcZEffX/7w1hfL
5wZaQ2iGuyLCNoyvuLOiGE8br/FcJaF5aFRtPJNY0B69KDdoHJUezOnst+AHR8bk
PC9gkxImp12QQ6jpwjpVU7YhNVVTWKzSaK4DYEXKOZcjax9Uwp2Nc9zx76KwPsTl
9sYGahPOscqTSkd2PIb8IO92fXG47KDfchOagSPhoiRPo6U039rFm6YjR0nnOskO
ok05ECP0vpPIS8jr36SLUumAggkOlbdwnSJd58GI4E+2Gz10BpIGkLSh0gtqFRve
vnyIjtucgNyPKbFpVDO4TlXIW0TMdjROUvCJSjJ7L9a8OnDCgtsNl8jEtyKG5yiK
0NddZaI7M8vP/J8ttXHxcjySMqOpEAnE7H/xTMqkg3EXwC6BVfUyDyEYfZ5nIjUy
EZrG3aS9YabjfwSk0ZdaT0CM7clsC3EIPVLdJdo2aQZR8vx/ZPs9W+a4OhTU/XCD
QdvJUfNjLtTFBRZ7Javaq5cUxjjaJVRk+GN6pID+F6EbGn4JjYSEN3EzbJo7l3hy
eLnFWLTskOr5A0LrdvBUb4opAHzbyrwpVqeziP8oFJdxUe7vXkzGeh2zITrBHY8j
H4cnirHAUX0cpy0hxHE25E1SLqp6naH0MhqEmd/bUXsulkoXGIcs5sfkseC7H/os
GALc8+N7cevdVutVLX1aVUz8AHjNbz3anV2CfzfL/yqZ2QjmVlLOd5PE6iNsvqWX
Q3TlZEBn9Jhq3vG/TcXys8yi/DYb5xD7o02iWIREke6x/RmiYX0HHMELg9SdwdaI
odvH8CvFfhlylOtfgR9pjchmz1lWYsqRgXx4dYyanodNCHP1mgz+hmq20QTXnPvF
M6t4pi5Mx+B3ZVqUqxT2+QGAEprhDmg3IgAy62Rr08SPzfTlE3KRH7m/8XdbNmXO
kg4JfsYAhCIE1uKRPDcVL0OcJzKPmQmqnSbUehi1kHWKq7M+pJbES4trAC4ji8l0
U9DBShqN+Gg3ENk1i02fnCTDWDgjPR6sj0Zmsm20zVEFSJK7IAyz9qL4iDueyb/Z
oBVziV6j4n3tN75DU9Juvp96F5aa7Pauz/aHFStYSJ8W4mDR8+eG7VACWUoT9D2n
H/dW4UqBgd6uZcQk7Xn0XoN3W9TKuWVhkinAvJx7UkXAI0OAn7Cyqvrf1b/YMB49
oPil7m4/PJJbsbxJzYCeFYnrgUb51xu8Pn8aDbJ/S4IItuACFFhY5GBn/nKhUWMD
Nw+/HPxPpFRgE5fDTEnqyuErAtJqVMlpljQ10x7l0y+bXQIimMAnI1TZNhG9kV3f
YILYZ8mFYipPeN8ckFF2SMdBdLRM81YEq1blu1bVjUA/8I5VGbIhhlTAbOgZpO1k
3+5uwOqWj7vE8jTkWjM/lrjCXGRjOKjac12+WHslKNzMQeqQghqiBm6aXp0CIsGS
EZvXX+fIruMvrTbnm0RqAX7Fbxf8VDDB4HDkflQRpaLEKejdLXoS0X8isQZj3xEY
WrVOMw6S//5xgGj9w+Zm8rcq/ThLG2ekPXeVwIM/tVMIiaDdX3/fuh6CoiRq2ukX
Lbwd2kZQMNzEluAvJNb8t+TXe5TdsiFE+x3Hg5VKuRFJ6/kDnARTyo88x0aP197X
FsS8yT5kR8ugAPY6QEZATaevUYjsHkKld+nBbwcFIN6bOsxjfB9R273PDKUC7eOG
+OwnVOJ1KXj31c+ZJmalIG0YRsGZXLD0UmaUkz1lKb2D08qhLEenU4XOeOjUt34A
ox4tKTX7FIAfbv0MtNt9Mi9Ogk3pVmPSm+INGvA1I5rAcYK9aNTdGEroH/d1pZL3
Q9/lXPHhQjfHDm896RIcjBVbzvBUIVTZVf1ZLvIiB8fTmcMzN0267Y7bsQBib66+
xQEOGEw5Qu1l07+FBJAYUK3FEdkT2XRJ2HjbCLbiqDfJ0dp+J39GkymonUBw7eFq
1v7owjDKYSU1nsF/i/pZJEH839CPBKa42TSGw0zUzgBbHXi6NJWfoK8dXMyTuoqB
7SRpfJsc0KA9soNJ2Jq++P6hFeQnel+9mA9yFHPr2Y/NpdwVTuzNGV9gPPonReFv
Kc9IdlZHHlP59dpIMzcTDANhtAgpU7oXs2F+yuwsNwrMg52JwQhyU824XdAL0U+E
MTDKYpgKwbJzvSgb6UDXkl5MeU/p4KiYmZxipFyT9WFnY0w/Wev0vjjt/gYhO4yx
QO4Mxxdom/IHPtZJ10LnJ2tFz6lckUonv69BvNa9dfsGNb07u147LJED0iWuvY9h
MWz11Gv/cG4oV1q1n4BavOInNH9jHiK/cDixT+mWkRgytjRGYN5wPTYLHv59EdPz
iR6SCJ2ppdV0h8+mYvDhW0hmDcEVp+qpuJDS6Qonb0i3rlPwlCq94TCqjkkfcEwX
8ryBMoO22eKieLSbKWGbW+OZkaoYA1VvT/RZTPB+yeQYjGQWKnphiuWNREv7UF0n
OHbKc45vsqwn8O6zANn2LiQbV3Z2P/t37oSSWvVtrK2g6iDMZQ+P+Ye4jyqOpqTz
W9/eBGY9cDyFeM2TFxvgFfz6IFAsATkia/Cqf9jfESHwQPKdv+qmE3yM/bu1h08i
i2kx9CEYK9OFuS+/yOE6cdVxgHU9wCFH6v+jhaD7fAQI1Ec2p8fjqUhqs8yBIkO0
x3rUj4XVVJf9YsF4HtV6OtX/uY/nfykSXkf5IK8CABsWAk8gRBkCX5z0QVxYmRt/
JjGtWS/mslVV+bJdNhAflz9wz2GsjHT7X1QClLAxja1mat8aiVPRgGMwyzznVhm+
p/DT+rj84bo8UdNp2MeTrrd//rh3zJaQiUkBjY3rRCd96GYRh0RkP4hm9zzrlsKp
fUmR4yE8iMMy3P2WBiNQYNSbd9sZkEOcPCHh+539MBtKcgA5F3nCTYQmcy6WJlko
oMhk9MIiVK/wzCbxeRc+jaqykHtCrbgWioy1O5RlFHK84t41fscerwzQ/7m1ISUN
TWDI9UI6pGPFnLKmlEy7m672MAOgNkvXUzox9EKxCAC7Ox2/0zldSa50GqGY9O5V
K0ipzOxx6TLCg0NUpaQO2kEa4y0KUw6gslN2MtkpHiwRJNgG1xbG+KrKKeVUI5zP
YMAMXBhqBhb7ULslL5If19wbLwNoktqZWsCHIWs0WgO/es009FNSN5LCdTyJ3aOl
Wh0z4/2UjtPcYxpH9BX2VmzrnhKW6AI+oYY0LCIUC9AOz4STd0M1n+5Xc3Qr5fb7
BH15/iNVm+gGLq+1dPpCVmQuMWyCmnnNzEqa5haL6FkWPC48sNmFsh7EM3u5/AEp
ZtSNsjKgLOJPRz3a5s24Lo/RU5Olr8Zj0XQwHB8GXcUp+j0+ZmrKJfiZ4hK7Xi2+
x4ayO9E7Gc+ciUOznqIzbMXvmkGf7oiMvntG32LQtMQeOilAAK6B4aAogwRHz2T6
5qGuPkPcvCVZsawhT2MWEmGFO61KoaFqMesgifhBcS4vuBgkS3gw8pbeffOutE64
hQkIT7oacAIA+8i4AsMXYcu27DwWV9ZLGkx/EWuCI1SEIJ9P8OLgCnQH/1ofwGVf
zL3TutujBbZCPFrJ4wRU5Ntn0AseIJgiaDKWKZ8Itb0h+LYMJnK1Cj9dFpOL+xW4
9kdg49EUAW6vdJSa6PEeNh7G9DYOw5becZ+NKpPsJreplqXowEmSU5c5y2PG9d7T
a29Z/AJoXvTXpWFciPERLNr7xb+z00vvVmtqsxz21bzzsLhSeaIe1yJ7Kads4TP2
dz4wt/x24Qm5HsANtMBsSP/ALix5+A0azhBkypJ67BoRwAZCdTos3TVHRUOthX4o
5tXhp6/fkbR5N2nammNOJi+VSdPLYrlgNwV2oGultNOP68twpLygnxpg9AZLAVg2
BY1X54LP/LH/3KampY6Sx0/dzLRBjBu6H2XAdZzizdzWqawHwGdpzKPRTK7nAfgh
/E7lRaFNQj04RTa7t4k2TBose28CLOVp8GSmn03GBGssBCEU7lHt9F47OWhy3Qfj
ZkB1LA1gwtTfx5vzmcd0PUsO8t8aIAXChyzSuXqta7QLG/BSKHxbaKZl4AaxqKfo
kR4If7AJRspWV0Z/OzAg6WdG/unswS7+ayi90h+fMAab/t/RiY1Z+augColhCkEi
4M55IdCj1am2KFQyLzULV/+VylLA75xG4y3xs9HmcMLxL1tGZZowBSpopflSlser
NwA1E3wuqjJoSaCazljTB5KNEkUPpRV7HCsQ8J62IVeGUNSV8eTpOZMmMSJMrsd1
cUkNtMVB7kFwVDxAXscZvqEILO6Uw1Q5cExyLSSMV1NwdqabF7EIOVchPlUs79l3
9z0J1n5nbL/jDkR2ZLXuNfW01WUMybeZ0inkntQqyaB4MdwTHv9zDhh03gsWQFAs
ZKbKp+mHavPNVWk7qAN35jcJY5urMGwYeevAywoJ0ovOu+I2hX/imTKsOSOgYPcp
WedAf8Y33NoFeqzAdfhiQ0S4lZlnX5NvBfBknuy+m/umRpk36etOWCZdPJH6rSvF
0hz9mdDxeR0hdLVZcLUsAfx6mc1unYhY8PaE/49E/11XceqwAJ6NixDAZqH/d5Ye
FIy4nJ/XV/jnb5FEzuRHxStPkrLBkgjwCoEavxxaMC0kN8VblT1J6I8wPzXVtJXK
2JjvvAjhAGkGOaJ2BGw1oDYuMllYqsY0hZicqwNWGEaMer+99hCH0ZAIRs9HZX/B
yNvTMLN1COAvjCpRpZnTyNb15kww49f4NeBBQS/mtqBISNCy97O7sYhrBtQg6VnN
rnnVeqDklwy4A8Tmk2chy5I68XdD/a5uXE4ANswrQy5Rfd1BXmg3R7QplEK3EVYI
H7jvezMq9IPGJJgzBHw4HZxCZWP00uVRmVgC4r5mFreWmDUpb4BWvJYoz1T3uGUe
gmqxLiz48SOemqXtUeCHDiUH9dHF3RJ2jUsJbr0WUROqLKeVa3W/4PbkBKJRFZqd
SONg5f6GroUctjYlWiurNKgDAtF5TcKAEoLS+aoYt7MQDpgwYxhnVwcVwTzzPVvY
BhiNmCwQO0n8Dzwq64a4i6mIz3sR3SY/9ZvmGtlgxBqGVRsUplO57XfaRKsLQcox
X9dJCp7uFO/BfGDR69f+Uk08xbvcEsfzXGiSIVFj87Y5+SMSWX4TeaaDIQer3h9E
+RtTEqr+AMriEvDVvdg1a7EFw2rksD//6vSw9PuwaO3hW1sTlARNbPwBCLVXQbue
/CBTwnv7ClAu6rm4ILBHdlZbD6DjPaBfvaRaYYML5Yjv1dA+H+tTs53/wbHibZn9
BtpPY9/75TCTzdHqU05zhWnJ25yv7E/BxswVTwqMuz6Le/HyJxbtG+XrKHXgfh2i
FiJonBC090NN1x609LDqorXZIqFQmQgwuiNK8DJS2afuudTSN3rxdMIDa1EK8jxG
oIO9pAfs2Yen75+Lr+CRH5pbTPpieEcJzMZwofUtg/Px3qcrIg9+OplzxxIl7+FU
wxjdik7bwgW7TPb3BVgz3zEfxNjr49PeOgUUcPbmkaR0U0aQg9ICl5CiShUgqksX
byQD10y4pwrK7D5IQ7POsIdSTPXWKYa+GqvybpKrGc8fzM4ra2QD3Y7aX8ICyxOv
PWbZSoiUJvw8dbHvRiFlRwDP6AbQej67e+n6/AwdsPM0YKtcuzTvqxnSW/TGtxbW
x3BWz+7B3Jx4+0NvR6qMrCDbcFz/sOwr0vcvRM//JrRhIbPSI8LAWSP2Leeb922v
HIeMptCHX3RYbFrav5clgHqmpGKMbIrgOVudgQEVdlhXV3KwpYq+8QMf60mTWa5X
hEcfhZTj2lTU66yL9wbnhMYysVWittPalU5UY+9TkJtjSFRV1nqOW9ztKHzn+A4Q
XRJxUJu1KnJeKeBpFegPAe4U4O64t6zlSEUeSwd42w6BOWrRY+uwEGgfkPjb9hYD
FsK0OiVbd5ErWNM/FJd6vq8lT/oifXPC9M7ruxhmXsNmFb00XoKgxSeKcB44J219
2TFwjTklYSo0iD1qM22QZ9ISWi+CzRvBCfvS7TDzJMCmSN51ayI/0JaYP3UD+EP6
v8jNAn5mrnfpPo958y0QivMFY8f+9gcgMIG8IInrzoY12Qck3fkIDcEsvETHiVTb
KUY0SOL/LuFBp1wiiUvd1q2BOwGrTEKBmWNuy+8WdKW54PXNVU7duDa29RoeUt30
KOYQCcnVq4wTv2pntPKXW2LaxFJa1dGPY0cox+VkcbmumuurYACY0o9DjAUcCsHV
bWzGEFQGn9jKrdADNts8enJ0xYYKBYitXS/aqjySToWMekOBJW1yQZfhoD/D10/7
eXPtdkHc+niIDkOed1XBmA5sVL6+GGjLZiNGjcR+8jo2D53ec/5+a1Io1fYzdEO1
HG9X9yhoEoSGlHQN8n/mnJ0bNZ1ZYmU8ZDaBfhuNafLjUvm1mQrNCoS5rojgJsTh
pYePUzlI98/c8tPZ56cELPwq61HhlSgxRxJKgO2YhkK7OR4AFEw/J2q9MgFmfKql
uQq2OTEE6h3zvvmCrXvVqqk5VV8scER9DcCX5eq+qG4GA2IUSKB/sys/vUhEyQ7C
rro5NeH9KZyEJFMEAQXMWhuQKnlemJZmXBk0MYs/uCHJM0CvNcBuHeBPdmy4b4uw
mKcSIK0CVWUYniuYmT2W7R2brVj8uYTffAerLqXFBnOfrwQ0gmFvvQk9Re5LxYBg
PKtE3+AEUEOCL0GEcxZMTiO/1NNr55sSmczJWdElBhXT5jWchsO1dRCrrxcmm/FE
jyCS4ORiEqJ7xwE1Ct8rol5KzoyjhNvp6QemYCWbQlceZJ3Wp/eFz4fQdPWwVmfd
XN2LUUE2ezbANOgso0YWI7z0UD6k/ziB9SPw9R3bk6Bal43T4udN8YmL2Q8xZuWo
RzVi6DcFx7Zo+9vTX76UKzl4GNmR1iPNNgW3A3jso/5yupTjWYGyGYlW9iqz7jem
p4cDtz9qcUUqeTqA8aUnZc9zaJ1PFQmnMMkep7m1vwkoG96Bwwq9RayrJhAKiy4C
ftOs9v3MChVIC51IZh+j9Iy/TJ5ImUrzAqu8bDMCG2uR//rswSGhouuGfIENIILa
fp5BbOHEITN5rjMYX2hpxnpDlQwG7urahSQ2dcUjJnQujb1Mf+NSrmnRyXKgFkLu
ZlLhSXCRRkjy6f7HTyfGA11QCRLeVreL5oLkOWJU7lzKvvXOLPrxNIOoxoVagOMM
7+Fn7x/jia8hWkSFhchu/HyE0oT/Yd9qMFOxVSUHWhp/qiEAfmZtkKFXwgGW1qbr
dbkh9+hyVPhBQn9PlNnlleT19WnE4/avx3uSzsZrBsoZHIkAVj6mSZiMOoxvfqVa
wihjgXoYCaSKyNlAlLvHewPE/UDsZvmBsYzfn+njQPDXja8Eqmn8ZwVBBDHOebvO
FFSW8GN51EJQoVVa/qshUnxlRw7XVYA/q94O1xXdVWBZPjH5bo0FRZm+rlWaElSv
kkHU4YTLLDnHOQmkgiOzV/0xtUO/9W8V4vzNBKyoIvi+Q3EmeejerM2CJzwlWP3F
U2B/XhjBur/rRMhMgZRY9inrxVl1yUTPYpYgu+mpAUJE6ntSRRaG7Wb7S7AGZWQk
ehBz0HK8OaAlCJRqI9x3b638S4SgeW2CF37FjxVCbK8LriLfOJnnA+YeFv+Irs5d
aNDiEZpAZrryQBpxFQslYA9WEJcJNnQpaS00Q/rwLZ4uxLntniXm8e/6kSIWtxxH
U87tPZLaCb1VSeB0/ECYyI2eRKGRS3DnjsC9ECB2TfluUFakRO4FHJ5h5RUDQX6Q
tpqbhUQM87Mqggymj6fGJRKLshRssy+Trgvi4+qxJcWC1IyydFi97oGd2mt86KY6
cH/48H5uEKfj7iCK2seDVqB1Nozfxh4DxBbIbr/18Qw34siOT+Hi52hDvu8eimEU
79UunBvKYOEc0AJrWjZshPbolyf3O+5m45hUuTeOcWp08Gnb2FkJOpfPhwZJHveY
hFi0RSMkisVwRpsU6HJhj/5F5+B2Ck4vcE1MJMyMapHL6OjRguTJcan9JHZLsZ6K
cGYCsoDQeU2YFSHdHpCm4NAiK9o2okx3B84KqvQwShCLQDiXDmp3puDgvEJkvRNb
B8LEyeVBnR294/k3AlKXG1n8KAwDLYfJa0UB9ez54fv6PNA2w6BsYpn1JhX1NqQy
XsBzYCPozLHQ2CuXyr9ZBBhUzmrcYSSjwrwr6+9M+/uGlDPff8vHlEIhr94dSfP3
M8R8S9qrNBdSSI3+Nci76JbMuSi8dzV+QrDo8hQxHvP3j5ad+6SRW3m/9E+m1fWJ
S7xnfuYXvygBWOHZpEDelHUe2gWeor+pkz0vEEDjgzeGV6mD20nlTsZthsqDMbwq
12Jm4yJeV7ZbY6SqsOm074C12OVWZSmg8qxpzv/h/YP9PhCG+Kg1HsTtgZ00B0As
F1UnetvGoFIqUvVP0ogNNKoQ/FSen498Vqgvt99NsjLQgwTFU3P6QNWqx/Vg4ZET
T2z6bwVLB1LpRh8oJrG0I2YgA7dzUMzx3TElGVcoXI32rZjtywSWIv/6wPpYXuhx
9nN9FDlbRe8BUk62lywxRS8Kn8t5IjTu3GBFawtoa32Cee8dUr0Ck0l1XC2/g38e
pcxad82RujDd082eovZ0h33gcqvKizjDo3z0K2tVlZERZe70Ycx2911pLOe/FuaQ
FelLiSF56Bv+Yeu6CKReBvcehqfB63ju7yxu1lr80W+adOFFcZdiZxkFnJOQlukZ
EJjVl+VxKezbHRzziMKmXY3qQQO74mxXzyvsxRZcK171Q7XMYhOZPgh/XCh43gmT
GhzKs5U6qstBPkvgbMxPdqiC3k+Rzt72Ti+lyxkrOToDo8tJlQ+lUoqU2d4gJ/EC
VuBol7zuW23JVYCTjj7Ts8aIXPGcKSRCoV4lpBsuutw/kPdGq0HpHDmOcrm5tvp3
MoSCqZdKh8ofbV40fwe1GD/99dD8W2cBMzPvLThQJr0unF1wwU2qUboW5zLsO4ol
jnUOXMWsbnhRKok2VSZXa5HUJqgTNE+wqnFuX1pwK3o0Wgu2Q6mcQpWUCFa9JEFi
R0ObNS1ivtEHf40c+Z2bJftak1sxoR/qspmfkBxYrIn5Wn05IWyy1wFEd2DRAN2d
BYARap1OiAlguKZ+V7LdJOa7rOHGW2jlm/eOhdXeMo9exXZDFVRqMlHqWDLUnEYq
vxqM/SY4ElD72XYYSjZSXNwF9E3SkQrFVqCnmoOqtiJRlMEQvTf3EGSg6ezUX7Wm
B9CZJM7EErhY0uG6jGUVgewlO/NdEvAauHhIGHgXg0/xPB7Iu2HOh/OIa77UtiEB
+ZWV5VdK5jqxIHzUbQa6E8nik4YMYBNkQh+FvX/sw8X8PF6ad0fMfq3sko5RSUPM
Ox9Pw0gsorUpmeL56sx2nq/tPwE8cZuoPjNanheyTWDkeq/kLCPT70X/gZXHrWEi
wXyjrcWnvQIfdYQB3LFjtO2PIlKXLHOngAUp7gMgGrHG9gkbHRATw5iz8BCYNWBE
wZ82UXsV287Exn9VWc9sICZjcGPfVnJL8s77WzHnDjv8Hi3iliK1T2PXPdppLodm
tWLT+bei0cEVpUhJ4tsFFkU2TUeo5mDthSoVupZfMtNkDs5zRsRunmrzUSSUxXjp
7HbcqyBP6m/EcDEcFXvnJDFbDduqytGvzM9JDBthDQLQSUAJpbCZlUKwjgRGHBe8
02PqPiLiKRbdWeoEZTpsL7IOUtNGETz98GndXZDRl3EAPsilmOlEKBAIqSXLn25v
SzrTUg8tTZqpRmQnSYnkqqaOs5OhRJurAVw2FDiy4VQn9s1BKaBq/jPAOZmexd7K
jenDkHnXW7CWqJ/sZRZ384DhpembBm8G/tljoiROcYENvF+j2V0YImjOgHBKTaqT
7XVJjPPbUmp2JqibQNIjcYKKxyxlQtbUyIK+aIyNKtbrkjbhHhaitEI1QLv2Rv7v
+ZJriXfobSv3C2G1wNSm28PjWPGr2hDNL36fd4EPoqxvGTMoaK7u9CJ3SYgyvsGh
qA4Yv9lwMgjJ8DQDoUEDlN6BQrwV5BfF7W5zybRfkeNU21SFGdJbA9GESA9Ym8PA
BB05Ehna71JGoja7rG18ddtElEHK3EnZB0PaRyKBOXWqV6owgf5YKrAysgQGRF6/
b5/trFo54vmzPm4HGcwtJ54pMi8sohJ//HkT7eS+1FkyfdQPyR6aMAV8LeGMnguS
OQj8O6073cnbI3KOtvXOozyj9dixjSC2bVVMHB43FHKKz/FxM0vLzE3Ojt8fTJrN
P92UVGqdILuwPttmttD3HKKxoJoVaAKfPzJgTK5h3AGpjmLpMWCslQG2lUVVZQ7k
G2xLtNXGYYT9S9bU73ZXo6oouhQYpHb+nVs2yQoIzpqG+4jk4x7+aNImFOlj9Mwy
UUAzhc5YMFpLBXrUxySwkRj1ZpwhrNKLiHqFWPqzvFB1Ayz3M2B1mxKTxWvshJUv
f2uL3gFZ9tF/VBC987CCEDVQB+AyU9FFRPWjKlbFXrcRu7vAdvkyRsCGNRfM17hU
265E6kjeOl8e2vwfFQwk3h14JuyliEjCZ5hp9CvrLnsAJYDhTwBdREsZTsfERqT+
v5zszVOHRw/3JCOaXREuDNZ4UWRps3mWlI52yTHUWV6Hh7wqSfIOyGQN1fxDuVDJ
orSv1AztCK4NdKLhB4T8TIhWLI7jvpFTgsn2jX3nixhXdf6kLKkDPgnnpi81VTaT
AN1HpqQQkfwQi1Vv/cXY/1/VhynVLXpgqcb7/zn8nTOfmTonv7OMkD37DoGJw2/q
xMkHAgGce5NYRhf8TtfecodofoKf8JHP+GC89adVh1oiayXgTSHs0ZZdVpP72vLw
5Vowxq6yrRz2fVF8alp9tjClP0dAdrfw3hQ1e3WtynIxIXD5WYZBtPwkc+3+07D/
hRIIaqB7vKzcSEP9fqnxmn/2eZDbJ4Y8Z9IQta58IdnUWg+i9teGS5vfZP51yBqo
cFeeXIP1L2IbdMInKitg57xniziyecZxvicLwPNpZaVv3TNS/CObc9eWDMp3sXf9
5v2ngQi/JNE0abFUJF9vGs4J8iDwzwlxb7AjjedCCxACjIilXw2ioXuP6J4EUhRI
PJfVGrozm58URwGqSHUAM7Wkqe8RZ5d95xFGnydR9s+ZuWEgt+FckZMrTxThzgqQ
kW30LXtX0ig6sexhZOy3IiLV3uz76ZYaORSfCuqoC+DVu82c3WERcCh1HO90rEBw
/+F1+nJtxwxu1JhRR44Dg1tfK3tDxTz8AApi+NKG5wgLzwL07J2NSfKYI1rDo8Tb
1i+MzREO2jP3MqF/AcgheXpWnou4qyR4WBCoBJQ9XveM7HecOLYAQq3FQk8BkhlK
DKEIUYVXCoII+2JrYO/jHXLsymXE5Py4UqjyMqVasXm3geUsPGGmKVrjo/WVQmpe
OyV4o7mTtSqeiXwc1Y02Q0NEelCWW9bjoc/jVanZd161pISgmulPfPW33ly6anQd
gQ8SWtONM2uvsmz85ayHUuXTUDH1ykwctqOiEXjw1S6NBhh5F3MTjVKH6IojYGrS
F++XY/TofP5e19kIctbleLj/1H0ncVhlzAG0Zd6NDY8wAw1pSbhfcrd+k2okuZVK
H5SkbpjDDBMu3MxqvyF9AXb3cgEMajRNWv0zHDb6p/M6HFalw3xZo4xDx5R7dZNY
wkjN4mffriYaS0QaI8u1LxD3sGwLPavnr1a92aSjR/9hpWv6GdTUzpTq0AQApI2i
aU5uiBIjLFftIig7wmyjoYsiejD3cCCQ+wxXUEQyhFy9I2RkifzbbFmFV4Uc34SC
aFgnccUq38uU9USr2JdUuF48fgNAxXfCMItPEpP7keGothDvgSDg9iT1jAs5u79l
gbfaatLLniwQ+0Vl+e1KOpInY5JEnRJOKSar5josu9updCEKPgiho7aJDXF/0z9y
8RNm8UyurMvJMb9Ydh4j2upaygmCiBuz/Nl2/QgB4YePIN0x8xjTcN3ldqwdEbBk
tTkP9lcoCFz0mhy4KBNqVraUdNllx3ZT5E1M4UR3AvLQ3wYSQYSctBnVAF2a28V9
xYLH9hfs+ciGBsIXmj3otTb5BoX7XggOOjspKrVUb1yXcJuP1MWQtgDu2f6RwbZk
imuhJXo1eQHEVpX4IEsd2Ojk98NWp/u5UBmeL29R1jeecGJ9eHpfY6zfpDiCXubC
t6OKJU1vLiE33tWl8xNoJiyZd4UMQ+8OqIj7LtGJA5KQgGat88YdVwjvPccksNM2
ekBYGcT3w0SUfGVtI7zr7MH1MAnbCR+MF6mmrfz0flZ9z3lPSHEqnI+58JAR5hIW
awSSOyIWufI2Y2OorsPVfGpreeZ2LKXPTexUmed2whz/YUDKPabiO9ZQKEG4qz6J
Eb3Vw0cFp8OqMl5xkysy6sbbnzqC1VGaamgGX+6Au3eELivTVPUxyxWYrvQnkV56
Dq68xubW4MmdQaHe2DBlvK2FzD9Ciw6ayiWCuCXhBRdw5Q0V5ySCUA9WC8ldl65D
ClMXiB7Fx+IQWZMVzywD2kgBXvVfaiktksRafWuIRco9YqMte/9t6g3JztI2Z62P
BGomLDY3+/UB5DGZv0zgglqmRYQ6LjaaT4em3KtfRMTxq4aYVU4rLZXWsFSasdsY
qs2/+xE7dHaMtWKvDUcOf35VP3xHxwbkwVOFDNIOkSyvNe1uD2e8089tzA6i1f4O
UbeNrFEVfM1dLs5CYFOUMf3qrtre3Rbl0430IYz0SFosEEROdsZBwE4KRNofUNPf
7sXJi0VOchjFCjr150v7MP2Tf08W4ZOF5OSOZJpCKpNibhJucQba0EMKiP5D+e8u
suUMT+qW1jwSQm9RxGkEs1lQBrvduFvwVJUmG8y31jiI0SlINR/1MKVQw+sLyrw7
UK6bFyys85CFjX19oHb+KTJASHO974SiXpF19CD/XU180xutCdk0W7x0aBZf7eg+
4R3vuhXdZkYhggUMQvnkeiQ677vA1eOWQRRT9jT52zvIZ0GsMG1hVztHcqHda8Eu
J9e+ig6jAX8ISP/oHWUy1DWCsOkf/yySnx6okdbcKxLER63AOXlHMKhYOnuwTvIX
5Bmu2H/k0xau24uij/9IBe19gMjLwmj5cGMg3tHf6qXinKRcOEN74b7MjMSt3Re2
IuQI+pSEV9s5brdGpQh+W1Kt3XiDMUH5O3C9t9RSYSYFEcenoeK/IDJuuP0Nfefy
eBVaQtZjD7IOJplvutdPouodXGUOfqIFZMv0X5mX2sOx8TCMgRdknvdjOwD2RR5x
He81LzcoEPZ/RS3VkpZbdct1O8a5BqmCKcsuhMidPXZo/rBzILxcX0BrHx+B2YPW
0Cyve/t2eb7NlEi2s2mVC63Dz6AXamQ9FXItw5KFqvk8R2agCCPqetjez6VGDn88
e7I9xuYe1DUqIx1KroDnrWcX4x4QGAir0eWs1ysWCItWPmfSdby79mEp64M69YtR
u/2WKLE0Us8YgI4r0RaTe4BPpSPMOy+95Q6LHFlznxcK03ekd2HpUrxnMH3NGD7N
b+4A/p3hMp+dER515PFtpKYln1kC6iVl1VXw9e93uV7w+8Nv+SYs6jHUphZ4L0Hs
q3Jy6tyio1noL8Fd415BjlQR18UvyGhhJjdOf+n02LYaFZngEfy7vYpbnbI6CddJ
HAlSKMRElfhF1HWuHDcmHrI+S41TOdu3k9CQrGiqwwLLC9Uu+8jJqZQ2/GuQqM6I
ygLbE+tEEL7IIZNqPcG69Mh+HWaPs5JOqQZ68FAUP0WJtBIFh+YbGnt6tTnWeSDX
K+w2CwYl6fpWVU2zALDaylktIaqxHmLBQ+Z3NcJFVZJswWHqAOTRHbOKIvhQoECz
bvvYDxUu46sw2GzuOM1dQsyAKraO9DRbwhH4lq9MG+qUhxweeHbnPTPiGVhGUbIE
l4+yWEPa5RBCBl9rRJV2xbt5299g0AzwNYEBi+rL0y2nti1S6Qyl/wsN/+kbN0zy
5NURMPVKmQDLPsxG8nvtrTrjJ+IYLec/oe7cKhf/Peu0CRCO0ZoIQ5Yk+E7Ut5a0
GONaKUhG+63oUnPwVa/O9FHwY407U6PX0E4/XhMt/zjSG+GMv+8s1ewybs+cOUdG
6DEl7utO7x1XyKo1uORkhawK1f3/Ux5aeCoZyCCgcMn1ChKopx013j3nGEu4nmNF
CS2PjKxJ5FkvTVXuLa5pJiRTppdcjBWtDRoa2tJ0d7w489eRJYLzxZ54szcR4dp0
PRrhAm+uq03GSiL8GEkvvl+vZKYQnQaNOXG9MCTSzydFkJJizk7asY+ww7X9/sAQ
7I3D7wH20onsVV3JGbPhBvhCNcUq5bQM4pcKD/hmSd+XyL4uicrPyIJAGK33i/93
A/41IHkX5A1+vY7wuMeasOlkK857qhPSxUrN3E2No955JI+i6elUiAOM7pPkq4J0
Rlqt+5u+9QBYUVTTzCdjaZBywEG2L9DPZhqfzlQE0CTc7+FPNPMeX/pZYSjrZjI9
NQcmF0la+ymmiJR13/XedN8Jcv4EhKwj+CFYLIA5rR/v/Ve8MjNZN7PEBtH3lGLv
D4OXeAD2wpaNV7Lw/otc0WNiR4CO1q1rMPjlQr0+HW9Oth2xzxlBDtp5YVyY+GI1
3LoXr+sK70KNxTfUfd9pngQhhDfrRHiUBcJn8vjSPVSMswyhWztNag4P5cGjbBVL
MG5zhM3xrDyUppC8ShgT5RJwdTLqDKrNVRgA9IU0clFkohaQ+XChv88s02EoAdj7
7kaqEq0Tjj6EENiwlUpsF/soFfhy3ASOMY1h8FG2ZmHjXlzLQu6tdQyr5jr93akB
IYauZ22lfdsjFsXecJfDeDJNZQvH2OE7SIyTkdoJLzrYF8hjOyL8Y4LqJwRhvY1L
mrqegAmRGHkd5csww0w04/hyyAVnj55FyHlecnVw0FZ2HOgN0nuVhVTNw/f1Vaxs
l+whJvw6uRGLDzSYF2UQqBPp1DAtkxvBqyYDmc7C6tEwQCle0XTL46wakcEb/auz
tHNNjLjOwyEB0V9dsAW4ht7fbY1o1Q/2cU7ljHYF1Vc/KcCSR7kGJhGt2pktKzlh
j96bBcYkyxwc1/uy34LqLxSkeVlji/g+ZjLNWgiS5ZJiip7IDHcG06Fd40QvurYo
dsi/f/iAI4MhpvEy5T+iYtoDloKtnyn/MxNFul+1keOcDBgBXozcd9aBd5dUEQYd
rutJl7PKsDzANlZI/WOgiss5CFyxv5UWee3rt7RbIt5WHvmQPg9S2yEKlXPa+zsj
hmaaGEG0fYWmpzTWNHdEFAITyohBQ6UM72C5WBXzNvkO4E0tifMlTI2K00e7SfkG
7GkbHSmC7ew4Uu9aoLMekVAMJ1b7o2iYrkPWq82GnoRXaR1NxE0rkZdOFvhD/6t2
l61SEsY/UqEnN8FZeJgEwK2qLWMRUC0pGlgFeWLyZ/IQeCThv5jBfbwl9g+g9eDR
5sEHNdCik5OE0NthnexFg1Xfv8wjVhsz4BmIGdVeYwGQu8/BKF59IBcdoDcaX8Vp
L8HdG1efcE9zYE1Gn+Ank4n5cGcQylIrGrB+A1OZEc3tr0kbFRktMMl/ETkGvdpn
4TtazHL0LvWpRp+9EDkk4kI5gD4+ecTPnBDPNvdg41RKVJ+IXI6Sri/9hK97MTuz
qZVI91KW4+v6F5PKP/fqS1bikECl0SquX0JvXnHAc+v0gh57fV+X9/6TcE5QA7ey
O9eaWihN+G7bb+ZJGDiasCie8lQ0RW/Wl+P6F6mTE7tNvoXNsP2Vyaussd+/tx5E
9t8uHb7CFbK0gNzADVJLLss+owoOPvIyWlxKhWPPlcl4HMBmx4x1rPlI4NK7Zqdd
b2kXsuPiMKlt+v5XvcinHWheiGuTBYW562nnFNd/of2MMjsPDRUEPmDfIkbEklLh
q2l0Nx/5GIsOCsuwUcNkdbey1nsj9TbrykzPTIka1NQevgy/KFniJOXjdKnymdKd
HAl3Bko9nylQzq0EYRnVeeQMJs1PthrQdwSSndZjheNdkIlKKNvdodh/6RaQf1QP
vU7whJKHzpG55vZitCkpPGbByWLRMhuurie5X7r6gElBiJwSW1fvGu0GiWTvGwwd
ELvL2fxpKOx2iMkbr9xG0kHS3qTLW4d7KoP5gXs+XRV3PVtSqOoiWPHY14pWUZX9
AVbvWkbaWirvl9X6uRwFjRZxoS436IJOnKX6nC2jM4a/pE7IlbGxxQs3TMXDGWmb
wIRAZORHAgA8XhifnZlk19CoB/BLw0csykckErg2/H8V/ScEF9fxVc4KSykP0F9j
0mURyx1VgvQAG4rWKl+u3KbT7IZ56GX+tZPH+CWbEFzMHQN2Oxi2jN/UvjpVO5Eq
dFLKYKNl7HsXhjur/QxXdQPUB+ioqi3n037H7vcsneixzP1TeqgACXq9tquEd5B1
4vkkiImCcJnx4HIGJR8YHWBK4Xx30mRA4exm9u7r232ZSWBz/m3wza8zvbkeTh4Y
6jhI1f++Jd5j/qIOaRXs1rnh8wUoS3Im5hi9si8WAWSj0fCRt3slAeSh2si9v/uD
Og939DijQLx87LU/eKTvYstlRto4d7IEkJEBWprQfvFzb1Hji+np6fc6S+br5Vq7
/QE7R6PlWJFhitkMZAHqfS/Ta0NucNvV3tYGu3uDTBxVj96vSDbPHqThSBLj4q0z
PkxNjHJmvSwii7cs1y9I78KHHWeH/v9p3HSN2jZ6wBF/GRr1n1tu6zqtRMSwYs1u
yQWsTRtiNU+j7JDdnR6dbd7g4VHHhSET8JgqrwtOcK0BuybYKemO1T/gGo3A7guH
MgWwwFYYe7Y147qerz4l/GrhwxIU4Ss+o+ESshWH6oQ6DNf1XtkyNjwi4zdB8qfT
nNYDIyVGOi9rKH1cpE6TnbhyStpSq4suXurJeYjhJK0pm0Xi1DlWVZxbU/PE2Hl8
65PbM9V6oCkXHadKZOCorDwbcFazlq8CfwDAursws+DpdpSjIHMw5P9+nJc10gnF
Cl8FffCgHuOivV0bLXwI71cu5j/32RVcxhjysTFj1P5Atsx/7dnFkvg0YsDFRMvh
SX9sQ+euSV2UPDvgZubYTMa+IY9iApKSERxgqvbBzDTpyIv9jULj/T95HtbmUO1e
4NM0IHiOpzFAB07GElDZQLNLigxbDDGXGvCCBhNGyy2+lTFVfUyK3uDuq6nQkKf5
/gDs5P9Cs3VYuREaViFySnCoB00Wb0LMJPNmr+6vpSDr1uV3fLBl7QaIcTo+1YPS
q2i1xGEyHxjzdrgb8EDrvjRKmmfPSXAG60kPNg5709aRiKOqxwWeOvv0zHZsBC4O
HIK04TXetl3TLknmGnDWhZflRoTVzuiS8Up48n7BcbiskdBsyblYLAfgdHt+AQQC
axYqJ3njFJsPc3rHRNUS9cS/lr4yuWTkTSEZA7sypXycQfwMewVceaOd/A43HeSq
QBsLnohE9sZmqBJoRgR+fSoJ0ft0dZWro0pWd/3rBSCTkQuao1Wcpm6S0aBvp0U2
EBVKSJ/F4yHfhXPUVVEg5w9XGmGsLxtM938z7NQ5kLvJ//7eBwSamWlLQK/j2Ztz
XNa0H/WDpze3oRDYud8jZ75KZVJfxxOHTw5ffs4CfhbYFoJ7ukLVDyGqQYPRekGf
DyKM7675ENwUgwgtTI9B3iBzUorHiI2HtcK+yvXMcKdFdBSkSYuXiw0iazKWbu1M
/1gXOa7h4JXNlqBhgbqOE7TBD85NNSc5vnav7+jiuoYtSKFZ/rZR7eXcxGIzbo09
YUwW2sh1DO+Zfj4k+RWLwusO9SnxqeNGBruKORt57b2fkymK9pJfUMTkfvN1HiE0
XMpaKCTUPQemFIygmfMZ6WRYBC5wIpLBf/Z+orioUlnIVlUzn+ddMA2E4QhNYvf5
Tn9NPNLikbAxWyht18jTuQxf3bbWLvX/lEYba0dPOfYwrmfgymNHEN7DqUPqwSWl
bkAqOQLnhQ4SUNGbbo1UuguoBxSC6OFxgNcADsG5lJUF+fGY+fMdB/FflOWQLWJB
ZJtkidzLGnvboTU7eYR8t+f8piVZz2prQAyoU61C32I2wzMlXmPsTdkJlMbjIWiP
GLKcMvDtG4Xuq5pB6CPAo/0ltzAKFBbsGUSZs/mExa8YaXhlWYZ1RjRVaGk6z9fh
AX6bdmUFPeaArx001oG880Nxv4M/DQ7pe+1N4dl3WNJtwSSWzZ80wQkaZhsYIbn6
9ZyUi0ch1w0sBYZVX1jJrHIJajjMjxZFhK4u2nqY59nOh7VIgvB3YmMOaI48aatV
QppPwPzStnDpocDJaIJCAssh23yh71jIHeC9+820OVq+iBzm7K6TgESuqlDN+IZ1
maJa4u7PHE5OxSgs0BpTKGndg6OjWusZiXDXS6E0buLpIixB+jRZYWxNge1Q8zzG
jtDVWuPNk3KWe3WC8miBdHWMrv21EVYsYmg4lErzed64sAFtotMDQawQ6WJEZrEX
PLbGTLpxZMYqzfFgtASgI36yjzexgEuBww1fHwQ6uW1CQT1kyA4AU4+YvK0/HhHf
WhnHAFShwab8Sdv56C69/n2VSTTsXvCS8V9NQihp9sUPIq7km5rXqFLO0kCm+AAw
8b9Y5qovGHIREfS4WaoBZQ3CUmjFRvDm/Mhqxl6RbVwLCul1wiJhBchIoBFyKrXG
FtgLig4SyPiwsb3OMV8FVgJlfNRIH8GrLGWx+uTO6PXAWvsj/tG8h4okj4X6oKE9
YWMdFim9Q6m+BAUvoRvtaMbtZQS95W5TTwmGEvvjKkmsRtKYkXFZcbms8vC6FVOn
KTpRJjW1wtv0MuDOpri/OihlhfvpKSh1e7kMG1Fow9aMSJu2SfKy1Qw2jaUiSVIC
YWJozun8SF+YQBDbQyl61mGOVcmS62GJlq9crHLPIAQf4NtrzM55IRY16z7rs3UX
mt/rqWsulCJp7O4/ib36W8xj2x3N89Ccg27DQTBp+dk8tiVopNOBE0+m8+Xt5egi
hrKs0z7ufcIjfNBA6UmwkVAG5QRD58g0i/MX1bbYv4Wh/LY3XoNgRc7SPNZ7qadL
ZdMVKmw1+ut+DiKZ4bpyf1UTs/TTzNJXkLgODByZvOwoZDSbrjlnDWFQqr7jO04f
uynKJ3t4TZhnst5kN9hMtLeO/DMX7q/kTwoqog5Ln4NC3y6LkeY/UmHajqER/5Co
/2BBHGYAFPThAxONWhH24mrYp26myim64noEKKRzORH1k8Kt9G/yI/nN9o8yt1eR
Kp0pGZxTlrXMk2DyiW6lG8dM/B2+X0xMcHGTo1ZruLGo4kIguz0T93zWPzPaLsUa
17Qk0iA5hO2RnJqJXBvXUd2g1rcNjLrypomvNzp78sQn9Tm0aPTdRL4cO7+HKNSn
AM1kKKHQClyTMUrbEMFFv7SByANYqF5p3Ra7M2x1bX7RHfc5nYP/gpj2SXqwHWww
fC3FN9ILaRgCrl2DbkxSkskYa15sIl14lMZkZ3XfBQO8PUfrqYf6F7hxwbrXgRA+
xsjOAezc3yCblG/Ugw7197PM/gnZDn9TuddKBuY3KGxH6Ad86/SQexqmKiux6PZU
EGNn/Tw/VxUaNg1A4tCbAYQpdVeTk024ToGc4J7qFCPEZPNhCJ9HAJ1rM2Tagmkv
VEqUOeq6AsSeLnyXDd6635y4+UbYi/acMqmFJH0vdaaT4Y6A9nRg9Gmd1t+C/TvN
oEhbWXMKfptariGVBVWPLF7Q7sogyKW+bxbNr0t1Bhwk2Fx30LhZfh0fIrx4SK/R
9/V6Rctcfr/dsv456zta/xZQWnTNeH5/8cULc2UVbgqCA65WMyNdY7pSK2Wp3L3n
Q+zXWyM5MaQ71T57Q2AuXFMf9FCOLx52XE5Ek20uw0TnKJr38809fKiomGgEC01Z
x97dQXCNMMVdFMZbyySuvQyReNBsGDEYQqVIL16oHo3EJcnHkC6KYMfIN0pTB1SM
8BcogP/+AkgDkHchUghp568BEIKTd4urWEi63MxwNUe/BgD6jb+aHCj/tC5LgfVb
462mfjQj0KX3cDwxb/Oc3lbyKu5sNszmBtEdHJspBDWtcJseuIWn1eIao3ehnpeS
D1Ib+n+VRHXCaeD320CKFdE7hFEBYJ23h+OaGoNin0h4HgL3l4t+9Tt/8DQt8z5a
W8QETczBueEcfhO8kT6mKFlKdUoG3trHJNT4213Wkm6k9CR0fxrm8SeP8N/A0lc5
1QSM7BPpNgU1XzTJkaEIXIByxqlLnRzYYY/lVfsXFmbXOu3AqZnQy3yZnyLBwTgt
H1RYJEHBjKe356mqx1zmbP/eVhvgzabwwQaZO7yfFCTD0UuR4dZjd0MHW9vdPCRk
rF5zVbzw+GcSy9Y53G1g/FEf8BsWJ4e4sxR58H++9roy3lnGUS/dbfCBN274zb9a
6zdUDdYHDFKbkNTY74E1DrBYGeQ3JOZHy4E+QSUpUeQZwl7DWASCcmKhNEl7H9X5
+HKTN68lniY5fxxre/VyK78uEIizf1Q9tFmxnHai/DD78b2FY5qeHaasCkZpn1Ax
XxlX9KUhW+VmP419PR/nkBCMojM8vtztUsEGRBYdQst9rIlJLYw3To3/2ZDnl3zo
Ah2dnOPDvakqT0/OjuTnjVtJlHSltiolAJenkImES82Hi6+Jc8IqbRVgOBp+K7Su
Dqtzj+0BYjs/lkVVUip0uIO6smsduDJmzw7Xa2kE1Jl+/0rlKaVWCdHqLshFHTnG
gDFaSHrqUOSTTcRMcVPOdszMKMiwtGe7FYB8IEeL7hEanfn5/yLhx10Q17BNYgAL
kM239XW0tyJCLnEl6fEPP+Or9DEFNqLwEmuitflG3oMOGg0KUkG2Zmd13pUC/U83
09N+u2O+6kT+h0t9volsTsrXkjj5/88Zv1HInKwymbbZIlJMqmf0uJV0PE2S5Fa9
wHYZnDO3rXpHo1saW6yqGx/eNNrmx5FzEf21ksGYdBP2Xoj9+i/jaWSi/L3FQAs8
Nl9+jxwOz6mN7ebAPVq6DWZ8HUa6cKSL3I6GXYmur/NNLZkYY0FPTF3dvOaU5vZh
hMq+gAhyHLTRLEeRyWnMowwL5cYv2RxgwA7E4MfBtXt1dsJWn2s8s8l7RsQCMZOV
W9xfZmnEZSlo5YfI9tpsxfjniZNvLFtlGP/M3jCbqd499/jO7sN0UKfVahHERyA3
OIhxe9Ay0fg3Ik/T0nS01WLTBxWCpdR8HqRsWXkfz/+l42WKsbyOzZdZ5RBDtiW8
iZE+xNViu62E41kHJpbxAAUI+69oxxUF8dVZPD6Wo0M5yz6/LKFGVxaVhxxNppaz
Frao44K/stO2EOwagNJF8xZD7J4kH44SD9aH47WOLsCRcyffYfD09ezg2COVgH2x
E8yx4XxdtV6/Cc58I6pvNn30Fji9ksx5gWvXTra+lwNeqlK8NBu0dTt0V8UJoMXF
SahhXesJRWbXyFEdDf83CU9jxtIGds/wgXF+ZpuCodvHT5IH9NL4vYfcEFV9cQAz
NinfysB0y8tqCuw06GWuKE49yWwikoBEW4q8s1bWJlN6a4IeBvBGw3AD9tQIG+j0
BYv9wjWJjPJM8vXq33Yll2k/QEBOMkDu6sIuN/7m/lIzc5s5RC9xk4aJNpoinjoV
ENR2oYwrtvove3u/02/zYO2SQHf/Rtq7aT6ZEaMzcracVl0fbcefw5AEB41yy23H
HMKzzWgiInSZWwDOiLUYtDH0x3o8ozHjbMyFkPeVCTJO82WRi1IAily+JDYR9ySI
+3bHvds5TT7KoSmGMihC9aQxWaUzY7BWfXycdfd28rYvJRJmaEgKA0MMBeb82Nca
go3BEFYUway1LhZz8/ES5XjuoCyq0tY+7bmFgQ2wz9DRiDZJghh3XWDOW3vSKMwX
3bM2fDpkSl/FqjUCyFhSuH2cqF+xvw2OaN1nm2fQP2fQX+ZOw/79R+AXU/zdf+9C
LXBEW8WPUC49kyeVvqX0fC4XzBTV/kreH3k5MZa/Z3YSZp8P7UwIy+G6i67hL5/8
RXOhERuDZA0VLSS1lhYDLjG6CLUYsN/O9ZyXD9FWHPBnPHaxr32Kb+OQctcOj49k
AuWf2V9SM8x6tdSAHQVxMRGjSyIGrwUz3afVCfMXk3aVqI/edXMyqNAo4tx20Y3M
r2dg+rxo1jk6ogu6TbJCilx9H+LDuWh1Sd1JA4vnyVPcobrAJa4ueXzivfEn0/30
BewE7gPVYGPzeExoOra7TtqcEMbqHZ0L/cwJKZrBiYHGDGpoQb8Pp8CczX5jS6m6
g933VClA+R9L9lXCXM8MwUK9aICLMD6py6aJ257mjbHC8qRWPLRNbvzDRANOoQLT
G1veOUf9PasU89unn+WNFkgEYV2lj0qiJLdh/+V6UyKcLSaKWpODZShQLCE42bGC
dvmG8bJ1NMiF53SBVAbaG6ALLqamrgIBQwt18H1HHt7QWaWY8HFzaW1bz3vUIFnE
1ZdgPkYWaig0XkW1V82uQealR6y0L5vJyaTPX/Qpy+fknxYoiBxppE202yecI/J3
7yI1x6dJOLriwW7FGcrPLv99aOwttfdKgRou7mB4jJ5nL7QA3umkE/z+uAVWsIgr
t88Mxw8yjpqPTqGNvD2i0BObUdi1Hrgf6vSWLXoFlguz7UDPHfgOvEZVQJksFbLo
PR6I3o+NcXc2ZgGXWjeSc9MCekiVSCB+Dsx3VZVd//qxu4NdjJGyZhLBc+UP98hH
wJPoFJtQxaYNqb7SR8DrXgiSNBExHOCCT0GZqOcD3TIDWyQ77f4l+L0dWsa45wQO
nRTW1dDRHVuYfEpmuIbRB+cp+t3Q1BseG9JVa/PERlhFSGNvEVOsnDQjPrVkE+Ta
kpvbIhksF1DLhrG75njbJDSSJSXeXZ+UuYuOXTXseuhVzN/Vbb4ammqS3t2jp/5a
afOY8fwIchrp02JhJahDVEr7YHJ4ac3zK0FWsG35VWCxntdGep9kkapOowPgaH0h
gqer8YM4w6wjtQpEyjrXKFPMXZUIWd4Qbu3+7jyY8oV7+jp8Aogni5EtLdwhMren
FaauDL/uKpjLc/YRv8NxJ71qSTQcZU0C0u+gd6F6MnG3P3yR6aIvSmPi3f4eTjuc
xAZyQ+rI761VMFYmcr6oCZW4FJ3/jjOFZMmU88KZp+z9ccq9qsw44CQrBV/8Nhv6
MymjCDi2DeKLyowwIKBVAGzfAgCdbSxxbFEuK0DesVEa4CpyjZJdL8aM+ILJ01D9
A10h/gE2wQCN7tE/6YTP/Ztr1gS5CiqbQuMAGE4T+4imU7L6EEkFdRLvVe8IKsQB
oFTYEXMh/bNVwnfbQCyvto6TN8j55tYK4Vz3YPhQWhnMKKF3luieqSCef2T4eqaX
eL2H3O70RzdJSqgM1MLDHSaVCClum7sTsIFXVl9Wjh+ZZm5mxfvyJ4Qc/SrQYstA
dS+i9xEUENW9yZFfp+6kCYMvXWONhFa3u6s9VUtjWy+WOqnBdFaaxB08V3mCUwFH
bjsdCHHxA3MmzHcBWS4ES4G1JgHnatbveV1tdwClxcQu97zZlmbkP2vfU6T/9av+
Bodyff/CeyWRw/a0M8b3JPD0dKMRKydoGOJ68fCim3B0xWDzPHq7C2cd9u9D+5FW
xBTfSeKbbeZ0fYc7TR/ZaMaZP3xFFQsHbUlm+6Thog5kXrJvFH5kdei/k4pFkGmo
df310GsJshiKdxRuNb9splBW0aeRuUIl+Xy4uP3IfCE34nIk8TNcZnMq+yUjHZam
blc6IMw+JJwWDcak3i5g3zGIqnXpAklWSjUDdtcRwI872GsHzuU2WyoBhbz7qP2Q
RUNj/EHNh9BOCD5QzKA7KnQrgEEXaaQDDhLZh0UuKGRS5Wq0w4SDIaTq8vUz8iPK
v366x6ildH1ucOVYhYnyi9hdAg+NJnXFAjeWGeX2IIpAY9MDPhluoncJR0NnNI/R
BgiGbHql7pgW42P4IB7VAO/3bgDKvKB6sHOjsdiNjKwRitZdXiax1obZ08XYRepw
OHF8H1rlNXJnij+VA6EsqLGNMG8PymGpUogUyEYWcmvsj1UbGR9Lo5CYk8qDJhOz
hL87Ln3Tk30Edq1L4SIarPbHRkrqzDXxCexExTcB9UGUj9nwsihiGXixOGSSeo/J
GCxNWnvKPEgK8R/iKGfDFtMU/56XbPTWjqgCX4XOD1P9xmiA6/ZaLaNYewd63xT5
Fq1IvIOLbS20DifjJBlbuy3iR2PwdEqyae3pgy9TMmTu3aanE9xhG4SS4ezTTdK0
kN61XprSXS3mCl3Uisx4mEA8jjgcn7Fg0tpMtSao7JHLmbjepQLxCgQpaOwQWdv1
yVwvVQj66T1fzfdytznw6LrfomUN3hnRbes1mdH0m5kQK4/FuLviz4PH8K2aYiT9
ALVeL7mprOHMBrK8/OShAHSXywZb+sIV4bTObaxO9Qz8od8DKAUrJttfXcG6e7OM
CbvKzNXO5rr8ydHMdzv4M1c8o8toAtOHrCHpvm3RtO9IWESo2VuNITs2/mM8ycNE
LQBDkdmVbev1l9K9UhUu17ywZXlHY/C4CDaUeUS9sqHN26sPkLqflMQ/3zu+Xj/g
xp0P8jiq3O1/zcIKBQHDdO9T7bS+oIR/tnMb8APIEHBewILR7Zmtr3WWsYtafnML
4xRQ4YYMbVWUNA+DhNTvtgEinY5ZIWQ3i+rb31eWOMvVtVzVVURlZVvhRjAt8zdp
/wfm+MWBMVzfbwywvfOfXHniav5nYs/V+emtdvGNQolmViqNIJ/eNfv2wxZGCgDc
ckU7i3ItgjfolgnVdDSc5uB4BeIvjWEAI6/d1DlAj5DcxEQZDo4n4XxrErifmjl6
rkRRrP/q+w3/UdWMD7fNTuO7gZBcOuoD4Ajn+vu1UCyePFYM90TLKxBuvV5WVi0I
ZFmGVFJupwJBD+2LcMwM7rZgeNO9nRhIo3n9V8gbafYG35GzZ8EBVSOrJTTwLEva
hGQ1wwrEbyK8F4MdoyeABNu8O3OUgxkBYoh5W196LdixDJIDrg/z4TpxQcVT/bEu
bmPUZdohlxba9znfHtAKFBpSLNMrlI3wYSlk+WkFu8oTRezvg02g8LZauuI42t/l
piv1irPk0RCXqn4d3MT8LqK6mTWKGtuKuQJYqcGwT2ZnEQ90Ajmw4sU5PL6ruZ/u
Th+rQGLUsSrJWVexVRs1Dky4/3ngT87x7DyJM8AjPvG1U9gBX4I6fKkPWSjx/omZ
HFAXkT/bvhSF4PAcPhSci1fbTja4hDJmUjJJA6feBetuDglK3SzrzX0Y+/nnNBlk
TLU02wihVnzrLPL5DdVWttnkj55BWpoDcu2nN7r9jubYtl7En/eHXXzVuroNOFY1
P9QIJ9piMomlCZuYC6J5dc4u74Za4iJbqbHyas9LV6gXX+lWqLnIP7sqIyk7X7S3
dAQBCe+HW+hF1Aq6406WGIU/xCwzUitkmcibOKB4+ASXCql7j1y7ITWIhCy0DWBx
IH1B3Oc9zGGcCGFCgCJoDor40/kWUlmK7jlmWJATwjiib8oi/vauOZDNk57Eyhu/
KHu/TtN47Ll0cDhYLKvxqKm7znoJsAI7hgiH6bUxIwThLnOZfKUXMmIaCBAwmXCM
dRGEUHODlf8GrCqTUfXcihZlqAWY/7X66NgmwsKL9R6RirHoh5tGRiUJooV11sgJ
e9ICJUjSWOhzyZyVtzz8SXH50O2Gi1pnkW9I9KC7Iw6AEcXxOqv6tRzTOsiWfDd9
vAu/23dDj10rAvHT0Vp3ols9IzTlfax32yRywlrZqMjOXUsq1sgY4wnScAT9O5xx
/YPXJf6MKTBo4WTFcA3ukDGi9KfVIlaYlr5ak/dx5p9mQRhj3YZAW7higL4wx5UL
v+x/jyy+bfTgLJDAS9hnVY1jdMrwtKuSKQn9NHcgH0m1eqAmTWUYR/2bI4nNtC9E
4/PJIl/pVO6+e7hhX0NPWDjfg/kmHRlFdPahuXwyezkLTS6RIi2+Xh/HSZMxdEjN
Og5zZMQsB56eagKPIUAEa7/m/ISb+HdhsDHMZ3i9m1z1KezVSlH6KsGk2aPwSrpj
OF3lmFqbwFY6vnq+dmNGS+G/PjgOz1a1hFABeeInNEp3yCJDUnQNQVmW6v7kv5l+
dLl1LqoqJf16Lk0+voWKKiSUn3VRHDT7IGvIb2Q/Y7p6AU/3AxcZpmzuQLuVEx/k
SWlDwltvjADj6918bDnYW7vrRjT/FymORy6Mv72tagqJQUUFC6DBlcPpchfee4Xh
BsBRQyamNrgDHoydBz68TXd13thdlg9Wvg2hOGVIivZrz9XEJpPgXM3/PQKmNfy1
yxrxLZQb4s0f4giyZEVvyuUnvuAN4gVguv8gTQERcMwn80ivLVMV09oFw4b/g0hk
VcoJE/gnJBVJzmYnuIJE6wZhUGPCcRyOiImc0Ni/Dp4ouKmSvumPEpdhBNQaOgNg
3ovZ/d/3n48diB1QTwzRf60WUv+AVzRSZ55INVdGOrkNppbnSYqm4ygLNUIrtHLi
s1mwMQi7YbIMAfVR1Aev9RWWw4q8E++4xGfGQjRtddBFnCf7dmTUx2+dy9XkKFhe
Z8scArBdVrSydna0YJRHEVJ9Y+1EAvaXGKvlr7kiJKicdEZP/bVr4Cl6QlyhL4yY
gPN649rB9NdTECpBBuBXFuLtuU4BHsFQJ+u5Xf0I8ggy6FyWEFo36BvkI6VMu7Dj
H41UZZI5NCcoAXdOmFKw+U6nFMhFQ5hMJq1Bj3cThSkK+suI+TxYjQwBtMXpiBLD
DSdRTLahbJRdl4iBfSEOgp8jhiRUj33/r9AjyjeXQhAukwD2ldBvUp3/Y5WJYfku
6jdT30AIK1iQJRhy/lyd8ZZfyvng37U9QkTeHHhAGQ14asYApeWvqKfN7ONnILa9
5dSmReDFY036OemC6DKPnWfrkhMbgL99J9saySCc1Cc9Jprf/4RhaklmH4idk/oc
VgR9nQJKzTCncx6lrw47k7OQ+8P/HBXkqanBN8b3zhamCu+Oca0nMMIeuYvPJYM5
7IKqIsL+y/vjyHEILoNlBTGU1ETvlv6QsMUF/X3UWexIvy5RvkWSKWRJiGQBUipz
7TLPGtMTAV9ubpVM3dsaxgeNYb4rkNLgh4TywjWDqYcz2EIcpccjQ5MLWQEgoP5n
HXtZU5KCWN2I1sBZPJmNFv7EqycA/HMhrKjKpTYuYK5MnV4UQudXRSHrWW+TlZuu
JL5hfbG2eT6WeGEDSKYBlclhlwS+bEDM7pa+OPaDxEAerrhbTjPieLdMH5XEly0m
KKNSfRS4+0+B7NELM7cQL+jRs0QwTAjP6tIUWSOLdw/PGOD9EQz6mwuoFcVnuSWo
4POd6HecR6zeBLzr6yzF8+FNshdzDTZ62lbFq9zNI/ZCTQ+M5sC1/Q6A/mYUsMQ1
mTJWIdeOxOal0fT15igQJ6E4HgcBoKJM/le8UcdI8kCRdxhRuBA+dYLn5EKBHm07
ZQzmveJBuiAgAy3RWzX6Kshu81LdLDzoVnzBEnqLmhfiUg+NAZc3cCXfQhFubcLm
e0Full4S8V4VeCCKvo/LO5fYLc0ZHHNAz1aTVkWa4hmqMB4P5FUH+pFnCi3S3l4O
3c6Z32oVfTEN/6GZXr4Dv3GrsTfUrPm8r+K10ZPa+wOez9+AR92Vl76gfNwZO1Sv
wMAExBcRdMlvlknT3yh3r5h30SnO33qLESClEF7YVMl7fL076FKx8YPhKb8XiXX8
52dVxShBrI39brHr7QDFwh24LP7I9O0+b2lX6wpljbF5i1fWFPEZL9BGtwiogpAz
jhGMwCQsZ3fCpmb06h1MAEl46yZBM/zRGn7cFG2UljEo8hEg1C1HLoY6FKjwXCL6
WeYUW3HWcKerkJO8z8KWNgoaDUXfVadhbt8OcpBbWOFtIff67r8WvBfDEo6XTaa9
WFXcchpUVIqrUV3ZEI4FCkI6JFz9T0iVOPLQAiliT7UeRDM6Ny1lKCnroxZdz8BS
SQyPDTPJlrk9lQG/+5+zAB2ePpbDR/ABi60kMBv9Yjb94eeBjPuwRNccMQfzqf4h
sxS0S9TaCRuXt9ou0+rrs+pFijNQQp9MsY59ohTWzvmwpduEMG6Oy2DYweN/8Wev
HMW1tLvTOJp1hgdAt88pwNCxv/R3nmXAWA3YSFAU+IllAVIPrDb/EPyPoYc+igEz
OWvaNBBgB6zuCi/xzkAGWcJQ7ZMBtGVIimKlgK4Ks7DjZfLMw2cBOSzdWJfyVcXP
xAmWM4XR14kSbQojqNS9vpXTCBqOP+Dz0EWQIQ3kLymf3dnRXtbOhkvqvSaM6HGa
3WdGKsRjOSRm3Bd+BLjFkK4amF13GeyU4v0lfN55g5Hxiv4QzywVUrHOmqVMEbIN
HcD3HXMB/hqLIke4Uh2zoa7JzHG9oKzfgQ3iJKf4aSzDIxYfOV2Pa7gCQOBeO/kU
937hhrhS7fciAocR0yrEnJwnL7Mz9UTshVv0PC2Ret2iByqSz5neSnE4bsn4QqJe
cDhmpir1mUUDBX//dbEaeNKvBmNsRItA3hp3ZUOJDgeALt664L/Jt6n4LNDOSMHa
eV/SRbAkEQATpdiicG01VkKKDQHEfiXtDapEUzobqel8L2/uQQWBtIL+NFCmevEz
peiYtzVa0JvnNdwdbCUCH3lIq+IxkmuIrKdxCvlYLFXSjL3f9vWy1xeSQabfTd7q
bwOSUnQIYF/jaoCVwl1p33IvBmq86zKU0RSxH1Kavqo8q88tLRntm/qsGXgmeSN4
J4sNPUDFnmdfnNWcgqTCeJmM2x0QK7xzVP1Q7yL368LMU2OyBIicDGwwo/lGcREx
bjbWj+98ue8D5toufPhmYMXi6np/zxn5pD9xbvRRr5VrzqU9hRGosn4TMVChqEBr
rr6Qun0owC/jNFNmVUZaMveZZieDZIs60MXB+INYdBt698ijjm6x1+oEvDlKeOyu
cg47wi4ejW/TPL+bOPWhWq6C/bRWzsyAayrKpOuAGe/OZGTamRyqI+ugLeYrG6aE
Cx2YUdVNpXtdEZNYF4HjELDP967tIqhkrnwNYGP+NhKotqAvRiR5RDn+U7KYiCF7
qyYbUNPmZUW999gzhU8VUDhdGMxRwAZPAHYDm7FqoQFHWWerQLMOWLqdY6h6Ej98
4xguvqoHOENOCtkEdxAVHbo6UbLJqB+hnpu4KQcyL7ymzIX4J8gAmjmdLebp/Pp4
yXZhG5LVEbCvMZ3b99X91xv/2VVyVgFYWBOjW/n0J6ApHPUMfER+oLkNPimWiCCW
tfNg8kU6Ll42RrFiLWINpJAtCVb5uvE09PuYoKiZdJlo9dfoPpa3KYk80sgXaRD8
9l1TjdNo5k/0EgZ7g91ELLSqM2SOC/f3bFTCujVdQwcewjho41wFu7jFk6HfFviE
6A3qJwtPqF0E20ROrdVoElF9Ec3pf0QpcNx//fgjxOmRSFHS9IuRr8arc6oD8pjX
4hmywrhb+CB5Ly/5AzvS1KCmwvNGpOPQWkb1VDUlmWp1ouJqjOvCx5jzqYYbxpa+
qSNQfug2yWupI4utOB07pNDy5zlMxIlq0T8mOxJuzxtDu4shvWp4P7EMKbTiLumJ
4YNXLJofRYlomf3Nfoy41Jb8KaLIpCT8zA/Mqf5x6eVytCxksQPehq9KcJFhqepn
C+tHusrw+Q6fESWMMyVTGdyRxej22c0PL6SU7AoSMW2SGkmcB0SB+Cd9FvYhdtOr
OVgNS12OCAZxrjiXOOxPh0LOR/cBJYRfUbOUgCz9P2uRjqB6cYYY0CGe8U7i38w9
fEtBEmW5+DKLtet++8Y6mlPC8rP6+kzr0EdKArcYfj4WCizd7eaIWywjvCC0NWE9
PCNapgokS6hIEA+gQ42PFMG6mqaOSHC+/ThkGH4VyLz+uzhjSOEhfNlSYnZS2tDu
kMJY/d9LTFfSyV7W9hwhsS2BTd60ZZwWVI3shYm+2TUtbZPZY8drPp+C557nvHzE
5BWuz2dE/PT+pTcf9PEoihmULPEYyHTXHKODd4sKpr8dg6TYHdxwwWLsvKijJsX0
ZmXPFARGcG8upa3OiG+nEABiW1arAkUKtzzjNDtgWjqWY5I0XY1sEcUMRIsYO7vy
4BE2I7GiubxLyODlZ0lW3SIiDUlJaoXLsEZuBb4UulYnSyZz+5I/Mz3asaB3Tt3h
FG8QjG7sb0pTO35NaaM9MpK2U0OR+3+pFXlGE9AK7HRoscZYk6ETmR/9R/eBLdCW
X3UWMQaJCV++bDcNvb1UbM9SFmvQhCqly5Z1VOB8/PF11iuMdiYyfFA32pOeuwsx
IL2QQTxIzT9b36ZNZB0qLVlev0z/nlk3MYMc8nIqp7VHkNwkkXPthEZJw4/4CQY4
ZuSuHGLYyYT/ryOm6d0X4ZxJexrU2eV32alfC2esaMZPmcmGBRbWE44p3JTJKjNF
BM93K9q9MMsHcX9cj4RQ73PVh3KdJuBAjn3IFbLMBvdCSCIT336qHwm3YvrtGixp
RBjjxaKGn7e7wkiVHkSBMuntT758Sar8kPz/wwNGG7dkTIK9JNqFqFGzhFFSi+oz
Mojc0oh7uY4tRqMZyi6sQ6AHkzqyxpy+DZxTIWV7tMaShvbruQxE4eCA2rzrSwdt
CwqaqZGrOFN2VJS51HFvyczH3LCWsQcIlsfpuVLSE3r0LQKtVfvtbDmvRLWtIVim
Y6qBO/JrqbxEnrmlGHy5qsdydcnEOK4CmNXJ1Q2Pa9sR+DNkfwE+t9FdgjdRFZVY
Lmim6LDvHQr6OTdoA8qqwK7FQ9lvK+HxS5kqqlz4i+KAFzXEXjbt5HY2G+BOhZrt
VPcIR1Xwg39wRwEvR7XKKJ3DaWx4tMlF7Gxfg4YTdolFIrvEHyrq91qonK5YVJMv
bL4nTvLwJFLZ74JGL9ht3kjpVYvOMzWmNxLFiOea9gf3Ek2kh9NlBjqL/M3YygfQ
OCiC9avHeQond7g0mq0psD+VqBDgOyKXevKbDUF2uAdOOrfjHBpWn8jeg9mwwUld
hiuPtEwYaFbyODONORebGsOBm4LMHylmFw6mBgxhyMSr9Z0ghsDshBTOFzQzonsx
El+QuQlpryF1mijgmkmEMdRkW+GOUqxejbMsfKDh4/M/DvsCgQzZbYJy4Vga6vFQ
tGWw/glGd/1CUwqwuXqHzO4M1T7r6JTD97bof9tf7cqZGuEi99J2WJrugjg5JFrV
WdKAub17QmSMkUjkjDeK6xhdLiJaygoMP1Jzpg8MIfN2Sh/S95UOq5LUc3uuNva3
be9T3dNSHScmGs/fCwg3EMAIRxTuAS95MDPVcYTsoyAVw7goyWe9wormlahi1jxg
QYtw7WkMbG1ngH+jIORHeOcs1VUco8QL9v725KW1SMxaIaIGUxJJzeFkj4I8lPS0
sa5QzTfvGoFUqrLYbTK0DKrjvxWLibPS9gb2D/d2cLEm8Jp48+5c53MwIuszpOjV
j2IjdH6EmEXU1SuUkNA7Z8GBbzpSEvc5KigyiU3xZKnTGnLFB71nbX/bJL2DlZzu
MkshYzkt7ofjb65nThYTmXp/57HM2psgKO8uobyAQVFHsQNluHxOAPb6tlXupnfL
ZVQQh4gZTrwwDu8SFyMOPP62lomw00bkyEIPfky+afMcYQZ5JvuBfm22OxgqfDJZ
utGgW0Oo32UcJx0pbUxTbg4/9B/xQkL8Ag67/g+L0ZVkMqeIfGf6oOaaSaTDPSsl
urbD97etVVZtfyx/AuhBjjn26u/DiUWP6JrtdwIzqPe0ygiXRKZ6kcqtjy/oAmE2
vPfTk13zL9IBI+WEOBQuAfYvptX2REBvAUj0S54EWIFt7ImybKEzyZiKhgGdo/bv
gFeGb55duk7gzMyfCC5c8aNYGyJtm1gsRf8Ldh9sgEz7/z3ClsLt5ApbERTlsP9K
oJPkeGjwOvZn46Pw1pJRuTmuZ2WY3ZPzgW6X/ezrDVZTrvzbMO7byGX1F0Bu1Vys
9k8xhBAGlM1gJeMi84aSMlMjbkZW1Eiz30a+KZJ9oqjTL3xdaMfxaIycpzfu6ItG
XF5tsziFH8JTrMUAn1fks8remE95VmJDBmftr7ZIBoNihZPwuQ+GP2hLW0GUC6TH
mLj8Ub1ziEXl2MA+xnrefL2iaJq10xUq2ybZKX/OV1SZn8147XOFNuEf3u/zYMNM
5JMmpVdHXvoG4Y2wpWzYaOFPQMqYR25ruN71eec12tJyVcsW+cWYysupo9vs8zfs
vhAV5bA3pcq6Q3T2gnXpRbz5IskDukS1vktcMihdXhMA5oSMHIVVp744243ApxJ4
v2HNCTl60b1tlbfv/SLomEEsEHKBeKqrCE4kv1/C0IN1WMv52d4RbwzQvlLXifj8
ENemtInn16PwBZ/Y91OaLl+BL8W0ToxlbsLp2/HMGsYy54hA2RZN8/cnSd5IMb8+
crUcl3an9HXWittKHXgSh1vFZy3+TuKcwvAJovHAZ4DnqEG74NZhQI3a5nU09WdX
befh5nRekYOA8rj6aLPH0lWsCHfk29vifo4Jmb/cHZcEEiZKwevyY7Z3MiGEoCc4
VV5hMpGshWFRY+ttNDXdHtedhP49DFahNWoUDwvRtyy3BMurkeJOqFB6L45LeNaL
EYvpOLKoKKGLsvTkn3nekKx5evVV11SVIvf3GYmvyzOUEf6REeCt2CAgv5h1/10G
B+CoRZcWpJ2Yhs+w7UIBTgVd8W/I3r5Qty38w5O2NVZHJP0A4oaoNcKMnCAuUklZ
ZPTe1Nc9gRLSrz32EJ1Rvgb8kA/a3tdYWjOWLM/u0hCSGXe4p15qvZ8b4Fny81gr
ACRhxuqPmq03dPMeyhXK0HF0BE+uobVIehvU5qhfqOuQY4GOCnNvrA+p0bGr0QVR
/YQwzmFOA7q6EIu6uLGvj9F3tDu2Pkt5W77d8phvfl961fH101SAjoFADhSlEqeS
Zv45uvo+4A13McUIr4vMvA0xh4XKCXMSk8d92fbXcpmt/ABQAj+8hQj+Dy2rBcsG
0+fn7PlJ6s3oThb+WLdx4/QrR5eRcFQmWMkh46VMTIa+hpw9RUOwfbhQePDrVWV9
DeJ7gR8/tLtjJQmG/sieirgF/zI3oEOEj6skDsedq8arqMIPISNEPvX6Bj5oBywN
s/yAeQmEjW6tzD6Kq5zLf+tE+xa1vHCUpd4gt16LqaayOaw9DcR9IgfhsS7KX1gb
RljLLKA5bWplawUKln7I9CMQBKZQXLDTwdUdNrZrxhW5Y+VQsBYBOSXc7DeFmGEx
Vbmb52RQy3B0I93Jpr1kQJulRWjkpYHv9FU8KnEkgCHaLhl5R53E5yZOqFcPCGel
pJi8HmKvdPvYhzCRg2CPPzUAgySK2lTcd3xTbofvJHG6CUxc0Fgs7c4De/dxa6bj
mZBacpZchKWmDFSAwFbu2Ky9j5FB5ZbyXrweNseR2yafyvCV1wK2IP743iA45JXx
c161xorOe1+Jtf05IqtkrNiWvKSJV0gW75Y+anno8bgIw8fBXuzAHmFNOGpM1iZ0
CAif2IqvnFf3QEknwNRqQzK+Yxx4IPYptCwp5J9NT43/ne4bI26QVl3t/DHaoGsQ
XF1Lt1pCgyWTxYTdd+r7sOdrbrnCW/wP3HhtOMMYQ0IuiyTa/G9FVdifvNc04mC4
z784VvxoXEIYOLYmsgJQ1O+jWhBaTruf1R48L6M5UoOV0yDp7ofQ81MIqPjEz266
19n1BJKoS6q5jCwC7sfxVtPK72A9b4w6BoM61Ecc6301pISgWWguZeFyysCCIZdN
pSo68N78Nt3nK1c3WsAxF+8HYkjuI5epOEha8vSes1ZyCzEVqmO6wndGtv0h1y8L
9LzaDb9Kv3JDhjAwk7M5RB9pKTF76inD9GK0C5jQUX44/ojVwlrF8fY5fmOJ7gf2
sVtPMHGTFtjovPZeIc8PjcLCkLUIqHslML7lrJ0OLxhJmSd3voEc3Ozu4wkdGWeQ
c6kbqNT88+mHu5e/erZ+DQ9+Gv52N6vMyNtRfbBVrmDPCLUnuLX83CHzIVjSj2SV
a9aQJ+GUl/Qnmg4VrV3KfvNmNQAPTo1dFYYDBcUNuHWBNlm8WMoPBXVUYk2vIg78
XbuUeVyyglss7+E1yTdpjxINKod3kU9zBlaKwARQFUNHwv3Hrhqe3PUsZJY23Xhd
9cTMYhlnpPJz0AhINCF9LmGWFgC8AHoRwQ4woHvpe5RAebvdgLoAld3NSw5Ca0vL
c6CZ3HOAE1srE38ItJMfS827piqTuAwjWb6tsbFyIjNscXEJTXQsVSQXtQt2nPER
hlEcg9WC1KYM6s7CrDvnp6Rr78Va1Qo1/9tKZ2pyJeHfrMechX/n9A+O1R0jW+NI
GnE2ZGvvZe0wGKjvRJYJIBV4kYmo+R+nPZBQYUoEvxir9B4Y00JFiuPcjmcJ8SBs
Pd54SfAupaIqClgM4jBSYJ5EvDh3m3ec3ugXXrzLNWnX5bXLFnlbY47Us39pGKgE
Oja23Y/f3+6s7DQ/qi/PHHkjC02QpWSsZT74ZWMb3sVr6fTACsdyAZdDSxNSN2vg
snb3Ovtxy8tEKlKtITVDleJSRom5OxB83804gAf9b4kh2tBmlEoJexYAtRK19UNU
xvZUzgqCwSbwgdPy76MVc1YUoXQmnntKHzYy/f7Wk3k8iBTM97nn/qqzylB5okCa
DZoPRcqvA13JUoE9RzBmvlvLT5aCRorISwPcuf71IFGAFdjBuz2ybR7vTxpt2Tum
jW2YvMdvcxK/hpzSJs5b54NHEQZ4n1p17Y7WIWhtgho367PrQCKmukL+uRvRvV6i
cGjRFrnzdyojastHy3eaSobCOHBx0FAKD6KdNeuICAZMbUL7BRUEvwAPC//irnK+
hQwJqWaIcb56KEphUkN6DD+8Y9x1N2VIAnRcoMmaKQjsVgx4Lb7PCe3S7/A+54Ka
EQ2q1tUzeKvdOCy2mdcUHkt68WjjkSptk6qZ106m6b99o95OpZ6ea3aTWfBmtuvU
2Dt4lawRvKTzIYKdigS20jLOIgHi40Ku+kvhhE7onBs5yjymKogvdRQTNHbfrlLS
bErdioOZcYxq5mEPyDtGdSOFyeJX+mVFmDY/zT66VcOxzJTKPYvKdBE6jeIpoN5E
MDMEI9XQf4EfOiXuIwgU2K9YNjYAQ/nrgUqddWzNzFDDTsQ/NIilWcp+7X15rvo+
W4BPMMf9/0QxkwPLBLgnL4S7pmtCRt9SqXEJngAqWZ4tOrePVAMF8XVuIXsuH1FA
8+GyzEoCiIfqtLCuNF3yANgY0ZqYk/6lPDX84qu1xb88/17omXXzzGFndK60D0OK
XeuyPXeGK3CetkJdZNYopCEHQlstBQ8l8i+VNiHbhkwn5CXHDhXUrvducz2qWjVL
QT5LvY+7PgYoIx+ZWvwAAkFbYe2NJNfg54Gi6H8YFskRRj+13IQ5sgjQBVrqdu27
oGvAcDeT8xC+2kWrnfa0gKtnVIve9mHSOYcyo6kcW0c1d611pFVqyJC+1cCO2T1D
iGMUn9AsWMI3qLtVf7nHpmTvqCTPvVBMUzC+TL/oS2DpBRLj5XajpjonxRyCFlaf
hrU4LBgG4EF44AKyqtS/epJyKDwfcA7qlyVLNIWJaS0DvxhktRf4AVghntRtq8tO
ULTLPfRLhtTMX0xvc3Rjtmxk/x7DUbk003YBaWZy+lRJOZNPUXIh4H0iMObZrrA9
+zL6G128fjrJV7SuVsipux9UgBVr4Kb98QdXrAHGIUZe+y5adbg0Rb7TBOX4Gd34
5jr8AEE2k7EVR5OrnkhDb6DCAw8aS7Hb9tJNaZotgxsWSYaUZ16NuxDcmX2O11gH
hlFSkVBEeXSMvw0oPYSCpt3wJT0RQy/dGYrMNWmsUB4jxaBB/9T++diYfQG0vG0W
ZJ4zgo0HafZ5HJpmQ8e8ok08zzDkeYK0ph4yuR6SrwfR6C9EpyhjQMexEqGXqL/u
km09JTbn0hhSKvDXtncOKVaa3kUj2/cbX4zmgKgHltawQ10/YGUQOmJSqmIZ5jvK
9dbQghglePtQ8AdOjQZvJCXpvkggavdxS9yOg2FoWu+9yq4bHgylCaR0ryYkMWcD
GudyKOTUJfvNJ7U8A5kKDHVrl6wt7fflg9dB0owPJJzjPYvsZ4j6UnzLsui6rTVx
EaFN0SjMG4Pad4PMjS7uK4patvgpZNwz3p7GSjod+++3phqSgDR6hyYRloO6Wwl3
NHXM/WQfMYK9pJm+N7N6LHkeQEPv2vdG5nqaMrhrYMW4ZRqLpjktRD1D5clmaiso
7FshraepMgAnbNKqC8kpHGcZVx7niccvnOKIW9JZSBom0YlxawbhMWaI9zlEdOvM
pGQw8mcEt3Mk+TXtbVdFrYxZ4wUwhQxqmdSn2AINxlLAgTJsp3WvijmNwPVZjH8j
7nCTOG7U3nmXznjzg/Gk4vT9sdX5np40XIvs8sNn5QHJsqMnoEXKwJA+8js2fbw0
YUFAWd1iWLQVdscj4AqAnbk+TYQTaonN7PFpxbnSx+4F/eON3Z8uoqZAt6s2bT2W
Ei8EAxeRtqeMUnWZeoDZ+3DFSLR4jib+dIuRGVkOlt6VDDxiQji7THSkqUavUc02
x0yPTm2pKN5WMbcTUz3m3oE4EF7aU3hHyupVRc3zAOgGA6CF0mXDYZFM1610sf1S
dkNisvOwnRtMwk2q4sJvSbhQ+SB5R3I2UjKfWMJYUkMo5nImGSx6c2r8FpvNA1Ss
2hXjRUoTIedozH24OwlIHR4jrFOm1ppPnVnZmm6YxULw/mNt1ZbEE2ul0UzaOW+M
nz/kzTj1QrK4vYBioxTDKqGVutwdKzRBPw8X+fdCA7AQxna9511ZtKs6LTXPGmIw
MXSUxMV4aMxsWcOV8mH2UccoU0R09vgqunoQu/W0Nk0zO/OoU7VKIiQc2NJl8nj5
6BdaREPm16WfwHLFQwiUpBa/l2fqLcisqQzyhsPjJ8oAJFrRKl7YhfrBGSTtwd5j
KaxnouHg1vZgqjq2k0gJffzUAFT0XOuTY/Sxv/P64kxj8FdeYfD5SoNBBbWgYzIv
cs2BjlsnIUGNNxDJrOwiwHz4mhB8fce6s5lTqzdi3nLNRhQW96R59I60Wjmk+vLL
yLbc2ZjnR6EOiTFxfqDuucsuAJ7unK4NMEaDmU81t/Eap4MQw7l1mo16hZrryUY1
5a9ZjSvvG2sRuIitSYawNmYaZMjS9DswjFmwPYMPQjVE2lX6gXs3pQY7Cq9jFj8C
TTy53Jc95jkAcZhJtveQW+xPHejWNUE7oCbyUmohrromNGJLYO/00Sc9hiJmEzxe
cYEC5P8tZ1hA1b0ZFWBza7MVeYo895XtnzkUvO6SlnZzlc9bYnk/vKgT7p7yw+xD
p1a2TC3ZJcV+zfeg6eM5k5P2HQFT8v705TT7PFjdbQ66WpoPJm4xqSoy7Oeisey9
3V94WR78bjsxoOxjqEtP9DgoEPdV8+m5QnttnFSw04diA73meQoRKxYfwfFj1HME
AEjnmZOs+fxQ2e1hTsJtunjOJJKCGRBwHkrH99iJEMRJta88SeV6/5MamjKPRsQb
Lk88W8fVNhWzJ8+i7rMC0P/EH23lInzZCYc0rntCHcfG5AFiq0Zkttm1KWFgoT73
F2yUdxJ5NJi0gBR92mBODLMidspelypg7UUeeVK1T7eYcAFTEalG6Y07fUkpe833
6VexQ/dbIv67jByUmYY+VlUriCLaWZTLEZ8qzQxyuec2JCx7S/Sz8w0gb1lxNHpF
zKorsQxKAo25TcALv8eMk/+kQMorf0zC2U/K5D9ZuSmtYNd461lMD/oF1O7G3GrY
JujfN6IpYJR/6+f95B4nX86uogTnoGimCNeKRVsHeEpuXDwd+VStIOsmgVA4K4sP
gjev7Yr/nWx73gMyxwTMp791MIjHS3bAAPDnvu+VjY5lwIiHxLIYj3jDe2Xbfnuy
sNDgElOtwZMaOEOPPvoEYEeL3eFH8KqKYtatial81YhAIc9F6FamqTV7Pk2jHE9R
CV5KLQbaYb7jpEgaZ41+XxFoood+O7qWq4kyzxsEaIucsuF9Ds0A5fQkVckTMZPW
pkj581lJ/uFKyhIQvOKON5CUPyMRhlMqU9oqrIvGpABYMhGdPpZmfsE99FctrJr8
cW8gb/UoEHen623iUi8Zl4+EhxjwdQWaypO5kRwrTKnk5U8oYwyCwD3ioMLfDjLd
EqffPDaf1tI/RMH7Yn6jP6o1vbK0zJVt0N5yRJRgmC2Z8PFmwDOwrpIPn0KT7DPC
CZP1yuqHEjMmLrqZLsnfdsSMAq/vlLMl0O93x8PmAEzY7jvNQlZWbhh8We78CNRf
JTy523Kww+rNkJDcHTgezSyiFT6WNkKKTW1JBupWM9Ws5xfWJi03skXNi8gr3+hs
uhb0eN8UctFY1jso73SF9qy2vRwZy6psRc8h6ktCYb/b3WIwhnKxe/rFrE1Vk9B8
cV1pAFyOcbRRVO+uCuBFhcxqNV2+wHegSATL9S92O+aOySiTdWj3Bax7cDPw7hnt
KUWDI0WKaSpWwupHLx8KaEWNDLmHMYMx3MwMZulMaBsbwzKpIknNn/l3IbOiWTih
9tfvePM+6sFgI7RTNQhHtpC3Gp/B2lnWZ7/h9oflMc1xdptNUU1z0Fyvi4QtDpTJ
R91Ex799QmJi34ICoCO2+jYNiKRheUA6IpxbLJjWOxVa7ZiWty0jeSqou1wj4Kr4
0+ZZWf9MeElM/ZdctyqOMC8Pj9pIodLgMGbMw1pM/a02O337ctrtO35uHekR2SG1
Aeulq7N5cP+Fsiks92az2FAHiQOhdkKZsk//6gV7Rc8kjwp26fJ73ZIGL1UCJobA
e+psBvhGdrgHOzQh6+cI0bs55AWgPrM01BwaMIpuQI0VKDtGx501pypj//U3PRYY
g/RuK7B3WqwvQwdYdVjF4lWZ7elGmBHGZcBdJwK9d7dQ00huOvjAN5Dvke/hJmYw
Yox1F8JVPzr85COm+/1Utj20ixtowKlhZUxyS4UXK/kVJN0rg35NzpaJwC7j5VFx
BGumMABNrERRK6RK+Ks6Sf08iaBi9FMlUTL2ldM9pf2F2q2Ne3ukBxdiyq3r27LF
NvFZUdenl85YpsZ//D6xKdsxJbbkb+4Y8toDXAHrSV0k1BOPxbmQmPrFbS/bEy4b
T4UKchGISWv5EsVsbYvBMHAqFrLI2/I1JYMNktlr4cOCmBDDC/5j9LdRtT40SF2g
UGC29I+wOkgbXQaFTa+FdHTIH7l2ER86pt1OfVWTdHAbyDFlfziQcyMsI1Wb7Num
s94vvnemmNSlELKyq1r4SyygZuK4rcwoJxNS98rTtvEu2gBTKziJhl0mdgKMr3m2
/8yBZkHu53rLfmiXUL+savsDBIty/NJRtBtPLB/i0TuOaxVAjMRO1qbA35i5pGl9
ZbDL9uyVf1yrT3QRchjAmMtUQFx8xEwHwBDk/AI/OCWwjGcfO/qpEqAVZCVTL/xX
IS5RksGOMPiMIOI9yrADNx9/Zhz8+SoffHkcpwZKOEtGgjDNoHc0ygE+9ESD6XRw
2pwIy89IeFK+Ga8CxE4GEZ5ZzCi5UklDYWY+b6i9Zp3c3DZ0i2qD7z6RMasyG/v9
2mm1YMzZppoeiWUn5p3NdLsXpThlbECJuysROBJ0x2+JHeomIvoqV81efNCFoY2R
6ZA3k+Ch9uwSqHRhme559iWTGezvhVbMo1qcGWoQpc3iuah1YNhTj5BT+JqAWVHp
g+a0/0FMdXyFf9Bxdh7O2mFGvoWEqTWt71zKz/UZAJ0unPwZDK1xiaHUFMkHBrKS
LDbW+dgDm7jx+CRyuJZbsagZ2PSaCrSJlv9Dc6vKXthyuAl5O6vifOi2aAv+1Fiy
TcnFe/eb8CjPwAds/WI9bkEu/2jOU4iQp7o5XthpCwJycwUiN7gIj+Mf4Kn30k8Q
153S2eio888bLhlZANwAozNulTOlwnGnanC0Qyws0ILlwNN7zIgnZotgSOJVDDqZ
rx55I6sSBbxhbl2d0T18bIgmMAEHhSdFKx95Su089YGn5McGucUROEQhEtyIRneL
1thfuPiEiLzWGyenEB5uKhMRNsTYO73SqgRCSr7h1PTHU4eDikhGSt+gG9226XYm
jzMtqPZ5pVRhySH3D5/Q9DoGS5jQINGULlAWFH2VSme9dRoab2vksK0NCFEa3liF
6J+VHxKOf9NmrZS+rLl76wOZwu1i3Akt4HkCyj5QMEqaILkjvR8GzdD5yOoNp2TI
lo5But8DmYBUu7QxGNdDEQea6z3hVyEItj2RULaP11MuqnT/1fO0CU3EBPAM+vga
rr1BhwOVvMGc6Lsd0il77wFxDEh10XpoxXVN8gID60whlzc5ClLEj2AKZzm52H86
UVyOxA4ebVWSdNegD6G94scjPPUxpro9M+DMJZKpTpO6Uz9SC7qBp5ycjsYCabsR
xHAsxbVUbfDcmlRg9lgVX0Rws7VGhbwYTIM6l+Ska7tSlcTOFBkorKL27WcnVIUE
eN9oDnOMa+OOjCO1Hxap4saioXJW/YMNCp7K5olTBzfTfJ3hWxt9Xgh7px0SPkWe
vW2Obor/GX6Hx8OpHaWqehRN6Ctkfw1+EEpJZHfrNIwQpXtDWv7eVGYCB0IO80RB
UXa5hrFdTc+KD5x/fEnFa8jUD/uNmqJ6kVhW45g34KC9cd3/YTS8Lor1QqkDoaT6
H19p3armXs8OFIy1x9tzFfNiI9SSrQIQk6rsz15dC0SC6XSsyrKRylooNbrjLIfI
d/CXi3V6r8buhAG6BwmZuIJakkJhNgbpR7F7hwlri1zBqh8KDYmQRaMOdSc1apLh
oXwMLIXIISuhXC9eaEwVxcgzruOKmL/DYJ51m1bGtM3JvK6vRvQmI+Ir/KpdoHeU
0j6i9XyAT2qkMtCfsK+7YMC814Xv7nAxfpwmRjcZXuKYznq5cvemuphkwL1FLvCu
UgQwRw78J5tv9T3owSQNGGSmWR3FqlWOEt5H+tTVagPcSznAJLoT+ejuan6T2Cg9
mVzAB4/0Wn2fu7z+i+/ip378kjb19/wm5J2Ftcnwb3ph1vig+iBtu4BfNmZednRs
jexlvXoIKhm/3vdRqhiz7NsFkQbv2P6lIdY/kSH/4+TEEKknFmhKk8idX2rGxaOI
VzxsgJcmayBO4zFqVGvIiYaPYK73tBECHb6L9TrUN4/i3JbGKnZhHxhJBXofI8cL
r98RdNMtMJFJVVhCBbprMuD5X9cwV6S44St/M7Zzb10SfMLITO2WCjOMR8uV8v2J
a/5TQJoyoN2CzNPjqxg2cijz/LhH4JuOGMEqZuS7tR8rOYLEUgeyRKz7X04LV6Fr
xeASZyipVa4p1d7Brh+ApP06Q74PMx7VTjcUGvj1tylVMzcQ2VgOTTvW68C/RuGc
IPI/dql2lpkVpqtdKeSOwXmm2nBO5Yboq5t4XSIiehDWiZlknBLNrXdI7jEwy8RJ
4l3UwbNziG2SJIwC0UnfhIltECcHcouUck1E5r+R01wpP3HA4PaLHr+ODQ36Tod3
b6v4DTLC5dZD+WjvpNTU/HvdGkDg4qx6p/zEgosl/i98Ns4+aE2Dc/Vmga7mzCVM
fjH1j9JywqaK57WA1ORwbujwREygu9ugQX66D6/FR3DTZh/7yQGIklbB8ph7MKQa
jDhqIUy8fTdka2WUQlb4U4x0GdRcZuBjBqwZAz5ChvuaEqb7fBiX8oot+57rWJ4y
LZ493TWS7Bk9El6kmnMvsDvRtpuLEGpitdIVWK07Oj7nhXnIaoJaX5wpGKg8Xjzs
8jBz2BBT6hNUFfWvQDzwFY5T2KwoQEn1MXW6N5bCoSm/lsbTxtLv4sfKPzvCL2zr
rfLeIo8zaY0Iki+zp2+VSRuZETxYyOSmFzRlvtuxchCtRMdJfrLOWyZTx9Lm6J04
LKD/Dsm9iopHcMwWdixNhXM8C3BFHhFjyngoZph3vtI6LEHsvR3WCn0InxS6pJYA
/kxKosisnF0fl7ZINy0Yd5MA6ylQOblTfmL38Q8Tqg+aB70FZtnszTszrAJgdtOd
fB1HP/Wjt0OL+rCDHyx9kRAgesX+F17QmJWEWQp3IkV2PnNmBApAj7DjFzSijVg9
yc4w6FjbSf0PzUIG0y2eX4jOqtFikr45nKhIF0u6cTE7uzf9r0vRqNu19qf1nbnp
LPHG1h2AIVo6m3puZHTkXv4lN9h3Q3Yuv+IMpF+1xtcXUcFz+pvaCLSqQBXuaP7N
AdrqAviw6g+3X7GvHHw3sfPb2qtsA4c5xSyRmKKyvvKdGN8vA5NTLs7b+MggJDq3
XIo3Of3pdv4mSy/nnBPvhGXLJHelrZQGwmN24X7DJMzqvh/30hKWE25cAeRidkVp
qLmkuPQeD5WHrTzCUlhxk1wz6q51w4lR/fC3kPt/4ha7wLCMGIzT7CM6tnk/RJjS
nKa0ovuexSPFdzykqMFCK2g512I/ovwOwQk8GKXJhlGg9FgOEY2hsyYhQeQFtSyR
FQ7X/2R6/xnnhJZ6g+1veL+F/mMR317Oh8UjCNVSPYY6fyt0qwF9f+kfvvwdf4ah
aE7azZkSC5ZFXo4l3WhunHV2un0ksmdsThvQUXxz43kLLQ4yQN07BNgUPiOycqc4
G6+hbJ3tXNyw9FcAMePFmDEjUBLMqcZETgcWk0PUu1swgc8W4v0b9XT9c4l+0EYT
IbcXxL1o+XXCHLdwMSrQsFnhARcdRkAAaS65hl7kiXiRfBD6OD1QSmwnVk+Lb0iF
74U7jgT/u4Y550mvgtfq307fCI5PCpVkPU9TGu8bCNdrdOtxAx9VYe01PqDmLJ9b
v5gLdJNTVeTNwJSLhRs3xEmPyobfmiqrPUzrznDE1jM9oy32QCivX+haYqQeTHTJ
ciFFmZXj1gSeyhL02gpUtBQlCqLCUnY8y3JYdBuwz2gJBTk2GdpCySF9t1EM4e+j
aRcEjEoeJJupQI2uTf75u7jZ6540kHHxvFFyWGIt1HkhJgH/2AB7vK1PZ5Oqyaxl
a31YqWhD5xwcVgw6Av5uvwLaLG6aAqWP2Jkp0hDi8JtFkV1CS/TNJH9RaJPRHXPM
vpH5VoPZ0Vtkp7oQmX+ir9mUm3c8cbzT+c3/ShgTdBkfHxDzOthbswYqfDvM5FPv
6mOZghghL+y1ziD+2Ivy75IaUjBtFKNWq2bXkisnQMb/aWnzmu0X0N4thwiRT0uO
Hm2vM2+3E+Svy38U5yEyn97lmVGIljT6aZhPzkuCzs4vDKVmVfCxZHYcn/gZAR3o
6TfjoLlnJ0llqLJKZqnCKK5lnUF3ZjcePfqx36qcjObXT7Nbh1kcMoRe9FC6hRgG
W/i06PkoMSxHGR2Pbtd0B+Do6MmmSsauzIgC0omjNdgUOJnftqsam10HTEWuANEi
HXZVnhGX5uTmRGBh8nk5PIMP+HVFlKqnQ2uBEQcmO9MAIdiX0xYVRWaNqW6i3LZU
fFgUANdaSx9BFB5vN5tkoRdq1jTo0qKk3tpr9EkB2TE73nO+TdyvA9u+PEfNlnA4
4wwDolIk7luvowIs6PDdt7ygVoDjR3Q46n7uCx5c8tfzhRFnC87XW0eEfElUNCxp
ysbssxLCp9DsxOjXovsn5gsMe7B1Tew3/eeXhc4oEEtkKvhKmolng7eciH/SIUdN
Sop9siR/R1HZpzAQ+ma3hURJQJBcEKHTYmo/CffmgNoOoy7fK0Dy3F/p+/ajTDHQ
S+yReHeqinME1IdjAXe6/qw2j2tOv5T+Qr1JSxPI2kfJb/2q7YX5r+DHvwPH2LU1
Z94DtZ6kt93QMHDnN7jIiXWpyI9Fhbc8nCGQVnAfzuS/SZeNF3JKgvTV8+K+GuFu
YRSyvgAloIAHnnoIacH+xpT5ZnG7SbPUT/cEmM4BWzVpFuoLF5AsAnaCKhjSPOIu
RBssyQNX5mvxOShsM57u3YCUJH3VsiLvwbTsPfHdiAC5IEpAOT0CtTzmgTD7Qv+y
I++xPwN6O8gfaqRzwUsv7lz/ouirGRzsWbvJT2p7VsHGmTSYUm0VlvkZe5sv2FhU
TM7RudZxUYbxRuV0mb3jA5JYvxKOnjy3aZVN29kp9gptcehWaKSbopaSDYkWgtQi
slzqdtyzh8NWL0LUwG2Zpa6kFNDyqkx11NPzHrbS1xkfR26V639FtDjToE0Vgfbo
Ub5GmZ1i65WxARUCi+oHVUWslNEQHeyvBLsWPmc1eEWmgJC9KBwCWLReX2zZEpFm
kJPwOUTwvZF6A6DjVjHYVIj1ClbXzvIP+qH6Qea+ezh9Hm/JM/uhVDW8I/hiWwXp
WQA9S9In3tAo2vjOeDMOc/xfu186xfq0+NbJXR44waXt8eMZs4eO7uQMaxZ9A3/t
v3zMNQiFWsF7usmUEBEDbwuHYT9yjI6bNtYcHMDv/vZxCBbTYiCuls3S+3wbBoyr
eOtzrBa9PU4oUywF2vy+Z+zpTLf1VWp3SPZm1Wyd2wdhn7XeV+MCulwway2pw6hZ
cq3qgqda1wow8ld8gspNNjzgkOARXRt+UOjuFH2fU38/Zsi5o+KvwMktJvQ6jfD3
v35tk9YWvYo2Wr6WkNPr5G7TeIrxKE0boGHiNyTH6DnADHdh0J/pMJIQGEE1c4Wr
GaQ/b/fusdGrtnpq89Y2COzINvlGSR4MJjkQOHwWOZaQK25VDO1yp5W9GlXDc/5s
t8ejim1nXXVx/jdPxouNUqTE2uYbPz63wQQQv1MFUIlwVAp7K74u9GUY6boNgvEC
/gNgneWDyR5A9h08WTt2/s3JEKneFd7erIskKt9zEJ5yQOsonOBMzNppgXHAYBpa
UBl46PABSRh8fgzefTTH01p4bM2WB2ho4JF+kv0/eNSkRU19pxtgOroTvV+d5LZS
VlWOYZBuaxPbdCCiX26lTA8vMUgIJ/R/mQD4fMjwXHqQqQrE/tq3L6ifxI7U71+U
8vVCdqED5JzW00BiyJ4BpEGLnLHt6uMgokGhsNw3vTPLg3T2vJCmE49mgugluACP
wSB6vU38OA3UmOWAfADyFC3MHF4oUxKPkDKzXu/JqxcA5neK+5CvSfge2s3xMehJ
HMQY2q+xK+LfS924bTMgK5avV0aKCqkx4ZkqkM18+tLkKh2ieGLGRjrIZmSisN+n
jvJBZXWp3indbKgEehi7UbThpuWoDovPF570otDo1hizCS/MBt7G2qQ/9XBHT445
633gfc5LHssrQRTTXUuCM0BahOU88YngQ5ZbZVgfeHk/TXv1PR00LSXG/913U6MU
x5muWqGX82eCCR234+zqZCJ1wh9PY2hnnyC3rgK+iE1tluVYo+aHwMzh209onBv0
R9y5IW2W3+pYlFAqAu47Se1Fk5OgnAA616pHX/deTUwzFK3/K0Y7ZaKcVnz8/FVg
0Pg8uzswLNndp6r7vbqWPKntCJmgJrfd/zkmS9AnlyN09vt3YDfTFwHWSzk+VhaX
QjTXqBs1HM/ZF2ldkFBIcYSCGDblrmge1hoOYVR8wulnTGCoF1/wV0d9MMjgAhaG
Npev3+J+zkGuMKyXAVFATVTpQebizq7Hj2wKZeNWvoAtiWrc6iDL5Zt28osFSChk
HICNp+IFIK+jebTj4loMStkMCzX7fpCSImV1sxwzr7chCz1GRlYq5wAxxnNYEtgH
V4bzVD/7ZqxQxOL3YVCQ+nsMyKsz9yaZKbQQHh51HLIuY5J5vKKgtMbGN35ilLJP
u+lAB1UjcOQiYdde4hUxl+bnOpfIzmnVZH0Bv8pkt7YI9dayI31+kJSXh5jsViB+
9pE3Rm8mdKSytXVGEdJ1WN8oD1YXRo4D0myOG9Uj+PhfidoCch6u7turtn5aWvRK
mybIuBZY24u8MzQdgN+CoRcD7odaWbC7QzQoOD3kjy+EccalPi5nbSF6ShFvnZmD
PosBdORH45E88WnCDd5GD7u9xZPPi1OQnoG0p3ZEJuxHcK8aB6N5zMtbZtJECbZ8
Kgap7eAK86okz76sRMXoxNojgX2rqnrjuD5VQoPqPAVqIHmo2Wmyp/kIndAkf0zJ
89vrkiAgkwmqHKuaV+Ci+lk236wU35T89NcZAK6TH3E96DKaIqLgQJwfJR8O+gkg
UVWCiUnQfgr0Z/xrXCC+9sa+SqoEkf5rAMQwOgDf82kKuF5V7FA3K7aG61Jiwyzr
dF+YYgLviJdxnlXp182U+Cjjj/HKqTa9TIcpOuQFxsOUL7haKoY01YC0cNjEUALO
zdZQxWurp/PlfVyejApJyD8rextuuo32LM0lVBAUvEeKEDiNU/UfE/mOjixB9ozb
H5Slkhqd3kYHsbbDtzYr0Ue1qIhM6gNtRVASP0ZJqEPWMrmSQglNXrMhLk4MaxeC
KxKurNXD+fqqt/ggDjNCOP/NzX68PDklVdEQWOBiK/LsVjJhRdX8QqFDTWnqn3si
Dz0cpM/0ll0EY6mkVHpmdujaexYyNWTi1AbGxdbS/2mTJ/K1H2szmZNK8Cs29JPx
lli0DF0nFM2qSZ7m8bJP/JCQacgOemZFKxvpmhHQVB9SrDpbBfqyzQXu5C6cn6dX
BrrOmj64CpZCAH75nYl1gKIi+yocWxjvov/XOZj+frq8LaUYpWHg/gzVUCqoT9fI
Br/vNoMbMWdwQX6T5rpxL6qSCM+PPoqsdD+MW8LqTAZqF0hXbhvASs4MDoDKh8E5
Gip9GGs/DzsebsTBjk44UnA2SYFtgANm0iZ5qPeatVpcy/nG3s9bK493TxqV0m6d
WbbE24YxmsWCKCUR+a4EbO4N/DBssZppubbV2FcCYn3kxKiPUUlZCXGT+WHGuUba
LsCVhNvz/FycrJnNY5MFGQvQlHsirdUC4mK6WtOn7/kWcxaGEGdRASPJpAMnUHUz
A5GAb/fGev72agKIkrpcSWYxI+aPf1dEdy0Cd2u7FSQbyR4lh9PWOxh2MwHDuvFB
SUAZaadnilHPC8DqCQmbCfgEaezjq2846vHOz2WyujPxKZQfZU6x3vlMvpryWYkd
355cVnmKaDybtV+Zt2lRI2K9O2RQ1JjZgQYhFBeJP13YGEQ8X7m5T2rH8OBfepfS
soA/noKtQMFRYGYccYcQj5OfS8mbANqS5sAeuamTVwFZBukT8VxJSlvJcbg0Si98
S02c9orBYapPnOGMRw25d5AAAd8PBgYxgjcmrWkRjDM1GvxvtaRh77SR8fkwZwP4
i3Rxtg/akXo4uiWbnXF+o+lV9S9M8Xx0XimdANLHN6RGzUY2N58gFiF+IxhZ/7pm
OsowbDLqVm1++Doz7PZ6oJSNswtqC4ca9ohy/1RZbzTUuDxEX2lIEopPe7YtfKVr
lWcwhfbDJX0XaV7hVEXwjN6LYBVO4Oi50QP4GPdSsbCWrgC7tkcTIpnUJUSaw9j7
toC+X7emfrkCOAhGUoR7UhUBk3mW9ntPULy7UWVhEqn8k7xgFcoAhQi3hW4S+RLA
axEUJtEiubXK2oK1/0OYRNUyyp+U96xxX3UIY1JhZgpUENqL4qeNXqB/mnArIhib
e3qd87aVfSziEXnaUuaYpzIZhnk9Gnf2/odIrXmOGd/CDPMu9klewvVDccOGKylE
yO/Uajh0Svq9IixrTd97zz83uT4odAedkwl3dvcGER2GKVAhUo3LuAgPt+FDGqqE
K2ybstx7Z0A8xZsNuCsaS0A0i9F2D9NDUcv+TO4bolbTbBBIeOGmikFW/5TPAAF7
rFl9mAygKm4YeKSR3q5lbeDXWD4X4AUKb+HYFrQvfGp8Gu2HfaSAuzihUYFTSeRG
k6AgM6Rqim4iJ2kUhvkxhVABL6bxKQDWC3BzGmGFuqEEcBSbksD3PjgVuOkpMq2M
Kb6RIzBdmoew4t65EXYrVdUHJ+f+BNb8RDx1yrl+U0JqyPkCKufeK66jHrwmCcPQ
pOAGmcQa1DlaCiKxxEaj9CTxpamcqEHxYnezBaOg7jBu8gdxDWvOfj8c6I+mxwFj
gOGHB4LhzbAlzPb6vj+bU1U2erAuXqKveEYDZFn4FsAFNVyNqAP50bS70t1QjCto
hwUCvlK+6ZPF2K0DqX93c6U2IzjE9Gl9rIbxKMDUYKRxKflbMrWUmT3kuKv4Hx+9
Z12XCdQwqh82sa5Uw2A405FUrd0gSo3NDQ0WYGZS3gi5/cNu3LqfB9cyU66PjCWa
BDhqel3ScIjnfVfkQCva2J6juXeCLQlIQxEOm9SQCe70Efjucml4oA7xj0uPNCbk
zC20dWHRy7EkwBl5mQOosiWFS/VrROF6x0qVrnhhNNJxY5vEACwHqZc1zo7V9pII
tjxjiymziLwyChfFC2pUf+jW0KUKBCix7wY4TPmd9uQU6E8GuRDBfrnYwmwWYEMG
bMd1MgNHXz20J1qhofh+GUB2BmldI1JmNnyzzocX5pd+AIFW7wAYSMpDzRKmAMuP
OxUCzUp3JD5f84H8ROVrd3ZiGu78Wd2m9PQ/TB9zCqZ5OIhQqQ9geqKTE1y7lvU0
rpLnI2RaH2pDXyPwmHpyaWcH9BF6kg/SVcXPFBZUysr9g4SLSF7QlzzIvbG992mq
xeN6fO4keD5+v5aSEeLZS7DeT5CCGp8KOUVHHXayYTV0wDYEImd4d1PVz7pQik4w
/77fSXtHUSBVyE/Vtdod8z8VQ7PwDyqxe+mibQrM7Cri7OkLOCwRmI5pmjegUeS8
BA3ISqftDtras7jrK9KRsQ0UagzxoEpBi4Bsucp1lhN0MpoSyw2J0+abgLWjwGPk
/02ZFtXj9/OfyAbkWm9EdrSb37QNfQLDHf0bV6xb6F4NTKTxXeMyWcYGAX3NYphq
i/h11wnPXOUz0CXnaLUwuPtSK1NZ7Uq96J1Cuqxf0ZqW79OINTD3FliQYT2+6kmG
K1VFhS0RamQq/pTHRz1Ld+sf/eCeuuZfRVLT9EQompfRZDhZgqmldN6RugyF+OZc
cIJ0QlgZClgRler2WZCqPETUmH1TaqwkzIumz8R/DCI574v8q7bvhqKpN+uQa08M
d+bo+wNnVM+vyR1p9Kt+Nu4ojxLqSAv8P2hMSgYFLrlt3kEu233XnbSdFbjxx7Di
W7bnheW1BEEooIK1YAh6YZs3j4B3O6/y9dNp54Pg/O1RjhKMW6cEDKVOl0++RbfM
tylR1tdwHRCnRemKzY9F4kLoCftieKT0Nx3cw/Ho/cVkoS9pxmRImz8WyB1iLesA
`protect END_PROTECTED
