`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pZjMFGQdx7r7crf0ZWpz12FU8NvWH7v4BgbsQXkDuKeB92xn/VY1qgKZP6VKjpvf
hzKPLi7zGUB5p20lHhLgCBBBL//SQ1JYse0Yp52OCqY9b6QcdcnCz96r5TLPuZfu
4Sep4X8QTIMgIMBMjGtKUwNOROoQWI9XTOiW3H40l4F+7kZp2lGaG/qMyAcHeFN8
P+0t9khLayQ3P7v23VXdBgchCNhYfH9NQzkkaFqUDllq+9iANO7fzA0ChNcP9CnI
HIGIjbzERCy7lxB+A4v6W5iVbRL6M2X93AaiofN8KOTTF3dZOpqzUPZ4x+ljVjVP
30zDq68GpOi/OwanDTnZ0ie1SPVLd85pzBxirpUvQ0ZSlvbEJMsKbhf5/pDqthcz
FJYNaQOiuK3ZXig7ZfbnyWKKfNKvd0blBwJCuYMU/5YvXRZx6sh3QliQ+Z85dhjE
dw3kJ9guqIoU64ZCJ2AwusuDf8qsmkrePq6c+CC8zPKMxGAvQxQ7635bh+K0yHBc
ou34CffP9wvg+okl4YQTj6ETDdf2qygQFH8Q7lk0AD7bQp+IrzUkIalR69xnsV15
R6yALq75pDOBj8aAS915zh3+HhdF4TXkspFTPgrHoX++9hibFL5brw/hTCGAchRY
c4piMOiy5u9JYbOLvT5iS/r02o7uCyiHETwKtDMarnp3alrOCZQXQ//iGEULf7LC
Di+RxIPHd7PDhYKo0tRakuXMVANtkCDphNoqpwIkTVlFFSTnHnUzFlxaoAyUwYHS
cbzN7yBpXG85hurV9Y2FXvTJZSRHk+G9gamJp6FrqpPV3bI+BiS6shg3IeFB7LUZ
/DaGof/A5laZw/xwsc0DRr8OO3OLp7X5hKJt4D7CSVztqph0A9jhbpHiTiy4q/XW
4RloqVsjDiewEjaseh7plJNarrsO0svXSL6WFFx202Yg45ueeVbTpb+55/tuDPf7
IfoYLs3hs1E6w17Efzz6LbyoH0cznI5xRq2Gq5KlOFzphk3NxWsyPe1lr9nRb9un
n4bkGNcnUOFB99MJp6CPNFozZQ2eWg9oSVFOezdV7xFkrf9Bs7Vb9dONaOEEL5uC
flJjRll0ggYjtCLHV5MTUdhbP/XxuRR7UzPl4MaMX1TmFlnPRefXF2maQRytvmmD
2I0KEWOKEgwlR+67qJyff6uv4t06gNmMP73NCcq/qOqQbhj4lHpsSUNVtfX7qOWd
eUSWLzNejk73vTHRPXOdDBZ7Wzjgz5YeY1fF4joqyBBBmpoAHUFaVB81uRbYnN30
myNhquBIV62mg389c+rlraFA1Wifu4wG4xGuzJqzFMfNtCtxPZOll96bB3wDFcE8
UQUNTjTUlyisPOLG/B/uq5JKif/YDGfs9nvYuxPf1Ap2QIAJJN/PAHaJ18wgBGKa
ebuhR/JN/sdj0ztweoGkZ5+dK45Ba4WxOkyCKBeHdzrnYX8rHcUixMVmW2lEteH7
tcxMnC9SL4/mK4UpIO9zeHibK9Vk/OGX/r9ordMjBPWbzwA/j2iesqxWjiPpGEhN
Ou/9Smrw3tE7pP/1bwwq0tmZPw2BcHvm4S7cLL4aPxfLPYNURGYWc39JAUD4feMv
lfjjhvASmO4WwJ9Wmg8Heb+Khe4+oOTVHVxoEf3caLAbhg2qBt4ulhxO6ZWv8SVN
tTRrBuL09OwPMfjFxG0/8XEIIRFC0CMbWewHFEkSNBn5dtoQ/OxbLpTGupOAJri4
rRKTdAeI5S60vT+GVMZth+BEB5WB+vziw0v08HHybYA=
`protect END_PROTECTED
