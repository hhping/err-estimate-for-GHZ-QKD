`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4COGZhuVYRMfTPjxCP2v5RLW4TlMHF6SI/QTsn47n732T98IiBIfzCc/NQdnRgf/
l7LN+XK7oxeUzSnOqRtRXdrzneM0RWPQDnxKb8ee6zUFGjY19d1lQDFhUYoucSZx
0jngnm23CHlLUE2RDqjbsi2Pf2v2IilwbPx+Im3dVNK/8iI6lth+d+Q7rMQ+Q4Fp
aWGy3GhaUrdLk9lwg/auR7FVPb9wv8pdvV8D6JF9qw+0+FikySqmt1OHw0mRMxMQ
UOmyQTa+Zg518WIoqYw6MkTBxC6X7KYWsnrJ8ePg5a7Ow2Db7bsg4PzLfmFY3bwG
7Qx3UpHjhR5S+cMUuau1v0TCEWdu1QnmhVCfpp7/LfHxDqxQPirr8m831fxU96zW
FmBB7YmZwvBSGQYujT14DgiVTcVGh82j4tYFoIwgIm0=
`protect END_PROTECTED
