`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKeUjzZeTyJq/X5IYJP+2mMHg6pvdAreFDYXK2YZOsWyP/vkkht5luaO0h7W63gk
Ck1a0hHDyVBQ19YeeIxWWYP8uVnTiiNKxjDAIAtLPPYZfLyXfhk0rw4ERHgDumPQ
evstmPODcDdiiXPMbro7OVsNhretrQHklQ0/SeA6FQKixkRNGs9GMVt66EPk9OIi
+3tLIpTGZROalZXv/BfkqDddo1mHwZFSwAYm+I1M3oaPdK3PGV5fNiT0oSe3H04Z
Qu2PCLAzD1B/93klNLFYkulJ/giSSavmLicT+eRXb5Ay5guQ5SeMjZ/lSsJl++tc
N2cKnX0ckKhMZ60/FSgGR1FvqG6JvB7Dt2NLHaNyZlaFoZ9No/4QyUs2+I1t19aw
sz9nlc9GQWf0/MmwBqIg1tMivrVDOmpdRYffVEcyChntBHBHU6zxFNHFuW5AVJ19
2kZhHF6WZQScB7shzf28D1ybOSGul3AaUQPUIXiFe2yzJrTmYHpBBqrDiW35GbtS
yvqbgIVj4rMtrt/0VhyjKiKgryXD4MYRLTPN2iUYqJM1k1WISK9OcrHgEtVd7nl4
+/8VpAC42CJ4PU1azybsNgQo+iSR0gFgjMpWHcUxLn8ljsm3DfZma81RRjzmMgMO
3S4VJh84ke7nV4L3bV25P/BX3Ds9S5E5BsvRwOz4j+2VtltvfMA8Dw8+61Sg+IbW
w4EtyJK1IjYJ8tHywOmg3b8HpTmRKpt2wv4v5TZfsrr2YsUhbeBl9qN/S9XKIG5G
jnGdEEOKCyvo7Qr28W1r+1QutYMMuC0CFLIL13p8FC6y436+zGpT0a7uq1BzJUmf
gj7Q9OFauseURzmQa4Ip6rDhTmfB3FYITwC+ej8XZCg79pvQ6ElPDbyms7Bq+mbF
RVsIHB6Rn+jGEpkQR5yedirZOZ1Rm0TlMwzjNAjRk//7N0Bg7ZcxB/sq5iyWIUrs
AvvkA81aSChfecrvnsHp08+sclbJN5WIfQrZp9Dd1hKJR/bOv2UkrW2ezkeJ00Md
nsjfj+OLq1vr2XHJ2GPhtg==
`protect END_PROTECTED
