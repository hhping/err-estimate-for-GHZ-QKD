`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWxVPsEytVv0x4CsqxdLJvlYb63diiiVBsa5HCyDMDUIAiLGKzWci3/FwsSwcLC+
wv2JAxPxT2EEa8grJVIQjbDpLc9JI4nATRVZX+DkrSHt1h5Iv+YbtR60q0lI2ILu
JE8UCaDsWvB0dWhei6E/TNj3ABGSd4a54lxu9KG68jZwRVmxarKa4gQtPVu9D/fN
tDFGR4U3RSIQSBZu7ZlAF3fDVrpAqeYspkyBIduHfVc1DJdhZaP+LTyhjVKptoHO
5g9xUJNeKhSVk2cKrLX6MlLEI/RvlQn3Iq8t1vCl2IyddDd20YPNr8apxWAnG+x+
uFHnKpAlzq0i24GNI4er5gV3mBSb7GwFioNyMz5qFAv80xylLsI7/dgXx4RImAtO
OZ0g006ghSO9cCbcyObVkX7tRb6G8S8rx9e7ik0JMFlNqh2B6GMHrMWHg98FQZWi
sjNJTatppZVSH8R8uBIbmWKhorfFaSQcfH6PVnn/o7LhCnty596GUk6gadLX446y
dP8QxF05s9yrNd1sCzbmzX6OvCZLX0luJxtbIFtRIpjXMXayz0OobZz7PGoGmx/n
tdYlN7lHuyXa70s6Bh2avhsk773s+htfktD3Bxsbo/4=
`protect END_PROTECTED
