`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qTwUp4lLIDu7XbOZvfAbopinbolwg4v3/ffUULi1S4BoZLef26pL0+MJfFfjOUdW
Gg3eQzJHxsQnJ+0ZQ8VS2vNZeGB77hw7Hmh84Vkvu7K4Xinu63mQmZ9/YOs8TXr5
uUFjqCPm84EA/ogb/MBTHpoaa1MiIy1gr94smXeS/T60yIACbPllqg/s9n3dSKef
bmICWZVnGu+BVKvNqHATjsY6ty1FBim3ENrR8EF0I35V00tCPedzjq787KBfZJcA
fusdEUXEZeGILvvIbMKT9nTmFz9PxpAkB4yZV+Ijz4en3zYLqqfx/I7zuvjE5Vy0
E1YSBx3+Osl3R9kTw1yswTU+gQ9UHDcjnvHcx1UQOHWylkx1VhfPcxPWPvn6BZWh
d8PhP/lrkH5pjm1GvVrMrzU3I5qpEYjOlaLk+8VAc389S5CDD0uXxxjkPMuWsacU
Mq+eA8cEKUSby+49yb1FKKfYzQTKwAe/wAWfy7jLGz7AmjdQBMkYiqpTjUhfvd1T
0G+XfF18CfmQi29nqz4bmrTKjburgNyB+cjG9EJ2kPOHgTLdvRKDSJavpZ6dwe0L
AhnubrIVr4t3jr6ic6EScGv3yjhGkN+MUtuvsgpHKZ3XloVZUT3MN1grdfRs+ZlR
Q9x0opWo9aFAtJWB4GzpifCA6d+WiGwefXbF6SsUXcI8GiPcB+SRwAm+Y4I0AqcS
s9cZ1G1+DjpUc/TezQ62tYA6i1uTdo1scjt/15a71++pX29mPn5EopYgqWCWAGUI
f7cxw5XiMY8PdktMIl+vys0xm4p3jO4b4hmG9jUlX12lPkWQIv9rCdFKRzO289NT
i3WNYrcJiBZJacqCrtusrwISDduiHJ7vjY+86gD622Btzt3HsJyThpnfTiP0Xsmj
lfoN3WyZ9jp0MjFpfYk2SRolLFZspsXZcgS4EeukXUhsS/Mg3h9gTE4KuiMgv8sm
5jnUZWLFr0jL/R18XUhg+xakL3NAQwPX2Rcz6/4Is7o=
`protect END_PROTECTED
