`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ru8VaDrmm037+N8W47GzrfX6Rk7Cy6q3I5toH8hKKZXHoe10aifU+pdQTCGMz64m
KL769jkRljSLJ2U/Gnj0mCObDBp7ALJ3Xb7km1W16hhWEWbDgkwdElc4aqXPlB5m
O9Eqedzjnew5HI9d/B9+XHzT1qRCkJoVViignx4mApDlIO5eImIkgk753duyytjQ
6xAdDxJHqWKVx9AJD1Loq6JYhdfZN0FrS1FtTxac64BUy6+EbnmiZpE8K6PRgKCw
f+ALhRk7QHUHyE/DjW8xJR9RrIRVQMJ1nWZMK8yHHMISEjFlwdK1QIgV0/iXS0wp
OCUEcCs7oY2Ajw6w0i10s6L8LMZK+6kfo/jg4ywCGTXyU97D6CS4lXBVVgZdBD5a
vOpwG2gotWQ5U9khvlPVEnsxfy/Jd57cJ6LtKNAIQs5WSXQyIXB8SNjfH5Rv8nGN
GE42sblexRHQSruualkG3lpIG1i5s3vw2w2UoMa66bzHKG0BfYs9Yb1WXwxo3G82
95q7ws7svPiFA7elmPHcKkaGaKFvgqRnWfkJig/4yJvPpxlQMNSWBbyH71niO6wT
o9XmNpVREVJfyUh9bR/SbUyztjbbaCbtbAbXaQztfWh5E65+S4MUBXBx9UrORLup
aqzivziioltAowSuWD418FICteIbiFOkgNj920qRuN4CzjmfD0SC45oztg9/a4yh
98ZIQ1Q5AanyJqKE4iUxMWTIFlNfs/wrMNWA8g/ykN1GmMu8/19Y4JdI/DjI9pQy
jVg0vclqmNDJTBjgmr1NVQ==
`protect END_PROTECTED
