`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Km0ijWHdDyxAsRuyU9vCfl5aMfdG+be046P8wy0vVB4pBCog8dul8NweFoxr1vG
pcwNUSEx466Xn0GG9eTISdZCUuaSis4dNgIB7k4Xh27eMEQNyzLiKhXAh62AWjiL
TSptu/0sZzoneZHQpeEeKATvTtoaStiTpxIxMxclfOU/9bwHjZY0CXUbPtKBAQ2Y
Xd+i00OAS9vkXMgP7NNFiN+kUVhVyA05+hzYmkCooX8QH/aqkn9l5a7iCrj0aVZJ
YjgcxSFPv1+MD7wc6npZYJnHekSZecUyrhJ5jmuHZXaRzpUUBTxTD7H7ufMLSAf1
aQ9yUfsY7PH9xwIVGWN2AuwtS/JIJgVBohhpz7iG4G4JrKjzSxFt2K6anhJnOpcN
nh/4IxbuHzJHIxO3Fy4hIYE4wISVbs5K7c3PZsHT3sQ5pXFJm2A+zx5ojd8i5xP/
FF/6FlqisbFVBraLWOPXugk8VK6PAeoW5bXNkl5N4GCsSC32qOY18TB2fL1JiJgQ
aG9ql0U9mO37902p12Y62TvzpiJ0NmYxUkYgTMmJuNfdsXd/Eov9z8CuStFIiSjR
MdOWrPUiA3tPiuPiQaHDwLyRcVRY2ZSHIwC0ZK/JaRW5vR2TPfnlvWQtBCE3skgX
UrRlM2MMCjtQBMSDo/QdUwqaqOmn6l1pTHen98rFZFw=
`protect END_PROTECTED
