`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpYOam/RXLQotogxvGOH1kJxGDk0rFPXScImH8W1U4RXAHcQeuZiQ9SWQNKPQuP3
SAgS5m7lMZTF6X92GqCLtj0n6bgtDpZLgt4PsbaN5gFgpzQB5ArkQNNCxCPN5u7Q
OX8Rsbjlby/kq1398XISdpCZ44OlA9apAQvLK2BQxosXVFCe2rbwsQKHk9Essyye
5MFvwzDf+CbtafufbEidHabrgDw4xjF3ZhXXkzvhpFmOv9V3+i8Pfyx+HAea5fpy
Zx4EciQYIjiyh0IKCL1Gl79lHEJSP96aRNWXVr0jcTAZZVIuJXXgeCYYreAc5Ro1
22nqQQ4L1j8xE+4WHoopz9moMtD34ut1yrpnYEXoAH+dxztCVwpONj/YBnDEJfZg
mAOG38l7smEWelM5cYBL/McHKycvmaRu54RNZDlnFW6u/tg86exBRVz0Ks01C9r0
V1JhoQgwBdo3gcmzHO1IUVV36Ruc8LZgEZ1Ff8dqoJNdOotIUOFkb/wGOR+SUeRh
PsKmWQB02ebM9OWIXZLOGnx2mSN+Tp2NFqOixe8UeUatgij0Ypgqp0Gx9sAAdZpm
JlyMSnbXpnemoCuBiRYm7AQqvpdFm5/fE3FAERKVBFAgGoVBSutNtVklZ5SCu/3u
WDyRXG/BATy5S/waHTkeldI4M1VkHJBHQEme2NagQD0=
`protect END_PROTECTED
