
module log2_fun (
	a,
	areset,
	clk,
	en,
	q);	

	input	[23:0]	a;
	input		areset;
	input		clk;
	input	[0:0]	en;
	output	[23:0]	q;
endmodule
