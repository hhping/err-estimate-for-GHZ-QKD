`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KhvKPz81uSVZFumc3Mw6HIT9ia2aHLaWv48v37NNgcj+sN1AmeRGL/DdZvUbYsFQ
kHmULrm1gU6RVZNmqCVprUqRyrIhs6HNoIy6vRSosRuQ6cUlVIIclvmwEvZU2oM4
rDLQ35Mbq5E8KkiF3Cf821P5WHQJF342vypfMrBo25DxdUjq+ibeKJNIlWlskk/d
dfjlU81NqfGKn82fOFX9iIsCl0CLzJHpVaKGMxqzsbFPS0mow4+bRHXyoPACtygj
1TCZN+HGwjb4JfmpLxc5uJzLHhXH9SOc6aUwjAQe3nMs+NnQbz3KLjiIYw0uE8F8
gl7ehHlXcYCNRo97mq0e5OpD7RnRW0/Fz+3pww7jCQflBegOXb9lKd1JkVHJyMXx
TP2Ssdjm6rA/o6iW7xJBsEhySy1zqsGKYp47p66VtNOnL80AHyHjMmXoksBlxW5e
IGq27SvTfZt7ooZd4rBYNg==
`protect END_PROTECTED
