`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxIksuICy4eYLrAcpmniKw+7SOxaC+tmKCD/FDx2s/zH/Qk1h1+t0rkU7gIEPmXr
Lw7KqYABXuKc8qgtijWdePePGj3GcDcJrskyhzT7Po4PE0jAYsOGL0BeEJLl5RB1
1QD00F1mPP+7wbq70JGi05SPP55bxn4zapr/UI8H9JKWLcZW2Fd96lPmgEqemWrm
Vh6306nhtXBvoeA0d7KYRK0J49K1H7cfmfthnz/2BOgV6+H8fl2Vw3gJk2ATZfuE
WPO4FOPmBfCfJ1RFD8JJIz9eu5dgIg649DMGDnlilF+6senMUBwlsWFGY1DKfTpO
Gq4I5O/gEOMc2t/wTeY+jGnMH0IWonFotBtr3wh6nGtiP7xYYl/ewLnO2Dog37uH
mhR8p5b4R51IPyYIHbVPgjSeUs318MLMemQf4qSa/IKIB031drRdDn7+UNC3qz/Q
kizR6eep1hoKPADrcGMFhTooqT3bEkL5jPM21spoISaJVv5JUDrNq71vZyYA+HD8
7HloByBhY80izDkLWhUBiGrhbAdvLE163Qg0KMVQYC1XVWNyT0TCiZH1lmDWIV2Y
j3J8hT2hnpqc0VSsVNd/nlO8kbdZi2os8UXlM+R0ygobzsicBhF2uLYwzUmSGie9
5g+wuVDS1LExfso/y9A/v3MvRrcxVo7O7ZyduTsaOOjkhIgHhljLDCg3G7J8yFCl
j3e1xfazrknDNWalZ3/vOa1CrWitXG84S9dCjs0fns/nbHj0eYt4+5Rw86YKqDHB
PfmNWWyqjrmFwjXNzuVH2DfbMqrD35lqxaUMtoch8kHHTg7UilRAmmcnuUORAPAP
4f1M6qZ4ep0jiXz8sQ7XSc4mBcrWs9RWvM/ucAeVLTHifWcCCTRykSc3GN0DjIg/
W2Ga0mcrVnEFUZbwSZZul69vHQeEYoKlpVdy8IYHg09nW/YxVA9sAbNzZXxrdyZu
Ymk1P9QW1dq6ewBNSl/Df5W74u9pH6Bps5PZD25vSyNMsTRM6lLfHgoCuxb6bHT/
1MHHE+tE0biZDvYIUUCYSPZkX7lgJLOSoCe5giYuT9b3l8MVCCbIsikOQps5aie+
Q76k1npukKy7d7y1tG2eTNR62SMeuz+Al14HmjE9+5h07vD+w9JX0grE73l1Qj5G
T650DIXvzujntxbrXgfh7C81rkQq5iXG24aVaT1S79tgR2f105eUSmQZ9khnqT8p
fv2P+9/HY5KIrIeyu1niYCLbNmD/LFYfaGOTTFHuNY7I9+ttHd16X0o8FZ/fN26O
xmF1Dx8onRaM8RAyWAMo+p7MWHiN8jodBsznXlDZk/4RoB8UD5T6BGaxLXMUHUCh
cspXRXm1Qbhy0bor7TVjHxcK9+qnsQHUDAiuXJ3we4hnDjWy+5ubyw5fDIoPpXni
dmd6QEiUCsHT5pylf+zlVKy1whZxbzJ5aAf67dY/qk+tuC3kdj2wDUME5LZr5FMB
L4vTD/7+Ng1wT0bpwwAwwlXiLjYG1C5LHLDpaTCaASMxogQJNv3hx5bB1/WbsBop
GqQhfz0HLVMSvgHLij2iaaA4H5FHS4OZUjibGDkrqM2cn7kb+xbyaPoMGY6rzkM3
98pDfqYZT9fZiTP9zqQEdNEM0KggG08Idyl8rmsJB/pM5cRqbmnKZdBEDLYHDhxR
YYTjjMc/FK6iw7n9JbpsCN77QWWqYnYXO9a2BHoLAVOFBDqMYN/VMoaiA2mIIhJl
zQ0IORlHDxpbQwpsJdYj/+esVO+5DDgQjHYVGParbJ9BdBXzFlZfrgIwAsTLZsT8
iHteOLKFAZVNxzMfRsCjhQr4Uwym/F2kJcY1j0ScrmR0KZq6TPYgo8fcsK8JzLts
WHVcVoGKEbFWP8QU3CVIci1tC+PjZ79+yMwIY97wC8/d2HnWBsNHNpdjUft5DlBP
bDuI8v5dw/wUhaPdNl7IIGRzt8dLSwQtG5kUekWdZ9yWj+K9+mhiEnRIi1Utkn7R
9UjENcu+usuxk1o2K9YrSV2B6bn6Hhba40Q3YUml509u35UGIfcuABAlz5m3i8Ij
nwQ6rNrVt7Aq3u6YkSX7ezabO2j/LefYhtP6c/bQfA2ijels6JeGUBEU4igox3zg
tOiOVxv9vUJKmUiNN1CPR/acIwZ/iiUN4DdonYQ1AyHO5Z9omzMn9EOLHY1BFRAK
Kb+nNlj7bsCCvBZIEu2FWKpqueHNMYfFCQJM7OZXam/m+8dWjyUXZV6n9ZYOQM4n
P/UwCcNEmAIgQPSQ7l9NfWTW+dQuhcxpooChed7lsBLG8ByVLjhhA6DB4rUg817L
/zDMUvPvtRF9BKdiqihd7xZKZMSCOaalnoa8rnP0w8XSK3pab/9kcPX1zc7Unwit
IJSPgpAje5iIWj4XH6KPOaV/1vi7sitJRyF3WMmzEWjz//wDWUliJiB8sc+oYxUE
ozSS4hiAEjmRkxJJCjGFz57h3NnJK5b6CvyN3VlZZl/dcqBdCGkuNPMJVfdMt7hT
Awp5z4Ra+CyRY1ijcVhwG07Yt5m84soqX994tRa0SFIw16pAn61I0k+VFkCKIWsi
XNxUecvHAbHP9qXkKpK1H+xlnlKI1xa6vy1ZG8o5XAnT6/Ezn5VgIaa6gMgrOS2Z
SiLE9P+R/cLWbMLaLyyoKPWHIgZHcBBMi11SLr0mIsgYIU47SeHma1lNIp1DzFBg
K2FCyX6VqLTxr5VtW0lhtOcvj3tQQNrEBOUNerBJkmnvNS7TlqDcQZOVgvH6VlY3
MTTNfY7kdVRx/eXClPGsYgiP9tvy7BkZr77Iq2jPtlghcrBO6FXtWelciUQNGm7H
H5rE4xPkr/6zAh4g660RkTkby6RqRAN4+uw2D9lm786ITt9eVLAGczDTLCJxBW4W
TBn/RMPE/wUbPGsMeOHn7Ewnu881R56HKcZ13DAc+YkRKyIGpX2hz6aZWKP9dA0L
35KWDnbxlPfq+e38++6/qYYaB5w7zXQmUj2lvJis0YabcZhvweaRaUL8bNxXYqZC
4YDjrknvysWoO8DsE8J7iI443oY2BPX68mDHvUhxTPVRSlityumSA93tR4ueoiO6
IRkVGKaS24ZyeI1IsP2oeADvoqh0ckuGKfDTkBzN7j47jSuJ3fYSk9q55PhQ+0KR
h5kYXJe/Cj2j1jOPYRxbNKmVzm4ej8ibkTqvogjTNDQtr5s/iDHjql/3nY+0j+Ty
bQJ7WYpNdTJnP2cXgK+2jTgheFr/W/4BpM6MvbZNknTigyTNE1huTQv0BIYAOv1n
vTjCB08mfNPwTp5tFwQQdgblP8EMLyI0EL9BK6ecu2CjnOL6LS+kLe7OS9HYbzkz
y3pr3kEx+9A9RR7MfwMnzkX/093r6+YSFnjqb3vQxmaQNkHkH7KlrjqNc+JG055o
3EygvuyhKaKKRFOZ4CtV/j7sCguK52ldpHAKZi/BljW9vngwk57Lis6TDG0nP4Rb
PaET19lB/x0Ry9akhjl2KxQjzJrptqLrjuOV92N1G9pCdTOBJYIU9494ial70UxM
W+fyYMfClaNr+3gO4XdqzyxTgSTY1/FZzmGv6pNY0M59/gElL35KmzTz53MRYlpk
Igm1idutu62A0T83NCEvmquIt4vd+yw9YIC3u9v84mSppiN0OSiuSemkhLq0aoAf
lzfmPDFEowztfTPUi1wnVkdQlokn9a4iA1dqa4tKsmY8g98xpbv8SlxqR01WzhyW
Zojr0Ba7nCIbdcKDuEQ4ijgfRK40RkXyfFZ2sM4jGqcRtppsRFciFk7j5+vfvQ8X
AMnrBqhjIBinWBaBD8aH05A5F5fJZc6Y6f3QpeS+r7S3ntH0Y8JfoWxn2w2z65/x
gECDz2CxhaEo5B25rGB1QigNhgMUAizae9Zb9lU8zyemK+iC+67rbDSpQyz8o96e
aEYmJzH69BsEKQTErud2YgWkUvP6bORi/gJsgVMTNEigPx25ey/CNrzw6JCUn0YU
BCHhnGisyTSAI+hoID9bY31ReyqEGNftk0D4yFjzP3yWLAl2lkbekaau3duXzDxH
KznlZ5hNCtseulMkOCycetHhTJl5EHHvPygV1ZpGmjQcXPJD179rODQzcRFJqkYO
uqSCwloEXZqySjZg65lgEH3PjJ9nZQPCoIGygb/kdEWQLpHw0JsH4B2vCWPOhHS/
QQ/pEZriv9VyAXPYwIH1PAyq97WdixHyz0yMpivrI5+VLyXfIhhNn6LiLXqzhScO
3auBIw/yb+vvtLmPIOD+uQqvil6aeZzQpBvuBy5Ge72oR3JJ/xvjGmbTSEiomv09
bFnADR5SYU+NdVVyayczg75ZAls7dEtZQtcM3R7eHV7/236klxRqkBHttc07KHHM
05l0eksPvf+mssDXohkmMdcRe1dj105ePBu5XS+XAz6hVJ3h9HNf+f953Zd4sRtt
hWNeDoLQ5Zlpuc6QWUCWxUY5TGaYu1adV31bsU9gCVPpKALxCfZl17mnS+3BJjLF
jeYUIOP+Z8/6I91AD+n277SA4reOfwGU/Mmd5B++UvWMRfA4VrgzKQRDF0ecAreU
7M9UEpC/0bu6PJAgNTH8aRzbYTqTClySwHy00qenApuwmuYeM/xrS6HzdRiuoS96
VGVNcOSeymTM1u3M0wTuiyICjsop73vh+XTm+xwdUoiaibLBWhy4oaeK2RxKuBeJ
iaSpSZyTRU/3es5ODlBJbW4jJFhk3wYjd+vSAi3GdatYZg+yP9lpxu+qdw3G9Ld5
YmrBrH9JqysI8fPI9weefx0upR2OMkJTyE59vb4wLaXs7ZVWlpn7h5n8nJ4U66uv
Q+Rp53BC2+t3Ey/PFRNAe6Nt0/RtTBqdJlaJlF8DL9FaCQKD/tBIDa2zWhUJWyyX
1hfO74LnW2Kqh0LYc8BdW4DuDsyZEu17gbw6pxNakPpv3VUAT61Ze9pm6evAHDZq
BZzdaHxDgiK3Aiv/SwHPBFydNNH2YaezU5wmyrmGR+24G4e16tvc9TnEvVQUM+/K
zGV5SpYPsexWPrhHT4AQNsWqwh7EoMAPHTlD7+RzK4EB1cF68o4xhwDPDXXVdpr6
c3ahvrSj/nJqEnspUy/olQ3rJagwt81vlBlIkzFrU4hn0BUdZ4zgdBbniVkQETeL
zuwTQUvxM9nBR5wVlfPnD2ydpeEODOlxHcfp2uxcEmR36dWRuyVIkjuJ+adYppZo
8TySPgKt/uTp3Ct0ZEAMu8YyhmEHj0ErouM73MA2sy0146CuweUzbAgBF8IuEFSy
vpF0hr1KEYVXuxuMGOI7YIUHzEC/oDMz3a1xe0VjmsOFT9iMFG419gkIiWQ3hKD+
INm3TTSbreCDZguP33lG7uTHQ2/gsr8glOlYdJgVzVE7hjfk3WidaA09u3RwGTHZ
EZ6kN9d8kRnpqIKKPv1yYjszNU4EeIkf48jzZgPWO1GZatUPBKRi/k/OhYch8pPT
jC8D9h/0NdD/xvQZkA+NDa4mw6tnXnvJrbuNhMhlsVsSPk5dks8IQPki7OHi62eS
+TNF6Ts1z5ZRGYbNH1NlCrYza+llHBMbgIqUbxWDmM/h9DgCVqu+mKjrbnJRQPlE
VvfSeowb9+28ztNMQjMaAhc1Bl+ELCcqromLeKY/jHzjWtjLGd5iKAtZ/qsnCRm4
0vSZNDSASvLNLjfoEcupSu1LqOfdnCWdd+GJNtXrgRRFVLJJ4XfVpLWq14eAlQxm
8G+pDTeG1xBL1I2yo7jHOyXSvd0RD5Wssitw4w9k0i1cGL6uNbHj4mJ/Tabd5Efp
+ZYvxL807k1wJzGIO2D6irHjAwam/yqB2a5KijNhYLhFYUEn5hg1I+F4Tbmo17r6
EcyxJjE64YA3O4PvAI7Kn0fr1dHiQrRYqPan6LAGx1JaAB85JQB8n/4eOR5gR6cl
NlF0FUZHpO46qx5T+GM9VvJpdAMUm6zBROqJyMBVQX5SHv/JIeqSnsaeXij0AfCJ
MHZCNM/53x4d5KJyTdUI+V7n8ZUpueRLdHNSnNnuQPh6uKhhJ2rs/D7q1N7nIG+1
H0GOEMa0h9qDY4QPugsHElhKZYQs6RpGbCtY/gkJGdIvJRWbxdGXAyRl406JbeuR
I6hEEPw78WOXF15B8//QnaZ1q8bwxgrTJhqliHCCm/FAo8KKW3iQbDC8lJRTQPZg
o4TrUQsNIwtCoybNiZ97mqPaBPWy3BTOC+9xjJH7/ypsXcz7dHa/HIcIF8iJpkOa
qrCHZ93HFc/67KK09FlNfbltAsL8fq5mY0e6zuYoA2YFGRcjwUM5iU2IwFA/1Iwm
/msOn8ag66GGRl8KvUrCZk2r4SMqij61I/vqS54SPv0m18NCdFBQLLy8EHdV/4+T
dPv99aF3wCLAmQ+VuQdi/BGCuKGuzTHtAK0XJlmgkzmAtI90H9Kpb6f1sojhjrvl
sLnDubyQRe4vyFF7NztYktoYAu+06CnsEC2FidEKBD3n9vPb6IQWzTgDGB8mcr0E
nU3jeOy3PV3NxcGBnhIjNbz6oNxmg9QWnGTIJ5Vo5RX8XCAMdMclUKhktTCgy2oi
1wKQ6Bmzbm0v6QUuOT3YIg2434qnXAFLBeE9cKzam9OOdvE2upPKdJbdjfKqgA9y
8nF/kEMO1/X8w2bF2PUjTy2AC+uE/WNeCZiw/8wYxH143xc4odEaGFF3OYOCfXBb
lp1nq2tsf1+NyOn6EuSCIozfy+AEU742mJ/enzX9DHLmNfCQwc6L5g3WqzddJXd0
QdUKdTnqDcwIRYa/I3cka3IiuAAJGjo01yFzVoh11JPyLvxXkPEyRj04F+qSwfyd
EGFnHjuQLDNtOsUKXxiJnph4qZONo9z00v+DKbafD2s00ZUCe1WS4EbbbWXeIV0r
R1G6QHpQsZ90e3lXuiViSIS3JHzSnB2Oym5U8MbtjwnaCspNdvrCv6rjIqbkZG+w
XUchWcG/jCo2+W1j0lEiYt/FPk5U6uBft0Attwuqg7PWNsF5OWR1go2vEoTh5LWO
vmT+9LoIAMHJsy1oJeeFF+BC85fYhGXe6/ojNAsx5uEl8oEYNzJRibLR/kOFbaEv
OwhPprGp6HISO5Xhz0ojohRVj0L0+gv7V9yHIibk+MgCR3dJMZZy99il0G5tYwr0
vtL6A0OEbFJrn/kFsshL85fXSK+WXwJGQMuwM6jnFuTvxfDfCIs5HEWQegI3Y1kb
oaysXAmi4w6QQAzs+FNKDuRqLOUrG1OV/IKJetxC+1wOrkKToPiTLwme4Ti1l3XX
Yqg43/KpEGjDPA7MKP6maBAqlmof6s/pWywk5glbOZHKCSMib3yhivltsRpFjw9Q
vyMDxRMOvPCqH4RdCD8wGLPLGhx2hTDC7kg6eem47jHmYDDKED7mo1JiX/A5fJHm
hgP31kwrQr2glwyEeWdjZesj5EQf1XyC/kmcW1G0h0GyP+1zBDgzGWa2bst3Al8R
ixHJzJPGINt6Baqx/jtklAGC85giZ4UsNe98zvgM7dhCkicGxnSeLq2mQyohOCt1
+5DnsJBTQghdFt1zk5jiVmQnMc0bx74oMr1wZ6liaVRJeO4TWXSWg8WEci/QgbpF
Wgy8z1es+k3RYTsDDH7xLTxXRudYh5Hxo7+h7gG3UrfRRvT2kj7wqRTeDOlotL5v
lsF/OoZx76ZVOaYd+8viqY2MkYuXvFRHC9ysg8nNa9CNzKa2o5Af6mjijaTpwjnS
szwVIckGs/7LsM5zAEg9hDznTob8XFpgBn8VCQtGhYFKAGKl39exg7jnaabiI3Lm
XiliOojxBC1X+AbQQBbdUuiRt1iLZmKLGcnzZmT1guR42cO6tNgMLYXvt8wAJ2S2
EKOUf37CGPHGM6JuckMvlKjvXIzn8HB0WxQc/O5DghI+rcxgrWeoTOL9dbqM4knt
bAvQUPTAY+YYC6OzFK/Xi+Q/vowe4l4SMyb8cMkPs8UlTyTYGM6bF/LglLYKLG6A
ILXDeG6aq1F236BFDn4nmd+r8unTZhtFUXMOP3Ctbfyj1IearQ3Fb5GHaEDE8dEU
nwXlZs2pplOTRsBol2EK/C6VUAQ8Oypy/I7GOUqA5MX5voky9W/3D87v5D9BdIWU
02ZAj9GCASbJbrhrVHdIVmo5m2lNTeEMs3qbvvWfQWQJ+jVpx+NkpGAlQJquVukt
eon1/0XvzdwZ7yV9fZmT6bvOTdc4feYF7yz5w+x6QjxjfKobVe/kwUJhkSC02oyw
wDnsArqbNKn7BNRmZlV7oCkZEdselVOlLtUUj7PYEy29ypB7GLvMTbhO9I9PSPGD
Sq5NdQbcXEWh7le7375nMIGWmofq1GTgIpE4V1kqEzJTTMbsK/vhRPZHHd9M6OL/
ZplWJ87nJLCF8Epk4vPVghEpl+RDIjAfKgrWchahDBbpGahoUvrK7LEiF+Sz7Dj7
I/B254aIhyTvf+rxzwtDjVub0PcjEpQmqd+jRCCo6HrW7HBqVdVpy3M1rj6BIvpq
+mEAkwMhg23IWsVdwz2nws/uMaOWfFTljrz/XZI1anN1asedbUlF/fKmPiI+ZBPS
yIKWF0edK4ji2UnpZ01Vqdy8FWxGpBoBHNBaCS4bfL5EtUEBYBnYUB4QkpeCeR1X
g0ZRjZHfZucPfl0fC3Xkrj+wlEHa8BEgAG7SfZDFgpWZ3oErseZzcR7+WzEVLGas
H/o0TpeOIrs+bAKx7+0wrxsNjBn8yH5hU36zkoCtGalTlMLBEaflKSNqkw+CEOdo
SYQwhUqVZV6UJjkp7CHXA/yLzMLdBGWO1EKyj7pCe8ETotN6Www4k+LY90JbBHTL
MchG9pD3tegm3iYH4HTDZti1esotaRYcwyMIT5YQYrMK/AnQtFSTTfcasUtF/Aym
Lc3dZ9IreCucWRHKFBb7Rodv1pilET51E9d29hYYqOgKHHjnELHegi+seoM6kaxw
q5h3v8Fb85rBLSIVu8KCsNevAVuLVDsoE9TUsdNp0sreWXCVHUvC1TTl98BCcWm2
RlryMgnRrwVWgQSnalHqSbptjmklX+gFnOoFMt33oshna4yhRQsaXWGppvrqZy2+
uOkdWRUSjgtEu/Fz8Yq14zuIwiOtcfOKhRJB0H2+WuzsvEf4QizRqmoN+ZnzCLC+
7ZJe+x+CHabLyq31CbsVYZcTD9o9Joo7+WDckgLsRlEDU1ndu9K/EdhFIWxB/eWW
FrBIR5MD0iA+JNmjKIRvifRCTTHz9Dg2keisP5LzqHa2LcGABkyRAsqjn19UyLuv
lxg9ghB2KSnHkyFyqHCRxLPoY8jOwgEeefK68ZaZwOPcfj/aCEjfkfHuYHRqeZLF
EGBVmLMZZsHhLU+PCH30Rccig/ZepTL2ACcsbVW0Mr2P1Gh3j3RpfAMUavc65XIC
bhOqQPrwnQxGf12f9slbkenSt7rB3KVJSW1rWUI46sG7lbv0Q+SXuzQ5tc8lnAb+
/XnnoNOZZVH4f5MzsXo/7MibQU4nUd8gQYJn3jNRLd+yzsDdb/1yOx/N+vZJR9Zg
gSHvveLdCuHzk3JmCO/FipaHI0A2tP6oD4kfCIBUYZcDLoKgxusvIuqbU/w3Gwfq
AZX9FStShqi+TTUK+4uZsZEXh0643Jaoj6a/wuymtZjXQtEqHe3zq6U1kEiiizV9
NJbr/sHnlJQDt4j260fc9M3BE0xY0K09zNR+vtYN+l60UUbn+ahqnX8hR9wkyXgg
QH50B/hm/Vof7u7r+CFBN9rmba7y0ofaO91tjHDoeZQ5JW462TYAv0KAjOnW/MRQ
x6GkFdLRMb0EZB2yUzMMgLL0PDxulAd3Y5u9wLPfohgtdwDpaLfXfQS24U8tFMgB
+JXKDXBhqIHGgB8p+4n0Qjc6mQ5B/TNcVHFHsolh97o3tLHC/s2Xztb+FMkbuPIc
t4QyCBG9HIDzaIM2rwzVpq7Z04Xd+0jGCEenKsTgeyzhj+h4omF3VOoFGXEaV3qI
uAl4HeMG1Vs8Rv+NX2xmVSGMBymo7nxFeiGW2Ssayt8LpOkUgi1XCMXcED+02iC0
PDCyJny/NlTTsy7m/+HiawvRdrJGVv3yh6uvJ4H+7pFDOApZwMx8ZZc2aMfhsue4
Oy3JInOb2d1ShtPE2dbF9FSWv9relGgVbobixLOI6JSku/gIfou5p6b1RYTs77jO
gsvunxompwmEX4jg4m6LwaD+ZmLH8U5+yRkbkUToECXpqTtRyCA9MO5mGTifznTc
UhLqHY4ZLykndIVvShTqbSmbt/tV8W+5d3peh+Yts7foMSzG96c569WAmFB+u+hs
KhrQCHFYhmUUg5IJksqLv/Q0oGg6xJtFLwSUPWIf4o9laRSCFozhMxACQtdOZosJ
l4DKVIurrMcPjMIxjtyjo4zfGoPvIlwqLE1Zlou7rbzPNKgZzTJwBgjRd4n+QXir
WRYSt/vqBz5g+zLjEyV5d9tCLQ/t499oEVhwIZRkYLJTjmvfvxTsRuxgzb/5Vztw
xkARaCk77Tv6p1POyPIYdir/RtGHWyMvwzu8J9jQQwQ4nMdhrd5OPqUfbMHgP/sg
DicSJUpIDqTuBanKUdhuw+U2Pu+ab9kfrSKLVwy0P8oVBMr5ioe2iozit9TgPgyK
mOO5BzzC/QzngFKqi72N1f76QA3jFmH8o+QXwfu/3LP5A3hApMdkRw9bUp3eH/6N
kIfYcMc1EjD9LiIkEdexHZ2vBBlIt1yV0QS3nLrmNLzhsf9saGnHJI48/zw+nknP
pgOs4kDuMPsmB6lN5yszdKw+fbswmqZ4dFeq5B+rk2vcGTtJbIMLpazEUU8pnRA/
LnXX7Icqa5tTtcQZHKQ94IK7X2hjU3igB8SH6GgLnAj0EmaUShiVW1GkUZqPbTM+
ENWJxR2JyWKUKseMnk+pQ4ukcNTw1R9j0DtGR0h66FHwZujun9kMK+qE0jn14qlq
Cj4dykVodWXKEA0XUvZOMGpi0ILBWW2ucKbdoIvcCUoE/4QXdCCTa3x3xxSFbXRv
a2DlqA0uvcwJqjnTknTbGc/rS28CZRhREgo8JlDnn4DY4KHG7+ZjSdqg796JAOhO
ol2T53CuK0Z4sWKHLakeE2P1dRcywcGL2CQdEiyTG42A1/jwUKOs/ZNQsfUhijmq
d4Ao2oVvIzz/fXCR1UA+34Z6SiXpHBKdi/OgTeTuQv0IC552uZCzEZhKK0dOWJTr
zhqfIhZNhZ/tjw8mOXiQcWLvEVp25c0eTrkEndj3TZlN69ihB+f62A/+LwkOunk1
DuqiUCo5lVCQxxNjYgSCppd8+C0/g/2NhYB5+ZYFXI7hHO5vmC1DZ/xnEYEpJCZ/
56EMICdRhOViKVXHm/ceEkj3jbWPQcKBHgkTPu3OyehR4aK82OFOdVFQwVfECR2t
hrvBRODAdo9MUbOKJ/JZDR8BdbOpvyaSm67WvCh4JAXinFoQsS6SVeWFYnKpRcsW
0QV63Xne99kETl+JQgyV7aEbPBXL5ntWTWKQEPqRj65OaMvJ9gJ212eTFM+T9WBz
6mRbcGgvdQP7PRjIydrNb/UCppAKf+4o5PqMW0MQqwSL6mxN2AzNxbnEI7i+e3j7
1AU0ul3+7cgS+NWJUjLSo+ITrSi5QxJhBnabqJ1z8UAOlV8RKfEK/i+rL4H5+hMc
ZqTlBC8cT/tQAK1tS3O1bSZVjPHzWtKDOMSk8HUZ52ADroFdZT6L9O/zyUrIyBVo
Qz9wfB/w4oITjIlmNKBGn6IcUVwD939o8Tlg8EuFFh6cXKBDngpa6vhiF13Nd4we
Vujx20gEFUOr8tIdybY/suUQ+9yPj8BD9Tnivl1Dv+P8qBGttLCRM9b7TmmRy4pu
SCbIGSBljdjk0pDqfoydcCmvgdMpgoItq3LHTLA0B7vHZ4eSFGsXuUtqHuTH8mrS
qyTZ7814Q4EJRCK4/V1BOMqpfA3bo43e8k6lElUSm+Kgbgb6Ou6FhhYPqhkMNc6T
v8mr8zEchVXJP97vnV2VcdN6rY/xEOrwFxFknp289bCVaQ5csbzVutw7bJmG6735
umGbH0eQ/giwT6N+s6k5I1uWX6KLhSLGrc0tzwUsWsR/agxzHzOWRU0KVMq/vCRa
HclI6RHZM0R44jd0XfOql/7hhoVTPAqMQItq1TcDYF7ofFQoWPfnJNb+M6t5ZBzC
gJOW9kuiI6Y71Bv9OX/J6anO8rpVIq5282eG7ywDSTxGQ2degnFRvSFWa8525eYc
KWBnFGgB0njq4Xn5/pZ0FeeL91D1OKweFt98+tB1W7UinYtqrF3QRiOWT9z0qG38
jg0dApi/QOxj+lLeot1nwxMAROB6/lfvm8MdcYPsvW/UJSF9Kv/jDl+CVPdy2RnC
25hQS1sJagA6jnIg7qzW7zOL4pNTM7LtS4hWJjAYVACnDCSqopkx5SmxP9v0ckzw
H2n9oVyxT8G372qF1W43Zgd4E//mo7lYxjCj0sRKTH0A792uIkG6cB2F35JaispW
++2Gv004CgaaAZ0CxiRppaadpdovyfo5a2C5ckBpaKOzRcFeeraOEbMHX+g1sL6s
pr+0V4lqF09VZx0mJ0dj1lTUTDbxegWZfMOnm9UD8aTzEjB0qKwBpCcwowueuoAq
nKy8BIBQNb8rfP9xfvv7RPxFNcfCj6CQHaQGVLIcLW8QYqwHGp0H3Bkd1gMyZPeC
fV8x/mohqAUnztm5JgmTC5alpulb0tQrdl8DeAgvQa7iAkmFgZxcXQKAdhideTPj
icZA3w0pOs6IcniW4G5g7C9QmilB8oQGlUiW6kH9vQwD2AMiePuE37dsTLFIEdNx
lmS6wnFO+NWBLMsEgMy3PmIJCt3QUcheGVjEZfwxIHToA+UbkeM9y/iDslmjB02a
9V5Y94ybTIPVVKpd/N55cfiKj1SsAOEJOmLHE5KMyXqWupvMSmmpw1jQJYn3s6VJ
j9WNjl2vayHqJ217hmqzLrNc5dyapiE/g6Le/qxI9DFblLgZ6HGnrc4U3CCbd5z+
syYurg7qix85zebqVXUDpkFQmMJSuUQV9Fa5aSyCGmZeaCLWCV+s3ptvOyHa9xXO
xg0WL7DAb+xjgit95AFildUkGQWYJJT1taFMd8zOrDxHRlfTt+ywPTRCch0vvSDP
GwwWQTr+PTUb7xKQgl3wHrkC/ewoI79TJ6NhG2N3CXLBX47RCyGe20BmHYkGD5tq
79Z+Fp6gSnHMKbRI1fZ6OMI0AbSHlGP/4PPmPotTiJfL1dzZIUm69anu3JSoVguB
yqn3w/MA7MAFJ9wJCZvB0QbtrpvdBZl4+5KwT11zdO1VTONP+NR/SzKb3MB4ljHj
FhbiQXZVcj1ZtNzXRjiiS8elFp9PuvfvpVmdY1tQId69rRBMekbXeFvQYGNLZEqn
vtrcIsRFxnIQdLa0Wff8RiNe0ElsIO+gztTgF7A0tsY2A86rhFZVz5nJDAFEZvFD
EZpl28V2JhajnRtEPZblLzQnOa1yTSTEissO9trXw1NTaKly7N4x/Wm/r9ZrAELp
gQjvSkQWJA3FJj7Rv8T72/Xkg1mry66e5EAQrU8R1woi579yaLhNhNs1nDGGoBkm
DiIpWQMhBL4SjaFglqERTcynWu7EdT41wdr76v2X4lX9UmAH1JSJWWsh172Cs9lf
XW/mVc1Z+9wHxgBV21z2cd1IRu8rtmZcxghVgR8dPWmqoZwzCBeb+i3MjR82KCQR
WzMIKbiCsAsQEh4tCFCjrpbtHc177+kI/BWlX/n/fn7mq92sh59uVw4OAfrliGca
eHTeTZDlpT82ZBSZC+31NPp67qkDlkp9Qf7LDLU6d9EA7VgMP/mhNwDKmSFdmTod
DAtEfDj+pW9AF0u+nsEZALge/sknfwGG0nPajeBRMsOiLYtmqXb/eFGe/UElR/dO
DxOlG+Vzrw9+8Lj9tLLkqtG5NND3LnfAYsrva9EeEaLm7H3XTXj8+vPcczH4/8BH
OxPza1lF3peOO0b1LcjFwwTMdDtp4kF8SqoKgh+dYnjT1rPSBDuoqWIr+0nk+W3x
7xE9NZGrCneGo1mvFYjjLDqVhWF+z+2498V6fKTMrzzdGJDHV5zN4si0b8f+4Adn
JTzbhsumsS9rytXQJOhN4quxxxrDjkggBtWZw6yx6eusaaxa+TVDYmzPLNA3MAJ/
59uDBaXzyr2LezH0NdoPqRau8dnwrH6ps1EQ/bj/hzDXzIGytFyRdBtJzIm461XC
FujgKmH02QkNSrfwetfZLxF7Hflm8IGIkNdQh6BgOOxoR46Zk2Lwv404L8KJlnGA
FhPew7qEJXnfL/KKDrFkVGXs72tVmWeENNzbxhMSabcPhurZBu3YtZrChS1ONaOR
NRS3SZx4VEJW7BzAYKfQyke6XZ7Z57a9jeev/3cCgYYtlERviOteMV+RJQZcWr2m
ZxbaHnjuo09EpQuqZiygxYCf7iT/l8fuqMHqr3BHcJLf9cDUVUN/OPVlfld0AKZ7
Nc04aiCW2gEkdsajRH0QLmvDQBiDmBo2zLGmbAy6p1yZPRNQAau8g7mgHmUOhUVk
EOvhc9h3yLLhubCSVD8ZQeP0AomkSpnILzwyRALHr/Nk3LxYZ9tDzvzqqrngE6iv
Y1JEEGybdQH40A4zq1tfnXq9dEvq9UCuJw8R0oSmXuJLDhlzGIKAUYkJF5Dpl36j
219ZBRdl91BNzqz2akcCP4pXTx4ks68EpflSCNqt5N4FKIu1FIBgihpq8J0eYAfd
LmeL3FqheEuIv69Gityli1TMCh4+2SB1G0c23YOxPvGRpwhmdu7yAQcjbFyI83CQ
p0gTlq4rDQIAwITbSNAFfqmPGK4YghcHANWA4kUU5kCARBk6Ie/Od+7PTfADwzKT
aDKJD4zIt+215rQEOrPw7ofjyNab8AldFJCmRKvKNQ830dk5HZAMY2UQpmUN2yL7
CgwI1L9a5ah/yGDmZFOxA+129FUZd8qgzhtMRSCqbD3pSrwxEqyh+ppbR9oXuQeU
eL/rNPjSQS6N+nbIKKfT8qqsfg0h/GOIO5+tWwSf/ETOYKgwSq0Q4q5GNCIZ3oSm
cUltKVZuLytg54bI2p1UJjPbvR0dJfjKewiglWYd8unixgUj+abAZ4lhqXxC8aqG
MnQL1xqe7X3tFyA/bPaFb0wd5ndY5uGHUCn/9icmzvbSxGXl/mygMwFX/1JJiHGu
eHGkJ7kvyPZW2s+6SqTW49bgkQxtKPOAh5SzoFYmi0EZYY+PKfyiLYp4SXKifWhL
qTgsFeGKsxaR0PyYPGd92klm2w2ok4kFPc3m75OxQbfwabn5FLh/5ZPDGLUSmdom
cA3pcKXJWSl/zpRuoW/3g5jOmbLe3in6yXcTaS8EtgrrsXpDGdjNQbrBmTW/Z1MD
E/sK6BsukXRN60IHMAdOZl0sL8AH0+SwIhSbJJ8hBQzkiaFnLJN+sa+AZtZFqCFJ
wsy+yGyjL0HcpGdsIhRZuvaQIgynrCz053jyRzgrxCWLR6sgHAupDCuYxnms8EmN
BzT7k60VH2lefkJX0i5tPl/6NUtDp3wJFq3YIB96HDn/KeYoJD7GPfuCA+Fl4Lj0
3/keH/8ZFGa3KG3ZaEmDrJXU0S0w6lxAOg2KONr0fvzYSSPFq02nHIxxmUJ1VoMH
L4tmnzruK826Up1iC+ixuxH1dwlvpI3t4gLGvWvuhF+m/q/VT6qwEkVGDIw44WE+
774y8mSIMLxaCbIF7OQJQWKvdlTlvjblb+IHUkC0y/HxVQrf5aIzx7nDoKRizYfX
5VHuOUyKlX50PRagfVzv8PmoxUWhvjV905edIWkzdTeoB/TT1M/+SSsz9pQkG9So
OlTcJWBRM6hnbXRtIIr6i0P4k5RPCf5YabZnLCi7xeNpd4I/5B8FG1qeXPDFkR71
Miw+zkCoFlh2wSzHGpGgn5tfrAmwmqMbI1POnYu9V9vnjO4m7GRWXN1qbTdDqRok
am31eZeh7bcZ9gTs8p1BckOGcMCc+bXgWgvnEV39vmaVvABSE7pclkyWOAg3HAkT
OGq1d9GMOC6v2itl4jCvK/7kYFtWf4fZ3Apg9Gn4ZWZLV87hyiGaYQoxD6vMovY8
FJmNdoAn87Wveom5dvRtjHEWqRgg96vwsw74V4Rdg4EE4jRezYF+e//plyNNvL+o
rd2rvojWzVdkV2gfGqeu2JQxKqUEQV+Cy1UHaOrKvMRTLH4Twf9Ve8GnlfnElmcT
YEC05nydbh00VaTK4Y5+LA+u4qpkCQbWyKITr1rY3NZqJEC7Cv/ZoEgWH8hDKGZ/
mgYLa9SZ1VdZKRDtLVC+vl6vZ8DXIiEgCffHpKoMstpx0hXCMjTqh/c8A+VpZe13
fa/tRivZOqU09kRVDctux3SNIHCCA2k1LYETDbVu1hEvzbrAoAIdJUFGDvVX0F3Z
SOSo7PL7J2kGpSfVwQgt7XEiacncueSpuELg9rsz7VlTPeB+A5W1t2g7cOAg8I7k
G89aWTtRpaXpHtPC7EljqW5iFHZC1cymJk+YdkCipM5Ows+VTTWOpnT9+hyLJTun
jv6KJIZJWnzWU1EAH8jYOCEiMxWwOXZwX3Ha5p4/j0ERvtoCiFybaeY6wKkJaoU+
jIC2DzYJzKuf1Wge//sFCYCj09ks+QX3MsBH3yPwZC0SA2TuK6VCKUPkwD/6MhYB
TmYC3Xc2AExOAle5cDtp7BKgwXymR/O4I4U1Pz9OE4odWkPU2Q96+btWcxW+iA/q
INfFbCAEdIO+E1R9RDTlDtZSSPr3cBrnnKB7EFxI2O3q7qPOBpVu0hOQvKTnPGO6
ieX0di35olxwDesVcNlEm4+hi7+DDScPQAg/FYrTNIuHtSb/xAoiL9h8IVU6bCnz
fxqX4nIzljZ5piR3JcBIoUWRgQCv6pALfG1enOLV97/3QOYt2Zy/7FfE35dL+8Hk
caIM0ZxQROjjI5UIpwz1MPGrvYwECS53Rmn+fm+6H2uG0bMBtxkypKx91kPtbbwR
Gdm5eW5sr9ASJinTltY7gHQ13/hiwi692xvRL0oR/J2XivXZdm18sW/2lZGp3i/3
V6SUIH2gwKvP2FoFuMBZlbLO7UmAvRPuZMoZrIxNtZrexzIvaGaFwgIT6NHf2NPJ
6LR4QqBDUm94dqIiHXr+vr7yc5jDNv/733rFDSP4HxCbwSDXHLo98Afu9eMMOKFZ
FaPrTxypolKJAtBPaTS0e+mLy7lTpRQsB7+mUUdTYJeON0iM+KWOhRXB9sJ96tT9
bEPBA1jYFnv0cEjGMmRRJLngeswu2GzVxaHXCAgVsBWGupYfRdh5cFqV5+sYNfae
RdnMxP1XvYN21swUuUHuFKyePJJe2Rg0o6bJlWADilVgMZn8ndw6NbU7ukcekQ1C
Hgmu4k6lQCkoTBcLcO4Fqv6mBfBqqBANSyODg/DGDXyR0cIL+7sTIBwN8z2YX3Zc
s9zQqe2/23eO/Pur19XJhbyaiwTYDtilSbu/TOjIR5v2yhbvZD+FN8fvqfFk+Zvh
m3FBk0WZuiruht3KNtrj91O7WpD8RfllhMWITuIlJf/sEk2GJ50oRlemWO3yszVx
ZVwFz3cs9m/9AXoEW5TnYqsjKMiY8aDp5tWnLnqkufNuhHo6YiWPYq8MJc5rYfcE
1YvOKOmIRFy39mHAHZVzbHai+U7ZZ8C8oZQ392zlcKw+0RPe6PRbG6crF5QoprIc
R033AK7J/a2QL6dc7AIVlQAnskXx2ts83ujjPJUY0hzSYCVVMNyX94VlEwKYYnjv
XB6BpGX8PsX8nakYpoBh5ipBQObzHpqmchluCteScu+TxKh5AGYBxbW4qNoB8OBX
pe6cL0qD4PEV2gg7YUS/ynhPN63OYyt8hg17p0z3R0u1BhbgIlXJiq5ZLlfxhqkz
VnRmCebHi+ssjl6aYvnB6f44mQ3TYU9DYDZYTI8yMHpygM82269wc+7tEG69Kqr4
q8mm3FFByYymnMKzK7d4q6SleePd01GTHUAoUbKrJLU8/AHElNGHRPqOJLMVusvc
JEbpuKrpAhHLzpDWHoAf9/tsUtg+I2DmUv/wSEyUb9zUBbp/aicGzw6uieGqS+Sg
DclXNvUithdA5eXy7ZYjc07v2BTeoxbmKdGVOwWDJD5Bb0FdEk7d+mQldDyrPlMT
x+dz+JOUxv3eLQ7KUdMPosAG8vrDDmnVbD1b3AjEGKSxRIPQJ5a8TIturxGJ6JPB
Tw0bcjLGicqbgs/0JjU94bUDzfQOigvxrkOH1n0lp0UXATqsiwABIwn3V7WnNkpH
DNxSdSGUk6DWns1j8LDR1IRWdKc2qXY2b113Yt+RsA/8u+6L7IOdONy2VBHWaNch
kz6ZqwXDyH//jWohqUb8kJqV5FyrADTNRyv7P0+pUknpn0U6yJk9ubx8/UkOYqLM
0I+mtCc+S4ZzVRsnhu4Z36/9I1RImc8MchzTAYmNvNhkmhKcaAwXWu+UWoSxDFXY
Dvx58rFVVn4OxDcdEhjiBBQoaL6qbT4Ee6EUIOdKq3UzSAGiobF8FPg8xfjXrT5X
pDCatP72f2Bo/YTYRqhtaKAxmDXe2VVz/bXfkYUHCbjLWyUbrVehhWvxY3nIQXUT
oX+1U9PuEUvKymooLOSqrNOCHV1W+ammhu/qjPiHd86NDNYRps6rnxjLwZQXZ0+C
SuFGz86Nt4BquU2zIq/tHWt6VtXzJKr2OJhy22+AK/NEZNtG9upG+fqlscg37/wx
LkPhy3YFyvw1WujX5Ibwl/wO7iWE5U/nGOJgweXVkXeiWqBKlLHXp+/jSW3xXaT8
LRRfMZK5NH+O/o2qXq/YG/qg0o3Vzr8aJNRbKT+PWGTYyajUNvOWTkTcXiH1S5Uc
Cg3VxqpXP0z+Y1jyLaKrh2av7hkrhbwTNt0+h8nDsiKFE+tA5eDQjAlO1P5vhOsl
f8Z/SoSNQRZXJYGvONKOu1PcP63b1qujtvo7WGvezvrvSA8Dpqn5/utD1lguyhy+
R0i3d79oLhTiccGIosE/3P0y5oIrmq+XMtNkNRZ8jf5QsrSzYtidC0QziFxeFILg
X+vW2w1Z5BemRtEPVTmG+au3ZJ4V4rnr60MZPBlgbD4Pr6tjue9UuPTjqLUENOU6
js2/NTfq81fNXojoT6eld0EcaktOFqjmtBZxF0OPcu3nT0XrRYG+a55lFQnNWqcg
leE7ckdsE1BaG407/b430dipKzH2Gs+PFTMtLOCahVlMX8BNDWoYnCzT0llhSfyz
g7ofd90UxcxlSQ1VNBzF/Tr/8hVs06EwniRAFcbO9Sol23dqlGx9UxJuF8NVHsTQ
NmuXO6coAHizJrvoUQKXtJ2Ev8CwrDXEzXXunCDRZGpF2UlJudObUPfePw/WNP2o
Tk85+uP/2WJRYzWfgEo2YAaAlLPw9yA4Dxat/QL/LcQPD7wQpX2GNG+qMAdnM254
WWJyks4BZDEvnh92VGm5cVTfBG7SuOZWN7iTE6TdvY0liUm9k3Qu78+PejlSkRkm
6G5GwCMxLrvafvecud+y/ZHLjVP9sUHhazbAkzYx4y+Zp21RYCGkna/6j5K4fxSF
MOvkSyKf8pyzAlaSKKWRn17VnJDhHdykS72GUdw2V3rKcgoGO+d7BFG2owXOooIG
MbSh09mANtc2Op26dbz//i3dyjL9mbZ7WbtYHqDwOqskLOKGiij2vrSa53kF3ULO
wMgWzMxP9O873PZNPCfWg4c/EvZdjXBHMasglsrNb+7LRlw7TeUSZRJM9xKnmiie
9AW+l9fjfoRj8l5V8d2LhQ6W4APo+o2wHEchtWCIdowtpZi11igZyO9/Fy7r/txe
m8omXF+bpAbMDuK1vkEtckAGlQDtCCnaC3DmoMvgJLfoZeBHMRCQ1in9YkZYMn7c
TtL1tX/TvIQNDnjpUtKNB2GP/sUaVmQUhM/oYgmaOKg1LyD5z8NGJyKg9o+JJyMM
lhOkXL2iQEKPcheBcmfWSo7j2oWKfUI+tePqoTxh+KD6w+1PVP3AvrzC2DJ8s78R
u2rn7LnrJuyKQ1wSoGwbSr9grjvWlv1/EOhRoH8y/AFp1LsAi9cPbXtu6hmhnC4U
9hXh+oX6ok8jCYpER/j1xAsgheZ2EBFNLjhD6A2kEGA2Y4kKgvSv5MxbM8tUVxue
cRL+rwwry4Qp82BZAEDMq2NLf15Xqil2Vbu56QZOwSJiGpT3MSpdgVwmbtSECVhY
QeHOTkNnKcM8QhIzUTZ2ID4J2B923WrwykJjVzbm31gCEGaxhXsu7a8mHQRxISSO
+Uw++rKz7vtnDGR2yiEUELhFH0EJVKJaYY0PqH564C08mN8r9jmKLV90CT7Q22q3
tbwWlu4oLbyjNj3lWhHaYAct7sNJC35jDWbWfk3N/MS5GenTo7N+WROtCIVlNNZR
02wtqa8kE82/4u7myx1TuCVXMXcni8FX6rpfl80CWG3+8WLgmny/SavIzy+Dyd9s
u3uGOViJc8n/hUpWusS7DbZxpfqcHr8S01il41comMK7VibuTBatdkJOtuVL7qdg
DFFLpHxNeL0I4NLPsaljZXeT3Q3HoftHHNpb2Hnlt2WomAau8wKkKbQT4aFXIv+8
tq6D+I+dC0pKartmKJemD0dAUpOE9jNLctqeSN/UKyc+tRTSl6vqm/6olhQs2Uia
33QN4AFmRlPVOarJ3GTHVhC0lmz2aMfAjRRRr6qFpjgxjs5jNvQMsFQeFeZpCDvf
bSC3/V5OsMPn8v5t4DVY0oUyewPSglzSg1KNQO5wVcl7sQs89ZETKT8tUrw7GdYE
LqkEicc28xlfZMEBpcLQ9MnSsz4oBTtkdrxsk9+KIMrH5aywtLLW/5nFDFMlDlLm
xP59z4smbTvafEpOHfEcG9tQxuH6N7JZccqBGLbbGgOLFIoH1LkpY4SVqphMmWhD
PqRM1PF+EFQB8EnX/pg/2C9hv3ERyTNHAnBfSEjejpt8GlyDWpp/4Nv4uoWLvjGQ
iS2NmXMoYBy8Hm2awDZINWZbPPzZI2/rtNkZc8KO2lkY+RjqfEuKq0MpNnhW8YsJ
7aE1vmM8paAHAIE3ZRg/on+PXguHWS3Y6sK9mb1cXiXBPX1q+WTBwVM2N6Oz9yY9
18j91xEBv0wXhCQ2zKeFSffYdzXoOPyK9bjTLxfYTtneeC7XxsWZrV2/J2Ixi/pJ
4L1Fw+f4xx9YqAuzgxB66UDDnSA2ho1T3CxFVdO2jsOirfZjoEevKS9KyZJK9V5Z
2mLzJFZlhtu6xY/psUT07RpP29t41tjbPWdq5Qzg72wBZz6Pbh70DwWuZgoEzE3/
BeRfNL/faI1WTisjKAFmpjYBkweYmpUHuu3Hfgp1PlrEJouaU02edKRBV1pkJcIN
hBWXUkV4seU/WIG9AClhACjObUniKBF42Z7U+kKMKtucVCX6iN6Px+vNDmW8fogi
wszSzxu0CyufgklZhKKxL/oxlVbYDpWmwAm+5t1uz7qF1F/PmQPZV4+ngI4Pu3WA
rNn1X7JuYtW5yeW7kfSe9wneiOy+G4KmcEfUzuuVlxFSd3v9Q7LM26qF1Mqkv2yJ
qc0VX0gvgvrmrJF+YIv5WKffgXO0qWDy2//7jbMnEJDdxgYXoNMOpDQKC4vjbZAP
3cadlztqqQq1LLYKQpUERlHcrKSL7cFeBZBNffVS02mAo4NT6PaeoGpzATfl3E0r
XvqxygdIo0rT/Ei7C6bkJlc+1fB11Nw8spcvYibqB1Flba9t4PYRk83PcFmy5BLM
zHMgaIjZFqGG3zasVOtNifrdf1q1xJHU7FS7c/o/7cypsfAEzKazFFzUIc7UhQaV
nPXtKwstMOgx5ddO9qAi4L4mfIPAYw4+F2XbEZh1Mt4TtuOsZf1R8HcBXBzfD3Vd
eVAaws4B9P4UlfHleb/RbeV8NrbHmeIvhniS8b3V+URhCtv2qsZdMPM2m8btHNHt
iS4FV93gZj4sBTXf4zdOye3C1jiJfqWoNKwKUZ/kC/CzasHQDuQUfN26DDytFpRL
b/rqJ6Vb+wYk9NeC1fSuEz4aqHmjauLfcXCyGvVo2ihIa48IYfZ/o007V0cW/Oo6
68wBgzIcbYflFbpNz8gP0bmavQ3NNw1v1IRS8u7b7XewQ/+BURznhDrUr3HcWeKm
lJaBZTyP6VjcHxu6du0PXOresYyM/J39fr4h0e0M9TRM5YkZ6cTMsKtnfMAFXbkH
giDaUGKBp43Nq1cv8E6Wi/S4+dWw0M5UGFya8tP+QSkm9NWU5RLBLiv7peuVEbnS
pjELAeLKKXPy4jQ27BqZwtl/4blY2CRTaqBH/kzkbxL7zusZcwC4H+4cv+/HORiI
7EkFobNeznV9FJE1MNilSsa2imUgGOUhThIJxRC8PmTW0u+qWnqDCUWcexCfcuF7
tWLalXwDU4sKfeaaws7+ApA3nyDPkor4+Uxjvp/iMKpSaL5jOIyFPgdL/wM8x/1C
TgfHTL70A/DUz8SG7VnSlC2EYzj3Uw8EtJjsA6rF7qkrf/qGDXj3QWMg1U9dJ8k+
lWcCKkV+cuXb72XzmL7iD8aeI8f/3UtwatAOhGsGhk8SwlH4ubJjxvNzeeZ7qwiY
J31XzPgTccooTfyh1mwinJI7Nikbs5nu49c9YmEq/gkzu8//xXAGQBSgLhsmucjG
th6yvIx3UC5dFr/EwXOGWQTFmDnOcx8UMEpf3vnKglXWTYCwdORUT6uqRkN81juY
1WJsI+ljt2/J5WbttHKz5g+egrip8gE9GrNNRF6gHHuB/esAo0dkEsefrFTD0Sfk
yGLyqL+TfuQ0ycdjbzXEdPZ4J1WCUgF70OElROKhaq5ePmN+4R5zLnAUlC0cSdPq
UpFpbCMJRiBYEnKlcysAFDBbw+rXN1TX91APY3TbTUHXZfavYb+456bO2+HFWBA7
Dcj9UQ59tWy3FXvpATCtPyRsZjbyR2+XyJVvIrZ5qfn8NXgxk0KHlDQ3gncyONLP
MKYxrc/WrtvBSyeXu1dUohqaCCV9I1mh966j7TyeyAtUlvbBjs/mb6P+6lwmEcTv
bpuFiQ0zIK15ax+oVJ1Xc3htSfOM/MhDG4RcvTpIqFZurbW2SfaJNAK9gkKyjGs+
GpUoY8Mhq/wL9Q8kRaX4Q7aUABzhN8dKTwyndsOQIf4zLqUCn8w+xr441Ff3EhUe
NlCCujZSh4ZMJZMGMpJallT55QFHdOeIWlLugQ4LJ1HN1NmPYDckvXK3WhbRpBwU
iKkht+ytoJpa7U21UjKeflWh+0U8c72+t6GeJbGwySPVTTk+TtLgqVhpoejhco17
U5GZs6gH199Ru9201IEuEcek9GQ47L2N2n+03wkkc3OqGdCKTKY6gCBzewb7gdsQ
7ts+lZrcK4IrryPKRlbCpg5GtXFiC5k6/OtporVdss3aNpKIRxt/jNRhRvzkLE3I
LVrOrVldUBC+nYTG4vch0Xy/sF1cBwtcLUjLaSR995iOLChfVd06g68QJiTG7qzH
DtACauJGH9nhSqCYkG9JRFucPes/CFQLFvTKx72cZbvVKTUCAuU6lp6fYeF+sRhz
ZqOCsXVECuJjyX4XWMt9vStPaXrfOI4fehysTqO3IuqtPu6dAMV3YiUv35exJozQ
DjMuWU8U9+5bVFwyL88T0JZ6YGhj4xHBkJu1uaIu711A9ywIWzN5ujUdLwYeXnL2
LmvsH859o5LGyG7Sq9E+BlaOktIqn+QbpwYyNSAwCJnipgFS+JfOKVHiYdISjDlJ
ns0RALkkjE5SINYxpzQTjSNoTeLMwfm682coUGReyjHq06bF6g5vYFPCXE7CZPrv
YeqfPjdYhk2HXOwT/aa25w7bevfUIPofXpdYpc06mgggLx2i25OnhIpYQl3cHkri
RQZ7FrM02A1DaBl12iMqugL6NKkCsnGUECOPIT18V/FNEbHi7CBexEnO32MvXtpM
LYZygUUd8mGwg91tSgTI9Z6cIcD6QQcqwzum8LTC/OPFtac4y9DIkVVM11bdwRHQ
8sz/hXVL4AIUO0YqN827qA/TBIjgkv+locrQ5Dp6EEvB7TIFeoCpyP339TrvVcgD
2NoeV0CfLcPUy9kaaz2x08LvcnTXsaOn6Z1LK5V+XIw/rmCZT0YwQp98xASrZyxf
NnHSHJQDhTJ24ssffIqkItLIvuEFoyLbYj1f0KKM9nyi7avuvYZlqJW4VEkrXDte
JsnaD5vrI9I7ZZXWA0+c0OoNl/aweHelTvd+OCl81zmBnRqEyWf4CXgYhiOJ9sF2
E+qBb+cmfDnA6q6EgbuxxHhx3lazwxkc4N1mKaOmDJ+7wiyuiBCQvikYuXmHsM7l
s5GWUaJTbABerbjQ5kkJh/pY1RHyuFtDiDmuI2FQ8f6Jqy8T1mcFwHjquQohHhno
u5+oh1JYB8yAtzhhfQejG1qIUK519GBi1eSZ9dX5GPqlPfNh13JzAiuozaNQLC2y
001GNq0LJv4W6jwS6KMevvGZbJoU3oh6Tpo0S/rdBFhVTFuZDE/YiiN49hZzoSen
/vUKG3TJ1wiVdtfsZsOwg4IZQeMBWx4WE6LtFUBd5ATucn0UOVs54k1AKN9TlmUx
qm9vvapZvtAGOSG0qkgrlxGWreDDyUwynFoRhS9zKnLkmMDFpaIJw+tq/pZFhDN1
vgLI0tb6Ynb9hXz+wII9oM9tT2LsTTvcCFMNXiFYUKzg/BGu0Ul80LScuQ46flgC
Ot5S3B8V9qDOTAhCImyrSST5X+j0O9dcBJIY5oK83gtzV6AFQJ7YZZb5J0T+7Z0C
bz1QtTEPUVhDA3f+yKNoEJXcxL835E6nP4wM9zExo6T2GR2qpPMlxCwgIwkjFe4d
2nBw4Wc35YAT7aUrlqL+se0G5mhGKp5jbrXBtOeOhTE3UgZ2xY3JFdLMt43pDvBY
o5HNjgZSQ6YEghSo9mb7vhQNjat+GUTKKdUBVu86o7D560hJ3FJVb0VMdSbTrdOE
hw5WjNFfm7ZTXdI/gZjK3hr374hsa+xLhA6KNeU96uywjUtjkp/VFR4QjVLMBAVv
XmF4L9/1cF62csn6AmGww+QDyCyoO+SXU5HYZGrFNvN6iy11ugu2zV+xb1AN9Nyz
uhiiE8srMrLOj3VD1GfV3wWQIxyghFKpvE7/Rpo7h4GoI2K7JVDrfWXNxoipjtj3
ayUcushFu1VhDq6bhNVqD2DdjU/Cia36efJe0NL5slEz0+TGGC7vEmYpmHqUmRNu
xnJrclSBnRSlwYRf8cKGZOlEaRW3jvgi5xKeDeqUzNhqwQndnYnOLSNrUUyKMEoa
TZASdJZ/nae7tuWJWVve+cBB/IyHc6LC6r/aWpkKFF+NvfEVOC/2yusvzzfILeg0
1EB/OfZYjjz6fsDCU+YRlFnI6uxhsPTaotd5bRIR6qjudInljA0HEBUE9aRjmb3g
VrMiE5PPdeT8yINtqWeuz4zD4E18V1W127ONRjzQvuaYZc3snprOmGHyKkEfQCwK
uZ8PSR5vhmEMMYzuLY08Xfzt9FbYKay3cSHV08pN/uJfH2Y3oF83CwNAmNElqKVY
NbB6Z2mDBsZCySyAF2/FwPA0AHDGIaNc5E1MZ1You5Jo5PxhedXfXRg1AIls+0Zm
fGgj3tX+JDGcBp6PBgzXCv/pK5Y4pDBPggBSRTKwua+5Z96r0sNfD+ge0G8Ww97K
+/nuj3a+jQXO+B/YecbnCsLvgvRyj1fJjATpH1nHHVJrTx+1v9Zv7QqRYP6JyX1n
lebrJlTmgDOGccjWbHqS80I71rOlA/K9BWg79xW/6T6HYF1LzgIRMR3cvUxhChet
wzpd2AvlzPC0bObua1QCSvjHDQK195ewiZnDioLShMwOcVrgI37P6Cxh7kIZth1C
w9ybz3xZ1L65DzYbT9C4nlxJh7reOthipIn18yzX4fVDhisiPvBptsXCZZdDeDIV
kd5ncy6f/XRitXQ/Eh/Jyu5JE/5YAzqpkrnekkl3XaTHHErXzPaKtWfB4t128cBk
2E8Npme1GT8W9t+cHlDRai70eofmmTBZ9vnAyfN0j7XZXtJ8ljA/MD+6MIyaDPoB
evBta7970EVBwFbvSa9T/X5uF03QCcgq5GDm62HoxuvXRLGxulj4FgEQDQUsFdvo
tdj78+0Y1r1s+8a5PYlHdD9pz9qNmuWn9aXWHeHZ4FJlq/wSy02Jh00dtMxeXCx0
sO5ScR82G/8uFnB4ux+8KDmXyrgn90KYSlEhW28IdID5NEwqI4bbHDw6QdqpcHS0
+hFCHzo0JTRTUsXaarWvpNlvg7JgEZHmT6JIommCVyu+UDDadDEIYarvr468DWIu
F1FFGLklm/mrQzN3E6YkF7DpJuHwEXI+9JepQw5+scOmqyGqYY1DarUaKkF+ewkC
QOCGq/8dRQ3JEwLCEOjol1LejlzCJ8lnVa14k5onANW/xabK8Cnz+CxCIcUwP3bp
fdsE9Mn3qiM7S20cdRbNT1rAEDg/d/Gvq5SI0ik6MF0BgyEVCOy3SUDJO7p+pf4D
n1XSJyqoVuv/qi54DK28TCGtlZ2x79/Mj/KGJdX1BUGjhENNeaiGUatdMduA8J9I
tsSkzGNziDgXSwNhTZDVX/SdNx36XBFC8YzYnIP7HAN0L0WLmtTs0BKWih23mEW/
wxa/j84yxmqQoUAgNdr3GayueZ8OfRxbcBH4Jx0g+27UIzDGSz0YE1WPw8oJeWd4
UZvrekQXcBS8I07H24m0iUoJVPBdmIdvnDlQybpk4ex61LhCOQXDziVMgpjS5D+W
29yPQib1E8vVRdrXBn0FxZCWBcnTcAViYibBwB7QGbinRZsX9T+fYUySKZ5BAAI5
KuP1OSTEV46bM0V46S4DomFYA71d0/IlVyTxTkeE0rDYcgCFWsnhgKss82T2a7e0
0W3UhcQArxF4l+XlTx+/pNtd55wOfF7HZ9LezlNTvF548FmQPFXkqjERd3ru9LtQ
CYl+PDb+ZT7dzbMlC0SvP4ZEw870Cu4VR86v1G7/vPg9+A4JMLRIHoXMI6FcDATf
uucOkt3Ufh9OuJ8FBxpb/Nds8+1D9Ny9b3eJ0A6EOZ5L17brX4ovSBkf5gxWa70b
9+Z+Hfiv1ZVXtMpCMeu2X8Dp1gPuVTQq6qeLjnIWcwql8n7uoFYB1m0fgOlH/CO8
Vg3EGk+jCDWylpMahTISh+puV8/zPIXhc6DYlD3N1hZeOTWm863HCXCTtr8Siy6c
nZCbjxtjJa/Q6tqGhtvz/2CphdQJCkF7Vy0ZEk7i0VfBb79qyn8ZW5pFLbQUdLQZ
g6Hbud8h6BBV0xsdysZEOZxdvvDy9wdBofYmuHLR/s4iuwePDRqa3wQVjNpyzESX
8mYlKq1jxR/HyJFec3IYSost6ZOr20RvNtQg2FhcDLBLTSNlrN29G0QX0/3zyAP5
L+xd1IGtCkloNcYz+uciG7+2u6AQxWznzSmozVt3LacGTW9Xg0IXmOTl6n3jkSDQ
E5IJxLoNkbNGNy2trB/eO+E/yG5PGenuNoAn4BJLDGitnQrn+tmaBPk45RATGNqW
FX8i7AGjDNIbnvBehC0MAx8A7ZX6MQl46osInS+4mbG8TAmnb+eCq1uZAc4YCqPS
bIwCT1U5sFr2IiwjQwwaN7U8c8AhbnBJXcmEokeB3gaJlbDYUHYCh5I00wIH5BWQ
rTcXjem8yBq6VJaI0jbbM7BgCDyB7Lk8Fwq6ScN+raDEZEG16c8HCxGABwB9u+z0
YoOqAC48Pxwvn1Hqe1/3lLKlVovf25xQ+T/v7zLm37o5Fwmt/OrQ/P7jNkiCtkai
NCAV9ueSCXxnc5ZhUYogH2Pw1yjXPshvbmYTmDISAsnmGVX2Yyj1NTfpnaP1KUuX
yVIlzkyRynfWaazBLQRlPp50du/pzWu9Da0OL2vE8dwaNyEteSRmlgHawUfJfElj
d3dvmc6flw7M0gkOZwfU4ejUZ0REZhMxPnZmq9LDQqNslogGWjgTnJmeUeYuSO5O
pIMtgFCzfsDLGS1ICtiC8z85Xfc3ywRxPhai7aOKLudXzTWDPWW300tSTqWBVBtB
2HDSjhfwGTw1MnRjVMoAOrGClWjK09c2eXyt7eJpTD714VCbOI1WQi0UxocHCM96
2eHZJAG1HivlEvbmns8Ot4IPJidfzZC7DxwwPqrpaWCyw/fkNpwwaAShQpWNrG6R
7Rytd2AJY8E4RuA1E5zI2bPryzsTsEWf8IE44Lot8T1/NEwTsFzszdXWS9n5f9ua
dBo1kRnXk7B/XG0fFgY7pcg6lLGL3x0FOHzPE0UrMxGz1rmAXrc+zEYTI0omWPfQ
BAoHi8a3AKd11yiAyYszwwqst7AwitpHb0uPEhPmYydrr2qh+VyIiz5EGHb/eryU
9LvUS7fIyV1ZNMXb7afdhlMjbZE74uAXHc/S+j2PYaWt6XB+pBjqAphrODKYaB6E
9aJfo/0ol6VFvFyiKBR/34t9BFLSmqRZel24/lY3+xDP34xXANOfAT+kh6YzhmtS
4QmilhNGfd2RotP2oVg+WWCBQhphxDCZubo0cIThDfbAbr9BPCwF5pZ2hqSHZ0i2
iJIsf7SddSLGjzI6RTO7GSZYiiVEURI2Fy4nAG5eICR+ZvVvh6ZNDK6SbXEwl9Ob
lkqbEIzHDuNa2ADpTdiuNd8vh6DrK9PX0CfgO1AKWt2AMaay7izNRdr7dbyoF7Lj
Rpfung1JuLsQbu0cP5kUmnKkyfWQdGuwbIOGmNBYtd7BKCJnbxDkz6+KZ3Bzl5Os
ZL48/vMk10D3/qaS7lPcfTJBdcdPaRihtJct0RHcaiVKZLANrz1KgjtcsPE+sGb0
uiVV+SoChPB1yoblBxZa5mEoZNEfoLCYua8UuyOvdZ3pvFk7gLtmZ4H0GQqiteb3
TM8/bf6RyVc8MsNzKVUUa57TMUg+0PWiY+TrAkfuDd/ZBD+5mSfB1DL4xdLcMsgl
WJiIpCfC2wWwJjElqaiWG6ytv4x4CzTBxTCW2SeN5jrfHZDVdYdLI9yc9Vej/MHn
S4kljnqgTJd1Te1gtQAFZYwbiwQD4+3sZ8KYX7cS7y9Hxia1z59HS/B7/Nmz2Cje
hSXDIFRzpTzusM/fehrrElAc0byXkgboIVHVHGlNlzfJC1YuG81hENEQKuYlwIru
XlC94y6X5VQmtSiWH1L+EXgwYmGrZSiq7HvvzWGbvVFV3PNT+BaJi2TGsEaRfwH6
SegPtSOinADQAgRPy19vtnaVADoHBs1o3Zjnwb3ermPCfIAh9GeajBgLIJQvKK7+
pz7zBY8xTyj2BQT44FdfAieKGkHaZzIKtGTupMiUNFCx+2YuO45X5LTDFyF+4g8l
c4IyzjhDzZtG4nj78HeBNvduOOSZwfh6uOxqlMr3NKn08sDaub10UXq2AnjInf9b
5Pbe8gTV/esCI4YPbtHTt5+btOSJuRGLrnZ3wqSDrgcAwYqOKdPvJMUfrP0Hqs6T
gyWx426qmd92mzzuHau5JfCxf3aT/ShnCNvnCiuDKnYA4fNf7olQmitzVPzg19qV
fNwzzJJRJZpizN917YV9BmcLDS9vdhRk/HnwPJG45SRWecljPGiCG4OJ8bMkv403
laBsHiIBHt+gj0od7tpjFW6B/KTbwo6y7MeRPU54vKJCLuU2uMvlsdof2+sH1gr7
38MTIAQ5YilDJ/VKnwdC9Wo2tUNzBcsAfAarEMZ/f2Vh+XImIM+5f6ghfhgPT0YJ
wpzsSqb9XNWzDJkjagLaKQddbjb26okXJ3jhMQ2cocC2eBY5YUBg+DJQ466++4h+
lNnzSAoxdajcjQYWLNZYtxdWZA9V86xbWTswVTodfZH3Q+HL/FEDxAeDuP2HyLlM
8mJPwolRToNHgkoGwu62uhazsfZb9X3oqA92D3tHY2XX6yj9RGTTQQCTTtvMxxs0
r123zzV3IFRWmVpieOecoyEaBkvmFoET3bVTDQP/QoYgIFm1mDSxY9Cpb7jdoADv
jILAc2gR20y5mzo7ULYx5p1m0TDpzjHpSkXiuPr2xt3uq7ZrqdhVZ0X0j95P8wSD
Mfk85l1bogdmfWXxJGZkB5piuWbMh13V2KPHLJu9IlmVnIAp15/Qzvo1l7QqPlzr
V/8kIGf1DFizxUILIrhpctK6uLhBSN8UJWVey6YMRJaF8ubHML/BCKHT5+MzP6An
FRM8XZLS6DrF6ZjGiC3G3WpESLJ91LX5H7Vsxho4jZiaZ9oo0623y9Y87J5xGT4k
HiASsxsauEjkSyQh6S5TF3ENe8evUC1IIqVJMtLOgKiok3e0Yer9DNEv90C0wTWR
jW44xXY0SAu7lhRqH+CN0haoN2Gx54upYk78Taf6ZMoniEtuRD3n7/++8WdAKHi0
FCIl7cdKU9E2ARv/mn/NnEzx7dBvuvP+FnAJi8StHFxHZeU/6XiEworWYl3kMKId
+Px2s1BaKO6meZg+UL1ABNCneMhDNmrYLqF3YbOEOBm+JuPLHnlxOMNd+Smr5Eyt
COBF/VC0z8Aj4q0lSezHUOxb8Lk1kZ+VfvwK21WksX0AfCC3gu6rZqnGI/4zAmKV
k7Wgg3h3kv9W8xcsu49HRJsLrVRkTka23HhA9lJmZf0oJYdOGwHK/latTFSQsxJt
QaCjCqcyGu2vKFFcaXiVaJzyKwfCO7wVtNKYWOia/oyH7Y4Bq8j5nVdc2gie+t5r
PjxsD3u3GjBm8giiQ5Rkrib08nuWSlTw+J4cNGTXHJCrz4BZl8S1OssWoOfsrfzK
PaYgJ0swdB2PpV9jP2hIPSTozUN9hM29T0pf9cNaPBdMZ49JwrqupItlA8d+FnPI
C98f2rmjuUGh5qNWEt1yyK+b0NVjstNnRMzKTKYQ0XSDNptCp2e+gi5vb6mWtQdS
t32jD79qQ4be4Hi8KtMV/wXjNb0Ucv5gyeiD1hCjBgKOGHiJ/jlXbVlLGvpqEZSd
oUntignJWzv4mJ63jHyp0xMnvIandHGL6n+Oje4ALOLy2IEzBYwSSoB11opUysBi
Ra9QBp2Iz2CVuswGkwy+sK9F5k4c3lySs3uJI9yQY4AsvlwbdMnWSmXCKbP7NBqs
sF6A6sZfz0gKR/yEVdrzK1m0b5PphYcUlk8T9Ekp7TRB0R7Op5U7w8+H/CCRJp5z
OssgwzDiLGw9DWRk/tZ+VO++8ugefdhP0VPQWnP2/5Ydp/kImgHKgfyxp+c9FLlV
Rq9Rlrs5jIqFb1AfKSsPLiwC/NaFzUPOgRuBh+Crqo4J9BYY50Uiq40zummlotiH
M+D26YW4kGyDV812+HT2wkEnuRWlHODfF38rtsx6iF3pQP++IjM0bcrRiFyw7dU2
fx6dFhW4+av6YDO+70Ls7sJ6sin3ZPVoP/vRDpjJ3gHhOwF+AVK5OeMfehzcakBw
Efxv1Uxbw0a4nayXHtov4Kd8nVZmTCVQCbmYK204IXNuVy5lRhe2e4QATpnL+Odw
8aoRIPBLWjBjikjrDnwNt5Pq2gGmga4hAtyd3RGD2AE/f07s0jVqVAksJIS4Uqze
kQBDH6F2mnQpU6+WrqxpW0MwAu93GLVdpdqeduIR4meEJ/ctqR6YZOBI6T/el9bV
9Xj5z6Dl792/EPVqmD1whN11fdZ+Np9kgFcQZ8ou222pY19jDTpFm6gosEOqyULJ
1bJZsio1RUPV9ZPMN9tjJJs9yeJGkbCyFetPVCcsG/Mu4z1O/yq/M3CI90rL+Ci7
VrtlZJZQoGX950r3iFiKIkyZxM5hzjPYg73O4Zd58bgeNpuG8NfyHnIJf+A2oVms
WEp2S0fx8I5H3sbN+D1isxtas+AqDkOhcD0nhZZGvgqe9Ck5BPBrBA6lBoBFy2el
yggA3gCcMTFL/CDvwVu9ED1yAmRXRkgcPUr2dtX7OiA5huuTLW1EzW+m3Q5/4VWJ
WIL5nJdoBLmQsDS5/kRZJRG4G0B1VevFmx1qPCDmN5k22NHHz0PLJ98oYrutkd1Y
uIel7YWMzA6jRoxP2tC1mVA+m1Xn+PFsI/yeHgLfF8vwkGqzkoStO1D51VnjQfla
5UfdxM5VIcrd1tKG9PgG+KGcEwXrtEZvf6thEY+43acsieVm17aK3MQgHX/uADHZ
31IQjPic16On6hhPhcYWwFt03tqdxzS8EuJBxe3LObApltAvusaLER60VummKUCz
mTZtiIkdtsobcG111G8p2dmhqhj1Tio+OWapYLuXDBFSMrHEFGODTXgBKO3rkDr2
d9MEOMfNQWizTvA6EHKeSg5I0nWrL8ztUNyALNGNz0qnp4OGNRw0cI5THkuaLbuF
BmX3J4yhaO3cpTihRQCm4S6ucnqZtLkELLHwY7PCPdwOPscxBlaaieYx70GqZ2iG
heeHjIag976HpkAoCRXz1HvjnOnojgaAjuPkp8GsTjsZIT+6HD1OGHgZnRyhp5/K
ViuMPVRR6eT2SH9zWx7XiiMu5aZ8upHhVIR0y36xVc/FPUp1biRimUHQBAzbGkR4
M2zA3wkR8b7eEox0AsurLMkIQ8B3fuRxA+fSwKWT5HWTNCHqAWDhCI+sDNu39oUA
zkz+LhughOwifCCjs45EGzNZ5MiZU+2km6ebG28bgsy5BBfVWEH4opPj9bVC2Nds
D13UUhTmar4yWBEDlve3iPX24u/xc2DE2r0AaFvGcl2eXTKxHK2BKbNWiHt+jV7h
iwXB2SNmDMNq1v9zjphGRTF87BPwC/0ODFm1xuvs0y9DQ+/e4OJQt94Hw80Xg5Te
WozSGpDrWCaB/Wrp8eYIsNaYDJLO5mm8MD3KoxNSPb7SwVmeggPgIiZxUrnAmQjf
/cRxnxMrr3qd9IbMKJv7cYcHFY3YvGGbEpRaqtwca5ncmyhXrA+7ex+hlZmoKgMB
mddp01UPL7YVJ8eeB6YYJ9bRkYjTWpjuNfVvO99248ufJS86LpSTUi4lb4q6qliC
K01OgvViFjiqPvvVIOT6JLi24d3RZlk0z6Bevcyukfy0WTFeK0kBiOUhzI9WPzy8
sdSGOLpX+nj7/PznMXNEDuDUX8TantFPMICapwD0+J763klxiYkvLPxfnz6AqPf6
u1Nx4f5kW9eMq1FB/Rc4u/zcPgw2IdsrehhDWhs0o20VxaolFDrSCDYFoTZQWFg+
DQUv8gh9I1TF2rblYMh2IvF44XV0jjl8lop1ul/LNBPwNllKgnXLPXbaJzNaidR/
5cD3APqz23rxDwM5vUNS/Ke3r7jucUwN7ghAqNLf8JW2PtcBYJtUq69IMd2cezeP
sVdSPbC60wI2yNulicJJeglS+mheiE9Z7Fmzr+lIxCZc5whBb+BqbfS6Xx8cZy+J
6P7Hb8j9EogzqpmYToOuOxwyghFzFPHdoG2Z9yLYfNHzi3kS1p6c6ai0IW3sxwbd
Pk8JJDhdTvRthNCvCjvcZzdBL3nSCvRZvj1n3nAzqH97GRDq6/qbWEF7ldfWrDOU
gXOPhdw9+Px68Q0aWxofxARyizyDgD0LP72nsersw7zmn0oT4yjX51OPOe7Pivto
YyUWLRBTi9xFwl5qFbC00b7wOoSx5h01UNbxNFibscLfbAsX9mHrHXNYC1N0OWEy
bH8eKD2Y5lrHxdJFBmZ8aoaEQglAzVnhNHkk/AdfyfXVu8BTsw63MWj33WZEqRHX
bob71dfn8AaEfxchW2Lp6MdxpVP+gX2LoMeUJgMH99BolaiHS19mJ3CItUsjGnG0
IlJz/GZgocNFOugBQZA+DwHiftyGUxtsQfZWokebHkTRC0bDsAgT7d+MoHcEucc6
3KSGqBU+mfh60+Cr3Fjs2il9LRaLScqYvmvEiw1BGH47x6YJVFi9BLwhUj5vWzO4
a50FKyCX4Yc4a5KTqjv+gEHCwd7IPYs4hiTvY6vk09OpYnLGtoAM4+NDm43ig/uG
PMhHdXktjqcMwPlZAR2ZF8BNLmnW2dwogIfAWFvJnOjTIcI7TEjL7oPR5TjvRRLJ
rNXFlf9BbDVotqNkGP60tIvuequ5hSO7fOBW1h+Ur+XtA/7s1hdS6r739pSG+ifS
1tIGhvTS5d09FhNf0w1XXtPQEisgh7ViZ2PNi+Zhy+MbqCZfFW7WhYiueEzGBC/H
PVkiigngCqQP8Lafk6nTLNKg1px7StpQQvbsvpaqZlCYrZ+i04i6QKzV2LpUeR65
dSXR1uv8OtrfF/s/CQpats+ndY0smP0jt+ZaBpg6VtepsR56/+wIlqHuMfGrAfow
8ZchpkJcTMuuBu/jxzgER3TnlypFkv4C4V1dRxHf5WWoLszLNZWl5QMbjdH6x5vW
EQg+l+HQElZWWCvJ5X+O7vQ7TJF1ap4fAGpTeSxGFNTg5hx9UJgwxrWS4qFKmRV/
iUwVhFJ6JfODh4qzfeUfDRA/OCgC5VHnUBX+pLM9l/VGToVR+0u1KLbwHm1KWcXz
qPn8jQpkPB7twUmLGRkxowCwWeMTahUsQy3znTtvrwLGYnMXIEd6R7vurjvmnxRu
t+2vNqHwYr5e5cNiRpWOoahDi/UI+Qu/2F9xoa5Sk/xvQ/bebiEcO3I7p7pQ3Cp5
nyKUQ2/uHz3ru6BL6DfkmsItsdnw86kWN5MoXD/8BFRu9yhYu/+6//GBs8g0FPla
u8eVu0VRADeIumMO2gtu7by5ADvS0MBgVh96XbzYC9j/ekL8CO1rvV8H2Lx421g6
9jP2qCM/biqdHOQCjWI3EC9P/up/AIKjbORabImkJf8x+FpGidIoLMtAcqu0/mAh
pNPJIBYYDcKpbA58CgqUhOl7W9QAPbnsZF29EpBnWbcxunVONDto7G7PDdGzJSGl
UfyB/fRcIdCAaUlKajhcUOg5Y7MASvtHqqA4NEEVW2uL9uUprHreJNHNQYbW77xT
B7agX6tshva1ySBSbQbGrVfDN1ZcfatixVKqejG/ZDqLXjh9D6Bv7jKrrTDPyBCj
Lnn/cUUmi64BjxAVTgrolZSM3XBD/LWQlmfd7AhEJy0ID3mcz/cNdgtpwf4jrjGp
IXb+ERW++YiBGAStU9wOU62e/n1s40zY+nYMLIjeu1LdSVQD6Gi+NrxhGYSNPQcV
dt8L+6Oznz0YoX0AgJaotApfIY0xxgIXHj9SfRMa+jkbRdMdKhzIgJ19RD8sIjGO
6lQ+AnMCM5RbGF8vOmhm6Th6U95W820YxmNJjZS/HeDWpdVL8lKkBr6rW+3uRwfG
XoJu8/98i3RNBqq8fIh9RXqNEe40jKkGAlpaLdeyoRkKYK0Y7rtZbx7orHM0AjDk
waI0BXBj3YmX/Mrz86JBczYS7T4Sptpnx9VPnZN/KiXqRIlH6gvLMyFHa5EQrwF5
TjWAB+BmgjVsaCVWoUF0dPRjs5aX2x6USeNdUe8kltYuRa/mURkP1Fut7AwuOBk2
eYKqeL4ojYXNY6ZGaEXb7a49kIT1bkO/+aszLBzPVNX2bwG9amk3Zbas2fA90eXR
GQMez86fNv89FRir4Y0SQYlECtA3TJyu57D18xP2vEIl7KCMwF7gVLM9YJrdlMUQ
9UiKNJj6Xb9Ucvb4oHiNsD5fRTpQsFO3FHdu7Qk83Od9x4fs2rOPRSZjf5DqkekR
EWqgUGrgYlQdTZqZtm2MfXyn/A2COHjSZu6B+r0/6OGbSTXDkJAKypRDf4Hy7gDX
7d7R+vv9VmDNstUFFJnUkLDiRPX3Xizv96oYsjoSlV6qPN8FuChF7Y5ha/qvo8bV
lKn+oAU+Gl9VGSn8N/MDf5zeKUjP02jSG804Qidz915Fs95Lv3uWSrTA23KGqBDz
wm9PSzzstdi7z3hKOUDGWfvuQZoQnpW9R7MofOwdDP4cP2asjlVb8ByMufqqpAzO
zrqjmoLnSVUbwXwr6IMsgBPSq5RS/vd8v4ZP+nbOVEspbkIwkMn1FBoNjoWruonp
SSkRcRzZElb6YDlzkC1FeLHTEv6U1JgWolQNZg9xgMBU+EaR7WqMi5wGCF/wH2pi
B+sg8bmTOe1Ydm038zAUwBybuOi5gXfta5unsbzKmkitYJuAUOF2DGxNh4Yp/G0R
HoF8Cg9D2L1rdsv27wkHOndkHr6pFlux7UWsushHlkaxSAwa6sRHYZ7BlKkYLU/2
Cu+/vHs8Vn8D2DYVRCoUSCM/9YfRtWjZwu+snQBdDfKeNAfGwHIxL1XpWroH5gq4
jKLCFVzm05zsG/RNyJH88ze7TVboJwIz7TgvU7Bxiz1Sz8d4pa1RcOzYI38Yb2DO
+JGBcC7KCWfjFAd70w9IH7/mAkEO945n/fUoP47bjckt+KtLDY/NPC0dY5wt/RK7
cP1Z3+U07kXBEqlLCT8tBBqjcN0B0r7O+CNWHLpkZS8R7uqItUe9wIAyNbvHm7Tk
mdv0h+3CEge4gLcKNODJCkoJ0mUQQ9Eh1t29KLyaTsZ9b2woJ5G0ZMT9OyYroBOd
HC3bMos56p3cujAYnzpHI/3XLZ1EHcaosZfuhbLrTbaeqP9hyRiPKAlDSPsIhId0
vZjrYFTLefXYzGbI3OscqU3Yqms/3LqwyYWG1rd07M3jIZ0oZ4syqMT6gzrWeHBz
TN8RJqSRuboVtP4XpC6BA8XinIx+LjPKdsajSaBFdwAbbXj8SwjE2g6gRGE+aEK4
UTsvNdJNX+9g9EUtRrUVnaAOHf2noJ20QbU19m5F9zWSsUp4zCM/kp09Od+5bl2A
cJKjGKq8U9aY9AD8gg67jFTlnXcv2TZL1M7QeAudnpWSQZWKk7QqFPSYK1dXJLkR
mIPknYg/+bKYpAT0yYK/7s+ZpK77dZDZNfxdHsc7Gj03KxQGTO1T9VnOJsATgUJE
2UTqxDkZD/VKlSlJ0hcYlwDe0LLBweaZdGIehex9Ism9nV+c2Bd446UNUQN2+7Ow
USdsrhKJSI1Y/WfKSMxEa4E3KODqWwiJRu6LmHtr/BlGVz2UiWXuvWDGiR/dE38P
mlo2qtLlRXQ6hzzaCaDszPkCSGQBneXkM6XmcrOznWqA6F/km0nOlJIkJYdBZEPK
Q/h+JK1R+uAECqosWM/+Cllj2b9C8JFhYaOLRrvY0W+UkeV6Ovo66iwg5vymwuSR
/ugcVdsZc3NX43IOfvlu4GYLoW0Fil+C1mml3ixbdUoO3cAithHVHbOv17g/Qz2E
p8yfFbawXpJ6379a9rbH6iWkeY8Sw9/4RUcWgec6SqGIxJbAKUIbApVzLPnAxoH2
dkPI3eOlK8pQ06Owoa+sf3Iik0QIS8PGMibT8dHQimwj1/gvRpsgGU6q2qn8t07F
TGjPRqfmM8NCI5+DvMgKUwQ5SdKoxUC/7eE+dqOiMVMEz2Aj6/Irdxud5gfa6oS7
PAG/yRv3pp+OynHLWJ4YbFEGLuAVBk2cfogYDZYw2wNYHlE1jSD3cs8MJenQ8a5u
9Xz/JbRMxuMPuda9sqlUW8BML/g2TwnSS3oMRljPbZ7bvqDmXtMNUN9MxKZT+du0
+gletIMV8djVFEYKUrOT8Zn6wAqjKcnbqgmBiIouBcskg9aajpnNtHU/E/OV3my5
CC7+Ev+xSrzqojk+6uJjJuYim325sYT3bKnQg7p3GvKxcrAaW4jNk7JDhS6tXspO
FgK5cpoamxW4iBqzSsXX/MR3CjhG7qOEpS4GJ+uOdeYzFW5AgAnytjDQMsYOStJH
jJg0FlCi/EmSJ0owPeHcPUdJyNvvliXmveHsFBV8314HXqXqm1C4/w9a+FoYymc7
OclVOtpnyAyObGYq9N8dBtEH7q/PybxB8oHVthLv4LIV+wnmZFa2Y/MCuIB7hgp7
2pQ+6y5C2QcjkGOeQ6S1Ljr8Yi5ssUYaZg3TfQWQpWALuKgWteHhCS7seBzWLquD
nPPIqYNEzy49V6rI8iR4yEP1DNBKzdzI5Y7YQBNK1NVokjXkbDJuWEuDC0ivdjBW
Nx1r/N6aGETk+jMSa/B8vaenRjpY+9P8QJS41wZQvP4TlnU4Zoks1S7y6bSX7VKc
pBTuzaysazxmWL6T2H+Jv4eIpH66qO8dV79OVH8VkoqKSEcoY7L3LxzWPm9BfRHl
dW79NadXMDilAEa4bVH7WESpC7q4EOuJ7Px4uON1IOt53l5NPmFY5F3QlnM+oYhB
0ixdohT/WYLb+x8PzWkIEyeAzFGco+DuXVzcNi3/BpjFKWUIDxi/lAFCx42DSpKQ
YAyAGBqGO0HZ4A9L7jeRrQ883+Zv8zwvAfhrQmU4QEUSeLYJnTafy9DslaUHv1bw
odpK7SPvGGgyo6NLVMsJtiGWGYZB/joez399EXyKA9eaU2VetktbpU355nP6YLiW
1Z+amox6GSfYx5AtZRagQcCibopCmy3AtiTJcqk39Jc9ZVKpBpmeeOuN8TGlwJWL
+m0UokUi8c8HNZC03HlaMtrbwTdp19Y0caAV+kpwDIpGhvcAnXchQl/rveHIx7e7
dos07YThqTtjNkj3KhPblPkHph4NcEOC27KOSSLTzLHwNGikNXnRwOrL0KKFe6xb
TuWCalOx7d0JWoNgMEpCztmhdGCmahaS5kXszysyvh49kCxIzyLxbC4Y5VGpYOYR
KnPPfPJ6sOM5f/wJcow3ua0jpj3endmDRucFu/jb2YDM9QgXQtqkFpgTRAb1b9YX
Xwq/q9gJjZDIdlAQObqlBOlJhtXTBxcHT/C0nwO8pwiNxoqKssbyuFmxPRLFJ5nr
QT+jnzRhw592XbTrGD7BJBMNl7/DHsSAAfXTl8xzbtSGblogMCQ7AaskJSb4Q61R
oUllczu2NOfdC4HhKuzvhhHsVLLYuVLJkXC0rKuXORV106xsPRhaIZPELtyd0Xcf
MFXj3iW/YyxY9hhjebqje2f77xUanhQCcGemUjkmfyBWJGmPuKYnSmQO0ee6WMKZ
t5uV/JPY0Ky0kFedtmFUGOvbxau+tezflza6xmOEWmo2V2rKPF2axS+ip4OaDhsG
y0xREvxd5Avs2AgMZ6XY3mdSAEuodKBM41HSI9owyKmSBMH6UbE06pwmmpLKr6vp
RYOfGPwe7Y9yYnDUiD+SosllDBgJwnEoCVHUUdLzQRQQ59CMZGEt2igqP5VDj7uO
JMVipbjRM7LThru8JvKoPQCUmSrFJ2/VrvrlwZLaw+xYZtx2ugoESCTMOvRdsghY
m5FmCgZ8Lu+/HyBYRH+XD34Ui+pIhf/i2ounqtRnbmERr8uraji3t+w1+TaV6xrf
oBkL6rA0K8Wjk3pydZhmijymvl7KeAkNxJWqTffaowTKYamUTr65uO4DMrsz3r58
NKybIger0TODqEn82XGHw3cFzeE8ozEu6ILXzDyfIfkPx+8QWbmnqnjQvTv6vqCA
k/CPM2wi81QgCNMv6IE8A3+29WAqk5r9f0hbrdoXkGPW9KMYD9bxhM7s6PVGEp7F
g5ddqluSNqKtw1mAFjoKFKFFTnRikDIZ+4C5fYraRhpsf2Bj5766akIzBsTSwc9x
4Yko6OkDHSpwd1g5/8O8fBfKl4/vZCQZMzxzM3ZHGpXsPfAXPnu9R9XUwlyIvy13
S5ecskIfTbzuT4Q8GlNCSGIaDGSwXLQZmofyhzCShdf7Ozzpqd4GfIqe3klNYTnH
ZeNU6XI1OUkyV7pNOf4Vi2dHruqbsOPehIkwQRyVAyVFGbTMQt1NOR9sisbYfeKF
5ruyRY3KL/vlFSl7zGKNEvuVacT5AM0MrvVcsSr30lK8FEObx8jCxZgN/UNQOTmh
zKELBHqOLQgJk47Zt9ibz/EGqcgiluMWyKJwOM3YlNnEmVu1OnRktqP445dDR+dS
6gwDUYEkzl340SxNlKTwc7txYomziOZcBPQ1uw7JwurSKseGmMaym17blno1Coa4
TkHCnVL1gfD0GTNC+moNNkWUYHjjYwSVMMz0zPVeH2o8FlhswH13MiQA3ZwFQfJL
ZB2jYA0QjU+i6BVRVF1krcTW8mse5HkBkw/fJI0vHI87/AiCSutzGp9vmasCmEl2
35l6dle+Wi7CW7EerJAVttnem5yeNB93Zg6ATCFtf33fmP250M2+jiH1fQbcio67
CKOytGMAD4XjfusN89YbLoL4zbq5Iv87gH43GOFqyYJD7RCtuazBfDYkaQBp8Yri
HZjtdgrwSmnRPLIFEScYCJ9UnmaYQtA/5Tz/n1ZEbMfQ7DqbuJaBaV6DRVBM75VT
WUktPMjkaHV7gqJghaBtHd+61HkQzvQpcksQdon6oA3VBjiqeUOdRJO2x+Rrsfzp
2ImZXNFBBm3bziG5Ra50/erdzYalC8AeCyejmclQNknphD/bJoSiH27oICnSUbld
qzHEI2Sz5Sl5ebYxrs2RJWJjyiHMZkGoQ0XgFda7ADHxzcHGrML3VhEkcj6fKCQT
vVur+NJtd4kQcP+TbK2OSspksSMo8rWzM4TmFKx7wAWEC5WG8SdDFHUukrqGNE2V
6R9LdZTU97Gp5L8RxDs2Fso7MgEHUS+ETXPxUSWkBso3of/qZdKWB9YB76WZeyQm
HBKRIGAtq8PT5/NDOqEKH3kFsUo6K7H7PiHcWtlo8grNpAVCZljz8vem0/7AfrPL
Cs8ruyENc5/jWtyn845tB7zsWnAS0s/wUO25t8UJNLwzFhz5WUnX1gT8mSBRd97S
wlgCZ/HVZKI4aRDgyhpPA6Tfs1Nbbp5WMnYoeF4uMzLCgmW29YiB3+AxRh1+FClw
20PjNb99sbrODr2SKnl9QmWsr3ArDMwc8Zh1KCnaAITvH3sm5KynBxEjDjfs77kn
5rOb4wo7qmFP/sl7Ps6c/f+ZCgVnh9hZZoq/c7KRJJ61+Gy9f0qe8NoXGB8oogLd
RwDIddjy0FSKGIDKDm/4hryFBnnBVzJTVzeHtxXtOsFX+G0OW9oZtLO+m2mkaRFi
4YSRNmsTeeA8lmc8bOpEbTtDbEJsGZO1V5Y9NYxb0WNSsV1DMefB/Yxl+Lcxsuyu
1/G1I8Cg9MvgNUpYYBS06xkwZIG/rgmufKfwcyWe0ihqX/be3ddso8r5x725ZTbp
9koKUlML9xYMmTdkHHhOWQrpvme2Y2NjldOqzBvC3z08whGjshdZ2AtFEEPpyd3o
/9CQ3+1aua80H8RMXSocJFa7xAFoM00KF0ZS2TeIoYFtYNnvTwgy1kwZ2bCk1XcO
yfDRLwd/lgePvy7FriBaR24r9AcgmuUBGN7PZDcuVcWsh2CSbVntGGStUZWI07GN
Udmnx+KZP6EfuLWZ1FeD5eWB9syc4A5Ndd4IrVOA7LiFjyQSOrlPfoh6EAG0Mc7g
gGEcy7JR44VFuE6k7o3/DOTT5lqeQSxTfM4hgM0IPsAfkM2xRH7/vPLRpl7Ixu0y
sbUVHV0YvpBG0mqlHpHsvdr4XOlvz2sii02SFdsQpjYC7a/oeeMUc0u3H2Cn9UXj
RtywknCar2zg+lPaS4NvVU3OnIYdvxMWsTdv6tca7IbP3t87EtHGXY2voXYDoera
n5VxmsfQ2EUWxk2AcyI/aM3lNJdOA3JBpV0B0RoNZt0BjhQAfh0O49EsZbxFjARH
tDDbGL46F8MKVl1XeOlZZvVCzJsJSjnsckIdg0D9LRXU+vTYNKt/8MBkyB9zB2i7
myA0hSX+Z33VsG0ne2onwndJ5nfKVNvVO9Cp12IAIJyJwoyjfPlS6qIQsKJiBi2k
oYAnlQQ8nGbGjj60wZ02mJBEDrgTlJWNyWpPObIuvLVrzLtogyysZAQaQD+UFpcw
QnAJxCGV2476ztRhRhE0ziWwLBK6PZcEcvn4Hs2jtWPorqabMcQFhRF5b/B2opTb
Oo38QZBq2IRHMmBxYJzKpDYseNqbCnI7H4btHvf+cXN/gS+U5/VAiurfYAPe1sNL
IwwjAjXU9Yt7Y0opYZeIdolhOGTQtr67FbqRM5bN+Ye3t4A9R/JaA+5GtRxcDSjf
qcH1Bdc95fDQl0JfHIFb9SRGDew9dLsuWAsCrQfs/3uXH+TMp0qpBUtU7Eb0OTdE
2TVDZrl4Y+V2j6bN/lVHp1axB7TZrii3XX8v2/u21y3EteM1oEnIuNLzgOsuWhAw
3jdb33rwUIBb4q51C6s/tkxEr/2f1g6DA5fIrXLaErg5NQW5LmHSvuIF/NJet7/h
CP5Fy2LtrwpfDa9+ZLK7Rja0Qkczht2MmxrUHSE4FrBdzpW8fuqX67BgyfOnuRh/
/NbmMGlCPNBr+IvxgPkfER27bPLyq6VODA9i/Du/hzqpFU70EsbSF91epe/5ui48
tjfZa11isEZ9MA479wEtdwvFWkq732yHFiH5ANFed0F4b+x6i6FlmLEu1ueuUEAT
gFBCq99sChgNAQBTBqovdadaEX69FaofTukWXiBQODRQ+FJerHzpi790d/3Ojhqi
pQzPL9ES3y69sRjXzoihO/hpbgUfozHOpgG62pgnF1ql+HYyKlEB3CTxiMst7/82
iIf91J6mWkhFb9WraUDRpvLG3rW1F3k8dxaUakoS6fHtIbpqTRdpkOmb4m4GxQSj
yCidKVNaBlTKiktp+gs3uKGuJolNcZqlCNb0zbVKvP7OMCxmBVRAiEgTM6djrpif
+jhV2KtzN1+P5yHciIwm3e6upsPQ8gt9AIeqv4MfCI8u0BJiCwcO1/SRAMJt5EL2
9gOuaG8N9MJP7VYZdZUs/BiK6Zbph8j9i3WWq6m6dsb5R25OJv0tomzTV+m2yFbX
mBrDE7KbP2y+RB2177wn+sq+3xOP2krdp8/ppsf2PZ7CiXPFXnv69R5XhtZtXIJ3
K32h8vd6+OeEwwr84ehVc5hqHbiF2WOKyLkSxwE1dYAe8DHgXiv2sSybg/DG9Dgh
GR6GGSWKxWGuwz+d8DAKPVWIAJ+OpGzL6JZfjVStQHepWYSm1idI0mWdYaaA9Dsd
EasEjVSCCUcuXHynNcbLC4J6XQzfai5pbbdnBBSJezc3DCkbw2ERdAdSpkK19g+I
Q+p3tZpcKfZZCBHgRGvgHhn3RPbNlepwiCfFmWAnwle9QEw86n3P02pA0Q4jWIP6
zq6Y3Z2DjZWZLlcnTHTMO/eZ1AX0lYSzIz8njKzfeY7RmT5m1l0eQ/G4ctlEGSzX
+exZdDt19DdqOBVMwbGhyGnSnw7R23dVXRwz6rU5E3F0FE36ZToRrNdsFAOtIfBF
jYErbOLOZyx+l2PTZRfB5N4nWTO/vowyJ62NK5Ie0a6TGVR9NCs9Mi5XxyWZWFVG
MFafsmZOLytaKdKMjuLXOzb7Yz2uhzmiqRlzODQbEjmBmvz9sJ9tmOatiGkLeiY8
1TQhKDTPn6VOIBRL01SHlBDPe3jlj+Ybh1rgSU91mzs3Ofh92YmCpyT6VTlbbZPD
YDygtNlTylzXa7HIhXgAJBrbjHq3desx5jijKJtEChOEgPBWCr3wC5GIRgIDaMUD
aFc/fR44bF/g6pDgeQoE1cf8NUUjAGaRqrsR+h/WbmsSo0sa0beMYwQsNia2BB/X
G4Dg0MsoGkodIbsygCVhj6Z/D9L4i04EWHNBcAg0M8ARaXVhRNAmbpCEGNq9+r8w
f4j6j6Nr+gFvS/4I/XlkLvLsnLC7iflpiVAgQIgdoI/5mi/AdVT6egc4tgEOpZpy
aRDZIgbn9j9FDT+bptnHiPq4ar5nbJZWrKBPS5zQ0SbWFWKRKBCk/67Ju9IeGupg
Jl3MPAkytXGaqtNoAiGOX3wDtscZ2HggIz87RQPPqVX3a+8A088Z5Segt3lxqfdZ
GYT/YozhgFYr5fJHeIhOg/kvai+6GdC/0WTbhbdXRfoL4Hus3DMOwv8MKF5tc6Qc
oIqcjDtItZ/JCTFnhCIBTUZl1dkoLQwvjsPIM6bZ7XoH9Lk+H/HvdmorrOqiQ+X8
xhTT6Rs8AC6IO4wibSApQ4RV/sp2Rzz9/aAIbxr4uZuTG4Tz6G94QVLHEiBW5yEw
e5fmvTdY+1KDtKwo/Yww6sHz3AlcY46kbvuSSy85ygzzFq0XuOpnGxJPJlSzyKgb
pHBYc4epbkqKYBLCStv5G6V5oVcOTxt5jPZFlOAEnGfTQ4BF+/4CKUTcKYJtPTIB
ruc1qzDdnkYVSJnC/BNoIkHm0osj3/pARJ/Qx2fvrmz0SgfUScLcV1u6uIkXLqJV
VktS9Ptz6SDSHYsBwhPewPxxpdY5IyEv9hWlCtGRVESCk41E3ViZUEuPNUgpRMM1
zbjr7OJ92panYQXcOpMkOrOlM8txrKpOEz6YDTwabuGKeKAo3gH8Wky4Q2wKKq8j
ITp0JChyfHiA2cVkAU/sJvk5iJ6wZV0wo0K6ILef3rDX8bn8JDFaj2BriieldH7H
tRvP8BBszig5vNldDCBgpr0f4QvlBWkBL3u8C0SOrslO0KPBAvDdLS1GllQzu/1z
+z+1Lg1pf/0E4HDwO0jT+w/pAG4bVZzVnlFGRz7jao1UPElnJ/sHaNwEKgi537ow
7pCjrVUJCpNaojuYfQ2cbxByDUuuvCfA41VF+Ksk0VFrMVHnNvl4StkQ/78INH2M
Ma5qxZ6DdDk9VjuX08BDvikwkfx3wWwfg560wOgEDhAzqvIUMaVJpAOoeJX4ZMUu
js5s6STjiejJe28pPOiaZ+ROuuf/4z5wzJ8HshHYEhWuRXr8mvYSgT3ljaNGUVXg
pr3hNydOdbIQcBwQZKUnEljkG7iJhYEHkFiTWa3s6brBDVdikAZsKOMYLDdqE1qs
S6kAb8qDP2E+T3XCHALDszYLqUFvajQuTzoBTctfZV0Bp9LTrhCsEPgcoeW3xVku
q5Is3F4xyJNj9ufRQ33wvRYKM3Tv2RC8bNGF0xiIEMPoKkUiKlYuw3pbTHZVJHNs
NQgO95Q2Jxo8+7UKPzAt9rGShTjxxbh837/VE0iNpjqmFqJDHkInPCYyw9nz1ZcS
qP4y7iB8p+ILfixjuDLsrKqLBehLXKDJyr0+7asps6YzcxJ416cbnTIPxxHqFH6N
RwICLuym0jr8/hvkW2cVczj54VjhGwDpGqlkI1UGMrPDpFMBXJYOWeKwYq3h0VKh
hmAuaayZH0ortoXKWrrurduS9z9tISCEwGK1ivo9zD1Jzte+sqCe5NrhKunAJP26
OZeF0N1HuYEaBjbbZUSj8ix6abDlTjT0Y5oPm/ZYhbc6gB1gIx3n3Toq6XuNob/u
zRVmduTlS1H90C/5mnIdXF3IEqjNO8ymRo3cDQ2M58LA6YdbvazE/cfr4F3e+Ppe
0mglVNuxIHtB8LqGysq/whZ9uOrC3pDD1aXktpyUpDMaF0GB+AOygBbTMKIQLjOe
BBQ0pHYJvkcZ1raXVB3iV5jRuiJ4aXqZCgcvdNbp6ZCiFGysrOso3QHv7GY0+Z5c
5dytv0HAaEf+sO9anWPPO+ZrusFvv2S+XgZHCc4EXK+D1U7wlX2417ZQbMmSVlzP
oPadffOtEOWTKcNLv4GNOpnjtxdIcSpuVQwy5pIp0g0xXv3/wGHtrd/MmvnzOrb6
DDkYUp10CupOBCEXFfG2jVMBnFT395oJKfEkarjIKlkKMJ+iYvE77Fxlf1elcrLL
fnb3PbvU2T3D3EMySZ9sznh/IGB3X4yU1DtRymhmV93n+vZEp8u3atq1jwpNg3Di
QJZSkA/sCIxhAKID16fCX2yPBIFPLUOJFpzMAwaonAmoaFQKzj+K+nixpV5EGyM1
ovoPPvUMr1NS7byXOGq/yToiXJUNxuFyhKGXujJgVsWBV9BVT+c8EnQnxkJDHjF0
eL0wWCR4TXajFD3Eqp1oq4HmAMDTOeayqgLJLVKRikloW/+yDDxJspy4PjIeg1mo
dWUE+yBQLNad4O0b2gEfVE7xlIc9uhHumq+zeJkKkYcMSVUiqEclZRIBTOJDMF5H
VqGpZHvwIBG2rkN1VX3zWxAKSwvLkXn7hsXkBfCB09yrZkJrM575ncDRliHnSQft
x/fDdhRdF8tEf55WJHN/Fny8ZeN6akoPC9RdebuUXACiBAs+TobQXOiKolStnYpN
pRckZo2TaDnr7MOb0icwBB1xIYeGi5+xXGoE8efTjk6noWrltPHhYvHukZ/aNfzi
puHQ95D93kapCQIgBrNsd+eVHRSPHxEiiegUAkUtI8r5hYM9fbR6hCMhUeJwb/fg
7Y4xGX6yT7ucJ4f412VcLXQprW6Ax19bLTH6zKJXCFNZJBGmvM3sHUL1pkhGo3GC
DBQZf8OENSinNZEUhiAu1cLMBK/mwcSkMrHw2NqYC4F2XxsGAxDvObDJOwCX9SRV
u1i+/ilDL8+5O3RrM/Yp1ElWkLsKMMiecMC3qDQYczyCaoo93p9KYFLlf+tE1JtN
lo0D637uw9HoL1Wq8qBmw9cDci2luImhSU3otMnRkQCZ1porfRdY50l+3k4NqdLx
Bp7s6CcMZr2PlWF6ZR1OgX0InS2853K+3BAIPlpBeor/7uvR8/ZIYZIaTMpncjXX
K1NpRIRV0IneyNl6T57FENgvcg2O+faRUsZaIVVTUSe9b/3Mk5p6Rg6TrYIjh78x
Gi0winhuXh6IAIAKyx6DD5MTD4yTdEzGP7B8FKrUlTdkGkYBvoo2iw7Wi82Q87Zp
MdDvNVgfvzy0wctqMRuJHaJc4PZYk120PqURH6Z7rLBeThVupVTzSwNOCdIVrZCJ
ry/JesKsgPwrqdEuuWdWa7fbAwjbp0kjJY5BUCq80l18q6H8y0Axn1eJ2gY33SQh
sxc6mWg5getDWJfwRlrtx2Q9zyZTcOhyMWHK/cwjFX7zSUYPftJsgjakobkVK96/
VV5EPt8xOR7IiDMnC+4ooepLcSQqi/FArMtsI8o1wX8w7yPOHe14iETuE7lMKn8J
UAau6f4UMIPvy0yGVj9ji4tHnRUGhCqAEQn3t+3rm17QTVOwh2y9SDnA09vROeaQ
CEYjWXpwJ2cMptrunddaTodXZVgry6N/YCmGeLL53kM4hQVnfmi3X8taEJWsRlIO
emL3I8czlyoT0bAAiFiVfS1MeNCYKpO8uSWDgUMa6bola1lNpBxIYL7HDV2Af8F7
XuyOgav3+S0IXOZOTieIRAQYMbriutr5UQGUIZQATVnP9v37I3CHYUIF97shnULu
eF46go8iXyug9r/jwv7bsPIaKq2QzS8AYZN3AYwqDNmjbjiIorwmwUPPKrJTSkLy
uvUNBTkJ2popFrhLIeNhCACuTcUcIMTg8wkV/ThhfEeyYl4ZgmLy9AGXXdZmCbEq
toWIoas8I2PsTcfkVRPxYL8kq/p6d8UK9T5T/UmDq6Wj7DkS9JNyT3+TgET+9zbv
j4KC81veEIj3MNnO7zGdsU2TyffpgOxRsMaqjGZ1QT5zG3uTnwNc97DpClYOu0Ym
zmfXnUfHl5uPt+V/z/An4aqMZ+O5WpH4vFHW0AHrF87ILjAs41AWa/+CrwGI4GuP
RsdMDpGAEz705RdPfFH7Kh1df4SW8I3Wag9BU9gYed3pMJlYYk3l/O34IH7B6fpI
L0lmIt2EWBZHHeKev3t8+U5ogi7jSSw8exo9PQ3WnR/vj7dwdfXw50FQVH4gdgPu
xG2syVW+KpHQPKvVaS7sjk1PkphH0R6CHsepF3R46IelPTZv9qJHNuMvA94Xu5SK
LA4TKxFJViIWc+NsRsljdsiNxxa9yZ0kKuGNzT0NCrNeTuozViKWQSpU+0iiDfWV
0pGj8Nn8cOFp2ciqRxt4z7V8XeJohGd64QHYUCt9MJEquE5BGDUK/VMw2bgTHSCl
QgVuGOkZIWYZULf6ttN5OV8B86zbMkzSmd70zZsdzn+D3ysoKgrkMYeWYDTvSL7i
y3qptolXBH7cRSjXQ59EjMhiUtPLXd0NfLqXIPQAhD7h69HXN9ySFlKVx9eMWmq5
XGRQ3KN6PEAyKPeGvU15jS/U3toDobXErCRP73wGa5Nx18FpJ1fuCsKXgBnHJiwM
XV2ztOCfvumedsAlci6aTch2bNdjv/OwDxhVkphtUo3uh7Js8iWMPnJr3cDouZC0
T/eAD2fRSMpJXmSU3baOC9h1VCLNqCuBcpgPCu2a7Kf9m6uqPN4oR7pbF/+0Wn6s
mj/vQdek+svLzGIIO6RjgZMMvw08VAiR0FpiyDUH1Z9mEwJ/Kv+IN7Uw75NvYjxG
hHxut47df0AlV6e7zFKXxgh8Uvgwmwp176Zd9fOqGhCO/PayW5Eubted7QgSj5Ik
YkciAX3TOioeJNq5g1m20TKTm7QuztGVqRgdbeAVXhdgxsl508T+HGB1N3kJ95E6
9E8Af4EN/Nt6RNARJpGUYoQgXK94GyGuinf3m0KEXkMlPGFEHCRDHFiCczVhZtin
VdRE0Xth2u/DYylwmavIJc3k9Dq81L7CaRByy6FxR0699OtvUgq1ZfpjS/1mruuQ
fUYYNhFebkeIo5SSoSwQQkJH5mCXoUOz67ki1or8mvc/rupgsJc72hCZ83JwfBnN
XSB2jk2+x9RFTPuRzNg3uCYM0GIxsDfy49+6wcVHz3qdzhfkkajAyQIGZiMoJBgX
htvdtccGwfW89vw81xlxW1nH3kHqPv56KfxMSIoSRHXdrsOozUXTLDV/3QmOJdHQ
ybHZbUR8sG7cXJyiVyeaYjcDVBDpxS4dlRMZXakRmnLAbcccZzRGdeerpSPFxjVT
pNEAIjDUHz9yO5FXjBimno7s0O4H+lSiQZo3Vn5LS63Ps+I/JIBtS8C2WSdpt/yB
jaXY8zC8B3q1cLXfpEJuzwPF7eblnKCp2M/hPy2HLocQOYaCtxsE6AjCghsvWX9B
yhOfPL80P2KuO7SecNV156IqUfi+57NF60Xwn+NIMz9Htxn4wUlbfDXpCZLLFnD4
cH3zZnAIcMCLsmWfkCY71gGqNs0F8f6ShZ4cX8Sxfm0yi2hocZBxJn/N/Fba/Rot
VPSpd2voD04qzs9+rDDfu+gVR5K1gzjWps80SLo+O56T+Lx7lwpE2W7gfLLV2eR1
U16/6qU8w4EKT8rKDQ2Yig1/R8+WTCIyCtd3dwGJ1BBsS+E+RJaO0ICefzyjSjpM
w2Ck708MNac1cKPmr3qF/8y/4uqHiNHoptV66+2siMMamKtqeE7yT8vwEDjsC95u
jXeIP1DG/DckWeIeA3pi0ebZ7p5HE2yml/LcNj5n+CnhHkxzHdmb3RmPdUfrn0/9
tZi66/N7V4beCtPiAbGAsWQNb1bT0ClmB7V5sE4rvK9E7i+BXuNgws4LCfUhCy3y
zwqjsd9ZDn6isXlRxWQ53ex4DhSPdVMDMJNudM6byF/I9+K/VeU96MIRKzgtClCH
U/WnvIhRhGDkI8sjCWvCsm/9n5fKssVx9w3RNjETrbyGDajBHFAjFDx1dSkvl0SC
DOw5JKxiabpe25uLQvzrx96BX3ukjgw+bwe2t8OCeHc6f1EW09xH36awj+4F+9XI
QJNNxbyrKSON9s6FU1BtG18rHZiQu0L4L5TwoSH7Fv+CNaIHkwzwoJa3pnRbx1kk
S/wHZW66VFxRmI5EY7uLIbT5OXvDwwH6q7T4X3klJqCphOxGiwJJqRyq3Xf5A7RS
YEC397BTp3Xoo1DE95AnNAMvgYM7/KN5JV6c9Bk2pZnyqeKWJkxq2EXuxX5Xl0ln
P6VlFwklmvwNEvi2pWrddizTOASC85uuzjJn6coBZaDHlSWPauIcXze+x5cYFGf0
yOwU5b4bKiYMdpGK7fNRvwmb5tyrUcOOWWJlmRSL9wiNFzUAnTdLmJlbqTJyGpUb
G1HViXHXFntn7NNizBV0snb5GrgPQtZkPwepvi/ilRkDXTmxJ6nmHewLnKyQkSVW
qF88kEL+nRun7EU797p1WwmMBYUbF5GfFTlzesHy5j9FwNrfWtFTjZIHDhKrNir2
Aq7qEDiIi+EQ7f8x+cZZ1dozXi2ebZSJ3dC8O0wwRYQf7qpGupcIJRSNGoADfOZU
GItu52LTnV7cmF8vFHfuRjMHqkgOaspQGpErRJsaC9DxwpsaQ9MEQTEGSP2w9TgZ
zvGNO03ZtWwraAk4Xx76IktI4sribcUEhjy3qMwQYChXbTZK0i7e9VAIExP4Mdcw
kHNgykFKi5ow8Z86DIjupKGArQxweFXI8GfzDHjDTetVl0mmpzjBoU4S9lN/2hb2
WxGPBhKRBPI0w8OU5VZPaP1dKHTjiRFGhcidt6Rv+0l43sKUjlV7V4F6CmfytPP8
nS+fCNrV4pAgTNsAES8CjlMR9HmxXvuamPqjMXadsBmykJccW8WjV9i24w2x0MEs
6MsQmmxLTvpo6MjSBMR6KZrtTWJu19bBK7w8Fk1YW6fyhVBDOZaXuqb9UjM/12Et
OmgJkOzQ3tr79/xDc1pnnGofAjht6MW1w360V2AeJ/tfystnvq/Ir2kZVhdOgk8R
/saBZB4ROsE8AunhBsjO3USx67xNBvrwXlwtQeegqoqC38RVI+5ZTX56yxDnWjNa
KAQUs1RY5EvkLyIxNodWFiCwh3Ip96Q2t6EPUFjgBUtvQc19qZnM0SuEWW7KFjL7
Qam2Ow4lzdQHvSNROLzoeDmPYDfojQH+vQLP2PSjGgc6G21IhU8mOiJzF5JUQr85
bm3oEboNeF5mROehlXPlhg4i4FLPJFT+siIhZ1WPukB0X54sX+4SGqfOaOtj3qeg
7ajYEKxKInhqun/7fi365MuY2IMuzK0Hud/hOD8hoqINm3tjfjjb1YNR3lO1Xdb/
HqyMpbbRmyfZ/w9psLZ/EhVGZie1YOZ3OqiGT5WyuC2ta3tUuAICssySjOw6Hutf
YT/fN/XjeqNn4qsNzPN6NqCgvamZ4ILXCT/HBfwK+6CLsIzhQBYda9cJpbbDqLgZ
HuO4K1WNkOhNruqZVLkuaENXiP3yI7HXvhp5Fz2Vo45mMrdUQQzELmTAze+HsF4w
A7Bj6QNMvDbc+T6szltShMiIUwudDfuhaBYWtL6ZXNDRdkKoi+Liwu9230uDZzQQ
Zoho1kn5dXJJJHw2jk+L1JI4t46C15bHBEZZQH/eDEOrCKxFynFkn6MEN7/igsxm
jMjrZ30Q0CpZHgaXRtnWF0e2lXVwcP2/clpDqKwcaCmcV3fZ/0GnQ/iaM8VevsLG
LBRUmjGWOQyvDSFASaOlV0rd14rjxnngiECjb0wLwpL5+vFnyZSvXWzyvZlzfWTC
VEVJad8d7cnK6M7NNFuL1RwGaU8ZMsJ+ENGbjvAlqL5bceWZZK4hHJR40uhfOvsm
M/9BbZ1Pe0mVMhNg6Bd2ubW5QKJqujulU81NEyxvJKeiCT1ULvRyRcHN2CMqvhrv
FCBW9EQQ1S4foqXRfM90aAHOy+cOSRdB2zEXtR7/L/ZHACZpN3I2U6ZXbyGFVAQN
NPnQGSdD09CFhFWmt9Pae5aDP1K3eQDnaeGi00lC9hQxB6J1iHNmk+v39PQGRSPE
0/KWzg2hFi5a82KdC468nifIzJOXSK/6Shf6g6V4e7Sa8eW1yVtr5XoYDDUDY8Nd
P/yCjEeO+U/9r3c5lwsOloa0TdXwghk2Q9epM+KBHjKZzwgD60tXbY6ESNKKCBq8
MAZQ/EO9XfoRUU6WupcsAYxoBf/HMnKT5xv/Gs41SS7A0EKYksFIwUVkSnwCZ+SM
dIThJNjZlcM70fTAni2GewSXkwu9MurFfS2SLwQQkEfJjjYteqIX3q4f7qZVSlRY
XwqeZsxPqQqTkTAYCHymbpvfvpwXgZdVViOggMxrhhgJgCfF9oI2ryvRPBXma3yx
XmGiV8aTliYEST35uhvqa2tXJ+RXosvbf7B6B46fBgQ7USDv6DnXafLST+lnm2VL
J6mWQYbcgbNfQ13I3KdY09chpt4Vz028wC9dA5XWax+gSWPjuMLyDZd6uNXfqWn8
0K+z81h7c/AAiBXgCfTg19/yrNZx9k8+kMGzg5GI4TbP+0iqIstVJdgUc6ovpTDm
hsJcmOfBta0tZYjsytjbh779u4fBkSbV3AUqkRLQlqPUiMB0Q+ss65thLWXHOZE6
2OSi4nOiHyy+46G8qI3vL0EnfXZ6Vf9qD4olLmmZwUqV8tcM9x2+umrGt8itP3Uh
8/pPsZc/CeMUI8XvwtfGsHFxWQul6G7u6vVxsP3oip+udi6KT+BXrV0Eh8dWFFrO
5TAkWmiG+A24B/zgQn/HfJJXFJYskDUzAgkd+C/ZVMY54WzJ/oa5HugTVA6Pjjzg
vilPdFSmEQzxTRytYnCxFNgnJq2GhCBwRMC+vGVE7E7sp+jxs0jM1I/WAHQ3NqvD
XoaRa1me0p5oHaBtNXu+kisyNw1Qe5XBtjKQGU113w3/XT2+K/HK0c14ZZ7xXkeE
N/n/8ZMCRva6+K/avgwjSbinn8Ei6Yde6iRaHuKYEqoEt1llhlP0dPq/5jhvzMQ6
kNkg1Ll4Dn5JM43KvhRn7zwkxM3PYAELG0/6Z9x+7AYesCCXS49wtChLeNTos39k
KIc4QGeYa6yWqzEilKIQ3rAG1RJOhL/K316R2lg3m6lNuYa5kXdHQok/3oxprPCH
o8C4Yv8XCqeQsmbejWRVVbJBF0213/J3qrOTGsci2udtWXc/DX3hhbTZn4NR9arT
/FFoK2ncFl1e2X2rcsWMa6vL7MsYeg2LETA2DltB0n/kQ3Vo/rsxJPXjzeBntjAq
gM5Tg4jR0i2E3SFe4Oe1r80cU1imUkEd+qFoGiPkuwG7Ac97glYNqH8un78pQrTn
CH1v/AO3rt/iium5DbMeBfhv+csVLEnua7XnOrzBcivlsEWyiy7DW3U2xZn0zxjd
dt9fb8aIxzUi1aDXJJK/Q2rcuAB1st9hX0rb1/lYf/NZmcFgz8oNanRu4c+ATaLL
iZbdici26MuQEq8FGAEX0aOGfkdB1+x8vTSUQwEq8oG7FVKxBvMbO4xaq3mSvS7K
QhONkJ/gihz9hmUNVHlD4UQAeXTLo3kAq9x4QzHVuB+fc5IvKayJIK1aTD3WShUE
36M0yNpPdZCuEHtkwp7/db60Hg9pejAlyLb4KQSovkV2Regmmgkq9RWx9pp9I02e
Jn/T+a2mSe07YQmB9+haQizzmZ20YHrEO/2ZIxKJRWHgW0xeVsfyuTFos+YhASo/
PKmPRq/vGUwu7BBCdbuBC5jIXaAJ671C/yuPuMWgfEXVgUO3R0If/5zCx98gcUSc
jM+kpFpPDVd1CvyWAe2nKR8lNnlUEQgeIPJk8zlMdeJ8a4IeGQMRvrT0ftx1jBXN
FMY88B22ZFhaiZaMTTG/zYtjKvRUt7/oEq/X689HEcJafcWd2C7fi/E5SbwP2DG5
GW++estvMmQb49HZ1eaAw9jkFAxvzJk/Bgm2WLhY86VswQo/amAx+EB6J1onIQ8Z
N5luq1/y1DsXsfQKtxJ46jxnIXg1t9q1XwIeJNZMuz4OCailK0Kmpu50KF23JhA/
ps6GhlSLd0VLpnUYX1td1SW7i8ZU2T9AaqpULPdmJvM72J9a/DWrGRB3QL1lelha
ygatUy67RzPUgXwCXy+OWt8+DMi2uhkufLKNtPa0xVve5o5L1ztkWv78BeCmPD0A
yTtsjFgwnnfsuWifUanYDaFz5o8LsHwrIDxui5WQl0ZU+IojfGo84OYNa3u8EWZk
nt68/BDyXQLnNIeib7TOFv3d2P/oDkMtcJXHO/XfZtkJH5C81KfNpWW/IiljRmb8
HrhTEDbfbcGOVHi7QUeQfKIKO+mIUU95j5t/4fRd+DlxaiDaDYfWjYANieiZXu0u
cYc7pPF7VLtSWUfVofuycDTgr5QCiKM5PeoBs6Vw+4hxDiW4SMlQo/ZPBHW7k0s2
iHp+27IymmxUcTsNlyllKzc44c3KN+cTFPNe2W7BMWBv6k1I0H2ZYmTg3uza1n3g
hEdfBgNxAwIS2PdqSXK+XCqYGaeMNbEmq9uNi9CcCkX9dCQSFhh+zthfcmevjKbI
EjGGg3bVtmKTg2HgA5TR7iM2x/mY4ugQYq7CfNUJbEQbYTrBBYuyhWzBXplqB1hC
n6qG2gjzz/dxv6aCXNfinm1sJWKMTREffUZ0AdqqQkG6kny+oD9AT0PZ5m+OHuh6
w7/OTtt2DNQiKZKSpaT6TRG/QtKKrG/rHXPTCzor4aFHYjQhrNEW0kgOTCd18ZLW
hB7UOP5uI/rxOe/4P0BaN3Xq7vmPX29cBES6cIonDLM9DRWv260tLxyK3g9icUcC
IXhmBbQfFjrfJDFmgCi4RXNSRgCK7tQ4o0dfhhy5qkfLVsfBc8FQ/yl9Iwz25KOW
kO2WJTGkFpUdLM4D1jWz97Ezv3Cln275UKdselbZjY3op8cgZObKzcEptlWdSfIo
1IEvpFGnHCi1StEW2OnuynuAxOpmWk9zay+/Mpy2Ew9rWZW/fa4IaxYMShvslThl
bvQ/h78Z2yIrfSBFAg8YAsEHVfjz31Umv66ECDqU7gkcqzCw8Jdtc52xYHZaBwHy
fsPsHWlGpeTn2a4xlkJZ4yQrv7ZOYizurPbXHcs0hpGE+UU+RKGLG3LwBXBwnbew
4UT1H0nH6TyHlRCsxiRlI33T6FRlFqgauTL+ezrN8zX+LtPsj1YwmgMXIJ552Sqw
dMu7NRcX2POv91YHitErODRWtBsq2hXFPvTVTjafd553DgFt6adAZbThz745+/q3
TBpdBneS050VEuzU3j1AeN2Hr5YnZ0jRQNtc/VeMM6T30yQycxX9hfwjxL17BgaY
U6+gMUKlJGfSq7LJX+Wq/Y8q9kgkf3nFAFCkJGYCOQUf0fHTVEmaJc7bFyL420W4
bCLy8hG/Slu+6y2QQ6c2nYIr0H+ifNd2pdsk0RI1eWUtJOE83U3nodg7/EDZHYJd
pXRbgk4jJSOXS1ck0WH6AzczEtH0NfXwCAWX2U060aZDRkgd4+RBVjb14NA/qI03
nx6rBC4QF43GbQjtyHgfFOwJs7PsRs+rq1momu/BVWefJcvLfOiPC+nO7ChyykL2
MXUpVccsg2ZWZ8MavMyO7zNtkeUltgCIlbNKgIDfZcLrBCN3MgKeFMopm58za2f4
KBHvtFonzAgR6X5XLxuMTYb+8xCDnNRrx5+KOji95g866mqoGdaP5zpTcYp7c2GK
hidtTNRkqx010xapmsIDoWcyga5fi5+4ucONSpYwPbandoyOQeaQ5I7pMIz4GOIo
jzsa5Ks3hKiHjpmDrZqOXgVceUCrua5wbwH2iRCW1QbjWNXEDL+pJZSJBvcJ5BaO
oHIPQRCvU8oIX8snSGyfOBQcPz4JTf0BaA3OzkRm07LYPoWng6/np2eCIXCy7ezg
odr7TsNxtbAAYxuGRfh71B0eE/k0OHjako4XGGchXtzeayblLBFGY9YnjaK2ac39
YQcr8HhfUi9WU3VQxtc///8a1D+tykiC6zZYWWOrv+dUjsrd8KVEiMis0HLwlXx6
4BQzBHuk3dvQpTOf+5PIcNQG2ildj2OtdopSfMflTkClnu8OlTKflLazitXdUKa6
vqpQKQqA/euggr9stzwwaD4ED73uiulDyCt3I4CJLH+DLpRip0S6O2NT4mjPF3kL
M5o0QOWd5cTv6x2LLIP7ftNmSStJbT8dCyTPKdN+dF2Ay/szdK2K32JNGKrjvhfF
UbGOKc75C0N7cIWY1ad+akzB8ypVAyQdCy4qFJxw6OCvIMNM1q+knvWKBxX9NEDV
C6FzOxkfcijn/wltLfPJxfEbEz+3GHAUFqC5vQFFoO/cCpggN4zFlXNFdA35njZ9
WhXo1L6oJguwXJP4+8LyYI2Il2DpjvTlCAkxSkLJrH7IXc8vUEvIPRWgRHo6RNEZ
8VRJESX4R1sJjomW1ufEK+ZGer4oswSEOgtvEuLt/r3DZ1DSz7BiSO12qTMjBd22
BX+2OpMh3IzRq54jWMpQJTtNCDyNUieSxCQeB0xlPlkOul+6OS6TGHFoyhUkC9fL
lGhlE0vWvyA+HhnNOxICS2oglMlC6Jq+NpVqH5bWlwG+NeVdp+GXF2VZkmaYsVo4
2IDP4YMEi8hOVS6Tb+Hk4sHT463TDPluaGKyFDGwKG9+UNgiRX9+OHnKcEUBtuYH
ZFWGt+qH+es2JIFobvC2zb67HNetueEXVFxJzVDXEixfG+t93Wig6cgwxjH+YbU+
02G1qHKbEpzkdJRHfwevZsoN7zOEzV5oxDcY+c2AmHQaPKuXUA6SBbH1TGr8HRj2
yCf/2SCYJs4DSxPs5SM/o49j21gGS1BZSVmaah4EfooEeIakxMPsgWyyTequ6BOk
5hCuEYy4a7yhjTIxztfN2nIaw79qSBm/nHpS2sfmhW2MBAPmHid34TRQ0owX101s
CFCZycTsrKVwqESnCCsh+WQng1cjkZb+PgATKWDmKEj+S///TXhRz5W5LLf/u3EA
gfpWObhJyk+OzqUDx6k/QYyHt+0TfTz821QwGnC+wprLpizaAQU3BUVzEDYAPVOK
fRC27BrVdm+qqDMUUqSa/FkAlZy9lrxI9umF5vKNJYhpeOY15AEQ9XUfwiVouKhN
/Bx0AWxnbiYqrIYWNwYDj9nFz3DbjgLajSwnBBnu6hd8jJDN5vkkV2yiDmG6efAu
VzpvbH0q4wVdJvRbMKpn4UGUrieeHJi9GA1xau5FcxyGpagBBDZMla08usbfp63w
ZVG6BF8Md9mRMxg482S6NaddEdZ7KLquha8AfAtqc+r7ue0Qtwijva+SXRSYUrYQ
eorC2j4dgkj1InTNdB9KYUyDdjB31qoliw3ZK+sEXB4zHoB0znloqz5NZ3liOjrF
D9WxX/832vSvNJm9eXenySm8pB4p1w6NT0jLFWpsJTjFcYVesJZNAtpWUkHVeGeJ
zRHBhHaMQiliZB2ddxJsdc68hn9WVwMe6Wf9BX0YRrnqkkohmcP+RGoKruFTpXhS
nRgB7JexD3uhBR8gLl0GRgUJVz456LpdXLEluPhnUp30l1122Brh2TG73k7JidF6
s3LR9s9+1/lTZgxaHTewOSR1PmmIhatIY8Bqaq3J7mjfUbmJriuKJojrTh79ldVW
aC1EEQrQsGDjDeEZbgOzrkYdywEzOjZzPVisUbb17fK5iK+hXS77NK4m5mlDaDVP
EoeupRO7NBoxFcKsHWzSMKKH4ZFvB4p9Xf2fFUTVfqkQYTYKuVzdZhmF/AZ5128D
1UHI26CkVUjtfuq7ssSsQCI4EzL5NxsvL4f43hV9yayQVyNVoGFUFRFFR2HA+n17
MIvUOOT+4Eh8sbuGmDBfybBVJ7dyoMoIPjmrbmyvkUn2cjJ5yBzjvaLkanrX8cCo
1t2Y8CW9LFDRp4i0HOXIwLiivpbO0uA4s7Q4o0H8JL6CVbk8FptEJwxB215hfFrf
fygILVFiDn0wEhuYl8Np+jSuXI0dQ5pNt+Twdph0V5f+LN998QkPaMR287zR6Mmu
m7dM9hf7Tx4I/xa/5akNcYae3dyTvB3bb/8n9qp42pnqYlODsQKnlpz6j3f/YtWD
blNOC7aM1k2q458ZYu7tKmqWIkKzCYhPE0jgIAWDnY4XHhqAl3K/4DDk5GAM2tXW
oJZj2N6qiYQk1cQSpFc9qqf9rvSCqmzFLfHNqzOlEL7XwnLm3vD2/8VwKEjjOvft
kTF9NKb/FF+Dx6tlkp2MFvxW5CUIHgc5nTgp0T9u09UYaQlNNMXwPiOqYlPfQro2
d3poHhIKMpfvanYRF9VkV+OEHG1MVmEOKDyjILqkPqgCtXm9vDLU2bKNSLKfzqmg
xUmTfLnXKaQNCvlrsPpyNaUkS2OETF0HLYoxy4jMGGaxqJ7wZ8z1+oSv/6vKxFLs
NY0OcKCl5Q7YCp3mnQteGaXB6BHFe1vrsfbT9xIVV54V+HQE22z2MSN2u6DzKNBb
R7KOKSgUwf99w66iA8v3xIjRB4MVlA7IrOLToZKgZIVsKI9TfcvZ+E0rKEUSQqSh
tX5t6Lv7TBh5rz0mGAy2cDaLtOsPEk3PyJKqvwv05ctIiegKQiCYYl+MiUvLR7Ks
KExZcDyIB2ZaicCdhx/IEOBIqKCC6wdB+IyNcoKa101mG/+mEoga6ULpvwpbwvSi
a3eZrIqyrsmJCw3yZD5W5Jnf4OlNjmDUbnPu56jrIlm75GyEq6WHyXGSOcWbjRfl
kCY+g3ej2tZqbGJUTCH1l4hc3AUB6nbWxAtgSVKfXovewr481hGp5RbME/kTOqJ9
AFLQGuRpHOSoAERcf2QUBEjxSQu3yPSDIoxCJayGrjzdbeo+Vho8uTHRvSjPIy+0
Wh/qhQQRaqPlhmx0UWJCnqXYtMYYotGiQutXy3YoPtHWFTbwaJqqAwgqeEtuCL8V
Kq8TabpLkqy3f+2+ytqhltcKMLAXNG8OjgbGbooQ1Pc3JqSldOrVxquWtb+WDAUn
qMqXxx4EWj9ZKYEPZIBL60HKuDQyjgMZZYRPI+zq9k2+wKdovky+wZ/wLRzYKSSm
9ZHtAfuB0ND7XG3xQ6qQv9eM8RV8xWn5d0wr75nWK7C1B4UbxtvC5mmimGpMyOfa
pwaTxIynwmvsmcP9MVzbuEkA2TaLnHCI1g8pkACTzH7fc8qYb7tzNJzT3Qo3NL4v
ZnwpjCLR8tJFMJJh1G/tkrAQQt6Jd8zLefl4zbi4YLwNrmHQEHuj0NsuvxBgcLqh
GO6FtgnFN0RfB2l8+C2WpF/ANjFJYBjBkmthTTAX1rAZ9yv8zVcqwlJ8nYix0iHd
MjqpNMtZe5OnsVDITjlqhS9rGbRlto1OmFjLupuskvbtBhKuHXzXzsRkRAOg/4fY
eztZNs39aIk1r1K+kmQLY3zob1t0vOycpCJTYnlNsSb0EQiidbEhwqVXt28Bu571
zzgRZtbs+ZnFcXVxA3cCGeUgglrkjajsvKRkpTNg/4NhXZsHo5R+V0LzA+wkRrtu
ybhDxw+VmApuT07ZCfI1+fqQ08fFxd7iDgMiZEuLI0Q11opF2UaTg5oG4FML6K0b
JNX+TeXcOCaYssEDzUnQdD4RRErJvEw2WVJ9KIqyf4AvjG8k0xPZWqJahrGBT/7W
eyUmtAEb2TnIt0OBOsu6H0r7D/Pf34h3l8rhB6FaYaUFLt7M/wyCMYqHHP4BEC1F
nBmedWs9cBjt9ypL2fu3wENmLnJ9GtsKqNlACrEgGJrCNeDAk+zScWrPeXIyByfJ
xnlz88sv4CgBF+mXu1DXkWDxmb2q1LPeWUHSzco4aV1UKiDxg96uQHuW8dppupO/
WQCVj1uK9rnI/rBq17o2MTrTx7vxRTM/q9RRseqcqcrDJFTL/KJx0TQppZEc/SG1
tCcWEnIVKsp/k2Elkve58upjf+tgEdWXrDZVhnB9UqxiROzhOje3hUQraJFhgCN3
JyOrPDsx28dK0twJcl319ciYsXMjKIG7YJFt9mRziiz/NrjWEpNFmvaxdUwHnMzA
Q4+WZTN33mPPpXHjf1im0MU7+fr+nky8J5JuJOJwmTyRHDyG1H1YzQBPvUUd9xB2
nm9KymglXPVUvR/VHxi+Bngm8wFD9r6QN4duv0ljymkpk+cZICStWWaR9wqVJ6dN
Nmx/ZV05jgi5d8GkEBqzQNlNy2WrQqOjNfIkyTTAbDD0H8d94CzmlEBckr051HR2
NqBmfe3QIKA1nogVl3helF4BQZCAPkP4lllhNEOqyJCOHs//3qA8DadgEHJCM5eT
TVYJbFMvAdo4naJ+Oy84V8edVnyOzPeoE2r/+kO5+yV2SzDQzsDwDX6GJcEVbpxN
dKPcF/wWpJIj1z+McTk+gn56TkutMwq+H6KogD7tg+uDOGmCG+F9nIn+2b9U2eZL
IrZigUpXRcOiVdLhTQFncpFXetYjWruw5ITyy1CGHbeHBgQDMOvIlpbZFIFkcH2f
34wKf3qrI9K6fvIIeMIftlTDORWPZek0SSIWbROUf1j9JUvzwjW6Bo1NJgidN3pz
mbJXx1ofvjown1KYCDzCYI4CPImw4g+e6qViDNZE4kQA1ZpzbcLHs8ncC298tz/n
nO68OZvn2tfjlituGCckOjwMivmpclz5JNdi0oAXMgpdfUK/FWsPwm/8SUxN11uq
LnvaFMGJ1h/896oCVPnPQoX0untpwj8sD7r72VjldrF2mpTaQN+vMtHYYhHUYWlG
4QHm1DnVyB7jSs9iFutmew2idA/Af2Axy/XZ8/HklURXN6GzQTm3pW77DjDSgpTX
nimKDiQ88p+6cW5+DH+YJRRQicJoaozXFTWQOWBZ/KHfvENvaw7e/FAGDruZLLf8
/zhaMMHQSeXku4iKkeS+7jCEeSuwjz2CVZo4dVbRzNic0VbCXhLdtdH5n5PVD6B7
LNgtkKCBsseqpMWhfRIhAqsqgPsPZJMJvH7RWLvakKUxzBqVSkaAX/+kRvaHQ6cS
GtmOGkm3w5QU42fNLsCqbOPfTv2ogasZzzUg9MUnmbR3ALVgP86BwPbmfM3MLF1x
WhLXxHX+n+TymYPw+XBIKKaswFJKwhPrMTvFFJlziW01Bym5y2z7QPKNs11JfoZa
rPw1rt5er2JCq0fhripZzxkVmTkO6K+rNSX/z/jFj1sdOLgi72KgXi6ruj46NVMB
sZLct+Yk6tmmjl8WSGp/kakEfs6rsrQq4IHbF5Cu9LMwVjo/9XMJJAuzpqVWcUko
8Vg/72gJQmhYozbw3Mah6vwyOlj5RohjIomDFKkfgmOX3lit8OqYUN5ZCy5bt19C
qL8P0Rau88AZFxKeBj/3DcHriRWOFd4LJ4yI28Tv8+ieRZzcWDCYTFxxd+9HMJOq
fYQG/IXxV1hahiY4FAhL2wcCg4i2y8B58kmwfz2JR/Z/hrU/RsbuMEhF1/JDbwh/
M0qWedP0mchCvVa+XTfxWIMnO1BHnOJxtJ2/SqJrtlAFN+BZe2w3BabAdk1ZUfc2
uzuuB9UjJZy307FlYSnOXHhjNWbwdZ5HIfPfSUpec/MyQGYP//3bgImv6+PbCkvT
9Tnp7g6FdZh484+7w/QO9FdeTVCxEYRYqUL7yzIkWjaZWuk7Jbnyj3BRwJaupLtY
znQCrn3oZPS2IUfOTdCmyhXzo3p3qjoSYYFAo9uDfwdRPdd6xy0ul+AdYquSQyv1
IiooTjPvJzeArX0geJSv/diFct/jy+vlVCnXHLoLs5U0TojNcQ8upTX6kLRhsm20
acsrI4KqLd9fwgQmD5isADkm8e4oafvg3OHEiAAjC1CeHEmLE4HJNgC8poQQeMPf
0EBFk5t4SpNNdWxu47QM0cu+NpHcn4+fFyEXOQRk5GZ0adzcxcipvFVEQVOz9C8G
gDL3/MLUFuRIq1L6Q9Ba+98/nqFURsCC0dzXMNSZ77oh/GCGIhXttEas4fx70Ldf
0dw+oiznQW6RhdRRC8yeuc4EPlNMJoZv+VO85oaeAC0Ni+SVN45Pvq2XE1w1X+CN
8uLHeNBfNpaIurd8bYeGXk/uBe6H9CqrEekXa0NBWBWA7fDlb0j2dEwluOc01sgE
giqGmEGm4qbryh82iqVgD6czeH+XzQ52Vd9x7omtg9IwnEaBrED3FYdobA3BVB8A
JfQJHk6iOYc2p0SC8HT68C2SGvnuAM0QvywkcsHvIMME+zY47if8JvcsmEtKhgwG
FMtYxR4U9vp4jO5t3Un+q+h6SspPmvnFqNj8+J/8gXIpSCV5/Aksa7IPAkn9WU7g
S76mehB2g+rfPkT5YvCHdeD3lHwtF1ixn7Y4HrSqYaTB6PykjM4aceQtNRM0vL/s
ve22FgyQoj2XYCN+c76s3Qyfg1QFA09gVdkmEEcJhbCI6/UlAJCMj+bga1Mmff+o
uJwXDvYlb2Ls3mmtVWUG5d9p3LbSqFRcnEFiTHCvLVsDe6DVlTar9JHDSfR6mIqp
qRBJJe2Octi0Vt40TbRvF9vesplLsuuZbvFYnKEBL7peO+lxH8yjmr6nvtOeieC7
VNdy1Q7C/a61CkXKXVPNBJu82DmI7dUH+X3aG/vMtEATI00TQBDFEbYP28HJtlfq
sHw/h24WcxOeDIi3AtRBHDi6AHgM6Etrw4fSxpSQial0HyeS3ob6/LSqHc7UR0Un
vRaEX1j589Vdfej2HDYjaOgOgqqtFVefxIXgH5qcgaazK3lgOhvP/Smwyo7lJHZE
3ZZ++NOdf4+TN1u8VZQG+tlsn6sRIi8cZGZcqfiV+mya9ktMzx1H6ZEM6IWbFdcz
RGw+eEHs1av8+wfijM6FexZ1SHG9jGkzCuNiNCju/7PTRJ3d/+ReEjQS9Say9ffi
iZzNgf9403b1awv4uL+mymE0eZ+Fdcn6xnoeAHuYss3kO+0Jqe5zYROtR7XVOn7g
TclJMvqd8k+ibGbyiY0K5DKB84/KyvsdZw4MaoRJ2pJIRvspGVNeR26hvuJDy+9E
Nz6hjpH7Sj1Xbl0HSoiVMBXfnwrfIRQjM2ytAjm6AgQIHUNPwxoHhX9BCWEHKQoj
HLLoDnhAcRgi22ain7wODnolHHorBBEDG3rYjZFBzXyseUITVWbtvt52dcOZ4vIJ
D7gr+O8lH9tWizNMDXFiqVTHrbPDt6rTosjPWTPsOvmh7l3gOqwdzjdaxQDaie1t
8okUjVn54CaIzy5TwfeZsdzEj82RN4F1C+5mHDqZDmUbIl2bXfvn6bwURj+0Ma/W
2sS372OLlaslcDamBa4ESndbAxqIyQSS6M/5oQXJpUhJL9Dbm2Yv1/dc1Dnvu7dc
+WmV16HDv2mAtY5vMqAt/EhKn6aX04NZ6+ZcTMiBGD2oGuHZL9x/yf9MlS9Y4Duc
0NdCKKr4yqRZ/zVRuV5PbhD99s4EBKly4hDFjF0mm3gTJq4QTiR7CQDhCrd9TQPy
VUHGtreF0tmR4bSYhszwpRhmk+REap2xwljoI52nTXY9aImrW+seKwv1Xza8i5La
wRhFep1L/yTDIzeWE7uA2733Mj1Fjgpc+UW20Q7p/wLXCJcu3/uZ2s9iS2zKsc0O
qTCvPsK/ljXMpFYwjZTfg76dvESLD8mChYtUZ6gYOS0N4eFu2KjDIIWYTN3toKdX
1A+nQ1pIAbTrkGEH9dIvULtsd+zeRIuR1p3WQkG0rq4Qb8NtJkgVQ34JZKRR99XW
xm1IAhDId3CRQQKfatg9ti7KrL08q8jSB+GKZEeaQlLBrW7lvAd7lSsos84AXDMI
nlLGV0VtBAzJc5Xgh8F7/PZeolTsmsQ5bLKi2UNztGVYIqUdMY6ntbwje8wuTST8
3NnrcF1k2vmYoyB4njC1PpA+JSatfglfvpFXpocq/Xz0a6ABlentHiVnngoQm1ou
3Z3Kd74n0VxpBFLwbcV7D8f1W6P3/k8IXIi6SyezGSdizEovdQRuOaFZZw6mWYIG
lQ/74HoaL7DRHo1BW8Iz0PIu/nGYW5c1MU1DvmyakJ2orKZIrbmh07e8V+NGR6MP
Tz7yqUgianV0eD0yaFnrkdZah8fjfVPutaIx/wESRsNm1mQAkhI8ksaUKYRqUDTP
uYsYRYTLo/fB1PWRe4CEDQWAbqEw2UvEtm6ex+9vhHvczGpMP9i7ommV6Za48ekY
vgngbHK21cRtfQFGTRRc/WNRcDDKo759HAAxqkf5DN6/8W1doQTLS7kO7Ra2R3kM
Kv+dC5LlMo/ivL2qG0gmEyw3xzbpR4Bies9K5y56HuEZv8wcUjmxlywjj30Z7LMN
hDfLiwbcl6J4PfYeLIT8mCN500JQ9MPzMKMqRHxDB4GGIXunZS/x9cEFHbwFe9XA
TLsn9fr7fde3AaUlhN+c8s5AyjYcmqHRcjZW+TaQJBUsbnWQb8fRt7iOS3BkU4M3
/nlly7/XfH0Dbl2FV7TNW+U7wM7DnXbdyrxxowZZuQQo3N9odlHKU90FJM61e2Ir
Oawz+3NIsYg70Uf0BxpKw0V9/DMuTkv56L/3MKZcZVTxlCb0zbCPuxgyfaEBakRT
UYJ50jUT4f00KHVSxxqUHqnAvMltk6+9EImnss1SkW9ZBHzhStJoGWLRUI657qTL
YYYgrY3kggZrOOVA96ems2sKP3Y5eSObwAFBtK+SnqyxcctxfU7jeGb5B2qTkuN+
/3Ce22KP13UY2F0y/73CK5EPx/DPRnoXkUydehwUGP2x28t2JOFfC3Wu9csyXlmt
kpSI+IS42lpe8AMf5bpvWTfg1ZV0ymFSHn2ujNci6PljvxnQQTFtg8ypAjhaKt5q
v6w9KGDKiYOQEqDP2l/YYeoFBQT7PURX2Khut9GUjWMmmUV29v7dwuOew6ipfuHy
1qVXbumgHt5sfpIP/9gcBmzsHSX1k3ww0EecqXgPWvXWHcqsTZ6K+Qwlc0bU6n4x
1sPOWn0hF/yWH0Bxj+ekiTFBo0oe6PMucgr1jyY5zaZfExqmDaSR19nSl4OEpt+l
wK73dDDKhRmnkMp22M4eupalhZGJp/vZ7iY0Z3M/oeH91J9fUrvWsSwUZxUnTQe0
g5KUnmtzM11Ck0OItVvoHpn2oJ7GdSrYn1cvNpqI00yOyHPV3pGHMs+OK02ZcFeW
xFppfjYkUqY5IpNEMtOt73d9ETJNheNxpnPtfxv9xKwZoK3HJs3Z+aS9DkgjJ99+
W9+zoVowUTPxvv5Yn7q520dm3/S3e2Cmo6RKqHc2E7Xy5OLd3YaI5xsYXQB3C7+Y
zCwurhoXQN4Dq7aOiGIUKImHtUAlH0QM8QY0HMwzW6Ur/F2JUdGmKW63WRLRa020
HIBM4CQEPvLg3qi8MYogYwFryADHuac0+a1yw/9JOlUvshhkJW0YGH2EkPnPU6oa
F9gzeAn9i+2wGbi5ERPinJfZNRdbyuryhTmgai78989m0Rw61UvYyhogxooEJcbY
ASS1aI7THfx9QIsEUoPXfxvPkkElHcOS9CUXiGoC8BRbk8wfVBngmu2o9H5nPULc
uxGbtG63iO6Nc8OTHAkkkxxsd2qCDNiYVVeNJF5pK88o7FfbwVjig9VDoY3+KGi/
HzmAdhp2tZt7MxzAoo/qQf6VFOPnUaOg4o0AQG8M/bfMdln79qCTDI/QKoo1PbZW
MPIXvXPe8fMKsM0MLdkQsjwaebqFmeS2hy5yb8c2O8H1cAd2W1soeZEBA4kpVARS
tsY412hf/fD0B0LKHaIhvNcfJ3YE9vTVnh+XeMo+CGk7C2XT99knDhg8KeoCLuod
+eRV1x/QRl8YqBnEI6SALe5AFy7KTkWiR8oNVoINT7xIgEncvx/ALqpakVqrFt3S
Yn1E/ocxYqD8cZwrJl5m5338E+Xjxx+4A8zPJOPYjk0ULVVNDpmM1emYrk4xGkF3
SUhLZVHzmQerHTQGvCHokWrY9AZT/nNXAwbNUKzNvaTG98PmrvKrPGlFsZJLa73R
0Y0IbznmrRW38xEIasIYxaPcfy5qo1y8wnPYIEqluzpUe9huDO9fZ4wbfGtCwa4v
16eiKvUrv7OBHHI1Gg2Gy1JOT9AsmOlt9SlevvNy9Z8x+A4PrQrm+A7kh+yDSGoi
qPruWLvPZYYikYvJvrhaxu8eMvtF3hTmZ+3BYJSWEJdF/lpwbB4szostICvb+JWM
Pg07CRwUVXUtoWvrN5/C0q0Jx+isCZICyPnoK/Fm4FH2eVwanINusFGpwytkrnEC
CaZJIQisyBok0QLSV0yWh13P3i2zicPztmjt1WK/JUkUqaJ526qd9AVf+uvs6h+R
7yau1V5xY130MvQiEwO/Lp0AVTd3E/doTbpFNwQJVGxsbhFLnH3eUilwgY58dApt
QW2zGCT7arPksiqBDADfGu1X7TRPM9Vp0aTxyoiww+u6zX+XORrgKt9l9+RVaisz
N2mQjJmvk4GUmjg0cBMgCrBo2xjBp2LL2fwD4jeiF/rE7DScjVxhIhRMQh9i+/Ln
QBvQX8hhU5lHh+fBk6jZJFuIbt851vSss4AZfDVm63tQVHphgRUqVMRZNv6DQUIn
DKmnW8WDXyF9L5SD2qNrYCnBgFZTxKmLqyuUpYLEPe4cwF7lxlhzEEYeg0R7iWh8
xKRAJgmwvDWgj2hspMEjJ0MCOUrJVpri4R9Cwvh8GEWl3tjQbIbYWND4FEw2eG6g
XVMydr1OU1HmW9NF5lR7Fr6sOSY7nVdHP2zG7v3I1ExynQErdqOjwut7z39D2qtb
+tquLnwcAzMoXd/oHxIPaw1RWm9QpgGnKLnBb8CBugvNaWerfcDJ/SlP5sowYViZ
rUxlalwLSJB5R5FbNJd/1C/jQQgVMSWHwDIKPp6+v5ydoT6zAWW4UwF0UfUKs0V+
KcEuU8V6xKgq/MtRobP4n+4jVNlEMLUCcC2CrSTbg4WSNUPchL40EWRA4L46oW9O
9sbEhCeX6jdqufgFdEIJeKn3wJ0sMfDwAYauYdIpu8NU/bAQYKJXsw6lbSgRadCc
PuKVzP57dPX43FudwLDhA4gxJ8Cdljrt6BL6VvETYle0otYcXyB2PbYpFoqG1cvm
SX5EvxgjEzDdqGfSOajoQYSNjXZjrqjQmoyoqoCf5MPyFdSz1HYM0kXWBzB6zWus
Fw9rVXl1A585mNWG/pYi514LYEEXg5VqcAxj5lLB1eNTyhIYcC3nEf7jg3IjK56p
cJRs9LbtHQyt0Aag/U1vJIrZVKKSF1fjcPYBwxJuy70GN4+cj0TbyvN5KDa0y42S
E6Q9GbwvxktPVFq1P16pyYpV8BaLy0SJjpROhGG8kxTQ+jcJpAksekvj4rncGnDm
o6Db/q748b7FC36f2zB/Y+zN/o3CkCmF/r266J29NgUqqj8sGgi+zg2nlUwMIM7S
V/OFG5Z/yqYCMWINYvGkNCsNdXvLL2GYK40Kj1brY9jlmne9s1VW9Av+P/1frSn/
F/DhLHaxLwwhOupGGA1NJGPkfZHw4HfJz582STH5/2WyOPH3u6SORJQliDe9vkMl
IX1qcRQ+51Pn681HWFoif2tY5ulnINkwpl1GQzqwu+O8H4sgDzrYMYPhn/cOFtM0
kY0gfbtq7RHw36+cTxi9qbTlayBDvNuhVQUtoAG0FLed3iJZ9/VoeiRre0gGSaIF
5q7+5z23awXR2aheIaB3FLiSWWAJ4/W8ERTDQzF8zjbr8GfjHIWF6cH6m6/CThc9
wgAi03ypGqVBIzDTfCyRlq7U7lNl6ELYklXXfSCMwp7EuKGjJN5jI+MueqL1touP
7f0EcNwuCH0tDnOFHGuOEW+X7kLH+hM4bE8NImpK1++9vrPbezBFkcBfAQmpBeXY
KZCyp3te4JdEI19VAKEqJLqTpboL7Ucfl+ERm1qcQ/Kl0vEkNYdqPtyYlHLTIway
V11PhPAvo66tweabarKMv/e4Lp1a4pCShqlJbj8b+D/uhQHDPNxFy1DM7VUXa1Il
zcZFXJBWnaEsGh/40TukAUDPfrPB8yGZNFqUmZCPT3StM/frqFUbOqLosBhfmtdj
PNSnQlKbmEF+hw/3LMKV6vS01CB7nEhrzjdET3UPE5I3nbQ2gY/QN6dLvPNM2L6R
37P+GFYhdkGnkZxb5q5tZqSTRsOIaeHGlJ74nmBdQ3jGy9QVEz9mLQcDjMoODwzm
Yry5Nr04AwH9mFriQ4+Cml9OYbfn9W1aIxpjLDOsmWc9o3dSDX5oTALvb+cLXc8Y
NombY/R9bp422l/5nu/FOXgkRZgXUp2zcqZnkZgHshGF/EieD9j+5fd5GwkcFs/T
bThuACS3iIQpaaT/4jg/l346/zdULj+XYq0qrzpfiHbpCxne4QpcM9mcXtfUaTzj
ZVsKTLI0fzIeW0Oo8m6KeojsBqXKrCdL3HRsYuqBjHawRIJPW/5/7UB3cQdgzQ1x
mf3vbIL0c20QhLezaRUcVUfFok068aaesBiIpT9pmGrrVtKzlPSzO9qJ1Hwo0SK8
WRGIFYH+OLHOE4YmnbKVl0zY7aQAfW25wb6/a/GPeZOdniRSqdWZ8Xh3JNYuOur+
A+oJP+bo9/biH43yBXieTdpa+CRj9Hq0rKkp4GdX6WmZXR9Zhm4PVBKJOUj0Idij
E1fqhDphcchQKqvzbmu65I9jfTtHWhxlOe4bH5xrdnTjlAVkWkPJGvIW3J/9XRIl
dIkUwGshIealBx0UQkPHnOAfslqFLRHQwCvFInkUnyEe56xxeMghF/4pWcOEZHHI
u5QzOn24ftV6bIXKCbzKgh1SptFBFBQQLLyTdNFJhZ0ACBqqq+SbfbsfldOLzlSY
2W0NAV+gn/YwPHoPTPtx+/19aCozuzbTvss01Y/HDsROVUg7o4kmnrCyk5az0TXq
xRjwMHFvnPIA4mO7AZevRxTgfHmrZ25zAME7522hgnakVL8uM6JodDB/aOr7bd5d
hFo/ASw0iCvMenHrj3wHLB9V72xyAr5imfmsNEnswnjveKUj4i4Hys2UYAAUuKfg
v87fYMgT2ITFWbo9AvTE1qagQzoPhvCzbg+zpI37OeKmaTnB0Z//scA+qfhqGYIU
5x2hjY7MLs4s0P2tA0DEG3tRs6QF27akTxk+H4APyQRDDlv7wSCqTg/96QJZ9r9b
U/Z25rvhDpnqbw5oUIa6Qr5Z60WTR4SIhkGSkyGAk6Ip6GXiOSPN4Kc82gnF1Tcv
HF0gLdAvQxx5oCDftmuVrTJVYyepbI5z4aMa/IDeNWE7ch+9y0MifUCxSWOWHJko
lkFknpcfLxmdi5sBjN0yED0dJ9xYan81w1+mbZNP2stFHGsb+1ehL0RdLsdRuBCb
OC2FGSGPnmcnsd9Fitwc98I06XNjaMupd3V2I7WA1il/eKgxykJkC6FEYO9DYzAy
2Pmna8nyBwRDkbOLAS9WrpuQMMcI+04/7+ohj4wRCmqntEIXbmUqWGjsr7CsJr6p
zpWZsf0JAO3FXex8XhzUJEn/JIcVf+tFenv3T6srrfg1y2hnleHkpnfu7llL3U+q
oRGvsl0nbkBrE9XId3CaC464L6Y0gto1FQrqA4O5f+1l00vfb7krpL/QBlF6CmCG
C9wNXYtDcarmxeuykwi90Ypb3Z+cbPxQsTbCXIvxuH4iZ/pIrbtZcLU24fKmUSBK
kFIWsPdYDkNN9X7pRBcJOYbp/CE+F91vuVEkSK6NHjnKiad30O+zJM5Ge88sYLWg
dhGCTWBGzmPW+cyDIl27UFi4cNsFygoRqafSXtrSirqwAMs1p1lr2e5HYwbN9XF3
ihiHxLOlw2qaWwNM82bFwMLehv611+l6MV+17Rg+MToLK2Bxb/5zQUjxoE+Xe4X0
9HmXvmLSNHVwZ/0cXUsCR4irjOmrLQw04cKqYLpVZ9gOcV6VNJfsG30IFrUobuBW
gPp6FxF4yWLZf/G/5M721z+L/feX8/S3gBxdr+8trhY4Txl22Ub1wfFXRqUUPHKv
tZ0i8xvvOR7VRvIznd6Xb7cmuWxZC/bh6+EV39GChtXb4M9TQNheogQqb89mshvF
rwr/f+2KZE8t53lcZYFaT1cYDLK03s7HWamTCXFZIy97TnQfeAFA5mdo3YjwWS/W
93SQvKrtIsnJWl8/Kqhxupy5TEL5Uxp+9urMsrc6IdLRRPovbefPlAwQYobUpDks
4gfLWuIwlyLDz6eXPmCR8DQPi/IPISjCOkGHbOAR+B5cokOXx4uyoyMcUB+kBF+T
n2f16T3gaz27LDt77LKitLpdU554VyJTAAEuOacd5FJs0eKHEGCFWI7+plPqHDt1
qMgjOF3h6WId3Jjjs6xPR9KK3byQpbtcAp4n4p6dIuZT15OEx2xVjb1imOMfV7f3
VpqMefvOvqwR5SuB08/moGrYVvsWabPcxdyzqfV+/VUNgGLSwDiehLjx/fNrXt1w
q3XF045It0Yi17SSL0B5c/YQO2jHLc71HvyLxD3T6wzK1S5jQEL34SYsD0DC0WQC
iJXpxDPE9chfBBkQnH9GE0VmjNVSgikIfm1VOy12wgrwzp83G5utPLv5GVNrW2/y
rXpFefMdQI90DXoZblgPqbxFN0lYCo7eszRZoqFFYEniHREZ0GMWkTh21iov6ICG
/IFbpy3x7JaA2XcSyxENgxEt8c4E6rXXnOIAfbVQnGEcgWTypg/Oimr8zdA7sEHF
X3wx6wA4fEmT19QwX5AGeDPJkLglvtY/oCYzZLcS73dnLsbTIMFFC77WeTnYeBDI
73BuVVz9SMC11rknMbmXr5ZcJb87axDoGJ8pe/hpWEe/Uy6NeaCMCEMqLbXgkoZz
VzPEtopnPqU/Cyumx2HCAmZtKyVZVsN2xifTG6hP488Hu1IJV9fKIWorSPEMYGZk
yr6dND3yfbuS7LYa79uUE901RPLnV0ZQVQRSHmTrBib3Nq86YfB3iK5kesGbR45f
ZrjYtdSdwQv71lIRgALpFIuxJxL8UkrUT8apUUOHW4NNGBG5LWoGTU/gapZI4Ntg
9z0HMjfRnRh1RcuIm+vDObuPP0s/IGcG6tdeXOdpiHBTtAH7nuxp38K2LwDOA6mU
bVPZFt8f4NBiPAARfUAFZKFDEZUr5b/uDWpZH12SewLFsRITKMXppq6hvVeK7IAI
iN2M0qXArllvThQJdHf9VEv3KHzpOIuKBUVFtciKsd995E0+QvbgfK92G0Re12hS
eNcjQPdLQZQlGEbzzBgADhV1LeBxVVVIXkX9EQXmuX/LYr4DbBKvjpxV5Tt5FfFF
XHOtbQ2g/IGYF27KzFNMGEU/csLfd9wgy9f/VMPR1IOJrRg1OibuAYCrteePw6CD
SceXbIycbwqVhEMFzgyb9mRxseleH1oy6X4kbbOJ3J8I/G0EOWs8eCnIA4i5U413
8GPktNsmXrUGsK4E8rWDT8SSb90eYILnOMOLkof917icnZsarMk4IL3uGObwDaDD
3/r/0UTLH8sHjGEE8xG6YPHYQvr7vxBjDBUIt6DTV4EPqGT5eeodExDx1IniNaXz
CyB0xFuhvvCu5uzU81UT58XOJlXqb0kg8JZ1EaKaHMoMnYvEGQ/1LGeC96FKD7+y
6JsWZKkDZntkvFK8jtBWaN/AvOEq5zYz9raGXzm0RBgAw9NSj46dnCIieVmqJyJd
umADyPlkVmkM31fWo+rLvRgz+JVynjk0eH/lRb1eC7VX543kfCcxAk3gRyL+3HhY
NyD4K00ae8vznwp+e+I7BmDOnHg75jDAGSq9aV+QSangvbNmZlKzLUD5+5Ypu2oS
AnlIirG++t8HQXvOT6iMHxpvsWQEIDJW2ugg+gvcloph1RDuETelQocvKfennGYL
Q4KBkBRqyY56U7ltJ/FEzKaIfBT8n44+k2cGZZaEh438iAuj/892qj5ydDNIx165
d5UDsKL/Q+xXCac2f4bpqcPIJkJ/3ZSJDhtlAYVqJIcVrYuqLsYsTiISMh4jXQTh
R+sbKf6gnczoUFiuYqixAAQN9bUU1JuUvjqmQo2B0X4++vcFFQMJGkAQfF9ctQDR
iO5YMnxSpm9QG1oIyExTtvWVhN/KtFYPzq9is8O3rsVO6Wpd2vPMDHR53S+Uy7aU
P5eVMghXEb1LaHubeowBOZyiUAWAzfrUxRE4XCp4Y5i0/hRKBfmSHWXxFouWf9MD
7zcQCrTqkweTizBQCtE4AUZgBVoecw1BjppQ24Tnz2zrE4KbaD2KEinrq00A5Suo
GOHbv2QuuKps9lXOc6QU6pyfkdmAoDxKzXSMbzL7GyboBK5BOXnsHE4BcB9PL7yu
TcV4aZy7LI8HONlz3JlMIIT9zREcFcxI4Gpf8+yZBDtz4UYWQdBfoPuKtgwTWtVb
HxJomKmMgGKcfvBxXIsb7aP+ZjSgJ/8TW0zjCPE3cmpQKXXMrN0mZw3HYkxlmMTj
bWKyoQwrp0kDj7jVqc1xBV43lsiyJFIHHtYN/xnM93xAH/VPtNi2jwiAfhcX/FKp
FOOL/Znoj3UZ0v4AAUao6ri23XU3bLGo25RCJWrAjL77FPSQhNYfe4oRREbFRts8
mh2r5da/lQRJi+YQZNWj6zeEYTFY8sRke75fEkl5f572R/R+3Y9PiUPQp3rPEaIg
Wte0IPOZ9LweaBKZH4EyFxby+Vu8oaQptVPPsiRvtEZojovMclmiRVA1ml0pOs55
DZwl14MTBdzcHIN3ln8zmLfRNtBq8233JZ17MUb9NSsXtmDRZy/ju2Raedvb5/o0
cgtgtL0n3OU3/NENGHsJ1E0GrueY9h4c7LK5uwV/GzN4N4J5GBGW1AHFwJmbzmdO
bXAvSdC1r2KKyIFcwhElbKUwnYWNhK2uPLbQtoribQT7FzoU/StigURNTck5aD1+
uJctr12jUw+k5uF0q8iM4PEuKaTVenNw36k4XdtzAuWALrXcU7uOWyJKjQQkAmpo
FpwoNeg1fAYhqdH4oRANMd+Lh+htPWTDHsahGw3N7/XK/gjCGlRr4Pb4of3ZTxdg
uE4G47yTqzLA64N/NUetV7o5EPvSwnNkTNIlCO42CvHyDHfCiqe+lW+NztXHzyO8
jzmNTyGJ8T9NxOQSg4opZrUV6kSop7mz32uUOCaPw+zI5T8F90lK9mHwfhTu5mVj
eaykUE7XS2v5LUOVhjON8viC4zflB8arP4sf+7KaggCjHezmYgFbzJ5n3/XDCpUw
3mQTADGKHHUhIoKLV/7Mu7fluGuYlChSqzmPjDDjzP1w2PEHebJRVe2SpIsXphcY
T+HPzTl0QeRnEImMEotTdGmOF5ok993stN2GQakc4/NTTGEQEv9P8jdj25MhS8Yl
S3X7qRfeNOrAvq6e7htU3mHGIFCkqNxJaZBhBEkIglm5khwCRZmmLdB/tmUTbDeq
yhCMlIiyZY54M168vJKWDqAQ0OQLTmwOMTqmIf+yEjmE4ePPSPSUPDGE1BrdgkRl
Zz5o5brAEXyNUNC3yL1BAxdShG9vkwsRVhdk+zoeIzlTiOy4xoGFaNSuvmXfukBV
SnomNgFTAPkFO1+x7vIcAreY7HzotD1fHizObv3KcRJD3zREYjMVYCl5Xu50WB6a
xC/Mu4ug4BISvN7an5XAcOALelTmrxvtCfA2ADSHlh3FXQCMxxeGfOWcesVSqhyP
VPhr1rNjZ3xzZ2nbnghQK9xJlI5/g3/l2BAkpuDhwbInXy5YG+f5ETW7yyxamXfQ
jyp/ua3vNeMmqVwSBpf/YStfMk4dAQVkzzJB9Pc2CA5p8xHT9QCNnI3baT6IMSqm
Jij1nLxgHJfv/ea4tFgsmgx+GmqfGqmk8al5iz3QuPY8RCgFW8MzQNihMNQiXd5P
G8+2hfFVyDzHDy7J+r8VFei5uaD38WEf3O4OBcHHeepzTlhTp0c1gwI4Bsz2qggG
joc6rEV+SYSX9Nn2d7DvM37wpBSDveznkFFa6qjVAiq4ZYbLJzjCdRkKiBCDy8SV
nMxH6ylIsr57zrCpLITBu0qG89Vtyt/GvS2XNXLsiJzbISR6b8QecayK9BEj/l1H
+MhGZ/xKeoSpnFDFk0VCd0q3y/dm73t8/zM2jUKM6l6miEdzW/PZogi8M418mGyL
nBFfvuKZMhN8XkFXI9KMvtX6Rm3dQI0myqELR59L9who3GsDn8uMgOA3dbBxFlvF
srxy6SQXtSbv6N9vZZvS7JxAl+q89rdcFQpdU5v3SRM1rBnepMSV9tfPSPWwc+31
aKBIf/9PDkJKEuyIVnN0r0n6n8azy1XP7eoy2yAoWQpawR2fT5ova0hYe8mwoRLe
UJn04OQPncblCDkeiYB7o+/Q4ya2aJv4lSYlaJS6TPeITSqzMv4SGM1L+zCwVbgc
vud2+o7+6kuhmuVLqJRgS7z2Vwq/bli3kcmQizHcij9sT8sloKA/5BAKcHuMnh7K
x+MQ/0FHiSPYpi1vWHG9GACB03uRt9RaRWyvqCX2I7K0/hTndGebRwd6hjS3+wM1
rkBi4UJ8WsG/guSg6KgxRCaiDuWrwnYxBoqlAyDl/8sp2p8jEOvcVtHie12M3tXR
JRCtNncFzjWBZ6I2cE2tvwX9C4WbRYuPIy6IyvgMqS7yBsOLE13bI5hpsUI0X66N
czJbYAgrqJY3jwZ+taW/D+hwhwRUo13zL4EyGqWreLw=
`protect END_PROTECTED
