`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jyKtdDt6gbUE112+A3uBny9T9HgdVQSmSQ/+pxxXvrrvBkheRbM0xQppAwl8JVV
A2pMNeK4CV+1gspdlcbNJM/wwIQ6xs17cgKUK8t/FbHAqMCbMYLTYbFNt2Ew0051
6QR+Z8WbUDYOqudVcxETmA67wpT3m8R8wJ6TIt2hAFB9S6ZN9YUQZh8n8MIqJbmL
YsbOjlSH0RzuoRg06gFACcucCSwxQoXMDSWQet9IJB8x/MJTL6C5f0sf+4ou1350
F4vfODe7hn/YkTBvbcW2ZHxMgDoLzwePbgAaD3USA1DRmM1jYrcqZUFM4iquYoDk
Q01E5UCCMdpvlUAirErpJ7vlJHkfvlKgSl2ReapQia1UZ+1IY+MjqFRTgiIHdYz9
XgHzhVwuo1qhktn6sLkGk6BWkgKAuQn0pNC6g85NhP135o3qhkXSoq/gB6WUceMC
65Px+4lbPnOhdE/XJUBdYZYyNet1G2my5j/kSAQSUfdZPkYDmuGMG52GoXJwBQ27
iLPzrf8qv1ExKR1Lo8f6+e5itgOVihcegp1if6/P7PI1QcajSGe5EQynd01/WKKE
YRKQB2V6htdav7GmYTAAtn4/acXnn0wqIdWrRVZLhBEKsS9fAE8fchqv3kC8jBZ+
F4YjKismy9bmLAwHntN79N6qLebGzFYqqnr0VoB+n1usCnFzB0j2/671QuJTfsGI
kBOc3jF9Ocw5nLt+YUgOYDJ03dxAvyXLMcLhbr0EVdwTwVgKGtjbX2xRt7M+v0Cz
HLkfoX7bVqa7diKYxqYZVFVcKZ/OM19NSET82IMBW3I6Xv6KLWrA0bleyFXtSHm5
yhPI+BqdfEVnsvFnG5z1n23qbOLi2minUx0Eq+xtNPD7uE1jGvCWTMhIMIWDeaG0
8n/06l4ZUU3K5zL+yCW0rLb97+jAN5rqmMj0KhWiyaGaJbECeOXIrPSuiHh6stwR
e9Yma14rXFFfbg6yCVHF+4ei7/M4QYBmImzUEhIK6yb8rwKJjYmcAftUNfKRZd49
SGgB7jdaYKkhEFtJWawlUnoTA/QKV/2sjFlQELUq4GRCebbj++b+ccuHrqxTRb3D
1f6+cimD0DLWbXAY+qb+HPB2MgIBMro36sJKgrHFDykaCIJFoCNguUcPoABhf7bZ
osqRl/GJQHcGDlKwjo2OXTyw5iEWJzg7Q0LXHY3zUQZ4pYaCdUKzuAVFJH2urkiF
nUCCBWff98ILHGQkl8NuXVCIOyGFyNm74Dhw05O8/712zMkcePw8UQvzEULEAotI
QnEcNJd1h5ZcnbfIutUDpRUGOIbptHTd8UoQIdvHk6L0ihs9nSlvZ9Que/dJFPC0
AZ4RkX4b1/aYprWRNdHQ9a0emhQLLLWIEyPG1OFUX7VFxnY5qZkTlE9ZDSkOQ8rQ
b3HAoYvcJ6OeSPjDXGo8nJH6TJmn3aojN8PQOzAHpy57Jn73w6TNHQ8pRaYJp+Jo
yqTvuzkb+h2JCCNfWFFN/oVT7qOe46JG4tDo6s80Imvd1cZbAVeeFnyEPt3n1lLu
WLusa0yFP9KUHrsqWNO3/mk0JznXl95d0XgwS3Ckuc/Ltv8fHOomLrauAYJVI3zN
62T82zvMvv0EEp6CK8YYVCcygbRkwFn8dxCvPP6ykoow12bt45rZp592FlOTRDSO
xHyFhcpoOt2QqqO42kC+6fr3RNooBvfcoAd8jcg7hCDIbiPcbNZc1FCCl0pSFXwT
GZKRdpDWKhy+IVr/yoPUj8jP+V3uGclaGPveKfb1/RMfO7EdM+uDIIgdzP2pMO7k
2FyUA2bDuSBzmfnE400QKvqnQlGo3tKgr9uenDdbLSsLdo8AOUI0yHuHRYmL/i1B
ZfcarJwaiT2Y91w1ogo9thEllFMxdfduE9ATg1qX7YsAz0p/ugSlBka49m55n8c4
s+WetdOSYSIHW6gDVm05UGckDVJebW5gv+99v//tksJwAChj0GaochBAKuTdV1k7
pRD0gWqLNUGc9BoFH4kpTz1e1ofsc/02dXY3UbitXzZ/qQ9XJXQkowCUKsgMK8OT
8piwKkkWa2zKmlPu0ogxWahFwpgc0GV3rdQKDXpFKM0g5c4DnTeKAfFXbvGTBjVE
BAgJhi6B8qkLGIZ3jrHImcWl26AtT6daGCfaJzMkUELGfZEfcWM2oNrAF1y07iLC
mR+y7TJO9G7S42MQt0PRnhfMBlGIOSp7ZQTRSNuLqdT+ul15Nymj2IgdSWTDzGQm
AoJYDagdp2Ou6ryW7w3yo4cmN6BKSDIA0Hh+CXy/doJHx9L2nDF+4kJ6fgHgyPm+
IzMSiVBbHwct0IOdpqdxi3cZZf7k9nFtxL7DGwPKM1nzm5os2G2Xx2bWbVljCTdK
LdHNEFFbttYO/1ynjqsgANI7HXVaCRI3v3Lu8MSBPunsIarqPk+vtzya/F9ZI5zS
vE82WWN3wAR1aKSt/893AXICXlGQW6+RTgbCyhd63mxH2VZepclrtodCyHs80WEi
+uEriZDRyDmQR0ttEpBdgywjcABt/yd2qJTZ+5TgB6jpTpICdDukaDyCK7SemHzW
rcVXVVudb3YZ75Xqp/63f4Wg0rcj6kpecWQ5NkZGNhrdCrHZOnMIdgE5TU7D5Fsp
fOZKdQc1AIe00cjQ3L0U1TZTW/+ZSOPs+iqQi9S8v3FeKo8ewjGnCVGqxG71FBe7
ZJcWdxBFbp/EgnNU+maanjZIQiHf+OcStYTsc5X5vaHqsXtaAVHB9VzUK9WmXfWO
4rxPavuxTHtPkkhmbdct3KseHRvRTEcKOs0fq7S1qbwQqZhh3Hy4Z0oVdav8IIV+
PlUeGbKsAEysoANq687EOnAn/72ase6V3sreHjPyAIhg2EFKWQw7A/f1PHO/JLTL
fh02knCxSJeoOUg7YRMrs+WZ3949DPW213n4lJ+kp5hB1Gn31YVCPAIsYIjTYmW0
p7IxGaNsiMH3u+1F65Bshq/Bu0OkePQTvkiSn89t4ndY9wCnjUgBXm2UIRRYiUE9
HCf/4qSgQ8PLv6JrHdsikszLzq51qUfRqq4EXHQENG4BbuOdkr/CVNrFJ2o9x3E1
Qfi870g90wIsC0KhUhOyWKklzmKDrDuwDte0fEtsS8u5MM9VltsNXwYZIOedjIkP
PjxU7aRL4cahIJvrmFB1gByeZ0Kz1YFNl/md8XCoLd9yrTrvzTlbyxdT/tZnXTi/
dePdWcedL8LX/Dtu0xqIFjI79+7mo4T3bQFa3etbtsc2Z3wfyUkreZYgLNPZrjZc
hPGxO0374KI+uiaTj1ZWbchyStFz0DYmaNEq9ZShKEEeWQpYheA8InJO4zPnOCOc
1lPhs/wyesmednTCN05kYi93rhTMFxPpB6RKsvBSClE0WifU6MAJGMS7R4u77l06
+TizcG8QIwNeKugkf71VC4yVFGR4Ql1+Fhclv95IGddc/lanNBY8w1IHW3YlE84k
WtxX+lcrkonuBMMEcp9Zyg59RbskBwK1JEcLHDIxmokePoJVT6WUY1aZ2nvbBdsl
GZvtFLt2sjRwZDTa4eEctoQPncKWZ7ZgA6ul7rNBnPE1+6sYzfMYfuBt2RnyPKHq
/+zanMzMhTW05CzX36Pa2y2EJdFv9KUalYwhiVh+7YNDDJkmdALvSETi4AGHFbNd
D4wrNOmUwJ1WV1gB7f39P9Qb53gmfXW/M/cYuMCy5DeKwZaRvV2PfgGE6y2/4j5V
LJnTR1TgtKMmjehFmj/Y6YpmuLBZWYbmHwRVLza6KFEkpucDmBLWQuwFcKkqTQSA
7mqDK+yPovas9R2BIC/YosYoaPglf6H/oKken57430GO0ZvnQvl2pWUPze5dtLL6
2DphWxKMej3ClJ5eFPz0i+6wPFWuG8ZdYUt4u9DQUKgcankC6LTPI9bSv2iJc7rt
H5Oh/ngUSOMiKiqzp8T6iACWmu5PfHzZAmLDsQuAMJUWcWWIQgp2gFM2o/o6n9qH
InBzrYAq/FFn2WJM/XZCYh9FZkEHIaHs9Gall4f/r9Tj5KJNiY+Q1xJmp6SswNjr
XBOUa/g/7SmdF10wXnp8336aK0z7Bh96Tek66OSG6YZHjPDST5NmKI4mAuTOft1z
wNK9hf0HCa4/ZhtrA8dGkBPPpaam+3e5w8luiKb+DpfspPwYLinDYuGMNAIqbnDr
44RJhdiDBAa/9301g+AyLpq4GA3Y84C/oaEDayYiiEKoNbjR3WOQ1QEojwShkvZ4
M5nfEyvJUm/SepkDt8KrW7skTcy4cwZhhphBlC3KdXiodGYVydyPv/puA65kxQLJ
Nq6tXuutWh9y5GXmWkNbGyy6bkFXAX/8nndw9F8WutmZKu61PeE6T7SX0VzHm6Yg
MZBQlS1YFSdNvdaG0r7w3e/1Mon1Pl9d5V1V+wm6ZFclqONrUxl6ICTeiuqin497
jrTD1cmCJFIc4e18+cjf++n7dvt7/UpnnrzfYIvgFQFlLYrzs6xvvVZRoL5IJE/V
8DrpTgXZIPdT3Wjvgqp1YsSr+X7zv6noSIldCDqzbk931g013TXv4PKG51Um79lc
y+ml0lv1l/iZcvdxays8fpQMawTxF/Yk3qYpIkRgstMXOb6pdbincmHA6Fqu4kRG
xs1RIZxWeFqfKSAoraf1eawVG5iCwHmvGgscfRhRXgQz7P2i5r1CYj6eXoAOenJu
e0SE3j77YEfeLaYMlYPp2oXxy9quPnelvHAuxvp8EYG/jXnxM3FMiV3GW2peCHAz
ZTz+FOZfn81cetYdNWha5FGkHnd+PbtES6S7+Byp/rkUo0gUEBhqUYPabd0Uv+7P
cuOJ7eexqr7Pj7pIqrKg7UbIcW626FBSzzYQmyPgcY/wp5aFrYN1sQRTN/sqys1n
8Z0q6l6muAojz0Fx6didP3yK6Xs26WrCfhLXaaxsy+Bjo9xDiW7faXMsppF9/P71
IdHJR04ui/7rV7crMm6OJ/StmRm12GZdJoni4XHsjlnu4RTz0JqyQVjFrR6tsEue
Th66HgC1wR42D1RtER9tW+O24axHJACgjq3wtDTYTsF/7nfnN+tOCKmR/ZJlLGgW
XkTAExJtA6Dzj56HHoKYbDnPCVdf1bTbj5a+eLqQdMLJXZmXbRoER9hLHIQXWHW+
ENff7ts4JsvMiHIqEclNamKPo28+zYrjwNIpLdWkn8bWMXcQUV+pIERGfH9ILfSw
tG5iRO+66a5BHZDj8gk0jQLZizJRs+wvC/ScEtomykastfBl8br6CSI4F3oquRik
Hez3xzP2cLM4tg0xdT1S4CnxGQIIsX+dhs5UZ1PctgL2JDFz0ECx/aIlouVheiuM
s1/cDFpautNtYN95FIF1duc8Y/T1dn8HNvTmXX4BT0WnXgsshYpMCkZDnmrZwuJp
Do7a59IHXnReW4qv55xWJ7ltbj7zjs+afpb1Ajc1NS7SR89Xk26VZxRMWJsaxAur
PQ3BT92nDTFx/ghgXgN5TEzC1IlxGAf65ZZ8X0CxDoEzR9NFyQuO08Vrwar0XpdQ
7nhohwNTlAti8zJ7RQJ6r3VBqcVpLFRHUh7RZPIcCBAzEUP53oOslzO/5cQZYUmW
/+JJh66nfoym2EKU4K0PY3WvhMgnt0Qc2KS19oPIUiaCBmMRCQ6pIS6OcbwyRUEK
lZXGIv3KfsQ5hGXxA0g4qhhZkyC6D6Y7vmvLskCocSQlmfgKoBK0yN40vHR/gKhy
VuC0ag33yKhQUce8nzfSVlMHBpmvtQhydXNUK62a+uOQ1NwpXDnvSVXUMtCET+yG
Yo94i/XEliOLXPRbgVoxlMH9Uk/3ZQm6YNZbpI/DT2/GITXGzmyzgC/LuyXHOlNZ
SDXhkKBRPs5Z3piGNs3lqmA3kLPYVZnVqXnI1FuRU0evHdc7uCxrUOdsvAF6lEb0
DTCbTqqBW6ozlv9BTEKEvz1A1AnkcB5mJYRr9XeiNDQdEK/h8vh8CtG7Q4AP0xJh
cNeAeUChaHJq9t0T5OLjYfH0IYeSFJp2LF+JWuB7vdnMjJrjeMjUbhXouZzUP1LH
csNE9Fc5VTV9j6RFykq9J8tiU+zFWzMy6vYIb99QuUL9f2lELxgiyOpKb5bmyWqh
QFsH/ArNdzUwO6iwXXuk/GosIA33QBCDMiHH7x1B1ZZJSdUE6i8pj7s8C1PsUM9p
9SR9CkAhQxDxKMTXZi/fo9whlfsHuDPepUBZpasejxhJh6LX32GaEf11DoAbL9B9
GwAxF//N9RkGaC7tEdp1Z6eNmSaXfip0Zr0retVVXhP2UvtzfzV53jUprRZIPhA8
QfiqxJYzHqNDo3jOj6hbmjAe4Ix0muyLSEf8Do6igLN2yRRteoZWALTD7ZbOpdVk
iUXhKP2Gxom4p/2tDn6JChv9qEyNBgXE0jbb39pdSgMdp6YQQRNQ1mDiA+o+/UZV
cQu3o4L/izBVEuZcHHlwVlQYUGpvhmsVyQwfRgxKe5ckegi37VMJe2bnsloOMWAn
jsPO3Jjdr0PqVMumJIZdBB19H9jY1b4MC88agkFSYKSVpr88OE1G7Pf9ESXUiHAP
f3ALPazAEEZPDO206S4gU6lnZzOx1Yptp/UvYUmUhYyfv8lP2P4ZWRFKn7zOfX8H
kUBbyMMkydUWkvMinNsLIPqi1RdjmB7gCVZns1RP0nCTd8o3/i4L2Jwvd5HfscbD
VlbdLl8wflo7VfxZNGKfUhNuk1ksn3bMsmZjEAR0sgGNBKrKr9uj+rpeyhS4eZa+
Fuh5n6Yfap9Vp/220fGxRJbvgND2o9k00hWiH5QY6fh6L1vLidcynCHCBRrYEcCo
PMmn8Idc44HAKR4nYqlDWyVJRQpp5SBDXNEv3B8HaZqzV55QGCrMMl6UX9+a3Er2
snBwNogd4Aovif0ap8wFQ6AV7MTMazFkRqLjOLu39iLERB9+RRgX776jJ8rPSWI8
sGDipAr4r9HiQiDxMkz/W6pLv4z99MG2GiA7xjQAguamc02MAdaqRIBCD/hRw7yc
DvSiYMKRcW+6KFpQZouuSB9oPQFeYFVfuDK8U2Wz791dL7jwE9jjWf1krc13ZFIC
P2IhbWdP4Z7fczBqyEgTX6KPjJ6uyUL0Ct9e1sseFWSDjPcmd7QjI+KJ6kdiz89A
GmQ+DvCEEDHF6JdAY7icoatHjPWcrEj8p0ThGteCW18qI5VgBOiHy9vfryUsC8V9
e2bEMABRds8fL1IvV9iF5lsOjMK3OTmcO0uACohywhaOQIdojo3SZxlUOtZxwnOc
jppPp+HD+n4IqXBUGtLXhTy7VvkQtwFxJwibxquOkL332gw6lJjecZ084kBK+PcF
IWckaFp7WLA2a2dfqkLI1+vU2fxwcyNWH7QyCZEcBfB65C1E3AdAxZIzHO1aCDgY
TqrjRSJYkxuZLztbmOL6G7WkVaOPh9/1DuKj/h+IB6Ge9nJtFsSgAeDKVOl4U4AP
ghIlwyfQhFOQVBG4/WFTpezKPUIxR3XQFBw6L2rCbzNaE3g44K5zmBt/yHZkstIp
ZwuCE4H9zsU7V8VrpZIlROx/ie/LoLsT9p0i3mHP5Prg2VLnDvq+x9O1W7JuuoGB
mAcotrxZ1nMS0OPa/JDULlh7F8VU/DuOQj5NRNqo/EfBqFhACQJwVfjhzGtcD+cZ
pwaBbz65D/jCsepj+DZpA6KEZga+GhCP0coGohjeasA7Hy1sbYpW0cKBb9ziQeIy
84HFLobofuO7jCeF157Oh3g6jso3nmdz4TPVQpS9I4g5MNo8ZvBd8bDosm23Tujp
Rr/bbimMdxY/RRXRUQ2k/7DMkRn7PrX9qPLpnNXwjrS/1xH6gtn2+xROJaLPydxv
1MEx6OWA8LMAG83YEC339hvCq44fBkPCof0xIEknoFDP9lnXSaL+RguRMKqODLJy
dZ3HEXc3AbCzO+t/gSHcHci7BJvLRpwTZnkMFEoty5QZDu2ZeOuDyr8DA40M36Bx
+dwccjh50Fjsc0ZE7MZPGahcOZvMYROgZlBTwcmSmPCUl8cg+35yyiemilxSzDoo
PGFbjCtcm5dh53IRWzU4lOmNaWNqbPPTRjMtxp5JKmUcUgOyC7ZUeTJEbIOScqii
Rih3sy+kj4KKKPrKLLEqZeChmZUgTkZDC0dYQl3/6IsmfOgYtIy/kJzpq/a/hE1o
v0gpNDZIGI2fsXr6xrE22y1iT8Qu1HcpXtYNzDJUlg0xbr9u6w9wfp9oW5GbgKRR
2GmMorkSgiByth4+3cDh4WMwJIQREWPukKpnTgH2MFBHplf43JTEZMQKbDiC5jRX
6n19pKCPFvWNIc4oa92Q1Rm1mDo5s0JVOSqqwWSrHyQ9A7NatybCYL10yjdO9BRr
Q0jOmFWmlALI/sJTbWr1BiABT77c/5Qw84p1niEd1ie7Sj/jucsFvgp/vz+aHMl6
L7UN9sqRUJjQTS0XldCDnb0Xr43p3cK0MjNY1rcaA7wz9bVmBdoi3Oh8XACobf1l
iNLACNtGtupboxJxWdLncqNaGZ9afNgq/OtY/KRZi6QP4LZ7EG5syBjuhTOKGrd7
m0snz7eLDBNv+N9o9J6PgTeKHmE4wDa+TC0Wg44vwJIHwK8yY2pT2XQwovp3TykC
eA0q8lsZMlw90WaqSsKmG+pU/dY1OO+CDkqh2exzy1oRdedTOdIz+azdDjb6td1O
tF9HcGTCzpao5UK/MgKJ1D4d7X19zdsdAdsLAcy4gMSIlwHgqoe9xpliLZnDypTT
qyIAe5B9V3YsDPrn1Ac3/dhj5NJaJO9Ix+hUeCcJqW2H3yWB/NytFCMGmJT1eZH1
+BE7WsoTiNTftsxZ9iLkEOjfYv7t9SIjH9C1vpIwt6MHYrpwwzPh9YriKklEx/6B
GR4B0gPg5wn21LtN0tB8GdJmldmiZOjAqAMUWOx8J3Zi3grLWt0EWFN1bNtOeVyT
JX8RuSXeQdq7wuZAtdB0PaImXa8Z0D2ZJdVrihfZTWUM1ZbX4U+gJNhlC1dVRSZa
W2Q/4UgnwsT51QhBPsoshlXaGs4so7LjpBs0lLR31Mj6stlGVCCEOKE/8Wy1JNT4
J4aWPBWcIVY190+6cO+eZldcxeycAzYBlTsae2/DdE/URzchxFvYJxQHoWb8QL9N
6ouR9QcORLwugWMu7Ibv3L7rSC/kW0ti9jlQ04PvghLtYlMt0AkRrAOcUqgsGeZD
fvn6pJx6ZGjxiG5Fg5D4hEMx+1Se1RjRevU6p3r3AYShnSh8dxicBidWSsh3JpbS
`protect END_PROTECTED
