`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GXb8Wlv5S0Nbwxzaj5JlUVQY/Orc51P+mTKK91zEUqnbyJao8oPYQp3QfjQQNE8
AjQISj28DXhYUPwiHkgmbjjP8mPTWgLrbd1Rmh5Q9vJ49OBRgfdcAFPf5dThFY/m
7if3uJbfotNRoIiL9bAY5R5TX+OcAuhIKHcSlGxar4aUjEJTaSd+zvyh4IXePj9c
sD6uGnjTH0dAiTYEh3lIGhm0xpW7yqagy8XtX/F9EHPHFHOzDcsWTMoUboLnsFc+
8wjpZ++inEnweKtr/hb3KzdsLK504JyVXAFI75FUx0XT0X3lJmOZ2jokVFrsfNWJ
+DfU/QlflDo3UO5DQwZmzYfbCw3kLvFOnHlSTYRdc6NJvpUHcwLrN0kw6FeEDmcS
utGIAZZvxKlr4To5lIKGMrFVJE+ZE28WIq9zCd7zPAEbWl9SopZoyVpNm30cXRsC
0gRnuzPgMVfiOiOvIYpcqtDeMrwQQcQcBx3EIJcs6P9r02KAXxSPfamjgyGkWCkv
C8ri6a/WygVYeg2d8Ji89jEBBI7BC/5IPMM/hy/3FpyzTWIucfL1jQyVsf71gMBL
SnOb8gL1fE29pHDFkWWh6cKKZs/AhQHNJr3kNlOLHPf5ITMtszkPuTpusBHwIKnE
eRIIT+uy0F0/Q6TkzPr0ecuGxKQ4fr85Nd7jutg3V1huY5Y3SrWh6vzPTVYktpRk
NQrb1d2UuN2VjDIZ/8B57TIRIi16HGU60SULnBLDZ4X0Da1zKZbNLftoe20OX5Y/
sUBcLK+EA4u4BAGDSnQJknpl5XJvd3S3m+tg1cZQGjI=
`protect END_PROTECTED
