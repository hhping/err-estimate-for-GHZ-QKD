`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kp+bXBoJwkWx5a/7cxCK8kfV6K+UIzOODoCSmxCrlcJ62X0JX2kEsVpVd66RQFvZ
W4cR/NkAWduM5Z9ekDYIx5eCGz3wr5euIGGx+WXXa2vB67iWwh3mpLaOS/gVlAiH
ouu6yZuWG6E1Gsx74RKLK+03PqdzL+oTZukeXqK2LU1SKMAsy7HhmOVlwvNOUoes
yRcjLx11ktq5ujmYsz3drWozprvsWBW3peIVX3KL/ASMZr4uP7mGfmNLmX2X9enl
ChjQxTY88Ny48tXN0j/pkMU89V1bzV++fiw+Gis2cBFQxUdd3K4j+l3PDJ//2XWM
/uieMg4/kQk1ucNlOJAEXzBFOVJKg4CIal2vsdH1faqBnQx3B64f+1KI4jIlGA3a
MIOcNWwUC+lrQQVEfDJKL/ahrCheglXspazzWY/bbeE5KGjEd+UM3EAvLV05se5U
mZRyVQH2wCXay0o+e5JwaUK1j+xo4UYgpuz8/e8nO9+t/64FnqfhOfAXdFYHP/+n
ZgpzfKpgQevv76zOy/FMYFM5iFLiSnF5ESwSLlYguXOaXfLahhXTebWw9fFQZ0wR
96rBAylQcIcemEH3pzMRWOEnBpi0BABNa0SX5XH4GTpFUS+BYeDCe4C/O9h9bUci
jZjqxrkcCrnSfeodHkcj2e4nEjZOgohGd1+NH4lfmmDJ2xJg4ijsMrfDaysO+vE/
kots1lgZGmFq9zh2zJPEYmCLMIpAzEXOlCiqYLDegxS6gttSX+DftMeyGt5Y8nuU
lHcDt3t/CFgSoD+0NbKwaHxKwZ2PIFwMP3Nubw7KUFjgqeehPp/VfXr5A0g19Qoy
rM/lWvPCS+usnVXsNY+jSrhySMY02RJ13Vvj8peMt6pWj7lDeXlJgZ5QBNYxsURi
dmcP+0HyGHYJmivGGMHqyMKvEoxcpq2AE42tOZXQ23uHmIaxaHX9liFSUmX3E2hN
mrE27jFG0Paouo+V7kZQSwrrAP83EebeGkgxjuGKwTxpckMJo162pok6fvSkmUoG
MRv4P+nIO3bVoKKbY0lIoFkyqe1PhS0fuz1J0uSfEWFLcrUJAuvX2PgBZT5GZTvr
yWUI9T9+Sr0OZtFkoqQKv/BoA6iDenWezMBjgYVnMF6JOW8Tz7G5yO7gb/NX9Mlc
bJc7zX2GYA56Ojn6CDpGR5q9x/JtfgbvrKpJh+S0UvnXLWIrm4QWKnmyRfKexA4v
f4PxdtNGVhYAn5+g0ef41w8tu5BW+OkD0rSh/jVxidnrAqcyYxEQsWG6SxEgVBSk
ONtJEelMK5L0J1DAW8rCbc4AjN9rv/zZEk/gk+LyuZO4RjaKQotF9Uai0tPxur3T
hVOOg5PJ/jYLs46iWfQElfOsF6pFmHyi7gmlTkPd5NOvXw/E9zx7oUKEZLQa7gBE
DUOLe/eAku0jUZY28zniHdDmcrd12TVi4YGbhT9uAdUALeJ2/C7GqOMZNvvK7dRW
5zplGWK4ksq6qaMv/DtNeOn+hgfyjZlrxCt1sFbhWhooVEpWBATQGiyTpJNS5ohr
6C3xyMw2JNC2Q1iDtyWtcz1euCNIZ1NALrGFAm6ks5wvT+JwMKDVKO2xVCKdl1bD
vq5VKZu1Y8PH/JMifdHwAFoqflzuvxokVI/5NmJgtKsNH4AoQs16kc2Z4uHKUaOV
tOa+5kRATdrh87VEuLay1QNOUkID0bsJpRxiNyaX9Y+cpfualG97RL4AA7xsWsXi
jj3se8Bjd7/dwfoyT+XdnouIq0gwBeU3C8jE0Ebt8mbMS0IBJLkmZusMIwvw+Tfa
QRbzrOFBoocmcSYeKv3E0dRcOnpkZvnspZq0gjSlluWCFun0rti7yogZd5ucAMo9
rYpceobasucyF6DzY5mfnXt8sMbFkZMd/KcqnVZRpWaZ2nCavuGkPJ2puUQk1hpc
nBRqyrh8DHZzR+fjfU0289Hg/Sa2oGoGPwMveBmzhs6TPvCv419v1zQ3DgUml59H
MbCSTwTahxHHIJ//1eJzDNdycVGSsFIqWNGOiTZNGvVyPVGZGUbXJkvQxFXc6P1T
OG7APSxz0sU+5hA4JmlW7xzlldD1VJ/7fRVKZ7lASGyghdPJVDDo//rIy2ejiA66
Ut2nBGHjHxmNr/IP+gjQr1OhYFePdf34FFFtJ6hN8wKdL+VKiWns7m3zK/LfJBHM
Q4DuKucTlMNL9ewsrsWO7rqG4plNQD2qO7NZxcTCu4i54z/zfbeuNLmKcGRJ9Rc9
d5Ug7RZtLOixGfR3W4ybyUl6vYpphSqt1rq+AhirlPACTOdhaUvIoP42k8EoC2Xs
x9zbjxFZCRBiUE5tQj4+b3iidmlozzU2/jfzf7xCJdKCKUbhXJucXR78Lsz3i/qW
KsOziOXdx2h4kbLs0QYlkF0joBAhd9d4+6o5Vi5/NdqjzV2TfezvlHcBQzSvV/EH
JpT3vIv0/xjmgWyrUacSBt9K9WNKc01p9aEyiGyix+LWc8gZFxWd86V7bKAEOybp
TWm6VRIvP62Efs8yEPIy07Oi8PWgfjIbO48CDGN25FUlBGO8/eX6jn7sBVmJ6FiT
e+vbgXeqP1Hkz0wsVh1H2mh+oigYeqSWe51g1ciHkbZhLK7e8DRuBYeTpo8lmjSm
T0CZo/0gQGPVT8bkmMSzXkVDnBKPKYbAT1t3va39zQ0EIYKQImD9kIBftKNEEmNU
7JxFLxFPcCs8s1nWfgKq2dVxLazFTU34tOf060rla7vCjwUD754FDILcucS9L/cN
Ris0dKDNTSy6Ms2EkHzQ1fRxJ+BtVyGqAkGiMYZ/BUUX57M5uL4JuCJOGpb+iI+L
z0XeJWXArVZ2Um1Gc2UugPhVgscyF6Oze5t37ihodXZmwEx0qJ2OvLLUtGNZ4z2f
hEaD5S7lylP0SsM1240IBcJa5nB3bFdLDQHz6VkELmz3C/rPt9cbXBiRxxe00HZB
M406jV7szw6D5anZfn3a+aHZ9e7m4YBRdz8lngifEzYP53YGCBlfQ4kvdal8skfA
6qqkIw6HsMIUafZrOnvr817Chy7pFq6M+VRwjm+EZRE=
`protect END_PROTECTED
