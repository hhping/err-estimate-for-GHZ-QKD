`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HUXOgzPxULvQ2F/TEpvCsOWZtsjerp9krz0tkVTX5y6XyNst3ejkgxC24wv9NJfU
P9RM6sS17mY9Fp5IEuaOh+pORN3alIzA2H9D+eQUX3R88bFnUs3SKOis+cs2Sb/Y
PhJZeSefeK784DFdg84kbQENsy7w9B59NyI9sKanOrboHesL9ZMQYU8QsbMZXpxC
NVZ2G9MenBuIDiGD9QrHXbAd6XApWTem+3qYnHcBIIqunwMmhMEoN38/eqppz/9h
DH4YPPjMboVPwjdqkYf/Wg37LJM0284F2F1iujEgjtddZNHz+CZMRsmh0kJVEQQJ
9gihNzSDnji2kuPtoHriC0/dF1/xdOX8OuZtHQPaE3JxjtrtqNTKR+xKqlnj9PWg
TbxFLKYKI3vWYK5DPtAwBwmF4txdENJHDK40Pj1P2X+sAOtINtFve29GynKwwwZ0
I/ixeP+qf7TZjunSwkg3ZNvoJshNOm1LXFJRDP0iNNrXVu2FcoYWlclnsrHja8B0
OGFvuUXZ/LxYibcgRu5eBAKcqbOdOPWfaLhpFBkHhhIWJq19kt92yIoz8wcGihzU
Z04tTekZbD6xcvdnkEz+0Q7dEl0PqR1DVU4+PrDbdnW4DjcA6LHCNRlD7ZjpxDGp
ESdCBg+MPHu4BOu/Bhz1E2AV6twsv6FO9uSOMeWIGXHyyoRCIZ5NkffxtTb9Yrvz
0ehvZ82Ci02b2bwKZ0oeXShDiHz2qlDbx8I/1G2o3PvujT0zV18i7oaBSTKcwK8Y
1RVvQyYNhorWDvDB5xQ1SOhoQxRWhBuqsRxBnTREM9CG/tiUUxzMdKNoqjKXtAHj
FGI8qPmxCMlRGPlWsImzcLwRcV7uXSf4vTSd6PfQMyiwOAkoviqLUgQWHGk+e9Qs
+uTIqC/vuW4VwTD0+aiLGDer5M6YigeC4/wCXywdcURg+lkSRXe1efuk36LYPGw2
007YvhxHZOtccIJt8a5JPw==
`protect END_PROTECTED
