`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfiilgIeKFdf33Lpk4BmPKZb0AMj8bKe16nWARq3KahET0ExzQ4kxlwg/tRmLaSn
ONxg9SHXH/PZbd/C2x334jumsvyYrsAehAo36MSu2YKY5IDnH3acSyOGB19EhPWO
FDp10D7p2oYvUO0NrervRD22vCt5vq2niuS3LqJ+nEQ7tMXrUAwg6KHILqAdkwY8
SWILE233WnIl1OCDIyfbX5roTMNUZ63pZNM/5Of+bYN/WaafkZwWv82UusaVSzcX
j2XVy5N3TavkKzh4Ge/vGongN4DJkGT8azz40QxOsHlCHnY4cMwKnzzbgD8kAcig
wEKuFj2ITaAzynQc3f18CFm+LmhS89IdEQ+uhmR4KosGqDR7BI/IgknRGyrPsRMf
0tLNsiDQGF+jAqfHsNfmCGUVXrWNoTIa4GZYz56oyyMNXFvmmN/OX+eODUJHgW/Q
oA/D9HKiyuHsBZagECgnWryKFg40PIzRIgU+/NmsxdM=
`protect END_PROTECTED
