`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRgHZN4zeuvFOoosmizht8u1LKaJ5GbxL2mT/WPGYKTxB8MgZNc3F+AgeKk6PtEj
+7vlk0vX1TmPYkYF3HEVe4EAASjlJujIvVyV2vHhqa5FFz2UTPMjWWHhKaM/COod
L2belrsvITPuh+u0JSluUwkHVEsfGM0D1ZEX0J+Tt2l1njAExf3KwZsHixxBxbZw
YoQMs+bSVZQujU2Ms1eu/ex3uyDTsF0riAa3qGC3XnV9y/Sr9JaV3/K7U2bcyvlV
V15WYqw4FfrhUAOOCSzSVl9EopJnLux7Odo7opdWOqU9FbTee+m83yNek9i9m9oJ
lY5aE2PxIeoVFP8D568YPD9vRp2H7B6IjX8689y2fbLbiCI5ngwwh9sfF9pHVYyk
oWg5yiaWKpqAcB120Xt4rI7tIJoOeeym5TAqQG3ySB8Bdm9ciIZNm1gMOP+5je7b
ns1QTFRtipheggrp8ONrYXgoSSGb1wHjiU2jTBWWSJPojfENfXCi9InybHZzYJXt
R599ASDrfhyz8zBOLL2gtGp5Nr6Z7mU9d0tEHMTznX+XIIe9PLX6yqtPAOfcOCRv
d/ypQDhLj/jsUf/nrtjGX1/fpYD6ovyrkC863OjI3YgKBcSqhejwK3wZjlmg89Hu
zA7LCjzY8FyhIqNLmxybbOHT3RMPcygnNGH/F2v5xQOxaOOAr5eu6YMiUKhmdepX
vDBIcn2vCdhhe4imZkc6magSy6sYnf9GIoS5TcjHTbd9jJJELcuDNobSkFntavJp
IpDPbR/tAGZhk9LPLLv540cEycri7sKdEvH+p22uWKIz/UuKZz/aMh8wUdNOBYE4
ppS99zpCUwtt4embkaoEeAUpLpqHGQoGBtOEMoTTxkV1xI6myqX7sMpJSMmNCw2o
fVBQrR3UnI7m8yxjvHw5pw==
`protect END_PROTECTED
