`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uwC7fBoYuuLYRWgYVc42lYcLo4aWpPcizcredOqkn4ZlBwz7H1K9z08AzA+iQ8VC
/4Q/+Wz0hcVqirSU4Hns2Z7jR7ol50Ts9cc2dVBPB6fBGkM6NZDQ0w+fvMuuS8Gm
sbRDxyICFgji/CJieT9J+CxfqokWQC0XXVgaef4HOxWkEtbU+wthR/o/MXd+WXOJ
5sYtYlYQluSAXcvS3oIlux8mAr+ScpvFaeuXZ3+W3+MaZoM4AAO4Td8oMqOrG5Vh
Z3uTm0UGxmEygghhdAw1Po/kMHX2mDg9wlSc7FWelOGyydmD8pXFY5amIbaGijz2
Gmq/574oUyajvGf421IOB2tu4xYw0VWqDLJ7zjr9x3u6wnO6aO0ILTozwwQ1MvPc
eK7OJ1wvQXaZdzS7H4a90AR7hNKzMSq8wS5ZBzhqyRwdWW/a4xQcBvL88Y2XU7QQ
INtCcQ6gL2QC8M073jQBSKP9xIodCnpS2j9NP5+AMMZfTKbeF8FBGyaRvwhLeJBW
oCumGnqiq/IhDvHuMWWUjFlnE2ge1+EvqsC2oL1QT9ewmdzOUwOD9+nnQ5LMW/yc
U80Wxzdp/U3y0NYZR3iUZtN/do4eOjvR2qdwlk6W7HFyPKx370j9xvSLBe4K11Op
AezkH1JHX4n2iAu7E3UcAGYRgVPBD6HICFLVXwih6T3pRcqFQ6A9pVbiqa45CkJx
hfzFp4KHWThPhYJGOX+JS/49vGoGuZM+d8wa1mgKN5oPE98bls9VEHqnKi5AosNH
6oq58Pe5Tgn7CEKBLoc03cAEpPRPauD6O6N5sfscyZqlWQsGAKcv4GC0A1zOOutI
ePeGNC2pudQLBRF8xk7EsG5ZwMvpqXveMPgO3rXxzXo=
`protect END_PROTECTED
