
module log2_fun (
	a,
	areset,
	clk,
	en,
	q);	

	input	[25:0]	a;
	input		areset;
	input		clk;
	input	[0:0]	en;
	output	[25:0]	q;
endmodule
