`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSPu0d6JEX4l49amQ7hgabmLW9Lt0U7O+2gpBAcbpCviroV5ZHXY7SS5LONJ5YxW
YmZOegefs3wOAYKjF4UGq5Gee267c+8yix97ktUSmqQMuVLM6PQPDnMvr9hjnGQp
m1YsHIfHrS/ihi1+upsKc3IduRUvlUnuroveluNsnKRSPyJQupojdm+U7DY4+sVl
3RvA9lJlEnQV58dSZG6vNAamHOPL+FU337krhd2+Weq4D5f3/ALG8xeq7s/DEx3T
UCtorarTkNj1ORzvXu6hhax+p7gKjVWkcGpdsJYaEkYx1LSEgJiNqxQ+l1/CLs/m
2PDjm9oSncdGHhGN80hcvz0XMvtGRRKVJDARoBPAAOcX67GSPy+lU54iPqtJ+xBa
iGCbFfAinxrUAe9iN/MUSxD0E4hUJamDWOE6rF4ifLUuK2vgGRyrInjkhO76tLPq
Is173aZwEIpsDgB4kuZsOnBiHUXnmzKTJSJteaZrwUXWuFWyMV9m018J46ieyDs9
y0cRws0SYlwbL+C6fEuPrFHJFObPCZ40/aTf+ZHEH/r8kPivkK8fd0JK/aoPeUvA
TThH8cnzZ3uPTYip6U7SUU5WdCOozpXkehixP4DBWzlSdsCnqQRw+nHdagb+/XA8
GZ2it8Oo22QcbFqqdZLwe5EfAvNyIU0m33bz0meCWZAMyqB+DPhBwUiFnn4jj85S
vd/MC2Aki7iJ3v3JvMEM4thNStMLujkLQsX0bgmBQYHcIijTFzYj7JJaeK/w+y4u
3cJP79raPSxWmlrqovBFkDjBOLmQAG1J4+AalPWSiq0IaKSvxubE3gxP5ehY/Sso
v+Dtd/RQvAvF0TBYHSo7n+5cSiPuLyaB1nnZbBFrxtryB2jUH4MtgXs4OhuA9puG
i6eyzBdvvYcNoTm8ZIMbLaIGo0cQO1SHlWF57IgsEvBlALwHBeUontO8G2eGEpNy
WdXwmlTSBUwI2yVpPtOf6ZpeFVPJ3PgZeFx4AQmFnLV2UUaOeJVAHqoCyJfLUz42
W8enSZzDrqmC+FSr9KWUw4T88MNWL2i6SuN6MNxsP+cl5U8nBcdpYUhgSYlTFJWG
eU8T/vBWCtScrK1MVy8MDbrL0fwmjxq6IDcVuFgatn7atn4sRc+pymUcB8ACz34e
tMi+Ph1TtQljgKf+6ZYrQX2KLSO6xClybtILQSukWZWi9XT7yKqLzIMxGjO277vW
Q0j16d+QwpjHcpBvCSTwOLL+9fNW6chjuGb7L5OOlpiDwzwor3m37fYArQld3Xmg
QNm+qnnL2gZz8DtRYJH1/813yE2bUdA18CVx0K7iJxF3R8LITYKAcb27xZLmf1Vy
9exJI9nGQVqYceNlR04F8R8zaxwL3KIL6cMq+lW/mdwlDYitZnQedjddRI4HvpZJ
MK2qroMlcmKt461R+ydSd/0vUacJh8t443La6qt7WzEaVIuZuBly+n/gNw1TRNB9
bLBmTyrvHEPuYgeas5sEsyHS5q1YJA3aq/k1120v5TIndZegx/MbJEh68tBeeJl0
eCreA1et/BY6DcgA7b93McAyZm37yksP1zv/bP/jjox9+9bzRPybwwfM7mG2JPu2
DtYFHR1hSZ9OYVxLgpR64i8Nz9glm7DvTDCJ0Sm35QMKsOZMXu+1hlBgrOzUgiH5
Vj67OrSZBcXXA1Ue2PY0uArFx2t1uRws0y0NHscCnwGYXGyHpUlRz2k6aDKV8Je4
cosRjBB5mxWMToA5FISyLUaK33pd3FdDbeT1/EN2UX3DtYjwegbUgitmNgHgrDxS
4Su2YrlIM54S7aDSF9y4eVhbkbDv5ts8sDW8q734Z0qF5FvBU0vMAHLNW6AQO6Ps
hJYT2jOhOJM0lwNaOEyDWnL8B8q4y7ufbwrMRGHg/8g=
`protect END_PROTECTED
