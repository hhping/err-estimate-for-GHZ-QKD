`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCx49XrF9EzGK+Ye0CCqIgF6fgVA9YmFJtyJ2IIynDuVwtF0WOBVcHUnG5ZEmisf
3pPCe958YbOIjeah/x1vYxTBKJHKVNdSmAY01YOl/U6WmdN+N1gY4TOqNJ51HSxf
YkIUmt9W3CgLYVkDTbwtYo1A/NiQfQhHSQZZGBBF0ZR/jT7r7XR3ejRBTyHd0Wdo
Lb+m+c9JU+cQr+z4a0K1HzV0J7cz75Ms7xXMq/is/F3YNhf3kWlqf9mCKgVcOVnP
5+SkKOLv1add51M0YyA3CracJ400w7/atiSFRmeyyuWaMxvCh/1Snnqy5kFqO5bs
M6N+xXSray7OgjbaM9sPBidu9my5/cKYMSAMLyWMzl/npXlv4oBZkAG6alT1OxRw
R7r2D/9yy11D8ZwBBFwNS+IkS811RRYqs8jFbEHknMCGutLxurwMErMIYaCKR+ad
PIPqkbFxt7DQY6HUEzSlVSYCzBumfu/mWrFlhKUJ/9j/JZaezUnRNAZXR2/tt7N8
parFWPZXr3+2NHYf5XWrOnGP/KA7VRxhj0d7fw6aJTn5khx+muGYk1kin48aYfow
sTf50a66LIgAaKJFlOxrfIAZxwVAprpEzPW7y6NE6hVTxKOz6L9lHfSAKBGwOLHj
7WwtofHhZ9Q21T13NOuH4VQhPpQAk5yhY/zHz+vh7pTu9v/Eo0MoC32AImVwdWGY
XFrPELafel73HHp7qqUrmC7t560yTFNinVO1wGMzUT8tLqaPDfkE8T+HhFWybTjV
TL9VRoFuOFoAEXgj7j4lS4FPHCRox9qmtDE4t2a9qNI=
`protect END_PROTECTED
