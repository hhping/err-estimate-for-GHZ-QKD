library verilog;
use verilog.vl_types.all;
entity twentynm_cmu_fpll is
    generic(
        enable_debug_info: string  := "true";
        analog_mode     : string  := "user_custom";
        bandwidth_range_high: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        bandwidth_range_low: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        bonding         : string  := "pll_bonding";
        bw_sel          : string  := "auto";
        cgb_div         : integer := 1;
        compensation_mode: string  := "direct";
        datarate        : string  := "0 bps";
        duty_cycle_0    : integer := 50;
        duty_cycle_1    : integer := 50;
        duty_cycle_2    : integer := 50;
        duty_cycle_3    : integer := 50;
        enable_idle_fpll_support: string  := "idle_none";
        f_max_band_0    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_1    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_2    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_3    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_4    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_5    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_6    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_7    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_8    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_band_9    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_div_two_bypass: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_pfd       : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_pfd_bonded: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_pfd_fractional: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        f_max_pfd_integer: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_vco       : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_vco_fractional: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        f_min_band_0    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_1    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_2    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_3    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_4    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_5    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_6    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_7    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_8    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_band_9    : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_pfd       : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_min_vco       : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_out_c0        : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_out_c0_hz     : string  := "0 hz";
        f_out_c1        : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_out_c1_hz     : string  := "0 hz";
        f_out_c2        : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_out_c2_hz     : string  := "0 hz";
        f_out_c3        : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_out_c3_hz     : string  := "0 hz";
        feedback        : string  := "normal";
        fpll_cal_test_sel: string  := "sel_cal_out_7_to_0";
        fpll_cas_out_enable: string  := "fpll_cas_out_disable";
        fpll_hclk_out_enable: string  := "fpll_hclk_out_disable";
        fpll_iqtxrxclk_out_enable: string  := "fpll_iqtxrxclk_out_disable";
        hssi_output_clock_frequency: string  := "0 ps";
        initial_settings: string  := "true";
        input_tolerance : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        is_cascaded_pll : string  := "false";
        is_otn          : string  := "false";
        is_pa_core      : string  := "false";
        is_sdi          : string  := "false";
        l_counter       : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        m_counter       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        m_counter_c0    : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        m_counter_c1    : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        m_counter_c2    : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        m_counter_c3    : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        max_fractional_percentage: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        min_fractional_percentage: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        n_counter       : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        out_freq        : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        out_freq_hz     : string  := "0 hz";
        output_clock_frequency_0: string  := "0 ps";
        output_clock_frequency_1: string  := "0 ps";
        output_clock_frequency_2: string  := "0 ps";
        output_clock_frequency_3: string  := "0 ps";
        output_tolerance: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pfd_freq        : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        phase_shift_0   : string  := "0 ps";
        phase_shift_1   : string  := "0 ps";
        phase_shift_2   : string  := "0 ps";
        phase_shift_3   : string  := "0 ps";
        pll_atb         : string  := "atb_selectdisable";
        pll_bw_mode     : string  := "low_bw";
        pll_c0_pllcout_enable: string  := "false";
        pll_c1_pllcout_enable: string  := "false";
        pll_c2_pllcout_enable: string  := "false";
        pll_c3_pllcout_enable: string  := "false";
        pll_c_counter_0 : integer := 1;
        pll_c_counter_0_coarse_dly: string  := "0 ps";
        pll_c_counter_0_fine_dly: string  := "0 ps";
        pll_c_counter_0_in_src: string  := "m_cnt_in_src_test_clk";
        pll_c_counter_0_min_tco_enable: string  := "true";
        pll_c_counter_0_ph_mux_prst: integer := 0;
        pll_c_counter_0_prst: integer := 1;
        pll_c_counter_1 : integer := 1;
        pll_c_counter_1_coarse_dly: string  := "0 ps";
        pll_c_counter_1_fine_dly: string  := "0 ps";
        pll_c_counter_1_in_src: string  := "m_cnt_in_src_test_clk";
        pll_c_counter_1_min_tco_enable: string  := "true";
        pll_c_counter_1_ph_mux_prst: integer := 0;
        pll_c_counter_1_prst: integer := 1;
        pll_c_counter_2 : integer := 1;
        pll_c_counter_2_coarse_dly: string  := "0 ps";
        pll_c_counter_2_fine_dly: string  := "0 ps";
        pll_c_counter_2_in_src: string  := "m_cnt_in_src_test_clk";
        pll_c_counter_2_min_tco_enable: string  := "true";
        pll_c_counter_2_ph_mux_prst: integer := 0;
        pll_c_counter_2_prst: integer := 1;
        pll_c_counter_3 : integer := 1;
        pll_c_counter_3_coarse_dly: string  := "0 ps";
        pll_c_counter_3_fine_dly: string  := "0 ps";
        pll_c_counter_3_in_src: string  := "m_cnt_in_src_test_clk";
        pll_c_counter_3_min_tco_enable: string  := "true";
        pll_c_counter_3_ph_mux_prst: integer := 0;
        pll_c_counter_3_prst: integer := 1;
        pll_cal_status  : string  := "true";
        pll_calibration : string  := "false";
        pll_cmp_buf_dly : string  := "0 ps";
        pll_cmu_rstn_value: string  := "true";
        pll_core_cali_ref_off: string  := "true";
        pll_core_cali_vco_off: string  := "true";
        pll_core_vccdreg_fb: string  := "vreg_fb0";
        pll_core_vccdreg_fw: string  := "vreg_fw0";
        pll_core_vreg0_atbsel: string  := "atb_disabled";
        pll_core_vreg1_atbsel: string  := "atb_disabled1";
        pll_cp_compensation: string  := "true";
        pll_cp_current_setting: string  := "cp_current_setting0";
        pll_cp_lf_3rd_pole_freq: string  := "lf_3rd_pole_setting0";
        pll_cp_lf_order : string  := "lf_2nd_order";
        pll_cp_testmode : string  := "cp_normal";
        pll_ctrl_override_setting: string  := "true";
        pll_ctrl_plniotri_override: string  := "false";
        pll_device_variant: string  := "device1";
        pll_dprio_base_addr: integer := 256;
        pll_dprio_broadcast_en: string  := "false";
        pll_dprio_clk_vreg_boost: string  := "clk_fpll_vreg_no_voltage_boost";
        pll_dprio_cvp_inter_sel: string  := "true";
        pll_dprio_force_inter_sel: string  := "false";
        pll_dprio_fpll_vreg1_boost: string  := "fpll_vreg1_no_voltage_boost";
        pll_dprio_fpll_vreg_boost: string  := "fpll_vreg_no_voltage_boost";
        pll_dprio_power_iso_en: string  := "true";
        pll_dprio_status_select: string  := "dprio_normal_status";
        pll_dsm_ecn_bypass: string  := "false";
        pll_dsm_ecn_test_en: string  := "false";
        pll_dsm_fractional_division: integer := 0;
        pll_dsm_fractional_value_ready: string  := "pll_k_ready";
        pll_dsm_mode    : string  := "dsm_mode_integer";
        pll_dsm_out_sel : string  := "pll_dsm_disable";
        pll_enable      : string  := "false";
        pll_extra_csr   : integer := 0;
        pll_fbclk_mux_1 : string  := "pll_fbclk_mux_1_glb";
        pll_fbclk_mux_2 : string  := "pll_fbclk_mux_2_fb_1";
        pll_iqclk_mux_sel: string  := "power_down";
        pll_l_counter   : integer := 1;
        pll_l_counter_bypass: string  := "false";
        pll_l_counter_enable: string  := "true";
        pll_lf_cbig     : string  := "lf_cbig_setting0";
        pll_lf_resistance: string  := "lf_res_setting0";
        pll_lf_ripplecap: string  := "lf_ripple_enabled_0";
        pll_lock_fltr_cfg: integer := 1;
        pll_lock_fltr_test: string  := "pll_lock_fltr_nrm";
        pll_lpf_rstn_value: string  := "lpf_normal";
        pll_m_counter   : integer := 1;
        pll_m_counter_coarse_dly: string  := "0 ps";
        pll_m_counter_fine_dly: string  := "0 ps";
        pll_m_counter_in_src: string  := "m_cnt_in_src_test_clk";
        pll_m_counter_min_tco_enable: string  := "true";
        pll_m_counter_ph_mux_prst: integer := 0;
        pll_m_counter_prst: integer := 1;
        pll_n_counter   : integer := 1;
        pll_n_counter_coarse_dly: string  := "0 ps";
        pll_n_counter_fine_dly: string  := "0 ps";
        pll_nreset_invert: string  := "false";
        pll_op_mode     : string  := "false";
        pll_optimal     : string  := "true";
        pll_powerdown_mode: string  := "false";
        pll_ppm_clk0_src: string  := "ppm_clk0_vss";
        pll_ppm_clk1_src: string  := "ppm_clk1_vss";
        pll_ref_buf_dly : string  := "0 ps";
        pll_rstn_override: string  := "false";
        pll_self_reset  : string  := "false";
        pll_sup_mode    : string  := "user_mode";
        pll_tclk_mux_en : string  := "false";
        pll_tclk_sel    : string  := "pll_tclk_m_src";
        pll_test_enable : string  := "false";
        pll_unlock_fltr_cfg: integer := 0;
        pll_vccr_pd_en  : string  := "false";
        pll_vco_freq_band_0: string  := "pll_freq_band0";
        pll_vco_freq_band_0_dyn_high_bits: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        pll_vco_freq_band_0_dyn_low_bits: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        pll_vco_freq_band_0_fix: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        pll_vco_freq_band_0_fix_high: string  := "pll_vco_freq_band_0_fix_high_0";
        pll_vco_freq_band_1: string  := "pll_freq_band0_1";
        pll_vco_freq_band_1_dyn_high_bits: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        pll_vco_freq_band_1_dyn_low_bits: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        pll_vco_freq_band_1_fix: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        pll_vco_freq_band_1_fix_high: string  := "pll_vco_freq_band_1_fix_high_0";
        pll_vco_ph0_en  : string  := "false";
        pll_vco_ph0_value: string  := "pll_vco_ph0_vss";
        pll_vco_ph1_en  : string  := "false";
        pll_vco_ph1_value: string  := "pll_vco_ph1_vss";
        pll_vco_ph2_en  : string  := "false";
        pll_vco_ph2_value: string  := "pll_vco_ph2_vss";
        pll_vco_ph3_en  : string  := "false";
        pll_vco_ph3_value: string  := "pll_vco_ph3_vss";
        pm_speed_grade  : string  := "e2";
        pma_width       : integer := 8;
        power_mode      : string  := "low_power";
        power_rail_et   : integer := 0;
        primary_use     : string  := "tx";
        prot_mode       : string  := "basic_tx";
        reference_clock_frequency: string  := "0 ps";
        reference_clock_frequency_scratch: string  := "0 hz";
        set_fpll_input_freq_range: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        side            : string  := "side_unknown";
        silicon_rev     : string  := "20nm5es";
        top_or_bottom   : string  := "tb_unknown";
        vco_freq        : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        vco_freq_hz     : string  := "0 hz";
        vco_frequency   : string  := "0 ps";
        xpm_cmu_fpll_core_cal_vco_count_length: string  := "sel_8b_count";
        xpm_cmu_fpll_core_fpll_refclk_source: string  := "normal_refclk";
        xpm_cmu_fpll_core_fpll_vco_div_by_2_sel: string  := "bypass_divide_by_2";
        xpm_cmu_fpll_core_pfd_delay_compensation: string  := "normal_delay";
        xpm_cmu_fpll_core_pfd_pulse_width: string  := "pulse_width_setting0";
        xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost: string  := "normal_setting"
    );
    port(
        clk0bad_in      : in     vl_logic;
        clk1bad_in      : in     vl_logic;
        cnt_sel         : in     vl_logic_vector(3 downto 0);
        core_refclk     : in     vl_logic;
        csr_bufin       : in     vl_logic;
        csr_clk         : in     vl_logic;
        csr_en          : in     vl_logic;
        csr_en_dly      : in     vl_logic;
        csr_in          : in     vl_logic;
        avmmclk         : in     vl_logic;
        avmmrstn        : in     vl_logic;
        dps_rst_n       : in     vl_logic;
        extswitch_buf   : in     vl_logic;
        fbclk_in        : in     vl_logic;
        fpll_ppm_clk    : in     vl_logic_vector(1 downto 0);
        iqtxrxclk       : in     vl_logic_vector(5 downto 0);
        lc_to_fpll_refclk: in     vl_logic;
        mdio_dis        : in     vl_logic;
        nfrzdrv         : in     vl_logic;
        nrpi_freeze     : in     vl_logic;
        num_phase_shifts: in     vl_logic_vector(2 downto 0);
        pfden           : in     vl_logic;
        phase_en        : in     vl_logic;
        pllclksel       : in     vl_logic;
        pma_atpg_los_en_n: in     vl_logic;
        pma_csr_test_dis: in     vl_logic;
        avmmread        : in     vl_logic;
        refclk          : in     vl_logic;
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        rst_n           : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        scan_shift_n    : in     vl_logic;
        up_dn           : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        block_select    : out    vl_logic;
        clk0            : out    vl_logic;
        clk0bad         : out    vl_logic;
        clk180          : out    vl_logic;
        clk1bad         : out    vl_logic;
        clklow          : out    vl_logic;
        csr_bufout      : out    vl_logic;
        csr_out         : out    vl_logic;
        fbclk_out       : out    vl_logic;
        clk_sel_override: out    vl_logic;
        clk_sel_override_value: out    vl_logic;
        fref            : out    vl_logic;
        hclk_out        : out    vl_logic;
        iqtxrxclk_out   : out    vl_logic;
        lock            : out    vl_logic;
        phase_done      : out    vl_logic;
        pll_cascade_out : out    vl_logic;
        outclk          : out    vl_logic_vector(3 downto 0);
        ppm_clk         : out    vl_logic_vector(1 downto 0);
        avmmreaddata    : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of analog_mode : constant is 1;
    attribute mti_svvh_generic_type of bandwidth_range_high : constant is 1;
    attribute mti_svvh_generic_type of bandwidth_range_low : constant is 1;
    attribute mti_svvh_generic_type of bonding : constant is 1;
    attribute mti_svvh_generic_type of bw_sel : constant is 1;
    attribute mti_svvh_generic_type of cgb_div : constant is 1;
    attribute mti_svvh_generic_type of compensation_mode : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_0 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_1 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_2 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_3 : constant is 1;
    attribute mti_svvh_generic_type of enable_idle_fpll_support : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_0 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_1 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_2 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_3 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_4 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_5 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_6 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_7 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_8 : constant is 1;
    attribute mti_svvh_generic_type of f_max_band_9 : constant is 1;
    attribute mti_svvh_generic_type of f_max_div_two_bypass : constant is 1;
    attribute mti_svvh_generic_type of f_max_pfd : constant is 1;
    attribute mti_svvh_generic_type of f_max_pfd_bonded : constant is 1;
    attribute mti_svvh_generic_type of f_max_pfd_fractional : constant is 1;
    attribute mti_svvh_generic_type of f_max_pfd_integer : constant is 1;
    attribute mti_svvh_generic_type of f_max_vco : constant is 1;
    attribute mti_svvh_generic_type of f_max_vco_fractional : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_0 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_1 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_2 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_3 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_4 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_5 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_6 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_7 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_8 : constant is 1;
    attribute mti_svvh_generic_type of f_min_band_9 : constant is 1;
    attribute mti_svvh_generic_type of f_min_pfd : constant is 1;
    attribute mti_svvh_generic_type of f_min_vco : constant is 1;
    attribute mti_svvh_generic_type of f_out_c0 : constant is 1;
    attribute mti_svvh_generic_type of f_out_c0_hz : constant is 1;
    attribute mti_svvh_generic_type of f_out_c1 : constant is 1;
    attribute mti_svvh_generic_type of f_out_c1_hz : constant is 1;
    attribute mti_svvh_generic_type of f_out_c2 : constant is 1;
    attribute mti_svvh_generic_type of f_out_c2_hz : constant is 1;
    attribute mti_svvh_generic_type of f_out_c3 : constant is 1;
    attribute mti_svvh_generic_type of f_out_c3_hz : constant is 1;
    attribute mti_svvh_generic_type of feedback : constant is 1;
    attribute mti_svvh_generic_type of fpll_cal_test_sel : constant is 1;
    attribute mti_svvh_generic_type of fpll_cas_out_enable : constant is 1;
    attribute mti_svvh_generic_type of fpll_hclk_out_enable : constant is 1;
    attribute mti_svvh_generic_type of fpll_iqtxrxclk_out_enable : constant is 1;
    attribute mti_svvh_generic_type of hssi_output_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of input_tolerance : constant is 1;
    attribute mti_svvh_generic_type of is_cascaded_pll : constant is 1;
    attribute mti_svvh_generic_type of is_otn : constant is 1;
    attribute mti_svvh_generic_type of is_pa_core : constant is 1;
    attribute mti_svvh_generic_type of is_sdi : constant is 1;
    attribute mti_svvh_generic_type of l_counter : constant is 1;
    attribute mti_svvh_generic_type of m_counter : constant is 1;
    attribute mti_svvh_generic_type of m_counter_c0 : constant is 1;
    attribute mti_svvh_generic_type of m_counter_c1 : constant is 1;
    attribute mti_svvh_generic_type of m_counter_c2 : constant is 1;
    attribute mti_svvh_generic_type of m_counter_c3 : constant is 1;
    attribute mti_svvh_generic_type of max_fractional_percentage : constant is 1;
    attribute mti_svvh_generic_type of min_fractional_percentage : constant is 1;
    attribute mti_svvh_generic_type of n_counter : constant is 1;
    attribute mti_svvh_generic_type of out_freq : constant is 1;
    attribute mti_svvh_generic_type of out_freq_hz : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_0 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_1 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_2 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_3 : constant is 1;
    attribute mti_svvh_generic_type of output_tolerance : constant is 1;
    attribute mti_svvh_generic_type of pfd_freq : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_0 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_1 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_2 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_3 : constant is 1;
    attribute mti_svvh_generic_type of pll_atb : constant is 1;
    attribute mti_svvh_generic_type of pll_bw_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_c0_pllcout_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c1_pllcout_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c2_pllcout_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c3_pllcout_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0 : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_min_tco_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_min_tco_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2 : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_min_tco_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3 : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_min_tco_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_cal_status : constant is 1;
    attribute mti_svvh_generic_type of pll_calibration : constant is 1;
    attribute mti_svvh_generic_type of pll_cmp_buf_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_cmu_rstn_value : constant is 1;
    attribute mti_svvh_generic_type of pll_core_cali_ref_off : constant is 1;
    attribute mti_svvh_generic_type of pll_core_cali_vco_off : constant is 1;
    attribute mti_svvh_generic_type of pll_core_vccdreg_fb : constant is 1;
    attribute mti_svvh_generic_type of pll_core_vccdreg_fw : constant is 1;
    attribute mti_svvh_generic_type of pll_core_vreg0_atbsel : constant is 1;
    attribute mti_svvh_generic_type of pll_core_vreg1_atbsel : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_compensation : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_current_setting : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_lf_3rd_pole_freq : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_lf_order : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_testmode : constant is 1;
    attribute mti_svvh_generic_type of pll_ctrl_override_setting : constant is 1;
    attribute mti_svvh_generic_type of pll_ctrl_plniotri_override : constant is 1;
    attribute mti_svvh_generic_type of pll_device_variant : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_base_addr : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_broadcast_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_clk_vreg_boost : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_cvp_inter_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_force_inter_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_fpll_vreg1_boost : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_fpll_vreg_boost : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_power_iso_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_status_select : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_ecn_bypass : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_ecn_test_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_fractional_division : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_fractional_value_ready : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_out_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_extra_csr : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_2 : constant is 1;
    attribute mti_svvh_generic_type of pll_iqclk_mux_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_l_counter : constant is 1;
    attribute mti_svvh_generic_type of pll_l_counter_bypass : constant is 1;
    attribute mti_svvh_generic_type of pll_l_counter_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_lf_cbig : constant is 1;
    attribute mti_svvh_generic_type of pll_lf_resistance : constant is 1;
    attribute mti_svvh_generic_type of pll_lf_ripplecap : constant is 1;
    attribute mti_svvh_generic_type of pll_lock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of pll_lock_fltr_test : constant is 1;
    attribute mti_svvh_generic_type of pll_lpf_rstn_value : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_min_tco_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_nreset_invert : constant is 1;
    attribute mti_svvh_generic_type of pll_op_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_optimal : constant is 1;
    attribute mti_svvh_generic_type of pll_powerdown_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_ppm_clk0_src : constant is 1;
    attribute mti_svvh_generic_type of pll_ppm_clk1_src : constant is 1;
    attribute mti_svvh_generic_type of pll_ref_buf_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_rstn_override : constant is 1;
    attribute mti_svvh_generic_type of pll_self_reset : constant is 1;
    attribute mti_svvh_generic_type of pll_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_tclk_mux_en : constant is 1;
    attribute mti_svvh_generic_type of pll_tclk_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_test_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_unlock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of pll_vccr_pd_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_0 : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_0_dyn_high_bits : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_0_dyn_low_bits : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_0_fix : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_0_fix_high : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_1_dyn_high_bits : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_1_dyn_low_bits : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_1_fix : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_freq_band_1_fix_high : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph0_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph0_value : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph1_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph1_value : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph2_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph2_value : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph3_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph3_value : constant is 1;
    attribute mti_svvh_generic_type of pm_speed_grade : constant is 1;
    attribute mti_svvh_generic_type of pma_width : constant is 1;
    attribute mti_svvh_generic_type of power_mode : constant is 1;
    attribute mti_svvh_generic_type of power_rail_et : constant is 1;
    attribute mti_svvh_generic_type of primary_use : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of reference_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of reference_clock_frequency_scratch : constant is 1;
    attribute mti_svvh_generic_type of set_fpll_input_freq_range : constant is 1;
    attribute mti_svvh_generic_type of side : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of top_or_bottom : constant is 1;
    attribute mti_svvh_generic_type of vco_freq : constant is 1;
    attribute mti_svvh_generic_type of vco_freq_hz : constant is 1;
    attribute mti_svvh_generic_type of vco_frequency : constant is 1;
    attribute mti_svvh_generic_type of xpm_cmu_fpll_core_cal_vco_count_length : constant is 1;
    attribute mti_svvh_generic_type of xpm_cmu_fpll_core_fpll_refclk_source : constant is 1;
    attribute mti_svvh_generic_type of xpm_cmu_fpll_core_fpll_vco_div_by_2_sel : constant is 1;
    attribute mti_svvh_generic_type of xpm_cmu_fpll_core_pfd_delay_compensation : constant is 1;
    attribute mti_svvh_generic_type of xpm_cmu_fpll_core_pfd_pulse_width : constant is 1;
    attribute mti_svvh_generic_type of xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost : constant is 1;
end twentynm_cmu_fpll;
