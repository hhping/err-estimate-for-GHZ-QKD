`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIBss5q9EoZVCVackYpRsGka7OfE8eG+ycQRSQWo27AYp9UTQ1LLrHMcQR3CQfp4
uu9zsVGtu+ZoRFr8YGN/5NQK6ll3Q597Qe0c+iAI4JG2oQFPQpzX4dHYlEtwHR1G
4U1ONznqzenDaUjBm9ouZqUQYL7/es1Tr2Q+gfXwMhSrwweDI0SYsKEC7d6HjqgG
Dl/I9nQbyS7ujWP9BN8XZro81eJxutmQ7EL9gQwy3Sxj6x2a6R0v/2id9GJSf97l
z31aLMeL3ui9W5C8wbQjm6aMTvKo6XMwcPqQUPLJm79P9HbC6ik2k4oQJ1CN2RRe
p43OxWsmLX0R+VOPjPiQrXaBNWb92d3Wqlx4EkTeEsXI8BtO7FPNaIHgIBIQKGge
irmwbKOpUCFMepnlbPK4teDQ83L8XSNkWmJ+6C90IsgvqYnlwMT3J2MztYAoprOB
OZIjgaPQjItKyMVjlATqMMQqG3Ch+qtucwRFnpgknxCENWkx7xgotgLK5JkOD/0I
`protect END_PROTECTED
