`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hQrRUXd6bp2ltfwZ09jl3RE5pu8r7rhoJiWa2l9qI4B4YZg5wZWCexsKJPgyEzk
xdF6nzFph7dO0D8b9LDnGXLtK94oPNYpXog+VnpCptND9+FtEfaKNhAh9bIKZGmX
HtncV7A57uN1XykiuojgOXId/b4S/3p05gEqRt1wZh7+rXsGXgEXc6cIWPVNq3ta
ErBJlUg3CNV1nqBJDTMnFhGSTu7MJxLloCdkBNY2monh9VeFxppmutxhtg/k3tdj
jyGRFNfOfvUxiCVAz1bzyAToe/5ZDhtU1HdUf7xuiFvG6Niq/FscFLAZ7FCYasC/
K+B6K7r0gYyyj1FyyLhQzcE9IsJ8fzkFHdFw+P2Fsom1ZAiZqlop/Fvg6WSOWOCa
yCSZyM4ANYvWitINFmqzrB4pHLodWuFPJhQm1qsJA4g=
`protect END_PROTECTED
