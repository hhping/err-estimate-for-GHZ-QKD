`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q0AMA7nTDOBk6+oop6e1Cv8EDk27Hq1uIxrdwNUJ0treCCmaw7eUNH8RmmJPuIDd
17XYvKz1+YrqARD2cJ2T+B4/knX4xo9PfWbSmsiRTV8DQGXoqA/qSlGpNYu61CSZ
cjvQT2pVb6E4HDOUaIaLUXnrQCORvE8CdybqIQFYd+r2DziS4J8T1oSGV4kJsKnw
eQznKCwBkRuctkZkdShqHDhIVY16EstSkX9Iq2h8Uj8pCqhZ5jjKeYGEL2gsUZ/Q
2/5UoDE4i0WlG+6Q05bJpKTHOHHpDHbFqUiSs9T3OVbZwR2FSfrKnsbqHUbBSM+u
s/gc+JQBu9H09B226mr48oVKQgABchwaHAmKirOTSGavNXSi3ZohV5qBhmbX5hn2
R+PWFDBX0LhmMziDu3C/Zm7g1uFtUyy6OamsBABB/LLD6lYhNYF1rJtbXY8M1xDb
b/6b/trH2JXcMvOgPv+JeYgXnR7W/AkHLgJeYox8ZcW1sHhQpFFuBAG3vy3v3JtI
haqLHN4BnNcwZEe7eOcaRc5QI9ghtoOqtaHFjVT7Wv1/7ZbP9jAGXQ5cUB2ApYFi
TS79xuqNslJdMhDAgbj6nornLkswDV5fXpFU3j2vVuuUBcYIcCe0RZEuVtXDReON
b/Gb+lGqvWWcLb+cZ96xoc0W9VXRDkoNYw2W8aP79S9sjhxGBl+QqBYOswkI57bw
ZXwBKOLLmh8qBgfekVLQsgUCRGB8eAvcQrQuAWbAAmYIspXpsuzP5BuoPT3VFb+P
h7CyVdxHztYjo4JHAhdnQ9JQizuK/DnPhY2dN56AxBmwlYIOYqpoFTb5xx/GHA//
JUWafEi9X25ZmbfuFhvNUffByMQnvlBMVb5e17UtWUPD7dUrzUCm4aoaNNbzQp00
LB1yzPZasJyTQgL/JZ8yMxponF6yIkIsvbD+jw6LN+QEn8LyI+lJSO6OjsclQd6h
0hHLix8uAWBUQTaJF47BUiE1lLJnqzO9mN1rgDqSpPmMiohZrrHg6ZP8xTXQR40v
UB+2rwxQAo4DOZ2yfgdoKZ+jZ8DFhUizN/atBlQb4F8dCj00PchUUObZbN2f7QbD
Rjp4Q7aA/TW54Fl3Q4za6WMh7o2lDRHp3DQs0WtIKUTEB/gW7z8L0s557rOdfZ68
teY3ZCqRIJ5m1eNe1ReCo2QMH679DKYLIdl8sBXx2VDjx11w+YRjsVK1MyAVh6BT
n/6AE8YUr1ptqbTGf3hcdPQfmW1MiaMelmnUFigVdi0185sMAl7XleQT9ysHDqyA
R/gZv5R3D29JoJ99w+m/vyp8Ubs/uR5sOM6vpLElEUr7U92UcDuHfIicHiOSGEQH
b6+3V8KHo1PG9wXRytjvq+jyt9gifanN66AZuMmQonHlgn/Aw7ldutnRJHrAIlml
e0w5xwmc2UG2Lqn2go9wb/o3IXFzjC6W3Z8VnATPZnw=
`protect END_PROTECTED
