`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hSfbIO8ukFO74R+xwxWIDzJN1yEzed87pPea0b3A3CYr8JCYGO8DR//eBJT+gahi
p//8LPRGAWrzWtWBnLsLDPvlFoAu82/65zHm3g51uldU+NOK1b9HX0Y7/5YVBpA4
GhSA13VXFzSIcu/Na4HyZbBAQFz4rp/s/wveOqf0fbhz6SeW87dx0u+IjCS1UhRK
trFqxQE3E7pedf35oFDnDx+XH61t2quGMTzmT/Dgzf3WxFhigtpdh5Ib3vOos3Sa
2g3mWhOJnOU2nCeObLVJjreTqLrnw1AgPxAc2s/5V4u/fFyUAGTUnY8xbEfGTYcW
RY2WxxWn++8PKD/4Uc0ZYExhJjAy39QK8qSgzb5oNNzKwNKzRYACPu9+JaEN2hOb
784ubh6z20UZaaXpT87Y5233Vl3E/H3SfKo6MBk1peu/K8TZ32duWfFgWg6L0zW9
vMYqutLsWWP2UH/kFa4VzQ==
`protect END_PROTECTED
