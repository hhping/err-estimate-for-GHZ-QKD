`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQfR9ahKcrelPB6pCOuP2wyYhnP08MFulxPxWm/0WiW6c209V/0UIfUUlsOGe/fB
33egp1UjYpXBofpLzD9xQnJDGI6UihllA+u4qEQDKkzFCGwlU1uE6ZsSlY69B0EG
DPPJKQYzx26fYtNIs2xHjj8tOCOR2DtAkyWMYckuuP4MLsxsYvIMkvfbg66zScu0
LWwQNaN9NAMiLO7B86eM4tg/bcqKtBN41LTwuNH+X+sClsWimb1dsYqlbH9JlY0x
XGHbWp1B5/zvBvyuQR1bCpKyxupq1t/Uhvmkkcn/RIBBE/T2z5UOF98I8yuuybcz
w9KqJ3Cxz/3TofCDXTWZKgq5dSq3tQllly79OtbAdQMzvqFF0bzHhAepK1bo3Lu9
syN+5ef7JuIPJYBD2ZGW0s6ZcqKzxlnd+bfvSjU8isk1IrCGOpqUhV+2umORAknB
59bqFkbhsDxCS6dDGcHO3BqocbVO61iMHyOPF2ephYsXL5/7n0gudKR93cviiDmC
fyv6Es6bgwgYVosE2BDX0EGO34JHB4TAKlmrNQ26jPyMd6FBha9F8SgQDa6GsXf+
yZKXVsygOVOv9+4RlQD9eOS5XmpA3l8fZTOBDPMUI6NNkaNBRIpCusfEWPa3oapu
J3A9Fx17OhLnHM5+INXAGU9uF1+StumJYRgYhzMf4YsZOOLhBtFpfIgIhwjJuQnv
Ymne50cHxdPU+1fAP2og2eWLUZ/W4wRxTc1ycl+9p8VqRHMhu/z78gZiB+F//luE
58juafViN/0Xj4V4eiYB4wcC74C/TquBthgXq0ZAI2IJYZuFrxK1uE7B1sNlCOjC
zEDONyr96ofsllkV/ZH97VpEEWGLEdcfe5OWO+fESsnXaURGQVus/zRpfweqqQNY
uzS/ACTS0RoMb4ijMNZf3pZ9dLsrfn2r77W62JxZVdpTqCicZ2AgrdVxT61zF3O3
zg1m67mgRgAF5Npth9iCk9fx3ujj+KV62XTHB2MPfrasChSTHkT+ys/Xr0NXwmhC
YJTgc1eHBUk6g+l0LB1zZIJ/Thjr+GrypNw+WnCRtZ7yb37Yi5kk808ibzlBSL4v
dlh/Whj5WCoc89YfFukJQUJU5NLjPo2E0Ee6fPSXd4uKYr1rIzAJrK9MYRKY5vT5
UJqNRHmzYC78RXcJuL1QOGEz/mId543pQUa2o80O6+AbHVSRrhkRytcG8KoZWicP
5z+YmcD9Xb/YbIXr0KTgTCw256kvOyNM4rId4p9ynIF4PNqJ2NMu5mOQ+9utsIg0
7Ven+ExpOAxb+eEeSWKsgpYmaLPFvAbTr1nTHjF0+cdqh6au3ItTaiEtlnfxna8Y
PWWmOqkdgWDxeQr6+Lria+V0+sJijhP6sTTL6d/ZSHLBll/B3/V2nNe9CGOWhLKR
zR2P0Q8YpwKX/l5b4zZ2uDm66r4cOKEmIV3bWPV0m0Xjp2uVDieL4KHu4xoAwgHm
vzqhxzFy3KLILpwEtAR62VxKkv9PcaBJfRuBxIt3ho66cW/4qEVkFlMNKR+Hg14f
ZnMHXiG17AIDabJBlqpX+AkQs+VoL6TzuhmEaRhZCZP09IhHFxYCvCPixzHzZs0E
usU9gO0HhY4bII6BrgA+bvF2Ojd4xEKsK8X0XZjZ/CZXB4RCApWJ89Dhl49MwVop
V1tH6hvsnDN5G+LLhg03qdGAXKkIzaaWYULSL9/N12o=
`protect END_PROTECTED
