`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NAsa2ixF/IKXOipcbpAoiDWqL3nGFY0i1v7c7IQaaQKjzTuFnv/0wdwCfqM+1e3
feKMzbG2GrrYUTGrXzi1AEjArzaQ7LyEbO6WqT7dGmXkiF/KaKxCB/esY3g/Qjjk
M56HO+ZWpGI0pIs+w5cVVX9zmjNRKvD7Yy87S0CNOua2T1ymed8oKcG0SWOseNh7
dXDkLmhi7FPQWYiNARxSPfFO6roXHHyr/X6iZYC7NbISlzQ+YEAvB6JJVmBJbEy3
CpZKqaLlcSAaSFNzB7jgkjVPcG4eCVbjscF3P/H9RzGrM/vCaKCaIeomr4TZENN3
2N9Y7KUs/JNTAHf3bvAc3oRGfDT4al2DxU/9l4BZI5Gadf39xbxpLPQLM6ed2X7t
lZXIwT/rX9OUlSTi7h9K+0onaB5u71vZ7BLNwF1KHD48fyslxoWMLipCwMOAUnS6
kFHsh6qzA/fpIXofWm/mOpTQfEgBA3V/uBbXPVfJz2YUE1lIpIyT3cuLDGyq2NtP
cNNo3HMDLWVEs3UrJDad+KWt99Q5wgZh43ZxZl1QDYeuTS3LS4iFbvcJ2xZaxpi8
/svg3MYj3XhOPmSmW/0wUMkjcMMEF95SLMmWbwaOesW4oC6t7U3KshcJr6acW6vV
PNYV42QXaGR/2ctNqh2OUQGs4eE4rLlJqdUAawGIuzoNC46imFvDJkYfokGxV5Z/
eRC1Qf+wTFdr0fH2BVUwCNjAxohxZizfkdN4WjFRKAO8S8fdgTQmvFFXN+yFZDhH
jvwCU3d8cLL5umfSGpA3WIHlB8J+51RKmKZWWapi0TQ2uUIkDoI7ohAvF/CXKAFg
nboLU55trx0wRlofK33hvG2/DGjihZnzaEZ/1Zqv3HMRHKBv3LCmQKBepYpCv5/j
236l2UXUtMJLIfEH2sv1nC+HukGvYG9J4ex81jEEh4CWFZLjX43FV35xnbME1UyQ
79So7XwToiF18SDjxc+QvYbBYQW+NyKBA+T2PENTaJxSTIvBX9fZg4+eYeGxuWdq
gY0kE106fX4PqKge95TtAzeZvXsP6lByh1Nd5bKW8U2tX2hkjMQBYoSBpCoggV3O
aJOUwZ3CkwuT2wjueRS+4nMPc49qUd8OCzQUhYfviJzbe7sjnzRr15OJPDHjNRcg
EgjgqaElsz0FZf064DKRckSWYSxoQmkD/pEJgHlnz8wcD/TsDd7j0S3iXxdjx/t1
htBptB7PZJISZptdrsRzaSe5Eq1OCfL1LMw1fEZHUkSg3Jd7UxzpFUVbkXJKzvbr
16C8pBI+oCY36Fsxq4MLud1kRprmZ97HwGeR3+3+NbAN0WrRNoh3DS2Vbp3kBnKa
oe7QQLqCl/zmQuAg2J7rEWRsnkzEgGVS4nSVP69yPegDZyViCqxd5hA4kvV/6SyM
HiCSEWnUp32OXi68dh1Jgn5WlMi0BxeXH/gLXLpBy+CTJnHgRogGxzVdOYNnBK81
yu5J3RYiKiDGCan5DjrTo8bs233O0JWnp5mMf9ELrK0XEjBfX4b2fkN345FWEVs1
`protect END_PROTECTED
