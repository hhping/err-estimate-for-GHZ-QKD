`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e8K5BNe1s+V2KNV+6JRbYoxavo5moSiab8DyG4b9bkY1jD5g7OQXOF91EDlrY7S2
8zzLQDGNjHZc6USbcr8IsZ4APzUBWcqSWdecRrbgyUrdWde2hx5k+pvN137Kn6I4
DuMf+E4mM/nir0XPlTIaPUJ/5oNfbtCdtXHjCPrOhPICh2nDu3k9FWYRs64z+78r
grQ56CarvYr8lDTKheW+NHjdO/doZinFGCLftmRXs027NYYXF0NpqZLoH1iKbRLP
fFcFsqBiKe7OMNNk2FzOG0cy6TUgJCGuw/e2NomVPpwXXp00FLF7l0XqjQ+G4mDV
PEWMRk1/fIXINc4EvTFTR7/Y6M7EmCGvjzqx3qM4cKiYvRGsYsa1R+NSIlQOBrcF
ZbthRQSXi2ypTqzAMglW1o/mGRL+6geVcx4/cTLGM8CcfoveOwhMLPGTu+Y9B+wP
rvNE7VOmFN/CSqChXr5H7yAYxf1hIX9Iqcs3tsGMTMls8MaHWLj6ZGfYcgmTAUHA
BSgwJTls8+MIxt98GvQm/3qmoa2sbFkt4SSs9Ukj8Ftg6dBSoKjvTe7+lbQvVa8n
f+mj82GxwryiQFiwq/YHbrmTtAsA/eYd4oAtlbSIaZ8oHIkB3bmHBqy95KVsnHRM
tE2F+FEtGFDGkbkGFQjsFAxL9qECWzCPepLGwtfI5fjQ5SxIqBJsFgKEJbObJi3T
f3YJbbggbTzNapL548UhDnLtBnOoerH9fU6KfRlRi9+S2rZVoZzgqNqIlPkWlN1w
2Bh8MmWnbW1BEOQJeihkGuROumvXvhPNvetYsFXYE2f8Jq3By3DbSC4nkOvnVhDQ
Kzq9ptNzdqpjdAvMy2Eq96k9tdhuayYV1Ka2PU55h+UFxsKxafiDUkZeSYe8xtoq
HcEnE4ukkCXv9uApX4n3/2DtC7kFCUTNHlxlLh5IZQOJONpliE4fpsG/G8Shxl2K
Fx4LjVfe/yyXUjCi7+2P/v6KseXU6lqt075WjOTadzG+NiMq5WmP7AGaqvjGPjpi
NZJZSnn6Wj7X03cQL8JTDbXixrHxjaWpZQ3uXejJkQRuaeyacl6eeC9JhpSqRdpe
HJ+VS9WEKAIuYVGQu6dq63POomTtWy8E3itJ1IqlVbOWeFdYnmz7+i+FJjLIKDT2
vgBD5IlDSTJXNydoKq5j3KVoiLrRD5JH5Ogd1w3jUAEwEpr+zAm0cgCt07apJN9b
+1kroBIQwLXcMqNqUrZxHZQYF6scub7kjtEdUEOYx9r6UrpVM846rExeqhcmstlu
axxhQ5OL89Lhez6X01/MRQ==
`protect END_PROTECTED
