`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1TadNoQVuQvV6JD9Gl1SLUs5rsvhEdLl5E9KUs9EKT8fKZxe4oqVVsWcebNI9BvU
drcN1JryIAmOu7R215W2A5fjxyfSg6hNE60E0npNWrKenKtxB7TLmbz4GblUbdvw
8T1PM+Asyvx/yD2BW+2fv85WBpJcO7MOUo0DyRUkP86AC2AbUpo6wMv2vtzJiSak
OvTYNgd4sNffDVsc3inKNi8F62uRSaCtMhfLLgb/F0Lxq9cIoojhKjCkAc9OGgV3
W694CSbQ41iRBW5BRK9c3BvhYToj8y7YE4zbyKtVJx7CRnr/Vbb07Sy9zlC2ruAL
isWZ+XU/pWyMuCii3tPNZ51MfC5U17kYLa44484W/LGGxsLQPtdxo2XqG2GnD5wB
0Yy4pOUCCLx0jDNJX2I98AfSxdtrI7Ra29N3hXaWWicysis/QJV0F8MTujkKFbSy
XBKsnZlz8SPo3YBlrCu2S+7O0k6hXsvfhbYlHw1SCEZfbbyMMttlBFqQbiQ9/gTM
m6P6dMOVBgu4H3Tvmt9yzhx4epIDcfs/Wt89Skae/Rlt+3NButmgg0lmgBkDZMeD
Ri42vO6xXVoRshzW51gEkRPF8PX7tep/bAVQ3tsZV3O4GnWrV/CX+l5QwdiLlK6I
Nz4lnMRBU+19t/UqisesOAmXG87WlkARdtKDHKZ/y+rJtAAyaJ7vexaM+xGEsNoc
SvKHgUzyZfzml3g+Wn9cPXxSYJJci8O1ySIEt3JdpVtu5kMQCfPSFPZS1i0ZUsch
2P8yygE4dopHXycJYtPPOPqR4HyiCvhvNTltj4ntI78hXjhDsxPRyxPkxq6Cm10/
`protect END_PROTECTED
