`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mL5BUOc9vNOAiLcJyKP0wr/5+N1wkKi7o5pqjJ2gAU0r+TCC8UiEVg3amUKBIp+0
Hsuo8+sZqKDlwv1WHwP0maAbmIDHHdxv3uxhCkuSohcq9Abs4TheOLKjpHP3XDgG
mzcBrY9BqdLqlFxvvdiuai3l3W8qPEzN3SC+TvcOskpysJ7NKSLBj50RirIVwwNe
EtoGbZPt/0FMMZOUg75vD3Mf1uiyJxgp6sF6XyUOcv94dpn1Rsymc3W00OeT7X08
bPkbsQrrWis1LulxQgh6Q4wUtubpDiOjaT2JapOf/wugiqrSH6yInDl22c03HACH
N8hlRwXwfRamsJFwDPCLP8Sj4IiS6mRnA+aeOB8geX0irLtWLC0WfSD2LJcuQLnR
h3Sb5ShBLIvVTRt8/JY7DhX88FACEf3YCI3lXGiMBOc/H//wbx/vkg0Og9yo9Oht
PBLcrCAJDttq+B1zRhI51LEI5pCbFQQ7BRGZzAvrVW0dvNXxj2KX9BT6+jSL0kA7
Rw9Z6m6ixQJlpzHhi07OHz/KPIneeOMZ5GbDmP0zuchPzUG2efij0U0IPBUot8fR
YWHW8oRzOhtsfqKgzRGIGx6I3hA+U7myCNliMoJTl7iWHSOGeLCyrUOvNwWcH5y/
5E6040uc2nL7Ga/bsOyZdDw0RJoTI/alZaaJ57mnN7iKsNzpWAC1VXMPnQUnSIMo
Nd/25jB6/bHvfCMChM/dXgQglc2yhaL+1ZJ2U3zsaAxW9dhmM3SHN9y8GMHlf1qv
nvu7d63qw9JPwRlgXwilt6tnX61al2s8QZhckf7mjgwzLS3OIbYzxCyyWe8ornfi
ehdWq1T1exG4a/ryIKgE9K5EdJJ0U7uvvx0mUat8b8lQJPX5R+Q7/6eiYSLZq5+s
2Q0ccK82rk51S/LpEgZa7HAyYTa5J8/uUFbZ06+54YcMF6cuiaXxDL7xaqR/jARh
xjM/iE+0t8L2a8Nc1/eD8KgmeRvJt8FwqiHWHQILnEpeJbJTZ7dnLVtYfxlRarsz
GikenZNyNgA/7Js1afR9PwKhm9GcAM0vvAfZJbp6IqerG4z2psQcSpfPp2GSap8+
DKpv1QhGqCuxF9Bb2SfMAQkSKX40t3r0Av+1cO7kJCH/mywHl7XD4XqGoBBo0X34
v8BrO8FvkCCxIaSLnB31LqCk37BMoKz3HMaAsNMcknPkRuK/HC7ZXpH5b8taTBKA
d0bS+q7wqsf1ie1TvgxXZ1O4hP0hgdtRa1dcEAPouEF/Wf3oN6so0ZWQi6EvKb7H
VwTNVTUieFG4WJpjHCdwGrndgAxNHzE4rWSMetwAGC/LWDvxcXdli3RFd02GHekF
P6N2Cm3zu215555wHctz+ersLZ1dvK7gxj+NgoOtSROwpLb3Ayl4SkmoD4RgWzxR
a37wU89OrRhfUAT/77C9qtjyZzyNZvTt0Jd3W1s73UPaRIAZ7NNdGY5DyrypkW26
HfL9Dwr2Sb9Dvuyu1k9w4d0IIBoYgv8JevoZb2EFSPKqEDT+98K4WZTAqRVjETC8
qkZ6M92Sgl1QBdw/2r8XaRDEf6OYaW6erbTaqnyUmcmoSKL6Q46k2M0DVn5YfYfX
3OePHb0gu0BdwLITubqHR4CzJwKNRheIO1aZy7bXy2aF/9HcIuFzBdsmzzwwupiV
iQu+yMM4tKEBZOuOkw5fTfq0pF3r1iJmBw/zqcodLWKriTt1lW4idKuYCQOP9gn7
hYEIWAljHhOGBf19/K9SfFmV8DGFg4Uo9ViI9nMIHtXYBrEADK9sF97YFqOC0NVJ
EfgbzCgtWiAeK66GMRrDvZXXJtJZWo0xIoTaYRqgR0fr88wcUQRjY1cS0Dg/es18
3xRucgSeoQLKHIK0XwoicpRZTEqWerErLLGQPg3mRZYwG1QKRTvMH4Jy3WMQ0rRm
3qHsHyLOTdbjdVMdZQ1jxZUrRlxPfRtpm/ANC7gnBlo4cGMyMcGV73bkaDlOHOVZ
FfTVyGTL6rExczgm8OjgE/I+d4+L2oMoWH6uMTv6VO3LBUfgeT3Sr89uwwgAwesg
1s+8mbjhchkC1o+KlC2XOx4tBdoltNlzSRMe4cunSYM1gSxf8koB0etiapSd1vZO
gEVsyrBJCCa2qhH0B+yqTH3xFagK6hI/Lzw5keQ8Q5NwYMwsnzI1NM4+Y1Mw8+EY
YwRm0pKz6GVvBwmxh0RF9y5hSwX6576vWIxZ3xvT7sNRvixxqf2jtM7jyQnHkinQ
K2ZU3aKC4mZxBPSXQy72NT+QMEdRnssQySBmnEj83Qy8G9bECrmwv0l2pZ9Vavg5
3HF0s30G6jI9cme4yqn8cEf/AEUV4pEPBnp55tpyfrqzi1UDL3mrmLJU3I9Pi4Gy
CYIfBQDBlVy1ztFWJB5ZU9cO4YB1KBOaxhJiZ1RE7HqrD93ZVpahIDbdWLljxWoq
7qjQi2DSkQ4cKUMy/UYn5zOrqYKcwoxJ+mOtIa2MtngDd3nqfkLafA2mCqRwX9oU
iuzaqYkR7L65RtMQFIFOWdtSI7oo28vFBhj2zBVIO0bUJ3dL5taon9rnJjmwd1OR
+cwudYSJTRdfZ1u0DtlKcFzLHi0lv5OggTHZEmDbquMzvgHgKK8dQfr3rI/jkc+O
Rq1rMlRQrG/ZwY6ppNBRTB7l2kefBpwLcmY1ouOUDziJkM9D+wIxsJ9y8H0iNrms
`protect END_PROTECTED
