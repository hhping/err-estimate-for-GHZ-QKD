`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VyjsTzzxPMFEZSJbcY8hRX8+ItHfh4cXCs/aAV4ut70eidfr+V389DGMVLg27zvw
gnmyectWRVI2xEyedt1krF5G3qKNj3wkyYajQ11roZ5shm3oan+h6ndhbXsOVTB/
0prITPxkhYY8H0nFSryTH48e9//FyFoVcmrtOBHwf+8+XfMUj5B6G3NaT+Y0Z39I
HYrerrvESPaqknnKXeKxdWhsCb/C7CSv9prCxYCkHTZEGW0CcaJXKdJ06tBK85Iy
66dySm1aYud1yyhxxw2djZM3Pturz0wwG8+OOPvNSgUVIDqfwbEQnc1Wf20KvCnF
sXoRhvveXhLN5zsWWeRnhItFzp2cc4B/zgVhZgGSnXQqYPWCMFw1cTRwh0IKk0vw
36VyIzo9KAXWgfswjBOJOasCxWvIuQ44DmKe/SVTHOhSmdLkewBuTEPPqPwT6IP+
N0vhjlWrfContp//uLZtg0oWHZbegGPHaru6WqjLgf3Cp59z9zrML9pfzOOCht3o
HSNWGfSs248GyKAEgu+m+HSbowhtYrm0mRMVTR/1bGv8FJ6bHjZ6HHqjJkrg4Gnz
kM1rgCcgA/kdjIx1KStXhqvB4cd+LQt7R4Z4Hd/rYf1gsux1VAPkJ+G0o3btuI5F
cs7dKbFpIOk9L1Hsw4LPLi3BxXXLNsT8TmMbBO95xO7szt4yHe1llvVkEAYEVy74
M8QAZRmPGSi7jVkJvtDhdqeptwID1Zs1XZoujy1seb67hO8u+dcZObOI8tRfuGi9
GspKff6ydhslSVfPGrHDkYPx/R28Ix0qZHXzfsRpZ5azQZdWnH0E8YmMaMADCbuc
3FKrMqJXE41yaU0qJ5Lbq3TJzhe/mEIdCOiXdcgi97FzSn014jEoUdgeSHRL3iHW
5rJfhW1F/EJs5+x5ePtCN4KVcpmtJHD0dmHssVAZYMoOjiBaK4SWjVWcsIrS8C3d
ocaXqYm8QWRlqAsNTEGDleUHA0R4nut8ctoKDcl72PaKJGv/6aCCf6P0XoA9X/JR
E/vle1fQ9JiJaGHFC5sKBUAkRmX0lgmPQfF37o92oEjmh5x1u/JxPAE1ChbWUbFT
FDw2gUk5GQLuyTJAuldtRZhWi8USrmaA4mmMM8HKQXVWBIhcMVDJodZO8wfOF98T
t7/4LFDxV0jz/SfMDMSO6WYPQQlKzihAj0GOjS+p3PRXOxe77C/tlVta3qXOZM0x
XBAgqNaTcaz8l3GiUJnMxNb88aImOpFUe0ZOAgQ4LR7JoIbk00Izn2Zvhx7VUAFA
doPftU3d0vcORJL3o+vJJCaF567M2H0OqylXRLwBTzFjHaciXcSal/YDbe9S5tpr
wauGsN/e5rXRtxBRNxJA/d1mbMulRGy5iY2mn6iXsn0JpCU4CjX45Q1gbXr88VV1
MnQiszrDEvccF2UFEhOrhp2eUOG1wb2JTNuQVoujYe9KYYCQaE4QSgDKPqaoaEtz
mtsJmoutVU1wuYSLii1GlEBI7l4ZcfhL0IQ22Hhiolm1jie/q7fHatfIzR3Gf+6R
`protect END_PROTECTED
