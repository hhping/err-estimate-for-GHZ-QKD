`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vNTZViQ4dVocg+O7FedPpKCLZphwB1c22oM+R+OGPfNlLIh2Qd69LQepb5TUu9D
UXt3pAv/PqYNb9+VJwc2qDyMks8kxPxx9751lumQFtTRBdDEAfsa1igq0usLZm3f
//aXPeq/Wdeijq+Xhg3NlH2oniL4lD0flDmaFyUn4A3YphYkeMfGnBgJ4aStrE3s
1PQkJPHXSQqYfnJhgbQZZ4ryVLHC/pozfeGf9ATCDhYUYRsJVlQ5ye7o6EcO+BOj
885R47xxS1973QwrCyEvNoYUJyxGjNr9AOtuvH5m7krkm0eFNcIx7VYgL3U/7f3n
ypGmVGJzJwkUMkG9/oZuiyHMYXKNkk05fN/BlxPcvb+bLAJ2hwPvnXFdLcCa3WIM
YfCNjg7Ou4zRPbimCC8cOWIc8eJdq8BYGu9D6WuxOCHKcbT6KJKWtKB6ARwPwPNf
Ai5qvdtVRM/iQr6u79XagMeHC9BHL1h7CzsYwosh4zlAO/W7722Jdh3OVzBj0pcm
hl+yAIag0a0cz7sYALjTDNIokU0izaoYEC1uL3NOPFCevI95quXpHg6ygcigjnnp
6Bnaf1uLmgxs+xtH/noczFecAvugRIz4iBAjBVUemZ13PQHYrL5wUIp/2+VFL+Ol
5QJVURymEIpaDwnzl606QqoS3ZloIS5U5D7BLc8NcJwPpHNckQQCXs8NxdHRPhmI
fMIyyh6uyVv05soKs8q09miNbLE9h6aHOYKgL1l75ULylliM2CzGEooOecmMhCNI
lZeaz+JU7bwxM3R36i7qyvyyS5bZIeKO039dOFl1XnT33Xgkk9I4n/CnPEQ/BpvF
FsfciX8OJslRAWH3fTDsLJxZuReiUFr0faR6fB2iDFzCbw8pMERi89NL2em1vDDw
wLxE4FHPlO8Ht6Og9emkvWpwlkXKfbEvRkD2wZHx14iIItEek0J5IMf3axBhm5Kf
PJviEUSVDoQ3KIo2m0+UZIyIrfKG6jWg1zZdIRhuryE/CATqxq1xG+zrdiVr9aur
5D6t7HCZeME2Y9cHN6Rav5lI72RjpunFURDMN9bIhXApNXyqN7WFO/Mzj/FhSE/Y
eT2KsMKajS3IAriplREScdaCoquddGQWUgHnkfj+xqXGaSoVgCTF6/ct0uCa4YeP
`protect END_PROTECTED
