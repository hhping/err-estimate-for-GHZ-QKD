`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNK2dPOnJYc+du5BBhjlxPyFF0boe/K91uaaGfCY5LTT+cmHDFdSoQD5lJGqPE+E
IRSFfJhOWHcRce8Rm03UtCpi5Y18B8Fv0IE4KAfxSQ2+50VwuGUvMaBinM387wL5
yLZRni4htIm41ljt12OALKn0czEFadW2LSiGgIVhrhWxX6tXdeJcldV0+MrH4H9f
sqXF8bf96DmM5PRHd2Pw76CRkWu2DrC0dgXRPCMY9I0mRbRvXYpHe0VZOxeB5Wcf
LySReJP4XLlkhXzQ0Q2ieJr0nw21aSncISFZd2aOpeLnTG0VSn55rDaWv6JdObD2
aY0i7KrcBrqUaUUwKvHUlnUhrl1kzY2B+sGS0Zoa2TeGojjanpzRpx5A02DUAZMD
HMzHnp5kMy6uYTQilXW68Y+egcNbaTx6cd67c7EYet1qSrHUIN/lhwSrsdNh06qw
cAKa5mSethk2WvUrXH/J7W2KpLeg1zQtqwK3fcEm0bX0zcDGEg9x4CQFAsKB726w
bHPxodcBgwFSaXESxUbYLm8n1izMnyI+o9d/lqq1k0Lr1W9c22Q4TkIAPwx4t+2v
jYYZSroG7GNPG/ZJgn9xgEOSnBRNduvzUW06eUkDL3Pt25isTij5qRnQwLFFYA+w
Zb/3ivuDkrJfSNTwl3NZaQh9Fqg9zYf6d/QYWOEdrQv7Gm0zcc8Dzbz8iVGpxBAK
ZDNrpoRm3Y27BoJfbjmvOESdWRBrMOs2qa7O1KkYcSynTpjx27c8ehYSjNm5likr
gvDX8YrtU0EqcOsV08a7A8j6MxUCsD2L8f7r1ux8Up1juJGMO4VXrayOCpkt0X3n
LHmc2nRH3/77rDHX72h0ceZAzV69vTdcaBcw0A5ujdmmn7kGn3kzZspWW6woKswP
dewKgVloiuwzym04VPS/EQwIHGBLZJ4nwlqfMbAUCb1m7KTZtVQXW3/ac1X7Wffo
V3znAAfD+RmqkuVAYFkoe8tLp7l56J9gbz8Tn91uCfvhFmnf6dytsUIjo8k9opJE
hL8ltTPqXc3c+5BjZQ9lnih99lJRBINE/q5lAl2r5DIjIRWs+g1sOnAYYFJckRkK
n4j1A1kX8gQH8WZPdCrwSXWPhv+fKvA2fzFuF2eK62rRIzoxX/LHPuNob8bUW8Nw
lQuPN9uZtXG9n0dMGPJLgypGytikZvbLWbXCAaL+OGILRP9L3eCwJhzFLXUz7zjP
3WnFxzKB8V0OZ6C/qsg/bVqSalsc6eisMbK3i3oy1ju2c/3z9NiSrXTrkcv2i9GF
T67P+YQ71mnNYWhDLdqY4vPrGZqaX19fJHpmZ2ABkvFY9bHHzWBF6hA9dJUl3ICl
AvxPcTy+1oMqdgIsTWbIglXFUafCirUscp9I1NQyXdszNzz3Xh3YwvYsDLribNHh
MIlAVOi9tOuWg6QJJr6XbSEhBF92ZTuehfgSv0ShkNFKP9c3KTbsIqof7emuWsxV
DnmoOOLkF8npLf93IUkSm9cwa10rQlh7bMhV35DYsWuRE1vodVbx1PSlzB7IqBwn
eeMUux0i9P6+LpeEBYWpcZl6QoEHWMvjLSDnQ/zIIA9LcgF+A6XgekjnCj8gCN6J
jSm9DIlxAFeqnAY8m6yxlW634Jemws6eDUmVS8MpHWTzCe5QEU9gsEU+5uIJ7zVy
7GXVaXvFkht8vJLWkFyor5rS3FIpfrNAnm7Ffyr5/nGr+a+WP+aKmvTFzG8m5gb1
46ii7SL0MpZJh5SV9RVBAAMtyF6RZL/I5/08wrFcfKFtZ1qFBf+AOZREa12jtGBX
lK93oX6cpUKHfzC5tMMd1o8XSZmXImoL9MiBENpA4nO9e9U12yTqSIQ+qQOSOiSu
yuAaVTyimOgSXWeo+RaGNEqBvRDiD+HlC6KJ4cNhqEwfNBcaEw0NkD+pmKMxg6Xn
2w5wD4aTUwGybIRLwvLe8bBAf7hzTzHuy0PpR0gSpqpyzYQrq8zQCdu8dFNcuT/m
sT9akTl8YS4UyyjL+SmmxxK/jN353Ds3ap8mQGn1kbldutD8AAoBjaHEFkiQCDvr
ZN9qDSNrPQGyaYVZOnqhHuofSx2zJ6Xd2+0n+hEVpdf4wJhtfSXEa4HclzFmksjL
HzRtGvO09UtgUdk81SAVIQ==
`protect END_PROTECTED
