`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ft0gcIOrGu/Jk+YvuWvHmekGRnvaxkPMhleuwCm5EiHc8DT1HKfRiX5t0WwruN/
hEHXjCK5aRFGMUw+BxQjcusaF1LtvOFr3Ph6NcsiqoP/sMEjml+QMkFlsEnDDAKa
aaumAmMR3mNdfmMkSbWGL4ShsrhGv+udgyCKsCs/ompw85bCGwurKLuLyv6OoIoD
uJJYj9oB29SmAJj+bEwLGURXAi6/3ioonzL419RW8hPULGLe9mtIaAmhtO7U1C1d
q/TXrYmOf43x3eaf69kD14s+P9pmxhnG+ZON7/5ShXm8mDC7OqwNivGuLydpljIp
nuUKmJbb84qyHY5WLHiGj5YsgBgAsDjfkyLWZPuqKyJT4uOKdOoUwkNHEmUctLpK
pm/GRexlDCoBznof0i8TAd+JijjiOnIjQ0rZXbrNEKbOrT84gCOio/gTkMsZUhBn
9KQ2GjPoqfzdGQf+V5HpkQqpi0loRWrXlSan9zYaGyFYWHa+aaz/fcPWHsBtxbI6
Wf9DA8seFCv+hlhcMHNvo2lWlsEk7X7w2ore315OGKYfAKQrrTycEAP8+THjzQq6
VnygEIOLGTYdMwiH0GD/Yhdu+JysrcOmyiUAMPzjHI5yZ9jBNUDPEboRjbqJyOMd
DpHjxAv2iAbPZJ2fuCNn0BbWuAEq9EFhXxeS77uLTf4lPP3wCfXYl/9Gh31vBC4V
Nfe8MSjVVnem54nGlmnkMSO9JL9k2O1dpN5N9m8NeQySZPy6hxT1Ir/HlXivfslp
mQfZKt/S47XInDBAueyzyyo9i3j9fzdyM+j7lRxqUX4zBfAuVGILGYYacpfMetsF
b959DnJ9KAYATfY2iY/ZWDWyQW+sam2VIIFpugsnF75/0zfEBEQGG8s//kW1CD5z
RRNVrg7A7i6WZeQeBjkLMZ3LXMQhEVGxkkaMeVPkvJNgcW7TeqVD7aUBbmNeVLLx
mR9UYqthMXxwFEED554/V4g+SBFhyZKBoTIEYbP96b1ZC83ye8+XOuncWYj7UT6I
5kquNkErH8CGqAM/4gkAlcIHF7krucfuVCQOUtNnerQLUz3vCTq6YgbU0rAZzBoe
+F6dwyJtg8+uDv4WEZvoFFm5FileaowDlP9LT85aCuDzSFCbG9xQsJ+yWiB+eKrp
Eg03NUoRSWYRDw0mBiXbEUnhTrtbWdMwc82Cw0GZtUrJCYEWnDNncPXcdhqDQBVP
BNV7I8FfrI3sdZzmcMBWbbpPoQiGtRBg+Qghqi/5xq8/Y7wnux5fsMvXTxucCeNQ
tin99jej04LXRYjgPddBZXuAUdvKCeiPTvPjqiungn119XUZkOfChr1u/xfRG8wo
m9eq6Sp+KswOvRhcQdyhbRdQuB/CTQF/zUV1sP0bl6KK/E/tJ0ntK/uePOqONuP4
AUoD6t66DbbBbkEJ0eI2tcII/3QOHw2tZVH47vEYXMD6zuDmkJHrYk5yqxHmpBRc
9NskhncOnG8yBeFzkJNNhCNrXuIzm2jqKJMtJ7l6iTvkXQ2ZAHgntcaVcVqhZCSH
qH22ZMfCrfSFR6BXJQpTljQ+3fBq1HvfCb7dmpfEfLi/0mRG7qWX4XNRotGC4cNk
J4h7Ll6VlAYSmNC5KJB8PsOldJqPjZ3PWvmWgZ+OoVm8wbTb+pndc1ygHIVT/xFv
D9iBhHdvzf1kOc9Ykn8JRtp33cwIElZ7UxtzfZeqaLdrisogjqEVO49Jbx5fTG3/
fqaOx+wbBMFp3k1PhgKrG1Trdw4ca3RGBv1kUueNOUQOgqXup2LGHwOsbiWq+7Fo
JuGs31acmCidGe4UTJrQXnCHOwx4Qw/9WjQ20OcxIyRxets+u58+Zh5R6S3lTQoT
ZJklt+hDIl1/EmOkNKPUAWGqvIXDu0+0SC00+zvWQWnf7jBGMIMe9UXwZc31ywWA
bnuhJEbywhoVOdeb5M2QA2tK7fBLpNkMshVqmrDQ638r9cDcT2rXtK8JwPmpasYA
7qPO+HQ8iN9z+AfAHZb5ZA==
`protect END_PROTECTED
