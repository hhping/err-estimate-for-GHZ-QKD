`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cTx8M5UUl2IYxEwgvCKAIipDcg4EcobEhmoi+injBWlq09fGgqNHluQ+NOysjTxR
lmV52sxhVDcxeIHzHNXhPqsEso2i3VNbVYsCwybxI+im4pV7by2updR+F5VR6OVt
OhgoCX1jVR15xicanPusR2wjBubD7vjdPjrRi+Bcb6Pp7mbxqZJOBDJAKCn6hDrL
A5MGcBPBIcD2bXF9UJ1u5jbutpzHWJmfnEPAQstXO0nELQwNCOLDc+Sfd5o5FHde
8GshuctU0xe3Eq443krkFpqo4e9IfZYEJyU4fXBEb2Y2g0Ji0ORMTvt4FWkf8ba4
WZDC5AuTOUInG1sbBGEDgtUvr9tcjaI1cgVdCDt9wpWT0d+/bK2mQHxMaiuGrqMP
nOMdmUNt9S+5xZqYPzdYZwKh3nnzNeXofLat5WqetieyKhyVW/noZchjaLoBiR+K
vVqn7De5P7r6KnE8wamGhwXdrg+me9bv6dRjD8vCLe2jgMLuL4e+s/ROO+Zm8BVi
bUnWcDl+xSCgd0Absfsa3FxfxgL2qqmv2L6tlaI3xyXm0W+01foVgoHJRohtlCAQ
0DSLAVW3LoCDCxUG9Gx4vsFjNYQyQTgP61BtI+Ld0R4FHd9K0stMT38gYoEJtJ4C
JkKk0XM74JRQdTfpDCdOOIQomXpL0Ue/r+Qy9YPwCuLPU0bsbNIee1i3LOf2MZ8J
/dsAVltjPsKm9nk9r0c6awg/Pr3A1vh0uEXv8CpcRPru5Xm6qfmel6omGKNFijDu
kuVS42zWHOFVWlulbmhiJ5f+hrpJFtiRf3TBf/Cy7yfhVKhToAaguKalvWmmnQxa
ypfJz04/ftbHQhpILbLAJ+QlEKIsP1PTIomAKr8HtmJsFCSr4g6LAt1Ya7dw9LXA
F+MDBNjmnuqi9BYIDw8oGOISEswXc0RGo66N0Ptub/pum5RNJZSLtuj3laviAXpB
SqrMFWuaxSeDdWAooALfsvVQ7jQEF3Tv1gRlCltEannizNPLn48R1is7r9kwtH8F
RJv8FSajwARYIklv+XxbabOp5h9o8QkxchX5KHtteXY8ZDEQF8XcgD5eWfgNQZgj
eBL+TW7wcqv/bjDKGOutn+03bS91NSBVclyw+vYcIZfaBZpMYoOM/bXdc6HnW24U
L3oTTy4dqtS2ByilMYTXxFAc+OQ+CtusBr3kpOKOy5LaJzPrb7m3UOHHRCiFQljW
7ZFKQPdxrjmUiSawjlLG8NNKjkb99LGmJha3oMnX4CPmyJuvsgqSfF7lNj7TRnRW
7wDe1S/aE4bJiMUYdet4zEUscdtcYOqgq4TQLQGg+VA4KXLjVu/WS8eUAShIJKz7
6CvpvGhqXObDo63cZ6jYmqTrS+9JxAefvXcHiIJ0tkwvA7YkkrHWiCOHqVclXkgl
FvipJi7o/VW6rq5TEPT2oaajdD3lqWBuFqXJ8inPyttlrbgxT4PgvO+rhgd44eGZ
844Y7nh0bAfyMvN+31X5J1+Y8HJwwTpaKdjAhmUJ66wIKTnti3yhqwcwiD8Xal4n
zEf3CUsHJ3NS5xJtWSS+EVHVTezTis65lR0rr8bwf/Y=
`protect END_PROTECTED
