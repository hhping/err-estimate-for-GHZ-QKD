`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
incOm8ajELxbAmWsXLU4fnoxlmYCC7q3Fl4bUPfedYTNujoIK1yH3n3fq+/tcXXo
z7t8vgWgosLhm5qHsyStbr/vtiLs5c1qDRWUWCrUh3q/k5IUVhnjrSR/G0bdHEQ5
mOY17ILnXbNIbtlEZCziJ/3XvAswBcKdbSiIBWf+J2WJYOLQDs7ZG8hl/FYLcUjI
Ba5CNcyrMBABDZ6TtEWbYvCWQ+17Ej5vveFe2wPKOYZdVLSCdiOuQzY3DMkIah1d
XV2YNZZpNrrfiEBamL/ZQiJiYPBMxIe1zkzRIBUrUm1xUbJ1szoXckiErAZlseSj
fUu8tIma2bZGyxe4OX8K1uFAvUgxtrAY+7fUD8sjJtl7bgj8ijuyNbvhCIK3113w
iI6F0SaaIKTUraKGeUYuUjCbGyDKGR/6FRWUaczGThpcqW1p9JydwJKQ14GVtBmr
g2gMYZ/hPsOSJPwuoVflx7997LzTMi2Yj9FAG7U6zoNXNXpUOPC20zWWQJY7fGgK
b7M6F/REYSirHa85IdUn24MHurGUWAl7pmrtYv/9/6+dImEp+03/y6Kd8vbXtyAz
lT/QhhGBPZYFbnJAZiu7QQ6/oT7ztDWvA9ccbu2Qj/rjw2QiViXM+l0qOnscxRaI
vdh3BXdY4gtQnmHlF0UNqkp3BaS1G+vRMIgWGI6y1bH4JpQHVWVklR0xxJtETlNx
GpnguD+1VdxKxz7VuHBW6AzRZZ/nIWnFOziJMDlRgxZWRbq7ComYXNN2cTfyDus4
2f+/Z3rqdRkiExI6VXeUkzCAriH6huAaMSKAM6/ApPNNQB61deI1JMzGtQvFj0zA
wj3uZoeX+i7cSC+tQPU56J56wyPGYKIOJ9kn2D7Ihs39bK5lMommTXlPP1yMXSRx
73bVVq3q16uIiGVu1w+vzVvlNzFAchQx0rHrw22tmWxefo4ldhXbctWVzWjB6ggr
TIcZICOaia9cUtWrdQvHfb8CIoDHeghE5frVqzetF8bvHLySWReSQ2nG+y9CxPUh
vYrA2cSLm9k/dou1apUDx9LRsambP5f0dmzcHhVNONdcOE1YA0sa3Ul2hDiNRf4D
Rpf5E5Z5PlU6Iu5lQTWmhiWkfXgXvqbgOrss9CKikNy5a59triSUxdnL8WDBY8aV
C9YEZ0r905HjBuYCXGA46aOnaMRnab1cB+eF9GDXzjiKoivDVOztryJYXWXy83UF
zNZc+ZFRnSSkiTDFzbhDmM+WTxp6vfWmXrJCsikx+j/W2/yHNOxcyefGopdr2bJr
fNAPDGwS1eHkWG2gX3Sq0yGxumqFdUG2r9HD+3SC6452V+WWEWHlG3+Q8t2Z7ud3
y9/AGEdeFR/lRsq8MVvWHW3OvqJoolJoTO0PGn8C7jOMxfk2CL0AmVKdZWeutPUn
+i1noTW5LNEu39EyIF2/OXa6ObsvT/SIGLpoC77hNBBXU9ZJCCR3V9m0VN9Mv5SO
Ouxvc2rbxG4jh1pDoAhqorjWsCALC1T2bviAOJJERll60DB1WLhyGbhXwcoN9Gej
HaUbQW0tIY/74uEYuVT282vrbSRd27UyZZ3b3J+Xx5L5iDHqPXbwSmu+uCz0Even
8jX2Ma/l3/RatuKWP5ogHjaoD1QyQCn+a6kfzqhcx7eYHFIgL2TEcosjZUOCNtbc
V5dGXSb1Vzssy4RT/NuPvwKTO6inx/I7AEptaFg3eAM5luI2WfAS56D3Gx2x2i+Y
1hGLlxcQljq/j1LZZDQDxFJIwwzyxgPfTZFrzOmzr940RBemxj8Dj+t+CGMVLQEE
l34uihXmYUjoC2tAgsjyrI8TyyxrLFGnpMaz5Fkwgrr4Jx5i3aa0rVNkTfOrI5JI
M2PnxkUqaGyYKYMalc+fX4pF1u9Ud3Cq+qcSVDZFWzXD2aIJ9Z9nsqB4tAXCVit4
m4j7ogPcoaWisY4yWcVk9JV6FbY4uVsMBIBt7ADN5b3t5//mf3lKPpunAzdfYCWQ
7GgnP6FnTr3uPVLRC+fD7Hhu3fnRzgAwEUSc9uY4lYAyw+OVTFFgKfnA1KPQQvLb
IfARvEaGj0wL8GS7LAxM89+1IK0G2LZlhOGZdomVG2C1KwbAKcg7HyrmNiIcA46R
bUMXbm2GOHVMzkySYojJ9YT4BpfnlZMG9FOe4QWPt9as8dvJmcGbY8TrGOZdMUE2
DRvHbLKA41M+wm3vXQBrw5r1RisC+5mP9Uxvl2gzE7iJ6n2ggiuJOJ6hfaBfEPbm
6raWYaRTpnK2MwLBsjeZgfJPS+LAAVoxgaGPu60udtRf83gG4ko9L1i8vXT/lvcz
rUuUplQyRDBTeGfzXo95XpVQjLc+ZGpuMlK4hDWKJyRsVqmspnKuPU11yjc++uCN
scwBaD9sV9ttcmSfUjNa2OhCQ+h/0zlY1jAmtKhYM7TN9gMPwP04pTPLAzwfmyiy
h2PHbhdLvsW4voqVdQTMAtLdDD2CXLKq0AhYN0oKTmhLVvS05v5WTWSiGRFU/nXF
yVpiB3rRBxRn34AKzki79Sel+52NOfn6o6jD+pTWHOnp5eSNE33ga190hZQlcufR
AstFIqR2S35lc2h1g2/ZXbskZ4Yts2UC9CzyX8k5AevR065ygt5jURulfiABmJCn
J883R9k7bJyf1HgxWND0KNZyudtK31Usfz/kB12Drrz5/MAA20qK7lw3B9paV8k2
k3N2yVvqujIrjuOwqL3lwDkewGhWu2uiYMtjNXMvW4GI+qBTCVQr45HB2rkjhQpG
TKs6fLBTGBU317+3rLgmQrTXvg0Iws2a2ni2t85NMV4jsNoE2Bh0jK0Gbk48jd/S
x0yjCzDeS7p8/1KS/E5MWklz3MkRGCrMrMtP9+j/rBtkRQ3lFBBCDaYN8ZIM52qZ
NTd7WHbL1vb0lA/bG/pLIQSIC7qwiGb03us5AAXzRWtAh2PsBuOFfDq7AQtfCXi/
vLK/j1k8lbwX/NrT1ad5YJ2l6EVbT8WvdSkFw3CZJCMzx2tUX3gzEQ3NiHQvBChP
AdUEoYhdEVK1hsQ/bJekoJq9xwipEy2GmBu4Dfo9osz6ke5/idPZttaVMZP0Mir1
xvAnBpzSt6cuNe5e8kMkT6pN7egwyQD4DT2WLeWdnEcxDG5l+LonswcndTRMLL+g
2HlGa7r5gUF0CdS8RHRaFeMFw4UR8n4bUK23dbz5iRi+OGQp8W7Gf2VCUz57ALhy
uwNp1eTpBNYeFXByCVl82KJv3lBdlJL6a8QTbM4UUa6F8stKaTnDL+u8mwqI07yM
RVTeWA06PsqVmSrz+je4r6XdSBTbATfC/pJxYN6nbBLiR+S+99IoZvA+qTTu2LSF
CVYOfl+fO33wvFDAVSR96vEI/cGKW79e64FRZlTLq1zoSOugvQ1eOkOAgaPsynsB
S6X9ikSGsXOn7RlFpiBB9VTdIfM3uFPFVA6XBCLQjct2hmYbKWhEEWMevR6slYxf
Uw0Ysd0JaRh9vPXWYXeZ/MPs5HSM+XkpQ8Mu9t/31pQ3luOIw4LMain0A11Kemti
/wTmM+i1KRosEXpMlHuuCFVSPBtz1P6iAUnHIh1ufhkP0kSl6P5U7jzKhsfb5OOG
vSDNWqje+XJKkv4/cKzzYatQqzppeTIhXB4fDkXjpJp7SP8xehVKs5nBTxqwPArx
qRGTgERi0p1/P9IjT3jVLUlaSsUZiLCgIc1SjFt4yz/MMynHqWelw4kTS+vqo7OS
puQDGRx1vDZduNnM26T0ZnGswX4T2DNnzJNgPQOhrr8KkmrIGwIRQIW+9IcGTmex
P/wOQEtEo1SvLmQ0IQEfVoqhz3y+iP+PTuLMxMBXrSqzrUHPoqEN+fqLOcxsoXAU
QnEhEHa+vK9HY0FeUHsJps8ImUjeAeV8Q13Iywrt1vNjdUJCBf9kkifLF6719mcy
MWVTF0Z3Eb0YLap4rmyiBx9q0cNL9K+gYnqznGkn/VQp0KOgFFRCUGlG793zj/Ol
2x89fuxRH7Y1UXj2fUN5Pj6nixZM3oDn71ScnxBC+z9VRLqDyPctzULuaxhRqFD/
uVZTC2tKKLCUKCaEc9XJs9YLci767ll/JhcmjdqPkD9/L4omkxtyjnulvFiLxOEN
DBIJv5QtVrHjZ9qOh+ywhZNXWXt2vHpaPmRPJuKQDDUhCTkB9kx25sV58zgmVjSs
L2E8kUJD+kumH8lq6xF9qwu3p9yC/nm5mt/i+N/M+HM3Xw26lF0gUn74uezCkXCs
F++hT3c4IbqquXWZetugXbjuLqi64N9bSQ244AL1T1hCnpYPlkWvlRw+zkK4scmw
jCIssGXg5Iup4E9Lvq+LNMcE8VV7bS5n9rB/H37PEYegUQ2WB3Mr0iwjZ4BXd+HI
OFzFzCfJW23yNI0mnwDvHnP3yk1fqK7FpLN+0hsOTS/cGrpth9cJtCNAw8XKypVu
6laKZHcwb1OvQNKDRdB6MWOuCjvJq+kl21KYWod0BjqdXsjRr7SVgwgDBKqAurav
JXvq/h9OQeXYylFipN31Dlai0aQ5Gnpv32JdMZkKTG+QuOJzzHEbBwHd7tvJiQef
rSck2/046N3QRRiEpNAhUqrUCs85v6KHrnOOF1+qZKErkip3KjrmOlioM0X5GZ3P
BivSEovWO8/ANSwc0/yR4tS8jwb9I4gqs6yocvmjVCcCTefo7jOXgzdYRZ/GAfeR
ZUdxkohVVgZNr6L7oBdAUt3G7dya6cU8mEyzI5xD4O3BOUk0FwPI6gQf01oS3ZFF
tRRjcUqzmWopoMbf6xpwwGsBy0XdtAgcqiekf24/6KKUJa3ANmMQkpyEv5Bw88XE
c7U6egYI52l7UeFjTlvih029HiaUbJeBbWCu3fHs2Q6OzMAYCYazAxeDq3wytIqy
9HQHSrGNAmkFVgh2lc9DvBL0LLmNZtnm5t9M+qZPW4dDSfS31ykwAwNmmj+G3YRx
ZkKJrqCiJ3umOSuhfpiCdd84aZOUT7GjAZ3ynXH0rWAMq+a6bVC5LaGR17p8GBw6
ar9AIpA/dNe1jS+S8qy2YNn34NaZIriGQSUKtbV60e8Gf5yRAmuCQueH0Iv/yf2P
AszQJ6p9aHOjoZyeQ9R/r4bWdqr7ZrtOZWQw2dhL31SH3zJGLyrPtiktug5Ybst1
Ed5TeUfiBrHK8wZ/P8tbFe+kl3ipU2HyJ4qsMzhawVJ1EdU2nu27QjtRm3kTqXss
36b5536PM6ku0E8UQzxrf918dTJuWpDF37RKagoxxEMs1+5DBMzXntBQGAqI8slN
jORsCvXAzzsLOnaJ8p5MZZCQenRDkV+NZjLpm2Z+Uo0wD2lfYatKKHzGpG+2PWgd
57jWGv6ov2nIuijTWBerVHj/2O0BZ5Yjou+DFUNJm5hY/ZPUXQFhldDrLAD7Gihd
ERe0NylXivGUdfHOPF/h8XYPso4KthooELYEKNqz8uUFoDP1K/GUsHqgkJhL1cnK
AqsGu/72Nf0Y1ZKXx9YiefMp1cZCjNC/BXc95uHPPcgD6hALj95bsRF8EzA3BO0z
d8LRbchoTYCPoUNohpDZt38WGQJUeeUFlDOlWvVUyYa2j8nDkgVWCDKufY91bfB+
806cFMoY05mAHeQ2NXDlBOzsKlgzpWd2i6JNh7JjguNz+HMm3t0oPg6ZvILgmGyu
MWiragG18QpLhGY/lClVmcm1gYYjeECmqvRJnbTEcm3TtMrQ7iGSjCFDpft2P/ak
GWWkX2tUqsbFO3rHgbdH3BFIdyBpdlE1UD0BEKSk9V71f3npRD8k3jzPhw1iRRah
DZyRqnzonew7/GRAatqtaJexa8OMKMFx3j3qO6C7cq+OabjDKr59u3LIemT+2tyh
SL7voBZnCx/JZxBV1o99nRJMuVzCV7c9NveTTHdcFrul1T0QvuiDrGojDfEyBjUS
3JvmAnfrHmNrPHhTXysYH52eSeDiu/ZQQ97LfRMkKgkRejvZgriVuPhg8ex2hIup
+U1b8xfJgAde2DQrv4RZOCaaCaOlO15XIau0FTrEpMel8kJMnphW7oas/1t7Ixf1
GPEIQi7JvW5wSl32FX+QAP8sXsEL3c0mR5YKWxaO1x52uaLNbnh+YErIDBnDmc2g
lBjwbF598w9RwEkEPU/H58Zf//9tTUDhtLh0k/KaQEwuv+OPHbLfPIDdykaheLsg
CaTiZY7gDFYhdUeA9Ejk94UtCuRT0vbsZq6qymkdfaxQvgGjOYVAsumSUW+VeQjs
G/5zKMjqFbCKLzfM2ktLJz9NDQ3TwPrFZrPwIagm6GMok2IG8sECYOiJhqbZtySr
wlZWBrle3ozvVKZAt8LoifnNDfdLZfocroyRHe5dfBFqvY/AmIXwUUaatYaFJvIr
1vsoeuoCSRrjaxGBOOdnqWH+moqaHR8UJ4RV6PA7tr8vg4LVGJZgXFb6DkJ75jQr
bx+22G5Wg3hItNQUaR2fheNwd9OuUaadzAVA4j1pV0EbZPlSngrsbho6Umj121CL
Ui6tu4dRXjuN2VsyAfwDG+zONhZGjkDgeOGumiTrLh0ojYc6tLhmX/ZV2fZY7JkZ
vOtUmjfruuOBrBgI6kjhegnAj4gQqJ5uOyXDa8OgiE2v9Iu2qXCrxC7EBm780kt5
7fc/t9w/QMd8A2P/bkU822mRUaavaRKH1TfRRw3wYJe0hKfucVRzFAMbds5VvGQw
bfeb6dT2kuHPgt2/t4HKev3x/W/E4kMcRTEr6io0MNsFGL+GPBND9Cyv1IO1BwQg
ZaHGV8QhlZvvArwvyuwncljdhns1gTHVGt6wZNzHHWI9NLh9Aq7RZ/JGhUTZJN+Q
qQ8H8HQnqIqrdS1cnVhAzvEtuNX2C4CwjVDZRCouumBceDaJ6vqG40S0LorFTwby
zDW8e6Tl2Wz2zE4eolHEn4E/JVf4uhHR8GBBa1fhz76gxn76QWeUrQpO1c5B3kvk
b9auNfPuEbG1oTpqVvhAjJ1Q0SWB9k7G1xj8alhVEVDX97KPNEyiHrTMX1A7mKg3
83vP83WhtY2llrmjtjreb+qLOOP9OiL1r8zKPSGedDyGpOQHtTYtDD/Atf002AFT
L8hqTzyAvXjDC7CKeu9O+RcdqAOHybfzv+5ct0GUhvWn5xrF3SHXNNqhGBi3O4wm
VVpS99+KoylYQN21dJnvjjgZsHyvLusmvbt6UimisbF7QkzhFdtgRjQgKdI7t6rr
BxBtb3Zkc8NHMzTmgUWiSEJyS5/huhvhK3eM5XbhbpZ/uAg/45/QQGypokKXyCNj
dUedF/Uk56ystMBkw8XGrq9st/PPeqUudjWjg7/8kce0W3Zybj4MDQ0BuEJ3n4XB
y8X31EFq3gyMJUytQ9TAW8xFmwMu3ayQwAmqPUd5S1YokM0PJo4HXK7t8DuxykUw
4GfklOyubbdDN9XPSi63cS6R8ptwXmJ4cOhFb4k3haKztgBC8dNuPxFSw2lgXydX
tBapDucYZOmhqHxPmd6UyyGHP2QZ3Kv6z+ojJckOH6grbEC+8lw67Jr83H3md2dw
M/sD0BSu63p/aNqNdL5sSrPG/Kuc8jCP7N32FMfvBs9Z4z+KAcpXMcLc3ONHlqlb
OGaFkDXAJ4Xjwqkdj/oCHJEpVFIqam1adrmvXhvMz0TTt7V6HO0DcAhlEdxFg4Oo
GDv7u/8ytp05IRvwxaCcxg02gL9snjHp35Eb5esknne2vB2sWr+KHB5ODP2ZHUfO
NyUVhW2Stxr8MJa+ECAkcNefVTC4uoWGILittYCJjWt1spNEKQrGTMyPLtfGRh6F
oHzh8Main7o4jHsZjyWO1ToaFuAspcrDIvj/RR6Sl9Xu510JRCpQ7XCruRN9OoEy
+0mWsuV+CRCob/6JZUHwxqydfXsQ8CMb+dCm5P+PV16Gw4/BnEwR+Ff0Hzz4fJvc
TwzXA21g9XGl4CCSw5T3CfB/NohokwqmUakS/m3NtqSs1aUU43NAeORW32KK5iup
n6xqarexyk0l2d5pVeVX9d15NxiNZuFlGSGd524A28TtETfbq1S/FUzE+OMXIdbX
Ld5l/FPB4iJIuuZh4IecYKulLUuf5YP4HmtlNoL5MGa3x2gejAUu3lzstEDOC6uW
Fsg03HrgLO0clftxYCwkRARAZ0T4PUiAUjr3iTYWG740jRHISMu2j66x+RatnLw8
NaFB4fVowaBcGNwGa6yfd8PPn83VKPv5OTyqBio4JZn2TWX56dHDmJy3yvMXHDHe
cAEx0Y6zx7o1tm0IX9RmLEUT5ST4kDAqVjPqnI0LkPtZtXA9f+nicoi3bYbDDvvU
kA0nOZ6B8X1ArnVe1vCeNQSqRGetc2p2bOyopesQqShATCsVXAF/333zJWWTjh1v
PAG62OcVD4eOU8quMUyiVOuXhjVgyrvIXSWmPqAacNmDlKL6m3Pp1J4GeuGBa202
WgcohHWmQf34cBAJMsqG+i12z5kXhPsjW/k/5GEAs4mNE8QbyO9UBmVgNVmOfix4
o/x1D/WDB9YHoVu5bsdao+21KYRDtDBJUKptYzYkYua63AYDKUKgY1R9RBdZD0rd
2DaNddc3c/NDOhGKBXU/delU4r6BEhdzJ9ApNaVUf5rbGcaOkU4duLz+CNx6kMpn
5AZVYHn7O9uYw8RLjukDI8mklwI2zI6bMawY+6kVYraf5TxF7GBlK0CVZDNqt46n
EjiAP8FeqzecQmxYraxgD20yLIa700MIZxgTbZwzOcShgX0SeoDRSY3h2AkMk1KE
wUP0na9T3BQ4CLMZoOpnsXKO1Wi+nxEEA72CqefMd5HgXCgfhbDWB3lpWCwIAZO5
C73NsOJt16R0guYjv0mE3FXjFkaM7AUCS1SUReVzO390Hrwgv8l5fIXZ+MVZLtrO
UCNncBARpWQsJfJwoolsdGEzszThXJRCcBi0T0EppX9SckZFIFUwSfCjBgfkyR0x
aVixi1Ktl4tRAxvf7JpMBN44QaKWzPH49jQxl3DHbi7yTE1JGxy7SjbTY1D5ZVa/
CAwwaFdIQKRXyoegj/vUidlcUKR3T2i0NZLiJ5JfM4QFu/ELlYzl/u6GND03CkLT
qsc7fYbAFbd2gsW0RxwpRDOSm6uYhBc+23YFui7Rz3XMKZ9Ait/PIprn9WvVmjTS
L3jpYPFExXRcoRLfNtITz05S0ywFM/sd1N2sMdh7jgxfxa+UKMVQeFZgUm7PS5c0
mD9jIf62n3c0tXxrvl0GmFEgq/2kAHnaQbWerV2RSqeqrbck3AKHks4N5ovGjkcw
txqKZBPV54Ob+ihz9LZKiCFZgCrNWl1FORgw210VTvQE1jUmSpxqNmBXOJO+rNAL
a3sq1N8B3XGLIGRr70nLPP5ZlROFiCiKE9YDBffIDq/cL3s/EnFYQLY+JWC3itT3
8M4vNOzFcHPkCyP6SQTEUetN6cycE7ho9fQRRg0xYkWg6bSjHZB2ywavTFXtb0sm
rygH/kYDyVdlF1GteCSVjfq6Mc8cKFiYEx0FRDzOp5AWv92hU1ZpEsIC9F+gyOXn
DmKEeSR0tIViSlPMYbT0pFk1QskETQbqb6bqxPVk2BbIb6VOEy6kaoNcr4G8oCdi
06HIRO+nCcbmtuczZBJz694R8z8MXvZqBMY37euKEGF4bODIqBlbvf1QEqvDPt3Y
IaPM82Z/VkSsGxaTCifxmDBqEyagELo9dyrUO6PrNkQvKwoCJYENYrTFJY6/Ojxd
HfpR5/zu4CWW1uyWbCdw2ev73neWOdhaOTY31Qgrve67ckZT8FU/wEZnu6T64nxf
2Mozs4Mc6DzaJJdDWZeUf2Ev4tJgcsdJRw7EC9Dh3ICk3zKS+AP+IdUS+z+yWZ8K
uwXIoYe+RQYm7WXpnx0MoKseCDxGTtY8f/s71v3ABPlc6YEkhjdFU3lLsncZci8O
5oUfuL/u/H3C7XfJRpXM4yQUenuJONv9fh5Uz/y+5set4hvMzyIryFBInn5oRBXd
AOh7/7M7EPN3YXgXpyQKKQVyJGbSrpMB7SrmQBObdnseNujeFh9h6Ra1P4olX1bM
7jtFWLxJGkGQ8RpwVaH5wP9nuGQzihQib3mHBikWlQd0l/IuNLhBj5VcRaG+si9U
2sBKt/gK1GwoD0EsBX8srnfKjFv8ozdaYXsi8AyiV92v7pHh8GgiC0ZSTF0xUUZ1
6+mmkJbU+2P0duL0rgVzGodPH3Ai5r58tq2mnqq7nFiiOWKoMNERX7MD/GWkRj6+
KsElXzvDSx9MRdoxzokPLDFkkM9cZst2SbhFGApDyyA1KAibdjubSMbi9gRIXOrq
QJB8u3YCaZKNEJQRTBHBY57u8SjD3sWQ11DBRGaSS37YO1KGmGRy8ZUNHpLwl4Jp
RhO+VjXckGMglMi3D4C3bnhsl0XLOP+RiPG0TKbzgDZPJd+/19eIbZ8BGOLznJmA
2e9zsGHQrwQNCoOm6UEkn891ix9JvbkndV34XEx7lUU5hWXhH19d+XOT0NPMvdlm
hXh9yqXkEffHeh9Q4Z0eH9BxS2dsK3/pjfsu89YRMR635I3F4nDRQKTZD28qfZml
mZNVsuuGX2u5QIFDAokVSb5EKKNu5d9H4Jf3ANeO/1Lfp1oGAIJyPDqGcwI5YmYp
AJ/fpYzY4WecjbjyG7eGyc9ooOma27G31tQ/M6BQhkVMbgQP/dYwoFl6pxlQd4MF
OzObkgLHJDah/t/KO6rSkjyO0PEMYU13RBPuNvy3U7fJ3SXInxS55tuZdit8BZt+
noygFAWypfn9tqlGl5M34f279JfLqCREBTRTO/qL192fQkOdpziU5AaAnNbvghqf
sV2yqNtspLUvXg8hAw2cnp1Lxv1UgPOZcqrkyORuDBfYsViWm8ecuky1AcyqToF+
0COmmeJ2gU8+UBTcu8GWcr9O9vzzc5Nq5fs4npWsSmeV6wZ7btGrdC0tCyBPA1CQ
gS2kCtd0ITKq2ftt6Fjg19j2IBZxHpWlAMwYYzicl0BEYX3cqWyRpAlaK17uhncV
k00+cvFZcmL8vo6zx7sjWsodE/5kCt283DX88V3GSZNcH7o2GjQVt0DIDMniGMpF
wj86vJuaTn4XPhH3lkCmFhpT0S/mpcjlfkldXY/lusR286eLzAPnSYsR/kffdg8R
CZx1FFc5dOXVI0EDFXZFoLF+m0voXeg3lhr8HABPAMc8VBQNATrO+e0f89Vrds8l
7aIqxLnbT31JYDTsuttPDcKk7Jd5VWOuC3jYGX+sCsrpldBv5RCSR0UFlVN1QLE0
MSDPHI6XbWEuv9h7PTvzaRSWrAljHhhamklEalO+Rd0fo8ArLAAV0kWPVZ8Q3STP
/Hze2rsxCyW1kAOQ9fN86YmFug6aqf7dLVPZ/0E2nFx7L4I/wN6xozS1+ZVgENkO
Ma1H3BAD//WlvARZk8wxJ0SbzJO3BpT3XJ4jlMx0JWxf/7UC3ez/xVv8jVGb5397
yK4XvV9aZFoqy6dgUUpKoOWavd4LgAfDa/FmjXsCyJQqcq2fPRKsuc0/hr7/7qim
3wyducbwHEi7YdW2jbH1zp9+pKbGoIUY+V9BH7DNLthPxh0Q/5h6BL7RXG9VH0FS
dPC+xAlh00OoGli8W8tcqtH7mGm0ShKl+dIjSBDQfW1Z8C3aZZvnOzJM8/XQVb54
pN6sYpw9ZDsYlx+M5dV4Y0QDogO8XsU04qbfke43FQgEImuBGXxujYw6MLCICPt2
fEAMuz9cLmp43Mfl9Y+sxqFxyjX6DsAYuj4AwOnt/p0dhJlCD+8fwsya+DPEQCJ+
SottxzFmsnPMPI0OpgNoaTiaCT08N4Coqxp0o9fytV2kcGWWk/x6M24IWhe3AsbB
EguQr8HI2SgMJoocn58Gx8RgEN5U9yRtPmJeOBA1jCJWI3XvjCwUSWClQJcOFuKi
knNxAGkhCcAVC+b5nqJBfIEgFD8U8Um8CTo9Cv9KYAEBQ64Tpu0ZFMgVXXQCHuNU
/WVhPw1Z2DqJzReiRrpPF7vM2c2brTdcBupnBKO1GG1hPdm2y07PBs/0myexLXaP
vJwm9C3HbsQvji59dbkmgbICUEYRax+d42KMhTMyfCaxsWiLNHz7nBs8UIQtWnj0
Nv5yrNg+GlE6FunpGnVtSZEm31KTH6SnBD621e+D5ntiLPBVOBSMaFEZAMsJUkVA
jDXf9oqcBy1I2xujvsvhES/vWfilGmqyyxuti+DAa2sgSR0HAVY37OFabYhcNt2B
LNt8KEattcQPP9ONFJx/1GO6DZ5HYsPM/jE4rUZ0Y1qjnCNm7yTpGcw2KdTh3dtu
ywwE3hjqPu7m/j8CFpgCocw+B3Zg9ou70ClVsChq6d8lYbom0As72wWgX6BiU4Zs
PI15PdYoEJGk4wazjjAKz9M+qY3IuMvgXdYkJEjMpvgMMmdlT1/5u51U8oJbZbFf
Njg7pH6EPhlkrPe9nK8b4RRlHWnZPiPJqgEo5w9kgK6quvVg5n5n++zg1Sc3lItD
OBhYXKguk1bMqa/BQENAewIlJI9PBWgswAMAIB3eU+xYGRSZB4rXDAZe0lMIuBBX
tujWmhvSxzYNcsWfCOysthx/Ubr21dSoyR/8Yi7mgNhkHNcnqR3/ylLItqCoS/Le
GTdHSYZgoqQAixAf0Q9FhFQV2WoB5xwVPc7V2wDfLXjASVZXXFWFNEI2sH+usTHP
DIqeepfjPyogTZkMDKoJlqpzVV3rJg5zkInMyzs38DhgZQwWTXo8x2E1ItrKwcWm
4GJuNc9901l/WFhkkdI97aC/dA8bTvHVwjVnEbW/BukmHp41cWC6L/weJ862eiob
E7qMSxZToK64ffhYPBLbIrTLOsrBb3Z+lzsUy4HC3F8gmfwMSfsdpp/XyyaRye2e
l1zh/YVafM3feoyzwLPvJGJb4TMdcvHpzkgQGdQM9CnwQNUFGhgrKMrc4HWNjZA8
VOzlIwhVkbmh0zJS5aWZqzKp5bG46tcJ/tzOKia702+LibT6+53RuHKWsTskcn9c
/DL/eioscBgiVvv7d0sfY0dC2J/7wSyzz3llqx79T88ASslAcCnfYWelaxu4PJ/8
RZqkXyluRJ+CYuuL7dtxjVj/fYdMwS3rJoXgHnqpbK3yefAHmGQSJ0UGDDADH0yY
/guHe6BCnGbXp2eo7rNmQYWciAMLKSU1l/foJZ2nSaOgx+GPI2J6V80RoXbpxVVm
cLNbai/orSdIt+XvTo4f0s5A9A6akqQf7Gj99Ma7Xq/pYgVfMSnGuHPnl4gi61Kj
G+IvGoNyx2lHeUCHzJZemg2/jyYpF41CLGhcuMrMRGYikXMVboFOV9r/59wIqqUP
q2O6xg32RqSmfsuxcsV2s3KVA6vAo45M+xktzbYHcwkWVTehn9U1Ns0JRgkJ43Z2
1J8WbisDPkDEdWTTrOKQ2zR04/l8NrkEczbKAphKynzYBAXVFh3NO4w2r64xx/kr
Xp6fQQ5pZAIMyRCt9xdQsrMagBZTJ/fiBNn5TQ8kN1QBFudivbKorbxXkbK9N4hq
mJGaA6qWpMQg+MdVkU+6lbrOAxTMuHJFZByqe1Qnya/aYf9ohtyDHW4ZbTYf9up7
TZH0nTBYw1O77a7ZwuNENgZSZIGzUPaKrlTJe+dhR8L0i20QaurtvumID3mu2GQp
qIIm1cr/bnsGA6W94yM7qkN3LaceiYWH9hueUN8xEocYMhbzoPkr1OqzqifNAeHq
O/4eFELV7b67PqrjD5kUgbIuabfa7zPmyLzYUpe+fbuTOudIXMLIFjZH4/aWKn0z
O7KA6unb6jGcBMz7OU20/R0NgablZybBnxYdiUu+7ANF6OnTZERiQROIMDN03CBC
bw1Cziq8QLqkGSnMNMfG1xhwdFRwVgV0BIAz+RYbYyFrk3gGo04wFrUYIquEGuQw
TJe1S7TLPmYNzN4ij7T3msBQo98/B+m1i4wfhIgOyN2Q04I5Ed/5+WAPCrHkTFmp
w23raRcOKgR8E28KwNLzLX+AbqELG0gmLCzbNrNkTQxApb3hYWCKXoZttcLc24L2
fLBnBMuOkxn8dT4qp4ni3IKAorNKRd4SNw3jHW+MRS0pF7aInze/IvqX9BAnLqFJ
wpjM38CXlUMI5/qy7LCmkKsOtNWkj8YLDprLfKJ1+zSlHK8LWsIWK7Pr+8lXK1nh
rW6Pe6a0w/BnUHXt/y6tP16gtaxD16aa4Ezs1H5BOr7Rxj7iCTc8+9AhxsUveO+B
K8rZNud+yj/7vHWyGy88toQqFprS0CFPCdBdwKlzzCbO39Jue3EtGSAxmMvM+ciu
8YexIzEJWGzw0QlNjsI6PYmDq2UppqjHGTy5oEw+68fS9E+SpntkRY+V/Y2WnC++
LUnfrBvHeluO3byP49VOz9v6uqWT3vjrf+EtGqkwyONeAby7pC2s8f+0Aud0eZIi
l9cMr83SquxCPZEuz56JlB8pQrOPtT1R6TvU6qXFNW77NYkgwZbySpsw+xMpOp01
Zkb9vwhNKl97PLjd8Sl3gs4N1eiGTvPuk1hGwJghzMmKrD6PmvMOVYu/wVe4Raao
c6Z9g53vZgygZyVtINap4G0wfi1N/I7cxEHDkVs/veWKwmb76kl3MY5+Fr1rbfyQ
IlAKo1SXDbWtrEoI9w9vjlPPuCDR9sLCn76haxWG37gek0+iTYScvnb/SU4tFV6x
Qp/1QDJuksk/Ijvo590pfrDxOUb00WGYGF/QnKI4eX2GIlyKvWKEV44Nj5y5vn3x
bEDdWmMOZwLwwOoXmKQsrsabIgu42oiW1Kn+ZOkv34mOaajTLp5saUFnut7agfdM
QPkfL+lEjx54uNO+cGiDZUtOacgPodsA7FcT4Tn3MMQqVVrHNE+/QskDuLHUgQyJ
Er0eOIpoecTkdhCl9NauElCazP396wI21yl6Iw7S6CvmsnJzCmLSG/yD/VmPjrsL
RRFL9BGUqGJdde72ugDIgEvTAwy/IZ6k1q2VPkd6FpZ8KlA44vsl935vFy/s++Fj
rWc43zBkt5DY8bwLZrIqvBUUNZ8kKjLblHtFADcoKAxCtmeZ2VLHPQQrKNi0c//b
t+v8rcfQTrZF+UiRPjWsyTsI1zkEFU6etSuUxfFmJqNSxG9lWFJKIAwOYogivWqY
V2ZwWEX+Zv9soiynIrz28VtEBdb0frL0Of0eTLExmn6UT0KSiwIblHQS68mMEc5P
Y28BhwC19Mu13hYFhCVPSbIfCNwexA70sKOPU4z+Q/th+wNy5k7AyOfr1GGDBL+e
6kOsM7NcmEyyT1ecipRLarF8SNVK21Bfrl6id1lpe2EGEdZhHm+zS0JaEzPCkMHn
ILRzd9TuqhEuw5UEgkNk5pCDaD7Y1F2Tzu/FKoTsn9Ko96zFbFI+5VsJD0cExImw
KydET1d6mnyZHnXlq8kQPUAz7n1FUlQ/aVr+qM2rc+KzdMO9cBW4Bf1lO27bisXg
FRavSFQ0XcKYEIUDtzTrNYoIa+4eURMdO77mB5IqCa8edmRQt1BqzkfJaPTWv3Td
HYXCdH+hCn89Vzz3M/4Nv4vAGvy6PZsZmClxCw+DSS2g8qBF+95Evcb1cL6Yeosp
jFmacin8uEFbv0lqmhauJvM+6pC7PDiS7RrFxl89TMwO2Xogo7cxhiROc+XbuAAz
73/3LQuiq44H7krUakYoQRCbzUKHnn+u0QTDZfa16VYXcHjH3ouGvg4Qly3ya3lo
EmKB3/z8axkd0sPWhUKWBcsErZP22VsZIE3a7ebpAVkAntK+Ahir7xJOQzMxmJI8
Ha5Ic79f/fnG0W8DTMNt/uzrSIYyacfLCE8FaIbxCoFcHDlhGdC/QsxH4BgnbU4y
Nk92vrmyg//5zH1mwa3/FhSj/xf0WTc+5u2iJFAFvN9LZI3lqAp1q0k3a/Ambk8q
jL/aZE7kKZjvDfO8V3pJaA8+rH/vAsPN6UONrkFI+IuLdRUYvnseNVhanC+pzrfX
+OAG4KPg2dOg1R5FUqVGg+K7ZgZ/8KwTdBViR0spONhoyQ5osQ59Yk8Hd455wQTz
31hTIc+v417qnbCgMJns0uRobELiQGeAvUmg9pejScojN3LuQbJ6e2tTZuxNPy6m
6hw6FvAba/B/n7T3cb8PqUBqET3r7bus4hYQUGmjkKl5HbDChNfpj7QBfIQXho8k
FBrM0e23JU0ZOFdS6QwFeHhx+LQc15KraIM2f3vmKbUOGTIg2m6Qk7ag/k1Pj0F+
LuLt8NeAjwAvQQAbUw8uB+7Lmt+hPzOC1ll0WoP5FWDjN0QVS5J60v76zVewVBlt
ZA3ObRR1+9y3XTM/j08g6YtRJ2Eo92UtGD5OYsYxIMDzG5RAuvLthUa1522OiYKf
ovYidvmwewNDaf5taz3LZoMGDjYILa926/LF1Auy3+Smlytp28laUAhoc6HTx5SA
qCGabsgHJng98yixSVGrjUThujQXC0f6P0430wVf0f9b2Dvcg1w2wu2+RGoyVoC9
bEtltETEOn2cwf6ndch9bV0iQwdcBVrnR0sCsmYOi0Nn1bsnGgZu/z+iTZW4rfmg
9FMuMlLTfcskHsEzJvFBS8JYigvMNUtoPQlr9zwHoGhm3VMju8e+ogxQ3y+cdMd5
jr4iuosMffBVg8z1qKaIFhKdUWovpowvhbuGgjAArA/gEfpJVSmzE7nSBcYZed+C
UynhEF1Rwr+eGxZRIkWPeMJnOozC6cLHA3RyHvYBWh96zcsXWheyv1EftiN7+m6x
NA80p+EVID3hVfDHDE0CHxa26W5rpPN6Hv9/iJAreFgE2F8vgx1GZoir2XTKE/dx
1BXn9X2k9ogcQ+VzVy83mXiFYrbHjMTDAQrn1duvxbzHyE6EVHrtopSirssMDprk
sfJx6JScEK6Cp2kkMiQ1A14yRT/7yXXkSUwAang98VnU90TmV4TOLwAP0f37ckaP
Ln72sHnCFTUWmaxJE6Hi4OiEzdg6lvz3MBSCbroRSsTzedV88Imujcw7A9tXdiWc
lcozz8Pqe4AmgIpgCQQ8hxFsJN5rSo4LN8TgoGyrmCBzpPA6XT/mb7UxW0FQ0EHj
TvT8U2AzBVJC8Wil7uk1OQCL44wjlkEst9JkvIt+T2nLa+/g9a3a4OJoe6DPAJeU
voEkJqBhPPF4HgqOKR+Dqz2zIkoag+MjPwL9L1TE/Y9bc3j6680rXMi29wRp5+jt
TIDNRA3BZYowW9uPZF73Ww==
`protect END_PROTECTED
