`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3yuRY5jxGywDE8AG6Vf05/dAlXvJPj9H5i9G9oE8HeGgRTNSQ7jJvinjjEj8pSv
xWM+jIWFUaTvqQwyDnLUTm4PJCLvBdl6t6ZEAiQOexTK+ksjYZCw3UqO3768EdiC
nk3LxsK+wPH/6DarcLTIfUvwDw6hgqT4izfzqtYoqUNm+d64SZuSD3LMxA7yW1dW
KizBRTUB/l6hV4gQTExit8icG2BLJQyBNaaFr1zcEQTawycZLWjHQ1TxlQy+tibl
byb7bnVRE+8xm4ZmcNHSEPoiGsjc3Dtd7WjXaP6WK2INr10enT1OiSpaZwwZDA6s
ZJKWjaSApjbruzwpXMLviBA+DlkZflmxzLgTyw7ha/TomeRiT+h+Kr4HdwNh50vK
I5BLBQn2mZ3hFYWf1407N6G9pbCPPnQy/hKbWrH3u8JUt2B+UMbVoOgNPAQ7QWVd
kNRiXRZyUoY44SzDK0wtVwnaGP+5CkBAmzh0Mg/2fS2gstSpXBF5cip4jk/4ld69
3cygILgtJ72xZtG2IAuJjKAzLfwdfeGccHhhYf9aLV9n4d82ZIBUZfGDsBXbiJM1
dzTw2EnWN7oAcJxKoMh/IYkwgEuicK0n/5/aTqBPR/BE0nejoOF6/kYIvUxVFylM
MH4v6IHvgpiZiKuUtR6w6QK7G4bjAoFxXWktzmpFewhCdREvppLxUMD61bqNR2xb
Sdt7859eWNdaS30EqWv7dgsyYDXY8m62OFe4WYd2bQtNPv65/DueKplLDTFkgrB0
9s3AOCXW7rIJ59Lb2QUUS/kWvmS9tvb6hADhmAgWGR+VaU4DW1Lrhk9E5oRr+pz4
QvaGIv0ODVWVT49y7+h1Ch+brb1mMU99KipvZX9t9HDTzwlsFwCyg+32ccqeQ7Fi
yhtqxYcaZGVUI8DAz40NTVm+LhNoDK4cFvisdpkb0yT5jDekr1LMaTYXO2wvCObI
Ubtq17QDW9u+iuByYfpCOSYIN/C5yOLawf13HFbd7wr5MQfpwUPEmzBzwEdXMObA
6IVk/g60wftHWKPqLq0T1PExXQ3oewf/QpeqyGcltXe8yNAbUyffG9vqq24mYJoB
Dxmp3ROi2irxn9QsgZo+ScJMbKUU2ZfpdDrtdaXhaRVyxFsS/5KpIsds6aIulnR9
p7WY7TcPwg53bS47WDLz6J69y5ALfPn278yCvBLCp5jWP7WHDuDWc15geYO5gRsN
S11oNTYZhwtLwbxBbnN2MWKTlYVYHlqQrtFu5ogtxc7O4PtxI7M0L13iJ+fKmwRz
B5OB7300ZhZ7SlvGrOEMe85I8PdyClYrdXea7q3bsRe+hLEPp9JHYE+20O3Jqypx
oVh+lEx+QzM89edN024lyheNkMbDa2AS2/OX4IP2drVVjIpwWTdxVVD+g8J78B5u
+819q3ZthLiQ2O/g/LCYjFyR/WJgQ6rr0seQ0qvn8t70qFdkNbSK1nnyggJV1ku1
8la/jGxC0ymgL7fBUTKpL0QBM8ehhV89Q66oyCodx18x9Jnj7Y0VLu97htQOpVQo
uoPjcGWQT0/rrQ/AJtlfBBtFatRfGQs+f53sgPW9zH7EXDtGCPK2C8qitwUayICc
spcGqmD1Ls6wZ9KGNznbPauQ6/XHy0fEZg388cFw2cvnNU1Xm1WnW8xPedytQGzE
zs6ZschXTsEfXce90Bxy1gJMhDJvPP2ND1QnwtaAjeL7iFyqcw807uQSxynQkiUK
yEmScPA+AgOG3aqYpt9bgosowbmVK2buMoWNrV1Qe535mQcu/YpxOnulkpif1hvV
AD7+DF3f/2HyN32+TBK/IRdFS+V0yYIhwp9nzLliWQp+C8ggZuq1GPEsjL3zB3q3
ZFnSDfXUNR2C1SKdIqey0CZgl8L+MgGATI2FgEXcNAmba45ROjqspcECI7wQVkV5
s/BHkp5X8S5aRjRehZC4DcD5eI3IgMgd/U6QIsVm3Da0uif1S9GnxLmNi/xKk/EJ
s2RT/IF6TeyN+Pj6QL/Vq+3tqyuUmYYhB4rzrI1Qx9xB0WjcO0/MtnaWaTa99hjz
UXayDIvtLjl/jJSTF/SrulTkL/3Fia+MkF2T+wycYkB3oUlgtKsYfiVYu/gE4TVM
Ft/UY1/wCL5NiD6je+va6OpbgLu7Epnbs2U/14Ym0IvGnqzya1O3XTaxrvnVr+oO
EVa0ND9GpAGpjTjrNTMkUeQVP0Xt1+SIFX7DuU5iO7VTLWvazwyBYrmqwBRrQqQ5
8D63lWSX2DWrG24y7RkwTDUp1AN0CqlCIhTVpZZb8ONJYxmBz2W1VljSl7/Hs/2C
J6qfpj4zjcN5rgNrGKCzVJNK8Jv3xvP5BV3NVNw0cbMSidxMC/jsRDLBXeomJA7q
7R6lxjx5EowkBG5rHS7u/WXmj3dQ1OBWh+00586Le3HgdxSVIXHe2CkoMn23D9nO
2beKxKQd+9J1PYxcypOAhVquC3JUOKqeFfce4fIZZ1GaXTojhheyYKvYGXs4zocY
8e+30ZH0w6v62djNheCLImeQD2FIdXTPjM7zzD3v212WPBt5RAS5uISQ9B6QmxOI
S3qiiiEAxJUSB11OLCApw0Sic2lZNTZFUeElBcac2etQQzFk4VghajqfibN8/NV8
//Q7LBL9az5ZNMJmjXq2nvmcRIKT+xnA9TUtEQc8Lm7wf/sEJwAj0G1JcPAWye8V
s9wdMlSdbSXIUID2YyTinUQbZJVwNH8+lzt3hx5CCpb0SZcJZYIRnmUc2UZ/F4Bu
fQZPA7s2QmMWN1grkf9D6lErYXNvoxGOqHXdsnN3KRhvpBc8WJZRx99SGY9nC4qM
iY+p4jTQ+Lv8OotV3Cx/4/Nd8Tm9fPjjMsDpye9rMflP5c0lSr8ql5ZOPU4u27LZ
kZUPEIBgJNfwHXroa93vFK1DfR8h/tC+nH0JhTpz0Nx1P655TTedrzH+d9dSvRuK
Vb7cAHFMyOPBI+scBEiHZ6caJ7vFM0jmkYVWpmiVT+OdHx2EqmCyql2kzgWuR242
iAQKiFzRGpU8nM7JE0FT5ih/tkh4X7pJieZXzNZw6q7ZdkAk5II4LC9z2FaP7klq
BlYg6ZncTaorbLoUjLt5RciFCg0kdEvyVfx3dAJf86BnCDLqd93iKR/17knyiQAk
IyHq96CZiB9ZqyH3vu0Kx2iNQV8j6KI/3xIuD+5GrS5mo6gu8kX7rVj7p87MHPtR
sXQ93j4JTi7omNpd0jatXJmJ8Kvxy5BbMOAqB9601x4dadmVGRxUk95ugitJ4hzf
OmQUnnZH+Fc+U1OybH/k/CAERS3ST6wsP+yiykdUhIk1Vw0WPWzIBxTsLgO1BY1j
6SHlY68fYag6vImVv+rQRkJqBGpdNoR0XKJy72QutpOSSsLl4LAEJEMkbxCc1j8u
AI5noYTwHRFJ8dB5peajH+n6TpJQIDHUl+S8nFQBK3ull8na/vdOReEgHP+QG0I8
eL+SsHruyrP6kp57iLHBV/hWLS6FLgr6Kopx9hL8YzBcPN9/8gz8Q2+oDu3k9nTD
ozmk1RY/TItxy1n+05B8xKaF/TS6mF3f2DfUq8fK7EjmT2SS3qlk6aIp7G4oKcaD
PNbX/frCCuuU0wI03kFpYKL5MDolZLqcjDi/0EZcKmjpLkGkfSnUD6iGFrBUkDc2
eoOa8/isWq27XZrWDXeUjFMXXxVLa1zyQOvWXsULUNLl+P09qs8KhOmPG1mJHcKx
`protect END_PROTECTED
