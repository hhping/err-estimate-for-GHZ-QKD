`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AcwTjy5dO4FT0Rt5EfjGPwqeqDbSjzS7elmH4o++UfZPyhmdctMbqYtEn4mLXMtc
i25dcnKpMxbCAZXE4BKX5vT2pGSQxWAY3IjfL+8XubS/NAb/bDrMeFwoWQzdPxNy
Mobn+yYbzCcIJQjmLhyaAyuNJwYTKOO5NpnJTTHoytdgCDDa7YtSPX4o5maDMUr0
i9uwlme8G1StpeYSJOc4PT9ryzMAoBrHmAj9tNGswjP/R0vBAkQefXgxckpmiAQf
6JSikf/A4oq1O8jJhNYqMppr2mwb/WJ/YLhXH5o3DWpjv+lU7I6904iCYPXGtp2m
X3UXr+k5nK+GsDRDwUMGpS2Wsvk7BiBpkQHiHUglnWhWPdRR0PI1tcgQKZWBj+v1
NMzQHn1lFMjddUFqkI8Oxbi/GwdcTdfC5khdtFVF63848WpWIEhBd6fGaCXJP1aW
R2QYqQr9mSW7mA8/afCraAQ/d5hWuNVnphMDDDlW1YUkPfVx812z9pWThxe3rZyI
NfVqQinsy7QjS3SjKeE+oJFudlZXhfRqIT9HFJ4fFtyOy396r0f3TWOkACK9dozm
fpIp3FEgw9ySAXzzHZDbVUNbPFRa7j0FRMtu0+cVTg/hehtmAZlGOd93Dfh4EueS
cO5WBHv5a/qyPXBcrW0JD9BJd708vzQJGodGXm1wrX3GLpPMBRsh5sPii1WmZBF/
aaJTd7ZT9N8x4iresvmU7eOcWgyHqTSUeZCdV/NZ9UbdD0IFUs7MY2xZPXw7iGlk
nHGoLhm1h1QHcUgId3aTF1mvyr6TH10SMBIOfrpVM3H1KxD+jB6Jn9zZLkDEp5NQ
wwMGQtMWoDEre6xz+CW/j3LW4b4wiKXDnCj9QubnyjbGHpZuuzyf5oBcTpTSCsf8
KMJgaVdPicBYvlVWTYWcPeik5G6CIWB3iC3rwkMpECPkuKQa3lmtK4I5uYJ4sH1a
oM5JPjMX2PniWuIUksWDAJ7AhgBn73h61d5Dv7EDZN9I3Y7X1qZKBH4alO4Le+z7
`protect END_PROTECTED
