`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wa+RIYI8EQuhfkJT8DgJ6Om0qafLMKDSRVOa+mVO12BaFgLYo8PALAUzRFVfr5Bh
Ugw9FBuyBaP4bC1PNgguKDrKj5vCgLnTUEyA4Ok/bwzuFgofRPnQE1OQc2aYhMII
vhMRE94KdwpjCPVsoRN8sZcsAQa4PAb9pQSYiTtIRpJBhRd5wbAX9oITzgpPNZyq
y5gOCx77E0fFFUFoyM6Bnr8aT0NugroaQZevBI3ZVUwn1yz0jQCWewHYZ/gjpvbd
YuSeq59VdSKjJKF3gUVNPPmdSS6ZXEgsfGUpRsh6cgjdU4xxyOAJLdw8wpAW5cmi
Jsob0raBcCQB+4fY9oAu5w1UGulT63yQlurBFYHeWx1c8KNydNUltgUob01y34dv
tCDKOODym1WCHHXXcJ2zoKUeBwIQAchBGrHLQRhwyfsBlk9behVQDg2ySLAaOioT
X5+HUpHsrTFqHvOwvdF0EgUfcZW8mhDcbT5SsyIa6yeeI9lBZx4W7VDxGq4Hq9Iv
nZZcwtZDi3X8AvddyrU7tKHwPPNF02zTUnxCE6p6hEfi3atZYgZu0IJtPtsaiz9D
MReJW2bBxOc4sq+21to8eEjRPhww6ocV8NqO9FiJmHzvZJhC4esAMp53pVm3/CVr
LOyJVeDsFBmx2waCcWB9JZhN8DRM7O+whblQpuCQUE90IAqVOB9AMEEaodqp8djJ
LP9PgKkvEB2ORyjPFX9eJRCG+2/ZJ7NQPwb2lRMoa0MR5Vfaem7NsOa/DSSDgyVC
TvK+FRWD3QR8+jx8PQW6an+CQaqgPRbOd2bGCX7A17yvDkUoEE59rtpWU0UBlgIS
u2ssTrDFjW0gBNyzHjRQY54CJm4LiBpSH+ysUpzgGZVxVuV7SP5FDbDEv6fT6mmp
zI9dwz/E/iuh0L0qSMoUSvQdGhUGa0gFuvUSMxuqomG3RrutAmNiuTWqIJZVouq7
COw2PsBgyJKebA+u7irNCQx0lbIkB3rS+/MknTu347T4fwvhmS0v2B8vJOrMtHCF
uZxZvb1f08UBneOlkbaSS1W2iXRQaN1buALs1J8bgrLZptWSYnGdJU36I/fPSTMx
zduVAZwVrRlcxJQlLUOuiPqg2nc3wr8IbVC1sIWMG50IQNc+uh7AgoB7OKoD0God
zkmYn9uTj+ZiiDVOlR63Zq40sl4XDlOfQoI4g3ZGOUPsbh0j7wL1fuOi8ofgcnRx
chQ3VijVzbMiIXpJXN36iFlfx7Y0OvQGdspIgbw9FgklSQGiPAceWXPXweAvgRat
X99SDExnGx8JB12StkTvfFpEF5fRj0LQOBNvD1asbvsNlkWJIrhvEHpBTH+O0g0m
XHWnhpIWnbW+MageL1SXjt9stMv9QgzVlWUxdrHhI7FWhcrlIK46gMHqgaNywXOY
d8fBGS2F5QqITIV1+8DRKK/JNRG1eNIJF2mHO1IOLJef5hpOAFUD2UxJdjc45VMT
eqLZxK1GNKwhDwdTPmvcnknonINVJOTD9vjeEBKkusGHkebjC3WzD6pjJJycqhtR
VmzYf2n67VjTJmXy6YgLziZxjq0ex1Ww7ZbhW4wJQlipbRWagvIreVJXgxOwilS3
Ws9af3WWVN2Fzb16xQyFgRL9+1DxfLJX/rnU7uq1rN/9QKJOTNKf/lopT76W5Agy
PS+3BW2w1eFpdkxyM+4/Jjq3oMuZjILTci6YXHtS0FmU1NWXnp0OxtgVBC31QtZD
rgJtcYm99zTL0Xrsk6aQC2S3QEphmTGckfXQ0Itpbeg1y1ZjqrvH+S/JE9GA/jkT
gIU4mr3VUndCKeFr7Fe3KpjImuwUMcysTx9qurbuA6yXU+stvrCtXW1n4qVPuO4I
z0hDk5U8efd2302+p2KB9XSzITSFuVCc2dTb7maf8IkORxIpkvGijgWD+vAdx/P+
+4zOdbaQRP5Wj8qhXBVydWn5WIps9WBMpR8yqHr8pAD4sf3JmB8YQVIH+ltg0lLp
7MoYqv8lgb+9S37crV+el+Pf9Co5fyGthe7RtxYwLU9My/0R48otq++eSRZmyB4f
8mRzO4XeILS63sDm5mh/0s0xORndhIUIspnKqn5faRKJvW0OkANE2Q315c7KBLlH
vdsAdYB4rELNscueNbcSuRRxRZq+EE1az4SW9n8XZD5e8lsF5XoOmDi8SybCBYcI
k9ieD01WYzCwvLxVVO0dDQ==
`protect END_PROTECTED
