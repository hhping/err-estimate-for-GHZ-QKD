`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMqoM6h3ESZH1oL7F54jFcC0rBxor4uRP7sSX9eEkH3ef7566yXF0Y/FOhQPDutl
rmg819if2TdVyA3dEyJt+UhUJja32FYaRBdwBpgW5Wrwo8yjkhx+zE5GMv1rKNFo
l+Xk6WOZJhiLU1k2e9xrt2tlbfZYWqYzJRuW1HxYTbX7+j+AC1vNGzueHLO0pWDL
vnGGzTv7W0MaJvf9MI80cX/ciqtwOudz2nmX5GdRMDWXPZCPGFFttKYJP3xnxhbL
lejYX8aa9jZPmNSOGWk04RjfUYjvhgjEwiGvuNdlD98MB14scgrcm1kGgroKzKBd
T7DAhg5Yo73NmbcSzCSXeOzCpw++tW6cftiB5XWBsPbyrkWXl2N5pcXPdhmEY6Nz
XLglXpdmTdJpV4HbaBEF0WV1XHHeu1sLAjDKCATi/BARy97wziCaVYnXRbQKMi8z
wIBtQpBPux84LpLFjQ8EZ0ocgDVItv9NqRbxblHOnAyEXFtPq/iRwCGY3xUe8Lg9
yTRumLIQx5RPi5SYQS/EFqRk+HYCrwqSaM2i37aCcyh8xWhtO57Ba+L9dJACMPR5
3NqqSFYNA6N51KcZvMdy1aj0UFO6SSFHqvDfBls1S0PEoY7+KMfXNyGvO/cpHmRV
IWU+aiCRWIFPGp3V8UlX/Ib/KwvX6EFSQuaUepxs4PKvEC6KMLOCfL130fdUfXyr
tQwOW7eVWXW9CZsQOdiK84evP/ejeZREiC0mzdMFa3q615hD/UC0MNV+prLl4Ige
i3VQZn/xgD9A0MbCkyIWzsl2OSbN58b2fKTiUx5yXU4ctlmbo3Kz5mzZdb9qtAjR
mPZaMghtp3TMajNrpbVkZI3UDGhBTP1WVLuoag1UuKsS7pzKdWAe6w/eJL/VBDmq
Ear93+k5ufvjspSYWHALf0rdfErkh/ZkMrwR004BjJk0vFsjmVl1HUOx+p/TNhNy
TAs8RtSOCMNDO3YxQkj8X8IBU5XsGE7BiCmZqYX4nCMV/bs82J/fmPvu/JJ3gki+
IYHAfWd6sZ75JPg+TY6HqX7eXcpL5Q8cUYiosa1khWX1PCS+nX1XUmThZzSfgnE0
45pfD0DtDF1GCnQ4KHLYtenk6YraydvqGAEQ8Joqob2uZlyL3/NKXgjUqRNa4go1
Yiu+f/4B9cL65PiXeAHpwzaXVlwNWn0QdyHPiCyfdWizVDgsqQh0G3sJCdC9KXx1
8ayM0Jsf6w4ch52b0XWAkjsTLdxTvda7U2t6W9mJuCzlU7qDIWTscM7UCOrke/Eq
+V1JzrPpasmUO1iGeKJlQT3eQFLilAm9601XiNTfuAcrBbSpmTkNhOXo6xbK9cOc
WOpR20qevLD2xRP5sfX/t1xVbJbHLH2ji2gpMZ1zHWa7Cgim2imgVaCqyBlotGMI
V0YKnLI0Ik7si57hNHzGiJAAinHsrW5FMZ2CVMyfKlIsQ1Km4tUD/jEoJbjnszzM
`protect END_PROTECTED
