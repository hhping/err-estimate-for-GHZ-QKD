`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SyAr/KqX74uUO1FJyb6C7BPmNEAISHvotRTEQwnRGbEsAfZdVRo+jeWjErOtPNbS
V9MoLYcHxBiXUxZLkxcFjVP2sjypcOxMavY/qcSjFSqmOHJ7ZWdQ9CBBd+5Q0oD7
5FU5bRvqCJ9BlrgugJJIDkwMm9p0LuzJr5USm1meSP3v2a1hchG9i1BUX8FrJNYV
3j0y0Tpv8QmBVfkKVmdz31BVuAB436YPyc9FL7F46wWkG171maRa7c7q4ZeC/w/x
bdHpWb/KUq/yhoo4PYq5ctnYZcXol3xVaUggj4RTI77hOX+g/KivR5vGUXi46rxY
0FX3IdPVND0ykIO2PQM7TKuX7Go7enjLuMR04AX35Yfakc8zfokMwgCgUmxP2qRn
5jCoEKBi2Kb3kREjcnysl24r8z1W4Sfx5woWQjdJuXmm0BpY8aHlRVNxHqbtv4rG
wfenHACAcOoZAGe2tQMcQ5i49IjxoXk3gLSl7afijLnfXQX2mLsLOW2KNUNp44Zo
SdJ7Bq8ofDXgX59LajXfDRKcfVP5SdJ/WshdyJE1toRnBahWk4Ivmok5ELrXvuB2
3e234SDfkj5ZZGzeZQtt5TH+a/nf3tB3miLNff3JaPmtOsMeXdLwyqdIW+mzSuSy
YOtAccRJMEmj+HHEW+r4xV5HaB9bIDW/RACiBr/XJXuzEEF7pMqJrOe704Itp5t4
0i1gfl/KwzDWnxkW1cZVAXk6EDeQZESkK+PHkAO2j8PdbuB9gPYvA1tRe4J5mSKt
EHmhUWTWtfzwKM7sgRZ6gAsyx63hfCgcLhwpyhdtzlBQX7UXdOdRQrHZ1RYupHFd
`protect END_PROTECTED
