`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSYAj3UullBNPxts6XvN7nFvHEbO7NTLi6kOFzD/M2lUm+Mo+nGkoiXlw6KGbz9M
J9Nf6wtjxvQ3XKkuw/rxAWsGMdzxxRytHPbQ9p9A9aHDAHXaXCY65HfBwM9KbM9m
5l8lx5yKTL9tVinvEpDa4QsvHWaxLG21Zf2d4a+YIV2fBVDrLrVtxsWLzSG7AI/I
+QpY8QjSzSN+SBZvYOMdh1WVdE3g9Jo2icft9tpyFtydC8HtagKzl6CVFtfgwWxw
SMAEJb4j6CJRFQazXLd66cfnK1Z+SiLXM2aiVH7SLJ3fSBXbbJtu6nC8qyT/1GQA
TakseiGNJgTNjKITh6i5MWOVic0sakFMSfveyhYBq6h8tZF1sCUWupJNQZa/fEQJ
PUo4aR2ofBU9/r59dH/nRzqeB0JRp4IMlqUqMOoSql3AXwiva83RmxE0Z3Dh7M9S
QLZfW+HkQfBtEn/bIoyLUn81VoQRL4o01mCoESR8UEZfJcx9F07Oh58oqMM1FR7o
yHHF+e1ot6n3TpCGzcEDRWHjxYtgKu0qO/vkihbkKvAsBp3B4yXjsUTUo9pp9udG
sE/oyIk+92G/y/JC0PPyJCyYWuDg5K8Z4FN2TfuBF59PSXVgjjxd8sBzyKBt3/bg
lX7acgwRfMf4skQT/A1R9f8xBXecE5PAZJFlvVtl4b/7PokeEBxOZeoPGCniCg+e
OhkN4lTCbxRS8LHiEjRRUOheeohAS1uTjxQC7RCXQ1x59A2ibluPQ2+OpT4NiT0Q
MPRGMsdYzSRjquH+e6TA9H3sDLVcrauJv5Z66IWw4ihlCMMY36hWhfQy5DdzkUgF
6qu/Q3s8RXuTWQ3ph923eSIqccPk00SMDXfFtz4+8McNln5iavo8Ad8AVvK3rIis
noA2O9VYB8vOwvhQ6aSVgtzHTofUdzjTWj8KgLCtiv2oqhXkEkrUldceMy0nHjps
QiBniNKPtCWijwEzJiyPDCMaPzhlEciIPcUJAziBI8xOmOIJFyLLF/rEOlFkgam6
oLCmsJRzEIJxK4q4E8zNHw==
`protect END_PROTECTED
