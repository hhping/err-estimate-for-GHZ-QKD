`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4seiVHzH+zofjHP9CqUnkQNkiUlVkwy6TOkaH8rs1Iy5NQwP9rRiqrZc50KKzB7L
FatEpibN47DjgEz9TgTFhyX1HST1Y++dWvdPwXmit+SLICyNTnw4eeMH13OVmQ4h
AjXu8g/i5aeXjW1yIEfeXdeDklvPpaqWKYVGfek0uue4pzOZc6QyUcNMJ4hD11a1
RhvU/Ws8UmAdMc5UAlsIPhM2eqc+4rMre8nebKSeJ7LtbZ6BdFBIHlF4YTBkvgPa
A8FGyQsBsy4q8fvdB1rl+s6mpUoi4fZ71ElOF1Efl3Tv9xu14iXo2KvKoDG2OTiU
Wsoh29yluQ5xtyFxB+Gfevlp0Y8l66QlsL925kgRSyg2G7b5yp4l7wVNNqYSoiM2
BB/IS+JRvyFxcjMAORANX8Iupvm5xJ8icHftl49CWdlSsiJlmDKLIXjYqSmkSk5w
Kr11Il2m3BQHEl3LniQdJaSSYxTvpXXx9K7rBTQpeIm5OwnrbmuRo4Whq6wotAIj
DPMM736wZQc0r/X2MReg3Ou0nK0tMqPq/gi72g4B0pfxWu0GAHNEZnTnh6BMiEHQ
MABdnQicmzcMao6Qj1+SusR4YtZDRaAQHioQMVDo/KYuas1/Nx+Ax/BGcQWkGrRY
1lUU8KgFq1D18FR9dg3zHSckdB9C30tL0TtSYperGNOLAKoS4iAxrzZO02/fiwh1
igdXvKxhlVZSKxYJgfOx28u4pdmRZD8Q1KgC760tOWRnQFcrRlF6EZKsJSRbut1c
bVkrrQiNlUnxTgrc1/gY8JpZ+8ktTsZD/IYzIEJXq2VZgVKxgD4qlZPjRVNzzb8q
1TubuDzqPmQvB2RVttPKtftr3esWTh/89hDGe6sHlrLlernspkHxNBkAxvO7BHad
TxjmRRV3y2Ijh2eWhU84pSbz+PuBZCpAv+DYJKQKPg4xY39/aBCCYQHvM1yW9R87
QrwM+uHW4t+z0T4bF81DNIELglSJDmF/+7KAgZEVOr2tQXTEIHBJL6LSo5NEiKMA
`protect END_PROTECTED
