`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaID2HKpIK9Rqwk+F2qESOJnzmo3lbsp2UQUm1460GqzgLUWkysGw1RpPryu4eOC
FZYXzmDP5XAmhAsTMG8qkWMD+e8N6A2xxHa3Nqj0iADyeRdERc7JPQWKCxChFIgs
h4qLhU+7ahZGydZd6k8dW2Akda+s24SaCt9/A1ki9U6fzi1pGd4yOT2y2XSoTwdR
0ijnvYel+2AC7oeGvuZ+TYT6ZOR7Wm0y8ZXGN/rCWYHDAA07zg5jhodnJTpFZUJE
c6pkbFKuBw0fC7rwEasvAQ86j0+PYYnQiktTgTrG68WFzF83IckcdPe70Q6+28bk
DVQ4bVySg3TwCkiJx34YWdL2lZHsYtcDZrfR2W2XIQAboJjpAjv3SMzISL6xMp4Z
cxpfvhtwJJQaw7xRcqY5D9nLEHfXcrpb9lqbZgVoQug8S5k9e+8qyT7zw9kGlaf5
Ca+yU6+CM5RIvN4LER3h4qyQI+k9HbjGCR0v56QvCO8QVQceuVFlYtgYWF1NmWbz
Ad4fG80aMmnUZGZbbYvonprKC2en4tkTu08dXiqNsIHyRRCmZirD7C/8bv6as8Mh
n158kuoYoFv8pFLikPJpkuC56/cFVEWWIAJOZ31gvYGE5h5igmFJHMhoPMS214hb
t6hKfU9MJv0pwJ7t8xcRf9bdGqq8CYjUw7cc4EaFwlSBk5WrqmFmjICMPyLtVhxC
ys03FShRULHcSaGwRYkCo9nVulRNeT22qKsd/tImZEO4POW1UPXwKtCK83rxTbo8
rFOU958iit3o8QIWkjjoynM446dKwFYmQsp7r/mfRqRhpF8LXXZD7/YyAhZY3iBW
wjz7X021sbf4IdY7xjHzJVejJF3E5h7FA6O0dMJzdcE3x6Azoczp7p85MwFxLa88
Rob6FQqc+hw0AH496kdD+mZJ6x+hZ2pHRfiCNtzyQHpYrQ/BNtNAxTME4PqagiHs
Nzm/h91S1sqT0ZSr64hmldL3iCopQuQTiaseRASyv30SvJ5EQHb1M8h0csYuta1c
hBsacIiltNXr4yyu84kNAvYjn7pWvlB6vBrLx0sc/rNSAmEJD7MiasDet1xN55Rk
npiTtY6jzoeyB82EMPaTvv5i5wd50h/XHabmgO+9XFOvVqRPt0xX8NblxFioEEw3
CVwWru0udDTePnns1gzhXBCnJ0TNIeFtH18MtH8v/IFumbKLIYHH/cNhTDgDvnna
CogT1EujVDPGC5PgDOqxB/GxWoq1JprTsLzV/4oiBA7lE2jv1Rbm/z4/WTABmg+b
5yFXlkod/+nLUiZhL/OQsi7iUZKMMzGK6mh9/neM3tyWygBjXZKeEyLijUMwlj9J
pRxsaPnR2UKylUbm7/YC7mCa1p38CJvsl91YlQm8U7lJntMn5h+VoCQH6VB3RQyC
tM8uAHRF0AzCR+3l8MBqDu75Rnv2A0T9PufuvuIo8KlHyPc3Esy4Zq5RG12AiW/H
F2cDVfxnu3xNfExZFix2/Yzcb0IL/yEwn6VSv0opUUDC0O68PWFJ3HdG2EC878Ak
h1e5GlEINdikUw/Ln78PnDkvBJPC6mBMZyWSbJTjUGy9PwmG7bn/+dHtxV0nT1zc
ZG3rGkE+lOOYtutMqLbEqPCu7dT8E0xKU0cl8eS7wxipcO+wh4rhfnkG0hEMcb7q
KnRPryUrz2U2A4dbZgLB9zycUqKpq7nfKh6KMsSaaZAAMH4Qyzc5s44I0yb60pw9
JcfU5ME/hXj6AasV6Mk5GDylfpw9T7o4oYtttBpuienWAjl2OWb4tu0uNWdcz8L8
gUSYCr0zwHMs8xm2hQDP4yAMF/SYmpbJu3Yd482tBRyMpZcjAftfRWtmQDwdrFOO
6YAKFk2A6SF5PXTjNeBPnoy1icLMIXKFmCOrz9hiSAd4EqHwMyZ0PswfLikKi8A8
tV5LhKRvKwY1nKY+CFWtxL1FT/70+SNXoLg9H86SxzZCCe3jmm2j/l4zoFKznHmT
XTKQz2KpaXGrzmOfYo0+OqpxO3ECMpqS78pvUL3DwHYsodS/YkOdM3lSjwI/xzma
UcODFI8LG7jWAQcuCBcvRVQcSV28b3CLi2Q4bJCc9XJI3RFg1G/areLoxQogY9Ry
5DxnZQhLSqvOHP6P0fg0ueLcVEOSqAZQr+OKo+EyIqcYQWRd9+vEq3lV2/Syzhgw
xQTYRaRi2Z13jlv92LvxKEpizhunBqPMnJ7mxQN6gZvz6zsUJgNvUFXJztetOTHB
YAfDhGicfOH+qFQiZgeYs8h+88bSj/5hEMWbRjHt5wq5g0RdjrUhVrDrTtCA7bF3
`protect END_PROTECTED
