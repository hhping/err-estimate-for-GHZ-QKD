`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WH+lz+6J7uO0lAT8pfe4dNli1tNNvGRuXQshwZe7FAGQC4cRDap6/2dEq+tNITDW
WbcWDRh+Fq/LfZvyXplF82Gl6mqu2C8QRmBrGcPJ5vPR1raSqbw98YSKWHuTumnQ
DcFJzQ0BQ0V+DwTVzo4gktFAmMpLEfjKxe9yKyrTtqXVXIsnyIqvMtfkSW8RdY53
Mvi3Wrpw6D2eX1aNTQrG9w30q9cW+gEbYR3C9MWPqkX1+SpMrWVQJwt6VcEYkU6Y
cjjUeg/+KkwpSWC8FSrgL+1fZwo90WDxf5zyplUh60kVx7FoGsRDOCfApKCD3PBY
ADIpHzHTXQSqZQgZ1/f25QUrTrDIQ/qi6jjp24c4czSYrdZx/gh3yxufYn8m+DLZ
Dsk4UOWYXMz3FyusxaqFkoAqTSzG6q81RhMKp5KLpNWMyNYsORzODF98ZESzixvx
ZCj4/1kIdtUtltd0npLqRQLNEhX3CDPTbaUqhu1lPfHEa6keWvEVhT6rEUHPn5CY
tIZRx3MOMrr8FuuuiXNRWOg1atW3y3qP430N2KsxkAJBU8zdxFQJwdM91E9/S8hM
ZIn0EitCG/AANOCSKXWx4p2ehzMrW4oECL+Co5pdq4geueqy93puFXESArdZJnt5
kP/Bkm+zzXM3NjDXfdCStVtJ7cWUj+kKlBFlyrcDzkZYuYYkJNGeYIuxZ97cwxzC
bLqJO3CyuzqlNMd+V4L+FWtn9j3Sg82vUgPynRxvRepa8eeHYyAwloyAVGLupn1R
i2O+T2EyzgJVv5sOxgghWGchi/yoeuYAKdjyQh3IIIjzKW8vU5NVYj2PMLg0iaTV
eU0wZ/QMe8v18tnyZpPTudB0hocy1enNFJ9cbSwj4nLrE5G5r3K1Gfrcj/mzyB1n
hMOIBp0I8Vb0dSa5I5/YalEMaNykEH+3vseC5eSIrHBthFdvUwgfnThGzN8x+JX6
K9AkmJtZc+969DAx4O985Kpm0/4r5aDtB8Zb42RXl+1clTnoAk31z0mT0xkZ3k4U
8TeC9ufIR88GSSwJhJMv/drqqIOOko2hx5+lAZ6qaWdZ+ps/DPVC1NXQ4Hpg6Ki9
tYjVXDKB0evUi2CIoYL7gfnYB/0u6cqLKmVe+wDEBIYMPwQzFC3fhb6voPo4Lj7o
fgy6+g4gwBHL853TVqKXBPyDRGEQRpL4EBf2b7q9WfFv0NF0zE2uvI85pmKsjl/2
BKfFcueD+b4CUS5jBWLgnVJ4oSSBnOFtcT8e0VJka1HZFrxWFlaWADgBxhN12jdv
FKjxpvUqE6m9zWY9ox/CH3GmXY93xfjsDyBfWf3lPNwGhgimvFm3D++Ai1m0ngMu
XGAgndcoxRUOkYmfuQN63Paiol8oOeySPi53AtEth+c0DwkYHzzGVmVVyFfwGYZc
NQYF+94e1Fj6CqlRvii2CnXkPKqGPrdyCeRuaL8Ro1nVGtBZr8pbPq9OtrAZETy5
Df2mkxyJsOmtp69JPcqctSVOUrAqWdfCau33lb/iIZo/wonl5FkpaYLEtGR79nT4
5d+h7mfGlUWTB1zFEXEwBcijCPlWVEsC8QQNDykK9mYy9oWKjzN3pj67N6VhskFH
Uo1QMfTUvY9RDr4rzPr2QOzg7ImoY8r1mOOWifpW+sD3DgdSMpViibwM2608yl3G
SYBCysrTuhGET0WYaoN3vNDekOlgSpvs6SkCgsMYND7BlCx2ca6iPLUzs5p4p+2x
QKZ+O9gkxVMskNs4Miw3cQqa4D1yaRogDfD9dzcRYOO+hOdViNvk3Jw/3ICixgxA
`protect END_PROTECTED
