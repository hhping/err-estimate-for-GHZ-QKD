`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvvhxd+SU0IM6Rg8CxDEDud6U6RYsJYiEI9l1LIFyTtm7qpMaaTe9RBgEzOpi607
VSu/7m6N4wVWbd0Oo/565BDHr9A+sXMCeWl5GDuL5BwUV3Uy8lv+0wqUE/iU7XTT
U04tOD6Okkvbb7zXXIipSNDpK5iljrfqkaqAq5K+HlwwDitB8zLPBTO1cBX7MY0L
2KzNWfe0jDi6TbLhHaiGe/BSKtEv+NjX6ZKCp83qpWaBUuFt/KR3zqlx6bieJWsb
udzlJAZIHRSaVNgjCsV/JmUGN0o6Vm63F4SeBK4g8pgeZe2JtLTgEdsPHuED856i
dMQQXcPX48z6h1Cyuwkaudvvst+WDy3FzAEeXSqzQaoTJcreXxLnkbQe3GsDEa8G
W+LNaeGv3xIG2Vm+wlg5r6gIosO2cpi87WvoeqzKRWFI63EUM1KR9Iauptin3rkZ
ZWUiILjl27om5Q+nwdMFUG5up4aingetTY6yEMlwFdB97NVBn0b+tArNO9Z8oTUt
ilkvQ0GQgndu46nRSY9Qc/pMzTXv7tF6k0QMLn3EC/0eHNjm+JQSbcZ1wPLw86xY
bnKF75pfm4uPOtLgrWE+6L9VSMrbwBMMF/rw+pM/eyQBeNoBMHdsfBYA3v3tris3
lBdgXlWw33yCgUPp0sgQXP+3HDLNke5glZZim1moghfPAGBCx+48jga1PeTeROL7
/HKK66x4K8LI1LS6B9ddWCYZadQngO/wTpKEarInukSNTbDTbas6n5pu1aIGm5OB
NAC5iBxOl5XSeRB+uzlmsMDRmtbCrWBUksFhlDIU/KoTMTvJTmR9uMmpFjsFm/nU
25SWbLhpLLg4E01frrbZvXPuBwkrL3B4yblnl68ILHooP33yLWST9Ar73Nogocvz
TrOt12RiLp+XPQb4cZ7P2A9nkOrzLIg6tide4dM2AT1mKUn7lzAvmkkeZ1yNJK8i
Z7AQW3xSTXAzYAxZD1cCsKzdRQLXQvkHZ4yslX2lIIS+yFGgh1CVvNRybJqFkhYX
v+ar0yTKpYusmD2mFgSeUvKpFZ83ZOAaZdaDj3619n4r9kcMEqOFaJUEeyoLPm7M
kZIkRm1aXdTxfTquhlWS4Y2QS6TiGjjU67xwiQrnAvzmsEt+lWVwEOz7vjdOVj2S
cittbS2TQMVG08J9wA1z4LpBX6fbjoiMOAodxspbTDnMHs2IngSrEkr6OT3jyyNx
qkIjCME+mFsmXsLCQz517FVSrIoG+FwCMu9bxfLozXYvh0GGwi+wGjyjYenKoQtj
GiPi2Ea+NgtZRcEdn9Cl8vwuwmiZ2lgWAB+9dQzapjoeNpOlABBlCHMLej7VixuY
MYEhBb7y87XNc6UPoXZlONPTH3FI6P0SwNeEScwVK3PK12Ygighc7OjCo4dXubTH
DxshXbCdab2sVWzqMs8Cr406NInpRVHaFrfAQ5F5dBTz2jZ6/41bAe8vQaXnqOJe
fx1qnZACNiILiTC6hCosU7cnIz7uXXbmFnoqivkn68LrHJOhwQc2SHst4WTEIo0t
ZuoaWqAja9ciSBrOjuJIcOXxYFLDoXhITbfEGFxmeg22j2e6WOkXCKYB2+oMvpHW
N/PgPMNT5C9AXhsOKPmtdtZpExriaccbrfxb/2R3jEo+YMCyXt19tO4oiILkbndz
hr8C5sDntVb6AfQcGdonh59iBRGYJkiWOZ+bpgDzbjjLlAM5wm6YSRoB2rmlfUCy
tomOYNZUZbv9d6CDX+XOlyGEoITguVei8YIpsByYe5D4vZ/de+tp8IL3aG/r6wOf
PgV2vZTES1CmEOR+nrIpGw==
`protect END_PROTECTED
