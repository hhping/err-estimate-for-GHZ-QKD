`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QS3Q0t3FbnsNehaTXNPxo4GHJpLq3Do0Fl3baL3e1k+In3dxNK3a7/SOKpeyCPym
3ATWIMJPb+YIjPg1qBMFmg9vau4jktnnyCZAUvBENs+s/eWFukMD3EIpoDnnsgFi
tiGQQcBeHnQfENSPQX8n9Z4qBOocuLf6LV5jVfp+M5bDUbVP6Rdzy/nTT8+D8dUS
QtuLXC6tQz6XEkJus7cExOMMPqJAk/cBXnLMVWMXp1z6Pcy1YnZbUaZYWm85cEy1
2CXbiqcLS3TN8JitTm8ME2JfY/Z3GZbqk9LWJRtRom9YLeN/h+tWyuRyfiEb0OFf
14Hnv/AvNEm71Dvqqh5QMrt3dbK1sPotJxHiBFt01o/8l7HKiFGHfcbNhF9TnghU
iH/KHpgl9bHF5/16SaD9Faj11foM0fH4vhUrtjflkYw=
`protect END_PROTECTED
