`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZF5uqsOgJFF+6yOAcwOcNeRsP9xzAs9zyYrncBFgatDe8KNX/qK4iGg5Bi7vZ9u
uxdMlNJFLHxKGJxp5pJxIIiRj1nOyRFeB4kC6n48oDMM3WKDF/+XOaa/Aah4dAIW
zJZGbcfxshBTjstciIzBhStjjY++UG/8wx1iV1FtRTd7z3FFDocqx31Q8Gim14Bs
T2x90X0Jf6HtcWDgDS9OgRU6EOdWmNQOgYW0VXIScf0fadOppNXHe4bnW9jbcd/X
8HVeT+wzBneUXXAib3dDZ6rg/FvgRSP2iwPZaAACtskaK63xdBpto2AXxF7IVq+C
ti6T9+OxM03IKZh5zEdY46lw0kSI7z8mjR+OkGPQDuDkFdCWALi7z+FQQWD1E3do
J+tsdf5KbqhtvdVVABPkeXDpbTW5XBv+8KidbVa6hRd+lSdQsQy5DpcelTuR88EQ
3s8yDhqmGa0hA+IAFLdfC8aoP5Gvhw0XU0LwypG7G9zYH3e/70ooZNZUJE1s8XKc
miXDbfxYlZGlgCamrFSJmlMB7fVsU/l9AfILp3EFXMukjdTwzjJdl+dHpKMX5e28
tEhcNboASGYQ80In1OQQI9YDpSaYcfKfIg7yZX9SfxslIjQADpKtIMPH+EajpD5g
ISyIbmnt7SiEJtWck1GoUePiA3HC1Ju1EHB3nuGs/H8oAbJcoHl3CbPpUqOFhGBO
JZ+t6jd6F+rMVkMYG76OVr/SU6Cb0A0AnkyEHDl1X1YKI+0bE2q4SI4gUIzUIneJ
YRdlTrE9vhr7kW9mqxCU0fhDarb61oNym9bP8jB0qp1G1m4CApm2m5prhxJ28lOL
6uyHKxvy38+MjYWTAm1C5Sp45YeNHmRxFflakFLtZZYlzqIR1H5yddgVqLoKjQUS
B/qCD11i1lIF1YDRwxWNiHwy7AVuAmJ4Qi8aEiTYNCu8BT4qXkQ5kLfbrK4UJs6a
2eVnaaqgW9OtuBdB8amQophIQEqMAJYrloFvWcC2z9Q3z3xCnE3JP9NCxKf0ev4X
y2J9t9lCHesEUcht5CNm61Q+Y5vmdi8iyo6vf0oU1CqhqUNXBKfreruhZqkvay6T
aj08DgFsAPDlWj4rxN4bSHbosn3qAtuk/6AXIeNubFk=
`protect END_PROTECTED
