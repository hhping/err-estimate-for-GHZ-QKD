`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dD9SB5OloWYiblcFLje5TIjpB9Xj8Z0sm5x7cCDXnNwtabhomWnGlx3C/R9T5xnL
lXubqGYuev6y4XWh4ON1DruNyjfqUvX1UD3MVWMKBW4HtTCPKnHVCYy/L6FYX0E1
HBTb7asxvlgCGIsfALk6dt6n6f6A04FsJIFjYpp7dyZNwvUBSiRynW2zyZIuG4Jw
N1/t3WmQdkFOiIjRTBmfh3M/6Vs7Y+HdNMHm/ObUUgknwKfFY+4wkMXhQwT7NXRH
XpgAKOv5BfXaNRFmeiirDc8NIeIqvsbYQg10l4JgzAHCo2bU5nGlhymHSUMIV9Do
lOWKfBQuuCf6fb8W63V/QRuALgU2enCVgMzcFnqEinJy08PeBwBteIVzl5BRc16q
Ym1td8pIbj7b8RNgXLb0J7UBSlOA7pjVkE2VvwFxcjrxNHIo5pDyj57Zd6CCsjDT
im7ra7F9cX8YHnZQW+ba0u/DAcZmZsvthxg2KG+Yv/xpR6JTYpr3Akf3HR+xDLs/
7+SgPRx8kQGAFsroUxqMiLrPBgFckPr01pvBErSzFRbYlr+3l8Hj/k5lWTOjqpsg
6AKeGf4qmtuiQtoxwxyl9MzQ5aG5dXZtjfGO5WhnQ0aAEEMDxwbMx8S6+3sLU5aD
J8u4flS0SLpayUXyRZ8OmUwuX9FdgpODCvHT+PIOII8+pdSikChj7rQfa3sWRGsZ
hOnbYZBiQZ9dZ4Evc6Y9JVvZQZYvpsaM9bMKuUILAyMMMeB17m8wTC1yyDKz5S9B
PHwqe9B6YTSAHe09zEe2qMi+mOXNYxXvKNftzrdkWDhJg729sKqFRwUqXhEVPlwu
M3Ljgmv8W3tJCFcGKqe6raFW4UOQrHD8GUxLWGbUd72NnnIYvyTwkmYTq5b/OQRq
aISOzF5qpnqS49YgLMe5yk3ALpdB6FjdOXqkbc/YwMhZStDL5ATmtYd1/YMKvnfm
olGjUbdDWgFDnEbDhRPt7px6/VBA4GO7vf+0qYjsX1WGr3Zr1/kLHQIOtN3iQsp4
n+1x6EP8DJrPG3RkFovNghvVXV8vT4rVntyiaGZHRwqWJmY23BhJjEWFZTUgjHvR
uqZpcIkx6hWgasPZMuhvew==
`protect END_PROTECTED
