`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqghvK74FOOyuY4b6ameg81Y/BT2OYm+hW3OXHUEtQg4N3bu3QFhhdUDCYoOhZBd
+zfwUygjyA7FbHip9tpebzW575h3muXPXG/VpPgWtQUNnYJSvSjnhVptctbKJ4ax
6FrSQ75v9ARSaxBNig84RWTxQMOFejYZ1VfC2Vp9zfJ1NvBvO6NhkAAuSU2o58ww
blGlDxvO8ZHgOxwBvWQpqWseKtmuj+cp8PE9VT6ZIiDx0gG3KWc4dhdSmY7xuXaO
/gIkA8NuCuStw975qoS9ErVFUtcYPMnY7Xyvc/9CgjsMw0S/jEEyMKXuj0PC3ZOA
enGPqPFzHeOVD3+1nNVBIF/aXyw5Vk1Yoqm+uDkzbA7GRp/rwgtasW0WCI4hjwD9
PNZ49Ksj/3NzjJ50rOHXZNe+iwg8e1AR3/DEdgTPaGoWmPfr8MPgPrTVh0xaagfg
yqFPD+H0sDABy1RtuIcNcx78WwCGbyAa+KSy4otDrlIVYZhtOYKBiydgCPzYmzvF
tg1gVkYRrHkVyK8luRvXqRv3Mh0mzjqnhnzPt6OaHWWltCQvubDZV83YkZfSGcPP
Zt9MwNRJrUQRwuse5aSzeVg2tUdv4BcRl23pVpwGM8dLBRszO0+L3ocgLod+qzif
R/RbFNkQSAN3lwqJQwKL2rNSvsZ0wFgt7kxMS25dxBnz0jvlxAKUHM2Jyj2N8pgR
H7YRjr5GiE+srJJwROU71shIAq8NP66J/M/zOTpaY+smCVITUKGB0P3m+KIxB+Qg
RtxPYTcWpSZfRQRExcJ+biI77S050ipZNX+Q53ATk+u37yicI3AzLKTzhEHg2Czu
rroZ3G75X74Gt/4JOmu6duw/OjojkKNp4HhrS83d26Bg7kB3EvLrX2OBTIsXBHgU
m9t4v9sf0rXhdJj6WZ0QJ3sE9Pne/3OwviIfyK5yMe9Aj/GopVuCGpykL9ESNg+s
w1ssV942+foCl5z0vzreIzjXyBWofwoY21F2KeDWe+tL0gYYo++Ly6Cy0MCmZCcK
bdbBEkldCelKHwipwJd/vGz3JcmvB4OCbd3kfDRxoiqZ8/VxOr5to49p7y65duz/
yDFMqigCvC9zlRIwsvEfyqI6ZWIfo/kYWa249Kt6nKuZHSwxNRmSVPBhgKBp4jDL
z5zmYe8JgqKOf+PxTvRhDf1ec+6EEqqmTwPuqB/3dsaN1++HWw98ZWO3+5cTbsPA
fcp9L5ezEW72+ixF8O921cO5LF4r99LxkzKc/DU4SlcZe5Hfg4YfSTAFb+bNCyQS
siCamsBhtYA6MMPcJcbSWtBLNNz+Sk30z1XfG1sr2zOE42ZR21fTdSLatvNtaynr
xHtD6W8ryTW20guK38d165vUPya96IwONu3Pw2gg6Nx5vAPpmH5mDdF6uzYimc3z
Wt7xt0KqimysYUWguDF5WNPhb+tlgXnevFAcYfpaqkR+AixlrTYAv0Ce9TvD9Bd/
nbjjwcUy/TGuwrupy6kjNdTDLrWgF4XwWWC6vIg40N8GRzEowyKSrRk35AsdC+y1
cAkf1iGaE02E8FWxqYf1dzbxfSxTHFifkTd+E/qQMwLblVGdWzlJjelPJ9c0I5fT
s6RWnO+Hj/8lIHgzs6EWFl9VuYUOzQ8iI7beGHWxneEFsNlHdvQL0ZRtqV1MKwJK
pOryVg6eQ4exmRHCWJcceL/5/kkc/G5E/qTL2zQp1/JRoDRrqs8UKghTlnJBVVj5
TIr//Lz0mkZ4lDQT74QSA2VjEcBmfoSGd0yEbLpgGhUnxVmhAUXfu7m0oqVUwiNJ
VRlQCKNxxvCo264w3+mUu3lrL6/3i9GocuoyvA7B6+yQJyC4UPzOrQyS+wVr98oa
hAOiMexKbnY2do9VVvllqUg9P5EjBq7Jhy/6QPTtrbpkV+yN0+N9x0s/eWzSrQ7E
wVJumqnQbJe4moANSSkHt+epvgWEtq/9opXJEjYvsbnqEB+hxFTebqWO4+LUSpxs
mCR1I9ryfd3SmuLQKjI/qU4rUCfOHkTY4GwcbqPgPk4kOYelCO75iATCi5d+4QTh
qSDTTrtSBYkUjXEfuf3oN59f4sjdh5/CsX1KrFqB085T6hWg7u5joILTWCeXndIG
/FqyxmDNcvzHUbsBbkA5KkDDKI040yx2q7ccWLfIIM/+QFN8vGIQGKjz0p6U5Eyd
3lLS+6Lca4EPsIFpS5UbaKLCTmAXwD7Q9V2pofUY/6OMn2FlI34N2fl2gJP+N4b4
S1gTXaNAdQgw7DuU/FC7wfDhW53pXG3T/ED7ClY+L1cxzNRDjOKhwVdQ7OaApUp1
iZcJXCAYyTcsPqLHq7YGKnMGIQsmYyoFlSHqWAsOsAvE74BB3VmORvzXntYkPBwu
jL2cgXkRkt3RzUaDJXw0DZgwlZEdwenawi92Kk4HDWETAMGMqVx6+Fk/3Qnf74OH
Q92GVQJBMct2DdOgMHLNF2gpB0zP9zjxVt9+/YX6e5E=
`protect END_PROTECTED
