`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tITBEZcme+v2fS1tN9RSGlm1d9Qn2FIvCDV8guBA+zuCHP2ZBsH2hEn+9/1L8uHp
yIWR2Fh3brBbEpf+ivgm7JbzTSwjd4TNa3kyUknX8kj4H71Nr6qvYJKzPJBjM2eP
eju35EmhpDu0iA0tQlNhy3Z5rHxOVaXsnFmmoufQ6FcooZMyQjsF6B0u0mqYmjdd
UqkyYJm0VbwXw1oJFMbcDN1DUbe0z06cAyK3Ma3DJ1+apcFYUs18WEuCIzXuv9gn
v9mtFlWJvxhjxC84NLE4o5hLFMxXK3Vp8yN+KzRKcT7y4J/GBbFgTviBfNpT+1PO
KFhi0/4ZvhI54JTJ/xAnPQCOrkq1+QLApL8NmXMgYB4cSAf2OLNQlESmOMjcoxok
QXlZmDD1+n74+2Do0HFcQRg5u4x5tMzlsC9ih3lsmtvASt96YEKWMCZ713uF00Cz
BMoR4cGuHor2bBtZODUnmYV9nZAErrq9NUbdF5OHtSGVrKLgng+6S750LE8pv2+b
NsX7mA/zAnwqTjOyP23Mk8cIvgX2vcvXoXkVyD21ru6jdcJ2uJu01XZiI/1D5o2l
oGYwP6ByNv0/f/nKASbK/63jsC1+lQp9bVxa6wEZMoDRhXNGwW3K1NClaV2tMooA
VJa5mpM5JwnfW0sVzmuRDvTaM0H/OY+YUfP9AcrRPRzPA2wHXmUrlUsCB7D3wwjW
QfQXDB7Ga0X0bea0dsv6IyLmFLf67kcDJMLe4NWb+kF2fbNmBE9me4RswM9hgh91
0f5MQj3kpJ3MtY655mJ97cPKMQIZdwxzLgnU+HWes31eGpmsFuuscMXzoPtWuObd
t4sF34qkpRzt4gXsaa0Ql8s1MrwS7AU31QuZgg00EnjqMA9ZyJCiz1XO77Zmz4JR
IjLvyAzMPB5DcrqE5aRuLN81BWOX7EKxWuy0EW+RPvM6g0+na0QM0tuX02CNONhw
2TtZaW7Gl3ccLnJN1p7GhxAfL8gIaSNSjv0YlkLVqfbbWh98r7taRDZTDyCN9X6j
NdxWlQrQXUKFz0c/TDwLvQ==
`protect END_PROTECTED
