`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJez3Strvbjuz+GiqSdNrbIFNeGBRsXiWpLb27SSpm+qvsZ5Fqb8VB2DN8cQIzN3
lwQ/2287IXYugQ4c6RZI74MKh/yzi2/A0eBTE1ihIykHqJE7iOcAZvyT1xREAOX6
JSoji54Qa4j06nG0syv6ySYqde4HGBbXe/+5NtZj3+giVa8KXujK5H30iAG28ZHo
RTKgSkNeZD2IeIya3u4sgH5kZlamrrxmJi1WoXgFlukSAiRBmZcjlxrLLfWGMrCu
RdtbLkv5lp5vSgV6MnFWtq+2WpWEwa+P/UhKP6y+bduBf+w90x0/lR1bFBZCcTcb
uNxZBDd6X2/tDNGcUQ8m5GiQN3fDdwcbcDZSVBn1QNqd0qPE7QvvsCw7QCx9MJZ6
G08UbUAoc5g1ffxxAab4UrgDE2Dc3LwntyKebXHgZp/DzR+I953YyhE5XhYmcJEW
ri6w9NeIRHUgEAZy0s4ZYOO9IWK5tVje5k/0a7owFf9S8E2CsTaZOIQi3kWUg7kf
humMRX1C39+kAC0VEGP4CtWzbHS+m0KIPwLsPcm3PH8WOq8IQ2Ntz9xDTfq2XVFz
l1ZONNqNtNkzCs5+OgZRtOCJLEvb/bGa0YBGjJTwfAcVHwXGeOPNXVslFPt+/bYg
UahL8WjstjWY7OWtwfGEOeSl/DnWrc+4D4SbEGtKafMuWgAR0rKo+y4rVmtWdS7m
U1dfLB1F5DA7MM5Dofg24hWOQM5Q6RpliSVrH2Le763Dof5+YuZyTl9WVm4UKG4C
GgJoto1D5HHRAH3u0QWf4Mni05xZrZ23x5Dz3erQ3e8lL70h5Bp+dcRs2HZjR3iU
a22eCzuNrx2Ee45+eWVq4zPNqE5j45Un98B80WxyramrgOztHfJAZ80UDmZfiEUa
l5qJQ5VyM7zoT0qz1f89wKsAxEy2rht+eknE6bZnFozkTxhBpYmp/a6E4V14ubLc
kWVdXYHe22+W0o2TW0xoEaCfiH8XnGcOugiGZ1eW3BFCMAqOIlxXq9pLSn4mfP5X
`protect END_PROTECTED
