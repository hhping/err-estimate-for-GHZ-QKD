`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pNAKgrMzlby4CMpN4s0GA32+kWct9DeVNQd+JOIeP+E+0SN1bxD9qL1b/xbhTylK
UPV15w7CmTTYgXUoIflOxXVHn5UVNe/Z/sOHK/OAZevaAvGGRYPDsE3IcoSVlgnb
uq6hkuJATBf1LQGkG9uAUPW3PjfiUYPAfutwwxZiOmAAR1XP7HXamcQoJGvO970g
qH6Rd+LysiQJ06pJWI1xjZoayEezwuv8ykTmNzxiGdEADAy3vdNhlVgm9vf2yPHv
eeK8N/kKdP1zt1TLlIUkBbZfLAL51haQaEjpp4HrpVIt1B1LsbneSZeNTRREkcCF
O1COVA1pXvCO+MDIeg+P1GjoWXnkcnrLH4lwhPVFZFtkMpvZMavK5AFLjKYz+jBi
HqJUkX0SVawWb7SFnhNx+LxzHlHdnZZhnd1z5dRRlgYm8/J73cPWLabJkFh/Vj6Z
9ArDzUs3j7nN7AaFzHR/B6r8MtW41UyLBKZyzWEPf4WOzWKBGemfYY7T6qhIFTkg
X4y7DNvpiPclw117Hb4jqtIJRHQXzSDJfTmmmeCFe6vJFUzjyVCLqyZxIf25AWWO
7UE+ZTwmPjVep/0gTf42cXBU37REkReE+BlnkBFL4E/ttEOzkzeyO1NKzUZE5TDX
nzFLb6Or1e20daiJzcAJadB5tdgcCIcp77BqZkVqYe4Vhw+NjFoaCHz3XZVwgv73
gJEhAu2W5F2Rwtt1Gnh1QJYlY7/WrGGILYuBcYB1VK5lCv0m4v3AtpbKTCXxjMaf
t0V2bxEDFmSSJmD/rRnci6Kwx6i8RVnrtbWvtl3hLDoNcs0u4oWUpdPhep+gJsMp
Zn2ZkqGtHyMl0M73iRyNOVQ/m+F1phL6flhCVBhKWzUZ6cRC3Iks/Brews/T/4hD
RssuX5hGzU1xK+4zbDTujkmkA7b5tMdYpJII7s9ErCXG46axRpMCq+0VMuoZYOGk
v7QRGt/f0KC0qdUuHSJwjGrsOOTwMtr5b8I/lPXCYRa6O3vqnK1BN7jnzdD/seDT
Qq6iqRDKw0avrNgKjSQxYVfIhQiTgy47EnbNN8FnTPc=
`protect END_PROTECTED
