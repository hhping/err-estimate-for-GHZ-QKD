`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uFwyoxitASfzDBZV1FT9mnuZ+QO1MefKSuZXFP4LjOmaG63FNoPjrcsFvrr5mfHp
FUgWAqDZJZHVYsCq88qP44dhy/hMT3R2m0V72qLrDoNu6OGBy/gMVnRHpFapfnX4
/qlytz/yP0c9p08YCMS5WUHKWhlLI5piPy5g4LWuV+ZPqJTz8bkTSDeBAl3ombwg
vjVhQuBMrXAiQPnRN8i1z/RceAejTOegndzQePpr0Vd6K3KAEzJSRKAvH21wvV3e
wO+CWtKM1lOV1RjgcpzRzm4ajRxw+mkN/9HsYHEr4gKU95jSppCEWSC5oeIP8ECb
ClMdlAswi2nfmTbRtYNJlxtv5onOqTnfG5vcKsjoHq31duxR12jTbTduKGpc19Fe
KkIzBDgTv9VJB192CyBJdC1B7AEJkIdWvjvFj+8vrCn61ZF98iaVH3BUkt6EadNe
IbqMrEQ5p9+q5aA0vMHPmtVcEyQ1cMLa4nx5yPNNkbVd+g+jk7rQQS5Z1mJRJU1E
ebty3kHK5J3VwKC9+J4lpUiVEpoQHEXCi9GwDM7WR2h8F5+4DAOL2csB8JKd74iU
TMIl6wz76CKxbZ64JSThU2L9uXqmgrrlw1v6DSk4rricscoEDPxLhFmDzHP5uRGE
p7fhf8mpPiUgqT7ohG1loerQ8Zcr3eA1Ev74BuVzNKUaZTD86H5OSnRH3As3hUZa
d7Mzy4h3lUR7qaWC2nVRNTaoYpm/y8cwxFOhigbqiLMgH/jpH9mZxCsV6S0ysxi8
uTnn+ORkWPo0K+cxgydB6Td2RjfJ7ZxAtLduaR5TgdcTIX3kIKiaoJzOlIVFEFvu
JL6oN9fuP6iWS/3rovGPugQ9QBcZSPwWBV8eDeB+FWd+vursjc99bAXkxX9jzduc
e/iyfKweZJSOGNeDYyLZDaMcTaGgz4FWI4sof79RNWCaYO9soGeZqLu97JbXoEBS
6t72jiXBSuX8jwWxsNenVwkW+8SoY0W7S/HgxERXEb73lqozMfvi6lFC0pjynP/Z
z9TgaK5gujJnUu2+RKQIRzuJvYIlD0xwbz5379vK1DqicpY4dqpjxsgU9kHhQOnt
FFVixeIrbO+2WWVVGuO1wIOv4/2beopTPkrjVegxUgaMoTSMmGUF/GbY2OR5Xzy+
sGs60WElZR4G13ZWreDUuV5uDTsNEv1gGqwge3KdrDJU+BeMlF9dBFXma7zLgPAN
k5c0grE5iOJJLGjFve0hfxJXKjKbdiqPyvwOCr7+MGKmSBgPMUbJeuY8XtGOLmET
QTZZXuLVYnPZmpSGqpgSvuPpVeNQrMSPtappW8eiNVQGZsTcDy+mPAk/4Kbq55oL
Ut0dgUUZ4mKCyKZ6HOTu4JlDRae6CITPmPjIU+8zpl3JFZVGqYGc7iXBIvG/fztv
Bupoop0KcMKv0deuqNL+lQ==
`protect END_PROTECTED
