`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A0JfeMmj2Vw5tYeHgcND2o7a9A75UnPJnArw4J645SSJ8aCcrOU9lvn22BGN3grW
zUJApHyTkGNU5271EDY5HEDDUYuGTvwEsD73ZAAzJovflMIxxOtwZYMvDwfgbeT8
VlHWG3HVuvwbudX8b2Dmc3GBJAONMT2TAopNgTBPAVPvFwd+HGEkmf87AhgFKqZF
FpsbzVa4YVMi0WhoO25iI+09fDXvXVEUtCrcLs96neN5nn4fJ0I0r1tsGIAvhsYZ
dNtvyUJX0LbooazvZcJKkryE73nz0mHxYGvV/aPe11uqw6m0LaGQWoi78vco26IS
s0xYT3HEc6xs5Ihw0ui5M2cZ3PgI9HqCKzmtSqTnKsn+wyYQaa983yjx6HrYu7K2
VZdJE4gvtpW2D4w4uY4fHjGm/W7o2a5N/ip1fOHs39WkTVAz5MUKBRJW8HahgTqZ
dscHqI73RMlWgYDL73NpGVkLhsOKsM/W32ACZgjyukU25XdF5r+hjmTIuNBevM3i
EHrtfsAHJvsHnIPwTPd4FuntJU6/blCrSmHcru4pkR8+y4kh9sACVeRU+n+e+XqB
FcL/eR/hwld14+6izB1EwaUmlpoEDlsfm0tc1OWLVzJwhAb74SLL+G3al5ntffRw
sADb+f1IFiz/7ppVZCUYxfsgdMljEKBlHXCrbVZGkKjtXfG9zfwFneW+vmZ9KQOk
vxnQIsZVwKyB+DgNVnswYOihTxUo2Ok1uX4CfjN8IfiGSqvtZkdHZ86j1HcHaixi
0DqBylVxlDu/YKoNHqDSpnGYiGB+YpcSYNQvUEcsCwQ=
`protect END_PROTECTED
