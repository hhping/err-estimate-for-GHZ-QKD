`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EggYYXZiHTISK+h28ZDE2TlovEZ1rWYzmi8+JyvAhvTm0uzBcZcz0ClzdOf/UVYn
yfd2hsbZ8rO4hGSMaI90YiuMw6tVkKrLThJ3EEPZ/Dh/nLkymjmYAPHe7DUh3m+m
xapKehlizVW+B/697YMYctGBxbkSwj0L/dBSHqVHkrIWiZlicqSRnLJp7NHJWK6F
g/azlg14OQU8zyKMziGkC624U15zMX26vw0j1yO5HE6Y7YF5/aMmywLAPHrdhnfj
8Dqomc6NPwVAeKOSEWNU7Z2H0Gj3GkkAX7nrbhRpQ+fCRdK3on8Uf+ZZCz9PYzrv
S9FQbVh4OwVxUcIkevW+ShSSLVZIOgswC3TpxCbui8Gc/jPGB+BSdxzmJ2dUQ+Wj
scMo7+6B+i8WrFtQ6dnxQyCqUOlAYKiEW8R4WcpXx/MpxcMjp15Emww9CI9wf10G
soJ1mzdtrRpibJ+aK55vf8ioMTSQCnMWva4jd+m/GLP5TKsvLJJYtzzXXOh5Hx62
Xxifn4jYKx0drVeY1UheHMRA19dSquCyI7Tbt34qG7ICrPXGNjQRzivDYyD+j9D9
JpDYQcD6hGKJ95JK3ZNRaRtIarGMLBlmT0iQmZ2lviaLpIRZynZ089YacL7iHWh8
Dt2jAGpHKEnVccRBJu76A5D3NF2ZsYU0+sdMGcD/GE4HuUN8lWMbYdMfCSCqdPUN
9QHnUFcNw/tH2IzJpowLe/7IGLic5CsYwGfogq/3QVQlljQW9XV2uaB/1Fb4H75X
4p4nsAVmuXFNf5RFRKZaU1AGzoyCCNHONruD9QYei0xJp/Hxv1557AmfWG89RqRQ
L1rAT9ZFb+KkCvzazb1JNsRVRRfk7iAZAukE342cXs+eopkKwgdDkFU0kRLxO1By
gCndcHPiqkXiEYEwtIL1mFh31VsPY51uM/U4Yt2KxH6EhOBGqI0JuOiApl59HX77
3zgjrdtB+2IkkqfNQG7R5zGFjMFaLN72wa6QiWpoveYiFaZv+w/t/r8W0QgVrqSQ
G4TE1xpkh3a/Zz+D/VGey1E6M/TrXYs14zUFJyaNEo45wBVkTl+Bh0faoAWLtUZt
IaZOUp44CsuMCcWHoS6OpRyTlY6bj5l7DtiETLBV8CKVZu4rCeBdkb7OcZgr3P7S
8DUuy89tS+sLHeOLdWC5BUaMz+x4lYxDCa16/meXWTZ5ER0ejoAkb2sm2NkDJe8+
J2U6nZOT2mn8v+KjltrA+AqwaIy53XAaNloGAOKAmn+gf8eJ6AIrpgza4S3pd1lC
AZajJ3NXnQSqWJDqkqkFXEkE1JoNnGlrcxxK4dScA99+fgLMS6XLFoLylgV/dpGo
1LKj4LerXBCXhLNkYvEckKwssI+UlXBjBV1cPnkL78+BhWbSxRxzui5mjDf+snBM
M6lcxa/UW7rYgTHn5Nq6EtWxn3pXqUAP06KDkHOiR/gN9Du+RvsCAIbPKU/jNAYE
6TJjvMSijIhe7qfpg/h2rS3RZk2iA0ZFCr5xwpdvdhVbiUMlOaoEdfLClPsNUJe4
i+7XQWC+Y8NGBVpatIi4Tyz1zxikSHafjLMdhOhZ0c2y+unCI3pi5DQc7VnyPqHi
f3tWWziF/RzXcFp7fZS1kmWtcdW6H9NOP8jRSiaxKD3OEwlceZ/y8A/+o+M3VI6/
UElqG2cWuxkPPoGNaYS8zMXWpnLgw60M+oBAC2S5ddWq9FYY9xAZccn2/k3QDlf0
2lvpjpwexeiW4/h+0wriHVLi8h1yGzgwpFB5W9snBxnvFK75NCIkzZ/Ff9pPs6am
1v9wlJskbvF+1WUhi1vt18T+m3ZmofoSHbrX79bmgHS9/sjxamERhy1haUBrdFBm
+5ZXlE3xbi7/uYi4X9FHLZrgpfjqCkgzZCeghu5nFn4UT92xdekBPqiqbwL4MLOj
DNQpNRfHu6tteRxXs/R5bJY48i1bIGxpU8q+W5DnAY9QnhM8WcVOZWSdSrD6Ub5z
0Rz1gvFe0Gn527ICHr+X1Pv3sJ6aDl+/+sVt0idLee2UrUjd4SAE4nak3zxTFHVl
Y9DDJGS46uTdNsT5V0A9RUAGBQUTXnMHpXzH4VuSZNNgXJ5jH/22nfQkmhUd4pvd
agroTBKaBDnYwsaZfnShZbfjx+zX0F81bU10g4S87CVuzDcZ1LhJr8tjNS+oUx79
Uaj2zVk+FxFg1yn+XMCsGnsSAhTfpT3xedBj2okjmnsrLAk2eSAB/vBXS1o0NFB5
ERdDxKSNQz4noTMc84GOxVLGKemqyEUgYYJtS9guwFo=
`protect END_PROTECTED
