`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HuGEcNR+zGW8fSlXiNLm93F26KKHxigcNDLYD1ZX62ieCCQ06LMS4QX0DdQ/HDPn
6PiLedDxFi+2M2Wg1H7VcC7DIXIFC5xvGOAteGHgtoZvQ4j2piB5GW1mO5tenN41
tKAvrgwcPfhxnvq157eL6zEK687xNUuDaQRmu1AzrSbuM8crRZBvQi3NbNVf/7lA
Rp04K16SF658WLxStHaik7D9C89D+hmUp3qddr+1gQveZdj9kaVAmEbeLnyuagb9
IctRcJkf+A0dAgnHrYK4uDym7snmvfo5zdOYt4LJZgdnfv56CRd2ZNCZxOrkGTp5
rtwImZD5xpHMdfTUVkdKHgHOz8KRI+EvCMi+c1M5SJsqneeSTTmMVG36dHl4f/IX
EyMeQMliWRS/EKJwTE5pII91+95mYx+Hnvj7LdKCf6+zQpCj0NC1daOUGPq8ekFb
mpbq3Z7IyT3L1mMduW7ScZ57akawaLBd3liHHjUBAZ9fLazWNSxua0OliJGeJxHR
aaWspIQJ9cmj4bQVYZqZsnK/pxOs2vT38XRDORfIw8wQ3DRixQMRGagSMHGTkUZ/
uvHOerY+g6SiVcsU4OWmeuVoi4+qpwjeySUPKtm6EyvsHaJe6hCjR+j37DgJnXS4
mYQ8pgwqVbxFjNbgZx36dAwSSn+i9x/IN3aAQXivvPK2EWQRkRu8uWSbiU2fcA+q
AcTYeXe0+dV1Rowq89/5joTKDf1OiKxLLgZhAgn4BN3+erTBtvXEQe88H8a/kCb9
BX5dsfEpCimiu935oMmJJKu7RJoVT88FiyjzcY/IP9INJ062I7YE4avuUyFMIh8x
LEfI2P+GLF2Shs/zTKJ6QNZbceRYXN//YaJVfcd/nLMknXmTBu5+qIkO7SWS4YE4
Bv7KtxMggFfvWVwkv9HuPBgcq9WyFZ3EIEwp8coMyY1ctFhnnUU5fD/FMYeU5BQ3
X5c921WzpZp9S1UE5IgKqDrV4DLQF62WDFBuJL9Mwc4=
`protect END_PROTECTED
