`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGJv68f4spKlrD+PZimL0QHoIRv8sYsAm+9pQDUO57ScBel/dV69Pt2K7WZA61mu
uysEsuirxvIzfC0muG1/Fwtx44SBCjoFI6hliMaPbtPuZ0C6pP3k+v5MhRVUO0Q9
NbcG3tGl7SxIb3PnyA/6olHQCxoEfxggYiIdeTGHAuLRSoegPEiuXlTE/7oZfBLQ
ujFKSRtXqIkC5PYMcbeQ3iHGhFA6khpA7sXN948iK1JppxiPkqT+SMWhvkGDP5KA
lBZ6njaDGaX/tmLa2eGylc75E/Uj62CBuhzNKNDwgzZ4nSyXkDAXNAINUxdYbz+2
3GHwBnxzFdd2c0bUHchjimoZPLi+Xdz2mygkISxeAR6r3pwJX+2PvugExjiwkvFp
eynBw7MqAG9X6IlfaCDmO7RHgo3eZ90uFipzE0yfzjBxWh93GKOFqrJgsBC7RHxI
Fs0t/93Fy8JRxY9KzOVG9gynVHnDh8GGo4mq/8VvPD2jQXTpKLe/Kr1D/CN/Y9SM
Fw0jc1ckjTqlQh95mPYinQ==
`protect END_PROTECTED
