`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uyj/LK4NSkcCf9g+JkxPfICoXbAJFBwTkyhNNDGjzRfUyA5S18iROuLOTfzktryL
rE/eNISjUJU9k0EMfVBYyiczk+GPOyfVeV1X1SzTwpUIq3Iks/tMjWnZHiZB0kbs
bghn9CyUHraRbXHqj7QV5sKKQMq9jXkZlpU1UxYznC72A85Xc2kJ0VpVRjLbx5aA
vB/CSJmC+/9tTrgjQaPpovCzA5HLyEZZ/uCc4qAGnTuVQMQIqKLP14YBe4zS8Qjg
q7HaJrYYeqQPtxJ1jMe7SbkmrtjPiQa23wr0tx+Ir8v+AEQ0vVA2v2pYnKfLn/tm
G4OUf7iYJxOPMtcuhiF/cZ7grBHqdTa+ckyCsIzcRbaQZsb2Rs0SOfQa+8Mp0FEm
/05vmbhgfdiKGFnXXgSl4kpEOa5+ukiYmMZw1SmNIdWtLuYwm+dHNlLhVteu8CWD
+FRQu2H+6vLuJ3bGR70BfI2Q1VicSs0KmdxZQtgcllXD2ERTgfTrrdbDdHA4Ngkl
ojH+79b1x0a6O7jPYcSWf8Wgjn6Kc1ZZCfCcVd/0rVFCaPuJG1L0PYyDe5E+WBXT
IFOjvOVRlKhw0hoOLfPQj0KquXDWMu7Xrixwhx5WfkJMpFaVMHau0XLt7UcfWTpb
zuMFbVqz8mggr101VSaYdz/vSsmMOIApH6KhZTphJydjYdSkO+Z0jCavCgnbWH0s
16jFKynx4TA13+o5j3+QH2g8w2Gsc5JuIiPQlpxdDGIqswkwIMm3ckW4gg2dl1GW
1AfQmNty/EAuWNuXVdt+fVRvApBafbz5nbB7ZkaIIMni1+87RE8h3G1pxTsGnjsV
yHUz1sYUJw6AWKly9DQWEsMb4gdpLWX8E8fYK6GOeMNM4dYfGM0Ygl9crzyRsUjv
X1kn+tZzeNxPfLYNS5wzx5iqgFM80oZlBIc7QlTrG3qGNyeHPzgp2MavDBqlrYv+
PUjg4aJO7RtA7CKpxm3c7W/c3OcWME8vzDxVitvBQo1ZRPwEjrm74MJ7uUDgsyFH
sqLrDYtCJ8t7hF6O5cVqVMgWUUzs1Vwo3R/s7oRJZ3ISVtkAA1A5/hj0g8DM/mbJ
am4sDc9nFMamtutRtqBwPsNfePXkOHRpBf4tKMKEvAHeJ5ES0JShUBeely5UsMQT
gscLEom9oEWoYWTJHW622JxuY5MzJM32kKc4YEsyIIcrBBFEBOGLG4jN7k/Qba3E
ic3Tp25P8JnmXxvR9+CQieSBR4AclVhf+pQOm4AMUHp9BLaKMv64LLMPvAfqKkTp
u3HjhV9PLEW/MVH7hRy53B0wJlv6zHv1xYWNXRdTteUtGbP9cpFe0DeclQgLEhvY
5tCiEUhsIIaAwEmYa/7whMe/sZTGf9EqBgXu2xXScid3Xm16KCSYs2JebZMoGMX0
NMOdoWcndmkjvGSrh+lTJf7NsKOD2TjZzISv2FeV7Tm+YQs5Er5FTBvlkyD4+e8X
s5IhKZtzd4qQoI84yM051QUWRj+2q2WVINP0/uTxTv1D0pUXPSDfMuLZG4NB5HkW
SBnnnkMz9wllLuP5kSRcv2wMULMpmmUaCz6EZii2pFblz84aHFJV7VHsJhs67rZl
QUATJR6Phr3PVvfst5AXlaOaytXcSxG0S3bknFLSgMVYFHQ8Fpd0eXzLpunY0kdC
tzJF4mQW3aMRH/kmq+1pUkj/SmHACDxIF+3lf/wxHEP9eo0v7dSiMkoqPiuYdNdk
H/h2/q8rc12fSNPSvNTGTpZ+DOBApYEBVpF0ooH3vc4xxsNfYoAyGYgJk71qt2uG
CA9rrtBAejwg+DoqMm7avd615sRgBxlsPEE5rjbBMRS1E6CU8uxgAr+b70cws7g+
sagzNuktcNSP1MaZveYNLrIe5ziGc5s0J+dIEXGXH1jINZ2soVO2V3FAMGg0f36t
GP/ahBD9TMyaAKyUm/FGFvPdxk4hQidt+2k/ig2LRwPqfV94ajmVN1+9z8OdJjqb
k58ywoN4m3Nkj1zxKCBz1JX5fWbCl2ly2LtMY1bhDOnTk9u/ivxeBPZ/wFlVj5uB
wc09jrKmdL9LlFPZjOOcAs+D5jWlyjNP2/+P+MLN0P5hR+bpR0Kdv2zR1v2QEoFp
CpTmZmIC3eGYIaI5qd8GGdPkSIH9Wn0afSs3pvCTOasHHEiOoWTY8Z9fS0/YGxma
rACXNBQSZuPcYGRRNwx3xidP5zQhILcxp14ukRIi6TkvSsvapPx2NJIiaoOc0I3+
MKfOgoh+7u6qnJvnwq8vv/GECHBRvoAUcq0u1Ngx/V8ixtT4NLcqCO5q/WXFBa3N
fQv1fxQ9nGNHLiD6+jVJyA5EzFQFhBvYUNIM1618E2DMO9XatODqnu3UrN7JjlXZ
`protect END_PROTECTED
