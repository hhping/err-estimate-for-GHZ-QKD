`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PULV437eDGJXYzXLG6MB1MoDvfolg9oF0TvvycteiZyFMtqKl5lKXTzHUs/WuZ+2
ePBAUU20oCgdU1Pkqxv/S1H9md/FzMPCJmCHwZTYbb+SU/kUqDE4InNM7NRnp3u2
VrTMU/mHWhBwFotFLlX/sYh7NarTP12a2Yy4XSIiZZvGQBglK4EBkS5dS4qb5HNZ
GcK26pxMI8OjwK/bFCLkD2iM4MgLI4YOrkgJDeS1Jl61Uzo8OzfaZqD05d5+pSEn
AoYFXfzLJHvSIDDMnKPQRxwG85e315VuNQi+VlETU1qdHxI2bPgcQzLd6LCYOAvT
KG647rJWX1NP78h9lEu5RPwt2r+MyqzIhUsSsAxnq4bLfzX0/IcfnkXsWDK1+Ezu
9cKaEQUvJhgwMdIp72qPzBDN2zSEpDo681oEBESsSHgdKkULg5OsOs0M3/B6veRw
LW4uKm4ZcOoOux01+vnCBgo7FBeLn5UzQzUV5L8X4i5M0i3rfNNIS4/aJD9QhIXc
g6mMjV4VpNI0j6e+i5zMCjEk9mmr+kX4EuXJDsdhGpmb8y9gMthYD7p6sfR1WX0f
JllZJAHP9R9CJTUNFD1bgCFh8VzvFUJnRGnssCG6tK0yoSXL9v0husSppFiJVVkQ
O1efDoSHUdPVglH4JXkkGvWkdaTh4Dc8gLb+4pM36EXdcJZcfa+GJdepFwWJ/ptl
UxSzCbP0XUhIH+cjWUOkel2BOe4Qd4JvGGHkwQW0rVR0lSCvFg1eFoQ8ILV/D6hP
hAxUgDN5VMVUa0WgSJPUJA==
`protect END_PROTECTED
