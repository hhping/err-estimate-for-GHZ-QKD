`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
okC0ZWyxN+0GNORKK2j/QHjC5Y363eIUC1ks896VfLJg5LBc+CBEsp0IFj+7RHU9
1lCp2OwdiVSjWtBhDDAzk6aitG6pBosavYleWhvJmffwR6nN21YH5BusXzoz8kfO
pFaC6dK52Eevszj8aoPq5cJquZQshnIVpwq8RET4SmfYJs3u2pQ6G6SbtJ8SIZ1R
Vr56FZIbBendulRhF9pmD/XW/Wqe4ON7nnRPAmyOgKtXpXe8LK2kJKY/xi/+bKvr
BqIEbrSL39Ki6+tm4oGXiMTNO6Z25/401/mcdNiE44gRviQjnTJfy0qJCcdtl8Z0
jvRQbNpJw/CgE0pQs9McuQG1TmAdBRA+Qffp+hc4V78x/yGNZfdRfJ405RFFni/i
tIn+l2QjKzPhN1PH5m2n2x+lDurKrvMxgLU93GGf+Ss=
`protect END_PROTECTED
