`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tk1YO3jnkjJ8ILdYwBphHGexCS2vPgd3R0WLyPMhClhMCcm7UjryiLITBRZ/hPwF
H48ZUh6ksGkMq7rXlTz87LSr4Q+curcTxLEhrKRxWI7i2/BvJwADtSDjdzcP2HCg
/41JYbWR0kgvG4aTx+iskCzRj6lQ9cWCxAHo448FQ/F1aXwZVwBx7gXeywE+gx3a
BYkJ9m53NLbxwzlnxt35H3GgjG48WrN3ZKJcQI6niSVPGtX+Nn2MYFrv2cWvIpXe
dbCitaWa6uDwylA1UDBOhYsCAPsRcGTSO6erSlYsZkUkHBlStA5JXpQTr0ty5vRo
MuRR3a2vNPr5OeAMRUlthJ9/pJfQsEcsuRuMQV7Yt1N9dyWeFb/NUdLr8Fs9MBth
7HblnqL/vk6dVuRCJmhfmIM60qOaFLaREXO0viR47+eJWkbX3kUuDARiPkortXiS
++lLpupY4mRux8gEvBXs0dlF0LtK9RA9lcuZo3Z+v1cEp0gMQtdG2McrwBGd4mKQ
rcgtX8wxP+j2/hZfmOHqkxWT5qrabBsxKyka3XuGwma3gTMx0KMeX6v8YAtntbdL
QUr3dn1BXpr6OvePV3bK9bESALUILEHMnqJr/Vh4t3sLBVQYRkqPZXDNr6jCAXhP
oTJVG0nNoUj/t1oJr+mXdplbWW1g9+b/Gk/5Lt4RNbyP1c7P7qV26QqPRAgTNO7U
kjnhPzvRgr6dmFhW36p/o2xxkiyowFqVyJxM5ciJCh/m41ZnxDTZ7gAutA1Vhma3
`protect END_PROTECTED
