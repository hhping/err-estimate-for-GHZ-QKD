`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0PVxjxVqWb+QhrN9cmdC7ivsa2NDR3rdPnlfIOYa20tgtUHya4+LE1UIDL3Dctu
MCVGxvcSRozoqFgU2qwz1aAST6F7Byhd9vqtuw1htIMI1LJ09A9joztGTYAdGwqm
be4BL3Wq5IAe1wVcFkZGAXLQn7z1Agj307JbKQ4PT1+LP24kR8BaS2/K8nSda3to
IPNzkQiKzUalT8IdMEq4ncG0UkLF1+p/hJHvTayVa1PNkf0RS1nRw6afcWwhAEew
tbKr4mYqWWCIzBfMBkh/egxa0p9hItweHl2/zcfQbQCcayWZ13J1E/IgSHdZN/Oz
r5fMhidA37XWpOhCCUe1i6xJQHNLx3lVw+i78fr9JcS22w0419TZcamLlO3cL1iJ
Nll3GiXnsuxKNCe01SOsbFgzbxX0zwsyhPXysCFY0fGo7AnKFw79taIUprJFPSDw
XmtXi3UmbtB7Hh86/T1v5FxZnpLNy4w/2GccNI1Az4RPDi6yuw0bvjpv0FPxd3mU
Uh/b1FuHR6dHvvgt/aqmT7tUox4lgZ477kq3m4UmsQgml+Vvh7WpDnSrVeGhGANk
r0JgGynwI8dHkPc/BUTxthqlkOjZU2GEsVausPDDfrDcawwdyd3WcFmOl9ZeoF1J
nD7XHoj5yFf8HTOATO66kQkFCtLKt2ZZbakm05HGNykievhn15U0+cPyCuZaPJ3K
jPdxa+TbMrF7Rj4r0xwF3g5nEaac2yZVYDpslKeJOlErAc+9qww2JG4nZLPKthyu
2q26Wz2PnuyYCrXZGlIqWLLkvh953cRuGzP4eZX2+G5sVvcUdJybGj4/hqHQKhU/
JGJcpSvG18Pfh7/idHhwlI8sAR0ZFxRhgq2YUQmVD5fU/bgmnUB87Rvjv4Qez6Pp
TlkWCR5xIOLY4TvF44drN5FbSrb1rOYjFaelSpffR5p8EKIbOVZYVCUGNdsnkVOc
/JqrXi2dI1HRmTJCF6dXW75eUlPN4T4blJmk87ZwCF+xnDHRFIC6hxOmmlq6lLUr
QzALZnn69Xl7kz9XsgW+oTZcTN5k25PKXUMnlFZfLaxfsEroqJu3CYiZJrzjZq5q
rvVhHyy49R8fK6sIYKbMYLe8/IM5WQF4Xhn2yB3FwRaMquc5Z12njqoe/6gkF9iz
RgGDIb0Lp0Slx5mpC/5ps2sL7JvVlKgSO3VCGYAGwkXuTuUe1jOGjvdEKjzCH2Vn
dCrz82rMVTViXf7aoYPPem6+nDpAmmWpc0xPd5DQQKqSSKmU2iMu93IkOn3R5Chj
ZzDJUjOxI1daTotWUqTUrcn/paqHM5v26UBSfXRWqMErzMerTbTFhDmnqdYRskeb
nOv38+S9QzE9P3EpYvmdKo9b0wxV+fmo++iujDlk7nz8YXzDFdmw/AoAGjGufEU9
3PTAKBRTIGp7AqCvUcLcJQNzqpr7VXM4AMDUWkUAAMSQJAoEtcyX84FiSkt0PfcJ
3qMbCoKWqJwDwUmjNfhMPnOiAyifHOfGodSHuhey0BatGZZ9rIfhkaIZ+0IFZCcP
uzlVfcHdnWIPznpEg7BCFJ0zBKOPtXzo9x8SvEo94HDVer81U9wCHArGLFgVI2aB
7KAtYacz1NNVAYRdvXVsfux1ebruncpVmMmhTWBWw+xJj+74vPXmA/685MEoF4aX
Uc2Ab+m/k92/qMF5rzhFNe33/09SaamBqIZHJAwWi4yxwCMWQtgPQK8Fkg/XLOEL
X8sGlZSSd6U4iKe5NFbbvb0eJpcAanE6EiJZbHqhBAP+mFcTVXVNM9LT3NFDgm/j
vanHasG+0KNBllL8+v+qFYaa2Pvr/+yjaS53GnFvVIlwkNzKf2+NB2MkLpK8v7EL
ETX78eYgwcHHhe2otBU9fcBwBJP2MAdE9SypHb+Hopwm4dTK+pH2brSjTWLIhvQ1
3wpewUAp4n46U5pyR1uj/VI+XTrHhb0YM5AzVKgDm3HNJqr8GhWWtAqHAikX5Emw
mpxU5uS5kjnOitE3GBaXLtMrutPUWGr8Qt2mJlqsNtjRSDeaDOfqqujT/NM7cgfD
fky2xB7Gph72cn2e/LpmpV0JnNCyi237PVFpW9KpeJnVl56JYouFbK/XvyKjH2MH
OnpObKsAPoUTBOlD/BKLZGrvy89gL/3F4DS8SBKF5dvUf4opdd+UMCUYOkhBg19I
nalGSfuFJrqQ5i9wfSknJ7uTvW37KuNFbzMXPA0PXzlIOVz44NgvZ6Dg6nT6YdWS
30uHr2fVIojFphTkRbPrnRJwa9p8j4WRQ6ZB/q6ry+TR1K3zbstV9bR5FAJqTK9k
5q7eRbKYU8iMzWHP03brfFixDsxQQGtWZpT2c3+oEBShqm4Ofmf9wh+iqy7n2y6d
QGdBAtBKI8PniW3AEVajSf1q2lGl0/prih5tK0Iovqa/PAwV/zPwjmwnpyw8ddOe
XtbW/J7QP1Elz/sqeAtfif5HIn84d8yCbRBNUVfb7R1YMviNhvXQ36c8DaJ08+yA
/XeO/tSMVHF54ynnuX69LfWVe2mdRXAvh0YgvPdV0RHaeybaJ1pNGjornd4kw7bB
or9ng0ZIOpwCLJY+WlGq7BhB5z34eO/5DdyOvBmh/kvibI3tVYeNDEmZEZeHB4B7
EeWmu85W2pZNvzWDFW6wWHAj0LIvhvmkS9f8ieOCkbz1EP9tvrSKRBSDev/bB8Vj
u6kK2wOsHNXUgUgHh8KFMDeTQWyFJpRZIIe6OcPfiGVZacgGWdgNHQ1AG9Vuv/RY
0sC0OjqjCgAxKXXLaUrlVKHrCprAGllvw6R8wkaku1OLMRryBGRvhOuGQ/12S7SA
ZHpdEPckSawJdy8u8+PeqcXnTvowh6N4jxjvkCptFA2q79qz01sxPzrDdJ8gNpbF
NHnuSdbxjOyqbbNicv2ody62wb/tE0U6K9bA4eBXCmmgAdIICFxKo+EF9XNVslfE
zsnA61jPJOGC+jXoe86AfGCcj5/+FB/gAjqfyUJU/05AhWq7gWrdEhuH5u2rvPjR
8H+QLvds2+toBVwUeN8Akv23Gx0g4Z8K9+GOlIdDmb3VNxquOI5sv1Z6SYPd+FGQ
yLlybBvkXRG9QtknJ7aoEI7lrE3a0swUWYeXCjyn9+YqBhJV086fcdDQ13AnXRRl
R7Le41IwmYvwd9gnrCbHTNLkI7FLxx6Rcy19bhPYMo3aMbLxDkjZWcSvXBrAmL/L
ZPd3dlOtjt9Vwug6utSKehZe+HeDWY80pqDv4O7C5tpWc7K++MpcsglqZ8rSu4no
wem/ffsYATR8U04s3NGBB37UVsclkWdQ/rLOWY/ljQeREUJ+2pLs1TQgsifE3Xo9
WjDO/ETf82KKePE4LkwYT0CqJVciqtzdy2NmAagna/6PDx0P6/9n+ONMCTHg7CI7
`protect END_PROTECTED
