`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bFxahvDvX1N+q+NJyls1g0EqCfmX0s3z1ei/CM7rECSC6Zh2M8BdDGzjU7KHYI8
ENLwUPEotKDil/j5Y+kuGk8zer7/LTp9FDfHn+HHNjMAw3bRNfEirPFqNZQecoHi
wwJB+PawXCMtVPetNzY5dd8nMEtWo5oYpgqmdrKx3FVI59OJD8efr75uGZQZHC5C
dexLm/ufw4IKenxsOj0jlQCiGQs0oVQgvKJRJoiH5lElvK8ijtdOwo4SOtg84gKh
wAu50wLiUajSf05iPzSHEI+TAFuyW7PfUvS67NwueOMKru8b4ZlGviBwOn1PpgFK
S7uzK0dQAZaMhYlOAdtGsnasDJbWCWW7+nRfctwUXEpyPQQV05BmDgz0DiBEffI0
Qq+oQpIuwcZjaf0KuCypbRwzOrR58ceRtQHInjmEhq9ZRko0456pq0t9D2GPOalh
A04IcQTesNVJuyC4gi7nsoOi2dftAlIe9Z3hreClAPKUvWmoM3NTO7sMd6v7LuxF
fZEg+x8Yq1wuM5myynMftWysVxvNSnNSIi5UBOBqQHS4RPabwlG9qyba8n6a2OXH
0jCENX9sk1p8Rm+v6jDwJm8HdScoQ/vHYMVJ1Q8zGD8BOlzuG+DX8jZb5eMqHRCW
obGq8umlRBE4qKIZsPoXxhG70zMTOcOV+qS7QADUahpU91Y4nzOYzWlucSMLHn89
6yrJ0BUFO2LvLkusssoaZ0757pIBLS4ltNe/1f+yZ9fn8htA4zPDHJnuX1vw7bKH
Sc3PR3DHccLX/l3GyIOITBsDP9AouMcwiNRtAJVRI0u9NMMFMzdBKPR2Ks0PJGN1
gCE2/L3cdJEJqCJWaa7MSu9ZccVtgm6bFjm+5fWpXvL8iX9C3RlZPFYyeeczuDsb
eFokETXUOIulAPN3GnLM5kuz2wPQSpKKPyqlCHBB4JUQmnfomDcRr311i70x/kZ1
P9IO9+xSvtPll+3+pFEv/Lrnlu5njRezNQUX9eu0tDs4N8Ll4k/i0iYbruOoemT5
CG/ZwmwOcw/7s9hPngdHfxDSLClYPwr5/B+7pOaS5SIdP9RwvRTwknZ/ynxcLEbA
SWAwc4O6HxEBGQ60+QLLqL4Eu7+C7sRdRwLflZ5iMkeXr+zVPoMFN+wFlAj/dKPm
vouiZo+h3DXrXtllD/BBFwr9MVnFVH8DQSVE58CuL0AKKH44DOHF7DOcpCtUfng1
kNKwPdQ0buBUm5LS3kaKOp3veG25UNju0L4cDK6YgmGCtSAsycbv6pvuWJGBBM7l
dXOcexoYp5uurLbcYOFIXfDxIYhBydakz2gMoPtfOPC/xCYtpgmYVKFRcLJLZaCL
+DPurKA2BtchjESXgxmHQBa5KnLM3ZyGIhlPFq8ukisyZXLvkl1cOgNt7oMrfKtE
sxIX9nYS1aXFA3EctZSv+3jZ1DgLfDFNahiDt0VW3eQKJUQQamT3cQO/KZi9BO5T
`protect END_PROTECTED
