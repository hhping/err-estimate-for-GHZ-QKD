`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBmnsGMf98Po7cLuiQhBgxAexMa23CoUNzghUvUAZo3c570YmJ3lCFba3fzRGmjL
WmZKKVh0BeZPMw4vA1u5BIeqfAY4spI6tD4997BaiLifTpfO6Rf0gEZ8vfFTgSzy
OZR8/86YUaJOcPR0gICSt/syW7U4l8+O2br6JrZvBMtZgZZekxieSLisiBXLWXUs
49U/7qbJvsAOv5zkMZQFaC/N8Xg3gEIiSzfgowkXs6ebi6crpBXQlX5PnFJH5kmh
BKbGBWWX8iKV4CQUZWXQzpm0YqevsRMdVQoPvBM3muw/iq0hjlcFLXVEThE9O+tI
y6eSu+p2hCAtSYSotvYyuI7iVyuAXLhC/0MFBun4eiW4SjK9SiszT2C++ESdn29t
u2rxBPsVK4v1X9KJROqcDIl7Pgw3MGeBj0BMBmbct+taDH8JzemGaXPdOf/vhAds
9mPhwf67BInvWNqrLS3GQX7T13F9Qehyxf/xdkTD5obhfpK7bXovkU8iOPbTVyVp
XXbyRniRwe/qAkNAo4tXztbNvmIxtqAPjUbpFqvYzFHUBVFirOOahI/84pM8K7Y4
7+i8BTJjv4tjywh/Oz/wmti0Rga+BlTiqdR/TNXY5/ajtCQbg61FDtH/wEjMOFze
3XxPDPA8Ras7tZkRR7FKrZ3aesWDFUGI+PO1V7BfvTxlW64BFVYtaHy+kp2bzrdC
AyquuTI73Pt+FPX8w4dNur6qKMy359sqnJommgtgKZv3C2nZVYO0JP1Q524EhgZ6
`protect END_PROTECTED
