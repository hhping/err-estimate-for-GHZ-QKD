`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ebuh5vXcRXpRX9u3JTJC9FO3rX3juOW4S6PtKs9GpTX6NNtOcWSEcQId7De1B9df
XFeUjzdiGqM7vvcutvNrQzBo+i1JjiknlFTvILLULpHTI4IrSuk7RzI05PD4sACu
X/QjmkmbAEbHKXTpM4RLBOYXZvwnD5Z+YBFj76hM5xlBz5o//fPc+kDtHJVpZpnY
yDbo4IUES91CIsRDofSnlMEFgHcmbK2Fr9gn/SYVQduoJQ/VqejQX2v81BI8/Crc
j1KnF3vHTbgCFn0/gvr/6LmZHaZU2D+P7EBZ31rxJJk=
`protect END_PROTECTED
