`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/QjBzU2v54W5c6jwGK/mA6qvr5NkZSgiLpbbIHN118kNLoSbFJo9EwQ37M3E/aj
k9+nQhRj4V0trcSyv834c8RVN4olq6Mq6tKJOT3wXqNGxkL8kmU597hmOfQPS3RO
IhwXpYPl+NKVceA773iRFPs1mX1FPxnVcHTVEQdtCouiMGCJoDFxKXIPlxYaDeJ7
G3QYiEPuUPWZcW6aQpXaUJ4l0wxbiV2gloqOaFjdL3m+iOYRk5YeXWF8lGnOvBbA
rDIl4S+Lsg9xT9yZtWfkdW7KOF1aaeTjaze8o8hMPZEnH9TmkawXwhEN71rP/Q79
imPPE6itg2/Ie9Q7S0QG4o3i0KgHPdv9Xvtrx/8vixPwZx6NiOHk3bER0lJml5+s
JBS/itSPEcKA++AE1WWscoOFsaA7yDcv2vKlGadWSMJEkpZ83Pb4dLVcG5T3xEU7
1/V77M/xjE2bGOMlKVr68XlbUDftbQUHyvckqr3X2TSRA4KVWJnjrjsGMcejzert
v9ZZVCIdU9fpyMuaKVZelH3kR7U9ZEJZ8wroidypewxXLGPd//UcNtnlBfqjsQgw
h223CWapAV5HT/+drJh9R3SUY+0RVTEdeZom5maWuR0hvdJvk5IRm4qZPhHF+kgC
q5U+z4wggNodkEYM2eDKSD7khcRcQeRL9UxU4A+Ye2e+U3O5g0HNkthlTOKmXIeC
l+BJmxDKMr0GD+KYyeH1t9M03ZGOANK3vA4OTnguVRpMVBLGi0FoldYN3hlMXMNb
RmjxXOREPKhdBVnZuPPLSKQnB32P+XTt3ouhlbua6p9Zc72DMX/Xe7vdBWBxkx81
rwtPVSpkltWW+fSTv4tROY5uEpxaohvdLwqfvjobHv45jDDpmoJfD4DI6ZOJaUkM
sCc2hwz5nkJUXteQhV/U5YZ/D18p4IONuW5Ge9kXDUcs3gBkU5nCUmUag+AAYfo8
ix7fulYR0JT6td/V9UhE4J1zqCelszII2cCzB0QqFDQpb1IbgXgJz7tBi7XKDWRA
ufLorXi3epbOifwfOSb6U+am48zOyDrKo6CIuLIcrWBKgQ65haOC0F2LKoACiEPi
rzHAYaqE20FpmFAbYHPc1XL0fiwXworMD2mzwRRRIsVC/sCL0p5s5+GkZ55OzOIy
hIKpB/5yksAZXUJI1t3HUY5zd0wP0tolFKwD/dEXowO0LLEtW5iVH1QNcYuUccqA
RC8tF/R+UrXXneKBYMTqJZLwxM3mvSGeShGiMrILMDL4+zSX6XAFyjKfpthMMDFC
XFYOGGcYhlHjz2Y5Y1RTjYduPE8SAVFBn5xlC+ZG7yOpFKEeIgmTn6xqEM1HEI5/
caAaTjMFB64P3Fq02aIWhZYG5yHW1o/F0efHNzoBOrZKcB7rew3InwzG0Hz53cZE
mVVLOjr2MWapro6inCM9ONNdxBuMUfEL9QZ2TXm/Re2PNKreVPlfmyVhxXBkEsL0
YnmDwYiac/eiF+lPLAaOx5AmtQE9ilMIvD1Z7f/PE7Tb6WxI3NVhDLrOZPLvaMWA
mQVaaw9W+gLa/himgbRNN0h3kKZZtQEsLrynUD/QBF5eugbcOtNCHQ7LaBhXQMct
HtmFcKAo7SNe1aFE0Z8W2ZCxwjABQcLgCW2MTjWzAkFYMnWR9TaJLX9YWmSFbwcw
AyF1rxR9J0v9k+XI3IL2rrM6nBC/ylOMTg/oC2cKa7mTS0p/B7UPQ1ufm2abEEho
9oCvFNveoL65OlScARGp9BWieEswdWtaY3jgq3YKb6pXjBYk+Us1uOdDAFPK+DJm
Q8TBK9sLMy7rdvgS8skTBt/Ts2YI3jSibHVRzmzDCVnVb7xq1xdrKnDtlTQ4aWhK
1ft8vYqU6eVBl4eGSDqvuJn3Jm1tvj7kVfWTQRbDOwoxFJe7tGvM3uhkcVstYuXx
JXLzHr3ZFdxhbeCUh2EeX/jPEG/sGYTYhdUsxxw8gEPCjX8qNGViCBKoQMnr2N3q
CWIEOyhKXFMZJZO4ZjA6kDTLAx6jSJmPhSFf7fUKTRIySQ83lL1mGFhm0xi2GKAS
sA+FF7R8ymjm02yxLwstsAEjIvyi2KbilUg3bP6wFd8LeuMjmb7jmVGe3lzvL/8J
GU2On8xYynSx5k/w4XNteqz51q8c8UeYb8cjQfL84gVDJMygm7vplcic66y60xtl
9e/ioYUKIAm7NeryhD6Cjrpapam1bJBL6p9mF3Mq4q3dOVyY/iw6TANciZsKsEUh
iqxr/R+FjBOliSr2py90RmUCUiHiCfCqWSYTgPjLNDnTfo7d+L4ebRx8OA8RITrw
IF0jPMhmcbyO2QdNhWh4W8yY+uuegDE837eToBgWjtusopOoEu/Yfs0AvFskLEFp
+djfn946DDQ7kpSR0xCHXx/lU3SiNi90PP8OQj250+dVAcCbzvHKAHg9oqY9WIUw
YxvKwt3eznQhVkcPTD3rh6cyzMZJ9C6+HfDFJo2aFucSL3xh6ZgPI2vP01NbhADw
0vC/qUjpM03bRA2X9uZ05euX49fZzPaceGiftOF8Y8SxuRKMmVg3GItNrfQZ31Im
yPqFrFfUFMravBjDniApXfciYyrv4Ou/ZpbyKN2lNDJy3g9zOa7xPHdzHnBzrYsW
z1nhILr9V0/p8NqlESXfuD9MZilD5EP1xl977mag1lMXvqOtqHQE6wyWev41oCVT
EhSH+78vFogQp5sdj7eTRRJbvCq92OkpnFNY9B9wwI1MpEP2JK2G6Pt8Y0zVS7YZ
Uxr7dgbEepgA537Y3800lLzXrsnGesWuZxDGpQpABjYmKgDAFaSQhky6W3smL0Tj
VGVUcaQqrmhD3Y/xHXPnTGyhZrTNR+WEbaZKAw/SpWR7ccridZZabF6Bkn1tzceq
Ruzz2v3zshPVDBFhQXUouhgOM0+LAke6+0rT3S+0YOaO0qBb88MGNo9Uc93R2j3i
/vi5pecvPcooFAlQCGfSIeGqFdCTJDEr6QYkRUJ0wBeWp10qi7xBGjAfMxFvZZ9P
VtrqE2hEkZtgr16slGy0J8nkV0HKUGVtzx2Lik+GasqGPuwemwJlLHR87n/Gef/C
wS7y6v6I83okzJ6cBbiFCGTUZOWetdNw6I7imYY3ze3b9hmYgf5xiG2o8Si9SaOr
fMrOKB54Ij11wwFvnMuG4mi31O9xfZczRZ7qVyvgbOqsX4aEh2WEIKeWAxAVtVVG
C1eqFIxYR/p7FpaAG5WoAh/z5L4XaM+x0FyGvTP1wOZRDZY2qJhOhfqxdKVlIk8l
vFkDzUYxMljquWCfQBJwKVJE6R+OIN8YlEP0vzWks8oosUFeXLaL4zurXP6+100p
wOsDyHBdRtLVF78OKUFqligZnKYyKhpM7j2nnOJhmwkg0DAwWGmGkQcA64utNbaV
4PKaDXvpkrdRpo9wvsQ47DwtfKDqdXsoOkrLL7qo3uRiU939AkdQ9b5ngtpOGbFT
YUIiB8/EdsEaTRU6qS/Y4RLKxlg7trAdzFITcZSSfwhjfP34j0/ViXTVMdYxH9sy
Ob5YFc9Ga7LoLRx0L53uTVASSlqfFbW4HY29Zf8de6lNTXeWd1zdDw6i+8gVxwfg
QRlVKqqIo8iA8f3TV1qkpIfuQJOmKqEStMWkbUP79ZI6jzVljpeGSQnXggxVsqRK
bZLVUi2UYL8Cqs+2xLvMsl3UJ9SZJ3ge/DZtEKgFSJrGepRT24EzlSRku9hAdR69
Wqb14my4z+l/8Av2Q5D2O+XBBUQ0Bp6wi4GWFxJzLw3gvsMXyeEjCD8m9NiPumNJ
YKQJ38d6MKiW7WyryKsLp9ATpFFXB+uZqJb81C08O7nLDN9rlDB8LfqW7SSdSpRn
aMK2XcC3w20cTdiNelImYNakGrQHB/Hj5irhmBzLDTo4E62/3YhMSfjjwDxxf/wh
Kq8pHJuIHs3+xAjtqMXLUx9Paz3JVk38nLKi3amY+8TndKrzwG3tqrmOIPPbYIyX
94rTJdtfGyzaaYgcJZNUQp7aA7tUjJID4t6SbTZItQmmfrOsntDtxROnwiKjeMlM
FHE2zRIe0WYi+LxW2fZ5eD0IGIYAOTYIHfslDQWdpyY92w6GjWJgj8lx8H00TJN8
H6EMc93CLbwUvX+LgSdM6zYOKUYQTd4wa+E8fw7Y1B1JvLVYpgLASGs5RK55Q2n1
VccIdXa17ukh0LMpCyuwayr9FZ1vF/3uYV23FuWeKqpKL0oh3vN+BZ9EwEsCOJvH
v8iDHYbg9b74u1xKhYehLnRsxfRYVN8wAAqFpAQMdaxoXuy0u04sTq4t2ATGrv71
9x3rQ5doVkgI3ulrI7YKJnS/gDLtELv628lId/+l0DaoPHlQVs3oStNMvTZO1x/8
flKh9YNMgx3Z1J2bM8huGonWAYM/ptX41fT+ntqKOd2d1AY/xQHAtNPZJPhyIse3
m2kAEB26oYbqbg4RUa4T06rGxye/D7L7E7zxCyJqdcMDiipYtKi1XqjnQrEHY1mH
3U0OMu57NVR0FpaR3EtYX1okRa88BebOxnZSUOqFAvZK/jyvxlZJsNJml+IZhyaV
pmeiF3qce0XOGmjDfL182CCKg+Oepibq6sZJRKCGAIFiFMCC1iY/1jrWLbSMqJOM
loWojp/QVV9gSwb90LFEPmIrHkyPKvKUcLTMhXSha/ast7JVVSUnkQgMsGPPIsnk
dz9wc7iEqNIH1aEmGyCw7O/1yhh04g0K6wRzVwsSws0/IZFo+gfA1Q8OLigR/5fY
i7Bv6URFJd0i4IlVxcEJ/iqntVpTzEH/XEsLVCsVCSRvYnsGTUPHLjvXDltKI6br
RdBUO4NaJzXSUXbp2qqpR6zb0DSTGVUcXuc1e0RriFaEm1Huf0UtcZnsE8bIKCPj
uCOztVshDYgP+ixwuOe0DtC1IaKon07DAhrUMoY1qN7S7ZtHyPEnTRNT5qCOHse4
Jcu7QQXZPZKSjafTcBJniRCLfNQECfQQKARFPj36fX4+vQx/EG6+KRFfB+/hOXVg
WvUkaMceyJJwZAqAexGwRSHWSN4tZS/Wbp3Mp8C9ExedF46sJ8GBd6AWVj6uBjee
pVs8312YZYR1jZlZdudR17+6wwIl3y5ZJCAqM4To5gQKKhTowURclXkSKtJ90osJ
YJ4Iz3t0jyU7Lty9JtlOPrQf/NQXpHC1lHH05k+LTcdJvVbk8vSgw0/1ARVoku0d
l1nTjIEa/M5GLx4SEEOChw==
`protect END_PROTECTED
