`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
anPJbnUncAZy9qshdUU6IBpL0cExRlalw92eL/+z/qFHmYIKKK5WfFIWuvc8RJYx
+Q8Qow71CvehCDTg+GbfDV1/WxykoaYzRIYNHCLjZOgB76rUUUyG017HK6UdoC/V
oM8tvlE1VlOYYUmQMJZyd5nSScWnNSJcuk67zlmGUVQalLvK/ZIXadGKO7VNezqK
j+7VDsIaCaiOlHaNbXFLRc7qjnl3rryNwDAzWFYQtB/rBvF+LS1thkLCsFK5e7BF
4d/q2BdynhapUFN+YaXSHtYjLuJ3W89hnXTdOhW5tLUzADNT8kfKKehUIUApoQpG
xeNBIUkY2kSWOhAkLYW5Xiz9XM319OrdQdg2o73hVMi9MCb/qmaZBliQ4zc3SnVR
V3L1P+SogplD2/ZcRGoPeAS37g5yvmkbvCNMkmg0FeVz/rcfgdWyXCD7LTycD+t+
p9tI5TBeuuWLbX8oK3EdLtthJ6fHVmmg/EBiVDT4mRQI2WFvvHKr7TkRaULgxhGM
HuPL80Xc9orbBtmf04EVM1JXWl40qsEnQKTMkq0lUhh8WcreH97yYxI8t+Q5sc0Q
`protect END_PROTECTED
