`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3OTJQLMTcmAAZVAx6K2eduI9FmD/1s5Ej9VymNyCIn8UEfRI2/hLOllSCDOS7PKk
w91lD5R4aLYn9OXf53p0IlJzH2T0GQMojKI3o7S4Gl+gHY2WlWGj2cIyXb+/Q6yR
Ekt/Eg7VKy/tTvtLt+bJuMk2YCG5glWV2N43BzE3FP/otOPaUhO3WjonTMoH/B+9
3MdHJ7Ph8l19eiK2oSLr12QHHKAvjOU4J5e7PGe93KD14E7mOwUvabE2theCMjrh
DQJAU206RbF//S8M9Q+IAErRi0hE023uXCqpz5fh1ApgZbol8DWXZ96sIbzMmA7G
IIWo9o1LJ7LTe+2namIwg0DwC72pNZ2b/lryU/scKVxgdUZTV7XcXoyulxqN8NS1
UUS/i/b/oYYHJPjSFciOreDLHTe8gMoyajgkCRMh5oFmPYGM5BOuveS2H3p/se6g
Dqoh+/cuWj3mMWqwKc1/Ahv/2JXt1ozVrqlmk19RDCEhpFIaSSl6irveM4qdSfAT
g9WlOXD+TxCX7c9FmvUx/TREOJsdaPu1s/lENXn0b+RJc11uwkLUGnO3A1DTnoe8
EBGiLHPtXH9pwCuxHiowWi9Yy+ym+KGrILMXTla+jI74qv+R6BgX2RNK+M0rym2q
KnxJumCl1fkATpGtsdB08Aw8jNrCRycsI8Q2Hthw9++KV63y+Z6gSG2m8gbiVR58
ZK2ZHWDZ1dL+cv/PKW11z3e+Vd0T3C29WDdMLNlf9TzZXQKMmazlmgvFQRlqfF8q
iNsyTUnzaJX25KylaxwwTcPYdiKRoxpuuLe3klNCMA2u7Mn/HhVw7jKCKuCoEY4I
/jNUmnAukaECkpaoOciuNl9+EghBIfHm1/oawAcRQQsX3RPVXD+dW2q1VaC6C5AQ
aEKg3pnZaiEk8QriaHqF7lcA/xMcTQSgerZoanXQdNRsDNGb9Lis6WscT8IgsPU4
5LYBZCJzpAkC9BiCLt2SZiVMcJhqwVRDwYzKbI/82DxgoisADsKxCTfUWbnijDVL
DU5ITEZ/yrh8FVPBYvQAHVQrF0lrkYf4hdSdlnMzzjaInYS1pTvQPubtQKvyqmHj
S2aRb1HUSJY+EKIJxAetkxJAXA+1N3QIaP6TUqWtDhquOOxD20Bo+2/h0NtWB40Q
thsSSZsV1fgdiBzxStn5sdO/IKhg07ZSAFEZ3Zjk0X+c6TP/41WZ0rI3FmaKlI56
MbXokzDhRE/CUYw7fAuUg7Jf3vAHoprL/qqilI4zgpNNIiDIwcJ8ek/nBJQGRwH9
8psp+vCL1ZOyImVLc/Acy2cy1MJuksVp9sORFvuy4b/f8hgqSBaxRK+Ku1AugLeb
dfJQnUIeRrsSjo+N9Kc7rP+A0SrWHOqINindpQd4RKMOJS6cS+qaC3ESXc943mfI
oxM+ZjLGNgRmS7Am+KRvdykV+sUtI7r1cgPPqEBKrL/TqZw8bUcvX2weCeHdawsh
MM98UHNheEa6zJ85XFj52P1Qy2Vh7WEuzBcGH8bINUo4q/iytJF+5rCwpWC7uOoq
r8wzZDnOUbgE3+HFM7CfdFAt+3Oi90/ZKf+lUpKUaqgNjVqDCbHJ/LV/4mOmbcp0
IGyhgjEwkxeI6dwrzKrGVZCvI2EeRWD7PYqk3pjw1nhjLSusKu3n0T3PTmvtdEjh
GmoMX38eI5foMb2U5/1K2QWAO33F7NP07V6f/JtnMwVzMvsGnqr++pS6GiwTaFHC
S7rJ2EE3LTg1cpzt2rBpysra/us1sYuvv8jINIS8emqBez9svA1gsVwUpsx/FAlQ
24Cu3DL9F5wLKJeBjFAcSeXe1g5/x6iu6baHQIaDEDc5bQqtEGhRy5FdqPdGeJbd
GSJDoH+MHVSAsu1VS45g8XOO+fwt4We0cuaga0nLzD9cCeP79u+ctkiMv+iy/E7/
+lFRMirNoStLndK7IPCvCw==
`protect END_PROTECTED
