`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNwWbh+4iiyjWz4jOj/VNIc9kB/LjSa7Vo4J3mmaFzFWqznjEAmyrhmkMCArjN+U
7ZhWx66IrD/B/ZFCCLJSqRYR2UrEqYkCYPAUVvZrPGRRhy1+mkF+mPhRuL7RAXVI
MCIiNtCIQ5dV/IwHTUwdCgYOzMS1qrnf8hM6k8i6r+rTKwo8F5ooxnH2cC8HFFly
2MznyXUwiZ+dIjqWZ2dcJnCvI1IxibeyN3bvGSnYsXRWXiulL6O9DY3j4+HDs5jN
Nrq5vdPU3qtFDWplV7wABURw2tQNdoQ5RlUBzYcM5iluhPTaDyyoHDrMMV9Dvps3
UHla6KCmg8Ld5PKW/g/PecyVO8WDW26U4pe4WNH3sQuieuoHych2fwyczHNp8+6r
TDtAjdMmMiIBjokxSkOSDwDt9VeBrSM/LhGFn68oAriF0kIUVaoOMrKw+qL1d8QD
uvdx3yT/Ae/dcP+P/4yBHg==
`protect END_PROTECTED
