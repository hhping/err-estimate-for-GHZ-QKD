`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqDDF+H0W4n8HFyELst3lP0/ss3pv8MnCYNSZS3U+V8u57zIvBc6Ub1Bp00yINcN
O2jJq1UBXHUll4ncvY7Bij3v+0dgj6SfFsKhpB2vGammXA6df6ONSM4dsLGU8l2n
qlZCnmlNzeqsED0BrPfEOZP4j7i6mjo6siennWTRwnvjFrIO63qmDQ8N9Se88sYa
YzSp8lgxCwZo4cZKcvkM6esA6RQHiAmgcaSq0PCqndkW6i3l6Dritvbz+4etQxIc
Inm92HkFimhAG/N/i2YIZD260319iUmJbpxOe/3kXTNfo85f6BUUbqzg9pbnrSNN
4HsCXb1PZnVkFdUPD8sbAxXp6Z867tpg4bqfHByCXSxwR0dvFJ6S24HibDIKDGE7
w9WJlyl0V/8YyTuXlzmdo9ZsAm8mjKh+nQDaKr6C5uPV3rXxc1m127gbWYaDsxgW
2ZhBieC5BLNvpjUHC4J9Jdnq4kWY7riGz/vkcKNDMmMYHnymPKxVcMj1FqaRZfkL
PAJmIWdKpn6BRTFHUaj/pZ3bci8/rd5VxX4dCMEqYyOUdnVScDxgtDPSjY5ad2yf
E20MG/xa1TQlZjHTRLLuoMmGK2pAvOt8T+rjPTkyk0+EhobSlU7PHzMgHZhNM8yc
GykghUy94767ucQlOgkhyWcEztUwHOi56VOpXJoONf6l8R78weA0uFMufE0ZeD/R
KFc6c0JoqnTdDP3riLIYIEkvBmrIL0eN9MZo5cbYx8Oj6Ut93+u2EWNhUftQGhoB
oP4SD6kb2jK7wsrIQ+wgCRI/hxZ//piDE3stOhOi5PTNJSxEx7tLIbzXKJpjjiTD
2v0be2kY3KtctmhBzOZ9BOAASz4TIRCsKj6dqQ+ogPuYbJF9M79MXanQHXcEjMEL
aTuW3o6NJFtxO/m9Uax3DefbCEIR+wPQjSH4nTz7ecQC0n0qA56++xmy5+R41Px9
4SK7wRc97X0l/chg1ai6sQYZvPK4xBvDHXvgZzwYIW7/WkLNcuedLjz/M+NiyZf4
ydH4Zz9tUpNcUDDHmuarBiC8k1L6YWfk2O9wviTZ4acyyW2wG5jFzSsjL3G90lbA
GHSFFsNjsPIDbJH2K+e7YsCazPAq5RzG9ootVVceDfsSf/mTI6Un6o4KIZ4uc6Ty
Qo7/GZ44rmvHnpO+Uc67dlfL+AQ2Yd3ct4jyT8GBWS1pW8MB4V6WiA+nc63tuH5g
YV3cKcbn1V7jwkrky07Ji3pGzb53+j7Ac4NCK3oaiS7/zAYyylqlZidtCUfbNBr8
tAG1r5S9LKi1OGHkpBhOJzbetU9dQzeLz4dHzHdlIdNNV0XHeVzlrFp8dPcjWz91
LAr6jONjbT939IsQ5Vje7j80hY0RIJAkCPsG6VopcSDo48zrXV/wVpXp75bI29q7
3u6JKaE1VTGpfOYsPwwHiw4D1lOo1MYBpzNu1N+D5AS5IwZkdObg7x6ABK5NFYaO
gi79a77xpbJUPgwFpBOt1g==
`protect END_PROTECTED
