`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cwCiDMa8QTBKERNbN9Gv7VqhjitAguEn3CRvZIfsnnRtvWyZepZbRZ9n3SH+wiK2
9NZwjyFSFI3g9yVIVXh8+rY0C9X034057oavmGUigYMCQuz8Ajuvml/ljqsJu1ZW
0I15Nuua0+Us+ZaSL5aVAFbtFELeoPf3F27A/cXwQbXPDHiSpSW22TTwKBsJTObx
1YAGhDPe/Dz1cYN3QPWOdeDu4vOWDtFVuuncFM3ExI5/5Hd/JcOjtxL2fUBTXiRd
CWMvDft7xQX1r9qvXkY9ll8bVVW6GdNrEfIwy8Jpdq/cmugiXmijXwSrHA/r8biC
2LZEFMBtt7UbWAThycz+S1bXa6FOyLUIQIk6ULjyH7xKmVCUUrPhmnZ4u1qfCEjS
MXvVLdZ1EONEWozfegli2lqsl3RUCwyKdMkJJqtgj/kSznNgRIckwbYiwIgwlamx
0c2rnk3LyC30V6fJyNpPymovnrPk0f+ihkPBX3WHt5MUgvB6t6pQMy6ynvZkHEG7
ndWorbmjCrLCPnh/V3rKvnhjSVKfEfBTb7WgBS3rmUBB9B8e5YeqXtVeZQnVWrIR
8GugpDa5q9Q4+cofXE+UY+AoRm/UKPWXv09Agls9UmTqw5b/j3hXx7sRkrkjDLQM
jYhhASo38WJgaB0B7eCWyP/6wLseTw1w4fZjMvW+Uqlp1Sxrwj0xG6HYGicSq+CZ
Svf864KiIkvvqqwa+lfsUiR8SolVl7v968o/NC6jtjRXNDwHzS7rwzvj1QjTzahf
ppxjws7yAwi04FbbmVn+xHrsPlxqQ9d/06t1ALQis19zv+neH13iaginTXxCpjmR
J67nIY6F/9G1889nC9ziRanl3FAvwnuoe7M++WJeOd1FCUlRpOrsCdCf02AsqJzU
h2OKqh0etUirlFCzrc9rSxE3lpRgMrJvK+PPzpNsAOthkDATlIMqjWl9aOCJOHr5
Plpi01aihp7zqYxIsWcAgS96yJfFGj/sY4ZIbaHN69Rb75WvZiutnXhfwRkTNY2x
fMfRS9XRT1KeQsyPxyVMgngvevp8t2NBYak4hhwuAg5Hg4vfccnxgc6r2LSzppUS
NjKK39lKe5NCyHvd7cyQDb8y9QfLIvd36GQfjmD0pLt0MhJ7anlj2izYIBhSK3st
4ZaHWA6A0Li/R4OYDc03hlKayYRgqNQDDoEgaA5O/pK0J2YW8j2XloDtlqP27uAy
Stp1vVg829H3UeHzZM91Qbsi+hbkLnwFYuPVpXPI3ijvBAU8ip/gBNuYkD1Ufj34
QDuyLCB6wv9g+Ya/TrFCJNa3cz3QXvXCmX3NTF5M6v+Gjl5qalQL2yapYl9J0mES
HAbRg++7a9Fl+ZgKKZrT4U1soPsRD9gMVG+BCiCPB7brG4kjlMJ97Zc65M9xlMLV
eNS0QmUKjWUWcp+YOTWHwY/ESW8b+q1uU/ASh6IDvuSwxklwLnmibVzXka+yW/dv
be+zf8APiZAzm+lFcpxD8s4VYK3v0jrcxGULZabAJDTVNtEevmbdh/AFUh9RknbS
2fOzyYkhTzlmxixTPNU0TCj3396gzLgOE96nU2zD9FBVLEE/sQYUrkifTkuwiPCH
b0HxLazrbD7Spi6NUP+Dt3osY1niqCu7fRSg+2MXghNoh5TfBbl3iHL7lfKOi3Rd
3CKA6Nb6k0gMZ1nTGdXT00VWq42BBRKYFDTRPQ4XyNvjlJXnbzrPtetMBd75fUlZ
AcTgkddLbWMDkYCZGDdlEwnXDGogNcfFhWuiYlrobC17oWSRPS4kpiaS7ElgO+7y
vcu7xn5M92NRIkF5dxsMTHOt7SRhsnT/pI15PRmqqN7Bv0/oy+fJA1bCy3Z41jy3
ChdfnGf7x/29qhfDCZ7EFGXC4PuHeL0eV7hgRy9liNN8tgJM++244kOekdP3uGik
nFmE2ncTJWCgDgs/+RQo5kbr7mqMmiUUagBcUJWT7yiPDm91nu6igIN4S55OUGsI
UvkK0pEalKvslNmuOWknPZg/zi9v8FzTDm5ZWIW7RVgw2OfeRCwmg+i0AhoytyJe
tmBGOEZ62crLI0ssOMSywnPqNZhLURXNSKJj0pFwtyUCkGLSVhjePz50zasLGo0J
KCv8UueFAcPUQKkjlesIfkWtCzJZLHJjOMr018HL20zYoAYGfeW3cH20QCOk1KgH
OFRS1IumWLBSvCy/QyK0McAjKr9YLnOsHYB+qpuIVsuRhcVZl6TULAUjKYZbtxqS
m06PBDm5LBh7DQpcURn8NRog9LjOQrVM3K42LC0Vn0mc1fS0ARVtHeUm/5zq7T2W
9ErJspyUi4dA+G3RcuB1Bixd/UectazFTiyCGNVc1O5F1w15LyvaWCS4sFuLrCd7
7Yi5oOk4tj2bAVuC1/URyaHvrb3nmC3fg6+10EU+RSSmlWdSn2jKSuQONexpzy17
Qt9sw2VrcIDfS5gHoFpJdR7QUKwCcQgFBf3v+AABfwT9GEesiNnxbJ1p8fP4VmLE
y3Y8UaSd14Ts+PXkCBvVE5Q7lIZyXvU8Xpbv8p+fb14g5PtYYssAjtlA6kAlEGCw
USaZLXBVJwyMMJiop4XDgIdHs0yU8l0b+o43kiXbq0WA63WS4tWP/MrLJgGpOEqo
QZAq28Mm5Ygt1Ez7ro3C7cUHP7nmE30B1KGhkhgua9d7wbseAIbOsJ2FxjneBpUr
eompDk/8c9CQsB+cuIZTS5GLE4jJ2jS7McPLDSCJw4i6IrxrwT6SohS+f+N3vepx
UYSSk0Ae5opyoEmd7bPFV0XeQ4WmTKgSM4YrUbA/g27Ne758MBEk+bQ/96A1n6pQ
h7r0qgUEii7nCgHaGMRcRjj9/HlwUmReVBmqMaMEHxmkr2cUccyuJjMr/fA4eBdv
/oFC2i8kS71uDeOGgH7yvv4ZWg/BQBD97yjWKnwO8dCkor5mk+JsXt5Ld/oKx5Rs
R0Yd2RPTdH1yxwLpD3F2kaHF1jS53ScBMEKZMgUHcy7sveKkvT6zwakp64aW8jPE
htqDHQ0LJb0n7Jo/1PHi4o/040EGAft3Us2slefinoia2kQTr7U8id8xV1piSkyH
KByCjyPMvNO8nzDJHaofuV72YOyxN3IaHHj92yfKvzctDI26/r0Vo3GiYVnxfWh5
KnpC9bOTAxdMkFGR7eeqT3OoZlHrHIAq+g4pjAh8nVsWAOVKwVyJowkRQrYJW1qt
bXP2/VGNdafPi3GaTS7LbS50OX/R64084SowFXA32BhKfnMvp99FxcluoZb7SmHk
K8trVsc03yOAy2fxG0a2VZ76zYMDRF2jvRJkn7Yscas=
`protect END_PROTECTED
