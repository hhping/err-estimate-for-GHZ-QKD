`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nl5MHkzB0VBPylePb1YIcor/Pb81/6QDVnXe07BG8Mu539kSWdiuZcYGjOSjYwUg
kkkzCPtcLZcL3SlPRYQLbELPijNBx06W/2ZRNZjAvcjpGRA+Po8eo0MEbkEwM3M9
Cwp91QvVabWu4z/MpPt/wLxk5wtc8dftLB8tqpHrRJ/wh2zYa/DFzA1tSj9eWese
brAoYQ5XGVfEmwOPyiBk2hfCzmot5gHiZdXiVM+DhYE6U8YA/fDooJZy5PQ8Xouw
1tCLR5o+fuEx5QxsFAn3PueYHKfVvCNYUtjHBFhrWcuH/DaRvjfK9PgFCDNCGYb5
lnL/WJMdcYUw2jO0N0RAmmwtNY+rFpScFohqBErxqha+WlUt5KXjWOz8LUGRNmjV
B05+Xnfomj2SwGjR5arenk3H7aN47tPkLp850pvEQ5zRMMClgnCyxiw0X6LXJhPH
QtU/wZHd8wrDkLbbMRNI+7AmjiJutSzUvKgitNtekcwvCsWSs7EFRXDUCqb8Kyqm
z+kBlsNJQ44YT3+uf64GfEyX8JuUlGje41ErLYhg7syIoDDjla7PqYX32hzkJe9/
dJM6YWQ10wzb7P76CQZayXPiRYiE/WDZ/tkgazoO0sqzmpY6xi5VSr62RISuTOFO
QacH/FMAeQw/lONk7gHprFUKF9aRVayhgYX1DW8RUUaHwSFiMxlSqPHoHcQ4vB4o
ItF9W1Rov71CT1pdMP8VHOVnoOJG/jgYvUkrJR2xDXUyKAx42sHyeP43motDO7mj
EZ/f5as1tSt6gFLBlieF25J06B9S0XSBfarfCfjPS4Wdo6IU7cQQpOKSwEuR+nxQ
qkrPh/g7ORg0/pReq4x8VQrhkuvqYYYTJqlRt9VBVyHDMd0ZtSl8dJ5QhgbFMtag
qr4YXZdGPNRT8I/WxerVzLTRq6xnPRcwteqQ/mvhZwVWzLWMrqNIvHMdHlg/VfiC
aRujZawHiNo02iXhVHItnEM/yK9J81RuT+Fdc/06qaCBUWPxVq6EU1HfvWIlH66D
w2Lv+Q73oFmSWJrvo1HLx1uUO4+Rv518jJ+enN32eenGfOljEUT9ljytDc+kPyEv
emoPC1PraybXydABrAevFtL/CkzgJ0dj4YI7I6mSpeBf5ztQ3Gtf+ISiFd+Uiekh
kmHbqQh3h3eGs883Nb6UO+m1UtsRtlI+NX7U6qaOos7Fx6DN8qOXDNgpX31AvfB1
`protect END_PROTECTED
