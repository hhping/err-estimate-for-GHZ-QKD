`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3KR94dlQJslz7vQng4600QTSVVVrx/a2miOV6hFVbi/49cUW0BiDzXx7HfidX4u
mV1USmeyAJBFUVrLPSsJDIrcAAk2KPi7wFDt5v+S67a48DpiLk+TPpN/jO9dbdy2
+rmzfc/0XU9RLbv7ip5fTxNVgZOyXP+RhSLXIOgZ4cQm0kZPYlaVCZWH0iVTBYFI
/Li0LUVQ2Uc4VX+tIaSSTdJGoSml/BNrSV5LF1gVhLIHiNr0+UH+FQwW3qkfTx8D
w4MklTlbgbWYnMjX7ON8RZCAyeStn7oIAPofN9wgTr/rZOtOM280LcdaS+HktPAS
nZghjqU+S18hywkas7TIYpXTPeLb3udaho+ZUrOoSY2e0He5+/zJI0dIjxqMsnIO
Lr4Ot/oe5dWrOPkxsb2wZb+8NJAEMOEXGIX4ebHBmaUtzCZTc2uLAWUHDNYuvfC7
v18DWxpBOC8Hk47Ntw2+/r+DxkOy/dPiosQo3vJNhH1favv7YamiJHd1DURe9gFn
UAainMQiGPpoUZejgM8BUOIhyAlr4azpaQCj3KDmwYL+Cc97Usfs90E1UsZg4bpq
0sBQ17MifWpDMfl86rsq4rRI/TJGbRecYT7zr5JeW5dr4J96Wy2ZVMWgkVp2Huxu
UwEtMxBiiGs3nw3pqNuDXgzfKO5IBkQsNcXgIKiiPtdp7ILDrD1eACtqgeCmuzBQ
yN9Ybh43a36CmELULJSZ/fVCdCVyckwDJ59mXaXqCFnfrgdC5kf4jFHpMvU3ytIZ
CaFqD7IlBY12sdwSD7rL9lh9QYr5ep6Xy/1OqHceMVOwh/W7ApWQ1fxmQ0AFxBbn
x51X53XRO3MWeW/o0f4qvS44sqs3x9BcqjJyiKj23gkPc+L6XQvE1Nof9NuS+qes
Mn55v5zGA/IL7dd46PHmUA+Ir8zl+RWi6UXxXZUedCxNLrLBHcPIoxB8hur3GLm1
4xqyxPG5mNM/t55dHETebUij+3C7Ji2KreusRM8i6LDS2BeaAH6jdjd2UPUZtt99
sZHG2QSm6/T2P4u/Yl0vRsg1TSLIkeFhkkapsntPXv8louYuzdygEu8eR3f2HF7Z
gE4lT6zqQEti/uxzT7LOXiLvOa7OBtUGmQXi/dN+XmPCQpJKvevZi3vcHwTPqR84
RKhGNhMMkdv3QHNlQtINoh2k3rtzuu9f3zZXWLBF75wrbVynsrlvqyPBBYEhsVtT
bnPxwNCyzUUBMR3EuDwYirihZMhzqG2AakymNNBFzQKVjxVN/7AmiKaffMYZHdUN
M4OOSQ42dRTSriAvgrlBOd5dwXzfb1FqDQU/lfSvheZCzRLLwG/bbtEgQk8KWb9t
Hoa9+8BielGX7AZZfmxujiV/B99dPJWtoPdw7hNpu2OwKnkrxV+ckU7Rm69dIeON
v+dfJWd6Pj7RRo0XsO35osF/KaZPCLeIDeFyxW2V5pB9TyXvMOJ3m6mzTZv6HAI6
8v94bqsiYH5i/2D4q6MiLnaEkfLpgVJmfhfjmtL8kJVp2GrH1rrCpInQYckzjEmu
p1C0mRU4pe7KKTDw2CJ8euP105kHtdthdPvMb1W9z2Y+VJ35Y3ecTuq4wGf/Nj5o
Uk9+/ihaN4ORApgt4+jDP8DX+YUk3JZBdnWAEpFWsNzZlfM+Eh6f/PxHdAhU2iOC
lwlhWU2jP9UJYEcjLIW9E2pAu8ktKsrCuMX57T9vwj2vVR/UbZQr7wMXkMjIFoV4
zLVbQVIEgw7gmAHiKNludvXHUS0hotD1PoTg88hHgg+WUAf64fY00FqJu+HSl/PP
Alqz5CDUdhwVwijcrp0wySCsDDG6jD5MrYr7iH5cA/IjtGctEb2S4pYCPFcDxeXu
/sR3taoj0YKyfxFuwaxtzeF5ORRp1JHHLJcq8pzDreiSMjwS5KmD/Z2dDzuH/JB2
IvhC+15Hct20wMM0I05ANe8dlGzbXZgVc5rE0mQXItMAvauWQrjShhfznm9et6Qs
u16MZgV4VFgERbaNJ0kSP/VIOOae7YvLU99aGtf6cz8+UEMmeT4Fxc0JioyQFxtH
1LII5zSg03A53jfweeoU31RyQcan7PeO4ssIBY5BCHdf8OLEwu/2LYA7yoZtJ9YT
fXdehNwBwtiljvm0nm5fJz6RCEPyuvfGBR2x1Eqgu7BcBo3MaLCLpOCnmMsGjs62
7Z79Ry1v6h/UOWhGbjJcgj9Q9OA9yGYt5Mcps/TfFQ+FeObG1hV3AjeuvPABBXy9
UG9ipbfbAPfqzwPMwU+FhLo+pw2sBJtEHaYFEhClS+nOH62bxOnQdbShECjtEERW
i99m4O9oFaoStTc+q/pbScYiVWFSITI2XK/0qJaKHg+7LZ4AZx/q5s5Q/Ujdaq5M
lAKAZ6ZfatgYuERbsrX4AGWx82vVHrx5KALhnCKDU1LWpIJf8Wqu9rerV1tjsExc
RYRkKKKBwc9/V+Cb+ddEAF3WXDSqoQwmtlzHNYwImCOVZsOaghmVTzfCzRqaH1PZ
Au02LWHs0Mrf4PjN8UADv56njel2RXoj48LjgoTl85U=
`protect END_PROTECTED
