`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BBbFSvonc/FSeBPtEk22IS2RoooHGW8vZSzFhXlXg/DvSHjQOOUGdATQe4oA94dH
hqQQIxBb/tHdL9h5MPaIPffcNGaDnzM49zaXfAiMNlivjKK+Gkywg72yt3c9umWx
Xdm4FgO/U3fWzstxepkuPtqTrOZhNB0EcdNcreVnqZlCQC0Ty9imuvtvtHtVADXc
TX4KgY3SgYEI+Fn39EmePyyxE+ZeaMcsf1HwOxrjujYQfbgVvg20144/ubCvQ8Pt
cj1L0VE/2nsYh0MJXKYiIYl8+1MC6bkMXBswl8FJ3Qoox0Az5PNNv8DAJeBWq5XS
zyHqbHGhin91WWIBuNMjg/tyOjnkx6Bsk01IzlELpyFcDTAUQJRA+gv8gX+3PruL
ChjbLVx65jKYI7Rn5g7Vo4q0dcTRPp+XqLHccSnwx714PEHfZTvPigm6x2qqP+YP
xDVZkrQMh6sTFc0UY70WCprfp0qugvK6BR6e55YQ9IZO7ePD4DcTz+3CpfoT1fEJ
cwN8wF91hKgPbdjghJRxFrp2VbdWH+twC8KlCQnh6xk=
`protect END_PROTECTED
