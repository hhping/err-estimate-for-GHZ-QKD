`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VaTXMB0eLtDhJQPaFpGM9MNg/x4kUHvQuh2U7loIkjkNJxiE0iYaAIaVxOcDoLQP
UsqAbk/5+8vdlHH9OuI1Vy6hbm521kHnpBD8S7O/IugRX+ZAZqyMoo4hs9oWgxxn
bZpBQA/PXSxnsM6nTlUBvcVtsKTpnHMsNjHd32c71r2/X8O/n72x4YrF65bDwo2u
fzaOp0g4PRL6VLUjBb8XM87CEpzoyAnviTHqLwVSB1pXmaJYCMy8/FkEHdmx/NsL
5xPx4L6GLyirS3KCJuo7cVxexJJaU6tepGAJLi8dr3RVPf9odJOEQDNhGng616FN
z59wWkEuiRugtrImEQxabaDuQ2AiOBp3u+bzI5JV7B4rGswE1yCK1DA9E4Vvifsb
ZQgxcDtzJTiZPc/p1c9aHB9q7aEjdtKr5GKQS4sGnXcQaZr8nNEuNwKTDCxiFCQN
a2GmKsrazGKSDcnvzy/LCwW9s482TPqW0duB4Fb/WjAef8kbXH/yIgBP55Vuwbch
wNV2bKtY9+QKbc+XkP9jniqfP4rI+N1HvcnFL0NwvZ848S/LPzzuiNhY5qkVMaAv
bOfl3mL7VhjbalwuY0uk088OVjHu6YzH6kfx06AiN6TAbS7VBlm83BXiHUMn9MCY
TxMxdSToalFP68EGzxHEWRj8LcQ6ye5qyBzvg/PYbbCZAlAy6F2m3dneCdvQveyI
m+zQmMjIMOpSjo++0u4as3NVIyGYZiPUwWg+NkF2Va5m02lkE0lw/MCJqzZmT4D7
bgFqmsG5uPpidxuOkTwv368jDcwZE2TYKe4Ugfab4elxdYTNXGvcXyEInTO+VU5E
UWQDML5SG46WvPz20foL1xCShaXELG759R1r2VLkepxZgBF58M03qQs8y+qYEXbs
mD8mAHZgwepWcw5Oiw7Yfxzz3srLNRrwgdVL9FYoJQKatyhG365tHh53umWsZgw/
5YVvbVrGEwdIzVNl5vqAjOOIdNPBex7MUyiuVfyxEHwl5O2/JcNxh/5RR/IVZAdD
Cl/GyPg75cqHwXwV2wgSbkAhM3Zz4VE8ZHERTaGxbh7zz6rdyGIRpJKvXZW7qDxd
DE9WCoLuLV5c/zMEaZq8SKkP1J6d/p8gXk7kmHgqdhwEo70NKU+zITuCMuPvbpjI
Unip/WjtWvH98REcq3N38mH2eUCHlabuCWtTreM2+1vSkkaqM8E8DiIxXunBLBvn
YUYwT140wKgMcwHGRo41/RZlzA2ffoMFDHXmy4P47Ydw9bYHyj+fZrJKSYDjsSls
8591qQ5iwgfm3KrHLIsMILmcnQ/gnK7GF4p42sJUrjmWBGKsWAyzO8VTLc6xC+24
iVQubTzgkS1h6RsAK2xxQBRnv67C2MjjzVV8NL3Q380j8Gwan2QMynjHr57mN4ID
dbqAMOboXrMfd/CZ2Z2tgUxCsMxGfoLbxX2Amxsq53E4LxlRFOtRZ42o+WWYAxF3
jQdRrhUiqKRLUa6kTxlrWw==
`protect END_PROTECTED
