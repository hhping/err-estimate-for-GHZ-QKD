`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgZkYGsqu9G9UGw7xqrO1+DA+LRYzXTKhxItEU9IomGY/wjL9z55NBg/eb3nHi06
gvTIJe377MyW0fXfOs1Q6mX0cc6lgkZcPzKpx19xbJkqHRCM//D45HLzihWHIj+v
OyDGVxHie1LsYOtKt/gg1lC5gkgGAXzdW8v4sw5xdTGvnG38V0bKvL9m3r9jXWNW
Yhz7Y18abn4d7BGEy9Dw15PxY+AObnQmVNW9VybuqHjvSlcZUVV9b0xgzQRDstY7
lSgfb+FhnYgKTtgY3xDv30asQXicvpZjrM45Ja5Yawrr3nPFNTN9WQVOmu5IDpgt
5vAqlrBSqMUNYcL9cVJNWZYeh8zibPUHTKlQHSjHI/S9KrGCXh1peWO+bES6PzDN
OwnrUAocg/j65LIydjouh81xdHeU6DMh287Fqy1mc1U=
`protect END_PROTECTED
