`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/qbkk5EF36CHdb7zFqwFd4ZWQclVC8daVhO6s56Cfncdgyerp8+NA6Y/HDGNHYG
ZY/MwsuDi2s1tqulVDSL+NGhuXd0Fbhmr5kYaBmhBtzHpqDQkR+HcOvutoFaFL0d
EOVE247yZALxk4c+UgyFhCZBDrzh103FqYsTj6lC2pN+uwTfRSGQG5hT82mHAp1o
9Qk+LZkr9tF69ay2s1f5SfMZahcu7cPyrII3KtQartF9xNCe1AR7vqRIkvs9cu/9
/DpdTkgoecq8H3mLCynDyIOoMowga2JtGc3QFkYLLx8VvogC8bH1Zxr4QMqwpE8E
Hs3vDKc+Ho2PDEziSO6BQL9EVxXd4/VCGK3g5ftXWu7/0S3AogXDvRhmEKkQ0GR+
FiIis5PiAmJxM41YBHJGTaUZLKoJfAm6kyqXb4oERnY3hjjAAgi3CZzLchFUGyrS
cKcHKrKvLffxhG/BPghE7T1CaOmcyceulFRNXFkk9l+6oE0nbpl5HP9ir7jEdPcy
EmVNgi84dK2MPBxytUjw4RpgCR3c6zT1GOaPpnyVD2rON3Su4UgrqrzwWceANR07
qUhj//ap8oTV44lIo73FRAr6tYDFDQdJa+/l321NXIee3pMLhyq8gZLGM+sQEmVt
cjyPzFPwevQi7P/BZQZ46O3E6QurLiZoVBvHMxcvtkNAnIuPC/7j/RNwAXNWoLhZ
UxBejPSDSHbh3tF8mu83UdWkXPVGjexQzx1kgvFQgDpOvtGm6cM09/GhGMlu/Lp+
Rlpcexg6mKXkoLNq+liajIf5+trJ9zrdkJc/2bvcJUwNIDcZolS3KnyMSI9eiYmv
A0fz6L/5nTTUEF2v9nOeMD499kbw2IJDPl2d5xZDCk6DhBuoa6zydhI2N7c49dm3
YlhY8oZUXhTHVxx05Q3bL1oTSlEqGjrxGS1D+tIrLj7AO6lWvlzxQbfr0tJ+m//8
Hj6mN8KOjAzYd+II7kWw9LkJy27jyrRvGPNeI3K0jRBH/YDciYWm7X7SV/MCjicf
XbLwgQbPBwBfl65BmvFhfb6Aeh26EoUUKxLidgQz9V8=
`protect END_PROTECTED
