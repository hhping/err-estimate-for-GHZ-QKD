`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fnwJKzvx6I4PmJrTZLeaJGAoa80CcZ6Bw19lA0QJbWDq/v4m1OOe2DFJH0Wl6Rm
jTxB79pK9FkWRjEOCDJn+Uu6A4KxDP7HooigZjJLl7lNeS0PA91ZIG9K0M3f4dCP
XqQ18IeTpptfTF3Hdo2jd5dqObHHrwhSLfegCUJfZd1OOw7LvFfBqje34CR4gVay
e5pySDkITp9+JS1o8GpQXacG0sxdrQG6oaBeoCspRONu3G8ucTyFp8LYlcnZqaGh
rSBSrmeA459Eip8KE5IClln9Tmo5QCvOmWcRpMp3tRIKpMFSKHjMZzBgy57hPsAN
N4sHScd48bFqU62f5nwLRdosRAvaMcnC7JiOmPOT6WychN0NZD+K9S63+fnQKL1N
vZDkfxDErUZXk1gEr6VLlrKI4lsa5L7/BmIkSxCO30Ny70r9yvfJXm78v/XAkvYU
l8lnQy0QZduAIpIk6i3thkoaXhrkvPsHSzihYm0w26NDrYTLovynZxwIXSY5fe6C
P63Y1n8toLi2YY4Vg4wMTnaD3NoRk2Qnf/lg64kr59uZ3u5LU74cNKlBV0C24M4d
fvhePnjEn7QH7CzQm/kExLtjiAurPcyNoRKxkIsYtIQtdi1T2F1WRyF7w6ltVUb0
3vSqwrLvMrXPYb59/2cmw22HJbGNVHQ3tfWCNHFUJ5B8KpvDwOh5sXDZtCHXPrpS
Q8ruNmX9zHztDlUBBg3ak9GlDGDt4/lu/IV19cT3gWrA9S+Nl6Jf7cURMsBMIEaO
dLuE23ce0OS2x7rDxbzsU01z78+wy4AQhXhJBw352dea1b5HAggQFUF6LZlURr+X
j/t7qOs7UJR0U6/QJsEw8NMPdnUDYOFs2QcHFw3ERIOLz7pmbqxr8R7e3uZV/blY
N/8a6ID0Pw+eWkxmEQ820oWjNNiPo3jd/1NURrsP+WaXwCri97l6DW9KId5OgcmP
bpJg25Ro4ay0PRHHRRhEItsoqvh/VoUhfb7V47K3Ftw=
`protect END_PROTECTED
