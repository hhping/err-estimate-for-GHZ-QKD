`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pb8KFIdqVNmiuH8XT+Dvi0F5WKTo8Xp2g3/JxDtQG3NuYVNBTnvo+/k/evUJ7SEC
Muee2OaOCU0lIKoLIguU1yLBdtfk0sL1KdaR3KhLorkIa/ALB4pf7L6BWyS/d004
tZopb4+8R2hYS40QLbJGVx92CcNvVFXHRaNgFZguTRwVpYZY/6kMepDmsqD0WNox
uPKnGOZqwjTFoastO0L0VQrCUmtjNTSfeFCPhYMbDzaaT9tmGdQyNtHsnpzRPfAr
veNvw/sddnyB0SN6uIL8jqU+0r5RAHE1arPYuJLY8YEcEQT+fwULW3R5DEghvxoR
Z7WwpiS5vveAVzkFU+WAZDCFyw6coe/O/uuOlv/Gb5J8Q9F3gpCXm3NV8PXWE0Cs
+6VICCcSMkT/m5v/gPlu2o7+k8K9+gef4jRJPVpsMfm5TdjQwD/anw9WOjfsqSGw
uHRzX1VBWuyaQ2gwQ5N9rSid3TrmV3N7WPY+z9QQj0jih5j35tNNBi4nypXY1oM2
zAk2/ykLzpoK2J1NQjgm/6VtckjIEYiB/0eGpJbY23aPFUo50U6Kszgu7NpC1wLc
O6trq0OEPeb9I19R7Pkk16TYfuUqX74smKqu90L91aW8lBls/91sZZQNH+G7lw6u
5qC/deSfoQdm9dig32fFDhrdMhGBP+oV1OKQyn1Z4lHu7CCzSzZkYwEF5rAFQOjX
8TcGKe8G9i9KOI4LvhB9UNcDmXblBi5R/Pr+Av8ZGvEUObsHMu7OU7VaOULDEg9d
cN7jcuDf0TeCl6DUmS9Eu0amLRbG0Um9UMfZq5dE4jqeZGHn3p3l6KGbDzcZ43rt
PcWhHaglIS3argFopcvOYAYfBpsw39OstLVEWBh8PthpYBdvIK8IW7dtTjzEsZiC
pzcLQ18gxhZV8jcgEOOL3Kdx0+7P1Eyx1etKzUkA+gWzB6Cy9M7jCqwx+Vf7TfTt
0UkjJDoyfi592/Du9l7ARbIFDra5LAXtq1zvDAUPcZWRcHeJ9pTR9fadGkhGf/3z
qfy2xQYSvB2k7cWB4E2mq1/WM/r56UKU5/aJZpxpZRQuKx2kwjfs1usWWtREPuWl
oneea4yL63nqCRmzyzT4pKcNMNLRI4TcQHLsmFrhJZtSTa5iXOhlSDWMEXl/uaTU
Y8zDrXZnoPfO5TZn8Pt3o98MjE3EWG5fiPTZAWDopNkrMwJ5s4qapikXkNi6qq07
ZTJYWRWxam+2Drm4cjlML5mh1bI91l6zzCs1TEmeWlabHApwABqFEsltLGgty5Ap
gVXNLrstn/Jgd0a629LvAT9KkDjeA1JIgUjudPBJ6ZxVDPd2q7KShL7QM2kmOI4E
OUKn/nwVpBlui+xVyo5KCLK1U5HvSvJE9CUlkVBZXm5HW0LAsU1AhQsyZi/ZtCoI
opiPw/vO4Pv898lGhQ1BpkN8JUqsJ3fJWIm4/BHdQutP9zF5MNgF7A3IFwU68Xnh
F5PaJ98gdMFBom1PgBc+jxG9+DlAQsa/q8XwInIJAGomPUvTyUzGxRJLDBOhHjLI
q52KC5rKR7MKG4Brz3NeGR2FpChw5bTBlqdMOvMemuOdla/VnUaYzqR62Lj0dSox
6TuPiluL39z0n+Uhb3RNsnROt8yzRA6VE/X58/Lh6b2yqopgqNqsjhsj1WU6nSQO
RoOSedC3wQBdxMFmzCNV4esHPFWwEPXs0Ts+2557HJ7UPbED4NH1m0D6Y+WMoTbw
bwdhHedYeURcTZ1ftvyE0b5w4XzAp3Mdp4hFx0XCl+MNWBYT5663zQ9D6jvyZ1Zg
n69F6+cQUyAuTcE4hajP8COBP44vXP6noz0PCmrPD41+GyYESzd9l3erJII5U4kx
VSr4OE2nPw3oOpNibhP3qO57uFoj3LmvITSIE4swMpSABSsEc6XPxZ/3PtmXYArK
RIPFYCmo9Q19MR3rmDAZ9TBWeoxZ1z6dluXt64urM3nHGJHafIi5BpwGoTgAg9LA
ZYOkWPKI0DdHU9bzAcv52L+Bn9yZSaM5BSglTqoSWOgkasNclfmt5zajkuqUCEQW
ToHgcnPOK/aC1XQHCiflERUhc6zv25/IyakCNtLYq+TVly4GOcxRt8LkreIEpgDj
3CNbZPdyqWIZnOXfz3WsTAqU2ffwg5rc62z3bOm0ECyma7en0u3PhddBT2iZ8qxC
OFcnV9YutvADUd6hviV6lCziktFtMSj7DKXZObCxBFd/vHGABwlG+VYDsUxYxwIV
pgyLr1bcrGHfJnfk0stEU79zcWpoIB8a2Ht5s5RjXAOJfte+sXwlGLyxp1jZCG5t
KElMmMvn9drWyl0siBXidcA6glDNC2hTBDoLLoXlSYloarUbDUkcPsN8bHN+wZkq
n6ls0qRPVMI72R9v2q0E8EIGNfHFpUWavpt5DhWj3LhqzwyriFkj8kx/6Wne9GaG
tDW6lq2n/CC4EJbnyo9z0ZAaUYwsY39qFwXpTte1Js43XFoOEGtb8OAiROt9foii
6ivD65o/io+nFk3wAQnm3krbmjRgJenphUMNb2mnGEJn3Fyte29XrFExADW3yh9U
UZ6k6EAeGX0b9F5DeU1fdTD8wQyfgLjLN002CmnEld59tAbBG+0qSfuK9Jv7sE2c
+ZzMj3ObjvyZ2QFR17nQhZy6dQjffDpfTl//adbzcGlZKYHEeLhtWcZetzIjolmg
kHeiJjbIblaVAZ5+4wC7ZtHOx7rDWVEYEaYPCNgtytqXyqzQjUjqfQ3qPqyFOHHK
uD55Swx9n4gLsZeoJo4njsK0bs8zaqkK04gt8ocWYt5Yj2kDz7dJHmM28qPjDllL
H9FCBYki2zSTk1A4ScTj2MA18JVVmB97fsqPgo63vRdSu4B7cozl4kKV08Vt6/Mr
h8YyNR+DAIe7VGRl4PIDGKMR9lUZlfzDZW5XpIq3/ueS/SNY4j6u9UWRdsIVWRHT
o+x9u+WCNFdh0aMT10aS0q8CWcApssE5FXhL3GpPIxaXdB0LdbAG3ER7+FotAM9S
ecJ2wLM9CflmSgi3LD6Cd/tAc++aRUmZ1Cc77VH/EtZKMLaIwNAuXrbFN0/8BXJ2
WuS5P53zbRUmwtN20G6ZWw==
`protect END_PROTECTED
