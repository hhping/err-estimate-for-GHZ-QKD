`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0Gpe+QQsyW4lsYuc3OcEzI4z95394uIxlFysGVfvKGN39JUQr/hDkiSmuENFnYW
xl7LL7uZd4WKfeJ725pRxr2hskRuzxhuaxPPtRlOKjvxtpvXXD7M8NRkSiYYzgH8
UPAg6nGJaimjR9jBV5tgOq33M0N9Cvi9ndn2v0HGuXrs7rnIHYrQ3H5EOAHLGEPb
ljdzwahapF24dK2XJwmQXev6xElpmQkS92vd6isID0Q+l2VVmu7Z8i7x/3Obj4Lc
tKf6J1Ko1/aoyx/VQMFBWVSggWx2g93sl9OPCoxA2l8xG6bEvG0MmkkRYj2dQOpm
sXu3IVvz97susVoE523Qxx0sqXyO1ZygopIgI/HK/P8BJTBOYxmD3cKlh9tTtH/y
nSxq2TcRHuPlYzPNfmz4nGCAHUi5vFqyHHZ4VoYVFim+pJlPxfGtF1ywS524gkd9
h1G/Yo+8+2DkiBBr3WT5F0ea8RFaDRwUL/c8O7kh6EWvs1I8BuJxjfX11cLJi2M6
ZHSTAWGWUUweKlU73NbarMm5b+oUW4uBP3AFPDhu6BfkyKNz4JSgLwwyFV8ibf2t
ctfV9Q0CGN17Z3SB7CgYY11y2AdRCSwn2GuU61fjCxdjMYO1WyyOU68QLC3mKwVJ
zIKTobjJDEAr1p+HBbxSQe9/KN3Dbl7u3Og7ZfVtU6GcNdLsvptnS4z/jekjBh/+
pOrcQun8LZM7ZiuAJFjcbiKeYAOcFZjPIrDEKaKvcR/a2hu9WpS2gqZ26un+Z127
5JpmvKlgTQ1n2uOgVegopkhcmYu1Em8O3s+dUHMkdHXFuDdwCC+C/TgUJNJxkwWG
yowi+Ry/BDQb1qwl6isSMU8SFK1TE73ZOebq69GNkbo8KhTX66geFQ/hgtcn7jeR
XnsZ6IWLK78tjlrxUwCdiZ0pdQUOd+vykTGygaIfGA9L5Q3snsk4o+nIgItZAiHN
Rs+UMSJlZwupFmU0OIoHAw/RgJzSca+VQA/Vl7pGZyv9bB3uvozaUCmcxBH+B+lK
IUPY0Y+7PbEnf/6avLqMqVIGuEWDvjrmhgAitws43zxX603ekSV3aTUfC3gvM7KK
/VybJch9tkaB5jJBbyZZnbxcZqBjLjv+jreJiGwKsfhXgmLZDJxo52FVgRitOPw0
Jzgbya57BUfChDDLspvz9d8ro1Ls3WLi75cj5nsDI7OeBhmGNktt3WpfecdLOb6D
yL3/S79umfkAc3o67G1gJVouiqnbYfZsIToAG+hAb3SiZizp2p5T4DRsjy6x++XI
BlquSD5ci8Vy95xFrc2+JNS55OYkwYWW7LiTSVtUjTCq4tZhYYf1fe+mJR8hxRNK
wBJt/MrUwHCWWdDl/kVAaRhNIKoS1lkShblWjsRIHsen5NiII6FrPU/l3IctGYK8
pWHImENuVr1M1Onnb+LwlHaH4CQcvul/mXgpl4mUN6hstpHQmxbUdg7otN/2C8x/
QTC6E05OFVy6SObzYEjsaB8/3xYLBHkE7N/0gbff88vt8CvpIb6k2LlyRxjBGEsL
yUFri0XvyzsnTgwwyvFNlIuhx9QXLhfUP+tjFVaMz0e8ICbAF4LnktSk5tEAgj3F
Y0wzr/T26+NtzRi2ClWkJWJnzyeXTo2cXTpQnoVhlVV+J03jQJAPOccoxdkddGvk
v3M8I0e7jsMc2Qx9QHQDspozMIvxrHWadUwH2O8fBuqG3CuvRbsOq6yQTgM6hHvm
j7hl1TemITZMXKPyrlZ93yvxGoLxW0Ay1G5pK1T8vv0tcEUGb3Znbr3HRkZV695G
HhQIgWQ+GdOmSInsLjJceer0CpTQ25WZPZdoMfV0W3vbzwLhmCIAoxzPz0kzvLG2
wPzZyi4tOBk8RfkPLI0Fdxtwkj0ovGLjVE84H5hlFS2J3WmKc/JxNj4MvaqGkYGe
nqOAEUUBSo/pIMVWaqCekxTPP2JYhiBPOMoIYUVUSoewDjm3jWxm6NyhDo1J8RGl
21f4fAElHq6u+6EX2/utqdFqTB1DP9ll/AeHDkSjWugdBjnZ3EW8WjJD5MzobXoe
eVnb3qeEjKYOrpUbUmBWhuwnQ1C18kkawS/eEQQfEL6+2IbF0ze+TdwPwAhaUxVk
iOpWm0q3jtJPmxwmOijuYFuVJ4yk/mwcCXeUSENnAV/tytjd0ub98B3VvKLAU4S2
4QbeDbEvAHgDrJzYxdqUuAFU6v7O9ZsgORGPW3JYwT+/KGF+gVf5ZqMPmx3R1Rnr
W+a96pClpFDCQd1DtijWYCc07srDARN+mFk04v5T8pbLEvaJgn+K6p+1EWrbnOKt
rgnkPstN4DkSCw0UUGduAWYIxk2FrdZRSVZoTuel2aScvgwKuK1IoVAE88va71qV
KWMouWZ+KUjwErkmuwjbjRYJomW7ryoFSzwRVA9q2hf0mLcO+Kyk2BV8vKPnJ69l
ZNbTtOBhYXbP/wg7KNpEObjRFgP+SdN2Zq8sjm1DzRHiUrs9BFqcZce4i50WCZKz
VHf8kuM86run33tJJJbWWEcjpz1TA5oJbhEnAnt9+TraPN8a17BmIgnCV3LVkCUu
7osKBXnFCdcZFkXesdn2Z+C9CZcHLKUhudWcrEcp7JXnilikqAnbYsVnZtiKBwel
aWhjLebz6NNslm31RmovHZ34CdR8S9YHqBR3kjUMq58v1ZFJxbmZv2ZkpwfNrEbr
nMEc8sMIgHzA8ZfHz/iQY7e/3CNm5WOBfp/kQ38NaJ5Tpi5+5/apqi9meCFDHv5n
/hGI2jltmq5c7ktaSMrg45TGpRiEN+irRSZXqZjFij7dzQJ/x4IZzmLHgcxYWgXW
EIJCwVXTK40Es30bs/n9pMLUZLF9shRLvxcS8iEgnIoFNxy8m2rwxU1fOTSzMU+9
EtWWQIZh+DZDg0/8usccSR9FdiH/0kkAKkq7aeNFJWF7NMeT3ZLYcl/r1YzKF8IS
qNNSkqdYHP+5UbhKxKOdfHUkRjWIjSIUWKaT4GMi9+jfSEHf3drRvvf3FlYzIGRW
IAzzUCXY9z82aAjNZuIqj5Fo6Fda2Nu82shsEH8X4rKaadJVQrWPsCMhn5ZvKFVv
9PD3ojhtiq34WWtiP9iRWHl/gI/C0NEINlYcN6JcsOponqFacisCGGi0GBX6Bfer
wrR3QhUgCx1oSPNndBTsax4ql0RiNV93K9xFwD+OrHFLWVKOqerlxh5PUXcCg1Hp
q0h6Tab13Z1cEG8BlEUNKrfZCmbcN0CyZfVjlOyNCZxGSvTN6Tz84rgd+GWLagL6
y9DqRlDKXTpISQILFDeNgNx7WRnTnDCqUUmLcYdL73lV7zLuj34bC0efMagFZQwj
F/VCqlKoADhTLcD/c/3xNudEnOjT0eMx0jV1CtBSNmc3F17+zzTb9lVfhyuDfmx4
hFgakohIJyfqoZ+bBQDObq+Ps1utoPz30FpctHghssOeFBKdGlxA1VcNRbuBsBnc
zlfm5pFW6GsL5q6t/6y0pv679bd8P///QRZWpwU33zglvCmxIBQvJghVXFPwwkg9
ywarAqdSq4q/pV48BrGQWBaguK3/eXL9IKpsJ1eUu0jxHA9h5fpghDmTr0pCQjt0
na/uOACM5iJaugTRkqQNbNELiLZ9HFAjmzNw8qpCV4b4Vsliq8/eF4N0KL402K3d
I+O3ngiH/EsetLJUWABKRAMkYTwjCRoeMd+nVdDZCLX895r/xYWTSOI8JeKN/uvc
TkE6p4wakCo6sCWWrQ3FbvTPlOAab999sGOk0AIwzRVizjXA25Eo94OCWQa45Ijf
vA6aQThPxfbXicdslhHprSsCUZ5/3HZ3pqWB6sNHb1Eyty9+7c2X/yLNKzB2yP/l
Ed2Ve1bcvCmNJxOAgkWMCZN+J0WkmqNCMKYBCZC0IuViwJWMZU1wsAbHETaOOmPL
1KMua8EP7wNiERujHwIXOLtZIG7KGAKiDIC+oUvITnv62GHdStoWWd+0FvCPgV4x
LnuT51bVBBxF02qsIWq3xJildtyb9X3JQnH231gcuPhuj7yOZwdbcGpG25nsfmMJ
KVc2hu5cqhXquuOlRbBz+/TM6fcr1yuwyUz+z31PJQ5iY+t2JYr2zKr2qvJHXXF+
o4xzCXlHbV7JkhlOokAxu3Tn0G8OcT2wChgEmy/ImJVdJSaBnIn0XxI6GqiOQod0
kcaYJVdjQt8CD0e/T9uInTfLQfmpqsJzldFb0czvb16AVRNGg09NQUmkAxmhrE69
vuJZ0DzonVcCworU27yJmxUwL2Lzs1m+tS9xEnybOmhTnQ25W+7MTZLZBvv/1JeO
A5crmVtclDOdHAiEkLF9voJCSEbDK5TwcGECLdLV0L+2ZRM7ZpjRKKsnM+fmbagx
zXH+xZL2al215+3DN8pBp8NOY0BQIJqV5lsyHoFw/AvoqxjJnJU7vte3eseh1/YY
S1QSA8edNjnGtcgqzwQR/aTGIwe2lNdTacqKsqzYdwSKEXAkntIXngVy1HJ9O7ro
PgWupWbN8tTuMD4CIrKU53w/JWB8CxYfUIfclTRHF1jF6SUavAUdhEi8CflxClKu
rakbLAi8IUXlHckfxMWMq1yv6ddcaBj40kq764QRmf0ZOCuYgNEzkEg5fNbe5KQc
NzxKmeiWbe9ZgmPi+p2a5qjwZejzfgGdysMD9jAhCk3FCVzpK3psMKNsVP6XmeIn
5mD1ztaE0DlTyu+YT1GuJndwoLPPvKPKrccu/b/6Sdg/Ip/+2MhhLsddLgNzJKeC
rrpoNUGWvLnpn7zzOGBBWyA1GCm/jEbYMTZupzwoIYIgxprsJUna0IFNaZfAKSGT
zU5G7a2KMFT1h2wc50N6seKVQD/WyeNnV/8JIP77Lr76k8/APQJpC2z0AAVrIDc3
BTI7vqB2cKUjDtXr49Ezzw==
`protect END_PROTECTED
