`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k2NWvSw1TKDk84zTWSeay9iXj1jg0408ATaMrRr2zFBYlXqAe9m5SqxBtGINRfnX
XtvXPK3XDKKKHOWpi0QQRiqdYWVBackGJH3+OONUOlTqjKp43ovgbIVz0KL7H8CY
gXrlnqjcqJyG2Jo9roYiPqFTFEXQai2lXy/7pdfGNQIaWjs/bFTVrKDYlIbdsD6+
znJ4z1VYfqrymaAKAkQLMjW4SQFXQOFwYen2x6DwbN9dE8ynmZWJyk1E6K1X/quJ
AEN9I3akatQycP6SQD+iW0rlD75OGAhnQ9maxSIDKmYWjLiBgNC6PUB6odOhyZvo
eVsOUKgmctPkIgBOcY1dTIoqf3krp22jmJmawktObnoytshrYYMgbowWMH7zMFXr
Yqawt2aCLUJnwHZf7Akgd6yEEf+AbupoiE34RTl9oZATPR34oB5iII9mKhDIqzrU
pC87Uu8/qYDk4eF6wlTSFs/7UiJZL30ZqtirB/U0ZNaPMV/9FT1nZu4q6INzuGSL
D6uYYhf9BCw7pskNSMIbf82Y1URGtCYKABY4ySimtW0ysUcIYPtXe+nL8C6N/KjY
ifligv/DCGwfml6G7zF6A4wuujOwWnkW32CqGqyOMTwzrwrtpzIA4b/2pPqszIsG
fuU8wxwqyXHE7nS/5NmYq41gR0NKKD3ozmkoyg/emmFWnYoY6Rpbgqw4E8nn/8jv
FldSxIQmIPvORbfv05DKgl3E4ma/U3OAJaSAFKDZagwWFb6HMpfjSPAXj2SaI3OT
OFgMQ3sS03tX/fVRnrhEjawHn6OrC8f7R6KFJvzczTV/6nbAi4dss6cxraaQIYmg
FQdud/5FkICSJeaXqckJ4O+GSebu4UPuX558wOexqsi+M5YQQR5sgmysLixsUWZr
Kx6dOyhdssJRAi9FWX6BV4q+iQTDencq3RmBiLyNoGsnYfQwYoqHlAyfR2i4YvDw
duuWeKrlSXHDjlohbnapP4UFRPB232jyYOotwRzsgMWPwMFY32ppT8MhJ+CIEheA
wKh2N6iDVmwb+oue7M/J1YhJXjnmpRk/21gAvoqBdmPhQp+ij6gQNeTGO5x+B6tH
P8ChD5SIlyDAW/DoOD4NDy+2RqXNFTpIq1f1GfmrZkSvQ26ZzA2PaLkWF+++Hf1n
FoQIpraubXecUrvxbmlbKtEeki0a+DZARPbaPlQnpysSxJxgqiF7WmZsBjGoOV6e
ewOQswqpEGDQxGrVSC8zbsVsnyNg+vBrp0tIgun6TiYPTy+paSkfF9OFCitT8OfB
so1fls8cxpgmVIZJCJhSa9QWL55n6ZF8ddDqP8GRM8F7F+WNoLmhYUBk6d1f+UPZ
GsbEA3TYF+E8bj6Zv0WQotG09ZKbaNw0A18iH3f30lA/NBRLqHiZC6sYv095A2hw
s8RMO0K/gPf/A78nRAx9GUrNqX5HODNi/7b8h+oRLGYGEmnL+RP8/QQmGmShJiwk
gfOQYxicbjwmYy/uxcDWofoiWRKhUSh9EKILXMCL368NmP6IQCr8TEjdd7bHp0+4
1zEp6JsK7cd/OisUwgR/IUPkEPevDZiweAR6oyGBMcroCYVY3FI47Ox5D2VJO60L
ZBiUZI/JJxEDTCybTZlE6ulLbJPyLsoTw9aVTea2bLwoBlSNWt4kXBFI8/+/g0KM
TU4yZjeYdsv2f6kbBFF85MoPZTSb57I7R68FLn+Y05ozV0w6KQ3taAN6AaMqA75v
GEZlLH3eVKVVR7wgjtCuzp2AS3sNroUMg5McldvdURSeaLt+Du1wWAHGqS5QI+Nz
hiVhhEZp9lVhX6yycYF2zGXMBbXKywduXwHnFzw2bnmGZ90TPRXz7HsSIMqitEqE
w616ndXzpHo4vWjG00ULsSoS3iEX7VbSX3yp6gx9mT8GLgKtv5djv0HARKqVJ20P
TbCB+/le6n7HyTWPHNXLQOUOZkUUZfLNmOr1z3eVO4rwtlcHDYHaQnN1t6TuvUq2
`protect END_PROTECTED
