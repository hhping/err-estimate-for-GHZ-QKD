`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiN05S1T7s+RRiM4vdx7HniJaG4ZexWtdUIeaSd/otmQOpXMbGeU3wDRygmyLRpV
qeGe9MLPRVSW0Tsnmd1tOMqNZuFX39R9QrJ4E3SvQ5Me0i5QdeC0XLYfwKf9L+y+
DY8PqyeCS80lB+8FgYr9bIhpdLKCkIbFuW+9p/xHzuQhFzU6jYsWigVg1UBtF4xz
5Reg0vuUEHmZ5gKGcs9/XLpYP5On4V/XFe1uRJhniAePvJqk0zU+Xtpl+wnSHJbo
5TqfMbGA7RutHoh0dV88AHBF9LhZqxSuFxCiZMv6k4BRpQS+3w72tgGGojQxvEjC
+nJ1XQJjWUWDMx4KWsZHvLV19Ffkb3t21SJ5mITQsEe0ebX/tZy5vSUeVmm1V3o0
NwId3aErNDIeFrCxBK+ifGQAp2wM6iYTUfifNNYvREnF9zpbaIZz9XguasN+xqFx
UHh/Qj0dwWTlIpVb79V4FKAOd9V88hVrPIITEFQFiXLqKsH0Othd4ZTuVKQnIKKY
dUOG6WiO8ZO0x4O7dyNGJQmXYbdcaDMmuBTW/AVTi1qywIanEZYyvpwTGSt0TuJh
103ksUfWx2irgUBIOZEwxidqoY3OKGvCeyg7FNtwG79ymbZTYE436w/uviWkjNJE
GPAW1elfzKuaZfv2qqFlq5KbPaJ6dFEP5Lq5RBnW8h0hYrZd+U02O+pw/IrVgMoN
m78OsqxsjdejlnLGRV4m0LQ5YFh0CFFJYSRrpFG6W5lECjZlVUhY4MScDFxdgpZK
kmmeedej72tLvnvsNfewdPIjoKxA9M3uyblNw2Gx402VSz75QLJIG4H8PAs1mGIC
PTOLj2zSLWiQiuFiSuwrFqjdBkS6PxChsQlO52MjBR01sekZRwz6e/O4rpi4Un7T
LxeVi0AkpfsOJnZ7kq/32L3Og7e4y0P5iWULujLOyZcuvq3f7AZuzS5jX70Vjpbz
PdXwQ5KkELoK2UxPQGgtAJR6o2PZWewec3bgwWV9MP4QjbcNtJnhEOLd+4pPo3XM
t6kC77QKKpx/uk9dTdPjMO3XrkXDnHZ23yV/T/+kBpbC1J/2jxN5KPnI9bjL7Heh
FK4mJ1xi2vVOcqesId4Paf6K0/zSggr/nDvllBoEcoAE+rsSt8WLnWYgJXqe0/V0
EslLAR0oZP4TfDBBQ0wq1iUeApiomv1qTgxS5LOYmF702apKjiIhOQrV/7aKTCWD
/SUBQCGdyzM8fgKN4lPm/DEwduW6diZsqs/EjXGDvzavxwAEXDceY8iGPWUvNNCN
mFOrJh4BPcQjiOYmN5t86/68ojLn+diDPO0cowGhKwgISeI5AAned2RCxcVYMA1/
nXElAcRcUJIz1Sua2p5yb2thjqgAO7t2gGO6/MDVmAtvrayS6w92M6WAVYY7/m/l
ptaflZPedI84vYoRlqsUv6PMQA4Jq9NOzkJxW9zrWCwCaMz9qcPe1Etf254ctz/B
foNLxU/fwZlcuYBvh3o5hJALnQX5bm81j+64ueGDm0g6b06PSNPR98OnW2nLIqcZ
1R+gg0Hu7W8sTchaM01WPkv3rlgGYuccOnIWFPJWTfps6ra4LF9HV2mw7OCjmZhd
DEWNTjei8qHoQLbG1YzYBBhNmGiVuBc9Fr9S6qSVpAEItk2d9Jct50vxhlwuQyyj
YculZ67A0qzENyvooi4zZ5DtdpWK88/Dh4dymwRcVhBWpyN5u7RpG8bEWAgi9oCW
jaKjczzmYdm0smMv35eSPruxlSDgs3/xD6fGSmI3Ts5rvCfWG68dJDLYT8EJnWJI
NOjTpx2sMBJPyw953BU+1ecEGYGKuXy0UdFHC1Qieuo+RZM3gVtFUMLUZyA1026D
SmUU3dTAOf3nTr0WhBIFu+ZBY+tmWntKA/YuxxlcPq+jDIesKN4tXY7Ta/mWL5Jt
JrJxL7Y2Zs8yBohasNbfD3WHlfcMfJP8n4VERrX+tqCPGrTp9Ks+TqVyXWFruDq9
0VlcFWbnQBhXs61/LimJiKFDXqPdbZCHBN3onDPZwFGoDYhaEiJDCKVwtWydFlbF
ponRzb8YD+MRph0rTDDVhFzmcyayYjy0Qf0iFZDL6y49GCbkPAf+uJADuOz157AV
OEnaQeMRBUHYDFDQuwEUvfI49rTmhPevQF2zD663JEmlf8B/xdADxV1MspIuAlaS
gNs9iyndkAvgO4HvNiykwwW4swd04P/y3YN7EfPnmBBPo60EvRhMA3wqpViJQrOV
4Vub/3u74ilHEMWKiiS1M3tkg+OdGrXClTHP2mow7W5yIHQzHySq8cvTJshLThp4
FdlQ+ZI0TkYnBXZ6clhuR4CRDzbnJyZcJp1/BRZUIRpM+0Ts6kpgqMpcdbBuCwDw
PntyHjLuxOeQNCWolNT8zar0jT6oniTXIhx2JtIfY9lbYy10PTP++MzB/FkcPRNy
rQhztR3kX32r059f00WPvhlXUwSPVInxctgBsf5jB8THwREXlT5hk8E+oINPadQx
zMAtq/Rgv4JEf01ZtJ5EUNtpsZ32qvbgzlaIFWRLWdK7zx4NhGrzSfOItWZSU6n4
+rYAP/JGbtIZahA9bGSrnfPm1F7oD3whSovvCEgIFeXfB+DJDaT4Mlx73/4TB8S+
Xk4mBKLoVzbQRbUQBjFGrCoLj0pQJ/DFmHCu/gn7xEAiRyjy7icTbAQA4EpLR1mE
t9E6/Mgprp1sAfIk8JTM/6/qUHXZr3EwG/qlpWB6OYGC4iK3ZQ/Y39qJhcJywAO2
y+PorU0vI2rARLpzn1A4VAvXYb7x6NcTYDtcLTUxvWxJ7QjH2lYYT45cb/KyQOpM
vYs271grQcTJqcA5n92eyzA+deNdNtk+9Ij3T4KlAtAdbZMLwA+By0rT4QfT9D5J
+ekeZDLPeaOhhkERj53/T1XLrPQHosch2QWAsOnp3A1dpTrdiuQSlOHnckmdNMTZ
ucCvV14k5neMp0cb8lxmUX8Pg239ePG59Ob3dqnYyZ+m2AQ1CWtqQnLBdsmd9QNY
kUZATe7jL0G35z4Y8wA3g10e073jXDfGW5lTFShSCejI/e3dDqgocP92KfKQ5MsG
SQxjuMQIWCfgXQzQGWvlYqiwSVBPrXf5b5z0CaOHd+CzJ51eMFI8Iwy/EmXBFCv1
wcYvXVx0dvwdwrtX/NKdC11mcDTwtGeme48Tw13mTeINFI0MRbAW3LMy4oqqIfmW
0LjnxM7z1iCOxfh6hzONZtH9W0EWmZ/LJ6TvUCFxEAitHCue+AgFdidHhS8ZaU3C
PG6aJ+UxAMv3jIWq3qO4VBS5sUnkezytwPXuJ9o+9ahY65R8dHDBafwMugyPSRMm
/+gmr8oAYhvcPpeKOHTvysg8S/bJQERbKxcmHm9LpC8O7//fogfsVpGU1VDREsXu
fRw+eNlRlaj7pqOTFFNur542I4dCt/AVa7gqJXX6mQsLT9vO7R3iF69C840mI3Ap
3jTTm6RlxHSsXe3oqU9hHV1FvWJVsTd6PxYYd8llcE4bOeaQchALLP3vAEx46+gz
dxO5JSIx2IeHSjwZ0i9BkUYKiX8a7QuFsunzQH2VXCI+YSkboSoNSDkB0dQuFh8T
0mjmNVV88/gHfZ1JWF/EVQ1RXmVL8Ks/aRWD650RUksF/J5xMdB2OzAv2KBkJIvS
yZ4Kng8sdeRwSCDNPt0+oNwwq6sVTxZqTOldtlctg90rD61s39MKzRDM64KvISl4
r2uWj1NI/VE5YopYHSgCdlaXKjb4UmTqm5cj3j323LsMX+gz8nze7RHJKLsFescJ
6a1C2VCX9Wxr8iSq6fbW3R4tgZnB7Lu8lJbPFvHjYoFIlYAFDmH3Dir6LNe4FbkL
EmMINRLdZ0LTdS2Ud63kJw6i3EdbJia16fNW6pfEw0VAILI7kU/qz/pTqsKVmHUa
Rr90Tj5RbzJhVKvxqNAEPTEsVItud3aIp9Eh9y0+sod5usx/oA6yjP26W9jQKSwd
Wk/WFIx/PrTHA6/Mjftm7n58fBA1fznq+ebLxwsXgY+AP5w4EzsL27dZxpFT/c5T
n0guJHDjkrAU7xNZyDrIGNKtJPSD6YIqqjWb2SzhNt6cY1WDIEcX2YZjdzM3W/4x
844oFT8tjZRjHNBm/kWqh1c0iF5yolUUTxhjtZgIU8cXhrqhle3VrUaO6BWNbd6e
C8Mbl4GCCieBglosXECzOZ2/7HYN2EsUiHIFBzVaQnhuv4WxepKbCHcBz/3L5PWO
9alvYUYPLDjmG9xAdPUk8jGnTjZyihP9T+pXFl0kg9rn0nCbM0LDCItvbb44Db7H
Aula4XWQ0lFF+cwhvkebSC08huqTTTCEe4F+GEavCYH+xr47JA3hQi6WvKKl+amG
EpJ+WEuIcUjwE0gjUKRIQVxQ8VMxZ5esXPHfNxCvNgCayB/bRBbjpvo/MHB4Aa9W
kLH3mpvaTxpGmEOgtnZ2d+OIKjkf+KUoKocNA1i2pNYT1GSYuETRJ5b57YFI/rbP
P4UDTSSj9GzWtQQ6d+2T0AGk6eikkabzJicKrt4IEs5ozkUe5JRXx5gz7aR7irKy
PwofTe/aDFKmjpLfO40f/o6hLxSAEnkW3bS8qysarFgjeHHpshxFaLPM3JMabM4G
efaY1dUNVn+8Kck0rk2ny0GkhTnnWzacoMkiUbb+zswlGR6d/6hUhUSph14Rz3TD
uEzZej6Yual2Jj4o+TKJYjUS89mlXSRbx4+LXoRJx4GrK4MY2efugXrn2HE5Pb+W
5o5C4aM6eAmcDZDuJNu9KBEe2EtOaVtXyqGvqYpVLHFxzXdwCuZ20x/eyZ2o1SN5
pIBTgo8tpKD/lIkOidj1w9AsEZu9HmrH2jUTH4JEHI6R+sR9nR1jq9oLcyc/X7+H
6uld6ygoiTnba2fAazSG1+/nH+lle4ooHIJe1sNarwHodUC+Rr1DcwRZkiGheynB
x9qDl5HHnwZRTByFT1QTyZ0/2GdFGA7IjfDX9ObS3UBYqrpz3j76jF/KOufsyjUc
lLScMkSWGQQtxW25h0Con+2ADbCKHoNC35wmuPFT7/n8ldJFU1PCN5eTA8+HOigq
pY6ni08OMde4Ho/gULnffsmMT7dvY0KEZd5H4nKXAzcBno/f5IT8OvLR4zjxH8/e
ml7E91SMSitEbYf9ZyUIP0+pUxxGXxSr+6SGBT1LjURyQLg0pZ2NYVyH12Sfakj1
fjTeFy5xPR0FX5aLlMbu1Qa//rCBKiNh//u0Bbug/fnL4rjrEXEIEsJkCKj22zPI
Ch5qFTh0l46xE9d63ZImwSmY5+N/eoMQ85oG7iJwcRrQ7zR2qUrd2kVsfVnQL1jA
IuWHz5ILccWJZcSXlIqgCrwku1JkaT9tm4g8nNnFmMoTLfNbXEPi+O2x/aQnl6WB
BO6EDtB6RzG1ZB1Xx76wlLSJtVfZlWs0uTGRv0gHobKWMUuWPhb11R4o5WOKO20X
7Yesb/On47f5NPWeTV5D5+eZghKh1pSy0ZU5HLHcIUX3I8Oh7/Y3VY89AdS/nCM4
/3niyYmFKV6HUoZLB+kRQ2bt6YDBoYTOYimKIXQsNPBz5DlVYuA/IGPBHFx4LDcD
RJBqq5U5l4Dg0tUaO1Ob7f0YFitAqlGTxm+/PEYn7Txo+R5duvYimz+wWyaHPOWH
sGg8J6dN5VkfZqapgOtaOTigHLY8Fa74ngpVuGCBtv6185HUg4s8OPxxXhV8aq3N
gTXm3qu24KR4Zmyp0/4u0PXBKR9fBCpYQ4x6aN49FlxENqsG/zpolbD5EMPSp808
M5d00VtJM2kQ0/2UQFwiVO+q74urN7ZARWHwN9jZX3MrhV01eqAamBkQZwXTj136
qC9ojbVLZU7kmGZeiap3TMN47/03LnKUSvCD6o23+NunSXlI2OmoIrn7pl9XaJYS
e+HB5q84KLbo4DT0CFMdstQxfXnZbejl24IiVwvoNejm6OEzvHaQlqUl8tGPR+QX
2Ajl5xdBnRrUxIQoaTB498PChz9Dv394GBo6feoydte1sKli5JEkRBTzJee70jyt
a4KGOABmwSec8wWn7TUbm4pDrKPkFgsrhChe+HvTRZ9KejA491A5Qa//Qqcprd4E
UrUbc5UPbiHm+vaho0oa8Su1M0sjn79ywEg+xkykGwaOz6bxW4eQtNb96kbcT7WF
ikhPkcwFDiM9RezejLI6ebaAQ2Kid7VN/w72fuETlnCrvulXJ0oMZGT3+PDzO+P1
Mg8v2h14kYSFbiLPOY1mmIjmBeL70e7FotVSU8fwZZNptcpzmfIecfvJ9jlE/nt0
h4OQnP1UkNMjJ/JPzgCUXDYlJsNFzanc1AvYVhQLFKIdH7hIUUGSK7CiyUth4lBH
dLeJFQZCOWg0m8lUeKw9kzqPhqRLUDckcK4CNVcV5c4v4S9YCq9njQPoQiUQ+yBt
USodhVzfnpE4yuKZh0fCaRMaKf5tqK+vnYOV60lBNC9MESKHQGV2tgmxOxKhx/rb
R91b6YqZQsRIj43DQ4x80H58Oupunef4Ebw2MC/8VTbE9CN8QauqSVi87vwV/w1R
/ZvS4aSwdzF6mMGhHLgXtB12JGG+iX6GutdGELejDvJYhHvLIYZSw0dMnMr2qaOe
fXh7f26JTW1TCbnUqF5VYsv4x2GTE4IhIyseBO97HBsqLi9t7/cOImM87JczmVe2
cbOVHFh4oNwYY0Hy+Vt+eLpIpLUZgNOcZe1Yr2aIm7V9IwLYzKGdwYyO+9OA+SbN
l4O/VDp9W2LNWG4twws4Xfccmdel9WgFGa5NyFMlmQb31oBnYMbClp2VfMWplZaW
wAhfjPHP8ZBvCXpBLKg283IZkv5NWG3W0ehkEaSsHGGUQJ1hbwmqBupzTK4IdqrE
bcJ4KTOgGA2aJNJ3ECZpMg1ds7lAuAtqZRQ/qbCZ96BaCmlaOxjuwkgbo57tBQGp
G7UlU91/ZqcN+p0ppicAoi+FLOXNR3GbX4rwFqu/usDlpt4s95mxW50krUkjnDkU
qw6MXwHIwMlrs63vHnr26N0i5YHYZ7rMfrhcJzeNGuOtlRpUQjqDJXPo7r0nLu+3
UdC9NqcOmEMhoc9IhnS5GtdApMkgtsaPVOQou5/LWdvZ/ZWhWAsW9yc1RRS/lOGz
MywOWXDYWmSkEAOHl8p7RpERzNVWODGp+muobrHzL0tt0/w2FcC2iSaNG75WZptg
9jP/YNDWnkRaKgXBU0O5RLfIetuyAHvTBfwYVBzf00/9eJCOdPy3YGrzF1n0ITMK
bC4XeHBUvRC5BGpktWk33t8rDIunJbygYgzqm4AeuSnJf7xH/0iveKMoRltkV7vF
O0QcDA3Yi3v9P+Bvls2BITTgRcboBvOBBGZM8qIXoY5Ej8szZpaV4rjVCo6OPSlF
WsgVJfZA+p6nr9FwplYIkcO5z98ITvY3TV5i5d5MZ/emTBQVIi3gxdu2TOorjGo/
dsd6yn7qBf1p5RebGDxIPhmEZPbkldLFeAcJAnCHAsUtRSPzKVhAn9I1VX9wiV8p
0ma2vdNQOnq/gory75R7tFbi61Io79lgPbDLMufgJPo14igu5i8OFjUEHxC6ffqI
go1Q+wa5Wi5ZJQy0Jx7KYp7AOPe+U5aCRhz4seQLoWYaSlTDs/iqIBcDIi+pZHjx
37GmKdHWjTtBO4LGrtCGZYzSahzAzsuiuq/vSf1N5+hbma930PJ9ado1go9DK9xf
rx7iiMaTWQNFacLHPwO/k7xkKveLmzZvJARFqnTQLPAwRwz0x3fpNyhptS5f39qn
eAIfdmJBWUjlNT7WLa4d6DfbCnx0K/qfyPbXP2fjO9g0r3a1MtYXwysC8Zm9PorR
ghT582Te0CY0Ed0R2Pfm0uSkK1Q/xf9OojodAaSJLRxTTZ/jI4lQ4BXt4DLxcti5
k5TcURcrlKsYlc7kA8XDbaNp4eoOnQIjg1No9UASqQf5ntzr3/8HIlWm7m57idmP
W8fkTukyxnz7Skf3tsQb07UVhG+J5uVi4aS3A3IxoB1Iop2vpVgD4hvJig/Qc90p
9/s7QbKyADDNSmIeWhPJXpWkB1wQ30wzIqusCqi0Bjvm8AZEAMc7Gq5L3gOUB1fR
GbTr95riKSkRGrtdUiuPLTmE+NnOXXIuXcfv08FeEjZcDSHSrv/FWKUhS0PE8/ZR
Ny9MqDlfAwCLVQiN6NQlv6rEGHQ2h9xon/cfWQUvRkB3NcAeyIe86KDrs0EsfjnW
wmPSbXHNjFeFi1tCQzAaRN/WXFLwjBDn4EwBFM4VnBBGAr2Mk6eyuqdQ97eN6Bvz
8bqTPkhEIAkFO1rwVGm101LViscPy9jRNKGng023Edd/vcEsyJR62yyGsNCk5Edk
p/6YXON634eWi7j1+butJiSR+U6DdgiJ748EvdxakzHBg1jkGhsjVhHck5pbzW9Q
FMwBX8/XlT0Drdjx3WnEc+jrnpphaD07khlggjfKAi6Nlcf0b+JaRU3q4izjBt0F
TimpXiAjyze5XFPH6bwgU9a3fuApyUwfNL+eaFabUsi1IEnAY+TAQss5nu+sp77T
cZ1IgfPgXfMfNUv+tCQkyP3A0VlbrEAUVwFfHSpwEcdDTcsJgAkJQIhh5D0+Nnsu
bwF85qwkl3UcY/qxo5z3mJJKY65jbCsnS88n5yqqT/e/6v4PY6N7XvXblzrhvGT9
SycZrpUwTh1f2kwz8QfhUJRdGDmHH5nmjibYkpM4MKE0tvbsxreF11lv9WlO/QEV
stJnLcMzQ3hDM8PYLLPJSsxFI0IwDybk8I//Z9RGFfK63uN6LJHnSkw0vsJUf8bw
bV/6xAY1mO3iePLdnkCdx4eIoURZA9GJfwSgFeu4PnGEFnY5zSzrAcO3ZHW5d1Hd
Tg69tf3wdxWSktLHcWCWz2cBoOBKecSMYqqACgOdzJXiKieThj4tRljtwti2QPGc
RDzKITTsZFt+SswLguGmWVAX87IzHuFO1CbR9YMBnLT10xLqRgxdCLV0+zgo4aJ+
nXnpIbSLxn1MVXAwclCFeB8gYS9gmd5zG5V5JZvsKm4DEsjFnFrZAJbVKiL/vS7c
BUmL+iAWIilG/yKI8rqZbkvD+VEzve8sbVGn7MF+PpQc3g3Dj78eIWNWx8hnFxBp
emBtDeTrHXLKjbTpgpSaLebxxiNNMlrwVK3xvqR0Wcp6Ieo/yzqU/2rPwUOGp4si
seuU4dG5VqFFZGpzovrQ0HwQLBPFaJKGs9l2EvLBY0d+6c/8rbe/UvUWjGXk7Luf
3tDFzcbSWUCy75580fiME+LABANRc838MfwJVhVsLJE+mRPLBXctFaLjBRcnEmeL
JVRHfKy1jR6tUMKz+C3vpMxjrqWun2HKsuvyaHTF7gal9P1/dI/aHIvFN0qeBytT
SMVsAMTx43n6IuEr5pRebESiVktvfAFe/k6n7MJ5PWsq01z3GWUYW5Lb1dp3+WKu
CYTLCN0tVU2jC6bmijqGT3Amn2dk9MqbkvQUzGlGVA8ozpCaFWrqIIKLLBNFmyr5
J4JNoZOwUZY6G+8LDvEKpq4rR65ksYtx8I7XQ4z+/Z4I7ht8XJoJtFsxNWYnF4i4
kALSIuIN20C9WkRIUMVrW/g3Ct+lvyghEzMxm75O6o8Mcg6DGalV+fqfx8MS6QoM
8+A+3JiLCfAzHgDgBo2Q1jtNRE0ZliEPNVvkTHzWrSOqkIV7yaH3an/ePrkm2slk
7c2Oot8QaNwJyoGeEeE85T0n4Qu565lSYmeBQXlQd7vwgpanN/3YF6tB2VHLda8w
hCp1ehJ+ksE3WWRe87uvPHd9mwwpesENNsgemdGH+1gRfnOyCAxMKq4drIC+Air+
M5k5lIcJshIHUvgTkHMO3FwPkYI4cpI6mBmyntE98HFdS3MKqFd2A6nvlFcJdgE0
qC26dVbTqRMJSaUyb8ZT9fiHghgZEkW8fCItRN9Xxq2vK+KIrL2tFM6qHgkb+ydd
Z7j4moY4WHpaOQzZf8L2jabItkpTLvbollol88HO1xDHs02NAkI1vMZERY5bmWjn
b4f3KC67h6cN7/0LXuAYYzTEYFTeVgyOuzPf51cJI6IfQRMAV0y+HsmLeu9kmT9i
d9r09Cc3CdpNJTMjKGOLS+FrZwqZZQ7tUHKUFswECPyoqlZN/UYY4dRJVMAdWbXV
LQYp4M4MpCmO8oJhaeHogw==
`protect END_PROTECTED
