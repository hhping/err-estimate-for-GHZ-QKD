library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_tx_pcs_pma_interface is
    generic(
        enable_debug_info: string  := "true";
        bypass_pma_txelecidle: string  := "false";
        channel_operation_mode: string  := "tx_rx_pair_enabled";
        lpbk_en         : string  := "disable";
        master_clk_sel  : string  := "master_tx_pma_clk";
        pcie_sub_prot_mode_tx: string  := "other_prot_mode";
        pldif_datawidth_mode: string  := "pldif_data_10bit";
        pma_dw_tx       : string  := "pma_8b_tx";
        pma_if_dft_en   : string  := "dft_dis";
        pmagate_en      : string  := "pmagate_dis";
        prbs9_dwidth    : string  := "prbs9_64b";
        prbs_clken      : string  := "prbs_clk_dis";
        prbs_gen_pat    : string  := "prbs_gen_dis";
        prot_mode_tx    : string  := "disabled_prot_mode_tx";
        reconfig_settings: string  := "{}";
        silicon_rev     : string  := "20nm5es";
        sq_wave_num     : string  := "sq_wave_4";
        sqwgen_clken    : string  := "sqwgen_clk_dis";
        sup_mode        : string  := "user_mode";
        tx_dyn_polarity_inversion: string  := "tx_dyn_polinv_dis";
        tx_pma_data_sel : string  := "pld_dir";
        tx_static_polarity_inversion: string  := "tx_stat_polinv_dis";
        uhsif_cnt_step_filt_before_lock: string  := "uhsif_filt_stepsz_b4lock_4";
        uhsif_cnt_thresh_filt_after_lock_value: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        uhsif_cnt_thresh_filt_before_lock: string  := "uhsif_filt_cntthr_b4lock_16";
        uhsif_dcn_test_update_period: string  := "uhsif_dcn_test_period_4";
        uhsif_dcn_testmode_enable: string  := "uhsif_dcn_test_mode_disable";
        uhsif_dead_zone_count_thresh: string  := "uhsif_dzt_cnt_thr_4";
        uhsif_dead_zone_detection_enable: string  := "uhsif_dzt_enable";
        uhsif_dead_zone_obser_window: string  := "uhsif_dzt_obr_win_32";
        uhsif_dead_zone_skip_size: string  := "uhsif_dzt_skipsz_8";
        uhsif_delay_cell_index_sel: string  := "uhsif_index_internal";
        uhsif_delay_cell_margin: string  := "uhsif_dcn_margin_4";
        uhsif_delay_cell_static_index_value: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        uhsif_dft_dead_zone_control: string  := "uhsif_dft_dz_det_val_0";
        uhsif_dft_up_filt_control: string  := "uhsif_dft_up_val_0";
        uhsif_enable    : string  := "uhsif_disable";
        uhsif_lock_det_segsz_after_lock: string  := "uhsif_lkd_segsz_aflock_2048";
        uhsif_lock_det_segsz_before_lock: string  := "uhsif_lkd_segsz_b4lock_32";
        uhsif_lock_det_thresh_cnt_after_lock_value: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        uhsif_lock_det_thresh_cnt_before_lock_value: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        uhsif_lock_det_thresh_diff_after_lock_value: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        uhsif_lock_det_thresh_diff_before_lock_value: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1)
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        int_pmaif_10g_tx_clk_out: in     vl_logic;
        int_pmaif_10g_tx_pma_data: in     vl_logic_vector(63 downto 0);
        int_pmaif_10g_tx_pma_data_gate_val: in     vl_logic_vector(63 downto 0);
        int_pmaif_8g_pudr: in     vl_logic_vector(19 downto 0);
        int_pmaif_8g_tx_clk_out: in     vl_logic;
        int_pmaif_8g_tx_elec_idle: in     vl_logic;
        int_pmaif_g3_data_sel: in     vl_logic;
        int_pmaif_g3_pma_data_out: in     vl_logic_vector(31 downto 0);
        int_pmaif_g3_pma_tx_elec_idle: in     vl_logic;
        int_pmaif_pldif_pmaif_tx_pld_rst_n: in     vl_logic;
        int_pmaif_pldif_polinv_tx: in     vl_logic;
        int_pmaif_pldif_tx_data: in     vl_logic_vector(63 downto 0);
        int_pmaif_pldif_txelecidle: in     vl_logic;
        int_pmaif_pldif_txpma_rstb: in     vl_logic;
        int_pmaif_pldif_uhsif_scan_chain_in: in     vl_logic;
        int_pmaif_pldif_uhsif_tx_clk: in     vl_logic;
        int_pmaif_pldif_uhsif_tx_data: in     vl_logic_vector(63 downto 0);
        pma_tx_clkdiv_user: in     vl_logic;
        pma_tx_pma_clk  : in     vl_logic;
        refclk_dig      : in     vl_logic;
        refclk_dig_uhsif: in     vl_logic;
        scan_mode_n     : in     vl_logic;
        uhsif_scan_mode_n: in     vl_logic;
        uhsif_scan_shift_n: in     vl_logic;
        write_en        : in     vl_logic_vector(1 downto 0);
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        avmm_user_dataout: out    vl_logic_vector(15 downto 0);
        int_pmaif_10g_tx_pma_clk: out    vl_logic;
        int_pmaif_8g_txpma_local_clk: out    vl_logic;
        int_pmaif_pldif_tx_clkdiv: out    vl_logic;
        int_pmaif_pldif_tx_clkdiv_user: out    vl_logic;
        int_pmaif_pldif_uhsif_lock: out    vl_logic;
        int_pmaif_pldif_uhsif_scan_chain_out: out    vl_logic;
        int_pmaif_pldif_uhsif_tx_clk_out: out    vl_logic;
        int_tx_dft_obsrv_clk: out    vl_logic_vector(4 downto 0);
        pma_tx_elec_idle: out    vl_logic;
        pma_tx_pma_data : out    vl_logic_vector(63 downto 0);
        pma_txpma_rstb  : out    vl_logic;
        tx_pma_data_loopback: out    vl_logic_vector(63 downto 0);
        tx_pma_uhsif_data_loopback: out    vl_logic_vector(63 downto 0);
        tx_prbs_gen_test: out    vl_logic_vector(19 downto 0);
        uhsif_test_out_1: out    vl_logic_vector(19 downto 0);
        uhsif_test_out_2: out    vl_logic_vector(19 downto 0);
        uhsif_test_out_3: out    vl_logic_vector(19 downto 0);
        write_en_ack    : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of bypass_pma_txelecidle : constant is 1;
    attribute mti_svvh_generic_type of channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of master_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pcie_sub_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of pldif_datawidth_mode : constant is 1;
    attribute mti_svvh_generic_type of pma_dw_tx : constant is 1;
    attribute mti_svvh_generic_type of pma_if_dft_en : constant is 1;
    attribute mti_svvh_generic_type of pmagate_en : constant is 1;
    attribute mti_svvh_generic_type of prbs9_dwidth : constant is 1;
    attribute mti_svvh_generic_type of prbs_clken : constant is 1;
    attribute mti_svvh_generic_type of prbs_gen_pat : constant is 1;
    attribute mti_svvh_generic_type of prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sq_wave_num : constant is 1;
    attribute mti_svvh_generic_type of sqwgen_clken : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of tx_dyn_polarity_inversion : constant is 1;
    attribute mti_svvh_generic_type of tx_pma_data_sel : constant is 1;
    attribute mti_svvh_generic_type of tx_static_polarity_inversion : constant is 1;
    attribute mti_svvh_generic_type of uhsif_cnt_step_filt_before_lock : constant is 1;
    attribute mti_svvh_generic_type of uhsif_cnt_thresh_filt_after_lock_value : constant is 1;
    attribute mti_svvh_generic_type of uhsif_cnt_thresh_filt_before_lock : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dcn_test_update_period : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dcn_testmode_enable : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dead_zone_count_thresh : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dead_zone_detection_enable : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dead_zone_obser_window : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dead_zone_skip_size : constant is 1;
    attribute mti_svvh_generic_type of uhsif_delay_cell_index_sel : constant is 1;
    attribute mti_svvh_generic_type of uhsif_delay_cell_margin : constant is 1;
    attribute mti_svvh_generic_type of uhsif_delay_cell_static_index_value : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dft_dead_zone_control : constant is 1;
    attribute mti_svvh_generic_type of uhsif_dft_up_filt_control : constant is 1;
    attribute mti_svvh_generic_type of uhsif_enable : constant is 1;
    attribute mti_svvh_generic_type of uhsif_lock_det_segsz_after_lock : constant is 1;
    attribute mti_svvh_generic_type of uhsif_lock_det_segsz_before_lock : constant is 1;
    attribute mti_svvh_generic_type of uhsif_lock_det_thresh_cnt_after_lock_value : constant is 1;
    attribute mti_svvh_generic_type of uhsif_lock_det_thresh_cnt_before_lock_value : constant is 1;
    attribute mti_svvh_generic_type of uhsif_lock_det_thresh_diff_after_lock_value : constant is 1;
    attribute mti_svvh_generic_type of uhsif_lock_det_thresh_diff_before_lock_value : constant is 1;
end twentynm_hssi_tx_pcs_pma_interface;
