`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HfyeP+EfqcQluXgmGmCZrif40PhZHxd1XzMtDdSnqSUHUSuENP+tzj5EiHqgDprU
uG5P39xmIvQRQ01f2/CUoHmos5j3WA4FjE9irkz8Gyryk+YWG8HkBirOQDGwAkXz
GqqAuRUnUbkKkpjbawJlhVdEj6o8GhCYp/G+CTrsjRAgHNMXkI9G+YP5IKIuOs4W
rlPCQR3d/G7mPON4fshwA4Q9VQCGrg8C2u2sTeAJjvNLk/d2z6kwOZwhWEzMbXgk
yFx+TyRmPQVtYtFsBy3JYlWKLq86GWRIIGFoHH4Pe9aiZ1PqkzclFzhFKbjST3oR
agrUyPgJHtjnvPBb8E4sCk2iszlbVaqftk4aCL+tz4h2u8EIQdp4mhGh5Cae57uP
liN8D23Qog9F27C96grw+FapH3YF6QEsNGN4A1qRY3zjEHEsmT0CNcAHfSuAxbcx
RU2JJEfXOloCcQRIOTdDxgZR7O00x9WPZHbHGjySlMwidwdh937s4R82w0hD6/W9
Qt989eCZu7Ag3SsMkkRGmRUxcUjYUqaPPSFNyfFPVF5OQ7PNpDxor8YuOSI4zF4O
23em2kmNg5EMvAlUn2juj7h6SBbCQ+I3qbR8SLgleZW7kgMEuXx0/7Pcrt0fpcan
tMBmBAS/msCEutSeVhFrEXsQ0q9Lw6Ogkb3ZyvT2ayEuBj71SzaSt2N+mFBAJwu0
eauuYs0IynE0GqI9/uDQSkZE+wFcbj0AZckAvjBroX2deP5XAJg+g6ov5Q+irB9E
9ptGtQAYi71jfhMGJy3YdZLUBKIVgdP1F6HUZscAilEMW2+FJ31xhEjUt4qmsecG
fKA0esS7swOlz8ULCBgCUasc7uHjhV73oOtsVM0gqSsCiOYYpV6wDbiKwdGRXnc/
E54LfvdMoj9hgh32IOvkT11Hn52oXOfoYYjuXGHFSo7D/7DVwc0jRc7lBz7bWdoU
bOWQeza9dM6UdgZPG7Q5Wv174X+JZ8SeCVlehl6avUN/H+2IhMH+tMgrK5Cl4hmQ
moYfv8SbWMPYvLnWfJeQvZM2CCDCGEbJAFN2Cyt/ky4jUEYsrarpr9ILds2TAN7l
3/8Hc1K4zeInyiBg7vdaj438mTko+Eqlp9knBzjIHtqAVdq4rSLZLAbafuCgiR+G
Hf9QSMFZaejTabX4VFXVdXqLHa7nCcjrRpiUPfyn+dqFuzwUX9t8kOtLxUPr0fyO
IgAiY18kODtauyCLD0zam0p2x3+drtB0o6Zc7X2HIE81kQPl6HPM/GuXJsp+HWOX
7HwzFtN8++krl0QndLyEeO7n67bYVunTxyaCa3hWGFDpbwMo+J0fLVECSDugRnbQ
XA/0ZVzJRhSpunnNhnx/iMX3qd3h5xuJGVD1ufbfU+p4TRx6TS7XtRC2E20TWXRx
XaDyVF+rlVl5FzzENtd42Cp+rMgcYfaiHorpi0+1WNMgyJhNgg9JO4DhpILUqp9A
`protect END_PROTECTED
