`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWcBPiBa2ytSM253L3/otVUfKE2gdc8LiIduUpq1qXzNzWmXoWJEQkNiZEMzSar8
suvfkIJ4Ta9S0/vrvBqtwXXYJL41EJn109AOwjbIAPtzmbgZ7audZECUGMf6Mpu2
ElBft1zHFfpKvjlAFnrUNy3xyCyQx7zc1G9qBxqGzmSVRHVixl/zZFycspAqTZvl
AmHikWL+amycy0S4LPABOl+CPaBr790cO560Z4zzNZ2naygNs6PtWVosqkvI7Fns
AajrRpGXkknmetB1DHKDlNMxgzkGHuvyhFL1yrIFL27uNknW+QxEG0yTKGUoI/GI
Ezw9poKe033OKrpdAmb+2jtY2WIvf3YmxBFgwxAbd9EUvWZaXUlqHNXirEF/mFlx
`protect END_PROTECTED
