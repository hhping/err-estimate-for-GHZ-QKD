`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CnHqLCSkRU4OE6t2MktlrICNilfoM3SnJwIIUrodetr5VjS+8ctHJwUI+hELALg
dnu4u/7gPmJHtgSAykOGc9HBvXE3RHkdeBaZup0OUHp/zedNO5VuL7zNaDy8ZPGl
iiehpQqfO/jN14qtHaVUaIaEZy7ygq5gJUDcmSbsqp62NoGAunrh51EHnORk2AvN
QNjnhlA+ZJSnCr5h+EV+TINya57d6HSR95R7YlHGBE7I+dmd4i40eiOexy4AbUQ/
eZSpfpcYhCtylw3AguZku4Q7NTkg/ueHKZ6+xywfWeKHiLGaThIBZu7qsv1R6F+S
+RzENY3WkcvgATz86C3hksbrbwpJB611iu70tTqiKphZ8iLLzHTk8Hpwr/b1txOf
AHk2+zGqgAcnDO4NM7nkPap5Y5oLdnIQP+8oD3l6oNHeIrW9qZCV/1rDyi859p1g
HsN5I5BLsY7WmRiPwTEqzlNk5uws1wopeLmhHRyZXj7yGWHknY9nZzOrsgS2bUdG
XxtrDeIEYe4DJ0qKHkAZx2UdEVz5CNl/RoQDDnRr7fJRzh8hL5SLe2RAWq2Y06IP
Mhinci1975SQ8BDhs2q8XPzXHcXBe75580rLyA1n6Mlk21cPZvTI1oeYDc01q2Qr
whBcMhIgYpqjYw98WhXYUUU5HcBzyfvZOwTD0Q3m3HYKrKbkc+2klD7SQ5FIc66M
czWh3sv9Bq+T6e+AGbLuum7Ibi4ur4b+XpHCUyCWsPhwmeORQeJEZnBqZAdz72Lk
W1PZDe58a3do5avfLytOx/RTv+Y2Fw7h+G4ScB/jTy36lTecmaondC8OqNS2EM8n
kRhK29sXdDNJIhjoN/SvVw3qBQ9NLBFL2M8GNwQkzFY1CRhBvYmdqKJSkX5Vfzlf
c8ES2vKloEYZqJOcSINvijXD8BrHoGE9Ij62Cf8Ea+i5JVgbmEOp8mLwzMo9pmxX
4ogATyGMkCkxEdy1LzsNQdNW0dvwBuwAMPavuHbhn2r+ljmKYjksTi6Vppx9XVSP
yK+bGWSmaxH019JgaNGWjCLsDaVJfhIdH37OzV+rZg7cbW5EdbTYhFqX4WYQteJX
1U7PI+D5RBoF9QTz2dKC0TcbG4egvUwKZXRMEiZMZtVysVW1pv1NLiIezfVUDcVm
EO94guh7snt79bUsnsOZknH8kqwSJHVJDiip0epKmF3bG9dtxPyMxybLCV0XnVK5
pHPub+sUrUf0yEHJUkHB7gnoLhJxSB1tKwDUg8TwS8oz53VIvv/RqZ/Uj0LERVGL
3N6WtOS66oCRhBWdlSo8Oa+kdj/mTyBvM0JggazFe0xVZeCw5e2UBUEFiomZo9Wy
C5KuMufPy0Ve5l2M77WbDyIE8RD1W5+V/XXkiOP+LV1hfYeUw9ACvvO4089zZRdS
51w/tJHY0RoDIEk3f+AEhfmLttzr52cc6PgUyfDmzV4nfwgyBurwKRs68PQpcUiF
jy/VnMZn4MuruCqAott+hIK0LQmUOY3/kjxMPm3DGrD72y7fp7XqEVBVrPUn79UV
Xq46zUiWZNU5jP4E7rm3TN8iA+esker1qpfUzeqepz0DK8cIdW5k1SqyYWxsT5cq
gU1aV3euyeAbxU/5+liUopvhbeeeuqzOnCRRgdXIaImhfI3aiwp3P156UBwU9glT
Br0jTVoyMmf5bflyoAFr7c/GafN1rFbDPPuiTQEsmD2wTI+lmeoFYQsUOKiPEG6X
TUVugrf2Dkd4Y7asL+PHcHmQxTWwq9YZq9/Ybu41AyxMB6MFtjGndFvu4CELxSX4
iKnmADreM8nfp15tANDHTGtNOtunb5mDXPhT9gPdQuu5tAj52OHYzzvLgQErZis/
ifcVbRVktsKhlqFiUXG/6OgeYjYvClnPcIwZvTNnlb7a8qSxHyZp6RXSdoSpsZZS
Tj+JhZSGtiv7IiqMD7+xEZsd1sFpij5E4A9oBXYUC9LHKrrUa3YTuwTrQDM8WQu3
+1LsZABbQX28HdWueB0DlsDs1CDTy7rQY/bBTda+BP/9p7bCn6xqZrLiPS/BtDRw
1BqJlQ/rY+um+STWbPpjRJDoAgt+T9MPxcfiwAuC/EqMaaRf6rdD0RqB35RrE0n4
LrPT2fIBzy3Rgsx8HdtYbLylqnrjIR3Au8kTAlvDwyMMgDFtoyx7jzZGC+AL5XMB
asl4h7wXWuMvEKAQu+VXhxx+dms348U0IXDZAcqSgwhUnEH9HC+4sRcOHzKsr09m
MGTTfHkB8i+RT8m/7at33AG+vkUNgcOEdv+l9PN1lKmqJ38oczhUc0n3xcTl+0IL
kI5wA8XtwUbMmtYBMnbULnTNYgnHb++md2dzm+D2X1Zhs7ykTOElpT11XkzekzvI
e2uuZhcJpglmmVT+Ps6ox6rNyXxkCtjR9UV9rmYzG0h3f+iAWlcDqO6Kr3tyMKg1
xK5zvY9klFb9jBbzE3sE7N2Wh5Yd7PWUg5ShKMSpzDLytZfTTOQub56LRcIRv2m8
eeQQfdsOFolmNb1O7QdyWMGkdR2qASU3CmBS2xTJ3YS1NzL8gUSr28tdloDUKZke
`protect END_PROTECTED
