`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RlLsWj58HKEIVgy4heeU+ZzdNVVIOgk2+BWFHqeJ2hYcIJIQwF2bg4YHeWiebyQU
o/U/BA+wxm3xtPWd/y087AGxk8yz7d+NTdUxZr2WbH2k7iAWFuc90662Ltj6jKXh
AZNL39SdJR7kyxxG13gYc7R8V9j1dOLmTL86PK1TbdBQrdrxw/Z2iDSs2dc2kqVS
VjQDp2xEw+2rpw342WSbk7kWjtzHywIJ4GVGcrQ3ykSUNhnuVD+Dn/xYZGOGgtHo
dcNW7xT9lIrx0SOaeSc8fpUunv9M2g3N8JT9R3D6kKGAUfh2QW+gFAsC201xLRyM
abappHJOlfaZw/j+jc+fQ/WDDbLYzS54EOkWIh6L8XAi8eDYPEhYMrlHvPQZrpZ9
IIET9HkCgd1zhFzuwPgQquJ/dOvTIMI853ujfa0CTF6JBHK4DAxZietkmPry+Aqj
SJ9GRE/Rz4gIjBsmhprwIn8DZbxDegXhGOfdABfT1MhOAAQyBRWVoDyl9T94uIU1
/vMbfyk3AufUZ4ZdJbgi5yxDaDr4Q926Y5Zo62q+Pgg/rKp/b7jGhNw9T+9xGVFH
qLnsw2sFez392av/aIFT4xpnVB/dI4XyhXh3aeFAxZWTqTPSz6ZGkSjZb7yMpqb2
53VLJLbaVXb+rKxcPWhZIS52K25h21DVy8PRfC3Cy+SOt4L+4LLc7djHXFWwyL0k
eDqyYH7JWdDh7Z5shi0vJnMB3JlfWxZn+TbXS72j+Yo=
`protect END_PROTECTED
