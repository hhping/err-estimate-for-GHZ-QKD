`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YKVJB8Q5QWYmB6ERtOWwb1Ws82RhmvMDHO+avHxPGVZaL4pmyZZRmTeioZ5V45Ot
Zfri3BEGwRiGYztwNHUQ+LS7pd80OiaSSkRpoWZ+xekoxx5RPBc19v+G7nHe5nGc
3zM3jkhBMOcNQrQfkLJpD5F2zYJ2AA7MSN4RMbn/r8L5X+OWd9mDeyegOV72EJ7u
sJnb9xn8CGx1rcFR4jZP5M3Jvsgby520acElE4aWBfyK5n4B6ixSCY7f2UOr5XxH
eAFaZ+bHCtIzMbIOwOdJzIkDVVp1ewXIh+weFaTkrWICsZxc74glLnqDRM/fdNbB
fSb5mDrEOxZQO+LAShfGDiziehyQDMGbuA/EtKBG5Hw7eyZ5j44wPoYKiVME/tJh
mNdNsViY+YekQBJHDwYEuDKUJB1gPuASdiCCCm3M1tq5/q8PVKfcQTFndwvF5GIW
Pn2RVE4IhEw5jutmvYsCdKmDTQMBerOdJqV5zWllOMkEU/iDKMkMpDeUJEZqxgOs
hwd/BVgEig6xDB5rpfnUIeiNytOzM60A8TWAXNXzFP4raP6GmsT9AYXuDOY1rh/P
OgF/qMAdj+cJPqZwZszbksYhRJCCU3oJgUy976cUSX7r9QQC0xDCVe/Of+rUvIDQ
xmFLuQkXVrerHqK6dL2lu1mleM0Pch5tkzxRu2qQTx2lUXtLT89yXNt55n/jy3Ob
+q9kkiZrsEh0POALmZ4BXySdPZySK+WTE9Nd5mgcWmRwxWijzJr6/yIPxJeOCV3j
oIlA3AkfWuiAMgkx2+KU2vSP0M7bvJFLZKcYMBnWpbkk2XwbewA0ErcVAxkCutYX
qpQpE2K6LdfcvRr/vvY2o10BKxbbdBIk3ILZ8U7YiIPUNpp5UXfUeHFo/W4gF3+I
42NAv6rrIaOvoL3dLDBD9lmKiSdpVJDFpYLaNwE4DkYXnAwLJFIRSglirKWayHhP
9iRWmic3ewhO9/rEy0LdkMQMkkXTzbCnsmpNni4ctn70FK0Dz0fQy9JPI+5JN2Ut
EiDg7dHX17SecPBNIvjWOJu+LT3xBAimrk6h/Q6TFfzblPc4wY8UPwVUMFTdIge6
/EArL6WBg0CXKe8strc2gjJFZj4qGVTBkNSh2qwr5mI+2BZasUkAv5xoPADcL8fJ
2JqZ4R4vLRMmV21rCRvfgDj9lK2socMN8Rgmm4pWwli2ImQiqpVTfnSwp+iWl0zz
ADi3L7leiafnRDYDB73awwQwzWZLZn0JToQANkGNo+hTgSlbzYkmxXZaKwDOZA8c
iTI8JSOjj+ry5NmV8P0s+IXXRRYdPcAPpp9/MGBKcrgYW3J8Taa4nWvOTlu9cKl/
uqddOjQUHBp76zR9VButbZ7c4sDugaiUXXA+kY0Uir4NNCrHZGA6MWdwCgdtEvGR
1ZW8MnmWVpSX282/7ojvltmMUKZBIv37ipYAEbRIiClJrkFulZrS9ZUbK8KYZC1W
DcL5T7Lq6qjMvOQsQHpAFpVE/mViCHUUgJb25CMyp8k=
`protect END_PROTECTED
