`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbdAvdo25rzT/w+cyXfvrCXfpwQy/c/ZCgpBiQLUr4xy+rI5r9bkD2XCx60dApoj
6GN/71stPttQD1MhVoOvmzWiAEXCgA2HE3KF+G3saJgjOoaYtffeW0ifuOEez7Da
RqwWyafZO9XhlBlfZv4kvObEAXWfbNjpfycIK/dnIMGRBGQOFnHy7bo4TJMpWqzK
M4XPJUoxooIJdHtixQcmxPHALmH2VNKugWfyj4ct8oYBqGDlJ1nM+ADtjDZRfsuy
yjqcc9YqimY8PGN1Ad04Q5oaRvSpK9BAEV7rWHjhhevRj8fmNI+ceAKQiMm3saX3
bBJiRyC/gT96fRt+SOhWjlQu4GeYVv32uXJ5JbruRs5PKCRwAIrCG5a/JuyRANf/
jBF+zKC+bNExD8bGQNinDqqPr3HyzYRFnz8VfwkNHhaBf2OYJ/jmETQ3rnHZrF0n
WbyF5rUuCDs2W50mNc533pUIG55HqoQ+iGYmr26bxuuSQW2C5Z2GbHu+stoCrTwg
Cakr1NMjGuqHLqKAwU16Q0/qP1ZhBBRbnIWmPE1744yjlL6XBuKZo08T+gdufJk5
br621snIc1SLyZsDqBeUVXqseWHI3yGI4Ow0nC/R5zkrb4rPsRqoX2UcJdbAr/fB
joOJU/+VmxnFqxG/xDe+cWrrvfDzBPjBX52l7XBZ01DXVCnT2s84s847JR22RGGb
CWna8bDIR5i3bhKUq3tVqPVv/O5+8FN14PjDakVvdRf+mLU8RljC02xP2NJ/8nXh
n3FaAXS8oVZI7zFTxmFq53a9zifGvTZjz60M7V7u+ozqUfwn2xcDZF4LkRQHQ+JT
QVI8K6cUYuKiZ2NDANWCgmJC30XFQktqOK/7kKZ42Kl+WF7rrRWF+X0PUAj65CRT
Bwwf/Dx63wDZHrHjfLxDcsl0sYSXfGDr+Urtbx+yBwO7oG0P7RfgxiIpZFS8/xpi
xuvVzXP0Dp/WY48nIkk3mp/y00jwBI3zdftRwIVqvGj9iOOAhcX8VIkkhDgQxACn
aNKmEk6QdSYu29SD1eFgxaJXIpL4Jibq48ASv6k6BBwCrdcq057HWSDcv66cmk+8
loQERk2Ocpt7MXi7jvgJgqNeTIiEgaWLDBMbAlTui8tW8c1Q3LOGbk/nblvPnTca
VHGwRetEfut0gEKCjGoBB9AYXzn9crCnzeDLrQCH7niVR585WnA1BFX186xqm7oL
/lNfyCMtXOZT6iq3YTGDnOEJ61m15KZW/MItmFDDYl1+jr9Ii8ZtVjc5MUc44Chj
No2sHXceIuk/n1+yr7oQT3iRUDoASoLuFuiBDELYYMxC9id5apSdJeoRBFIBDScr
N779x7AjkOvCR8QOg24GcyMDKZi9Bd4AuVJaB2R15UzxfQLm6BF5vW4mu3fCjTJ1
f4PwOhaIJ9Gb3KnkIj4iY0k50YZZ/KaN/imSCo3WEUdBoUOjNHJbm+GRekbMPHBL
Vv9t3s4wsTnLO2D2ECvRDjmfjvHl0fdga7qkUnDeNMbZ94aisk+/efR1H2aKtxnR
dGcnYfLfvWmgwbHnonplabqqUckku+znYz8aBizi7uQ=
`protect END_PROTECTED
