`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NazRXf3wjsuGc8Oskx/mLySpRxNJEzFwF4JNjMyxG1lVZYgn+dXuKuzuITNj0A5S
DO0/TIufw2UTvaNf2prO9lksLuZpFdEtYqZKhf76ZKIpNEUb6x4L94002ZO19N+/
4GR/kjvHEgnCYH0pdr+64n4ifViEjUQTze0WZzN6IGq5PMAxrlVo9Z1xYvGo5I4J
8LHICnN7Ny8rf0ESNZ9n0+T++Ppmys7icaNe2jOwd7v2O3PiiR+pD5qjQj08oRnS
B3ySxfJFdjeQGpDMiKcuq7Cu0F0mnBY7XMHbY1nVS7z2g/ad1rmfLeAfCtqUtnZ5
skqQyvINdn/CXQ8GJpKeq4om9m/Q6J1fewLX295hJn3YTc7e3DvFNXV/SI8WiCyH
mI1UB8p5GRd3rq1e22/emNkE+tRJs/Mkt//BQXjMw9G9JVvtfiliL0hBneEoatfX
WovAaOK2EhpVCUc76/67WfQKjx/xiGE49uN/dh+lqLSgmKOWDKIS9MplW0qNTkHX
3O3jQhx6nmp3jGjWS5gJPiaiYG7h7UYJZvNSDjdxdYqC6c2gPB/vg9CjmwXohpEm
ZtVO09Jt5v4uEfux9JKpGI3TlVQsm7HD6d9atNM2IPUQWTEjhqZBfkXiEsVyAE1M
kaAcqlv1kTjon0suNED0RSH2wKHSeMfjrRqL/E8hHWKxZjGg8/IPF8hpsxNktTCQ
CVorGXzW7N7xM5xXNn2iKrdObxzCSoQRG2V+Aa6L/THIfoCPBMz0l4eYWRKvtOwP
vaAnLRMoy+9Amb6rtO6w4NKd2LjaGczsAc3UTge9T/1gQ98CR4vxtUypBREt1ISK
AF/QGkaFsRRNZDHJ2zznSTP86mqQesrlgcM0uRjSOakMKk09xdgvTIPbciB8d/Iw
I+I18QrIh7vBXHJfDx3cXdzsO8c5fFKdiUzf3CzJHfjXHfxpIH8+Ik8SJEntC94J
rV9HH5TGwi8tkT+qoNAJZJY5TcRJ5pFHCEW4Et+mvEu8hLAdrAE6uFChy4GMON1e
TgCif///8i/icMBCDZ7fh4eoZlkjH77sKU7WNCPa7ks=
`protect END_PROTECTED
