`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQiBLogoC5ycFFI519nXPfCdBKAmeFCrfou0xkEkYAcbTBbcViuZtHDSvThihBmt
otlLmJ0dpma5fSQuV810L4UE81Kur8aI2iGZtK/vq1yP4XaMis/YBIGLke4+Zkcx
xtYWORNGoY80uOdY+qRet7Q6zMkGOqpFECwzO8EgcjU3ymJqtNYRXSmjyKbzJfwP
2oYQShWz8mkEQ0h3nzmfsrJyzGtOA2JWb8T8yGEjMU0XLbBO6EmdaIfQlafVrRJ+
pNLO8ovKUbY/KZPsy2vun+FHK50ZD3Rm5h9NlOZP13Ucb9hxP5N6i/OPwQa2Z8kF
srErsSJpWBydYIfffFcko1bO7vxbXui0rMtVkcDtCkTh6BV0E+WYbK2CbK93lNF/
twWAsx6gYlaYVBWELTIeMu9MerRUiOot1a0oAS6mG9njE8DMjHH/mF6xhp0oJct2
0hdbDNeifUgGPNXSpneQTUXM5E8puzKTfTfrh3HzGvatk/kgTnioszO1nXu4VQFB
ZtPLqdUHnR4PegkuvwGEo/9+DFNNzo2V+V15LxefA1OX6ucdrEiM/bHwLIG8Bw15
NzHEdFThH/uMKPOzxe46l28BljfNJFL1uCW5vOOxOiA8U79oKgBX9caHb4gfZSoF
YQ+TUFQhAEa1PjANj6lV8dVJJoPGHB1MhZMQ/ywzgXpG7NDn9xbVNyiW3PIkFXWT
ZExg+ZieIzg0Nxwu8tRdl3sqahg+yURZ2zDy63oZNP2LgFill0+MmG9PvsNqFMpL
HDnYtS2MqUKEQxdl28ZtxD0c8YHLW1CDIODXZVg1QMZ/DFhVHJKBIgUCQ26gw6bN
6O2fnxeezJYnR+sjABwNNGG5Zbd91/b/5SAap18CJcadW6QPxi520uolzwYJG0am
xZcM1etGDc6rVysZAnFQNVVPhy996HnvoleIA96ln1uUZNZkMwiKOhfEGNqP9PG7
letwaxaRYeLuTbW0wYt1juIA/V1KgPpSeyy+KVE6Qi4z25YvN3XedbPQriIU2nap
JLMSGkYefocZ2J30UrHlucxgohQfzXRoDCsf3xMfqIKTLFKqY1RAImowvnaB+DIE
h2eg0iSPX4Ts76hVxcgTHjdCPy0lL164vUGzzuTZiy2jqmi6utUHA4GYQiLsSFEQ
zeqwSl1P83hpkrztLSCTVaQXIYbvQqTR69aG0aeTcVb2s9pE/Xikr9OQjfII4Sz4
7ckLBe/oxbuMDjk+CpDEUhfZDLcEIa4h4Aw6p3j+gB7/4lZ8mSlVyeI4yzwr9MUz
XtzRrdYl2AsE4FytfoU4pt76mvOvrYZdFWrmObSG8wO3yY7a/BNmjXOnBOSRPIgi
fQWmQjR6tH/TX0Eyw/ajK7HKP1NL0LCv9g3HD7Xd1wfNfGsorBFoSH8hcfOT+wDS
u/24rxkL/F404T68KmJZ5NAZA/9wvLqdQy3VskeV0thmjWglm/U4iKLAd/ttx9K6
hEtcoeafsO72U6VpInXdepCU5DGPctoXYqX8UNuh347RP6kJ9Kk9/RQ4cGENB09q
pmhbKHNnIc1EIMGOXblHjL0eoVXw/O42UTuX2DEuvVMln/1WU6cYzn1CTe5pwlUd
VIk72g9QNYk5ZzBhtLyPiKFDQM2w/Ff6SVOB9Vz2oVXNTFMlh0M1i/GpMbLMq8kg
SHnECFY7OIpAzaPFwIT8X6xoZppFaGiLw49hoYkXftfq5FonH6rKVn4kHgX7Aqv3
85svDPx73JPIpI+myWcWb6NeQ7L+RCw3+8baRYK6SnCPAWhltNZ2FIGbpYabQjQc
/6EEqyXak62/GBzMj+2E8oAc435Giy58VjBAsS+SRfbJiZsi3Y+wenDiX7xsRI3P
RBCGaxIrJ4anE6q0grvHD3fe/ovEBraocWPFzbPgxQXbhsSlAngtsmHXOtdiXJ4N
AxeQ7Pu7UO26C8dA8Kqm/8R5Z3Idzgd+IkOKHVhslEL71h2Olla7Ghkq+pDKoV+W
gat0oY9OAJ9zDNwuj3Qd961vj0uhP6hv/rb3X9WtBnEf5jzzQapkgPIxk3ghU1SH
TwbfUAE9IfrJwsOMidCRKADMo3Gn95wdutTrR3szGw8FylLmPqYLIvDyOP0pFNwF
ugZrMB/aa4cCGKZ9UP7ON38/dkGpPVGfWh3JiU8I8Iy43PuZKth/eQ8ROeAkygpo
TFRQOEMPgE2z5IDZCWrucd0y+57+Pc/3BlG8qXsCz0pmbVSCMkmU3OuN0O52rU/s
ksA1D6kYLmLYVLXnUSBwDRebS2up5ucELlbq6Hze0iTsWTQIqWsH2cXgBRSYcUWy
qs1nCR6/n2c/reWEwVlkksCN89L5neizJVxxYQTEwRP/lUxpwGrVn7RqveH0AJ/a
qRZdgVlwG8gQyV2nXoc+YPh99IJxR48dBCwoj9gxlbwho9CXe7sxIIKBCf6X8gIH
8zXI5QOZ7aLPZRKmn0/BXApcA5xuIc74W/D+7NyK865nN5s2Sdv4s7VLDyaswc2r
Wse4ZDv7d2zaQSnR0EEOfjLOVSnxdvjPMjkXcrpmPtgkEzqhpEtcupYNU67LZZm/
IEtqe2goiV77hJYFMQC12HoqNCEoeO/bzd5Td+mmGYYtpPPChezq5JjqnqkQIUOk
pGNKYksj8uT5NsX0A+n4osJ69vkBkPDPu2QRLlX3iLgKVR/YOiqARnFKIkN5B0d/
36HTvbI2aTOdYoYJlDc7x1bCeJDfTjhyQo+VK4IAKVOK2VBaEulH59mb5og5PKBy
JWOrIWdGqGJbUnQrHFke6ZR5gsk3wlyebNs4zRObBPjDeAwMWMo/A0HhoA8vB9iW
7tTuJd+qOGwD99n4eUJXRUyklyFi2XZ+GYYgj6TSQy8B690wzXWI25S9Z3n8MLbX
rM8NP8+vT3fURLNOfefFI7uqUojpN5+TeWN+ObGLzCJ5F0BZBaPIzetbfxIqtbmV
ImaxavXc33sGrCYB4L0dKA93qEgcYTTA2yA1Rbyc0Tes8XqWdEF62I3BeBkGfDoC
lGWEoD6Q6+WtA5m4BQ0UAyZDPTPRIWwGqxlOEXWKUQRcbup3ITBOgALT76/tuyZP
y6ulWnPb4DnjJKP6z/wraPzoWbh93BnN+GjfH0GBucx3alSa4LInkq0Ho5Pesbwz
Pp4EJUoxDuAB8hYJde592RCSKd7KwQkb+QjpgbSeLyESNgPmZxf7EOxwPKyI+dwF
sSX4L7+NXfJm1ORcEC55JZkhpLG97qOeB2GQVhq/DgnL+A0MT1h3tUq9rR7xIvfb
uwo5QrLPH5dWW8dU/zCfBACTIGdO3uQE2K1rRnQypEE9Twm9fuY+7hesQ4F35cQg
vkbRQ5lgtYAphAN8XgxV7LRlDiwPtxqpumrrB+YUZ0lNF7JJEardgf+SOB1zqfeK
S/HkKswYu+WPRUHY+KjOV4hnFWqxwq2BGGvXKIWj29quBSCrjwymZFB+vtIVNxco
pzPBWWjiukkptLbBFJrcYPobP/SRcpV0WMHqtnWT+OHh03SGqt+uoNCe3yDas5f4
WeLlUorRPSsd18DdhsB9XUqwXlwRuZAXztqKWQhAUFilVaRkP+2QSNojuI9XZQJa
/OCqJIHca2It1SvHiXRNVAxZCmWA1fyTYINIGpkvTwwCRXebX9dMX7fLtAZ0K65H
BNyQCUpU4/XEwnjeq/ageJKsPLvbLEZITbpTjYopekDhh4ieHM6sGZLhcZkRKxwh
1vGX/lfy0Gr9xs/PFrFHGiMOS+qxWKwwCyrr/Ww5ipgNkNRLnuSKb7gfrEQcdBd2
qK6Lscj8dA1/oKYsOVlXEy2TAuo7c9XROtrq3zJLD+rItcyZd7RspvhCv0lD+xvv
jUGu7TVsylMqv6kh+/YqZx+AVfGuIqNXLvttApRg3nzSPmedHzxKYZcPkqIq3XuT
oO5U0/sc9ZjW0FgGN+veefgbqPFMCAPXYrvD+8ltX93Yr2VBOrVH0crdkSTDaQ3s
VwRwNKxhtAzlVOJhZvdAViomn5gBCQctQ7/6CT5X1cLUfITEp3MN9Jx4kMqSF82w
6IxbV41Wm11PqHzAETt4rTjjZ/s1hHQufC8cIJKbHId8M4Xqq8rkBayrVtSw/9Nb
bymp5dp22BAv/KhE/TR0PCxFbJUTaQ9XMw+BF2gplN+jGTHPLtMTedabmwD+NyL1
E3AbgRPMkidf9LgKIBR5gXG8Dcj/wzwrIe21L6QxTWdS4h4AYrpCXKDHwnn07EvF
e9Gm6LOSwkYkEZCQZBx7RZU9vW9/OAyrfzCU8agzZ3Jf33IhrIstzlmTWvHyaHxg
7Yjs5KC9wNmmDaaA2I+lylFBnyXmhVqNFJUt49kMNXWCm96z2IBOO0j4pw5X2iZx
p3CWsTKEa4G3T5TriLboZWNxz0naTZlPTvF42CBV1XcjCmW1pQe8rGVsFo+WxbZK
rO5P1pQaB7k7gqVbFSlSFLCAWOiulpo1Cq8VKCoG3zFZZazk6UHMaY8xoZx8cSh5
2qRtKJbu6MJQYYFiulwVHianJbQuj7zj/dwYoulW0lYJXYp/k5i7U4qA+qbZy+ez
g1Qw/voIBe7Q0aPY37nfFTFVzXencAiGJvYeAz8TqJ//Jbl1vHwJpGl/jZwzrhGY
OS6xMK3cVSPHpcvoqcRupVUyE0riiXGKtU9+xL5vgsT34KTWovKuWlOwmUJO2gqm
CEalHU1XyTtBY1BJA1NMon78TxSYEBDUeAu0zePCbVaG90BjBO4ciDqJy1jnlRCu
ma3Z7g1oJ7aDVnoECpr6pX346OwRfhwLzf074SkCsKX/pQ5VRXIC88DzKh+Mrir+
ia+qWHl50E+vApkGrkrp8i5UWbkR95yFmZEhdjYjaGfOQ0UY/6mqVACydelYyG/y
JAl3bIvK/lRTAQ07zMOCaagl95abxWJGXxdpZ+kGjghLMSLdi2b5dktBQGZDOjwx
CUwTwAbrb222AwzFydUIo+VLBZzRXEGdupkcJA0kDY9x0ek1IQK01QnbmlIadjNd
+jomNo8PPWilaPtAXe1M0MoMDQu7LcycFmQJ5FO5cvokNN5IYExJBuASuN9uzwf1
FpgEzWWEXikAWPYC6/bMSmb6G9FJ33RUd4YHA5UMtDS/QVLfQSs0gfD6TZYqlq1G
78IGh/33TLTcmCASj3IecpkTDxLCVNJVQTWzvnSrOQuvId4P2BEuSqcQux77wXl3
r2Rl2jMlCeUW0BFHjktANq2rtN+ulZZzRHPPJpk1WgjoS1LT3pJkY1ZeAD+sAs7F
duu+dgcknwouT3IqCIQMHzk/jUhb0YeVI+R9l4EE1MLAdNVFC2H316PPJv3Uvbmw
7zNRLPJ0JvOFRivh226B9nM32n/Kw5hqpjycHnaPJDCEu0hIgMr9CaXClYL3JksM
iY/VCNOaPn8bFCZ2uc5Va1X6e4uCozjO6zM/W5Pbgb/wP5LBWm8liNX/D+OgpUni
0ZCfVJUSOSG5YaIUBXw6BlJafGp1yXjg+EgDA8bXsbWiSaemJPkPP9Aq54gmQdrb
zK4NbJN/T5o4YI46GTsvVebphsJvrRoN2ymopm4PQSmIFyKWsC0GCH4Xo6c4CekZ
HQMLBGDMhOvf4Nos73uRXXAVzh//Y7QPJ0Zy1D9Xa+I4+E7YJmLSmM9aFyPMdkk7
4ncpaVwZlHPc6hfIslp27dGOXdRCg6DbHjUeZuI6o03Wm5C8Iiyr3Zmi8l6Aztuf
vm720FIPOM1i7fUSvF5FlOBU8M7LsEEiRsjKjMeo37fqhx0617Uh5OO54nMqE/2H
YH5yHm7D2F0jR16TgL/bKOkpBQD3P6glqFwCRVh5Iq4lV026qu3rnzgdA5kjxoG8
VQR6u+FyEjBE69KszjDse2KIAuWEM3PKtYPbwxoQRcCFOSvTacXzQnpnC40xpxfV
vtNTJo1wZNjDFOcvMTUv720bVrqnzRrP4m7ygYAdGk4vBtrMapuV6QvzZXKq+5Nu
rWzqN5EaWdYFn1GlrQ1+gBBZXE5hz1IhLoV5W/+FpruDqr0r53lZqh7ecTn/gF21
5GS66PFDFbFofWSoS1nh0cX5pzXnDHMGaoFZs4BpFNK6d2vQq/0m7nJrItve5JEU
KGKkBMY8JRB4gfH/GtEt9ow3pZpZVRUNeojZKDwqNimK1/0acTZRtPzA5L/9udyQ
0sG/YqEY4Vx7fi3LJi/JFPMg4/Gih2TRumWSFJmU0NjdvHq1BsVCGz/2A2N0oVE4
A+5FSP+iKF9Iy5ZIjkY5HR7GyBzWWKGwgy84QxJqEsivxt1TGu62eTZiYl58ehY9
dozyg4G7WDkdMtTSIoCxHswhhedntmTNcN8/3SBep92o7LkSkQL9/y3eZeA+sV00
M5d1naDcC/pKvgkYaknIljuDz7Oh4Q6x4VaV/9VVfAQuMBxiAE+q4fE/RFg01cIU
FTz83ki+UavHkJULg8sab/tk1CdR3487886dhUr28TEZ/i9/P7VywndotqbEOUra
xDp44suLPNXnZUYj/nAuJegZOF/zkGJJ0gQ+JF5fDuxcfyi/4Eq5Bph+t2RFyfXS
B7cogHnzVI/8ufYIp7V9znZNVNmZbn22d2jSOZ3/0GdfBDSdYV/12si6Q2j2F5DE
IfWuh4G4CENbvjxIe4Vah/iGhRIYAQ3RKei0ZixZCzNWaLs/y32WnKdMQ2BcMshb
DjC/0ucrTqdZxO0FTtO7uFlvk29tM5plnh5Xhej97fvPC+nhwKFWgRFtDMEDwsxa
TtIWHj1ORooumdKYPCNt76n2LqoE7l/Uv6w+E1iJW68dtqwxSpmmL+gn01ycIuVx
jK/ax9WhfgB4/qr4FoJKc/NqV/KrSJdCm3P/yzgWjFJmHrxfE3uQuHSCryIGqSE5
y50eUzDs3utI8+fhahI2/Sm9+t1pnwp8jeaJYJjAirHgcME2ucEa8UYyz4EFflJo
3TU1krF8rtbBX9DtCbbCdyQ2vG0AJXSJK+Lh8bWfAe9wztK9c0nj6XnsLqGQTSOv
EZUT6jILESxiemyzOml4OS5INP3BhPLSHPRPBtbufHX4yX4p65KiRSCvsSS85JMD
pWzA4nlwgBz4bobdEQ7fd2zuUwYU7mmuCaOMd4plPIkPt5pViqzkecJOO2wpXvFs
WzqyVW1FGdxb/EWHoBxrbpTz08HPH+Tt7Y8z37pSRijoyDF1IbclnuHAqiqTDwTk
zQVPxp+5Ky6WBB055LphrywbGL5Z1TokqHZqGAaVbt8KjaK6B3+rWv8mmkVVy219
b0185TeUHpBPvT6q+pSEXblByWXY3NwEYe8pBGmMPuz60SZlyV7Tmbmiur02BijG
iG4jp/nbj9u9huUzkhEdNkFyAOxgiRkcmZCUNUrok7PYrjLCnMiXNIrLUnTe8bJT
DqDCmvLpvQbZPtu2u0F5OgV7pJUWLd4VKRzFXtHwpUXzgY3+yhQyKm9ewzh5Bv19
dL662ZcjUp8ucMG8sjvuzwH50cqft0Lth3FYdj5tC2JcNYqE7Meupyw1TZJIPFLc
MAl6x+qzyiB/u8K8fuakty+HgMxFlfc18xwCK4vonSE5F9PEFwCuJXH+HRII2b0y
88gUDwcG9A+QCkYFtylhACk1UPkCN9YVjwablsyS8J9Vy8tQmixVam61qpiV4/ZL
ipqz3UXWWb2gQ7sBobwXfoPsFrIh6yQdGDWvwfj/gsPBU5XQHXtO9ugW5mCsiqQH
zSPDhgJNUTym8JYNCbhZBqtYu310mAWlkGlsL6mkYagtP3ImPg03rQkw5DbcL8pD
/FP69hTFScsWDMQnAnSWamZJ7pVbJYsVNNIYWcAQlEcg/8v9D9/TKt5j3AbG+hsr
nQT5V7c1nPfdObtp1OXFYBItQ2vZKhleb8PuZ0c7BHcJ8o2eiA3iekK6D7Ua0Fgs
NpdUgd5hDT4sAPBW1TjOirw5mquf8yispG+Tils+PGSmR7K/+VTvPN7D99nn8+aR
FQISeFDtrwaKIG2mCGVNWSTc+MOPqBfHwXuESXmc6pYzUkDU6m07OdjBGLfUJhii
qD+9GcpvnsIcex+hoXH189hlzU657xLFU+OCxBGMAJqI8grXvQZ5Kv3NG1FsxI9G
rtL53gh0gq7EB7UzTctSTO06edzCMWo0vYoQ8oPQMWNFHEo+Yc7zai2/mo1ib+yF
fpUEOq5DVnvLLCGUblLw7gr/UkdBXOB774xZefbz1Q4elQSOzRRS1b4cRLkSaNa4
y1KPU5aIuXFoF44jmyP82kYebb0q06tcv5jLM4tK0B0GfGiHR1NxWwoDoWahlffx
+8UyTO8/scaRPaeVlWZH3dlu5JzJ5bJiC4ozb2jOmGbzpQKkFIphhJFs5HqZnKnO
urPvJnEg5ZGR5+UtG8keHCTAhTuuNTpystKjovjGfkopWJA+MxtVTBTBrbNzU+zJ
TQXEN/MyTU812J8FwDI30yy9hjRYaKlu8X8QpID8ws9pL9HSjknU8bRNRzLbnjKD
K33TRo+TyeaVX/AIWzaF6LXNJwUaSJIFt+XXQWENH3WagO9hAn5VegNmuif3RYQf
1TcDZ5wz0+N454z+ji8+wIuck7Y9dFjKVVKg0oQms7sPAuSDxShDp/vSvet3DkxM
niFq7qopkzWUfgpfVYZBatmgIKy3r5lAmfXjyJGGuA4tJWGjGkcTjSqmAd3Pv8rH
k8703YpwJmSEqdH4cnoWMwRN61IgCFetlWWv913gEVtxXsielF329XEYuLVWAVmc
fndj8y9qDy3Rztid4INH2d57CdMV0aPQ72WvM0X0bNSfyvbxn9mFNkWQxuVNVWsf
XUiTb6ZbPwdfcCdj2USmQpoSbsNIyxCek7ZtiuI5RrtJfBFRLCZwsfFBDUnynBzU
2sn5lnZ706K8sHLnQm1/Sd3QpC9uSSmJDdV2CtGFF863y/fby56WUjs/jQ0HuU07
vKsNtQTGprWjSpF5qW76rkP60a9hQ2xOAq1pzucsJpOVr6t+g/m7Ezye+cvdXlgF
xfRMdYqTgTf4HEHdFsVKlxGjZsZmOPjmV5IE85UbZ4d5kjIB8MrN+UJSv+TOIVw8
V5DsG6reJJq0odeeYkmP+w==
`protect END_PROTECTED
