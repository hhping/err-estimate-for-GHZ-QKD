`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SxH00S0gQxY6S+Yfo21rq+w5GRQXpsWKuylf4wYIg1MiLoo4EbM2cKJjcFX9i7WE
KfrJv2PrbdtiZsldfrRlJstYFVz+TX+qyWmA1LWfRExYKfoQ1u0dBBS+FPcRw4fX
hXV9YNcgjd8LgCZ+ONyg3FqtTTmT+Id5WpjWhoi9R+sJrlqkFzSXfOx49aCsTB8F
B0/r9y8ZmK84VxxuWHMtaPsI5oIP6BMtwFoN0kKnTQtDvrGGMu+WVZcHrArqUI7a
cwQz0I3eeCR5NnyUxK8NHNiJjFuNkzm+QDUG0R9YoGtAb9dWYv5EqSMoiAji18hq
05ZbUnVL9S8MLnA+/YtUOExdt27sm4w6bNI6vNgNzuWp4RgR2IWJtDm18trwyP3K
vV9uUv/QuAO5WOws4JupZw/UEsAgL7TyZO/w71dCjhKqwssiVvGMkkykagTF8BJX
wVrfhSxuvcfKFcvggL5Rba64cQs/w7HwQw3nbusJ9efgykvwgSfYy/yy/g6NRPrh
fug+bLBTvVNuFiJOG5vBKS1w3UQQ+QxsYYOebwH26UAtgn0j8jmGOYZoZgM8lKTn
9Q6h+XGNQQ21ydyvHL8ZOtYmEWEBWWi2bBZKSMT8SzVop/M5twJ9l9+sU/zUEe+H
DexxfoBRi6GDqaVDTolcyhY0AIgsL7zd/AR83Y6Vl1YgVyCjxYTNdc8RR4Bjo/4m
9cv2YFhabbL9nmsMdbQl+9Md1EmoWPz3hTdS+imG5IoXTYcHx8ASvK+rmdzRLTkV
6xM0lm4UN51APpgJvOVTDlO0ccE+ScVr1d7WdEydry2t+A8T7w2HvVFvtxEiIv+j
/6fDpM+rq+50nlZRto+w1yLa965ISyA6qLGbdkmuaqF6MU7Cri2/oQdq5KwOVivT
l3p/5ekH1CSfLipYXCqgiC/xTRG6Cztaimto4PDf9J38RtrD0AtToGMYt7Tabl9E
Ux43fkHLguc1QOnHncl6brT40D6mZbp7MN030BpeRws+VPFMRSlX3mDgrdhrDr++
e4tN5WBwAA9GRaxUTAoicorTC5UoVRhZLg/+CarxnjMQib+yV49JtwaM6KHTP/bj
1jclVIkpF9D0stOWug8tnXKelo9CHaArxwE0X7502TgNFChzUQ0LJW4C4g1Y86X8
ZfIxGeIvD94Cwc6HvEqrEd+jYQtRMc3LfdxVEqERA7mTcYoTDC0foi1e7m+LSVlq
rYU5FPVciSE5Jz7ZfjBg4+DaObU3wmOVK7c1dBmyp0O8neta4GaMQ2ea369IFWTt
JNH10030mRHtrvPvgB2Lq0vk9IWpytFWq/DW92U8eGM=
`protect END_PROTECTED
