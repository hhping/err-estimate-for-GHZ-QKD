`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ro5FygFephvWI269U3qYN3W7w+eABqMK1jiuEAak3aSIApT/wUEzkNtlHG9kpJW
Lm6/dz0CRDj/DhYaNbiRARuez0wKEzPyiEtsmtIVQW77JFq9QUWxBsLTnZWCbhFT
kyUAdgElXSRAO7mn3vQVoNZwwc21q8EHSm7QSzoB2X2TCBzmku0ptZTA+zCfxu1F
fVCEdO0vK5BXTZNe/cOqYX2WciVR8eEyuC6zag7GFb5K98dE/ZO5lFADfMscNVqx
i+uL+USOIN1PjOt+h5ovdlw5Crgos+QqEcDLZ8D4L9wskLWkW4UD/4chCi3CjWSC
ReXH4Xbk95/bfRwt1s+wTsVcPaJ4BfSxvEP4WHF2+PsSQn9T2HPWm8xlml7g1UYH
L8DyX5ZqHnBMUD2o61wI1adbDblqPsscTBwWAn9SrTOZbrtgng8/q9xhDA5/rZ20
rGTdZaKlY+7v78bFazou7SlQILQYzitxgQB+9FKK8mI+5hIzaFWB2syicaT423QI
ldqUJzmqQGA0bODQBP60Rdnx/Q5usdy4SPnCB8b3J6WLioRDDHnb7m7sJMzCMurH
fK2jAsiJGU3Qf+qXGT/hOq+RTlp6FNqyARd0oPEi9bXU3LMH65mvT4e2fycgWkzS
OioNFtOwUoloNze5mlOHvCNLR921BQ48ELwajP1RNFQIQX2NzAUVfJZuj95cIjWO
WlOQOf622GSYzVyuAK8YcvtN0FkszEeM+chog09sLDMiKwcp6ZqVU0WMRtDPupJh
G0NCRSzfqLn3Zkcvv99fImP2eXKWVRe+do6bM4ATgi8eBObXcMB2Viyj1m7+IZiQ
xi+XQQDa3r+8hmMZUV7cL2KGuB+ved+8CSX8XAlx8UyTqi7xPzH/4RSK65gpjw4l
skz2F2mWf1Ks2KwXlxmKPp4BoOGwsX/URunCSDjubjlHsDhFF/kgUHTsnodHP0iC
r5wjeEmq9BrLHXkTq5Ec8a3MPQMAIMeNMuUkYvtNE/qlk6d74ty1Sx3m2LuCpooF
DwpWCj1GoA7lOc7MhSD2Zy6+eRoDM86XCg8FmkS88g7tHZsuXGWcwg7ZnKB43J9R
m9sY/Odj8mbjjTvzXaTFsHvZeUGu86Ew99tXtdS13viB+v7XcNGFmkBc1g/JiEh4
jmpniQrz7nUTee5arKxUeMbz7DgQpmRN3ESHudLNJykNID5zlgxy7uMRx+HxBGL0
yxAi2hmW+dxbeIglLNb2bcBENzYHiw+ILqHhOvH73Io6/o7eT/Y7zwjfKukDQH28
BB+ZHdng1+owOd57jZFQTqHQexdVIEuOlbaFrbwaZ7WZsJiFAYFSlCJBZsKBsv3M
/9ZJIpB3ny8NxuG2WMWelDpCsennCymNaGkOpZiwnz80OjVAXwqwodbdja7WuhKK
LTr/2XsDBSJz7jaBoZoITZxkpMc+CGGhXnALJh2nLvRTyP5fH0FjOQI6EfiuRGag
GvnrQi0reyxIeu41RvK4w/bZPzhU5D6F/QAxnVA79ukVHdfEDn4aRj9HZaGNBwB+
DShB+k0G5P5xZ88VUPqthjo96JE0IqfYpx+8R5Ms9oQ45yjTQNOWBLPRfn/RMWPk
MvJcYPDY8Hthv1HfLPO+QmyEm9RmXrTWBP9zG22cuhDE9VHPReVvRnY7Mb67/1s4
NruSB6U+/m2emm8iLo6Z7cj/xQlqQeSeSrUj4dFAe5AUoO7zdr+QbCwSm7KCdoBa
jHzyfpaf3aw1F9uhGhLcHzlYyM55sxGeclhhM8I1V+3vDkv83FacufK3VIE4W8fI
WuSEmA0HLm/z1s6gpP3M1eCrVw3qBhZYPHjQZvi65xI1TfGoCM29lmORYKodN7VQ
AAPZxrdYiFZDNWIXjrq+S3H+lQOKIBX+6SmHkyqr0xu71tbZP6a+frTIVpnBR7pD
wCCdSOZnNLOTRE6N06MfZnsruUvE2YJvTJzPtUrLsssh2HyCESAPbKzLTspM5607
HohvpAuBzS+kR6GAbMcWwDfy/AfOA3zo7HqTySqzyL/hFlhLGe+ABkOYddii9K+6
1UQvMqBfxlPvVa19avAM+7h3SHOk0DzZo50TyG8mRfR4aOOUYjpWYLnTycwrFFvO
tLdvr/pC785OJrHzw9tfQMSjfHQxnrgmpdCU5GuRe2GY++JZ/DQCZ17VyulxQsiR
YMMXydBydvHnFjMLmpHWngeKbdKErvGtERV7uDcXfFJzoVKJFFyqkAgOI5cCh3z3
RJdSqlUuZJBgUuTwJdmvcVTWi/WBYJrBZffBw3XNEClA6F/qQgHRWnO9nEdlmiyC
OyuFu+4XCG240CQrAXH/I+9rXMgS87e3ID6SJtMyVpytzqYs+BDjXBQqfjOlG1MT
VKHB2Xj2qvnp+hy2Ysl4gMNa+kR8RVTuH5N7kAhemkTcCxHDxRRMrf93fE83xpo2
CxT5iyusTX50sQcoOKLF9OeSIUoXpa/ShP50H601eprRcC+OyaZ00+DRGV5YsEU2
4X9TPuy2xFhYywBDrHyY1dC7cHeFtSEilpxkRgJVgxsavJsuNC4/pBBpZnDN4uvF
LwJylwA+J9+PXGqG+7S3pbuFnGYTBm1+92cqr2c+slzDU+gvCQaTa9GMu0MWMhn7
VIoOjTsz0tk6oABVQSNvVNS+bUqWfGTGpeMzGruhf+r3n2iWbI7gG+tqCNhAgU+2
zyse7YbxgynEK4xcwgJ7b5f0Pe4k4GOdUtrQETCoYDvtrgeSjTyAlglSAstQ+LRh
vU2T1S/P4mmAPI66ghtaAUMIzcQAD9Q19KXBBI2MKkY0I7M5xlftqEXAtN1TFEnm
Yf8sysofonJ5SkvGJWTnOymkAeObgPDuuNaFcpTWhkVDEme83PQyH+SoOaZ/bSyk
Srt6X2yIgVXrt3jMMSe8IUQ694sea2X47hxZxevG7/53LhM4nQJh3xpQs8FtzaLv
BZc2JCCtkz5dzAEci+h5zT6oV9kT6dCQfAdhQtmSOZs67Os9EkhxcVy/d1Io/GHq
iYCVxmoQCUNZOwoBWFlh+et1vg2w/29eF4z89OcJHCFkTU1w4SxoiLlPWzg3L8r6
WQ8qsx6e14gG+7MmzhvsTNJIBTuqOG5QO/kNTbK130Rygm4QCr0HnTyToTCLWts6
k3bVm75KaGpKRmPzAslv3jol6r0oWgMEr/vqUnX5pijCW+qMiweN56KhDZgC2SHO
OMhi+WFgVmOxgdFq3Vb8aRfXAcMbj+diE4QQBs9+KoULQTtfgHzyEuLCwyx8CosU
4uVjbOPNwwozMMvMPAwHnkt88trIHXJGB5AsAFwo17wUaSs/sz85CrpXzpY6kmGc
sBrmFslhuUf2GiU8uqEcKnSNX97k6Vm77tbiNXw8yjd7c8WcgsdDobM5ny/VC27D
jds9c2HRXWhCuOJ1RMVr3YWGsaDJ3A2JEXLZtIIPZ3n3bspShhkzquekrSbZcVUq
T9a3KiQLyZGbf/KNd1FDQwC+1F5ks0/xVINwhD/6Dh0mM7WDZRYqOb90ul9nyAxX
M+88sS8+L+bXm9P1Q+O2ySLda35YBL7239bOx9TahJyDubiMf5bU/wzGRe/Z/wRK
gpFkjjIENKYIBf+ZD7tzig==
`protect END_PROTECTED
