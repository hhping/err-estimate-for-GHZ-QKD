`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKGhSv6PMtNd8RN++jgsiWeVXkYcJvuhZq1ce9YOUB2DCUXdpi+e6b7sQDZvNRnp
ovPgLssDjUHOwEUMzfqRU7aciIBGt902VR2ehDA83yQtp6D/YOeaaHk4ysMvYyUq
8uLL6XSO1ueeB2wTTedSygF0aH8ZJXt0pOFE3SHFYaB/5+rXu3d2drwWmWMV+gdd
P036B1CZUeiQ1rYiwlmAIjagH/wEMakAf6uzfNdOkfp5RbL2swe5CMhUJo5HeQp3
4EmRhWBz50n+zfsz1nHJYoXGhuZOh/ePWl4r/8oZTJPLaVAB5u/2MpxcEj1EIywO
rXzf6pBvbTPJYqp52W0Qg8DaTpwpklauVwCPGqEah3NgZt3O+TfYUqprP/rujBd9
tTjV3BMZuE00RtL/HDE8XpyiUrqtRM8t1PLeJxsk4XXc7CeWDZX3nGbwwgQ2fskb
JDcy+Gztfvwop2cQr54zOp+Il3fqnRLvAGwMXcBwsM88kVVYl+bVoMBJQGxl7BSh
nUns4u9+I/WQawDaGH3udR7mEMkOPMVLk2ApYB9QBeg8sHSTaTL6PMCF5ZethQ4R
TXNMHR4Ix4ih/gt9FMjoB9oxiNrcN4H9bFc7RHFmYxKyApRaUB8O2SfCTeyhrUYA
CfA2Hv6Un0Vld7dND+ubM+oGEzO4Fo7gcUAp1g1qZPBEC6KmIXS1uqZn/vP+eKja
/ld3ZRvaMsLflltt85fxp+2CB/MiPKjumd8gUDXfuqbxoqX/p1+R1JR9E8hJwhZg
tDGSfoQHAGEXybhDM3MjfKiZ2Im20k02UJe3Wkosr9b4HVPZcFJP2LV9dTCK4KZv
B58cZFUnP25bbH7iHIHMI9j8zm3HFIRyZAUiTotrp658Zw1JXMe7uWD9aLJh/OYk
HeY9XrFYlhHDOmgqITxpxBxWDvQeRRPwvkha9DuUSiie+3qBv+iZh7QwS4RLe+PI
JP6cQgPb0sA6re6924HzJlm3LoSS9iG9Lkz3MrLzpqGaL6Azh4VduWUwsjY5AYun
9ESliU5zhRXg+/+aoQjK5iH26tKVyCrHV6yGliakJksBJ1aIs67836YqUZai2OvV
QKgAfVvE6Lzqs1GGAnn1u3ZWHHwivxb4A2K3wUSeJTNt1L94VWzm0ks1bwZLXApD
3N1/vHgOb4Lc+ls4FdUwwZWzv/g98vx5lECD6lXtPBdpENsQ5ayLtu+9xuTubR6l
iL619mnk6XiZOc8kcxvI3cFojG5CpKmfJ+8LWttYx3hwj2hLLYW90+BAxht3ydOe
HEBAadBG9tXtUISxkR6ZQv6UzE7XVwVCNRWHUNeeKhYJYZcrcK/vsIMPq11WWN5F
7q/6YdgvLICkprxghgvrd0IPNmFSuIBVtNy9prBlxSAK9FYfvva9N+ki/Lm1MIP0
SP5OqReJ8rJUjXd2uidmCmpJ8vz55BeCrPc0O3UDeL/Juo6y+LvZIxFNh/dMY9Fn
Pad/arXpRpXRGD2jY7FOJXOx4iUPIMs+4WSxAp8j8+YYn0r6O1hiIuZPyPTjOMdP
yE6RYqhis+QWel7SmbT7Ts8r+5qnmlQFKIbmrRe+iFDgs0DyKHvOWlLNovR2iU22
3ZQksoIuTJ0RHSScMVCcv2I47cFlOMyxAJBHW5i5fVSodInkohWZ/jy+jAn1c/nM
blUYzUfUZl6weHBx2LAe4IJLsAyBzHNbefw9L1av/XMxtP+UzrOgWKrTALfmvBPm
DSz6CKwkc/FmDtM9HU0Jf/OxPB55GjLlTJb2YPFrb56H1TifDH+RgEbw+LXRF0eB
yTQ/hzrbUb5sdcNTvx2scG+Z1G2+ulYk7GvNebxkGw/scHOH0IFTaaRQKJNkDLN1
ADDhYWh4oDf1ABlfYsOGoIz0vAzu8sUyUtJK0G8sLjJ7yCFcdMNfafvF1NhofmMD
4oZuP5CCZnBY3tVFXZ1Ouw==
`protect END_PROTECTED
