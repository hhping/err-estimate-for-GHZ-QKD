`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44KbmDHPpxgskJPPcRZ+7TtFWsRlifOiPURh65RdPHycEGjKRKU21J4ThfWpMzLD
YdW0VRUGMb2XIN159Ms40hTK4rPYC0FyVL+Mdq9569EQHtRjtv7wnG04NIhQCmbi
66b6TYyhONZiG3x6zHlUCG2OcovlLD79T6M+eq0i3pMr+8B8ZVpNfUzm9G2ZgqjT
wZbo25fJFR+DA18vNcZYDOieqzbxNTSTKLkBOt7xSVJwAkgHSK8WHPvf9aiZx9ht
zs4XCcxs8QZ2o+PjpBj7BYDwyGN3EVkScCybFXfquzCKh/oL9UFt5rY+Z8uAWvtn
rTXjlMRLiB0Di9IG+pA3K/tc0YqndzKQsnPnymuTRlZESmy4Z21qxakaAK6hWGSF
ygQTjEjg+ZUxoJoXHEvCDyNtVzYYEqu6pCSrZl1TdNbQ0NpuubslSggo1UbBOlJ9
MGeH+2tC+MMOdz6/V/bacLrwgRyGQI/SIG2vvAR5UAhAwWOV/W6DJ4GCzYdzyKa5
CGw7iHFKUIq/UyaFteniwj5zQVISXq1b7MHdFgZHeMIOUTat72vlxh5i++qJjOmA
K9ir86dJWBqg8jYhM81ean7CQpFSYwEkH/F942UYJE89VwcoJh5lzMRzk9pn+72t
fqlJYJYcwL3GkUB+xFhfTGafUSOen4OrxTHYp2hx1n4=
`protect END_PROTECTED
