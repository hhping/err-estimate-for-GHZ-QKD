`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18SaVKiM2uBYYhojSPRtDQ/9PMSqP5yUiR80ErJbiqxJfS2qJvI86b3VFt3rSjkW
Gu3zZdJxiajMGjcbwxdculB49BkwfrMgAqcdcpOK2I+4IlGr87KkTpBT60onETmb
JG0URt8nyvi2df37aJR480B80f8MAtMZ8f3Hc/TC6FhU/TC3+RJbozXK1UoqskGY
Y5HSVLGAcltE7I4KmNF7K8tN5oc0N0/IaSHQuMHjc6QfrhAeXC8tKzBbqPDFrgT2
Lcl1qtSPcNejFIF1rqAmVBtu0VtdbREXGXz32d/I/SByj+bx8KUaERG8xAkPl7kb
zEbKc78Pm7QIOoauxTj1ft6eKw9LV+V83XJDNb0wQGYQF0Hn96Rg4k548c3Jg5tJ
G5bPpVu++IKdXtt+fxNIQM9oXTUO1GpvjPDaHlli/D35CTKyDw/nsSeon4VDa3w0
8KHfGD6N5TFQO+DcDMuhb/iq3Fz1tl14bsrT0McV8PLPNfu109Hkvd09SOyB24Lx
VcEGrud3zhpINBFYHgMWPK33OJe2TqGuZ0aP+LNNBGJniyyEBnSXPfws6qAaH7tm
f89IuLdeWqSJXB+WB037sx2dPPSJWIaY2W969DVT5q05JuAMCTYSXC+QDRQWPvOz
wJEp8Cnz/3siQHcyHXiaNJm8yXiQ4ndzlK4lIlE8drEvUiyD/H2KRFcrNPdDNZzD
OQsOEFhbuprGIUwHS+8FUTw1JH+0b8DxKbYNeLw3W8BOGOkRmYF4lbBk310AWlHT
QS7tk2g6l3Eg9Mwn/kuAlVe4wwJnZiV0FcuDdjmcS28DrC62am5VMlcrSQ4mXEIL
8+V0UaIgNT9g0gbHgI8IHHzAGfetZGnAy3jkBNc5gX8NCfVZiiD4/06iG9luSttD
0zBXmqnCSjynOhYd5zVxJunGez2euqgkJb6ZFQVrO3TWgoz8QCKDOz6//+nHkgyd
FoM+mXIC/PYPvp0/WnHIErClfEAova6ul+/dj4PktOm8e47BNPgBhps74VOIX60b
/nLUJXrB9XSf0yNM8qQYJ8MlCYv0c2TYSiWB2PHxB+WF2kJ7vO3z6ZNuZ92XZOZe
60DrsqBx9RikKzDEukMAdcGlj9W5G9+3vCwHAkOsOFw7k9j+1r1x3BrACw8HPsPQ
vNBJHXfgY2WSalAImRokizI4y3LluMrVgpUdDOO/kF/Qv0ZkVAvWGswlxEiobT7F
70h2iR1fMT7r7fktYu4+cPt3K8+iQD/PqOlQycqbmUnraVBBulbdxUFwhYM0PtMn
G7EE9uoDUydB1a4h0QRit8Hth6Q8dxqjuG6PF8cjQm9V7vV3wK+5O/tTzj1XG21n
AsvsHfIvppTFCsrX7a0NJYfYrw2Oo8Anln7MaRZB0jMLyLMj3gZ2Wh2XbXKHXAbq
eo7ApI9xb1JVvr0mGakI6iw0uzl9C0N/MwDxoNS6ecQi1U9v2MaJzDeO4+0/2T6w
UXORJygNyKtdFqqHZ/3JHdySbLC4qPACfDas5oxkkJA=
`protect END_PROTECTED
