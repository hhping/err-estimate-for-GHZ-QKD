`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yabsHpJZ3zH6chAHia1uvd69vkA8yx+hupWGEQkqGQxZW0F5D3Yc0uGZMB+4iLyb
7OOxEGagpayAxw263EmIdNd/Gn329HgpL9r7khG6BaPqe4pJ054CtpECoHgi5Iqh
U9iZJ5JO3WcJRt3q3FK7ImRWKH3PvRWs3aDBBif/+6d11Kp1xi7SKNuXnWN95HQ9
t9p95ZGq7eAAZz8LnGnRMNm6SrtL0Kvgp4Dkzf9nHIyIvkuUQ2SFNhes13C8MTgj
2p65D2NbQ3cMvwPtGYQhwDQF67+j5aA1LjrLHfYEXPDcuPyboa4cYsjaPu+aUR9S
ButCC5XJCo16YSJA8394ObERfAOS6C+2Npv0/Bee0/43lPqWo01dUPzVlH1cTXAW
6xrwVZryTkB6LHT72nPMrBdL7PAdjqAlhiie/X6+cJxZTmcN+VDyG2V9zzclmDUB
sooU+qqflKbYRf6ddy/QRd6ITdoZglhAtBqI4KQQSKHWHBx83INvsUwvamBXeNGS
`protect END_PROTECTED
