`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQhC06hmS8zB+O836IVeExaiE15Tq6SrB942titmPFD4/GuGdhfXX2aHJM5WD/Qw
PkEX96MxiMXz8Z/JDAf7Xjj9tTaTClcGG6VMwv0zrnAbWp8LixmVHi6iax+3EoLm
7f6ioE9Bz8i6eLZoWx6PMW3OJh3yGVe7nEwhUa7xtuBdyBDdMICiIuiT64JjrXjp
dzRWNrSCOnb3W7cBH9j8ql2G6hXHh/TepgBCslV2vpai1M7IAZb6AbdGnNQBp/CT
/6ZygpQjw0FzNQFi/+eMyxYfpiPXJJD6bGpAt+otX9/Yx84NgEuVjfR3AIK3TZ2F
91uRLOVYfL/TuAnbRJS+y5MiPUDNjUJNGwj23e5XAMBSidSqkbufX18RjgQqUSCM
E0de4MOLiPsJ4hnhKiFPPUmq9y14+NJQ/7llfF59ycRGv2bPwiCvPupCa0qCItKU
iXS0Rcx0incxVpKVWcJO8QVjH7gVtRhaMrSmDwRGGDV+HplyCz/rAyv27HDjkkue
qj4thysjGDebR/5Fd12R/3aFWrA8tdrrnsxLpbQsJGow//CdRXbX5bth5+4268lt
NTF7IHtS/pi3r3VbNWSCCdJrci5WSIf44+KrTgWgY1ItYAKmlaUzv36l0F0B/Rpe
841OAx/xUuX0O2RGdKE8TT1UGAGeuNIy32audD4SNrRb65fxqdqi8gPbML0FRwBd
zu0jry/SUpDiZqfaM/wbMTTpEX2QAt9WGzSZKm9ZwrMoTOxrcO+L7tyrFgSo/SG8
lRYgMd35HapXLVDSz550eUKfDhgHuT83hpe5WLxnmsw+HXmB6CnEHrXMmYHqpjoq
zCGpwS70HZZZi12cSMAng9FjJCS6b1Fz25cAC/0r0VYoo3mKA3rzmpPrffM7WiRt
VXVgxKfS9fX5K+BkyqIZ/8Oy9PvJRoqxltGztvdnsCVE1aDkVTBlFt/541Xh2qhJ
/C/Gx4eeQRfb66wTBHSk5vWELe/N+PR9KnqLmrbGJOUN9G2SXVqP8rVFt46cxLR2
SBV+u8TeCq8I0NIwh1eTyOemwZAFaBQRuqVBkCxR1m2CoORovfSHs0u584tMHNYH
lRsy5YpE3VNbQ+Db2vfAkwp+1rqaTHhxcRMPC8TEWOpSaFonJey0VARJvijkZhxX
wAvpzZTICkR93/YrJb+9BmKkH0G2QvxCadUQWErTW5BwciXtqRNGGKaJVWWtRhtf
C9X3zoDKzUaiHEFHqev8Msv/FYF63pQ48N+AX5by60bKzqeecq5HOExAMm3KGAK9
VRVi28GSMwcduLVjfnWvRUQvVxjSxY2RSeVKoSE+3WtBd8qvn8HONwr970s31QhC
b3LeHXIwHKIEMxp4kh7RyvYJNTHQSSJj8eAetjg+iL6QQ7orZD7ydGHeNuoiEaDF
PBopjhjcyHssbXC1HV6OTKuwYabK9stQoWd7GiudlMMvLux76uE5IcyI84dJ+BLi
8eHHnZICaL2Ta/uqfHd5CTz2v4VdrrT4OCxBZAY6sgg7B+/CzZ8YWekuCByZsq1z
weP7GSfP2F1Arz2zX7LphI1idjEaKD4XA90MxKuotjTI406StTa2v0gyEYQFDQgS
5od+2CD0HCLULOCcHBSDN0crJs10vmVkVBFopPqs57T1oK3z6YWohtoH9pl3rBW8
N4tkbA9yd2Cs8Mr1PUQUVETlsD5uyuVlcu2F20EACHZWXjxa5WPQ59J2SPN8nm5K
oxxtkRlJr0jMNi5SEKgQmA2ckjsvV/nU70BiGW87JZDfCp9UH1bjxNo7wdOK6IVs
Ps7JcOSEWgwoKxL/4ZTp8mUusc5BMdhWLqQEFi5Oqwog/vseCWjgWRysrhCb4rhj
C/S+K2oTBQl0qCXLNXXOzdl57RP9j3CqtSy+2I+PWCnVM+O1wMUO0rA4pVPwAxRS
Z/eyfnXvd1YswNF5iko5c6yXTt1kVoKG/7n0r66KWDM=
`protect END_PROTECTED
