`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEFt4QEYch63OQcmQOvVxeZ7c/COSg3L14W6eJryGGu8a4rM+3HhCWHKy7Tixobd
fX9qCHVUFP8RotrC0s2mCVJUTuSqGysIiJKAbRj+00j2ADxyFkiUxQ5La/pha0oL
5VUQOwMWnf9qzCm1dPgUjoVd+yRr9yDJXuEnzDryLYNWVANy5lwbfnGxykMi0uHz
bVvqoZDQ9MBNWMXXXCc5OmnfDc4OGneVyM1sL7zurnBM3iKV+g97mzs88wyTPQyv
9/1ZGZeE74CfVzp0Qyh9Sj1V7YeePph7djthki874z/MbDAPjxShQNsIGvUe7TH1
AxY3qUUEnIrK369CHXtbED77kBgkcurprfsoAec4j1NC7iMz5iVZesgx0DNLdHNj
DLswchGFKY8cld6iIyEfJjRtQ4GYBiiSkB+DP16oEyDrNqonB6RyfcTtLG4I2Bj2
YpTi2qW/diQRSqdV1rRBMGaIUkSm0akK8YuAPH/NWKoZB0mLR9k2UsCStvk+C64J
+zD1/fXVhtC/o8D5cxZlmONiwF6bSVvtk2aJJ4PLYVvU0P2kDIg7WqetR2EcjYA1
ZcaHnv2qKq537gi9pFM9an4isiUsrKzeLuIJX5+HD+HamEjfYdjnK73gIUF+Bcr5
DJBy6fNHYItejvvnU3eAu+QGmErm+rz9C6mexj06uGyPEB6FCMMV3YW5VFr2+GpN
76DlGu8q8OjQKqyK+k/QCwwwkHRUNhrpMy0ms0BSh3SLw+fGQJLSGaoBCt2z2j3U
UASxmvbB8DGtv7qgS/tvIaFaevUcpd0cin6xf5BkEMxeBkmMT8p9ekV4s4vpv1hd
GUGHGqDSNQlwqJ1Nl2ss6LCYkuF4YtzH82or4JieHQ0WyArhsVyXpbQfDFMnml9i
cn39zqIC/iPeEmGLzcJMH9GRQ8ghBR8DxcJO3W2c/F8+QRUMmtLrk8TWQFrxq8l7
W21pwFdF4fdBsOf/hcuRD/+yn1uIzEf6yy+uB2XLnb5ZlHQNVqlqfhDa7KAJknzw
uTbbjLRzal5fOGMOOKrjpjjYG0CSav+E2jrsTVm5sD2BDI25x6RuI3lOCRdCnhNO
IEK51wJdIDtI1T5obwVo3+IKiZSRUXtOdZsFz8DHQYHUS44XXtYAthMD2HcF3dRp
AUXSa+6sBT+otepiK1YrDAGdrWHLIW245K7fM3pkm6Ht5H0E3TsEaqZ+tCrAjPV6
y3a2Dx4sPFMKnDwbup1ICHG5yvh0Ycc8FX+Lu0e9ADO3fstE/NPHpPSeHozPW5Cz
xBdKJ074FhUxgMZpLdafjmuBNU0/d98gLxJnVFHJKjW14GVYwWViAFdNOuMjhKoL
5bM5SCCL4+prHR+1pTRaq5v66+ykOGTw/XaqT/Sxa+4aXhUT0PV2rrFAo6+tmjKJ
8deOkaMSjjegitE7kLrMM9/IGK6KOnV5YSiMjxxQm3qZzyZZtFSzSV1My90WZRo5
OoLak0heEdmN8cc3DnLRHWSFexPcxUQ2kro0+GIl9HvQFLd46WZ2oH5qT1O4xTlg
RD0H0+UHbO8vEKpK5Ad20Q+NahypEM/ZZvR/HEzAHbeimsWeh+CCtJ/t1UJs6okm
QhZ5Emms4UZFpvjMm3zowJapkypt0WuT5A3Czvh5DUWh83EHg5eYJXCLpm7ZtQTw
P2VfmJkkcbAmv/Jrjj/BcY5BHi9fB5480nLYfp8989Apy2gLC04M4cR8M2QubICp
fH83IM6bIVwZHZrLYH3eFNc/h5ioS5XVuQ7V7uAdKL1bIIPGPcWYylbtuT8vwA46
fLxNf9c4C1i/fZkVHP18QVFORVFpx8LJykDyRZ81gh28atwtApq4I/bIyNVyrogP
0UpUXSNNuzF2pyX3Otl/tqFtKzodKkJ/QaNbeULzop/WQW9Bf1jhC4czhlhrVqwE
xlkLcP3mxTA9UCh9IahqlpAHUgeTeu3JH0VrwxlYMJR9cVblJIb6hIVav56yOvZJ
IsESbZoWM5NKdwgsBRxPIt5UoE/821Sc/6dYUW0OH1oZJxokgyPG+YpOx/BW1rJ7
37UYh4q7n7TtJCuv7tf0rOtbL0esjWN80cMqH9iI+92ZRDWRpXZ61iKj45uUPupC
RTpGPpb3t1x8qXNk2CfqiR/HA4XlkeS68n9SUbu0oRVSkTxRv/WZRvKM80TIxYbO
UFx/+Yciw6TGc9szC0X24qa8lWhC5j2OMdN8KaHXhekBgpYrD2E9chjYXP+/5O2z
sc0L7fOND5s9fHkUlVa8b+0m/p/Og3P47J46kgZKn4lJ39yhXVO4sfNXbgEonI8S
Yc+oReVN18+C+zO9mynccm4Q/VEfXZ3XSw2Z+IcOwIcbZntm3MOIdTLyT3hpIGRl
fknhidI79Gfpq4Xw2loJnnVJrRC/v7epUjOU0dYnZRL14Z06a84+PDp8dcsURs56
1M3e8NhNKQBtwriQ7mCS2g==
`protect END_PROTECTED
