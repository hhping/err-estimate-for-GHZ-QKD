`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2VFAdH6WEwQIO4hAYNOG/EwWWCH8jcE7pEm2UxR0hdGpbx+G+MAhdQZCWl9xTs1
8kp4lcY+g9ZbK4K6lVagq/vdHdzKwl3njV4Z+uA8Y499xd/vI8txC4I+DMwYigdO
anp2RYW3iFsXNO5dWz3ltUkHeYKZ9OS1zPCjcM5k8ESGWqKIjYBtgLfjoTxOUK36
HBluw1gz8GFeBdy6lqC12xoEDeKQrIq25s2RRe+K0oV2AGjOND2KjkcVA3D4xAgN
NdI5wtv/aDs+iIt9tJTxxfWyI4Zcbt4y3SAMoh8Cir3Pp3ddhJfjEy52/iHUcpVW
LuATJAg9BSqf24vpqzRiraC4mWPlQ/M9vxmT17IGX/+SKH64TjXD6wnNJD6qTt+o
yJR2+xKG73NkmfGNGjbkk0noZNALHchV6gIcue2l9ttIwaGa59X6ezH4NfuGSzgt
TIkjAZb1YrxHjdAH1aDLgx41KFSzOfcaT1Z0syaEAH2fAdSLLRXDusXhDUl5ybtb
x4QrKZrZZHDIvXg5Gp0VBrPqQJRMbtlJEg67gP3zW7JlXdwPFA6Dhb8+RxjtLC0o
UxoIJ3deod4jXkYZHWfMJB6Sq8iaqYHJFvp++PECCI6om2+8fsYNTDm90byhgNQM
CboSIsOO5eHyvuwzniULj8KK/oQBeu3tdmX52JFDxlGw8h3LBZQBsAYJBIepQ/BF
XAbOYLiexb657dSqbvROfn5yvoZyrBnifEnAwDCvnCGka0KuHsVa70PXbNql3p3p
Q00d4BgIBX5oWyZm2MqpeyIG2yKBtodpvvXtelIT+WU82KCsiT+wJxeROh4pgic1
Uja8NPVodXP2FW+58aE43zaJoCr1ht0+ALFvQ/ttjXLQYgzW+ADi6+nT3IS7PN09
pPpRn/xJYx+zV4Otgayt0FuM0MX4A5emvPUBtLfOm5toPGPfj3DLTa37dm4T09CX
La2CbhIk7EVpjvhs3yO2llDnruvtuPtiCLJX18ML7+UxRvxViCZMY3oWzHGRb2Ep
+k/KsC7qJlyjibHIoqQKqJj23oxcQRu6lsYPvM5Hcm88dMKQDvRdSM2Z3ofI6UfM
lD1cebnZBQ6a6RGe0JURYFs4wf+iyiTdxr0+knrRn6X64OYx6zKWhk2LVqVm5uug
k6LIEb8HjpI0oyGWfWa/SNpIwQa5CuiX43jgAtoWGFs5WJf2g8Z5p9APTlKXj2ry
yl5MwEDceK7Re5qGo4JpBFYxubM8Q4bM6kTstFEYUd/JYd7SfkeEutnXioJr5MAU
Kcsw3MDf+EYidHBZCzphZX12jSW2dxm5hLG94AS9cBfrSABGoYNOayLBM3uw0FCG
NsopNHe1kOaNM7+Db7DlN1gAGTywaXzPhMt6bEN2W8CS1QEyZjidh4i+op6OgTLk
GWkIIBheeQIQbOiaGN1rw6+cLPp7oF2YesD7fVVkNAS6X1OjOMTFZL3JAFQzIxHa
EA+fIc5qMO9imWuXVOleUqcKSlfdyoCYY1LKwVd4KRVsG1OhysQkSTTBBd8fWAes
ejLPBElx1uqClsz9+0SODlxUdYS4/M6Ddb+fCAyPzDekurIMWg7W3eIg0u5niFwf
LBp8yJUxpzHOGywuglJWVr5TGTtfRiTOZM5crDWZIXkiiVZ3YmH7rMgSGi2LYKHT
wrHtVbqtVpSQGR1Yco/8uNK/RMiLt6EXWf/j80wZShLT9LHjnFi5N+/sXt8w6fz9
IgPuB14pvIbrl4pJJBqY3vIw3P9wbT9cAItGu4w6LZ3kTKyT2ySGtEeJ9MdkAyRC
/l2q2gL0M6Q10Vu/+GfNj+81GlYoJrsvAybdBQPaIB7IwQtHAUnFEEidqW1WLHp8
4VibTM6CLaZ6IIJkZ+bfAuwwlJEhBN9HlE3fECamrntypLYnr8O5hCuFW5Q62FlS
CzMbTWa+pi+saNk88ClC10H9IQ9xlg+A7jkSVO4X+h2vt1MQORMVukwuJ6YBGt+r
s5qC//uM/nKsB7Q1IEPgg8nf51Sm+5fckFuXHonHpuYzAJpzXvyrbuad9C/CTk5z
z86yn+KxMwazOR/JVSwG3FxNIif1JanEN135aERKaaZsO44p+s8ocoxdwmWZ8YOQ
2lHzl8A9IGCP/Js4gS9SwArHeT5WzX77FFPuLs7wbDryU82yk4ugtLm0dOdkH6dt
aOFCM+yxIIL2Slysg3ia3Qfjp0ra4NY4HtQpjJFKxbF+lC8f3rqW5mNQBOuPncGj
68xIUKxUiVXxI8+AAzTI0lnWyzVYFypTaj5TD0Xf4AQ4M/MPBRTVBKAKqSkG00KN
YH0hX1OLbjQ1cguo3yQ4ew6hKTYMpibA9kcaS+5VeMba+8UrLpr9Ob8v4Bth49QU
KSEpeAtDyj+AB8pN8CMBHYFkYeinsrGVxmJTYQJ/junTLURWxKwxMpdmYwQqlOLw
rovmf3zvz8ZiPWypUjr2QM17q53LTkDA46pD/svUDX71cu5eBUoOb4U2BwpmsOiP
mk0uGs0eFlx/iJBk0SZGWylFjXIKwaRxpViONhQu4UpoQViHyBlWEcwqU7ib3usp
WlDVkGxZHwEchPpDE0ClzM0Xw97hnV7iznrgkDCmM29P/7RNEYSs7VUAvxEnNzAl
Y+L3qL9gyGqZ8jEO1BSZFiyupAx+zTMETYwiv8ZeNqvBRZ+qHG39JjZqf9zrGIKj
RHpz5pL2mpTRvxWA3+KlYCZKH/87Um80QF9ii2bgE+CG+SRtacQ8gEmI1UakWt9A
ptcVg8A5v+gmZP73jL2g9HRDseAh6iJifG3XipA1UsIG5sv+CN99+i/lJqqZNA08
wa/kdUsM0CTIeIS9opj0E18lSRX8p/0KBGt8zQLeXqjRKYkYdeE0/e+XCPAMs2Kg
XYI4ZZct4DRUZq5OQwIifrgJybtKMVpn8gcwc/XhJ74k6JM+wZsSMm0qTaLsbkuG
uWvu5mO7ZB/ipbqPNIGJGvnJDmJS6kPJ5jMBqaz+QPO/PCfNub+z123PTRPVT8Wp
JDy5eS/9aHhqcIRzkHSnyWxzl8Qn0RkZcIQwjS5Y09RZu2Qp1VOsciwTG8GuJnXT
IAmVSDbTxB2mpHikDKQNyYrFKNnEeitSGVdxy4D86oLiHeRY7iDpPd1roI9r9hpC
MSvH0aBVpZDN8q2wqkMuK8+HPIENIKrjqOZHn9zOmajBQ8OhMqzIjyDz9CER+ag2
/eHuoj7t4t/wKR5BzFE5KTAjXHSVT6H+zp223+QPmcH+SafTc6xtnRzZnlamLuzI
pLEX8iKC3jPuHqDSPHCzhF+DUTNNJPcEnpz+ZS7Nz5geXHJB8hvOGCLunORYG39T
2PlzCcqnav+gJS+qnAEau4i8d0Njl4pdUScW/to8sevVpI2kIpFZLIPF+pJKURiy
SQbEgAW7cALvK8/PxJ5Fb7/BQS4PgGSEDxZ0INxqt2Q1R6xxQGhRvBgalSgML+Rh
Ad0rqvqGFkz/tpO08po3PQ6N6v/8ohzk6e9rZabm4KK3ebPwdwRoxOxaXBdET5hV
9EvOvMWsRAYyou+8TqHPqCUDUzAFDnqtiH6D/yAVBSCrk9yiOUeZogCIBqzXqiH6
dRhciZVB/8DkmvwmuLgjOM/sUJBEpSLwH9ZS8GQ6EHVs7T5ZNEcGWx8CJ+MVmqxe
ESB4Z18p/tfjkwPatp1wxiAkueVcfufxDjdGtEAyiVl4iWBKjBouLpdX2K3garGN
O/5QXTdtR5oaqrEjunBGJ/xRa/QdMpjLoQzalXVTse2lrZzGBpTLRb6o9nQrHQsP
L6Pah+7u6XPD0tZr0yl72g8rftM4ubR90CukxBWHb9cNHXkxozA9FSYFu3NoeTun
TCa1xRvCzDTxJ+Me4SWxvodPn8aBxN0/uDwyKf3ihANIeZbL1uKu7mRm26MnpPL9
ciUrCXPhQli9QniIhKWDa3gqA1DL8xFmDIinMjbN2XQuIA7py1jKQ8lIDg81U+g0
VwppM/B31HECYbLRQTaUe9yutSDut5GUJb+ZoI0Gx/YwcU7QpmbX5AUTZ58Qzz6Z
NbT0qo2XZKO+xBMOixGrk8LLaqZXyeqG+9eStUHm5Tbmlqw4qgfIO+JM0S2SWGqG
Xf1JNhCZSlUHeum5o3ATjoRCYPBP0evEJ/fh+PSkgSmpH35UBbc7vw0QXbVthIXz
068fTjA0FPvjNc/9Pdmd8rNOERbHzURK7Xx526dQOalo7CH7JBZ0J02Hxu//oX3G
hqkv0zcI6D44ETfA9ICvxLh5MSB0CQBSERButwY4iT66NQPYpaDp168yqWvXk57v
f+0i2f6NbG4MuPdDJLvkwR35SqT2XqsoenDGM4M4/O4QySDWp67J5Q17ebI8+LqA
ZY315hzIeYP7PGbCcF3Vco+1I+qLtGvfKy9ADg8uuWNMvOwwVOUgeDEpMeukHRo5
7GzPUiA0dEBPpTFq5u9ODYBLfcSMGjTwkWb41fz49N0=
`protect END_PROTECTED
