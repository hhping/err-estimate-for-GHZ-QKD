`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYvPjffv2cmH6f0B8YjCvwH0iA2+xDLGrdI/B7PYKtmTcmHCpMca2ZUPcLNYZA2W
CytL/GEFv3kJb0vfKrlDL81JEatZLw2cPP0lQRWoKGeAPMKeDlyetGFYOtn6sLd7
6boZU4EzAYPngeHaiBjdT+PCkvAjoZyinAL2TtmXEk+ws3lLN/sVuyUVgPB+Hzh1
`protect END_PROTECTED
