`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2wm+YSRxG8Vh2oIKC9aNnpAjAl+VL20Cm8gbw1/WXjTr51S6ThfFU1Qnqys7Qxzz
LOILaLuIkiq9HDDelGkGDJzJnmhITmOqKIwBdm7buIlVOsumtxIGQR+m6pqlxNFC
OYP1aW526Vz09msptlIIKIrRa4yYsipWULWBDGcG/MtjkbOItmmKI62d+HRjrW/c
SSqx+fwuvbfcHIkO9V7/QuK3xnwCLrVbvxXOzbIJyzFW3cbt5g2o4MDRFjO/4OIi
DF+q8ZV92IVn9Edgh8FMQh7G9yHF4vorayrsaO6nwwoeUleu82PSEkQWFYVTRgfh
Tni1d2B6ZFlncLE4aJZesKnqQkx89PLpjzAwaCcVxHjPa4wcNXJ6C2u1ekDU8jp6
NeApjjNzNw549dU5O4TRs4g9R4Owi5JZPcJYeFE7S9sHc7j9ZU7Hxh67NMH+C9Bw
AIbcNEjyZAT1ahha/rhT8AhG6GoPABOwRtZxwASQJQGau3ZdePu5fxj5AoOVhHfv
2Ngzvu+nVsGfyGVFekI53npOKMXBusLuAT3KgpMKorKs/SZFO8wFJdddQz/PjL2Z
6QJE5m5smNsvPHNoflikk0rmfg5wQCYpMgHTMSLEHIIFk+ULODNmc+P7yr6j39hX
XGMyQKTpuQjcVeHmbKKP6uOCwo1fSZUyDxdwlBGCrzoWwfNA7llItMlkN814s3TT
JLV40UF8x49xK8Ln+Vk9LZ3OQscPCBJBH9nOAg6MCtAtbuG/XKSRQ2Lre9Jcm4MW
AQEcFSl1EMboFY9B76uAnVlvGQHMquWo4H2dL2sovmgl2V1hVeUlarroTGNMwtRa
8i5GvzhlhalieGFX2vEHtIWKHk91Q8lqM6yO5DT6seVKHBGBkAK7uk5+KvoqG52x
8UKclVP2IMr5k9tHIC6M7RCVzSaDNG4E1t4pk5znrrcFY2Z1Uh+RZPNERFdIcAv9
1D1aQhecq1Whl7+dsALCYeYhzwbrzMlDSRh0r5iAkAfF0s/ksdKdedAdnXrrKzXB
9nzQKs2he2fM912/8Fj6LEs/L7nISd9F50wKHNoh4eIFfpkJ6Ss0Tk8c1S/s5J27
RMpv5F+GMDGbgYVghAZ7d3eJbbAT14DT/k91XEwUmN0bG3PMAfF/KTWpRCwSjmm5
bhKxoCdmAjbDQ0Pq2RYiLoCEE3HpGP15B+2zctT3+5v3NwmP6E7iLuJwvl1WdGrz
DHD6bTGscVfYOhhUyNljdkmWd+bN7aRryaFWmat+bqAqOCfTws+Ofx3nXaQ0RZSs
WsaD/LpxKGIfdeaLMi7GGrUiEmaxLrybXGTiKVAyrOJeRJbyO6VaVzBjTEZ3W2gx
4tCFfSdZv8vI2kTfVQ6peM6sUMrRLBFZZNsMzMoi/IgzD/ilttwPHrgAomuac/YE
6fMxMC6RtPfM2gM9oCxg9Xd17QgWFJzxobdglS8MssQa2xIQtmOCF+TonFMbQqSl
2w/xNTEjhu+5kuUM2pR79jLvqsIm3xIeMCkxF0HIXihV8bqCqHmWzE0XDl6n265N
ubPfqxjyQ7TfxnIXlxaQdGUDWCZeqBtQPlWh0iG+sdZmzFweyr23EbaqIygRCVII
oXRqMmDZQR8xsDvynfIo/4FsOho/LHrK35HM9DcuGs4psW44is62YX2WAss3oOA1
bBrE0IAsz8bPEAOpcMlOU5tlgLJH1mMcWQGZ9/z0gmC2MmAHZJdZNIFCAwVgC5QQ
OMXOX9ywOvy1pnxDaAeZO+Lfy9Kj8skBoGJMPfNvZQfdsgioH/LMeCfzJ/FJp6kn
kyUE4oT9n/zw5RGSq8DQpcgHy/DMYgmd4OPbkfLtT3psAfu4RJY+9TRbRAon2SyL
NOM+YgVpeEfTMj6KI4j26curM2Vj11MRXlNAdqOc3q+2rLK0gnyZtPw0ExN/WJmj
3hJdfpBtlCM/tphqGs7Z0Y1t5uFSzSiT8GkOLlhZiG1RKusWqMpPZLZfdSA1Sx6T
+JrEZHdff05sYfpp3RPJLnl5SvSioPqVK5CJtpmV/1Ae1wZcan5af649C2ROvb+z
1RTlgRBPoOWhXNtsb1YaK4gEqqP3U+q60ZAM7t5GnwkieZH9ubvmLFuIyElspOBX
3ApsCKmC3jSJOhd66CvDHOYBeWpWDwMXgyBgCkD9JX/irnqEEDW2r4tBAWcF0dQu
iWx6HkUOL7KZKrQuICFYA/TllGORbrghXNltiJTV4ynYBsjcQ/xaHvT7eUoieaOw
zvl/Ws3hdKx2lJytLXMI71UFWHLkewZFxad5NJGs+oc=
`protect END_PROTECTED
