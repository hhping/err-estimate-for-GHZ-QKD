`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98K7CkuCgDLeJf6XeEc6KB6+uTKQPBvbdhtiHxXoZW/irslqTon0guDRriWC4f37
W3nFAYSBc21KVhrNSHDt30IbHUAZyfU+Hpsr0ADe+koq9tNKP814o5x20LBHkhEN
r/o3Mi2INFJqvHLv4DVnckUJPefSGcagBJq4JSfGM3zQlxyvBBsoOUh7UeLiBJiA
WrLgl/C78eZCSGw/jcIFbytHTYJhDgDPFsAy0DloYJeaHL7A2Ll2JS4DzGJIud5X
LdmOppPI/sJ9NBtXQnEOWdE44y1cGGKZFqzSuFLkLF5lULZBvWeyBrcWW6Us+8Xa
2mIlpOIYXUIz41+ccvs46baq8p32R4EcvkL15L++uUq7qDLajQkjnTbkH6OPmUfq
LuYUqEhtMmhGFEmqrvrzUxP6EjYuqXhxA93U/YREnwgC++zfcO11JZ6cMxKHRzy7
gS0yprA8kwxG4nCodgsdWDra+61jYrBm1RtU2VdfReGFzK+x7AanlNMNsH08ssD5
ggCq4fALFjs8IvU1r4Ujw75s/fmbJmmnPoIt+6GZgM2ZwiBLvAI4CTPUQyf+xpYh
ksNkUk14RBgnuUhigYO+1E3qbZ/WDvYbaaoyWi6KxdNocHPnFDr8gQg7ri2MT4S7
9ZJOj07LBSZBmgtV3OUvGaiKfZBbiFN+D0/8WTnLbDaz6y2hWt1O4ranCupGRJ+u
xxG3vEall1zM290Bb7SOVQ==
`protect END_PROTECTED
