`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYlKB9hxb6hqotNJqHX/FrZS+SQFhGsBnRxbjPuHrlJULTuX43UmYT7LKuJVX7fY
4XBMDOFy4mzc4Rj2G9iakN83te01rlF8TEIrn4Yq6jy7odsMt6K5fj870WGVqxtv
iNMlgvtQaHkhHuLrjwYx4GClIGCm9MaZD9Yb6Brxb52v56Mz0IPKbbdUy0JaMSG9
uKTbYBeRgK4ed1k6OyMoQ85y2unDFU0ZdNUO6iS/JioS1MkCm/BEKScXY8bIc/l4
tXb1Nk3/2/xOk5Pa+E8Yk4/PNoYaRK9KrimM+xtuyxw4LSsdCa1UHdrqfVT59KQ2
RJ1IuFfv+2IYrM4I1eu2/0kcj9HuH7g6sBZ1tsODR65/z3rNQdjzP5jVHj2KFECk
dfJvTJrxGB6j5ZTZEu/flu7R6BTfGnbkHIE46pRgcind8RTKBVEkVuahAdlVKJL9
WjABjK9YQSf0p4u8BZR5tI5ws26AkwXBEA6qds+reGm+N2Fwa6r+mh2al705yKm3
kGbUvlfQ289ucGqHWju8uJJ0megPGQlfXuKydHCYtsrzi2lFG4gjbdRzgK0S7X2+
QmAKUVRRN5XUPpjYScj9N79n682kCxMZhPKzmSs+/8RKNTOt4qfpIHIg98RZfWHJ
La+S2eOLpmnyI+64AfwjykG2gGKuSXabtyK+bm2gJFFwTtgVXWubCUpquZ3PGwDJ
Fhva32I2s+emRjl1j73q+yNERb/LIzlATy8J2+EiZVmxC8G3CS0D84qgRLRnhl/c
kQJXobgT25FzTyfHh1beJp9054Y0APOoLATNJJTg5cvtU7VJg7pLDF6my6aBexhl
qbMdE991bbYD3o9h52B2E0WItZ4joUb5mJPS+S48OtUqrVBqrDOKTbSsG7LCSwMW
F6xj6ZXDEicu2opMsfRo5djGlBrWt3TnHhAXKE8zfXN9jp0lTbe6Ll1jCBTl0Kb5
Fhq5zkZ7ag1sxb9vGD/OgX2Z6v07uakep21lhUx88y7fnHsDTx62fHd7meJPkrJe
O0++yN2dxYF0SYMWbu6lDOeauR/0ifOC5Vdx46a9Tz5c9aKmaAZsgRGQcorfyZEZ
4MA8M7JTz9D5ntbZEYj3cMNwKIMD0eWxr+O34rPAApdUx/XXSZU/7PrASDi2DQax
50qQUfCrpUCQD8QajBwCBrpSb0ZH0yB9jX58FX1JtOmTDyrvI4WsnQcUp1pXjaJ7
SWm8KH51m7CttgzAYsqoiTdBqI1gkJUwVKT3hfGTUngP4E7GdFqmMSftBvj+8kHV
XSGgRfHHMHycU4xqps9oyF/Z9rImINterNBxBM7pAk7R4TbUOscgncTd3JhNS0ek
5TJHfMUXiqV4Tk2svTsS6tF63c95+jj7ECmZZCjOMWfzxSjq9ffDMUCRktvtWNpK
0qRNtGEDMLjnh2ikn1E/XYuA9S1JpB8gUpMEmU4tof4D4lYRuoadQVCaLr1jJl+g
qiWqCgDP82HiR8OG5AvedVFHcsOnyYge0F0Z6OLABT979c9vhVixtZOlK1dYPUwX
U4+TdOn+nE6b+fTzgWvsOdEx9jiCVAVwhI+bw6ozu2oNN3vrzD/oAOKTLY81Mdea
P29gdolvzRZam8nzYaODiPJk8BF/dkRyw3nEJxVffMMEc1MhBDxXbsoDt7/C+b2s
o2cum65lpb+EMxOGNFlcrAMv7/MDdaAd0lGRt43bcuV9K2BmF1Ste3bHtLM6YEOq
9yWCW2bXd3ZQ/MqQpemMlw==
`protect END_PROTECTED
