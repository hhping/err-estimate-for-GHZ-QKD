`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgv0LjBbV9aKkJFAsYDf5QVs9L8e7SQV9Ph6iVaiBDG3+y1dcMagr6Y1Du1g9Y1S
jvplxWvg8uBU09lmkiTkaw8/hl2xtFuW4+OtfkgIKwhOWn3xwNW1/LOGNeiGFEvE
gKfhZmFdYZ6DOIJjggBk6qrtVnw8tP6UiijcbjR/IDc7r3Ww01nQvstUcW8B1UcH
7G8xCAXLEdP0/KA27dw6iCgfb2uzIlnMtCDLW8FruU/M8JAbpbVKj6I882F/4KEB
PkUsDsdGr2PW2ASTzvqsKbtQCxP5inERyhNLyaB5GzTH/NuBpHUow+0EbKWjoS5R
3yRU62CGSW5BoQOJJYCb5QWcu/bqk2ilIP+9cSRvbOrxqCDbI6f/h8O0Zor6C1RZ
7g9zDiQkOfD8COajnQgvCvhXCsNcQcZPfmIY9HKviYsTlAX4NtdHBr3uquFUagQS
Q6ZAsZc7Mg/JNsAFf6FQ2V+5YdixOFeQjqeGiMKbOCGMHZWrXEHUg6Uu2h6TPz4B
7m5+uGVVEzYTJLyfn4R0siw1n79gm7W6vC8EjQWbDcw06ttbYYR6bO5p6M4adEvC
wezgK0zYlpW51GePXFm4ixHJw5BdQefYVoZxf0BOa7sNF9nGf6Xmk/y4cFIQEkL+
k+FEFpvwbVNACeAp/0EN+gOXzNLQC3A0EQNVmjyxq2tnW7c5wHglhM6xPutmX9KJ
pJUmyLZ6Jr2m8Ix/PId0saSi+aMFTjpkq9vvmpzgMGQX25RWizWxIgsNIwM9fhTl
yczxDqoQ0/vDo4MfrFiMFQQu3OOG1jLm3VuVfjyPUlHmbYodhNigRXTGaPjt9KbC
N5zlicpv/wRZh2fkMM1jIN1bI+toj1Pzd2Ug4C1SUCT4Wiqpn5EdBOAjvO+U0Kxq
PAaulNPGh+rTn9VEF/eufQUpR1muZ29GLXYt6O+h54CjYjQ7rWaKutiMXld9/QZa
QXzozRClmqE/OYA5oJF/dhl0xkUoZwRvxtxWsPkjngHeP0c81e2+HmnAgaMqODBx
uBDvhWW6Jqjr2FVQyag8Jn5NCTrYF7gahG1EU7BMStCgIUqu9HlgLspFBwRO35FK
DZCWc+iZqGdzYbVArMMm+qgMVnPiFmfi9acjxCt+Xc4mwSB4p1ioryMxl3EsJ9f8
ewJ9Q4WlhXE6HDr5sfe1NjxaQO8rC/qIdSbbdn2mYTKs9xEZBJj3WuEw6KrUsiSx
cQr/JsxEuyh93ax8WeAVE3CRPCGCLTRPOHXo7eoLQ/qv3hms6p25jMNlyBSdwkgZ
QbGElz3LS7rg1gu5YmPuBL4RK59D+dcqn6kCQxFG4TS+zKncaX2+Ig30Lxy/CkhD
90RfxKF0E5hJxHEbZZK9DdXeycDErFOn3niq8zSpRAvPuWtoqzjUfYsa1pCAmPMI
Hq7SSYu8kn5RLl2rmlaG4M2k4JclSQjRrCBTHujPQjjEexmVBVeIy+7XBSKjF1o+
dEOPZmXWvX+cI0duYB5WXfX35bwpDIqx9HdrSWGGHy5PDu9lDikeFQOFiJa5NVBV
VpyfKCpSSVxmhSIb7IgRPg==
`protect END_PROTECTED
