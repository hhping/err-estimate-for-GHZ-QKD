`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/KEuhL4r3+B5j/H4zdp8ZcJWgFKuG5N5LIfGNw+zJhXD+P4tYA3m2Z9+CIeHjmc
42lhps/HHg8VFR2x5gwuBZVQ0Sl+4FCUQCpS6jQA/IV+pbMEMQ79UXOtaypiHQTR
UqW8xLpGZPBXeZ5Xg95Cf32w+RxQrIKOAO2UWLzdt8qo3uwJuAGZJRPxvst6bSlX
7zVlVRiPGirntAmiGj7cx6/Asufz/X1EiO+uUduByHfs+9WM8ZsmMY/4G6w1Q7Ze
HUaIFYwppDZaDuUw3U28cDHxXv8Yb5g64cGi9HwJb66K30E12V1r8d8mCf1UXZp9
0LjXagtP9YaGjtxACGus4kzEEhfIoxMN0sRTF90ncQ0u0p9+EfqrJBlHvglPJGX7
d1SZvnUzpdzqj2imo+rTx+3XDyQtn1l2kNJHgyd3FcT97EOPWxdsi/YxbR2JbORn
1lOIS8IR6Ul+Vn5kVTcZvf7rInUkCKb016F/mW6k+S/X/G5Cur9pzD7aqh8Kul3t
iTjj7gjKtqXRs4XcjBRC0v0gGTr3//SsD4POUey1cGj6wzXrICORpd1Lbwdn0Tqr
q/+aRLmwxgL60KCdEVVUUG830QyA+741l8XFZuA7ThZInQn3uaWTD+FNNLGnoveN
80U2+FacaRryTQdE6oeu+JFVzRNTdSONn21Rb5C4OXbXd2DjXgF8TZ8OrHhOtW9r
NWG84hiwjNrKz4ydJKCZJbfdM0eblMEIxuktwLEToUZtd8QA6KW1OknD764MMUrt
bQtipflZIb29puyZ7JSMl8cGe0TLPuSo03CCn4myJ4ysH744ddsZlHTPjNqvFgn1
+dBiU5SnqJl0pBpZlFRpEDgceduY4ohAWnZKOK45iIz/Ie/5bvpLDtZiC/va1+R5
K9n+tRFY8yRqvpFeYdgJic8/7evHZuSr00O5GtIWQ4OzYxuX6kUEWU99X5UAZUMZ
d3LVBGEFkeWe8g2W63z6fidTRDx7H6ZMnIKJM+HMCz9Uqcfki0aEpu/zYMLvdwiJ
zmAdr6NNpgXl4pUGSHkGZFHE0QB4jLt1yfUgnkYDWgKfEf2Z2NDOL3o9ZUfTaP+j
aZ6ohY5HXlXJmQ4B+QxRjElERyawygDicaOw1W+YMtBIBHElH2ePdeshaRsvydHP
9EGjZ+APP8cUDuWCyvzZetOz0y57F1yCfd70dHI4YDXhzvJTxNTy4IvZM65gReTo
8hRaS5HMNVACk/vkBsg96V395LfQ16hUt9ut6wQPP9TEMycj3PtLhZjrMBcQ1L9+
cOKLqtFJBlraIq7AizliZTNqjEh93SNHJQ3h6NEGTfSIN7w8ONLcvhgJJAm39DdT
uTofJL9WEv4En5r4unyADUy0IlOBcsEk5T4wuiNnZDPYpe8gvn5zGf6Um9nyV8JO
4ilqbShD3XlZvPQ5vfzn9eOydtE62bkgDmyvsmvjgo9cOwYEGqCTttN8hDqqC4yb
pG0xaawOQtOIvXTD9OWc1+bmsA7B6nmdYs2qdVmedV4JG6BO45pdt1Jrf5PDYbaK
JV3eEv1/A9gyn+iqrJIr+7gse/o641ws/InWzuXadyiImjUHDlI5TyByV2L1WQo7
5QZY7hvkH0ZyVuDo5X5iBFSDtHOKhggXfNqUAJ4HswdBsRph0nFFWGW8v79AounU
RrnxGsmsFcqZGm5NY36rp96d0h+BKCygUkAaFP+G6kFb29aZPzyfuiY2ooSzr6J+
ecpSNquupdpwXIonzhz+HBFUAXqYqSbSxGsLK/ABxC9A1MqeP9z605uM3xd1STgS
gIl25Y/ciCw/FlbrrWtDtKGppVuz/wj+2hEdco93e/Xh0GHkG3ALd9PFjXvW9cwG
VzcF0ou0Wr/sC8rx+oPVcPkXllWyGJgV2PhrZAva9bKkbkKX/ZwDk61nxRnop8nK
LBtIoBrBNBJ+NmMgi2C0rL9KHngvlaZHicxmJcsSxscOVPf2b/XbG6YZInfrBVyy
cSrHWD1iGP/2EbfW/HhoxKC+BpKKdmGveSj4X2adu2ixldXxrzwgfWLnKmy/qsh3
F8merVygD0iffPUkEeOEl4HpKC/4j1FFdFdXQ8gpLocG6I1QtR2/HxOm/ihryFU7
iUFqF21w1DZn9QUrIKj2vd+ATfshpxJNHc6aU9GjpUPR+WYZtSo4/8PAKG7AHvR0
r5UtTPExGyesmxe+Yh7N7ti1Q2946lIbCuG5/2e3LCCJq49Eo7/71R5zee54j27G
Ji8D7rq7bsmzpObPOcxikSgQJcUEJkJCh7hGcYvw9l5yWUGxJoPgUiJKCzTDS7pg
rM8bWFlZT+7ZWzVs42diLDHYxoXVYRGELAuusngtuWrmY2Go9Nl4Eg0pt3Hdm0sZ
jLpw8HlY+dWp86Y0o+2Q3FC03Rg3cOLw3Aw+qy6fpfQ5UqhmpJZg/O7GPLYZ1y6N
haT3jdG7NvK1Dx49dC4n/xf/W7R3UFn7/OuwNRFpudd9DLIBATLx/i25VTufTArK
zkF2N6GXkc5yjmrym6dhuAm5HsSGgZs3Yd1c54+gkJ8PFvOSUwbOmYENsInTuOTJ
1eSa5/ck/Qeb8k1JRZrWkOTuj7VRNY8ZTdsjj1PfpqfZ0PrFA+tiQ28omPHdN26g
RyZSrKO9epFpZ+REsWhNx8SE68/0DTuemc7gHKyzUlmYjqOthyfYT0+75zoQFnnQ
8ZpstLD0JLDX6WiPy5s+SX9DcKISPU+QgK8tp/+dqNhGxDYWqrMjBcZJWa069XV2
Q1biB5QRCHUoCGJAcukk9a3H0Odn0cZ42lI4nbQA7zv93q1MMPK7smmSu59gWdOl
cqT4Rv/w3Jbc6A6UhQs+j1H83obZkoyjhtoiGfBfJPzUCMsjGiBDPoJm8cqZ+zXb
IEWXUvobCLFIfLWKvSZqhaucbYBEeKUkk56zX6KFlaJUu6A9zGEcQeYlCSBRrtCQ
/9fE+rUQy+LRhv0ClEN1gEMJvxKOlGAdxhyAhMr/QOtecl/tx9eowNHTqXmWuTT2
wBvWtJeZb/dCawcwSaPnUJp2hnMfqxP+ubb6DWEom9a0nzfS8B4DlkyMvPo7Eg6A
S415nmBkoPbe/KZgg/AwsK9lhFB8HfG1sp9iVfe50jPJkJtwemjySzkSb7yFg7uk
xkkMP99JhvEcBAccJeJUuAsZdUUvZs81D5KCY/XLqJBsVO5uxJbSjOvQ1wYhd6D5
/U8flBjRI7xVLhiPJeKDfxXNlrYnnaWEmikBbofSFp3kwQdEKBqy29df3sRplc3t
UIQtY0jcCjtoP6O/VMP1OOs2ToYAXZaa5M39ra3fzUeyLkil40q3meIWfX98rWvi
rAwrtp3aWmVo3W5RzYdHiiWfmpR+d5TPTq0HXvczplyTmnHctlKoH7umwCnO3aES
Y1SFKDJ0DkpRu91YFtkEbWk/sx/EZHYIK8hKqwimiUzUpZCz+5JVXnWzOiEE1CF8
mLMZ8D+9mDmWjczhtmmMfypFGIPm3x2QjQlV11jvd5sh735gznWrIfifkl1btSM5
Dz9nTUamPep2e7b1hmGu5kPeuY+2odlqnc+GekLRGQW3pNszGNsJPVcbbE4DRexS
U5FYqAHwQUtbk8Vc9yMhR/kdbaHrM0HNn33DeckJ9hZcOKwf1xw1qwORRFEJw7nL
qDTrre8+M+Ro57oyxZOOopRcHVWofuXIuayLwfFFGfLwvoavQQhaDEXA06TF0AI5
e2j111JnomfYR3Xv4QxGJjxm+LWnpapAas4s6FDBei3BUWD6kMrDVs70MgldBPZ4
EUJaJr0bBRZxjymuvYqtUoafOG023+tP2OHcpXkcJOY9xGn9HdX1qJBpyzX/Y2tX
e57oSATxcxA3uZugN/SQGwtSwWXz7OfLrI/BYbw+A7LYyYTwJpu51SwCBQxxkgaJ
8lvt7FKTwWa7FW/kjEHxCoUJSymhraVJLkfOfQyn+6dr5mLhS068N7ifDd3Gz4w4
7NXU08DOB1QQuiwTVqaLvFXfHfjnTe9m7/nwBa0w0ftwDK6CxAMPllA+dwHdmvng
6ZaHzjfL3SxERSH4SnAFJ/i1ufN3JTRa8xqcT4IuEIz1tZcAOJSj9fXASddgcyVM
Xtq02bZJhWGOPJV0NcGFRg5ajom534bgilW5WWJzLrpX1XMqjSqsg8TwPleylwof
j193S9QooXLwgZ2eJfV4HU4LeB4Mzc8catrVFoZAEZVnItqoS1NPUiHXYEvL8SAd
jsj/HiP6Y15uRGjR4vz96kWSubS6NDdWkjLpnKs75ptJ8HFK7ic/be+ufUW8oXfb
mmKbjiGvNS3ErW3nHoCzQVlwKSPrtwd1p2pMnRxdfBn1S536PFDN4EUIvfe8rJkd
afgV/VhziOsrlUR5lh+UHMKauc4eWTRq8n3LsR84N0WdXGxR3IrrAeZEJoEREOqr
Wvg30LBqpPQtbdpnnVpdvSQNZBQj4bE7AfmmI3JkpQxeN8rPlsR4VLKZscZo9LXQ
iGETjQHqA0hr1moL5DgKmuXTbgXpVMdTX2RXhjXsGD3NvouPal62oPOvbMn6ZRIe
+FujqehVSf7dMnrK4sixLQhy/zYZ+rrAjC8QQsOS0GIxlAyPtGAny4jdhYONBIYe
lj8flKWe48iZMo96bcfteMKAz9ZAwzKjKuqO2/Ygp4qq2Xfjcc6TazD9BJBvWemv
e4gRK4qSulrC0xkyU3r3GunPVd/jDG3HFVuRBemLYQcwd4SkQhj4CMcWkSk2ycTk
c6odoOA3MYuEQBi5gbguRv+P4M0qjqiIkyS+ub4jdyybQ+7UPDgWXfvxi4FfzurZ
IN6qS/aCeTKJBVnLmBhi+hSeurTxeAJ0Yf4SCjHpBVM3r202fhOVI0kpP1tP4pXM
7rhXXocRJb7f17xKeNZprR9+aiSknuAAwVaqQ/biBIMuCTgAyeCROzjJBmkbWZGX
tAUL9eRrIZcDzQnrB1PLLbGcZFwCAfYRLJtSGKd9hn1WaDdoI+UWbzh7LLY8mGky
mzRbe1+Ty4LRe++d2SGiNJskNHsnwqKwYiZpeGvnkvUukNJdkpAPkHgYek4GgyES
lRWwmd13FSVSJ1f3R9HvgkXTU8kxTDLO97NfAE5DKrla6EblGWJKWSp7UoiCcyC6
tdWT7rph0VyB4iqTT/hTp9k1CLoc/Sa3Ui+QgGSFczaKW17vMkC7XSqsbjrP+6s4
JcAhS2qxq1Cs3yU7tyVTo0zsKF9aE5l/aszzKw8NH+lYgVeJ8iziGK2oLp6g0uxe
d+9iOoxJ3Fulo10ZALfkKRWt1uvSs/S64L0g94E7wAYUFEMj9fOjjiZEMKrxVJqf
79bmkYeB7+BAVZYq7WovX/KXLcpS34awoEvMR5yXJy072MLFhYi/D1sL/G1VM3Wh
7alpgf6CQ0NQIQJYUHVL6Wwor5AVEaGG4rkjJYV/4+iC44k69sQ9WiZYVsSMvKmz
AXzik9XcnrQP6lMJKIpVjE2j1A4F+7xI3zCdGFGN0kFgkcOXbnduuFYz9C0c6bqf
yIe/nbMpBW4Dr78OPHoehkSLlqBpvCiC+c1tZQzpFEUu9fqZv201wqie93aIZpd4
nKlTEoZGTVah3COn6IUAVksgItqKNFlU9+myvy/Ta0oXpgiGjU2/Sk5U2Q6QOjcz
SEKA+QLuJOJOh6/ALZIcIf3HR03XBnk77SOVbm1ybtTCFWAhSZcZM3ec9R9Gh3at
1VMmVED9b/fbkNYUG/KFdoFa38V0xmEjTxYPWUNU8sx2vtw2iLNndePfMFHOrpY+
TWVAvEMZa45hZZL3RzeC630ogypps9xK53yDQPZK1+gz2rfmz+JkbeLQB23clhus
gWdT6Aux1M526lnX8tAa2zlCYsUbHUzWKhNJeyU/EWWM4mlddjiXep56DIhaafwf
8FlhmbO2qGs+gBI/URRkutjLkUi+tQUuzrLNLzRO37bZI7nH349bM/k6E/1hf8Rz
8CkGFI3DuxonLb/o8fyhbRbuXumlJD/EQiZBRuGsHhFWp8nsGFDplexwetnlxkO5
/DK95qle9q5eYz2RmxsvpacU1daCgDxQovG2g3NPoldp/HDW2kUusquqMJ0tNG2+
238DQ6/lhCU7EDFqGSJgy90zmWDN54Z/BskTWC3lTgGQn2G6Gw4eMCVZP97sUh5G
t1xVe7gGuTECkNoYLkNoTp3qqhyLCmnFlclvV7Wq4jvQGzR7S7J4HKALNs0sIUte
ES1HZ91rvUxuHRq0ZXYoBWtln+NyTfax+YXYo2gRuQ7PgbfWe6GEaJX8g/bXJ+pQ
Ybbx2T9OnID7S/luodNJ/FI2H4B+4fJCzNQFa2mQw1wIQn+KN9kM1X6mxmjeHjs+
vYtbq9ZDYXJ9TKO9Ee7xMuRd02cd1flgw14XXP/MstmSNoFiP1OX0VGyjfopYINV
524xd78eHN6xw8qrNabrmca427VUZhCPeK92nWUGIvlfTaDj0cjaN371bnD8M8Fd
3BDScgL+f8x2tlQbSkhXlXmaqbKiPWsd8B56E5xqdLjy3b9CPNAlvcV8bXWCoNAB
OzfeGkSJPeCm3mSLh52jLs0FCQxUi2Z1eCrmNQpHXOLZRtgej2pmY3ux7gQOQCiX
mhV6ZohzLnfLHACfQ2lDk3ftEPhLYCiAK8pRp/HpbQt5EMnP1ZjxifXJRFIIVtxS
7UDvWIoWFlxPm2BVmf+ECAU7RuYwWcxaX6qP4BJLM2Diy2oEhh4z/glE+r0dPz1n
5oU66L/TiC8Lul+jcFIcSCe9nL/TPrAlL5KytChqS2e9txVuTapR5UnL3xzWEoTZ
1ShlggtC/YRnJaztJxttheQzsnk56y6vZsgKDQ0AdLtrqJ7VsE92A8/Kg8h1aXp9
Ij5TcFLyixXZvbQmL19jPkdl5SHb3y5ZBZ07czHJ3+7XryBpBIe9VE0vFSfXA5yf
IuBDwr7k71yCToz5KmycXSpjVbKbLJxtQmQlsf8KmYI+XLBk6QJY8SI0Q2ZMtsnn
YRt4s4emrJxHNMUyQLbPvEv/xTWsDJiQFa1DfGQpIOTo7mb60MZ2etItL/Vi5Ipb
HuuoRayKEI+qcVxXpSYhlDNb7CeFowF/v9Pa/omJXnUYtZ8qwWUXNEwJPdiHUXn6
ouSoUfQKLg0lQPwyK+74f5/jZlWhzqJ3EFd2CRqcWtmXPcE/2pY8J+b86BKuAE3Z
QHlby5uyiBYhGJx47Llous8PovfYCdy/zDj/eL75CRIpu5eSSYRNRZFtAWvEOE75
HOwvb3so6Y9vCc5EDQUXt8SgykG0Lwq4TIw5muVuDfRh2rrH83bYWAuHGF9u3klP
1UFT+MC0lHPvIM2YufVFMCnvyFfDk2SfTrTOGUci+XNlYGLlkIvYLvGDJ7YfR8OQ
yAj7mPYlygBiscEJlmfCFmTJLXxfastmwlJuRTRKIGa3PEwy2XPfNaDuGZF1dr2E
FHxUZFFsp0HJ2eyFUKANjwliD5DcTH0OHFXDj5ZmY2oc8LGyYKPrHyzdbSU7XnOm
afeDM4wNpCPFNUAJ/xVp98iDkvrbZTfwUE0Vu2EjSUqZYDx9WpG5thONZ5x6cgCP
kdzpgghd9Q9u4MfOYKKZiFhtgR6wi1BJbijXpM/V7SE0Ao/7WmySnCnzCqa4oONN
A66ldSr+UQL1CHd5Glb0NkxE/10OKpyyiYn+mlsRKrWcWXZ3MK36ECz++bnSWlP7
NMXZRfi8dt28U8CNmsaccQH2bs/hOuCbD34PBWH7uGUXnIqtXoLq6L366/QxwGpH
kcT/rypcj89jFY7AOnLEGNHDh+vTImH3bxnIR1zNOIbddBpbOp3xGiVWOo2xMvZ2
xrskD4e1kEc+Cnp5jhKxXnDMFwFR8TQXSPdtzVL0XLQknVV+IZ4doALPEUNtw1hV
y3+ThBlX4zP3CY51FN3vFVIKyliUONWfnHzPLtmQVn8wUP0qWKHvpdgknC6hUCUW
dA7fuFODcWpeGDA2DM+tJsZRQaPPS6rvJKhj9G4Cka6IvSp4fxyimeHCOyhhNoD9
XSzfKUSokz1BGA3igABpUuuUQQaPP0p/8MrpqDpZ1K5KuRxC3EIx1CIXohtOd9iM
uuR3QTPUia7gfHH3hL6nsEs5AencGREXq/ddEXfq3K+06ITfbKWoFCYt7AzalRES
y5DHNf7VSCa5t1+rIKoo4pwvJr0oruR/mz5xRb1fW3YNel1Oz3pE8Ite54XjMhbs
H6YHqouazkYWuSmtwJeaEvzCJqR3T0kCttVJJ2jjX/FvCMQ6oeEQCEBv2M9kJ88m
R7ViEbIELJuZzuNLa/YnmWk/CWEdBX7mNKO/FJxwGYFXwny5fa5GbiFimM4bW06e
dLHw677AoMwSypCWHrAsTbA5V8vmIC1LND9ygt9BgYqoH6rj3RnHVSctuWG2T2C6
rMuiYcFl2zg8yjufS8dBB54gLFN+oVijuUp3mwgnXnvXfcVkW+OxdIAWsklAf/Mt
hMHo83K9L28IR+TzufJW1ThMOSIULoxqjQpo7Ip9TpxUXWfMagrvZstYE7zstzVN
nTzOLjef+4qkgZCuE/BD24Cl0PfZlbiNV/jRzr7a61SN6+QSFFouLOiJIsEzaIWe
iWBY7PotDFtQLfMTYwAQQ5M2f6ImJbKMa24En8QITHb6v5mA/Mx8H31QcckaxlMj
OtCw+cToYTLAcrdJn6oGLt+GX34wksaDadDDCOO3UOQi5G8mTifFLRHp2aNfETf/
aDtGNYDVpF5n1HgZcucq6vqsoAzRgtIZhB2VbXkOc6ICq2kJ6C9heoVg0FeXXXAm
p5hoDImWh2ZggC/SICBzQq7WGs27YncXBM1WwOeOlsAiO+8GPDKSFNgwqqGhTBsb
/LxP/erpM/Maq+n2qRbOnOkvl8FCInhDL1eq4IDzR6A7vsmakn+inpRiW7d/neoX
X0UGsUiIXcoydVl7YekXYaqP2wZxkntJp1PWfr/+pqZBu9Tc9iAcLPaeRrVJANDh
OAC16SCjJ7TxXFqWsUTeD/GkBCFX05gK58o4U1wkccvj65e+p2RjJWE5/UNz9XNa
W3klRRjPTYqMQFMfuabIls++bpskeE6D/Gn0UZNyf+olbQ/CYmH4h7xKRXuZp7tp
eSj7GEVLlBfMgVl0agqwN4QyCuNJLr6F66xl+gabNbna/09W4Ll2RBK0WFH9GqXh
tUyFlnaoJSBwMst1m6F4Fhm5tmT5igSjs98ohCTNP988PLV8rBTvrAfmelOqqHfc
WW3frHHToOgvHPZ9uNFhdPgyh1WGCEZdbwwwISuHMulWvWgbZsSW01ZWo97I33Au
iWVWHAXvrL2w2fyuiXHb1MhpLEh6vMo/6ViH4yxCALcyQgBJMU0KtP8rj5YM9yx2
Y82GWHsXIR7TsefZWe02KTKJGqtfISxxqccyNRriKPX4coOHb4rvmdDXHpwBz6JF
Ypm1fjFBgWE2RWJ/cIWyXrABTxsafZnw2jCIbgAQMXfWCJ/s9SliIAgu7ROv0xTj
NZDAfZ4iRnUyVRrAUbU0c33+mi2GbwStuQYW8IkFdDa2gUnpMxfIi9W34BIdtGjc
OlcfwPnnQMd6w41KvrxAJf5ccgw63vKC1wc0pJgdBDvIqJvd4F5uQLGiJ8iBj8EV
NeMOexYykowZDjRlR7w7mPlVgl618a47oO/iasBQtIQloz+yc3cmV+oK/91CVq/w
4ALrJpubyq/83qwmB77Pyrt8wtbQ0pZ1aTnghxyBDzfg+bjnVG0QLRQTu0sHZPlj
E2Iu6l+RHC2CnAcVp/edOu5Q1WEl0rlYogtAeoDzlSFxKOlV/TB7M74KDGGa0X0i
v/8tcmchtqlHu96TmsHRpveaYi30b520JVGVjVmVbJQzm+gszM34Sis33nZo7dUA
PKVxZDyzilXuyl8q5RkpiqVCRadrNMl3xjb1hILvtKJKalhhAvNoRcqWw3PxKwzO
OLpKi/5ZfCy/5zmUdOTQ2E0TMnYozXsbMVP5RMji1CM1kb04RTBmgkteGSX0Y9hX
6A/ng08ftJjNIEOdM7bIysX6VbgJgkSUAVwYTT9HODN0KOKX0T/mhsIupzdeybHN
urzr+G6uxkD5iHH9TIei9zcgzX262j7ve78+EJknnSaH8Cfytl1gilcKl/1hrZdB
DI8Gnt8z3xGikd3TWCTLOa+2xoAk1yWJI9OgM2q0hGRdzMdOZDOHjuF0zKLJyepV
UkBmyTb5qa12YwjcBvDSnhxUpa7yMDPudk1QqzKlZpgdWV6MwJ0GRYrrDzF3uTRH
+fGjQO0j7PXahkIHDA9+6D/3HTqAzkot8+68Xvuk0r6S+92I5fPAcj5O74NJxAl8
GKwue1HMIvbU2lDXC4AQ5t3o1g6SN7N0xGC/Jjw0VjMUYV6zAZOsQs90S4QtIJDB
XbdZmPiC/5ws6oZy0vK7D5VaMl679HUioER9qswQAcJ8vlbiXOhdqP1ytWcvrGcQ
T1NDZ89zkZDSDRX23iErEtWB3qTk30nRkc2noYRqVbeEcVLC85MPPg4I1Gh78OCj
01KXLrXn4SRT7ZfAFZ1CAo77zqyzTr5qZWPBPDbt90uvNMuYOsAaEIBmArc7SGSi
FpCAnV/IMfvSSfodJvpZrXkGmlnle9C/XIpQlha7WcH4OS2DvuKJBWKT1QC4+aqJ
0xZxMHnn+57U/PpIl48w3L6bwuha869CpeqDrOtFqful/3u6fkoY4+BssK55H/Z7
fsEb0OmTXYAzqkLT29abNeOfLfPZwmNGClZIUA0GQkz//oCTyaHOY6BJkC+UQbif
aJzJ9sA3QalzVzEQj+JRMWQaB+cll9cMcPhWbBSo5k75UE1jlzx17q3KPqt9JrBJ
jUZ/IR98esXHBV0GC7M3cfNY2RGnSD7bV8TEs8V4Bl2Enl3KXTYY+qPaPtnriHlW
mx6Uxc7Ss6uWbv7mBmOqF6tCrLFmkwIxwBWHrEqfMDk3y49bpdiRaHjoF6qB+Y4B
QNo1O4q77Z42i1AtPi/+Vbz38+9/Wju0fx3rvsWSliGFc80ZjutYs3axtNS24c2W
d2e36zCz6xVULL6BcVa3fLM4yujQPXHYkBSGlBSHZZDsKTCkuQjQGx9wfst8Mbru
RT75fFOMUaTvNtsL6ikc6nMkDTP0tbq5kWKrkaGF11UTyQ8DqoCFsYP9EnhH5aX4
mM3Ixpxdhe47f+UBh8tCWP7of07EhsXlfFbY40svET9cAuem3xinScurZaE7U1eq
4kksbc61Cjr4f72ckSc8J+rYcnCLOEKJeuEbLEyt4RheztZH0DNFFHZGUX3oc/3L
8E9+qeyissoQHxdc4vw47H0tG9tUTQxkRpj5p/2vyZKRrRUGzFx6zpfM75xp3eDS
lY2Ka4FyG/RBoUTQlJNbLwokznub9100Ug/UauldBSdm/6hZHmFzTcN+An7SgqmZ
4B+MolVkYBQL6exH1OKboYTXYSVE+NmHScSt6mUdjKSSDFQ0ueQ11Ywpki+YcJTD
XewfJvP6fYi1D3qI/HPqIdqgWgnye+fwKcShaxBZeAfBXrX4CP5qy3v5mjLlcNBQ
tF+vHaJInGCyY6TzAvZqj75IfRs7PM62muD9z7HglzZ432yq24RT7DaFyxE8BR4q
R8mbOCwRpVU/OZF7XLENvB6yLfZaIpYxWb4HaziBgvLOJJlBMVJS9yo5iH0zsmYl
HmsUaO0LBOt67DCrVdsBczC8mfsc9mLqzPcYE3mtON5qM7zsmdIkg4oFt7HwZ48I
Njb1jYD/rUZIDf5UF20kMRx73zENhPxG3JwRMppCLa6gg7pcJy5sg/6TirXDe496
+MVe0jgGcp3ziRBenibp6PiurbQrNMSWPN+HRISms2jBM9x5kojEIExdKqCeTlu0
EEEtpNm35SbnTFKSYmCvzGnC0mcvsnXbafo0bpDIW4ValrJcS5EpSbL9OwqRCY/A
+Gi6GPahNwImutUMT64WrR4SHwDOHn3y9sz/wvyqA0kulbUvhhUSH/0cTNVr56h7
nJx9coE+rTh700tY43x55a6xk97MzUvOAX5v+c6UsmoIF5rfYa6ws6pjag1D3Q7t
abk/6uM/uATkOze/IVNh0zXZ8PTDXVF7r1EC9QtrdRcJhqUEghFmL93Yzd/kcdKT
ybzKRVKLR0j/3B9vOS8m10NnsrFXrDfanJM6SOdsSY5fhsCQndftfEN2G5lRfMEb
93q07yRen9Tnig7CxUvap2HIJD0N9jCqPxJA8S/A6FqhmTjvW4xY3tGzO/H1LNHi
QgGxHe5yt8IyPMBhqFGNRXd+kI0CWePy7+Z1usVz7kNXW2/rdXT7FTEdrtkE2O/3
88ePWRtmNjI5THrQQKFrtrgn3ZYCy5xt2E9qzPdsERhkDwU1ttaXDqqtPdjroEDg
xFuJVgJuwNSzBVhpPUphAyW/Pso6aebw3uG40g0qA4O/ONi+iQ3sMe8ZmAC3zlwt
k3iiyx9o36YEWXxXQp8QORfWYM8lIl16jj5FIQrtvTJC9gtNdiNezut1W1t5blOj
+ln3BNCpSQS2H8TIZuVA0AMYZkYwml3AGtJFzn1VyHJDgUT0Mli+hoEFQq6CoCVx
YFzKDEdeteRK+neWtICl+D1HJCYE5whlMDoul5+i9LjjJmuBFOx1lFi9tEl5cpUn
Rwh+5QcppOSRleFloWZr5dX9eCh4IxzT+3n8jK6zwrVNlCYxLd1aOIrtaR8bM+9Y
gjDW3e8B4l4Zc6Djb5AKMSh8A7wP4g27Vc0MHSO3QRttV9BSB5ArcELNiapv+fW6
9la7VeRC0Pvnd02zNhys45+FgmLOI60TyCQZ1W111yxIOt4SwvL3n2iZ1/JbOZ5s
lKHXFAuDuNfhgI/Um+7+86EyJhA6iFvVFmn2ke5LC/V3NtMC0BcpDI48SA7y/hS8
C+33uSqaKXWeGi3uJ6Ymls+lxJAkVT9+nlVRFdgx4G7fi2Rpm3LUQ35QV1YZo+V1
GCvKWpsmzJDFcErThUZzoxJHDLulSY6IQ0lV3jGNUkqDKpHjBz3rsxQR6O+Qy3/5
jBWBP3J6zrq71Igrbf4t62uYYwx0buEbQhmFRZdQhxCbAYyuFDig1SjejG3lyVjI
AW0GCuabViLwuuZOSIJmxgga4uF65KHidSZJtTRgRYcj0+De6NvC/taYwwMXB2TU
OQL2BLgbnpRn56dbzT/L/OBmqo9TPQw46oL1JVorUjD0lNm94uUxYtnC6Dn74592
+y1sv/bOfZwIjBBPW7gnfVBORsp1yPtqPxNi3Qj9Iu7p7B9WukDGa3qGkrf9Pxk4
sEtuaAimRAsctumz94fAk8P7ayq23JH9/D12zrSmhHIOAYIs4yrTp2kpo9JO5WRI
w7PqkprG1mm6+cPKezKWwBLwhnRo+0xq4BuKh3t9juEduclu+ni7xKu33qUlFkjU
h0DTzSl3ZRgHoa6pVqT6WE/sUdUA8Bhhmu27tAv3yaQEBag0kSKPxCSzhWEVsN61
ZwrL2dIvYrepUZcO4iGXLZtudVDmtNrqO6lLsWzGt1fW01S60908S3HWiLhHiFnx
Ghez5M7N6cx8P/ALoX52Rriz9wRiJP0I6x7uFBmr9jkxMMnRJcl2zRtq6GrvSYmS
YCIxP7BJrmiiws+3lks4SuQxY60lyNRN8V78JP7IvLsQo+JJu9yAciO/KwFNvmcI
DOKVT4hkPWAtu1/uqEZd1UBD1RGhM2AwfnXf5g2yDKooRKwnIa8xrq53nO1jfar/
EknG9CQGKYKLtq/Qc90IZJGg1sdliuSHTuHy4X3cmWAeonkRgk3lVWn2smTOPqWx
4NvlmhOZhsvC/QneWxcztfPolKP7q78HfbDctLYmq+jDXDeUgIr4MFmGsPhVa7Dk
LhFmby6DzkxTjAqXCuwsr+sVzlFsZsalMpZtlKAL/ddheUi2qja6IRhUu0jOElNM
t1ae55exhqOrT67YqptLKslPSfNluFifVsoBZzY6YCy8TAavzp1A301FBGfeVDUz
ZcZlfgaAan6gZvRI3p/jkDIimO0gMg4YEd761oP4pNZZHzIE888GkpERgewDnc9P
UMnKzAAf2TzmaeXimqo7HbxqBKy41tZWy7ZYeVv/LAZdiHJ1TYwvx5RpPj5v+lW+
J25faxRR6b2sqPytTNoJax84mqX6HXtHyTNVXwjHxNuua/LFZ9BktB6LGraVprGN
zX2j9Z7GEnmkLfmEB5ZacTJ8vacaemwd+/Stl3BenjLbSMyhV0MqwPnijwhDOH+7
ri9P4S3Zn2qr7qUBRI4HspMuDKmR7DLHyLvcp+beqd4xlJlfvJQJrJ3l0tR43xRf
FwJ79EAxcRoru4QZPyH2dsi8M4QCWvL5gHeCnIFW5cz56xINdBhbb7KSt9UT2N0b
a1RPQRJn/hsGbHzyJUpYWkd81xIyCQyoAEQMAIvNP+e2AZmm1PKcsyTW2vfd7ViW
KTb9mhmymVUAgQMFUs3O7nOmFV4YiKLlI2jt/X7rqDO9je95QP7ABCarlJtbR73A
Sk7/hJ/d+EIKCDy7osCG0oOWtvqgWt2bFVWQsL+1M/Xz7Uo7Fpqz+2Z01c8j9pnA
GK9zywcCKpACPgmCYkNyjdWaB2aLX1hEMmr3s3OSV1iecJlLWl1fYfsZz1bsOAzb
ewKsobCc9LQnFRCw6PE6bvDiGXxa1DU/6nEPdyLiRCMVIGWRbFbZ1NbKBdIu6tOa
CyUw/b4V2Q7+LVvxxrmovOBnnMQ9GPpY1C2gnhHH7rAVMYVpel2AbgnQUfRu73R9
V7FY1DhmrAlXJKgTH80CzQ6qnRacXXscYEN4sBeTNC/i+T9decbcxO2wXy+P4qsP
J3ulphxSQcaqs5dmLJUnAz1D2lGxszOxsXBP1N+3Hxt9yLh+bD3mKI3ux+Rcf9qj
zwE4Yr+pF/io4YBdCuKMDrQNY7ofUITayscXGvKg0/2tREdC4icGUH/gqYXDcE5/
V57JTJd9i2PmMuuvAZFkBnLvV5n4tMfigJTkWHX++dz8oCxR+J8NyVNQ+shmMiUg
v8tcQq/PZY2ExVmd4eG060gJ98G0yVPqOAQQJ5FLp3dVHmt1/cbLBpobCiu1RKvR
vxA9jBvDfTWUmUgLEgsCQfIDEXW/mzacV2ns66TfbGG+JjhsnbpikIOt6m/QZ0/4
+ZnWoDnGkuA370Jg9QmqDuKQBsm7C1e/k+XmHNmBGXi7j1OEEAjQWfb4+r5d9NoN
dnIalvyFwcYMtk3yUNhD8ql8rjoznGIhocW/EOZHq9HRgdhysTk9195ub7Vakhri
M7gyMpmkmo2mqdeaXJOruLuIDj477CPB42jiAWDRjbyDv/V7tjMoksurBNoamxFH
Fq6m5CZVJSitmTJt0SwvUXnnYQAZ/eszNkO0JbDOEnRsm8v6bojD1PWb91Dg9vqZ
+UDgHI4Jkv3GHQuOrKQTeyPa4jufHteWHOwX7PJ0RfVdNw2hlRpAkZKVueVt8CHY
GqrZ4SbXseu0sQyQn29B+qTLY5GoR25QYUxyKYID7mOacAccit4eWaraAtMN/U4C
hpaurZmGh0ubB7b9+Q2y9LiGvhiAa3xAn52JqdMdltrq90WkPz4jSe+KWBMUMjea
3MwOJG/xPjO4EqogplJbUJlkLTEN0a86xq4XJfTNEaOv5j/gKTi6wegiz8gzSLYA
1EbEym+H6aL+6OzClZ/0aerwGZbsgr5YnjLsgWApSaU3C/SiVpcc+QB3I+8P+lwK
8OYZmxBGQr1FqxeyQvGcZnZ+jGpq9+LrWfVPMvFXKLhNdiNkBxP9MNCBj81PqlUL
r7f11vV4QZi+iUs3ERDNVYtqjG0ZZQ+ujbQkipBe7xHZ9roAxhHZTTocBVBDSTkd
qQcFLJ98A+bHs+T72RLL+R6n9UXFNK2+otjrsxJik/eNxHTcpTknKqZhmbInqzN7
VTy7x/sWeJ7pghHGvNB+VVIccTkipYGfNs8AYzrkU31h6UIWnncS7E0s3I20Uopc
IIc0EKCWPQPd5DChOHW60x3TP2fwwxSU7gqWWRa9oEvU6/8wIRoiFn9BqCR3lGkg
TLiwKm04BMvgNPawizz4wUddzgIAc3JY8Q2+A2VW8Aru/yZ1PCCC/KxK1hFDAoP0
i9vP+C5fFfwOT4E5evEx/tV9bjpHzo9YwisQZEgo/UPvcAUSQXUdC3TrcNxwrZwq
h1he5BCrNyKwMSV9EwfGJVbS7SuZb4ZhMq7SsrKifNA01vl5KwMkWZfOZbYig2c4
9qEkjInazOhhimGBGGTqxN/krSfxfjMZy84601yo481Me7+0mpBcV/d18sUAACeD
pIP4YRcrlvegxeYRf8KhuK+o5aC+6gFV6XEz5/1yalx7LoKn9pbmgIUK8baVqslm
HXU+Mp+Hx54Dml8md5ulb5tldfpNR5Zx/jKRG9JL/QDleoZyOO4PF39+Y+doir5o
cADyBwi2n2B9puHAGznqXLpElvSISfpXpHeB1lW9DMACXK51p11HuqgP0pcrShPN
8PHrCRrjAr1AE/KQt4g+GQOyKWbFSA1Da0HdJDyOHo+0hTSoNPZxk8Kmf5CamRLY
mE/UlS+Fsj36brzIr35bV1sgH9eLb2WcQ9MDN6TwDrtJ7/zOakxpOvU87lyg4IPR
t6h/+GiGuZ6NbrwxURg4ltLqBw/g1HHWPWisSG7aj2rczwFfGeKnnkcJubGaVPjn
H/nx/Pa6YMwupcNnUkhF7MhzrixglIMCaxzirC81NALJhUsRj99g355Gu/BVR8CP
Z5TamvkNyT5il11pczUPNsyAl9Ghv/4CIQWDIfWDbhDShJFXhhUJEJpJwH/5HnHN
jJB1xSdtuo8ayWsCatF+rpezihHn66x1klmXx+DEY2Qi8sCXzn/ozzSbKet5NUqz
+v9Lb0Ot0JWB0f3cyJkBBhk/jXPQoyeWn/5gs8HLvvL97q+7YEDc3ZSKFyjIsN61
n7LERNWWyEwOI87+XEU5EPJ2D9KM9HM3XISgjHIW2xY0LL4UGazqjwukhZdZnZMY
pfw5C/K0VM1mE2xmgY+rCjTzyndQpbCG3KSk3Ysv24sd+RTVBC3U5gnDDNrw7zAa
uQNdNqYjsgfETdyuR7xJJiMv/wUl92eBp1zUW99GZDIvMMLz8+caSJCnSNlm44x7
fIa+9GGh3+ZvxuBADz0N/R+kWyuU3tvATTqgsfvAkJ1b6R+QZouVgmz0m6oJNQQE
v5wVMavZpeN1o6xMhdzOWMkM8KPQrCNCNrIMhdiACux5PZxpJR38uFS/mF5bXWFw
dU1Pl3UJDcXQlPYl/ObBHGiWBxYpVBBqN7/XfDL9oRKFK0TEqG1r07RQgagW4hc/
HWom77CnohgzzWbh71Zi04t2RIm0HsztqnhFnADyha2RBRWciUdRVaHlD0Os1bRF
rFvUyx+JyAVqXH79aNpivsK3PHUFLSfmgcjfvA3spTOBX4wqJ8Y4pCvZqKHDWdxq
siqBl5Wn77LrVlVnZEyUrPmmcKJGRd7P6QZLd93pnKdgO1lcmRw8cKxcF9hvdgjH
NTsVW1oFgwPSmsHTaQsD9pF+9XkB8phpzlF0RTew9usxBrroY+mdujXwSQVffqIN
a6B/T7e7hpPnqTtsc9af/xwjTZrmgcGZNj20uMeelgVlIJiJvUwq/fRWm+r+sbVs
JL/pDCe/TRsNDXvMmnlXiOyRKK8cf8PZw83vcN8mdJwevUkCPIKZ8shvcIdf9tFR
YJ7GQtnufjxOm7SWmu2kVO+47YY9+2X+N4NUL9qUexGZb+roRGN+bwDvMl9p9yqn
zNjgq9siPcq9E/1+DJtgO5Oc/UEEfbvHOSnFyNM3Rwg38e9LSAF1mEwO2TlBDBds
l9yjfERWiAnYiWuz9BWezvmczs2nVkNjNupv8sHtaN/cjhy5x6DRDdmWnEEmiUSm
SbfPH/gyRmOzgeDEoO3rDiogFgLAvzPkAmxYhW0kxVptGGoYqOFgZqrOMCw22IK4
3ZWB8Nf4QIf7GzBZWYKuTDBCk9jEMHHuzJbeoAqxmfoneS+P6OOh3gxFEXXXP1CJ
OkTZ1ncvdmgm9Rg5KyK+Lg880UDm1mHZppJRGm9T7le7H7wXqHsaLXjuhsWqGh0n
zKHMw6XjLkXSfEbObuvgD2/M3OMoS4Gld8bF/K8etbEJeJSpR397wntyAFVTBHzy
x6OtnijWch2oSFUxeDkJBQtzfiq+2qSlp9JqJHdVrNkNCBynDfjJL+hlXcs37wFH
RaYMx+giCRDcoxv2qBridCEL8Y5MDnrHc8CktUzTjXRpA0oq798oH/GYrk5nAumY
6qgWKhT5LuZYSyle/tKBouxWC9n0Pd6N1FssuAjoRdx5troxnWtJud3mG/oqqxtW
b4GJrPKxfDNQyNnSKWzGM/Ct+NtaOThpH5LebpA1cEwud7mOVHwc8zRMGqQsObRu
dZB05QKHKyGcB5pvwuNPBjrci02lvlQ71HU0H0Fljo3eEMn9fsAOBYQW+bbH1q9J
5v90SbECoVRfVmEgfWun5bttdFZFUe5jLM9qIgSj1+gHEHW2MnrYmW1xJNXvUaA8
UYCOz1NZp7bN5+7TyhgPbZlX4luE9n9OIcRcI9OvqI6tyZP+ho6Kf8Mm2KWtcmrq
/nR5BfZskiw1J026cX7csp8Ggy4FCc5un5fX8GhZzSHHOLGQn4L12SyNs4mRrLnc
b5y0kzGg5njq0B/eCCqmRUZ4pfmUdHQBO+AOxu5EwK6xtKfaMrm0dQB0eGbQsw4D
quJlt9bKWM7T8cqnlk7OtQ1S+/mMdGEmdu6BZJDv91m3cd7OPCxRZq0bSo48gqR6
CdGVA9plTOYe9+UGiYcCz+26HYWPSRY7YFSZCXDbPqAkqBMYhfe1pcaFfXDlrecx
ZFB09jt5BxcuYUSCWDB8z6k7WPCDIxDKjWVNi6v1y1uZ5cMCqvjS6X7iftKAhJC5
hZiP6ATFrM/2HSxR2gqYepQ0orShbFkq/x8eklHIlMg438ZnpexXiNFsLDeaVAID
RY9E0tEmbfMmSGr2bik/8Fkt1gOdtIMT7FB3esZ8Kt/1Kgi7/mX6/QtIEx2iWGXx
+8Y4lF5yJ6wPuL0KfAOSZk0LjhxhfJWc6s2e8E1Iv0huqkxTFJMYJZtVJSb/lgDm
E/ekWlE22MDVH+E32WUdQuzvGXZT151ekyuxYIoZe6kGL15Im0CuVthDuDZluNNL
wdJFRhYN4f0mY1Kc9mkG4BtzszP1uZkd17GCH3ropA73hPosDmCoY2IMQpovIcsJ
tGOVwaDkaxOO5a1R2q6xXe07iSs3O/SmZ7M1lD14hndIdQExd1XxxPEGZiWnyul4
nw4sRXmuDn6lmK7EjQOBrNNk5IlnEjbY0DIoKm+Xg6wrlbHlrG1AYr4grdTkrSyR
Agdls8fnzOyGwJXh4iRlLdndbin3EDpXQ15tvGNou6eZzU9vShaNr6myiNkPITLT
F2O8AIIWFR7I3gzGmcxD54+MkBe/1bscW1lAq9SqlEcLu4z2RvanXDzYOrsWP8HC
0TbmkMnuvV1GAY4vyPvFKejkfqxPyYETzNhUi6siyHtRNDiknCJIqgTDkhKHI9q6
LaYR/dxR0nTtM3UjBstVBBIRuZZY4zhKpVaTIhVjztDi9k4HV5KikhFhuU0nvSJx
BVGHdfZkRWnI3HWA5cLSpUSh6BJp7Hnhw2oG+PNSLA3bCjL7LcLkMtn70g2lsk6I
nKWQrvov3n0L/rIExsmH04+An6VvywsXskO1z1waoM7NuiXULniUEMstjH38UyKy
1dpri7c8d54ynAeJZA/KbJoOl1c84e8p3qt+ZHnkymxE632pHHemJf3y4glsCieW
UqsOPbkhHNmmXDWIwUnGb7kzXXNgqypIlhnbKm5wRJrKjfvfItAAD0nHEtj248Ux
lYTnR5VIdEtaQ5kpOV0Iwp/bCvqWwmRgwvxbVWhrqY1JDGpObO5OB74rwkV+9sYC
f6VnQvd4zEI/UhUsww3J8FH0DtsJxvg3Y2RBZFizPwInVVsDPquLYjC0yLS1ilau
TiL6aTXBlZN977XfPKB6F+kFoUyCeYLP+5dvoB8W+0Bn9faPhjS9nhqiG8bK8Xab
YtMWufaePx5bmGBMbZ0xpSqfKM9zYN7kdz39+0xGsOFWi4IT8PM/h/8CgdUr/Ix7
rN1WjcSgBuLGSpyobYcJEMTEbtJ0JmxhqRRDjank+JaVM1HM6lmL5WKB1bbAMRbW
2WcxlZ5RsJrIlwx3iT0B3I/Z3vGALgG3TDPgNVKCW3323X4TD1BVM/tYi62zMsFZ
pJ4xBPtZlMJSqhJp/hQInlY8RxIwfC1b+OAzg9FB7nvaHD6ml6RvScjx06OnTynF
2Yx8VloURpnxMGUXFgcCvmOoxIm6WztKmoVkiZMBqFynWxtSuCgKO6hr26xNt5DK
SIvlV0xCTWtLN2jyF6aJbLkIx60qM/uu/ggCU69m+ZmUQdy7u9rTnF+7jhokAA9z
dtw2Iaympp4GEUuMGJqpbnXxwmGzuHq8MpLKEv0jfwdDeioRSdw4mS52hN4ugOp3
C8Q3cTPhz+fuQ7XLL5sBS1Itkk3/iozkuARKp4E7MGe8bF7K4xZlGq4bPRZJq4Ue
s/C9Jax1X3MC+eZ/LodGiv4jNlfPgbU2lA5uaYzWYhtSv2ZusuSRfPujO/TRNm5C
KZtKVngyky+OCdyBdYqgjgHphez7yGKj/+qt78MyvOYiq7z2zBqkWmZgcjnHlVYs
IwXxrhxxMlMgibWRGQ2796UJZC1TGhB9HpDm8T85C7DMWK/fyk4nh3btwGM3nYFW
4Azqp0Azs2HBCr4RjyXZCC105M/AFiTa3lamRjx+j0cRmayhWpXBbhbxvnYasO0w
ewyWAJSVmYsbMj1PD/YRqcbYLm459kQEyOaB7edvTD/7p8HgiOLPNhH07oemLKEp
HHSsLWwSiicLBn3EP/AjEJkR7DNJNPZiK/Wec7CkzHfauF7HIf3lhlMc10fy4jLj
h62nv8y+0I09wfZhMg6tlu5L3eZOaXAtBxevyM0J2dBEqltcWuVRHoBGzPV6LinM
s1ntZUhibJdALVaQKurAeghNpLfAKwf/TgZQc28zqy1B0zkdJdAR7TAiDanZWso8
ztyIpTyBBRZNJu1X7AZawrTBandL8TDCvQWlVzSkxGF7aoKOHXJj+3ByrOQwkZrT
RREcqR7qYRzqSf5npvOhC6+TIlAG1dAzzijXUtZBSpr6QErdeT+3Uy7z2ypH7yJx
2Qu9x8n/rmMJq5Dz2joJjt4eyx+YmNJxZt/9DNKnA2w4lvzACEaclGh1eHIbn0t/
mUJV2OXo2riueiVBTLaahL6rcDWB88mXjGhfVhK6kjR7F87gZAVb4bh00c39nOOo
U0zEznOAZ1HSp70xielsf1eb3igXiIedUkA2TWKk/pkcc+eAOFvG3ScdS7yl18x0
NaEFY/ZtmSaBusk/4o9i9DGeRX55fI4ekfyBQEgqE9MNtlcaykfjE8iNJhS2WVjD
6ELdeNM8q3zHg3yXZIkoiFr7UfJrf5eTZ5pp4+pCO20b3VyOrfRoeV8T0abvcTW9
Y8k7BEn0qqFqLgCFI1FYK2nBFuaUKly0FqnwbTHnnV+9j4k3kO1/LDjN+tFZAPzV
RaAKZKHs8fDn5R/90Kg4tXRngxNJK6SiMk2X3A6cm3h/HYrHjlh85gRXo68oDArY
u7evrS5dxv9BiKDt3GUREWp7xNBMIVy8hrKZdghkIgae8q18/pax8ldWywnkJNjA
jdEW6BmVudJ9EYnQDw7drkGR6rIxD/DFJtbFdo5ebkiv7ZDroeYZhDDwDqdSghAi
liHiNUGMpkRt3V2T+EMCg6eZKeuVx7Ddi7yo1ivIIU0P+le8C3rTbPN+4H5Oos6O
l3ll29Nr/ycnd80YKRUBnVvEUL5Ecv6kRxUgNb4HUwzmiwLM8avzkxE+zMVBCICs
/AYeBQw1qlOC98W50OHLS4bFUSbGeZNWtoydods5cnKO7q8wa5V7cKHO5NUyhdeW
A+rwgVU0ZcYcIoU5heyj0n5p38Gpo5Yz2FR2xTHXmt97rEwo7pPn0yv/ogU0rNd3
qN1R2tJpaNILoJVwA5/EDGlaRqykcGHuNhjrEearukOGIs1tODBrzqsa7m9ylTaA
5aT5aWVVsQWJtLBvR4dsk5LVTiOhQ8WWy1roNHHELFRDfZ24rJPf7VPVpcNB0yOs
Yvj/R712ie71Y9X9gJqsOj6fuP1Akc/LDiWHH5Gf8nAiZ8PsMB30bNF5vWDkCeln
hA63ktDPlF1ccaoR54HmIDMExdwVauLWi8690r1D10MADFArq1OHtYFeOMitmx1y
pMfljZ5GpY9kCQlfGCo2BzmyL1U3vqnym1Lyl7PCUw6TYL5fq5OmtrQPqTucjgrs
vOikxd2Yr4Psv+BrQDkOBbCvz+e0wadVD1xzy3omrFGFZ0UjUCSb0Lp7KZ9gedeC
InSsbAcuetR4695ImPUql+F+q/6gB9W+nQaMaOZe5Y3HTON70R8CjEhKTK3sde9O
b9m2JLPzqlU1yMeRtHpNJfssI4DOqCKd74QI6zH4OOiaeg/QswCnju+Zkcvi0uhg
u2U5Ssbiq/n/g9fRj7HLUtTdUh98ZgeQqyKiw7FuWUBnt0SBRRU/S17E89AnBYFZ
AvMO0xMOnauUUzWoZ3VTBB3aJeHBMZYeuzsoo5G/8YjEB/ryq+pcB7uBlQzxIIjY
TaOdnSDSP6rj7rjvIwx0pZ3mvEinvSL/Fdy3wFfYNYF6w8xgqnWRFuUAKzsKG6v2
hWV/nXNvePU5D0rhCfcD2YV5ZQGZLuO/vIeDeHufpJdbXlR6W+WiXkxaho6hqclG
BCF/5xvB9pKqJoN0V3SDJM/xkYs4xrXOZ79cp+VlyGd84rfSOYhGiltmZvOx7Jcl
boM2VE6nnlIgXy37v6IYXHSAwiYkz1J/7aDEEUgiuLYsPoVLN+boJGE8E4K3S9O/
XmuwQSlyJjKkYwqP7yT6d46766OvV7eXgjVln6CRfg5V6u4LnFLDFDMNxAk2DVA8
nam+psU1lSjAHyqxECpkK5nCXHWdhslYqCYzrpbQv2KochuexUYpd96tLhfctybk
2LMjAzmjwhlElxWRnIudjrcXOFGCnTQcESQGMFM3El2ji2ihzSlGP/VLjyVCMfuV
+3I6/qXRkf8Jrq9KfmgYNFGnP9//Jg+ayslbsN+gI4hrqIRutTpfwJnfaPT/9Y5D
SeE7W7WcVnohJ2TkdEmXFkNYC6duydh3vcQNolZhBuCzU9NYK4/+b11qh1jmt7T8
UY6QDxofx3AwH10DmKKXxdHAvUvdHiwunrgt+y+w4dvN/VBPT2CcOWMZ37s4c38L
8JJlqVDyIh7gga39t2HNI6AB/YrEJefTWVYZY5lIUJ/ennAT3MxUqRCoK6ct41Nx
6ImVnFySw15w4mXe9p6oIUGNR/WdqYUuNBnGWBGaWUR9BFzSyAYX9xsxdXrQhXTI
1V6ho+dOWSTfxhqwsGicpEgslEwGUFifV533Ko4bDxxZKS1XX3vuSZ9tEtWb7cK/
O/RhO8aHyPtnkgMUDte3mtVmKuMF7hY0z8YGhkaZKNqnazU37tTFLTKTfQykNbq9
93YDjH0ypkBogVdQpbPkBs73DLpdxmBmSojX+Jypj/RPHbfSneSNEKzTEKDubuFV
CF0Dp84auEtkBlRXvizO6DtmQIjBc/pLM+efvfUHi4rpI/+C6HoIpSD1HIzeg0TR
GqkrYuPmfIcFQ2pTfWE3A6F7O4YzR73+oD5+0g4XN5947ZI+PO7nto1FXplrU2ip
eCh27rXgT5h67XGbiP/QRpk8/7FSLdIhz69wDj9LiirTti6WnzoHCM/YR8PHwXv9
j8D11s4oc6JFLW3yMpxnFx9mFMqlPf0lmUJuEAq9ji2YDlovDGsLmwcsF7a9YZo0
FD5jGuM5mUSQouBwC12G6Lj5afCxMRDdzGT5WoYqxY/CLjXws0B6VruTihEWj065
xg6JU0C+6H595hSzSFJoHSI1UaZRXz41+T6ntBPWZfp3spv+yP21N2Lj80im+p4W
n++C7LOXybSjH+shGg0PoYVcD1zw+Wnd3LAbF2l+xSXYlCcrVFQnm/LWmCldEH8O
ZzZ1KrozBY9mn4Z+cPNTML1DIhpzxqWDNS58WETDFSKGnvz63KhfDVx9APW7/cNp
VJPHt3pX7Lg9y5HXV/o+lvak2n/jCspGUDg3zCHsC7zjLzmzLDQmaQ+H/Mtbc7GS
LM2+redTSuhEWXxfvCnFzRFG+fU80BdW4FU1uMtzbBZcuKTFjiKXYIYFFMzVJRmd
GJ36d+4RgI+oM/qYjUnwx5BA0+QmATJ3YI10tJQnhXe68ELTVg+STOSWnG5A4lNf
k/DGTps2GEmDbrGrVz+BbijuocM9MFH+Z9YTMhO3SyMcUQHOkZUpG77dTO+kPDf0
PU6b11xk8G9Bsmx3+f51XYdk7ckUJ9uBPTRz1BsK5aPO0e0hkHJJMJTtkNfNVlCZ
1RTDsVbNTf0ToLY5J/7VDDgZ8es+MEZ1WTmkm7Zi8Vy17Y1ZFINqoYKUHsGMWyer
S9uXZwG/EIvjz1ZRF4Cd/CeKgERwB77K0yADYtEtox3zLlVDgdU1owRVdEpgHERU
JoEeFStfIn5zxDDFAc6V2N1eqJo1bqtTGib4ZAfUdbFux4zLb0X6b5XmdqdiYcYk
kLdWLiCZHli0RqhHsuvpiJjCn86FNXiZrjrMt247gFN+qyilPex8mudKQvc9F131
1204y2CeydNv6JfYmBhTG/49XSMxkVcpxyIw4KCa5znUEXo5bF8EiA1OddWw4CVL
vtsrk4nojoHgxeb3Wfd+Yo4an2bi7EjU6X8TGgjhoYFBXRleWlZTdAK/hY6AzSHE
8BVPOQviW6tmAI36OH7V/BJkA1N/GKcAxvNzpnQyUMEy/hu2k/zv7wMO6TKq3gCq
Tbv0zRwauMibf+QK9nNI/gy9shWRMa8OeMiWVb556slu06fWaw5ZSIoZWLd68D4z
2nY2E1T/ZhNBmaws1DEt00BhLdxvCaV57yF7467ymGk8Y2xWhgk2IdruRwmwvC7i
UQSYny7c5S1D9erDffs0EPZblDJBbsRhBCoqFrwi054gx/55JLtRhONtQ9R8umMN
5KHvuLbj0A5MwMiXU66BKu3cUop2z5KVgOXzegeke0v1X9tm5uPVmCh61aTW6hRX
W27UrqdSaohkhmrDqG0HlQDGb0emH2P8ars2V5glPYvBmwBVxAQdLKPXlQHEZ9x6
jD7aKm6N+VD4gOJ80BhKQmOjrarDl9Efe5Fx/BFhg+FcVZw8LgfR/tdLtIN1wP2k
FSFej19Oz2gEDdfA5bMA4IjIyzECbXc8CLkgzBcdkhWNUuWOfrYdEFC+/UdxcyTT
ti3M86kGKyLEn+WRUqAk4f3zdikr8SeuPBJ3MQDo9aT1yzymTx+k++zV3oGD/TMC
cJosML89raMIs+9R1ZWMYTo7lnd0jXnSWj3YNc+hPNt44nkk/dttqNF/5z64K+zH
bhegm4nUKD1/yjlBq5OOwQsIvupybeFcwW5xAdTjC+wRzirkXcYFLdfLgniNTAky
TP8V/tIDrRYTOE8jG8yuhUpAP1i7QgOYvQAew+UlWvNHtJ3cLxCoWczkxjWCMaae
0inQ+OvheCVTxdp7Jd+5MU6E4GPKPAQlpEzmMkuyGwE2042TSt7Pdz0gNZP3qEUI
iUi5RZxA/hxa8U0E46zrIyBCoahHL294GZZvYqYxVmQs0/Nr0KJW21o0GUF3a5ru
mjIP73SH93K8gxsQBoEmg25jPBjkuSSUIWr8yQZWlZY8uwXUj5OycT3vH5liDx0+
XogfrSJl3gmWEC0PpSd7EVzOLncZ3YF5DG89OcMAQl+gUrtYnGDqGvQYJ6/hihQo
7T46kZorbjYLXL4SjDuE711CHV6k4CoRfe+JSIbSplyYu962MTvWo/3rG2zFVFig
5iwCTp+1Kc6M9l+mhEB+Uy9opztFXobq9YmnXg8/Y6FSPoizdRJhMkINDnvDxNnB
Q7rwjjnZkclNB7JqT2GvIE7jqPU0IpMgjPj43QGGgeGRTugT4siEkxgAT3Gh7bAi
ohlw7YyPOkMUQu9lfRh4JlLTmkdMqU+h1N//agqtXuoSLSrTnRZBZdMR0OuYatTt
q63sZH6kyQVWneF7odOSYSVF9LuJNeCn/XWUc/61HRvEGSz+G9q1ILQRNEz4UHSp
tOGnMCdG2EskvME0zr+aUgDJVB/E97jcdV/Yoa4EfSYiM/Pxh4v92IyFxG3QEnn3
2XWasuGTe+mlDeybqcEtgI6rjka9iFn5kuAFQkcBsgL4DAzbnh9BS3Z0xnB5JPiC
gVrKSnmxtt8YH9qCkKitD4t0SCU6il0yxARqmDGqmIo0WhN3zzHYQdE/zlcWEmKZ
PDetArofsSpljcdhvTPgQFNgJxtYTd7qtnMjvH7h/UdDQaeS9XZ9YUhCyB/FVApj
PwdUyzIcPIqUBvo7cC9vy1gKeC646p+sZ0raE3Kzbc4WFKC1wvxPZpHaV3+Q95dk
1Z/qfLLmunl+GMHtn+5uzyAyRNYEmLD/hPB4Vvxh8bPk3zVBri/PM3QWWdbimolh
fJ80lnwcyJkHjgPnqIreny1oBUfdvl1bEPT89Dhg4CvgR0RMg+MBrR8ZyvlX+oos
5+txLhbT5hoorBTo/VctE2KpSaVdyzy74G/tyJ+IgZ+qLovMyuV0pHQZLIuixqXp
CmFDQmafsq7XPn/wsiFSx4UGc+3qArWIRHNZ7XoM5ptEZZG2CH9MNqyyooLGeqCq
bdZCwVj2T/b3jxzkYzhBtKTHXfQUne01kx9vSrtM/puxL0lL+enzqtw0Yc+fKy7T
6q2cXWxB4pN1iMUkMiZgaWz+uwAkijsV0C/TV7be4hFTshQD9EzskOyDzTZgIP6V
THpK0jgHmyM7D3KWWWcb9Oh3koY95Y6yHGvOV/SY4xuVa9xL7rxU7yilVKkGvpUo
miene6AH0e+nwEql5Nqb+wwOKcj7Bjx8t2m8Pc13/HVTNhE6hD7IL3vrrI/O+Zw6
i2Pgueqq04DgbFt6tVckFmtnVl0Xh8CpjgRjg662P0luAaWmr4f2HxqYFZeoKaHE
4hdnJRazM1OokAH84+JMBONNfEKFoGaUD5xQGkph0HeIH9tNpgPANB27UTv4erCh
et67fb4CrcRmtcfD7Gwqsg0FVxzx0newwULy7fd33iCjxzVc3PK3OVk9c/sdC6eF
8hXqRdvgMmXxO+ew7Oa8otxlwQNRaC/l6oUwdK2LpnWdPsi3OsQwtZqPu1/khyP3
SjweHXTzqBwAqtESghbJOrJFFOvk0E0fnqriN0gegjt3Y1jN3ch/xjedOUG9PFSp
R5iQD5QG1cQQih6MHViOWWc8CRn1LYGiNFIUkWxOOPZyUqDSQC+jh3zqCFedHuIC
af5tJ4xzJqAbe0+GTmhHl5Id0l2fio4COzeHD06o209kpFOQ/BX37wOekJhl8+Iy
7yyz0ghRWF1VAMQo972DAZ4TqoqFmBdpArdnzeOt6oxJLo1jAT0V+93RSlt7/AAe
AawrQEw8itU306RJDsflUohXg4WHSGd0Tz/JvhACfHiSxEoZcgeybLbjlXbBhKz7
tJvJxPQazdaFPi2re34RQq9yB5fzI0z3ePUCDU1AnRt0A6BOw12SN2lg65Tnp3Oi
h6fe21Xualh6v9k6OXiZeZE4DLGd+fDsnO64GfnK6AUJkTl/Crvxy6cXOeJjKe2H
ps6FkLHAxi96JwXDug2euagoB/MT69t/ZoNrjL4jPkFn56KTYsOXEQXg0BQaWKDF
POr+aTNH6/uudYS+DMNtlu4nqgtBi0rSS7sXP/3AraGJkny1N4IbC8Hq/5F+Laxm
a8bjESZtV4Q/HiyeogvgzJs8v37ZorCwh2dTeb9mbHneudzxpyk+KHUw8V8Sc2u9
YxZrav5wj09Q0spDHiuLKh2MaLkTSMIeEBjp5fhAQXwjKLY8VTWvQpeTsT13QCxf
iwHtboCnNkr4H6Pf48pUatNTUylj7MNBXrm9SOgcaUL60MU/YeMCIDP1I4LtMABo
C2eG+QL4juxcKbmD/2FV5Op3DE+d/E3F7iRGXfbnZdF15QiNSMp2LudqgDb7B3pb
y6JDUj+8Vj9KSZVM5jFjDdmPQ0juKXhSONIgQKAyqOGea/uUxPTBoxaxCblRW2FS
AYJmydERRRJHlVYHfyTDXdD6sqRTyH8Myat828XohEaDbHgc13zEPOygs7YfxBTY
u0+Hj/HbLJ1p9v1mebARXlaKOhQlc0xYR4t9ZAE6+jYaEPEkHYUp9nY/6RuGDVI9
I9+YKgRZ8YtLKSy0j7TvrUFUv/fkdHEUlJn0Nya/ZdgDk+sUe16NAszFHnRuuFr/
lY/7JBt7PeGDEoXnvKyQkOqTQbUEVZ4GsTfcNTiYCz0cPrRh+1xxHeM4OQSj4nEe
NBiPBnTnj/mXnSHIyhOpbMd64NCA9eg7MDUeV7pNFShnLUIzQ5XWHfN2dlVYJXof
UhokOcgOV+k5vuaLSep9koA8htAiHUl8NvkM5EHvJXf6urc8iA/4z4eGlS/p3smO
W2n6erC2P8AyoyQ9niKDAppcMMc60jvszMWDNaV+84cZmNaOIZ0mQvPzdxRkR9NA
E4ZDyVap0lRfcMsbo5hyZnofFRCQMSdG4oMBrDlYGv/1y8nLxYCiqbxvOcErn+fR
WZVTnJwCt7BuAwUmU0hwtZ75CMCdjzO2dJHB64pTFHx3KFpfJMYrKJk1Dg+zCNvk
0LF03FgykY3Xi5ljsUbBAxrQFmwTiOGRko484x7CRvubWcprb5oNqh+g2eOkF987
yqqvTv7TzJzPPpp2OFn2H2TjVAbFqBsdzKXy9p90zJ2rtykTDNyxGJJDk1l/zj/q
QD63ugCRbhZ+o3AqGtG9RYQLFPJD9WcD+yRYCmyBZHjJxw6qzz5jdARFtzExw9Jc
cRwIVI2cWEJvyqq56PCZbRuCzTtCQzMnRpCamKNp4nVFIzqfN3girOcA+zUPg2R8
8m1eDmBvFPZxJFOvSx7vvIdhzaUiulUi4CIEawAnYm1pwxuTvm3RIiZzdUDkkU23
9rRmGhxPVYSMR3FNoZCNOa1CO9WEt1LMH5PoItaqiN4TYyA942N0SqMo68MQqTbV
7r3ZAWV8MQ5Xv9iUUoUorAR6VVqIOfaLseGfapWjJB/2kS9RVQKMP+qEaJNQ/PlY
U7sbQho9tV+d+hRG3t6Qyt2Z3XhR98yAbMe+1yczSKXUzeefsW8zIReuyDlxG2rN
LKX5fic8VnGdsC/cIUX734JbOrKtiGhxBxH6KACXgVkmByZyhqIhrc03Z9syhImz
Zr57r1fg/a9BD5zCSkYjSa3SPIABXbAbACO+eLm71yNz1Jnx/eiGBKqDGz1s154h
EsBPa/b0NpVAVvJZBNmWoaepmYuOKU/hshbdFO1eT+HiO297McAOEB9liX7sKleZ
Ydt35yxs5UkeTqGvSuh4up8sn7BBcI5mu7E/qsg0ppUYA9hZSuHQopz/ohiUeANo
HM29/W6mzMUnu4i33K+1nZpMCnDa/uoQhWmHTzpIeZUtveZFQdnbylQ5v3XgifqW
w3mbFzXrBAGsG1sgB5oUQC/jR0X4RRBm6jjWDMYFlzHj1a2pWLIda5l8wIqz5sQb
WI/sREIOyV/l8NEkFxMjUP8LXRZijEpW9bUjleW/r/NoW52ipKOqrE+3JJfN4co/
l/wg1q7F5RwX62VbyqOdMJ07IobtIwkSWCb/IffRpGnq35kJdm7/mGy5ZB4SDl7a
7G1hiHCP29tCFxqioOuCH9ucIT7GqhxlvuU+IUP9vQ963fJVWh7vyvVWilpolMYS
V6vRUUoR1CGeqdJm8gNjwl6Fo07Tlt+CFnBHLdeWwFXb2RhLHRdZTSRcKLohAHSf
sKGpJD37nGePAKh4hUGafVm02QVFItJ2sitsznShIclWz48uGxEylcH4iPNzcoN6
S9ximAwykKJL0YnPVO1/VzMaf+k1sie6aoLUih/KlJKXDdDHYaOYDKfYqqSks143
iqQf/2e3trmhRUNouVviUEVHl/VfwDJcCh3AE/b4vW35dyUByq4ijx4l8eVM2hAV
GGjyBfZKUryc6KC3KmZlmV83lmrFDV4EV3zv1n0NIGQpIlxUdTrBI6OEesOJbJ9c
kBbU+E1+e3HF1QBWgWtRQQcspvlz2lkPskItSDuNfiT4pMj0eH7bf6Wz5Y4pdOHu
yOH07MktpHgv7tCFCohOgTkGe9wWndtnhLG2nQKmCcp4GNnSwsNlT6pE/L4Kogtj
5iYIHEhSkbFxtQUWYl5pNlm/CMVnv5j3MCMT9HlvhowePEH2RZFb+oGJ2OnSCS+6
vQIIuaaKT9H81RNo83mcdpbjN7y2VzAaME5kWIZDupWQtnQUYH4jSceJcuAX9Zfu
D4ur1pffMZqLFLfNRC3BGanxIBx5bsLF7GUPQPw5mHdM4g6HmDmHMq7Vz3jNJjVH
whTPgr1cnqbf1TKkMzMnVa77utaKMalH9NQ9+9i25/Z8/f9ZtYtP/PEUmBTCVZN0
hIcg7S8A4eZMdR14Hp+2eEIF0n7k9UQozu1UvaU1FwiwkOo4ceq8MYFm6xSP8ogy
RNOvJpukfPvCJniw96z13D2h3pOUCHRPSVCfpI3tCpmiTgYcdFWMfcYIALhB3Ngj
hKTeiXPkDADjFbyfTUo5APerfWdoNczgah3j86lEGFJ3UAuLJC4ClI1bVzIf8Pc1
5U67+xJgSsjqVP0JsEeeEpbUqpj90Ypdj4VqwmwDjTUITCJGsZixQ/B8sHUe3eI4
HEf8qiv3PTEJ7L2vJZSxn4ERqBM+iDMYF2yiWFyNwr5OHCrgFuMmRrHTwIVBWJJo
e2dYUFIoFP6m1XUoYkDkCxaLR+/bf6Gdbobgef8DMgxhpd4VVUul6KoaJhe+bPgz
vxpDlg8thd7uobYjxx699UwlZhDtwhGW6aQoXga/aqcC4EqcYAk217XWB9TxNLzx
0RL4ypxQSjPUqaN0jTpAOI5DUzDpK23i78+POL5V6u9TJNRYzCeIibCzIFrsI7s/
RNeNVmiVK0bi8MqjalMYtUKJ/8rF/BeRXA1Jueya9u2BbP+hqW5bWyVkzzQhuttB
qtxgAW/w0mrhQY2b0D5APHQLBZabfSl+JTwoEVfK1Jd6Rto7kE9egxlsCin0MRhr
gl/vsopYk4TMmi647jBi4yxGLWxM5bjMOTjyAy5p/hqQenNuBOXc2HoSZrwEsvGf
kMKgB5nV4pX5TbJiFK2zWfHUIe3bnQDQSxDWtFHehRu2CAa5iTW5BdKPi5HczDKB
mgh7dUPcJAe8R5UACnXb9H4aeAnBqVZ8K2Q+nUAQ42sUxu2erPIYb5NJVa6Fz/P2
aKqqM29TXE1r0gN8b2W6VFDRa6vEYg/fK7Vh6QNodNc9hUzFY2flzKj9fnzz8aZ6
mxt8GkaObVLjRPT1hFo8pBbFeXY4MoCL11+yx/wvKfVa78pXcPG0lX/MHR9iKeOW
x4Cawdn3OgYkbHj9imAlOHw6xBB61bQi8UU1TWnxJgxWensZbnZ/bMWhrzpPennB
wXJoX6rV89Qgye6VcIvBzTTwcUYmQ54O7LCgGNTVzG8A/90h2XC1X/Gg+K+sbOqn
b0C5WoD4JlamSrOYEchh18cXY/vicVQnBKSAhRGCbeApRA2DBRxQS7qF0vTsT+g0
beWVoFkAnUC/9UoriD2+r38YWal6yr3r3skR1xXt6lS7vey7wXYJjh+5e5tPPBKQ
SFKp2KTqXO+VWsbsFOiXz9SdfsIwq71F9d4cTnLMEbNeB/8ZONtSPIV8r+R4/Eeg
beLLak7mPfSCVti7A7oscKYJhmFpHkEtYjsiOglFnQkZjJkt5lsW9j4kbiXV080M
8AiFBjrYn4AlCh+ZUORGxuP60zWA8sAnOPTOrP/RIvkrElfOF+FDWdR5UoGmFCbW
VKeNgtoR20D3nWfayoHFsRvfTEHqxILp5cJ+Q/sbk7hFVmdB9fk2th6OrEKXcyG9
NwfccLm9ANCWFlJK34ILtT4EzEycpnUHNy39ENKtYmwPcyna09iQBA17ZqDu/bUM
NivGcFkJXFesK0Rv0z8pxN96EXoBLPf1EIg6OrBOPl7undEVMpd6qJEktVl6//8A
iSrZe7+h5m4uL3ri9iMRIGSGYFpXZls2wiEYy6hCwdFgSNqhNPV5nFOOWa+b/t9O
G7X8f3afqEIVSjejYhMowix88RfMeptfp0D1H6sLv1UBpoxGS//9vkzb4wrdbJpu
rNNmSsnLxO34M0Kcu80KEVnHcbpKgSBDyrwfYonNot+ZUlMgqttNc09CWcXZPSam
cW2VcQEp0I7CnqgS1Ujd8eGSkLZ3p42TyOmpH+tO0TVD60Lc40ShQ/RWHore3YfZ
bNZURRAvaIK3r1G9sUbXqh20gSOrY307CSXPlBLU7J78qQbEVQICurWQeN3eXXK4
qjkgVwa41ZaHE9WYgMRX9zEuXC7uveuyy64djBr8d1QSno9KjMD1dDpiUBBzbd5O
x986B50KvIJ/ATHSgxD8eo8fX41jcKg1Q05XDNqknRB+A7vKdMOMVBAFqbtiQSgc
rObpCl15S3v8yhwB1VDqUHdvOxj5zm9Y0sAeSQ+8OFW7I1Ut0xTsDmyxsc/1YIT1
mqVK41KIldzgGkjo9YhkNoSPZrlifFz1SUXqvG1FL4Z8ZtzBkUyAl4dOvEaeplTY
ZkZ7CsmhTAuRx7FLAW75a12ZlhdZwZxdR6szHEKwVMxxfkYD/D+WG2UFGTTv2eqI
+hvbwGtvVJzP4WdAW4aEsMP46z2GzK0j/mdl39YyMYfYZ6vqUGTgIl5u6qHlNz0W
JpzbcgGYJqp6h16RIUtDyv/bugWY3v5RJkQx81E92zBBv/nmgH/hZuco91qAV6CH
HI49ULuYz4nOFJizVTHzvVoCZuRk1/F0VT/1JlVJX8X6iWzNteGVlDw5J4j1OeRw
QMRtBlG42qlCpdNffYi0Fs5gY/fzGMATNnatiH+xSh6XQPOYhirdYDxqSD/9jLDC
r+VxBDq34x9BJJZ+fac/AjNGo0Bg5qC7FJbNm0+ngjjlQOzLb1W6GXicEdBIygkh
bBhtUDGLhY6GRANTrAQPfGK9z8LepuG3fY6rp1x2L8YeJ+F8ijPUv2EmhWJkgphD
dd5j7iCWFIZUT+CK7NZJeMbpRPlSNtZCXnilqS8p9x6J+JCahf737ITyoVHPTM4S
UNTPL659/H8vGg+QE1wNOXibxtWgB12t0c8no3lMeTyGuL+cPu/taJ8EHNQk2CrP
PWxnHbuJ/PBt7TBBt5E/qxBQWjgL4aale+Bu0/HUwDb6Whx5Q0nc8PBtkqgilWcz
1N824tZyYUqagffuWI+TUKxKunzg8LZT4rEU+eNNz2gNLuDgDsJmKqDeimb2DBqs
lyjrgBqdI/wEIvp1Q2NGhlTfWUXulWZP8UM2f700B28PlzSdRr2VWwRSHthnsoI5
3X0PnnsVM6SVQqqO347YRVFDQGxxfgqjaBOtmLbBqN+52iocQvujI7OpoNmvpVMI
hu9NLdl1XkPayriL/RkF9qeWtfupjR1OA/URq8M4aKalKg1AXJ0Jraf7dlDEMJul
z2t1kMhMACQHPYGRsbnvM158q/4Mj7ohhxakHpAN4mNasPou2vc3MDklocGRTa3u
ON0TqrI4eIfTjr2cnBHWyi9of8zvGfm0w1LpGSCwBZ+yp1UcXsbaxIvQOckwW8+l
2JgqQjN4QELBWN5L/Jm1ZLEdyUrSQDvnav75vJzPyGCwqnQZolbrvOfDvMqsj9b9
vK8zJdsy6B+0d0RqR9/YpAmUoA0lF0j+il/BSkjLZNCwUH9PGrxWWXq71GRMaH2B
OFZ/W+raBiTZm993C1haSdocPlMF/0ems4NJf3U9P2rXb8la1+dA0sNmGeKe2uR2
E5nZs81l7vFin1khI8y53tgxmWCyDKxu7EFuD6wom4zCMm7M8J0MPXHfKxMVFree
mNgYZ9dpzdpoHZ+FRBVqUBQMRbCxCX3v2jeidiiEwZ6FPzY/xRK2y7fLajru7eSt
ucAKdlHIivgToKWgdREAHxjScG9SUrVChcXy5jzSF5q/U15I5RwU1NHv1HgJ8VCx
br3DrQetA/y9izyBtQJA4GS4eYf1nATyAoLaVCN4lXHMNYh3FJMdjgHv9bHRDOb7
zRLHZ8z0A4ZZZY0L7iVKjBc5gJ1tXGDh/yvOwJryVxUWdzD/LhTuMBrPDRVKbvB8
y8Qac/1QkcCEvYzArr7BoVPU6P5du6T7EBUxXqDHuV7GO49RnnGMPw9YRaiUXbkZ
nsLQRfJwyuInP2yx2hqUUGc7wfrFOsYY+GYnzSeBIDlLV0Xy0iPzQ7cJ9YiAjF3v
/oMadpM/OgR5HgHoHzZlknlShtlhPTnG6EphdpzApDY8e+pmS3NDM4wPxoqtV4+2
MHgJur21LbYjb3uMpz5Jya9FvWvRRTVmpN1ECz+f4PW282X050mWpkkbHWo3ob8t
HYYh3GlZjl3q0yIFEhHZiw6ZKT0zZUs/ckmZQSHRDf9BxqaL0ZoykC130wwp8ntM
eFJF+v1/xnZnBBY6gaw51KC6KGv4JdyptfIUSrqzSb0tX/u3nkZLXFpoBCKUZETV
TofLZHwfO/zWK7eUBBNIHWIw/VCMPRTKHZhP60M3nqb8EUcc1nvQm1K1/zqSedDI
EYIpCViP5gKexJraIc2v4obRpnZtG+hGpN2iiItofvOs0u/RyCHCKGcjMJspCbP9
jLmITrkwVKIRehcv212QcNwingqyLbFAuZzy58KOvbm4a1FS4WU9KVyB4MbbDbz/
9EcuOSmUF0BvQ3VEIrkLhksG9g8jgJUX5T5IK1RHVnPzbQTgiLkRnSHYVjzI17wn
za+Z2B9GTvHE+NvnJOxq2FrO+PMisO2/redMhT8MwemP3iZaeT21OMnIIXz8XmRG
6RP0wnNfdIfuokOEtyHoKIsizbR/lz+WmM5/whVPe0JRcutVNTSEBPXnk9EsN6Nv
OfG0A8FEYoZsIuve5zijUIlUW/39qfW5+SDOMNhzmXnQJbudAF4eGI1oV+XlkL3M
1apY3jzpFuR0kKG6rOTMe/b9iAZsckl7XdWZPzlWafhnFNLWpBC9ERsRAkYjrsAZ
e74bt1yk6IV4BoGNvVYckj2GIBbXuYzIdt148Nq48G9OwDMttuMd2XJtHiTInDa7
hnX3HBTKpvPaD8zm0oGevaQ5pmnbvEvRpyi7fi5OBe0Gaht8BZTRU7PizUB2HstQ
uPf4Vo/Bt8s2LLoSryGfzmGBmXLdD1MQx6oevFJkGGHGXKlWSCVXQ/kRxRtzJYoL
xqDOusc/ksakz+agWFJD71XpigjtwJNqOdR6reHlE4W+Mpk3oQbQxeIlGCOAVb/Z
MxM2N3YJKLX7hDTtp3umNokCg77k754ETgcIxGHt7KEXuFUn8/9IfeEjlr7QmAnL
WEyYDVyhjL19XasCVhXW8Zix2Xtycssd7BBdcMHHrUuxyJYpiYAe44DSQz/yYTT1
HJkQuJRbVrKyDnWIBWuP7VigeuZUG+EJvECDMf+9r7vrOocbEHl/YosW4sZ99Uig
I+gQs2AtuUow6POj3aS1SB4HMwMj5iH9k8Hwi0fQ/LDmS/9xs2yaO+UkTJQzUo1m
GHSkoAsoTRrktSwTdVBSGxoEQHANafg63iDDtqweR5XwD3d/DproCMCniQ64VJic
NgNARrvtQceWajByrJJJPaEoIINxi3jAgjQpghzcDQuyReBbX9bwh0X4mAgmqYgw
FBnuJ/gNv9zA+FoN+VwNNT1Dc7qRsWK8PRkGRzcfbb0kF/O9+XnKJ7+ekb2Epkzv
SnwWdQAyXi+ssYtMToM7NjGo/9/SBX0w3iym3hPxRtbAqongG2HLoWk9pNMCxxlv
IaB/u1GdMV008c6ir0B0KJFvtUAbbO9R608+lrSEQtQuBRR3DzYl41f+ThTEOxPU
KTaZasxk0Is6wP20pPVnh+3ZzU3I1wtMb06Z1ToxmkobC2nmraaDbzmb9oCg2eFq
ZhZrunxrFvQTTMBkX8IlzFBj6MlINL9J2WmW4LmS/jo3gyHzpgMCDGz3rnit4U7v
FC5XwKhB6M5l3Z3ZObJCfTasss2aHx9U5vVJxr8H/uzfw6Dgxj+0zEvqQvtc6VYm
l0ZSjJwueuUTjC3nHwmZZv4HWraoIZp3yDKMQk8gDujo9MUpUAfRunWkPC9U3Qrj
R74NKvefF/Oa137TBcYHCeTfDRnljW54MczE42Rpv4yBwdOdipfCb+FKENLUUZWr
cFvf/daciHJ9ITrswWomeUPPZygerlmEAlGw4l3zZ7oZXeSHNKfcmucVefvHJFg9
/UK0TzK9fLH5HoPhxoFpEGWgnki3nTrgWGDPKbFsU6DJrpwB2tTa1NPZHPQQwKor
qkSZfMGdR0Ybtu3hNFazV/VpugOyrihfGxwffElOZCihxjq0LuQUsThQO2j1f18g
3iQcCHk57zwipCg+3c8ZdHqabDeyu6n23aJOWBOjxuGFmI5bbsMPyP3bpb8R/QIp
1vu2wa2+ChOAb0O7HyDrGXE2wMSl38alX/dHesA+zo5hpTVl3MBimjBiiQAHAOww
tN2pjhEp2r11FHCVkKc8G4E0m9kZW/uOGTHnIfnn1DAAKF6q1DeXAu6uJL6lymno
+B9m0VnUDypzn1tS+vVWJwwxyBOMi0GkADx+2CY0WTC5vzt44LNcYDO1O2eJIIsF
jwrre6srbA/KD1Xgf6Udu/zetfFI+kCg7Trrxa6gmnsbLyIM6hYZTZ/C9tYQZbiE
2CuH9Cx4QPtB09BoAq5X/1ggY8/ThHqg43l5thao/FmJSWakMPz6hq87IE3bN1hF
dLBn7fwyYrIKTitbkP4NXyJyWoUgyQRNSe4AkGU5KItmpvmpOa3BmS7Iq7vPs1EG
qTH2sgVpfotwOROvkG/TxAeB94NUe+EWFV1dTeAqUA/FJxJLYykHf7jXsBOUZeZB
/CsRSE1KaFF2Uo1XKFkLov3vY/8NtAnyuG3Kq/MTrr5sb98pwzNY21rkEha6GEkk
oLAjqjyAFgmH3sOC8HpY9vLAjcvDC95YT4agH0wFZgWJv1fCSdhHkO1l+jYe5lh1
x2hZvWG9inW2MUH5eJc6B5xMvBZ1kkAjr1VI7bgtdZ7M/FufIf+4DTH4i3mKxMh5
7mh4Q7tH1yo60faaXUKwMw74XGAWu1DXkyItKBVT7sjoz4lBLyNfKFM3OnfWwLHu
nLP0+107zhTwmSf3yOE+Knfhyxe4l80TgANTrrDy5IkQ2cl997oCmsDMIU6fccnz
AjGp81ddJhIIt0mXLlKXxf3goqQjcm4fVNBoHWQ0OMdoFNfDvzQN7BP+gTVe9xXm
QfUZnfPIlaW2rr74Pb9kADhX1GK6yhwenFg3JlSjbZA1oJPTPX5Iyrf1O98kkzb6
15DeL1Frat8vEY1SktplaWVJ4ZmO3QAWcxYT9AgQ2FJzKQBt82sKFUK/0Brqugpw
ZoWFXa8Mkcd9Gqr8u6gZe+JJhiyeM4v9lx76Gmm7LzlHJCCXQ8OnSPuAg2SSiym7
afP/+5Cgo2RHAJmEwdyKzc6T+l7WhS1bY+8OiWoQjbt/IAMGdiasrnpMIAuJlmra
T00icJP/QT9oqZYfaznyRGLX5E8CFh7ILplZXyqbvkbXgiCRwfGFR5gUzq1gnvwe
D9wjhXrmYFz+DEX0srK4HozQEXe+P28ylajkorEpXwmyCj2WgwBV+J/A2GytXFDw
0or7CsOX2wpQhK34bC8RuaMfQBdxjVW5unhgVDGOxgz7Y4zJcOkPY4QdUQGDM/S7
Zi8GIZ6vmgj9wDmqECUHHb9z6jKvHJiAVX1yVvXPrSd/7LUy1hSJ8lF8So3/tpG6
BbKu7GjxN1ZynBSLrM1lDhPXAS/nIIetMEvRKkuWpWA79mxEgiHA6Y0Up0MzCimv
7TqIl+qjVvu27yCExcMpxQF68p11gEI8MYK0m3RXF5yiSSVi8rqY0BSAUMzBoh09
T/tT1e6C5qcta9aMQ/pkVSDbycYMqr/8QH2RDhbk4MqDnYvszIWcdISI+zTCfOq7
q3syc0RHX+xM+VVZfZDRqpeymmor08qCoJVfa1hX0yGxFpPiMl3wKna7aQRj1khD
CRXSXddPF13JAFm7+6ZuyRBCA3whik5RLaS8u2Rq6kijRuZByyOMUCX9JSQctjMV
H17M3wtDYxEwqhFs+3jgJ67P1mYxCttPteT2ay6qH93UEFaxN8K7Fv3/deKhny0e
EUCBFiZoybQznKNSvX8x5/h8GUgu+e/mGjYc5MP8uHtVry/brhWnzTUsqOt7IEa9
HH8+z9IhBj2rO7x2AjVeAgYR9oMppxvFQ5J2dggsudMe7TWYeyzkVOIfUzsHwF78
PW0i8BrfKguC7LJ0pXf1pLT63ICT41otsjRLuDHT1m5hWWmV3iLoxjuAJEYfzUxW
ogYBZ/tcETPAnXk7jDg0QIZS7gYk3e86Ny6ZxPdtwWTpqHhKEzPaGO2Ktsxza4IR
UkT3uA0LPt5Z+bTVupOXDbMqWrL8or1KujklASdyRzc8D1AvdNxeM15y+5QwP+tl
lkBLEr+9VRI4Qcz1OK+nxu+oX0FgBv256glgL/bWFek81YMIrzQFN4Nh8PGmnk3F
Sl3Dp2YnvhJ0/7aaqgekei8TyAWB3gm3dlYzNUuB9PnagXJY2AtHCvOv59ZPnfWe
Hn0h5YlvlYM1aGF4TUA5e3jza79sV0Y7q5zKRzidBrCZ7ojQJswoItr4ritSHRQr
RXIaGeZsUoK89OZJPyO5CrQyooGxjXVja6Eof60uswaGKIRgzgznR3O5AekxrPyH
2JT+jqvAgJZrA+qWBCz0eVckAbs7npflA55xTRPpiKewV40fZLmO1qLDry/2wQ3s
OOmZ9XUJqgSu/V+BkEae/EDL2Czb9Gzc/l2YxqJgb9PxRO8vUnCrk7DarFlaF9pD
d92Y0CXoayZpokU7XxUweJtPHlKf1AtsXpL3tBED6k85T4O6zfz6Qr4sKoy2Um2/
F5ZYkFbFblaszq8uWEQnMXs8s2VQwVkf3hLoSHgUEyVFae0VwwbqYhZQSniJZGi3
OV6Z+9QVOiq9vdcWP2kNvmftM28AuZVH+LCXYENKqiMwQodS5UKoPz/fVChXDuVA
TRoBCBPsYa5kyBw4j03WnNSAuHL5Oz/vX3mFyNyp0r32n+d5KY1rvCcd1A7KYXhq
EfCN6Vteacni5/u/UYDIoJ3E0lVoXAH3TZLTLoifuYYXcJNqe0+i4SN1s7IMVWv8
X8+xn1YV1w8RlnvxXytOVYnrbJUqQuJvNUEMv27j+1Hfi41FVdX8+okoZgf1RGG0
w6t2QXKBrcmepyDmD/dvR5ZpFewt+BNT+TGrHOx1lMBgFz2Y19Vrx290Mudp0zmc
rNNMbcpt0jr6/Ko9C6S/UCL20v0MFl/cpVlUdresg9N/Cyw5HTmw5Mi/44Blus7C
097N5h4kZDuvbCVNlJc/Q0pyRNS+/boK+hprFpjRcek5oLbL9xU2xy3tEWLc6mNw
fJas7Wp/GfMQoaN7IWAFOzyT5XuT0CYLZmcTh9tAuW2Z12w6X33I2W/wwOQ5ahkZ
5ELVdUGvNXqye9DRuXMB/+hTwUJbGGA5aNsuI+MxkW2/opSGjiub/x+vYb933J9y
Rr6DjWDA0TF9ODFKUA09jzsf2mKFrCW4Y3BGxD15PJvQtNm4jIkSRK5xgVYfFY9Z
youSgsO4ghocPoQsc94A/W33hhp2QuoKZ0HfoUf/0F/zvcAxWgAlLQ2JFLcRW5X0
q4FRIBjYJHNt5bGEeOOb2WTFbKjcyCnFU7wHpU45fYxfUpoEY2yDZC46aW4cqUTx
UWlof+LvS8EpgAx0+ryY/5ySEKYr95J48olV6UB25q1hosjdNij+F/ksSZK1MCmJ
Bx0NPGhBFfHe00wihfD+e9oUPZxqFpNSCQYLVcfQcOV3xqqRW3pzqK9JskxhSky7
Vs34xIpbEmhbOqClNVYL2EWXY4e855uJScG+EJ2QCIZ7++3Debufslud/itQ5U7h
5yw94WDeL9vKi29d/kuNRYW2J3kONCrYTU1rXVEVyJkexmhC+AhbCxMwPJZVBWOf
zeLy6G3pq8HJf7pf+5/CmJfwPfRebr17Norz16HBjLBIrmb41gxHgTy6ZRONLkhM
8m130bWk0FbzFl6S2gbP9JcXMVmisWRnkWDc57zUY49G5KWYEmKs418cFArSLLgB
zgy4ZisgIboFUtmYW3begwHsh98VLZ6mFOW7B6mQWc0fgANoySFrV9l3S+L+Hqjp
W4DeF8ExwL5BjMSGbgcPNWHVTlX/oys/+JvCIJ+mwplC7k+Dquxuq1yC6g9cXOQL
ROiAuurRnEFyzQg9Y1emAbw3o6gdJJ6iaNwFNbgEMVqfwV1QLrUH+nVgelkikmgi
OkEzH/efDnNFgjERt5bJd9Vfm+kod1XAhIzjm40IiP2Qnqnp+c/o68UvylA8CWhm
OKhO2uzktIvlw7DsaQJYsCHIQwBUFt4KDYI+YoErfQtTs44Fooy3VxGx3GEYsg44
NupeRcUXUuK/Z+zPpDO4We5fuoMhnWOi1ETpNWKt0WXDNSXHiHqNmIn+DXZmcvot
DtjBCQ4ibDYmQKCgcesgJ4EEWqvmBeZf24w9ZnNbROwubiGnNc5zDEDLGbH2V5DX
yqpMEP919zzMfWL5Ua/VO41nzqzJr24PzGOR/YqFXIBZcATmRsLT/v/WvFcsARwu
ulVPdQaFuxIJf57M920AEbfvcu0N5v43kyWmHlGSu+XefyO1dz/FbqF9UetMgHAj
RikPRusWudhRrznOwctagCpuWsTHa+Xypg56fj+1JeQGyMqjeKwrNohbMv5iAiAg
x36EB8CByTXbXOmBLgQE2/9ugG9v/BEt+yCsFNbh/lGZO59SXnPlkLVM6Rsjg1Dn
tt9osU1Yr026G5d3Tz4K9AxoboVcby0lbHhd7FKkqJZSSjlu5P5bBY7WZ8aWukLC
NIL5BeJCGl4fAWq2a6DwQq3XrqoqfkJF6m+QnCnViI8hgfTR/PreCFnccFqGmhxq
aIQdtUj8ob5aIoodcxTH01Q0aPewOfWHkXwUSH4/6UBDqipWtsK5f4P/g4A9U2yW
E4Qg0EyyjE9xX+xB+/F1V526Gr5qxDk8opaS8tLBXoHhwhCgaf28CF6aMXJ5Bvc5
nRhr2PDlpmlM/qY9eLtXcP71iIqIDadCGYh3yQ/FpKQvf5aTDIoW77QKMBvn+gLj
lvWJ1js6FB7zwDwd++wiXSUE0+V09hChuZ1j8tvCbeapTjEuniY4ubJHun33HVIj
MgFXjpLPzYYoEKusIz8cQDkDrUhqv/ZdI+BE1f2GHHKgnXmyIEeHtapir+ApJibF
oAwipadM/pna7ZA9zZcnKrAxoWsqAD/1sPExWBkqrO2JT+IGkx5TzDhFr4xYTuJW
exl3LenED98uFWi4mMWi3DJO11v53argSBUMueO6bNY3uBrKANGWZw/YtpvYXqLC
RGM1wk+yf+tY/LtYW/Eilyr22mRG+GRmJWaWeF7YRCTfQqVo0YRS2vZYGDYvhFL9
yUyOkdU3KoYfwKnlzi8xCVyzSfJaBLzGWopRCK4VTS72Du4EtYMxkcQ8A61UPI8e
oDYuI3LlS7aXaMenFKTAJTt0Mp5Eq/h08ESbn8U7ch7oAUqnug4B4EH28H1P2VAg
uHh5pGhqWV8OTARmBCat0Kc7NXDKeqUcWbk7x67eZc5mY+igyMKlisTl4r9CLmrK
Lv28S9HT5lXagoRgNOE+fAwvIJks3d196MxK7Vc0t8oY59rP9XgnmnqvMzdXP/0D
9cHAgiPOSqUg6BmlMzQYF2AdZHgzA2eR3pIVT90uFLlgKi7/aqGT8WYm4tGMSLsE
Imh/nBdYP+LrS49SjtpLELAimqTlMdZ66/8Z+FJBJNir/hbhjZK6OI2Kf4AHWWM+
iV9RHYKetEcppk+xZ4PpuNI0DY8LyXQlpCsXB/Pnb3stK05wl9whZcxhKRfvaCr5
R+Z5zJKU+VHv9prSd8sQ9I7pudwG6ZJ2q8+Zjy+EhFEeRED2Fai7BnCVsxpxSP/e
72On8ziaTLw7MqMk1d39/sIxUGZUzg/s8vU1jWa4975Dp8UsWrnuuB2S9wwmpQvG
aXNK2c5ahoD/gxPlMQ/gRk/egCUGEKYdTh8jTV4hKhnFvYkCzwB7/3uKR6ZfTVai
Yjd92Ji1rSvtQ31WxYhlRSBFYL8J/+MsffF099wH4gccyoMY8+Aa8jQCV2XTDcho
uBM2YvhfpqnebhvPMbVIaUZU5Zp1JBdbG9hRHMmbzHoJ6CHE7Xyp8IpVIsGgyy67
m5WiMy2r5SIjolUJN4+mvtZXsfyjBIl+rHWMhmzAJlttWNr/M6uzWZKNyrQGUPQ1
4N1ud9a4K41ZaW5KjyWhhRfNp/H8U7B8W54L57ndz6ENG+HK+AWixOG/IF7B16Fl
05yTE45UC6tTJctM8Wjq07YwXCHqtCrQeiJwv+aEPvGMkP9fWakuHbhNcJGMZUlV
f5r0hrr3BgRyeUQX5E5mti/MSW1ZTv2EbiEFbTZ4bqnT44VviVNBQp3TdyQah9r4
MnXTo196d96tg/9RPystPRCO3v+vXDytfkRwVLoBGmtyBhLsTaqj5hFQ36I9mbpG
phwVJprqLPLZjVrlgJYtBnUmLzwg/rfYtxKL0hx4B91qzcuT7mgf0tX300zi5yU/
cZ6QamtjlVBgxGTecIVXYmyHijWqipAshXBtbjzoxz0x5l45GIltp5aWy5TcZJTw
/ZEfbhMU2t8kAeOpat7AOSZVhDXq2sA2/7I36bhCJV2XJRaC4yr3SXDI3nlwKTCs
Ldh4+IKVGhbzJ7qmWRnfEO6fUJclNauGXa7AyF+l3aWR8TigMbFUIAbhhAgjREzQ
gXz/hkFm1XMJArQQ14UzZ7Cf7jf8wtLhXAAP0Lv5zb0nV8R5tKS5q7GXhh243SjD
fvCSLw7LpB+jzaoEWF5cOYy7MdiABPIJAZsJ4dOn42LYRM1abaZ4kgpGP6ppzILT
mulM0h5wvXCVMQOPdv8kwKRcvzA0tjkyUhT6ogsIlX03vWpeJ+YaA+OtbnLOq/4d
q/EBQKXpC8cyayZBN9CCM+ZXbv3c7gZhPk/9BQhMLKDNqOPMUAl+Y0+mU8ndZ5Ei
jeJQENc59EBfUtlCxrjT/XTzESey2tofehuqkaOdc1qljZPud9F81bGl1dAr5shF
DUoad6HWdi0wN4uCfgnaiLQ7QZ80fD+pN0ArtyJTM5QkHiq4uaSzrVYGHPL/B/9N
ER0nagFPT/NwofhMewGJ/w5Aiki6a2xia3Q7PpKNjMYxRYlN03McmAzl5fzmOW16
MpTNEzHJiWoDuGOnyGL4PiXO/Dci8hd2p9qSpCZk8B6Y9kaF7R8s1AFRvCBhIeq/
lEb8xJYPz/9ZnFbufkjeuejuXuG7e8clJK+Ew30Lkfb11Ss3uz8eKIXs1vIG/CIg
OB+ZQ9Uv1ArHfyYncgecIsFA40ccpVhcTmmx2KFldnq96OLeMxZc4YcRFOLjm3mW
zLB0Suk00AtVtUwOUO6zDasC9mWerxrXDEKcx8APT6uNFbw01SknhQdZCiyMDKRM
pxk7sKK95aAhqCkzCdCMkH9xL8qb3wNjPpkWJMQlaC2ouUQogdICmDOl3fBnI/pB
j2GFKOGrQW0RJLOy0b/hlKfmJYyrswYbeMv36AhxP2IdvCbDZdfUtX+/bx4qR89C
wU6yr5vPHlAUcRolBLLGClPeZIu/nsiarWu4hOBc1zfhG7r4c7Lpeaydt8HqTnY7
uQpqo/LyLrqYC7PAuKW5JHCZbxJnFyesDlRXSwXMKlzFr99PCFYn0LLDhJ+fbDvh
o6sY+M/u9OO8KyYRogHzYjuVTSto+C63W1AG2oVzvNMgGwwBW34ecbZinibD7MXB
1hCuXv3aBNF6nDLjIACjBnUFW74m+A1Y3dTL0IWJzb7gXtFu5TrvVD89EgHbR5gn
pAMnqG0i3hi/ipOgmpDGB7BNelVlxpv9mIFiqQzLXaGH5btDxJTpR39KMiDeqCT2
N3p6sgeXztKtJ4Skpgr7n867v5Ckn/dHTL3bJFnRrTQZnIZ8qTxqeXvGggjPd8LV
5Vwj917g75tIFBUsMm9oZoOGeNMtWlAvzBZcZERuc9DlH5DE0goV7yukZbp/Cq9K
UHagtZmVYhB3ajtUBCGViKXRBXX6yH8tuJkmtZxz6tadO/IFGlIHYByvKe2KlWox
rBgBqcgPHyz4jWCoZqcl4P/iwiqOm61IwSxKwM1FI4sjHQPvWaQEOPvNzD124mN7
c/ZYqFV3DzorILn5031/EuZFd3uZ4BFID4OT0Q38HSbWWfjix14nVpd410fICTqa
Sf6bLVKA/UFeRu/lPE1WzYylf6B3PTfKmvyLA0MEwLj0Cee0UqtJgaE6PvGNOsvv
ROFHhuXIdqT4sjgj+XQwwLrmg0ZTU7rZMk3Swxq2MJHb8AQZC7GsHWMGGgrhhr+B
OaXZjgSfeQXUqY6H9o5F98oOjgvVazzNMVxWtoKeh4doOvRVOky9KO7NnoTtHx/U
IKiojSpJk5bLcB53ob/+ufxOsg1VUsD6llohoBzlghhOl2kPMn79fHMVGLyd3BGl
AD79OvsqTkVLraKOyWfM4E2DPHG9omVdkwUx58p82CZsENvv6wmIATLOLkQ+1Qx8
JqpGbWS7Cn57xM+NjU/rc4bhAHFVdBkodMGdHeRszSliNkO3zwRU9FEf3J42rJS1
YELNBO113eK7vgdgyXwzQoFm+f6QDhJWharl7VULbIA3mWnGekjGlodQvttM11Zx
jDQIPNj1PvNUouzmavr8+NdUVM+a41U5BgBrTRfZse6fK9Mg7RrB3mQKvdTHcFDJ
tnWa5SpObxLlfZvNU9Au1dW7qVeSG1sRD+l/9JquK4x/1MQLITxh5bvWFS5/YA/W
h42aFM0SlBHbhlg1RD53ZivGI/fVHldHcCMBnWGaBBd14eCMYVgQpAE5LdlXrGGo
97nmC6WvqdLUNPc0NP698Llba3LEIkDL2ejTihHLJdXZEnL63gdaO/l5E3OBCxoJ
NZALTWKslwfZJOzJuE6wD4QrM/dKdvxR64U3v+MNVvLpMjb+pV2eeC7iROG7pe0e
dIicZ10yl7+dZpTx9hUolsXdnG16+4tktp8kqSTJmThYbfPeNtuDtjZbWBZmjovv
2zttUUWLhAUEwgzLFiJsDsZv/0xA4C5CcEXMNuyrgQ7htv7jm8DmJsm7XZHQM4MJ
pEGDlTT10LnZjLN5x6+5pIqFab4qmvBIhCCszROIeFEIHmLDddFIIAYCGmNPubCN
tgCTceZmC8ppeB5Inj+mYPhSGTYwnDR/v753mFRdpNexAZAppnzFasJYyjBq748x
TpxloRpFPTy1WAsHlWdt5i/E7LAWFqWDz6zqlbXpLmtZHFD2rdxcCW56dKPQquVL
EBBZzS+9DeQFrOsuE7oTgK4Ht+4LR9NbidotoNtbXaD6Q/kYCIF1HSiAeOFEoeF+
AZr1T08qzGwLFnV2yJeFISBreX5MxNd//nNWzXQN+xeOQfurA43HiMQPkXtV/5/G
gWV3Q+v9CF+mcpSBLv8lCVASnNv044bgKIdCLeoN+iLjeCI1WF5vmAdhuRSz5vNL
oj2L9RfjAKygc0LnBkVMGKf6lZVy9i8dgKwzRozoti1NkT7PGyctDpex3M7OKkeE
2ZXlPq4cqn4+asxmWq7w7GVZSueZYV6bwI0d99p+PFX5w2nmn++w7Pd5Be7S4Ezh
U0407JPRfw4kMrjSTkRNQcEQKBTsapmT1cLvj5i1SL2iDTakOtZUVJ4PH5NHDudp
5P1lzxQu+DsNesSpx1SsXYEKQBdJbCqmt6u1bYtE8LklHGtLf6IoN6Jp3P2+dMP9
8gphrEIA6T+EnuQdgFZP6jqe3G1x8bh3RxTphqycmnLggmqzurACr/KTC0Jozl2J
8JlH8L7pwX4Lbk/hFz/RrvL30rl5OSc+cAZVjdAVbXixOK/Otd0zCl2TqCzmdUQs
Cum3Pa4Z5cmgftv9SG03LsWTOx5gZvvBQ/XXALomSaI8P4l7lWa9nGt/h61h9lG/
uuPhsesWOF8Hb+l5g4rNhyDD0aiXAZtu//D/eZmNF5PqNSG/anDapABilSOyZ6Sj
Uc/4QnL/z0TLBSJMO8IYDuHI7G3yKvlYAspx8LeomaACF+JQ/GESuw1IPhaP1sCt
aW05hEBSCNpnneiQeO+ZRYag03c41VgicCZhztkLO1DAW6G3OkJH+GwSrKWcR4xz
JUa1g2t7hNN80doCTZFY2J5PJT7cmxtug2HfT05zmfWCI7atBPiEv8CH5lWd1Mrc
lKopqIAZGqS3OgvCpFCIk3KRHkFQip0h+9C3uC43YrsC8BpJNvD3hKaQs4KQ4xfW
uh0h573cO1OCWE5QEJY4q5PKO2XN0Y8UX2bFs4dSTsBidE42uxieLMGcbPcE4X1T
9ePkHEiM+Or5dxrM0oaeORnogm/7qBrwGDPHhMRCTt0P8W8Vua4wpULsdycQH8b8
fKjyK4y8hd1TAJaUCNZMdURBwVPZkfdRqThmwFyTOabWoeV9x0ORXmYxbXbPYxDa
kglwCPgsnEx8ZQEaYe68uc6WP+nY1UoAO8srmjmzKYhFu7wmKSW4bBPT1RQWRBhR
jYVw2uGf/LhLN+RLH7klxMC9V0jjdyqPBy6WrLwxVOnbdv2YnGz05BcYfsDC3jMc
YeYmbdSuOtoJl14hGhGWY2EZ1aa1Cv+KbsKI9cc3qh3kN3EeIxCt58Hgdq4OCYVJ
RqYPWXHPAItmxFHPjstEAXfPfYaHT6OqY3ztMBskdYRIVihulb2cXjnv2mVTW1Y/
oICLLTdTvcto56L/Kn9AYpyzNsAwBAH+6FICq+NLV/3IPz1N7naI/DRbenakTDsr
+Fxm3UBDEqO4QmM6qg9s1W7ICHyV9gqWdaK77Z3PjcRn0hn3UdUBfMDBaBgPCRAg
VJ8nWvSjWPG02ihp3EaBhRuEnwawW9qitLLRVbd3oUxk+OemWIJNmwNYHt9UwFDr
xNfY8WTfgRu29hECm2MuPLAP5XGrQkhDitIHoLFOtSTsxigzhpTAYvyDyswxCSk8
wfCjoyzhvt1y9uztGV8ETVY5NrddTIZunRe/HU0q43xnidC8ks0HrCme2nMhBHg3
0Mnl2wyfaeMxRd8282mbdBuVWJyixWWdOPD+dYqp0ZuvCeoyBVYJxITn8GEXyMF8
GJVlB79Gp7u8aTDsN71s1f1CQYa9syVcZsKxhkdAmChV/i1257rXdbqQhZ4nj3wO
Z0swzSy7zqgIeXUKfEfKqW2u/QLVzS+hHopYoUSQuAYDYcmvhrMEcbK/Oxiwj/0V
5ziQAFFUmH83EOZqD9SBJ1y80s/pqA1k5sQWqtfkaAucckEnJ0/NO71GIQ5PRHbF
w/u8jPHk0SOMFLLVlc8yJ9CpcHQhCdldKB/tsaBOukeQ/Xuxh31+ddBdTEqKQgn5
xl5/KFPW8DjsjB72cus3FyElzttmJhyJ+85SMUSGvvvD7ynpybq8G3oN59dnoSdl
dr4+dudUPrdH1xahN7AS6NLI0O453SFHa3/m08onyl6ezCxn8m9DXGIynBJnOSNc
uyPTbtPIwfJUvlq0ZxBGwFV/Ncb798jE+iNCVoeDrnC8tMCMbJw14fvPP563PJiw
kBn6BRrzTFdrPuiOWpie03+dQP8hhDrEO6zFrumN4OzbRG+cbf2qbq2G/H/19dPM
JfPfMO6yK7f7c2LgaY5PSiIWA3fASOc89Ru/KpqOnmCz+KlNN0AzY9Pu+Pr+8DIP
wrAV8p/jnZzxhb/uoBGzWM1EhsRFrjNNxNetsGSSR53gK1xyAIuwxo3PoU+dZO1k
V/YtmKHqmfI/m0tngt6jpwbgr9WjjMmdpRFfEbepEyf5++L9XIHLukYlt05oVMLP
wHtowSRexMJohzhq6AG7n/bPXrzJ80A8BhotRsPGOdk4FJuLVt4jTWvnMiLqayu3
eaaM40aAnyLl9K8uRZma86N2AiiZz4cF8mbN1CEu1c6oreOwEswSFO+CAum2KisB
cGbXKn7fu+BOaKj+ZxZbifP/tZs7mRxDypesq7J52MpwBp4LpEBzU+lqo8ki3N/y
mxCziqhrl6hKAe27DgaGzFhcKw/8aHHKzTDg6F0Gg4ihDr05uYoeHIZwjqyB27UJ
jCvrocgf74kEMz8b75QJTJUAB0EKAQQy5t8B9fK7oO4y1NFw030vPZnmQ6pgFSd2
r/PYrYZZX4CG1KHUDl0KZpuCLI/rA10qte5ZmeWNntUPa7pe04DpqhEhW7mkoXYD
WnXJ7xBgm4kp4guAeUEY08gnWZUHsvVzol+0z2ivrgiDCezDQRd1Knei2Q0QRTAH
f7f5/wbg2aRHnfWqOj81sTlKCnO2Ub8Ss5lQJ7ESFhfurl0FryJxJK2Eod9oL2u2
dTkw36OsSBd4Yw4OFW1aXJrPhfM5MWpkS/O/ncOugmL3YUe0hBwB7mzyaembMQ1+
lUpXMOd4NUUh524O2qLS5d3vYyWPaRcYzupUCh1X5rOUsdA+cT92ZXZyX/AVKl5j
XVQAMSNtrymaIAaTjx43aPmQmDKjZ6wK5t7EP/YnC9cf6nkXFUJSK6TkBy7xSRln
KxXwACbhf2qI1KlLhisaNacoh26Moo2iKSKMIWysMx1Zl2GJAPn4hhfXIDeSSUTS
4L/2Ieb6pjLaH7r+2/PSXoeELIknLobtK0TepXmtVYIyVGLL63TGwWQBh4Abmc21
oJffeP2IpPpCHr1DxgJZsIpW5pAHJSpBTStW8OEPXpVJwz/H5K2GGX52AbdnDNW6
lTqKiVtdriZtCh3MuDg12CblOIg9PTvbAlQYggZkQ3kij626XcnW5jF65u5ps8am
xwQjX5LmGmrJtUL5RCt4+BkyIgdjiVVKPg8cOfbNQOi/thvWt9xSvKWM4CyDsC0y
3oMxqDQhpcbU2Bd+35RL0veet70eUDdlttpl4imTpR13tXaUYRYWfwC/qFPrnrRC
WVJ0XMOthfzn/ci5zg7Zn88fFfrxJQVkFRgEosd7NyIlYuyi+XdSQftQzKZ5isd8
47f7nR9KCAy0wQIaO+ERVKUgK8UO+a9076/4KmJELtTmhOPVxhCjwvwzwoZKlB5T
PW+UBWHMJrYXM2IKjEWNlRERIvagrnbXZjoiVfbcUr5IyOn+q7TVicKBF6cvPZNF
5hzRQiJas05XJhV6zr5Ox0n9vPnj612Yoa1oKL+iQLXbbYINl0ij1WG5g0JMlNNb
OBa1hnfL94FJy4/DEkx33ZdovUcFNsp1SbWRjpJLZnT96X4E9bE9fk5SDo6Q0TS/
HG8yL+54oNuH/tsmffheFvgJ/e07BfhlkpljTocpVCtyVsaFnpRb6gyXCpz201Tj
enjIVQ8qo1sP1u0+27oERlQpyKRt+bpHCnuVDNd+QMRnPcCwqFVCEkaZMV7R2Btv
p0GEFEGAZdmBJ3nNpPPHVr5AV+mzjmiHdSweIQ+JrXXvvvcMIJjVmvXgRRQtLcCi
ep0SKMcURFyAylCAJuzX+xQhxugg/WMlf2WUoXRYIXLC+GsqKZKjWfJFTCd/cQhi
4N5lqmF7Emcd4KgynxW1fjRcgTtVk3LLqmM4WB0SMmlBNpwST/t10IMfhSL+Drvi
Q3OZN4hRk55IyOb9mPnAJvTtrzFvQltkrXsWnBZ/wjYmlQNVX7hheO0Uw2xXqd3t
mz43u0VnprUA/8axRgkDqhoGQJVAQUde7bIchkyW+u5iQhl0W+WbasCiEys4R45J
RgYjAzzj2k03uotEj6HGGCqTEda1ZqyCRpFrwrhaEX86Uk4lY4vhLseYcfwP1eKZ
NVbb8EF6i6qxsbww+mxC7Q+2iMjSjDuHUx0v0EXUTdhfT5x+H6r5Xc1StZ9qR4gD
PdZNZMKtOtAFafEeCZ2aS+ND9gpffXoL1SuDkHQ/Pq/sCt5qO84OmgebM+2wEoRF
uXHBJA0lVLrW2a73EIt08dWhZULUD4HK68FVbcuUOPvPR/9ycBq6udufVcR0I1jN
eDbATACCni5zoJVtlIKgwLgXU+ajr8LSM79ocLFUe2q16XqMAGZiuNw1gEjnv0mb
Z4VJy6UqenrnTlVDq1YlldrZ/iagFH+tk8DdP/opc8YkHDadSjbPynz0+xWZZj/6
zeAgKllCs/xP2YfmBZmIqPj1ZlD8//7y84kCjLKvvNbh7k0Y3fSAzVvqSQcx0UIr
AKaYS+IBkIAfHMhenaEkauY5ljBpCu4VLDdV2Z7PG1Wqi0XPFAZttWdHxPhEyEbz
Zl0AMQEvnH6Ay8chpsbDnacZvzx2jrixDhb7mYDSZUtJBUsfX+avkSQX484EhVU9
YGu9usU3SGI8dFuEwmVgtBblZ1ewawiBC/fckgNFedjD+qy1/3z8+zCxEOM7DP/M
Z4820SfUann+RaMf44jsL1fzLTya7m5kLKVKVpG4y8wYAWXecHXXQO+WH0XpS6T6
jVFd0uVCCYDfb3m11VvMSKUYzTqZmQboMlVxgWt1V3CwdtFhpzDlfsopCklIv2NA
o2zSF/dKucVFhIy478KKUoN1RXd/7iUlHXl76ddtuILt0NSz46V65FkTxxdk7Cg5
EIx5SprRUpBW1+9dkbkUQVnfVZyusd+LccQ4c9mjb1ymfkI42vXg2BFOmWPjkg5a
tD7Q1XJcbke+F1JjMc1Sqy2lDCFFlG0RuFMTWMJdG1DXhsa5nLTrHsWLQKJW7URa
UYA1DMdEpfC9FLMwoRlkSUFZsUEHo8lnphCGih8LG9AILMkbQY6qKjjixcY8KxrY
Y7j0JEq93wQGvKcZePqqRC/93PrFAIKFXHv7ZFBkoqTCqc/9D2nltiOXtxif5hPX
UDZC/VqiLnGT8je8AXPOG4mVIk3qURM016Uw7ROAHwO2Z5RcY7EnvtcSclRl2Nx1
c6FDWQiELxzO2rqoBStZ/MpugROhJKcTlbuckHoi0DBpsVNIblnVyZyV0YbXVFjj
TjqPHOZOVwfe2UnjsiDFVsqUIhkRjF96IW7/RruNOVm/8a9psPToOeU2SNxs332I
eZhhR22o0syQxXmFCJ7kOYG81AZD28Y/8hbc0V5Umr0I8N/RvXNmxDjG4uad58IQ
eJO7a7J2zPdYuRiN7aYIdU6MkVaGblfKFxaSvzi9Z2Zjujq2sMvnd9k+/YoQqSpI
ubTzI2tLGrQOVq3Cmd4BnILYA8AMjnHME/tEZ3wup2fEksfrZ68z2TosMKMO77lp
OqY9FvthduJ63CAiMq2izNNqve0UXiPAHbhLBDOpUnXteD5ytDF9lU7IH0vjfw8T
ZSIMYxr/aepDjbaff35A9GKHgmh1Ji5P3IOUEcvybmtnxZxkqXJsmnyKlmZLjn8T
v7z/0+jjWTwrtPDfMDi0jZoRw9CCpOuR5Q3B3KM4O7OehZWqSnf7kQi9JwxLCf1T
SX1q6bc/iJ7Eq2GlNH+i79+pLuKlNU3E0M8noC9XM4WnKC1BT+5GWbT/Cc7gk3NA
jn5JJrZND1Vg8KJatA7BoqcUYzCpu2n5IxKvzQp0wCZ5yr8fxw91l+GIiauBAE9D
sJ9qYIsN87KtJ+0pDVhfZPq9RAn6kIwO/Oq5m1RuzFdmSHpgQCM73HUpWp5FmpAI
EikJai9NaEab24dUj7C+W7uSYM1G/40PfzamKdWxdWVhgSGwEP4GRXWBIFrwhYd7
aAsx/Zif/m6VJKaJEgYioFL0CYeo3ftE7U0tZW9pY2Y6O0QEH7dk41ZpZV7/jiwg
LXQO72zsNeAWFirDX2KyMiLX9cTu2ALNkEBXoQrsiLv15SY1LF2ZwYFK6LNDkMRU
0q8ft/4nDtI6ljPd0XzwBBDhnKFP25lWDd+5SEyyv562bRoo3lriQdAWMOyFddiU
340YhNloNSRTMEadHY+9IZMrLfGaG2v+sx8uc+jmK0mEwlNDww71ULaJV6ENt0ot
LcBfmC+gUzPZ4v1NsCOcVpA7J98ZWWJBj3uoE5leZFVhQTpk03s4VTJRy+NZ1ike
cfRR7Zupihng7URIdOnO0FKoL2LRpeJ/+edSmsvbqc4HppxFpkqhxH54FNVuoTma
ZNHPYoeDGOvEQly/0jT7dLYTzSgv/GVPWqdw+W85xelcaDpMeEcLH6w9s7S1kzt4
18nlZ6KcrKvIt+JIbKcDg6tEwu0FS4RrfnbxvSr7ei9iI/1g7zxX7zrj10GQkbaV
e3I9g900yM26dwabDtQlmfXR0dd96s0NpU1b6b3p/qnoQQSH/b5IZHArj/E3CD/c
MXjewtJIdopcgp3/KYOmoWJeb14Ccy7MbCF9g16++DSZ5ALKEyR30UqjmvmLT6XA
S5uo0pE/Jel8Aq898cA6qUbO9fNrPtqQE4LiBIUA9MEAlq7Zvu+TT400dN1V8kRQ
2qvTmx73QyttYWc9PVM5h7BCcthAY7YsvclyzbVojifpOhP8rZcp8kp6TG9RDNbQ
loyW2Rj21FOdQiUyVLZeoewirEmp0w5oVTLcXUD8HFF2heWT8gro+ptVH6rQGouL
1Lmry0twxtTd/zIQvTX1zJIJ3sXm+Tz0+drKcxIQtiJLd6ELRgAtiHjgFiL87Dul
F1Cu0l7JRojvbxlm62iKrnxMG9wueKf4LB3cK/2/nSlFnBzo87dX0gJwBmTHNjHH
N5mc++pS2GP74gCbbwZybzMQ7SCsxFkzvzdITzwSGp7T+no5uOvs9ECTHZHb83B5
MPN7Lvt/pj8nCnZ4ellwAGrRd6fRZN6Uo22Zp2ITWVbrMiGSfIU4NN/K6kGpslIv
bPrFIz3TwX2tbRydBeqEJSgXQgtNhtxjyOipNSYB7zh/W/iV1ByHrERtsL9HUQ93
6s+UdGCr5shwSboEpROVg8WR6BsHNlQfOof6aosRJ5idpnUwvXKoKpbHEgsnbLBN
sshnJzeOaCKL+4jyoXdhieAcyFBFaIrd6oVh71/ywqMw1FfgeNF35iXuTNh0ZjFS
60LnLuvayzZGteAKz+mSuchzG9fth+S9AhcgvXS87+H8rlMSgGHoSrMH2qzRu131
5NNIWY8GpdcIihf6M5ScTWRbQgrFMif7RE1n/Y9/xH4dJE0giXgXC/GosD7rbIte
oVu94RtLqXFFbeLRiukZeIGYxJByI/St7yBqFGqVvtzAq0xHo75LDEgo2ydRwLTp
3k41PuI9EoXOFr9p6Bp/2xwS8Te4Lrn24t7M5tSKLwvITcfYGW2HwN8gxZudPD8o
hK4uf4DMN+xgc1mt5wyyDM/GOKHEAhOSaJYvaSrdKeVRDQoqUQPU1qHMbGuZxJhe
2cu9FU8BBy1n/YXmAJNuOOYg1SKWGfyw3A6MOx6vDjcydSN0hJJERG9x44h+I1FD
+WZ/QtE1Mwug48EeaXDLosdk8fupiyfKscaXRc0UvlqGQVinlOIo5rncmTdJ7Wp1
u2FrMuDjKpvLstL9714aksqDngv9vr9I1nK9wBcDpUwc8PoHofuWSuiVIX9wTqbH
4pT3ImsX7VgFztpJF4clMJ4amxSEAPXbCMDMr4z45om2TPeTUvHHTXFVUWXmLb/v
JEsUJ7HsZ2Eaom8ptFkbv/kCE82ieGlHAgXyUcyJZrNJd9VKX3hHyUQsEmQXuna7
mfhmde3voDXKzOzAbYQH3jNetb4YZNgQhWmTuR4c/21ooPwzsbQ57ozddo3tol3c
BssPPZLUokCCQb7K3Gzt4e3UgGHAPFitMk78Zfop/lHmQ6jFztNLpjPdh+Qepbvu
GeT82zpdcrMdW+PGYcHYLZl8X1sP7C557VJaSOelgT1lNQr9/QNLfjSyiiGvZAGI
DKo+/aZ3XKesrZZoQRkp40w5kFXJS4MICmxVDcTZGRtYlAbd2PHM4682hfNVDD3V
SkRJq1mEGLCh9JEuqc9H+pX+oK9IdBhKuZotVaIOVJ0Cu5k7aAT+A9gruRh4u53u
b1pb0jG1jM6rREXXhZHpz0jkwrSMEy/Eq9oTv6FBNYDW8UvsPnlbgqLrXnZukinD
QOOq034l+Svi7Qg82imikmz05ujPMp1XJQ2yl19nHNoDgtergmjiK6KAJS+6I/Sv
+dzCrfnw9BbKjJX2KqZ/WsrcOjuxWT6rzJ9Z6G3WFhcomPMtum1T1O+gSXFJwude
n51i5EFSR5W4Nlp4iA4SUxUVWHLdVySq7Ofzo0sK93Qq8kdndAqL74g6zvVgFsy8
0Lu9bU4yDa7NzBqE4M3UEv0EoBOJX0xKxBJBQ0CnVRu8VOM4rQunNxJWqOBe7b5D
4HxvsZk6vMPTjNzpvdn4kvsZaooAvNf5i8BCodiAg8ki7hUogB3N64k6VVXsrRjB
7vGAYiCMKz/ty6xiJcJABXMiA/qHrYvmdvm6u8WWw8h7kuN7QafZFC68z7MTGXNC
aa9nozBXhYlIKpwVgbuxijQ19hUodXOedYKyVtcbDi8eRNug4qc6oI4W31FJEv4p
etIGLxtQl3pNHt00fPo4rLcUUsCXlMGzYKkWCMV2twbrXQChmpUcrgFwS+VM1YF4
zzRdbdaU1w2UvbLzFnpoipYocrGJR64W3v544wZP97YU9uVWmSx5vVHN/MbgyYoe
uA1Tzq8ZymrHD8+rwcWvA1wwe5kM1A6RqMfE2Lzzo4UWX0VesOjPrjWv5zXtOess
I/sJg639a5ktYFM4zY2GNk/uW9UCeZkGaMkW5+eE4llZWuXs0iSR1RnUr1q5L8gl
GkvWXMxZL0ZdWUTXqFTgdITebZYjPhg8mjy74qAYe5PAN7seMkENpqm6J7FQYR5D
26327aeLiGQGYPnFMdcnZxYT2PlC5xu2b6wR8iJvWfAe/v2B9inxWEp37TFk2uQL
QZuQL+vWx3dMhRarEr7uSKoABY5pKdUTnbzn+qSHiIraF9b86Xr+TmXaJYI089G6
3WSX+i/OC5eqvdkqcYdl98JOcbkqPmRDZobj9sudCMBANUu1nQmsHcSSICp2S3zG
VWbptWvWVJBcl+OGRyMcrHhY9pPWRIMLctQAoa1oWGSHMRGfoRwjbrbsI4bHPLPB
WFN+eWNyDNTWfJxK2V++o2MRR+dCXqNWiFh0ewIoS1zONPT3PNrWaBHQIw10pvnf
jX4fKurb1UPJU3P8Qvyy0jYzJWNVnSB+WlI+55a58jgcu6Fps4+4m7/ffL8LD1+T
lOZslt21QEoLXX54+tDOzsS3/FbXXKBUUdk0g7fV6e2YcxuNQHHUBFIH+XfCh2kS
/Aoi3tYB+VNX+3jlxPWLf/Jbja8rnWrGtacunk0w637YDI7HhgMvtw5354PTSubZ
Ohrhmi19b2owtp//Ec2/WpVWaf8e4B8afKLZsAt8tPa/4sohMfHjp4k+byra8pKn
T3qKAZOSpuqKc9L/4TqT7zeV3XSlcJ080u99x+1qppp1NHgbe6HRgOzdhY9jNcrw
U09k3TuqvbfbIuWXUlvuQ1G+PifCNkZaijrHL02GkhA7zrzmq3HPqtaHdnoYmyWe
dXhpQ8k/i9jYA6EluymdZ/mxb/MMSwqoL8hCQw10PPLwJ71fuw/4KV0jfp9Sc5rZ
7xhWsfj31oj3e2L4Z4jn5qmRTGUMeJwRwAapFKCZRkihZaj8AKuS7rb3gh18dL/C
mbQry/8dP1nIyWSXJXUc8ozw5+ynPvfBmCO7KRGzrtKlnJO0611llz0/TQXEkNEY
f7PiWLgkc/AO50Ne9E3RdYc0MxP+EApUhngBCCqKzkDuiOd036dWbFgmsFFl450Q
rznwYhDv72PYtBSwS+yZI3EQkBzv37DxIpHjNXLJSK7zO+wz5IKtC9undfxgu+Pb
xDO03JSjYay0o05TwhaXrC/6xtF1PuYobGxZjm3JQxiZn5kqJfe+tBe+DTU7k7BF
X1TDDL/MgsYQ3Ox0tq6MVRbLV20t7Z3RKhiOclpTCB+wRzPpMzu00EmiJ7Wz+0wa
hIxBoe8NamVjMKZVpMvNiszE1EnNVRMpCt8+lcQrpI4UhPnhrqEluH9m7XF8nFVI
PVCvtNsvvhNa2zYuCg+zUo/wyiHAEnWXHqHdF2VkQNJK+HulT0ma82iKGhlLS2Ky
4qx/Yskn+Ke/Zcf489B7d/2yS+hi+rHBQ+7yKRVNo+NvgjLefgVEFf+eh0mYe6ox
YYxQu4MO4+94xQDpIMoxYOJ176HfP/o4QGCcxSoHnW0ZroA8wpR0u0P/d/yHT3Vg
4Y7X43s9mByJyMUCanm31Uswgvm9sEv99pmIGEPQyw5db2XllH1gtNmm0DPH/1N8
/tkGb6stzmTowqYPJnSY5wleo8yfNCyX6LW5QnkYC8vbvU46M6ToAlZcCTdoR+Fn
5rG9mt5pPBM1tqI9MXV2cJ3qXL0lYOlTf6Hmbq3IpkcjbemXrXFAJIW91hrRZz0n
vAhQ21I4hsNDHwcIE+w34+NyxjQt4hGZORAUi8jTeFzooLhbkw6/f3LT80ceSL9d
4qmZsmwhzi6uDC6uLuMKHKrJpPptC6JFi5QSjHuRHOtmr/bGiW4h5lktDVvyI2pa
dKkgNwofoO76BSS1rEsBHBGGXYFlFD0uQDekDxEltTmo5D3Sg0e385w3RAAUL0IZ
TY+dK8vzmJloWGiBSrk9+P05Mmql2OrxhhMa+g1Ypvle0/gO+IPWeg31Fl870q5u
DTIrOQgGjwEg4gI3AMQSW92dc/aLAL2Vz2naVemPKRtC/inNSnVFYE0ETfhPaFC7
JHjWHC7TOzZ5+/j9apxPYUTOE+rJuTSrHdfshmnGfBmee78yneDzOvngbqjUEsnf
7dsP9R0xCN0X+HSfXAoiJ0wBPrzq9Jdn2q0H8j1a+M7VE3O9ELAUyVr+gU/GFcsB
VQDthJN0CyQ+/y52up7Pn5VOKLzrfTSQb7ySUK1XoL7GKLc71B9Atp7cZcxu9uKy
F9XqUBhFWK9Y9dOmuZ4hZT2OiM67ALIdOrrbL2cRLT9WNqoUPtGez6IxihMy7DJ2
dN4lZWZQFGQ0Uc68egn/+Kgv0nK+tVm01bOMA8Bntrz8/XcEiTbkSUnAVPMiqx4Q
VLJE3KTEJDxTTRI2hfN9vFl9FoQq/QcrLM01awcO1rZz8Hwf3C4HjIDzfhzgVdv4
cZxQmfl1jMZbbeMhwqzjWy5K4KbLBRILhN56Xe1iJ/B39wEFXfud0/IZ54HRb4TV
fvbc6+aihWnQGfuJKQ/dYUwcWjc+nT8zxjED/+3ZEmvc/vWpK+nxSzvILZkNE22E
tV7jMl40Vw73q0wG8Yj5vYrfAwjPKVSJRMbnaX4HYAYgDIbxnN0fWtpx3NP+PpZu
t31eRoR57xHVhmhr9em0aiyzxLpPY1Tf5tPFNtaUf+61oXa3ITBjjSDKUQ8EBhgp
C8jHCCU/vAvXuq749byAnvfjGe+5XRdpd5ahVh4tYvJbQJFMBphiszdcc+c1T3km
lGVHtmexCHNDHUtnOIgHCA0CQWiIZgCTcYIGh7YNgGaunWlnUOxV0VewcfqOc3oV
qVFIuLvDN+lOGF2O8aMWZ0oSfaK5wPwtZBZWQMt314QVKcaHEKD3/FJ335zb6ZWp
lFH8cOtMmkKziJLfbLvbF8mRAw622iVoh5tJgAI4fTw+b1zw2IbOm6HNEtdUCit4
VFYm6maa1T/6cjz5VvnlehO6xCte2INqN97vovBdCL9JGQnAznswlRN89IEblpmw
o/PFjixw4AQUwIMUWRRPH0d7fs4Q2rbkj4laktJ52Ni0igJ4AQS1uNgAq/Vdo/WI
QK+5CFMnJKhjuxusDVZYESznFMjyTluu/97ltVVHlDE+oSum0MuF2ErxKXsa7Ir8
PZ7Jj1eyWXzShHXFLSmuAtuUz4i4M4VM3PkC3vqbmFHHw5K+d8uo/bMTJOxia/7E
s7yS92QYgBj+K25TtbUOmUObQ1r+QrBGzcVX7hTk5OgkrPIdsaMt2aMExocMLkA2
Iv/75LPi4PKNMfAaTDXjwdwmuzX9TOpb/dYXRLpPfjvPc5fbVZTkKu3NmO0WUEex
FGrVB8RUGzMp4s0RJBsFEhofJLRHSJuK+2BqbAol1aTdih0cPV/ZpVq069tGium9
gWeToxjq025oLkJNYtrOlH7+c0ZMf9EQriiomW6ONFx2S95L5KIfSNDaLqenkPXS
XrEMKTFLrGaYEYAmtPy8PXOJo7r00+LulhKa8FkLRn7KF6q/QLk/j2t3qMembepD
+pnOMUdtPlzAn5oZCCND4fOKffPBLmfv1BsB9Qt29/smHuE1DyY0fa1nAtDEJBqu
+el6JEg2ji3xUm7IzY+YBHSSipQeCC0kh1ar61EZarOiW4de0aYWanNQW2UsXgzL
oJ9j7XypM9KK4ZU40PKkGQuB1IX1D3tk0oguitf/F9hEKu9wvNXWOFRAPkJ7P3zN
Y8yjvQmyxOgtVJ9iJRTlvvaI8pDpPK1r9L3aRML1MUa6KmR/22Mgwzga9dvfQdyJ
F/3qRmHkuc+SDteW+DE/V+TlegdK/axWz4e/Awdh+vDcLPOG3IWS/UMRp5xWYFXE
DiYPjY8CG9TwkXYc1LEWYQ==
`protect END_PROTECTED
