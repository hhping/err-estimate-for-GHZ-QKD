`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nLdeXFJzhwmn6lcAcKF7EfQtrVodNYEkYEtr0Ak8E9FLcPK23T6NscUKx48BGvPP
HPpGkao4VkmxEamDWvMkxkbbVJ2O9KW5Y7czc/qJrWz3AY60B7qrbGmyUo44F5sg
RwSyI03HiaOxBTD0Z7eotVH+jkffuFUJRgxtiB00qtCoRqbr2rZlm3QPpj7JGLLi
urEzIa5j/NwEjFP7295ptIEDwfLHJBghF5xSW/TJzoiiPcBPCvCe7ZUArhwUUQBj
esOZ7Eh9HIjfGkY4yooR/yabHNbwH3GmAi3ImAvLIENSY62R7q3gEMCDBT+ivh0k
jHL8YpJ/1XZ/pySAVJjIuWLokaxqagjmHO2WPiaAO4N+NhWORko4DCb75msUtit9
ueVFebU/4dOwSROJB0NGWZz5wAwC6CVegAn11bGiMjEj56w5M+ONWi9ktdJeKTuA
s5syJPSF8cZq4tdj5zzq4z12sqoLily+k1SiO1TQruquLMryRvHIPH9cy/EAfn80
Uj69pRqpjUVCNpsakVBlTy/BlEt6DKDaOGG4+oWr+Dh81SY+RnPwXJPu8UFy33t8
wljSrIYz5dKFhj2gS8QmD0kSm/RJ8oZcL/eIsyrgB+rfe2n9LgTxldyo0uZioR6g
6/2sjFXDTYYJrmH+e9jQz9gfXU0fwgv8KroZSOXFUX9A4BC4BaAnxf1SI3OtmQgP
MLStywi90rdcHbaMICi03qi8SWwbmSaSHT2PSQJZ221GRR8BGaD+YUY0ehwuQHtD
akpsqVA0F1TsaPaMckbfK9QAlOmmcU5CAtx66HutMiRDEvLKO+gy94LnInCH/9hQ
CckukugSA/423iOkoVPwvA7uq8nOMuB24lQ9WFtzVe9j7oI5zwXpaksxRVGJ9vZn
7hFhFV1quePel5726ZloHNf9D3P755dOizN3Bc0QHN2NrfbFpPiA4dLWVByuRZlS
1tlp76vVW7czmXEKekPVHyh3Ca13rBjn52TRWgquRWbeEXhVlN/BOQHacixIO0Mq
pZIvsd8P9dNPs87otj9UQ35s/pLNnX5a4y425cfstfTOELoxeG+F2jE4zxtqEZMy
T3gvaUaZYVUTTUeQKfnMntfRteu0Sehrh/KbJQgS+jKGgJ6exCbh2+1VzBewmdOb
4eyMe/+aCMlNsyCZ2p4x9IQu9gRVo6uS3fcouU1VM8+ZnOd6lAaP4awJzLXuuTyb
4zEdDNXY697bUmlW9OxY6WKH15DWdliK6tvXbE50eborI9jJ+gV+h+A9lF9RemqN
Z5XsmNKq/2PbGpIwwPXBYMW0C9RH7FLpk2xTrM59K9NRDb7zJgOjmqznMTI6B97u
IIjRwcKJezR70O4xXuQnMsW7mTmLEV+OD1jaL3HnBS5RNFfcXHERbZ9eNcduzsr1
+5WuHgRjljVNGoKHRKVTUkLdHKmNPZ9xy/545oF7qRjHgZRghhwuV+LFazjeV6Cj
M8A91sBbJ0rxvJvjpHEks7QJ1jTum4161rMlsdb4MubMAlhgKttpTOfdyTkf92NY
P8IDE6Es9jBVdcdfA1XnsWjKl8kArT7weitqqo7Z097qV3bkl/RbOav/IwOa7i4v
ivMQf7gkDA8JvIJ/136F/+u10fyYiOmHr5Q95x57FzyxEHPGFa7bmtju7sOS2Lb+
atvUveqAj8iAfoS4iCBVGuBrIoXa+p4jnUu93buXKhbntNpTupWjVHCRPtZYJnwm
RCqLZEbHlsJodyS6kwoFHAJvRZkgQtMMKcHVMU6ZvQnTAX+NRBDXzwcKUycZ8jLO
3/gjx/eAKFAhgUfJVhxqeFV5VUaJibv6J5rQEF1kgal+1Vh9XaiuOheuIB6dSHNJ
do4Zy5juVf5KgEsfkDWBusjlq7wj0iszi6uKI0i3ecaMPK91mnFj6oKQAZdbmN39
eeOv/lp2OWRAx5D4L/nk0SBDpB3vid2NuDszsXSFNW611Rm/RN2Na2yjF345fYed
f+gyeBcgSR6jJ1dE9jgMeCXH+bR7ddfVBYiHpYI1Z176p7V6gSIYw5HOASAnwfxo
R8GAHehVP2zTMx6a2GRDx0eRPS4XhglInM2pePJIjBnffSMRqXDmHY/shuDIXsdF
At87xJ1nvQrt/w7XiUqA/Vbncf1jGo0Ai1jHkfDsFQPJ1dyB537/yM1+YwY1xjIa
eCxJRdyRqelACUS+/qu+5dy6+xu4n46+4aJrSa0mgOyIx3kZxV6P14t5X3YM10kC
jlcXLL6KudbhygJAVKhQE9Q6Gf2ETpACSGskxzJu62vfUzy6A8zQEtOIbsvm7vpC
8iNQU1RYLOtd2z3AOA9u7g+jojTPLmL8zLHckt4pSANXI6C2pLZrvu7skAbGJgVH
2nKtNvje2fY5imvB6BATeh4j+AiYK2mJOW0kD5OTorHHX40aeXewXJdW5EXiftCA
xk2+0XpE627n+RH3dBn8A5Y6RFPnOqbLZ9XtwWrz3AIQD4JMf8PrHiTew2zr23gm
YuevMBjKggYi9iOQVOgJFlIP0sQWtqkzTUlQAzLuYPvvDab1HrltC9+O9MTc4Wch
JGdYdXf3uy1bZC/izVPDbsCYhwRCHOASeEfpY+hsy8sR6vSzpNpy4yxcTcyfW8ov
89Ymtc4po+iTklWgrXg+wXuhCRsDD0ERfWtArE/k6r9koKcn6x2logJEIUsH0phu
UFenuS8ZgPeYoUaMQJfRISGUv+g6ezz9/KTBcQz780BN6gG62DBlBDolENu24y7a
ukvlwG7xAt5SBoLlUcRSjnt8AG2D1EKYLzKyo1U91bgBg8tQcdVti97HbYNPdyqA
ttS+VGV0i0l/PknmzsPRweZ0CCgJVMEpJKDsTakLlm3Ow6NpB/pFa8R1ETC5ubu5
TJBs/NgMj6xK2QYRN1vwiWwfxp9Aow8chJs3kK/I+PhOGYVfalRuYWKq7lU/aJd6
khouF/nZIELeCgrZdwWdIDWHxldWd3HEUokR72okKrE2x5egZ8YTmhIivCuLClxt
odiP15MoNlXS37fPSrR2k9BavkXSaNYRq6KIWhlagEzfnWyJ7jdGH7RDUlieIz2m
0K4CCCii5e3xLHKej5RVEUJNKosgEdGDH831cKk4wdwYMKNGwFBC9uk2dGR50alu
ZouIp35qAt72lvvFXigowy2+bd72iwst7dIFiYs/fuFb4MC0U/MT5yKeS8Lssn97
1ALlsWpBveJk507JdxSfO2nHNn8NaLKsmFURl2/TIdJSVYk81pu/w7dezEYePfzO
lnn5sF8Kf2e3OHEQ92TCpYSCNc5xdtm13bzX277erJEYQ+S2rat9oVhZBrs/z/TZ
Tafkndbc5LmtmgtoP99j3i2CPn5/I6uYdYgMC1m2ptnxFfI2qGJwY3meLTPRijI+
ZUebbfMIn6Qx+cT1Qtc8fzLw1+1j8H6KLZE+YrkWWWaVwgJHRWFrCeNMfjCtrlrd
maTIFFnZU6VrMik7sdEUY+3Nb41hm3Pcx1Qnt0SIlP2UqlQZO3U37t2NMsg17ICQ
csTp1F0EJ0hoChP30iw5Smy0VKG2M0E9XZeDNXo8xgBr1z4YBdbOWEJJQQTFKKc7
hgjSrlnMyKpOjfQe6o2/sIrtriNS3CfKXR1LoSOhKJYju1e2W21VwIx2hVX60mHA
weZau13OQ0z5TFA+E5TWihbd3j2rAad/XXJ2HGeew5SvMOwzkeYgn6W1J8mI313n
6gktGQk0y1MN8WuJD6k/zg1o3h4VO4GuHyCq/JkWIGLEVaVt4ExP0IaeZPtWGuIP
v0AxjHh0LfcD9I+mC8ya+udRzm3BEfRlMeVO+8jArsvWviiUZDxnu3JSKcfoYe63
kuOChD9WwNq3BQ8/b+CTyu+2FhRxyrTjl0jt3JdlGZs4ZWy+3QV99U/5UPZZrV8I
nQuBXW5F1ADQkz0k2OwCRTCPBZoHgczT3cc5Vnc6FF2/ochxhFFlMt/4WtANm7SS
KMoGEniDPztZZr50QnjRHJ3cGijGkShCowGI9+4YX+L0eJi4cVr+3lCQuUwRB3Uy
nBBtJWjjf+7nfOndOrNXXjqxJT9plDvFXyXGRF9OjGF7dVdnQjoFMb74kNR1gRNf
vjgi5kq8ku/RD7pp/RAqLejJRkl7KhVZpPaeOYV9yAj8pK0vU5Yl50/wM8jx++eh
h6VrRAFg4Y6nIIClm4XKT4VT4zfRDE51gjrq8elueLweokV47tgs/JzF6Uq8HjvZ
zyJx/FpKLFwGNspymcZ8ME5aXX4j0tx/15K2x4heK/rHtzQeYy+8ZqL/FvhPMF80
ncu3TZPurRPtl/cHkrqcjbRwthMOaSQXKE+74n3Ttnew/vP7SWS+x0blyTiFlztt
hBASGjgP+obS4v0quj05QxV2wqtXZbdSRL9qSgfrz515xf8D/6unZIzkH0Ah0MG6
ahwk52qQAMH90EbSoJXfY7BdWV0TstCD8FaeGrbVO3uFk92fSjsaqxk0hDUiJrFS
QySzyp1rVfUO8AZx8Oetb09scheGcapc6GnsKeVAJZLX+apAyrKlJt63DGrb8/pU
nRoZx53JV4MhemObn9+pVe2JC3v/0Yz/EmRC/4wBIQ7pItJ3JgC4rZiIi6+/waF1
TETHnGnorOTLjB3fQse9oiKQargEpCKc2yiBzMWTaEYC2RayyvMw+H+Lmxhw+yqJ
KQD9D0QBCNpXGW/9MOorKctIfBVOvq7L7LvHSH6YEg7ikZZgVpk56H0bXfXYlew1
mPJ5RyFomw776C7HXeOA4AEqksG6IAAVYOkUkrLn92yqUz+7G1Sy6I6b2VtMS0Ak
BQGouRMsOafzYYz7z/KfxRelTBFZVUmsA7lsscn7kASVLvZMGzwigYt/XEyyqcZ1
wvctRTr4rAGiq/4ywBh+8QNX8Dl9CiJtWynXdqlnYcFzrrtcbosdxP1yqECJtqIB
dbOAqkG+yNrD3TEDTvb/0sZxJXK2ueEoQ7ewqEliFggI5Cjm2rQsK35cMn0CrCS5
Rba7NeRJnLLH/MVI6W7Y648yelqQMhMKtTMeaB+Cc4v4ZePPH8y95O8oooeSH0OH
iUSdgU4J2yXyEh8Y+8RdtEhHEi9AvQfuSbIdhFCnEfB2Eh65HEVgaXYlugI79TTr
WcS05pprlM3MYpvXOU1cvLvVVNCsr8+J9AOEc03/kCNw5GEASPDDGUgL0ZgEpi/P
m3RASG6YjlHjyVdu9syow/hKAIh3GgKVw9AzaG0dCU6L5X3bNoR1Oj4nPwW5U3v2
oIOF7E2zFNppVxjgUuj2l8n07sY0bXiAPtS6V1tfs6NoCUkFzI68ashhhx8e/Wtt
rzbbEO2yEYP7e04P3Z5tc1+JBzkL2RiDFI5qa+isszrFBa5DMWCg7GcHTMIIFHBR
12NTqtiL/yXr4fBZ24Rd0ubn+SiQQ7tiYaHim3NvSxB9AZi96sI30BZT4QEeC8NU
om0b+YHC0/zQISVm+R4K84dR9UmswIz+/UYHk/DFhFv6lj790hwRjyuYBAgzEcZI
19dbAH5GPUPexqb9Fxk/H2Jog7ZZD/Vy/sZM0aJm0rjSIItk49zMHHosBIJC0TAg
29Iu1lL6RAe8wSxaEDMzMTQaK8+lltG4LGSTVishd0SlDaj4CiTSQoy5VBwcjTH2
obwU19Af5FvwkNHtO0R0IUtdXv6wllNz4Aji2na9udTwkRTSYlzXvfKsQqYRuuwv
U2HWejtOCFPCcLjY3cLFmwTa3Mfm0Oke9PMrXqGu3UTArwq41gGaYA+1mBeF6k4F
fbyugWl0KsZAQA/D5+o7JFoKCch0udCK3t8okJHUOBQlV235RsyCjWfRoxrj0Ow5
5PK/RvFU3Ya2mg2eK49de6Rl1YJtKTmUI2hI3f4uHoUoqluIjdi4gsC8K38iC3/v
dPWKsekAVPtcfZGuwAVksS59UJ5ZvhwZNJuGXZJeaybjTNDbvTJttBGBpThv8xR8
TXd9Zs2AOei2IG4blq+QX3YVUnK8FDj9DrAQrG2iSmqrcJV/sQwHayAhvrRtsiV1
orJ8kur9HJRApzL0SCc0ofwMk/s/s2bd/ONGM50Iq1NeRkqbBkVhK9Q67IAGDW3k
viZeV8dhrIL5I517E14eg917m61DppJXmW5viXFGpyGuOxXPD3528BZGcx4B01hh
QBrfloQ2TcEc3WMhXRHKHG+aM8N0rZcYPGvlWO6Nt5lywOMitlXMtkYbBYbSyzl+
pYU0QeKWnPeTwLZaXpA36anW7286arRam5qw7TSiXiMQUWeJnoe8jHfxQD4+VJV7
JxNnCUQlgur9MiZOWr/sXCvV4afFeX4EZvp7g/M+XyZ+TFb7bxOTnEPDDiCvyEmb
SYJBS7k/CieYHsDf89n37QCeWTY4D0yYZCqn8wyD2iPm4tKOp3DmmvvE5/BBJWQ0
90L+1eMabg2Lm6hpsqZfHGUbwodE3v8NvhcWNG3fNMGt/WSZ7yAbIGKJlwiO+t08
ihceSFvVUhwtSWfQNLW4/ALWDeNiqSlBoI+VY1LhBJsu/HJkIPuf07F7B1JRx0Hw
Jo/G3z55q0xTPcdAMo/vIjZy0d10/JH6zugz7wan729GtKNsDMI4k5trNmhCOYVB
DNfhxkfQVkLk+YV7LwQygSIfke9aWdHMK3EzYmwrBuk21XHR7zZ9uhbizzMmtHcY
TpmBcnHhE6Jg6G+JMpoSz+PSR+OExoYo4rGN/2assnhmt74bdGoZauPX5DEfVVID
KXo2VUm0Hs8Ol6OgCnK0fqQgEa0Ml11T+M429rxk8KeJWZ6nvQlCsIUysuPc8urR
Ks40mPG2pLjNbMyPCDH2b6KNjIKdUN7/mney/kfM8zdbp+C9Y9brVqQWgQiJDRKW
4xOK9JxBTUOJPsUbFouq7C7JEdgrJ4+cyiz7C/yrfWJKAYgYbqEVeeMV9Y8RJzfr
606YCnCIr9kTxw9Pf8gv8Khk+b7dsoFt5VeKyuV6zQ6fFjQVldtpgV1gbNXGR6H7
ArjQFCgqhu/6jyKZHDTAfVuqni586xGq1gHVGs0t7Q194gHRADtYKzIokvxf4Olh
gIbrbok4hbDDktYDDS6lqDUM4YAXdC0NTvLe25LaQuF8X+AC58IsmGDyC2sgiJ03
czQS4NDbuGlA1eG5bvY5czgTE7x9h0KvW8AEd6/PM6xCKm6vhEGjVaEWpAqrOazB
Zh8KbH0PZdZHUY45w9H9f7KwMV4jAhKqn3fL+oThruHdyR7uPL004lJT1paqVxhM
uDROZjSPSMA+zlQ+u2y8dBDbqGgqdJcmfQLy3/yG1mgVpOjP3gI8+BYFUL7A2EKk
RCUFqnJ8Vq5rzXlXQqKpJCof7es8jFcCT7aQ9ChG1w0uAbhhYx8B4v21xnRoFTV2
H2++vTG2T0xTUNGTNVS9clw6IL8eBJLF+WunClXerjt6XW2Ir4u2HRGL37Gi0Tgd
ylSOqS1vSY93g9FxxvMvON7rv+28RzcWnw+Y9HMAEaVfSIvuS8zI381rjzoIVoBY
Aqi91uS0ez1p68xoYF6mwk6/nyFr9m6oAS0H+8NbWBggY6SjW+ART9zaJuRa+OvY
DPcv5J7f9llIXkhut+IcDiu+tIWD0bbO+XCgQ2j7WhVLGldQcsREhMPYgIqdURrf
zXohmnx8Bjpl5XwGPLftLgrFx2cUXSO2P5V2V338UIZqQPaj35os3+7T2vWsdSLv
3umDzOFJMWSm8mqMbMU3P//gm2clbXYdIj4PMoUElxKeC2E5Fbg/upPA/x+Ds4sO
XsyWZgt99BAN/WO9aScUD+F0stqoHJQvi2vTfEvOYRfV9gZ7XEOpqtvE+SYV1fv4
aLV7NZKD0yWlOglzbYS4MGTnmsIlwS9pL8aKqzHy98UvhI4lC/TjEA7wmrGNdRiS
9nf31nvqx8O/+yoXVBuex22pydjLsi6umTvyFnOecQR6SBG84rQfb5kGpCdb9ZyM
3eE/JljDUs1OAlwaVIy9g1XU7lx9o7D5CbaO9z9BjCx4r846S2PJn67ihE0zaiHO
crGznUDsgGny5Y0Yinl/Y4SVtrzrh7foPQp9flXGlj5B6PH3NZ3AmKEcP3DVgYv6
yewxq69zi43e2mXux9jsRTqIa2HzDjWHUyhcvipxJ5jHcVjpR+LBqFdx1+XI5qSR
+UzljT4m7oQ3Tuu+FCPtqi3r6ahQmFzbJjuXVtXBb258dKm1xItqTrdPCKOqhCEG
lGfw1XFjprUxTb31rADVGqtdSERB5xPz850LxwOgITpRoKdTymSFZLXJTZF+yeff
UZy9dOXGPeSLRVEF47bY8NY2zt5AxdzBiSd5Dl1VHmRvlUMsD6VHkoT7WLhxyERX
O20DxNWWeYI9tAYSTmC/coLUNfXEQuckfJf5YPJU6cocllmABQrotyjLJJKmrwQI
oup8daYu8W7Jw0UxsnzUVHJ5rDelfGabdn44tyukMSX9bXKYire3PskXyWWEJUnu
ciDVYcDDnF4EtEmKLCl1aVgaKYeIwpHAXKAZZ2oxckRMpl8blZzMaFNSmsv8wePN
R0bF0R4ARnQLEhq4VAlrmDfzdkrZRCi/8V+a4NrbgyqwzLx3BCnRTFFdPBg90Mg6
2Uqm4aRxVArYfuOHJsYN96CiMrDmhWPI3D6OLZHOYy8OPmi1bCPHoOhfPkvReigq
Q7yrI2qRP+PMYI9ngwlhOa8EGt2x/goP1sPgCwRQ8qeFeKEyvCL33erZX+3kyhuX
WQ01O3ok3eAYc4MuwHOgqnD5dinCx/DtmAY/1cFtsEi5oKYoDzAfwBeTo3X9G5Q6
8IHAkt690I15DfovG7gjqCXNo9JEbQn7Do1dIcA1uQsiiHrOuca0QE1cJqZD9JDi
3F2mURRI11qUpW39KHXuD42Upa0R7JUUO4L8jFh4/IVvnHFHr/4tT2QjptLQTIJN
tSuQtWKChE0mNolxxYrZjoM0JO+CkeOhPY/DjSggYA7TREduQgp77ez2dqwY0G4T
KDpFZhslWkjykcKMUr0vhmx0wnyGvuKBpVezSvG1YTl4NepK+8VgP6Ar+njY3JGm
LDf108CzOpFAzTClX7uWsYE6NJk9IXJfXX66xwjfozIVvzEE/rUvFNf9iXwr9pYI
RxIJw9sges5NFj9dpYCZ1Uv2HxRHZSnnmYAxOqfSjWmWms9cAoZvw/ltrwhwW1BY
gEJptVTD9Nu6Dmf/s4eT+0bevAdk/cef+KzOhiKUskqDcn0VY8fzKGBZu6WpEdyx
st3uOIRH5+X7j+GnlZ0NyWwoIr1+KNRTzGaZgDgGMIiAfdLe5tPjvekxamJFY8xD
4Q5J/zstyfd/I+4KLJdq0JqMiuO96MMQuQLUgFuvTesMdG4z1NEXl/NsJi30Fmh0
X49fCwZ3ZyTCNHWK369KzIunGzAVinw/rGf5hzcAw+FM2NVA48p6Ni2mDXi7wEnY
0WzzUZaQ+/KwQtMFWRcjB6sShnScO/Lymisrl35XSVps7DJiElr/3YNVQOGehu5M
s+jiitHjaR/B+I3pP2X0u5eXqhTFxHmEevPe4Fh2eBGg27uVKy/DIpFCaff7L0om
AHQP8zgQpt0+EO1N3HSYQ9YGB9ANIkm4zGX+FpSZz/Tm7OSgVpcxMae3rpTLPCGa
1NeVergtrrkP4KAz4U3+He0CvHpj6XsKXhirTj6k1noWbKVcSewLj8/hpYzPgqXT
Q2DB0qWHyyrvlSm0HwKwxqeeBAzZZgWhFMtWjY2Ff2Cg9OSPEjfezVP+pH1++o3T
8yO6hRtyIw3+RkcvUoWWG5x0DRT7d/my/McWoRrzA0V/i4Wm/B+KAFNtJR45mzhc
Y3TdSyiD28aqSqMk+FI3GPr6iIdfo36WTdrJcs84sirVQEpIukjOOE4u6GdDWkJi
SgaiEa5JKVCUZmM1cqLKs6LjiYrCQLop6RjYj3W0BAdH0Fh72Cvt1BvrM3CjoFc5
mYyRCx0dyq/HIupQfDuRQfv9BCbgxOMXCVi6qSJzQUrbfaqRAJM2xh4+GV4kgdRC
iY2b41X6K4Cb/xsdTNK3X8TAYgpDQRIoFpfM6eAqIpQcG4m/V+q+YE/GC5OLCWZD
crWe0ZqhSaGkvhwVmUYjr8X25eKT1kOlDfQq9sXRP2RYvlMenNv1goYUUEBweKI7
OPiEqbEW2d+i6eb3IR82UMrriT3p0vG4zWeprWEkNp5q7i2XYuAZipS9N7S98R2J
/Btz3G8oWu1PEm95ifSmYdLRyHV6RZoUKARCKSFtLWuNlAp3eOqqwD/ACj6SaqlN
I2hlur3sxgyvkW7pDCHDhWwZlX5sfQS4NhB91wieAEIfu0wNp3wxyePmZTLGXyVB
z4aqd40Dj237klcnotwhGvICY0cHVdQPwemvq0zL88mZ9oAzAI47w2gSnrujr//l
bQW4O7WnoNLJK1raHBCT9ERoujYrXNJRrZaN8L1N4NUwPJbwLof9V3uLAg5nUE5k
VCmx2FlAV/6sDSLada2VY1ah2hCsXR5mks479fVPHa6OfCQ4UezHCMTXZBqig+O+
1WoZAdy04i8cb2DGL2ECt6RbEKn1ztJllATQIo1pYO43M1KO3nvnWhLDkB2FEVsv
WYz9Ihjl8jZSHh2aAAbnIjX4q4wAd0iPv6RKHGirqC+mtheryRY3iYo18/aoLKGa
eTLsrakeASGccPzsK63Eo4NY1nbWGbmBLy+vTjtrHZ8DGmnpmebVoWpMqm0822IO
VvQ1NFdsOssibHnAnmmTvYVLKFDvaiUDGNsglaEVFU79Go3D+kFAQkBLH9alYaSJ
exX0Wgapn6AJyeaOTVgsb8M+6ASAON+R6vRyM7srjSOfcp69UI9Fm5ruPw90CBPr
eKn6iWXx4iZqbjuCIukQ+k7qkep8abLrX1SO4wISI1l2MlwnXXBpS/juI9EYGq7I
ADX/ToHj89coW+4TcWZVW+R8nFNFQLs+SrscWx6lLhjgidPzgnDkUYDE0btG9Uuy
P/UThIn+Fv7YW+FkvwPutkAsKTNX3pHI7GSoQaYFPWzPb8kEZM+7b8th9pC5MOXd
ftagkm6o0W5hFgYv4/Zyu4XHjwXOGlzrftNdX7ladYREHTpNxWa+2orCVnkKlg/C
+emaomEt8OwSRxEKA9j6QXk4mdBGOJqjR70dZ03h3QZl5Xi22qGayHG/LbNig5ic
AGVKQwDfYqC+HNo2pDZ1GJMNpZDuPXoErc9/+2IMrAoqG+wbEYJUGS2fKg+DksgA
2iKMs/i6EH+VSqo/+cuorWG54unJRjkJiKFHM5dA60tzMMqcy344GVqVqHbaEgc7
uOBFlHNNVvDNSdGBYB4Los5SPvelIA8aguYtHV2IoAV9tZH7MIq7XQadEhDH/b+w
tCH35numEPNOCycvbb+Mfdsje7argmdSefMh2WCjvngQ0IYHWsNbaArHGpBgVFQZ
E4Tl/lYYDZrw9X5mkZHfmPtRdp+XwGOo5PgvawYFcVIQTgARkMVllI9v5ewifgdQ
L6nahx6o8FDAImrMdLHOONzryNY3KDkfVvok0WOk+uG0ePIO27ESlubLVMEeDDJ/
ucfvvkN/aGyjyKoFlupMB6iqDnEkmiGRFEKaSNGEfy+Z7vs2K0e3bHOtFvcULE2L
Jaem/5Bxj5ydU+zjbgkF/BVevcKDsnFaLT0jcdvvCfDvaT0R+LaPsIAAEfTDCktI
Y4mCpVZoZ1tO6QFtaxm8wtns/LYhIWKAXsFfZEXcH/rTbSt72ptdyxZNM1eeP9D9
y+vXfPFu66zRzlcdP2asrx+cm6foUXet14ZxibsIxsDrwDh3AsIBXTnh2Qr/1oTi
5HzYbfMx/7nbLI6DqrAD12oOs7XKBi5BGwD0gR9AmsX6JNlWCnQJh5fLsPYFWDyT
RwsB2obMKBFWLQcnE1I90zOcoYStCLM+7geDhXUqwZcbG48EJdalHD2VLdcYZLZ1
ArqcoCfP54M0sfv/wG37JtBIMdn7ncpx1g0b3Y0iKRWJ7Jl825EYQFOSOb8/hpmS
Q1ICN8KaCU3YBjSH9wdKgBy+xp/klmZiXkr/W1DHzcDHZj+8EPAlPxJMZ1bJ2h3M
MqkN2IpDvh8eJLOYk+V0PVrO1XFL2cnss7rMBvNXdPJ9dKoSZJFZ897sWNEmdl/Z
BUqa5dvNlgNI5bXNq5Meo+dCIM5IqFa64C9KVQxtenbPuBUEaPK/AkUd1divyr5W
swkng3kn0vHkCI2/qPsi7VI38Fd9DxP73vrk3WlKc/TwpFQVVz5JJYxVwhP0SmY6
lUbo2K2vYOw+3AMfLmjQwa0qbZIQJQx6zLEcwpvConso115b3vkUSEYPH5A++aeE
MaX1lvi5oJDOetPRBKlHX+1ziIzvW7t8NJ9U4HV0NiLuR9oCKXz3dKG1VpK/HmEt
dEKmVVvyO9uzpJHlxnyf3b4BglLrCZRTSGRsdU+TERMnDehWfns+aC1Oj+4AMlqT
rb05HNy0eR0y4dnIPknxOeV9swbL4sjlNte+iD7Ib/q+Dc5qac0bluxRHz/RhyC0
gbzNSf4sKzYFAcqGnFr0/umijTXn9D0Hid+yyCmkaL+LqQ7Naug+YAyeiOTXIC53
O510I+V89WpJcwwHHUfcxfu74KAkXTh1uiiQO+r7LXr7qSFeaClB1W55H+QuvN+l
KgXFBIvWwu8MeQWX0VoEEw8x6R/Th3VbdltEkcq+6NwW9fAKrkYFBMHVL7YdE2OK
FXfzt7j5iVyMQRwoZBL+Mub+s3ZN4l3bEE9EgKs71SFGM1kfPoe0fqAdY5PSJovG
ZvrmS65MppqUYhJRjD8vSr32Wlq2rhdEbUsF/XzXUaxFjG7AMFrzA/t6D8jWFnIX
PAANpPCSHmFIKt+Bpjzj7le3U0PdkyyIRYC10rFdYnkRFIO8W/l4xCB4aYWNxN/5
EiIP9Wl8WBGKXzrYr6J7/osILtRlaQByhOaPYc94I+79VnUmYVVdag7WEyI7Bcuv
csq6638lC82vtE5/lXBZ9nnJ+3/jgG8KXWX0hJVrNpQ4pPj8Ny/nFnc1BN18ZxCq
diFCsB37h+G2i4nk7ykrPqNRqORAt2Ua4chhDBFlr/rqvGBrrpiy5amWL93GXPpq
V/VBc/OIPfr9cDa+xVNT9yAE8JrbkoxEebdyv19HAmxs7ldLKtJqAAmjyPBqngPt
dL8Nj0K+3uQI4RPAGdJKbBKApaBEy6WwMcQIRijlmfeQHcOZQHGo+mU2pEU3D8K0
WsYAB24yanLm/96qDwa6UIntDFy0btIkfuglzwWBx6F+fxOLXzDLRjv9SlSY5+mQ
PZboYrhvz9RD0yebEAUUMff9hSJkg8jxmnGn7pgfWSFUxprXKowDH37PvWYNOdl1
0TP8HM4FKQwC6lmAPsdTxAm7pf92PHP+ELQ3be87ld6LMXYnBGaoj3hwqIVFi8SQ
dYdoePC9fbMJGBnX8NtZYSvnyFovR/LyLRo085fbZjgU7ph3EhUIPXq9ulsaKFc2
lf21hgNqnSTU8D9UeLiVgHC7xF7LHEdR1TxT3WWAoxEyCR8Y361rJUgmbsEShR9N
cina1H2r39hUNSDHiupFsqqs/XBRKCxHf/QxIDaJFAoU1eVQRmbuBz+k2T3L08ml
v2X4gOaMevG1F5FdgD9D7Okcfp44Roxzkc9O9J/8cCx56c88cavQCqfFAC/wi1G0
AvzjOraJH05peX/BHuF97pGaFS/masj7GeKE1wTjs5Ly7C44ykOLeFej6jg4+z6a
5m+8jg4HCz8Yxt5rJFQluQ41OUWHRWTABDpwovAvO74WIyzGZV0ddYcOLc9K7faw
ORc4UBpyE0kJVMU7dhdtav115Qut6dJaLU8Exm0dCNMcYlyQXMVoJ9bh3PT/nJ7z
iqdSASMCKbg2suuuRvlvnRVAv0pK1FRYkdX8l0Bhpw8B+54MMW9iuMNtTSz3UbUc
SyY+ooosWmFoJPEMeesiSpKbt6KjpXUKcKsQSvfONbc+p5tEOU7z9brUQ8CMoifC
sIauqyjzoRMw4/H/UoHCYAGwkSsz2qz/ca4OiLpmmi+pyKKfMw6zXDMLU/ixVNdi
Iew9J3jmRpyw7SuN5bbi60GAF6nv7tdmO8RFPdWwnKWFl/xbHq4TavMnj8r+e0i2
VFqhr5OZAjU/Htgot/PpUbz81AunF59IlEBhdCf5ssn3DI2MGA95tds+axYnNycE
IINCxkAo+TeC++lCfjsZ0dKHLRxhaKU+imXD/ZPQnAuTkbbPZZd0IYH0oiDRFbND
tYGHZlDNlCGbZINyRkbJV1j/jbHdbmYX2zCuRr1jLWJ6GiRQkikY//7DXbm4Y+qp
TAZlbi+MDXG7aNze+zOrduC7tz4ZSDWaWYmuqzh1VXmGCrii4SEg/u1RqLSH3Fkr
3obAisjP5K6II7V9WB8diFbEctXQBlwfdDxWHDV96JDYvXZVT7UgLEwW0e1x+XYz
EficuXL9F/GM89WRdXtfefXDjhyf3CYoNwATiutp86ZTvfV9KxDtooHkjTkR6A+z
8449wxAjpQ72D7t23c4wJ6OhXciBfDMSxpi1pX7n6BHVf90Ug4oquPZc9w2SmdUt
3AKQpV1uockqehx5fMOLaz1008Iny5f6c8ZCHhEYh7/ed3rtxcTkszMh4iCncujJ
LoPpttSiDjL6cOdDz2kb+w2ZSv/TzpYlpZpFPh7BCSabecu0/6AeGEnipxooTeAo
0i+oB3vxOqU26Ois/Bj6YR6wS+V2mdYNuLFQOXlkVEvFMmUKX/JUN1UPqbBzfi75
9x1bj6kU1c1VBw8rJpWQNQ0Y+ewq6L2V1hvsgkzs1qiXnf8+LjrV4fcuHLUeFEBb
FOvxJYIhRvJbt4LA8colpm4rOAjOikbGJQYqGFFauNEBo4MPtA4MPzoe6LDeBVon
C+OOT96SKoj6BUDTZAUUlSrtjTgb/DHYJZLSoCVBCRl5ZcUKMVoq5RB29kxGd72D
s397xVup6ldUm84Mw7M7rHDjncq21q/MKJ1PHstxQJN77xKPo04ZoR4Xl6+eQE9y
4BAkY3SlA90gvq8AD62RGXqS7roQ6bwWTXDaljCSxQIhNb0M+GQhDjrv2IxEiO7c
tj667I2+cVDlqOLXZLzH47wzv55QKConOjEEhrdm3MkDK6DhiDi+byXUshu35reM
mBhL06yXzN6U0PFMMkWSulv/9sSuA2KBdjygSrJe0+8ZkBRQD1yyv2jhDWcdOyCn
WKbGPXlk6v8OphjNXdOt5hgWMNIwCTmFDlLPs2kG0WZUBwB17szlax+rDtJS4SfZ
OlwGN+D/M28fh8hXpPiVOYXFcY2G9OfBM0+2AmvQZHThbIKQZ2icL9EVo7UL3HXq
XhT47AFDmbZZBIAIXl/Qxrj6JvXEK3cTGs5xigXOvXUNK+/xsaI35n1WSVTanlHX
vRl9Jav/amWpRx9MTEF756yiPwL8fxYuEyz0xhIj2vca8GvD2dH8AS9j6i4yZNbr
gvs6B4Ec/Fvl2BeWzVwDXak4TKGtW37qFZD82qBAkT9xwD62yLQeOND2GXGzcP9o
PakXKz8oP6PnNHeEHvJ82qHPaaN9MUQ2fTTZyWOU9r9co80GWgu4doD4bxZqZLls
kwmL5tUUpiVomvkIDPmITWhBgubR10+dVXrrdY7pttGxzDeIWX3ZsUKkWg6++HUD
F99qISZkWDoJTOtt4R2WxemMurEBElzkWDjSB+MqZ3/Nq+xJN0iEQbVrURamvRNH
J0fTbO63DWw2XynyAQ3NMrGQ5OxYFsmx9Twp6UteUzI3rZrXdf0dE7pA9GPwLvmR
PEL+k7szl/Dmht1vG4u9dugIjvpM8xZo3ONqu7xpOfazflEPxO/iEuQ1xNDmchbg
tIciH2agHysM/qzqUIRlzmaCXT8lSrWrBXTpsSMNL02otnqKbY2hPeX4WrLziMv7
p+JS+7Vu+ZkjAjU3+tjJRkDtQO/DBhVgLEyC4x6Wc2Tu/SybeSEYvfSuBxOD4nJT
9APOwVs9HSbl4OqyRXfsdfN+jENA/lCWH0IzloLPRmaYBqhnf98ikB81evb/OGeI
9RXN3wF+7BX1bLWOlQe7ooyHLCxif0NBXjNE3p2W5iiUmqwQvs8xaOpMb0Gv8wyC
V84ZfSqvoVp1zw3VrC73+4FPTPgpiurjAfRAPXrera7omFJbhS7hVYPx9lsQVC61
F4UJ6VQHKAKe4GHV/pylDN/9gAF6+bT1O3sf+N4F2NzvgIFrZcZcGsmKOf4BcMww
vk9QnWk/zPEShOFX1EdTXf4vUERGpmwFxLPDO8ipfvJsa48Eic7tov1IrUk59dJr
Gg5L5WQBELAXFNla9YJjPWlTa2Mh2lZbN8I2mWYEQlbUJAODtHhimh2R3j/xZ8Dh
H2eb2beOIo08phGMYbYdpNGXV6kFpEumOuZkeLsskgubO9YtLRh7CvxycPxZz7Fo
256vGJoiEnMFivL15VkhcDHYLprKk4mX5srHILMhFHsf6ZLGqKZYm/gvfpgUSdQ1
PqJXJ5TGWaVWp93Bsm2Y/V9hzx4WlwOlXXt73eHwqzR/d4ta9bciHYrsJ0HAIhOk
X3JEi1AIPLBoTZHT80atu5opiVJMtnwFndT+p7FCTvKMo/0Gs0KyCK21hbU4tvpQ
FsUwgX1nCzn5HHTQlRpBvUyWdMe47YBi+ocUyRek5tOVftcgcq6GQeibUhfj/Clg
pST5avlyRZm5eWD/xq7NzMBuFtN0ZXoztGYU8qsr8UBFMpM2zzanx9OMJyMHT4Da
EhN7cWFw8zvtmOTmzESpncSQILj4SEytpyZF2qoLWRG8bHHd24BjoAg4w7pvyrkt
JBukEABFHw26I3FTXZb/PNG82IAkqBdAqD7b5tBYxJpUydifzO5OHHLNyQnTs19s
0Lvf0ytYE/U8eLNHD4zX5PYJraKNAprVyjeefYCMaBSa92FgiMNGl9erb3ACtVSr
Gc30LHTiEa3BJ1GVkNG9cAtS8p4YudGILEFXCGzGaL/17H+eXCrnbGNheRYQzEWS
vAQu1BeVmarG1njBj8/hLD3xJo6L8YWe6Jjiiwqnn2hgVz7F0s+aZD24tpwfihXW
NYwYG+d+MIujdpovvGkR8VCvU59MYjbOVBM0SyNsZGHUx9g1j0B+pfr6lHSqjhX/
2FL0DoDzmPH1ZLg9ZWSfreoDGtkiJIy8i8ixqnAeGjH4FD3DBo3eT2YpK0B2G7e4
r0uEjAvgi2C4BDbFWHlQwUsy4/jx0WYgssb4eMKIpBh7OwcGq4p4c2GXg/CiL2BA
muzmdrD1f9G/8M0q+1qBHxC6/0uciDRVwamp+VBpKVw8yq71M2+krJjr3SR9WSN6
7WlFgT+090CossewoZvIVpw0KDohBpQ4msQqWPfhcacUm7AUO2tIXenl1OJkGl04
YQbhsuWd/zcE4kU9m6N2Dww50Pn59bqQ+oKTq5utkYSUIJxR8BtLUrGi5F6pkhr4
Y4i0jTnAQByvq+HkLLSA4TTpAeJoUp6sR7Uh0RvQacuGAI0CPyunb8TubTDgyMZA
IbxGQQkzHcS6tb8MSzIrX+bfC3aWiL02gdFyUTsMbtM38hlf52+TXRn1qMBSs6Ey
flGfStVkCcU//S2iC6ecxQ1J+liyL27FCQnR1oO4BexMnNdAPPJeCaFJbGf601cA
psc/dY6+u4YBcOptlf9a2paruy4BGZSm8PKZkxZ9IXjuFK85U5qCw3HJIAeVV6Pr
1065ozuEsJHAGmVdDI8J6ihwFPRR4XaOnLLpPEVLX6RDPspUkAvKVDNbCAxy6XC/
+XfrlfBdFlNVE6iAmbD7xaf4tUAZKX04PnHqJilHh5dzH11RqOpcbZE59BX+vXVy
pJfSxkD/pg9pLa+TX4S45DF9SgHbZSLlDFO4NQ8nXjRirqa/9PuQ+NkVflEjjQTb
hWmamFVcCNT2vvCRylZa+VgS2bzYq4wADt5GFUl15qzwm04LhoTdihbX5QDAnYMD
CjwYQFtsUp3zI/b6R7LYn65yqoidHRZz1JxBv7jdhW+Zn3ULPtl+U4Am6vQwIEaH
oM/FkD33obGpvz0Wec1qpiziXL53g5DXAJLAel6F4bKjfZXj/0rMf4LU8SoD9DYH
OqBA0SBIHAoYzWVtMaKRYSPdHbJqK6gRNOagKe3jxRXjhYs5bYxRLU3Qu4PDbMKf
NBY4FpStTh2LzUqhxYT7CDg/yG1YIYceyIpNCtAm02bis9hB7lvejmcirJtKnJw+
OSxHDsvd7Gkc0VHga8avV1aGR9ti8MxA5WkTUmlevzLYv52RPa0IZIlzZffxuxpc
+Vcdh9YzjBn2igZxSiyZsFRQ276Z18Rr6VJpDRvKXNrihHCLhW+H/vqDqSv1PrLj
OMqtKWr7x46rkjSKvQFANTS/9YpgBBMJ8N17OVpjxlKxAiuNS2epXACl0nTgjiJh
h1YwHIjcIU7n2YCPWEZyo379DSNcRn/SHZL0VbRQfuKsl3yiohNkmYbz63OCot8N
yGcFtI1tJbRSU/gn5STodlvNwNMTF1Dn+tpKtILVJRjK8NO/PQ4htDQZlh3Y/D9C
qPLWZBd2Ia2dzj0jfe382yq0bzRnkUesdevH9LTRmLV4WWi5JO6jqJ/HOHhvW2QM
f2RhwYNTTW/c5pV4dPaocBg0CDk6GboOs5r5O0cgK90pjRXoyB48CBISkKKPB1hr
lUFE1BgZDnpJjqEoBpGcthRk+3t8f7YnBIn68D8oRjqdWaN1ZuF9ZO31VlI+IuMv
rxFRmmKA/861kMgoE1o4Y3Zt38X92B2u1/XTqabFnM/UBSjkNeoBtosgGT4a8wTl
6cgt2UYRvmrACt7aiYR88aC4u+PqYEUW3aRoZOxcxAmsR0cUCxRwsegwd8O8/XxC
IvPudfGLrc+yuN9eCbd3scFg/eJRB0yXYKvbViNOHAt49mSGKxP55hmRIweg3JQc
xio3LmExu2bK3QEkAlFkksiHN2gBcgtQ+/8q0VXdz/+Pp17dPfROxfGHuOMje4tA
Ip/sQVrnBRscFEcFLQL/IebsbzV2+qmx4mj7tP7l3RMa1nnplSixRJSFVL0zdim4
QO2khe4IR44u9v+44heNW3aXVjVDYuM9j+a7L4nLmNZw+FYqcozqF8SnXTOQ3duO
094HXpIBbwZ7bHfVwt6N7FA/nWM7jr656AWsX6NxNPJz5R2UiWMmKTb4DG11a066
GoLSs3mVhPvCUR0/ffLJU2Cnx94l2e0vgdPEfURoJhSeVb4Jc1lgGLS7y5RR9GtP
C9EO6/D1N41uoMcLRVvds6PeixGm/Yat8av+MuOlD4Xl5UVY8HbJR5BaBpEsuiCX
c8oAbHMmV4Pzln2mICq6pXAC3NAYfkatNbcXly64+/3iCkB8aY+Fpwl6SKHOl79k
aqyiamINXKZsym1Nd/EvW1DYkpWyOZX5KKEO7fDQpOp5c4HkFIab5xNl0AAKDgND
hkNZiAyv4DDAB4Zg21HEpVeFzi7vLUhBgJCnfOdff6X/Ajrx7vnkNiuCkgYcvv8d
kW+3jndx1zw9z6LYYG7Shtjwls1NpiG6l3atH/z7kwmDvxcEymcWdNdFflzdzRTc
xOhXyJIXNZN8Z7StKa8P/EZmqXOfsx+nF4YTAMaCwB+WnxJPzDOBtkALApVA07/y
2fYQE2THO6tQg4UxX9uSYyXC46xY5cGKpe2sjNybOww1ACQBxULHPT92Q1XnhvCN
Aj+8ROdwzcM6sviWeyYq2ZzRTlYGyHCTtKBVFUd13UatPcv5+Pf8U3feNQ1ZEXqv
LZ1jd4jqgnP/1YYzS8Dl1oHRv1koHucH8nsunh8nDLw0roVh5old0hiNYTMDyZ/a
6RMcfUvpJA/La8PARFeCEMD9g3iboQZG0E3I6pvfOCRoOajYAktbit1d5gKq3FPF
3q/b+9bCyjPX/nhwiYQQsJhEoH/czkJ7z1/AMVB3jLorhQZXloeWPd3s7z8juwzp
YxerCJayC59dFbFEMSwByWM7Sgj89aJHXHfOfYQ4byr+5BdwukZ9vatav2iKIK3M
ZMl52dBj+9YsUNgJ9ukVxK7qZehIS2CmRWVgcivcabJVbqaTaF5ADCzrVtBFTXFN
tvBkOdVu1uyy623u0p2GmXqtPpTYLXMvP1DWjW/YS+sBY3q4MHLctZKTe17lKh3h
HM6C+zSxkoaN/FQLNeIi+3w9mNoTK5/0GVoTL2gIvDZ20rHMjFBaLK+n+CHfMUi/
ieWY1U2K4wsapgwFWDJOMF2Ai49W9mnfVgSygXDRib8FrzPTWr+/6mm0tv+Uxfvs
Q56Y4MQtChNwY65roZJ+zJwDqW6JiQtrXVK3+hGfak3zBqq8xlRYUz52sA5/TGOW
WYiztgUP/LFcntjmV0stBcSgToZDY6b4+z6nxCa+ECeLkBeZxzXGErg6D4s15WKa
sPPjcHSEONWndpZu5GV+EHLIeSXfwh5CFy2Qi1FqUzHrfPB+u2rszMGLWdiypzoG
NGh+v9SsSJMiBEDfnSHyPFrBJUa+KY9+F3oKqDfxVBGSM1ZuE0U7UBPllJ23FoT8
1ULnbwbY0W07RmclrD5c7qKFq4lrh5uw+Zcw2jlymdFiQAocj/vwCiHfDHbNzDZN
rAmpovXdacKgsNb1Igl0EtLfFy9GeFkCQQhpz9LcKEBmrUaj9CxzGmjacaOECf+M
KWvH4ZZKliSnitmANVcmeEKIFmgy23OHyDiDtvBSazDV8B7PH/uQqYk1qI65BhMA
BogL9gKiVguu87eWqAZ1ldZRftxkHXUFMW1njNn3U6Y2G6qKh6HVjT8s+XoG3XxX
5/ecTmrInpx015ubL1KrY0K0eHowHUL/XRl1iVr97LOxI13Sso3URE7xSY3tmBE0
2+rGo+GvsEVa7dCU9PURO+gRIQUTDmFYpahrM9dBPhZLjG5azXPy96ycyhC4siR7
1gbeoZd1YzTdiFfB79tSzgJhHykreE0+F6bph8jTkx5OALFndzI+s8f95dkVZGRf
nl6FxNTiQhrgg19oHVnNy65N1ihtWmAe3/q29iVZH/PA3G/nqF0FdkZurXC0BBV3
1ZRbC06ALQ72JZZCxJ3RAYL2P0dT4mJYL9GzdeXeH8RI5qS9laHHFZEVHc5yV56h
sCplDRJARf7h1OECVxdO4E9QXACEPmHBSACxSjwq+LX2HBmWRwmuef7K6yShy7xZ
Nz+wXSD8JnrBB2WS0DxBuQkhBeKwUOM5llQrTtPhxx0/r78llmDkdmr0hSKBA7i3
R2mW3m9HmyR0vH19sTXI2Dd0j87IUaLPNwmsAAql5gVUyK7j7RcH1Lx9vIOaApcn
WIy1C4Q+w3BJIHnALWXEGHwQjhOU3rvDtzK3xz7Ys2nC9yDqRTrAmCDko4fLkorY
oXbxmy5zO/d4wlvwJ0CcE539MxZUP2W/r/dgWGBvX3Ud5oQZaUnqcttK4qeZsgO1
OEFRE8tPUGBWhLJw4LKV588NHc9lm6CKIlLHfR3Ve4rzFCkBJ0F2fWSv6HhVyDed
/w877l5EkQxbxaAxcQmg7ircUJ0dw+sQRYekH0M5Gdlw4T8RQPIDuBUx302MYWcc
dw8VqMl8g4WsiOCqJRazHpE2w26lH2nkAQ6vDmB7959iylgEDPM9uH6CPE82Y29x
5OleSoccIf9bHEpawZCM0OYHPoOtFG7bhMjeW0aryZwGOuYsciNN3Jrm2+3D8zwU
X4JL7JXWlLgQASh1lcH0PGTHpVAqeJbEJDfFFGvzqHN/1iNyuTFSbu+7IkP3oLR3
z/QW1hBenRoy+sOicIEhMAY8IGwcNid5UFDYktmc6+DdeThGHijFamA+ywWvCreH
LU61h6TkLoxQhieMI627A42ypMrQc8rGLcSxYKQbPI5fdW2ibkZa4vPmtpJaYfZ4
Qs6rbR23OmwtCX8cFBHU5fh41Akf4qtN4UF6EilelYHYAT6PrR+KLCkmTY62SG7Z
x37QuLq4cfRwUw9g10NBezUicg8Ih2T44cVqKITYbpdUHdNNtQjDt4Q2IqkdNWY7
vYBbYxSN7rGxmz1hle3S5x15yQkRY48zyneB9iJomK1nLQ3SlIkMmiNoaLkgP6ju
MhlV643gG7tGgjhTOfYVbbgZQWXc/uKL6eZXixxih66Mb/j7zWcP8CNtddgirJA+
uboR1FaMd3gKgv00rcAcgB0q7nLiZML4aCR+8lUtFpALhTMElilrwJG2FL0yu6JP
L2zANtiNkO4arjoG1wz9DT6RITcqBFt6tPhqWYTAVBpeUXp94ComA+H96n7Doigq
mYBm1sm4rvsV1AnaBJldsdGjPTBQ9mle5dlkfT/u7Pqx9OY1fHIXXRWAbM6KM6gl
Q0mw4SViNfCnl82ah/HYcmqNeX3trTvwYdde6iDu4v1X1E9XuNvsdFkFBDK26tMv
U0hEEnH6nXvPGI916OaS8/tOiOFQ2aUWyQy0w76r83Jid/dS9a+5Wzenjg7MkZhD
x+Jv3RDG6llP+iqYgRUsobKX3CVG8rj2zq9aTRNW9p8UksH81T8jAVssgf0pI/MQ
SWXf3cyimnPMRkvUNZVPqHvJI4+G8z2S9zjwQYQEYtzYJZXnYAwmlkr8beTIvXdG
LUfOJY1fmqVEe1pms/T6IjCc/dM76VZJxxd2OcoqV6nsSsPRkdkr5aaEvDdcI8or
NiKP2HqQb9uTBaM96kYLaiT+wdxmCSirTrDNXuc+DN9HcMdLrA9K0QB0TfIHCkoS
1voVzL74uTL2yrU/QsPiOYDvLLsvCAPuW52eqk3ksVMvF+0iwcjpnAj0kzJliGOD
EakM0NHQsn3Xyf4Bp6QoVLCMra+OG6BHHMI2zdndv+3/GwxooJp/Yp6oEcVySEzp
rN1i/3iRsA4ybE6ir+YcOyL3P+FWZcrvERC7wxAVDxgkFf5FvqpYlQRsjHK/qkyE
Im7D5f+uqt96zjpk0Qzu/dDv2+e4KftxDAjCCUOd5dhCkhvfW9Ji4PH9mP1vHmwR
BpREsJlRrQ3OWZ7sx8YzGALsFKbrOnC4nMlSdKZ75MxStucUYhxWfocCK/Z0f45e
F25ptFKOSVZSKdiKS+n7QxTqdUCKRh29vr24VFmBuEvg8jE/kmwT6ynLrOGCRQp7
c8/UIEaVlTKfBUg3c9ug2PWCbVV8sx48dq8nVw2SSRoNz4XuC95q7yO+Z1VMjz3z
RFvT1HN6eWzvWcYGHkQy8crr0FGWGHW9RNOx23FFhQyQ8ix4XP1emnHS5Mb/ipK4
riOo29sElNIivi+j4lkYbqBgGQihO1CywN+/OAMW+CWEQkZw55IZdVD0sM+UAiiF
GUvrr4pOKwDfR7FvCs1Yfi1QL3WLR98y+Q33C3ZCue+0rAim4+H2ZXAtNX47bwsT
599MdSbYE7yqTl5CyP0SEwrnZkpUn5tu1z6PlgY4HrUCHWGmC7syWNCzyRpqYM6V
HDsGwn5uboXhv1tvbWqQpkw9/dh+dYjsmYQFGbOpib+mMczOew1tLJMpEoXzWxFm
pzAbArkVWKHgdt8NEO6kAyM2Zf9GQGO6zjDcvqKpvqQm4HeC0pRt/GjMqla/gRoe
Grnie41cWMY/WidOFkWPicm3MFpVR3ca9JeV/eggKa49AxqwAZ0s4r/ZEdd1SfZL
3ksWr696VAY4CsuDm5MGdJuoWpIKe43KUp3o4yRzLhaj9mNRukfA5io39ZC6zAJU
RPaMWbvxq0jEqn0tq2Vq/yTPDBhpCTEtsY79oTn5IEEexHbwNoWp3f0xmOaGYuLk
G+dosE+F5japNj6pc7LtLspX5oy2pmcMxLx8XypZ9k9ssFSQdMKPFfoFbi44hgIl
wv2amabZkXA8Ipgr3VXsM7I0jvqlUZMaRT0SOKvgLaRSi4t8V+9UMnyN+b/l6QRn
UhqMJYFSzlAOjLyD6yln2W3Ya6heiV4o13yYupApoPsJpvuD/wIblRVWA8CV+ry/
PLc6NylzT/kEwReuzQ0WWl/lzRCoX/mUh/SwHvBtTw+iBSss8JOc1rztUeb7eeRu
imPgjNG0YWt73KYd+XpbimbIQudLBCABURvJrBN0drhdVRsWY1HNSuSFbHjyCZb8
/nqRvOEftjYG/+uTFxW5cgZD5pDRzrCPPBCorwdaHtlgWUGO5mhaJrba6omJdoNr
Kpx3ImWKMl1jYbqLXe/99Yl37RU70jrhbbo9/ruPpHr7t4AWDE+3sEWmxBLQGZMX
I0NQdyGsi/fsebqcsrgj/UL8w+/ByKIvykgF2s7g74bEdjyaaL5vPSG5Mn/AK1EC
ea1wVbHu2GC0X8sRZulctji5PV/cTMcAzP8V7U1QZJYyf9PjTpcJT0Nla1ZVBbrY
G+Hhj1/leKHkTtv7d2QOMw2vbjaoTPBe4JBKrwh7iSlLJ3FhV6L8MQegElbDZvOr
pApHOKqRP1Qyp0K7ogdcY2TpklXN6IPAHARuEVHbmOa3LyzCQFjLTEzMyg3vJwb1
XkT47GpixCXsICARP4WinLJvlQiM202+LryR8nPAZS6kOGlRw3O5S7TITITIVZgt
DOXSqGqFZdvtSTq1hM0ZHcwTqG9PyWWNPbH3ar1dDlHnRYZ4y9ZFphsSnY3DUjkN
MuFvZFRdo/znijU6B5k59nsp+KThdbTFBF1xJNWvm1e5pDrh1LO+OXzxnWXi5+yQ
Q3aBj4Hxsb0fszHnrjL71qJ8MR3myYLekNP+LDniTbhEgd93bNUVVdfHlc+3Gn7P
8jHODXoLVoCEqpR4EpBFaR2x8c5fqVLJiFr9IGxKul8rdhAD5O1Htc6E48tNxBzr
DYRFII66mJVNcccnOI+Aan3+8Sm0L41g/9u7LAxPBU5sZqBIHRDwkMqIdP/fv+Ng
sPoZwC8z/GuxjG5aCEOYT0Kj3VFeEPR+GDmmL2JX4SS9Z0eK9tHXKpW9gO7VmuEe
XHGOVE64TttP1zD9m2NW0AwI0qc3k3VXh0WXX57dZH7mO5AupCi0EJiRdOaXEG0Y
FeAJfdKqthpzdVz+UvfkzfirTYVJUzMk8gLa1Vz2nzaaIRCWZjL3HrgLvUaDxPT+
1qs2xask1SV522A7xubWVULddak6FOuCLFJrqL+vYjXtWcsiw1QtLc9LWt1Klki7
XvOVGwz5ht6Ujr6PTkgbjnN3afTOrl934bZ5d4b/sKfUbg9nda4qUo0pTeLSBsT5
HQwEG8Am4fwWTqITpByesQoZXGr41eVS/Ttx6kM934UsD11Qdt4wVJ6lwT1HE9sW
l7Edlio3DZF6vASybv8/KEqYgRut3i4c9p40KeVV3YRFMxD0OJ1g5DUPPL6WGG/N
A6dKJBNpj0K9gwOMN6FYV4EQOfP9dCpccodsn0OX5ZPVgj4lwQtnawlD4kqGY/zv
V4HXjYAD9QM6ItTk8+eJNR/r+7NmQv2i6jZZMdcwKhD2w4pTiu8uikxxwjYLkmTb
aRY1QnJdYf034Z4QhQQVU0JpqGFlsLOjuzO0UxvC0yA+hb0NCaE428lJvhjohBx7
IC1nBmJve/RfUZeZfoUO7TDxaW1zK5bdSG7auTOu/S1Lmikx+UyUMuW/lI+va5iu
kUs1hCZWVUfYz1TZULuzUusJ4v16+AUvJCBd03zCRswFZzzAuSf57k4b+nSML5bS
F13FGC/8A7ZYVOhIHYpnXKBwvvB78uKyy2+Z9jy5Ws3iiekf5f5q+8BGgZ9euQoZ
sh8fwLY80TcvUOfRzxtL5M55JChWrmwoF58YdNjLSWs708VLE9MvSoPru6jl0jt5
g6oZzzyKxJO7dFXmjZXHM/mXiTSxosCgL9OTtvPrl68a28jyVfG6v5bobqveh3Fv
pfK2SGE1ja68KlZg5OBkwyFiChD9ti03ZrX1h3+7Qz31W7rOQKR0uJWtAS+fZThp
sOpAGRI65g+sa3mu5QKwDeUFIVsorzGcrWJuS73z22WhOxWrtVdvcYlgbxFBZEEq
7zR6k07TYoQm5STwMldHGMH40tGnkA34+xRe7mw3YTS4ZCdtd2rg5HcZ28O9TCTX
IP4IhuuydRr434kp7WdNhn+3vnV0AuLj51yf57HLXk+tHki9B7Z63sGUwn0oPY9w
tqRe2o32BPvLT347YsJ+bZW/0Gq4RBsNskFPDFn5XxmbFNqOwgCuYqhbXKQSsAaI
EL1Zfi/v4RvK0TSe9hZeRzYzLxSZQFLtf/NPs2RMDoOu6+J1qUiZytqJFUg7aHHD
iK6q/qrwiv3PptCoKcAaLosU650Es0OQnq6CaBL4LpK6uHDQWnrX2lOf+Z51IN4n
+N/K0XPQs3gRCjLMTiEPMmWjq257yX4hjuE5yvS4foyzq1C4aHc4uIr9mR2kyVcp
P7b0+xyPXcE3K/Todf6Q33GaL0uoEJStgpP9t/IcoLX08PNyPmbAJcHC51PxUXIN
tVU9bvl7pfoN/DrMsxc/BfUlzJFuYsbPJKEbudL6e+KI+rISWndTN3mZ2rGCJM7E
z9etLiAnEORMZX+TDDMLB0i5ykugOs+wO+Saiix8Zf7m/rd0bzilqpsy8b0cxy0F
kfLp1dUFVPy8T49dScPEHVD177KxJ5SHJ1SD0AwSJ/WY4HkOcc16JD+DZLUW096G
LxXJD0/1MTKWWZi69mKcOmwSR9PDGr3zW7xRAf5W4TczNsQjpdVX3ft63J7vY/GQ
LkhBTV13+sQDwmgTsM+7ulyiEudwyZA4h9iGL3hK+Tz7fhxxy1a76eESFI6xV2pX
Jdtd39oU2w8aqyQm9qCQxMZX11B620+JcEulDYiytZmUkfz5Ox7Iq6E/2hawWEKv
Z1F8HGUTpy63KjM39qOnc1Nsx48RFoY19dAiyEt23Vm/fEmdBecp0jTXyF1BiMEX
4EXXixaWoUbqwjgRj2ZL75TnyOiWH5QJDwkrFhUl3U+rVtbRdmBQv7YAB/6wliNE
6NLgLm3y4k9OQKTrxYKNYrDCki/WjigCEVL0yUHB4NBXm6Xvp4JQd2UE9JsrYol4
Qenr8QUMG6BCcr6MtdmpLT9nghBYA8acNj6kbt4OLD1Wlxe04WZ/N7ZHd3Jr1Qv6
xXYkpOWvradDUpdy18uWVS9mFUDvz/tVu5uBK2usm8TamFxUQ8dceZpsm1/Q6560
qMZRU19bvAkOrNcRbNvLHF/E5aHMxHE+mzHYZVDIMGj3wY1XWjOGEiCtEYkBTH+m
BLv8ibcv8hEyynRTEEGzimUPxPoS3NJLlQ4LnqQXI0O/tRRbhwCyffv5s6WJF6DM
vGSqfkJNJbIIXmFMTFWGO2F0TJSCedjjXMpUOKsHO1Re5WfFnvTntkK5T5cM3sm+
KEy3RMfZTU4sJ0FVjkyYwoqVlTjRiSpwMVrwfzuvZms4Z928AS+kK9eJLux10HSd
QeMOcZqWkipFhGK4W1nrbCjhTnEGYBPzftKQXD1I30K1de2RX85fNwZM6/+uffR2
izOZ9sV/cnq4sc+AzNzHlGqIGz/EdMBHNn12xsEAkYHF55Ry9R8gjXYRQE5v0GB+
Q9dPbwXwS2NXhkyOhxj4ROJN+yK4h0M5BUirfCvGA0xlkNSsOCm0LfZ46y3n5UlP
ilObMbw/FKyp9s642+8PMOTTFxaTgLZWu8VnyeaIklwsfRjJIXRZJ+K2CbQsS2Bp
7ZjUY6Z3b+FpBi4ApcHYbu112ZfVOG0Iy4lXSSwc1mGXLBS8Kb076dpemRGoEwUG
m/6d1lFGObm3HHE/i5YuhQVdPpiTFSHF9g0/sD+P2ACrXMm60inP1uhiv6EFbqcr
Aqc2AI4TtQiXwRR2jl1vFsotG/wneL4oxGSHT/YJBhK5qZSBXJrpx7SseUpddMa3
ZDEDh71mRCHsrKg+dE3f2vVfDK/9Plu93LkSRJkE9m0i6qgPlqtxn07PdMrWQa/x
Rba2gK0216u8wsshLHtuVlfWeOcT6X3O+2z7bkxYkiVBicBNyGAUYtXkgo+cHOjY
3vBd18pBeIwBAHnnV6mxS7o8X6XFoeollrgg+GH/Xn261QbfOc49iFDjyIIFaMGX
KIFsYJzov5q7l3pZZ7EowqO2cKMVwuGtLIc2m7ddy88vUzs8UqQBkn01m3OIYqEV
dpUw0ucyL+y6q6MWO1NrtWQB2t/T8VnSPALntQM+F402BvOLr2aGgO0RXpA2HPWf
Njmc4ju673iVAG+fraNIAOG8QTZbieI4CUSgIRrUr0no6qhdRMaEtlRRKKX/ymDI
oOxzZTfHStjVMfUi6wJ7Hw/NNOResYFv/cra1EK8Jrp3tYtFr99L+8HwIhhe3ED8
mvCojeNhWIvQEKBC0slPjyUGgL1TSiXRRy9Gqu+bT7bnbjSylrBpz8wwfL1kJ+Yu
4TJ3jxcfiRAr8jqKoH8LHBTTtHB5pceJIizDqCllkAppDN1oJzY1nrhvcW6zVENO
aztnWP4GEAfzwmyi+McRcHutpY5i7LbXdo2qljMdty5EmnKWjTsGmmVQvWShbUkI
fBfwkHKWGdxlyoINKNAn63r9NS6DPkp5yzEWmDfqMBD63Dh4SmldVjanyiTsXAtH
A0fQWktnYzcITieTCwP8//M9/+v8/gcEQ4tgyU9DQacB7QZl/YopVsbpYLaE59OM
/1C83TRhMwHTtoyoEvU8IN2XsH9Dy7vEslSgtmDIckuRkBNDykXw5IqKubLX5ecJ
lA+C+CxaZH+gcHt7nFGnKOwapVV4KJ+bhy7hgBezfbM4U5V64CdJOx/uLvrBIKFj
zxReC2vNwB/KqJ3/9yevds9AY944z6j5kJhU9v4x3I6bX167ji4u4w3powHk/I2U
GwzUr0habFX1tr8hWMaeTJ0F/l7Ycm2gZBK93Mddd4ZTHYS4wHMr7gX+2eyzqsau
T2PhlCHVR+hVNegyvMFb0OVAWswpvoI77i2n35ogQxxp36VbmVpKu/7mj+pQYmzb
qcg7kHzEbUMJ57K7qjtrzmCfC/ZTWHZyyDUamu/c7YqQfHFNjRhpZCHwrAlo3nbe
qPRufOzrrIEebP8I7bmhl4PsLe4xBHcWB5XfsBcCAsSwb8PcMIxa+O/SYO+A3aIJ
f2rzbEWipHINSXhd5AmuJEly5aK83jpsIMpgGD7H/ge1VQG0OjaNojOL37CnQ7Pk
mWaeIM6gHGvUlwEYn+tvejryxTJ0ZrizQ8uFCrmDuRE6fZOS9P2pSw15AlPt19Bm
uhmTN1jRK/a9jekQRgewR33Yg4NI4r8ic5Scor1BP7ImXgEtZ9bqd8CfHoLV/czM
sqR3l5ITq31/kgdlzvJ0KqnsIW1zQRJHZ5LQBpM+eWpwL/LIzqZa1Tw+Fj/bEZaH
IV5YpjUqj/lupVxzWAEV/IozBYHmxAy2fobbjgiaBpW/RoCGwIXvyP1hK3cpfxbH
7P0xiC6cJ9dvJIfbFZ94UprwKxrur4YMusO1f09Jpxxv1kq5Ta318N90Kxxn1EBJ
78hQ+95bXApte9+/RiO8f62mETZ18F0Q+x4QIva4cdHPXHORdLKlu88gnt9ayGlO
2ABSFbDTRaOhwXMVEtgxyjrVnh50gFBttUNHQuo9Qi6aaSEn6i6sAtH8/WNlo3K8
slqAcb4BTEjH7miKJ3QmPack/LPCWoRTtjVTjCYKevFd+xsKYpoNXEUPQiY5TeFr
fZ2MtiV6lgERczHkDB6588ILeS+5aJC+u41qIi8jaVT/jC8lfXUVkKq60brywK8/
w2o4KFWBVOUoRH7nRt/U9onYR+MElfQKTmaiKhNT3B1xWVdNTRy4EGf10kO9xumb
Hj71DJBbKpgKC01sU6CSB4bATmGY2fCwJqbTXUflWfbDc6tTlVOTVp/rEuvS5fSZ
okYZ8wNxD1/y0bMVMdvUOVn59jzoFz8qET2Sdfc1AzpQ7SGkfF0LsJuRBrUv+7kj
BmWc8U1NrCgU4VWtsRrJFw2M8Br3CarI/FAlXPMaqcHHQBhjOTCdd0D6qHoXLPC9
M8UmXlV4JsTbPOvl2c1I4E6HL+7QO6qG7a2cjw5AbJfva+nwyYHP09FYAt/3dlPj
C21sY4lQzSsRMd30oegkA3KMM8MdqZxpXU27X9hrI+BXYMLv/VTJnel1eJ+2ZsuQ
dhOZ7aFkBWsdcpRQ8Cybca8HLEZ8GfnD63hnKxgHPY5/BePEiVeX/rimRCaRUXLy
DcTh+D/u5vQGcm/HNMQexrZSW9Hpr6CM5m5cqJh/syczZRp0lc/zejEbPUdiNQu4
hh+sCZmqVAway1H+BcyjPDOKNvEAQ7JtQmEBvQn5EnmE5wo2CM020QGIMPYG0T/S
rv4MJxUOQvbhlZhZpAnNASKnrE7WsRvfwESHV1R86I8EWS2s6eU1Z/+lmMqjb402
PYmQ8tpiGgDPK+3lan6/Iz8lbtvI3lwWsijZCWnzd973H6UZ0wnWzBuowYLFihWA
X7LokunLY7MQsz8M058BctkVI/o7yzmMW1+wbGVKz6PYNm0XK7W/eJA0YI9wRAoa
K8m2SlzRtHmrR5vyRHi3L6MLP4ORaxc8z8whFgilKkUTbxUjSMQeeO33UO7h9PCo
5Iwt0tBD7wEs7TU/KAFwCk2xcJQJGXeFKKC7F5zWFu59TlEDoq4205/NS1jgYROY
X9y58hGjQz3Z7xMZlodswPlbh+kiHFqDSohtXPmgtvisKUI+6ec3Tnq//AmJC+4h
kK/xj5bxulSwVzn0qrrV36+AdCjF5M3NgDglFf8sZegA9/moagioYag7B747SopJ
eXlv7UgEbYFs5M71x5Q36y3Y0ql56cPWMswLmp6z0iE/wAuHJe3j+qb1SU/YzPGR
FhalplE2xPZsZJWag2hc8aLROwpNFFX391oZbRd71xnLoYHo9LtqI3yRVMDCuago
EA1JvNJm22pU5YUBu+d6zI9dt2pSMy42d7RIBQroH8TCF8A5iR/6nRXZtHIvDTqv
0UPuqKi2Gz4jJ8s+Vu/f6CDv34GjibsCaR0EZHcTI2HJK02e6rrM2vRzmzFoMKHy
FO8liJ92t3MaEnCnAAk+vELlDfcrzebSCDQlJIqa4atLwVXQohPLsfrE3oBI4yf0
/2e2iT/3OwH4lVudXhEehcTxlIDFNCO4sOR+InVINDTQdFdCegEtq5gN/qeR93bD
ma24Szda0UCCDcNQ2+O94Bt2+bepbMtq/wNJXA2QRweQI1D1hD7QBATSlQMMwPPX
QR6RFGG9CUZgsk/nYC4fbbddjCtvF0V0mz4+/0hYtjiuSdApPRr0nPpJzoEDNeV6
MYs2Fijz1UsVOzBOSrXO1q3Xg87gAVI7TYjmoju6RJ1vLY4py/9HEsApW6NWKIid
wKR8R31Y6+jn900d+YodZpR5gfs49Y1Klx5TiCJ2ALLzk4/M1YoZ5JNM1qe/a6rn
RWZGABvPwf1QgwjW+DpoUAJ2HTukuUg3Fxp4S9Jj14FsRyHp65baMcl/r/muuv3U
AvUwIf9kBhgBXn7jUt/pYM1aA+SP5YkJRFOPpO+VUnX3TRWpAxSiobcwMQpCBQPV
nwouml3F6sQLV0FLBV01FU7+Ux8VKWD8mSK1+tTEK+ZGWY2/Ewo5qxq3XzN2XMFI
1dmzyHs0ZLGhtBmz4gVHFKgtbH12UrbHIFmH3ume+0j7f4Cpuv/UhdJSFWhlIUcQ
qfggfoOVzutbplZOWTTEAccmCFBFT4dIx+k2scchwtuOefix7wAeb3dvKm/CNY1y
ICxtnTpTKT75Av73zi1EDryjCdLkb8QhMzXJmaUCY7+EQjMxkzvzc8pTboDeeo5w
yPyyxofOB2g7fzw7LZ4r0bNc7pqtpL8AaJ8rPA5MQKDJaka0Ln6fRCxe7tvHnfVA
4EHdKdf5i3ePXJyoXa3vb+68OcVMYMeG8SXKReupH32X3NXd5+76G8vQIz1x7GlZ
qlTDfRyCJYMP8TaRrZNcGBlyn1zmD1+9eAlPNrV9zyxD7VQvno76G+sBeWVo7NdF
OiCgBIbC0c0+2rhDLPXeUClxCNa0cujaBif44lz4/7bTMZiUDyzMOkPE54biOJWJ
MVqu4dG5Gyi8FqklR61beQA83jHcYqDHFVaTtFRAzgGmLRICrzb4HVTEaSBpeVDN
pcR4eZwp3gTjg0MSqDogeBZPAN7TGlLqQGoXc/+GBf5I1J9vy64ef5Ls2415FKFk
L2kFD3NrnFiqXr4j8NHILrW/CLMYIX9NX0VXuiX9yYCuVqzjhJ/c7vIzraUq9smM
sirFcz2i9Ihb6wyvjmEFEerLuDZwZeqv7/mv0V5DvFZ8v9HznLkZUzaVhDrC5G15
2+mYvDZDuyD0UxBlNeFSeKLkHNByBV4G87kRr+ew80APB0IHGJE91+yvACcJk9xt
HvON1sElh0pr5ptqe16hLAvxQ8OSwYz0SALIMVjN9/J2HuDVZbsy9WIWYU52Iy8O
sG+d7m+Nr4TIGYtvLWVatPU9WJab8E1EHnJCXjh1BmHuFMpZdOE3vk5NMfvNG0hy
V1QAi+qRO5dzTSUxGWRbzRvVW1sQYaP7yQCgNh03km68VPoKMOa8VTL2+3gJLjzC
OXUjJb6nJY99ZtVVrqWdUlXlGLaNvPVkU31sn7dwi5eNYbpN+J6rlJc7xEhiabiF
Ux0cX26D5RXtEYga24P8kpuSsUeOA4BvtuHh5OyeUF66nLirg2EHj9mcme21WhDW
AaRcyeD9NgZBXqr3uKNXXUnadFlexXgj146N7KPtqlhdPug2EK/MZI9PjJ6epJdt
UwGH/BQnVQMfcXNvakAwk2hPscjrdXbotLOQX+wKgWg2S2oR4jalyACZaq2SAMpV
eUczYUdwZ8sK9p99C06XXbM1GHJ1R6eBGdOAjn36ExP2uHDWnW0ypF5nqAVjfJNQ
FUMWK3MtHEIow8zEpblb2IP1BYcLUWzG8xq3V4zwgBmmPnDI7bkJdlOqNMXRf/Kz
3zWUAojOwrMQCXAVpUGBHoOxhTqrKz/w4buyUKDOzdrUbmMviGeonXvstslXCwA+
5AQaeo37JPeaMu9yd9NpRsVjL0VDkQAcjAgcpwHWl92Sw5wejKM7dLHtiESZGnxD
IeZCleb6EdaVhSKO7mlmCahJ1oyAHuuIlXRI6C4YxAhHnIrAq26g4CTZ+B4EuFZx
vYQCdeUmhJY/vEC7ie5jLgtG7YwXDKnXCuRXNySzBec1kw9aBO7NbwgelnRRhlSx
TaTzmyRY++/buKJFqjApmJRbWKzkPnnTU9BDTZG7OqTTxZ8nkwwaK1ki5B0e/A+R
yOUCi8xDaBLFi3wwkwWFDEyj/c/UNqn9DRYFDONDLjUm62b9s1gHGU7s0/w2HQS2
ixxXRiyZMEKt4YxuQG39I2XkRUFgcYCEou3So4WHcyPW2c4LMxlE3zQiSsad4Qyc
JZBzgeNzlcakqbGvT6IW3x9WXoT686YMKbFJe3G+GR0TItPz1LbZ2YVEWa4pXHkB
V7uZLsnSOlfDY66VtLu0ZBVzfA7J+xpIZOY1Ufb5vM2k2uvUAIiMaov7IkSsGwpA
YK7hWvwxjniQxXk60ecaoF7dYnOx9Mw7yVN7AdYMgxkmq+P38+sHZ8JHAXNFXu93
u7qM0KSDclR/AfnqfAdu7j6+LCgstwyYVX3ge2/4FOdBcuUXNxxxl84/q4iWTHda
kCoF8CujcgK7a9vrymBotFBhUGtLNZvGVX+7QMORq3HQv6i9u3lC3EE2GmxXsHym
ofrItA7kEoJKd5c/hG7iyV1sBX22VJQV0yOIR0O/F1dQOrQhZ3pBsw782icrERqP
ugZ1xFsW2knbyvKWcHAsMiYlOFxXVhVlEt4a5GHpOTS+mH/n4usm1MxAQ3WQftsT
vQk7YQbBFi+GL0aRbYpD3SWRPZZ/RVu+ctHZ2nCQnhq1PhFw6pHSettXj4GxHSDV
nL/HUqkQNCjm4PYAOafCHZDeu5a1PxIe9EVCIfgZQedwPF26RgVaExCxkwQVB4P3
5e7NZKZq4HaO3CFHSx4rar3TH7FTjHMTtZzE767tSnKYCB0SFwFKn/eSfiQbvQha
LUtBpvH1PoPnmoT1eh5Ld2er+K24anGD3nNxVpU0XoGURs3Qen/DAFRnp4xG9pZQ
OsZocMF5EY020PBu6ICFHMvikcGW0x/cWD65jIkHInGrZwsCQdn30ghAv8GSiA2u
LdyNxxtZW+rZxvSK4EVj1yQRidGoLSLZSxs2t8s9Dc7FdZTd2y2Cy4WhR+Eq9toE
Hef9OD2w9yNv9sjkYjWf3Z/yh0PCMJl9EThjTLZ0qJ5KOsATIe0VTUkVrLCEygbL
Vnt6pq+HHK/YwE7uynnRtizJkJq/Cvn04nkntUb9ZG5XSSNziMs9npx/lN9rPxt8
f6G3E/Tvq8hRZtcVOgJgnhZLPNrV02xW6HEsXIWTdb8WmJihryKPJacDcBuxZHgi
1PMUUYl3gp25uS7fdIbGbZsduts9lftRS4jDAG/3+Hqn3h97NgttrUb4KbMUWQQ5
0vYxRNK9E4goH/BjpV0DkkGgbOblLmAQqFt6uF7f5z0exuuSEfkMOegmD+kXU/2E
oouwjDDXxxh4ar1Qi5EtmAjqLS5tbqpdXB+kKrTUmnjBYdQY+JwzJZvqOeCzONhL
oOAgJMyi0CQnebgJC18XqyuT2K7gM7SfztfjeP9nnTOh+EWAktUqfY6Cn/GmWy01
PIoZQTsEMzxM0E9f3v3Ua6XDgkeqVYIHwNW4D0r/h+v0RdsU/D74hp5XLFYpcHF1
HWM5cg3mEKuCpLgs0/fpPBfd6KojTYMiSgAVwwzenq9+iItVRlGIRFXYV+tS2+MJ
BuwMBsPQ0JiMrdU/JNfLTSZIPaEZu99zHZ85CgIisJvWlGfJNDJOrv4R/qj4hTQb
pro1KwRR7WCj2C/EVtsnPc6r2EvXDynetvtnzvgvg5QzfAol9ex6Z9jx+Q69vC1J
kSsDW307++t1LPLUcBQ3/sW5fXvLk1DQxmpyksoEkOnepPCfdD04jiWfjYkpvWvO
+RUduL1FxAptH98hdeqAq8ee2RqVL6VQfk3TeKak7vjWbBLVAZRrFSsattndbwvk
7cN73DUyr1GXn1HlhAUrHtq3H3+Mt7fop/LwDti/Z+TW5L/oaFswFNX0XT9FBR5v
HZQ50I0XEAjRoL4zonZgwT8csYrx2CHQgW3Qwf+aVIOuLGgWMgLMvoqNvagwv1hB
4HFSYnjLkTalYcNiDdm47tNQEXQvmDjIBr3JPBPR6J0xI9OKgsyyZTkK3C+XijEB
aqCR+yDL1+kzxirOYMe5aR/tPno9R+ymn9pHbAXt2prnMiBAwZjigdQHO3AFZPbe
baqQypjTZXRPkWyMsSJL0RwXMl0g2cgcrBmOjAMXULOCumxTNo0CbtI40y3bOd7w
Ci3gqTUmUJqiTgBaHy5IMJTL85uF4ahAKFNnu5QZFJvYL2TIpf7NYsnDM4zsQFmk
unpWUxt1smChJ882EyqNDkX5t4PN6a34YLXpWJWYW5QVJp0MyB4dH86cWaDR2Pfz
/QRyc994dh/yXnXxMWNCe4/b7bOucIvLbfgKdxoQ9fjw/BgsikokZyP1aSzEw/4v
TcRktGH/n1AA881KrPhiFwwOJ3oufMVXhHPUc691FJ0yUrgXMoZnFf/xA53tyUUq
x4VBH1g61cRKGJUJtjkONPwbYHLs8kvGh8IY4xdqskn9KuUNhxQeOrSrr+8tD67D
F0HBNyTJpy3W4d8h6lj/bjoNIUJ5JuzYy/VK0pRRpVf8AM8l6fgbplm7UAilAjJG
9X/sM9azqlOCtfV6CuDZUGOfDdGdfHbsCr/oxKsa0jnTDzqSw1V5163AYxVUFRN5
0TIxVvsexN4V182VuWJzW0VQ13MAxXUxYzpUB6Z8u4eYpF6XJRd7YuEjKY+UqgDR
m2lVxBdOzZq5RCHsxt4MPa8acNdXmIcD1H7jG9hmxKgatL3UxKQCW5NqDPPrsAvp
da5uAu3k+zKM4CjyHxdXhkOvyJO+TYOjalwifzJAcEw0/FHMoqqTQmmima8Mpros
Uc7ip5m8kHUFP7dknSpp9BLiF5wyAFzulqeTW6WuoH3KoZ1pjxYFInl2xXzC60ov
ozVkOMCHz1D/AFaFao2k4AZyh9SPU1Y12kWaqXJwZ/wCW1BkZenfi+FEGv0FJO/i
uKkf4Bs6hE8OFHlSrFnswob/FRzk16/PJvFAm670XAb2KeyR1MZyQYRbWmTmUbU5
HihCwpIJBV0UKvi+MhBecsNQZLTNbkmfvcMh0Dg4JGxfSwGc7xssnl0aHW8iM4uO
G/36+IsTElcjz0T0PvuH7GTVlTFvpJlEBjtVbhPgVQ1/uvPxuEXxZQzoQrlizYKk
so4iuFWyAruLF7Y1eAHYKXexEVH7sRC677OIso0hQC14D5UHX4Y2gYogeYgoP2oU
0FTCz8rB68qr65AiVxiovQ6cq18hwivyLbfVxQX23N7G530iBzy7NPvDmMcGfxWZ
CWobVV5Q1ZoxVrJ28Igr2urUFiyvtFrT2ry4ZunJmIb6Putq8kfKAMpsYy4y7EDb
mq0N0xzja7aWDKD2IOHNdNrH6/sf/z4D/jOM4vNttHsepeRi/p5MjeD4Pq960urt
xQAd3C7GrB8WqiB/d1eIiguKkmWUa7oiLD77Gnvww2sx09s4Bwb3b7s5k6EB18cW
A/qA0fwPxlD/nWRFHMb5j8S8HZ8aSlnGpaZJ9PE0LPJRzgXVF8ya2VT9PAKM2efM
UJSzM1kEdtbBpMS+gTd3RJAulv0IVmyqqCI4QT5sNMseV+KgHBaOPu6OOtCnFpBC
wpBMYan7+73H58NEUQnPHMuGPUZfpV1cS5xLtwgADH4Gvp6J3bnJzG/Zc/1kNcvE
8lw+hqP/bJu2dsBmmcqm5ko7PofweZ0RA3fnuIorQal/BnqarpqM6Wqd6mP2teqU
Rvlmp1o7O867UrT2bSqi5uB7JowgsF4EpUw6lb6BYvrXMUSRTFZkO7B7V2A04UGh
vsclUzQyThJeHMMIr2xJPXBjHJCKybm9PVkiHVvKaPvzxhtnjez7kq16K3J/mK86
RmjUfCsAu/H0navt8MT0o2NJHXklwRYZDZJwO70bn0rqb3Ke/71e4YPrweEC5JSh
SK14P8Hscyy+3y2Uh71qQ5Ia5vhNiW27EeEucE8Saa2hLph0Cc14oqDJ7pRkJmC7
gIr1wahILOBKL3hC3NEajA9HmqTqXZ1Scx+N2VWyjO4GO//qWL5Ryju/Qe84kBJP
r3FnBDAnrK/dlzcID0E1GvGipeaW5mXUsDvl48usqB48CAmox1JP1ce2c7ZrCFf+
qUeAILEF9qbUeU9m09tbVdNtnPsJ9GCU6mN1BgnuNP9OFXZYlxYyil/AlRjChqHY
UfFZbjzdeZHdPdcQkMQZcWNJojgrCvaIHqELAm/2Jxbsg6Vq8OupYu1zFerNXpSi
iDoCjWhRNeLYI0e9QeAmbfJl8ZP5K374NQ3wyd3qlTrQlep0emrKwhoN2XFlj+bj
sjWY/Ijd2Y9e4AxFHMTF2OS5z1kk8djyKU3TsWzHgJbekXT86liDEnE5pFAenxGZ
Sl1ZtO4ioalVGDixVVEhU714p4a2MqS8jQmFXmjS3TqJ3vUT4eYfHw7gtCfuaIaF
i8vP3FYUR0Sd1mB7P4ab9GJb0ndYTQqiXLBgH3KSUNkHpyhnX8NGoqhnSdDrOUM/
F2cBoqybGgU2OYwKIlEpZu//dKzK6XGNSXWMbxL/FIonU51mmgZ0pRznIBowepCG
eYQ53B3OZc7bOgbekQDC9F/qfMsbyz54sr4piATlfCFO0RztHshExrXBea38tsNE
gHJhlMyDIlPjUwb+elXKxxi+hHQDH3rfDV8NdiWYtjHe5EGZ0mIhcjwFOl6DkCRc
ElRWQWug1Ho/B4unxi+SNGNwNDWOpJmDFsxmVBfcbd3DdRnMUGOnvNBVZaTuorMf
eegTtykIDexq7nXGSl8C/aZrRHOC/6oTpAKFRp3WP/s2IYn9PJUF7fjqUIYoubGP
QUaFFqVZNXULq+9rbhv9VCcyhkHx9Ec959ZEUCfdGh7hdi1Vvuyn43ux+ORgAzSm
Dm0C35U7mBAgCqGdFBbI5jigl8rOFP9vdHxXjSyNEC/vow/zPOwfJt3YUZips+ei
LF/to4Pf/+hWIsn8GQpk/rDBPx7s3jEc5VRlkPk+8xv+zJ4YFcuCYU1AQKs1+vli
gINYSA6cUzvFCxYeNsa90pbsOTPJVtzZ9fe/g532h7eeQrGe9mDmnS+YQ1f4vdWp
jFZoellGu1HT/uWmYrDRAdr+aXGQX+I3i1YRSM9Nmd9x+pWeJFjwpTBvXBASlEv+
9Cuiol+13Dhxj1x9/Qng/NQdS9wYNP9r09sb18N+KAvCzc7LV0BBH0k5MmsLXaLc
ZiPtbuK/SjQ/F8WTTK9u5qBzzqzzlDVqYRYi0HYHJxkLppy+NCOTauDVrwktIxnE
rU9f2YmOeLtMdxhLQhUnblvJlnMrbJJzJ3t/Rbt0f4dLDx8gTpO8wREZkGMHgJyB
hixiX94ich/4UD876KkxXMsoOhf0Ue2Pu0wYqpMkN7y43/4SehIPUNKy3rTfUiL+
joCGort5kMh49TBMK6b5OjIRQhA7lT6RgAWRSZTSJXFiI/VaLUZzumecz11JMlAc
VNFBRo0wf/Z2WWEzJ6ngB5Ga/F6AAYg5YkyR5GT8VIUgmDFmoW7TRAn8RDtysKCd
kZdQGqHpDJtmjClQGmqn8DbsnQTDJKqe0NRD7LgKhtak7Zr5jBzSs0xFGyOWJ1od
vUxr2VcXbVAeBtb00AsmbfWvW5IN1QkSF3MfkpH44ViyVwMzQNVN9lzkfCIGhKs/
3LcrQOhjcdEmvLsW1T/D5/WYukNffr9caWYFlm54gdiEE7Rcm9MVAdpq4N/OK31a
OJ3+XZRqIyk/ej0RdZaxQ30nxq7ReWVkxao30G36zrxyM27AmVvwxEJ7o3+Q0HWt
+UdUE2rK5dCMNEEhF6nmdwjyR2SI+1hkg8NCz7QgrBnmnGIBf+Upp3yDlV5nsgRp
5WKZHwdkK75Av5W6Oy4ga187wwry3vr1UzAY5ihIOIXkHXoEV0+slPwr7eaKRW+L
6mqoABsne9qqftr822yziWMfgKSXoyYI1T3ZsQDND+RAoBChlnBP3/GZWXTYjemb
IDigBMeq9jO6AQxVbFyNPb6QMoT0NIqUxTSr22PPs2zABAFKEmCprCdk73/ogXO1
8kOmwlQ63eVBZhFsyk2+/Mstx8pqa2b3RVa0rzY2ksQV+tIB+m39czC0f9ze0PR3
Dyuy68Df7VzMXroMrwtA4kmhljOYRd36fAO006jjaA8Da2neYTNPlevRE8JgFrjH
X92DQVL/bQON4FGmOT1LexhM+0qvQUS3qxpd99lU3M3CqAPWrwFFMxILz1/XwILH
a0livcKTd2aCFL15vR0asmnVvWS1zC7Sj5CE64570MNOocipf9Te0b45LD+LiLud
YuCJSc7Pcp0yYBkKeZrXRsJkfLYnARovIzu6bgi5qDj5XDvsPT/2BMLqGpsDGaDo
31XaBXSXhY1eg7Zqo2B31URxOqaeFUGPWMuRlC+D8JxM5a7ot2rOA7vbXXRkA8hu
hI5ZkBhsknaYAZknAyteNBKIwDagzfbPz3M62CNLQTwn4N5nMxX749ciDsx7+ZI6
+D8Vw8FultIw+WaStX97gYRNDqgpyPneUxpPN/ZlXLFDW5DPyr9y2xatqtU3o4P9
C0a8njvEwGk1xfewD85JE76FlAXn/OVzoBEABPglQNB7+1UTMjySUylOxUoIga3E
RELCaGVGAoHnOFGv5i2gLtgu1BqGyHfh5af8wGzd3Rvtyz+bPhsCdIM7p943wteK
KxIFrMDqg3zyQMOeS+o5MyYtADefOy4NJgov2ra23GCwOznZL5xfFFeSEfAck+ux
TrMoPEbNnbTKxUcdv2VWTCJspvIFggBFeWQNZoAql6wWyE7EN/Rl5tAo92BMZNCn
MGa/ijY9eZZT2+kcEQyz59r9v7Wr62LdNPbGjiHfPjWcQZTHvBjQxXJoAsmNgojG
xKs9rP1YTZDeQUCLW1alOlyHNP0pgYnN2ElehwMhSFUx6pIUTra9ONbX62Dy1uad
bfCSR44w6gdD2oDSOQeFxQnfXB4V1wKdm+9nTuao2kZ/UQKBiq/k2oyCPt7mhiUZ
shK1PNezwEgIrVYq6U8aPTPnGJD1NZs4ODpftdPLdfSkqP3Qyb1moTWikHfSfyFG
j8yEdkVmahBmwRXznosRAdyoZZKEI7Xt9X+bvZACYpXYopIVuv8z6ashWadLrwc9
G0hnAseEjHGEWo4MW0czXYqCqX7NaYo9HsPN0wh3f8ZsQHU3xgiEwMtUi/72pesJ
NrzCWA5c8MJOAb76ncwPeoO8YZopMc3CqKaWsQ5L9NSQbS/c8QccwmqIk8K4TF0Z
UiFJ8P9x7iPUPG+WD+wv5HsiRsyOF0ixWpEnJCRtILAhuAnKhGisbuZCyYVlFMuG
BtT2iD9v92Nfb+YLg5F8p3Ty9GD27FT0E3N9J+VGZh/JORfcRh1m/9+EheKh2HUK
d2sK3jFffTc8CNQ+Z7Hm6ZJhAGXJi+WYAF+LYiEUSReexskn41qykDKjeHAyRo64
Ny9KKdHzpEFys92inLoaODPaL+5tn0/YqnyJa+pImkrA7hSF0VxQW7K3toiSOQxT
kF8fuNIZwC+OCfnoBrrfOTQlI1NE0MVDEpvi5R1pR7GP/hZltI2JsTb9gwWfQpve
eDHi3Wjbdjt/egJJXKGvHN1P6ic/k3s9ykgfrVjXNVzLLxlLdDx2edVZJK2jA11e
+fyNtXEitU0abIvDOSXoFjk2+P5GdtuagDPCqVHLxP7tSd/lWQku0LYlV2GLlW6g
id7wIeu80S3vbIOgMQJGWdXge8Fy9kiKIe5w/PIyOFIXjM3hDqnBgY20hWIfjN5P
UMeCuVjwEilRYKGYHowkWhB2/JOyrZcl05LREipAFz5LLW4ubcKSn3Vt2foS0lud
TSN7WuYr5ZDJOMH6cEgYkXhJP4Lvbx6irbl2iB40XNs4ZLo2aSpYcOIkvkvJi+j4
fK1KrV3YaP9yauJlLJZHWiWOKZxvlZ4ox/Y1razwA77TvwjiZpawEQgCse/jinmp
AbySaj0yCdl8vW5fBp1KwUttKkLXg5glT05WG4zQGWHNonpUVl75EENsoTEMPZxA
DcPAoaMT3CkvqOcOVDYd0LQEATJzyX1PxPqZAL7+HPvaOfHuJqIWdb1gLnEiypG1
fjAGi9xMaT6F8CaVY6QnsUOZrCaThtcsHOUPEGp8lpYSdVKi7+GNhxSwidh5FYfn
axi3urI9cbKbrqUuelQ//Kr+I1wSESIp9CdreQPQ6e92c+pFbm3wS//cxfUfRRMd
Md6qTUP/zQX5TJR1nOB6AUHYLR4eA3Zs1R6c7ZDOM9WIzFHXJhzXsbTnavVmZIsB
f+uqRs2VLG9CoGCHaj1HYsyF1M/cTeYbq0/PY+DqGft2ewYrUFLimz9srh3gT/aq
85GQUzkljAv4LgInXZs64HWve6IxNCV5z85mSmJ+l6KOJYSQq5wwUGwv8Dab6yEk
jwCy/ICctfHfObySlOTShP8N8mFOag+MthmF/7X1IxjUCjLvU46G8YfzTYxEuJsy
2+g0dy+6mWIcCfAMngcKji/s6t+xcAURcpskJqNYdD2+5s7oD/xo/MksYn5z/Dgt
V7AOqyZpL4U8CWNfaMwtj0NL5zjTkMRknz9oBikdIre4aN1MTgaVq2YZdy0jtcI7
nMMjRaP9QjHqrFWojKw7CUdBPagNERI2mhED3emOmlt9DEnNGOREujCYszJNl0SV
LDxTa9oOgj+LWULfS+rNCB0uweziIuRoLrx7H9Mp6wLIBb9SCUKpo0xr9Q8zQuAv
j9P6IcdjWDP7ErUgqbzj196Fde4vsiP0pbBBogEcC4r5Vbb6DYKsVeJ9nch59JGA
u6T+h2XjWCquZGG0aR5B+/YJHHkXOMXYNpEaMDRZLTfMPD+mJp7JEaKdSZeyyKDK
3GuAXZXY7vFBxrcvYucY26VFQE2EpmkFCuNH5+ZAPfKkxy6/pt4ZFkb8chue/VDr
Vlf3vnL3XQO9eDjhyfvYQt72ybvS0kMwvC8mzowZyrMN8pehX3PUE1VDfs2vzkBN
OFpOoeW05Sr+0pzS+VZVfx2gauH6e4HM/J1dGS1slH/dAOVADUbcIyf1+WV/NDc8
d9KkcIixGydnhnqlmGPyLci93sr58Rkpc+gAMuCd+OEFBkwmfNQvb7o3/srOoy2q
gjy9f4YYysHzeF351/xz0CHsGNdDgWMJnTi9Gthpc2i5EvdyH31+16HMudpMVvqi
mPaJIzRt9dVk92AELda5RiZw3NusCYnJ6YdfOj6U/vMUI5LX/QvIIkO3K8A4xhjH
wZOAvwmy5nSYsPrSb4QeHpNtMik/YaxzjUC+6asSDMZ2CMsjkVc4vy6fDomIMlT+
wW7+vYgmCb2MORslduBAzWivbiCDHVvWFz/j5OjmdoS16mxCVm6qsKpC4ctIsP7Z
6Z7oFfzVbhUpUIW+00l4GwpWu8azeoQzNg1aUpsv//Oo2wAUjKjWEqB5el8tY3lj
NyQLhObin6stax+92XT0VukTk+Tem2z9sam0u0plyjBwcFgvGTx21DYhAKXHlwX1
gMq7hXgM4mwlgLzUUCktVwtB10k2ZjlCNI6ctzwT1r/ppuoE5zqW77rRnFoQ5rD8
Es6awJKF2GjKFuvrHkMeO8uGReZXKZrkymrlsZI9LWUA5oqkqcivZ5lRtZPGr4so
IPwxQZkBt6YBTxsnvUBvg78Jq1V+RX3pRgqd+mz3GVZnGSxAP5m7KKF+Qc9+9K+d
tIgO6aHFhGNxYx9RAG2dNsaPRTEsU2/hK3bFG2uHcbuhlsOq6CKIEXabqATwatW8
7w+/+Pbz8cT33PdnF29/IT4PGN8WRc2f1AjY/jNPDaWd54kQlNndE35b9Uekd5gW
+MM66G9tCMC4umfG/rbXvcm6VQEa0+Y0+sdNW2Hfnwa+hCXLbH7g+NPU9FuahBD5
rhK/IsVqV9OhG4M161lgYkunpb7F0cvdhyitdSS666CiNvoP3I0RBZ+kKLnhahTF
BMC9JYGMVc5rxIQIXFX3w9AOApz4fwJIXeJz86dtAWc89C5f9+wgfrJGBvyXtisW
ziHirGowGx0VtmQ9l6dfBAEhbqrJlNFVxWLj4f8Q0oZHVMX0Lc7wFVVWduXAcT2i
kJrWejMNofawEoX1x20ft/3qzNg6dfDPxBZ3Fukr28k3IeyuyvxgR9RumMja77/M
IuwK1dGjZ9oJe4Pslb7WFLpwpumtAnrmTKqiDW4SM6IIu0hF5Ny05YKOlBU1qWvA
dmLxLGEbdy8x7fwMS7G65WR7o4iojbACMlh18JwYSB1abEnUckgfWbAX8AusgehZ
HafaJ0SWhGH4SttGTbHQzsNh5Mxim3tj5Xh3SyWKeRtwpKiL6fGi+sNW5F+jz7K3
ARlGoDHSJZ7pt50Xng3S10iVeZ61EZbepuZ0cvyqkrgFT5tZ9pQb5Bl2S0w+PnOW
u1W/qO9Igc3dnTdAoWPYeuGb8AHrxabq1oWLQWDaHf68XicDmkWQ0w0gb0URhK+9
TGu2/kwObbsj5r+Zpoyn2Vvg9+bC4SDYaYluJ3lnVe42ZZEb8SXCETAHjCpeLJBq
1txLZais1USZOdOVDfUMfQls1r6GIzYfRBznVNvBVNXyJcLMJ6rpdBLhGcdl4jGU
cBmF5wfbnn2LrNnqrzjy0dCuZJqfISXchEMhGiuvnLYt10VIx0cj1F53NxDtTO+6
fG0wjstuFiAr51B9O+5jUHkmK8JoIW01sXG10dvh+/53QOjsRMmkvj+5aPHwEbVG
4zE9NtrF80cYMnImsnR5Slp7MchX4CMsOd/4fM+5Ge8Jay13yVJFaCX9aSjvdBjz
nbl0XRb+9cPOdjRQUtGKj6rQBZzbh/hEftRXhikwHdqSaX6Qd5mrN8zlVrNPOASX
jhfqQqp0JBi37RTbcztyDZxmKZbOmkEeyIxfDG0Wf8YeNIrTyKeD+iCs7+eq2Lo+
BOCIIQBC8qNUMmNGFbGeE7ttpphxMfl3KWm08N1/GqSQt8EHCpkhK0Pkenv+sxRR
kp9/MPt3oxN20HGjZFtiRP+PJ86Q1ssSW05iRgKn9HRz1D28zusOanu+qA/Th2fJ
I495+8jT4nS0/vhMoqCRq3olkq/nfP9FlOzO82C2SaHrzQ3JS90Cso344hKk/Ymq
dNHd5Jwjzy15BDGtcBOxa+V9l8+cma1VMXFEHvsey+MD3w4RqO+0SL03+ld1BB9d
2pxwbrkGNTB+0sWQJpmEzIAvnQq6V4Dvtxs5Buw8Ws/WFHIl3ZBQj4C+tHw9YQvh
xoqIaJ/FUFslBmFb9X1coVjWnfVJ9QstsadUBjA3ODyMl0rEkQCAI4OKd+6ZRmLQ
fL21y0Kci82S0tAKGkSf61/Xx95+ICPhHWCj2DAzf/I6s9IwzFrnG+Z0jXrL+p/g
AWeKUTVWGpxbGF2vlEbyg5Y7G9NAk3cItm1jT1J5CGJCPOMWwkMz6kfoglbTxXpF
JCjMCxiIi/hDlDCMMrb4mUrrIfAB0tdZNRVcIvtkaGbmktdgLMAsy+VzUH3ImpTx
JWwS0ldQf83LlKT5Fin4SghG3/gUGOSB/rn527JlnO8F5BSbthl8g835iwuRsu4i
g34NpNlmNvabls9V2VxyFfSZN7hJ//N5wLlmcJzTnziQGGK1zy0MTO7nQJ+dQNuw
0Ujdr4FYDB7Nq/AJcSVmBtJQXW7RFhChKAaqDeoV355eanEjy4c8zRvEikcyeZQW
wlcZHkAm0ukakBlZxgqpxIf+vU2i1ypus13i5el7N+2ezK31mZcyCXSHTqmwzC5Q
qFZS23Xo5nU+jndi3f+95N9KCrYOjZdwYuiaEu24Gyd3NLQUmXM5QPcs+TbspUyt
bfEg/VvHQzkqhdTc7mvwOzUi53AoRNcSQTmmeq8H4ZEmIwTtLz4WcUh5guQ2j8vr
Agsak7cTuuC09iaQbpO6sJo+vcBrPOgglTIykeb1a7N1pLz2OYNnaUE71rpYAKr5
u83hss6FWfEBoquEzbPSSIkziH8sfkgfgdyCt7vHCUBaAOTT3D5XbtNLm/J/Suv+
QGJqaWNFcG1qfVPAYtcEhPAtqxrnE7TI48Y3Jmk6J9D7C6V6T8s6b3ATfOMsIEd+
XOM9Rl9o5Lbcgea4RvW4vxVJQHRSmeNgvhsJsrbpcFrq+zwB5MNgwGL9MBSGWHAX
HppoXrh1Q7eg69+U8wgrWaqSL/bO6q4iS3NOr5Gf1Lqv2yOCMXoC1cmCPIo/6VtC
KUjNROnPNMhn+TjH1uv12FSoggnrnufXdeg806Au0wKrPDeOpsB0vWlxMtTjzi8V
RU5T5O8qbo4/MQB+GZwW2L89d0sns1iBUcmtYn6+rZBAA81ry4/x+s76gMF6HeMi
asKVQWh/sof5nCQbT0FW6rcX/g3UQiPgQxYdsMAC2tnVKThnZA6zO7dDhx/yWudj
yz4Aeccu2JSrNBjJMgAUuCKvgRzCoRTWWsAr9PaHg+ZxpwCWOTcOIgUZoQ865ZPb
KYgQES2apnB67eJw7akBSY45+VkDQlF2TcgLTU2aDhnjgo11SZKEA0/ec0yETaex
WGQ9dBl43qqgQarL33V4gYU6u1DoVhyG1AeiPyOSK3l+BG01Kfg47LVulyZNvk71
6F2vVRnyPO81MYVDEsxwcPVbmeDpR1xGnVtiiEHVCCEwNiwyume98XKcEDu+F6zW
aeej8yiJUr+PQL1hvyzyJZURh7JVLL95rd0lcpkspRj7BS5DelnV5wcFlNx2VXxC
Bji427SopDpgn/FqwITt5vfhwh9NQC5558krduTkGGiK4XrByj6GnaEYaYXoZA9V
RDuNDTunYIKaz0FLtl0ewM5xiKNCxY50tOVWF5oEpJC4MhoEqeXMLNDz3C6sazkj
OUu6CHIQ84Sc4BRn74fB1H/Of5ok22cLqRZvkGOv6WVGe8mplgPT3wwwwfUVkGkQ
JGcjz0g6YcB5bIZt20JDSk+kOhebgFFUEa7coEntetHfda2M/Q3BjMYcleUqWplg
1roL1ulN+p10JNyIoQRI0Fu+h5XzktmC+nukNRsCRthyXxbGXj5I0dp7GHZHLn8g
G4kq0FtcI3ylrkZquNUg3naGuNyPr2vRtII2sjXcamPdf9zjp8UXu6YnVOJEWigX
AR32oMelsiyHgzVyzabQHckAVkMzqQgc1oNu66fvgDY6V5iYFlNg6kFMRLDnO3HK
wfzNwfUX2UXs8R35kqPc+Hd7WBnpbnN5SKorxSVOUaslicbyeqXQz/LPkhJokiCT
e+WaNjmY8mkivbBw9vJsNmGzrQr3kP9xmi/zv61YWega4qArn+kFggYR0G5BHfr/
b/bubbz6wjYWBGPNcuHRSW/cweejFYtCUpq01rXlnZjnVhQqrQ/k2B1nausIEbay
MuliPz8P2f/7NZ1pRln0rBfUhH3EvYhLQRkEbPcl3kr+aDXyMaI2+pOt58H1CvUO
FIcVYe756Jg8xb5nuE1arVu5sO7/vvCL9KY23xmEtmgF/lHpsdAE8VeS7wDh176U
KnoNRsFtXnZEuli/AH5w0sH5XAg8974xbtA784nzHPQ5U/ySirXY7OB/NfBxwVO9
T0j7iT1iWEP1sw9huZO5gf8o1B/1jaEmZfOzW0n95zR6McqQYwXkDLznhu1Q6LRa
BF+89sE3QaJJjMo3U+eAufDIZXYBHyKELUINygQetgDd/YqF70SF6AQOSRf0a7sj
OCLlGlijMR/fX0Nc0T1vop6hTraSnQUI1tnChqI+oXzaH5r4N3BejrmoPrcZN0Qh
RaioKuJVMMiEKrdYIvxOcDKwSC8ZL40mWcp2pbi3l7iZ/i1615q9AjMjb7u25tls
4aH2IrteVVGM22behvy88j/jUBcVGSt+nmiZJlr8bzhAN7JF/8eCLwo+0TTRBUaH
t2axlHsTkg+RSGQYGEDuImmQ8xk3968U/nOEQrAyT+abQbO1TEsA4XPqqsGXfv7f
AFXkmLEXaPDRo2tgRoWvffpcIoyU7oC5Xk3x14/rrnZxuoq63452PzvMnVfdt5j1
zsMxmpAUvBR/xIwc3c95hu0iix06bt00coXlY94LGmlDBw5T70mPhivgrOVCbrKx
xkFzNIYXvikupAuUEgzN2ApIJBeByPiJMDKkiEKMrIOplVn3fbw1ykI7wL2ZRIJ6
k+p3RaQ5IOVGNeIK9AHeBTgqojxEsMDt7ltxJLxl+QW7nKmGXmDH5oZsOBJDoGif
v7t0xzrQ+R4CIBwdyVyWFGN3rh4jeRG8Fa7Bo/Ba8rEOyU6Mjxs2xniXCiC47G9M
yWIsZEPn51WGOh3PVbF9D2v4RbVDHMzXZ9jUTsKDvgALc+u6KTNb7jwqcZAJgWD/
5K99u83/ebmgGFZLZBm0Zy4tabj6/zJyM21YZPXNgRkDhI8FSpvJdKfJczD7V/pi
4+KEZxIbe9bPCypw5RvtkqI7WHPQBptroBzEwsJWQ48scrBPtQgaJtgXAxAKZmv7
BjQEsRkQyv2pfv/TQJzuI1rH+PAG3kEGuS56AniLG7IWw+BpSTYeuPzSPMw1B4se
23hpmmVx867FSw/HqV+Z+D3rcqZ8nfEzmjOGjFDEm49gj7s0wis1CdKgFrwrKPbR
iAwJRxDW1bvdXi7Q3BDILF3MUJG3HPukKj0lNtt6F1OMmipib9ASQFHrYvL2l2+A
YmbCwfAbd3bWYG2Q8HMR/MJteq3J2LLDXMHtxJ2hh3uyWyMDwxAXkDRJqrmMt0TY
aOvqvr1+JEKw+oggvJoxZ10OWpGmO9esk9kp8arlgkeJpHQQkPuyf4PCG/dMdo52
Fsn6RsUSRRUeuz5VUAx6GyqgzlHZFTx/+InX4RAl2nPmtv3Dee3LAzsM6U73nufG
sZKMJxQviS+chbk3cPn6X1HfE82nq+dK9B/hoyFpSCLO6VlJL08ifx1qgRCttKQ2
7UHvhXoDGXEC4NtV82SL+itXYjJnofxccTjWrpeoeiwLG/NKbgbp7553omOTB7DM
nCu5V4lGiLb1wVR3w84gNTl7EWZYGAmkAcSn6chupQrTxVBu/ydSOToQY1tYPE20
rJp8gjzRCCnnW7M80oUXQnRuw4yg9Ta+j2+0wa290pofG7zhiqE8gQVaXl0gWeK+
DS5Rp2aeWhnx4NtykwiFIM+ZTMwfwEpQuh3BhXenEJ6MonKw4wftOMJLX/kt30HW
Jad4E4BCitXVfAOC5ogbEeXAB6Amqk+3WTyl8vljsJmolq6suowKmPd2D05wsBTJ
SrAwErrBG4uoI6HK4NXUVmEWlQkbshXL//mJKaHeCqSGELKRZCwACUZTKw9mP8gq
MRABSqpD4PoF2h6/NIVIN4YxH4mOAB4Gj0mp4WhTBqlcQDKlbpCA7KkCmw86bcRP
07jdGJNT9e6Nbpz3XQICAXHXBGL+dfquJL4Cmg9pfz+q5+CSpz28yFrzYNM5OT4p
H/kf/O0zCLlEEGSbLY621WxZhiOaQMDMZE4nE9jCjqSaidyDB4xGCEaLY1Ch1VDh
bF2zOtGXB4Sh1gyEQUNT+chEzAsSg0fOxDDJ+6KSBHO/nxKKCvzSZwfWs1GDIBBx
ZNoCJsVDbqMvi0BDOT7fJsWFlWbV9JSmS+V8z6Id+QO81GuWNsR6Aa6K8nEw4IgM
Z5yZh93CGB3BM8X3PS1KtUz7BlrFqu3XQEWdubmpvopLzh4hLDh6Qw89VhF1I/49
ZMXW9uC8iyxt/PX5CtDK1NeejhShaTY48892Rcp4uQOJwqzvTfK12afz3QFbh5Pn
jZUDXRskTk9W03btMGNVT7861I2GrIFLvlSoWxHrTS81r6KHzz2X9CiXdu1HRW7Q
ZD5J8OQ4BQFR4yVNYZxpzIQzwaRYwGRqibGdLgPWrLIxj+FBPKj/VbnosxHsEFBY
nIm2zrOKOgkFEiyfdxdCygHazgSAXrceL/zozXV+pDz3inIFnJFNGSyPyUkWbVbS
hcLRndwtE3HO97nNOX73GYMrPnX4LMX6I7faqRYown7G47uFHmoSgVu/gwR+sZzH
zH39vAXHLEjszOt/5+znprJtbIUKjv8l4C4xtV6OnY9GronEzWHejRMEiGXRB9Tm
HECUisajaUrFN39lBl2kcE+xH3X0Lsvw0yYOHZ5MV7h9niq1rJUpE6IqYkscVn9K
kfn07k+BLE2ET7JZCV/c5tzWhFRb7ApX/2y+vIiZqv7hW1Qd9LGDqRcB/4AdqZmM
k2ywaj6DRd1vU1SjKOChWj2pCNJzyEwL6U7Wgt3pX3RjTc3Py7R0B3CEZQhazydt
PCgBIEPkhgL7jlwqNdqdmGMqU0sz2zqoHMJmHKzIAN8bmjbbX5OaiYNyWb4mJpGs
91BiTcYRc0Y39TG+MHft3PbCaKXaHjdkWd9dudxTshUjwia3lFbKZvMBxN+Kd+mD
esClZd44z0E1Du4JDFJZuyIgC8cQUqyqRtxSAhS2mu1RFQB4KL0OokGYBAmRMlvl
ecfjczQ4kCOqA5PfRJ79APPwLax6OxS7V8QIVad3JKiYNpjSzTIw+hIqORKq+rWz
bxIwgtpxt3nbBNco2tUjYRXSzEm3Rrp6SX+iTZMmEidDCjitJzOIyfDI1sOdJ+93
gjrPW7vC1m0EhcpGTADTu7mGFA54YuQgir3ydscl7+WV0h8kFCJ5t4U512fNGsm4
tBXTUqvOVRhEh2Et1vmr2TlKNM0kuzvGmDUFROKJ+zPTqUpbna25I0yjvljK96T0
5VIT4zRTONiboSYOYKPb/4u7IDNoVve9EqeL3f42K3zWedFNVLa9tFfIijtDuglv
3X3QeBFtrGIlX0P4njgXnXMOZ6dKgNoexS7EnoIxrZqNkDcyoRDPZ8FoQ/9cOMv1
J5brRPNS+TFGPl1gPBKcmBtLLdKsjvrdlDGJ2lIP0vnVbFYaRegWpZqy8yF2Zbdn
PiDfZvuLKclwvwHeZNi9cdCJ36B8BrLeMPZE5SmR22T4GebdaLJndo3D/YxnxBeg
NJ2yA3kbWQcpZiN98J7Pr7omIz/bK4g7LZTuHPduUe4DQtZ6CLzwFL7aWJf75Rc9
yMUuVSOZzVl7Bu4Bg0eBfBxBUfhGcFaXmRBYqMBn55CZiUDhkiAbQFpJcq/Vgy+6
g8dFCQF+isz7i/P+xCdH74d8tF8i159PxZ92G13VvFmDv7iTL39X8DeOxbwwLDMP
rGViEH7yalToyKpDR/jWUyOc5PEZyfiWd3xWrczZkwBNcGetTbEOlRXR18gef1OW
uliZfNcovTekGl+eN2zNNpro1hsvEbkT6Bf0FwOSJCxstXJhh5PobOHYOT9PAAlp
TEyuqbzJdXq2s80hRVI+mgUW1F/NEbXFkHO/o6M4E0E2G5ItH2xB+3ei6GgVC6xB
djirh/I+lalvcNXEf0TvGOmIZO+UiDhzt0v7pCqQeLjM0JbhpUJrySrVHPIoqRcN
n4C6cELSxguRqdvaKUcJm4CNtQg99PLYZiABZyK1n4NvW1tPmHQx6mrdv8blUh7c
IplCaXGERbbXdFWGCkponcI6DsOueNUewwiikGlAG5BZt30ROCIYIG4fwTSNjQsi
GHF/FLQ3Ju5qDLqQIPc5a/f4J7J24a7KJrL7UvgijScJ14Y7ZHkCvBc2uUwIqvYj
D7EoZjxBYJCzzH40YN0GzbK6wARcM97vJ7+fQJAxkdTISWNlKKPboVz/lXBSgAHP
E0uiNFFIAPB8v0upEY8kaeFUreMvrHu5YVbmIwMXdLi6/5e1U/4i4UQa8Jqw1CPr
9rOggmJ+XMYFvOQoJFX7jaDMC2ZwckuDCewYDiECg4BpvMFrFwMkDhv16q2DADMr
vvuPPoMLwexaK6M7Q43ZFAhIL2vu5OzHqi4l0G9tSB0W0MoJVDt2aDdDXCb/ZHMQ
dbT9eifx8jOtHxrXQhT69sexqNwMfz3ldP6jXo4UczonQlB1OO7s3OIVIQoKa74T
YM2+JSuXWUSZxZtz+G2X3Sf7vmMTX7KpRHzf3PRrZDC96H1X/tQZQmZHqW0jkhBX
COqREZ67tRjLhdlR4xO/sK6t8T67YY+KOMDLbzCMkDplSPe5dDgtM3mpg2hJ4Yqv
A4GmJEetxJFG8jzU9px+IOVPMaW3jWCcZyQvWwZ36tI+h2LNsGJtlFo+1JXbwZQn
+hKIQXXfVvwv0Yt81ECUsZwHVOiLQSMqfQbj2tAZA3Qq7V3T4FVAIbZ4T18EsMiJ
n0hEN2/5Ih4xMgfbqsa4ygDdhf8GjeT4c+2/n4TwzYDDT5Af4/A2tY+D3eNl1W4C
+7bQZPe+rZE+d3mnq1ZgSpGv8VKXYTmWcTdjLc7tMVM+lVklgO8lxW3ddsWRr8pX
vzOKdpbAyrc8NdfjW7rp0oBWWL7brT5bCLxU5ulaX7Zw4+A+V+mj4ukQLgX8faWe
1Vig4ucH5I24zhA3ksxD7NP18NOSe7+jeP7VmgFAL4kkWhooqeHSFlcpMhT7fLbG
aYEVvn4RYudGH6X9ZoSyscFTweE8vpu4RcAb7rfTLJYAmZHxtsOhAZJDBxX4pAwT
7RohBj1sJdTRf6ZzrIhH3t9jGYfzryuc2blWOyI4z+IEDH37DfBar/rmwAhaLGaV
inUNxworPRlsi9zgB0U5sG4hba9sJyirqdAts3WYkcP51xfX16JC49+0i8udZNzO
LzAEJnj4AdfQZfJ4KWhHfNCPaJqsJ+hamHsB4GpZ3cxpWXrd5HEsgdyrcgjtfO0B
ANRaT4sc5+knPAvwnZcVkNgkw4oZgmciPgPE9rLOi7b6vTTRE/wRLzujE9KgRydp
TMu94A1caBm4l98MRJIrsG3a4gnGUD3t2TnGpAfdVFacHQLgXKRZ6enHhy90O8ZC
4X6C2vn+65DiOGjxbm4Ec8NDk4IXW0KsuHwfdtU5Fxng5C8SBMP73zXBNDREP25I
T0LBNnaVS7r1qezQ4GfNx3SzsZKDee+YdoNke0UnuyCixVxNVksiSahx5ZT6e7yy
FhxsxaUzoci+s6035swif1F6yk1Cs/gsOOOUdb4eXYMDse9XLSiAzzsWt+8jcbd0
x/TGH7EoYolNeWDjE3QtEieN79kGYWDVMHYFtZsXIjLPVus5KnPy6jayUCBREZ45
kYqED77tUVOdNGuzqBZetgRpeRkIxfpVVvIUQa+mYVSfJPoAfH6VBQmk/Vj1wWdH
U2yyzWG2qOjSaAdGvF1lLGmQhr28gZgBfstITaJUbkVfnDAJyLAFNRW241qqywWc
cbYIbsRNgloR6PByYCPrq0Sss0oysbAqjDV6vwaTl43WfUn6UC0UcRpe30F0Sn3z
pk659HdnIDGdoHY9Xcg713R9EoBUXe0ZgPa9n/Fzzk4W/kThFvaGaKJ97mssPIU+
0+keDS0YifYtyBAbUn3Z1mGdeBTK+K38+RsRqT3FOS49vV9jbImbu0QKKO0ATJGG
S2XebcbCNHCiojnuXu7lpjVOIbi+LdyPgVN85wqimCkYOE/H6z7MtbTYSyeonODD
F8C68uSRzI8jr0eFPxI4naJmFIZxqdgr5+ZAYLwsx+ddi2oQLp6m3/OD5Eeqczze
ATOdD8t/G2kFcExrt3vu6908qbraaxP+XDsj1Ya5MjldinAnjE5MugbDX1t/E43Q
qmc5cfAbOF+NeQdYaphfSY7heQvj7gPzkMlk+lW/ae4dAYaRZ8KzjShk07ry0TYa
FCWvqaXUgVADVtgOg0vdoOEX9+rEZxDLV87v6caSsDudS+IXtJEucVKr2LxJserR
ovEccMgXZqWPQUs1MAqn3t9BPNAACK9wniSM+ZAaukMSvIVOmGg9kawQw9NNxFHh
3dToMSOsN3FR9fpRhku3AxUUWdIRh1o8JV9mgMI0FbguXSeuZnJfosyr7QrRxVYb
QrITvIPD9D3/BYgqSUeuTToX599w6bUWCazLtt5Gb1+LhNdnh0J5PH2KuyxjynAW
M4LzneKo6qti7JbCcnK4CcoXl+ZEwCks3aZBwCG7526qVh7i7Y1yPMSJtEcgXRoc
KukFBx47siqfcRqvRUIozqGmyRTAAVaP/gcJnGtX+N2nqtKVaXclfN8oVKG0Hlkl
L7cwvlulsTlhdB9TH+BQ45LezRgZjf/rDafi1gRl4MBaADuLiVcY7bqjfmvdOTlH
ZvDMEXTKWf2qmZyAintQ0QKWCYxwufZyTsRLo1nzWUBm9hhCVt9+/y1SQ9xqsaCB
w1qPnKWdAoxpNYrdPTEc8Cz/A/dc1C0reh7mFyRQBMtsxL00nTgwiKyxmNzAZBeP
KiKbaW0YMANeRho8+yyt7ZNQGBjyXVkkS+1pYAiQ1J0izPGoDuQJy77g7bCmFvaa
38IwME+6VZPNngCx4IDrJOxFmCAGwArGdFL8X/xyRPyGHBe9Ho/ZlV+W56zDeCil
GEDBmQEyG+glMJY73903/AN6BBXt2lGRccEEwKuch5OfCNKjhfEHX1VF2e0DpZNW
/uDdDP0Bd+YLPpgRTrPfpAAls16wumZ1mVoPfg8WwlfAOva5BHAII6PVv1zxVJhS
Ul4Io/N0krHaYsxsqFylPTnHJAbICpva8yRl+mPkmXmyov2zI63QCrLGPJ5tPFds
8sOPjSSrnC6ycLOFBfawKPbgJyqR73tYBXD189bzTWSHumDc9+8QN2Xf24U9USfH
i8ikTOx+9mTWOWy8TTtUoEN7jGsPC6sqhNwWSsxomqWsPO/gjAq2DAOISMHTnA1g
IgEiOPN0m/uBbiJCickxpfnvfbnFzuGdOobFvB61zKequUal3eMwehVYjsOm6X01
NZSrft09hFWAjv0vytQIyUYh2+l247Dp+cvMHyRBdygNPs3jwOLubkwPzJ5MTExu
on64y7EUxbTTONgwPv4zOSbilYjYFgUatFwuTlWO4+YMEI5ekuKI/JVadxKqkHC4
oB8sLlNAFchfnBt1I1DdiVbv83OL3xaZ0EkaDZ3Enrcz8cy1tBlGkbQtxrgcff4V
NncJGt3KiWMWVVO2pjIrCg3l/ffhF6st+9pDEvLTZ555VtJC6epBf1BCMzKijwcH
eXH816uGeF+lfXziwT5rcfe9udwRDkpyfiN81PhzK48Ny8s5Yiy4CPm6Wmy/IJFN
/QCfTEDCmIe9pxGZaxwpmki9WeUlf+Cr70Cb8pvUDnCpYL+Q3CX+403iB5Pixn0Q
uV4LNayPmV8hodNEVdASr7LYEfks29KlRi1O7QOFR58BflKXk7mxrYerrh2/qZ9X
tmXjLGEUK1eXtVHxUrs1SQoGPxe77HQhQP+jbQtZYr3USrECRwj8VCJLwGawtR+Y
oppixrJygZjOB7R+IZxHAysAfb6ld2pNFXBG3qWdB2v0lecxLy097xPNUJd2SHuU
07ZKpHJ8bcW11dsWx6ucJJ2psb7krmwQjwYNSUu7FwVVYyQDTXQeyjUL0dwlq9tK
i9lTtWfLCRHy4dr5DPzWIteetBUgRajDU1uTXOBq8iFFcCQrk+poVOofgVmo0EMc
GBRwNguj5UE7EVqwg54Yfr/O7qEXwk9IwAHfWExCvQvqNLohfIy7HWEPgTwIRVwo
zUCDqS+guQRO6yRW8MGbgHN8yw2JlPnKCbRuIj17Uwa121yvSizlscDp5v4crUL4
dF0YdN7zYrUCM0bf6iZLvjAwKP3zaObUFXrE+oM2xwOE62yVWoUXYGZVsNZsoZUG
XgidfHoCyLSsvUvhOrmGFqbTAgeU7ZFrzQu++QIlcQFycAN94ddka+QXoguZ7p5M
rAtqEBZkYSvqw6rncC7hi8hKj5prqzzUQYaPWqaND8ZOfnXaiI5rniBL1/Nua8OU
MKeKhvtoUQ9ONYktuVjNsyfkhbglhxht7oGB/SgUc6ua3gV2LrKLJHjQPK/Zyji+
fWxlOMiD/kUMUuTwHO+nlcwQn7Ww8llnvwWIAXyDrhG6Ivp4qq4IuuAXxBoc3pRb
mrefguEmDta0uHwPkojd4qrXt4bUsnPzXlUHi+MdKXBDz8IXSPo9Zbj0MNZrOK7V
xJzdzMOqxYSNb2oM0EECQ1GgCbbRIflaxU4R0C8UFqU15eH2+JynsaZKPPR86Jfk
HcLNC5m0de/v4KalQtzHVcnHwDR5i0DZqy8/qJZOzY+FcRn5l6gM5UOY13dhoq6E
Y4gr4OVppmql2C9fbLkRLj5JoSe+30i1mM/16taoCe14ViDBmNzmm76wAvUHEQcU
9memKXsstPiJSi1UklnfsXjB9EOfI8z6/E7JE0t83dtjhSyPENlqWFGyKWFPPMLr
1UnKf0HoGaTJIVNOIHxMy+7ZmfvlHMNfhQwaopYnP7xn31XEWdX0ZzAH6YmZGrg1
OyGlSUDRMQ+7c18z9kaBVcCUCEoRFVPQ/Kf9Fw0I8IWE/ITtJAhxq7MyBxK8SdVv
TgpgLKoU1Ir1HMvbMz96uYbcQ9GFF05Zlc5UOG1yKQz9RlWDpBGPl9o9PhuJNLN9
hB81+NyzmtnK4qQ021Qiuz58lPAURaTeLUXexyujiYUyJ7Co1WAYZHSHZSMdnhKE
UEhIeO3zqmdPHzR9YCNkRyw5mtHL14Xhaa4Dgp4USA3M0046rGYZSeEH1PoQuRQH
K9gQSC9wniJalJ88C8L/W/IAiXNBQ6xxp6uDcH6A6wvGIrH3uBa2S1osLIZZ0u8Q
Hqw0KvQ9fEkwxjW+mFT0ZSY/hcoOPIPvo3hhexVmPoAeY3s4JpsC3KyknKHnLiiN
tPuf483cG85o8zpr1kPP3VFdHuQ1XOXKOqxGy/Y4oQ9JATOfgH0nJk1LPgnThrHB
/jUmPBiWrKADxQSve6IHnoNgtsNmNptWox3m2U2LrmLywAJFIlxSnv2Ns5cn+y66
9tj3zBByr/eazVotEMAWjfcAB1oMNcZbZcRpQvYkIzd2V4OzZFVBtw2aQST8etqq
/bRqdsEf9Obj0qZrbKiJ9uBGCYo6MUb0mjSnEg/crP23HyNUtbRk+mUfnuW6SYEp
J0W3adG3KJCn7ag9xlMaX/pn//dWJBThIpSHBFCP60VG7ejHjHoezzw3JLm4S/+I
S6Mg32/2GCs26BKZgK+etZzMqOAoGh9hfk0YgRVt3KpqISwUc8aDzGpavFk4ltUd
wT0MHa21yvUWviijCWH326AgxtIk+llQHUFBRYwxosI78u89XW6na3RPjYF7Uzau
Rgu3I4vHMMCS2BXEI6j6UhWWU4SwklVsWriFy6/aM0xfucYd1nb9O76FZjVQlIj9
uA5ffYw9X/LiRgN/eqRHd5vCUBWVBOPUIRZsRVdux3ijcKEHqndL50gn4rP3ajDn
YWrHWrNYFrXy+DZ2davICJdzcjcJpdW18ArcS0tCXisHE/w1nIQRycj7KHcqXuwq
NBEwPLxDBL2nSbWQEAeamb2IM8I7J6rO6Jj8esYOrF3BZhWSUIwv+s7JM2hPMmjI
JB4ivFF2dJoYGDO7YI0mhm/HZ8RMjdwzV4KJAb/FZSAl6YeA6BVGwu77EpBpOwaH
4wOMmxEP+kGIkAr8zVv6tsF/lQstWjZW+byzRr8L5XS7FaB6w+kofmidtHrBvdgS
ycWFFu+nF56HdaOPD6qhszbZ7mAsYJnoNMmO3u5fx8QiNDVPs9F1HWTc/fWYt/89
swfvmc0BSFTiw80cLXufcVyCzd4TqzliJQgAU4t3Ge5CtfyoT738XPlz1LJ5wEqT
DAAUnvCvsAL0JvqoiIeXagH2DcK/bCe2x+w1hrDOE2uR6t4f2anr18HXXGILUYRs
9ynkQcT/B+ED0V2M46aGlnW3+GzjlnRlocIdvrk5nB6bRrpD0B8hzTxG6ooed4Di
HGnQEMYFGCBvIafXkeqsQE+EK5ISsSKXRgCAP/tjFKIIfN5bzK8nSmIyaaY3mMDv
TVQLD78WjFQgXAIstxdBNoIqrcewe66j2oBS7H64UduLtcbLG0Xhcu3rVwUphjax
UWMhYv5FPQhGxHNDDMcLtB7iKvnPrt8PYc0Hb9wvkTZ7iz9LZXEG0RoRzDDHTS1e
nM0z9SuJrTkhnmtJNrwKWNeRCuyERzaRcfKG1oFac9B1qEXDMtA5RUUAgCStf9TI
BxU8bFQFXDWu4cr5WOKam2T5fTw/iLlfvt8ML+dNIkKKp65rt1bLLiXF4O+hrwCe
IQE4I3V8noEYMiu5j7AaG0p1yNLBpYKkGFHOGQxx77apzInf29QF2FTpn6/2zvhH
RHaJdSP2MpXisbGr7R+tHNUKPgdUjbiFe3zex5muIbpqaVIKd+ykr2tkcpS44USg
hiQ7VbRwgSbh10G+6ev+hGIjS8RVuOVAHYaiQHP3n2KZYy9k6KqJygb5MlR3NIc0
W7+MC//+9rTA6lS+ZjkFTTRHfhpczZUCkPndwAGsD1i4Xm6UO+Oc9vBMAN1GFG6/
Qal4mCRGJzsrPeBoB6DbgR2UGXESelSibYXFU7A8mr1aGKFWKaXowQpe+AIbFbLr
OYLjKxWAGQYfz6DL1CIsEFn/F2+RkVlhWcqHA/Mh6TTYD9lG/Bl8/dRhEa12pg4U
H/99SGBFBwJFfN8yR9FuMrp2GKMXiExc++SIpIca1MbmSFNWOfHkVLkWPedhEnHO
22PtjEdLUz2NMWAsAEX76W1CGf3SiM8FxZXrfgp0zgAArATYHk4NlGsTo2YGiZem
VP/ZapMBgqQPAkhDxgEXbNaU7q7z3OXvxZvPfEyZWaghErfU9JrK/gvPG9SlTV94
DwQUV1Laofu/WYJ58eEzoSlT3m31nwY/x0I53ckEP1GMpcoSlESzuIMAuddERcCh
AmV+avcVObdidAZoc1FZ7k6QJMztM7XYWvvhIypwerIK1Z5Pb4j8pYyBphxcrW3h
P/FN+cRGZCzoMyW02WhLOj/W9lZIyGpS7hdEKmgV0BmTgnOkBxVmjXbA7iah4iXf
/0OzeXq1dbcH3n8Ka0fWHnD8rvi+G/Sm9c0YU7oXiVus9ZhRvS4ptJQXGYoeE30+
+wHHuuwizkCbmRM0mkgQpUVu4U2HZTQk7iMlrmsgJKWe39YgavxHWWfZ1HBhV6qF
GirpfsaCTL/zoBKqifJJv8t/rhFKDIq76zOjWv/zAC5/pMxU8SMGDar+b7d4JHoH
z0iENjOsVGW35GEgpeUR5CyvrmtzQdm83wFo9svjg0cCTeGr3wtY+4PdeuR0D0/C
HYAsLOkt3UgDzccma6t+JYKY+LcY/+TBQ77ndT1UDPsoyxvbxd6ibjzcz9VXZm43
4RQ3dhsX2VSoQ7vVUReWoHQSmwP1QXm17GaG9SMGNRDVnk3hLYJ3wKVEZ7zD5tNn
Bvlz3CVfVu+xwHXNrmxGXg==
`protect END_PROTECTED
