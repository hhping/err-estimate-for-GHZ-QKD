`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbK3J+4kdXdveAAwgsJGD4tnFYb6RnTDzgS5e7adtdrITxSq1LQI2j95vptG89uc
oHfnkslw/oDAc7BkcJshldDrp+InZkw0H7A8Lm5HAvLXgW+QBKiu7gldJdHeqjX4
PPFo0mciVy6yP4C4juxsqs+WSrVmvN6+wgWTDQ1wuJQxXRw4zY0hSBJXo7QHcvK6
T9mye5Ticgof+79xxcW+OTPU3yj6FZ+s/3J2os/kOCXMM6z3Y98k6EUenmfhIOTA
iSEEJHWK/SOt2C4QxgzrUuB56tJw5dENVOEU9qaPbvQCIJX/fqtvVTn1tyVVRJC4
1keX1wJWkpknpW4UVsNSrkAs5dwcHDIMfwsOza2kzd61AQqGL5W94hVqUK/rN4Qf
/x3ITVZT0h+fluJ7ZZvZgbjEvxdkXLBL5waEtBhCq2nFGF7L0vG7aUgRuxzXymu2
qGzXMR+zyAE1B4eIlx0F3WTsOm8sKjASi6dJq4U+iVoZKpeZiQoXJdTX9CiNQTmM
igTO53LORllzvpB0lTOQ3vkCtDsLeCXxuKFUuBPvBeXG/atuC18GAplqAu8T14Ve
JF+BN6MxGT1rxNXFvt/kP+UkiT+zChJF2TeA6vTpZoLCyGYCT6+Lwmfaz4isewcT
Cu6zjlxebLy4QxfErqvVj5JlWe1lY2BcqptqXPOLTfpRF15Y1ndjXtuNSKbOYn1C
zIdLNc6f2diV/KIoRi6qen+p9RoiJmibC/XQOHxcLCIH1M6dM3JIirZHhw5Uz3f+
jCREgKTcSfUjWJdKUpI+r7h2EY5Zl8Lije9kdQeuDEFuH8pBgMeMrO1H/tYQbJUP
H+4CANv3iDkipNhCXEEfaZyDktOz0XwrCQaRcg1U0uEFDpXEHmIuULAhehxBLrKc
bRUHgUnvMaU0E1ZtsrKGZzDvCVp2o+4fF953/LbWqsf4n7qY/G37tHfCov5yh+M1
B2sB5UVfc5Sr28Ksr6UQoJ9l78VdXuA4g3clu49OydKCuy57Le6kOW+DcKsk++Br
4lSkvhxFGzTmz8THHZd7IVEQWe58XUpI9dKYdZG112LeVT/3TQooqezyIQz48TMk
Stt57gwD9kBgOKRhjDiIL8m4ZWJ3tAbn4VxU8kZ9GROAwbbTi3avv8k4MI1QrxZV
tm6K4vo4Ho7Z5TRbbcAmWgnxKbunUi4RVV3UwOg/Z5vnGmEGTpuP+vP5+9/XX3gZ
pAGeO7w4+z4eGSvm84aVPSFpVupekc1c1b+uffMeIJZygBAPApOQOPj6R4LDM5lS
YGxKMvLCGWDFDJty92ck2vwiop93wMCjHEiAYe0GyZeiUIRKUnt7VEEq54GJSiM3
XMxHPfZQFbQYs6YHlxVENg==
`protect END_PROTECTED
