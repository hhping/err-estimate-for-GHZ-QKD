`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhK94ml5p20Bcui5EB0NwLpEgt1WNvaZGsbhRhJOtXXrfwRtdBUmtmjrTDOAv5oR
nht/lIXFsxrbMgVNy7ejprWS7eIbYDe0X2dYn714TEMf0qe7jM4CnJaIs6W9dJ3y
p/xdkycZtumh/a/JVKyTwnUCQvqQmXeMRxOiynlAPthvqHuQMa2pVPLNbQX5XnKr
jt64xQuSRJ8d4sbVpAC7RFMnrOLSny+W/JedNopkUn+QVp704n3QMSV3h1yeBHga
k3UGRX32tTs/DJNIlax9ns5/fNSzjb7UCBq3T1IltyY=
`protect END_PROTECTED
