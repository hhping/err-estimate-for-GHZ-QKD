`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/rQuhr6REygIrd8IdtpnwpxlgFf/tWQTf3hH/o03CuEnnGcuL7nyghtSBlFnSQD
E6FabSAeUUHGSr3xLI3ioo4z9feWCYfTuObAk37RH3FGEmWRqcsk75m87KDKJJt2
JBLSyUcT7OZweICDhAujuP3vCVZcbCtIdO0H8qLc7+8hRVhVmgBXRnNfQgz9I7Lg
oG0nXv2a2KlOBaGhkzmeP941YaavoZFlT3QPnA2zq5kHNS3t3gNDOGM+2Ltj2NCG
nKEvjBSLI3iSW9u/8xeLLHvuhApobWM/jd35AgQ58dIMfKxDOf1gO48Zkw4qi2Bb
+/lSbQP/XxAEr1L4DSB0TR1VXcmQ55G0hk3CFByP2Xsu/al0YQdjlreT8d50RIli
TBNBJUlaf0FMi3oXUYt4pvj+kRlwumAmDeAOOGtk5M4RRsJiuBT3VO8puW3wGdkp
8g16awRXJL0SsO+3ZW0KAfG7ptNOKJVXecX+n3xhR1NFD6Xq36g7k4rWn6/VYB9F
vxPUBhoeUox3hbIDLXEJ3L+v6e7CKmp1xMovTukqeTCn8p7gsFY5Gmu5QkTM7eG1
G8ML9wpsAxyOMOE1QhJ3yeCjedZoq+HuUohQFUxWq5wbgpiVqQsCE3c15KFHgKwB
3LDkFc7KhIel9RAditc80l3LZg1UNB31hbH5oIwiwKPicU0Cu/+hCzBC8xnGcb1r
3kZM5Ng+KvkgdmLu7PMb7foqzYz1mgk+y0dGjAbYRcC4pV+bwW4+cD/MNAn/fF72
QhsJhhz0UMBLQbPlvqub3obSo0UmOXWuQzM9k54XYA1nXzc8qP1FzJdBxgvFpA4p
Ndn2kXBB/eUQAHswbZBe7eNyWhAAtl2vrUkIcNO4gyc9WTC8fIUW+61gxJUz9Kyr
EuSOkb7ooxUyz80ncNoO2eTPgV2/OK9XBHpzP3yBPi/3nfzSuFnGp8ASv96jNJy6
0w37UvEtz7sulB8p30BgqTcZUVFtj6iceeqddLaGbZuB3D6xHL8Wqs3GtgngPKat
mXAPyvataTk0lwJfENcVE2V8KPyzdGwUElFyl7bLaVI/SF/t23KGiwIwLBAmPb9e
p2inh3dSTNsuGkPY7JPe58s8i4+s+S4K3/lfumng/KZkDRzhXhRkuzFjKeRRIbe0
tX7N/KYp52fx/efLE6N4hTzATWPjj9N0AcGkxecZ6IP61rsZvrm/nBUQWn+yKORI
3k/1Gp16YyirvRDOJsYZG/gjNYFXyO3iu+73lpT5HiU=
`protect END_PROTECTED
