`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9DIDO0zd/YkC+ZgZbVeREBdXCSochJlvYt2QnNmBPU59Lp9mOhdPVnBG2/cFVkL8
dLOxV5VCA8679iljm9B6IGoeWJIFaQ6/cUlbZY3E5Sr3ISv6tx0A1ueZ2kF059Cs
m3XyCoCy/fGLqcMh2lgMMeZ2WDj91oK4YsHrdszlr4Nvr3UaI3OFr66DlmmNX40V
O0HEc739QqfUu81OkyLbotR0byxMUpOlwXmfNS/kdv6f1WB2p6aWMvd0+QijAIkg
OIFbXGxta7sEIGsQjSwmeSNEcVg8WnR613vshgqNsUR6zNh5Vz+dSorhBLJMgqNP
0yneHm3P6NQ2d1Qc7qIOLm6cbPrUr6YtXGEw+0nzkYUNkbxihPCFMhWP1V9Ffe5N
`protect END_PROTECTED
