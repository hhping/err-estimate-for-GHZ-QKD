`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0xmA2zpY59j6EjtxokI0RcnyDhpZN+AB887jRoSJdYvvEppdcvV5w5Y8RWGO/jps
L0J6JXB2iVPd+hwyadYUg4nmDOGX9DtJjpJtgBi6DF+U9Gs9FvYhSacIv7zqEE6s
qSzwQco4A+wMqd58aq+9MNmmBmhvMAGV8Bd30RWDxlsDq+R6u6Og3XjBehE6qGuD
5/seTL/xuU0ndeGfiviqe7UxAIedwVKvl5nKg2YOGvLmgfMbidmwiZkYKhB6gJdW
lnywXHG7T1lIREb+1B82j2ibe3fwpwN+TWKXQy6S0q4acMq3feNsOLwmVPgJBH5d
Rf5r6oWGwJtjXxnvn0TKol+DRBWH1shST4cQmhiimi2PIMdDS/FiPnlKkK/u2k6H
7zBgW4f6SQmvXwqGkFVDKw6duvIhkpmYj3Y6ZkmkWkTiJQeIpdh4gzKQ0LJlokqP
wgAwVE0eALYQSw1hca+M2j1CUIS5BTmgNKSb09HHPCU44XhafnBmMwckXCBDOhg1
GK6iGZT/UXiAARV4/59HRlbvX+eLuPTDAxD01Ziii52zrDdw3K0aQ8k42xb5BFRu
ChX7GWnZ1yU3Q682wQqmrdMZ2Mq/rghpamM6gOAhvmrxqedmDAhTCTF63gy6z6Zg
v2xXRuD5rtFycYqFsR4yHYDpoLwHBTxCjyH7luKkyPY1IDK9ZAPHciDI6Kr7DFXk
lSqhk8K4qgbCfRkCQzj6Bd5cjB9a2opZ2aLBZGY0MZ4MmkLURsTgw2I/2JcOxhLH
3cYbTOrveP6WB7396D8+8jnR9rWFm9cw7E6Kru7iMs1c5vZZRPHEbBlXmU4Bnx5g
SYPeWDJSo9l5iwjp7C4aGyHwpZBeJgXjziSXdekvMsrv6vYzpx9z1hPrrwV8RJf/
vrdHRaehOM7nIvwcsiixvnAHTP8mtHtHHBzV2OebRgT4dETRXEv82UPAP11y2u2i
cplcF/eF0Hm3SZLcoY/KwkGwHDJIfA14jP/MovntvFDP9e4PNTTlO0pAo/Mayqw8
LhsdCVgaH7KuCcWaxCgCvTxwPh7oiD/RMdGTSpqI65m6HOH5cuwZZzyCx8de5CnX
Er9QwW/Ix1VSl7sis9wIpTa7gn1LGzcq/KjZTWyQ8Et7Ak36+wZPvnjfNW04r/5p
XrQAET9uoBHPMzYg2q5K5dEQkDnL/OclvXi1yoR1b0UFNMs1dThrw2tMg8kXKJaY
aj0XuhzSVTFIVHO2VKRBdXLbB3FuQ+SjdR7GDi7lBUqy6rw/KfAIHHVd9zxmo6dG
We64GdVt48df7Fpj8xk+afIbSX98WnY6xfR45WW2OeJF97U6tY10PmQJOv95ezZA
21mpSgDScitCSxz45AFHAm5DjcVSz86EwuhVBNnYwcQcRj/TWkWsK9TjtpWJbOUy
VItz896P3SFPNyKl0WNNp3nZfSxzcRajAVAZoT5M2YGbTsXkAapWtT9ARAWHgsNh
aCmIfSNOUW2fbtFY7znY6Q9KL2yopTjbMAbXRS7GSo/BS69l6DwtsSVAknfEKkpu
rp5BQPs1qK7+xab8exa9kCZLGehhAi5VAPYSEr6Vos1c6m3EaOLqEL1ro+hcWATu
BCBJ9xyefVd7Iuqm+E0y9b0CouQDOUAbbfC0z6mxu9I=
`protect END_PROTECTED
