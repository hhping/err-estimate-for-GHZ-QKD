`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzdvQzkPDtTm5mfRRcPnQGngA/bFzyWFgR3H2G4f0qOsaZl7AVRfCl6oeO43y50T
IxSrERyL98irhDiqip2/bKPyp07tZ7nkGhPzkmuC1Jg2wDmuP4RxuSlH/1SjR8My
q0DpN2n1BzzHWpQXc9W0/D47L32BvoGZVnLrG5Xax1O4/7tIRhOWzgkxCE//2ruL
p1KwaCAm1cBxPnJZUWyNr4rlhtZJi/h4EoluY0AFTO0PcZusyUlwajbDHmVk4Flz
xgb4OTTG2f0LEoW4rCGdUcxKhZ+S4zib69de7Y1Vnf2NRn0MLJrPJEf7UyuOj4Au
xFACDL8DA5vABHxRW1VFXaMjhM6QbKA41eR7U3LbLoY9LJy2kWawd8Mp6lEsIhZ7
qbE2c1o+y8VavOnZ41CtfdGX7DZsiRKOQWdmjAfKERfEBzey1UFh422mLTIXBOzj
bEky9tJ1bUBoAtjiDCAiz6PqFFMxbW466jrSgDC1OIXszdPVCl2yWbHtv9/0t6XD
F7HJkd/ld/4LOUP8D8tdIlxV9+UB456U6wkI+AQSn9OBbZk0nIVL2imC5wsf2j/X
lRswEcJ8hkJeyQS0ijb5MD1wyZeulO0cMDI85VRwnVV2uUxVNFE56VlZvt71xg3d
rrL8cMGugXlB0NJ8WEAS68PG55b9CgG+1k8BChm/JRnNaDXxwl9ddLMcCO0Cts4D
tNv7TnQRC8w52PQQXFSl8lKgjN80a6kZ9uzl8tnnKaD4oK7l4rhCaiuvJFGiWteM
fd175vJ5GhVv6oEIGgVpS7pB0PkrgKAsxmsgLPh5nL7PiIV6lOv/SSQ4V9wVAvXT
hjgVEN+ZVjbjlAGlpkmnnA5zBFl87Y1+8plQLBsNcggR4mokTPB2nnA4wYZObSnA
95iUvJwDrUDBehZllvvIvSBTuAgJoGYFVNx1a3TOtNp+n4A/KtBmTIqvn+AM4arL
U9oqloVTQ+nqaTo0MyMGgvUEmNZXURjhuvmOD6/EprSE5/DVmCQkNE4oVHhgSCIF
uxyDfRHuBhVwYntyj7ARpXYD1RS3p+vZRXIObr8l/X6bzLIYEgKeiI/QCSTW7VTH
IZnOmCZUvLo/qKhujAJJS6TqSO7fmjyIyKkKnhGwOemHjxMPQsmGRH2PpHs2CoqF
cXouaHvfDzjI2p6QRVdMaaeMTqcgXBb/B/mYV5F3ZwremvTHGhFL4CBeAszjWlYH
Be4O0VvRNfgMrtGvK3kuZsyyJOscDCz9IevQ/8/iKUr0zShUfEbElofeCiSCIQ7x
T94ydor13AVEkvPy+PCR8A7msX3uaN7ZXAMXIJ7KwmdIwXys7OmDYLSgTIZr/iq3
HBGKtu8wqN3vTyYOLUpTHWskqgrQfCeeVKT0kR76pA6TeVIXleaXgTwW9wW2/zO6
IGxNOLRDqsxh1dlDJ4vvQyaoaGfdxfKppVw3KROmPMDPTFLgh/kuU6BDl8wKXBvJ
Ljy6tKolFZRPgiD0yU4HCZdHCBUxcPO9t4GXEvzKlCwGE6UISsgL/ubyKqjnU0VZ
yx9D3xPkoR5IVVB2tLpLjZpNBeQ1Jodgym4bg9TTb68F/fD/9J01CwMy/xYcI/l4
TtCWiNNlN3rJwKAj51diFowM/361SRW+BzJCbzpIACDVPPalbPug1+Hvkq26cn9m
T/VS0ab3NBtnsy3/8LT6DmzHKvvxr68GwhTutq06ce4NH5/BNhnFyF6R7eCfEuq/
QzKVJHhNDtiDy6/cN9KeesXwFWd8jWGfnUqIUxK5lqR7yguBaZgfxJ+8jLn/aVWA
5o/dLj3Qam6Jn14Y86uXK8/xF8zSSQyikAgbtQW1cLTqVDDIqlaHRtvvTBRvXHIP
YquImyXC0EE9A4/pZ5NIe+YsdxpH5uBMzUt3aoEMKrDZ1GHnHOP25Oqzkp8THedS
7ApsqV77Dl2ou2Bos4PJb5AffyP22Z45/snze5nseMjN/miiF9JhvMCWrwOrKfNl
Sv5aftsVnzy1lLxXQ2APjM9BnUaP3g1tQDf8I2QcVYj5/7yKZbEcuLQuUOldfNae
fTq5R4Y/k7Rg6lDuEZ7v7Sc1wmxu0Iu9YOTPGA+UvSVk5fev5WQoA+5NAmfqRfML
8NtJsN8oc+q/C18K2ujSYbUDamgcB2Uyg8M54zdBd5dYQNpuF6e2l7I2QYLcbWgd
+m2kJnIqsHyF4j1dN4fzk2jpYrrIQBzb+YzLLrmao1vZYoiauZqO9q8Fm/FbwwNc
LI9jmqM6GjRiDMaVVHXAfSXnT1Wo7v1MdBQ/aIr3NTSPTHJbUgRSm1ZSnq5XpDvQ
0Rh4q72Eop/EEQRZs7HFQCBaeJ3qIZRVaSlRUZmLPMydp9/oza+/o/YCkPIF7cvC
1WwuzQ9AROcKMeahnK2NjTxaP4WTpgxXGeTzmKBrMq2cxowxkopIcmOY+wgjt3xe
tBlCn6RPwooFsbflcHUdwi9Wv0qx63xl1zUg5QXlVr+vfTjcfxP268KzY1hkbqA9
VUa6pJtBAMy70DKxe0BhbU09QIc5VLd4df7jOYi5mDadDDeyWKI3oxSq9XtJW4uo
1DnZGbdV+KRoR/H3kaSkPWjl6R80WUVfVFF4DtrnxkjOKpb1gVC0qhF70MMxoVwi
+UrZhGatqIo09xW1Pn5hUMElpUSqwyfFxKUz/QNLK3zp/cK0JX7dcOD5Y9/rTHjU
HY/h+ZxWBm3KIadYds4IN1TeAMNVg3CeajJXBV0u50/7/tN1B4WeD7Anx9zYLz0t
YsK0zIg7WdZEGIZK5qPkJF8AfG19JBeaRW/CwqaNeJTHsv3kFycz63YM0aGkXW6j
sh2ptHafIVx8shla96kTryWjzeUMKxlgQ7k5Qmfc8arjPSVhV787pR/Gq+3+wRz+
/a79YYYCz6cmYyv5t66rrv5+0gEMOZ2bcr0FtSHkxlJ8xcLgGw6VYDYKOR/+rbKO
KdaOkeSMDCSRcI+ovNSw4Jq8D9tS+RPwcQ5o4s1EnR4cjfqa6XZfN9mawnyZCjSe
jnpHYFnaPuAb8WGOTXUZk4Ak1zG6rXB61CPL6sivZxGb5abAp/8ef4WvURk+72RU
hXSi71fNeY8V5+sVKmeV4//K1jLmCpXtw5s9421mI4RpWiPW02m4EIouxooiuAdJ
NIQW6o4lrBI1TOf08i2XoYnjiRDbx6BZuKwyKj5zUqq1bTJ7Jty+oCldrUAIQW+Y
lCVXKs5FZTeO2ZexFGtBFzy01G04i++1RE31yYiYqnUWGK4floYPtV1kOkTxdWGu
1NgELL8pu6CvGhmbst5pIxbcvzLqScFA2xmU1DC4PvOF6Wx5WOa5YasdIQ9+nwXt
qEb7+umPUmTS9nJkL4PO03loM6Ff/hi5CwygkonDD38rrHsQeqYW0sTrO2i5UqgY
gDDSEl3jVuZr/H3m82VPO010corUZp62JIAxpiL1DDswn/onDB1T5GcCVhHycHsM
RTltWPWJh15PHheiMgQNMuWrtOtNB8XEPHfqO8Wn75RTmbiLRUGDrWub7c8xN0ST
ifxY6vrr1JPV8UAkqjSh3Exg7g7NQpAGsLTL49j2IxOid5OY1lt2fMnar3WwaEnG
PBijkI8wm0iezG7hv4TueWznqVqF9uH10QKrzGBLsym0dNSAqf8hF0DYJlpqjBMS
G/vVwaTOq1qeOB/xFvrt/Ng9wATJbK8TtFpCJgw9uMVvVvQw/gnTGjZXxsyrCkAQ
gznH3CSk20cXb/BYzQrVdRQRSdGH4o4LMhOLvupoLfbSHbuinMTjX2B6KDp99Jb9
v09WhupCMoSjPZNNq0NPD1cb+pNqyDVPIu22Mk4UKb79GLzWFeGLUCDCgtdEXJgq
CLzZzZGBoBhxkQuvC/TqRAkzyHg9ADxCkGzRiuYrSB7f1sg1MCqRSfMovH6xQzED
RyxdYOnY8QvYENFnMr+/9D02emTcWDEAWhippG1bdPZZltDbgOoHsv+xAMVan/Ha
H1dbHMK8T8Cwp8ZJRo7iX/GomSh7pld3kgKaHmY67O5+U9EkkXwKnzUXX3vgmSm2
3nLd5wppkoyUecebBJBjLT9IzUYXQCq8kJghCCuva8M56hK3csSC5uqMbsLQ49z7
YrVbzdxsJcu9Xu7ZSOC6PaI0G4x3gDk8gqa+PUxjVot4xmKaSCBn9FSPSzfCbt1l
enjI/jq2Fdnavv2w+0yVZL9oN3pbL59F/ENdr7pWMUb14qhaDYkBXb23EUPFTKwr
4RUhV9yptHIirY+3GLrGFZfkAs4uzvbtCgNtkzyxzoX44t4VoGWbZcnKrzvPeuWK
DCFdKXFuAw7WqmaNPEhhDUi8fIlF16yhky6tNdbRelnPfVQXMFgatvX86iACWxiN
X9To5QRX8cCVs20L9fkuz+Ykt7UtU4DPvVvhhTyfgN2hE225WLO37coPONZ+TJdB
ADigrZe52QTmIKxKcD+c5RLY/jnhfnVZ7hnlWqpjK2d4g/jNXe5A3lVUNHol9xfH
XW8IucAyeihX1ZX5ke8vlYPcd6Fe0oK/qgpqlipN/1EuB2XfsvdlhgfP79HexwRH
BGNZhMMIE+NRc9aK5Gxn8/KROnKIsnRXd+atX6NleMGTOfGU7pmepNC59+3aqdqp
/F/hWZwUi0y3bLtxCqSyLTg4jyv2ytjL1JqPHdB2CRll+4Q2J19Bsm/H7ZSv/XuT
J4xqQhNkQQSye4FTCK73TQxKRcOb3eiknAclRZdSy3JHW5iWmoaYccyRvBFlvdOj
Hz/lIDtG/mDNlLEY3ql0Tp7NRB1GJ1DmaFt69v3OPZzGi3yiPvu0PCsIGDQOOfAF
xnl1U6RUroGJU/rSy91hn/PhquT1R5wWftbaBW/evR+x+bJGowwO2fqdfBJc95h3
1SyH23+Eso11vnTiGGzwWnpTtO/wZodJnR/zsLYJ5Tu8YTeaFjZs3yVGhe13YIrP
cYsVAn01RhTioVOtzpTSgeSZNAWQc4knV1X7tqJMuLy4Nk287RibxIZWZ2zw9nrY
oSIvcUR5jFzry+auxVrvuj9A1c1Ad9iqpyTdavxrGEstOvrkaB2io/818IUHPP6V
wA+i1FF0aA+dGdr/gFW7bNjYfrMvEcqrd9e+/YMvWNp3/SMO14uxvF9Ip7z29wio
+BUbafqidwMEalEvnPs74NEdMiJhhs9DsBfyRBpirgflhg0Det4vPtzaXsMRsXFp
4lq7HIF30YxqJ6HA5pVTCl5AkoqBLhdHxXuq0CeavbaUQX7aq5VcsIHVdtVcf3jn
lleo4kO1gMX9E+WRsxdbuFDug02vtae/6mDVnsQkpX7QpyXVJHoGq35+Jrp0hHON
r4a9I86xXjxxRoUaDrsfcTtC48aoA+5cRGr2Se+lous1QNVkGNaBc5rYF1VwgF7S
hRguTgeMRl8TGoNvWOoV+3ShniuZv27guu8+1PWtTRCXOiqoVKC5xo49vI1sPmRU
nm0gh8SG2xXyJla/zxwnRQNsO5ST3PuMaZ+s6EMsfxS4lY/QZIuVZzcLTITfZrEG
TOcW2NeXu5MBK+TbBlGHHkkARlE5BXygCwf6r+MYET77K+IYZfg6CyftJWYORGxH
ef08rrUSgBwOpZ2P1sDmShODvVh8wodYbUc85X75obH5yd1p3lq97ubiuNaFBBi8
17audDonavS011clG8uGizX/T528giRzMataP526wh+T2SUSTB1tcjXJ6uTHaUBM
IMiiQSyvDhA2i5mu5HmioLDU6f8aehuMtosC3JSOkn0XXEmf9A/QplGWBQYEnXXZ
cZgRH2aaK960klppJwKs6tjhhKhRys1KDkbkbbalzLxMgJ25St299f7HuOWM/y48
vV96dizvwRwEGy0Fhcam12lT+j7iSrpKUyjB744bJDQEaG7/f0t0NBPWpstH76aN
s8PxsPC5wEwxuo7L6cvDvK4lQ0ku1TYZk5gVf4XV0f5t20cHbx5rrDlWGydH9Aia
lVZyuOvvIDz1sk1w3TxbbSH/X/52zrb6qT5MHacVXIjm0VEW8MZUGIprymaaoowO
oYnzRgW/KQ9t1cq/TZ1/BVbAVW4Y+0L/pfn1bFqg0Y39YoAPwDe7BJ28jQUJvKkt
evOMTf3IoWq6/XP6xa5MwcpM3phIdXByloO9uwtwFpcsEWzpvdm0ok9H2p1M4YA0
MybTh11csiOo2+wK3cLN3WDvtQEm8lGTM2qhSvGA1/TNpkaJIQEN9pSOuBWlEfds
EMMOvQmvn0awvn8OD7fp6oKIi00Pkg5Oix5XUtEOcLb0QCExUWybK+opJAGz1EmD
wLvfHdhTeq4cwBkw7oVULiXxjFAg0NUF4cUg+g2OgWrroaRGhmChM4rJXr1G+5QL
4sy2YKBrZU8yV/ySfXxRZKVzhBpbesOiYfHrjS+uTxfSAX4Y5/UL9QSG3s6ASh4e
jceL3XkICqbmWHdTjwgIjRneZpUsrdPNRLtRgLIZehNeJ4pZSmQZ7Dn2+Qd545+D
ief904N1+O4917i+Zx427NIhzd5taR12JfUnJ2VimK9tM+OJ8grhfTLZzJbgzg86
ysbXZvLpW76LjmBoBCMRpvlACojv1nHMGuqGaj5RujNcirG97Vl44InkYY6pApkX
zbqCSbvDvJO1SW4e5w98BiUHbCh+rucNxoeP7PvogPX0/0wIDh756gnKthkFGkmU
B5ywQzstOh3wic/iVzyCduUMJ4yfE9dysTN8O8JtUa2YcLtkRWpVfeVkHt9gmtFj
LIw24dI95inG0Skutme3DF1axJks0IfafFV+JxPpWQzFf0PXYXo6uUz/pgM150nA
S2Yf5u94z8OEitNz9jHdxNwNf3NzIf2ReoxQYxwkYchGRcdeMobkodLwwne+r71q
hqayJqx2+/d1XhtpZKGBm3yeSySlpaIDbF+zRSC1TfQG6FrwryDpAiADmQIJ0jLD
PG0zIB4dB6Af9QgbRugiU5iKnZVbcpujtH14FyyNHjwo/JwMEDt+FCYYtufQvEPG
00pROXwgF3G2Ez8x5jH7fj8JLb+IX0g92EUUbnrB/TuGcQ62Usv98x026XFg7ESG
6nBAgWdAq54grzRso5e2e9Ca7qbUAHTjzxkwisciEfh3jP/rWAkK+ZDq6ISsbTkn
3E+aeHPPFPT4kNN+w5Wq+Xb7VP2ko1UneJ/qbenQR/wOB9OEVf3+yl/6/9Dave35
c+6Tp1eeciYoXBWxbCAY4dLWQW98NK4SoS0BlVDlaQ3cJJxPZs8zDJfB5fRXomaL
FzVauuwSp0euW0I7GF9XG4COA47vAqEyuwXcD2hGs+2I84QvxBQEUt6dgVpjyrMR
ehfVGqEd+Aaoa6IIxtm69ft4mdcPcQ2xMJzR9Urk47z1BBR+HLH0Nfkc2uR3VgYL
UeH0H8PEdbfXQckh6Yka2Bx/LTQ2nHdr2+milnrlyKRbFosIZD/dfxrKit/jaqxC
pXYcOadBdPBES5OaQvurm1PMWhARQgfvUtl3Ls9UhFi465Sm+84ji/TPaydUbrP4
PCwLq0U+gI50xk9pxL2W0Lutc9TdaTl5Ppxcb2FRD7eGG3bt3YFAMen+CqSTbjJK
LM3W6hzQTnzMAHcXRGIgT1h9095I9iJjh5riRtKre5LOqScxR2muBtJKUKK8Lv0f
Rc6xz6+AwVDjysijRUBVg6J7u0z6jzuU5+yZsgrmg7h9rZ10fme0zhk03EmMz8nV
ycEt5s9bfshm+M3WdfKxsY48W5fm9LZ5i+67dVusQMllBHmDHpbYmX/teB/IeOKf
GenC0HuupMOYPR0OX4NYPFkaU83EdDcZiOrdbc3CJTPeHU61ZbmAeO1sc94SaGE+
zUk4LpDdpVZbqOc1piQDIc1wXMUmhCa9In1cRiXc3D0QikrNPvfkdbz5PfTWkvGH
3eVGC6K7LkJPqOSNxA0afOS6HQEaBRSz4/F9kS/btYJMUMcACcBNj4EFp0S4GOSW
sBQICtFAa+NhpZqwvSIdlCsJAkoTookWP3aRpU1R5EkuG0YNtRom/cz6a4fooS/D
M/tK/Ul7vPWQbpaUqiyt1yC3vPQ75rvOTLUmx8TxuuDtAcaENd/ISe4cL+3uLa4/
fwR0AIBiK5ALx0S9mG+zRpyzquv875JZDO8mguIEu8q0gZhsEQ+QYCMB2hXWlzM/
K5plgXm5RX/m42158CKyOANX2QTuJVgQvVVhu0uqfdEILSImbWlanaXp/vKy6vtI
Ka0ErlAS1EL1B4f1w1wLe9i7OQWSS13JA9OS450ZbdrJGB7tKuRbAV34O1yfvxHi
Wj65Nmnt023z3o9IFAa1tsa6U+bqIkTGsq7KQYD/Udr7Ow6/1Af6EC/iFpUU/f/c
mD5rE/mvZoCwc/gmzDMar8doRtDOwXM1V9abXsioTcn6KCRuOyZDEuQOXJYsmHnL
LG1bB/1ikLMJPNYYRG/6ihmfybcBDJN+vvZEA4SCSBarCO41jaQoe4NHWcC5/Xof
CldODZii2F9uWDONAKdHMktGYjdu5lOYHVTypuEbH/i5p7sbHSQ+n4NKx5F1NrgU
L1h7mqy0QkbK+KXMFlfUYARSnYZKRUDyTvnYOIYlyLUblXsZbp0peGh0EKFZjLgc
mkYTsnhzEv2ZutiCVFI7HuTn4BX3On5nakfzgVMs+YQ8ivOL/JUHwCM59kgIhY0C
gSf7wTfV25/w8Pbps6VCbtzp+tjmDtj0Oi3je9ayCyxHfT2tVE8NApqm1VbLagqd
IO5dRRfHWMKuHHNE3Oikmbipx8HOmwNwf6LY4KgmNqfYniN4cNi9YXlFiJ/pg37z
6fsXNqxq9Xmym8Dmf0Tcihb408ARDsEE0BedzQmGXUhQohfF3BU3elUYfDnFmN6e
y6rSCpLsYZn5cuskt2dVyePIFwh5hBsqLvGs9B9vWXbvhlH6OdYHrqym8aF0MzVF
2sZs09kl55UpblPhfKmdWeCvwJKyPN2UsOcqUFrWm2lEA6d9whIqVbSZicq7BDJL
drGkwDM7TktitFfgTuzPrnunW4HXAJ5iwbV4AGW0JoTHAJxmCzc/GEeTo9/3UuXf
wIO6c498OxFzsfKPBXFxiRbAgZZnYPpyJSgR2Y43TKec0tLxQfRX8nWm2r4Yv/Y2
4ETdYxfFzYooQMTXizMdY53Ly/Oz3AqiNjFsXVrs4onjAn70o9CghTBljhEk7BX/
k9pOP/oYXSMK2QkFaJlDEAozkDvFusjHtLu/UJrYnSfKL/kYyVVCuu9EXKlp8W3a
TV3p6P5hdL5QrDhQK9RxEouaKt66AZktm2unHrQ4qyX1jMrXb8UVqGLAWzijXHyh
+otaFl8MzaTGYiIUcHmIn5wC89mC24vjlM/ch33kWhfgkCOKTvczIEPb1EllksUi
G31aaDg5TCfvyrTkAP5imagOodt+fYuOEfe0J632P9mOaN1RiRf1Jit99s2E7SNz
IXel4tLmOBgtM3pH0K15vDjTLO4GTctv2Ob3oVme/gdpT6zXZhp7ZIiP7LeCuHA9
CzN2ewkvnT6FCnEbhZBC02T2j6TmX9DBOgAS0wSqKN9c31zHwOymJtU3XMIADQVp
DgBuahM+N6WqSf1HRhl44ryeSdiEqGJbS/jbjvk9UBDubbkjYwmu5QCT8tJySzAO
wqj5sXrsJ1Uffj6qDLGacRmXkwUic1ulmWw2c6Y0p4xK1d+tXWurFFkw5b/2hCDU
gub24ECtk95V9ZM3scdP0cJHP4uOlRT1tbcXxPeBT2QGmdGURCsh9w8eE7skstRv
i3OuQ3jRy10HDjm4g/BpsAweKRlI3htmApbYQOAPLENQ/X8dkT6E3OaVQSR/3DHt
N2IoFGb3A3f0CofvVyQ1ddpogQ5jV7/WUaVXglCg1j+uQ9iPH7giBY4PICpbNKwJ
xHsaHVK7vgesNCx4RRuLKF1GSNS6tqboV0j4tZ37Hq4wmYuwxyNBJ3gRXy1bo1Lw
O1mGVI1l8VV56FTaNYQSSpyMDdP2D38NxNfiaPX4QgiSp7OYNSXlmICRLhMCPgJT
UYJbsLXv+/6O/boG8ozw6RRg6UYbuKbMbdJAvkC4AVEo7oQO8kmzR7Es5Qgzcw18
UoYotJDSfivywz8wCbYIWExnsdRhb8Qtgn1yGwcdX7rOIXd70QM3giLMuGribfSm
o4of565oyYooX3ZyXb1ut0ftMAo4qt4sTdx+mCR3EuQl8z/gPoJLkTopPY8zLwhQ
VPsGqnjC/6KLa7Dq0O5e2x/MO4m3FBZ965I3bsuCJ3Vu+xS6yPvFdAS3EO8FNIg2
DBZX1PjTgssDuEH7Zm5bdE0i+fv4UtWVHFcVzO9ZkWZwL1+OghriQWlFylXnTTP1
R9qn1Vo0DXRt9ubzcI/H5Zld7unDiHlIKUjcSXNrDK5z2UpnQRbdYB7X3Skbof87
5Chxjvorzt01wbqnbvDCBqkBlFPHP1SXkKrAu6SWoGXaSFlrqdyI2uU5UC837HZI
LvaaqgPe0LBFDlK3Sv9/UUyDFIpwq4ppOgQMokoBuTDlvHJtUZyAp9i3mxqpRgFw
tBGHuR4MpRc8rHjw3aWl/8gTkJhUXR9QZE2E1pa1mWE2p/ax8pEuB+ZRQwl/nntU
iIMPSfWRtLhSQRg0PkuVlBmZp7uq0uiayIU2sHfinYxT7H2BlcJ86b4OLthp3EBt
uagYb64cuecyEFKyc+OH1jLw6+Snznw+/PVWjaoymdAScwErrZ8p2698XDtv/Wwp
KdiyzOOGKPQwMFUZ22eBbMVDIhtG/VNn+ObgZ5d3Lq72xhqWmd/pmHrTjfOBVYXT
kpmDzrMcCC6uKHfeA3/Ok8khnIA2JntfBGUcn3Q0sMduGEMKr/NEjoTnDhYvFzIG
HwJc7tCyg7cCgrVeR+YpQs9ahtFNPfXeidhrkXxQaGEg1w6BQ9AJhS0WIA4x/l62
NyiqCrQxjS6d/UnodT1qkY79G0MgJrLMgrm2VPsLx50jkAf+lN4hGumEm40/JZjN
ZbSDPOFszQmpeuy3MXL569Vlltzypljk0vlXuVD+PQtI2XOZY0nXnuSCwdywpnnz
4qCoKZZtU/xIHSGn20g/8DZulaYTvL50EbVURdxfyg9F8MQ/EjRUpX1nutMrcf9F
UNY/9/FGRZN7NfQPjuyHpgYYI37wx2NfLNf3zPxIAVnwpGi2g+ISW/EEOB90g9nH
0Y0VkePdQaBgNd2z/Nqaj30aOHibEWQTIhN6AaQU1+QyTWOTTPiyp19Tn/xxhTrc
14C8r9kEaZcvOmzZFFvMRZNuecS8xgqfqu1culNaNHN23npX3cC7xPQ7GWIMh4lG
cXSEYrKkQ10kzojlBUaO1GIRGcltq4YczUeVRV0yTjHu2ysQuFiHWB4YNkvlcyxK
RNlJMmIL3Vw8dG2c2P8+lG+p6sp3VMPUXZA/wfU4hir1S6GVqv+InbpB8rwvnug5
GZCkpoe+9jFCgCiErONbnxpfvkbZqP5mtRxVhuA5FRJ5apuQz4IEY9b0TtXn0vKG
o8iKWAX2y7EFxhR4t9uUPeytT1/jQ6UwLV9jDE9vC5TGa6AG5/2PtXej50giLbdE
6YpH0Ew308R8hMP4kyEkAt1sEUdSCoWQfPxlOyrDkxxT14Ffc6KhYLwD8t5sg9I0
UbV7eWG15qv7J+GM9Y+6O7I5J+ROMO4i9NxKbbrJzspXYTtkG0PKXukKLQy9sN/x
6FItuMmcmxmgirjA9NGPw0YNPgwvVHnwZZVIr3O2wvLCBbt9jw8zFwqauv09N7qy
+wZhnD7pyxOpDN/QQdOa6Rb+xLdoLrr5Njun+wlto4jjB9NPnMSJXQJq3lk+jJ6p
pA2Z//gNCKzjXwr40UHHm6zdx1GS5Gf9QFJLvw0a9vrCzfKjx9PYTSO4sry7rH5X
O001DtVYh+MmZlH/FJ/OumG8B1OTa780MkpYmrxvgQfD4l043Y36YmQOnFXZWTEw
TctUskYQk/EJ8nESKwC6QKTZ0bq6e2y/ZgPNFOKZBDcW67taJIqxkqK3qdgZxBUH
QCoEthN/dNh480DKOWM7skE6VwXibjBNgDThWwCybKIdjEVuMLskmCG8KXJbZSNY
9ebOCjNwE9yx+TozsYyl+QYFXRjEQ32gmXidS6W/FQjM0atIcVrQ0Xa+FI2Ow+Ra
PHWsfhCGzVgQfG+bJbe3m90umY2CO+/E5JGPKo5nphk1V1cvCDFCvm9GLBMWIEqQ
xIVud8tox6YwqZrcSxHOZjyivDPEyonjm1kTDOpfussohtb4kIkaozcA2AehMSiD
yY0iQtZ0umUAiSRTci8pRbtnzlrU3qT1wKeGL48jNKo1N+qw19yL0Yf52FiTmUrm
KaaGGxoOk59ybxH16HPFeFloC+OAzH23Efzid7ekxWCSLOFLniQOY/Vpjxp91drs
vJ4Yoi1ALHGNlZa6ptjssQK/TZ0g3q8MeTA9dKBTZ0qo4tpvJFIsWUAKC9tIobVV
AQ4+dg10t+EudWk1FxRz5gQZkvvnHizTc14QmwxRQgX10EObS30xCM5vfAeGbaR1
dtKUoiW5emHZTQY5Ou9mV1v18QJ2/7adxkLCws6jifk6ZTsxRM3bUQxctBA+ml1P
ahzlre7HOo9dwEAvS5gHlSfuxarClQCg8hvLBEykpUQmA3skj3feGIWbePLZ2913
8YSBcInbMqqS8Uj3LoJ27eDZ+6LEiQ5043mphbXiS51670QAhwdwxS4rGSl72+ar
ihXRUw/9cJUyyK6K6ACKJcvtMSKAl7H++JHKluj6CA430wjSXtzK18AtvOQfH3Fd
XWA0Q9qv+WPSBgHlK8ov3EuX9Yv3jbaHd2Q1rdFvsQtk3Y8xKmrF+CnUJhKE0XQz
i67VlLjIJHXH0X+taOlS6cpNd2xD8f2zUUfrETjl/jkRXyB8QNDJaNOYNI6EDikB
T1ov5dDWVwdAVvLxD4iHYfWx8kpGhDo4Bsa1gvlzFDQ+HxSOxsU976/+BWUUHKJz
jrCO3HjwCipT6rpIm9drWLpshFpQaLZwY7TwUNayuE1UqqHdIKV8534ZdU/rvK3B
iiNLgLc34l/265GDtfgT/UgvbywEDcMnKMRWi7dD76ukdtyYcbkJZ8ZR1ao54jr2
UXxyi1Y2eDZqTml6DFGudnzDTufjvYXphTHGFhTi7dJlb2G83QitfrmbS5bl07/T
qvaMv570+pbFz6iybCUzOrSvSxfolekzBkibOPYTzcxOEE0/tbOERlT6IgFsIiyF
MSEPVvhkOYAezROBkM2wkrH1OMMpvt8kkvvf0k4PLQqkQmcWuzGQOhX/Ov/otf8f
G7CThobWlmizDYmQQnS5D7HhRvE8yReXyUpFubw2hQwfGkFi2jaFtwbGscL/Kkn/
wxxs39wu16VX3FVae9TzWSyRGt8Mtg9m+uw5hMMvvgE8k4AmNOaJKBqWda1QjAKz
i5POf45fVCko0jVzYeXJDQzZ8Es+on+g2NejUdd6Onckl39zQdF8TxzwfvoTAlZP
y9xJ6xSBzyd0fwxWH7vgwqqNYG5x8LwPqFJ6xYLYLzen11vSQ5g0DRpCs0D9BlVN
ziQN2hYSolhHXUa3iFWm+LplQf1GYXAIIx9wH/BhCHRZAxCK+4xh0R2UDMjGGzVj
aJ9nfJxNvrPZ9Z0dQGb+q7OfkkIN4WZXigb0UlZ6U78eW5FBvASMDdMuIWHO3WrD
MrLMbCNZQ7OHFjA0mcKnP5SNVCo1aUDViPBwn6Wnitgo18PQLY/ubvbqYE4lqftt
o0OqrMKjcb2/SwQVFLaoXgEVSJPPI/o4YhZFunUCGN+mPqFZGM859UUzOyg2YKgF
BEEOINbPb9wiLcrdbmCyYCt+7U3u4kRTfIl+oUCeKZsJcg+vo0k5ZD08rcPxCbOc
9MGJddqSeUPUMzpEvnLMDas9p6xvrqE4y723at5sui1AjMe4mPlP6dbLe5dkiata
vSc2zrGFEUREOif539SAcM13rBtRxXGdSwmnVXV1iu8eflmurPOrA8A2nfBnAXh8
M8sGkeOdNLNIjx+FV2lys21vJDzYW9fUUnppdU3CQa4tqSFeeOtRFlvbMAAkGfaZ
N+coKbPn6J2e57WGznByi0VdJ6dPwUY6JOds5Xy6G4lxlsSxZ52JciEdv0+xud0I
HK5iE7HPVsTm841DRqfrHwhAt235KHRpbaHQisOH8AryOOwnos4L90vu7cdAkbAR
ahTQB7ANIJTUfP4Vba5TanzROeun5Y52srSkL+CfwYFk4UmtEZXlXyxV9ug+KOye
tnAd/Wyakaxh6Fy20ZU2vp7G7O7dOeyGOwGkBFp1bZZKVuQVfdcniPFoYJ2irnET
joph0/n15v2rMpA2qeeLUEPw/4o15HVBAmyyLQspZ1w6jJJ+SBM5PB0rAIPIlNR0
Zwxzp5R99G2BoOSaGMXMBirERZQD0icQjJjmPseULXl91qgps6I/5XnKPIAnwR4/
V2hnblS5QlrvNoDQCvn4dyDtdvKX6a7WhBdGSsu18Ol5s4oqpVCvuASC5Q5b0pfd
KFRjwxGD99YjgdfvsLc1WbqcoQBnIADWBfMUxAkjRswmCWdFRYV92XbXxdrm8j+z
lLngu75MS+8VF+MJGl7OReIgC/xb7q96XOlFQp/dWdOn2QEhd++/fgq1mNBbpJgb
xxFipaHg/WDB2AQn5N28HdMpq3HtLQkh0fslKyYQ9RBcMdgDFrdBgNISq/FoQhdb
Qhu3FB5l79MvfC7Efh8MrdpagrX4aYsJ1kIHMWsO+XZZLLqC5x/8er7rtaNUkYep
CPhTA35sH3T1WnL0X9ryzvmarM/RfoTz+Z8bTAZKpfrUeH3jbBAENZPVLoe0N9AC
3bquhpAYZKhHUK0bXKdif/j7ZxuPtELEcFjDoZxr1NmTxQIXgindfMs8ZEMXpe6e
KpiwXiLJxRlNDjIRPqNyFv0K2sMDE44XO+54Hoze9y3QcGJ3FReDWwNdgKZpY+lq
D6sGasnQ1K8zVJBgBBEZdcOAdt0qcq90SzKrG8Bct7Aq3ZwFRXfn8t38Ek6X4qX0
bz4RcAkUNsQ9J5N2c6aOxdFM7eBaqE9T1GgaWaQF8aPBHPG5BcAbRiKtKFJevOMT
QVQ4ApKC0rvVI/RsgD9+oCfsjdMBorLZD1nv6ymurlDYRxil0iI5xVS6FTIkhYx6
jb7H33DhI+aBfwfDDHitC4oKsZ02aNmzww9Ebh5sHG7+yXUyTSPx7vQRkal17tLf
ARq3WPCwnAjDa/ON41rMvAJUNUL80Ws8Fn/ImqmzAAUYqHPysMF1D1UHAhlqO7Nq
U6Vvc3H4NBLH2LjG031JiW8BmYcfNfmiHlkBIbPYYO6prqjkjl9xINBkaHuLePGY
j1/XSH4nOvMH3y82AWaxGGVzFNklXaE5m/XUJ3DDrJXsQfhcilMmja7eF4ikcx8c
uDg7g+eBK8KwRHBn8pS3vipW2ZacbYYQsHryZ49tVdgSP44Ib+MkaDd8N0LwzCQW
ZZvCBtU+ncr+RgJ95qmnruNQfNMIoW5ca40CYY+E9VLamGy4wqoPjYbHzF452kuB
Cq2N78rjW0FrMFG5+mJQBbxnShOrwYEWLg5L/zihddS/WBSD29zEPoNxoOqILd7C
eM41Wxt8j5DJlVPkdam9AWlcQesHlgGhTx5K0WuL3rzUADarzF0itQh/cWJKSDCN
AKRlPnY9EiA4ssl11LGpCIdLd+6VSiFLONV9qHzEZm9wtXH/AXp1kSAHFruJYGaP
6dbswx3a2jo+yk8Zn+HKU6zQQL4oakbzyJi4aDXQvMtyO5cGcgKLYYRw/QOm4Ec8
el77/6oJV4Q+oKA3rUTWpptwcDhtHddt/MkRBAoI7L2BeeJLsNX5ee45IhOG0PXN
Z3jAC4ah2Wdc9sCCT51kt9l61Sf6SkkuI6wFTDzv/FP3/j9KguBEGKkEshe3duRb
2qvJ4zQL8tmrKucHmJjJkYzPMA0rZqa+252fBih+s+xaOlcVFOjKx6awdZU2Ckda
UHkEYdgrBMjx1Ic4zzbo470za9QJY+bgktc1DnTbh2MxRDU7ED3VHn4CgNzYMDbY
/YqFZF/0/HCa06akWhiZYeGyzd36+0a2JcmXuQugISUEnoOU+AZ/ec2c79F7Gir+
+l5T2Vn9b2WljSc1fWi1lbsjhyN/CQhwrPpnFdsh/dq7JPo9k2Ubjq0eOeI3abuG
OGhGgd96pLElWT3EphBKDSUXAJWBnZ2OgBjKwdRuVpim9Z5TS+UW66upcaKzCE7U
YNP3LKSs0ZmLw5LV5VzQA0X9U5nrvYcSPf776b9gfBfbw4Q9tODCpxKZuhqadPI4
sQTC1P8opbnXXkgX7Jny7/h1Nwht7rtDHskszhOW+mbdIPck3ENOoSd+LlolTYlB
jgtKrjv6/pikHo0vnufruNg/ewfQCGK8brEXkqbKTlI00LCz1B3220ktOXUd6tgK
ap0eMK5sWqC0HYNODlcgU8N8LwASXDN/DWGcgx9lkhM3FumNGz3BDeCYiiTc1l0w
KhseUyu/+NkO+yQGimtsvN7oyuveXAmBwM9CBeW0eVWzHXhUXMTvgda34/b6AIhn
WieIEUq9GplnHQ8lOXNRCOjOlsFezcBI1NVP7L+b+1PgEvxJ2y0sRhbUFcv54x/m
DuvjEjUKPS+wfjUoxLfgnTJ0zaANoJWKQkWi1y3ktEf+klUfKLB3vYKHr0ktKo8O
Cb3/DbXPQNn/MJrqmUvFl9LCbEm3a95G+y8p2/sPYNH2EKytYKdAtNMRPsNj5d2y
JqPCeocryNs2SiNTt4dLwN9PwqINLYRDD9YPJx30rXZXjXU7mj898BZynpaOaZDb
5Vpjw0dXZ2q9xZ4KislnT2ng+qZB+ck6k+Wde8lA5ikTqgtShua0YdEcgLZdQK2p
9L0Tw+QkqOLOmv95ZcnrTODwMETTtZUf7Q3YP2QzoOR5lT7jG9D5Od1SgKtlPoWB
ywMR4EoXLUaZ/2fXtWMNDRX+M7g7aLwikY8Yc/YHD8OhRN+MjqQdufG6utfBJDHc
64ARpqFYjpyGxMDyrroEoxHUeHWJlYgKoXkZCxSJRxgiLi+Ut9BT+aAvWNQ5dE1j
drTuptJ4Mk7Vp8Oism/3/RORxDCBXdU8KMQnbJSZv2sdry1vp41bCRfoQmT8OCWk
yYggHvGln0ST+YvJFkEwKwqJa5t0rc7H7ZMoR9TEawj7hmaVCylQMC8lMbS0N6Eh
8e49ym5ahgvDxMp1hSIL3l8Tq8KONihsCPb13a6dTFH5ui48SROKdZdgS9EwTwz4
GwZvhD8uD1rJm96mCJ2PPyfP30M9ZG0sIkK1Jn3JxKcx6044p72TNMzRtJEgVEkR
gTplBcujcZ3tmaV9b3BlfUh3ww0YbxNMmQoRuigoXLsqlHYzT+OXAtWchaKTnPX0
E8h6i0AT/j1AonFi1TFtpop5YvuRzPEUInH4F9V32zbos9R0pWjNF6vuJlx2+WTj
nZAPGdfPC0DcYA9FT0KrRJ8p9YyOaw23zxly/P6PFd0Skzh1BLpASaYARqa1pMgo
i3e5x3WeThQlZbVfL53WhsBuIvPwhpCxvnR1JM6WPIVmNyClep6f530f4is/guBL
FGv1N50UgRoEE4XAqBfziDF1YTpeEESxA3Xg9ZEME+IjiWWoDvTldr0M7UlQjs7K
Kg9xnmxpq6CkbbIbll4j+USlR3Sy6gag/1l8qmYsY9r+6JxLdxZsnlgHynJw9ddr
OotXtmUXP7ZHgD5lbxPWO1Mg/rFiYxM+qtV5mIjJUe9hreRc9WUW+MftkmtPFoIu
TlErotvdDF9Vwu9mtAdnP6MUjL5uXzM+tu5BhE1GxSkxspDPtGY3r8wa2I/Q8VSs
Epq272XOoM9UjPjvuDWjKaayzZCqgHN83S7tS4HBc1WTBzgs2AgY0N2IBKg2voOE
7OIHqysAM/M3GXsTDFz4l+YFLbMLB1cwFC12mkPdPPzgCz7QOEq5VHJvCL0tD4me
BLH7qBZ2FkL6Y40ttAhZ97/3ekaLu6X9OAKk0lYSO/J2AGr++ssTel4kC1SJ7lNc
CVVaWOx4QsbfDNjY8R3/SYZEDSnp6RX1kRMdRumCEbiUtHXx3T+Y7MEKyt/FWVPV
y22OvS/tXu7nVMAgquFLzyuQKJIdcvy+cvp06/0ysqbugBhuoG8B8bCfjjGggi6k
Wua3b+QJdweqMuYxlsAvtUziGRMz6qHM5uQ3NNF3aK/5dzdneiOIXC/2vYX3r2mr
cCl0lfcpxMpdX6Q4VAEMKJkSMGBdgJ71O/g0GiyAvY/9ZPFQ6HKzzRhtNNCKvERJ
dsIQz4w6eucXUtMWVEbdwwIBfwxLwBLm6qsvMcoxL9CO3/aar9Iog9kORPpgqV50
/yY9zMaEZxL0J6ESo5JpfTdUjsicsHb0cQbCIr1Uh6oL53EoLY6NCDwsvsiF37Fa
hIAu83JtopuxugFQ0Am9NsamwNET02T21lrJYpnxHSWoG1NkCGgfD+10xzcIzjf8
jZs4OmrFn8Zaa+u2Fz+Q7EkA15vGIDOQFUw4T81l96sfRJkzsiSqHfNEkE92Mn2P
R3XygqeDy6bu4LVdkybFoKPVV6bB34gjkl2N2eCfyBFmLa2YCGR7GpfuYbwDgdd4
9tA0jhIN3gxPiCkMi4/QE7s5XlPttcqBP/doGl6Z/m1dqCYh0+XHiQK5yT1ULyK4
/HH5cQe2rRsMXpJOMJRonxxBlL4fNI0SCs8KX1zRKaHZWhquucieINJu6gB21hgM
W9aDdaPIg8au775kFpbHS/nna/V/SYTkCxcAygUo2sSPEO197ofPuGP5Ke4oyuam
+kXw8Dhj3uFhIveirFoNgAMJR3jjlKNej99RMkF8rR6RgvNXSFk9X1Eztt61CMxl
Ejm905zl4/uOcgoMiB6bZGaEtnOWDEoSFUl+F6H/jx5SfoMApmIjZ6A0gekmaixH
EOq/SL2ErVkkgbjk0T9DF2+7a0g7auo3xNkpmN4ZTSXtndy1pk9BcuS+jKm4Wk2t
dhROVnQ9+jOAckHqnpYoGPaB7pV144y98JT+YFqLE5c6YJ2/lmmvQ/2EVW7M0BoD
jLDN/1toGfGjley3bFuK54lfTWMKYu3bcGCw/SVHCwLp7wxp67Y4Scj6cinj2uLF
NZ1bEDEJZm4Mrr6LFE8MP5r/OPAdZPcXE5w9f9Vpomo/qQwRbUz6OB8gnkrkPCGY
zJTVHX6lbH7gg1N5Z57mIFDSpcg1EGJpn44NEwW5xPEvOEF0FqYtu9RkSBLQHKcE
eZtodJ09MaImnQTVzroJfQ8/szTZxI4TNJo8wInIzULDJ6KTYzjrOSNXZmUOdQaD
Wx3Ix1crSeD6axVHCRIIqDqdfbQjCwWPMkIY+/+CULYLFlS55qfT4cCyfBy8y9Al
Bth7k1Uhp+ZUwHHza0+UgS5ONVuePuNlnyXSKJdW69T6PH7i2V/yz/bdPku1nmzJ
Ew3oJHBiWk8HkCX/tKJLbwQ2CpdltSjpRSizh2rvZau/7DixaThS9dza5J/5OfIU
Bc+28iKVtSi6e5FGExYHeCxLIYMj9lI9Ux96yNLnF2g/bblrka6e9UHJQannG+Cm
FUG6VjHs8ENEXOEeIdxVvoZM8SOOik5sFyoA3T7kcR/0Jp1YcDl0TyFkp5jRlBBX
ogt0qiluRhSATINMn42ViuZzkLODMOiXkd7gAuUQTvHegaRmfyzPvP4kMm7lJEpM
9fHXkVV22V7DmnBzEdPZibNOG+Uvl/XDwpuxcbdA95d1OpZHbopWz8bor9JkoJ7L
/YPuH2qWuTJD3wbGD61o4nHZLl0Alm010KmcDBJQHKXVGVD9gbCQQxx1fHiiWwx2
nPcn1nM0tK4wAhlkUG3yZ/fVdGCFB0cstPc6/gMixoZEALJW538vvpaawX3PVMGo
lceCd6a15uimRAUcRTYZHqUynkOYIhzzFnEnlGJ6TorENkmAgczAEPj1UmIkWamm
JGrfrfNFbJAgTc8V3fnvkmS2ENJLnYzyyZiTBHEI0weoE67dvHyi9VINFJknVX5o
hVapCBrYDg8N+ak9LGBdbn69T75vlpEV73iG6cwSzZHuWopyqvPNfVeXhaSo+mAV
3Gd4gzg4f8/dnEj+/uHNsWaZS3TMcxbT1csoBhwW9QWfbPLiMHH1UJAGjMxZWK0N
hy7DyznU8nrDdTxBEpxfp7VL5qqRYgncLN2BbpTPfOmmOQF0ZT7cGSbFe9B2Y6hl
QNZBF6DlH2pWdKOnGMSvBzA4s9tpj7Bozp101eDU8j1O2E7Tr+La5TEapOIL/elm
36fcncLuPuFqGCkDRl/x80KU1Ow9+sgOPA4xesWMYoKg4F/e83b7l4AgTSXA/HF9
jLMd0zbDxQhozXOGH6gkBT93UMdTz6Adf0kqKjdOzxJUivUpgEyPfz3AtTZwQ6Sl
62nsP0VO6NnUaWHNLFIcPHKTZbiV8V4Xgx/qdeuqJtSy7VUEhuUm5L56Py32bwUT
2iAXZRdVUhWyL35tVSMBpfr7jFfJuKBGHVON8i2SDh5yHGNWam+jgqnrwaUvI1Gl
e+cwtAQD0BnrmJz4JpcP7UmaAOaBLZQkxsK7AFRlPh/w+VB9pASg7gNFq/5w9CpQ
lxitPXU/Yfw5a2MqCos9KLhoB8dlPS2WxmCDvE9GfaXIztQyIwNFo6ZhJBocgT3o
fI4KhjREzPYB7QPqaZuVPmDPvm0T/DardYb0o0raBlI48cmJGM1R5x/es1JRnK7Y
iiUjcGztpPffpQTxdq8S42UznHqbQKHwjGwFHqg0VfGLcjfm6b98xpQfE5UISykD
dlEABoDtfllDVjj/5C/pixwuVkKcUKnOZFZxFI5uuj1yVTbQWzUjOIzNnMpRr+bN
SqEEdO6bn5c4shvWK/CJlwZvBXd+okV4sTcQndZAvK3iGJH7fsuB9A5jqZ+zrUZd
dFeWzD7Ax6BtThA67CjDOz3RiqOPQGm5Qe++PGRiWmIl9MfMgvM6sTONYAneX+vM
e1G2vjiKufBw2lrJVLzpb55KlYEqNh+VS87TPWhu3XMYMO5QGoNZCZhB1K9o1rJz
8Dn4FAdHvdZL0gIQ5PJ4lNKgFOnTBJjf86R2YV8d6keq8vNl8Lm4sjPfnsIiwAz3
NBZhXTFxKGU5Syst0BhThOqeCCuLGTz51CXriFigrkNwgdlpGaSR59+Z9L0QPCfE
V3qi+qZo1oi8GlSbni4vDVc5CNSd2Ah2gJ7SYQNhf1S6RoD1hvbbNBCdQLZz0lxH
nf4EkcsKVTTUD3LBFWcJeWW1cvBYmidOqT/BTINj0YLRHCLdGCatt285F3enKjmL
D/F8lzSSbmRDi5TNnNXtDI0uxBP9Ncoh28y6w8YBDVfWDONF7a4f0S4B1xs3lJ3i
X5dug+WdVTeKeW8rvBmqB4RYiVTTySIltTzVuPKJwFNfwAyA205/FB9XvWbplbC1
XGJlxaRP06WChlUxmHC+QWCXtxjsDzNuBWVD99EJOJljEKI+cCK8+5LY+HVpmn4k
QCZ/p7uF2Ldd3NLXtjvbwYy4Tv3rQ79JHrcXXV15dCooii3wSNjVAcF64uARPzAN
G6Sll8QGGLBsNs5uGol2I6krQeTffkyKjTGngbn1pDDwCkSTXnC6gO+V4swqmrg5
Wte4O3OMsPC90u6pZ2dfuqUX/G+XThSSpqK2NW6MLob3iHqrN9MWzdYVECwWJ3kf
wBNvRxJVJXaGbJyrrwQHwjbtusGVcJJ6UvwgvHxBtqoaGstlBYyB+rKjFsoggYp8
nONPdfp3ErgvqPxwAiJ928ROSvjeBOX6aIZjK1vDUUxlnN02awO95GTg+4MjfKSh
007zPkfP4nLWUFGe+Ji1IivfKiNY4xRyf7JEcnZjm4eqpMYdSuMsVetpi6O1Vraz
ITAC8731BBwJEGey7rXuOOdCIFgGUE9zxJ+hWgSW6n9U0nL739N1Wt3bP99TmK+3
iz2SoZ78gtdBu1M4G3a+P4/Qxwd3huk+SzPG+h5EY/IoJ8ppBzyKzVGfw/k0hiIq
T64W2hp0aBRI7c5Qbg3YPHJ24Jq6cVVWXfEPyNjH5+08stw2D1kfjLt17pXKU2c2
3hRDagQorluFRK2P9+3q4LUjEa/BTZ6DZAtIiijzfIy1Xgn8fuIpBwBVlIagfi0R
igjlRvjqnLH4+pvnirp/gpVMtcsl7EEAKtTOSLIQAY3wVLGCrvMizb5UNZye9hN5
f/OYOKOd3c1l70P1hBFx9ffolCnpZ6MrhZkuuigNSnfXroTvfuJePH/sc5JQjXnl
BXT6j387TU9c2sklt+yi4GMcTpNDehS+kx9pvPkfa99EvFbbYJHjTqWe7jsiVArY
f6xSxteXSj8l/xYqxJCG1qch1x97eQqC5p5gyPISCrFmorr9v78Z89k922OfuSqw
k6eqloFJPCMK/oNzxJhHoL8qJlPlWuCbbJnLNHgR5DSdw78HiR9Hs0p+Sg84/3oG
xuDfO+Nswo+3u1doHDHzceXxFGiOte64JpDESQtsqyFlkX7UPsy9/+7CktZSsdeX
rZHZg9b4TV0aDBgHyfEZ/p1Uc4116Oc0VUDIhUS6s91/LPjykNAVQf+WUr3U2rXv
LP4jjZseSS5ca72eIZQMsmUJ8uxn3SV1VhoXp5FUsrL3llZI6Lt6gAs+ZIEjnImT
97AJ8KC8mkTOGl1qICNJ2vAOsgQ6cYa+cp8/KVljoxQdyVPHMttfprpH3fo1q1Ed
OuhYEpkZwiSR/CDKYSBuYH/jSmviDVOO11Fjjfzii7Yr0sBjHBRFUAy20nFNibJf
ti6qvUrFYged9MJzLtN0MFpvb3wqTMmf+HHRKjzA99w4/KeV5SnNGDGOVy+N3t1l
2qdbq8oh4hIQzVvAJU3bDHTLQxapUaLz3dWQmxHsfGW+yboBEHD9zQMBYO16D00X
qsV4w1PqhkKGfmmLa/r9Z7mXocixkEuF+M4qsMFuC3FAzccAiNvFWCMe6QrBl+B4
FFMyrBu0CzIzD9mSDKWULxyZlvU4Ybg6cnPUffA7k/TFM8L8x//yRWJYd+5teQrt
ulssZlNHpRX87dU6/ieqiey0RD96qyLvTBXsSgWtU5MEX22WR3jIO5eLXhLVExBL
QzhUwtTvCvVqAM2avcSAvG+RlbdCfSx6CG9GQjtJY6pSovEZmijgmoTDITPJKsbI
CmUxUzFAbhzMrht38xMWMkM5hR5qHJcBDdJJrfuaQWiLYNloBwv0wOJxQWfxwOjc
2PNNwbIuYfGoGVzDuwsIAKYrSXIhohxQZvrdB15rfB2pawfiXcRkEdBrpSpo1ab+
+bPQx3XBbY2ihXumypZ8JmrsOJAw/API9r9ZXYH1QJ7V6DziMRVETO4NAokxVRUx
8UY3uQo5Vl1C12PlpvtJvWnlbh0T8uNZiP45dEFGgQia4gzIfajysglcHQwOwupw
1bC3bJtu2oR9z+MI/h4Tmogrq9H1Vj0JDfAdaxCW0FL5uHn3kLxzEH5Xj9XIcVNJ
lCqBLvyxXnHjl7QT2Je16QnQdRX4ZAsQCO+l2jmm7+k0Hh+T1lGp4yoY5EB6vqJQ
KYJgXDTY8hKKopTLsSmDf/3h5XwsxnFb8x8q1PCIxl9Qnros3IoASA1eSaRdYnwX
hW/4CHdKNPPl1ZMs+ndI8kT2nD7uA+tJmtn/AxcrjYA5Y0fTxD9occVn+nuwu9V4
0nm3oloJ3gUyhz0985jMAZxgLrBkVHfPRnQEamtG85Dvu6B2o2GOY95jMpj1W5QR
Bx9YHTpzl9aRn0s8m59yjH5KsN1tOYOQbhNnkORnOKuFeL2IWfGpo64DjLGnJu+O
Cqg0Ejud9eHypdQJ1Ee8ZQnwTeN4JpyeH32uophQ9Z9J1C9mnKFW/7rY1t1FPu/r
oK2HzrZnNFQBHtO4ziu4bhQPkGyus4z9MMNDgd6dK+shZQ7XMRLvAVSfEgwMuoSM
y22UyOVOLJ42cxXxbGA47kXFTo61rpsRbzI3tqYnfrtRPZAQ6nqF2juz+oJkJ/aI
bcLO2wfwy2tBY4dsjsHfTlH14uSOzNLzQryEypWwZutgVTtJoSsjMiPYvbY4cyUF
w34kVFSZ1yyslYxyFrOjtTEvfyDj3e+1YLxlK8valUTYLEkMjAC5qxYsPQR8rkQm
UD5z48IYlx3PPvd2VoO3QrV6jy3pgz2JCnhUNyHhDkLoCbJgloU7iWzgmpY56fZ4
kpLK9DmjU5Vwl2FCWgax/SaNCn2cU0tDHwpbws8iysT035tNJVQfJu7BRpNwo4gA
8gS3FPzZzusRDAz5vT/naa+yhm4JkqiT7W8bcLlsfGAceZTmeKUd/59aWZzvZUDF
Q1TJx65ExdR5qvy9tBTOCFMFFiWfnIWjGSpWV4gC/HSGVi9VjSjJgc4SjQWg3gz4
Nx67YN4Rmqpxl4TwhasWHt/VRgY3H4DhnvrWp1aGfl3v3Iyho5kXPMIWcq/9spTW
oeh7DsoQykgBHVoQFrL/t75rBz9Ns8XpL3gAwy4WaRvAFZM1aivCd3rG6xb9Nayg
FTXKGqaterE8j6voPbZ8T77vWajpZJ5D1oyX0z25kwDadIq8zcpUSvTYJ1V3zTIJ
7dx2PHGfuItawGhZ/rfXQJ5iTG9vqGOdiN8OIXAqbP2Wqn/KX75wfjsp/8q6Glwk
z0QY0ikhVj+OZjzwb0onqpSelMGPbKHCIA6d9ogCZyYZHOucifwTORmxfpkjYa8K
4016ixhciut3Vov4vwsFoxKeDHkuMcyj4EEnSOAfD0U5mwpyEfrsdQXSv6oWUGHN
dYNvgAUa+ekcyiUYFHNMmP/Ky+2l2M1hAe+PMIEPlvwMSmRQXJIb+7Lj0ewBPxqR
RQNRW18HX2enPTvL0BFQ262H7w/XFBiR+vJ8QncW0rkmwZnqkkz88anSEM4onxQu
N3AVdCmzpusDehFxhZ6eqi5hUobHW1A2Os8823gLTx2Ao3G4/t74EjNxafANj5mv
ofxeoZQSX2CKgMOgVtRE1O3urZWz1W9m81jMfagL/gNH5RZu47kC3FAhA4Aye49z
AZnAbewDlU5W51tUiEz/LQWRpKwXjw1FJxqOOkpKYKEwtJ/9zTEDJ4B+sYkcxrYV
QFIDPXQK3IvXDl/1Wuib/T01Ni7oDSV/4ifn74N8oU5BqCvoTSB72mRIZ5ISV1ed
b7yob+BY8crX+OrpXYpN1w9mMgv3iszR9Kia9pkzJ0mFSafczGGO1yIC/CdM9tWw
w2AozN1oDkyRGV5Z1kFHN8c+zkfLvjHoiRQgaTu18PRuMIsKkJ9SqcLykCFuCswV
oxTxf0AF5GD++vb775zTu2aK9Nc2tQFXpvh/X2jIzkVsz9rFgv3iAz+kQ66hWZ5p
XxkTvIdeaLLvWaOo933Qy94L+ITcAkbVb03wQTid2mQ6ep3ayiqHEtgdN1soAIem
nfOaDZb3BcVMNgAH/DG0+xlJqlW5hyaH6hoXuJkLT4H0MWiopVR7Tl7L6iDTVDwb
jQiiN6Zz4mLDgnE7UWoITQlarzIrz7tCtT7q/BmJjCt8f6F/9rVVh/NkaMSGDvRd
CLcBrvj0R/dnq5IRUbAqaO2lgA1Qzq7B3x8EYONeDZsaSi7coc7RlZbGjllPLGax
qRi4qCs/c7Axwesj51N+cseHR7R+IzZjChb3cBNswWFHqM8xlJt+2ces4SeDPwcC
pe/ejfOPaPxBnE3NIJzQYWaZqF8jnxfHvcUYFFaG/uMvdEld9HpGrDmaAeqGf3rL
6/mk/3ecPN3vVfsYQ9ZPDuwY258kRy0A58OLQGsFxkwPDNUUyBXGHs68KIHGk8Nu
GZqANoAiZS0hVmZHNMPIfVyEZlow5kf2yyuQR6+VtsX4Rik05HI1uGdcEGoA/JT5
t1rc5EQRBb9d0y+zymNRbBx7kFYjJOcKuFhuLLIRCwmbLBJTe0T0sO5A6Z7R5Umg
9MmKofCq7PeJqGIMZZMklH4ovCJDhhVv3J9mJzb2AVjmW33OiiaMuoL7fq0fMrBw
19+PKiwasPkHWusaLHkuq95lYoAHci96ww0dbEW3X+1ykA4EghvOwoR8e99MzaIO
PQn2mjyfPzr2EWvIOSBLNh9Q814FF0BhEfwawxFtoXG+a0ihO04xhirxfDxQTzaR
rtAQqk1bn1tQKATgq9OgF+NUbr+pVdbtY4gXqGaWB3P2GhSuSDc/3E3NC1Ij8WQ4
+SZrta2N8V3NYgy8tIDtSW69lFX8bUxzqVg6mDEXuIiJf7RKJ8jtA/+b8OEOBeWS
NiPvjhlaNvk91pFztGhil6tTnwN6evRPNCs6ICm3fcLcK1XKYguiG0hyJpCCZ7Gq
Nw6d4x6RRWv3Pld5LhfHEmpOJNPrxQutINk/Ilo7rsH7dX+Fa8lTnYgM8Dcamyjg
mJ4fuzbNUx6ufVI+Lk6zp82wmYk0gj9St2IBf5wuQRT3RDwXVdesvweQDce4iL1Q
+b+W59kwitXrbbsflCR7ZNOTn+ho8uvaiAUctk0I2fsnvG+xEVjhnjoyTiscs/rh
Td6y1ApN4EBDb4P80bmmookZGscpM4dz59g6zn/65e0yGOwwRSU26QiIPBZM9FWH
adrSQL1ngZBCuHDeS+F9kUO9yFRBzn9exoC+ZVWuqQ4NU9H8JhohSmQ/v9yXouGw
re+26ARUpkVgBw02GB5UVrQSWmRZDRSnwZfgKO+bWt/SthOBSTv1T+hBbqfriAJa
aKX7pX/p9MCjM7PoP6Io3ZzHMLMw4IDD7tHCrmlElVpnWb7QlpbtCBhBIAhlTpAz
eVRuQyd2kGDIPjTHUhzVRbDRUNK1KAUFWpKDhv0u5xX2kUb1hpAW7pgC9EZsF8d4
VYYJFU5GYewtpVLIK1TC6RicrmSGwnTFN5LP1nu+ZRIcgG6aQ+f/KcXvxtriRvyD
pLSUOA3T64GNSg8zJVAXiFHmq8OpYSBkQ4MC1qOpB7tes2leFhwOJy9I4ValINxw
5TKX1QUD8l71M8yA+3blToGS8bTnrlA2k41NjnAmoBYQ2h2OIEGA8JVHMtkgtZol
G/cnqdd/LMPHR1WtJHbjSNEqorlYHMeyjWH3OlkzBNUNkgPPSH2RvHLzOK+rzEdh
P4eLaLd5dgWgzWFmpW+JH2byKWrrKGypvpHw3XjaQFeiS5BbGirrrwqGS7epKHfu
keRexSe0Yo6zFVAJTC8LMaUWRsTxBrlGjI8vvyFrJ76sJakxY1qhD4WQcqsKyTVK
0XIPWq1yt4ssIASEy0x0vNP47NfCjH2NQR99gyH6fxFb5rpz88NJ/Qo/R85qAqpq
AUnwwtfKcDOIBNOHM4G/zpk16dM0dsbTRUbUB9bKezhbLByB6GuAJ+xtlrGJ90FN
ybrxV98LIvvy3AWUCJq5IOShle3+YW7APqMuXTi8uupwhRKuXv38DF3nhn2hQNVz
qfUAsbfLo8/gpgZc8bagWGhubpno9AjsA3zdIliMmlcqK35T50qQPkx9uZ2Qc7cC
ZbobSbpZyQzU4djHJRoAim7wrJqLsTV2wnc+1x+n94zBkGnfIx6BJGiaoQLDzNg4
VLKhtQQ4IooP/W+NHBuswFbu7q0Z8eeIQ5UHvZEFQhm6D0HmjW/3bQjisaZ8N6Vz
rTybWFzXDfs7j0ArdsiQ5SRg9hrD3L1KqUWqK5+zRgWgxhQOduJ32bXARtYxLL2i
vLZJqvSg4m07lt3l5FOBXCYFw57li2emkA2/ZJ+ErNXsai+H1utqxXG5Wqp6EjRO
xm8EpqoVge9LmdgkH3M0xHdxoX01zEieJtLuA9CmogqLpZ8ZKwkeZWt1EyHIvuTc
hYLDww6XPGWB42q1MR8uBLEHpekrqw5Ch41/LrJGlwY3O4FZXtoeY2qu9Xz/vtpL
59TJ1hGTJWWHAADujzNSiY7mlj2iKxOLIcMvGVMOcLxmwVKSzhxbhc1dSpBTXM15
f6yejFy7vLcuJMjwJ8cWcDmRS3rzccd6fwLx+mhRPwYUoMduNuZTg5SGre+8gqlR
gYkw4Q1le6VTkn/ZIl3pkyAgOwEerzYTbB18U7sjD+gjaajLx9oGo7lP+lqGQ/Ck
7ZVfsDYfYKUfLYvB3B+CB8qq8hwRqudPLWWtkihn+CvL5gqjgwh8GpW41K8GQs7Y
jp5dBusZpfdNJXKO52h1ZleMl5AALamIfpmFtOc0frBw81xH19mYrcNWSwWtCclk
xl8cKG4DT9TVF+NIdlsek6H8ndcLfvIzdWAJJPcQcYVWhX8YWDQEd+hyckkKSZly
jlxKIrwoO1zbMcyW7vXLYI3g3VcDfVYv6PuwPQgAjp6IK8cItzbYiwGXA0ovzeCz
3COt7U41kHZaCv9ANfotJoLAIx39uNJKepSzG56LIHAy9rWtQbESSOk7a8nnMFgX
tvEeOqNjKacVu13nBaMjl21hrJrR2hxZiWyOw8+wZYxJTvUyPTkKwU8Oo3GMvqI2
g0UZtE2UzRKGOXTht3r68JHH/170NlfLKp410kXLtT6yNyBqZ96xUTChToSF/BBR
PuDoHF5Cio+MlJGaaGK/aLfdLIYLQsY0V7Z4dezITltkgNTwYrpw2PjDQhsCDmIy
Y0L9lTAcqPUFcctp1EsTrku/A2mijq5ikEBRKa7WLXupg6rlZCemMW06W074qsZO
GkC/e6rrtrNO+zQjLurSPBbtuWlvvNB/CVuJ3se6lk/74a/Ex5kKRfzq5PKkqM3/
P7k8G+g2bShJSy0hxBmmJoM7AiZdHb6oFgoGdTFt5zgsKsEUdfNQa5dcp26YEpCE
+wd38QSVPTY5R4hnPEPi3UvpJts8SUjbHq3VR7nk20Cr91cUeH9WqBWbT9RF+tJo
jp/nq6WfHu0lyxmVErt7IUTTe+69YCmm2Ij5415tM6jqYK/uQkJ7xI9c5LWXpWEV
nIgIRxtb4U5sqvrTuP2nKxbQ65CTuZv5fhhU4vLjFa6HcyWLACKJDHghM7WqFTcn
JQmQm42bLjYYS9VsQ+JpCWYTGAXXWdbN9IhFf62/Wn+fgJm8PEphXjkDbXfShMT0
94e7zFYwRSdlPffMiPx/mymXVYhOmSSAlKGum+ncxcYRtSDH6joLnqR0At3c8ddF
ADegb/0/r3pkgnRYskmQzFxmKPmIyeylXQgvvriuGobkY1kdY2CYIYx9M+ErHxXN
l30eRaRKFU27YMJKCmztX2QOwur2k0iDxP/lfQmG9uO0Um/ybzbM4wHm4aMOo/6z
Zg2tCfHaHB4uW+7cgJf8IIfqOKkkypvDBiOIGI6fWallGgFoEAWU/fFh5hqQ0eFh
1wmsMu4lE3g4Ugve5ZnfD72Pb4QtgLFZWqyjMLojsR72IEBMxDiONfuaTdNykZkM
z+hOWBDlJBS90BMEKpltU0MdCGQukrFk1PDUB/C40VQkdjYJoiuM8nopXYUdGnms
rhpM7jhkdb8oz1pCi6kCoXKN75R1N1gH5BCPw3PW/2JAHyd/4yHIuJC8yyqOvhNh
sxFNqa1HloubDqc4yfdHvOLt9lpszVYReXimL47giWOGeJE6LwFWh13UB6291kQO
zI0dkiZBA4a4UgD7l4jcht2JbMyIr6LXeHQHj/ll/LjH4f4we6VwemwSTwuy56py
3yCLKsV+Nv1Dt1BfSPbPQGUamkOk/at3hlMlW+re0rykIT7rA9a3TGTGDAvmS+Az
XajwP5ltIOu4zDEKHZlSBctgJrMdHOH/ctREX4E3Xshy/iyYRglCN/bX3RHdyHvO
8zU6z4OUIubGq96GlVmwgUx7OsQV5HJ+17SfG9QKdfx3CbJE36LvJ6wXMkIzOzbn
laGCCSF2F30XDPPAiIwY3ohBYfBotgHavLFBn72qjpkjhPugph0F/whgtig6Ted9
dVkdOzvn05Ms9SfJu+YFYrnjGE7Gmn7Lxn2L+I9PvB1QjiM8WrkyjNB7A7XXVrIg
h24EITNbBqhqSL+3pm77qV8VjoyecIW3P/PmOY07oSlrVB/3SMtFO8j0VqnddPjM
tH63WRMiT2BK3xtzBg6UeA76d8537qMr5EvLif4E42W08TBzNC7c6yRAWvE7HBVe
4FuSI0/fcYPEbhJwxR9nT2RIp4mMW7iiLC3ayIK4ftQVBmGr+JFXfbF7WucZPujN
nhMtZdicGj0465qwFrlyYUytmRmvwKtzJLXHY+1gAvQwi5CQC3zegMzjY0fS4JCg
fpHGUdaBZ+dbJCPo9iYiCMooiHTQU6U4J4U0fsnhutZVJKkaORN9iFnZa/L65Guz
mlFG6ZVrpJcSm7ySY21mClR57BCKG1aB9XMj3wb2vc+Lvh1S3lWT55djmD+Nudy7
WzOIdLQZ9orN9f3TAtiyv7GUcRpgaxu7VVGwRUVc6I2KjYKCVkfBz1ewrgZQi2k2
rf7xtIzemM0BTVX5YIn9O6TjDtJ5Wa8zj3/uNL7N/G9A3HX/rL6oN0XoHOFHOQyF
9p0RxA04RYbvTj6+Xx71GIyzp64tKWvHPaK3Hh28fKXlY3WI2qgnGzSVk39KdfWR
8VF051UJxrZwTHceimb+ECTurGBaah3LYBMK1IkjDkK8xMN1CQh4cuIEiPHPFc3V
xTVdyQLQRjqOBlB5GJen+KIaucpyVjZLNS2iNmiv75Hj9kkvJJYDvITevSGDuRWZ
KlTu8UnEOa2JQnZLSwq/BuYCv7QGN1EKrRqtoXe4pXvxdD20T3SrsMAml+2a6W9S
SgK/5t4OuoW+9Q4Bci2I9+oAgOGZMjfyPekA97TWa6fbp22GErmsPktImoHNH9w+
JUFQivaEmyt9qNIlwp+4az8ngF82d5jJtYhwdCj8x+kwVm/OMhPuqIUUguzzZIxF
AQ4Gk0pqgtqIWt59fuXM2hcgIujXdocwCdSiHsF9kH2OG4IRmbWgsZid8lS0mOVJ
QprOb5YdufEHovvv0CnSz2Fdtzqy/uhsu8RbpYIu+/DxmH9oTWq/3hcRzoqWMQFA
1OBKthqcsWq74xs1ycFhN8vzEXKVsK+bRsYeETJH5qslZp+jYkXgkbxvaAqtpPIP
sDRrDCx8fuZvmnSTQf8w2nV+KSCveyS2FEFzLiYsr7oBPkUJ/5L7oDqbEHDJRuJh
UXVyREpdihg4FXFR2w5nNia2QKG6rDzRtZHpFyzYfnuU1SFa1krBRDE/NsVfS1sU
50OtV2Ra87jF2MF7v7K7Xc44EytaxU3DBVmdjUs66Jv0iJA4O01jp76y3REDxx/Z
JxtncAZ//aXriEPcaAqWF2dfN1xbwl8hmkaN341dNMnn1UvUNrQ7edd6Omq/J+bM
estlxrS3jV6YuJdxU4VUARxtW05nLMktGyStheZ7ToYj9/L03fvUuH1wUKUMiMW7
Ab8ELBc6pCxej1ueXuxJi5hMPmka2+OGm8BHeYo41aH8DHci85wQw8PNdzP0kg7i
dXyEp3Qs+ELR8YA9zeinST7D/KnNzQVszlTQZv65GNwNtgy+ZOpuWU1oSnfYJ0Ba
sMqEPw7TAjMrRGQnej4eqkHPV9TtInXxdamD0sjlYDdLQQnhPLE6k8XKa4G7RXvl
0iVbByckXW6uRRov5g2CunyYbhT2rEzWMD5bpjpzA6Mz291Vn5+o4x47Y21uCdqF
Nh47KF5gVRBbJkwr2EbLdFx85GGCQRvVaWV2WN2bZEhHW9JsJB0yskzlAgGynFZ+
E7+jkqp3/p/w8uh4Eb+woLydiKZncTswSF3gUq507asE43ZCWdXG1t635D0p2qsR
Zcm9q9+p+cTVNr/YyySy0CH+m1qPygdNDUkzO40DcY+JUVK3alyNClp4ksvr5qMT
VKUsHmGds9jvGNBorEH57edD5at3kwzx1H1pvzRu/p7BRDZGwuahIx68xX9Bh9mH
tFdVhuT9+RbILQAhHKOBIyOlt/Pt0N5pBRnNghgcXGBnpOEYXiSoxXE6PTs6W5Ph
EKxyIPMfW2iJXRzGaqBzOp+FSBmnQg7JPgHB+I/ec+VQaljcCfyW5Hrv8WNK4jq/
Z/4aft3XF1JLcyo+lZpA3wZKHzXYy3dfnAosCxtaKG1Q9kwMcqlPSR6LY+vXQcBN
jamsNkZLYeuPMpH9wlyPY5fneoWops6lewldyOA+KwEemJffSyL+/U9DJIWrNDAY
isbvBRHgJhOWgiFTarcynXPAoOtLQymvItpYIU2Ya6SeSL8GjkAqarYjy+eLPfvo
7v8HfSNKMJ/AJlAWs7EEMbD6LlMBVljri3oL+tHvilgGNmI1XYLHIb+ERjfO9XKW
HCo6k3rb1/LutJ6ajgo+nC9rKOY7fJ3Pl75IHOAfJcJpRJYfNAqT9C4GcIhMHvXg
Np1qUXD/2NZpC2vAmVD41NLwlenQl77UzpWvqQkG3Wf/JYtvSaT/eDlKCqxVPIL3
OJlJ21lr3YBXdyqkjG0a5pwvF9iPuUbGjEQLwlHFQjxkMqdF2qMs1wsLnqlYy9JM
44l0Pldoi+dB7QrZi9kICtQbsvcYCSPoqRvEgWhkgGEYZc5bCAWh0M35OQN9C4rz
7ynP0u5MilTHsayE5rcVokxHwGGqRKbL9WMJNI+n0viy4Xh3s2lMe40Gn3LzG6fh
tUBGkGvYeyTDNbJsmxq8mf0kNyvtwt0u/Xa9Pl7SGynwzrSJO/8WQPdqgskKanEt
ZMlGiageK8plMMvsm0unFtO83v6NV9c2rso+4Uyca4Lq5WY0e0aEjWoLg29rLvUh
uDJ4Lvgjms8uPJpGVWxH+jC7e9d9kE3cIJytUny2g/bt9ZqUV8dUcyRiMGjPZAdi
6s1LrHAWEgu9ZZlE/JS61+gk9yIR72zumrDnig7urxE140EZALiUiRupop9xKakA
iZWDBNG9UBLdWJQd47FiYFZdgliyTYCDNsmOtoLTZQ6trlgjuZ+bk4oo3vXFJOXc
N1j1qUz53zerHjW9FQ7OYS9DeZTo30rfNMN4CfoSgQsrA4U1EvHlNidhATx13HXq
eUALR07atkRCfW+G0fE7viOb/r9KS8Nfc/j9gsnDiCn7IA0eAZakZ9WyWCZ+bHsY
1jb5HebtS0n1FszMcGa7apkJDyNexexFv4JHVgI3Exa6b36ZQsWfh9FotHd9Jg0u
LLXAMBfv6Ia25MXAg75fk6aH13vpglpbQwqXCb63KzZA95zjVvTS9dCQdrfwZCyY
MO6wsaN5VVeDhWaWqWaOeNOSeEWt7YKk6gz+kXMUFqcR55VQuBwArGlvGLpS+75M
FjZvxFToFmw8DdhiB5Qy5abR2wbVS5qQmRTdCOdeaEcjHp3b35AZ0KQ04GgeXa2m
AOnPiIidXKHVJemC2YVWXufImCJcBsCHnk/XQLgw6oAchWRLfizXkYsddE4jjMhN
J2j2gZLaLgrj/cycKkZ/znAViGEz3tsi+/XeKsrp72Xfp2wDS/gkbES5J0AKsHqT
qClRqfT69Y3VyfcTJJJ8RAlvoR7HfIzGAmy8jYGJrVLEXdz6eMfMbK2/m/FPFm+4
wxyQKvUkeCJ8abrK3jNfRCSGbTTzgl7qdL5gCUz7AV2QkOCGkFxyMWP4Uv/uXeBs
PFZ2Pi/jiVmuE4R3LA44q8cMchJPb34dXv0LOc3YSsqcVpc5BtLAIFrx04wyvCUi
3ryW8QcQTOtd0egXEI7T5JP26D3+UVWVSZl3f8tiAIE=
`protect END_PROTECTED
