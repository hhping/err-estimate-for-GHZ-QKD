`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2pr+dddTWAMMETQXEsHeFNGeqmofyQdqsdPrMwis4IUVu3PVT0CtB17lIZxVY0Eh
Bw9DJnKswNqWRLZVHvVHoFuOhyou8lcDSOzRco27puQhUTM1V5ScRnYgEl426xT6
pJdZa4WDp4OxkaYE/JpqklcivjJ2xYFu9bGTQP74gyGsn4ZR6ERQPBa7oWXH7q5o
DjBQFMOiruC+fa2Cw4YrnaqQukqplkBYWkDjI67c/GXaxV8ObeujcEcASYE0/W5n
KAe5tWeDB4kQ/ycqenszmXTLTwTs9+Tn6SssqVv4KVS/cyBbAkxMfl9QsAIOiAnS
B/jyG0HKgk/QcfowkDXRI1YIcbdgeETaIFTQML6G1VRXlkeMmRXEH/y8yXqXDdXA
8ZHKdPssTaGojji86UkHHMLOASPmpKTViz0ArJxMcIlIKR318lk7WpvK40+f5c1r
Ua3IMywrTKAavSQBW0HkBI8APS3AFK8E9JC9pfg9sU9NMdOZs+hc6yFZVmODZGOj
6Nvm37MDdQ3ZQHNHsBsNCNauCnaoISJo9SCDkCg+v+t/InVhczZItPDDTs9gjdLX
e36ocbgvJVA9QA9GvSVDriCgB3EmU9kicXbTBKOeBzRbMEh/wSWjvDg6yp/pRR1b
O5HZSPSzPPkFzeYa1am5r8vxQ5/7qLCwGR9afWYSuxKFkLlR421DaWx/FaIsBA1q
3TaFp2E5qld+RpeKRzB/O+xYSMlzewz6SD8/lsgZMpjvXN+/1tbstB/o6uCRR+Qq
GFcRmxQX9e6+qdT6N8hUxWoaccbPYXqxPZL/j1KboIlM9llNe1srVfeU9iixVQ9Z
`protect END_PROTECTED
