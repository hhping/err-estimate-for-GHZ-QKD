`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HtRM/4E7K0x/ByIObWPwI/7yewPkAfziW3EYcOf9isPPN/0hcftIQyT7HkylE2i
qEuy13uNxAw9OXoUq/4kZWFOTzMivLsr1hNQTnFUcdvUfQNp5zavICoW6rYIRZd6
Dgd/5PJHq702yYyQ5xrSSsrGIV4y6P33p3UQOGlx0XJFLwhfZW+TJJzamgnLJCtn
1s0v35RhWB67LYYrG9dhIjX5hdjAX5eQG9H+9ZCHu7HL5AlcPxpC2kx7E3frBYAo
SDw3Xjp5QkYtJAgPJ5Lr8kZHD135Y0zHbla2DxVVDM5L+KPES7xBhg2IFKbgvY78
jjJoh9ZkUpH2eLQv831EVns4r90w+79qAiSRTRLUW7TKqvELCVQrt17DPqgwAXb5
L8EEkHdsfefSrcWFk3c4bo3r8gcWJxk+egc1TrRr/QpXWOTYv9LXcUYmyEQ7cdbH
e5hsRtyKVWmwgtFUsCzaGnGuvFsxt29CYNP5eZKN4At6J3KOpSza963mc0v/K0v/
PpZEDsAi7LDi9STW4BGExW4b1yRMROxYvN2R5q5aYf3bC4wwhAhcHJGKsQE3oyog
zxIegrRYjhNlXxXbbe2mYYSJrbNADgSC7ETa18RZ3piDPRTMRlt4BIqbnDBKy9VA
kIz9BWauS8G+lbj9OvEEKKJoJMMNN/qVGNy8rHON8wsUc2gz4dqOogXdnlhxUxe6
b/w70bf5NkNGWqqoDSPw27Y7ejtVA7c52ckKqPTcmnS3KLmZwRFEnulmYlsNQR6h
h6rUQtGzOqZoWZ+irmaFv/KNOjBYptzdX7sdwnqre07Njmhbt4VsYlkT2XZib2Tk
oa2rLHz9du9GN+xNzEc4+9K0J4NzUTUEebw4SH4If5aK93ovtzvtPsZcAdRQztbY
GF4+WLYj4m09PGRDcVhr0XBmXaNZLQMBFKX21IfcwOQxmzRPa0uhpYS1BpuAxwRp
1a1Ijf/bRr/iM9k+hKeKMJSJygrAAEHdxhYe/dOE9ciX8ASEVMutBAMs7fANk9Ny
QJ0jhEijRndx/sW98AB41TXqYn4Cfz3Tu9dN3yi9hvjgBMoX/Tb0/uzdkK3HxYwp
b7seMqLmSL8BmN8sJ6sBZOAraLeiQe1abG726dF8me8/QvoWoErKVR376HKY2okZ
SxWcLBEXE0v6xjsy5EPfbCRsdnGXTHO5PNBfo1vnISLpoC/gShKzn4n+7RTkz5I7
XGyZZ8Z3bKOwNvUZyM28mvZOtc89j0dgdi5JkW54LpMmKjALGf10UqetkGh68pTj
FSSS2k9nJn73YBc5qBjz119dDvG4DTgPKSwMRiEKqNFtYDjOWvaqvmptvJzJchR5
6tpfYjfv+1Cx7MjkHX34Hu+UMaohmfjUwFCziJLlcdqvY+Dkav6U5iWN3fF5m/zl
gj/eKhkhCNM6+aHp3lBpHG/4GLNa7r5cmpd4LbgjLgXAirsjgwXFmFwBOHaozj4Y
MKO8PLmGQ5Ds/u9VIH9sYbPTH+Gnf8zL7D7Ic/2zhw4Um/OXXu0FpTV1wTTI0L3f
0Y5hKdrMgKvtCtrhYBCuacXlJwnIWYK6TPHhx4IW95bo5pbYVfmrELcFlnPiJsBp
c/eAN6kS6XV3WO7qbkmzVkvdHYqO1EussvRQA+pHwafuibM1hVqGRoUDsgxntA6H
WnX29FT2HxzL+Ha8SD6BhNovDqiaaN1ETZyJ0sSwcUi9ElPaF+6CZtTRa4Rk9q49
oGc7uzjvpeTsrg/TGOTZXZOXkUpoPGIVP50TTGqe1HwLbBKMB1XNgur+1QsydkKB
db7Vk+TuubV1qZAsV3rtCdXVQ3lz/VtEgZHNjpLwgEp39gWVa65wpvuQFtfrDaOT
ahotfj3fv+B75WeqiSQn2vpL0CcOCHqt7Rsjpd675IvQhFoJ4va0rEm3BwV4sXRP
wxBmXWql8CR46yy38s26V0EH06e4+SGdLylc3HQlmYQhsKjD4074bCNAbzIkddrh
i8LatGgN64Q+j03gf/pKxaJs3MhtKOMf/uhb5FZcLgECkFOblrUtaZrGlPnh35v2
8glbzDLGV72pLEBqCNEhXqlgN/3M9M312nt3w7vpMWBnD8s5KcGHR6fNBM1hnSyM
TJzPBXv/bTFGFvkapF1VG4Z1SvZn/IUVcDlEMRRP/g3ZFbsp1ENCtCank/NMZ7B2
m/m0rzPEvoVuNSTdVifjxhcsbD5x4jybTChJ9yms8AOxtvVjkJPePsN99JoI6wa8
xmCtJxM1kq8w3Cji1w1BYAknNxJ7lMvS3GEB/qvYRyVec3sSYwnEP/iFHOdHRzGd
En5SLsUGkHgLGvxMQWTWliQ2RrE0vINIK3iflyp7LWdDDzJTBmlKYou1qlYj1J7U
3dr5KTOTzC5vRGs2OBpqURBJ/zbZZT7FQEtefBLmPHR7EkfVs76tzEV8ll47BiGC
rvQxXMbPIvlX+vkenc+/k9nJvHUWpymifng+2iGP/tbLq85W4J59UYCU99Ynx2E5
mRzBDfi2a/CHu/s6/GM0+MzV3kDeMzQz1IeTyIhNwiKrQUj2zxi227L3R+TC/8fo
DxQQfTh6JS9qgtW5htRxA/tz6mzgGshg1B9ffF2s1CJnLj3KjYX+lydEW6kHLtz6
7oocb8V9dUByPc2t3mmAekMbvOZqwqVZ2+IfCPVHoZ3HQsDFtaHk9/2sbl+TgnXU
z3IY0iE3JPEfqRhzN3HbpCZAwru4jTw427QJm7Alr+vVe8J/NIVRcKkVxptQLjTx
H1SstZifLf0610kDVn4BnqnwWVxloOity13tnpgkSCHuboZMDJ0AxsV5n+CGZqmv
I1oHW8Lxr2bmBNL5c7+V13PXCl1VdJUCpBoo9QBEtBAQbLjP5to78Y+pKd/S3xMn
4sVu6Txa2ksWxx1DZQWMMV+5oYbw3rlImUcEWCa3+JupXWr1qJPxn6gIJh5LBSl4
ZPVBXbJDY0XnNDRML8+qanU5sJOjCq0Jd89SYcv8S1RPejrqKYRxIkVw0J22TmHZ
G1ow06Bs20OMBx/Q3fP0qOBanXSdaoYKJRmh8DveD3DERiya79blFgzuRDznUN6w
7q5o8iaSW6sAJzNUEHpCwQBcQzNN91w9vScdWOfteC9LVPmV7LZD1hIGDxPttpMQ
sb5+1KWC1RQpSIHTBxXJRNb2URDrNsSepWQB0tsmFUlOtS4ZJrfjabfmWKacw9Sx
jer0IOIPVgZyVinWcQjSrNhZpeIzUzNChrXntMjrsPEO2RI+lgLf4avl5RFugiVo
SE3hEBUo7FDHrHSH9yTev6SYdno05wXa/DwcCE5FrikOUtGgTnfQ7pqIkuljI8qD
/vV53M2Ua01tMrKJHi/KIdi/8XETSS+jezdggD1DqlX2IVQ9VrtkknBSuqX18RoZ
4d9GAYdrBnZ8+CxBOqz0dSipZ/uXmbjaUMRsYOCy9l5NPdc4SidNkTGIKGYoErfz
NeH66rJcdX5HZ0Xbk9IHc/Xt7ETkefxPYju8dvAFVszE8sVaItHM70UcjCHGowoY
auj4vuAlh/CM5bmauWrv4GqWgHo8l0dJHZY1ZPfBBDqJz8X/gS1bVqgBWSjnD0zm
Tuc0GfPm5P8Doa7xwmheojn4BfgdTktH7Yv6qLxrG+KCVzGI/ld9da/0ZUoYOVNh
WVCwdGuVwuDHzDIaAig+Dbs+ZiOxwVjxziPBaR1+ckZPIp9/GiE/kl6+nksEmeEG
tVit9zAaixzIozR2G8o0SjTqlQOGJDH7hzRjhdIh+f30EO0ddk0rmg61z84CEZrU
bLdY03wX326Ka1fziusQhgvzBmD0X/qTmKsG/Zy33u4J25flbOre4Exbq/iRzE9Q
klJO8KZ5YVrrllXzIV+2+Ndh0/wtXhYStzDMizGyXez+ea0sRhW9Noj0PDqQjJfR
+UwF3+3BfQy7KVG0boAoHNxnnwbAMpIU+GGhhVVnBEPYgHVII8c9hgHmb/nJhN1K
mnABUcPngsiK78MYeQ41qBTb0UbBGZ1JSzbLOBgZmZQFLCpRHQYB1PtjVD5I/585
7+yYxgnu6Pwj1uEjV6zu7Ll4Mwg4qw8cKrUevLTNQlQ8SmMFwnWltjh2FKqBMesN
kG1DcMA1YRItUMIq4veUlp1uN4/DuVoe0eGj2JQo+dOOH97QevmzwmgWsDdSO6wG
4676SUMv/ghYM5eZrWLRDX40A0Wd2CTLojrgmCQMXJkXZjRdmiSG1yxHA3GP/TH8
rrbD078tTEjLo+sRrAfWKyKD9ZoWb/w4LFnUx55xf1LUUMl8BIajyLVn/IO0B4tc
EcLj1HN1z+/0z9r78DeMwLSKKFC78zXnblowf2IZUrKGnSUcutCvboDgkRZsQNqy
98ZEHHFEPHc4i9taJCnAPocEXtgPzylWOeAtz0avMNOYGGxwdGo2zxjBHhCgCjd3
jFug99zDsAxLd4NXc7QCs6+J82I+bQF3Y7PLP+lobZJUJEIjM6SYJPrlkbwd2vVa
BveO5IDqV5CajH1IM3VVS7Yz+1XDi3iEH1L8WPVR5oIqzow1vyEkLmhAAikA9tXH
Qbid1NuHoG6bVo5qCbrmOxRm6rdIx2baAddYHcabMf3k4tZr/qfx+P2PR/5UVccc
gHaSRrQPrJNgE12iARIEX5K7VTZ9pUmR2GSd+fbUQKWjFfnnY0W+k+1s6de1qNvv
ZNaDEiqF0eUD8cz3ahWswkx7LGPz9Q7YDWdGa1VmlajILEcX0LZjYPVWQC5EWbUV
1Asv8jE6Q70dPz0Fb3xj0p4EipFXtGfL4pmcjTxI5AX32e/UE6NS6DSGIcYI+MB9
Jh8skJnneNqzKoRqVR3KgXavYmMZId7r9JKQ8t8+R5sYJwg01baZYET9TVV5f2ov
wv0uqtOaA5hqEKhTFoegRL/BILMJGVcBJB9FLzLRHfZur9VamRbcP1Cc9WzrojXb
k3VQca/a75rim9I+vT3lpFVmoWAQ3tUPS0CkCyTLnnXS2tZSTojmQdTGMwm1A61f
CxwVcWY70pPsPN8Rv+lxnZlC+YJREtN3lby9M06ykqSf8qiGPn287+J2B1drA86j
PI9mxKDZswVApfhMm+NNxTTSvYJHQotZeWB87VsjI/N2Ws4cL9loV4sTrEowC3uC
8XOoG14Bh4bvqCgHZxhMiPRU1wx4cCElmKno9CV+19j+rK58Exe5SNaYWPmuSlo3
F/EV+sHYzmlj9otqSUOAh3TKtHKbTYXli9f8jI0Z0+BAPyacf9U7V+4YLKidyY5e
Hhcx6rOtqycpU3jGHkK7iA0avNJTy8bQ4lf7BSt0cGV6oq0vCiVztwxrp/AeXhv6
2kuY966bWcz4RsXlf/NR1XVXNlBVtm5jAJ6rbnem3xUcW9qeTOoQ0KMagf4AIvrG
YmVEIWGeGyeqcelthdRGhfU981Aiytytigo5E8bN/lXYbML5/aZBRAabqkO8FYsJ
pEvPDDggOEFd+R37i3Izp+tbbgkvH7LhODcYVem5ktbjyKTT95elT+bPSqvJwGw4
Tn4eF3MMyYHrOdLvPe+/yWmcWts332ecAzAnIE2gxByISNj28OfWQKNLwolc+Q+n
PLY1NSo3gvHfed/5aL4ynNLlbkXyirpATgZvhi1pFQzJWbNlFR+HjgyQyaGAhj/t
BrVPYmZXpJ4J0fzpRCpNNbCuXEdfBeuSuCPO1rXAOoMSgIlCtJoALj9j5XsVGQGY
Xmm7UULPsSbrxO0xtthlPgydjjeeS6RVuWOBA+zMg4r/SRsPk/iTE1OvQY1/jxt6
AvDW6ONaKpmj5elsDbG1wtOOsdL3F9XPZablpMceIKuALXHpAj7bjisIIIx+q64c
OVcddsgrkn/pX4bnF55wKcgKPYYP6e+ZXzM8YXW9TLJSNybupT7Iyz1+JMwKVm9m
o+ViJcaG+/+W9TqB3axjHlrP3UvC6g//BXqqlDZeHouqctSSqmPu4+/ESLQOmp5s
l7DbH83X6LzXjNsyqxbYWYkz3nv8WoVv1Xb2coJT3eAankLRo/JY+ud5CXRGImu3
wbnNHxam3zPV2XiekS5k3NciX6FIuecKAntVS7XhNfxD1t3m78jLzq0T0DEepPRl
v15ZbuCXJktbT/6ZCq1Krw==
`protect END_PROTECTED
