`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNRvfpm66MyMl/L8vSXp/oaAasTuTjnhzo6mBKWoya1z129A/Q+W2CT09LFnE9fL
uDtxBDMrPqzoI0RGg106NdX5Geti/J8MdMGx+3KsM8sx8BJP0FVcwqDPH2p5fc+F
DBVKQQFR8GCFoXE4FdSq7FjfDodmbk7LELQ7StaUOHmBi1japkX/nr91hVOPNyeo
maCwbs9atu1/D2CQuuS4iUrjOdW2/PL411Jc80ca/3+zhBtEv1Q+Tu9U1ZT4QB0m
dmOPewTPKOVem025S4b5g0On2OpvaJxLumeQVvcyS1blwJP2G8v1oM+B87dSemdj
/ryWYDjkFY5sMvmb/QXxJ9cfhcghyK9G26gfBvXDP6PbcnTgKhVZMcObYsSCW9fY
WlOfKv6bj+VPhoBwhxoBtMnLynbSKqenuAi9JFrW3rTRgG8tsIITx/oP3HeJsDRB
l617XMJmuWe7Ilc10QSm8Din6bsUzSYc2VCcUE6Qo/DJua/9iUy9/OsymggYBY+i
YPamH72Mi8GCON5owDMzjAu/J1xgwJNHkr5OmY0fM5FB9VHaJ0xcrI2AZUm7RuIK
OWFV09OkGDwG2syI+Ug6fVY+oPsKYpCiu1jxYBmgyvAlf47vDz9IxybkgvRJ8yqK
q7MQVjAxx+gFVX8iO0gZCEniGFLW36lo9i4plIACrd9esYr8CRe30Mg9shkyCdmD
V2iklWt+0zhtubMTHOcGvPRG9/FWtaMJ0W+qWkmX/m3rxzEyN8/ZI3zOtWdt8GHE
WuYr7mgjhC6hTWag4EsYQKn1cEXbGAV+lziTapcyF6Tw1/uqM94gZ8DQck93oX21
0CCr25+BZ363vi1WYDrFSGYTdRGblL+IUxHG7FiZr8bom3m2OhKVkMyDLWE6LwHy
rMs82tuD+5oyg15uB/M1AI35A0VY3xmn+IoJ+Umnc6mDtln6d8WiO1LTCOydrPGd
Qxzl0GVKSJkNLMdK+EJbqN6yQJEy0l3+DP9S+jr6fLOr2a1TrCihN0EiNLH21SUW
xq0KtRzkbUrthVoaMbZF8sRTps/dm/w/NnVIS7SJTG+0JvpOcrJvFvkfgFhmYhbi
ajYqPBZQVmD2gmvYMTiWW+GEZwwkUVYvNJcppo6njiBHFHS4FWXZoHrRzX3p/714
ImXbgArtkheSWZlCYGC3aaCcpf/462ou/0iboGRAK2zato8+vO1pHit//Rhgk7oO
sU+RdzB1Fo3rdaIv7gH5qxvgLtCyzekCx0IobO6E1roHQ31uCt1NL1H76yE74psV
+/T99OLxhJRMkKxUSx5vU6oF4anVghhvwi0S+HgEMP6MLFpTggnMNuIbb9RIgFG4
2MoCZlMAhG9Eg8PIuLm8Rg==
`protect END_PROTECTED
