`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8QG4JbA/Aqmb6DIq7+u+iW/jz51b2nl+hHcGJTXWYVU4KOjYRMn9TBWOapYvCcs
p4UxqBt09+Ftm/PchNUlDIAaiw+hMW1NoGmCEG+OntGuvDqDx0o9N7iLyr8sXnn5
NdTPxIAw4drqMCmUvz7+FGHPF10O39znnX9BXCCMl/79e4p3aN1/rAukemXkrAuY
fG9UKgJmo+7h2TXK4ks8I8waKOgkCmj3Gbopw3NBxReWYdxWyhq1xjp5NpqQYZ4D
yrQhMTbdlg+RU1cAphJhIng00wH+qBODHF5flhWVfJTpsZzMwtSCn6Tyatpkk7Dr
tCQUVqg5ozx09XiF5zSaGsE25vItwIfIjZYH2v/hnyPhgImoRaPnJkOZDNFVv3uz
Ksx35UJQ4dWaHaEJ1VaAo40BHzaWHDDhjXogAF22k5X0hwlvyCKP9+ZjyA7+i98J
nOGWBDl3ccIY5Y6sAz/DUls1Fer1nPH+0eVa5v7NiyVvBYLtTuogTXeKDFRhivNO
lY7mnkv/YZYKwCGx0wefH44PVfWUo6iuG+4tZop5hYDZBjCY/QO4e95Q5ch2S/yN
VRvJzUucd58YJEnWQyr2dZu5LdX0KeN8H8rgP+RcuO2kDJ7oZzQ/6ekFZEaJxnZn
krt9GjONpYMePpg+DEimw2KvOK1/emgjd5HTl4q73Crb53bYBu3o9xM3GyoViiBz
GoyoV3hbglwdiyyqbt8uGLr6zX3+pnZULZ5M+ULFwPp6BI+psd88KaUd43nAMSZC
b1Qt1cNvbd2GFlMptKB+vv2DGkkOwwrw+iopBEQJrC581yhh8PSLkBVEabKIA5yI
xS/xGa5vWF7GFsJAE5P0edBA8XuVjijsUp/sd0LkCqsXEfARwyso8M8NBZTNJ5tA
ya2ovAH3TBkol9UaFj1XO8Mr1c0LUv5nC21D8ezQk+LyvqIsyLgVE8xhiMosR6TJ
UyI/DoJVfNL3pWKxqFoZ2XaTZhFyiJNVf/Y315RyjRbgtMor6UnolCHGdMLfiqqs
NwPFqG7WdwFGen9n6fYp2E5B6YHZs7BxY9hWIb4QtTh8snD8wIcvSLqTNW47khO1
HMvne8oCURNxw+ThAnaNck8FzjS3F0cDsY0ZDN1pm9cgCHHlRfNq4yBV3EHuW18x
Q253j/eQSVTjlRCtgwBId6XI9yICrZRlIeb9ZdlHK1rqmaCHRgGNRCJMDtNhNjM5
KEs8fFMFcet7U1qSCJFWjpcpm0ncZ2+6vYCVEvKAyND9G3pkc3clqlfUnL/bgyaZ
csFoROiX+eVrgDWMHa9Lq5avA+1LZN7hPbCxhsm/AwP9tuwp4D3WqDfDgwi29fyX
iEeIoaBquTHoCqPQCygmxFOKVOy4fl68JHB6d1JgPAGfj95Nn7/o8yXNK8R7U2h6
Cqvup18FB2ABlbA6rmqgWZzc8ymCO28P+ihSOkjsWoA=
`protect END_PROTECTED
