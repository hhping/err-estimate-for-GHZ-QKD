`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/FcHUG9uTUauQGUljYt0ELrJak7bYa3OX+NrwNzxTeTcDIzaeD1lEfczBNP3Me4
lPzkQ+tiYZBi0pwp+w7BMR+wUKPQ3IemMKi4yt53DmMAsvmX5LOAAAs5adGr5t80
CM1RPl2IcJki791Aeav3LoqEFBpQCzHFj+nVU8F7su+eB+ul91aQxdon6g3MxjMi
puCasJTMwZDYmComFAfDnVabk0NrJFS0OJ+ral5hJ9/+fI2lVa+oPMDpIOBzMaxy
s078DeyoV8DIhzw1B9zPyC+ecj8KwngJA6eceTU1DO2Mh76DApFUXlUXkEVC8nIo
LPkRhNA6OOO2SAdsWKw8keRu7w+CmS/J6VDMHwuNzP4OAWyEV+Ksp5mKWmmaY8VW
Zn5PeQGmrEbuVbc7s8g9IKfvC70R01qJ9VD0CWuzVZLUJbeDVVZ7B2egsQV4E1h8
sknG73FP8NtUek3rX9KZNEE9+VNBVpdIoNuJFypqsbuPR4C1oCXLRY/a8j3HHMzC
AGW4bgmKXMgoWatuFBJmM2IZDiQX2Z25lzJksSbDELy9H6J74EH9kEd+c3/3sgBV
ENdcPORr9kZmYkjNra69WJcEIT9/ePEi7cOZsLPKNSj5NfyEHk5evLFx3YkYyL33
RJrABGdtDpgs9fwG1Qqh/9PWDCiTS/0/q3UjRD+msae3jWSZUGgy1pYhEw+z1lgX
uyIhQ9EiIjjzVohOCPeRczwx7rD7iOnO3AgiS4WQu237acuH+Nliowpn+NqIscfj
WxmgkHySE6nTY+gRPT8lt5/IVQ/062drJw6Zf+Mc2IMinqdLnLX1DkPN/+0uK/qw
P//bbzTu3tQXf1d4rfmrpgjWnG8y/NO78t1v8wrVmxdYRDYCutLSc7agdVaaMgSk
Y0MJImi2uGUmqgE0B6jWR4aNR84OHgAZfh+i5KeKqchhZfMxqUX30gT+0J7bKic+
tGennAgbwfntWxsJuwiMvVJssclGctWzY5ZUX2INgYrhBRAVhIFRULgjf6gp+q0T
T8VylouJn1GmdsoLnJHpJgrECm2t9M5nWKgWxqwvaeas2sjqe4heyrz7DiGiQK4h
r3bqeni8mEIFMM9q9Muc31EwBiVCxCKPXL2AjBYGDmWLqhHx5al7V1huqMP/c17D
q+zSpGCmfC+a57z3P0mz9BboGwbkIuF5uMcVMkkgohQhKwoKc4DVJvXV61JLjArP
Xt1kNhaxMPGdCcFyrKbqH/EWDB7EpsBKrw7zw7zoHKvw9DQh//KTRI3HIqfspJ9F
ZUjJJ6Di5NzJ+mLBw6vKy25Er+YoI9puavO7eORDiAlqTX7PmISctB1GBkyzbuCI
vaDWb3tg210YQdtX8OT0xiso4Gnz8rXawBDV31mvEoRTAB/Tctk4PgYfQQM8Alwc
M4h9JO3EO8KYa8DgpYpT2YxnpIfO9q/5qPLL9o1+chLY03d+gVmlUd8VYxvjXppU
wGZZQ8f62LlKf0dk8TFbURG+jML1YVwIfGfC+mz4SXguX+AN7JEmP8SUOmdo2fJ6
Gt7rl828IeulCkb2wNFYFQkRdeO/dwpLRP9kXPL+jKi4IYpe22f9S/oA/jggbqEx
lcX352+W/akBAIYgUHyUVgzE8JhPx1yfbX4xHb6U5t/8KTN7DUb3yO07jAPhkRvB
n86f/wB36hH9NUlCDDmbBa3JhPwLWkgfLYwwBtHUezrmO6u7ppwLJrUcCcTGNqct
/AAgKKVEOyPRMqAamoMXX4OGut/gfzTJB2Vhh3bA4Fbd7e76XQClZrpmtmsKUTId
fzbpYN+t9mVy26YU6+woHIcbGSxyNyR8cU5FUBoYm+HQWMzqmndALAIQQrLS7/Ix
JTCidBc4S14yjV2GXKa4eX37iPlgx+1VN1KKflSf6YxOrchIoY3AQQv5hPOKb+Ks
GOkBgSFMyIIdqPwWKzmNMTzWq7Je/dH9pRWgRnX+PblSU1MOLkKkt9GCEYdb9gTF
GrFmcNX66rkG9XHz+aEJ9s2vg0+3BAPzzC/u3qHSbrjBGx/RaWeAab9+ciu7oHd3
buNIyHiioFkWBKxGlSNolGQNj8kdi7oCA0KYjlsz22oyLOyTnppvCkxlKeCmAlCG
JzHDSItupRsdlX/hpLESjdRTMACXqQuwJIsOH1YRhGASNBYV3izdwtrXVpXxLNfI
oxXDgT8hNimHdqXLn/bLGsr946J/2epkC3ZBE8xyhicFMSRMoa07kC8LdR4A0Vow
KvvcMI4WMhdb9kFw8hQe+h4geIix1798cMA2srBmxvpjFVJzbln+a3NSNlWqQsdn
MPd4XnmBT+MlwWBS0TXWrEM3CGoCzReqJaUjXzO3qJJz+lpgfsSe1Bl7WOfgir0W
Y/PNi+Oxq0XwDmlleN4m9Q2lNgM8MBEM0ItWI6uTiiDwdO+osIf30jSfzt/ZDmzZ
vcIne1RH5NkhSGsmxn+c7abcSAIJ2d/n7wa1k2Pic4SkVN5R335OS6U1Z4XMqQE+
FJ59vqKeVl5G0Z+YQ6sxTZA3aXtSS+F7yS6olSYzS+CAyLNYQ0+dx8GYzFF8EUU+
Wu4ikiXjX9U5/9hU7rL1yRC3XhZndp27IvwyxuVRvBUCekHjxiwDwoTALYLZrHOq
ygQQDgb8GaZFYNjcZTokVn7kE3LtFqHaQLRQ2L43ockhH5VJ+swRhsBz67Yk1rkb
CiCZv8SNre8F9wjtLH2fKPiOnxZR4CHUi/z9Oc9Cp1bcxEXSZx1GMCibpzDuqJ2b
fR9RUow/vbQAtIQ2dxFRSm516/1Nk2HP6oFwj00C5WSE4izbV/UE5eTR8be/WXuc
h8qkNWhVhlQoTzUjRnAzkyPWQkiEAgZLeGBOfl1KaPXC2/glZxrKUKAzVrgqGpb3
KD9fafN6ES39AXnBeAerLRZ+kor32MoZw2dMDFN/+gpWYIgMAnQyAG4D1x1AGV4e
v4l2H3QjSBIYz4Ap2X25R+9iZekS6N6bcKBB04O4uVFyQA03TVv09ZQeEO27H47Z
CID+Ynx5Hg1eIbZbBvtFrnsweIfmQZ1M0DwPVyyjHR8rHx2EeVGFLcafOG4mWEkg
RecqgPXMm7+Cbg2+iySzvY0xtzyjf3/T2cOFcwA5mGtrVTgyl/aVTClhbH2S4KRp
BPKxyDTBpaO4ltPA5Y0JKFeYrynwjKwofgAP/+1OSpwgmQpaGuvJ+pMKLo/dqkSS
SmeLIfuSGN76p84L1z1xDe1pGcJXG5iXzriH6QigMplhcy25aaOebpKWM2q5a3JL
W44Gzd1NFdzbeCs6U5thhiJoSQ3uzs1srjrdWoxmRnZpCPZjgiz+wCwYBd5chnKJ
swKtw5hdcksIlkhB3evTk98THi+vy/4KtWi12+DZ4zEPUQshHfW5ou4dQ4r+6jUK
QhqDJlajc0slwBIbsmQ2tP+TY8VyJ90nxH9gApOKQB/doQw9pm1fJwl6rlhIq5BU
9H/ncailUONt22P6FG74/vl+DHQI0YR2nvDe+tQVF1Jk+6J3NtRzmao2YkTbN1ph
txW/rDXHagXnjXTGtAYLM1xpHeVnJVh8Qn/X6VRPfa1Drw76prAikjuzEQqzYDqo
zdoO4AOgDkFrvFV77mOPulAMPPbDJzUMDsbxIQXhmu3kV88VIyvbgl1P54qLLuka
etu+flNMP+eEXHQMDxy4RRgEhTnUfr9uYib5AHf3yHi2zZxFiVLnzJzgB61ltFEN
pbVoEYDmHL2GPWI+LBdDCqFWp8hJiDUBTzJg+TKuXxcCLVJma3/ZH1t0NXfphCN5
P6SohmPC7NG9k0cuTGVpQJrg7HFGgc0548g4RROqDLzmEf8hlB0R7seHTqKe0aAl
z9ZROOa0WTmg2QT8xPDzzBIB0+dgaJflq6caGNsrHD6zdYxSoTeDl8cLBJ07A04w
R0IG1PpLVsQiVxNA/TnKqIKfdXEvJG6FdQq7oLcRph/l8qXU8AGS7+OTUi0BKl+0
rAA3LXKtqRYZ7Nz+ZA7Ei53HKQwTsPmhuYB+BquSMXVkJkk8Us0/OIinzwxYmeYz
Vk0C8FLwpcupDhWLCw2SunbZrMYLT+9Hv8O9oEzfjdwBpz5QXYJ7fPscSJqFRXLx
tsGoHgNopRjwag4f7lDcp6C8+3NWj/fHM5yHnWIu8JRhKiHDc8k6BBRRuVJzwG1B
sOhbKyERUn3+VET3gDhVY9yaEgheTk84WVhewMV8Is0/cV1sHcpx73ahEsbkcQPa
qRChx6ZlVms3QOh6H/u6Jg4vJnr8aNRjlvsOdj7arigGcU6tyuX4BTGgNGxCDJi6
3GOdNcmFu854+F2fRiwz8K5mexIw091w+KJQpQHo3q10YPAdwbppEsPWqVTEu/BX
hmQGOtARy+A+Yjx1HGeK34wffRI+nwj2m3GDbGgGNkjUXNgFeZrK8rZ/SUm4QMGU
ytaOXTQfrraurgCZ/CyA21wAaHsLyCext4RqsuTUSx1bObfk4e9wLGLLq7uxF2wO
qZ8CQDeJ5J8oSqdlzcjp52NsiP2niOfx1bX5rvxTqxmOUEpVq9NDiRgl4belRQc9
o1QNSfXN+C21OdEZtj0QqwrDc4yEdbuGRX7mVMinioRBIrepHQj5HGQWJ5GcDd+u
AQHk1jYwrq55ykJ/ZzTtsLGo1gZhkW91LM2pFGnMtNUXhSzKtxXzpjlZr4UNU7+3
O23NqqXelNxrnxGQC3/U0zJt8HwTL245s3/oxkmXOnMiQGPmZakIJzi/nFQfQS/q
xJ2jpMlMAjHe8CGSWGsc1Wz1VacRqnVXRSuhVVe4FoCoBB/KtHNxt4iffo25LpsG
FqJJQWUYfg29TaohtWYq1Q==
`protect END_PROTECTED
