`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OOIzgYCsM1CuCsj/kr+sZHS6sKwvcgxULM162iyEMRshjbb6VllgiYp/NW86LMkK
6f9IjlZxgWo7RBgd+IZ/z9S9HURNDDxvaxr4ZmXsf4p6rgU4BIxrFbc3llupsFJi
4Cfl/Vl7F0wFoq1G1U9qFS9nd8aBeMSXu83kdT/bb5gjecJ/LtUFYiwP2wqSTcDY
tOQe2OSSRkRqugKH96jJS++XMduBo7vk8rIu467kZsa2hnWTxDHe5zCpl73xsPvt
yq/XmeJXApCGskBuVXFRlD5qYBeWirK6VHF0Slikx+ccmdsYNh5RhGQxgEMS39r3
0J1SHaZcJMDniABttoeQY2zqkuB7xKkywsNO+orocc8VcO/wgXiQWE84iNTCtVCb
ryTZygpycLGPMaX4kB2scQcRvvlbVd+6Sxf/cTKvbQQPjOrnbrPNCBZosU6V+Gd2
b1Gg22RAZg4kE/yKuT0dx4VCwL29uj0d/H4IcJXN/3MNwvIJyypKQStQ3Pu7HlDQ
gOWT3rLl7h5BgBpfsYSr5uuxzP209SsOf6DXxpis8AVQrLOYfSkJUNLwoa04+Vhe
Y9iB2Yn22glCdT1wMQ7/MkEEqP4zEvt6VzdKkRxrzVxF5z9lmflQiLa+Snh6gHVh
IxOWEV02hMkhjp9u9f/+77AD22U6OexVn6dulV1TK6O335Pj6FHWWNeCv+nG9loQ
9r2Cz9y0ydALtHC1h4hS8RPrTYSrfu8zR+k8q8BmKyxxxDt+y6JB185NR2HpZC2M
Ytp2a2v9G/+bx2093N+S8pzJitrwOic7ue2rsb7xxUtxUx3obVE9YVYh90EOTqYf
keFWJALjOhaRE45N1vkBxEOcUlKjz3iEmnNQqFvK+DsC7y/bIGQDeebIdwATZx+6
2BK9j2quV1dMkw72rB/7L1X89+1isZCGtEt1jCL6G2fOn1TFyDt+V5/9kiCia77i
wRLnzyKLJv9ayTGn1V5yFhfyY3TrZyyuVomsP9auWpjq0/ShzE6g0ckncmgcasgF
4H/lxCfeA/nx9RRCA1MqoxrRqicqQxfli1hh4isFlV64Okx0Ah+YHGCzDKeerB0a
X9d9iqbMsgG7CY4BXPtV1XyRz1HP6pRI39LRJe76/Dpi4GiPJUYSRtr3dNJ15JKy
mGGL51iCHFM63rjRQj3RBj/wJrvfZyOaG7+pU8dFblzmLy/hc6pQyS8JFuB+9CuE
FdIUgJ8mKTfoeyU34G1vBdYCFr7bVHIe/2CkZSIF43ZwU7bLxxg0IY30/9yk7I44
gpeoBryPZz4isZt7NzzCn69cOyqAuV/m1ew4Dx7RpI3VPtxMxg/QeunqjHcDzFv3
QxTf0pZEZUGCMzLli/l1cN9mLbTR3U267d9pIb0vHhZ1vFSSRAc0L6Mwax7KP/GZ
dHusaZcOwj75NHdTPH1plVCraJsN4mHKI149Drq63D9xbDDOlqMMs4pR2aEbb7d9
Hbv3xXARaHy8I8KZOBWAzgDl4KXAvFuRgXLPu5wOjEjf+paMBabMa+y06QLOyPUs
0n7smA892uNekxA+3dD1O7Ryj1coQcEraJkGzstrv7j+4WDXj5kZbBE/o9CHCI8a
aFLwx3EWg0jTjyga6/ur7DluG6xTt+trZVFejTY5g1ipPnK/tgNg9mtbqCLgKoqT
EN+OeypJe+0CAUIGnVGLQXw8fArXjyYXdsNd7tewrXfdvRJEaDw9J0ESl0H9aypC
4vb9++/Zex+kRBy1MuY10XvS0h/iE+oeNs90HQEfSPx97bzGb6oAB3D6RWb71xL2
hnQ/4c8g2y67wlGws6GK9NYRvjFQx48Ge0GOJXgRMplzn9S98jU6PCO4pcveUBrK
MQs1jPtoPFQh4hzFOhQ0WcZTg573F686dZDA+V5vZD5ROPQkP6F11AGRueKSuYMs
3JbbyDQZ9TIH1sZBLveYOsfFML4sgZPT5Wkg1PlOJVo5U2cAzqM7ntX53GTM71Kj
5tYvmHQWehoJWCDZcXwK8KW+8mcVwjeAyw/KuGcz/g2xWBOeOcBj4HUAdI//Bsmm
zHdtMDE1EIZcTXJvme5U5ldXfWGIBwOcCAJ6+c9U4L6eM3nHV0MjBdwgKLFu2XVM
9OUcBEAUqibGwhA6OIbFYCDUmDe+mVwOYDZrMaTAkHFx9/mzo0JUPxn+/gdScb3F
1gZ12Kkputf0UNmVnXhvKPdodevEvfg3QV1k90aIJXfhLRLlDFUfLsoLX8iSLu75
FN+XbwL0J2JXqoVYNUY9ketj6OqgYiWQkZmX7OkCwmAh01cwniV21gky0bP6rklU
i6fDSV2wT2C2pK8fcspz/uFx9/BwgcpHFv42PW6B52ZgKuVLwYjm3j6NuE8jbXuR
PlPtwAuLO+RP5kZ59u3Zf3R5pM5OYWyuJSOIn75xjBXksxknQWJbsLDIWaivPbg6
k4rWPOje9pMvgtg6RWeOO1wMBVjpLRJQUIXIBsy16nGnmg+hBQA4lcYm8K3ElVEk
7AVCzMoqALGMdwB2MOXWvD7ilzYNpPbqAGe3nnaNrKuhd+WMxG33rpzpKr44CMOE
uHW7Dg1YFtMtqMwwkbWpV+xSxGUVOTz481FphHRpMpFN4e2QCp0V1OElK0AUaWv9
alCIG435ORyc/xy1dI6UhZbeuTDECGuLOp8JZ/P8E72B5zDp5bTVY9iObA0PcSBY
oGw5SjANZbuCh0/E4cmAh06zTeAUhYylokXzMs66rvH62Gdmk12wrQqKZUszRYdg
`protect END_PROTECTED
