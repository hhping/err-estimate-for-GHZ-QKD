`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y9zi6jUl+4PrDwOzihp2mbWDkHZequH9qA3tOz2aJLRHKVY7QePPK67OZJ2SjBM1
1LYePrAoiadnPGHBCbTFF344KMqhQCJDijs/23kvJt0X2Vs26FslqPU34a27sSZp
jbHMg7weuGEvTRY57hare5LpuPRHX3y8Q1yannMyGpE0NfDtkgCZFqFVQ+r/rCGm
fck+jWfkzhOWIRm7FuJjJGD9dzSXLc0rxPkyA0FiQx9li5gM7WClQGANROLQbvae
SZAvSmsAZedfE9Jf/oFaYzDamN0vZ/TG0Vmfw62zFoukYcVKP+CaMYMyXHTqmdd/
sj/c5gGsSY/NmBelRfCc6fi9HqeiwY5IBaSKQw9xqlCvVHYrjbUN4dRYNcAgj3C3
JoKpc1LvpYKVSw1W6JC/Rg==
`protect END_PROTECTED
