`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6kFXcRdDehP8X09xPwCF1E1F7XtGf5MmOXCJNlKzs7ypy8Mbv1P3Vop7CYHS3gQ
RonA+LutfvkduTt6MGTF/4OdaZ03ShksJ/SIaYd+H5MuimuEbWpyF7QtKnVX7eNm
hTNZQMa5AhKQ8dmCQ242e9Kw05DvjMi2O2Jh8et6IaUCQNsfomchniT6vLSrNkph
EykyBIvuYEFUHJ0QJITdKNKPvdQyolqjYmjft+83tYAII+FSoH/FkabIt8t65BKK
QUk2HJeneb8C+LeUE8gmWPGHc98Lg50amQDd1WWOJFJRWta/WHmpMGVQrhajoIhl
SoNvMWgndO9RkKwKnNPFMOJNwvodJmP16u6/mCoEuI9bGavCM/wURZCgeeCiZy/z
NOatFi2fMT/dsya6VVjgvW3zUYCoPENhsYl/TTeXVzqROWuZuCy59hdyDxvAY8iI
4Q871q1Hp9ucc0qBOlbNp44t2mdZ+0F8aumYkhD7DZ+NG5U/nMKV7m71x0Q9MFav
RPxWaDGNfh3VTZZ3r42zglyN3brvLjqOR17WRtMePtOCQRVxOrxD54Vc+Vx423PT
a5q5webaOpFkxd9QB0HqLYpAgZ01iHkynOXkfjW9fKQ=
`protect END_PROTECTED
