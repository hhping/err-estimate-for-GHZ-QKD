`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
saFinrDby+F0hUIh2G5G1ranDH4/ePEPQ286yLH3rtN9ofkSl0W/fRuMKvVEnaFx
rtLG1Xqn+0Xh+wU3A06JOoEqJFxLvdBzPaHmRqIpHPp4jw3kUicIhbnPPJMvxEjd
FlxjZLuhLJ2gTLtNxg0tJGqoTKEHxtIOGsQq0MxmIv5btYTlV/DRD5djr15jLqix
jx46iY8A94qcYAzzKYaej27QKQcGkoadEyZrpyImrSbBNoN6+O/rI3AjiBGAKp2J
phuDXrZf3WHW431rc31wBe2xugf/Zpez92i6k0Xmif06tHv1kyE1d1Os2wxnajTQ
VZqx21CFCUc1FMLuv7m0eSno2ALp5j1W4Kk28LVz67HLdO5VgOQGupPRrzTNpJtu
AS1TvEnbc36IXHrU5OEIVbL855eNjOcI42/K5pkE6TwHf6JfyhVMq2s4WtSuBll5
7ZY1NBaKDkEoWnF1pw+egQnlpy1PajV1ukNMNcTWbkXACHuZo8FoAer9Sla1B/5H
dbE0ARetHr5GAn5zNYY7DxcZxOqvvZGwgQ42nrvFigjfGqO7gfX3zftMWRgy8Z7h
iyrkEuiFysXa93UuV7VAUme2RAbLrEOrtCYMR7D9DxvHuqApUwSe2FQH4IZDWvKk
wMINs/4PGXQOW7H+vpm3FKFV437hyoZ3SulqF3bW/zB93WLBKxW66T2oOqTthAiq
uOe9aqfcGvVwHXjRcFhYdv4GzP65WFNFS1mIEbezf6Li0chb1/FsEIyp0EwYrX+6
vMZ5+6TG38xW9taUuf/6Xe83nT36DM4WDu2kV7MM9H96U/1DBqDo9i786kDys+5a
67N1wt2meAeMk954BXB4G5EMU/LEpx/xoHJXgFLrU4to7NAB7AQITTd9CHh6PtQ9
kuMlGB0jizSwVwReXKfKPlGu3se4QgOR7cFvr5z/nwcIft+7wWW0Y7xw8bCL+D1y
L/iCc2d1p4qAT66+gObvYmgx/aQ73vXl1w38kGnoghSPe8uJvAf696hrUbFe8HqC
ODkGtdnAxEYK+4HAWXvinht+mWcxrUaagK+S/tU8U7APqaYowRl/XchUk2QkvGlL
QlwJOag+Z3t7Vv547GNvlusbrON+KPdKp6e1Xl2DhU0Yxr7AScm5SpbJfLG0vKfG
5mv/CFmWzpjaccQwkPNSUjQgJPVoNrYh8BWyjjfasTSKbXOSndRh/VAnizA+Z4G2
Il7x6cfV1az9ssvNM1wX0K0MdEMBIWwwL0MtJkKCF+plLTWqQA9W3D5JEkK8ircf
cvk0Ifl1321r5KrsSZ5xC10MfeUnhPernHJwQGs2SIdB2gJ/R8/iDIdL8iHq5mk0
CXDUlLGU9P6CAsibaBO96CMBQdXz5vbxC7jY2j4XPSwsSWma8UXrX6BWQ1iGso/D
sTApmND7CyBZBzQFsy79nVCkXi0G0gvPD259VZjHykDHAPnPvseDNkP7w4M7mNud
ePzE0oPyKsoTzFPXRLt1NvMVn/z3H5OXuDqUTyFuepPdVeUz5ThrnKlE4A+tMBFL
9nKNDNokxphxk1MzXpLejJnUTnCD9jyDEGgn+AbU/QnqONeS9aYajq5ME6s1BJHI
z9dGLwvF6iMURgDdI/5ceWFWgFUr3anZIbZUo3CGubOIHAajUe9A+9/KVXgRWqX2
Y83v6ZTYui5L0DwASgNw3+tWC3h8rQcAZSCaHIbPFim2b0sRszCzA+BInTZ25mLq
Z2S50Wk07KN/3sD8VLa6XMux/ER8L8yoieNUaFW55VtJ1yy4J7H7C1LS0CujhXUg
GZPhBXAinn/hlXp6b8e4uZqD+pF4bidxbUEjrKavqTAufeTfQF+QMJAUbxpRNbr8
K4M6IAwFS2RX7OC3hcMvMj+czX85KAZ947VsYabser+BGj6lNGt2CkOPhLTazEjW
mblwuIxYfnXGHnMDe2EQHj+KLvRhoQipi+DtubuTQ+Yloai7L7VPYW8SvKUV7Vj/
YSTC0wWnRrl+ULU9v4GaU/WFnUDhXJzilID8N5A16KrMquJjUWmXOXO07P8R+nUS
uVT670yWIqL4Gdb4jJEutkYA9quAuU0OSUQXyc5mAudkB32StR6tVyWB7oqLe0BD
/v+ZqL0NV3MzFEB5K0L4CeM/uHbslp6YXUO+uugB1VQ9KQNkbzjqZvbbQO5P5VaB
uNOOXb0QeWPTpWJgSpQBU8wKIGec1tq3RXjK/3bxRSUNAre7z1CTsQXgjX1V6oVx
QRMRL9wK3dbOLahRKWT0yajjDIrmL4BW7CigYFV4SDmrZ+J8XxnIyLOdIIq2Ilkm
t829IXF3GNp6pRP3Mji/gi2Wswp8DPe1tsqNkitxXnq/fy3A5n0ioWPYaAk5qBuQ
bfbNqwHddnIR5fMdYpnxChxbOJAzVZBjV52m6g2EONa1uRVoNkaLHTMe5Zkk8P2/
yWIXW6h26hd+LpQWqaJYXbYtKNeG8cZfYn1vFXvZxj5ZNvkTCbs3QxleXcOwisUl
wiw8/FJTHynjOXD1Rs8JOkOYec7omTOIqYcmA1tPCBb0zl/f5jxSbBuuSMfi64+d
+SSEfoq8jRYwId+JVj8DIR/n1DhOHhBkwwd3vnN0RIBZ7kU6GpmBq7X7pHfkG62s
2qg+PFugiQ9vbSde5m4yJIJYKnDTsYUYLFd9/hlF1ENNF3WkI/94cWqsgOWBOG8n
yRRTf/aBiOnGYYJo+k73GVOnpnqEWpaw3taIKDrz3fyIzqwRG9Rg5u4gQ/3DHhld
zSRGZP9+/zKriEKv6g/erQKh32VIpKAt0tiGiEemRhfeR3ebDWPeevvDbQHeGt1k
5HSMCT95XDBp/sXDTb+KEGmVe+BuGso+bAyt6x99GpDXz+NxqTAC3lPsFUvRavnC
dJD2MOL0iwYJDdcM1PHYfh7TiGdbW5Ri2tXIeFk+BBULtjYKWHvbPG0mQZJlelV1
bfpE7fZpwEMN1sGR3mEZtvKmygsyrI+4X+D3lu/qvZ/J5gLexs7Gaj6bWg009+Q6
ful86PkltlFEcHV2TacUrQ8due/HRWqWee1VaTAqDBZR5uDbenuB0JuJlFc3PQZj
YBLfcTesovy81wN1s4mMkphKMQBeSD6Apyw4/7BJHhawRF7BLQdcIVTygA68fRUU
+NuIZt2pyJbqvvbK1YeKHqM4jSePP0TRIAxX0aHpjJef3nzNaO+/CuZL9hgBGTn9
CbpaTnWLGBG7Me6QQ4aJtGAZ0vykBpeL9Am1Wqdp+4PfBmrE7RxwEBY5bUcvv+42
185CyWvmwrCuWSG++jmry7pDUSQV1ORDG53Hvlinm4UhA15jXF0pQh5KZ5omvD6J
wqx92pSMJRoQxS+8CjENmBsB797dpRWCeJgnebL7ysIlOoBbFrFWh+q6EkwH2lLC
WEGK7MBR+7hwAwj8s6rYiZVnXxptSCclK/E7kkp7YvZpMO2oMD/TgZniI8HVrh3j
hHScZZCEVnrkYTY1NiJ2msD53r+B/aYOIAp6gUxzXikPI7ZtPVpIB5nRdm99EYzK
AtW44yl2Mu6jAWgVeHvRJYGLwtdPiWB0hAGZOkYPXD9u0NvaHyhsWZI1C9vb12nx
780Qfm4yR2fLa5arz2C53WFLqxNkYIwr384Wke1byPDt3I+LO6qvVuAUMmf44HC0
mJ+lbGgJYF+ARhUpSRNsnbB3k9bvMj/j7iDUeJGbgXEgSy65GSMISBTiYbq8U4CU
Gnwer4BlFGtWqrCyAks9e8vRr/KcJryCYcDfY+CL4iOVUjDXHc6E7qt9erkpQOOn
6NPESa59SqCUHS93IwEPikvXV9LcH4kU1vd2Ehruo2a9fWmUjI0Y+25SMhVQ+EzE
bXf+dylWS6CIIz0QFmEVIKXyn9gJAomAtbm1ng9Fp+nnSKoaVgcSUa3iUHhh+s5z
jaU9/VTACeSCkS/xBooZsn9nRihNda6v6MS0hHTSKMvPuVBMxnUuaa3TpBwm3enL
TqcBbsOznaDUpGgocXzjQZcCHZjSLlY2hqLssLw+4wfDiu0yJd66s1dShiPZQYya
z/AZRskZXoYtH0uVhRm7FaveE2SMMVlNFbP/EXxPwdFfYpQF3GaPLYdN74oLXFGI
c1EMhddUJUyKtVMuFGWrQ/zFbBNbI+09wpm0eTRYqIF1zF3Lkiqm9PtMYJxOTQXf
r7dSK9OtfUu3ZPhCu9lC5CkBmuM0j3JyGJxkqgnC4XAtUyaS+hzPO6Yur20Uk9T/
F2jeCfa4GPk0uJlts1+TLVgvIrdhMHKlCyb+zZ3LB5Sisj1VS+/c3zXcxv3j8SNG
ebxmQ3HKZKV0S1MavH6V6cHTX4viYrnG9eJMlfrm02GHN1XiSa+JclAawpbl86ab
UpuK7/jx94cyxaeLfSiwa0FCL7tHPKJrnT3CtGrPvCOClDUw4n0YE2WY9UTUq1gp
8oqLuoyxwqApzLOym0YpThU7zOgYVI7z1B0XyjkzeLBE8VHbnaYAGJMmQmPgGNwX
tx4X87dzB3Eyh+210lHXABupU7QgrnYbnY2lu9YD+ON6jfmXZAsoUdMjj5cCIPLg
99JbfDgQR5ghh2bWfihMWUPf7ftaj3qCO7GtnuKvUp1MKxdRk+UyRV5k/K456glD
ppIPXQNxVy72PoIW4shnezOk6DEliR0zAUAOoe8ohMQiAJH1QgyWnpV87M/jrHxB
hqzqXzUuZz2V0oQpNhHibLDHsrUfosEiA02ZBGPubbpK7ov2/E94KjM1sVpbjCgK
pNjOrbj+s9LvhkiDo2CHmhj2k3ChCV/pzCVgEBZTlOulDc3pfecqwOdHTAzGR1uU
iScV86m3cyTjD2GObZ1mGX7KU51GIu2WKg6JuB2FMlFuiEwYI51C8NrMNKsrVsc7
NAMDNTIMFzGTn6F7jNVbiDSGvLLNHB34reoBqs/cKonAYL3oFhmEGiZmhJYpY8or
RIw0H23szRNbR0ljLnl/Wsj5ST5CrOVmizdnlpGKzrM=
`protect END_PROTECTED
