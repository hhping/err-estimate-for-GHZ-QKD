`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9jqgbjXQ9I/1f4XKrVWMEHbNVFLxsvm6DqoMhpwJoVkzhrScJv0BPOkthsQ53vK
SspYRWOd6BjEZnJm9qtmBlUPAJFOFmbLET1pezfdhrGmQf/1VWb0+5B+MDzGp0yD
BEz7XCh+xP0PJQD5Noq2DTAMQNDX0fbubS2ijZb4IZNbmgiq/Ddg6byDpjYBwPTO
FpOYYhqXeyt9IPxOjiWn6n/MwHsDyNnRMDDhe6UwkTlomZJ70AZwYYXrbXx+m+Zq
rD3eRzQmx5c8C6OXTK4lric4jX5b02WofmhMfeb6Xw49UM6353E/PVf6wi9WdQuP
yKasjMyJAXcy7SWZw2yOxG8SmoIc5vf5MLYR0cQsOslsjrnTDq5jRZH6ANF9p1Zh
OWu2ULPYnKAJQvjYwoFtTBA6pQWswIf669FY6ezJmIkokClyNxpGLZNZxsGOGMw9
6b1nOVIHFC2+IASz4qlb1gs4jy8fciJCuk0Yr/D+we+r4JL8RF51yQikds9+PpO4
WyAUsqFhV6wqWEB5CrooLFc+axDm2IUBUCCXgRVFkGTQ8puBzcf4teoOCcG7T4YP
ro0caDD9ppQPFvdAr5XKqtWTo8h74iOXvG9p8GNzLzVcxxr+4rgJ1+oMkIP3FZET
pL8UOdAz1Y+6bFaw8pfQSbnIjS6hLbKaRozJLa/FJhtIydxM2mtdcvUf34xzxiFi
gVeN62YMU4jNwqtf1aMdRLc8aFkm/nXRqV++hdfCjXPPFhGNF4Xcxjv5HTUanI7E
n2Bbt7PqVCyVR8jq6qjne/eo9y680MHxON0HgN25z+8C4gY2asVVPhwnjuWEOtcM
nbm3uZLY+1cun+4quG84/0Fcawes/dlTIHR0mJVCOKIwB8+xBY+AM7ITHS+65THP
EQjGbcVyDWjJvguexT0Er5LUpHlY1trXAQH6s0s+W+3B1UOY3hLFV13WUScHJI+n
0AAwJv+7TDGeQKCTPgB0WNZx/niWI4V68U1fMwjZ5IPXEpxy6kYG+EySMuyaMH9D
tj/cbgzTNMrz2yNYcscWk0PJN/RWhjc+QWsgDicpTo9R+mH+Hx6hNKXbkWU3SYoP
WCSJbv45feejhM/Mo1oZ6XMWfKpY1Uw2VaMzoBJiAtmglqhKuPUzMn+/0DEaiJ8E
o5utmLJNezvSslACAaXii6gwnmEBgxaMlvpV414ZKiboQc4kllRiTpnBd48tf9/v
r0O8KWdyrmrEzNDwkaaa6PcAnqu+Hm2haSSg3OjYp+nE+ZHeXwdqbWJWmNwa8e8W
IgyryN9J4fHra4uYSbKSn5p4viYqXCfBa5+P3IVx0Ryvptzvcn4pEM+uCXXHsp53
/tyhfW0qBbM2Jl+e6aQfBBI1NSr9VnWt0DV8XtvzS6uTVYSUxKdUPug7f9zrycp6
lyAx8DIAd6e3Cw0kC4LLT/o6UomlruWKSH/bIvSNd1/b1haCYRS3rNgDyFa1nT5W
3Lrun9epNpIhpmzOzioiNe0tF7qpFgD9GenoXToDpTXppdavJrju/YKWRdK78Rbd
sI16aX+xqj2JbnouN5co+RFW8p/OE5tmEJpZtw+sgfurdCg1tAyFov4hDgkJ6NPe
UGUZENT4Vg9sDS/wjEMgrbuGxMO7sjYbSCs0wD0zslSwQ/i0pOGXrrsiRuZ8Y/Er
RaGVLbVkZLkRYbGRu4iNxgepEEif6fUpdB9EM9fno20QvkTT6Te3cbCo+sCViSvm
/9PKG5kgKfdzYMjX84fX2BKK2gwk+n8Yi4igCgJWFZCtni69i75he1pgGMe4wcIx
Lj5QMLF3WdYOAukNC+yZHUnptYWIrQfKmGX3H7+2PqEfiPDos1GfJUDcg29WO1OZ
WhsiXk1+Mb7xPbgNa2c+jeVA9J7JFuNeELKVpwdRwhcYGvkh8U4cw3ulw/O9bR3U
/hElWHxhUUa2zl5lCBrxDIIhc5XXb0pgkBW0qRKvc01Y8CEuDPT0+NnZkczkhMcP
K2F2uVeo1dQ2WS62SKbBCa8uqUPjp5V6tJv1TmvmXsGPO50y/fCXatmXD/+Yq9vB
M7Gvg2IqIqsdG0/gTd5/bvg8f7ykxkZnD4lqEgjh33ZwBJz9/u1WyxyG3bY6BKCb
azczr+TqKRppCgN26E5C8IsUZSMbr6y7RE2I1W1LSDT5AGAfiWU+QTnZUIgifes5
01qd0zNcd2VtJqS0VF0EGsmOXkM+Kr2PrmUxdZRy88TsjfWDx+CVzkog7UVppPzx
T1sHFvDUoSz3PuA7vHHqypnBJ0fisvVGb8apuLglRCkPJlTmPAxUi4UtjfYqbJcw
90mgvBpYEYFd+X2JB8Re0MS0rAW+GLv1XsbKdeGYspoTliMC247/QxqtPnOYQ8/5
w4kNynEbjUY8H4yz8V1FHO41u3kn2oGhK5N0TVA0B7IRiUa096ICMoPURTyvrRce
ta1H8FsP4mzEPJESm5mVM5Y857aZVPtpfGVCRIzTw2RBIDXwhWQ47XAW+w4ykJxt
iJ8JaibwD9FF+klTTRn+WtOFht2ZAraYj3MRVCyNrdJDsnnTWCC13JK3/c+TiLOt
Qfl64OgNo/vrPAYrMYENOrjiwrjBP84tvV3M5mDADJERC3Qs65piYWRZevGZRwHZ
bC3i8sAm2yITnrjc9Zm30YOaQMI7PLe4pV8KUubPuaI+GAyjaPbJIB5gtpamuBMR
tvXigsdAO1Nq2dqyIxhTrIHqGEDRazaBjcc9EpbEDvSO2+nKs5DUcbd6/t+YHbh4
TJntVPJsTCQomI1MVgoIq7HbYP8np8kECLk3OWVPHQbxD47jmPjmnH4TxR43I4Vu
XWDxPasSLneAKi7oxz2UABwuQfwHmFKWH2LM3aIVT6XMH0Xw6TW6/VG8MMqWNh+t
W0vZ5KjaOr2gXA5tzxYpWTxv/N6xbz7HfrjQCmP11SJOzQLolOGtjXd+ekEEk8+/
fFfisZxtDgRoaM14ZbFMBnJ2vm2lbM5+4hDG8zttJu1ugrGp82kbXSDXyV4dDgU7
ncVROXNwyGl+0xgzBLqgaA5rLnWD+EG9DjGxq5ObO4dw5NJ24GaEFOMXfa2MmzHj
CU8irHBhfuNr2AZlN5mhj7XS5v7wTHqG0KSD9ZxJBTnhr/atxTFhqgR0rc1un8IR
AnXbiqF2STH+1a6VTlu+ogEqahxmpOsm2nc2oXHwXnnBmD5d6vJCY9a5+zpcZbPW
a5BS3wrMEViqgdmcGk05bwZcLD4/1X1gmtmX8XKXLK05AG4LBYZwzuY5UC4sZg7i
g04tvHICS7EeGR0C3RfhJ1o6q3d8hxEUTjI1hff0OlOWdTDJ51VY9iz2hNOCS7L3
FgI8iGB0lGyS9kv4RIZuxWhMTsTbVJXghU2FmEBAlH91hGo85SJ8C0jo1LeGYAak
E/64EyOxctdatNUuv17UQeVlWzLEYiLh57NG+5EnQDL4M5818O4Mu7TzdpL5LMkT
HwA1dS69TjRaoJ0c9TU7WkEFtE9utQMLW3D0IQTx0RAWeOh2+xQbRME0BFre5sN5
NX9WLLK4MzIlhIseOVjAUUqbMiEDopBvHcCha2ZqQGZovemsSptaRacTKtznD8F8
lsJbqvzx4JoKqfvayS+WulsSKFmzrr/3tLhsBvA3mvU1SVxeXJwWZnVBG01gEHXE
RdMv4AGh/tEkU19uz6t03iZkyEj1g/gdTdAJcj7995GYoMzqf1hDXeQjalZEmTji
pzCooNKJYY/0dQ32VrfBBm/hattc1HzmN7Gda9XzANE3EuOdUwV9OUgTJzKyhTAa
lOu2pg4gmbg3DOSjEqyuQznSz1Gp7bv5lAs8o8yCfLX6hr+EmAB19KB8VgxeX+4c
200x67vhLxABnq+EeMtDO7BT4nI/0UZ7R8qo1QLvsOP0bLCWS/jNAPuz6XkZoO2u
FFF2oZq+DZ4QpTMGzNxiQDIG9C7ZATc2h84IbvCPSdhY5WBIss1oo7KOnn3n6KFC
KJEMmGmNvgYHG63gT9vU9C0V75+K6i8T1lImKakEG1+wNA5nUs6UnAGd2vYUGW06
ZchKSiBytEGonxqn6T4behrK3QLGQCUnzS+I/ti1gz01F78vpD2QfVYrrOXRAc6X
itdjCLdW5svtqpwMlNE3pkXtv8oL260bcMAb8cM9zVx3AUOeus7HmK76FTdjhaZa
q1JMoOIl57xBBUHSfanVQtdLvc1VPXZ4fJHY5JiGJjcfJkcnWeXIfAzFGxoLyo0p
QgCvOytUyvYLfIfevcyx5/avWoxMW2hrDexvUZFWQmFlLo74RFAWbs6TDw/SRzJJ
4/5sV9fGCB1ReYptxgKthA==
`protect END_PROTECTED
