`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3aC+OhICjdQtzasAho+nY7fG3yRCVFiDI6RxyKFG7V9Gw9Lw9R7B8U94meKO2a3+
vHXjsW0b0Npbbh38BHkKj2Og5jHnlq3omd0ry4uNz88MvG6evyLxnfHbIZoxPlgb
H7Bbev++6gIRt+8NyKrGvXo1bkVqkPVzN2a5iPaC3VeA9MGtqKQjoZ63IEqS3EFb
FfL5rkIHPzvoq8m872SV6RT5LJyZm7ltoP2xdKYniVJvnORcyaKPsgrJa4HLNhH4
/YXY1auzcVHLlMNVkU5MX2xcDXEdEVwLKwmXpwtB5eYENZD47fJUIfovS28FZBRK
8SmQLFY3xHpvMF6qBSc8fVHo5RFhRNB4BJjSYn/pzXhqHny3r9Dg3lf7nqHidtnz
heiZfhpMFDQd1KdrlU6z1kgGoL/xMqt/t6a+xtrbxTo4JQcJoJ8Khco5CsaqbG6h
2bSIyjWgF1I6prvCQcYLTirFhmslX1Ajv/GeWZ4vEyDAGij91sBSiYFdUPdejYpj
trfb0za8Bhk5YCnxYzyrNZhnCPu6Gxcr1Toj1xxN3a7X4uKNMC+GFwTJ7t/FTMnm
6XGolNyUzIvKApSRq8eLRMYYvrvYt5zImJ4RWwAba+rGMLfVTF+BfXVfY+fZCGUs
GXZ9+CF29wDuT2dOlpCzwIuDCIY7KCpjnvAxvj/Mhk1X+JJlZhgdoFc6idQsaDYJ
xuHY0jFXGxWgHXC7E8Zcp1/w67n2B8aMjj0yqoEM+/X56ry2ivHXCTR8OiimPkXV
/scOGwTmw7tNiRzPnkZiI2JdsZ9UrIDvqoFmqchDfynQRJcvYgxnOXThKy2/iJq6
5EaMZNmLcTjQktnijLPpw0GbszUg1+Hengod/EpSYPmBjrlxi4a5HclSKMJU/kHO
FhppmhwQ4UnXbxoZ+Uq8Kbp0BXePmI5c5Xwg54e79aJ5NppOysTcaaOPszdDfPfZ
dqo2afQxspdlDAt46rgpJqga2eCEwURm1wPudyeWBAhmL7VMyNJzYsQpJl2lOubD
2vlWDD2gd8U2ZfNUYJZsdTWe9H3+gGpYl6dNz50AliUrakPGACtjSDDBTQU/PPaA
iOJlbZTfCJf6ej90sWFSyVvRRXlqWbW+XiLj41rb0VIulom3WyD8yqTLU6P46FaP
2vSfWVzMVjpensjwEq5qPnZpzUpgDU0iniDozbsavU2JLA6er7zgFyHDtIMxj4CN
0Nz8jK75nSNLESLc6Baem7U+gIfRC/15tczKPnhYWCbmgGzFZ4TzwRur9byqWXKs
yPqr/DJ6t6xeWNT2kRKykFe/qlJPB+v5g9/pqERp8Hb2cPzCJlp2wlIk4egeZuAX
kl2MkHsB35EsUA3SEx7Si/KDfZKgn2zg6UgBxv7z2zQAvqqZmu5D/6abtcVaaoq7
AFj3v2faXmdZX3Me+EViOusA9pFSb/LH2sTaGoafqtou+DJMlY0GchzV3A4cZUn7
uXg9IzbrMADDA90thePQeKE3O4m5/6tWa0mNgUG+bgnK38ePKqEcd5D21kv2EvHM
15G9gVwjR6CzhifJxTnL9g==
`protect END_PROTECTED
