`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tN1RKJakI7gJTXZGwEUPQ8NN22kv+U6T0AEbUAIXBcv/EH3nS8/uzvgvmvNqnVwM
dAuas15wdKi9n/Ml0EckfSgol8pzSqtqGtMnD2YyoJbYZTUzHR/99qO23T6mN2Nm
i2RsAGv8hl61Y3NOA0KOpvonIphKxWBbgcrfwqjMCX/HXD4Ng/t3K5FDmZ6lClK8
qgAAvM1yzvaWFwvxgZuJ53Cj2lzH0XHDd5xiWc0EFQBeRCO/nhwkck+aYl+vf2Yu
qFAiXOpJZB09qx2iAkknRbSGhz+nBTRca3uAXRjkULWfjaLVIpyY6afJUEGuzTtO
D+aikUiJvSK8LKrEkUTD3jXR5WppapPMKJKfgbGS7IUtK8nsRsAQgsa/3oq6P1cG
UeJCOpxtkHkjoxKXBTwdy2v+j6DytZXn71mThecjgYnI3O6u2enu8bqGCr8TR85v
fjv9EAU9RsH//nhOrnAhzTbO39DrqJAtG2+bgIflo7WjWWoULAB7dFtBaC6bnO2V
K7lNBBxpCQBIg+uS3NWW09jrQILi3XyhCBporbw6ChgyAYSTQfOeRfOgXYfp7H7g
N98Bq6C11+f7N6UemeFm1ofSsTXE6kTx9RwF59CwQblvD+ryD5h1Fk7F0swAT9nL
j3QPMGlSVwDVOXdQ/o6ZC6XoLFEAu2FHtP8Q9rESA4CFzQnU7jwygoRe4e66yL/m
qLRLS4JXV7NH40xs+pJveam/B9Ss0gUz+Z5X53k7noaCKg66CrGKrOEoXEXn7E7t
koNwI16h+vAAkzuzb9hZ6YBpMWcGUhoxScFsM06h7NOS/c2jdEbL0p7vAjx0pxt1
k5uuyhqBUprdw+wYfwn/aYB+tCiaPcp0m3qBZMaYNcfoisO+MbLxLPHSnDt4HhuK
NQkPXL0rpqbuCasrlps07wKoEVTGqEviOwngKtPbh/gloqdQnzn2WBsl5F/wgYk7
0t9HIJ4ODKq0cTd5NKaIMlBytIfMIrvBeZrE2N9rqK1TkS2TxakwJ3AY9RwDwDH3
A3JK9kOrMMcni8IdhRilKga1Q/zXZaXvDkITfXG1q76fAdhASrPxX5Pvc7Yv4WQY
ArYoXqS+kf8LhChHWgiz4OMQ8bdxkBL7j5627eHFOFgT+2dUY16sm5xIl78xb81N
Ee5hxOYJPUr8CI92A2VfIw==
`protect END_PROTECTED
