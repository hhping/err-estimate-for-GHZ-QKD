`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rp6Gag9EbRpVlZI19wBSs2c4G/TvYKbizqF99wQkc7M7uDGalNSr35u2xpzCcUod
w9TKMSkxbsK5upS2h89tfGuNCzWAUzxmLmZ53CEqUwgH3Uv03nxsW2eEPtVBoWY5
IyIW4NNAn7J0TxqgKH7ELX0jK84vqA1+18xWNL3+BhDdix9HfUhQRPw6LB5q1ZSQ
7DYZkvTURC4nQjE+BrUzrK0HDqkWzyC1IgzQTKq8VDDlwNSgYZrL0upPHMq5mHBr
FXa+41JE7jPGioyoq20Zo1yBhQuSdobKE42LBvmEwl0u6yf4yuUmHpgP6FWocwtg
jQaPriQXNOQr9TiNLWSa3IVRuXCKlA4Tar3s3jITheRdKZuLx7mdFPRRtl4MRYzo
QTVU6l8gXOA2KO2tgEIbzCgxM5YJ1mbJhkTILUINCHGOclbjoo8wUAFSO3q3vQpe
FEl34mv131TsJOXBxqyd22ZD/f5V/H7PrL/1sZQHKPyu75JWBhsi92p+JwnhXSEq
LL69kdSdDf6p4xdqoM6croFRP+pJtI4VUqyzmin1fqrr+O2g3b1yeG8ZJWWx4xsv
rrjXr9POIDHdypqHKJB2zj4cVT1unxggNWBrpxeMrsBRBN1N2YZ76Envf6rUX6lx
QWpm/itJ+ht0U9u1yij7CRjUyX9Qyr19MppjJ5KKGBBTX/OqqEkxcaHOQ/Hfpime
Jg8CZ4TVmYhvfyUkpIMnwYRzrRINLkaF8NbQ5Nj+Oexys01sQNNvI3dj0MnNgXU6
8K7r1pbuAeBIDoTHjkaMOYXT7rQA1NufA6VP8ZyBH5a9x3hohh5w+eYWK5fxyLSQ
6YYijNRKxQcVMqhCuv+G0SZDciudGkDctA9qCV68ddEYyPJKMEYhDaVh969P6d60
wE+36I3scTJeuxhFcXo/sfQ0rL8vs7b9sI1zqD/x5dbQX0qcZbmQcyNkhVtRkFkH
kFuZdeg9i3HgWPy75PBqHYN+3dhKHOXX/gkN0X67WCJg5SfgOgKqSdQb9L6YEBaY
Fkfeal7iY6TTJi3cot7cXUbCOOLpNZzP5zqR0O0/IN386k2VIy0c6ZuexsJLIk6y
rdGYZmzgOj8A6yfm3pvXGw==
`protect END_PROTECTED
