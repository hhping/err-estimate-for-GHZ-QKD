`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYlzYxXmoX3/5YF5vAIhb1y75tAawIJKGqCwa5do48FihFk+imzjo8TgGWdJWPrQ
bxsRI8M/nbsHNn5QPCleWxltICI/cx4dOnpTTATjCAuFXUrcCnSeKkblX8Qr36ZG
sfGC8V00lAr2zLSx+mne0ZdXS6KePNMgpywb8/i0zE9VfBiJs6dinZk3vvxF3Ub8
A9eFUl4rHOAOG5mFE7gEvUz3vQCsfGuqyyueXd3XjYQOhhFKch0xW5h7n6X/kaf2
FHp5ls13GqwMR0a040tuA80VX5NA7ra0XaT7GLgWFUR0eM5U9XQRWn313SXcm9BF
ZIMGxkFa/Jbf6YdeV11ALdniFJoEFTZ9hYPZAo3Qw1nvaO06pCLZ9uh2rtzpXMSG
JGiPrZ973+4U7fWmVCfB0gNXebhJOxJbbh9NnUe7p7YTnfbSlkGL9K2dlqY8uRnT
yFDqb/M5COaaQ+wW2j5z2WlNM6Vo+qGdpq1gRKUbSR/WQ4b74kefPlVqzPzUYwGp
YWVjXmlaKm9WKvt1jfQoQ4GKENKQ+0ygqDoQTYVJyClVNnw8HdhUtKVg7wwTulcC
Tqx+CO+CrSex6Rthhb1xA1n91KxOEzWhsez02IRSdx3Ca4Oglr3A5zSi9Ep3bNhS
p1wiE1+rTVfqLiycfbYTkh/KV95K7nOeuF4ChKxM1VjsEkfyp8lZVNg7nTm/c663
uYi1cauU1sJbek1oXLOkes3dG57JT/y3YCv3vRweinHyrSNMTPXzZCjlRKKS4UR5
PXPvr21V7Lv74uX1FD4G1mhmR+6OtJXKVNWfNaTJEBPUYGuLCNz+vb7wvhljHe0s
iOmdzKTSHp0G8NvQRBBaS94ijPhVUEXUqQqvJm7AsIAYGtCJpyjeRaVJu2QNPnTQ
YcAlqEhfVTAvR/QreuIe8Q9s6P9+sv+OnRc6hyD55bbcfj1DqO0n0SfesEUxxjCg
1vZLkozbkBSg3I0NnNUItMTeal5p7gQVAiN1gGI68JDbVUDEAUSdhuH/2RL070PH
39AlUwC0zd6iI0EcJIHD0FuZE/m2c4soGq0hhwPzuR0erybBMfoXwmithh4HXeRA
CjgJlNzTXcDbKxCPXaAGM/5Jm24MNzOMRC+gfHQwhHSEF+dYbsGXTHac5yquACPw
nlzPsvhgBaN29PuA8WKp3FKKhpin8YQ0sx/PsXvcyciRcrRUSMc/KeapSIGmOTgq
BW2YbLRZue4R+qp2ZukA7A48tqxIUkV8Xqj/nD7hqwBw8QaZrBoO5kQaM39A5+yl
Wai769BhRXcwGGY1zks8Vf8WBmSDhe8c4jzLaMQK5SxWqY9Thd55W1gv2w25yOXj
qMWNb7RFIWvyERp4aMTw5dBwBN6vfAR7UmaNg9G2WMgatgF5B2ZDnbF7BcbcP4rk
GaWJjK3vKZ20E59xUPaKKWngAqAn4eUZPZPIB7KESpepR09B2M7GSmxo1LzZRTho
YhSOUv0oKwnZDxzBbHywwanOGoLvnKt6R4eGXy6LeUhpP83cWb9pOcuTB72H14Vd
palruSPAGC2IJ9tvt9jIQncOiXY30Aqxc6CKuAe/M3M4E0UrlHlZQNef30wBqtOl
JxRRiLCybQLkA8yECW327ZQv0VMU68tNuDGNqvtJilZprxShLPU6cMDIeSuuU5lV
Bew3In3l8YhpAar6JQXE+Pt791YvZ0UF4K+nUcpGY3/VZcPlpLRUevMmSErlaPE2
uZ5EQXDdzxv5WF62XotmsEt3uuqSo4ysGPoQa2Hy7f2dzM4WqUyCY34xt4DvvRR2
pBczAdW07jwx0JZgRIZyO2v0dhI7abjpKCiDtTyey9l/xzj/1fRiA/ahFnDiJS2W
T7BUr6l2LbtZCR2Kin5ByltTVXyGTFC/tWniwnMOGw6Jwd1+RTubdHUeKi+MoE9x
cIOAA2dDekg8V9L5YK4lFIFqRgUMZUSScwJjen5Xwrl4TBtt57XHyuQedDe8UyJx
SpugQCVpN5/48v6mRYB0GdaxXyN7Na9kiGzJ8YtT/CIx7sMWEwJArgPIKgSb7VB0
KbyBTD+RNi1opRrJPU7qz20etcmXS5qU414aeu/j9olWYH4oTGxq5+2OHg4ShGSc
74mf1JZ2dYM98mfJv++o90XUsYWWNj9iq2TIY7X0FDL4nXocZR537eMk0Y/e+ZcL
IVeh1DRjOQ+06YrrmlP5Ju+nkklNibQpI7InHqC3e6bXsqEtAGbhXdAwlxjft6Js
tWipIjDymCuBF8QqtDs8ws8EeweP13ZqymxhKEFH3k4NUn9EcntZJcYJxB48CMtE
05WsIz/hJhkGN6xWmUeR0PlhUpdhM0ZzeXArQO6lBQgPyhnf7H/VWR9kgWrWLXOt
iU68J6yxSBYfsYIP4tyASXBEqXDwER5uTj6KToX3Q6Mg85biL0dbn2GuZZfRCkEc
CeNN5bbmlS5l54eA2j7SNACvIxGZFo4fPfO4+xBfsqmGFVlFBsq5viaR7ZRNk/q9
WxptfCDsAafQ/csJewa8cpbaS+ZtN5G1WdHAVtmVRBMKu7NiwrkTLV7a1yGMFlpr
41+zymX8/EthpuxYim4hDJpG97ByK8PjGbPZ+Q6VC1b77z1ySaJHmb+1KcQLXooi
fAjQ/ZiD/7B5yTo5woyrVPfdoORE/PxEvOX9sD6v3l+beNE58z9wszGdUkUaJ9UB
qkH1NHKjRgk0IzTGxZvshTRS0emia9yn1EAEtzjhyR+fFLyJnWbZNp22kSO+m/zM
QxnkaPhtA3IgJTnKn9C+zSpMof+BnZTOkG4+cRgqyFzOejlWjai04R6G/VNTK6Dx
XuNOx6XrSMGJsNQbtrTYbYmqUtYkh8SMw9TOHYE3VGHN9AMtVBlbOULCo/C1Ut+7
1neTKOfY27Vh61dAW/kYJRqgaScWQWdSxVF9+t5NY8Eu2JGkpiZd77CmK2+xMtLS
xmOP8pAH48bXEgBrr0GUSpp9MavzQlBFsa/Wd/fwZjgeOXWYWWIjmzL7UCU3hTWy
RU5ApbueWuMt4VH2y05+Pp6fDkdQzvlY1a5QwUcemvOi4hWs0Hr6ejP/YITGkCau
u8xJ/SnlKU+w4jD2f8T7GpgcuBafy5XycxwlAwMnFolo9PQXLPiyIY5mmJDefYdl
JowGSqgk5ONdp8CT9/8sLFby/1L9l51PY5HzCxJmTaaFQGWTCEoqkrVtVFrKzjmc
HD4Tq8k31/0fV2PITC29seNb5Bw7/uCLzC2pfilMZAW1T59Xr08jEzeLQqE0QmyT
iq1mp/GTCEBQqME4yQI+PWjK64g8hfPcxUT8SY966SWpugsqA2RCZBL7rPRx4s7v
vu9WYuLlUeMng5vGDysKnEiH8fl8NwtkNX+RbITvz+Qg50R0/Jq5M+JRJscFflgB
pFoUB89BNOfRDUczVsAcDT+77PEIenYm7/50x7Wxax+SZNa6uLO+qnT/JLP5k5Zp
B/PmHxb4WhAhMOhxF7JfoZOzAJs4jCV6OKva8HtExN42IlSmcwVgpg8PGj8+wZuD
FFZDdFvq9blQtWHOENynoKcHoyiufFCau/avPrUxFlkQOm9OOxSEOr0dWBzE039d
uVvQ2KnTsbGgi7xtybbNiP/6gBP2BXjuvyBkcVsXuyXTTRE48Lw7p/5vBfuk8LuU
Vb75SMfjHupKn2f1pVUT7BWnqAcqOjCRKPpFhXoZNiadfSL5RV0W23jrVGDEu18T
EO9sbCovBcTtoELE1k6BDEtqNULbJEj5+hle5NkeWVgBFg87X4NgODyzBqw74Ka/
Ut3aGcPcL2Kd+wGpnAer6N2uXgKu7W0+a3Wl82cmnJ3PgBzGl+tBz9FlloEoNEjl
Ad49K0K7Fvj91mJyu7kYjgF8LoFSAALHUZjBjFBEgSduOMKHhvbwfD0juwAWjfV2
Zspo9qNAgN/dvtsD8yAWqRFOi7vtgd2qzLhmG+Sga/v2K36/GfMdeJMvlLvrNTpH
jlVjMj+XyLBQZBALvp8kaz2R9iCRBah/AL6om585NtDgHf8UlTdV02JZ9RWy6oiI
2OTIYemjOMw/ACeihSO64AtLZSa3Cr91ehZJF8XBZK4XQS1O99rfAhrY7uB8gwtU
A+ymZEYPRTxSfaGQqwnziZL35dYGz6oL936VoG0wcM541QD8aXdEJ3RJqxvmyekw
wCu/n65Me/lMENb6SiAUus6/dvlxZoSSTvNt0oJVResTiTujV2ISGC8E5ttmf6nh
nCijYDPDA2kQJ4dlXCVwZQ==
`protect END_PROTECTED
