`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0NuAgYn1oj5Hzyu0dGdIRrqxuRMP328kSK+4R4rK54EdpCoDFWU2Pb5imgKpBqBB
Z7+HHcYnjOPZ8QtoCiLi9Viq3F3JHxiUc3i8OOkwI+jeiSav8/eWudS8+yvXE1Fn
wPvLH9EGJ3FA0IT3mFLaWqPC/7MH32TAZXLYR0b4sMCvep7XyCQab51n1iCrAm6D
WFJnstQsB7jlg6xh9esZ2JkiCUkZ8zXx8nlTjeAK2Is+mklwlBih3EqYwleDOdsy
flJEPJrSOnAxJNzbo/kVfwCntdirgQ+VubfXiEdFsaYxH9Z0iuY7IYnUNRq04mmO
EInhPHCRujLeo7D3feYcmYaHp5LYbaSFkR6+VbB/gHm5+2LFOts0EnAEVQoVNQwY
hi1NMxlASqsXzoDB2kZf5LRUWjHz1SnLkuwrF+fDTD5dpgoOTlty/Ym8sY7C+V7V
mLE60t8Mb7Vz43XgGoIzlvyp7EMr6oDn7Bb0f5f50E+LP+JDCIc8hoXqJpp8i+CC
Bm4ERtigGwCv/Prk/1zD17l6rdn+fFUKG/N9EDfwUwZwe39/ZicmpTQHUXj1wmYj
6p4F49x59fVUaSR3Hei/ffDGW1Qcr8UykPs5Q5YFzBwvrmYtRHN3UQrzz5x6HUqi
T4MKtRsJJSd2qo3/tlGU5Mj2NdfMg0e4KT+e7o5TC/T/JweOtcWZMNP6TV9yVi/3
PZH79zjVfOxeWETNmlHu9UkHogwecwdsbrQ8v0m2uY5h40qp7Aj8Yi1q05A3lD8b
RlUMANIQY4gjybuguntD5DcgzS27d6+P7++4HGzBThf2ITgw6BIqgzyK+8OnSJ9o
af9mRx0hvxpMShlHO5anyESDjKdm6xIJajfPMmTa+jAS9mLkvNVYgUuotLU9juBD
mMy7LMD9ISMtP82IagCdcZ8haZSSRB7Dh33citKieOZANBmsPDhB0bCPX0KMI83z
N2W2gYpl8EYAM5o8YQynsdYWTQGtlCAm6VaiJ5LY02RqXTuzvoYY6NjuWLLBRd44
37w/WnHniFblL9GAbihuoKxNqR+9BQ7WxStj+Za0zz4RWP5XmX5rw9vA/qvGuf6i
4OcjvHFakj7v3NEwyNvfR3Dx62Lb/PjMwsnONHo8JKpXtLKmtHTtqdE/B0TnC+/4
XmvFVOR2JPNXjY9cVFcrfUo6z8LvRJOdJesLURqHAQLaxMqr2mWV8smD/1RTPVAH
o7crK2p/LeAQzVjDOWX7lM7O+p+QMV5zq7tubnjis1LYkhYTK4izgrIkIbJoo8P/
XMfa4CrN7KC7WF26JIoPUvfEmFaE1tf3KfKKaNbEvLrET0kahXCCOl+iVr7cK8/W
BS7f77w4zvtq3ZjL3Ksv55/SXPmBugQeNNIbCgO37A+2A4qd2RDl/xBmTWynFpLH
Np8An+o0Al1dHbbo1T4h0rAoqpWhBuiEJUJnep9Z+HSXSQAVP93/pJIRTuIlsee0
iAJz7C3Mi5NcEVdjMkfoTKKjDunf17yNiWy1O8T86a9YwLNC2Bu/VQLRXmJOISF3
OHwEnasz6NCji/K3PPVLSN25zuQiREIo3jYH2lq9zRW9w8n3UuoiEi+rQCJWqsQM
gQtAsImUBBzsuq50bcoXuuquJT+RRGXt+3bYI99f1anREf8swL6smG71U/lSnr0P
7sGvGp+5G6JogT63SinwUaF3smtes4cLDMBiPvyU4kzI0SzuGDn0dL/UfsjSM1Ye
hMRrMjCJ0YmlIRQJkRDbOtNVGNnjnjYKWWfMso8PbCLK6iGpu8w3KEwj/vrq9dUt
+PHx3aWFQwGo7aiZKUy6Lo11Y/quHkUJav5PI2v8FW6irs7h4E6sbSCLEROWCjyS
V3AjosrB+LQeb3p+M6h7Hw==
`protect END_PROTECTED
