`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ywMqWqCWnIPZ29qyY43OGEOJsGmRuwBfAlXoqpX9TwTjIUt5qfufS5EKND9CAUqM
a2Jjs1H9X4ueQ6vSfS8Z8T92ipyWV/oh1aFqqlAcxG/k80cqlJV5lu3Hmnghhq7t
2BiIi2QLamvPxshzDoGwUcW54AZcHqvsf/eTwmdVmG8thf/cKxavu5JcZamaP3Lg
bfFuHZfvglkzKZpRZVP3eoB740SjsVl8PTovl9wASMWOiK7QVmNGhCkFZDzG8aT+
uZ8HFx4btEtttilSVAbUx+4ZEKvyVA6Fs1xk0pCXSVgU9AKYP3IFcPOb3PBst+So
BFemldH4p10YcXwrTw9LTlRlPm7vvn5/OaUtlD29SOEVDEzrRplKzNgGIIDbokhp
DruZAK/95jI3m8V9R6E/Ow==
`protect END_PROTECTED
