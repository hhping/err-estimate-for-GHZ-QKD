`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/52dCSeItcGWArHlHfaA3mDDkj2FFH70hVxZMnFKf5Dvo44I+tgqd6cAu/YL3O7
cuPe4GWzSOOxMmBA4RiRe9MOhJFd07bGxTAv9EM2spuaxQrl2H85jxOTPtZMEB6W
1xt9tGfRNWj0a1trcYuk/v181TYC9tSkUMmqi2KlD8DvZj7/WDO4FMfy/Dpz8De/
jme7shP5Hpc/LSJ9Zz5DpOaHfOs7XvZHznss+V24VZtnPEPBa9N82KHHQ04wc4bO
ikH/pisVaHASbg33krew6fW0LOuiiTC/SFuguCMDDm249dvbGQkpnqZ68UmHwlZr
oRBthi29QTMkZsW8/w3Y3lDY1stdHR9Q0DS2vU19WKLtAd9BarhTZkC9yPHdFYpN
/g1NfU/q9w5261HYmVswNLtJKuwDH0iVVTT0t9MMbWsukXPJlEQMs/NVq93IXaBv
7HPpQvuuPJWOLQpriYT2uxe2NCoUZgxxAtFQkUsqpdQEikW4WHbrc3KtxP15v6/i
xc/h9bOYlGak9wUtfI7QX805EiadN5BR0b0D2DNfKTI11RRyrjg8TZXrUDEhrJhi
GdWqFBX8ex/48IY9PCkt2YS8Nj6KqBDPKeQHOrPD0P1R/YApQWU5RywB26NxEziE
4T4aiTa0qVqm2veiGCvksaumbqcWpqb39xEJaEQkFbYbFGfX8bA/F2EC99FPnGmX
ydaDt6XO+0if+qalutdLcwWz8wXaoAvolr9hnOaacGegLHzJLxVIPi84rjl9IKuV
IaUTY89MXJSXvb8qV3v+qAs9fymJcOwFFQt1oehGb2ZuWCajJbKDD3TYX+eKdtC/
dLwEIUwb+Ur0CBJNTrl1saOQdFzqTnVa2IDUrZC3IXW86wdw9WI+lYHaFR8CDhfZ
3D+qIH1bjMjxvlNotkc2+YVPfnPYtBzgwBgI4xAf2gJ1c3q+OIsd3BJbK8dGP5Ek
6bao/O35jsh/HL2uapzi7T7QPdhDxZtEW3aXwk4dZPsPpi51WeSAFmNSwcjOldYD
neBnS/V78Peis/DNW723QNpBioL0n0NcX8OFkLHj2KWdXsak3775BvP+wiMmEJW7
UkGqdg8pCBphm/8XdPyYWI+jAJqKlXkswqogrjD1m82WTkW24DKrG34ENfrAUSn2
SHi/FMylBVa472uGsUhx0+tUWdrTSkwLfD7KRjpetxoMszJ6HJe6YeEezRXhLa4P
jpTtZzZORfEdc91WuflHk8EAEUz1MSgzh2IzH8KfEJDyFlEC7paXI+mxOPda0gw9
l3rEMHnqwmil5UP+1PrClfcDbAcaYmXafDiTfsf3PzXdny4qjCBOabK+r1J+M1zc
iWUXuIhvJoG5EsNT5VM72mbsdwwDYbD/N5h/IoUObALlFIX++HXBMUqhpp3QMMpk
FD4yPzLcMJLEZII/zpa62hZuNuo8Gl0gEh35KBVliMZgha2hZkbCVhEOYMyYoDvg
7LBe418K+G1vJL4OBqTgHUUeMxqmBxY4K5q8cM5E/Lh7PSee7vWGsBKIafeW/fEz
m08h4SJA/susRQOibdNYBHoNiFJKvG9EEudvKV24QV1WFFNSsLHEjhGcV5Fh4Zpj
9w9ge3FIhCoXRMApUSAWrv1OUKhE0FqUtduvvOl/eUoJVR5fQYzoXEfbfu/SVA+5
Euu1B5odY1nR7z7DpmluBRWqisy9faM0l1teQXu16iZk/Qbsb2SRbWV0BOqlVncL
dg6oOvNnvNxbZ9o66faNWdHPnB2/BIs2CtyBHttKCGwdeJ/9jR2CKBklZ0UUp68e
IwQhQNZs/b3MTDd7IOwKxwZhD+4sHax5/MydIlVWl36GnnlLrRtH4HZ+CdZblBEV
jNUIn9TK/kj2/cqeC1JCdUyumusrxjFAruQ6slFyp+FS3OCSjTMnqYVhUlyvr4OB
Pd54zXdTOvUOkAr2rXGjtUsUzeBQ1VYniSEr9/+hxCRnjFMea274E+wWeUETFMv/
Us+qhP+Lkrd8ZsOZBsT+HlwJcLduzQ4d9QVMvasUSTQixvUKkzox5u633zIxl0fh
PWd43tpI3PWRM5DinUv51xiv3I2F85j9eqHpdRg+SJJTNhIvMHbi52W9Me+DeZs/
qt+py21Y0F92ZXCAmaKwDg==
`protect END_PROTECTED
