`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ttVOSYbhiwUbRQ0Imqq1ma2eDKYFtq+vnDh4AzaRywO0FXAVsgNn/oqiGWYh2/27
+9By7GDScJUppD2dPg55M3tMeQJzrriSmTjB1WXddySi4DscIBTKQKOMk6UxmvZK
h8AikOdLtE4LBJADZkBC+7GZKMr3WKb8R3KZn6CJUdcfMGj/KTnKghbgU+Dby95L
b3UVrSRZ3ldmU5RJXOT/NiUX55GCC1BGy/klYu7xeUOCVp6K8qO3isaIWNb1+Dto
GIAP/5hBFCKSBqAvnVL2RCUPqT9o3xrFhCKyCuButGHyuWCIk/2Dcy2Gd7C49fUg
rLTttk6nOzWxzyF6xXhclvcYS5MmwlcB6T53VAxOatFv4Ru9fHQ6hVOWprGA9+oZ
ThVy/AU/kt1uEdjjfTWgD7gvsfzn8UiO+fQTUoHQ8MZwWXxJJzDTQIdazGcx6JEZ
gK9uiWXRAql+OHBx8hhwmwg8ZvCBhvYITAOCz4u56ouDtkCMrgSbkbnXPoATLFR5
L/cCZwJZdvjxwFAD80FNVi4zjZKjBZuYKxIFQFb/5LkI9vY9IPZcI4vhNp1p0P37
AU2XENMBPXZaFJ3aRJ4iaHPXxpauPaJ2/kCm2JpetMGk7rvJ+GY3rlsXF9fm5Ayv
VWy71FUVKG1ET12d38cQ1nlFCIyb2VpucqVak1z2obCW0BMho7gVjApO57HKlc8H
`protect END_PROTECTED
