`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BmpMgwQ2pPH0r0SpDYXdeUZXHNAYYvon72IooWuwbtuyZ0HcNu8UI45izHg89n8i
XXoRqW3dALh9tWww8D3tWJ9SX6dTnPd1cJNX9AQmsleilqxfKZHbL9uh4zhCEcAP
FMt/lRvXM9FameiOUYPSJ/FurfdZzr5nA0lgWk++hvnSPU4e/G9fiYHRn89ROwcv
7bV/A1ruEMXwHWbosZsynYE6YWR3ZhZubBXH/7aTEAVqjI2RcJv5Fbb6gYmGE/pi
zCb0CsnKYjxzgVudo8/AubLM7lHrzMXjBHsBdg8+OoJBHStuJzlMPj7hDRjQzd7l
9K8IiWMpqULvOT84NMVgJaSjNybr4rSCq0NUeM4T98rSWF2fKtmiHCwAlCKOY0BK
jn1ouDrNulH3edVXANHL/FD2Lm+moOjWWSFcl7XJBxnrMXYjGGOFXg36iqQdX9jN
972ghUx65r5IBx5ZQ/fvvR2N9DDkVos74LIW4QgF2IyJcU18VwqF4mVnx5EjgX4i
xnCj9z8UjVgg1VtUy8Ol+yy3xvFTLlwOj1W1b8DoZYah72xuty3+lkj6OC9jSD8e
G7vrxl8gIP64iPFan4oHKmPqrDZ/+SgKWQk9d4z/vrYLBWx03s/qG1jzNBsi5W5t
v5EooAv78Zs57q6NQkX24kzA9AdZAOczRTisbg7pMXsJem3QQpewUxWdhx1sGVGH
LTELH4YM43RfHLXwBKhdZ4fWSOcJWJPVEVYtFzAB4XVKRgC5oq7Oz13eOkpND17Y
y/hn8c1MpHlxWPcE2fkarh6jcB244n/3cpbKu7waIid44wOgy4TQOX2k6ntdqlwt
oxSunKn4zEVG4bxDSwT3FfFloOckEN6+oq91kqguRnc+T5QbG+0qC96AN5Z3CXos
IW2QeKC6d92SDIFPuiUA2PxPLzX8G1KifhPbnBP5h3hcA+U1eqWii7dkXMDII2SM
Xd2TS8QgsvAwZep+Mvsxc8ImNgNJGixjTF60c77UaGk4iy6RKg0OL031hXgYIYK4
8TnE6jkxUwlI3E1eKUWCocyejzy+wenPfIDU/h+/MiFIdDF6iSomZwJXBAkgEOsT
fFIBLkUeuKMYOmiUOf0t/yrw+6SUscd/CgqGg7sB0gClhiPefJZ07a6WwBL6euJD
Nyvvk4/eQ8IjA9VX/yek+rxHiA9ZcphNff6f+jGDBMN6enVf9yvK3NF6ZzGjXBD+
p+R/nUlYNoyAJDox3DIEJdaQ7CjN2sEdYCVtkD5l5VjzCPVbCf4/GwSt+bZ+9zv2
PQo2iMWN6hedVrzWxCT/BA==
`protect END_PROTECTED
