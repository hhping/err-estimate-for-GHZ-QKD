`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KyPbuoUQT9G4E9GpdtQ7PcsqqIkBOX4PVnfOdsMNLbcdWKPQWMgQ1EGk5SQP58Z5
aW0syn47NS8GoVIiVPNjS2VRx1IS9YSkhBCKUn8TiR7f7WW3liDsOuk6KQPNPth4
MSBc+1CCYQSuf59sP9XrEsHhBmADZAUJgwschHERUcEtYY83JDXz48BVWwuLy/IR
dxTuyE9jtni9iwdDkAa7CYFu2d3x3qRWxAKLeXqnuyLSpsUet5/6dNPkpDtZBFuW
wNxO7WdQLT5rxRAW0MF3ZLqDHI6JDLSofK8xI3+Nqxs+t9syiRpPfOrEQSOjqjsc
Ibf5QhBV40pbGT3lX7gxQ/GryRFq6kn92DmUeIDgt1HY/4y4wpyVvFlHOo/6i8CC
1MtLUn5ALeOT0B5IaZ5MdVXIKViBVki515zABr63cazkDUXbJRGKGhnIFT4RWAUc
m7/GWXBQB4nmFlwOizWEqE7ImlGs01VncV1Bfq09aCFrZsjTlyfgCgTWLO0w6Ka+
yJ0nPfwkf5XJOqHHvxwQ6Y9Xu/yHWUNAAED+S3n3DcQGk/WGqXZlRoxahPMqAuPk
LMusFbqLlokfLzJj5ZVtWGNUtRILn0fXhs//A7GPOTLVaIVNLN1NhU4xq7DRKGNm
gLJZVPKgsgxjfaHcCESkOIOQ6Fph/BKcTAiCLctUOK4c4CBc2Iccbpv+j9aFLBAe
+JlSEdQ+LlMfMacO/A+YQgiICQ9yZrHPqEJ2yh/rnvgwQyM4ns86RFHv+O9YjQ3a
3gJwCGATRun7yMgFWrKjFXRUHvc49C0+koPnYL/rVqz+SBigYEXZYEWhtcgLRSUa
UbQMnTlXmohtWN4ILC8Wvg7L8fxGUBXXp3Xw6kIce71p9j/E79PZLVo6kanV/JMk
/Whl3x1pr66QMqP5NCTJn+Izy1jTEZAeDGk4W2saSOHvbLytTcfBpQ3/+Y+mzWzb
2PsBNyxBKfMPtUetAYpOmjfWvgZG7XlmAAcYzsjUAUI9X7xsIji7yDy7K+bD68mk
2s2mzpOTYf6E4+ss83pT0sD3OJU1DLpqrE1pJpiJrOblz8TNy4PfStjtEDYAZakk
2MMaRQogQihIt8JSd+RNe69eo+KS7JICFKLK7B7Lr5LOy0V5p94eH1aOcwWLKSZZ
izmh7lQiJeQPw3Vl8J+yneWFMvKVMdd9DN9AUkV39np2xz9WsRXcDU2OwEByHOZR
2EpBLSc0ii9SXlvWjWDkHTPV2JBvq7TyOCjVtfH+fnckj8F2KdC1x9L2yH/JAozz
Oka5uHsjml25AKrVE7W5W9Qg7kvMTXQqgNvNKjLnjnZ+4mjGLQzjvuLXl3vmtLW/
zDq8MURcphvLjMwq9cVisTaesuDWZ0aPKcPzb7PnN8mZdS33ubr87uDyLvpQ9ON6
3MSJe/zkYDS3cZ5Wx3b7DXIGi5kLau6q6PrvNJy7PbYpky/dCLX3eowIuMxuDLQk
fmdAYOIWvdkzWQJmUj2QRxZlHj1WQ+ZIp8STETbxAyBqQEtL8Bd3ETQi/+X3h3wM
PlXJ73EWsvAdO/7ucoyVj+MnHWgt9GTnQy9g1qT0T7MJpw/caeninP55nZ4OEztP
1tMHo9tSQGIv0auyuRFApkjVxC5FY7f/kd/Pmi8bR5nL9+OhI/RUa5+8LXJ+TFfU
12qdPmU/BX+LzSz7QG18jZatrI6lsJDbszP3AHmq0m0X3sisYAz10t6OPMyIBh04
7IVAyTdjFcRiyusus0uxCB9ImsNRTPoSu0RuPcSUYkFT0D/umhyf/KjuaTsNpNfC
M8J0lWWxcNlzYttOZ7HOhL2h+TpPQCLe1su3LfRxYL7NUmM95JosCNA0LS3Bh5KV
sTzttSbzhy8pcrbmxAFQZjPGFWFr0ATwou0A/Ox13x+nJaLi10H+RnFIPVNpkTwg
J0QZ6022t5LZpKn7339aATBhS73Qh43sogCISakUg5a31az9V6eaD79tedX9HFrJ
`protect END_PROTECTED
