`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6ml26bhZ5YhOFwn0lB7IZ30ieGYrGQent0CqZnpzOT/eElJa+O836f1OKG09vcn
7/RZ42sAq+9+w/tGOc/NuHghReOvpu9z7HnwYcwvRWi9kM6AmkSiLP/Fn6rQSWS4
yvx9A7M8ydu2SmaVOr/islOjyHC2u5SlybhKGVwLratNQxlj2HVSgaSUJAVbEY0z
bkiQw45YxB071qZ+u0RzzMNGD2V06pDfDQnXu72lHIPlrKRrJBSb06cBWZKJvOBE
f9rLiQeQ8j7GMrMIy0v+QKwuhYqq+6mb08TxvvYpBU+hFvs8cK79xNEUIlngmg+V
uFLaazpbmtrYkFAm3pKsYtFX2hKdMmpY9JjNVvTZUESuAskpW3G/c8F8xBRFVCNm
nQxVL+tXcg/zey443hewoOUGJ+fYcvkHdT6VYZACVg9ldQCCqOqDahIGBvzcePsD
CUHcgfzkTNwg0cqcJy24FdR7/M04uN0s3dW5Q4UK+lknMx2onbb1e0uOtdNI7nRu
rvC0Et6l6+BOpDCrCJn09hqHONd7U4VHzr63/yGfh7A79SzI+oOhVTguczgcGjKu
r3P78FGM4Ir9pM0a8WvBpievAVljnlrtTCsPSNZrFMwiRTE5Es4nti3DAtRrXDxa
3sGvbqHa7Fuanc+u3xWcJjfOfzwM0DSmbMWiYsI831MRPFZZjk2D1ZYAXujgtnP3
yjZR/UErTCHrcrKl3ewjeMVWDUzueQMQJDaM5fOpGYJarZD8EalMTUf744yG5Kqy
bE3UOYJ9QLmGEdlpm4RHvA0HYexYlGHD6/jMb8RQR+FCsX4gg7PpCyAlpqHzovDw
SJRrzmlU024qmv2WDf5tu5Rqt70s8SZP+cHUhCXw0vvA6HmH2i+xh8lhAj+dtV8t
J1nOC4e4JSYLrxMiUlSEEF0RnUKOTn0v7fejRFs+Y9o51hKRALQ7rv8BxuVGXAfw
EcTtP6KRdYxf9/2pq6Ox8Wj7v7NxTlCbk6AKs5OFYwPKabraHuzdWkAVmGqMHU0R
1lR+MsT2nzN6A/qRlxwatHO3UyfcTTWUQBTA/TDq/r+6ZQWzch/n77cfEfkVX2/S
/x+TI3/u6ejGBY0dJ/MNiiF7/NqjT3OXmgrc66VWfmBZxJhowj+JnSOzoBlVEqKj
Edau+EwNF2oLHQAKGZcEQA4qHPVPHfeQ9LPgb4oHXlZASvnIzBEqlE5w0LMSxSUn
aPcCQA/llSIYopbb9HdQ8prhsGR2VnoqotUysRfJpt7VBBdOjo5k3Te3xU5J4EXw
vFHO86RyajsvUTTtUFdCNNL2KgURmPfAcezFrVlljMpmfa13MGm7iCdA6HyakXJ9
VFGWf6CMi2Jw14kG6uaAXwF/JJ0OfNaNMtArh9oEVOGiEqDZW7Qmjc+JmEcKKhwH
Gp3j/IVnX0pJT+Qe8T+66LAmWa6pj3SVJLS0cdasoyS1fMvHJCYxKPViMOOe68S/
ZNhI9UZLBHZGwrD62BGv/bfXKMnLm4t320Q/eo6zz8l701b/9OaAO1VuSAwBsAha
n3QZNiGxb1Qa3G/NkOI7rW3XTsf65yAe/NRObb9YVC2C6G5W6E+ej8wUKzIa30ye
zbd4mOKJ980Jr/w5ZfybPuPaH0alz7hXP1b/i8U3Q59kvWJsK1lRkmZ+/Z4CVs3p
SVbErI9yfw4ThX/snYGCACf8Ke3RqPWHyu++E1PC6AHMtoEhC4+cFXqm+yZAONmP
HqRH9XpTuZmJa8i0UWm6gvRZh60BjRZDwC1RZQpt9DKtqXJQKJtLWa5vSwzXev9n
0xZEidQ49dnV4ksX88AIwXUP1R9fuMhl+lfIdTZJF4i7A6rYXXbTs8O5g+PgBlWY
SLPvUN8/7NcAiaE55fifH9/UAenZINJFmaTsEnZRKb0tYd2owE5x1pATaFloLkhj
JPhVjgkSDsW2c0RFO2LHLZ+tZFvqJAAG3SFBESecXLBJTJ9o0E7iMTBA6czm1nPB
xb6yscnJ7dAKagz+Lc3WCijmXI4FVzWC5Hol2Rz2jOVXJoRfEV2CzVy4d12qJ+gx
ppRaQaWHo21f2Xr0oXEJrqZ068v3INHVRh5lyUYlxAbozUoQo4iejImyBJzvdg9H
nHJP5FH0Y651pZGTZZXZC+v4P8k0eNkBqJXQuNoIDUgPE+aBUUVVr/QRTgVqLIJ/
x7I/VxhckCNaqpfJ/MCifLe61WcdfrChpAALaMs0G9ffWXsrQsRMBEb+IV5oqQL7
WbfqjKj7w7vYhiGCj1gBMiLz24uFhzAqa+zHP+hLxd0qDsDbkTG0JKKyDAuFWezf
tVAxanIewGh/xsdIyo+54Mjqgs/+5GopvVb5vUCbRXzgoN/me6vsuMgepc2qCxlO
iZ4Ik6Fi7ITHGhy5ueuI3U/Yaxk8ARBYvtv+3RHUGrrgNm7D1vavy3zNBokK7Fv9
7oZTWccPD3A/lehpTKWnudo2YZEmbt/fMoKRXPRBY04Hy9VUJRI984zAEDQV9s3/
trX7njhRpL09yeuiI7wIyp1Shin1O5UPOj/JmnAxFMIEg+HWYLuHPNyQTEFSXvtZ
hMwJgC2IUS6/XfDAHiqoNONFfr0poLrOUH9yS1oikRe635L0diU+BZHKX+hQOZN3
wlgLkdhOjH+Nfrovsp/0h8f47ruzyOWODwWHHu+N3RLrQIjP9a9gaxNiCp5iqj88
nG/azmWF8lU+j+69CC8QCxlSsnxjBMgRJtsmVOr8uCOvHEtl8SsqApZ6ZMZmZ7OI
pzEGT4qEngeV3V0u5zDwbx+uMPesP80OJfLwx+9R5p6jpS5UvoPWq24nhsahH7N6
za5OoDYrxlL5LG9nPbgAyW9Vw+HJzSbTCbMNLGoMfBS6758SBY6E8YSnunuh0h12
fgOu+mrVujqP84NC+x3aQfhifjomyWMyONMsk4JYuaOypsPeO+ZAgkYO6q4SBZzA
XWsej9M07cL3jHlFAMiTNIkWHL/WcIITeZ58aV3bE0ypctgn9cydiX3XdwV3hYbi
n+QkqD+oilhZOADeWjjPNHZ9bHeG8owtyBjuSEO7gZKYFmZkZb1E8QHt+id0/+Pd
JKtzQ+N/v2CUwn+3IEW2AmCtfp4aXV6EnG1Gf7VKTvs436S3TDWFC6M3m00gPPlM
l6I1cT5tl8Fx1yCsHSvzcNvRYKn+58S/5O8Axs3wJw8T7Wr4jFuhe6ez3bSOQMBy
FIR1DZ1gmZKry3Ra1RXgugV73lIeTVBw5IBHQctoWPyFLdNFa79OQTJHmcDyL2S4
w5PdgoZH43b6pELwW4Tfthibwc+G4g/CqeKcm+k5PRNsjyMyuIO64rGmoCg4WJ0X
YbAt8ziNLim8jWfLRZmuWfwXJ9dpiyxnaLFfo6gbwrn554DE7fksUlhddxWwFMwB
Lj7rlJT3rArglvD1VcSvfPe2GK9G0PvHUZJ/4M7sPFAtUN4C/62Bag94UUNTts5g
uE7VKnIyq44WM1bccBew0up8vpY94Nm8B5orttWJ90W1kV2aORVjVS0SqC3mTXtp
darV8sTXXK+FgJn0XrhsTC/l1vPkFOvHdGjO4tEBWC1p2j29MwuDEKENf4NO3dWK
UPx9B9Yq4Ukyq1u4Axz9TgIIoKa/YUODcTM+1tL1jDhchAkqtUFO1H3N2FHmbmhW
/Ryf/LtcP4qxvIDPPX40l1PWmNKjHehwzmcqQE3uBG/KYCrjPCDxvDYu1BHi8kE7
AAdJfYrEeuPdEUYBUiOqPpRwL2y9jQrjegOuz6yP0oC/C30l2wM55pcqX70fl2b5
yxdVYzIlxyYcmS9G6z9xRGtEqnU5VieGkCJiz2NiJ2Uh91JwVjTDE/TJVS80ickM
wdeKiqjVhd86SwuVFJrFIue6GWSWHVvocPivoIB7fz9bhdKjnOyUEPhsP7ImrmXJ
S8GiuZjMXryy1VHqifxfOEtn7NOJwuh7A2FUZJe8BI900FfBDQ2/7ENRLdwNErs5
cmR54qE1BFrzIzt+QgkTim+f09bfnfNj3gN7aq0d4PnHqcb2sPy1VXAGkf3+1Q8K
dUn0lybXVOWEnK80s5lJrJi91DLXO/w14bIkNDcGAX+husT2a1r4W0GbRmG9bp+r
xq9HrXVUveGzL3OEwDOkugdKxd8JVSD0PR7r3UCuibyjNIXu1YlQBPDGMbhr2/nB
C4VM+VKr8NSXBFhH2wLwyu5Fw712+IM9EQVirbB6rMu5ML73cjoN1F/Ul1yJSGr6
Xzs9dbqYN5iOTy5YaknGIf3sbzaFgtf4dpwL+rzbfOWCZSa6iEFyqdjyR52hUuIL
2d+/qtHxc8uRU7pz0UobXxNjWjUCeTM0mIi9FoBhGB4=
`protect END_PROTECTED
