`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdoDra0YTPE/i1dJYXc7V8KzsQzrrBGoW/jfEm3rHoMLjNd//zCtJ/JJp2Gc9r1b
MO2hcaMT6Al+HRZNGHT9tUXh76U0vabZzZC5ZCj2PpxZ1+HxF3Ppu+YzuUpAJW2+
iOEE/RUsouErZP1d2/svfFpAzE6CDEzbLefM+Gffq4eED/TV1a4oiydU7EO4k5rv
khxzry0TedVFYj1E7DkMSDKckRdP9IbY06gWMeYt5sF5BDuAn86MnW+Dwe3APgke
kdxOZdnQ8ovLJdatyb0pykDX81T8T/FPPQUjEbG8kSJZL07AAqnKRZ84tBAw7gXn
hGkILN2GicSh11NF0ihr3aEW1CRUC+hgr//5QS8WBPIQDnlx+knrEA0k3SRWYbhW
eKiH1suW7wNGa3hnpW5uBTR/u+2RLIFY1iCbTN4D8V1IJSER33gdD6B4a4uCkQcR
fxf+gh8weTXWNEqx10kf45b2gf5lXbEYQUMSDxMpaWC13ku6q86f919gfce+vyLB
U37sIWxzPB669MYmwtMa32fXp2cWzjCAR0zW2TzVanNFBAbmOZpJAseUR6dOqM4F
lzkZ/pChCNx5BD+2mQIUHLHQyLwRcO6eMYyeF2vUjYDNIHYunYWj6L4Ue51FQgFn
SAuIOmvL5ar+h3AyX81uUzTxwM9PG+9qDmSiABlIxEUvzkgViDCw8SoVfBtGmv2E
2Buqxc7PuvJVP1MO+tJ8OW9lCFRJT6uR82KmC11GwbABRKq8/mTPrzdlZuC/of5m
eNw3gyXjCOWynj0pLXNPP4iTLLMIM90A4eIIab+3zvokJBKkXrj4FicacNljtIiC
NNmqCfyKjB/hi1THFvc2FYAWrnsVjym2MDgDOOfbwlKA9AZ4uIhsdq6ZZyZ87anq
+hy1bOGkneUY/EJR2SReM/AIOfxf+3SrnHfvZKChgf0IrAKiNrNsljFbGbb411d4
1vsnsnlKQ27S3oM/6MqEl8NAnCjIT2TmuYhAbEF59TCNXU2FAcGKg9HgLRgbMmk1
hN9tK2fBzqMKgw9QPo6Pg1yhn63oNvOW/HtXkiOV6Odjypco4bVzHTJXUJvY5TKB
bc8Q/Bu5Ugrfl3bYWyVL9nvzOnNMiibcXVH6eItXAq769phlbn1E66va0zCWYOw6
3+05DJcB8OZ6L5M0AKcCSx1if+wuMF7zONQYETJnfD3dKOu1mD4+r3hv8jwrJZsQ
XOm9grTcyaTlcM73ag5AJflxvYU7N5apeNniFXVnlMnuSKb9tTrR/oN18NoKXzo6
c7HXG4fwLSoFPIDrRlDoHJ7wqFVbWM6F3+UmFAqNe5jaaT+ovHK8jUKP85kNipsP
+eUoFS9zAeGowAhHPsld9MZC2UGzSdN6IIgQ/hOXdCaKLo3xOi+jnznEteohiIQG
4q7DM3yCCKKAf0ZnkbfqNjSfTWDmBPVuwFu3o5eq3h4v3gwHO6Zbstlsm8/TQBji
fP19FxDRflqwFHTZr9cHLf54slhnWDG1XJfZ6fbpQym2RIDMfgXY0/fkouWXYfjx
I5wkdnrdr0hxZzpFPE+xrrxEQHj7mo96f7P++CNp8+FC/euSM2MfUqmxu4NsWgQz
x3q2B8ivpvu8wul8LdPGJ/zOT5hFaCekzgrntZzGrQk0tFIU9OBbEEc23+MysVk2
T8sPycWht1Z/ZrBKqCCXHx8a9e0cfgaINF7XEuW6R+GrQl4TUyF5fqnDTsqQFJc1
ifPxvqG9mksnRTLKMQ0PJIezjJQ472h8D5gaf6wW61TY/yveddOuUaOBa7R30erQ
y/Xdunq4tHrGrBj9KImhfMdFUz/qR+bDTJpmD5lwtqKcU28fdw9sch0Uss2Rs6mP
/+mv8wSm38YZcaE+t4mqDAQQrPVabbQVZLjtWMwyvp/OnxC+wbr8H7F8s0yYt+kR
01BvOWJ50CoMjf9kUBjeQ5MNw48gr5tCdxYyl7FB156/I3sC+O7+IzFChmdvZ30K
xnYeF3JCFCPq6tvoaRf5uI+7Rg5imP3ZHKPlL4vZzqBKH4thr76P0KBLcm8l9qRt
phKyFSDqX1+xJFbx7XWosZGe6qiM6LM2i4/4dhdfFnFv97vVVp52Q4n22AxIa74/
VJu+1oGPH4X5nkai3aDwl4hzVc0IHZ3HqPQKV5evrpUNVsj5ebOmLZjUs8WSGrvn
`protect END_PROTECTED
