`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l4EkoU1KU0BBhSW2DxGeo7t/zsODaYWzktkCi7xNwBGccIiNpaiNnQU5mBpWnNoJ
qFFL27QXqUhvCB+sJ12HQoCWvJBDJkaQActsR1R6ahpHGkAqZIx2ofjWEGBqJDBB
wWjQGSL3t7fo5SlnrVQNdq6lZ+3dDBa3vXXXNo8VKrf6gmz7eTWdnB9mROxiib1v
LyC8aBxM3NY/K+tB50YoDcX3qhUS81w87xsSs+Foc5/vM+l5lVtcQkMMiVl41Chf
9brnHRj6XttUFLJglPh88azyoV/PO42dGllYXfAreyZpHRgb2MVQzVrkt8MhkKLW
el7IWRXkxMqStmFLBXMAl/MA1mX7tRdSylMuGb+UkCy+tqWpaVu0uF2nYy3hqvK2
3ruuIcNlX7Pz/x4J+jp3cV6zGq3PN5KP5CXvR+hTIrH2nfYM2HFBoa7WzPBF8+Ma
mt1xOZgkk5An0nrk04kbTccQCEXgZ23eVPstaVKsY/eN32UEZrbYu2TwO8+5PqLm
+lLSwBYf0XbCEsD6/YHidcghGMLGJ3YbwmXLd6MF9xZhcIeRitHvCYBdSdSKUpOc
IIpW0hbVmJKcYbPcvOs4hSIOB0BTC537b3LhS6A9VEuQbm8jgkrJhkeNbTo5fFvq
26o8Irb28CNQ8t39UxhAmp2SDxnYpnj2X3SF9Ejkx3p5AMndJl19mGYxXtD3PjEW
iXDPVj7MovcHUZtNWjjO5R4f0WTJajNzAOHpYuGIamjHPrXxhdUFAmmC5eVmnMPt
xLRE1eLuv3Rc97WINWKifm1Hq0jw1DE68PvOAFckooLPbhw0e4nOStQ/mEz3eMfy
lteUSwSXy4jzTE5b6W/uwhc1DKVyZvONtSuc9m0Z5DHGEwpPMrak+iAKePnvx54C
lr10maLnNqS+cBtGSyZ1uQ/PaOk4hpfbABb0Pvwb9FfNtznrcZF1fxd78FyiEmAi
bUAcvtCrG+EsmQzlCTwnx0AWUrRdMMrSCGwE6cnsmyEFxtXGNyuvFdfmHe/rOP+W
JNzaNX6tFB3Erd6CUZvVTJXs6SxB/2G4VDwPfVuQbzMn51h4g06yLwupoAU/kaym
ge75/SFiu2ET1TPY1v8mR8JMRTLOOWJXZj0+Y4SHX+DiHIDLLTLrlvH924c17GZC
HYsDbS5RckP3i5dXYmzR4Jtd28+5u3Rkqe3gSqld2cY=
`protect END_PROTECTED
