`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lX3I3VIB2U+1io7Vm7t59P/fkS5vt1odv3bkzwif+3fWuCO0GTzycB+5XeT6K1lt
BbJ/IvBOeSW8QZ/4c9O5Ba6L1owjBokiYB0RTIgN1jz2rjX775NEUGEEfPQkjLd2
Sof/4N+BX/cYY4Xr4OTb7c3Mq16hE8otaxsgR+ZqiMud6A+mt1uSs1ZRbf0+Krbi
a+gwulp7wZbDafOvdOx9W7OrmbWIBq0L9m6ztaBfF5DSo8/KIce01SQx90JbwS1b
Q0gHRaFVp80mffM+v1K5bJaZlTzkUQM3p0Yhgpq2R0FenFP9gbBZn38P6nFvdEPi
QGH7EHptuXd+0UAn2ZWGwSTClz+GnNaG431phdavS2fLem0sp6CgA6Irt4ZzjxEK
Jjc1ahZWGB1uyWHdXDBkE2NBzGM3JtnazIzTb03eyezgnXM0Sr57BYRECsLuSRR0
L+B15ABGUqHl8NxxviTY1dnpVpqXwPLUMVkYBanP2TK3ClrSfzM48BgZ+PmPX5Ky
zFRm6tKVlA3KgvxT26HKsTxBTkCDWc+zYbfxNZmnf6Yd+80lybb/Vvjl09bsfZgL
`protect END_PROTECTED
