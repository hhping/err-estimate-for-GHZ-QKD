`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h19l01Ns/VhAAc31Gx1ebxDNzXx+uBPl1o3PanlfELNmnNDpDrjCxBtTv1CXrK75
i6A54DOFn5FEFHBRdv67rOT7oSHPGGZtNgNYfk5LQyVVZb+YyZ+UATIMSJASuGdM
HKT4rWg5RiDLckOjOT13gUHslB0dibKM6xlm3JrMvk2rrnri97FXuhajQR7HQ6G6
9g5q9QlJ3lsfuWPGzK0+3137i4uvz8uyoEUmmp7jZQk=
`protect END_PROTECTED
