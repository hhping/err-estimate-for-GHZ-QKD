`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PT9EpF+RP9eykLMFY+wyDW4iUQt8kQuy6U/ztvWA4Gu4F50629ExpHzfONEdegTF
uCyfZOFTlWn9v3CDp3bQ+pPaGvot7Z6ODzW9LXhskxmYwaV1j6Jokhw45PY992RY
/ahrbKA5p1i7xT+TsO2FUbiEGGpjZfPYMnWufl8H+9bDmLT0AO17QuFma9H96IVD
XoTSFn94s/ZhzAD4EdDQh4BNI9ZSMgZwfdwSLyiOpIE21TaMWAI4CSNOc8uuyOLs
ojMG/IvhBzczSdkIum7RlX1dx6GsnQwBQ8AWQ3P3QnexFK+IymdkHZYEcxOKJorW
wFCLMWIZ+EuJGpMDLkkQE+fjX8z/i620sg+OMe7TJG2YUnuyKYx7Ame2GQNdmyjO
wPNR2D6Zmb4aadxOrVXpXItFetqXt6KQ6r/p6KOqFpeQu6DQOblxwGbOKEGzZiYv
RaWDBzwud45hP05hx6csTDv1z8q5DJwceJgFiAJwLq48I5Scfi8H8KK/YpWHCnA8
9Zb2GSA6t/9rWOEL8hKXd2JTzThZQlsNiRfOfz1e8zpT9sdOk2gisB8+MmCYrS5u
shDVml3SN1VjIO80GS5n4HNuSP5RlUFgDNFQ2UtpqDklGJESAHM8JVK2akE/fyWl
yYwq43/ObLWlOm1zdbEc25wmGAoyl9XKb/ByUbDJU+i5YEikdKi3+UBNbkEVhmCz
qBIqRGO+qt9ahItFNxEi3sF0OaEtNMWFJ0HHCwn6GCWsHcNNXjDUGSNF+XdBg4Qp
YdPtokNC1lM+7SEyCm8H2du/Fsuvh/BJA91Go8Pjyjiz09kjeVPx0GrSIGE5s20y
PEVQahXk29x24cYS8fsDz0cuPedLCrUAVsukYbvfUSjKmRxEjzF1oIrPiqfS6ShL
3tlauZiePBb8JSlMgaMvzQ==
`protect END_PROTECTED
