`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5a5V+9Vh6I2HEpP8oywPtkUvvi9XOeg8Qx09u5ss1CM/RCxI9cQK9OV8q8nwUpi
fwLu5oziDRY7EsbkGHFWrV1OZ2YlfzU/xB0a8dF1GWPIW4FN1ClScVEJB8FPqWo6
PsnM75+kzgwWlZS0Tt0nBlHv4fN6FBXcmzJRE4lRrGdCLMcMQpoYlc9yUL6ieiVq
zoaVFA1A0LuJERc8nnqbhPz8wSaZ+wdQeLf7H6sJy1LBFfoZ2MEkA+L7cVIheQ3l
yMrUp+qI3eRB1KtlpAHPRNJDpsv4rGIUc0WZ4Lgz+QZW3+ivkW6Pi9nrPbgP2c1A
b+bc+g2ToTFx3+l5bIadK/m4YDG9FJ2ij7OFeKScoLV3LbiY2cfdX6kPhdwVitrm
BAUibhMWjCJnYG/McedsWSXiLTBmMRKfvOdX4tvJZtBt278C5iRggq/DrFEb96rh
vujVKm+CPEibQbHpVN9opb9Ij+CoobNdIOUXYOxaNyImOQAScBpzfN6/RU5tLEZq
YtVhNJx+zsLjiqHK3fuSbO32ybgY18pigfXIRCH4FyeXj1tg6cjWNx2HXjVCyhgJ
z0S44X7hd8hb88OLH5k2HriDcxqhjW5Ih6mJfiO6yk8ClbHPHYpsL67cPviW8z+j
pCnBv1bAWJ3ysphHReZqtvvvXafiaw93c41C1tuHkeQbMtf6EbkY0+OKtr0Kg93c
c+dqNcZs+/jhRJouyoL4IS1R9LBCporqRjRkQhGIyxAGug6uWLHF8AcnZCnghL4/
idnDFzM5fi+w+3w/IvDp5AhPW9/6Qvuo7qzr9aavldhiU4I9HebzAnLxHyhh33/H
cZ0g6TNDc//yEKeVfrabTlr4T8Nbb5m1RrS1JZ+tYO01/90jdOMwKGflDnOWRUiR
8vF2tNuyslKYiw9V9DzXjFUROzps6jtvYyFr3MdY0UCha2+/OasFBjG0UN9K++cG
owx4Rg8d9zzI6hEsC5wZOQVezvisZBa+GXlrug7mjezr0kRvh1wEWlp8G1Yvy7Kf
QZBlt0iPRALPgVigkrXOwJb+H0lwJsZS6Jvwc7usn6FOu9u3cppSk09MMHqaDJ/T
HPCjuq5GkSmbvKwHdBThPFWi6Fm/Qkl3Rh0Mj4JbR/QjzlsPcnaS93yqTuQoSYTD
onLCgr94oks5T0/MnVEKsU7Ps0dbC0HwaYs7BSJYQxwAoAfUK1MEtKYYEcYF4c60
5pdMKepxWnOPat9I2SuozlwK2Yg1XGVGquSPRjSZaZhtXB4EOiMN0EwQr4zx/czD
Zk09qYY/guuG6iubK+9mf5D7qz+ov4ScGTj4oCfmMTAxhXARjkJPxCnqP9e+HjZR
PVFw805QLB/g6YTlOkmBWFN/DqPxKp3FMacTy1M3+IyV/vKhyoa1vrwV/84VSHCf
t+efFz3WvUcHn3eZ/2s0egRLMUjF0WwEj9rev/G1Rgzmif63LjpyPgqkhrjoyu2/
+TzUXRsslo+CXyoa535Vwl6bbGfDivdLvQ7V6Sjz218b1cgn9dQiPBDq/L4Rjikd
4aLJD7WAsZB6EcYOsLAJzvrIdQOEaGePb6QJ4icyXYIt0j39RcTec1KdVzAmneEd
FqwHi03Pe1/Yaz194wUAQqpI5lqRulHLKfiKKvhulU7jkDGl0YZdhxAIyhgbH6aW
kGB/RbsRJFDYSSKPPZrCVEokbwfs70OXA1V1pOZSFUxg/nij+Q6SuAHFC1/tfmhe
JiEvNf4v0TGEiboSoSFoxjlNNy3hcx32ttm6NIbtcowic28kZldqHef9qxQsj39r
cIemuSN0idFGO3nUJDjnwtYC26bBlYFSMMLw0Skdbu9lJJcyWOT53GG60YfOSdty
Iu5+gIwb5w8Tt6lTUUdizeSG9Rvp9a5AVTo8+m6vrbFL2ipiNjBF5oqe3agcqi6t
zmWPDxZ4fdedkJTFieVGG2WM6PMOSctKUPXLD8vHlyCOz2GDZ7b4htHRZtYM61Ty
Nyo/iRCWLMQv2IHI0Sq386KHYMZFfyevA101axRqBwr8DcvmhsBs/P++t03vUr2w
GRpI9WMyW5b6/08qeZYx1IZka1MYMAy9dd6AgJpeWg00tKJFEeuDp1ngfnN4k3z6
J/rx5vvc/HmNFoiHR/ttYGu9UZDC22uZMiXV7AcBptR2vKoFMLBA32g0ZSky5npV
q1os8Yk6yJvmhLUdR9e30GolUI0axv01Xff/WLK2GDyVboa+WGDD6aBeUAaE2vp3
bmOBpi9WLeqh9WmQG7AJG+qd7QXJ4XDoSj4I/9gJNciXgnmfHy4TgN1li3/yFmZt
XwZ++SFsecYG1b3IQXthVjF687ovcBvVhaB8hi3Dw9KtwVjbItkh3OKUKNSfrPrE
MvOy/rUxL6YsPJAV1Sl6doaRHAtxpxAO8nAHXDyPdnAq8kx8kTlLGi92VKd3971T
qERf+zhVsaFN669S70E/n4/GZ1byeHQTx7TtopmbWNAhGrnDupqMUgWkHhRiygYo
dSegAZ+1cbe3/jym7dZXU4XNGCwXwZ7uutjh4fNQcSZobbP6MtGDmhOC2BTq/vCD
pIV2x0wHLy+vQGo2zW63JM2ej1t4c6hl+2kyzgEKe9LxejWyQm/nca1yemNFGoSy
qmNRJrFc76w/GdgkjXE8JGA6/gd0WnqWY8yCk96iMKA+6oA+HDeh8tzI6u5c9Spn
EnMP5/wFOb+QbFYPrwmqyLc17YkECcjZ+5bj+VpUq35/PtoDmuwSzTP2GBFUyNJB
6lJNXEjb70Vb2KMwA4Q73PxtwTCMDD0cfkaAy5VjzloxbygUd9IlztoYNvN8A+Fz
i3QvmUsKSLp51nbp8rklUlyiuef8FaeHuRi1gOYeHpvTIFqMzknSsjsUlX7mh5ZT
bttU4cgexuStZVQeGGLfe0i1fc3WEnmwbahWMUH0TsfqM16YF/qxfnwLp5JXZwZQ
UJ/5iSq8ZkAihjlQ1BOebwEOhu+Msm6602jyta/iKOoTufDegy2bhG50culZibeS
V8HOVoab9gmktPY7TOlt2Bbjq+cY8xsjA2GGxxhoi+Mn8QKuO1XDT63QfEkhoFua
3xBsDOAeSr4Je7Ke1RjnH1ubJ8ltdZtwOldCIio55mrYIHQ6dQk24YExUnwcnfiU
My7KIKsQSAcp/8Gw60WGUArpi21D70IveEauM7+J2yo7d2Ljtc0DV48DWRMpCQjo
VFCaTeobYfUy09KNGyBFpWJaE3kqcsc57Bp2yXyVcO8=
`protect END_PROTECTED
