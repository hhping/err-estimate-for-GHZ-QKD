`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zWT79vRsTTyKLAaMzS06JG11/qUDN0GGoWGZs4lOdUiFOgq0ybnOc7ykUA+NNyvT
6AzJZFxqU+u4ZTocuAT29RBWAN/Za6FjD67+8n8w7P23FfuMsxEaChGa8NvaI8YJ
m5j6qoWRhlikD6tctSMDjKa4rdjXxnGS9gkpUm7Lx/eObxLkW7+gF7svl/FIaM5t
e7qBPnRp8xGJwd0lrB+DMqDKFUMLgjZIxElwIm4hX7ts29MpWw2wHAhghdWBoZkQ
HF3HKmbhkO1oCbwiMwnd1wsvj87h4MilEylQlChnsFWY4QwtI1hI7uh6y7o/uz2T
sarjbwyllYVwHSiaGxY5DRQ6u78eKidZEYN7Dd0sqHblBfkMUaBs3PiKL0MVUs4G
yKE3etaI2XFknexQve7OOI/4fjUNcOb8FHVxdKlv1FAtvIfOEf+yBn7ki4uI7RS+
8BI3730+ELMw3m9dw5tDW8g3Dq9DVgbWpziigXbIUT41QFrbCgF/e40AyQjep3Id
k02xW3yTnEOLsxQZfdU2HR0EIqGZiS9hIgKp87/NmhJfOrlXjek+Fl6Jp5KTI3jx
LEavpfE6p4S/VxzWvBmalzhYrpTkreDfDZpGYTbVJAzys6sDTDuUnNU69HiuW9K/
+y7WC045890sBBeQmmZaAfwaxpbzxTEWgKpnpu1X/Va/YfIMxBxX25ABZrqeKYVt
9n1OfVrfJAl5EzWKT7td4+Cv+iv4Uh7K5Fgjk316EAmxNXwdqlFZKVoDw+lJf4WV
sMqNwQ/HoAdQohrzmMzajX+LlEMJymIp20QWWYv1rqu+q1jbW5hOPAQjZ3XGrm5X
t1WNhsgkYS1aMmNfSgeiZgxsM9E2wPn+EZRXNla95mtR44QFc6oibYrRlSXZ2POX
0dFWlbYdJSqb12y8yy5fbxRpOFK+aVOMhpI7U8nzkG3KhJRIZN1xGw2/tPFyLIu4
BqgDbIDNf/npR7sve3i3dSlNRqfJIwSZHz6RUEECD6QBfLYoZ0+kECJYP4CEvxZr
2J31E7kTpN5vt5DmfcOrgb8xX3dsVFPNT2X5TtKt9es0+fPetC+vr2vRXRZrtOa+
cyJGiC86gyZ98dN3j6JtHWYH/DhOEVx9VvAhFv/IyP+QCQQYPWxhtWUAq4yGWGP3
N1xqKkSlxEPe1xOdZaUpamDj0S0EESNlQyonu7zMemf6RgNZt/SIrz61sZKCVU7F
YR4VQunPmrcqR36YH9wDDxwLC9My8sL5SjFKHMNuTshaugm994QT1Rhv4PrqMvkz
iqIa7kIokXrACehD0Mjfu3WBTQopkjbBqCZae/zOb+BpiUKMKZ87qbghsqHoeIU1
G7LWBGYprRKOEJ8vJUDKgpnZ05KeREyYJjjH6UCHiPIg2TStXlG/K2u8OKcs+Lau
uR0MGP1eLEADZYHiB7ZlN0v+Nquuk11lAaIEM/A4R1T7DadtmxNYXvg2/Ul+ZIyB
vJofHQ30KPBf86ubiwtoFdZx8ub2xZp9G9tKHjpzh8Jp6C8C4eViJKyazIRF6ip4
FaFKHFdjM0domodBhzxRNlBKGhm/4iL9m24KrGJhpebMECGDx/Gkou6uICOviuM6
7EtcCWVn8tLHCRvBIChFa0mZJfG768tKXN17T90kBl581f3RUcRCqS++++2o8fJb
ZRpEsIHCeD0DYneaWd/zBU/LaPbqe8vNIXCpvKvVljW3C8a6HhZ25mrv/FopY9nh
784F8dDW3tKnBtgE0/xu4s67hIYNvzEGfAom5q3fB9yOEbz5OwrDdSfzqDzaFYSj
d+6LX4XyOFtUwCsu3vDCUa/QK8xUxRy0vz8CrQt5nd1R7ERJmbRlJ1O6VT8R/Qmj
J1hhn2kDaB+IOngK2+4oZHi4NOFY3I95T2/aXJCbr6WaVNrjeMM/25asWXpI0BLm
6X8IqrxZbyYfDuKRJpCD1J3pI0J322/OJGO67P9xAHypoCbiy8J9OSOND9LL2koC
WghoGXYUP1ISf/opjAOBjTVCqXOwoOUWBrvUoebjKT3hklR8mpWOmjkztT01nEGM
VY7fPuD9sRfudY5QnwAExsOr5qPh0xeV9Pyv2uU7sbuBn5ZqwLthynACPU2BX+bb
WjrJkMUNciQFGVjkaci69IOg2u5O2UEvj50wHZG0KyAN2IL5qgk6Ct3lAqdeBobP
BKo5MzUdy89bwkaKJDqyC47F6vy2MUdOWOHFn9NDYbfVJz+SjR9rm/kLS1Z02BBC
7ODiYnb4QXhW8UrESbGpPaTZAt9GUyLUjFKuCV5/u7J8J5fRvg3dKSghKWeoDZIL
9rDtrzabV2NONPSIa/FJTF93efVT/gGlPuSznfq+pFW2tmqNchDBxr7mukCa2ztJ
SOq9yYHWEfnkgC8uy3mYUnVLG5J4ZyLH24puWKAgzMil8/5anMy1JWsY9/qbf/sE
wtRf+C7kSSfvoNiczMTbjcMDIlYKnYpYKOlTOM7cQvp/UIqYN0OR9tpnN1f0Imkv
bTBFT5UhMaxTmbu3B3dk2qBvpTx42gFlrtQvSJFAbo7u9yKqYO4zp3ZUo3zm1K24
uPtRnG1maj8oE+xw/Th4exAxBbHgrh2OdIYW5zpr1JouL3MgctNm5ZHYxuWvkqda
shzvBG9WNEE+FyM8wI9jJxG5VG0HOmLJCvJJY37V2PZqMa1FGsz4xkHpUrUx2bNI
1kEHF+QzfuWmro/gP6/4PmVgxYGBg9SsAQVSwcREjcXYoilue1u4GISG6bHJp2wq
yfY/eiYBiLRoVED+AbN1+CLr5HGjH3nKDpT07qpXLymDDKkmX16W8nywOXiN/Pld
5WZyuZafjQ1E9VKFUrZjVMhc7eZBUspyaiGD/PWsWGneUm0uKyOWEdxAeKYl8EMT
HfSp3YERBmT1xlY2fRFmPDD3X2N8Epw7MzWIyBHxulpf7CUrOokN0IgeNRn/B4As
VxDpAUpodV/Q3UJcCK9e0L011Z+yM9z4qD03s3nK8lTs51IDVKHPSDynaFO9cBzf
a70xx7dh6o0d4gvMXKUgI4wMsfvAthrtRWthCgtY3M6RV13dom7FksYoQlle/EJI
51zUuaMV23bXsxsqdjVv7b6bcYYEb2aCffOjMpSeq+s9ooDgIq5Msg+qg7e5Iyuu
zwjGn9eRfw4XT8YQlq3wTa/0aTm935RzooaXH7/PZx3Y5Q5ra4DmErB7xTHkKdlX
SB0WSAJSrDWXcg6INq6VEEu32UH+4M9wz2LRGc7TQCu/PK3/bN5LFARweLK4NFwD
mdRYnGrLkpwEWZJYyQ1stjrKqlw3U7AJp3gObbiQ/vySNaP7xc3UiqlHzeNaYoY8
db8iszeXdosE1lmsV33Gz/ZNL5doFkeuzm5wk3/RFLYBoZS3uacMIMABEjbyoh05
BdAQBwBVgTLKrm5ttcVLkfQ+Uv1ZmEb9D6IFADIub8iPB4isX/TwTDbVkB86CAhu
bB+VkXv6IBPAgIZlQ725ommV4KQZ1pcNuhtxGY66fk8+unZNUhzTPUfaG8Ixlmim
ulUFG2KWVxyzcFqTOlTKoTeYBiBon1RzW/RlBT2PREsyg/pqZw9gjObLFQhF3+e8
9YrqfwKdvXFZM1LPHp/9pAwztbkePQlIFYPJ3eSJCp1oHmDJTlXZyGQK5lMd4sTr
gDfqpH5QO4VXZ+viFp7hz66rn18p3TlI8wKvVgSCMbtSkK0OVjzA13bOI9OVVFhj
kcStC4T7zqn7xmAcAXf2NGr7OEIqwWaxoNtj9BqXrwR8pCYKZ6+TmilK3wHEoA7L
NapD/eQkJc00mTLIWpzS9l0Xcs7geIf2ZVl97yRH6Gm8wLmFd2LhyFDlJulXwQJb
+wQKddreax/ImRurZHCNWjsuP89lwnX7Sndn4jVtoKrUO2OjQ4DI0GRSsNxbiJdn
V0DbmCXBEORhdzryP6uYqx3CqQXJdZGqQkDbBV4++ENy6WESZv2JvualommQ6pcq
J00f6HEUSkTipYEjizOi1IYr1Qk+qjGIquzuUsiAtzD+/N5Icm0HM07whQerJeWE
hTawxEeJEmzLfMy3RMGCV9PTHE4SK8OrJ2Shba024/n4EjgfyYzpDlErdNHbsP2h
A/d/uUEvrQhU4VMYTfwp6Iumu8+QtOWKgmQNgJ78TB0DZpFbory1Evz+ZUI6jCa9
FlNB0k36o5QVPwMDr0w8cACNRvYjfGYC1zA0T6W1PFyN2Z0i3HJjk0SZ64HOjx2w
AuM7U9uKgzwp26NoL6zFn2l4Zv5SO1psDtEn+GCCdZSGer2nCcqlf4wL5TW/LFwE
7FkQXMibR2UipGYGzA6LCTfMWR9LdnqY/AvpwxeoRbR0KK8EJDvPBuXqFrZfX3N/
yZDZoT3kb/ewLhLlgA67egyMKo67Q0lMh5UosuWTgo3wMxrnkPRKXwXZgAcKxiKF
6ivrzW2rkSqz4fPomdpeGXuEBlhx5QmIZB6p1Chhu3arzfT3Z1mLzwnxz7s+EMLR
Ae6G1v9l3/7K4r/RYaCIBvfQV10wSlLAa7J/kQRlyQJ1kfEma0MS/T6jumu5AcKJ
c5cjK8czX0ZWGmD5Ol7Auf3KFo0XGr6sVQTyvGDeT/WZzQvJ4eaqvugI3HKidDAo
zqTT0NYcz1q0HcbUfWVPHH/VgZJ3ZISRbPgSJAa2nU1tl7Xhz+8Xhk/8BrEe0BxX
hHVqtIHxZiS5nGjqBps/ZenkG73XHxLgGqGKyO/0/CMWjpU2HzSOVX5LrEJvk28n
+yur7OPucqiD8+B4j4OgpMvBWEXigCXBCQWxpePzqJJgsUe1K78w5Ln3qPa3HrEg
kRWi6D0o4EtwBbFeL5o5eC1e1slT5ygbw9wCUGM86qGeVav0LhngzC6QLiUVe2gW
A4Uib3I1atpEuhmNIkogEhhProdGzAKan0OseW5yDJyFSopwJHZAGsVsBtV580vU
r2w5Iaj2jE3F8dK/TXT9pfuL7PXeQJPUdoDIr7YeTEQuZSpt9rJYH8+xn+fRfPhX
Z9SCYRGUj+lsVF+mTR2gKYkvHRqplC4Vrrcd3YE+dF7JzzggZW952ZFNbdJzY8Qy
7YGqmX5CTs43HMMjPJu3Vs0yHu68aBFz2W+gZpdCA4JuCeL4Kyn+0GsSyd+LCMMH
Hhc2yzGDlKLRfehfuTl5LSFGklCfT7+2s0MqVVWZ2Yeu/BIWzhsTjhr9eL/0pk3K
1o8D+q63zOWJ7MVbvoPdeqlF/OMFqAh1cD7vqm/TnG3x7GtY0rDdajHlDyX2CAk5
NGnLyjkAQrGVjL5dmY2gajfqy9s6Sd5BAHqsW38Ncr6+N4YsbZ39RO9EYwZTri8G
/R/BY1y/YeNkyv9ZZbhVSCchO5EKGzoONvuH3Vp3qohy+zx94olcp8eNBjFC4wml
69e3oc0t+JeErCams42x3O/8rf15oqcxikes4fDpY53ONYLjkLJsi8aoQE2RjWYo
feERJHyX/pAExE4OPF6vZfrG7fQbMkXaJHQp4PjXjDMuX7TUYQ+UT8rH1C2IHxSV
sN89uXzkM5VehhbieD6iiG93lAJxbcpfZTyQh2N36KXWAcvMalnGzAOvFyBXbvbS
sueBxTs83y8QRhcwY98kW7hem6kjvzQjJv09eB3e9qljX7hVl9SXRBLRsB4ZObmw
xCFPXivKLSK/HwH1VutTY1JWKnM+GrjCSbZjWYhG9oBMjTbGiVZhK6JAuxCuLC7V
Zx8Fpjd68CUKRWw4+dEPsYaAttctgvJRWqQgUq1VU9rhbexnT7+/3ie4cJphkUSQ
6vw1evIXWMPgZwZgGpqP/BKOnb1DTdZh61EZG8bLWgMafoqp4G+DK/+fQXIAFKa3
nF/gSbxbpgshI+xKYpUHYoORC1nqVSlpU987b6zX7CZJpYDliVNffu28GyzrO+BH
hBfTyZ/7zaytg83m5Anu2TPG0Zekyohdt7d/bpZeYtzK2XufsPKCz74ew1LnQqTw
RxuynYA14sV0dX1bdVFMTxl8RB3CvH20jeIj3KEOtZyOpRj6tDJsB3ipvaTT2ke2
iLG0SNS1pfpZ3B3X5jKxEy2g6M0CAcarCRXdu1dZtvPAAdoUXTvfsiks1x9ytEb1
vataG9akzooMAx3whI0LayJhH5zMkp22py4bhrCfuaEbGBCwvWgqIJPXj1yV8WWB
3e8JQ9Dlto9tY61mex92wIbBQqsOtm7s7I6yqfR0SMkG6bLkK3JtF3mgs7dDMdVn
iJSjcNaYW9Oam7xNclYLDPVnwYe0CDc48WzCc0ZszS5+9HhL9IVHx/hUiH8tgeOb
puRWn12oLu/FBkIPVMdCgGE/qA7ORIoh0bPFzd0tew6lMq/q6OZucDiikUNxxyEs
/lCRnxENdv+gwfmZLxy17Hz2s73r6AV/sRBI0t08WH/L07a7BJlBKEy05vMCkcYt
EDDkXMqE4x1G+jTZZwgs/URYrQJi6w6QWRFR2aIoMuJykCPjZR+HVwLZdiBxStEz
D30qyE0w57sQiCMD88fDvt+6FEXW7quAY0dPtvIDtsa9EVAl/VXWfUmE2GBLe5KT
s9qrv/1F+4zylILDv1A14sCmm4DgzWySy5jvcte64bZVZeCzkgxfyOAeQzcX03Af
jrv47CaWZOMO5xnCJzemhXJAz5fF13fVvI5c1V8U5VpDNn7py0Ngh1K/6oFuns5d
IzHLz2YAKDGm1pxfYTcWldmtJ83yqjoRAb7sXnkVhD+quEeZDhPjGIVNb13hRJqV
JLv4eqjSIZVRRElpIOQsBMrVnMKzylE/0PJyu5w/Rbs4UdI4Wo5sRsNPDeFKdjlT
AZUsOcxfeih6AOXXcB++n3GTEh8FUca73RgGmt4io3mX+9b2RvEL0rcBv8T0SBTd
wVe9DN2RAhRL7Sq6hFYYMOSQwmoC9/DGbb0NlVtci/PgIsjd+Yf6kBUWwKIons2l
ReAfehrrE6dRpeuTuC+OqCd4xiobU5zLyMelcy9EIFZBnBwzMNOJESSXhC8iT/gf
TlXdXrq7xeAfT054s14FEDJj+gUtWp1w/j7cop85AFV02NxG9t68ewpQbthGSfH3
2m1bwpGYLKZJfNqKKCKkGGq4WOQqO0pUqtFXu6BuUC7yHZKlRVSR05TNHwT9SA+2
4srCxmPdbzKLIlNX1aLWCgEn0GI5S1VXTMofIKmixAhChZG7PsXKbKyIeeKUosE8
MTwfMPHPV2hWrSWMSGZSuQey8eyrUQU4+RC7Yjv1TdgRP3O7GXkEOGFLGfNOJCKb
qHErZkZzt95LsnUu0sjujbU58Uv0lk+UQm26HGCG5pRqktKdeFPtdkKwjflK1AUU
gC//o2T1no8u5mPFJoqtocTKHFpBw9tDAJC0+eWSHPIF4zsuyEUDzXV4z28tk+V6
6dVZMsnpFvCkfZr0woKvBHfjAeTHm5XLmZJJWKaFnufrP8hfTZTytqNSA+Z4vnjm
l2g81+mbx5NBqUHRCXSReUjPEwDh5h7f5Eig9Jzxc6bIc3Uu23pJ7KEWhb+ztN/u
D/kKdir/RWUCc7uIO2U6uZDYkEiUj3rIIn6tiMK1lkMR3cuXFki+WhEYdLRwADJa
sT6QC1k5U4FewLev5rOdz8YiUnpbPvVj6+vbIYPyBXmQKI6z74ykb1Q9X6jU6CWe
U11v0skcVPzOsJBj/DSICZnuhoKiRu0Ac36u5LvHXKoyU9CwrhmGeeJqwTRYuDGO
ZntbxAcyQiqh9db2f0cN0Hrj0fF3S5NehrkMnvjqdq/AvLM0N57w+zjYXeKWitng
Lr93xodmO4YeaPYV8+vFu+PPAeouQcxrWrFY9r/QGD5UQQfotKy9zBtkz+WdHvGe
UAQcrDT7G6SATGArWI5td+BX6i2YZMQ8byje9ufDc/0gcpLh3RDa9YMWX/2AcWMs
Iylw2wkbosJEAt5tGIqLhh3FqoKu+IY+ltSfTZIevj7cddCcIyyoZ4qdgx7uOO+f
3kNMElOe6+R7ycO4ynVmGWfds4xck/TRlkdO7HfEjSxfq1zpXgqC++N02WpUeH6V
689NzLxA+ZaYQcFvIZHuWKCFCDxzOGj39h3dqNzgNg4lXwoADzmOr7qhGSbES3iz
JXYBTUDtR9eLHybg6SOug38fKGvFdQSdBxh+FUgz+mx6R4GLcG1VPyuR34Bo1xls
ZAxoDl66/FebV0XZIWjC185kw62yyVdTI9rfycFKlmnXsMaMQqs83IH3dau7Zw4e
mxUzvCzRNuW1uNqw9kJuhoQwP5uqp24EN2h/adET3GDDOc3fJi2pLm7LP5alwmX1
DZe1/rRGrMSslj1W2/5m/467RQyp0wiNtyNJYA7t35SbLeZkwTCFGC9gauUk0HRy
Joc7h7/gZNdXEPEAxoBe1QiV/pTiLLNhv2wmwuupe077TCSiKHragHQ9bYkHJ4CR
xm1/kMkADWyutjlCQqs8g5mf4FWCTIiR0R1okyx/fUY4sajl3BrLZuCzRie0/aSu
Kb9uQHotY4b8z1EGEygYatoAcey6CDaRE0bryucguVZaOWgdcWWnfLO4Ng0i0RfL
0I60EN9EeB3AKzHNNdsLkuWZL3TOfORPgpMQcEaR3zd4doE1qlUGw2D4RNNJqm55
1Jdk+485M2I0wP/bPKaIFHmLX+iWzJgz1ORPJtlVHnqlS+A1p2qK2Ok5Ud07Od28
AvX3ySZxpPOm5ZgmN+4yH8i9zZsg6t1+gR4fypgkevtjCrvN/fUI9Fc8HNCS8nLY
gSS9XbuFs550Pg5UxDuN4rKw3iaFUrd4XxliEA9BpiOiA4qimQq8XzSVorfUNxrB
T/D/3oDaNkYxjgyg/hGir0BTQZ9KVvdxtUwz0EnQJOHYlBHqiBXlv1CzuXH9uIxO
SDOfFYSltw46h2UfPciqYRrephHqnctw5jHitRMkLTqzFjZbBBrUQdZU2FFX6cSQ
DYYx7sWP03xP1AGzdHoIrTclDXdI9SfdAaJ3Lf+4Ba3kIM7KVfiOAtNPoOu4FK16
JZkdf9NkGKRzer2vOMGGenGT6NwzW9w6QmCyzrPw0nlHw6iArgPGKmxok6c3tAGa
us/wamfX2HXHqBHCpn9+X7RZLipAwC+qZID7OIhtPQwNW5DXfVnSN8l1/tM134hy
3FzNiVqW6eyRVoQ85/vhoHRN6reVhLP5W2bV/hs58zqwXT9/XGynTvSOUqAHCRt5
8F7kFhTYE77RkdqdjyUj1swL9YP1IEIgk449xJc1g/8ITgYDeE4zDXdduKRXADcQ
R3Tc6mXcrhuCMXR6lfCFfOXXnuJCESZF/Su8G5De54t124PHkDwUR8s4msBaFCH8
Y4p5SiNHQIv+6zEXdbu7ForEQGbN3y0ADBjbq1hzrpqeElSd200XsZYwCMyDgktm
sgS7hecH6rd0TOJa4Jd+ERi3SkTVKvgZyWIToqfFctxjs1lMm96mrENrN+Fg1Y6q
IbpbgBTpEdiY2yBWalKQ0S9Y0377o7pgk5u+7x4pHXR7KMEdAV/CdVky4wUEqQEW
5Fe99/uNfPkfKPOzfIM22bbSYjWgFQXYOZ9qibNApqg9H/fXDbHnZNJxTC2JGMeE
Qv7UzwecUjpYZG1/93oC+Sq8XuOJTIDbGdvPN1QASHpBDVgYPCE/L5wSTL5ZvgBF
MtXpW91kH5vgRgs7C3zQui1XxisahbzrrJi3Dd8LIw9KHvY3uCr+B6TSN0tIPSMo
+TVxP8ZtdhBE2TiBMd7TGjLxA6szvkBGyq5rWTej7ww3O+ogPDS8oSCMDDQy3IMM
HfxWC05OMAitRS44SzXpFsXt2sx8DrYA/uqo9WE6OnLDG7JZw2VSCXcLgAdof0kk
3xPSQRFBt2qwXo0mHo+56DsLd6D/aGTCIZ/ciBbeoYb/kDcsCicM23dSNzPqMAb7
C0o+jR9EiL5cU22Hfs9iIQrlUXL9n2AtNb9pAmCwV4wtdFjt3jfDBqCJc9aLB8i4
T5CNfHhMqCOv/tpEw4x1syx9/iKnENC2iIufiOXT4ZCssEm0jOmTqajP0GDWHkc3
TTtm4WjQnw1/RCzV6+P2vNU7m/NkeKqjKgsD9+y1TA5D0QJ4ER3XIJDMTbWZ78r1
8nUmLIA7FtJX5qj2/cLgQF0Z4em6kXfdPmsL9tVnyc+BBBA0fiso1d8rRwnL5KzS
ZGWYXg75yVlq4miuVHAfYrLgQoEdi3j5H+tTQBasUy6cA7MDgPWbgwhAu5gSx3UZ
gZX1WqVEYfUjmExJzydJxoaxMuFlhjP+NukyFGsmYwEsd1yxleE1KiWcCAa65eDA
OJ1Ys/R/Fe/+HWTis3SMhF1yAXuqaFxGROE321wiuxZFVe/dxGCYb0keAinMriib
Lpb73e6A2FqgtN/Ys4oaIwY8G+EeG3WHN62XMiqofMD2wN6+O3THkz3lhHspZGr2
lKyQ8+gDYw3aF7PasIR+mfwXvefa9uvrizUgCJuakQcBEWyvxXZV/hABtU/ItUQ3
JrlHEUpiW6axw79FBcU2KiXCbq+LIxwN368Z3AaWDct0sdWC/amQMhNLtFT8oy59
oTIiwtE0D5iONcjyRw0geu9wOG/cu0vpqWxhD0Yx/cJl8/F1oJE6zh1AkbiDJH1V
l8KZ1nqn+czTV8C2PzNcfhNyOx/7et/JHRQ9c7SXT4+5QTm9jjmsUeGeE+tpVprR
SajPMzV979LTYFN0ZVtyHHsVuzP8ySBTEwDyn93o5jIBRQkq8/p/d1hrjMWkGZau
8wuNHtMo1oNFHJldG3zpkQ+P2Z6CRobZbuviwJvQQ5PY9d/7ee30hjgflAAQF6qB
Kj1yiZKUhxzCz/Wc/9RJzA9Z6DkmN4vxEA789ogLC+MGbI8CFT0/2wpZdcpWEC5/
T6kYbjocyCEnmqmCSe62z5BQGhxV20q5mi2w39H9+5YKOLGaatkkEqYRPUHTF+Hx
rR+YwcFE353X5L4e4d0IqO693cznjABtFjm6n5w3O//dGukGa8UO5KUdx7pgKgij
urTcluCpIsCc4f0O76YQaI0y+qNybONoiZNDGQkT2/q0rAZIPfDXogzR+34PybxQ
gif0ejwj/aJtBWs9PkbLytCKYlbC/qeqvE48ql7tX0iSfeGui9FLQBpPd/lXtQVr
rfxtKucFxDOJPUyaL+BIU/lDqsDVqrpJkwRK0mfTqXy0v+Er0K0N/gxis2tisbwd
jptF8th6BgjOQQ8lfIRuOV4eWznh2cZQl2KDp0kXAwUhe4YnJMHbeCba8aL/AYIZ
jBeydrwaWoo2p9JldLviRlOU/pSw/fv3DEmckqPXYdBGHJo556aUtcrPmFQfcsnZ
iw0k3AvoppfGM60umubk/fsxld7Jdwp12EpFITlkUIwxx+xN9OGtOoIWF8CkqgoX
Ofhg7MnKCtIC04euLLR+gALAs/Z1lr8pB1Pjn/FHaujO2EmO4u5vF47DP3b/Rhad
Rf4li7j/Fd5JMYQEJ9oxGeO8DLcP65YQEKFGT5gteDVmNIuJk/nb6WeEv8yLP1va
vHNduVdxj0dyrEX+rJzZGsswoAA8QoBWpOUN8psevTatqj/aYetc+WA/fQAttg//
VtLI0zjCyj8Vz8jD+k7brPFu2kjplBJQDf/cuDrs5pzCUt1AsFwFb2pr3HZV25hf
1SL5meEbWtqQBz1sVj3wW6yu1mdfcH4Aw++ubIv6lSRMYh4iZQx7QapgY38QWhWD
w2kO8YKb1J8lFjro/ruW2Wr8wSiRPOeuy71I+fal5wyUG9jtFd82x+W5X+dq//jm
a+Obubu03Sn3XrzuHyTbYEFaCjmJf5ljP5Bxy4rMSE4sbTyo6fZr4R4bPP5BoEIT
ZNdMrMz802Seoi0sv+wb+EPOvc48w3MAakqLhfwQcBlh4ztFLamtj0fL5Sfyayd3
vQMKi6N4YGLghDEev1nJt/ugxznZxflJq/Ki8/XkR4h8hhaRIHdLalCrT40Ttf/s
Cz517c3Id9l6pGWnI0XhNikfsJonCkhYABAuH5fERY6As3l5JB8uVUFpkL+0JGhK
Ik6hF94p9v3hxmnR9XxlvCLnuOCSUTmjDg4oeT1cXOCcgX/ZlMq7pIqvJseKgysL
3hfd43KsUU18X+P4k6pY1cPbIti1ncahEOuSFstYdcHGMeMBVdTSlEHJi9mChhiV
IkAP6jL9WpAeM19w2yCZiVJRpl0jqMOq98uyeB7bRiMtLoctoElCMdxTEJKahoNO
675TDr4iljWN3sa4OwYysN4wlb/ihEAku9d2Yx+LJ4LKHrgSxQFuWEfqVexmG7G2
oeDHDpuo7usMOm86Ljymst48qADT+6S0N1y2Xl4xj8GaF8pZlJXD5nDpe7IDk1kJ
9t7ftyNcqv8arlH4Khn40jz0LDDuyI63QloO1I67cLHHl6sLdLN8/7zlIAGxklE6
6u8N6kS7CTsE/60e13hv42+AQQ2Z/560yFD2/FSeMacmA8Xb0QRUVUD0OF8kMSyU
2ZPOIVy3e68zBJcu17WE73Ee4/YD2p3tHGfREaPeU0pz3Vt54LMU4Mzoj0VsEodf
4uNSu0aLFxwgtcgDIw922Eq/Q9nlNmdnHL1ccotmMG7OX38gAcTsM04UPMujFSsu
uay2YwXdp6CxOxhRBgVM5cTK5WoZCSAUY/f2oCxA4eS/E9QaHY+AXb+TgjLePddH
DELhTuqbQVrz6fpn/MK9ECkdvjO3JsuygvDR0ffNU9F7FqorFQGW1vBY8xmzZtwF
+zS9Ao/uKXgDtUlPNv42ixULCjbM4uy6fzK2Mk8OCbHqaDHwiVCIDoCzOk/BEBrd
lSyeFcR5pTfFjNboTKiVMSqe8cc/6qaoTxubbWGx35Hma1WzRdJamVT5vvrJP8JZ
4ic5/3FTuK2pkwv0/GZUp8tZcxqxMU7V/JBcGOrNyBrwfyXeEvOjhx8JPZsfWXa+
ng8JUzrSQlvqox9EgROucYO8jBe40jqTqwKOb4N9S4Fed1U2fE+tkcmv2OhmqAM8
vxmrTP8hAg1EUbw1vwTzWMafqhhoOs1bjcf8SDLPPcSg+bbKi1I6a7seqxGErR5i
9yDHAg7ixFQ0b2XHm5lPlZgFIM4/ZW/jB5/3Kh6o9YK4ng8+mzeHkqAMkTGuoMxu
n75m2GdjQT2zRIHrFDvnisaiZCIs1NKy8JpSVFI2T/NhCw4FjFw/EyWnz+GmjlGc
+yLbEFg8RFkFRN/ynEFAbYroWOOPn5CbrXyMvFnADJkOzJ8cd/2iShvWFHx4870X
zZ1UeiTmd76wPxjM6CZ/9M61/uScHKmBYg9p2L3HosT/dPyqY1/en/uxTJw3cxU6
JAJ56wk42MHRisXSyY28uTfnY4h9/DPMc5zcgN4tTv1pQlsastUFuH/eZ4Fr0LtK
GIo5PEWE447ITsD+LsUt9QdcMLIn5kPpXXjlU23+10ZWHH3ojv9t1Ohm6484YoTy
eZagbyYSJy9Jl6u2eTpsuE3U3/y6MTUVRo452Tyrbm1Lxb80YmophpAYJgGmlMBa
9K/tJzL64JqETyT/NoQMcaSN2AyzDSVQ3HzM6pQBlYbWVUWbC6+XvuMGImfBAKFu
BKdz/bcEncmZUlxt44xFtBVGExTluDu96BbK0a3kvy63UC+YqJBWDW8eV+QY6OpC
HXYFZMXQ2+Dka2lYu92/niUEMta+44uXLurn2gx5PTKCwQ50ElTlwFoLC+aoYb78
82CF2st2OHnkjXLX/ceKJl0O2gtHGrC4sCBKmCK9C26U9LBwJapm7chSDkYdm9I9
yUNxfpAfpYDhZCxGkXuODJ/hEVWwtSvVOFyB2XmHEfKRTLM7jp2qgNY+LdQbtUpv
X+Tav98DSfE8Air/EQf1Qs8t1idNV3zoO7lIpeq7l7YDDgssPrsb9L9SgFBZtIlJ
DHXYlMPXjP84PM7jP57mRgcvjJUNrYdnKETmDAUokhrnvgraaZ/v0JCOAGxIsiMj
VT0u5U3KA+tlqp/0Bvl7jK6RXGp6TzQT1ev6exaw4Cmtcym2PkzK8iy8f6dv95H+
P/aQ1/SHZliBWOy7c0eFF8PGABl/qyrzNaWbJ6k1Mf8e5rxLzYPiLLq3TVGv7+8D
j0pTHf42pGO3h40wEQftMhriRlMdt4M10SQ+y6bdsqq8psEABGeew3+qeHz4iDTB
zfmMEy2rxqkbutDUIlueiyQScCiCBfYc6nIUHy9NSTrefynFW6N1sJBlNU6J0Xb8
7gV6K0MxgT+IoN7o1AvWALHChpdfXdLXAyBXJ1be8vKc8YyP+0ztT8GifcSHSZf3
peFQwh5GClt8TR5ZOiPUk5cOtbHjtHIDuUULjRHixk7B+8Vlb4fAHySAnH8fyWfu
XkFRiXmdHnypI+dDtZ1zlv6wLXjWxGvulUbKvUL18a1VRtt7wZAvvitL4TpLKcqO
b3zCxnYvmBVet1YSqHTeto0OTfB9pqfEV89NogIu+X2797I7M3yef0VOMYanI7Gn
xsLNiHTqz58tUlv4fKGIl/NsIKqYpCAoxlOjqISybXAi4xbmSaqw+yEcnaGb4Q1N
B6+mzwmeRYEoSfEO/ZMhX8apo/OWffCdh+EM7rAv79Dk291Yh1WiVsSs/cVSIzP1
tRXEB67meOOq+xgOhjDQCVwRrCOcVrdUQ2JSFX9oBAS+PY5ZINsWay7J3xNevtii
u77304DMHpmjvg9z/gWc0xbelrHMMUec/SUgI6mZTqjrXVeJ0aQlEBUwWs0CBb89
Q99pWLK+F58rsqtO9stKmCOrIphaF67f5IfTunJZQEALtwdGUZWt0nJFLmTOc015
CBoPlgQk5FQuwpRahYcnO11vIGjxcOLxly6R1XPyy3AZTorCWgRDDexi9O6J2eBB
Ww+8APpxrh8c/mxWjFzLG4Kap6zSgGldc9La+rZb3NVTQSUfjH4fDhtV3tSQWsi6
Y9niNBEfua7awc98gQ/lBmtnI9EFI7RkyJav5BkProbqSpH13QdfPSfgRXHRfSKG
vUuLQUCsc1xNYxCFhpTFAs33q/Tl5N8hSE1YiKriVWW+pUR5L4EGXYtjhWxLR2r0
+mNfyNp5N4IRmbIQhDhRfrQMrwjs0MKJey3C6aQfqnKmHeu3aRCrvhA4GoYKh/cz
Fr04An1Qc8zOvjLuLkVQQL8awd/OJ/sg5FIJIjnb5+H8ZS64ljqPxXFdwcE1H2Y4
UF4WXhtrqgTB7z8j0fneDx0eRxzkuzWiTvk1scUqgnAUb2lYw8m9RUgzhzxXxPI+
lDIK8tZc4jd+MTYU+GfKjrZ356StBaNmDlkM0YGdc5aWJohlVAKPq9ZpDJV/aMES
J0dFMcv0pt/bHtmYb5H5ealrQQyBBp7ZSnYpb9hTnqtMfBB9mcQd+wHGIVw43FG0
XVBijO7N0SxQSZtIXy4lV/LuXV5ZlmIFJwNDdUg77dCG89gZGkiVh86vfiEOfjkW
juYEKF/fNYawex7XMyhS4VwC7V1Qld4jCzWUQw6HNKM24yEA2E5P2R2igdOvIrIf
oCGvIIL7/19TiH0jsPk8kE6sfsN049xCmDqZGoKYkwcbaG6m9gKTBCSgznQj6qD3
uCRP0Mre7xDeW4KfCkYBgzqsESyFTCZuK3iVjiXKgV7QmMLRf+yqQpafHAV0ovBU
bcH58nSyRX73rNyu4ANmuQjtYuq69Dg/2uq6MWB7LbxsdAB9/YHMs1TqSDkrbg3v
Cx+V4VVosOQ1tPWuAlulhQlHHFkYkrPw2G5ULHUJYirFoD2AZ1i4sBhVx4XQEyO+
DlUQBrL/+iziatDvfUVvRvWrfygVSo5IU/38/Viv0F9ypUPeWGFKcAgojLI18pz+
9T0zRjoxl0GzZp+LitekOU39Wim3Jigyz63TPIfsuNyg8OPCbIg/SFbwjnht/SrT
peaawCM6EYXGPEArfl6PHHi4GDTezZ2/BcEvpslnZNc3r43T6see6yTUgsDbg0oR
hU+ekUCV7cekz7PWJ7hZVwmC7Q9LYu0mjvz3A75kxq35WciNAT9l661rzhnbV38F
Eymhf2x+itwGygdP0RCbeqriYg30QAEsd4O8rh3cUjCvAuagkMss5by5+XX4y4FR
wBt7FBGLTv3kT0x+LnCQL1+dU8fS9Mb3chXxSoNNtgFSGWFPaGq1iwT/mwzghRa4
bLFvsg75icdR1SRpVPNWxUQFKIYrjjgM/8fI7ufGcbiIUMWVYvEYxGf01L7Fr0pZ
8RFR6iQJidWAxFKMtBZ9wQPmLyy2NyJMtxkoursW3gElcjCeSCMbo77BK5svHPnO
jLEceC2ODBMdNJqrxQgRFkry1sukLWc2TnGytzdJscfdL6f+yoYwd+7LC5JjkKbW
x4egheBWpUsNJ7IXtosmxeGxSWNOJoIuUFzRAqwPXH9K+a8W/DcCNiTW/DOzDaAH
TFnx0Lqj1tGVahM/cUQPiOylcvy7ubZoEB2TFKNvkXtunfZZesUqEomIR7M4HbYH
cUyNyaAK+kbr14+WBFWFa5CvhsG64zWHC0foig9CjBpnQIlV26/7PYVtD3VfeB5V
uqUQRv+muTkcN+qgtfDRnQNpcUTknOd6+M4FNo0SFySq93Vx0FCFGHJ6zdJfg9dd
Nt0EwRYGbof8BOHoashCVR1ssXsErEh2IZOi8nRyvFlRT9zkhc4HyEfIzt8fzNR6
5n6rtNqFKW8WZlzBgN4yIyoaAwPnig6JQjNaVTpHfWovqQjJLUIhxNJ8SfYtB14j
jAOGUPUpbC2+jjQgMyZKLEa8yIdsF60b8ef0HGfs8UebcEYI822C427NwvFm2NSB
5kXiXgowjkjqheoCtN7tcK4Tcl9sMfUAin7C5NMaduF6nj91Nq04zwlPWUnxYtlH
O9ZlUSCH+6SEpsavDqWnHYSkm/yXlujI//fjDOuIcGyHLZTz1mcLf/V+GYgvfmmf
ynQ9nJjjjByOsUp/VMxc5jiLAa5CQ6kvDGXyGBLewDhz+x16zGwYgSEpvlhy3HWA
KuaEZUCCJ670W5kkp12d8B22lIgDMFR8E4ybg77+IPlOve3hRUPlDAo8c47AZszK
tfLH+ItFLzhhHnlCqFVA0TFHrNrQ2H/qzQDYoANiFNJ1ZRiSgt/rTK8RrpFJr45j
x0bLJt7z+1qbSASObopzIfOLpedT+QUWiICmEU3mwRltDc8jnlQJCzPfsMQdNrX4
ml6nrvfQe7QaEU7b7BUI0TY9GY09beWaeH5XXsJkLok/1OMRxerQnUrhAmGUFHWe
aRqk6PBRt/GLMSW6dtU/Q0kNluY0+MyYkvmaKjcGCeRq365LO9DtdWfojNG+h+Iz
3W/7PtkOfDHosdrmkk+UuLeEEVIsL7GKJ1hbl+qXQSGs0RsrhSCVgaRo6/nQV9GO
w9SrE5EQ4KCuPLweMeAFZAKq7sLUFzSvE2D0Cblo9KxMjP5eM7mBPc1w1RIokCP/
SS8CUR7rJgNA9+lEpfczgukvVH1HDMbdLTORqwhXpIGDbLWVywZkxJsGa9DbBziw
7+hWM69lRd8rmuPgJMR+bjnSK/AuK6wbCWJvKZDBJQL0ONGrvhGOspaA3aOt2uEw
eR5OenoOaCbsWFbZws4i67O1W46cEP527IG630Y14F5idZXeWPuunjlCVNhTUJUe
LgoNkf0XNvoWhGfT9qCX3tbzdM4yG2wqYVz4oVxwfcHe4ePvgoawxsnn8PCKoKF6
EFd/xm2yNCxcO2aCES2HWokggOYJC6gLffg3ZUnLd10Qg7uZcyGA7q+tqoLxuUbw
EdML6EXYnc/GYP/AWDjCoPkCFQj14xBmYGXlT3dSc/VwPIBi6s3cUU/jh5DGn8oc
jT8ETXCYdjNbsVGthWpAkIWg5XB4kT5ohd4uXDsAFy8OyhHcYXxAcgabH7mWNskM
IpA2pedMp9Z0PhPZAQTzlI10wQQHRY2d7QTXUfG9v7570RKJC8aSvOc93hTW/Cp/
p6S2JiZopBaDf+EpKISDDV19E4Fn8KHL9fwZoF6TPnOSP3y9cWITFYYuYffupAeY
a07AL4e4uNfp20s8kO2XWbBYOGoYNVvnEUIfiZE7Y2O/0519IZmHppIC14KTUnT/
eILoe+ePZS65ClDz+51UbhRGTZ97EVOTS1TaR2To5YtXDg1C4Enh/JGLx22WZbi5
Kb4gnaMbVQmUZStEEIFZ21mbfRZk1AfHLoRyoGiRMvv52xImLjZFzOU4xwkl6ADz
Ppgr+zZgZx+OeOwjpJFjozScfXRe58Ay2Xl+n/Iw6YUw+GWK80RPdIDheCHOoYp2
VSezXwmHtpBRGDWWCqAJ0dZxfyx0u98NRhAdtcoscNJN+lNOXYGQlTQqmFy+Ktwr
bawsUelr0ECiPff6OhGhXlaXLT3Wm/PsRd5JDiRJbn+iavQQxTCxRSmxdfjgzct+
5vRIaECeSoT094+n9ik/08LtRFbkmm9Q2nDDU6S4q7ZG6B3R8zhQcAzg2KbmxXFi
NArS8qFahbqsmSXdpWUe5pCiQR4fqNI/DeMAZ4jQ01zhDMMr1DdMOCHHUY/jIPBN
1RC5sX7tBYFpi5S12SlCekZsN59UhFlEXxGB3Lpyb9uC0Pcmvf6wWlmgcFvolYvb
tGHAO3zoHTi5X99Dx2DrY8X9sWRJaa+SI7VnKs6CxAsnhdh+h7ztx/LqgymRfP0f
I7cfvQM7OPLkqQuL8udCv2n+pJnF2IFq+JdH6ScdMHpvKMshUIOjhnHtaUOOkVEr
+gjGlO2jF6xVrJ6PrguZOeJoYmqH7Hua4FYZwIdGeq1mMUAGnWyy/8lY2wywLXB4
FDBCRmUQ7GrAb8DQpUV9VSmFoxq6/jU7xu25lgQWUymr+cHOVlvXFkKQIPHNE6k6
3OxxIoYBYbFydWZ3+3Zvspl1/xEv90GXqFBQajY5/Tr2R0pxYOUDjT3x1bmnK5wy
zNO62Rc5ZFCCaA9JY2WVeSHhToxtiRVOBdPX1/Ux3K4xSTaaKVEPLCd5kFiqsp5W
aT77fLotvb6RsVZCh5AAYON6+xnPbJCaYbYOu3a3WV6gE5z3i+B3lnwJtQWiZAsH
HFfmpMnczwufYMYUE91JaGzcAsE6MnvOFzKVOLbiO9eGo/S8z6D/I1eJaOv3zVH2
mH8A3xu5/TftgQhYKDIZkMcspy21J1RUNXbB44p9g33V4zYWN+RlejLzBQqnlRNZ
kdfSJJZ876dhWGIx8XHl92X1N28vOseFXN8Jbz58bH66mb6xDsXmf+tai6zDKOsT
uNe2Hy96zoyaHjmuzN0DiAbO2FxHDl1I5eGwcKs+ptHdVuuhR0PvzrJFa4p6cl0O
68M61HBJdg/XHCWVVj8DgenchYMt6IaUPCV1JBq2gjDEkFMxcb7G7cPa7rj3/lC4
+CrVKVjVfMJWpk6n/+AeLNiFjUOt0fO/qV/TpQN0RODc60zlJJ2NhjYiFXW6bYbz
rnSj5kkK4X0p4kvdVbNMoJuJ+yqdyuEdU5QU+TMJn77iFzhLzggGV0zDW87dyZd0
uoS3C71eD3aBeZuAOgcPkYjybojDaYzOnk6zKxO200R3iV0IlmTM8UiSx9fjr5Rn
U6NQg8cyhCflI5PJTX5X35dC0AVgHZF76vtJDSZrlGni0IEcJigFAymlJtoKZIjp
tUaBS0Uxe1vUd8hI5eSh4Ih9CpaX/9aP8HWX5rQ1NB4ehWlmEG6ZU/F56tTULrWt
xKBzapaNQZaKp8bTmgTt2VZg5izu4jlP7jHm/o8vmTvxfQHiOZZV3MM2wf3J7Sxd
d//Ba1vAMiwwA/CIxszWp7GJDB3s6Ah2Itn0CCfpVlk568mjbcu2ONO7x01h5pnc
Nxpt00S5QNM28B6gYl8fHd3JYvjETrcY6OgKiJcNpfMzyPiRFB0wYJdinfe3tZr0
cRuIdhN0GwhlC7n6MboOcTSO+3LhJkOfsfqr1hrXwR7UvgnjBT3nUFRW5AQ4Tohq
8QNG98rCTCLfZkc1gX/kJvcDRHugERCxrK5dPk9gGMVv1/f5uQEcEcLTJg2Ffdfm
qIXN44qzIFcFH1McHkbKaifpy5yRhZDK2CY0eFAsz25Fi5ebvfERVUXgMZvFkcSt
65Vj4mxY4Wocu+EKLwMXQJk7RJAn+9iHVy06VopwLwkgofVZB2GyAh14wp7ZKmI3
IaWgdcSVDlLwN5Xix4UlD1sxbBFSb6oSJ8FVdUkPZ9anjoMmWqO3RMHevEMiLflW
tCP2NU3yy/qHQDgj6kjxgmcR6uTuGajbmues2BwXjjgyMh4Sz2F+z2syOXUGjV7q
xf7CN0y0Nw9+wSdzjCkPWwq6vZw1k1Rm+gvvOqG2VO46lEQ4z6saRa/feJO6HVrB
PH/90BOEdL9oR9JFJLSLfy1bD3Po+i3fAamStK4wwkLJWYKleDyJaEYYlHWr2RE8
LlKliYv3zbcKIQ8008dUVKGi06T+v6IIFTDNz8y8US7lILm44LN6+kPWZWyf8Lri
loejUtM4ymN9LzjypmHOkFKGQ9qlkuoGzXhVrM0ZLIZJxMv7esTWGtvM0RtYV3JO
bIOTurEqAPkSAewl1Sl0A7wz6zgKfVbcppZseelmeheG8whuGCUylXV0/BRMXqfG
4D4aAisASZd50wMcEEbbzztuJL72oQRi8X+0mreRQ0Ou079uI4sPTNUrnkPMeXt8
npfGNwQX9mAFlrKHMcDOteZLZG3acVL7fAoeknL2KqitPTblqsb0lHVCINxryI9w
5RsWTSq+4zFb8CSapxHYYbx2k65FsqWI5Yda4iqD/X7lf/jBYX1tFVbpfnKAwxQF
4pzn6QUMvb1yxrwGkHDVJzjdm0w+l9Jax4Ol0H0H78uDI/1sHGzrTQ/h0qageDt2
EkSO7Y+fAjaPydJcPa+Gf5Xc4jXhnBkOB7EXWGYwaH+BiyVuDAGM5cI65mj/fSlG
ckD3SBrAuv+ZAriAAZK25tPSkscoQEQUVxpzwtjenovYbD9JPzZF2HY/D2LtNH72
vghj6fXFBIGWgZWieHRKRSqEQnbKU2ZOz+mubCzmakN2kqp893c3Y82KRrXldraj
eJpLoxxm0tZnImjVOwwe1+h/LJMsY9Hqscr4+7QGaiuB16NHO4wwgcDoBbU7GJhp
XFCgceb0Il/b/6xdtMbLxet3qGkODAAa2LxuNV+H3t1CyDFY8/apCyMOyPDlNEa6
R0STPRntlIL/+O3HRZWWzNZMoF/jNLWMX3+R6Rd4NnKYGdbk2yuervVDLzE8PtIo
nX/My47sEhZdqlVH+oAdr8WXfltj0hDe0h9zrqDc7SNcX3fX04tNtURNw4kFWoao
zTEx0tK/DC1hD8zjKkHDoUDzMuf/CPXmc6CwG+wH8klOj52ff79UBn18juwoutP+
aLmaUiVhFukYgnUyuSabLGHv99FvBR+Hpiae9ceT7kgl1p6ZZOoiXw1ZFt9yjL4U
jtZYMlbSKJ1IQE+LmWrgjEzHD7l1X0eLHIAVMQ63GTr9g7m+Jk81+QcBKN6aESA9
UwE3iUmnKGNU2P21xIPMCxnOtRfuaGizYZPIJX7+3FJo6CXhW/Hy6P+CQBcCHHfj
xqJ3V7SGG/0pEu9Sc2lE98Znct85+eNjXlmsfZEE7PKxDd5P9hYRNC1WJuoT4kXS
6ef8/dtkjxcvMNfiv5XLtEq9f33Obmuit6I+xTttV24QXz9pErlEww0VzonYLvw2
xZB/udNThQYPaNsIAEtUrnjfmuSZLklcl9H1RQmTFBzGo9a6PWd/C+UbYZ/3jZYc
sY9e2CgGL0YNcYLi0CWCoBVItcd+uQe2gem3aNxC4SLponLRvofKPXjt1DJfMD/c
aJHA39xjHKQWSTqPrtCqCzevhADfOmWq72IQxfgaAGIjTzdWj/STjpX2CuGvY3bi
ysXFZ2MlJbS9hKx6ZcrRcuYhqMMDWOvJ8nw5b1lxmgezIc40fWcJ407O9EW3VPHh
b0RcA/HeSicgOEG2rk73ZmU2Xui3uNj4jKokhLQYqW+lbXMdYhIGRk6uhzhDZPd6
/o83UuxDp1VdExWbgT51VQ5GtSSPpf/Pm38tevDPy251rRWPVWo194+KjjsTiGev
fOD55VrxpTn71i7QzCvoXkbIw4cjWu5p1CQn4Rej8B8h3uNphPqHv2icyCXXC+BN
mTTPaWNUU64p2STzfnKmuOkepDebzlVKrR7jF90J15Ld3HejqxeyDN0lg34DHcD1
r6AtNG3l2YSD4yNghuL/oqjzHKllWeCQRssZb6Jkc4mMITG536oamiexIT7hEnCj
RnfG8IF99If/SzY5hCsFPuluQiCEokQimi++dmoKVeR8epKwDytfts0+ZWtUzMdt
fIUOlBu33GS48v2LL+02v3+UFA2eJcdZ2mzPg4j3cGiEW/9JZerxZcB6WwkemzvF
tHK1z2Tvxli9hKIgawLU8TEtFhyDqOtuVVuIot6mWjQrFQyBgNYwjH+MJV6Fero5
YXFm4X2qAR0mPqkR5cee36bN/KELOGQv5h3VPedQ8O4BSniHIjNAyr00brlT0EhH
KMhZM3HUIzq9Bxm88VoefkjbmuY9mEzuvt0qYlzOX76mkPR/zbQZUETN3xQ+WZtx
sGlZPB2tZ/MZP57rvTlxquo8ncsRzsPJW0yQa//ZquvJDHvC9hiLeG9aPYBvM0y3
gj1a+DzS+Y9oVPau+Job98defmL9aE6e4asUGh1x3Yc/k8wTOS7IAlO2OcD2+xoM
oX71UfKCb7bEuOlE9/V4qh/nmaSa5FuKzoYQzdmJLfTOW6BVnWBpQ54MdhOALDe9
rdaMYylJGSE2oNR6Nv0kQ8ejmX3vcQ1O+fBe8nC/D9XiQ0BhsDf3CUUwMmQKf8kj
bB6sgbMGGHTbdAxZmrh+uPlHdiKzeY/uYdispw8RfiSZ6XYcrAz45VmzafWS3jN2
eOTn5hTmT/j+4WOnxZhBGeqQLI+7RIKfAFNWVswx47MwTDc6D43FYHuWFkGLGD7s
jTlNtSlc5HGXYLK0AFaCVpMOJGa2YAR9CJc82Sf19Pai42JxijXpWKEraOCjkim9
N81Wk7NsrLv0Zi+LTKaazB363BOFR4phqqG+ZHHpItwmSg+MH4wgfS5z3jwQSXhv
MfPCJmxAyEHT1gPCM4YJESG16UdkH37wc9LMkGyVzy6XdFF3MI/F+PGIwn94RUCV
vKVm3w+IYwWDvcAYcMx3O9EmpaEQBFmRE1Rtyy+uxfqs5aHPms11MR0126v7A8r4
K3UxNNuhVx/q5T00D6o2NdYu63AaPUZ37REFNa0Gf5ps8xRYgOWgEiu7spDJGYta
klaIIzK+ZEmuZIgshBUB6W3P/EWQcE0gF8lgXnzOPDhFu2k/YdePrb96rSiqUxtb
9WGf2jeGAP9NU0A8g3d4nBVYAG6O9MsFpC4MBLB7WdL1Ka97dWYt3rHbl96N5opa
JxMI0KMiv2lmGRw0zIeHswVRPeuiXinmSpNCI13hpMxf5BGJFfLvwewp0VL1e4wj
bYsVQC1Z/V4SN7LzdCLW1xICWuB9T5NdkLsRyK58xUb09vXe7PdOyPflYV3ZNLNy
H9SUvVHVLG0azlJ3t/nkHyoLuyVUsNoZgMymb1XvkWWbmGd7ykxPZgAuOdqRq+QC
5+18RHD5bjMLn3ytUKf5gW8RkSp6A4sdMTyXGZvs1oEJuCYXKeH92wutqM+6dK+A
8D9T/1BWkkFylwPUlfMhh+clzN6qmbk9/+TpsfnBmHW5576c2UbWbjWacAqjgLTs
SNmKTN6eJRBjum5QnZdOqKELaPWIa7xy1O3UqY/7G9SRewQwMHUPwHQ7hCi66ups
hfPoByOdMXiYVXjH8KbdnxBC/Yf9hvY6o18flk+Kk8dpdY5ZWvedQmB7XvwpbtLu
F+WRN/E76Sr/M1wTZRerW2Mag7fT2UmFBPlzGT/82Tgl5TgwQyWI0Rrvor1JpCZp
atqANW8/iNIIsgKbhyFc4kS8r3+dAUDRByYE76osLbj7oyixtgzqgS4NMSUZa1gX
4c+osy5tzUuElLCnEeXSKks6ZzsIZObvZlw073IyfTsZ/ORflZKPrnGXuhtdka43
UfReBSkFRWsynREh3h3yacr+ltzRD1Cv4LWsJRE20R6qEcnuOXInfqKlPkScK9e4
tSNU4RR5i5j8anf9eLKaLhkXZInXSD8KDmnxJnzS7PiresskGMzRG1zo7vpe+rdF
FMfDE5QGA0rvjlkIkBmvezBPwGLG5gbo98DUvVV5b5wKBCu4Ud5sLm9/hPQMBqwk
888kCTznlLQ1zvvRP6E0kl3O81FGnoUxwK2V1ijR29Gnwy+2BlU7aMJMicRks7HK
FYx4N3nVhCYLjCkQqEnKT+eqnC1oZ8jMKmASRUIB38g/iw17bnfGl4F8rLAR7MoH
umb0BIpxpYAxZB9SAtMAgf+0APpinwbRZu9oueqmoISVw/FRWDM3yEP7MWD7vkGf
vYQaVv6AWaVjRLEAVoNNVA+JBRCHyIwKEdgnA7DAeckFl019hzDo48ACj+6X4xNr
vAIc9EUXWVet0riPM0IRthDhzjl22Edh+MhiljTrVdTRluCGw7mgQFZUJsj8Mqpe
jDFnrIl9wq0vyQ5+SOHWwKzg1xo8UNOztilnSqcYYdCmfhwbtPMDZBRTYBeXhx7M
1TLA6wcQbMXTkgyrJv7atDWXK5b9QKHqYe9/6MYuPVzPfRheamsg82MXHP7sQYDL
t7zr08vDzJ+FHpz/1nPK9xjDD/89jJQS4oSFAEWt2NMHiPpGvbbKuCGE6uCnbKKX
lbZWbt0i9y6Jafb7khghEvyYi29kVOoraI6sTo40/bADIrOSXsp5MqEnuF9IQxZK
Ts4pd9y9BBIy0c9zFKUTWK3MZgkVZiEA0lxOkXhFcOJWF+XtCgb9QJoLMIz64WQn
2uNtZjD70SSW8Ant9iBimIaUtwFsZssJ+yTVODsI2reT786JiPjTUKotGzEsuk8V
Ni70csMq9tEzWpE6AQrZhzie2XMYqKlTW7F9IMBktwZn0y774zCW8qY/r8rnJtHW
i/usZsYNotHxUFGAByIaSXFlc0SAFTWC04mqDtfIIHFwAXbMoeJfObfO2H1NKBTD
dqmGnflQGMgsck1GydeYRv0hEprVTQLaTUWi7/UTUmprU4EjP6AaRkRKiLAsQFxt
IwdPWGk9wyQcy4854yUO5g/btkyBL1oUyHVwupGvSWjbPhn7sdKCUXKbtT/jL2uV
riz11Ts0EIsIHVhaasTSHk+oP9L6jt6R13UdTELhCFv9tWc+JlAxav/tUEp1VIku
fVzC8MpkjNYS3+p9ynfbHquY4oOpm8PePW4RBx9AolMLm+sNddyUhFmkIEwEJoHW
tK95UcswlR/rigc8Br6hkSEzxoBI1fe6iJMToVgGxQJdE7vH+2z6jHUu8GGPvTXS
k+Aiul/1aT6Bs/6nic9VzSxX3IVGnX4zg+/qHy90Xd/rdC+ZoO9jDgSzPczbNueM
4I5XAqJmbPrY41TFTHz0OVJ/IJCHMd7XofpU/uZAFPWSMn/lYwhTWoIM6sSueLqQ
4qZEFqWRIYnWfChaYuqD+oojC/CviRbWyzIh1+k0QRmgjHzdlkInr2ZxQIJfOYj2
i1+ZSguMAOrm6ksfNaKyIinnsI52hE38A4SMs7OoZ4/LlXwkVL8aeGcBDs1QG1Xt
Uwe5sOEZUIYzU+kh1LxCF1ZgDX/kx0BHtf0qDRu/JBTPCZOdXHikZdfJQIW/bPMF
67hdtcsMBGvxfop5yf26QPxRiqkUM0AZMWhDVjE8hISqAYGyesmYBOJ3PFBf/EwT
jhPqPgbtXB7/PObb3J1h18ISjFiiSFkCXrAnEBfwtG1VnU/dM5n6aWEv9D6QwRba
Xl29SWM+q3DiEehmKikceiRuf3/R+xEuKKxswKiBqNmCcFHcBZTiee4nbhbRieUR
zFEaHbcV27tl9sclRnikwB4z+OWT83Zq6Ut7NfND06lVaubbMHsshr5OWy7b/FWD
A2+uzOxame7y+GAtQF05jNimqTw5wZILaaORS1L1FeBXOi5t5k6mVg3e9DgKEcKo
cf1R/o9qmLWIUSp+h7ksfbQuvDMsqLlTEANFciheQgtLkK22NOqej1wehS7hhftx
tHFTcNOW4YqQg6bmOFLkUx7FjwRuEcp1ro/8T3yEMGz+8rMWTEjKjaUL6OBHqKmw
CjAMfjT672hrpyMnGrluzWJ8195X2s/nCwaBTmCCwq2MECp6nnONcn1bxOkzQwoq
OjjWfWuCc7N01m7AsvIXGlU680YCu/kZJC0PT/qYjt7jG8e6G7BwIfW1GCD4egZG
sa2XdFmxJuPXGGl6pg/+fio0Rf/VWJmOi6s2klr8HJE9QPShQdOSXxuUXjns+jtC
T/oZ3uNd3bIA7wTr/8CTDjze1RVWoKPr5BEpYfpwYukGArDe1O7pUmapjamLUoto
OORmpLZ7WkTSIpHIQL0rRcE/BW6yMHcyEUpUawrjdbFNIpiXybsczuxs13YsSmyL
1eSgbIzpWma3XTk8tpAD49E3ju97OKwqoW9SFi4a84wm48e6OR1qbCIYw5+nUcWX
zEgiAEDwEx8YSe8g3OjZWVhpXwJJ4pcCAtfzuk7iNUKWb76sS378jFRONuapzNag
n6XFD3wR+L5fMMz9OXxuRdKHRLFAWSbZH4RNhi3rp1jgR2NeFG0fhmcs4DMkgD6o
TcmsYyjR4xnUr0bBhvCyKHEr16Imeefoduf7MorrplL3aSRWsXSpKlSWJn/GduLy
v1GfxFY9iH4ckxSSwGrqiR1CRwoyKwie/4ze7B123+oDDLgGQ1VKZj69Yq7s5Zw0
Z7N4me9SDIQogbJlDvf607fQ+zlju8jInV9/3f0FRR+vzgNIircMnsS0eVmBQwjV
1cWOTg4vCIx4V+xHnoK06Ti4c7cHz3Nf0wNmCetbNn+dDH86+pLt9bXaaM7FFt9f
kzNkKZU5M54wOycTlICckZvIsE69fH9sKU7rvkZ7LnbWuhVs6l9HATgk5fdbpYRs
d1BZ+PyjbY2cYsUTEnlh5YtKDpjikvWeyruBH8Bd2ouf8X6ByYdzsIq1YdVEWsXs
KNzo2PXLdSzUP0JWjxMxvHPQglhMWnaQGpjqkRpF5G8lAoJXc4af6VM34CtvwEO5
UikGoYQ+z6n51OchU6ylBzNHmKtOhLGUN5UIPNri0S/kS1HMQmf2xE4NStMKaL/t
Buut7wNzGpIRwXIOiN2nTlvvGL3Pbra2/EytWnob2SsCmlh/jruDdlj57OgYJiX7
CwBZhSndyqi0fKx3n5DunzMSXsm4VajK7O4jo6+6zm5bLVp2JNGWzuCe/JxZ5zui
cGINZikaleE2dny8qePWWY+TtzBl9kwvzKUKTxJX77KIERHYtsd0pTncvEZduMW3
uN656gFJ8gH5McoRtQT6iBWbRyWmBYMQvRWas5A8BzM18nTGNXfOePlpDmlI7FcR
Djy2/7q6ZtHNiENIgwgaRwnXO5eVnNiSMeBut0xt143sO7wxGiWOfoh3JY2EicX9
9+dTU9wuQn/Ft4tfTpNolBjNcTWW6sJAX7WKLyFgHyYsy+fGqRa+SQPTONebdA1y
Hsz2g6lkp11rZiCjcsNLedtYejBtc6d2Inh7UXok+nLQTjUCHcu4YzaIr4YzY2d8
7zm6frJ6EVLwBXUONm/POGcNr6+lwJxo452nZQpbzr6oa/V5cxMcSSd0e1wxKT7z
UE5nnyOOa/0iWL9EwZwG8oLAZbmupPD+t9oi34ei51dfxdYt85GB4F9UL7W0qR2x
/AHAoCOSyMPmH4oU0nNEgJvyD4y0vuAdwLsYW4eKri+thjDTfKrVmvZgRjtfHfN+
dRiSKFFcUAxRniJNpzMYmcHwupomOrg0ltKLTSPxTUa2nu2OYIHYCxKialXD8Jf2
oJZEkES1bVjLdPP2vb6fPWlIAFWoyehEyGa0yfaj6WND73tP3EXU+flO3mFkRln2
CNSCZbjZHzaDN+V+stKfoJsXdjJtn5GZOi5/vBjtHGJ0YKvFF0ZySIVOXf/PaKxq
zFmZ73pUUy6JqkJmuRYpDuFL2cFFD6FhshrvmB8NindFVuY8zlWGjVhCUdUqDfj6
XjCjmNCw1nYguxHlBMzIUPyM18hh1ZUe6w8c8TIXz0eE+30rKL8yCqSifMgQ9PLm
zoZXY5NGbGC1mDLBCst4WuH6G+BQkCA6o3UG3/b5UAUn9RhzeZznAsX+yRUhWp7d
jJIYJYCQcspKDmQiiw7AhFU0ajZp2DxuipsN5a9W5zeJbu2zHqNemDg7fImHc6v/
Wt+tDrC2CUyGHEmJtu5jCAPlSI/J3N6pTxVS8NxhyRqRx/BWWMt4l47k2sFVi1jL
iwX7UNKSW08Jj1eHTUuylkAGGNwL8UVtqSBmSSK8UBITuG0lyGMlXxltPsLFLMfQ
BriY5LzwQXNXVr9Ubk/o1DlU9UAzTio2beDAG+biB/pHXJG5aChtJpYYpUSue9dS
7HgYFmhtZJXChS/iyTk7OlWZL0YqqYDMUhv8irMYOJr36PaBgYLtDeqZjYcEMc+1
RFSuMSrkdMpb0ul1MwdJP05cDN1hF0QWwMZWc1VWlWB2oSHBMJch9Ndr71yE5gVP
5TvjU+/dCu8k5cx9yUAniNuSdQ6hOk53XuXB4jORcFzgt7A8UX+mW1dz5WXVWEML
cvg9Premkk1cOs/oEPj4BUNsLUlkqqBTsbisj7taW9H26ZYki/UK8PYdoDKudcXf
wlHpYwFifV+22bLZKUaDchrBR66rDvqu4bsMPWkhyZTKZLAAA5HswPWFtUlLLast
5gz0Ha/AJqOhgEhMqybSW9lpC98h1bmZ/qI7YJseYZs85aWDqW+ocJvP0+bMLMx3
ndY8OhdOoYcJl6TxNWu8AU+7csxQVNEFiwXIil+dX8vpIAFDcOXr2AwYtGt0OgaL
zAgrPAG3avAfYiiJNZx8yxcBLwId0cmW7yDYxYyqB1uRP//fY+6oCNhlgXHOv872
w+NigINWjWwk9tb7kydWBcwRvy5SHnHPY5lahwPChujYFIU+BObQsQWLtDHHwD9o
YFaMfZ7OalAyWYTYcazlUF+3GGm+p8OfPyCSek1wdUzE8sRuQ0Rn1tW8hCf2HvGh
LAk0VmfGjCGz8sV30nsJObZbWJQQM5PS1/+gAEMOyGCjqsoi9BpRHG6eYQ0uvfEP
00u2QKD6ZYyR/R/Xpej17lMAL1j0bfI0k3YN0xxhC5Qu+XabzXinICO2TTwv7Sml
e/wB4GFLc0QXB5cnNW7C4hjK1NnOZ2wEMdmToqqD5OOkHIN+PjDc1HnyF2Hxs7MJ
pLk2M5+CkySFD3aCgBiY5nDMeGkSH3Sg44VRxUjcKVEixfwnOzYd7T3A2j+LnpjJ
ZeBNsiy/xlod3KiMTqb22iYQbAHBh6TtxVXLWfgL6c8imKSGGoHIUA8uAz67ZB3L
JfYCRpHdDrYT5uEcccwbDvqmSBzd2WXW5HlCpenLd+gqJiJUxC7ihJlv/z9WS1gS
3eSTmHt22WAyZYEacB+ijEpsXrFv7N60GA3MxNy78N7ktVqJ9+RIRC9RNQyTLJR0
tzwl7hkwgjUKeTxByu8FWiEyrzNKqgD4DQ5bMCTX5O57Bs6rTZWnWBliOPHr9RHz
xuLgee8qIj+zgISbuOg4R1xPNRQm2G8Xyifsp1XP8LtQf0wsYRZgdrafi3KFQhJw
ukYs7ve6Xwm2iBLEsqCUs7buZ3tOu+NdgS9KeuaxrsuhHSTpTsWWZ1Bb6iLt2BrY
Oks+PuFdmyR18A2biikkO+swV+cmyl3UXfhb7QCjP8OBURvsJuigF5kP1utAUEt6
ffdAln86Wt7Snlpu17EhtGZNJUbOGb7Z/r/n7mJd4hSyanqTg2Fc9hhWsJ1RnhXq
eLtCXn+DgZAVshpG7948Owlpq6Xjnp+hvrsbtc50frh+Wv/122PmolQP86mS4hbW
9lDxo8xJqoFmc9mhaPjN7ysx0gwgkwoQUyfpkJorCXi5nhZ3tnOGqLfBC4b/MYNb
kPJlufclo8RO1ew1JRkjegPBgMOTsNOdrsZE2SUdyhuNEF2Nm1QUaFtrDz9g+GTr
LsQ1yfUNaBbwTvA7b7eI1B4F+dMR6HouPfWmJJLCsOpOVw3dzVRt9PVK0n6/DZlh
A3YkKY1/TBwgR7VO1bnYu2ewyQ87+GViGcFVBEyZc4pKKBsZSyXb8uNXnE6adk51
/F8p97YXNsEz2sJVsisSoeV2rGnSJGPi6KxPs/YYehxgak0TfY+xBx/ZJKcJ+o1l
NsYBYtUNOBdRaN3NA8tjTbXK0vjj0is1IhmNQkUVxn8KQgvJSVu0W/JCaZolzNXb
qnM5OpDaNHz/uqOhuXcRquMsf9xPw3/bygFG4PkcRDniPhJXpSEf4nr8DEjvXmd2
C71nsYfXxMHddFwl2BV47hrHQLrlVEgtskC6gJYmMqdIMO6Uj9OVpvqvuEG0e8Yz
avCupCVtC6nhUSq8muanrAJ3abQOSEb92N7NrAi4o9ZXlPcWPQJkhtoUjnRLaOYL
u07I8ApRL+/9urMHxF191keiHTYg4G3cAVyFqVaPVbkvLGb/GLY9W5smixmXMl2r
S4DU1Pmk06zonWpnQEx7YVBJ4a/co7ZNdQMeQ4Qf8T/1eelePnh4tVoHfjBBR3P3
n2Pqzj+yJXKQqMUf47haZ43yXIG+6E4yBwXjK3+t9WcCid7T1KA0SKllQRA/XIDD
kkMpWXvcWKlr/5NVkSDoMHF5nglLh12SbMEHcBQUWdZA2ilAsLOnf31rbFWmcpme
eKE3m2/3NYTMYWaZRco29ZOcScexW6HpC9CEAmcPDBozGQPuRSJonItDm2/NeVFm
OtOZuktGNUbUI5yG9XXMavwPU2YItgNMPlJjZYa9H2163nC3b1TfuvRWa3Jp52Cd
4mlCtu0/f6gsnjrCNF3vpmYc5rCdpXcgo6c6TukP6vbMeweytQ19I7J7KGSaUW+k
6fGds3G2rEmPsy7t4jM602A2PE889AFw4DWbG2StcB3bJ9qAGcBR/9EVK2FBxDxp
9C4BsgKyT3G52mG3mpoTISviWMkzwk8Yf0ZTiRtti6wV/p2ACeCAtSMaMXjSdus2
Bpn15yMWgfR0XK2rFL/pQXunJ+WEbRzey++Dji7li9qyid3W43GJBDlOZGBlfq3O
FEy3OrvUWdyb9R3k/ZVkWDW2RMQ+j/nZ4EojMEM5TO5y3H8xquBLEd+R+qeaihpo
CcSj5QQnYfxDBZZRbmd33j54knfnWuFlcgNR4itAR32U+2bAOLeE+QCxV5jtLAv0
Nuz04KgSD2X16ks98lCEq2vS8NuEUV1zTaV3A9VbEe+YZHlMVUuoXaOtMwwB2zci
OR4MCBeQ78VQhAYLMsYm1M7sOl/0dT2j7NhorAUl86Jc8vClcGNqDPMHpW/TCNW2
nRE0ckmq5y2FAeDW6VGtGKCgQvtu2ptAZatSRrzZ6QW0ma1tx9I0xcf6MtLBp5ie
sIv7vVeTtMaYA4cmWY067k6RiP1AhANArYx1sVhUxCScB05CkY735BhdsCqRes68
S1M8A3XkN/BB3TAYBKKQWpxzB7ZIaQr6rWQ/p/av6AR2C3C23F8S9JBdw/PFHo9q
sCw1dT8qqYaHjZ9mtQmtPa6ssLxjRUPeVsVi2y6vk8Xt9EXORqiocDgvzaOO31Yk
NZ1bTSf/U/3cPE6IR+4+WHFmc7Lundj5tijm65T7dhx3n0TtAKzmaLh2vZE+y9NV
sKbADCHqpDO+jLIS5LavCo57MzAnjTaUK5OR8MIVNT3Vr/yhTXvQDfmrBboMCeev
PvUW71zjaC7Rf4Vw5wxCmom06KD8/QFEjK8AtbHRl/SI0bHUNH6Rh21EhBna6VVH
kQ3HFFRr29XZnQJc54KqDX5bH/4XFSX5zVhUUSqXPSoFvWP/CvNndAq6vbCetWEE
Cf4lGJRnFE7ygFkUZltX+e+nsSM4EhSMcDO80A0T4Hryld/OF0wMQ5IubDf7ByBs
Uwrh8hJQuUGjxHOCP5jt8ebJPcYeRVpDRKb4zaqfFqo34Yq+NFR4IemwIechfJSs
76htXiJ6OKcl8a97+F3rUmkO2ZYXUT47jHjPT46csWCNOjB05E5f2ZxirFlR9Rrf
+ZnK9ZlWoN13tgk9PhUHs1h992ulYdzrW+kT9FWH9LDa0eKcietPD/XBWCAEFmF9
cIVfMk2wpfLqgiWbW4QB/AZaJIzYLynfpIk0i4O1Z/7YTvJZ+bVx2ORaNEWZ6RzX
FxFtFoDWyX8K1h9Wq9lVPTh9lj9CszJNwpda9FDjkbL8H4EHSrwVBVeoKbcPtdTw
iv66HL1ONyuguhIG7L2jq2RVTN0i6ZoYTCjtIxyx9lAgJu+WWX05UQkFRx/7lFkK
1eFUe5PJyjp7m5TZpgiG9bxssRAa/HtQQn+woyskAXutkqrbojyPyMB3TfJEfz6F
pyhyGgHozZQewt0afM3bwE31wEhT+pW3wuXs2lcb7XxIUaZb9QpG9Vo47FBaJUHC
484CLhcSJMAaEK6M/Q9UlVIBdmDlPddKTUwhqydoziNWgo0q/rImR1pL6nipD8vl
7nyJJ2GYpDA8WFxk8AFMo4TQQAGtD9qy5ZFEwnKwmt4OC8viq4oEQHrVC90UEGFM
rMin7loUmJdOPOB5FEr/oSfG8uJQfyfRWQfc7/1lefYuSbx/jjqM7E//Wnhs6yCm
nKq0R1c6TWQrRTT3gbaYDCA2BeNS5JWdnFTzqV1VQX2HFHygBLAi9Nk92hAtHmtz
k1urssrZnQA8EfWP0NfcbbiKIHryLaNlu6A+zjLafus1N/sRNZ22icisu0YlZPH1
j0IWtzVtIgV98bkAp/sM1dlpDTYDtKExNK+wvEmKv50G6rHLawlsdiJpGT+puDaL
BJk21lzdxTjQF5hWOCbvxqHmWmLSYwMhTTqjOckzW+vALFFawVDNgJ2Qqd3/MG8U
thplO1AkHMpvaxVl/FaG1LxZHNMc5/Ky3MgJxHhpfm38qVj9P+Ri1Y+e0t4/T7H2
xsp4rMYl2q9O+n7XGmOk6dnwp944oitkoXsePDvMlOxjBanZePNK2vCdJO6H9Hbw
aj/qzrlWeS1h8beC0r126PmKVd/IEo8T36b6drMdMKxWRlbv/T37MCsz9Ni5khfv
6hULxsrkttjZOYM4izPxKHLG9+8ZmWuxZ4Tl9zuX0SZpJmBQ1mfE49QmsSTUEugR
RnpxTiXOhbSBV628pSMGBQadoD831prN7TshUGV7Dznhj7cHjHEeafzYtVHo4H4Q
Kuiw9xnSrZoK18ktBp8/zKRGYFP4KCrCwyJvXGpmUrmhXoIHTtbbDRtdi30ql9D5
n7KqWBh28Txs/THgcxQaJ/k4mk/UJHSykW0VYDmxl6knsvae5fVDNIY57Y9hvk83
U/Yaif9ZstkI1CeGJk7B0r+R6xhakSQRTM12QbUY7FeFzWJaNApXZIhOEY79TEaK
eaEFBhLMcC7mXKfEL9EaBKFhTZdEypWuryckofjG2rrpcczWKpHvWYxCfED8Q0OG
ku4UjwHK8WR6CrIpzMNyXPFcb7eTzzF47yXClRcegc71dhWtneYV98LiGBl5AQau
C0mux2YLMMoh8RrJ3wFrR0gpaf/JIHknuBzPPqWFNxuCZ9JH5/FIUHlb/JVHF3Ds
RYEY4NS9mgF9vsu4zrjpdiYqIGv2VP4TJN3oGibF2noF11tDH5tmZmJGVDyGsdC+
siWNSloUoZ4PTQ3kemzx/aCeDVWnDECuYY/xjGtUBPwXzClquwzcLNhLByRKk5aU
dj9k4kf6aEUGvAv+UEZwc4gdT06CSmnb8zAPXKS7ux8hlMiU3A4FTJvghYLR9xM8
ERXDujbm5ZGtCa85homSla0VDtFtUnuokUDpLE4LJZhWD5hi81ksMHiXJdWCguot
eQSqXDad/q/gzs7bUBzSBC9vY6069F04W236xro9EzDYAT2p/B8z0SiupWb7u5am
m/G/XnUw2Mqrr9LRmVlbGXW0zELHvB0hSSDnnk628PieSSYkslU5UjvtFpijYUcj
+auiPYCNyRvGD9/s6HmaVrQl/BpVdyx4YeNKeeqZKQ9zUC4AIe5Kr5ONxlxmu69y
Kid2wNQxzFJgMi23v54pLWstZpmIdrkfwbTWrqFBNv2P5rScUclhc4kyEKVMhOTm
6FHhj6l0iaPfqH1PhhIqRk10jql8kCFGBj28SOC8tvMZ5gagOpyqGpW2l6Yb6HwN
1WP6mHoVGsLyO3N32vGsBx2KleReeFN5KZqm0BFrRfqBdvveQc97ZMvmvKAQZG+C
sqRMx6SvSuqXRXq4gsaMBwlDfH4l+2wfmqtyZdGMfv1J35y1yZKFXpi8M9jIQbSX
80Olowt6imH7kWPPPvK6xy7RRXYNbnU3govsZ3KcBi2Dedpg5RGWfAwdlgIpaIGT
fCbzIGvpl4Vmy7NovJ2E4BAGNYtMfjt8UxcgAHpFLzZDi0kjKJDZEiOqTElJ1+X1
2IMsiQ+kE9LgxKymEjpTxEtCGYkX66s26sL/5DkHxrj8gU4ZdTgrizzWL6Hghwwp
MhXRgvePNwg65v6fWLNeZB1sg6x6pJlZ55lTHdqMgZ2uS0GLZQTRM2VD0HaIVy//
5wGf+31MX2ay7rs7BCt1rJc1lFT5vJNA7PsNVCVIsSWTHz5feWa62tuLM1kops8l
3syghn5/JyoXV4Jx/DSD7xv/kT6Zy282HQiAB+HNtBHllkywI3kvJ3pXNKr+KG/m
k1/gJ4bndG1U7MXIqBD/XuzLdLEJBP/lBCM85GgOzxcxgNgt06lxW2eS5empZ/eg
B1W/ARvmsH9hvuvBTexKxv+7ZhcIOoCw3z57brNcbkjv07Yu6E9+hGnDtO7HXBvL
ekDtlz2RL7hKnA2pL6CG8YoeQEafpZra9q/nuzZx+wzlaTILV9nQ7QaEG5sVNEHs
B/P0kqgjvCge/HLa5hgwO/RFWc8RfOBsZZI1fvfqPl+WzDKq4iS0yvGMkZ9PQYfP
qVL1bRr5RJ/a4D/bx9hUl2gb4IFwQRhb4aAlYOrjDhgUBknf0YEieCoAfLtEeAGw
6SKjk1juF6jZ6f8pzaHn5rOy9rJGo1cOg5rNBCAIjofBM2ePVWwkzwGSnlz4Ngwl
Waa10dVeOSlrAOXAJ1GC8RYdDmT2wfaemr3nIvOdhnt2nEzrfTe6BDvqN7M3d5ZY
06xUGbVlnRV6nfDFA5B7H5m9vcJGOfLuKpyWWTnxpm0pkCzx0kEv7n5kSA4w7Az/
fPFfagHoPh7+qoFhf47OzC5E91vqH09tiMrCwMn0MTaf8LeK+cvlEVdRIrj88Nei
HAdrdwQatBjhtXoz4iXEJVwrTWjiaBD51PLwqY3mR+Dw5juKGEueWbthn6KsjSt2
uZ1qC/9QWJJvGT3psu9c9xwBOs46cWa88eQm2u4fvNLFbi/XEX1LrJ+xWRAP1McC
svuj1AmF6QR4eaiIkmi7n0HS9/CVWutMR/TYSOLLCOzOPuZEmI6WuNOPf/uN8pHc
WfJIJx/WIIm5zzE23yIi7WBS1LvvKiEsEWatQaJvDEW4Lgx6vZ2x3qtfdekjIVhK
i29hDMU0oyZwpMbklkToKedWncD9uZ+Bz4H+3dPtZ/MzdauC4h5Or0NKKlCtE3Y+
JhyKXefHP8OVSHeUsOrhK1NAzGzvkbjeOC7Ako89RgIxhuk1Y/FpYs18/5RvdiKD
TOigx71dz+HKq+nVlcNbF43DIQTmztsO16iyqPS0YD72Mxr9Wv73N7Rl/pkWzM0i
na5CN7ApDmfcZIlV+50pZRkR7eRa75PztBN3YjvbrzEsDvmC+7l4P3b0zhDf6ScU
hSNh7J+smyzrsWPC4MQsSooKkWGTQ7U7CGMcy6OK3aDWGxYvF1B/DP09Cz7pCh4O
7N3hcL9/82wihm3A4720k5wMJCV7Fds2WwhJcxtrbiv7fu9EpYpru/Hhvk1rBCJF
siqiaRuQoWOTXnG0oEMtm+GNEXEZK32a2wIgaau8dCrp8FITDJMEOou2SqRG9pC6
4BI98PQq8rE5YrqWqF+TKwJu6wpUm2tXvVIQkG24tRCwNJu9O8pgKWfPE1TJnXCm
PfWeUFcDvIp3sL+cyT7jOSgTw2yl3WrI4/BGT1SXJrfojCfMTk6jlnxsyZYpNCTR
ooa22/aaFxonYGP9sWJH1/Z8eFKR7jAEFqFCpZG+ZX0VJ5GgtfXOIW23dZ5EC6Bg
2wU+b6L+FYlnLVUdgGai/uyj2n3rK8UotESLwEGuodhJUXPgCagv4jJORfTfOukn
5+TB+6zeBcYpQjBuxrPpHw4cLxrMbCOKlCkrWcpHtK3Ftu0y1IjivBN5nXZ4I9yv
g+Zmk/TI5ZrTX5cyJ040DN7AG3lQpMckHDrOvf7VrMWsVFb9Pc8SeWCx2Wjzfyen
ZcErg4X3vqeRmrjbFZoe5KpBNo5okECvhsbHeaytt1/oDkucPGeADb/msoIwFehh
FRzTLCH2AO7ZmjFj2NsV27ZvrJpYP/y27GPk9FgMN64tTGKWhdqwmq2rM8kcw3IW
Pgv/3XLyEgbyPjk753ZL2XGiLPG6mOU6t8zeiXPb3CZUimPEjGmTRMy4EUvc47r9
YTrmKSsBflu5ilV9UJ47fAZVIyqPxeqid+NXSUMJbdStpdqKzb8TgNrbzwP6KPvO
BZKaui4+IR119qRmcWXje63z/k19E3bpHyA3DpszLdBVkfKRT2K2mkSm6yBr4IBE
8K6U+/ElxNBr7UZnVHaUypM5E9EGvjHr3iEvhmi9zFlrqIb/h0Tm+dp7XtxHBi4/
TNZdEpJDqygo8VgtvSXQzzveUgryqjmWD6W6XKG71kYrltJbSeJl1dCNsS9WkZYH
82VQF5jFilY6Z8vPq4OXBJdqZZcae028Jlqr/CCe3uMc92HTZZcqPFhtGuTtHeOI
y9DFvWXpR77BE3T5wjozG4xJ0aSnKemnnsJp0I7waz5a20FJeC+yqP31Fo1riH9Q
EJFl+h/lL4GJYGq3nVo/Qyrub1yXqodWCT/vyKm1Wwg6+Z2v9Dqra5amcaH4ko3U
+k2loZS6PoEDFzbGrbgAZgH3wtXmzte7FxBf44Bi4paW+aXclQLafudVLXAlP/Ga
HbBB4/BxQXPNElr1FYaJO9a7NIEIpnF6lWLadROtqrDnhmehJ79DjJ20x3Oyk0OW
HtMJRBXi4T4o7fOLwjBk/hnLbYyG52VDvcU4xJwXjirFQf5ozlFvUMCY9eX1iN7X
HDB2Ia+0/UsOGNuWkOtxczN4iF2RezxBpB9kq7/OA5MJY2NFeyxNY8hKV5AROJ5V
e7EnX3ArNIHslL1GWA6sp7KBsM6d8QaPZ6zFg0xl5h3l3js9bJ+k/0EC/4PW7l58
2CZAdXT84KNBiYx2i1JNKevmjLirP6X6aaa1Ig++bXhrCOpJ/A+qbqcnOo9pPd46
Q73IHsvizVSP+NyAvNYO/dt4WDLmejBNFMO/NXTIREcaAuauhx/ssvzNdKCqMqIz
Vpr1vv1qAIxmFhT6WeVl3WDnSFVasJkBu4BP3qOU7REaMWfJSsikB3Tb4C3AzRCG
V9MZgJx4PCrwAzQMqCDX+bZ2rkSJdpqKM36vqlw+i24Ytqb/fBeJiz7SRICXauFh
6z3j6j+0cbOgFMZb4txBF/IMJfyWUURmnF1BDhX0tzWyjl4Fue8SgH8g3vReV37+
jZLIN3arNPvGP00FJIlmXDZ2EduJMdRudVuASYbp0Fjh0PdyjM4bqR8W70B/OCxl
jr384stcXCmh2RUHn53Yf6vXqLwmxSTkHFDyPJ3FerSPTSLtaCVjZt3g7HdGJh3P
Of3AKSRtQ9SYllyIVRH1boOZ4Idj3snGHzXk4pHMgd9qVA2HSNRD+H0pZdf6H7Vl
It+O0WDzRdoDjw9oz/FG9qKrFaEn1tEJsCCxc0Zpu1QZ4BUY24270y38yGdPoRFZ
kLhVLCftQZymYnLha69szZoRyCXoGFglMZQYOUr2v+Hp+Lsf8Fj5KwCOCqKvXmGc
Pd2wkFWGtgqapJZ1rMXuf5rerHE3lJvodwmraacMPP4dq/MMVEZel6W3f793nUlm
WBRekOPXQUC+D69OmNkkZT9zdxVre7WHt0VPekcgk5Pkjk/3F3WlVasFbnDtFvzp
cEkrotXV72ye7Q7aE4HcuKQZxVZxn7hDyD+mcOa0w/Ek6etWwMdgG4BkbBfNbr6a
Mq7yEqjEkJghyO0dQXtpgP6FwXPY02uLThyravT9Dhg5vcWtI96XRet88JzaOpMz
DEIBZHM1m7APR3UDrB1kkEkAB0iKjTscXMxySnPjr/5ZLO8D/Wts+bvET1icS8Y2
e9avkoyq8T+7S1/ekzixiN9YvHj7KZc+/GTo3PMa93sk3bDFZw6SlIEBOV1wgL2i
aR0RtVkNMuiuRGG3ZluOU+XspeUW4HvrNijeVE24c9wBGGpi1KMbefWqOIwwyfLd
DPlsRsLcf/qOVsRDG6DVuHL5iIBxc+1j1Y2Odx4S7RcGKUGi2Ncsv6uRM5MKWCeE
onUT2/SgAMdEbdWreJwrHxsU64dWYcpNZ8mhFAxMPTjipWy8sfTDSNRsn68lkqWn
GwnRPpEhhH2mqC7gyWknAZMdKr4RW1oZzvAp3C4rmfQv7K8m24o6huJaLJrgncam
3Gcz1F7FsADvtlgmm3IEZZ9UowaEf6Zlr/zf4UU28F49VIc2x1h6MOTwN2VLXI6Q
zW6uQddAaxeWIeGtQTA+xUT9M92ILLecAbwRWhCb9jGVzAmJF/wZkh5wZgyni4UO
fakHhxCR+gm9Ukg46GeRJ0OQqa1v/AFnzptf3jcrXowYtbItp3T8ar11ZoZG/S1w
uFUow3+nSRTzDK/OeRXS+gjsl8sI9nU1Bz59LZR/6HYjdyh6zSnrrslVTmrSz3Oh
8BxvayZWyxw9/3ZvVA7adIIvA3KdI8NMYCLYGbmpbnxR/ASGa5wYYZE+rWwhUyct
wCGXegfQH6dP1tEqmjvdtoDahG4lBAw6jb2/T0LTtq4zW1JoGo3nwBa4+YoWkruw
OWWParAXZ8Ddh2lU5GUa/POppO7uc85u3Na/cvSliIFF4UZ9tBnBmfJr5rBWJOMa
CcFIpd6tqqmXdNAUVBX80r5xeyls2i9Ldm6LTHo9+DDNzFX7BfEbhLuWRePuNh3/
y7HA9ki3QQRqGG90UNP7Pi95hUVM7/EhM/LIuR0RCbGM8g1f4PyYJ81cJT1V52ai
hVoqtVEwCZUj+LxtL8zf3np/0/9qAOKvYd531Gk972GSH6GF8I/KbtK9j989oNEQ
I4+ljyYnBYdn1mVOuD9GewH1GC2Zmlb/PmHYIphTQOzstBdAvPrY2uw22Lomzp1D
/aeqLXV40jqZKWfYTjGOOaQJYOLi4nQ/k2dJ7UiUvm4Aw2u/TA73f+gCFC/ERFUJ
+Jk3Y7a3+DOYv5oKKjCPlKu2Zh+m8srmT9F6lN7SpT8WtRZr3oyahHvk9/veN36R
zoO12pGFYn9PAuQOZnvdcaCV3Az1wM7A0OZnePg8+2QeQvyy0hAaM3gzU+KQgv8Q
rOEjotUVT2uAvVkbrdq2vtj+wKomU5FWeq4VUpStUUoosXq9+scoyU8SYPNUEDAD
`protect END_PROTECTED
