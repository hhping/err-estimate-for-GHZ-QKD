`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiuTIOMfcPFqOP4OLzwasoPpE2b5krC9httDz5HJDeh04DWpsgaIzon1RnJWtL5d
SUWyUjYOCJXaV2Q2Xzgk9WoPgD7/H9RwrvStYNX/eQsrd8g8lhrcqx1OUPUr5r5R
p7fObhZ15+NnK+5i5BNzGqKqyb7zLIePaybnroFPMX4w6chMejW+u2Avc0bRhav4
YukNAmLx/49slrgkfu7cu/e/AM5aM2Met8WIkzu/ovylzRJUzlzTzShGrVGr8RNf
hskC+RztK1Bi8MU4viuCZOgPKxeIdiCQy81q9ejuSMXnq91AVJeneKg/MQ+hOR1A
6UQ89FuPyczHLxnxsfT2OZBgoJllzCz6i3SwVwUJ6vXfC/jwGgeKLxZWe0qaWoam
i5j2f9FlgzjfQ0ZN2RFW+0rnrZepwJkIIGQyZwGvXJIFtEd6joYYvtI+8U6XecIV
yj2sgE1evCs0K6eL3hiAhPPrTFeM8g9qix0i/gzyj8CZgdR3pkQhF5EpRYmDM0/v
kQoBU1Nc0g7WvBhghJrwP53bVwrEoF7eFEtxIaVxfEmV0oKnoSvtGtqkP5s0QZ+y
/n5r089vVfv99xLN+BONTi9Uh45eGWQc5ppwe4o0x4i462Czfs2/XflUh7h8xCTF
efMQVKEom+BLp4/q9XEPvhkdL34jQvzVLofJw9WMZLaDpPZvIjjyTtmNmTbe4nhB
cgMvOjgR+ty/vGON9zkNjpesAVQQNXjJxP4Ef7LutIdBAW6y5HVkMHxGCZBXydRN
J/Veaq9gciJokOgcIRBIew==
`protect END_PROTECTED
