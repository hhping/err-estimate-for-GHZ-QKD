`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jX1C1W3/Gh2zrH48SXEwdomQHww12/xVfpTp0bebuT7tQ6gEfDnchL/axIeqRCgx
a6QlgOpNZKzNb7RebX2Ik5bLsjhQRDrp6KzgY89gMmdjGVA7TN1odA5WWKw0IUI9
VW/Mdzz9geuAMzOEIzCBIUOa0FfoeCvcDB80fyR92ERWDMpxzFiW+Odlm4JHRwm2
iF1ogV5u520GL+CPTDb3k8QCvJYouafxaofxoHSny9fNe2hArSNZX/vpVq+jptjV
tkotqEfvWFJynLeK6HYOBIBK3Qjg26O4VMiLy/laUefFzIDlsp72hiaCbEReojjR
Y59eYVwVj7MYsYWBzL27N/fMSy4KkJ8A2GWTnNT6r5/w/xKdsGk80WNC9scow5y7
Ezor58HcsITX7AjYlI/GutNNmYAlQ7BJXMvuyre9dQdQiqSCWS9V/79qMknn4nRI
vNYr14wEJOI1x7K+Zk0QXWPlf/QOaNCAKLFaeTTyWPnwV11x6yJ9uOf8yug9JXmb
35/9qUsHZzuE4KxZkZPPjc29gWriIqFXjoQR4JmPy/zR5ft23vtQpezDtR7Bn6HU
upjv0GwZ7VHONsZm+wKagpfawd+tjyjWR9m4xhkNLR9U+yN8ey1WDnY1PuI2N9sl
WskTmbVb/B8wCFborcY9pbOTDu+o6Hm3O+L9kAa0Hj9U4jtJKufrD38lPmUw4c6J
SkRytWpbxpfszKlM0m4nlMUcr1qvxqp3gd78hileLHwtRe4pedeOX6ruLsgZ934O
ZBnlRUQTBh4rdlOc2f836cvV0vP4T5O8LMa31EPiVyPKsJh4p1I9BAREFl4r9HA7
c1tL7PmnwVEmMeT63yoSog==
`protect END_PROTECTED
