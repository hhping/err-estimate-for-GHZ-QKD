`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54xYl3K4nB5gpaQhXhiryCjkGqbji3PkjAMAIVMVP9D6I/mVTAx27yMNLbhBAnXV
LnTGhBhcpu6F2K8ie3W59cREDkzG8lenRK7F5jirHJrKCsb7IpwdrCfxKFYhQDJV
qDqpol49LtXVX1NGIoaNjv2kMxTLb3z5VO5WFruywcB3PvHD/URnzaSSCyUjE9Vx
h9iiwA93LmHB+ab2nFyxwiqAnD1EPHUDSp9LAkKc8x5xmVg16WdFbuzl5osqLA3+
430mqcLyBrEzZdHcke/w8j584cRQN70yzXBhZodkW28hjaRh4ylcHaly8Wc9DOwa
6XuN1fA37qG9dIMGdslcpMxyUDnR+/aF6E+6k9PDZyIpLtHPrWmFadZVu08mVc23
4yRhSEfC8oJZtPebXH5fsDTBcx9/qsgOccMyCylrzSAkryFBOq6XhEtTyZgJouzd
q0gg95IFSICL2rxJ8y9eaDUxQXtxdQj0ziUtfudj70irBNFBDMkftcssH7Vr4vIJ
r+YtoyZpulQIoli3U3hRR10EAOwQDHIiNAQHkFaq1ItmGJZg2Oe80h+/T0t/Uwiw
wdrqTdKPh25jCOUNA2N8LecX0B+PdB2R7HT18J2N/+n35F1oJmEcu6FWMTfS4Em0
cW1hEErZgw2C3h7VBy7I1ckwWGYy0+o79vFnzKk7K0lIvKO5bgFbu+GK7VG2Ld3o
6pit3ICy0N0u+FDTVtRXTNI8PD1EFRq3pw7p/g1pSjLPQaMyUUV0q69dPyZlNpou
`protect END_PROTECTED
