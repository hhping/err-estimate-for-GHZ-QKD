`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dB4Vk+3DqhNnBK34rPYyCMkgoBlhBZ3NihKHLbkXzytENykFB0Nh4qMjfrUf6BEN
UAXsT5KzjptpzhckUlxkTo6KWAHQGQdOzAyqSum1fvtuxvsCgp/EZ+ntrmEtqSGi
3OUk8eNhGaQqTP16lq/et+sHyPylZ4rzz9mcbphcMAn/X5E6QrN0NxJBbcz0OzZK
0NwIgWHXnNe+vcr4vgpuWzOOfaQS4xjht/FJEzWvXSo=
`protect END_PROTECTED
