`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ztIKtchler33eKLmwJ4qJtodGrGzpi9uSSH9UZ1KmNMbujbwhx4ZjCCNOr2YW5vS
341ay9/OG5H4PrSxcDIeEGf3+HoIUmSMTyCYv//9vIVwbS1H3TpCMlILbRSZOwz0
PKyocNaYVL0n1AhMkUMi8nHZ9pCc+tqZL/7dYJSkzK4FJ1d/Yubuis/7HxnOkuF8
KWcCQjoSvqSd+h8r7rVUV300oR7HaWG7mv4XsWb1Z6mK8GutMErRYfhkbCB9dwwX
+LLcfmiQXHlyX8ibZzix7KrWy94brKj40nUwUQmgowcuyaxTIngmLyIrFPNwonr+
Eu2fT646cyBQc4VEPjk9AqRIQH6ZFC4OO8GpvWuXj9rYhnGhD5vMMw/I58I1ao3O
bclB3GApV/2f18Fj2hFXx7FzkCLHpjqt/RVr3t+c0KHsthsThoBNrPDqxXiCfwno
OvjRhvkJHmFIP0ekz7gq8/KX5qOWHEjc554JRRyXNTqdRXBkTEFkhkEpmMQMt6qu
PJgABeCKxTWLUvR6+va8P5JNWE6Qd2ObbQRHSBa/vnWGZgcYUBeOkPTMtVnYOu6T
ekJ20XFGIrGbvqZzmqnXYQRdu70FfIvRe+W6ukn/8JvkqhUOY1oJIwpMyaQMmDL6
iW4LcxVinVevpKHs5yqU9kI2+uLYvNFRdVnoWT8UAC6tBCa4ugOzi3ApToFbFQtA
kn29k21k1GsNr2tfVYuLjkDp0IQcOxM2VjXaREVntTmfApXwqb/iAaEeZ5Y+KRaw
hA9GidUW8SJMwRrxvhHJjMfn9XW+hFDojNQxTh77uQosJxg5ecU67xWmGxDkvwf/
RwyiKR4wMnKAplUKUT/brlCd0rjxwoHcCMQmHC28vE6WpUqM2/AtBeokWrPqzNQ/
SBQxd8mV2ND7z68K0E1Edr/s1HcElg4puRPwRVm65z6ZBkcJUuJ22S2UytLAYFxQ
M8Y2HK6P6idFkpSMiaGcR1dY0hmtb/SSnP7JlhCaajGonQZdnRlqcqhe9NSEuq+l
ySlZcBKtGoUW90jF5RWo2VW06nVbKiuNxf1hpZPF9CyrX0WwA/9SCaZ9JhE9vJpQ
91vrrJzoYE6Ki0X4CCLDbqE0lYLlDJWVqykWIsF2qn/wnikYpzeCHHkSYGnhcEvT
ORNOqvZJOUjohg3m+xb+slltB/2If7YTzAguEEMr4gKogo2iE4iZgQC0Aqs8N92h
PvdJwWW4gDcyWX3RLendBoY2qwasGsidQqQ4kZrk5AhGRq/UBA+OTWcO+jOVNItu
OzFR2wNUxFx4XG8gUHqRGNCyNxjnqoGgFP3CdqvvRaJznydg9zf/IItZGlegZHrM
OIO+4bz/v9e36ghzTK3lO0uiLmKVL7JpXiXBv+LBgbRBdRlfy7+YK/NgQ2U7AmgA
XOMOnmShK8iscRTIUh4GNrsf2Dw+sR1CfnbgRYr3X3wokf6LNghq2o1Xy8hmWjoW
DEvY8df/X9rzaKYODeq/brdQQ4fnhAaQVB+G4Fed+6BPhfkkQ1DBYKL0ihGO4wF9
ErD0Ucp+YnTrWLscTADJExysJY0PlCCSHb4aw5Y6zb+NKfKHS+hmhX+HybQ7KrT2
90ECKfJqkCGU5PDCMlcBYufBgpsufUEwrUpbgdukhreJIDm9+rfIelIQMaCmWjXW
r7KciwUzyxGW2bjd8HH1vVq7qRhf8I4Wcscw3Lh8e1f7XR2Mt+GxZiwz23DfWlGt
//XYTPPeW0qM/H7oRBtpLl0DK9oh9Jte14xJoxDbNXCisCRo9IMEu89qUGj7iKNi
/Y9AxPopIYpz/jIogwrfi+6qNoj793Gnqpz3ygKN0JB0m5P2ZuXV0ioKI7HEpgup
6m2GqAeseb3ql5IvTVw31vC5HsSzZ7yvxh/TLTdKuOlY++2EjEAHc1lLj16pNZ6Y
1avo38kSOm5AOn5QORGacTF6FJw+pZ6xonKeyTWyqi8I4nSwUX9IHrW2XlEde3De
M6PLBOn8ZAWxi/TAn1Kdo5PrmyHnw7PFoDRV3kWskpkybDd6FHgRgJa9qj14PDv9
M8F+w3wZThpdBLhtaHNYrMj7+RtVkMEDphkKoIyJap0BmZs0Vm9A5h9nwZRwknUX
ENxBlYCMqhaxVUsjyGhM9lk5eFNRS26n6RGse78RjJaxBQWj616l/1jF+OeMvsea
1IJod/cAEFNFgfKOBFntK8FphLbVSMwxWfNDCJviRp4vh7mCd8tWfbovzh70pFAD
daDP8525OAw/KU5bsHB5T9NTXQn/NsVWimdRrPrmdJ4=
`protect END_PROTECTED
