`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16XzO5XkJYXpTrWnqP4HCUuTLlRBVBbFvFKEeMwfzLQuHhFv+PlrK0iT6/B+G5xN
M+SqLHbyxCsyKkvu97en19m3QlDIFMg8OkECmIEKs59GfsYGc5olNWvcaovtVG+4
obJDOOW2DBDfHwyd8pb3Cg5s11r2HaZupmeudAO07dqLCcyLomLKYyNSERnrcFYu
qlhLb1AIuTSsYEHedxScS/zXSczvN7FjqJBSpVMenpcVagUktdqgMliddOXwXIYr
mYHno2SEDHUqIus15Ju6jk3LTzfRcOVR6O+3dMfQtnwGdmYCcOEgjgQYEP1+Rgk/
9tnTCNn+sXnommnzy++bI3Z2nHXlc8E8TJnkA9dakAUqNHmhZJCBLsbYGtosCjFN
veQ18lgVKOuqw2vCy3TvlFtdJylYdOI1pyhYigUZf6yfPPMKLDlaJAJPFdKnZV1V
LBSX9UO1N4KhZGpftlYjkfKIhD5vef8+uMs5j0nfZ6FG7vacRJSji8+vcphcZLrM
AV85aFUomhHGydcf/CiUfOO6MmETHgdFT9U3qN6PjuIy9Ij64w272fU0rVWm1s2e
44VFOBXmOIRG7GaA6lpxvGer4hkxOLOhV3NEcSVr/zDOSEYP1SCWFNilOJd6LJGU
YNuWNwloQVxi3aa+QuPA24tWBEvce502GLD0jt8l9/Lfey65ZDASBT4iEK+oFH8D
rIsRHhbJ55xLxRzd5Wkhw1zBJmM7oXO/+iua6QsNltN79Ic+kqwNAqhCDN9NNGRn
GGa6SxgskNuApU1HyIPMEt2mAxWASBzSlh6Q8eZ3GjTTtya2Ck2G/CHLaUhLjSPe
Nl+Pbhrz92NOhIaOks2hFMNm40nzK9zkeVtUgLYXf2Ie6KGc0fAzPXidyanXp9M5
QD9XFYKlpobI2C8dCAvZYyCzmNItFMRNdOd21LyUDQjZnik8AqbdLFLfgt9U2m3/
M+0JGh6u3cHqaKTbl62aYct3/B2nwr+XUYKVN4QPKj/65dFimiSHOf1fP+XgJJtl
PqnkDy55+GMkbvH+Gl2Ee5EHfs87xsP66LVe0d9JOFQr+TKm4i6Nmq1JgnDAhxJg
BljEdam++ZsHO/lkFj3ufSHz2PmgO9YJ7wp4UJgw/kZXOk/8cte0z7vMAGh2B8Re
A8BiC9+B969e8tH/WYlddZtegrATj8Wz69S/hpzOEOHggy1Jke0p99tGN31F+Ktw
9EfQ2LPF1TB/Vp6UuzdDW+d0IHNhYnwhV7DAmOu2G3cY/mk4Og8GKjeTxUtoJEwd
8gR5Y6SGBm5+3HYLL1vilwqCLuyl31vBu5XoAoXfgGzwgiRFZfoMYq+q5bWZkYY1
mRsf5OhOVFpxJB+r+7tgLxj+hxIlYlMa5b3rRTi6pczFudfZ68zdXnixSZpgHavF
EfrqTwRuFh1nDlLj0enihCyaK8A7WQeYygSAHkQg4rCchlvw8c/ChJTcyDNwPMC0
MPX8g1ZTTcZi/99Hj2bhrkA7Pn/58dSustZNJ3glvrUnq/j0UMQh00j9Yo1ZiWCW
h46Y7r+pbpQgWMRRDuI1LqOHbHmpL/0laiZd1Yrg0JPAiTVsIUHuQgYv3KDomkhC
GHg6hpwG2GixjJaueWBkjtIWBRYH45KnBS4LDAk39mQnoMdrFBO3zhS/coUv4UM7
8vyxj7gsmvfqmUoMQimWT0K0M82xPJpdBHBwS0SjoAhtQ9sc7N2egt06opScRAHO
6BSLMwXRpI1+ZyjxRCSJL3tBfnxEU77uOzR0s1rNoo+vZx6fii3yhuIwO22WSKZy
2It23ruwHMT6OgKwAe81fS2GpKkb/0TnfRPE27e7aS5/aWPuJg0UylUDLhVf89BQ
I9Zrdz8tscKYKrSfpUpdL9fOKxuNku2pnsZ8ZROeY/+b5yBwJ2c1sb0FhmBeCB6v
5g+Pjo4kEGuJEU5xleJ5ZwI6xqQ2owj2h1aS5CerIjd5lFF36FVLgezriP62Tpvs
RBOPfB+FmONCO8tj3WUM3Pxgd1G8n/2c8Sm+WZsoqgBBu4x2bJIUhQH8MLifoRhJ
Gls3/znwZEBqRwpcpKj6aSzo5wMJpKOKJug5jCuMmR7why+viWcWB9fOFXQtx4GP
JOkJLHhXjkEAnjOFNPtTRXxpwtxa3Shk/+Z3QzpQmeJrDtN9peE8XZTtS+zJIExS
fIA8DAMu0qx0NBDMWTliEbwkTiDLbLWX1bV7xOi5OqMQXEBcYunn+P9ao29oZuPw
DcqScSIWIAQ2iEzCQ96YFdCZCoIdhllNHFwXnF/4Kc95NOFPi3jG+mNezRjKC2BV
upm5Qt6sNFqlcWeb/BxI06zb3M3gdFPsq0V8agNo8Jjwt+P+acZsCbE62SmAl6tI
Fd78YAcfh+MvpaaFvgNm6vhqEG1OAmHG6OpptdpJCDXr6MXW8DVkIyzj+govtMK5
LRyU6BD0xW4yBVyiEz7H0SYOATWgnJe4lCLKasnlyj7N1mwbtpF6Kmf4VvuWL1V9
vhi1sKE9vxcIs/uoATKfUZQTOR5NBxjsPb2NqdZrF3Dt1/86XKfhVmrbXxXdIPVV
dOYN7dZMT5T5c15H9zxkNFqd/87VUDmGmR9+9iDIln/PsuXX1F1zEEEvztvzCjqR
ZSxIUG9e99cLBYbpcFPcPq+ZMvqEjzA1+FbrI8yx8pnlkVj4VnE0vLD8raZq6tSF
kgR+lPRmdydeUu5Vp8JQr/2DXCy+g/x4YNwlzCRuu5yz8s6SMzN8BEOBpMkXVIET
gXVV8RkveYQiV/TD4Zkhx5Tg0UCy8i7kLVDkCG61OaKB7mnutEnBG08XHzSBjrrV
OwAZCDAydVbkiTAvzj3UN5eUACus8GCWGyXLG3Nmpz8QGiT6+8dAnqXovL9ysdmi
6q2t9CiynjCTj7/Es/eK0gcoAOwX2KZZP9jlhpIh3GRAMnmBAgxchpLxzbIdhaUS
HggXle+S0OduWLOWNvLcDbmBE8B3ZB6VES1zti7ipk+A0sdwHf9Ykq8j6Jc1RMXb
mAi3d8jt64304L9TdpcV24QeodlxuR6V5qr6C0SkdT/UtpYifbpFoFwhmfg+elL1
eE87e6F/DU3wfR+6sbYI6rPzlYfYrqIzU3FkkQ/bcoFLcYy+R2jrvOXowDwn/NM+
L9pOqlcK9azl7WWzpgKwOk/FAXrcziNZv44Buiic1LDnENVl84rygYqrx1dTtXPm
pBTjXRQ3NlXSlnvza5JehHerIkkGQx30E/FnskITsigCDwHz9JFSxugl7bpiAOCV
cfIcLrw4Zf4rfL6ChYaer1Qcw3EeL09rgBV6Po4XmH5TW967WiFAYVv+jjgztPzE
teJLg4mUodOAeMci5nRL9U09bWVsCxkf9UkqPT0yRaFyPS06fLcl3ofklDvgsSfP
z7vE0lw+7ttSoYc4834cWP5U8hNpWCjMCv7G9SfJxYy1PfpwtzsNw5NwP78MLgy/
LXjqo/ZSBCwwi1/Gst4yQ2de0+FQgLPg7+QQkbFLq4qeXJYXPQ0I/I76AkyIXmMa
LudDajvmJbt6lQpRADhMyAke6C2hXxr+7e0gOIFuAP6ZacAvtr/jgXdkdlPn4Zwy
Fk6nRm+fxWoAdn04l5aasAL5XVNSqEmgwiDd74VurCQ82ZpMDxCMNFmNkbyv1D0T
XAat+ZdLI8wo0wYJxQxrA07OzhvStuYmf02AoNLkMBmf1wkTMiX5IARQYpYhpCGB
NgrXF5wt2nSNJ7CZZl3zT33CcWd29yGRvpyiaLZi+iKzwytc+ODRA5w/Ch8Ga7kY
J9eKqUlT1F7m2imorAYroCINXViDeJdiFlxBsKtFw5b7Igjm4iaGQU5xNenXMJVe
TZgih/X5L+c/R63+qsqkl0UKqs3PozDVLaKh4tzP9Dt9tMoI4ZfF7UJep04zeSBf
2QjVCMwMjkiYP3tmSGpRU+aecls4qmDy5hn/NcyNbNpU7ulYViH3lKxMT7uXzKFX
yKL2JZnfZWGZcWL7givLDCmG0EwLnjLUdjLOAYPQiLXwohpr4kAW4W2/E0AZh1CQ
jGeSRXh8tcDdg4y4ZCgxNuGCyrPpaqnGroco2G0xuQv2v6fnwt+37XsNd+qgaNqJ
nBLAxPN3zEHjpY/x/jkvR3xCqcofPjhOAACmFWsbKrBy2n27d7R26HNUS+/Jx9Ss
zDJZmmkcFBhyNKpCjV1k/t4k/kXxfO6oAS9q4L4YxVg4ub9d+Rixj4w7inIfumDy
5pcu9W7CKy0xSkawFGqPbBWt8ukblbOevTue8axEgkbUlD1t+LEy3RWjVl7Dd0YF
xbtK3y/NRMa962hzsNvVTx87IXt98+m0RiJxGFJKUDWrNDEG8l1e5toRL0mDoOxh
vATOj/C+dR+7KEzohCpPnG2UF9gPNVolMqNdcon45HPCMDtmfctn2xsPz/3RTkW2
ZPF0jhoCIQYhBiXm14M02zdQehSduEJ6GiREoubhMFsGk8W3VAs7hquxDzkDWsmm
Yo0x4QA9nc5Np4LxFaYpqMqvyJ/zxHe0ynSxXtW1zwocVE9kqMFK3HMhqsVI8L3z
lyi8C2TPzoTL6Qz3mey6of++Q+W6ck0F9x55+JUau0OPKdNb8q6z2FQoWyi+8asA
2icbxZUjJKbdltfW18KaFs8C/K8QHSvBla2ox4VGJPKd3cZVN82BYV9kc7GO0bUD
KO9tIXEy9/d9VDUEPG3DlHe4SefNmp0KiI7RIaaA276H4T2GB8OlEJsSof+Y7Q5V
KwWkqeuljiO2blLJ4qqEnibcoeK7/cMhbFVxPbAiHc1PjFPBE053AlXX10F5D1r5
mc0p7uNmVZOrYSD9H2zd/cPdsTjJ3HmFmA3B/M8vTFhLKCZHXZJUSDU3Nebczz1T
HqVMRUj3m+O7ZAHzYll6o5GZWKC2Pv5GWKQNOz2bbZy9mEmuG2YxlYPTJNpucsKK
+1Lm5EnWemdFxb3+1rx21+z89eZYgzrV+5e7hfaQA0YJKsFP2XrDA5Apr5KbBjBj
WN5voTEBqQNSfxqUM6uqUCl3XT8Q6kz9XYJyHHAKg+/0yW1Lijn93Gr6UjBB9MnX
5E1TVX5vjW0MJr9YaW4H0kDhGkiCBovyfJ1vIpBmV/V3fJgwANiD9Povnb6SUTv8
Gx86kACBxPZpdi8LRycb8lX9R4llyvoerzXsl6fk7oQpxV2WXMGccykfQJxabRyn
xh21dpcLNTmRDeewIqegk06EhNiuM8Cd0MLZxovN4QTn568A0txHzYpeaDHdpZ5B
fiaSQW97UcjQ/3AJyxBAc5y9gy0+LkHuPHbJDNPYGLASwFP/qewqtpx+ktFBm5Ab
SOjoh5RmZ30ancR1RXQW2wMneuvGpKNBkAkhspciPO7tBeWD6jc6o5q2UUUJOuEI
bwt9NhTyK9RoFKeQ+YcHqdkpSozrUYgjmT3Qzl1TOXzIjZAwwQyYp9gASvBZuSo9
DlhRr7/JyHErlKPc/WV0t2DFUOfdLCm066D1+3K3kJi8LuhKDFH5/ToFg7nro6kt
3NkKXeWxUrLOXt2Mcg1NcoDoWTP7LKITr/d+Gzcs4JSYPEif11BoPDuswI5f9Yq/
RLDdLVyuPu1aZm1otqUifqL0KdCZuWK1DpSv1WczLQneLYbsH8O5Ry5kZbM3X3Gi
`protect END_PROTECTED
