`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kn8nHowTgfSWWCRQ9YvWqOqoZtSDGCcWkBPik9jGRfdEVcq/VgArv5OZybLcAklu
yA9aaxzCN8c+rKhiC/qsBV6uQgR/RI9Rn1HNf0p5wPlFAtxymffnFINYrZSi1V77
NdgZYAEhIrRM6uIOOiMwisG+vXJGPqfKRVm49k4D4PqMlonmUrHRdMBsF9wQGyi7
cSHRC74T1r4gwntU8YRWwYE3QWuqh443GLWUuzQFmAI0pdvKVo+WPmGO8g+6dn8F
LvZ9MLVIieLhdxAO7efN1JWQLV5pYz4tjj3P2Tje7GvgkjFsJRkyaSn3oMU8+fnx
1SzrCBRLnNHwuy+PocLvTN5/FNw8nhwGk6kHzYfwxfsNxfS9LxtvOCB4Drp1Vyiv
8I+15DOmIWj8k0NszCXdXMgEc8iFdwqY+hB3iP84YjTuCiBuikEHsahUkZ7l85QZ
iujed1fHFRD0pDufKeAtsHQxgTKzeYEZdYJTkSWZLsRpoN5GwhSChH0pw1D+kiB/
D2RCqmVhQeCJHkfjP/E7hONrJpjLfsnm1QyAs9SYOyYKvAN7n4HwQz9Rhce0inIZ
ASVnwKCetnUcPzk+/LwaFwyZOAULex9lGk+Qyx3veq0FNSBHtr7M+BuopNtBUjlU
wjYs4F9t/XxBQdeGhRwqPRipujGf4IjHsNLzTR0MG8iQO5TBxnSbkOyWk4dheNbB
oTmmdkBK0POcZg/I7Cpk+q2UnRvqq7DQR5KIecqBwNymzTqJ89xFiAmQVOoBaVSk
A6nh5wlgIxnxXexF/1xC2xmZlp2cIdVcwx9r9fnBAoV6IIFwI4LvtFctorixEsUA
l5AFzm/UjtgYHBtyqn3ZUDapUWYnfAFqN8vfn1nWI6tqc0lOumL/sKW0YJJ0MJPQ
Z8BITw0kQh692kXn5SuIZnniSHgT1q2Eu0QrV+QXkEg4ZAiiJplo/wLt0io5BYgB
hvJYzsZeEpSEF4iHRajzTZypN+rYTYaFRJ5TqBt7l0k+1g5fSSJh7nSezJf1anFu
E4mD2eCtlSfxYS09aPB4M5co1a7i4Q9XLEE7EZDJ81h3SxZWvFxgWk25t+y4+6QJ
J4IkmUV3PMQE7kVB7Bmq2bLf7gTneM5LoCq4NHQGrX57ti6Mc+5YXkMKhLOeATWq
yqHMKbim0a1T0HkVdTkSiIQdQgjkCzHrNZHIKIzMKr8w0l38gzJSIhh4tAtahDgI
9SzPQR+fjOP1+e/bzBd2Fm74eS9ZQqxhSEVUpSpGcHY6CUyYCwZ4OQJIFws24gKx
dfCmr+rfNOpx+mYvGcjenr/TQTUqMeAIcuRrs7pC/CPqizl/N7+Ly+Aadshq4GF1
uOjfPgIK+S5BW7U1grfK/4US3ktlDNcYS5aOGvJInNznCrQMe13dxuFwHkQ/DYZj
yYCViShQCWWUXeSu8/umdBEs83czXOQXFwg/8Gwh8jjZUFqnpOuGk6Xsl2aLxuyb
+TjckAbNormNkCpowmrqJeF55xmeBgjxRmdBGUVQufRCnrX4clQKx1i+QKxeckLl
OomhSTC/O9MpMrD4KujhaqXbUj8lFXf9wlPWAd8ZzlERwrbxetorHAqlU3jt/DaP
5QPfrJY2p02JxCHFz3BzZmj6Sf/hjoVdnRMkPcmL3X47qz3aQEweF+HVtWROVhYu
H0GkKGYOofjgiBVyTkY1/w1M9U4cvjrorWVICGieB96+kccelSk71RPnCBj6WnbO
/ZcJYu4oSE5xJ2aVqIdhrTIGJ7CAYg6Y3yP3NympvNgGePyXk9xDPp2aD6JuU4KP
DyjuEJbSHLKpXw68QDQwchf4JRs/OJCHxcPJlbQNKW53n3b0hGiu0OXkP0XEqc2Z
NP11zZHD44h5VNa6eXkwbAP1Sz1X4+1VvrwoKJAj4BN16l7BhtvqwTuLAEvVPiIJ
mcr/VHMRHLkdXdO3uuYD9qNA4uNc939HR4cW/CtadNldehA2vMDzxBNhc9tNBFzD
JB9HoSunq1aGvNyUNIce4FOzLiu/TgttEb+TV0lDcNuemxsogNIflaitFYaDcmbX
5jwdBX6UlB1DPjK0Vq48YweP0uQ9vfxpK5h5p1pv0iJ9+wd9ZWEuF2n8u9fcgcPE
TOdgPGucR2Uu6s0s8B16/ctybyVE2cymWNBiyoyrtrXcCuPahJ3PfrGUZWMVb+km
rFaTh9UagNuT9Mom8L1ZxKHo2rPhsAnPE62Y8rFr2e+HRFZQ380/4iKi6U7brXdT
rMYGCJ6uAPt+HmkV52jmvLmeMGKpKOjPQ7iw1Q92xZVFUSK6Z/K24HmLRuMxYUfZ
oXClPLRc+GBkpx+Uws7mmcsQooZjECZRP7sV2bNj4BVo609g1CyiwjZxSkO3fL0J
Q6YfcO93ZSVJZg/jIa+p06UvuH8cA3yEd8vHAuxPO1xbkDZ5/ybzJ2u/uoJBoOcI
6I/rgFTrrdrgPbW1hsDdOyHqZTrD1HEMlBFP2WRdTb66lyTJDAbTzKgLhvpdt0mh
vimzyk1mwaTn1VdCQwisw3wZhKTUZIT7hpTBnInMjZ0r3DPJZ4IPPFXW4fyNewak
vod1mLKTbAvyvQuCXS6nlzqm9JjBkl2f7VN314IR6gwBuWRryI2jfogs3dcZcKlW
nNDe0bog2YdRAk56CW9Gd8wd/YON8KMLruCRgyPd0WWjaBNK6Fsg/uJGvtt0ONZI
TfvlnmpmhG2fibH1VwZQ02cSnrZUMwE95wiVCBx3O7NcvLMKrl0mLAn0X0uuSv+c
bB2Tpp3Kc+T9+vkv6I8KcC3uX6mcA2lmkfavPS2i8PhfnRRJVWUrxDXXrtErOjZr
oiWRUSzkZLiY1IKIKb52WMO90bg/5YAqbAXsF5DBWIAH5HaBZTfMdhCWaJO89LoS
0vxeu6NKbkPB/aIsFMNxPlCwnZoLCRTrp0ra47eawv+S0tcFk4REFFX3r6Qbr6tY
usFqj9KdrJLWpP8J8NLGskxJ5PsEgZR7PkdRcNnqG7opEc+egIr65Mzk47QYrACg
p8U9ELZUNAuYioHxlpmobfDjbv9GzuSPkbUBmM7TtyM=
`protect END_PROTECTED
