`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlheYOEGVRotCGZyOcZ2WPM1KEtfQYA6AvDGcZkIR5DRRLjK2tyLdqToR9sGPc1x
IT1uHfNOqKggjz7MkwZe9QZs8Z7awryJlnZCtchHnW1xOQ2XsKyDWSMxMUDkbu10
X/3JbZc7tDBvoFA7rilMHyx3VJQZvSHH5LWuSWV97Bc6pQxKaTccri6QRIAc+WP4
jJbWvh5LkDuEuQ1KPxiGx5G4m9qi9VHganV8ClqoA2vbYPRe8fMivPU5NVsIrGYS
/J4Em1P6tkUtJEybl+aQTKOVthJftcZr58jrS+VhFlkGmtat4oKcLPTaoWIYk73A
8XtAIJLTxatgPlCMGZWZSBCQkGSyDWmKkI6B8l3/1xNIpsRSexhCXtEcTypa6852
Lsf3n48RfQ3YGyfFlfCsnRC4Ob63FuOL8xez/NjxAQVsTUicmd8zDPmatOAWRCWx
0h7wfmEBDkME1YPfGUbo0qg7lNFvGvWwlIc86jDWfpMK1yLjpcfWyp0DKnwShiHs
w68juMF3zlReR2ZPZe6YfutywvgeErD6Bkdn69ZjU0yPLm/kaDs8Bf1QfrmHx4Vw
Uht7MIwKDcvjIx5KFrwEUOIWKBw4AXA8V+KTMfqTYMsxfnKwsbJwFUHyljFRRMyA
QR+gMuISjS6Sz9S0+JzHCGL8Ke9A3r5G/rg3b8dQiFxCpYKNY0cfDdy7aNra0Ps4
kFqnu/6zGqeoaeOPF6m/NJO3d6gIivaujcqJRhMolDx2EA7KozC1nLUBDKTRbCAe
uTL6tokz6jP/imVovyubvtdbeqnHH6iapTh8xXgzICY6CTWbOBes36eCkbwlIEG1
ni3iA62TDnJxhuEqVq+V8JJGBNp8WA/J/HA2evC726kWwI/sou5m8DcTcRAwm2b5
WyiB3/xWyIda/u9lFpO01Zsb6UIM0vi6CoLQsi69Bjyg9GS8pbP+qpIuEGkLFaOi
/e8WOEBtHc886fEbaOmILrCSYoy5fTIZiIxqLiYGbZSpzv0/oMfhG7MA1fu2TkQm
GXyvSJM/eXH8YzPrRx032Lo+evmaXimOFbKjAmjBRvMBvwWcBB7U0qcISfXfjq75
`protect END_PROTECTED
