`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pMrLHl5kZ/45IDCzWVONdNc2JfXJlJUXHzpVrcKnbx4M+xmy5X00FrSuIMPVZQr9
k0R5gC/pj7C4FEI/JdXnxZyI8ZSyqKqBsx0z+iVftL9HJDtsBdEfxTnJ4iVPMYKV
Xuoco+1INjPCdnj+lVAQO3QOsVdCPZsHZ8pChoAim6/brmIAoMpIdEQoPrNNqiHk
PVOioQA0JD6bsT6Z8YMXnDmomzK7WmY4kOZdlXhqdOJEPWKnFd6CFdVH7bjC+4LO
6jOTIrZurzcpPrWMRtQV575W2QjBWdd/dfIYvBDdZ4xSGhyQi2MqfTXa/5VnttuT
oFj1ryp9ik3eLxCwtv3BM1CMYnhK51zEWN7XWua+FIy38cMUmBRm/C7QME+icQ+8
Ma4UZp3HSYvuXy5anM3AQSWxI68yE9dag3MQ8IWFdwZEj50GN2x7j9qr+5pydRxv
3s0BSAknzqvXukXS+hMYPJeQFi765G3mfm864ZX2/F31Q5ne26ZpRxyGLo2cLKvC
e6/PlTPfEI2u8+HRbsKDVs9JPScaUQVq3hZHZnTmpJ8bWOKfLCmWMt+J6xQwnGnd
3vHzUFLYuidSyOwlwqpEv10kmv6R8//vfvuxY7LhnOcYhZLqndJ1W0GdhCyasAoy
RMn/Vdii4dHIgrEDlO1bCQYOwWEk47KCbsN/31p2opMKojbgZrmsTh4aJSHw6FgR
q/ErEkQiEV0OXJ5O07K4YgUdsPSC+5JHf8P87c9tx8LJlV34WX9beGvenxNKkZO1
EF1ZXT3xnrxM5qhe3z8jMU7t8r+Sr43AaxT78c8oxq8XL7GcLwfz9DY2cCnfYzML
HZcdQ2BuXilngagR4s64s/nrPv4NqwuuAo9+yWeIf9elpXDWYDDyKh8xGoeMU3bY
a+JCn3hwzK6qyImg/4PfQXXG68a4SReJxcGLtcovYJr+3hAqGMIM50Sm8+vQH3jB
Qo74EI9Ve9TOeVR/soqB0eviw0Shg/6lpaRJPQ0gQX9CQ5gh8hsnve5owKR3sL2Q
lC0QXwVj05gKp9FU56fQlawclkxlyCV6efpB/KPHNL1wSsPd8GOhYsgC+DhBPFHF
neb2NMmaT0uL0X3ekO294L/xsNTVrCOq4Kpsdch2MrQgjr3KnTRS5+U13vu/eJ7i
b1ZdBDojktz2ZT330nNukuOo5w+EvZSsxWVIBmQKxIiJV4XCtzxHbjFUU9+CFRAV
VCveMnEqRi7xakanC9cfrGItgUfC+O2BJf5ph2SiEH4F4C+BMQ8fdTIzQhU4zVS2
SR4kWLt487JYGJVYDTUwrBjsFlHB/qyCdy5N5lXwEbtNAWs0JBxIjCOOSDD3DmgZ
xfGUop2aXq5MMEs3TeYTe6nQO4eQKqJY5Yx6c2TtzgK5CGoxjAdH+hCA3klvYvL8
2YUwEmESQlf+xLTQedddTmkpbs1c1IdsxO6WLozHvdN5FQ+aFoDq/UNgIsyuEyYJ
s2H1VS0N7EL224AQQB1EKg==
`protect END_PROTECTED
