`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHM45UrKYa8j+nxpl3ICS6iXQgsuiGADFaTnqjlLs39VNAe9rA5h6iIMCOOcjTmH
M0IrhOHjl6LUW0U9ANCp8s0ytqR3WizgSp1s83kEEyKvpRREGz3dIJrnmFJu1G3j
6omZikZ6yFx5gLnJF9hWUysEnBosJEum+6BVYUG9HqjxBPZRsZn7D1HSJiRZNCBR
rzgf7dndzZxMkDZMGUlGckKhFSWJh11xaZR/0+ZCBYso1HPnTCWdWfYdhI9V2dSu
zTA8B/qda6XPJttdGeTXqadXUVs3iQbkqvgSfMDL9tOoXLJ0lVZfYZPSwoseulkE
w3cBoV5EQSN+ROHYpluIhF2KB9yqOrTBcQLPwveFg1OV9v3e6dVDGgv8ur1qT6pm
oWV18OdOPFfoXQTfddEbC4T/YE9FdBclvzZvcfDrUIV99aBzndsaepwFCp5BfGvM
lW3LoD4M4lBSQCMGr860CYb/mYs8g5GwE4wXx8SNHMcxTTRr1DkxXS5u4suLNUYs
tUmgJhjVeRBN4si8rVjvrYbKPhBX+AdmGOJhS6WATyV6iTLrHQEiCVR8Z4Fj3fFA
AvSECHZwyI+mDwBTlulYqlPYJxy2CwKEmjH4cp4ULKV93AP68C8f/0pOBBKELjGr
W/Msizk8dkQtot2mzSFJhQvT8kAuz6m+8Y4IfFmuym7MyzsI20Q3GjMpb+mFCApd
C4Mnfre6XJpTB2S5b2w8K/wy/3u+SwyQ3hGCW7IX60HCBeyTbf0rlm04+OXATQON
CVxNnBobxiEaRfQEHZEWww==
`protect END_PROTECTED
