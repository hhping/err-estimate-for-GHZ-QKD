`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXZTIOnPlacI0HyPZ7Tcto9vZ4TxBNxNxe8SEpb57GCEKEZXOcEeBeGH6OO9JaUX
IU41H7OmNt2AdA9lDCGHBd0pBsWqTRjBYFRF+Akkig75NfiiKzSupfNvt8Xv6+Iw
ehCnFv7KkCCYdAlsKrixzWKDxK0KRjZm/c1l/Wg9fZ8C1HZqJRjirzcM/yu/QsA4
icpmCMFx2Q9jhOizQT8bKXO0IH7k0VSiJ5L/u466eJl8dcaSfeREZR8j8e9/pCHK
zAwcdutSv8lQChoTJHWQfe83c2LsxMjard8M82gOBoGBOeGRdOlnSqS6vKuY3m4t
eossjvNy/vNxIWhhoG1CX9a54PZz0gwdmHEN/RpLRJI=
`protect END_PROTECTED
