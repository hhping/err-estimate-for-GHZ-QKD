`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1dEgY91NSN/ZPdUg9Znvi3Wt1ytHdyPKEZU4H6SsbhtXtwFMqCzSPfJmZ4fA/Z6
aPOzob3apBeSYKjWMuKdXglVgugB44F/XmIn71jvByaXkZUzDAjqQ84sH+SM38kY
eBWoeZuVGQv1MBwQkolfgmEJqldep1X1YF94UGlEFiGYQwJzto60OCgv8O1UPAZm
G5XE0Tkd2ZNmACfOvo5OBSn6oEoHT/vIzs3a2g53SBLoXmEV8bv0V724SDZTUGaT
q79UD0Fh4SL1yWCnH/+m9sc93/4P9UAZc806Oyue+rEllCiXsZqDQNTdl+9aLvEM
kmbQp4eL0asUO7Jp0vQ3Tq50Ka1CwJk53zcClnUC866GuTuRQXA1KjTM9polLvlH
IHalic/GGp704ZKE6G6SLiVvoE0/NAwPpb4imJetNYSc+vGEINUZsr0KS0SAJFIL
LD3vmaJtmLBFkWhgiKy9kSQbS5iiV4UMOmvCHAfTKviCjpYbckGBi0kTA5sAPC5Q
RSb6lQMjiNKe+vQ3uuKlbRpxXCYGqNDMT5m/a9zPV/xMZ/3gslhMJMphwhZVwimk
w7CAHfddWAdMMRBm4g4fLCPRdcM5B7PjOkR1xxJwG2M66JSzzxs9JjcY5deBv3jP
`protect END_PROTECTED
