`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vf3Cad/icg338oVKcZ+AfG1N/PHPToFduht9nEQg7X37jMDKnnZIJTxsHZv2sJq3
Khl2b6j0vv8Qo7C9gm/Jvqaihs9z/ACFnIVTIc2Hcn0XBN2jx0sISmYpKeUHqBZb
d/4k7Dykp/Bk85x+5QEpGqYzVBfygF15EOuvnu/45+IuAz3CB7X1cJi4P7C7EBX+
8RYQ2Nhrr7MXiFVh4qTX5uANYQLiHaz6hePJzb9vJoAAumq63eZztROXf0RhGeIi
thpoh/AYjtpQO086sY3jIJjNQy1NFdUt5Wk/Vnf7DVcis2vgsU5Lb4x2p+K6YxrX
mSxQi1fTYtf/fv42i2ADaEubAkZoVtWNe3Ew5AOf9gzhToh5GSMX8rcolmv2jRAC
LRVJyiE0KWvtNxNrpzBRIeR4sSa4YodKJdfdDG0T5xOZ5/+qiExkZZcMRwuxC/Pf
lIsGMcmEd5P7tv78qxDtBCgosaSesZE6YmnP/oS9pGreL3H1yc6BDqJKQYyy7Cjo
SMUTLSjpgx2e6aKSr0YIk7zdzomKTnH5s8vXq85ffM9cezUUyV4PCv1dbU6pUa73
DDDjIncgqrJliF5lMTGqXVUP5/dSShOqh65N5XZsTxYbRVPIsAtNrHIvi/OCO6XN
8jPUHtHqoBEd1aC3mFQ/dlPxOa227jLs2uxuy/s5wrtOuxYAZi43aE0wBqfaY0R6
I6g1GPcf/JqWkJQQUVjfHXlL9J4Xlyiu9Yp/AaBcDeSU7Z7+7DyAX/81i1kUCvgB
grrOOpn+QCuio2xwVYB1t1tfS96JX8l/lG+qvh5WQ5s3+UKumxaaCRmncLRbAVrs
hdGzDSf87Ca8cVKalkQ4L7X5AANu3hQ5L9wSD2EMzJpZ+s1EH1yNQP2/ZM0tIUFD
8zAbii4t3yRhllu60UfRUM1NH2WbfuVgp+lrC325tWaak7GVJSDmRG2gkcyE915i
m8adVH5wGTs4vKM+plId6GHbh3fGMMrwImcURtni8ydhDJOf7kaBdvmvVeN1Os1y
ihpMs8/En9jq4foOtC/pzzVVn2DvJ+ekYzby5O5FeN981pbUzHHvLkA9zD2OlcqW
NONSzinvOXOJSlJQZAuIqn8O9EJB5GdP4pT/gCYUEF4Z3C0gKmW5Vv3BG89C4bUv
+lvCOXY4kYCZ0/bant0lnXNODZk6VoeZQRu1cY6SS2nc0KFoVrGhUz5gf/R0k24S
4dJEHDPQnWPzamhkZQDkqzOOkG3GB1shSdw5RgXUxY2qZDfgg+GOJ7zf2/HDUm45
NDOmHIYwBFT44IszcdEeTk3qCMs25K/i6cqm+r1L4R8bUkNNExkB7I2JGSlLDDT3
oX0+Ec2t3O2Y/i1Yvlu2KmAGniDcUXwL86erq2dcuF6/66fRXQgRrk3yOk7t14Bs
`protect END_PROTECTED
