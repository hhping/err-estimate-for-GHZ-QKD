`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
omve9y2lfGGtKz4dNNP7tfpPQfawhpCYoGNs+v9zKPvVwA7kJ5kPPO1x73u9VPLo
/8PfWA3igtoySzfqk7g9xSTQZ/Lsdabea5tvstBpSUkFFz+FCZj9CiWAcYqP2Onj
ZKUYUTiUW6YJcB9lz7mtJiOEoVTvl1uVaglGBHW8HSvtsdLociumIfCZugTClRqG
szw1PcQJhxgJBKb7w2vB4nkD1INfB1kPKftkx1g//D13IplQN0tVR6dkUr+trmEx
EKifTjh7WNJuQoyg2juyf/MJvUc4QcLw3vt2KG4NIZXmp2JmGRrgFxZo5sEOa2rh
WMD/mL8KhiEnlVsEghEAmyvpGKs1ZPmxlRw6HPdS/77EHyJtcPKrtWgKDCyFGAlG
433IVgq1OwTzIOlUTkTSxIl07pNMQoKggchG90FUpXrBAkRcd7LdsY5H8SsKwPHK
grsKizrv15cNv0vbJ0gVLnnejioWpBYYb/7kMx8h0aEsbIw+F/7rpJ00kP2TIkMT
w26/6aw1Hn98RcO1KBOFuCgQ1vt1yFPJWsvnEiG40317zeZ0cMFvbFgYjApY/nTZ
58ycdEKs6bBpLhh/fjieTaRdPnjZr8USNFBJl7T0cnlBNhThbQ6kqX9sL8m2+8pO
wCN4ol3opwTUxsqto1CcsEHx76xxwfaGjVs4El+/8BWmdjM1s8qVN7xQK7B4CILe
kvk3rC4+uC8qh1faDegpzVpCkWEjTImd8tw9HPRdlOVt2eg+H33nlXiwyW/Zp2OV
I5aSQbCK7VaPv82rMMpTae+2suPGvMVS/0aUIVRbLMYkv4gf55fSd+wzCCwhnPWg
uyzmXUShivrhyM3Ea/g8+LVc8sk/etKCRNterD6EL71hHeNH1cmizymsa/GRCxhY
74JaO7QlivltHbqoHMeTUXUKUF3jnXFYqGuc18fls2K9B+ibsRzctMRWD9S8MZ1T
sUyBYC1w+iUqmOZGHcTSfsrjB5sZjRlIos2h0rONnXg1nrYva9MdjcWe1Bqh0gYB
o1c4i/kClweEY3LvvKFklDUz4xBe+8ijm++dcaqt3Rxd52dlpoEi0aL2aQAEe5yu
e7OQ+mdT/AwYrrQ/JRUqfpjHYOucwteBa96RIM4k/aW45WdSTXfpueqlZuuw3x7u
/BMP5cSbx7Evnt0E+63XzcC2bKAkMN7Zk+Kbt5c/VZUihtIEM63E95PPMbmRlUTz
bv92puKYtVAgx8XclKTGgb/P7vAhT3pCeSFy80UheNec9ILPSuonA437O8F0+fMA
uRrdeWp2RDZhh/BTE+iPdh+KUJTg2JfH2U5B4pHd9FH77JXbQlyei5K57Bd9ZKM8
NKRyzxPsfYHtKUfMwvQWEQSnJGj4Vk+IzUKmHHugeR4pSNghnLFpXjLsjdlx08eg
HphLf17QbZjqKgNpR6cas8lGZhdyU6VsM1QLBWNRNq/2xbUDkm1BofArHnalImtg
pylyelkpcSZjIZKVniK68V5CA8twj8A/Gyve5LWSZaIJrkTCA8Ivk9LB1kIt/U/w
RFW758WqOs8C5/vjfTn5lRbN/yMb2dj/jjDn0CFpcy7F5lnGTs5cwASSZzJ8AqP3
IhanhiHic+0CJ734DSxrLhbfIKuEmnYXsQvYnajPHEc92qUukfykj1yc/PtNwcYq
oq6Rn+f8UOJawQMZDDBqJjUov4mwiEScofgLymKMZ4YYwmFo9NZnB/s5bJmEOdQa
7A+tk7EGDmSnOel4aFS2IoVINUAo6wfsFSWSogWhNWAE5afQDo4VyBCNe9UvlXdh
efRGu/V/nlFCtEBt2bnQsse4CxT3YdQsuj2pUA4LNNbORrryGJEhfn9c3MFBvBpu
OujZG7B8G2SF2ErYCs9oLbpzM8SsiNUqH6JEDD3FnimXwFHIZqSUcPci1rC0atO6
6D2k4nw3pcV1yOj73axQXeLh+7dqnRAZQjeaiMCySjIkOMOhYJsYBcrnYc3uEhKo
MbDWR84/x5ezVbHVUbLNF9OfLBDX7hXCo3StveEGA5HpTIBfaKdBkJRV9H2IYHHf
JNi8r06yP8YMD+JktMtksauLIqgNc6s26gNxq6FR3bIOoC+/65aCWkLRMB2tbBYZ
d0/8bBN0S0SFkM0WkS4ApT9XJ8KRoEXIH7v1xrEwMGZ6AQV4o+llVirFAABLM45I
6fKZ9i+6aMummnAJjhg6ZJfJIWGMzeSAaR0OSjxqMEfybOlNFIWL4ZUzUYD1HF+a
JX6gfwkoz+yGKD7sUcMr8TMkT63k+aYl1zsegEZ0DRWTSaUU5fNDoNLAUn4FiMUs
f3KizRvEuN2Yg7ltPQkdlHHfn8o3eyIdje5rjiKuUz0OOBb/WVd3nKR/IRYpTOBh
VtL2okDf2w4f50x6yHik3zqMN3N4f6OblYV7t2JQwl4WxSidsOaeTm/keSO8PcxW
kKA3DZjcVxL9DpJ/YJAegKlf3iqNbOPyR6y6/cvqKc44tkvAEljf+lwHaofX9L+B
ISCMHpi4sjsCQTvL2QLHVJY6eScESlvl63/Mfhudln+oZONBnlzdm3lkZ2Ve8hmn
F8tTzSbSquYJzWjY+m87CdCGCw5X/gJbIiOMOkdYojWf8h57F3WAbPlHes+ROgRm
oxUlkCf0QpApiUbRbRDiqizi9jTvdpSG91Hqh4naekzI15CY2NmhXorSKtBt63Kz
2qXONQix1JzZoxIEJXlIZuxG7odwTgBVUxBxSdui8PJMukT562V2/kA/hfDydgg6
/at73dWlQCxQvS6YnyRmFNx0U09DxheDjKBpHCeb+hlR8ssIH8zVwD/Gs8WCIMAh
F+jcDOMotgt1JXzBhtJOH0CqgrrHQnZxfEa6dFYA39/CAFi1RqcshYPa7UUoBQou
QCgAAt9BWr/i+HionOmQ2qtJ8Jl3cBClCLg0XBpxBK8KOXUH1/HVU1MMh2TDalPz
JL4LM51DKnrX6cEoxPTyNahgybuRsi2cyKrf0QiIK1+0OZZ0WVZ6bkUY7+EHgKLv
nebKTWR4LSF7kxRLp6Rgs+M/ipvbyCsNAwiAwi/6MHjiWYjntHb455fOeG3i4CKx
uuslIpm11JTxHchWWJZx1sLPayTwFQj0efBTioN0mRJestiRg8tlwqU6i3PfXUUu
rxxtY51FzZxb0opVNhGCH+dz+bMIn7q/QBQfYx3sNjKwK/pkIs4i5HgSyKPJCO9D
oTDUv3MVWCwfdyzmSWjUtIxDHgDaoS9ArYoNo+NXxWn2h8P0nM2IK+G4EWP4h8hD
jhAAj/erm/kynv+Z4qoubbYG9FWfWK3YWO8h0BkVRjjIDyIdCJ7VPS/gEasDU67o
mOldWL8b98Oh9tZ/FuWd3hjBdgG1ryrIXhFP8naugr07nasOSUSqpSkaMLpQO4rE
vuYE8/hcULcWwV+ZOHXAVligDMs+k2dmgYLniYQpFqqHswGyhgM0XxkPLg5fCQWL
zcqBxZGHIksMVs/HkYFvXKlDMHF37UrcM9g0xcxaR1BuX9AFg+OxJBV90zxFNL31
X3xtdrELE4nSV9hMGL87F790awEErFgCr4v3SQ7Ec65yUl+h+aE2vPxSJvJSBeZP
5/HdJNRZZeoz+QMU5REKWacuHhPEQa2CKROIfGRCCbINDDJd1A7oQPTwDNEHtcsE
JQmbNzSl0q2S7XSaEaOyYvIj15tWtyMGsahq1sFzRGl1WE2zfelYYZESyRtjp0g9
hIo6SKmvGkEmMz2Zma7h6zcDfYWzslp8Fag5PPVu5F9M0Qf8H88X5EgBuj5PjVFW
F8i2t02cYYH5CaqJSfppAym4nb+ZkzFxOaiLCsSULrjt9z39Itrg4kTBV7nctgSV
jRysHo1FJ7TMcr9W8+fgE1VEHBw/WP6PwtXczz+dDkEQPAcLncC8K2JpjCihaZh/
EwI5R6z0h3YLzriY5/WB1zZ2YTkDgOmATMKu1mnop7Wvh25qcqjOmlPR0UDs+ev9
29ykH5r/N1t96F5gNRQDqVKTxJfnFf8RD1+Cse0VnR9iOjYJQmYYw6Ngbn/1KvnV
5rm7ci75xXCbPH2C0dKpfNHrlWJqiOJYyvyxwkS6oCppVM5/HeZcE10nLOKi2GLm
fL2/kO2hMVJznp2o7+egkmkqUHoiZKz2LjfXbiFpV1CrlRs5wmddeFs1kSuYrPHB
B+EZDRLkEXFyFmvUH8MayQhQeSZd5aH/bvcvLCvWJWnPTyZDSrP244zwtKKseeHf
YqvOwfuht3WetR7Zb/Z860iJdqffuaOb6mfpen584zjdPTdsSH2kfffEsjE03KWo
hifRKcJn150cwDX/4DstvY4D2c8dWrq8XU7qs1vqOF0RjfGU/cPXdlgax5EAxRT7
7QOhWib9nV51sfIVnr/J8RMBVoivpfPz8bXJjW+7eSwTNilv8Jf+xHDwEJ/J+h6a
MzK2X70jso2ZCgS55DXRyCT/6+uxC/o/ei2QDTJsOWIz1D4p8ctddVUN12vrXdQ/
8/gtbE02Iz/bGthLzFTdoUx+vkJvGLGL+NIxyxAOnh8NGOfv8kUQSxn5LxeB9fkc
/rQ/0essNWFzoa1gHc6FVhjEQv22FYtlgRuijk+ILYAvHrRCzw5QF9TRbhsL7VMz
S2ykUryTzI0j4xYkPUMNfdLIFCVVVplWwQtJmUU+CFgjMKzwXJnRS0Jof16/wKHl
KLrofk5RYONG8CovjruZTiksg3FUvT09/Vd5hbCKa9PnXXlumG8CrksM5hHNYrnG
1iusrIPMwRyo+3tg9MLFHZ4EYCY7U5ayiyevEMCb75iZ+uFdwEfFEp+MBn9iAYM4
mMAWNANY0MWCZWy6HIGZXEfWOhnim0IPgg0xVMOpyzxOO8lAHs+mA1O8Jdm1aE3U
1p56IpKwevdKd95IDiQM031hBYt4dc7Is+blCoWvjSvT8Kyy05/iW4maSsCiBXyy
Z/VqS9naS3HNO5Bgz0GM+t6lBD/l5sGY9XRULpwrcjJsb6ePAUav1ERhjJdqVE2K
emx3J1Ko5XC7eA7CWhuI3V2HX1EYxovvasXutEBRq8Vj9yDV4ySs+sQK322O7pKC
GRyxPyEqLgHbREn4LOME+yBb8nOOzxajo+rSbq2239lDUJnUgWwzcrjLqE1MOOYw
pis8f4Bi9TLd5uJ4FKSmqSqnCE34X5IEB+N77mLmQOG9HVlo5aLEveiFSg8tgnSL
vYwUPMWt5shT9QU0eZuetKBfBEjeVtGiKltZgdAKsqEE8scK9pE1DEX7ODEScElk
kU41MLUpX2y2y75bNjCf+7uiCfUymlQapJCu2czZLIm+WzzhKwMb77nSZe1jvv5c
Ux4jlXjM0Bl4NDaHH2l04GXn9ZaWbN73Q424phG7/9+DsVg2SFRkn/9jsK0Vune2
ux7Xm9JcE9w12EXqG0z0Ct9CW8ivmcG8EGgZy2mYSTF8axdKjZL9jIsAQ+CHriR6
NaqH153/XJYrSX1yZ6q57bCd8Wxrw4VPBSZpQnxtZS9tcMtT307i8IwpU70khujs
rybFb4G9PawuAUyC5GvQqDEJdTChukI+nmyVAVPfxgv/Z3CQE37KgjDT+hmb1U3I
JO1s8QZ79q0e+6/NOG0Bc1XmaRJTHnfUq1CpyhuWPUayHYv3g/RbYuoNYFZUIEby
ioAVnYDnqtY5vE06A1sLV9klW7skFj63jIIQLodhYjdBvqhSPZ56FVa49rjtjUBM
R59mJahFFzB3I7saQza23wbltHnX2QtC518oa92oTk77xuWP1RBvoElpc+eM51VU
gON55jdCS8WAVIebXzASP3nVzN/bSASuCj2I+r4/Dy5bGxd0VNJFX4eZvs4mtJ8f
TZiizHMFMVbjiAG7QmqUAJ76wS0U4gLQTmjFKJ9G96agxam4bkFZfoaRoEf4HkWB
4iCcHYOH2A08pUxvRr/plLru8yh+bFtDSwNPUjQlnmWSN5JjwVslCfyA9oTFTfM8
HkYJU2SXQb6PW/c5qVCRWO8qi06QtBr7SaVr5lWFgIpinr21aBLPH4lecCIC58Sp
7F8eP5JgO91HAIZoQj1elem1YGBRbozzodsQShdZwKKl92IcmigywCNeo3MOOn9V
U150xMkdfJWydgD1qNsPgPWlZWtlPyml7rVI8aOs4zhLbd5GKLEcR1XDGKHUM4zy
k5/GR6poa5uqnNtx9duKz7ruEwDkLyJ9VL3gJNtF0HZvUErzhsn1+khrbN0UdlRh
FK/AcDJN48T8MX7zxzj1tyhZQ+WoW+28w9jyZEEA+Eb1llHKkFGIo8KQXVsNACdN
RQU3yU8ogY7FjGcdHcGJSSlliaGOLT8i46xC4lriqwrOFFLMbPg9CNVY/Mt56Wcz
3gZEPtwmo066QYTnWChitxgSrxu53EYrOccbgWmLTBxX/YEzzqtI5X5WoLaDGjir
skcRw3VNl1lzH13tRIXp4tzrgDVUXqhGJprkkFYM+PbZeUblozTjYdQ3r20oS9kV
NTXPAF5OPll+9GDHnuAto3FjEwu+RkYRuVir1WK23alag4sgSNoqBfdH+zKTQfPe
69UwD2Dt2nGAdgZ5j/r4JuYnfm29n6miUvzGpotJfqwy/qsx/RlOuIdAu9MsUQJM
T2PvNf5144KsxEU+pTvVw12vCrRa3aaplVt1AkvoCLVwXD+BNu7stD0JXQG8DMHX
ZtBEnhZAfItmFX8QBCBgeOVLgmNm+jM3PjOaw2A8Bq+lfIRO4cTtI866RQqRXYs8
jU9jzBHzGiLZABHGKyQtqLYr9M8WqBg5Mvd/6BLz9xKSoA37FEnr3mkSMVqj8Azc
LXM2ooZKgoPmofnxYGNbiEBAzkRQyipXYsIpoIMtBw6AgGqmgOzLpq5aV6lT2nkO
czpKGKcsrhbEPbkyspFqWc8Lvp5uWbcaMUPTGQEYW8giQfx87+7A3XJDlLjRnBsI
k8TKbWDap47Zze4tg4SNlID7NR3iyMKS/69Pb0en2dU8oEWpiMTYLLzuX+qIUJir
spJbaqg0tFeteBnDfwUo3DKg3GUPH6hZOxHvKDv/lmbOZWAzxQ1Ac4wVCiDNFoKn
hZ41XshsGm/zCKR8Qa/sqOEcHOzpuj3o/hiJYUHsh8AG5au8+MqK8QZX1eHWjKYR
cfPyLj174I9Eu1iRoUAd1uIG9Sap5rWaGKsGfoLW5RLHTeTV7NoTJJSRgc7JqFyd
W6ZsUE2xHNSO2J13NTT+0orJxCsZf3C7SWH2A1+FLqCFMErKhNVMhc/ng74pXZPf
dBmukAmd2fnrYr7t/PdulDr9x0dkCCK5BNZJUy6gAlPCkrJBahYZBqCd+IhZgeTm
dsr4cOwbFHMhTzAVDQjALm8tUoEy1vfAqTHQrC4EASRAQKsXAf//KVylZieeKpQL
KKPDo9r0Y1PVPVOQ/WRzk5GRUtVSGOTuU/u2vJKrJt+CEehnczm5j1CaElqUtf6R
4D9smwfK8YXgbfZoI67ajJv+a5siXYhqfzDf5GZjDnKa3QVP/BX/llWo95M6IqKV
ek1MsncyJhqpab09031lR+9oWyaR23KIPsh7i5L6SHPpJinZ7RWZUQjF4+SBYTdG
krNrNSoeOXHbFzIWlnSoRXKBn9ORJPhHaXbs7NSigr7NYN3JZ1b1j8zUepWOfSdz
m0E12+cPY4fpdF+8nEMrSPY23/8t3j2qPANxq0WMrSeHmtA0K5rszsAsF9YXaQh2
l+zkGZAnGcifchJg41iVp9RHqssCl1bjakFVnXXaaBxpZ1k6xqzrjCGNyiewgw9q
scVBQGy8ewjZmbsrZ5rRl1bIDsUuI6nRztxAAwMkS9T+WqH4lM29tDGjDB/MguXX
yWghQ0QOCKkyLVQ6+S3nXWj1cPtOtaP9uh4GDeP/VAUPPwDlF2xB0WROrBhm27yQ
FKX1bHIOudVmLw/1qwZd6KOIhiKlW6b8X/bIVi7GJOmLRYstWZXdPRIdm8lN/hkh
CeWqF19D3yezT1jiujW4Uf1ZOT/eLs1UAKLWdAFZjEvDDAHothMCMjEqU7rLxcq4
0WYCANLvoPiKDkmsglLLlhUG9+HChpVHkWCCiDoSw8G4swext+K4yrHOYSB8RtSB
GYlqu+w/wWsgXSAFCZscfBmLphf6Qjo7EPIxbGsLRMZ+EDDcscL046OybtwVd5uU
sSM2x8OMkKQGzEgyvzweNNN+946Ub7fENS0dlel5ARH7/jENkaw+wEP9YGyBLGrv
Wj0VcMeDvKqfxagRwgblYnpbfEH+bMRhmriTNhDBptE32Z/C6+OuFx8jVz4JAMfb
8JVi2KJuzWNqW2v8dX7WE2pqzM5xoGTcf5Ayl4+/Xs6kYiU6MeY/+jrVKdQPtrxq
K0JAP8mahW7vLluKZZ/A+b4qq97f8bc4wJ5duERPu7kJjNYsHGWJJV1caVDPnYE2
ofkIdLsfEtGYAdQ+2J2aiChGbowCoBONXuzkRMhn+VPyzXNvg+4pE5yU3/iFORqc
CngpRVvULFrY5JYkXTJLuvOXDU8gbbLKT5s1tUbLDiyJyOsp6NCPrkLcaL0kJRbS
yo7Codid7ZOSO/cbq4jVFfDIqP+FopvsRgnGykPYj/UhFWwAL1MdEiyRekjKHfuu
gQ2FDqyz4QdvIv6eJSq3pNVreBZpKufDZPe4Ybvx1Dm9uplklzE3+ucUNqgui7lr
qJsmDjgWQSFzIqifDinyqP3WR8mKNvWrDJz01vQKORedro9WrRBo3z0NWSdupziE
VGftnaF5wzc2ah2MWinoZYl9w/THa9EBOiYsaPUUiZJK/jVkJl8NTTsgTgRzTmLp
yi0kgYO0jHVnkKGsvIE0HgMhdluSdiEOmxKNvKi9F7qjiCnpvKFjgx+zoddwgfqq
x2RE/B1yh/5ykuewTmmabmJoxh6rq+s3poU/9jxZK8STCMpZpNvFYTqAnJtfidYp
SZD6xeaCoRWf2Boul0ofRjlogR2IJv1ooYaBLTMyUQuY0LwoxWe2zgLyRJsYSib1
0BQKf7xmG/syyCsa+hw6IiS1oITR9sJ+sgieIgec2LS6LC7mPxnmcWBiMqCquERn
IlujhD0KNzA3w6gcMJMm9GFFJ8P53B8ypn28yyOzS7/jhaORlsMG10xqffUkT4UZ
c9OCMWHf4bLmzeWrXEbiPF3RkifXSE63rHui222tXdqcZzNHFP5LndnXXOU2SBcY
03qPRIIS33SDvHIf2mOQw7LZ7jIrvbFMCDWPQYbWIXaDfwtdJBanJA7ndxislPFv
q64TMEOh8gZpu/i8GmwVymo+v+W7nlWL5++uHva2eutsSEyScq8KhCG0SoP9eHUd
3+veaxhVSYCyVp9pi+hQeHmYKVFU8wmPm0ABNVb9hxfAgGTlu4T4C/6lVKkDtPbK
AQVXgaw14DhWPHSwrokW3BwArSPsmYpX5wKN9rRh2ISRhzggKxd55TgaIRF4sLaX
n0aq7J+u4XeBUkQ4QQaZN1HCnuY0vJwrFUQfhPcVpPP6FLrsrPUlDENQdr7QNEtf
xQBSKT6F1gJtX0J6OFlK1NVs4J7nGxsnk/+J3gtNJeekdrQ6RpNZR/3JjEPI2xoA
QZQcJqNZJ4TWkoMvfO3vpMOwUEIfRzsxg1FYWvIhCK0mxBjw6E8tVvr2aEmNoqmE
uaAgau87RgCUajdeIeA/CXPKFoq4ePJTkYWl7rtPz0ni68KVp1HvNgC7FkLPBajO
nqkq8ljuMvlsSLIfAlbhM0L9NpNU4joxm+E0DvbzrPjK4OhGhTHFPZjMBY7bdIrV
zxCk6GWHR9eKhchYzPVzmmhHQd4H1OCOHhN1CA2wAZkdlNVsHYmXmjwrq/gtDtnx
EY+HvGQJ+prHEFSoq2DkiYDlB5Queh+936h9++/OGKKxaXB23UF0X+s6dgXsgTZ+
0jmL3moo9A3TShs8y/WLRJNFIooqTx5OWKMBfPGJm0zvO7SjhB3xQNV68XBbpBd2
Jtv/t9gLUBYd5TvN1LocTcJJsRsrgf8ALKt0VeiYUccbHaQ869224y4qpB4D/MSU
zuT95Y5JTJyvbP5NS1tDEG/8E7JbSx4NNgHnOVZt4f4fewj2EmlR3NqbJksYsSFt
dsdTcJiuh8uv0p7wYML4jZ5UGXkCV9l70QYhmJWBfDkNBf/gxMG2GqcFpBkmcTna
x3nK32ACkf1yMdATN9vRv5zi8vf7NGNqHL77QVHB9Z2gbJh4pzv2jXNp7d7qHQgE
OWkSXuKlojNJIqbsCYc8AbJ3rbdcEe5DdeqAqeZYsctXbuURko4icnL4WBbhRuB4
4ZO9Qsa0cgaYPb3NL0e602UvqQfY0+4lu8Ucoo02X2amGywV5ossL5qHtwkXca2R
UNgkGbXyhwgHs9ntOPmfIs760zxTIrHmWwlrMhn8fk4JPoCLLiK0lUkX5ggyJz/X
IwO7mzo1aT4WADFtkEI8djxqOzonh4jmWdCz/gGUAU9XK+J4+utcxwXElxThfP85
5jzfi/DcOUr2PnMHAF7SLaqUiSYlxIjaOKKwYLXqdlkBGVLjOf1yM2PPwEGpeKzJ
pDrsLVNCnOQyc0OxGctTq1vPkGr5VzWdng47zilIx+qWPOg/XG3eyINoGgbjCbsX
5oz3kd2DOcZzuHshmq7LRtVQ9vU4RnFY011knno8ZwY9Z+6ZcSEblkI8wZCyT3XK
7f1DqHuFazWnzUcqqGXK5z481Egz58hiZq/xZ1cBHRjBBzLSQDuBuvdROvlvW53j
xjOB27KeWKv5q0h1YVl7Y1zEPIuXALVvQ1aUTvBwHHD1ZjiT1Qqt6ZDnGKBDGKrK
sYG21UobJMaaC9CiKl9QiVu9a3SHvXTXFU9f5UFKNzrjd7VBCCXhUIxsC2G151wv
ISX9D3IoaKtjAe3omc98Qq7/xgle62aFytEOmq8jVj8YyEINPUcFhz6Yf5WORgIv
UIZCgGtAfmzgYgwYiROBkad+36nCiM6kTQYWnIIYbEE5mkxlgryxSu59XTEcLXsx
y2IWORqD7YU5yS7uyLrLh5VrP+AJ6KDH/qRFi6LVOvM4sCYH+L5nuu3RmnW8tnes
UJEG6f0wPoDsWSPpal5po7I89/Hsgd0R3pB4vC0sAsZ4CHr4JpvZFZlLvqVUQzNY
OZMqZ8cSQSMEeWRDGa0esmQxqS64Wt5g1m+ejiP573vjnMjXhFiVA+Z6zOELDYUV
jc7+b9fjB7afxG4mTpc/mnonJMDHoBoyjOiyPblkmRrhfZm0zyDm3u+nCneIxJjs
Ws9lXzrubltZmYhP5ODQu/eVOKagCn6XH83Ck7WN1Te+MDl8QpBT0tp8nAUY48lK
MJydzf7Qo29jVv4UvWxuqdQX/uRHXYSOvXvbMXMJ8HuOrXXeZvBKUfplENauP5CS
kzWvEk7dH/uz45YZcpq4Nc5a+djfYhsksclRs604E4+2h/v10EX3RQ+kMCqhh+Us
Hkniam0RhSN9ESanMWRy6zEBC1peEeC7MiRGs1Rbo1JZGfi4uIrbJG7UInSTzDVS
IyZmvxwycB9oy+K3iFawVMTwlETD+jMvWA5O+BgvjBUIOyYWEp80UsGC9q4zH0BC
zyVnUFsNsS0Nzj6G2aLIkkDAfxcLWxAdtfs+Iw0fxOgT2HirRAIk9/Oe1rg8UOGm
SqRlV4KUM5Q5SnSi1Y7GOm0YlWzje1qZW14gGT8VqhlxSsKLwXLsIGU2hUAKRkHl
bLJfy+dTYi0R/qDyvqMV1AmrX2OlupcJo9vjAu07S9IaJd8K93d724R9yK2L1zri
sA/QuGzvCKDNWaKYog/e3/HTp6Mr9pRnHlEtZT+p4urfECSEN2Gt8gPe0UQGA1Ys
pn6jABF4ORv+AXNieBSvJ9pWVyLaKjU+T/VP/ECk0GjG88Wr4vZbOwSg/2CTD9ND
oDiETjeuCtMLOBrX0NK4n6OOer5dPf/mnskVXwx4E3LEWsXASWKqAJ8E11pe/YiB
t7Osa7F1lGeFiduWlWgLrRhlMYhV00hE5Oq96z0giUAX9zMrGkyVF34zgnRM3n0/
tlIZ91IUuXoOYN2stbwfOau0Wf3Lzo2HXYSjaUPWPbfToINUJ9U48Y5LuRA4HckA
7BWVclZKJpYmMTWJrTVU5EXH1EL0E73YSFiGtVxEFsjwmmPXs6IFoh643rHBr/Hj
SGAjWQ5pDZyWOI22f/tmhaGzur5nkaFOaocQzEkzOLzHXmgfs/gE3izXuH2skbUz
dTb5lwu9tv4WO9Mbbd1yYwdVMTFT1K+rrq+ajJ2NWt/+bn0ZIaICkWWlepgAjR4y
pB2l09dzOlCM/USvW0iB1YPb7MsGQhDsvwqcJbnE6QRVqLz9aIVtNsiGqOZHfhNK
milxnEJ32NT37uBT2WEo7lS6aFA/j4O/YqLnIME+yHV3hjwWW6M1tQztEZAEQq7a
LJ0TCQR2JQ1NGy8EVULJpNuEVU+252k3pCdIF6C3MuStA9fhSEEohsjT+Sn77gWN
5WttNwfXp2JDFWCJdaqna2QsDsNQEjwi4JNZLUf5rGsCl98vx7uOftlVHAR6Y8uX
HheTzurwNbKbu663C/fEpUPBUCZpZfYDjEsc6hD2J1bhCwDLDA76C+KSxe73wqmd
TLFk8EQRYz7sU51howK3inEgetnQB3sXgPSrsG60g7yZ+fYeVQybDBf/F3IuLL7F
OFvOaiormEhTJWDtj17vId8vB841nSgbFhw2wa0jJ3Ck61zZkzdSNXVsqXtZ7TF+
moWLC8DkhNCY8o5O0XWaLrnHRxh3dwDpqLVlx1rd0MrUKlQcPTBMI9C/x7ZeENvS
bCEi/id34LGu7mQBZ4bLTlni1wYb1+/OKW7XaWT3hE2gKpzY6o1ep5HJJvlSE3X5
CBKo1rXF9nn2A+PDb6BaP1BOEW4rLf/DuzFUQis1ToeASDRBwwWjBk/c+E/CJ4Rn
3HvGJ+HOb3pZNf6HYDdy20WNW+lv1pxik/d7+C49GyAGaJXqpP9t83OGE6oZJ0hA
iWDfLdsi6M0dGGygUDgQE2ywEo5xv9glKBv7ppTtisy/ANTq8LrDO4YldRlfmGpS
+RSp5CwDIE28sAkE9scWR58N9N6LQZjAjJJgl+0yrnoALFU/nNvYyo2dpjpamhbk
ux0lgYm+ZjvNWo3lqKp61ZoVPtpkfZcUvhSDhO2Jn+hcwJqKr1XJirtju3n0YqbE
JE3xPScM9Q13VR/iXGL/e2kWnXi+2BPJgnWGS9Bn+VdcMerYbCeeC9CjCuLERmLM
3jhTfyFD4Gi8uMojV+z3vMgOUkXTCvPB779UB5VkXhErpgwmJcSbgDlGQ0a7MywR
PLAa+mWDdVEtGgvRiywB++E123UaImhYakfRqnDUOKn0VzSCufBqTn4ErM86JYor
Y6KoacZLTZCu/3A+gbI/b7EVzbGXrxMPyY1gS4Q0Z5+7n+n3KqhoK1uzRn9RDT1g
c6Nes1rB1wfUwpSeZQw9T6UrTfa2T27zBLrHN4UyQAKJqMoww1uaecFtPia2R6sF
cNyotuACdS1a1AE3toX+3cm8WC7igxIWGSGioSvRRygGbSHXHcjZ4HC/PqvQqBEj
FJrxEtxKj+FxH27p4hsp7hCk/VugC5SIwGB4SBc8R8BmtI+ImOyY3wMY0Si913Ec
lJJRcv/zfuPyCX7TVDTupPlLQszx5yOIDt9RMesNiBDx2xqDFCuaS4c9eYwSWRVf
UbUfJtM6WQoSXEYkSAZI4mrbtpyRnw+xTO6W/goIKKAqNGG/CT1fGGhlsOT2fQG5
wygHcikLbx6+Nyjm/pMitM6WBHVkLVDw5LgloJEDTR6KpknU3Q9A2b3l+ImBaqQ7
YUxSqg0Rsj8MOJy6Qpi0gtbXuVT3f6RhaCjmI039cnp4oWR8N4iZNtQcHa762nU9
GKdIA75IyHiAPpNfd5GQtm597cNcC/zz+0DhqnftNES8QIXoNifO3xs8bAe2FeHk
293taalqwkdyG8LRgHAmU/kUCLMeXAUQPpdeEJW+lIwEOj8+gED7FCqtVIfZ3jTZ
P0dIE/pgi+dD/NdUnXIu/oiBfcy7AoGn9pSJ7pgDVN5s6UL+DrjDcpAkSLRuvbq0
NIKIoW72AHWdP8lgDoRqRU8F0szxbTGcQBB0v5RDiii+cn+gVbFqY3z1ECZz1Rtf
3rNGB0plPCydZE8YqbYcrkkAT6ejPr13p7gqs6ZBrhqveASsAJ8OxmSrjIhmnG29
Z/z4uR/bD8unc4pyUJ+d90zmAST8bByngiqemfCwvvdt7OkiBDxnikgSIOMlXN8v
esdKdDNRH/5c3kyiiQKgHhTnMtRXpxaaczgmqTFHI1z/VtTuXe6iLqENVe+z1Pr5
LSrnGzxJCYy7frspYk4lSxOCucfLsYQ8vCbJsAucWYZy9ButQkRlSlxgpTZryBsA
sBf507BVONtgdG9GLr/fvAeQtSBrVGghT0T9/5lVYwJbnZT14bob6kOq/xYnwKO2
/hmHQWA6USiROl9jZfFUWDx/9dZHKGBs0/xaR7W2lOemGliT1oJ2Jv2MY7dWyvmM
D8LcQYzQ45RHPa13fEFJMkmx020jm4oMN9+csjMS381C2rTS+NKfokpEGB42pBaV
3xtW1GUzaTSOG+3+nxDhcDZY6urRhXl3zCJ7tG5t2drxHENpJ7ULS4JrOtHmaHtW
rV1IuqDWBsykvvLg8VbXtYfg1y6fyPeplWXoW3EK/MThgVdqy5Kn8HWQyO/2DtLS
gDagP43YMjVjDUBVtNHh4ZOwGUWSuEWRhGQRtWvKl/G0tAbINGmhIIeT1XXBTQ/O
XkOdAH7QFINSPMT3jow5yZTtU2Qv+nI3PwjqqTNU77Cip+mdAq/SVra/hKypOoMG
lSE64X7gGdJa6iVextv73nNjWu/XNTie50/gX1oyGTMQ7b8TklFAkonpBVq7xbf1
Cz1ZLOcM6kwQ/NPG9s2XimODMS6nSFr5mVDzqGnxcNFYaN8lxoMXP14JjuhW1bDq
a2gseItwNJMAhYOxi8/PLyINSgLtIbkZRQidd4SKu0V1JW0jgKOFIJPlz9skS7+H
8nd4IFM7FdlZtrvXh4RQ6pEmYa7AhbYYPgQu8C3t/nOZQw+l711dTbtvK5txwoIB
FsWvAXQFWH1mgZCeNjKSc91v08FkVjBQ0a+4zvYGcbQd2XDz3gRJQkYAX9k48mMM
xdjQAeW+vl4eIC2P31T95rQ/45h/XP/pYoAriTfoxiFS9Lutk1OXEoFhUiZZ0/ci
7iigshLYPOWD8CxhEeQp4KcopFZBTBVnGotjz5EO1MKkgVA8OSbrY5d2KbO13dWY
g+Wm0dTgvbnl3F0JUhH0CvwXlMVzjesfO1EzrlkJtjyDBzOpEqrSx59sQg6lYjJo
gLqUVoP+Ekx7rou9pGG6v1gntCnwaNJtGe67MhJoLV8eIRgyyjqda7Gl6aUpD+fm
lzDN4mk2OH+m3QJ+C8UyNjGHnL61xYNra0wtF7QATqrXXcfxPU60hzJYIFe8UIhS
bJEKuFLhPOsAz8eGOa4OZtdTlnnvkbSRX0kMcJDok4xYkbspd7LdnqKI052Qrub/
l6pNN6Wy38KSkVuXs7+JODflqeFIxv5Avt0hJx5tu30PK/pZNRaecIvSdabquUR1
EzTGeqillqliIzctViqEp6GmRP0ZLcMm0+PyKr1tRP+iLX1iN9BX+R7UdIp8Nbzv
AEf7McO57kys5c/Rnr4GmzyE/PfQxnSwmZYLKJDrYYlEkomGXY5x+jpjhEiaBa+3
8YGlqOJYHkx/qf9a0zDMex58NSsFsL4nlxQf1AQfRdnXnhdNjMdF9QO+kKhzaLUV
/tMvUFvyl6XIM3TX02XXDuEAeYKPKiIZGWCR8yWvDIdgUggGVEMpsDsqJfgfXn6W
TeannRch+CxJIzQvpJPSsCnH7ilBQoDNsz/U1jwIll1rp0JL37Ms5h0Tmr4lw40I
hQK6kkRag8GsSM39wyRGE+xaoGhrd5R2eYeVCDXJK5yGBx0ipP9B8/DKCiCmlNxK
2BIuhORWMSHtVC3gPoWr2LJQkXU/AEJSoBFGj9M94ej6NE5MLXHUCm9sU3ZppYql
1nWltIrFZvxoLuLqR4oyjHzchGyifSnPP/Ya81cPgpZfqe8S8OwyYzJ/ijwRkdRe
bAeWPdeYqfws3SjiNqC+3Y9sx+bCMn9s+UZUZSJt8Q2FoTP4XmLRLduVLW4MfOn9
rX/SDwWarPXQDpF/20O92q+uqcfOS/wKdIi9R4onFWxcoATXEVlJGZH9H4VjlxMw
ZGy1ycfze4PnhrBdaKl7VH7MYxJ6DaZnBubfX9OtovTI1aQirjaBMBcW+jONuIZX
dmi1K2gGUMdrx5bzIh48JL/SbqzvEwqSS4v3bb6fRq3kJzVIYg+vPyuzOm3JGXNr
AEDAgScITesW+QoqQLrXS6u+tXMLKly3KubuUOAQCbHtpDrutaTw9OhrSWpwKsVv
4Yj8VFqopRD+KOyog7voYbjDARc4aM4vmM9/t5uf6IlFRcbSwvMGPIhnLu00Uzqm
INv+lsVdp0tMrH8IwP+YlSIETN2tAh7a9ojw3kEuD4VplyRIC01erScQX1B0sraL
35m4zBIemCT5FhY/z7Y//o9aM9KR0JYXTU16tRVjbd6Iztt913pgU7+qitmoQ/7f
rGmECR74HvmRnDpaf8pT/b3Kxxlx50w5Ff013PVx5Lpj7M1zWKeWsGSAk3s2qC5K
MgkH+ZhJKibTNSpdd9ohsLtVgIb9oDPqbyJqx6jeuHokTOPqtbTSpquk+4hNmXqa
n5IXXPa1p/BLwg87ULY41GKu6LCk3vGr1aeisRL2S2ot9EtPk/1vDwj/VG/981qS
2mx1p7xmOE9YBAQE4nHuLXaLr5kOvKOHfRTige44DUoCVtCBWQ5nQDvJo2xbKdt+
2oRzq/ORL2kwYrInLkJS0fPPY1iGMlK6wJvLDfIm2OZ9oy7vpR509pyYefHxsMUp
k1krrMxCUEd3K7UjGUEcvJL83Xgj+LINAmxCPwhvfIT7v+P70TNDd6jBcLvnhog7
8VkYK/JSAFMpNTOkVo6ZbtXlmWcFG+ZipewnGfksEldWSlrJ6dcO+/aYJYP/M70C
GjR5hOyZyc+LlRRoIszadJYHwuCU6NkGLjhtYe8WraiZEuF+XWzwo/LekE/tzngl
54Fdf+k4FRrmqydXGiMnyhE4q9F3cnudM6fHFHELehT7InoZUfHwwVGHVLnjCnQC
C397o9kY+cDbxP7FEdSPKCoDuzatLtINKWFmWb5YWIeKRIyDnUa8iWK8aKUkzgR8
mVX63EDEs9LeR28014+qlYXnLYPAw9SmRhg5WfYbbCs+jUC4JTDvXhSLHb/+B+8G
cZfXTPAMCQa6cepMzG3a1N21bc2Fld7sowWfKbUPGTEaz4cWMp3djB6ek23JlGnD
2HB7Jsr6PmMgCKcdZbVY4Q4z2KZenzBjXwK/7AP6KlxtoM5EfYSyXrMT9gdwoYQo
VkQCxVCiz8GFyZ76pfl4vydWbGQWPWP8gawjCOqrSB8s5ZetKzjQWStdNXqBdaOa
6glgvV9JQnU6RbJPt9rH05JRgO99zkLqRSju17mmkGCmHTVim9mg/dxchILshe28
wlnYhUm/Gvv6UrEPQy9JRxzqGwonEmiaVW74vYiBJodyTL6M2JjhDRn09W6PQCVT
zh77YDG61d6r0p4uUeh/6a8KhEYXGzExa3eA6zQWTmgVNrEN120Te8CiXVTrtiM7
ON5DrMhJuI+/+RDOoniJlQw9Ix4U3t3lf0RBXCXEmsdrNt+Jsiuid0hchSpABKY4
Yb7P0MhysqsxRk5sN9fTnEsUHc0E+rF0MJ2JllRv05R+KRvnR1KatA3VCrho5/IM
Hbv+t6o20d6y8Z8aL8JhV9ezin/4ifBHMLHH4OquPSkcBfJ+0Wa+Ic5PRek1zlSl
4iB7IGGC9VhLdZ+oURCsWDbjHBZ0uygwddW7ISuD8LJ7ZVnu2ooWsC4rXSwO5UIj
8mLkxwsGrqhpo560zEq5bJLRJzgTf1Om6pNjlDMdOx/wrxXHFm/74D+nsQgxkQFt
IrYA81syTVB0K4HJTXDWLMMIpBXoiog35kEe641hFNty7f/HXVtu7OjaRL6WjSv1
EAfGhbQfYdDcACYprAXyCPSDDY2E6jtvP+0WFdojDQ/HRucBWMCYHw76e2AVhIz0
+FQDuQi2HehSoPKonOSQL5LcOY/TvdUIXYrOVB2/YfYGRqOtQEnJe1lmp3tSY1y9
wYpYsiBsPACHlQIdvDxVDKnt0i/h7wbhl1xhhpB0tr1/WpG+GRobkDFqWBxRNmis
1bT/qYQ3CYFTcUxHLgVKVnPKmJmfe494eYIUwHapYAr8vOEfyzYy5CkPwiOOKrEa
mdbbEO2rf2Za+XjmSIB9Anwa40cmDgEsHEdV2+RVweN69y8HTdkYN9yvYYxlaS+c
m46Y3u6E4/HgpXMatpgNVzrGTB2p1/2o4kWrXzrH+/nM1zYqF572+ss0Cavbavo0
f5oHOF1Kn5FjAN87yE1+ZWAMc4/SP6KRuUUroXY/uhyuik88csCQcB9CkituSbNB
EchSmAKTaTH1mdf5abuJMsGKuBoO+eAM5bhOz+DrFlfVOaKbcfgqAV9lbxCtGQrM
P3PhPKkdSTmBjHsy9b+hMEYVLQXoUAnLg5v/7W9naONutOoV1TEB79yKtaALdfmr
pVyBFZ396xnyViPRatD5z8egknkVp9Tj9bmH5i1hTlVjcQJR9y03eTGRcTLDfjTH
FNynmRwmzq5D2zSDqgY9O0LUCejTtRJyMv0gNgNRireZgboxBQk5hNtZ9tcztf3N
ITEnoaajN5yNthNUU/TMGFQCfrKCN2ASQ+deojTk1UnFVqKd4W5QuaoBMOtWuoNZ
oNF+aWi9oO/WLGAnU0fLbI9H38c3ODulTU9DH0yV860xgByKqXAmnKtWaVjwqJvX
Oxbt+GF05kLMLtei+h8OtVAVQH4r+ryE15gdK4hMQVrCra1QMQrF2J2y2fTaY671
JK4faa0WBLAi7b/h8N66XeHJWP7LTjPcrbkZYYR6NminTdhN0UivzF1SxCQmezLP
pbEFEXXQds3p3CoiRHLe0JcVrT674uIvPhXKvmeMNVIQBW3v/zR+Zv7Y1a2v8E3l
RfPONoruEnmXyYmFg5A/R63CQUdi00rLjc9OF3QABYOS8jozjWRGQNrY2uReLCwm
7D7JWNFYgaVKqRH6BtQeIbJIzpo9f/bf1VH9cDUVj9/eLX6E5N9bKBDSAeLFtzdb
hDvbV9G9xJ5WrFeUf6JEaUO8GiYIt7Jg97da4fjpLHnI07crG8ZFfDtq55D5UFRO
EWkCEjbCPq4njy0jv6pArr8VWMEhQkTo28qvOmF9rgzlikBQc/Z1DZp4uuwaQkLd
O17WDhUxdCAFPPqP/CQcyHDk1ZPec+F4ZLHTcb1F5t/W3ju9OR8BgV8Uk+Y3Qu4w
j+h8TJ8qfwyk+mIDiFqhin5mYy3vxm64YyTs905Dp9Drfzi4GLr8kBqL5D/E6yOc
O843TPgCeWRz+w5OoFSTXwGuu4YoZxOU1MZgAchHmJEihcBq/pKw7VVgmoDMktpy
b2NlPRs0q03q7/az5QD6k+2X+qX9RR2CfX5+5jeHE2s8qmxRMb2tlA2xs/B6BJ6U
rO+ueQx4oyL45oL5uJGxbaUeywpiDMPKV+pd3RtYUjktJKf4nRE2bS9HW/ygd9E0
W5JTVKpNSWlgQw2kDghVIOzVMQ5wTgIsh9Gv1Cvf/cT9FYymRXS9lQ+1qjiyLvsv
ukrE4tn9QJYpW1bYoDBWjy9x5120SdrytN5jFpWfLi149uILNdCxnq+jjCU6sLLa
pRzWL1n1hU9w5YJ23S2L0Kt8vHqJsJ2TghyfbGfiz4H3dyoCYPhQDRebQMtM4u9Q
N2/wEYLw7exIMBkg3PPyLY8KtYuxhnTBAY4Ol9p+KpDnqsOTrw/nGZ3SwJKZp2hk
IhOQjlL8qmhT18JhIEELDAmWhQq/Wdoh8+Y77KqA0GTvSXghE1Nb/X7c/doyPc01
gGs/h0iU/3jDxS/GIZsxcP+bCuEZ9NB8eKeDpZfQtEYxq1yE5eo3kewZZq/aWzGF
+vbVPMMN+OrpnG2HWN9JlhJIQoERe/+eVN/TZIzfkv9LDl2+xWt1i+wy//lCiZzP
7PAS63zhMEfstUJqKGVDT1QeIug1eNpe1M3Uy+o8eBJC9hrW9p/u5V6aZuw3jsQj
8qVxf7/30iPk3qSji+P3Yyr6ZtYGhx2/pfQ1aZ7CWnZxnu91bqG7EMGd5TTNbE9k
oYRyjZDvWhIgs6k7Ywamzt52iKck/ASNuTcR23Q9K0QVNCA7PkX0aFddjlj36UFR
zSMEY09eYJsqU1/ZkcY3ePLrFDV1fqwzrlQGeLG2Pb6m2AtawxRBUUpE9daYk1DG
7npTNziKRTLyB7YFV9Il4UMVM1cITh8YJmYXrT+oR5Gb29Y5upPtMV56m27GmTlY
UL/VrhTLjjhpBE2MFTV/67oisFFGl7agbACPPrP/D88wobsiwl6qo+DvlgzbhwMl
YKXNuPAC80+qMLXyqiI/sT1/ywlrgN+GpXLzM2w+oBIt7M6xAqKfSf/szIXKsM7t
ftL+hf52YutD/bEOoLvlRtW7Rj+VK19OuqJMvCI/dCfyieMB8MKsHwWiKEca+1SE
FThfrypR2l0YVLC+Q4XdqsmiKz5VYuoEKuVHR5e3gB5ZkWuqGnBI9GhVYG7q2aHb
8t6ZEtZqCz/+JjEhGObrSOh135zpWCvoHPnnLR4O8W4oX/zPMz7gzQfFErDFlw9E
Lt5Fc0nLotp8K8Y8dKE14lS8+bG8taHRwUUAUQ/IMwVTHQDM12BTPtIzXXAx+9YG
zOk4cJ0z8sgKAq8AIi8dmz64fwwpo7kgGw6+tsE/NhslQZwU9BWckZsKlt7xrPea
iCRKu0A1SFxxkYGUcux71I1iHGeLCi7/VNqUScbBCblg3Bj1zODcLGyfByc6xR8U
gPxz8BArllSCcQgNzyNfenIZrqrRZ2QtAk2uV4YxjxvD5NVQeX2glqMNUMi0HVIE
pZ12tksq5/gyEEYQ5C+9gPSgf8VUadqtRnhS75JNiAKZixudBaGi3etaTG3QpGjS
h5vbHrbk2D1DKnsyianp5ng4RrUI/wCC/sWCENoaKdslihKr8Arsr9ddFPu0G4+Z
nbDSyWYc06mIziAZaHHh/fxrBaS2P2PHYvr8V80ubaWJQjVlWIpOH+bBGIGxc9L1
RxkBiY/Uz0Rsz8Ep2uxrkTgppA3VuWE05Gxm0T6HbH3IrSZSgtWQhij4JXrpx/Li
HJHc39QRIkbNtjgD2pG3lPeSYoBuZkvNgd9r4+pZa+/A5RJ/THfQxa9Z7jZ3hvqL
1r2wkt+BcwZjs9R5QAmIT6/3x5w524IR2/qihFyQ1hejboAI/daOCf5g17RtZ9rn
LjIV0w4pdqXLvHaVlkak4CI1RuXj2YilODBl8j284sOiDqRtp2Qo0fSFrS6uiXKE
d0Wok1YTvW/a7R2whM8Xy1omYUqX+qm+HYUhn72Kjr8foLjy4FfCuanCOUhE3LeI
Z3sXb9epcTIXF8puDZeHjRXNPeaUOD8kHwaAFo1SG0DbSO4T1nJpHWa+3QkwvnPa
mWkO7gPGdXoKcMpPhk1pa8dX34O9Dn4XSjHnWM9N/beuciUDOsCECD4HjBjuAmN8
N9h23XaHfOArJHdE2p5yfSciss4Kj0BYGRZtwUw4Im0xy/Vtuk4U/R3Q45EaH+6o
5tVYtcJcnNJ0MqdZT/aViZG3sGO3lsd670fEQS1BVZNsZHDNBQQ/ArWM0zRGrfJs
1pYKx9IJJVnvgN5r7PLBDPQvnM3wzK5CslOSctphtoaWXMf12aEODAgW296/ZfKK
KG4o63oupyn9Ujx8V0Sxo1tBcfJTbSTR0w6HgN3arkRUC3Q96T4cNp3QKnlMBYqm
tNoMsx5B9rD9FE3aaMqYPJISxj3gL4R7VqMUEm+2JFqQzAJNnkeZyE146UHEkC6d
lXHkMdqZuOdE6agOi4IdivGyyO4irThFu0KnF4At2bz3V2StT8RFDjlhmcX+2kxU
TGVTbAxg2ZSnM37a43xzXMncmx5zP6ERhtxc9cSkR8GYs7dvw+UUVc6fuRcRwMXw
aKDzr6K/YYeKuH0JXYdzTZeBSORyzGIWque0WlHvlo2GQr+905yA4yTbgyiyjaBM
pfy6s0DIVDSeegvkBOw9/vS7MmIa0b6dYUZOj+9seipDBrc8vJ8Z2tJil68Ezd1I
TxHon22+N6XpeIedfRlBE3Oy8M1lPpAR5yfOy67rftAIZlN8zd9MWa7tbnDqzu71
mWLjA/RFk113RZ9vWyZxiaTlKc4KEuD3duuCyW9USc66S0eCvcivNR2DGTsXW13h
uP7WBgRq/hixp8+IBkiWjkXv5eU6XP7DF/0WWe8EO25wNLgj/A5b89lICfX3kfni
F3KKKBdqeJJwF5CJxOLnetITkCqQK8IGtoCXSJ21Ca8WDvmJ1DotVtLX93S79KsV
aiyxcUcjMsddeim3k9lwLh0C5FZg7Lr2kqRZn7OQAoJG9JMWdu4mIEsiAPxwG8wm
x07FadNrUilqD2Muy54Eujw+/QYMg0RG5odYegA6yVGLVBTqKJsEk7O74Vztm5IH
013mAotjIIH6uiD+LxuqkCDCGAi6KT/WlBvxwDwUCWZsbBXSquc4yD/dQvVEwHIn
HKZ3YazajcJjOIuvdbEr9wh08vE7gNF6/7IgEtQm9fTon15DtEhVgd8hnVkPs6eY
QWkY99RrC3PeploDYMeX92+Cajg5Qt345yrGrXetuodR8HIYRvoSRUUND2WoeqQ8
qTuy8gT3Z9wjekLOgC4qGor/cfXpEdnsaYd+PfA2+ttHNk6lVUSUHJ1fBmXsgnG4
cgMwxSLmZhyEJ8w6uYXv50lKx5Yw1PZqqWhAW2FCLpMv42nTge4b2Bg0+u4exSa9
Og41PvCpGQ0p1gEFK/mi3KJdGk7FspMhUXw3tKN6h3TwNVVNsP6QC5r09QQu41fG
mI8QrUgkoCKjmbVIWqugSf5zMXut3kWU7wxeDU4ExsHge8ksCvzXSP9yn/D7Fgqm
1lo1xPFErn6w4dWyFFfxZq2p4ax0+q3m5z3iyDaUkRRLlSPOrnAa7Rsi/rDbzViX
zWzrqUjA3SrLbOTMIbW23ts3qcLebfW/zKS9/xZFuJvT5An8EAQLnOE4UGxjpXhh
Ve6V7P5HfROQeHiyacK/Z8ofJCcn5ohQ1F4gzE2rDt9Ni86K22JVL+uLfMdge1mn
RPu85XM5gKrfxlld7smpgy0x5W8vbAXe76mjeqlJLEB7YXYHTFISwXyRZnzr2m6l
bxWEKBBfgSZG10rm9JkyiNaEOPFyKfDdCY8R8yLNqzJGzWU9V46r+r32/HnS6/SX
ktTTbOlBITh0gEGXJP45eLGPzgD20wwmxSgU7QFIRDARGDDC059xC8WNDYApxVXw
gEoeiboKcAkkLHrgsEaa5/xQtmfaKrndX/XFhGaR6beE4/HMjdCmhzfMzjcbfcCs
qZ74Mb4tB+s8lc5whZHVHRGVV4G5ia9us3HbCNCKIQocDY2Wze1IRkUTXy48DTSB
c+nkW/nzcYO2FELDWUZnjZx3R+R3VnmTurTv8ON/KqgYW+Yqbmk/aRfnNLRM12Qn
ryQBODEX6ZZCGVqvnZKj23PGUI6AbBkI3O4OrQj/SbBba1RCI+MIxcCKOgBpXyOW
WfASWyUvcd5+J3f79OfvJp5T30YLqq8wkse5NeHxdE1aD/zTS1GO4YPVAssHPHbg
Z6CfIAWy/4VOSBHoaxTbIUwdXf2C8kwGkgcWd4hc43GnO8Zfg0Jx8motHlM+UgR4
Gd9lSV0TOP7gTvUmeSalD+NpJnX9x1iFAKTkMbXiL5XCRaTwV9uOGRz7O9AYd8dd
whrevP/CX4OaS0avjPSZ4kgPJui5SdXwMFhnCjjiSwbcOH5ivMEEmezJE/kdeHvn
SLMaMyA08JlW9Tx0qhPhMUn7OfuP/i3UDNyS+fMvhKJxOsHtPaKOppNuQzlXaZOC
MwJuH3dOwf2AYcBSMoWqL94Wxn9/CFuGWP3HJCpybJ8LNC45IOObEs++1SPsBffh
qcSyZm497O//Y5vYUnEncUy8IEbxBukwJXr/lFtZrAN7NK3ambCu9MA4LDaeiw8l
1iJ17xQ6W6K946NfeCA1Sv24G+L5qJccPGkStSS5/jbvkbF4Fxrx57sFKfDhVEcC
GUNDPUOgu05w9yU9/+a2aXho70HbTeunIYqKYKZHtLfRLpcTAqblrQXZL9nsqwQ7
9hR3DIOkOk3pZkSYcFT2uMD/wJxJWST7q1nKwTmZAp+FgGzcd6r8Bo9axQuoP8t+
+QMt3ld66/u56N8VYbfsZEhQfLa62kvkixBfyRMDfWRzoWyqbfvU6PaaSgG+y8dr
zDwiSxGRU3cWGmATtpp3CS62GwcZXL2GbVMn45Jd5xf+w3rdLCwBTo5fyPmHuKN4
neCYVqrAOk/UwpUxvgUSJ7RTY/EINk2JEyEoiHUr3bQX+W5gSoTBY6Oeyk4q7oj3
9QXkPVo2pUB2kyI+f8EY++lDgjoO+UzWzkPfg+I/9Xb4N9eu+IGE/hZ0El2Xpi6c
LN40ZOWoqXjhJ0EirgzHSIQGNZtr3u1o+AXBOMjo17UmOib+YMy5DjpyDe2ks7EX
EbN3ZbKQPBVB+FfMWCjzRH0Qbvsceg34c6AS5L1dmKKCjZJvuWt7cPptUMap4Jnn
A2R8zPJcyzJlUER6qDvpWbja+SC2XcmBml4+Jx2xutTHAxwPontU2fUANnZJ4WvV
966/7Obyn0g+uzxMniztiXwMTSis/pxyGj98VdMYzGduoSMRY/YOo92n4oTLztgl
9luTPSJqGmgVBgoG5k4PIpExv0ijsYTOUGZtlEeILRPX1mSN4h5KkEj1TIppUGKc
aI+amy/t4jFbHaS3xDjA2y3JgwqiUaLPINm6aG8LmRpQbtZwF2s11hhwTkC1hMqh
rNHCIWgd1buyY3sMYkqFWdLFbBFvt3ZfUun+KV3kcZSb/cG0txmc5NhaSkOYDfA1
vx4bU8LsIPeaorqQPy0+XzobqC2HogDEovVnLXG9Zf6AzDzn2mOq2K6H7ZM++zeq
Cjqs3qneb9gClVsQ9+1FtMMtMac33LG4V/76izOcLvWsKKVbQs0tqkedxS7EObPD
2ze8o2eKFYBmCYeIOUom/H7PiRON53i2bqwG95BguoG9VQXa+CdLPb2tgltESAIo
fliZsI2VWAPRtvp0D14tlZPiu3bj//VVj4JKLGw7jcQH1B/0FpFPY4PYzg0FDPOz
kf9Cq5aTOIvay6sP1ggPxws5ptfuyC5ftpdokHzRYNVcSLgGoRO/QrcfKaLpDhI+
L/wpXzGkrgUCRneEba8DPlxnasb9cQ+kmueufkTuBqlT+9xXlqZf7Qx0lWP6Z7bP
IaaoicqRmiJzMWk8aIBA55HeTDO1OTcxQza3oSYrQafeaR6N/4KwryOnLbtXowuf
uWiXYHieDcLHoX/tDxUH9DiTItZwC1G1Lgd3PiJx7OK1DOzGrTWovsixXiM7VCKY
vWxdYKC7IubmzjkkBwtqlc+XVyfkKYDiIdOjyque5VZS4XNqTxl8sCNB8XCM7Ya7
L8g4KKesn9ZObrTKPtUvT/qNqwhwdw5IhqJTLFbjXoaWE8CLhCjjlWugVRUTOQtD
K3PuH739KLb30wdTZ8E9DNQb0vSRszwX/UoJ5VUtltUAF0RzK8tnO1lTGCyychsB
EPEh2VNyhXZpM3zJtYdPta1Cbq73kb+gyOd/LNK4xIy3B0aKRTpB2k97pCYhTa2m
KV4fvEf4LGfTi3orntOjyYBvBVO4i+bM5ICei467Yy2k+v6872EzNdK1neGwl282
Xai3ZETRNLRo4siOWafKPqPjw56GUWrwGlT2CtKRoNe6yMoU3/7PyMMHXL2KG1SW
3FOLw+Jmy+G18rP1NqKk5E8XkB7OFDdT10dO6YD146tMDS5MN8kavsS1weNq5HuI
Z+ILh/R0Z0rNYnJDI34Jr54DyHM2M+XfYaw08Rw9Bh/TxbD2uPFC1RnCY28ph85z
acwAhi25joe/sYzSILMXB6MUXOTo7ijo0hGYlMsAER3W0TEY9F3Dd8RLY2BKY4Lj
yQJFmg6ZgpzMi9s5moMcwv39VjjignlpgYC+fvifCj13Z0vGoHequV4MoljZ4kkC
HKSdWynVMKphiGKGRVhXBpuBlQUCLUJEFdveBKGPrFiEe1dgFeczBEkkQLlM53BZ
3UdxtGRnfE3VsS9EpV4z3LbYR3YK/6vs6cjBnkUw22uRpccuayoWnvEnOFXWU+++
ud6GizxbLPbLU8ktxkSreoY7rVeBZzASJAvN8ypbQVmHLZtt1HxfngPBc6UaWxZ1
XjKpuFMdOjTrIbcxGVMbJA3r8tU3usILrChgXNPZh6mcbq0Xk3HX8l0V4Z1mxmp1
3hK8MpXkKLL8RuhEQbP3l3oL1JsynayGMlnDdfrQlrl3BF8jHFyz+8WFP4gFPuEL
rD643IYQPjWom96Pq0rSRPygIePlDlCMrieESURzAxRk+m7bKpIXODFnd97Z0Fq0
PHsFXsDOu6wj6ZVDn40CWN+VN22Lbv+x1bUTFfc47L8q8zxmALBYd5xCH1coJhsU
sgdjJVF7g6SsI8wrYi/f8dBJVrrT/Kn65lUiSSe9oVrGLK54L8DgPRfTf/Fi3P4P
l33CrzXBWpk6YrpUp7ccPclLSIdE7m5jpT0JGKd+uBnQDj3GhBakQaiQUtA8X4js
n2U5InwZ3ySHa1mFvPEpAPDtPmoNmhh4RVzlCE0vVYmFQFHuyAVBJCRU3exJ/YuM
HD4WrE2GzjxUpTjQ1somogQfZPibvCl5sJV+1w8bj/Qgw1XQqIxarKjws7masEoV
MUnDqPGMtMG68zP0f6LjFstNFz7IOeD3+KG87bD1D46fQd/Znwl1AOCi0nYyyBU8
8jKSc1rWeuZVsCOeWZjYO5rVl9sTSpxOZxShGjPuVyVPdspoNUeMISkobJS429dK
fIpl5PeEXisBPqdyG+I49SPxL449g1RneES5GuPZJ+4JcVT+kOq6LijdSuRkjnDa
9m+iUJHrAAC3LSs/nW7i3YnsJltu7mzGnW0W5LS/lZP+ty5N9Z2OvFSLV6FWcGMa
ubC6/HvM+htuoDTXXBsfaVVAebcsAM/PMMjJF9/HQ2bJq6OcI7XUg44yaR1tDCWd
ocAg8WN1MnKzAm4s4ogesM4zvwxbvsbmfIizjt5ZZSpEn1ywtShhfv4jxkwVm5cM
If2MqQ27Qsv7MVsPPDKUgwvCzGoCPeQA+urc5wRPcW0eaUz+Iy4vqNxr5I/pNS7C
dpgwE9RzQF9M7IsztBUWy47Ams9kB1dQ3ZTuqqcg9MYB9wvq9mVc3MkLbMPpQ77X
L8QRsrNzFDhduPJb1XBLuAuAmBreYSboqGy4aCWq6iXrU25uw1kr4oVfHO4zQpqa
6TDtPeAgELkMrp8dv2kJebutoSV7ulaJwGLTYg+Ov6WOXSBUsThFRAKAFW61EM2B
0Pvh1BzpwDjCjEoKzdbVEEkNUzndiMkVn3l1jCVjnUF1tv/JzQXULqTdgMOXF558
7N49/YD6UXvPfMw0mtyT3MRWVKCx8/XsmkcVO+Hv/6MPN9HclwbVpj13XGPVDHkI
R46MiPKrx2mY3RwjvuTIVy+C01gTRkw9FAgNcbt3+Dd2jH/CvOURtS3mopy2QI0s
TDJFO3y89/7L+CrzXFLbac6kTHzrizH9qPGcbA84/wYrFppHP2ag6ewf05MvkVH5
B6OfKh2G3SxAw1ghogUH/GJmion+Kc7kSIGgT2omryZ1J5Hh/4Zmstfj8AloOwhm
NkPEYwFNyZ29Ag/Tv/YsoXUMiD2WrNjFHSlDDrnyANjg0v5id69SI9tiIaArGEMO
rhLLG7yWA/KtwsfV/BX74som9hlxu5qZzw5WRwrP6Tir7rg/XSSCHNa7zHpZA0+w
Xo5z6G6G5h1uLV2GLS2DhFb4Pr4YzH/Bu/c//bBQBXkfwBM/AxYuraSeaEwO2bNr
mgraEB7g4ShNm4vhaHkB2M04CPXMjF2d2EuTonuN6jIidDsDEoEHJmKo3R/o/N1m
ocAX3phr09YDePGgSgQ9tjX+fD0LDFGYVLmZmM5J6zg/mGoJMnzwsjwlk7e7G3zV
noACLu11V5L9G20pA3rYsPn01cvkU5cLwKwIrafgcC1mSHfdWsiaKZfOXN4M/JpY
0OM8H4OksJojii1wPwJWrvzzSZwA3U8WCeeMHTTq8/KfxQiwAgxfb6J9ccOf6l+v
jBw6MEM3TkYKDoXk8d7FyIVWgi85Qf2b1p6gZ3pzswNKsCCShqHYC+XrD1+nF/Hs
ivzlo5xEFcWIcnsAX6/BcbtDD9/UBRSiqbC74q36+aKrHu0fk0KxDfginepFs/H2
3loO/HQDq5XEdw+Hscqk5v/UL7qvtJ3HwozOYGdQa+0iku3DqekH4lHp+NBJgiXJ
GOxZeCWMnxeSZ0JU3Ab3zzx7XcfgSze4e3mbyH4u8lLLYtb9MXFT8b0cvEFjO+cU
bQXlkTo8OvS/13HkV/ueioe25dD5+3A6VpEXQVKKqFaph8LeaoxAC1llMLV4ENpR
6MN+JX0wu05cfuetmrSsdgQehBz7bCFXHDTD/Lo2dVqwHyQPjvh0PmIzha2kyHqM
91f71uZHXecGI2abr2LnZPodPtWkc9i1trQcGP/DoeSBqYWVt1ReUULxNctoc0mV
0jwOz6WRkwYrlhDTvQQYe2R7q9giNZtrxEaEdXZvFQN/Pu4Er3e9prmdwzpoG/nQ
Q9kd4ahjO24YIUM56AT6DehaKVpiRgLdXAUZ2Im3Xkz+1iPzaaT0If1VR69yQFb2
AmryRl055tetHPQDGa//gDUCalJ3qQnPg7Y/tlBsAFcfUnap7x1YwIdnjE3nsRJU
bVo1zuIIyoySoQ38kKn9wFzdun5u4CUSbu5lGmONUtGve6WF74V58wsyjjzs9/I/
8sVjWoV8r1qgCsH0yIWseLAcSd9zGPT2guBzKtIFWIt9yzfDC1NHaXQ5B+HjMGnP
M7KuMlWxFRx1zoesuE4qMgCJ+e5GGQoyTIowjjGWsN1APVujp8WiIYh3EHZFtDj0
p0rSf4bmEBWR5Qo0Ru5AhsuO4vzKmLF0UTmYCq9pZPNxfLKYyWEltfzl7LHjEgk8
SPeIoq4JoIXSPlxtbn1qKM2qKocLr9iaWujygg17PzSdi+kDi0/CZYNYyTiW+jHf
g+siL82ThysVauOo/MCRcsyUl2i7BDemu7T/uBOX4+xOI3Z7Wm8SdUPX5066kfJX
y+2YcBPT3OhOHwlTb2hAuqLssmpNLMqEAHNVZcNgG7gMUsRSscosYbEN2wdhNBZe
ve9Vwlq/tWaM2V973su2Vw4CuRu3u2W/c8r7LnvtIYLLoGqFOxnF/+hczBFz9aPe
/SGY2sl1BRRjJM3xKOREIQ7FyZKjHyBSZ9eE0cOF8HpmmgQOCcbiDMBX6g7glAmQ
ZoTx5NUOMXOr4R7OSE6PnM27eGSFDVZR/s42QSLCYYR+gGz46pTWNSoeRTHqxMfG
lKmTYBukaj9+e0gosOqIOcW4T6uolFKMRA5OqtYJdHPskO+xz08Uc0EZduc/pXWW
j+OQ0Gl7vZnUnp98YmGtFwrviDqE+tqLzhBbRxnm2K1fT2HCGfDQCVIL7uS0wKMP
LeCusU/ee6tys12hQH83HL6ZyG8QujI5iD0dYmdOukcfKBClPMjvuPE7LOYsQxK7
lhe6ZVWXVUiOHAhUulQJiaGdiBaH7kT5NYnjr6q5YVuEX+J3HH5OeGlW7y1OOpY4
Eie9TGlf/NSYr7YkW/V2CCtoo/1Y1NqtIlT7c0KMVNmpV7HY9SfpE/9i67qkYAbp
54JTn2jT+zYOSxm4Eah1/dpsauo6fcN9Xm+w7/Y4S/+inS29APT7MhTImK7so+gK
/Az2N1VeasIPkW3s29mzWBvK/Y70ZxGdEMcdBPGKgio/OZqZuC13wmRFPH5YBOAS
EKjcnegqT5RlHb6Vss1Pc7iR7iQmOEmaMxPo3uGZEU3rd34q0riB9eTeCm0rmKz6
aU3mpjIbMEcNE9Gu79jjNBNapbR5Tc8wrJ5yIo3026BxdGd0vH0FTtXb155dT/tX
dqnrY4Y50f6utkWGWFdkTPZ106Hwc0jmirIQPBm1ts5Ly2qPGOOMMtId0L7Lyxyu
lP5QklvHMAipvxKrpjUPWBvWERKZ7CoK7YoNQuW1fzaiK2eGCuoohB/qU4td43iP
sN7Jkoddw9FKmTwDesUzSt3x2W7/hz2RJj/QnJT3kKgdJl6xLoej4XLAjTff6zur
jr3fESXaF7x7PbnZbt+sr/eBNWek2UyS77fxmmxlhpxjz8SsxClM9Arp3qcKdW9m
vR0Q/0+x8BNGWU7irLhce1ZGR6cfDlAp6oW+dzjcaC4xt2P4wT4iaXjGRLfg9g9C
aRLGQ2gn1wgtgt7ryghvncLiCBwKsGTOoCZEWGo2mdiKuvFDdwUkDnrt0rIptPqL
6KhLdxMvqsinrHJavQSdYWPv2t5tQjr2krkHtbiH9HYJfOqJVGPieAUszT437Eh2
JozhP3sYzdUq76jihIjdxzVT4y+Hsu8z/WmMDAkMJJS1lBsueDdyY44tIW1lRa0d
fpdfryCyGi03YHWwly/7VghdZWmkpSdHc0nGdbm8gvQpAkgf9/49zKnIW6xAG7QO
AjTLA8heebs8igN5aKSh0Z7UCJSqneIgkOvvTBXCYQ7rT6xIjrb8SJcjNwAIK1AA
NjeUTwYU3FN577PG9hwWmUf7T+XDZ54R+5MRztKHlKXMva2ictiGYcTa5xWpKru5
iDnxPJlrO0LYO79blvig4F5xF2vq47OtpeZh+5kmaF0vfCPQIwL0eUnI1LBb+jXo
ZzJ7M3ueZRsCNAXOF/3CxWqMGuWublBZGF6jD2wwCje+PIWId3cyAxvdklxlz+1b
HlMBaKuSpw2hbZJHeOPRzzNgC3T3pYriP9R+inrUU+Mbyrv2Vh0outKSeq7z4iGX
FZcImoobTuVNArGX1UNhRB9S4iQTAXWfZFJwWdUnYfoupCAEqPx+Fa1VfMcgqVTo
Diqb+LvoyYOJQWGrYVgNm3tJZhRYI6w6W4sN/u66bGyDnJ0Dk357kqI06zqLKqud
zevHut6w/cavlOzpUpkJRA8vuEIRGddUr6EcOBnDZWMEwrpr/vLQeVlwQGZ7M5gj
oCXeT9eb+NChAGBEMYJhLC20kG+KOj6lZHwEGH4P7kLcyrs0u17IePScl15jBq8n
D1TF7Oz6pqRDVClKAkX5C8CDuachcrDVwcJzAls5vu2J+kJBndWWZl5Ga7eM/wIB
xoxXnooEs893QORYCu4tMKS6QgVUijdfdLHIRW2OQldmgDo6r3GoirnexKwqEr2y
Ruogg3al23kqTNfdWNiNzMA0Sc7tEzAhfV3n/RuYDXgrZJXPPXBo3SmnrdqUB71O
d2xsqpLb4qzqsiLgvhA9n72yK8xjB+JAEbGhVJHB4uHQBJX472OstIdVYQTZM6hT
2PhJk6CGQ149zAYhfxaXDbezEuUMzqBqFGVozpVuiBbFaZxgfwjIr8CLMdXm32D8
6M7kIiHGayVYiNkWKFV4eviItdY4OhR7/0STjN4EzDSx2kfPtl6GqASMqvmMsY5b
J3bALGV0vApFWn/s+2BWzeFzDLRgLRcLgb8fkEWYq1CRCJFbrLsVemPyqDO4p+Fo
B9ZCp/OjEVOy2WijjTegqDb9gP66NcE6Ukp4nLxF3g6rrgRLyrxM+NYBkiuGp08G
hVo0VarEWcRRmQXQ54lYrA0TqY4lvtznZ5s5FiFm2asODss8zYEsVfhyPZSX3LBG
zE273Q+TCzwnpE4qk2rUaD0RCtgApLcaadQlYq6wfEJ3lBAZMp+rkeZ57wXl59OO
NpAmnT88daD2xQGdH/Q6HSiUV/dRMXLLlMPNRum4ulOWXv/jJDXKIVq9exLM6lZD
UagtVV4PtYKnnZl5xSM3Jp0BnI+b7pWanIBtVGZsPX9fbC1o+5pv5OncjaTst8Uz
gizIYA3jy5ppd0GfiMi9Ide1stJPTeVaMGg1RtUbDFrTR2koGTPwztiEZiOR8+vZ
vEsS9oZ2Y90FhUVMyZcPS59Lw8lWMXwkgfUpYZQcvnQ6NxZvwL2xYyp/52mGBAP8
RQlds0q/TbBxVv15d1+ecBdFimp5fC5aK0T4U8T01myvLNG45EVBgEG02fHUwzgE
F7jljVIXcaubgocyDeq9InWcycoGO44tzxJd2mlCZiSga/6/A5DoWdhXLGPK5uaF
ZVnx8aOwmZIo5BcU0ZpAruEIpUEWVCyA6HRJLAGdVcDjwru8fogh+5UjEA7FnI+x
VZ1l6CuyaKb0asd9EeE37vFwx3rClKKYg9DMaIYTKBkNCHZToJrQQrD00s6tZ190
LJgXG2dikoXfQHcDoNBIhVCnEKIJRc0ySuYrQEPLWo7inWK1giym0EK0Jtb8U/Sq
9maYWK1TqzZ9pzgQXXqdO53zXO8Un1Xtlj+vKSM0z1lnJnmNmRF1XmIXTPvtzVbU
PmmWhI5aSyEVrYfxla9izsawfkHZHpw8Mck7F4LC11pwKYbRDcqzENlAZQjUe1ll
ZDq4MCt9ztd+lZ4lFrmisxK9pmGtXwAkPMBisK8uEkjvM+5A4ISlAtrrAac6lRIV
+xao0rAVZzolAU0S7wNmb9wm85TeHdfTn7gpA8sV7JSAqtYnd4EfzWgLyawNRy+6
mIwoh0IqXZ9y8z6Yb9TCePmI+YVLd56lU5fG6cL296yvYs2vMJnbPzElZ9Vz+2LB
dSA7TMEv1iVXGj6y0yB2w+ERqa37HsavChktnxTc+VY7VST1KOMBaap2H+kjOihA
XJFRHT7HNvrmnf/eIXEEQF1pfiuYWkmpmepAgxkhSsHIMml5Vbkj42Z5M8x6oeDG
TbqXnkwNqfc/wMyavI9DkiycbhCbAJkMVX2lTdFgcMKUuM9bAI3zws0+oQc8z13N
ZINuOWymNZ208YcjGGuJRYSt3YmpcDekCOVNPJhOtZnG5F7nEObVUbXacIKV+2JF
JPdQcqTTMxqbIwO9w1sRsPLiuNDAWnMFFLzUQxhWuwQqQJYrs65t1yKvcFWycD+i
Ry+bKhgw5pYLuvaJKIBMVOaVJxHGGQhh7NrAgSlLk/Zgq1CQCbhZQjRaHXxJXldg
pDVvg1vgEjlbxVvoacHhunwDN0u9nFBbsLA7MvY3Xx8DQBsOBdsN4P/oljYfIwII
iMHECVjSheIpKqvv76gqsWS0RuvoXl3ETqbWMSWkkfbqQ3v/+I/DsNkP1OT6hc4U
NP7bKZE5DWRzBnsMEDezIGv+SalA4RxQ2NLGsa+9Xo2W3sj0kD8DpCW4CaSANdNs
r/k/eGbe7NRaw23zSqrxXmiGkO4x9P3tJf+vCSojdrmlpYCHhNBlRyJnZ41aurmS
KHPvQfnT+VHlbmwbUZV1chEwAVy2gwDlp4ZF0U9uZoXfr8K4+K2pJzSj2X6Sqr3y
4rz1fqp2/ha82ZVYqrTCQvptCx4i9ue8cVIuUEDxiWGFuZEOD2mdrcDP54BRcMM3
IQIY5byu62Pu/ftzjUi8skq04q4CqpwFDVtkCKgTSyaLqhy0/9Ufe7pNhFPribFQ
NjqD4qukZLmJZ1nqulDUKwRwvH5G1WWEuPwgarTeqTns+NdoaTExebb3ldlqpTGX
xvTmsYSVbfg/y59BZyzGNmH0LujxRKf9pWWTD7cM5tem7YQ+LgWgRF5n7fBWc9HK
kOSTCpw1QmdwdmDka7TRUVn7JJqmj+6PLCF2vpq3ejbc8h5n+vLN3ldaHdjJN5Nx
PnneSxDkannaZOvS9oxs2CAhTRNWFzHAHtGPbXjd3lLLH2oEcoeCYQ/oiNs/2H0N
7Y9MVLS8Ecz++i8wraRW1GMagWqh04VrqXP7nPumn088ZqngA7yAa3zU8BiP3o05
QwYT68WiPxzJqilOMS/KI19cqb0eAL6uMA2qUBJ6aY1hI+/16sJM6DV1ZdtrlgAm
V2wjQ9AM5G/V4f87XfTms9vMDt0/HvSmy8TAA/daaDntazDBPoJc9UXMDsSGluNA
gbMGEeFtFd958c3jUFrf6rQC/pDhLhan1p+JVKp+BX8uTW/Hn+6c6xQHB9S04RXv
+JSjCeVqzud3Hg6+i+OE5sfJwn1vDoDQotR/FZQwnbc7MQlfxZbaWYcZThhyM5l/
wsr2hOyiuv59eSs1b6SdNGRIYm2hJHdeV0Aa0fj0jQxUwF1UYsq/RiMiw6XzrBGK
loFVHdVcrq1hYKHddarFGasomrMCKJsHqVvXr8GYwdS6F7ULcHUjy1OPUhqY8cl6
TF6TIeFD/vu/2b1pCpUKIU8hJXZrCv02YnvBId6cH/7u81a/Q7yMK4AF6+67Zbh+
udlfybJBMGdbekkpHg7I57JFXV3suVs8iryJP2K0siHFgUkfNDsBkmdl+4075HhO
TnIL3chlSDpP2dikjQQ+wTD/lOgpwPgTzpXcKqVMQrTMivE2H1z65X6LpPmYPzoP
6FS5yLSuAOSPFltJnqXcb0eZWs1KS7m1F7sgC7QzTgJa7142uYR5YkzHgHxIZI91
+zOfnsb3YWuQhv/N45KXSktS4dnDEEwuHjg9QCgczjVzexZPUoICYtAMxOD48++/
CVNSrFlM1lbaH6tlMLrBm6eGVs8O8UKjuq0mNb//ZeGZj2VCoPCvS6aFvWzEV76c
Nr1V8WBl8w5JLumslXS524HH8RSfrYo8whLZr49vROMQG/dmB4Hhnp7zLuTJ7xPz
oap7eeg7EbJxWQUz+FOlf0S4kNKdPhu3JC9sSDlYc0/vy1jkJ04kS/QxRTwq0GOB
nbNrOsCiidJmhc5fkU65cuA7Aj+Wp8m/ynrCuR8JyvB3uPr80Cv+/2h3+QUSAZhN
BYRBrJP7oJzJLXjGkCZtUCvOSHXgtUGIjmhve52fa8RidS+o1ct22osgMiWIimEd
els5LBPWXiLo15cXPQM8hUq2dz4JnNd3/IssmhW918WxAO/JAfaB5m5lLaroS0dB
StJMoV7dwdiJlDte4+qMV0F34IEQr8u3gB2U/FLDykOQh/nNs7SSh/PB40gH8ZrQ
+iGzkW11B1/mh5KiAdn5Y1vs1Q3fZ8Hwwl9+nn6agQmFfs6hKZLY1KH9A4c+F5eU
p34HPamx9OTX3n80hSsefQeVdLnA4Hh7UpW3smYBzcprRMnlLULK5xl5r9nadT/x
OBvwvldSEIThPOLqyi458XAPcdpvTADpXKRBq9HMFBRSkP6TC07whLVXQVSyThXV
R1LopH+c8ZyTCAe6+W/X4b6iHVN43Y7hcehtn8WsLnL49p7ZxTGY/WMxZ/b5B7vu
Dpg8C4MLc51tIC4YISnspeat/9yM3QCoSw6xgXGYKQ+Uww1NcwfPZBDe/zkzfq1N
+uhcDee5W59VULbZ4PXGr2P2pTxAwxvUsXjI+Mj79DZ7zQoSrPpwDwDV4bHcFQ2q
hbFIIgJ2MazpZa9LmlF7n4f4w/WUz0qWPgLxarF55vlhyf9H9/VoXQlPvy8UK9xH
on9zjl3wNq+IcMH8+B3D9oRf3vMSiTyxk4zTjV16TR34Hn9vOh1GMr8fD2HbyAMP
xbGnyjXw4JWyHjpb4/qpBtg5OZDcCDyHPBGUlC/p+wBiDR71fufsx5iOuw8OpvA4
Bh3PVDksKs6GJ4ivdoeZopLXyBtOg/vysRXzjpFIv9+ge7aUjO1UaWMjL/9jMOxo
bGFFrHCWptGUn4+7CVmJHa4hu27R3qbVydFDkgp5AaGrfH5xP0GX3iNRhuDARXq2
QVQvbbUci4P0Ax/gf22yEpb6bu0c51B9rFvwH0xvRh8cMPWvFKIw/t83RiV1/grY
a0h6TPSzoqXN2KVjPvH+XbGFZe42nbXC8nclHrgslZKx0iJ2HztsZ5aBUoFKzWbc
RLN41hArlr6nf2TRUEVrHouFH+hn92BHROFdvW1u5t/iGOSDu+4hDLa7M99wC+8b
2Ofg5+IythGi563n9LIHxE8gk2oQY9e8qnpaKTSo7FXI6YyGn/s8sRNa44GSXTGX
zVWPHzDUGcZm+7L3+l5oa9iflrzbr9VxK/1HX72A+r7iH0Ekj86q9gWeUGE+j75M
RpB24wjYgf5xCDv9CdRWXXXECj2+QW518yCGcjv2AFsCC6V1JCXap7bYLC4iiNTj
bjTxatBBz4TH7ECTRUsEoyXShzMWBvz5HKd6b9Vw2WS+nbxNIrenGHDKLLo84wlt
h91wcxlt7Mgs2iL4R+d7mrncN/53+La5zpitFwrqzy2ndVLr8NgPOpqsKodHpcwr
epbKHDFIOkmKt0ZFp49yfghhkqo9QXvG2YqxhAGpSrNdIPfJWL8UTq09xY5pgYuE
fDO7BAgGaQLeCVy+tf/MPslFaRzsoFoZgcjEtKtZEUVeZ3FfPi3ttpBMCyeW2d0m
18KTQTMkD1e+ZGZcs/3ZTq3rTjY8TQZ0V+Osrlc/f/Wkl9nqIa37egvMfXz92jJj
e5A6BbWLOf843+HHvZbz22thJLTIWY2ToeKEZVuuImSrZsR1QvUgS2rRhBM8VXPa
SYvyi/AE9JGwMaqia8IUsqw5QriBjp76hz8FaT3AspiIpTPnBSF7FGgio2CAPDu2
Hxj6o6skxpH7psufT77dTCPf34+f+kh6vQDwYS1fH/y8x4npHJsY60IBPunwh3vX
xfgQy6MHv7FFt+c5OVnIyDmbkFXj5D0AB3b7EdKqTzkMKyiOjmorPm4854nHZEeg
mnwbsMYo9nvGKvYdCugNFURtQeuxWX8tw7D+yTVZE/uveLcfDKQIc+b9lxObNjd1
00u2kUfW/LIBIelx/wTJux2PlxrrKKnwkFlMoM6FAe4qp7ZLUmh2VPhB73L+tqgz
Ovx/gxFhl1cYigT123cWutskXxDFKN1QiBR9Pm7BHxPXra9T6wlLCeAyigilsD9E
yboMLIUd9yI6LPb1f3UUmDlEAJhRQj1S2f1bnr1t741j0HkAuFXGGX9Y1+e/k7eO
kGG18QMepyzW3TuoHEbOYm3M104Cih6eL4mE+qFp5A+7TX8FUDG85etfOjS+yIbV
9nrjlEsQ0OzIq1op2uqyTjqsZKQ2TrxCTA1fYkkDbkbYlwwZPNwaH44wHhacQDpb
dDvXdr4TctwLaor4PeGV+YbB3KFTDGifMw6riUnxZ3A8+4H1yH0eAVJXzEi0UA9Z
qEN8bWWimAVBsdk5nudlN64OqYHIKPaQPT6XUUikfJ0lHlI94dFR4U4jBeaKDWhL
wJvl3ife32y0HQ4QZR0l4y4d3DDA8tZv6tXJ/g8RL/AIWNxeZhawwvNaafDnJ+Ct
VMYv0m90lZzHCSTOLENtFxwJ6WJkt16HwJc/lPlr3lcbeyGnhEaT+LH1YsysRlYK
IlDVmtxlGnBAHb70xW4I/+HloqgaombaxI4j2oMBHtEBBV+yMvWjVJKQnM9V+0S4
u8JTHjXaqHt83ZbfAdJg6/X00j9nA1sQXdxl/P11GhNJFb8ZqYscESVstuYYn8uG
GCJlejmZiMbKz+STKBFMRORWXy/rrvmfj+oDI69gjfZ/jGfu+jh4nnwxD31Nl6RE
oyApWI9OEqrGzCopzpkCiCUjyQ2nn8EfAMrkPwN5Ni5S4j3nwHF6Bf7oDWAA1xDL
l5pFX2ISn3MbgzWUfgbPezVenjCeUnLBb22vsmYqJNwSIC+9zlgEADoKTNcB7QzS
QNkte5PvZPV5qnDJt38WfjKSPbSja9zluBv1HiF4pbTr80r69fQvOaSbaL2fsFUb
fCd2pADHInlkV2MXA8fgajF/Q3rKqp5slqBXiINZNbHcrem9MHZLpRKWOSoBxejZ
aYB1zesFDv821VGaHYGlPH1/UM6OpPtg7YRTEXVbZNuph0XntWx9MECnGv2nWNPo
KUVPmsqjANImcaM8/aLgOtTXSLUV9xZxO+cmNHViGl2rmbrIWy96WTQK9DK1cH9n
OuUnYDXztVOav+YWQ1OnWpzTk5/fCi20RWIhbE69mXHTpda/uo/5jvK88i4OCvM6
bwPsXKS/vZ8gxIDXBsMgSE2V30Wxg7NOlkkgjcKVUA0iqiJKX7JMC1NMb8+TkH9P
syH2hPII/H/kMoy3OlOSUv00sUdazCipOHSAVGs26WpTn4kAnlUCDosecgKpihpf
kLpL/y3uNUMDZJCE/gEJDF4KBBfILo8DAYAyZvJ5dIEJ9jNV/CnlquttaLSSj7T5
kUCjxEBlAoZJvTkSe1qQpfklvNDgbAxMoMcO5eAVtcYIaktywSa/1NvL7XZxAUGb
ad5l0uZAn3hAG/xQtUpmr4rMxx5jblx0zCM8AiY7EevAFttOrxiaQ/xS9S4Awg5u
yPSYxCZOsxLwUSqwbEtzIKBsONdjC4rY5Hay4piX1pQ3Ca3FHUkCZnv7VBB3Tcyy
s7OyLEivTm8b9KxMbqcfZdegr8bFzo9P+zCO2lKBddx3r4gOkPG9yZ7OqUWw+9CY
RozNnCgJRSdtUGrami2fd293KZ8SrX65pHJWBBqwO9oy0R35d2rvKrJxLGF3NKOH
qTOG0l3jLjvF/cG7J+D7xOLPMsipRouz9akYagdtkKAqZV/ZXCf7tAMT7lqY6iqN
x2PoskLsIc9TJ2CFJsoXfG0dbmskX8CfcwXnn94MATRUXh5uDT9R+gcqN1tgGScS
vemR3zaeNwOhQPK2ikDjS2IX9wzEU063CF5mliMtmrK9Ayd6WpNDDMM/QcaHgAWG
gJV6R7DI49giYrk5TCckDvmqT32GP9XdAK8soD3Foz3UTOR0w38JoS3HsPEEAknm
hw96jz21KaS65zDC/mDET/NEG3sZTFpNgnqexmbX264xiKIwMEo/NZNSGfIYNEoZ
psKmHb8cM6DLiUOMAZGKUrfOmA1d2W/OI9axf6CoceRyznvdT9sDaWWVvLbZXhG6
v4RMHSYAFN7jylcr+9zrobtATBncS4xg9vEDIJUiNh/Nn8JUhwgcEDpA3ApeoIo3
rAOrnDU17KzOTDb5PzYnVEAq9k198G8i0tTbZ2bF5Z/Z1UJzlJ+m+ctUA+NUgv0X
r6xl7NHklWiHkPZqLtTa+ZWQdlmp97cXF4+7uGM56Yp9tVpsEi5PO8nfXlfjOazp
G26INbwBgU823sjphtciaEEMZpF9pQ40FPD0xfQW97/oLmdNbXV2CnzBINMXuy+m
dn4UF/hcHVTEO8OhKlYY2Ul1Rgb2dI2YoBSQJ+exMvp12mopNJkd484ZomkFaJ/Z
tpKikeIr+9IEpuyWsKANdDlO3GLbscPY4iqW6DxoQDubmfQdM5lp0hfi3/1zHBSX
tcaT5Epp/R+l+RPbSPEaO/19eWMmDMiDTXHFlMBJ0utHh5LfNSryAJzhuXLrfeye
dgKDoB3lrZXLZ8WP7w5DwsBNovgXlXy0SpApE8NhysHq4NLiALQD+/+oFdiwe0L9
onMfRXw3nsuVfZtl6aZQPa/shueJZSw6Q5NGIUsOxxgJ4kjBZUl5nkDMniwqNIsf
dQTxn0TlO5pPWHWVdYXXQ0uNCf32Gg0kDzVXerzOG47DChZMh6PjCviFkvrNZtgp
iNeNLHlLeAVLBjTDXIwTzBfjZJwP9qutU4WZ5tl8y61A5rfUqezDyGoHnrqzggQX
q7mkYn7hLz9oHHMRyCxkuB9fn/gEeQPmGjbxF9itTbGyT+iIfEvPDDyeJ5qp8ZaB
035E2KiMxHKiK/GNYBL4xFelno82403bEp7a7mUWwPfMRKPiIN2WGdqy5cZDKk36
tiPQrGy4HUQfbMb0P2O91t6rqrsa5kDxhL7c2jdy7RkNlA4dP6ASVJ3No6qbeQlj
vcqhpfGNlr+d8dZ2ZhrM16hewxUlFRN4sYDf//Ocp9Tlonm7VeVkCKw2sdRUfSQd
urmWL0ZD+tHfIbLZTF9UjMSRbEbbwUYXk69BsGo6/vGTzz9hVFjRpKbufMmkH4vW
bndRJkZneZYC2sDrEEJjHw3ukL5VVQXWWjOs0R1ppnkM9wYzQPIv0JCCGJfy57Yh
LMFgPR3GA8xskvPxmBwLObl34DaQCDlYMQjLjUPyTpeqBx/N07E91aR5q51zdTu8
5K/BhESdGJOtWEb50TvPErzAwKVhkMKzJXd/kHa1TLkU+BaiFkCWLEt5CXAYeusb
b4CGUbTcPOH/QvSUDBJCdy6ZgRa8+YBGJ/fKbHNylRAdluI2bZ+Y8zDu7WjRvbxo
h3Bk4PhpKqmCh21AOKgQu7Tcx0VJYd7eb3k+D8ybniR/e8TwvBsjCKdqXvw+dcbp
WMCcqAEfDFI+XhbH02cMq1kDVHaVBoW9GmiC9fW0wRsyCS82U5vQhm6c0iGBOvMj
AwSBg1Gm0b5dU/JVUlKDNUkh0Cfu2ou93gBpku/1oUzaNzUr8LdHaoke9J1HlvrX
LFIXaYp+bvwATfFnQXBQZoabEd1FOgBCMpn73UtH4f0EsnwzlA6eRRFiKzsZhrvp
qyA4zONQHqnlb4UnwmSgLxY0kUeytp2IMokRL6dMuUCI/X9aK4S0n/0L7LXr1Oxs
q5ABBNJhUzN3BvvOu0GuHCS4s/NSi3yo56mRkGXs5tyuE7t2036ha5x2kyP5lNEc
ZDmaR4JFT7RnClw7aMawKB+O18ZvQzGD9E6xmn49k3na6OwVkPpwtAAWaphYrV43
A5H+kJuKPzUPWJHE6xauMCYzT7JbdahnFoOJRYiQwGuRCsv1oDG2gdbLvXTnV1wi
SgH1mpRLd/hr2grYfeM4ISZop8IrXD4fR9UEfYeaM0wYiMoAkN1M/DlGmmOgx3XT
Xwwo3SnZ+G+BnYBcgl3Wod6cpqjQfG4M9hBiczNkdOxMpFQewP+mW5hdplSh/TCP
mr8H5Q2Kut8kfUYLEdDJ7VP60xqygM3CHsZvMNGzOkVD6ZTBKo3laQlOir79T034
ZOtkh5Cr6Am3/6Yxxl32fFxLjQxbTGHZru8sSMLAh6+aYNcdK5D/9almICXa6bya
vqB7uMiRLbAWrYpAzygNypIkBz31yn2nNkGDvUBinQb7F5Ym6vnPFQTMeAmalsQS
Te0Wcyf/QA3X1umegTpWXf5HMWXDv0SQlPmMPKUDmu1ukhTGd/v7l4M+pVYxEzoN
JAn+/zNz70iZw2CjzdxDfbFUvPUYaztqCy2X6zrgx472Esh+iXOOTJm/izBortkX
swy7SJjHQ4UPwPY9WKpqzQfBlUwT/6Ttf2hP8xnNRqfm/ZdK2A0lxjHNhYeKVTR8
067Onjz3vsdtx9kPQEmg3Ao80Y5Vy8tyX4swwlyg0Ye8Pqy/JsLZuW7qOpYabFM+
2CgKC6TwsWSMloa7hGqpB0fDT01XBDAJMc0TQprVdlkCpTAJQ6Oq4n2MIQtxdzY+
pW2MWQh0NYJ3iO+dEo7OeK+ACjUYJAaOjgb2h0Qhlk2OvZVqHY4EHqdVJjqw6EIR
juOru8D/a52q5HTIkyukqCqxNGresDCIW0+7W9LczTA6zvTOB3lgPk4sZpbpUUpZ
rIfPt//WNdCx/u8Br4WMU+Lt9b91ct20Yq65LsF0iDk+jMIirz8a+6mn/CKf2gk2
GThY0Km8Iw6ylL5Pbt1kLb/OmTcanxZtypxG8O1qZCypjDZBOMtz4oxTviOgrV8d
3pJyNa/WaeA8BKiqhkPx36ZG+Z+xUAY3/7KvUx48Yz+dTpTxkno4vLj2RcQi7Oe4
rcc+zfRo1iNHY/+LrC7GLk1XlosybdiRAmSaBD+cg6/tomIS1+Iglk/hcLze5O8K
NmSQUzbLd75eyK7mJzq3yMcEqWvRnORQ7PTuKUC1ZStWeJHDFXcmf1bM1mp9wOlN
AxQbsoI2plxMLKGPYkq+a0Uin1SKecuVQclV2ErcSmGFYx/L2AfSI2BcVw0EhS1s
/UvYF+eL+A4DYClaZYdsMxFZTnbz/vCf9//jfYVAHpf8HCSLU/cIBXUM/x/ypK5B
7auyD4RAcbpfQTYm+7n8155NxEBUkjG7xhC4HiffsN4Zxh6TG6iUmBozMA3ZNjy1
kIWp4omEZ6FbZ+HFhHt702Y3IICRCSU031358AbHiucn/d+Sd9WL6W2QyoT+G4ul
lZwEmWf7cO2bWAzmfSEs3S+JsH5adNTo/Jw/+3UHM4DhNllyM9+TSEpO6glfTtX4
R/seUpPya+uvRhgqKEMU3Kb+QYIu78CtpNg8SmGWY18rxTLLbuzFcIrA7FRaYL+B
GdtyZsPQkUBsiYRS/9EuTtvAhhdcgrCshkB2tJV+L/ggVMohLndqlPUDPeORRMW1
ONW76+OM81M0gK3v4CJVjRsLnwFC5djmJp8b9wceywlVfoibsQ3C+dcO8YCsYYs0
8yWoIPgGHbwZer22Zs4Yy0zyUteoFx2dG1Ey+V1hKW7SSzkvqAZp0w25S6VFE7ho
HjM1bNKcuEiTZ+3EgsCduv7i6z60uN8SHnnYBl/34w1aInXlCLTI8ene6ltBcDyv
HAsB2OetV1IDb2e1GvUbBIuwSu+Rrjbtk13nZ105a8z9FjSqxgjVx3nHlFlceUwa
Wa+kc6uBtsq1j9jCVrcVyF2joOwZNOPDbZvi2Q6noCzrbUyVtfet/4BZa6M03NIt
ngxvny1g9yw5UegyUYr0QHUgZQP/8f5ToyCnU4ppGm4vEmiZWhlmzXjo6xqlIt2n
GL57IzZQFpNEaXZ5HHPtg2N0s4NcaAFIvdj7jaPIqHxR7e36XqPh6JEF4J8r0nFb
/fGL1c6Qb7nA+FKhPHoD2iL27yiyH7LgvUTqZTolsmRcJAx5r1VbDwENwuWMYD2C
iZw2FOKMy/gKRr62ge5XhKSrgtwsGJRp4CXp75VeOnCNuRamKuSyzraJ2o0/mPmT
zfOMGFVVUKJ6pc29svXP3rIdpiewk+FTMjRPRemAnERnnZeKWAjQadRFpI+aDXmH
bMElve6acfgYKOnukx5FRoJ/xbqC33zygbuXvAUK52KEJ9viJiy8vOM4hPaW8tHo
zK1iA0pqEYA4s+R+jW+0ix5CbrTTRNdeof4ieW879jME29QN3LhxANEg3dWzNbot
PGWSGTgISm8VS59NO89Lg5qLKkDfWqX1tNEvNiiZlhdbOeXdVsxLhHlJI5b3ZiSU
7OE9gQuV9FSm+UTUaMkPIlyUxVvDZ+9T3mamsEAwGKlrXeBQsU9WuM+ffQiVxf5Y
izQs/kOOMDbKtlwsZjCxmwIsdyk/IVVQVV4XAWQ5m/g64lEuzlH7RtyV/MmsfAaW
Cu8jmw0bULqjIVEIWl6lzZXWcfAiziz570MMmt0FWegKw8dV1JkcAm4OuUu7uV4J
eRaWCgtx7LshsbDCP90zovLhRz0xGKsuvcE56hMtOCjvHbSmkibtNJppXTLU6Em9
/rBWWrgJ+VaUKpOKxdKJYNmbtgCH+cc1VXvlinipMFXNzhCRmxXIpMiQCl5DHbeP
wm8ngexkQCKSbJ4xmDarXkOSEL09/23DroAIkdN26U40DvKE1TQOdpVDGjFw1SSC
iZvGehOo43Ob9bZaa8PlbfYjtNgygcSbG2Dq7xc5d01F21CN/0rVA6E9rtwAP8/x
d+6xaZGRkSaBMAQyi8BEnQ2kNLDWxtjzsVU+ubF+vlY7cyl80gBLf68KDDrPzRiP
FxktedAfwAL5dZB+QWbl61hn3YVYqw77fDXVgkaCa/K3kEg7lwBJIEYs6The701m
mPyezhtUcptpy/wSWgYNI/e+ewh47YcvWpsvz1qU3XFFdQLuZE71fKEDCJrLlrnB
vo4KfIwCOi+PTehRbk3xqpIapuZCo6aLtVbgeH5xFclgChx/GkMhz1YqowbSAyZ0
6oJb+PmECLVFdXmFPKAc7ibjPfYb4aYOhuMIdAdC8va4E3NwAnagODAyjU0Rozi8
CD4+U/3uJp49I0Vl1b71/djmVhBQYi2RbHHmBw22fQtYCQ6S5xYJkP4noY0Ysjnd
P6c2NvHj+1aN16IDIgz0cK8eDOpqrpTWB7aEldVafzZ1gm6dZEoQ3zTM5PSo1eyJ
+yG4pm/EzCkDWLvXN6xes8x502QxmvLrBH7S+NM0acBCL3Pttr2nYQOgadpIi+su
H/w5HRt3O/KMsE1BanTL5PObCSgDgOdrzJ/iO/cTbtxyuALw1ffgDt7wjF2YizWQ
wOs/BfXC/PlHdcRTdQJpR/DO9bnqIXx7+rWYMo13CIWceBeTqAK8Kb8eUrz16Lx9
X3DyFZFezVoBT2tCjfImdSRfV8R8pANrcAi0+wkuKg3BvZAJSk76qwEMljp4w/3U
6ihHQKTOnYdThSppBPi8T1j7367c4TOG5j1nLgbOpAkCmFjQrt8p4XafnBGUUlxt
2zd/20V8Y/xcG10EMDa79E3unrs4bLpW6T/rB5NiDe/yTaiqoC3iY8M+577P6ZRV
XERhRqMK67uvEWsmFvwbOKab4S2zItHU0iqryWO8O5g/mLsrWDLG0OJoxP9eMEyY
eoSq2DQ+frd5bdAG4CdRjPpOPcuZ69ZQhM9g/jxtNmBafzXNXq71HnZHozfZFkIX
g/2y2z66h3lth2r2C18ot5XzS/zAY805QWCGIsYBpli8ZKR3jKFKbu5/3LMN7Qj2
UEXPB6Xw55pGb79AYhrTNspmLWm+TESl5F02ApaylvCu2WeC/T06DvN8iBIpcn/w
nKCelu4/+ILBnlnk6EbSQ0AoOcK5HLw+qllkch9WXbhP1NSJ4PbuFz2nAori6t7m
qvQzvsSYuLhkRrZnkc/ezp8UKPTDjKbvIfDhwOzRUlDOaV0x4iYz4I3XP/Ch78Jm
X6aXI5ZZShXy4tKqrDSqqT1ggwhFyndVoF9YeAd3xzZW51tiOJ7PAGaq7NxcdjEG
g0hNJS+lzhE/E0Fnsqdwvqbm0w5+JkiuLPZynPpM8zXlfVHhpovsl0wpNK8CGS9T
KqSSFqVRyIwpe7Kqc55l+YcvJRJVXreiV/IKKCNp8FIfqtfHjjaF7fm3A+mH5c8T
zHcOp9hNUThi94x9+aXdOwSeTyzZ6UCU1GT4oZDHuJYx2KwbZJL0lD9hbVd5xzpV
E/00QN4MT+Bq6wo5YoBgwd8vgxfWNetF5/sf0tjRZSqAV2fhJ4qcEv+5Hma7qOfs
nTzWpSTAWlstBrcyjTAoCe1haaz81n2HG06uHmEVihO5GIF5+4SWQon1bcqeN4yN
uvQB8qdatLFh9KD75jOLo9nPtxyNZc8jG+TFxch+bXdgI7yPoFp2ced7f6ttjdJ6
OIuE5ISEnNuBn1ETlmzHWIhjHLVUkhIwteBFhEripegyyeHEtoXJRKlU1ZqdB5fX
1vrMxNtfvQPkuTl1bjHkrPvU2zmDtek1gbb4QWHwzxduHZB46blTpH0ILdWO0sHQ
yBVrnLwe13wXXZgRLLUfaXguC6RN1oa0SFSoPimWO1KRN822IlNFZPhHU9NPWyEl
nYUTpumnkvQxsdrf3I5BR6qwM8NkYhWxu9WRNlCE+k7lAQO0/pBBck0UIaxQr4Xa
kJ332zFKmDVsyJlnuHpXms82/RHr785QwXIYpVMbhs9eYTvTOYsHm1lBcYgU1VxO
iwkH4MUJY73VnRA9cqIAlVg6AKh9b2xKzhrE7CCXCCrB9rupEEivuNJyhFMaLcmc
gHI6TTRi3Ej8aBZIDozGVrOrHE+q2UrhEp1Dn9g967O2FLUR3KnLEzA0rbh78mpI
a4BtHC2YLM0QbwptbIpYgJUDoWnpeDanbGvvjFEKH4Gr8VU4NHi6jF/uaFHl+EZ5
GUlmy3QB1ZE9CbJXC/kT+Kr+GLYA7UqlCOKIaIWO/UMAU8/osv2hzjsJ69np7yLL
RS05EdGFTMuGV/H1n0bt6C+2g/VVJN1IPKi9d0UHwHEJbPmr3gzNQAf5KprDunV6
64N/Kle7wU2aV49gkgyrIPo5jd5GMBb01Y4vt9WoWuOI84dBxI2YwOp3hFTu1u3E
nbSSuD1RkenX5+A8U2z0doxRyzn50MBBjH6PrVfKbgQuhSQMjCp5JhsPSH4EcZlQ
4m+QeFxS5Zn4iZOkZWHGN8lWKVULBRatkPb9HAmkD/zRr4v1ZJ7XyOz4lCh5omEC
h1qWs0YMXRuQ1rvnH3kRskzJR2rCZjafhrlcN2yFW7WjrV1oEW8QpVAvYPxSmrdt
QKa1mpa5APB+jyz9c//3thqb6prRYyN/lcp1GHVbABSgP5SsfrNcfLI+RaMwYKv8
zEk1uf8Xy6LVwPl/2J1P6QwWdj0fe+2IZV43Q/i+++aoT5owkgGk3PJJvQR+0Lts
z1VENFZzU9YXUCcacHyU69Eh6yMQJA4nrMooxjbSdqkEDBUQSNhqLG1GxuFvfoqm
mkuaD4X6uFnZwGNxHA7jYEQG5ipAwXcKKG1FCt6cS1YrQWFrBmzdpq16/bVlT6aS
8EZbYMzPoDN44GaoHqDn7Qk2IZdfQ9mUyNvP/pBMr7Sd1a6bE1bbdbyDEWMpMPgC
rM2Fgt7PcGaY5qyuW8jp6iDgzE7h1Bq4l36Q6J3O1C57OIkqkPNJzWKoHujf9YTu
rvyvtDONpcfGyd7ebGWdhev/ZZzVg1YYrMFF45kmc8xlzigFliUIxE3K1gpUIgIH
NfgF8ctULnktwTEU9SrS8L3mZAvj+x7tn6dDyni5SOK2A4Wbbm5OOZ23FnfZvegJ
5khAqII/a+Zt08JGmwP+vNXra9rb4SqZmAhjNRj84xYW+5KYJo1sZA9mgi1Vu9Ev
EwaO8hMgsCYeK6TDMM/lYg6k4I1Nu0z3X7Btxz5NI0jM0/qXVdXBNb8yx57QNR9d
YJtJlSLK6q6xIvyybMiy3okwhKq3Jmz+a3VKQFQhxLQvynAsLz8eT7s3tm5P4F9c
1xLDLSLz+UJT0DjqJu8fBCFgZu/VBO1k8BJv5AQ/2mqek2V5u223N0HFdOhcsmTx
+YWgiKWGBCStQ5Q2+7m6scBw4kBSB3nCVDpeG0V/gMVS/c14kJfzIK9kAq0J0kyB
oLana5DasbSi8e3Z4Xp3WAwKgXE4ZaSnuU32pqVBO8ewGrflfDwrtdwKJzQ8RVZr
5hFXlymGdS5uFzXjuV9gjeR8PRtub/u+HUEtJZQLMTWRNsmR8U0Leax0rma+2/8/
AaEZW0Tx7v3BFn2vphnA5mXW2ZN+CA8IJbCOg9bMTX+XFemZGviGJq2CBKarCcZi
capkO/vPW3dsJ0/iPgmPN5uCMRqto0tUB/Gz+T3rjDRCyfEIEFfWrT4gTvSmuN1y
gGN9yrZLYY270eKuDSXOBv0b5GQQmlyIvtpkJL4FKJu9zECsOkwDrBYvneDqrCSt
jN1YwYd9Yn+PlJAFpydgIl8cCe52gECO4/hMmmmxaVgirYpgDSDJXu1PPUGbdsxO
ZznLlx/EKyBiSQl98anQrlIZQOv7dSZTztIb4gdlH+6m9CT/8jLGH31eBBvJx3qg
lrN8OPmyGdKsIsb6iqMd0fg8hVfDh+c9Eb3pZx7qVbm5l2zNv3PbZ3zGrjxMdfyr
Ov2N6qGL25D32Naj5LnPI2lQoKVuZl7VAv2lq5q/si2TxF23DVDIVhUqPRrIux2D
lJTYBidQdnBvV1IaaKIc89lwdGqPHdUj/cgVFo+TBt0JjLM4UZ807Zb5eaPKoila
H+azW5+/PlBtGBOh69bIOPJWiVyVfbYZ+1DXOqbgTFTJrjNyzzsbUi9XZrLiUO4C
5NlzTDw9GPK97ggY0acBxV6uqsnCRYj/4zBIAev/h4Y70zpvG91/A+6atz+yFmfM
/qfUV3nAqTXgbCz4UF9BfRjMz8zCvbgph4aojMGettOI6ChFe+RYVYLTUhsrsHO2
YU7YNJFqq0o/Pk15UuiLmdaUIcwVb3qBMWz6z9D5CJRrhpDCDTe2IAMvIFq3jAqu
ZfQhu227q/ZBSBy5+/XoR3KsR0rlyMRs9k/Il3KqE9CBD7nwk6hloqUiqWLSxmET
akApJPPQLNqhVQkqlibSmvEh+HjrDUZYh3GBxZrKtCcFwYunuoYJzjeo4avmyUA6
bktbfcVbrfcdqL3Lt1U7p9mTzADJv09/rWXQfSMi3nKzGYVwX1UOi3UctNrqWtRl
tVyyyIHZXosgIxdxtJ6oHN9izMZfQlRENPySwlO/DmyJkqUYO1HqWkuVUtr5WjJI
27u+qPCRBRlEhNPi8GVok8zqGV/CDjZCZ7JbpcV8xBV8WDTGpLkdb0y+dSSjgDY0
j2YpKfCWZ5rkmN306X/5j66IAxuHCr6J3eZ2QmB4UfxV4XBbjMiESAw4pCj1qJ/P
Ovkw33SYVQq1AkPwiZ0Ef8A/lbWCOFP3a5ZGeifo54nNFISICAgBuLjyhsJgTNJc
Qqv+wKvZm8Z53YZCDN7VOsdW7nQHMFoA8h8uA0mqkDLl42SYr9Jqn960oANF/kad
e5ryUsgEjyrpp3heLWpUCXMLzFBya2YbbMlFTxk6ZLJJqkCf1INaonEB4LfXf45e
UnwOAvQWjwrEtw6xNHIrOd/7RcJBDyK6fOHHRG56xXjo76OiCd8clE9fNAVYTcs6
cgqT3fHyLQL6Ek02Xr38lnb31hYrrqzOcttV9Q2yoBstjodiq32obSOJoQATZCac
nOJf1UFl3OsoZMjmfOZO2udOGVgtz5qO2OWfQ2JwTtEpZWukydKa6T2+grkpkaYA
z0p+CZbvNfcW3QxLNq4jsFxVUwKXw43WceWG/NPhKeLxu6CnIwmc/coVl0bXdGN1
afV26BwVXbNIGsfmQeZYl6d2jSTLN6X+H+YP+DndUgEPfmcYG9Iz5Eva1Vd7lgua
v+Qb9/XrCIX/VzEFm+Wz0JmQdvpiivxqVH+AzdTrPPolN4oEazZ9GaKYD84uQXO2
XaBiHx5NoPY6gkm6MDCnY8JGmz/qJPUrJiderAvFeN9bbBJM5GpiwUvwiXtPYbvl
IAgWvSo8gTXW0B7bnyoDfDBScTLqlO9PHXmc29KYCtniROUcccuxuJr+KrUfKlVj
X+R2UfCpHIYhSXqC92KSj+gSmdqfcBAkof+qUMl3pNwyxlPLM+NOG7TuyhZu42gM
Q3oeNHPlkKE8UrYDbECk3VBqTaHyGq/IA+F2ArOY74a4hYFHO77CPVzn32/6EJOz
U9qn4fAH9XkPB/nbK+eXAqBtDivBvrL0Svd55gKYJhBZ5v7INr4Ji/uRRDEC/X11
ZPyNptnsMf+i9bkflhQlbIBZkfSd+qWd/G9xT3xOb0CjWLV/rTQuwMJb9s39LR9X
1SopEdhDzeKxiayTkoyEDiZVTxYU+W5z0Zw1BZCaKzJa/KZUgpzYlSCW/LspbrbD
S6JfFZOAHPsBYCwwjy0Ny+pwUMq5JELVxKYA667WaaaMfFW0CL2MO+O2J1YsbSu1
XmG9VtusSYgS/neZY1Mx9hxhtaqQ+CixRrmLG2whBqvDR6V95PzdTgyZsErPFGG8
GNKF1wNponJUepAoH4U01MyA3OgXEl0Pr7ziEnkXe1yVDzQa7FydeZyHaK5jISkj
Q4SNiwhSVzaqfVCirISDC4QVW8WiC59ueSekhC54leF+AKY7hCLfXYxJiyK1bPla
1GCtgphwY/b0rXxEMLdTwcNhQG295/8zFwoYAKoKz38nRWpJL5axTRRMGunU/aSo
V6o5TDQrqaCWgoRDx3Z9Ew/dcb1diY/cIORWG0h94WNGS6Vw4hNnz1/fcp3frZak
fUe3hKGpb+8SPDzDTVWm1HXdaJDoAS+zz8iRAiF33Amue0GQte0yWJyjMvEKYRq0
AUWdyKj3TB6ygEjXJBB9Yzq6i6af6/diRgzlUxW97XBWPHlldUNuCVw63pQ2ZCw5
ko5rpozbOtHITF5wyIWtDCt+/lVwto+L+DIMEAtNIYrRSSwspiQLwrrZxAkg6hPq
zUOtrcAM48jfQ/7dx4cdjwSI5YKAFiayFF54I2qkOl+TDYNnHR78IWucyV/BzS63
13MMa+8Tly6cNvuiZTtrDvEhKckPyiDx+sBDnlRK/zpReLlzzeekxE7IANgGE96G
BZzeH2f91g7x97vOhM3+2OqTduQS4MzmwZPIdddWNN4LURf8nQ7qRIBdfn8j4dYT
DgtTPVW7Pbki4pGzlLL9UC5wKEKQrTdO67A8Q93i2Ljjeio4uZlxtF+4fuKaomsH
hw26YO7ZZ1iRrOprOoGlb6G4IAABa395dFIIRWFdLbRi2qBqvxXaiRnPux4ApuBC
+huUZkV4asRDqc3zkWXrP2rPfORWkeMXFSsilNCKAyyXftIAbfyvIFiX9An9zhdD
2CeVZBB9IToQECqwj2kr7DeSQppH23/PX83znpsY/iece2ZIBBSoVXtEjJ0CSJRL
dUr1UdCW8E4vvWD3PBIl2V9YxxSOOts9feAX62eJavyOW4zVcobbNHlmP3EW1wED
Akc7ltz+eweCh6q+ryqCbxMYo4WmKs7Vb5cjO4N9/t+4ZxHYHWJ7bcnsTUYMr7CU
aVjA2Qf8AmHJTHdezNC7/FnX9ZJUf6mWKyBahtOTBHKBKUyXeEmdgE7D6NoSFyxM
WIGY3ifcseDvEt0cxnobU/zROE9VlzZ99/J2wNHLqiZUfCtuG4ACLkkgvxgM/OAI
NRZRcXrdUhnaaixGRHBiFT0b8vyh19eUOO3VChOdiLYJCDDJQwXllYJPbhxpmXf+
Hzxu6ipCPE6Kubs4GHHkMtRvQDuFdXujqGqigWFk6K0Q3TCjTwCc+TmlExdJL9dp
tLSZB0TdYElmP0xtdAzrJ7gDdwzcyv+/H6POQFBvNSBPcuFYdQDWRY11+MLD/487
G/JefdKmiifyzaLgehOS1KUEylw8mgRaMCVkL4mF/RLy0MzDmLtTBfy86ouLRTgO
EfptZR0uO8T6jGAKehoJjI4GaK+d2N67B9xx5diNPXy0sj1gTmjcY7OZqZvrLlmJ
G2eiE58jhSRcXbI+mMCsDil8eIHC+W6vRkKh0YjPVYQQuaVDZb1l0BWthnCvyLcz
eptEsgNDS+1myPgOHlYyAJTya+WNxeBnx9dnp/Vwbpa2qLmorG7jZkqXeM8smkvf
IRIMYamGwbPSlDsHlwY70r3BUDcnmtGTT3JuXODQAUqCRC7zFknTNeyY1usGd1Xg
OQ35w8QBSIx/RqEqQpkxWYBHcOJ52UkjJn0r90JBxt1dvsoI9yl8U8QC7rvRt8WW
L9uJhVsTaVrqNqi2mj6KDqeLJXdNSI9pR1AUYZQ/kdSf+2OZ3OeMSHjGhqUi8zK8
StOSYkfIQ+xnwFts7Ijh82YLwJSDEKev3UqQK5VfSRm7KIXBPXHYFnptcLdvv+Zx
hCGwHpmKFiZ1hj3REn1TqsL2Rqv2c0AYQM89SoiXlWIvqWJfEey/jAxPBOrDM7vo
+1arxVfG2Xw65rw2GLB7OAC36xNdpFh/DOo2tbCbPUAtdQWS2RdcfnkJZH+XSD4Y
hQME0Y92wvE/x1x4mxEglbiD3hKZdduhHjoJdksTZtV9hB1aVDEDxAu5udTe6+Oq
UjB1U+GkA2ksQqSsRX+7nrj+b5MYpy6cUvzcwwaIEIIIFBmkP6A0F8KwQ8FGUk4F
VwRka+oYM08JYxh+v51wDMEXlyoaTcr4MGf0U9wOyUz+8l6srALYND7sH5MPonr4
EOD9WRAfYoUrwxy74PVbVOoF3pGgS+8OlRYupUiOBVS/1Lu3OdtADQMJwAgMDNmX
h0pv2y5N7qr4rwbAccD7S05934cng95GidCvYXyP/qH56yCBOzxf2KBizhjvC4xr
zeYj08y4HUaR0Wiekx+Pw8HobffsXZfFI4c5pD502I/sMKeExRRav+vR/MWYj1tT
afFj5ISwZHnd2ZBvoNgtbfVZsHEnU/YxeygLJahJvRXGHNYEBQaKqIDyPKWVorNl
wslyyGcS5GEmSQmA6pYTKyI7SLnS0iriwIzGqotAAmmBVugloMovSgxk2SkUSgMD
9byaBdxfqtbu+esqF8mSUo3pYrRHcrTSbOBRpsL5RqyTN5oKoWUG7zG1dBpIELTi
xx/3Yzk9KoIbD4PfxV3Ft/sU/mAZghjVZW91y3QmIHCKxLRjkb8OZPAcpbw9BEqo
KjDVi5SsJapG0xcavK1MB+J88pLD0aB4rixAM6Onjybjy9HPNmy/mQJF1GN7j04w
M4TdRkQ4wa0tePlxYNjpkdJQGvF0IAbmxgSFpW1GpyS8MuPip/XF2TaTOzqO/Gh+
Ab2QvcZb+RqoGPNINyRNfZLkXeRb1aiRVPq+OW+CqaCqxot2Jf7MlZXzqceTULEx
n4WvHtGu72jtNCVdsX8WwsVlRe4A5J3ZbU/h+HE312qiJ80Hrpw87UFBlDNChbrp
PW1uLNc6gR3apyX6IZ0kVN6eMRCEteygO2t+/RKoC/WKHeQKbwca2cImWOX+Mg8E
wIwG4UyCaT05Zb7vO5ImnLqwkYIU6Lr0OpiC4mgnyqjZT9+upurNpZbdXipvy9ho
OVcdMKaLuHZ47gWn73guVw4j+NxLG26fFvcB9l9oVZKx1CUO6yRfNK6vAJ7xSqwO
dzJIY/zO2wWl4xW7BNeK4V04+HBAP1DcCmjyT82EpVUiXZ84/B+1sqxYjomkFEv7
BZeR+ix3q/k0c8+Q9LzysjByDlA3reVyitpjEc+pgpe9SxgsVfEzD0ySd3Ek8m0e
Irl1U2HmmVTwcmzoTB2mwISeT05GYiicWv1Ia0Qx353bRHE3ii9+VN0PbllpmVFj
kQgT0hIkbTZ30i7qBBQ72ALe87rmkPlGdF+ue5iUvHfiB4Ghh7tEDJAjvi04qyXl
xCL8vUZXprA1sCVbRKsSKsauF5dQFRVm0aAJN4XcIIgzzKGS+Fk2OL8NseXLtJTA
699xw4OTDlOp4t8yyxv+1rnN7VIUDbLer+ckzd9sbbM1tHJykAEWMXgTQL8Y1XJK
KMdXVQmKDsNtCwN9mJ2i8pkO5sh1Xrw5iNJtU3iFDbeA9uOm2Rh3pByJPvlisp/T
9fOd8QtA+c87vKzAYsRUJ6usRKDJ5hoeC2e8Y949zdoVmAV3zJgRzQpsrT110w7C
Nbw4be8nWf2y6Uiv/xsaJT0aCV1s+lZ3iZyHHzN6r5vbnNmI/LO5tw17j1DF7W+a
PHIfjYxYsmu4CSualae1DN2F5AiD8jLuQXA+2oFin7sq540m+/fyRpvoVOyZ+Hp6
VBx5TSNLqbf/mLMqIvNSwEWd/xJTIcNA7Z0MLBPrU7HpeQzOzi1W10cTkLwfbPC6
wJ1BsoXeldg2f/yZbQPLVqRRkpCmPtAHOgN4DC5x1HlYFr32jwr3Ur6/aEbAM5Lr
nd8p8LHwVX1jZw6bXelcgO2eJVwrnGtvYtu3WK7MjR4S8u/+wgCzMXuyps9ADNGm
Sd7zEv/FjdpMFPD1eR0ulnqdseXKKAdnxq6N7bZbnANnSmYcsh61S269sO6xehJN
DpyfZC1ipMMD50l5LAWroer5u8kXmz3ar/NRJ0feEQjHKK64noTm2UGIJ/FnkNHB
AhTC2ePdHPOij2uBgn2U72DUQIYpV6x/yuW2gewgN8nADyn7zJNfnfXBiBXE/pEI
dSYYcqVdWj6SPOtACQsMY3HIiFNcMALXpJ0kPE3U6AZERaKJ45jr5HoPP0RZhfTb
92LtPSh60OJjG7GutF+USlhMKx2dsHiZlyvsjZKcHSjMMyg8U8fJZm1ake6+8pnB
8FJkzeQh79KgyzNu+Vq4maBiRcBDNkFARrw768nIznGuJekwWx7fy9ISDeAfk8xu
+yhZZ3/nSxb1ma/7sbE/Iexc5TO2epwoW7mWKqeNQbu1rv+eQtRE7wxMn+6YibAL
SnVSxXwT1xqAVNEbdrxDRew4FMYoU5sbCAZh2Q/A6t2yhKD0ElhtXrpqVKr79zWN
HPdsi69US0evsxomS0RQLM+5uYpfAsqsC79WRRsHtJMHmCVBGHLFnFfUjz1GfYMO
aXSk1NqsC46wUw5kGYCqFhtZVcKiS0YT3AwDCs8+s3l8r4spmOOsiHS5cmDd+6xx
2owWbANtcwEAi34e5mzoDWWAZu/LxoOKdDcN97dpP5fIImiWGpcrU3NVWKYDukyG
gT3gC0Eo5vejQEyh8sQ2oAr4Gs7qfitDN1F867SDYC03PZVNm4H7FKp5owIHc5lx
pjCzyz9Sb9cT0IlS2v4eacWNcgD5Tu4pbHkNW4QyXTavDDaApH6rCxp9SftvCu8h
RROUPH+ynwA9bAnGwYRTR0aY406dZQ9ofwIJ6NGr6cogaoMcACuXEymyU7rDoz6h
1014fGpOHj5p3hn3s6Jsaygq4e2CMwVUzcBL5Sonm+ydf7CbjKEjskobhDdk0tDV
3BIREiUHkk8PqDynHy7qlVkf72zBYsA1QKzGwLPPSv0WPTP579KgOvf2BeBBnjJc
EZ5XOvJZ1IrR8JDC2AT37yhTk4VekF3qFcfYvu2h/8uoKvrCJc+NwoEAiGPImyCc
rn8/BRVxOZxIpholUxpxWsMxjer3jWNwGT+JAOGUtA4psanIDM0uqgVS4SU4D84m
Op1aNGizQLhHqsKgXowMxrUfXe/M+c25ktLjIo8Og/Yve5iOP9I29rH3kNav3TDN
j9rXmcPzKUJE7NaTEfR7N40a9pIZhLiSfU3CqIUbLtfSLfWJGGpuC02B1tVUxUz8
CyDJq0781R3rH3m95JjACSQZgCLgx5+Avyo9WeHEOMH5/Z4a0ivzlNdWqT39R9pW
JyJYGTkB+BSK2OslDIuq9gCUZuxAYKTyNeOxhrKuCdVpmCWr3Wa2drmhcmFQC7m8
0Qss5m+m9TNXHDVzPSWhDPZl7zqW9T+P7ugvAfniBa1ATBsbiEftjqNfvinr1wyY
HlfFxVFquJ7IBsItM0lol1AiCldATIad6T67VK2QUynjZRQiOoodPzTEsLrToWHL
Tce09mvqWpWDaJn5e6tvlcix3XpVTtecYXYteOkU2APBOOn9Si0rxQsIyiOr/6lR
Nl+Tivs55mC8nXkH+eON22SfFY62qKMS2QCoAdh0XXThMlSQZFUlCkcXpQIxJ++8
rRVitloNl25NcczGEvq6P5Rod2lOiKnzDhJb/sowLDKqq+wz+GLm8wkG8eChbi7Y
bx2fw+qWpCAYkcDacjjw7ZAVoYB4c6eGRpnHHx/izHds21fMcajhtAuBdDCNxYhm
QblytcYnMgWJzTvBIK4C7H+mhLGwmbs9Zwqm15q5MJvdrg5eFZtZxwRdcnsBI4Mv
aDnBZ0Reij3/eXwUf+iQsVJkiuKmXcJJqQUggePezGXNkgjpJttltJlMPsdbmSsD
0cvaxJZW37dOdm/TUdCKrmCISNLbSlLSyOTFxTig3bOFRfyPHUeTIOnzNSlOS4SD
Pb6DkhNIrgisW5RhcXQoCivqaov1zlaAVQq41/3RKH/iOSMXzxKYY5ghjgLcOIFD
QFKZSeDPSTjXr8nfdq/FbWk3PiCIHwZMEcgNLADJ9mRGSPVaIZKqPVlScRLeJki2
Kp/ZDQwYg2N44/WP1UI0MZeQl8CudsEoVFdudhMDQbX65yZetLYmM3MQTf4qwi13
lRv9SX0YnQx0KrUIMfj8iy/F45augO9cFKxomuNa9dFVPPx37RGCkLoK4MpDxg4G
ou51mwVX+jubzBBotA3Ut5yzN774yyEJIA+9TinQvCdhnXa40TTvDYhN4ogEtoaM
k//UXhaPHJJM+8BOK3g3RHmqEmTtJpkxs02ijklLxj4sMP3Hv+N9dtVeApi93TzJ
Jx2WoMjlXtdMWUY5EDGy5o91cMrJXljyfQK4swY2LgDh2w4Pu/UGSzF+6KiRZJo7
oIVbVvvCtK6QeEATPFPmQCSgBnl6sPToW5tG07rA0/BQtme9CLQFDdHwkQ8nsev4
lFk26KsdcdAwe1UYsIaEslmc2T77FVlOY6dkLcw4RkHQY24gtam5asRbDcuSD/rb
wsSYuanWX30RCiTXyH7D+s+H4DBdGHMlabayouGSE4FIh16z/b5jiha9KyLSdEQY
q2wK+BhE9Z/BHoPdztrlN++h74btSgc3gIu8oYTPiAOgUfu1LYu7PO+8iU3VrgAG
1dIgpsAUZicJE6Hwra1nXgYcw6N3/Zip/Yv05Fzels4bXdvI2fmeKQXAeHonh+od
lqOJPIuXwS496CvNG85C5dGtCUodQ+90W3sAgmJobDR0z502RUPUiF7OBJbSVS/D
TdaCrMj6zrN18YDER3+DPgbbD6JhrCQHUHRYmQ/ziehbnZsoCg3Vw3eHqtMukMRo
vZliMldT5+vXVehvTuiXlN4SXzRtou36AJJwehGYgTZizPe6KtMyuup3PTIRfgkx
X+c1i3wid0YKljS8DaTmRcPe/cqdcWalvAeWbvkHMgZDAmXXF1KmIjXATmzxAT6d
tMJ2y3VGJb3bxeODX+AG3rvvHGWYlTVplrJ6uXYppH4GLF36CdUIoHRH8jm6ggA+
JD+Rnb3xFNfDoCdzVNKiKiXBACYfmz47WpeCYJYaVxmS1ThcmyjzoRMwsYQnaiJf
6jVKU7NKaLynWmos3RlGwVh58LR7artYEY2QH3OzcVWuVHTfp8yv2m+US6FuEkbq
0LP8qOpdrUFIq3/RRrNRcs3R8KZqK/fnU+iWxGCx2tiQ+BEIiSYgMAxvbwChzMcz
mTMp8F6NpRhGMpPgd2igXAKTRAv8xsKIZ1TUowUIrLT6lYI4zDEG0nPQucNe8fe/
nYAM8Q6axvtA1ZwzSK9OrIBQFvi74QSRajyJhn13rIrn7t2K4YR9yfk707Apmkwc
lyIRNGUWgHfCKftZTx0UyQa84+WcYdohQ0Pchfa4+VW/0g3mIkOAomvTqScXP3qb
86ULuCoBLmVy0A9zDWKyE/lIXIsapImS5syyWtHI6QOa3JZIOIK55U99Vq90Fjfa
R/9aTSHTt0hA+yRK4BApN8Ai4agaZ/e1Il+PrPyo7J8GBs0lP6LkqaYbhwzxnDdS
967N/x5EN+p0PRzau09LRzQtS94UZhAhgsyT2FKxLrCDMs6BF/LVZbEWWah4bkAT
H1w8+InxcT1NGXhR8mkTNlz0kHdEwGh0z/aqBLausgt+1Bdrh0LGDVAq2yPpatS6
hqElb3wXC4DPCIQ+/g7DFRGVbpDrttAd+qbruHC5cHymPA1GuJeeWGywyqUdYg5T
pL5LyV9C1kdvPHHMT7uqG38bgLgvKDBuI4IITgfEcgOxOgWhDgtbDQt3QCoRzdwB
KNbEHb6k20LQwx5xWWF+fkUH9kIDXowEus4i+1aHPO0/4kta6Hm2ULHAuH7n4Nxb
1C/jIT0rpbU55JSR0BRFlsdzpZQMb0Ag1F77DxM21sOBmw41mLnemA/5UsBMscyF
qrOYcn+qUrUBMWNSFAu09ZdRgU1fjoByZ7mVOQmpoWGo68LYRBOSbkr2uvOq/reS
qEJg1ONx/T+pA2T9jL+EJZ3CTGJqXkCrcket3YRtmS5CjLOJuvcCauFyv04HZG5j
Ge9DmPnAk4SwCf+0Z7xu6NyLdyxxh1NkWqS/csNxMmTg8xzZKxwIesW8he0M4D3Y
NAFOVjDhhWltPy7gbQ3+e41a9JqTY3+sg4QwiuS+Koc6P4B0XRa7zQ8TdRJocZPF
0Lgz72J6ZIw2Zeju8cMX4BVo6uc5gq7KjovCSn0ziTU3BB+RnKUBVySROl9LUc5C
rKX69qYBXFtLnGw49f2aPzaJDvoO1PMnetYjJer2OWolTZoTagk0A7FodShmAoww
DxrRwYWW2HNOC0+pfTxolmiztvJSOoyZ/vjxfqM+Dxiixofre/kYkGO9cK3DCqv9
A/LSti5TSss/J495hE09V2bFq7aWpH8oeX1ZoFUluHyulIzOwF00zW3BKWosV1WZ
bBrZTdlbbjFepOdlgPFOxhK3N1ut6CnlHL6d72A5r2vU2mRN9tne+UfEaJgvvRe5
2YyLdZy6e4vL/wBL84bxhMc+Jv9bZntRMbM3uPTWbzw+7kvaPzU+MUFvXhnZrqzf
hBGeVQTi60RwiXpj2eSU71DWIO08x6c5spkBtBZVTxgrIA8+D7o1nc3aNpb9klX4
VdsUTWoyeYdGDEbq8ffG/f+trWs2Ykezoc9M4cGWIYL21pj6p9nGZm1+KyNQ6LGh
8uIVeSJvtsbU0zBzSJ1b15D8qj//mt/JsiIXzOU3aE86ECbn7uw/rIAUtEE5QMMy
1VBEsF5tGT/Y8DoaD4nFppxjZ1evfc6JpLdRnaxv3AViX9UmqlR4/wgXPIr4GDt1
xXbN9DVHdhjGegRXDljec3riYi1TKb9rFZS5H32F0xZIF7n0N2qjXbrJQ0YOQrSH
q/SsAqIPftzoVsGOJpWQwXqXSie2gXPAKswa51oxa9cyPqrxxuC8gm+pUe47qGGF
u8keHLsrBUsbeuJBAWg7Nhp+6m9vbteYC9fqqwH/S6fJRq9Hy5lwvJDOxbW64GO8
Go3HOKksnS6IQ7+S6qvH7YSxK29Meghma5FyRTzJOzY2aT3pnHou4RixhOCxetic
nmyGF8kPZCpQ51m1v5Dcd3oPlFaOg8zSqatoF4PGKMkcNwVnhg2zLHase74dpHVS
MXbFC48Z5iuNdYlTQuy1kDXrpyIt4Jb4NNAQXyPy7bM64VLAz0BdVODynYCQC8Ie
5nuhxUTF/BCoG2YSQtXFcqqT+xtMCoMMWPC5lcUoUxiVHfVVQ0aE74SGeAecW+Yp
MQWxWu6glE5DD9w8qKXIaC9g5JgsfLYtp8pElkZ0TOcl15W54XhwLkNdU+MddhWK
5+rlKLsRIlgksGMnosKxVzCrz0TTG1LsEwdKkNK0Gz9IxltJ3BHZzoWC+wUn3mjF
fFxpNzqSJVcBjWsMLWxAr2J3R0S0ITPfMrb+8H4jwId4IeSnPOleU28rrtM17H6m
k3+e6+y2Tm2mjJemQj8b3Q6yqpk7VyebV75TAvDcwyNEvCuBvjxOgKjE0QkEMDSX
A1/7ych3qXjIunowmdfbwQ5Uj4+vXciY1kh/uasSE9xGXteTENNeE0OK1OK/WhhT
VDNJIa7woYHigqgQd0IziAcwZ8h6jAotbxkP0nQv4NJjBRX63CSAgrjhVVJj30Zw
yX+KnhkATRSZkyXyEvAi9BAp2CnIY7AvWZmiB1eGMY18LnKVwsJQdMv/BO/bpSCE
5/UQ/TAYFuVypytMqC4T9lg5xLbBD9N0mdOjUjj+u+zXFnlyVZIznJ+vd9/0JEpg
bBkff8rxuVsEbgegeAUt2QMERxTJtn3vgncBUWub+brZjyg/2mCRKU7Qr1nChaAR
0UbB5Z6/zHggJKiOvcD64BWU3hDkwpsTdPb2TTFkepqI8LKIl2xgWe83yWXyjq5B
QTRyqsfRIZnewg76SvFVrZrbx17KoRymaUKVNoJyQXTBZ8sQ/WvQOpx5H4X3S871
w2ZiJr7/rMOGamCEwGTYaDAN2yS1c9aBybGc0f3k3MVJ1n2fRLc0RNsyYaliVJN5
IVMy5C/mcgloCudyeL+DHhhfZWtiF+LOcZHF0h4KFLMip9JtcS0+zuAjfKqnI6ej
StrlvnjP4oWnp6J1+c5stSpK3j3NgQa0Umytvmaibo8cAeujT31aCK9bNoE9Tz6T
4DRJDCIJMLp2xcWn99DnYTEOCTtVaknPPiIEJ+/FuUmwCs/00MmsDiCIs6GKpR4X
q7LUBYLHDHN3NjX8VSY/GfpRBEQM4K/XaSxrtMrgFNSSfCzHQiuOXP+HzrDSxepN
henWSNhfn84epbko+blspn1Xh2I7QeAOVRSPd+2/gTqpnrBDZRp6sx8jFLKCwo4Z
FS8k9qSyrjm+ZT+LeHoQLvmFCDBVs48jCbKZRDUwYxQth8IU/yhO76ihw85S7nqd
dn3oRIAa9BhbzH3Fcjjrl0ifkU3QwqjNSKarQLx/2L6nzdywAAGYVJ/YGYKVwPkJ
8Date4UfMa8DExz/JUhVqp+ppMgNxzTRenie7BLg9fTz3vqKbUDzaRqxnA3yVBvb
sMXvtC/m4g7bIwlMtEkdBGXLTrWmUFg5G4W9/qfMhWjiUyIeMwemKIL1HlniMQ/c
vczqGUAnPcSs4ClTDxPMcVcMT01PKCo25PAOOJUPAEgFsBAehYyJU9zWR+Pm+UyX
lz7ot7Ydl4PnIsgmhuMem05pamDIio/Zm6zleVPHXV2PAY1Ey0fAHIGSBW/sd+4r
f4cGhzMf/rHmomrxt+M6FELL1bmG0JYiEGS/2SXYhWkAexHkYyY3i4KU15nnzrF9
GbJLDlL9HIxEzxstphfN+fPxqahXjD87ESn4pvTpgD6n243HC23pKZF78Prv5hB+
t/PQDEzpP85eTQlsKc3M8/5eT4DACEnw4wrQ2jZMrq/d3cTLPFnhzk/nrkR11dkV
6TIU81NdW56d1W+c3H9kKlgemSSpXHOs8wtELA4W9X9SkD2CCvXVPWuhQB7dSwIW
5kR/USPdyi5MgzH4HHaOnEtOIlQu2u3xKWd1jBHHC0zFFno1LgEtTEmcN2r/EPtf
Im8dbgND4NPP6yfRfV6FxsPH1mjGjzmV5N7UqpNbZ85Rvvi/0FVepg5166rPS5CF
3PcV8T8OfkHM3+PPHsLNmFmsN+9Sj93d/Ec6ZY0pELvSodL4qSoRlnXYtX+8yMpz
f/ONPqHYyTt3zrsYrRb7OSozpElQObo1BzLr2tpebMWI5wDk1fMl6hfeuPLH+fpz
3QQRf6c6Xyi1RJSxyupm3TsadvIMFteSLSfa10YvfsG8c/YVVs/9sbldKgcFtoRr
VXp5n8q9sq8+3gCESdUgPbpSIDz3b4HUvygYkJxYjBKG6wtMgy8Mt7JLo48/Rw8s
gkZh+VsJfQesFUpssYmPZQ/va8sYwMt0zoqPCjzFFbUZN+nBQDjwcgp7HiHG9H0C
q6pKzN1c0raxIxrX1t5tIpYi70BFHeHFYnsJruCmZ79/6wsVhfX75eDc2NduppKM
lRZ/3TjzbsFVgkNvpLPlvGX90Bl2OuG2IJyH8fPEyXfQbiySzEU21/RkIfK7S262
niK7goshDI1jROBTII/k96xf2keOuceo8z2pWdr2BjcJZh3ZyNUmtxFxiACvMbAj
3pXV8XVzllAiCSi/36nJafX17jDOEOlygHn/ttuin5Dh+uVb7X7sVd/H8eFEHYBR
dJS0sPVZaqQLJ6GhXlH42JnefWQIJD6N6YRSL+LYTh9l7EIenhYC3ihRXknsPV7J
0OeIBUURZZH9EPnGztNCqVQBN6La20+nXe4kxOlWv1acjjgeWBgbOHY9m8GcDqeu
7Me1N9OSJng61zaKNAasU3FYykf8omIr2rQXYqpoDaVfZO2Ogcwcerw2vHE8darf
1hLvvdwJsZpl0rAyyE2HBYrNKs3Y/n/zGlDz3psIhfH6Rdli7vpD1FhL3WF1t2Fw
A5KpkrNQtuDIaQ0pNLLfX2R4s4KBLUnTD8TRu6AxX8UB2ei2JfnLG9kmU1Fv+Jzc
uBw4XzNCk1s29Swgs6ly47tERgReYbnV0VEVRfxu3QdSi2rXMDRaW0w6eF9qNio3
hukXigP8/dMvG5XTkmgDiDVOW9e/F9CsGtmJjKJsfsE3mnfRPje104AZ8jJf3xO4
TiE9+nJJCBdtfCDL9JsKpqTi8nI9yb+lqYyYtDjrDSSitIXezBXaekPngF4XyKX8
OQAXV4mYUj3voksGle3OZOlkPrgT48y3zDkQmotygMWVR7K+w4wuq7+e6aLdlpMt
T4euuRVdsPK+/O8RYtdpqX1LxSnNdRuwW0viA3DVSjS3ta4/hnSAyAvmsnB+AVv+
KE8XWLk3938IjptfvUk39hY+iZUInSisVZa2DovOSqQdgLuWqlQPY437+ykYhGiy
qvePZdveJjIaxGMTf0vGWbWXZQanNzlu2zYOJp0lipArPiirQT6zNb+lLK9xgxif
p0OCla5Z0s5TxI3Zafh4IkZEoW+c/KGsSHSNAixFQQw18faQnGKiwkhn8yO5hiSs
ynQ2ttOI/WZ2c6xpFjY1VMHUrpkno/iR9SdaLUDC1iuUumK+u8ZFARh0aDdpWEnv
8Jl9wLWXHQAMwi9haNldnlYidBYvAL6QGqdOw2q3dwnspd3U4L2fgNnqg9Jo5Uv7
zmAB+vCPIaM0YQX5llvb6UEduPXIZwlxXsE2QyR0rieipEE10UD/w1MmdREXBkfr
FbF+b34rt/hynyiZYFZnOgZFLlv53XcmfEF9Sv2Y7r0e3rtBoJh4/qia3JhltZ24
2HA8WjTjsZNoNpPYn/djiUYHA0T9B7AplLP3uanM0fTXyMZRjycphIypgVTSJSQA
i8BZpEB/fiuOVJxOOiHs2YBAmZAiArwtysHpfxDJLgbYhda87Ot8jHFFvyNgj4Qw
Jqgzabs470M/3zSnLiAVpaC0usTCek59UTWAvqMG9HD4RJHVz1idbWiotlGDObG5
g2ZKfKulaiHROh+QMa60rJ9xry00dXGmJJX9QXoOlIzU4JhBbGT6sqUfeaEeVvIl
RjtRldnBwLaXdqEGfAJHvZ8G+POcSAtxjPjylVPILg2nHWWNccJkFBblFHgLKkQG
HUpoWKEIXiP6n5xTaTA1abC+8Dh9f2H4eqw4Ebo+pb3P+giDrH8Tbs/xqT8jtkPP
rTS/npRCqNolKz70POFgCWpDnGs7m2j8+VYN/+yRDE2MzlDKvq9sc9VlGQ6P6PNB
nasC0dTrN89ARXb21BZvYqozTAsCXbYs+FT0elF0R6kZRW6VC7Q1bR0qTyTpGRlO
49mxu9gM82WaqtEsDuFsTi58oWgn5+cop+54Bvs5MBUCSl53qIj/gRbTL8EKUzVQ
T0iWj0lF1sze3NBDcdYjKbvsyIVl6q7W/mIjr+M4d+tQ52MJk9tQxJkgNMMpXfjW
5Pj2uK093GY+6qp2jB6Jc6gB71OqJV9C0W9czeeZExuh5BPpG4NBM7S3FqAVK/6v
UcHVtEO81lZ+nSDzOIDAyFFcLbDVtsIiDoPX5eMW/M4U8aDncvIlsTXJIFmx4ucm
pKU1gBpfHPfi+gMFYcmG9PEk2/q/3McaQwmd4XrNzXcsfwoKz5nveST/sxw8ziQ7
BRdbPCifrwDdKc4aQESG/VHG2uSx/QWq8k9Z2sGSUol5qcFPryiO/ul3H8RU9HEv
3FTbziP3a4TVF9pk0vmtQYGaLLaWnnRmGIiRZIj9XDVTGL7kx+uQ5UPAc9AxF16O
16Q/Zc/BW5aV+SvMkEBzZ68O47sRJ7sgSW/1gyuqKEUm3GwDVicwjNxbqnyUT3lZ
wmNb1x9CAE5e4tvMOtzHMTU2skh6Ymf5dfuJ0hLFc/hTWdT99UOfpph+sw45NcIv
r+jPQkHulNCid0snxRhjchjV99GIzNwqTTki/nWAe+bjMWmyBx6cHMJPDR96hMXF
JZE9IJ3CShHLHGUzHGPLBI524SDbKw2rlKbhlexIkBIkQartedm4jEZulE+Jrq9i
w3DOSZ1F8TKqzocNeM/fmkb7zeyrMjKjOlmAfvoBxGIll8aWU+7g/WIzACiYaKPn
c6V2gyqt/6kFe3j3+Sq+E6AGTfc87aIm9KXUPcaYtkBsJzYyIZPrHBMqzPhTtA2S
EKM0dZ6T25wMnVbNY6OWScSx2K/hIDx82TxzxmBXk+Oi9DVX8JnVt/MvTZsMIcyi
V2QfWWOgqA1fJI7WEMzo4KHcVUaSXAXFqunPDbIItwVCCqHq/FocFG8ND9oAAGWw
EqeiJrS9ZTua5HNqjL2pgv8Gds+xHOhpcWGP+MC38W3lNweXAzL1slJgZK+W+F9C
i+0RjD6eMgheyUrBbSVKhQd/AwqpLHNP6wUTLjH7GpkOwwSxgBY4j0k9F9YGjw30
WYsz3m0nO17MfWtchio5HIycOr+Nqvg+zKtXOvplVAdb0SEFIDj9e3GHqcD/2VN9
FZssItLEwSTrhlRO8kjENiUB+E1/tFrUtC6V/fALqGUtnW2ujc/0iMG7xwL8ac8/
mS3oX5ZM5oMZC+f8SKkvoM52txbHeYpw1TdL6bwi7Rsbal7ds26is09WifurKZH3
gpcOqPpIk8dyMR8QVBm52Stkv0XLhZ4ngQ9l1l3XmKxych0bLwrj4h1zT7EKsaME
7oE23Xgm5PBlLAq8IPgWTgmsRfkaaGR59bQvnMX6Q9KU+N9ZZmijD2K7KYZI7WTO
CvIJimeEawwp2w0bqL4K/aDEnv2m91kcnV7LmRNyJmXIylQjauN8UJPofPaoxeF6
etzdHb3vVbjpj/+rx99Nx4seooYdYptak/DNq4BQgL6scgaiDzzhQxT2uYmEyhzc
+KvA04OoZm79xcg3MZVQVry40Xhtqv9DXiPN/ROjOIYrnkMfEdfe4u8mmwo3LlcD
qrYenF5TwunG6evpdbUVq4PPG8yEN53Hrni0EdOE0C60AQ/acldDCgGeIIBDlo1k
5Qby8k8xUidkKWDmWTAsOmnUCSbYnNG6sasqN15GGhFn1jAcZCqzeGYKqLfWH0a4
leiJiWxH+1JxHhi6Awqf9UGB1xlzbq/US+XgC63cKcVcZgymvJiPgg8H6WQDUixh
I09if6swfvVWtMeBX7h7ApZ2CLzY3OIBJvSXbmY/7iO1IAqSbZRzXZGrw7LX1GOA
CK5ivViI12Spys1p1s1xvdKQZ56biMk13dtHy1fwKWBiSGiu5qIQjKm9wFEjPM4+
ty78EWmiQXzs4pQjp+0IbcUwnYPhA1Sr6P6VcTilskpNvoYaa0fkBxkfbGl8uWYK
/n4e5KqHiDLWKmjw6B9Z01CwIQOHgNyLnrbaDfZ0CFtubrA7mHhSv+pBq3oEV/uU
q3byrtQQ72gHicz2kl6nzXwWqdLVLvi4o7GXkFq1vj6C/YR/IrZMREFtxqxK4HPW
M4yB8IvWbeaz9yfoCZzN9W4PEB8T/xiWSQq6PvgVq3vyarmJDzUuTbrgCGmD3kip
yG/x36nlOIUNwlGb3bp2nDWAmQfogBA1/R1/FO9EJfaFVgXithp+1FgsdAAvflRD
qAe84iQg2akFXRBhokJWOufiEQEWTPRgHWwYiAZB6yfkaCawIzZF5vci+d6f9LZM
pZg/sWHaTQrFEXmNAUl6YyK4CsYC6aj8Gm4uAyTxIcfBpEbfr0vKTOfvWfzLZR8M
KGskxuQFcFii91Ja+cC4UXUY8OOpmwQsLIEXotEcpmAqDsNLrpzsZNPZswRLnkl5
GXSdiubBurfB0BksBvCJAgbpgKJEtA0Aob42vvyOqacYE4d/joe4i5Aq+ZYxIiTL
BPQK00AqTUMtRXynzXTgZ9nBSUOrS25wkqMNXH8tH3q6MfRWTrbHh80e57ZcXw5v
nSoYiFQl3G5JafrPHoU9at1GEirl83d26dXE4/BtOFnaE8ZcbIelejYt1kzDocsW
L+UyynZtNJ/ySK7ZMVbEkOMsO5cY7Z/9em4R+zCReLjLJ9hGRcQ7wb+hBUQxSMTy
PZxmhGM5/mQ+KVYQG6sEB0S1LAM5sI7hWjHKnvNxPE+EngyElXqW8DL+hoY7QCLK
FRUHVquTIOdK5iLxKaDx/vWetp/V5hj+kOs7t+QBNspOXd6wSKkoDzrmF6EdErc+
G04eLuByYQ+Czv0Do0S5NgXspP35uhUJxal3u5bou8zmoMQA9uWph9SZKcTWycaA
n+CD72YXDeYq85FPwCz8pFBCIx9deYSonEPdJT8zMIEVXCkix+6Ghdf7kHX/ctEz
2NldixpQKkyJ83qHjqogj8oKdsDqtg+G5cjpww8KzpRlKVx+IjJ8y6Do7sssL6Jw
ySGMgTlDk82lmu0iWcXut1vdn18JMh56jO2eHiJ+TYGDsvajymQ47U/U5XaglP8A
JbTGploBCgpJSlpvzXphPeJyTY+Rr+PCW2tB2zqe+MSJONJCLAU5isL1m6M5PP/l
erK5SkELqQuQWMS+lPPUqtWoQFJkzuoESPbZAmzos1n8q029RMRAzR4UfM9X4+dO
bVU97cwBegDgvgwtkULjbczvLnX5mu5CfOrVC89Bekr/hmbVsbVbb2bWxqcuYRwm
Ew5OpwDNxg5jmXve7tBuoJrotBX1Tfuw9WWvpGu8F6WsGL7xz5rpHm8xoYMyqme+
tKK5trr6Vgg+TPqHWBCrQ5TnzyoxOoPzLvF/GR0ZViRA/RTi03pkczNJrvlxpyXd
SrMLbjwu982gDYLyhRP/iKbTvptz1nQpjzl/mwuh71Ldy3O7KT/pkRqU6pD8HzBX
0/K8U7dVXAwLWAEFPzflTzog3+qvahvvu1Jfsnk5vf3b/GBOX6o/O2e0Vt1KbYM3
UCe0yjsdBkngs8E1grqjjC07oe/mz3jdXcZX+7CNM7t4Yz79tcTQnVAsHH7Nt3ot
wHhnXJbb92VaztQnbPGfSCIP1+JFeNw8fjkJEyOJP4IY2K9Q3X1PkZY09OeESZFY
DqlLXL6hJwrysIes3Vpi2doYhK+cJu9Sz9Oj08IReU3LkHeopWf8W2eGxefWBU3x
NNo1VwzZRqCaLm11rUr/mPnUMA6h45TqW2T++/cv7cewh6BVK3HMKvnR2RdlTN5h
nAso2ozF2g1ADb1ZCTYov/NsuH8cSHb2qLX8OPwLU66EUK2MBn2pTCFCk2LJDYSe
j47B62tU/Pt4w15zfHbe435DDp+SERJl2sAKypaY89XwT+LhHbxwbWi4JD8VCyRQ
f7MCyxgmfNMHjJdEvtj/704qn9NJB4RddIKc0DAn6cL/ONPjMJvjVr4t8bIHZ2rq
DzMvQ15ypQcu/REQSvuaqYuddxGHcDwQ5sCgIS5rIErQulYWo3tMOlJEnSfdpTZW
/PX8IJp9zB4Un2ks8PH1FPLpIJEGOzdhHFoaWJ+s5jmeJXoPig4L2kUpECKLDsbE
RXU/VVbJgRBRNBmBXsUhoWXuDWB17alJcIlSHFWbNbn4EzXAsrd+/+6Ihvl4+Mdp
Jk6sQKILSTG0hq1W5Kj3txs5UGVL3wLIDiYw/KlivYW5aDtOj67qiWBQb4ZnaBbZ
l4HEdJR69Nk6N1yX77RVRoSKQ1smzXLm6NiTOQwkBYZuJGQ2/WdG/8AIrZ2Usf+D
02p3eoEyZbVhQovq+02GDj4SZNgNL7fGbzofhFSsI0mJZMIemNILo9C3nns7+W44
m0xNqNMwGc8c+cb/pEWe3qJCvCadqVI3KerTKWmGEBcicoYgKTcYClJ5pTSqgeni
1oXekA/g0OmBgzgtnWoOigzQUqWmDEtRwziQEb3KnjS7BrSfV2uP9kY5KOB9rZvg
bFofQCwzA39BHqHf51mOW0SS/YRiWWVwtKMB7DFfLtffgI+fC//ByhRsYm5VKn2w
uB2Bff6nV624JVlnJdgpaSzrYXzdPkY+68ODZC+xgYLEBy0lvHrQLbslWIxnqpQ6
GmFwYOYm3QPWUqdVajt2/FylXei9yK/dfXCqqvc16NniNOYWCl5eVKp8GEJDzG3o
AI+/CVcYqwOadnXl9GILbiHleOe75ws8OEtYz/2bU/DX2kQILn82Q3+bqUEyAzS/
LpoauEBqeeoBpVnLQsNJUzG5j6UjC+MXjIdZc8JJaia+FryuJiPlZLKGZJbQD4j+
2Nj6fpuRMqzC4YrX0e7n/HyWfm0eE16LP30ME65rgeHCumQftBfWlQUlpuOFDbu3
lzE5L322Mn+2/iBxcoS0TUQHJs6KNxYqo83+Ud16TNRSBl9GghNswsw1K7aSW74u
5ydTxfH5sD6plGmXLV5yTpZievGV+Eg3vBtbNv5BEkygbnPe1KprnYA52qJh2M/J
1czvC9CEpsPB+I6QCnL4FHJPnMpZoOfD5M/otFxjtzORj735vkwt1kfhRzddFwoJ
I+7P9mBowddZbpQNIYSCcjrs7OOht6e2+7ryUHv95ABaWSwh/UT3ZRFvZhgkh2UG
U7NSlTBG2MFLniW5DtGJ4ZtVb7Ep40HKWdcS//eWxqDUBxz1RxFnVxh7gYKHZ1va
LWIRh+4sBSDzglcOxAiTKIH5owlXTNue1le0+aR6r3mUYeRYo4j/sKO+rsVmYOQW
JniGfs8nA4a+emo8uFx5J4lnZndXOGqqCmR+KWo8gPR2lu2Hv77Pofs9Gj2+3xxz
LWSBGEAFcldtH8OjUKysyVcjCs2RDBp8TANifnxvSm6udvWQzfgVcqyY7St4Qy1u
HmTUv8OquKdsorTD+4eYIvuWHFkeD60EtjUNZ41YVBcnh7y/CljSyUuaizmIufVE
csoDyspUeiWbM8qzJPYbauovFWY2G0sb1UOi3GtjgCSNc6LDhGH0j6QHAgejb1XL
vBMDdfK7jcWZuYDOV8ecmv3WxjvyA4AQnGKlDHi+Yi0JkhH/JpokffcqNjJAYG23
h/hcHyjFxTqGwyvK1Ytz5/T47+9pRk0kCtQeivI1Xhu74E59GJFsyC9pJTtZNvqw
b+KzSTVzyIviHZ25ZlIkcG8AsIkgeCNy1aAlOdVzTyrI0WgEo1BdJL/f99FOeIrB
AON+MFIsvzS8IbgtCq3M+o0hWlca36Aflh1nBGqGcrFudOfdnGUJCr8fXGNe0hWU
Qqgw38U1PdHks0QxueY7Moo09KxXR99xf43+VEJ99qtQcNLDEBG3nLpzPAls8hg6
eR5UJYGfMB9iC3e4UHFgR3w8TxrQ9T9b3Rh8qGzysqYG2YCspr+JagNi65Poo7oY
YrpzxE/RiRXNYMrYOUznC2AI3YnXnNQmMKDYFvsS8AEQ0MVVzoBXmnOqJs8VH7Bs
UY8hk7L5ClW0Z9lSuAIexgwJV47BrBcC50VmmianALUokvd5GWER9ZYDdT+8FspN
2qkWToUly1j79mmWPFWOqJ2MeYGOEuXmp6jzUdAEnB8Yg247TztYPRvbRFS6HUn6
HJOIB6VTyzrjgtH15G5XYlzsqUo/qBMTjvO/QDUHDVaEQWnRhqrBU8Tio/Tiqi0x
bV2VxNfqdOzfiSmkkHN49lw7lhwo8/P7wI/F1xyt3NQZ01smBZqwsa639cAwL4Fb
AoJJH+6NTgX9HgRn/gz/QQuM7aK19IE1p2vNxGB422CGEXEuwGBymv1gvAf72LAH
mk6UaEy26Y2aei+JVX1gV/tAz/+inkcyG7yQuwPnZAu1ieEJ3DWliS1zLPgd0OVN
pRZxAPvW80oHkCswWnB63K/Bs2cSGc/bqklNxkqSuQCc2YRl5dXT3l9qwlwRehJt
eqxXSwqLOvireNawy63jd/l1RkvN6l7P5E+HM+p1Xau8MbXziQpJUcMHYm5lN5i4
b1tBgBMYaoeHfIB7GPEuHwaU1iz68c3UhXcu+DbLlpWA9CT+tRE8mlCHSGdIoYus
RQ4FMGOL0LVw/QIkRJ6svdIujBV7Se03vdK2iuB2spwAVH3tgSAaY0ESMUrVaxaa
uhb6Jr1iBKnpbNi/jDag2wMI0Q1/5kjfBs2F/1ZvFjemdimtsFnOvmo4bcmgM6oD
u6gQB+Li8CAXXzekmOLRtUGHSuaDhAo7GqZ0j9KJguIhoFKwxh3iOLjDOhuw51Fr
dTkFG3TXslI6h025zE4AQY8y6f4mWvyJOOzUEInYNEY7Z0gGdRdXBSILITrIltoU
HBtfAg3psTx0Jjwn/xSzE2YO25Y9iEuG3uE3fbr9zQsaiiWK2QH0Y/bctTyVNfKr
L1pLJbAASkMiCoOVp4gEvlenhdt+xIOTE3ieNhTOy3JYcfoOgAQ7EtRIUUMR1Xea
WWYA5AchTBDuHUbewcz2ILVkRIMtQ8SMQDrFwA+Lt0o3jqp4e2vxD50V9hitj/Le
dijnZ67jBIKAZcQr7NVIqvpij/K1HKG9eTWmtUwPtuEtiwvSlEvdpZgTOyQepJ0K
N01/EST+1bGvujuEIGFHt6eAzP7qpL2MgTOXzuQF8csHuYBpyU/tGPhgX1ykvlmM
H7U1pUVcqE417tI1vhYJsAlxF2LjuigqGT02jWFf1tCahjFX8AOd3PSWj3437Fuc
ZRgo3dpHcNBB68GOqygkrU1nHkjOPp/8QIqD1A2Be/E68+GU2aBAcagAOg+8Sd5Z
lx2hE4jU8LdVtzt7pf3AOZ3WwVqV+51WdDGymtTJjAh0jugkzjn5mA6q6G0Qht/T
RfpPhaLrx0jZl/CfrZyPhpbnSG+k51rSyoqPv6EtluEcPM5l8Xg0W/iRBWpnSTL6
DkHUoMd8m1qTEBB/Ky6bbWSmSsb4JX2AJWb+LraL20G5FwLfC8KQr9o+PA85TBxP
y8MxVIIQy/GuxH12C7YMX5c/AEN4WAhpSVTNoenXXpj1QFWw2mbbYkLfpDhCgeYc
FgwtUr/7fKXaVloJHX9tEOpPRcMyO/bkgkWGiTupowH5uJ8jdUgFFQw+lzb2F3UE
90C4txJxLVXIvN/j4iWWOemWaBZf47pbibAThAoYggBzA0Uioh4D/7YtnxGTLhpx
q/rvPYKVItGDu/5kpWvD5RIdUjaUUNg+dbbL9nssK4SxLyWuliYYk6b0V5lYZZ1x
K/wIoZ3nqPUtY/g5DAlN60EK8aHUbpasGzqKCWXtT+QLsppBFm2ZAIFEgDM7u3+k
qaIDDONhKokTPDKYvId49hvYAS7lYYnUie3quG4DSdiJJY04yFiOPpULWbWUPGUD
LL7JBlK7/me4GwzMe9CFfabvXnPXlYVN+PJ+piCXW2NvvnNet3FPtL4Zchk9ZqAT
n/wvV3OrdUHAsnAxiWH2mgsCWRJC6wT88wTSo3JsllV7OnxCD0bocav3RlOLg1eY
n/J/OjVWfQcXxH//ORDM+NK305l+jQ6vDICqmtUPM6mPOh8vLxQh1y/z56im/XVC
DcO89xkfPJM2M45sb5qcXe+eFP7ybaXC1dAFY0FPzkkM653vN2dpV00vTlhvYzNo
CLr11WSjZ6gY8CRo7JhdGhzDq5PS6LfWxua3nz0Iuo0LbFJL86bml4NbfuULtSQd
pALKvbrUSKalgNIO5LyCEws+Sf0SqZpb+bJucM1p6/Guc5rzxwwsKjPWO/6Geyi+
MxMG0dlM0FEgBK9Jd17EINroiGvxPPYzHVEto2CIJvi3FvshUxIz0q5M7Gv/E1yJ
V+FMo56F9IOZZpJdrWdyEgTQfz6ZEaZNzCWrPhkyxC0Bqs51s1h/mnOse2qNuM7p
4x1HQXcycd8uu8rVoBxn+JnPHAHg5sfAd8GedRGCQEm9GMD2W7x6usqEyZrmPXj6
DOS63C0VFiyldzItyLE6M+7f0aPtjX588Y4ziaaxqIh1X2DZEsQHVjPutc2bZtpT
ez46BAJD3f1O+6kiKGLTQN2Gylhx/DK4850nCjsdUL9g6OE+AFEhqFQUfEHBzfEr
eJFG82Ivxdv/NSSFUfmVos5mSaU55PWQTKJ/EYgTOvV/UbRg0TjyWdLLHf9X457U
vmQr9DjDwXuw5Z7vOg9c6iJL+hYhn9DUPg641+l/oDjZGxmZ5UE79Gogs0CNaEAY
P+8/8FoE75q/Bw30KwgZzvyYnqDM+FkVhY7LE1Sb3uh/qrzTaZoZpPy/9IWPP4E9
Io79RHWwGwkEz2NBSuK8xnQ3F6qWwYGly14PrT7SI9wO7GGLnwVUITjKErq14y9w
8BY0G9iX7ua2ep8N0QWR5D6UPw1+TlD64EoQVK/aL7LN0ocZd7B0dfsZNbJ+BAnm
ClAuT6PU8iaJ2gSq8SkI0j1jVm3qn79PXvI+ZBWAaMjef+R4UA084psoo+WQibMq
Sgt9Tpb/bDW5JKZtWD+102N/ekUFujfdzCwl8IddSTC8pvpPiTSO+28j9QthoXjM
2i0tXjrg2h8yLjpoESjOa6kB7SDMHjeW+KTMKOFpi0g6IHFKGN+mFmkCmWadYrnV
bAyuhEUvb8mluRS+lZTOvx9qsjSU3cBDzQ64WgxKNvvs7OtnT87eYPpYNak/l8Be
SLjcWPZuCm8mNvqhQiC9+ZBJTHNPSbahRsXpqoK0Tc0Y61oR8/bhesb5UfUcGGWs
+Tz15Jr2iQcRBsHLU9e7XGbrLsNDDFciwIjsB+uQt9zBCyQr3B83gKU81nvx1JE0
/F0Qaajh2p76IEObR9Py/ONkmID4OP8SifDK2InNLHEp9B0Y5bZRj0VUKORbroqN
DdjOqUi+vW10ludweLmfCuTaEFGkfjaQfTIdSoj+duaB+YwjAFg5tuWj9/Tkskp4
gVubFtU5k+0bSyPo6dRHTAZLhsb9VYRdXy6vPCQlgNQFcRty1WdNjvLVDgpCpd/0
lIQKM5KA+E/FkH9/5XX5iCYi37hrKz+TzfL/80ShnoVg6MjzXPqOxZDwy/LZtA2i
z7hOBWHbJcb2yWJUmwfqGy251wU8+DUumcSLVWC/kQ8PgcHmSXweuiWzEmHV3bed
A2k47DsXTBOjRkYOrCKnLq03KfZG2itnB/0KOqCyL62TWwQ4v9/EyGczGEKef19I
/3Cctdj6LGM3o1JesjriOcnQMdTs0ZFgCC98Fsr1ttvPeum8IGM/EAb9HbtZivNm
0sR1hHkcx0AIywwIjRb+rzHX18dczaijdUHFEbyAxvtjUe/ZBdRXx27ThdEpjdhM
/qIchjXTWOWWonREUQq6QcdimCuqfW1THyuuJRoRi91IfFIB5XqURSlnlvxDn7Sj
faVvvzC+TCtxPRp/EU9wls0PIUG9aEE62NjVxhAR0h0htesblVBvwaLRvKkeN10p
774z/XD4mwN+vCuWFDnueUuMvpd+yGqCk2jlWxonuTQXkfdk7sqpGPEKxpxpAJm6
6KHgl6di2B16Mtiu/WI3n9GfKG70xBSIAvjqcQ8EWgPWv/Qc+qb2dInjM4m0+GTz
XUwBmM/mGU3NfimqvqlOyzbcPzwUFZtgdqvA0Z7WpojmvHy+zhbryB75MCA2O60z
LFLQ3+Xt8n16YXHmYxucuIu6lLAHI+wEJE4BhQVyLxoXVf/jeEDPca8MJrh0y5ha
2G5uNU53atHAEzyC08LOqpUdaIi2iwKpa7rQhx9vRFDJb4M3+SNBO7QkDk+aOC9J
GxYcDfhl+rimDtt2I6EQvTSC4v8bDPN+gjnO+uPl10g12Jo6pThMSmiU+z7nwNet
31yDGtY+Ly5q/6eMPgE2kPdaHpjx0ykx1zs/Ga/3GzDnlQ92/PPyXHREJ2ouyG1J
iuRr5H6mLvDFyU8z5P17DnDQW2oWyNBgzo+P5I5iQbFzPA/nx0jW6rbiYLccb/C8
SkC1Rd9Inls8Qmzb7qVI6lrpQZeOpQe865YpuD5bDAkgdKtyZNWlzTl44iU8Ead4
m2KT3sPHdvn7jv1ZsxTqgEGr8GLWcRj4r5NcPB+xhW7bDQhB8zSsCDnPTcUPLhHU
t/SR5QzlUSDENYaeNg3c7K+HP7i3wlDjZQxhTPoEW47+fzrrKlS+5Uk1NMeRxKD1
/fiXa3K8bLS9K0qHr4nHKSfuOVcRZYaK4Kws2doHK51IClyRaoeYrEZCXuKaT/KN
abYhacpXz4QSqq7b+aT776qIxgQEk7iBMw7HaLN/0evhTK5O4Fo9S4AtYATdzoPx
WOekGGSyeLjgjnNZqG1OrqknYq0+KY/cK9jEzFy2EuFYN3IbLnO7340D1xBrsY/P
svu+JHuzbEdA23W/nu7Vz1rcKgBoZtTNLYKM1gUiUA+IWlmhMjutbEY9Lex03y3S
UVAMNhjPeagR0Xe5u1SW/WLo5HhiTGidPUBDGyilPcRMHAR9rsAi04ULmBh49D96
P092ElP8/gE2ulhFfxTLmhT3Eb9QP6RqCVcZ9lKlXOfaXMTJqSi7OKi7MaR99YW9
yYcD+yn3fvk7hQGDXYRYQ9ttb8BsIygbZWDnsQaiYZ5N9M5ajtaaBQKK+KAZauqm
uVti29CyNgwSew+OOMxn9+WPwS+vEIOtFVlYcF7tcG7PPaNuJeJnQSoWRR9qHSgb
5ddkKCJ1oV9lBTSHiPaRcPjTjHhwVqMs7eLHQAJQny2PE7zWzkiuJny7GRC21PuG
wfAFSSFy8jCbpto5oBi7AWS3mpf9Az4YUrroY0ylHBJAdSicDlq/j8jp4e3OmS6B
/uMtAc5VDI5AvOLfEVHvxoEpgQYvhG4PyJq2UXcNxtAdqKD2fMBjjObVztS/8WXk
6P6B+W+cqXoLm8LZCMIq620u+Dr7cgapQIVQZ6O9bH8zsfEVCmbWzjmyj2htYZU7
uJ66/HGNGr2Rs3am/FQQTH63JBUF0TW4Rbf0UyP9W8VemNcAUHvUfgTmLJVt8hxd
9j+qNoT64RGjHu+sY4V1k8/o2WGU+utPCVDcH3ACfsVwX1VfxX5VsFk9VLtwfdIF
ozY6A4Qi/sN6JuhZ5ZhAUz0BauOkLB0cRJQu9bC124cK37w/BTnxPLIs9c2s87OL
ovvpecFI6m7yKzUiUoa/FgcDmOWXhoeb0BO+qvQhmPYY0tnpzB92wLNds/xtyGyY
/eAC2emPz7xEihuqBWg1/EPTSpW8mwdt9xaa8Aqanm2B4laG8us2aEYxCLJF3Z/R
fLsc9ZzYD6+WEtytJoVE48eq1S5p0yfy/WjDRIjNtSUujpO+SYpOShC7bKtSPFQc
neTf0qnHxOvI4zm2a+dBiDcTTjaiX6zlmiZy+CcoBlcH1nQaCK6K66jfkKQrAzVl
hucPL6PNJ36F/e1m9nJL7NJ8zL3TsaT/3mDdblwVZ4yHzKaN9MaLLPiaS7l9Npjx
sPDjivzmpxnvk/ogYNgpjhqcKrF00wHaLlqnjXq5OKJ1nbQGmiSy306LGVaJYkI/
NZ/etvTfY0wFVRCBT5HFBZp/fAHANIhQSbyVuSrQbRSd6hncJXcXL58e41fmk6aS
m8Gp0a19Gx6wN3qAxbeDclKGSFbEntwAd2BiHerW/A6T+MQab9YeiLs9znEDsGwQ
khi+mRzuMlzmNoAgElCiiLmf72HOa/9uMliHdsuhbdRL0NfABgAr50xRcIVr37vA
cu8TWmR3UM+BN5C2993ALkKFj7GnN7i0VhUtSutrXelFVMoleF9iB8fmvDW8YSho
QVxj6vMRTencI2gCKGCmng3CnNDFn3U3AHlTps0gsX5XnMEDubUUOJ4o59iz/Ml3
7ccMFCM6qThHZSbQb9kmrQKgTYu111WprH0UxFVYL+Sl72HHnktUndBLPThEoW7y
N1huS51qbMqif4qonEk5VXyxw7vMOFHr1lcGPNxTcJ7BlHY2DO7uAvsP9RetvL1d
1wVkw61jSDa2kpH2jd6ypeHRellJJBa5NQpK9Ve4e5ldOGSs8y3MmSBtuoLLfUj6
HA1lXVc10LrWKvv/eNv+4Hb3VEUyjumYCQZ+XLvPxYdW6tBQwCr8v2nzGgNupqX1
oDRG0aFGGvfVcQP2WP+iznHYCh3eR6NXHFbdFoGAV/XvwHmyOVT56WP0l4/EaYQA
0BZt/z8tfU+VVCAlyv8i+CKOPrqycrpJzBE/NLQ7Fj9Kqt9uYqKKr/if/Y+/+XCD
R5HTzwYwAPwDLWa3jAqGXO4snf9madHVxw3FzH+14NzOWBOC92pgXMnkaBWjWyqh
/eGENTFQeITIwpb6A6PCRW95AEDn4oD6NmGi+PhLK8xRzV9zN32oKVuq5YJPQaMk
tAaO8yh5s3bCqqf1/eghFPejZ48kJiSiQaENx9GBZ6ADytZkpGPaN8Dd4rFX+C0N
BrFJAYbckzZFb9Vye8AKIi5AWVk9IaXeUdgCMpf5XzBnaSrd2EY8vMZXfrVL3giR
VdIgMEEo/f7SM4O+cc7fUQzwbIB4h66ybYdfuPjZ181BRuSIXpm55ugrg9Ko2+i8
ULqC+q/g5mN/3htWVs02RzuQTU0XWeGHiTDz+A1eqjkX0RIbDnm7narxivj8sndM
WuXNjwphzIOMaDFYj0McSGN93zVDNmOwurbm1OEV+3l54E0to0mD38qFKna2sEXY
RZGL7t2vYWQixGxUsUSItCOPhhmz4ynxKTGFYfkeMO8SfuXvZsHKnsnM2tAk9Rge
Zzw7fkDN1ArU7nkZB9TkP0Mxs6XF6/4dbDpdMKsR4L3xpH3rV9ta6feDBrZmNvVX
bbDGfuHSSH0F4SgpZ3A6qoNf1FOhhypXEzge1sARwRXGphTcGDYzctP0kULTNt3A
zOslr8RvkjOUFa8G9q3CH2VsRUlljorDKSP+NYhJWgxoC2bduq8bv4EOx1q72L6U
7mkU0+g/jd7B7g1eAUQT0X+KVCeYnezL+w46wWrYkJo8rL0FrjLbqzupOeFTg4jQ
/GJ/367XZhn3pNrUxX9g6Yej/VsZ/L78AGt78qO/O4MTYUpC9U3vocrreFRm+a+7
21yYaIn2+rSiA7C1vWfZKSoEOFs9x21qv7ar482BPMInd024UQMvjHz/Q0/lk/2q
BZrf/uPyEZ4YgIgq85W+HPvJyPM4xW0eQKND1zBtz0dOmjZ8D+97MUjz1FcBzoam
LuqtGXKsh20HUpcWMIYTH8MaYC/bREGU+dy5tfJG3kQWjtAhGJgf/qoAjzpkP20d
nx1Me5rwkdIYs9OPunYqQzS8xqWUvzL4mCNj2Kjx2IOVRFvtFEBdAfQbRctueEkE
u9pbr13At/HjCLRGH0dm6Kxdrx7dB1PXsP4sckwDvy/XU6yLaabVudi6C7FFYoDe
we7+f5v7GBGcmaAmgByrS4+J5VuWjEw8ydB+QCJGkTpuRsW5ILANf2wluCtL8z3C
5X3Q3/c5xvyWG+phvqMuES8O008oaAKsf0pSw4gulojxlgsm7jvHqd3hiTXdagf6
cn0YbM5JSBcny1UUj6JarUnZkYLUMOi9srdvUpPamuwlN8A9RqZvBoW6nKs+n3ts
JUIDD7R+2wnvZXsu1QdcvwQUEKlLNYoufO1P4EnC1JRS9kItODBpRExH/h73jH1e
SmEVs7Fm3Rq9bfGmN4iNxqbWckizpSt7Xeh8yn31b2/l3n/qODESjYfp+CS4zqRS
k9PoRoIC3l6AMOO/0HvgRiviWpBk6eAq7whk6hhY2JjLYKKrnbnx5e61kFJbzj3w
F1Cz7Cfo0nKFt8HxYCLKwitDSHQ4mV9q8duBPrJaA7rMvkSHlSCv5SpWl+fFkhXp
6Pid6G2gPWPe47sxz5gy+Bf/rbGs+VxIWpABbr1x6ccQpQ5KGqUm4vtsfQ1H8XtJ
B+tc6ov29TUnnt78yKexoTO8sq8hz4aS+eXaAd4hHmldolQoiazxzlE+Zc/oMtpq
CepLhVn1g09oe7HgTQqXOvoE1xUW+FBguxvkkjcFisggPoAKRR00/GSc9DEpquOk
fJ1bkBf64YW6zF/sP3x7r1JWBWECu84Oc2m4Km4AYU+7+r+TIgcuPB+A3yqQnZPI
vhqeLyUt55ehzIe9gywBDUGIxAYQEK78dy/1kZg+6Gq3qArG19TlW6ci6bqBo2d4
4g7mSK7Rk7Ac7BJvEOVvPgFijuTJWz6TcgQWc/mrHbK4u/sXYI2eeu1VOydjdEau
OorkA5SGPMDUyqmiqGPkDYo1xHJBFDkTq6zfv6nqjGajYj3oOlW1Fi/DbprTp46I
az3h/FOnJILtSe9TbGs1AyQuDlTV7JVJej1wiEPDfDK0kc9BpNWLAyZpv958qkMO
wrNw7EvHVaK3EvzUTjck0+6xVahafUngd0EI0YDl8VIT0RmVcuffzNNCSe3ZlwUs
bBZi+GGgUDHGK0C13Qhz2utALTn6L9exfxmp5ayNz3goLZa34V3ZWtDrrt30fyLn
An1XUSFsZ1Mj0+1zvxzCnIVyolBm5M4H2J0dU6L9J0sCGI6mht56AuYLDgs64b0f
u1bb6qKuSHzcRggpjs8R535q6eMuwV4mIkSuyFUWSfoloLYyfsWhXdODyZhe1Gf9
V14RTL2IyIicgISTmlGdBJ2iofICfCfG9grZQbu0frFcwqcaXyjGqNUb7g+Nxl0V
gFmuX/9SeNC85uz21ZqbFOenNEVlMkAmg1YlbN/BrzO8U10NYCWp40vBp7r44Lbb
aDuKOo9JpJaDwTNNU/CH4X3Xo/NpqD2l3wKUl/J+DGrEHaxyu4r/X5f6gxrDfh6l
ZJ/WWota/j8R70B2o+1jCkg0eJ05kqATiDpyQi2J3Mn+oqeWI/I8M1QmHQfkeCBB
6GsXMpuiW99MyybpDFEodkgBrFJWuX2Rsp+POsnrqLywN6+CZDHojDs92/lYH7NZ
0R6BwrpakMyiWip5gH7mEWN+wjlCuJuciRIIxnBZG9OiMeazZ9pvOfM7vLtPXRBi
BTc7FvY48YpRZEf5qMQ91Ap7t4Vp1Telg8LyrvkRT83C1CJ2AWUa/kZUJFdJqeMT
FU8iFawRDPApZhh1Q/BWLjuWVufcm2KNkrW0He4P8SGpkrbzfX1YIaRkwx/8K08x
A5h6OI4odbxA7BzQrsTAsrCDr32u2QF7FSYXEKLLyOpqQ2frYwRuv4SVcHb2LDVL
EXC4IWxOV3/Kz/FGY33fHvzHZcLxe/Lt+y/gnJ9SjYnabXhCIpQ8EHcOMmL9Znu9
QcZWZ0kWK8a+2i7/wUKfnI+VUrssHijhAhO1WZaPNDy9JEtBQNRlyLQvHKZO/sYR
48J/52TljxDt7YcMAjEzqmR3gcKXAQaQu0Pn49oH6SlVZpEYuNajLnsNfK8e3pBM
EUpCgMDoreChRdkJJ0QxbvyW52darMq0dq5nilQ4VlA4OXzhgQJ1Owm43piYeKph
hkQC+ep6mKtwXYjKpha4uI5rUDOurqHy1vCo4/KRawwMzHCkoabeqPXMtZE9HblH
OXaG4U0NNgeWK7udUxsnKkdsKw4JjaoXIedGMDXZKN0P8T7yIV25Fh3Zj4kkv0OB
A0cztxmjuOgcW8NERmbzVcXuRTVCEVaU+FTgBcDwlP/M+QYzbrEuWtYUVzSkyHvD
UyZpad1AViHnsp8vTu/bozyYMnyazQcU4ubHFQnQNrxIxRksNLOZzfa/gcjghprD
tEyf5/0wIJG9p83jvOyD0NbAJJHLun3FBOPKSSk/6vxb7/3mrKaIzk9LtWUqvNNp
iOhQNyr5fXzH64Tnee0Z7nc+RC5ucqUC9ikMsrg0d/+3UvQX35qNtjk3UmXzCWeP
tDCo47E8/J/3Uk1JBJ8Dq6WBoijGo1luPZRQeS6j7An2OaIlxAQsmBL2jdHvLD2i
L/1LjqCLO7qBhlZs980q6QFDic+xxAGpgcnU/sq0RbI+ywo2aox5b0xk5xSSfhBi
bPelYSYLnHRxwqGlIVxIF2U3rRR89Hqs4SvWkSMwOZr4s9gXlEHPlWBo9E0j5VEB
s9iQ/qAjkL4RUJIyxh8xMmwM0cE7W82wTnZIpIlWUK0bpmYU1AJ+5LpHn9VFscZK
uR+YuMq3zuThtaQosE5LZ+Emcp/N9hvS1vV60LTUdl8+T4ZuESbPV6rLK/CnI5tP
KkbcENQP0mDz4t6iAhCsbPjXdEUSACTPmT9l0hCRzSjaaAwxIQ0YsL0XF+/+upL6
3h3sdwSMk5pomWgOnzkXuBpeajUYV4jZJONQ6eNv6fMEAa3mygHIF2p7K8kZrDWY
eKMwd/FgA7x9q6VZyM7gEJg7sbRkoe/u0alb/BpJqIq+wgz00xRHmCU3d/D66WhS
c2o0OP4mLmXJZcaP38IOYLAUYkHGijxQZFhy0C3pO7Q0MJW8ALhv1wuYRwz7ys0L
d1ZPUaihMnscWmizCOFEp7hkO1hmRRYBG2lGipFgtIc8AYRHu0/tHcda67SY/oWV
b4PUNUbyRTzoh8GMAjVYQDcWfAobIK9wLhDffFCsJSmACD/gcOHTgFrHw6jCkjru
MJIIYTgScsszJYlyIN3hM3WXM/P40rWdrLnKiZC6pUzrZHU7enr2Ku5/4iO4WBjy
h8dq1c0/vypt7SxyNh0Etp9Q3AnkgStyCDzbkci7CPKmnWf8h4tJVzM0tW1efBJV
LsGw6EfrL5VAcFs+uglIFeCb41BRh+ih68G2Tg668us6Om4bXupqjQiLrf5nJq2a
XL5XwHQJmd4450Pn/CFfB8Pv6MZ2tTvNvOacfF/oK8n7qliUmvdin2CJl8PN2BTM
GknmNOvQR5Wj9ZqPa2xET4PTHyIbkK6TC6de47Orv1DV5x3RcvHY/Vpo41y18sF/
kupP4Qe9H6RvB7fz6J3OybGbp+D0vCzJZfRAqujzgPZxbF9oDLDckSizmMbfgcQ4
IaE9pvD+bXYWlZ8UTCVhLeOPD5Y/GUo9oAbKDj/wBUnmdBRyE3lnVZi5b7K51iKw
v3/Ex/RNemNDbOqHiq97Z/TPhKpJ81tere0tTTRKRtcydNnpfAu42yy9BuGPqgWX
X+3mJzWpm2AXfy22ttVsWpMAtM2jKxlHScJtxDakjCjRlPGZrncOw6VuH/YXa8db
cf2utWTiREnf0dhUSJnBNKZ4uuegS+RNK4CzJ2rB8iy7++9ZQvFiogj09yBUXekJ
DgbiSmmW9La8xEoxzZPq0pnBkTITa1IvPU7UGtrYGPN6fl5sV/ChJT2xFzU7Hk1j
kwJdqXc4qhxteIdGVE1GIsQn1D6xSxc8sUVSBCg03EB0/Y6ugYJuMFVQ6Mf5CeZK
KII1KS002pTg1nIEB8fDrk55U0eb/2bWlnpdrSuYXC9fX6JLcjiYqghcznR5Fqcx
r6OkeO3aihA88yGJI0RdbsPfOcaqJsKCmmW4URZDehC8Mkgjj2fntQTrkQ9iJBRL
T2uXrsBwIQKZIqaYf4rPs7IqmaVV4rAFV/A9p0g6b2VMfXjfFqfjxlcKATieubry
Zayi1wgr1VCcMPX4OL14AiADb9ahedOUmVsjjnuuLzK0g1dnP+uHYlB17SAOdQ6h
DbAKHUKFjAIV0/wzjY0nJB+h/E/oAiEKjBYPgsgN3R7BKwDt1eEPHShLjwnCusN0
QuwBS3N/lnoZRKeYt41L8nXfle11mFostx93QkKClGbAANdqwI4KizO/FeiondHs
kcAQPg75rLc8FVv3EfKY+krCNoJef6Sf/0AqNhelijQ5VlMTsMKSCXtIyqJhIapW
FL5nwBZFooUyMjmPI9nMhtO6GwQF4487n6QT370nrMOA1eJdVAFnhNBUkHWirCMw
YtOVVwXz8/JOpMP9uC9sIRjuOQdjpniJaTwDdOhzSS5DMja4kuWIxqhKnNgtZx9u
j/2lMk6s0E9NZRS6EAfmHDe0Qwp1j94iNReIYhUr8A5aOCE1GdK0UKj1Ib/8IJ4e
yN2ezZhaeJ4uzlizUye5St1Yh1RNV1NUWonnT9WAjYgakZHm8rQ0/f2AcmvhjW63
/eqeYJe1z2sDFFt2ai/lgnZH3/LYjr/MKbIjE6hUPaaIqXvsl1BJNu2/5ZeZEIBH
RSUeesvnoLQHB/JVP0NT4IAGvkYk0YaavOwUKn1utktJz+XxhvSazfSenl21gad0
3B6+QlDhFmChuQVQ08BCekPixdK6Smo2ZxhUOJwL0h4yQa3h9U5oc/FxHIQtDuXd
zwHG+N9+3AywqnapaD1R23Peqq/IQmOMtf+ITOQjj1125lwK436nw82gTcDH5now
+5DJPwY+N92ue2RoemK9D2FFm0zmoyYZ71kJWvGzoJu3WjsSgIwLpkvlDeq2hx4v
mCCInZcDUVlihCjlbleBf/eVT7CoV8cyMlCi1UI1l/1jQhFHKFDNURTWfdsKkX9g
mxg7yC8L1ruGSrTnTGSM+OP+hKUsWZE1AKPPPvUZkCNRhtmWY0BUfBG3tL1T2KDP
IUwmSH2Y/R87LOG65P+ZaxtqmuLZBhSO1s8aHSY9vK3qyKwtcNpakD2/6PtcC8Ay
fLzs9JCpEsR3ppJg5Y37nXAh527Q9tOrNekSGzDQ4Jyh4YC6qLQCJG4tQM8+HOUA
aEPCj/wCGtxFSkNc+/2dWDkTA5/1KG/zDsavPSyu+47wYe24JB9oo2ls4OS5Qg16
e/zaZmZ6hp8oHYhqyHLgv7PSqzaMRNDqZ1+xyZ3iAEv5oUy7GdhLFnqIH2cNxbPs
IT9IhoHGVbb8WX9JlOKA57X0G/AJRkL/C9IZh6IZqbWfeR+xuuhdoczCV+oMY6FF
BoqU70h8wN+w826VV9FLMT0bhVFD8fSdLdhXn3y+Dngmj/9FzErs27fFye0emIax
jjSle8WxGhkyVw3EUaOuzOyK8SgO3VMesqZppjYVKuUaGEUbrzkgIC8s6SpXSCxu
5ILmgpaWeAIoi1Ytd00IK606/TYs6q7i84CPLacPRHWOa39R2APgtnHuq4tLy2fF
qWTbhW9gfcqPi9Y7LpiBP3rgFFfZsyaort9FPUerm06Et5mNsif0NpYDwnRWJ3dl
sZ2ayyqlDjWzmxI1I/tieNROwiDiKcluSZXnxFniHupWj/AU7B/C18331VPAJL10
v29HkNjzJY5gnllspbOCnr2i06Z+B7yqf+u7qx/MiokgJHclcgt/C2/OUbXpLCUH
9Kumle9M97NCswIKOMJbZ0SO+mkbCE1MUpWxG3G53sc7EpXJNKMUhgsMk4vcR2l/
oDDMaWfwqLDevNOc0IIy53r1HYEhNYeGsXttYeZjHSvYrSjh3Yx+pkN/geeCGE7r
6cH89yQGrOKUct8ga0lU0r+XJspGWNz3J8/2myf+SiCGYhV2aih5dW4D3spAKH2j
tM69ocJTN/WHRQUyd4APuD4ORS5ACQu2lZkR8jAZP1IqB6ZomyZByk7Uni9Yh7PE
HmH7dzbChLyx9wPkt6DI37tcoFI37jafkXCGmJOqvnTylT17rBSQo4ZayGomG8oH
EOR5gYp4XSc2WmU1vVoOrERmdu36GQWMgUkdiWjq5p+FJBbrRobeK6dVzxru1+Rf
seZDRKaq0heRempPWlGALHigIqYg9fCS44CruLjdX009J0rJRki6/FaGyZtYjRF4
7SDs+GOWwC9iYEL5Z5gGiEXyCfzpz7sa/ijbDZtcEBnO20yTGEQB62g/kYn8RhDV
WqzYM+jge8/Zz442tW6QigTrEjHccDujvo3TKxv7IcrWv7e7Ao8h5GibADHe7OoZ
9aw6Jmb21DJl03xnkol2RrlH2DwG8uySNgmS79SgQw8jjmOQ+NwdD0oHhnTK5MIx
aD91e2NBiWpJKu3axb/McZBi8+xuY7cZIUI2cBgvelPUtjUlb+eN4pbqkOyiGvUG
2siRG7uu/UgbXuwpOP9j8Domtfe68E58e29XJT+AbIw0x/wgdgynMEh9EA0z2V95
cU8RIo1yhZVIFCKG0iSkzJqcw93xVBL0TwPDYzz0M7tKQiQrINnM9Ba8i3XDb+LR
hd+1edVRimzHHBD5UWTbjbRcDlgDu9Wfrp8rCiMLID/6ZAL+me4MNFwjaPeU+lrG
PQRJnLezxlPXM+xkV6o1MgI04VfaLw6uATOMbGtjadxZVVd10c6266MU/yYtG8Zs
eQXOUBf6qjUOGkdfvOqi1f94A7b/BASZsUoW4jIAJQkhk6akLkwwS1anV8FmUj/X
VYOqDQ0qjhxrCIiKoqSD/yFeuR/VTxUYz7ZFCCHUIFUKQYJsJAq4oxS3hdpBRpzi
jRKxI1iKT4cOAyIwR0oq/rOYXlUmq/WOwzActPuyIdbYyGT9lVRqot5a8YqVUJCe
teY0HIOoc8wpaiVwctKpUOuPzhXSVdwEtVZ3ryM1a3rnlQAt/3MOjlWJhZa0joZ6
mOSQ7/UJbZzi4TUpBXYbPqf2EUohJz49Zir7grJY7hUVWTD0mgxj9MsdizOGr4U3
U/BZwW/oQP+4tAPWsqLa11MolCEHqYi1YQPwg5+rAamBcmpXbsbjyGorNqNPu5Ub
lyzQXGSvIZsFwUpZqki/v7bqY1S08As2HAXCCjoeaTdtrNrFj2JdITGYaDGJUs72
HbO2hoUjvbaUPfb0+eaE5I+SBef4hVgQdj7H3INSrCYkw+RbClrwcfORGASVKS90
Zd4JzXzbCAjIjIHd3XcJmEyO4l0V36ptCcj1aTtv59lV0HmcdbRB/LJEqySST4IH
mvLYLgVohRszlK8lnUoL6o+2ba1Uw0OrvS1o71k8nnkOi1dh7XRzRxFBHFUNFTde
JQd20u/xabHRNXkybvP9QFLPZ08/KqeUOgr+B2FzimWELiWiuBcCcI3vX7sJIU83
hV5p+ungtoJQ4Vt3UOFcZZ7va2m9CU9z6bY9Naxye2jALl+WHTBx2G9sI7K8JtjX
apzKw1NHfRkku3h0BMVZuWHIw3AjTP1201yLV7xMXqK/mAohJ7qhHAP72autpoOg
uq1xW7uS1+3kU3uWwBE6zq0gwKFQUUr97C7DRQJduaJsM2sJS0uVE2iT8FwLlgzA
V0s/Mbjqn8fsUzbkcNZ4RWQ1yVz0wpclccaqJMxKAdjQNmVLGcJcZCc0K1+f+JGk
VtfgHUbQIcq6WtHdt+f5zduFE1uKd3e25XdaG99wfz7e/cHV9Y1RREzCM/U7xFPv
IxFc9ysW5qIGcieiea6Ie20x0NSZey+l3cf9tL2txtcd+L76NAY9uNozIYwDzvQI
8Akf9zxJ0/TpihAke97Xm2lYjYp3+RrHm/zp0dQ2fjVvSCuV+fCwBe9w5eS+gY3h
OvPwkQyLrxFG5Vl709KQBEbY205rPtSyggT/8qQE+rdzxXCZx20O0Ot8dkWt7QFF
R3bUIEe8S+N3aEjB2QyqfmgpKwqBO3oN3YMTqc+ZCko5gJrU6AC0dLMEUqz025gw
4Un9KdQ9ycRXrBKVP714jux5wl9jhKEEq0vuyqFBPEZGwn7DO3e74vZ1F4F9A/0T
Vv+UNS0ivCCrsrkSXqlikc/+5Q8z78mzlg4Yzv2kijMMmhRFSExf7jn3LI3MLGnw
Zugr5xJ26tIRV6UwmpsrZmffC3rI61EBl2L0O5rjzhq7O7bvbSd5nDXvVCJZExV3
RC9Cxm5qdtnHokEo2ijUXMs7dYRMIEeZQCNva2ecAC10A9VPTsLuDFIH0dOpRjxp
oTn7GNkDH9NFfRNzsFUIk4ML/LpGPJAJJVVBJTLZbpnbOZmT5gevb4uwn9Aeonqs
qFVtFCfXO6VVhOVYppwVDNfkzT6LRmBVc2ukclSG4SRXWyPrTw9imp/ubkir0vJG
4KGIhe9wh6UtEb5S/EudWQH3BtW+ppHmFfFI5x5+MJltJU7N0Iln0vBX65Tx7WCk
mAim2OZg3HBk+2x2un/7Hs9opQOef/2Ei1zkB+HaEbgvYN4FjgjoZoaL/9QyA/Wl
+q8MzC6Ma0hEOAJqOAHvi2pUnnKuHqVfTz6Ad6mYbDOgb9pjJ0lbUqeli71fCk4C
3YWIdaL35pnzNP/wmikIHtd15K3VhZ73zX+thovgj4X6xlHkvm2ahAioBQ2ULfGI
AzGbU+y6+9ji57ves53YkRtLiNorp4GpiYYrLn8bCei92V8zljtEBdsqN00COeuy
Z6DGlUEW/MdZ13n5/joFk1npRJLuxE5m6UMPdyknRosmKod+LvXiZM52pCgN1CbP
QBmZb52idQNypfRxk5Mpp8y24CLkkero+Dmf8DQXhGp0tCQkdbt+4j9JBlQsNadG
Xqk+3KNx0pT6sIBDYlIHZkikxSCyU72f07wFz1NeeRtGwtAxmDK+5AzAvrj7r69s
aQdiIcHCZLNa3JyaWtH+/DCu+jVeQOdoITSSlOYzhfrOW1GwYao0uJUEZnGJ3rhJ
LVwBnn8gCd7Yjp6aUyLwyqUBBA2uIUNK7VH0IZtE4R5UprrzbJEKO1gWV3JHysiz
IioRge4HSaWI5rlF1a+bjk7RGqRMDT5TmrNRBB+EhKh8g+CSvklGk0U17Z2tnhNN
Uo8DptFCFuyqF5i5V+J8XAfePnHOil/omD2VFqg2jo6BGiZqj3mBggITB/4K04Hy
IHwtCQ1Q8M1CyINT+/ACMM5umj7eN8qfBUJxYUJYx500ahXH3tEhf35XT4FBZlpi
/2XAG98sMo4GPjfl+oDTknmsQh3rzkv7K2basxamWIc68YRhHjHepqU5tPZCVZGT
AnJdb2PxxM11O2auqDi8kt9dnT39BeAeF2/sMq2r/3zZ5nYiKV5I6dIMQtsdaGvo
/Fzn90ZlEud0dkMr6Tyx2Xz0yY1/qpqr89KIyr7eDpTlpBzeQYu9WpU/2fS0HjP6
Lq17hPwIebzTMGYnZrSzjtxvZ/1Q2CpkqMheRac5nJtByoRERWv5+B75raEOVQmR
VWWQ+H+BtdRFL6LUiDNzZepzgInXv4EbAj/ZZEzp2K6wForcFBEqYHCyl5BhpKJN
MT7s8LX9li8kcIRRF0rPRy2HHZnC8iBWxRPmB8riF7j5W4ab2hKyMSjLXZaeeyKp
2fQU+25LArcXth5uc7KmMwDkeKweHDYCB0DYZoa2FEIPPiL56CX+H3+BmuP7N9LS
y9UOlneTg2Knloy7sCgvn5y314WdEg28gBLgg7WlQL3lH7sZ4J2Ai8K1jljG46vy
4BE6nwZcUPAQ2ZaeCJTeOPu7V0PF9+eX41ief1IxYfZIac6pjaJ+S/IklmsrhOhw
4XuPlSTyO5j6i/pV+xrALGLVvJzC3bsXiSQuRbWL3K6ZZ7smpy4gnkW9UmlnvlJM
TXgDfdPe63NB4pjD6J81IDYCrhrrQETmWj88AAk6jD7H5wmgvlqEkeiPPfHeTXiN
AiEW7eMrIz8OBPQRWFKf+ERMUoG8ydeSJs53739iL3UYxXel7hBSZniFWc8xVywB
8xIXJsEZRdsmZh02ryE8zW/wGlzfOmUiA3jSmovgkEhRG1/8MaMbyA+zm01gH23B
excVExhcIKf6qGzzBhKivsJHNCWllmFmzXco+WHM1OV8uQ0sG6rtezByoVsPRADg
DFYz1ZzXDb2QPNqve06DCtR7TInNRevgKmJFqHN+7tVHu915Pa49sTnK5h6o+Hp/
3AQ53vh2OHpORgYwJpLhrmy/mIY+Bd0Ps/+Crt2/61wQ7resZkY4amTtMbnVeF0Q
pNJ/1DNj54pqUXoDQu+90pjmabqTslwJzVOUMlpUjpJrDb/YDQ1PuCdzp7Z4c/Xy
o6F87XcYht5/U4qQ7ZLNIcEVXC7WNZdjdxkwCuq4H2r0X6DXvpzs6FPq1LbSUIkR
XH4l1TZz0xS3s9xzLRDJQiHu2E7/4j8J7YjsEE9eooRRyoSLikcoQuxBsmBLQYbp
yU6yvWRTfF9Z5u1Iq3RKi+jOFZnr9gXMkODrg9U03wxkAQaUpFVdMBineRSy1yfs
q++8wFxYZ/8fJhdaqHgDWjwm9ovAFxzctYLZ6bqz6U39z/aM6eDgMzlROPK1Bavg
DLBxhyaw5NeENSLbjk6SCTori6pRCNvjbVCLe7wvVTEoO1dbMfjVsbuURReuPkdW
9+9Pcsn0+CSQCFcRZRz91aq04dZWU780hH5Hg+6Mdf/6vTiR+tm+v98uLYkJQ7NG
yC9KsSnda7Mzv8dxJlk8sRN9EnNX5g30YQ/jqOImyukQPF61/pO02U/ZtiIE3NdP
BvLkl+H5kiv/iJCkrsrDyng6rdhpj02+nPNk+tMXlvVdACIE4DALIrk29/F6Jqqf
4xt7P+Xw7H9q+K4949tQtZQ6IAq074sNuZSHa97ctdDGOkzvyvOs93/8r8YjQYT5
t5Kg+8FD9nCRfQNHelSlvxGNRKTbbpMwLfBTVgJD/NUXnreJZzNZO8TQ1uAKdWrs
ykUPv0J/WwGW4CHDuui7elIUPzrjndHR3ewcl6JZpm3gFP1zSbZDI9Jr0LbfNIsw
Cjeqakp+oaqLJHXKp7bftzJc6soKD9aD43WTifJgGr8yO56fQF2Tu1TeOMwn0BF8
LpAgnn9uFXzb7ejhBuX8CrFK9RDDJ2N1zb4v3YuheLZHW/+XuKHP6pvJPcG1D8wI
BhQlODfOL8Dra6GH/jL7aV6dOl32L+hKNaEOgS90J2p2kMbGgJgkpSnXllOchMO0
wfpsYy/7YQONtuBE/80IpKiSHvqydGsypy+LDQ30610jl+Rd3FW43ZPDfetaC6oj
as6yjfvX6eODm9qsFNNc03SvPPjGEursQ6tmnif9PaDeDXn04TNpYcBG61HJARLb
sf0PIZDjToxrH+q7M2+xMci6hUnnuKd2furs7mFMBXWD3bOH3NSgN4E/B53huyw3
9mc8qCLkHaVFhbLtrVfh9ysrpym/nm9+EW4JA+XRkhN2i9868Ikt3zUtT+qKfPpc
A8y1wX1LRDD/029DUEYVjJedMvVdLV5g+enUDK2TMuwsQxRdQQo6d7kFRJj6ZGiT
X6TqEafNILwaDVXOyXidlEKxNP9zmybog6IrPJOVE7dmMhJzYUR2CLIL371bGSds
XXdyJoA3oMDllB4PfHugrXWDKGNYw8yHMBKqyVxJZk19a888y0oA/a9StKXaZxmJ
aa+58LZ6/aBFxYhYh6rVXfXdUpiQCcMLr0NPzG1SxQfuPGsoq6/gDbngN0AAVpwc
CWPfqlXznLHpZ+MKtAuJZ/HyJaYNCHh58T+IQA/eEwkQ+EvnjVwYVQQObh9MXm8t
wJ02bifEl7laZTAr70mTgJmilgRuiSwr1FjxnixX+6aFVn0660FmYHQmWh6zIYjr
MUAKINO4iVSyK2ZkANqcS0hwzce21Xh/ABM2tRjwWuvPenByw2FC6VpsRqDb4nfI
LJLWMsL/zyUku9PiKiTixbR+yIY3sJh7q6rvw1CFEJLBjnAfdTeJtxzOZqXaIZg9
TJaY1UIwhjzwsEHjCeu7UFPc7rDCp9eKtM2tyAh/vUf+M3m4AR/ivUuvQttl8RvB
irMmv8rov8aKxzct1+NsPW/RSN4R6BEJU2AFRUYnfaMKJEMyZRJx0DB89ujbB17u
3wehngRBArH7dSX1gloKap5QELH2q7Yh7iph4CdZuOd9ycTXdgsSKSGtjkOa4H7K
fGHTs8FVeZG/sWDsihNeJ1aYRDnZhAApQ6Wg2ognOfgILxbm9kq8ZgOfpECZzgky
rTVoPgcun/d7J/TIc+iKU0bLW15smh9G3cFkhEXtjP8RalVYm6ZqomdaztRw+I/w
mCWfUCU43/FdNoi4NMxwOGGrLNvHo6SD8DCf12JujebEarryTwuN/kjabCjCOY/k
d13zpTCqzShZXOU0a9/vMoQzNyR3yF5onplpqZ0T14GP03vU7LAa5j6wDTgfze5H
TZfS5kyC5Y9dGLYSAsBrXSWo1YehTBWcONZd+23ApYRI7kKWd+G2SBa8TkpSWOYp
l6ooXOWiJKJVmQORcFVVpCo3dUB75/LQHC2JlhBtRUQhn9XwBPhZZoHbiXz7P7We
GYlv3wydUv7HHgD2awnm7aCdCu0coz5deGgbDw6nxMrEr/+68z+1bcgQdN8YG7cB
4PWipjB1CDx8eNmvs75/sQtn9K/Zxapyy3alZTGaJU6TAwtbtFoMwYGvslHzNk05
gQQBVrmU4a4s8C5s1BLboTTcmFQjV0bh7vd7YURmm68zFYMRgOvEdg7K181jeG+O
g+QKnyd0IAZm3bRaY+K4ajFDP9jS7EiDE6FzF8x/SyYa1/IFYcLRtmA+KdQ/Ypq2
+simDZQxPTSu1YBTHisFPt6d7MbIpJeqURdjboKMHqitv7+Cl/bRier6yS6jaADw
DCEEPiQ5XtiHma3u48wjkw7fEOsvT+0o5NZBwgmVHh8a7P65/caBadHJGZxOBn2e
jqScGWlMh/IkhohAuvMDe5Ugqd3AFUZFm/kT7dDwM/IkHLZS8PC8Y8vYo3F4UGPB
XSm6S9CoTYZKeNDBtfDQPXvNPDWnQDfiR0VU1iAiXFSdq5jR0ZeVqjv3YCSRKmg0
sYPDpVD+HzG3o0pwLhjZ9qeWHySPHc0AEDjH/xSfSx5kMA60INN4MfDT/GoifvYM
Gsmjw8DJ5VhXuIpryHPd9opoX2jaMd+NeEfHAbTVboc2wDgvknFvPc7Xer/vDSu3
x+S/SMEy/6kJxFA5V9bSKMLQAko2QW7tK5fveAIX55p73yp5sm1AMdvK9hHoe4ti
hNyFrG+ER+B8HOFyBCcz+Dm0BZvPjFqAVUgz5MUK/7a2+YpaG8AkFrKKbS+izdJW
xA0g1CP8JR7Cp7N40ZAK/r+A0b5UJPQmGBYG6u//MQTbAA+uO6gYpC8KDAzdnuM3
Yce13WK4r5J9xLiTubuJCH3y/YOrq/vd86uMKlygow3Ckpxwo+EnuWeWQyEDNPkR
m+cvGLKM9TAEWr+FkXt1WWOpljqwMtrljojnCdwlpr3GQw8AA/JmkNmHwAipAiWA
Z6xxeiv68AUkypoTRMxhv4mJH0FTvRPUMXqER6Y7fH7hWGvBCnJzYn5gVZ4grpvi
Md701uKvMpVDrS05mdqHRhwPbT/+dyCbEsXX7Rlu/0VLHTlMlvMrHh16VOhgP4Dd
Ps2kzCW6Gy4S4SUxGtma7CoDoZRKDkh1Hnkuacv7+uAu57l6do3Nme4He+wQah0B
IvlmLFBtGjGUhg2sGxU7N7iG932eSrGUPRf2sh9V2Xei6WQIimshUPDCca357Sr1
P3PgXwuRYk0TsvCrKGbav1uxort1SgHtiNNcyQoPZEcRYCtnsx30Kc4IIc43Lffa
Uw/CudEl3OyVHA+Rj++WIv/tvpP0wd1WtoE6+g4yUJh58Gvg+RDvJNcStXvlx7LK
YUtOPrlfeQ8KGm3cu0h992JE68NguZSvbrJ4Bxrq+XN1+3ux3SVolmAB6wbe277v
O2DxfxmUSKSbzKK/MqQYBWw/y5DHew+NcXlZiEkW+g1z0xyQFR58hoymYQpdi1Aw
N/wOqQhviEiy5ycwiJF8QgSUp3Jl66lVusEOhoBATsAWJs8DNtIvanpcg/UlVxLt
wm5HJCid/s+P+V31B+TLXyC9Sl2RJCmhODwj6e2k3I9W1b7frnmJAImGJRxyNAL5
gpgUOapLucPwgaFmdit4AExpaGAU2dIg8Fyu/xtCHdsoj1ooMj7JypxVxXY34Y28
2OVwpo5SIEuRUTxWlFIA2TB++QoLze1V/NHrx0Mc9A4JVK/Ns+z08l/wpODZkd3r
lnC5rVm9n1dq/gYw0BaGuYZvMArZ2AwVfgWYEAZlj7dK8SWUzPnSaBrMlGAS0QJd
uNJ0IqGz3KwtIfqwYzFMvET5b1Oyq4hTMWR55aerywbqOuZyK4t+XWy4wdcRqiXb
515ks5NS/tmuCgJBuC3AnRY4JlWNjwbySlJfnQEfjpHFU8AG3xEoHF5+jcgIUVu4
RSAmDjFLySqq1SdV6WivD+wPeb181N2NNUrBprQJ+5WvLsdUW0q0e3Gpc84dfTpH
LYZVuZjsc64dx7KwL9p1EmtXCodhZXt6H47OF9lPf+Za9CWnjuzs54K+t6/HVr20
zBkNolTy8HfB1LisPJfaKx2Dbh119nQdFpxoZaSq6kcB+F6YYJl75477igXSvwG5
jGCW5Lh/J41GcmD8fLngc2YEjgOFWzZv15d1D+uM6FAsxzUhcV4drfiDO/LvLa22
7gs/aeA7J7yk8m2OYCJUG4lOnBT+7YmIacwQyd4Ki3zTOugABUujw35YLK+7ZX+f
PV0B2XGZ9/biS30/zdGd4+T4VZtNvvkYMadxP6YkMgNlztif0FVvyh0AVpZ4sA6n
YsB7NGdZfKwp50fICUzqdILNSwpkJFHyaFe3pnmPc29+IgkVOs0pOE6J6p7LagDm
r02ZTzwv1s8ls+0qbX8F4sJYRza8z9wJvg8m/TOH76xvAW6XQg9R2Y3LjYqO8GPa
yx8wJfkMib8WL+XqNqBaNrCjTWhTXv0xlyXWGjAkDRq5O3ZRhd18pvymByvD/5ms
goEuraNEvDqXVN1bXGehMzoVJxqCulmgScUbAHfGQ88NX9BQWqHeasRpziEdF8sx
GryCxJ4egATguwTzE6DX96ONzW3DLh/MzdtfDgx4wOrQozybSYUyjtP4cBEbO0ZP
uy2lOjmp01Aa66ZQyRY/con9nv1wadf0ZnZGFb/DCYb1t8sG6GdfB+QagDpEMjuY
nXWzphzniVtJNKz/rpcKRRyALLJh50TT3x8a/0D4TILrRXeEOqYd+B4AUGjF2Cqj
QxlXRkVPgo/WrI3TCASwLzzjBxuZpWU3dX4Mt+JW54M5vif1RfelRSk+paAv6rup
3HLVpNikMGPl1hFJr4+MZhmuo076L6FhnqkUwX0SbcxK7PS17PI5NbNiLwB4W8jU
ny8HnxJiC8ePAmnCy9OvxPcc7VGcKHjXO03NamlUjvx4C/ne1gYnNnU8I4ZZN108
KGLB9TANbzEUoqzmtxU05Um+0nRWYHk5zkNf829mc5SSv8edHrkqYX6hzGJ1WVam
Et72d36VMTXxT6T8xQpBJkzSr9wB13L4oeh0wpMOZA8nEWkZnvX43YEn+/SLssld
micvUP82ljknwHMoG3UtQ2Mky+o7SDEygh3rxinnRdrcMqWPRGnKwi8+Uvb+oUhg
FzcZFpzUpAGCSzkdqmQ28HHCneGOhRJznAtWwMAV9Q9tJ2fijzY6Eacu6WWbx24M
dZDE71bCWDv7fxCqIB2Y5pk0a8OYJWzMI5oSoXxJIcHqkmp7d034KyuG6/fxXV1Y
A8lZzL/maqJ3hzf+Nq6Lhn6jDoBukXFuIDo4cPnbGvUjtXkMLRkHlFTyKzgma3H0
aTxU+ge+/RLTXiEOA2QbIDXgiCo4H/UcHj8dRnlTgUTsI77/SOLjOXnsck4bqxjV
BYMmd5kLtWXhX9y2mIUcq6QT/gAH0rbNvJUoKmnPiEfvjJzpKtw5Diy3A+CUGrOa
4ZoXhYQwdWQ8aUqauEIX22bvqAJHuMcyh+G61L8uAqmWxkCqm/l/YFqBQ5GNaeQP
9Nct4MHoehwxAK+Dy1cYkKxfmT4atLU8wTMfQ9OfBfzbuIbavZCSDigAuBGs/aZT
7DUoyoMmE9aBQ6hMwCatqZ9yviFX7GZ23sFkX/y4+XlRrl5u1X/2k/3FCXb3ZRKH
cSq/8e8Ku6JfR1jHMzq0f/Cx0bhS7sgwQVusO0Z48HxHK/vaPBenvh3azBF13aVt
NoJjDVcOnwBr9CX8NKVWCAOVfDCYlfhqCuxs/rfwIF7yeFzxFHTphJ0Isxv2gj/V
+s/yUHmyfi/HLBw3dRl3wHmF143taJimAKGow5EwCrOQM6AmakLD1cBmdlC21yB4
silZ8m6YOwpRTOMCZY09tL8tF4T9/lh3+YeIl7U+1uwBTu5keYoK09eUOu4H9G2c
sPNZVhCKmLWhdjtt3gJcMAiiXWO659h7pIXUiekKtjGML7GSR9B4RN4Iv7kzuagO
gGS9Hp5KM6QXO5H4D5CN9fpgCDJnjUIHEIVZjWFCOxT0aNMNQza52imLonB9h740
/9LS3A/HYc2+xbWknpwddKXUmfzZlOkBdJ8MRcI5VBE96yhaAo8YPabMy/rgT/EG
oggDwjXovj4VDc5IDYQ5hFRB5NqC2IL1Qhf9fhTI2rhx9VZlgW+JWmtM4tjP+F5L
c18tTAeRwvIOZDbmBg0rXVR3r0aBF71iwbX8WFD4b1s/Lb7iWpz6WQA6U3R4jlI3
+tcu0Z/aZyvzAMTuUI3kkPBjE5FuALKdeA2OpZV0nWw43HL6r4DYa7jYWZd7u/7P
W3BNezJCrF/Rid/Fez0SANsfOeL5YzzjTQ2waZsjWlNw6Km3BvbewUcKiT7z/Ixh
blCzH5BU9002CH0FU5/WUHLDA68aAU9p5WYljskioz144MO02dqiL23i1LK9hR5L
V3cUU5YQY/98DoNL9oF2lrZoRl2Atg2cW4qyLjifgC8Kv8+wohLCqq1Q2FrUrCbM
JnJmj+c+y2P0hsQPDgY6oHBI8RaCmoaKXLP4Zm9igu0va6Jkl5kP0idV4rjgl5xx
2YAL4RnsIXX1/LLdDVWfBD1bWzPA2qrIALLvnzpK1UWEP0833FQDErt9Q0b9vQuC
6Gv4169KjJYDMzkp5VhagbDK92tOYMY7d3MjL9M8sA/GMXid63Yge4c6vIrBqTw8
vonF0vf2ZFcnWFwOdXFIy1XCELRnHQtge/Gr2NTRjTT3CRkY/MHoRPiWvaVvauMt
FW8eCfMw9lE3W7yAFhVlV7VoCe+6aLgSwgJ1u3pcMYoQPOQxc7OlK9nb1QoY38EM
wEdVE2bfRRopz4i0gRbrvxAAWhLnvrTONujndcstWfSHKcrXsquWrCXT78SVIgNr
bNytbvTlCTQKKk7+tFi9FaR8K3ErgoTY6k0CdKzQXTDHjkKprSw2YY72/2Tvkp0V
0BkWaavRaCpfgyuj78CvYsufgCe0vzpU94gmHTwQirVythG67hMHmXdc4tTmxbK1
Txi60ho7CtSKqWKpHk3oDmVMIxHLk+raDVwStD2tKfEPyhHejIY6IGMOx7XvdC3l
uWTA/+HK3JHJ/KqsPMhZ9oasuiOq8F3rIBMAUii0SInXU8629S0sDPrd6j379tBt
WWrZbhJWQay+6Kgi1Yml+ljcWSUr0FMhxQk0uh0DxqU1IsGLyX/LCqBu/vbIlJ+j
jwcU9uTjxiEDKVHiGy1s2wuqdx0WF/0GxPB52VlbG05mkY5as3UATO1vfFKlSgca
DjhIyN+EkQdqYB7pDM8TLONi+3rKTLQ12a2H5ocqPCWXudYoiSdz4K4NsXq/nwlt
BdnWdhVnHJv+3rpyP82Ub3uvYy1NACt4t9ETm2ccy2xqjPrruAfQ/E/okjglY35m
HrSxa7aMjpVQyITlpFSMDmvXwXvOL2z50kE/1/GMZCfPO0s3iGz8GbFl9RsHLntg
CpHlbfHGopP6Mj+88kPATU9mcPuGxNErLyu2rwlxwwy4Xhzt9EIWjUXcek6v/YLG
X+oPgrtnChFxpdBrpRxHvjrATh1/HVgZBojsz9/oCcsGogKIQBE/B2504VNaz4uQ
og9gMj8dmoDCDa60zx22WwIR7/oj8VS4aedLJuDjJK4Y1ypqpy0CtSrKUEA0JB+A
FW5mlbUlbJXbdelZkKrgn5vBgIDS6a6wRdBIIsxTYr3ovyVs7cVdCddtSM3Z32FU
s3shwoYZnXzrd0fjHb3cN7hbQyNbU+FH3xKJv2GYaxZVhRGMkhrOirQx7G3Zqqel
tkGvCHN7vdy46tsJXy/yW7gffA8S1pCJanEiKLPASTvMMmBX5KchXZ8kDBmJ5pFy
ftKat6v0pbvzy/eQRJNbZOuFWHL8j+7uIFG/YwHQeeIsr0BV7hr0vLPDMDV9JP8Q
PW7js2rEL4x5Dg/cD3vzu3bwdeZGN7NzJfmhE/EvO0iSxJvzFMUFuDFXyhMvivnU
YfGeNv/tBdlmkXgxKhOkOxeNZKVsyBid6KHTrajkIDvtPA/ibz+qtUeB/wNg7XcI
VP5/8nLc1BKx8GpbCJeNPOKHNl5eTo6nWW6w8rbIv2lNi3UGjaLDDOnZNnPtm6Xd
uwuw+WJ3GdaJ2JvOJYTMItxs49cR8rISYTg8cnHwC34EGMMJ2kw31lDWKvU8gCWN
7dn3ZfvCUbYFvSn1NKzN1cM211VQLNTSvhTAAqGVQXqRVBlL3Wu8Z9MdbI9/+rUO
nIuvorPBsjY1d+rIAgjDWC6PqMSBjKcXeHYDi2LjqTwWzA0VbnKtegR5S1sm3RpC
CTf2pnsSjftqYc5jFtpbKDw9iXKrV4toxLEVL8p5eCLTguHoUeZ1ixnItRZaDb6q
o/yd8ZQpqiftcUUAnNUjgOBcca/VXRH0rSqn3BTwuhiJ/Y3UJpTaqnZw87LTqmjJ
QrONSSmtZHKoIR0SSIfjr0XSUpqdI58mMZrowIIGs33ekr7pP1N/GeZComMOvGvv
JufG0R4WuleIta99JcJ1PnlPQv/thQAFTMuJ5OBCtYLoxrd/wHPE9YkVRKtLCOLC
1AIeKwQ2lOTUEOvX0gtqKaKGQAgOOTxBWI6bBtWVS2nuKiJgENWzxKQlwsu1uola
8240Zs2hJION6+jKvPZgoc/GAW7j0mbC0VpvJ0YCNLWZFMKdQG9W5XDLAcWheB5J
YYNDJH+lHCdawWC3GQ7xjVc2jnhILeG/u3LH/dN3G6CrLyIY/i9xB2heLXGXhlcU
racyzw3/U7C//hvj8iBUDujRpRyh6z2JNhcbFx4JczsLkpSTgNEpv+2DJcEiRGsN
A5AUe/UFv24YUVvg6iBHPyUyxcb9y+UWLJD0ptoqyZ/PbJDykemGi02ApdsvoBe+
lbYF7S7Vh9bSZpVBYf1tvGYlRknqGOtd7lf0LU5OW4UegJSuuQI+s3nZnuARrgQg
SepPFPzKUIzHeW9OS72LbJp9pTeR3HC6NrvUMN1qExid9W2Y3X5Q5Nnons5SCWhA
E/VrPJfKcI+j2/xpyMbo6xmJjdxQh1mDIlIEFixfTG9WgOzp0IqRblNkFE2XH80m
nLdGelzPtlsU4sWe9NQ0e1PkQ82SqXIrwQUm6YRL8v+cwGE7KN83DNmz50D9WhLe
6KLMXDBdiCKb6GYaGUws2rGF+7xdDXH2lAVKSlWd0KYtc5EaBMMxAzJ6qiRh1GxN
+aLpcVbCDbh4KNDcaOqsdg6q1OMLtddj+QKyYlO2ZfVww7KGXPnIdCep6OoGnqkG
bxhtLjUsdhGLjZq0kFfk9StlU5/a4ehofjFwXE+UWHaH9bnEUkuVW0rbK/UqHYHr
lhUZ1as9Gi3VSNFB9lSSWZUYnFsrV1CuZNHf74C/p7nu95/uD9rxqMGA0Dfl3Uqy
FJy/VPy7yrlPd3TPF1ZOnex1wtfEu9Q12ksGueVQNzeFi2nr5mr9dlWP3eyB8XVj
XhAspXL5RZDaGkVeqWUTbsmIsqNwax/SuQTbchzkM4pOC0lHqeu1XsxaCNSLBpHj
6M+rNVq/exdhQnYDCFEzgg73V4OcepRS4xQchgpHe4y6hQcMrDw1xROw7w6cSmgV
5s0FdV/4rVAPasc4tKC9512NGW0pLDFC77SxsxdczqoHoPmEApJ357gY5miIgbxT
2WA8IJ5koy7anhbQZgWHoMSzowkIAL/I+OPzK6xQ1gNNUhYeD3M/0V3G2uIUj0Bf
gVjX+Tx4cGSu3b5rPjlbmLrMq8KU516GDpgOPCxXkQYLzOn0uTZj6K0bF3lAAEfz
itUO7YPHphPXkm1Z/87iPyOXc/RHFIEL51tGdKd6D8iIUISmQChBykNrPKKW0DJ/
RkE+HmLGLgIehXmDhRikk04VhjRLw2wbq9E366V3OfuvAGoaMNV/LxPf29LiPanV
L0peIyIYhavBw/D9gxArXnjuDp1uWGxgXHeNo3Swo6kcY1E9YAXgwddI2b7g8SE0
VDnpJApbd9X+U5nnXUYSBTlZTUbZn7ZDlb8/s0iTJ+qZ1kTdqm1RNjbhVGFc7JbE
zQYbbNIaEy7M59xlN6lC2KAruiaMBDSHsvnhI54GhUN4C/kvjuXrYIGXGn1K1B/C
2mUCIrkvXFVUuKO1td+xsIrLMVtGjlOoeGqZOL8jJn8EIyZ6/WKW14R0hOyPCmvH
OWzcNPtEg0g7FWYn8UIrhqnuhxp9NBc/TJLoBjhsGb/6tzdRUZGBG5YiAALKzHyJ
pjKip7qHA9kt/GFHY6dEpEXd1ZZNL1O+qIzPSp5/Y7HKTWzKpH+SO/9TsBLPa9aK
TksCynG4Fi6CpuyGNhEYeHo/dtxrU+SNFhdWtHeHf7/STMhFcVnIfnecVeIyxSUN
YsVlOn8GAjcHCpcU2ISZ/sWEt71rB92D7HFXZoqL9Hc77k6mP6VyrNkS5J9qWWZR
Q29kqmiH99kPhSiTm+5RuGAvaBhugbUkcaOlHXZG1TwWf5Rlcta8aweZCemxZbtl
Ht+dzgvNt3Ijko64CD4Puz7Js99zr0tnQAr/sW/6h5mUVbPS3BICkWOQ+9Vzk+lZ
0gIY1xhXYAURgmyApVR6NKRnAj3DhlQBi9SR3cdtDQPLiLJd37lXvuy/VPrTmdmU
MuTGb/dylgusIN1bu2O1tZJyPbwzuGkjL3bPdo/31gIiuxXM5u8x25rBGczz5UOi
5wLwZZpEkVYqYZaBYOyymtONyHcbf7j9zPTqfvtMttcKTBZJq65BesF/snHXPFdW
CCoxlK6J2+RBP1UPblF7T5eGHKw/N3oef5Q52JyY0lx6K++gHAO6Xx0Q3jgFVUVr
QQw+ipoEyVBlNPbvnmRf9i4wGK1RwDwdJoADAgaPHopswBpe6F8918KjpRXQNIvJ
1mnMGEMK/RjYv7ByEjHwbeVIP4wTwwf3SI15U9dtznM++ySH3jo0yjICvycAtIGl
84NbCgduftwfKdDf5+gJZiUSRnU0xgBx04EI7bZc0fBxizn8E6AO3PPaJ8PKs+DC
zAGiyzCOVCw8z2LRp9sK8Gpke0z906pjj8gfRT/5xKttApbkBGzOFOBdcgIhWXpt
6oB5NDaIT6jeyMt/Hs0r+aqS92FqZcyBaKngsHfkFS5XiJLf8fxlZhDzsP4/0TQK
BtsbS9gxYFtHH+OiMCdH4Zuj9nOFj27Sh70QvN/cFUj1koxX3+e03pcHFF6mNOEQ
Kv8wD7PdqmNIHf9ETrWYy1w18j4/cphQTlt3XYy1Hjl7qW2kcxaBC1r+BYYpuEAQ
nfjLGtdg6//CzwQH5P46s4bsHl030E4YLG0PVBoT1iEWXgixmGmgt1iYxIKkpEOc
P829PY3VA2kK+Yr4VlSKOUY6qf95e0gWmhJyfuzkQnccVFDw22tJ56F5hN/c6m4l
RbR7FN4IPlMexaJGRf63lLHSn9BZ02OSVehRHbTqaXSiIpdTTiORt6zVgzutbRh9
5UwtPMcHDQfUr8qqWJ9miar4XXS7Br9QeHnHQd6feUj+WyHuA2Jee0bwbSo/j4Ym
GjSMLwjL1/AxIE7V9LDjdAdAbgrcFQGZJBRRJke4s6hSHwM2oECDaAR2YbMv6hY3
0jfHl8bzf9M2ga6F4aJxLdeht3w1aLq0hi33S3I8oLteTSOHk9Qe9125Q+X2YyP1
bCIzfvIosjG1RtAAvFc5fLnZ70O9lJl+zhtKTDrXfD6nGvEtW2pYJf1sAoCg5d9S
BgbyGShypxsaZd1rBeQlw+51OYPT9hyfekVpY+j3cy2L+fgoChk1TTLYHABOQuac
I9kEwd/vFrY3SGLjHfr0c/krCYBx5Oodlcu8mxzRP2ovlnP8e4mJUUbWXrLCiVjd
LN4Nm9xqr/ydUMpVMidook5PJEHtBX7w+4Pru5+/JcLMqSTXSssQwQC0OnADt8PO
qieN6hQAeq7Oc1q3tou8E+1zQmhcz00XjE/LVsEcy02aT6csu4/6G/1rz/zgzXwE
5jMXXWI09i9wLJYGZF0C4siGTtvmgQEpxiMQjGes0VPpUiFrrGwq72o83AtHhK6V
we2elyyYpr2uA8PvNo52o80JV7pMt/laUkOTTSt3r8MUk7esSPFgMgk7pdQc6pL5
igWU2gcCcY5sN6S0v8V2tY5kdQlpQ6tQxulmOL6klxspXuJHetuD11MYG+fBmMl2
IcrRpD5vs/xwtDm74oSnDT//Io73stPOpt8ODlaEDT5+VVIkl4zqcAmMJFKz5ilN
whBz056GinyznyXMD/2uAoD2Dd/nSBAVwcymoDe20QdIUocw/wwRbPjliMZE9sEu
m8t1/7O6PENL6AjQvtp+7hxPYjd3TdALIzX9XJo0yKplcUitrYL38eMk66L9VfTw
3MEaB0qIqTgc+KDl3Dvo3OCqF7/GfbZl6YDJl3Hf3JwcP/HM7crHWEDAJpB/MEdk
mF8JvS0q6wxktLZhgOLjJa2y9jfUAREUSxS9D2aQ/8ciyYvBT60+ARe7e6A08qPX
OxixkOM4CyIftkDtONV2Z8Uj91OU/ML/XraYH277KAGcZXueuXLJCrRVxoWHXje0
3aerl+4WNKBfg8uNzcWbmLO1UofVkjSYnmDKEMZSKs+rMb8PLCDCM5dEu7KyNLCr
/0HeCrNx3lGi4ApzB5CFlR/1uiALhCI2VV5eeveOD3IrRH9ktaJFbdcwZZH12rfq
6eM1WlzaAM74WCMyYSZBO+QKKOxk61wJ31p66if/LztLgrlbIME+Y3bDanmU7lMG
+SmMJr1DEvC7tdzXs2k+GoAaoUpF8B37WfVsDT1elHfPaso1d6/BbXx+fjC9h4Ab
/uDspwoheGG69gyv86py5x34a7XwCFzMCEZMYPBD2DGuTdUb0QcZmG3rTMA99LGD
encnJFify6XdpH1CCpgN4tUNOAqAybJ6PfykzgbmqsESB/JCKX0S2v4273oi1hd/
0k11IuYanGNnfu5dheDV2lIALCCZwZDF0att9rR2x+M9MDyGAjh/lESuuDmbzLcV
9PEW5sXKaciwaAiZYwumDi+KdSjtgD8gm/X8FVRp/hTItFXZFinyBlNrdluoE56/
0kHnfCNBtElGevyLc31GymDrdJSi09f8/XSN7GqRYAcsVMqoawC0WCYbPa+TEJCw
DN7vU5XR+Yz60oWJkBBg+GsCTJu5UDjZhWnD62uiqL6Gk6xOm9Kl1NDYq8lXl2DB
S7vNSZkGhWQ6yM/RqmBUk7550sjh+WLn35bzFePWiw78ckDonWnx2gSqsBRVd12e
R+x+zHJn7tUiiWfM269cnbUUNx9Tagw1zyajOxXYuJrfi0MHBDu/8hF2uMhpmDQD
8GtDktWEpx5B6XguL5JWapBD7ataq5BKv3Nh3M8mb+YCjP5F9S3QoMPpj12MuguA
IrgdE1cjxBtVJKnuy2BkeVfbcxXnH3vBh2OgheIb3eRiaMjWP20Br367XOqx8Q3J
ZxoPRgAZ8Lu8fAvbkBlD8jD0eMjbVJEfV6GB/hNzclSv4bjksvfHqWQ7Zmj+Jr05
/0G02IDSG+plIpRnOPHd8eKX1uWK98X5vX5Ko/CCJCb7LQsIxatERsZ3ktWJXbDU
9QM4xLB+3C1hmG7QtM27algwk6qSHxf95DD6nG2WONYs9OI0IZ3FlKvo2B07Kbz3
+Ksp/G1Bo4Uq9BJ+SaH7fUE6G4wOVMhWW6pvXiGPh2QBwaga/EE7+6eTc5YzRC+E
oAIB/cdu4nmmg6sk1BX5PKI/v2QdGc88EvLrPncAafhOSNU3yj1ow+D4tCY2oAiO
gOhLrtI9ClZjGvDcG3PUVauicafUSuaomvWmTaQ3kCbPFkhzCxPjGaYwQlKa+aDa
xZ8+cxMJUg3tkQtsJ5kjzJQrJHJlvI8h0VJf7WUpOaEiColdeNwgFbh7SVWZBbNy
+VDRg1BcO9jYfIfGLQ9QhEZV4YiT67KsQ0sErg5C3CercxBJw/orNS4dz7Wxr0Tm
HAAexLKfqX+p3ok1RZzfpWcrtV3hcyB9E88NpNA5Shwbj54TLgGZ0UM5jPYujClH
nm013Yz73oU8P8qvVAKIWWsIrzj80g3hPDBQmdFMfqInNXXrXoX32q2c8OQUhQzl
Mno6r3qIC0aGZgOOoQ7HVBxo1JBNtDvv0kWdIvKqDd+hVWZfhc6ufP+KEiovhTdB
Mg/67U0xZP/wdesn2TGecKdcN8y2WKSVgKhC2NiJ/yMDeS5z/bCAGZ5FZBzOyxxj
innTE+t0rC4ejmvp6Kfwv+mhgAaWtxNSkmG1iNd+3+ImdApthY//pEi4SHTIimom
LVDIen74IH0E2yLm/1Fn9LU13otgGbiGtSlrMnT4V1Axs4ERYe8E0Pmkuy2CR6PE
J3KFitY9enCfY+XqHcmJk0bHGXHHk0N/208yLhujuWlEbLSKIZ6vB9R5rsMZdqEL
h5YXRIyDdJm+johd6oAJJg5jwH9Q5pnVppzpD+xjgtRPEgma6tui9RkVJtZmkh4P
yrOu5WyXR9KFSlSuWxo19Dp+4k+pGbEJpp2mv21u2exVC8o10BP5SwqmcyM3nj8i
T9Q8LIsU+60YBAuvzX7gVt0BsORPrunPk1xpjWv+p6IZUSA1707HWUezfcjiAyo/
yIObm1BPfhJDzKFEl0PpkNusXzJ5ioaTVJJ+NA9nSqHOWUpwyNY++tbd4rOOVCDN
J3zMoAddUlE5tPAizrwKsL5XM4O54B9z0jcBKyOMqRwDio8vCk4X7qMMwAWcr2hS
yOiOBtJN6+0p1/NSxHZKBO7yOtZyxLLA2WZ1MRG/LLmXWjbvfs3bti6Ed/uQ1/1B
f9iK3KFwTETTQFlX9oDfEZS9Xzoct+u0dj9631WVUhSql75b+uNktpZ4xUVjSSLW
kE5jIIdR1WHUI9uF0OiL0CQMvc7YlwyQffgq55b6XG/ntG2s8kfUfkgc0weeADlc
CX9wivL5NAon66TYQYjdFBEj7TqHkgXyGqpDv4WmtwrNs7DuKJISLmTKeIHPo1Py
i2HM/naa2foHDaSEr0YASn8peeZewY8Nv0i/+PGv7tYyy4pYwU7ruLdNZ25L/LRm
NaghNToKRb6sKVxtyT7oxpoBmd151vP/iGKY7GV5C2QnLXC1sVDpG3dE737BpSvA
bRm/64hmTPm3dZgXTLw7ZYAm8TVlpGnoozOJmfH2Mp6V1BvKGs1wR8M0ZukGq3W+
gEzdrjM+LHJpBeIMDaTkMk4JBowLCzwO9uLOAYlFHhGxMmOE7cSaqvL9TgzJYSiu
Qf+ybRjmzlHnRbf9cYQQXj40rzKFmIXivY17kamMY0dRUENrkhFYPeO2BHY9LgfN
JAja0skysmEmyhi3b3mlsYYBPXTps2So6N+1e8uxiNMiaEBB3E8af1SRyRwOJ9s6
eCgiivNRh4S0nJPl4BiLs+NDOi0Yxebx+1ttXnSXgCKIf4Lpdszyr8+OhMjuAG+h
3ZXSK5KvkFDbgw2YcUkmrFU5BtpYoNRia2P6AbOh6i9mrY93s1S/2erbt8WH+uJf
yAbTmt7aoTo6qVdLZXmy5Wc0EaQrshe655+3thot4sNT3q1XcEtmTTWn86Hiy1C/
MwPPc5UunlvSEoySXm4RHdpwDSJeHGVz6/t2JwlcKimwCe7YgaiUvxtTP3S2udhP
hjZ61ijfeNU4U9wp/vWZnTQEpb/ZKCfq1M848JisrjBXEUAOb8az3buSNtHHJDBC
5VjT31Xfa9qDj1hT9ohp1VAWHghX4LMgH99ylA/ukkiz7P3C+jWrSI/mIlNG0MtR
Ddn2RIwgZYbti23NubMa+GokG2oYD4OCdnAkOy8T6EKfoz5EmaLpMhfhkwHNTDDU
SL2lOBFvd148a7PSFKP25V93tvCiw77ZE/zzRYicSQvPg0oUpc0qd3iSApiv1GnE
VMbSBIxWyH68iN5ZaoTtr5DY6tlATpYujhJ1O4j4osORpvC1bZgnrsnCTLZnaYy5
WfO83GhSy2fVQEuEa9StPxwKuCHRtfp7/3mtraUH5E9T3nPDxMPGBLrjzCK8LthO
Jt7ofYwOGLZq2OZh9Spl68Cxn9XbKc+SFnh+FGhetEcRHaHiDNbCMFW089+EUc1s
eaXKiHxOIuXHGylcWWcOG8jXHfsICgQQVPQ6HKIgmMMIl/OYRKUAVkbXKoymg6Lo
FHd/QXDJtIYC+q7DNpMiJKpnAOjFbUk0ocW2luMNfY26gTec6tFGvwlzU2fl877L
m8RgUdwDl12MTwORk04AbL9zeG3PGN4wUeGWPMjOejuVC7rZZUUMEKEGJ7OI7Y0h
ybf6mmLiPSntnV+qKthHgJVrM7BdX5wwdJ68Zan8fMxtuyB81Rtv/sg0DAKCZVSa
HGUfBUe6a7Tkaaj0c3mjVinC7TIyXgUwlAQfGRrd+7dxaSUdctmTOQD1gi2g1s2e
SNZV0ZNIh0K6NZ3ETbw86jyEg9Vn84tullDDi2f/OS5aLJMCSuWSOkDKxbZ1Thdl
9Qw+KR1pEaZqxN/C8syNVPYDTSPZX9lJyN1H3dFMb7ukv0lG5n3XfKybZU0aXMWF
khINZKHviKKEM5a6MkUjNXLASv+dmryHJ4cXF2kRWabXxoUw6oJ/TmsiUwimG61H
UDRpAqNJG4GhzeKPUdFX6GHDweR51i58ZxDSLmSSR64KdROkvRjlCSz4GxDfL812
tzOsCnxBGtVdSUNsEgpVwq4MQkg0DO6BPB8R5vm80elqjCM9NUyso9uTMmFuD/Rv
NWh9oauChJzUZ7drCoLJOqc1QBzNMDU37MVGRjFO7Z5ut1fN06af8GtoBOfbK/M2
IznCihpNXMKhHZAYKHomjLA3VRjy5lmgJOZpF5n9Hen/soYrkn41DNoASW0my6xR
C1bQKxeJ4UqrBTLKA1mMw2kvNFrAerhePVSkRzeg32tpmhNpxoyFUCM7Jl/5kqNX
4VgrrW2lbWHpQ9U4bAqCokaS4RXNj9tFsbtGCgEX6ngDWY3MMd1GsrH3ETk82vHL
rjmnuYWq43t+yBkMMjSBvTgB9VXlBSV1IHnfiiOxQxM3Xa2cqvUKNT6AgCe3fHkm
HD/dWurpAXjtynzv9UcAAiZtEscpV9J1Q5pPA9bheEQaneY+G8DhKqF7OKsBwFBy
zmbF7kiMZ1f0EYUGisJe6EjprA0uThYbaIC+Qb/mSqxggN5LKMUYD2moUCM1cqzP
liw3krexWwbUQNUAbajxosc5w/v3Mfj6/vUO1/AQoAbjqMkvljYFCwWKLEwvwqcz
0vGjEzfczojGthHTknDchzc8fLi6ZN3HU+e4FJ8PI+0qbIfRfzhM6cuXPqy+peIq
TUFYdrzxDtaGE3vDR8H0abQC6AIOH6opLxKO0/ofl/QM8FZXt8V7pcYIb24Ielwu
wYaSRI2jn1wWe1Hp0SIpElv2JHUMCk3MBitiYIeAM7NSaNWCKnDFr5odXFzChdOH
+8uCUT7uZqVqQDThSbbZ2MP/ZWC3FeIPzXu155bntiS6wTp9AjUlrYtJGvYWjFVP
k/478n9EI7huOr1l/1IU8PCnwc4frxg9Vxh1NnCaDp+611/Xhsd9pKEo3gEgOgPy
6WHKRMf6l2pt2ej6igZ90GJ3HlDalB/7k+ElY9CcbiAjCIJcxGCb9nJfG4lNQrcs
+gL95CTa6AcNp6ZRVHx282F80twr8w2ezqFKu3LzfbzhLBAbcvKZP9gsrtosPbCo
9L9TZHtEB3dI/1Oj+WoZCsZx++N+z/etFv7Jn6ZV5nlZKiEbTq/LKJbwiu3QQmuO
bLzbwfAI0Vn8Z7IQZDcK1hRKqX8GF59UsTBUiKCDEZgNt0iduCg2iLn4AC6Eu/Xw
sW4sxcI84IvcinzC1edJhubNDVeY/y0HaMGOslkE3qwa9nBKk/RxTPQD+IRF/m6B
anjnqIfucDlsLgyEQ0Cuny9s2LRY9KT8yCwSM8C9fOMAzm7AfgfY4pZYPMUGKVbj
B2u+vM+RXgmJlUipLYhVOuWpUUW2UKdVRh1EkPjDmBv9Qaoenetd9wThdrWC3aNb
UasWSWoi1i7F9+Yf4xg9miZy0n6b8VaMvz/H46IZNWAJyn0Xvvx+BqsI9vZz2GrF
LRlC7EupR+JcHQqDkGDMHfUea6NqKgkzINKUOJY6p+vXtKc5n6wUyVPFkUhvtobI
1hDlYLlHPOwA37WthZbipczflkdC0voT6XIlsDysk5vVk+3/7uSkpF2YDb+Gyguu
hiithtuh1Jh82DO2QgWp3s+WCD0X6X8rFnYqTeMZUILYV8A7oIob6ltDTaJ8acb5
QtMTx6NZyT/lIQ8bTTmHGt1G8cXBUEYSOTYRFUthza5qXCgUQT5wGOGrp8XnyoeO
qKJLu4TQwY3xd6IdrnGtSZzzb7smCZFi2ubhQTsrfUs1ZxvQXd/fe6yTRWK/qq1j
EGzI5mx0qu3v/fxmbCTrcvksJ8sHfqONuM3pIj3vMUg5Y5qBKJ0r2aEnomg8kgj+
bPV+F+doafhhi5/iU4SHZonm4uhWqBrl+wjlXu+2Qwvbb528+PBir/sctbnDz6P/
vxGJ2yeayfI8Hcwg9fkAa8TnfQeBV80RIf1oSygrIOoAcYnxBJF4fGOO5GnhABUb
iTSVLEfgSsWaWiVLOyVtQ7kvcuiJl8ucc7jbyMKSSY9NLCA8yJlFgP0qLg38gR7G
nYOtwW2IFHnQryXEwyHcS//ZtqAReMeAbnVLhyFh2Zzk5Lx4AF+uVfG5UyBOoa4A
CEFZu1NOW4WQbS4aNdnA6mqkeHYRjbbTY7OIZMmSiIc6lAGDAHmVkpTF934gqjJj
NM+H0naBHs9iZdqtlAvWVFhvQ5h8Aw/IaOjnZCSEXk13/f2bHN1irXt+u/56uwf1
NLhk9RnGr96aJdtDMBplhgfzTq9HEKtEnu6DHfqYGp3TYCotoaQar2QbXjuy+Xec
SX095hOz2jHU3z042F0tc6WuO4whA8L/JkpqvUQnfzdmNMr7P/PiL5fGQBG1n45N
wFfxEFeRMZZiFzMSLFS/XGoWq/w1vgazN2C3lvsXDn+r2YN36bvZBnG6rAmmG20L
k0CeKgba0l1PEGKrja0mWyFqJx1nIQpWSfVeBhWQHxKi78VfljNNT8UZL+mIcZle
84fLX8BwBeb4yvr96j4mwJzjF3NNsLe7xbYv0Gg89JKmJmF/+pKntEH/t0zB9Fjy
qqTvB3/nEpHPZj7xwsKPwNThWIEjL34CGSt11TK5cvJqGv6jyzLUzFn9kHZ/bg4A
r3iuB+adPUSUJKaah44aoDMNY8QIYw41fNiWVhktF3wiC5FRZ3Q6T6uf6P/L163M
RnHCeFNqmEbcaKaxZBit+tjgqM48pYacJCOqKZHlWXPrUCe6cDVWFO7SRIyX2NKn
WsibW4OtFlP/R/U0ZpWNFWbhzywRbR6Z8aumBrkfH7rb98ilybLNxGvoXdA2cCyF
CqLYakcRuxqX0q8atlKa83k/WyvSqselCBa8K0zhmbqf6qwo+MQ3Uf++4gWYuySM
L6mMdffpx4db8caRVaZ4lbibvuZCW7PLWdZgF+NNzHx4aXQzR/sQvxFUj0gLY2Mt
INz7UD5IQYODSdVrMvN3Axzla2pwoHMan9knZjc8/eEyR5D4argD14MrTV+yUVY/
8bMqe5wyTmqe3yZ/3kC07uFXWALnLqMjyJGoF27I37Dm2l7rszrKkxcCVtss1g7W
E+1stSJRNlxa18L7OQGIE1CdsJ8TB0ulRjdBsj45y4VddesoGNI3g7enpjFegPn4
nnczB91Tdjk0KbJ989b1b9uVUZT70NX9cKY52vd6ULlqonzDj/NsxCaOWWpJovem
oDCC3dfOnVDFHqy+DuL7CC3J5uY6pdsyIbaJLi+DvDrxvYWYdvozi5GHaz/t7+p/
G7W2xQ+kobBUBjoDTCw70g81n7Qca+G2kXwvTNH3yig9fMVmYY7MosYaXBqWJzhF
wXUrsyMVGyzSBnPATU3n2BJmm7NxUEeYX3MebT7x145hUk2jioaxClOM81xGSOm3
hcfhCB4GsTtoWliXiQE2QXfGkCUuToMUI3E0rCBoVjpegdjvUrbz7njy9gFm0BQh
nP1Ob7IVomPMR+bycBEXGXvLyD4WcKrKkwTgv+UGh7hg/u2AHs2f6GYETXg+qQ95
P9B3SXmfcxxujrCN73pbZb36Dizh2eUU/5YxKuEqrIpfYrqt3wha3rKSayC8G+Y+
qcHDUPx6fHf2bdCpIIp9U5T//yi868Vm0wWvNs1mID+Q9RFYtEwBaWjiz7ZbJC0l
HDAikDDQDtTeefkkeKeIuyaVlCD1lTawOucOSCNucGvLqjkKBEGDkw71FZR3JxqJ
nnYyY1blXradda3vFwYJ8ZHGpxBXpyaz/zETZz80YvGqz05okD0or5S55t77YZCV
ZJaUh1P1sUTTHw32Jl8oTfWPG+s5DAD5XkpRK5XVd0Xg1v6PfGekfNlrwoZ1eWjr
Yts+NfVTZaDpvKiOMaD1zcudn2P9OyRof/7YvqQYOc/KkB/h8ZQdf2RQa/tPywMl
CXuH+jYOIb1QZerWcnY8hwTpbmx+WDgE4NZUkmRqMfA9i8x8UA2Zhvfv74maOn5V
g3466FgoDk88MQQ8bBD7wR+1GLN3XR/92u/S6lSf2yHngmIbMD2cVF5TJI7TkCGl
bpDkFD2L4ga0VpkA03Dxb4ogbNS+fPP8VUJbMw4Qv94vNBuUexayw5nj3ZSKL1Jb
48XpQqxjFy/vzsnuxzrgRsE2Gz1R3QjP/c3I2Ds1tIc5csmW6vKG/5YyVTjsAY1E
973FJDEVqmXnCo4wc1k5zlrSTnyFox8CyZ4//rXveqZqnaViTgeVk1htu03WE+9u
ki3mywtA8Mi4cGmDfO6VW9UhW7PZYtGNMA1xO6PvvWNI8l/l225tXp9DUaKN31yN
DSIsyoO2zEnS1wzLhkCtEaHjiDFhWuc9WQLuPB0CYgbtY6kOleRQQen4C4OPXW2j
OB0b6loGTO5CEVswz8DN99ZrOdS42UG7Wy+Gv8Z8po2zDQONwR5b+DIGi/W+pdqm
sRd2nevyjzB7P9FdgIu/mIFUe0msv8lAH1Zt1teH2wURGT92woRbMxAly1beVmh4
OaRRROqK58UDO9MsvkOyiCJmtOD0aytwnqm44ok+ANPIz7e5nh53/jmGo5izl0bj
+H1BUbXzl3KFQXhootoWbXfzyL/khrsVy+oT/BXQaOTxgklGSTxF4PLkJBcnBULj
+OEsvKKVicOBnJn0I0nTCM3GTpo998DfQDCgUZZOJmf1FA/pg7dPlgSalC8PkhTY
Y8bf+IlKfDZWo47gr40rAowJOkqSRBfzE3nObqocJZUfy60Ss/4XRiIx/Dk2EIuK
5hSnFZrusU+n85BIwi65cOCH/YhB10HAnTeDxTBXmmwHJ+XJcQbBka1r+T9KMILW
a9Xo7x+JXsmOsUxFfaHk4xBrKex+1lyLxCBsaYUomAUYZVt3MSeSl8ql1mb867Wo
ggNWocow3uayLgD5Yamw39rfTOPN+W5q1an2Jw7YOZIzc7uYlD4c5N0M72JGuuZG
1fiTweCW9rP3QjKBdKMMNDsMs0d73QNydxtCVlIPICNYPE3bj3nxtfdgJPvaVjGO
bL8GEUaBBOW9jRvk0B4S2TTC2rV6bZgH6EoqNz+VkTJKgkmSh2RRltNwpftZ9bn9
/t1+UAcWSkJd5fpeOz5Z+CWeHNze5RfMAVsKGLuZd9y6EX1ftpRgM4RnPU9fYUEW
paOMzMYKK/aHd/brXQqt37H7YxWpUUAMk4IJVcRShmNClmoc3M5y9yDytGx4hXEF
cq0/F8//dx9JLM8v/czno87SXv5jFCony1ZqhdfeFyz6WFrpIapTMFJvUC4pY2Le
1RMkt7KBcSl+HU7qaBWOLd2DyG6p3MaHMbJIMlE5OxS0F7cNWAO1rMu+u+0z5Coi
ykqtInJ84ZD0YB0VzILjg42ncKVsCgQmGzAhlBVVtrgWvDSKT4wSGqkXSFd5DPUU
UlMoPI1E5B/u0rb7yoYF0EGTkiDTjR9OJrXHgxpiIuPaMgvfrYvU+b0k0vHQvwsK
Z4jxcw60hjMyfNRDvvxx8TZfbt7BQ7LEnTGJRzAoGxa0U0AQ2FYlJxpG98zaMNWg
Tf7TDxrVt18igkN0KNa+BVicZx81m4GCwGKf8vBy2lEXQRQK0Bz8BfdA/GMfPb0W
eqmjr18EmJe3RnRCo2fWhAAk5+aaRYbeE1Gx8oallXn8Tmh09/I2Cz1rgcjLtDPO
qHPFftcR5lA86LGcbiI5Fz03/TqjZCLBZUqIXfcO1aGRZ8c8HSbMCpzD5QcQbb+D
KXTrdKNM2xB6NNwwo/8n/H1CeQLmKQgMbZQ3NSBxL6tSPZ3E/txip5g/UZ968jwc
pQPvN3Koo5LWcWYpumQY+ESpsNzYQBvlSP1ncrsyprGxBnitBWS61wvXc1HASrFZ
iCkavjCpyRfPqFpQJxPB+vqUyrwA+rlNnjxO02Ei9mLLnHzHJUTgvu+kZ6ZXt366
qpUbiZdIKziHjcUu/0UfLmPNd06P3OJ77PGcOF6NaU/QsgZ77VjLTaJNJX1cp2Bl
TEydC6azg5wgCtXKekm3v4b77FN7tU5fkBTCsiNj2+Ubku0DFVxeun3Ypjq9p+Kx
le47ZjjbPTvmTq2vbbRYTsTyZG87TVJVyCVZkzwsJ5dA32QTCIUug6heEYoKKazf
8n04s0WwnGCBegohVmCYCxFCboxa/3r3fZgHCzDqhcSnsfFpQB+PlCD63QyWpNrT
qCb5Im+DS97ZpBw7Nqpdmi72YdjpZDN6Dp5FCo9Bo59OGjH+fzbg+1ZixUNjJyJi
jhS/UPOBmkGeqAS9fgZONSmKV3Mv4ui90wJSH3wEdRxYBu/4WpqT412H4A9dhKl0
QXIC7E5Y8NtLOFh+ITrPBEz/My0mREIO6asLxACRhGYdM+w03OBHJHIsKtOYcmis
/nVktS+ymcMGun/6WSRq0tmVlpJy8m8FAnGQGSYAKI+ZjjzjgZHvKXg+gtm0KBes
CrLYj2ewtEKSO+7/P2IQ/44ZVwrIgo/ETV91yBYPuItE7wz1MbkhSglOEbxkG5AW
SkbxHIrrVFUHMFV9gJ+UUp0EILpr+QzxKFk2T8vCQNK76loFugUt8h+/MWwrBBXg
+piABGVDJoS0rysyAneTJdto2uTOPcnhTLZiUS4ubxadx3NGIZgrdHakjZnpk5b1
H9Z+UyPc/X7CMvLz4auAKvzqrUy00X/kkaB2FoGtKoLEEx1pHPhqwtTdSPFWt0fr
bCgZSApPUpp0MRUJ1J2OQUPpB+Qe5AKVjsER8n9tBw822k/nJKLYo2MBrseHHdGT
R87xZuGYkpu2rcIYBr/vjKR76hFyXDFHdd9zW5DRlytB6IZVTg8IwMBwjcxxq+ZI
9hxuBYPEOAZN1pKflW/HD48usor7WSc2nfZkb/5vpYu+EPQZ/bTbu4U13v9v8nSi
63VfYKoN2njXozHuOXLvrcDDvCIUI8LkbhwcAWrDSop2gqJjiBhKgXz8s4dVYORm
bSVPfQC7Af8DvZKM/2P9MLRVQZD4CGtgsH6m+Y9iC4SNNY0ouCCeQpoHeEEe07x8
hnbkNa9pKDfPZ8ikuhU2e32scHsSd6ZXekms3e3WOfBilpzUt9hGt1KjfmC+qe7c
kfkRT3FH8s3HiBCcDc4qKGOK8/FZQNWbPP7W3AaWwZYei1qiEHeTxIYGMKscVyzJ
lqX3LAkpUwFhTs1Kd3u3kdvtr85GL099IuLqEeLqqeOirb0nyo+ZvX+dUKQ2pKEf
xbw+FnN8XfNMLugUyR+wprWKc7bBRuAuCz2oh2ovYp6gAKr8az2Rq5cKIK3cCakG
d/V0Txl9cga/yHvsoFnhiasKeJK2az+scaaR3QNi87E123tymw2g/wBkv4D+tIbU
GAaJkWDLAukBl371X7VChG8F8zAh1AfelVCuL/jxeBZJ4ckqsaa3yVYhppVhEEYc
vqSk9nSQKYWxh2tZoSyW2qiZPMfOi2p5mJk7T981SG8a+dAJpw7MM0IayosVIvtw
dzYgDSyHjTKv2rR97NHsdfy6N7UvzIuZgksshZYKnXw9DPdXE/uG2pfcQEiW/fU0
V2mHJqS4GH/SLcU782nGxZkWLSSoJ0xd8reNNtybDhGeX0kKLGq0adMHLQqz+Ko3
j98DCQdpxM+i2a1PKEhbDqnuRAmuHpuhPFDG7cGiHPMFgTpWrWrBkg58H1zbZkNa
aGi8OO2NT8lT8p2ulwpDGlr66wq4SzUBBxLRXXkDYEYabbKsCXWo7P59sV5SkbNL
lDJxm69JAad3q8EiP/5Qff9XHmrfDtYYvgla0bwcNfpSoPVqrVsbp7146kTN5qbp
K9gZcjxY7bHT4G7JxqLGy40iIi6eifY1QbJnWgqwxnPdVa/9FEKvitMTpDWcmzrG
xNnc8H6rIXrKKJ9v8SQEB1ytqIHQQ6YgO5+qNdmoO9fHDeGn/TZpc2Hyfkx2JHK5
YjEId/FIwHNRCarFIFeGUwnPM2sM10a6wtYZX9c22t1VsoHncfqyAASvmAdqcsdt
f6TCI6/mo8JcmXNxodW5T9M8A0ejVBHbYERdF5ZDjzRi8LRDBl51gXgykHKM6zgl
8wFIMVyl4LyjI0cj5TsZcSmoOGWRJqMn3SRE6LA4eQ8+ovxKX+PpXZ4LZ/HUXSS8
R00KUoAB/sD5eVQeYj2GnEuCkcUnZhRd58bbQrugrRNKqT2Aj3H41ZuJYjkWXlKD
uLuTpOa7QonoEyCN+2fsQJRO/oxKwGKtJw/g6N3u2SchozcvkbNcUCmPou5GIjAI
sIbJLu1qA8Dc8EBpIP8qw4lIMwSbl7nFzhTNgTMB2yoxhAy79kZQumxPscXhSPPT
/jT2GTauiC0+MhFKDzRmTagly0vkaNeXthpK59NzkSBl+B7oQKmGFbndJzIdKUrX
LZlQsD9NHP3qcy0XK+FuogFT3R/exynuYHrjk7g6lu01Z8212Lz6lX+Bct19vXcl
WUZk6Ak+9by+/fLb4Xhr13AhqjThqOvrv9ieOTNGDKoyaY2d/8WQBcIby+MMrDkD
wmL82kgpdYly3+uK8BMtt8NTYd0F+Td5Ed9EjmoXCzQsBEl9N1FSt1fQiwS/gzrn
2kWtLXrX/7RyuWkn4ek+Wrp5TXizH2w3FOGX4XSuYgn54CUHtuJ0ZMzNy7ssV13C
Ifngd+53nOWoCgHOiugfF28GVBic3gdSVqPKKFHto0QhR9dLOGkLP7vid+Uq22wI
x3zyPKBroS+4Ezgfk4n7rxreyDoNZIhfBgrNmm5F1PK5BweONMGNrfavKn+EowYl
5bGwbw2fcC9mFjeC/lsYemhgRevz7F4WjkdsGZtH+5sGS5b4GE2yIPy6SpsJvWrS
CMisKiD634rogRgyFEsz41AlvZN/qUg+GSUZazr1Hhc0NLT2wSCMOiG3u26jiFWO
lf0T6CkxfOT6z2A5nXn7OlSkMml5jKIGg6GuoiSeqz1e/safwGVMk2MGCdo2uHyx
dRnJI7+1NqlCCXImBl6yzEtWG6j/y7neRXSqHiwPiar1le/qwbwWclIsR6sTVxqZ
zf0UGSLQWY+BObQJE+SS/dKggg87acdhmYElAUxqkp9hWjoBsXgFmbj7DXpyt/nm
pKJzNh3g84G3SL2mTU46wjBeU4Lzr3RQefsWCCQuakiU2EZG74f8vXrLhHd2j/dT
O8RDGTMMt22ixv3dwg2iGGEsfBTD3duScIAy/spCFvJ/lijijdkMFPp1UfIo8Y4s
KH1kQ4QsGFmLMVJ2bxR6WkwtETo/EiTGnBeu6fBY393TJDVG3wT4n4IXndREEx0i
jVWJmaDu9Ki9pXTgaRzXevyN7b+C6p/QWwPiVUcOJ2HwSo8RclTMalKzzxeBqKc6
/8IgnX3xeZbXtkArb1eTEm7FDIIo4I8cXT/pDdbLippdo+Guu1KkhusohNV2Nstp
/TEEOsAf0d63N/frr9XmCcq0lPxRt1AHuceItqL8WRMUol24t/ePcUxieYobLfPD
vaFShmPf8as28l0jxiKnxM6hC3W2hlSUEPsXosS+pXx32I9jBFB1dpCFGx8W5eVU
2ozj2PikIgC6o+RztE9WsGg7x6qUmelx6zZ2QyJ/rYorTECaP+jET2sNauT03MOT
v417SPRE3tHTxijkNzgXw1BHpEn2tEQ3sDq9MtJmBG7c+/l3whEcMbz1nyRedvDv
KkL8Xx7KdzaMg0w2nXs+n1AxRO6Ihg4hoI4EqSKt6SNiqnnbnh/hEErKm1jd5+0R
tq2ztdmo/RUODIZ+MahLVuDrFTmjqAsPDB46C7kxa/8FBS040C4qeoNauHXk1cuC
GK1M4j8Pxq+aW5RTDAdkqXhnwqnL6dQqHDIC8inDn1LoRdXHs4/YjZ6TkI5bTF2S
nswhQe2jK8KoEhZXzKZ/9uTAS/FvlrL966HM0v15sMgis5xcTDkE4BwHiteAp8hW
jVVqxOMwh6ZlrycCeLKUfpj0t30l20OBdKTp/UqlcNclYKuU7805OAAJKZ0Hex/9
sf5nD4K58mDfgS3YIUcLHn2Ei+38Meo8wYVTcpRXNQDLiKwzfrtiz7Rm+Wsx0HMt
OD9RnYLJpKdrxdY3nXPc7ZKdRxgIzULIBKlbvWLMzIYK7uIVzcQ8gl1lu+bSKwLC
u/4BuMkz1sR7u4H5S1oMiI5bZdHtSc3ows0CfMJ8yQH3IIX+fRFCeM+i3nBBfL2E
ylEnQHlxxeojeK3OFRgU6sW1CctSfQmwDncpU6VPP/G3WIxv/ybvec8hMaWBzEc9
yDm58n1sSNmQw8/JOMLBbaaK8/9yy79EjJisd0zlaAVgMGswI+ltENWRjsgHOyva
qpNdQViZ9MfqVbK0XWcy6K09aVW6I2CLQvLzlMUCxDi8JTxLfkM0kUxgkn3XJEDJ
PZ8WFcRP5qP2880VqEquUZvG+zmJI3YWdaOE9aOAfF9b8iIH9dDvCS4YxpbqTUs6
+WdX4CiS9caKv9p2r0esTCB+hqhl+r/Ew3wd9W7wWKB49JStKdU61Lziz73kKzQ2
v0brdVNJUH6LqEbJzWR0O492993ai/fztQSp7QqNF9CoNNUDE7Va7L8aoALNppPq
iVbHA/4hmZjCFfhph2Io+uky/0D5VKeB+zp0l4v7CWlIDaNvnPXnjSNfjskRVp2q
avgFG0rBD5CMGiyeDfM5YtrInXYFMfqpM/T35zHI31Mc77TS5uoQiKsAyB/9oXLP
cARe4ckPdaIQDJsYaVaX0/1FMWzmjslskRlbJmebMIv8kVZZTeawVWqf3yFG6UGp
EYN1XRX+SACt/0qPSwXW+DwiSorAe6EpOLrYTRpYZnSSlTM1XLEULTvGfjCHIf/3
nKkiGHCXKBlg2+LsUcCTQ7j3pNhReIa7zTObqW28qOB3XZijoN5abScj1swBCn5d
vF9XslXKa3XaZvXlJYJSkl3QL+syqENQMu53cux1vb/vQMtLP0KyRDGww9O+Bqcv
2wj13L/CXmo6wCljStQDhmL478t4TNc7VGwd9ZLyGFAqjZXH7mhE91BZst68m0ND
IOLAuMsdz1Ybfl6oZ6/WTm63zPEdVQuGbgjk8g8/7U5wFVcf5TcAjzoARfWoc0pc
jr8Xth6oHkGGABP8XqdXOoDeg/doHJVF0X/OGXf34cfIg7AnNQ7pzg3zriYfgcRj
85xLzvONZtWQJ4O06No95ZZ3AhggfjY067MPBIuFItGwrOF4GS8UCmGbf/dXUisL
DfLG5QTc95fHHVzKfMCvKwfpIT9sONF70GxRiulVzpFOPp+aILhR4aazVz//KQuO
IGg4uia5rlL9RwRNUFlGOU81PH70kGjzeuJ4EFM0wYJqQule8CHuDVlOC/oQ+B4B
xO5oh6G/EcjhLTO+gkdvaltXIVs7FMoc6xui/LcUUIxPIJW0M+hfH6uS2VEMQOPG
dV28iYUQGPydVeZfbsZJ3ogVhFOvDbN1gtqhc2yg79GDpeL9f1ww+lnViPJpmaJ0
nJ2atnlL9tSnh7ksv/4midxG7BEsdO02bK8M0TN0Q3vn+xYpdpO7AOxsBSU12YMc
chBVCQxHClAYbMwJ3SHpYFU26A1XGaKgM7sW+1feQhSVqcxsY49yFONe2CrcvetB
ry5u/z3+81J4lJxioIQxSNUDWEHtuQ6U9EFXN6m5TSmiqtMDbF+RsYr96atdQCrO
gZapbcPY7NGWzEghVIRDb+zE1k2rkmsaQMiLrzGTq+ZZfZwzm9snuO/YYr0wAdoP
PAwexCrrN2Ucnfab7LQHjjoxjYLqybsrpTe9kqdijdpRhFdClOIvYTVzfqQku37q
uvF2fC7PdNqQQEADucMIIwlhfB+Wysjs1xyJERgHuepggozTbRF7Q2IBbM73y9/i
htMkzLuXwauagH913jGly6zbICEC1MWcwGvTa9EnhLN5wUT7S3BnoX4xp4FSWWRq
6LrFmEPm/Qxe9RG/TmgHPhuNEmBPAgCUVuEdH+x4Btm3XxcQUIeW28xaSm7shmzl
58diTNVLvu0JqlFJhBlpiGL+9KlDQ4CXiXtVtt82r8HdQGAMLA6UxwvDF3ML8i/y
qkBmKTdPOxP2DukDBmNI437DvEhCyQj75QWqSnJctKx6FHOFxwjETgfSh1n356aV
SfEjrVVoMYqCxA6QMB/5tMQa8h2330OJsPqqUDflpCKNkxx66izQLq8C1Zld1fhI
647000ckH00r3IRa+GGA9eogZ+8v/I+LVqhyrHuCb7XrEV1dgsUb/2XrDDfudWOz
a42JAtTyJsz2aSaZpRGF7WBWM0wgvzNxf4p2J35zOrVzkfyrmIDURCZdHz6EGJrK
Qvh2QjyyWQdwQyFj7Yznk1M6gVxPfDBlR5/FeJSZPyn5vjabvOMtGfJp/r0vCyQJ
OHzIZQyUUtPrCpqmsoHDDFKpQFdQkHDYi+rcZLrv9fDXSPvQDdcNhkHlLnk0PQuT
JaH+qbnJYvNCNUMeL7f4pWFk9QO5rc2TsZ93sd4slZmpK7xPaO8dXRo5RtozyCbF
DvpY/1dJAa50q/BvpaJUF5JOCCam1QfQnBhNgSuseZ5hRnGUFX0zLmF8ktqA7wKJ
BDrmDP4EqfifvPtOfQcEGpDO2b0JkAb/1lSqqmLxHZklOUzslTsYidH1V0KGaL5W
P1uXffZpMU1jxSDR6DUr1lGmhgSWnGchdIKrsRWwA4BXo5NASkO7/HBfypzWG0Mz
j/aPlKxBt6bqrptOw6Kr+meBIdt0igWtqlumJZWkCIW3wysyPZYSl9cY9BlFH9DB
xT5asnQHo4jkcu1rsESQ8qYOiIAgfBZGflGV18dOYSPx1qZr6/KzssGBC7FVm0Xf
7zP/m79Q/W8JDcrODFL1p2fUoLvGe2eQAsB02tUQ00s++scB3sqUFcTsuXWSzBYg
SfU6ta6Y/U1e1rVaBUUTgG3na7rzcw1BxY9AB/4zBo2P7wr/1ZtuCUgHtkpyvKdb
JcgBzjczKWxYLUt5NcEmZCp0blZIhKT7pnyRDlfKO1n18nvX/3eK/7pLxPeBZz22
SVqcb3bYfsgbgkWG0+3/ynMMqKcwLJx90y8SkmBLPl5TbyVTCy+KhKUF9H9aCAjU
aCsDnslMn0d9AGCLrxfuzHwd0W07yDLS/H2P4G7CCo7bKdrs71yhVUG6rNUCCvLI
x2FIJz/JbVK6lf8DY0zqptiboHy14y5VdKJirvzxBdU0KN6Ux5TDDRrrtJfl09HR
+cpFrvChCif5//5h9tX8FQ4ofpyXQiXtPauNFg7UY/BTO6otn/xhey4NW0IHd0O5
bhg4hN3L3ewNWnUxAtxyg3mxDv2xj+IHl6UUwQJpqvYTyCR75ki5bxzojyLz8VhN
ANUJ/9ALqktBftiTPdxeaVMTxKT+jh/YUtWBBZh0lJnnGbPTWtgNwuzGNrgdOLvJ
m2d9yzjLpotLHWaMQrDtT9EmwFq+9+N+rJ7cLKrLlxAt14I1ifcF92jGxOJauoKU
E7RtnGs6y3U8KlAm33/uIyahiCdVodYzEA3dECDCFrWf4HwK299YFw10NtOexzoD
313JDxNRiXeLXSUVFnWdiCUuhCZBIbhM+Dnt305P0hSKxPe15bsvD3MUWWtohfWP
30HpfldYv9WFxDCnskMWcE4Vt7KVXsjGzEg5wmOJmXku4fUSG42CKd4A5HW5UlS/
2TIDxAB0GoYtsx5OBQiLflPjA38tPKiEj0rPA6DA+oXH7JQt5jMxpBpgk+hgPihB
GsD8jYZ/RoG+ab+08VXanhZEjkWmX5Jk0iXtN/6Refkr4JZCcUGTtyIjO00eugXG
jKX7KT1NryZpRQ0RPsTugxhvObDFes5cnvJpCAAnx5PwVTHaFjIH6kv0bXCnNuDV
Sj4rLkHxjsYjUfdtE1CRwBtl2clFvOfDR1bJxC2Cu1yUEgAnm3cmkoz0ZLluW00X
TK7TK2E1Pken3O7AU9KiI1eyCMyW4NLAIPDUzls+e5eTp8YqMizi6xxkENUcQQuL
xCS1frSgEaM2dtKARnWK8d8J+eAeH4zSi/KC4WOh5EjluIYbADsks155aKYMFiLk
GG8HvQCCKOgv64CqcvqLkXjPrusN7GvCPiW7zudun9PJ1YEkgsJ9VBXEyk8mBYff
mCPZTa84GpdS6BX8a2/DVSJXgfBDNCE7c8eB1NYQa+sF9crgyZw39cJF5M93haai
zce9RyuCQZECC2Lxm+zZDADBS4U3EoCmz7OLuyY97A9dsHji5O8odR90rynrLj6S
1I40C2VJWjVAUc0gR2oNfwuup0d4OeZjEZxnOVQ1igN4AfI1Wop6muZICL4YwkhT
CannIKGHUz8bzHhTcR/hX69HmO9nZUc3yTKZW567Yhkap6YobgdqYs0AXDHiZqOk
25uOeIARrkvMhpi7+2JrSffhMT/9XMA+HIa+6yUWf+IW+eIZ5MaRF9cB5g/XtJO0
Xow64Krxj9IUBKt+UuR33Zfem9gtmsgcwrYsfx0EsysdPWPisZo8/g4FNcycMVgk
Sn0I/1sKPqTFW96I7OF3+IE28hkX09yZX9U7DzZu9rooHMjbwjgsRbTZCsxuaLFz
mH106vVTGsSKdBO5b03sL7bt/p2SSYf+9OWCk/FV0cPchFngnEKUc2jYXUxbTc9l
XS2x5RcBlYLHXpC8ZS3P/GHAGSPAJxZEkr8+CuvMolTCMzwk41hbxH2cD5tn6Pp+
rnTVD76oNOSujoCQvT+kUEqH2DGWHT8RuGdQuHV5W1emnYTwN76ptvaQN24FaS2N
BMnfUiGrczMJEL5PcJ9nk1voAo7dhxjtSgznyfnHRyqkQLAHAc42n4qenDiJTwqw
i3QGlNpScjXrfh4fuJzauAEvwZhuYOZ2sEzgfNzlyq1k7Oe9PGwN1sK3L3yH17Pl
+L8oSGg85UUpTr3LAh0RwOGD10hJRDK02vHtZiPdRnPZiWH3oBuDLuSEi56Q/3b+
XNpMaRz+TZJ8lJkZndADgnXPoYQjfsqcKMwiILdM+49RzuBhMRaTlpu/LWPrwZb4
zXM4KtmIE+i7kEyMZeJxKiLwCsx6KE2ONCdZ+tS0fgNby9lYS/9hJ2U7KVMDq79d
YhY4cv2bgzjYVr1I7AWDLCdBKVpKb1qCqCw2rYMI/eZXkJNQnqjc0PhG7Il0nWRz
uBhPvQmwBhzZ2pdKW5FcuKuerRBqgKLtq9uNNHfQtzeq+9VZz8pFCXhme38IoW+D
XlRgKMs9bLQ2Numuvdqvi2n7/Irlg+Ji7bJn7WodkW0hgTPj8StFoPYNaBK5LzxP
Nu8RNRP24q6qISL0VqL2XLCsQJUTgGJhrlZTWVUc3mqO5ik7Y5iu0zB9MQ88pq9n
sMikKlNJis8ub8pU4n0iAOoDN3o/BLk6WuhFare2fQPFtQdAtFXiBN+UWpO//2SR
Oqcm/nboB4Z5kxqgDal+4te/MI7hGVnztR95I9bKZ1g8ldsltN71eDJrrhD5HG9W
QhwI8YGSItLpwwKEGmBOT3cGo8s+RzppVSz3Y48obsvQhLm6mC3KCA1TzRJpsQYK
pQEfWTB6X6F8/F5EAa/wQ3E2gMyDdNWNstMwJwlcieC0fHyAYsLHyacc3mke20Cd
HZw+WVVHPBwW9yCRopD/0R5uSfc2XDssdVq+JKPHtmyv9kJd9hJKFClU1qhcM4bm
kiD0tjFCUOuOen8T1NcY0Xf8tRmmMtjZTjp6dlAWMRuIKP5Q+n9e4x839GLqXJyh
OrVoKWgr4t9g0NHWsYLaZCH3rgajs+TWRpRiatNGhMi+l6omiYfwNLODgHnq0/Fs
r29bo6pGfaOWn3yE9XZq5oq03ZsgAG8skFtkJWnKD4Qqi+3xWRNpXoqiXuGBHCP7
8aiKQl0N6qDcpy0l7/2kT/keqo3oHIcWjLbmM37Vaw7BYPMu2rxL8pH1e7nVquQV
+cuY2OUC+I/lyfg4I1MOIfzJJ3BVzeFv8Jt823i666VDcnR9lyczYafmfDEuj6VH
Aeu2SQgOwckLaZeL1McT//VyCMIuTOKRAvlasBgZfedPi3zVDEqK6jue3doRu1cA
nYSeVJxKX6yAUB6adS9jhamS9kRzEeombaiGe8FJu+3vHvdM0zAOAfeaxHbQTbHC
JUguQzBMd0Skk5DyXt8CqGr+3F77DbHkTETnhYccoGXjHQHzOJ0Vur9DTC0sJjDX
mWtmwXlAwNAFwp4om2pXglF5oBiqP0i5zybhwxTxYkR6ryvYfdqDgz9mTgyXn/pE
/OKggvbrFqtBkc5ag0C0eP+qKs8cANoPLFrwh58bSVUax3dFmVl4oFMtP7wDqUmT
T4sZ2n6RnFZkNNVRzwkGeFDlkvUItV7EHrMvueXCV+h04phkVjJIE+8IHjO2vJbz
XcivpffLYyUAxL5zOBW5MO/T2iQcAejamFTEC0QHB1vFv7G+b0muDu8KC/HhtQHV
CuL7Uu858Vyru8IZ5d6SYlG9Wz8UnxzJNjRy8FF5zYFIOS21C+G7+d1j7jOW61Fp
F+E3qOBmM0rtTlvcz92+yQkri5cZREq5w4HXLcFHuDISa8BNbfNswgo8cuEavdxF
YpZLaCPOFbLCM/VMbgzGQYhsMsUIzgmpl+PvTh+2ulIXWQfKZRA9g7nvm83sIv37
eOuB+Hc4xJuxkU4+VV9FjJrsXgh5cNFkF0LhtJusOWDQZ6hlPjUU/yE1AoX4zzuv
zqBKljIpTTHlxyYMMaMV5VKNnuGyPFTK/O+DsW0RdExMtekHv7tnDu/f5ImhcLLL
GM076fEVxz6wUrXiZFB6wtC7n01a3BM2qHnMiFVdjfC6QGvPqC9W8Ruqo9UzthmV
S/eQtS02Rr+WT0Q7on4H6t6QK+JhxLp5+b+Cph1JVgB2zZFtAFjMgW/a7KhzBIOX
APn8y8ozIb59fjzGhux5RxaguIE16J24Zi+qAOpdf3NJ4xPcKbau62AKZBjE3Fdl
NzJWDvv51Lop9I+PAGIXjaT9ItqYZsC5KbU06CNzcijsEjh8PcgZQVJqrPO3DsBS
EoJHtH6geOfFUMszCpP1lxhyzYQ7bJBXhMff0mMklesuX1uvSeWvgNwxv9iww+iV
yVqn+kj8c1VjS0UhaCoQ+PV11tRr9AiLdJLVwtZpZBMQKua0D+i48oLYTj2SCQ5Q
RgiwozznrLfO1ObUszoNbhMzq6aLTjDB07lI6v2wduDhbQj+QKw09xmu/aZUUGf6
MHIN8tspImb+IH0p2nIz+TUS97zdJzi2RQkXrSizTb/vlgOe9WhOF1DskjPwIO2w
SLfYTB3vK5Q3vOopogKiv7OhKzutGUCh9ivOE98xtcdb37AzymOwAOW5snUX1Tty
t1VJgFGItM9jB4lxPwRf5BxamHZS7N1zuVq0Qk/+K+1M5/6GejyuGh8JZnw3YtOc
Qj7myi2qKDn3C/0T/Y5ElB70ttLVwT5rFNWoUSCjSsPoQ2oo0n9PJaeKaIunid4S
cFxP0GkEBAWh+4hp8Y2RPyavbZZXR61dlavLZ2QgWG3p76qAIs9ieRNxaysIchOW
40YqjRE9JbXLXz3WabeJewtLWksd0NClKd8OQgSA0MM1ypVZ5YC6g6vYPMNepe3T
Rtdw6xmf4Vfqg1AsS5JkjC5uh7bAkz66yswvIULG9lE0tTlz/pGmf/VgsM2EhSt0
z3hTINfcLTYflB9RFuNMPG3HE0Y02iCxsvJHF/sSDHNoub+PrXpvCLGhIoYON2X8
eGGtBTVAjG+VG3tDFe/SV107Se+16uxOa+oSFTc4rOs392i95Tivv/eF+U0q5K+6
U3/SvTpFL2B1EYtjz0dnJ2/fngOn0cY9iSZlnS7c09k8Dk5KvXI1wzRUFU9ZMN25
fzfr0fVoz2Djt96l3Tuij+3VJKxLM1sBltXesESIy0QOp7sx2FAt83pztSGaP0Bn
ktKoeIQZbFy37vkdxvyE+OY7e6oQLDGR8AIgvoW0p4bCoUafRx1ixRWX1h14Pjjw
elZYX2bKLeVLuQVXiMM36MGejmLPtdU7mOYZHo/JETEVAob7CaydJm828rysiooO
rUY6ubDVUtsgC/r3EO6JglNM8SoBiO627prkg+mY1Xoh2h7CM+apgLK5dJi12kCp
xgYKLEDYdHw2RChs4dz1Wr89ubI8auInc6YV6M7QS+0GPEibTag+05+ZxpKPr7qC
bA9r/F1ghQL9ZrcmRVvVyowjZH5ZJHMEBCr2ILuJZ8RUTv1qpRHV9A3dUPiPxqpB
J3Cl51VBWtkZmKyWC4bNUp0RY7MyW3RtvllVQQY9soPusV/x2DQr4bz7SzUy/Xu2
JmVqA0PuZq10AS8nWJJEKyfqMsV692X7CN9TwIv/ruPwBBDuPiuqGEZ2rfR9M5Z5
0jh/tcXFd79zaZLJJnB7JuO9lD23LrvvqxGdyBEqP77rbn6JpooOt6sbOwCJrtLl
gECx04qo/rqGCAIA7qTQxQQXwVTjhwv4MKd5fk13EtFZpOFPm/4Um1g/fP4RkRHX
99+SBs4/lmz5Thd4wOWMcyBCXPKgIbZFOWKTUPLEV0gg3txbznTh/Utky4fwwZdY
N+MSXI3IFK94AJNRdjVLyVZ06sSEUKaen0RvDoTn3WD5yGQNyPHcHfM0pNX/GrgZ
ztzqNkCcMoxwcJzYe2qfSnMQC7zaEP1bEK+YLhAif/SkMNmOT1UQnD+JZuTzyUHu
Wmc2pcnXSHvLTxYfFeUATMU4po2O/4PbLqU/3BIKUzKXxmmon/SmRNs+DAIIMx1A
drea4q7JHDi8FxRQOTOVEDWvfvgN69c1FV0GlMPVPYcczbjll1KV49NXVo7859DY
fVdDjULivJHM0PPdO1TGBIKXH75W8qXCAl8GiJWUciSmXWMbqyKl1yXGx6OdyyfS
pNfHnuQGZZdFNpX5Ot0yWrAyPaoRdquzBHpDALBUAQnKPa3hT8ceOQSod11kQbdg
coWm9Luon97Z9H3KScmIexnyChtT85RGDfzyFse/HCyDOmdz39vqaPJYdcx5z6My
utIsfdcd5zZvD7cVZLpxVbUfu6y5OxHhAoM0b2mG8X4oEFaSaO/saDMcd7o235Oc
c4qREhLeTYYuepDH5PidKaznNkVgNJbYUZRXdeOycV+sdpiDyEAS2YYKgTdPE6Cy
Ir9ixadPhtRWr/389TWF1pcPeMbbMhZJRGyrYDOrF9YDW8hCh+azx/uBgWOuol5j
RSrOkkfRW79C1FKfXgk72j9OJfy8n6g8fBoD4r6GL/cG0I+fDkUks2PLnXBaWTZB
0YBx3eTAmCWUd2aB97yKlbazXq4u4ywbLli5OpVQsf9UFi4gQeQdf6eIk82JCoP+
PuNsuGSSDI56BY9RLbVHWnfKosT9m6sTmkrSgJCz3JMF2vPvYH8ina342BrJpkFE
X/pP+bbiSzLkNKguybr8Nd8GVsj9iXSK72gJGd5At4ZGHhJwYSl630WeZlI8aT5j
fFr/a1w93Y8a2X+6cUBN08/JOQHRk1i3GeEymhAmL5Tgp19sv2zqn7JsRclFjiX0
ERZSTJwcfS89K7E7/qgEGq/221omb44+MxJa3marna9ouuomkDPQU06Ix4Dh1jnj
Re9jL4g+c09tinbRl8JgxBkXhey+7XtJrUIUSBN3TeBPrVUma+LC4X9w8aK3QkqR
1fcoM79WtHS3/O8w6LsovYluI9g91uZMlA8XxXoJoLico7C+YMug3ff4SLUh4jdy
6CE/B7uW7VTk6/CKMXa1pqvEM8UP/7Z+gy9xWJltxDNyszhhRdmEAvNUNDvIrtZP
tysm6TmqHc9zni4Yhe0/nfHT30g2sk6et+86PHh6JIRiJ2N8gARaYSz9CAVpKN1E
3hEBWQQlCO2KZR6FXdQzomsCbc5MxQZZV+S+g0MkHv0yBYi6FJJoh8K8bhpzhHkV
tJu4xCdFt8+UkO3aex/7iUPXN/pme/95kHuqoNiXqhxo5Xu2OrYX8PUpCCVOl5gI
aKjgC1HERxwTq8ivy27T7gvxAAyZaxYdX7fyiC+I3dE33woxsauHMizsnwLQvhan
nWflI8XdnOIIgBjTL3uKYoI7NsdnQD7Eld8Ir3oydsrTeqIkRkmoMoxOdgjuClwr
o/FEjgIQ9QKx8a5E/SQmyWhShMuJOMnxg2j+gGy+Bdf63amBf2BHE1xClwoqD/dO
FlPHHBizH8Kk9cQFvQ93HESAjvhW9puUVkIKaNoTB/5UNYl7kIbNiTZ+3/S6gTDa
DVwo45zj3LIBprib0xOHkWkU998VeP2EWoNSwkmZ/KD4AAQma1Yxq/dMhcINHThf
I4kIm6FhrXv38qme8O4YDch6wvWxjigvthS+7t48H31Y383jgtGYR4Fd2+ChxFLC
E+Usrra6nD+/9mDuROJWhIKvjtMevonVOsD59Rpn7AJj+IvtPR+jl9cQSCE+H4JM
kc1nx91fTNoxKjVZthafkzB5aFRyHghBtdVcf1KLiDvyDtGytXHlDfPwjUGBwz3J
LmUBbYnBPDDsB+uc7KbsxSjO5GXw8b2vdKeMpQqoUJPml3OEjMDV3rmDXQTNC5mm
VVEvAXVWYVsIj/R7/afLOOg00ERPx/wtztOgTYCcFSgyMfx7j8kcVz0h1i7F4XzS
6Y+RryiifxjMZs/m4rNNpJi5VdCqFubHEGqv8gg0pvZf2dsOV7ithOlsLBlg6iUn
PVBrtXC8JMyg9UyBJxsOC29n+S9aREWfAOjU3Xy8/xy/WO4LYw/BoNLMcq6N13Vg
iD8lv0Vszw2bc66AgsGsIH8s8UEVz3ec1KBAY8VvWBTGMHdwKaHVVD9ndIipyXI3
YFpJUUzJRnR438OFggAH0NnLiaXKs27rhMX9d6DxlguX/PBAXO2O7RWEV69DFPKr
i0zTYOWCxJQG6Frw91e8grPnGIDq/13CpUpA7bepURXwj61VVrk3bZUBtFuY7KzT
kVKpZuFmmUNoo4qdUGIDofZybCCnwKdtFRgRfaUqMvoqkbzXYlJE4bimZB7F294G
1caCWjLPqmiWFK8swT/3ZoChG41eLOHPZZUlB/60QW1t+sM/3VzbZrp62Dgzt/hi
A1T1bs6Mx7+k/PSprtr96KSbcweSBUpd51/9NF3OQhx+9nhNHxc9PDRU/HhfPXnN
hTgITcBDzpXiD1V7XewXhiXABySUe4ox4RAk7RWoPFU0YJEsSQvEMgYGSScRBg3O
9mzZW95uqQQXsmDt+CuGOInogpoWD2eTmqCQag4L9Wx8nBb6NQctaZFwXSU0YPjq
nwsFAiuQ2YX5ZfcgMdCVMW4GXdPOffkA/wjF1CnEjrtkPfoU6W4ApzN0Kiqq72r2
UT0vZ3+B2gFAOgCXfRelgApVyjASy1SRkMJbCPq8tfyNxfepvmWfzO6AAmdy1Kbr
Mt1A2uCDWN+oKN3MlqiXwIgrPti2W/OAtsXiWBHvKchNo0WpgE/4nsYC4QoPMaYq
mJG+7dRF66ScvTREmWx6beVHxSHBy5NBsjsdSd2ovSWzrQOWr1QiBN+q9hbm/CZx
oYrbQjIpuc8qANezSgLNHNaYmL/tBB6u3efthEslwx096BeotKqWGnv5jC7/WCA4
49HKjOmPM/Bhy9bHwEJDAALXU/DVTeHAeVc21VfgCthv2nFhgRDGfjoBDDxksnVO
L2X1gK7kUqgMhkerxfWTC263ZUCDrRnH6KLuIvJYhbVsmonJzMCRh6/XmxQEca9h
CuvWlnoUg769tuqdtugLc5D1ec5lz1jPPt5nHZlZPryMWRdgqqf6+y+rH4LVBLIa
7khn7POwnOIyq0GDMQ3yC6hmmilfGYQZO3mp+v2AY5VdDDmZ6oAMACV9QZhB3bpu
gtqqITFSn6HBcwmaIxu13NmmxcnmhO+zoXNvsXZZQZDeFgf3RXS51jztflRMsDCT
OAoYbglTh94LD2dXqxB1/f0ZpZxjmIcJJPbqCBuL4XGUHgALhc09BA6/sfCKjM9C
k0DXI5LiETSOgVgJVGzfKyNP3NlRYjDJfj+o6wLONpBOxGbeiIoAvbZH5Ztil3Jf
1nK3ia2lLhV2M2BpIXcNDImsVywP2J/uuDylT7cRg8NEqW8q58zif0uVGkTJeCq4
fAPBQR56QIfU2OQ1fCSzBzms+/XWRWPRQmZS/jqp7fz7CfuS+BYlnbgozQ0OSX9l
WYUSkaXRTa5M3agOGsNGu69LsQFU3BHhGHymRvU/ChpexpSAJbSeQgyBFPBUaDgt
IQVxyWVlEoYBsY7hsPFTilGa641k6suQ9ZTClgUMK58B3i1WTTyisNk/dxB3bUmf
jivTACc1rqmMdT0ng7ZWBAYfXzqcIYmfs3+6N8a/Nhn260LLdCMwwppk2t8GGs4B
6ByhNI3jV6iYaaK1gTJ85dzQpwyUQTEq4Ftlr8ELVCeFoUSO/JMQPvS6Tht/Mup2
44gQJZ5QHLdofLpNrB+bLQQdXfeC33CVDwHjZcOfqUBegYPO8pZz9nCnMRsSHw4P
hv4ayWXQwW+JNCvbMMZAQzKkpX4GjdwUjjQukrahJsL8HMT44LJGWWiCysYViPqO
c1t8O0q596jvve+2uJM6vBTek0btD0GZY3hEWbQt9njVxA+u2GnucuLKdrUOtF2m
xAElyyAiZXKjxEPmNjtTEJV5kC34ntdSqKwtj14G6c6s9J7hroj+bBlugWsC/dEe
gAHn19DqYuLF/KKcwGBj3/P79UmQHUfSrGA8hfuww6++U3snZ/hnlnxlT3Q9VJm/
+2bVTXMFah/6aYhijzOUBJ8dqBPu6raWgZk9Ge7qBI9hKn72Gff+CLGCOq4WlH1M
pC+wIELLK6cpr71+hj0MlkH5ZMypP7pFEw/TOM9tVHLitim2XQeDsuMLy8jrbCNk
ZKW3swHcJvX+VL7LQmDhn02kzWAYjl77MeXmehYd+8LutrpC7OQz3KYsKs3pSObx
Owa3OKgmBoieqn+X/PV/iBu17ynQNlsgjhRAIdZbq4p6Q9OZn5lICPKyiF6dKf1c
bOKUVmI8nh1yCfGQDaLwl1k2QqG1bAgfSFVJFIR1PdMPI57HkRnKYix+ZgZG+85F
X2rWRtgc6uEzi4Ke8o3+dpz8Lebz0lMBjtRyO8FdGer1pxPuu8CLjz1VpueRoX1p
IpOXQHkseKfyZkMN4GrxdB/Sp6kGlLrvF4kmdrvd0PZQleD4Tu5OQTBeOUNdG7NN
f8tNiu3qrWzr52QcOTM+KFrpOJGAIJ0XceVCkFKkOJTkFjg14EGC87pibKeS1xbR
8nRt7Ubd+bbTYvMWmWlcPwv9soKQHAxy00/i/MlKSJIDft8Mshi7zwCPz62IKAo4
/K6pS5BUqQQlosHhcKUDxMx/VZrahLH404fnqpoSZ6pKT4JpDFRboeieYTeHyyoL
TgoaRheX38qrS6exGpzKS/MMg2t9oULpJ1o97MoQlpTvxI738e3wCGmLhJi1nfCw
+X/dYWnodJF/dPOKrcoyWdEHFHvuUdnkqDXiwAF7tkR7/NyhlgqzV22NUcJI4mfX
L09tzsxXu2oRZlMpJ8LiZ4SIfLMzFPuLSltX8bUiYvFn8/bx8Y3DfLHCW1BLntxj
pT4NzJu5AlIRh9jyQDwa1L5w+3Bf17LompQv0cArC1Suux1OMWQsHUB0fdijRtSQ
ZLJ0O9omJUEKHNUnMDBdKJBOZBT3Q+EW2mh4qbqCADBZXww9E9k4roWMvmO8rcHb
L3baqTNYisEzHMgdxAHmEzjBtc8rPaFq37M57KJSCIFvBQFDFR6qaaOl8rEWzjfa
AOE39mFUAEOqtJYK/ptTvQ6ddpwqcPvOxiH+hWLjbs9NMRZmteOcFkby4/1e43pK
aQRQEptMtwbV8R7ktOjE/lEThUoVRid4eYgVoJvjOf41W0z5qPmy/ESpkd30cZ/s
nfjbJvLWa5MIaf00yx0bLZDf7rYxlPgfyaB4IP/9SJ9lDWoalLjc8Cmz4ArmyTp0
CIwgPzZVpXPO3VtNGyxaSGNtGMJXktLrD/Al6agl5sAzNHhYHmHXPQDt8B4lUWtA
sN//RvZiuAuov+K0XmpgD5gpPHluGUcRtqXst5c/i5gIo5puTe1yWSp1Kv4wc/NX
qATlSvW2ZbINZO+Qm0UrRaoXMstVqIHy0AuF455O6W0stySs063B8ROJLEES8CSS
+moSmAJ2rsPBFxgeT4Vb+a5xiX1vB1t1q2PaVC2Kj0GfRpxcfTQYP+Wnpf+tGKDq
i9BIkKgXujg40TTdODQI6Pb0Gjv5PTU0MSheQdrVwKBjROCyFTBuPlgxHBhSG2Oq
0zOmajV09VIAL6IzRBtOJn0FHcQi0O/M6CcBsa8vplpjv6n+pkghOLAYdXME47nj
rdLbODQy42k1JLpKZr2FcPN9pobpV0dv7wiM/Dec2sF64O5OP6sSdNtRWskTrIGR
5rS5PR+ngRj75JBjpR3TK7dHQoecIBNnP3FsmRjkTzkZMkSaunfuXluZbLpfLplB
bRCzZR9gsgllLQdia6h4H4lrYE7XIpFzbOdTEqSPoZF8d9u2bJ0R7iMsZPLsm2aD
h+tyhUvSJa1Fsv8MPDOyAsFp2knaqJOBXoPeFjbcksoWs4ao0k/XLR6/BNBeLRbp
xoIXUjv5aZG5Vh8G39VsUXYjN+4sa1kJfBAfghV0g+FTYAhXkq6Ciq2qugZQGq94
klubzMz9+nKc6xwhtIoLv2Zx5lQ7cIJHpH2pG+4f+RWLuvzDQHdK4Ht4U3Cu+HYF
OcglnCVuVNJC1k6Pxr1uDe14XJARZAw5mpEBWu3xPcE4TVUsaIOQj+D7/tPI0v8U
XEXkQIzQPIR9snPJ5orY20TgRgZI10pHO9vZUCAOQDyFqJEVplsPs+j8g0mUxgUx
21ST9R+/buGr59JDgqL4u5nTsZWysVIzB/+jXUV79jL/FZccuPq38sV01O/dp2vx
n/i2Tjsgeco5t02ZvmdJM/BK6ed8qy37gz6qfp+amfraWeZ2cOD7X+rpI/dZWmge
WrdPDUOkbKYWtR2o2Fn4ljkOr8sLOiSPj3aT3Tol2hM+mocdJspoFVDT3KLP6842
0mun4kbQ/D69j4Wxx947iOVIy06VFCQLffJpZ3EpAhOOYLoF3ui+gvxp1SzqfJOj
tj6VdTzyIimC6uJU1c+zaFDsQUcqHV5SxjjqoFwhhFJ3eyyXDr2OGOwz1/P/0ykd
hC5z7ZUUD7cddEheoUUhxj7jiyMwfFfm9/iJ3WfnosoSoh5D1npC43qCPL/jXoic
1oo6cSFDk8Nd0tzkUPr9XAAqm507nEUxBnhTOp/ut9Yp+8RzZHBv0YGgZP4ZgP5d
rOhBvqn9tQARHbWYdBYucn3fFnAEP0iDsTk7+bkv+dnpBzK8Gxf8LOTF2Ec/Q7DS
FK3eo66SyY2Raeyc1NU5WU8r+BGayfFwmni1kJz4PemtbONX/oSh2zPAY8esc2kL
szL9h63VLGOqfYv79WdC7ZeLon+cnCguZ9ySyduBymxjs8GiYcYin0SBMSyzuEky
5HYbRSKbKTR70IAxfsIKErEsG7jHFbcQAs/3l/DLN75OlaUUV0enqZJme2UnuWTB
NiDL//61XS9T7rWKXFGiECKHaB08g+hRl5Nu4fT1MX7u176qeoPmtouhIF1jPpxc
u9tG6OJq7wdQEv/DWLoiBmmz0VCK8YtJhObQs58rnne2bZWgEEg7T3LgibNBVu//
wRDATzCurPVKzJYjSWLF+k64vQJAJ2P5lY0Xd9hEtX5FB9/W9zsYeJAEUcUZ4Lgo
0av7fqDTwwjVurkSO849Rh607ug9htyhzfyBXBL4V6PNEOTOMxZyU5fCgMlVTnLa
VOTvbPXJm1Z05pPazRlKVvioQ9w6Rh40w7ZerbmOT5BHiQcgdSRtYVcGpbOVtfo2
yZyLS19E0wU1Fnw3qIbSMtGPArAT7AGPuN4TeA2g1z83AJO2ZFKg15KJDxw2U3FA
pzFE+ct4iwjuo4vpNiXnzmyMKBxz3C2JmNw80uu+HkmWa2AdkWMMXATzn2Krtx2U
vYHzHBFn1OYSHZiGBvIsrgSDpEOAzE0raepUeLi+YBmPOfmYe1RCvEN9VUAHo2x/
dBjjQZbjwhRZLNOu1MjEkcCH19zFCuqEi1MHEVPQKF6y9xKo3vxYqA3kAxDNQD5H
dPVT/nn5qtXE8sIx1uyFYAy5HqDT/H0RTvsqOo5PoLqQUwb6InXhkAXXereBOx46
eH6qIIx5mUdwh8YkSHM0/0mX91oM0FsWq4biQEsS22Wv5xyQWNPJklhZqe8Ixp8c
141ErBLWsFaK9Ls5SDhfWJZQoJl47CJq5vI+w5FsQWc1paFp7EwW087rNg6a/kTp
rzcP+Y5TVeEVgSGR5cx9dMGhSAwlQw8v2nC1T6sgje+wwYV7rK+kbTQL/yTXE5id
8Oidx6n36FmANhsHFwY2fVfxz2gnk1Pim3WAsFp3Re/Q3RU4NbBK7tYeRX5JPCQw
Ax9CdNZneqaDxVny9OWGOt6VrVm5pWcfylNEULLuQKGBQE8e3LXNsF1XHlaS2gvw
qSkenkRlRDrPEP+oUEF/MkjZ+n6EIaDB2hFBVgnYseka+Vtapi3UL4ManDjwDiVg
d0/XG98U4EQ80TQiXvEhs/905AcyZNlel9VJijTahOHmPIYJkXZvearC+OtDpDHd
LsSEFRAE+D2jwtBXXWgPUTkZMDQFodQw/Vr2iSoF2MnPftIpXw+/cAWYVGKGhizu
Bva/6tdtU8Rt2mMiX6icpj1yyYB1u6LEM94KXpsY3E/z3fv4NRSVr+dPQT0/p0Oe
RdRDb4cGHjeQXdqIOTU2oaI71uV5Mu3/H6wtpOG3OQE6wheE3iOn05KIg7xIc0J3
MInjHfR+CASQ5enYabEHXZQ0fSyJkRkXlTkx9N6WcQb4zeVTJzEH/YbW0m62RK6a
vRFMhuaKQAAkl3wEXNvPesQFlMtqi5Do4pKA7TNjinrezeeGgX8yV0I1Kj0UvAAW
0QZ3h1wW3Ts5VduajpKY2Pzjlw332hga/HoZnGwd3jDkCGpJ0izaRxPSpLImBOwS
Q7YgYWzzshTXpimmdnli7aweAOMNQx3FRXnSb2SwfdTBc+f0RqlVGHpSChq1du2B
xQ4OVhZ32GKSCl6dOy5MBI3iXbFv3sYqfsqn2t6nBjBFE2EC4piVldwVHggrmBaK
5hzSMb1gB53bFxKfole8l2sp3LnsO1Vdtoz6ODE4esPHwgIWI2wKABXj/36T1DgE
2ybuMGgDVe7KqMCTRYLTRDlWLGtc36cTe/571tXxZ4OX/gzlcHwz8HcsFiF5lTXu
VrYHHEv04aRt5ZyEup1PGOlJWEaexvIvWacP9UMu5P2LnzVN9VsXa7VZSv3/N6L0
EHXgi6ZdG24Vkpisb++EHYks1SlzjyFxu3Psu4AibAUAuTjqJXKroL8UYGwDeEq5
rfS3dEBsTXKzkVWP1QHrv14uEDLWhdkWDLTNkaGWHNsUlUegBCk5XTALq5Mei2W1
EZnU4my5iLBgBS03joUmlHFQWLXV9JoupYY8hy2gdNrS4IABoM40FWM74lq+fR8o
q9oFfzDv2hi5i8Q0kIw3tcr7UwzaeoCVKYw5zcTXaOmJVe5MEunnsoB3FvvbaSUg
hPjk+hVN6ic9roDaiRU97FOM7IFxVuWT5USB8YydWnOaJWBeJPgPJ4pO0HoEYcIG
ycrLjL3judq3yvTEiBzNMjziEucR55w9u0kbPNlzs/UXmX76XTbL1VPFjy4NtF4T
ZFy9RMFq+QC8YoC/vICcBJDI9SAuY5w0Gfak/vKCJTRe1xafvnk6um0JCVH9sDUc
CEAvoPiB2w2QFnFjnFZv3qvAJlo1d2VF2YwWA6JnuhuhzYgQ9C9tK4xuJExKQZt2
nFnpcHSwUz/Jhs1FQzdJpBaplMUmYRN0dafdzFyLQ+zd8GYC57wr4nCwULobI6Zw
/vpNlbr2UOyWQw9Ysvo9vTfNYC6sj8tuQmvlRIOWB7E7PoHtuy43k6+LFNS68/KF
nFZCsMxJV/NzkfgOmTQDW113N1QM484o0poYYHaE429e4JN8r0yAqxorKG8Ljh4Q
bRg2lAgPwOa16/bQNHQ540h2ByaiYELkUOlgOOk2KnKVc5F1QM6GLhdPFQnw6YFy
WiuVXvglXtQKLfp8Dr7FOG30RHEinYvQLoawND0blj9ETAZ/POCDuVm9HcD6IsGU
2PTXFMLzgkMfg9RmrdyJSiSoYNSIU7jDpWIdn5t6Ie9GXqrnYmBk+TwOtyT2T3op
A7t0FPSonLcT1O/dOE4KHjFs6fpyFdB4tySJiBDIPwLmZh3CI4mnfZWaZ+6PX09g
LvYIbjGjJr0nt22eJxDHT2KT3vgNJP2V2I9EJ65cteme3TtBm1GyHWdUus4Nkcd5
3S0a9vvKuB+nMNiF/ICjpLIdvRNrgXerWg48fcqSq5C6m7AZClgHeSmS8NDvtu7W
XQDmzSIPmA3jvIOUSFZKN3swNRGX2cDsyWXVqO7HwkGbkUNyKK4rlBmhcYG9IyG6
BkrEkNUUV0xXdTSD4dFpGbh6GA4BwqQ7e6G+NeWaingv4fWWM2HLjnsO2TI5Vikq
LvjK77KGaPxBXzMFq+i1YiKtXDRQ8+DmICV3tYYEpUukzKJr6XeoXQcSZhU/Ns9R
OvBoO3rp7Mji+XKnfqIwSQiF9ZOMC8bZJ4ZAmdaaVipR7RPxp09A1OeQB3wHWs6e
oIrEOiIg8Y6wGv01PCELpaZQ8gFfju/J2JW0eR8GtDOkMCrgH/G2K1bA9/8U7IsW
dkXFgpihsJ2qmoIPyUrpGAO9NyQBRAdByk3tQK1l93eM9fmlE6T+UaSaPYMsNT4o
+ew0Nr/4aRuWppNKFxLH822yDri47+h+nqX120ZEMwYmC53TA59IcVjOWrCeTpO3
aM7UttWE8MRtEVu/6Qp9trRvwVi3o0FOx0IGG0TS//LP5POj5J+fPgbLRC2lpjaf
D8sJtE49VjPRkOdSL6i9lYkHcyQq48PPX53Nj0SEQfz4fIe3pqk6j9IsLwOfY9+T
YpZ5fTCZQywVOScuBLDgFwzRFvthNrvacVoPOvQa0U2RnEROs4nJABET7amy5alU
Gy2/smXdBUUR8MyYGS6AJmNeQhQCvpQ7UXyxO+ouMEshKh4zt9VUkL8eDyyH1Aw6
mC/F/OLO+Nm2TYnVxz0k1LUpc5RmunxzYZVhUM1cP1HbF1xzaVUOVRIshkqBFAVz
csbRpbqqVfzkLoMNNPYuHN7tkskSjwhLL/E7pt5a+fgDBn/7/8cSTM7kW1wsf7pq
9B9xEcX2KNuJguUbWurDMsowU0aiZbvkJ3W5gyaUU8SvR9zsblLHvAuauY4rwLuj
l52QP9yl86vBGMEZhAMCW8EhCFkY/QbX4qFbeSnMUs0XpcJT6vt+nEt4FB6jkN6e
EyRPQbJflCC7MQaMT5gO3b8HySn42mz7IQROALK0jd04d6/tqzw3twotEK8NA+d1
kmJiYueEffPtY+uUdWKscm8WHUPq0y+SE+AsVGqy45KGuUF5/xF6wpDkDlLg59qE
9nPewjkD85g4amPvogN7OMl7cBIGiWXl49eqMh2+qPkIUoACcrL3qmbX/jnOVn3W
QH0ZF4+bVUCLo4MoBjB2EVn0H87l/aAmdl4TQY1Ho/JNkG36vCKnn3KAHTRXQwcG
2foycaDJfet+pX6mNF158JXBkGCovwYErfyjGMiiMP687TPW2gtTqo1C5CaJuc/e
U0vTDEPN6J1gnhH+7gavh4ArcGZOTocTcliFL9SQ6cLKPv2MGsl4jaJvXYZU6bDP
yg6ikEhCwzVRMfxNt+g3e94qQUauqu+LpmzApCkZscCGlCTbe0YzUzodyFtArfFb
b/FA6FU95hNVS2ZifG1KTcatDC31xo26n8ZOHZxHwH/WV4NXFmM++Us3XqfMExy6
sK2HmR+NdwXhCEN7xm8ILQil35bK9zFNQeu2Ob0N24dRTHmAwvulaxYXfXVfwtRQ
FnOIDGOfqR/nhsGmnvphnNt4lPw7ViHMiAuswnW6AjvNtOIlRRFUlKQ/LhLtawxG
sd2uTafdbS8g/pPdsXHgCAFADqt5zzqpiLeJB7HslwNvfW6u/ivyfz+KCtrSdIgM
1LTD4/hz3Ireg8l7r+LZ5GwvvluO1WvnmUfd0hRgPvI+9w3GMV0Rex0Y2Mum4RW/
GrwnMnO9sQnMa2x4sbk2RYrTgZ5cpjkUTIWHkgYKciOENBFZd+9bGn/b8zO5o1pM
Rj/K+sCZWcY3Ht/r1rGFj+J/KmrWi3LEnjkNSnuYJkUZG6aqMvI7ADNThNQMilvN
DZT1zOFANm9oLFNfEeD0pmrMUW7BHUpMKvOaHowIjrkx5Fgj6IMZ4K8ARhrQh6g6
FKC9JvI6c3ww/8hRyKo8Rqa19nWJy5dT5lSKYfsNxnU/UQbEhavk/kmBdmizIysq
nOsTxSkGPCAWv71qNgMqf0MYq3lHxWBsbT7AxeTFhbgQKTnJR1w9c8NjT1kNGaaB
pcYekaKcheeHIWcfM5d1mDxEBqIm8SwEwP5W4dTpeFIBf106qoC8lt1Wd4NCS+pC
3xQ33uTIiVEBgA3CwiBK7SmNlB8TgZSR/gw1nfwvCF86lsG0WpG5J5MGcDUoY/q1
du7Qx9biTLlI/00wdUA2QgwsBeJENrAv8gfJeeQRUeT0+eZ8v9o3cxUuQ36J7izT
RnPfh1nrD21QKZ2nCVlXXko282ADJYwjPRAbTmwknniLyvB9hXc1GYMrXlIR2rTZ
EFh1NhC3k7lJcSIFTtt1z791ovYMQ+E86Cqk+VwO7oqxfh8LKbjiv8oKo50k0H8x
Q0g6YoqT693yhfO4ZnfZUDHLOV4QYKrocoRvIfyb65Chez+u4M1zTNTjAaYn7S8E
DIWnOYGwj35LM0VY7dpavMPcnwMim64fY2YEJcpeKjY3R65p7rX/oqRw+msTzga1
UabosjtZapXvRJbFS9BFSaIraLHyUl5RMmKr/7QSUovBASWiLYWbN/QgDHv7UHIj
TgUnzC7oDeiLYZGMFdcTsrqOrwPdjsi1bqCxd5C69mJovFGGAHmzb4YkNtoYumnJ
GGGmDFA2TZVov5LUOVGBDPUjxt4HfTywhNvHOM9pVu7iPpTcoHCZ0aXFLoyM4mcR
yBXfI7dvImB2tRLsUIAg16P4l66V1P6fKBpr/j02GXsJ1Q4NIP6xmPDvbfGmpRcK
RnPSdA/X0Q44oQkrDmv4ISFHRc0v9Pqlcc2N8BvSSZ7DCyJRmN/pKEM1Acr2cUUO
WB+33DVhfMchZZKaPlpBaeFmaVlPafDlhE2SsMwSjA6dJHZynGWlueDEMiOt6Fa/
H6mwsnRBwYzXkw9SQrhDeMkwFg2eMxq0N5gKoIQgSf7chlTIBGw4DJ7plsyo/Ls3
cmTKCWA3yM/Q61pDLS+AyVhED4fI5gI82FY9Nl3DGS7mluvIT+g1Hxy2I8eZ0gGv
PUuPqcfasKiaWDOD/o5QaTkpxgmazblM8Sxts1Np0/UtPqUB8/U6DZyasYGncGzI
IFpvLdZnz1X9H2PypD+WfN0NdGX3moioSwYmIMMeYYfqbeO5QM/4c2cXz5digvux
Nn3GQZ81/tCpNoRw6PV1GNVlF+35TqNpwvrAcFfbDa5vEMfRT5JgWj2/DMdjUZi7
72+xs+bU/5XYr1X0shZqEpDsCglGvZRyKVMe+yyIxvqCnsfWny3HTwu8xVV1pOef
6gGu554owv/GENBPOkqMga9i44QvdtZJjDhGie/bemHP+3UoG9iXu/m7GIdojHep
6wRmiPkheTCAmBzrCRfmKxPtjGbyTAt2xmssack6AJvsUxwxTq6h7r8R9vQ0dscz
I7PXpLfhxPgyzxG/j4yrgr5/8JOjnvrnxMps2L4G7+kdEw7RxSToun6t6ZbmYJi3
9jAPYjX9qh58bzXMPQPCKpqqP2/e8pMofqaWKD901oBJ5fjgEPedbql7kf74PovK
Y3jgtzEo/SvoNZQZBIYefR90T6d+/9Nvow0CMxXl+EgdSdxtOB1ssr+SVPEmXTV0
wOxkF+/ODJHj2X+hN5AlAmh6R2F5nj3E+xcbdiKKIou7vV8kpK4KWrCcYV5hiPZ2
H6iMTuG9oPDfHjjYhh8WuucS1zmEFFZdfYwnfoAB/7guHr59nsckksYWEIvH/4n9
DSHbouqJae0zi3MuR4n5LZyRSTiBlWEf+Y5ondryLQpi58GXfKdAAtDmMQ8uHDDR
U8TeF8YmVuVQAGPGwVnIjb24OQmP/BdazDRym8zmPGgoX3etGlLCC0Uj8nirn0M3
8FglompQe3o/q1Qi54359yON9tU85bzW+18hHpzS5gPiwZ0JvbChemzTI1KkF1P+
xDJHBVxXzZ2DNSAZEYkww8ZtDG19/r3QIM/A50O05sI1AvzZeq4GfRDfpWG7V6FW
IaYXgrs7RKlI+rTdXC9EOcBLDYg6i7RE/koj4uA6nC5/LxRNIPGe7Aam59df8mW6
1XIGqIyO4nCepnsAKjLmeZltSZc+4cCzQ0t99iXz1qYjvFU7ih857WiYq/ye3Op1
lVpEGzNwxlSDqVPOtyRd+1lqL/JrKjbj9lsCNnZsllkJU9yz5/Z38V9sRKMxQ4CM
gePNQwpJBgdf4B42gz+yqy48g+Zu4uIzSSrMpwpi+eMJr9y5HWtAncpcSpVTHRKD
T48w0lUc6WwQc9wJVtPi8FVdR/0X4IlH8L7mKxWe4JoaLo4kJrDgxtFcVdB1qgMN
0fyA0XUeacOKhwqn84nOc58VZuVwct4dui57vGXev83hyl37vhjKkUeP2KvMDd2T
CjjhZUDwnhuppr9f4usIN37k7Twg6PN/bWnjmsRnq0/Nx2fOr+Jnl+Df2zMelOKR
pzddpQv96nX74YuLuHNTcKQ0jDPd5iYdDh1zN8agI4GKFIx7Z48dGMT5fsDEYBLD
Gl2pu8pOML0hpKWDelk/KXzupHggjm2Vh14vkzGtv0ijvYxxJQJxv0SzNRKPUt3X
adr9xE299K79nT/S/USpOzGHQQHCf7Z2O4uePhqpgI4enw/TrN8nAnzE0G9kgV/i
l1r5bOHhHwCyc5G3hZDVgXQucKISNkbEa/+PFrlJayZ/mVtNVaY8PryAAwj77f1H
RCXX6je+zP6qqVR9Zyf6M/HpMBZn/D2G+WIrSVOTtbOF4AXkN6NRCaxjRI+J0Uwl
d8JuPZRGRA+24/A1MH2iI9Wdj4SccNmdv1HxApgsVvRmMlH9tTY/t2UnSoj83bEV
pFikjk1E3YyzENlzV73SlCrlav7l30rJvvT7ryqFOtXIH0/gMu0WDcpyEIhvV1x2
OsEe3ooGlVgI/QTm/2AHNP60d6as9/xr4paTNvLQRz0hQnR4V7YcQvzfz9dKf/u0
RrzF3MP5XtSRo+9aeaszCRg+Y/76JhTEfNoGQu36VLaL6vuvSHVm2zn25IeoN6nr
P1ccQ/bowJ5G0Y3qNp8ar/GkuRnhnw1xRoFxF6xC3rH4M8uzMLGbchHChz6dePcW
i+Nh7MjLkeeABWPg69WhKIiqdG/B1fLgvjVn94Co7jRHVklTWt1fYG7U5QKC6Ylw
BI7803crgL+boIWf0HqPmHdGxFoy0zxuXEJhJX/wWKwuW4+D74BRKPwoza5k+xDZ
qnevLheWJtfRcvcF9TDdx3/Hu1MM7usEqCyFPgUh9D1W97Po1J/YbmzGRetE57Qw
bAcK7DB33GD7mP9rvyuYna0sM1JREOoWiyYMmbfrZkNDaWgbBzfuK7QHimP+VY6j
wpHIuRgeTzHjh08wZwIIoRwzASEzh52uIbLPvddIkAGSuAhoINJzulp0UC321JPR
tq3kkZmbhLXnAEv4/t2bStV0gSWFWNO/zhm2+O0KhTfzLgiuXpMSD8a2EHYjYDyc
BYOBhKK5XnFQbo+1g8qpiNUsAOYTR8hEwOWKtDQ7lysZwOcW923EAj7CNk3Yx4Kb
65Nh2T+ATVOYdBSboo2an/Eiu3Ja048MapqD/29HYMxPfRv7Ed+H/0O/YbakzXyz
4nwIwm0a+a2GDXVRtybIoufIdejd2oHBL5ejXzxDSM44MmdaWXqaPXMBxOvwxARr
AESfNaZm/8IJC8S8yfgBk5y2a965HqthsWHROJtxHJT2Xta3tV5qW3yP1+qk7GqA
CkKljb6BKchua0LAHtL4NqT226Zj9k7PvaLIzBkHUg/mXtXYD+JX158RnW6fzd2g
dGZLXBY5HVTBfg7pckCphA3QiLCilcSkYPJLCtCh/W9afIM383g97n6xacQrqPzy
9pGJx18eM6efQXaysDZHgD61ZAn+giRvtsncFEs7DIo6y07P+OSA13AXLYnxKpqT
ax+LeVCSckWMFy86bsCj/Z+0Wcd4sTReo5U0DkbHZSkYSQtIgHaIb3XgLIKfA/Od
1J8lRCMdCkoKuPgbL3ntjzL5ZS1F9qK43nb6gf63+f02g6Kf+36uPI8n/YZtYkIq
jTqaTkdnmEdMbMHNP0y3EDYEtZ1AeLbReWTqRL1kH5oYT2xCwS5o31o0BOfF7Hj+
DedfmR1bnSILYVBchqQmOgu4kN1yPbtmm7kGBRpl/onuYkzPgLb4+9XboKsOnraL
aGLoNRwVWbHl08A8wl5/8zJGRgIL7R6KuPa/v3XzDKPX6SHksyl30M4ickWzSgQb
ZknWCjRp7cx64pI+f8GMhvTBkv0cMWjqGgiXVGsKFjClUeoMxwNZ5unABgtb6In3
JxHpsQ/SAeXOwSePHl1ZMiqySRJZf1awFtDv+SrEA+rZe0jN8HWfZCA2SAoOhM/y
7Js+3v2gIzrktpwEY5LbU/LHA/n0i9PwZry2wSMAd6QoKyhOW6AgaDinJ1qztWDI
XfpTL9XggMF6rV/jzHsTI6XFKv25OFY9QA3XWv2iUnQ865TDGYIrICQKiKIGA8YD
ueuTomHAb9zbaLT7H1RW2DZrUdj2Zi/u4f8GE1bAhkS+rTRtbh4y9/X7UnydcC+I
vkuLS1cn4XROjD9WknPGRTr5RtaCn3JoLNdk/8se68t/j+MHtyfwxO678KpXQBsi
SgC0RXtaH4V/iAloUjPBm95qc3TK4BbKNnVbP7M5k0TP5SPh+KQrQEoBmKxyGVuZ
nkEqK8/STAwGtSdqEnmSsa8Sma7dTAt9n+w2C++44pradz88povznkmbQlk3B2aw
vZO4D1rrnqcDTklrF4U5OZRxLMG86tMGmeod4Ieex4nLAo4TpObYeqLAUtSGOAFH
ZV/dmEDvjdQlfaJJNWhj2hleAh8HZHnTOXOexgdCLr12qPFYeQYG0ZEVgGuOUyq/
58pTBtjniXO1tQ759VWnA4ECiaJ5xOld4sCCA09Q2NnVJIUOA2gZ8BRzDqYb1Ikb
bvlKW55pytxt46kYv8T5Ii9Xnx8QOSK0qKk0MtLJXYsh2wW9QthVkyV/5rkcv1zH
18eOej2AiPdEdlVw9W50Zs4SMrqRo9Y451qcDbpUu1fK0hGVFGm1rkM3WZV4v8Iu
3mAIWdtZtijzwfY82kAJisOhNSekgDMI0+9PTV/dwf1z4LdMYACPwgwtzxgBuDe5
32HRZs6+0iEn/LQV97ofsOFSeplW/xVIaoLrV+Ja76I675TnUo4qz5uCWZU9O4LD
zLTRNzABh1DTEWJ4tBGGSvh+/jGbRHgl81kL6u0+Fvrct9ldrsX+V8OxvqsJHjN/
zKKU0zfWhyrHNVEo8l8cSqgDTb1lEDlFsqPx1bWEKO/oQ1PVPNYdqkdsBM6bCZhE
ac4NPkINo4lCQRXWlpUTu5mmuBOXVf+xfNSieU+ALIwM23zgH9VMgFteiH9fM2NJ
x5rkDH83GjSpzXhyOGX1Ero7/jrf6Xkbz+0lo9E4VFaXCKskTncf+jH51eLCUAik
l0WYtYdTXR8RGntiIK/ZCeHgaCeDK9THzVt8mp5nPZrFOXRliu5q++mJAazaaRPN
oRbocMYmISxYflB8LNiyTeJm+XOYDOZYBm2xWD6IKivKRm41WTFn1L2pfNjoUS24
z2h/QaTVxtgggj/bdKgGA3KNphGsQqNW7gvdtpZNkWwJL3OXCzYJSL09Jk0ocg/x
AAG0RmmKZsi3TwUGbGsauhUzTJ6c2Wad8AGTL5bOZKvaWCk3K9K8rEeF/e5XMdU4
76+ILu5i1BGB+H8N4g7Y/dl6l95WFWvSo1maZAWCDOMjmkQmBAyjQz5KmJD9eMtx
MZ8PwdKWsy0rxCMIdGcIgefXj/KlROOxEOBn8uKGEaDBe1EoWJi28JV8yzZ4kayR
Pzqf/9CP3iIHRDmg1RwtVVkMRAoxWs64lgCVWOK38pC5Wfw1HVlsoWkd/R+k+1kX
SyqY6e6a7Y6kni0vX0GP7JUC6V6p5sPUS7i/3M0Of+F6ehXfumDdQKmVcIOeMZ3q
4/VzuLMvRwrbA20D3LUeK0NXGbwj3Zbi1ZGbI22XdrlI46VQLZLw0VJo8SMwCtAJ
qKErXdyN7sUZ7cutiq20N+far7cSXlZMOptV9rYCd/E72RAE8XlXFUrcb4KL0Wf9
+t/8ninVwfWBxbUxAnkxXQ1icGJReKRS8014x4rLbIaoy693ALtikv2SJGoXIdPZ
wJZlVkjrCMaEVXCrHhFGAhYRd8xt50UOK8O22z2fzfuLSv2GsZ4Wu88A3GnbOv7a
lmbflOTmrSY56Rc4eXXil612II9ur7MG5CHRxlREXk/bWhnkf+EHj7WqRnbgAJo1
mfOtb1SxQRLTvuXAdLkekmd02np1x4PJUV9RsFHA3rkpm0j8i7xHjQoHJNIbV5QJ
ffpnMg+rDqeRoyZMnvO/uqZE0mZWK0OiHx8cLV1xZOH0Oko7zzOhkpX6XOCh/SEs
Vk2Yu+v8/L8ErfifPXuCjs2quw3sGuiwRdWRuUOZpN0SrIkXJMvs+xZgHTJPCKLN
ZIMxrmXZBPSk3+O52QaR3BwYod6drt5DWJ+X9ly7F+qWGgcdXBawegdgcAPPOXtW
3l9fnCZL8dTugNPNG5sueqDArsJB7vGS0FVkgcCFGdW4PKxkQf3DWKhMY4jcx+Gi
8VpIIzOWMB3mjK6o9/XSCKaClCUFrvaKHitj3p9lzQk/96EOaQMcFMTmlJieqXWS
av8pB3TiSeh3/zGJBxHUqPZtL2g68iRX4r45IszEX26ukw4QLoPeIPY2HrqwAKVR
5ANLLrwCyvFsS4cuX2VGKhkxeB8Kb83Ah4rOWTlaxl5EmyiNbgFEX6YYEuADJ3ek
k0Vc/Mr7skA5hfpb+wsI2XNgrfTOpbPzliTz26x5NuJ93s5YDfPagAoGIqPlpkYp
2QG6Gl4kIx8zJUZRXFPReOkFeM49k/PYW+YfM4P9/Eck0N9wb2noPJkYiZxHXFER
qaHv0DyAMnfngbz1jOZFJK70Nb5Ym0J/MMXYUW3+e1qzDgppOT1mp/qVtSvLqCqn
9nnZrcbA8qNQLikQ9XcX21V5xzGpknWeJ6GGiINHDWoITyBWrz0hQPZvNT1ddDlx
b1tgO9caHbKfrDqpvrB+dCGEDbwYUxMEM5Wx3vdd5ZV9qNX3408AOJK/VcVN7pO9
EcjyCDDnLNl9TB/sbQVfFwBHJa9WGV3kLZ9R0sgzyewiQcdNcvVdPdCcY4th7vMU
8/rzzOavSMCjaZXOuFBXae1xqUPrcjkntFr3vsQ8548mks2YYjXOaYpLnvE6UKO4
7HVQO98TDZUDQxbmzYgwiKePeYl1pcjXAzzPdLp8J2MHCjCgxzFa0jbCudb0/Xdf
sBJ1ar8rFq8rldn2ZetraO5I+WcSFH23rIzC/zpCKfvXIIYte95xlekY9vzHzHHv
5NO5EQCaAlIGj5FHlDgNWDRhr3c6PgfVpHkDn5aODmZcnzzucvupa9HMrMP6HBSb
BnLck2VDBqk+3vTAXOKnM9LOi+7WPeVIAlymmKywbvi4jwERtCqGs6GAFpILCw21
c6JGtEAxuupkfrLfLRB+/pnpc6Q44jzyE2PoHi+QU4u98f9X0uIcJuq4ElmoHek9
mH8nMnwBBEipqpbyo7ogzhCp4HN+sAuWR/HQhEAFLmA/VAbw/XxHP5+fPJnF1APg
kyjuDLwznnAxCmDzjtQ8P1ksp3Xa6rx2kXa1hLqXb/hyX+LS67h0jbslp0/Xdbp0
S/3FDyqvSD1o1+LCxqiW0LMC1nsTFoJ6CgmA/TniVmf7b/Imwm+s1UO4mCT6znUj
qH+FCBfypTcQAz4Cu6ujQ6zN2GE3gDAba/kFkunAuoOlV1B9vgxoCyU2DhCZYiga
zs+28U5CxFzNtMFFJtxFBOc5V3Lp3SeVGSNfY8s6RQSl6YEwQMaAa9FIq6SFrb69
9tugWJ++k0oSk4SaPtF2571SkTQWTjo9hIV3P3tqvcctxfd2rf9w3tCCoXQWaWQw
DiILA4HJK+BXCBkGUSOXtcK5bktVr7Ls5xmmclfgHoZNtLtpXN/YV4IK+UbJsKHg
HGRRIxDAiirlxKzxHV2zJA2qPyQWHO/1pWBesJNye0pGcqve98lhPvwHYjETOutM
7gadKOrTBT3q8CgOsx9aqRiY/pLcrJQ4Jc4i63kRM0iyJrK3V7MnVnVN8KoGVGA9
prEl61OVUCWmjDnjjCCpkslt6UuEFhWyv2tOKSMR1s3nOdFv2e+HibBefaB/jFbh
G6Wmmi4Ale+RLW7t7jLSahn+Os4ls5TSTzMZXIUrSWVUkXpKcKjw9r96xOLFkgQD
ar+1VfcyhHKk8rQuFvXjZBxLuEBf4xd7uCnFbBBsYvka6T6psQIvjm9QEMiWVfCR
8Qno/sDLHTOrZF1/EBgD3RqjuSpn8R2WW/4RnkLvcT5HvAEcsUv/IwxEgZf9FDVL
2+MQUQdj7sXeDAUFEGXh0Lws8aB7VslHySn7Ygsqn55CdUnzrTqZrHBaa3AvxuTB
lXl/ClyUCCM0oFPNTcxFJ8KH0kOrnDuSor3UGqlzMvySUcBqeljBLvqOrHU7ixXb
u6Ivw3MVBAopqpmjXcdZk9WWDGdL8uzljtD92xGKX+5jP+EdM72LX/q1hQ/WMMkO
shXRu4JRj2WjE9yxws6FilsXTFmZslBkzWKlnBOxsJhWcRUgcACztazc537PUuWX
37vMe5fW4Fu1lHITqUTK/IlVKKiJVWcDAZKCe/+ZgSj9oakFs6c6ng0AAsn76CSo
ADI6j4O2Gfb70nV/3n2x+By6DaLukr98GNrZdHrNtwyO/YdvcYvLhe9vplKYYOtf
mcFPbbsyfTtFWM0NMWAruIwO+242cpfz2dbdpDuqzdMZSXedjsh+W6EvvKEy/fP5
eeg02jofTYgUtmgTF8GCFZ3zMC1ws5mAEYg0PFiwgfVfI6op0fO2FmyAfBQxDxzI
kGQcfW4zFXj7mJpK4f4K/lcPzz7NwE47L14v9njv0TUhf8ila4owGc+zyBo0I089
SLwSVLKFeHWAv4EHL8iT8I+4UYVdA1jgaHjAlMo+rZH0Il6GvNykVSxVt2y2f34l
P9gx/yqih8FQmWcuUl8VV1QgpYxv3cI1e3pLcOkVQDGoJPSoymRABmiVbrkMM59d
5k7NfcQTEyYV1obqAJp7ASVzrdjizCDqftaGnh23+sGpxkTlxrtvJoEg+ll1eEQt
FEVmkPbYWpSaJCRvhb/izWgh34+zBe0U/SPhpotyIHyoZFtwslPbhMZS5nkCLB7n
gzsi856tW8twdKDW5Si+dbKVX1jofv30KF8utA+FXV0cOYgQ32Syq9kpuDuV2gLm
fy2PNdS/xP6uBufnmJBnrsvt1PU6wjh2fCn3MpI/lcyHFgTZtD/oHpuAao75wnyd
FGN6M/Xb4BDmfNZ+cQAsHE1CNZ2YkmE3tPwv09EF6MLUcEH4lZ0KFS965zJoXJjv
hFVpqMGV9HQkr13+xZz9u0Fa6i0ZComUWVns3XkL4jDATjX8Dcb748nN61lxrgxh
dceKMr7LsSq5LLDIjb80kh8xhSMfOQF680a48dDREwU1goMGMXWWuZWpc7CJaI4w
RiFQaXn0vHhgn9NMrysBprRSaToQjWSjkADcbu25timPgShgZ+nUCb6cFVpmZIfG
c/zx5nr5r+1+bt/43SsLlHIDgL7NrWHPbBoJiZIhi0qsHeqUuVXVejF7JKdkSo42
imkcamJN7hpcjpKuZLUnAjGJ+91I32jrFOAeJ5gEBNojyWJUy6Vd54YruZXSmQXD
VRtEcwTAeLrE3VUPQmBQ2o0x2HXpQAk8rY+7puIY/aA9Jc+yW4JT55xm1CTIUnAx
j07JRaHO0JfSs8c6/yNNuPLLPtJ7hKOu69sScF2f4eYE+ZkzH2wngjIZuiyqCab2
a+H6mfTILmEDLZCzvSmPs3xxmr3NvUy7BF4/hXQGbBNIjoQMxjaID5S6tQ9AScJA
nFm387g+xyPuP9x5/zIhhuMk0LWKI9JTBSbVyoyaIUEaeW/LW6/uGekfpONw3W5D
fNreIC1hN9JiiJt1OUj0z4EN+RRPT+t7mAzWRlq7CZrcUzlI8Co4rfTBlJ4G6WEp
IPqQ5kKnOBSXitu8mRJswZPZc8kVAB3wzBUCokeAkJT2S8AEEVm1hI5UdeWYE0Kq
itxK+bO/sEImw+yKPjk6ZAXa7pSePdGX0MZOElCsKmJB+kHNPXovS51EjQkzdxex
cnkCpSo6XpXUYoDyuPzxCH7RnfaOAJmtJQbNbWe1tzHXqsIypCZg0ygL9jkS+rEk
nSqqcTLuvcZtwsJtCQ+A6N4ZVPoCjWMc6ERqzft+uKL/3FKF9QDFVex7h5qsgzV1
JyGyjDT3NgtdNejgpUgOHSBml/Oy0I3ulw7CSInuuD8RED1aLZt3Hy0SqpFKwMH/
WQE4ojV+Xlbn8dWd1DJsrHl8tEEUNTp9//CfVsSsR7h8kvMaFqueiDDEEGJuBDJr
q6imZ61C5Kd39xBEfblgsUAOl5WCueMOAFaLiCtnZjmvS/IUkXmB+kXOTPQNrtin
AuhK/kRybgMZUWfzP/wZTLtyfEAlGMNIw9p0Vgt+ATQBCnb67BcljndrDBDPsV8q
Vc+NegTvS6LjYbeo4a0LyGMeifPqqr1qWf8KI/zCCJtKmOct/Yx/74G6lGrKZXU8
+WKyiJ4Aose74xrvN3nhJPuR8cFNdlrslgkXhrQK8h49DcWtmbzFgwyp4t0Whnmh
Po03hGD2raK7SpZdHyg3guxD6zpax8cGeaNdZm0D/zF7UDYLK56ip81+9o5Wy8Jj
bGurr/57CJnUvVhLInNZvD1Xrp5zFwYZh2bruOQa+Nr4Cg/Bf5ASGXrxJndRFZPL
1Vk9YJk6u02MM52QkH0VHnAKSBYHh1hD1jmP7E3ocdM8LUwqVC5/P6l3QXzlUbXv
vCiKiZEMt3V1Xj46maSILI843O2eWMhhaGa5hN8OARg0FJ3+cEbPRd0ygKv6aKnZ
avKT3JolvysulpfSVFvcoELMhFkgZX+UhgXi6+2/2/ueXG3fvJxab7/zh01ch1C6
sh4J9xmgoMuPqTEvSvsIpH0XdSZkOcO5D/pYhU+xqcVnRWsCCrcrk6jGxyUr1A/4
ynv8AaWPKVQugoqqRI24roxRfzAqx8VXSdd8JbRKmc0/vyAbNFhCsdR9XrmuD8KO
yFXqv4uhjTopg2eY74s9zG+dJGWiYN8A1xy3grhesI833b1GxTXSfU8rE7p1aiqg
DIfKEHjunK5K/wLP5as8VwmVHA7Lmd8p+yQSqJSmoHhh9dTtMc/2VvwGzFShQIqF
HIGKrpbVrOvGIg/drab5AEX60ZfcFiRuRbM1MkEMz+M9NXr9HSh9DJlMNAizxAlR
0FS+Nr2CbwMQmF4tsc8X9KZ24jHhX8UZAFM7bBDpj1xOb7KiPve7zSqkk6P9hyo4
Tt+5qrneUcOaPpBlbPhJkoy7lCdfXA1W93hd7RxNLMuXubqx1M8a5mOzKF/7oqH/
uagZDDVGSYpI8NyV6BVL4DNXv5vSDnnEe8TtslT8qhoNJx3uyz3dYnDv+AEXh/DO
j1IuSlsDkiTdFXCxG6phHEkvXQibBBJ49LdhFXH1xE6KbrNGXSIyhzI6KtsTSybr
+PF0UOL0HjPeRl/d6P1qqDIt0ggmK9ihIPcobviKkpH8KjCe5od+ZbbPp3Fpu9q/
kqJUov9cIUA8BptFm/oSL+bCdlDGY3mEP2HsXrn/YRItsXOiPR3KZFlqIIIDDI/5
TcQBv31y1FQ2Kn9EA5TaviZ+cICUuRuD4JZCTsXPbE6KiH67f8TcahLevb+BcvLI
GVxT2Lajoe+7cIP7BNxIp0e91/rjnurn2mO98FPTB5uR11Wn05KmV/otn25R5K5g
i1PG71cTSyp7hSvWQO5EkPj6MTKJP+KkfDFChUwBC5XoVW2Epfp0yzwJud+cdM6n
E5qNknkdkWu0aX9CfpqI1F/BNPJo4c0TjklI/nb5s/jv69tM69Zi19Imhc2nrFmm
0DmUcBrXY+YjilkB/e8TloyrZCPUphJQgap1RqD/a+ssg/qbr7em+ZP1P/Vr/LyX
gEST+0y0QHZRBMhnxQb44Te2kPD8oMiv2WU1hKMwEAC6MLMFoOZaz9IHd2ERXSaC
mKp0As+ooU3xzccldylVjCb59dp1OD6CGuTznBVQSYcTBeLhVtcsWNY4TT2rgzfu
KxXRFM07LuWJkQqxNJc+7M8BycJlDzF7QstF8fNK2Hxoiy/173Lz5zJTYTE2Zf90
YM/45LLCmtj0YmSrMvec/4cyLadhzIQk9SXiDW56tgIf3Nk8xfhqZzIkcaR1T2Py
M+ntZHN3SbaUa0WvUQi51Zb93JQ31WbCLsv19nvqmm8Gd2wbWfTOy1FOcbb+FkS2
JNqgDOB3bKfLCYe/zvPWxEHz+v2TOslzKvwsoizgg886DiglvHUhhMuklZJeYpfn
Hk/0VOR2w+kQhFmNvNQdcsVrs3NZC1ssmyvko2Z0sSSk8tZG+2+6vHBODavfGX41
D61HV3+90zbQCd6sKWaNafgr3NhKwQl6vC0qbZlyrG0CevRnubpqlfnbt0wuSCsq
8T7xEhOxm0E+ntMjT2izJw1WjV2yqt72l6u1AzvfPcm0ViKuEfWHlzxI2DDui37W
A/wm3f3G3plszP6UGMM03EsdM3HbZ2CnG91FDKZ6e8pSbAf3jFoeibnU2SERzqcI
Ztl4QGW0B2DoTiQxBnduxeOSXmU5PGvi6fXY6OpMXqfzg+FhZ3Foy5HOZWX4zQ6i
G7tMJ8rBXV0n3BoJqGKmgJGFYHPp6i4Tp9frZhViiZoVeq212LxMsgdV3C2+RHeo
mHB+9QZ0t1un+Q1DvqFo0flMIa9VGKyJN6o/GBPLkrcJ1dS4LTO7qbwC3Z5OSg7I
+rrXA7v3EFfMH+dSI1o+kUWnAEH4MCO3OTT6PWZVOPSgzNJWCW/WYfb+YMwILXVQ
WCQNEF61Sunu7fhtbkd2qsINQxKddNaPtJLY4uAhr4W6OFfcQp4HC5r1Xu9owKJC
FG/haRq850RBSTMNYUUBEpqyMvJsBu0RYxcEHaImU8jQWYH9jaNUoc5emgcKoNw1
5PZORV3CaoxabDrhNzaloY00H5wA+izHLFZ2BhE47nOVOLlsu+xYb7jtJuu7Y6Jf
2jMSkE1Cyc2PxOsubm9W/65p0vPNOpcISnDTZDa0ioLTOzHTahhzQxMDdPxpMYhq
AxPcKbX2/dmJh1rg0a3sCxBSR8pEJB2iZIKQDj6Zd2dPjCVA3j9/GnqNaLPchAGj
JJt8qExSE3oZjJJZkbg2+ce5rwGToxh2i83j39AY2xoI0PaNwG941p6Wat7cDncA
mes3POYBZLLfX2dzS1CTr5djWMQtt+gdd1iAsJrUKBFYwXLqpHyjUQSt+Xh1VpTO
wEA6zQueLBHsQNcGYpiqb+Yb7jwift2qsm2vTgTnIPjv3eUMwNSGzSjQr85XzO6C
TSk9tfY2gX8OzLhPW29HO8PiARDkYbvIlBnf1K6GIISLxHt0IrURwUwuICwUnSf9
6IA0hwdyQWzg91tkMWdl2tFJyBhXh3iQvg/+Cg1bzLvZ01iA0o66krwkRNglahW0
/b6L4LcZntoYBua9l4CRJuDfDWJyxwWejFQu9u7jFjfyMD9cMKLYSkVjuq2E1n2p
TtEiLv1CLAKrheqI/MhqfpC73n+cXYUK6K/BpEbOtu15F1nxtNHipB4gCex5LDpn
x9sfBJGiWBiXWLiWTARUOikkgBSapUxk47TCg2CG4NnkszD1J55CF5TLkUKMJuAJ
71lTMaZj9PpQu3mf4drbPs/Wm1Khic1+N1nYS9lWDHBaUAEYljxl0tadWYxEdPhN
dxBSN9pKR+UPGg1ZOKc7ef0xtMcrHHNXtOWJo39V2tpG83le5t9Ycfol1+AylkP4
P6w2SqB8+m2TnkWElJy9on7q5CvLdi3/wx8Xd/pH6wT11TYY2C7TahUNwKfouK2p
lpuBYsBH6dwsv4j52VzX/Y2/TpGDWOnFTC0CKG7nqA29xBddwKErva/A/cI+gkyA
LOMpalp7pWiD6+v4C38GaNTn9ls6UT4RAgVSOtwutniIXMmcDMD/Jc/8bkpSsH++
m/6hvnIeCCKuz4HmnVOUgycjiyutuElX/YETUNtJXKQLm5ZJlCEN/RV7PVYh1p6i
k+4axaNqJJe/UODY2JgG6XYcjJANNNdKvppT9ice/aYwAvKDQjzHxs9iL/w/PMf/
nDmYKWyid9dMmW2t2mOBBGhrbr8wYslkZXygm7xHGjQ4Wz35jc0vHpWuB9uSV751
ImXCH/JiSoRik020+EKkQdd01AcgS2IidviFCyjZjg5JP9TFz6mJ/d1uvkYWgGFI
pTQ+gdGDd2ml7QzMtH6N1SjfbPi6AIUUj6jnt1NETVhhZ3kovrVfUTeRPnJwg1QY
Yt8Sz41NUJnQApXC8CufPRPB+t2lyX0/MjuHxGnB3HZ7UcOguWJASj3usKodqPhO
aWqLyCsbDTmVGrqB4fiAAu47Pm9Qk575kmXqW31t+YVwnikmZg6tmBrTXJSEdLnH
xEFVJn/5+F1FmeH4DnBVIvPmfCpTUsqsKuy3/ZxVLaXw40m6rcvEw2EiZqmQqNh0
KUkJWcGyNDfwahp2lOE/NCL2EdL+ZB3ABVoewlquTBHBvoyy0OmGjcvqiNnQHPlg
fR9fC5v4KYSowxqFoMX0sF+lbjwsPF4gaxW0Rtc8VqDnz+eDH7tEgr0uB4Ekxj9I
uBEn/+gAfgNl0mP6rPbW78zvohoMLjYTgHzIPF1s8jEFNQwTQnD2UpZFoQkr/is5
EI3OM0cuEQy7Z/fAh8au+4zMMMwAiAilhrzesLtoGF/mok5qy6pZ3Qh3pIa/J5sQ
+zkBYzqTFjg69YBDbeqDq3xtczHG1yTvD+dyfok80nCo1bA+xYYxt6Oly5FbMXqM
qoBQ3uSJK4ZCPNDsdZmeoIvU74AWDF5N7V9/R95NunEs7n0NcpezUuAEnHdT7Ehz
xS0FYCohxUAQywKIXtx9W0fRx3U1WOM0+Nq+Vu435WXG0V4GMUeGomZ7aXQZdvmf
Ctco1EjtPrq6xqFrdQZehFreJkPQDVXtcoSyJptkdjFojU5U1DT4SoRVAkV/Qf86
ikluPcKX7Ys/Cba0kGI2ZOwbZ2X6SlkuIxt+eoCu6hU//llfv/8IPixEv6vPHPRi
iWBUNNG1r7OKhJldt3UBzt3zuPSA/0R3XQ6rqlVZQk7qNszbar5Xi/BIItM7tljt
Aa4EaOZyQLD4rY1USJA7LefVga2UUKosDXDMTswVFd7Zlu3jn2fo4+JS1SaaqM/9
QTH1n4FpuuKBAVfz2nAf7t03YAn0WOrpOl3KvXr9TRA9pPkHyLp9PzWcI3DvJQza
YJq6ZXXkaBZ/8OQ2ZkuIdcK9dwdsJ6BNmsCppgCXCTfVIWhc8olohdVgptmb8ojd
5n8sfEQd/baukqx29kNZOZC1svuqcIWzkS82WtQPEBvnrE/Ct0q3a1OSLh8nkqis
l2wQ7TIMiDrL/2bGd/kM2iSJXIVXP7QA/MlbMv2L9AfUpDVBTky6q/yOJ19NS1Gv
FMDaGW4uprXAPuN7Y4Y4tr30l/z9bn3hzgEAK/YM9WKybN/MZvOa6ylzxwal4/0x
hj1YPN6wcEHnCIoZSNjHS05xnnAppTvHHr2q5h4vm6j6m034Ef9zrFPLseGT++ni
yzjFJpvLdK/56YeOpu42NAsdw8wBfEqmDg4Qof/GKNp1SnTYDgQOTkWjl/YIeL6u
+OHhx7FKiFSiJfXxVhDXtjiIeE3xWjkzuYBgFKCTnqpFKckdIhC3EcIvj5LScGp9
U5/g7kYRu2+srUShSFhNpl+vm1MIyx+cSNs1W6NWDX9x/9x5POK86AgQKzvYvtdL
avmOMf1xBSH0sYG6Ct7ogACWrMviVPC7MG9P8Hyuu9f2TlldYomUUWSN9Yf2eHUR
S6PXWLXBSDRXUZvwUdvGiLVRYP2qnkzN/t3NQOuw+qkuwbiz6PcmBfiCm9xxj5K+
GSsOjBJw+6Z0PuzwnDj1pGQJ6ugbKkl+cXX4gITBfRPNOUiSTEEykk/cD5R2jyqz
+5UzmI40AaUxHQrV7pADYUOel+pBmPGT1+u5zJusXIp/SxF3YsUbV0GRAr/GzasD
9Y1hsRY37XUyIMoJuBXIXZDIdQ8Omcez+QJtAgphpQ8XnaI+r46rsfHkZhJzX2bM
6bFU1gQkqM2T8DsQfsFHtpLuDYpjwoKryqnwdmcvK09eDl+IqhEKA6IuWDK4Z4iN
Fv1S0pfeG+0czvPgXLzCraclgGWuqX6mfMcU1UoZVFmWS/l3LNP5DLZOuB10hwXw
Rd14NgNBIeDHTJ2v2vwMbB12QzHZrfQM1aalYt0j9xgaz7Kf1iUKe2RJ7Ec0BZjr
2KK1Sf5rkBiR9S5vV9N0KIMh6U91YIl5tAUNQ7KVQ8PpTcMMJkiPyWMLprYzSLSx
JzaQcgwfbkIpbehjeXtsqMnbAwsWvWNPVgj4KEPlK8MArDX2Q/jLiRp2jE2IlePx
DfiLgMA23EhdO0Bt0HNr1aBYjVhwCQKy5f1GUol7M9sNgjC1iz7neSywycWLQ9tO
4gXDMxMFj0lmP7aBdqUYzmQuLTTI1BFA95P0SHjqoK+/eQtiHXFyeTkGEnlQjv73
1TDzEmS9SRkU4cBL3XIFSQCD8b/3ZICdXPunNYmEPA1zMVRFbE3Vz8WTJnr4gP3/
mKiRgkyc3lCVGKWWcWZsVJmQs2YyMKZ6kPE3jjP4vNmQFJRMO+9+0dv19eRebQl8
SkYyDneP5g6fT67c69Bt7yDLjlTlWsVEo7YbccHtLcfYMjv0yHFZVraJ8WrJTECb
40bbLg6X8L/xyHP1+NEuFRoejfrazNGT3kjAiGe27S6IHczJUbWwJxCAR9Ot1Rv0
nMxBxMqJ4Z8lxBCzL+eRPlaveu2elhsVl1cQe41oCDMzUtP9N2yyiM0CCbz42eIK
1+IG0WCDncgmF/+Kp4JeIYsw77jEJRGREvxj0PD1a/1qXhWnpLlKgjbfW1VE8sVd
0J62qw55jDBkhiv1ib8cM4V1Ymm4KHRbyHfstSUq3njVwp14aRLet7G9GYEucwC8
iJfN8iWSJYKNZrFh8ciaHTbf2aAIpKjrFyPbv4HL61gwpY6e639fU8FJfij42ciE
Oz+3CNv+UqeHfKoYFoivJIX6alc4pIDep76k94CgUJT3bYMAj+Dl1EJpBon0Wih/
0kS6UxKr2m0Uh/vIWK3rlXoHDnCqJkDwwjJ63tU+joZ/S+dG5Q+8VJDMfxrnxJGl
0l4THay5v4NllcOlv99YUJhKCNpgLplva/3NOorEfGa65yeAJfikyJ0dxeelqmCp
rNo2stU3LjvIvxrYSGfrquWX7AScwrggB04mh1xCrimJNijFdGtzh2316G9avlpD
KChT2ZDJWZF6YsLzhsNRVg2mqRF0z7rzdhPOpSsnVkkCfQcKKIRgd3Dp0WFIzE5y
4Nmu179xebtAimtKaVRJgd+98EGsDPbU0fDvaOu028YsceLIT13lrPDj0Bui3Y0F
LZiK0LR+FNba6IwhBvDlveyFMpo9ih6fpClWXBxFQ6p9SR3Sxn+ypKTvA8pA83r8
fw/0R6vBYo4mO1aD4D2CC+cc/BByBwA1nTJdp26WXeyz6B+Oj0E7FvDxoRkQcRbZ
HAcHOgP3tMu1gF0bV+pBstgnksMiO+cUVse3y7vdc21LNe+ZuaBSdolUz5ZAwqKA
yggLidVC9e3nlK5sOp8ae3QukrlebZBrLlx2/hzopldXsYnPv7WI0qofQK5Ze/k5
Okt5V9OgiOd3b/CbEdWcq/qexkf/ygfQ/FCEFbVXnlN/JyXXcxH4JbCIgeQHSxqf
zyBAVuLNDlWURVNRhHo2+xXglV3WrjB/nHHrhHdao+sG/WwQZDXVtnLmM+dwBgA6
iiZPFde7ZlP4EN2S7uDy2XXRwi5blsjRxh0yDQCqbmgh1gcxQwLHTuZttxlc/LY6
4wTsLfYvHcN3iv+G9KtgLOuE48EqldiNVjLyhxX7MR8GymJAE6oFjMvmIb10LgTL
fIgMFSxKW6Lju0Lujatp/uBwrbCeow7BF3pcXP7Tppnz+aH/N947fSHAeMysKC/4
17UTQ+WzGzZPmWI9ZfLrHDu6paytW/05IPdJkuCprTGPgTrkpMIpCrPmUQdmnECc
KkObM0SPLhPL+zIgHUXrMtHeJpRB/5rpSyEQWYhk89vXo8p+yr/+3L0O/fzn+twj
38X9MGwrlQ8rkY6HojL0oGw2zu3AjepWgQ6SMvKJ/RGfJy1ZVN6onpHzYMXK2mDJ
al4lX1CmEJhbQOJ7dSMc31X7jZI77d2kr06OkjplDOrYZC6a2MHfjWru1DXD6VSG
LBh5UWSMeXkWFaQk65fPQKQwBGlJNO6f9guSIvXFa6n+Vyg8kGdX9wH/sMW7Pxvc
PAPTXs/cNZnQySW/kiDipyeET6PM/TFzLANOfqeVXpVROrFnGw5cAw1XCTSQwXWB
pvVLgsfM0a9UkVUEk5We4db0/fobyp+HK1E3m3aKSu2q5PhZCmlCmBXdsphTPe/0
BvMO9lDCpHZWVt1mgIAioplEWS4U4bzMbKk459p1OLTC1CVGG5jtg1MOuriwNlVX
HPOlf4CaunW+3k/DwIzCAt/HybH1j/ivxkTvbahRGOzpWh5SAlU0Q+JPmMWMRxCW
/mT4+/isFtsDuWPrz85c4mZ1Fz6mchqW0korpzxF9DahTeXWgZsTIhcoRgVCE7cC
qONeHNslDsFquWi8FCS3CvXmkVqI8kK2nisOxzOfcXth3FBMFWKsOkVJ9MX+Ql9T
k3HNEZbkglb6rOWmfUH+vUKT6yTmW8gl1UERt3SRYmaudHLABwKlwmaEccHfOkpi
kJw6z99GB/zby0x0mqM6l80reZVwozwSiAGydIF4qh+Vmw96otch3A+qa9Zc3558
yDkwQICDpzV1fsvfEXsErc2OeOQXPpCpNQixF5zRj8TWpu0GooYtvcKFw9Z0JZ0B
lcjLkpUu2quAZ6jwRnCekgkEBmYIFfRsE+04QagR90Ae3Xxtj0FZqRtBHY1tpE0r
X1JvLfGh37p55/Sk48CO/u944EjZCuyyNbS8t5SP5zFIImURLc2doKKJUM6mWaf+
NAizOPPgaPdx+LjWAgnXQ8jz6O946Q29kFq6whicOJn69nEV6SbfWNKzx99kqEjR
dXo+Y5JGs8ogAN45HVn2aF8m8SdLu5E+ua5+K7cfP8ZUpNucOtal8IcT8zgU81H0
PWVFMkm26FUU94lmzSgc1doIyI2CfDpLp8WZhBvuIT2kj39UgadF/iiYtp0lf7HX
SwIaajsJmG0pNEajJGpOEAKQJbGkPFihVqR9jMYMUSxQomp1MXQM4Nn8//S1eoeZ
3rVQKspw8r+EmuLO5GhW4zGAkx4oEbjJ7tOLagV8KJkTjRw9E1bQt3qpkhYK4tH/
vLhaWogHWOlXSNlWR0exY+1KJHRHltmn7o55I5G8o1ONB4zeMbGlo/wfZbO/ApiQ
6J+FipItb5pa0qOwPPKmkzQQw1icYHbyFFK4YrmKsVT8fzm/g17HAPDOpUThDogw
kY7P3YpttjXoQGyRw1TaV0DleiTuZpKUlIUNFg6HgWAtpRgRWr5UqJMoi0VG+wnQ
mgv8TYph7pGJdld5gYt2sl2f/Xw20/nE8R/2KwBP+fAbeRqa8QWrp8WPRJtTb5iJ
paAtNmBfWT4dZnACw2WjqzCyLNQ1aFrundsDO/WseAfLTUi3gCXo5/D4q7nMK1fx
ZZ9yBvLK5fj44+LL0Hg/0HpBW/AKUHM8e165BOGFBe36K03obYcRhAJULdCAnUPL
x2j9QW8bAlow6ZCdcd0ZgwdjMX98rj6CPYk374855klGwOc2lnSdkqKXPujkGphX
2JTh94R52G+GgOq7NqJrGG0DRZelorfNsPl9/LGrmSman2VeSXil0SBsMDJREtzk
1Q0mnd/F6hNx7YfKeoBZrQZulZPsimFsotrMq0Hqa+frUEp7Y/HaaP3IiE9/QsVQ
+nzDtcZ05rEaiI/sb6MlSfOUhkKLU9IHOYtLoo3RpMdWG98CI8wcrGpGzB+efsCJ
LnIUUFZW/KS/2400m6qKOlOXAzm2hY4KAb8NQ9J330KGW94EbxHv/2KZGm0qXi40
s5x9cMRhxL0UOlFYCIBcGDyVjnTQ2nCJKO3hW1izilgwNEmVQ4AuodAE530fQ0lj
EnwLCnn791rE5834GIthvM16SeV+qIj9H37ishP01+Fxt/Sa+EOMfOHFVVgKnD0G
h6+bWMQNFNDVs2ZtAbPnL9gXMK4+9m2wlegLaR5A0LQooLAYUK8OShFJiU5AQjL/
tfJYVTqxuzKEUyYRJAHb1+P32Ue3ILYmc9whmUwaOcW/4X60WVCVio4DcoIEU+JW
Slooeb6QEARheyeXWVJJZXppaKONgTzbGVq/cdgmWmuXaE1D5Pe2k6iRSd4H4NM8
xygPGUGvlvUCxQydpuWVYvvDdiCp5SWNjyyTuZKE5kl7Qx8+tIQy4hmYEmBL+4gS
PO0aI5YlAqyh8Gzsr11Et3hj4w5p0mQdvSUcKCTsLj4K/Cjw3gSQWLTbSRdlDqzr
9/VPLphykz8IqmzqyTN62iOWYY9u3ViSvRcv6i09GpoLHVRxCiLCc0TH5ZQbgarJ
ltIUAFjOUP8crClIcBjeXM5Czo08wvFIeUw+xaoWBaxjm8QBd5u3Ipz0QDmk6J8A
AerRAUN79pXMQUjZssxQA+zEWsb8uqVLRFcFuCawd6kLY8RTnSMZd12lM4IeP5VL
X3ZlZ2ne4BLGW3m4h045Jkq4Cd+LcV5hcEB3w2mDFKPQEnc0v3fRH7yY9ZpflpWu
jmF0bH9sTMSZf9s1AfbD9vszW1ynfyKJ2q7AqzhOM7oQ54dnv4WGiDXn9FHiEhTz
o4jwWaj3L1yK9P3ledJ6tZ17KphAAoKQcnyWVe93+EHed+RONjW8t+cIrkGId6rP
U0/mM7WgJx04LgTCwkGb4LTDvlzfivU4///p1osvUu1A7W9Opd8+W9OIW2+auDVy
kE+oUam2Nu6354Bnn8ZApVhB236e0+BZGSM1uG5HPfwIA4N9Ott2/XrH5/e7XzDy
9cgvDbqciTkyJs/2OPjhQ1INp5pGMHj8NBdbjfY2D6lniCudKcX3sL8iSxf2z0s8
dTkM1aKKfjiTO8SiWFUT/9RGmwkuU4DuWvSHe9N8iu64ps7eBOpseuFP2taZdgoZ
U15PV86LmD9g/KcOUD5cz0cLgPeGUjkHu3B1fW9DUbHrUCF8/1miEZkRS/DbAG8E
coMkMnqFD7Mw2xPoPmwfNPFud5R2c26FtJ4U44BYr3WlAEiUKoYpAZ72mbqF0QbK
VBAKHnryjENXoAg1EevxYpYBma6+QCKAKVGza/pttPC+eey/2hHbGdzXyAh0IhdA
1juuAXsw0QPEOtA8+UeVhkK341aHkYtVzSH9JdrLKuAEIL3H16jyFL73g31M87iy
GAsuSOKkPEOcSLLIkfOa6vKxaFx8mdFFY5KbmSqXT5kL7Sau90sMvOI1/0ITZrg2
0+ZCR/eqLj58xQsCi7vL8yl7coyD29Y/5qqa9PhCu5s3x3oJq1XDLO0chech3xNa
DkGLhK/CjQDf4j65DKNjEv7r3JUhF4etWwE9udgtW0tX3sJOiCjhoTa5igbG/mHd
vkRlEMuhtp+fpNNKqNuhTDyPV61zBiUZnYoSBNuHE2cKxbW9G+u8OG46EP9Swj3p
7IB1qzdQlOHLqNqxmvTGIntTTPFvfcUkDdg8ChOrO4kAaJ7hSrBUdc5A9Zap2UZU
doaY+ht5P21O7PoIadpNxTBwkbCw/4jJ6sVyj1Jcu6ODhluasad4QX96EuJgW5ua
GOqcsjhxqmsXc3IyB0vf5D00ftNiKqKyPnRyAGn24tedJXLQ7PlbaNQK9AwwwaOW
4Al2lFDboJI0fr7YlSUnGy19gW+A2Jzq/NRC2XEIX2wUCuQhqtUkUXYAW4OrxSod
6VtYXzu9B4h+FhyiDdgE/HF0rC081VKlG6HAXW1x6DRrbAKoQ7wUPbjn6G6V+JOX
UvJc98lqAcqDBUeqOv8PjJ0QHGdY1TjdLkDIJmYcYBY5ipWEbGaf56+jBxgb4OMa
VVpSJ5yADX1Lw7nhzDUSvDGo9Gx276URkcpHtC5l2dV2iOMOtt4VqAkq7w1HQEct
u/xbYG43R88Lh+vk9/fAh8m/GU1+zQZJzgJYqfKua8GImNGn+XdY0lyv6aSZVyOS
NDuMrlE6D/hYJJStrzqTLWwq5Zc/w7DoGCECJ8vAbA3ngWBXg4p79uWtVhlruPTO
fumBdE23rUns4A3GAqUj+AIySGssmSNuQAbd75CXSZnrEIjog5fKliqG/6t9kgAi
JeLdLhc3lAgYBJ7CyaapUb6PE0XlWLVncuxS0JO5u6MIbqEuauBz5gFXwF/HK1CH
hM+ohAIretLDqAuBW91leLnkYEURER4j3q0zOCHdFcrtTpQ8PtB8ZLnSLnkvCLu0
1E9XD1i5WfoKhnvjt4U30WpnQ0OGJbHOCEQCVL4NgRDPFxyJgdv4JHmVGshOHcUW
MmTgiMnQ9o7H84CWED9rov0uM0Zqko55mofsBlQcPJwCQO+/tTIwSxthdeDWVm5h
5DRoLnoLo6pElh1QIJ5SEGbjx00xDahdm6YzZOWgEzn66OMVDsQ8WvsxT+d8rjim
jxP8PGUoBx+Zgj3/deHOQrRQ23SuqRoPcG15qprHiWNazFGTOTAJfIf5vtpgC0y5
86ounPFQpX9KMAamUQrRMBcnD8/QDi77Gp0nBwo0znYkAwfLQGT+l+cYOKMvqlem
nmnSxpN9KGRtrtsNEWjegx9NvchDfX+/kFtDqlQiHox/Yvsg+F6uYZq6W8GSB+7S
ioA2eNad9K7V4IYvnN1aFEKwkR1ZVTDzsWF9w4SY9X+Xmlmq7lS8g1uznLK8vpJP
frY0BJdNpOjFFRhGPvciXXBw1wICENHuQZlBKNROUS52ohIF09X7endiBOv552Iy
SHqVsLN+8sgahbpW+13SSWoeDBSdHRoUsZUQWQfWkXjRICUMNAF+f/xtqPcDlYOy
cKnn/rPe1LNuWLg918Q+VTKGuyB3vSroyD1DXWnyXgd6ZUza+Sux2GvB9dEk0qRR
C0ciHkRKLylT6Wp2Z/oRay5srn+D8qZNRH+Nma5GSfdCshF9efeovvp5wYlK1LHU
nmv7YduFx5p3MgkB6K/tOhIhU8+OQH+f1MYrWm9o8D0v3wdaw0Qqp7KXq05c12iN
auL0JPfGCncm23KH5AaWjmXJgMa7oKJeBqKBz2UVv//UeRU8VEsFgTo3iaqFeIq+
puAa6KlFzFI62oRw2RkYYKLVQEF1wCBbAvGqI6sIX33KUwcR4zjKqI9t16MU/KPS
h5pk6mWNXGZuu0klx4yoYkFPdLREJtrjefJ/7gxO30RLKxSJ0qOibO1dFiELpFEE
PRPi7/jCCRsqGYb1ddCuOAImSdeRsL9/ynLYjID+8RbEwbCOAhGjinRbYpuMp6ko
ck7+/SNZaqlw7UGl6+bpJUBELL376lpR4fAvflD/mvGhXSW8dLTfzurFuPCEjsW/
gOyR/zl7AfPoFSKzndWcSxHbuJWgIsI9tsx0fUCORBA3n6lLW423L/UbaLdq/sOw
q/55dafgnGDEaFeLZGuMg+AYg/0T/ln0cwLr9wXZhMk6utzAYYZqULFOgQtsgMU8
LY5huU3N9eiI1W15/MuQm5HUSLOvzypDN1ztYNXqLy/849vj580Q7CeFxfEeB8fl
a1ijmguW5I6Sjdxm/IeA1FUPYjt+t1xioVnGE9woUj2ylcwBQpaY+USm5wGFxJyS
KW1L380UIBOOcuG26LV3r+AFLbPbh4BYN/I5sX0KL9eV7cbpNrqUiSFUX57M+PZD
sGKFJ4YmUkfFv9fq43slgEPlT5zOHNQDdV0jS1OW51kIj5e+PzfOa/FrlbMABus5
GosYgjERCkLZksMmCL7JC+oP6/k2+PZUytDc7GCkbyklCTcx72Z1W78oP6kSHUgw
lGPSEFRvid5xiZBuL/ZO5Sh8KPmVppNLdX7BwAYr2pAqvYOfLoeEKZlDWeAChBws
zbRkghDfZH3QkK5VvaOhCuvf8LC0mKiNeQjGonUetvycBiZ/VaO1NeosaRcQKBaJ
2MpNM6etw0P4UpSCPD/vVhoPQl+7LFa1rxuBvSbJeOY43YB0YK2qN7JpPmopoQzo
c2+lpAu2yVhoBcIHZh3ddqasMVPLEgm4qXL3oEwSTHw2OsDZX3s/WwgA2S/2scQe
Q98OYYAQtmAojOXCM0Nce3dyV5CShogBypgy9Ldz+ecCy6tx+/LZF3J/+TQ2S9By
o9+kfqX9d7ztJdQVpi98XFtf1azfElMbJusN8jdjGC/aWr7uR8FnPk4LjIB2XqqH
s4UefTOG5tKpiGPVTquF2Acak2fPWmnHY8Ethchl5JTTuJ7EO6aAeHIvLvEsAxwD
yZaEvq/UB3os7zgZ2jGuKqfI0fa17ITKB5RUg/hQh0/EkfHdm+dewiV90SqmqwD0
Luz+NCX8qRFoe6DgZQ+PVrD+ofur3bkfuRvO8+pURymnYSnMkT+8n1s6rWZmN3W8
gy7K0tz/bFCjgjxmNxlTLFxLs9p2yHrUWfEFVA+nTQzWYg+o3AO7cosMKENj/fon
buFjjTaGRRPQizFMS8UvfYS0ZWhRpghNAuDmeytJhbeRGUgkusacrXZs0FrLUKSv
YS8hPw/D+n9koQILDuPgQJn+3Y615QfnGB11HCC9I9aNUr0sr8YJYrTeoxHtlcQT
pb+7Q6OYFAwHEEmzQQSnT0BpnEsVHulycDhI/1hmzXz8jH7yEhKP+llG56UI3poc
+qgCBSkTYM2ciFKMwwzS7WoWIcpFETajfu2RWzzbnS0Oa5BMAwNQMFVTtXnQ/mRM
ZYPSdt1vRcjVINf6ksoqpIxIwGA71UVIfuL7xwmRjXcNNCKsYYG7nNUUKam8Wn71
a2fdxD8hvF7tjxCaLq/xc9leyxYItpbGpIxoq8MKIguoZ4bh2eovoffHfyuiOGpE
rYKSZd5cnIucQKXjEoS105NwGpyP94ZP7Eqqj1sz+b/Z++F+qeSBR6GyYsfF5qtq
mrf6eRpV7z7Z+RxS/XY7/Zf2jBrM0ldtNh1pOEjjFIv98lB0isQio9q2HoHPRAAm
GfJ3CR+h+9ngSr+H25y0N+ktFXWpZoVHIk6A9Jg59ktI8H/xOfFANLc0SloHA+WP
VfC6g2SnB1DQldTQ2eb+DWJWdryfbW7Dw3Ir+/QhaEWvg9DezuBqvZKWqrucUbTM
LUPRl4Z2OBMlPwocJX4z96pz9Z2zBQSMbrEzRulrbDyINfzgvDTjZdGTZwVR5DaP
zcWXZuS6/GnjmavokpXkGT5eLPdixQJgzE11xPdm9IkqT9kMDm3eCnD+sEedysNT
u0acfzeuu1mBOS41AtAgzE45EBEvCFTqyGYm9KY8CHhoh3KZmzzbWVlqNftl/wrJ
rudpJGEKPAzFBRnLL2N5m3DjS+q9oM1cCYB1Tu1xXqg9/E598CmBFQx1A4HjXEQQ
SbCFRovrOk3VHr6s8LzsNhhL+Z9epG9lEugPpSWWhM4GEHrFFCSytiig7lDVnXZo
YbNOUdYCRwywKw8lwtXOJjz4Pa2Y2sicGwb6Xqp0EFIc0ioh9vaNpgL6BLuvz4qI
THQU3p78SrN0WLuYJVZ/BAJQKoVZsHAPVZfXeL1emFG7UNw6IlpqqydqpXY+OkTE
FU0TUkKw7cCuWxgWG0T3F2wGQ1wwIaZCGY4jksm/4H1SJRDtHpoOAWqyv2MxoJZ1
hssLW0EJGEWKv6OFL/4X9mhCH/mbw2UW6QrUK18yKU0IjmB3cqNPXGhOQLKOijNt
LtXCL93ZDkx4BQWXYcEnaQ2o7mBKkjhqGX7B+fRc8sHmuxpOwGQPG8qobxmH5aH7
wPqU2OkpNfGfI96qyebYd535R3ghZeoShWhrfu68Qv8XDAVMbslQ4F76ZEIu7IKf
sT9Fpafss/k5IgR97ZUcnnivrd/rnnZe9JrJy2yO71V9FqWi9SXqnm6KWA8X3bsb
dY4uPcGa2X7QVMkucuWCKrP1nBKUdVLHez3k2CjJMzcENC0vOQ/Pv1A6+tI5wXmJ
oyTyojZPdWsBzqSpVHLSvGq5J8G1rIlUiCGb9/nNraHo9EZK7fH4TuC9OQkcY2eL
qXqxPMIHL2HWx1lMh1Pzuy1qZo4pAV6amgZ2K2ngTfhXO/tTn8ig4sx6Kp+fmCUe
iXDutIw4qFIONoyMOJnN4UKA7e40tLwAUQzH+I/KVwjsQMsVcFylGQRvnL1lsoNS
AXEJwW6IR5LPLWD7Aw2uLmx2wkha0wWKrgNiKH9tRlp2AKluuOj80TD8B0A6p+lE
L6GQ7b5tgVO1pcAcTpgx0g8/qIXWTxo1d1XvjSPBDRewIz/QJUhKrusLWOZPP4sp
TDBL2/TDuknduBHpN/Y590JGl9oSdBZTRcJz17NXPGnc0P74tO8AhOjq3mGPh3mr
mxYyVgX7D2CyYHMl9KLsu+Sy2GAET+cAui++hSgAC7EgZwdzoBtiN6TUjdMyNlz0
TVbpZTmpOzhi2NODE+tJgGT0X5RwwDy6cfMIjhV8RKuXjVJcS+JwD8OgPwI3I4J2
EYW+1FrcLwFjtsGQTOCDLQSFAqYQvoYURaTl4rMl3HeDaEzKkPnFyAzKnJehVC8d
XRLQ+IEYgE2fbzsiAFJNyjoQREFOuIFPSEul8RBpeBBbodpCXQQNyX6lUykfeA7I
8ZM32RXdmgYEcY8DdczrPsCXfAx7tCRNZsE/Y+dN7anlt6lftXKvnB+v8bPZD/Gy
4juuW7+CNHbe3+AQsQ4+6LwZ/K1UCj90ZwTdb3o+pVERFwOvAgNWAHJEfazgvKl9
+nP7MFZxMKXNMAh01VuMXmga+12i4WO2TaYB/wB4DNOPwu0G7kK7uJ0k4UELQ9tn
EES/V7wuV/IFYxHnbf6JUjKiVAWBP97GXA9KZSYfXsbjlKtcazVmwBh8i+JLXYCK
tAYMMUKbJR3ykFuqJCvlVnYXU5PcnBgAk523ixpFfZgHjL5wMbW4k4w1BPLvT7Lo
v4VdjQYLO10vuQhKsS+bwzaJEVJ3anoF5Y+LvaqSzuOFfgpYWP5j7klGO7u3iXlV
r3qAxSEboKlciIMXzpOxGrsnCoGX+LShJrd59skptx8xP22HRc+/nr6fCKIh/giJ
7aq3Gdh7n9FLTrNRY5U0kKE4Vh4R/qpGq3y2w992g1qpiHqzXi0Zf4OgJuy9h1g9
6i4v7dqxlf/SuX+LESTUXFpRyAhCpYK9+LzgqZfxqE38mtwFPcVlDHEdRFRHphnz
6SBA6dpAsje+3sYGQU6ucY2TUqE7fnWebSDXug7o8Ds7o0f5luAdJCA/tM8yXclq
9/hZWLMZzKv4ZtKZ8pzoMx3WrHeRZ5xeoBIdib+XNJDZKAV2jlJXKDD/fg8zuK+n
xfO0d9Fd/mLL1YT8UQuP7y/PuH8xl7YdNWn4LL7XbofSxnI0PFTaNs8izDzs9WSd
BaxPT00U7sVXVxbx1qFFSihorRdeU/zzsurOHliEJZyjijKMR8o0vtnDDOrHQdl5
Gltnn606OkKr//qNlWeuRs76KFiQHe+3lnZvKyHxg695oJOPpe4SdfWs+AhiP0gy
7/rPJmG3ydrb6YXK9BZuoUyDKTx7GKn0DqXEruxEsnR64d82dxj+OOtx8tQsT+Br
eVsUrIf3GOXKsKdGFoyHf9I1HscfX2vInJOVItt3GHOdJ55GyIfyGyD326y2qUqQ
lnAvbROfK+OAJYwKEyunNh7LcdRJG/aFTFVfept0d6q/dEX8Ae0zcq1FZYJCTb6d
wjNUrPle0pyBBMi/v0Uwl4Q33iyl7OzyN1gchzJB9Fzs9PQ3SxksfjQCxDFUcrY5
oUUZUB9qHo0H2VcJNNEkFFFgTihOZhmpxOjZwfZ1soqz0pQF5UCyjLKfnCvF5132
1OXb3+JSmEDQaVmB4qA9hYv/LZZnBHw7ZV0MCp9JLE/LBM4eXRKeM/iUKAlvCzsN
Pr9w7gG6HHzUEVo8ovXhps5G6u0GDk0uio0aSLxI9sUDD27sid80qaR0JnMeTenn
EW4ABY6rVie5tgG6Rkm/3T+MFJaEVVUGcJI/iosOz9FKMRiefnhNxYfqggnUFLgq
QqSDATTcLK+Ox7gHeqJmqSte8cPMa+YB6DFsql8Jz2QfWNj9m7w12xEgkXGy5WUA
0CA5jil/0OdrYCB7j2NTuI0zpFNo1WCTIzN9mWtWU5USZ1nWDTBQcg9IvhNJpi6D
uOHkXYxMAQ/pcIqJDTaa2cTQidB923YJs2EQsRKPB4aE8FK9GYqjqlaWSUz74gtw
cyRhbeHO3mQQtt75qe4cm5YFlE1n+Q4ashpJ5kF3HFxMotKGuoxvHplIXU5qjcoL
KuE4IbFuDkxVbTyhxzmWqvzoLMAXK2/FEO6i0kj93VjBCF1sj0oeKJXrbrL/gCwv
ihB7GJtvmYI4EvTEl0k2dqpeb1IQuv5fWQlE+ZqwKgqHlHpZ2wzdlkefaaUR/GZZ
gurJ2MJcM2ijlRiXmgbnDzMfO6O4xv3UEkE3KB0NxqoiKSJIBA2Zgt1oqeKyvSSr
CvWwDElOOAMb3GNnUKwKYwLAwdEHcZV3jVDWQDEfIpoGG/zHxrMEXtiETqTfOOvO
mqrJlfLHIssL7D2/i2wKBI/KWE0yhi2Xl+81qHkfSkj8F1bWHGnmF+A74/TbP+qg
stUF0VCboKpDnHa3RuuATRZ2zm8uJHPlgolMmLzEwgODrPrZY2dfOLmYj2KLGHeO
KAIzxWfnKJb5LGYSYGpjUgbwKDsAe9N9CXyVUY8DKNYGPpVnVo2R/tg5X8drl8wT
qGt3YxLGhaMNVmzMGhN+UN6TcpNYNHp571O6Ao6piTg5GVAtxfpUpZjQFez3Wrh+
CQ+XFc6slDtYUIArmxxg487FvtFC1EUDfBpMfkVYt00F9Lbxf4COqUFtlcoqd1ue
kgin+/g+xle/Ldqknr7cMeiJ1e5Exo0fHNyJdh2VHbFm4YEawsgHz1woz6p4q21W
puauyxfI8u06iOXgjERatVv1tpbwcgO/WBmURFwJ1ca7Is/tFsXDTn9U8BupTbWg
SQ6NArGthUOSlNvKUgQ61mz+BtJrauwQQDa+Xg75FkhtpFHgbYV3rkIiPoLVpNXV
jFy6HX498St8nXXv4igQ1dvQ1Y23FtSHGRR36Rlw4IPt+VQO7kLFW+EmQiM9Nv1Z
ZzFLefwyY9C5bIXyNZdHa0auWpV2xBgtmBcRdzZ/YwH3xZXKtElixQXdNrAa2VS1
tfz3XQHFKqqc/Ceiuzsa2mA4+LkKllb/YyDIoThqCJRtYtv92gQjO0EF69ydw//9
iAxilwQaEZM6O/9cf4nio2vzdKhB4HNLzPSapjbWap48s7/chzg9eNQS7IpeyDzI
rWhOZmGCtuwUW9jWGQOJPBOqkscW2s1LpyNGwEzwR454OIAh0/tK04vS4JDmqYq5
6csv//+yd0Bq/VIerO9Go7PQSsxvr7eWcHq8I+6nhOGUW8hXZLQISYxmDw8OloUn
bFB6ARRWrn9SAPQ0zvOE2Ljynd5YFvKOuZl2wMk4ns+fyJCyZrdwcwQipC5MglSg
PHrsrOO9lthyO6lnJ1S7cCKYsyTR4dOqFUss4LrfJ6VCS0naCal3aN48LtpI9ZfO
dAA2jyPm3jPGz/UdJ06ILWTYzvEeHr1rqfjmaHFRzaj5zs3hb6o+fQGWbNaOnU++
enCE3/SX2a089zRNwlPE4poeu+ic9c3t0mGWtyhlaf7F5T9hqBPkkmZyVwZaddHB
bcP57SnIPV9z6jIxKcJT7fvzjkK1y2DRDDXHqdlzrt81/fZ/6GsZ3RH/avmY+WyX
IFgKlWBleTjQqBlbzDeP95wBOgusXC1nN/zWHR/WgD3VHHvs5Kb3dCmyiELe5pQ5
KgZh3i2n/o/3Umk5yvAKus2Tymzk32W5O0a6URJDOckd0lJvseI81gpjqRRSkvyw
1ezcK4JwlBJVWXeg6BKAF9/t7Sp5rpPclYxRp1+8YWs7W0GrDImTrgX+8od7cmSO
9XPe+uVALxpLvYaCyrA34I5/NabMBxYMOGZKsUWKxS48XFnSgiylWVHSUXkbkz9w
ZXcGu04IoRjdY5UF2r7L25MUduJNyKApqKE9Qneyo+qKaOhlM/xMbz+cJdEWHUbK
K9yGpRWzE5g9BkuIotE/gukjf/UROdGFOYLMfUC9C1igEtF/n0wA83F8KyNR2QJx
UfxGsOlqZcAMrTy360SNmxQDC+k81BBkWEcY+4l+s++JjepBKPd4HkHdglFLEA5T
2W6dYgEtAZ5jOvx4rYa+Rhl7RuJyy+V6z9YNUyTC20iv7gR8sgt1RpM2dTLXlPu1
IDshvVlOeOrZjgHmOPoi2NbTtBnOcuvbtx6qgvYg5VRgy3AasxkgysSZ9vxroGj6
4S95FthjLqiRz0Mfp23yfXjTJfNyHIjDm0GeTxJecZTZFXajIFzbw766mSxyjLjW
CSj8W4OqORF1txZ6yoLB40mdoc9b7IkpdqSGQqHgAqIi4lwCMcoUezQOJ6rOHY1O
CDtMvcuEFlBJWPsCi6OCBnbftHq06pmXHxaksABQzU69JMdk0ttgCLniZzpllV8u
9bj9QA2+O9d9I4k2Lnc0pKOiROw8jbFX2VyrXOJ7dUQke4bw39spebHsXF/LXmtP
t/BvHPpCcX7vrRYfOBNALUj3d3eLKr92sdAHfDLVFbRpe5Tx8n0z8PXgdx2DGevG
26IeHYXU/PP+HUZYwg+4XEDjoBsLIPd0I/kFjtLP3KsoI59NbQlTL1mbTDPgIF/J
2h+kXsU/LhWRPaOs66ADaqyErwhdEYHovn29V0gtmUlBIVVKfXmkc9CsZ3drcyPr
759sHdOCF6MDEDjVG8OqKIYKC83QZ0nY9Gs76rceC8ndFcijzV6ZEyQgjD9FXsr6
erQrntF+V7jPZf0G0tWuchX3W/R4s+w+GemA3w0wUR69f7l1HutVWFU4mRuTZjWj
SB9/3LTDaCIJrpKHDBBk2XYbVWwkdELmraZUXLVY8asLIBQNmyQyMXjp6sCsFBmZ
aBZdx+KegRNRWRMRemMWlZ5I41FYoj3wE1l70H6CAjRS9tyLZnrI09Gu/1SXzIqJ
EghgXRU5yn7L9mPU0XkqC6b0lSpi70ged9FrBhhXWK55CmgKtrsNQkAsL5sLeC9/
qZCN3fHbAc1rW7h5J1BVNWzhOk9rn8X2F+cvaNgY3Yt3Kd7JBv/okV1hCctshode
54bkMmExTFaWLTyJryRy4yyax1msibBkQvDbiF7tuWkm9qAD4oFg3NhcbrwKZRrE
6MxlIr3diGAjJXwKmcn6JYis1oWZ6O2AtyTguUrwfj/zP5JPjxmi0axq9bWZ0w/0
K4Q5ZeWWMmivj6yc+b6dtgWwTVPG7RFDSEhf5EXAJNcCw4HNwmkZhtLTr3K2HcO7
gbTfYp+X7NhaLXBmrbwGKPBWQ7CQHQyenSCJop6R8ZOt3i0dsYwVVP/dFpBEQAEf
XgiaoNb0n/Mif19uKvo6v4lttpXEK3HzPwppwhl5Mwh7czd7JnlwwMs5NmQNkagO
J3gwX1ErRc2xk9UHKlzQ7Ekfb2GmT1YQLFiwKWOo1gfUfXf3y671WChpRwuoJWsh
LkLlQz/9U4EZcDDrs5bFH4Hqlz9NRNppNUny9PLd5nEvJYOxw7GplAoBW+KXB3sy
vouv+1c15zTs7f9tXrfYFR/z2NccAPhe3iQDgolovAqlE78VGOv99yR5GH4DkoZB
Bi5Sp0b/ugFwNtVcSFGjx3ovXBcaPohWYDKjQJtiWNmEla8gi8wwYaNIbT6IqLva
LUL0sNZXHYtcsIkCwsSDJ6w4/FvpisY4s2g9B0FSneSCimw19Mb+ofYpmuo6BcB+
fU3nwW70q8DYL8sFxMQz3Td3MVZ73it6HGBTpRAAKaZRtPA+sozykRe6IiGyKvVY
WIQO8alZqjzs5VEhnsg95Q4gusApmrU3Bzzb5OM89fJmZQ1DhNZca9soOhtFn6Wg
oKcdlJ+JxA6nyGWpzioXy8bfj9Z5karbgI8DVW7Zw5cso94SIpbVag6AMuOCDYj1
tlr9PH91U9ZYJAWZIPHl3eWnAO/sAGAYw8q9171JAVpMxjEKCgIptr5/XRLcBunt
MH7eeJ23g1S9uRigRvWTAb0YDSr36GmlFbtxTA0SO0F3Oc6CxsvrmdNdJ6fGsqgq
VUMhcmvWOSyGmJUZIzY9e3+9jv3NhFsFjf956XDFVXZyZzgj+jVLtzmuZHiYZxCu
xYZ9LtQInygd3EoNk07UgMQzf+wew8pnBRMzSIdEezjQdEQXzCesDuS/MMG/DuZS
+YCHEz625XRLNMU8/48OHsXRr+6VXbLld+34PE+SphCnJSX9RLDx76HG/iRgpm9k
koRbRrnw9HCepDNa4vgW3fh+wJC3v6rYRx0cuPfCondIKou2XLOTN1e+GJqwRHl8
2wqXQUfiT6D7B8BmxHlMCQl70iJYBFCmDczKGmq7kh1chdVcqedx95Lomhm/OVQI
vLcfPTSowkaBL72PMVnLE3BeaFLy7oaOumDY/7+y6ZdOyMzZWKc/KwfWV8DqG5Og
7QkQgfU7AhfiEzIdLG4DohdmwCf2DvBEbLOen0X6nRZ7OJ5m2Nr9lmwG0SMdSbi7
gU7iweASa/gF8mJW+bHu39hrFRH0Hc0eOpACAnIXerjwaZvu7q60z9Yh/Nm2t37G
INfKwJdai9Py2EUlOkON7wSmQI0Zkvj2Mno3zSSk73R5KHhvEm+K7jJVBj2PGKXq
vQxGzLIYDax6OLIoixbXpRU1Mf8H9kbMeQzX26eyAHnR9Pn3/ojCHP+CrcI0/Xe+
ErSlMn8o1+A6mlOV7aQeoC99M9TXVOdQazGzeuYwrGN0i1Z3gpaGUU1VxuFoNL28
gKcMErRP17ljO5BvxA+1i7/zGzwbkSBJ4kODRjquv+BMHxHxe9keonlNlJwQgeT3
0HdYRDv6fUFWYRG3lSiTRQ4h17zn/+3KXCWm1Y8ZLoX038/abohByqZ8U4a3b56V
0UAFPVfdapgHz4tOIaoLWJFamSOzfinUdQpMSLLdTGTizwNs7UVLGhyPYHr1a1eu
OXOHBzAoA9LYJJXtQULvEtDBC5zuvrErBD22wPgvqRewSjM6yDEWrpnaSMNF27ew
gQCysL3UC/6wUl7Ib5vaIC25+4iiaWG0fCZ9k3ZIntjAzYSp3RabS28Ecpwe+O6O
sgl5XHbkowy9s+RKPuZdsITv9oe03Fjq7jBjw2lrGAZ+5U6n8Q9wHzochiZP3E35
iGYbSYLtlk03BF7Bod+FZRwExozu9hpWQ65d/vH//hzSh9SQ6jOB1wFMDlWoOSV6
9TAxxXy+pwwrMbP0Jnw6C+8DXnFZrE6CHk0Ng6cIkWVdmM56H61lXf2MhWJLtzjk
gTStB6IpTTmjePL0Qj3uzMi24DyAMgcUQtTgEv9tDppqUjPaRkyFFpZQlWFKdlrD
NmWRkF/5aIwvGdzkaEzrLe32NuhP1OhQ/nmxXemlw5mqLbEVAH0O6GpA5qcTeJj+
M1qZ5xFlZNqhSSKIpjmoE/u06W5LsFFA2GMkeOJhUhOPFA038uQEP/DA9II8rEOM
l+OgI7dV3RLV4Yz5jRl3Fi1nkerT1e9EiKh1eKVk+ZgxCNGw7qV204Fz6t+vfmfH
2eqKcu1Oo2mBoB0TOzbh8AljIF2MSu8UrKLXIBxj19Cq7nxJQMFbTRKHR+zeaY2o
lWxj2I5TFYxFGmSus5Dp3DiOZiHaGaCKIwD8MATuvtlTrYIgkgrIOQFRl5sWKLoC
WmVgHR60wzrJeeqNmWwE4qDSGADWz38qK7r/uIWy+a9VCoxKTsLatGhZ9tX6HHQy
ltHIQKRpCUJlxZxmiyJE9raBUj0W42sqaQmThD+EEWSdKjehMI/g3Hb0a5toqVKo
QrgDNAWXL5WrXTmvPUBLqMDtNpqDq534XjlUyBZDJZ3OjOHdNjCu3nz8afL9KWdv
2B9mf1nC4TvgVri7UW38ilzfzcWNdJJx0TcPNZ7FxH5UwqPkgzZ5O3or5RNO7Hpv
bkBZFoTRRJxWHgrEgYXRv1ZFYtlyB04nzlKpoz3Q+C6+6fgQtBh9jKI2tGmaUk07
mkKqu5eUswhY3CDhgplHfQJ3Ko9qukduXPa8yXMbhApxjoQEA/AZ4vlRya34NjJg
U7cwGRZKLE6/lY+3N6+H7g0XEhl4py+ZtIqKU8l09sHfAhAqJbYiEJ0ITXXc2R/t
3dnXTlLj1QWz6pDOLoYJsZ7wyAmIKEWAmSPivhrAwUOOmbFdeaq1vWw6SyjJADg4
OyWt9u/KV90+sibK0rprnr1Ol/g7JFGvRJb0+7dCNewbDp6v1FTAbpELekuepp4R
M5vBKJXxqAxcVrgPNJ6cSnt39wAj+NENqW3csmd2VK1tNVg5y0OUwIUoByRFfyvI
KulyqeGVRmXtQmIlLcX5p5llKYHiCre0JAm/K5DNIDTVNbToQEQSvfBEBlP8bbKc
ZuoAZ09cUoneKlnqcOCc3CxJb+YAaCtdNIwLqVasI68ByhTvN0Amwzs6dMaqB3ix
sPkI9aqWRDWMg9DAGNtqtx0stLuTOxXwSsTd4UmR1FuDmEkCwmMtFrtlWvrjPSu2
0sQGK396rQfqN5WLfBGSLhjFtPyJ317huoQzgtb6TKo0zi6T28N75a6QdJ6GFTzf
IS2c0qnXbCmjBUFl/L5IPMoKKEKMkbLZhNhrBb+WkXGa6jvCvmrLkO8YtHvHkFSj
Iw8C8xXntRD1gVXf+I4ZDXBKkRFhgnk+SYpWeSTtYD1zeQxMuMl0TWKxFbrfZAzo
G7Ugc0rDARwun9gvCzmL9f7b2qi4cGp6u9Cth99KZx0xgPlFZIvpyX930R5yA2M8
+WsOEntvSNHLan043TznCxZK1a7JGrfzNkEHlgbXkPqzLcOVufHYNH6qEf3aA3S9
CZAwVDv6Y3T86KO1CtrEYzeUemPaAoYmYmy3U6XTuIvLEn4uDzUAtYrliL1EN39W
HXNlSeRzoj7QVjMDKfBKzRBekSejcV2LFk0VGgkLqdGWvlXJZbu194fuJy5PEK4L
pCW+G3wg3asjmXiK8KgsXNc7WFgEc5/pwR665ceiTbEAElBi7pPt35qd7bxE8qTc
O2K6b+4rViiyOQ9LhwF57UV+Fa4mprlW4AgRB/YPpMqP66ltkbrNoV10y7nCXjoU
sbEIBDFK6OhrgAOGWmKdhtleIrdrAn3OfRnu5qDgEYmogDPZNlC40nyN6JA0D0HU
Mh0u86vbmcrkT9GfIAkcs6R/GT1eecFZTi27mqXcefodcHc7Phq1bDqiMoOuNHjT
tZlgZT4/e/fXjtc+dfWXmSrZzQ4u/v0kS5pFCSHJcrjRkZgOHp3oK0l2D/LUGkK9
4dkyHhqpDAKiax7Ylz0G23Jn4hvjwXfhNMpW1ml8NIxdl72wQ5xpFv47GkuDwPoC
c0tqPttFCrZQfD3clq0cjk7b1UKPBoj5YfIPNaN16tQZYKzxPSnugVuou9U+m3sX
fbxHEf96lXif/H1NNeOdtC4t22JDmaImgKg38B69Nqq/tRyma0nc3yGQMOTR+utw
ZE0f5G1zSWxk5VUORXySgbQpY3t5slURLoqQM0EGNG1JEtyNjlNnMHSjd+LEaUR9
gU2KaMFKf2yxqfY8QFbxfTvmMWRtByrgWdbZcnKCkT1JPdTPPHeHiLBimXjYngkS
H4Cb28L5ZO0n2U3qifpbw2xdIlfg/Qy6W+NrNChz4bzV4g2VjtKxMabKhpZGdAvC
xR6b1lP6K1umlGaDVvbuPCJ1U5IR8Q3LGRPv8D7ArhQcf3P7Un4ZISIUdR0r/drc
Qj60DGZx9oAF8g4oAT2EK7h1o8xFrp/Ws0GC3YjrCUVPVjlhyO3M6iNzXSrl9ZJO
VEd5azXf4Wl/sDLselExL/IWDzBt66E8kvBLhdd8RhQ3byrpJnmfAWhi6NDXpi0j
v6Byc8HRejRraSsUh3rJhSZyNvCZUifTIwDnhBveoXsuk8H4w0HFU4u9C39z533i
pVuyUdDiGooM14eiBMakNIPi4dUmoXFkf1lZVSJWmmRZVm1Wd3a1oSGPonoXH+Bj
GkogZDCwzKXl3GQSBgkDGndRYBUQ8gKea3mF/aJr+pdd2alPD8jer0WNZXMt4/3f
a/VuFhkqIua+20d3o3Ae6q5ORI0GEmuOp+DGiZBY/ZM0HWwQ06e25jAZcBCBxNsn
9JUEGE7Dnqu7Xw7Ik5B8ofudvfFRJkdv2m+Uu7/M3TXYJUz24q9FOUGgCmikQ2bc
f1DVlc+R/kX8h+T8Hg6MoZNEqum81CHS2Z7PehH9i1GKD5nfLkb2sglVbUmTbg2a
D5jOr6aosnzNCJCFskFa6sKw7EAkiVUYC8/G5qCcg8lZ+xNRHamQfeuIvhRIfilR
PlTWOzZfQcJa92hkpp3d85A85rOQcmjR6eB56bykAByHSi18lU3GBAmO0BxYzxS7
Vsh3G5iECNbnnnl8RMTtZYA3t8QLtFBGZxel+ZnX3ubVw/bxyfh/oRLP7DWaaHhX
B4EkLf8lCPPrQ1bjuSaHZ37OB1sDwZNg3cYju6jFk2+oTlb3ciwAokdXgXGLNgtR
VQqvbkZAbNz/Zfw/Zu3S1frMdsN7wa5y2hYZSfAD3bGrwagSA80KgjOt2WnetJ91
7sdBNswaHhaI4VlYr+z7h3IzbEKSvvr/NQ9G7XMUTYWAlALbZFhUZTi1ruV5oeQQ
01ON0mcsmrsB5jpuFOxydnx2BAYM9kvhYaW+BIrUxh5R12hPo+4XRmBkGw0zJS4S
uxbvTWsj85zTr7iRG7LYnfsOQkik5zfm9KzEeRls52+b6eoVLau70zRFgNlx4I3b
8Rb3cMC3dQ6pr0brfiTQio6MbpT2c+cKswvYhNS83kN5W9nqwpH9Y0jmlXl4rz4w
nSYAE77aa2+RSQ/czCOVXVsaSEyNbIjp2IfYQCZtbgMf55yAMB+Uhj3fAbypKNBe
qITYM6W2YLxQ8rHnFYYlt5R2HqCoGtsCW8Py5VV8vNR+4XdVSbQ27GpC7Zf/DRjV
NpB6qNX/NndWZltieYBSH3UQean++uzLT8voX2QE7Mf9TtfmkH4HpZxdu/Fh5Q5j
BNbQYwd07fmduHlenKBabEV5J4NZPU/DylZODVjZJ7D6xe7bQeD3UkVzn2r44zKH
IRH+mqogVVqCquh5+xaHtgGVudUX9PA5nrR3F6oQ3CzLgvCeaAFIlb3l+noYx47S
nXBhFwGWtp86/xXBYB1+axYKUi6FfOBB9ljjjXmtK4WihktnHXIvtbayJf6OTdgp
bxPIEPzBXFehhVaf8MR4VE6z9iHLoSBaM9J6y8+VQDYc1vIliZzcRpEPQhftvGWS
O8ODIY1ckZgmHON0hA9yTqVRUHrJ/0LBnveiRVJFQiJ6rmFHfGd0LgP+cdAaPfLX
NAG/grkz2sgBz9X5ZqEBun0IeYfPyujQ33fXHoM6HnHYXIhYLjUdRfVTkl6ayFjE
ggv5B0J00hXn8zzalIYqyyGJZsn8B9odOHUvN6psgQEprzRvVJuC59xo8GnUQY7w
yQJhQUpME9hhiHRszbR/Mu/yHSa5jstQYH/ZXC5LoxnvEIGcVPaG1LlHltnyxnph
Hirhu6nTXwzmEvx3pRPMJkWJGKcbLwc6xryMxHG84wtD3C1LXL2ZS2hG18Ynkqva
/fke3WUlwq/CEOFvPW9jirPj6qrdTeX7gys7uYFVHQPIs5zj9t+Pg3TsCZHAwHBe
y0vOmZfn5sOfbJF9Yi76YPfw9SipnVFdT6sdP5W6ZQxa8Zr4ePS8HvRrxggj1z2I
C/M80Dm+g9IxxZnmf4rmwK+4xxEHoaJZHn3rapxuTPZG6+Hw29PP2TS1dQEgchna
4Bhb0Y2IGerMM+6byihMU3CuJne3eQaVz06olgQ/s+nXj33CxJITHyaF9TZxDK9H
2rA1HWSd3g8pIJbpz6PJzCWPTuhKHtCQbmcyZjGTLETmhkXAcyxdJPctj4xLhHXw
AeByrVLGndNn9B+AqNmBlWd8MbU+r0tZbCWenPdBgHx3TTt8nFqMiZOKmr/o6sy5
aRmdvY+p+Su/cpwKm8LiUKmEp9My1ANv38bPIxD5WkNik63wJgQmW2mGnesNZ5wN
uDzAFhKl1jFJvmhJKP0H4mWMpStJYL4DZHy0Slb1S2rX3kbflR982m+7GQMp2RpK
c4lDWD8HwGzsqvdQDvgjH3MFdOjKZrjwpGeuj+Bwr0LxLTNZTx5rPbWmvqjvRFQh
MFbttSnN2UOv566Xu3hg1dGoYftYv5UZX7FDYYgTf/BBYTtGkFpDXrLW1B70D8DZ
sAQJffpJo9YIKCQjstcdX9vZblD2RGRrT45ZAumjMIpywt/rdGZXnh6bSHbBt8A+
1LGJZS4YmtQ+i4cKscQBYVflPaGLiaJrIJlYyjY0Gn3txwUot+MXWvOdHzNQ8SYv
Q7A6JPluG9ki9RsohycdDuNEFyCCZ3M4sD3RSOYpzB3OuJaLh+8T/UfP2rrV5hoZ
0PBlXwXL5TXba5B45FgtXgpYHySw07h/Wu8vhgqMd/8sGxNmq9tHWt9ZXgEQ4KTB
NvKgiBdHrruvv/B1MZyQ92bvPQlO66sIvvEDGpzjhKNsOy8cKriov6ANPdZfY70v
0zPlbKUCJ5n1J1cXSH30nj2fZVSmCTv/hDBkAZacZmrevKBjjQlLFqqbSVgPBAXT
+EXbv3pgHbxC5ccJ6WzSvQlJZ5dbqcR8yvxY/HrR3Trj+ESJ3EjajtbX6xWaPD1C
YKk45Qx6+TqtuxovyMNH1gMHBO6JHnlB82AMHTuIK4WkiihlJpKJRnKFgbnRp0Q0
z88V5esNGL4P6+wkNyFa8KJbSlFxb/aX6OXyFiPE2AmvnXFVDgpG6tMFRawUxFrr
ZpGfSJWDWNJIO5/hiaoIeQUkN0fLq3JK7RcaboUMtqR3GqkMJ77aQxke/k7EYjMO
GTtAe9gEtmGgckfboxRfzFyN9KuynsP7bi6MHoLhmdWFCzu5bFGt7Ait+hbKsjZO
GS6M75o88QDZbV1tqd4rnluZyp1LCBlRelQtHLduW0dryT+E4be3vfklrgAH04Sc
XmHcFBT5sizpn0pTPNjBS43mK80LdaZSxPswVPQC4d7CKqZDC60uzWwCPfLaabBa
G7zWExjdXgZIyL86qcMBz/tEevRcIKHHUF0542fjzbGXWnfnMoF+5Ceu4t8Anp5Q
slTVgN1119l+k4HNWNE1fzsdFMUkskev6P4eOo6xfzBIbS+nye1WEYRnCVm2dbTG
jXBszFZjpzrIhLkL5uFveDcqmfTpuqOUJuZYfqZudXRa3Rp48j6Ee0rjw+xYXuQj
EswVHN6Dwqt8M/I+nBubc1/PaLr6mbrO2UOl8gQ0X07IKJ0pkVCTUvueBXGQaGWX
nEdtPSYw3lwUNcIfL/lXvG11Q711Yf7ueEp9Kun6rwM1wI7Hf30+Gmn+H3pZJwtz
JdkexCv7SyQKTbW+w0ZfkEAxY7Vzf1zCg2eouGeeykOgxcqKzN5qkXklwhowIaGJ
GjeHxfqX4Pfe6VeS2Woa0ms3SnchU2tz05MjRJlFKVoAy7ZJIDCZqwiBL0MOGck1
zv5TBQBG509hLFm/gS2bgd0HF3nbd8F/NojaZubfjQkM6zRp9sMuLHjY9N1cAdMW
LyKXGMnHKMdu5z5f7aV8BKkON4lF1x5+LNk2HzkV2S5br7thrbHeTqtRmOHDpSeK
6y6fhYcPTFPdxxk8JCx1cKX53tkfuuCOJHFOULARspm9kZghCKWfE5qfqDBgFKVU
jIX0gDhOHADAOLkMMD6992Ydoj/OYXLe7dN3mXVj6ihP/vM+5oqsTd+7Cv3YtVpk
uXsdHPvYxPUt6dW+pQenOV63j/PMut2PQ2hKLSwN17l2aMLht9HteBdUyfdCmget
a7y4UdsmfQOCkkGdTq5qNbiP6C1MqMrH13bRgi5rP47h5XcUqqmPZmnPhRL7k2/X
VXs78YMzHblCEukpM8daT/vP0JPfE49FtmILJaRDY+rY2N76D37fz4+jvIROXhhp
jVLQiIDb4rnVoa9xrkXD6Fxz+mTK9oDtdqXbFMQYqWF1h8S2Hlw9IE7jzQmyW0E4
6E4IZpqzDVZxGh9HouOlLTYboe9hJCErGtCketVHK7lwipS0V/6J/6M3g6fbRkeJ
b/1dY8DWr/lajrdbVRCWsDfXERbVKYpc0SewqiyWg86xd7GA4C2TM6Ntx/tpBxU+
iEGllhUrpZjojdd+cNVtM6fa94Gei9OI5Usz9n406v3dzapkNTekayD29XFdr0QE
vgFbpLevCDB/UDJxvkF5KzHx022NSAxBY31zeu7d/eL65qu8jjlLAbkAkYAb3WZM
U50MGscANMtlgBQYthIkjcIloJ1MhZJm+MRaky6dOCCglGgI6KNDa6hNfBzoJcoS
h3vQqIyykMZYb1NLwilOg5SjnITLdSndyp4UtDbFLDT0m9p4EeJxz7esi1hruje6
D5DnyPecfvBCNyctTi+R320gMs05US2Cs8c7b0s9YO5WjcbPXX9WG7yXZqB67+9j
0L1Nks/xVCiJ+dlYDjRErSgRrCJwnDJXF2qjAqNeS6yjsfxmuaTpGAALYybzy2dV
ODGY0Xhr0/lJiTMetVqkSFhej72XcK64Iuo6P4Jf2LdSAk0aaB47Um2haFXbSbTT
oQKUMWSgghbEUi5E1g4gbvRCluByxzh1c8Ld14QxShxlRLyGLVeCnTaxMXtxytum
ajZd8m/vs7jv9HylTTyhdAvM19fZYjNaIkP1yXhn5RbXcwFkuBSnIbqhknGMpzmV
ecvUUV52o7+kWz70T93J9wVF/4z0qM2/ahS0j9wE+TFGO4Xr1EaL6qXrAapu+DfX
u2/uV5p+nHfdfm58l6sYEbIoO6kox4iKsfg70Bdy10J/FJqyAWv5nP5x+vaAWkCD
tQZcWmsqgz9RLdMxpg/VcmHrdwAczkH+g70HvLLtneYZ16T9d1YoY82TdqPRYxsg
RjdVPZwNlHxJg5QXz+uYr7cvj1yBxJbitXcpFoToN2JLLP5jvKIMfXZkRdN/v94+
wEUV/1/Ze9VZHJj1qOJy205E3SUkRPvR+iTQwm1EpY00drnHiRFOxzxyqjHOc2V0
mAtW+B2Q4gGrLxyojziNqz+YkASS8Xz+NjDjrnJ+fVdW/3HuIe5X+iHCwvvxUAam
hnZBdK+5yNNvJCz3fRwNHrThFzJkI5rh0O4Shf+TnclRrqpc1ZHcx2trUJqlKKup
GcaG7gwetJx6ycA0iJetgxkccRLPB4JrZe2VP4hiRCXh9VbOHdnoDUvnfEPA9x+Q
PpGVIkzqlYQeuE5MICT5VgyJGwyOMD4cjgL1jl0Pt8asmPb6PDoD3qkEWhExmuuq
fEhefOvx/V4S2MQtrVrA5O4nPtbC0cL2TgG/eYauQqyAPa9H4h4/6AEAPDgiVHU6
THf96o5ZDe2m0zpsTr6C8HY/opKvtG1qGBmWrUI/TZNXCGj8rJsbApj/tUjXwkrc
hoi5uLHjinFsQG7jhxChb6nhN2w40aEgJrySJhQ+tXcotLJIZWFdCGneD0fWiO+B
GhXE8ycQNa5wJA1qTHGtHpt2OAUOIV1Vu30tqDlboMNvtjSsLhaXrtrIVvXKB8bW
LVwjEGkE81wAZtJXlNenx53Gsc74COZDOqefAVZJJrBL2mjqsEULcSvkaN4BCvY6
OwCBNJkp4+tII8sTwZteakDZuIqPGwveHzz/sph2rw0ktBSkJpWiuoAiI5PuuvDv
vExNX9vWwS9Ty19ckdSDcG6Blg1N5l8DmUIxt6p5KLa5vs5D4BHxPvhYxIEyjfUQ
Ls3ImkR5cdsH7JJOeUOvWkhTdWlHevevt027zdM0qGUcb93kEZCKClTqgvaEomeM
JugJq7oCD+hPpxiwoXG5Mmf7GQMdhJUfv8Oly2enqBBEyUptnXKjB/Gps9aIKfoM
a21y0HlAsxUxTnPkMuuS1RkEcIFFkYUpKX/WLgUbde1HoPm013szHVI5URFifZTz
9FqJmN1mQRVlqkVRFoLN1pDv65US+hlDcAfOYigukpRplgJxbwsS1A1Dx8klUiu5
+iiSrYf+p89ZiU0L9uQ/Xa+LU0RnD0CqVYsMTIJezKXzbeWAyJFiOm4zdrgXzvyJ
oqu40B2DmSAVt2ez6LTtoIKTaFCBeWkT1TSs+CBM8E3mSSZHLYnvyGJGbkN04z/E
V7F6zNv3xlcLGVdkDX7ElKlROx5Qaob+6tn7asew8OeXTY1MY6jDAP5D4NpDhPsU
C6hsS6kXymD8fmOcQny2Cnrkf6i1mpPvJiBhPFVgZuimIBsikENQ1t92YSt2BlIh
1beJn9fpJTqR7tcaPpMgcfGItQg7vXOLRJHYX4PqfJeSTIRKuhl6LQsNRH6NwPsj
izAqhfnL/xO1OzJzUbDmArKRCD8g0XQByk0V8pdOZNk3JnpmOQiPcSgHVd4qk8kT
tD2uU8D9cSTEclo0PSKxmpzeF4KjwEbIo+yw6hbW2Q4t0ZXPswRlUYMss+slU1Qh
2zskC4U/v4vx5o9jx92/DxX5WA9sApvVgF58uuhh8DOFGjDXiJVAplAvr3QApkH3
Ln+EWT/aXDW8Y1UWCUH24ksUkoJARZLzpMjgK/v6lzGH0gkmzJZV3pkJoJpPsbm6
Z6FwoTHffnH/wAdgKUVttDDxEATo7WZr66pg+rne/apCKueR3eC3lSYABgnHWnYq
Ghmrjt/z/Ct+EXtKDoHJm6bRAJXsPT7RBdcx5eLKVPTRQ8NRovTGCCPgBn883+aB
j/su5YiEpJRKLBart4eAxgu0Sz28VSICxXLkgJwJ+T7wUyIIIVPjWodUvncoxhzz
y2zMvbJLIbNYC5yK4jcT59aqXhj2omC6l1C7bJUoff8gKHJaczc7FXsbJncjrKhr
9HpT1zJ5xUZ4EYWyDPT+7nECXk4nwf6WhhLLf/bAMARAm/dzTCLkjSoe/28c6goW
5mEYYvE4GTgotHCrlGGBbCRwIcbABG/uPxehs4Hlm+6bM8QVDTatw6UEyTHZcmtK
pETzIz32pqY7KoiP24s8I6g5/d0DoNTM0qWI+KouLrjyWnlowZvTgQMZgID+g/J7
8+8tLZVzgIhfs6//3UAwQMzVmb6eel4zzpGtoX8v8cb0S0iMhGeZqKWwgRyN5U+r
30FUKEeWgrusuGsHRQVj+sBpdngdf3rEJX+u8jSdY3pC8hxnH5ykk2XWv6f6YM9D
lufc1Wn8RbjcoHMFi3Y4PAC4NsqryDSdWiFjC7KtqNKWEhpKkaAiJ5K/28OS3AGB
oU3QJipjNBqor/e2+CmldD5PoieeGMihnA8cCT/zcs6YGn/VN7NUFDfjCXCMdwGu
Lrifgn6db8Ps7YJ13h4oaaiqIUKkMlLSW1iht3YjaWIJhG1kiQaMpl7NPricQfoz
kKbF7luOo6JbOr4lk+3O8EE9nKTlFOdsUhpOw7M5ugdktsWJUChYGM4Ni8FHG/60
DNj9Y8L4/rrsvy9Quxnzs2q7Olt7aFibhLjz8+lT81DbX0etRt0yUfZZnG0dZioH
uWY0Q1wKklNQIc2BlT0vub6GBEC0iiwgBnlGCnQkwqDAaa8sYGXlIjiSsF9/W4PY
TxanO+KvBfblIY7oYOTriSa5nwHo9sVUFy0HHwxEgO6tLA3NsbO2Qf5J5ta5+Qsh
HNqL4el1KaavBBNWsm1S66OyzvFV/9SnQCjlkbXEp7qxZt4l1q7VmoGb+7yviDXF
eoY01LgT9WZtXiIFImguhsUPE7sPJZ7nNBR0fycGpByXmtIOOqQKZivk1YTUyZVA
I/SYtWnTjR1LXvjbJTrJSlwOUOgNCL6ssofsP+wIMes8cZD4ZpnNk7tUD3OTNBca
x8sLXKwVNaInUMSat9WJkpQHeg/IR0ta8Gh86ss8v/o0LJTLBkwo1JW24xw25Ye6
iSMqbwjubbsaN7e1TPnh+7zZabplnlhz+FTByDLDyGXH77w26HKNWol1heqpYXLl
7P1pCYSwPU/4RucyzGAg5wCLsPC5I56TpcRQwB0cmJsMMfL6AKoCC2zJwOu73PU/
7ibT/6Q+gWy2UwufJdNjAih58LCIaDxP7jzOH+76WD0z6aKZLCjyu73osfhVNUxl
btdsQAZnnlfIFm9x8GwcQTMLBtlS7gmRAbnroJfX2p0y5x/vvN/sSJD8QloAeXhK
I5a74qNc1byUZ19TumT1yS4MVGFYdTHxvRxo2k5Q8yEkBa/A9dLwsrTa02956BRP
3l0nq/tmmyr+Q0Tu61aa3J8CaSbYW4tgT1N+6aiwNFvZ5lb/rgmk9r43nqPv/XEM
+8J0afXofuajL9+4SkwMecjFFzLAzMw/iiIG0xsCiJ5Ycm3rBWFXhgXIAp2CngrJ
q31oXZGD15jT5gsqCfGen0jml2CTbf4xz2m4zZc0IbCJWtT4hIOzqH8Xw7Wux/YP
l2xwyYQLzPfqPWX6iDd45L6eRX2lP7VjHQISR3bdOXSc9EElZoFauNwAsSsOm5vY
FqddmoYGG2hmHqUuOLB8WJGJcKVsj+BPdPDW7bESei/tUG+E+N/zZAWYDMSgNwOt
EqDQ1NsJIApB3Z19kNegRcbxHAfYTaeDxqW0434bBZZklw1gdLCqzgM1KqXW8dGi
bDwKHza3kY4OUTfd25Q6gGtJqRQ90QozKQpbJgUk6mM65DOFHP+FzbmTbM4I+E3g
niNgb3NahjU5hqDyMmRQnPags/iUG9IPgCfsItHHF9jqI+SyUegv0YsYLx5Z7FI8
Q3G6soRh9eyoc5689nsmFgN0c+dHQ2oyMIc9hbpE40RnAec2Z8lK7sUYncEI7kcs
EenlZc/GHhL1KqKcATzB0P5P2PKaJqgBxWG2PGaBEaa7BmeVvXvwOmaYg72rnD9h
kIWpgza0nP8nvjHSYSTNVYhDj7EIupBbTHHswiMNY5FlhRhNxbo9tKv42KMbCEVD
St48Sr0lvomhIoo29PXzJ6XzeFBc/buu35oBUQX86HWBXTW2INQ2F387xcXlhgem
1juY/Tf4FZmJa9gqX5HoBRrlaI7MTRH7senSypXEN1hNS/U5+hKoL6xNsm7f++m9
LLNUy+PWkTDFNcMkSVnwaKdnIIFA49eGYCZLwQcIaVXycadCvCTHxrIiQieJJBJA
2of7JPKmyR/WWyab4KQ9EY9ACDJFSaA7kT1EnUfTFCi8Nl3bNvZQxyKz9mvvMZuo
4ia62S1vQ/PqHDbfjk7hZ3JJ7FMME9CO8yOlPhyNJtitiZBN412Iz/FsvzJcmrgY
11SBYAyI/z+6tZl0gbzoSoIDOb+fczAFbMBLAlVpNnk5ljIA5zwXJHvqfjfQwGx+
sUB45J10LzONUzvdTQ8WE0x9FeG9klDY4Am+JuCARPu/97jX1yPHQMO09OyPg0Sm
iuYWdJ7rqN6whHjGu423nwWn1Q4RXlO7crplTYOftg4BMMHb6zFe7IYUvw7w4boF
7GAj4TyJOZQ6CKQfve0TuA0pgl9N2rr/jlvOcRrGFGaJEPNCYrj3WCANJuxdop9T
GkAsRVal+tYa9UHnb2EYrAnmRKAdU5acOPrNaaFLULYijQpV136VdpTrQcLYYslv
ut9szi16KO3oQ00UsA5pgeB5yxdLlB6vi7YJtiVL31u/XemSnuuLQ6zo+x4UsAVE
gSfKmDspHZ7NrDjaGfX0F19LP3v3aXEo54aRDRYkMJkYwQAJZtxLWT1HzD1xhuct
Ev738edunc0x8rQ2z0eObHs03zUZALQBFQ9JDe8Ot736yj2CzsGmm4Q8izxoQs7k
XRy7P4gs4pN6qbBeVjFF/w7V692aACo5Kc1dlXsjr0HGXGTn/MHGLixift+skUdO
/P1DYIZfZKVTDyAzTiLIYcyLfr6u7fGD0+ea0/r2P/fCAk30MOgDNDCnHidEdLIE
bXpbjgIKPj9TMKxVva+aTIb+/7KtBM8Xh2ILMcy9tjx8grNVtQ7jttf7QK93k7hm
3SID4LgYjoI8Oy4kT6RpX91GXdC535c8RqmdnYHqreX61FpGOgnfGoiQyqPRvuMG
5flCorgqvE/ZccRlFWiEwqtsJVMdBU7uvAhQgzW0kMVDt3f/kHm1X6FrBIwnlEDN
f6ycFOmEbKle6v/F2fb6k1yxATFg9u9+7/jHhfXms2E9tzaY7t6dMMxJMOz6n3QT
Nx2qAEVLZz4e2v/Cw/utB0CUyXLNmmf1mlQTJQy5ZuO5f49P8yB2gzmdXcQlL8y8
RK/bGGYbZn3ov+nsPlFRd4Ntgcle0wdxrwLSH/F2fmjIWwUXL2c67+OqnIggrEXb
mZwIY15FZkvbcezNfG7+2v5WscMBv7HYzRi8cwccigvmLFCGWdLCYnfcwR20AHkU
pfGtNzZTsdJumXjJL8KIlVKY/jz62JhIo2wE/x2f4le3U1KpnHlNQuwkbuMlPkfV
fSkaM4HHtWgvEE0MLPv1bsA1WXF0p9e8XH1Sm+IwJCEW/5HXssfKtTxe0oaGSeZy
kINTIFzkZT4tHMTwrmaX4AL2vja5BWYCCEF+7PpF6O6f1EvHZ2iwuOoLEDZZFZim
5V7bAt1hiaIk9Rzne9+H1rkSiHLPkZ8qapPxJw2hSR+b6mAk9irTUHGEQhSRmeqM
atlQV6uCBo6eygwHsG+vYxRdIvGh8uNmoBUROCMagqeXmih0rwRwTf8HnRPGsJz8
BkhxKFugIEwhIALE0WCPWhTRtm8MxpQBcN/9gpwWAtNNiYNW+AIspUBvCCM2NY6u
uQhqieYfgtjiMjKqCnQESQcvCzNQKQWhOhzqRP1dpXLY8HdbvP+Grt3vnpvVnPlF
F17T2JueRYcazw1ysLenpoiiemob27NFjMnR1wOWgrODw8SyHZdKzSOeYhKTAvsy
U6KX+0fXRS+HDEBmwAAmQ5dQNYhKdeq7KMvREwwVl1nlv9WKWjPbqnrg0w8oW++M
WgbAWbpKVf1u1e3IRKPtAr9sAj3RYTTc3zbFPXOLidLQS/2KTr+JuEQvqwOTayAr
6Gq7gQhUcXo7h78HyLeSDsNt2FGmAwlqJphf6J9kxrusFyyb3QL0j8+Rmj3HRsNY
aIFkC35an/uYwPeOKYumtzTjH0lGHoDjOmA5Bn7vdNvCTgupq4RVjx3SVDkVRbZ+
DKnvZGsra4cXLPctyxnU3W731Q5N3qMkG67XiMUdqyIYGeQ4+krcS08lLb4KzetK
ZhTE6BcRedQkd1vReOQIGP7ktlXMFfOw7w6UhnhlK9Yyab44Zn/AB+qhcMHW1gPM
iawiaYfbREr9DLusYKTxRynli3JnYtRdhsgY4MuXzRXlJYpVJ1E9G8G/v3NNb5/f
8CrfppO12ZAnDe6jrgtmF/KcyaWYxiyiVat+5hUKhryjwTYzElJ0owkMKDbXsDI5
E0hzBYU3IzoX1kuWOrHvyB1n+RGlwOyE4eKod3eVy5gKYQy+8oPWfSbGIKth6mCi
0of0F/YKxshaNo1ViDc8pc5U+ux6DcdTBuP++9xKDaTwQZFK5ukIalb+eIN8BGeA
EO6g63KZRUykOQIWPfii59zuWWEdPUi+SD9HJLtKvO6cUnxATMZd250E2qtvPQug
jLQSudWZHBMWcViPdpkC2DV0vHyJ98t1gqcbQWz2U/gZUWmDz/w2HZ7Z/YcJi/A6
Wb5XV6LZbqvc7nVu2MOrv5nXQFPgS+wXOGHG58vx0CwPfTHmBnQu9F3dFv2RHuTG
kk8/FU2naeAsEeohCnrGI9rVBrNQfF+pdYVSoG4GXBZxF9JkWmrughtk6jnSJqx1
tc2XgmSKUFB5VZ/QvoMqWMwlAsL3KtFSgkQcfH1xVnd9aig2sMBHssNhMpAmUmBx
DG1FM2wTDbPkZSSeOG3CPDPQe4laDnADmbU1YTIgGu+S9HnQbpEZucoi3CaMK9S+
iJ/wH0PcKKHESX8Tp+kJXjYwkTu60YrUi1AYqf8i/2mdzlKSw1oCHS3rOsqvga67
i0b8bFvtnFksuMa0u1xgi4u3GDryGEQTqSbBCi16r5dBjiLb+jK9VYmo59N1dDhE
OUFuBUmQJvAKotXvcgiTLpx9xAI5Ylsp8tTDci4bWlB7CxPHBedFJME5x4CGndfM
wGjB6vGaTHsy8SRb13vfkMbjbDvm5u8KCpDCipVWvKfyOUeg6mqeoRdSsqC/D6YL
2dg03azPWHR2G6KjZRpBE8P9WqJBGnTf0b6X5Z9YVCDLtiT5N0UAMlfKufTS8T/3
MLK1p/r1mHHZsdQZ7fVyFbw+EsdDy2kPShadBDEhluMqvfY0lYYggWkCCLtKKy/E
QHt3HXZo/56oj5G96biE7PsidXJArfFyzxe3ASjpPSIIBjuq0kbpwiVSNk918hcs
KGMGXKwQZj6QUXdaHyt4m2bRAv0Gt3WLuYQIvTQamh31C09xIC0q4u/htO8rNeOW
IUrjYW5Crwl+Fj6BRAFTQlCwZ+5gfgixlBrQPs2GO65M/XFtsVujZaesHu2eh+3P
U91P1iOlousytBBMWHymNsgKB2Qzf6OJcXr76Ob9QY8/j26yJsxOX5O7iy3tKEoE
VIoJUJNCtVk00GAAeZhKg8n+cvq2BB6vXTo+L5ncQziNoBk2NMmIupLYGr4xAk/D
+MsapzdRA0LwiNNSffgx0ddEoMGOwIFxQ68UOfkpiV3/WcD5Nb0Vh60bIdyCs9tX
m9kIx72ZwZlR2YWiZz8PNXgp1ie83qT8OtKmmVrnLkMnDAVHEzYOG5s9DLthW0X+
dro03GWTo6qonJcHHqDtnt87HmrNZP+LPzU5cfvOybgvaUbEpvl0tRw8r4Y6HE8Q
9MB9oIwNLk3aXYelAzhsueA9ExPSX6/2xUmCN5PnwzbcfZao7uK2Y6j2xDKqFRwq
IRek3NwEHE4xGn/ML3IMcJMmkbKFFIrePLKTXJrmJdMRTw9e2hGVlxer9Zca60H3
EjscKXIp++ZlNCOj//cDNs0BOUAKjmHBouZmLQBnYBqf3XhJ/oUdCG459Ir25fl+
EqV1ZIjc2t1slk2dfn8Uaap1jBsYL4Jbfqn5Q8aytQqxhg1dSr+x9evV8prxFmLA
C61A7B9duzEn7jCGuI6sxGMsozeyjC8ySU2wtPZRqD/vt28lFrHTB/TbQvSTiaFF
A563ho91PP0iKKQyXix8/9oFURBG2XpjhL0ikM0q7Gt5R/b/20PPtH2SEroJINYK
/TiinRYv/n7XP8FI8iCKi/vFLVpHSpdRn/CSKCh32T4oPA0C94lOkyoeFf7x4LKM
mhthMjo58eoC81J0V23OnALx6THTnJooWVQNtffl/dnRUJ9YArd/hA+mzEjVmKJn
GQlW6SIyvpZQ41W2JYGiSAcuPNjpoE2/b4F+aWlzJR5OtlU6o8hISXHlCOmeEHDa
1CsMf20FhExY4MBPjbX9vKTrx1OE210FwUP93+H6oVuXcD4YsS2TFuUJ92khX/p+
RGWkWk+hfmKGKYFFPViuEPhWbnvvxqY7l4k/pkv/DkW0mzyL38IJxGu4XMi9dZWN
fi2OkuZLAiYUTNa5mMJIAHwEHHNr20/m4D0/e+ZGbB9fnaq/m9dfduxWaX9oZEbZ
GFsyh2hiJhKpci4EnF/CwFUPB+wLhCYuokBZAfVeq3SH7f65KB+HkBI+BeSBGbqE
UKqrkKTrnT/YgfXpTO6ZQ6Q5qq5HiU+vOJE/QK5QOvyDLmp1B3Ik1h4pfBBN8PAq
XjfLEmtrqJO7RDxPxRCY/DJtvYTFRqMsVZ2P45vjJl1a7/3DFADuRR5IZWhY9c9Y
sugX/Owd4FM5kj55vtRQygPrwDVC9nngow5w+QJFEQm2hVbMO5Is1hMEZnWB0AQb
FUyvs3hfBgS4lIySjxehEx9AsLuxrOyVxLouOgEfMiGUXPFtzJ7sUdZqgvJ07pzz
cu7ZV4b3I60BZbY4CqXvHYvJmIE+Aq40Qqe1Ci2Q5cl5JG0tdW0qo80LcJXEtSf2
lQFf7iL+fnuf2JDNnDfaNHW7bj/GcDkx+UShcim2hOQGuKQ+YTKrg29/52WsITKG
uyB1qMoQdjJ1Ev5ZDMrTSFO2ocRouQh33HxLwGm/dGQkLZMRJtCZ+UrUjePsXy2B
+cYnRs5oIJfAz5RACmQlrN+GuqxTJSQ2Khzuite4gQIdLrYsBAjkYaDkH/ty0QwT
bdHezWwZNWrylqh9q0yLybHzmXGxAunmSrY0tQ5WquYr76mLw7n/vo1z6uZJFJTq
zIigMeGiEY2NYrTa5skEwfq+NSZPN+Whkb7VGj5a/rtsMtiqSuo0hbWTeqN8ryhD
YhqDRil5osuS8XcSXMvBhXPHBHCbCqCdMpdRwztTdEZMFB7/9qQpy6NQe5TzT0/j
Wnl8YWSnn+KszgSpGDQbZ8EoBu60Cp/FDRQf93uVg93hI0c/WyG0C3KeUuWJVQm7
boesb2M4pPDfj/CvG1sFaKUEgAMBzvCmzt8gwvxT9BVRfQbEwXOS2d8k6cecBV4D
0JosYkcJFNS7aWSy5LHuVzzWZ3OImSWxmUSROcIWf9SKizb8iL1vKkOIpgRnwoJ5
oabEi8577HCokYN1MhuF01HZkKgo+bfptWEJ/vF0pZvVgDczNhffQvbZLFwctYya
Ng/d6LdhLzLqJnTeHSHo1casJUk3H8A2grHXyWPOBzkbRTKz9gPXtLQEaJFypDfq
HMbeZtTEnHrrUiKtMO0v4ezb6UzW8lp1HjTfDPlsD+A0I5hwc0gwCRRCLxfGRB9W
Hs9zEYVsR9vC+PEzBYvm/JQnT/dMzYWkPdWovbHsoNF9feJGsRxXuRhM8z69WHxM
y+jaBDdb6lIXe1TCTl/vZyfl8MFg2t8Jtc6sHsc9c9VOZzsLug3wAnSPYGomUle4
ZARwoMYd6wkvCgwscaVm9hWdXZnmyHSUQZw5uiDT2MvvogjBjU7O4U8sDi2I0Q7W
WYANoFgRchs3lNIGsA3vOwQcpVF7X22rSrWDTRQelpq9JvT851VrGHWBxkV1L/9l
wjjxluYv5MES68jbPPItrjLAtzgPh27L2xflR7KtrAUB/qWXB/B46KFFgnhpFwn7
lpGVAHljXydxK9DzLUVDkGddKMydckJsW+mrJk7yZaOSPz4NaUWO7N2fiV8ggEjN
CwQuy73tVYKR26jIfiHZV8wE2h0d71by1IiBquFKou6fuL7ndEcJfMLv/pdoe+0A
OxTvAmLpeaXpCw5eNVl/7YelF745qV1THrKnNVqNXIEUXTp4JxRrDZ7Gd63OKesd
jwg4Gk0mX76xBaYxccEuJOVuYoY6fSk+MU/xbmTtxY6/RMIYeF309xm/MuDg3R/7
qPX1rjFrfo/XDK9jueoQzqSpBmvE2Q300KDRzRwDDqHbW/vvKToPKhBd4r0YadGA
Eu9cwIPI4LPYr73rw31u0KBWO9toe3HKHJ5QA1WSsjvRmSNJTqJicLcsa5i4SfQa
5FNJ/SPTmZe5bLgbRLPkdZqSNsC4ELL1X6S9EBdjLGgWGvnkvKEn996Kc1QK8X6j
c20wUz7JuF3IE4FxYzBG2sWGybAYL5BREVXcL+vqN9t0E+m/oao+2vJusM350KCo
BstFDl3WKOj0YkhDVTdAB4FT/P4lhY1W340oyF4A90swYztmYWa4LcEm5BfiiDTs
eb7fuCbt+7FqEl/93q9WRepiEjMG/lqnG0xJExAQ2gR/uui+bumuBsmTIrUt1YTC
qsdO6ynIw59hV2yc42tB1NFvgYMVec6+5FAdX1AkaYmHY5589N/Jza7ayr9IGk8k
xYc+30oOxmaebdx2Bsl0GdLEke5KUSr16RJxoRJsawBbotAhgJ9bryT432h13NPi
tDOlQPdevIrkyvpLzvxRgjOjeT21AMc2X/+MnGhcmxn2BHN2pQfCV+uIBzs086mp
Oxdk5pl48MqPpMfdenCQqS2ZGarlkOV4kk3TvnMiLd31CFzEAJ+DNwyNAlBEXsc7
Gyv9XwE3WsKuCr3L+RxFZ5LJWRjen/fbqXW5H3ONSvsx/1h50lil7aUsJ+lFqjpb
7gGrMAuazsBmTqLbuFcGV4QKJ0hPQ+e3b/WzU313E3C6uvHGBM1ubKzajs8Ql8i9
ru0tLOct2r5ouuqPOBfscm/NvxlnCIKr/rP/dYQ0QLn+Bxyh6aFSWX4IA/Ft/XkG
NSCidRs7E+lrYyh7od272+HckIaEl/SUV92C/TLjQy5IJX0+gk3E9yg2BiCP8ACG
hHH/PdmxYKR62YbLQD7LwOmC2D89w7ErrgkaSUAgjDiTQR0iOBV2uLl8S5ACkP2X
JjtMZxYzsjtGKm+ldp0/+AQizPNBHnpC9cls3H7eEDzeoQC6Kwyr97eHbsluYjGj
XfVxEn/E4uV2AARqI9KuZB1jyihS45MEg/nWkXGHizvex1rxHPijdoWQi19XBcER
SBxOnGUHpv8vlGD+3s0y4OEm6BqSpxdRcN/ZCHq5Pi/1MSfRfVMEQ7ZWlK7J42hC
dBUnu0OD9zcmCv+bK0bFWr84DwGsabtBlsyJ9ztRhTK5GQsZh7xUKiW/flyEzPuz
b4sYQ8lX93o479Kyh7o7K8MiKxweAzPygf4m4p79Yxe8hbzOpFOEcWDm+Y4dmBPB
bMk7Lba0e3l7hGNm5EdyTA09OYJjSWuM4IRSUNqQC/ujirCIJuX9Mfm1KF3CMJky
XGOj1prqoFQxDwS5N9jdpHq2BIBG9ixAnLztZofREgTXz/M+AVvpSX38xeB42FEi
ApKoK55+omnguxzBRvdZrSt2NJ8cj0mI93BkK6pEuOzcJVOeEOJT5wlK9i+C3qM3
60TIiKbd/Wcm1gOGoJOodN+cVHlySEYDUq69aTIWU02c4xjWNuZKow8LrSX8Uq/M
9Yu5vhVPmYi6Ed0sLbpK1Fq5R5FsXag+lZTlLDz8mg27JcBDvaA3EXUl4E4uEwHm
FUz2+BZk2as88BazitVx4oOpM0dMILa3SORKEM/uap+L00F+Har3GfQVJoY4FBPZ
jz59FNEQTuVdUe8U1jCXPo1/BFm7Tf1dcAkBhSgipSwZt5RbDivBqe/I9pNXyPTt
kSYzkc0c45RjGugH4ZJGkaH5l6WW2ALriFpCNjxHja5mSZGHMZMQLST6UU44NIS5
IXbW2kCaBbEnJ4CBe2XTGdXV1PUZFZvTYt8eZ4Peziq6ERyZlPuUEbqmFH/W5SOr
WuaoBvX7AP8VCEN1bw0f8ADvnsDRiT9W9CsJlRbZJbxrum7B4C8f100NHw3GLmPI
WQsWcvV7DkrbEEb9TwO46fc0q2Sl1Q2pZGwDo14B4HHdt4OXi+Z7qUMfc6/ArQtW
tWQZsGvt0PLHSQqBYd8xsTW4YGFI6GVJbjrbtnhU9geBWovJZL5PN4tpXr34hnQe
tyV40MwYz7Jpn8tooSiQhMz8+6OEc3HHZf5HCsEpF/QE0T3DD8Iy1F9v+boTCoSF
VFBjQQJ+uMilAV1H37s0zG6ytThT7FYSYGjDUwouJ00jwKkfLYy6DCuTvDhAW80T
IBdx63p0a09zLUgdMsovIXgJtTret8IxLCmW3MdQc7vme8xNULwJn5rfp8DW4/hF
OhOQzYygBm1cKZ/GiDJiJ0Fcu0ThuxFAJGtY0hxTdjDyYg8/u5PYo2gL7PkjYV9v
Y6pgYQyl+WWiOwNc05RRpjH8nLbJw4lPhpzhO5DoFqL0J+RmH0MUJ4BNxDUEP2Dj
ODEDenTwKDpK+W8APUjDgz0BNopv8yPVzBVH3ds2iss2Kw0T4rPiuFNYAtbL1Wrh
fWnevvhex20FsTU8Zm5MGkMgfK/OJ3mveolbYF2x3YhTFEK5VgMxmG5J5qXEhSNJ
VRRwfOr7RPjawrykqkailbOKJ0LZR+gL9/AEoUVq9LCgmT1L8pw6sduhegdNAaAf
sR6AZ3rba073QAWhZjkWyWEFn4iHypF9frFFL4W8wOZerBEjmXF2Y0h3bEuY37UK
LiROoxCNYz2D+5LJpXII71KFlx/qe8Z+uri9tG6/76z9cgCUe8Slm0Z6UTTCL7Bu
3T4UxP/i34/qk7HEEUoH4A2xwcMWJnCfdnd1B6x+UCJ5ej2nVledSire0UkuwIS0
I1W01KzO5i9vt3ZnPeLHYtwwQD5xzKIVnZreBu4VpWTs0kY4VjItrcwHq02X66xm
FQYlFlUXN+i49KrO1wwKnUqWvdQcRi8OEuGvst9KNfMb6IT9PBjCb7Mp/G0xdQYz
JkUUfW5R+WHJVQzkoWea47wN6uLvLC4npWRnJi4WkC1HwYf0HEtuF/Hb4j4USnjA
kNF1h1bYA28O6Cak+450GRTe/PP1Rdw8Xaa0dtI4uNC8DMsErQHRCb5WSZIfJBrD
tcWKQO7BUl5EZ4h85FS2BZoblUv0l+cC86jSI/LUbRBAMJ9L4Qq9SW4QSzug9svD
vYuJFUtliJiufbjfMliQgYWG80iLD2zUxzSC+S4jEIQfHZgNMhQWRba4gDxxmgjz
PqVFgQ8A/TDzgPLu+6NQGpOjoaVqnM3e7QfgHxOn/ovGIhCwAX4TNb1VTR+7a2xL
1TPyDVMQ72cXaiiAUw7uPqQBe2sV4Avofx5Gp4HkdfZMVpbSrWayG+I/Zz0R8QFo
OqXSmtUrEZB/yfy7GqG4aSjIvsP3TjGVZyuyVK78nqXDrM1Ey9Xh+yyKX+T/eGf4
cHhQQrO2StAwmFHXOZyu2z8oJ87MQrFO2UYVoy0RIM48FoSvXNITBe15VmI+ziq5
k8aaPG7Cys8/ob3HTKEsOL6RAxTaf3nhddKwYaa4DBcsEVvmFrn9zrswJhGhkrHt
oC58pIMM36JpIVSw3oREv8B5LEIqHqCv8qglTae1kc3jtrZsbDXhHBrEfJj7C9Sc
Ey5JKeH/i1NLnv9P6FetxkRnR7+j1O+oa3IG8aDOaydQc7Bt5MrnUNIcxmH0Js31
7nBgPUq/T76izN5rxWNzGLTBo9wgo4QyQspNRUctZfosQ83LexJIHzIlXetuUVcb
dnOzlCflyQwiN3XgDWy4sBwIZFtKdU+9Ey/pN1FTYSnUy0GKpG0tF1Qt4L+Z4Hx8
bQk1AIudNDa+QIMyCUexXJDNSX2cac3CHPNQwTWAbBIQRLjfGRmm8sVc2F3cYHwL
ZtQkoO4GwPNsqetBlzCTX6hnZIp6wcVCx8BIXTwf3NZrK1pc0QxGjBT6hqpd3Bzf
dyLU0O4NwpyuvtrDbzi9zojACiUPuD2ZPz0X34TZIom9Mg7N6NjVKxQfREfPrtHE
vvEUS7xjVlv/B5y4VXDxonJKJoRBTKzFn8E+uvbfFwkvdi6/T6/Xyis09l34cs/G
n+a1crRoNW21OeZ5j+eDiYrZWzo/hN8vVbWMCcvnWxuE5aR7h0VX90wIxv+z61p8
4P1Ow9i/6EBZ/BfRPRlmtQugdizxQSOGtY+qR0LyWWOHU31S7rf0YvzCwKEiETOo
4OblH2Q0Xpk1ZUxgXnBHWAX3KS+zRrj0QYyjntHn4R76An6vYl9kS+tI3DyaY5zD
z+aA9sIqLtOwRSgh13xGS2rJp8iCfnENLV5SRMuqzHqO2Bo6ZtlrMF95RfSsLj7T
UY5RlOl30edKHMt6i1eA0bVBBX+5csGOMCjCqN+I8fZXXMEYhiF1un2q66sZagNb
NQ4hur3YJA9IhmMpUOXecjP0szkVvCAzcAgb8KiFNMDNPQUz1lQDUuyqQPkLXCjX
M1ESKJux7Hk/tUuxp97DTcYCj+WrjQ6lIV6p2XRc3RXletRbRUzoAb3684HUVo0i
Fu228BkZlvveQLwwKm9TsVX8vOLIpvcgSBzRC5q87NIxyCvNwC6waiBG6AAkS3+m
+cVe9nzg/fo/E99cW1oqD/fXNRGiRjgNitIGUW1U1OFUK759c3U7idsAeXFzSL/B
eO4lCbduv6asvi89oWGQ+MP3QeRd1OEzLUe+GCRSEV1HesLTeDT7EQH98Zwxpou5
AQJsIYXJsVU0u/Oh8w9oFXiyzbT7FKQYduEHxtKhNJ90HA61fNnoweuOesOcz2ub
aC4RhK1zdutp7ALHpQKvYMO0id86ImM9I6h4Wu8RZNKoBm3xSNVbioOcrGZ6BGdR
y2jDNRcGd/npPr2E+31i3PnEfybLX6XhDETMlgZrAL7Ef6KhMFv913U2aSASnDui
ZXRbvkuGoXnJL/y72jMtWmYBJymOkqWnQWk7Q1Aw/ljRIDdYPoW0gGwAU/QAKjLc
PW6uXD4FAVmVJvZY9lM87unFLZFNxNJLw3pbWlZAuwnO6nNiiBaORNaPi3kObX6y
C6/rHPLbjQotdg48N4LQ/9MzSu8HdKs/tk40dwjUrPIgaGqDgJjz1AnflQM14h71
xzS+tSvIYRgSdHGkU0ecc1cvnAGub8P3riGNC8tW0odw8o+jU0fH8pxseOVKu4dQ
bMAPKixIr7hYp5wZ7TzNnXCud047LZtz2DXzYwi3AqL7HhWYf39ojwI1e7QP5z23
40AeFCumISpWyo/DnN9Y3+3GjXArYByUpFLoHbygdz+6FnZxgdPN+jDVM2Qe8toX
YrFrIIdWG0u3Uh16tXFa5sy8G2uXo9XOLTmO9gzlcQJAOFLH6DWYmy8FK/yQVzmI
Ofktxj4Tvr4U9OO/93npLJbrFSzQ2DY4BNy4HIPgnENsUVcNWPKRzVnA2UPczX7g
BLnlmkMVdty7hqbNeoZV220K3fhuDcNW9fy2XlKsqmtLNhuaKIpXG/nq7VuYGqyc
CcmDSGfGNM+R2jIby0dSpwp6VVeVN7MlPnlKuU1nTauBH+eJiDfXOpUm+2oLvmhR
XZCdj+4/NGwWfUVnebUS350LOdTdffSCOzN2cTl1UA8G/Mdxm5xIqcKzh/qQH9oy
i+Wk2X8vrFemQBgoSwt7oA7eW58ROHatvshT7YHql79TrAUnEjC2DguW6DVEfmPu
hR7BrCp0vn/rqy241YDd1GksT9Uns3AWpp7QIJDZEs3o+7ay7Ev2dqCumcg+Z6Pm
ijnfSv3NMlmSr566ygntJfwFfDoWzfrIAnqNyz7/riFfuLbmbBngCM14RQMw00tI
xONNrFQC4djejpldfFuAw53XYK1Zg3Epjer4QSZLaYUsC0ViuqjYYXp7BVoVEPym
JiVMJv/89bhe6uMTFpqqwVFEQw9yKAkuJ701FXef313OdVKklj8SYpS29QeTgGMv
4OQCsUuwRq4iHDH3fmr4d+mjagpFVay1f7wDWr6Ev/FTUzVU6XN+Qfhl9cfVjJnI
whh3kDCXZvSP+er7ED3A2lXpOcLSP6IpSYWle8khVFylKr1Z8we12HS0njUgAPPU
NHYFKO05N+/NRN45UqAiiHaQm0QfBBuOE/f/FUHm8Crxhfu5DdZYh4zwPrzF5A1K
/XJ35QKfaAJirys+ZdMvt7G5yMO+utmhrjdC+I6Mi6r5GIPaBZEdiLVXTTBqkhnN
HZJadvnnV1HRWGVqO3jAsNsozuRLEb6gSDkm6/K/Awo+pByU3iVpSZA/FwCsQmy6
2IyoLAT7d95cihf1QUEFmZ71u4dGtUO8VlQJFRUPTNxi+S958lyj9BENRNAjLVfJ
YrLknHZK+YJugyhYscIZ/Z1UM1Bfee7Dimts0ckKSTrefU3UPReDSjshc0xo7bHf
CQroIOrLL1ebE6Cl8ZbnIRGZs1zN/5PCKrQqz1GpclRhT3AC8jzJiw7FpfxHSamN
U+K2HyzSen71rOGnGAj7vxYfv6hm3V7Q6yrtHccxQ8TZqSXbmFqt/AUCx30SXa2/
hZXix8W0xLIFeJtbcJ0jKBRsulb1oN3VYCek8nBLGibC71YVXj+59UgvvcTjl+34
j4rAQUcdBkaawsKbi6hJLEFJ/Gt6Y9z/SCcLpD4k1aQPM/ig5ZDNkj0aOSPwYVaG
obUng39iRAZPs4HWHbJ+OMmsL1pm2dXwAHG10gRKFx7FFBTTMo5EsMwW9NHC31ma
rFNlvqDCltturTUD69+JF8N9BO/lxjIOkBbNvcvHUFi/onHdznZOzKJDJjnQMkEy
C8oNfLgoiwAKNjjJgKdQL++UchM7/bf1tOigYtSVNayQU8rNOiq7AnP3HyKhflF3
KANG6yTDHWGcxQW80Rl32C784FNmdU3T70vW0rIPr21B5op2HaJIGy/FkI0BNm42
xfMho7TPJGR0/9li4KJdOT4M9RCK5vkSCHS9eILxP23dgFMkH5CgaBpYW2fvku4n
EAJXrfdGMxv2KKahzyRvIZSHuV07cwPNbruwa51PP34BNxKBQvW4f6f+XFISvyg0
VkfqWkvYsDw0nmmpID8yDeo1djK06oEQhWD5oXwWuxcCGcpTQvwRcgiIV8cJEJdf
KtqamnS9Yoxp3iHjdUouCxb67vmcCXzjp0HkLF8Go1iaDNzCqqu9JrCL94kyCSE2
1XWGtM00VPHjUJ3Cxt4DN10aOYxSq1yZcXRsg7Pdlt1JN6lAItp4YB762AXb004y
NqSOb6ihhnL4k6QokMv1ArhI1vEvNBjhrcjW+OST0ugUY7g/VO9TuM+jckf5TOz3
0xo9XX1wC/27bJmy47nFjhCtGyC3C8OMSuFvGp1FEm0MsvBT51iTmtCQKI8LRlmi
iEMs0RhxMupMU56jpMvQWB9CbjKyU/StFXfXERckxnFEwE17+u3N1tM7SGUf3j2r
OKbqUVW+RB2j+0pOgH58vASW5R4y75BKaeXtqav07fZFrWuaQNi352fGRbUKclzs
vSKTLkavRYGY2BD5FRhjhfwhfR9/v5OkhzEB1o5WZ2fDR1/024Aq7f/HucnYW971
YEMyE6rOSB2nr0s1uyHWnbhH8zmjDzjqdnBUicEqkYLSEkl8W4Vjbd+Jr/6nsCtr
s/Z+dzPmv3Zh//gUqwljzP2YnOCm3SteShXOHr3751plven4gymtxbDvVm6+HRHj
67Fl2DQJLbVHmFq28TLU9re0sVHgaMufqwso6dAR6t0kfYz1xzeQJSheBqYVEq9C
TAzhtIlh7fp/MkwU6jmthzXuWTfbsq5mRKs0xlAk9T8nVDD0TH4CQrY3O0BsH971
UWZg+L3l83876+KpTOFGM+viGkeWrS0hqXe82g0bt/vEGegUYW+oLnkUb2rIFUiL
hClLcn8qN2bPN2u7Jb5VV1roBirNAxjeXZZJ7du4tLn9P8j8mOuL+3Il5ox2wn0h
xdRIrNcoSREBwXWMLygJyBY+W/VPS84vPezG1+94GAt0IAub5VkuyuQwQCyHsI5K
wmVysewyT890zuJaUmavqAOG6Q2iPR79VW+6oOqSSAPd9cWlu2iqe0AZRVYOvCEl
VzT1odyLZdWRGIk20td/tXYN6idJVR+Du7D7uid7Qid4dkL2hvU5lGde0gzH3j/r
ZUWHBoTQMrmCUevmpBTgvM14und/lGsNgNO8yxPAvLMrGRbfrA/Jb6UQ8He0EJX/
i5jG44JgTeXFGoOgmQE4yJuqf+AgmmhvLlWCo9hzH+siixIyVvuFoP2jsV0k4ChO
9DuEN0KnpimWC+BMiCXblF+7U8dXxK/3g0KhJ22qc7nOcDrQ+v+e2NpA4CVz5Xxo
7idcPLY1a/w5f/jdilqS+AC3YJs/+v94TcHgY73kSotGzqQWt/TdycU5GLUrJbcm
rujV0f3SZJbbx/2R8HEILOi4qxqGjKKIJ4Z191ZxLA8gDD73TmoGHhcD+hSykRB3
JxA1JmevmsY7eK9DXlVwFVdhb+3H7bSR3DKSlNHn4Yds5LofpPRruzM5S0xam5ka
O0EV3tmrYb2XmvekhwNVxy46XByyXuLC2FWCtTRQRoC2G+xYftBGXZsWX4mDYIVG
f6HJTrgV0Wj3D8aLORa/vs/T17bgO59HBEWmNh5U0ZDiWKsWlZpTshGVbRMLEwNk
vAp1qOWtkR3WyX0XhAKmv0L1tb9gKFWQtOKBStpNDSFDr+XR0K5WE3FWxTWK2Y5A
xl/Vf8N5LaAyJCNvPPfZekqIdzM7TaVEO/Taug1MxV8FqzzFUFI54rLYanP/sj+I
0mNTvAnxAkeBNTL0RFnUMCgZ44WiAv9CEqmuIhTlJY+7p0vFywBadnXjXLPbvYc/
NecK/pljSDognF9xvTxbA2Or4RYIpIy82wOsxNeNvYwD97HPHVc+k7llmjQCbMDB
DFjjdEkCvy621/oZJ+FcfXw6YJKcsK0dXq8Wp/sueXcl6LnV4fDhgx7gkum/UbP7
dYh1uQBe7fjJxVG1zTXsB6UUNcQwAjUyxUhvAZgsfiUPnQFQIa51XkD5QE1tpvTq
XfmstO5t6j3/S5iAsXjFCQraia73XGgtL1AZ2ns9snIsYm+hL/EQMYRk/lkK3n2v
KQ2j+HY30LIoTTXyPvAC/NeGH2rwGYbnu0lo6mYSKhbdBoCr8TGqtRUKLknL7mHQ
jjZRKhirgnfZA0HwftrmghpIXJ6Tw/JoUiPCPrN0k1uXUR4iLkOdHOtqTJNyCtpL
v2zLpQJAKzr0ivgDlKmMQPTReE11y2AIavmcl82bPQbA4SwIrg9wdOfbLjpBLucO
Ih7usEnqZaX4g73OWjF4nhZ/LljiQ/TneqTJqChiIF919L6gw17RPllj/rJ1um64
uZgTKVFJqpqsuxRM+CgZklx+lOws9PXJg6UStQMrR2jERWrMY5D8/sQFJldmBfsI
JuXkWAUMbmyCWxStz7P9oA1Oq8LcgQd5fEEVcVT9Im8gWCdBPrZREy6R4xxRHiud
fGv4rjCqKs+rJn+pD8b2WZHf06WgGSU+XRQoMnoMO7cOOVArWsswL2knoEigUZTA
+8Vvuf4ukUsJfcIjtrgKm1TU1WczjbRThlmKfTfGgV3tJTMfQmV4blbTr03zu0iX
JG1r5Pysx2Yri56jp7ZK/cwW7HTVGA+vgYdiA47duJ1JzyYYfrQeH5VuSTQPy+8Y
KG2wXYcrYRpHtf+W4tWAqzB9SOW4Z6ITxiC9zL3i4JBkLY3bIB3MVMmbMQVIOub5
wUwH8e0ca59M8hy6zwHprOgaLccTlVoPRkWZWpKuCY8fJZzCO0WWZUelBLpuD8nA
EcnHjjE1Yo75nDk7LPlGXqb5LoFgmnDIOu1U/7iKtKGY1vSlsLodS0zPEwyueYM0
iCE1kSrZpcw6fN8AODbFSgj9bUJxCpnRJBmzcSPQ9l36Vw4LSAjDZyM3yIBhlqSN
aUX5NpM7OjJ+dCQvVEkejdlOnUp5GP4vLkoejDk2QGLuC7WMZ9ksPeLoFyObTFZ0
lQTmeZxAjXCOQwWkYFFFaJ3Fa+O0cPWrYlpH+8J5EI74XvsZcCrug/ZGdh9upa5x
S7lM+51FgQ+jOLV8vJ4yNcAvhBU80drfr5cXUB7WixZnRmStpJGDQiYmwKQCUr9i
07hvdVIpMGLdGr1zv78w2CYagRtDbSpnBjkJ9VtbliAfO/ZnT6MSikQcBaqins96
KuzfPeCEEZdt7HjqMvBYjQvXzxaAol/lE1VG6MvXToOmj4ZRxMTtzxFso78FIl7J
c7VXn5CNx8x/BCQO407X81iKXwglR8ZLW5ESXXHXmUT6Xj4xpF5D2thHBwVpo2dx
pXEuLWasy08QclezJidEU5/o/06YOXcoiOqMKqYBrwj3zSc18lrKFitbCZv+Mjjc
hhBVdQ/clQx5KlCI1K0Rmm8Fp6vnsCxXt9g1cWQMbTHt43NUXApNQpAZ/wR+vWTz
jbw6wzagKsL8VY+hPiDYvtGe0k9ovcxM6Jt9SMc3qYjyevx2Y9nuuDxNIuw1+nSC
Jc0l7hqd/sripn9J5FsQXpSy4qZ14Vdr26YxEer2S+asDB3mxwP19zvm7tBnzCqb
klHJfZ0Un6gRHmfXR0da/p8YYDyEOg2LJvDqztnWjqbnNBfRxwISMd8fBPG2hFG7
v9tP4BSHofiXjo1mxOwUgp2uHZVx+HLWSwH/qk/MMezSjUBQ8r2h4CXvL8IuR3Wb
wkgU7mue3H+gC+VfLIK8vOdGzJLs+T+ezyLRfoYmvUFB1iYl7HH6PE2nBmuq3OwO
ix10Y0Cg4xW4uEpk4W3lwXfGS0v9pMjGZoihNGYbuIau97oLuChnIH3itB7FMrGH
c/9/kFNBIAB1yuoAMNH1j/OslNYVVRWPpsUPrdgivrrhm7W3IQdeCDqguKzpNvSy
ZPFFnwIBhleHIGJoOkx16s1qywPLabhGuHafj+ruRBWSu6FD0cz4kEYCG5k+Wa9k
pZbzuBCxDs41N8XBuUtuJ26f47dnrb9/91iWxHUEinMz6WulfkGKmWe5YkfCjzav
WCJ2rYLbRWvnRiUP0n/tX4ALaMpF1r1s2kO3f1ZvQSU1UGrDosgVK0f189e5T7en
60Xliob9iKGLVySVGskUS06NHflD0XOm/Q6WpP5ATFNM6XV411hQ0uQI6HlcxT7y
wuFP79zV5SWqBa4PPR47ZbmWLn3FCiVF99IIUHH9SNxGSpJ0cs77pKaFu9yhQ/4j
ISBD85oWUDi1gp2+Tjwiof0qRoRuEjhP3l7ZqiYkHAW6ZfxE2bB4R0D1kmVQYcUa
gN7G2v2gcbkMDKUNzzcj6kgHvA9tFU4BLnfrcnW80ZF9Dt0bdCSX/JJq8X9lGI3b
jahA/A3v8zVjjF9TIV4RYWrW5FR3TXA4sAZN0JS1r73sINbggaRxkhlPqH3gccjq
WiRvSpN3zrEOxn5Bcei5TaIQtcQtHDzbpb44QlsA5iRg07PSYasERXemM0un2t/R
0oF2w/8iRtvaSNYY1B3GioJsH5ddU4yV79zu64rv6X4o2nwIQ30VQpdPNe0954RP
EvKyaK37IaNWrvBidCnZIaCNojGtNSldl6A/T3NvfhyE5wq3Veaya14ds/JNBUKq
7Up4pr2vpVn0CddXN6AnN+OVhcXw66aXLeDhHJ5U5/ovaVJfJk/v8H2YVHZ0mUaY
qRZ54I/2+NRS6Qi9tPowV4MLFTfKUJu1p5U8fTHMPftJ3qvJvx3DMpgZTM4NVPgy
faZmAUMoxg+jP6om235pYUXh3vd+/BHzTfwZH0+oXRALgp0HYm6WEBofo65jvbHl
3JfP53fE4wyzKtMmpl7UGnQuAO/vaeYdc2v2grI7C5UOZ4QH0NT06jFQdO+B2CJc
AvR2G7CHce1cqMs1K3OpkFqkF/FcCgbDsczg95B8od4uZrXPe77gzcc9PufamXaM
v+GjITpkiM3UtxFfmOFprs0RUAgueKbWdBDdnLhEEoR2BKxAeZnk2sxr0ZF77UnD
q4Ec6jCU1q1Lg0ikZGm75AyMl/0kabsxvKC6ebhq2E4BKUhNxaX2SvCDFi5IGNKM
TIzC3kRAqPyvEnNKWUomz5XktKMGtw7iKrqc6ckXREpw1PhzOggMQgfJ7Bx6u9pI
YlCFUB4GI+M8eHBzEeubsK5un+Nz4HSz/1c3e6w433RjEbHbALdvfzJASIL6xZoH
cWLh1rjtySUzW2rDqXAacTxKVPZaKQORYB1ypid/7jXHkM2/KWVWW/m+1Yoq005z
w6HioURvJtC5ypeknHQoYGEL//QT5MpCvZJaWm1Zoz0NfkognExD1mzR0QzXjD5/
7uTlUY+ZfamPTmhjwKh9glT4QqJ59wzwnmfMfgHAIQvYbIA4i9jqy2S/BnV00lhN
dVIOXInEH0FhIpt5W4qoIPWHMByLVjfkDJQJOuWGRnuMiYFeWBxjIyIQVIsCo+5F
qb9zO9G3UE36tweL0zMLMV/2mXefj7HeDVMLJjrU/owqz/vN98yn1OdQGSDOXAAE
4CfahV64ECYiPIT7lT8/xINTYSN1cnYMDSKYCGNRsiElim2BxlmAqUstuvBih4GW
KRDHYYeJnOWiuiGc3WpRn89afgnpdbzO1eaHsulu4mtCy3hq1hfVQdC96Xbl7rTx
sDkvii/5Km/ltfRJqwg8owwAjizuf05BCscxtt9fEYapYcdV+i33e+9iCAdli4oG
r5XOyeE3i0pCccCBMTdueiCqCGKEcsl619UaR2vvdmpQHTV41SLxg7E6BgLV3Bua
DpH0OE4SJ95+mVoFp7EQbs+ogQFyHvBI+5g7y6y9jHv8xEF/QHRQcLzHZJg/We8X
tb/S/bgBipZU15YlMWKlooyz2dP4nFgkeJ0Nz/dzS8d2RQULZR24tb93Kjn10SeC
A/FnQ0fJEJ2PKJwBKQP/x9AiMXX24DsFuYBfCASak0mHQ/Von/VqPhq8lA3L3itU
wOO0jBp5FySd0WfcaJLfU15TDm6vgc5blE+gm9cllOvN30vLBOoe9xOdWwAqiTWc
4gDHDZ+lo4f3z3D5MF0TYT7+Tl2dujCwrQbtMwBcLNxGTFTUJQEamjWvYnoFtXns
PhmA4mLm45WdcHA4EG513C5BkR0+c2GGHzcQsviHXx0SDEz0qZ7N4yGx7ltuv+Xq
klctPvgQuVm4nIVB8Mj7gx2rtmqqr74kkzgMuDlLqGTJB7S5eZBxVrOyLJFo2rUS
JmqUXQ/C+CzJiIoSH1YP7UiOoXBUj8+6we/ajblpBHmtSyEavHumfaPgpwfoPE75
E2ldSACnTbBniKZQNzgKDZz3GISrtxcbOZwlH9K1Mi2ERlZ+dvMMZVWvu7ww3OEe
V+y5/+mjjqAU0XO0kpMB9+uuL8H0MsTYSRS+/82oTS2yEDX9FWjTNMolIWNaFhRe
vE2dzSgkrcutpIU70SEIzcoD2EtithuqautHHwL0FspdlYIF6KkvlgFiUuK8GVgs
/bSQrzUPLVvIhDa9ThYX5Ifue5dAZf5vadGbORlipqZg+omQEhEpPfoXv/NVxU7F
kLGS+H4XmX9drny6E/WJOZiU2mmWhNcd7Cwt01WmvjDla6sO/c1aoGcUJ9S1UeTz
VbRuiYOs93t69y+Wvh5ibSSrG1MV7Y8RmBi0tucOq0Ov+dXK3q9ePdm9kECRMQag
Ede/Yr3rHI683Xs4pxNo7kcqLVSHYsnj9etFwBB1/jm7vlPFCIBKsGDKZI5e4MKl
5wR+wPbzjAouN2T8mHqFocU9NLxM4sFaJrSsxpefNlbywEgSvSciXSXv90Pn1Msm
zht2WPZN1820bMiS+SxCx1xFYMNZq/lwGJE9IO357Npp+X1xh9xASsgzACTJM+Mm
7BK8CF7zUQ4EAAUqGK+zBmJh2hiNiB0dlBCS+Ia+F93J6hiHXd5yj6vLgq4IKr4a
dbZqpv1JXN9zwXP1B5BJ+4pnaqVKdT3t3TD6RZ1FPxUXMpRztsPEfpQ8hvZTndlB
l9ZCObLNWVbhvFHNVt1xyFPTZUd0ZmaPuNe6tk9TvcUBJuXBH4IglXIG5mB/DGYR
a8k9ds/hK6iHleGSdosBDIbHl1DtdMGpZK7WshkbbzKlw7xG/m+Se4qMEz8Nt7zI
lmWZnxpkFq316dK3zx4e2pE3x4gR+v4Rmp8qwyJLsYICypMgww52wFE8vQCFV3dr
kDcC1wZHKfDCbEasHNMA80MtLE55Kb4xtx/F7jVMEDTkA97pgwvnIYjYrfTGm13b
P5ITfAJUF5Ea7XcoIhKiSXvnT3xl8y8dkhH5Umxn8mJumDS3c7BCvDwXFsTYGeYD
gKK1PT0YHJntC1SM/sn8BvxuB7U6asWeLpJOMyFMJSBRUv4LRkyayWCF4Oy/Bl1Z
tHti7bcyZxR8rRbcjcsbtXoHKNE/Jh3OMQlNrn2nGOz0+F/jlqOzcJgauMqd9IwJ
jKfoL1WnEqJowDpI1nEupT7bV4fJ5G96AMzYXQ1GOaY2P737WTtGZv9csJuaWGlV
W+DDG2O7fbt6qDI8fpGlXCfjADuCBjUGVw88rHf+e1blfvOdFymXWWmaUOa19TDv
ajYG0155HpWBaTCOse8qigJqGCMmOJh1VL1aO1zUvm6sCxtEczZCCwuXqm51AMAr
An4nB2Dp9/aLNTR90CRjSb2tJTL9jCWk1nkpZsiqcM36e8JCtA/N4vt6Rf2KcyBG
r0SvNrQCvi5+dPFZ8Mc8Euu4PmaaWdtVGT0VDZdjmscSGj242hn2b/VDadTVu39b
9AnMEXBUXf5JanUeVjVbk/UfzmryATJH21se98Izwf2u1AEYGW1UlZdXOohbC3M6
UXD38InxFQH7A47o4cxWYilTl9Ga/JvsvswXtvVlKP7jvPlP2t7Q8AZHZ553Y6Z4
uQmregf/UibPm8FyhrwVXt91iujPUXYyoY80xIh+m6X1HrVjbC4qDS+p41xN2QFW
jSr06oOXktkfz6Fo4XbWBrs2mowhcP6hHe7+4STGMZzWb/Od1Ml/bRPDmGGSDYzi
MSxih2b2HEQadSorNPtSKXabLCFHQPOXJY5wpBvvrYXGo293nTCEchM4T8eIpx1N
TcKLQMK2xV1ChBaaoNWRR8C6waaHFb6/ZvCxqHolJ3i0ehyr6JR3Gx7uYV/uSbCb
Y0DAk06L4ET4PNbwdzgydNelrhEXwy2FP/RufxHDA3HNNwbofAkXNu3kUjBboiYu
PEuhQqwRrFb859n/wjInqhU7pwFHRjcx9DpbQu/T9G8yXxyulwnJ1dDygdU7sZLz
eEOo8PDQArg1MrZVFC4N+ptmTBk/6bBQMp5bYVT+Xwv2k/DMFen8vz5tgu1nF/gU
wReGefdCU+k6DFwdbwgIDLZv8WrQMFXTEmUG3s7iBeHHVf72jtuwm+0uh+bEdQEI
r18mBLzXLGIooPvVSFcwX2YtKK1scDT2KbdVcFSuBDeAinpZ2GXlsXUb7RY53M0r
6ZDWvbtVtlmEnU4nJODaOcn7hMKnJ+6Td9wC7ZVIvGW3nAkL+mOUzFdX/7b+FQsk
NEHuQPyeYj95y8q+NypPz6RgCHI0Yf3SthHbsHj0CioV699BwBkJw1YzJ2PgQQdy
BUYhMZoLVJVCM2/DLBQ/CNz99GW0J/BGv3/L5VUf4PofNmxbuZFZjy7ZHaeHPGid
JvieWN8nlXKsNIHkBmOXu/bb/ynTXXy7vCwNOtY/a4TThuROlRR3PJgzKnyk4e0H
jK+ctb8WxYm0l+JCT0kRqSgyhPduinK1yU+Wu+uEvEcaywYVCRkizCPiMV94epew
LeSzw7A61VcJqUaF3/0oS2dk5d8EkOB2LnuyTZ9Cz3eydDvJI9Q0IoPd5MKHXQbc
0RKdR7MbvUEKr8zq8eWMMAVvxHRYfbOASqpP3qN8FLl/eN958+X+jBCM6/iit1Du
bhLiT1LhZWS1ZIGADwrSYrd3PwCN/tsSCmJQ0Mig+CX8K1K6rSxqxDe1rD2EbLzq
VLoXlN/8/rDz5JNezYdsfBfJSPpF3Sn5CB0j8UxXRRsBiy+PIjMBBs4O0GXVWqHZ
QsUIP44VDkx6LykCyZ1s5D2L1mPPHuDebuu9L3H5+KYaWKbMWIBx1rB2XViyiuPQ
V2XJH7xs6K0zuY+rgoQFUAvIf/UGKoanJUfW34m46cJVyn4lpO6xxrkzaIHr9T6G
UMVM379awqzzAQs21pyC/OTU442R+sxk+64PmTCx6MLbrWW6oYLTmgmxTHTXZiIQ
1dRGhnZiv0wS7JTdxQHr/WS1ZhKYru1XwszrMbI1cCr4tVZn9klzVQSIQKLN+Y5y
RW4oPXP2QyUF/s8YfgQbjOi0uvsVrwcx32hV/7htazTOfXQkm2FkcMqqT+EoBRP5
1p2T6I1YMCBqoKQV+dYkCBN9xbChsfAkUKY1hShCGukwEUk57G8kD5djECk6ZUQS
sUoCDJn4lrneGFeEZfbNhMtGxSCGMNA4hLmk9TiU7I3/vGpLlchPT20n6Y1s1gLM
OO2LHPqoaYnozwPTf1DBY6p7FnOdL3Wp/AF/4c5g7Pr5oMOPT619BU6khWXcOKqd
L47g3W9I17QTwtL3cZ9j8cDeoQsO93q9d0WR/YVdOLhclTbhK9xzVt9fl/tAMo3g
aFvMrUzqxysrhO4QTrRXkvNKKO9fsrq5mcI7leVaGzmBHC/SDu0HGADhigpryWgM
BLl7BAgW0yrIN6HktPvTe+SD7Vqaj0OvqaGtS06y6DmtO5fcZSYVDFqCHl09YVRP
IVhWSJZ/sZ3YguuYu6FbG91oLbzc9hRRG6GOJe4AGniNIKqOXCY52X7wnTKYJmRC
WzqfiGQaesRaM77HRfdz4KNpURaqoaToj+AKw+ZHNaSSlYaV0qs4/x0eE4xxOLA5
/hLIPlAH7O4h+YH96RhEQAP4EcvFjUxB6RebLrY6jwhfjRXN3i8Yjbl8we/+NPjU
kIU6jvhH0uCHy932Zku3+3k5Md6HXk6v3nlpjo2f4lCfqKP5Tp4r3+PcyQXJceHv
42PSD7vA7xHEMD0NFi/vkdQETfES6qL3DQ42PlLP1htNN0AkkesKrbrRZIwIjoSg
ndYpl/DThPoiNIfWqLJrXyCJ/kf6b6bRRjMHOzImBIfcr1h6/tekiFL3cRZiLEjX
CwykUGMW7h16jMttLM+cyLgw3WMjwwIbmIv//bs+TS7IiXur3vNDC2jc1LZmhQj7
vRgjERuyoreTvSQuM0pR3nXnIUFtHLTfxF0X1uIKEnc3z+UAIDiJDX3+MEAQfV0C
41vb5B7P/TKTqxFq+yEdtFYJHJ4WBzpvKo8FiqE7DQ1kAqHt+RRB7GkP/dFiqxGs
d6rIE+ONd+eAM/VUDi05R6abfFwEYLGdfq7KIkSnyCHumf29XqaewSKjqYBpYtxz
W7MITxU3cXdaueQJDKfVxyiSB4IMP8EJoyLA0o8AKiCmzeyQydirAUhDKxoJM4Xp
qqGQs8FUp/UXITORAR64Igk/ArktCF5kuK4Wk4Yjq4HGGfZsRH6TLtB5tRLRMmaK
VNVdj7spSgxjGd/1JbRkFCKJ53sw2dUctEwmW4j+9KAP0HRwA3lR25DkpmBsXU8n
yhuWdnIVq8kVqKvlbxncfKqC1kDdMsDIS077J4E3X7k30moZeak1AmQSMHKLB64D
X+yl/xqRAL7wr7Dxf0UBf4dnDSF08HEXt+0R5v2K3cpOtMHkGbp0P1Ct6EMzr1cx
Tmf4bRxdKH5JgG2kXjoAj/YiTaBy02/qafvzb3+BfXIBmBsBK32cgTfzYMWW02XB
+ydBT3cefnautkLNRhrdSPvT6UV/wZcH2jTGbjIC36JQnRt4KqJt1/LZT6MJH0PT
l9PhbgOk0cX8QsHhgyzR6lXkoxHgYFUHe7MlQ/4ygJRSFpi63Veif5N9F71u/LNh
bWwG6S54o+2EEkd73p/sNLAUis+fwSVTjQAUNZuWnZWLrAgBZYxaSgx6xCP4XW6c
xjDTA2hTY4/AdSe1l6Bx58OJwLJjSR6ojaMMS53Ll1nuYfVZIs2VBY66YtEKC3h9
J/qCr0U7lODy0JEL6RtpX5WTRB0evxcZ7tZ0Ec/+Y4jDOhHIRHLX2hH6HKFRjsY9
ec1kCp2fXfgEuC094c0/WhzAXwoeI4oYH2R4m9B6Etw8Z2y/qnMEoA370D+SLuU+
aPAqQTws4mAwPM60vHACqHXEJJ9yBEbxUImC8CRcDS6LonZR/Vp9LtJ4OGvDWc/0
G7wazhZmMCD5dhXVzFQ9ItqCGmYcJ9V0iQryb78jlLKw349gjxw6Vq2kix0KiTja
zhZjD7GepAyRyHsFBOIDjF7keZ5aPOJsm+Yo7GvoUOp8c4BXsvDYjyjxIdjJd5YH
29QEL5SvY/c0d9hUIMNpWLvx8YqKUd/ScCx2lorfDwtn54YA8mG9XIOYfDvJjnpS
ghEtH0RLt5dSkO7oY0VFrvYyiFJEX3teg0tvd/NwjANJZALYxOUAwUUFu/Os/NBK
CHTBFk/sNmSVYyJobuJAI15xUFfN0qBLu0Fv3aBXSaxYCkhnCFir+yTbvm4OIq6T
2IsWWh7Z4uPNdvTEzGNnbvtotoV4TeYeVYIkLb/L+Qgakd5AZJophgW3pKSeFiy1
nQEYS/lhpPmxLjmu7zzdzhb8NslYPyECXPLoWawnec5EcuFIoRhpPX71SB0jD9Rf
fZMngGJJ1EIZrwhpCoZydPq118udZ6U9JypMbG/imZIrUKYlTpl+V5p0O1eBY+yI
GJARP1o70ZpUhd7bQKvCtFTG6TAP5PaGOjUgBT38zvdqUWN4OLFDSAPAFca5p1Bt
4k6Wa6xRSiCRhxgX3/XTAmFEd9kTHAxzfchw6c17QpZxiRH8Sg6mef6HgW5214yF
/deKX07SuXADrQpoHnwOSU4PiTZ9jMbQG5f8pHlYjicuruCCC8yuSRqCGWua4/qk
3xIlQEhPOZVJ8qdSxCIUtt6cjz3EeVbMWZH5xtIbv8AIoL9YVvxGR4Yt5sP2JXsr
+6Akr85HWoDmvxBd/OwOkSR4On6w450SurORKI3raAZLoCO3Jm6PQy+qHHqKnjks
uhlq/5yWJtHM0YUs0TLaN8295CpBxw7fES7g7ZQJWKIS3qwBmikkIj5iCBn1AdPi
PpEiIVPdrZimSwLBZHJeP0V1ooxWORJToX2kNkUJqPInqQ9wcoGXC15ZhDMIiKfz
0T63QoqRBONc9NrywmE1jWxoCYd/dwDYpVe9EIvt/odRLSgFCz3WacI2dLc/PVak
RDzkNGfxGPAvJpZmndLWjInoXOffciaBtI/ZzJOBZ6FWLs3oe+20Dpr5326P/LBm
O9UtzAtgFWq23K1XU3G/7hXrMhi4DcEs5nKYmK/Hra2s0DXH2/2UpIfWR+EL/J89
G0P2SeQcArJssUmf1w8CZhAomOxOzfKbatodixjchDfdGufXyCk+VsACwdGM+2vC
cuVt4sfss+oqyiS1O+ObQHvqb0qpKwEw/HgxSSDTNE9OfCgU65wbiRNgVnUBdrIc
CVGrUHKNECD3qMc8qOj2rwhfAENuy3yDpOB14u5+QRFVIQmHIWZBOiPAY+ayO/wT
VZXE9eUUKwjBrRhwgmJI2CGBCleuomwQihM88Jkld7raDSIk3y7YIfpSn58D0q9b
efL6RYquEzR1j3+24R0cmFjSAWFZTwuDlmNShAm2LY+ZSxTEWGChBjTL6xZDAOEG
o+FnHy0+DHtCj9nFNOX2hfwkpoX+L9h2J8DzqsfSvA/NyHnofqKl0lQ1AZzbjLbk
vZ73utx6l2wSrOXj+9BpyoGS+4FJCtS80c4DQjTst2ygHtAQPbrXtyXEWb+vPUO1
gvMeFpvweCJX0l+LoaP7a2fTQ3h52t61OCmcOkCM7PzrYYQoRN9k58S1E2UNql9f
G+1d88VO+iE7wTyMld4Zc8mqs17CLGaZlOlYl+KHh0upIeVtjh5HtCCmo3Eff8jV
dDlWfjOMt/J1fOQcjKu5VAZV7CJYQlMUCFMuWX/+nUfkje3ld4WF9IOyDLIoxx7t
SR8iGOf3YKb5bPvs6cYgu5H3GXUh2wWnvn80iUwBAjOcogvgP53XYFHXmk1FNWv7
zDM+sal64kTgDx9HC007ytIVZNHZ2ceEBHA4Jp3zCPKvAvYLXtrVk7e24G8vxJM+
IgHjo2s4Qz0ibFfTYr2X7pEMPr34rFOau49jDjflfFnIyt8mtcCYtXnFVZOQM48u
jbMmBW6d/vcSa3KM71v29uhUjftdBwg7Yr30jkBG3sZSp4KaxbIWBdjIsoTfJ36e
M9qAuVs221YWADUpr2GNVJQGmWrmWfR7z/n2tDRk5lFG5hNwTyirETINFkW/x3+L
khjWkSCcYzPrX1QOxEfG22WPYHx3KIc+3LS+Pa5d0SMlHOPAD6+0nY8w+WjsnU8X
bI1JzCz9avI+fm/lg9K7UaCx3P+C7MRSmB9xQhu0D5ffP3tx/u9HuCpz4hYKNNEI
R/Enacns7OzEaDwN5l0Pl5KZH5g0zP1WrWr4DBFlkREYIrjiY8ZIWIGdXqEgRlY7
Sf+QLqx7HErmP9fD4whyGlWxZRwigkbzgTKKYRpA6C0MewC9EhNnK6Op9tz/0law
NqMVplQ9XNQXZImtqIBEV6QabCWka0yEpSgXHFFCXxP41V+nt0M0zikxholH/UcH
lOnYfTlpH6RZ1ou/gpA3WQ8BndGbJhJCOMtAqaKinhb0rdpb/R7gPHfFnXMrmffG
kiSUBCVCS94RcERfTQ1PNzQJVPtVLqiiX0Eho6A4zJ93S+6R2BBqvOSkxnVr4IzV
tjzUdKfyVQws8QEBY/h7HbP3ppRiT4ToeVMElLLWSbn6dnE0yi8qICblz7a9B20b
QoMV1vXsYymPzmfyOdzgUbHlC1MN29Lgq335BgpVrCFhohXowsnU6nfmMDhubGsr
WRCKJ1qPCGyRTiMXLeU5EswoeotGrhqbGCar/QI/22TZiQM+Zc/qgtFrDk3Eo31H
KneS5hsUfKikKzBEVB7s8wpvibGCDIg2wjBLr0dKvF8WUyHefDfl+HfS7bmWEMI2
aNLDtR7u/og3U5MDTnHrmpMoodlqh9OpJRw5pms9QVHRm4qEO5F6tmEszD4Ph3Dy
/Jn+wKTdURCzx60DtDEmU9yemJdwGe79WfZeuIfUhdNs+DcpCHBQ8660oRxifWdp
71Cee4JO5MJtU/MgHpg3Ob59rwVwzg1lNqZ4ywFuNR/63ebEViXhxJyCBOTV8mmQ
QL752ncmnCF3AgfsPTKQCI/vetL2FTbXdlHi9AcYfI6aVeHtTW/prllOj9Sc+rVc
NHNqQuAEoBIzRG+CYx6hkVwq9ce8H+N/st5aknvenMFRZ2MD5G9AaSv/j6O/3rxC
OGMePH1/YNdEeMGJYiKS/bcheVfCPDd+Fb7UTYeLMDK1UoTztEOUKU5x9Qh5DWgi
NAqImEqnUvW5z1kifLmT7gCAYnxmo9pm70E8r8kZrbG6pC9uiuWCFYdkUb7Jt04b
ZXvXj7U+K1nZ2KLGadAwPa52Bdvo3cYEkYNpTzLjM9APf5/zQn9Dg6hSWsUNMG4L
XPMxLwnKYCUiSSEwNdMcLm5Nc1GCdkNaCbRyqV8qauTgR6r0t7hyIyQ1ezvsdvRd
s2xDC5XYk5Tp7ilCEzhA2lLcH/xJtALFjPD73p99C5W3CpVLZechdMiSS1XQHONa
UBJ6BdvxnmNd6HtprTktFtMl3IYiuSPQNrX1EgbBsjfBLS8rBfv4QZxrj9/tsTA+
e6LwzcXVaMzLIvbR3OapZ3QaoLHga9ApA32rV1MV3fKwBH1t7izthT+evc1cxSfc
kpZaIxoQ3wxOI0jzCiY674o8ivCX8RFTYoFfi1bmvAJiiR32SyGTZup0IoJU5bvy
UbTRoelKl6Uu4TibNBJhSfXVmunN/WWQHaBWzi+gU7CxUmxPUn5ScGLwSenpPS6b
/pBJOpRxhjLrKzgOH+AAlzz0lnnrUUryA57iaTCcyR6b5nJ9yC/4Hxcx6AQEAPEV
1TwdkNpmhUPBg+WfaTie0x4UfQ9bjOnrQti16LyUbP3bkTtbLocT7BOUplFRrgQN
SXIe1sTseZhkLhycNipCCONAd5O3zVHfXqjsUxvl5fgWyTI+JNdyuh2DQ653qGVZ
Qe5XqDmSivOKgGhdcq+oIzjbCZkT+BGJQExMlkS2N6yL+icjgBUQU+Yy8qKVUFZg
Sov/VID3coVDB6APIwakQPqKwL4NEaFko+7MSxWZqmPtGqDBNs++ife+L+t+jrG7
tCCtGhMsUvIwFV1/oJ4pl7oHMYtylZyPIFAiLN+YNu3CJfIy6+Rjw6VW87GHTHBy
SJiWTq3un199imKkK70tygpih591k594HWDxJDibcN45rUBOZF0q3gfKSuNyqzr1
YKBTQRIFoL014PAaTPZQRi1N3528VYLPanOhMaU4K05WCIV4FcrpBHCN5ui9ZthY
pIZbhOvfluI0McU3WFBttHu11SoRE+vPrnC+8r4oN3D1PGwDfPTLcwAUh2kJQ7rG
Sm5RM+mFZB88i/FVylmOf9CPqx46bp73gWXGQjhmO7zwYZzCIaeolg1GXedj8yKn
SzJ/kodITffVhen17NXjsCb0Qbj4N/PQQ9MTkFDtRN8Ge3d7v+Z8MAOaeybGsois
AXkTOCQvo/K7mTncRxYQY9CFw77B2rYYlfyBSpCTIFBKck0BiavGo7viBHRlnrwG
b0rbegyEC3XkX+u+4YOoysQGnTMvx2V8jZJmACdGX5VLbZEWMhD3qe5MlsLodeCv
bnxoaV1UrwGpOIom6JD6W4CGT3GkJ6+1IYyJQ5swWIqNd2tmAyFeIyRsE8d0OaMh
hi2xN1Dclizo4WZb54dS19Hk+bwJWggmEEDxi2XTrLeL/AD7eIXEdPOrC3c7+lf/
A7USbBlHOd1Zd4+nD465P4YtXmBi9jfMUqZCoqXXWk+be10EgRx7I/QOr3tLunlS
jSyS0f13cTjkeMa2fAUlJIhM11emKEOPVYLa6P9gwtvqus58eFc5xJw+jnylV4HY
mSWYvH1zaQ2DJ4Aqb93YQWCOUtb2Umh1UJ48svtGfeHupXrjjyhNmvPibLgj4/B/
iOhGvRa1OLgoo75pLX/gIveOgXY3gpQFZoHZLoS10tnXjkc0mXaFe2Ie7ZdfL2nM
8aHkl+uN18IUFeS7bHBqPmDPwEFhLiUI+Gr4ajAfM2VjIAZifixJiTIsmGbOsgcS
pHmKBoAUgWg7USh+jy+vcogysrQI3hYZwQNY5/P5sPrwpu4FwbIxp8FVCbWw9vcl
W5OLF0Yx+AAJ9ZED/SXJBH0WSDrOdjKQMvbXwU7qb5PVoeEtWMw7RxgkkipizW3W
weXyQfZdIexR/uVy0oQipB1CXaQOgBQ/rfC0tL8zsoCcTh7KbZw7lDZ2Ceri1+Vu
W6vhMnKMIyM1J8UqeJUJi4vm+dhN8ZOQw9LE/qp/pPQH0aapLn4h87X+hvF7oC/J
fOxkjxpLITAx9B3HFvTvxZdl0g8aSkywBM7HQ8w4qt1BwzxifUiaAqjFUuAcM8MI
0wRaIyIUe56B2HP+0Yfai7MOzX2g0wU4vKepd6XPPxwdUzx2kErqJUQzkYHTwi8t
K06yAOPfiyQRtwucs8nX5/3kH9mjME0XWjarD6qhzVspU5EVZRscKIHfpbYuHonK
77IHMVpya7txvsofLNxKABl1flMaWaCJkHu9shOzHHUJmO6HTDfi4JGDcn0MBxe4
Ojby8c69k9Y6d0Hn6oatriyRdSydQ2J4eMNuDd+8PXL4frxXCVQrM6ig+Sx1CuRJ
28QfcQho8xoyeGpcSOnH7HUJ9VxgiTMZChVzdBqoGYT2ZcHlKAmnWx6D2japLIGW
Kd8tRMF4eyhgUkj7Qq2/xeMAO2dRFKddJ2JF/hDmMCTJag9HSyt6outT6YIzv8LD
vGDJABW3Of0YJJLCYUulQWdlVodDpxPKS6arRIeGVds7TaMQF2ErttQnyCHNP3S/
bCxfaci8oV3S6srGSzjEmcI9dlTjyM2sErH+RMalSbr0Ae0HH8IGMgob9vgX9Fvj
av/0AhEnkgqhz4L92NG2dYf9tppDqCjax06CleAQHdjNNPsoSQoTTDrGiGDn0k0J
NxXr2usMvjBEiDsqxY+s3IyDqmvgfdEf6mjXvq70nPj404gqPvH08XH9zHXS9/gk
/9LyhGZfJKTEvzh9Z1K4ebjCcI2jdRwP18w9xz9RAr+E/Sv6z3jhlf6r2gv1GYJs
0/zqGBzmHWpO+DNH7+DwOqz1Rai/lEMyB4vktPqc/KCfk9PLSCRM3ZiA/VmSnGqq
CCkJjsl1Gg0nIjUR0A56lHARuvCjLfZaKK9aB8NL5gmRi49apc6KeBtRM1+ta24S
Y6swI5bIin/4dORKJnhaHiLn86RWGHeYmxu2KVP0KQN/y7yDxLWN6XcS+ZD/eQVO
rGhdvOKTGlnwnHkXQzNKJspLgdriag8ytOoNFUgFajI2DWtGDJjOEwMKWEv9pL88
Qr4FWMHH4FNe5tAzzHXUC1oR8yWn2FyvwYivGU6Apday5qvX0aBrnX8VF99fzy5j
1Ur1ygdpRSAzG3l3cR9WGE21/1Dju3N5Fl3OE+bh2TR3khH98UVlvBK9AGSwLtrX
9MFsCnVde9hc0Ml+v0TI9KkyZ4+xUsIbE9DCA9qK4spb8PGR0SRs8ADx6DO5oskB
AjXDSxJ7ru5NtIgP7TsE4y3rdDKlEklkkXdHbX1Ni6gk0khvmVqGxe/aUq0m0EBa
JGZZ10E2mzKPL7tRZ+I1RZW4RfRZvjQdyY3jfQ11SrqAEJbkT14jNbuk+OF8Tv2Z
qdAZkcvBAAdejLK6JzeEbh4T6NMYIRNRbI5M+N2bWzZL9pNjkqINXupR48jWQj79
Av/ILiecNXaRXaalzh0L2CNJMwN6j9EzIkL6Mjqoc8OURKjgmGiI/SWck0fHmHUQ
gBS4T9g9Sv/GISBERKpCL1Q41H/itFCbdqJ/6UVuIMeGaOcnFX1/Is7YJtytcqaZ
rO0YU3Za+wyrt4JUEaN4xE5NmP+mUYNG9AMbJ9CBAzh7gN8uqPgkXIAGcqSkeqTw
Tgp4WBxM2Vv2cuEAzzrM81ZaVLyKa/OomQ0sPBn7xVOLyj/I4l0aumNk2BGLwMTe
BcIU22nieWWG65YxPAiLPtcGoFhjA3zNP4pb9RxYDQmNnrc3cPajV8HvGDtbbtw5
/jPk0OHgPf8SZddUVFXyAVlv/6IeJIl3XCGrvOMIr2nytk8dDWMrlZrb56ptD23H
ZSK+1pvy2wS9cNcnY6ggMJ0NkeEvZe9AVBlqql7r3tSyv9J4W5rV/xoQ7IjAQg7H
wZ+FhPyaitiBc10UeiLTeQx5BJ4GehGmozzH8I78zKc1MzrdZukk4Yp+5fPm/FE5
jYNvpnpi+oXWCROeH8bBnBhCwM0L5+RSKdxgmragmeIbarVz7IKNnZyUtuzBzZeB
33rYhymlLNeyf7DZy8LpM1A5tnJDaVbUiyHDKBIBWpJArkszw4ZS7MipO13ePASD
uiBXjC7dWz1JGYgzBjiOuLWlRXOUIYJxICWQ1xNVJcNKRHMSOSalXtxSduxJ2DIo
O1mv6180A17FNXlLnNo7o4/JR1XEKq9vHHbwV1Y3U4BwZT9G9a48iiIB8zwYQtc4
N5ydYyGQMLWgc7AdZVoLWwH6fHS+ngE21hPmkwxgEMITVaNFioRXfp8fj9E7oSlx
C5uN789QLipFal3pYp2gEQSegs3gFLuRwxmSGYzLyhua9m7AJkZ2mFaAPei3xI4Z
2wr3OyWaKnSkSYHJLvRP9OFSXQK/cYlUtTg48uExL06H39YDPsSE6hweiBRSz+Fa
y415jYXQLCiRqMErUux953LNgf6VXFIFMXTJfgaDMuLzy1DUk+KoDeZMa+BNLBXV
AFa6NTdFa/16dRyKEIlY4bOwGcEdNWL/jZTWnmWQu81WkIPAvdWxLasoJVUhiSlF
r1Bv6eNtalKSEwhRdBlE/LXH3rnxgpvLDGhVzqL3e2tAnTacHwSiLj+TiSBacMBO
qUo7YLSM4hjMsM9SODQ27S7tA3HfD12BDXv6CeCaUN0Uv2efJV/Qu9+UWucgp/HY
pMZPZoe2e/0IxTQ1rOEbrELe1yfldj3pSXtDqnBad0KDBtI3XXJnXeiM+0qF8ITe
ZrLzVlzuX2cCTBXkxKBqObixAsnyyv2EkllVQYmebokyuNNju/uIzIi14Rs77nSD
coIbA6l0oydrFI8cc2JAMnunKJp+zMIoZUuqGwrnDkaWJDEcuh1/OBQFlTqKGOCu
sZ1fVV8+9Luvge6GuCu80yoBEXD4jrXMsLlsGacTpxu8O8BckLc2JVcewKtb9m17
moradX7dtNKGElX1cVty06I4XLNQMVwTES9Zwj/KZq1GC2xOiMUT3xYANUsjzorn
tFhQRr7S10pyAEFB7M3gzF/+n3i6I1ENO2usJp2OUpwn+Lzux1ZCoRxG012NjLeq
URGbMwJKpM6TSlHQQHNFkg95vejp84ehJbBrCqbicmHROqH8PNIS4qxUKdUxeTN7
euP9Rt6xfaAt6MVR9UjATDMVlB3e8FWL0Et8v9uuR35O0piFvlQPPFM95pi35ZDB
jQcDCXzgAb91sQkSuHloTkHLyvNbSH3GYXnJa8z9/cf7EelMF1j5GZ4PWIwfJ2vB
9xjMSO6Cj/LB1KuRG7EHSMmKNHIrhhyuwgp6NQ0U7vTvko/xpIF5IsNjSEMoVvKC
UQNmR21G9RzSBdIiAzaKGlDJgyn/FdKvojp98wDosA2PweU1vtqe54aW5NOiOQJF
Xa4PX/t3gv6Hm4AX1yQUL+Wtni/x01MfYW4YpJ/DwcQ1ZXyqCu2HHtDqRPAuhxWa
ELeLtFfqxVLjzBl107fBuYVdvk9kLfJwoRK2wWo0cdcIAOQuN/rH1tzlchHJAbUN
aRnb/UgDNUqmkYx9/19mSbnPea0bice47el0W11YX2wsYzr7DUR/JTwK2uKX53IG
PMwLtqRAEG7Ys8krXVrQ1JCydZ2/ufqeJRRSpfilPL+junHfUNsAp9YJLTEtbz94
063zcc8BsO3+FDA+bnfJDSVK7iF3Nc1DOeI7w4qFsk69tcfsZ3rsp0yoFfajUPb2
b6sSrxuenlZlSLbvXeKdIZj+/R8Cp1grom8ToUjR+1efrX9+Y0WSiMxA4+uVdvih
mH1ai/G74u3EVY5WymKZwxVP4zsY2C1qyq08ptD1C8aTJlfTiOFT2X/WnrwgLBi0
Qa51kmwIoCs8YpPkzlA0Xg0mMU12jtOaoFZzxLuwYtNlQgT9LvfYofFaS746+SHd
Lun3gbNCDrP9HHq5KfZ97i8jqZjr8iPsMzqbKzlhKrKKkHrcynA1qDVEUnC3ZI9h
xw/JgjVNCA0toTh9QGJx1OGgOIPSa7fEMEbmOkCgEPgEH3il1vciiJhm5nle3whC
6FbiITMagXY0wNesBk8+chTYIWjdJUqes3AamX+ynwNedhzNLGfZn2M2cuaO+HLx
lLmIEJ/5IRcsejgzYoQOzcIegjlVnM5Go0Vl7b12RHUY0kaUQ7llNLQ0jrb8Qn7B
+HQiXSRE0mUdbwjKAnX4Rq/obXTvsKk6qmDcDu1I2yw/+R8jwZlw200lv35Hv0+2
jgj4dxA9cDS86QTev7j0LXu5YYB9q0g7ufwU8jUlgnWwQh5iBmnqOC7JQsH9gBVh
qaS3kGRmRYyK7VW8Zy8mHUXp0EmFatbCnhVkYg5M/bGEXhT1GHdg/UI76kn04CFW
fT+kDu3ff1T2tGXLeC6njRm0iUpvpsNwHqKiDDt6v/bDAxPaQGCmh27bTDz86Bu4
yGNTY1109mDX4wD7f3huFFfBjJTq7oG+Un8wr32JrLjF53uGjpqNo0siV3WLE8Et
qLHaG89ZbSizZiS4zuOT9uc5PvC5PaAdd7xyNfcrpmhF5XMRE1sOTEvoe+a0OMuV
nEm6OKhLfyE4nuQzlIACObYHEB7IMsGkqLVQ9KgdJc9za6FPk1+WIRr58oz5owqL
n6EzrY7E+z79GMvJJpXvSyy3Kj/3/oFgB7PApp/B8gabhXd1iXcb7gDM0QCNgAM0
ng2AJKiCQ5Fx58og6JGCro5Y0nyhN40xgj2+/B67MiUWB6kIws0sIgglcXeuM1bI
tX3UdLCTKHcBSmN/W18z4GjmKRBkHt/NBelXT/3j1NQ/C+PUui6WhMT8knTCFIK4
bRunamp06BY+NE9jTAK4sKCMDGIHn8T6L0nhiQ5Qwtn2DwVMUipDoQq4UCCC9Kn7
6GelEAbYXYDyj+OTLBiKybQGZQk9Qx8AqBL6ydHzVkVgBKCWpKaxpW48z1IYNi6l
6brrVXyatLcMA5nNg0OEocV5oz24vGx4UEDbxqVSXMhoHJm0meWuseZFWo0YiQAr
421cJ4kHzj1PyJMl5NjzUoXWP3KeU8Cam8UA3g8mjS9KfeLiZFZ8h/oUFS3P/jfa
Us/dY+PfJEr0wBWoQTncn3Xr0a4bzOIaI6v2SG+9rQEyKMrXHa7g1hZb8A/uwx+R
2EehHskOHDbT+2d1yz3KvQ2CeItHsOtg537SI+1jqVoSlvmkbIj/W7cQ5tO12rOW
qOOmEObjXADWROdOARxMggChERjc8bVqq03NP7ETlpTe3VE3kr4SAMjT8J7tdFsX
atuP2tcfm3NBWEzGt9KYkUTpzj9LMUa+HoFHqdTfSHl1nNFm7WRsHrP570usuGWj
3HzIybttGd7xHL2lZwXgXn+8QEBt684rolGVg6kSYuLkvMnY8piEBHxMbcEGyPZj
Qlt116gOdmPXyB1rDcG9+vcMJRryj6vGngHt2PJAkFtGVQ3BDEohy+V+1LqPidrh
dqay3lXJ7yFkIAV3DDVZSaRlFtz16HRPD7BNKGPdfrGzJSoJd2FSFhqEy5dIfC7N
q1KrT5yG47ma7g5bBSEympjHE5EyjInacMQz3WhQ9mGp5pX9Vxf59yraNYfrQR7v
f8keUP/TZkA0SEtn6wd5wCocLNPTC9BHw5kqzR3i8oQZK5Msu75EGdIQWi3ZketX
a8kY19X154ndyOFhIGVFpyXzb+5XfIgspMOKx5KOJLB/JlGhipNOo47bXQJGa00e
dxZ6H+5WSZzWOfkOCf/23dCsRyPvpcswPwh7RK0ruN2Of1MkqTaRxbmZfHBWhnlu
suPadrqSIlScv+CC0YetTbobGdv+AJrad+FGtFIHuJ75oqj9/zP8Ys5yyF5vOpoC
tkTBdKoqxpb8RHe5EKgqZ3VDqSCz2JTP1Ljn5uv6GaSlUFLKUu6VFNTq5IlZcQ8T
POkKiAn/xMrUyF9JuXiNELqIxa2Vshh+JpwDd8T9SJl8dXi345MRoQu/tvKt1dXP
fL18Qrdh5juRglimtDn9Al5NsdxJeK39Yte4TVrfKswNv8T1OxxHLlnnIejj7TY2
1APTHBIkWCGLkrXJttbIjaH6KFOurOcC4r0vhqtWF2s5vCK+EqMt4GAjumPK26fO
jwxQOaHzBkb2YCohtgx70R+3FltGtL7Ur+nNY99BK41msi2VsFprLxECM+u7jgjt
DifXH67BYrOqxkATMx1Ivb34pZfzBHYKW1xcTzIzZJ1RFOaCss+fQUYq1kRudfoI
+qGdIFOHnqnveZDhVrdxF3WMPKt7PqxZt3SH62Oilhdc7O3236XDp6A7WjlwerqC
9DKV4XgvIERJm0UcOMUjwblGJZw8ZhmP9DRaTQ582JZreIOKM0/d2G2HA395mbx6
fd1HiB/zGQDBSl5t6FCT1wBnsVEfQ4fXX+vQz8sDsBoxGErduitWYSSEu3XYJfGr
CEcXeMnBMCBfCrGxmByyqS8AONU2N7ugX2h5sKl/gVIfk0ajk7NxO/KiIgnXG3TR
Gim7Tw+hn1J1qkp5dqXzRx2dHmdSKJ6fLDDevblWuVish+cOkPBpKr4oz8iYI5rF
WSXQHKy4B2aqkAU+z1OIBrMw88nNByZln8pBHF1eORlKQiDDd0p1WZ6Cs/5OM6Fx
katHkVEzUdZ77vHK6k45IrOS/GxHvwszKdcElMrTdvH0oNdfN+cFklpHzrmKnTdk
6FAs0Elw1+uT9kNrlJcdY2tyclV8rEADnHWRfU+rUHr4CJnjBCqe33CNotSJocoV
531GEQQ1E1rVGrMUa7QTOTbga3Tlh7haaAxStulOEdxFocfWPfkU7/cp19oAsszX
3X3lkKsxgPDCizf1F2646I0v1oz/W2kgSwlcWR6FRyesniQoVIgpvPwlY5p3AD72
G0udC3OgsLGXTbph1ky2BvDrltiy1hsUjoRJHWZCuwaQm7vLtThm3fBES4Uf9e2D
AkzIZhjgdVH0DpxeWDrZwhv/OXzfz9fbYiNOAAxGgtNSEfUpN8SjFSNm8/MP4jJy
QUYdhASlRkbbKqno5oqfls6CUJhZZVoagz7AVNIx+0qmsCeFLeoMQktct7uOo1kx
35UKclULexP5ofbcAEt60seIiQtVbt0G2dech0JPredKkJM4DQPcNGaSTtlN//5x
KU3j14jU9sOgEKF0unz/TKOxPxBEFZ6WB0dXlZU1Z3+5dyVLsnZzD3vcG/hMC3qc
hP0x386XVHuewzIAawx482Hl5PS9myCUKrUT4K61SBmN2CCFF/n+8joS+fWDjuWV
Z29xwEIhd6C2GVYLjznds16kF4muwjvi9ZtuB4nOgFTw10efQ61QHspqeK1oqEUY
/3vA6Ux2chzvPk41WipdXXUxiDrU5Ba10tjFnLrPttuyW2Xg9efjFHFs8DGB+WWR
0cXTsqpj/v6A+Bbd3mmOrD3g9qgp09zqoZy61K0Yo1G01ATBnnbCDYR7i0Dih7xE
NWudaPXtb1E/bnQw5EcNSrnplh9hX3Y3qrJxc64kkHGAoflo3Dgw8i/lUD9LH1Rl
6ZAkx/14CHiBRr/dx5LqLxbdi9cAZKOjNzqZIW5sNX7J4yITdttV1v8qIbuHO/yH
IuvIw/MQDR66rhgZRZRwNRhsjbdulhRb6mDlEuCt4y78c+Ei9yrW0MPKXmdBDhzu
92165omwqiqa20YKzFjxTrVOFaphAo9nrzIfb4+cWy1M7PhLg+6YXsrk9O+wA/Ls
XiSAMn715w7dfUTZd/p9YBpoBp3QvBFtTVavKd6XKiB9hOb6rRjedfYh/yjyjyFM
2gq5RREvJ0kXv4zx/dGDehX+1vylCDJVvja5I8zINSN1hpodLI+5O6nwroRM5bjB
WzeAhxDwtNK9JDRbQGhxq7Bek9F+vof1ORuoovnPj15y1tlX4BgX+rSX59uMBB9z
4BVMsZ+e1a1C+1AZ5bRFMDaPXXXWF3npf1QbpGGpz5SlffI2BzM73NT+ExmPeOqC
d9C4wpKjsoLkvHrFk2u3kvFxnkuRltmqEfrh5JRN8vF61OhY3Hr+wCp4ZLu+uq/2
JkiZvcJn7/bXsI6PSGSIAcSGLrKXJW6pzEkS0qfuniEhRqdx+z+tXVY4UTf3UN9O
WaobbUDQvGMvGqe5XjJGFj3fpRmYL9EE/oKFPxUukvYmyxn7L868tiqykmuKDKQp
B+KsrRwgPrryRWnd3ZTIldsbwKTtjiEhPyLMSRbkxaWu2WGfivDOyt7Jh3kRRO5A
QJ9AKLQgdTzmPRSk932TmpnhClJtzyC/oKG7/6rXnfb9Edss8QEMI1IzozlAuqTL
MxyTFunMDWCV9o7ProSF3ErsEAiSyCEIZDShU9m0sFQEPEx5Aqm01wGzXv1nIzOb
6VJh+dgI33NSsc4P4heUwzZtM+o5yWXg5vUbA1m4CSCJX/xFb5umMqrDjZhS1u+k
89C53No8HcY3JOQuY56+8MRd3WOFAXScxy1qU6vS71cjmXWsQVXO/PL0tXXc2f7u
Q7+Pj0hkC0x16VlPvMkGqzoVnuIAsTnpzG8EZ6M1gppiuh58ei5L1De5pi+ffoh2
DjdVZt8Jk0AGOwZzfiTLZntz5LcWWBn6Eqr87xatlzXRRINRvqVq21EHSOoqBzHu
rZvPXSfLl0+2HiFN3gNqX0cREousf5VUCrgUYOOZNvTuzNIhleRnjLtRPl8XIy99
dWOeIP4FeBnG3XdH7x9O0mTi1ore3EYmLkknIm34ooYKMuHlfkeNtmiBq9bzgQo+
uFVVDkSCwRbjy/FeW2p51qn17DcjKdyrj4lQx1YbZK1Y1YeBwxzrnohg0XFl3rTZ
UNaNk3R1mZrLdJM0cs8s6uxZPM3GC+kRO4x8/YwKm+icqtgIEfITCjmr7rwDONBo
JEkBGmNMyRz9zlQ+IaGNFhPHJkVqYFd11+ffDyhz7Y7CMnCbOWzTjIH5V9NfWpgA
dSgXIgnAE/ZUDhLjt7bHN9aGxcfJmszQ0zl9XWht9uFeyA+168B7y7eS0Lhhgan7
lVLkR5c6WwrqXbKyy8wCNgMFSK+EfshPZDSPFZohuZZe753YYNVvkcbddZ2TfySu
iF1baD6e+wnRKMAoeRojCAbBT8YqUJTxESAjWUaXDiAZ20rdoEnJ6gbbj1cz0Jp4
aeF4aJ6AntGm8ccJ0OPM/dXLSMMaPysrV/KN9OOxo0Esv+YhGA9auHBZO2zICojF
vCNQjCZsJ81aBIhLku/bySob2ZEF5mFY+lIU6NNqVe+SEJXdMBhF75Ulgirc+XAt
V5KR0d/8uipgSQWqlu47UAkfzWUp9QRjhu6guOjg81ulygsGAp5G3PC+BLTzcmPv
vbZK/eaWfSR6HMsQCfFfwwpd5KAq8dnVwKujLNNFsuXeQyBxGj2hhS3ZZGptqAFg
t5IhGHof6DYIuW/Dk02t1wn+B9Q/a3lE49NB1k4B90du3sssFn808WzeKIu1Cva1
8KanG5WmhF/hk3UryNp6BJfYLY6X+ZPH1xsHbx/58qhmJKnts4wm3FD/1+T51Oty
l03L4+KdG6/zPZ5borhfa4gCtfae8QonZ8XmFoLKEnAzTtftG7HMpeic3ujwjPH2
YEAB+ePBgfirykB4/sK+SPRtd5DDR1SmmJtX2yOcT+QAqBCszZckRhu78W5Hukk9
dnxUK88S3vcQ3dKeD9vQvQasjz6iD19B3HHGZJ+OIhsXz70PEwrjTEub+EXx8W5O
EFy4WevCgeN4eu4rQgnKgCo9ObXkasXa6ZdIbQO1HxvM0L4q2nhYd8APoeWn50KV
QiVG1GPmX8gfCAmLcKg7IYs2sjYtOGch28HrgMijzZ9lukpx8BGtgHJCJokPLgup
EgYHfxKeFYMEi9J1JuUMd5YRIafsvB9+bk4VjSyo81ixMx8FjnFjXuLzLD5zimUe
eXsL6nnyt8LAKPlPXGyEXC5DckEv0/lPNwggbHqQQGZxSzLP9gbboRGT6hbjaURu
z81i/q/5nAG/ZuKU+xzKOEVq7IEBz4uXAz6g2FdbF3bj9UuWK4dAa4LLA+adTEc8
hZ5a1b0KxdxxrNG4cIJ4Vc1BlEm7b5hf94LYj2cZb3XUCoIACe1SbPDYJpM6t8qi
GvVstVKRjZgx+Gf/u8Gvirqa9DVJqSAxckxKngZW34SPZDZQj/D8sNibk506J2g9
2iwR/5uCdozPSjF/ncDmZ8bS6yPAjfN4fB7LpfO03k8eycBlVAXthJK0Rci0cd3+
vpiZ4s54/xH1GtzWapwAn3W2gxrvcLDuK7IJLmhkNValT+IwSzAv9Vlea2w/6rdR
o8X7NloLixYzmoLdQKO9JqqGrE0S7w/116lg/uObtQpZbyXg/mDzt9B9+qg4wAcM
H6VGOd2B+DYXgCDp+JvLnqD0kq7axPjair5SHu5kzl+HJ5cZxKK63qBBlmWDcjMc
5v/HiLQFpLQepMGD91RSZuDZvpmXGATei8UBhZQZi/9w/zU3mHZA5X7nD7jFfJfK
828muiy75RBL/qEVNawsaoQg9+argQKGvPrWZRoEQHpYhwDOpdQssoQtRIn2pxnZ
FMvZX5NWjCz3nKvdUkCOjaLg293QwnMHmiTOdc7HNzCCxNadSemrc6a4mXTOOvFu
ZyQhQRvX3pLiRbIwXaqHHuhPpLFrANlCGLrJydx9JIhC0gQRra0zAmCnM+2D/4/l
sxhd43vEpJBxgcHfrk4Hn3Io8EKJpOrRDI5x5mqBMgsf0zFIqKyvFlzm0wdsofmM
4lGQ2l587GV30xLklMSDlhyjAF+QFeDNqlCF+AdktwR5Hy/amdzw2ESvlY5ABLa3
MnhjUx/o0m4n0o6+JRG2ukM9L/cSeH0jKNEvWqxDspBK2t17pT83MMRRRvluxq2E
gaaMbdigWQz/UL8uA5HbflToXDNepCt/N/banaT5BUbujQZ1GXigSHsbbUEylwvV
i8tjOxxM5a0HiDWhOwpqedhW9Uzs3RLwJrAM1mHCsKchfXGeYDkBgUxB5J+Nz8RX
PUEFxdb65bIbJd4xjSNyS2yxZk1MPSvqcwVxPQJ0iCGqXwCP/r7tV4ZHfykTahcq
QXaEZLErgmvX/Oc5Ec+ZvSLGtRdQM9olGegFBioUaENJAf5OoRDI3a9EVP+dvzKo
Ol25DpQqj3sIaBXjstEw/RdvwA1saZ12eDnO1O4D7BcJpnbN9k+csRkLwsKbUWDw
s83Yba688cFGHCJpIPjnSv6xl3z16ttcx/RW5qIOSWBD4FtJMvSuU2r5iL9OZIZl
XUFpTF7vEtBy27+qY8VVsWYp4w5vZejI1kcSJe2RuzkxpdvxYXWHWyS6/jDhz/Rc
jE6lpKuS9fJ3elRvMpOyL0n2YUVg2uMbCMiPYF45yHKx+cmPkbWCWhzT9xRveGwL
u1O7g9wCY8MxkrBKcsc5mPVtHae6ONHa9CIQbRlFi2JeMI/Pl9VzkSBGoQuFOw6F
fpNGkGfdcX735P9G9cLOpLBlkqpFQgAGD3RLGbmriV6FDOgepudqrxsnNWAZiEV7
mPsD/W0ygYgQCou213psMa+SNRrsKeuw5XVXN5YjJO/dw5lj1xvOTJ3yMKSE3+Om
43p5+TMr1YKhF2wYq57gRNZaC3HB74K6cIh4HY8QwJzr2eWRL5WrCENLqARswHGf
nXTBlt8YfiNz+qrCAPbAnMtErUIJsZxNGrLVaaNp1I0SRMKuHR4IMQjnB7sb+J3V
gyNqeTP88+qnaNb3MK5wfoQ66Pd8FN8rPxD1xO+kcdPczwKSRORnuoxkc59+DZLw
3jzTlJ4hszgrmMKS6DCNesXUcTaz4c8aIi9vm/8gbQU26RRU4X1bBL07HC0rX6gK
tKbV4N3fBorveuhDIAn0BW59Mk+1xelqVTk3kR5wU1Dr6p3TRvaAfjLm9WGVtmVa
xYSyxWEpXMndViHeH5WWPeg65pnz8CpN8JPiqPgVFZXpN51D4GI2lREruVnaAG0K
fiN0JIP5wRhKVwrkI2PGLMwoFrVGC2lD/P6SvkWo2/5/4jzNXlOWLzNQYsJTmI/8
lVA94tGa9Hg+KmjZULEWjGPjt3/rT1s8tXE8irUOvMKF1gjR9ReDKqbAXVh62yqx
KSVq+1STsZgD0BBfU4R9PzgLdlmSQKZcK2NrCFlmCYJHaVRE4ss+Irp+rIB50DkV
wDpaX/d5F0R7HzHZmsOZMrNM8ehE0vgkcQ88yyMkvITfL7EIsFM1p7FBIPzo56+Y
I5NA7Ege+U2GKFdy4rMuLA0klUg6QAEIPwe/ENvWJr5gkHz2OTUikf6pWAL/kdNY
u3v+JYfRiJB1mcQKyv9aJgOeJDSplNL7VVrnanCJ/u4duwvlublHlUma8s70j92B
h2X9m//3WGjGTc9Dq4vzupPgHRYACYxEoFlCa7a3S8TCbVKCMuyEdcmXKsmFsONw
Gxq/BFRyIZddx8R/Qhq5swKPBElH441ncDMZ7UaTxf8JF2RG2WPihma2dUrVax5J
zD0My75e4FZkK2s8k5Qy9wAITgqblsOdx1+nEHh87PlDp9GXkz9pgYs1f59zim7b
WCG4dHOZT/4Ue4a/zhglsRmPDRjzgzXhZA9ov+OcmLBeZa1WB6p8Crj76KTccLtb
vGmSKy7MoOzvfpwrkPkfdDkYzj2fLo7+n5zg4T6lqWz7N4bQV/xLSy2Qtt2bZX6U
DmOz5S3hROCF7O6jhxL9OpXiNTM10GLGRlSBCAKqWP4JpEJOPlL993OBmpj3Cubm
s+MGu4bwdDyleloUsOa6SBxnFJkJrUEqb12f3y0LiHS6K774Ipw9mhcNKL3aH7LU
e5huMdifqJimLu5oAGssfZpel9obhumFtewOg2CLsABc9jd+YswwaHUOEH+bs3Jn
PY5w9txVJFp0BzHTyypw1EGNCBFfLDpJ7YCP7mhFP6nZiQ3/9yETOHUJXAWy+gVb
+FzZAwwI0jyUCL8PcNUPbWAwWITFneNvCjayGlXFrOfuLtXXsFfePd7s0meAafWI
3ev+vq9iNbiiY+JXIntgi0iNVmSZ9LIQ4yjw1d7jsGb/J/mEEweVuqU525UXTPoj
RRVPhhxl4V8S3I2pXfse1qFCWphOuGkyJ4lwuWeHYoH2yZLQmenEHqsbm/UyAv0e
gjI7pOBPLhzC/IdsxzJmnvS+wHDMOm1xafga3A7kIeBSuxKQrbW7gnRlFUKTI+hI
+R47g4cTe58M08HzOyqBGnxxdNRwv+j1Y17kWwmtxmEgP47sg0NcnzCUawkXT5JE
xHy2wjk1BB+Uqq3Wygv5Gzw/2E98NH1oErFxbno4v5ysw0CoZpSP0QpZajaCK7QE
xAFt7rGWqOkcU1zUG8au+l7uYu9AQf/GhWmuqTFpsJxBLXzfmt+nXSa68r2Byzku
YOFFcYr+1f+prVQxv1npczZMqruCSTSz+dyFjIydShwimvD911LZcoAJ6U7TywzD
q9iOJ3LwQ1YWbwKzNAhf0SqF6mT7mjmdJiZv4sq/rf2xP0U1vc0WUdIUKoUqTMOs
mhVPUax6Jl2QKeXN9PK2NxeL0vYAB3sZv3aKz4a1SekRPozD4jSBNk0M6gvvenDE
RcQ8RsicgtLrwjhegUbYwkL9nI2clqP2A96OsOnEu5B4u5F2QplesndceEKA+2GQ
Ku5mfIwYshxRsUBdm4Z6/38md//8RGuFcv/W/NgEzDgreonSOIwNJ0KTYu9mRnKT
ARpPu/53JQm2tpbC8BbexdJbQi8lgO4GZgZ2EdD8Hx4gYlLvLzbnBK1dJi9HupUu
ZCnf1FufTupK+r9tEIljOFqy9XBKE5+EFdVTdYAHTtYk1O4NSQR+9TY3FY4hCtQv
QAICx2GWn+ioYt4Tx29ZFp7rSuIyyXSdmD1V7famlYfq/udcOpMyckss4jtm/4w/
JqOXlJ0cNMbAg5JzUg/Z4lVyctnshSah/yi2MboZZhdn3l2xI9xELkmGWUGbdUIr
IZVpFKSFjYZC9uJH+dXvR4WKkXp7OcI+7JbPomNGgnFks2yoOnj352bZ8ku0es/G
+IKSAHI1JC62DOg3lt810W9TqueSyTm/Nn1St/pzvifPpQMyrsh/lgbpZkUU2G+c
ujkXOFTQKAaWQxYlsFbOMJDNqDVDEMwiJqmNl1rRrrfakXYRirE2MCns5ifWqSHZ
o+6OCc/bWrbwnRT903pDRh9sFifWbB43Sk/c2FbAVSRM7ybDGZeQn4wf7+mMgUKR
z0m/DX/+p9hag3DFn1oDG9wI0fSzXRvZtvoZzqthw6QMMlM175Uw1NVEAm7g0JYA
p8Ve4yJPefmExmzEX2CFNUJ7hq2sSxkdVQty1HhnIe1dwYt56IdJ1+qMcaBUn22G
IXb1sMJvGtOmon76WWv2lPvijKz0w7X15scfGgqErtx1NybPMXA6XMevE+ypUTf0
b88XJkHvCCZQTxtphk4PQX2f5U1CFXwxH1HWYdTFyH7A9ff+rd44k3ZpN7d4x5qw
3B1NRG3IV2Gm7DG9kwtmL5g4u0tAXGRIcN6M4ZakGd5iM+Ruhcq32kc/xsXPouy2
8UWz/M9zz+pSF/aRiqyNVhLAvkbLD5FaoF3jXDoxRSLhxKZjkuz2Ni5+Q22CvXxx
uN2PUP1SlEGVWgeHngdm+MHYdTPe1216pTh762Teemg/suvMe6gBEL8y9aSaeuh3
+wP3r49SAE5Wsf7QWA8Q2rbGrEcBwbelf5IWU+jEYgCTdiobV40xOuq+XofMYy0V
fqzduVJTLvg0RRCYupNQU/W+xwgj1/moGQOoy0ye1JjhlPRoWYbdrNWC6Mapx8Ib
YYg9U9EPW16OL/Rtk2XgnhYr0LD7KyWDqAV42pnq6qGUp3NBlBIljzXal8/b5eKc
icDrT3OlXJN2nN44hVRPALdroSdKdwM5L5uOTfTIlYK7UrNRHkyGw9ts4xlbmazr
vzo1rmHStx1NsCBTfz5QtQA7eHhxY52/Fr/S5odKnt7PAB3NzRgV2AQEagTVRTqO
UO3fLh+64nvRuxJnuFkyTobtDoI0PD1rXLVBdX5tdltWkfxWSme9Z3ITm2WOidjD
9jITIFnYgoM5u84MKmjbJeM1Js97Cde3qfmae4y8ibKeQe72V5jLfFvJoGlKrLIu
ozQPR3zjje6h8ev7Ta6sqohmzp0QrkIsMFiiJWD6LTty1qYsqSCkafH15zEMA2LU
N6iLChOMnxqgY7MBisjkYsohlEX7tGvYEEXEQVTmpsA0mwlWgArOenSZKqpdrRxq
XAQTvDGj+JjUyVwm+SbTKl0mRJYIx+Mhd1tvGhYjVFJ2jnuDmRxcB90lMuwlAJie
/K/e9KlalGqrdU9gkZI59IhBA4xnsVO4zsWHHndHAzwmUUhng5A81WKe16PKQp8b
vIN5GxZBUBYr+dn7RiyGy0HbOuH3gteSTuxu5D0W1P8rrPSIPw7rKmvL5/06cL8T
thPTf4ejfjCSxTvCxNV0ZoZddgvWD+W4W/kfH3dXL7uWpuSay/AeDDSTeHPPSQkQ
hAQlV5tj16eeS7FKFuJnzchHMFT1LljJNWp7wttmyTjEwWzDl1RnG+5ug60RoMbf
pEmX+r06YA2QytIinszzCpoW0Kk55lQK5RV3DpwhZJfrC/z5zgdg7+ecSjYUgWNm
0kRhZZPPHxg/JEeuPr+Y2mRncpvqhZb5ZPi93nzglXNanNuxlL17vChbc8XaB9S9
JSiv/WoMgl/KEQTyhIqsHJBAPHIkxDBRrgacZB7nN98Gu5JYSAvO+12A2Qsw42Fg
uPtH6sZ9YrABgGGpU3GbsImDP8jm2Oqrfj+IjRILhoJPfoy/ITuZz1zkzkalDBY6
AZ5lEx/TRh1JCN4KBZBpItI5TCJ1yDhWnfgWS0msnpZxln1AQp1Ik9iTuYszpYPA
erd3u8weAaoO15P/eDAyvUOWdcW9UWRHapL+TwmxEhhGyZPbkUkGIiKThvS6ceP7
tVbuLMjlP9dbbzi36XqsoimKHUz7G4ARG2GL9GrraPTPXSUzRuxdMc1IV2UvmrtE
/401aeqDgmO6QEjoZMaa5UQhbUV1ei2ohnaHlSzqC9zionHTcjPBB2vMNhmpf53L
Eyt2Rho8605/n2dyeMZDx2M2+4/PmpPaOpRh3owqGv0l2RDwtiIoDNoYNw7RfBj/
gFACrxBJLJD8m+cdRtf8w3/+3L5bqyTGiUArs74RirAT+dUOk91RvBUdOW8qd8KB
Fpuh5bWBFugwelOq0H3umO2qaGrkFR4zG1F/6djN6BWDe31f53g/c/SHguQAGzq2
KQ7lDxrcYQqSnANOsL8Rr0FT8KXgfoXqqZwSaERnucITqbSrLni1iyWbB4HM2xk9
YY7lhx+oQv2aH6yPB2Zn8ktgU2+idlmZHL4sErlRNaHMLGcvYwD+qDzQqzC9X+P6
nUR0AfL2JHZcfOTPzdN+9IZwSdu+TqhvIAhTb++0hS3P7Gi1CHER4LUywX6OCQf4
EyzgL7g/x+IojEPBP8LeXeB+98YgfIGEiL28xtEQEYj2+TyedyXEptvhWL+Zt7FL
JvuSVC+6tKoMtt30XMO+gk9RZ5/Nm0lN6I7hYooFjrTUjSQPw5dTGN5HuNUgIbvO
WJiZKrQ1oqz+5cn1ER1fx9M51Dj32cg/r8O7Vzt0iYh9b7F4xvZIiUfOysL9x/b9
Hrm+zJKJkBG2suC4ukZC/X0B1fTCCdVctF12ApGgHJbgJHXsGnFcBiaoJi6qrRpb
W2yvmD69Isn04gORIs8wBdHcbdUh3NAFHg1L+RWzViGqLleHWZqZl+QBaQeZ6sa5
TT4qUCgqCH+9AXkBoo8rajULKSaKVhLr1/UF/dacIJtANFpv3/avMoK7xY+H4f+U
tg7LqSC73CcVhtZWgJy09w5eGZnbMY/LjXZTTgPkhuNaHJySUI8/RREDLMu44vWK
3R3qhVjl+9Gy5RKP5SlXG+uUMy5HNXqcxDVk7BQSTtLs+aQTzzf3u3m1I9HqYmf4
uKaBOFpy3DpSkajHTHoSBB8oUJgkmfH5lgOAb/a7Zvr2UUP44kJOr98wa1NDcWbW
D8rnmGnsMKVYETFt6tx6KaViSc4VaUUk3AIQG/l+U474hIX1U7PC9xeB7WtPtz3+
/qTRB2OtHMyJwT3dnBaMp+gwz2Pq1FJzG1qdYWZr4XtCZXqOkT8S2i5lRXBWZi5h
OJAnbxlyxtzlXbeACyS7yazpNMNJ8/Oaz/3tsAstgmlg/IEGTNlfDuYuFcu1AVwY
oJzURg//Cv30RF33aJaCnPY1HQJSjjT4gnoTP7T41OHtNrwUqG1b4c3KNS6yRAaE
5SHp2kJzn7EkmBpOK4FMOGheAFA4zfSIJo1zpjFTjcPNbH8lPV9uRgDnTePjj7T6
BeoMcWDFmHfovPjOhHmu+hOEGkZPwn3Kg5DUKMvLvDFPaKGpovNGfo9x6UZB6raY
K5DhkQL8VjmGuSYPO0c5Qm+DlUl44wNTrEX/XxjSKpg/MwCAXh6m64D6SFGlvxVQ
dFqiXUeGy6wMbbicQIcVTPvNRmw450G5uLBQXsndFxi1AdOsxLgTNiIggRFor5eZ
V+zgXg2roLPvDgEl8UK05TT2cA9Zt1Ghh7jXOWFeCRYVPrNc/6DRlpmZdlmRnU2b
PnbXxfKy5Zrwj5EjI4PhoCWd52GvSepeCrqY4MGpoYlr8MDYJnOR+i6nLBX9uuHd
JGBVj6+TrlGK2uoEY0eIlBNjJzL2JPBPufh2Ky7WLlkMmwe237MAoK9MjJx67o+j
/K5TBs4VHub8XM4E0iC2FWdRn7S6ZH6cTDYQZXEbFT/Dc2m6OKCT9Wo78RUJX0Jb
SHYQI+H0LXz3kaXWjO3Ao9B1Oh7670H71xIGv8bbS2lVDa2RNOELI8M2JgBtVZRD
7ojYLD/gJdgFoSdHjEcuD4E1jjYuH9cqhHFFV8dx3d9vvPFPYqrLRD4GQXEKfO5c
VRDm57v9Ip4lsEaJfcnuTEJN7ct7vaQqQ1iCLwPOFEct7zsMRPWwQCluzAVnVtWz
u7yMI1fzSJPokv2p/nI2vdeGqLHf5yZeN1SpP8vHLag2Yuu9hcr285VyVxl4Ghbd
XNnd8ZQ9tvXrLaCYVGw2fKUBddxfvL4Fr1FFijFEKSkJmfMlLM7VVsyJuO7xbn/W
Y3k+5y3u7r1Iz/3DGwm/odsZ+hO/8K5/lSlU7+x3WLqbx7SoQYMYtzOJjucXqey0
VzUQzUViFwodNaBE/sCwnuFWElN7fVlucZ6VstxTB753skd5MW1oBwmB/KaV7reY
8Rz3sUl0QaK2yyR200V9uPTtY2Pn1srXIaIBS9kKLkZjq0wzMYDl+S/Txuel8mQi
41AWI+60UgIO8F7ZDd1muwPoizD2416WUtoEuFArZWObQPx0ZvZGPGAfXzjdOCsh
P9TZ28EO4i4Cg/o720MLOzlgB7qnFbeJaMWt/0n+FM+BtURtvaB249niW22rnKzV
7vE8giaFrd1hGQ+jIR4Z88vRdqZtt1iyTAemmZOowXctDkeB9qKSQzB+pDUtjvYR
CXFBLcXVZV3FzPYOXRuOko6B89UlllGU7l3fbNVrldjCLWJ2IgmaFwWN9zRmmIPw
4BSJbaIhIehy1BI9wDsZ9Xr/6o15rgc241OCpWLhcnjy27pyDhWesHC4qHB/GGQE
J4jau14+Xck68PY6bHKC+DuAzTDP1YSKHdeuG5dsfPFiQVyFbk1jqaHZB4Hqsori
MUUlae5sSrzRVduL980LFEFnZUFEebTpqCI4QYYl0VYfnbrvmHWUrAJECQW1Os3d
tCOOeJJO0VhKB2uvc9tOiChXJ3RuIN6AdDL63jsCBt+JluM/DC642QRZGXVLh7Re
p99vG3qLdLAfDBhbbnrZ9zcjxGy+Ca6jhEl6I7+CMUJ+zX3X3pdfRiW2wDz3mR33
K8/o7KTQRv1MuAPlr84cZ5+4gXYsC89o05zpArWgdbcxluVELQGxa2w2/V6xVvUa
57TmeNzUNCv7yXhmtrbsexufUsT62p5P94yPhJDcaV2u/K8iCqT8pHdtSgxrmLvM
NjKRIgwD627+YSttDZptuTdbFvjO3vBw3fzzb64A/l+ituqT5SXGydNSZJbgc0Ty
D9gGybEfjZMz0FmsTu5VdSBRFb0XYhnfGBk7u7V46FGkYACvVgDVrYAwjUmJFJSa
cZxA+WeFmYcNIDXvvfYxW+3RD1mdIK8qnMd9yBTrkr/RUHF3iK6EqFfPinNj+Jrw
FmduND1DyiaN8eZd7TEQ/55c3Z1n1x8L0eItyE3osBlBK/AZ/ajCS83L96RHstwo
I0lsh5WWSAGD8yBDBmqCKnC3PwJ+5LMMJ/w1FPyaB7GkvEQHYu95FNGt7bU5iNUl
CZOEmh7ASH4agOstHLfFnBuh5AU83IIM6da0H6Pq4qw8IlR1bc4et3sCsNY2SjqO
l6x9FoUYKTqwNtn3y0m93dtjpRenZFVIuLB7k/8xCB7iixxL69fgpywH3KQOKN3u
2TEzqVokMcPORjangZzNgB1OuQ1+0XmMcZQTK2WxDOTSyLKV3LfjSkdnK33zOQ/a
I9KUkUyFvmh0sPOEVpeZ9YRCeZnxuUmFR7zeo57bvtz2Lr36nS50zHX4kgaSqQcY
AeavJc9sa4L2cLPpl97pmDmrTu0cTekcktF1TJqp0GsbbyutgpLOTvlluqpjrqII
L9vPdZhmEUzrbQC5V3FhgeXeYOg4elgdBZxDxOTntdsu3TlF0gWcD9TOxF1/liJK
tczbXR/59o5RVK0UnmJkh8zmX+O89rKrpbQumWqKesRu4kbRuumtjmkls6sB8V88
RdyYn4l+dKijBASR1r4MpB4hx+IOa2OJFmAPPDPrMntwvqQN+WCN5irA5t5zrMS4
Y+5fUcbzm6pZdHgUz4NsJ7nvdyqAXrlq9TfzvCAGws/I8bc79IV8hJWh9jiS67cr
01v5z63/LFv4Whw0Jwo7CqzSA7nGgXHMt55XvU1H28WrFrkRkLRLy5cGS8yGSK2x
QQ/dGGd7QIUCwTyYbb6ZD9rYV/Tt3RylOOq8fUbHNvPLDCERsvFnAYHBLoURglyS
MNSLgtXC4dbtLSKW7XO9JonSYj0wk0S7llY0dt6/+NoxjixQP8J514PV+En/Wr+1
GhJ4N9MC707HvDFWH0O12WP09sUrbXw1rLQuDR35RELBSfjG8bVVDgHpVkC2Mwhp
qxOEWKYxx81h/YEaROruZy0w7+r8rrGuimrVGKRyu0x7kJvav4DBaSuSBSiikYdU
NF142PwpPWdSYIm81dJiqPb6i316/K9bPQTqO7s+PktVkz0Yd6zGldbK8dwJVk6r
W0234BIid7T/wCjyzoiBq0MB0V5fsHL4qYjVwaa9a8ya+S/NE21ufFBYC1gLj0VH
jK6F+E+OM5c8NZBzKbAnzrtsN96nU3n53mqBXghHlQSgcFsAo8sf4UxT+tF//4JH
7nTk9h8A0nllFRAP2QzSSzThwbo2t9Cs95xrFe5rylxUV1KEPQEcXV9Hb/SesGuV
2OxHHg8yVGsYfvc80GYUVx0j0VQnzWxRYJHmf0PJw03+Lt36kBHEj9e1byX7VYbd
BOP7C5Gq8X9DAiOCe5oADXNOc+rU2MjL8O9M4IXsAWW6mDi/fUPZYJe/OiZszIbD
Qnhl/rIW0TOOwqqPfha4dRT31Lp71YLugGOnjnl3jwsoQVyuzWC4LdxINBxN+HAD
NbXbajivusnrsFNauyPe3aGfjKIbOU9BgSw7hygugs488YjswKebHIBNzr3DJHNG
V6wbsG69GOl2c5WV7fHviZyBIGorx9Fw8yQxUjNTPkC/q7l5jyHLdpcLgv4ejsMZ
akj56l1AJmn517OUeyMUWdrhAF85HGDv4GUsyNte4F6ZJDVhdaNBcBsDHoGAwzHc
A919CIPKAiqgJ1bZU5uqJYnjymwhthnlW7X7yEnLPQYGAyUQclY3p/WlqG+bpv0a
lA3ocAgsO+ZceoXz0fmq0ccoUA/ZEpXYgETtmC47osYpjlcvY0hmiMy+ADA0UK3p
f3flvVlCjhJiacEV462r4x9o57tRl15RGll66NtsKkFv4t/iGNLyWunTDTEGHGhB
GZ06FNRTLqbFpBDSs7QgNTmEvV9bcjxkfomDFaUcz3oJcsetNIo1B1J9N3Funkmp
1md2mj2vmd94ytxWCmTMUh3Xc0O6uBpQvNDK6uTkBw0osUmB11E87MAa+bqXPHN2
ggejxtFk3XzFhyW4rdDiDNS+LGaw7AqE+Qh7QCJRaz4bZINlptb0eSWOJmHXLdJB
Uw1wS9FuUAO8Ew0XGVMM7AuhwSAtoCEio0ugB+5kA1DttM7CfPob9JFmn3BtweiT
caQKvWIVMT8nZcSlfyQZdJGg/RSd9zFEIy0/vyD6QHfueGYVscVxQEy02YBGguln
kV8OK0TFNc5FgrcSbs7rUme+7JV2P1Mx3kgidsBGEgWC49ITphZlqCtl3/UytNcp
qZiL6zuxrhZr3kX7eyShw0lB0R+QEjp3PyxP+yn9VIM7B2JwulgJDWUAYUsnFMv4
GKbED+yxxcLEfY53GFE+k1YVN1oXUm9PUcf79ralCa0I1pJulGxivZnCxCG/66ew
cArI9P03XYX4gADymf92TCkBpaiMot5hr3AyLAuowrC07QOJgj4ItoRYb6mxr+OF
t9ipg+3g3Raib3AlL+N/merk3AYB8kgyPQI19nZajIRTIMnuaghFuYrSv97tIi3t
YKd5RCQkpIBkbqwq2HSMQKQUQyIhmJ7PKOJCHX/47C1Z0POmvHlm+lA+rekBTWMh
xyNQPjJ+HHjO/6ikej9Dp1B3wMtnpH9Ibht4SmcbbwfTTTsYmfTil36Pd1fcVcje
+qYQZlYRa+8Ky38UHG58dS+dCLhLAuUyvUar6QPBcBUyEZi7Qhl9Q25EOFzWr0PI
I5Np4/zMt3+i2C817hKe0U1UySs9E7VoXj6Kmy/o5PftGJGroGTDvmF3vxWZt5R0
9V329aQdm0kQr7mubanQGEMLX2IewhcZlL8e9TEn+dNz1k6EBjwd+uEbXpFFiJSG
Nbb7tYcicFQLrkLOz0W37pcMfxQ+UZ4kGilIX3+lPiur0NGGvdxm6k2V3lXEhZxJ
GAEqo95NvQY//+dqbA/aNn4n8fehzvWGiMee7oOpPpu9hZXOAq4TE8z5iqyEysvk
CPofKDNf+Wct7g4T72CbatjJXDoeNsXeVLtt9zCkzhwIIHxitcO88jOhwjev0u/0
EZdzm2Ji25GkIh8/Yicc2KabZMkOCCFgvzbFti0AthFMh0scdDwIQksz3p6qsmaz
gAQNYOrEAw9Q8e/zBuaPDSEjBy+zRO6uh5/nWzjemkOoWd1bTX6cRhrouVUO8HHM
lQQrHS7cmgX6GkkxyhSaAMq/Q/wzUHCe9QOm2sgNCWXvYdZeNwxWdYdydgROnFOT
gOmcssTiiwbdRy9qhUw94AKOrEXVjv9Of3KNg4LNGcsNLj0YnY9ekUpW3yRPMVvD
SSNcylYt9tVDo6nhkOpI8b+exA2yXSbmpY224PhOAEgUglKuehz9fyhtONlJQpV9
7uvVRDkaYH59IXO3n+NnTmrv0gw//bB0wkSr4Qk+Qp9jfLLfhsUYbHMmeB3/NIH0
kwaqMsJM+W3xRFqnFP//SsvrDJtxmlGTIZadWqEKXaEFcC2QPT7/OV9kgmVCvHFE
AlKAvcN4MaJQDMlxdc0i25yHp6vjjEMpgEBj/9DWlb8DPsDR5zXbE+jNvadym9tX
fjzCOB9shNJHDeLeOO64B6mkoS80ImA2mcRwTDf2d3fNnRGklxzITE+rfpYp7TnZ
AZMwOvGkxIDZ5VFWLbZjSGNY3Sa8Z7FhI83YOBjEoKuRDAfCd6lgt1qSDvwjXm8l
jX8KZ02mwJDXMHy/OO5l6kkNQAaJJb/GgPCfkoQC0fB7I9vsEBw7knKZiJGBcnmZ
vgBfC3Zm0wSdHUvn9ijrkodcvAVYIyqtItEUcCJDVbMwmkMzI2szW9tTNhifLgPN
9izR6eH0OD/Ah/udTQg5nmUes2hEq5XnZ/okcyYhFh9MkFzcgFv6yZJ51ojEZ4JI
ngPclhbbaswmTzOV2PHehZ5xgB4tCC/GJasR8EgKeoGV5NK6W+MXom+KlueCSyE8
YGXJAV4wq6pI+TWON1CE5RdfCsBgSwZgwzDq2PztlMmd2zvmoFwPiRKininVcwrV
qSYGJIgAhmKTB080oCZA1Uu3IEd+U/J3rR8rgXAZni7aDF5DgoBI12sxR2mRKK82
9YZ2HYswTuKHzdZfa4M32LpP1w78WXcdhnp+uHxTgDjUy5E4CEMZ+2GhP3Y+IKm8
8EslpM9CYp1ferz3zuzV3PuLnDwTYL8ULB5RS657zsVHQiWv96zkvDkcFKPPQR7o
Jodtb6AGn6PjMULcrhP3fUymXiKRbuxgfW2nJx/qOCXkBZZ38rqj+Q8AeyWEWFZG
MF2JIK9dOKuBo1DD3od5b+ih49nqScV0mzyWoeg8OJ45LR4Q7qrTTY6yyx58qOLI
8LyvzSWp9f4wcUM8fldmzojqDjf2VdViHkyCB92sjFAmNwlAxlOMj8zhhV6GbWOS
vC04aHHcxmgGe8tw3+4r7F5Bdb67UA8N0sHLwbnED+3+B0c2G8fVSeLFRFnMYdWV
43gOmG98JFtUpbDGYV8kqnY4w4DRlFptd/+VFzQzZ9UbuWUwzQ0fOm/IA3aOYtLc
EuRAdNNgfwMxrJSm5k3U/kkXzlx2d4viEOTpTnZSsT0IY9R7Iz+rkFP6CXIi7C/u
hVw4Ejpk7NTDZy0rkDIYuTgiFYNorEinuQ7Z33PlyKbzw0Et6C/3RaO/sAPl//o5
B0XGAg02kKR620DA7kVnHW7hOg0gFzegYdhgDPMlX8WXhi5sqo/o7mgembqxMCUA
gKQNRn2XGOVsMp+UCdZrhiPx0KAgeahiZmmFQmxAAS6qZWmylF2H8cjY1UQAFK4c
IzvEYhNEsyNM6cdxjtGm0lTIl99/fqwG1Koh/QMTfdUOgMaunvIxy+1oldZvimKt
Dk52J6+oh9A7xJWl3gRK3mUsaqcQIu8iVV3AKtgFqmyuQaGA/RreD1e3Ixy/3vTs
Sm60UNiWwsWW5q65Dx/S8LGOommbOuO9sdL6U8/y1UuyLQBdVNcSx1qLQHeMzc81
RqYo8nKSj8zJ41emHFL5NXk6lx1tnSnuvLtOA/mn99dT+57noHMHgQ5FRxeK/L4R
QNXGh9/SnJArNxlDtQLK3j0n+ueWrlzZ2Yg2PWHS+g55xDXkBSmPebTavDRXHuKr
tEwImODMkWp7+l3iZXd5vqAkbuTbeWSJhA60n1tStjhY9ZBsoaDdikCSqes7eB9p
OMTSNgDrCXqWB+/BkGo99s+z11N09V1SmAusnsHASXQOYzQqbrSU5w8ibSSqU4FY
Bcf6H+5Rv4P0kUw6RH7/iygSSkGl6wz2PqZzpHNsLHBfXSLex9ORbXrOQ1x2cyae
d7kUIiQ5RlkwK/hofsv7f+k/TomCicBsLQO/JJuebv4xfvRTmP/gy0TzBzOBWyZN
911B+XjS54nTVrgosQheX7WSqMOA3DDylR1pbTq3xlXhQp8fVjwrULSnaX1WohzY
c8oj2Qg2M1+HNJR5xpqviyTkQ9txeTfEhAwKiLNUXHwNZbqpCia3HGDo7H/A2MYY
pdWwiY0d92TXVM77rPQGkfgp5bX2ZHqkWwzn4LXW48rGKAnh4/cge/dUlpj3No4X
EEEI5bu2CWDes5qdF9Se1xuTgmKN7JFXnhVmQfjze1N85V6tHOR0S2MtLYWT0k1f
XebLUtS6ExTb4IHQjwYqH9LlzUW9pkO+AV5qG3tgVkdZ5AVBnXqWAIF/EOvvQ/iM
FDvZpmo5/HbDmOYiFxvCaVYJrpx1HF8Hh8J0a1FoLNMjJbddTYrksRFRZhPhOJRy
p7c7W+VodqH5dslAri5byNBmwOkh9RS3Y+1hsUl+YSFW3+RtjbDJKP+0QN8X2blT
hwjKqSn7dwzc417VpCMiJCRV+GT0Es3l2gz/muqgK5vKroSDS/13uCg+zi0YRcuT
J8acEfEGOtXGud8dQbZfRuI3LP4LEQhqnzTNateEQEYNaWA7tSTS0TgiDAJeSu5n
/7V0vhXsZ7gyi2tTAt/hMhSZvM2czar8tv9lF4MLivahKk6srC/sHPUTb2RHFqDH
+XCTqlQDHXC5g5C9T07w9UQpQZLy6lw3OfxOQoTrumVJdrs8CVZFIOQZQgRzH0wO
FsJhRqo9lp9krzSuH4EN/fxXW+c+xkHQL1t/pkV5K/0khv8+0utaOTkN2t0hSwRC
kJKN80Glkqq5IGQ7w9rfcnrXV5LInKz/5acktHJKWp6v7QclDNA4JVz629jvX6hy
UnJdTB42bVStOZpqXEOurAWo06A+UjY0+IVB4uFP+Y9GdDOSNf0QD6RQs7KI7Ax+
dn6sd1xGAXxW/ktY31VQglB6O5hhwIrH3mTLhro7vcNizLniTRHHZpnmo3c6ZYna
f4ck17YTESACSXtNUhXs00+Rl08lvcdftjsZIXXYsIfYYfNNgm0nngfmmxIdU6t/
bpe7AO945oqOSoMYgxQ0U9iylPNzUVOw9RAEPvIQn1EKoW8wimzn8tb6G4xPjfJ1
9G0MMswo7eaiz255/liwMtoVC5FQG/FaJg1eKI8Zg8Gt+488a8BmZkxxVI0TFvu6
vnfzAkRBhOLOAIfIqeTI0z3nFpcQU5OnmQ/WqqDBw8gjHHn9LgKEFRuHyyvoSbut
LkLZDl+rjApa62iw05TjTJ/kjU+nMcjBxbMmXglwB6Yyx6KgmJ+pB5Q+3O/PP1yH
JsSSTKNO7Eg53PZfORggpC2WYwbnpuESl8YXo8LYCl2pT0Cr1npXW8hWsAH9DqG0
Yh2nQOJGPsCCRNc69EZjtTkQ8C+YaGJeN9tCcZLtoTkA/Wyo6heALHXQ8EEGX2l/
UJfcf9Upe47h8JYw6D3IlO1xG5Ir4xn4q7e7sJJhSkUYyp9NWm0xlFqS72vlTo5W
yW8LEKDfUQmkHCAGki4lqc6kat6v+2MQOnX/r8fz7J/hZazpeK3637vo+nVHLpID
nPuiQl5EGgkpokzUNChV+qxeAyOH2rGbRnuHUDtAYleMIxY9sAfQNn+lUs42FoyU
WRWtiHcvbo0sx+XLIrwWOyfgJ32PEORN1iuN5Y3ArRemSJbe3McaYv4eIoP0rXuZ
ZomlZ1bbKUsz7TIvK0bYrJg6V5sCGRAbiedvFPwSq1+4+cKtt4/+xOBcTDNsORJ9
OwoCrKlSzJwzNYX3X8iPJhevYwWi9XCfzpMbAqoVmLQ2wT1ebZbW4tXyqZyCmbDH
WRlGrbeZL5kPXN2VUpU65ioNNBXNqF/WWotcoJBidqiv6WGppV/V8paMFuoj+C4V
3HepCTPCuSmh1teybKYxrUBvhwLY5Ln+NOn9CASJMckNENXovAF9UnhOv7G1eU8v
n0aT1Jh+qIyIdXcx76UOViYQwh0UoF2/Ccu78jjgyO0T/swlP10IgCjq47YsbSe4
wurp/5kA9VIQyWC+vJsTMbm+JvRQDio1/0St4fejNG+pCCidRrlsIdSjyxhUzHT/
LASPdEYLOgcBnft2glnTGV3YRUvP+wchV8Y5Q9nif4KvCE5uENZ4L8bF8DbGWyZy
uR2JPeinUtTBwDdDjm73R6QkOLEcsdU2Za4nwghppiRyLvTS7ZacjDpJqqL+iuu8
UkDu+JhiJNg0bzDYZd2soZnPamJUqCtetyh0rbbUrt+vyn0j25xn1j8NkxsrVizq
P9NLxwni1nyYDxMKYpkqsDf/ORIlshz3g6WH7/YXVqBuT38I5l7HmJa+5pNqFU53
ZQfe4azPI+oW3/jIvd79p/aPfuL2XMpT+AxnT2ydLt8YS3lwUnTfbmuvOiSbNGfJ
hwVDPVp9Q5t37w3AeBg2p2bWVmJUEmV4K/Ktj+gmSRp8WFuvIQ1ERwjvfxT1IH/v
3V0H/g5OS9DIbftdxn5oP1DTUjU30AN77DP41dMPjsOuUo0t6vMg52iivjfrHN3i
Jufupl6HhL2HUNMaOlBSYzoAV1iLNxeaqQFGp/0IZgUb2ik7ih5ctQS2qsvAiLfq
VOHJfVgzkXu2NXmmNYAZl9qxEVJufCOuQK43ztH9k6AOVQ/iyiQPfwZAdYdUwokP
8D0cgQG4xuR90Xf30ET2kQMRcaEfTfV/BtNTkAb2xUsTOZXq6K2lH/SmV4m5F4pn
fHB8Bs2Duh8je2yhXD63bRKDb8l8v8KBLshphwRkknkpZm4H5DDGKdOvDx3pEHIk
lme/QwjjCYhffASXhBPZmYfztXFDYlGpTxYOB3u51jcp1eDC88nEmNbdIqq8NGOE
tfd2RfX80fdCiZqUAc2y+YT/eDgkd4U6FdFYPEAPtSoNs4tNWMSPT/vPogpEIk1/
z4OgYxDJRkw7Hawo38XmkwpMeWoz9/qqIUq1Ggqgitif9kj+8fDiqTCqubI2WY5C
srUWTu/NYolayrN3C05GqGO9pwc56vljwBKuIbyDTKuD90N0+p2VdRjunpGjKG7b
N0F5Kkbv8M6sD2ZC7rei/33XxQFKUcBAYqZBKmzmxjEifS2QolEnglBE34MhPkWN
PMu3i1+Jb8uum1HOY47H/9aLLcjtyyBbs26yYVCK87XpyUs4MeJulXxcPUaAsZ13
DDnMD0GmZ5HYO1Ds69hid3uMm9HoNMHJINA0PGz5KTBYcD0jU5D6q3nbqBul15jW
lBj3DRrAtNYXTLvN5Xz2zX2g6vAYrmhTbZdJeOn4nfbZJ6RTPiQKV/LVHW3/1H0u
m39kgSHluqnrtVCFzZxaRArPnh1viADRl3N6rWaLcLUchm/qHkWPb7L22bdamMHd
FnnVPsbhc7BcCVekNdPfyu1MdpHoRZjlIwlSWlKOHqifqgH6TJWCp7XDk+C7Rb4o
J7rpaR/KlR12goB6BFaWcDW99cS4KEe2AkFkun+MSm540ShnksAU3GkFvw7boyVI
1uQ8TB1KLT4k7Nm1nH7/sYMBIgSRmpZR6uScKW067hLaWAHmi6kaHu5ISJbrzcLZ
N0vT3kjt9eYywgGnvI6tjf+MvTJ1JoeDgeIe3FZBD97GgTIgPPpe3uz4rTC85/BN
fJQ1pzKo4aOcKQfj6W68DmVP4bazPCbvVLeuKPw3a2Rm1wO0E1UHFCLZEpYXVo1P
tFW26EVczxdHUaUDTVGjv9pZoaCooE9Lvb/50lj69wyVsL5k8EsRiatUCQwyj4TS
b5WN3EbJZJ7XjsOpyn6yhomL7rz51YvZzT5vaLkWlHruNGxpRBo3cHuSSErhOkUR
TWJ7hpfNpWJgx5zqEO4mxA74acDsP0nSx4ChvoEDkT8XA4pw7AW43IFpuUdxNgEf
7yPLEZnQL/8PLbh5VhOEXb2YezpFNxNDlAVn888wnc7hNPMP8CympumHwBjmIktT
oqKlVyGjJ60pzZrx95ah8ZHhT7Iy+X2sgn/NPgCbVlBUkChTyQcp9/Q0uZlgr5Kc
LoWaOkRLJjerRPB3mpkAUAR7L2WAJCsrLjomz6JJ2LeSc8JKr5RfeDNhnW/mp4SV
IzZFhc0kpxgDRjYoIbzHRbPT4JP5KvQYnmujkAkOqFGAGECpC3KufZMCnEtUGaRd
BaXXlmRKJr/GmZTHdwZmjPl8klMyOkTqJ7LUPsIEPryDKE4oZqUeP6boNMHiBI00
H2ekfRZ4e6wEXqzQZ6qUebgqeAC8F0xG4zlLgdtS+aoRJmfYJuRj73WSTNc3qhqG
hqLfkDxQZV7V1vwKdF97g7argV+xnePtOBNGXw5EdRlZMv68jgoqA5BCj726gfkh
TAS4NHifnQmhr5t+Lx69ioIjX23AHrwI8JrFjREfm/KpSpkTF2tFrHhZcJGyrLCZ
Nt0s8NrdRgMKQnW+xOVJLkiqwx0nDFYzL57g6+c3sDCxRsoTtDioGjLmu85kjthg
u87YKw9QfbT1z574SeziHeSYAArhKwT5/wF3Wz1CrYr9OkcePzEYnmbMrntp6r2a
iWwm2nQhJZYowL6aE1RcVN8Xgu3I/4LP56eabjFXrwpPhSgcXQ7oqj1xt2CpYvN0
a9PlDVebva9j0IhMKq+n3VscXCUsTghVkSpypK3eFXfPGOEx2tBUIxKKg1P87NXP
cdzXN+NNpYyih55CEPDJcJlBwNzR2UjfIzRidhxw44V4DEFfiNTonvaPIoKrSCT9
p3wxY+AP17/qZ9Abg5QSia93LsGgI41E+bkdkYM1K+M/zy2mt8rgpVJSgdhQobeq
TkDYtVuWOn7q+3txY51b5h+3fOSHhgAJpiwSFJZZwQEYRLbIRJ2Vi2Wdb0Lg3wAQ
D+cna70CghL3nJ4ks0l4+j+teqVzpZ9WdZucJmNPkCrWcSsUEFRx4E6UMT5+N7ZK
3ZpvnBHTiufaYhqw4OGH+RFuKFAWV0k7KPKrNLbAgCe6dACU1FHd6k50+s8qVMv4
1blK3SGCuRbQrylVYJ5RWty8/HOLWxeTuqtnFq/yrVhuUQ9yuCgVZqm16XDwzKy0
dKSO+i3E1cjXRnXnwB1FdfOsaEiXncQ8fKG9OJKrxF/eGut9P0SUOFk9htkwirb9
sd5DZVrx1h+gewuWmX+I2koeCnAcJJmw16JGmXDkKtn6DyLU+Y8Rm8OnrJmdm+0Y
nHEB8bzNe2VNaS54koAcPXsUCH8UUvATNUmRTqBLvaqqu1Qb0q86l36f3xMF48rq
QohqC6HlfZ2r0Rt3fqCC6QZ80zA2zDV/X74qYTkNkYCSHr5on3sydz2r8rtwYao9
8VIJw1h2hR9RQUCimhPjstao0g+ggmTwq6C6ppr9KJ3uvXuMoHGv9pw7N9x0+lLM
cCntfjMwuBVNgQlDGdJNrJdNWutQdLSKU7M52p+vrbvsc6pZDm6ZZaGR3+3ZECAw
/bN8SyXz8XqnpJs11mhtoqKdiyakQdzk2nP5uGnF0tcrMDzHz6/XqKP+VWBpSpzi
XROZOH0HiEpNk0C1WKBW1VkgKoG3wRkVjN+e6SMIPOtBAOBUfl5mSCHAjoV62rSu
SkAvsCYx9gbo9zYElILNhHTEIKlLoa8KW3/wiiam+CAxkMtNaqe97frkgrq03ZBs
gEp9ldZmBiEBzo9/aqG3F5yWo0BWvJ0SMUh8egpcm1zMlqoLYIZEig6HnpbUwb0n
/TCfQSgEDCy41lehiaNLxp8PLlv7sVARNL2t+dyMsKpXqwra5csJlZkZghq/fs0v
eeJE1ZpVaArys1NjJtINCKYz4ie9XJ/s1e4KkcLyW+gJes7i824dw+Ikl3WHJ7zK
3uXJub9lUYQEi5aOPDALC5EdsmigxyC7FR8/GOafUPD1CX2oQhd/JwTI8dILmO26
ay+uAjtz7IeDY/fHww+NUWgByLHegX2DjbeV+QsePqKkhtaQ40+gSAHboT+6bP4B
bY8574MCgchQ2TJTg56lWB8Ly6etBUQpEgZ9QUOx8xkxkuzd/Wu78BKDCPd4x+PX
7CePSH5g7h15fuS/JMiTwL2W6uQgvcOJhvLKtFc1cR3LY9SpEd6k9xXC9k2XQqgs
wotBB/3y41rJ5CBLKhlzdVJz+amfG+s5zEWdwBM725eDvLPkXsa6qeQC3BoB1yxd
8heiGOgD5lJr5m28jliV+mIs26C1/Erk0jh8nKQLeMcP8r0IjKP+7arLEi9CzuKU
1OE0ZS6TaLaexH52au/aZcrMOzaWP+nVyD1kV3Rj3P/GDXmpLlRJwgvvJVf/vHxG
qAd/c5+N4lL1DkFXGAs6pE7B19iafLB2YFfGDhXxdGC0GvkBzVBUHwfGlePF+7vB
rvKtbZuLu92NLoWVJp1BneAw4o+MKwHiqYZa+p2XgljOISNFp5lYA7iKQu5T6aUJ
+DjulWLMT4/fokON2BBn3keHrF+a9vjCbdevrL8pfZe8u8H32+c2qCXviWNx+kqu
hEAtgcNuEQTbKt09DnL0kIIJC4CLj2hiVrGnAVepcqlFEIHyjaPqwQDS3O68CCh8
jqJ5CSR1jC/2GkTTaOvGP7BECzb4jzC3Ntd6MfiHBO5VhJ2WzGIPTBX7TvrcA3O2
f75PDtB/TwpKLNLNWNtUjAQwr9sEojpQkI3v+0v+NMVk9FvHWOdz8cSD3gqWjZqT
1TP0fzZFrYiMwyOBfi5EHxtGvFs7wc6nmCk/WFM+urMj+nw2d5QVJkrHkhijOquk
GADzjaXtnqS6pw/chhPNLSwxAVpshgALtzyXqDEfddT21Uc9xnbBwdV548EXfXeg
hVm6GZIG5aHvaI0ceE90rVYUgaXN0cd75rHdSSPk+FGCZ0BS9ny8uCyHfbzYnX2C
XBrHkK39NccVOFUhRTghLvysjb6S7TVMAB0FaFCwf0F7EVjvoRFXE/VpphK0XuSU
MBrppxt2Cqsg8EyskY31q4xMCtYWsAFHkft4xHDebbj6m93KtJOht5I3uc2PfPT7
+q0jSkwp6caeSBAohpyS8ecFFQ1jN5oePQnbMQBeprj3RmTdEoe8lgmLRE+12zc9
Jsyr5s/i3FloP+wpKyiciBksV2HXxnS5CHl1KhMnRbQNGpwKP4rKs0ltSsZmMdEC
1ndKrooXYIAiZEZM2sEPOTlnQakCxhwGG6geyT+cFy6mSeKXKGSvw3YfQTjFAxg8
yfk59Bbtc9Qf5MQGBdkws5yRUkLEeym/ZKZG7zOLXZ8oVqpBI12ouOEHAEUenEdY
2LX8XP1qqsjT5d0gtsrGWRjRKU3FAo7QqslhdV00vaL8vpd4HKF9nCPMsdv6Ucwp
qBzYbJn7srka/eiulFPz+6/OzhCyI1qFEJG6lX4de70BvVoPveZAoFEbfuKIBoOw
cLK4BwCznvV4Lv2rf7OVua8LS31wPccCNrqiF3vsP8u541lEvg8LrxH1787YLyqT
Pi13R9jo/RE5cHV1/a8/Lk4OGY0h79aWdLJUCiTfgCePHpknMBA30hk1TYeMbih1
mRYIc74fq0hswJZN/SOtnDF8L6i0qdg+IX7zt8ydtpNx+GoQvKD24V3UpjncrnST
ZR7J/xnH8s3+z7V9yAKMkt64F5bUZZCNLmRjO4w1wuTqKGAyepwjWOnKn1qduSFM
yCxWPmQpACpiBpyEV4jB8+KIupWA+r2NGZGmhpWcfI9EGsLoXk/t5cOEtZRCryYk
Akij2MJTERr2V/9MHtIBdU/eiS4Go15b7K60eEyYRwvRzTM0iHJJeuJ5shfOY5pE
7IM1a01VQo9pCB/P6VAPlOKvV8hwua8KYFOVI2eVfhF0lUENmyHVORlEz7XlR+4T
s4Iw9mAiQqCUhIWUW5j5rbjZtpvvG5n4RsLGb+EAiuSnvjrpCTGdx+YUfRJb8hFC
2GPWSqQFdk3D9cU53cYHkAc6nX1+JdhhwSCCZ395nPKSPLKjaUjFS5nyeyNAmFkM
ezzMPe/K+IinSBBlt547m00Dsvnp5tvOvbTKT5eE3wJW2uxrfAaiR2K8L4F/J3VX
Q/debqJN8NqcD6Gf4NvCWcwpRuzkB7u1/KqtnOrFrIIvHEjKcpDtT5H1ekf8KVxt
AvCHQfEsClen5Pq0FvnY1L/8PXp7gtSALqnzdIVyzVBCiTOLTYGSeyz2+illEVcy
o/4WvA8KMi5PBCfAS57YETF80gG+kdBUPP3m/jWNlOEiDqGg7jGIqs4YEF5Ks9yM
z9jynqvUnJjwa2zciOh0bwWJKYpoNqd+4EatuXnD21R8B3KUlRa4EkZpKzu3DBnW
NSZ7Nj2gbZvrWDKd/DQ9Nu3wgQ4Lx93wZ0PjVgfwTEuAM5tDpM5khidBJ6CyZ1OF
S2YgSHsTF93LH7Q8KKsmJ44latZcdiMRpurWQpN4mmyLS8F+GvR1RZASaLYge+43
YHfbtWkF5gYCePZSiwZ22RZijRWNwvkNjPbutD3AGTrAYdeMJxccKErMEbkBCOxw
hmbERYK8wn+9kiZ4RFgfBaB1mbJApoXq+zC3bgpoqo+YDpfGymv+i3WeyVguwngJ
UTXmPLFnSsOI0vip+aRv8HHkDST5e4ZNMxHhW3MswryqM9EID8U5ystSJy9m373W
QRacl++RBQHXP7RwvLHZU2REiQDMGMElXBuq25m0p+EMpX4zJD5MDDSX72RocL1I
1yqgSUwWpKbWwhoyIY21Ms9bsqwoNajbinPVg/XxtTOZCeazIUdzatlpmB2pYZO+
WpHMIBJVzGiiMNJZNARjwxpkabFZZi0prhm6f7/2pui3VpULL1zAVEPIG3rVjKZl
5MOA9uA8MVZedhq4Cw5IOMERowdBkQQRhwP0oU/J7SBGXCeKpj8q9pbLF/msKQx7
aFgSyYKloxP6jd6+xN2+C66Dpkyx7C7SCa1psqo5GEqdDCyh0PDIRgShzBAbZHQq
QNYaYS5aZI/J4/tWWWXoGSYu1BrJG3t51/oLGgBOToSrFcRm9SN9hZlms9suOaPz
SvE1ynaNGGcTMT68hYeT/Q+1lSDZgCnnuHgAE1g+7CbkBvBq9jEZqb2geoQecMbl
yiHApJvY9TIiF5bFeoNP1wdRfN9I6zlHlUjm32qNqYj60EQ4FlMa1q9UeIyyaygv
qzyATiCNfnmCv6JR/lKZUtiAHJHYYyXwBWkKgmSv5rk6e17fXKAeSxVBR63cUcJP
PbjLG4EMY10ysH+PIsVeUASxyNXkCYGbWxHOUFMkDuoJr1LkwRfDOzG23fC0O+rh
bte731dpEdt405czfftzlo0883Sdl/QNWUdR1O1LJ7naWFs/AuQ5tSyL2yvc/idG
zSvvAaUjpRi+drJ9g/ULJb2ghvXC/4XIhUXveqa8WCBIil3+fAKvYrepRmrw270Y
STgh8z9WxDBA3P6un3LO4gHAFKlGImnY4J4YDeyxGQhphD0XcTxtbzYPwokXYu3u
xnVSulaP46OB3m/XMCoXdR7eN3TV/AViH/uib1EKraE2gataDQFd/48nejaeqWT1
cP+kPYEiNiCPLj3ROIZoLkbyWUacQi4kk5RJkYic2GVcgJCVeZvStjMo+NDBZlIQ
oq64m/sjsoQRuWg7uQAaQjw3gKAWquwdg1R9wchMBGheETFpIPVv/1h7o+2SbSFb
9bYzThf4C4YT5ydnCYq8xImsIMwRwYndqzxv56Di04jmb5znw5ZgqgGWsgp+mEpv
5YoIs5MT2Sq/M1Rc8UJenAnVB1Blfn3soV2Ynw3icBZ6gCPwXqBLJINPOauESgMC
vdtwc1lNx92ZCYFu8xjdxVcjow3jKrYK4lW3114rbia8qVrjE47SmVP0AZkqzlvd
QG/easiiutAb+lMKKobzb3egHMnX4+AeO1ppyhNmNtGJYHGNEzBmngtOvMjOK3D2
QySdZKzvLSbIr+cR/vIe8ZTdXprmvtMeRV9X1+rqksA4nqBQWFTSTQy1RHIV6iHX
RK3pMhnHfap6pGzRUrVzPSqYhWq+pf4GO4COelAaymUXRU3z74oKCr4zCSz/+dVM
B2mVTPWFrldz+lqfYGdNHY5b0X4qLUCW9Ud3mg+qqUZ4e5S/kqikRfoO1g2Aeh9C
19B1JvpxIbUrmUE7uaKgd+zBk5d/+8ni0vFbneG/4N4JMpjb59OIEDX33ixqkNdl
4kIN8sqJplin7YxGaJZxoAa6vAIChjaZ21sTtVEnD4p6p/K9+2DfDAVe8wbKWipW
Ths4+KpN62ufncxrcCUEeJn+bScXXpb79beIybhqcRa1OESEYsxeQh4FEGRwd2En
ZWIxgVAR9PXP0joNL9DJrHi+RKNO72pf4a6x07HRqIyWsAADzLIa3Tut+jnJzuhy
vn3UjDwmmZ+gjClnDn7o1EldBeZ1y85tKCcOTUTvEIKD0uT50dCoTBmlfCjKbhno
cn9f2NOJAEvqxAkWK+60WoMfmgfsWilLnblkPdLYAChyRO1rE1O9IZW1JBWPZDHx
p6Zw2u4wPElDEApaS21ygxkivZgqhSbg2+Kbi/to3i4L911Jxu4BpI6Z5LlPGdEq
dRgmqnjPTrf36aMvI+JGMmtU+/p33hh2sInTzvpqcdVifIZOESZCbex2k6Y+eDYk
GPxvVe1jZ9LMb8jc1N07gfSAm9uQOavW/TnrtGknD8HoJDrnnpw74U+D2g+nSiuH
mjHuYD7FppG2M0l+MfWqfpEAw2daG0Ujv5inKVkbS2irVPWyY5ACH+/vM29+VOn/
H2jyPN1bahDSptGXS/wXgBSllqm/Nq10YwCLqEk3nVigyogu5dctyO1lQ4o/58EM
T6xi8nzAAYHLviQMf+YlVtRq3Op6KaVMeNxdsr67VoPA17o7qHfE+aPJMi5+HzzJ
aDnJ7JHOD4jMhjg8rLKZ2hImBU8c0GdJ4mAJtsskZ8DKtm+uvKdaLsfsCQjMkrqF
xnAxTxrKzEPT4/NXD/Zhlfk/ZHYVNpZjLyTLuzAIKHs2v6i7/fdf1DtKs+WCZ233
zRgdsN7yMQsMCQS/TW2AGQV0oGkL/f2E3iKxPb48TXavVa7QJpaRIAfPIOcHnQnn
LrU6rc5xyG58ch/kbKhBSk1qMlAKD+2Im4UtUW9HD7VeaCjWJy7vMRt4gbNyPn0D
/sTMLIsCcyVpBVg+aabduKtuHTpR6kLkHWdcAS46FD8G9V8e4s0N+iTdqDB6tl3O
7oHTwUpgAtmb3/pCaCdcEJ4/LY7PMIkWS3hW/b+y3ULBWZFbK+DokrmZOEl2wQ2S
1qcu14Ys+R+FpqYqwCuX3PW3sXvWAfl+W5UVNYc8ZP8WF9CB4Jpd8/KvYbLRtc+z
p1npbl1pwle/Mx2l0vjRlpq77uK8IKEfL6OHjKcr5P1GqEo0UTj8Va34MbDs4SYD
ststfcuv73TXn4nVECSCxO/TlDxqvlILlOvkEqCe2lilazWZGwPRKHQzjO6I2DQN
2+dUPV0eDr9HionnQFqsSvsxiUJ1XN+UfRJuasa16mNFiedz0VMECCvEmyCE51/r
uFZNbWTnXlANUoXMJy/waPHj+7FB2/4ucXx0YDUZZ+ihV0hv/Nicu1XdHS89xuG/
EavTgtkR39rmoYhhQFalxNre1UkCgUVQ9vDQxBZAvWizNiRfKFtKBRDYj9XC61jG
I8LO3gbwMRc7xvfylNNzSlftebc5YqdQVMoY6Oa4/aguyoUSfPDPkK0ZDV/O70la
HyYGH1M4+c/S9QcUPsRJVu+9ZxRMCctuJGXyrh49lV1DGvxyjyU5oj4vNOWNxHbF
QhPoafftdetmgSZhaMFTJj69MgdCQP2vYhneuByER71JYxsnTE8l5G148OgdQkAh
T9uPmEVM7gH+7UFe1auj0bd3zHN39OnNVVj8b3VN9DLkxFacT96uPDkwmlQnRmPk
8RHOGumPaIAFqtNZQcAPKDF7AGZDEzuvV1jRrMPQJrHk/ZyVaE6W2CGgNWR+eH4W
GkAdsiYYpB75Z8fJlhdOlgw8PqSqrbMibhIgKfFLT8yeI1NRRfLbVrumaFqNgOd+
cYrrd8j/NxX1fMmf+BLrbEs4qpgnpMUoEpeCJyTx7xr1YXmPVLg2SUQtJmHjlvRi
6hVzOIRF3DwHZm5ewn5mY6yPDyiDmGnAOZuhcIu64ILAUcX2K+RehI1XZqx3Dy61
RQ4SUzqaPo1vODImujJMo1ezoBt8r8OYeUsptqOFOBBuvlm2klQJDShBdCmHqJz8
/EQKu2/VDHFPGnufflHvVwVUHvKlP704E4jiX0AU0hg6CLcwd+A9ZJAtFKTKmYTs
wvJeZK1wuE4ncMLrI44lO5juWM2gPr6XxjV4k1F+TkfCtbrcMsueJfz5rRL6Vw4y
JiO5zwZYu+iKz0o+2MUmz7fDUqOjCQT6SJgPsQuXhi2TzsRRyNiFsUjCmVsLi1Mo
7NmecfShsselonvlzkW+ursT3W1pPEmztzNK5DPfR0Lopcj4WQlm3ngyFoBDGVyq
NPZu4WkWViGL1R5M8nP+vmhbVymCi0J3rj5NkQHndaDtkxnC9rTrX1xQFeGXVMIb
KhSTZTLNvla7SoBnLO6zbk2LnvrVKQ0U6CzciT45g2G/73QF1+wevnVhLboqlvwP
IRUkZnmnSu+PSeLeAqS5U+6xBwaMX3aLZD5l4qzn2GG7VwiYPzjS5UCKuWRc2X2R
9GEssFEXizHxXQEalC1kRZYxgi8Fecs4zU4WClUo/09nPVPBGlffCKYg6ginmGJQ
wCCQbSEwp2TTUC8e1rfoDJzFatuCOin0nARxGdMrdCr2+ID4vGcblyXsZIed1ehB
fSKVYuoL4CnTxGrmn1J3Uvwf5AFFrN1aLXXu7C1iTqz7QI5sHnxwmsrXfmUe/Y4I
ulfKmK07mHv7zGPDaGgK+pXIGRJCan1znY74cIsR8a1IDPIHYPRTr10xbwpc6eUg
J+e/J1iOdbVaFS9L/8R8HYQqjQsgDq3uZ1+YKUjXhNzIPuZS/VKaV/JlVCf6jlGl
fj8c522GiEKG87rVBJ2EwfX+quBH9HPJulWBlDOfc4LmsUGmV8m2+bqcX6OjkrJq
N0W+tNPkxhuh138GTWplnLhC6MTE10f0EnaMGEhcgetEGtljJ/W0N5vvY9G7uOt+
eymDCIMNUGSI59yN7Ry3D3cxwFIevd8sfHmjOIAGkAUSVSBxviCikm5EgQnVYH+j
vcPFiSZDusaiSdPXEF1QzCvhM9E7x94OQMzJNbpf3yPmCHU7boWrXd1cLolPIup/
ZmW/IIOTrkrCd5zAGKM60sMQTmmocy6RHFNx5tzqmdgGOkAsu3POKbHZlLPLa0yK
jf7G+X7Bogxh4cHxUmboYXlVhALfqkEkx8DqQXZxW5TRjNYkWCTGZV8KYG2RkID5
oAPF1kGatBS8EQM17TxzM2sIIEqwHM0xXT3sKuOoh8ho7QTSr7PaLic6OQO/HcqD
P6S/EfT39wAilmsLjAwknXcVfPNsO+i7Nnm6Zdzs7y2m6YfsnFxxkkeKp7QlfCmb
HnGwt5oZHro4K3X7/XsG374Ctl5j09NdcB5Kc/eR/fp9hTdqEEtMcFRAgplgR8o2
t+LQsNDEXUPHdNgb2ZUY1UxY59uORHds6Cjyb2Yo/feuUS7yepAQNURFXMbIoq7M
ZbYSR1scoW/oxbD4K4Jz5tYw9q1S6LiiOtIdNV1ajvT7Al2+FUXcH/z3/bZBqY7O
O4czc2qN5y4IYX4ff84xMSxStbNN/pgidxUXMRmHbva2cL5breaLT4rHtvH6aw37
VHWYQLE+nXC/9XVbWiL8U/Ug7tcH9n2sOleVmSL9ZeAufDsxCcIOoybOkBCtpGLc
iXrjFLWFR92NOblCMU3KrZIkPdTw0Go4SUWMdcDCOBgXajOG6piW1ookcgGp3Xh7
K/hEsf8Co+zRmbuv76oSsjMjUsgDC4aWZi/dprGT+hb2Kb5xPXkYKlGttzdFi2oe
ennC/CaMkiwMKlvvEGySiQrGceK3l2/806WAMgZjkTIeNyHhl+6jnZCRedzx3T9M
a0Nu7wrr7B8mW0qroxpStqllbe2ZTlZDDQqdXoumLrg//zfGBwrEDp6HtHBUK/om
ffUEt7wk6uYUO4oqzw14eyQ0VD9U7513keOdN41vJOD4dh15jlau5Cw7QBgVK7F4
zxYiGBKWgu1hBPQsha+WbaEep2qtu2viMWmaHWSxuf6fICMRd7egXNQO2kbfNtLZ
CV0K6N26x7NLIRf8D2Tymp95rziUivMjqF9+LgtuCHjLmwHKD4OINY6AMNdBxrXr
w91OHIfDs1811LBOwwntwTIYk+/kknoYHMYT6jv0L2Jo1Oa5fpxj4xc5KYIRgG1y
FgdaqnMeYpOWptyxWBNuGSN63tzDG4uAmt2PUp9OzLlNRnlaKe7o24pLkJ6sGZ57
zF2G8kvRldlGdsjb5lHUG+/MI50L7F7uZszANpJn4qLowor0ILsFX3eHIoEUcleg
8sXjf1B+ipr7jfe9sIareWlnnMD0ATqMctWed6o8jJCTwtS2wGzaSD0xl3yPcP3W
QYZ2kwoSQTCFOeYoNBaTGSCDhmRZYKjuN5GBQz38E5bQIy+2FPTiDbLc8D1E0IJi
BbgxcY7tymqWzsUff+FDrASsxacPL3P4zzSidVs01HfBOwVnJ/povYw4eZljdTaB
iSTsI9q4AumRwCxk3SKxVyRfPDtHB8R52uOdfHJKsaKsNOWrEY6e9n0PimOe0ehQ
+uKBcUnWjckWWNBDQuwS/0rWKu0OQ0djtuQyM4o92JJLDZaxaM5IKYHC16yRf756
6+vnI8M9H51Lrk6Nrz8jdseCr5/CqhbzFv5lQ9yxhlY+3QZOAL0dIDKcAmetGTis
GP/tyL0vick9Fo4NZnWidIzv1kdAK0kSNoo3dP0OPL3XwrlOCOd0d1dR6ZBkw9dZ
/CG5dp7ALGHWgyJDBFPMEf4BBNSFhAiwyPeLsiKMxC4uEX+VOkUx3UvvpA3I/uCq
h2gbjMtjNzG7lXdsjBDx3WjzD+7Ky8E1WJ8JgfceTMEkNjAnSmR0i4gicykNqfeh
xKvDGVUwFliB3LjhYvDjUhfgbcR3oRwfe6aM/+1AeY1zQUx1BMTLaHRIf9Hm604u
Dlb4+6KJLTF9bZLym7rOIgnE7fC4yX005qZ19nsNr0QvrGB7Qaf3WapilQYR9FzN
XDF7jgrFZi8qNDMJIM1XRrsbebKMcMpP2fvB0bSHJG8AjG25+hXqlLNcYWVfC3JL
V3XEUH51//NTvrWjlNKIQ9i64aCQ7W1b/mjKUvFf3OrKThXsHF9CYRy2Ajn/JAM1
ZNNUQq0XDKT0QtuRx7JpPay798S4az47MRloT8jmrTaxrMRoniUAyTpuUscKirF/
vtGYCMjyXGsSX6SSfxm9d74X0+j+PI0x2oz8W6zWczHXRcgkPCj+rD/Yk4uV2Qeh
Mk1n3TqRcI7Yld2MpUdpVsQVj5pl88Jn1hUgggT1Fbu7RRfPy2l8syzxS9pP75Me
PiFNd/XA+gsUy/xf9FjQ6PbRmH2LD8+gPzWyBr+P30MFMRFDozx+c38xZC4nVr2M
Lnai/CU05uLvZng/p+pEqFfmqi1SRREmmIvGlLLXteS1y4SCBhXj0qyCSKsXNXXX
f9MMHFHnzKn/a4oXCth3g+9wEsMbbOoAwA7uE5CPHv/KBIgxGbG0ti+ZezcIbAhV
hqPglIK7UDp06iSxJBQADZ4CDGkXHlv3wfm4vWhLJLiHwWHxWUNduN0Sejlcfpg+
D9grZdYTLhLT5Bo47XCmz8GXRrTiz4NicxK43crUSG7TvNL+xfyETvisISHq/vHh
3g5cNaDrgRvm4+T+fWwug/3RescICl8rSn2WEzSreEtGArElTAi5dRKYZbWOAjXT
rcyzi/DeZ2rbZqxkqtBnWNrVImyirLW4b0UBZ9EdOrc+yHQqZ4BucwCgon3Y3V6d
dp4+rDBQl24FSAfC7IGKvl4myId6au3/ivHhztNEJlZSiJDij6Gewh+E8rYp4xKQ
gEyGpWt15xKSjL7YYzIFLC0kpriYNCO7PqH/KqzFZtwFUq3ER67W/fMHXkvHqwTq
I2oDsIpkTChLFrq9szamuyP4Fb3fgbeo9XFDHs5TA0NPN0KOfMGHrxR/NkgFSo0C
Fte2ZfDOmod1RiYcfT1JPGMy7/fnWnopAQMATWjjILcdkmeM/jW8cK/qwK14kCRx
44JKCo4WGhUTr+6Y8PLclutOGDM2FPmr2hSU22mg5O9DfVDurMsZ/ebjzPvnYSZM
AFjZSdwad7JYYPO++IRKRxQkY5xMpBOyZ7bdm9+FMCDBli/n5ekQYkpgTzzrru1p
41DphdXakl7R5iucq1E8qsjsst8/lZSkLyXFtr6m+2zRTHEAZFw6R+zUuBCjTt8G
74lTQMLQbN0qU29GXBvU7QiH8gIWDBtE2ZpCHY+6WNeWvcAYXLTda4aPsXR0Pn+z
kjg3UNkVAfEMKCj6MzB33MxIwEFS8RNxRYtIIy6DjEFgPo1FU25Z5GffG/drX2hz
ebKZ7es6iiX3PLYlHMzDo1kZCQasb1d9x6D8OIXsWqlJHbsDKdq2Wl4/1dBEvTOp
6YlJFCqd+HEmzQGBxwH/PiltbwUNUzVAvMofuLn8WvWg28+IL56Ez+XNvHR4+kbs
lVAcb23Ow3Gq4MUi/vasjeeBeB1rBmS1hxkuw66e1wXQHdb50RIvOtGOPXrLMclD
FNfS3AS/ylmV0AQm+ywrNvFizvUHKAu4/dQvYnRZVLa0PLWW5Uoq5nYUyghU6o4T
s8DyIdkMZ5sp081/Lflg6Mmijf4RdEog5rJb4PXmH0L+nLX+zzv8PQ0UKeEnr/nA
RAAlDj24FVMpSHB2cImdmZ8nWE2z29p/ew4sV/EJTHx3IEEUJif9QFs+CrD/dOEE
iJpyF9ofv4tSraJwBfbZJv6sCRBpGz1U9JE0GE1Y/YAM68yrEMNTvn4+H9p/qqTo
U+GfPL1XRSyY+OJxP0AfcNj5WvgKLxwa2Ph6a5qKlhKVir59ZgfflofbiecoGNzC
wtZqUZCc2+q0l1TX0I38yJqIOGEdpJE5/VwXlv9PuZXPktmbmWa1VJWq0Xm1L814
SzFqldJWDoh1d3WNJno7TeDPqQfJgJOMTpdUmCJl3F0oLkM6YXuradeoAkY1v/lk
vwksONtVIE+6FFlDo0GyD77pjvFt7MbqhGuw3YO0vOnAlY2KHzxxUjI71//tMaZQ
tzKV43HyDNMWOkgK3HtQUrKCX5IYw1WEZUdwunhc2sJ6B6JQQRDSGs0PSxhaztoI
uMLKOzbMv/0GHlIi/Yl3sttoPBFeLy9/un/EOZz/wLSlK1S70aLZek1Ejatl2XsP
ic3LVwNhUHGtKkQd5nir8Knby6XjfjggZD2B70ImY7UojeBLLX+AofBArM7VJahx
tjl1q20m8VsCALfadHDcst6DKUbVPhZ6g19A6KNOe9EMUbpBuGFoZI9kxdlexZcY
LyBSyv6BDwudDX4P5H4NMnyucuYkLDK1zbdHxrgciZ6Fn9woqXly5Pu0LESyC2ZL
KdxJu7QUYvYDHbtd9xO1ofhCLyGvNWNt9xG2h/L6LLqmbqyWJLiPLaslcE2ThUs/
LNdrPU/qLQ292ldU3atBtYUTM6qDcolloZ8D23p8nZeu0GIih8LBSgc9BQ8l1tP9
K9DSmHzXJ0H8XvU7zeI3sL+VmV8lNWgHydMZg1ywexX7LDpKTyFQkABn1g/7aZJG
ingCGdFUasuZ/u64lQKAbxVGuEBIRddxPy0KWHvnXLhRfH72Ck4ouV7G7LlbA76d
GbABVcT2H8kto37KGdc+1K/Kb3XIdqUa1yamifTshXguOw7EZ1FgGGOwNS/0bHI1
bWbphsflTuvXsbuALJv5pxfE3IszlYDX1MYUF9cM4bj+SM2GbPs+Qv0m/0j7b99y
Vcp4oMVIJRTUjmy4zIc/p30HvY1chYSybp8piRwblMEpXUyTpuK5jxAIC+9o74bu
cNcrf51PGWUqttkH197vCxteGBWBdfYSG6GicFMdx+JZrKWE2FBuJaiBN5ginzgA
IgLSMkP3YXZh2rUEOCvYcj+xeMyVPDFcqN9wubQO7zdh15c1up234nQy1nehkuYa
Ozc7XtJ+OlYpUrkwniyMgUAuMhT3GZDEaIG3CdZDZstLeOtLu1hpc6CWyYOg8dIV
3d+NUXQg6YimOIg2u1phrE7mMkTkN1JZHKAGzIyMubgbXYJjT2QCjgVCMPYG5Ewn
fVD41UQJEt8diofpoAdKkjiBgLwTzSYW6SVvHDQ8hUeCEdANLFuyhnZPcsPsxAs7
AHk6BiCZ6QfPCsIDm6EhCZq081wWVY1dyeilteCSZcgRJKOd8npKfHo89KdNVZQk
LsbZlpPa+Q0X4ZCJeF635RWf1eEMuAGVyqFI6LBOuXbCKfMCcYWlAEw+2bOCl+2y
bHjIPb/q+86rfPrQnHgZt/NI2j+hliE4vGfMWfVlm9NkJUB8q1g6DnE0FFph1rrO
JuC6axfbVIvYeLCPwGG2K1PIvXPfJkVOvhWfMfQujng5Gs8jr2Ya7StaV1WwS+JW
9dBCAEC5WTkMqp+y8nPT7YiQqb2uWbtItbFTkW6GviCiY/xzv83+NxGQ76HXMBft
xJMdf0JH0oU+cO1IYrKWYdIfH3JG+qZC2pFkIu1LiT/MgjZSvdUD5VjsRT0GuBFU
bKscKjtEGEp/JkWaPGwd45z8UP/LQAOZsC8jdvxILm+9hnYjYIMk+zfS7mSHEaIG
eqVxb/T84bKaRu3vlHhnxcW7koH1ONVDqORe6PvRsc2RfnmrooO7PNOcyc5hN0Pc
pgAqGndVtv8XK0vjGy7PPuWVXMu10V/WvlWFmEWdfB2OHxTT2E7BrAC8cDL0RDIJ
qlAckLZO9V5c0R3/GdXVTLi1YWn/HYLbI2SpM6GuTsiVxIH9HuIvbtRAgzrlHV9H
1+Tf3jkyuQXUqUGdjPjs2hJP6+tgJKMb/vdmr/em/0s776rumyUPr7ngEn3lMcdx
H0o68uYOXaW3UR+11+/QAdrkxnE3E6I0RtwJXZLLMGCUeu4zHsdZikP2MCdo9c3p
U9qAAZYAapMeInHBTTz9Uaw5PBGIUPPopcoFh16h7mit5bW1esfXDvqqGzHn/Tnn
u6pqfChSvUfl3ETfwzez1lAYM8xUgEMoAf2gkAJZ5IKzeGAQQc6Vd2D1VDGcJK+8
me0zys9Iy4C73YJVgx7CAGnPTB7TuOsYtR1r/uEDDiP8qni8kYdLntw3cRvA3Djj
T5WwbQC9uQfHfGK1nxMUR8kE4gdlDgpLeDV9VXv1t62IkzPlZQBVPEpf50o/bfh7
Vu5n9mtX6j2Q8+Ob6d3yWgoo6R/yRZ4WbzkXBIvM73RVmoQ67hBavGG243dqK8M7
3kmxTEuYHP76VQcqav5BlWjihEnc7ECB3Ra34SQ/DXSDFwbap0K7EoiqbO7k/MQm
F8PzKEZ63ACyBQxvrf1sj2ECE2m69K7sOnkDpoQBMqkQmWwjwkIOiAY7SnOnRhlx
KE3xdEAPnxyjoj0AsXvrGyCY+uKdc7lqH7hGLW3OiV+SYJShxq7BHhPzUeO99TT4
HtOHzkgAVj1w2XzRlFzd1tCxXZnMnt3mj4H3oZcJCcflDYOR+KJGfPmd1xa4OfrY
hg/wR28YgdSczGBFqheXLvo3LT9o2ZgorRm9FCgHshq2ZLWCG+l0Xu9ePHxKfDNs
IiAd4vrBj4qpPVTVzByCvLPEuXyoCinJUJWIGsN1ijfF1o9F2fJniElw5nb1yNeB
Vr8n2MoXulCIMy+czVH3M9Jau7Ds4h5pAdmvfAwq7Ds3JGDKV20anr0qCt24DkUB
b1NiH3xh7LhrigOUrxvF3UUCaxAUe5qjX3Fc+mjfPzDwFu1zGtvbIRshcw/vsBFh
lx75ivFJNKajpD4ActzA2MvZPtG2AuN4XdWF3WRS4a7Dzvcr9vBmrUUa84wvRpWY
vV5cD09iH14A65XoapmhcOLn5why7Tr25SvB6MFsRKmzlVG9EKJ/Ne84gae7qS7i
DXTpagFw3riRNgdlA24XP84GBjROHmx1dMknryZvvoaGHyKwIA5fnRSQfFHCEOpU
N3evlSdspWzDaxwdPuuZZcA/HG1ezKIahblTOODqZpFrEVKeLpfczyEbyZ7arYr5
2UcmH6ahwnUPchF0Qj1eGKuiy8wRdfeoDGzquslgX7chdbixA0AAyRYBqpbIACbo
1zRqo0NXPPcoJal7RHPDGnaY1sA9Tc+kULUJ1i7aopcs4oFIbsrnnIBQ3ahIzQGY
9PIZb3fEdy0tfHoL8zXLRri9LgqqZMvq4o/OaHrwn01eUBzi/axsKbI6jZg/4Vz/
kd7qaQXGkwajaIaWpu2hi6ImsnAAqFA0TvRGbyihOBUEyk5FyV6/V+rRKdoTOpV+
szhvORlDuAKKm44OqVf9mQ+S1D2MIEkBlfCOZ3ZyFRz21DMS1hgXs6KVA+aih+Z4
fZQ4elpDlvOGo6bNPTkAwaMKvHQLJtaE4FY/bcciGOGjU65n9tQdpFSlGt4Eqz6z
UpZVejtUBnpzY2+IICbRNgdLDu7KoiWu8L9nUTZk9UGK3CKmj1mlciWkb7qji2du
UHUKXkTI/CN4f3fWbGbY20dRsaTEqiLvLcsIBOjW44A7MFs+WOtygcIOSjdSyTVy
ekh6D6d2HECbcFsbk5//uYcHhDzlSerehhTuwCB3lIfkf0WAs/Thmy8tjx9Vw9qm
P4GTPzIYNuckol9HANzPcb1nh/U+5Fl54V2fooASAsW1uXiu2tg6xetNm4yOYlhM
lmWF5P3jsc3+xUnT9DMJDOhNXpxPgjP/+ii9N9tEzoTtO7uRrBG2jbvAc4+4uteh
U9MEjWiaFLg8VMeOhhcklziVTcAjgHFkhUk3pNf9DZB6ugOgj4gecmhxG1fSHEzL
RtAg7QYbgLk9+BLYmExiXiraJx46igDLUJSTYLoWHkvQgySRjxD37imP/+eteEMV
AOAr37zDjERFbu8AwegYLVzxntrXnpF8Lf/aza6r1E439Rk7Abdmz80SjLgmRJMs
wCFOXRj7qjOh8COqjVHaOdxxeDZa+7xCf222awV2b0rdxE9eOKiZovKIQKMpPDLT
b+G7JCGw7NVXIHBxy3jKZtSkY7VTGctKYxIbbJSWSl+GD7HrE7ZRwOmtQuzAPppw
2E2vO3hkI/bkYUUA/dc45g62Qnt/oy6CObaJ1iqVYBe4XpfaTgiQsJNaMclmC7++
PyuQfc4Na7MOnW/bNPd/9FLPHAoNFQRvaoP+ZIDo18VMtSL5Z2V3yDRnOWIFN4V1
/4RPYg6scEp+sVYgDpubnd9Sv3biBuNow3BnouktMgpU+AfRvxQLvG61V4z1OYsG
ub9HJ8otQXH2tPkMIN/43/9vsIAZJ1EUbgWs8tGKor9huRP6SuZk+zzUdNqTAef5
il0PMnHDr9N9BlsjV7Q8XtJHpnMdiKbxr5C0ewNpuzS0MzVzEUyoKUw7qHI1WXQD
cMYXOdpxubDhwrmc7Ile2S1PzG2kK0QiPpixk68qeplKjxXBwleAsjTS/oAqD0N4
Ye1ihAdYmrSuvzngzo4Hn191DSo5G4dMe4zmkJ7vvbr8UGY4A4DHVHKOgge41WC6
ZtWWWpFZESm9hygGMe5OnnJ5wXUfliPKvgHoTGpuy6GFa/WG6m2FxuaaM4ZvQAn2
dOFCVtp9l5IYbzQFlQ+Bj2BT+1Baa9/miqzQkn6QPpLKXZLHEZQvy2MEUR1Qi2U5
7HxbEXIVsg7lDdA/MVePLgqlSxOLhKKQLUE47KvCh4q7wVyjUyfaabJL1Uz39c9Q
uGSVIJbH0aoL3ss6MSOoabi8WWDGELEOLZV3JglG354omwhX6Tbggka7uMn/pLF1
vYj45GBTnN/+u06EoblmcFA+8Q+eFFG8trG7IoumsEn2idPdyUjBCJ0uO4mq4Gce
kC9Nhz8ieQmwzRJqsCbVlKAJqNc8lgdeKBSqXs0moW4j151RjOpVmSR8zxqfP1db
XOUSGzDETpMQ3cHsb9kP9jBOel/IOgm7x79nYboeLKAE1cH1/tlWOenv82M6m9Tw
y0ttp0xKmG24oBDVKchJXnV6/u9DCv/IdB6Qi/Q3E4nqD21ze1Oonl7mbksnRgPD
StNqkfq3Mup7OxBHU41sSJhVTK5KULjqq3PFxW5XxCYd47edJBH5giaIyxriwW/V
LUsS1UQ+QFAh+ySpuK/NJ/QJ4GVAmGgTXYjkCoB7EfaWs2SWIj8CA9woj1YkON5B
YQ6vbDUpUc5+SUeXpn0enFenWXLABzd9q/M1WuBPThAImGM7jnCxO5oFKsJ3uHcd
DpVDex34CwJGBOwmjQIb9yLb3nEZRnjpk8qLSbSHLHG+wbFjO6OJUPrpu/H2uj5o
cwBdy2q4aqMsrKEJLAXo3afo3lpFM7mz8qNqMUPHwdiRagfZC6YEQkq5NrkEKf4t
M1QRMEIfTOnbMah7ljw4TeE5HY1KE0SirR7zo68q9lNP8RY883V63ym4AnJrQzR/
qvUtsy21hcFIfJs2Dc9TDIkSNcnHosMx1rjOvnDbonlG0PFDnn6GvNLkrXsOcq9G
Ej5p8BKSwHYHrzG+8VJHNc+5pMMZncJKp+8EOwEPDv45+5JLFgliE7E2t22kUHu8
AcvN19+Br+clzO3brSp89gvpl6o7PcwnXTX5kfjqm+hrQ+TsCxlSy/ZvKon5bsdK
FhvuRInOwXVHsQvNAFqlp/CPESftmL3gd5in6woYwxLSNGJcoOzH9ZLi72o7XUyf
8Tq97/68WHBEgGYaZ1LuQ2hXYwEVTcetj49Y19D3B6ZSAIR790wNI0w1xD0GAo9F
NOAcROKCH/QjRdbJibwb2246QSeEAITrTMPK+ZRaQFwL36Kd3s20DmRzpXVY9rA8
pIuydlRjfm01cPAV1Vh9Hw2cuzORP28/Ue5LI28+Al3uGNqftwC0T6HvS5uD/u3a
QbDcdto33Wwk1iUMG8azfdP2HVmueT4czDnC9C/8C++Z/25yMW+Eop0rTYOLKpTD
0xQM5routqrfLznhKysrTdqa+4xc1ydQRhO4diJm2QzdxDQ6RIVFVNoO0nKoQb9X
SSjgQ0wvkPQyeUBTXd6LaTdMvYIAh96h6nvdikTy2S0dIHzx5yQCHvuNmaPD3FLO
iv4W6zbf4JBFbEceUasTCR4znV7Pe77GCJzfHmDLwRm2t/bgKne7yUx7IRW6qW4j
rv8ynHU+rcH9paDHvVUowXQotnHcz7VyOT3q34Wm7RNGjDlJyugG+LhB54drIBf5
WnuJnUT+tKteqGALkS0JJvS8ErQRH9CDL7u4D2vI3bFYGQPe8DPYktNZKxG3hbpC
dJgn+Jhf43bxS1LN0JZG24j0+Cx9ZbRgDZKBc+sqgyQ79ukeiih0GSLxBT7AB4oi
6aqT1VyUfAktTnFAaCD22ZY9u9q8gu8/sp69dsst927/JGp1swCBeMwYlMqcqi5z
l05cJSm2pptc/U+pbmHorBkP+Rc2Dn+ec6L4dJxSb7gz+cC2wOFTj1WVjg5kWmgA
jFgI/GhYfr7uQPzbIIYIBv4nRKDMobfnYxjc8IoywieKsbBeSjdObFe4MJ+08BNm
xbWrdQ11rk0WxHEYXEUzJ2oGeO2l065uDFyzHTPlsDFwz8qbXSuzi5pMYqidtfJM
a1GLi92BuaAtpbBjaN7rvCk9COXEdhOGs1M9+a+OW2LAH4Y7/cUyIbnuN+DuRwgL
rpAVm/isjyS/MFYCI4GJWXD91DY98Dq2EgbkKd5JmxcbPr0W5Vpzsem2fkTkdoip
WroNYxlV2SiwTUgCw1/ExTHCpI4keDDCKy+mRnVmA3NfIE1kDotUeH4/cbdumSoX
iEOW5O4dxWsJk5WvwYn8UdpjtjCSsV+42NvH0txnycLOF9ySD7+jsSntrvYnWclX
ukOU45y7GIE2Rhq3ySq4Nh5kCZlT1vLnlvv4zjYFk++TLjf6WPGbvSqrNovQZSbM
CpO6oYgeu5PDgwDbVV9eKyxpZigz9rC3pS0ADh0kQzmMZxLHrIb76xpRn9Fj802R
HKrFlXgfgEqr49IHcTmTy2G7ogO5MgjuMGdLOFODM7reW56fXRgUivKEd8Xa/QBs
JK246pqUsWRhM9y0wriUETJOu38Cu/pNR+ftfhokgK8T0+6H+gFXlSkkqmbyq/BP
IQOvdckSAAVcXDn3yq1BUSYGy/HYPQ+Cu35TgF9oBINdWURud//xEttu7WEN0djR
YxiPC6kKwnw2PY/h5KGpiC3gxpmqQMJEBv5/zvPobsqX1EiUlBLQ0zyxw0FRjofJ
3jmwwPoCxN/XTO6j3sV4lBGjzGiw2KyzUiEVrE7RLhuSsojglbeLkZ8AN/Aj7prn
wA/xJILfkjPoEc1TaTxF2tghqMYgqiDzvoPQTEXIIEnYg3NGRllonLLdzqOWgkul
yalfXomvpF65UBP6HmCzKXtp+XKfs2q0T3JQefZXymL9WoAJqlwv+qcfFgsjFSTa
6FWiKHSImvXAgd7MgHAyl5VIKsI08fumIZU/BLPf3dS773DTCd21TTGzWKXn+zm2
1W2hS8dHma3gtm4QhX4qx7nmZjYVtoTNDpPymFXdopbr885LRWzbQ51MP+N/kVaQ
gP2mSgXGBzpTk26Mz+T6SO+qOmzXz7xtdaxDrpJZIcw2buAQDjcGP8yGNzFJ5wfE
q+NW6Asupe79e67xSttjkkVQhD9Mq3CU6EFv/gZFhTSp7wYe687BYE06XoF+MP7y
Eb/j+YE6JpliFbCwn+aGByq8IZ+a4cg4sU82re30PWAzPrOt/rlQZy7ONdjUEelO
QjMh8uPpP9B0l2fZH9BvCaFEHypTQC8TJiUdKzI0cAWGtmOEE7SULb7DAqQfOfhn
6bMhBEsKgw3gjdulWQ9aznR1nz/lBFPs3VBu+2Z4SjqHQBdZnrFt9P4Lr2swoaP8
/i2J0oKiWAROagscWQpmrluQB49wVowjOLLvlzKd7nvRJzsFsbWw2Extzb6Ywyky
kxp/uUeFQxU5Dzrw4ZLcOcBvt0at3DmiXIBvoXkpRFW7i92qro3WhaHtsMIaSTqF
CnbVckyXf8ICsF6IghHtTH5UJ9j+sliRdx1DyQC4YfqhtVWyIeA15X/sm5eHrceD
K9sRJoh29wRmd8U8914KbTsXi54TvnAp6AO1MJtjHWce9IPbkbzdTAbyjLEFZBL0
vBmzSBIL2Je4ng1vkzA+45L9qYC9cyLX82711uc10+70bNYfG4F0ZWwAyHHZ4wV/
4TZwMgXmK5E8MC5+ovE4I36LjLJk8t6/24zil15h6a3xUHVyTIG36jzAHRYfHKuX
c7s6ox4bJEY9Qj8u3yaFq2JdGrmFo0rMLLVOay3szWDHcnlXfpeHjHIn/ycsHiBm
oZ0VZosr4ba3N1wHwSXaevrZ6oC+JkevRzubGMvVjwtnwbWFxb0pXXe/kyY8gUmi
cfJTs93aaVPacPNVOJ/0ME7mJo7Bo+Jf/CiCh/8Fhd9LAahUjLIIlIxk87Wlcl4D
BoJlsREUACj5OGKDKo7PxKbVy4K9iInDHikZngLMW763tPD15pag6sIcV8aYJ7sB
OhGME0XK5k8Kr1jW4Vh4X7+fsN7u4Gz2UMM2jhkMwdQ+XMsrgQCHU4/vnkDug3NQ
+Px6XFjcOYVJYnImz9ofpqiXlVGSdtWoCBLXqWD/KP0VYshZ4/aMyQ3EYrXM57mv
sb+pkPSSUqA6aW+45fQy/gB0dnoZUkaO1p92a1s38gn5ALyAJjY6X58PvLF/wCxY
IHn5MPTPNUO+T/3h7IJcl+ZEQQYR3BU0zJW538VSfaJIZ9YahSSJeqlT8i+iuZll
AwTOVCup3gNZkfkLOOxkr1w6BQvS2qgFC1a5daRWBkWhW0JfvIRZVTG5IKbEEQcu
WgQTR2Wo339W0wT1wudKQNxNZ53MTex3rZf2XKmVBmsf9MBirlNya6RWsJIaS5jn
oY4Giye2U8NDC+T8vl7cGGmRqgnHON7BQwRD35AaSWP2Y3+BVyJEZ3BKwczPIeV2
ADtZqCRHZPOrXQthYXI15kJ6t2k3coE2aY3h6DAFflkyRkYVdteZwZZ6FlBOGcxu
W71wUzuUUzOfn9Qt78U36X4vY9d9FMWaNZ60dAbNVV5m1hPK1DQY4KSAhWXy9lEl
g2ABgnlQZ5T5b3qRkq1BjYGr8tXU/eRx1A8AYW/LeOXJd/jJQFW7funfkCp56Yyv
z7WPNbRcWJAPli2NTmUlMxUbvocU6+k53RA3Jq9R3gfzHpfINp4KjwmhvtTQKA1k
x38aVBfmYH0t9H7DKlm7cbtA3ouGlo9WxN/c7JSYnxvTYDdlMNnTsaK0Un72HIs+
RTDiv1zmF70iLnzWe99dvvDdIJ4BAI7JBGb9ebZ2U7bh7MSnXzT1xYkF8+v4xN4h
P98doTG1xPrp2ukmdZpWyRLa+sWAnovygix1oXaiET3+f8Sua2MLmwjxdEytuEBq
5MgcwgEttjiobNf/UbTEBbgf86JZHEWNky72gGnTO00JuiIfuWd5Qr4+3BzwonFC
qJngNuweQwz30n8oGyHzm30CAKBnQ81unU8FH1c/Cd30VoyaTbOmlEPS26CGNdIQ
qPYvYB7Pi7ebCelKNTRexZcZuof3b62t/aF2GSqCf5YxtPfskfhFGE3A83E573dW
mB/JOPUjJeQWHmBsIsi8pXAQqQjFIDJU/wtGgLapHPC82ygOVhctWGubSY68NJEe
9RSOXYYXhlBLuK6NEh0NPaHb4xF/EBj90IkUUgMVIQmKWqEMw3FcG5RETkVABgMs
cJRwJYWw8i10jfOvS2Hjq0ZtXKCRP5dXxwrN5S0Kxsf217WiMfEzYrJZww0ndW3U
Xd802/+IdjPONLlWBehENMus6V4UbJql09SJfjzg6tS2oaaPas5FNvuz5GgefmCx
oeyI0BYvUtE7tH33ywA8BGranzmxVxCEtrfAbVDiDaomw2P9gkCzPrpdmTxjKsoW
dh1NUUEGL+c4eJOogUQUm7nDXl0gi6PclVIMnhxRs4CnGpU4xnSnrCE6kTEPF5MK
nftPNAN8FNXH4ogEgvmIf+6Or1ZzJSJjyU32Fe/UUfjhpFQwDFORXMJDE9ARuHWo
9L46yt457b2aj6C0nvhQJkszMibR7ECFsf+HdNcAl1Gi3c0ktuinqtYJ/6jZr8Zr
o0eF+pK4ltzSeQpozVSeObRxytysdH2i1c5p23ULAyWziQ+IbQXLys1Je6LQL5Yx
HxEd1MDgw8xZN/b3fMjANZwLFmjF3o5zq7XSIgBtkwIObS46AASO7sU6wYgThIaD
KsmW/j/p9hGFQTF3o1kSYeGFvnPFvrwPXW7+GM7Bz+7L5apw/O4voDQ1qChv7Mcj
d0IG8j3EjqndMRL3R1WoECadv1qbRw66iXPamviXEk2yl7b2czxHqs5n9rcnrvAq
p+QtktX7jQ3k6fvuKjTpHtVAGUFDV05KC5sLuWhzCRZU7nmdwuU1iex1gXns+R55
gC+hOs1JaBeNbeDua/DE1GtEX7wDw+QiaI3pBucJnVRURe7owFfpjleRcLIVnWWs
zzk1d7baH3RS/fp5kCX0G4MyzrwRNeic1VAsB6D0SIgLtaNj3i0RnNWeGtWnqpYx
DoMDRKTpRJx5MNyZtfoiSBaJ1+0EWWR/vlZuCADLKafXzuhy3fQJPmht6dGjlvqw
QxuuxKCCjBRNqal2nNJuTFeO0iKIC1gOohrJKXK77yjHfytfO6hvboCUPZwx2Hp/
Ep3CYUm29vLPl9B58e+Lz9sjk13hFwbB1InXik4QBZcLqyhqoJ3eOBTCHohNsPWo
upd8+ZAsY802r7PRAq3h2mYRUFx8izxh15AbmX97o63XtCIsC7aGRQvBAxA7PJlC
03T+sQBaBleM10pTP5+BvPf0wN0xyE31FtZg3oaxEehWcNjZ/0+4o7R8ZGRUiBhb
cJTKuzyopfVc1afneeuTgE811l3NNFD/yKtKnUmMkCMin5EbX67Q4lmLNfosIM04
GeUDzib639KLtuxV+K35M68xHJtx7ezW/9utdmgsqzuCrU1BEXPqC02yEv7hoOFB
a4SFjQYcoJP7a07uu1GHHTWClZdVeNNom0gO7VnhSXX5FOOdv1rs5wpKuRVXqCN4
SWPNuOAsq6M4bdazKWORiV1tlD7lyYL+GC2h+HOSKZgUiqOurOsHRcIeLo3GSYPR
uyv+REh84dUJEKs/nsXyjo4x3HA/hSy/efZ2qaH86CrQIJ9SRYVeyZjPXzr+NB3I
xsh+kuUzw+USNktjRVmYqIqMRI6NjJck2MpPvC4OPBjlO9v/KRh3jFbHlkB59vEp
sY1q87exDk5SF2UlzjVfBqeM4kSLHT9xMlC23cUhDuY5/WzNNQuk7BuDpFpwyqwB
Xp8mU34216LCZsP2IiMsatpBUW1k1+sXct8Dkqu8H3V8uCQSbUj9ly97X+Oc+Q77
/hB9jrhDS4XbBJvHWi7KaN7vapE9WlZJJzr3L1rEVoeXc9XZhaxe5E7hi4HJrjm+
STaEYBzO8HkpmWUSvE1mPVS0g7IBdmrXY/4JCFsVeF0hq4J31W6nTMPB3zeiiCou
aWBX4+DgoctjV2Lj3tdVSHEd82gRMGaZ6Teq+1bCvZagj2W0JNQxnv5wwz72TTjo
91sQFsBBXl+sa49cS2a15LmjgQ6aqE1PDyOn5yT4bh566O2N6cJrQ1wZzaMHTpyV
FR18Z8ukSzavhaevnHmATGRjD5ZXZW9WNuLF4Bg6goVkZlGBSk3b+MykkqAonL3J
dC6He3T7TPauA/aWSGdwRcWJ4BXKnen5rpp3c+gikV6Fu4Mo6LV3qMR5u/hZs4Ve
ukyHPSQjruUVZzyD/f7wWV3GdYobIvXekVzaOoTuIh5NBJyGa2mFg7CX2VhcK95f
2DzE6LmlDbqEO5PUcIOHiMSQ8wo3sLAMPrQhF3m5SIpmRFiHtfjtjY4lO4YHsq6D
0SaafjrJMTpQCnJjelfBbs+6Io2xvxre85fovwqntBv8Jzz4Au3NlkiJapu//eVQ
t4iQN+aDMAD77GycsJJUe+igQpDU4e1uKUiYofHJ7ZoMm9BTQ8UAUR6bcwILw3F0
yYQ/utEmnKGiof1rFuuyIDlAPxm84bziUJyHfksA9EjRv850DmDG5yHR/Tu8Atbi
Yvk4lr36Ife3St7O03TXQnWi3M0W2BzWFeFiPSYeL41fvOCih7gGJWNG5P9mCPoF
fMiCyVe8eb7K9vdON+401wo5t9n8OhvzZ0bRlTiCHV5vUPAkniBRK1HAD5gIm7R5
TuYthSZQ1fKBNWsLxA1HppK2uP5PE/YF3jNqOAG9fk5Fx/33IEjKBlwra57914LS
x4VqsgOZBBVYxtHed0zRNufnJInqaF6qSzokMmkBwINbISYCfJuDGw+SY76OOHFw
XBv3OhIXK4n/lRlkvwj678XI0dA06GHJiAHi5dzalF8tCFUysWsymEV6lnyrvjue
RK4pbXbkp+Z+fXNZ0wJMdwDm9tEFgj26EAQ/7syyOdDX6ORdHk/AvAwAsFVwWigl
rT887k+m5MVws5qI6g2bXcSTtl9SJAJQcdbhLbtvwCE3dE4qoA2QCjQh1k0DPRuX
IaAB4u+iUCEW3vLc0YL8LO3jWkzcxuT0R795l/BxCe9IqkSO+4cQapMBNg+e/+Qp
o4mHEkaiEporUpJhZuYzn9BVL8EU6ctm6uu08ipBrlJNZJFLRYBKuLlx1A55kc7v
5W9Dc3b5LXkqp8U4BI7U6L3eIkg8TgsMMd+wWxtw/eWSLckSHNs9YkUcjmiF1nXg
u1r9NklgbeqkkPDT+guSuSzRnhM7UKzkTDRtF+BYtLd0iqR+6acK1JGeNXCiK6NR
bA4e62HdXpM3mkYaDAWdpfGr3OW5nMcbrqxtFkoLtZG5JLi4YViNyrKCiFMfsAd4
qN2zo7IW+7pCVgyVpsghNp/HtDD9X3pJEC+d65OSEwitxrcULc2k5ozYnmJUCFfr
hOCx8mLC3XPuPRn/LtKowTFQc7bQDjhP0nl3dbb7UAKHQTTH3C/FWIINm3Je4GXH
Wegq7589FTJZJyq1mJD6U9rvN9JMBKCBd/TqjKWlBFQ8Xyv5Yq+ZqecL+EZSV/VP
GCPC3W1PEvAQAUz9wiQYevFGUj7tRL9DUPtbZjxLWaUegTNkCLeL+ZCbo5vggc3r
WwD3aOycyFbozmHNONSR1R7mLQpgA25u2ehXtn3H2j1TpUmC2f5dR+7P8wiV890e
u8cVjoXrHupE2tBumFuQTEXl6MGyHwa+JgWXSaHhv2D4xblsjFEKKLOojWY5NmnL
sOtyp2zOA+M4culUSGbNx0PG2zFXxRduK2uaNGj6Mo9ae/qPyKtwv7aTY0nD7PEJ
FX5OOXQtB50AE+pmqtj2jhbJ8ZTpXIUmZIxdqMzAl4lr+vqzt8vw1KVA8V6h2ADv
0egsO5dGIXTF0Ve7z3gSPlaYpsfURwI096S9yKFeZAjPMVkw3Cgyz/vHFl8KHqLX
R0jtnHIfGFR4GkNkdLoVEc69qjlvfQ4gPEpqfNmX2HL5/HLykSjtXWVlw1xKYQAl
YLau35dWxLmAE5GPVtQRQoZek9lvMegV6tKi2tftnZ3533Jsl6SK1Rssy6j24yQI
BnNdJorC4leFqB+t4Yq7Z6thh0APz8knc4E9mVARoqFsZhanNvktA1aGLPlvo7cb
DX9LeDMtdQx2SSwAS2CP5vOMHJhQir/wdn8BgQJeslyw5iaVdJtAHruVq4L1gkmR
7XNt9nCMV8V8dpQz+OkXBQV8JAbAUfe77Xq0POHaMgbGmAfPRpnesR4s/7ky0TOn
G2cEqrMfNzLJVgZxdOCzMAhl4OOj2PIZ5F4Xf5MUUrPof/ErqlnYkh0MCkQBkjuV
SokUZ3tyZLFFTEntzogrk74rAU5AmnCJljKc0gK9NmGEchupn+4nLQ+5AwruAj8b
meo54uB0szxJdME1zBJmqMDjSDt3zNjw8FRJPT7c6YJPMjvMf+fOHGmGJXgTvVqv
slP7wze+pv7H9bgSZwhGiScW2G1/2l16MHZ3ItDhlub8nPffa3YmYrPmoGiVTCMB
cCw4JTyqXtuAA/S+FQQ22Uc8fU8m0P71Rb7cYbZ9gdF9sh7XOjxyuiQSB6cJgQtw
HJV51/oO7+OqFUS1Xa8X0HNtN2uNSYdI2A0vaDE8YARnRd6XWWC5e8qGogtAdVlw
i0roLxwP6TTeS95vRLD+ORKTW5zHR7ZO8RwpM9lOk2DeQmDQJrJU/qklCNBKUZks
OEz4YYJ+A5+bSR+jV3xKHvlKMULzpnnrn8/A1ipksNe/hZTmSCWFkaHn20/YU06E
rSyrxb9FSNnEoYj3g6inAyfM5AjTFGJfgQIUCUF3Jz7E/N9DX2FE9pCskYqyoSsT
5/q/XuSLZJbGRjr6WRzVZhN9QO0cLj/PDiQ9tuHyhGntWpasLVAcj8lB/4CGNaDj
4WpFNEyHO++UgrzyificTJpTN65qwMw5mPZf6u/bBhB0ndVSvgHRy3fpfX1+I+RP
3Z1totcE2CiZMlswmu8ucD5/a8Wt4qwN/X8Q2qsY8HNJUC5sK71H+6Onocbz1+JM
UB015JoDcinQbO2RXCgLtfi2d4WkQNTtPnCpPMz6an5n5epTwE4VBPQ7q8tn2X3K
Yfk0ycJ9dK1kF62BP9dkBb5S5DpGLweWi17UksMcYZIjMh+1rGrc8xPPmrH6qu47
pEor+92P9F7HySlG6YPi3LABt+GsYjOF2CzNQwsgdkHO8aoVEZepaCJfVRlgJshM
9d3HOeo3wfkrdFxiudTwVcQ/pZ6Eu9D59U43JDsYnnuISNj+726YnZd1UE0PDgZk
Fy6ln3005oKhf9dKv/8ckQrCGb0yiqFE1MDF9pX6mmEjBjmSNh6Q6rLYj8RvdDgM
vkCcyqEcdECXI/J7fCI5GaZwHlxlED+M2fqmVURWlJ6AXuWbgUnBgtDI0XhDYKev
CMu5nu12VoFvaSkDgo5VlhtIcZL3K0NX8XiN1IGldOHbCpeyOzFGBhbU46DxBr9M
JJyZyWnh2x+Yoc1l89y3PFTQhwHdligjzAGN1QIVEKO8vULDRUyDxHIWo8vAUQFX
fA3ZCMQ4NzXpEoTDsa7iYJuYTh75x6B599vVwvKkodN63QH0OugvZHHQarjoR/WQ
ATKe8VdOpNUTe5TZkegMLWlWe5zG6xxDcHVIbo16BPQF7TcOeOgKCiD48ZRm8LZy
GV4rP3GaAVjNXEdo5xuwn/zdA/wPuXzmHqfRJknDL8OXedy5Jf/+gjNx73F1f40V
xzmgj7luE3lE7HM8Ezn7gBHQg0Z0C35k45BPNlk9jhHTlPe7OsWvzmfy3nBBeTmR
LE+ZPBEo5Ovj1vxquBP1sAA8xRiEEsTknn/PS0JepjzUGbwftIM1tDggnJeq7ly4
LrxyCvJ3hiUFFjOshQTwjti7eVHKZPXam7lWBsC2rBx0erMmvdWXIGVbUhmk1JV5
tSyULccCQ8RaufWWYdL2FqTryny2QwVRefpgo9h91heaxxd/9YDOe322h7oAiHp2
QXUh6m5rcdE3HKSMAc8bsOK8XkFi3gdTzHBRlXvR7JS820QgCM2+uxe4qah+vXyG
Ut4dNRXPoChmIHH6weTtEHWQ44FqJWTCiuo+RuvkHNO1WPkSGQfIEmRmn1TmCGbq
Cu/JnN0BVv6IlTxHgh/0KRsxDc+wZf/qauMU7/vEhYmSQguHxLqeAR68ycxqrOuA
4L2Ujq5nDEgiRyJPIJsw2xsj3yJl60LB0EDcsS3CEtp18KMpIxVlvnNc/i5u7WE8
GmWnndZdWzjLjNkbvo6yGJwP1c7bZYHeFkIssgrw1BSl6pBQDPERYJkI5EgUdZMx
5mKRYHNMapS1acbsP14Y697go0gueQCWPE6x2JRF2Jef146NwWaaSsEsjxKm2Nll
RS6d3T6cGL3PVHxpjELdxex7dsD05w7/BNKUpK6KnLVDv2w9GcsICt48d0tzZRpx
dsGcRAw4+TQIY1XKpBXxT6hXPi8yN8dzF6NIpxU9cwIFLtl2Y7IsY4vUSgaUkZ5Z
z8JjkpvWSrgpDtuQoeGPII5dfRCk4rBrGcG5x76265hOmJJ5KySTJrsAsdwS8OAw
F2Jd3G1q8OptUaecOpw0IHLtv8XcZMKVYbttfq42eX2tLFnC7Hf6XhdDMnoFTzwL
EypBtCIm4ZuCg972hO52pl9t2UWUDeBJMuELJtO2cq77Mz12VYJK/6ZOdgkF74MM
NYsNRzMQiFTjzcW0LU+fW1cCihy8NMWmpxII2Km51KzZtyEx0xoKepEyIfJc3mFq
uyDN3XWpFRDlcoMiDwKwdd5YGIfothfeTOBITmveQ4NcEfvWHuXvBD7Z3h+I6D3X
D6q9DyqO7Qen04deJqByEjIoB7xTwgOF2dRnG7VODQQT0X0ytwNolzLDARiO094Z
QBNNPR5/lyPPU8KZOP/gafrKJeyd2Q7Z9Tn4pa/S8YYv5fCYJJmJKpwRzgUQVDqi
IF5Fln/4Q5x1evVE53s9v4w/8ymfbCEsu9+n0hbOjAQruLbfAsgrXSI6vcRv9oQt
D1aiZwwpWAMTkn04hg0eaFHPVX24SeaoScmzEIe6WjdhADf+IaUxGgE+p5q5SY45
WJH+/cN7blTNt/CrYdWoYIMlpwuA960/j4gXe5rrvCAO7l1nhNQoQqczxDo9trmf
4J/88VveemMRJEm/gPmfiPJaiHCeNfLLjFwnNyMwomkcnjdNWI402TmFHSSNZ63u
wFwe83Y26HEHS/f94hsQUa2UJu75Uc6hSF3FNMWf+9hkQAB4O1/Di0EX1+7J71au
/pP3DV14AEk6gLENhy6sdhiSVClbPsBcbEuIbGhG1VKzpyXeYxQpx2nqm2Lxikoe
Rk4GFhLXAo9x2pKYgYESDW9KCdwznADxIjsoMh20+3h2IUbECkn/GHvZ5s4RTmMM
3oPfJdsHsTlDSnOEWAfXFnNX6Rlp0VuNkmhgy5gTKFYB4gW4AnaOHaw/2o6I4Jym
W717J//iXazNUbDIYS14umWIzEGXPb4/8erxvQUaLIS64xrj0lSG8Y+HoYysdHX4
vmTJ+jIKUAGmkVXsPQEO6upS1DnKiWXZsqN9JHeQQYmXPMIBOT7tbPTvgg8lnyLv
1Ynv4ZZexNkoz5Wafqoxw8qGMsalV1v/S/Il5S3gBYgGI4pUVI6oW7+b/6HfKr0F
oN5TWbyvGQ7UvcPoMf5AQG2rB7g8nS1atCdsf1oJco4k6LiHdiZZr9v+xbah0PYo
nM9AwiguxHQS4+3wrpvcNZyCKaAbauyVHjEwgbPjX6yzMazCISIFif2pmJ7nNnE+
u5Aowdwa4TjKuBRhUX9ghSEXrbcMG8RAPaxMlI9qyysOmgabyiSIRoIe6b9nzUfT
K4OyUYeUaMsu52LjcCU+bJYnfjhL68jQWUj3O/fwX4PF4ClH5NlRcHW2S/ZHmWEB
RJ9NZXCLNbR5jeyRgn0Sxzyo40aU7Z8uZRmR3A9u5/4l1JJ+pfd/YwpZeC1QfEzF
91hMb1gYOC4oz1C4+tQqwSo+WXbDdT5HRCtfQCbsHup1DeiT+bxuZVXEc86d8eTX
oPwvDnXxWYeC5g4lUPcOsoTxy2p2XatBnnSraLnn0blgQM48rOD0JSLuhpvtoatC
/1SvT2L89dVnNKdTk+Kj0Zx804ANGNH/w8mflaPKAFDRTzR8tbEkBkX+hNqBoHuP
+KDrRsIKcik/BjGFpP2kN/jmmR6Zod6zwa8TcFY4AmFkqKJcb4+bQGCjNe0Wv/Yp
eI6w2W1FsozvlzppKFtTRiRI3/IQ3kMjSlQ9405zXbobqHoCYdu/i2toC1lRwiTY
JbaajE+tbVJudC0mGRtJL9GItzJ2p9V+SUme3B+JLgCApL5z6sRGH4R/n3a++wfj
KqxbuEbaYIMlLnVQI/itSjoKF/RmWq0yCZ6qf1diUcZ4MbPxoaqnntXHL3+iYNh3
jgMjwSGQJpY6GXez48SH9O1/TkopXfEeA14BO6J2xDC+rTnoNwaxuQd2ITwYSAlv
gK61VKia0E4b9GPRf6cn+L+fXa4aVmDW33ryLWUUBG2yOJVc03C6+lqqvaFyy/k0
4ZiwnmIHniC6geZ1JGpTOUK659Wxa7pziEAEt1nERA62PFYGziUOYaCH8wkGy2eR
c54u/MRNi9L3s9HNR8agc0oKnHYbfQsS7AiVJgaYl3k8WOVeRwZERpTeALtiQ5ge
PNwmV1AE74vWdyYDQW9EhswaYZGpkDyoA2FDQKzxSb8A6nJRES8nBIWynN0/VE7T
rrtZk823tvWNhYsdVp2X+RTAPmZVbdWjxwvIPhXWnPhZxtdS2wvzup7zZqNXB2ek
/fZiQE2nxdhxxXcl80A2PWxI4xEN5tOpgMANMXGelqUDpZSoUoWu8Ip3KKySjVGu
YpGCp8lf6nO45ydcq0djcAW2IxsQZoaRudvLXqZfqky/S+5OFVkHjdWo8p85SJd1
ZsIAn2fbG04w0/Ba5yY6q9H3Szcv44LQ0LC9annGuU2BJfMQLrbwjyh2t4/+ynQ2
+okJh9aSH0Vw3+g5lgft/l9GFpo0gzPfKtZCIzlm68rjvVy4XUQMPdl0sSqtOdo1
essjfp0sxSlPtyKvtYktpYENJorvGwVp1XQHxl4ZkkJ2gN84hFxND9qAg1bsrhCH
ZSXtdrOaGBui47Z5d2ywl4EkJznR1yLhlcaukPYFewMsCnXnl9WF6LzXGc8RjLen
4naaUo+J79vD/GPhf6cl1e4ah6Le1aLf/TPZSwvyEpEyp0O5BfuZ34kxzOGEmuwt
TyZklDVFSC3mSII7LqwMlqkxugHJsS7ZoFQWvQWZblssTBV5IAPoMtjdbJ1Fut9L
lkQp4q22BXikwm5j10679CAAL9rQqhH9Ov/ZWeOPbfJiGLKFGcch+EamxN7WNJvi
IbwB6SyZGzN0XsO5YLH01yQGT+mNKJQph2sjfWipcO6fYo3uqYKM/F4GDL63FMMl
MmQ0pWmGs/p4nriIr9f9mhdGclK7cw3dACuY0/RMybcTPFn0EcG/mP85A+UnJLft
jHalN1oo9H+Zff1gJQAyaBwA6hKUT+fI4Pp95Ud6ac320jhFHJKbUc8SbpW83xfb
e97PJmPhSoK46LhPP1H8KdAGWjoB7LZdGZKRSkDkhgAZk0bcF+h/jTKlEEGrZR7g
obdjj902jKvrnEuZBVho12RmgkEovr/krsk2fJMm3TXH1fIdEzvGTeyP+SCxQVZ2
gmBGGOqA6zLeSt6ZmXIntMulu6rYdmvcVWEqMk48lepP2EjM+u6V2OIkjJ/a9nV3
Qp2ao0LWRRB/9lK2aIEaUsMsT4Uibwyh0z5hh2x0tptMxSwY/zzCVTUj9MRK1Dod
oeTcUUiSpU+gBObgm+2rSPT2k+xe5iQZVdIfzPtW6i1cfsidYDsdJZcf7BqYM/fB
SVxGk6dRks6km6oAxiyEPszPIhwRt3oZnlAJVtAXrwc7mDqBsEqN2MqbmlGsL1Qt
p6SYRdNjc+32XgEl35MWTWoNxw+0zOEeRw7T2+8JkXm9v3rlKgTqpbPpNzIDt+BR
dGgTASwsyxv4kazzmcXW5mnzBGqRh5BQwNwpGXuRKMC1e5dttkBBcumC1bXeYo6g
CXIdOBuD0NzwVFxn1JNMiQejX6l2lucB139vwIUDatlMP43OzCAwoy0SjfkpLnSJ
2i8t/Z/Og/jmdwUTW+GCvClAuh8dzld8le4UzAcu4EPhP+8e6B4/vPodtLfkwuqm
l1mA8Hwujr8pbhjtL3NnibrW2RTp78CL+KTmwH57iDWK4/e2vIQtBxU8B1LqlKzP
TKdXfz2nXPUoyyx4HpKv7ROBt6SCgun1W4zh4halADUTwpVjTpqg2A17s0lA2dJ8
XogEaNmGrYOVE7nzkhPIWt9GAn1MD91gYqAfbrObApmFTHjXtFY4pPs+/0zcHoPt
PeGunddDitHidZxIwszZdCXECPbpftX4sBwv86hcBsVxBG/WivoBlixrbVpg/xud
y3WDd5zftQ9ijrmwRs96tLqQHvrmgAfXrjHWNyXcFX3vTkpciJAMUgc1F7ZCOpqn
YV/vnOcKsuInWpKF6xWxr9fjYduLKHxHcP2vEOMGhHiUPfk2I+mXCTrBEJA/r7Vy
K7p+qRLn1eU1UXZns5Y4iILOTHzmtXEY3HdouowDD95JgCEr1iV/SRQmlZYREftq
RM2uJH43JsT+rwCrhoLxS2mI96BubJoT3fU3SgTb9usIvlMRBFybpWkPu3Zuosyv
VmGLEu7zTfwkfUysGzbhIGglW7KDsB+uXzqgwB9pWe6zSmjXmANOVFefrAJZi2Ca
Z8bOAC90rw1gD937VeUtrO1fOzTgRn4NkPItwXJ4AgTCmmTuZ8NPJ+eRZMV9nwhE
DId/+HosUOdGlt0yeeuSpP+9Y76udPlgKJQ/nx1NMEMOdVNdxYzaAiR13vUylVTv
JhWEWQWQkEA6NR7/PfmMhPJu7ybvZd4ErRSVf3hZY8VCnh3mu0MZfPsUTinK2qNn
YCLjsMGkJzK7LgI6mxtipxyiMx9Txw8kDAviXNalgoqFCxTLN579PiHnc8H1fe0a
/D9EI51F/HKsQRud75vGypUBnDYug44Ilu3bqLJoMyCX/EOwdz36FL/j6NPBgdKS
nbQhSdJH/4MgxZuj7mXZc0e5zzlXTqMnaKllB29GDu/tTxKkTnYdYd8xo/z4sbAd
9kb7iCXCamuzZdlipP+n1V8SLhpkbBDT8EwtqG4eqRzPSqJzIHxw3z3YbIeDNrhj
5At9ppv4M5Nvdk8GTGxYK/6eSvt3HvRFR+FT/sz/xgZma3vaxJg4hOtiaR47zujd
bHcn8VlZgGpV9lVlKm31ckA6gzQTvw7bwUq+rlccg77CHvNZZoVbmHimCk+bFxRa
1Q8/E5j/53k09A78M+WD5hZKEyEpudNJPv+R72DIbj5rRAMKzcpNw3DVvQvvZfWH
hEY6CuZ9Jw8QFdUinPlo4NRxMG63jiIY+y+4uvZBA6fRnuNzrQRYg4bSe8IJifQB
D/qSd2rEm2XG5/JLeckKuauZEabOKzyHJdJVlDMmwuMQgdyexVvf0PmPKx6nIrNn
ECI7CXysqwuyocj8nEYeLF0aD4q2ox6zth09u8ik6HQZCivEKIoYgPpDljtNSm9a
VbSVs5hz5qGt0vTGEpdkW5NBtUyNOvrN8QmHHSegEdZyCNIN9TdF+GdOi1TVCf/I
EBndzgQw5UMTtkA6r3v3szoTQG6mSJpDnjYOo6q66IvhcSp4QAXfNJyVT8hHqbc0
qQKuoYiT7FT15/cFgNetNUxMkrKR+PVjp5r1CdBb3+y8hDvqqLbpLw/CMuXGWAZU
A0HOcdhaAoYCaXiIMdAZB9AHIrnWKOLDfqAO6gGW7YbDkywGfm4WOaHXXpmBnlzg
yBVvYhb4heZF9ZnP65MK68DqjK34HErMzfVYoLoshnNIlQjbtmn5/KyLUPUwVsPc
d2HOgatI9eZ3UKy88kLv5u1ZRmbhcFF+YuDi11GHunbN7M8dCKH4QtOyHC8rJEiK
WXEBG+5j91Sne84d6osjbMQMg0CzcVfzYT0ienLKVNeShUusdTua8UYlHQwf238f
6OkaOsXQYfqhwe7u1Aj+4h9q4Z+aod7z1f9N01r5pdEjTJF/ogwI3oh5qRMQ2F/U
7n/PO3yBveNAXIX5nYt3BPTUtY8jIPT72ryynbDgHY4Ngww5VekJX/o3xqM147As
K72oJWJhjxn+8EtgMuYj3aJIZrTqEIKJJlhqVi/EtPnEp5kMR/IHXL15/fP9WPWV
bWwZCviFXMdmAxvSncNPQpKILY7CKJprPAjz83Cuayrh+YaOUs3QZmM9hrINH9iG
x7imeeeDezMpQAqGDT8F8air4ua730JP/f0Lo3CpNDZ/X4sfsRym+6DjVPoG4eo/
kkRjiA+a13jLrrxEFWl1Z6860zbig+Tez+tk9jSpQuzCn6QEmZlLrrVD7QWvmqU1
w5jLSD270mWzoD+b+6mOA06wjVKmmdo07+GrKtRfOL8KOUij4DU4JsmR+6e6prhi
BbMtVxwf0zVYXZIQVVKfkumfdPK/yk/5dhNq6zBDpBfTs0PO5SZbi2UCEbFEVusS
BKbm/H0h4XWZ5U82aYqcsFAS8F4GFRGg7FKw1xkyPviT6F7gSWUtIPZRmh/Z+KSh
5+u5t6MUQtuwFStiUT8nbJNzsbU9vAB4CSk6rbjVIaxJH2zOaHgAHuI5FH1VuD0L
EDLsWwMgyDOxb3o1gbhxfZlDexi83u1YhWLqf7sMSNr7u7cCVkSHMbXSLZOzPbfE
YOeOyTKixZUvXxiisJO5JBPhWVdQ5Z0fVBaM8cBhWaP8fk/iW/6ctBUDG98t/XaT
SxYHw9wzo15KoyWYY4cBB/eABAEyXZNaTJLCbav+XuBy3VtO0ApXJSwltxb5CVet
btoaK5FIjErN8Eg6C2K5BwOpoFRtOZYK005jIdUOauAM5yTx8LUWDx6g6GuHTgQo
0gD+LPLrRny1oWuDLkrxx2f0odE6mmI95PfdfXfWS/6eAT6zNYiykQ2kh5qPkmhs
33QEBrptt+PJ2SWxU5O4CBd+GnNXxTDP8RUfULnvkiWJbfMflI/7Ahv+KvKC7adO
2XjAi9OvPizrd2p5Sz500J3lQPaypWpeUZ2jUzKuODdFoaqtwfw+Qhs63s332b1Q
IBrVeZPH0UUcQVRvLefVg3PQGdqGsG6Lk4kFozHNxiUZU4VfX85y8WiWD42fyerf
riu48ac7xi5AEVrO7BGqKs1GE9rqRX/oiIae+b+SHtLQ30H2brI7VcMBA56Dor3o
rjmTyUASVAa9Acf7lnsHzsktyd99cJDV1E8BJ/w2Bl1pxMP3QHIMYL4ed+yDADZi
cuoOFUsO4LhA4jF4qcwH5ig9N/gUw/HQQr63z7XUlS5Y7wdJUfo3D6nge8Ox4Lmj
mev5w2IMZ8CK3zx9R7UKJ2jtImk11srstpzR/3JJSm+7acWrSWqTZ7QZeZqV8V7C
2IndBJLnZpuqXzUApL90XYrdBYKAAAKIQVg7HcS3gSfIOvvrxOy9JZYOQneHzZOJ
0/cE2GaXhEHneIJp2nnduExuK6//17uulS+tiughGD1kVz4JvTFwOqqPrKzjf7DZ
f//3o0xLw/odQmoDVV5eibjIvVyztBydDLq9jWqkxljemv849AJ52nEGHJ4Ok1bR
Nj8yGfdoywj7MRGp4XHAQMZu9Ag6LxHzBR0PLA5o+exRtf9Qq0m6kWxeltTpOsEM
AXlhcL78kcZRsjDF/SmwflPs3caTd5DMBIYMuUsWVgm8no+2FH2jTEWXdr9kxDgB
JgHwpZjodY4mnPFWm6D845dtXgI+/Df4TELGOtil/pTICwIedWw/zWeE+pgrk9sA
dh0+hgcMDsbJZwA40E7t53CyAibbX1wrJR+MngXP5aD9HLYOvTc8izh4jp7PCSJg
lpEpmfPwdavq0wkpuVYhBqVirpJWBnYrZFdslYnrJAeOjwHT5nXu8HhTPcbx4tWA
FQosSuPH3zeQAZOmapKziYhhEJyoWDStuJZS+JRJDvQpXqmgdaJb62Cv4NxiCo4h
Z2c0e5XfoGOCJtzSVzZQSCOcGbC+cY2PXsB/qIZ8C7/NQcz3hZHv69BpdZoHLbmj
dbAk3vr7QQZ7ehrAPZN049LReO3t4sI5mYRvMQFMjTN29abCXMln9YBPqKqzbmum
62ksq83TcjfHyYHN6LzHO+WuHTpvywKoRQnwJf65H26K/wyJlg47PTHuvFSPhEcO
gcYdj35aZhA37iurZ4gH92FqeVB8DIBbI0vzRaoH+TRPxQeiN4VrjedQpCVaPFT9
O2OF5E8H+FkJl/6zEumoKNaWqJf1egLXtDbG6VBGHUKmm9jFYcE+QZsORJdauOqG
+79G4U4ZF0dIc70g2IbymmxcsPrJax/WZVtlTxjb2nOKVEw3SNfmIsSRlb6Q8ggO
pNiPiU5UZ2+h0gGncfwiy972+DEM35Ig6U5VdwM2llDqc6VZsAEfbttukkc97HZE
RxRLTjH+zdtCnecFDYh/w2kED8e+7NOWtxzekA6yU3yiOcEjfq6RkyMD8Q34QSmn
A+ePLqrIE3qk5zxQfsOkXXNqzW/R4NB/NiS0J3FaAzzteadyjD9J+hOxr4M5LAr0
cBS2zojCo12QbNM9p7iSzEksqhp2+NuguYW13IZ28/NY2ig0j+wuzGEykFXFBrhO
1Yc+0qYC7x1LLHjpzMZxoRyn0UqQcTY6OJBvYLwYQXVUBFv6ltdgGECV+23LxoWK
NkS2XE5V6RlHPzo4ke0bSHTR79JqBfnFpRyXARo1SoYocmeQvWzC5JodtAeYAi12
7MtwbvshJEybneE+/fowTrBrXmVGTAeW8Y/MGNcQ6Zzg/Ollvjd2rxp+X68efvng
HS6GSo2wpe7/EVm0bCiqj3pXARVe5XhMVE/X1r8Dw5gE8nwbM5JRB1CG5b0Cebkg
qds15qZlOPVXcp47myw0wd4Pap35M7s9gFIh97sDikooQH0z/zNu2DnB7FXHrZzc
UnJz3YR1sZVdsKHWX3KBqw0xPNp8uBYV9DSBimn1UIxuEv0IMWlJmIPIth29r3fQ
0rlbuUiqeNNg0Ld1L1S0hZmuFgzFIwHz/4gud8rrQ8tDflS7QNDpiFBPHVvReGMi
UMaw+Hu3mTsaJ2vNQvKOmJH57ZKkQ5dcwMPcfIeAZ2ElIbMCqRgVROdStlclEr/C
IM9RmiUmS2SXIlzvaLMDgyyZQ5W4tTuqRwASlDjCcCSCNp9gh8ZMHIOL+CPj9xlC
7e8OV1GvL7pRi3tqVj26FIAuTIXqLnUJbJ/VPz+0ouh0PhU/Q5NBfSq44m39TlC7
xwk2Lw7SCaNU1VD/4KI4iBqNHkVkGMxmtwrmDgn2mN/gsGfOV8CFQDGK/8B63gPd
iK3BHPYHlSkkvum01MdL4e+vOCdedre3Q8Kcx9lCTzznflCs9AtL+VKaFZ/YpqfD
W94HLWLS2JJ/5zKM2vqwig5M88CnfG2j/4bUi1dvLO4VXWSHTQvRJx9U7wjcgBfO
zBXQcmqvK00VxOCmIPEj5zO1noJZgIZfFT2K8QJK1Zo7rFTQMcjNP6cieGQOX8yt
WOLL0hda0Lnbpr2YhQ0+M2Obi6Ptkb8swY/OTQDPuts8fNfEdKiNDL8kIPPESYBd
QadzZoWh2HoqZDtOrpE1Z/B3TYCbV6v+20XXWwOJnZNNrQBN82fTX1kiSR6exR4k
r1LCu2F3IXxAQSi45BKgv5hcFMoFqsQwKp2+t6R1YtSOqSy98aSSL3nZ1FHPzymr
Gi9zV2sn6kPRIkjL5D9jN4HWWROWTTJ8C9LGNac66xDwnyleyesJEWWPQPK7jCrW
4fV5kl/Xm+tXVf3n8kZP2/egRHF4v9x7KV94yyV89kZg9Bl6efvH8YLuRVyyegdC
VWwIr0IcJAOJkLNgI7KmNQCUcF6zlszlQWmiE128vFPEADIbiHKlmOMtRo5IGQeJ
ADIH7sI2qPVh5sXHtXa2VGW+CesL9apF+ZPmOu9yTJ3cdvnTYAZi20RnLcxe7as7
kRS0kDHwj7jcxTTiNklLqsY6R4Ca9E8b0avprqchiPWK2xKYeJRVl4YV5/U4Sh60
xixijbcGgY5FoOvaulCQQ9vwc/xCm8W5bvs8F+1ub19xET+DapOXu1cCJTzRn4a7
6W3Xq9oZlqcTizRfEq07Mkz0Kb0V4N3ByWfmdlbWkBuIhyVWxploEYWRf7ZnuNfs
3HoIxt8HRuRhh57yaNJGVNXrqGUXOvjmyIglUx0+dUflB8wdn+ne55d/BgngZh80
lvZbrwM6e13nv1iENbwQQMxIs5Q5D3NAKCeP3CiLpL/9uuEgh8XeXvNFPixchPPU
SXvL4RjBLFXuKL2cRew52rmG/16JtZq6ry+l4LF6IuJnU38nYr/PUxk5EtEaS8oJ
/6vpmiXj51hn/0UZAsO5rnxvsuyIu7U6knIGxt5XWL3Q3iTo6OQKGyUqwSWaJVaj
DWRIASfDPi5mC0R0sTuPHPIfjFB4bL1ZHefrT/QJjiklOshchNGSY6YpGhmGvBxE
QJar4b944yphXeqk12KAyIeQcYrsR1GS/ByPi3f+st3ScizxkcA6hiKGthv85B3k
VnT7V1U/mATQflmWd6FTQe6Jj6bEbVvuibFztS2BSD64Dma6csyRuIVSLsTNtcbL
nen61E9CTnY8i0rrkJcrxWvgE0FMDBFNpitmiWNK/MYAkX79XaJhcZJyTuTkB50T
+dPekTfWrA+4TOvZDhLnMubO0QbfeEscpbqhy71gQfzRd/C0wU0Daw9lb+0fUf7v
LOr3wNS6O/6PPjA+KTRreGXMMIAMWGshs6t90s2c6lO7/V7/zzrhzpXFMddcs3Qt
zO09jQIzRwjw52EWG4LrTE6dPNU5wgDUm3nTO8Zk8kUxc3jI+0nGoSwQUPaMt0Qm
BFAAuH0s9VqQPVguHPYeUMxvh01uVdZiboUxrcfElIbLy+KsC91/TEtfoobvD2Ko
Gv0TOJFccFT3efrAlSm993yKDAgD8e1GCrhofKrFKHwj7KC4DzEk73JBCaCMynsF
sB+0Y9ABgOAsqVgu/mzbXrCG6hFJ22dP0EkmoMKWR8Ux75xcj5f9VL2xqGcF4tHh
igfYGoEHQR434c82ObNzFqfIDxmNsjCOUdPqktvMsWDO8Keg2tL0cqKuyUxyCoG6
GizABmHjKlwiLo5NK0QS0239gr8mGnoMCrx6EYTwThkcvX0ij2ohtyC5PLp5PW3F
Bsu+mt7iW1i+FuWCK7SFmetE0qj0If+D/wOCK9KsdCVmMjsyOYwfA2rfKZzvQcZ3
w2C1ciuKM7RmdJExWuANoES2TzLSSgIooA5jYZBEEc6vVM/1KzIh1ZgpWCInYIse
vkdXQpK8x2HY6ILGDBzBwKQqtS/pX3YXGMM/daGOZM3G4OqoKleKhNemCoDCkKVw
M/J9WGJpVWAtxDSQjvTCjZlYCMMoDlsF2FUOCGLvgJEXNygVPjClnYUnS8n7SPT9
ace8IwBGfhYTkgE4oiW3YbvkzaBcQ6DPNUZBeogaE7IqlhK51d770gL+nD9DWMpY
mKt5AnXZnVs856KkikBvXFg55HWPy4RldD2Q+5s3bnAvClo5+nrJii7+RQTUKPWs
9I9IeI1mFEBy+MKgj5HNxZBglV1LSakwuQGGmnB0pgyQ+5B5mxlqv02gQg81S48j
gBu26j/Oro2aWKPQ3fpx1Kzi0uMpE1cjqCimlwdOYc39l/4clAwErdrUumJckr+g
tL1lkza3Vyfp8LSxYoS/6ecECRBzVZ7VAZRcqBTAUnUYQnpgEbdzooprd62ABG1R
BCIflUwm+goyD8KDogzFSpEFk6p1MGwPZ4tW3y65W+9IUMenlC/acSfdR9zjmhAi
R8imc+JCi7+tdpFrHqXinCH55lp0kMi/KxD2OM2AsOjy+1gxFm6SBNpPvRceWZg0
l1E44JOJBNSQPO2XcdjUFBlV6BnZT8PVevyXJYCJz8gSL++Sd/KIFfA/XcX3PLZ5
5th8ooPMCPYzvnQcitan5+9KmAZrwEbAxuI8kDsAZR2XaqfvtaK3ihXNe/dxT5D/
VwjKu2pHUjyGYe2CMOfvE+UwOc4rixJygkzF9djspW4vgvRWfA/WV017VsksYGZZ
/qr8r/lm9/AG5vd0Mwk2wzibeNzRgGa3Uqc2LLumtVvDt9PLMtVYKYHXvZHH0tOD
FFSEAwYUPBXOwp9IHrZfpo7iRmlk/t52nzgIyAmTToZRDLKL7ZJKr1EZa+IsswgW
ILoqB2O+RgJOdhW3luMTUs/SrBHsw4uBv5sL7zZGyNt7XcMXo4bNOjr/2Z/CHL5A
EkGC8oIbxI9RfWU5GT5TUpdPznCU08zdnCL6BqYAWkjP4kxLTgdbIDZzZ2QVS9zf
mPVFM5Gv8I/rQZX+tPYAH8nmCzgeLJWsDA8FNLFh3sGBdUtwuTEiwwr9wbTCVf4Y
OOePX78+a+emiZneipZhCVEj27vy5xlJAO86JEh/1bT99iiFZp0WiQOcDPjYto9H
nhaqpnvo8GEHw4HW0jKbBLPzdrAoUsCf33E4yho1SClmsp4Ii/SHoV7MQXAWOybg
6ZIBdIfcuUt1VvtSavOH16q21dIdwZyhVJGT5plFctX+kuJTtba6Vg7HQD0l+9aP
HdH7ubioBfQm0z8kRVPyri+LUmSNBPV5RAuEvA2bsOYimvZViplV1ShiK7AqtpIe
GWrMGJZ8Ez06F+E3W2SudQ/MQLdPXYG/goBsj3JasKFou1NHwSY6Dp4g3f6/LKUQ
IJOf5ixccrxuMmKSnp3LPRdvbOYRfe0BlsNseeceA18+lwMwjF8tU/mutyIU4f34
aPWWS2TV8UwuXRDUThSH/ERbvin+biwTeZ8pE+MECv84yuj8fwQszNJEor4vNEvM
KpOtJJhs5b+PNahm0R6FSKFKpxp30P0689xbbD3PyQsdkvOBAc2XW4DBxs1gvHXe
HAmXOVElrHgO7b0ppkHzRRxSm4pVt5wj2nLDaZZIMn7DPK+hCLQwSbAJ75/0kI6o
Kz7yHEaI0tCbpdvSCIbpek9uNOvVDQl/Vi5+ptG4gzDvyAxGinbNRUCRinZcygsK
9EtfzbauoMVXMORSVVyW753wzxe0cAcEFKVAnqnbxZceIs2302T4axRLEScMSS3t
bpy/rpZwH3nx581KxCLhAx1aaCEzfofOAQZaiBGnaUPsThFFvtmfG03dxow8M0+n
3UJlQpY+Tj1gTziM5SgiSCTD6b1s3gwG+XBAwI/9HiMQfX7vPLkWQ7ljl+89qwx6
O+FH4OomZWd+d9rZdEALUpThXBSHmNjnk+hmdruR76fPmgg7Z8FQS2BLz65zJwce
+cutEsP6Dw2dI1UcSDzh6uu2dqmY4Gd3NZOCp3WuM5gaFCXuSZH+/qVv2xG5uyyo
dO8s1CEtuyZVm0duoRErBBIIYwwZraJelnt1PKOz7khIh+ElZ1i+TPsNgIgCp3KC
AkysIgaDZea8EXIVr1rBwVJKfIzHFeZ04UxNlO9KNe/AaafmdUltfo9BkVkyYhuZ
0CjB57T49OJQWWvQ+CM7Z9CW7palmUNSXPx0EekeY8EoHWaUvoUd9DWIWGkZQuBe
S279b0uHEabFOV5E8YwKPWImLog0bRjmmXr5sTAugCjm93LbS1X8ew1kcj0g0+hl
0u3VSrY/jZM/dUt3ksJGMRle4wJngQseNZQ+N6Z8n2AJrDB1ZmE5a0R0a7HbH8NN
M4c9rAnESP/DzNhNbBFPTSya4XBSqif49MTIRf53pfOytN1NGTOZA6863KfG4FHN
xAgEoVlD4TsPD+J4FvFYnqPzQCqE2RjjQOxzMOR0kdN8XMf3wdPPuV5k4b8MUxz7
ZlQTn3SdM38KLOv7E2fYx8LHL4B1y2wPovfqwPCA9OMx368OAAfdSNhMJLykG9jb
meRXXmivNA0Uf9tNWe/b3rNg7kj/6zSS/iDx+uBhWAQ0IMMGMkR6UvaVUzBbe2e1
dfA3/IxFLcpuH5hj9S9cvf7yA/XjtM3PdXyQbyyKETT3IDBIxUC5ULbmMDf37Cj2
MJtgXq7bmRREFR3eDbygM8102KbwW4wGkx9wn1GYk8mEka6lBay7HKQkZrWwSHL2
hZAyJKpN4DgEOI8nn5eSGItpR8QKibyqr1HEycBnYVqZ3uvra2i8sy4ArUvLb/Fq
AGpymU67rBj9ixE43d4xKKjqNISx11D3iIhmDSITCZh2PBBEiP4QNsOz10Z/e49v
8L1hhci9NrYVjdT0FvqBwWXBBpPn7fePtJXameYWNSZ4QUrXfE6z2ACVRLfLeklp
EP/rn8CbZr+000qrpr/m+cIvvwXaWNjU9gIYWrAWdkq4AdZvjB6tb1Lo68kw+S2l
ciNsjBeQlAXthHH+Y+eUof+X+UWgl3812RKJuiF6k7I1J81yvWPoM+JIQUVL9rkL
cJzLpcui9Xhp0mL5uJqk0vB2D5chDFtuM/Mqm7V6rb8p8IKrS+t0luGeRYkJvo8f
qxp7y0svDIivAGafbjaO5r2NUoVNb9mj5KsVnLneJ6+uimay7BlpyvXeohd/lHQF
8PVDqL4mt+HCdVXws5oAtg29x1kVqiZOlidPsfVlcfcUhqmcWOS6ke8S1j8yeuwr
bLTXyXkHVJrmNMz9WiKhHEYm+EIy6zb+RoRjedAlZnYJgryPzM6yCBwV/ShHh+uX
mNLTy/9pa3o5wlbG093qiIr8cWWcHUPtB/jLtXJbpdO+w/yoNRKZwynX+FJTwqcl
JcDLSZ80xJ6UpFG15T+40gmvZmhoeV2QsaSnD2kx4EKMeS2SoWzZD0RgosFb6ffE
mFiicMGHVKQWFozKwloIfWkXpKxVFz+HjccrMqZewtx5pKwfqxhkup5v2V9dQgNi
RJ40Z6LRLJpoyVMVeX4k5R8EpJ9JViB9hoUB1RYmIIPbNMw5mGtB8UocPA7fa5zY
HQrpve5vnnoIE0QNglHKQZzQ1D1XOg8N6uPpI3YD3KIgCB22qB5EE4ULpgcg++dZ
vrmivUwxoQGgQyHgItEBDdL9utScI8NpcFaeJoZ5oDI0IJAfsN1auq+nmwga6TH2
GBnFAn5VOAy0gJkUlaDmSdaSllPYSJi0WBrXwUlL8qZBmXQd4uw1PqxY6Q9NIiz1
lV0N7/1zhb6U0dsVuxMyNwNNaRd34jZsTA3xnYv5i3e199ckVAXVFFxEiDYs8Hig
+4GRMT3lj7M5CluNWIZ3U6IrLLQct++miHRo/IKPOYBD1JdLbAa3NE0tDAln0iqJ
NpYXhzKcpAzfKhNtn17YIoSmyXj1KSwCyHDwA5YcIOCpOnHPL/m9+rQXOQ8pOd0e
u7CW9FjoJDOQhqokV6DsDtpD6BSNPLuBHtlNi8aIVzgUWJK+MC5ym+LBrJRFHfww
v72bQ7v0wdSVL8XGWSvvpJnP0kOthZl6FA9B5fUMak2LacxZGjYdmDARB7SIldv7
dAKYuBGpq/L1QY5UW5X59ZdF1JUJPiB8rDAqGKD17Kbf8BVkdqXoVAmBjIdC76c7
YuR/D7EKNo3ZT8hoGvISgwMJjdXGpprEhnTUeI3XOquYbgUg32AHLXvFkSCovtKZ
TYW+bwwpk8roow/fqfeX0xxRHVzKdS66dsz1sst6EHgC795qWfMTJEMJ8I4fmmAu
51EULPESmXQXlTSGIn5G/9ch487NM1V231GiV/ky/ixNS7gm3GwSBF/BNepjs+qA
pAaIy7m1H3RZvs3qsA9zhMB0Vs/qF22uZ6l2kiS9bvk0s8VpEN6Rtyuheg0MVyx2
4hxCB7Dn3d9ggqqZC5jPUC9Hljj064/xF4MrZmSlCDKvU08K6/bcQJkBrP1kjNp/
pSr3lKRs5sWVo6zo3nds72mTQe+Cd2qbeln4mXOTsa3hIEe81EKY0+JH/HY1c6C+
BTyt67eHCho44GdbH7sbBGZJwRhKrPE5SGm2WaMmqelp1y4sxtf3YbcJtZsG88ns
HahmM8Oyid/xIVYYSwylgaFHAU/wCWDAv5ttTYHDom4Li8s/i2JOU2QfwdUWtY0A
lwyXa+YoLymOitFqbQ71G20MU+bLZpmoz/eBTZIUuZ/ZSnXogAjESharM2OTMT2k
sU7ELNwrKsltZdBWLcRpxS6hVDOkK3/yMokNoX/EApIKAFUd2L/XixgHSqaXESZ5
VvQPqlNJwNmSuXrxxEbYTwNvFpk+FTOfvSTGSnH3PqdARW4wUT8likuye6A6oL8V
vcScF7fhAxne+E0+2KRxaFL3QaX1QjgyVxDQIh7oy9K8wNTaMs1qKSgEiFd6KzjM
qCqfqbQG4W3lSgfvNH3IcDOOn3O/JHjRA6XyfL/PqBiCLuZhFIgKIJLxXIuF12iJ
6AV8dIJMVU1mhxexWzlubg9Km3bq7gI3e65TR9RP2DzUS+nRDP7TvDtj4rJpUYFU
VCa4JMX86fYevS6rw2Z3fOT7nSa5fXNXB1dhdtlTqcfQC29ixgIsv8P0wD0H5vdr
WyU7oQSVIxxwvQDDrWDkWz+OgdljTFiMXT9TDkqgqZy45PylX6IbZkvcZIT300gq
EyBFC0QldilpRvLMGXrMX5rRGLM3yx6KF3DwH+VtIWVjttu9egJBQHOACnf0r0eC
EzlRggJVqIG7Lgky/cSha8we1BMKpUW45h6NHbcAG4bMOzXpdceom7pf+XOc78+6
5N22F9baYnz9Nq23WL58AuzAp35CU0z4nZMxaWJALPvBtb19V3ASkDn/fyecuHpt
BlalHGBoW+L0m1eoacccBr1gZeRl1erBvZBPDSTBUpEDbAWMrNs/Hw9l/hjiDEAY
Vu+1pQ+bYpY81uQn6szLg2ZLQ2Q8/pGT+OPW0uSchb5/ucKQNFBTwBLDhSYDV6lK
GN5sfTA/DhMVUN0x3cgbvb3LGQXj6+TFElw4z1zrFdSToKlw0dmOo37w4px9mhD5
QS63LaTY01MyRLSCygM8xfWbfN37DdjVqco1pLtnPZ+hIMEAf7/0/0TkNd/fm/I9
nNOU7d3h6iiVQuWS0vYf1Wy8G9+PpGMMs6+bDAVpG8oUbCyFN4RYl1u00mI59uQh
hs74AnuYEkdelSKznhzynQg1hODXnVpInuOF/155S8NFLiq7nEc5al200UNDcttQ
IuEawZQHvognNctXcRhXYmtg3aVK6EBeBd/QZn8pP04EJUgSMhmQZvBxh8fyY2Un
OhGabwIIraGHI4+Y/XoNNZ03fSvKNf8JAllfAckO4tspCWimMrG6a9Rx4tL/Opo8
QMvplmA0i/c6rDaue3TwMUvi4kuKUnzgCzZnllahP9QSH8p892WszYXUeru0qSyb
1SvAl/djcjqAPwdKNSqLed8Q8X/RmvfthzSWoZ/Uunq66HU4c6LxnF9U76Mhze08
L1OkJoQVEHZfp8/Kdwg5gdBR8ZWQDUdyID3orNs+z6yo7V6wVJVJXjvc0utZhNbK
2V+G5nZNAiIVJDQ3RL8r+to99tbuEO/RFPFotJK8cikfgv32eQ72fL2TUm1PNqPG
dJ0xR9zAw5atZiG5sAGBHDCYRkY5LUGufFBhgVaufu69eGKQ1KGX8AHd1qCRfGBv
mtN8OENju9VDQarAfPR6yZjDjhU2UjyzxRRv9/e7n5EEb296tI9M9SDV08G9G/im
DYQUOE5UnXKY+AcXk+b10XfoIkDIbB8wtUp4PIDq+zFlsi/PmmYw4bueSK0AoHEj
xg34RyATbCrwKNAlRZljBf239hmkOGw0i//k4oE8Zjb8S6IKqzs1qkOk1wBa7PW7
U0um41uFXKL3n0n6GU6u9UX/kB+AcPKw2lwLjBKYzU8LbFab089d5SqTBdvXc5d+
K8+XW+urSshS8UM5yOhindOn23DZr7SBXvAH6gaBtgeN7CWZWlHBieC1F39LRg5V
QlU6wR9z5DoSMtpiyZp+ULYZs+5wdf+Yb0gsD6Qd0Zw1PD5SHT+0+C7G87iX3Q2H
0SdsWeQsT/hbt3S1zSzXiDWVTMHJSskkW1CHSNNZT3wPLtF8IOyD+LzhYloq4NPH
VlWW9m4bWw3+jAhLHNdfFtO/bphlk+zRAYEDHVawqp3dt2sUdMBWuYDkYzNibqzE
3sRiOBAajyyXdGGUB2YGWSFypVGEBexAm/RO0xYyyGoR62awH4ZBnL+NPRdYoCmi
AEhgyL8T9ZECXhh1ODM1H52hbQLS7DxEi9HHwqdnOOIoGKiU0Q0izh61T0d6IzFt
+DpXFJs8sU5x8OFNcm+GhVdW/bfJMsoe5RZn81m8BPqOA9Dh2lIpSeeXuHr1zmzJ
2MZUI6uU3QACyFvJtaz6H+rNx69B9pkd3D196WEb0Mywv6vOfX6so6+/Hux3IbBW
XGY878PQcWqCQXoPphaI61ShGJKvRfgprIb6qa+wtqLkUnTDeGHZda2ej7hdaepq
dc4uDdIXk0C3LwdY5v2ndHjwlZnQ7Pbsu6SpffEUZsj3FVTMMDpusvkMnJNfAjiv
eH+GNLlrjWTN4hG/9odYBSQ2ZMuv1b1ka2KIo0OoflEF5Iooc6wH/ko6bUFsdOvx
bxmG38VR8tKZUWHX+dtL6AS8wWdZcUKOfBXMZUygGh4St73L0m8TbXqA5iCvjvMr
Ixe7kVEzmY60GcE1yMgdIhsTGhT1EnUM8DibK/E9xceJSgunFr5uDt3YAmu303gi
CQ3RptPKlFhrq2cO1ZhCyY1ubVWInGV4AaJPTfK+z8PBkgZGSrxIFYIBXPaF/ByU
KBaqVI73lkt5GuM+Z9kWWvSXAEsEwfEsh7HsbwiLsoucdBpHzzUAEeC1FNcKXJX3
bD0GMZ5q0D+yIgfYkI4xDrUeSvhOSmY+BtOLo+XYAofw4uYBcROp7DRytSU+PneT
mpEp88PgG9Rp4bwBCAhp7RbYzV7jL/xskVX1OLAkroDOeKoU7d+93+sNKFcxc8Qm
OpMeGYWFw+HC1GbcqE2ItnnuvgLPxdg7Ltq57Xaocia8UpcLaxaV64QnpAKxaBPW
hJQa5W9ydc1NGtTwOHyBxI16UJFNpTderGJY4QxY6ZLIJUVDChsVTuGVzxkDtjpc
1SbDNWyRhUKOGtjNBXYIeOqF+KhK5mlvbju2AjJTj8kasAI+wMWx06mdxUNcMGiG
P9H2ITJl+2Vvp1B1VPfLsISDAgVP/w18OnAtta+OFSvuyDESF0E7n9x39iKc+aTJ
QUJVAjnPAMLGnBuGfEAPnudVzFjfZ3drPz2W3q7x0CDRsGphxRS7bm2AR+7noXB6
k+yfZ3yfzplZ4hjK18V5ZXlw7LnSPLZuFA4zxy1Z/tH5NCzVXMeBECBXsdEXlrxq
v6QLdKMaZN+yigB9OiABIfyG1Ryr3UHAhshAc8Xf0g271CTEkJ3wwiZ2/HerPWlO
Vh4DfQINsTkn6yhRB+HRX0+4h+wgR3p/bNfmVolCeO1wYJcCmBSswKDjsVFaE5iM
v3AA8CxuYuvWoaDQ+qO3fCthtVto7D00X9YRV8IfAuidV2luh2EZpsgSDu81VUke
c4AGtQsY9n2nprbeKjsI8v8LuLkIxXL/OzVQZrt8JyUZFHWXp30vk8TFP0rQ5OMi
vmMwdPp7lnYrmpWLyKXko6SQnV+CC+WdGgbr9Nc4Cf7J22ISBuUAlDprcWhWLRW7
E4mWgoLds4yf2kYfDv/pbPhnYrdiKX5+BIHNqhNW6sDhTMDKgwv/iX8MmWwSCPB1
L6dDtsIbh4AkKLy8HoDWqyaZPKVb/DauwnvwzSUH709FcP9tDqbw0xU83E/BnHSk
A5Y8hXcyECr2KmblNdPyUcIGrEDlOpExDXdJHWoKbHCX5T2d2x9FmK36X9E8Un92
keJTDd0PW9dmbcHwVIF/frzAiAnDBFFY+IJzsj/TrNzYWP3KHWzWa365jvjL3oPJ
d6pjTcOEVNYKxNGdewt1QJjtV5uOREpNYSN+tBqYaFZszOU7JqEE7GigorU/YZgU
gobXcoC+a1VkM+/bg5sVkxQESU0hz3f6jXby7Zp9zoHJopjQbgXfuUhNvEKBhE3g
QQVNERxYPOCwmo1Ya2JyBbdyOYFjvHr3biZ4wGGFUwVNplHDqw+EIgkllffgEJrD
KiwZrdOMlxkGglLls38tQPWSJeJOaSoveXMfrWuwTbzrUHbV6uad126Esi9YLBWU
PlBBLPnb76ol0FO/jJZIWm2B3oFufCdhTt/bsuqmSYTi4w0sv4iqFGmrVIrIAxwk
T9lIdXMaqE4otnrI6ZKYRLbpreKzllxNypSGzd2l6Z548X+VNZ+FzENCfNMPH6J6
OGi7ykbhJETrNte3ysvhVoo5Nx6BhL9hirm17feMRnCX1uWOlJROhmPV3b0i9v5f
vfEAsMHPjWPkqKYrendoPNh+F3ZRq9lpqfL6b/6+MLczbVBMq85z1tq9wgWRfiCp
AZg/hhFkyQOWoKNLm+wiMYb+0RnQ14/uvR4oZ6wPJsrxHp19LTxtIPoIIUbJyhVP
Y6rRKy1Upz7ri+gcgTrakfDOLmPZWJlojU2F94khFRBZgKOQj7/CEgrZwvY0hZPp
Ia0riFxlz1cEwpNFAbJ8MZvyiVW5HZx/Z3HctJpFky2qLs3KlwSqEo2qzAPEKbIH
V3KNckvElKtRqen/xtgmMVTyngq+7cN/0n/ECuds69usKAiknKfXasrxoSWuWaXq
F4TtaOZn3OA3kqUjwLKRUjVbCZwDnBivNXf7yRPCqupdQmoaie8OWv5Cg5Gvd8Ek
za32+XOl5JH4IFLhJW+6qBvIx89VzbaZ6gH3deotOslP2lwIR/rnx6pHyhxxJA4m
zzdg7UwOhpRErJlT8SYiEvOIXtrEXfaHMZPycY1fqiv3y4kJDo/ai9VryxtYPqcQ
wLI+I6IT5Yvz1PWk/CSsBOIrc307U6MeuVLH0/gQdtAWho8+CvPYq52CeIyhi7T9
LUt71Lrd4LNyrnulrFE3zKz2U11W+o8Z2+Na+zG+/7BMmEdFWwKqu0ePDFtwOU8/
wGWfSAbZBujYfwOUeeMh/cOhg2eFFxYLP2Y3/HojSJzudZdpQad8vMwCQuCc+MiK
DhtPeUqBZsAVz2cTN0HP5QM6Jfm/4dh765bK9TT8UTGCnhl3WScbEKlYPxbOAE7Q
DDFebJPhfhdYf08eEFASOKyxXBHaUXU+a4hL3dulIcI8MYrDLzju1g3Ets64tYnm
CRRoppMIOw1xl0SQPQGShKX0s1mGwCDbh+yjaOxjSk4mpjh/aOvQiSISjZrOk0xV
lFjYqrz8I5FY5auvIORpprk/sD4SYzqWY5rxk20z3hYIWLsSr4ny3kL0MOwQgiRS
tQJAMwdDES3ek+0I4daEl3aQFN04q0SJ7PckykwVQ5f/0Rh2m8FUlU4afgP2fSaZ
HlRTzK1LIHEymAAS8qN5L9E4Wcxf4geQCa9ep214HNzW2ZhITP2OvaD6Ud1SlCXE
mSo+ea+9xczRX/6JvZgQusJn9UsjLHwH9b2yc4Vsefwb/5j28OJ01eRfIOWEwGRD
8c79qw/qgDs1l8WNxZlcwqmFyGT3x+kJBJyQ7fQUu7b6msWjNfMQOuFi9P00z9Zd
Qx861WM8d6BD4EeaH0xAvI5moj+XX7BWDjBfKKnI6o0/he+C25eqi2IfGVqEH+mM
//CtmcBroneD0l0hCSN3n7ZvY5D2I0Jode87MFhn1sQA+28eBfCtGYO//EgifAS8
e+ZQdR7a30uANLXz70YK80woWb1ObS5lmkDzsnDeWJQW4jDoBa/QYLB+J4sToCwn
oZMtEjcaOmgdmPlgJCrH7hFvA/tKtvd2THZ6+jtUknTck1VH0/t/opEmety+q86n
HKF0QjpNPktT5KcB14XxoVI4mA4AJsEJojqNpkCUOI0W9/oGZki5TYp2cL5xbhcl
hdSup9HIIl7mU6lmRtbyR2fCAK932qZ47+RzYj/ib6dv/Ls2a0gan+CiesO+SXZe
tHsrDugCu6w/kwKUcgQh5A7wrRR2dJbgoyytPP9i+NwJUB/0cYLj9vZLzW4wbOvl
+cPjnK30npFGm/tTS/5iZyMi+SJVTfLAZcYh05N+WFf6/7hC4hR+CWEfiHio1XMG
jO1BIjqj95afgPvjSrCrcC45nFR/H7TIOL3s1HwNq+EBSCXESptwKhBRw4T2aIo6
K/TXazI7afmDR9FIs9xkPQOK9+cp28lY2pB93Nf+zsxJySrzr/bHy9tv/wqDndcf
wiqBOnkROR/NwIQU+1oH/Lx8vgxfJ5CRoXmU5+ywk7MLVKqeJlHF0P+kAdQVp/iq
mHBOv+oVjanZAhklV3A6Flye9MpLqOYVtuNjW3Lmh60Z/bzGgXJvv7QzX8mKTUvT
VbSOZ8kkrks0jRlplbHeGTMFHyt6+S7B643rcSbR4lmGT5YqzHCr2pt0DsCH6tZj
r/p8OoHWHr2QJDmH7vERzBpoDj3L/6Jij3nHd7rg6XLh0hUDlhJUm8FGoBO1z75f
yTMzLCZwNrOCwkrbF5mbVU/GrxXNiU6ve0VCWLSybwLCUc69j9Mg37fOO4C0CNiv
+aNI+p3BvSYEVr/f2iuCYAnq78XgZweojS8d3/xq+bAAnc/5dwH+HMYLSL0wXGqi
2DiedgBYwdF2TX+e28ZqCDlc6wrUqbuFlfu1g9q2HwA5u/cloKp9/8hkYf9VSkwA
EJuJGfRKkpj3kerVLfGOqVzJhLa0TT6cCdwcqkS06OkMmnCh9BiTobyXJwl6nKvj
0vxNcANroAlsmskCAq4tiH+EBnuk+fe/efXWkzkH7QT6Tr3YaVxX0G1P2kAQyl4m
d52WpYHavLGDy9zLLGnGDd7JFTiil0HFbl2S4eaRRvmxAV3e6g79nOuphBtBaxwc
vGYfHM6GAoydXylrDkfUU/5JKwRwJx/Pw5V69mMs/9z5L4rtrmC2nINBiaaMzuJP
U2oZwn6RCqn0SOmpHU0JOiTR8Dg5s4c3qJyTk40FIhugUbvWW9Jpv7CzMn9rmf2w
7N8Wv4GP/MWB6dFbnPxCHTLi9DbiW3yoGImjjPD31QVzHduGW1B1e+RLxPta78Fl
vNVUypm9nh5tsM1OY7Emf9KE+5iYKrla1xC9R2sRwwBnTzrbYwXSkzYxhrWBVcyE
fUV5lJLz89897yT++qUbZzEvXyXMAYoMaroNpSIlLsW1hy8e5i77xz8OStlUoDwb
CASNmixi5ANf8dHe3pUXDF7zPGqR/dBcFbJOftXnhylYR5/06G/pDQqUFjZ9M/KT
GahO9b4xcTjkTuRTIMJe4H9PeaXlV8umSL2gzaQ/KvzPSuWUdvgYCKZ+np0/skH7
nUUhRHVISH4rd3vZkGS4HL6a+7duJLiW7FAGRdJFy67cSmYo6f1jZ0xO9nvAtEaW
pshNIKd8uIMV9qM80i6Em5Xh0uYNuIbwNQxpq7HhynA1hthh/tGnL42Iecs4ZNjU
4GKw/06QxkQy0sM6Alvjpv79vzhEF+RjQaoZ7oE2m4R94lIwGh161IbE+AgLurky
xfRAUYh1tD26Q8lHAz1OFp/ugXiupJ1Ks4eK4uoxyrM9aNwYYiGU3TYJNJuoHyrz
E2CKhWE9ZltyE+mW4h2FaZhCZ8CqQzUeEkBCQi0DpUSzV+La7FuPHcebOeybkX3a
/jeBauuTMh5FjHc8rwD3HCArv7rdhpUK/2c0JWz3yDK+/K90Mysz/ZTgh8HzQNKa
3fD8M6NmKcVpmGnRzyEB7RxOZLr2N2Np1WQivXl2XD1Im+LsRIGp3V9hM8E0PKxi
O6s7PNzHUi/euXlnYza8jy20HnrXPq0HIty8fX5YQVU15/43S3cD0lreaCx046y+
Wk/p3Z9VIZBrzzfiv3REj+SXHOkbUMCg4wIECwTo2Z5+7dQuIjx2bWBcvR2mgIt5
IsvoO3QB/opYOBa23Pvi1OxVmOvy0WiRhNYJZAYB7i1hbKcEPXCe4TI3djqWatLU
eK5IXMQHW38AhmITCHoJ04HDb577cR4wmQhGhuz/p6Tp9ee2GtZyFD4MWwXNzsLc
Ok4FmjRk17HfLNg14qojn54fykZQy0iQmr6PiEF/OT3bF4vR7vBdhpo80P3XI71j
XRSPPOaZdaad+dwVH7nqw9V36xgxNbP93fGDb4m4VjKfI7cKnt0OqTzchP77qyuO
gnqDz9nRREyNXuJjMMeWlvl/27FuJiXAUpZGz7E18g7m7zPSBaC5b6pg99fgbEd3
j68gYIo89EK6oi2y9Ugto9a2RLYCR3NwYckbsemXZLv5/Th0Rxn+1QVL9vUe0nUV
x4n+NfS4+sU0HbU5f2kZsX023qNDjMXGl6tGjKXrJYzBN+rB+9cbneQFBPLrvGk7
kS4Adx0LyNE45dadum/xXaIDviKQ8DbsEcG7k9MDMWUZIkc1iQ8JQExMqVh5OML3
cDRA4siAiaavmcPsP4JW5dop1Lv2Pn9pAOLTEg0paRvr1CNtUv73Uk8bRb5lOyv7
reM0ihCw7anQZZ+Xte9hxuyd4D9SKjDg43eCW15mzRCDEofUOgu04UZuWeSZZzp+
nYukFmAVA27VM/E9JdvHUNyAUQ3C/StKfbinDjY6phUHaF1mKSfT55pjJRXei1V5
ppvFzZxiTUGGIm+n/7YUrh3yiQMu0pfYmydZYD26/Clr+4aA4VAhj8/G55dW6MFz
55up+6KYrYpqsJQ1tIATXfuWXyCTu3uhw8aELvZplbTHcLLYaZ6HufRCF8qd5WUu
wpYt7crrUfZQJPEAch1bSJePM4tjQF2UeVGsVF3NIDpjpm/xSQKCwljQh4A6ZUA0
Kg5nNcLdQFjWmbVNiZ54sp8rB5UHQwyTKEz34PEiYHfpDJDxnGFBmXk/Mlsj12fC
B8djs397jWs4XRGPniOlqxOeDBq3ELb7XiiMg0DadGJ97Gifh0Od1nZ+JoCdlBmE
fv9tmzP715XaPhzyYfejYeuhI+KPiXs8UFpe5HDluSlmlxf+B60/m1Olmt9DL8VY
qfowubAw6OuzRT+Ml/JeIS7+h1J60D3OW77/j82nkM4YpOshIjMGd5IBC59jMcHU
28iZkC1PS5bPc7CKxnSVdKrB36XLyGHG9pF9osm/3T3U3+qIVisnQ4ye1NeiGA0g
gAr33IkYuzhA5n747kdHHVL3cfS2awyOP+yuX55+4A8Pkm08cuXlFPvBM9ZbApGb
1rmNUucHxbCB2G72Q4n5tBI8a8+OwdUHhGyhllMgWQF/SkAx1TNztmWdUwZIqplX
s9urc36qzkFNaUjMmYn8PJMO8BYms49V8/Fo3l/9CEobhG93t+RnihnQlVOvQ3tL
N0L+sMDXLV1jzk0R1giS/IjVmrHHMIpsQsQYWYhnAqr2jIaIf8RSyp0MWtayp+gh
tFtrBJmXovpgj8ypJdjLBg5Eeb0rxlPWK0rtTVDZDKEx1Z4Qbu/FH7f7PW0WetGV
hEkbcFBoVR879w1sbuws1j2Z1A6ohE/uSbX7DnwXte2/ZNegsNwAtva6DMtVsQ2b
4sPMAbRT3UrTqI/zsapGFwbzf2WXHFnyHUFaJrSpswJU0J6oMu1nfgMEGMg65YIg
pXI8mP7ZLSRiLFiqT6SWK2bc8PMUyHf/mE16DiRhk9HpdZJ4H01s/yflVJt3r3AH
FboV00IqCVaJl5dER7AyzmVM77PkG0QiPrhPpe+mLCbyV4c/ZPNLU2649GtoWEfy
7jUhQiq1hdihpKRxhYywrrUpVkE31H1u7+qa+WFDotQ+x6n157eU+Fj2GTdzajMS
zt7AOp1Adid/KTedi3z0zC0hYds1712FhYMFxl6VWR6qjzQBMfKHHvNKhRXJ5R2i
z0KnFmXhjl0XQq9ljIZwyE8qCH1a2R42i6mx1p8di0fEL8JVIPjQPp2ptl4fexl4
AU1niMiXGguxWaTae+axpsiHSPODdpTPkNpP+KbVd5T1gQZYm6Sd6Gn2U7Kzls6L
6XqNaVuBb1GBIo7q76Rrxa1WLbA2QmUI1F/b3Ew4vjF6cdmYQPUKZYOVbwSY+Bb8
nvsni5QH+ea38pGLQZBIBFDPkYtLfIE3CIWgrXPhBwxlRao4z6VYKvFWk6l1183Y
rQS6uDnUf3q2wU8/FjAUCDzWreGOK4fusmxu1x4555vIyJ7UfMJkrrTp4SiLpHa5
cTAB0ahaNADu18TQRldC/jXbJE2nithhY1SBHRRvjWur1KcBdWxG6i1qdCeElHKx
EOeFyzeIpRq1WOz0l3XajRo0B3ShaHNx2BvPb2tCdN8wIP2WffCrwF2VVYha8Cmj
CWaxXZBCDYifVFEF6CgRZt+zJzuKjKhB13QcxRndpte02FpQRQNlYCfeItNpp8Kj
qzsUz8XyXQCcObpF0zsI6xUlE8HCFU9CUaUJ82uk2qUJ3mGHkSK9U+7dmkvUdKO/
BaBpGeHPkbVBwYpLRdwEvkWYO99sLb6TYzECum3iWGGpJTmAki5kVKv+DUcLOOcG
+v4QRSuNGF/coc5dR7bXtzj8q/ULRRAjVkbsVhL6mJLeEKEZDen4q0Un4/j03Ca1
AwZNZ9Z4AnuS654VZqE4meHRL3meuvZsMZUohMPrllRoNpXSFWsi7aA2g1TzjmDq
0spxPeY1qu2P4Qm2VrKCtoKrgE2IdC5gokvqU3eWiMp0/SV3f3lDn/0cqfpU7s+n
aJer02qSeO7fxntF1x09FxRtUmXwyRCDbTlqhw2Smu0vbVXItJ05krGwSpDvyPgi
h3bK8uEgyeEmdyxor+p5jWdjmT6yZTOyLcsAC4eh0meuNtQUzonFQvIJgEH/wtu4
6MtqeS4eETA3RGdShyNFbDf5gUNPCah4qV0Ljzn8Q/y40eK6yTYlVe1mNfj3pQsn
BpNPkhxarJdsftzQulXz+zRG1hGkZ153wXBDolRbotxxKJbZmjv13G9F71Rv/oAN
PCfsJfcLtmaPUIjLDzv9HBMusFSNZCsXPuJCcTp9O4KmRxXgKzNeuU6BcWoDa4FL
vFBPOvkNeYQh5pt5loNO99k3hJ/5jpLFEvTmtr2EAA65XnXinhL/23QfI0dsZTBW
As/Z9dAPYfXyKhulguSLkHEBxgiKBCaz0OU6hv7XdWEuVdhfz3LaMyQ6rMwT2Vrc
Lo70s0AFqdtgGfEMgHJq+RoA8eL8cXrvrg8uoVW+x0Zy7luSZs9x235CjMihjQ5m
aJ7bL4oHD02GgABOWIaNhl220ecua9sMXQ/uFg/7xGOyZ6eQGZLBleiGJRh+KR7C
qJ/Mhl64P+GxzOZ6r4HKiZUrxzc9WyuOqJrbSxNa7GAlt/f9YjGWhHizR8VaiIgU
Vsjd6W3GdnEdPk9Abzg1fS9jxUeI+yuPadfysPHtf3udUiXm4YIOrCyd/EkfGgpD
1KNev483RbIuTII+u/fGgouXeEg/g0jiGfwp8yDEEK2wpyEezinct/XPvDPWFmM9
yeGndEbKgqs4/GwviZf8OWkAxTxhsxQ1hspnbduywepN+kamMrVC5uPlWXYSqeRM
/wRsjioLS1JYXz/ypwoo/MRB6Y0/Af+G1IFQJBtPSUJ1vbNBzK4fZKbngVAeoRym
M3evP3ZgBhwhtHzxfdE6jfDuKQZBWxBj1yVg20/5ExIJjc5eLGHsxyn9SO6jDe0F
RLdUf+b0ZJL2FRQk72Tr9UUyRkTawNTuNr+XmLzu2/BAtWyt8EULVTeoFkKnseKN
d/xhDAQXTPLae26xxtnBjL8/iojEckKzZogWQaeZ+ZwAosBp5NXoCR3xn50RT5kb
Vpd4rx9zJN2SnThG1x++KKdYAu5FAuRXU4I1OCoeI5GGt++Y87soKQoe4dd74r4w
tLQXXyNdnJtUB0L+H1bmL8fK9/FKHHdVPG9xCldErMUf6cAHuQ5sebEqlIAn660u
UFakMrDOB6KW1YjZzlltOwA1z93P15zCXysbA2ofFgVYA8Qm/Jxnw7fvhDvyYuJN
u07Wb61KQs6mA25uAI9Dfq/tOok/GxwVmnnM6ZVY+241gKKqpnghcYIxdgVZy56G
+Djv9pDuvZAl5eNPW9hjaxL4RpfQPtmntgeOtEU5pnwEJ4hYtsaya5wrobQp/Stt
2IEHdrQBihwtglJhTgbJp28m3MOEX/cM3PrxRGlodzkbDvj+FscN5dNtUVZlRCwn
8FJ+JbrHMp7In8UtuuHmwLxGeNjy7BY5570G5cHdh/2iE95buLJ27wmdoi67MSp1
Q+57zHgqGiQ/IEVpiANdg1SQE6fXKc73WxgIhh01xbXX39kvCeAFy8N4kOlh6hJJ
6YI/M0whFhclPrC1/qtGQWdHksDMIlim2iA/JkCTOuUAAQx8VpcM3IVJfVEXeReA
Q5ycy/qh2/N8WhImbKu05rOwNwIoUznZzDxJL0uvhrpVYkhZsCPexm4rxWw2MWfy
/4zAzxH3WgFry5a7uJFBXGbE6NjlPdpZG2EpYnZL2GDCs0quACuPyi5/iEDLJwg3
cvmgY3CSV20JrjhL0rBS9rmGrwjXYzmPi4jVFyvCebHR7cEtqfBwBCqVERMPtFT+
sPc5La3LDQIZFGXbdLDcJvsOizboYncWD8E0cE4nss4Pa0SBrtBChH/yj+P8zAv7
Z7jYb6noL8YTTLrCQANdb6z6EzwC865J4oJCLJt0Aj9N63r8naZzLHLxkkbv6YnM
tL2xMKySFSI7+BSAcCxdssm6tEZGE/L8gfuV8z1bf7fdVmGGDsPX4a1o+JyA8LQS
Cdu0VjMgatweMbATGxlFeQ6/q/7/iknLi0ucGcIBCnOALaphs+BVMAVsOWuQ5dIb
slRHpL/kY16mszR8soEKaloUuc5/+iHsvlPkYZ5MFuNDRigtEARF4UrfMJWSVo2m
W1xwq465f3RJG3ZMuxKSKG4JzD5zRaNPfmu3JUKTap/f3R232qaspXd1vP9TSX6Q
oE7AuIfRKuRU6xmcjiFHUzwiVkRg0tmviVPMSI3TEQcUfAvCV/p8VHgcynoo4Cfi
Qv+S7xlWAfQvkIKdu02kWuA5UX5/hbeZSI5IG2MTCTmdbg88rFgwzqFeYJ5z8w/N
Rbh2SdHdjeQpMLjs1w4WUALcFpwQdZwjhFWbRscEvxLG+w98ST5pYseWyK3FOXoB
mDIswcTKBuKqKakQ5a2rmbi3qTYqIvAGuHNzUfK+kNEw61Dr5SnrIngGvjf8ir7m
ciqXLl/oJfewVdxw2ufavi818ReqO2Sa3+9luifBmPOfcGA2HiFdhu9CcecMZHQi
X0gx+i6ioP4Y1WIgohxTTT0zYgV8KqTU65gy5LL58QhXjEKTzJBtbOPvb2BnZe8i
ld0q8dMyT/lQL2DWmRp1loF0L6U2jzwQgQrMOIJsWSIJZiuchYD7wLsauvMOijbY
I0C07yGw9OiTJ2qtfitleX3Bsx4WnLfvha4SbGmXNmOt/4lUwNEyziT766kXYgfG
aSoRikuRfikINrEucJs1V/W7sW9M5SIKkgMnagIsMoFO/2VOL4IM25AlyyJ+ehTI
LTl1DwDENu7NVYhUsyBO42Vf5DBFMk49Aiju9VOUmgp7LDGBh/V7OtMSG7W7497D
dSgPmNs8RZuTOUdDJygnYzVtSUbAwPyatQSmaEQNH5R1mb4+xwVV5REAyrOYaWND
60p7kjRl4psPsfvultVB4TendofMGCb9ze1IAIDR3vsfrWLDNjfZCV7SkOCq8DD3
krDtdnRt2oYbPajfTNgIbr874JMU8eQwU+ZITMDXBP7kSOf7ZXVK6UXH3wrNveSn
ES+6X21gsAo3U2r5XrBwC/P87zs1Jtd5AXvMYXUgzHv/tXsIj9No5T4WCdVIxOlt
P/rLj9/SNXy32wuuL7S6bMn//6DkiOhThvvPA76fteyiVCeHbFNKjqO4iMLn2U5c
yUrwVbYee0We0WQlYEH8ugMYkKagrYRrbC4MxKOAy+Uzwtql28Q2oV1g7TT55zHn
aWz4OhCdaMLd/wLjnLsO0zTQdPvA5JWrIj/NoX+Tv4h/2UQixEVDtHrHKqHZMrsr
CyURirl30b5bPMeIh5FVCdqbRjQdGqmFGv3jw6il16eE/IQa+YZPuKA6eUNErrRd
rDBU9m0cibifmuPerMZsM/7Z6juCxbLVNy4yAANjZUAkxZW23kRCEN6DyOYsGK9i
JwoL9ccDKl47rHZvhj0V71dgEMACaX17xDg60j7LIl+T1767Yymf22G5NHrIyzuj
+DJsS+yS9xbtLPp+AaaOshJaOoyozr8ePEa4W0yBhk30K5FhY0wx1m2r2aKZOvZp
RYGHA105yPOvo4yYL8v/qe6/JqPQ4awYkofeN6ytvJNiO5w3+/KV8FEpk9bfNS6O
UUXBc7o+cPrQAXbLqj3ytPPeG4abVSsBrA77q2C4kWHAjkCl+IP28ypvxlJzRRxF
ypaUY5nTXwItykSndQMf0/omHGZY/MrMvdsvr1XQZYyO0d5Smx5nAqQN9Dgmp5Fi
1m8/hqWlkdjnNXBNGxy5RU9uWOFA5UluH4+NKIVozbN/xNTCa/NQOXTqyX15Ilyv
eZYb0CYgdL5IhoMZBAa2jF4JXiBnDZCnXQW15AJD05B0FI9GfhOkEKp9/MbRO8ni
sXGJuGbid5ocd8TNwh1QM5PNYu1uEel23mGGlokOoWylIzgD8Tcwb7it4p7t+7+B
mm/HIqw5C4QTVYOUxPdhFHr3Oz8zUbCjuviH/omAxgyshH8jpEzVEJ34onu2MHJa
j4MU5RFOuFSfNegIyT5OOfIQeKjnnbLWnjLSh6aevN9wj89YQHlL/3nuFAIyBW7X
RsLRqHpQQ/UWP7AoFf8GvuUdroEPU4U8+2bsc+0bsScUiKAgwYmKYENlMYdnmg3p
gzSMejbRmBoJxfi8bdFG6UeRvI+z+ou09j7VPOu3SiqlZGyVBw8oS9slxaYCrdeG
RsuQCTNrkTxOu5BXY9NZlAVPtIcrINA2jzeJ2r3DbiMvjkzENohi/MtEOl1WojtE
T8ZF/xozF4Ee7dXILxDKOh9Z6HHFdevK05xfADh36NjLjcfGhprkDrU6YekdyZwk
ufUj2fetDhnGP52o9LMeJf8jahG7Cp7kjE5rl376VHQX7CkxUWDVwntiDRuaI37X
a1k0nZP929FoVT6USd3pEt36YShVQkefnsgEY4WHw36lsX83PaIVT19Kgpa0YKll
J82RcGyYyzTpYaEM1XNCBGBB8T+3ObJxMATn8CrPdxbq3Ife3YLGFw6hYT9K+6iH
dG6uQX8l2FmV7g6KDFCw7GLEskwKdb25sn1fKCFRusVtA+EeyzU1uD2CrPrxDcYu
zQ2yfS6v0utBVrjrOn8l8vAM7untEsHaX4x3oOlgg7KfV0ESINUKttZKULqjxOez
4du8S5tQ/5CO7h1Dxxm2KjgZdQ/xsY2uaR/TlWdj+du/HCYGwsP2mWq/rdLMLvB4
TuTZYPYmiIkJAakcGAmt3zyNqypitrHEaDMjvnFFpqsnTW/yTDa4c0B6+iqWTLHe
Dyb0u7+XX2UMPp+ZkSUo6VMjewYqVajokSRuJRinL34H2dBxeHXEsPTUGNwTTPkE
Alb5Z2xIsce7BkSGq1WZM9VDDc9eXsFlYhnWRAZB9aH+ILzDbdk+hILjgStKSTVC
gktzS5ac39qQ/eIQgr2zBlAb0r90YbEjbUYOsOfblJcbwDDyxpoplqDm7+bT5wzM
HIRHoLGwxp+iNUPLxua4bIFkxO0nXd6NeTYhDmWsMCtbeq0kXUgraWhdtqmIUExc
bwaSCJfsVP/mrEyz+LRNlAXuvaqe4jerpuilpXh5XRHsFVwomU90M9CH8GhM3+Mu
dokIh4W+hQ6HE40u03WgS1c44SIQpeYzgZ7ZnYNov0XVF/isVQqrz4MKACt+rk36
pvaZluJh+6k7mnTtD99vah2yGLgo1UDXOvnrfhp15jWg6NXDMsfuwPa6IrPR8ZJn
6kFmqDmB9OD4v+H1FMlwA2xAAJTMj9ncZEwzrGOuSLhN1xpxDlsIBEYPXE4VXA/s
WhHcXRdSU9WkihtZCgE07dLQSkdklhdwNS06yOxGIEveet3RzJ93YB9yPJP9amRA
j2tSK0tHmkoghizbuqw9zAfnE6twNYfoMWytUwO46Ol/hB5ni+yvV+WcERNy3E5E
nHUZnkXk7Hwu5YHftrbbiv4zToAz5DEEUSwZoz1xvyVw83Jti7bdFhW6ntiGpTUY
6DCQhFLvjDEJY1vfrXTtZOVVklpZYtqnxGKimVOv0lMR8szeh7gTSsBa+ocYiMIF
KzLIbjcqc4yAlTBZPJQFOcn4sSRZyhLt1dGbR31fPCu8QWuxn6s6wEMbtzFDqXWB
ySn803ckck8QRDXNIgp7UXphSztbD4RVm9yShvOVjQ4MzWY1MBhg3d/OSOaMAHqi
hbvFd4I9o+oIIQA4cFKqBg0JBc6wt4MrYsUHM+h+KPxomwYjazOwJPe8Eie+jX2W
t92KrDg/Vpa315CB9tAcc4F+uVUhwZ16y/El4qhQ6a1YpdQLT9TLLk+CTSLHkl9C
mSgwaGn2wUsVtvwk3vqz1BOXT5eJMsrVmzFR/NjiJXlMh6ucKbtc0lpy1FpI2W2F
y1gNImd1KeSG81n2fdOKRMOXVvRg+zqOr8OdUCYQFAIByexAPSyrdvptRroB3e+A
yMpWnd9kXt871XRg1qdRNH/iFMWd5nBT1nyQpkDexaqL4deFjS0HA4lPT+gKYss0
xQm0S7Y7mIoGd1+Uh4vCls9j34jt86WlwdqRtRfnud3Q8Y7V2PPm1J8Lo8Q3jgbh
mCD/lNz5tLK11MfHip9PHSsvlYsxDoEL6Hq+zeCI8CSBrv+XbJh50HNXQUVEp3AC
a+fmDnVwagDzRAZxPubOHoFjn1dlubwZi2C5uN2URjVUrPSWBKz4VDalWwqZdgRv
vSyUF16L+9kZppBR9w83wqvVgcivkqZp9HzbfQWzCK+ySKqQGIjEAVsUpqn14BBm
qK8xDWv5/32Gn3azOkfC9oECL7LF3IgsOirQisEx/34MoT/sCXINa+EopYJh7ZpG
VHWlbg+fB3yI549em58wCpK8DNPmTBcSKL/NmZzcsUF9wAZLHrULKRcczpuXaGwF
6+HFNu/Lb1cjQbal78CMtMYnRlyIbFmXjwYVwLwfhNtL9+GS4ajL0w48/1p7YyQf
Bs9VpZioiBrIsmqt10UXZsBgN88fXL0otU3Klk3z9KeXeHmcsqS/SJ+YnLbRDOBN
LmkdGGMSWR45pDJGgXAMekjc1u9DuymEj26hRssacmJz40vjOBH2cEvXJjE1ov+U
q9Nbciy9pFY5nDsGmaYV3z0Wj74oR/zhoA2SCh1lqAGOdgSUz77w7BfRasVKT1w6
YeP9Dr0ho8XsLK03/7UMQniqSJt6+eIRiGuztyYrs8z9xNz/v1yVY/nYNcWnr5wJ
wP7gY5m23K2pcSNlXiOZ6LrCZ1hWrnjGsCoao31G+J8mV2lhHInUzMtMgM1nt+2F
4zbxPko6T7pyXNha68UPd/acdJRR6Mn3/BMuSr4DydO3rXlYieR2mirgR9RAsajw
4+NIL+9KhP8I5c0uJ2OXk1cCyVrZrXJUH6OHOakKqpbP20zttQ8ZQQCSFrWk2A9b
evPIQKv+a+yNv/CBZeYU4P0qcPPgkSXFyPTTmgVSD9VGr8F6OiHgQZTu0GNHkcKs
vQMQqeCpnGMWbG5gmCgNqAGnoEnBEAwmb7rXdEqFgGGZhoVdxf4N9rWoO19UkoDI
y2GOBiwLJ0yZNQi7dKdt/WiWuUdzA45pf4Neqe4f+odi4rAvcjI2TqzmAUpB89AF
nuslLMNCwZusrXAaE5FTXz68B+vPSaWaYJbWy/Cr7ShUU3+sciLbxlb0ofbvMHVt
Biy8XEbDx4WIBVSJGBoAdSLQdCoWpHKmh8Jx8cePujqt76svGx9WP5OyoIlZqFVr
YmYPWE58qQKMbNB9ccvD5rwhhE0V0HntI8f+Qf5BPp1x/NB8ZDHjJ7eqgrkZ/Hr7
XEbhTBPhYle2bHNl5ibpm97ZH2OCAs6LC83+GdHbCesl4f1sD5G4SIuqe/qStJul
ZWAMdjmgtpWLP/go8foZJYnqCUf8R+/oUSffFxiPfy8pQ3yRQ2P2RrpcA1dRyVSU
2ws+/kzATmRUMn7poU9UsTwogarrRGWvKdg/QkxicfpWwsMki0dRfOJTIyjE61wc
p3Unr1lPyYVSwRMv4e6i8K7dLSyWQvTrwl9igVDku7yH2AuhlirmGOloUvrRiPQZ
Q01l0q5kO3inqVRShz0ahapF4DgR6XS25/RkLx1bllD6yYXZM1X6UNGFAah5iD7L
h1fLKirzi05sJ6mSmkylXmhmChvZ/6ABcVoPtCOpsk2ijqzTNCDGE+rnOZ9d7QBe
asrJDlE5rheFl2T0h3VgtIBdvPtp73abKoHi0hjFjQG/XTk1wLHT7ZKz7J9vUGWd
hLG9OYAl0aHI3/lGoSfnXWJlreatbLNGMzJj/RqfuzDK62SPX/PR9POhUJEJmC5A
G5C/+kWlD7X//wbfNl2Uv5p/XZCpUzd+1zrqIbzBKdP2DjVlJRTQHUJ4LBvGttMu
6LlT8ZouRF/KuKyARxWQcnm61iK0jROzzCrzQVGrCALXlGsHREK1P4zSEOQ5pDyl
UuPHMTRPu0xr5t+pdqYvwVQHf7dtsu4WQ8syc3gmTP6u0GzE2ydyEOrLw5eCt0nK
2wHZOoXMewKIKMOW+cib7z3pxB3T5sMdCERqT8VdAj1V0OjJ3aFQdA4VuIEI2uEJ
arkDG3YEgLlSsnm8tCBTY3q2EN8cztrICDfezRAPClxNQOxUnAjhC1P7LOzfPu/i
I9uVg/CtfL5f1eu3du+hucMKx6yC9Xln6psAucCiFDPYiJ+IQfH/H+VUZI6XzAQi
jQi67eiVu8rtMH+PCfEyf8wO5WIRxYtJfzYgZllAL2t7yzKZIxsopD1i2Yik/xwu
OXM9K/8VZs3+cusSoRr/8vX8L06hSSlYqqTEwUFWdgHbvaUB1uFHTnAfk55kYpvW
OMA8G913Cnz9ZIxCw77P3nxHEwxewLrd+yoRiaOBl/3tCd869fbSEtb8pkdNpEXG
ja9oUWEHSNQGd0EvXlx4i+LrRl9O2O3CPSKhb7lBwvNTrSk6It75kGUYqYmetwB6
Cc128ZbsiB2nrnsY8IJjIHmaDzyhkj0ufffx+xz5bdWUUdV0y9hv4+kaD1XN0Moo
Y6g0+rkEkfNkK6fVJ7zeIywdgyn+TkeFqZPdoVDWSmq7mFi7ORGG+Koe5rJLCrdO
W2Nq+sy319SZHMbtO4YaP0YCzgIGSSCCxodgGDHNJHiLK+0a/8sLiNQb9oUDO668
MZJB2iaIWo6FaLh5V+mG2cG5A0ISTUA8t+NQL68ZM5cjrjU90Ozm342SMU0GXbh8
qfD3Yf4gJXrHVpGTjfp/qqb09XH5BJj624o3NiBGA9fpNbUXCCehLIHv1wXRyC0V
ZzSmg5W1lPKIZcKDdwiKgSfWjlIpVB2eB+M3K0Ts8v6Mf6783+/XrB858AoSciwp
iN7m8nx7iVRT7O//KjCuD4ehAFVrO4ByV/DmAoo9gU80QRYruElw2ZyX0AqgLxY9
duICHtdK+4xAxRMs5KqQ73kM82npUrOXbgSm9rqP5bqhuV+fgOysUPi8DJpKVQm9
3vlWjxJ3SWv3IyFV9DsRF1Y9zqgGtguZKg2KxK+LFITCCpEKMZLtpTLcLh1ZE0aL
7hH4+mK4mG1CYaezCipszfsv/L+ahzp40M0hjiwiT2xHHZxYyPMiuJI3bBD4Ej4M
fKvYNT6D9Cd1Pugbi8xQXuK15MpmBwXFxYnwgJXC9cSc2C+TX9364tpnTA4FOgeq
XlXwe+elqTmwQTOqqinvwLSpN0MrnzbagzusKyopBrY2inD/I6W2pPibZW8CnK1x
IF8K8qmeBUnx3Lv69+kfWqx5bEcO69PiGuPBQuUOd1XLDYBzbPcwVceE+L13mcv7
i9IFfiN7qiP/ya2i+ftyRvrEFOsNBp5FN5tLoMFYjBuJISH+K9y+CI8IMjSLldE1
vUtdhW5B3+b+e1zs/NyWE3kyIKf2iu4wIcM3GC1M1bdXrYfS2y45EUjqYNhn0vgs
Mm833lyCh60hCeXQ5y1NbHKgwInmGRRZV6IKYZykV7d326z6m0z2ybL3++HZtqWX
Lwm7MudmcWSHA3UDq0HTFbpi9TNnkhaoGQ4KF9BFpTpf9eV1huYbCldJrs/NEIC5
dWq20uhwwczKjvRSKp8T+fFEZgVwb4+m8DaxJ/Y4vEV5ejitSnDq25rN9ZEIIv5d
msGNr4z30lOgfHwNMBjMtqN1LCfN+4aiaonKHu9T2IZKrIXFsujgvtomCD8Y8Br/
gKVfn4G88U+pRs3/BfuiarblGwnOk0y52GNzLyPFmVhzxftDkPbRcvaQYPf6Uc/Z
qyyyeK/wlS2vDF3YWxlzTqBQ3+HqLpCcwxzr3f8jXq3netbedMky0Ald3DrWNUMR
9kOBtuxF7iOJtz9ITFyodOcdLU/T7Q61vc4dWLFTP/7VOYe8/kSmof8im9PgYSvK
vrCiXbHUZIDavW6lU+dvB1tQBT4wb/pySidqekiDGPeGorwGiV9J/tVo0ZkUc/6e
QlFrdDKSaIxWDMgDAnx51JY6VXqD771Jkm9O8p9x26dv7SJmczQ1pa0C+E/O99vH
JaV6j9G2GWWkrBZhUqmWgXb5uMPetDXaVWEP3Zv5ze3mqZ6lmfTIWrLV4wBYvPjP
ww1i0gppHTVdZwfMX3O9zo1OKABBI4QDB1YHQoNZZ1ZQ8nd4kXQ+nRclQxyjbJ9n
VciE59+j8Z+vID9wPVEOHJoSXUtql+oJFC53qccYqK94Cm0l1+A/RLN8eJAJWZPM
JVzMtK7V879BWrZ3T9Zwk9filBYftU3YNDeFiEe4XqmWYbEKpiVO9nNQpBBHjMFt
suXCfxx0KTVrVTy+EooS9wRz8FvShtLxigCwuwS+pnnoVUvLI4F7ORZrAicACWdv
fgKDqmZoqvRyTg77JpTZpZt9jhf7AaeIwT8FIawqytxLejeT0bYz6PygkiNobX4F
tPAgkQnpisK08GBTbUU3opAgqD5iGsC2rKJc0fjtOOegvs+/gcT3V/1CM64T2ty0
HqxUtMNBFG6kavX/I6TvcqerDivJ3eMWMLi+B5qsxPf1R/mU+nk7SZHhrLiNmjOS
SMmGTO2uaprvt505fPA8S9X4Dya7LNuQ0e+ZQIOzy6ypj5/2pERfiFCidw4JTIJH
0YJiFzaMt/tNjgDAdgL4mfaW4NhA49GTAVE1SBlQn2NG0Dn0lg0WsqOjMBMKQC/6
phtr8CRgLZIi+kbn3VR1JzuEt1rKJuW3J6ZaVCFAVJfcr/oAUluUk9xVGjyZQ0Ja
iYf7OphcVFBaorEoJX3hiBulxMP7Mdz614ct22n3symtpAKLEXcBgJ6y8dBYSIDU
o8TDUBAI/zqd1NethqZfOrVbrUVJH1T20LqTItJA230MhxlQbRvRZ7j5DYRvDo/I
gNWoslQNRevGbIz0R82EOvp4F4RtsG/B5o9w4wkNp4XjIZrD+CKie7Ot0vqwQj3j
YpZenKFSLk55N9mUpej+tJ7WrnT5ImsB20gJ9Nc3omgOmkWUOx3sgN1cM4A6Eij3
2fl+i6ycY6VuoJ5KEePCV026Jk4dBo6Mm0qdG7CLq8Int+LWDcCvn/oLHeGI8kLv
yg0WaO1rLBhwwBOQBr8w1KBdUadfq3dWLE5wU9qfkdRw+5rT0pbRFm9U0wDrc34q
i1KYt8Y9uV4yGzPwCmAOWg/xgc/8dU/Kz8gwQRirx/TvqEMVL2C7E/xwNAg/m3FD
9Gm7X8T+fAF4ZNNHncpdUZLnje4fo51l2kvmyMJkNd24vo8ybUagdfLqEm0h4abr
C4XB4bwI71ddoDBQvUqzrMBBcXV2/kaB7Sx+8UecdQaax72dR/pLolvbeCHlEgX3
FL0OOcHDe7Ka9o/mkm04E1/u1t2XIyn0W/HP9rWVX9F0XHzVmL/AtDr9l4evhL7v
SUmhrJW7PgWmPEQ2VqeeyUxHTCjeVpdwSKLEZhWQ/Puthq/8BRxltbp8/FpVwAnb
+CTsAeT61WMqZ2eKkK5pn6AZQKXYJ341Hu06YljDv0UugiEIB5//eAR+MrCtadN/
Sagx0iv7H+pg+aKse2QRtgDZEyUuAdUBUaWJeXIWzzgWvo5RxU1va2CPQar86gja
P95hgLsMlPiwCjvtOqorD+e7dneVGTo12aLIROb2FKcXUjjStBmnCt8y2187cexi
fyU7YpQT7p//xq9OBiz1PT6hDoc66RXdxkYYXjMYzU6dxJbOQ4QRz/zFZqA81CSF
3G9UI/dOQYLLYSNx1LDdjcLLWdGBZ4L3zn5BbwWGcby8lPTE/QsbdDRnOWFbl2Y8
PbUIjWGhq4Czp1/Za8FCnv/y7GShA06kiD4D1x+yx34g6Yu6A3xM6ng8S0VO6owN
vGSoCFe9mTqwlIdwdSGA2e3p6wixllLVBtgm0SOR0tZYyiYN7zKyVU8h6wMryTVY
HIjB+rswrzjIWIz6WqyEnDV1g/mXkrF4v8qwClaHi+m33VEwi/rAN5DeCGGCwR7K
hKLmgYOrBU9W6+E3wD82HRxKHyKy0rzAVSKODROJ9uW4p/9kXe1shtQsX0Qi2Tyt
9qprTZxXsEGrO0pdBKJYVDJcZhWY2YrAC9ysyOmIyYoGxUQcQETthybIGlgKLy5d
zOFSasRNkklQEzHab6C1emEfBTbWnqq9AnUeH88a7OP8EYz45A7r9i9Sxb8Fkeju
WZ0PXQ1CbW4CcqDFrC5gXL+YRWBn7CEdKTviAsF99Jg542ZJt32vFZz8/v0ri4E5
Isddp9QfyAXZfgM13ANievum3C4fE/JevmuxI7wbCAF0TfgWSbMl7YuXFGcQVLUP
793TNQ0oQ/Iluq3OtEMOKjzgXfNT25BWO8+HsxpJjCskLq2O3d2FfjC+SR/UAy8Z
HE2kbHVIHY6l6J9s1DdAw+XZV1sUi4T3N8ULG+E9ltWVsG5DMS8Ct50TvMG4VXTr
cxffMbWYhC3+ABLoGOnM8H3bPiJCzCEerfDeNNXs7YU/RJqwGCafjprSXszJI3W5
8DP5EF/PPG0MclhRiFilZJ70KiARSAjk+0hsDhsHDHUd/RnOHy62aLQWfIK9rjZ/
Y0Y3HtbVKAEaWhOUa6ldtcgbbjBNQDYKt0r10KxOn7gm6cXBOKEYicFrUZOX0Yx4
km3V1LWRnkcmb9m2yk1DFra0WqrEWJ8W/3DefRJjEuqhTDHVAPuv/DoL2vLMKZlX
19XFaShA2StbcEJwilTtXq0UGK0HFEGZ0e0GSb6/ZIHrxMjOh+rbSfIDIb06a2VC
Hg/dH9pUheJOiYgaHXW37o19QV1WNSUdJAW15qt5BqluJSTXAldq3725JX7ZYkeS
swKv1kzj037q4hv2KRTHltcm9KuOm0DfEvz7v1wqH8r/qk3Tl9xzea9Lhk+cMOqX
ph4PLThkokeADHQwb2s8Xkm6+llgWhyv9HO8tvgUq4/T6PweoQo6GHMWgFcb4Qgj
vxrj06UejtXrO70wxkPyRMcLYBw6i84+nbyEmDM4dgomdl2AxlyP6SDrjN/uFTC2
UDIbE+AREjggHNZK8QVZ8sQozaPY3PT1rV8X1JcCLUM25jnLQkFNXIrgtt9Qdso+
zEpxlUX9ZkF4waLwRH8kvAJRZuQ5CWac3888A7DBkqF5MyfylTdoGFz+vcPy0SCw
Z6P13aUQ1IO3vw4oihftzgELg0xEd4CqRwqPnJneMjQ9iWUz8CBiNBcBi+FXYTas
7E2hDUxqowpX/CvRqYhPLUtcaz+Sqtb5PSim6yk9im2gY6XGHz73ipAH074FcX51
5gIDfECc5mL4Zaluhh27fHaPPkEraMX2GT6+ITYF6IYpRsDcjIBjm+DP4fN1lgbe
IEczfGUkxbgKo6cRCS30uEXo5IVFrxyJ9GrWJ8oSNCQ2cb3eKl1zMqE/1l2uud9s
rSxpQy492W+/JmQ27lCy1A8pdKHtzRDjoypZrREZZ0M7B4HBIf5N5laGHx6Wgfn9
1UkiZ9X9hDJ8PQx9vol0VjSmL/Opa+kVnsg0k6E7rbdimjuvxKmKr0/gT/1Gqybm
UiXfLWOS2vrv145AzQZzywYVHowam7Yb3ZQp/sdTal3dPamrkjyFH4ibiaCQgheF
Qinnu5emowwODyVfqrVLcrCB4+jgM/3hbAIly4kgGewcMBUMf1djvuvrgBw8yjz+
UgkjGE9YEFbs2eXe99S1CL54tYgYZfAe1qdzAP6PguxlzRV20Pp9IUig8iAHodl6
VrpJICxf1ZiXogLQclIrmR59+RWPwjLTZPiKTprGj4tnpax1i8JAQs2Eckt15K1Q
0Uk//4n2TASx+xpYVevmfKgPjlqz+cS0/FYJRjLjNqaIHu4zPbYhAsL4vJgzTjTO
K2pbwUXvpPFwL4/EgAJ/DoaRvaj3VmPqfLjlCs1/bJqpEOqJt4G+57cjUbi5Maq/
KxK6VXyxryriveuZ1efINe3JbYqL08bUXAMZzP5UMY/bI4IkgHOqulICRp0XAP+r
QLuVVetC64417+U/8KdoIUBLMXb2OkXT2JglOOKxCefSyAN6btwnXUojJJk3lXE2
nXdbjHkdfi8K0aLKhTThsgDhA1CQhBcPKmd/l1rHVFbCfwCe54JVizX3Y3w1rMNk
zPcVza53WJ1htas0oTogJezy8t/meA3eLKwWFYL7CS9RTMG0DA6iaAIVuQxrRIFD
w+o3iHzzBa454s+mchpo2L/1wBiL0cVV7th/yq2dOpt0DhPkewrib+nh9GlBFiw5
YGJI52o+b5eRZWfLBFiv8LE/vOCd7YHEcHxuaiMx1u5KDnAWdEb1S6Qz04m7Nham
nOrqE/kt0W+qxR8ekhDLbPcXTTJYbk04lnda3qg1yp89uWAOFczd0cExEacC3tgH
o058eKwEeh5QvwzU/Lw1KFeduYjStT0LGHSwgVQn/Ycd8ifTc1RgaDb1aLku9Bnj
H/RLp6ZQMgoSnyqSwZWzWyZx6xJQGCn5qrBIzkZla1TuL8+83z+2vcPYFQosERWX
/S+BgepWucxP5rBj/wimNZXhafjPkldJWRyatTjr0jeo0s5pMDvE9QavmvZkElUo
+Ocof7i1LBMp4kjkbw0tOUBRvlKF5qwLzVHf1uLbynTG3J+x2rJtAEqE0EoRERPA
gGXkAnwGsovZPxlu2bVLVlcmclIKUnuD8Yhq3oh6obUnfH0CAte8pIWlkpzQ6ICL
plYnZRWLg+v1X4YolDsXFS33BhEUxN//ti3D8MeoucqXrQaWotd07muYI8swo8j7
QKiR7WGilw8Ys2RfJ4xbUzdpv5mIAzTVo4DjIT6l722pmP8ln6FL6sh+TacL3yro
JkGOYTIke6AvJoBxYpRaSBjAp7AQLcBQ/7PXoLn6gL4zF6xGVICtYo8NCZnV9rBY
bThp/etbENMVfgH/OMQBQCUvJCRYndm7UlfDKPJF+pOu9oJT707svqN+ecgLOz2k
q2tFDFrouCCAx8XDhtW0KRIZXA0k00nYvFgOjlNiRGpAaBaQDTA1jcv8/mpcMbQw
q+x9gFKkJLtQaVLZjAOkEdU2otx9Unv2pA1lEXunQ+eklXYWtQMio1deAeNrLzsX
FREKMd3YtbvjuOkhD/fVX4F5uwX9+LnBvwKiGxd6Nnah8HPQfClJRz+rEnFwKyB/
B90vXn7e+EVWI4cvtYw/ELTolBfJkzR76k2vLIlKx8wsD4BvbBHyBv84gIlPE47Z
SQr2RUwCMTJ7isqP6D4NIOMEqst2Dc/8u0jSV/lIQVYKSDgpeg9VK3Hv9BaNupEv
yfOzv/Du4jAuXlzPRzSmhV1aJlSsVHjCy7LuI9BbWfZYTb/6j2pBLHfMeK5NRW/H
JE/BSwK/2kY16K3qV5wtcqDIhOAFa3TWjYzD09XBQxGmusNulPeOGYegFfHMlhZ0
WTbIGQBfF65vhhhmsVzNcn3dohgfKu4PnUnKdqo3Z8fWTJYj2yMSW7W+GXLmRcTJ
WtGmQkHOZVP6RUbtGgYoPBSgiznxCdKYB+eTpcrsHNLarfigWPqiyL8ghxHVxgY7
8DqkNqSvEqEFiM83Mrv29wg0IDvI2NqjFxjWLTb5xGUBXHM9SWKe2LgEqdowG5WO
VZeNbxkuNoyycgTSWHVVU2Daga27C26dOwaiQx8QeWMaYtWFFuIgoSpMQT3W5GPU
V2J+vLHxzM9ojFeP+t2/FSRMtwGAlWbak8R1gmJkBwr4fkiIdcP0DJhSKULPqYLm
mvsFScDQFqlUNsBvz9CSHPCCyRMAnQ1UnO8C67VTmCEUQBC+to4Ox9yEy5ckOJpx
Kxb76ImQ29WaMHOiJ/DAbLESSEuOdDMZcVFwRcfrgW5ktGcoizyHw9je1EdCDCHc
e/zM7tR06lKg6lma55ytfejg5/3ZEHRB1uh3frazjwTEcCFanx86td+/eTFxSt1x
H1Hf53+0d3hmFlUHVYngKjOho2VaJXiCVSJsaFySbMx0mx2hMiNaORkaYmh0Gr3N
DT7oxRB11Ylfp30B7kEKEXXcOjHpDr3SCFbpmtZH725pKSYZPqS8p+PPQ+oSfLAT
hKLfVq0Qs6LIIpl2OXVRT0zMV+F3qaRQP9tdv15VrLRXyJb0HlpvHpwfR1Kj+O23
LwwjoaipI8LfFNtmvTbd/1N8aFEwKSRFk6OAwMBjOnRpZADEAiDO+SlmCollULBi
lbeZGrfg+nMgmshcFe+ePIxS9DjCSxFbKtWSa0VvsHd/uaAsGnRmlhxTDZ+qfCIE
g8WHjb7CUt5KlGb14Zs4rhUXswznC60iokMJMRIAcRkKeHINnKeIg9veGlBTXCib
Ou2Q/fvCuG+eWvokufe2VjquUmpiDZJo24auC8v+leMB4wX0EmkeWZmilPXUKlEx
Bo/nYbcF0VRtb/+DRliIBTyxhj41Bf0fgG4CqYPj0fxtBLIoZrfvTB93OkxOZgs+
HvPuaqgItQu6wajwjnTS8U+EmaabK7SbnuEzLdcNcZ4BhSK4Dks6ZAv6cWimqalf
lngy52a0k0MUyCTJd0mnzikraw3k0PP+Ol+rX16IsfpJB7m4jp01A9YyjIuTYwUX
f5PrK+9E1XIEU8EcwM1R9ECrFUdvm2pCJ5fFVYkYxY1rt2JqYHXpUIy7dxe83IuD
g7pN99w1Dfi110gJicw4t2l1rf/7GOkPDVPUntv80FwebziutV33KgNhDICUHlgD
Ba99HNTsc3wC3uJNVanXAnrBbM1U+OJdTcZH12SIa9J7BGm52yKGt0DfXXN1HOvy
whSV7VlFUEcw0C7WTO1TUb2q8A53hKirBzlWo/MUBClXmwRWNgXlf2vAaPA9npBj
V1VZVFOC88vuTbxoa9Ng96TV39ZNTY99l7J5LbdcCytFKmwbu6cfY7z8BVqp1TRu
N2UtfsPEn+IRgIIxNEI6VWtaWcHSEYGS36fh2CFKjiNgSyM74owiS/Jdh0e839dz
yTTMrHsbRiUnwcIlV8/HOZZ6RqvGCj4X0gBy3N9fI5NHouUH8iODhG4Jxo3FNrqP
S2uCYfqivsU4cs41hYqFrNIS3Yc2iTtsVG/4gdTeSB9lwPRyaGCdssws4/Xaw1WH
Dbu9IO8KBPSW5msPsHP43dAI4wWI6NDDhQ1L7XSBoqq2biZSAuZjp2plAK8xgk88
GKLnLyo+2RhUB69Gwmth8YW+lE2nDsz5FibpUBPFDBJxfCikY6VQ8yLFALNUmjof
mdYKLm6tFcqJzZCgFVkton/FfImn5UUrQ5hJgmBFSretfss27yIxVZGcIl846qE7
2IuVqMlbbpWVZ1XJV49JwqEl3QR9q7Qp7ilS2495EGR5dIxWUjuVRzZ93iLQOyCt
p4dl+AG1VxR4ZJiYHkZjuXV4x/ZuC5rCAz3pV+7RIhA40o4eTqEr3f/Mw8MEHW61
/OI7XimNTp2u5yze4r64ZOVczSIg2DT04pPABdlH9FmDiDkFudvwCiRTXcWVz+Pt
tz/DE9BqTJsTgXzwCMbqIiq1UsKZMgX3mwWeo9kOGI/isUXg4oGnuFu3XhtmuORG
mZKT3fbvevacIh5IXuj3YL+lTrmsAj6Eo8JSE06vziYTk46ZarTQYDhWqplUs6Sp
V4waXCTzoJxeU36A9aHjGK12y4gd6dXKmN5ULB7goToqkRBjnuQeSYU7PIY2Ffw6
8AdzkO4YCZlEdPUKL2EokE4jyrJMiDlR67vZIVOC/11FIEOq3E6PFJsJ0OoBZ81U
N83C0gcZnogFqKe26phztorp8fB6Rf20wZNp+TcMr7Td23Vr+dU7KqaG3wpmDBe6
hQzoEd/E9yGO97QHxtGzwBJ0kSCu+ZdwdxbItzJbY2bK7RxW4tv6Rr/siUsZkGrB
UH21RMRo2CrRvjcpkRAE+fLqfaecuT0a0DKET2UpLcxrU5sRaxZhtIXbaFCcyUro
1BdQBL/962RGgR8bZwSWXkNxUd2jILCtlgPw60xBt77eh5/Z686UDFsghNlqQadt
6zNEi9KTk5Dm2mguVbaT9A+1FvYeWMV7GcrCRuvyc1twnHVplvbfdLZCcUUjQ5C9
40VFYpsn9o7+GUHS6tD1dpx0hIFspyCI7z+bwmFQYID2CGnCFluIvSKr+LUVZ1FD
mqaD4N6kr0b6BJfyEftnvHMqrJKaSV8eKISGVS7C93E8s4PG2kgrCiz/0lO9idCh
BrqIp+WYSfiZbBEQW50sn37Atw1sxt/v4OUJUtgBDkLfNtc1s0VJI2ynJlseTz3O
Hx/Gw86hEZPtJ1NjvwVZ0U1yZrYkO9ryo8ZM0qQEgEM984/k1EJ01bVJoyXXyrAA
2kZKR7WwbNf2D0NfGD2Q7izmnsCmg7u1TxqFVrK56oAQvbuOpxIYsupQmNK+9cK7
X6g8FEuoBVBZDIoHY/bSiQIkZ/0fplDO4IrF6slb69SowKH8uJcMMQytxrhvzXQ0
9Aps1TqVl9QBHMwCRT/0MtuYBoTLoUgH5IdB9fLkDvp2DSbJh3RJ6BVQG0eNndFZ
pnMA2L/pzY7Fq9Y5VsO5stnyXOLNO7Gh1qTZq08PhwlUKydsX336dOFk4/kwMxr5
HxQ76ndEFeLIj5eMJNu80iKSbUeOl2xm4JwmHu+Y5M0M6Qeu7mb83ItUf73CxZbB
8Ph05E3PajsRqctF3I8uCxcPpZC6cMFcER/AKGnGq7EmFykJbOGFRpqLWLp7FEDT
gi/sFy25rcKrIChVtejwsLFPDD48BVd01uXVIwezW6fuS7vc5K73+yFRusGjrG22
zMz+4SOhJxnaDKrajwDFrrcHDwwvHC2NjgaS0VtZ9P0NbTJPW+eUw7hUPUId8enO
TDrOgvqlPzz65JAV7qCE1pZvsGLk1UXVfyCfO8TOHjFRQYphzBgEZm3YrUGkzPuW
ZPFjIOF6Rg86tpSW072IqnoG7dNAHt8ytc4xrJZtKEhmSbrG7TN70fFtSGWmq8rH
2qnCL/1y7rkASK0KmnEMwdeqxVKvC3a03fY7fpK617Ava7Tivq8VyFW1jejgIFIm
AXqkvraQexoLs7+P7WDx2yd5bnDRZuqKQTIQog8u+w5aJPtwgvS0MqUA9MRPHmos
TGOI8ymxrTYgoQztnQkDIC9veSI2xcOaE9M1oR8Vh+PCwqvmruHmkxa02w2p5cBh
sKVLz4MSep+F6jxlzwhBZfHgwKztxYWIQMfZqK9A6aa3qTXPjJng5EZJRDUDSJGH
bviLJm9q+F1vK7aJPiGgnWFPKlZMJSvRX+iKN/yUm1+Sk65VEnZ9bKdw/CtNWFS2
5tEYmNyrn6UIsKfrmZDearQK3+K+/4jwvyL2uLVLVEJEMqwB2P/ayCx7tAcLRse5
vjkpZWqX25oK2RCojJ8NWVZGoGnuGK4HZO+/ghM55nQqz9Ot0E9FnmA6Nt+zVeT7
P2Bjcp+AuhJqFDaWFGJBTY9bUiF4FnM5/pe2ZfficDaS/uuhQ9em3Fe1Si+lhNPZ
j9AvygojKZq5kx028N4V5I85sTa8HfFzbJktDugFI4TkW9JAqelYOmXC0B3bOfTb
F8aRTGdow+yOEc0eUPIzhYlp07RLNx9eBma0MJ+xIEsBcPhgbEGbCOyVrj3BY+3T
a7kZUUB8bdrKqVHkVdic13SRWcgZbvPFr6WGveVZ2VhbMY6S6hPMM0VjnAEJQ83X
3XeyCO85k61wEmNidUPqqm0c3OkKzvh/DcixzqQTjvt0OgyeyaipqH/ItfaKV/4c
VuUpbPy3PX15WNXzQBVTIVLZ31SG2/5LwBasHAFZlf1UmxvcHN5EvqC9iSHnj2Jw
eBbknivjirVrUK0eMzidXfVfEnSWgHxwAVHQLSpKI8KTBE5q/tNBYAtqogr1HewH
F0diPxnvZLhbcRqGOqG7xsQO8LRG9aC8JZ5CkCMFf1fQQo7aM6o5/LjR+y71FH7b
NUe8e053hF1R18vT98z6fRtv/b7Nzx8bKRGYmez1+glt+3DKFc0+MoS/KgGsoeLQ
p8Fzav+g0jZnOvy1wDi7SVg7Yb3nKWUkJUENWbT39OaJSZ0olV1nwNhXjce6a/GD
df5NkL/cE5VTBHCZuX7nrytTe0idyz7KjbLl4QGKsCEGxLddMd8Tt255go3AYed0
D6aoPYUWOctKl2PrBtAcpwyDlaQBpuakTw3SeUwQr3aiEf0ETca3ptyavD5TybkR
3jiGpjzKraNyLh8JNyXtZkPTT/a3i92KX0cbKmdMhsBjBIi7mMZffWDEHDoGcyae
s0Nba3iTqyQTldZR1BiQjeyX/gVIWp8VbfoHCpxfpblSeSbJmSnfgUJSC+G5bLUt
vChBs+fuMOmEDvE1hsAMtqeMhfXCiwy2T+9Q/3KgMbmAy9xZu5/EoQF07lQWj/Ij
APbOGFiL3L3rqLKsJqe41VhwiAuxavO2a+f1Hd1108a+uegzAYPY8I/e8YcTta2A
Zf3cU9hLG1NJzbQn6T2HbospwwXUFIWHqIDTbSafJIJGefyqpdRWNb++bcShqw86
YNx0WMmk3TbuTW5qbTCDP+mKNPWD6L/UaDgruoUNOJ2zcgPJ7TIChLZfplg82+3A
3eRuMSbCiksEezc9rukkt5LtQS7XlXL18IXJTq0YSJuasNQOwcFDeJdzbpqLzf8U
i3DGPWVRYak5vuWSwsr16q9N7qzxQU4IF/9Or8DhvaQo6+ZQp/0U/6KvV7TTZ1ZY
p4Z0wLRFDefa7JrAfqeBfCIilV08fcSD3JANFMDZTtZmmtdaUz/vZqIv/KLnMOH7
wh5+CrZux+rUOkwsDmjzwE479nUtuYxlaTJ03uvo6QAovV8b7Z9ZoPw6wCFyDQug
AbVvakyHvNh3ECAeuKT8gxFjxaxqyxN11lU98DqFvsTqlQK8I2EOuM2vwU0hZxiY
h257MJzj8M0iFq2iVFvtORFNa6NOYucLH9/eC0aKpmSyHgWBwtfWXZO6dazmgbOW
FBS8Eee6lJTfndJktrM5YiussKi3jvKuRozIep9bf64zUzQKCCC0DwkTr5q1Llk8
/PHRtc9rmpxHmkkaFcm2AnfKqQE8up8NVZAIgen7lho1Wpm1QzufLjy9iDb14g0g
UJUFspnrOGx52ZTFevN6YC8Ele4QDPEdMUVwiaM1O4iyBmMOhA5uXLObF9YArgSZ
TqAG3GsYJYZuPanGxObjIVz/gMIIdSMnsBauh0UUDHriVwlNKRKDb2MrSZLc0K5D
FICNQJlsvcHHIhMDd8XfLhev8j554Nq1on0LTTzqwYkpX9M3o7pU7UDOGfGMTdEw
VR+29qnRp5q9yD3KoWuhS6f+d/LIV2n5D0Cl8eOySv+Fuxja+cAERCpzYPo4ZVrU
eFv10K8mNTxxXHl2IDlPDalcuFNfHVVsjpWvh9Zn5yKGgUmE9+hhlYKxo+5pK/zs
d0iCrqfpkT3OSJ3YXGCfuFinugx08P28e2en6O5pknryT+yf9+1uLax8v0JFmEgN
+Ly7kVbYD9m+KWleyz9q3pF91SJquVS+RqSeNkQ47if3HS2HOGe/kvVKx2jAunSq
Sfkvt6XsQDAhYZHsriXa05oCh/Jc4t54Wkr/gJnS2S4wSF8Mx0eE5d8ENPUWHy2O
X09dHbqHhfzvkXus6wQxRvchZDyd8+3J6HQiXQWCc1+DeOLKV/dYeTCT1Fpmaa46
hkAQcYc8ePQQlqgkBnIU5kaLKQ+7swSY8IPuZ8n9hOlUpboJzYhSDi9k3IKssxS5
txOtBh5tfRaV9iCFJlHKraFoRQjuAu1Nhwc4B8exTPoVzQrBqQ6AR/41Yw5RbnO1
LI/XPHezs6eaBd4E4uM3etQBxXLZywarTSKFVhy4YzUSg7ZB1qFfLpfRh/gtkMh9
GpMcJr85FD4+rNXzPH+Th8JO4eV2RgDQKjv8n3r/af+d2+IUYdE5f/DuRFO7gYL3
lLHsRSGlDhfoeDhwghDizb297lUdYAUNKgocCC6caKFUkfv8XUztN2afImSt4dEr
C9CfWWbbltv6Rl7irfFBgphmDW6GqSMuaB3+4irLUt5NnfA5C6oCFogo9KP0fEdy
2zFLexSFQdB0lWIsv20283w2MUpIifOwsaEsek94mUf7MVKUC6OyOilC4yE611G+
eJMd4WKS8EeAn9jXMaeRc2d/Yf/3a6pCblnP6i5w+7S1zLh6vQ5Rp5IAluEZtW4U
DjbsJZxX3rsY6wgrlKN1LGO1vyIKy58dGgdwuk6UFk0KZFuG0wbxnX7ObkBZeV1X
TNXeJKx8IHXEDJMGxE8EY1dJtaqIl+3NP3EKGzirNCDx30N4IF2cAVisrhWzpQcy
w2/Lwgc6N7qJ/cOzo+DxG/mVidWTdQkxAtQcjUcq7eccWT79ilLHgn1hJH3btRtt
/W6DzMxh7Kub9zYMCL2UojukYt6sxBzbu3b/9ZsnorAFGvUVxo1HQ9R0cK/FZfx4
xVnwcYXSOWxw3AuFL1+wh+EbuaQ5husxxwUqwm4cPqbcXbbht9OP+vjeHyT6qtZk
TAyy2dRBXtStWV585caaZ6kRM3nmar0+aT56nQA4Nf/WErYrpRIO1OpO3HMkR64X
mO+Ojdqp/VXNNaD7Cu80ry6TOJGnRJjTWxlNU/bcYMTCy0kH47+H5I+TAU/gbODg
yHFkI5qm+BNvPJwv2MT2u9G6p1V4DDsxU2EWIB9VQTVx7GhRMOfZkKlk9vdhnQdy
qnY3f+SEXpqgHU9QpkC0XovlL/ohFojTice7bfKnzFIc2aXM7urwmWahQY1R1Vgb
K6eTnWLUspRaZ3xSwOrb0Ycj3bEgFOiYrJlf6yIwZSHTNUN5u1Oo66urfWA2fEfQ
Lcqu/2MN9ndfDXNf/pMM6+uEAHrv2v1izeOIMSOWD/jHwjl67Ob3VHJsMD39sDR/
ddsBYdITbSfPMtbip9O0EUOpqrPomGgq8fU5G9coymFRMN/eUFTY5VZx5wwjbQeh
4zs7+kYZYm+kWazFANvhInAyi+IOOAPdU2OumK/YQDBC1pHotSaUyuszgkqJwRLG
/ib7lGX4GutSzBrqHR7l15RrRAwrbqdNlT0ww6lWr1DxXBIRkYA98HdoTo58tbW8
2AM2//U5PqJwP9BUoZ8L5Ks1Agxsyuwh/XJ2HoPg0Y2KqiwhJAPtOHl3qly8vK7D
H13UT539ancQmwn5GstkxqV0UrUHhuxvPTp8LYjuotAHHhwSLvUE7pyWpOc0GkHl
uvYiokNS2h2EnZDOKooWTDe+qEamHWQNdyCmvylO4FOMvRrg3XFfWZ/cF8mx2AKq
+Y3puiXdZECUpdY1vlfVFV30FpVitNByab8zSqTdhnmVCNDfrfn8kG0SFc0Jfef6
2pSm3zJEXYWcVrgsF+yO3Tk7X4AuCFtY3/r2ukoxoE4FTTr8oDOlEX9zU3tGY9/s
q3ijndUjUaHTC4m3Gubd6A/d5fFs4v6HBe4RkrDbCoT0guL5opZJcggNVm+ksxOQ
Ko0yNlNAQXdGMGCNYGICpcMRDI3DgOwXbNZp06SnEwWhjchdyubB1/kCrl8ZYtcO
kVFu2y3svimqveQEvaJmk0Z9nniyaPFNq0UUw2abpIoCCWgROjgigEBdqQu+lRcp
LEOThDaOx3Eq6aJmq8n9UGWavUklBsx25WmO6QBRSmo8rCgaa+PM7M1GDJkf/QaK
r2gxT4CI5TOHqRBN8B4pTBjMaXjlyM0gjKlOvWFOGXbrxPdVOuJ/v8z+mMjWWKyf
jMi3hE23J7dfmyPSDKZvtN0s8yLxSEJEu/vDsACWh4VjiAwPGmxo/gebNjtytO90
IL7TVnpz1/Cq5F+vR2FeF0aX5NsaG7uaa3xEJ+z1ndfTlVXQ0LuVexo3Vg57vFEE
KWczuth2GCUOA+eL2cO/OVTgE4nxYNJtc76D+yW6KpL8IevoL4lNd+9CXRsH0ACY
l82w5j4j0Uwu1uvi88g3/uLHlWjf+bWb1Vs66GI8wdlM34JAtHWENYWklmpyBfox
pL+6QvgdInY3xq6NpcEG5VaaacatTsUZSqgjzl4kqRcL+E5EVGITEb3cM1ZrihHQ
SJxngzD5Y3qaxm8+THRQIkpB7RODDc+hQO5Ua4ZK+a33j+UuI6UIK2KNnPn1WQFZ
TBh13o5zomNOKaG1mBNJv5BwY/rq3BVSSiwv64rrcNMaDAete2qcIVGBRSeSQX01
6g1KFkH4JiDsuKIfekKwPsjngOaNjhC3Oq9NwW05lizJdHfbhSVQaNezZw9zGez0
+hRYJSde4tUHrsWnexUNKVwxW6lCqu3LmcWwu6ahLfgbctKd8pvbEEMgDj2jcZM4
fN/hVQsJ40R3msQNT0w5wFklFPWJFH/selePzWKOujvkedwgCaP8k+ZZI0roe8HW
NyTzoqX6VzO5MSKR9+g2t5OsCUtBA8lLyXpGXqDoN5TYu8+4KTr0ew7NqSvDrLBc
tMfMZeV1YHm204iCsIrLD5lPJ3rCF5DERSjzev1QtdlyFZT/jzW6b2KaohB62MRF
+VDVcs7I3CsnpZeZVHkLuw1w1SskzpL9xfRTtomD1oOYnAUxB50GRiQqIzwOrFvx
arADoopDjgO5aSisxTAf9Dje4Nd7asbGC0+B4xxcWNMpHNPhC2PFjTrQA+OgUo/x
LTKCFF/F0v2dr7/fpmQkQzxnuk45jQ0DjZYPyq8Mix4/zQ3yvv+TlL6fWmBGX4N+
KYNCRR+6fqq/ZHailxZ6l56zhN2kHSj9pg5tGmRk7sN/brtrstgk+kJggVcWyI0r
46kYMQ61hfDS5KYB56ajd9lEIrcM4zz6GYwWzQ890aRdWdY3P35beXNIFrWDAPOk
/oR1BEB25LVLEhzdNv5opA9SZzm21Cq4GJfuiSCHWAwhABUWEEImPZtlImguR1uj
3Hi5pai80477CTQZDh5DnF9oUYNIl1qVh2CXGfKuFLnvg+Te9Y0Q6xlMK9AM1OMS
yDtd1wbN9tvx+2A0TnhHj2uV2YeDD2FohNcGRNkHBSzyBygSQdG7c7FOUd+yPPFQ
9jmhZRh+N3RG/ocAr0qBNNfXZ0amzXDj29fhccaBXztLA/skQyAq1i5vT5rGYUSM
ccvrPZ9sA8a2nCacbfe0OhXBNpl4L4hHVgCqrhkX+4CFinu9t2kunCVboxtilsCO
7CR/C9Q8S0gGWIEBQE8leFT9WP2C67XG2rvpMjtkB+nXlmsexi/PdKF8YopOfJ6X
EvAACDn/8cVNvYp3k5Gy6/RESTJj5S+WI7SAXu/G3pV2Mq7PNouGLpUjPx5g1JIy
qzBmKVrjRfLEekUY4ae8eAGK+pe4l6YW6vTOfwwpoCo9iuDKu1cZzHcA9fH5Xrxd
RdydfSpNEgQDKl9Xy6Zuw49i1FpIJu/nBfdiUUFjrILQoW3YmJ5yZmsPwy54+2S+
GAzAO7KTBbBD9FNKU/YZ1xSYkTzseHVX9yvAR5r7yQrUmkj/WyTZ3njcXm29HX+J
lsePaX9kNqSFIVAS5MGr3RyZnTrBP72EIrNOnVY203M+3wjakWww1R/9fDaBhHKs
G/dpMlgbkWEsslCfnedckfz0naH+yHPNwvaz8n2WPUxxM/wprI4fbUteFOrxdybd
KQt5ypWn+JMxynt66+QLDpDZFS6tDuifipFyV2C/7jCBFMgHOb+M3SK+fTGs9KGv
txDwHejd1etX0G4/ug7t8R+wjfL30CPrFRU+lCq77gQrbhtF3NZycj29t6kvFh1C
uzJXJUuvdq82SXB2IcQ2qxBH7i05hQS98rg7Q8bUrWhoMxtahL4jtQ7TsCH1UTNT
HfZruzx7PMN4PgU+WqIppCtjqaZhL5oLmApv7Edh8fSwN+e3ea4osTXeLwiBC/lB
SATcnVtBljy3dLmJUhNZwuq37Ol3lQIdEswz3CB7rLHpcte6xPf73ehd81xfWOlv
IuP8i8Qx/kCIRgdff5MjoniYsKR9F01JwXx2mm/y/+FUyREygusp7tkS7aw47i2H
LMOlOBwzsZfoiG/fsnLzOIhDrHUbb+uWJINqhtdvuTs/puRmyeWIzmD0g6DC8AvV
jONnfA0M5NcJ3ox6Xgh/uTPWzlFmXxmbETLB2O8HevNqfbqccKaOLCBKNuuTiEOd
wV3urGHWALS7c5WqhU41L664xhgZ+4tFExeTe897mQQ745XdPpFhaU5o9CEVFHhH
8AQQOC4uapjamByd1o/3DkfW2OICyHHDyrxLgADsZN93rZNnuUhNeYnR0NuU2/qM
lvUrtAr10VRkT8fhS7qtLCyrITEpi1pOx94Vnoz5WUwfFGTHdjiKeD2+Bd/H+V2V
4eQF3ZKWizUDcnO70jwySdTqx5V2/lI6QAKDITpCwxY/NnktNlaM3foV8bWSJFZD
6YRAak9ph7l1+Iy9BK4kPLulIxU7umiO8LjvAnoi8wS8k7m88TnHRkwtIF8sUVtV
fJHLMSTEyqo4G2tevBulruM4K/vA5yDfSVr6cgEIbTRwESjnyA4/fOkvxxGyQZHD
q3ntc4X0KS7uCE8xlEFQZLx4eI7s4sw8Ed82Ci8IA3ptgD6c3p6pt9D328OEtf8z
CDr4SAhm7/Xuo05YjnynmIB/kOSrYpUkLjmPqXVCMmfpk7wpgvbEXMwI1Ey/qJI4
2zrn0cs5ruPTMB9RQADrkh9EQcO1GlgjWC5sDeiTidFhVQqzsNnkqAOxF+lAl73B
9eGTzOaeu4WO0Hre5jHe3RaMKD5E1A7kYPgBSgXuw7GrnYowkFv2bZ7F0Z5roaic
pJd6FGzvKNHB4qPC5qeXLDoZeg8Cx071yW0c6OwntpvcX0t1hs7wMNYKiUTvX2ip
+051Vc8nO7vnyVGzU8qRwzDmS680NpyHkVmt9nU5CleJ/nTlwu/qgES8YcGP4tgH
SOhwFxhVgvSd+f6C3l0qLNtreZnib5PLvd+9Q+tpo0i7tWGnEigKzEWjnLwfIJgf
xS0+o3QeC9Cjeqm+ShNzqr7+YgQvBQ0FzAh8YiBn5MQ2qnk+8np+fME1lCDwkKeu
umaKOM87CX77irLgEn1GXqwMe8scyA2PJooBQ69I7MWrOtsRGYvxU6lLsP7vuJv7
NLRnOJxK5icLkyWH9aGPEX8FOmhK+PLXxU8E4ZOUJ+8vm9DDuxi1xIrCkzIYrcaR
/wieMhLAzuHgK1aPgK/AhzHJm9V8oF8rk/h4BIU91uYUg5LCzbhQ5HWwiFuhpBkj
HiEsL0X/OAE8aj28h4KRgZQTTnJTNd/KXeP3wIieSXBP3ipfVm6tyujWuMG9jIaP
SQ2h13/F1mQCaiuOtKoaxcr4Ihn+epwSyWViHDKt95iXW6GCrWG+GOPrL6aUlvQs
0Te8xrfxbgf0Xh/reZREMN4OBIfrzfOM09G6wjqsZ4rCp0461G8I04Qdgf/SI8vH
vPV9UO2XsPfcWzD7rUVFuhomtcrudQFN7d4l5REkSypaVg+BL8p5Hk/tOOkKkM3q
rcKowvJEdluN/49ajtvZdoaeP3Pxvqt4SfITbeoOIcyMBcpozU8TRl2CSFMy0o5z
U8aKuryq1q4ejpY7zg8rRBlusGXtgnYN++UYB7WjudA8a1WrMgTiUg/qS8xoN4Kc
BhzO2JUO7Nk9YV+BbTNU8TzhJJUcAqzAzcn6EtHAuXRf4AhdJDajCF5AU/yz8eUp
dCXZ4ZJ224qcrdIzDIPA3hJGeyxPZQO9mwwUjWz9BR3XhLTRgXQODfTT/9mhMaUc
A8ETeYpoyEVGx8qw+s3Ph/ZdDZiflqKscrB5evTzGsl+JnESwu7FWcs0GgM5PJFN
qOV+X383V26MT+inOwPP3bF8yKe6ijadm4SIeNVatwFpwnVpNvjNu1pHq+9XAAP/
Fi7YAGCxmRUifpOhxbx049/DDYmD0AKj+Q4U7fM1aMW2ljTZrvpKW9aM3XmxgRI/
zAUnQqC+XkeYSfpKpQHZG3ZlU6jgni44wrSJXZ/gueOUjCWpljukrLSJsmWDSPso
3/s+FQ3I+SXy8HTiHpEfQkIoS5L9evCOKzdstqISqERbd+ReLSCgxjbFHJ3QCpnV
zZArD9CvtvbNSD7BfbLBRFjjAtS4tgG4v2PNCFKVhSzsSKiCGh8abPzQmJFrtaKn
+c8DulQ+ImUlFMw7tkghdP3qE7lr9OZdbyG7mCfctE88WOqlwB5i716LTvWLlE+S
zEA6cY6PnW+fXnGHJvggfzAohaQcT2tzPeoh9sp7WdlHCV9Nj7mFmpR4JNw8l7sR
r59zMfEjqxMeKwphpFPnhITFo3FQDo6cb5IS0MvhzEMCH+K6h06hwub+CnXmjicL
Mz1AuCIEk3OzS0SPCy27oC5WyHZ5Cdn4vxpbEuHhu0NxPjKzbOnRDsxu0cuhq1U+
LIasIuu0JWbHq0ZYyyJQqzampYbIqqiS9Sty/YfklM7/KDHhVU4In/CYz6sBXmQw
5nJKm8gH6I9DS6hgtrouyLaVTqlwoV1NpSt75y4UwaP0O3vXz6rgAtIwitkdQb6I
Ksj+vn/Ac9FN8d7j/mYy6Mz5LkHcvKpTlwpY484h6rrG4W4PQERK6Mf1jVJW2RJ/
2qBENT+sUBeoui77PBV0IWKL17G3ebNKLSavi/rJoFfBNwO+oKZ6x7PhmE+lGkfu
LTvdw306Ttpj6zilBICbeUBBJqB0PobCCCX41DyKiUA0nzx0nDzXn9cu7HhKb6ig
oodupx7XRagf5jDKRUG6vuWbpSv+n0IroWJiEVtyQ4fQU47ZKehAxyBylT9SRQNP
6gzD2yVtvxKXOsZ7OWnFp7YmUv0OMcLSvICsGZfcYZ+JQ9igPcCjU/3qqbYrrPhK
CQaEPZMNUicXkttteFMa6O9ukpli7ZH2GGYTX3OOu8uLrHsTAfV+9c22RauQ6yJ9
caJ0Qx3A3jwy8ACVwwBgVvpZlUWQrPGlVCRecunaLrT0Vgmb4oFY9kbKAf0sHdrG
7txOlZjd1IpJLklo1aR4Hmqh4nCp/aQsKEjs28Gq0kxj7zH7C2sx77iuZllgcwRk
iCv+snwf3gvQ0SkNfeDTlffuVlfLWie+41M8Oh2dfkIzB+C85KXV0KGmFgluMkd8
j1dg+JSbe9DrRVEYjKHR0yQ9GUQOuLx7UvwE0AjQWqtiWvtMrXDMriwmYwWTM75o
qYBg1x6B6wBQCvJHDBV1OBfLjesT+7TW79CYDPykclsnRfpAfrWNnY9qGo4ycWHS
21Rx3EXa9PAAm3xKDoqrcZBXDiosbBbHFrSl7Y6A01GGSTmgH8GUX6picIuaCN62
2Wbe4sFHb4UOsXCD3zCU0btRvaOzNh9m6PsFxwtpAnneL6hxGkSQqhoV2AdsJz4o
S5KyAoPp8sdNs1tg352XQcqH6KBPtzASS5Fhgfbw6c7FMfdOYMF0eQmDMjtbTRU6
AaDh7qPDeYjcFGv0JHesoJfuY6A0UOIbwctvn1jtYngV87Nm4mKjo7NPyqwGDb2Y
AREnzoo+teFn7PfCwZKBrMYMPZBeF3r45Gb2zv86TqXi1AxRD+ht5gumpsp00F7L
GhgdYEy8CAgSopPm0amT8fX4R84Dg2xXcDK4FmCncZZ5u4udeKD2sb0mL95kBxvu
nfA9KSIAVGd+Ho2Y/YKllTcreExUUunxiVi8zdlEhDgDY+v3zbTDX0KW7aWDgmsE
mjpfLzTASGN21m92rAS1sqbzHwDVkWZkgWLCO6CKiToPRMMji65cib4DUwMw35rU
VuLupfenSN39to869eoyPvUNVpEXCmk2LUmzV+5aabkkoJxTslEj4kvz68rHJdFm
gy5F0Zzpya1B3SZ2i63vQQp7rkrCXtdY9O9jHHYiX4SpiACXtnl5DMfceMgQxEGz
8ZxQXVmfM/VTa7oDs7GyHPhJUn/3kmz1LXSBG4Dxay3BFty3vDszfaLueuFcqAsH
k9t3UHOXGjmg85ymTek823NakRzOLMRZckMCaq7egzryISLpAKUyxgb42zPowByE
F3RgpGo8ZLvdWgmaeyQbFSu70r7jtzsWS3zaQHywXnUTsA9wVePiV/y3nXaoMvUg
yb33QagGFZQYfGYC9V1n9UCgxhl8AMxcS2A1AsUKbzhHGitpUbsjoLeWjKWdaZlf
14yhy6UUYkwkgE521VzlfaDE3bi7wyZ+ru5aKN0rBuqO+2Ldi1vlVuugOwls3E5h
gfdf9T1bqqF+H3YqU0CjYVu+1Sv4FkR0w63tIekvdeYXJQOWcd8C0UTeePWr5Phv
tTeVA50rRAFE7FNS+FCY2c7KFeMSNnbUNbrVdFPRWz/IbslcXxKC5q9Vy1jCNZqW
YMH9wTwm5L8m2kC8WmIxlknB4brcWTH2iSBtVkf5drNNTxAtNn4awjWn79OC9GqX
axOY/48WDgOxkd7DlHEaweAeq6GF7/igdcMNEidVHDlhES8qGkDxVoff9SkvHht6
wYlc6uSvYx3vdjitZxTIFp+QIWD9EiipfftuJ2LPtoIqJ/BUaVcFxcBmPMda0o8j
RJt4MHV3N8N48BnKgPltp9po6vUaX8f/DGWONg29LFLSRriWNHD3qGMbvgDq3wgA
GKEBgfdNi2e5efJo/n41q/lZBKRrNOe9yCZqH7LmYESL7ecNI+Fpctv5sREa4PLr
XW9xoEeHTMJ6VuUM9yny3gBj7Zbo4H2GBBOZ63OOxCYaCV+TCCDqN9McuRcO8OOp
Wt0cenC+hdmXv2GDQHHpLeP6ZKQ82aZke1PpyMHcMnKDe8tFAzQGcbKdvdmZbCkF
USbN+xCC04c5M0TO4UmWjrz6QGqk1k75V4J7XuGlixgm96k7TBoVQDabZOCiz6GM
8djykV7X7MhnMqekuccQv3+ye/baFHjmxAwpyTdKMxPpBl/7sgY6Fl2Ji+TVSs5Z
5MNn8KcF+dPIHT+CleEpU314VxA1AL36j4PbQmhyS31jMjifZwuklBiDyDv909TI
79M5QMDVyf0rMix7CAP36LJtZLZSFtzJcYzG+GkGQ5lAXEwylPpkPWNlqP78P+ny
fIgDM17/4CM2NufFqhOY1MPZP5vUk77kkU8wD9wZhHNXcaIJL8cSqZUiEpibFiDK
xuAhDGHUiNuLlgL3uNqHlH3bn0ub3LJWL21919hFpJFbTJAU2vbVRxvWGYOSUdhK
jjx2CuqU9xrMcqSr/pAEuAD5yDfZeVf/1JmFAMvo51yaV2z0FvEywx/1wk+D8C1O
yBwTjxLBIreZK6s8Ydb0xBMvdtskFlUzK3GmWYQhOlePP0DDNjyF3vwqJXc2w3lK
UnjSljmzSp1vQasrNGmaVs1iRtrdqLy2Qe9/9yWWey4pyxOgYyatzH8HPcset1Xn
Gx9B87yFqO43niow62iSD2T6Hyo979d5zzWETURNCyKz71fQeDtBqAzUvQTR9fX2
ltfN/59e531PkvT7dj6MhAQ0wpRLV340JQmqp6I4263ZyYNDWP6s+J5XpYMk6YGS
j2r+DkJVZhvG93VlnwgxjRF2f0kZBidow+4BGoCK3gPotLFymrGEqKMz2VWJ7mvE
6s8bMwxgdJzqbhnQ4qYo8TbFRNEpz7ZUu9kp/ZnhWJAYl/UqMnOZD7zom8WLYVHK
1qV7wp19d8Agf/1eBLq/9Qf1ZVpE4niIoSGHeF1A1uCPLcRuy6OTuo8tmzkMUhRt
djod4rQ+cyLPwJ2Mb0t+0frqOzwaH8rFVTrZHGmIBfu/7BaWs5FmVchs0mM4TFrv
Rai/MLCxISi0Fak0LKzkTi0FWIVu+LPtPM0p8so+x86M7i0+GWCjMLFSvSM1h9eR
0v3lWwarCgDaSUICzL5ekg383YlWU5evTsrf9jEUkQ94m1PKLTOXca3xYzc+9Ted
dVhw2tuihVjAI9BjeiuRfzWTzn975CHrCSdSwxhPhzSDpTsBMeEr5VWiqeK+aixR
ZFgc4Qdt9wzHnQHDaGmdAVbhzDoUHv0wEKSdSLhh37COnkWpLenmRqBvR8nHYWCg
VdkjYFp4XCrv4MTYhof3yALy3B7tSdsq8B8heBKd9wbOJYD3G7AMhFdsDnYx+cf6
gGO4WtVLnLylXAZaY6ZJOH3jJ9L2uGNz87SITE7dL7AknveDTQFuGmQBI9GYL/Vz
gjJ6qOWCzN/QxQTf4wXH8CnifaIP1NxLyKUHqsovSeljMCWQApUO19BAwfyxxmKs
BWnACXc5TV4HW6Fwmkq9p6BcPtY0RHO87U/Ccd1she8OzqqmB5gcWG8aq/dvFE/+
GsbwoHj5xVNrAQ2ntnsgkaKJmBCAmbJE0LPGFkMSAn6FcfEvApCLur6GXn9+1oCI
Ho1D2KDkAv+362D+8UohOAzme0kiRKqP89XTV2/x5kjdNoQL/fvpbUkiA+ypcK5L
2wGl30ssGgNJ2expfe7h4fsPt2jeAcE0+TjD9H9IfjflJoR+T0TVXZEBW9A3J+Yu
tumE1qLcAWc1s2N7/Hd82OcuBG3leBctl93nk4iTA93Y8HdXF7+G2Ov+uWlxKvfP
aoukCpgPL/QPOIOmd3pAEGXMPbiVgVyH0UWGBcR5Va5pjvWwMwnr/a+/P4EWg1v1
eumpGQdsFc45gtdN9Ki9X0x2wRQ8KD0l10wAy9TkZKUvsKSvxXc2L91ae5MY2HF9
b86YYw/QomLkG1sDZoJexcjyw8fpEIRtgZpF6tm/pewqiQw6GvcTsVf5htFnh+cc
NoCYw7oEhB983u2rzWRYWwOjmepfLTJNOXQ5IN6kFQuOm8M/9lQxohajKxKxzXAa
dRqkBQCvMXEYMqRUil7bu01gQnu7lhK5e7IgHk27CKhHl3Z99FwY7Dekv9qRXa7J
EU6z7wSYEZEGXyvya9nkrFZKQbeYglmIVcb7UlWLmQC2/C+0gApk5bvcMJqv9Vcg
mGdZ7M9//9fYK2wDFCoIl0H7wuM8bWTuju/S62daJ/F/Vnx6jH68y/2TphtZhlGG
eDaQPr9QYS/OWcwDSyRAsiT8UzywDlVngmnE2FG4gGnMSnkGF3wkL3CNcFrX/k38
ebTAi1hqTqdsLIHMKePMmv5fdgiDk/ElPg2betXnWuTnV7GQrEFflrcsa91EWdnz
949I1/F4lRbc3gK8YHgMaiA4CnMAElmfCugjevd1Uvlp45GtAuTcH8jmZ7kfO2aW
LRJA8qODSxmOmF+T1UAaSXZ3c7NR/XFNRhyenpn1MZiImmAiMXDbUpP7AYuaPOGe
NBDOD+ne5wTajwoIyBoQIMc2Gjsibf8woOELKzv6ChsrZdT4uzoMjnkuJ/TGGyF8
eyavCJZynx9siGnJoTuiU0oEfUOlbjydWIyBV6WPzqdfS/Dl+M5e7CpOACNZXeSM
J0fvKtkEr31Psyye7FN8jXI/NRZoRyAbeAjSb1Y5N6K/lxmQSl5+/uPPzR14iAgH
rFoIGG5NO9Fdwz7HmTxA4AqOseDELFK4YCv0yifXiSTW/MRSDCZmPW5KsPjENFZq
+PW0XFULjxWUn7L4UaYvUXbfn0QF83A7OABKIWOVOqfzUL9hD5TBzBfr2colGoQq
jPujBjx4A2UVAYLbajvw7cRp1bj4BR6F3H7i9RzaMMp6YnJ+Vkc13aAPfYmBBtEO
83oOJJuwhrv6ph3ZzmlW/MmDKFkn8gM3WRpHPnh8rId5VY6NM8lSRc+TOezNRa4t
fx+2PCnMvXYKR2amCaCKH4D4q8SB7GfHd8JkQgESq7bBXx+ex3VosfzrZUMlC0tm
mkdC8UvrrtPMZZUqhlPV8Cm6NMXI6LMmmep/aILTByoFLPpikQgcWemoPQkkGu7N
BCWfYTO5poJdWU1FTWbPIuJIzsLrzlp/VIxLrmhDlbQsEvs7GrmSFtpmVso7jHpo
/yW9yhn1D5wUGcgmqIyaWeiJBTG5mUaAE/yO1IXm95zrO5o5IkrBgc9Dm0v/ylU6
dQCBSFuuUexRuCFNaUPU9wkAkT5bm8E63g/zrz40270NPyvxOTAbRjeU/vx7HMEl
RtpwOzZ735N4yG57NErCtOWMCzCaUVUuGrJnkPwGOzCA9miP233E/KqbJElNu4Nt
miqMQLTy6eEvJwbnfk9v+5QZBpMgIOOWXTdm1ubM3h9+kcMXqC8X5OOAVDN21Ki3
7K0J454mbRzjBlST/jMReXhoJrdXev1gVYAQfKrXrZ1nyjrIYddUZo0KXMdW+Xrg
DBzFA+Zba1K92WHN9dayKalmQ3aW5W0cX7Vim+bzluCZDSeHXF7sOm9hxScdhV/j
yvgpg6vFyhN9FPMp2iCtJeBLnN/pjl39ezPhdwR43mgjipws6ymFDfsnKSiSgmnU
bmMV/Hp7IUywUIj+sycE+idi8giFbokGSSuvxoHnlqHRkmRGCKN0aUemR7nEDsc4
9JdF2ZChb7cQNdCe9exbVpFJVh8kRcflwek4C8GnGyuySa2Vg+eCAgy/rJ8MRgRY
26lYla3rAXrTlxmuXE2gUvgShwN94AsNvpwyLu9U7wUYLDLBsTWtr4m1AOVBJqFP
giYe7UmL0quAqVNZ9Ew+Dj1XQqv9B0m4XYpzNh3UO+9K2uvTbTWXlYgLkcGMhDb/
mVqJYbn/V3LoTfCGGHwsDBlmxPnqvXAFQkXbem/ntCJxqeTUrRVPDoyTJLfnm/3E
VS2/EmjmdY31TrmtYj/697HnLVGpwK2F6qAIqSr14f4Tp5OVq59xzuCahECWRyMl
BAIvpdyl9U1gzcmwkKxULKLRYrtTOfXQuzmktvY22CoeSMXlZWa4MVIjLwm3+FYQ
EHSF4/rPya2gPjZCWHDLkfEG4qrAVZKwMBwC2PJ6t04pIq5KfKyRcsn1yw0mBicI
RjdHfzoh6vwu9lTPuEQk8a+yYLqN0mJWtqVw5rWBSrWNfZnzmy4/cnm94efmtE1f
/3Cj36G2femtd0nIq6Drw3SlO9SroyNZqURlFp203mmybDkXwhqUWwOXD9dYjAxu
RONPXA0gUzCjIXHEyk4genUFMgh1kAsXEQdXuMTe/LvNUEwmgYTeBnfjAaBzsWi6
xbeXdtGN65w8RVXHh/EZUbdNnIB3VKf0UGJUpSDsZJ6lDrwtPN+6FnJkaQvMEBPJ
2ACTx85n/S2Y4oUa/vrTVE/Vu1lAK2Mh2Wza1xqF7nfu7ljuxNvoyRWX9IqE13QU
1SWF1NbJFHFPd8FrDvH2FY6E6ItMqM96074nB3h32WsVo7A8tCPsGZa1+Zfe/FDj
3oPsqWM/Y5x5dRoS5WxkNV508ThbrOFK5Oz3+6YMNvAujRxWHyarikvLciNb2hfG
VOHS+O0b0neFZQbQxl89hAEk3VepXRT9zNFrqLWyoJh2GtxImIl4/LkO40SSEOxq
gCxiOnBkVLbLQsfiCkUT7H3gbcQIYjJCNa9kvrO6Iz1WsaN/lBuzwYomaQGpRZH8
5bcubvQVNBAO1p6pHewihCMB4tdTH6GrijfEOlxR9LPSCtj2d6CGgOe1zYqjkG+6
V22YKrL2BH0zTU2cfWeezrXGaDfL60CS5HWnU42ulEREI++hBlpKL4tcLA2UY9bN
bQBOsJkoI8H7NjpjQquKgeOTvlPhVsb4SN0psYNDaFi+TglmbGO6tYdn6ZYdULHz
nwWI5WqxcBx4C2OXsdgZ/2Hudv6OLMMVEn4fidFNV6bAsCpjX4BFOew/9emJJC+4
3AggfQ5dlmm0M3/+YWAYjz3nVn3ahhAXnzBr8v1L1I2+tE4QGf9yysGIMuA2S76q
+beoaES1m3ZlbYWdPUfFusZdu70wkNKe5uUQNUQr9INCW+7ODDymobuH9CumRQwq
IlcPjyfGRuw432TEpa9PcaW3ZwqQjDCK5UDnO/LpjDnZgOr/X1NMSBTVWXL77KMq
eYknEythbGYmz81q+KMxfsBOaMratQFdIPDCrXLty3tIcsiHAyyo8t0BwiFwnysa
FhdNFaPJlxpfIlMnpBLc5bSQIEh5jD/0W1NONdDcscL5NQLXC6Lwo3SwBj4jkt6+
BcmBEsY/5FsS2Axu8mVFaBsit8FYIYMgyow3j8c14+AOOOvDPK76gJNzmcz82vwy
VgxIQSBFZmJ5k5anW5KfTilu45gG48NjPSKgBB3VR7kcu3x7rv3LBzsKIaoCoRkJ
sbujF8oFS/TPEa3ipt1VNA1PBAL/xVq2AUXtcTcS1vqBcx8PaPSm/tDRLWauoV+P
IbqF5m5UY2VzXnTPhFNWh5EU4gx4q/Mmlv/BBgO7ItKY9VX7LPTKT8zVIj9HP9Dk
n9Mclc5lIewE7LZykm7r+UB/mIzL8bqw/8QGqGSXB6nehXHXXMY64l2voYk68qCf
XG3ocBm3zz4AkRuYKb9vbIizkPTW8LxBCaHSoPsTlioHWBRW50fFfMf1HMSz3UY5
uCaIk5TVRjXBttV2086naIA3cPN+hGr0YIQWyjXxAVnkJbokqubO4pNQ0JdS8jK1
8EjXxXy993MaEAV6drZJnTDotDz95dWwyZ7xlmtrRD1yiWG9S8r+KmqcZsONTqko
NpH60Wrdb9f1WKYlL9VvIj1SS76xtGQKtOlaEFNgU/DZ8hBeEX65dDB7aWosIsCz
BcMKLyeJoxp4jfEoE1Tkwe/JuA48uMvma4VhiP95iBzMnzAgvZmqb8ChgY6mt8pt
xbmIB8Y4HKEmKGb96k8yGS7nnxVUxCzYI6mARFhpuRbaXgVp/LBw/g0hzNPQAtht
ADqtwIN5D/APj/CYiPF9GraTlNzahuwRFD09DY2WtHr7KsYxogavDoceB6QDK8hD
kCclwYnbAoYkouYLBo59cfSC2LA/wIweCBH0bNzYJMZZJsaaZpdqP7GOM0EIYnHr
DWa4xM6x07RzfWB4oLpaNy2JQRK+nWue3dUlPnP59oD2lL0NBK13Z6OS+N3T68WJ
TQ6vRjK+WaL7D6xq2oa1faWqfOYcCpVtNfbxFeiDnF1CuC6m/wHwLk4yMTqIVns8
xCYFmKfZTUjfT4YojwT6PsOP+sHiNK4wMQcxHZVc7A30OyrWrlBN4gDgsV1r4ubx
P+LOOZyeChTyKlRx6WBJ+4UWp41YxjdbI8et1yNzffT/E2/+3wdUUVEBaiJcRt9d
7xaExl5RSXyHUV8Pwps83inkiBNgH67c/3++uRtHdb3vLlV3o/InZa8bS3EnCBKv
vbYntpq0FH56RFIvkGDpwsFPz6Ka2L4Wzoq5RaLIhsbmM0bWZy4mdOhfwgCWXErU
gY/8U/M4YhgD1x9BR6umHVVZSR1dA7hHKF8ylvdKWoNvNzFN72LrURB0k297Fjik
IH1DCRUBDVz7culCUuvg36U4uQN/1DH2xcDtrBqZMT3+NwzJoH378dcZ9HqvVRKN
BFMz7AVQp/rhPrHmUexxUgwQZ/VQzz+ahOlEEguP3J9fpDucdGmBHknqMlvMpvcT
1XKT/A8TKuU1aMcHVl/C8yGA6ipGiJUXO9+vgjD7TFK4HcQ+n/PYxUuqbJKcPryO
LN6xvl5gdrTFkEin96ey5sg+F3MtPx9ePJW9HDZh+7zuE89EXDmuquWG2wQm/ZDZ
BhkOpULebR5F3jw0035Aa46StNkSVJ+2xZITGtEmx6ftHbfW1YkmHjUdl8zwRLIv
CZTQPFbU5FatnM3d5KyeojJ+VTbUXMJJ3rx5vKbE3QUvvnKLCLtfxmeFuw5F4Dv9
hYb4lKBif4hiuLpoHTsbYSuYAktm9y9BVP/yGrN9XKDw9eXn7lxK3qwfXp3ruhwt
JSayBCAytBxLAY/G8Yf+5e1IcPQYQFUT1ntRJMuMEGSKLU2ttLxJXOzEREvSjxBp
1SkplPrzPtRynj64ujyoPWvRmmxW5TDguYUkHCkZPRVW21iDLbEF3B+E/X8UELq0
/J3NyxwhzZ0TbGMGDJg2CbjdZ56Z4Tuc68IKRFRWsWXt+2ersGMocEeJ0jxVzvIU
ONbpNm1E7tL4lS/Q34pnZVfPIFkXQ3bm0eUQdHuOdTb/5/an8dhHRjGLQXRSr7HH
cK26iR0X0Uc4yG7fsV8bCkjax4GW3soEtmpD2dC4SXkpP54s203whJC8cchVuZ1r
LbRpQh0jzG+NgwvBumpssr6qFHLS8Ig+5LWTCilS/Qz40Hp7tyDRPDGZ1vrjSWVM
yFgrGKQojZT9LuN4e/wlo4wQ8NfqX1aZEIltVOh6d2SL3sTb9wRrBeJ/ljdM412G
LWbzSLxHcy3cfEvR5thc5HZIJKuqWD9bC+lG0aSKYJV0nUxaEMRWo3s6wJ/S/S4f
ONG++geSdCbA1mdtrKnofJ3ge2LVJLHppydP20G9L9csQqOhGWd0NLxEMo5SE0QW
M0/Kq8Su8ptZiGqcO+wgowbW0asJI2nD2dMxPU8mSypa88wBw9hAwizJ+7JlvmHD
27ppw061cZIOyxeyYB7V73COyoD2gcZi/OpD6Ooog2hPycKZYF74HK/aMRQXdT+i
ZYp0pyKSpfXlKFyKF7ek5DuoV7/OfUhJHwUCvpGcle73X2bH7wHL9Pr5gbdl1mnH
Ss56xoWiKNyRoXAutEBymAH8qOIHeyTIDvyxKtwF2ulqihGRy5fEF3GBN7uEkp5y
k96BHIH31elDt+zkycq7pSJWpGXjQFRxOkrat/Cq0e2R5EcV1o5cp4A1H9azETJr
3HPqeIRGoPsHn0Y6D+WPGLpu6M2aQBcq4X00IjI2SdXhDdFBv11Eywf2qRpAIjoQ
+mkQekgJUgwiE7YvbLfq2gXFFQjIk/qI85qCVL5/wzoPIJmA2ZBlP57SWTRSjhni
csQvCnAaLo84PKAcBA8dF+gfR4Pven2EccRA3MUFhrwz7zxwzXqusqWFIt6I/4a6
8kfizPzW66ICOVhT9Qmd4AN9ZCNb2cFyJNBAaXp/hodVGVJhndaQancAj6rlf4Xu
9OLf8t3UZaQvYAZHR4CJpSn4aB4zDMebC6qUnMhHWnCmr6krgxn2dbaGwKku9nhe
pTIUWERW2+D+PlQY4LaEX027V6ILVxgeRcKxkeYUsSf3z9VG3Y+DDYTqGSbh2mIe
JS4X16L3t1uvwi1UpB53XkESSVhTIu0eKSgfEvAvSB396R9xbW4mTOIuq3jWWnWl
mqO1MLwNEFV14eA2gnh7ibfHaZzopaVAiXxsUziFNQf2nD/E2khm7stlqIUuTv9L
g/kcm664hWc3FG+HGNj9lnICrSu2lLAe6V1L3L9Vo0XvELsAti/gJO2ej1aR2MPA
kEDHnimZITGJulzVjFZV98ZezX2lUp6gvvfdkblgShMMUyY8jzBpBRzO6Kz3T5rL
XsJQHx1GM6YdFHhJQSTgQ+uh88x+BMS8YAjo3RXn0kiL/ZRtPiiYo/9LnPafSZbe
RWe79Bq7HG1bgVR/CUWXoM/PdyD714ZIZTBaMHqzU9FUyN2yS4bqx9AME5M7iwcK
cUA8m5aUl+0RYplSfyyIoGGxWcmAPBde4WTf0FlngfulvIjp0iNqiE1cBixVWIUO
OSgJilL6LX4AtcA7fa3nLvN5EaRuCzH+HR2mD8iJAHxwKFwyufC+tYdjgBsUPRvb
hE5remKvjE6Cj0odB5rk9ArmhsAOGJz/bdvoSHU3wKzuwraD4k9gxfg275gK3N5V
UVChcik58HEAuqH9OGBmtUWpi+CgPKmjFzPV7ywMBuZgxmVmF4s/XKTMSv2t1i61
pszWSoH8PSKD5Xugu+otxtpZGrOC1ZAgpA2HMrC2OVrXEflwrcgY6q6MLmTHzm6d
wnYPu1Ioc+JOAuUbyrAr6kdy0aerw7C4h1g0ltI1JWtMKgEYabMo1xbsRO227KSZ
cHkiPQ7Bg5vF4WFew6fTMFNYABFneeOVsg+HlVaIk7iYST39Mujpcz3AwrO15LXf
KUY6BB0hLLLQSEB4WzSHBrsUyVY1WKsMurfsekGSH2motHsl51OqEGzwekHOKS1w
DuI/RO9P3Z41FeeinZZ8Q3mN55Jakiyy1LH/OHatrt/wAgLFG8V+0C4xvt0s4e8I
r8A4tRvstLALpGBE3ix6f+SiRUZ2bxT2+qWbiPG5M6gyKvKrAyte5iizzcJJ7irk
Eb+zW2WTN6LLi+THdTPJJfQ1SRktKcfk5tLC/CvVmlP4B5OofhiwvAZba1aUZ+Jn
+s2U3VaZ4cMHvSCafJkOxWAh5nc53D9fOfPuqC5OtW67xBBLTJgGS8tiA6RW8+kn
qrK2Rj1C/tm+4qCyBeez3cn57oiJ8z7OfpOAK2MIE81H0yU/n4M6GvTt0MOcroYT
ju/o+Ti2M3Tt5zfnDQp1nLiQlGVzs2AxY+XcHvvvO4+xNOwVL1cEVc8o8R2augSs
35ZVNAmzYuJ6V3UYmdHBMDsovXHHmAsxhgEnXZx1en4YkFd78dOM+Yi8hgjujlks
4I3xlscURo10VPhJ7QHNlKDtomsHO3zC3ZqQ0qsOAEfHpDvDze0IQnnB0TyGSFlS
6MX21eDaxhq4kTNP40YRLsg5z+1K/T1c+ocZ4vEdp4AW3OUvwFA386Nojue93m4p
o/R5yRn1Cb2/5k7XJ4TMz3UBrn0BAqmd+hdY/0Zz5gPxAnofp58mJqow7StuoY9R
ie42XKqIDwZ773BucYlLmtcLNr1T6Ei84bGae0pNzl5J2+HnedMtcUpuEMnSi+Xg
FDC7wEfR1qnJWt9FlJ9J1wWzxdmuDBhMvstCzq8INxaoiN7qJmOZdsGh/dlwn2Ve
ekj0j3qBPk4WM8exDuxyRFZXvkFQtff/rtJwsxLBwTcMK20Aa0mPDW82/guNGGtR
60fKesREnJr3+qs8RWKnKlUaxJ8/7DfC15epMC56ldu5QXz4v9zQI1KW8nJZ5Bke
Hi18Q+5+SC85LHjMAnvUd/0kzLCs9w1X5WUVuMP49Cd+Cl/xGDUlMywNFigc8dXk
XyqmEK7Pm/hlkSKfnYQiXkH+VMSm18j18mv32oclBl9gp8kQmvhAEb/KBDjSuE9X
BfueNbD2XSXVb2pBL2mdS5ceVgaV4+26ciPKXDlYV6BJMhlDtNm0iP3FDYyx66+s
/7UtLyl/UEwday8Y5v91CyZv64SfqG4Yih0AcevZnxWQ7M0eldSpZkmgL/MYqCif
15ql3+b2THvoH+OjG37rr21w/l3/i76e+pQz6xwiYxUOO4CsYTv/dmD3bPd4sjf+
NlNP67gGNWyyY/JegpPSpGal1EjbCNHft1XpIeUfnPfBlC8PbFtXZt6qdyVtgFEn
TYJbLgL1h7d5TdfGCbtN1FhyyaPVm40/35KE9hHLKy51jBa5SGjo03nyvtXapAon
7aArcaaZegE8wP7UduSvOv7ukiXB/QgnKAYVFQ9QRGZ4Hz2GXulyXWB7m9OLf3MQ
7k4f8Y0Gm7hguuJ9fz6oE34AQ+aUF08hI1gIpztPOKUCT33zUD3LKceNyXDg7Tl/
tTV9SH+34RgvZSl0mJfhlztrlgjentEK/Pyko/q4oXTpYwjfDbNWS6JYz6hyn2Yf
BTwOjYnTHUwFqWOnbodXbwe3uZYBG1cyA5kFNT0aZwSdsmyOIlENO5ra9Tzbm8xB
YPL7UNEOZLnypa7y5MBs+1T1BekepQwq1Qg5hIJs4RTNM4aLiNG/jtftMBH4F6tC
BcgTC1W0pSiLhFvEORopCYhlFrknYLMub2G7ILqg0+vLH5ID/6xYj7MyZGBGuWfL
ZKl+zf2sgLO3vV7wX/t3iv3/1Jfcos3kUiW4/NvBuN2hEMj/Yn+UEgH/hWetElxc
xlmjlBD5LCHYdWS6OTbjPYqoUHTeloQffEJK+NZGuUNb9qGEIXL1liBlBIad75cb
zxXiQgbpX9ILC5oLrbPlePxQXlBUiFi/VPn4gJau8ODawY9r+kx2jROEJSVarBBs
GHCAz+zfjTrBVUeSceKiUOy6FrRv1dFIOGRJxCaht8bEaZ8k5jFsxd9D9F9px3Xh
fRT1UyTvbWUJQUymmUuvCX6oBj/OMuZoVvEsGFN5NFTryNLNFN9MDwsFtjWEJG98
9Wzw4TMituuWERQRPtNqiNpXEz1safdmpVhHCfCY525JLVw25I/WDr3DUi0h2wbE
QmHbMBZhZhqB40stpq8/PU3KTiUTBLpLd+dUDxw00sF9w+5jbnN5YCy7wHQ+OofW
Zuwsbrn0iopfkYDnAHvRw6+KApwZiDdbdoA9jmAWh/jzlzR7CE1MJIJlPfW7p5WA
ZIeLXEOf3nwmHKvcCHkrW3gqSR5gQj2VY9Fbm5lT2/dm2sX8fZTbVmOQ8+J/mory
PvcLBdQ8uvOhjeVnZlIwXcmcDPWIZRTsDKZQIBycMJZdQ/1i9i5xDAuy4Xg8wcJd
nPPmrmw46aPSAq+Gk+ZXQti4uojfQ/+MsPEf7JJVErFbBpuMnbqltalClXIsowof
cb6ek8Xxi8FfjKBM12GNfsf47RgZQEwBQIvMO5oWbpNXG91VkHprWhspsmGgcDWY
sHP34YaBr5+xbBs4kDp/CRXxT1hLj77YIHDpaSJ5IYvTDet0p8LjIK0Wrb1maZ8g
Uz20A5F452NrM78cIyVQW07kc5pkrvTFt4JePZXt7pyOma/af0GMfKXJLqxGTBUS
Aj6gX2hD+T6rYXuDAbFmeMvBphz/W1EmN09R7WlojbO5U4G97sD1vAT3wtrA9S2Q
CIiYJmyTQDIdLP16H04IST2fvDrQJEIMrF6x9snubgcSF1vrONPuPgBS8yYY1Z99
MvulM85r4XkhxN9WglOLs56zaFe/+fRxwSyA5Bl9eG7dZSsL5P9WQWpnG1kbXUBH
J19trVARQo4dzrLfzX/1YjdSYWk21sYsXcpda+UqwvRqVtnRTzA7HAyut7bGL6UR
OQ7K+PYbTFc+FxQRnD0VQ/fnr4To7BmBH6oMrn78VHbmY/0c5C94ERtYaxeHVM3+
O30DKtL2FsFntQNR6bnQrl3k+7NIbBV4jMS2tBQOF1eKUNEXtLf6OyRsezuQ3UTT
T82aAp63Esrj1LZNEC98XWepasXqN5HvQISIpgnSQ6c8LvAczznobgQi0QfAY73B
xNkw6V8yCYoIOIGM4Xru3261weMyFje6smInxAk4IV5pLWy3KL3MMsA7A+PeWzBa
F2yAHAEijfySkWsYEGyHeJTPPL5mdM/EFoLdX0QTIbfJPUcD52gXCYyqBDpd8/jT
uTestfVTQKpHcyLL2ReRfw2JdpFtpeWp9gxCqDuWCP/9QWLL6L8J0ATgzfDzOUNF
ZIz8f14U3qiWtpY+2lEMqwm3164BWCZCYdQFivx+Z8wEYEG15dbeJB5f5yo7oEX6
zARpRgtOdWvsX8rDyh0YtX9UvS3GbyPSI95t2sTGax0gxZdhJhdXHtxBaiQVyCPU
zfG4XqBLtaO6otniAHVuSSjpjS1L0ceooc+BchuX0SYjp1xdKdBjGwqsRrxFcgfZ
BlSw/dP96jwDDtqwfWjxxhp8UFu2tzIunNa3tYPXEGe+X/1RdJH9ErtYaTJcaxYe
gXT3iXWIWzUpAGaxo1wIp4tEXGSxcBE5oGEWJ0tMvuJd0Xk8FNCS4V6mmRznfCMk
0XEcCFRiqi5YwLvopkca8jkks3jd6+U6QZDSJKYmIUEBe139ui3iKvXrmSAQ4TGR
d4OFghqzqHwy2qAPpDWb1aqak9BupWcFSbrCwKGQs76n6fnVDexow+Z8lPsZgzrq
NyKGCFuXF5ZbX4aH50tvkHW+qGqrl1jBg0301419m7DYhLQc1e0UZgJLd01PHQBi
E9L4q7xVhKOXa2/DBSkmhtsOz/hvbyE+EiZHnlnEctFhnC1zrPhxUkngNQ1NNJ9a
mxj1WDJrHoxz5tpfcpaAn/R7Jlj/bEz+YL5THuj4vDtkGBAttZJMSRm4at4e4Iid
C8H2ugDoYSqeBxJgql1d4S3u4xey+42s0MJ5jBHPbq7nbeP80RFCELMWJKmi6WgU
Rl11voCCnSK75L2MyZpdwBs8bh7RLMwND8wSg5Jk6J9e1sV2G0eAxhndx7Dg8cYy
sbk5UMSGDPYrTZ2t2/+J3WhGUlXQnSky9K2OV08U/LRpLWULeyKSidTWIzJZthJv
nZX7CJBCIOcjNyY6TWHtUTo9zAZ9zKbtQ0IAFKwe6OjdV4YfkdEa335z0TPAZsVP
Z7GoDVkqsnmjcs5e8XvVBzk83npgSNJrzSkdTl4Zohpmf0hZye3FQZpkqp0SVqkw
1P6tjfLocqqB648XWXgcgb0JkiotFN7g9jmA2bP7+yoPOYwI92491v4BcgXuNBH6
mjlLUEi5xM4WOhnnxctUH4ZFSaZr8NSm5J1OhFIX+5wec/ntxgJM+UuBkaLeEOj6
sbTXDqIaFN2R723MpvdrPmb2gvyX5rQofIPQX3TAEexQ+4H8hB6EqCcUregEV4ms
G9ODe5dKPU55LI7In9keJ9LpZT/g0txa4hT0KA3utLFh2LcD0X82098PnaurPLxj
sAavgzt3KMQolbmAK/T+JksKsIgHeOUyR9L3tdgt9MWl97fJBZmfb4FN/NDXQkQR
dG+OJou/SNIai+VuL2UHzWuziKkh3kWhV1m4RMCnymXvLdI/rsKIwJ7Pr7JfGOLj
hoXnzd7kLoVMRM2C4jhcqT1YEz5FjFzX8U0nDIs2Lv3ykGC5YE5g260hr8ulnNjK
PzddIo3OJgQpK9skkjJEnpU4rzc3FTFCb54W7WRg+mw0UdKwbQnP8fAp3vWEAlYi
sv5FQ6hnqfeGWDo3v9/uNPPVjL/CUk7adgGUzDZAs0tLjhqHUEYl7lpBYNs6qtyX
P0W65Q3jOoaKaNcim0EICKbEhQyUM3bJP50FCAewTcwRrZHbU2NLzL2gySI0FyCv
hxygwSYvtcu1hoXRdh8pkwPf1T0wc7ANNSbEt6fihW9l+KvSBafNZSz1BJL532Lk
nfdk6F1aSx6bCr4JRMFK4MUqGW1rt7MDP4jHUCcQZIGjBCl23sFPl+poaMDgV23m
PRXO0jDg0GB1JV2ZO4hJ2Cne2YMIs7RnCvEdLUJBcsZ1b7dyCDrxXjgpuflE169L
9RSWuy/Lbz7lfXLfl5DmVMcfnnQpSZZHyurbpx4vznilYjDox7Sp07TRiL5IgAvZ
sF47DPXnz0PYmQJ3KrvCiyegFeMuX1+9/YiOwDbVyhhUI269VJMKooNPO/a4LcaE
diyGgmNjzv//EOIUwSsDkLjcj0DdG239I6LQOB0hhvY0jnszwOT8yqQSJTJuPWOW
EGR4YNuwVp56EnkbisKkSucSv2Ys1h/Gounsy2ub7K7z8hyVX5F2SbOAIkyaNpI2
4FJxKni7w1i72Ge3icvta+Pgs8xdziwvja+3B+5Mkc1sUPDap9BLNS8SmjKm8zQi
AHC8d0Z3Q1k0PEzGeTmNTDVh41Bcgz/WZq6TyScY348Pqi1BnK/p9LWjLPW4L7uk
5ORAUY/LXt77tfYFxNo5BTPd+9neqfolSnSs1MnFU8VH9orMR7YMcPajduWooDHr
xe+2S5SDpw09Tf45kHocrG4RWLoaR1NGMMyKJIwoTkcNDPU7ilHUV3eGtxHyNOCc
19e1skIlsyy1knMYqcjYSs2bV7Fvlp5b8y4s8OqZGndSfyviMG6Pd1fhr77ERikF
kwBq72OBh81y0yZlrzZKF7tmXAEVTX2uf6uC76MckFyUyO1+IYabEvQFJ6Yipa2j
yJEvh4jyF5SJoKZYW4tyPFQfhT/Zgj35JGMQpugZyFE47yDiEeEOgEfLRvyCMSel
pUxneSqLQC5soPQe9wgsPZqUAiJZI3Znzm+j00QRYzqy0rybU7J4oOvHqFlpzlyy
NfhJaiokROdqkmf3+CL+JUJNrHv7iqdhDXBHPRYpNjYF9MLy7iiQECSbeDYQ/K92
eolCTKyUdax0/Mf0Hk1ZFuuJW9gjPEfC8tg43VK/6x2FLycFbK7PHZMRkgU3HmtS
kgx3xPSO/ExRXPWhl96HPym86Xrr9S4VQgy4LWXgp8dSHjuIwy0KNI06YVcnGxfM
2YtdBUfZA/vxnAtDn4oBZgs+07IJB12gacT4cUYqrOEUFCrkX3Ib2nJRKGdnO3Cu
VMbjXsJykuZ8CmdwkAB7NA0qJujHmzBPqlm6XDl8VujAmhHoTxabxhLLU65nsGSe
kVx1SycUZFQDCj0tMki6jeI7+SadFr6Dv4rUjFIakgrjpvNRc3kDF66DzmlZiEUN
M2DM6sNgiPQUGY8svpzB5u20ur+R+9iMjJCBv+byoCXDLH4gJI+MoLcQUPYmqcGb
aG3P3jp3njXEVm+TnlM5PJ9t90J0UoMmD52Wa09Jc5h5UjpoLk68EW+zEk9ArnHE
lyJ7vRDK6EcfsEvLdtRxgYYOvfWdFWnD8CckQry8QyRHdjzE/ce7v8mudEDaOf5i
OcREaY9GoIx0OQdf290zh+1EAqTTndFTsSsCnG0DbvZSRdlY1sXjGPttMGwjrhb7
yPucZZqoPjtlAlzSQHFsLEc7yv+2zDVxPFMucEK0kpW8uW7ivz9GXZztOEaPO9OR
jqont1mR8QqH+0hOseBuW7P606gEGAB/SP2dDOmuU0HMpiQnI7cvlBrFokZiE9js
NPBHolSgBtjniw1B4QSIt508cnyozRnltigM28VBOZkafgIHQW3QJPV+9o1L5H53
1GTHAdkUioYSrXsfA0UJVy7u1uGh81B0aCLWKVJ+eCC6bweNoH/IODU5dJoWCQi0
LRJGgN3Bz4ZV9Yinc3SU0okZ0MkWyV8tTuB1F5CHUrBE18FHOgvltcgxKH0pSYsM
ZK9d2s2mvXfVugjrla7uk1Y7wWqT5uamHAgJOjpgDXjo6MoEM8GxFR2HoHPqUwrW
AyKlxLxyqg2DXx5TZ7m+1z+bWzabwJWgiZxRoacOkpIOZSByvYSEN13vhKOXiQ10
GmwtN/BkyTcvZ5R8/29TjG1BHpqvtKE64EqnNiUO+awhMEfYVqKb4ndKtRjJgJtm
KF1iXjYv2vmOhsddCSDPelMWJwq0oFcQrSRDA5mXIXL5l4fEPooSZDHFobVlJN2/
moylXSoNz4NY0zbheuATierDEn6nyznPL2o2jHMNfhoYsiiPSQpKtHTecAykdk6G
v+1zcXIVvtaXNeuWJaMcK2YAugIX+Eahz1qnJ3Upl3A4PDKqkLVG4ozwRnhKDV3G
QvKX6jl0JBsz33axq88OkWRjuy7hljhWsiErWU18m1reXUhfm3BlvfuLaK1R305N
qfV6c3ZH0AEldUl7PMXRfQvJ15/F2XBaDQfBW9Lj4A7JspGuoCkMBEi4tI3ddCWb
B6sECU2AbLXPpuCyo34HsQi+yaDqHSuos8IP9nz2bTfLnBrOh/Ee8kCA25bODbCq
ZfiU4zgJHsrJzh5+HeGAMTJ6Ua0uBQZpWxqgP7/13sm7w10so0TkvstZ8igKEz0p
akXrtd6gNtemuKSwSLG17vgypN19cMcA7IRbnVGAUmo/hr0yeuvcIBnFxsZq7OMe
3Njkoe+wdzK0qyXwXw7fTXePDdktVbOkOSabYHVkg1KDPgyUc+mDfWe12VB450dY
/XNEsRGxIBeyobYtACf5zKXeFrtLUb4UuHzt030gNkYFmZv5EPwvHdNldW1FGS42
w8JIyo9h3qGvRWBeUYfVeLfC6UIdMbmYWX5dOnX8Eqp2cigrvSdGILKcwIjwF7iG
K4usa3WlhgH42fg7FmzYgkadCJ6qtaKwkxoalXN2ERszktJUmNRpUbocrh/VTTqL
bSor551Y3C9xIgwC7IMjj6DepmqDpxIxCwqrHSYK8Oy96eLaSQrlYD+Hx9KGq/zg
BrmAAEXPGu0mf1kVNjHeIDBKbavPpcwZagoKJwnpoOGBBHIm7F83B8u/FwsVkeEX
BRJnW6GObDFoJl7+j4GsR7nK3298pcvTu5yeh8+5cfjD7F9mO7YwOXEji2vPQw3B
YOOHlGy6Hq5Rd0tbkn6ljE98ulFUJyJFNeYur4IbbbF+qTb4hjtXHnRf3+7696QK
02wLNi+MF6U043k8DsfPPnumFkY+YEv2Khy8zJUOOXUzKG9fbTQ1qEOADfBf5tB6
0OTaVAMTpv9++fhGaEZ6GVWPtdBMIXkDPWNUFpuSzMkit5CTp4Pwdd/jl+1uqpcz
MU+R3ZxYnkKDu25IdHxbhGa071Df2zkVtS4XgfYWisnoCTZmcUD0nPi8OraRWpN6
6zHwn6uuvmwtpukEFAnskOpKeXoN8yAV7caPhX/c1v8z6ljl+LktNaYEWXVUJDya
0kT/epBXryOR6HfMTpy8/x3UHN4AH2I+IkwNu+pEVwNJgWPo2e4mh6mFqLohmAxa
6kiyL9492kzhQSHg6u4sGO8y/4jzyX/EY47u5nWkVOGwnOV2EUaV7gbxEi88ojXn
QLAxkIcIlJkd4kjCEsCz5i0V4FvJX+FDdZIgGo7bQua52PaEji5Kf8kaasXf35ww
X8ivpWvmn8PQy4hb5Fzn1KEZ6rMki5w6ey0ckcpuGfgXLtEvjXu0UNADgbjFUcaS
abR6/H8Vaou/wgBVyn+GyV5L3vLSK9Ldl7v2EeN1Y940wTCkCJtBdt/VphN0nPD9
qlpJvMqfKun9glayuGpFzOaZKCB5J7Q/NbjsxM2RjNdYpYiBrwmMkHqkSeqdxuGS
Ed/HKkFnhWyQB/hhcCSqGMN0CToq6mE7xgsBsRjNsyNDQBZePcjRXjdJTvlaRuSx
zAgS13TDPjveHbVqe8WSL97TXaDrdqPs4nLHyFhYSDWl5slRVdbzWOIBfc8E6BpX
0tGY8U7NIDcyqaafGILN9+n/UIbISWnCs6RfnLVulmOOKoEPTjW3DvK+jqkRKAIV
LT9R7fnaI551ZPiyHYcad92JSFHxzrEitZD1kh72EMADDuXNV44kMm26xaGpvw4B
cSbqzePvZVCxxUfqKetrVx1ObusRU4KuJMMjouqlsGyc5GKeJiedfB3/VkvhatI1
1pacjP+TW0GLbOlNeYbHYkiufkoiEheW9jeUUi9e4TWR6YWz7Sz8hCAWEYo4ApmF
McC7SChs23TVJOlgYz0CgeyNusFf/O7NtXQWEBIkJd7thmDyGYOr/u+ky9wllNQP
FtDTVynPt5k72SncMJJvjmKfM4BrBNK0z8/ACok+x/UIEuaFzUO8bNzoWuFpLFe5
UbZDJ6jE86pUiAl8dcTtKICyw+thcepT8rpNuRc4z6YbAiUVxzYiBFDZN3ziQ0jN
z7poqll326l+P6eiByUy8QoaU4E0TMgWmwLuizYaHfiSxx7kdmFpgWUWBzVVdZV6
iGdxpBQxl4R9lIIBImYuGyFJVivIvOW3koKErZz+95aryxdtlOtk3rQO86WKnP0V
krXLah/5mwIQ02Fj7Uo3yRkAxsQcgzZleCmYXHrb6EmPPp7XvPSB57BkPUYtwHLk
pEQqQspxWU5MqS4UScixIb25QeGg1PAi6Eh5/PCUkjX3vW2tsZhUwntrY3MdXwmI
WdrM5KSn3vjjYjq8PLDLxWQcPafIDDqyws1FcAhoF74hzWSZMP/T5qGcQsve6eI9
wjA1RJXR9seDzaHGoFpt1y+29f0sEA4WcgdHcyNNfFQyM+A+IdbHwea6tNgnogl/
cpgTlBGPEwZdZhuTPyej0MLa76Hd42B0VZiDMxiMvJ8bfeBr+o79TDW4mgTKNhgb
KCyx0DeF1g4w4XjPIJzou6x6gO8mV2PC5J6YJrIETllKekApjCgTsYPazBV/FmwM
PPG0NZ3gL/ThSmIqlq5eeZ/yBpeJQ4PYd7z5yNikZ5GU+T3Ufvg8cr3rAc4klWZu
bNA1kLJOBP6KG4rRc012kFTFQoZXkRSZO7ncwnQIX1l98KBwgH6HxGObdHA49G26
WqwC6dGAhak0AjPJ4/p8PRFqGW6gvjdi1YXb6S5QDT8QgAYuRzfC0Kj49NvmYfBK
jguOsxKuriVUDwTlLCQ6Hq2xBbGFZsAz/Ce28+/T9eIz7/dZr1ZVa0SuNQ+hnCb3
qHdMXTOqJLuMhdF6AKmj9YDortC8oh3qwqrTn2bMHqDkdK/2kkP7Z7jIQugdRwRJ
4GZtgUjkS8jbSgyi2KUNT4s3NyQHgcksi+LHJQ/56NCzJ/15ux4b4DUKDhMCujbL
yCzyoBD/42eBANgr+lA6CuisHknjUPmCtceblFWh1qEDZrhn9TOg64NMqlNXLBvV
yVUZS+SZ2jTrmwagE9fin1P8OGtUE2IDst1os4vGKWY4J+27y09kPSJRX1XoVfXx
JDxICpQL/gxeKbokvpRERwXHINP0gIaZUzXj+XaD1ldaDVUaAGuKoy33IjPfCVVr
/Xjw8LiPFYyX6yOWIEW+tz7TTd0e7rHrN/fGZF7sPcVAI38MwKbB92BuJC9wgCnC
Baw35LJSFZ0v6SfptSdQoJRkq4ERCEuIbSBWNEITUpERNG8B4Qszign7h9YjtCxf
tPr9K6RBJEvFm6n/sEe83zA8GFrEzwkBRlhB48oGBKYAPUCX5KrgNyoh9/b4mOwT
AQtpyC4kLCTy5Bj6mKWv1aHQjrbWLarOWb1MGgVdjFoczyJ1CX1bctJAhVXpU2KX
jNAmeOfqb0A7ao6DCCFDUu5sPkIzoOCylUIFoS3oCsu1APHOLDo3KO9zaWZHSW5H
+2SZ2KGcNElAwQX3Wgcuvy75pInIGw+HPwewimmI0tIvx7w13Dc5qiT6/wNEfAWN
/LbzFk9lP8HgqkY6upzN/t1rZBzy7ijSxNcocfKzrEE5QTxidJtZPtCbHw+K8+S0
2pjAyU1JJdbsRdTQAJoepQbsNcRWodoW7i7mQ6iZjzKchPMHYd6WCKtR66GhnCZI
8Ci+PjMOwYJYs7+C8wGUr5nL5jgThVv8KigPf1mtb5QhNUlYNXa6O99wnIpLqAG7
+h9tFjmKdLQSexWvkRIbHyhL29R0r5vmDdvtuvSdmtizxBe/WbLkIndF5Nf/HzPq
42nIKISRvVqB1ijAkwZSsG5sqHP+am6iPDS5jw2P0r6U90yWOIDY7hrJ6wwuWgIb
Yg09xe1hgxhOoRXYfkyHAZg+gTT8APty9dGlVF0Hpa9dhxej0b+LwIUrHnQ8QL8q
uXpmamTE00tKT6nQpK0koE7alvaxaBVGSKU/B5oosgHy0mYSnYhT5AHCHv6GToTq
UuUapfUBx0A8IUiIhbCzdPHNs5IpcbV7Zf6Wt4upoItg/wFcYLn38b2osTUn80+5
+01QNIc/Dxgp4kHkMKwvmzeqBxZ2g76pJ9OufPOjrnmBfbIjl6s7SQ7hGzY2U9tP
mg+w5uQtdlBCEKujttRsTB4EV936e4XLRFTyLxzysNtiyVEjIncNlwO5CBHSSttZ
bdDN9PyzalCK6UwFVJm/9b4uTZHeZwl8y9cY5bSxYZ8IGlUvyfgu9arDKB46k4GV
PUjJ3YLldyqG1qGiTkH7UGD236hCtyfWW87wJz7lPMpOOryTDEfYnSiY4B1hK1oI
FTax/OLJ/JbgYh6f5u4GFRrz0d4lZQjN3+A7FCvQTcSz1/A5p+9vj32qFAix0r8/
XaYAJK0Qb2+0cxb/tbm4xBV58lAhh65JcVotxuZ2ZZ8uP9x8lr5DcxZpd0WTtUB4
jxVL6x3TyZzGb/C6iDdUoBr4UAGODeDYfkrjcTy7HYGxdQ/mUNcmWScacmgs9UFq
L1w1X68c4n9erKTnrMduY9GxvTgIFu3HYNURqEGoZhpNyw4DVKYbzgmt7z7Ka+9/
U7vO6ZVgEA80YRDE8hXIpFeHCouioKNe6kX7HrpTVKEtDvWkq6G+aayM1zWiqEaJ
Xf/tcMrrciA0c5PwmNegKBKBvzgmOWtQJcVu3A7KOrxIVBjj98v8L0HcHhfcqY5u
9BKtxue4MYZWM0aIXHHbyoX95pDQvB5gWhrxkvuYeV3kP3ksMR8RD8IaNwWnya+k
8W5se2WYVb2gvEamOA1xt1kJWF6gg8wkue6z1z8mMwVW7BNiPdkOWbot7MfAvfq6
PZcvmIgbF1WEl0A/dTNmDRxeMv1NZvg+G0SzqhQm9zWvSouKUJWJsgCdpn/ieW9P
VimCpZdjLiO1QECOZjHI3NG4HGOnGMjJg4gxWEqb7pih3duMy+3rJK3+PsqcMAe/
1oSHX5hnMX78RXK5YyUPIiC2zwugQW5Yptvn/iSwXxAyya1UaJEOPkfUtmERVYFG
cLCaOVnLVUSDB7+yCO2LLcm7GZ2WQVbdQMcJaEMtBtQido6GbRuvAvDWMB8sqvld
Cx2Sz2aZSpm5WoBGZLRXJj8GEwKm7araPvbaXrFuEhRWKfD4hTU4w36Ojlp0ZYxa
drmDNW0XLshkAHwBeX3iVUWuBXiO6nA7dVme+2wpH/FcoK/0V7Zf1ZpxkHhH9Coy
4dOhM/qK0YbAY+RfmkVw1bJFMoJcLvEE+d//vHQ69RZAp5d2iaY6xVRQWjHbNON/
GLEsB/A3kOerzJVPpzqB9jNUgpm5JGonjC3Im8GavtGIsYk+9ON8HYEiUGqpC2Fy
HBeJPfBe95fo/HQkkUtvjY9dhviswtNshBnWqIidYKk1Tsq1p6JuMuLQLlzVxzgz
nsObNUwjE1kOuADx3aL8MsNTLuNDZlskTUma37AAXlaobeaufE09XlbGKaSXT6eU
IMe7SWpnnxVRQNzbh6ogh31o7C4fNUZllYxYFOWv6Z6nBuPCS06/h9+0CyWxvixD
T0BU9YGLOHSi794XtzmZcKfn5A+s/zb4M2IOvBrWeSAikzmbWVgK7ujW3ugCoOQm
cdDKMl0j7qiGsLLvrwuzeparXixbgLMte2K/wxY8WW76cy2V2NlZiY114I6nwkSq
sQMN13UxL6f8huyWGArGwRSrzkUoy4kGC55iXGPFl6JtcyNSKeopa3eXT5fN4l8f
jGGXCc16y8pz/Zdub4oNxcuA2Umk4ugfO368WwZKkcrUjl8aJIapsOb/VyI1cqGu
HaSw2+W49qUWwto1vUeWPBh4AdLak61kz/ta32HKC+KUactoqbggpOlgvZ9qDwJ6
CGO8mPQmObgU7El4NsSR1/vAUS+kQUYwR+qsVjRwtXCjAhOrwc/5PlXEbV+X8vXu
4geqYVpo8abZNPfV/S2wDec0gVHIgAuScJQHZwMKNN2peEMRMACMJ/0a02Fng6cJ
UYan2isfxY44A+yWYgPyb7PFaAGyE2N2y2ddC0r+x3VmG0/6TiLIoRBWZT4oDlFW
sdoIS6YJPaMZMUmwbShH8X1g+r/oUSFS7TGp/giUwGGzejkJIeauAeQ9TB+pB3Sj
lN+sJ5SLLekGwSD+KASSs1yTAhvyGD3HwZScpJUPF+D3dbmVCsZVpKuUq812tLfy
6uAl49I4WUGWymvau2uDb6MlO8vKChWF3z55M5JqPTjj+qLW0amseZQ1iCu3Cqvt
eVAAFQnwEXbm1P2h9zt2XfaO/FlW3yaD37KzGMH63+GN8VjCOykgJqWjTTSCKsSO
sarcs5kQWa23wa1EjYwCteZ3Q/PPeYcOgbhQ+5bI+QFbb9SPbhu7JB7duCyHt/ha
RCwt4PIeUR1ku8jbdJnyfeztlBwZzAlBN0lSg27S8u5SIYm3t80LfuQ8Ys1mfJTw
42orodPbeAz1MBPC+LMfHCA6dE2NUXqUDNFpXPVtmmwIJ5n5foxUfwpmGVo4muEd
Fad9Q2sIqAXc2+5SCuh3fTxe3eeeruNn465oYw4RK+aTWfz1p/MfR6Bm7CMy/Hx/
9d0MQZKEpzu/cppWarU2QwVsKUQ+4OkYbWNqrnF5u3K4w21Vv2LWRio6LJ7zGlS5
JuvZbbPJwTV2tREMmdsKLoXrquht/nG1ut6CM02+W03e28qsxJujhoTZXM7Cxuq4
+uqJ4YSj5VjsRbxWpSFKLxhuBtohKOI43XNNKXfykmHMxRdeCbH4riqoohmHgq9r
cRXMwjJjNqFMHudrOaNjDAhZ+SI4w0cNjkwOVY2pE30wpFbyqGbTM9Qiv5DNwpT2
cu7ea/L94iEOZlufU9Kq+XM7x8QRtk/Clk0N604UoY2FLFuCGs5ZE2c9MWW4nF5H
RlULGXrQ40sKZ8f/R/WD2eJjkpWCGKKsSKWN5bTohuoqCM7VBfM6CM8AEwoJsfWz
mkyZv0TnqQimx35LRlAPPrKDOLSB2EaxtUlTp3mK2wQJyHbo0mab7n1SZB8+SCmz
f4EcilzV+c5+UlW8SlHRh/8FacBDK1h6XS/VkinlgTO20tc3FCWBz/jLJGMuEWmk
TZOGX+nbWN3h7TERkTOL0S3ks3AHb74Hg8Xm1XHWaEaUKLSWNrZbQa03N51nI5C0
u/IyHJr52r36vjIeMBCh2CYlYh/7rkbgj4ra1eHNH0R3H+HKQSJ4+Pu4YVdptqzG
3wm98zi1oFOFmoVa8oxCdmUQcBKbHUqOlCJz6/RfOQLa9JEETJJyxdOOBM//9Fiw
OENzwVyTIGiogD7FZiPzgaVxJbbkU8b9FctClTd35NpWP27Ml6sQ8FKVXIdvNjZh
VewEXVbHmAbA/KKRpi+ae/jCVlKf7yRjYqLEb2Kxt/HX8styiUg/NuiruL5wXObW
8A4P44XTBmUZtDDtjyVSpv/q+2n4mxzerClkFVcCeZ4YOYfDGKTkUnr7KAzAXiKd
JR6TsJCRTzeO/P2myPB7iC590ECnmaV4F7WiZJmJMDCNlBLriewp1gq8fHVSJEzq
1SArhjkxhsrKx+xHZ2XkY0VBqxkY4g+phjNz7uWsofMq8Lg63yI5Sb63niY05LBK
0OMVyNVmGPdFj2vPzh3bd0oVntvuvCVR87BOTgJgmuGLueJRDm0oCfMost/kkxBL
S+Wphcj9rNPvZd2AYwQXF/ry1OWkXLN0go3gPiX3sZ77UUmv7E6oIjTMba4rA+Hf
2m+o++mT/r5KzmAW+BQ5oU+bGeKyIjBa6yJUgJNDEmS2XDZdXqbQiDTARkSM/zSK
mG49J3y/JNlqTvF/Jn85MEKunkdUwbNCph5hAa+J07xbrkF59QNgkc/WcaGsYeaD
KB7cpXHXQ4dnTBYL6Lc6iZAEVB+JsYIV4JitSU39hd+aQJSG/DsG7HAdRtZGHzNH
7cm94odBSqKN8o3Q3cb+ED6WPORqfVMAkRVCbAmQ+FhF/qshz0HC2cDVcfC4q9+E
6lyeRUOiQ+Gut7FhrpgtdBVtmpVNeZTO9MvfBfbW7SwPQO5NxuF5yUf58WbD7IK9
4J9W5GRU/dfL9WhGtmfdhMxzv/NZw2KInVWhpUsHGtZEHvys3XLZXrq0Xtm55LVq
5ptB9x3KBP03ni8rTYrPitI3YFTR2Xjj8POSVie4FPBQUCUoz1YyiMLxt8MWQqkd
oF8A03vgbaPjciCbpnqCAduaYJUxq71TFqiIjWW/ogE/rU6W3nf/7AyRZH2dkhPL
26nbdX9tdFitshBfIDf4nB9doeDAcFd3H70LIEcAIx6J3xsG2inXGsx6kUFXZRsK
VjIpwWxH7aiF3wT/dTcClFlTl72cy8TYT10SPZKNSw5urJl4QuCxiSUSBindtFk1
lE/qtw065MUytd0nlwgeJKMzX8podssNew+BImDOGc6/KROHMcbNAXbyQUK+ocqI
6ekrkoYT+apf+lURknhL4c4tfTYlzyTxAcDQwWKt79T271Q9tiT15bcEnCFNkFQq
W3dzQFI9VzAcmL6dNJuF/DB1thS86w7SBLRO+gGQ/+4Z7lGTZSEvastz5hFpQta2
eS5EP+ZWlPqnUwJhE8QEhd/qDgoJ11dW+Fjl2OoY937DmWL4fQad5UEAPJvAPDJG
9aiI279TuqgyL2cXQxxtyFof2HVHe5WrTAXBzXCwSLAkgnLUH94LN/9Bo7TjtvVV
+/DOSGBT/rqC6bO4WddTYgLW0G/7tdeTyiy+5P/DQkFeBCQZgzkCOHMlOwdyV82L
TH8l2U4H+eu+dp5wpc+sFWDYgwhyvuoNo0ZcsfonEBaIIijzak4rTt2WzAwU1wMe
ORIfr7pi1u+2LuLhkTmeO00IsX8puOsu/2cVKn/BkIoc3eZd8b3Y9r0LMvoIWMdS
5beOh/KCyUt4uTjWDOKDVCaq1KGfEENkzn7QCoWJt0gdc4gTgIdHrc9YaFaMQezm
Bmzqlbf+8qWBeB/yXk1uiCFFY6XAE2KleheJk1n52FbEqpr+Hp6WTDONjfg8SPPi
XxiGlrKOXfMxD2IqYNgxDP+xu6cy/hRNWio7hLGe7D4qPAY7st9QXFLLsVaRaC+T
1oDA6lmUSrgAftTYPhXB/V1t943a9S5X+rBg42zhPSgga3OjAPPLg540T2+t4P52
Urz+vXql/Wi9vbTdpupjqvD6UQlKM0VtZ/xUmvffV5aNvlWK8g9yixTzn6Tkxf6t
6WvOYeDOO0Fc9NbvsXCNbjLn1sRrIwC3yyIkcr1n47tm2fCrVGKIt8L2y2D2/I9D
Flcq9dR1UDwxMymnGzkuMckYH2yQLQC/fx2ffvdokaWSULL9DP0R/ZM3jNYdiice
Qf/KSejwFHgORWD004O3c5ntS8PM6/7VYIM1sqyoDZ128iou87CWYQsgunzWx0fA
7wi0EBQf76+Je/RBvtd4HoITHPIjFF6gTANJPbemz4RsLNlgu4UFQkIrM7bhgu/w
hkJb/SRG4wB//gAHclpSzEE1sru+h/JYXaklBDOhqqDdYYSUOtom8NLCKKPC6ARC
SSCYbSPwhjmbgdIYIlqzStrEdD2EfLH1SuGn0At7UEiBJNBaPYmLIO+NgD5cZ/xb
LFePEkUhWFU6rfsnt2f9Hd+PfwK/tDHDBjZ2TvOR2peRFxgW6vR9OVAHxYbpPhX8
yYDAR5Oo/rIPK8/goBqGHt7Nm1sg8Nm0dNM3vIAHjC1RElOmubB5H/d4R2iZJJKR
IJYEP6iAwyICDdO42yZzoREIIBTu1tCFJKDscybDv1k5R3hrwrbQgpSknDjEE8Bt
xwPSxPHluZZ5IOnffyWYuolj+mlHbjJa0L//r8I0G3GkgAafFxuGmll65/daE1Lz
kG2BtOG3oNpJEAPjCUsYLmYP1TAlNAZvQC0N7ta2D85XN1BDWuNDT7Cf49qRZLfM
SybFGokOx2HX45Ox+PuhCMU/oHXdyQe4/O0a7sG2CpzGVlWD3mVwibCyyuY6ysJM
Ndva/G/yAOlA5nE0WAY4YTJmrYRuHRxOToM5QO8+2PVWDUWWvrI2RY0nNij71qL2
dA/my21GRmy0oIEiZhV3kxwUf5uu5LG/nAdJNd58b7dHSljqTrfQMuTOw5XTwuai
cg0l/Kq/Jtm/ZKUBwFTrR4raV7HA1bF9HsMkSGzvUruWAGLIJQxLQQFnY6Fu9qzm
00aXmvUpyoMba3M95rkqVdSxrIFV5wCnpd3fB2FJNPrYmaCNFkImwxPXLE/NVvkn
7ZO9iQTttZWnB22JaSPTMrC0qDlKo4C3f85jc/bVIRI4/NVvvqTWrA5tJaEHt20I
mxMpZp0vnXbiYfMNhsEwJy8w01VhgHMeV6wyvRhKm7WdQOyem0CEUjQ3GO036aEz
yCexd5fUIjhlloUP9EccjfOIbYJCxJ7mp16udR0TNxKe5XbUB1e64oMVfg16yfPM
MV+b4ksFD5lDlmgOxx8YJjl5FgXWFDhoQdw9AFFRQBVw3+1JfBlDDHY23Szi4kyW
mke0p8+w116zwnmA6UH5vTFz6fwHgg7eTZF/hV86AKKgNl1roIiUY+Q4hZZgyRyp
J7rdICYFEJ/24FNBuQay1ZF6ciFNXVYtKamhfjn3P1RCgfabZtNoHXhNrZ6+JOHw
4fqV0kFRVuKf/34KfmMsC9DAfhVpyWNh2c9ixkfZp26yON5MZ0R5jobY67QjI/6G
tkLWR2/uQIoRxIIA93iwxhr9rKPIKq40TnTaEtIy6noO8m8vUs4ny5GDxA09/M7O
ukQnve1Faq/lTLEzQz4gDz3Icr6fnYbqqc0jmHDpSt+EkYW7S8pys3SpAzbuUSGc
mNxUsE4V8ID7YkyMLqaBEbXQtEuEhVd/8midhSPqyx1t4AW07pr11vHCgYGHzerV
nicpsv+1wXOWlH1DNnRLMf8ektOb2iyFBgN220y/Qp4VoWfVDS2GT0YMyOKEshXV
F1lfy9EOFRBMpDqNcqx12ex+kC029eknclNJXjnDJUQUNx/5hNjNhvXEue8E8DT+
wj67ct+1Gq1yLez2OUahbkJlQCBPNjF3FPAVy0NrvnfBXv4t+ZoiCfJI9KgFC0jZ
QWsBl0KnI4SiDm69RNBbvDigl95Mpa+vRRPTk867Bs3whOzQNPleZD3HILSdrJzt
4O6P9vhG1r9Uxc6eX0mEu5Xci0qXv4BOr+dm9HEnCSA/Q+0dGfDaDzsOl1vBc16s
LIcBCMr0KMIZeFReA8ajxnLxZUDT3NXUtzcGlCbG46hbzYsz7rqEWRG5IgZNmwve
6NwS57nAQvmKIWNKAJx7dLpEXpKYDmPVzI02c3FgXeJKs8ReacxagWeuZqBjliRl
m0IsPYqMpNTEGyhafI6LlUWKS4RUwpm7wUtu0+PR/x1FHNHbCnNr3zYtI7rbIj1m
AC8DUUsxMNYwJt3Y4ceGXUHZlBS20iMkbDN9gPvGIwSEhhXr0vFcc8xRkyDHgpJt
TLmbwi3g7f2VTLaWNlRgfs1BT1TrfQBpgEBlpaYIJYsk8ONiKvdaJirnr4BwuvRR
uiVEenOGwFyswYyKCrFk9xd+VfUaKxNAQSbyqGLkAy7L2TCSv7pJ1rrTIDFrQJQV
4fsUw2x8zASFLJEf4urd6qetkmbJUpku3VqchfwHGk8sX31t45lz2ish88t+JeKi
H7rsM2b/y4NZ5wIJLp33zty34JK2slztSg04DDPibvHFz6zFKG311lePGZ0udfIh
xYxl0kVa+GGwgtKxgtFBztG4BBvaVUx0bemDd0UOuwpdJTGjoVGzYwJZTapgy06B
CdV8xbqqoH8mVM0WHNYZrT24Y60dzwmkVStfT6YX8dE+sulJDb1z2I3MVSO5ZfK7
o7nhlDYmwIY5Jya2OmGsDnJQbenGq3V98sHfjk/C44tKJUq88/oCGrEB9djyXeTN
+7HaHtOK0v8x0wEHGoMMwIoOvg8E9YRNpvMFasQP1fQ/q23inOd+6Q9OOU8yrZte
woU21WYK1qAf8gwgvZJL2LuvDsGv0WyKFCdmaqQRvsoNSzV5ajV9ruvG2MjhyE3J
hJmdb7D24LEzhTHh00Jn+vaNfjPYJPRWrAiB9kZRXUhKaDh0vo9/LlTVYVTljY/X
FLZ0anaVP8flsCQVDF1T/WSvotWx/GvSE5BmoPJTCCrt75MVZC+L5TAnSMSHCs7q
FoA4njGWaWsqhUd/6lKGZvYGw/9gO5Eb7J+me3Io9xpXDKti8ad/7QNWg+ILOT3a
CdUjsOKiZLEYm11fk4uV45FmXIrko0lWiIKWpVwsD54plF8GudKeid/HKdsMAkkN
V/qqX7esUErbwui5pnT5tLz5a6+Zqku/D+pfwQkrzcppmwlK0uIGJ5yIoPiLtSnI
unhmc9VvydMX3r4MPLTHPPAFmYKDduOpSQRLzkKsDuetGp3PfVx3KhtjMAV4nDy0
rjCxTOWRfk0+1zrLyiDcw8XmeP2U5nJj8TZhd5MzbIAO6JuB8cJVGHcWV8J74Xm4
wmvkLJjXNCUnKR8IhVxD0DwQXhe+nosJo0xxdDsQJ/J0dPHCWG9vNIeIdieLlFXo
Ylzksbdhmr3LP3XxFSClPvhFU1+GtLv06y9Cl521BRko7I5quGtqUrZOV/g/51Gc
HnmPoQKuFfZPcJsSP1V2l5Y4lJ/QoyDPXmbmtqX3SwsLI74WwCi73h247V+1l4Nf
KitYk5rZ2i4lD7gS7hsta/AnkYD4WvvwrTtN68lmgrbDjuTmcDua6JXcIv3mpa+s
xVNO5ulZi4S2Q0wEuSNnpaBZUhnmxhj1F4FsldYPAyiccU1n//dnJeTw8yz7EaWx
3S+3k4AblhgoZXfvBD+icq3hPiNwmVni/uZETFLWkXYiHfczBL3n3PI/vfkkLtzB
HPbJ1we0+3hLLh7hogy+JSE0Gc1mnqCa8+r6GOuwlRKeqPh2wSaG8+R0TCDhNcTN
ksPNHnmnvsXvgiZTqvbeQSO5+P4yLxzz7HkjmCVZq0HTaKZHKuSkEPyUHZbnaTE3
X1l9M25Jn3RhMYpmYLsz+DgSdF3/Zm4HYko6n95BD2sNE0wnH6SQ5cmZb3eOUpCQ
8HuVve9i9vqmmBE98ojF/DTaomxX+0bz42AgFBevss3DjIZU8QU6L47yAigMQNNK
MPWSxfhovFiZ/UuBCSdTD/WXl8v4RqAZ+AmGvCoBEXc8jgzZLP4vW7C9KQepZbjw
9OUjnEN/zYokn7BybmXnBXRagM0vkHWG/igeEknNNId4xN2uZSfT2E9ntf3luSSm
mZMyxYUoKeMspi9Xocz9z3nhbiQ6VJOKTv9mKNOcH1xLTLHhjpVlAcyL+soBZ3Xj
cd8m+RXdcUIzZm1AJpvA4lAt7qk9XGa2AfCztQ2grcdFzonF5jt/gfAOYnBo14cc
eNZlB4eiZJyyzc13xPEAwWUHv9RwT0HX3Y6WMiMUjhZ+qqw5nAMKYwt5tLFWPVQa
xy8QyloOi6Zx8RHnb7quBpMQNw0EJf58No9L5zzsIMdb7vgQ14LoPejL/4tGJJ/f
MxUHjQAVwXxGSM+mdIoh/4AT3gi6PhzLVsCsRNz7UNxAcBnEl1MeUnHUGerAn4eh
euEV/Mi1ni72SFdTFX3geSoXSNKRqq0cG3+gn+liyjgBFA25u8UEL6CKOfn3Fi2p
8jL9DcW1584gU0dyHvVTH+UNexOCm1XO00U4D9lK7eudq/+OAmgNyggKebdTt8am
bK0RL1lmTzGOUco4MK2z5SuXhmsSIbwsWLQfib51tIHLZElDh581+5zewGpvodcp
Fs6WBLMNUiBADteKjlvRfZt2ih0LrQYJ3yr3FLdAHYTMUhahf4HoTP6iEhQFyz2/
KxWFdlewk98FK/hq/NG+obwhA4yTmMG3NDAA5OWqgnTdbcQWlYf4JVc822Ax/XD5
Qji+VetxsoFvPjyhY44fA4vbj18MYgmdv57UhC/sXoJEvw7lYW8qF4DFp5jbPjZ+
Xe9rAsl77mbgclMKMY25YikNNuBrxMw17sT2lOSvLkpKCeaL3tMMpR0xtsGljcyZ
Y+L+Z1xS3WY6FZzS5jYg/hBp9tpdgpLrrQZLY/fkK5vI5Kepfebrye6uqvg3Gs+3
+ZKh64qZqOMyaHewNEr+Mk7mVBQhrCUWL2wWUmiALuh+yDP4YQfEjmIBVOWbzd9c
eDtcmRZWV8polHi9XNHJFcFD13B5hWw9JLrravYr+sdZ3x0R8lBjrV/n9hICAQE1
pAUAp7CVY5Lrzl27U1eLEkoGwTf8gdp+IA4zkATTu0Jq3T/S1kxIwIO3O1o9yrqm
GbCg6dTQXEHXM88mu9XrwejqqcDayi/sEqAuVGRYlXS5jB9xxsg5Lgh7Nf9mgsZu
s3rSaL4g2NJOfpL9D9b+SLyYRFk06Ifzf5vGOeFyW4w+/Gs8oNGW6gg4xVgW0doJ
ZQonxlVSIKPduanW7B/vjV2YhmwpphoXWpLoOmJ5F3/J9dHLHNQQ3rsbyDXTNfuP
p3cuDo14tSt/CUuNcp0KlmWsc5con1G08ZBv10rjXp/jMMSXpg5OiwM8WUjUxVSB
Kc3tEPnvCNRvfJQLXwNfENx2vNSktSgSM0zqQ4shph6RkVJ53DEVze8pSSvxc/Kd
W8jfcPDaPn3i0aMChiwUem1jJHsKXjlS0J0KuzQHL4rYYVd2epHlHl369uh81IhZ
6mxkPFx7U/u9QRfoEHwtytcUaEqy8E4512JhDTtic4Hr7RrdXv993dASXQXU0ZOI
EeMTjUJ7Ng0o+B0e5rxBuuNlIiDnnLjHvbQ7rNhk39rWsKcI/eKYt2crCQ2GBv5U
cOkds27jKKDbJXJCxXm1QA6iMLPw2oMDNkciBM4CugouJad0KD50B2wBZIvGdBOQ
s1mFA64HKeNOe5t7/c9ulNv7XK8Cj1IrNcmgbyPSw1ZWHUEwRXuRSfABUsHbHR6K
s2V1J3PWi+dt8yeGnB5T+ht+xKDIZtEDk7zMjkNd6nSXC+T6N1HwjkjQJTX4asUn
Wt+1SkGIVApS9F82PsPcu3FpZfHc/iII0Z6YVrgRWSmdOkuWs6dwfzPbyN+vHYuk
ornvAthQsKjha/0vLG27gS+eic409ylMbfBqP/YKiiI0clu+FfxaVsd9lCKmXTLJ
dOkLJxP6AyQYn0/VnPZJi08jtnL3EkI9b6Sur8vRRXW1vTMeQzPLCGVxWWZG0fDz
vLKDDV74DEZD6KAH9380wo3gOiJ2//twc8gGtJPaVWZtXmuUWs50MUFo1ivDlDv2
8ilYD83TU92sMPfbYQU2Xc4Zd/ibu2/a26HhSTK0vlUNt3mT2cvqyGHMib/jmDPH
X5wJtlzBFzG19VDWDWBFW6YG8+MsrayVp2yMLvkCZgqkrKokvKpud6OlxiXWhJsf
ccxjLYSDyl9tfiP5oYr96lhJWQQzh+jRiVdLanJ5SUC8wkhYREhmCEAt5+d8OTPW
n9Bj7KeMi519beEzNT5fgGjuSmytLecfmiv97tqNzx0fyHLlOE+4dxrqvaFYp8Ao
wZhrDQN9y2HT5iASZFnDJy9Jr6JHPV53wXMIw/yZpnGeFxd9P/lGNtV6hlrSj4Ht
TL22uhNFouhXhWNzW1nOLEqz28rIYrmgueKoHdX8YM7g4NY325FTkSb8HvypJ3Fn
015vWwSAr+5uFLzYCHw3Hcy3B0gAT7iUDoNJDC84PAoyN6xil4/R4BnBkPsQVPjG
jui/TXTZCvAb78rVSNY8+98Tc18841DRpT4hTYV132TJQOtwnUQQcA23T5OyHUJP
7YHc+2W5PXj+0CtoZygGqFhoElNc0EAftPoCJQyKZD/PukE3bCFYoQB69QNcCo+j
H1a4kZyczE1xnBSuz5EiK5U/FHRY/hhmDPdSc6uHgWAIlAnHBX07hRKdms44/bWz
aCzYdyLF1DN1hnJhSt6AJcco0UxNxR8YQ+Ii3zySRdLGl4q8UX2E4r8ybUMhE9LN
Do9RaiiRsGa4AbAYXcaYzXlNpXLDJ3XGMIBpAq8vQvWAdSjCuOHnI09+MWnZdBW6
gqBOG/u36hLmi4wzLBanQ2aKOIyD5uUYZ7bI3pFVJFMqeLrW3VAILkeNWVO0Opj6
64qCdwoB7OS4WY7LVVKySEcBEvnwOUf7BRJkufAyR6xvDuHygrPxi0cC0IkFWnq9
HjlCQiJTsDZytTWbtLClEFm5u3D7NMgCLBzVRd2QrlPre6VhN5HoSlflVykadvx7
gtL6Gv0vyo5urJ+5tTgl71VYdJlJhseRXIou/d8Pid6mnzi6iM97BTiM1NIkfeX/
EdYhCs93SVkBAN9wGwpaEynnziHJjZhAzDMqG2AaIMoyczSHmlj2SQqAAAUEE3iK
JTmtGy5tkKWH71xe9V27ISo51OWZDm0qL9BjstfbG76+8b+JNzXiq9kbYwWsVGcs
oMSdThOXwjx7L/bDXwNLpWjBj4HLUMbPG6A4SXkb9w5fy+lxlJBTyUvuXkW4JKg2
fJWZeZVXlahXF0NRQgTjkv/B1i3ZT8bLRovtHXXSzM4IUfguhjqtCg8Ov683OOic
Bw8s3lKEdTGymC1bAVVVwBv0rNnSGBKReEtIgWVhK9+RNd7lhJfhA/DPfqzOB/1p
iEJDh9ejPHK1RMY37Ypjz/+EfgCEVRs6uPAQU8DXlL6kBo17DHvOu8NKydE3InBX
/WKc8LPugdV2Cqq5oQ7etyhVSPi8n5cDKXHBr25PguPZy2hPxOpRDrgSENqVMunA
HO1CJXUDHz4gbRwgOCpP4juO+43aVePT3/P4Abe91sc8z+GRJW8xt3hv0ive33an
phQRSpfz0TJzr8xg9Nf44Qy9zs71k8wpS4NmZsBczK9Zb9sSiFMTyFNYXTsAg9gY
KwK7EOjutkI4rV0KP6zTSqm0vtWrP4h34mfIPUvEaMPSC3TfYG1SbGN1X9ZCMmP7
T9Q3YNUtdYs6NnH4yTYjZ9I83E6U5dgiHTaQyQ3qSkKaeUuzJWVq6dfhixKF4mNj
7OfTlHTcUbgWZA2p71Whnzqj7zzFKsevGMSB2JOo3nLpzcLbWt2mCRjqA2qP42EK
KSnvFQ0wqE/uTF62ARMLDYK8Tg7f3FVq8Rs5CQstm3zV//GQpD282tkwEqMUwySw
bUA03WvPVLFF/NubE1LixydzBiXKRXeHNcIWUQ5x7dOjDQqYDKCQlXoH7nttvNoU
vwVyQIfHEUjmiX5R66/vAdgKO6AxqLwduFW9iZKN/NJKVwi0Vy0LzSp5Xb/6Ndj5
dpzhLcGvYDFMi0e0Otrhm7oIqA/TebGdnUGpNO0dvqu1RWpIsOJEEUhQ/S9/bUVT
UXsB1LiR6Nr7mTqa5gEUuLJPbfPuBK6+kJn8ClSTA1qr0yZRuJx6fcUgXHOfGw5X
y45VxXNQQPB7Mjy+lkYPbAMG9gVfu7T32NBa04oxa45rT3Ojj2FPS3zOMtKknfp5
EGDeS0YfGP/ojXLxYY4jjmWQO7rQ1G2Z3JHv2U47TL7/OxHePA96q6XDJQKr+WlO
9DuBQLTPzmSnNYhbE7YGMXUekwJnKTKtuoJwLKuFbngs4lhYu9J+ur5rDrZBvkAo
P+JKUx4vOfUAroaWQXsQpI+Hr8s8T1OgY9Ri/iqTlKksTYa4gKO6fgCrzJlSvGSl
6PP/VkZ/N/hTYKRomc9Bv2EC22XExng+ZBovDGyTjB3aHpaxnnDHdBFJ8XURiDK3
PRYYIJBgKF9ffbOlYs1Vnalv0yDH4eSH+N/7FNFcqUcI0De3XuyXWsspriJ3i74p
8OWi0C+vNg6S3dLT4Zy8woKIuvP14nm7OWLmqnRRrKQS1LyFyCHWj1iivjr0XM3Q
Ruv1Pnpz42Bl2YCVpa8YuXkaXcDDK81h8i1pnVU/xyWC8zhghuW6kQwzO9QquwQu
HxDfTToFN4ZWQtGqcrAqvY+JksurYcjS17hQmyExO+h0n5b4Sbmsra0kfshpVkos
08H7ZCUZgJQZXB4zATztsA0qV6xqhpNDYFaIdWPPvZzW8HAol8pcCsKuy9DV1Ijd
hp8bqGa342QGqYtlHt5VZpNvr6tRDkwqNM3/qOJhizGLEgsaImhy2bdlKrAvBOMM
UtwSOKmrxh2eN9wwBJj9jxt/ZEvSaI5vgurWuhBstUyNQiEytUCIHqYaNan/GnI0
c7Skd/UY1HVyNOnNMuE7M4D5wdo/HSM02UA1jIAVirZ5QnvtcP5d8FYl54BHbx8c
xWy086cclOigiyaE0nnmUqYp/GePL0EwvAcoSnzK8uZEp6Mf0HIElbV/KHDG0ePU
jv1HypS0Gl0s7gF9VGjTMrcgVcG6O6YkBgLKAnHOQhOZWrFtqrA3Wkz0h2Cf7QtC
PRjKOHX/tY9jlsynH51Nx6CJ7qAe6m5II1SlsS/Mg9c3QrYOCn58KfV+upVLqEPd
woM2xeHqV4hlJtiy0ObXPSQ1WHx6rf7Kq5UBolT145WA+vVzBX2uY3vhZ3L+EOjY
FBR3hTjPLXQZ/JhZkd2mTayuuryj/YRN+Y3VcmEN2ngsbN/XBnLvBe3s6f+WS4A2
hIaByZlZ5GJdIGY+LOn7rIowXff90IEdDQI1sIepm1yFw8XTMtf+1sm8qhq4TyxV
vlIBbRcjxbTJbumGG2jDbqiWbeuzwKLYJNKmBObdoAv10VKIXd8zqG03DYL2Zlra
UlFeMIbeTtNmOC2+quv3K3ZvtCbiz0kFlADW4Gjip0mQK9TT2BhZ+ujxxlbDqaZq
mqj3p7yDw9i2yUa4DkEdTb4eZIef54AUP2m/lTD//EnIYyPJLk3aHLiQjC0SUp6A
589mKDxxb8GmY0Z4pIxcUnu/AeI7b0Np2350PYCWlNfh5IL406fb5TQFUpXIZ2O8
4MIi2mlOhAl9m5WUV0oj1xW8eOfT8UM4JSfY6GCLEgLP9X0b807qdfVbDFPpCvqx
gJ49Ty1dPxUj8ATi6lCGlXtrugTfAaT2OmPQ/GONhOjynxeIHIJQyhrqWOxMVcKq
8dnJz95JfYO9cqiA/dpOvneNsEkT8m8UzqaWmTExWOKqoKgSKRaxNSpjUVaEyHQS
zHNtMMKkA3Aoh0az/JyA2pnIjq7W9cr77FsG68bEDwCgeS+Ksrg/eOc2LwW50mHA
QWrK5R7MpjegEmInnLYVdO82/GB9jiA13GgbQGWNZWnuEreixZu9Xc/jLbTocTXf
87VPAfuksy1HkyXAYk7iFSvTucNdn6y8xSm4+9kNCYkKT9nvBKjJNXjmh1Z1cIkt
U0DsihrAv69bosFl+sLpr6oJh83skj6+oBZ8ycoQQp/zwiwkUJaJW0FoEKnMCCKF
RsVNqlqe12x1IezMMdMTkXGFuXS160gmkkT7CAXfz50Grfi4t8f7j4e2E33YO61f
4Y07sY6ZNDuvkYikQSoqqxI+GDjFrq4p56Zq2hm+GUnGp8BYALHC9L99gSwrkife
WRcyB5uTZdUsM7moOl409P0jHd5gVkRwKYvXdTA4jp4Ata5HH4GDNCAQBCbdhL1A
6Qnuk3KrWRAtPiIBYodp1YCB3+xZAKnemCLW+G5awnFZZW+yYtaVpauwAMoLSlE+
2tFcHZ0Pc3qLF/QMsLBl6xHpx4OvDvoxqQ6lVicRmf6Xhc/Ryk2e3G4ua2S5ROvJ
jFUxt32QATkVmhU64M7NtAOE5O48kAGXV8++J7PemvGLj4iwtVGl45jyyyTyA6OP
EeWi3SsfTjA+3SceCMaqnI1S/5MVcM56UOi3wzjMGJAkLImqz/haVugr9GVaJFMq
gyXb5EKOQJqLDF3n614trCvWTPYRAn9pUtiddjprErBNogRBDdKQPSQOYLGZz3Ul
vA8KAWoaD12tNRe+KS1oawroH+eQ29v1QR+bJsq9xGKWJv5SNVMz6bxjHjd/PdBx
LwAyyMCIWMKgTHSsfKmrSjJh0ua75MyI6cZpFSbTa7jNsyI3THmQw/7qRsyR6mPY
QPYLpl7NxN/QcahiLxDyP+xEg9e8OqiH+zuvltKsJMPKzRRTlzriEftONwhTd0JT
fkSTxTwZ8jxFwyxQf6ctHnQnGg9nsCtdJ+aeVeaxXsSeFX6nOXziQLBnIo+qjjH4
XV2mRBPqd2ALDmGSynnGTtLNykJY/95W+NQGSEVeh2baXSC6i73DxSp+DK1jFZ7B
e4zUZPC6aBrXLzi3FPvyct8zPF40DlpkAvXRaFrOYDYVrksubb6FJHWyiYnXFnRb
jEDnQAqeziBCR5U6onPn1ATWyRRG4IaWMNjurwkxtm4+aHky2JihwXt2b169en48
+9t5A9OGO5V63AcswivepDRRXy8a3bq8XSGIOzda9S2dR5TDeSpWLcuo+SrLaT0q
uzssnsV/deFH+BIBtGROXl3mUejdtzd7xCVwQzSenr817W28U5cqdrKh3t1YUCU0
ofRr3GXm5fJQU37lu7Fi3RLHcxZjESpiLIwIp9s+RVuE5C5G++ggRyrsOiYiBCbu
kXLJ8/B6GI87TTJKomn0mz/s0nXj77Nl6kBbFLJjWpsQqJ0dIYzsW+lS7JYLsBqL
Sd2ov1jTLTYiLBodRuRMqsecSFEt5Tplryx9ua1Xid8iXBjLEggh7X4lMrLR9tKs
KM348gsu9izpVXioiPj8zz8uRhPHCd32ws7pVLgWcQQgjzSJf3eX2772fN1TMyfv
b1ooZ1TzJB+XekzGop9pgONOxInsbux3WfL6zXdfsUXkgfdgHacQctat3lEJkCNg
QdfDPrccr66Se0KPsfL1yYOHni5uh6cbHriXWnd/WzFuNYCJlD8z7yrpmfBXeiRV
FKI8W5EJHaUmX8gZJ756A1UaV/pE7tU8ZGUd0nCDA/OEx4w4G2LYWPqBqN+5Il3Z
JqC8QUnbGWKs6z492tzJK4OiTUuL0ieiwjPwIplGhP0UOoLwSN4MgcKmphH6jhyk
irFXPADANBrEr1gReSbTTCG/VhQI5KajXmYYUmmnU41fpusPuckNKJBjE6l0pxLn
v7waK6vmI1RBs2u5ECG9E87c4BRFpMZfWSBeG7jwthRojW+mReCeURqDw7QC09Tw
hGFDcr/ViAuk5YXQ3G4Wse4vl4YcLq5PaN8hTuT4XyvkzhTlXdF9L/OMakXFuap/
vcGFMVa72xfDn5kfZ5veNv2BhsdWYm6qlY0T7NzhgxYlgOj5YRAk6Jvsk+1Z5mQo
NYG/FdQO8JRoUSS7ct/XtVIzRd+7rDdvcx6gNhf/eVRFcpVU7V217i/x+G0wq8Hz
ewN/ZcxASBUQPr6bLhhPyohpb4Qwpu2NELiaihL9la2wp2VY/hgKTbwVmgOHmoCg
I5hY/QWAvBGaEfj4z7V9cLR0HMpfUriRZ/zOl2U/+4uJ4SyN0TXj4Mg/AURS3h3G
9xJOe2NYz4mGfEH7nlbo5do7YAe4CyIP3swvd5+8SDL3YSt8+RjGqzbLPZmqUrVP
swdKq26kcGyA2GUVUE1WRRaFDFuUPRFlp56J+n7M9UfuTg3TnoEziAEWxsHGQHvG
0N7wO4R/mWEDEfEUkPv1/UZx+qY8V1dOH/son6GCO3iTD6ojK0tKskdR8d+tNveo
kKSma9HW5+UFYuiHr6cH3V4Mp8NEeC0m/PQsei/8x2ACJNQamwBR28HPF4oaaIZU
SvBPeVmD0K1v9q3yQ+hHa14dYKr+RhdQ2ju0VcsddjwVPdH3U87vg8mwFfoi2eas
6o3E+HacY8qxPLzjzYeXMvLRqHEkvC4zBytKgemQIiKsnpYi51tuzkWamsXsM+/4
4To8IWPtFScB61+QXx9Jc7lEG69mOYoQyhtnnbA4fReW2ny+FLMuMaXnViA2YmeT
O20bvxRCJXXwem5ITcLiGrAP+S0k0h63XE9EVoHvBDj/4ceGIxxIOLIHHDS4bJ47
Ojix1PL1hHJzMZdh2pDlG3A7rK9VrWxv+l2RNGJWKPbCNHTBgYCOaSctxOeehMGJ
9cSiZY1lnmMxek9vzuA2ig7Y+ERgK0hENviFtljighWWyW9he+/Q4+PbforFoVBN
drdTzojBGgVVoHQYKBJtGpLA8/Qo8mkR5bxPQP61YtVpIyj0KJMZnuHeEW48VhIf
USUBH5xQ/6z8jz4THkAXeBxJas0LR3IIXlboIux7YBmnvSr+RlWdAFfLP3AM3SQ5
mqsx4FxX3DAk9gKxp0PaGqb0J6eaZfFLbP02B7lJ+RD/4fx/PFuamJ085DUCUShy
qpcG1RdHyvOrjlHGgaiZ+d/GFcuYI0a7uGZs0aYPhF2q1KVZUcPdaRCmKNVEN94K
hnBQ22Dv0TaGqPqPggfy0foNBoHd49AxQXBfLuXb5h+SYChdpCnG8aoSF2kOO0Yy
eqZxfOM8he/zuyLXVnPS5FDqk1j3Z/ug0CWMvWKpw4y847mPVQQLMlLnHrhZbLoL
nThOT4YBIAImMpDDrMdPfC6NLuX0wKdeULhb9ZWZ0ZD7cH5bJ2j03aUsA8OAskOX
1859d5WXv/Z5JZaFlf17GlUrn23/bkClmh4q7CM2UCohT5qS5qBftyUStAmtj33y
83DPE8nByZLkDs5QpxQyDkdb89SEkVg8PzBVCa4aoY690v5dHYGsq/JKndjEYxMY
iP1wJnVLDnN3XeePjlHpAsnufI6Qm4TRc5KVCiV9vpx3IgVdM11uGUfqefdcDqip
EHivcbd1ITWpDTChUVDkDKnZy/ET87RZ0QO71ljqD+E48n2SVhpFWsiEaKeLvAhW
Ps9a6d++dObdWH0np444mCPkUWGjD7Ai8k9AzUQRzaZBXQDnlXORqwyWGAwcNBEP
Mx14XsIVp1TrADuQT3Va1mCoL375obQurD1mgLWwV18oT+EfxEKpl+R5G2ip/5/a
SwCTLSYGWu9tYLwukLJCkCD+Xo3o33NEbWn9OG2uUpsrJHZYF/JY/y5FSGwXaV9k
tJquOYQWbXW1EAqvFzxZGLGT/vI759qf2zqC4r6/3Y/bPXVsQyhAckI6zbJw/m0w
U8/Yd6M5YnlYTMLu2JmVzmnXk1sYFDCr4qE0fohsuZC6iHFguh6Yb27DCa1jXJry
Oau8hcXTwThxw2yWtfjS/f9h8pDlWFe9uorpB9W6FD4mN1YprKoz1flTb9ZGPwtl
U9+BFH16z3KXjj8kk/jazM4jx0KbsYzXXqS3nBAElKxx9w8PiqQQIr0/Ud2qsaBF
O2sQe5hUfSHn1tqS4NCcXl5Mr3I1DFZEFiMrWCmwE+qLrIz3/ZRbhAAAfIaPJ3oR
nZTdVf70T4/jS/tYDCVbQHfHGyNI81ZvkfWedy4FBfS9SiRp6Q4lMIVtFfznLZDO
Hpn3La/opUKoeLjZPhmQ4+uIrL0pI0T8P2jj028i0lPYDuXBwrsy8u3gpbw0jaxg
bmbO3ijMjmeMMH9ypjW49gVyjy1ffCTEPgIV7JxBylGSX5GFgb+2eQFLeQ9Ut7U0
YLpXhwEyP6v8Fxmw8J8E+VIJpPgWVDbiheueyasThpqxVl2CTptiwR+5gG8d4LRu
nm+E0t1MOJ1Kk6VdZaXOmh31C0djmoN71XW7zP5592mEa/1Hc+NnnhDPedHShBOC
dQzCl0hz6E7zi0KGb5M1GtXTfkErHh/iF8oJLsc5baI0XkpFXKcsYR1MM/Ywtzwy
DxWJ8ZXcDDMzqfnG00c/wAKlnAJ37re8JVARW28PGpji6pJDLoHuoWwo0ceaPmQl
BINWQen1UWImLqUkOYY37meDAqBArh3DNe/zP1m1/miKZPee//ZoDXg3U+7LOnAs
olGN+Ik9KMhmpssZMDWeS5ZiirKwDbolZtjbsqzySIeHfT6pjm2MiOxkoH5PYt12
NCd8ovZN5Ug7363OCiNPPGM303tc86Rteiojz9ywr0yeuo6gKyKDdvsAhPwFFJet
X5t9oF4shFndmTzhONvHXGAhLdByPy/MdyFXmDFK06wwr5wFi5jeXJ8lvsArcuwj
vGYcAl3u29QJ43X43hpmZnNFRP5mPzIC9Bf2KfPyT+E7r5Z/aj2zNRlCBH60NJFo
Nyqiu7IDJvGbAnu7wIAkLTJPHYP99E0iSz35UtHZXvVne2p63oeZXSXS8sVdkIyV
Lb0IHYZu8PaN5UX/lkeHSFsfss3uetWMk6S9DaorJEHB7S7vO+/DX0fFWbUP+dL3
YpaBxesJw/e8XIqGXgs70voeecizrL8GwurQh4+byJostx0ijm0EHSAlozyz5htb
0Xd9b4RJflVDMQxk3Dnxp9qyYN1hm6pD/4MvxJCMmpk62gVukUjl7BQe31R53V5R
Aoav/JeLy3Ej/s+IEiLnFlDNWz69NNDg8xFnjDrY7BCTuyJom3lu91nB/URG5/Bh
Xde5Z+s+aCGRgPcGaMIXSJaGC6rRPynUBKCepJ+CO5CF+oQhjYiZYjg6UZ8AbVOm
7GjgbFIRh1I9rhggNdaNH2jhR9n0cpqQ/Ruyzxo7jSeOHyv03MOj2RGJiNOMvMC/
NycK0hZjR2Z3e53e9+xcCFbdFjfbvRInbYgJESHrBol8pKna6JewCElXMWGu8sgn
GeEDrd3AmAlwIMooKLLbJTaz5cSZ4beBezqO1swT7qNkhw1b4dHfjjzs/6g95QFp
wCyrjW7MOp90BqEBzBRdBEwlb/BIDgHJx/T5ERJZNxqN/veyotmhiqxeMf4DhHTW
X2daKyXtmTCpRTNdp86HtaHVz1WDWy7lI4KTPe13tKWpLntftrhNiLCJPcTzSDbH
1IQUJ5N8a/25nOHxnJMbnP/2UDeO6l1uOvm2z0lE6q/eVPZXkzY5FN5tp81R4p/i
JdBz6IV+NGWUZicive8TwL9oBaXc2MsKngSY+KfBHizBhaMVF2Am9WEYYW9ICB+2
fTT1musbF2iL9xg7SutpZSncwRX95SQ59Tzn7bgcOzfVXy1F4xyxHhmyT2LmlG0Q
EBJtWgNtZgc9oZDCSWoCjxyyv4h4djxO9wSIx+oqJlIsvEpM/HSK7ioFT+zeSRBd
QO8KdBL0XD1olQJz4PUMAZ6S810mpuZv2UYB96vV5AHh7S64ydVPYKBYrJgCkS2j
D8s2AoMFFO109JRUo7biF9BZ1V5r/GZg9W69eMuiZKpL8xMwNaAbeanOF74bdrgH
HP0UtI4+8qiNWQqqANR41sYD1tLchiQe+wy8TIbMKkcEjQjEzHs+/QMFje+zYp1A
q3loiHtFpY+CKmR1DQamuWj/+ap8K2La7zYO66iMFOvgKsGrsDGCzQ8aOyOfoFWf
TlzfqBRryPo+5W5VvKjuy5CZJmGYLHbgu0s58l4s1+zsP3HBW+/dykXaivI5G8/9
+EW0ujGrAxd19Z5ZLEiAZP1EYvl/XKM9WsLqlNZUy8Ov/AXr2QvuGMo7VlmXVkxw
BlOEOL5z0InpV86o6iLnhGjLiMsj0SiYc96NyPeto3egKb36b1Iwh5Hfuwz4S83C
ipmujOXKPIa7Jjcta2BC0vJW5SESGB699M42aa1L7cvMilgyTHxIxOhlNw1fek+/
q4CkUZ4Ek5WzayfSuXS79tezNkrkOPcPO3oHl1EP5ltW3/qYefDr84C5J9mAhkQa
1HyacSYt36QDIXee5IllT3giU8fGcrw/wvAmTTsE9zs5WusJQUUjGjwZQQ/dh3T3
MRCkxiVhJH3e5Pwf6r0u/MdZGJKs6vrBwpNwfmcGBnMZdVP+qP7BOYlDaDkcC9zV
53awQYTkQh4GxZc/P44tjoZ9k+tDnWYqxvARAWZvpwTaIsQHko+XTqt6rr3qwQ8F
lpazL6fCaOyl74mxdciHw2ibB7yAL28+Ad6Eb294rIk7XziQ0IEa0DKXBCbnMPPQ
ymFdQISAOXZaKHN3GnPOMOluMcR8TisQyqtM1jCgfMaN3WhHA1IT0+ESrgH8rZ7J
5ILq5KNKAt4BL5GCjY8MLwX7ncBwN43pN58JiL4Q3r6Zo5+vGrThJY/WqQa6x9Xx
cDm5sn193tplMsYnepNUrhi6DC+575aDzSO2l9pzj+HVmGg/VXjTF2xslk8EX16T
RdVv8IFyeTeHomJVTo1qd7yw7mtPy9eECbt2ycp+oc2QFbD+OE15ab7QrxcD8pbv
yMuS6x7yClzjyZxrcW2Bn0ktCT1JtXfzD6YoN6/CHLdPSV6Lc985hHcPPBJM0gzP
FY7jt1Cx5FwPTlYVk/yUCIajXYfmRQMI+6StVFSdI5EBfT/nZIBIIUA/fUvysRk2
l+uacNS8dn+EplnYRKOIVLzCg72cw5RepZtN9Td6QcImH/lepOjtFUmcenU8d2RW
SYw5zhm5CP3XrV6NfEX0jxIhIF5aQPOH5nM9uJ+VeO8dryjI9XNaAXISxbPTpCvH
kBOWVfSvrw7FlneqnY9VOE479rj31ChkEAEEiEd6uKrzPz8XeWcZJZMncE/dIVK5
104ghDMOEzRb2iQ9BzmdNA1yitCk4tQXlrsQETEKw+Cm6miwliq6pk9Z7X3etT9z
UNCKVKypwecWB1IpP+aSpjaV5LPeQTiw9cHpNyNVARRVsQvIFFJC2B56pCw+oGC3
qevXUPBQUtRDlCl8WY5P6Mv1ODEhIPzLJYwO8SA/i8MiB9j4xf/2kOdKX10KvHO5
enWtwWhKe76I1ZVfgDcFpL/IoqfUfNyxQnsXwcGAPRFVastfSBgqzQClJlEIFKkV
3pvD4kVuTYfPdDbLM8C61TmxhZxz9uNXNutUweYNUKKwRNaSScUw3k8Rn/CBKIQK
5LugVTsAZBpaqTBRxnnnkB5xK9fc8zVp5rIdsCTdX+RMuSOM65joFhjkqjK7pbuN
ha1DKnUIhG2J0XQlndPSEtbQr4NaZDVV+qTqOthj8jXC4jXQ4XZ3GEFgh5y9CdXd
Z7F+ftJd5anNwsE+9ZeT1l+0Mf6UAsYQusNrC8IUosJS+V0eG8dc5ot0TgP7Y/p5
TuZzLWA4Db3qGV8k415pwwsuYdhRUXj/Eed84GJ1HBq9BaUQ1AGLY/bv0zdPvU83
E0Gxm8JcdBnyM6UAUn/BJLKKLin9dFUfaO/YU1T/XxPFaKVHSlAnzBZmg37rPl0X
fsbkV91ovH5VsXYT44ITxQJ5xvZMGgkdKjUWFaWok9HM9rFFGRIvnCMCew9Yx0P9
zZ4ZOsQOjSDBx176Zbb9lBE2nyNRAd5bwhDlxlZd7+M8I6XU0dT12FogBeEqkkSX
dQkB3mtdNVCgGvFx6J+dTUQF5glH5wMHT9ErpmVwmOpxS26XmMIKZMpDJU8YPEpd
83RbTks9NEetYmN1m68QI3Bsz/pbo/4gu6409udNT6v6sz0FoE0lvj4oD0eE75e3
VBJrwoEOwPIRpDo+touwBxQHPeCCJbMzIOdfO3wJb404TyqdCnABjvabKZduADfH
7f1yGn4MgyCcIR0FtScbL1lBsw1Rrtzi882QiRFYaBNZY2PHl2zZsFRYdSMoPuwk
+msKWJQhbj0HByLd7X4yTRQhZHIG+L4HPN4/hrQ5e+4JZWfxdlTEu23qKP8CZVig
DFFnfy0lioHrSS+j0LSN2cysidxpNg9MP1jU3sCTpEYpCUrngEFKSKgeOK2Lw1vO
G/Yqg4Q/J3bDUTlbnBV8SBY2azpEYOQOcvqH5PX6xWPnEN3ZVVwyxOOtE7of+yeU
yDay/DiG8nbakJoqWZqIsKCl2M6HeVYxuU7GNmRWpPQKZrkdwQc2XleV7FswY9J/
3T+XUZygz+7eJOu7Ap3kMgwosHcKQ5LcaWmgfc3D5GlqyTC9zhbAmeM4aHScXCP5
/2jYFh+xvO9MShh2wZq/KNIilCoB7s55ltkBJWbwzm1Uwf8RrGwPT3gI3icbUrT0
KjtNB3MehFMmAETdBO5+A5l+m1+ogy8h/5lAvznctnBgJ7P5FHU542Ah2dWs3I1O
hXY6WV5IQMgSNX66GyKU5Yf4XN1JqEn+dCHGvSbu1fVDGtH/M3EI0LgJCgdLG+UC
E7mN93TLplFtdNLklHDwHXZp4VbCUqMbSfgUotPjb3W4SHHR0EaIC5E19oiChkts
az04lZ/ZQUnLKodZQ8sEirZZsqHMZESWjxaxDoDLGmdT/qfoA5sl9y0TnkE3sjUi
Daea5ZGBg404ZOaLU7A/GXMtPAnWCHbt37WQ3zMH3Hh39b+tJ2Ln50ncaRCfYGK1
2WbZj+xkQvkd/m2jGSWcJ6vSTMTLQdEZ839krFBenXC1otX6KQDdJmc27bbDMTVC
EEGp2qE2vaVg6nMMaXlXOtkwQFZIFn8nn2u057B8Toh/3AOc68aYk4wgUR3wSWtA
40We5T1lKHMYWaUiKfAPYUi39p6NJKpkGljKpTDHpGOkPh1j9XUYjCTwb58eaWAa
Bb+RLLBgTNhdql2SYtCHDsaCDiZ4SEDK8snoey2sOoP+keBcTIv19bJH9LXYzVwj
kAAs25J2ltZA2w/6HY0zhX68CNGCc2E79Y33UatZTCA01Uiqairpp/EIKANneMg+
jvK0GN5uLKr/VYoaKZ1XYq/6hMh/CNfpCuRiBrDgwI+s5eYqrK31CrcpEfJ2gqiP
owrJiWAVuXbrMFR7BPYGnTgPtOZsGt3rTXHLfxsF1w9OwVoMtEIPQfG1GCYq10fV
vDryPWt0hUG2AkpoTP7BWRLMPYW7x9VSu1EnnMDvjHKGdi1A3gteDQOq+fUADd2/
LnrMVbitXqXXY1KbF2pZR6EvzxP90FvfdCcr8lR4dgaGblgqVsy2DB8+E3hcqSNL
P0jozz0YTVwyjcNuNUnqIazktWvcH9Ivxrolzhtc+0gs8/sTiV23s2lBvVloHoTS
8iR9iYV8WpByZcf7laKZkx729dy1bnrd8SmrGnDMoY9e84zJFoFf2avtjXBx3T9n
cWVTqmpHsWqLuONwmbwvBnQg4SIwpLUIYm1vX6Gjsm8KEXyaXce/ml80CFUme9rR
ZAGQ4H1YdW6lwtUBNIplY/CDbwDS7QnVuGy9y1NlWGZqBrmUijF7w3g1Qhpb32uo
bieg0a0yqNyuqcwMP+2+d/YtRWPv+zEBhT+Z5xzf3t764qlHS67V2aBZC3vRf2ep
vwYiPNaMnxdo7MbH5i086Jao+D/U7kK4HQuKRL4vj9NpCDewvJG9VqdjObJrhuu2
VcdS5SQQh3r8H7bmZCg9rmvwrYwbcyCdHYkYb0s1EueD9dcRsbb9j84p5ZgNgMWG
YBjlgv1W+JuurWmioeyNaVLJqnyGN41MFt2FVPSEfKvYVlSLkffXSuTQ9QZ8XKqY
QPkL5OFzwQtwcxbmvY0Csb+2cCFB6Sn0LD3qcveRXemZnvNpCwUDUyNqv48Iquzf
dmp9/4uxTh2y8Ss1emjYmy/78hjAGXlrhlizUEgLIEvDW2FbmNdnj6/TAO9T/B0S
BgFpBZU6bpTewHTN/Sm0CkjppXxwl1TTr3HOrBolWV92exAZcJbgrYJLuYPaCJpu
N9kcfuXO9veN1LHsZ4Cry14AJi0t6rEy99EDqo7zvROvjG6UH32bep1LW0f1PxU6
HSCnXTgXMghu9tzf+76qxNnKIuGeeGe6nrsq4acBLTT0Fd/1nAVlpO0tx5GVRew0
X69UefklNrX2A2uaGQMMXJYrE9JlvtdnPH30g+Ut5ey3x3vZDYpNYtcdkYjUglDh
Qw2NVDtsVZseF0i3qCYsUGeiK5JJm0dVVmLceXXOuOtHP8X10/PKJtxBx2bYm2Ry
ix0/vHpU5d8VFNp0VQpvBHVQyIZEzhG3oLB8jKklwsw4urn0COp5o7v8crolaun8
J/t/4fcoxXAgCIOZDHDetdAC/OiGCBbzQk08B39NvMt0o39LFNQkOSKbz1PJOy4p
eo0OyzXWFHZkQcpmtSMv15FbQQ/v+DzOVwXDRjftfialrBow7H6pCQe5XXJKsQW4
XIYUeWSrLKhPpqifvOboFz1hAvt9j65TajitahKQ5OKQdHFRIdg2onwWF5Yxg9J6
m8Ju7LrolWVH5Ei54tYfbQ0d3vJees09wIUshCEw5VwXqskTW/vTWANqFqEFsABC
c2NblfnYfKTcRMqJsFTY1Rp0f5vhjErgNZi7OzvPqhs1AaL4g2yp01jrHOQVJHD3
/I7gwhx/0zQo6yjyLj/g5fvGEOf6Pbg1AHZWprcRlVOkB4q/FWRvedpuAwMp4dOw
TvgRm+2FH8SpQ5j/Ggv8+RaZpjEaGBuR9aCVxiJgLULgH1xKMw1A0V07MNTKQ1kL
Waq8lspHBScHNCyD3q1eTG3U5bhlLSeV6ekrxLf5wQOdBpLMfJK4SH6R/Hp+iZ9S
MOxvC0mcZHXR7c+Z21cXjPtVdH/5p8hBra0MFDvlmeMY1xSS7kl/z3xYZFHQqvgb
oX0l8c8E3ibUAYWx6A7pQPAUB8mxV6e4uIiPzBxN5uAfR9TZYRGItnFt7idZQCC9
B8OG0oq/fkwHTC/dK2fBm1zZI6rd8XnnkALGvg2noXRXwUSv7P9eZPkgHis8O6U9
WRyENRybw7LAKIWr8ksu3d42rsXXWriA2c+ffaNyIOnj9Xpo/NDU3ribnZUbfhUF
jdlooYHW2JFT7IPP+bwZ6g89ekRrvk+YOJ70N5EITe0snfgWnZCUqVbj6addWV32
gzhPD1SOXrsX2XXrfuvgC8Blz0qPtHCGVa1HGAky43e/+8KFCQKQguqTIGhgaxZK
6iy9UPVpGO/8LhM9RjsZ1sM2JRrE++gXyrEkYCTC3jN2o37BkUQscwalU4FpB9xF
jAw1MvXiPbCJMA6j1g1vk/d3ADxNm4YALJKwycZya18avb8qKujcEJad6kfrgt9D
WC/j9hydAADv8P+k786Ux8DIMMFNoWhHr0Ya1itUds/XFqGsbZriHU1xeIxUjIdi
rNiXO8mTT595D1jzqwjDyoJwqfH6QNMVATrYT+v2lVXnu8VaqX/g14qpV5b/jjEL
ouPHUhklXz9cVLLfQViAFMZ3XpNec3iSzYynZHkUZYuK8RMnNL6cjvYfaCDLlMHY
3j5GIA5vWuGJH/iNmV/bpLYEN9diODw0HAr1PxHi6zMNZLuphH19rO8eNZ84gj8m
X9YcUneopPrdosDEyNY9s1kwdNddqy4jlhqgpWFdrH5OQTFDOzKCVU/7FJpj6HgV
oHuvo1+V+FPBjdeXehWQkV63JGeVhKvxLwI5KNHMa3s1Cf5vZbJ/N3R10J5IrwAV
9KpTQGGo/AEbn5XoT0fRzNX2h57VgTVEcLGRonbHGdemZIjsGUByQUbBypvzDpMS
g9L4brTl1JI0YsoJFf+eoO6WuB6/O4tKSfjZh1glxMGQI6JKy4/6E8narB6ApJNd
AU+t7SMPZ4SfGyFGqxyVHT2G+25bQ1CjGECg8A2/RTIbtp9tDnvC22wUeGs0lKKl
6zN94IBP5mYLz7jt5AuIj142LhBkuDrNMpTp6vHSLpXjfD++lmHPeHII3x9c8MEF
24Yk2GRygEblw6f/hoAMU0SyUq0zTN5cSflQgnzsHTLN3WhXsydfVAMxEcq7OPzf
aw7t3zHtiRCErWnmdThX/FchRnk37KpM5fywPr/iYXc81iRxdNbWIS0O4ewH9AAi
fbNCQBzPct9oJvaPBR0uLtqcpCmMLf45R3j/GZ1frriH/WMYi43mkq5SWAA0AQEo
gfZ9UCKca0G+mEbsNgPWUHCl6t7yuChiwHavqm1QDpmCcXqcXGuhKZzZVLEkQ+3v
priwIcC34C7IHywQhi/lIVeVexLaXtuD7vByKn31EINWl23eJs6UiORY4tVzyM9U
EcBB0ykJH2DjhXXlA4o8EtNhyUInK3VLjfh0htRhOfoW5iuuB83NACxEP5B7O6Sr
tR7VbL7Ax40VMUewe5Uro9gTVGpbuSJPNjg1KtAZky/wc7FIYrY2P98FU/T0fSMQ
4hZxEuPAuehnhi3A1rS8V9LFyNVaouzzkgEQ9DiC6ws+ul0x0Y11UrG+28oHCGr2
QTr+Vj6VgLE0Li0O1m2JuhOn8xXgzJ/y5gQ7gZZQOaq5TcGgmehOKKjTh/ZEqqBc
TZoLSy3y6piXF3BaU9rEfjRptsGdFzp5Y2W+fLpKBCicQA4CiDPG5XBWzSCjTDDk
OnrL1jJRDpgzSA976EctDFxEO2nA5efcrZ8hnzuQSjtmm38g6JoVp4O/NKuxjHK/
BfDISmbwarZKCA2vsNH2vS9YCBNUOH8iPoT5u8YrlHNgLiNhMoB6NaaAiJbDnPl8
InnKXANRyfFvM7b63Sn2vOWoixJEkembuC651uAJpkmarJiJbEMr7WhRK3EblQAn
Oxg+fdFyLaP6+WpytPExd4bZQVcFvFHoxJ+RE0aS0YWjNTvj40Gmx6WVxiDcAyvR
PP3OezbW6jMH3ImaZsUDGmOq5+eQJqqOh6jZ6Kvy9JI6h5tA9GSZd6/0HdCrjo2I
+64qpkoC4QIPmA5PernlWdCa5Ro6LLB8i3AxgZH9GRzO2E2QwyftHHhnB4dnvOfW
HupGp5Nk0lktJvep2GL3ud0+93tdCnLd81epx3q+VHbZT4fdSWcZM4kuINeSL5b4
fF5Djei3kNalG+1p8ZeZTgF/l8oTEtitat7BnggUO4L66tQh1LRN7RiBPukC8qKi
Pe+PkFPuDRMasS4XvGrogyQlfXVy9jK6hNvB+p9utOkHCg44uI7DIZQnQZIufwBZ
hj55+KrtNBjFBHXu6nRUw/NhPd/W5gnaiXyw1DJdXrYGMV4LP59aT2m4HbUP6svR
msj8IA+Kir8er27o4IeEC/wBaBjz27oYhGf9j+x8M3BNB8kLWxKkw3r48RVb7l7O
/0ZzLQAUzwYLFBeMTDvp5nFF/fnQalpVn3bdjDRGYYnQXZ1zdpF3zU4t7dBhYlsN
wruy2Ewq+m9iTyzN4AarroHSBj4CYQVJmsgaqY6+12BJ5RdRyXt6dEu58oVmAJoa
6DInixri9a580UVxLUk7RZOulGGa8rtsfPPv6de4BErY7Qn6vTd/FkYk58t8LXgc
Bax/TXYr3TqWdC+Re1W9cTK6KaEih0/NyP+nDT1Y7AxwAzgTWIUCRJpUeQAW2w6H
kJg0QzstManTOBZmElo1GKBTXJ2rqJNh6K5V1OcbVK+6Ll+bJaT4vJ9ZcNu4q0li
QqrXwe8/wpR0KDfPQJiM0UlR0FgtwZcBh78BhkeyIi1eIJ6pFQziI6CQq7uKXF5q
AVNZ79tsUOaUZaZmNXq0xUvjeqYZKBCxkKTKmhGhXYqGz5XyQA9o9nR2ageeAQkA
uFTdNq0B1WUJYcLmsetvDsJ1Qb3gImzvrDVJGIzHnd4wm2cwbaiZmBnka/jXrrzS
d030ahAm/A3tp3QBDg5QU0jb0M20uBZRygY2zPE6xgSHyTm96xhyY+W0HuGlVhCa
hkbl5DmTWOik+0Ckbll2UkbOa3moRdm+7XVH/bnDGnxtnbFyNDu8o4ARP0IHr3g1
OIW3NOcCPGdp1St/Ci5n3/5bN4jB+h8cMB4R44Wnf5lM83XdTxC4IY+QxJmJXff9
Yw6VMurHzDmyIjTpCPhQ/LSrlmsoWP74jvXuL34x2Uvd8csHB6ZVgtcPenRUaSS5
n03qoCeX5+8dKxaF8g5WCQdz1gd6INFaVe+0tRCLp+UoFs3KroWVyrsUyJAoJ4NG
LjM1EofC9B/7OrgGrJuaqTk8BRNKqAwEyezMK9pErehu0mymH4sTlPvKThNWmbB6
e6JdUsmzzuN+V/bxz/+8BYfNQIyo7BrvahQi5UVsD+Y8cQW6aof5PheqpeA0YLZ0
aPVoBcndbulj4dSUqkmHY++jOY0KpH1CFUrm+rC5qvhyJcIQ9y8XS8kXKk+HImhR
dBHkYz+rcvcSbVc/mXQ5+7/VaMfH/T7TyxEqYROuZGYxuroyI91VXkOP8Roll10P
QORkoPq8BIE9PJwyq7lx6Md8l2scJZ2yz7XIVCHhABssahPV6uLOLeJoFZ7AL3Qk
QI2YXdJ0+sP3WCPo8H95FLWpuVSTBS/iqwC/we53fCqQEuxdlRk5eSUAucbVMvMo
BbMfkKhMd8gwgkTXGo6on0iph/j77p8YhddSpKFASj9juLKBo262DpkfOUqVr7Dy
3yDllSQhK54iMFc+EJnRyXeBCXAhzRQ6062DPUU9l24ad2e+jhpwRHpsEL4XWWSK
2LxaFKTuLfM52J/Alm5eOyPzCYauVIUklUDAcd+5pTWqJbr0Y5p6WH181n1iTIfa
Glg9rnD6yDVVM0cPz1I8x3sGnYfBPrZc+JswyA89fF8COP5XISa65/TgD2w06wxa
sKhpET5rbLToCTQMDUtfPN+vadCo4ZF5hi3bCSZrKF9svO10W4oGFFizUVOTgvJX
eOpr/WB9Szwf26qEwP5PpTxvcb0rmTEI0RtGrnJiN/ZGUx//c/M1Rgp4kw2EnQYL
HSCO2JKOgj4kMO2fkTMQbwxXGIbffjWpx1J4j5870l7ArlfjQ3KAGRyi/lNstvBK
3aDlGQffdUl/Nh4TUhGE5EpPfOW2Sz4ycs3bEmXqZNva0ZL5Q4rhUWoAAHx6NLMJ
b/QgjyCVVTqY2rcGjEEPLunMAzYYf0S9BdVf/wj8Y3Sku3DoqmgvFOm0VMLPvMBg
b/8x8pfX/xQvYxyRgyuzdVcnIuLYUMDLBU8e9DSJc6njsSK6rjwYfYjtKasUmz0c
a5wSMpE+JlSzLr7RgBpTPnAqvfDsJNjIzphjGIJjtArN07/Jod3q7V7iBBrmEvtm
kb7qKd6sfMACKKfgUPt+lG2xaqPTn40FepzNBr6gaSsX9Yc+euUxdjwxNTqYJiWW
G+Du3VCh9Z3gPmTU3jVx9rZ4fI+V2MU7bOb97cqSFUrH3wiOpzzCw3kqgmrWonDA
XrDccOB3ix4wjjkkxRt1WN6urd7nX5sKq/7v1TVDiduZ1DstwWWZAKvGQTVBM7Tk
gvCVt3XKmWD3JiwHno15a7nc+amM6mYHJ/CaOalMTklNa9vrtZ1DcdNx+4cvP+Nz
ELZFlOQ4DyUfqzj6PaHDUCAcvSrhSgqc9Z8zOEvrn6POMh1Me7i1g6I6Sp6Bn+Ye
yxoOf9uqrts+wrbR9k7eKEyOd1SxOtADb/8jwrwXvXqEMLSqAPvYVg91VbdYhn+V
VkMBBZBeMeSarc/0mvYddGazWAIqKJ0NdQF9PT6oyowFQDvkaL3W4F1S2B+D2CcV
cN7Rm5MVedUllg5xoXqEQ2XVd+gRABsMh1UMnGkFUohsmkb1ST6u5BewWAxZEE5d
UXlx6acUFMYsEhEv8T1xO7X/dnkavkGfIHg/rfax68cSZhCTwqg4OUCj/Nq2SurS
/eY0XTsUE3DH4rpuW+l8bZMvjpqqN8nuAQU3CHZaEr0Yo46+z2gbQgUpYYtMlvVk
J7SFuzPR5k5q5eCGYqF0HpnDaEYJ5fiBV+KktzTMmXbQUO2qHsoKO134G/6LY4M1
pET9R+oNTFCXLtddpkU824tAEw2Ne5HCUlJF+tJfBnFENCGfU3G/k0Ohevi7jEaN
LXJr0nghlSTCwwEw7ibMgL+vxcsc8BM8EKRm3vgE5Qycz/n0nu5BLFikl+hgIXoy
DB8yhcvqicPoSKCT3BvIXUCJ/GIVZc2KSJ0CngexNoOvLworUUPSBHElR+pwoOmi
nNbV3HOLHnoMw3k/hHgV8Xg+8k7UtZYdVc5iH7nfeV0jvbVaTtBn7p/DJPYqHxfG
Y78rltVUd6moA6jhowdw12G7zRMdEqcq/f5fHDo8mcDgYUwbjHDAEV3B5pL2Uoo0
Ndtq0Oh7tGqsE/qcfzHerUefBBzeYFu1S45L5W0pKlAM6p6erAEzgrqsrA3at3tP
77E1QKRW020E4c//9a6ZACc69liNJnfcCijAV1FtWWUEgLjXwmOqosKaMlZS2Osy
TD6efXcFJjhaXgZxvL69kceFO16+y0PlP4lJGijCDxbtSpc4viOrW9Z449IrPAbs
SlUMzyEzM0SlghCWL3CKhvIkHFWtngRMGCAHOdLAFc6GZcINAePDPd9hjAZqA0c/
zcDoY5jsoKLBw0twcffr9HMeBw2xJrzhboQt/VSF6wSCgORgppRiDktgpeIT3xZX
zkJq2fhD86HI+Yz08AJapXjis9tQW4fUvG8bYMLcGG0yP0zufWTOpg8G4VGk56bq
vd1OdSW1m9oyC3Cxs5jEJ2hI0G6J28m9fPUUl0HvpsPuod9UXcAdlUUwO8P7b4TV
z6Tw5D4Tg4xdl/ku+A3dsn3Uf6FF327Wal9WrsF6ANvgMWHWYcfwBP/Cqcuu9jOv
l3BDSJfkWfSfXhVZ5V8hLYucRkzQ4FN32ycJmPrirzCP3E09IfQif+M2cANYg6Ev
Zs5ha8yxsy4aq2d6HRdZDFhV21g1ZoY1SqJ97xmjFGf2XHd/Gz+1BJqTMjvEfaT+
HRz6mGU8x5TB5HRKuzLAFvHIM2YRVjRrtuhNd8g4HIjXX1KRAToVhj4CYCO2rpRe
vIgESMqMVohsx9TeWidyEkSWjeb8AEqr7uqXrDatV5J153j/Fzn+zQE0pLepW/sK
h/4+U3b+skS1out+etRpnXNhFFrC9HCZ3A7drLOwoyCsRaRl5EXi5RbKJjETnA3A
OuxUNm+cgam4sZvuhNiazmtEHjBrHYsRG8WSvr/AoZzuraMkc1OARK4nbYYsEFIo
V+qFS/SLS6Lopk80CMn4L6SgyvaXq7p4M/W4H95eoqiN+JD4UwkKGWaFPJNEObOm
wVmV2ShTfjNUXesUrFU/iRoKT1I/fEKzAw6wmFyKBmmPXGxKiilD3i1O/02hci9y
2O0ynaLgt+CCTTYSdpGo70avuR+Ly7wNmKUCCbU4bfwuOKDmTmonCPAIuL4yagcI
5808pUFj7rceeyG1UBe0GE+xKDtR/6zlDenoAmPao0nLHYD+v6Z5szMSuLaNRoV/
DAtUNctcLyf4hTPp0byXcKGMCnHQUKfqybvW5fckOa6pvcA5iNztry+ljRoiiitP
1B86vAIeXWKdtWWeu4ybNsSwXlvrKBeC8Dt7qrLZbQW+GgM6aU/0InF8xJK8s3bQ
26ppFWoC4nQFF2zzweF8P3aq8b5EzqseMirRzrc36b39IN/d1gqd3F20vQeMvnNf
3Z1pjiArhqpBLPNfXJIqfCZWlopNvBMHvW2+XYwSnBDw0vTyM3JSSKiXGww5hGyF
2VdoE7PQPPItRdpoh5g04qo6U241t+6+54XSX0hLU4lWRLrhjjagIttAYVfAmINp
5feFxEmIdvo133Lfa8dFK7vogyEvBf7QHb/15Q+S0vxAW4xeOeqq4HxzZqctlCgb
AQ2zBMkezwqw+vKXl8MyCmij4jiWeHMEnJij4iS9amC6Rwcnl3FtCqQr9CW01Stb
8faM4gH588mFHglJ/R0x8Sd5o0WVm+bwtscptz/XpNGtdcTyU0ZnvA+p7kTIhGNv
om8GANi1/uXchfV2+D3TpK/2AHC6GIaE5F7FbcjbGyZQFaw0hLDHoi8QMdHaldc/
Lj+PPOcff6cbD3GKo0+c+3KwAMyOmS0+Yenf7XWPGXB6oiTtDPQK+6za+48M+sNp
5Lawh2r4wv4o08kJz69TxoC1rrNgyLkRvZlOhm3E053w7WAqtF5rcJHCgKl0R6xK
3MBli9Q6Mj6KjQ98eZx9JQRbAbyrFLOWahKYCkE1oBj3s/AR1H1iZBRRmrnaeq6j
kTk5U1sBzLpCYgmhCdwJsCDvR91zgfh2Mn5hsfIROVqqaaNFzKkLdMLr+m+C3hZf
uvjRiBom9Zda02F7fzVPGtdsxoOzuQ4FNGQTppIps1cuL2J16KpnqV+cdAao/gL1
zWqkty+3C8UQrRQHd5bBaxqwsRCQYAGsdXvQy71QeYLBPk0GlZEPkHXIVDagkRS9
nIYNCWE9zI15v6uppGnaej2l/oRpf6Yb5g9Eb/yCbMZTpb1fDIqrGr8KM1NL2C+a
HAmrMZBYvR3lJ6r9F7c2sARsdSBVquxXBNQsNS2ZMk4/60kMkBqXzKk4qF8oIfkb
rJaMMxC0HGWdeswd2S+uaptKueoIhz6j7SDdHlBiLJAIPO2J3nEk+LWZ1KtG4WyI
yF401i0sKhD3382oklc1L5HhG7Z8b/jgO6TzMrXhDFasDw75ZBv1OyitqCHNVVEI
klY9E/W7+GtIZpF4ZAghXwet6en/bMO7tk4kueHPBSJiS5iw6bM3DG9iqNb4yu1H
dmgOIYo5Uo9ux6x/2AVIRnCiIrt+DBKit0gKQOiavDsdLrHoRdc//7IPyj5QsthO
3wF+w0U3fD8kqvoz+O4fvqgNxMMpapkpmI1XVyvvBTNHm34ORNp4M4XCT5ElZ261
cqUbgqmlmCGtcVNW1Zsy6SN/Z2gkCWLc/slBg/dfrcS1e509mG7h9Wv6MGaGoI15
E1E0Dvinlis2/3zS/+fWTfo+bdlWU+Om3LYy+rgK6iFAu2NC44umOuTsiWMcRhVd
M8cRqAW1+Z6mpasfCxcN5xIjvpmyjGauV3FqNrskP2TEM5r7rptI2zlOdw1P0XBt
1T+gOW7JS4056sYVmf38uIEuTfuQ1LZfIW1eQvHogrE9AlePNoEEdNGznzEMyGkF
qiIiGFiaOLU+s1pmYvA1LPhyLFqVSIZZ0nUHa2aYPtnnhDa0k8Tj00+tahkFA1LD
k9FT+YlEKushbWwPjVxWnZuoSr9Tq/BXu/Lts83WjPXUxKJB+33CXiZYgX3Jt0Az
l8zZi1MxRmZ4sN5m+O0JCAkEiMzZA6kYVFbuBfcGU1YnRxuuK//Rtiotw5dzYgUT
Ck9JRbKsHdMuq/7fziyqOZug/mDlE+DbRkr1XERxk7EO4av0gIBsdjqoZw8YPBpV
4lmeTZhVU8d7MU/wL2C2w92aDpdf/nbruiUbcSl46aJg73iaIBPbIVWYGimauyie
9b+EOm9HuAnP6M/m5UZ4SpdJeDg+eQ7CpFJAd3lGR8px+axYl1M+Q2gkh+nxmTnx
fP6ZeVIpERpc1Tg9KqCTUCV8t+mwIiZBsNWaRwutzaVFeFrUswnrl/6fFEUqf1NI
/ckv5CXJ2I/n8jLfoT0KBP/V0vivOnUkItvsNUqBrkAHo4xQfXkO2AQASvuLaPvl
QthvhO3BLqlkc4/tZtXSBFxmmTaXbz4eZdy3b8d9NMLVONCgl/cKkVCTAjHEzurM
hMYPs89PapNy6OHi/tiN8ylazzQyWE95Z2vdrDTOT7YynJjVVBg8ooOiV6eJkegs
tyrTTOcluaw3bwaiBmDo8QmCvw4kwF1lrRi2K6VHwYY8/IN0IK9qiD0xH1n+bktD
kxDS1+HS/xFADOYKJRUotp1HiLeJ8zFMDSziPTsI04jNzixb2yKhA2S5N0eVOaVR
iVtHAP0oWO2bJ8O3P0GI93559OQNE+fLLDC6BWvrhP6EQZUPfN4/fds/XDAtRu0J
UBaT2Hc4mR1/07DUlSoUfsqOpJUViSA2w+UcwHe520b1cPZ7o5BGjmyuQXCLyZh+
TXqdcC3hUjrK3GG5LX+KIGqfXwa9Du47ZSdH7L8ASPkZA9l74HUHklkUXiBfqglD
m87EL+aDwZKWqpXqtweQ30N1AbsZCNpc/z7q4hpRXBZtYe47eSfvEDjDgLkJffSZ
85iFVGb91NfTvAk/AQd7vSe6zNBYx/zQnSco5uR7dBtT40I6qcl1oTkNOko9ne+H
+1tQOa8z57UcD1BVpFMj1u51pmdaRhBjFRC20AKg492RPb9gIy4k0Q9esFMxhxCE
gLArriTHmty9BthBHHZXhn+dMsV/qJby+trSn/2W1WsN707Uwc2pcNdwJ5gU/xI2
KhMfgO27IHjcpifl9T1DS6VwUmscbERUMoJGZkVeoe82wP4HSgRDDvZrAEmUmGDi
zfWwZTQ6Od09qgiFE8dp9sUnOTCkWJuvLI2IeASuLwacb9WOaQxSoPOjZcTTUypk
q9wZl3vWARuxIOsNgvPsVZfTFzHdk5Ob4/+or+HDlFmN0WeEB+o3CZzG5o1dupdj
hMeP7X59zXWfXyVGfZf64K0KDTNT/TgWG6U+TVBS+ft0b3eXVmFsREJpQ2eG35xM
d6TBYwTTe5WNplU6bzaDRjvgh2nPs26nnsjTKs27DjSNHuyVJVo1ZEEsiI7SFqeu
oGjhTmbDZPAlQQERohz8ZDpSzefm6GEH0UEIls79wv0e8xTRU/72xczKy1Q+FN5j
bkgUxgCc4ninBNNgm0dCF+1GWjqdXfVUQqKE8HN0H4LuXfZMZvRlpXCM6lp5f6sU
yNWpv3gKOJD1cSnoVGCPPcyVf684OiBloZbKhRhCAxuVfyOAJltzQ9Mw/8UuIdAP
ZUMlb6TxGoy2iR7P7VT2QqlimYj8PL6zjMWyZ7rChAY5/dLtCxMHecc6rgJH+Gnp
mNt1zf3etiHjmodzT+t7v32Ps5d0lVl6cz8q3rrtZPh2IQyfXz4YxsN4rVOzTjpL
VUgbgmKZPrub4GcxCyFuUP/fsREyCiQowkg0mFvt4MH/5xu4ko5bF9R1dffx42qq
RS/keCoq0Y+oTzEp3dqeKZoi2bvdHCaMMqLc0PQeUVcx/sIAjNpGZi7ffY75zvSE
P5a6tMm68Lzq5oU2EDQfchoE9Jw8sB4Lr94h5ajEs5QUytdbY1VNVpDmqa77WPko
EyLOFQ6TuDZ18Zx42jXXnsX/Exr23Hd7BNdvX/Lp6ahokOyn57Sw7mGURHT/4PwO
2sQ1wdZcqECQvtRkcbhxvL2SFM/zr1ICXyBVQSeOTXraJhPZ1pVbdP7tzku42Q/+
rKuwT2n9iNMx6PmhlGLvt6AEpSy/FdyVcIQOKxm1zGC/nUpGdVcujO6AdYRWrfch
C4yQiurm7eikSbCP8DnAFzsMcuZrud/ADJC6y7fkGCp0ugB41KPn9Uvs/Xpc35DE
EWvVVbkkUE9Evj/WSE0c4SPtFfHQ2+fH960zZH9uNXXnVSkZDpiWp0arGabDCeV5
voPJpplry7k4FYPRbR2Ksl1ljaZ6oZmrTCZb8uwFpsPjSej20ToHRiZ9Hpl1K7Xk
ysuv4NiOmCOUmWA/jh5n16W2gKV3gL2hoBGIoLe+fVz0kv6ysMwZPxBDi2nWULSp
TpbVB3xUUc/tvJzVVKcpbS+y8NYxZqNpnINE7JoMgkZseHgyDLnqn/SbeYDcXcw0
pPXvS3KBCOS8qlh6ejwRErocuHRhBChnFRrhVVtqjLo3X4uEDiBbDU+BjxFXff6R
6UAnIpHhkLUfaQzUbkPGuJdVD1o+LoUrNjUCtNPhS8Zz9j1YphldW1H/ymCu78g4
/7eEynyNg/n2lsOT2gVdo/MpPO7PBcxrQpuEfhTBbk6mYHxfPo5u95tg6p1f/GeO
mfT8hcCbyOrzDJt6hv5O8pJMzq1wJiXi1ypnd/wJ+muJWGBWLA7FUmQudX1lZf44
FZfPnPKhD3odF4gIjPuQJd4q1bgmHk4FRxSmCfcSvknpYPX4UHXIVCk8g+CnBM8N
SJJ02DEmKI1pJ3li/f9T5V+kVD0lEmVDLsE1C0007ov81JpXggWH7aNXDsjdDZi7
FYqBnaF2brgb//Rko5oUgfKc/ZVMgsuWCAQCVsdeW+HCHIPkRszSViP55sXbY6JB
gIAjm/w5JcX84OwtpsWpv+USq5dWdTE4/UlRErIJS8yN2my1B4KCzK+pvtbyBU0E
SGx346E+tkbElUbIY94NCA3Ub1sbBL9WpUXN8J3HktBRyH8Ec78Y+tTdbFKfMfGL
Y+MqSYsfJjBOoUG17IGn7rlkTaAPV6Szss6xeQfegFBXu4aQ+a0gmggNQ6WqyL4V
mQrJQdnY5v73yKDLtCw7PVdxvkz6nkHgCIAcghghoxcOq/8jWtZPHTUDp/qIJgNb
P9hzTDOEfFhGe5xZ1b+wxMEjCvR9bAemJg6PXf5egI1oef6IOXQSqoJzay5IXY2z
p7wGJYkjk9ZH2FmmEddGwPcdeHX7ZqCfslzE5SBkpI0Yhu+tiNW6eW24sQGT4F+M
ogrnQD9DVWtl78UzUiwKSsZSP+7xxM+9qVHgzDzBWEHUECzu8CXTaVhtBw1BNANb
uihKtBqWgiISC267J/GjfJIPhSVk+W0y3WgWXckRyriXRvaCJ7y6y5bW9g7jbGG3
MqU3NwRJaHEokcyZEZXzOv+HbFHLx1SEhRUzyqRH2igUc6C/OkVTeM0Epg6R6iHN
N2nk1G5xrevK4JQHwhASDfg6it+b+9+RTVL3gWfkdE/nrIZ2AXxrSkhUL8xujaeZ
jnl2t7OI/oxhH0kyao+lrh5ErEDvD3w35AQBrdZB4ynIrS/nFB/IUIsOU/bLDpi1
olAM9E19rRsVWAzOXR68KGVrNMaJiaoahib45RfCTLyqLtzpVPV/gpV+SeYcnpr6
hjc/KHjKyGZJCklCVaRskzq1MpSwF4DAhjZ3vsM2Gb3pHXTjycuNOugD0qDfPk2z
altB9X52M93mzJJ4AZFLPzDsdZU1LuzdgXEzBG4wFDFj4/1Z1TPzCQBxR2c4rJ8U
Jy8IPVFtYCKSIv07T0mwywHcavTLLM9wqr5HAG5q1Do3K1ZYFarNDkSZi7s10Stv
fnnhHU09Q3Cs8Ev+C50V0xsMdUm8+JGggi8mHuK5FBp9Na5gzpkpd6FgVkPZ7xud
Vk5kViJ+TqIIEI3aYnVNNJ2Rn0u0/Qf5/GIU2vXwn93W9Zdo+7wkTvvSCySAfurQ
zESYbz8SsiuSqia8TcxLOtaAkxOBm29IfVdYYkFKH9NDz1Z77xsVy6IoB1OrHCAV
2LDwF1h6RiPMM/nIyEatKXf2koHYvhujQrFIobtByNsSfBW0IbOcSWtiEErF7gFi
vo9C8d6Bc6Fr3b1+oKzctRDHxVMCHWo0eJkn8KQnHovyrpsBawrvS85pdKMvnE8z
sZpIunJ7XTCBdQhb+a0/kn6dd1F+7IQSa02HNsGhexdj6NUnQgDgvHkzjY8G2bjC
gNVU0KY+OcJtTGg6+Y0iaZNpKD+f8mbzo9X5PAviWLgLgJyOcx5ZouRMCYjfmdS4
1nVZv7IouGnbTr5QV/Uia6C/esJOuhf/cSslMUSFloFSuIAZLcW1TsHb+gm5AAcv
KFZherpQeSwY19DMYKiHEh+Twjk89PrEhiAbKBr08D0YGKPGTDhLbQdSV7ovXb0k
hSKQi7Rv/LGpH7sjD3yx/osWTER/nIYW4cmUd/TDypjWsb0chCtgfK9xkjJAZ8TH
xGFoIilDftvLhkilgqidVxqjrKU1ifhpKhvEBaszgdHJa5lnuUmfqkMcP7oZbmL/
G/gh5vdP8RElzZHdMduR8vLvOFBVhna7BDMCD2Mlb4Lf7yyjvMhQrqZwamxnC6hC
WaRV59wKk4leRZ0uQAJogFi76Kosa8c2DTGAKp59EGE+/c586OWCxqL7FsXzcpyc
fFb7tqejEoVRlngkUzBn84bAd1guAi8E0RVUU/Oxbxfq6uoc8HmNCHZCEQJ5wcIH
Ba2JCyt4JjYlKj2S1LplIf1jd9wbJ2axAnRLvySCSOUuk/CSLmuF6SdNPNmNxtM1
CVrUUkMgJonXW3/0sL9iBBo1QrHJRfxxkI6a+DThdubCZmRLtI5H39xjEEF5x6To
arMUq5IeH5jhOPO0faGafXmBv/sw2p4Fq677M7pUGgyx2zy8mw4tArTW0X4v98jy
rbl4JCJ50VGE29/mndCnvBMFcCHu9seSFpvR+LApE4PXdJsopPoV471gVWmsXcV0
a0GfSJdZp+VyPLMaVyx8IPGckAp1JlnrKqEPwP1f6vaiin3PJF1yws9gkyLZ5QWi
JK8fg91UsJD+0xupp76MIe6RMSCopjgjSb/GntvKXgyYD5N31hitfLSVcL/H4lQk
o0CC34aKSEKYahkU+d9zoPVTrOkTO/2YHj+KpqTplkSZTaR+ubX9mdshRuevFsLU
y9pc51K2e+oTbF6aZv45+m7AfIg0g2zsz+nGI2yly4bX/f8ZCoupEdkCZT47PlFo
tCTSJv0GWJFLlV9lYmmXhGloiBRonK/QIBSfd4IyndMCFJ4QSlM3FZKwJ+HQzjQ2
G1ak/kdBf39BSoBWZ89rlCMX14OtAB4iJ/BIBYNCC0Yy259NMrWJofq5nizd8Lzp
2NrG379Gu0V6RlnLdAxhtWS06EqVijldCzbHneqCGjuONTi+mW1iAlC67Q/HbHCV
sjsJN31g67SXVgDIhupgLDkaMHf+TowC5PjZdg9O5FsXXTr0idlUINCwhsRJ739l
pc0SyLdu8kr+Ko7gS1ijmPpnVxC2HfTX+rxW7d8nq2UU60J6wTJ4jpZqa5UuATcj
amtzH/kFFZ4SwtUYTcMb1SKKGKDmC9HvHQZsMMsbnEDEgC6GqKStzELVSolOK6cT
F4cFjicgV8fMVxZKrK9XFdATKpjjMof8VjigAk+Z4/dfNYM3/96KEiII8Ej4aE7o
sXfd/oC49Sc2lA+T5bZ6LpZQ/Vk48Q3bZCXjz4LV+jZwOvG4BdCLuIKE2JgC6rNP
Clh+/alts4ZSC5Lfyae4rqvVmAjqOmmW04tkba8kbK/Ct5zvngDqQOLAY9hl38wu
zqkPysED5DUH07GLTmO2l4elgqEWl9h31lDf394C360Fmh/2L6WJ8tkKcTNDfNYo
LROCVTyUgOZ3wtGkwflrTP/Hov6PNWIvGD0IWW5jW7+2x/aA5RlSnUbdMgdhFi66
S8Eb6FFAsoB+MhmBSQNdN/TZaKLlXUGwC/DPQ8LZXKNx30QlWa942Vs0cF0uFDy5
QNjcNnYlGC0pyA4h0TSlytFCI2lnz3sMVAY3Oap6x+LC9l0FpF8+F1ky5PcqAXB4
gdgl6rW3dtbLWkikLsIL0MJVSNiZQcbuuKjZ6qzNBAk/6IgllJF9x1e7ON513TJn
a6d8od+xrXUyqiAMmjpBVYhmPn8g17MIkJdcSCEH+pQolA3QGH8RQJKFfb7ICQst
B2PHKNtIvlxKyBL6ZVYzq5JREt0t7F8YCzxCQnHRjl1jwhenc02bGDhhpSgQuEb2
T7XX2cGcZH2GjpcL+rqrzbFJcwam1UMOSlq7Nf7uDQuHEDAHBFoNrcMQAyXn60Nd
MLlaxXxhIuI26OlfM2L82RjA0WSPwWUGDLYUjUZzHapxkQvoBuoVmaxzQcbs+Eon
chqq8oSfCx5zzjrSlbpJqzQ/yGfP1OZIksh0S7ACS2jxMLHoRMz4IT2lMqzTWYTq
XS7wKCywvi2zpgmN+1zHI0FMxoLTVNU7jnPyQjtwfE9a5nHffZ0q2sVwSlwGYubg
5smbdlqGPcwVVFk8gTX9Lwvi3vYfg5VEVf7qwIMgcXDbPB/NvNGYGw0IP10vlM2A
inZUbLNKfBWiE7RrLTmEThfXftnEJvl14EWlAwX9b5IpJYoAe/owX45C6NdxAW27
TwrQ/AL0dQbEYkzTnO/mZR2Pm751fqVj5GJAGWXF5ZfpS26DpL83taIfUKWZhpZ6
7GqoQYQDiMIY0Mrii2jf/lPJEzL3LRPYJOq1SzwQMdtB+9Ll+DfAto1b0uJjq6Kr
pi19WZEe/tv4ignmuVj19KaAAYzC5IX1dGYfcmQpc2ueFLwhNSXLtSwJv6hXDgJz
JJfQkinh3vklmEtHz40NNXXS2YFuDT8VLteFUlf/Pjov6x2VKpPjbdoJL5ecq/2t
Er12W+mhyJ72VvGR/7LAqr4KVcdzulPOl1c/Fpv2ZO/2P/I/jMAVS6UA34MOzMk+
CYI4nrnTWcFesTyCM9s4/T5P4WL8E4V/JqXoEGtrxUZOBkOOeYLFhPE26yetyOH+
ciGY5RE9mlBk1PbqmV9mILqgWO/hv3eAFSBa+Te2B+DePMaT0x2oQjHYNJ4mnvOC
daQKluZW7jChS4KV068nw9qTC1MrgfFMnXolU+iaYDajofUY21QCvV78HIzPo4WD
bmRyO6iVZyS0N5yDrxx8TvixAygpMAzEDtM87U1wyDZHU7TZQpqEtm53UISN51rS
jgOYDFzGuu5CdYynUo4I8kTCuRliKtAksqpTK9FnUr8PNj7LBkyptXw+B+eNfhxe
qzV7hI6UpScCqJ1BtjfUr4/SMK6y6vt4UD1FYA4/SBSGf0NaUABINZYZdma5De0n
Cz+ibAHbvOjMbkuEp9BaLy3xQcRF98+Hoj277v5VAgAjJwM9z548NTpzqa613JPo
W8pVoLzPBJGe01u3mn5ba/3EIPDfa0c50o3O7EQXBGCnOcaX2GItNVtFlsTzr0qF
HHHS1R1YZu5K8zHHGdJVZhNOZ4VKGjDlRnsGuBERrKmIPi+FV4bVV3/rma8Nb+2J
wm3gBx9NixGdqFkFUZnEn7KhKnJmZinEp7ZJMCOAo9wivP6hRLsYX8O5rh0NYN/C
REhrQy3s/nZxeTaUkw4vt+044IqwrauCT2poAmoVqQ6swLg20jkdUla/W56YxAgH
6XnIoOrOGwxCTtUBQdGJLQOqbe5YKCZ+NLh53UDtmkrOD1ErpWP8cCPEIVg+ViOD
Ye/wQkcYOQ8/p7icHxonXjFPyq1QWtCOhG4rcxUX+LDbVhShtSeB7ns3pdUfgC/e
h8NDUPGbATrFi2gFVoqKfAtJgr5Kg9f92FcSyrurabk7gl4xKrvCOWBB5Pdctoot
ImJ3xpOZDBXDEZCvl2OaRIyrKQIAd+smPsb4CdPWn6dz+4Z/Ft9U1AnRfDi1y6sY
DZHTCFwg2kFlhc0DazYUXx4tOvRbLIxfwRTOy/0+b4ui4g2ZJBeVGY51m7CUW0ZP
3JGiu+c2sqFlSyItRpD1p+3t8umt6DWvrVqewcg4hU4WdcT5FuyDUXJmErgnP8jL
rWbKUgms38eblAj0P3Sq/flOFetf8HWOhAgCnMz71LyVfFE8fwOHg3fxuYyXfbdJ
BvKdT5O0i490NT8Mm92r5SCbOpRDQKjJfgTO79uKJNDnAkivzxis0vKFXreGHkFC
rBIU089hrFzUFK9iHKSykcpckILh6Ug5lk0Ww5RbbHFuFaq/vBqqmuPF1BpDXSmt
I4TUW4LJ3rdKPoqWG/b3DsEk7aBWRozNsjFTOgVSi2CYTtxiPOhjwYsx82v+ZRII
4q+BSC4gAGwrqAYZGSsp3i8xl1cHwgAR8ISNeqaYE6Ecy+OaraJAv0FVqpKyEDC9
/Deh77AFtKRGlw3hRStdMna9yj5mUz5SAm1FPIotHLXPWSoUVTw2BQj9H4GfxPgu
g5GfsE5Bm+cfMOAbHknhn9cathT7A6v32rsueirjrmQRIG50nkFkFZf+4Tm/1Bv4
vSZPkR+ukF63qgMxPTf8f0dXaR14s1r8wnQXLk5FdzsDGHTBEfG1VKNf7/0KERl7
CSJXTZPGo2c/fuW7gT99uB0Rtq2m1JYmF/mxERrWyss61as0ivn8Ls1+UPRh2290
7n7DcIbUfklW43+bmd0bbaVJEGjEjRumj6TiMKGB3raRH4/ap8+TtHYfXgHruJ42
WMzk2yGMH5K9cYmUuQUH5P7nncCZjia3svqB8qWxJImM82F/LMY+ZCFVoIHNh2xp
CyjXAt5dMb8hAo393XiV084iK7IhpJ3b/k4woy8RjJ6J8T5eKq7TqXJhgNHZosGd
R9Ak7ZuGde9/8vSey4ori9WJP8pC7niqyW2VwNSvw49ap2qpFba2eDPzHiZ+UUVV
IHDb5N2c30WKO3GE+WsXtzhNqfkCANDG+rxQGw7kH4zl2+OAjuAw9w3R2rNe4eJU
5iKPvJ1HGci/JIn2Os1vt7lZKgOI5gTg9281ragaTEMen4be726THChuCDu1ySr+
Gtic2DJYr9PARm5HJOFOn37kASys7TBwmISCt3QvGwSJJt3wjA6LjdmsqGwbdZE2
eYioghCNz4yI5Q/Q2T3x0V+acJkeYmda7UQC9s1UdAqzA4VFNZFiJ97+FRQkwqnr
WLxJxIdFLhgdVvMj4Ss72sgUwWyBKr73CnXdVSvnmG2IV+gKz1tMl4J7YuCqMI3i
0RuJXC0OsZf+nJ+VdqiMIMGRIvV3+3a2lENbb89mzBX9eenSVQ2tqvL4rOypDMeX
X5GiG93e/Q5GTNDeTGb8Y5Xdeuh4hmXP+sdcF8PgstkvMMMV7D3o6s+t4IDcSFOq
JqA6mK5AVWNFcWIvyzOoWghLKtWMQolVKcTWNtsvpCagoXT5Plc6ARGNe8hQlTNA
CxAjDDGf5S+LTBfJZdjK8+h/q74jVfXDk1xFyYP6HdiKhz1RxOTaM8e+5ue+pPXX
GVEzaPCPLoVP25+rn/aU7udI+bhIZzmvz7NwqS7ke/uXQ84TWV72RkvXUIUmgR8w
rsZ2kyidEaf++AzMKvO8QnBBURzoiMNf7jU/m+swTb6p4rwpiBiiDYTPoE+/b/lq
FD/hO5Z0Jfe8wpXEMxeX08GaGawPSFMLQ0yXcAjIzSgWlOU5RhBmnVAdZcEE4vDw
VqBauF68k1320PnCUfT/x6wul4/4IXI4RinYMRkg5yh2HFuK/0WKcp4rEIJz1YfG
6O2xrsi2yfHuAiT6yNFe7kbY58ymnaSTAP23mjE+7EHc9A/FZ7UG+OP/B2dVa1/K
GiWyL11wTjWyHPVQnF6nJttzqAF98Zqi3X155gSLub9Zrf7nvtLytDsoReQZo3MN
t6cVLrLNSVFnIHWWdHC3QTzFnoO0uSIMCXVA6aS1F4CT+I3pc6eLyMrSiGyUYnw2
acazc1rqm6HfA9sUAueMCogV4bum8CItLdDgHLdAtARk3Kf99n7gk76OU7ZSV8v9
3murougZOcd2StgZ6aMlU+JGbsd8tWo417/Gw83sL8a6vfaHPwyDVYMdEpllzYqF
EXpQYt2hKlwxEs7YaFJ5Wl5OpMeEgEqLbzmZWXLNtR+7QmGsmarPb78zvUYnxjQP
WaHDRvVJOStDz0dUjoaQohE9dCsvaNXk6cucKiYxYTU4R5bBCd/RBCG9Xxl4EYTF
dgj8qnreOiF/G+QMmYXVXWwXbCAwIFsdbizHwdiQm43BcdnDfCK4j8kjhKw+4TC+
2AJBRDVM5YceHB2zmQeNUfdJMrTXHG8opAlgJvCh6u6+x/aqPFImWDmtedalmk9z
yHWwplnbtm3hwAM2O+aenl92q9hrlLBClkwv2ljE8l+Elat28Q7twS0ANRzr01hC
VDb0peGL9HJvgtmjVB5dbD+yb4LzM2mFiek9E/AhugasJsSprlV1e5oasATrl/7A
nu2VIsIfXAVsjnvnk7ck5+sdNqNNjjF9CGq+mMCfCLK2M4WopIK3gfmGQGo2JjVN
I4lS1dV4pdLH+f9J7zaxvVTCOaBmEG/CB1HN5TNX6cFVVhiS/sa6Y2YLXhgv1NvH
lrXSazf0CdGT+rxe3y4mtgux7j3iRNXoQKput5/Dw3whfJIY58uivlYcs/R8ASp3
Wc5SPncUd6dyXAO7x4o4QqAJhbGBz3DsWIeh0pY8brwUx055yshm5lMuBbRAoJ0k
hO8Yyr0aoqy5N2iHBZ2JyDMs4dN+zd9cHIoCxgfckFWx4q2gtMDjXgqzmPge3VSI
J/CPqHbWbihr5mXOHXlN5jpWz46inb2o57u+JtUCtL4zKn7bDCEnrT35e71prnUS
iy0ioQPgW3v/+imdC+VUdxFmZsZrbd0eqR+acC3cT+ZkMiS+u3mOV5QajXsbyT3f
DgkGHQgqSis5NEualWcy+zd5MileBddmDAMxFGVYO+rDnNLQ3Omf3e0O3t0hP/fe
NxjkVww0oX8HgtJq4JpNXwK7kSoBL1SbGY/1iqCSRVw/v/93PIgnYohWPc4wOR4d
ELquEmjWL5ocLh4TifgIblqSx3nO6WxvC6U29EeMRbz3eRIy1cX5Ed/erJpVCums
A+qndtXOgAKi3oYtdjpbmGfAq2Ax9rlHKMvb40d6YzP5BFYrR+DluV1MooftFkmn
W8ij28zJ6DE5TfbBxwyNdJaulvrhO97xVlg1rD0rHmftnE9wx7g0g0NHyPat6FeE
huHyjc+errltL9gJsh1lXoEw7Odmi4ABXuwRA8QtgwWyb3ZQPLgDvxn76Iz6UgH7
A/Mak6qpY4RWC/g7BKVHeBC7sXZAP3nknInMEWMhDHMT695y4hEx6qdCVHFWPaCo
rOumaaHeSX/f7Gp4A6t/gm2BQagfTNP2gaC2kVKVw8L2WGHHjL0DK3Fc1jQun+ym
KbULvZBrbex7+79qrJYX7TBu9VNp1ykosIFirky8qRzc74wBJpC4iWtROWMLszAq
HTqzf+N+ineLtkZwW23qTyxRdyPZZtBdReypHyoVaZMyzShy7jrRGMnCsF67Ov+1
sPlPHl/aTRrVOyb9L+UuOcmWavMWJuBW0ED+myr8dNKvLv4uYr5WNcNgo7QPW6tV
Fv+mbJGgzT3ZS5Vk86uJyXD+2U/M2hlyf55EjLWLWIgr+xDsoZ5oZ4tn11SuJ5G0
coamqpAnxziTaqhKYQT/zJW6WeRPz9JagKY2LecQA6D0lkwXEngbLD+3wEv3ZINs
pR1PFs+iuLy1dDHDxECj5qwwDLBc1FhLv8Z7il1v4Vwuu31sR6jzziZO9IRxr+dm
8Ai3+3TuVBbPPiflkke/w/V+mNDA+9zbjgniZujoWj3BOBG4sbVZ7oU+y8yf0pwi
s0fEHuRyN3TrAI+BNV1vDl+sFr5FblkQn5gMtIcLZh++LWLOP9E1gZW727b7Z58L
pztNFr1rCpWZYpOf/Tnc/ashafBg+W8BXB4H4+mQgXRYjq6SjnvAa+9M358EHLCu
mbXQRdmzTf6ERC4Rg3PhGnjODHvTfNpjVxeR46QbiVZ437OBfOXOwfGkK4X+Q/Il
aYRfDnUZs+DGzabtUvKIWvwhk5SlQioYdGmWSFycZ4Whhbm0H0vOha37I0KCXONB
fIgtvuieCtOUE5b3R2GdrmU7qFimcyU5T7jQrFcGrDy4651/Exfnny1gEEdX6vQW
f4erqwdLe+TEk8ex31q9gN2qbECX91VlPJWlukIa6VxuXIdwT5xbb2P9sGymWIQN
mrMfg4pUYTjFA2NBgXoh4FC29iq3IGSBU7Qk+vjGXCWvvxXwm9AXKhY6X8oDPks6
e+B8SmbYFhktQJfX1+s1qw11LNUBgrjyM1FvUAwYnoG2ENlf7nfPq8TuiQBKEycZ
RKCcWuzG+m21WhpYRoFMD73RBOKKJ4zMIQkCDt998RgwRbvcUfRxHJZBEgu1HulQ
WTW5+pRZRkivs7pTVbxU10s0vlrX5VVqmtE0cKs5WpTICpAmY/CadBkg+kUNesBz
2yL9i9e7q+JuPMiGOcn5KXMJNmSWz5rBX/S8n8M7isaBf0RB4aCO61IPYF0Ckfcc
lHmh3yytUQabhDWC8UCMGDUITFP5pdBLQ623+oXHnaLlZhISEplMQpVqewGXKsS6
fObADatyOTFN/6rjrvBoVXVEZE1pjT+CemXFHQg5VsP08BoXuoqRwU3fUzs2GeOE
+4s5zzwT/ffIaHv9idJW4YtUQXEpJ1u2oAteCBoirwgxZass8RCKs2I0XHQuOEFQ
G14y3p2njU983xz3EUiYj9UGyX54ue/lGqWhqpZ3JAjSN/QGscn7eA0Ydvip1rfi
uUEO4yveT8fugb2qDoetfe4vVDUZ/Bak96ZJsYltge286McKFR+iLTj+weQZKUSn
TuKDlsvT6QUnRfAhUJ/pmgXSif4YW5URc5dYm5JBZwSOoi+mogwj6x4Iz/K0pxDl
xGh/5f8hzTSy1e7NaeatMaIpnzcSc8MUKa2cwGwMacZAXFQEHTSCYxaFHgo0QMH2
/HODslOq0byBmiUfkhWfSXIFGwmnhOnU0NyOzOxlVjWK5QdN6OOYIVVYA8r0FZXk
9EHQsobnbNSsDPcEwvoeltYOBcUefLvnygG1Yxe9rPjRNh+l9gRE9WiiDYrWDmoD
rlErGq6Le5r08XAocTtn7AVbfTcI8f8NNN2HipSQ6Mqp+uqyiBys0irBQFPu+Wqq
zLE72IhD7DjCKpN8ZAqGjlcL4/fA7HVEFWAtOEBbzXp86E7q6vn8UFPwLHiM37bI
0btrRC9E3JMxj8Utax6rnpYe32D24dWKgHZiY82Lv7Z30n1OlGmjvftLKIHV37hd
FCsZmCbcJWFywg9vhg9/AH3yokCi9w0iqaVosPglBQ07NuJHQ+HnBRDv42RaJ/bE
mjj7VR8/empI+ZU4JJfh8wG18RDZuR/ckXACizZS2GEAv/GNk1oTCz11zelOHvho
8qsaV/BisYu3IQFwuGtzw2AZF672IVYkpOMgnSQrJbqkXLh11VqCfJ544zCedYKX
SQlqir40t93wXMNrDh1XetpvVVNpVHEitTTjLPAWUNFpyr4zQvXmTQxJmjCUN411
7slbg5Q1ZyUm7xBVMGNebc6lNDjjGJHPHznADQxV4PeH8o+t3wbWsA21rSWhAN+K
7SixixubGPFvMDACX3ieXru1JNKGAHN4sHJZgig7v0G+SXVhSzdV6HFOpYSex0pF
ehnTsJoJSaNaanIEMYh1XzHEmIoPZIGaKmvk4cl7R9ZWGRKUCjfGvBF4EKG5BSEN
gm7kIT5c6YeMM70Ni51cun/JAbI5/b5k3uJHdc8ZWC6RScfNVAc+SEE1QwKJmSjU
F4LvOy0BmJ8ined6cC/rPIak1SSCpWO/ljQyIum0Xptx47HagLsSBAEGmffiZmKG
3WgIjAtyLEs0rZNokbDHXY1heBp9t6a3iJiqQlnM3SzzgsfpHo4FGAqpetjLQS53
XG8W2GWTEIPAefdr9C/Fb1iFIvDSdKnUJHSCpUtGU8Z51TYgb7wezDDed0g1URhW
OLN4aIJVsDwCQBvNsvKfctn37CZqD1z9xce5h2xoiwOIL1t8pOGyct7aNG3XufED
YuUCJic150aKV+J78Caze+yOPpoavkPO9TwyigrNyvGKoMUL6HyoE/b/LDru/7WZ
lVcQKUs8Y1J6019PY1HaXsBwuwa6hEIZAOq1P0y2vfLfsRlb5ucBHxLdoP89cBdy
9dtWvikGpB/4b1vd/eddwkPv/D4ysHiewcoDnn2oPvfBIO9khPzRk6yuSFQ02QbV
4Ac6TZrSKlsNZhMFbUX8B2O30WGxpruhhVxIl5n/LwzCde4awa7YzAGYV+UO/tfM
ZXf3NPb1Z4amboikRV/yZACf1+wWirVSdQK8doNS4ZZaL2+7l8wZgYTdnPDAqW8W
kH6DzI+f3a7D2WCAuL6AD3844SyLnr+vkvCE/PMQRSIcqHdp+JJiUKyFvPQOF2IA
tGyjlkTQvUmjaN2yaFb4YxSCNZ+QrFc59UnMFh7YkNjYfs40q/ku9Z+uPFaCftQ5
g979HM5fjzzS2fUH5F1rjpO9T4BpTdVE7stF1LAZJv0nNgqCpuSEiusKHGmxc9zE
wBZuefzHtuIadAYlQaW1dH1rgDT1ArQ5nZhxp3m1toHSshr28HcYr8dRED/0GA/8
2iI/xk2ybI4FwAjDov24QFXDvPqlLTUFJpMuPZwFSWo47OYmmpFsxdnduQawe7gr
+NCL9EXUoOL1J10WS0rzHaeJ7TA7So5wauOeeTvyB3kYU7V0aMKma1LLnjfrxjyS
9i5oiM6a8VQtvRstfJC1iRnBhu+kqHthA1LF4syOGRi/x84TTl8Wxr0s/bQmcFjG
cO9oFifM3B9wSpQBYsvsQLSoZZ4uWdvGa6cWvu11d/wOkkEKor+sVfWzsVIDXc7T
8w51X7miuij2+2HRMJD+2fAvu9buyU9Yi4Qx7Rlg6I+uwyM7LSi9jcp6isDTcckO
fvs+nAKTqxDpOuaSC99UwRLyRoDLgY2bdZDgXGHR/xtwQ/lpAuAn1cJgor5eKocv
9af9EGrC7519YnyEcaTo0shwMn8IZ6Ofe+ezDm2Zh5/GBj25Drk9lkvlb5ZAhZav
cZd+b5OtFSJP4hfKhicwGoovI43wRM24n2YJKBv6XFkt86d8LqT1UKELF/KV3lPj
CVCviyH2ZhtIvMjElhL++wVQvPEkfJ1AY8Wvlc1NfEvrhSFb1N7H8a1rgrlS41Lv
2zHLeAoOhqGy9UdnXkXevYhxgDgXgUoe3CWL/fFvXwoKvdx3tayDijP6M6anhKhG
2dARNEXarFWVuU1TuqbuYYClvPPAXckhNvijx/oLrASf3z9mzgNLkR1qakPpNVoF
T9DsdkTygbQR3iFeqW6Fk7OmduK/DENOPO6giE066cRRkePpxXRCNFYF9McX7S0x
FwsdHB/TTb9G/E3bpzo+67W2cqcXsHeyTuw1VRIgbZoNSFk6dAk/pUzqT3sCp6Ot
EoUu96BmTwdaINx0Y7KfUN1LkyddQkDMpflR9Nae2JWYt7TTtDWFQzt/GWWWnGge
vE5ozd1iCX8wm2U+Uw8NAW88Od8pcsUxVZ0RXGSqKqpZDuoMBNSQZjixkpC6jkFT
DM5CJCyO9K3ER59D8rp8xPntaeQkhQ1FrgxtKdC0jlEmafzWjldJtPw0q9CkU0pA
72tWlNWOEjkzaJcd89CTLvcwa+WjDX33izpDaLxX3Wbf+ohqwMrnFhqWcbx4kFFO
aTVOUYJD8JiucaqEeLoP9LGLOV8x1PyJOr7GMtbfakYH8mEvGp46IXqIW8rRJaaM
WfsmBWO0dSRAjPeHRIVVLrv5ujbpeqQmbUxUyXhhDwefJbZPefx3ALQGABnT5Cdj
1p+tv+fxE2qTtGe6M/GRKfCZ9WBnr0us45byvCBVAoECljv8K+bbmRzHy6mHJOiF
A3Pp60y5pJqJCdnzwiTcOo30LxuiRPmWWG+/NM9sePuE7GV54/D7rfwTTl+/cgp0
bdMYYouuWSRx81onrMmix+ulAvXt/VQAbQ33QSgD2UD2sR7bU0KO4ebZCZQ+DxnJ
e9EaF0p+fV1N78i8IlcBBZJUHVSGRRRVRSRNub2hYW6TAbWklOYRHTZTiku4xzgo
nXAKjGT0vr2gUUNB/dl5858sl78SXofKVSPSLKqdCnC3vxGhdMBA+ooJwJmp+upn
x/Bn5j+2djSDbSL1i3ISOZcWjKpidw9Xcl7ibHnUtxjXZgjunL81KxUB+/1Wq4g6
1VsIkYcHzbPmRB+vulxB5j46Az0x3DxP0YrcN7o81SkLZGvfwyEs0uxfbEr7Xwgz
OkEbBrF0SBeONh6JbAk+h2YlwBX0wAJkwxqXA7DaPoe9kdcMQSdk0b5rjPa+na2r
ThlEjgatUBgf5BC/ghSXPqqpC4fmFilPiV3rUygYH5CUzQ0XfSY+uthR+NSPr1tH
hYZ0YpWgF5uvqxJPlAWEngxrVhqr2dFPOAtzT86WoDc1Z5mzRs4AOqeZTysdycA7
/Ru77bHDERjC4806IO627r8niKOMtm4vKvQoJ/PXtb+227dCCqKEgN+y8/ygwppL
qh9LzxsWUwmNOMd7UweteTnDKagR5UW4DZiBmDNrpTysJM0b5dnlU9z8BwjYd8p1
lqxZ7chvHwZ7QYRsEV975z/FS2GHlYNIMV9X5s2mFxmQYbRl7A8LXC0GoxiFjHq0
x4qfzSasZVTGJi3xne8byB6O/tneQwchqNbIrHiqN2PkqFLSbxdBbSaPTZUl1L3e
6Ch5bjNo+/F6yWqLsaHfJBqt9nkRmzrMaNKIymTT2oqkoNHwyDrI7NoHDDRWNKkb
f7ClbVDJH87Iw/aHFv3uYIKwvAbUs00sUHSg7SaFKO0vx5s9aczs0Vk5WqvGHoPk
ecJWGZzuGxeKWInrELILKCjcF/aDg5MM1DDaXQfE4B/YEwSCcwIMe3N2crInZZwM
I6OwHgnowDX0KtwZkcn72xcvGhwGbilA70pLO4N/oZ8YV9zY6xoZLCnmqm9/tVSQ
69SWJWlfziuwpTwshekyromZSOSR287rSqN0dny3aM/j+anU8/PaRU+AGvxlH4f/
T4KLkVjbm7swKlfGSNbVIWNClINPcUWimyuqiHxbnn3MiBMebF56TygTSVhrO9p9
rjhY1pOx4Z6cUD7YHwFUENB8kvmO/O4sGNQ5vLWIyJdkjAOEOaj5NXj1q6U2ZzXx
yhR128K5VXhY22BF5EpFO4vGLJSPjaEEeTpBJbIrTFiHcp8O9/aj07Q0QjjDfEjd
/W6OMYx3IU19+cnMOR7admkej3ADAIoYrPivnLEOPocZua3+QKwIoH7NKf4TCIcU
M9uTqmowaJDwpc1mJ2NIQb2mlQLu70R2D5phjxn/GYuuNOzobVRHLTyujiPWSnS1
KUYWlnfTDWJNObxNp6wm3gosxzMZslCZNbaUAQc3njcxSHtxVT1+9CKktEnoRPhc
Co0U8WT6gLy24YsMoRrc2OJ0iTFz97ALedWV1gTO+mMLN3W5eL9YkYXGFC3Bi6+k
onAb8kdaZK7FnZFLsLMWAs2BFr1kNN23lPk4xfWp0k8QDVAPJArreuv21RJcgGEh
Ahy7vUbnzY3a8kquT3X9lA0RkHhe5dnwK05SJPNDKjtzD08uPWWmqsU9Xx/ijdjA
unWOB3yh9ZaXE/7ZhW9hOEBKEiZsFRILjraFLvo5YuR/66Tw9XqVt0RahCplVAAU
7ylnwKFVtVzQPA9EwPfWpg3NoFvCi7fNPKQGsfDUJbwWVPZrm/TVtvXUnSw9FpFI
HRtmVcq13x2TL/rhKgNYHAqxy4jrdEZXrNGQXPRm+j+CTEz2uBQ84Q599J7Q3470
3IuuT5agf2XeC9hs7R6dgrjUrMndY8AlsXeTXOyxc8qm/UWJNsHjLDme3hUyJfZr
/QF0H9iW4cKnGFxiRuHA0lCe9zFOddlXRa0PT/L2aWuyksxFqypsc4/qOcnnfWKE
mO7lJq3LAijzyc9SMpPKq4bv3WrQPZ8WkPSMCynTFfEs6biUntwP4+q2w3B5MdMO
praR6NBg4r1a0VdpHdiH2/4b/rS2xsaHC7J6Yipft0zQvLgfLM0HyWI9yziezltA
4z5d02u2L5CxhVk1LXoGKDIjdBW8mbOsq0cqkrHKAXxloAg2Z8gZiZK7QnocRskH
HWWgbsTESC6waSu1dMam976uJf+YSSdeGU/gafyGqouwFso4lo6q0ithTyyahtIq
YP1hbH9+4ye5Y9dUisOwa5ClgeRrs4+cjByeU0tQeq7J1ylnW6ddZcsJSP0w4P1y
IdlX3U14vzb6uUwv2PiCp0pZj9eEbLcMYoS+Fk2z9/2uF6MPt0inC5hqV96Dur+y
28lu/YReYgAXO3ZOWaTSrg3gQfXO6pItdJQJ4HC8i0UGWL/V5IukRnNI1b1xOYZU
c/N+EDcetUX/oep6ADQtcVC0S3b9A9EaMjSihsLvKxMwbajP0jxRcWBJAg6hFtc2
VfiDWXM4mvRC7XIhtgzEf3kB8PDYXtlDqWWe3nr1w+OOKsCcqYhnReRLqKUCll+R
4IPTUBCy96AX5cH6wZ65VmqffIH2mWVpPg9fMzU6HlJdxTAaQPYeOuRe0bCX/OCK
RVf9B5dAITRio4KAgcdIBsSOjIL7pTaUO94nzilNnHkq+qqY4ymm+QY20o4oe1Ug
Tn3dtj00AA2DJvRheuHvRz7Rvoksx+QRHnur02UZW+mFiz/G2RZUJwMhojXXaAXQ
5j5dcMNBUGHfPh1L4Lcx3jGzXoi1mvsPuTnMF9sjUUBzbV3m6vkoJ+8LSfOoHHjb
nmG9t+Bzss10Kqov5iJZotjsF6o0BQnHpr/8IQPCStSqBCu08JCg7xm4YsUWUOF1
Su2zIpmURRHZnWA7BHB8Eua74b/v3zdg6sMvyUB8JTffSAmiK1YTdnGnFUfll14u
dk/NF1AeNbpQReo+ejJZFWiEVE33Js5oyPTmbwmXFcC8t5W528F5JdKpWXN715La
uTOSiyVsbDG6YhvII63xe4ga2yj55R38z/YF9mIhLu9nt/unK5o9yTSx7rLLQ2zc
9uHrMbss49rbJwgKjflP8wHCpOJCEcWEO7lwN/KT10XZUZNOCUuktjewqzdgsC5u
/kw6RNsdPb5ZPaHoQzqndcwIxEcrn5CQKRv4I2NLalFqMb2jBgHIfWkePHAsHo7Q
cDmco7S0SeQx/5OEKivDIhdIGbi1bx64I6Do3QnpgxlTehEccHojiZjZMi+/rjzC
hZKHvxdtQrC8KlQy/bNGRsGCgPSKGMU/bW8vuDyDx1IyOKjGs9qUeUWZtqOScycp
I9Hw1Z9SNGev8QCuSAjKSOapOla22NCu5q0dpQQjBg+f+Pq/FVvtgmISeopPNHXG
wJ27+R5LR2tSNYxSS/XGDT5WXiGeMjkM9vCqKbbBYHnvC9nO7yvP5esFX0nxzLKk
rXdItgFu/veGucH0pJ/VBfsQDzjMpyxv6IAON8wc60wjazGsvS4kwUcNB/NCOBEn
dzw7T5jNRz7wZbTW2zji62Eh33LM/ADObRjV0kZBRwdyIYkFeN9ywpHz6TgGIKjR
MVrlMFx60kzeDgsILkFw5vCDOyo+iz8tOYenhAKB7BDD2HWhgUX0qQ/+l4Z1g5dO
i9MIOVd9aTu7C5s7widr7i8r6qinpzSSk1fB63WDQc3TLasfLRY/UPl3LJ9pLU8Y
RwoXo4X2ggpA8EfoInG91tzJKPtzqlWPyM9bbwW3C0VQM48kv1hklTdXhsIOpvZX
qy0CcxRwF7RzVN6cOiJi183qt82tweKWTAyZ+i7Cc7J/fb9uWjCiE07wCR3IKRAO
jOm6JTnGvvvn/itE2l9sUKyl6nc6DCcLmUS6p/Tf6l6hoMkYZieljOjMDzh6Cv8E
wKF+3U8ejHnKuV4TCRkSEUj5xMjfRzaCbNy78q+IWnJZwwGENmRQ9DCIgxsy1Zt/
aHdruGWSpnnvoff5fccWKrXZO2we/WAGNNWZhPNm3PoGJErG2UglGHYTa6byCQ2x
bs8oJyb1gQf7APrK7AeUK4cpQluX0xsXOgba8TuLwwSH6ot/LNJtIrlY2q6kToTd
SGSTklFIsxh9tM5Gaxq6pwVGC1QkzuMe9kuaG9Jfm/qESI2SjMNHEHQ2a0jfpx/P
/cM11HDiXKpuPIFBaANSMJIVRhMH0bprCDmmUyrRy0tTPjwZWKXlFnBX1L4mVEIU
UDdvRuvWYt1FM2Tf0+bBO08BXIki4dBxvLBNGtHES4N6hZB8sAiCrnshhFteR5lN
LbG0xxm3Mz8JaBx53oq7wwZX0PaZOHHqH0wCCf0rTdyqWomJuxpLRy6FrbTV7lDy
MAYvzDlAgmmvPqtZfXd5agr7f92Cfq0YBZlR/TQIqsq5V/eg7tSrf0yX5t48K000
0VDKDlrEwTiVCV9O5vTDV3gJ4/QUgt3YIo2eUUBXvAjrBwSFXmoM5bySHZCSXcmr
r70VvjriYHtaPuaEur3xWmAAHxISodm0Dzf8ltv4OIc5IafjIbylLi6S6tm+g/g4
4073k3JUqfcDp/20ffKHXxF2IOG4x9TKB/Jg86LpAbZZsM2eahACoWgm6QpPh1A1
wYWCkhHZkoAxnEvphTX1ywFi2C20252wXZ/umBHVF1h8kNRcLo0P3+MazOLn7ufC
+bwAY48aJuzfzxy23Cn/8TV63RGPXWj1Muc/9HYe8KlDIUAilM5J5yGRcs+ONzss
fsjZJRm3AV3eYrE5DTsQ1LV+r5EEr58Z4sh5GOLP3oey69WNIm+e5cda/1dUOAJ7
NYZFy634l1deVVuXHsEZd0FwL/eySwd/X1USyQwtxMBRv+SLH884IqlOW4ObpKea
8dzBP4K5jrtkSr4VK2RZl/cZGXEXVGKN8IQeVcSNFu3abUA6KXYSRrECIgaI77EF
pZme2JzI7L7ISZPNE5V9Z977EY2R15TIUUuvnOj+GTKu4yie0aNVqqLKZLXtPPh/
gvnJmOOn/c28jKJD/eKU5kfvcoyYgPeG6Ug0Kh1xUK/787BWKHqCpKxjf40bftkK
fzzHlGgdeUlXWYuEdxNwtAHSAh8aoSeTiLNWzoTGYABAZlUoEG5ha6PheMGHBtnh
tQlG2a7FYcEPBxIEuUh65h4inmOo4AEL7D9+jVCXT+ghi7cJn7MpJ2xA1S0jiqfw
U8UvfJZ/gAJmAX3qGpnFUrNqbtSuiJge/O+MkuNC3sQmVbPNBSU2qChwLTMFBDUb
hTLAChRjaRslPSyJ6wRVRw0xcFKj7UFXDV8XZbHLoP8qmrsk2SVwq3+1/K50qtQb
9DvbGKmxX/FgUjrx44/7Jz893DTYxfDX7VlzAW5lIUB9PFDMrQm1Eqsw3ViG0HoP
VhPxLTpYBdjIQrMmrTsRETcpv6dPCY94OAgHnyufQVJZ/wbzcjWWFRz0QQS8WGr9
BXIUNIie3rUxgfH/IGk8PIyGoqshT9HzIPS7mKcstcMJzrQoldyVe1EESCgZDTAG
hiWWGGu0biAiuxSgaoRCkDnlWdfwsGYvdZo2EoriVXN35mN9VWODHh4eILuOy/Rk
fEa95ghqbmHXGHc+GP0MdR5b6ZuU2FWSVqeRFDRZ1KUBz7FFQAjcZjeQKnXkbi0J
1NMfjx8Y2ggtLkaDWjzYEnDj2UoxKIq+JwKD4t3aooRNrNt28J0/cwhCpi80rq1q
6lMkYnmyQJvjgFeamG5V4RU35sH54zdJCwE632CDSdA/XNbfxcr7IDUhT69ZMJVa
cqsHA2RqtdYPrCu/+zAgS2k4utmvl10GO2JjaMES36jMz/I+I/An0LbO1JwyQFIP
9n2husHeMB4TXBPsFPk9XJ7/vH+iHVcprJA/KUKKIUO5/2MT0RwasC8OupbdZFIf
LJr5Tfhn7J9kjABjGJe596Xy07eH+weniNTmv0+F5CAJvcg39PrCAj+ICH/e4dxQ
ezMUm+68jY6CbM1819ALeJODZ9kAs5H+zs/G/yniOQpdcCfrt9UiPIldUQymTeJw
CcVYMygGZ3oJO1TlkdVxc3iczmupVykffP+03pHSKMXzIk41pxqt3Nwz/OTqtIo/
wYRBcnaZO0ZT/sQ99bvgxvEmER3La3X2r9Ha+MEyDIpOXjMo0JBXrN8j2vVl4NuR
DfBUZqXtAYXPtRPoeOwf72nUgn6erN04Sy+yFR+ThPk+LNKEIU2sMb/SF9DQYQIH
7Hwuh7VjHCXjUgghX66vhuZtF10DDXl0WC0Sex0K2DHj2dnJpWHjXSf0lYmRpswy
sFWnezuURpIswvGQ0lXkjv9N4QeTGAfxbqPPd7LdPZX8Zog7Mxd0umInsmt0a4rw
1jq28RlJgNk9Evt/u7iEizOxvDNU+tqtpDJmKtm8zXMfp/3uvd5uyiCKViGLcIYQ
/XejJh6qR9TnHfQ5aDOYXW9uhostxPUS92ARLt5tJ6shCcd7Dt+SejAX+vMLYcvJ
v9eVrrOUOK/3GLd/ZE/XHud6b+owarPwkO4N8ptE7MI7XaV7KHMJZFUpvZPauMho
1L/a7civyiRqqv5HYVVNYapwV+wpNRtZh0nJbFBVYa7hcjCy9jIdsz+WbReGJWhL
jsRrJwCkl7iB2bPMh5I4vX0/zU9T53wqXaaXaP7Il3x1kzh4/BQ2Xb/aGqd+I5Un
bh1xxUZK7w2vz2VFYjADq4ZkaIaVQfR9r38sy4CdIcls5P/oGQGE52nks3omLbdw
T5j6oir2V5lScovKqW+qztsYmg0+rW+70Rm32iBrSqBcR5qJtTNImh2FkwTdJ+7/
rFn3Zi76N84blm6Ia/dGpc9PnQvYUU9Egg525LsOC3S1ZrI6EkDad6FaSZmxk0ck
qVVUja3BqY3HL0b0T6oiFH5FAULUUzhlBa5n2c+jugDLzjeTtQjvK0pG1ZRuP9NM
JVJTMtt+k+gFDmrcZ+nqXiBgComi+7jQQGwhB8tZ/GnIGHn/tGR1ujdpODK+JXwI
ByLuR5UQ40hH74Rqu3lpgnll3bZu/gTn30QZC1CYpPf/1mWrz1zJg16E39BFmYNr
imB3krnCKSlmRHZBOxxVXXSCs7xommEI3AzZUXmqAP0Oa6PkEvm4X2Dgsi6zj52Z
1JZ/7xSVMp8BqvbmeuKcp//srttTHUHT7WJW9DLNMat2NkE+zcyyEtXpnbsNUBlS
l06dbB3kz3fXZL1IUmZNaqQKDqt/ZYL2/yc0q6Lu8o9iT1HBe3qdpP/kvFem1Wsj
ohsnmwcnFYyE1b+MaUUZuwBfIQf5PJsxfHusLTjmAN1Qjkyp+VJa4LqQg1ALnvIV
PG2S/W65PdUz/+R7QhVtL9fc1r7qa73fgRFtgmdBA2sITkHZxW+vZlSc33qvRO6P
3Je9AmgUlQjkXeQYDo16uZ8BnphmHjwAtbLUOfhW0nmV2wVFuZ6lII3aBC1KFAIY
n0TA/t9wyBCpm4WAaMVeq0KvWyH+Ehm8ryPcHK0Qyn30J1aPgEe+FMU6YVejmQL4
f9Ur7cDI3IuMNBFHeL9ysG5bmrWOJCa7EMqcCTHUtfzBSTOkI4hHfbVju5LclCK8
wbpnZqlQjGRavNwD4rtQuHC1L4wvzB3B3SvDNiohy1bnQ7jgeeQZVt7DlqZ3QMKS
CVpXJqW9sDXgPJLS+1gwvE973FU50/2PWXlVvsgbJRBQUnAzph6sT47bZd4HG9le
De7XeXBS4tfJu6lG2hwe63bIWh8MK68zA5yyHvTQii9a2d7yyBaJk49Ztquxsnpf
FZwKxL4OsuKUJ1IraxjDlRZHAqi2UhETywys5ri5GTmxj5qeqzKwFPAduE83kicf
0RBlvK012GYNUH2jEB8FosUd4N14FsI4f7ZSFNX8A9AjNNmhHqtYtEJgSQ+/5mwl
4UZ6ckIT9Zpt9izlWhR916X5IqBtWl90frTu8/W00SDvWwJGzvncYHIPKi7WySVf
LegL7QGge/xh1ggdAamJmwXpNmsDBLL9zm6nSPt3tKyY2hUkB1037IQkCM6IoBSU
UgJE9ARrBEu7Xd7u4fpO4iOSkfRg40aCh4N3MXSFA8h0ZGXjhDsSuxF/Ff+2XlPC
vPV5A4jrKPpEK03OD7Ax9I3qPaQbwJbFPFQv3lRylkzGSIH6XbJXrHeyBVo+jTlt
ar0McL9NW/rLwQsokTtTnEDCDRp+m2qQBTFvZ9HHlmtePJVWtLU3Fc1e6hksBN6M
4MXQVcfxt5gBmeiFlnMexS71jL9nFHskHce7xaOvBDa27GAwCscf4fQYdCFbXjGZ
XQDxpJpgjkApLvdMANkLV4K7HbvP8lgvU9EHpJYnxV0NXPxdunJlbknGON6l90YN
8CCCKc79wLavD7/FRxH7tyhejy0P0zdAZYtToUr+LDDQH9fDwyvyFGnD2Mch/It9
IWqZdrYdeF0f2zH7mokTJ7jNooLCxzoei9YLrP4zEWOgofMM+yhf3uH4Im01mEa+
iWmOtTYxTHwlKiTAiKudqo/JmNO5lW1bqukDEWlJnpdgmlYkW1+/FAuzyVR1Lsf3
38U3yFjeWfI2YHvtHxvWvO/wQGSZgW3ZdA1Khntxq7nZ69fnrMF+QoD0rLp7EnM3
N04uMgMQWdkjB0217YU99SP8H/qcuQg8FMs5mjEmcE+dIrCQK4cf8qOuzBGsTV67
FzGiAatu0ZdegopPYlN4mAtIuLjMOeoj2yej5P3A+ibvgS8rXzz3O7yiFHfKT6zF
FZfAIIMZAw4fm6k1mHqJyF4R3GCyAma5d98H2EOsF1+/7TRCz3RAv5qB6rd0P1LU
f14sPeoHAcEilbk45ifiXrCaz+hw3DcnQZeiwR7EeHBVEAw7SuT6ZykqLmNmFBsk
Ah98+lK9z2oLQrjnNTKPNjiopTaUrfb3WN1c+OWUArdYIegD0FbEiRcidPsQbB5v
hJn621macdj7iMQWASZ2xWspPFwisblpzpMwOxHZdQ6UYJxcchWMpLxeco87Wq1J
rjIOyp0+C/gve3Lqn1z/LWIg4BioFVXNFtcUsnnxFJC8+44gpp7P0uBfBecSRkFb
weCKuFnWhaJkkHU6EKc05s00g2stSdGTO1lj9ggxWvd9dSQ+lybdBmMXJ6j6uUQC
Io7v02xOkvb62Sn5o6BfTN0ct6lmMY1tC4I0Vk25ERGZowIPA6WjSbj/XNYRsff/
4NjixXS6JrdyuZmw2RhThzfSFkjwCvrPYSDamXltWY/JMJcEAOfvb89YMAW0lguv
crJDcir96OuQFyWswrZppOA6GhxMIo7FiOrOgnH9yJM+zSwLiB25Vu//WxSz1XiQ
kbxzAO8IZSOWd8oMVNOquRAWNX6itxNJOBsoqCLUygwBldeXagDHFzB1dddVeK7q
yeOR6iqaKlH3Rdn2CAvaQtm4uc3PJ2f1mtUlXL+oBgXLH2JppcBIPJGclfs33I3M
N5MRxN75tNogd73HdZZdQXBheP8LaARTb0+w1BwJOdlwJo3TTF+0RIpcnkL7AOOJ
GpWRgZPpF5xEEpdxuYfEvCN5uFx+OHtX4g+bIro5x5qUaiLj4UIxX4n8ysP4jaNO
Me10dy3Lz4877qI1oX/X25LIPzRDShuEnkWbRHnwId108C18uJsafASu2jyO+PNH
VEM8DieGc6dLpGcq460/ohVEnJyYpJhd9NBPsyq8tlY5KmueGV3V6D04z8zIj9MJ
hzrGmMAGTaEkKMf6RVkaLL3z+NSXM9n+XqMPvi1hJu1i0kBwV8rRJSDZRaPS0ON5
BUkePac2MbBIYwy+lDWToDcKHsIfTfqosWa3clQ/VzxZhhHBrGeKrqxDOVTAWZnH
TBiZz6Mri3cYhj/ceTer03byFmg3X1uNstjFG17GI7638k1VK/RvsIOezmh4h+bV
y0lYPloq5vxe00cSddxVrMwg54BX9tsBkPeG/Q+iqUaoHB2H10PiJIluRDR/oyp8
U1zJj+jR8uTEbFxGQDcINraOFHUd1Uk+p6XaqUxHKWZpi2aTqDgauNm6BGKAwT8A
WH1HBAYWTIZ9Cp9r+TEV6XrNq8mc7pryrdVEjdPj8VEYWOT4CTLDuDq2DAQzziN3
mFs1Brb7eCU5gih30p6zyWKb8kswS3b4ogdZhoK8H2HJW2ebxQFK2obcp5rGlCl4
jDoIJUv4AkmOka1O6vs/WNzV9GVRIuJhmn1FmGsUbYoK4m+LuKl2Gurs936TEAZr
0TNLb2ehOsaPB2nBWLxfngyaRdw8wPqYeY221MSPCtDBu4NDjUae8UaJ+jhwzvKr
BmuvTXgNIYLDSiApiDyb+AK0yQoRdNlKaqtm3K6QOqeVH8jF0Igmu2g+hURt6xsh
Hm4fx74tEZQr+sgLeCbyIp45rGppFZ42KKW7CmcpuGTsmZ0DenvE42LeYUi8c/mu
2gRLlMWvogtENmNeGFPwRxGaT2hisbqp+XjEdmrzj4xptBW3YvJ0spCjNdWtGg4v
QfPDy5jSp6NRYRFJ3YVHlgqgCfxJfF/W1hrrZhXORRL2tHI31Q/DvnPa77S/MWfO
e8lKNiIPnJo2xXxAqdvFFwg6F5+iufyh78EtZNlgizyp4hULB1nFLcbLcokIFSz5
1PZ/LTLvTyH/BMWWNcBdXymtYQta3rEQ6vtIcXDvuiYbm7GHq+XSwDe/Y6nproqp
ZggR5AFpoZX4xMB/fA0PlHfahhpZI3qeA+O8DE8iCJWjUgizlVGS5BGj4VAF0xo0
gPVCriwOjxG33cNYxOXW+nJDoHy+TDPZmOA3uwCnjyRVyK6zbu37Yh1NRphcbCUQ
l7vlP+lR5WhHuc+sgzKLcaTu1nzR0txrB/Pg/1d9EQRTsi/nFdgM6Eg76KFmGDdZ
pnodN3VUWMbcarg5tjO7EmSlgElTDaoz+EmmO2MY6x1XQ/Va9V6uSr7e78e+x4cS
LsrlVilgfiWu45GCb9MUeVCRNz8u8VQyzvf4xQgM3wKHNz9iu/EMQ9oT2gOlX66V
vTze6wWfHFT8yYs+Ocj9N3OXlG8ZvHJSSRhrhZMTsf10W/IzJvuc7x97cuWQSYIS
lBNF0amBQ6+A4Rwsl4KHdamZbMiEH/IZZeN5qPD1SI6Yk1Xbt7/WmhoaQceavj+x
M93IWjMfXulROY/tmSO99ul3t6j99YkbKHQ114/H0c/pQxhK9bdR2JDr9jSNrwPP
I6a1/xyBgTz3Ocw5Ky99aiWaPPjKfvcWMzuiJJyiXnwicpIi+GP1gdXpLEFmJ/C+
dL+OQf79dwcw7Pi6L0aUhQvSUwXyt9MvsQgG/PYOLxxatbvWtxmHuNWaHDS4xgQD
S/lgbGLeW4t6JOKfclW1JDw3vrTWPxDrdbUQnNPxzeAwqF6TL/oazTRBNpCtn65I
hqXofv5Fz/Xd/flKW8P9nOiJSP1FE8FpzywAlO7iV1/vMBNsQf09XzfK1Cjh23aG
1FA0OCzNQWbbXf6tT2Y3Yrx3ayExoI19WsIW5pY0eHR59uRS0aCVCEhusVu6fmqo
d9s7/6KH8I6NMiqFbGQF9N3RYV/ZHPuu6TdsLcyuB4NrfpdFsqWGKZ1bjFfCeTad
ABVcIEThUsBif2Gmiri+dzVa9ms0qwCbxWnHBPZpb87ApKuSwtCE8V7ZJOAPF4hI
JTemL+po5JZBC9i90tldkxP82m10oX2XsEWjaN2Gx7q0noYInsvcc/nnV7BhqSUg
IpG1XZg0Xv3YwxyB7ayFYvhSJdbavPlDLSLy0anbrPzofTmBDnY1haQsUk4tY4ZL
dlsBI8G5iO/YsFioyLRwED4l1wZo3eCDsfbSH+QjSh06YVSxLUDqFhSOlejccpzO
L+4ksN+ARbA4ARg3XZ8ogoyjiCEZLQ9N1QrFLVnWkvetbokLNynhJiWv9AIJRVwu
DEVxJA7fC3Zpsq68U/1yfcfKL3WeiWJAOjoTtm4Co0lBrjKtjhN7RhTLdhUjCE0U
uU2EdrCg3nSFyWEYcgAD2skOixVUsntpQl3gMyUDoJ+xSvEyXZmLkM6ME24JqhEY
+uQAHljl9sGpMlY6POPnpgVye58zHYUBHtcEO0EEsyiv8BPdkpzHwu9maBAqCMoJ
XSTRrIWOKwwhxMUUrZcBb+dbWh0/pxiNoW+sDRNIloTqYbGmQghUYejRVE+zqIXu
gz+/YJIfDNQafnH6c6HkpGENRZTGWteaBPKBPXWdBY7QUubmbx+8XvOlaF1X99/k
ISZrIk9Iof6YuAVaCB6kF2IwGVhOySpBQHCsYx4bONJzuWxvI5bAHfIStd8IuO9N
828RqbXOxkXtrxYQ0RbN668jpT1S3tIpCFEWSDcJJW+zy2yPgfxC0MuGNvWlFe8g
u/kKQXUAqt8CkhaHMspMeVS4LLkY1AiQuT0601ByiYSgWp+xiEv7GWpWQPTBH3wc
+DnBu4ofwn4Qgmx0zxWK/wLfeYc54Ncc83EybWSvF/WpcNt2ZqmAKYqZxPi6V13G
n0WQFasSJC8EHFWQRkefSy+lJaFh/E3V1gu4uOqjdsLh339VsY/XepshhN74/ENH
ECFKGnAGPSk5uAOpmlrzX8W6i5+Mpt05THmVHGw0y+ot2s1UIsC7ABW/92IvayEb
K8S8bl+L1yYdgbrinkz7b5rQZi0HO5QxxU14A0u14wO4+DpdEUvclyUfYCpqAgJJ
nskUrKErxUzoEhZvZ1l68xZ0JdotD+/C2NJi7R6W7bIb72qOMyBBtKB5F3RvbHj/
mj1uhv54VFoi4lqvNtUP2aueB2fsFcxBYigc8EhH4oL3auRVafQt5X7X+6DMa1ds
PWSIfavYxncqEg+FLfsCSmydGJkq1uK2AOr4B6YwaoXafNzosaw+6T5IDKApTgI3
TNo58Ez70x7k7lcL+Bh0KFHyijud1ThErmsW78uNLL7NY8LFsY9gKot3QaIieo1E
ed3ElON7RVCtQqcZ3/0r7sAxeYefpivLXQQOr/6f8RRLFsFjs9vVXp9y4ElEkRKf
bv0K2wHkiAsxA4aKsGFB2fFOcMKvqLYE0E+/eLm4HK4ayCPNOoWeE+F/lNRJWfRu
DEmz2CNrAmJVoI4UwMXSmyEMPlWDEstjfwQm8qGC1SpWrWdYg3jQtSSHNFMWfUiH
uSiQwvlGVuVmmNuW9jIBBEsJ7gMJ0IN5ntRhk8ltztlo3QS8WRkyIAnzZ++MyKZf
dZwRR91aMvFVTb2ue5SEzigUaYd/KWsGpLZLpP/IseuU0NkmFRVG+2IOYZfFTpx3
0r+MrnxNxdc5+xoeywmsQqr531/o2uxn8xdlz94EhkjV6VAF/AAbTsBgRTG7c40k
byPFbk+PDZ32QYYYax1vsDlB399zgim3eFhv1OL81nFta0f9/CbCzLHvW5bLnJIL
SBONTSRZ8CTjSCuA0pLHpnalganZfaRFkkKvJOtscjNkz+4X7tbMvqAqgGA3HJf1
9gl0tqUfLOAFWsdkUhHns+uKSUcXgT8gopo+m0UvkGhiZXrochJPEwN5V8lghYlC
ge1/pw5KiBmWK3EQxUjhckZnjEkZXDATTAWETRDcrTTTaHMRMaRwa1gs7m+kHvTt
OmDnhWg4RnHSVS0eIHTilLYK/FXyfEMQ7O8bYJ8pvXysu3dFMtTVEcGR7GBoM/qY
eCTqjSNWZQxSUUJtZzbT+CLUqFLuRjTGT8joUvWSbr3ixZp//XGh81+t3CSKiFBI
S02YtHywjhFtLwyfgpqv14HoqzxWxCKZmGidmT5maCLTnBGaRkjkO8t7BUnBUVMk
SXMXSwxuMXkY4CagaHHnD2Fkg/5MxVjcTq9eKJc1di13XYvLv6v8OUT64n1zpM5n
pI1IGom6acVugJZ+R1HiFbrtAwAW0N8bEJzFvQHIh9Hma12LnyqWhQpufkBhYBBI
32o1LPpXShc9I7uBYonEyuqNzpxX2iyMUC+egmCOig3+uEQseO4RuI3XO4DnNC5D
LWoHO3L1wHqxoPQKtwt2EJ8saGqn7bvxKwAkswyvMagyBnkK5bRvamRJopQLd17O
2es4lXc9vyX8du8Zr/GzVmadwnlIR0v6/O3F6odGsz3DbApizV8SOIf2Oap9gq66
HN0hT9+dbLA84H1K8Wz7Ol72L8tS3dRW7Uc5KzmN9Yf+3H9TTJHzj0nFfLqmzYIP
/UbUQFwa+luNSPJ2wswTuIiuVzHs6H3r9UKjGg4z+pJrxOEpIz0mvmaO/Q+NZQSU
cC+puJ5ncvbrQoaLwrtut1mMykbSBCMssLoNBuEqzNDtHxtCknSbGxEINWGZAVBj
1oylwj7jV0KOpLwt3A+C86mEJ9IcBb7MK4bVaxFCV1q8PaPqvMTg2slVKz332wo4
PGAHkrAnuJOHyiTCljqEvYhIL4r9NYOKfbKSGunyzz7q9QCbSnhFKgrBXzv4TXSe
FiD63AMlr5duT27/HEJQBK0b3GxV+1qlfucxtrSVssEDfCmQRpONJQcOahn/cdlp
3dUpwsETU571hvC3uZGQuoFj/sdQ9gtVO7TTB6JCtuF6x7tsYZmdxHA+VRulSEJl
LT77ZKNGXrw0QSMI7Qu+aT9HnQ6l/S98G0t0UlU86XK08b1EOHGe9zjsGguxvOWg
QJCsERYdhC+S51/9T/htWY5C5FR/DRgPVRpzLNTqcjHs9bmq2/qlS3QQ4bVcL5NX
iZbt190BSaSFzjKe4Olq0oyDW5UBlGc7F+CrwJlNq7DCsJoA6j0VB+mMnbpvxoDB
aGDnss76Ch6TypdBC/STK2wIvAgaUKdsptABE4UKpdghcARUnjsUblTCSf3vjLnf
iTsStbdGQisjiXuV8mcSTrNNG5kzRu0c/H9fMI1AX0+BXDvJUSpypJ901Y+5eNxF
hcrruDUw/9WmEmb2t5S9WaKMsgMT1HXahF0a/iuVWZpWIrDyC6TlaVT6+xYs6RLE
hIOqXgQQPGn3n9JM3fIi+Tnusn9Ip3c1HplTIDByvatgCqsRCJcPRcS0wnybUTMP
jSfALVI3CjgSB95MovR5pCr7zsaLBBZ1FGr8tdmukbfBOYEb/jUkADD1vIVE0M58
2dT+AavLNnMWNDpNv2vhEjrS+AZQU+kc4NVgI2rdDq/oz9KblCuAj/eHo2PnYuQq
ZftXWJMHcouPXXLyvX1o1vNVcBl1VGq+PHmKoCOyO26lmWrPPhzOiNq1QJvERgl0
Lwvj8SjofNsOcsG4MB4tDewEnAc/7jgkwKMVBBsDX42A59y5o5tuOoQbKVYN0B++
H4mGzGw+EngeV4KWE4HEYcVKgdgFBwisGWMT+hVD3/HvtC45Antuko8wMVLs0kvY
93C1U3Ow5TIk4732Cs40D/QxMaS/iZ/Uy6uwb8UcUVeKVw0Ny3p4Age83M+PhpFZ
tIEc2Be4udVwyz4uOh5gCnAgV53OV6uKB5q58gDM+GR5teHrDNZ9ExMbjoxDXRlg
bwLuWo/zBQk+BpvMdJCPeFul0dqfS92kzYXfydwU1Y4mexb7qbGiFP2RiiS6YfhJ
LylfMubRaXTrJ2kg+Jzvmbi+d8AfloUVE/mUOy3WE61uEbgtEMzoPyb8M/uAlbKZ
P/p0WiJiwQRlP5cLTw2Qw3ibpEX9cnMr4LT+WuP5lj43UHUQw83U2dgZhR7mH54o
l/cTKDDxFHer0cg/y69Lfsv58/UcdiIU6jMRHvSMhDFVn0sik+bLmsPa5gd11MUu
y5oJBlHz8aL6TrZ4kMYqvEVNPbYx5sqKPjKUISnpK3JEWSVVyfUmh6CfXQBkgqOt
TfaYcH6lpl7xA6scfmq9BrIRALw+6i6Dv7mcKK67sJWohFAjmGpFGsJKOWpWcFYl
TaQI67C1nBMDovTIjQkFuf3B9UyeHvWqR1vKKlCcDABl6IAcI6N7zT/ieuCdajCr
7zLAG+Xtz2vBWtjj93mZMUYDQ1aXjZbpzHUd2L7aL96EEDqLzc4nLiEgaKmQHfn/
YNynw2ygPT6TM8au2K6D3h1f21SWhkC6GlJ/v1t8SxHCDnqQ3HiiDQ4Nib5ElYyE
PVe6uong0WW97pl4j/lzPjPak5ugRvBdi0iqt7KhB6AcgXGHZDeF0ios/BZwVtEj
zRInGkKT2XLsikL/wN/Pl2PGWZoy88Fdv8vY7pL/jBTi0EndCLg/hoMEtSX6lHcb
9XhDGdSeAdaHb/xEkiK9KCd8AnGToArGTJ1KMikPvawdRtM7lVhFJXd/wc7BeS+T
1BsCxvX43yP6aG3EJurP94a3DvO0Mp9WyY6XtxCwDyOG7ueKSE/uWjQg41cbrIhp
22yQiYTDxt5DBflHsIrYNKKg+YKTkELItnrXRmXzfvdql62B1Rb7NrwHqaL901lC
vhJQQd+HQN0gphb1MuXgqae2EGP8utwvOYdkiJ35U7X08JmEn4AD8selZspsleZ+
gicR1a6W6swmglbduToLnXjAUfOSoJP/+m9OrnpgxPdNV3JvRJ2aXkKzoPjSCPwU
ij+XOKA2ltQ5jWT1LxtpbPzaKoKFKNtjzQSXdFCvS0XciGvacslT1gSMdqHsNEK3
I6epcAsnZWKq2hdIWEbjEhimdCBJaWpoUy/d38Xbkp79HskkoFEN3leMNW2R+LZD
OrI8qWiv1qomFJ+Eg7mF4ZJbjryODK2yb0aswHZLEVhf8zpWC5N5JNZVwkl8U6dD
VYmFGJmA9op8jS3Lfa4KJptzfIws3gYja1Cl2qkfa1VuK7vSbbFm+Uxb53wWL/sA
FXeKV5xSSvfCsZb1p7iBRT72H3Ms4axrjqVw0WPc2DAwOW3ScP6yx8+wvNDwrHi7
p56qK+gAk2K0BRT4JV2X5k9HCv37atV27fB1S0eSZ0wTX+V29O3hA5USJAA1qVJA
Z96/i6i38xl+FtldPA7mCNnONE7P64RQJINF/9G8/q1YwgMyWQ9p1ht34hKXfNkI
X6KeSqQyiY7XfQqwoU05mnvAYh2Kzez7McCeMYdD+KJRAhIuHN2hn86xzxSnBIyy
w7OwvxrOj57hn9rXe8FE+TiOOlcIKJRErHcRLV+FcHU1LfgRBv3t1wUntng4gMLQ
qTwhHBFDnSw17eHh4F2Rb3mzZQTzJJCuh7zNFuCK46Atr01CDYPCzHpEoF1H/ELJ
2WtpN4cgAFxHcBcyN/M+57lsyHkT393WQANc4GA9KQ1U2DKkw8PHJIdDNUILhHMQ
a/7BnghLcqIAQrU3R4eJERQZQNtpAnzC/gaaS3i9P8NDYlg9PBwkonqLIoYiu9V1
YMhyj0o8oVHFU36ZGirz05iPJS/BwZa4EVahWTBX3XWhYg9Q+m61qZybFY3ENTbu
daoFNhvLmXq3HMZlSwWg8Gic+0v0bzwp0THcP0bZD6Q8jWXuPCSivsAijC43lCdH
86aqW90SlnVJkcQ5MWX++6jtHMPzL8kjZRmIhUiYeD00w4d7MBk9qOtGU7ZMsXoH
V0vTWB/CrNH/Q8U/3ZmSxtf7DrSyxyNCBu9BAWdS8dKJ7wz23D+lp86e60cs0W4z
DWnz3C7yfV4FCEFSm7y+OuTIvpnQvNL3tpwnN5i8rcO6j9/ud/VM2EsdGAYq0qia
NJWf/RaTcj5qR+VSRTsPLa8VGqTE3kWufz8C6EuvSs0yGc2l2+fuIIzUHuoX1Cnv
/7v8SjpU6hL8m/bYhpQdYNbZdxBVdXm262tvHP3X8LRPFBSmXOd9dS4ahoAGwJAd
yWv/CRcHSVaPzlAEol3uyvXuPTQ59XYLy4wPHF34uGAfEvZRP5RaGkbrwXmQiyIk
L3fRkWNUnO2w7lZBoi52pZeKvF1XuaupUGM6L/sFyAZSv/cl2QiWm21Zjzrjk7Pv
+PHNDfhMJQHQKcuSm3WlwghusxkHE2Z2gz9b+zRR65DNpmm+XWEmI6E9bX/XeYaw
Y44haT7gLgGlmq6JHQI2VpirJ9kg3KmZ3bAFX1kQtaAVkUP8FYi9ivAh5ta7jOUw
OoUgByrpdgl/FgJBXkC9KbM5jGkn8jgXJm7O2bZ5VU4kXF6zZBAjUdo2FMLU1gcO
qIYVybeouQkfmlJw9Xvj2C67+7nHMHDiMwS2nJR1Ze+UR7+/FcsuFtVHN1xddtjG
HaG0V3hxem1WR2yqBRZ+Ftu+6Y7i5aB5eIoTCzueBgh5SwVR4tagl73zgabTFCPG
IxjYUvjwv+OJ9pcGbhS1sTwo/YCaLq642qAljI4M72h3fg+020p4wlAPXE0bkfKT
vePiFq6b04TNmSwA7GZGGEnKhEr4gY8YH8WHTB9Y9rzr/SOxAX2bozQ3Xen5wwxo
Dp1kYCADsPmjnXE5RZ3awBYkks7B9Q9/jyi/MW8K8FfDNyUGlu8vHskydtAexxzH
ZcN9Uv20P3NXFtwJjOfJC74234I/IRcxjHJFjcUVUPrvnDXnB5KyioI1LhLJQJMk
bbvzgNHiYi2W5wlc4CAlOkz0HAhFcnz8Dd8NwjcJJW/kGMRBelMPBN4u6aNwaUce
kbjpLrI/u8+lDGttZvqtoUi+GdUHDli8VOmUTRnqgvwQzcbPKs97FJ2asF1D1ToB
kzrwKa86i9dKbI30iP2zub07xkSNO3ryk/uRLlF4o0SGyN5s/fSMQxAVwLEylF8P
jZo8SSxm/kwFWqiA63As2rAmoEz0BzdwDOK05fLu4OjNkBLjR1vskM+t3qC/4byK
emJ+TORAf8J48gfNnR2MDlh8NnN4jXItt/S+V423SLRbEWFf6EvxwaQbr4NRk1N8
iEAz7d6qxLwlupL4ubemQV3ICnhLVYEAHT1/60gWVTnJrc5T+GlxKuqq1JHeH2z1
ighZoxxLU6mn3KN3vKNrwi69qVL84xd0xg+8ijjshY/FmGJKLQWs4TCCJkPoAU7J
h3xdIL/T0PM9SBr8PPXuncP/yI6vX1L2qGNTkU8N2+tazIiHxRnjgv0rM5LANKOC
GtIrUyVf5JFLQhDV/7ki3//J3XeNslNiWYxeyjKj1l513o8iEnynGuujjp7OhqIX
LDpdJ0FlVqt4Id9Qsoiz20ivffpn0wLEYILjkYkCOcGbqh5/Za2aP9WaDiXDRQFg
4htzrqkvXBZIswNvQI/xG8opgK5C0GL3PZlN19UZzXbRGjJnFM4MxXaWdOrltKzW
1CR/MM3nvHYwXTOjkoqAUbks5n7EYuTz6sAe8f6qLx4IQNFebr4b9qooDt5JRbjc
n1jUwS1NAGlY/3ptnJ4Vu6y4ZNXo7U8INKq8IDyFShxFHL+1YdSK4t3WVa7Va7ul
KAHfPqy2TXYcrHliCorGr8PBs7Cjr9AuDY3dxINc3yT5Emg0qoowQOj/lV3qfT3Z
KtD1X+fv59rc5Q/MSAzk30aNCQ7vhE5m/yqk4xNl059FDyh+caOzV0uavxvlQlKJ
+iK2TyIibH0MEITuswj+hRdAknCV3MKgxnuQROxsKpPCk/jb7P3V1x6qffpcneEV
7goia3c5tjl21Go6P4jrcpbDXohBxrWsGBT3rcndUYqL3BZ2GBXmdkB8ZAZ/K0dV
MwdArA/nqJuj+eGZ97VyQL57vZV+8tFj6dDt0OEWZt0gsFhQFP/JivrMZorceHQ2
K64YT20k7ThiPX9B1S0mwBrtwDAdmMNuDKGlZAEa62fMLHSG/C9q1jZ+N+z1kdZ/
jKajyMBpViHV0uS/ccVkBDoPisMUAghX4pRPWyRy2np34tE95G7h1GpA80cqYJnX
/DrWjxYk7jO0vRftFN3Pt2avuNostMajw6xqMX8ms4YlBFBrrgsWz3yuM7M8P+pV
GJFm0dGd+QpdjWSf+NkkOvucZhv8iTo9LJeuhT9S/BcTubnwhAiTkU7eCRyS7yfV
zFM5E0Yzgu0Cy7bafhoSTj0kosrohMJMDi9e9h7LeDEF0Tq/zdJg9O2ZNtQYZ9EN
jkN/Lh2gtHUSbvjIdjPEpd4vx3t4pCJfdGDInROOmtze1mPLN5BpOtN7c7Gh+sol
m/1L/sZDLwt25Va1BTV5wPUHKATAhd4k4m6yZfJAalg9OegyoqsMrFgqxCNZFF+l
1igl1GSSx8sVCKM6Qgli5SQQZoIf2LLGARirsGbIeVlBJRPLzt5j3bMtukj1d7ha
rayJjgxZfDFac0ILd8OkDQhGAdrJKamVGSpIC96RkWddX0ZdDhOBQPLc8jy+HdOn
OO71y/XDUwxYcsA0xltyikeAEQhfWc1lWQz4Ip9UfUFc+Utm6/uV4JhZcuenGwbz
2GDc/yD0MWt04+b7H1sMEzd9gUMwTF2ZVQBgWoRDk2ePNBd0j8BcJBgyHe2TP6s/
rTidew8C64m0BIzp7k5tPXleufehtpjIwgrkqIT/T8H3oQkR1plCR+ekTfY38vHW
Ey4wo5dRBqkQ/FR6XiqsJJsiS/7H9o9p5bTKcteTjQMr9t7cUp/2q0sUz+WlAl55
1Mku8rIA1opCjRFNjkRT/wGaN6XClmyJ4OHNOz+BL3OdHj0DuDZVQDxl7AAFi+Ef
Yoa+Hs2mX/8rlq5Du1YfcLiAxlUJnGKBNG/1G6Z1v33Q5P1CimidIF5HTS3vClDF
p/O0Beae1jyF2CprmuGZuUoNgJLIPo9Vbg4M6jCBoTBXOZatPLW7EeQUtH6PEd1m
b3/NgPyntNqTfLTX+oG4rr5S0eTJF7iwmGtA/wDw6hqaZwpKWKuiwCAKvlpY3KYL
NkzQL5FzuNfB5uye2O6R2+VBRzY+ZDxfFId/KBxw0wBQzUw5fuBeD/q7NVIG79Yo
FoNJnh28zvk9AS5uT1IDeSUmnCKwdncZGZ+PJ0O5HMTK/RFUYfSHncUJvH67W0Po
XExHgagTNrXzZhAloyNU5ro5So+iWeKBjqlLWPtqsSwN3vaT0/YvFWpw1YV4jEA8
wlhzIA0FtCPoV3RzOa0Nga6znvJ3Rxlca0dX2WA86Y4MPVitw+c/KRGRHZbMMssn
HzlJLoCiClyItf/JxhoDPrGx1FNdklYDR/v5Oy7kHGHiCyJO+D+Q7PLC6BoD8LPg
+kjSPEsDt3dCy+LCJHRP4dLR4BBtUq5ylF54p5LbdmFJf3pjDlP0zMXiZjp1z5wZ
SCcJ4g+u+Uzok4JvVEm04kh+YybDIIA9nNYVFCsoMFJSlTzSug4mugVzlLlcmSQf
51FDlKYaIN6Lmbfy7mPUo7LXWrjeduPKLkGUYytuciRdTCQ7gkyN0OB57g89c1E7
tqP2cC9OK8Y8u1NUpFxqK9tzu5KpXdAoGzORNsXPa63kBNFlGd35p0O0yIIx39fr
9LyiGB0337rqWXx378kRhbTZIOO7UhdRtDXmJr2VVOI60miplzuwEkKIKxuwIO5Z
zLD/FNaBx477yIF8hRJ3E7QOIaFxJ00yBFrIo+qOXsDiZFy36me/txGa3Gn8slZK
Q1qx9QHDEoJQ1g7asWdc3RIVzYgVnmqVhMsjcyir+OO55ey24JuIz7ytGUEvFTb1
O2Jm1HHkTi+KhX+xDbu6rbPIKfJLmQjAVBpbcamgYgeJtNlAs/w5rEPmYd4+VTRz
J1ZVhadQ9/aqObPi7CEVUx78B7QvTojyGuyRl8KS1sWykqLauGPUCQtEGUGVHIK6
JhV2QEFxN3Ia0ZkbWyfwZ5NV5IVoEY680Mf3lTPzeblISNP8FFtf65C0vdmyo/1y
um04T+P/T0BECiHcWcmL3hhba8uOMw6ZKsj13JZINl8k3X6alDyo43WfQh9dUmIv
EFhYZrquac2YzBqTKQCPfr0m/jqWs7dvSKm79eeg0DhoG6rHrrE9lmbnGEHBqNx2
xCiPEJ91Fvw0br7ahcqozd8fa44RqKLjUnpQqYx/NB3k2l9x8YbJKBJ6/VIUDe/k
zYAjzgT1KwDZtCs9DIRtHVP9/7U1XHE6jLJqpSC9SM4Z9XhGMPu1voQzC05Oyeld
mqkPtAXaYRZLnUWn62ZU+PsAooQby00rRP3tDw73fjsk6S7fDvVYXl4ZEWN/mrjo
oQYMW5slfXxpbqy8xa8Wst2GLMw4XLPnG4g5WmGoRsDDs8Ruu7ccNdyyDnLnFiy/
dNIpWwcC85o1LCaaO5tkpSRgh606l9VB/3BLhH/qQXxX8P6tWHpLhaRd1aTLuQHD
0qVNSHL9j6Inn1FUHPf7QImywQjh2Bsj5Xw/eDw1gRPRLRKN28DXAnj+s7D5iCtf
kI9dQEowj6Pu/v1/eUA3WwRtwla/HaKxARW0R6+7O9SKylKtSyXOhAhLZSemNGPe
3vwnKDGoKxPb6mHZMYoPz7tPAboq4Rj6CER9Hd7bHkv1zdo7Hgyox6hDKkvbbEDp
+zxKoRuzRqav6TTwxppoj5tY0gFIKzntBfXxqBG7wi/a2VuOBWWdiRnkjxPfp+gT
zRsLAHcBmRFLYkprQhsdMfb/zhlJ8b5l/6Unqc1CAPnljO7+UBcA/UtF7vUvp9NN
dAZWhGQgo+wbA/22RsDl9KrS3rKLSwPHkoU+psUxSrNYRb4X0LAuwEBAw7eUJXhn
fKv56/A/a+eXbEG5LhcYi2TzKlDBcp051OPVnSDFiQetr6UiPyJrRUq1GFxOty4+
G1ON0T0R7roqXqtnrNWdIEDWb3lrkfjZKAHNJUuZ9LTSaC/u45aG+ckuOhAc9AFN
pfBqjw1YGLBxgdh5KaEFbJkpGtqJ4topjwtbKxzj5nOqckUm4SGF+uOsrEg/cPV8
4Q6l+MkWCQzWpVVwMLfyW3ifu+hynzHfdZwqXMjlJBPqZyGx2iZmwL9T5XxELp58
gUUsaCnu+jI1GcBTFvk0AAS1ZtVojTzFOcTt3aQUfR3lpYvdtjgJ63pb80H8Qh3S
6FWOgMGi+ScOE7iWt3gParA7SrZ0O8gGREGnlggdIX/vBs87OObVH/KQn5qr+c7h
gy4K/oaWfq9BL2b0uwzVcjR3NoLrOF1oMWxnDm0Kkf7gPsTAa7h7EcccVGgaIpK3
YKxGB2U3lzffrvQrreXx1/zu3WXTUY22Cnjh8X62GVK3w/sZLtAQu8KrX2D6Jjsu
GGC7ZHOMH5no5TtuMEmKyzkTSLqfhH9FobRgI/sDjdXsHHo5f5QiGWtYFLBDt79p
YFoYYrrmDfsCumwDqLhb6EgBHfUB0a22GwC5u4iyusax18RpLLkdx1REmbMpz+OQ
SNZN7hx3bW+8h1iAxRf9LC2S87axpFwxutVSXSk6bF/szMYxVy9zXASoSwF8OiFx
5/NFmj58/RliSgPGUQ6GjQX+SKYXF0bG+yIi5tMS0iCf3+rPLhH+Pkleme2fIGrO
U/tmHa9tZmidkoiG4qV5H86//SDyGRFsLF/3G+rKBgHfr+RKiEWGadtjXRZEwRek
Ypo16cUQaw4bCV3Y3LaNN1e78qfGbH9NtK8AuEjHkgV+LySQsnNgwbQhgB1jJOLq
3dvDFFakghx0L8pdYHjM+zItbwg+uNzmpyfb3ZWteOFBUKTlCPppplZwq8zXXmMZ
s5pQG4//H7aclLTEFR2Zwa8kKbYszuvyuVrj0ivQIRQuq5J6svQdK9eBdnPFYB/g
KhDmlspj2HqPGRiWF20kmD2eld0J3p+vs+z0T2OyfT01FCBgS0GDLbZg+hBrzXV/
wjNpT2h3zBWf22+zyB2DBnjVY5iqweoM/RZUEKL/pJ7ZfEzDzs3akdua5EDpTTFT
Jy6u4idZ5LITI9wN9XALuseDG+nft7LQQM3A5bLnsuTewHA9eGLIHCTnlkhHAZhR
M5fowvU4R1wDTb0ynUScs5gXTGEQwBZEuEK/z2McO12EJ0Rlc0+yS0eEZRHBftFU
mmiClcNOjkYl1Iu73QP49MNWtr1AESx7+VPaXneFK+d7Y7wazGKkxRiSsO9AqNDY
dsj/sl9+vWTdTnCNkM78oTP62FnDB0T3cyKOjuD0zkPlxERDwU+m64YlLWSEYkds
lWPhRkinqmR0/s6Zm43aF/ZGw2YNmfPud6wC3baTtbLaoz3Hvm5rpip4vF15zCv1
lT9VTk8Jo5ue4/JcqTZgVeLEKEwoFXikM8uoZPsOlt/hm/2UosnviNumTIEARFMh
ilgmge2VeSou80vqjRl9cgcFZWIpUGmxM4nH36Z4MSHYMG5JQEom6iYofchckOdI
B6HE5m8KdSY5iQ3z8rTi+cO9yHeyAvYjc5kenRbnYdELBYSH4Mu1PAFOZQtYnLTL
WE11cutQVK6XVPHTJrGF1uKgiWjohgKEu9DyFQeXQHPvvlZSudNW5K0ZKM0rMWM/
YW6lo7PWQINUOBnpSDbmGnuSiYa7wWTIBofgTxT3gTZloNoH+pRAiqgN+xxj/di2
53vCJmB71fZ24wdZiK6h9Yl5n54ocGbyyfP7daGTxUWx4OcdFHrDmKs+UTZ1EEJL
Snm1okIkZE/wMqVnDW6kpI2PQstuACMxZYqfEw58LgWowIi92JOyhIDQxkxY/ALi
Im4JXnWPik8obkif190IyIUA/oElmakQwDC29ERs9mWsUY2yab/slbZV36mMOIHn
UHM7cwdT/aPHWqoPK62BRxk2n0fXcCLDMpGlPOs3Sf23yWZ4vzyRXWl9kgQfDvAK
XrLT0tK2k6Qxz2FPJj56yZxDNJAaev8M2kVFhJKdjqQ8rws+5B0mbskeiMKJDPVs
1bsGZ1e+pQ9uBK5UkeyI6XSzsqKYdARr1UIWrWr36EaPFB8Fn+SNbxHg830pBw41
/02jbZwFM06qAM4RW/muuJfVkockco6BjwbRC0Y+ilNRvdR8JSASLNkSdBpbBA7O
II+hcHAYeeXTaT0c/j9u94iMG5zou6HiYSeglUGH8fvpI0Fw+gn6iEMaXLH1LMS/
mKjARbaeNBNnAD3uIia8PxxZ9ybfJ2xBOLF1mrqenIkhMs7bEMzeSWENz1nlllKh
4PKAzIFkUD4J7jVDQTxTbK+zWN3Hv0KOXLIrWkv7573vqXtP1oOg9NJ1XlfpE7Hx
7vOpftS4mQ7sSJrMBPMkKbFfF3xD2825Rm+m7azzNWeqKJ8jkGEyPWBbQqAJlKHO
oPGuC6NrUdHw8bF7l7fIJP5Ry6Eu34j7hMPANgIjEADTevNhMLbio/ilB9qsmXVL
l8HBv9PfF8tsFZFlk+CCv3DSZR5O0kTaBPc1jCojOyowYxXCjjXlCGQT9sMGDWFD
bp/Gev5bJewtdSD2ue117jdfdfOSyIy+Ig+sUhbEChO36kQKHAjAl5DB2Y/kpMau
Em+NsGmBsbJ0bGHSegvVNlnffDpZShX5K56ZP8XnRwoVda02JbH98+JkQYrGDpQK
IeD1a1J3MaXtzE5eLvBcFR2SIivE8z4HLArGb/Ceizefyrk+T16ZvNzTjfS5z0IJ
Udsnwbz9tCjzbo1CDibsJAou8O544vVCTPbUKAzR/mSSMtF476hYU+/BvvKJv89M
2HLkV6r1EmOc0NRApYrDBaZKi8hfMv0ZRbWjd+Wlk+PLjd1f9qBLyZAFeZSDIr/6
6tKQ2+AsxIJRHOy+GvbiJCQXreGgMqOV47sctUFeymyxIDVB+uMi2SMhXE0NNo/S
7v1gYyxrxRI1CMSdH4MIubZ9GBO+Ax9FIb274QenYdvhgTKV3Vcv0o2UrBd/Ocvn
elDashs2wj4jNdc/0fsRBHl2NyE64Dix8FKn15qLG1+BEuct/CmEqpcOCaWbCrqA
Q0jtLJv2NsOOPfNSUo7xEZWoo9LLBdNKqklD7x/rDkQ2CElPCGBXAMWF1Bju3CEl
RQj9e2wtN3PQIfCfkK7V3+El0xXNq8jHI8sUw9ScS3tofrw2lLv3MTut3Gqy0G+U
J7QVnr41YaJbCYcX7txFOGWVwYVU5W0zcXUNwOycxmPPPMet5qaYxncQDbyHVyv7
RwY1JJseJDgx8nTNCHV7ziJHvs0nA7e3QXDsykbccnMS3Vs4gJfEm9ecunsAL4bB
LIl7+wR7AgoYw27KMPH+IA771G9f3WDutKcrlwvEpz/u3gKrU8atQPGXkm2yp/GU
j59w1Jk6F5coZp04pm0L18tfEIiEFTBi0/OWzX01OkzMUuudX+FLDlREWg8m0Tlw
uH4iT30V3+tXqgU457xNJje3cgRoehYKIfomHkdfFy6akaHaLLf881UFa7LXFPKO
cdQ3erSLYqfnMjJaQ7kcXNGaQpJREQrv7k7sc+tAGYq/SmIBQJNwx6ovV25WXisu
MQosWHnCXW2kVOxHSd9PQW/XjRZ/Gv3ExNqb3dMZCWMtWwkutZmXuSo17NcAWzix
5G7SNDHhjIdphdRrABu6citdio49GJpk7vD6U+SM+B+arzueTxC2Br+qVR7Juvpa
usJub/MTmN95ACfOWChqPglVkH71DHYi7BTkKKMjbjx/201TigU2gO6LzvAVluKm
HeQoEzWPHw5t343UKWkonsxDVHCTM9KRTB4J38opxkLspvlxxt5uzzx2s2YhoTa6
D7ZWF6hzZPuPpwU0MpearMZaKeytxnIBm3kZQgKBo3jbPgkuksmREXTW00tF4YUM
7rZaBukpVSytQQR02Qg2iFfYbOkSIXeao+Gr9b//pt0uxSnSkYJMQBPa/K1rRq2t
IBljBthvWNP1d+bobhCdQvZEpsXYi7N/Uiqh3wJppaSvx7Z2jYtzaQ5IRO5uQN1R
wUoFGzXwyT0aqWb3szfUNzzkQ/cArQFweRgqr+K5cVaTfInoTxMxZzI8XvXRNxWF
rO99MCCG/01jiQUe/Ii3waWvlQHh2K5BxSaAnLzZCZFPCet+awdiNxjOHAz8viQt
YSh04CU/Vq5SpZP0LOI85nryi95RPjhVPTGahBNWkW+wkdL+S5pq8AQWWWVtZo68
qQ+29/ZDKq3z2cPglz7BjInU7IBv+wHqmKfkZyqKM8fg1t5Ew2SnJ0IAqJRGdV4l
5PwqGNjz4c5SzQT2wfaADKqKKIyzyx+cDT/U0yK4AUJCXBfs12PI1Zw43kHr2Ir/
B0F+ZX+HQcmycYQQIdBLL2kwlEvra4x46uowQd3M7pRSSSwfpZ2JZfcfY+7/BPK1
2Tb4IVxEkmP/Eqr0XUgz26oQpBtX0uiicvzcMbe3Vf4905W3OmyiZO936e2B6x+x
csgwCHTybpOUyGL3Y2MIu20MaoWIVMFbcnGSkIuvSREPsiY/6hRVUupZvg4h4KRC
MX6P46M3B6aENRCq/ZwOKWw/EUxs64n/LJpXAbb1LXKrScnxO62YD2uSryE5ayRr
LooqG+GtQL3NGDcViOuo2Q3qVaVcMTzro5F4UUDiReVowh9r6TuOWnAGs/JhJqOB
NCb6Lzht38lm2ZfNYlyLp6RY6r4yeuKr5RxErb49UJG0brwiX2IaEbqlu6zgUv6P
v271Uyr3sXE3f/AgBcEcSStRqeUrIlqtNcQwwzlRZ1o/+LiNjBQOoFou6qEmqnqm
JAgC2xvnAyr74Uk0T4On+IbrT8sKKwg7r++EkZYLGi4+4nG1vh+Af0o2VSIlI+OR
MIz1loq4jC555YF1azYamEjLi8YrzqczeiDT92YJV7LNAfsCwhqiuHqv5mN5F6HS
EElJ/Gt5nWiNCCK45UrnnZTTQ4qn7JHEueUxGPd0tFEv3j//l4o3DtUruieTaNzz
ViVCwo0Xp+A24ESfFRv8VxZg8PCYNf3dBgaWd2Tj8WKVtcX9ALAcpEVx7qBDKlf8
XthmZdjuwmhABQMBBUcZVV1p7ViXDUkr3VdW6LU5/S0dzjxWYX/wCfx8a5rBkQLF
uuSUKhGJQ/dppW/Wl+16rLf2bxmTa24HzsOZ+4KGYCdHkGeVGco5jDvS9HMo4jX0
Nua1382dGZeS7eAESCjp+ZSvQTwynYUlRYWD5DcHbDQH5Zye2Q47NY2LgkHogWvs
2LtiG3k0h4UiTQ0CKCRqRXt9rQBdJ7tKKi/lZvHwunnjCw6Ws7nY8LTExRNIB/aJ
bG14Qxi7U4W9hmTAYRAIXMBmdkPp6cNmsRBY5jLChCyWSGqQo4QsGRO0/cc/T0uX
v14SmXhHnyRyVOaWGoq/BFh6HOTlVLdsXUvB8qPcUL4L4kiDhm6w0EoF9Z8SC6Cf
FSjbdK7z2UcShZ8U0csRm84jq60BhIBFHES+1weNFam8LlAQ+uWpER9M7HSOA6Xs
knE1nx/GTIV6gkTopQ6NkIdeFdGnn4UNLV4DG09Fh6pEnbpJw0FUEW2SZnPAi4nR
2Yxzm/xXG13el5RDfdGuY1ClDkrs1DaENQGD3WFwGpocLLovm1tyOPV/TcAE5tB4
id0uiGC6fo2zDH7B4vR1yCLFu5pmtTDa1leW0RnOMnF7F4bfE8qLCIDweerczBlz
7mdHolHzGRKdNeKlxsynlEMsazLr51FTsOCZygLWWPXEY+GaN+vv92FS0htKRdqo
W0Qs5sq6Ys4/nLNpnbtDScd0FJM0nnoKFEpZQuo9j1k6iQoYXIjcqNuuR6yAIfx/
0DgfgaxZDTZ/IqRzoLmxpDWVXMxhEYL/5RUgoTs5qx2z4KK64WIqfD1/W8j/izNw
kSWZB2Nhk6JRiGjvJsCIpLvzIfxkeDntEfPJXf6zk7DssKfFfR1lGsonwdeh/Dfq
QxN+zvSGz3e3FQpCBnvvqln5QG4eOA+6jpusu26iEU5qOHqIqaHsEe9qinowgpjq
UXYH1Ox/JRxj0DkCC2J7we9xV5AUH1c5QDzWXbNnGbMROfQpVDaZrLooN2xXOJuX
R+r2drzSi+yq9J2hstHPLn7cTioIFuPYTUhhbQ5XQdEyZdl7xH29eLlGwZxW+O9f
BTkMgkOtT77n7QN7jbQ5erOjuEqXDqFMAEUShNWgdPhuHQO+SOO9JyKNL+ZliiN6
IBih7Tm/oLAaUrw2IX2y1/0Ud9DqlcsSDuFKtgTn8YmhsB/oAaruPrKDO+gFR+8t
hrprqc4J3f9bsVEaR0TXwh/B/JlwxaG8dmVMMmdpVsgE3CpJjBbpgHysMy/XMjne
s8M54189yZ+YPUudGcwk8fBWBxJr4lj7mLcyRLWiOv1DB1hYo6Tx9xjPwULUFVjY
ed7d3bwseSmZbWzRGWRbwAgjiYBy/Xu+v65kqcmcWD5VYBNNGL71jlBxEl43szTz
ajBDAArmDHfY2/y6LJ3Fd29fcf+L134ww5bt5Fuv+VpNJdYlS6S2HChqMjpFg9uo
mXzwypY8YRth5extmNzEE+5hnV4YSUFIF71meedRQ87k+QcZoUi/cM0Cr5Ss/qGu
1SeAL7OUDv4rHgiMwt6XPRxckNHLu+I9+RvmkmDy5TWsZb1hE/mncOvEMgzSBCgE
46TkkuBBj5WhqB1cPKg4MnpEpB1m1pLJIy9FTPbyI3su4VZyjLIbblUS4EFrJIGj
4FSZjhHu1/oAvvH6/Oiam1uGpHTS62uJAjMybp3Ok3NGZjw5ELisaPVU3O9Ul/z3
zxYf5OxjZOrxzeRH13RlG0q2aHCRCrAx2SRV3Km1WITnMeKIGLvYuEHv0trCoQVC
JO+Q5E+ADcAymECcd5Samz+3CXhHorM/Gkg7/snh6hoBzERxU1j3MkQI/sD6m35+
ewxk54zVU4zkov1FA8dyUe3rMilYv4IIaWzC61x++byiC8jpg3/VqON0+T7qCBtm
qE7qISHJYm4UiS8dcbD48dbCAJlKhxQI1jXFRP4O6XNkLjoTue3Jm42qW1r3nITI
54lWU+MHZujj1R7+R0ozcc86BlWGwXsMOVwoHWcSrmOWQFZFx8mLOKcjlKJxp0m/
d3hj8udoBwIxb0achqQGe4b4Q9Q3cPcAio/UfJbrD47Kl+0pnSiGH/wU3uoq4bzB
FMiaQnDCW2SUCaDeFPiR2bsY+8GKEE04ED2k1yb4/K5JBA/8iBziVQKo6OsZ0LFu
ck7UXLh7qTIEcoV0EDimHUfbI47QLBl1zftxVhJzmUy1Toj9z8FiCb8c+G7uapC2
waqyIDp5IkXBHjWdblimGqUi1FDREXvAvGWAxas0e67Alr0t4ySwHmXdkQVAjboD
zqchDGefYvQpXAXix2GpD2PSH8lneCdD1vO/uYubE70Va1onXFYT7y25ruBJUuFq
1NjJ1BOivNMGeEiLYy8WzTqpQYmKG0KnPs4yoaHD6wS+w5Mnl03RxwjZtqVt+RDl
0dvLOpT9L5nCso47lTnO5Mpgu6T2alzvGE2Z2xRFzOqh4hNL1pXxNfoOSBi42mIE
B2QwBILmIIGlnhCZXfnKCYvE+GRYZYVpquVb08YjOAf7dTzg8y2NplHSYaQXjiRN
lhL/qpzyOga24fw7I4OEDA3R3IFZ+8sbZe6qGUHL6+5LXHcorG2TUdo+4wPHoZP9
i2A+tSs1/NJBHQFNSpDVBSXd64z3PCMk9luGO/tuL5oZMgIXVVxE5gkHt9Y34aTk
R7xwyqN77anyEMAl4iCLbwZsWY0hq6FxRjegrD+EfN8EOZ4sFRu+q1FFVoXeHF51
+zTUzdW7edwhYDm766sHTzYdJthyZAuWsDAATaEk8rQj3ARGONAyHX3WtBP9+jr5
rOloOJUVRSK+kLnixigX7vlIFwidgim1rEmMAqFqjb0Wo5oTLHrfQA7fuSIVdIci
4/KnMMOAGO+f1O0+3FEjabEFlboIp238S1EMpwBMp97HYW9pfG4BN/4NqcOTRWQk
kpHxpKk1GOSNxVGXWTKW238D8bk5ewYpBEFOxlQzMRQWTLQyKdgGcuNT3DF7jrJN
xCKMoxwmGqj9IS6XqfuriejBAkSsFgiy/TRGdMYGiD+5fRZAXn0YU658jnc+aq/q
8e7Cc0LMWA7AiFb0jG0WRICQLqKX6/p4YbJVFlnOxhjaRcQ1Ea+rc5LxszjcVF4j
1SqlgJl4OuqHtKyBKNxp8tpFd4Lx4/nVFekrAHIw0dEBrs7IwrvgIMXQ4NS2XGi4
1KYdNeDAlLnuCxOnS3R/eZaM8UmbsL2kkzO0nJ8v1Cus3xQPktoG2FG6HHUAFRys
XvPOfAcXZWCZsor8Bl1ABWWD1cae+fbx9HYQCtGGOVlqDi1leVzaYZHaJT8wnU2f
851Rcr+8UFlh+nPBDtZzXC5hgACvP1jI7X+l2iDYS4DTOaQTUN6Sq/Tot9eOK1tH
HP5EiH18wBiGYEPFyCfsY+xytmJ6nOFfpWbYHfV0eReUPoiMlOTQvHDzftf8O+04
ADqcAsn2JemJRdNKRRMNHRy6D47DBwFHT1l+DaRKagSqEUKJtuBzwRAP2d2xkQhE
qVKQ+QF7Hv3musHjPGpsL+yguDrRI79bfit8EjnHtvcGHKIWG9k5oLnfLTNEQjtJ
TdaS51YpFPl6yn+6bQPPGgMSZxgcPW8c0APS+00HE2ub1hajqheWrCsNxqdFc8nC
CpZqwOei/dXDAbesP015D4X/W9ofBftbEH/9CHtTx8keJF2KP0LySLBDAyxZK+hS
hg2HRRAl6C99WYW+J2FXse6SjZcLuimbYMcfmURlDBffihuuOxfBe3pxN/Id7f5C
zA8bdn8pOi526lwk1vhCEh+A+f8mrzpySOYvj8i3Gkbb1LcvFN2nySKu4HUXcm5m
I3RvGR5FxomktJStTXUsRalhMI0VwaASB6Em8cZK9/H//t5M1tP+5l3+79ysZlqf
RYpoxiz8eJYMqtMtWry689dPWeYIlCYEZUrykRNOrn1FvIyJvkFKtrAaSgmaCr5+
kOhXA1u8NEbqhIxjjFU8IuihuMBFpsnPIVOAc6sStbmSuinHIuod2EzTvkFhroHG
FQ4nP/lJ3RD442R41i8yEI3FkluBJjsIRV3z7eb/bTK4PsXGECJBhW6YR0L8FRBi
a91E9HeiJAPihQIHAHXhg/965T/K5oYWyXFWhm4NkPs3/xoAdpsNsQ8lCe2ZvqRi
6nf93+tEUqKWcTSzQMwcyO2UNNt0YpfpRfewxmLxqhOBfjWvX5Xb2bQ76d1bnGgX
bS2ekzs7AwK6BDJ5B88fzJPID4g7r5WxYBZRnOccLMTQouG5MeQgha7/05nWuIUx
i1/h44MJ23+wz7mFDFgla0539IxY7ekkif0SscWlBcQGMi1EUFHzlojTxQJfGQN1
4LC0ZBoPwlU/xLdRzwd/vHewcg6Tjq5Ts3358zsTXj6vne9WXlePZjQyTz30vyBt
3hO3jcNiUmKV47uFv8NLFNEBcILSBoeAPKv3oHqNYKXF22Ee5aSvSoVfD3VfpS51
1xsPsJPiuF7ztQetA90ssgPNzdT9gPYiAk1MvCFINYceFoT4YipW6l5iQm4NZJqy
8Crbg1NQWteqmE9FNvfLzV2o8d+GKCeF4jLRZHru84hAU+vFSKCo6OZN+5NCz/jT
cZ9nych3xsUbldJP6gRv8OWJ2BtvnjOMhAh4yLkaAySzjeW80K3Tv0BAJO0KMwx8
axqAzgUKk2wxb7evWuyvOs+dnjXXBgRBa6FvLRwCtOQHdPca5nF3MTPZf+a4ifKk
nlQZOHfO7I6GJIQRjdEOoPV46nb4iyptYBthTll52VMEIfhxPxtJNmFrAlcePXUt
y0sVSHq1LRaMqGheowcyAZgvn7LWsuivvIH/6tGXaCGtROJ9BZZD0a5s+k8RiHa1
Fdp6olzvIfKkOLv7F/GXwMTYU2RRkCDVcyu0I8pa5AWPM9zHsF/HeuSYEWoq4lmK
o8H2/WAz6sfhy9Zz8BhPxhnTil9obO2HgEmydqLDB49DUvNAv5UUCfXMu02akBfq
wwikAdCGyEj7IDrEPhO/aWNOsSvF+IbyTrZW8YJyluRYjnrl8OvvB8sWuJx29FnR
2Gi7AN4UZj9SyKbofaILhZqFvjc4R7KLEN761i60h3n2RlEBoCmwXlW5E6Pdp6j3
eQNqlNPUMtN5wmSYUW/3Ejep/CijAHWGW+YbksqQSrhT/qahxeOGTER6gQM/huYx
Ub4lWR53VVNDxGKsJB1qCfJRsE14MmvPhH5HJtBDeQc1mw/YOX0kiN9unTjFh5Ep
lAgNgAch9liPrW36JOcz4X/KsYzsLI0fBC5MPsoGe4nH9dlJ7YzvHAKqrcpewDfl
GKaV6MuPlUSX521zHJ9phG2zzaaZ2EhF/TLRmiqsc7yRwosLKNsnL/ZNuCFh3mB0
bhaJZWXPm6JMz22juGFQ6juqIbAosoo+f5jzFcOadohWwhsoZoUy7bAJf2E3ojwH
MafXPNPmewz4HZeQYKrWWHHb5r/ha7ElwV64NKiqieILi+Nc0bnz9eTm0A3svQWl
q7QYmlR+bAKNh4ZtsijOS9Z3lxxivbhXg8mg1TIbCiMBKTFuan1Hd49GTK5/kChM
43bTtcQ4D6EBNnVpxrgsgqhMZoyhYDeP2ZYU/o6XdjFwdbTm+39v6ruqDD6QpD7o
wTj187X1TmEtb7Qy+AQ6i4RT7zU9e/zVophoxEtUgjR9E1S9efgyPH3zsFnoCc5a
PUL9IAsBNV6irqzipPTmbT3hkxHBz4H3KMQ1xisviB+Ud5MddgRMKUH+GZuVCEMM
DQ13L8C3CeD3JWCv3iFlbaGYCtazDpaDv/yX0OvZK5G+DFxvUGTQETskZk8jnxdB
EDXu78CFirXejhXnJWsGu5B5FBvfDOwlPwjZP9mLNELd5hVgrXpcgPCdYEcOHmmg
uMnGomW2sKb2l3KxgNFGWCq5PRGsYQGN+O5OdjQEsWQjd5ZEyPO9wHicbA6y7omG
7+Javq5CY2Kt0hNJv31ncIz6MnpvaE8IAAtlt/CHoBUEcuQRGioOl6gBNaiRm+mu
AIdHSkYu2crQdK0HNW9PZC/EwJ8BicmKGEo+/8GxOzlecPp0u7OqGdZvKNQ/+FRZ
bC2BKwlTKKHRuD8vMDBdkeyo5K9cvXo+h0kx3HQmGk+6GqhWheCIKX6XIYBnMtaS
kiKC/3FvWcF3vXsffw9GIV0XFHtW1tcM2i0faAfucCwb/bjMztVUprWlVkDDTs+A
nCGv7od5WuWceZFw/7XIUPGw/EHpoW1akfxMk1//R366Iiv1P51vfoi0nrPmG/yj
x+G1emBVFa+sDU7kVl28ovykFH6sqqFT7HM3LlkfO/qfMiL1dC+DfcR9FzNrxbR+
YpQ3GPuXjFKb1hirH6w6gmft2ETnrj/cZCwi6cS0J/VbmTN6yDvRTm/p82LYJgsw
UsH1b9h5t4QCWIhh9SENJVl7qN69CUXjSrjsbjhjcFlvZqfRe1kw9kXCXbJfEkrU
twscfjRAhfw3LO8preLUACWFdm6/M393uO6DmmxkHP2QKHDFR2ZCfmABJ+b2cISQ
zyXquLkMejvAHdbKtbm0wCk+leB11FmYHciwrbuFTpb4JiSkl0opLNPrqz0oTB9Z
ufXX+NNCeTkUQMvF50lN4hiqnFz2h4Nbny3Eq2uI4Q9Nl0DY1gnoN8XQrl2NJuFI
p+DLKl1cdU232vlnPcqt7iorR/2K+M3+bq45TW2ZtCMtgvZLH7ojGH6LK/iLG/yH
ptzQ+N8lR57/mZrTYkLS/BMhlsam2yzbBRrp9iDs57S1o9JCNx85bqOz7/z2sX9f
MKs2LMg712OmCzKW88TQfMmn9OfJ+BToAkChCoTQyfIj1ZwXDsVouLRzCQ4KUlug
OPnoKuELWarGegYFKnfEJ7XnshdP/ALxrcHCqLlEtSyjR0lqFMxj1UHKHlJvlmOQ
+5acxxbAADsNlFUUuTX2ICbL67QE+FlbNcxACdXPxli6tQrSaDS6SvHlZn1KtjEi
xcoUfXWnubwgqJTN7RJXS4khj5o0Rh5mzSJBhyZHoVnUQ79DakRzpEr7Y3799TkH
2FvvlriiFdxfrYCUueHqxpFGCH7yiB5nIAyYXysrONjq9crbytp2RsQVR5v9TfRH
cZ2oV5jkywl+nzhPOX0QvyRm0vMH9HB2ke/uJ2NgLYWyeiP+APsiCCNjRD8mTVBn
yt28uR/f+mc8FiZDSj5PSe5iT7ueYUeQnvdF3wS/BWRKlbJll7/Tme+Zgk+eWgl4
xh+iDKTrWRRN/dFVeIWUVpKoYln+W9mVdhBfRWLn66lJjrDbV9v5SxBv71RCviFu
9aVX1TnPvPm/CamqiKeiVIACD+mTczflSE2ggIZC4YKduiOcxITWqWQeTqAfrqwA
hOQ0hG+x8L+RI0qBln61QWAoGNfB1TgdMzjk/XxPc93pjhKw81haNE5PUUe8SjkD
LoM0I2LHn/uQY/aMW5P6Qy9aVxAsqSR33pM5sLpPMxjbXCO6Qa40sNtQjIaBI1TS
xt0JuUu8FGUV2TdyrqF1glpfjF4V+JLYrFBtXCgFUsEtwu0+tvfQMUmalFnu08nC
DV4fWMH2d+hf/P3u9WBc0bqYnMadyU8ksE5LgRIw0rnHABoiRReLCNo/12pgNrh1
BdsPtKk2KcGQEZSAJjJOSXUTZea+12ipdsL/2MKIeH9teWXj2YxjsJ6nqjp4eQO2
V9d7L0HlQGyjbamQP2r6wk7p1+Gj4uoi0vfHivzxuPQyRM1I8Rf+6vnRW+Z6ile7
03AHApdUmP7I8QlriHwjCLFjll/ldj1eF0B8vc9V59u5+8c3DOMiQPzj4z1An2u+
vXxjNH7fdUVE1uhAZwHqW/G/sWFnPS+M2Dhf/YEqgnP0bIJe4Ol/ikS/bS1l6xbj
p5V0TpiXT/PxSlI1Vk/U8MdgcQ9L6029T+SWLtfujLGv3xH+IW9wwqgQvm2F86NJ
wYnDEqLSj05ZyD8VJllj7R1YGpphH3sV1wRnQWq5y0fMWeg2UjKKd3veqQxSKnP2
L0SkNgHPjbJthBYcxtwSV95pTfW5OsRk9uhMZDR01dCMz3IFtkdPh3TGBjkMiCuL
SxaO8Q0KNkIU8jnF0xRbqmtirmjnY3xTsJsh14ipCdQ9vMMTiWXAbpGtIHaedEKr
jHS+ILVAUTGvq6qfpt482ZMMEJDChiYC4zibx11uD5LNDJIbpmThZEGtQNKz1JBA
jmZxpkRG/JOBEws8l/gRTrnkvh+IPNbQeaeAXIA1zq464QxCeY38RI78GIRcIQYi
ODIOKiLXwMMjsQICPxGnZzqTDWY4bFWPAoMB6tXFmrAxq6Z2QcMu3lX5ttV4SraS
ODyoYDB18f0iRG/YKzr2VD1cLCsreB90Fmvr9uBE60YO1EUUtABgV5dOWDSlRTlh
lv1wfiuBTlzm11TorP9OLHPMoAwX39nUOVw/F/UKJ+XKjE1EtuknfZuNrnL7wDhd
RE2f+pBsJ8hu/h/H0vqYN1WjuSeOFYydT3cb9ASEaLMh6KdidS1PchU+X71Z1bYH
Bor84isjrPzmjXP69m3cVxek20i6fqX2e1BDZweOYBBot1tYWwT2Yali3QY7aek3
3//003vRmWKymblNAAvqvxwsujefpXfKX399Mj2QxmXZz+A81P9k9rK+JzbFdEou
ZWlsTKDDXiYnL892SOyF5OxsIePaQbOcEVDqZltpTl/WkpaLgszrxO4WBhV4HPC6
JfJ4QITSAMpxRHIOsuApC8sjDNbERoWi/k1JDRnVBBLdrCQO96htZLEiSO7972H7
XMluWWmdUGeWHBaDiJSXyF25xCpg1rqwhF6zgnPokWBB5397uaE7RZChrubP1GfE
ZVlzrWZbNqye9qb4L2Ggll61+awKzZQ8teyYaLvziyL3nj9vnTClRmX8PeZienkJ
sQ94RWIIl9zUQ7MoD7RzRTKW8dOk03okExgY3+tMZRhndDLMh16ubvw7+nEWNJF6
LxUm35A+O4IPOC11U3EtNAmEnXrHtIo7dzVzsINZqVCJFVNgGtYldE1RXSCAN3c2
Tt4YjBKQHNxlgNSjPiJWZo1ImYOvSIKBoAPWlxtafDdt1GJ9pc2aNKdPYrACm0zp
qx5hkxy+W7h57QFXCSmunvQ+uV2idHvF/NNNg5UPqyPTVNOXTwsPace8WOH5HR5J
bgYjZYoDIXm99318f5XDuVmdV0MX5tEL3sgSOdj68kk5YgVCI+/rlQNn9p4vSN5Z
DU11Ewmx1/sM36VovjdBtiw4FEUbonlYD+11yyGRXp7ay5eu5aLLSH4LzM+GwGuX
PhUKGR3SJLmE8+UmvoecXW9g/LjyGYHIDoZvytFijr9aKwioxm4GH9QKYFwDKFSa
dEvmUsI14PkfmBoLWDhDeD7Dsl1sLOMQwqAk8eHG40cu9pgX/LPc64BuxmsNTRlJ
YcWcFEe2CE1+O/3/smzXsd82nV6rM8QMzXyXNWE68PwhyF7oqI2ex/2QHqIE+l3E
JvF8YImw+14/ix+O+3ZYkXb0qm9QQtvx/+c7tKh1zzSbHPMBulSCDrxDfYPoF6OT
td4eUxhxZ8HSf0ejzKeAr9YHzLSnJcsxNi2DiVGrccQ9yOA2KqQYi2h2rDTj6tmB
b69sxDUnanq6GfPZNW0LaF4TB2i+WC0dPPakObZ/QU+icOyB8/Ggx6Jqin5Yd2V/
MWS8tfoS8hUvrD2cvPAvoYPiqh5K3eEHpxQGCwq4IwKtIaLffNBj2hcltYf3LM7V
bYEB89EkvsDsTdq2WmWPSsoBwbSw+BkarNGfFQsmg4V6QcfphrCb4wSeAh8tzgf8
nWz72OxQO6iryyNsa7TjyhDOL8N+uswBaOFnO2cFCaWQ+XitON+yOqF3pQV4F+3Y
wXo6BvDvNgToc6Jcxb77/EYzCDmSzf4KBDBmHYInCawjRiRnTjg6w4BD1m+LWCGh
74lNCWcjibaLu/BFZjVbZjvhX3/kj/6TYp9tf+hhKQ00N7KXiG8jP5mOdTEap+OJ
WCMUahEh1hD23FXF8aMh7+C9X82L4/B0Q4YCc1eWlYoId544io8YS32RldezgbFB
5Qash36mFJosxgledkr213cobTPxloVNZ4G33nkhscx4XJ5Q3/pk9xK0ne0srCqV
q+mp8GVIcWCmh6owAseEJ0CQSpefacm1VaMInFZt+oG5IUb4NmnbnJVB10VYnEhL
8ofakJo1uy2QkcHRccS9ZdZiTZn9a83Q610JmsLiXyz2z/h6IyBdFDgjCOlWlwxP
u6OO5ukpPjgG39AckLik3xVsQ9i9rMgcaKIUF0WkX3LTLAMvoYewBLNlPr/Kl6ZW
E+TaNpMkUgd1e6BvP1QtVUIKetWry//pHjRkFe+ZbBz/xIJFPn47yrKgE3fc383z
6iR0mcruLEVjVt+65rpiUa0e1WJ0cnLDi78u01VjMlEIoONoY2n/JcxdhDDTSq1/
3xRCkT0fxIXarqb80LyJIUog/UgVGoQ+aF0P3PwGf523AMUW6l6RjMhWTPPJuqzU
FBhcXovndr5cdY7OaZPhbtNWcSWftQKvF2WiNrZe/aBmmsmT3txPaE/Xd1TU2ckb
/4ywkR2Mdf+qyRuBTgAT3h7kqnnzDkZ79wcWKyoT8DRZq4NWnTtRsz8jLLIOZDKI
w0CNY912RsxMxNYxGu6/ulnTP1097couWTyfg/9nrUKmFKbFvj5W1wEkVfwXIu+D
olOWJnCUJnIy1NCpfXEwM0oxb73RQWGz+UF2NL01sOelgGa7TyHvaDEWYfY6GzoV
uV9vd/GxQXfZzz3SI2UXxBQAyc66MMWYMvchsn2iSm6mPP+1MLrDUIURZvcJ742K
MvjipQY71JHn85K/4p0OX/nGI92/xTrazNMfhnGjBdFCGj82kUZFepYFBzKbWYS3
zF3mAxmXFs7V75sIvVVOqSfiYZWtqyX29GxmN5pnVWpH4cYPN78EJvIVdT2ffuU4
Unfvlce7JIkUhGcs0mK7Nd+nT6O6fZh2tqys+MaDQrp1ljDwk8yB5LzTsmgyhTsq
d49obfLlVp2rKctWqTYVODrIniWD/sY3ZwxSH3ZZsciq6guJIsOTblzksvV3pJj8
DAFSCfwDEvzdDhpv67PfcvqYSJqGmumhnLv8WuIxoELgRCdAa41BB+zXJUA58crB
NvkU9zwsw/oziBHJaRHM/2HprG1u8601yc9FhyBd0WZl0fUL1I4AkJ6VvedJ2cO8
JOdSeRd9ys7GXx0/OiHDqyABS/4MeTGGfgF3lHXLQW2cfVNgxzHDKKltKbrrFqn6
45OhqhQFEvr1SJrH4y8+DOrc4OTL8vUGFAwiLTcYdZA/HQELEBX5Gvsr7R16vnIp
sTgEyn1//8/4i4dNRzAo3LuqrIXVoLgsvjdv16XBVTEfryLCM07VDSFMPBOF8bhx
VSmiQWKgOIQS/b+msWD0q+vIcLPi5Tt44EYczxQwCyWQl0EedT5R3bZWONi8tWb1
PD6pCmmwhn6ynGpdQKFL/rS5QSASib/AEIbFxiHyNVqpH62lXfOQTDvAaJ4lE9FD
DINh7ZfYXX+ifUGkAuidERvnywYzK+XmkEqjOH+uNSpxI8HwC5iIe7u6IyPV/mhV
HIsaNiQvOYA/RvtXNVZ5Tn/XXikNNduOGJ8Wf4FO5aYFEcOkbouMXpVYkjTT+yJG
ck8uN/wJIWKfidPpfNIoQrE3PH3aEECsm7h6H7qqAuj2hJnOuzQA/0kBdUQ0fp9d
wNXjUsdbba4nnthWbnqI4t5sqcSN+yhl5FF99yjKcdBh18vvkuBG5fH9X1WwSQyQ
RRMCacBx6QKi/Eg0tvv5ysmhwYIVe76Ru/WfQYkqEB6gSPU6oH91hktdqHJhW5d9
Ie+lhqxrlrZxybWCz18sJ1OSqsupfzWa02Dq360Tvoepc8MSuLLg57Icz+0XtSBB
N6ylhWi5gF6Y5ODgczLL8MDkH8C/6S7aoTg0P8WIko5c3xBZL3EUP3NdJmp1bZoO
XjIatV3zz7Au3oOHnt3h9sKPYlrL899+IFq8iju3vO129YVVewb7ISzrvtkJvkHn
pZ+w4UNhEnhJNyO93GOCNIpul0A13/Z4l8GQm8esbO5lJqqYuVlrA7Wz1sz0nld/
8GuQKwCLRuapfgEBM75OCv1vkEfqN3lIalOoIBZHu9kNd/ex+CK+h4MyjLC+WOLH
zJjx9hJ8hohlfNsIGARerF2/JBnFg1xnEWksjtVxUK/DUsY7y/7GvK/VD7j4y24F
HdFpAalqDJikK5W9bGWxOpJR4ySvGUqFSEzGIKZnzELCbnlA3nPPg/Ypqo4FBrgJ
bVpaSc+E69ACPzNw1I5QCYbIMzdD0SCFlbVGNtStO0ejtt5fPI68zfae3eosFhsC
BP2/JxOU3qSNmFLqr+8HFzX1oPAwnUOWr5c3QL0Jtnj3NwML/LUS+1V2SpTm+jTp
po9x4S2svDYpA/JP/fvjLHPA8Dbcvn2KPZMyn+bI9zg4F8dLvR3OtT1MeZw+/fIP
uo6t+BFSqc4O0Zy63fxBgM7MupUO79ssbBmNNo1Pxfc7ExVQn3XmgV1rLp3M0A7c
62NKXHwl7jUlDESHBIPQsGOaXhckWiIkt5kKpHUFajynp4TsK7kX9IGUCrZ1u4mO
Z7bj0qOxHUX0ckEtr46AZ36suaTtiwYDvBLxGBGO82shOfe+bsSPtPtzbKRjz2k5
rb0uLXKvbUCpggyVkxpmZhaKloi721KMluXi53StJkcpcFV0OwaPrWN8+ndu3Vc8
FBFej41Me4+OfUklfiyE6ve/vhge8D4sHfkLM/4AIb2V0LPFFrZNMKrpbbEPb/bL
aS2TAs9JNfzpa6HEgM1OFVdZHdbA1WAvmd8eMtSCFxsamSjH7DfVc3zXrfZam4NE
GyaQWqaWm7x1pPIu1+3tw+i54Iyj273cq2kmLDOj/cCU3I0JTgLU4/C8pqRlvbeg
dUZPFO3nQiO/WDdyxgFvR4JyLqAY7GniZaPbS8Bhjkc59PEB8TymaX+lUbUy41Sl
xfbgCjKTi6GgB1hXJFnt726msJsmgSLmK7/blFbrtfYncdnzJIrXb+FgVH3hu1K8
rGFxI6u5f85Rwh7VqegZcgqmrYyc4fOiHdZqzutuQs6KC4K9e/3T1B1cPxX19poM
cZfXZ41HfSKBrwDGpfJ2RDBda1IliBTGrpzhr0hGeJMU25jkiN5mxGQdbp6j/Y0f
KvKpGUJTD4mxCM+XBuxj5JPfh+H7aAzlIzekh9d+uU5o+qeaYTwxQOswWXW7MI8e
8MCUEkNLlq9W4puyFqAvYRTJW5pEmK2iYn/N+eTeMbJ1mBFHqpacCYNGh/eH10y+
Vmn7vAr2o4LeeSc3DkFscHC5vGxPO7LAkW55IkOrMQ9Q8D97nybCgVVQRabo9gLc
dvUMJLLCGXinBOIsXnsnq57MUY2CbbFLl4Y+L1E1WU5shZhv3oVsQ0lTMmLwoNRT
xJXrXSSazbhHOS7OCAwxlYVPNMYJ+BMbTs0lwr6q3LfMn+r8SQlaT489wxvcFvw/
TRyve+kgOW4os19LYIeDbUbIOlBxCZMhRi/FoYqEHXm1Pv7Atpy5LZsgaFAv4cFW
Hb1dP3IT36Jn1sjcsa2C9y4dWye4j0rX/vfEqoWgXWAm5Obf6UO6sRfh94LkOM1t
Mb7qNc26S6x64nEdF1CSKDAOFNIw4dC6gAkp6jE8qmIux365B7TMqXBjqOYVxP8R
inUZFlHD/GBU+nmauoRWR8MNhTEjWbycGUOlmiP5RaFxQocbrS3Oy4IZczacmRoJ
6V1z2t13OLXnoGi+mxNT6SYlDTsYsOmEmUl/exbNJQlhjRTszJq6GSMzr4xvS8vQ
wnaRe3QNQ0b/986NasF2BHioamVon052LkxYLhxuhhlTnt2nMwvyeQbvC3Wfv94R
V20NWfodoQt/I6OEDDs9KWqQYj0Rbm/9FwFKDoa54lWpYuvm1ttAL0qtDxTPu7Ec
DFUY4bEtfjdrNU2KCwNn7McFDDf1PtZu7c3CG/TTmGJrFUnMmazwAMDYr7+/xCJ9
7EpdILqcoaub0MoDOLUOInyN9ly1hoSRodLx93JLFQE6bLEEi3xyP3urnLJXBDs8
ni6GqueWRn2qptv5yxBVhAXAxsTZSNzT5v+GAF+J9y/gwl5qLi9klD8znipFknI8
gy59YpHFm5VOxnCG5KHBjfp3xhyhpiFgPdl9Vps0djYzHOBIHzIA4z5eLa+wGQqR
PAYo/WYdRe/ubqhCaV1DiaKN7YqFnotqd1uGiX2HKnCWcggcQzFWdvhKNan27p3b
168Id1pu52ua2fq35XVHSvI6FYNvoxF8qEDMbynwmUpxH0O+dGDRAtjUWguNMDSn
YOAN3xXz0MNICNAsROPrduzq/SxRz+Rf3keUYcES+FJP//8/Yr/PD3vENeU4pToB
Pc0x/wJunMVIxdMNuJYrp8r2zUQC4UwBWpL8loiK603c079RlsusVssgNGEUNtw7
mX4AWVHxvOdwQZyKAlX8RSzWXPWFe7qimPIZ2F65sxkwgwaxhFrjsHf+uPjz6qZw
1/Q/FMwZNYq9djhiGG0asB9CVnrWCRXpgbps48VDy8L7YETFMOPCe3P9/m2B4hIu
yphIxuNteAU1vtdHqzhtIQeqiAXZZ51lh+sbwcBLwqzELhYiUELL24PzV4Ad/reF
DB5zVmtoup7oV0A70KwiH8qopN2lomWWTKAOhDvyrX8nJgOncuqo05rbuk/jeTGR
+dXHgmNQYE0k34r/K6nzpZGDYTKwRdFzpPfswEuZVtsziO4gG5imkX4XNM35Wwrh
0NCsbZ0apnYxeTaicWTI1FkIwdKLRYxqAO/D3UNswSMJdnH4xgJSmndroWErypZh
sKrkwONgv6f+v9N8ge4a5upYFO8JOu1pNvZMoYTF5olVufpxB+/3Ei1hzh5oMZwo
vWnxMVYL3/H4xET7Hev3cF5fNrUDgQq+CxWRqBsGGYsa6N74E5n71Bc2ZwpMg//c
D7ir6zPdh3i7L8TppEMMbgH1XIjI1ExmcZAZ4FL7qkLh0/f/8YV7iwMNqUe+Jl+R
l4dFarPExGD2YZwNBFJGOMSoU6xnEa0UWU3BnHoz7J1MyeWVrLirdO/A6ORZ6+8a
jWaOcm7sQ420IBsrHlX5J8f+bih8u+Z1PGgK4pjct5X+y/dItWKuvHSB7FDFZq9/
KY+s7lGCKSR8iZkpOvC6NKrlSkK0NCLdsJUtq8CzVRhqLyLYubbqW+Kygjz4ns7v
ZWH2qSaK3MSCqIBlUpirQ5zfqfUdUiLEabuB/ZYR3tFQ+tpzLut7N0g16mtyWlM4
7fc6fsaGl8IQ9BqLauXmDB7XBbbwg6nHba2nAsrK+tB2AABPueSShehSIMBPocHh
p5Dwe3PC4YstjJADctGbbZRm8B30BO5z+mwpXUPFEVAeBjYGblPacCtbjXovVuwz
vd9DCBDWLdvbB989EWOmFUXmep2WWfwIvjhCu5yYR7wBq8yWrPIxohRueX6WGSdt
WsCyRKSOWlTNT2rHwdSHWEAyK1n/O2cZNxR36vY9knTDlGm0RnGNlOyrMpJq/GB1
Zw7H6M1AYzWntLYmz6bjSJLXBClNVGwsUokZg0HRfA1kkxahLLt5/XuOcPv3bUcB
ow+XLmDlHjIJK4Uckm0/Fpbk8R67U1Kd1oAeSjteJdIpRtllzTM0sMGaCL138iyN
WkSvh9CEtsxF4LQU67SQcIeuE57v2nO6qMiPBWr8fHljv4N6gTaqxAtVW/Vl8b5P
mqeSmXg4/8x334NQnrnAtWu+pb0mNelRxzOumzYsK4mqy/zwKTU7N2HjvgpWLRgV
Q3d5g3jMVVR66Fkyk/H0tEu8m5KJELADR1x2123bzzQ5UkicVbqfY5xYWkHZWiXh
jK0xetsVnlQCszOodM/OR5E3UOYb5FLo1w7Y8Wgu/iAOEaZHkHGA8z1iaj8P8osq
vGR6niWDjHU5mIGn9DCA3ZUjSY3Qyt4PL48KGWB8fNobUMHHo12koZXJlmqNvTjx
9mzWArCS5WdcA9Jcmmj7Qdy+WNv7iTHHwFX446Qqnw61yHoLPfpYZYOKISVNCtmK
w/TqR2u1iRU8qj91AYWjcgIj99Y3aZYw9ootZggl0t4Hma1TIqBC5ptplMPMv0by
obOhkoX+7PUnBxZjeAaun7jQz0OI1YBA/nYQsd1IgLAx3SMI46b0z5LFRCrNsi4v
AKqlQ4R2OT9Stqs5LKLFxome5wr5ZIuAk2OwOsnhEmYmow5HQYbiqg1Nzzmv4IZm
/DSDY8eR/dW+HLV+QohirLwWd9k6cX0xn6/IbUhbUATVYVx26mdXMWpi0wqnSmt+
KjBLrGEXX9VnHrpLvch8gxG8dWkO+l6KTCmeleNY1a2gId09N4r7+xDZ0HTqNSIk
4tJa3djAMoA8LMI8auSAepHMJsdoIFsoufixuLmXIK2QkFV3LTzPhcDAUF0pkR3B
WVMdnhw6uJyK30WYfaYismjh//l4j4lhb5yxH1lKbojUCuMb9iUjGebAalNsCnQd
3Z24F6b4SnOFBtKUppUxLzY9ikVKs5/8CQXD4loe9D3CxSlluBmm0y8HUE8I0g3s
wyvC2AtrhJlx7+OnG6RCiUztCwX/nDLyj8Upj47ykZBxy5ZrXu5YX0c0b/WryD37
78y7mmyX6iddQ+Rl2i3n5Aj6SWvgSsveRQPl59Lm8UsVzQmcfG8dvGvzavrKxp0y
JaRHnWX/gPIlxOYMivztbY83df0e5bUb0Nb18t9EHxAFVlx2NKRRYogfWQgUy5cK
WwT3MA/dOcYgg6mIpxJuzo3RFpkI5Nvk0hY0MxrSIHwBQpc70RqnxNcys+6Qc1Ld
ERtt1+mbtKkvtDDwO9+uijYLrBi0ULCjgHd1zllDToWWSjAYVKAt3ea5zl2qkf2z
jyW50nzdQXxktswb/lQtTrt2n9r+34RobrNj90tEbLLZGbUz9T8E3Zf3od9+gh71
IbYD/q71vRwB/Y3tEx+DFw2KgJ+6fWsKVdTE15vbA2hzdrFle2qBEirZr1bvf4F7
u1eV5e+97uxlN2/SjrihuBCu77x06zqeW4AiMjSHoj5W8R57ylv877G1OUQ/o1GQ
lJoe5YVhRVijTtknnxXMQe0apZHBYnl8Gc2x2lxPekpSICk3YlXbnM2pKdN9TLNJ
BdGy4+Nu/Bh8u1AXCcJRUVFBe7Jm+/Ax86po5KnOYXXYhHN2E5nFWelX8KeHrJKZ
fHZGLAp+TIvHRlfQ/Sdu74gHwTsP4bfGcNPYzUf18D2/Pos9+E5GS2Pg3Uic4hh9
pKbiKMKmsYf8a+pFFd7pU8MBpZy9PstBs45OYVtoVlXnjMhQN7GqQViUsZskawd2
263uXjVqvwdB75LVAOCo9OQ56FU/RvaAqm8EF1Bhlnx+YyLKAYxx0OPNaQOvAK8V
kM2sRoWq7ECG5Ioum9CwDVSZfqOHWddU4YUmiFYequrCO38M/Pi/bgFrX9S0882R
6km4pFQh7cvmlgg9j9AMhHpSLQHExUFJH2jFnEs99p8B6B3WVcNCv0uxlWVfRVEY
JNUwULdFYpHJk69chCF/GIGanL1nAxOELKBCTNg54zg26Gi6og0ehC0kFsRg7vbB
HIBSnMzXlr5GsvllNtVDHJUJOU//UuRgiI51cK8G+spBPIk/wCcepaBqM/G/GZfr
Tx6YijW8EpV9sKrMOqPObIw8GOx5CgJBIl7H+yLfv+nOEcRY5CBbbaV5t8qBfnTm
eOxjy4tLvf5ahav9i3AqqY6FlhJWFoecqgT2mOe4VBV9lxMIXc8eSTnq7PDU3l/h
oJe+Ol+mNcAWXRcW/mSnpl450QwtYB+cu6HHMs4dMElK6Ed4Lfl3OwxZdzh0DJoo
J99g9Vdq3kdBgQDRRA/pbFBRXWQRY3SbPzZ9FzmxEDOR26hE/ZKtkZFquFXDokTo
RrLL8RoxFxBUD6AZQbNNXvRxl1Zvk8vulSsR1T2zw9RSbVZuUC/eJU29HKFoge8+
AahOCAHbZn9hpWIl4R/cFGwpOn/mfMBBC2Yc+6qYH2G4buzPwXoIhU/F+JZWHcrL
MpRYP/mvz5QLZf62axHDh3jcH/EpGKNWRu43pieE+fsZF1EsFj5V3krXMYj6xSeg
zZcdISSc37sdpyZ0j+xbg1FQQAASDtR0Y0PBvliIkckq7OJdW5pnLZnTS/J6t7pM
zuctTWcKlJzhYiTqBQ9LwK/DeHiIGue3LOfV0xUqSqyKMlqrnmAiyD+d1ykD1IQL
f4mL/TeRTRg2EI/lOZ70cX/w/fkNZoOwum51xDWuY7cmZ4XLy2y5udmOnjcKM0lN
Lwqi0waj17eNleNVxs1nwOp1D8dbApkMJmQo73EADgJLD9/ztq3q4tgx8DEEBfan
1vByNk7xYJOM6hMpZ6W0ctXFySsQJYQWenFKljHS2JMcx40uTq3DbMnQtOkbTmso
WnhtQ8c8HnBdzZPnMUsk5grX1u4fgf+Dj1C8qei3fdAkAQiIFcgx0OKWaB+TFUPP
c9A1NtTqJvl4yCAbeHZOj24Pr4ZrwOChEUgRIXsv9CL4kS4ZkG4A8DzyF1D4VxLd
bI2k7+jYEoC48VIUFk8evcR5rsm5s2SNpTuqDjvYsEMVj1NAiCdFrjhN/1Tw/JWH
o99hCUkSfhFlO1xvBL2bSy4AQ5FlkSZtS/ULIUWlI0c0GlpCQGtVQcIqmaVak/NT
8Wj8q2Xz46B61Kwf4kdB2BzCtwu6VwxLq153Ql4OxlB6yvuUaNgiPGVr5aWTV0rc
Vf9Txg/qLUQrdilh2wviIIZm1s1828r4xMq9K/FifsnENzbRP/F3ethGrMMleu7K
mhe20UFuTrjE1kT9bXa+rI9O0WV4Hi7wXv6CMNnWXst1AVGQiSQ+hOlQN4sJfPj2
jYR7kTr6RAeyFj3yVvZhNfh/YA9tX/CzRt+TZ2ZldtrpqEL/AMxkumSMXatt+D+d
dYfU2x8JOLAqijeHyeulq9lQfw++HjM7ZUdD6TrWvgOPoz7dtego+p75A4m0ScFi
PwLjsPlw5d1cDmYHQ+ZBDALHJvbVsaDk6ABsFZioDOfEnM7aAEFgIcp4E0Ps48Ex
f2AzkrrVaczVSHfwgOScZYPJk6tGce3suBzPNOKa2nIBDSG0INHE8udZkc/DB9IY
KoHLLteYaQYI+vGM/ulqUInNfxY2GPJgZAGW62dbYtj+7LloXc7mMBq+BB5oi3iL
vEmXwv/H0R9PVIHD2cVvytsP9CLJrJPaszzT4BtfdsE1gjbqaB931W7MSlCUbMwc
FgnhcGP55Rb2uUCkO2Q5mTS24Bwpk+/49sX+/6pbEp9oG/vdoAXRdycdw8m2qcbq
E3EtmbkzHyYXEWH9IbclchGev8z6WjUzZGVM51XVjeJj3grCHvo3Wm/UvOUQkK+r
5MioxAz9j5vK8EKifRSiX1+zo5W0yc/q5vmkR5MeH8B5MVYp25erSytSwGxAuttE
PvvoIvbyrxnOs6FutQ+HI3WWK9If4iVdMsiZtEfxBmEQFilySq2G/W85I1aVsTMC
kQMQZ1OG9Fm5TNQru+y0+2sYpPaTItpDo2paRNBg1tVGa6oRGvhJQSS3DEMPBzd2
2wqBeNutf6X8T529k9hDyYu6qvQm7IdumrQcFjVxsHAXfujemyd73rBOs9nOGgCL
QtuCu8I8tR2qMbUyA5Baftky73FPxnapWVeZRrTKATGewIprQZsWYOaF2yB4Vbi0
oxoyekJVZaiitM4bt/nIL3J8HiP8VvW5IrJaPWmelP3/QkKCY7PWtfIptgoQ5aNM
8zI/+Xmdu+FlDplapi37S8aeaCSe4KO9NyBuOieegSdu4v3P2supAIzzsG5u4QNz
4rnwbvpaCVlK/pNA/uhS9SudaDRF5D0NVWzwmSupIRu/JvkDl6unnGIWIevoy5HS
ne1pA+ABBfsvwFsUATmDGwQHDabkzhGbEWxFiM8LNsMGgCWfX12LNFbFmHYf/fJ0
TVsuPpB7AE8ahEipHDPTPwoOF1JbB1QWj8VZrU2oEZYGew7E2KHNUJHWROwRezaw
2uUS0I1oGt9ByTfdEi5GkPlPrTTK1pBtXTXczpwf4AO1My0us+GS9QPsu42EJCrf
Jgprz102NcIc8CQK6uey1gAIXLhPCsDhCH9eA6N3Avz4ZMK7SWDXibh0vF7J9uB6
+w6V6SjzHG65hGr2yngdf6TbQjDsX2QyIDYpvFAfMmos3Bw9pWIwBXLE3cxrPtkL
wW8ACo79YtuG4CveHpaTDQxPVHLxwdv6JsbS2BYHrWA/qm16EoBJiJV+lWSFuUzV
s6dh3dKuJOLbVrtUhXeetxr4NLFS1TPqi0qw1SJ0TBTRaJaqdTFAosN7fFncqkwG
QSQTwtmdrMvBeWGXQ/hZQyINQyUf6WUuOjS4qKJhLS0Lv/FjLEueMciFjsvJGRa/
uiZZV30Vr+YiK5DCVX50TAaKLzBw6/8s7esvS4/uAf8gra9i3XEMdndUwIo7wA3L
6Ei+73EBUdCt/Qw4n9gEZ0haWL93foc5PPa98D1LZaNYWL8a/6Vp5P/KXoCmk+7L
SRI6u/2Lja80Wee1ALyt5BHJRpGFm8lLsJIDvlVZwFPRsi6L+19d94iCO+ASjRWz
apcBpFmvXEOJ5gRH5sj5leIxXLvyxrQA+Exj12dof9X5Cu1jwjj66XY4LmNZdpIu
UwZP41r+/rT8e0p/JB/1Rib4xuN4mbO7MAxU+74JYRKV/30TL1h6Z+oSsHax3SBx
3KeKaRjcTgG4GtE7c+SHwitC6EG9Pm0DkXxRHdZJmrDqCuZjoYgxRMvuHJ/sRkcU
6kM6cHYRhD7X4YS50QmgVIADyTNr4ZmK5YlZMZw0ma//Wmsfj48wyWGAFUHl3FUY
HXT3+glrrBb/BjVLzKd2+FpDFwhVcAOog4hCGYbK3TpqGD6BpbPLRCvazytUzVuZ
JNs4P/IsX4lXe/zZRA+wXxs800EXHczfoNQwfFuNzO2cW2tRL2c+17sEr9jW7lHU
nKF5cBM+BW6oLMF4jMfk8gQ2JZpI/N09NUBz0jHiHT11rSH5cIv0ViUE2kMyz3aA
6h2lHHDQu5Up4ODsUMqcnDJzYwUaAxPn8SOXq2/GnF/yfwsaAVxMBZ0B1G3a3/44
iGrmCfjYI7MuPDTjnyAU4xyKPAMwP9fp/MePt5NoW8LpKEVcimJ+kJjgBs7rIsjA
hdhlVvkrnw3UZ8lMrdq3bAB4JXJFMA5hsDU2c3mOMvzNGtSGGQ3SthUaJXqDJLej
HkgGPnWFJyr2PUR6m6VKzIK9bdXWsBmBYHKRQSlHKVzbGPGo1w6jLHJk1ykcrhf9
jjV5S+8JGJXh1tNn42S5/oiuml1LymSVBeYpGYDF4zV6SVvicaSLk/FfmmxbN1ID
1Nd36HOa6AY5ZQflwUdtSrWbge3p6904mdxr4ytYGtYyLhZ7cQOf5C/87BrSYj3N
+t9cTEuPF5jMj+/e0xessfsQRlYdF91fDXnUNbV6PUOZ3u0699fmOH+vQe3KzS+o
vJKUjIRaAj8zEZbvzAA7U0xsBoLkcaOjsVJkj+CIAA72TVnFwDI/imxXPl/ipegV
rXJ1gGR8toHTA06oh+21sr+HP5mlhNlAROqZ51DNiSR6klxd4B0tfnmePjuLEhW3
igErP1TU6BxeL9R8bOj6WlyufqSCFrcinf1Bc2bMekItHkoSVEtr3tx/amvEJzI7
cM1ukHb3LMdgieP/7kw4TaQKzuyD1IptBTHkrhKC/oCDZRQhcRZAS8CRdxmeAvRK
Uo7gLHp/+ri4AtmECUJxTNUx9AgYPgjuhcUHT9I50zRKc/0Q9QySku8nLpBdMmzW
wcwwXphKNpB36VSp0f5VbdBgR04u/VupSMgLjkkikCa0OPof9R066/5RRLHCrPi0
oeu43kqMWh7HnqSSNinvye7p7sN7Wd/DVZlB5NBwDbu3TfHmGiK9cSAnNTXHxdrJ
0rPuFy2JWMl4F2GzTyAsIrEKi8vrqY1eFre6t4riFaH83EdkpLYyzB93cFEOBRqC
wNSmxFg+kJ7onGCe3ZNUhFrzIVZ2d8JpdRuGmMoJePL/2Oh2715mX9Gib5xbFTdR
y0egd8QQtObeM2a9vBD2V88XeZSZ5DgoMJcP9JygoT5qlWRbLrQsF45EC1VokKS4
GgbH0mh2bEMxtXv8RGSsF5epjiWZl3U4Q0c39lI9Nl5IiB5qFucTEJ3K2rO/fQy7
oMb2/FXm/erSfFGNh+GIcUSkvvj0KUFXvYQerFkmwNe50BxCmDG557fFcVLOXfkS
yrVRh/SaSxDVbh/aY9K6hTU43PZJELuIiPSgdEm5THyHkfp5lMLCklQFpYaFm/RY
RI7jBTABZkR9L96OpWs06T7Jaq7Y/L4STrFszd8HwIGEOZ4jJKm1zg1P0venMbFN
GmE1F6NloBX2wyLH7aBiVmoPNrnxEdfPNTEbmdE039jAIWKEi37TwN/WH+KijD73
QSXX58NrcxQTihhf8MfetfcW6dAAIx+DImFIYykvJKX57NPNfBPbdN1nwd15wdgI
UCGTF5ytC2by+iSV1PA0zjeBGDeBrd4jQlhia63UDABxNLj8x8mBcJ1opMqUk+HO
gRpu6y+OxJMo4je1qPjpMVZVN95/lOWbZC8C0Yrl7iQKu0Stu59S85UH97x/CrZv
A5ufELcyIUKh+kw7dGQlz5ChXu5dLrjVyYIujtD3vErWwPCMmUlrpemMt6ynEuii
dci6Qaju+S4oZHOo6nmUJ7uxhIEd3CshZchM7+7pwEqJlPdrv7Y9+9E+PzI3oFmB
i7TcC0UGOt8r/AuFBi1xpGj3pPQgLTLEPYxIG6n1wa2YvBcHJO4XsdzH3duwSQh8
1L9ukrqKY54i//gjPYsgjaCPrNx7Mvz81Ep9EhD8yscxX5hRxFJif+uNMW0pV+PV
3PlOYr/zwVwr6mMnqU0HDVr5Q+ECZ3QxqLZGx93e9Bm01oNuIRdQdgdsdiiWuUKZ
+DLVIGWSDq3cUzvRz7cgWlHSkg8v8xnPYNOwAwUxEsutfygdOtID3INqThwrrwaz
lbZYT6q2Rum4ElQLhQ68i086hwOvfeqkJQGBlptBftHN9NmLo45RT89ul2+SPu1G
M6w/Hinpu/uAh5vx7Z+77ANEDBauyUPgTmABL1Mun4fvqa/LNaHIHZdJrLAlideE
Qdt4EPO/ACsBh06VkSLLwC/oVnIlPnWcHTacyWAdCwPpyUmAvu+YWkAjKXJWcLRc
kVhR9poNa4224IAbQtutxKpDMnJUxorlaA9P6A4evXoDQICF0XjEW1w5aYDQ3TJI
E0Wr2Hh6SSpliv6Elq4Ciuc+41Zgb5AZEHXahRKQCX55lVq/S5dqk02Afafkrj1/
KooVJLplVx3lx+kqVm5aRcFLPx5p3vXGUtvCamjjAYD0wNcp79uOku1+6CzOJEK4
v1a4egGpTk20NxXmIM66WdlSN4boe86IrxiOrz7/gEdhse7rtYUqxV8fIusThSQy
ZDfl91I0qXTkjAXPNDXDjGRugWg6UbQI02AHwwz6kScscGbMXz5HKGXOtSq9KMhU
U4G6oeDeirjIiWEbM+tGsvgpR7ktva8S02AIB9btvGQx5y9zeqewbjvvxsr2R8EJ
l0uXtPtoX6SUhMNeTIp1IUWdn8StqvGVwBVz5EfRVvgrA+7d2tZsu18hZnASvVta
Vba1Q6g0Pq/C7d8867u8wdIntX8s7kcWeBXsOQGgc0DAFMlhUaF2Jhhwdb13EV34
w/UWdx3udj0eZTR1VsywS4fhQNAhorFp0XWmTFaJXIfBKjgsfKIjBhVZCtu+K9i3
WBplVByrn4U0UWfDqC9u4vzSGc+PWp7ewz7VgCdTlH93jDcT6VQ2tI2NYg/OK8os
2TyIPlYoAF+vY/N2SWNb6oTn4P8cGTK9PzRIBx/7EKXqICKYMtYZy3gU0CA6S6Uf
BX1bfhN3gpxJVgLDvcCLaHOMc1JlFbIXXaPZzTN+vcEBN7Zq8jzQvJe4sw42JNzl
kB1I0KVJyfggI/SNHkDU0dzfwOGBnZptG5K3SsLhSbf+rUnVPr8/drKlVKX/5qJY
XzGuRPvfirbUCvJerO9KTlQeIVpj4qEVXVPyy1meGdycYh7inxtwUxM/BAdd+H3a
T2yddJ+W5pqhciB+WEagOfT5DNjYsKl8t0YaqzF5U7PVB2jku52wHhe8FoIP1PgM
RpUeqv2JQr7Zo5Oc+afMEiYtZBawlZRqQZ10hugqC8QoL3C9ILMbIyfzMp4mbWSZ
WeEQVfTyNh35cqlgSYYJsoyPW7GX2HrPnXoNpqVLsZHzJfZBpl2s1hBAgR7Jg2HF
Fr+Pygh7wYcMRe2uRBLSYwHrDFnxIyFoE2daMYuVfwp8V5uX5hHJHwh545zh5LBy
TR37ZjNuUH4ig63O8Z9CDkI9F/rb1P5WLdmEVhujC0+U8mZVDHCLPruBxrMqSHQM
UIcn2zweAzXjfRnlvsVtrwseyTb3TGK7CzO9I/Bo8pHJ0XantnH589EXj2Z9UIrX
ZSZXG38xzG1gL8QigTp04AcRTX3wmZMNkgUfCzDoGDbIywKnhTqj8Gcok8TOkF/H
pKHLPK3Q2sBltPl4dVOIBdijKEYt3H1XHmrBrQQYeuG5zFx8Z42GNUylbmS+JPEF
RY6Uv9MwwMYfi3j7ywpKLedxyyuo7zAfm/M7PJMJBRARrGOa9nwPAxNGoODA7qZT
X4dp5q310IAT4HAqzQwgPH2ZOF4aQREXFkiE0TdTehCtInbn3qJDsRKxj1V6hsVq
3LYGUlfCoI4xZI6TLQNy6LLDLOibX7P/fs117XzruBzYUNgwS7OPZmgiARa/RyIU
Q2gAIp5JkfY64HQeuHFcyr1VHtV4r0mZVKNJZ93GdOginyrG4s8X033noNve/c+p
S0BQ/WoevABmL533IcdjL1NvfUadzrORBz8d8BWzOOMzYAH9NSVQ18AIVeeq2eQj
TRNBPBKHRsYbuq49NM4BT+5fTxgbtmrou42BOSXe2KfvgFuL8M7JAHyVB8TeQZBh
z9xXd0j8rmBytwoS0UTbJ+UFOo53J6uU+jecavfqiAZpQlsF6fFvtOYo6VIurpKW
px9goWtS4OAHs6w0gGdXqOmmEkGC1paO3T4BUUpKI84hYkHIESgDHFAK/J4HZVHp
3t9kj8QNaN8vdFBApWVPQz7EhVQRAM4rQeMY/NoQyz4tDWeCBzAYqp8KtBCZVvAC
UdK/RBexrJYtzjN0OOb9vZI162/7nAwhc7HRy+hVi/eEjYialtcP8KIYiDGwpaX4
ELlI8dHuAjJN4Yonj5iWIrvF5Mqts0kC6ieJzwt5ERBNeTkQRPOOnxaFHwhge6Mx
GBjH7niqFc/Zrq8XL1uy2kVgXkQjkbWpV9PgXoFB4DdYabZVIsb4n6hDvQ7dtgKy
4A8JWEAiLhjYkC5XOVhnERRygG4Ix76ki2elyypakXhFGOtNi8qyX+cHku0IgrBq
nt+wRNaFR8lAKP5K9Gje/IrHVOibu8fDstgkU2EKjGxyHGM7Mjdsd7WvKH9d5YFE
teuPuYlM8FM4/qjTZbIWkbKipJ2BiyxOxLd6ENCV81tT7Z4RIuFvDqGTqqTVDFOM
fXghzdlbI0m3p/YUVp9RXjOXALgWuFy3U8nwt4vxAMbVDZL7nq8rC9aKzdA4IRo8
e35+LA/v8kKW9iaAs/jW8I4lEK0doZ6eMcLcy6vl4faQW7qyXCaqYTFGnuxqJPBb
hh43VWi8n0rk5GJxASGpXdYsnNE1y2P3+PyEUHSZVPo5HOBdC6St/6CtTzgFkr+5
Fe8qixbqamJyqkOmjfDHnmN7Q/xEw5cGCiG8t8ku1kOLLpqzOYH5P1wUcmtTdFCG
t9Z+Z4HODQuGUrYk26qJc79E7EMqSLr1HyyT2JN3FEcQdLn+HJUCtbkMpnEPZOtG
MfePAcQQf/PmUfjaWyRDix3k6Kat8sWsEv4o6p0qeoJyhpYma1cioo4mv4cIBnQA
ErDR3cJq0FQwTP+5nPawm3+P2EQm3FIz29I+7j/jXeB/h7Z0hY7PKdb8PXD8RcX+
sm/cqvnlua2c0ICXUJDic11YrCjRwfV6hskekauC8y1BBe/yzS1GZJjzYJT5FSfx
Fl0zeNcq9wRzr8vjTp+1IiDb/6mm0IsEFdnmgZgzaD61h0vfGH+Z0OOLuvwCQkmZ
ac0QhJKOfm9pFPyK1moqKbAcGfjKuyS5bNAO+nyl/tYxDx9HSffHd086G9CQgYgg
GF8iFqkIqyZ+D7U6RwW+XEiT9wM5VpVvtefZbq+mD6K95/rZLG6r7F06jybKi2Nc
1IwHxM4+3lKXFjFBQErLVuyzU/CUwuVbyU+eueVmDgEpiYugCGcBn6559RJ+s4XI
sxDIXR/VSzR5ldXVPMZVzdHkTE1FIXMuQ1ot1eUD00rCQDSlKKRGHNFAt7kx0Qs9
nzkQMFwjtA6IyYfmiuo2uuetuKplWdzMHhG8+UeJHw9VpkMvc8fbJkFuEays3Zfu
txCfr+S5vVmpGWlfSXOb6bPGzFcrMogxSQKfQz8bPY5nQ9cwyiR7d7jtNPe4XPm0
yGJD3PiF2nX0qz+MV7ifyRktUbyc5H6ne5YVBxqBxNBhMD541HpXwhtWNe3BWw8U
Gl2akUS/ekOQHS+8nTqjrtQf/VL/0majJkqxYmkLGszaX/07inZ9s27Hjjcm9fMx
nAnM7LlzHeXN7bKslUjEp0Lt/eJ0KWpAaGroa7mmYKZKhsvPvKQv6+Ta1nxe0Nu0
pPWIPWwCS25dU6CFyM5K8Zwe+xu9IoS757VyaSoObe6zZkLEwj/JsVLw0Psl8XX2
frletVBCIsqbC7p5XcKaF/n6bZ7S3YUBJctQXH0rV33cJWOfZ5ZyudGkbIaq4dsE
+u0pFM9bhg7QbrTbMV9JbQUzdisMvSWeiccgajLd67qjSpWgKRyt36nRRnsMwP5m
ETYP+J1ZaG81D1fonubdT4yZXHjRwHhEpnIKpRyMx5C/4n0CVGXdqPbrgDRaa3eT
yWpkrxvvHcfo+0keg6gAm3P6VBI8d3/e2PVT9kB1gz5HdlAP02pJ8/QhTxlQEnYd
QKQiIuBWt8TXbbZDhnF9ra7fW5lB8K/zSc3gs87Umopd+pR88znvaKN2yVd83rHm
dDWRMLpXaEfq+hawAeF29+N7mS38+Ox4VAvxHqdqv2rwPj5WNeu2ed4KRubS3Jww
7dHya7nqvmp8DmdDqoqOLE9+JrM/A/u9pmbibIyDEXmuwmBvxy2Z0kGXhno2jGM3
Y59fc8nsWkTokkZ23UxP+Q6bpBOA/u/VpwI05In6dL7LFvfG5HUVgchwoS8QB6+q
XIe7BWF1q4mEbf5ah9SipYQhBYCU/qpAC4z0sPou9l427/n9yU4otGaJVU643ZGc
dohlRqp8W5AlT3y93RtkxNaboUAWxg+ub4UHCe6H4E7JX+uKQEBAfY2x0w/Tg2W5
rrMe6pAW7xnmw5PhzmJ4u3suCceXMJfnnTdVzsm+iiT/WdulcPY+IhpSrSnw1VFv
kK1Q+RoW7UkRgDGn6J3xNbSCFnmoH8pwscIDsGDcN62T41j1YTi0Bg77p7giTzjB
zuKaQph0LhFf8Dc5H69mTj61ApgSDkxRKFrFG7guYRq0A1iB3a4+ldKsqaNMkIua
dh2i0TDEC0nV/5qiOrf+YDbJpkNrK/pYPEZt3p9iP+cmaqEvJUIgfqOQ6OlCwEDx
Il2TT+ZyXQrV79eLCz24WmTwjRvpN9q0mE1nEBz3ucCqoUF65zW22kEq29kcp38o
tcfgYaLyZThOTgzG6LWkVh+27F9DjZr3cDuO6Nfsx22/YMBl+5NWFGP5QRBgez4q
JbD9KoNZobSBEe5pvN1CNUQufhGPnUp+TDOZ+CihkATrudtO4W0xS4qNbX6y98Kg
rp5demYR38yRcrPC5Qmojorh2Bxtk/xR7kHbwxhwosDbUq7jse3CX/waZymXRwNw
y+GGX0YDTvq+XQg7cPcTFtcjHdUEyH44Gg+rQNZ4/z523izD8+UfjYGJwLKg7EjC
qlzHbMJTiGLXOmr1Ge67a+lGuioxejkdmBK5SKlGviimxPBYqx9fUCaWpKFE/Kf8
COD84fZCQC+wjX/G07EflzmR7XUYsyuwW7jqHBgguZe9Xi4z0umlprzVavZuYmCH
M1N34QCJ9xdSLF9nCxIkZ4jb5AVV1dxA8FCZBROe8cfjhpfEGfwKC0Ez8b1dnn4o
3O8Byluk13BDtTgFqkI4ctKlhYiiIu+R1KXtPhSjW+7Ng3ie23DWlRLf9a2Yl4pE
hKADhwOjudasKTLSu7lsDToeo2BpJ697JMo53NvLB/QquQAzC0yr53BsLGzNHH/8
7K/HzCsnGaft8dQ1WQbQKj94nqhGLhRAtjzhLEIpUNQBP5YvJMv9R90u/owRu8DD
DNoPzwdCrC8Ibp8KzabBt9RYhu/R4aTSVL2lqOjLGpwr3O7vp+IBwq3zTkkKZvG/
IzngfyeKRvNJhhPvTQBKc7KASIJnoQR0n+TGHRySS/pjGCDnkgDoQZohJXy2iz5w
a953R6zbEPIY/WKbGOIezy70za6DeMOrimZzakrDF7D07nd9XUo12zoORVlmqSl5
QITTs6vIA529NHRDE13v/VQnjDdfAlk/4Bx7j21OTM8lLcfQMnM5v0mqjdemnBu7
ZxrQYCaDgj1M7O7GIfTB7RMltnoxTD2KgAXVpSa8OQZdkfqapBzk+1F1PStntb7+
g+rNx7+zdjCoXSG6QixWnZO4HMS4Cl37iy2cjuwbLNhoMkHl7mOvnpTPRvohNEGo
0AEhLQbxecJBY+j+V1MO4IrUPAS4bnI7YZhT633vss6jmKkCa5svgr7DyJfXosRO
dP1uMbOLW/NOWdWibHyFcPQDd0rJfVtWi3JDnCiYFPYhYvtgb14jTRChgnvyRCaK
EbJF4rnTsPwhgA/ZH/RDxSqb0awIygutHyx3nDpgbrk4gM2u1x/w7wKojDzHivcB
Lp0Rm7HlOFnrUsg9a6LmgrKfoUBBJ5RRJ8oxy0qX4JUIyktPZ+a8KeseZjQmlync
OwoiGKVQ5pL0r/CqpEhG8IAbNqBvFhomnSOR8B0wFOCvx12FoKwKt8CqLiMjyzn1
uxIH9MjQb9f9TOjpnuj1o263VUf6l5TTvxtJuRmbYcxfZiwavvUEGTZHcs59cD5p
1WUIwYMaltIZk3vscDBk/TvjNCKSkZoaVkM8Ow03z/3z7Vt5Hv9JKqyy5CmJOtBt
UcoEI2teXqOg8xJdyuQLDh2hGrJWQ/Ehpx1Zc4DkknecSrAP7vIN6mCqGNZ5ozOB
X+dBN2BrMNwoiEX9A1A38vo+E/CySNFNWSNioUVsPMqP3fi5eODLKNsYuVop9Czx
UgIQcHY27L2cgVoQujpOiUj8j0Lmv0ja7S8LiX20LhfBTgCgHUccwdCyULcE9Zlh
gFsC/jPTjJuEjOu5GJ9CQFT0cK68/Vlm86GuBx9BG3aU7T7N+0rmIloPHXnypFk/
VoTkP7FZ2D4mYEiR0FxawAsBKZWE9ZX0+OS7gh/czpR+6WOpvlJn/PgGqWJ/q13/
LadfTJR+sQcw9cHpAa2mh/3v1fLxh2Lsr8IUXkSTHMdbfeMra5NQAXMvc2zs/QI5
LY4OaLk4JAivncbr6I13MP+CkSkNan7MqjMtz6OIB5diAVE4/SCzEwXPeQo0qNeB
gTfcvW5Qyu9yye/EUlRpZRB+8k3CLdVZqYnqV+BTv9+c+Gc9Om2WWkSwS5jxATO1
GPO6ycvDLgg3eMQr+WWS729YVuwYHRu1mU9qOGNnsEQyYAZeMS+SjP/uuS6pPZ/z
1r9GBD1zjXHc+K5aXxAk5O/keonfc4C5tB9aQb/bHj4qkuqiJVZxCTTJyJChD9Nm
dDi/Fkxbfpvqdc9uFoImW/IQ+4ofGr0+LRenKymNLlMYYcxzKoCbQfAvraSXfTte
iUmH4J1r45mVfyXz+uz2AVHAJF0CfJD5SEak/3PThg4bbMH58QIj7w+G8B9y/rhj
rqAQJ0aXKZunkPZGwOU8A4kDgCYGEoQnLz/LntpKszl5gs4P0g0GXPlm3gbZxoEi
dFPXdpceBuhnVGhKJ3MS2kX0JXpVSqtPOvGc8ZlS3lHghLY3weydSp1Oya1tcQL0
gMnthFlOP6FPO3GLEMQ9lgXc2KPeQl7K6hFMo2d6wLnS/lZbgX/VuazhWR/D7Fxm
31AMqvl7t+qEk3foQV8uT0PtvcvpvQa8Ovv9p7k2GEMeDhw45a7bl/7ujT7jl28C
ZrR7kcUJUkSHSqlcapfOXE92QOg0lzam3+TIUzIBHAa15q7XNSTNYksbihbWEn+p
OmUbt+VlZQGgyuI75o2dM45BzzoDXBBzHRcrQsWVLdG2d9SSo6GMpkdcsccdVYYl
Go7mlZOCm1qncUo+iHbovxe1DF4xC2+oZF2C625WCRFe45TE4RCwrXM57wtx9MeX
L4xxUdLkd92LttrfjD+QRD5JnGP6rjfyFz23Hfi0E5c+pd6ZueZEAcce1x7d6wDs
1fNLceUdl4MeBbfn4gffTH9NyWnY6zBSUQU31KBCR4t/FIBYocotz7Ykw3rA3WaH
aSoZGmObjSGHqRaieUJnRo1q/JFFCJ7nxuu6cy9XVm0IeSOAr+FEN134qp+QeSZd
03g24EbW01ypdCyrD2CjMFLTKhJgxBeAczczTtbhq4hlDwp3Qi3F0L2D0lrCvW4y
pqMCUZujaqQ4OacoK8R2sdROJpcsGxH04LonU2KLxK9lBML3mAQ5I3/ADk3bzqUi
y5oZzuvxeAjEUuQrxv+mbNA6zo8jMaqU+uSjMi6m75D+UqgQVbMLpnsW2bxF3L7U
r9Rc63F+V7bF8H8w1UrALCGoD1sQm+V1sOD9PiioGdJR4G8lj6/dsu7U0TROdzf4
NQ6JJS5R6tamUGm0P+FelpwX0ATgULDpECPtqaDv2fKL3gbP0dt4NqMLAkI8tqQ1
NhvMppcTGAhvs3syR2H5CF1QX2PtTN27BtF/ZTE2qmFhaNMMkfING2mfqKR4ngYR
Dc6i5GO4jjib8rDo7jeJ/hjTpodhtWVCAgFIzVr8r1xcjgt3etvm4TiHDH9JJT+p
qCmZszAOEPof8gL6kPZTHp+VRttj5J4GpQ/9B7aRaCmwJMGRNnbg5ULzr7McjoKo
gzfhCFTN8NIAyLQGummt64FmIzrL6TgIs4E6G5VAQvYq9ZX8I00saG7Uotcm8jRE
2x8Ruev3vQ6gQvybskR9gsi5vmRt6Ly9WDRpUheyirgFSk1nUZA4dzrsIgNmBhCF
IwLgeTU0RtwpuOoajKL4bShwxyNvuQrAGGboqKjooZftudzboYKZKnwGnJzwzKTA
lERSQwH5toCsPAYSz81lOiDQ3hn2Ae4EttUESl08BmbSKqUi2JvFL9F9fzzzfVLD
NajUmaNBXy9qFuw5m2OScNSUuFdmqDcBXdmtAGd88zPXj7MxI2slF2viorH+dT8t
T93hD/tvT/ZSB9/ofXFDj1q5xxfOAn2SMgzkN55x53PFWUC2nCHB5Sq7f7pv+7Vh
ET/3xMYNAW4Nv6rVDhNYKlcvA+5KQzoP0xlwyPRVMWr6wbdkxGbPWM8mehUh2DBj
8x1m3dsawP2I7CGljRgNH1JQyEmgRPyN6dI+DavCFdZYCPCBM6ktXHf0bsN5tHCT
OD5nJaVkoXsJzZrppLH8P3hh/c6atMLclo60Bk1aG32Y2XlYk7bdfDP3V7xl1wWD
6OeD1DKELkLtSCFzkgZHPJEwZUNa60hYVDjLYw0eKYHViBFRVujobMkQnzStC991
HIknK3Lz1lGgLdvvNkG6Rvof/yth0nm4HrVhiTb5Z7xi5vsJNv25AN+mT65sgtn1
pVib6/+dF5n0BkyIAbxppEeAgC9Ln2omj3DYE8QyUu7687tvlllnp+sWK4Q3/Svv
NwIkZ5S4P4lA84DuosN774PtGIJZC5QTvVn/VPMy6hZDup2r00lv/089rFwzhZgq
GsfqO3RZOJyjuHNjBUu/4IbHKUT+undYRj7Ysnho0rzEKi79okNqJ5maWBTgiW3V
RZQCsIEzA3vrYZ2Eokz+W9e+bgQtFyqPZ9P6Wv3+XLf4JEkoKxWQ4+5xro2TxwNM
aQgGU8+d4HL2rL2ydlhFXpuc6us+H/rOvvcle/JMsewNNP1mNYJQxMy5UlrcfIOa
oEJcSWyOjplPRSOL4/VCPRE6sOwlIAf2p3KLPGTvf/7laZ5wyVKsGtplGLm6QwLP
vFHW35Cnp2Eig/7G/QlUUlAmKNm+++MnbxnueFfyl3KC7ZqVtaFWmqWfZ2ArbYDM
Vya9OHhaXn4pNxIMJ83+34e80x5S2Le2HTEWOiaCAIpLQBR0uEBfmNENE2SvO2Sd
OXYRK0xTGtPfhSkFnqL40s2XYiGUuwfWEIWwL8Bqu8IPXXJe1btgHI76AzPKeixN
6tUOB3G+fHv1tP54MGVa7UVOgOd1qPnMhgkHKwbgdDbRUnGPBXhcMvNbo97BU4Ey
Nbzf/JlU20Frvzod/lECLyjBbjGoAVO1dx/mDaLmnHgJnUM9tQxj4DxRXsXsLQat
oizTT4CZIuQxBSwdZKT5+huLl0za/HS7rV65CjNEpSb06Yr8JAwSfUp3G7DR50jy
OPU3cIDV9ED3b4lSjZdQo6t+JnblFd05GHy1RHD1tIeTtbgry8hHf+y+vfmoXsml
jsDMsAPdsWWEcwocW+oBRiaA5a/olAt6NGPzonQ6mTHd7yKh9mLW44vvZEIBsDrf
YCMwipl4UAt3p+KSWLMwRmBemnpuoPAGuiXE7TtJHoJlR8ON1pw4aGFyLGpNnVOK
/5MtHjHBM9eZOfbybsvZbOHNa1gZx0lYLMM234tfWuJNOzLDL9GTYwTK25gRkntz
2RgDEPaR/B2p+fTSLWZrvU3nMwA3en1jkm9hIPhxG5wTBSa+Aj94GNtMAy9Iuwjq
5D/lm403Hres862IZEDUMQC7pkSy+C2DslMsRfpe0zXjsBRTcOTTpzWCjqhdnm/K
+fM5ZGKi/9yWZtNK/FpYAHq/mTmxYCoWmZ2nBgB/oMvW5ERNs4OJcb+iQAlzJ40I
40Gfoz+GFozxLaoGeqTxTzT3gVyRy7KfyPwAdKJN2FLPEOZgsyjuG4+ZZmgVU8UC
dhOJlxETY9KbQRP82Vkdc1wIOzE+doxRtE792yvvsdrTdorNr3KYgaAmvPpi/qLD
NDXA+PjxLnCukXHkTTgdm1nt/zUTmGGzsT220z05mNWS8yC9gO6qCY7ZxRLgeXkY
E7XrTynjrpobiYKALgegDqz5lBvh7Sorn7TaC7MoR38UVuSpOmzGJpjTR2sd8VcM
PQPiJXBKG1d+I3bVYUC775P8UIw4MV7lPligW69qQMmxvTEIP8Z1+rUtltbJguFw
Nz7I9YHoJsVPHFi8NLqd7ZNpURaopbIqRExk38yVsUMxGHo29fJhn+wAmozItp+6
/ihnH7vtRcxGIuQ6YCYZAsrYQo8OOmVRh5RBz36jY32j7WtX7lVJR8fRSrp6U+XG
48Dox6dVlVOIJ3dXKWbXMutYa/3lelNpG3hX3ebH4yxCv/XyiX/qV6tJUj7EUtsJ
iGRqBiYNUp01URbEqKESy9rJYahCyF2FRWDUAZWXnclwdZLcXzPwug1nNt0vZGOX
LB6uLAaqQAExAsp8plhij++LFWb0Ta4Uj58QzHVsfukC3FUzHX6dZ+ehZ2X9ohoj
B4pKHgaja42HVyey5vPKtRLVXeDDNmxSknRlJT4GVjt9M6+pgQOORnNuTY3tLt7w
6aO9XNoxpHne4B82XKtNY59CJWsPGlNPmtYC/0K6oXI2LcMBWJkbyIB7o0NTaZMO
z1t/NYm4uuS+GztyXgVAa/oHyvy9m7NfnU/TBPDjimczzh+FLx3GZu1kVhSFE9+B
u5qO594L4XuEt2tl+hi4XHU4XulOtrIs/lHfRZHyOBEGAhgCMXr9EY/XXrP3VY4V
EgYhtFZhbGkRP5F4CGb3cyhetA1YVOrXF9dWZ2kR4C/yqhCJqoEdA+3X1G01jY2j
bSz3lUxNfeK2rhUZt9H2nvQfXEHI4LHFBCkGfK5xOMLMb2FzV81ufjxx5NGg9T73
JRD2sTAHJuxqTY9sW0BfrupvrBKlbkfUczqdN0VZJJ1M7R+MFCyW2WMERdSy2acB
8yUiUuTQ+Z+FQ0906MIUdMbMFsnHPnFw63xsFII8+dXXGd4MG+yd54eCQifoI9OV
Sr6FZCzs30pq3RfU6JhRdkRSdyXfIkXJPfHc+WodOvge6TamKpQf4KbwIpbppCgD
9lcVm2UAGUpJdBnM4Bc8SmWv5iBPD26VpV3fOTMjuFGNwEylNsweOWgbsCe8Fa8D
7b2/vp4X5EF6wGDe+/wscEPxbpmnqmiZvxwmKBt1uWR34oAVV3FC8c9rkcahxL69
eTv4m31qnMDlBEiwdHzPT5olLGo9AQ/ZbrHUYWjXmctGE2JYvzqvR2yO5lQDbn6L
uy+V8je9v8p12m6EMD0V+1mL7vEFelvBtMflOwvtmwnob7RcBET3WNDmK6szUpHG
r/ZXW5AqFI8krSVayIMPM0Y5inHs8bXSR3GmbXXk8CcCTMqAT4AH/UjWjC0hrpAr
EJYMNKB9wMiJlVP4AwCwDAqlEi6zeg4R+mvhbunNWzAYtsrQrEXloCAcf6TwbbUM
VcuiFOW/O8rcgcEE99+N+taenItDD9/+SU3S9vQvbyTFu/IUC11AbAw11j83l71K
+SyGD8O32ghbIqjlzchyVaAt58k69CZNnT+LCpj4ohkSl7wDLcZSpSD6UG2Yx7Lr
Wrd/RdOTlj5GSaGAgg2YOmsN7d/UhB/7Lzjmo2ZzZjn1Hz0CJNPhzz1SVM7kfuIu
LiQCzIsL8PgKiyuevpkElWz8GqsWmDvZHrVc2EmJtt7DIizTSomSXidfGEnbPvRm
gBsG8GK/b5hqK3nbytd4Ad7t8lVtO5kGLefJTvqwHSEx9rcFqAJ83aIdpCpIM6+B
fea104M33frFo5ds8BxjvpO07MJN/zMUAQMnazDXaKk3r0XXSVcCKLEW6hf7b9mH
q1bvVpbSxLanPC6hmUl8FALeUbybSJ+fkibw9eFmkwSJRrJv8x7FC57l4JHwoCsj
TATZdPn52oxVrYw6OidaPyy0U7/WMfLOTZQME+ofqsxqpmFRHVymvxfJxH8ylqSZ
Ita9x2tiugseyR6Sr+FooRG0DLOmjrTrOAYRYtp9hXcyfUzCYQikOwZtIlRQOqjO
mPXLP7L//NiYuzL5VHvcnn872Zkm6t/bmcJbZ0JU6BbaB56TVZdvabMq0VRVHCa2
MZHP3B2tU81ZP7yLvSzxS9eCvMNe8a/h1i+F+WrefOsUIwZBaHFqgQlmIM5U5BsG
t4YESx59b6EebPy5uHFzEuhnwaPKpzUmMpW+dtynEN0RKyXZbAm4Kj/EIDzkLxk2
daZh9jZMqpSBxOVqhzrRf/Jd/8hyCCfywgpebS+NAl8ua5udBVVsA3ZFkJ4SKOpf
5rZeBoLj0H7588cHVrdIfJib7cPMEw8tjbHh0vRl0aYfcS1ZiAPbtKn4/5l9gri/
EeZOLcMsdGIAJO1+TgeCPvnTm0vFZngP30OYa6U/7ptBugRlJXoGgKR7OWiMnard
GZgSxfGsmldJcSTNNCG1NXDmNI2ss3ehAjJE9XKSIfrDfv9WLs35tv/ARaxNzUSJ
/rRoFxkPT/gGNCvGX0wbuQ==
`protect END_PROTECTED
