`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwyVR+S0OIdXJiuF2ddsfDUNZFaMtCtX2MfgrLYxtBTFIs1v8pUvb5BKqcXM3Osq
bBaIINRpxCP5Fl5l/yR8jL98g95If6QMa+DNssmq0mncVzLVhpgh71fAR8Oa/nh7
A3SHE1RryrffsyL0mwFUiF/pVrqGTlmn7gbtXVjTlxCi4wg7U0CpHobNfbqKLVg/
FvZIV2/S9jeBQf6NeqdAv88gZydB120Rx785Ri+/FPKBLZ92gopDuidH4ngknNlQ
ix51ess2/EwrdO3/RDrJB/6AAuXS0LWpHO4bXbSJGIzOEqazAgFs5Fh3Hl7n6S99
M3UnVxICq3vluX+K0nqstWydi3uPRlRuxfZk+Gp70MN2xd6n3R/2hvGKrRdiaq1i
l1bQZmY3dgZsXnzJihHFd7F5k7jwuuujqtDPgzyU204UrvKpO5zW8pAovTm0laeu
g5QFDcoTI2O2ojBpgTpUTnUgBGBUlBY89yj1OqbNTgRQrfCpbn/oJDbkFX8id9ty
2Ze2ydhSFK0L6EIsFVCHfffIVXQkLDFmrpAHQL7WRnpuFYGdVkezdPrO0yw7qzn1
zaioBd26sYKrQZdSH1ljspFeil+kUPZmKFQ/Zq/1KhY5zMpqwz/jzscSKIzPJxA2
LKUTI7DS8k8QwFNG4JxXeXc9BpsprJetaarp/UNBs4p46O5htpuEl7x4JvsRCfxt
VdkeUQ+EYj2boFPU2rt1liA2feKNcdX6C0iXb4l8Cu8=
`protect END_PROTECTED
