`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbqOWhrwzJEwbcIwTU8TR6usbvnatYQXAsMkf5xjKbAWs9z+9TLe0l/Ym/JNVbYT
U4TJ7C7OVOSS2NVMQ8M8KBLLk0ja5mcL/zt/Ps98zoGDR54eHQnorEHcI6T6K4ZX
7TsH8Elk+fAw1Nw37EIF9ZEyGBNMPQ68kvM+xBbXhc8bz9wMyLBuVsM7ATbpPUKA
qQZITAQgcuIpLLluxuwst7JKOPAEQ4KMlnGGYNF/E0aECChxQJ9bUR/cbC+Ysnu/
ckbDs9yUhVhaB+CEHMJAdEFdNi5WJeeNvXKYC0bennwb+Bswc5vBbDsIaN7Wb4Zl
IruDHYBnusYonDwsqA/BrERe2DTZi80i0d3FB/5S56T+3hF8nuwGS4IYIDFoxDxP
jtAoISB8KMM99g4elgGTnKy0aP3WUl5QdOE08lvpo4m/tpUsgDLDWueNEolN9Hhv
ytLUjfINE2taKtIYqLLMxl2ejUQ4Pf3TKjexi9CjI8lsGB+3XeQ5xxceo2DSk5z5
oK3edesDN4GGg95vWtCbzcAi/E04t+7/6N77xMKLJYWV/+SS7UqkQ4wN5K5prGfA
UicxQ6wkCK48rLKm3vrCGLNIJg4woqhE9vnLa3qtqrPlIIuET+RUxeBDm2mG0CO0
iUuOy9Yxm5fnqDBFphnnNRfAixdJ2V4bnoNCwBRQkXrBV12/AMsui2FDJDm1+2ZI
x9Uvqxaa0yocbkJ7sT2gD+w3X9c2kN+15xiyplhgFJ5/PbOX9GZQ2o6A/pJPosf7
7yIZ3kHYAtQBxHFB88+yUMAmUOXSrMZbTYWCaWUAa5LzNheCH8BJBLR0564D77js
b9T7l6V8CXCkgUdasWE64urjTIBpGVLj3pqvMig4onTvBEXD0wKEAxNXJFZ5dgxB
5CsCkQY4W8CMPEtAGXwh9OExIUD7LXLY1NUU5/iH8Qn6Zc1VKLJGOmNkuJVBwWz9
aeOzK2vs1vUJ5PtlWPbeVkizvOsa01VgVHTxA1A+ZbpoZwxSJRsyRRjjPLa1o8X+
FhC7clX38ON7u+SAKRCXZu7qk3xMcLlNoXI7TAzqtcFSjn182NtnKwdgOoKKXMwk
f4i0NyXf/AUym72Z8rlbYMeMNWYG3OIVV/td8Xo+7FkAh1vGD2VlJyAqoEJoaF1D
ZI/afCzrX70DcKrF/6R8EMNEVXxy2JlUGnELJzOqX7bEdIeXXL0Xzix98Vd4Hh57
oELywrQSMA51+w6Irm3zvDsog3dc1J7FNm5TtyGO+PZYS9YzaBaB2MCxuYLB5hFb
6hqSKyK+pQyk5My9gJFdANxBjKKFhamwc+hVrhj2Hp7uPgctUgNdukYXsXGpiEGU
`protect END_PROTECTED
