`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ja0zpOXctiZitOEUoLos8UB3Sg4A+HfqNzZZ0zLJ0EGfZtkNlN100cv+9XroiJAf
CE2NSNRbvSyKQruCxCamRMu30fD6MorNxQR0qDt5eCAXU9xslATCGK2LsHKOktEB
7hF3okQ6ds3c6z9DpYp3sVEBtMLVlnqewYxTr+yBc6vczmh/+VaPqX27MLx7pZT/
dPtjJjEYZQNQpITjpeSOexbycunKBe5N4HC0+7kAVJ4vRsX4L/skXcbcNS2cFis2
fTlrpDCBPWhUP2Eapzn7wYEWgdwTTwx658f+YZY7xfqr+10KXFnw2UH7gwEjTo7a
UBS8dNBfs4YXhv7QzB72Yb3AuDCIktOmS32gCVhXB+Wq98NZOc3r76/nCfmPVZ5X
hB2uMwpJCEAjRftDY/m7HyGVu67TNJ2lrRqzSY1mO1qn6Q8zpY/hqdOndlgeBPj/
EPyurHyf/h5CBd/5Cm2/xc5n0/41518Q2F5ofTCQAmBv8xENrYOXnj6so8Kv+f/j
yW4D88OEVrqGHQGbEiuy87JHbXk+irQAops6rRMhjYQnYWS4pdPp3iGlr9yseHk8
Wk9VbPd2N1WoHlKBTxZA5nFyVCCT/yOteygx1dpwlbgglAWwLRolomtfQvefLzYX
SoLZggzsWXd7Pghdyfh91FIGEb7upxzBwZlIRDhkrNo8vutI59joQPOHgT5JiFbJ
ghUzPeF17mCCEoFwY0gkH2CPgsHICG3KlCkSiemBp12fKhP02dsQpd9gVAgwyzhn
6hAfkiflVJnxG8qXbc1uTwyB8pUq8v4C6D8bcrSAdIBqfi26Xjy9h0gLrQsf4pTv
TN2C2yS2OuJ/ykcP1qNSBVxQJjMGthn1/crRLVql5SImqUDiuGAaap7gCsB7uT5c
27tgrktGCHenkgl8plCsBmMHiRBJF5Nt2vMomxIXBbe+XKuc9Iuk7Ra5i/qdnOqn
tTLLpecX0PpAs9tlOOp4P5+Z3sIXfF6uILSkjYNQ3G8=
`protect END_PROTECTED
