`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1JKnCtZYxqDgHvTQMe2mmsoFbOL1jGlZce+KxfKPm/cCGifA6XT9ozz+ZTeewHk
F2vIdk4EO8CmpbJPoCZbC3vs3doZZvND7C6aPjH/CBPd3sQ1lsNtvmjdCngM5hsp
RImaLOmwmQ+5wJXHtT78qt2ShddgkeqDCEfo56PWgIXS9QMH9VJLO+WyyuJXp1Mc
8fk7iU4UIQe6VTyxO4MbsmCGH8daJdMFWPD0M+GVBtD03bJBMd+A50nVg/hBRjoF
pqZjCRbZpqnDxeTPf0Ui4EHeb1f4C5S2K3XOvfk6qM+2u9JPqDsh7lNKzhumTHDh
Pe+gJTJP6QZJTdBh6I33S4qdeggNOYln5iWJgGk5luc+DBC478svpQApN9J3l0iK
hNKCciXwLEpo4q+h3OTwEDKMXI0WXVkIAoX8wZp1eW01gDWz/ZfIiVoeGKI1gz0R
llqdop/1hbZWve1ZcNVJW11RYgvWCdAWcGh5Zst6xTDIVlp97ofvZ3p/3k8eyFhj
IY+vneMs6N925h7Qw3Pg1oqJ7X1yI9TRYzvhAEdmbtqn4PEbnzpmzLSOJzPheCrB
UWT0FX+mPGJP30yOZzuNm5wnpiidB5zgDliN8UlKGk/69X3DIH7Vf6LazlSoITbo
+P9S53AvYG4xPFj3Lvuh7tkDJMpKM9JTulNmRkfnnMBPZkKajHGScW3S1IkurLrK
ihJtAtRHg88ftCWVYHp32fSKgB7Aw0b0Tss/kmR0xtPb2ot7PYVbr+VGvi7Ooc0Z
pnSSn5tkxSVHoi2iZ6wLK6ldNyUO1u1Zz1sW+xuDpS2ILLJ2Lf/Dyx4Z7/SCIqn2
Z1+Xe+MtXJXc7uKK29TNSSejZyDL5WOAEqh2sfNcTyGlaB0beJ7km5RzHpPJTJUI
RUrGLdPuuIvwW0lOLucMeYkfQAXhQ8rf5OxgZp9WzDWiU5v7kYYNF/Kj7BL4xm0Z
qIIiSOSPcwWQMKNhyLEhSf7yPDokegfQ919wqibxr2maVeDuPXvVTnzix8Pi7qqZ
UfSYALUXC19dGmz0jLwGxzwxS/6smKcWqsBEm+aLPRWZLm1ENBgmlhGdv/S9N79B
3e9sm2Ei+xtdOkkZFb8czvPITxVgI4EIlar16ySjsae9WhlYOJCdG53aBP+IvxUW
xwofU+1fLH108+kxvd6d9AxDN/2tFqnBFv37LwmeXzgx2NYrr0Zu5oF8msk9ie2E
T+8ufVezRNRowRdMXRCQ7oKvjjUHkPbjAH7xCbH22h6oKrNCnuGL6B5NkXEzOw0h
pMOlj25A+80qek2aWq0mzEfgaiHuSRtbKpdc6zaMT638p8gnGOFegCMuvKdaj6+D
+u44IcUqG7G/+IEuwCvcVP6QjafA66sCo71zLi6wIpKb7EYPg6nGsjypENoBNwSO
ZsxD/LdofX5mnOVzGgbolHOnomQolBEz/Rj7IgrEClaWU80q4CHrlQ3Xwfa/kUw/
lUTnj5PWzHjcvPm8k0C9HLmnK2B8GxG3nIO1BylswTrFReehfEDdOPpQeN7c9FPB
9pNIJnx/8eQGV6AHvWp/NVykH2wUWeEOnqqRb+9HTRqGX/A4wxbUsAcRU+6lCVjq
9U+u0ZYGwaUDnZ92pHmxrOgplLsAOm6XGocT8O3uR2z75PEDq3FpJ0yznko0QcDR
4U4dMdTQ3UfABIzdql0TCnZaWpD7VCINkRtEOI8V8H80T67Wxq7ettz57viSOBgx
3jgEotfhujAIMYQQM8XMQWnUBbIGwcXSbfdNVQg/NRvBhmMrsRdETUMsRPBX8ATb
15QpcZnntasBBXu19ZOhDOrwsxmoaTbkmn/kh3F2EWZ6OqQchUlJTXvsAepeUd+k
HcJ+U0mQsPMnmBflwqQgTAlcJpaMuubKuF96DYRMMceVsemXQb0aCXnKbp1GsLhq
nKOl9xp8gk9ZcoAUEbb/9o5RdwzGEQEYT8uy159p4S9x8ST9yddeHSLINtjSpEcf
pjZvu8rO1oowfApRE2z9e3D44BpjPpZpMT40A1zj96/keFKkDGGpl7Yy1SVnXkkZ
CZhD15DIAWdQpb7IttqpWu7Cj+xMwoN4F+volXUn2kkQy0/iMJ+84mddKny2xXvS
4IdY8/RcU4te1dSayDTXa71m46nTlFpiNeDOv4LlKrmZ6cfXs13VHVcqEWHAWrPu
f4te8Sd2Hrudh09GYn0Ppa+4tumvDOqQRAI7ajDw4jjJxissOsSC8/zsAkgCaSGm
Etm1usWE7Z/ite7kUhMyOPdPay1Hk8oaDpTAqaejtb7zi/atBYR/m8cI3Oh3gVN2
pYcr5XJiyMgnb4mSv5pzSYrWE0waZEAMkyw15rkR5e/19BFgtO1RIJ3Ym5lDVoce
a4eVE/R1+/fMGIcb0nmAQ8uqLDfsxGXnU+bzpN4hcQ+pmwKggdhJbtODQpFqjf7e
Wq7Xv2YviqC40sN6rdeZDRLJPV6iYOFad8t4FdUr17UtEgv3dTYRLHAQ4z9vAr+P
NCEfcyyCbl9lzdJHVwX09F//6GhMO3G3xi9yAVaMxlKx/J461aWd4eVnLejKQ7Rx
2dvmdq54ZOA+kSsvI3gTBkMEzDIZpiia6W1T/1FJtLphhmmOUTOoLPkDXjGMpRJ/
6/slpFrj9bU7YeE2f84D4189xxJKwWSG+V3yIqCL668l4E3S7epm9kVB+JYtm0iF
3ZhTxYfgXSPaxkzNXXYe/dHSQdNbwrZ0MrnMsTcKI82lL5cs3D8p6L5vlPG9febd
5FZPxbEC7wwIZ6Ksj5LRA8RbHrZVH9aqv/ZDYLoghDWDuBASgS5l/KAgabiCb6Mz
`protect END_PROTECTED
