`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkI7xeokNoMq7q4scZJ5bcPYW0jxARaIRC7oDTN+6ExsPbjUIyg+rsHbNYz8eb49
U094lL5LFkrmM1qDM8uBzOc8TnOxlXIkBJcdsrosPOQMa4txJIt/SzsgLcYcRbpg
qVOrG/288IJPWWtzcVFf6D9WC3qKdT9KbzZUiKytGDuQ9wc8vDlaLJT7SPkFBzBl
9EX49KjvsFds1GhSSvsOSEffeb7sOw/mAVBYMymGyLW3i0GgslbF2CDnASPbr6cy
trBCc9UR1BaDj+3qLn8gsGaPxCbAeQZeg42hnDsX1sdU9CwncsvgAcVI+LI2CPv8
u1sbax3qB/+9d7lRwwe7xVZ6gHAfF0L+gW1q4IKj/XA3ah6lyeE0pO/f6O06xPYK
3TWQvjK9Kn96lgHBECETxIbbF5JB9WE03JzgR55R5NvKogofRtd3sIvJ0c+b3Xks
uQ4zibhUbP3RLD5fHp6p74TvWpyr6ZH/9Dy37mcXoIuweBB/4QqW3TQzp36Dmhp1
BA2p7pY4EgKtMpzTh1/sIJ8KT0HpKYO0Zpek4V/N1i5tB2P4Cnh7gJt+pGX9CaTP
6I1BK5GDTFScElrnK/Pd/VT7TTv67wE7LkfmndlkNomsysDlM3v0Q6qY3G6ffT7e
WHvuXt8jD6EB00VSzQBYX4pf1yBaTr/GuSP4qo3QQ1TvGQpv2Y07vdsxVil9Zzv4
7Pk+BYASOO6F5u/Gtwk/qm+MDRse+6TM92nJzG/o5Jp1gWO5sq+zABu/yx99E6Y1
yrcPnXVHt4ojOa/D02LH6v52RCAdhR4i6+aHCP158A9OmKmmC7J4Il73ezpyvyxQ
3uFhFfV3d2FoIFeDePuck6KVgDuWCOn1NVSJusIoHlp/QKSa4WMbr+lFFMTY53B0
nPfdjAWkVerJY+iGLWyRfULzyp8iTFBqbuiGw/qO/jkXTHeLHwsHk7/URDfinaKl
//IA8vbI1pyeJaImj6xZ+nqZ/uQif8yTpwLuA6H682xzE9vNc8gPa0XRjv9z5tVF
ezRtf2ofWnjRNVDmR+5KevQNzaPS9H5FPxeda56FbAXLme/pscW4SjfU3fcws1by
WG0YG8aFZURq3+qgVNT2nwJhhuj0IpDVYAdx55JjkIQX2Mh0NrEXCtYZwJttFMmI
sZcCB8p1pwiZQmnuyV3CdOq+86a6thow0BH1IAArD6zKXxyMxljdAa43CdWaMKUg
Z6mWVjXTzrtTchy4krtyT9XiGfq9Slgj4AvPgWCu1bAZy2Jk9DG1jYylqVV/4PdW
krzBdzjj6nceGyZgV5197kJ8mw7aHrY4kjfKQjaTgos=
`protect END_PROTECTED
