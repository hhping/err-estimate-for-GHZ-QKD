`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
25bWTlSqVEAp/L/waR2CJaDNjm4kF+vCoky9WkcOsl+6IHZX37ypTwHsL81H4AFK
bShrsxcAFQOL0QmduuZpqIOKeeg35uWpmRBQ4p2EqUoSZ1Cw5geRaD9ARKX075Rl
NQPF4MW/CNoRm9X5VhSNi2yO3ciPpSsKiC1Z4Ud5YBdgAYRg8/WPUTnP5mf62xJQ
Ah5OzvVufjre5qcNl3WXAd+feiRe4fhtkFPx1PRLGkiu6uy35oE758pHVpXPKo8V
riO2UeM5xyc0riHQsxBMDIovhXALIwt+WOqrIS8uIcbNhLqdVimDD859BqkdfXiw
6BkOJwiGZ2mIttvqiqgT3wBJRWunGd1Ga4xa2lbM4ADwcBnOKjwYrHbuDam8G2/T
EZgPO7A6ubcewTOqSeEdfw2r4CZXNptza771Jje7Ke9CxyWDfuyAVQaRbtv02Ut6
7IsETSkAwOueJew+6G4age5Towgro+8IqtQuzSI0x/fJCdF/m8Z8+u29iOfR4jBB
WjmNZXSxyQE0zWXY+uQRMa94Co+EhHAa4aS5TXz4kBisa8SKSlG1Rg5fstv72FZQ
fCpLTA6FNiQPMZHudFiuu+5XEyeVMWoAgdBv+bpEV5mRrqmuls7oHserM/A87uyd
vKvm5wIQPrwi8gZz1Xuoge3VCxc6fWl87tb42pPUaWO/73ZE8+c6tsn6BhICxFgZ
MS5KfjYtEacu9ikF+QgaiiFKxtWJX1L3CpNMmG6QDVfqpGcyVsPdBKJlt2K+kiU1
8qUV17b5p/GKNEgq4wi+C1jiZTiLxQiJrUvkZIDp+I2DxQuH3RD/mrlz3H9rvGgL
pTs6glrfAD31qkHJC9hK5uC0w7KehaCR3bsnJqvNN+0z0QMS7OvXet9KwMXo2LjQ
iVwD7H7qauj6shR3oSr/QgpwFyH2AhVGXEzluCBDqbdcYSpAKXKNVofnV1VlB64h
cEYttTbwaN/zd5rPamwakOiaB3bz3wSZA/0BQ0yqFGEZv75oGUr/YMTJ0S2o4qps
HCAMtPUTwTU43reQ1olUKx1D3dQaPUqDUjC+ln+wN9XWdnXFuQ71sxuQsuushf9x
R/r/cURuqgl4PUklJLXH0+6G4uMIeXYO81b7Op2n7XngvV0L4kCUN9uqql/KRgV8
Y4h7fq4doX4XUEticVKi4MSnqII332fiZkNeAiXyIWAL6sSHOQcz7YSYcNjYKsJM
guv94RvrKmwMpX+GhiFDmHOeh78HqABrppQhVskUnd9F4o/ZfCE6tmwaJI8uBp/n
v2I7AjUeDoSKrPDhrgkrCUC4Wsq398EyosxM3uk720xa2IxST6WPmhZ6sP6nKm/k
lXX5bZYvH4YW9lUg2i6F9KwfpdMt0Hbkd8rnCxrSz5EXeq2jIjg75F6Zid0mhK5P
HQaP4lSK6O46nFVYme7bJvxbVpoWFqYmmiiRC82l508rS9KMNC6TB/r1BZfQfKRi
JJJeK5M7HH6t0RcNW5mfflLOSubxsPsXqfeWbtyAMvd26pLmxhtTSv+ji8ppcQ6t
nXf240Fb9Ckp5jAzPve0LxhcN8Jyg4NUNQfAqwNRoJskYrm3t9jdXmKZKYLa2u/V
F7ioacsL8ygp2BR6SrY37PLVlTrXVEddwZSbRBNVMr8aghGDWryWzPLeWKE74MGH
nivy8QSdj6PqHH0RdRPzK25MJ+UQf0tENPJ6zbfOjySsHQa5Kc7M5kei49GODzV8
aGpE87NoKnq/VZwzlAQdkHsFptH7DTbN4yc4uN/RyFk8Yz7OyTBZej3VJmWSHCqB
`protect END_PROTECTED
