`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9gCizxXSRq2DI+tv02rcrQWAyItQXdi4xq5rHDWsGkutIxWvHxhe7OVzkIi4g2tL
VxhH3VUNOOsPoufI3acH3VJkUesn6dFumlcLm42SHfpWb86iO2/g6UelCAFdzPaf
qDhq7oUAVWRmcKV41MrblzSfJkK6gld/ZLLRG+awgJJhD6hbvYaLoH+GS7t+U0In
DI8cgJMqWfLlRNj/coXEYQu4kLQGqWz0Ci3AGHwNKKmiOvQQKJCoF7ucA5FKOWgv
ZWQ8ov0WGTJsXHfstWJR37YQri2F1stkKMK6t2+UEMKGNEHC1xHpCpm/FkKUeIgR
Is/RB1s1gW0exXQG4hkQ9h5OR+AOMPs5mgcnVcTyLTKRho8kzHjL1DePZbWXcaUF
uDKvCmOVZ0rpl7orbkwuTMshvQ0OqyZa98sG/u3FJxr38mm7wAL20N0QepjgMHnW
VBcV/MYrEUytD/C43b3QVVvqemn6hguBVip6zrNTzqGUQg8GvjlF144Zd41Yu2AU
BG2u3Engf3e1Whub9u+uSouxKu9wisYED0KjLpmzjKmA9Pw2qi+nhFCOPrQ1cWPG
Wy7+0ViowkdJQkgpwYVtye4BrPwak99EtdKUq+l7xFcNr88TQ4+zXv9S7YntuwDl
+EMUWbZ0MiHlqOp/40iig1Cw0uxxTpZEq+qbfEBtYzXqcS+8sMLtVREZbwIrFKJf
vxaBxKXR46vjvovsIVjnd4pO5NeI+fB3zuPsiVvtii1cy9Q1KqLcR0ZV3XBKsxI9
PTGXJs8I7XdTsQtKH7FkszY4rcVDxl1CIcy2cEPim/YZeE1hexbJXv2rIHxedqV+
r8hXjiVJpXU/WmPO6tEU8vLhVW+c10m+mZ3bQRVDoLwUi7nlYNtHzOw91euU3BB4
TAwFbLAe6WyUX2iDiphh0eu85GSDG/5+s1eGEXHIaDbHJFFxVqPzE/VmFNJxT7+M
ECuOg0MtbZBKG7yvBL0pKMYpchNPMgxjtnk/bmSEYioeJ7qbdzKzfDNCt97xhkqZ
ZBFkRKST684R1XEsiPKt21FV09Z9IXk2IPknDRw1nrlSVxWSMZYSvlzhsRHQR3Ps
ZR2H1NMYC+qrKFXbDBVzzbflkRpDyBoU86bbdha9Roe48bCaw9fCbGabBs6pXvNt
J5cwJMqGGQjjThJlvzNak00cnS4Bcs7+Clvgsr8a7f4Fxw9hojp6wDWOZDLn1AX8
AgZ/UZ78Q7X26Nmiyydrx4WbY6ZP9SiIcrGPnm1wiFTIcuLTOMcuYH804C3a1u+v
juThiIupq0vgMYJRGpf56Y9fcPA1CSj/AsGNsS6XnZYxlmbhd07sR3iTEuqOsbWT
swstmCleAY93xO0gIEDRJYuQy/LeQqJDfulNILwRepK7zOdT7ByCoE91loBf5u5k
q+SWh1rvOFOep3BtNKby08rfZoPoiJWhbnoPgJhtJagshfO4bjSFCneBub9bzHiB
5zi8Fi9eV6Yyy4KipqfChwaesiac2s2/bx6U5g45R8zUy/IzBdtcOD8ritNhml2Q
Bffq1VDcd4kAF4VoK/803i//oQsQ35twruOxmZFwrKWENNPYphsFofJRNi/HVrkr
yz6wl200+vPNxZ1J9NMTqvzoddCtxP7IYhsEoFpUZhBf8ARexnEfxwZTfNPMSC2J
eig9qdsa8ctXpC/vxpAyr+51NBu8uHwU9EeZmFemIfWjTzi3bBwyBW8+nHfVqzix
pO8PIF0fSULEBekLQlqSSx67hFYCZyVn2ov8gdFIt2syUhdmrk8C+wplG4b5+Lba
wDbHtyzteIMViwqaXge2bzxjUqMv3bf0MOxFcMzWuslXEPclgIbTQZUvzdE/Ct51
r0ndPEyo6wrQaKKbprS6eRv/6at1CO507zNmt7SvFA2P1vWuyjjY4Gt04O7q2nvH
+Z9Tu37M7gGusqSlfhYEa2LYhg4kUl53Dksk1wmM8tj88ntuA8FcXYCFKwPCDTh4
99zOYXJxjthG5eWyb6esdRGfjubWPaOkMjKU3bmrQ0uUSgDBTCUWurS+HDBoA3IV
RVQ7jhMEUYOdWjcy8snjn/C2OErny6bQx+ga+o4+FbIkscz2oVFPOnQiaIEfRv0e
l+BflC/fNRgmXo8yZ1bxiaEBprQizhxFPUcJu2ZlXndFOT0qJqRV6y0RVrq2WTJD
tlU7G8IhtQLgtXC1kEDaEbCI8gO1kotU6Z1Y8HWbhcnXov1Dd0wCBTERG4yE4K69
9rCUqDLCc1asW+8ks5dUpidG57e3ITzZ53STg9Po0OFljETGIFwwQxWdz3F179cL
WDAfXouEXfsTc/8lCzD+ET3nR2OPmHqicXk5E6DwnOG1KGu1QlSut+S+jmPH+2rA
fr7irb9KmvVGSvw8ILtvvEx3RSBSHmpSSd1ZeRB7qTX8rPhFphD3dWiuGuUhGNOL
qmmPXOnbVU0x9mt2/iAbeXiidus2ebF18Ydyut0qK5D/H+/UWmrtlM6Cqdeyqnmx
v8vdB9nuVIrKC174Ue9VzZF3dfMIkg1vl6ARlfh0BmX0VAF7LdmdDTLrY03sO8cT
kiv2hDWET98Pe47hrE7Re1xwGLrRZPA6GeOFkHxexyDgchC+CCsV4IqmtpCuhvZo
wswKOeLE5yUsOD4YZxDVbpRWzKRZi0KDdu6GlBLNU6hocfbm1cxfS2Rb2vmJ7Kez
Z9J8EbNeErC4puSK22Xf+9s8JKyl8iIP3iqtTuLFQnnPxoUMT0fjZycuGVKL2Rwh
pfMnDbb847bOAmMurv5dB29mxjg5W4LGi3ZnB8JNxgvntoc7p8H2snha/iOaU7cp
fHldjAYD3x8c8SauYLim6IEqE9DcAJuU1exjilsL/IVy1gcmPNiv+WBgvxdHP+xw
Utq1hq/F6xhZfaZ8ZMc/YdW7QXUW+o5ayeoI6BIZ8gYvGnUZKyEwpLz+oUaFJsEH
PzstcoU0VS5TIGHNZE2okmNj5VCCQaHjn6jXizdmHwZCwKMyqpEVmdUPJMLnNit9
uCPf8l0YAwVxRH4pl72JFclghhpb8kKnGDlT6xEgxa0rT+BCIiTTi2eFQFGcZrHE
c6HKhfb4/5Oz1hTUJHWoen8DNt00JInoLvC2C2l5RubMkSxG+huUg1J6sjN1EgwQ
IIW6IPtTzZieC+YmCIlpUFYEBFGdH704WAx3JSYMY3TNNot4sYJDnROErAaj0aH5
ZvglEs88R5i7gevwkDbBWs7+4+FMeM4kkBlusiSFZUA6TX8MSWG/v6bGcd5uoPhh
6dsU8vBMHXG0SwFOZQQTJs8e3ZOdMIYaT2lk4wU+T0jKsb4WLHQXuG2C5eEOcr4+
8LBG0ats0i3ANa71aCki5w+SY0LkDkimXLmDjK8RkFa0vzGQgteRnOhuMy7Hy+wE
IdBw9cv4VWxi+ewjE9afRp3AeIHzAXzTo0wzNOMbQvCgqgYG/Lbdb4GVx7NoP6hU
4vU9trRZJg/mPw3NX30o/sP7L18GYdgcojche+QTF1PrKM5mD6fjWpNbayaOFhp9
TFmXQqLph6CtgaxLwjRrUjFd5CvJYtKv3DXozIA3nPkYwyEvQ0H34uK0nTy5v54/
O26Atvxxfh0s0pkBEb4BrRd4vGAnZYeQvYeC3u10oFn4BxH/PIltigOtxffrqsPX
jquDqlqj2II8np4JK0Ynd+vv3GZg1NYsK0PUGVmPj4p4Dx8WrJpVBuqbhZZl8aF4
9AfJZq7YUmTFbR04aemUoCWqSY51WrK3IGUxYXgFxQOGz7hbvPyZBVhnPtszbww1
ib+5eEokNlF+qkyOw9wPDZxOZUbaYk2kInmDaZgO9vibxFM+j3dgaL7Z2m0kGzGZ
MDPhqVcW4EjC2NI4EGWlpbCceBA81ZFVgAWZKbydtjFKLaMDwYv4ZZYU6qhiCXcE
Box3dtOa+GV6MzSduD54UeAD+Jhm5IraQvqmsQI378Cagl3OIzTLKz23GDhUtioa
/1CLcSwuaTOvCvGBKODUibaYrdAz2PcEAEFh+9W1DnRyvn8OmO8Y9UaxuB7jKuzp
dp3gzPDZsNkeO2WnU65VKniUXxwEOqNT2icX0hxWlr1jv/LIIa39wGsuV5UhJaua
ghbjUaOHKz6a44tCo8Z7cPjtd0jLRoXWnlEX8u++76EU8lWaxEVyOobq2AdRdc1S
BV/hu+k4ja+9sto2kLJHQt/8Z7P1okeJXpnKwdhzXlGe2/tV3BidIQVJcLyZOMeE
DHTV3uvRao5KlpiCUVKwdRkBylMge04SVQ9RwuSlRvaSnINPD/jZoVpL5OPDbidY
eJCtB1eLz6cZfsLEv+RRAS/kyWaKRJFukYzFNMRzKoAziN3zpUHHAlo/EiiSTdFn
OwWvXDiyqJDuSjA5eY2l0ASbWzg82Onmr9T6RdloH1AhtISW0XL+aoDROsxxUtqL
VhZz/BM6nBH0v25fVgLbRKxhkSs02exT9q7AvOfpTtTQrWf6CrnDK0bYhHyKs4TK
+STDZ3ivRo8O/jbZWBvVRSKlNxPsvMvjCXw+izDDY5OQghlUOabrvHzXtd7NZl1r
LJp4JRmAQZzrCrwvnRrRN5b5TgcrlWCHBTZ+cKj2Xbz8vqtdB3B96DCDlPuUY5YY
5haTl24NVyQ8Bzw35BTO0sJ93cv3HBiGlVDJHX05od+0ERNO8phgv3NX9z+6wowM
LIUA6m6VkYt/gVW/WTojIn97QEs9oHCPlPKL1vELGDUN2Heg4BfaZkeoapfEO0mF
txq79neOuiIvdjYvzMgynsftf94nSUJv2e1YzAK7Xzmzd3+blWoKMRs7JGjRv4ZJ
6jVEhUK5/NyY8+mW8kP8W2jri+DC3Aw6VLCdnvowUJZmIgT2ryqmnfeevXD5kxmV
NwigcnsxsJp57THkK9Xlm61eNTcpQxiuRh4Qo1Bgm1OgG/C4P3jnJ0lbwlEKiC5d
fWtu7llRv+mZhwT6TDPMgP+2itcTks0sGYCZxgAqAF0WVfEoyAnsyciLUDiPNUcO
fTwAvqB1scLNtjWxIeCmUKeYz051E0ElPghGUR8aXeVeHEQLqnzJLlDq8b7FlvQa
tv8KxeZzFcTdmeW95s6cTKJvs+zxYfa6yKdmzDAwjJVWdbRjX93Tz0w8wgq0DPJW
MxkefPK/RNueticLS/HuyGaYr5DXvBOAwleNzlkPw4rPHeN7IUMg7X9UjLWEnaMv
q7z4+Fl1P+6FG88ls/r74fdnGGcFrbY/+YhO8G/qEHUuHp7sM3IB5m0mzJFQuscf
fsH7MSovZ8CNFzu3KI/43ISfauzgkTkx+zoD7XxsFxKBoW27/74Kswz/fSx+ZpAV
V/1w4n3ksyocFKQlgv4+tn0Xast3/lcVVb01sz4XyU/4MeGxWSpodZ9R+XqrrMCm
dtSnR4UQGVQqObs8JfZ1k0HHfCDP6u9tIlezesGnBU+6AHBwHW92x9M1Du1+h+pw
ZG7S9brKO+cW4h71IUbOQHSHluJHNDYtncNqCmMBIQRCZpktG5lPZT/SIQT9/iXu
rh+OYemJkBOuGXAOvm5pWtbQ2APxNtMvkfU/Txg3drbQrbFDyeeqf7awkhaCL1AC
H3kwRyZa5KDyKRZ6PQxILllYw8Zcf9eX2MQZiosVMl77c0CUDabc93IGniCSOx1D
rH3wjBB6qdxk/ARJBbc6d2tiEstMGEE92HLAAES1a5or+Sx7o+lrqNZ3WcI+uGd+
UpX1VwSsao89yn1Kao+CdgGivdpXPdr3yeq/oPPUwE8ZEYV/HrIn6aizRN5zrtg3
G9hfr/XPeQk2+Fd9B53+SA6noeIegxv6rpCuzgQhg/p8Zx4P6xP4DdqoDjI/WLno
nzkzk5Vsl4THO9eTkxr3+G69Ne3MNKFL9+RwIfMXMcudCUH75QcG1LD01s5NE9Ep
ACLomPWIIw95rUlrunSKLGpiZFAoc10T0kZjqyF0DAOvJkHwYxTJOeMuyYMHW1ma
av85YhRs2TzoimxmmE2WaqnP0jvRT036lKL1soR2rsgeZ5xxiTVeO3YQLkJjbt0L
8FuzIrlhm84h2EYBpuFaAYnBG/IL2FSnSHfoetFjcCVd3sJaUeLrvPdg9/gep+kz
Pb3KUmOaLLJEumWzcnUK+3vPRZCm7nJdEokMPd9uI9IPkjl8rIvYL7lHqbQOoSEe
0D34SU4cO7xOnddFoyvZOCsul9x53im1NmzMcsQ03q0xwPLJfwAD5+XyQVtjL4L1
S2F7rMIIO5oXhDMGHyUC31TG15igqEjM37KI5zM/zjMn6Jpj7CfFQFzrfbp5HNQe
tzAYHj6zec4PhuEdwE/B77O+SlkZ3ViFonjwmBUcsCxCk41UKZlFREWWwLoO0XlC
9MjJgT0TVU/NxFOqPzkLhUQirAqnSbt7VDSC7XeNao1rnX6hTCGcIaW4YzyNAT2Z
Ki2enl1Zaky0G8xYJbGxH5em/i/9e+R4r50EFdVLSymkzpoxedzj0ci2Mor94j+7
4h+8SFmbP15OjLUmdDHG5ow1XW7FX9gae4Eo1NUfvsPEqbJTAMDzpAwEG9S4Mmta
A4T+EhAZGSdA4iGKqA6AhKWLuxjhKp6pd3IhIWXGPMXLFuOfmbB0PL2MBQx+7ZuX
8FLOdMh1bF+aUA8ucIpk6zKHmEnLGMHMkoUHJqRsJ9ITQliJugtQhBinOVcGdf1m
1K3w/P4MWDh4LElVZS19Dxay22/XzYPBhJKuvnnXScMM5S0qu0o61RX39yYcHZNZ
xs/oW5KqiREDKHVNXckFt7M646UYGO5Lv+zm/TxOfKajvq1pUc3cH+WQ9UpZNPdO
Efy/7Pbfz63yqYC5kYmiHejsvZE7ndfPEsV5XskGVV5foCFvjqPU7sbexQavmk49
Tak3gFYek0gVTZ7qL06ap3PKsdw5adoAr6yX4lF3qPVBNQm9G9QcGPFeMzb4oeKk
wCmkjN2oQE0yIL11HpIW95chYyqg7Sq5DfvLvAaWgoTnKYh+dAxss1X3+piZ/jR+
SxzQMiJlUBFmeXNAPt1yZcRxWta40bX42uMVO5pnLf0egaTl1aPyaDdqa34g+oaT
lYhP3ZnPO6SX9qIrp2m0gA+pG1zkd8mBSW03DBXy/arvN/Yf9usF2fDnZUW6Q9NE
+BXExrTAIhqHcxL+r5gnQVS/ZapxfmYSwPkQ41A0yoadwd+hnKsEd3JhiEdvZLtE
CfK37oCd0UIOf+wAzjoEHRRNqHwFQ3x2K7EThE80vZHd4P7NEvfd3EOcAfpNScOR
YtGwoa2y66TTroWBQBRphglfnS1cl/LCqpEwvh3wceBuWAq4I+XFWOXxWm+CZXXf
b/VMj8nn5dPTNjWQ7IvBNyoEwsk3pJG+xEXcHNNcMTdwLYjeP0Zf41BmzZFE+92Q
i2JAxGsoiF1RUWeZRSqevHU4tzV/xAH/OnBaGpPIXRhCqZjiK0vkRZ4bl9J7I6bO
hMV+IV2EsEt+7kIf7gwGFxo7GLfT6EJq6Yjft/pb+eiTTGhmZUqJ7vYQv6GnTIuB
I5833sHhpHNVZDBTFq2yTPT1Kz4p43E53Dcve3b9SfYjOCPVr8n4hn6qlq0/aE/r
15dNytpqHGHcGjPkTzanVDZXETmus395OrXVewaIBg1r0cR3YqBzw7cZ94T1fOIy
xYEpFPBAUbkNy6MBijTo7PcnFJ2NmJgfQEaikcZ/IcCiVJrFnxYAjJoG+Aqamb31
3lrySsoV9y0pS3b5r6fWZEvKjYAPZMbDsRJgKVvhiK8UgKUae+OFLckD8dq0oMt2
0kda5dutUiUDY/yJEEIaG5FnA1CQ8iLT0s+V5iH8IeLC2uzPYGNqAda9uRd5pyFi
49NUwl/M3TU8+MBC46pbPypYCeGnRv5LjxCE3E3TKpdWWjZMYhd+6fXsrg4YMRBC
WC/4Eyp5gVx/ilEIsZlE6L7LMagSWQmdYf9yrvpbj+9dgGRJILKCt5XU9mfkH0P8
3VR9eyw7Pgl8r8Aofvk/deqYq11bmweZ/IyQvBlGve5jlybBZpHj7oE9sVtLMHAx
CcGCMXq/xtfOWXxLzjq6Bi2nPDif2j91mXRCX+fkOCeRd2gC4PmUjy1wmD/AnHC5
og09AeKc+7JTj47biAFEK88SP7ay8YLlEXji6UIq6H2iVtRMbdE+usFdRZ6+jkTH
SuRvQhU7uLL9FhnsLnHLh37iwZlVyugMD+hmjtVz+GVd/kcWq7DGFVJS1laKigWH
ZjXNtOLsnlvfFc3sWLC1xDolm9RqSVbEL8mQ+fmYHi8EAW7Mpcrnjhu8wAGBePD2
Wi0gZlPCkcFhiTye+zJRaULtND5dgZ8pt5BujMKmaFJLK8K1jAitws70rOWC9BnO
7bH9y16HWIPbDN9pObbmD32vSHzi34N+AJFDmFTH/SR27AB0TpO/sYXzs7Q8vzEU
/881rp3L4aYwkLRQkJ9hc1VNLLIM/gkIjS6JRu6eBbTwDxuxBePnuaLz+yxzp29t
QGAUnmLfiXFtK7p8FhsgHgPLPiNpcEFP2WwoPnUScyIlBu7TQS0VtohA5N97JRff
UQqGe/WEEreBIRxyWpjkUaLjSI9Ef2rgEiD3KQNQ8x/2oqhOdkbQtZbXsZRDqbJy
LNkjouDOVzQwWteJ9oGIqh3e0YnvxE8flHaUs/wlEdZn1nBT6x/omO7Yke0XQYfp
k98ibxJXfypNPYX//bnSPwsGvLqkeZaNirDtmsEWS0jintxr8Sc2rbazBe9m7pQx
KS/vZViQzOBIcq+/mzqB6T2jtbyUYrhm8Nw4tjlpY3AJ21gG8OPDndhgB1kM8saN
ofkq/h/+ulsJqrZdCB9n0NbswcSgp1RaGfCKnMf5xlcaMBlgbewadfYuIBcJDFud
HAhdT8eUXSlnBY8Xpo95Z91ZgAZ1NAPzJYogPgH5Ue9WGSAb+lfmNZcJFmXY3BLp
rV+bo2PEkG1mrEsKFqmN5ySTCoH4gse9VsVFaG6WDXRGzYMY3U8Lx1mnVDLz62X9
5wmQu1iNp+KsALQV9lXSvqyLL3kdo8OJL7bAX7e9tioa++O3JgS3KTvAqHEX+cBh
20p4EcOlGfah85HP65UW1GIZVc+yU6yEZRs1xmnfXzkCqQdrlw4oC2YVofSKH3xc
gF6dnEj8izOLFdxgFWwEsVqVQpJ6i882MB0Arml0mJCDC6OoACUCS0Pk/9V3r3ZN
IflhANFWqjfboqcshICOOOCWArE/UvXISK5EOqdapeLUVXjR7n6KzYCZpGavf0C1
XA0XGhWlz7IAU2hWcqeq2MXqIICNSESjUAHTyLg6SCVrvDIksX9lrf1eCoARJsAn
584V9MIxL4XPn3h+hY1y5GNQVTemy1F2XvHdyw8RbbXmvZF1cQOF1uppFUuXoLUE
/3zu9+3z9bsW52AOfGXlrr9fv5zMy0fZ29KAm172qgWYJhnkJngziHsmRCyu3U81
GCZ05KIer1TB4RS28feHvCVze0B3WEnFUMulPRfbsgG1YoyVDVb4EGH+Tw942WRw
mwrSJj6ywQjgYocvtPejCxa/bvov7NiaD/EwIjQXvoEVTpfd8XRCnb8hGDGCAh7N
ywFh1JDZNaH1ydRvTAj57lAB3S/eBwmtoYpZfOHiYLjK80GUDv/pylX8pZID5xWq
hCuH0bezAEQn79v4582jpg3JJCtjpCTUzFR9CFl/qBCEhcUQBhIRugretm0tBHnK
UpPO6DiZa6phd+u95hSME8NOxELEfLE1CBHuoGfWQerViao2dprfZc7Sd1CB42ZN
sKqa/zgALyvVNU9ilDpkvC8xqbHh5bmwsUAxTc744m1K4gchDI8m8JRKuPcV6ltS
uL8Dn6V5C/0EtLgfNN5oa0WyzQt+INy5dWBBY2beTe2zvQNnw1OvoIUg2YouqQoq
pZxrRJnAOjpyPV/QErdLzznzKZJYctJA++tflHcxLYC4t4gwgHW042MaRDbvRvKC
esP/p/cc/g4u6vAx0cWWKTElibx3Ie1uVjBEIHCQZWJ2Lb8nifL18oyDjL8NVbBl
R0ypG4AhNnOvy4PA86o3iU+PtgA8bpiYolTziN5yzjLdMr0PGdai6Hz8qCMtbezc
gjTqeVQBAjeLDBhgL8UJ8WbNI3eCX/DFGj6KsBeJYQZm2gX1k1xKN0Nx0EYha2LU
qIOoxm2T5iGxkOyYusiGkx9GbkiDt3lwOyFmI872W5ycH1ZK6bye5DgIWpXb8oC4
KrREfCITHqfZZeoKZqhNG9rF8cVow8YOahoqi25U9Vbz6qf4kEEY5hbWRBKOcU2Y
qq3yJUUUX9kZg/KRBNaYV42ojMhRpRedf7hqU+01Jj40MCZxcTOV5r608cNNaMC+
0tI0tGVavSTuJDU/Kn6TIbYGB6GIeuufC80W0DLCSu7rJqkGon464E6I1a8goNgE
qqFzQDvAON18P+BUcomy4Jv6T4AbHisM9A4IhIgc4KRxAotIhagq2/wDmqWZcED6
JasRICyELcdnjjCZMRQclYmQ14eJyW9KjFa1gjpJXKH/iAV8Tx1MtOr0DREf0mlC
QoLeDxKf56ay3F8JPkJVI7i2AtIPG2MtTw3tJL7QcAFKMyJCPEUMz9RyexHcf3pb
Gic6+YnqjKCJIr/EX6PU7YIKiAUqVYVhhIcL/OT6+NEegxqHHaJCSAeLJ6sXQO3g
iSOsUHP2KPcrI5pAuxSuUUHUMacFYyuq/LtyVDgJtPXZnt4fu27UKrZc6XYk/rZX
fBsho6+HaTytj+uRKQip4z/8EU1PNHxRRYCBaHu1OI73Yiq+l5pnjsCFRylH16xq
VOOwQtDQRKCFa0rv8RNIH+D9/G66BFWdJ/lwhCUHmYy647c0y9ujt18vi/j7jYdx
EUR8h58ADtApVB4gAxB4GA8uVYP+kwzmJM+CmznDSlkIxpIxsFEblKvuo9mgEA8X
DWbKkIFgzaEVeCjrRHBB6nJQp5fwJpvAw+KvUOV4dkICpBpNp2Uy3aD1FGhIM5it
9qAE+4dj94iCcilhI57VdI9WDpEdKxf5vU0Q6NcHIQRNz35eb0E/G0IO5Wsm0v2W
zjeUznx4a3xcJfGlXidsKMBYOXBMy40z2XF962TsiJbIJStUgvHm8FlzD04PNkcN
K2sjsqyXGW2E3+YBd28ks+MqZlRU8z7JWLWY02E8A0P2Xmvl+FsgjAfA564qrgk/
koxiWWpkYMDMhupLswPbaApwpfYSefKmQdYakSB2nf5M5bY3DDjNmdYJShFylzIZ
vi4pS81sb9/bp4+quXUg8agQ2zr2lU90xixPhhjAH8+Vj0dSADEwvMfW3Pskmael
nPAtiKTHxR2EwGskrtuaRguvV2jt2NbsYvF5VLiZqwHBuOq2VG1xHHPd0uZndQSA
fpmlCZmjivODavlbaS4Xi8OFuuiWujK5c6zD+6cI1dVkeDcK5n5axLa4UGL6uwdH
9xutESiilTlLxxHg6hPSbWQ0Z1FpiIvXy2BtFX0Visfj+MMSa5sSc1V/pGvO13LW
r4u0JYis2q/dP5h1eU1jfLWC6o7YvtDWY5OtPdmXs7QxrrEyHc/oAO66duLbnOU2
NbvKaO03m11hkCAJgDTav8X+a0ysUYz0L+gKuhB+XGE03mHICcjN/WO50PfXIxCi
hIagqRinTlnhZhjhVUi0htUvNIRb0nOBqbF1LIZnIRNjz8JwRkxE2nutDybGPwKE
d89jhrxNS6G7F1VVSYwlhESfFwRlxNLE7Nrh2fzwrdaBWPHrnt5Lwb/hvKSRyisy
u9fiR90HZ1EagRwxYswuhbCCa4v1ushnyR8vPiVi6A35PJ7oIZjAG1EODlFzq9Tg
J2a3NgLAa0uaHdXCyhQiFsoD6nqiAd3JgT7dmLKIzzlNAD6lv4kA59nwZNsXCvYp
VILW1Q07BnWkGS3sJ97wQ2oRHw4CULlYEMvHzkdj/iTVX9NG7/tsanWjW/1wPjsY
fnw+BrQyw85yJh+B4u0aT5O6tSQHim6FDkVFopht9Bonfx4RBmUEvYR6MtUccHI8
A+pSeFgHOOulGIcjDeK0D+7gJ/7klQeHJEsiV+k33ByNyLmcgBxzcqgjkA5tYq4U
AcodIaYtnRg8vy0c7+7bbZ9mcI4GNBBT3GeiRNzBLgn1LL8nvVtW8rMIjMInEH/j
nWC/jovFCVk3Z5Zc4JYudcFrEBebU9ghnNsi/6lujUnSvhqdMpjl3jF7jmPyDpPo
y8g77i5HP3tXS+ceixuOT8xa8Vca+9dqJi5fAx6PRL++Y2eehpRTbE8w5gq6OzWc
De3E0vPaglSGWj3dV5Y1bNZIPm/ncZxKrLGH+DYjvZ2rGIzXBUWpV+ODr8F5OCSw
5P/zr0eYk/mUYtOD9EcTihLE+RO3VqesTcJDhnISr8nsYaapXae0ZtCELaaymp73
U+cOFm9hZLQ0FbWG8feZEb9d77XzrHpjYqGmUCG2kj2nfy29WLGYbQQX6kuTGZM/
J2TcrFmn4vVgj7FslDjHK68QwPbHFN0aFvFCUGw1H49JSivVwSIFAupDnoXXdLdA
6FQwRyb+1iywxMdJkBA5a8iKJYVGeNXu4LrbfsqP3in+q2IX5wPwkCa61MOaziqF
kBLdh1cComYMLKw1pD4mlncXok96lrR5S+UvvtCeovrC/zdpem9TDopBZeceROqB
OgnT2kJqEzfKMoKxk5SqaB4MiTUrcVnnDb3dntek1mAItKt5a+CkaQ+1s/2sWCHf
O/+hx5wNTbeHFYw1Pnk7yw1WjnzdKIwLrNUFWX44zN+JjjOrnikYXGKSXGaU79Cl
Id6bbN5NHk2UtNWFv3n9CicNWSiOGrbWEkgiADxXNOHJE20y+N6oqh0vrtBlsv1k
SjmOqE/n8hoVtI0rR4porx27vS3t4WKFe6cnY5zaKuhuzg3QU/eNSiud+1tBiK7s
28G64uREfcLDmn7rp86rbCE7G3x9wzxCub0vq1PFf48tFqIPzwYuFU0tOz+ZVRxr
Y19U72dj/zot2VwPNx2ascu0f1W1cPbMSvln1cTa1flHSu7dMSi1JJ8yTPdxH+VJ
tp5g0iHRAI/4TnmaLVe8L4+EurznT+/hJdTGZzeCMLF8kZNGEYLluo/xdcVeQPy5
W8sXffObcoLeOTKrBUn+kgD27DG1DGXBGOroNlrHUEijikDDc3ROeXSl6I8kvxYd
8BzbJXzcVFkII6unq5sGXve5AM2wzPzyt+qw2031TSKRCHblJd3E3SBHFZXMc21S
yQEa7AwQ/JOpC33VxkoYWVqlQ1HJ53IfoWWi5kFzVeJ6bf9GHBtBzTdSHs/ms+mp
gTK3BDAhx4SC75mxvn35Px0Cwulu3tLWyzuzG6pD+yIj3Ra2+YCICdSF2V9iWe9r
0WllNSd7B3Hvbkbn+lp9S6sgmD7Olyhu3GQDTwt72gisqMDr0zYqCqayYq3qsANy
yudzF/iMVK5IZStuDsAXuLGxaDxFMemqAElNzGU3eKsPE8Y6+DkYTQpX3S4mll7y
2CT8bQ0GkTNDF7hlDgX1G3EKsGp/K6DgffNU3YKjATs06pZklY8ZVlk9kiFGyi/m
KnOC6zxXPkr/Tbt3otB77d8doimvpeGJAiv/uYP5S0kfD9kdOwk01U8Uat2HQ5KG
S7xgM5guuK6I8OU7vxan2pyPYaC2gsHdRicT6QmabI01rhA7JOJtt+Q2vYZu/8xv
HoDZzAKBJTCdDfBbbThiUEIwb7N0Er+BHhHD9g3oFg7bpIna3v08JEYyF8HPaVNI
IAonGoQReagOl8L+yT1v1MD6spTi0MAtIHgoUNUDKy2+bv2fNCg1mMgGxZCoraC3
/tD1/OtBw+TTlg0KX9iu4JdvBLhyKafbE7ywe4dFvdlgfRWdxCsP4ZXlK6hzgQDZ
o41ircwSHuGMMMa9G0BWgF3PMJRLhN08yQ/8Tp0V0vWj+xKc9Qf7TvUUytQnJV1I
T7UUg9DSQ/RvOtcZdb3Gw0fYaka+LF2xwkWB9ZBZMZdY4TPXHZyx5DIpfYKjbKHY
EyuHM7TrLFkccUPMJYpTTaVNTOLzNFO//ehvvu0GCHaDrZz31x3LmutNR479l+hJ
R+RdZM3+bIPXJINdfpzdIHOjk6PS1s+yg9rKQyIERRdYNksmyH9hUrbLZCShMoJx
36g3GLwZYzKAAy0TJOiJDvNBu+/IJVnf1zIeyYaz7Gz4ytEhIrtNp7chrYFsjPdg
tRVDE74wlaFYeJnr7T3Ch/cCFdfELU4Y+HFPGnWg/7mhXDEnjq2qRvOa76ZjqzZ/
Bj3U5pn1iTYg9rUz2UVXFOJCMenB/b7oMjOqPnMfKCKHMn93CuX6TxleQQRxcG+T
WjSNn+yANlTvjetfngYpWwsl7OrCobhf2HeZV3eAUv+Zf19utVyRjaF3LRF1Yvc2
ZUDfLX0dnRPxUb9VaYzZ8O3EhCDd+Y//YsgFC0WQ3DyB8pM4W7CcFqpgZiZvPMJu
NJTEWh9tazqynB+QCYfDk9+g91yKRUM15D0ZLRchOaRhDKXHN9Owao49GXv2X8nq
RCg4Qw/ggkow8lY9PMFhcOUhRrcuwzLpm6Zhdm/dfAqb2HqhU0Ayba4oAJAsnFDQ
BLBEXyvep424GmEXyWDRuec0cA1dAbqxM/NeA5x4RqP/VjTH7/FQhZ+TLrF2ETrx
ZjsdqXu3ZcEGI/r3zX4iAOJhjA62JS22XGH21ZjEf9aPogeWl9R0i+jRv/w9rqa1
CatP1NHb6RbaBqi45QGLoITzm9ab2gkJsGpN8Z9vnHlTQaPqnaMqpDK4s6MigZnB
5N36FL20X2txRV0iC1LjN400qKm0E38eR88UYY8pewtGG6nGZTB0o8shE3V560/l
8Nv8mCDijD+eo8OgEImB0arPAiJB1+xdeKIKrUZBwLME3wq4vQh2LxI7okvIg9yZ
93pTYQXwxEsLKG8YVyb4wvsruSSt5uAQ/flbI1D+VJmhO2VlobH1Tz9siGbhT4/E
m/wAtCjl/Cv17DnK5NUzKbzBNwF4P51eajeCqerASaM9VuQYBZCWxmkRJkyO/oEG
Kb9A0XKzV2p/8icfy6pCwHwIQdr9YFjUuLiiHw7/4kAPIf1Uv8BWJ7MskLdgG5+i
ON99ZhooiSCOvLzZM/rgCPQFd4D6dPQoM0pURV+IvvKCyPPc1iiXJqAYTvYhgamU
kBz6M1x8eoUEDy+bsCnR4MCVOLfOhxT8NEsYa8ackb4t0dhMhjSRy3TuHvXllbWG
39rR1rVvNuD9j2kD8gwkEr8aR0exMqORK+uHG2vzEmIyb7k5kU/yfbuT6/PGqimK
ItHLEm4WOXRM7awT31Uk8kZbITbD6saxCG14kRurL8QSjCIZMpVo8KEzHCucUpQX
I1trWpYkPjkg9rXzKASPVtFmW7swTRsHdkDv1X04XhaVc8YHm6UGRZdPESU2J1FY
JVVEBDtPq0poC2Ekf4GXgLUheJPy2Qm6XoK40HFtnIY35eC3xKgT1nzy6KuHScZr
leq003UWpO8cc1HcB6iEB4uzE6CUU5FuF5KtDmvwnIz0UEtmTH2S4rtAvcX3nAHL
qeN12qStZKQYi8YV7Y0RANTwjzR8uTwFFbxpepH7zyRuvYjHOe6Nxb3pi9W4JS5W
Wy5rx4xSL4hRMOwvzbsZeELggSkSMs9tNdIkaj49nXRScjrp9qdTFwGqG3pdGovT
5DuG7SpVM+4JoxyAusXuvmHDeVQ98CmOlkhwohExZ/W9niFs6LAUjPAYdAXQlxhL
yi/M4J13HIJ0tU9IOEeAJC2iWONeHRQLYDzDmNy9pmesmK4ZI0uWaDapDBL2a2or
RQH3IhuaVP7S0dwAA+M+1F4sjLoh5cWelMSIEcrkcCmzQ3Kp9ProHXTBnbUV05EX
KAbYtgV3o5pgOzVxz3QG0qTLAxaXlR258Q3vQvU+vMUAl8ZR3PloqV7Ae//Ma57S
4m8fUsCqWhZJ9fj/SVzwsskrszCcEHTX7PFwRq+G4x2yQjRwv0DdknhTFhJYoQa2
lxaaQQHfcJEn2mkLkGjB9FDWOoauArD7P9PalED4xEbuYu27izAI70kr4wLK3PGo
/aGd9i7XHltyu4MQgMm7Ctv+vm+GkvsazuvDDGkDtZW3nmX52v2WxIEG643Dst0n
Kb4h9FqFO5rmUeOLRww7SUyGAb1bd7FoigWN+kUrROdh0Fv2mYubaGmboZV1zjxq
5RBRw5fuWpbmM9fFWFpj93+9wZmn/IvGzlKKq+SObRWNk6le46ln7rqk/4ROYj9X
/PqeZq6/g9SnTXPfabLQvLDodIc4DAtL4QoapnxTB7N3M3+wMyFW90rDMiKj0gu/
QaXw0FJ6s243CH6WGRwd2CjxdEZqPPztHKLI5MhhOoHH8HtYGgtm6S0usBcys48K
B/KiAJJrbdsuFpbHOKjksWij05AHXinqumgXEvD/eRCqHfq2Q9pZfbM/sNFOA8MG
ha4YSoifuB6SZZSwrpfLtUjAWVUEtAzbgw8a/bFFCxiXLc2U/pRlTukUVMqEs8Ux
zrzqw/bDRf93IpN3tW0rHOIFukGIu6YKyXcFYBPNY8pRV7u55auqEM+vmAqyl2Yk
MZkd9CwEWEEdvJtm5YwMH3HdpPyTC4LrsHeaAeIjczGHxbcuofyuLaglTDFqUoH6
KCN6pRBN5Mb5fF2RYOw5AuS0iNidSyw6r6Ev1SlZiuomTZMx7UTI1VmhunuciyhX
yowrM0ZU4zbDV6AebiAbLnDY2GVVrNqpNDoOwPzq+0sZJtTdBPYOcfKYABX5qNuZ
Hg8pm/SvaR8fft9iuLH+mESO7U6RWdE8TNpJ7myvoYTQ43t5iP+tUs3gMld5waH0
7B2iH11YAh6cvkbDD2gtrIRD5r7B+OWeT5ByS3wuQPlJS0oVI0WllGSxkkXeRWi3
nYmaU6AGkN5QGC3eM2owWE1emowA8cM/tgfNO5LkDVdp8/EocFxu50yTYeJDQHJm
cQ8SGOVWx3aSAfQoOemLLzbUXJ8NbZI5stCzXwVn2lxkEnNfhrbJfLxSeryjSZmH
BTCsuX24J//OBIpF8u0/txMw7PFwJA/HfW0LfH3iwbiBqDnNihpucxiUktFKc6lu
7UHBEEfb0YUPJDJ++fKqHOHIow3kao+KYL7bvqbOnLsVHY9GZoOqBxd82zN0h3Ze
CJpHOpZw2y8KBu11qYVEedpIStbqKuRsFkATQEXi9RzT/pn8tOw3rLFcI4xWCnJ1
cW+yPVDMSZ+LjCVFGG3r5RW1xI2IET3Pf4YEzDo6AFbDV2UFID1eBz76nkpzUoIl
WicoX98rYoMxmRU295w1KDBh9lsQaLgXlKNWSv5lLRc7Qb7wcsEH8m8T4TeHq2sw
0pFa2CchSGXWnAJwFPNGdPRvXMb/sj5psjSxwyGgh9jd58klHcuZ9igw3NvBrOYB
He2Xz3mwa7q4T0uSMIVPy5A0O+4/aPEr6fOGAC3PbURfUqdUT/II5C1KdRlADJb5
WBqukGOzCxtSU82ibGmrcKq2UBZlDd0jNmWTCCplWDtUGY1AuqLQOfPnJG5b1OvN
VtsNpbNO6XwA9dkKiuSMuQoNgh/UhmcB6xsrnUz/Kj6Nw1C1gAa54qFpKmmhFb+Y
Gbf+PreBx0IcllNIMvYJOBYH5OIWC9MU4rV6W/1lhmBPQiVlND9qs2mg8N06w3cC
mIQBaCSjpGTJ40K4j1YWphMukMqLcQaBWvWDZfOGMk89MXata1amS2cpy/muXyFl
oyIt4/iSav2wbs+NzMYY2pVERyERIxDprn0kg1JenP2sjGPLeWyVOSbxdcW5Fk4e
qiy2ou8HhGeMPYEaKN2m9EYce2P9v+enbhJ8/weFYsp1nHx1nPcAu34O8xN2Kn9R
v8DEkmGcKfYG5Gz0N0e6W1Mn1T8O//OacZPY/7vKJ/bpB7nvSw4+KskcBG06Chiu
m4cFikZVQ/EHjhcFO6xrtctPh3YvHgsT3V3qyiQbXnSLjXFO0AxBBFZEoRavlR+r
Uag6masBO4SopcDTGkfkStVDVQHTlih+EornZLoYV8bt87W44gjfs05i/Ne0LAGz
PDXSet6u0RkcFcG14YOfAIaPpPU42rw5QVYDgaT/RLFlzqBhXSBS9RpkU1VL8MrN
T2AZq8vbY+GCO2tcl5LSnZIM6pjVnS9k14PTmOXTSjoPRSF/Df3R8hnrld9m0eab
R1Y++JrFduq9dn3xZ8Ilvein18y4oRO7LEdX4PJ/HJxnO6AhYz1oJJBc4sRQp+lw
lSQ1sqjUCzXdxy4NpKEy9Kmu5ceg6SXwedh6ZCE21qD57plBkM45PXjtSYa4rCGe
9WSIBg/pzP5lN3aGHeK6vWJOYS2j1F4RtKZaeO001TfY8Im1VwSJb0c+V7GKUsLB
Apk/7EyrVfND2xnCMqDTTga7/eHnMOb/PJ4i6iyDIzDyTOsbqOa1RtCQjkUJIVLO
bbfPyW3I7v3lAVCy5SMyJH4dkv6w26jgDCHRy/pGsSOxdd41GwFS4yWIckkiOaUq
in67KciGl+KpOYetvsQKOJrjYaA62taYnFHWH13D9W7NfQuiYsjKKt7csEqiVCy7
UOKIMpd+j9q/WE4cPFb3HbJ+g7O8BvCwvkwesqA1wNOy9ZyT9BoTcfF/dSAk4hxT
MY0v53T/nHo7LE/LLpoYAN4fOPvGn838FYCCar5hWKCgGtBwBdzeaO56iKRBt7kA
ycJ0/dkzJBoupuEv24OLkjmEdlrJAdnfo5gnGAVTuPkmX9AnND/NHXYh4AFaglCJ
Kar1Jz8Kt+gIuvU/pDGEdeR1iYUXvHQLHeUmAn7csDiDrgyix3UkvXcshZWU/EyG
cPNRUdwa7m99/nH+l49/XhqAqbccSJsxzQwI8TeRvjKcSc7MdyU43O/8msZHjgwt
CPBEbsNjF65BFtFRm7QBp/QA4XZcInltvTvko7emy34LWEareuja3e/OFMOKajbC
vpOuz5RZS9CfeAXv2qEyLhWQ0gv2Mztc5vjlABiiVa5WbBNHudwgi3JsQKAYS6Oa
KkFnGWffwfcyGPdMxtUcpECP2VSvK2BPPu5Pk148KaOscEdt1I6qoatk/fJQy4fn
hS45wupVK1hrH1XlmgNjED+S9Es7FMFZu2D+wNDIFuZ/Gaw7W1T/3acwqP63mfM3
6TV1/rSaNDvYo8eD3Gc3373zVeSzqPgB5toiA0/F8ilgOsinMkalRMyZU7Hsxk+O
7/nTp8c26s8eKb7PycSNF5qU3S26WgADIKC8D9ysIzpAj7jDXmONOy9MKeRedav9
q+fhoZrn1H2lASZPZD/tS1eGWjoJUKoYKR6ZyrknSG6zzXNUOSjLw6Y6oZxmovui
l/raVWRvu3VzvnJMGdDUSvBmM8XoLjTYQqycbxclmkFXXU6vxq9fuvCrWZmWt07I
x3xJjWsbL9O0jrU9rj8TaFExPcw86mj8OPPJvRTyk/a2NBRZLWYD7uqVEmmzhj8d
pVbkDu4y8eRjlMuoyXSK19my163jJqSMQ4UjVdbef2Z/BGakIYaVtrrM6TlFQpuq
1UO9CpDJg+0XifXp0Qb14r5gV5fpHKCmGo+pqHX0iZXLb2nUvMlnjmn5hmnhI9JI
aUqUSObFAkmYIW3kia5GQltHY3rz0noUw+B61++aH7/Ae1yuJSyWvogsYVJk1aRh
SC6ju8mULxgYITp1d/loNFLm5jjG8Vw/XkQFGvTbERPCbaNdWYT/E/dDpbh49jXN
yzg/enxP+tI5FGZ4cNn2FA+iN7u2pNflvHeWLkkI0JD6/PuXp6327zc8RfL/5t5z
EW1M+aV+F5vWt6gEIEcHSqwt7B5ZC/wXBpe6LoBNXes+zwLmRFDY8ba30CIKIm9+
dG3qJUcntYQFG/n//F2+jkfciIXrEQSbPiU7fhvyr8v4oEM0CYnFKvp/eVCHpY/8
RZnsYEGCbsZxpEAPMsUOSKhXgA+eaelcbmfld3EMpXM/PNdWkvKvfkJIVNMmlQ/x
FfKX4+ERpnkJQ9qWzQ80uCb22Hfs37HftZCXXgzncZcLt/t2Y1bqoByb60bIO9MQ
kEUEyFqCJgvIHQqrvnTZcwFfUdNpPuE8H0SgwZ5M03wzEvGKv8lQTo1hWugpY1cW
RybNLP+2oj3EJ9tJFmUVhoq+OmGCOx99O9gc6ufhjUBUKaIthDA5WQHJlaJWHIVW
GG5qs+6G1nTgRTGmtDv3mtch6TPttt+AmtU8eny9Iu/U9Z8oCcIVPqGog7lg081D
fFYYyvBMklpBN/McFtIsBX7ozv89LYGs7wMis/vur1n/TEDe7UlM3o2W5jbIzpcV
DMHM4SYFg6WH0RgGrK9B4E/C72yGuAiZP7RkSFhGBmqkzEHwiZ4Gcpntyn8GY/n1
pIeOFb/VOFyOLPiyDGsqfvAoZvVbZCpOHxLQVPei/fSQuH4ImVFL9k5puqhB5+4p
WJU0y15z7ukqKntqbR5q9LeV2FXfH1n9sNqkBxXGA93c8/jQuFC2DIlrKe4YWqAI
WwIEYh4LzBkwU87E6GKJ+LcMbyMddZzu0VZKx9hGYGCv9hUBwXPlw/58WgywJVq+
GdAL1RtBgecTECfcgKEydo/dXm5TKXkjz7AkEboTYSjS+jIsoYr4R7xGz0xFIWGm
g8BWJ+86h77RnfQRx7wSXpkiQSTB6WBjNKC8sJ6uQECuGb80lu9omC0hTnVLzRau
85fWkzQj8GjQI7q/ni3guSbINptJM5OnxPF3hOqDiE+Wr3mjI8hP/73zhaKNgRna
iqT3iMJu75dsKpDoebifMkDRBMTGxLz/9O9zJnUjY9/nvZAWFnZBPtAvfvETj1nr
Rfrc31HbiTrXBApOScHlriwR5PGP9mTrbhvQuYKBInGVyf8w7xWhRXBTEE6JN0Me
xC2XqbX5VnM6PbfEAkGCCYB4wF88aBEMAh7TB6MyD21AXaplzIYmwRSCpLPQczWN
Lg1uGHzdL2v/i0hyDLlOvvdfwivfiePzk5uSBEJDV7J5L/geAI8yn7aDFKMzajTX
a0CUkiZbYudFfHVyLfaxa7ZwUQho+lgbz+upw/gM+agtHucH7Wo2Ox7P/ENkkOAW
HOXWbzXj1HL9N9rQvw2Pt5isbJ/s+h6VQpcQM4mvCGCu6mML0+4qEvB0xUNnPhD3
9eJuuUZoUrSf8nSwqYXCxHOfpmbzGnF0jM0Y5qzRnhn/hSbLYMVQ8LEgXG2h1QS+
ulNz6R1v6BuGbc7A6+WSLDyLuy2mbFloJPxQ+7dm1x0IQMOl2mGxgBEvlO22Y+jS
fHIuAruWvQblU++JpN1boaAZp7t2W/Y755s9AnqtDuvD3A/ovRJ1xkUgf92cTOq/
OtJYMU0+SfodLsXR09Q3K1PZJEmIgwnqtgeXfabltz2kB+kAm5nVomGrNP6OriTN
Ai3UBgYnlDd5O/zloHx2Jm8akv9Vx4JX/lBkdA/b4Si01QbPuk10A9SvzmrTMyEs
8UaBQHmFMgqXQ6GhgMegEhSbJYndXISyYZ37cBrQmsf9S8cfK9c5CYcJTZ8iFZ44
9/DBZUTcH/l22SqYO7mYRu5dghUE7eBDdSk466X03YlPkPMewu2cPSUupDQpO7Al
tIkWgIMA2naxV2CUx8tnI6F1sGTZF+v6C6zKtnowDduhGV5jsJhqggUGAXAHESbw
nv2BqGtPPe9mnLvLWJC7JD1qN2khmS5jRR44SlyNqLqgEF6I9caGaQhr2FGLPYVQ
RrRuPa+eDYqkKGLSYncP8ATFUH8khm/pQkS42rVqSfTqL7PsjwOc29sd+fYV5/ym
uSxMx7NuoyOxSpoT7gW/LGCvRVMz7BMtUrr7Xdp1qeqaWPYAZ+MFiKo4Gyk7gK2F
hT6CSThwtVmhQB2RQ1m2ECboDPAH8SPgjs6hocXCoTG2CwFWiTnRCLVxUqi5EUhQ
xp66v7G+tYOW86wbdA1BBYowOHbcoQp+L/Cem+v5upDS9PvwjXNZlangAAhiJVqR
DMnCrlRy1LBj+/Gn0Bba8J9RfnnCDLRKW7YTWvjK3ggeRXeXztmYsb2tD1K6bZHw
JHhczUB1oXdjmKx9744gd+tru9rFUuKK1yHge6s/RZ4xUEtuUeYQERn9dbJY4zdL
EoIwjm27rFNadapJChvCFs7Wh5LCJ7rzV1AFtJ1kVzHHxGceuMadDy2cmrGAV7+S
euOw8AF733ik29S3YyLqUAP1OVPyUAgaR6624yj2TiJcyrN8uaX5ApDOb5HUQtm5
6YdC9IfoP78vqRM22TqDotHW7y+hC9FC9GsuEyXMe1z2mIZZFLCQpCb3jGYIZqkv
3EbcO7BBIU6Uiv1RsP50WNYQS2rI9lxHmFD4YmlU6ko3MGDlEak14xOVUPwz+BSU
QBfFz4t2xpzhzleb2Jwvhl80HmDZD7tZB6AuvLXmrOyL0dZxtgpIuV+owoHHNVN2
Cy7nVJmYEfS4t9YjrTbE+WLwtjTxhamNVQPqiS0MFE53frUqt8zhDdvzSDmTLukL
zFQrgtvlpuLz2ZpfF47F50fjsnUh0FcCin6u9GHjKnQ3Sht0Q6KScgak6Xd52ui/
cpPGc8Q8OXE24T+HdETA6ocpUxEmkCc2Mb7RXnlLnMQIhUp1aTfxAQ95+NFJCidi
H00LBbCYOc5c2UrwKWrrfrDaWE1Hskn5lnfIVfIScipJPPH6qt0/020GWTWJ5TNj
OPsurjtZZ1UDNJVi5+2x+TC+0fjD51m0C+vogQxyBuOeuX3Y89Cw1m6UXS5MMEqW
fhrrJjBOkcwxMQgTu6CVV2tZR0QttuqqG9496Op01KWbd70iDDvW58X90U8HRluf
9xNH640EeaEdD2cZr5auU215ZXUg16JKCns85xZz0gceQ0z1CwIjkNzg3oarwXR9
JCD00cHq9hj4/BFazYYNC3Wuppa3+wzLrNHlU7e+hEZuNp9xT9Kpv6BWacQ+BSIc
DX+zvMb75JGz2KyFiDdTtN8lrW2eelFDiuNQDhQudGmHWK15NCyAU909YRY7QvKf
sE5SU94cuvWJWwmFc6syzlXA8o3lgWcFhyckZT2BaQRGe5hyJphyIrDu/IFwtp+7
nEwGkuxML0TY8UyDQnlcgFsj7/ezVEnMc5H+3ZrPF8faKoP7LQK51H5zMlYSnMXn
BkyvZIupPxyMnhH1WZtEuoRB9tHUrq+SS6cPoQxGWGg2R0r2m8rrkH5x1dafSHK3
COfmFWqbcmZw8HGSIHNGecq9zza0npjUnk8Y8ALFtin/HbEBRkZmZha11BCaQfUI
j7WDjG24/gjeytm2s4eXCUMdPafRZ5lmyLdfZ6wArqUyFSPBEtSZYEwjioYX1LHG
OAI8uPaEh0MkcgnFQXxGBVq5Z7sVpCmSYYK8adO9ht9T6zwfoggTWMcAaW0GLhEe
aoRow/Gm4SSmH/LKTjuEZwVazOrHo7QEGE2v7n1VIdSt4oUyTRwTQp5gNJzKk6wJ
htxbHB82WBvCMvPuSzNKS3rDcGL1SHdIANsRNVoZFSIHZR2sio4ouo2dUIbaEL9J
5FDBK66icLf4+dZHIUZiQJMV1TiR2icluj879mzd8Hn076EmjVo+njdMwuSqmqjp
u1XcyJNxvPnx7pYK/DZsiZ3z+IAlCtEJqiKkrUszLGg/2bNTIAslRmYEIIcmbE5l
5LKsq4dN/NZQSuPKxbpZTKFXrMw38v3Ae7RQHyKJRlx0e3WVXWsz0LRBkZHz5ZTj
CzHz7LOJGTVGiBKEW5d/kfcznys6/TSfM2qY0z3Zk4093XeyK0h/d3OkY7AjETBJ
dXQMg1wgeN7Mepb1Ao3oqm2oW+BgvrCWXD0VhvJ9gcdgzmPXbQnPYVm3dZKXZ4NL
zqTwAPQY1KCgX5yTCnfgNu61QJ4bxE4H5lmIdhiyyN+oOh5Sx90Wvx0D9PWzKg+7
wfh2WBXXe72uPy/BUGgtaLtGL4YnYLlQkpRz+NUM7E46EFdx8lEITj0vz+O1LAZk
HCoXYWFQYDRJmkgIAIrRZubpDEcSmodmsAt70VfNmD0/CjgBDys73FfWoucXZaO/
ZdigOrxBAJbkdknQUYNZkh+CV9vzDJzlBMxq1Yn+A4uiAsqdyX2nY2skJG9xm945
GLD3eXShLHwJGyPh6ZMEl+qxUP/ZrwJgQa+Im1mb4mmI5RfRdI5eSEUgsfp6gFrx
SGRVqQLA1PD7EA/ynF9AyVwP3WdHPawXgnIT9f5Bdgk5suY8OQjyd8enn7geVLDY
mQvsWEZfbRHB7I4PMK5xMC0XoYuI7KUsp79qvPENG/o2xRtPwiOj806qxotWq7eP
wnTk2NVwrujpXcFL8RExMSWDD9M+D9XLXirop6h8MGq0xGAoK0TSizBpEDCjGYu3
JMBJ/cXcJXnWsDM5vNFhvPZRSjWM2RmGHU6axpo9K2rGu1aRXNTG1qAm7QN6UK2g
pJPEAsSSZqhaVO26dtQDUST63E76Qc17jZnf3lPydUaB3opi799TqIahe6ooKOPm
mWrnrRymeNRrQtV0QocKevyN++DkliZCva4p/wNU95jvigtzpGLx4L5xpKP3exK3
aC6mTMOwv5JdjfZlefL2T5R4cuKeOy5Gqft1M5VfgVzPFGsxCfFVQpJ/tijFzzls
KRjRkxDpjG+KFTGQPaTFWOFFNX7q5SshUJMi6E5yv3vo4UOgKIN9MgasHSrTP3qt
iTWsZpAqHej6JC1BHV9dJW5XJW53yFNASF4ynasKlRqzVsBFkp9qAoMIWErnkTBR
lsHB4hWlZFE+LjFdfFEZABeL3Es9Uf/zfoGpd6jJ5hJDkg6ej/fnlvj7FmxOhh7H
SnhTtNT91MOhZZelPBhMOXwEovfhOlGOv322r7aHRcC4LuHCMK6Kp2/AFeY67Iai
heNuoqjwh2PIDtjaeuMSRsOYipandEw3QlXRHQmiEaYi5xEmE6PnqpgWpa4jS3dd
PwjtFttxP768v1Wr1abtJaatOUvXZnTN5rDMk7w70EILGRwJh7zueHFH+9BOU8Rw
Q5F3OpA6XjJT+tnOCJRoObFVHkiouLBnGe4qIuqYW+rdtnvN8oWJKWix1U9Ns6yZ
nsezs4lMZG9BKYpCnscLdbR8tpQ2jHricxVxV34IJBQbsR8gKbyWEkQsPeK4mToD
wJBQ4WQMzhdryM4uxwCzD9deCFQtku+myCO+IXQB8C0xug1aXabiWmTaRnVNkjga
j2Z9rbOoFNCs5PsZViIcyLgGemUTswFeNPjHd2brbUaFtW1GN24dmSTYhoGWNYXe
a5Hk2XEu7prSHfCg7bV477A//glH7jsq6zJbOhTPyEKRCnnuWAWKQywObz0g52sF
qKqTKpBZjCLuo2K3+66YjFrJIO+bcX0ZESZEYGmUIlvVYpXfBFE/yySvg+AAK+W0
zG82sN+R9/3UdnIYRw3b8ZM3HDzZkI4nvjZrFNytVNXgEqSFfix5afpV/O8ShXW5
PyqAB51QSCsjok1bCiE0x+5Gj80JsWlEAIfjfhBc4z42rNOxUR0LieVnwMwJ9HWu
4gZD3O9G2uIpxzqTbFN46p3iqTSHTFW0dh9eLzLy6WdMvp8nucOkEv/YMSTV7G1B
MIqdJy9YgVV4fL/jZFuAIbYGOgb0KHWQlAMZe05+MoLzWo6HrH1bxTxq0NFS+UYo
47aQ+EjdNmwfrD4b9lURB9qXL15Vp/EFgbtKtXl9QsEzrUG/wqYFIH3lTgdkGYMJ
A/LHUDghg43VERST+pYH3ZNaMe3l7aSgmvWoiJQx/zToAKtAjUNWIyQPClJFUcBI
doi6bU7eOgI3DLkEzobvA5MwcNzeEKVuhRZUgK4mzSHi5LSj0CIgNAJD+OA48obN
bZVx1StGcGPN7rP2Buu4HovAB3t2NmA5oocq1cxr9rF1OL4Cn3zD0Sfwg+s3HW2R
0cZNhV+RfYcFa92+661mxMe+pSJFxWwEvXRMBZnoAhW456Mp3xNE07P4A6DqImeg
Lm1JjVJ41RyOauAUrulqhWVru8edJJMVlgPomJUf0GtuYgGWpenB+2rVeGhcNJHD
S2dBiH/lFlOfY2xNXVs49mQpexM6IwqUmaTkf4zAj7gwaidcsntw+JT+spTEhx1B
aGvsbssOj8r7YS4Tk0pj7AkS3Yh1O3mN7ZrBm5/wi7DkYbvvFuTk/RKApnUpcTIa
JgwhiB3Uu/02E0FfDPti6gxVx8cdNOL2h94RrcxJIZVEscfffgj71c0NMy5A9KqG
VKLtOWzcQxbGFkunLWRdBwN5A8IyxfTi6Nbn2UGoiOgUgbpbQSCXDh8xHqGm4XN5
G89VqqzB6e1VZ/2fo6xFx286/l9o6FnA8erC4/GXDEmvidUii9sUUz8zO/Xx/v3f
xcfKh+AaLkkqt4DdcquV0A062HMjBnpsbh36GgIFjHVd/8dEcraySOAjYMqMQtn3
QyGrdQz3pz6Gjx5Bjb2IzWRmTXycNW0h2B8qFmjQZSw1ZSr8KVliXGO5on1YXEio
g35J6BFmMW+IOx4fQoWVgYZjmblZn0k3qgL0r1pQYxWac17Ub+jIFIsWR65mqVoF
xJc26sLBj0TP3RNX6xQucf8mpZ4iEtrYVMgqsW9Yf2SZ1vWvSbJkeQ9YeGpgBbcC
ilT708zvvqXp2SE10ptmz5eb+F95sTPWkDFjtDtVQssLXBEkZV6+OznJnfXSAonC
hkGF6rAkJMU9p2lIROAxc9KftFaMn3pubytQI0RkpQAud6BctTXNU8mgxmfESnlM
+BgtE8jPWxP7UgvKkuiXPfFOdDfeqSg0RAqJMf7B4BOYenqsh1UmHMMYqMgAOgpG
v4rD4m/sQXRLJXzn4fn6zHzPgrmw2Ij2FBBaAwQRNBfyME9B2hsxM2E4TUp8R6zL
A3zy7YxughKV/VtbomZ4tWrQ01Kck0N25FMvn+MWqqTvyiBEzvsZmijcQxsTV6Ef
BR8bmZr6NUA9cl/fr89nPDkW2QlBixkUOgv+iHAcYeoDZGIA0m1hKogkvdii18w4
fEy9MYMtH5YWCMGiE/WDjg3F3hCXA3qUNUlhM+Xv5NANKufMImwnGTpdr7RazJQ9
ZdkhvQ3cyIA1EeqyjK6gOyHGnZAPAThbi0i69siMgInHy6Zis8ndQVYg88993iyE
EvYCdaZ91NZEr6SDa2e526bcxMh0VRJU+mAeORufvb1cVl/qI09lrs/3iqeP7Z3p
f0Rm1sLA9loHwDJ3YZw9RoIFIoiWXOTnadRejcjnAqfc8kD9k7mgIRG5ZbZJNjmw
vbeM/1ZgtWE/iyKzqUNVwdj0uzDuNkkEvRVCiZHmZAyoK9Awl84XRzkuG3F1IvrQ
CwkRpeR2G5Hkp1aH+JSECEboj0yCWg3LruwpH638G/35q8rmgkYCrRxlX4EPzm+e
KkKZIdqZMw33Vznk6c+W+5UO2/MsNl+13uE+yNhHuhPOrdtqxisnJbry/RDf95VB
Lue8RJui4eRficTW1EmX1NCwVoQm8ktlQtYovyuiZyqG8yJPNNOcKmDjN8bJrHmc
XXuWAXnVI6SYH2XcB7n3Voqt7g/FLPdbObonLlxrEQ8l3RTmPjO2DCtNQkQhbzIb
vICEtE5Y3ZdZOrF1/IHlOuDKcjohB0loLARwzWDt6XbIkQCOi8l1aoKvy26jeDAg
naDQn2lFicnzh/vKF0Hm4FQl1Vnz3B17fqSTrbV5Vtfv2NdaJxdI6H8IVEyefiKr
kwf8mJSP4UowOC28wa8gUDj8KtccNeMCr7Lcw/O6gGm6NKxhEe7aKwOB4t5WvGKv
3hBV8bnoaCMddWmYTeZjBsN6FXicchVrlDqOSd3/1fo33tyx/x38dAlRjHSkMa9b
XKag0UhrA8gxnG7l1yQRJ4LOdCzzI+PW2Rd7xsB4UFqb8KyFwEj4o3SJHQBY08Ng
IJY1ZuCmfA7w7Cino5FbjoXbCh+razxPlwyhlOXZx7JSwxdx4FECcHS8mzlzwzkB
OO+Ra6EsR7morpi7C9YraiCBVzB3basVzsS9LD/XTy4GUrtJNp0ny8b0zYDu9nXT
JCx/SNd1FpUSnxXMvuADD2zKp5GiDIqOeRdzf0ZlFbSkmGFQqCCB/STz8SqAM8CW
ZWcsZ6NkWV6ewmCPdWCSgM/ykWesD8kPwXEOllfpU47IIysKBf9eGfcD2wzuUd21
M8Mnr0TvpSWGxbG8iQ+dy9yTJdE9O1MzOxTGsRUVe8zEYVdaK8SKzjE/b0KvVyAV
BF535TyAFRic7lGiJTi9ioesqOhdXTbYzLcpB0aTarFCaU0n+nj4oSYx5B7vVeVL
M80pEMURraP8SqZ1tYq7UkfkAFmTr/aFdhetOCJNrJG0jo6aR205mPC308gjwPMu
kx+dvMm+o8IE5nSsQZuKXYAM+cBDB+VlZ80chDvLD6Vj+WHCrstXS5sJKBomVQBp
BBeEDB/+4vCdBGqV3ad53lgIVPmC5fyBm9oWhxtf80X2w1y+fHWZImFaNojPJVZE
SRjR4jqt+v5hNIpBz+aWt4y7DzK23ZdNe57rh42+h82P6l6Q4FTb175tk3js11l8
K4PdVL8WKRVV4HNyo1XA2Kqf1dFUFuJA28CWZ3PQYA41xo/8EIH+Nw2fnGwzzGxH
iSfqUEthYTVZsfhiMeKRiLOWjs5WV6sm772CVnaocvMCW1JavvnvnipATkNQEtiC
Yln8nwjavCO2H0nIw+cOfBnL7F3dktDjKNpArEPRuMZ1MBovhD4CwBW4BfGUe5f5
72WRG+iiSwIgBUvMGOUg2GtFkBDT7JjTyQvhsmlRA9psN7pNVq0ukP2FRjxTxSmV
tcXYLn8qhpK9ogZZN/jQ73nbjY66/p7KcOizEraIKET2fZktpAR1wKykQxPXcdhM
B4oD8VHy0bykx5wBYxZj6UgA1b3G0DfwCLt/C5NxSkyF7/vca63MEjonvklxQaDw
QsMZya58++Q2sA5eG+keHpom+9XorEUgSeQy4ZZ06ezKF/WfzGjjuuvoqO7sVyGI
nBeuZMyQfWughjACp/k0kqgSdrSJ1dqcHkyi/i43UXeX6spYkL0/p+xZTS1NV9tc
3REwl4/+RqdtGjqnQOcS0Lm2Set70eGnJkwdjWSLOpGoPZYIS9hYmeh1ZuqhQ6d0
zsoy15tM2g0A/OyjZT47tn75zmxiQxHfLiaJGZnOq0lc590l/atlc8oa0P57ud6s
2t15Ji3t1YpbWujng6Lb0thVRJ0jW+eIOSr5veoXvBgbvmFn9eU72gq0O9bquUkl
wPfdjr3uqicRU9L2qXnErP7biAJNLxeSgmrBOGZSX2LIHdZ1xj2uijfvC6TfgiQi
g4c5Goi9T+0AXkUpwE1U6SxHr47YZPCji6mYLNnf+aQla9h/ZPlvrB5wjJk094c2
5nT9cHl+Ji8EYn6J5DvypKz1DhpmalWZhV3JCaL+KPQC4ZlwhijuSJbvEVUizkg2
Ln9QbGLlMdrFeXNzl9jjIcQ5mUBdgDRRSKs1WP8UsIcpWr4QBD5ilh0XJ1muHGVX
9GhKIWGscPgxiga6etq8eMBwDe8/k7JIw8jt2HEcKvimJ8+wzT400NCIyeu8WSPr
wp2WwjYfct2DHBU61+1ifuSyE3QEtxarzC9ZW8M9o9uRkpUVpyZ+LC1X/Ndip/Tv
QKvX153NOUeNw1BmO555Ar2od+yUAWVIW9vg4abNTFAH0B3gCXoJqf39cJ81ffQA
R/Xe4nfZgHIB0O/hhOjcDfyRNzGeAKXMQuM8uXkJNpu+vDZ03NAGdJwJzZGj2dN3
W/64UR3rgz7QvhQmu0ztjv3qcwtiDseZ8Yr8dtUwQNTdB5AntH87C+V0U123pxhF
nwq8TT7uZjKsIRTzHv13XZ8tpXh6cFqwcOhbnPdQcw9tqlEXQCSJ7JBJjfKcbAKl
/wO2I/lOHTACQ/5Ocl02gymEa0gqOZUa3wBOTUhysvxrlZns+aAhrNWJlHm3edtt
gCbrMd3K6Z4n/W4TPOmJa3TCjmsFbkhj84V9ChEinUsu4WtYZIG9FY6ioh4sVFhK
rdU7LvRhEL4C7ne3u0w0FfXLncH5Q9qwpnJugnaOOhAnJuM11R83VC8cIi2/UEq8
toubI5tY5A+ZJuGIJuijFe4vjDXerOtIAYoyrTiXkYTeKzXQi9vGPObWKPWCKEzh
4rKeuBR5ax3PTbeTCUNPndIlufyLKIWVhMEcZXy1zGNIRxzJXNfGbY91CMdcKOHT
4yAaDBFu5HbGodkAgrrOUhet/g7rRJzYSk1aLyPqLyGhDTNt2zJe3fClMl/GW+pM
YCOVQK2JZwmr5n+urLu7BzRExPzGtT5qr8dSIxUWqmJ9keJjPn6r2+Pr3yvB5988
b/Nj8PW+ljtiW6kexOvBmRT7/f/HWDpMA8J1kBJSswVFxMjesY/CwTihCKnljKIt
ohhlpypTIrNebikzBrJSY+pMClGU97O1rBQwbKAPJTCQkoEZ1c/u/MRkBzFPm4F9
F6H16dboLLoiLqhbGVO0KpmrUHCkUaVrJIy3eyPyVXCl3DdO6/DLdY8hiZKMBagP
tqHe6YRbe9pFgZo94M9Zig6PEXcfw081FvmYI00gs01qT7Y7OicBmKHbl5A/nRxa
x5lkJrksKHGkYJT2gxOlVsZBOOPC5Zl+XgHfF6js1h0LWzRxSchTvSvC6FCCySOL
LUgFfrCZWsI76AMUtBLL2l8gKztOWh5MDpDadETRiczho5eVlB9cT4/XDEStkHfo
c9KOFeb9EtKjvOEeLOCGdWelT0VgnrUsQGJ6Xg/VWmaLFle6v4KSCf8j2vXlNiY1
YV25XhZAxVRUk2DQIlBCryXpDv+Mf9Q69WVg2vayNlYeQmXcssHoaWsCuzbu7tCh
TgZoOX2faoHFeQDgnF9GXoxrfy+jVdfuadiUI9oNSqOsIzmpShKSbp/6Bnie41pp
sL9Mj+A9OI84h5SP1gNQX6QzvvOHG21mRLE08q4Z086ExZuz3WBMnOG1/JGCN5Fd
oQwLLFt+6yuAMci6GZ/HL6zHJyRaUOL0pCp03hc5+7GhCQ5cXPWf2K7onGOtACP9
0bNWsoeAVXjWbIBL8LXyNmxuHnmZoA6qQ+TxbPFVFcPSwNpgipiKSP+mybYGQ0R+
GDV1rOIon/kT8TxAyF2xzXwvfVI4KVR4Pyn/mK4ZKSJiJzU2jk1ixZ0W7l2ywCsl
Tly0rW1mKMmxfB1fYySp0mEySOhlDJzwmoKwMdAT5teDYU8LVIhMzr4phOVqQQ2l
glQOgmjga8Q3r5JTzcW4b8ujp7xefLn9Xk4MjiohXj6xlqhMBe5m/vC2bbNR8BG1
gEfaWi/5GxYUuSbAqSHny2ykIV7z4RqT7B3xrkSK12woz6CPvxlx0Wym6QOsMbhp
TQfiokVnQV69rp3ybWI8X3fdDUWNM2frKk0ZBPHv33YiyNmDBubgqSUiWHIzz85n
zsv9TE3RHjYy4RljS/4iFAfRZFV/5MsBzVQ0X1T9YaYtX/tfNdCLXdf5a9tED59W
w7zAeJ0T88u/+pyvleQbCMoALLzNRsHoacY5Z6rCDNspYyzai2JmQ+dcoCHMmXry
ey5sMXVvqVaHT+2P50wnYq6IVfp6/BgWR2uPct29u/0cxL0utQydgE3ZiuU4NhFJ
2DqJUXe2Zhtwcg0r2oz8Rgr6D7XHcvhLivqs03+OLupyOrjG9eTvvoGkX3ieAdXD
vuhyYy7wFtDjQb2RlsU3p9dLaA4dhFvEhmcwmwFWeqWMNxeDlyvUIM5pSwg9eTo1
FHIHJx+9f99MUYg0bMbcX7casdnmHKLdHC2QeA+Wq90nKJuS7OFXsCaqUx93p/Y1
d+G2l8NyyzBjUpW45OLQJOLZpr//jyqD18UpWGd3+JBNLXf6KiKj2REhwm0R4i7j
rCEDq4ustt8acYo8CgOJPrkwu/U4AR+qHfocLBIaB7IIo9LgCOcllKGqI27J81mH
1mv2PMD03MRXd4rw6iwovGjp9MB2p/FfvQKKazKRlBfUT+7keqBePGBKB3akcWh5
VdORhlOjtvRx1wOeebvFE8El8VvH2HCoZP1KyiPFaY4NELxQB+z6z71Y6K8HGfST
9W2I4yb3llIG+NDfbL3zFo/RDxpMfwg5ropCJEPuMk1i+w/TXFPP95uqyhQmN3BP
3DLgHEFgZVHtI7XxltMsDl/3hIgwwkN8zQO8iOkf1daZYTRf8frcSY0f8+hVx8dV
ky0L4VKSvWmt0ywQUkNU3tfNSz3zAnzfBpxPvEn4QPdtqSh1M10lMJy3ntq0gKyl
+EU6F3Ehi4CSmQ+JZa/xW5K6trD+zPFqnytpWkcawM7YEYk6AVQ1dk7bYCSjA+gM
vcpBXRqso3o6ZhUUXuj98PQ+zOVALc+J9wBBWTuXw0/OkL8ZdXCNTEg+rHqVXVVe
9aKdfrt+OXoWWb70MtGR7IrXlYEE3fI9XVm8Jbj40GRenkF3xGAfa76i3Dqv8kfR
HKhi5MjaaAK5fkMALT5ZmxRtG4dj2ytOpq8jiimTLXaZoRxXJ/qB4K+7VAW1EqZ0
cy7EOmJQTpU+0bu8Z50yXE1SfkNnt9srHcO935U6tS1AtLuL9c2bpyE0vbrvw1UL
tinwm+hpO559CVZ47RyeRqV/6cAckSajX4OM8F6zCK5poJD/ROn2U+Sq4v4JwJYC
yC3CMnBGPQ5i9MHJ61cFcCooHSR705mNGXBqHCFvjZ/RE/ZxBur+twIwhWJ7ui18
iP42hMGl3i20cFAEnqhNQsSvLrsRgRVJEhKZGh181jnAaSX7U/L31Mix0qVEsWu1
JiyXtpBx5PzyukVDaNDBgajGAVCbyegG3fb05fDQNrCs2tURQ1WtTjTePm1Qkjtk
8f2lANbZnP2n9D4tIQxWNNPHsH9KijD03nvcJAwH6AfpJvtRETPLNFWQEVjuzEud
fBvoAwsMxDuBqrf4vM+vJF0njJJrApmyX39GrApL1FcPQ56JPEVrs7Aa5X8GRrUR
idx0Vpcfsjqyaez89kDDlB8xXfsuafpa6GQk2CqlGfTdeo/mkczt96Pn3TpiLgRl
7U+jL1JsOvEs9gjhNi7PBWbUoXzASiehdMyYlFZ16u5yESlyxvyCr8fESE1BLeQW
J/Z1d1UeqAHEEfjnUlD5MhpMBhdPH/v/1trrv8MEfSRak8HzP1m7T+VG9Lzffxtd
frAl1Xc+aMrusa/HXcJDPbNY+cz9Ny565F9QNb3RH2SpsMnpqR3nJgr/FK36k2E9
XSSYxXy83btIDCZYmmi5n7RTB5ZMRUVeUVzvdZ1R978rShQ7tfqEfpYAzOCbwTRC
bP4J0n2a7S75YUSvPRiBnoihgg1vkh51uW2eeAgIKk80twPMd5qwRgUeMfPk4ijX
/2o4fGxYpu/yvvjatLPpOrY2EzHR2N9ffLew7/ZyfoQoDlEmz/eF+6c0jGWusd/M
3gRe0hl9kqoLf14WBmoLcO0Uw5cMhj4wU4xn+wI2D8RlH0JHbMLs5aCZQiPhmSeG
R5kFMsyp70zXLHT7GRcgeorUuGR2oAuZBrHKRkRXFQc0z585UjIIj5Dx57uec/Fg
/c1fWl2ipMHLyZhc5a18NrtFmtu0VFGsTxRuICWNeyCRK4Tt2Ec1jZ15hmy3Vzxt
4C+T5R9RgGFoNPhuG67yycxkSrjr7pN21CIOGjk1Km5+GsyA4rarcixlcaL5M1P6
CqUhmyHG1q5bV2OVsMiYjqL83REGF65H4hf63Kc5kVRLJ6R0rg+4FIpCZShN+ACv
3+SqpwqV1tuJ+bc+iudc761dlZRJnWiEn+yk/YrVxak5yYrbYA21fI50acHnNLtf
5nNPj76wCScepEEdMXj5h6CGG3TKOrd2ZNBDf0TqW8N6bcuNd5+CNPtVQk9fEcg0
3HRnVK72vv7aOW0gTC9DKbYq+JsLFn4+spe/1mhcHt8aWRuZnpv4JPUVtqsAPkw7
S9BY8HUjnyGqVg07IBuXjz3ZejD/ge5e8KLuHgALAzsG1fx4t1ryA7Vt9QOemmP0
SoOQgoe6wdXpNn+lfwr7nvhvWPEWn2nPdBoBNAqrYMCZL5Vh0/7owc+QqYx8Eo0f
KSXI/cAbaS5nqKbKw50sDdZUYjUeuPyj75xX4stNni91RYG5X7j9S0RwLMo01EIu
PBYhcN9KGylyRDYDwH7GGD0oFSWkORlHpF7Q1OYfNUZwO/myPz2L8W9B8CYyCmIi
+a52X8xsyUQleYrJ/vX9aC5yt4QVSwydFpmGdC/B7YQi12Q3cFUhzFer8JB0wxL+
+5dtOWYD5SEa86XM/bF50WFGm4PQnU6K+i3xl5TRgY1n19SZcMdKvh+8JZU6Wka9
NJvaShCGe9fk5DxaLHWOP6S4QilPANVYo1Ob2bxLnPZGqzlx88B7OroxTg6OM3wm
L6D4CrHqFhgHm1Jyu0UZZHxQan7Ui03mgSsSp877T98eZTq1Xy+MInE9pFjKIARH
B0H4w0AR2+cURKiUO7zZQm4WELfhoTpIZaE4jSEPtqRxoo5obvdgQV0zyXVh+ThJ
TdjmaGxrxIivdHoUZiNJExLwEUQ/ug/O9qkkMBvTloISEzVg1vAYbvb+Mr2h4PLS
DPNeD8hJmHuca5a63ojPGr9pvKZ7o0iWz6kDL5eDa6hwC3fua+K/dps97wk6Nrvb
l/QK5s96OLaB9sV5poSlI01L/6EF999JHDck7VY1JATCR1fehwUQpgYtdNICxWMU
aXpXxdzM3bcLJR0+B0glCCje3CR+fJflpFom5pGqI940cHPXD3NgdjCh5JXC12ua
8TwZR/jh4y/fWWIi+JsYv0mXjj6sFXK4YY+g6+P7W/rez2qbii5QDnKEIE1KYBZh
3ResWSsdMl4K2UJrZBSJT1iHKPiquCtzVXhj4RUQv8yXbQTAWRRmC98B7mwo1UDm
6z17rbMyMGtFCnBadgTnN2/g5HRgsRi8Cts6zL39XY0Vchqy0I9Y5by/ar31PLvU
zh2h+PzuQv7z82dHey7Gg2KVFkZe+Ok1y5c/3BCA4+hkS6EEHYgEsSk8R83fNk0L
nGyPtOqlbZ1tXbY9O7Xnmrs8g0D28dBZsdElSv85l3gNm9UKZPIBJOtJxyQ/EdDd
DuGaN6zg1Kh8gtx6Q+Lf/BuDoyPUV4GddQdx7thpHgehXYi1YLNQuob6C4n919s+
2cUfZBZjA5EB9A8MOd24iWN7Gskw7wMG90LVKNvURJgoGrrzIhEGU5DwOSebRFvN
5ihIvMa0WyT0LPyjzeg9n6zg72KVQn+5VaszbzoCs5ZmeWoQabiN8Au+0X2QjY82
UofQXFh31afgi/8B+BONR7ToE8M7HvkfvQyZBpfmE1xBCiL0kYmQtPNInjKQ/Ajw
ltzum8/dznlv5vsu4ep8oBUGlCvpZfxZRE4SCfJvjB6hIEJfuxju6k5qGodm+aGk
33gKcVCNRJCbFW02DG3HfaGJNbjjzWsUlAlH9I2EYwRqmh5a2kktEuw6bXfLqkPt
jzcLyRNMJ9hB7I52/8RqjrZd7GMd69smBjtNt9ze+lmVFP62IchXWF6dv1SaryKv
Kj5agfL9PNtDWsRkN23hRhahoot5s5y7X51p6o03/WVDuH43e1L98Hb55M8uMGHA
hXXB3DLfMrmTwBz5y3LOMSD6z5ni4DRRKK5bGYJnjHG+MfYgWInF/iUGFNNHebDp
qMyAHwHDPoXUdJ6iGPESJXViGRb0aTMs7FVFn8V5sYjtBvNUh8HqAiIHirPMU108
Coa6PiuNHjljQ2Pm0uOAxvfUINH9QpvNgtL4AwScdftxQ4JcaJ+XD34fCyyiUYVY
sinyONVp2HlY6l2d7Q8EDVFukjKY4kx3aGbLVzk0EnhOdr3dRaTNaDMFgOXKrkCZ
GDspNXlS69JYyWFmPwfQJ0SObsQFJJqbcYaNHmGweUjpdlyM0f62ETQVO91zUPCY
vnXApkQFTnTYjixtQX+b0iRUN+AnPY+sSSRjFwn8RLhIBVNRExBNyJ9bpxmJEFxQ
5h0W9tb7uOgLgkm+t248grn0Toq3c3sR544wVcSSgDsYu8MPDnAOR0irVD9/KD6g
6Ad4cQticjLIiAKyip0f3yP/GsU20pmodllVCBDYLRJKEJ5GOuIkDoxLyC4ipEum
bz4Jzt5+euvLThAFIS07Udfg2gCOnpGfuXfMOVMlLDmFKNaIhn6tfVksyK2gCSlz
bitR6Y7D4NdqVWS4Z6XVD0lnG0jrWdutg9WiSXHRBQEY7DxHca3xfjPf7PDEKns7
F3RMFreUS/GC1Jp1YeRD/NxRo/5sAF6kX5dY6TkRnAitNdCCtRMnmaHSAS9NAPf9
gyR93TnSDoDQqiyGwr7qLiL6kvabXUTq8QigIm4hhmOADmKwXZwF9oisaMR+JAMg
p7s7oNxavDFPX6vifbAL+PVmNlwtPq2E8rtfUHX2TmWpEz6os+aI005QF2Tcmuyd
jf7OfvRlSyhttQrh1xMGoV3GfybLUWxs3FtcF1KhkRvrnSo/IxHHrIpIrhR7bUg0
vWj8bw3t43rXFzmg9u+Fmu/X5E4SgE3AU3i/KKOLAL8YADX5wXH5iOgaZid5NTiH
hAKO85zCgTeLBCUnSRLQ4Z8AYUxSo2wxxqUnr+LuGuBXdyKDIy52IrtiyoWHD4U/
8SoVPswV6vwjGRYHmwb4Plj+dQM22/x5pdrYvNnBO+hsu0Sl04LbaDiN7srmP2/P
h8i2oa0+jbWYD8B1Br6PuADMvJj7wJgT4QxsI54Qq1BnC8wr+ylpBObF/2HlrmBy
hP2tUOizTP6PuK9tBMDf65YwWTVBQD0sCqg6OWN+jCp6qSbKGTP3M7syNJixFHwX
QdlhrKFq4R/QtKay35WRGoLcjxQK0ApuBwBqCO2bC51F4Iud0nb9goDwlMQtpsjm
OV4IYuedM9pjkCu4mdpQHDZeuWhQ7Alr7Vld3ePYA3jg2naNZpwqAYWqLMFv0tam
vrqGqoFuhOQHwmp4mLRVGVhmTthPsWW6z+4awfTYPq+d0aKNCXvkeQdL63rbujxO
b8zgap8ly0X2uqBtR2ITnaXpRAQscLFRXkE8Lv0mhe9YZt8b72KbVYN3nwBz5Rtz
NoxkyOgl0AeTw85LrDxge02X2SHubPSnRCFq7ug6/zhYFrYkGr2BP+f1iaxUP8b4
Goth7MzTEGSrZKmlsmt5vTwBU+Miq9jYn/E2Kh5wu5hr9DtPUEwpoXwgpfZlQ5kG
6pnXb70vPbyA3HaY6lS9dy4iv8ip8ngbaRNQ0Kz8eP8qtRmRRiSRt2Q3F/sQGG88
mn/5Ms+8gewjuJlyGoTFE9ctGt53bMjEsjZO+jaqOf62aSxRdhmIa3v80rhgZa85
NVhGzZe+pDZtq2geVfX908ahPF7pFUYRNy0k2TaLh8Id/z0BqiX92diwLlebu0Ag
KLCnU2p8bu0ApAcCKId0LcbVNIIkdzt7jCBBoRIlOkmU3CwcyeZxVwmp0U9T6MzJ
hSm+scqBsVs0icwJZpaaGeDykqxAPF79FwrQhqSYmd2SvRsQ34F97jyYV36PP2jr
s6aw3wYQraq+y+p1QoaEalB4h1Wdn41ZnUwRuybvvaEMvRDyLZu2cGeB6IWByoUd
yM4QOy+dVmHBc6tzqqcO7561RMNdEWCDIEnQLynuFNGuoLfcyf29u/V0dVuDXylm
qvaPvQXBLUhGIrC8f8VLVJtkJ0WLOo+LeqhwYj5PMfIt1O7dht1KTxZCTh/crsYK
mvT0KBVs/yzvQYmEcUrfqKBhd9vnRE9aZaPbXbhHPLBadqTlr/bCg2KtK4s1o7rS
ZDYnjF4Zo8FZTJlBiS7BihYri9j0DgtXrNdAA8gfJS4A7azkLgYhpEs4rmWaOB2w
BjO11sF+W+3vq/b4YeAkFK1jkO4JCCbsZe6ftT34ho5m2BWL0FIxzCI4L18kIy1Y
vXYrvzZZ8AmAp9RUVHgyKb4XZDWtVWxmobMptejRvrredByTQSpAds9/SG3IZl7/
UU+ecAlHnDmvRxnMmf1gvd1zEFappkyzyk4V/c/ueGOSS7woezCv+AXVRC2+lWvB
3K732Qa9sOfk9DDttw33o60BqdsykcNj5iVHmLBS+0Lgh0K0+XyCbs8xp7BSqdEE
aXuxEv6RfRwCg8DlQKczTdYFVgQmdh9P3kIETjeglwYMFzFk4/jScvir47UO1MQ2
bnQBeS75qPwLJSMfRtRte0cpPTpe/HOlQMl3LUp2mu416OFfupoe2230AwDjxIUB
RuukxbkUnrmf20H9iTPfLjqpVEijROC1+M5VGamidHbf/qPFCvpa9vKKgmKVLiEs
eMXu66R2EACcON4EzCgIjfrBvzGGmUi0bU+eDlnNlpbIyGzRY340dI5xATatwQgJ
dZbhjWJHt6VYYJIVrK8tJ+O9q4g9EU2ozyiDgcbAIvdpXgd4sdsulpoQsDsXrH+z
CI9KAGXQy6UTdnsp5B33hfXiEvJGE/oVDUqeSVhvzfx6NJWPweXD/aJn8FzQyKV7
ZP0JpXb/3vf1RifrJ8SNdZkH4Uskr2Se1WMPBGQnqIUazhwWXJQ3wMHqpDICYK6Q
ZM+Vbh9uAxK3aaOsBfy9DHD6O+94Jd1S1/8Jh4NgvgXNboImsQVdRdDfojoGggWO
iKKfkHo5UixP7U+EDmsiBeKAqxw5GwPFp140NiSnF12mygpYT5Mpyk47dUJ3jmdZ
QZso6E1z0iQBET7WJHvnT9+jT6J+2wM2gGxLqV9vseC15WaKpo9dMsqghxKRAtbT
1Re5PwmcfD2en7y912n5E4CWZRBxe99gdWTWCmCgQo8vNJCCiRMdvRN5NhymLXMw
kV/zrnzmZRpitre4I9c/znC8a3rvvf1fTq8vJ7PwDKnJ4fkPQkEg44KMSGTM4MR1
lb2J5ZtiXpKfqpxo64JYOUtXigt8MJ0hAHXuzpnKx17JmwdZ7jOvKU649i7kAaf2
8quvsGk3u8hmXjF8rtWVrlumkAQD/F2ZdYMGBm0NQEPEsURD0AXw+Td96HZlAO2T
LUyFlyspwZSs10V4Jt+3E47I2/F8M4Wju5Tj5cps4kvpiR+WUTYDPRZCvVY4ePDU
zx1IPRLKhUT/+edXz2Hzk038wKaSuKvrFQIHN2D9nAVy5xe/RRjDWClWInFSLnFa
VhqAvZndDCzcO07LDkj7u9RVHQkCLu5lEPW/7u/TArAhEmf5q33P5BsrzzG44DJy
0yOHXkWtJJiY1vKucMANobJ0YfeKVsWjeskOZMzwK0tbXi94YsiCxFr0nltJ2cFv
Ct3Fm5px2mSTnKIn342iJ4e5mVDBikjlRtoljGaml+gq6KTX3BXZoywLalLooEcd
P2zI/U4BeNAM69pIgD/zsttHjPrOPQMpnX5w4R5dlGOocn2RQJYgcWQHJqG8SyxR
T0X/bwzk7F+aQuOkKV1qf+7xFsTG/XLPKQlvZ4t5QzMUQjZWJgEXJ/kb1upRI5pa
xt+4MsIJk+Kyajzt5VPlAXMtURkuMYReH2aMtpoSsjX9RHJFSEVEorIS/EZ1LiGG
3oge3XXcSfpWbZ1J+W+FROz+/bk55GGs5NkyucvPZFk/inZRhSHYvcGKJe7vW1Yz
MRRcbuDAkmXSnUKqt//GuG++eYDx1CEVSe6ezj61hIO0eYKt0jwG7aB5Sv5UGpwT
Rf6cTWHBRmyL5KGXA8q8DPjqsRTzIiWeypwADLJtdQBD+ENK402r4ysElgGSP+D9
dRRFG55mSZUnyScpqZkRltSyvaLno2egABq8js2BU69AX7Ix/dnLkx8F73hrSaNi
w/0jXPa8sEeGnCt9YMZYMF+talkro1g6YX8SLckkjZdV9JyIRVhME3uDBhGRXF9R
A3M6OGIxAzClGcuX4mgD2Q5NmhMv2vNXAy6iwthQ/PaGIVPR2aJy3kAfMgyd96lM
ETNYa/jYWpjs7HL1AZGWSW7XUVClj3U/2zAOUlopu3uRgPlp/awsiGrVkJ5Tj9ZG
ZXoVm2tmLRAE5gUIYe1N4IFnt3GaBpOrhWPO7DtlY3/l2q7bObPCxiHsQHZj7g43
MN1Ebf5A9cH75jRv569kEN+GJoaRz7rVPpkAJ5fn2bp15YSjazFYz3FIO4GA8tJc
NjEBIZEwucabJ+C9FYB718rpr5WQl5KUESP6ymhlpZARjWGJ+yeX/FmJafCe7MUH
/hcIFZXoIxFqFoq5aztEZX+OPGOzViJ6wuNj+HGACcEVFEjFkM6Dyx9izPC2IJxS
j6G1eo2TrEph4L/mbmRViXDo6KnO91IfJUAAsxo+6G0QVTj7ulZXjJdFoI/RWpsh
AtWHMrbzRwACHf4x0/05jPQbdIIu8uMpwwwdkWinpTKoPfT4z4+yP6WeSo5BjfZ8
sD+cn+wFmjVcTAfy8CmnZOwOi1ziL/Tmn3muW+kWmHFFa464TsQC1NVCM9gyrNLh
dpkHseyjnTGyBrw9tOia+tG5i9sDUI2FXP24HftAvAQNrXe0lxNTghe3qN1heLhy
uxD0IHACH9iyxLsNFmjygTcPbPt59PU+peQo72mc8AinbOrpZyDdKm9NTvKP7JtP
isvmUM/AmbOgbzQCMW4ayNowYPH82NQuTz6B1Jg6kL4RJ87mvG1Xcc7ffiOKO3z9
MjhpPyuLBp7BDj4qyqe4HBBJG8FxFGN6WgzyDm0AFIT3FX60IVG5q/4eqV1+UJoo
Z2JJ5iC2fEdGYfvdpBh6m8RoRTYiDaiYlG12EtOwmIf0tgoH0GX1+WxQ59/lwpER
GK+24GOnizyDUYOOTMdNUb+UjXzX8H7DyZxnAyLScX0zn1LvWi52VpkDtH1Wu6mw
2/tBTQlX1KWSYW3gIjmoUleQQ1RBV8c1s7RZE/akdCrn5XSkAvnygclKMhQI8GFd
O+nGAC+Nc5pSfqPBWwx0yyruYlBpcPSQaD9A6ZXnN9Z4PIEBGmfPRpSq+trtytLN
a6Mkn26fiaNp1urhL0l/rP/UoMwd47whgB+JfkeEbGXnugDbaRs476RzNEXvAU1S
hSEq+GqIm8hjX6KZGaBn29Z5HUc1y0K9YOfmuwS4ulB/jk6+WrmOeP2fjpvMLIM3
EGBD8L26pI7XnoHrp9WW7ZsUrOWqpWEycYVKs3F4SfzkQgjFxzZ1B2EasbLSg3Fg
JF9mrUqmQeCOoD/TgshUjsHTkbK6zoAXZrRKBRACe194HNh948xKm5Ql7IVZuxSw
5fq61JV6JxB8oLDiSl5WZ0dK1EmSjlYyHXEJheEdASbjneGNruhvbJTXzaUHbvV3
qZuTvXV4cc5nI6tQfURieSxK6dgzJC/CZjpyXNcxpFZEvNrF0lPQbDcVZJqIy87e
zUSKWzgCkcF0K8jbV2cvCDMfMCELqkyiNQ53DjRuSiy+YkTo8Fqv84PrWHdUxBte
2wKetUDMygUcf3Sor4H9kJjIdwYXprV3IJjOtH2bs+Bu5fqys4DFEcQnfWqLAV7U
L48c1J5K+NTrnChkIoVraZXzNdl2loWKVnCXPHZAfj0n1hA6cLST/td3fFa41z1X
HOTv3J0IqByQh4GoXCTYQKLI5rvjt2lzZvgcWRmp9fJuT/QrfYuFyBP8KLs9fN9u
RRtF5kTV9bUPZlJjANVAp9R1lObg6w5/hEwf8btU3Zwn1NoXuN1O4D5mK+lPmPdK
SKOuFr3d8W8bMRHqUzhcy8lAxZo/1OUnhV6d9CKJVEdWbZFyPmqgO7/Wx1toYmYd
bCjQdXXx8tr+btJV82+PglT3ZHlbdTFiAKjS5utdgLL2MkMBSwY5FM3PuR/IuK/A
mg61OUWLT8D7E9R4Awqrpc2ORlG1pGqOM/M8ks6kXYy+PH/+vHLeFKUsVys0maiG
VnfsAskG206ZqDJ/RDwTPxLv4St9DI6o6vFf8ax9W3K1wGRyagcz1MG609vldCWG
1aubPb9AAk2otwX2G58W0mEtlXILwR6q3m04vkTMfQ65vaXV8S8mZZjQg0qZ3D5c
XH3YTZjwLTFEqGtkT43dmZdfU6E1YA3yAhiGVUo1tIgMHSW7EduVktdZ9ZSzC4ST
0v/KTAzPkQ8NcUQd4BjCxtbv3miEs3W3jr+mAwvN1tGv98lHFrGYdAGG9qp4Lqch
3bynbmyBejafZHabAGshNelwlvShVfkEeMKiMeBgpFrO8D4a+u1H9tsceG8m3YBI
lLZPeGy1e2knY/IygNzORBRNrLpkLbnrCE1LXv3aTvgaOPin5RMJxovweu175U9x
9Yn7KIbgCyRGb0butlqH/qvfgkYRxx0P14OrTUt1B52L1pPamSvuGaxUXOnH+QZB
kbeARhk3+TZbd3SDgcdVlX6sX6uTOeLS+idO0T2e0n/thsoYc0fQxI24YJ63yPSz
01QtGm0KeVPf3AxInwmpO2Bscn1MR8ZrDZnXWaDdkrCous68UqYIkE4Pxlldlb1j
OsyS3TAovxdkZ5F6RBCu0WF7ioTzrkvNpFkP6GxLKc1Oo4zxf9lNJTonVuHvwQDU
mv6PelfyjSLPMzcMtn/2VgG7jk6TjxP9gjdbfRrp86DT1mqA7S57cFMyKwzPUvvr
VhuvNFoYSc64j5BO+DtVe/xQGy0pqdmPM1Z+hBfrJIb9LbfesLEJM9DuqXxIeofs
Sf40JEJ5XF1YYd/GneKPH1NhvnShI4ZloAoja2eWZwrW9l5L5KWwSDAJRTp1Yloq
N+fF37UHJwXi7qS/XPa5Zx1BuJT2KG12bN784g/qrtSpnvFEZ0VUq3WcGtJ0jNID
UGxjEmNaX072lIdL3olzZNCTZVrVn06zjfl4HebCZlk8vvZtJZkETDIUc3YudiN4
T57u7TXMgrI6amJMN6NFhUfjYqQqhu7BdNEu0GJtfrSsbvJxV/cKWCVRUz92g3Q8
ZQDKihppFHCyxYSTfyRBwre5hOTBpZu2ooBskoaz1z+dsMPKH9iR4fKjYM8MRVrU
9M9l/0ddM86n9O/tc/F/TbTkEkHdq2mXiXEoV9/QWunG5uJ3MVWhZStUj0obmjPF
Pq18nDyzivSKmr8TZT7WJPKY73uXbAy/kO6Jrl/KpX79CMu4TIGjhBWMiFTS8jC4
utmx6xBtfFQhQbjoe4TjbC7qgKB6yircfst3wvdFtUHgG20ZnivV3tGkHsTR75dS
qrtVpdoJypGApTluRPHmVWlcMlduP/UexpI5ji1g+JbT0vHb8vnNkKg5tbcGo3ux
9+VoTMr1j3K6VMEvg2A2rJGgD5bWMairyNBHJ1VdYQW53olBBLKdq+xanfL2LUFc
EDijQC8v7swcSwGogclaH96B4Z1jX69B0SctqXsBDVrC5T7fO+zmGxHHJBoKDQDV
rvjkEoLbqe2kGN3o8lzpl6v0arKX8deQzqkKdc+g3d3jeiTVuqkqXK0HIn2KVtSZ
RfppWRZqaJ28/Npl4CcwUNWqovRcwWY1fAn+xjmbjANwf5TPDcVjcr5ISMguGfWD
NdxNaxoVv8Y0N+YKfIwXFPg493hMkO4IeF4apKb7HSSScJ0+itxIncAbLrlhE74S
oZX080wnxBvhEs3lRZBXXeOHJ8ZNDICUY6drudt64b9ghKQBPQ1TCbU7AiRobL9v
4woN5q+3MltHgggYTKsz44UiWe4lOYNMOwUajIk3M+dGP01PKruoe5spQx4iXScc
HJk8XOhtxKaVc7AsVJMdFzAgYTs9IhrTcUaF1VK+p8PjE4FBljTOqMnpCWYbGVUs
fiPEoGUCueSIAS7yQHeoSF4SVZTVDyEof4u/z7GIkx5ZLdLdKslXcdrlp9NocW1S
xghKyrrMz2HpzFoCpZQ+lDwnd+7s+FV0aGBZ3j9CLDntfTfgfQ+AQuD1PoYISVFu
z6j2rricJXXm5NaLnEpk6iBe14sGoZumhZKSMRO3CvnpawRoi/4Yc/XdS4cWTep6
2XzUbYLCdqLhXq/ki+5JiV3rI3tkfkmM6rYExYrcjaUi2ZpQMc2fgCsOfadpBUzw
hlQfxBulCgOFEr/Y6sr/V8UOWn8ou2SxnobQXnG+VUdunBdobcubYb6wV14UlgRX
1CaC2deOpPuFf80cAnMIVVvOtAgrzIShVhx5RG9nxryn6TRTM4fAr0pRKzuf/0fE
4nyNVl6XVH+is5SWrxvkxaoSSn68SisvrmQdtKPSmsEeKCU2/Hm9jC4JRvMZwW9y
HkCcwH0cLVocC+8ou94HYgQVSpvKKtztZ21W5TeIClrADWd/Q0vo6LKYZNQfUyAq
2uvKYTtlum23TCd3+0KDVO6npkBZhB/gP4J1HUbFm/6SOQeXKeVW9C01Zu0fmboh
pktOl9S7tyDKLSnWYODdo5TYG0m2CZ7NH0yDcO4FeN3nwnIbbpoM+K43CVcIhyMq
Gpmro1Esxm9GqNh4encGpLkOC6LNldaOy8JAn1DeGEeyn0+uZd7dKAo+07V6yNtX
RxM9G1AubfuVxq5GQvmXz3kF07pCXvEYfGOj+4PHNKtN6DYP7baCmA1bJXbtGiSz
rbV1ByaP+sm5PP6jb1Z8Swo30Z9Zl0rKW711c4gLWdZU46lngqI1wXWXQ8JHIivk
sFMelkcgYWPp5MTJMfFC+MSdyLkqA2Lw+FBM5ktFM7R944Q/RAwzFTKssWyOd8BM
kgsABRiYjsW/WdkVOKkhyQgOYzUDJCIBhlDFUvbrTNTJPgG/96UNEh+bvB271EGS
jfdrYbO8+QFmOMJKT488U1NG3KjDWQrrBzTEXZI/U2GIZYQRFB8vQSpQFxrNa4Hh
tAJcqzeJSFVIRuPpX9oQkzQPkuysCf5A1UbWpagMWqfLGc2LH7leprSbOS9W/ZLb
x9DNuj6XbPdRfM1wOyTgdrScZgIL1GC+uMG9s50TMDCNDOjx1WRfh3+t8AZeBP42
Cyb7C26ylPP0gARgj7eJ1z2EoRvgl7cByWPd2WA9oIlGAvRk4Sy75CnbBDQOkHA6
6EfUGmK9fRlPNsF9KWsizLrhRw1zRY4UToOcOWsbbkb/TWBk1a+jZ7LfXXGG6dMX
1Q/e3WLMhh+Nc7mgfemoJ4a4xXnaWEY+VAA8+LVAtC2XKfmGQh66ThJrVkTUZKl9
rqIE8V4UsV1HYrtmNlPfq/B27ut2Hx1KH7+4aTKYXo8/kmg9L7e2TnhZHUbKZXV4
0araqjozZQumJPEmDlJD27pkrG60DZjGPpwQilya74nvvkkj4QP3RZsg73EN7JLk
xOFiftd1ds9Mk8RM18CLb+1QeSc3KSGOvaxOjdlZlSgM3blK1OZoBF33x0oASAi8
CYRab0nl9afsSuFA9kSPY1iHiq413WMpxXPs69kllnbF9TlbrW+S5tffl34bO3dD
R9gz97vkvqaZBZArl68uU+lzGH3Li7JB2HglzYKVJRKEQte6maM6DwXcdc9z4uVS
2BeUW5+twwmjIFLAokKReUUIbTINTrTwQpGxWuzHJ1T+AAeZLFzMt8Q8V+4rQfOw
P590yr+PJr0P+Gk3Mc2S/sFbteQGshKHMetcyQW76xQKt117cGUe11uKUxOqM51m
rjuGYbvjJNKhqkXmq+NYVpArXlycRkarJrNYgCNuW2/9FFoiXQEpku0NnGKVBQtK
b0J6vgZ1N7VspqzElgKm9qWsJcO9uPlW7vbpAhW5bQTISLK5NWJ9yGdhJb9Dxphh
KjEx6arB75MFM59yaOvViBmBpEfdD5d7qnqjEp/5/iZuqot56rKbywO6gy7IGC1q
i3tmI6ErTWtRSactz/WE3EIkKDHdLmApH9xh5jEDpUgGQcNTK6XT5NbIF1cr6wKY
lOOIJNAw2wd74dF80rrysmuWGm06kHXfxJB/FoyYTL7dfF+lHd0tNuwDa1mNai8E
RUEPGyMXzT8JjCeroznjOZ0rXXAwZUuaH5X9kT23ZdgU3QCW6TpnCSsL5Ki5Maxd
wNkIZ8PCTqNj4GQf30Pb3bc4iV4RQSHNz/ipKWze5Dp35qB97HkORUiSinc4/roV
1QpofFA7XnAb/+owwOd8jw7QNg47pJ9yBYmnJZLMhglWJasKI2FLUexBQXbJ/mem
ihC4HAckezYgB5lz75dcIeaXeMUpByl4sxKdC/Zoz/xK8wang2O/L+TqLilGIlJT
e++DuXb6GZF7fI3opxdFPoRJTef1anfl2hXerNvrEQBfbAN1GEEc9FsbU6aWGYuQ
EeTpaPOdjShNVCBXneTJMb4oC/2HhGMKLRnNlDRSsZXXF60atXE73Ajmwkqn/ELF
ezYeOna6nYayxsrCm+oNfSPdR5mE67Q8oFFQ5eJmbU71rCtycbzSrJCYf5NLZszc
pVtmm4NmjZ0tO67lCyYOhES2PpsFeRPEwSEPoRGB9RVUhwzM3gLle3lm9lzny6Aa
s7aoEug8CsbaX6y1+gN+N3HLD6AjUFb/rV4+xvidku6Pm1og6iOqi6hObLsrv33S
JYFnZv7NdOGI/fHeK1wAaC/XNFiF30U5hPJP+cdF3e77KimOuA+mU6h14/95Uhzh
YF/bAaZY0n3a3fb09jILaG+jSLGL0DEky8KH9cQI25aw3usx+FXUzJKcZjSA1Ta9
yUC1V4G0GhbatQv8hD1fCkkLORCGrRYe4i2ITY6kYiL/n+eS1qjaiOSn1qyvjYMC
2gvEtj+WvnrUYCT04vLarepBgdl42X34As4/GolIyoeag0VKjNU3Orqd+vXrMXDv
nUS0qXXcWgLOcSQIr6e7Q8qByYaMrJkesv46f236g61jtJQH+YF/1tNobxIb4jkX
AwCJJ15XlXCtL4qecCRdyTdAfCJ9FYqoY35jbGkU05bOyg99P8YwhCt2LYYBM/r7
+GJ7P8pMsquVXfOX0XgT5X6nPSYyUJhbAzK3Uff5LdL32ehu2eWuDQG9SofkADVx
qAe8+zklODUQJS0i4vNE/ID7P+ppyrPLWgev5y/8heAx9dgx2d8xnf3j7EpCuH5l
JpIbeoL9jyHNsRx5HS1A5LSkRia/zCOX4Nhkytqr+8gMms93loU2JbAkgxSd2J5M
AT36EkJW/LNvCb/CVAefQfJqaHI6qZ9C6l5a7UDjng0khOrbY3fiov4RiPyDE3Tn
ARJNSKa5jMVCO+rSt0wNi5rrkxtDrnVRNwlvRG3hKPY9dpoVQwDDmEeV97d23QB9
ljrVuLALvy7YwHii49mlL5bgXxoEx0y4VxE+MTM3KY9Iz95pQxwG6s0FWctujHXp
WoJ1LGTpqw2Eq/DlXWTUe3GtCJzJaPfYBtk9TiE8n85CE/pV2f3PV8YfSPwPLh2X
RqrgcDAjTsTEC9PuKfhZZ9++iV/vVaXFlDwaALG4WZWuMeDMICcObZ0dPff0vOkM
wws5FSatohMLpsd2YvXQU5lYgUxdVUirAY3W1AZWEBJYwpZtt3e3SO9ITHYStDLA
6F+HHOHGVIPAMwZWtJtEgmXox8iNsgHBU2Cpdk6Tds7y1U4ZsjcEmaksJ1bHX32F
Bmez94LP5DXck7t3dpY0rE0H8sR1nfKpdFCqc0ymyS3Bn42xhcb68WJXIMVMBAyG
nh3261+bACXNGF1UIhhf6aJLzF/oAXMNhZ35pgewGjWfKT+vpq9BVqUHppcC5Vnw
2SnbZOVNT0EWJIWwVr1I4BBUnUp91USwwACdXu977mpwHjY7UwePiL0kZpfBGO8t
yWE0w7nxokz0/Mzuy9u99PWp64ZIndKjnu/8fxa7mSddR+87aT3BILbHq0yI8y3o
Y6STpm9R4eHgQi9hhZCWG96TnPtxfnHDT0VulL+64kM4O//+6Ohf/DRuwNExp5Ux
DmP26E1olFbCWMplXfDYQZOk5r44YbGyugERS6x6jxpDTNIgvovsWrMA+dMUKXRK
Nt25Ae/SDTgsbEK63/TmkDrom+oIywIPYlrndX3zjiWdlSyNwbTKisyAi1iqeOJQ
iUMQPP2Lif5he47JF8G8vy5Vn4pk5PnYSATUdubENiM89cMXKaMgy/7MMm75ouWk
i1rjGVHQh1vSGme3JQWqmECnAfRrsHsddtjyy5p2EP75XZYTD5PEfXtjfHKciTJQ
6xQac6ne9GRXHKm/HsXCv0bA131X5zaEi2tUjctjeNmdAbkoihF3s+8NDfcCdYSx
962lwFgFjBNWkl5EawRkh8RUK9WjHj3UxMCgVbtWnyQEGaN6fCoQXp77RJmi/IjZ
0LgguHl+JlLW+0S1GjdJIxuOTVlUZT8vpAmJDUVaMRRShz0NeIvn1bfXsJsL3Kg4
Kx+fgcgzdlJe/rM/c52B4n6U5KT2G9MWVyoKQ8jzkHEgiEP+vh1i0NtaMu6NBxnX
osKxwQjwJ9YP+bJK7+gNuCSDGk7Nv/QQarLQ9mvb0I29VPK/Ms3G4PU6iJ24KTgW
d8a6UcvpoIZVae+SiGW/ze6typoFHCLZMctAbDmmBCtiKA0R3Z02yaiRHCa4ZtKF
XnhseupigrVZB8/jP9YeIQXYelzUzq/kAb5JDz2Vh2D2n22qB9wqy1nZfcYBQYtv
8cKpBG9GGZezIovzTep8YFt0qStOUEKslNsUWOZzzQW81m3dw+tYU/lkpIAxfpxl
9Kt4FZwmPLNW5CJ2aH7TZ46uvhkbsyS3qN9rr7Ctk2EJ2yQpZ53ucXxwOlkTCute
zw1uDDksojK40YZmrmsuv+c5czTah916bx01CBpaw3SkYXK9oaWzE5yVY6dd9zCY
gwKUWrV5l3YOq4HfjBgdxpHyqKNxocUjU8+A7zFk79KnZnKVI2VoBcEHpcSCi9Ff
fBPm5koq6QEX1jFHBHzQycU5MRFBrJ9tJFFL88U0dpdnK1gvgvSBB3DiWu50PeCw
OGNc4JwDWAJiGMlwlMRP4tdSPysc3Ktz4SOw9z5TMEDW8WRmH57rNEFcZwVOQXKX
RcVGxtwabqs9wJm35VZcbQKkfCde2CFYiL7GZQKSqe12G9wV2D/q14Xs8+/kO0Cb
PLblb4Cp+eDXHeXs4m0UBaHpR8Z3MU3Zq7CnEDrY9RX2AmeiA8P8ls0cSuzAvNkf
7drhkEt051zAXQ6SWWbZRUU4vnCSHCvqNwYSd+jCNg6FWwFA3dnEmXvAimQGV7ZX
tFx7ydmzVIBupqZop0IxqYQFXqj1Ks5bMveW9NRj6XzvCmwHCjDOEH+d1uApUiZM
pQ+mi6pWigNcuWl1kguZte8Oc2S0C5YzNj/McB0Mx52F5PuT9/zAK6SkMmCaJ/jf
kDCDy3qlZ6Uk+S6Bxoqm9bVcMnkXO8ay0T0rxmUWlMtW/TN6mj49WKP/0BJW319q
mFPTmZylpfQ8R63D2/QcylkX0E5oFWIX/fqbvXdJ+am/g9jU9ttdDb/Nk47JdRoZ
iAouir6DGsw6sG9XZKheR/UKMei6uope+74hPpfGDGlJQIqzr/nEml/w1gRdIfNA
gL7OcUiQD2nCFuNjxeeVJA9arJ2pU+0lXgxbTZT7mcFNTHH2R48gkDSs0T8ORPT8
zsXKjvLrJX39oKzCSh9rfm23GmpvhP6yJNOLpJVy53JDoDskFtN4QOnN7GJaF++B
P5K+SRBGZuuWxZy3ED+kvUOfOktMmPa+nEuafZP/4erZA59kRjJwVl7nQ69LJiG0
PJZOJu0K4xJqUJQqKQ/+LN7TsQUjMq8za5jV8iUES/5Cuortz8rxj6q8EvqAL0JM
s6qP8Id6PB6K615P/etcJG27NMk72MCJwf11YwfbcEAOdkMyVksaQ/4TEodgKeUM
bLiFxJJ4bOnptGJpstN+VjfPc/NgfZvPBPTDxrzY3jYRfvhGc6NJ1f0DmgGN7xwg
0/IOhgpFB/SZTfehQkFwHajLzDNCHxOFPLmKwH61tjOH9p87+ozJ+/sL+o92tSR7
J6v/AR/x/zCv4h2Cn7nbgeS2boTkQT/+WBFjvIPk9JRtqowzB1uOeS83QywWBJBh
4gEC3tQcld7ciHkAzjhIoKwCN7ReQbnYaQyvmtpOYFlv0uPupdX7XRZabxa2hzD4
hgvq38CV1vVM3q4hO3oD7bwk2/kk+25xlUFtnieSBy1bnrQy3eaV9lTbawGSQZVQ
LljjGSuVUNAOeEWEJwhu0f5VozNZ+pf5QaVoZnGlsh94600avIBAwAXWsXlSpINZ
IXRvXr/NqrXBqLhlmO5R9aUHXyof0Fo+VoADRBxBi59C7z5gavg7vaum6C4Qk2Tt
AIZLVlOa/AwvHq5xmnfDnVh1qWBrUQX7iBCsTkfLT2aYLfoxZ68f3wlJWwsmXX7S
id5f/DndIrTBgV3k0NNQCCZkhwJjRkdgNvym/sgho4sTBPS1OA2o2zbgmtC9qvsn
VZi8pBCm4bhsy066roJkRvIV9VuvwcikGnejo7sCgddNSlQtgM4B5oM3k4VjGUXV
NTzNOIBEkYQdEh3eiWgSzy/uMInL+DTJvWEIeMuISmIwIMSLb+rdS8u6d7tcU6x1
1CeRcOKzJEZ7FYun8aZ7gpA9d06jJEWdtn3MRs4IQsPx5CRT8At11ymmyVYoU9cj
FxiztfjfEqBry1pK18iJHmKsYaFK3exF6GjsR+PKTIuDvERF0qvALxyFkEEagVpM
S6S84aNVwFqQ8VNE4bEz26Mw3u1RISoNp61oOIZQRlqluT4uvp1JCl9rx5Yg+oDm
oDq0TVBqR+mjspdfJW/4vC3AK+U+QStHUGi6h0hI8AOfmI+Q3s08fDZIJac8UfkF
dPcbLggqQY8NPRoOR/nl6wN1AKTP3exkMku8JfkfkWWD906GhjoeOeGSnh/X/Su7
yhkaSEWy4D2sfkf6Zpoi13HRBnwayaBb3aqC8ZfMtBFWYKYRFCQ7g+LUG0rKjCk7
vno79/gy1CRsC/42jcacZzWGZ0D6OmICxzkx3lUsJeg0M7gwdFjI20q+Se0h3bIZ
/0HE+BvCgO3gEGf+VA5igoIcOIRQcxK73B+0mnOvlVvg100iCzIlVQ98Wn4vg5AM
P1jIbKvMDvggC4NvrolBUr9HU4lkgAhOBFEsYOGCb6COhCTQfWo1BbtNQvBnIv4G
IA21RmTmqt/GL1reCQPD54pndBfhZzgg33qEThc5t1qrWfXy51AshX6z2v71V3SQ
ZKey2heR5C8yPNxQZKHW4DodRn/5tJNj9kuENkXZ4o+gXeAXURlDFM8S1GUuQtdn
+GI1NOpiBRTDK8O5dbPfq/kwBSikH88XHYgYPFkLGdFAYFagIPFw0Hp7RujjV3TL
aeye8FTxaMhn345EcX+vEi+c85iPZa73DDR/UxSPooLI1/noL5z2bpPXL8rYKcQV
TmpjqTT3Tt/1lSOAusiZ15UI5tjEjiTjZ4ErbSeFJa5BtdXy6pqcHCrPhBHxWyDP
/Fsx9WRqHtAhDP0FsfMY2vp6SY8dsblKMGfaL4qGT9RhczUlGCYDCYdgb5fX7ocB
v4bHlY+0BUDfcz+WiC1bKElhmAN/Z0oNLbjUYfbkJfARIj0eLOYEvtOFS0GzZpLe
ji2+pgnQ4IS65elaK4nwz6Wh6zsvZ8IU+WWsQ4wRnrAzZ9dUcBeBSl8JApgw+rzn
w8LS+dCmlW9ztlKWkoEQxLk/cz4XKL3RZR7EgSaNFwUOW4ZZdA9i24Qn/HuJIzoJ
aqep4dQSiueETqUNwFqdcP9+CPAF4ve4S/s4Ty/E/tM5DxaWTTDLhDhCXryKbzf2
25D1acQ0Gld7Ho8AA26Gi6exxlKQH+h+msRifQVlakrj5L8eAQxB/77IUD0Eei+W
+j2NpXfIUAd671upRv4MPxOcT8Gq1CmTrzhO8BwCkxtftdAp0TYUWore4K6S5CLc
xx0eZZ8haxxZyEoaZqzEKhgCIK+ue6gXmaBfLyER6Ked6fa0TEL7UbbZt9KFWbu2
fRxCMrIlwZgEa6Q7u2/CpIASMWJ/vYlnpqWJCj76aTy5tgcEX/IvYpqw7Oq/QMeB
1zdf1Fr2nRGS3j4yAlE2Si+zUqJ9Pahx32cKi5OxCy63Tl4AhCA+0e1MKuvqPkjV
yZl2skIDuRXAfauhAR6X3KOuXWHC862d22yla8MkZcUlWbY/DobmF8pkbrQsKSJd
wO9WUXIKtM9i8kefCLHDxps8/NQqnbsLgpZAqHSsW1E3dzTyD8uNBFgHoLAStOgU
FD6+z+bbpm38BRUxIFCGBNCv1evbK35JX0vkQUkTtg1Aq85dx1dVSMj6biKXKFba
Bq3rpsBa42R03yEsPLgnqzZIubxgg1yxeyyA4xk9D5FXoLavreHCeo+6uQBt818U
6iypuLnCF3qHRribU7p+tzEgCF8+OeUqFcl+iAp3YWOfQ13vSQnG4x4y1nZ0/kPf
By4PlEaN0ysRzrozi4H8OOn4ZhBqfo68r/OylzkEMIHU1rWZaN3e+anXHrJ0h2vg
gJdKT5v7NIb7DZjh6cKQV/4SlWUnNTa09v6qcsPWtrAjDfIl8MuB7NFGUZSs4EHn
bZeBzItMAuya3t702nUSvtKwmb9h9aPZvinY6iX/RQ5hP0z4icvqNoJfmHcMdJJh
N/2K6J/Gy2YXt3Y/vOX+eSK4aneGbnmilkr1jaxy/rIDykyQhE9WtQAX9yaC6FU/
3BuSmSGYc4yLnuwWWPGVpYgG6PkUpZqf9CQgb+pNBMRBAJ06E8Jmf4GZil67niDV
rryyVZqwOLX6zV8aVdnJwCSPaoRDFHRYgHr3xGYtZdYcCn0QOUGoj1Pv/Tj4P8d6
E0x7Y30q9uZs81hlnhjH8dqT5ZTp5F32MkChEA9y6UpBKB8ayPADczpgMj2Fde8d
3p32rULOU9A1Q4OPmwtAoBENBjk76kjvJGenRWhb+RM+p21HAE77WBMm+WOcQnm7
YS6xufnUe91U4cO4bnUVUGrJ8YsOzDYPA25nM1yPvEldFVRXByzFgT8gdMUsjTNN
TqJhruT8wX83+5LwCct/j4DL1bLpd9S+XdorVEeWgRBoBobq+Gt3nvlJrTZN5elD
ADXhlXxEfsvNsvg0tqsvYqETI0i0C+rA/vWUC9Lg4Zbh3Ccvqt6E7jz1hozVPLvs
E4C6ygkzNRRNtueEYD/Xin35u3UOwhrDkMbX80YT792vHXjhel0Si8oy1R2lnqLe
P2MUorWkmMHIYs68naFF30zKUzKQ/h7+DyyZxEM7XfmM8xE1XL4HAYD2hlIQ9Vp2
AmKTw8hcDL7JsJvHjRuxnPcBhEKlpmnc/rRoWZGoZJ6bQhFrewyef9zPQGPpVzJA
+DlhNx8vUzMhLu63ABf8QsHukeuGTNexGLdRqgHJQSlf9WkLOEb42C8zbk6PiF3j
lZsV0CS9NR+CavdM9K5T2ojXhNQ/MoyBnEzx2ZRJcQqqs0wM2AaXAO5Wd6gKlnt3
TvwVsM74XKxsMcfOM4soZWl/U2taIQdUHgudazXP4ijyXYShmmkUMBExkVzJeB66
Zl6kGRp94vKOQKdV7atMEkQcWl8XhBg5Ab/AIfzGtJwgWHdXxHnO7Vq0/bjUrpSK
ud+m8oeV6RHPI5xMCEsyYYhZDB+h9v4y4ekELW+mBjG4qL8708j4Jbqh75PrHmda
Jw78mF6yVv6ZNNdcQ7RBr4cuZcsrVsoDe5cnv0y/xrIw1EuFNVEayyRO6O9KaypE
isQUwk7AcPe/9Cc7jc3MvfxymVW25iFba29WeAG2vMa8Xy/N96z4M9T8SWrlV7Zi
j6VB0knW53i9TPEw2I5pwjD9UNnx57suBEs+Cb2SOq0GVO2bpVtdvDJBkImDQCv1
37rZuYn2v9yDFT1rT6+wlQfDY3unslyOCSYrD5b0k7RiH6+qindNgo8EAr+5ijmB
/O9LUoWPxo5WusQyFCnlZ0KeJlHI8CTmuq0kFmDHwAbSYQrRaLQNXGhWtKESAa77
Rhpu479Klf004pbym4/zaFZXyTVwL/Y8fOjD+Uvc2XUIGLqWTqOfheUuo5GDqlEl
4CLGKtTi2wafPmN9zdtl73A35YhVQeEg5VAgP/I291kq4BMSkfxSAJGGHvL/g7Ay
4WA3rIvmVck8NV34z/rFy/D2WmDGCYp8u1jmrFjgAg6VK/DmmEs0IiKGhekeoXAN
ghzdqB/wUTRLozfiRpHabs/+B/e7zPzeFOfxbNoMsQf9o+HZ+GNbX2Sy717eS8Yh
Fd7ty9JJrbmwH1jaVEKzdmFRMW2L6r8n/TAxoQfspbmix5qxHd2o2/50HeI7YXFu
69SgG4fwyfEa7JrVVJyClKYg45fH4mJacqvs1JstWv5cOwM2ZlVU1+XfiE1qNzh5
E/17Xn5LcCdo902XVpVRCpWrGU1BrKx9ICdF8EdhmDa811u2UY9eROI0Ksatkr0J
F7S4WDXMJhjVkUd3IJxmvQiJB0OSKZdK4C7QzgHC3fwkPgKfZJS2eSrFCTWcOM3X
s28H94Yarr6rGw4NWgFtztjJlGU/voFhravx7LFV1vXhLBmYftioJGNxR2bX32yr
fRG7xu6dbx6oyjhik+vSE2lrDhgZJbYFXf3CZSADpUSt5mliGZAN6ir81eYyThUk
J6GsClhgmO+KQ61GLq0d32B6E8EznrQm9aRRZCKJjrcmuyrIB60JeeXWJw0YZggZ
45uk37FKY1NEI86dfRULpg6u1ZYNJY2fl63y2CNfFcg2+iQDD9K8JuaSmqywpAOy
Re1e+etl9SDnrc+KP7pOnWtC4poW4Ix0qiy1RupLMoiOEgM80ZY4b+hCydaXvt/R
9CE0hx4q14IMaLnq//weolpzq0CIf5Io5pscfsrdukveSpM8iI4zhLs73hDEALx8
NwvsH6A2TibM05v7QnjtUh4DvqYwOVBr91PJk1Yev0WWO/387OBH4SfKQ5GdKt+q
6q3GPq6MzesssfSXWkUXjTLJVTjS1wgGv4ZtfBxW1fAgjvec/8saugw9uFYTCN+U
Qu4OyU2czDUpSwX3b3WXDf/3xN5JYAZaPcXaasy60K7eT2QXvoyFxhwdkHZrt1Ao
+Ne7PCs+Kb+UxcdppQKu2IVThiJTNbUg6qYuEdw9jds2a38toaa6P3LxQl9guPB2
0BJfYNONMDrwmpDX3GWTTZP7za2qN2X1OsKyMsEf+uswwilA5vSIxPoyiqiU+BXf
jl0srvWDPvZfEjPyA5lhEDBVdNSdypFBBRqN27uNnBSj8hOBJsLG5AA5C/kNk5fg
GOpiWc2Xf4Oe6qkssYnuv5G6+BDZjQpmpU4nOxvNZVQSIqzi+BAJBV2tFQtOKZt8
2pWl0eFFFZkif+NyEN3CIHCNsyi8ymRtt1HoUgTgCEieC+Vw3kZc6aU61+eCTu+P
169T9ot95X8dq0I7oKiWNpLo/W3ssAEItJgYrhM4qnRhD/ANSGbLxaC1As1iDAWy
Sa0NOXenNsi/18CUWoqO4uxQF16B5vN4FKN01Cv8osrk5KrUvZRPyiHtj0YCfxj8
kMNnnBQ7pH8/4Br48o2xMR0IBT0/SRRHBDfwjciS4elobp88eBqoF6DTlRmpax+f
1wBaPrNNpnGY6TM5Zf4egOH0/V6wOtHKhrwvNJL/fX1/FMaJq9gNikoYbAtSRyb/
/TSgzgrmJY63VSi310rPHxGZr1QQL2QjYKpr/yOWcETbLMOyJXTlE3UfGHnxKD4R
DwQ9C+4p36p+VLYsy8pg1qvgrV9QgcBCBns/U+/vAZihyPWJtdB61GEULZ8yk4+6
rCxhDvUtNAgfxHZRcE2WhXiq7khtKpvjuq8FtFQ1KV2mFcoWWpM/xl7DV/DmsOL0
0BgZDCShTnBYvx1r7h/Wdr6vB1y0gMFJFydR425MldPCJklkCNyV29pq+PlYu3oH
PAU0TTXOZGOma7nEyQnDbC3hfL6jVkHlclhbV8KFR/dK1givlReZ2Elc8tHbeURN
oxvjmJ6vBaDrc3055TakW8lTog1VXhnwI441QIqwAttDlSwtIBrCw9bh9selCgTH
q8mlMilaNqO4N+bENu9F19O2WCRKVpDt23ehaxT+9HNSFHVP9DsEKmxoOJzsz52B
Em9h38hnOKG419SgCbYOjP4KS9V5Iu68ctQcQ1YOKHi9HXNoEdUKLibj4RL1kdoy
8vloURgCTw5bymCfHWK1maw7ddM84AqyKzF/J9m07MkNAnbgQoWKpkg8qVVWxLLv
RDjGd/abBtLv0iwhRLpw9tpXU2ORwelOaOD49gJRMuuWkN8k5GWPkHK3a1zrGgSR
TV2hHSTSQh7M+VtXcNlpOorIpQqFimFYDjGqmfedUyYQE3RuDZgx9Wi0hiZqdwos
nVQXVFVVRLsRhEjkzz0acxw32PVV8X31+k+Z74pzeFxxC73s3bnJ2lhM+w0TgqZ5
3I56gOH45991jyjHXaOUGe4f4ZEXa//29iOVFRxsA5XRJtuhauiuvyjI7qn3VC3X
1v6YbcwYVMfAGjhPzD6G4Cf2WdGlOkmR2WUXcdDJdtsIDKbFx5lS+kC9zGdQnzgV
D74ZmWsmXW3CMxpc+QDV5jOmVwJZ822ljEHUnUycnPML99inOQ6iZ3J3HKtcrtPZ
zR6+QZQqOdN2ApaYLUEiKpHRwBorIEJrqsVeKvgcMet8AFmXQdnOiQdZ//Ph/j+B
7pW5Di0+h5wXzvKzZKywUJSXB1So7RyH/lWDL0ZI/OFbka234e6hpsIMvlKNysLO
wP+nMSKMMPkF87pS8BV+pOtRRoXsK+FaA5zkx69zA/QZ6gekEs7sbZFAAuidAway
uRefmlTValOspKH/7Yq/o7zt9VzuUlJ4lrLwXa4465PaWoaKchSQ7cKaGpVXxb37
uzvEaWrWEj4hPVZEuE7lSB35v+EAi4EWp99yQipx+xmQur5GyP+jTL/AtFsMmKmA
JPC640LXmGRjf8+VUc2YN1NYfdURWFYYBFABpwMcnO8+Vt4/i3KRM8W7GpwK6Jq4
1Z0fv4fVQKF/yC6ml55/5ZXhi/x6JZ4WxI4cVzCET7I1PSn5NO3eEQVOU71hh0C7
lMiNhOcPqBKjyWkGKT/TypdPegQ2u4Tig5Tay9oksGiFSCtfX2bfScP1nDBFhjj9
+iTGZgwTWHyXywHUgwiUoPRDHojtPGj/F4ixabCtLNKFmAc1it2Rv11ZHkSpqQEK
h93s2s3oGTCwKlQfx0EDqSrMf80HsXTI3uoJa/G4MUjV0QWiv4wrFySehrUuaOrq
Q1Q9rCALFNkLoQlAi8zeTYqg74/2KOkMDgcF66V7d023cfuhBjWppKR/R6MRXRJc
nWDYUXbQEo3B47cugcuOG7wWoDzm/DiQAnDfczBOj6gGiLycCaIlnf6NWK3mBOJg
yN/j6FwGqKvKuIxi+L5pzUUuiqq06qnvyrbLmsM7rPH2udbmWAUe2EvTUN8M23Ue
C3uXdcEYndfN+uyanfXkqqZJ/Tb03GHog+09hTM+WqkrIxNMXM4Jm2jGsyusUYWU
/1xD1qKBiq7andL89Q9s3c5NZNQ/1DMhs97yYYtavDX0BPDKb2ZOXderHVlNLJb/
iDHHmpn/NnbN4tlX5Fd3UNk1ulLI0RDuKByHdntN6adXvI59atI01neuwIy42R4D
HuVMSIiPkUFRTt8XYxzTM43lCNhmyOJxLZGe+iCEXOZW+JYpY0HGmyuVXU/FlS5W
OWsN5v3BrTiTXJW4btfpahn2FxBBkQ+dzEjRY5faWWzEsyoFipzY183ssT/HnR+7
4hZoL4T6qYlUDG8/6fzepb9JnWPI41tOwDimAvvH0LrpoU9Gupuvz2xAO9LTI6V3
Qn8Bb4uukvW3ZlsrrBqOuQqSTmilC02vNzDvURJAS/sYoTjUrHDx7Jh3SAkjAbjA
XiPNkRC+PWjalfguj3WtOnuClwPhzzGqU6srYCT2wZQ/JCKpMm2u97E4rM+ma5q3
pgNLzgymjoWswSCbyD/Go3KayQQ+9xMDuQbnhKkmw42GHieLEOGsp41aZ8qZujof
KpiVVkgyw78cwItfS0C5mg86bdGJI//8rXBBiTL02PUAjfTFi4PsnoWZQ2LSHhAQ
rXjqO+hdnpARpn9Ih4dsgZj26AFMYqszip139KZpCJ2ib+3Vie9ZddzmJkalUPlf
5FcR9DfZDnQqw+C+RjW5iWUHm4lY1QYE4M+/mvxkTOODva4YFJqqABC8Hn+S194I
pNtxxTGgIprjAVrLM6+YHYhcuIr5Y16E7lGszGDi9P9pbdws4+RkyjsP81vRiVCX
bROe9lvlf/DbBfFTk4tx2KZSrdJ2gmZCUcwU8TNs8viIO4+zflVyYd9oOuy5+tjM
RrRnXzDDYhSr94P4P2oONtlxvCapfaeZBReYKP+RwOQZWUrFlHtzu3mu6JVOpM3D
N1hKmLBiP1itu8zegB93flATwmixYon0/jwbFPtdULiT9QDZdDddj4VOgNGReZwd
4uFQQraVcUalp9i852S9MKQ5Xa4qWZLtPTpPnEnmX7Heq6qIrPiTkcD7brLdK1Ta
6vo31kDcQQsUskYiHWP9jP/Jca2zKUFYuG/vTAH5wgpXSRErdM9WRiIDSboaJd2Q
HKmyaZKON1pwjXuUG13wuxAxaysEfiqNO3iX6H5CSLzkto0jg1YfSXHrQC2jyOW7
2NnSk+xTAQAN932xj8eLVg2Kt/bUjS7PtIe6Uww7/Zr2z6pJf6aSxDHEp5xeoS8E
3KUJXn1BGGtwkG23Z6t5vWaRerlH25YlhPfQNPKXStjGO1g6rxTryF6T3YP2YbOP
ATqqTpq0aoCrQ1wV3D1Jhzq1UnWH2z6Avqqr1jXRzvJ1RGS4aHfyZ0si9h1CpI+k
XZgA/T/BGqDgIDxpRkKMNFrgoUUR3MzNy3b9ehDTIuYapEe8AE3Mg/tccBKZSLf5
Gv+m1FxbjWV7uix6lI4zKnfh03kCsb18KRsQa7Ps93C//zNWq5Fui31zJPwMSfc+
mHt5IYByQQwR1mRas3SonuHm5/Uupr9uDTN5whV40t2PXr9Ja/u4YFTttCqw9QPl
O6jf7nA/7CWktZ74yKj7a03HL2hVrjxVJmjZJVgUHZlYj3AQljbIo3PUuym5uGXB
yzbI05mdnkzFeZtQ9DWRGj8Ep2j4+Y880vuruLE93z+D63ARvKSE/n2ETC7uZjUv
Q2tlaqpxLqUFYIv4YY6+tZRevVoUKMnDvUSWfPs3sOGXnGpbMw89n+jlk7k2Eq+f
HaaU/mlBvL2J0ymKWehoMwrI+oGNLNI7l6QKqxtZ0tqtgM9tMH2mN6PF/rtug8l+
yfeIOKA3UXULPi//b66V3UtUqpeOb9QB0qtgnjD6ukIm1RcvAp8JiKdIP7Zz4rwD
daeVlMz8njbYB6x2Wqf7q/IbopwoZI0Lfo9+I171tx5TiHPNfo6x1bST3WCIIrT4
KGqq2VcKK49WFKnSVzeKEgXrWlJ6H5U+FbIr6hc82w0cCaCx0VxHR0HnrE8z7s6E
UR5PDKmeQEefZ9yyYm9FGgapRaJ3e6cACmNowBcTdfdUAI3NTgd35dh2wp9j83lB
EmGW3gFv+Ol1W9x9TNl2GOEP/I1uN+qEvef7/F0MLBTslUHYLDIb1cD22IZAGnkO
OPp5Gt/h6Ypci8fND+qxO8AM9dY+TnQpIpWZ5qZSW8S4leVYyPu7/aLbOfKkfcZy
LHfJQfHfHWM6lRIMoIJyWBFD4D0968GcWsJ38p0XzKuats1jLwm4nD9OUWaNQHbB
rneX9O3VIDrFFHUgkQiyw3eJQak7MA6+VGUWSmKuRWKxkSEU6gGA9o9AfSF4CqmA
UXSRJVb/0wktLZg0WdIeseD3xtjjsXSdrjt9FvulP5CmfuMxUKOwaXLDpqsgQAaM
xNU3bzSEQT/hfi8ytz+AiAZyDNi9y8QxE22fXeSXr1U2TMLQ5ds21zfdPOCTTT4n
sZhOBsN4TGGl49mOhXb64xb0AJ9RP1am6OUfV/TFKKJGGpe/ikjmcu4dPRROkyfE
s1JGDSdfD/G2nxZjGn63fjCqVkf6gGeRSjgYxGPdCPPQKKoO0Sjng9wIca5aj8Bb
kKXrZ8xLVCKh+vvhAjsx3d7rM26+b4CQlTAljoGGbtBiBSuDZvVfr23k6SRUkp8z
V/WI6I43MKLc/9isl8/lGHhaXXIkoc51MX6Yl7b4PUiLRTBoWlxvULhOIXbrAcLB
0OOHayDITp4QeFCOj/iKeighIfuApoCthc7OoP4m2VJbuw8edH3zHdmK5btRVNGV
7V3UuqY8/+ZNOGpUk9KwPvygVLMXK0XWx6proqdJel+qaiZ+pr4Uhctig9Knc62h
vewR/irUWa+Zu6370X4LeNUe+tUXLtDDYdGTkQ1vZ1TKJ6BlaZn08c2yOr2k+DUA
6N3w25i+lvmTcUmJr4JGN6I/xuQAP1YG5FO+Norgi6EO41Wi/9S4mN5DlSMFMkDS
iELtWgvL/V9OP20CITe3UqQpB3OkDhl/XEDdIneL4rVua5sW+T4+gNGcdGXRZpJw
1cwb5y0P7DmQU5N39Me0O8h9r79V1Rxo/1RFCHu/YhDpZ+J2MZmkv/fcRGb3JbaY
BVwhiILLOBJfn/HrKZQT8fPeoypaDVg3Oz/Jd1e09MbYMLL+Gr43kL3FQIMGeCNj
E3xtjUN6PmiVOSmULlA9oT586ZyABkqpf2gbSdMX08p9BBZxcfTS8TQ8lqdJ3klZ
l9AkDEfuaRH7EZcbYc1OEgNP3urQ81xuezGvABiILOKr06XHbInQvrUcuz/Z4+zc
7L0zbO21I2cNNQwfn/q1jDhELowjuBPOtjKUjTBjVYmUQRld99gaTL2prvmYT8Sy
ulVIsggmbZn/i7Xb2M5YM16jgLBRWZ9o+sR264YD6mzkg4M5pu3EjbPL1V61JbWD
6hWOsU7EhxZvtxVmspc84xitowTOLzsDYcrmqROhtUHWwLyBSIN6Eglq6gxdVFZ/
lBkBxmKeJKB1nUBhTWhHClOi8NK6Tx5i5LurN3qaQu5JD2sQcvZ5Cf4rk0z8GUEG
oydfkL3JdZaA+I+vH5LpjdLtnjx2BxvehrogAtGVok442d8XuYNWPdSlqkTV0D+R
btyjT20ivzKPhblIattTjcDB7Bf6zeQoweyhMUeh6NS7vHRd26zO5BSesGQNCIBl
7i4OCdXXryeq5OEC+zh27O1allx1wwPjDkYOy8LWpLlo8D67jqx2aN+fvp+4G+ln
C3dSAhH1kxx1H3pvMOxu0qq8cwlOhi+Pv+uWMb4IfY/PScjdNVRKhnSeWPEaBiWJ
/L3IYge5ITg+2hHjUEj45PsC4nnk1r13pXBDJwRoW/3j8/0ntnwufdvS23NxNVZ4
Xeac529iCo1OgmNECq6ZtDUZ1iGf1ITlCNZuN5s3uJhOguX7i2kvQLP0ne2Wgcju
mHtVGb80BDMrwl6I7p7uFqjgUq8aFReuu9o8V5+AucT0MB47u+Q4rZhl9H+9G26I
FTzUWba0MmILgZRmB6cWJyJi5/W/X+6kCYtxkn9qMWPlIi/GeAwj/jx5gndugpPk
86F6nOk14flDh6Toj40Z4Y+cSU4JuXeYn1JJeeOYUe0ZnDbQKdzJtyRVlESsqN4N
y8u/qQy5JVll5BmIPvQ7JnJt5qYXBWBiPvbe1iXOLq9+pqUeXWfftQYYX5qH8+y/
uazCJJaSclBZbQ7JoDAFi/VnxBh67XNNMdWcQhLH4jqlwaghpk8WpSTxSoh+nYBj
KoK7XunJQWE49Ncz9v9GzbgNdYbzzCggo+FpNzF1tsntiNonKL28cJeFGtowJiCb
6EgW1E9fIXWIDdXALVmf4khhoeViWtR7Xmn/OUQlUPf3WuugV2BHc0eGfFrqhrhP
cENjeYixqK3BK4kVqOp+5e7+PJj97HLbyUnebkbKplDomhcO6m4hkR6VWuoVIj8o
0qNo3QCz+a09KcbQLYoY3Gr+YF/uq2roNAfNYIBKM+u8rP0Te+AlGjPzUrQRsfSB
fGm+BbwpL1lh+4RVtQDFL41Y64zl2QHW5TB1xgrTB+UrZkj1GgTzSnFFzlRjuNKm
4+uR/ra23/113l6cPSntHyqKihVT9AkEuD2Vkdq5grfY5eEbxYpQGgud9jAUdoj9
FO1ywzv3YUWom6sRTcdI1mxir2wL0Sgy5/mkLnirMtCjhwMcbmOCBo5dF+Hu9LrL
MncoLi8WnumSlPTKlqvpkbtrf1rhhtyX166fRXPGOKeRxVcWQGvxFa6s9Vrzbw3b
yEi4P2MvwxejPsCcQJwZbDxGgWig45sFjW5mwCHKIi4dq8i7uQP1vYWF+epvW6db
D0dFl3e3+BsSuNUAmNG747hGfyi7n0TGY4sUP3cqICrh4IC36zq/k7V0mIwzgPjO
FMioR8ozUMLcF9iqkt5xkRO1B+fkIhynWYtfc8c7nnIYfLt5iEakbP0/YjdcjwnS
Dw+LH//zliu+ZhTmGZvCsUMlQzqkqBM0nDo3JQDP7FuRqeXdJE4L4yzjiZBToFJ2
ogd9cWqQHu/ad3utyTID2PnAoR8yQBlKgPpcXasiOTzlg7OuYCJHdnjL4faVjNx7
HpHLHxxo1p2CKYwEOXbWch4C73oqpg2yllBuxVFirRMeJp26WEGU8Rb5bXNvf3yD
tcC6P6/E/TUpEKatEp2MxpS1KoccxeiTzp7805iTnDcOUiKooNfbDZ157TFbD2BF
75Fe7idA33hhGHUmNOJBA0kEw8ZA2ZNMkS9Bka3ekXyh5YJP85jfQWFHoVNe9Rg3
bKciMDwUTJ7SdEuZM27aCMs+YIDVkdbFYPRxMGUiW7F/RppXBFW3pR4OorHZRcK0
LmPaGLUFNN9K81tU6bY7LiQcMYE0V8BQc6IT5f+r79zpijyxVvMW+JggQJ49fJct
oc/POolMUqrpbd3tSqAAIW75jScEObrV/R42MoSfspxSErZzqYuJCnjnZiPMf9B3
O045MppoG/VPBVh41UK+boo4JNcU7K2D8JG0uNNPSRYTg3/fM1O0sNqjv0pW9yhM
4c2s91GnyYrOqqzGNTm0L7p2tzfmoV5MnLrYwViR1qmyL0q5LHTdcAATea2r9//1
8/Yegu4UkbkYTB1u3ABbw3cEQl8i3YogkcW1H1Qs06g0IK8jcyMeEljQDr3EEh3i
E6HImobgQ6yNxt6zHYmQ4yiGcgoO1PlL3sdSynr1nklhV7nnsKkHopCbJ0IMHCnV
CjiLaCu39JfngBmfaj/73/oCKyLytrI6DMOQf3M2UaWkLD06TrK/9f9uVSrfefi3
t8pKFp/6YQ5mz9fXjRYjPhoc3AWzjEPZmrf186cGRQWcvoAAVliWD4a4q7LbSi1w
6AWgJjFhGy+LAcDQ5LABH0sH+TaiJZhOwwbqHpo8mOsvMR9ok01Mn8MiY2zA6Jpj
qYCNfz6cO8XhT0Bs+aX1ryramdSoP/BXCztNZqK84QLt9U77x9+V6MKGvxx/hxKs
DTciGD+XBo15HyP3xHU30Z5kwlUz9XyZNCcQGNQS0ncpfFfN34x1rgma45viKs0l
ZW5ksWf2zbEuUzPp3DoR2GSQGKko5LXww9t5ibX+O/9BhZIRO907LG3DdICZpIgy
+ZNhvFpOlhYIsgTtkTjYRjPjR+hdY2k5CRmvfB64lIoMuYRGI+L+1EYYieCmtdHb
ReH8S/a8I0pDtsLtnFegOj+daBUyDZFtP3x/NYVRH8NQrZ52MiZWNUCL8KeJ10Yb
vz7HIwkvDV1gTjgt6z/1jTgSzZM1JAWrRF22X8d9qBV85tkivFvEYXcX9fJdRxgt
DMh1bSY4qAlwCzMCtU9kZ/076nf0SmVo7Pfca9WMKoGLHn8FYhRbgibJfaV8lm+J
FjLmrqeTWkH/6KFtvbfpCoCu18d0x7G9i2wDLdUMr9RvHGQlJ5Cfn24FlT9RG60O
N/mZ1wmdSHhVQpA9IbPM9hJC6IYydM65/lAgO7sgCHGG7gwM1Z+tNwL83X4Iz65K
nUmfRR5cu8Vx11Lfk4adHHHoS5bCGfAkr4wPr1XGiJsENemw/4kR9Fvac7wvjPVY
cLH447qI7ss0bjSXnEwKKZz6KxsELV7qEzQ/iGXNZOFoByAXRXIyZBEyfbLzwRnd
ZawL10086nFwIa2SqFjWS0L6/KFh3KMnBpejXzzVDsr7FemvzerI5A7ZkgrGOdkD
F0k6C03dtYY7xfkXgwxjLd1xXYI7sO9cZhhnK20bW1dP4ITu2S6If7aQCvSiKCUu
tfVVu2ra4tuYsSMQI/dwbeaWsGSEbhZTWLx84cuOkm3e7uyDx5f+dQ41TiK1HDco
/Ah1W04I9Za9eKyhW/QLEVq1y/nwNbc6wtnWskue9AihTmiJ8Omhp/xXmybOrvoL
5H65yniaX67jGYIhLOGewkyJZLoAALczu6YlQh8a2dT/8QFiyxHQ5LbYk6h1Mgvc
DMYnE4+JOl9jFKcmgi7ONNn1r9IoOTf9yU8dSNrls5Np+mznwH0cF3zCyYvTNUnc
3zD3Ilr4PpIDGseE2PrQPOcjEe+rLMXBYLPfRLoq5uKAJAEPCjQF7MetPlRwW/IJ
7Wwi+3QXNn/W0wj5X8m1TX+gl/amM8HF1m0s+CmguBzjhgnlGA/8wraElNw9dV33
eDq6vyMnuF+qVUJSnzVg8Rf4TUHv2N69wuTk+Gf6Vwr6DctDFMZkVgkwPzRP9ppY
l4jGzC3fHqS6diOFDF3Oz9PO4Sff5QvVgolwZsl+2x1vgcT6dCtJKl27z8vsIDmL
7nm/ycwMO1fV1TBUbBuHvw==
`protect END_PROTECTED
