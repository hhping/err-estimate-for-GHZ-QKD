`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FeDSpAxPMzT5Un/hcJMnnpPud2fwTH0vjwMTbwIrxgXzvyZirwgNoLTaUmW+RVl3
t9yCT0VqIPFuSWw7ZXlyjF8JJ45VlxeHrXYDEJX6zaVdAMQ/1S8Ww5ReIBUaQ2M2
4Mrd/xkPTgEWnXtUCQ8kBEHoOAwUe915E9CmIpcGJR+eLtiYzb1rsuwG3F/VUgoi
BX+AaMw1Y4oBHLXPSiQj1rl7xZxB6d5MdVLUoOs/aUJaK4ptehhr9hd79n90e+1o
NZ6OA2Lq3ygkmszXpub4rutFjrqNTmYvO79vPqYHJ/XHF6Yu2IsKSyt22Dm3l0/N
oNF+zdwYQLwtUiATJ6Gx89D9+EYPzbzmNT8oq+k9enLbrjd6EigK/jXzLKCM/dZ8
6xhn0qpz+tUzzE8y20PHLIljcW3ii88gPeEKr3neWPQxrCSyrbCkZL3UswpmprLf
K72r6bvbccFyPMduRmKP7kjgq8JZApLm/JvNFrJC7Lf/bjHHgSAM2dZ8uQAMv/KI
H7FM2PmxwVfpvOIVdY2QsivraCjTiv76d/pjB/cneYppL4ZtU8F3KzPfZYyF9s5c
Idg8g7rdAzlG6jkbasGyoVKry2WHVwXMNhpgwzjd4xaMi0cML8x8UTQC9ispGwqW
GxNldneq/4Y6iKMrAFeF/SXGDcbbVEoqg69gql4H8msdKfeQMo6nuZ+vvrcbMlq1
oNFcy2HqgYKXjYFf2MsiyTaWcGhv2iTzWkyJzYd3G7JaXd83j5n0h/bFUYnWg4i/
w3Q4BtP9rf6xcCH2xsIfPGQmwVKac4C5xNUpt7o11kIBoYYPqbVuWwODY5M6w3Us
/gyKHpLNXgjjnf9X2TWXnpYyMLD/KSzd7rOsShETJjy7s43/+G6kjNk5LLv6RcV5
fd3ipb/5RgrRxC8H9vlWuou8QjGSOQcNJ/qP2liP8uCP6roTsVlhKme9DjyPOLkH
Px4dcmHRjHVn9R3L+SAEENZ1kBBuqVybXYcjm+5qo/z5qgX6UkdT85HwW1tSVhVI
2EUI+/F7DJmqBoup3I6DVwdEs/8QlICikUwf+NIyu6xVcDtfXWAmuyMix1CuYYbJ
/NLHoaf2MGXcvJb1fWtBIpkXSV5nkdXOoaNrKP8pibeHW3/+0aIk2Azgj15Hjdxe
SahTXRVih55BPC+UlGYhgoAMH9/NtTmDwogxPJMstqbqu6uozYkJ1la1Rf7gOgtb
ErCE7X6VQ3cMNjwl0bV6HQwKrZ4CKKPCNkjd5CWRIalRk1ttNQ4FhbrVDPY3PX8N
3datMAmEKCxsNmykun2/Alu/oww8AfT5SL7n2UU6hjyXuUol/FA+Wntod+bJUIVl
3B9m7hA4Krm9tjJIlrjrCHfxTXiqpqId0xUxlYN5KbeYh6iVNaUhXDAX3nqiiRKJ
Uqis/HwIgupfQ2n0iEmn3E1YBZCfh3YIYUI7J8so9n23k8g2tn/Qs94KYlP67mNK
kcVJ/XXBo/+n9PHikilIMMR7OHpq4LB9ED9YyKZWOg05b9yitNhgfi3mc899l0wW
itcHyNUhQuXScB8sIaUCDb/qyM5lp8EUDt90y4iFKH6oTEMN+L/UgbsVioz4792p
qhia6qTefaeBTihr1/N940xYFhLmpRa0kzv3k1Dlag8DLn4twMcyTMhursU3UVGu
YqskYXUHB7EXismJOJsgPyMOjCC00vntkDywY2XSJRyyQxJ7IIY40hHG5j0X67Fl
/BB3FTSu1rijcCDUOq5mEACSNLPx9UmW0t0JQ1fDxs4KXIFgvUbONaxUTuXrWHeg
ch288XQAzHakFFe1vHOJHMaxMwK/rpEUXed6WZJIZ2EHOnx+cRpq0/V5MkLd3kIw
PdvCbRk/QC+rVbtHIQJxOnjNg1GyJz7QPoZZ2F0HbHzqQlNAP+yRhdu8xnKrQzcV
6Jb0b8m52qbUkIudKhTc93FBibQ+PY7pk5n5O6s9J2EzRfX/KCzgVOAwrmvGI87K
69Z+cGP7P0DQXF+YLd13E1eKyM8eR76Ncp9Fv+UxdZ6yxvu8zbXyBUA5Llrtz+Yr
o0f1dKjtw3xJ2BCOaMondQ7cFEqG0MWNlV7HFr9tahwHua0ffYEf3ZrBs39/eTCD
pb1UEY2GgJZaquZRLj8ImaxWnjTqXHyb3InvJwY4FjkB3moSp9RuUYMRT+QTKsz9
1DhqnnGPD/ORX+3j9qb7DQWVfmBXZdy1rpNQwCyyOfHgkLjjSTtsPM4q5RIZLpym
DvZyI6v4KzJyGSs7w6qgp0Kk61nPZjqtNsENBH1P12OR5aqawwy2tk/xugSAgK9b
m79J4tpTCfnY62XSVZI5UO8tQkq3pqo3byWnMrlIyj2xxewylWoPh1xxQ2JPQa2H
tQUwSlBXaljGxykLnebYQ1ApQnwgzMSov0LUVWf7zihE8ogcigoFD1G8PtJh60lu
EwuPVIzSVFDL/IxhfsM2SeQTRdttJkLZWQBmJu2S1MxtIFA/4JwMfZk5+yvTmxwF
pDNJGIJRNkOsngGNVy0EA6JdEGzGn4DDbHQXS5Lj9zemiTP7V8GJdTKwyCUQZ1iT
dxv5lwziTnwPOQ/tXfmjZT7Z5poQEDdA4nLs7PmrnT86+z+B80MhZC8zD1NVNFhx
pwOalg+5bxfmp9Kc5WA92cMoszTufUoBWStUix+QaBfOSKv5LhabThc6yxx/GRny
G8C1vdGvKYVlaZ3/+evnMAPlj0Fc9s8zvYPtDB7ZMBzx8x7/6l+fd4JMWPM7d6Zl
qEfiPTLD3OkwovNyKnAJxXmcPwNdEKnJZ9kHAjLE5bsezfyFxfZ18G9GkBJmZcJU
yZq0MFWJzBGqwUMIGAFXA6FVo7aWacHL2KaHR07TCFb/DAa6Auw1a9sl9kBCGvKt
EmW2m0x7ILFd054qR1NE9EGzsVqiXNcyz80xg3LseLl3vy0CjgvSDW7rdfIZ4NI9
5mAE4LiXRIsXigm20AjnZ/6iQC8yCOf4iMfV2Ums1LuEScHVrfmS/e837LOhsjZ0
o9g0nUoIbSpR+prARvDgUjKJsmvBF5j13uEnUbYPaL0SF/fkisLmd/puiYi+QTHp
2P6rKJjVw3foJ1EPf1Q4WJOBNOj8kbJYk2T4lPoalJIrA7ludRqmG2FE2bkeuT1K
xHc8YvvPkb0AHfg9rqY9TPdJxF06Xryv2niviDZkOGLSwkDtjopg+qSqmXJvoXDN
`protect END_PROTECTED
