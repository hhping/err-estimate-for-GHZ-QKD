`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNASRr1tTGGj+GUpOv0HLixbvV4EmKj/MDfElwjzne29rne2KvCeiF8fPw3Ie/BE
tJJuiRldzmSpAEyvqtiLCBaGALZreCT2nG4MuQduyb0TljaRnnuoRyySb3pREI9v
yoh9Qxn7yeccfpcShRrk4CXuMBQJ5tffsdlYvy2YvQQRruF2wvb+0WWXAb6Lh16d
YhSn7rWnAisFJJLdlH0aZ5u14cdqUYVhHZVfawjafOsrLfUMnlwHR/QwQKlrRKaI
RhZjIY+PP+/lh9S4u+bMJw6kiyudgc2m9JyW5hU7ckQsATdUPyj2P5aK5BWWpyjr
ad4dILTPYIXPFb7/5FFVlpkMOgambsarS6D2pIbRwlYlhqZJUHdmUDibW10LHRoN
MiNxicR6B3zPWKAYW5yM/s+UQpppS5j/9xuuTIA+PPsOh0kL/EXMWdWrtecCFjak
uftrlyp2kWtz301NY24bdp8W8Q6vUaMKK5iyg5czbWrh2Y6uVjq6UmnMf0bHpvln
98tpvgd0nQ/pzMnBgKW8rsWFW/nYzI0RqCegpWLHu1OJq5V7AVhgzSOY964TXZ2w
kwVjcst7KRff+wzDjKpz8m/g6Ybh1Q4zv5Q7N+Rr9qmHMi3MbH0bw8HVIG1MigpW
hylRg46wlBowUea2SMa2vveFuKY0xYSWT2RuYyZQDaNdXhNKnmNUvu3Po8TMa7+H
J/NvCkv0tcHilvu6QJVV01MkgWuuxiThXj/swxG6q0vchKMG4eZeRmYyQLAZraga
/knw/fyURyAD34hiKxXJtXQ57/BKLk2eFCZ/be3dersajdPZOmfAd+vZzODn0506
7bS7t/niti5FI55EF6Ftg/JB5Bha8evlXU8qh/OEePfKk61Emfmzy1yx75rKo/fw
46BSMAyEFX8MFX/OTuRHECetWggp9SMw8Ilh1dkvzU9EnHf2r3ZWGXnbReNnjHSx
9pDZM7ocup5DbScSWQSUu0xt1G8Q5tbJO4oxhmA9KWSkjwEUBj1kbUhP+jMrAVbD
NRGLYa3jLlk70xJh+bAiyfJ72Ml7H8zk3qAnp0SkLlIOQEIc+1osxVEIF3JIGqF6
kNNyOCzf3oU5PMVxEQLuIoDsw9acTFsx5ThvDzK7Yh61oBzYkVoCb2vfE3FjS15k
fqYX0uETeaNUYJc0k4tOjFqlnEz1nzMNIhk6ye0wdKvaxiLPhrV7//zunegxXquZ
sk48mGLm6BqEaxsoDZo9+Hw+EMFpcSTgFIIkum2T4RBf9EsmVXk2wjJaLGhu6m0W
RZ/4WUtbkEF0kGcQHnX4uA4Qiwwx66XHXa4LvR9reGXGs9/lMga3KjjEmgGH1xdj
K+vYphjEeSyfixfoPK7nzg==
`protect END_PROTECTED
