`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2pHN2vahrgfrEYDq9C8eIaUn5Vqv+rz97CvdFppTST28ddbf+oOATDDT332GLJp
KqXrA6Xf1BLl7YV1S2dLxPbU1THcx0yDbDIhBqNep+5TNl+NxCDZ/2ryEYb5bkuJ
odtrBwq0lwI6eJcLD4HtvGLTBq2qujkC/NpPOjo3beTuGAFUC7didsCH+ZFB86Kf
10FpqTaIq71fu6R0Obadq65W2wXQqwgs2C6dNLLjI0+tSAkK5SaTMF2t8hMwNI7C
7MdUdfU5Rq/EQJK63a/jPzh8oubWM9q+LVyNskFYszF7R3gJwkDeP5hZEaxfNMfL
M3FuRMPFu40f1ZHdMXXlJ6iWScat9OvnWKcC+X8x45WOWKmHgIDD4FKEdznS0Ni0
yIclAHYtf9Jq4veDbTf0vlgRMhaWwnFGktJPlzedxfM3U4R75PDGyLgBojWB+JoZ
Pw3/XQLzfMW98LXQ8logHPq/5ijAs+X1I8DPn77zkGhXEzO3Pms/9TVldgzuOKFU
73lSoqpF+ge5toy2zXTo0YRA0t0zj929GsuMHArzXRRmgwz81Yc9ekNEFYfIK7eC
QdUcRuelqFDjP5d0/9hI+huCsULrQryTTPmZ3xVNYHcFATCeRW9xkmP215h+PDl3
phymTNxOWV7x3EE2d5X79HPIzvfieOyC2InrwMInitnlXiT6A6RjhF4sEn7G+GBX
Itj7TJJzC9b+VHrvDHd5nnW0ecufwECccBic6wOJC28=
`protect END_PROTECTED
