`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpqx4w0cOYLp3W7No3a6r/xQVFnUna72IpCho7EJsFC27FtQMTb6oJyin/zyDXCb
QjliVrXf+9iE1o4uy6MvMB57o1n1an7j34kO4HhkDXahgE071sWsBtvTxhEWme14
RV7WfajFzoLo6yaZ5jXlzIFNeVt2NtgrAlcfJMrd09iFbvH9bduk5AqdFwnlrKy6
O3jq6cEeJwsKFjV2U4gqnY9+FiPzDEObQTuz8Opwx+94wg+c0uiYaoODaNQE3Fg1
EVk6yur1wqFhO/P66zgG76fyDtNT9RXv9aXBvMBSKa99HhPvXKkP4gke0NpUTiXy
koeItUyUuRwCNyjiQuL0AX2xj/gINqmKy8DBf42AoavXsmpfdheCJBPkAQmGCqp2
QKzVGheuzsSpWiGAqsRSc7V52vAz8Y2UXcLSGSnhyLhuabZ42LwWMMQGgj1Y87sw
h5pX2YwjgGiJqTS+3SLZ5g==
`protect END_PROTECTED
