`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kEQuK2272vDtAJJ3ltWTIvABYyn822mGux+Er3lxXQze2Sr7bHh6+bSR3yidVGCl
9OoU8rbJMALragM/RFClK8W+dK+oZC3ENHkpDwDj40sJw6/oshvkKyWDSJn6zX/s
NbRzbvlsRzBE4PSQRUwpTHNsxaKuD/X90mLSKbIUXzqKLcnyoBKKFvDuW29vKWJ+
GoZJchW60vlai9/1hx6oJnllYkMGfmVvSALsNtGJS9llC1O3RIA9CPrmPC0ihNOG
44KkpFguvHUG9sOURdG5eSbifM+B9D009aIkO2XBt1Karg8avx5nbb08TYGM6DXl
0gNlBWQtwmvORQlICQUfyOAQvHs92QGxeYVsJh7zppe8HBE/eHtZo0LoT666gGmi
yxab/zB6BCxg0ZwTD4Vd0NKcttJUiWWqVm51ZLpBtLAYYMRYIhAbsuBWBZGNkmr2
ubW93HiQOrpya6xdPnQHFhXQJUBtAlgbQ7x0Iu/VSKMH8NlPLbQt1yyKv5QBlNUK
n8t61+HPn+jUDIp2T+/TI/ZmtBguBEHJn9C/NWKSqxxF6hH4gSLtZdpXdWFaJ/yp
bHnzzjctMjJFAYCujPqQ5Fd/EOEyxSMpnqN7JNJrtBHb4gWV+mJqQRsinQ+OevCi
56y5K4W7IgXb35l6PrMQNcH6AulsOp62kjAPFT9wy8DqG/VdusGp8dQD0BxeUskK
MiAEyTxcW455ArKwkA3JWBl7uHfie/31W81qekdsCkllFG+KoYDHIsSD8R2iaxm5
SAhL7taGccfLN+X/NSJn4ZFlx6I36nBdA0Q5BBDvwAMRBvdto3RSlmmtvjcULBbN
qshDl+E7/0vD0glAieoSlqlC9qZvKNnmC4JMNEJAsa7VxRP5VPwUNNlyWWC1sbgn
N3uZGvU1fNz7sTMtx5maQsqxbEQ+ZSurgXh2Vap4nEamwzhRZU1KOwtWKxukZKk7
dAY616+yYh4ssKZhavB+UVZay63zZhl1Aov26BPUIEWEOjfAJNHsAUjP4ZMz7nkh
eVu6dFTZFoTHTftZjbEkO7E8dXw/mUxItubkSaMKoEdCo+7k32t7wrn9pfzODtaF
8+QEugL9zaVVtG2nO1YrZWZ36xmV8RZ3oJWKxz46wGvJ9dPAIzgmPlbiABm4blPe
xyZ2pMWzeG1zT8nBSr7pvohnpZJZYwHKfmX42UnmqoEYfBCDdH+v4JFENY8DIdMM
ejBwPfVPtCo9vh8ApF+gV9YYDIeH3gmwtZk9A/x/CKr4o3HOe9M7sXRweq3lHayV
TxakfVickHAFCdn1EU81E1VdCSXRJevQcFYZ3G3AqBeNi6OJaVVCTJObOLSOZKgu
T1Blo1JRjHz9pv4y5WepnKZKp/tZz2XCmDT56l7Q9Fc9vvvACrrOCyXx8SHbpA4Z
EY30HXHPYoAfpbLqnU847Ou+MjFC9Klrd5lqXCfGF98ooJFkxEYiQlMzPe8exHpL
AFDQHXhm8YoqbEHak3SxXoi98zckT4vCSbEQVi4S40mnVVAnyDJP3ardp+kUaeGs
GzPFx2SFVDZYUkUCjdoWlagmHqPY1DoayOszSrN3TDF/Tc+cfkIx17wvNFeVw3vn
l8JVWLKTOyMiceWosJStv8RKY5HbhkejYc4ZEHF6FEnAFC2ByxgXs8SiaczdOpd7
w0Tu12PnVy3sUOISTUtEelop+vX4Vmg5tETT/I3hCH4j6o8G9FihZli8pe1dI8yI
cIlGJnlMcb6UwdarZjQ8A+p7ffgCYusG/SIXuiOT1bmDQ26Q6NFCrwwFlbTnqdX7
hxIJvlRM2BN9w1xL69h9WIO7L8J7Ob780iMzAQtQNp6GGRUPyzAgaMDU07QfyhXp
C8GK0et8HarpGvl9dBIL2Ldg0DkHZNblB8lUFhOxMJ0IgNt6PJMg9BHAFWGILiMa
PErZFpvCDJdJN2NaNk9noZx7NEIgrdyJSHdyBVMXvxkV8lwvQB6UjSsJUylnI31O
tQv8e/rHdJ2PgnpvXVeIey8N9cd3AO26K5ZBev23pfnIuBwHXazpq0HGBD/aJjSk
nP8VdjIs9CFetOZrWAksykKLjh+/OGs7p5yuUzLgEGXVARzhj/G01SFfATWxi8lr
F6lXiJuajAYtxLYHVUNqUzZZItZ3kt1Ashv7rjZuj37T0xBQUGQyEbWHeOyDqdJo
qEq0PHYY9XkMZvukeYWSWcbAQg+MG2WF5S6r1jOTg04ELnT5Z2HoJHTcVGMxijbj
OTVhHtFHOBDd2fINnqlmO87GovjkgZz0IZIhRyf4lQx/7QAdOXUhlhRFkirHDzi2
wNeev/eMQwQPn0DDNuqLQxLHpcUZCcDRNSlcV6YzbvEXvnx37IYl228DqmNKyPHs
ImQv0NbpTCPPA6g2PNWWgDNtFhvbgzHFpdPoGXOcMhtexUXh8v3bQCLY4ISTZ7Lg
2a37LjG0RYayWfqlOh9qFtCN5a8VozRvL1Hjm7LkMbAZNDEJWFzZwz4lr45xZ2T3
kZBJ2vdgJ7w+qXbMxAIfDz9re/izMt0rQQXgh3SamRc=
`protect END_PROTECTED
