`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHF6OwcbZP+vZOqjImTFPB9wU6txy+y7nPJWV40mgl2wgib6KLdRNoYM6iB1w6dp
foEuAujzk2K2EUq2Mu/xRG8GJJTnR8GxzkMHCvvBlYXa65+4tuMs9tQD/1P9p4Xr
Ywe79RSy1jpnHOz3cCYcPDYarxJDjPlb0un61G+OhIv6s1sUbfH3LC0HUxr7QuqK
ke2R8gClh5Ww9PqcBDyKpyzaoARteQrIo5T+Pi0nMlvlWEjRf+iKAe3ov2PwcKIR
Xqs3TeAjT4zILZPpoqOe6nLW7Z9juyS7Atr38v1wG6/88qoco3pSk1Jw9GwwHQUl
YMwIo5RKkHwAqGrf4yvnB7NO6kssy1YIkuAJ3msatYg68VHaxvO6O0+14KszVbhs
x4RubwLfHsMc7t+6YCXf2IVrE264v5TlkAVFxBkPMUhqmA5rvNTXCORZLWoqQ0H9
LcxB3HMytKmQZNtxKYV+8b7xNg//maBkIlB02GPXei4jcEZBIsQ1y3pryj5CIbz8
xu/z7hUjMn4gyTNbDzfJBkNK0LsuGrhfq8ZFLvOhq/EqkGpK5rhNvf1THVKSmsWO
J7kMIl8Xo5M56TRaK6rrI5zYbTKbP5V/vJGcNe5dX9LsNxLfE563AQd0hZ1ZRkf7
o1Hp94EwDreI/jvZOxpQupzj6jLtmPAXmAMawy2Eu9uMWR8G58mWsJHDWJkp+Ptb
T2aIQVcO9H0RSrjckowX0kjwZoqYseawuObbfvh6QGhpXFJZAjTpfQnEuloMg84d
C8D0EH9fuMPPSUg2akSVKBV8Yykaxyq091OIcTuDRKWYPgkIZg8IOdKf7FosFCmU
IBPWxcdC8zrL/h+WpIs5KeILvicYIPWiBTaG+MjlAMHNs3mEb6xQjBcbIgPpAs/O
MHMosOIgx4klFeZWKoYmc0m/UJFA0tMwJkfwyeu87sN3wW3ER//pB9a0MTT5hKOP
`protect END_PROTECTED
