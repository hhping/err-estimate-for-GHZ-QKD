`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpOddzBvQhUSjfQ6Qe+6VcoE/2vMuKOf2u6TWfP5QZX4UXFBki3T5AGr8XiWKQnv
NmWSxe3quCWV+mysupNa78qKxZVv+YgTRiu3xe2roy1/ol7MQc/jUpLy18k8ef+B
xEcLF8HoVioP5k+eh9NVcgMHXUzcjU7ahSkT4LYl/jUeWXiLwcJf7rKIVN9XuD5I
RGKsQkzBiUQ8prmZZK53KGvz5xAa/FZ1+uORr4pZaCbq4e2APdDTkJSoSG1JMeXH
luqQZ3///QIVm9WYJaMyHHl28bUZQRC+fQQF3/52RpPzYIBpcIU8MTCZdOBxyTm1
9SRziqPunDt7FOUPy/7WeYa58D2gtTp/vsrlV3RRthnjjQk+j7pNDqzZq/vkU9b4
J55z2HIHDQ/dXi2EKYrUdUBUZltYrIhLV/buPbPTK498TE0DxS4ynDORcQddwGkR
IfaXZnf22rn+bhLHNoVMGJA5jdqv6jrZZMDiJokrXFW4uJ432DUoKcKFciTsPOfv
dNNobQlC/Cm5bw3R74vb5At2Szlbms7COy9XPEexdEKtJ0Gl772vsTnpUhdHJ76H
CKnuYoYQLaKoFt94Bzif3SJODHSQhrz8zPOKoZEixonKWKvCxkWcV4wd3UhvHvro
Ou7lAWI/GmRbG+YPEirEVDAyiSkPoEHNcZfX4Yhx1Leptpfn9diLLxTQb56dhCyw
+hbwUs/eghglReKEKh0y7oUJdkdbUJDTnWQzYWpoFpOoLo3S7q23RlzCyD7v+kXf
36+K6Ae11OHjIg5jJjAXBLmDDWjuqxuP3T8O29TFjJsLesbIHB04JkkEA6+K9F5A
jxl3Qed8hbP8HkhqDuRiuY1Ruh30nvjFqqdP5zgsIDi9XaOfUHtOmMaU4Y2wdUOS
5CAolsAwUNpWtYPPCjdyuG2xLiBBU8oqcKGr6lCVxssTg5jCOLI8AAKp28VnFFK4
T0IjFPdPiZIrqqrxstbC6UIpTTKYj9I/JNMRyXq1n7RcicypVSiVZBu8X2OFYT5E
NNRSyipMrH01f6owZHh4uDpfrYFFXpsEtCU51up7eAFNwIU7n1ca5gkumgQTGGQd
YzKRQKmhuMWyYarwAzxntUybDwWOMkNdprpJ2ep2sW+TYuY6eW3SqYb6fobVqPzY
KiC3QP/iC43e1rE7Z3xkC0djCIu/a9Tbjjz0InfewiiB7wKX9qeXim3sl9Kgz0uc
bZAPlYYBcZ2kPsKyJrLO0HTqbarsWeV2Jfyp4yo4ArqWth0d8gE+X7vPslGwT4lq
h15IaO5wCsMzDGuVw8T3Cf9BtlgLjYcVtEW6MBYmvyGLntlYIZFfOBZz1YIAv2S3
oLDk+HFwcUQkl6IN48lFPOjmosz/pS6oLKQET9/keU0wnBKuiFqQfo0cnDeZj5yA
Nia44hv8n1Gm6PxJoF0yrFZ6I5SyXG169bLRJ8Ck0FUEkk3nGGn5zqVJGt2SICDK
NBw+sUO5qweuMZ2E+83unJFbGhAQikaJLXoYgV0K9zGcM3dI+QM5AcjcOpXZ0C2n
sim3ihJMsxv4rBWSv1CVw/RWF1ufPiKE1X7LFgekTgli2Jk2HO25X4z4l6Z2XHvx
FADww6GJCIiJBIYNtq5n/++8HuGjoeOs1VpmhBYEeFAeL+HWDLqyjCEGvH169Dj0
aeocapEd5Gsnrxv3lHrut3/NJwN54wtNB4VaVBXUnjIBkvg7IzzQdYCt/tjJC5fh
zpocIh9AkUG8FmdY5T4cL09ddcJJiIw8vk1k8TmSWCFhtN+z/7R3Ki/FFsI/ZH9b
Frj+BgVVg8KpeyyTWZzjp/Zk+aebAbTSKER83JL8fPNb8c73RUXpRn3lfPbhJArq
xfAyPFs8WeB5yxz4u1UPkCt3VXcSvQtL5+/m6jhC8LLkbLh0nIsMb7r4lPd0djDu
gA26MJR1f2K1CpGuzE7Wdb8Zb04O5VoiXWDL1yh7LPA5PuoEfyQEY3BT7pkXejUh
Iw5PMaG7zL5Qkl4sxN7ltU0dRPtXtbpUUoHzJHX6L/C2mk2W0+Sz86uPLuk4vD8u
qYx8aduwI/m5hXs1sUdWw5u3NYXxiVj6Pym1yyqGVcTZ9vHnleyVJZ3+hp7evrEG
bxdrUuebXfhFMjvgD1iHhb4yCUk2VPoiAULynL2vw6ZA5BlD2cWeDSM6SDdPJ37r
hldpXHHvgz7ZS1ilXxYfPFq9jU0DgP6OOVwxfaMjT3wWZXj8zwMTHNjDYnCAWAml
r12JrH4ZXlczp81XCarWXHEvCy94Aj5HBj7OQK0b7NuNaUg12CcPCBmCnYuwu3dL
bSbWSlaCdERyeLnAqhwFXODJT4CFH6u5R8eK3xOTiI/rLFoQvCNnMQK0KafGUVuZ
hKAG+UBAclEcstKPDy7nOXrH1ZQg9QgMwl5t2zQaF36hWW+ocCYHMx436KnThVp2
rJs4RD7xCLee90qCc0xoSjwb4MuiZylHm/pYYmhR3T1Lqh/mRZm9bGvHWZcbUayC
R8THWrY/YXnK0vK+P6Jjntdjx3uD/fX6xjQk5G/gL/jgrWU1Bb7C64XzVLziTWvQ
SmHw7maCmA9nFLr/XZ1KG0huZyJ3Jm93dsdUbNY+GnyIxHhT4HYPiK86s8OguXD4
xkVgkXStlkAUJ99ztB5xomRM56CwzFY3fbsZg8G6teSdmAxerEHSMWe/2JhZW3dx
VyOlqwX/+sD3OeHAnPx21tmeoSpNp7KrvDzft9R2PoNQE5iRxwUMXGjYbo+0mVrz
ZWSer5EJLIECMc0g4YPaBjQOSEYidz0szWh0tfVGUlip8uDG3SUAL09cZTyeRy4Z
p+E3R9tEhPh4ksYh/2/11NKpv4Kb2oE6Y71YHyMmtDH8LRrqDMLEnBTToQDxo4SV
XVD/HocFoMPkqtuyrUx8kIwBVFbcBOh0WY+snbIuXsBCLxQVsh2pRy08s7kt2IjO
8CEPHb5KJvkbYa4ZzhcAP2L+4FajD436q8aQJprZNvuYGvBrf0OavqWXTUfMiwlx
tHGSkkWOieTGDslVmP359IKYmdoDHdzw721/7zv72OLMNQN3efjT6XUCfRS0mpWg
3MNvHh8r3Mppo2JtupCV+M2FqIRynOeV4OpB0KlX7GCHbMIOScC9cd15SspJZCab
tZDZZVKJ2MRBYZPHLLx74qxz9eU29NwHv65AJ6I0D7ygv3NCykY16iPtnyTGN+GV
F19DJx9lsoinZ/CBXQPp7i8040UdYsdZdRpr098fghoF0ff/3rn3jx6SeXr4Rt71
3MLl9e3WWkDXg+i5A1ilua7HomjcVXx72BV8nG6ne1uNHi5thu4Y4Z0dYZXviOB8
s3QsCEyIH/ijrrTek7rBeslS2w01cvlO9c0/Rxa7Jmv45uEh/u1QgtjC7NBM56Ra
a2nUta2/RTvrSY4sVG1RJodEGInjQKR4hdgpEimBxG8Rja9e9nDTaRDVIo1LDL5q
nSYekGPPMYhwBokkx4pKluSk0Ix40TNMnv47DI6zB+RLrq2+7D9fDp8oV+5yGPWS
f5IYBERJjZbRh0JVcoKZaPk/+bvfm7NFi6O6zKkRwXgFv21bnxAlrj9KpZnaMClD
gRxJ9PN7uNC6JDOU/g1LpBaSO8SEIXioGwBUSrPpwp6/nXMdRzCVwTbL3J1bM+4e
D4F1vLVSEky5ieiS9O1beX/UhdzOOQDGhzvcOLPfDV/uABSK89flU0unCkIFfg5W
8dq7oi1C8JsEIh00oP+npOSYiL1o4oY80NpHIAKbDoV92v9o7uemqMkXsStMb6gU
DPgVuJ/zfeMwEJ2aKfQGFTUASHPjXyLqURYAoSmS8ME5Z50qppP+Hb7V7EU2Pmp5
TwZ6Q/xhwtYbbo/S3lWG0SCeWoqKemt9fbcH+TTdJOLoHfFecygjKpWkmp2BcX0h
kPi0J0dAZfuBrOHy/0zfdQ==
`protect END_PROTECTED
