`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPPCZPv7lEuvWG9Wna04ssEs+8mxDwdc2JGCNZ9nhDLZuUNGnhO+9uUoowm6mwBd
HsZO1sYHi9HtYbDgPuCzGS++unq+leRAXfFU0vWYVyZK4jjbU29VYqiAysbQP6WO
/FeVG7LC6jVWVjfBYW2cAkVwK/mPqvJ5O5yvHprLFrx4IZNAQK/kQVkrUbtLKfVk
qNHwF8l8rv3gpP39qTn52KMWZycErIgy149JbGHm4wLe2M2oyGXHORBiE5gMNzxp
vFHIZ2nW4MFk1nd7rsvbFIr1Do0geUa8FshFvJpP+CzhZ0Uincde04xiGdtyQv4o
zrZPSXxk1/KGriNXLp4kfxdMxwu0p4mDE60ZA1q+C6IIQJHXA9rGx18+6wmo4dtW
G9eZM446+CwfP/8knQf8tlXuAMSef5SL9SESEcnQqNQH5Nv9Kcc8d8V+ibuFJ2FX
ssMIxFW/Kg4AIzyoslUY8GcQrdqQvMfadfV7oHLPUfhE0Zc6lAz214iUSwJP4zXw
+RimzOQ4Jv6DIfUXYwTy+DVbwsm+GgyXQFbhed+nAOzMBPFQG3dDlixAXPObPFQq
ngNI654HCkOAzH/a2fDz7dvnRF/tfeyj9gEdEkvdzRikL+mUAOzaW3BkBmcsYxyV
8bHHnsAvrpo7+5V+yJdA1w38bPxhnvc9xjHayF19uZ3KdDKHboqeFeZ5Sl0isxP6
adiUWyjPnTSGq9a+pjN2xKJ6qLU+nCApZXtHDBle5gnjCTZRkB0tcwN9tiE7cAGG
hbKtB/89wdmhbQ5KpekQJ4jxBIV//sVIDdwaD806L9hSBlT3CNgn7i7xA+QVE/sr
+YSInkCuj35ELhmoeSMciHT4NaAR/3s11pCq0WABh86rQxkYAS/TM6ZTlVdYMXZj
gfho0lhSN3tHRF+0x6oAaa50KNDm3JNBodvsi2X+UeRVcOShcYmybHIh0YZfeEX8
kuwdd4PzWyTU4tjGHeLt0L+WSn6rbPbfZqDUdG63FPm8jmGco13IIGNfKi5yoijA
+loctc67R2mzna/+DgwS/qI2Y0Wy1wUmVmu9CwZAGjbj6P4JtNC5F0vWQwLc2Ktx
98y4MJbV9w+8MZiAZHbyJO0+EVI+GhmU7kEiyut5/LYvBv7UJeOZFRaaoHpyZGNh
fG4FrmjGWog3pHG4s5wVxmzCAylIFx/rAJC0xn3bHj+XZnFb47p63vXnwBgkOX3g
7tRYae2c9R+NzXXJBl5uJkSNb+V1Mt0UOw+5NGL3RH9dunuV2FCK3QOWWcBt/jQF
YqvEdysvh/c4hMGbRllCyI37YdNC8r2d3mygMHjGSd9TW5itEuo3MiNqqWUTXsaL
w5IKOdHCMeo3IkQndCATs4CW+5zDqNnDSX9DsFd2C38QeoHq+shTJALPRqLcxjrP
lwF05Xw6fi5xbjAo2mh4+9KdBIxghJM4iu/QfRExmx5S93jfIB9tEnT28Kc+55Ar
/DTLDkH0srXHKp4g4ymrpa5Y+ZelhRKFncbKGlOdN8F5lhlv03f0j9X5R02Pprxe
dFcXE5gUqiy53QmDdK55osEeG7K3fiFdxRuC0lZeyJp39wQlEbtnzhCepyPzydVM
2yB+stjLYrJxWozQR6OgIhQWpeuSjTWHKdbLGBPIGfcm2z+pzV3VDN2dro+6JCa3
4hbBr4j8bLejn7sWBSdgTH04rqZ//RluOKsnCuxBMsz6kw36bgNn90fRzWqwzo+7
2uoL8z6vIykzDr+bzKTcdHxCh4l7mb10MfdEVNwhRyn4lyhfghBol6PNHAeCVDbZ
Tu18ikuprxI36X4e6xGrjnHIL8FufSQPNZuaPG2uBC2sodsn+16u1chXU9e2b84l
x499kPWp/elyGmo1gPB4H/s6TaLEf1VqbegwM/TCXVGY8yhNYNz8Xb6ukJp6JQqJ
OnrjKiyBjHhxI9i6c/HFjsRRoh8lyo9/xkvJa+rL7NfG0MqCmWILy50bnKkr0nKa
cJBxtv7FyRctUVTxPdD4ILKadUeNREvONkUz/fEi1AROKI5AdQR8iBqUjJbNYqw5
MAMc158dBZlbXntFw5FC5wDW+azARdw/IE44qkugh5MyaR3bjOoIIfxDm50G3tzH
XXbf3c9f95+fejv7xmOlKPhXseRnV2og4PlrluLfYJEfrsomP0SneosRwwrJOf4j
d4Gql8UkjsYd4pb67Ig+0gZjGF6vUFd1JO7FbkhlJ0okquNaWgg6bKSQdYQKDI5r
8XJBMR6ia9VR0fjmCEsZ+sweiBugjNK+zQQsMOSVOi/ixyv7nmRbyRLFmgVx6gMW
0cYBbGxPB+yttp1l31/CSik/IswMrJp1Ha4HbLaHTi1oJuSLAbDaHBgXTIrO9ofG
iVuyYGbBD8KrGbMTu9D2VeQMlhDK8LcoQVubC89H768cXKK0et1H0FEpcl3TT40Y
2SJyaGz1xDW6Nuug/5D+NHLXx2kiOWcIkWDDXB+D+9smJ/g+s4XwEH3Vby9we8zI
2Jtg6PvEObr3NPlDEVK3zT4ikJDS/GkSa8APbbVs1kR0esx2MLB7loXcBTWcy9/8
iifGVMsQQsFKmObZb1ow92GJsxOFP5Ka1L7O0vFfdjbWVsi7hQ2mbHJZENeGDBpO
bc7ClkeMG3Lr6lCKpYwyUR/dr1Dg+RjPd9XLEtHpy/oKczAh7ZzarPng/O8RI1Fj
G7ZhfdkxR7/h/Jfefhon/lPkX0WeVYEvzJrAkzxqxYc5rHIrNApkiHBjpfTDXtPm
WHujUJtqlfqIJXaiUrYR+NnUUvSDp2iHYeEtJZtM/UedIywm38bzGqzVLmLUe8Q2
CHsH3hL+L4KTT1NpRir+AvbiFaHLe3CB0TyRhBhYSgTA/UMi4ANsW6nqSdNvqwax
E1W1W/IZNYSesx3UKTKPFgJT+Kw3Ikgvnae8fYxPy/wWEOqwrd5qF3gIyVGUq49M
Sxi92ym4JcYKs0+vUZbvnB3njfTwnWv43CH1L1LDJnpuG0hcTgxnaTGbXJZaQbcS
UXoVYn+1xrzqH7X7rlIfCKt8wJVVGhSNwLpPADPznT2N7IoZYIF8fvkV/ujIv4xy
YfedtEOglWhKmgkFbNqMlUJtl1KzG2IoodAqTTbq37Y4og1OOej5uXm7dB6ejEnt
jvVmGZIlc7Wrlx7WKs7ZXWnVNryHmr3K0EK3tSGVTOAHO1VNt9WUkWMXK45V7zep
9Bm9JqWhq1oU2npO6fjI61R/BfW/pIvRC/PjdxyZqlKs0Z8AuYvR3reTFkPSi3rp
p6AfA62qopqmpLklJ4Xh+1Cl+ZUYxMLFLKcK8SkeIGrd5zAKN9G/gXQaUeO27flU
HUmO/BjbpBT8go0mJYUYRyfi7RaVlT1Z6L+/K4vfeiPawXu+2j4DMdrETNyZAirh
fR8NPQeqbeMdFBV7HHYMr6x7QpxVpgf/g4xrDBXF350fhgxVtezCUaXR5IVJBa0i
45BiafWnhR0VcScEezk0KIvXzNnkMd+3sD5dLgL+F01nczv7CgMexU/5y9NXouWQ
6bLmZ8Roc5Jr/fOta8utxx1LHAzYRdICf1c2X7lm39ZY/cbXXY4pJp8uzqKtqPOf
xHi4vgDB0sdC00Bth9hAxQ==
`protect END_PROTECTED
