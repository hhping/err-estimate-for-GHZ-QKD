`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahyvoASd/ONLirFX0Lj4tTOw7eDRufcGQXz8aN09kFx3CGkAM1MHvhXho0iWecPe
CqztG/j+SiV6oonIx4D3W+eGUZ9zS5zhajpLKzk57BH59fLAWyIyo5B7bGDJnsxo
7ZlFeWKYMg/spaESDnct1VxBAgEvJELC8Vl3gljeWEzbWkw3jaAB9De8jBP3bJ38
YiAUK59KtEe6PoPeKIHZ6Ou3aMsuJe1LvSmlFDgtou+Hyr6iwBNIszhZOHp0Pcd5
QV4OuQki2o7O5Qgv2q7fX4SaAp/2yqH7FZ9fInKi8RtOGcB86JwKc4+DKg2VcWhV
OmiL9OY5nTKKsu5wCCnPVImL+Furn2svqi8h+BIZuAkQZ7db3mNsUgs7uFfFCTW3
dfPqoLOGQTq3sxO2BIs3NFTtX2p4im5HQM037SIuqUaj9um4UpboKRv9HJ0v7w2Q
1okpC/P8U/T8icWKNMWTCDkvRov3u8l/BaU2teNSf5bviUoU5cpHSObxlGzFsEwq
fvB8JmvmdOZmitVBE1qa8yYE0QWXLetZyG0a0PoQbLtU5sAiE7XmlJxVPHtDpdow
BtP0xEjqsWpHNQJbZQ9s+S6Ym8TEsRxUfbfxpzkF5OhOMXQdTPIwPzZoVuiZfZRE
lbjQcBN/TdZaUE+yT8MH7+yHyRQTaElEJSKwSiTKsqIxNaqE+AHS2HIIHmTIVhN/
yafXAX0wSwYCFFu0ZLl8dX/FItPm3W4XGCdKqveZsCmvb4NabDdNpPLxy0uCsfXf
dn/ddCMOr2XrasnN603TJNJQF7+GwE5LDDyrjspy/MWTxx/i+06FbmPM3cdejM2z
jzQG37qaXpgww9CERRS5E5MUThCe+ByqzJ7Vk0J9LbTO6ukz+eSZ6NDB8CoQjtNa
ujAKS6zXqA8u1Z+o0WSgpKmmBAEP3OLxVnX8EJsZ2D5NxC2EIQ7n3T1ZROxBdxjw
HwK8kSjc00J96J1mx5EKka3qHJgmm7U7Vg/7kc0okNbMYsihoyMIhgMv9QVU8bEL
KgsKBV+guw3WpJO5eT+q2hpyli6zBnWIjr4C3wCOquLme3rET1ZG4knHoY7FqmDw
pwXeQ/pNsbXAMXpdduOCY9CvGdNhEuI25u6EJlbBwYgZrL6duxDNnG2gwCLhrbE+
xXVaN2P0sRp0qA6KD/xMPhi9u9WzXF8mmczbKOC1YzDF4EYUl987MB5NsCpU7RpS
mhWjunLoAQFIHj0tIdF7RwBjI9kdhx58K824O057rxuFN1K7EudYEr1fvltPfNyT
AfjwVx/N4NASDeDBUAkJ+L4uH+cz33bK/6NoyR0dLDANQn+kvkiOaKV+FR6gmnH9
h+kqvfqJ4K74wM2LdfYWX12ff3uY7TzpKlm9AOc2Kw2XhqqJfWRcCL3X0ueLsDH0
1QOyb259s165xWmFOTQuJGdADZI3FcBpRZ4HkiUPRrO5xTsOEERYdEthgYIyDC5S
MLpqCF2cm6h8jBxknz32aVbbktjFWjweDuSRNJ20+YgtMrfpd8dDOuWGyLW3aeIc
8nUkYQdbLK6ct4RqsKTuu3zJNIqIM8u+oNgZQ8ZV5qk9EKv2POEi3FatpTL45l8y
juy0iEGJE9jIs3mIJOCiPbJyXAlEPxBUtvo1poEZpM/FldplhhDpxFQolgqRYWbp
moCnopnzTruJJSPWOpgUrAY2XkitWkIyOPP3a9hFm8unWLqaaKAbAUONTzqJgAC8
2UvcaKuMkm41kOKdeyYmoFpBM4AiYfmrAjdlVf4RIzxKBKVumocKypyItnj+xS1C
TeHg13dIO2rTRq1dLKr78yuYNwoeQbovPpS1oLZXYZOb6vryvMq9b5lnQv7pHoLc
nT2cR4DrKg6WpxGifnUIABxfAPWk6nIDwU3lDRd//jqvvOjm73KLAsA93V8oqmai
V/eWtGs3Z1QEWRbhvMZW/E5mqIq6ziluOQmk5WB0GPMf8kEvw9E1YiByoLvU7Fqp
Sb9Kvns28zeLRD8kZEYwRQuNRgo1D1rV7Q5BjqfvvnefEp8Ecycf3XGKTFLmWQW9
wkOaYr9EukHp5XdzO83TEG6d13PmddCShJ7j8ZwcRNGUtRI6pZRGjrfL06KuDkb6
Pb9LRv0mbBo0lnWbuFdjofhwBX7e/yAOOj0O5Im1uLDjqEn+DNa7u4id8tw5gTZ5
hKxLfNlVZrEnBB82TFJmkpt0KEhB11Kw3/TNR0SOHPNBugEcjxOSQTzT2nEL8abv
Z4QtapZ6rFHvkUecq3VxDCRjXAV4FkukB4YUdWlKb712gXDiny65O/7sOuc37L7F
c5DBF0RUQdtVL5lhp00SfCRTDmmZ0M4qazF30FjIHCZ7RyFAq6fk8vLDWtCowFC7
/f3+YvxRkMj7d9UCZ/50OED9EhaHLXYrIYx8ogvbuVFHa+AkK9LJwHpKo/ojgMr5
BA07B/auMKxoDCAQZVXaF+GrkGYXCJDrW+qmuOFCSm9x8bZ5Zec9ALat9+mZPHKa
Gr3x7QwM4hc8BQqIrEKYpZKfLiPA+uzAukxOpsVRlrE/HNtNzMWdikdaPVsZmK4Q
7IlV6oGyXszjbn7FAxh49PGss8ARgUlpxzffNE97bv8xqwkOnyVKmEajSaLmjKDS
1Tl8HUj8c/GtJkkwtl/WPkl220XP4z3sols6yCtVwC9QNdqfaknL2ErD+AZ8MpOD
WwrfGR/OOnGJzxK2Av2yHxqWJaMQ1VFYXk36ePp7ToNP1UJxLgb08XWDEAzeKe8r
/5VR0NEtMtq3mcvjHcDfB8PVjng9xnmmLskZ1g3U1GrP2BsCQu1zsb7KicY5avmf
RzkCpU5NF8FrScsT7M7pzcPxEleDwt0miBnpqjZWu0abhWxL+/thd415wOLr48wX
uoDcNRCfw8nl7pDoQrfm4/a6als4puC98zMrVHtoUZg8MNX/jc9WxmgoNfAC+KeY
6rECeyuVemmkR/3JwzbU6UCCvGSv64mmjQ06+OS0k3Ubc8IkJhjRPrIuG8vQkx7d
HjXTLXNhLs+oS37Xyss0UxwhDvAnELmWMtSQtwKy2hQbNWAlDHGsYKb25n+3a1/5
+AZwecUOmaOUFTFuYloVsZx1pYuDi9NUu1wlfAZB8DiwbboG8xkeAT82LS0nYmyU
872WXrYvBSIXjo0Ypul6Ho79eCacltrHaQUl7Ym97TXN45tZV4MCnQzqmjP+epBR
gkIEl4lhEFdYuap5b11C0LSXWUsZWXdx6DRXeXRZ0u6mvlHc0s7fLJ64gAJYh9hv
myhd5glLU4f00pogYkPz9Sm9DkuNikyrzkwkk11cY5iQsJPYGNvkcnbKcPeMDSsO
MiFjPAdQNvj6yi93A/BE9fmXCyUkfGXQ46KKZrZiMtpGpEghgHP547VTy3/fg4Sq
R8zTBT+QJyIjhzHZPEUzgUVeehRMg0DCXK4diFi8trbaFaYfawd5qg/oeg2jvgpA
RqZnqv67X84YBw8hoZBaBxkSviaVR9Sr0mYflhDXVYbSuBNiCi3Pap6nZmm8wizc
P/fXzVTIy68kJndacFZWBv14r4P+PbeSTlHSMSUEA7VvOMTxTgcrY2KXVLHdMlcQ
sS9lXCLFoVYeVZVWqtiPYC9e17Cv6MPYYDEYnN+f3C/2xyz1HXm+Bp70AsT3aJYB
u5CEOnyKh5f9epu3f92tjV4Mi3czuHGtCj9LIrOZty2JSWO4lNPs9v3qOzd00bsZ
+f2P06N++765UOEpJoQBYWiwvAh4KVg5QXsYgSs6hASbQvxzy7Ydxl4rgTfZoGFT
GHTFSzabtLhYqEi+Q7stT/wy/j4t7OFrLRCbxEWZzBS387cFMDLs24tpMmn9Xr5T
BMyGxBkljSh2xkRYLWAF7Hua7YfiFoApI32wt1MDCxM9PAEK4/RKpd6FhWLPin6B
BNgDdtvjAACSDzm6F9MyDxD/c0nGKPdixlwm7q4UbS6lHuJ3fCixU3f1MzRCWG1l
9oRpbkZy+Ck44YXwSuLcsZ28XTBduHru/Vyoc+AkpulK+nPvpQ26LpRGQHHN/kHa
amCJbC/YroyaIfTR56fvIoL2W/3K3jhMIKIGI6oATr3Ilr7rbcOaEJE1nRQwFIDL
qZQexDmemvQYntwz4CfFPHRfcJP40nGx9XET9ujbDQmKDHhT5tkRsJ6Ak2FoOOo2
o1Ucggi/x6jXHf2aJp6zHDHSfV4c/lVQoqHjvos96yShmQpQlZyt0LF3DAnN7zes
rV4MTUyu+smsySqKEvZxEMo/dethP33NVvSLUDqhXcudydtCKM6XWy2KXYsQ8gzt
TQJ9OJWASA814Whn3i0eTBP5yHo7Q9nSK+lyC3ButFojI21eGj3oz4bcqx8XrUMU
D0tdpRgzrkOpDrsA4Eq8ydP9RcZxbPuFccqcaxwXqtPFHakPoFaz6er2ATf/HzY4
JaMqYla0gNnQKvbs558fyKSZPHm7Og3UddWnWjPRiXRT2rLuEbHZpyI5Qwo97sc7
F4Z6mQYBB7C43PPI/5LjxO/Ss+K901yw880GYoSQGbeaJImwy/VgxOc1KKXkjI7L
dOM0q6awSqwz3Z1J9HcdS0lTZscMQjnimtrfHKckwXlEIdhyEWrmPgeZKaByBiEm
H6wiv6XgBsUHp/t9xVE7uz1Fmy+L+Xnv+duohKv5ZX9THQRrLzJFO9AZPzAyM72m
IsDX6gfgoxb4Jy3eGDnb4cxKvImDYUzXJaBnpX+jaJqdTsBqAIXc7Oypx+/Chnx0
gVgeoUBzo4H204vLsgkkvaxyTyXT7vjx6CHqpIKvrbuz5yfWoQ16zlGMw5KGe9B2
lX65Itq2kjncMsajw3ru1Xq7IY4bBp1vxr5C3URqH8ASsKbo6FvPcV1xUW1kw1AP
YQkINDR8eKpp02x4doEcG3w3+UTSzFheuCgu6TktsbeZjt4PJl1PvdywJl2zoOJ+
Y/aC+0kUDWIcvcm3FGbdrNUOAzRekYnParQVp37NYXmuZfW9hk/vQ8yx1SWaYG0N
w2BEcsPmkAxTJuqV5eH4qWn5a3+FbZbTPL2X0XMdOg3Dmwva3fERJkoQEl7RUtOw
EJlOzbNfgFVVcL2HY4kQ6lhlOr4gFbOn4mECJPexDWCscPa1L9bUrez2r0GnGKzS
qp40NXfQeUu6WOln0S8swff+r70gASPl8n8wfhNxokWDxaJCsp23zXHfBos2PV0U
XutFPuyE4v3e9zDU3jFQFHDabyg6IEjlP/TN+ulnjs88Rse/I/rEvk9HTScl7i+I
8oSVuryLAlBbwBbujOf+slBRn+LoJEeTTZhpzbuKogXGf+krm0Ta2R1PEqR7KG7X
lZz6RaxGDzczslrqJ+ayyTQHwGUeAlQt8FKqzuYNtWvb+XPWxncoyuEQidUnbgg2
aQmCckqGPUy/SGIGk9LtnMYYR7S5g/E1fmKlgXeUxaQp+hpV3zOgeUvteGqNB1Cm
4XBr5aFNuuIJh/vKf72XnBB4+RcZ70wHkB5e9ZgO6yc=
`protect END_PROTECTED
