`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frLnDE5GyX3Jzxl7eBvu82guztFQ8CBII5RpoNsZIJ8F9v/ccVBjJ2Yz7EhUgs9B
OXmBPHrgl70fxEERMAzpjzKo6KYAFvB6BH2+q6vs5cbI0OPnUjUiL5ZvkNZ4xfx8
6MKZ+5ajbfrWgM8bORNQ+0LRfyeizJToCLPVG9Y7+v8J1Pd/Dn87z3mdfk5KVoFj
gUaYNmXyQdenjZzq+IdcPcQExJVZXn6jyXJBhtI5HT74MGbJgxWqxURNHPs0iP84
C77xTJt9cY0HV8YhOl7t088Z9krWDFtMSqcv4JMw2WSvjRH5xdIgAD2NDN/1NFah
TpfkLzxjzlptZ58ScYVqB2LS79awIzm7M1xcLxpOmNeLzzUFULpCbeHfyqg1SndY
EjS0MnFw7OnpzO8kqnmorAh+ZpCRt7QhRM5DX89n+9ZCisHP2ZQ1l4bkEIiVCgVi
9DXgvk6UfYISH5IckrakzkrCzTX4aDmMoy7nrkDS+PeDcQSMWJI+/NfLduUKSTCw
lTLJ2VbAQZIg2KuB9rasGDsq/tYJUuFGlNBd38i5zveWtVueMPfGvTE/+p3wdizX
B77lwV0KdqEzi09FdHsz2W4Jq1Q68P5w84rNZjvc2sldUSEPYsKeMj+tyoNHNAlP
kueFYmU5u5ZR3qvUUyBSiaAp8FEE7CulPaInPiyhmtZLXa09gll26iGIbu33AAXS
KypNNuUpv7C17WIxeCsKGFiHtNghNzIJ9dD4P3Phis9U7Vvw30fZDnEYyXD3nkDp
gU2iP/Tun4bPNAldA6U/2D9Ncv+LJhMEZx24yptH1xAkIfJnVLxW8UZUod5FSe40
itux8Y6gCZzbM+Q7gxwkUVBC/580+ZrKEkVPOrjNE2ctw6OD7XTI+GKLqjfDswtS
wp6HE0tebszZeeonDhc2ciIqxnVAY1V02MEhxjIZGxahyRxhiqCoOZ7VHdey8Ai+
t0l71dQ/bNUCc3UiLdSvFe07s9PpjQAalADyXJvzE+usgXKYblOx0bqpfCDXbbz+
oSJGRo8n284HIHY9Gakxl+oyjNVru/c8/mxRbsBuSWrSnsoKE5SGZpi3myFy9UXC
hCegkzAnr5sxCQJGNlo3JUHHkS1tZcf1c3/UvCTZ7p/eXRlsXqIQ7Zdzz1jm2U7i
g138e71KSU+1hnxreq1yj3jZ7aaa7yZRKwJy8TSARx/JjxFR+afKI6mv/EbmR1kU
Mq2KvjCZIY6/w583EkJJiS4p27JFJVVXQJJH7V7ReSH5DFLJNGC1ZDnA39leMiLs
fzMG6KwUtjoOyMW8Uhm+hkV8lWZkNMSWf6NQvOvPCehVxq+G24VjvDMIUBdA5xwV
HRcreyVDWfIavxbKVIqiWVGdFcg7s00LEg6ItRd5Yq8S07K37Wc+esvUrc7pqGrD
fd8p6/3AEygRyPdsH+IV/t4mM/QS3QhHmR9vVknS9HDMzhL+zZRrNzDPSKWa4QRU
1EJJBtyOduzoNBz59z3SqQgLl7ks+pGOJg1eCAl+OT+T5Zxi/VZQBDp5ONlLwhen
XZ0jWIvceCA1V1d8+TVHibUraHAMoOLhezDA4gw41769/mE42pcWgODg+RtNGUxG
PujJ8Mc3vljQ/IKlue8l3I/UfGvz8EYv/Vv5deItnFUz7BRAkqzNkMEoD/k6H5zn
Emd2jUCWaTtPdO5F3gBjRoMH+VYHAl/AmU/tgR4nhXZkVhuVYt0wUhIFJ3Tjm41X
TLG73VlvU50O0J0G8AgMKmPhsBUaI3a2KqBvuUDplbaiIOTPvbRzeOyOKfAE1AGs
cgPjB3wGzTd8QTuia/DQg7YySffKXQPZALgbyLGLrhLogiuydvkbweTWfu4aYgAt
h37TSoaH1JtH5xGfGvaxbTxAokDoCebJXc7rwW6eocXis1bBaVpxd41bnKxixSvJ
rNwueQU94cUjtKiD+JdZmsWj2CtvU0QBffT2aDFVrwkY0G4TmLTg+wNt8KX9K2dN
gcrBbPqqnODM/WnyjT3eqscu/aVe35FFR6Ke5pe8W44lYbS190fjuOlF5msS+yp8
hfA2EGoArW5WcK60ts1ySx0ZwivOA92PVG7+gQI4UAoBo7j1PhRvqfk8eyZzGEG5
sHBQc6RsK48EDxe66GDtYismzgRsFWHgmuVg+T8/ooMrzYEdYdUQMgC6/y7gFJcW
i2hg+aULvyLs28TdmFA46Bi6qdgoJoZ0fSR7RcB+LdfDIykcGXNDDbUAkiuV0YnZ
ue9Cx2cOMCcVSZeT/OfEqu4R+ARkQdc+gwx0Pv2+a1urw45n3aCp7j14W7pQ1PTo
VoK6BrKFKgw5VAMZe6UB7tyBQ3Y59AVucEMh0cNo11+aZwWN+WBH2Gn3nzAVi+oR
i1WWyoXSx316lAm0FlZA+0o6lEL2V32H3jdtL3UPoZKEuLubcPzNKSQwuYksh0W1
yo+ZGdNj506YlczoadBnR52MLoLCrg9um9Q0wZGu8OnhCiwXSJ4RZTjemnyDbtvz
ZEEE3sVIOCXzyg/Z3ud9FNvJVQkK5oF/5mXjH1iVRO2QW22lvIRmLud3jLqfEuDO
/O5u1vlktRFGs7BNgM+N46vJkeCxaJRCiGgksx2+hxxY7EXHcfeVbpqrrzzAa6nv
B2NRKoie+swRXUNdE79ZQg2nlkD7tw7Dne4ulmb3FVrLxukmcItZ+7Ad3eSbwcg+
SfDEPsdUUpTtExDtcEZvdKazgNoE2W8zhGKI/lfxjACfVdJBDOzXGmnrGxCMTI5Q
GvFPekK4EBQGOssF3ngJ8TL86GSeHAqeMv1VmuOLjxpFvAXTy1nopUCbIwyRey2y
51Hu18+y26+ZWXjE3E24Mphn5CNwzFCUw+px7DZxyZ/4asdZJjqH3PpOaArtu+kl
OBK/Hd5tmxAhU3JPDzOMxy9g4yuJTEWsRQNfzT7exA437txXvZjHC22Ii52o6qRb
QiJ7UA2xJvcMN+M3K5iVnl4P//dSroyj25MEsjdXVerhn3nTnaWskiax0OQqyvKb
33f9XLpp4r5/BdKrMH1icO5k+MaJOAgdOKlOUhll7ZSQACbA4DeENQ6H0ozLaT0L
QbaTSbtX/+DvdPlwLize8aMuQ/lH0dUfWPG6lJQF/QMjEiQeT1U+hn02B2MSJzSM
xGLGODjY+we8EqjxoPcNjHSyE/LbK58HKs+tU+fBGmhx93+HonBMX5ug3+6zOtrx
JeXX4hO6vpcFjUlkM58Kg3xI5N0j0gJVBvu024pnHRpvBqVX/jYphCpyNH5a80P3
eOin61EYlKVe8lYX7FW24LKynWaEanUZtcoKdm9QGysg85zqr5ZQ+Jr1nK8Sz1qJ
YVHumaXYFok/GpBHHI/EcGsTzE30an46RNfKk4JRK/4lM8RIO//GCyt32l1EREgv
1QmpMZVq9I/vVyEAWaHz2vU/bLRF+eM3XmW3ad24Xv7j34S3QWc/3D6CPlCvS6/8
1b+G1jGi3/4a+kZPMB5eH1ZGMfsPd1iakYJ25J2hbKfREPPccJuWVZJjbW6OM8p7
gFK64wQDa19ISL2WlQ8gIJSvLuck6ADCd7GUBZqNjzxC6OoJ3oTREuE7wgkB4yKq
pREH+v3WskvIM8t7+RTd+BNXMlNa5e+EdtSe92rDrfQMwjMG2c7CV803eg1uS9EA
XfXWcOYW084/zU6uEC5/G5EoQkTgYl/7Q+O0DQoIV5YkW3+jU9xGYJShdGAu7DIk
ai30/K6wOiCK6U5VPlgFyml0XpNu7Pmju5RAqL/nyJgfNJK2oMXwA4A6gVVK0qov
z9qiyUMptytdIr8wvJ45ADIIukh8IBR94Ul91heUo7w4WaEhgosP/BDPt708v1Sn
nOerVbyaviBkHoNChiUgcUwGeHsH8Mgc2PCpWmyc49Ttj0wRfHPgtOjC9YcU1OqL
rCuboyq9Qsbq8Rd6OiiTS2PtFkDv+5PvCvnrbxe9ea46PfqWnMzafyn86ea+8mtD
M6gmbAqF6IKoma31W1lbKPPlHpvdu+S9I9r6xVRkVEO6zAXA10AvOAWoMl9Agcpd
joB2x+TtCLHqE9KsvGQS4kHDzoi/lelguYLzfdj31f5M0RoL1l1vClW4Cj19nmts
Wlu8DDG56uv4vxPtwDkfHJkZQGKr0ziRWRqh1a4P1RrkQ6h0z5b4br6xKXGRP878
dtfcZhIFvXKniARD3bn2Xwf3159NXDd6eSbHL8PRf57HFcp6NN8kZZpJam4fIDoP
hUQjibaUbRyPcu6AGmWex5pqrx5NZOer86IauWyKnMCPcb6I4vPzYszPsg2iCsca
hIQVz7XR0eCkSrAlPVxCGUDX05AqPHrWoMBr98N5CvRpb93b5AdZHobVGB15TY5n
b7LuLcG9dNIEFTs0JTyeL/yj1F7BSXx1MVmOAZbLrb+nzdOFpqfSInAMEPo1TYiy
fw1wJKgcml72Rp94CAq0/ZgVIm0OH6gJr/yIlw4jTZNOCmj8bwkpr+tSXyqFLF+C
eLBOD4U+sv8iGP77LIfglupk3yoxiMZbuSr+W9GUHifUA9PU+KBKO5tTARrH5nnT
GRKRm66Mfh8evaso+j6YJgU2P+E2yRYpN1b4JC9yHNbJVHduXX26ZTriDGUD5Ws7
9EpTbRKPn9UtVQdi7NAEzbpv4nKqsfEHJSDAGtG7gnVB75Ro+aQ2lte3H8s9l5sJ
DZ+rym0CwlFT8v+qSDSh0xDXOD+kv12R3iUEYqrGaomHW0jW7aMbzQxGdiFbZ44d
AzWhcZR7CcWr8NLtelVd5MLN2serX5aMGcwyrPOCM0fuVIwuP08a5vBHjvy3NJtM
i7lk8fS9nwjiahVssER/0H4MHRI0oj2bOL6IdPx5L8YDM+PdFTmiTKH9tU8SWcX1
ZI+arXDjnCKP6C8GJmsvg+kK9BSeycIxxQ5NbkB1rQTQKVlFTyq/kJ5qRe8kB41y
/iR13ew/cNP9rFNCMIbnovg64ruyk/AS7EJ7zrrhGsYbgSOFsc4FQJ5hnlQ12U68
FaiQvxT4ne/OKImKEX1IAc0dABc7PgXPBDUxFhLPY+z41v0B4fE9zM6n0A+mIv4W
16S5Ms1t6GR4xcWUH9GHkwMq573yidFJFCC00reNnrwRUh5KGUVcQHSMop6tG3Ri
3phvYG58rIn2kgZo2OyTsmJku3Scz+wy61mbrB5QNQNVuzwRVf2k75WJ8lDIVCRF
M6cCOegVUexoPseiGuv3sYe+Ec4p/CHbw98og1VA0M9n5YjTFFyptCvuJT8X7tF8
I4YqgZd4Kh85e2ZRYLjbbXl4q3rQfFuDnLgcZ9foHGwEWpBvZ9Ccv8T5bmDnn2bO
gXpam99wG7gR9ZwPsc5wn7gDLSYf06EltApaC/ObicKyNl03AP4w5eGTz9ws4rix
q60AhLl0aMq6x3+5XJvm2PW6Pt9zYrmUP8aYcmUDnaQv+1Gq/8byaxtYl8CXFuAk
uRF5XbaT/1+GJN41JfCKAqk+CX8zmYmQF1EFeBK5J/sZ1MHMDid11s0AoFKPpprV
sXXkTFsDgkesGF0JTZ/o9lbIvjKuzw/l/mgl7LhTu7FntSsyJ/0mfZfQiW6aWLWJ
aosDI3wAsD9v1yNJY8159W+lNRuF2LkMVzuZRpN5ZNvfAzyc1a2knfZZRHN86oKQ
EH0+lK9cjn97BQ21W3NXor6JoXgT156dKPv8ShkVZK1xLYGDDGpo1CdA3EwzFIQd
IfO/aSlLHB83e5OHm/wXKrBoiZKkkaZtjmckNd0f1AljYUZYAkdi+WAbJ6PAOqPQ
FPJgYx2RGLGQB+V8o++W1PtJBZ6BDzA0LqLZyjOg+SoaUKDaATO2fJ5P91Ld2dIx
Wk3y5Ow1qJ5OZdWfvhsiHVVsGQpN6q4E7BsH4CGvflbztApuRF8tluT11iS65WhP
YW6VOhT80rga8suwukvJeG84Fghf7p3r0BwazOQPwCuUTCMeFrBm6/Kr4erS0rSS
23+OUgkXCZ17vXiXLYqx4j2gXnI14oJKvpAie+X76GQIKtZ9C9w5AwMjTusPvuuy
Y727IkSrZTSwQ2d9FHVEXaeatVnNQr4Fs2i0hg9JH5A87Ldps09kyYXkAxLy36VH
KtSNbfhQ3RemCe4xRsbh2n/468dSbUVeVKiBJgAB2YR8LsXlJVMmYY1EkxLbc6UY
4ccnCG+ktXhm1JlXzEeZggKw6B2H7PFnVScNlF3GIgnFz4kLJ2qC41EuZLG3ny+b
ZeGkNGLANX+DutlCiK5yThVNp/QijDmUs14PVfWlRd5pcdx768ny+0iC/yJguuCU
NA0dwWON/wni8oaur8M/89t75aYobb9Y8ct2+EHhH1cJiT8aUPrCI68oAckdmNcb
4UC9Y00pRV0Cg8kuiZwGwpPuI4qXZb8VuRQe3M/SI4PAsw6KRYJsdtCtLms+85lD
Kf9evdWeK7LmEzibYw0vDmdYZHDPfI6j2mb/y/7Ew9bWkLt5nVX129zHcsAXpKI4
D7OItqzZschgNcMrzqvJByuurjr+s4JauJygXX0iDfg9Ec0ntIeR/VR3is/B4Mus
tqUFwyVlcWCWuZg+dMZym38HIdxqqZSli4g6kLHloQq6rffdRRFd5Pzrc4zn5LDY
QYegaA6sNNjZrEg65osbvyqLLFghZ64IGMv++vRd4umYCXIB0j8EdrZFyBYTKTUs
otdEHudYXSgiPpzcQEQTaGsFcG7I1WWd5s0qovRI6dwbQH1OlO7QXOQ2sQXjzBEm
k3wqBv3a9R2y3VV/JqAsKne6sF7LhSTYEZAWrCv37WJLUtTdRl2v6de7kUIgIhRm
HY8jwxiQq++btODuuFzKtRNuvvTl+gj+6j001diZHxEB2x27lsiFtMXi3/Uhha1j
oRImJ/DM4PYkMbTO0F0T63Zcq0tjLG3DRDyVAVtRCG04eP9SeHJ3f92I6c6ZvNGF
BNkigJr62RNB8/8roXb7pvnF3epkIEfwBildOXx2j54yzV+zZywqmn9hax7wgfo1
ENHZiIwJD2LNNJ0tqeqxOpCuzhdBQXP7flMJuV2dStfAQjZou/NMLZnGB/e/hk3x
QQ+1s0imQqyrRDilI8BUPMUPcRILbbnbCvPtf7kqa5yBVMZ6CniTYL1Y30m3TlcI
yZ10Vh+fHIpCWRsvva2CcyyLoatsLAGeReV8f2GQtnKgEQ8384/i2b/apaEDuoZ9
IAlk5s+zwxVosB+pWIuc9wBbBaZUZ5pVdANo6/1d/7WaUTdn3XPpoLYPUy5YANHZ
tDJioe1bKk+UHGo6zV4idSAJOx2tC69X15hDqv/1j3cKAMRghv6GpRPLU7eyY2gg
zyO8vUx31jGYLXn6Jei3ABBht3acKqz9b5JwSCV6RW/y2VvO4XdDPHKewQopRQqD
HfqzEOIcMq7e5uUjt14H8Emy1T/2xzsiwdHkI8yiin2e4dRZ1OS6kgF7OlA8q3K8
tDq8LzjrXBRNmasVXGTiYTs0ovjV2oGGv5mbDLxQa4RYHUiYrXN8j/z6S7eFE1df
fgQmAPZl1bzTZnSCNn9fBsyV7OytRJe9SSUHSQDkT8VFRzPlneVI/I6MxqY1sC9j
QHV5ud3x5k8GiEsJegFu617/MPN8tjm+jkhy1rZ9UYGVIhVx/dpkb3xFQh95j+JU
5CJT17GjuMHMYZi2va1XsJq2x7j610xZgUutSnDSjeGINoiLyKWvdPnnLkKUPKea
tYwrbFupFQMosKcnZ4Fj88SRXJcpA2F1Og4bBcvIfAPdxLvl/u+Zi4VTxLGWbtn1
DzQYvAX99fMyXT+/1bINYWi6zY5qqgmeUTFIJsnsUBIQ0STd2no18m6aYnxreuuJ
QxvtMKffs0s4HEUGqiUvHUNNzsTo9jR3a2QYrMovQnyTLnsHE0eDfFhZzQ/Gs/F0
PbxhKC0+onJ9gQSLBO/YY2sRbADe6w0ZSMY8FImIBZOnQR15UqUM5alHkVKbW8jn
6r6o7tVc57z0on6Udl8beYOMCowQH4dk3ntj8qyypL/Bmm/Eg4OOIksWR0fMso1W
YzfGptxlPwepQJPqpbbS1jlbgaDymQQDrKpLrhBo0DOvojuM17XsyvGI1RVngm3u
ZNO9Fn8rjj42Bm14LoaXqhma816n+tHu0ZE1Gl2NyGoxNVBR4qPfx5J7tF3OTrwv
GXIlUuvtnOcnoNKAuN2UPikf/Lm5jukNAyf80qgQbnvefyPuZ4MAOiJ3WHPcM+tI
ZvCknQTfQC8q28CbfjMwuz/Wqm8Vrtz/JfYwtOGNHWlf3OUtyjw1OORq3SsGgQ8E
5dTWt1VorjMVkXQ5OYQQBhGuFdLdDmVU985L2XC3sI2c3lAqmnynD+hPKCKXezUf
sF6yjd4UXTo4JnuTRh84LTdIiR2TrAZQkUE/rOYesGO5XiHWJh0Yfy2ms5K8HGYe
/CyqoyUuQozTR0BfeMBNZ+SsrPMHQiSpjSBF1vu7jKtMGO9+gOQPvqupjNrdOvqz
e2EX9/lxLjAhrwzvh6XVGSiJvqbgsdSt747aHZ/5kEu1+xALbHShXq1tS8NjPEnu
cUkf0erms8vcUNG/VmB66E06JYW/ZWvyK2x7II/ea/fM+NaEBZY3oSOHTfNQlmcQ
3Vp7aCNK9XURO2RGITjN2sUsw17p2oFj1aacEfmhlkiUGLOji9Fke8CdVZgW5k9M
42OKROy6bb2SmmvLB/yTUHC+yhGqRfIA8bBmSW38SR81UpChpXNqB5RxhHLkkdro
xrBdnplmxlsqmNZMx7/JG6W9JIaTy7mlgCBGERMzAVQkqhU4ott3THKXIutA27k6
w5a0xoKG3S2Yb9kDsIVSr1oq8QkZdaJJ2pTJr5nwDwHH7S9dLaiFTHJKzBAbnnpP
AlbcU3kFVF2c3kcIpH0mrj1pqCvjRLnseVuY9BQ+mQVebrCs1NShGkD7kU8rfkWE
lzp4nNrPWv16Lbl3o8/1lIArNWDjXo126vST5sojnn6Q4IbyectQ01NCJdQlZRSQ
1SGMHM4iZRGM0nbaf41pEsd4+6q7Nhv7KEltSxLQ0HlOAFuCxUQS/Okd0vTwf6AC
SEbukVdm1BXK/2J/aLY+XP3cprIuwbWKstPtsUu12GEI5HUYlKe2W0DnYDdRNaiE
ERqK/otT7gIleT3CWtfw8v2HZb4KXFiHGexZMTlDlllYEgWWgW0OrY5KjRdpYoq0
fmFWG1zHD5j8r/LaX1Xdla8smpUwpy9HXnpmyM0bqv+BNlb0wwyL7FBd4QKVkuiW
HatUXlpdmYWeTcYDRWgByz/kszLiwWMf+hJascGsnRUMCcKL6opaTJQIMjiaZsFW
0HApNprXsvrHbNMB97k1dJ9haCxJxqHOlW6kYzRn0TJXJyopvHI/BP7u/VGf2N7v
ZBpqEU75eGTaxTC+gkZWPWaCZ6bRYena6QDgywRm+8zPOOsHqZoRaMvKrKXM/Irx
nOALwYxcSueQo0XmZQx05j2oUSROtRtSVYf4ql4CTFv44kOSi4XOiltk6yk7peDC
NQeMB6MP2307JoZiT8dUkPA3jmywAnQyiEQfrK0ONzxpLBDFiIGHX+EWu8h6Bb1s
wUnJpaeMrMq1UMjdNhwzVmAoP0vKskbBATy1wMtX80odM2BT02lERra6NC9nHWyX
iLMtFugFOh6q1M7kNUbOIpKt5r4KlC3VcuOUIM9T1nFSh+IOs5g3+XP7ZRqwjXC5
zqQhIVOwwtHuARY5Bp2PVYwkaJkF3w0LRmRAkNPzCaQyraJRaw8TUgnNTuOqxppk
1WNPiktT88Ix+R6gVKZ1ZDNP8IR527Q7f2Bq3p0lQyPJ2hm6AE82dLebQy6XhMtw
jaQuvJ95EEZSufL3kx7X/5Lh8eYfytJJX3RxO3NzYQeK94yalO47vYKy63fQKijO
hdHToiK7XWJRkAeJx/cElXwit6rs/T0BgiYBRZNIqIKMnvFB63+CZYnt19sdRDJ4
BA6S2xyhmf4ugynL7IVVFPHo8Lv+rTQ/rrvgr1gblivtI+G9/eU9QmMrShUpy2vZ
uWxQIKl3FkUXUuq+RSA3hEqZEV6TxmrNPg6Dxe+JKJ8vIhwjLn1AFoJyx/SaWWeV
MVJTod+i1iueUwY2MIrdnnIFttPHmqWXTeFDkWCWABKHOYRL253La1z73u5ALqhv
TagigxLVnU5gNBJF5OZOPFBM5/mWyVsYF2vzqIEhnXhXzyQ926KU/ABDfOJ9I77Z
+pkSJJDXJgezPLtSY701ictrgMUtkaAC7RqX5YFczrJa68/1PWM8TyYrBJItrlKU
ngXWu7FUTr8hridwPrvKj4vtF57S6TOPomhoQp8Q65EptfUkHtHPDv4W+jublI8U
bdsuwEO+qJoZelpBVSmXi7GGsQpDDgLpALv2iBsTSgHKVjrD1/P2mfazAMmc217b
PkD2Dw70UgKsehX9dItOa9r8dKzYMHknJjJB7mSaRxYyUwATYUZ392MIsvM6nfDo
9e+2oFKdJZ3Ciob/htCUzqzKXcNrCKnr3YVJcdy6SuANXKETkC6BfXji6na5OUVz
+NjI0j4YS3O1aCxy6Q0ALj/1OdApCeLIkNMEGwV/wlR1p1r7dkYYcRZr4eewjuUh
VKGJzxB7i/6FqFpPct8DzugDYOBA8v/Prw9cFMtl8LJBA0oLWvP8IE0ekhpKeeJ4
j5WPdOCP7CnHQkGTaq+wnX265g22ZSH+t+9IVAfY9vBtP0XMPBcZbeh76pAPHKuy
e8AZ930kk0Kzv628/C6b9TOcdtJ4D3kMNhGTa3i74ZujUZO4cY+E7PK3ScDVHs3U
D80zsPaTpQzBGJl+gpdAX/Ko7FsKTm9BIQR5z5aUDExj3exuF3FPPGo7NV9faBFR
MqPoDmE/Qqm44mu8SVPj7SZcziqTBj6N6mKIyDra2LAXzYiXiLy2E6oep8EawNYe
8AplLfT3cc9JSgbex5agyyTJIHBhat+j6/0MEU+3Nx2TGa/CP7i02fJ2M7YqenHP
hn7L0h9VyvIySo5pHN4yyMQ2CPiQT9uzDPBRtGhoUT7Py/hcE9Q1kqBnrlR7tntX
dFIWin0ekN3n/t6jf8u+lUyjNv16dfQrUe9ReOa+zZ7KVBtr/E+ZDa7OKF0OwWIK
GMc6SDET/RG8ULaCW07xdOM+xriI7boGTx/qbR8QiQ8tFuLBWIphpcJbVI3JmSJj
E4p4668X87en7RgiTpCUDBAVBwOgzudtc1kbSP/aFDdeyEX2ieZHNYiKzz6svaaL
2LtqlFqGKWchiTENpucahw1wqvKzbeA6XVclr5h5QooGMC2Ae87lkkLTXU8gvm10
H1I4SI9GlvzILGTpduG251so8W1HUfIjePym0x2HoiU3uvWBNTJTL5rdElzuuPIX
Khguw1+/extr7bZ4+fDKnIayKAwZBMlmJjxotqH8NUVkzDM8AUP54xgTT9YcpEAx
EtjUlSvCHHhdQETl37EjrolXF+tATYl9pLnCxzZZovJ9qFoRH1dYNPmpiKq8AoQG
2REeQY3YHJLuepthlIRIjkpjuPMDm4mMn6khbCy/pHcIc4Dw3dI3GQFd9bnDd5FD
urp29g9CtqlzkDH8bNsQfZRNUTCMl5XD2afRWFyS2J2ep/Fo5v7wyfo11JQiPFkk
t5Y6rUPsPVBB3+WEBRlORwHuawfCbrpZzvU9+vtP77IAJbQNWyypeTTvZOhNTWup
TTfVdoD16mStYCKFkXqA2lhoUEF/09onUrbz/deeizhP6rANuEGp+5nHTJgAn4Xu
NyzXf5fYGFaFI5L8JP34pTq/1I0kW6bz0PZSMhfNxXfby8K3tExvoR5uvqI3D9/m
qwdQbI3I1xbQwGjIPSxRKbZc6lNCjB0gvjWJ9Eto/eJjhe+LCSsnC3QJyAUnWAtM
oo3S84lnlNNW0cdIh0PiDKXsvXudWAwpYM4L0rRcabeoYGLqOK1e/4VhOomQCmBr
J8Tcldg3W1Xov6cqw8Nf47nI2agTltKUSZHzcoRinmwEfS+JmArumKiRU6oKKsze
77uLtc1kkE/exneEr+PooyA0Bs7UZqbvZKn0lWr9da/4RAOzTuqQsnANsRZfDbR5
mCzfykQ5j0Sq6hzKmUXb50lgfQpBmfd1tF0s9CGX8QHuRaCMRt7sfC6qP2byHVtW
JHoV7Fbz4rxStjkoVWJkUhrZv1hpwogt9xhiHo3m/RpPqtW1nG6dqcusS/rgwLuY
UVXKfRCFcz1We18JIVIjTunpn21JZPxwinlOCSudsaPfu5KNP42ukNCvir+E2Bww
9K4ZSH3tTYNbGEctR4efsGXKMrmgWXrtiFqHZoNDKDL1cZUJOrnSSBpeKgDWnHIj
TpcSqjBmtwHWnjNdYOwHEpdAS1DO0O6yHUAlqM7WhZ/XwSru8LuWfprnAI1PIevL
UZ6SNEolfWFgZ1YMAueWLQDdiy/IDemp7MybuYUGH7CA3hQpklD3RIU2n41rTLBW
Zl96KTQMn3VTW7mGf3PBjmip1yHyM19CxXayl4JcwiWz5C4FkxIJnecveO4avrvM
hhZQvoG6cEO/RyjUvr7PvWvxgNoTPBjUqX9Fektj9XtY0OBJNIzct8zICf0duSVF
Iv8K1WBKxo3Pz9IxoPnM65i0Hh3pEchidPsKAO3mS+128bGCZ8fZcdniPoqMYP1o
7+ejQ7Fbnjy62mk4tufkqes7ZUUeWmGohO4kBa4920VCQhcsJlrQQV1X5h4vfYCc
kL9KmGYSEGJoJtYHi//T/ei/HWSQvmwVoojyl1H26M9eRAR5xBayQVIyIZF2LXu3
3YeciZtv+PpREodZs6aQPEqxuhh19w6lBQ07zE5JGBL4DTHg7o7Zcvbw5+PiMTYq
dL2PTuFBUXeWCFjDYM6/iA/q1eYMIst1bfLPHYy02d5BI7utxrYFqEICmGRaepBT
dh42FiFdFgIBD49fQjtgUExU6Dy3czdEO6b67WZA1gACQZk5eSq3R3Fbv2KrAWmR
HEETCzxXw/Ml8bGaDIbMsecKu9FyZzAQ/p0+L9zXdULBffnyWg+sPcruNDRaa6RM
6EtVouYEras2675pzdcQCPtcnT7gLPsidfnYS4dk7MWUOVId9u5v1I22FuF7Tvxx
2BTFRCI23dtEYtP3tudySHM1tAgQoUS95S0gkIGfy2bfdXx7OQvD3GUtwIqNCL98
ygP9+J+NRJx5PmfG5HY90TkFYG7FfYiVn4uJS0U6hTq7zyPwNU/1dS+Fm7+0iSMi
6myIKFCOlgv4aUhorpIS0ut6uwIUBF2DguiqwAWLbURCD9nIHCnF1KP/mktMpmmV
TzaQmthHdASB7g5QoBGfAuEEL8/MWFumjtPKPxi0+AvhE5QkS2ymlYsPQ6xyNwr9
fpFQaeq2l9S6qnqPeZy1Mg2GYohbiOclaRW9W56rijJ/rlhThHbVnY35AkUS7aKD
9iHFtBu+oHHpIBlb05vgcUJQbFg/SmOs46jufe7R1MJul0Bs/ww8DfFGlvH9V0O4
TTdGSEFIv9Xi2E+HUIX6HElLJmAp6P+66jgrVUttjM8v6x9FbMl4m8a8xm7/w21m
ZwX/Z/4Z69Ubfuy/8I8xk0cG9UctfYRmjW1Zh7ClZKb+/MoYGixRy0joPtlwpmcS
QmOsYOb0pZsLXDf+5c44nMAbOw+p4FplvfO6ZqLDrvrva88ZMAG5ImBs0jw0owYB
8mM3StB9Eqw1j1GGaNmEemuTxbBc7fyUdoH3k+HWkPplpKq7Sa5e1TEPk+jXdX8H
I5x0hGSQjJ1/+7ccc73+liTOs/fECM+kAQYVANwYncUuBlKJ6lGB5bKqfe9E15Qf
5izWQgcgqRFtfHtLByebA2Z8i72MDsun1nWq8wkjEi+nhrpJKRP1CuYTZLuUU/ug
WR8OsBhpY6vFXsa3xVC31pi35sM4UowXx0t7TZ5nWwfDk0NrPnT56GuIq6V6N/To
YkxqIEuU4Gzj4w+R9j9tWWIuJ7nS+zwHcqTldrYVk6IvGofzXZS0l2vLm/SYs08P
spfFW4pO//KoB1R0LjeKlJsIT45BwT6be3ZgCJWdCnWQGAkie1/71igV5xRdTSb6
vLVVp/CYyqFi0+ABzKF0CIQ7slbM1FvAsBoc2g/GETF8OiclOQmTaqSF9Up71+zO
wyyBAbve3SDj+WwvQzIWUm6vRkCVFAtpZjGj1ydWe2VuP6SB00qPCOJZSz1fH5v3
m3p0gRcNfTdZ7yHhoS6PlJJuFdsjqpUQaRQRiezQ4Uxk2nws1X5wcfeV2bQwlxc8
SWGv69Ii9EcQSDJ9fsBxlo/LXJitgq0WzAf7o9GXneEhFt4/7BW9oQkgL71vybOT
vMy4fk+F/8Tv+T5iWK/hrueH3x+Rt8XAWvFliEqana3wg8FFhdGnw9kuzyDT7KiE
QMe9lhZPAq6oiurxFnTkjJmapRp9eu1OZKJ+/SqZt53el5H1kymF8RBlLEODAqpC
d2+CCxGPPM1Y/K85fnSGeyp+tE+mwove2+kjDlNKE+ry0SE8FvhqWUJjetA3FDpC
eWqguXqVkCZvWSd37KsvmSloLG/lzwyQMMEZb0i1qMfGfygM33b0W1e7ql5RaBne
i4VE12Tbuyag8nDTX3oNZBsR9LV3ky+Ix80sGSpX/12fjA9/aCD5B0XjdUV4WdC8
MPXu4/CRFnuPQr4NEyREaCNpWN7YzdcMCosGGUO/GVTrqEnWBpGmei4lM0wcgIu+
q+5vdioxCQS1K04GP+dQ8OjYGgZ9jU3l6uzFcow+KixnYlV4C9JnUQGOlpD9/iCo
L9Ym2du2X8eE+3eZ9l0LHM/yb6ljjXlA71SoWrnE2CWJJXq+Y17diuoD6XA8JEyD
XwaLxKJGNFlVLxN9tKqa/ei0FuQQD1VNJ03/k+RnaLHXkoHymXHF5yc0qCba/PSa
l0ZWsujaHYwQf0Umby7RnqLoZ20F0NZguJVauBksm9Iix8IQ/MOcKxdWCLur6QII
L+kxoXJcyrJNa1jyMK6xPLmK0+1NFv/g7S24Uhpo9PhD53QtaM7m7RR5X/3d5bkq
g5u9Xpnuorlg8es+8e9HUah0nZ1gGL53ZXVZ5OTV7TCOf6WnGE+K4xGBdw7LzyPc
DFepZVPuwXT9h8+mt9IRb+2Duq81DSGD4rmwy9R/sunKh0eyOPo+dhDTmaImYcw6
`protect END_PROTECTED
