`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rePZlQ+YHAG57T8l9O4/5yNZmV/2GYDgQOJtCTPHZbn+zvolctTV25yJARWVa0Q+
K0aRyfg9sjXAhg9aHRtU2Bv8YCGMLXnVgE04AWpA2XGhl7BfIBdZJfJEVoJiL/DY
zeORuzJxDBYBQ1GvqeKyEIsxvJBoDGqFRC+MkT1Uw1TsxytNeiuInmf675z1+Ycz
3XrZOC8gb37xzM4yw14+uzkQzsY1tzGYR9QuawT+GEztNusDJXTrQwVJyGSEckw9
Xzc5xyWe87xOxRecCB+9HHLFzi8XPfM00j1F/UZI0DuKd5XKHjJjzi1Dd8rsMd85
607UKIHxk7U9ByECpCGdwKRHwYRA9Vc4fqrOO4gbAyudqzprOfRbvhEUXjC8LPmq
meojG5UEZPYIvmIXJMf6yVJV79HC/+z6q9Fj8FUqAW00HWsRfRkTOahJKwBVOHy5
toi7tLZmaPT8Yt+kCbBn149nmFr4FKEQFLe0YV4fvSOAXweGCSCRSNWVoRc61Sru
52+pzxHx862S+rpiD9Mpyq1Dlsxgmb3wGbp+A1hGbsdonXA77+o8qfdjf/uyMrvO
IQl9IkMh9xvz5ZzaTW9J7XO2CsIRw0KAEW9EBbZuKV01Jq8VgKYXHRrcaVVDo462
2w7rQsLpMUCFnsLh4KS2aUjRjogq39CcMqiO1/c3oW6U9wfQ0yOuVNO+B1mPN/Qr
foilm9Vg8XKw3BD9aEIWfPmPiB/txLwf7hebEqH//hZhFll23n/Q8IgvKhSHIuvQ
gAG7mteZb0HYc3TlrkzoNxPpZ//27wXAnQuzApXFf4SrnGLxLdgC9+Ebb596kKrh
9isTUwlx7SKGJFYJenX99q48bHDFb5nvI4W5Knky89qmpR5FBQvHrqCY8LS99G/m
dkVqjoLfe+xLz8R0C7KeAzyn1gCzwqGXOOZWndBzkp50K4o0Rpr/BXVjcIli8ZyI
kGW1BffcMkwh6HTobe2Gfg0C5EfISDZKxcVoa/0TViy69Jet+FIvK8YlI3yAReYX
2jun98X6GgwXlls4t1AXJsGtzGbs3wEezHg8867ADYmkTNPkQnnuGu5K5CMwEbHO
2NotNltK6rfx7aOkUAdNqVHuLqs+9viOiz+Yu6SbbhHLAyK4gqJxxJJznRdCciUW
kJuvJI8FOty+XX7TFP3TojPzTO7dD+qHo0ZRFFePqzNERfnw91KP1mPaBaOaSj1G
ySG2x6CoV0n8kOM7lSs2NzrcCsxx7Qtii6c0G0thscplpwhm0HzlHg6kMW1nI0dx
7c0nu5KRTnIS6hsBkoeeUfkrspVZCMzgEtIlru0HBVn8MBcKXOudR+seECM1srWO
HprX4cd3PpRWlaIbrzSfi/LCOsqEfjmyU1+r8uxCL6TUoWyQr/gLco/tVjAfuyZk
d2gpM28zS/87o5nVqSaz8D4jk91QM3FUQ5iu/rY/p+PnsNTeVjUPPgmp8O4oNl0S
hDS3AX9PpAMcMrFuIE0a9a881qV3+DkRCgi9tnhmSh3TohuyWrH9JZYoSsBI491F
J4xbIIvN3xdLV1yWUxTt+sAppZ26UDGmSuxMwxRfPYxQ8sJc5ueyHjZRT4TkR//F
cjGeSjW92T2jkATbIVsIG9S+TG4qv8X2zwLGVZk4K5A7bTheyN72md+IvouhLipP
yKlePcSbrl5OcFZVb+u8DhNJze5Bd3w/Yh/D5IbXdyh6A2EuZQSc2imD6dq5CL1/
99b+/Zj1EOW1o4MjehTg5tkOaIP5kRsQp5OMGjAQa7Z32rWdfF3KqAmZXY43ksuu
Z8HhmEz8rO/OnKXG54DWDYWzmGwA4iWSVHsGjfJRksBvi1KrxnLpfqwRyTaNibIc
eHJhu6555AUIg0Nx3QwiuW8aq2oRyPpztOhTSntRPVdk8DqYy9i/3DIcgaLNm9/y
qWrPCMTTYEH2VIROduu1Otd4K3K9V7J0E746uHnN2TbOJEaTvYcO0Z2inKCurzUw
iq2x5SaLs4HuR4ccwfHG/RKUDVo25NjmxjoMrQzmm+cijGk55zYYa8TQRUvxGWBN
1IgKpdmz/KZlK9HtcAwpzX11/MWouEaqJ+GZBciPEGQ7ulQJAuIELuLXKMNI2jo3
bucyN1jW2HbkYQmduhDl3/OA+78l6lkin8Ns83+u1UFavCZhMCPnjY9fX/y+5OkV
viq3AkXMxHUI06/GRgzxQWhyKJsFcFGSiUeswc3H5AeipHlgnX13u9w1/WT9zuIH
jC4bgkSItnwXwb2HHxtmaraJzABGW6ffqwi7AZJ/H6nGCrphygPQTId+cm2TcZbr
CJj6LjGaDLlBNhVepaN7pVLvnp25HC/YZDjhm4lpDOlNjDYLFRZUw9I2VYT8xUlh
xFPseJlvUg1w1X49QVJkMGsTkykKld3iyVEMD2SVYQ2BEZFek1RtHRbAR/55L84U
pQ3SkVXnAlQKHoC+ifD5fsJR28rEZKOmjkeXLWV3QXchw//hqO5MWMmecZIxU1gX
7mKz0G8yOxAUOJxPJwGGJO+VDWPLLzwG6hd/IpZjG0j7Z59xZixPdn45xFU1YjtN
/k68lMboa3gUL/p0k1eeDM13Ombt6wSyH/ChIIFtCBQ/JzH/OUUZURUU+7IATH9A
hDZGlAocKuYf/FxGVTwvUvP86f1E/Jy+x+XtcSEh5DiGpa3kWSeMcexMf2fkbtgT
QVmPYg1vCll5j3lQuRvNLU8WBP78YDyTRdLgfYQZS8FiGIdQHMg/YVN9Lr4plpAW
z6HZ58KBAKYt2xFg67Q63r0sw3i9ea1WaK0cwumYXjjvZDChl+O/iyab/F5O6T0p
Xc376CBmSlgH6ZweTKZ9+g84u64ptqXZRchHa1F4+IJUKBiuJL460owZ2V9IV4CI
1MoZKKocappSM14xLvJQ48epiepLI33vMykwN68r6Qo65w/CAiedLu0hOYNKbG+Y
8S5QSNR38haGByajPmOswtTc9cycT1v5yWMXFwsotjrGko1/UbOxmmnMCCtxvlHY
PRU8QXrPoglb137dyyeeCsTY+28vP484S2bzM2nzSgXmbwOaYdtjEwgKkQc9SD6u
Z4585lFbGXCCFCLYSB31r7CQB5subE9HbzTwzLhwqUlIM3MvN8ab9hccEMBZRnbz
g2AN6B43E7WVc/0lBa3GjSti9Da0fsDRc1Tp2ppR8CnhNaQfKkI1XpNxb5TerCXJ
u5ZyXjj/FlH58RRTuE0e4LRV8Uvv6mcSfgDk14VT8EXhMdJh14ZbyerWgV2C+Rup
sa88OpgFXcXVyfCbeT6AxQGpsJcnvWB4NceBz1pDfPa0mZviPevtcA97gAXbkzgu
8HNgAm+kM1ThTAsCJPD6VGrlGIyQ0uzB5PhvOYjTYDzQciRZBe1C9/ab7NgdjQqx
PTvzB3uCRVF3CEF6IZ2TiQTnC2y3HjvPp1Rtv/y78vNxfu6E4bu0Z+0kpv4dY62l
aa16IrA83E6kj+jUBVrebhkYNfRGLFu6iNIUaTaC4PxOIuuBFxQkQdAgBEkvEJvZ
fW7HkWXSgerBLP16xmOx1wBhhZpLh0x0P4MK2BhUnJkC8Tnq0TsAJZL0uQ1/D7px
Kj5idjy5JM10lCTfBI4gkK6LnAnwqM3GtgpNTYhf8NcdZzJ4n9dLaGa4AqKF+LOX
Tchd8ryQqFzvM8l94h4GCCqMGcMUuvE69z19Ipy1cpUKE8XlDEiXn3kaZVHjTUzJ
zJZ1G+Rr2CrKBAWWZouOu4w3UBu7TNpaxF5N9BuLXK1Tj8BYWXXCNlbSGPcdqnBc
LwmlWD0Vs/pT4ZUO8TscdhdpDpSRIOGoy0T+VJ5S2uD3t4f0KTUxCLNxNhyOzCfv
QfZ1tV1ZlPa1JnQI7dMiBY5RP3dXYf9dS3NhPGxlK7VpDF+MHgpyCoMKtnhcFzS3
G+KBjY+5qD5TwVSts50s2+EF0TMyoCB3ZIetVTCUMOGGri9Yd6vljz+M/S84Iqvs
tRDIjwtWnI66fXe+9zZgdJeRuGvSRyMUBjgo6LN2C1x/cpBLq77VDVhUTupCszP1
RvL864e1Ej2Z7yafgijsaG/6cDUntb6KB1PK1bg4Na9TRIgvGdqv/hLhW5MLlSpO
QTiV0rWjjaOZXRfyW17YKbTGjFVMzivS3y+Fb6SsnwZsOSo5Wum4F5usEqHmZqKA
VdWxLEXd3uteMvGI9H1jElIIeOZvoYJewHgy5sI/hXD4N4uUiZ6sP19LKw+t6/rj
3LoEMGWy5XsIXg6+LYLm3EUfVZyLqtE6vH764trIRGYMYa+dol8zAGPSUvJIfUWP
PEobVt0Wsmd8VPdFQ9xBpB5B9DZ07HfUOr+JCepUv+ZSRFYyGhnJ4f/jloyRGYwH
dWj3OGmLBN0lPN3vy0nXI6/zP/4Na6ddvQAuRsM82ZigaLN+U1+yQ5wLTlHdtXrq
v/5E7xxa57UGOT/r40qbSsjTNwxZlroBjaIqmz+2DLivtCAYZvK4tTGnq5WQqNw9
iXuOaWo6BeW1XzCGbm05MjYjS6ZGAmlgqrPPDMgwYWmILYahHXXelWefOsxOjXOm
e/W1kKjFWa+OZo7eEznpRVv43K7ap9fZ6YDTD2XXs50yeU98jqQ01yOUOwgciLIj
1Q8Hp4cSvCKWLDAbXWEhYKe6mxu+eiaQvwtTWOWI0MxRk32Oct2XdF9BpLrLZCfw
+s0dhQw+YqcRdd5/hDae9TxTvAqH55E38k4nZ8cCMV9FGscfiEIJMYwMAg7ilW2W
kRAJqHgi328W5eqRHqPf00EMHDzx79Zs93QE0ADlyyemMYQwvXMr3qNs08q1Opel
55gInF0wa3Q0BEJeNviuJdYOAhd+kxsr15kFAbM28D+Lajfz3ZxQ9iyhIndd9WBF
9Z/njw2rWipbFjS//LAWEIoDz6cwH3zOZ1Z3fVYjjMNm84StgHNf1CtmY532mwIX
POtVORRvD5PvFdWZn93WCDDbFZCy4vZonISBXHhk4KfN8zi1W6J9YOt6N+i+MR87
YRW9o2edR58fzBy30rHlKS6jpTiINY00a45Z4QJ9GkXRrKu5txT7KFnGeflpc2Z9
tiVlsgwgCMDwGiFmLDDZ/dGgmVzCNklNTSLqDKt0cz1HXiSjvINQcB85FsJw+r4A
S6ltHllYpiEZeKgupDkm5JYqq9A77NA8IGidY+exT6BeivnPWuxh41hjtZ4E1rOT
MVjqv5nZuODq3BQimwuN/ca4yfF3VRcG9jGUunk95Zyve3LoALBsvVRce83OfP0t
pHYkIKMsHosvvqnCzBNINInSTkam+30uN1y2aeg/o+NdNDUGlaIzNWsJJ0WNdMk7
EW2/yX25Yegvs8HMD3PkhV7v6l2tZANlVsOLiI7XP12tVx0X6SLNVE371Fj31mPo
DyHl1eIf4Yn74hsb4J1nHrd+4dhNo/570UBB5dOcr79sb7kqJAefHC1C8Brn7KNl
Ak4wbzp1dU/S6267HaBBq+M/tcuGzGe9jZdD4CGhQIBrC343zhanh8xCVrg/K73j
XhXyRZx6WlcygR7eNkNQVrHExIsnsG8C65TnCs+zY3deUe67mv6BtO6FqEH1lAbw
SlQOr91RN4eGJ8oA+Okmw1HwSmiIv7vetNQDJP6HOjxeMOU90gBqFkysK4oM5IDU
QYj6XypmK2E6vgRWbsYLmw+9TvrPns59GD1vckFmDdvvt+cfE1pp0EMwtWIeVdYk
jGRZEfVeGOxVB2Q9u7DfKCjNLHb4pvYRApMtQRasR2Od31w5rwJhwHdBp9Ov/Uvn
XnmVHiuISWB0oPswhB/HNobbJ3jxkhJvutGxSRY8rR3NRUvAkT1Kk2RuFWYiyPhh
/Jvoi22PbzZIxiprit6f3qCy3y0tOkWwq4EVjdntVS153RwQUN6Jnu1Aum+E1ojL
gWnLSImaW7WCd1RebP4lz7IqejsbN4p+LSvdOYozYpDTtcHw7iGdpmY6icfhlb+L
Kgk6/QqUVoeqf1V3sz5ZPzmURLK/kqkG8svgOflb6xfk19VEjdnI2XJA0bE2qpZV
jdHnVVgUeafj1P1QtvyCKio8CkS0ka/qMHhBTs0/q96cGnRFaTsXNpckmnVmKja0
b3QdiouXQbQyV9DhW5WrRqJIoQGoB1nO5WFPvFrq4lR0xIQuk0cQcpWm3Xm6zrZG
SxJkfStOrTxPXPs0ZaG760AbUA7Jbqk/WxrvtrtTOExfdfxtHvrUyU/pAx3olu+Z
SBPxS//V9N/oeEPRv3I1coszFBhXodmqPQiwIB9TCVv7/y75fKvTBY1b+v1RlEYR
TAIMZX3ZjkqukUpgCjkT8nrv11pykuZwvI3EIKIqjn+OwNINWNiw2u1V8tuNGc1l
l1h/Yj9c64GYE4D58TFuK95ZJrjRVgPk+Ic1bhZgdHOwXkGRdYS7BOSsuiLwjRsD
j+K+l6GCXjcctCHAFWBvvzgL9SA9B2TDTcGD21lA2pWtZojkpVyg0eIOA16VbsQj
A7wDuTYfd5Os0dg24mxN8ndtnyiX2h3PCgbgFLLBbKEOaCiOLsUDLUqlYHnw0V+E
BMCh7REQ3s4+dy2nM/PVIXb2gQxt2eqPOWb5eDLiRe2aLP+6hvGlfZHlC+fG09Hb
hFlTxTjdakNjsbZBxQIkCZRwXgCD5jVNO3W7x6IEqdarmPyqqLBoSxVsCwbaf15s
jmhtIHuEQroFGX0VZT5Bm1KVpz4xfAFKbeSBy5SYhyTHwwhObbERolHUsnrGHdli
gJ2op+puxdc4B0m6I2ZOyebzOwGeixixY9pr40tIXAe7C3zjoid+JaL8d+xnngKS
DfdsL/+TQwiFQt5LmWjKPlNVyKwyC8go2Qqr7Br7/DPENs1fsFDh2xlvUVHNsLgi
kZYiAlZ3dwrcuyKLCmLs4SrVbwWTn92TK0Gac1Di4WWIPQ/fzTM23A0o4Ft5HVjG
5+zbHHFGgN0j3LY24Os3yToT/KZnHsLoLfa99102W/kbsDd5ZsGLASq4HFc6it6x
jh7M6XpILhHwD9lI8sn7fgGw51nVSbc1P2NspKM3GTn266UL3SnbSAHosmVGN6G0
eKLOQLenhLyjPccGnaBeCOAXJ8vogQCQpJ17DaHHr12JiqDHrOQwExCv8ROr9BEc
23jJjjg3YPqsoC8cY54Pol85u/EVAdKfkdAqbVMsa6KPj6P40j/dCofqJUJBvntW
BKluRpaxDc2dQ/X7t3k5nRSzk66qDxSECr11IdIrFBsn7B5diN2O7Wxo7zkog+cj
3qFvdfZEIx8BJcT86pT7Zg1n2cVkwbyU2UbEquom4ySdU0LA6S4OEzCuNE9oheDE
2nO8BnLvEuAGNww8YkS7fc+MsqAW0X7pwM4lvsiTiPykQ8dlT/PKA0TpUPIhVtR9
PZa83WeaLiaOfYEtqSkcza752UajsGzUcB/7bm+kkLOkEUPSB5XFpPd0txSB3p6o
0ILRd8hdZWMwGd+tYu9FzeFyyjaJxpPzzHc9qMgaIpU7l5r1D/uF5t6pB76dXyXL
LCzn8wl6eId45vqPtVwn4/o+IEG+t9GUbZiLKrEkhqLQOkWS5XMJiCLURxOFDxWr
GqekiNigXY57QdDpUXzNroniGgekTnM88v9MkrSHaD/+w4m+6Qv8eScmHD6kt0yK
4tsBSC4TLqi49wtMuNMFO5OJajp1BZGrdyElsizHJ1Zm9ubqG8o1aUZKd744V0O2
kdxEfEIdYAJnWx/EeAvgzDWzM6IzYBEU51gVhiePbVbL4LHchalwzU0Yl7lFbqMu
un4KEkJt3mV23Fg9hsHkNLLAKHs2IqYbnQ4CPEMtATV4kqD0iHSgPXvAykihlSkO
uDYnaBwC/IdbhAcE0AoQA6YVB9mUmZOJzBgvRthypDOkrRQ7NaSgXiwM1BIFxBLM
XbJqjIkGCVMcqJm6vZXzzxWj+Zo+Mc1ehOZFsHu9+jjlR3mXCUUV4xuf889H/7Js
nGXIdLEq4McNJsJQ5UNTLs6hSaEyj0qJeZ3YhH6+7JoR/WXFLOrMM3G4oQ949ePq
p2z0iL29c7TVBJ52orWn6WliJo8exCdsZUWOHEARPpVbuylQJ2NI1cuG1nCK9H6g
o7eY3ZoAkVYEOw5kZhUVpH3rNBR4b6nojEHETjyNRkLF8rj2GNMfARAUEK4/OF9h
4ZCPZUMeUYUk5tlgcAE+/RKwo1ue8bcMnlQoM9uPA70+5JxkC/zXUyROi7sl9fTa
+9wfIDLzXREYMKzAI/V+QDX+akoyhKdk6YAuy4V0Ux2p8GwmZSn53N+YmG+M/Oje
sDbxMJHZRVgkIEEyKuLWopNx0h2c2UWiWtTAgZmisvqk/EB7rA8onx0f6PC5QU+h
vAIS7kdtzy41NyKvstYMxxa0fgCfp/q8UjkEKbvNK1iDhURaZ9yeA/bJ3UN/k8yv
mnwROynrcglyKJO432wu/vBsuW0BUf4hnQZPUL+Nso89Kl8cquUQHhNkLn9Jb1dq
vhaOaApGLPJr/EOoqd6+9e+XA+vmK/C0s2+o6X6KhNhwWnZV8VYJRKGGky8c9Kq4
XqdRRE2cESur8VCQv0DI+TPIX0h7INsejzZ5KGke+XPm1Mfz8CIj/3dZ1YFI7J2e
SxFmPT/u2V4XrrdcLLoemspGm1vnyqIz1l4Dt9eGGycLfiPQ5+ZRm0CJT1DWVutR
Ay0AcNwwRmQrOOGpqaxe0EDh3tDdY/goOnl9KXB4c1wUjuGPPQUMMGlBK1Y6FgM6
R8FH9YkbpAJu7wimf79fdPnDNZ5iAMP/cLD6GbY5Wz/rQe/Oj6N5ootvIg0WDElW
v4Xjyr607/OFI6/zF6bTiyq4bj4X5fbac6Wvp3rDDvVeASGcG/UPaZIE8hr0dLDl
RSmJCr0pQZ2iRp2EUm168FlJir20eP2th4fC17J2Fu7deFxo6Q8modEfTmIqgdmA
AbDEmcUeja8jEfFPvVfRle8E5hq81X4siu21/M7S9XJgiGNQnpd/nFyHFjmnIor6
jbnFnbaxcDH0xyHkIbTEC317bJ8JjjC/8HMx5qmAlHh9asOOnkDGuqi+v//HF1qK
MzfxA6sszXF4nWHvt72DUhB2RW9yZHUrL6syAvMM51g0oujVyCdv2Wl9H0EP8OQB
ZHoGmPrCwg7zXkPWvzUHdvJqIG6wBYITi551Dr+9AGp2SiceAUwjCrUuEE+gjcHD
lWgxv0sjqempKM501or56RXK6P9DMZE0CMJHhg6qo4dq6R3H8zW5w6i7FI+JCCdL
eoW9E7yA0Y4rNhMupcmOr3pH/d4pnThRVOTcKOih2UyQNIqV/eSPacwRN3i+x3UU
e+jvohaZIURna7KZb+jJnrx43bKH16NKAS9CqAOFG9i3cgX8VIH9SvCU1vEqWBk2
9laV/tgvq3w8UJzl7YKmwKPgWpvlpWSNYje8jVPi0/XiNEyN5TBBE4+3UqfOTi5E
Z/ixpekkYN5kxK2fq6SEoxV2D5lVU5HSTnBnaYH9u5UtpbOypprDP6nYyp1cUYkU
iDoxvMoq//5QSYEAwCAd4c+8WaFLigPMoICJf+j48NqzZEVRTcsV1AndDNJan9lq
ts9iVNUtGIeCG7QrfNQGEUyBoVjYMC4cZQxIEZekVygI1NbV7c6bdrBBuBYhtIlp
4RySDXE9LCabsXyZm71ImzmiYlIcLdwEvIoTsRAYprwOop0aSVh39lIw5nqZ67da
o7clPbGhhgx+fpPBQidtdikHFqWc6FogR8Ew5gL4ZhkHhirjnKfKoUckjVnJeL5e
B8+5nIvafiDyim05/d953PqFkl6SC086HFYMbwNqJ0nxPRCrTXzSkTsoYBv97Zyz
R3SM5M8TXvgc42H+dZlBMq4xZMrnUcTBFof22eOey0DCOdL7kXFNPHqvXR4CFnp9
Lr64TpTzDRFC5DFS3RD3+yI4FdQdwjnf9dalSBwG602YZ9eN0+H9grdbU406crY5
crUDyG5Hy0NJ36ugDqH4C5TisrEaxJiCYLD/iti+1nUZsl2Mw5VoUWyp85fqqnk6
AKZx8SuNqXu+ug84TtZ7XpJSRuLKylrrp8i1Zip8+YhWHpotN63R4WySDvkM28IZ
co8vijxiIRcInJPPUqSgcqjFyENjCBo7AW6StOnd5NO13ClMbcpjLLCme4TtxV7x
pDM/dspfVGGDmH8Z5rgmMiQtP5AEq80+xAiUhU+qDw5fMpaKYHshSaRlDjM0bXhN
tNuxwGT/m6mUJm0Fu6bd+FiEqfneeDhWpqc10ZWrPpyVQtgsnOLu40NVaDwiYddQ
E2BplARaM7EfSZOxvZez1PDmW3CDde1nyBt+51S3Jwuh6sesS5082K3S/5tSsOec
fjmBOA2P4SGkV9kHP+0Fr7wvxpT9uKhcwHLwzoH+MKGByZ1PBhxYn+QvSZolMveZ
9Q5Nx1xUmS158gtEiytBF3IZEiuo9d6VwUZ97rJ+cGn2CLz2pqja3pJMEeGYJb4M
wONthVuP5y+Ui1PRbww3To7Bi83/KNXPQOKq1iuD00lgfUN2sSMyDYM3PNEm9uaH
O/NcwxZXD00r/o0O5xowxslun8Hmfrmtb2UV/ajgIQ3MahBDrh+RzaZPV+NcOJzj
zbIS2HVt4TjUE00+GeRAvTGXiGoNTN/u5aXhJMjprKoakz5B/CQswurm2NYRysmo
X0gznD/vUhKL1gQ/3KJacZAdXXXV6rl/oZZXX+7v6xb53AFsm1R5I7EczIAKK5tp
VCQGGxWAQS3pa0Xw6BBIEOJw5EUa7aLtnY09dcc9TPZbFsK06avZ52H4TfgWgIzz
4ug5mpBRFFXmavCMmQIV8Z5fcugvZDgxV/v9n3tBdcRCfAIxNYiWF/TMONiUNJI/
NrQ+yDAruuHT5vHz3yZDQfnmUOzP4Vl4qNh5xipMCgGNjBTqGNTmhK+9AGBWAPVa
CaPKbUyIoyunClO5g46SdfbT/zomtcb0jaKoPSdsZaNH9WHHtqslbE7drVVh6shT
97TAj/NbtECghZkkLcIMSGGE8QdVwwb2SW6wd/UrK3cTgFeuPPcwrtA+YT18pAu2
imFIhOhGouBodUsB8j4XsqVjwR+Hnr8XGZq3X7vyefwnzXW5X6hKJhnZuwiM6EnS
65f8nGYt65g5i75dt9u/dbrpL2nnLmOhtHxPJU7i4uNMqq7QvC8Y/XB7YthUAlng
fBV952cd1k5E/3cAar8ZidnSP4D8i8GQi5X79uhm6146DnnJL4xkw6zY1s5R+RA0
OluF78lXq4hScmX3troyPwkLQL5xedIKYFP15RXBhLgvNYtV2eotRbhGHgY15Q4M
D9MBhf9otCz0D9s/HpLhbkQ2pS0J9PnE35xWGLjhE0P876ITptWkQuZDvi7e4Twr
bzBiV8iPY63Q4L6edmODp0r1O/WvKf/Sijm45whh5zQkVOy38TGFVPQ96dKH3Nwp
vuajXsPDiVhAtyzmSoWFMp6rTOrEi+mz1P2eVpl8y7ZyddbySeZtFsYQ8hwdSS8g
eNlxLUnL1FxaeAKp6uwpHmPkX0CbKU7d4X7dISZdPQ8rYfFqDFKLbycs15J4JcS8
7s61UOQ2XX/UASe0DPRLe+RUSpV0bDHfcRoBfw+SHI0VJaNLiVVoIuBB1cJRiCEY
hf38P2HXiAs1x2hWJ44KYS5vBBmQegdktjh/b+gG12qIbmzXdffSiuNUCwXMHFSn
bH51UnvpnR/D+ZfZ9XEACAkF1InPWIC+/NqH4IqMZmZknzzvdrEZAxstTTp7TX8j
xs0uof3QqEMYN12Ra9CleA69EDoL5+KgeCC0G5aDfTtu7pHNLtRgZqmMx59/sOTe
lT7xJB27uCm2FaEyzCuZGs0+HM8UBRQFnYxjp2x0bnf0/+f/YUAlDrj/zKlHQx91
KXCg3Lcq3Sewppv6G++EBxnEOzO3X1vz8earvZ86iHFSXKR7//0xO095ERLTG1z6
exyAEYcpfbwvcKss6xuUwJlqrE1Hk6ezfI0xKnPLi+wLNxGCqWoGJnCTHMO8gQ8Z
o8oZV3O7IZlz0ko8WpE6V7+2ghIgLzkjzu/k5KKNdSgTH4CWj9VBDk7Ot08vbsEP
JO0lCBUJw5y2WyFqp5EHzs1hcLOan1J9ceQRP5bInzDpEqMlccxh4xQCoM7ua1vf
qjMTTuM0Jau9va0clfdA3YQ92uY+nOYFXp0CnZDT1qHPqySvom70vN5B+zXZG41C
uMZjDJq923lRxIyGA1/oomn+ZxL5GvdVgqXfb3jjJQTurPsuByWSipOngQT2eff8
dKQxCD6HksOoWZizPs1AeOehTed2KU9XIE3XcvxHr4TQI97PBOyYqrtvXeDQ/zAU
J1S3VLf22bs8TFpJAbLEmHE8KIQsgkRXOb/N8FXhrD2INH9Vjgxm0lzzaO5xcH8p
yYHl7NL/XEW3guFRBN9EdQhNBCio0Wge1ocT4W9W0IoBMBNBbPNNHw6YSzyqQnPh
bL360EkLoO+WVmfGuics+rlLcgkrElEw6JpNjpwwqlOFKmpis3yAdmWSFsE5JSOt
w0KZkTPaGFxQ8yqgViUn+rVDpFToRXa42h/Op82iBbmeWNX1hK/Jertm/5SnNWrJ
z1vNH0D7jsuavTwJuiOZxVXo3YM/0ziGT3npNkNQSDYWTLYfrpEtzn4qdcnp2wNs
HlAw56udBD+QtMUcHC9VlP9v2sprDx52+e9QpSuKZFpL8GFaIMEbimz2Y/9rR/M0
RGlAJZ8wPUCN4LN7bAXsB+QdMCNVeU/fk+r5FfqesWmHqno9vNbmLWdGVBqYEXCA
48WfGscXl4xVm4W0yfFFpNjm2CUq6gSFHzIoELe2VnlAX0dIsq32/QHWp00roZEk
GHSuEqzg/cLP4NYvXCWwyWCg7EVKfWTa41Ld0MMd++fuUedhthDLajZKRzkM3t9O
NR5qXhGcbNbMfrkwALp1ZQJ9f2IBwrf/4S2rlC1A/jdxh2SFBGDKI4CnZRXps9qI
EFi95XI5H8nsSmPinNoXo70zNSu/I9i6ytTmm4oZdq4c2T0wcB2TtbXbxlYexQYo
FIXYtypLZKkvlV9uAp7BPGMSooIhEsolMC8UGpRLBCxd980imTrmOeA250DPwVDi
X6TJOc35cbD9IM6QgKdSuesg401TbKSlDeN7P/5iCXLFZG0Pxaux2ZPtWeAOMLTi
2uA5ifEW3OZVF7IoZdqDOKZzlUrILUgEwiFkaWx56+1pwT8VDhVUU9GwzrlA+zzt
obQqaA1DQM+ttzk3IBXvFIcRuHwpcrlqrDlKudo2txGGcPkgNSI3S6d8TKirVfeE
EGrC/Ri/d8HVwYMSssl+ikIyCCHiEvuEvlSi2SQJ+N/Pq9m0mQZHovRlyyltyiRR
et27G2TZrMwRLqIgsan8TiA4/8ZU+Rh+OB1nGw7HPRBK0tInvKV85P/kc5olliMU
P7yWn0OYjQJrdorxQSs0rXzY1cmOyfGA/QArGx4IG7tPgozIqOZehLddC01KBTvB
/T2mB4WT78ws+wUS1aI8u56mWdPY1KOevX4C7XtO9HloqcuOqMNPdDGaFHQaVkeI
IciR5yaNQC+WxIGh/obKIUDZDM4/oP5hstXmtMCfi1OuGPGDdynkwd5UjoVNM5Pd
t3UOhvQoBdSXthIv6TYCjburZeYP7dDQzqO9uyaQt0rHDmb3S0+NTJrLXVyuSC9P
T0FJXMpU9vCcM4P4WkbLo5IQO6wd+7x/ZRvOTndFkOVIZeKHD5kGwWsUPfRe1gwa
8DAsZlduYPV5uQY0T9sPKXTXjiCVofnGUwIHibk3lqcRKVYMcxG52bgZjTijSjZ4
5hxWYvMClzWBQNAM4YTg46FDQiRVDtU5N2SCYU6LULNd3w/IgHUo4WP/Fj4pALXO
ZOyrGi4rA54LaQhuZMqXhc1ZL4stdcM6T6w1DPyaXzDpWJMnvML476/YataGAtRL
UGbWX4fwvZewBMxQbtEj6A4YSWNPmcqHzKzpy5+PmsaynqXpjtyms9O//GTBWBoe
mt+bsTIdAzbyby1qX1Zj50Hu+Gdd37xFfSCnfBgCMvA8LjdDISGz+Y5aFOCP8AOt
TkzSK8I7BFym+5ZEJREEPVYzJY0Z02ZXHn+c4xzI9AbuIS1ZViOF7ihCDdyaUvZa
KPSs15XYg9mhz0Ef5A1nD/BRMPf2FDCQSF1vRebI9sljjGP6nfoEwHDatylHtjqs
O3xtPwpVofeKB1m7Gdc4TwIjunV9pnADfrKTzhNZ9EJHzwWzdvJW4S0pZYWLhXe7
yIhUCdZGuUQG+3mms7juXJs5mTq5YenHx1B9Z/SdqRJ4sWMRcacDRGw+Q0aUILpT
FI17AceIlYuVM4zQ8zE8KjUeuwmNHqTK3bM68ZY2K1cCMctH7yK1Vzf3o7Hma0Y5
7tH03FowHKiKpry+yy+G32RFkG57/oHbZr4jTOdY4yf9+KhF5ZSqH8NqI7Yiip0H
T03Cj8w2S+1rc4weRFHJodz8/9fTH3+5LF15I/ij3Ivoz5HKyjOtmdB6W+fWu24s
PDjgEw0q4FtvZYESyOQjeK8JHvzV2yhnzv037f4gi3abS5nfdpEBtB6L1QlCx/5Z
exw5YuRpaqfqbaiHZ0dPyw==
`protect END_PROTECTED
