`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D05y3A2s6GTE5nQ1Lk1qnL8vgRBjFrrxSRYDZjC+P3+dSqJx3/6ZVKerVN9ZOPgZ
HNF1zDnbbuqZQVxjKNUS5laHC9io0hxA2BIVez67UP1syunysm7+W+Q7Mov4bMJP
xUIClaVnCeN1VddnmFvhwmMn1OcEZuYvk04C6wjozzXtOP6yK1tPI/84eL5iRzKX
WsrOzkVs5pjWoB76ogfto+Ak9ggzlab0/2SEfRBQieAekTNZtPW0j1BF06PBdF5B
MhUBitS/5xo4fkGYegKwD0YCBwP1S5kTOxl1hEBRq7+1mRlzNOKtFWMHmeY7RK0/
JhKOgGJlZCGj7I6kxHLPBxUzEkBeoc42uN2Kg89qkd2XjdQrUekli0YDs2C3ATbv
5kDMiLmyWZd2PJPQwhFTO/mNTDy5R5RUU7VAFkVwXRv6wAfKGfe0k5jVZBvP8D1K
RKgm8rbr2mb6hbiWKwQ3/Bjjjk4mpEYLpQrpfZ3Y8L9s/TKYU0EosCgPDhoOVau7
u33tMwd5meZBNjTSaZlwu4ozFDK5u4J2LFBQvXLkF8zW9x7925shOml9n3Ni2Sfu
0OpIITGyqx3ODYKx3sML2FPLCdnFlPgZdy/94pmr9mXH9FXesZc43dC2JCxWG44M
lW5UpYz5EbnsKUxFcdidX7VeLWlhgSiiFfSP3g8nDRw9iyRP5mN1i9svGVbpp0P/
GGZ4tK5EyYw355eU1n2oiNX0htgLN7Wjq2E4euMF31nS4NP1fKA1wDIesitD3hkc
YHolpAi4n6D6u0CZmiWrGwhP8QLOGnCapkYRqtP29b8JApc0T25bp7uupOI13MdX
kJixVH6VzOtfViA6OSq2qmHDy8HWQNC9RYu0suaUoOidFS6DgOiuajqKmMcgaS3x
bQoGFkiqMfcGOvV5X8dMWpU+m6GzU5dg5o9NTeyLPmJPk1BnUEyyEr2zVR9ASxeQ
CaHwW4yGQWOQOV5wXGFjkfEswvUDDcr9/x+GTAKdSuub9f6Uz+N8OFe909f7bF+B
aMrI6lOz9vABXcBC87L+eNRAQICLxM3nd9SLfwTD/PMQCVqdep4bMl5oJ7mtIvoX
xKWSH1/NOdoy8WuEtwJ0os7bM/aCHD4ixHCDgWKHNU9z6Mo8DA/ySveyQMQUYfHr
oOfbpUSpQrnYl5FoKRDuxdGl2asasDbUCPX2uYQ0w7LVLGEglNxVKJNPoJOzHVd+
XnWRGa2cnnNEXzNEnsbKWpI0x8ZC6T8dps3YFiRoAPlk0ojTHPTedEu2+esRNI+M
5SQZIuIF7pZYcBVme3JFI1HNLhqmQi25YoTR/N/uNJ9kOUkhuYB/wxcVWolX6R06
00RRXSfV5lIlwORvmv4l5pZ/67OT7Qd/LXd5mDGhjVt/J7+i14G+BjDBxTlVtAU0
e741qnW+aT+2tXt07FTlyajvVJUr61eP2LTPesCnHTNeKOf4nMgert1/kUL4uzyt
qmlyUS8g+yoMIY1KgLWr7LKdLvW1j5tTYufiBBzmZt2xs4UvgeE5TNN2i8y7Mzwf
zFZ1+ER1xzJsD5Rf/oxLbVA6Cxmyc+CY08S5doMLKSqIjCdIkF29Z6lMJPU/Zdcw
EzNUvB6yAF50OP9mIr97IS/eiiqz9VOHV+JEplUjoOzH++O94eJMqt80ZYSE79Bg
6zrgWwHyGGA2KdWPvbgqDDekKI3EVngmMdg9Ci134I/lKL31ieV02dL10KNeddaS
LAwj3FxPhBlWOGSbGEUS0Q==
`protect END_PROTECTED
