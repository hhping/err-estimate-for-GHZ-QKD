`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VWKcFBJthlPS8DB+y0+MS1RoMnBfKhT5qQxGwA87POOCqdlvSbb8ji7PKgvtVqu
tFJVYh4q2BPjUeCOgSMTlYU/do25zOejw4aCM7KNsA5/4rNnVnwIHBJ96cKVd8o/
P8xZ0qlX9KSudi650Vyo6uFD++hmbIOHXXKpXRAai0lUxYgzlejH9N/5KDPgz8Hj
ji+jf/NRffZoCh8I8M5DfYmF/IlPdiuydTKdLexLZH/Hza/7fCye37qvYy9NJOj/
5WttctlMy5AO4EiwCN5phxwt007ikLCttMAyEP3aHIsJ6o7qGL4mrfeiTrcNdajc
sdBl8sfqqb9V9iEFWWMBrc4Bln79awk5dkcCTUJlYPGqvhCp+KwqHlel4w8BItNv
Rz/2S+DBll0mGzo6EiHeAUl1Dxl3kS6OTzjD9hZyxAgRK53QAQZNQ/QXa8QmSRgc
ohmLT3PLSoOpLswkymQhKURmCjIZqJ+sE7K/7c5UUUK8YYDjlAfjtyEyeJtHYchj
MZRCy6a/A0wVYM3U9fgzu5JWH5r3dFZg43b0OiO/vbyWA6jJbEJSBJJbfih/g378
3DQ8rJ4tGUPb/QJj4uOMXj6dU/ddVPUjK4q6LcI2oZtz6Khh8gTEuySpp8OHIlAD
4nEpBgU8RvOXmuJ3IlZDix8slxWuX6yOp3OeneeeLmDvxfi9dK1U9q1oqqJ5bDnq
2myp0dq063ZaNP4nV0ob193WnRO+OKzhFf1cJQaIzI74hknoCN/oqwMsIsSvmMls
O2sbq3wlpCtTjtyjAM8VMH5Y4a5SEhfTWXpjTjQpx7+UQxFJgPRv2yVr5zPsCimk
FpWHNpo1LhKfCpnorgcic1lBLJQV3I5abk+phooKwcJLG22NQqwS9b7EdelVP1BV
GIi1L0YhQV3aalP/Fpdm9SAS0Jp263IR1cSAq7cPWDPp0Kzw8aQxYQFhG92+VLtb
X87q9WubJvkomBpkSf5TkZpn7m/mt0oHeI6HnG5JwsPMcGFl1/9H5EGnqwYhQujv
dN6aA3yvg4L+P8U7meRudUJy0WmaAL8KDC89pxorDPHSJQ4bMT6LsAAF8gDoLQ+C
cKC1CUNmenZ4kMFCPq37+uymv15AeNe6QIbYEQffewXlCS5XIAodizL+FLqFUj2o
VacxkVHNVgW4CRTfClZ6oywPkE/4HPp64CTM6EsYOK4yhKnTJqN39wg4xopNW4Ea
eRfFY27z+A5W55HUUCoRNQ==
`protect END_PROTECTED
