`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7r7gvFwHzt5ZtmclioU9+1LAcBIRdEA10geZlFuuBYrY96LrsdMkibv8e2bty9k
uHQ+V7kGGeiGr3yew5pFFL5QjvWmo39oIGNmcS3xvw9/F1Juxc5cpuxbPgNZlIgG
sYBJhnqq5EW1SnmcZ2OaEBZR5JtHr3fFNx7+k4tfGXRVP8jM/dktNdzmxJsRnZ9S
jFy8YPKlOrqGMd/wQtYPlHZ3QHCU8bAWyYHhWccQu22nG7OEJAE4Ji6y5jBTusy6
Z1s7I9sbRRNTnwVUlKQNwJh/gytHXx+fmByQOA1Hj3zy2QcMQi/uHbeQrbPd69fY
8JG8KGNEYJ3hb0qWx6HVz/6p/Y+l9RvtrC5ztBp8sqMkFATIs54i6QUh6p8y1Hvm
3gxFyMxwoWYRt5j08EoeEaaId6iln+KzOpThOQ8JBu0jqclAfK+2rlC5ZBmf+wsb
nlGL/9jPKqsg7BTyeuvBQ+8OuQpN1/VH/B4Q7YptcRlUd4JKgOKMaSmc2S3Wm14v
sITWRFA4JhVvr4f4Vf5fjd26fq+phoJ/IvXnuinxbRgAYPQ9aTfV5BxI2GG2aN03
DVKNxoB1BwCtHNRnQfg8qMvqmspwzGIyodRF6+6AxV7fA7BP0sTnx8L336WVLKEu
Ou1D+T/XPDnB1+iENrUIj1VThDKCg+m5ANTuTejIXVM=
`protect END_PROTECTED
