`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YD1GPvNSl8wpKZRtTdRNxPcj2gNl7kfAxlfWY8N6XEpTwdTumo/n4wWzodif3j4E
rLiS0X9e2AhqWlfWP7bbUnh1BvOU3bEO0Wo3N3HpsBn/bpg89UFfYRv/Xt5Ro+vS
1XcedlEzkax9004OKIoOFLrnd1gE2IZ8SHCAs1qGVZW6IWjGkE+V3SyF+76SZuKX
QqCrooMbQvTJXgBecLK8yrBuF3HwlmbnJZSY2vULdF1j/LlvjNGpNKICQPqOhxo4
UweaFJLC26iQ3XeIwCpSyEn/CcIdNooB4dim8NHDVrKWxL7W4yyY3LgnqdTBrGde
PQC/4XoNQ69oyPevn5bYsYZGwwq/IQ04SAC+jg360iq3wSiuPR0CNIiZQJnwbSjx
15ZTF43A0ftF+oOnxrCQutcpkFnGdpZ3rpq5lqmYV8QUWrz61BphDZRD6m4pMU4Y
br9la4f5OwBICBpFhoUJqeFal6ipn1fPX+1ArRHsGSG0qqZjKor+fTYmfot9MKFT
tVXPp0W1QqPwzYXXANYKolyMEw3PDkeuuOOicsDou3YTGvkt+0j2DhRWpNDGm1ki
A4azII6eP/edBjYVI6oBJvezom0dgN5TAMVqjJgIBFeOlcPj3ez9UaUugQsfus7K
mGA3Tv6+FC0ssQn/c+QtzwIPOmU7wqHBElEsSVZAJpUDjfA8i3PUgpUAyP+cSCvd
zwN9qL7skqUtQKVzQ0EFjU83TkCdxYnN/AB+UoF4v4ebeCiD1dpIt1QK8sOlBUhp
58eWfsJjlCinlYbRwwYQ5znMpqaHu9rUeO8pVy+lx+ArEhKaiG8sUfT1AW7rRbVL
PxZ8IgJ8Lo0S1DqD7r0eHFEOAcbnjegOTU85qQoliKZdLNeyGqI+KRH/VtCe6YbT
Gb3D+WbGtiY35ceDT6IXi1XAfNdsndDnUbt7FqlGZAl2I5MyfAkRHgPrA2fCf9bR
zAHR7aQ+PYi70pQJ7+ryfY/W4VUqWzRlkP1rYdSTu7Y=
`protect END_PROTECTED
