`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjgSJVErSXKjCC98rtonKcElsr3KU1Yf6CXAph46zhOV+UpXG2KsgPesCnsR456z
qJF8QlhPKrnoEZR9ltJMrMakIm3t/wytzq0deGYrm/6Bd9rJNCduC7Y677N2rr5C
h8iHhyvz4J82wpsUfassVB47/gnVr5EcwWPmvi03zm86XXqwjXUcBIwh6fRY9OCy
ikGhZxKjFIAqv30TvoCwWdgj/sAh+w6cpHOVQ+TfIGPHwbwdZRxKFcM+6/QJgUq9
uE0yFjiU9qeVcjHGmhXpcFfNctoGl2M2rEuTqY2PrEyX1pbhteVhOs9hY8vBBc+8
tELYmtVk4oEtl/sVk2q55t2gmIACBp8Wh7QBfosPKJrkEF4tfd2EwKqNiFSc2Qc9
WnUXP8cokIcPM9//7NlgdyTFlAq0b8o2yGp90eL+s5cILMvXHSTqufNguzS45mBh
pmTiT7PFw6etvlJimYcfeGEIlbbHorx4yi+0vHWl9ayX9Dd4y+CjgcDljK9Jay34
HaiOtxWrbW8v+8ETpZuGAuQs62lSfGSbELmHjKG1ZTyYyV8Ep7FzL7yxwMjjcPYZ
AhBge1gcYk4EYfw7B3SqrJmN+ILtOWpWVOTGco598AprE9Zj0dF7I9H2rnD+9pIb
bbakcOdFONqE2ZF5sHLb+mfYJBqQkt7j4+tAb8sXM6Q9ZtZh6H480APGcUPOSCYB
CJNHLmanHWcm6mo0bG3CvqZBhKGi5eZb+CuA0mMG2okx/WF66la33P2tlSeB293r
rF4SaPvrqYOhOKuvRn0p++Y4c9CA6OpbzzZRmTZmeYGebzwzlXnrnNWyEyIeVsvt
QdmPpPrDbkx0c/bmQN8Oy8XV7oj1UqLlysfuM9tb1SAd2TqMitxP5AGQ5gD8chr1
vbMMkbo5f8omdEMwO3DMfDh/dAITP7gwOdi6hrJQc+1wiRPNXII+xCO3m2ydt+Ux
WN93PkFtmgr2RtQXUSuDekIJ9nIG+HSDRdU0GGhVcxPlf7yBmUvkAc3poYaa/WaB
8IK9m1HjDbnkljZvGeaQAVI7/eIaSVQ4xBfJHwFJSBZbWtnSXMW+OImm8eECCm/b
++FuaQIIgv0VdlSVJXPGbLRx1wnSmzXxN5hVYuZW7frzvbdpbtmemEGgwq+G/ukU
LW1h2Phq8mcZqawDNCNP8zBUf+16/Z05ZLwEBYW8RHE+ddezqHnjHoatFn/a+QKD
2TLzjOlmpU0N/8+y3HjEFEwwUTkE/8eaUBkEQtQY3HooLGtob332WZVE+HRHcvnq
GUiumxr/GVb4Qm3DGgtcBeT0fYZy9o/KsTGa2/IvXpSIXB6CU14T9RhPKFiJ7sH4
9Cnb94VJgBghMM76tm5e5T9HMcll2kzEaNhzGu+4GG279rcLUnfVNIC9PdhDC41i
H+7MCxFDXLsDi2q5QhfrJYoSZAo33+H8KQv5nn75wi7oXfo2LOOMwN63c19Zz80F
hUVf7jTaWYCqZn08VCdCO6Ev8VOBzo8r+pBfEDFru/8RKFWs5yQINJEw2THth82E
Sm/HQGtprzZYpKtoDI3NumBWFWw5RkuTW9xMhE5bWzYiLeEXz1kPPclT7lbryFCT
VL8yAgBd9i49O83ipYEixcyBIC7wB10YymxYRoLXj1YmxdSvfe5J6Ra1b6tRTkQB
LT0KIrAXQyulM+Zbl/kCPVqfnlxQbbcA8zyJ+c/AAwo6gPH+7FNg66e6e3QiM55k
3gB/QBkVjlAWsT6/3G5tZLWLbZwVMLnaUq2eHG6/dfI/jKqlSBRq/JPv+g46k6iF
N3OYxs7L/fGxH87Ld3kkpWLnzwFPvLeo+cf0RTLJoz1GZz8J9nklQ1kzetOKetya
WpEfdv6DM2ZHgZezf3RrieEGgg5xOnfRrRFP44HEWIbKMgIdrg1e7qhMuFnZ019z
iOD+jMk6woNrcsdAPGD62AHMCQByf9Na28kbiOkNo21QQJwb6iNzR7HkpPaLBURi
SsxdjLvTNK1lynWdOUbQwHB8cPxIZWSc0cgbqEgIE2Xs3k5dyvqlTqCkCfRFhfrq
U23kSGvC9hdnR074R2lIzPSf9gpX9MvAhVPhaZ+ysosZd/jjufA/c6klxAsJ6oU0
2AbIziQteIdaSOfV3taZvw1SzMGn/Qsn7i+jSOK9RBqY9lj2nklHs970E1e3qciq
C4ZWOo9EEFdMIHdVvU9lmfrJ+qeTnFSNmfz+IPM+VfFDbvNVjSRTdc48RXfOL4s/
ydtGJl7CR/O3AJAdTRynZMzFWtizaxkMRNOqBiZnNG2AOvwmBypODpbNucZNrqFI
KZNAXp+9OkFewhwKL6FRDLcGYx4543N2p2+/D3UXB4ihT+TJzYWfqokc9M/z+Haw
qPeL+B3yOK53u++eBEH7EOC7uinQbyAk5oC3kDkvCQ4yDGZ1yyeDxRSQTVdgxm8R
Mxf+/4oIA2bjmlokAlf1YEM/0ZCndGCGddFQ91JMBj+GEKr+Ns+w/3vLSk6zCVjz
4kXt/0E1EqwPhZ5wMyspjqb/1d4jn35DplDV0j5FUkbUSFSAB5b0hI9pHteqBy6c
Rbfz1F6quzP4YlFB57RL8PT07neqqangPGLzaYwra2Yc4O+CHCMBZ2n9uG7vhIm7
+sSWuS24VMwhF0UyfHHFhzsubUeBgE0hRLcrhlRp1yxlAG2KS/orqIHV36Vh8hfA
XurbYXB7GfwiAs85RkVOuVy+GiQXPWgvt/yvzSqLJpzMfrymtH87yZcQ/v+A6O15
m438Xd2mquDJpmMbKBVIo7qmm/j8C5BNeYsz++FMt0MWgJI12TQR04UIpJuNfT12
Vvcanv17U9pYvzOR9cO0tF3nKoTpSczdym0aQVti2ZwtrUbtF5P7IcgwztpqS7H0
UuhE2SBA1CdEB3uTx9wRFEKICJyyvsZJryM5aAuHwQPuNpYM5LpIN//k1Q19xDQm
V3+1JftWbd1eAQ8Qr04R8jFqgB6zbw2vuUgQhSlNCDcRpv7gwOcScr6PDx9avfon
sJPVxaYLr/VjhiR0UOEHJu6kuqq7pCUyHcinj8COFRiCzv/8CNtIUFBsxYYU0Cvw
yXT6IywkL6/oLlRKQnL11/+MEOVvTmTtKL6FDjoc/4uHC7Oml73pFB+OAf6a47QU
SDjeimVzNl19IcgNHBzk5Y21ba9hQYbcS/r3/2kgrsYLI+50SQFkmDhmhVUKYKpi
ojRKDNFy3n8lOmeI5+tOip21Uh0wzLYG6f5dbhnBWKNBAsU7MAwBPSoCqRagF/pS
GpXUKxtXZqiIX1fo+EANYE2/2oRUxWDpo5ukAkwppkzjykx6SMEPw3ixBlPdhJsf
KmYJ40BPicYTx0ta2RBWaHjcSMycJ49T+0Xs+2dfTrgEPVmZWpplBbzy/5RI4OCo
f26eGnMflx/I3v+DdOKPiPHJld366zgTpYUfPwuIcSzG/XzCfnAZzgkHnbxDdJFA
XTlMNKlMhx1HQQGKl1CCzP6a1yzyaMu2yZa3uFyjMmMtHAbjhb1QKnx1yEYrwvRD
Oq1I9l+6liPQWnoz30NmYhaMQZm20z3z+J+QUL1x1GTgLjFSiQsOn4dYlyyfh8yc
0sCanfKVWkvbQBGbTQcrHcJWxP7ugb7zd4/ZV3CxtMAb5nGMMxHnId5BK+GSrxTn
+kb4r2VLUM2mL/vbmjxuJAJcADmFPa+03uOUW8xwslG5G50mYQxNynAO6zoW+LzF
O8A6RZy9VsCvTshzHawE/w==
`protect END_PROTECTED
