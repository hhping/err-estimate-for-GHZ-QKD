`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ozlw2RiCCLGIPpQmX9q/PzVeiLkh/2DzExydg8bxC6E1zp6h6Zds62LUOGvU89v
J/ijl/S2l+o35rbDS+PGUxz2LAEgMEDXcjID8T2du0umiUUm/ss1uB7SE+L3ekAm
yi5To0pjnj8KxXlCVVA4BNO1I7y01ZNdVUKpe5ZHCBopK20kPDSXz9eYG6pExlqo
0pmQVIyq5LdtM3zRdWpSeIbLJeV6dRXlR69nMniH47ZSD2ZNcrJsh3KofDHSO298
nfMrxoa9Cd1UBIp9kAQwotPZ0lF+eA33wCFad9Rr8ivJ0ChZgBYejXi7Fu+PIayQ
5ucPXwd2fMUw8QGOylFI7aaq2SZ2ra8Sf7NBSX49f7AJ9F4KWLN4ULhpmMi7XZKg
hLcfH00faNoZNQzPUybIJNROJLyhdsHYS7qf96n3CFww0bxccpYubfOren51wRUl
NiMNATD++RekAY4l0q3tfJEFTym0jMIG2x3kWDcn9S4bD58HSO5X/3+e7Zp77gtb
SylVEuF3hozMpL+wz53E3SOdlkiIHxKVOa61fHTTp/M=
`protect END_PROTECTED
