`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQEPZVlRL1gRVhsSYXACs2fqWE3WWMy2EJuxlOPd2ZEgnp0x20CzaViwkQA5bX9u
FB1FUnSchF8Q2dx5Q2Tsl4j0i+cOTA0UCMMyrhOYHwv+zoY1+3LQ0BBGJvKRlVAi
dgw3qlG1sPs5JJHpbALkG8dpcxMnISsJeO8Q9SbEao+1UTwdYiEPq+ISFp6vzAOh
gQCwHOj/mQ8vPmza4JA39DCk1gtNVmTHcas6XkfFBcMOSKyPuXcrb/vU9acCxPCd
6Kfp9cdGvGFsko+n/zzYT0u+FD3x3mDFwWzDqxATdwPxBK976Fipw7eVoCrw1jlP
z7qoYBwygdW6+goS0YwJjXZf7OefeH5yxVLgy0l9eCk=
`protect END_PROTECTED
