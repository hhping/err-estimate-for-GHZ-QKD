`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CoWV2dVhi8k07Qasvma55qntvY4yO14iKyz3fuhKrgBK69QHfs58zVFCHbgp8Y6S
Dq+tANPRxzGzaoB0NhN1dgfGWEUJfwulI6tbo6595qcmtjqhV9nXQ5A3EXgBDNXW
RL5C4/w7/i8j+Ly6/fWol9vec2/XrrScSyQF8wE1d5+pLtPxStBRvFGtvc8/FTDy
bKecXzscvzeoYNhZRhnILxFfxM2/8Hkdt3uAxEm5EGv5ZQN5XelR8xm7T8Mr73VI
JfDfYn/rkEsxM+9XRpnNKjlyVEO/y5x91egAXPH6dav/TU3eu4/2L73X1+0Psjb0
euCulkNFn5t1OvDAOQsbit/n5lB9fl2POSKZ0VBlmJP8DFrmTzeqwH3Ysoa3yoAD
ZXjkoTbQHSq9LkeoxbyqerfDvZq6tV0A7lNBytARODqASbI603+kPaHrYnIcL8uy
569dhM4Hf7rOWRPtYmmmUYfwbb/bsZZ52w/WUc6TS+6OgOHjhqsqeOAtpWgYfbOw
9rUwQkDpeCjBTvDO7GrVejaIQr/ZfQgDhvJa+sTOevfWgJclxZm4JLb8/t1TgZ+B
c+k3NZrSvr5t/TurRzuWrm5Orfx1aRqpEJJlNetE45EFHnLzKkTTdSpVbD4ToRKE
yjAP+c7fAypZbZWFsOY3hABB4Q+KkZPNvOrCqhWimF/PSqaXw38q/gXTmc9+CBWs
09XaIjHUk1KTcTs5bFH1Rwv7kRznFvD2Vz8bcRih3O5zUsd442N/v5KbSx8ylmP7
BtTeVSdI0dH+fvzpuFotobfI3YK4S+GmYzAjY4l8eIJNYWb0rcoDgIYepnk3yCEm
x4zU+31MJvS5lxmceCKWntSfWjiz+Aa6809hFlAHo+Y0m777m+v8HedhzB+PIVjx
p+c0v5HA30u2XMB3HDDv4M/o1TSHeti6t1zzazp3QU4W8G51or4sF/NvJodsfU2x
IxVgsBlsQdUxD2gjDzH7udzmASAaldo6tudXuo3OkIXe6QhWWWV21rCwRqTW0xhC
uUMhTsaWnq+PS0eeIPoTiiTOR0CsXI7uuExsonEdtQaTrogQl6LXX89ztPt73rBZ
D+CntmhDye8rBnnh4iDstXAQtzRaL20xBMxebPyfFXnwwxGeilPs/pFqXxYAcynW
08yfPY8BYo4cQfcWzno4t5atbJm9BpURWMRdn26T4pD+t9+ghd+38yuJ2Nlyw5mf
yqc9kmkAh2OyxdcAJuF2Xugso5YoZeL9Gbip9XE3F+uQsoLznwenl4cIh1YKvPG0
WvTGiQdJr0s4KkmvEGL5ktmMqb1/kylxrn97vD+OqRsUbpJXHiG940MFOB+cE64h
5qc+rFxWggU9ou7P47nOoYdFgLEXA3EXa06HJUiRzm3O5JEklLjjgfQxvIuUyHcb
in6Ba8ARm02d7L3zE3R26oJeXAsMxEHkx3JLX03Vnp9Jic5IOMi9hzogOKsRdv7y
ah/XGohBBd4iWL+E6wrTA8XomnMcwLTpOmT12xAMvgusjTnEGXHofB39J+bsWbJq
pVSbl0nAmXc0mz+nGywhxUADhpREOpdn4GJXMLNbEnKf0ct82/Joj3/NdqKRBvk9
wv4AKjLUM/GkFudQyjuFBLKt1/An4lAedKTGMJveePUnwBk2Uvh52nldHvuGxvmE
hLKJGg+CjZp4HmWqjIzBqUUYqD+G3ZXCWHT834zOzF42lA0c5LxH1udCJx4qZHE1
nH0ORdizjIbP7ct08hGXMbOQ5FZv4wrjAcqLo9uyE9mjo5EvBLi+M1WCuL78ZucO
aNDwtZFmYuhZKPQNkQo4Up3yTkbJqZVA4wDF67tJf3xvt3wbiImgVpKkMEqIuClp
QFftpCYeRXOy35h6sc5th6xaqnkrpCd/PYKAYXoxuJMLOvq/SR4QDtVtVhYbVU9t
Lm9hIdZbywK6yrLR5kAKkm4vf8sIMrZPgzCAzBbsQUHEE3Wm+b2/nyu/7abPiOAR
1fTbhPqJSX2CIhOv5qOVJBqwGL0Ncdm3XbyJPqTWNwaYair82X/RFJAD7TgmFK03
PrYkp24OZq31Diroho40lL0mgfoJlVAnna52LLtixGEwNHTy1bFiQwaRFg9yyVZ0
7MYDuduOcldLKboGCFN7OB5vFw4tBOOIgI89GjHW4W2MvgVgaZ7exTjbQEaUsC/W
n+2/Kdiz2iTqAF7oxttWQW4a8Tcak9ivP+Gxw/ozcJ+UMuNQFiz6eX4J7hXLfoiH
I99H2C7rCPc9e0pU3kLKHAYPkeDuKTwNX6JJ9dx1fzppYFVvQs9kT4abr3YdiRz+
sxRR2m5TWO7+JD3lAKwYbOng55k/yAtxXPOqs0w01apC82s17lIWD8E2WaXm0hk4
fxLk0zjR0RKLAPhlcGzSPdczDqld9nFoVhEvJq/A+I9FleSUiFO8c0B7Rtl/dENT
JkRd+dK94IE28Tmae3BfWK3cCtFeD8hHkOjoDZEcqw4Sa9WrAeQ9A2w12H/a1LhX
coJu0OQu8cYwieaN2thh2A/VO16A7JcvX2Y6ylA9l7qsMFX01lMIdfN2xAwl3CAR
`protect END_PROTECTED
