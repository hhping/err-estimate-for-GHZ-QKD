`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBDmblQYUOsvN2Bq0bK2CjkuEb6P9Zp5bJHWJvvifH10K2OEHzfVAovNpx+pGp+9
cWsELrPtImaJknf/meyqCybnpsRIwwclGwUJalnDUI0x5VwyRML4nA4NAxEskAHr
8cYVpLy0WvT4oU007syVvU9Pp+FT5TfpBnW8i5w6+KKrmslXJZotXhfuGPuj8dn+
F22kAWmdh6Cf04weI6ujmmUFNNdXsGJFh6cMveFUTAWa8gFEzj99CkPMnVwRRiR9
Vlm1yqL/NHMD7EXUT+wI/7lB14ONG/Aa0AJaZYNMudz89wN9Lq/zSUHFzKQOkaOe
j705t5CkhRO/+Yn++8VqWx4bGGEtJOO4RVpDuH9Tt4onj6iVS+3CQH9HqE4SuUHQ
72rqRXodfir62LgFTXgnQdvAV14kHaDZEVW5qSe9t9uvhTH8TIypzxJOQ2AP4j3F
rErpHNmMkmIMlX3rMu4/AtUh/LIpAlr4hvIyzN9OZps/w2SI0zpGyS0w+vj4qZpi
6wHsxRtY0yPaoeXNlibYM/Ucfc8HySPxSWmizy4xNBqlaH4kJWreNTz4igaw+GbA
Raq/dAnhNDyqFN7H4qt4HWcFzo0fh358LAW4OWWcYednb0TXVizLGVFCP1b16f0g
vc99UNi+Y/PPA/4vXwLKxvDS6hoigCPZCXev+O/KcF3hGkBGNBv8gcsjj8obz6p8
1a3f3j05aYjW9aRqu3bpfWuJ7rkpjOJWbt0prv5PyrZ7p7XfjXzEppKq/BvKksj0
f54rEX+GYLJVAoPP6ufElsen/RsTAgaPNOM7Yvv82zV9kYsk1p1C3vAuzNRQBPuO
EkjflxSd76h1XLmJizvn0Y51NVNCvcgdx9P5SKiG9WQ8ZoEzAbGQoXGJ0thodNqI
dXpRgIbQ2GE4XiQ6yrMZ8rfqzuPFpNiRiy7E1Zc5qsSwXDLGJCOZDzdU7oMzKhLp
+JfkMq08loS1Lkxu71hL2nAWa127K1pQbdN4YqWaOT+2aAHi98iIF8nP2TOVpr/a
sPs8coEGvBSoT7HysDuZoGd+kVK32NdfNP/ph2cgEtxhj3h5AwyYaJlSFfQcODY1
TSDsMyMBN+acXQTflVZfPIF6yntlwIZX8dwPv0OGr8Ow5f9Ynw6UrEIlBHtauhFi
DOqhDWQwkr6mYSp9TA/9nHjpOLVWJZJAL5PAWG7nGTiy0Rzn6qZ6P2JgjaAQU8yg
WvAefg+5/mKVJCJ7XRAysK9JmaO4LDZBB5FgNt96F1PkMpHfeXeZmj5R6ug5uyeA
9rrweWEVqpik69ZzL2MA7ZVSho3umgf/ZjFNeRNiVSIFqrBxL6AbfsymLi7wNVrv
7ySY5GiW+Hc3BKVN3j/KARYvWA+qozONjjKUcMEkkGVEr+qVfgTDPcOdznGDdfdg
80/SnA0gLcmNVNhXXoR9Zh/N3NZHSPeNKc6RgoVX/IYgTVNrKbtkM2P/n6pfVO0P
4NwfPcJX+g3K6QenP9ieFkcZH/mCQTcBow76DkcPQoc5t2Et3B2OTgJM8UKQRcKO
X33XAqUxW/OIeuyCWvMRDa/f/6Akl00tmB30ujNODouAfO8O+5VbgnjFMTf3HXv0
/4RItMpC4BvXW6YO5HdE7z7x7H0IOIvQ0T0UzNDJcy3GiPnCD2vDXxyyTudAnmmb
OVDCWTV3HxSRdpfkETOTMCi1r+8J1DLLgJcPw2ryb8SPEhRRGcK0XV+i8+BLVJlY
JvYXGwKMRprLo5ugbBtgJ/rdmyjCWz88CTETV3244hipvNZye4rDSf7f8yFTrz5f
Qi30ENHzxm58xG8IOAmsBdpBi4adKNkv/dCP8jcrVLZ+6ABnJxW1IxA7gNAKLKzB
UEOnkyQmQOCyR1UA9JUwV8cwX1/NI8igu0goEtupVqSebMNRAfoieaVUdVMxMaZo
aH3iq6tIMIMOoWwhoffyBLIJMeVKb5a5QdWHsYly8S0Y5FoI2mEj1Jkdul95z0tE
fLyYhMA9uIGfDXfwx/OG4uRpeJ9Z3n4uW9I3gjb9vi11i/3zCZZFBH4LYf2NmGyz
m/2m85201Q3T6AHNwyaRFiY2oMdRIigx8F4gSTWvogWtYTPKMR1mgxjvZ008yXwz
XiJQAZYSX7wlsgc4ckxyO+lhgvjo3slYsjaeN9IP07grcKBdiyl+wcw0N9VRgQxL
rL1KQtS/CfwUS9Qe1FxhRrZ2Jw8CIQEIuEMjYxqPX20wlwZijyaJdtRE8uE5Qwln
7n1g+utcZBqt1WkJWKsDN3BdrrwY0kbjp1LJu8/GYts8q8Vfeb5VHAOk/od9rY/f
yWPP9h9IQIZ0/iKBDw+YGsbEwTkzFO2O6sQdE1dBEA+/mrC8NWSHVjTdhMX6yewY
scaIOHEUfh9H5Q2VN5F8IKGBK7hGaUmXbDOM+jqd2qMGSru04tjwEsDOc5KWX6Ce
S5lnzw+KjRKbTaxnkxcdo4CVQvvR60hDO21SWUQ79G/HBwaFURhFzXgEy4C0Sk7N
BBULsf/G+G4dfJoVMGjvhqbHa4uVkWRP6DWA/xsOkMFSeMah7GtJ/rFrd8Dql2OE
aXUqHzgNZGdPOyYDvJwr0TBwsHsrHFU5nz8yc78+HBqUXwyNJ7mOajg7aMV6tfQG
L6BAiifxo4/88SdB1uJt6UUB6ltzEdOt6+FkZaFxts16D6WzymXy3TxWB9+uZeh2
cCEJkeKRj7V+YGHOm8twUaZKRYXVhBqxBGKtPY0fO6cycVvpzHylbK84oCM3QNUl
8rXpzxCXKCW1rdFa6LtbBEllo7xrQC+NkzwK1YgZmFYLwuqIyDcWrUYHqXMEPHTL
MnyFsda2wv9ceTlLRp9lMTvwQxc00c1Ov4wMR56bcUc+opQJftKap/9nyF2wzvJ2
0AnLjCe+BGZ1EIDMtPduM13o6+Ub+DsL+jvzzCIl+HFeMiaGgzUw3tMp75+d4wcw
PocK4T5htFExxs+FrE0sfxJvOJT8UmuI1ii88GLWm0tKvcgMb8dRLpW0at+AT0eG
pN9aN5tcvmCrmfk30alVFBGbRMRJXnzAMQJsqRILdJ3GeHWTy0elkrMZXjPSPcNx
RtRJ+nDUYxJ1R35NIuqwdpMpm1EV4MHGIWBA83nr1d3YF+P28YzDnHvJXMEEQQeJ
cfp/yXD92FXxcSt8OV1Igjfr6BptLUDosF3zbkKCCgbEwLHXo141i4rVr3G3SyWj
ik7Apx92PlW4+kZyDySM/8eJkK86A2X9ef2Bs+HG3ysa2/CO5PTDuxbksuTZNYgw
4y6DwAZAy6lLPKNqspD/P+6RThIqagVRcfxhODmZNgH8iURm/piLYwVGbv3NgM1w
1blU0fak5ywzSh3QEOKG93Ho/AA84cjNDnU+qUIz6xiDrZn6WOEh2cXrlGSgW9Bt
fAwBDEdmXDLd+BtV1O7aiCFfzEzir3gEAF0IP/XtbulAxPo9YNahcqu7GFY/q8ai
6f7vET0Rywdp3PpJubGUEYmJ5ZbBpI4aqyR+stgzSBv2r9p6rTh0Litpam1T0jmx
y50y8vYj/qWrs0RWnXh6xS0NgvnPlr53lpzxZzIeNq+fh+GUz2dpJtUr4dZChQ9J
OI06cOLA/fmma6J9oZIneadtsh79UR+1YjkDNWUEvmImnQAFfEVxX+YxCXfQ5kN2
ZfAIFwRbs3P0+QdLBKXcUwvjKWTzC4gFooJaD+tRA8EL2JK9h0SOkS8fMk4dlr/L
W9bL6YFnR/saCU09X0rrmNz3sS4wblXI6uBNkXLt4n94bhhts0UloqhPwOzlULO7
ax48/0sI9qbR52taAKTTwvTEjO5PaOQ1iGzaxPLkBvfeKipPhP/PmAIh3tAfobus
qnglZWUiEr/VAubn/xSsTB+ZXuwonHTmLTUsZJ+XJUTmq3/PRWAANBzPvx+Sfgpt
dzdf7CcLXeLuMWvAFmyAdli/1z4NLZ9X9XWvb5qy2o5J2U2yGLVA5n0W5FQgbyz/
oke+2khq7H8rdZ+7Oysh9Wn468vZbbPYf5X2Lq+q+opz6LO31omE6KgKgiekLeCB
86b8qQ5cjlxbLsfSuo3YoxglcIAMM/jhCUSUQzrksUUQ25rBsxJVYYlBTq2R+iBH
1NYaKlBmO28nq618Oe0tPLeuNn8MzTp0yXMwjB0VCAuAw9WQz7BxVkSsN6/CxINU
TTb77KFDQ3IoILpa1dRS9rPBQcNa1E4xNlcLlGxBMHvoSxAfJQ0OH0chjH4WzHaq
l54sUnq8xUHoFrHGnN8YQk3jAQv8JKhc3YdGj+GWNPNDQnwwjQGTC4pHcyXZbrrM
IJchP7eFTk2/MJKlMv8Ais61BDuL5dQEa3PE8BFclp0=
`protect END_PROTECTED
