`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btHns3ddHFvxVZntlCkZjoZ6QkkxNclbxD8pOzwzLgyghs6SGJrKdEasumIcARQ1
QPjdRaRDsc1sOqJ14Ju0goEqU4OxL+PCXbpxQAWr8yhvMGk93uiDujWaZ9duqqu2
ten6eh3u2i+9CAy1OOFp1xilRxScX1YSA86B5RL5U+avSVtkfw5omJIdrEMefYkb
73GPXQsBJvcNHmJFLfbBzkeXYh9phoUqSNEFgLcqru+NMgtW5310Ml/7ertNmOZs
puhycJ86FYo7ZNip0KTlWbHTPVT5pGc+cmf0Vl6TDJZtIAyn03PBpHhIS9ZfNATF
hkJRxIEKl0Ek/fqbFwXX4z+SlHBKTeUaIcC1k4FarupaacqR/IGZcvZ1Uj8YNEze
S9EqjMiQo8rHkaJq1nTBa+QvlpkQUIv5MfhX2SdeGhtH3tPu14G11hgMplNkg/h0
6J9Zu8MswABsQ4NfQ/dVwP6hfVmeWjHh5u8bmhRPmsRNMX1rEXaadSlIAC8HNo9N
MdpznaTsPXZ3G1ZPMORd75hfBJZB9dh/YRovWfAc/HDBdEYf1qV4Es3si14s+DsE
5eqi8cRYLmdOTWx2vqbArjluuvQ8QuJ1LURUbAOI5r99IPrGe2CZRef9T/aig6b8
i0n43NJq+0fXk288fxKHuXK6TevlADyG0Wbm6ybsklvF3J993j9Z+eolpKG1KrVb
/2LKcjV8yFtaROF8I/+UUI528yria9zZUbv3J2E+2thIItsEsAj0ZFie60wZdj/G
QH2iHZWAk8VPAqzQa6iKf6OlWWWTHQUIq+fI/h/5prXrZwypg59ZH0iRT8Ih5IIu
fsb0X3DCiIqdkkhm572SR7upHHkgvGJceGNW1UtfBqlpa0cKmdGvr/NmkNU5PH6H
RiqHzczvIZH8hMws//99/p0x6WeZnZ+i8Dmew7tdhSY4f4WvMCBFnglw5cMJE0g2
uVelFXmf7LHGJPLG9lxGccBAzWNRIpAngB7mCvL/xbE1AAvlMhAz4O05uXDU5kLX
4z18uaCFWBCwpuzL1YipFGJlxlNUnmSvWWuZrftElxtWpR4l0xOWdY1tU3zgwKVb
8UBaO9cdXvaye7mmGCVKTiUnbQhHLxJN34dr3LA9Pwfievgf7TpSz+DDIZA6nco1
ys280WTQOAYSMUr1xipnR6YDiPTbcNdZRVBXEc6NjVgblDKmTaIwncskoIm+duuM
LGZGHBb7HdelD8Isq5V4wR9Kls374KLL1zEkujsZIn8o12Nxu2ZhXrtnqiMFa2Xr
XBCL9ayw369fVylz4XZsoM1aXqzS4MM1if4HLz0KYbu4BSZgTDUph0jB3OTr+xhN
`protect END_PROTECTED
