`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a79KbcFGpzpUncUockozwYrOSZIl7XtMbemqyG+FnOC6Z0De4GtHLuxyq1ezMl3h
XzWs3OMeWeb30HbFiOQSv8n3D/3sUpf9H/z9J2hyr9ognDeOPMDQdzBYhH/fv+mi
fUQ+nJHhq6RhMCTO0589j8ANGYDQ/Oap3RSM8zSDSKTTlubHA01CFhdpVlty8cms
Lp10mehTeDAEtUq5sChQqulgGXCmLpk3JhWgvu4ho4RRz5Q8cObD89Xl6oxXQK1Q
xPL4j1f9XOdm7Sfk/H53zY5COEAVvjz32EYdg3sXUUNY9rVoXMg76myJe3gMWsa5
dCOT0DNIO0Ty40u3IvRpvxNgaUjARJ/8PYCRsO0GY9W4eBfSY9BxevPQtVANH5EE
/RikKdrz/RsBEGPx8/sm19kCNQEvvjBTj/cyYyLnp/KxvAYDVnf+EyjQuxcGmc2Y
pQr2OpRQnyT+6N0zYtptLVpgHt1QryVVtvKC0Mu55zcnewthuGb1e+dWCcNFSk1f
kCHWHSoArW3nniTHpEC1k5Z6/08LKNGEKuv9gcalHRfd9GhTYZn5cYEMfhiS0B15
iflfYA/cUc7O5aKeCpNKUUwvFYUjkBMtWqA2qSyVz4sGKpgMK/RJJLNHBVIdqFzk
3QH8pWDfSP8Otz3x/CA2kv87z7GBsmmxA5pCn+qKYKaKwp/SdRysrA+BJ6oQruEv
jW4Td9MWeuCt0mKD5L4tfHd+hq2yND1XoPsNRdy593ZccPJYv3YZMLmRGZDwPoi6
`protect END_PROTECTED
