`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PSOJFISGlpdRoLmAbkEXIKfrvJowP6JQQSmhSElQ1YzwXhM0MxuOPl+CRrQOXi1C
RZakH5hJmWO7F1j95DbyJIeh8kMALg02l/TXEuD7aPI7+OI+la6+Y0bCkfm/TQNB
rmfcmQ17u8SKiB/nk61I/blpsiaT4p+Pbmv+9shzTffP7EbF0BCFxgXukTFvCTlK
KWUGiUvORN2UvblNfb2Ge5mG94eQb5c0WF1zdCWYDbU58+fYGsSWnRgIsMQuhkHL
cINKbTWWcdxIOpnWKGggxRrWc6J7EgN9ySU3O8KGU4l0LKbtsExSrUTe+Cd4jOBP
OOORUmoLTNHeUacBdeuQwiY+XYzKaZtvlcryexdpiRDdZdfdXRwTgBI6LBxkOywr
97xB3kcKX5gQVNzUOlxPP0NNCAZIXFnbiIc4n1Y3qKI1nB9kxoZ+bQCC/SgR5Vqa
A5bquzD8iELBFd5yhS4qwFnQ8/9b3NOeMq+j/679IMOxnAlzWcAZgwqDlAlzpR+N
RnvXjUWyg8tSWKfRWDrZ3aBtf4Nc76gptluAzsoeJqSNUCpvOnaQZu3LXNen7ywI
k5Ij68AxLGQzhyWrkeCkXKOgJrQ9lFYxDt00blD0BoGB7Z5XktbHxdBMhkh/X20B
y1RMPPwcSNiJneJlc+8/IvwzoxzAOcTqC4w2xMqz7u+Md5ac2dUl4hwjvRdjAcjR
tHLWPA1h9Ivp61dh9Nf5toie3EX0kJT9L/JMOa+DOMHLysZWglBkyvDdDr/wdu8F
YlN7SpQEgOMCpec5anyKCT8Egt+zlGL++LxNH7aCSGTm6qiNQOGKEw72BGC5jO/d
9x3dkRCwNFwG57o/8vHph5q0AdaqiPrEq8yxng7F55w1wevuFRvPIoX3c/0L5t7c
REaw6tLRMJSgJ1e70JY8lgKJK5fZxtK0xjkk/Tkxc4YKdHN98gbrtuJMNFdsLiaf
liJatcglDiyDn26457UGDv9LqxWyV2C4aF4Kn7cgzOzK2NwYw/GNcCaK476gK+ti
SnFMWCNuIFcPCRvlY1KT2MtcFfvYhONK6niuJNtqV9ojEXIs3suVJDdmXLSZAqvz
LjJelWDs9NnyoIj+ukWPJIkh6f3pvvu/Edb6z8A+9KPQHmoTFz767HwjY3TPV+6K
VkrWaROzYRxxCYyI17+1/DYCAYZBDiFiAnFXBbmQ8inY2R+k+HfbwnDKzJUnD82S
`protect END_PROTECTED
