`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XWiLREyvXlc17Ts2j4m0j9ZPJ+vHDtdNyUP5QC9apc7b/BnAEybWXJI0bBt0Gyd
NDe2RFgOzUxlO9hKG6BViAztuGpYijuGxcfDra8/IaVR81lIEM4qhF0uv/VVi7HE
nFoNYyA0mhuficQ3Lp8iVfkxEY81bozaKvCXnQh5UWjYAXyP3DRkjiM2a4FAWqsM
9EUkYe9u3FFaph0DrCoHWk+jkWraL0TvxyGWggZhtPqe8gOG/WX1GENIDQBGe4tx
RSsd0Cigp9a2CB8AUh7b2X8SxO8tj/c9IHfIH3FjUf9O/b6FfVYEKzwz47qOAlN3
d1c6v4eTgB50Iv+Xv2DqiE8q4KY8JdOeDNsbA+vBOFix7gI0W0H5gcQmCVBv9u0b
CdMysMfPKV5wIX5gB5PPLq8mB1Y63ZAECshHYAp/MUQNmoQuhETZKGddOGyqvWII
3MQdHauytos5ourFrnz1bn3MNXY678EK4dYycmhwO/VpQs7mSJ5uIKXH12Gyfvo8
9S17bnRo8leqKIod++fKQnlWwZd+BC2UodRPCrh9m8TerBivIt74sicjSSt3fo7N
FH+GAk7e9OZ4hdh5yFum2oySIxgfLB9YZaYnhq3niyfYITtyNaEaR5OQFoFlxCJC
8BxGcifT6rPhJXTdy23wRKNWC9Xb8FifNIfcGGnuQs/aDWgSyit/O9rXSGdQl9KU
hscVcFnCFw4iKoEsLylmv0vThky1DtuXHJs1ICxIWnW4j7c9NYe7MHAxJQBPZ0dR
sQft7sSG5i/CTwypDqz+1Ibn2Ldh7kID6tSWZHcGgGqVuYnYG9vAI5n3YQP9phZn
yzFsoaUDN9n95YjEplqHidMdPGHh2g7egGNeuMyh5/TOQJfSxTunI10dm4zQfqta
MSQYmfoiz3YE9B7CnGvhiUwwapWHJxz4vPKgtdlo27+x2e23RSeDao58NvFsCZoi
c4LV7vmIRXNlrBf3eUGjbEbZimDRXUbJz1Ai9tRmGQwKYN0c2029ytCZShgGDAOt
5P6KU6rfcu52SrOXbySo8h4tVgxMELBzlzkcZkJ++Bexip7TVWbZXYE/hUZxotqQ
e/lAYa6OL4iFxOVIAPEBxuiSf27XSzTk5m1dqrNGWEWS6fYwwH9hBmFLOXzG8UBD
wyJTX1gEO9z40nzeAE9OkQAOIytoBpoPVsVYjBeWMrdThBwtdbZfHFiRT3C5Q6So
RnzZ/2ulrBHUvxzYWmUXt0lX00vHJJd8x0EVdPtTOZkGY9tMHXvSDETB0HBwoZ3g
wVbsBryQOm9JT9lae9PaBxlqP2Q2wQnmLoxOpEv+HL2djKUKy4tkmjzc6SQPd0uc
`protect END_PROTECTED
