`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cQKl5sfdmQ3t97vHtXJuqIIDpRga2CASIK31NiPiJLLZgHisTN4c2SqGXsJbQNK/
vne9OrGdutBrTmVWb56IB8dlNAChF+/HYX3KrHYz9dvlHMV7RLWWiHKR3UzKJrlf
DwDrDCni0o8fwTGDiihB0T2wwKzg660dNdT/3fEC6PDtMNarj+n5uzwb7QHQTnde
dvclPcymggV5MubB/Nl/A53OfkqR5eOrUM3nGWF36jQQ2A0CqyafEBPVFYTsJC/9
4dzBrf3n6admi4sQrJB6ar1qic2iISlAzeJoW8dhDJC2gOpyj6gsvTtFL/6Ysy62
2tyYUrFgNZR0uECupmZZG9ovLiwKNncAGkcOiThWeZzjHEq96rs4kFMPHeBguuks
+ylO3xXG9ZUZ+klvXqsrQFzRBGluKCLgg2mZmH4Uf+0/BwPNxpNxFaf6SPnLAoYw
lPI4UWRqzqslOeCGXnT35vpbirWaPLCEfz4TKhCcv1Dk9OoKHlM2ARaa9hXFDNq/
2ujdT16+sYMPIVOrGEdI7YBg6ij8gbC/L8zelp4TOmRvBEEJ/SDYzmBDvN9C9fZI
ggQILwfowVzW/LYv5r8XTzdHbTyQPRnvrdOm2pwkYDb21wbua+rbnJGNBPz2ZE5S
pstGMtxYdRyiJX4lxfBgPzjISGikwrd6gZqpQ9M+8TGuwN0cPourfw325JLsXlAB
Qs5pB/tORmIUxB5nEhNesuPU4N9+Bo5T6iY/VU4ilJx03dM7+dep4ttRFbGC/kCK
Fx97l1A5G2Ne429ZPNyY3jPPYsj/QFRdAtTBbuuoCWKvLauqKfbCK/bfEJ/SGH1E
c8hLVMfkqI9hwequ1dw0J5rajImsSzjsz5OSh6odzOD8iZ2ilXv9F0eSu7SYeROl
wiagrvNcgy3XbnUE62arXJ4oF9LiM6lU62ByKNP50sOh5zXLcoQikWKYddM8nHYb
P5mQi1XNphe3iEuoCsdhti6aKYRmM8YqYSWiTfl5mVScyWNUsCRCR8PucoMW/rU9
jg8Px7I+KOhrlcoaAcMm1Yd7a1CWbKowx/BFOxXi9WnBJRh24hkxr0IJb3H1Riwu
1qxpP3OGxkzE4bPykkVIOdOF4uG7fGCdgFzok3MWC3WuSTo9xpkYZfDGoy3msrPI
bI7MRoGkilU6HHVuzGw41/Q429fDj1UhLFH3vmDoUGHtRJynCYfGTBOP5PHoWt3E
xLUOgw5De7MOmLxqASjv+bG8AcV1fn3NwwbvBoEKeWJqRjm5VBMltuVr9Zs0v0dx
k9JCixkPVKW7/1opQv/Hh0Q+k6tJQFp62ww/S11YSySbFWs3NGjOfCtSjjx8wnH3
cpI+NfO2pcd/8Asp+07LEsGVK91WKdgC1Gb4jClulLLxmOcbigohvfeRsxVCHCrj
S6nyGp3tl4xyjYWFbjOUwijogvatzCNn2jp9+hIIn5O/NMotTNEeBr7JLUooQuZR
`protect END_PROTECTED
