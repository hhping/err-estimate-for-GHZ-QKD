`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19ue4uedonqG6YhC8smwHNT9DTkVQYy+WTybkYxAaBBNKi6Rr/ghdNf4i+7TL9MZ
4BLJHr7vEkTWTGfB8fJtz/HYtCHyc71X2W2hX1Kla85E7RtWsQXjhu2VeiibD3ZI
cBC4cj490JoRGsrKf1vGZQ1S4cSn7mlTVClgnloh8ec6PkUgqfQLh+W9CQ506XMJ
UGxk8Sy7ikRKDlhe7Kfn3TeboODgIR6An7mFZSpGDUE7IM9CH+lZLfR4H2dah0vw
JbCgfztBPTTkB7VsYeklQWAc6P8Pl4xtIECD2uLHfJbwqVbjfLrrPJqypLqdkpqy
nRwKjJeKg/+xN3Lv7qNSoL5hC6dyOQxBGrtTx1JLaMNpn9ppGXXZ6leKBW0OT8vH
TDbtTT2Xct6CX5NI869rwclkPE9U/HUWuM+E+jSnkRxluQvLNDj6zituSE5fx/U5
1CR/Zm8Y2oxSkywGv/rmmMQ/Ka5gtSwHkW+Zczso3akE5Po03rllhvIfMIDqdAat
ildM/tDWG4HWwDjrLoVnDTt1+/h9CnNl4R665WhXGKnbvXAFScra8D2v1IJRYKUu
qjn1Yw8uEc68eWzGdfb4HVvskKnryO7t9qasuzhcE0u3eeSQooQAvHl8BMQxZDrs
PnCbLg/i0ybEu6ob8oeQMDcdisKMwiHUUjWxDJorA3Ijo9aBKXwlGNnkIFfbkWeu
RwhJePg5fEkosRHJPEwTnwhTbTeM54rm2bW7xwhruUC5UuDsxdPVU3AKNKq3IRzP
rh3CUgB1JE5om17RMmaxssPSDP0hMsauVzn88FbBf2OHf9p4IQUU4qVo+PoMEtVs
TTHyPftMiRsuOIfBXj8LGA==
`protect END_PROTECTED
