`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rc3UGPyxlJEBk3aegfn647bHRAShe2p5Xz0RyRfRZgvqSZkEYyUEMKdLnvrjSuae
BZlXOZyXcsG19ZBI+4Rhla68iYAzKmd+nbYdbunpnIWsnYYjtL9+eD6NA4ChF+HM
RZHnuS1s1eG7Htz1pD/T7uclEXDbOOOKuCD6WNXhw728KDvdUoqrUFv86KFsqcA2
bNO6nPbmjus+G3OfFgGFp1auzOPpPFlCY7gXdaM5YFAihM15sIfU1m0ZqJpv6Oju
NUSGpAHQXSW569uU+VlpYA3g406c9qRJIyM4xnovsPVN8lMvANYx4JZRq9OlVRX2
AXZSiE0R+uzHpaNNZx7j6UvZhR852CqnO7PMJYnYnZKzcTay2TJtaM5wk3xJ2ytL
fPZdXlyLzOuHycu7DxJA73TEpvcm9B2+yoyKUXUcoh+gLN+S/KkVWi4z+wQDXiIB
`protect END_PROTECTED
