`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYACWMVMhxu8Pvvbs0Ghss7PQQEjVI+fVgToqCgApHRyC6lFHrwXzqmEEu9P53zV
W0bTHEa/zsUGOdNEKSYdB3blkfSE4UIR/8KC1GAU94yOTe9PvQDsfCfcKSKtuHeO
JRunouW4zyjKsbaE4eUYnZUMZPjOR1q4M7n4KNU6eVzOEU64RwXP6vvdXRwq6pvu
26VcYdBa27rFo+QhzSsZJ6qsOxwjMiZQzuUqyqTSiQDOpGyTH6pqBfYeDCIgNSQa
feHJcryfx6YI3xrlzj019kFYQQrGbmeJ3fNdwhDzgXMtYA+bnakGhhFvHseAdSbF
biwLgAOzdjCEPtPoLcnCBxwwn995RSLmKE4fvg1/2JCEsNeq/ZsuoXOpJC8LLnCq
tbjYAi90po8dXR/YO4QJg4TxF6zq9kTmWYcJR2ucgclxHocfA/2lEAa1d1ECR2cB
uAJic48IlICN90ymFu2che+62Z7MB1ueYT111REQv8rBVKQ/4cX07w4JTH6Be8DY
XxLPQ+b4auhhcEE/0M183wr6fHio+7X1ysE+C/mTHrJoXemPaWQKrrMUO4/KbhnK
YLM5jBSA6tgi0Ka4ddmv+L2xd2EjJOA++4VrTMu7BpIcGsd1lWhwt4eMo2jm5tYR
7/fZ7fm84xBM79ATUV6XYxFG2GbBUXs6fUX+LuOoiDQhr30+l+PWWImSagIOJAqM
z4/uZmLYy/hnlghMuNzy1xlISxw3W/sUVNlO/aL9ilSd8/QEVX8D0yCsGDtpMvuh
YPnkamEZsiXYEe7VcT0HujGPjHW+sd40KMIWWu6xDM8NO+LunZgQTo2un+h6OYKM
Ficyv6JAVl3ODDgGhXKwKtHwQ8RGGwKAo8ga24Absmq5bnJI2kLVJUSOOJiCdfjs
elcW9LGGxOCYk77i+bZwhRxEtyq3wwf49bTTFgDsnTDW44+9VzU/OxO4AbBK3gLI
TOsNnE6+z07K3p9N7KPEYdDv6DKBz8hCazo0oPiVTRtEwrb1jxpBM7UiFp97O0UG
O/MZYL0CZzMWvrSA4oLpZvsOQhKkhP8GyXrBHVM8DrWxqkUp8tkkmiuT92VQwp9M
0FS5qYnLjW279+2YxEZUPEwhehUBTslUP5izANmXFqHSuPA67QNeUi/d8EBZojFv
ePCYdc5OIFKBjBWjbh5vvtazM3KoWePJRgYJjOvEvHVIeVJAmZ1KoU/+f6lOTq+r
pRNj8dmC7mqFMb0TKXNx7Cs3eDMswHI8vu3nS28lzOwRFveCe40u5+ntmBtJEAG2
4SLyv3A5eP45k6EP77+lkQwG8gZCogeecrllNwDIDp7TrvsTUxVgm0PvYe4TqU57
CPsf0nZ6TQbogRShuKhDLIJdHMc9AUFIYiDm68PlGuSfRGdJeMT5rolsxAc4oHc3
y4AIUT/3b7MoguLFv1VkLAXCRha7BmvIYd1d+iZ2E6fUCBKySoT7HgG7N2U2rsT/
tXD1ADjPooKGB/RCouonhT+Xg+Rue7cOTbNgcXAl1uVByVHZsR4sMg8P21TK8dgT
Q2R//4IaOpAZfetP/36X6L51v/UF4JuqCIYnch0piJMihj913Prdc9Ocn1Obsj47
i/tYfjbcKZ2Qf8E/kW0p2m3URnlh/rKILoYPR+hcdS6lon3/dz8//bEAuw4mlZ6d
oBJ0fiAGczjAE47evQTYGVf9PGVxcvVz5c4KAlLdy6pheZ6DhT0Cv5FdTQiXjzbg
xddQWOJbl6JlfFxaTw4vIgCZiPbi+eCvM1PX0HFU+KtTg9rfr2SPeNuTZiQ8Y7TJ
C+XqXg6uqUyVv9jR3By6KZ+4OQkskwKnf+a9XhL5jzHWu0xFjOgpEfF24yJX+SSX
UWP0v/R++p8mzBX94b3HRfYuzbBzlQJ225oW2A2UFYPQgvD3bdXUXI8IbBEFUqYm
FLd32FqCaG/e9GC/xnxIegMyrO9U45qxmYclKTQFFhrG3bs+OEIoMGCeTn3yMe7B
50VFBzKouN/x9ekgU3emGDvkaFPjEYzzcQGbisf490azb09XlLQTVPx7PIpdkLgU
Nn4r5toTR07aaucN5e/OoZ6lshWKdxx+BoRQX9v2ZblKh5P/zsAWDCqGaeggsmYG
0Y3rOEHPUxONgA2F+18Revs/7+ZRoc74tSAKKtxe7/rdVvh4oG9TbQL2brZwCFXf
UpBBHZ3rBhkOzsNLAHz+USVfwN1tV2OZvdA+u8fF91bVEdSPl0qF++ygclfmSWDB
6UL5floQGLIetyd/KVVqGEGOsuO0Jtzc4xyJ6ECj3cDcERSyDuUr8yzGUI7k4FIo
wmcDWgn12ZHjstp6mytquPHw8uY3/JZZoIKH1ANrit4L65JQzo1bqensKoLHUATH
hfm6KqnEKIi4t9Txi8E0s5LuKwlV71cAhYopu35RruTjX/MEcFFSejdnLytwfHym
AfxIkBCB7qQLvhSB7CJqd0Md/TZFmBwzrsdT6N072rdTIkRbjvoEgvkf/MFnk458
vTNW1xDzxE9bVgwZODwdb4CFY0t0uszkamo0LBbmSjygx8gpcgBjWn/7fdbwyEu9
`protect END_PROTECTED
