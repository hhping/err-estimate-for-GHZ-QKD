`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2L7aa0DbEfMAR97LM8KsYK6JlsqKbm4MYVM1nV6/tBenh958BO4lzM9yemnMFbKK
mJhurjV4zSQgt7QKZ5T0rF+cciZ1Wqe/TXbsuFZKOg52zRtbqivD9Emef3k6i9K/
oTE9hDhfkVrl3HHcijHrJ0aI3Q6SGqRKYFfq+SVH9UkTj23WPJIvLM5gwnNBu6jp
2OaXcTGDspn+j7jjPSPLGCdDTRzLw8SgLOsjM0q8DroKPS5F98jLyU0uXTIA+Xcr
vYurCDxRUjKfdT9LshUsiu0N4Ia81iLiyxTd3xl9GPMJFvFsMZGIEYSu3nMgYDxT
SazsMnjNFvBg8BSG8ICIZmD1FQ+5JdbsTh4g0giqo5ihl87J9wQMLPrJlBEimnDH
`protect END_PROTECTED
