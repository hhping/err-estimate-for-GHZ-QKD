`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBfUi1Ab/LUK+Bf+pcFWm2Vx3j7OheH+2SySenAeHfwPZwAC3SoB731yPbuDCQD/
5iRNZuuBjR3Rw4fUhogveudOQ/mYUaYuB3+pFCtfDudkT3j6MbumJvwIqoMmTqs6
m0yBApCM8MAHNNmxSWw5rpWncXj2EHUp8BXOhyGd686YX4hSWh/PMHDFEAXXC2Gt
Ju+qlDcfzRW+jdQLjElRxDzJv5gNrqDCeuZedp2j3IsWAKgtQt1toAJAykcGkTIE
PTuncYqjNlPkB+muplo1g59nZSIC7rqjDCLYI1qAsejqi8VU4HDaECgkZ3x83b8/
6wmJshi5RaHpSKrcJAAmHvKAZT6tK9UxDXXuL6heXrOmDcSLIaXV6K99SPUh1VmJ
8ZR65PwaC5fj70frb2i+1LfPZf/tk5m+lGq62nn7Ih6jM1rKBr4jXDeWLbyHmhgn
3dKlGq0wDCuCew73kZMbmBRyBdd4G4Ib20MOC069SqKpFLDYGvXZYQJGErGFYhOb
Cy48uhWL5pbphvYf67AIox/oFWdKYQC4iUN8wTj5Foi6AcqjzisdmC0tW1ijA2/+
Qaa7ulagSknJ8zW1RPqHWEEBsrPQSa4mn9Jq2UjAd7BXNC5j5Ky7FszNrP67FK36
uOcw0YKhVYoB5aPy+1/qv978dektdVK6GfDZrc5Qpw1ojQW15dve5YWpuHlMwaDe
cb1wq6O3Rhwx6A8yQxMiMJXVz0vx0VXUHU4q56neLQtGjLW48S6pMBMqOWi37Kc2
JENEq2kyGEVl6Gckjc26NBfHBSTTqLJcDfgVpSczZ9DtNDF0gmdlJURdFxCnQlAF
pZ2oZ/q2bNrVarODbexpaI8Z6DKT6w0CsCpoiTZC4O0xwfmuehG8K7a0pQgCXbQ6
R4KM0bdO/6h5PyTm+rFhX1zayNMpGg40jJRHT1WBtA4eQ9W1Bil9eBL7wzodEKJA
UYh6myjVRvgL3S2oBqb/KxDJCQNjzb8/NS20+oeS+kYNLqNEf4ub7ywCpfF28RWq
sMnHnrorJxkMdv5CrmAloVwgSH0yHiZUe+5d0vhBdl9/PUoC7etSZv+71gJKgOMJ
PlG0kp1NxjnVsHfRqttx+v5Bgr9oJLPkn7xOHkY3AW9LJHKDUib94I1AloZE/sCN
oN0kmZvgkGuM4zMGgEH3PFNWqYHh84QxcPN5uQ9y1WUGppmokdasGlEt7U7fhrDz
57A4urBlnU32hn+RinIWaFiDw93C0JARszPAHSDjtATKkLknlUt8BtU5G4ESivWK
tRG8DmbVoaXcG+XsZSwi7wD9AIIdY1GhgWtFxzzCjexute457ZYmXvqjbuHEih6a
AU9w0+hQTO/ag9070gD9bNSQFzhat/EN6CQXE50yudCwa+dN6H1UsOxd2CkLVNlW
f1QpfR2gAvCU3m9IcFl2Gy6sKuGD7SgRn2QhCRBZPMykmMTBSemU+6YyFke9aRcU
FPZ4jX5MuiPsq6JnOYn8cw==
`protect END_PROTECTED
