`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wd6w62WjFfU0FyuDqtWLkVpvynhydaSvAubW+eJmh9kKbaKWZ3haaUqi7ASS8zYx
z2WAcuotbl4KBZ2WWzYjgLzN2yOujO3k74m05vGfiSVMiq6CddQPt576miiqjEq7
d8sYiK2arnY1+44LCfmwS345tEJZc8pdIrPXzFg/sUX+nwxbZ9pKgv4cVCT0m+kL
Ps/AguWXME7fvfb0ZbOx3jzGWOjIla6aTDFYQEGG8Vw5J+qBFzikFwM6csZANCvh
thbzW4vKDKKEcRPAUZp/A41PSKFoWrkHJOAaYcmT3HwN8fFynalqYNLbLcWRYFRW
Md314r0Imedej1XX4R/agxO6jvwpZUu8rmy9U4SZ4OBGQcs+X0EWCtuFcxRCB/c4
aiK24E/kWDJH0qDtYiDz8EvkozmeDXK84cHdTmmJJltegjJOVfSUOFfCXp2DPwzG
gyteKmGPD1yremIcLljEt6u9gWSJEZy/YryrT2evzd4Xr9V1ZUsWaU3+PzmAWouS
Ql63NQ8gT3J0Rzi5IixVHvXn8lzLbWZzrHivknSLIgkAun8y3N3/Ojq0OKNSb7u1
iW1vbuvVbndYwCvZzP9qUsi34Q2ZoEs1ihoCI0DXsjl03HrHvqI2tacHkAT5Lalh
kRqKdUE2k3iIRrVlOU93kCAKFAFsEejEcQR3kY1Z8bKbMykpjTeL3JnRaaxWv/Lb
WYw7T3+OmvhuvUZfnLR5Ma7zyDkhJma389Fr75mEg0b+QvSIExRwUDPch6naQnFn
9ubMbB3aSJDynGYuxJLg8j6XW+3yNosXKxHDNj61kc7i+e2RTYxdGa15jj4eo4/Y
M1e3ihLP0mpoU8qe66fftw0IdsEbq0jcjdHop7TtOSxxZMkTA1WYgWZ4J3oKj3x3
yNnfdagQA7RizxrBF8Y86EDQGYUZiK8oD7TTwAnbNZDx4BIJ9SNaPMXypRlEE1YE
E2Ja4sJTwUSfGEiUKzorbNy22BBmp7gpDxiGoILZnBe5ot6kLqLdcrbIruUEcapc
zJBPXncGitc92CPuuxfrO3zssAw2Uq7M0USveXDbm4eh6CaE6Tr4VG9DACo5YrpM
k1jExrM/hd5GAyzKbqHZDNjTJliVL4zk5AMMjDnlQcwHIyZvmqpUz4PEe1DJCJJz
BOfyvqJfEz7SFM/qep0Iy7CxDrM7beTupVkznp8SVVm5cyw5fSq3aPF24gAHJuHu
c3AEse8l2NPRQ8TQ4w9XK6zeNhnAoXtwGVcjZJsVtLqf+qCb38A+0BZadzRwhb+n
qOsOg+mKNYuYPJgwwJedSDotjoot8Hvt6qjE4mLTIiY9iZKQZf+/lFJ8xpQZMgnj
mrDbeUYqNrjjF2YHlxzv/TCdSPd8hOUwEgLAkLokDyyPs2MKu5u1M2SjWhSidJu+
165w11QbQvKF7V/hL2Z0AJeoe2RdbjDJMr9/C2dwmHofst+ueOfzJ0DL16IZodhg
wdBuqPb503Xzi3/mS2gGK2Zjh/8BwptwKPVqZHLLPKuGGurG0RLkE8N+YkdcfNfz
UPHyl3G1H/gsx22MUfqjhI2vZitVrfqLeMBBu3UGicNkJKk+j30cIE19LGzn6hBH
ZNFyvZqWNn7LXunFGRZEKjE7cX5FFV/t+qJ4BpP7gbMRPehEhVVOF/wnfjtk42TC
i8cgfxMvgKzhbFi/otXKcBY2Uq/jJ7P4HG0OCmj1GoUo6myS0srOlrO9y/ZomZL1
BEz2SeNXfvWakXraYk3DHmPcA7argsIgOcws0xJK9o/wc9RmxsKlYhHSe+CWP5QS
Bu8bKzXbg8+InbJmy1Z8jpOYZbjm1WO+Eyb4L/19TELnpTxzup3GA9VvSmD7Mgo3
wl1it07sF0jZy46cSqgrwPedBkUzASUxerjGPfg9pwKbgwtscIoaM0DskX5BXOhJ
uIefEj2vYYJkXhJ6GNxHpvuB/S7PeEJgtBoS3m6ghR4dLWoHLf4GV7I/TmeTI48/
TsdxhwgEm44Mf12FDtYwFJn7+EvHt1oP1CQ1nZhvnXr1MX4N0H/CB8HbygcA3J2i
0bb6xPiqYa1IsTzvrXqj21p/TacEk4celBQ0CxUTBu3PtGcjupqAgqlUQgx4liD5
S658Jt5iWbS19ZeiDKi9jycxTFC4IrDQdOIRMBIwmvckyxOMrKp9fBwDUbZZtmEK
2jYTWwEV3tyNjZUGo8vOaP7EQLvOXUWq7lQZkQtS4GMLKHTWJr3Uz6gn7cyK2dFG
lLw6Oe/MM2agf0Kbv+gA5QcucBzeC+UsHvRpqscihHwRcdstAF0eqmoyt0OA7mvw
DqXXHQoIe9Ojg7usrqnSR7w9j/UON+2ixXVhEdPABiT0FyGwaOsuKQZ063jWdJEn
qenkJav6QHDGn0PT7hM49+0MeWYJqLH2WIWPTBYmOiIlVdv72JswRTZrJZApz7nX
dOYD2GRPWCZbbNC4p9D2qPJseCoQngsAmimAIY1Bv79lEdqscjNuqVzqJLCmGW2U
dBTYgwYFTj4K01nr/yzTfinxchYH/u3Jffj9Z+y+KvH2dI5qNhLIDRN2slLSUSKK
rFsW62yoHLlmRDXTbWDgVKa239FLdcL8tBCUWtQ9dyP3Sv/JigXXV9QyyTR65BXx
Y+TjuZtn5LTk3mRmZRbxFP4tDwloyrkFgsX0IBGjlnytbuFDdp6iIr4Ncb+ctOpf
3a+2cvOhG3o60K3XQ27AI3InPm+LRwS2kk5uDgP2MqplxEwCE+YVzMAjOy18YUCQ
jA0R7s15cf4TpISDyjEMjwOKG9P5oJhCaH1S1PZOMEBfqxcVyTDzJcHYyeSeev1M
SuK7NTXG7vPCNY4frijOCufBBFSQFiVqWtUckLXpAPW6nRGf9hD1TQivewLBhKlY
8WHiaLaPYs2MmvWkKI77Zdcfe4YRf9xPws1qtg2jF8XEFZJHXhVlQOMxMciR88YG
NR2ACjCS0WU5YHrTdFJKQr/dyrVxLYBdH7CbMRJZV98vmk5bfHqOTVn3GbY/iKPa
5h6L9VQbAAHvE4fdDQ39phZT/jknLwFOZl0IztblVb13Wy2ULdvxfFNyCDaDkaAS
HBB+TSYOnGcFFXR90/5Sy1fgH9QA+1aDD/+/X86hisvnkyC6Bag60X/e69znFNzy
FStBVVuZe5eeI2+CU2D1kaVARIkVYcZZLsQJUG/AwxgCd8DTEC8lerU7DJfJ94z2
jvluYU+rE+pgKOymlNF1qFPlHCR3uORQ2TYFuJb4+l4LguR+Vcb1FV7QSJZIR/Ps
SreyLjVH1LDN+6PgVktZUdEJb0xTNMdT48HDSRjawRpdol+o1oszWFGvwrj0QZew
wRmJT/SzXktsDggufseNGpV6co3cDoWWWaR3h17Bldy9vPJg0mYsivD3GxhStzaq
Ovp3clVx7ifQt9LpPKa5/KOCjqz9tLj6DsandZy9FOwUqZCL+cl8fgUaguJoCdLJ
SFNt6Hj6DnzeZFtY3rJBjGiYzRh7pcJWHupwujki/Fbmoc29m3LR/nUddwcaAa7Y
QYZTps2G+ln5OOHBwSPB/nZkmGArV9gpYUUF91N6zWRl21zH5GYFihK4To5P7bRw
poQxsZdXzXvnswWTxr4jMYauIfB5N0CYyZ0aSinVbu4XVdIp4JR7qlmwJLbbn1Sc
S4NaLoug7l7tsJLWBD45YyyC6AYE1H0cjpyQjiKRyNkiGCmrD1QXDgRudu8+aQnJ
1eO10BS/7uhwaM9BkF8WGwaPgTkh7dy+B8BVaB3+AagHLjA9OUBuRjvvMvvQXKMP
p2TM2J4Dl/5ir4r8w+MUSzMwKAEHOFxjNFXJNgLavDufZNagw7/Dd4dLwrW07Jhb
mOdNFXbK8pRbaZHGZutQd96sH/RQaN0n9fZI/xV3OAd+5IuLJ50rNUb3uQ8swxl8
wyZafkmajIsUO0GiRytUysihg3oPwRmvYYe2E2hi4mEP856L2v3T7RhfdLeqAgMk
y71I8ETyYxrkYtiZvp+WTcyNDhmi9KRUfPNvo0pTAlg7zZTy8clyaAx81xdYBMb0
FIxuI4rstmcoX1ES7xE6qpN9KK1XyqKAp8xw4hLltF6qBg3+R6d42v9vioAQetYO
m4Glj8ra3OSYW64pVD6I1pJsBEg27w/oMSYcB7J/uAY2Ghn3LQJ9l/WX7oDOJsJI
+IhOEATZ+2Q8zd6/bHBvZNJ03Jpy2Rxwq9fyA9CZA2Qn8dCKzJOAHT7o5K//II08
/i1n8xVw/2Na3hAEDnZdgXaS35W8CAFEJdo1UY/nSwB70FRqjRjmjZ3RWhPIUGDX
WW4H3NoBCwt60AHF1HkJ4tKpGtNvNe9P275zwoWVzX6DI37janyTTb91Ig0Wb1rO
z+L9AUiv6Ol2SBN1L+amxmCfy92ohLu92Cjst8zyqm2J0jpAxURsrIb61LJs9PeH
w1VI8OyOs2ER4L6DoE7MDIwc0mxo10/qJWasC7vByr22YvNDqGA0lmiN1oevy5Hm
K59KuhSHI0yjUxTcB9TRM2BrtmUk2YdjEZsp2T/rlHwyL6ITZqVpvCQ00e/q+xaX
dvX/uX8A6vCtvIfkMrmyosV4PVIBvyGkoIGDHEQkLtWFbE+hsKq2zq/ZbxFECQ/0
N8KHU5wEKSX3wZUozBKRI9O7PIZYcPQLRIImNLNQT3VWbyPpvI7D8cncI1ngkshR
Eu9svrjecwXxaoF1lB4vLtW1vUzpBfl2K4GgsdIx/G5i8pG2BOgxKT7eKhQnhv4q
BKo4MCYu7dYS8sJvqPlFfoFCLBDXRpaDWsemUuBIDVPjn46q2dzM7kX8NLERhEqO
pQ7gUNS96hOAY8hIdbKsHLc0aJUwXIRzLbRJe5tsMhd26BAS84riNAuP1dlPY73G
NAwtiKLMtYa+fuhL2aeiC5pkKyLJTa3JLLuyG1KHrRTWaBE/e7CXyiM+m/oMYONb
/HCzAO2FBAGL1Qr6SsG/Kq2DHz45oM2baf+qxdejDng96wGoPDkPKKu1wJOKlUZJ
RRBrn5czdIosBnjVJWzz4xOX8g515lZtq/VTizkU8rULpIXtmB8J1kse55lae7ka
GoBjgHyFoxNxAnLEF9HJH7dNHfWtMOrEnuVauMxdI6gPassjdhIASwrNlmNXkIKc
0d/M8lTFFCYz3usah90YgGRRD2zqUErTLry5gvzgGCtXoyCZHQKqRLqc36wRgIce
b2Wy4Zv5SccONWvmtESsNjfEQ5siHcfX/K8czP5INGD68K0aWhKoDQ+aNzWKi+/v
WV1wAVTrXiMPjGV6DLUzy4H1K/rYJkPEN3gJngf1mRvejmsq95UaLzHYFLXop71Q
VPaEWCbELGOqD9rcYJXofX1XdM2JQG8haR78iAh0AwjJ9F+9QpWfp/GHlSaY87YJ
qREI7TVEv8JrCA35vDFZdBRW1axMS0EVutHJj1DcHA1G1jLfLnffLoCR4HMAtfeo
qvICV+wkeyp1o1aojvQAgJXWFs3tL/l28RJ8qcPVNbQsdppBm2Q7uEq8rDs8h2BJ
Pz1GbHV0dPSBSuTS0qZnmLeOVOvgI/B0Otq8fT0dHY1nowJY1xfAgdGICXRiYMKQ
v+LV210j1peN8MZ+4tzaZ9EqivaxoGeWp2Pn9rmjgV3aOUGHVSn89F9HWiXtpM/O
RECuftF/QokpHXs2jnABaTTYi7YGy7xTFV2z0Uwvj6BS9szzaK3TrFTcRW4lRQGZ
C1MSQ7oQaucapsT2MNlB/JH639pmYnIRomBr2BPVG445FYWS1M+73ciYGnhtX1I9
rdHmvsGjX3WORUUjSLUvBNzQqdV9bCceJ4U2NmXnnuDfnBGHyBnZ9IIjBtMgGhEo
TXWS1DYGtjlLuXJiSfNbcbxsQ9T9ZvHs741uJ8Lwv09481Zeuf7UWssQwJwtPKAG
F5cHV9UTENLdWRAbj48ZfzksrEra97dLgyHTWt+DZrxpDzl+7VRLWXAdZQLpxVxZ
G6j6YogomR6ELN4C5vnFLSzcymlak9ZfItvB4VFJQST4W0bbbCDjFNqrwn3f2S6+
KS4F+gqQe+KcKQviwWI1sOF2XJMkWGZN6/lvh+uZ/yCNo4nTL2tm7UEdrwhkZhm2
qelgK4tSIj5R69jEzBxogmSolLnmrbd2XZjxY83m+S2gAy8iJZII49JBsG+NjZqP
Z1K65wzPL33d89nkLMrwpwDMtPmM78t6AgxDpzcJY8/ysMV2WZMNFgDIeEDLhxN2
/Q9IUl+zII07vXfk0gGL2+Ksj27IApZ5vi1TKurgfv+P33i7ql//fa1AbdgRvnyP
H+2DS/9hec+8+SPbiQKyasTZODxoMQuR9BnRJWEqs1jy27jdafMX2uOrepvybPfs
zJHJCrpN2sTv2VV6/mhNshIqyUQtMunwc9P+UNcHaz/uiQVSwfzvol0QMeLPTcMm
RXJ/bbU5GlZYOM0NxQTkPTN912Q+jayYrkiAHb323IzhJuCpQNwOKUv2R/IhLM20
KZq34YViemwaJ8U4ZBZPls3nglcAGYkObKwdP1qwKivMor0ux68izpzAZmYfHav6
oYzcIKOdFhhh/vuZKqDQck2JPtWA9pbblqOAZWGzp+HF5ihR+CB3AQPYVd/Z+YBQ
HNzwRdJVOBoo0ZETJ+9Q/AIs84G3XpJL8+wNYL1QX7yJkgMeSnpzCmVVIuUfvDiV
8v6AP5RGzw7xfbOTQHXmmtuvlpDISs/hRdCh0qrJm1Dq32YXz8tam/TWR29++B7F
/pOr5F7Fdabdk2J4L1Ok1awAQ9xZxDYU1/Emfmxg27LQw5xc46q4oPJ+1p5DaqFU
/8wd0VLAQIF4mpv6sh17fvnJZV1IsWhJaiahz9Xqce0hBgoKYqTgV7XfK6risuPu
FO2Vtnji4OlvzPQxTfwJDxj560ptSPCFQRm5cbgY5zH3bskSf7rGY8Vn/G8q0ahG
wy0BkkkAEMXSsPee9wQS46CrbNF3bh9yXtUgDCAIiWOCIAeK16KCdnBvH5K6qjfe
f6JKFI+0PBmn46nPrXn53jQ/W4tq7xYEzcbvVTDE9t9Mf8kOrRy+VL6qn3grSjWJ
75QOzQ/Av21uIHw+EVBEouWjUwaNDgjeu7pMixtfL3+W1Qpx26hEktakJPnViRxi
mvTyN56wSoj3Zgi+NaP53W7hkihcAQD9vSDsp/NeQPkFv1BYDr/pjH+oVsU2WQZK
PQfp9RvhJCWEiHIySwKieyrvJO7Trfrn+FycrJaBMrvdLpoLKPqtT2Gr5R0ROlnL
qnXI5Dp2yyNuf6gg6paK1ge0MZ9z7sOhepcZaALRS03bE8s2vh4E9njLDroIAA46
0oBxNN/z9x6bFC1yBNNm0w40EVRjTMVCPGuNsHihOnWKAkq5gRfHNLTXlMNfywlM
LaXM62D7TLMJLlvO8YicG0V/bs8ijLlIxaCAS8DdShIJQ/SZb7a18Tb0RNUtccec
GvFqSka0+DNeboclB0ogIFZpeXbYxifsJeZeacrN+AMWZugizl4pKDt9O+UCJSAW
Ebz3efwMSAwji/8/nc9+4EG4biQu56ZNX2fpvFyzxbH78s6D0d7LoHSBi2eSqYK0
RTmuvNOtS63RK9+c84olsXDC5MpMroD4cNJMKRwk9gXNdbuyKPFMTNZkucnl1IBw
+4m1zFF8xsPzz5VH232JueQ39GOfZOPB7qXJ6cJOJpOU6/YjujyPv7yZFLxCkiVF
4Cscj4u95eoabChwRLbECOAAdQYxtren8j/oLL+pMBpR2LTHn3hIrGaF45Gla2yW
j4KsAiBuBM90x5769xmKbgvlCvrij7FO+2EEvjwfW4VAP+Pxkk7Vb/eWN+EF8gd+
jFeBxAbMGbuvsAtUTONswOVYuj4jRSZx/TPWw9z4VoMoblht8O++uhUXPV/UBMJc
bPTJ2yLdupxy9xqgOhxuUtNoYWuqGkDq/ayp6KWVH7QjSaxnDbWFNG8yr9vX5whN
cfdL1KTzhDxhPZ2GdaqMORC2LTPJIR/HMK0WT6UXMQU42CzAU99M7voeW4mMgowT
cu+OvCGB7so8PaZeTC5YndzQ+npliodV5tr7JwRKMf32XfcZtw1N4Ptf5GZMnvFw
4k+kE6+0stziVLZQGvrLm9QNGkhEasrkqYQVJdJD3Rq2ajQ2jC4Shm8zqaae6pxM
K9lWbtG35ZgYuTZUQDkcIafOPgf3t0Wy0HNcsPfwIEEw/E7lsIARG+cRrJmm2oQp
9eNJ324eS948n3FAylSY3KaPkLgD4Agvu+riscrnfFhAV1+D7qjBjhg3OV+lqSSB
ug95ROJ5eJnVpxvmoftKtyei+HRC2HcWqfX8B47JuZKw+HMvuOmmE3rUlhzyRUzr
ova0Zr8T6hkJhtDClDtmU2vO9bk08SSzn2k9PCW8rG9F2VK4OmjQuQbuzY+4jmfI
BW/4t9V4lPKYGymT6n6LASTH3GxSYTm7VwrR3GmyeczxewI5//mFj7LYe0UXk34J
tGhCQN9abmnkd2e1tsP389I++w6GJhplEDBIaW0N9iH6AXH/2WD64agUgeHsYAX4
PsKPT+S1S7dMmDGKcQMQfNejDmjl+wqWG39MVVUkArv/Q9L3P7ZzTriTECYURV7N
nhUT1H1E0z/kOrR7IvQjYsXsxX7UEsS0DFjCQcsYOHi6V8zv5wrGDCiH2e2Lz7lO
nQzsjc1Nod2IYbkEZ8nhOpuKKOTgeWoJN66/WwSR8x/QODDtoubGn+yNPVMqoKai
5k7J8rb9IS/4vCC++TNTu1x5jPyBNpjvm9XOBgawX7gVueRN80ydPH1DkAhquAnb
5d1ho+yhLoy3CfuyCc/LuNW2sAidJGyE0qBXVCX+Sr+Wu02mndTMXe5HndTzmdQL
G+6qNYZ/fewNQED+JlBwrkkBwGZGCpvYmxujRaT4G4+bDxnau0LV8uF2TBnYxqcr
Fz18PnZ2erNdOy3q4T5Nl7R4+VMPAc1x4S6Td0Ez0QMvIgrtMYJbNUiEtk93YLwg
rAuYIcvQEQvUK3DO/2g5ipj3vAu+QaCo8hEHduOs133eZdsXPcJ1DBFDHT28EAIX
Rydr0ExyGtu/tPmbfC3eR0io309nSd1zofx+58HTayTomH5nNp1CARBKIVqkupsm
jW2xYQ6kUocHdATPIKUt5Y8MPfcsEA/jwxX9G2aqU0Of+o3nRnGwlFvfKRUm4Jlk
fGOkrio9UHpV+DMvX08YX9CRrdFiM8AHjwEcAsRY2UC8IJi5by4QdMODoBnQRHJU
qwzoz/+eFzf0M5fLfakOfjx2PAgG0aU6pDZQ7S0cQZbmgAnFL95LSBhHAxiWV/Jz
pjSQb1V1pQn1EXIAwU+5my9eHy+fpwPUEY3rhzNFHRH//9TJb+bdf3aF04rJ2dc9
XxlV9XX5YMEtQuq4R96qRXRag7Wse6phQZxKfg6IUaYqZywnRrN6vPbx9Xa86Bi8
eqSL6/tCih0ecVwoDVBarA5f5Nd/PK/hPncUYWlcIqqmFOwq2tP1He2KfD6sEj+w
RFl/ea7UoPu86JDH6bevS79jt0wgGNKOxTt5LMCU+sf3iJxskniZt0655TlwLz9X
h6a9X/i5IId8plByw9dgHgZswofXY2Y3keNqC7gGI+neRaIGES93+mg2gLNodPww
6S4/oXSzdiKGaeLh/12Gau5HH4DbJXS8mjbqGSwbwI00To5gKsDznwUnYz156EGa
I8JO2N+GRdQ4J3yKS87Ll9ea71J6d+jZhJw280wu+znKcPNVxZ8Bnhj9kBY3g+Bj
KsGLZjDhIDSuVBgrpggDHv14+R/Gh53MsyjmM1l2rqOcTtqcq+Fy31/o1h0rJo+R
YEZmOfnuQnixg5BXZBvkLVF4/D48y6sCw/Zia9wbNREEbIlzsfRITKwapJS8uBWb
05sBzqaxi8gn3/tqMacZTnZfSSLJkVVPcq0XeDjxpOJayYT7m70JAwdTjD2279A1
JphumbCdAysViOrS8Riz56OaBaM8gPucpgt9AmRXHpGQu57pWDyNIIICZjGjTNFP
B4zgozfHeY21qcgPl1qWMPkGc7i3meAEIaJUWP9/HjjdBsR/Uw75AM3ckPVXsBM1
q0Toe5NHHu+vibU9JJzPzlI/XL/vtgYi4hhtWfYyn1O899M1O76a6pB/W1gDLtin
89vdWqdZV56Brs5KD27dsDS7Y3Fq/U1bBVRF1wzqFxBSOfoHVgFZprqq8Z856Os1
G/3w1R1CqJIHaiO31o4U9tHxO6/p/eSp4B8eMOlAdbCFzK+/UoMt9LgTH7w9fOdM
U3XjifpWmvGIEb7Jjkiaq9rzT0NBL70M2FRKT7//hQXQOZnQn/b1fpaUT30w6Xb+
UV502u6+NuB77DT3BTIyKum1HfW13CG7igmB1r5JOXXun/5WlexzxXeNF5v73le4
oT8hrQLG0CfhaGyoHz/q04429+er2wH25WqQLfrqxAXWUCk6/Lmxh6QYZuBXKcBZ
/MlKHntT1csQgXoF2iCxfWbVGrRV0q9L4OacuoSYXkCCK3qB661CEv+yukt4g1qP
amOWX1PAVTAfbQwillnAIej1ZXcZN7FJPbDE4RFKIRhNOrBjBySj+l3CRLeuCren
s9G9/AhLXX8BXzO1GrKQqkk6mKls7yKFgu7qnkrUMlW/P50TlKe/rCcwFE6UmwD0
3HEvPrxL2j2ZJyKMLGHPPEzrxBGUW31In9aBVZqds2bf65X26N+ooUpCT9Psiu3w
NXpQR1ns9LmE0pvkzJDGmHEyEyYuZhSLP7CaSAZcb4Y2sHL/IEGHwGlve1s8/Sfj
dSvdm/nmiaVkKR/mtzdPPOAXiJ3wZMRfRjprk0wDTUjNTRObHPzvK6cXIjXukfzC
ttlncA5XknasK/27y+R/by9d7SJkn3+XDOUq4riKZ7dE2SrLrij/DgNKzAvTSrEo
sAYx4zQeQksC6rrg3YjWQM7QguhaG0QWgsSQ5BMcwlxUYWwpNlI4Dj2mxXktlFEw
V0wWFei6HijLw+s05Rr6KinaOcV3I/AewIL/zYbVc/bou4feaU84DfGKPdv4toDl
E/5PbuZkYsjKPQHFJ+3bc5nwMBRYQIKb60YgThBoVw3J8/wvnHo0yDpskcI1NF15
XiuJv9Sb3EdFPPYAkiA2Vuq1MhgsmcgaCfJYHyRPanalgebq9oN1w8sycZFDZ16X
kpejTYGEM7PJvhKfceGYTieXxmJ4hEI+RQZp9jWB/db6zs16T0MoMicS6CbLM2GR
QYSb046FVJYL7AYdEY7k27InbQ+D+iY41NOzeqDoSiZ8djUnN3+RD7E9v7QhLMax
bMCJ/r8y/b+KH9zatVhtIF1Nty0VlU9hgwYuCSFUBp/m7tisNKJp775neLX3Ef7r
u09JV9i/DQd+f6jJzInH1EQTV/sepeMA6LAdvGRhaORwyPSlk0RBqnmo2qCSWhhv
d1tiEf2OEqVbvDJiLwloqdR5Bo+MzujEeVgt43NLnShAJJe4aDOaiKhDlw7mKxRy
R3IPcvzs4TQBNC4AsS6k0LnkyPjpFU7N4fuNUoQNuyg2qFuGYvMnp9GCDPd8Pv6B
oXbFpXb7jAQstP4w7YVkRzSu6ngwCLAS2Y357jE7qnGoQOlWO4syNIMZRCAEH0F9
c+YGRwiGsp2sMegjliFMknfWOMLuBwb2l4vjkDKT4JrQJMOjMArRSeawolfq7fkX
7kYwT9AgvIxjHAASqWRmuLzjoWS7/jb6kS72HfPvtwrbD7+vsOWaKX+TqDGp4pSi
SoB0ccs8CjupiDiXY21wE9kq66RlJ57DQeIGJ3nYjFcWNL88BqU+wvVLI6Ky3rYy
wITQ6U/QfKgMadVtNttnBRT+IqIp/Zg0z85o2AhphL4s4VDqvnX+rsI8BmwN5BXO
yDfv7DkomSjum282Q2fvjAkMgD5FhzZmT9nKwnw8hg8eJXH/7ISdST8dwKTMLx0X
tko3TYpny8ES21TciJACcB9c/zFnb1EwOiV9EeW+an9t/FWmrXIRrIDYDbNJEILG
gAHPElO1ej5zlVWmDkEMG/TjOdDZWUqfu2dURLG/Ph4UgrZT/XAxB43LMZVz7/RA
d1ViMmvgQz3ES4sJLigGb0EY+sUggHSyjcOoeyMOqlwxXasFNULn5x6K95H3C592
aQk3nKkuQo65+DXgS1eg1wkYwOy/OjbYLVeJoyQUkNaYcNBzu6v98GYSzqGUuBqm
61twqy645g9ijM+Rwxl/oOhg8/Zp4on2c+ZYTAfSN63Q7LbGfpBkLgkW5fLJpwEE
g7uihyjb65UsSGbVqAiYXkAkxieL1pTcIXr7A6vmplJ52/cU54/koA/22axgzSBL
wjtZviI7e5LWb5bkcovrkgj0Br7LvjyHOPna5EeIL7hQCI6X77qoydlvHoguhM3U
jkb1TaqYz64hR/N2bGoITFUCRpMdcKSrSOHt5j/KbsmMbrnjEjPg8Ov35VVNOOfy
s3mii1OmT98FnScXsliNgzCmZSov909N7XHM/MbBmWQpEkGgHuqQ/Pa9DH/GKXnu
rBJabHsfigaYauCZC+aD43M9hwmrkP3Nu6U1T+EY24BN2b+DzbjwrR+IsZa5ja15
Bg2xhGlZA3Vhbd3xwquqEZnoVs/ZJb/AsU6ZaiKrQjySbNTektYi65XXYjNd3vsj
XOFqHqxuVw+Um/9G0KbPsqO4o9mykFFgfHh2ycvoybvJapFor15x2Aa2QyB7DLLl
yp+8GS32Cuo+mkiKBY115URntGUlJypdSh8z7tlIOwgb/bcr0ABsp37qpce2TFlc
2NHUEW2dwejemre3oCdp3yxlr6xr2bXIJ4jvxAB4RharPcieagHaH5KX10JKKKQA
jCHIlz5qG3cFKrPQeIJg3csGBeIGPmfqdtHZEq+p7C01d0ZNzl47jwvGZAoXQco2
OVnSWoc6Ex0upaQVlF5WuomMSR2RPazNgz7uz4o5SXEIeYtkTvGlRKkL4BPc1vYx
agZWjH5kFu9RZGlMGIvBAiNQMXiQdSSr9+js3aI7X7PLj9CE8HkltcuReKNJinIH
0mDkEpRjAtoXYTp8p+Yxf4T/HFMBhkyTkbngMl01JkL0u79gmtLRBLcKvpF9Yxdd
9K42cZdLMyexUhAzwpMv6/A0NvextrDyF9BEYOuW7Ehzh37gyJEtlJuvJ2X6I+4A
AeatPvKSKrpH9wRygIjxgwMWAx70JCcW6rUp35fm1jpo76fVywvNZYphoBD94jDX
B1P98dgTN+LdfVBHVRN741Fhplg4L97v2Qxn6Wetbpne0yN/QBnUnX8dobwR9OxA
U+xDMj+tpv2IE4pLKiSA8o+7mvYoJ5k3jANfwP6y0v/N7yPTXxd9EWv8fTEQQqfp
LcyZEsCN7+4euA2RpwSjDeWBmdFdmQNnkLdKE7vAuzEiqHI0xcCX7uG1ukrJXoE1
BH1OruWoMTnkWXPW/CN5RW3yjgTVG1uRubblBVJZPBccl9c0Gu8aSKNECvaJzgDK
yDvDM2Rf5I+KY3sNfuH/ENaIcdmKBcXVtnzsLhR9mg8p5oKVfsGYhDPtUbF7THlO
rqCpZaoJEu7yvJvDaDCp6IORhkMvdEmWmtNn9iTvIYBlRvdnltll12zXY68txZUi
9F6DbCEGYDi2O8mykuL8ktMOTo6cTuLwI3f4oT7O9AiPIW9c0A4MHigIIJaYRzNv
OuGZL7rP5PVz1wYmfd5ElAbIWajofw5loonucDCcAvkEOQcsQwkkR5s8U/sXbsXX
NhsD/EiTWz+rCS0fTSljTGbw0eghsFp7wefoB45tkvU38lcAetjNeNJprUgC/QMs
rJt4//2pvAoy9v7YGlO5EhSrXyUzI+lwqxeAVDSI4XLACPwVQS9okSJM088SpZHF
mox6PKBHEmtR2kj6QAlWpe2zmjh0eij1D45PicgvHluPqg53ORXqxirSoicVZvcf
RftCOzyNEkveA7K3iu3ScGfEY7wzo+Jzu76HiX2TGYrJJVr5sl791HolWhXj7w83
QieBAeu07BT/NjUfj8i32VfTzlP7BqP7hHl+Ikg9U0nQ3sV8oY9XgPLd+j3t7UY2
ZZo8rK1CEgsrm2K6yStMlYDNgoXMEhhdPlnzxCumRJysRnNQkGr+fb/WbkaoiqKY
hDReo9m90uKKHz41/t/TeAv8GuTLlBvSAlSFliA1QF1NVrOcwcwaNJS0uBF4J7yQ
0VoyRCSjYJqbIwe+9lCyxHSsoJXOR2f0kgtCOF180k9a21WLTfgWC4lVhn2epFaN
S6PBdJWwg2cPJHr3wHxSxgh/0KXrpMcKe4/A/BnMhFY+rHu2YwREdG6DJA+dcDt+
IzELH+M5ZNRpKUla+XLOrYxPgWZXBR0XMGfS102/RckxT1W10W1sNuGco0hq3y1m
teI2rRBd3OggEJIaUmnaInM/zd7m2rEJ1M7UrEB+f1UchiUy8vuN2jt6VHQfEhIe
dXXobuPOWJz7z0LCSTuldXo8G0S2aR80xNtYgDz3rqnylxR6nfNNlbC4wAEooYE9
h8OQUuNRrIweFkr8nWHhhGHqhW1KeGnp6WAuux4dSI/nbslXZPL3kaNjKwH499JW
2yj++zrC8f/rYflPoKxBB0NGIPokwHvO9kBNSXnOMx2bKL/ngxBNPHQXCKZCqN+g
SVyt5rcu4gYJuU7nyVvdl+fASfDEEvzKFxvbKhxMjATTvDc9bqLxkSmEp1GQJbQM
kx4HzB6mh/8UGtZJhQ2oaXOsXoEkrETNWobU/yItjIg44Mj3FUC5jhhzp8dn3WHx
qe8POxsLxuLJwP1fHxyFodtPmUUgR8gOZHDW4C1H8JDURbGbTs7Zjp4nw/9OFaj/
g8+BqP889fFq1Ndo+p3VnVzwOmHisZzAQyR+tAxLG9wa9IurJsIAeEFEgsDEcm3C
my0pxNayCW/+ry6tHCMM/yKiTBAy3gUc0jkIZbeh8mtcluJa99Q8vHblBbP9tsNN
NVOWEyeEwtfN0mDoiY6CjeSW7GeWtLL2yGbhRt0mV6NisrXbpJ1Bix4eUBlBF1On
q9fVeDjU3P0F415EXS0ka4jQNQ+yCZJPAWaDB0ZKhgIBCkJgl4Elc48uScCcz8sQ
cDdaY/PoF0cQ626GHW1n2wmD2A3S0ZDtZQoHr9eFm9MUlzVJyWsubCe3CNgoA8Mi
4NjHbjTZ5I0YBT09gm273EjPd9sdbtEnY897eCAcxw6JOHznpYENf0gLc/pVTEe3
HoliiUdmeRrm3D8h6p3h2ClR7d3N8SpqErINNBgu9oWdPGRoxD7zG3pSKvtWRTfb
BPLgyY/JdxBDH8HfAIlx48F8cUjTTZB3/7XCDPHuaeeolZA+i9v0XvmPQ+JIG0fS
Xi0MWM3rSbWtyz3PheYvVgJ5egnrYY6ctaMZYUfCh6SbjZn4jjVMeKmx2faFJdud
dCIIWY0WGXC/ecuyQAj3pH6ECB0UCqhJSTrURiNamNGJaMJEwjhqJiX3zVKueIF7
yQ6KG+W93nWPjKg2sSpuhGNRUb2ZbXyhyrngTIDPad1DDFC1wtrq1dN8IUJMNJ0L
pjYyRBFdnz1IMMagUMR5AThlYPX1Vl7zcDSw307tQghvAsRmaDST88By9Pfurh3j
jwxDgBmlUk7bO6LMmdaG5HjWArnKq27qC7fhJ1kt1L/GT/vDlPRvKnR/NjFXoTJo
p9eqgDBXcZ/MPRwM9G2dEl1TIvNTOtMeQw54z1o6bxoG89yBZYnyVdU1K9pUqXeu
D2jbwstil9AMOConSRSVV59/EsMnjS7xfybCGE032TDAK/HXHxUNqqQMqFuvyCy+
+xG2248+A0baePsFtJneYv6ED0WjymSdkIOUjNM0z/VCOnNnTkTFWIB4px1mc56i
0Ku2CaNGHS1GFxQDzf/1Im4n4EuK1NhxcUgN/YlD+8GDiGT68zWn5kw3gdkyH4YD
jWMNfH8EfR/jXAP/k2DXol75Cbl2LASwO0gSPZdmWV9RJya9Piuu4fWgNcx2lp/v
Vtw9lehMkVrkgfQlNFVktFHszTSEv7TDgqmK0giPENzvAVv2unEIOozFYRV+wdok
eg/D65qEuq6gjtk+VoLM8tjj4StXqggifFsC0//3CqGErQa8IdWTvn0nA0usilYM
DUDElJeYIGFYr5TZhuVhDipzqIBN8cdH1QwkXb0xNJ8ptwP+XfVJ8qqNIla9ofa5
3FLTxO4poH4j3ndNfPBdRvFdRfju6+TS3z/suTjP6DeInVrMLWg3jSGv4kHMp0aq
dGfdYkK1eMN9kL8Ujc133XCL2OvOvXPnKHDRF2OWM5nw3vbupspNVA4cZbGgRGel
OadTrBpA5XgjE3MoOBXDLVLnGsjXDg6QVO7qfslOZs75Qiy14lFMaB9Cg+xvaega
IFfHcy3LjxrHX9PdhlzFy5HOXpdPEbV+OlnCe6ucjeiqRtLdYbBjte1OpgRjGocE
Mr7M3h4fAWURyrJ8OkSOai1pS/fHtbsILYb+uyUcyl8C1yF8NGkCMHHOwu0dcJy2
vqu2UGJRs/ORT322usbuVFsQ7OHAXcX0Xis/xeHVw2uq2ubfEHY2Y9g5yZGFkwKn
G9f7tWuMcr67tQlvChc+1Cvql/HbZObjKod45LxiY2TYI4WXRdMJH6sszPTV462b
gsPs0BJr5K+zwhSOBqWmPDeMvRYIddQOIh/3GFSKz1221GRrMJG4Y0xN58xEBzMG
Jmz+1X+UiaxA3Vvdj0slCN8KSsciYJG8HM+6sTe5lOQkOt2b/kQKYn/nMccmObtt
oawFBJ+lvP13G0Q+2KmRhH5gH7b7e+gn22Ph4/zGKiprVVuDiUjdlQYb1R/2Cb7G
AR1P5Ao+Q0yTKBXG1Tt+OnPRjHMlDDvW5O9hBdyZrM8B47g0ezc+18ld5Urtk2Jx
j7d3KNpMUQk2zkgxHR4dVi0azqnZPhFEkoVSxST4AESD0/Aes/3Bnz+RbNlDDjbJ
TnvZhm1POhBReVl1smr/Pu1gupeKH9Vptu2vEdC5RMEic1ODPth6iBSBRejKe2z3
dbVCwKhP+H96fjJUfZ2bQeX5f0Q6svLLgPunougUkPaglHzLOZdfQ6fCHG7aDpVg
GLRblig6qW7uOoXRrsnKoehuioFnsaIJGLKjWud2fwNNT3PjcNwa12X8aSC0Iag8
jT5drirwinDU8gjPlsTXya2er3rkBX9qnivG1VlEU+n/p4E18Jo5ebamxNXJvVqo
ZLSCXu3eVLFWZu2JXiJU+5mbfaiG4tZBaanVUHm73VMrALAO3gOdZxZCu77EiuB7
JOfystORrn0bRzh+D7xmZoxziJXtdDL1ExOCAKGoSnZAOzwRoaxTwT0TeKTXFB9k
UiHDYOdh5N2cP/qsilmVipeuB4cnPHBDc8e4eKPEAGDAkolzQg9Nbqh8N7yPjVe+
mYtQBJRlyAGpSv6mZbtFrn2rdTyonfrsst/JdjZgagQIACwPENlUkMGX9ZDYzkBo
L/19LZ0KnHKpU46isHpeduIBCobJeov3dOEXb5tHl6Ei+RLVS1Ha6r2/e8VS6qDS
Pp5WJkd+KjqZT1k09Ywaf9B6qbyGQS7g0QL4cAWxJq61ngeE9p4CVEjnlog6Im2F
cUmPWjoU3XCHrz4Azi9evoARFLTLCyCy3EL3J9WhQ6J10UaMaijQW2xi8XQ6ajsp
i1s1AfwcWxaGNrC6u84CCL2yBeSdurbgZI0NHgfsSExAy04wnpUq+/nqVjotn1yE
kRT+DrLSD3/3plQZYFecWxcoEvvcmd/SQB3oF+TC15rF16Vtw/4L9W7VjqwVQVFl
V7a/hM07tHFFEFRGxef3Bc4Igi35JGDKJ/tVZkJ3+ssz+/vFza4C7B1vL1oduPPF
mb8NF4aqMXge9zKmlMFWX9byGdE9e2xL50ChcefmIrnxTEte8psDZ/XJDd00JVvx
kglAsDfXvxZwZJ46I/eGs8/wwSpZuOGXbuyPTt4ZUg499QcygOYkFpluBWrFCa+D
7sDLuDQkJ7iBJjUDYl0DiPZW3i/QTZ5pCKnjWaOVdTVg//sOdeO74k59rFUTHiiD
tZjn0BcPNTIgq/KMczZFdGrSZZwFASg+AAj8iXFYAC/rSrVSENygW+HZT/ys/e21
Uq5snjpvoLMggCqqeL2dh+eEb38o3tyLgkqjwOo8btwcgBsKsixLkkSy59TX1cxo
AaSqN3q1XNGSWE2jYyyL3RE79Putips7wJG3AgnNUIT52/AL1qlRB7xjaMs+xEQF
U96EyPIj7CfcvesiJCV2YCEWV9ljcotOjDn2T0K2A/x2ZnXInQteuMz63UVibl1u
eovHSQRW7Mo8jI0GcetVZ7bPhADDz6OJP8yBLnL9gnKgh/3zARLpkPRsJgvmqZRd
ytrPa7M2fRBnbOO9JAgQ4+oAId1SlO7CDcIJvy5s/hWeMYl62+F/I1l4H62SKw2T
ZU/B8IBf6n04XRDQUAipKgifp1DjTdy9FmT554yLH968jOQ4PDT3DpmFVar1c34K
rtdjgWsE7m1dxgbgwp88bkPp99+AFZe8Q9fgt5MFmzJD+GwHSPVnBlQFLZ5LWhU3
FnPnRCBPgm2rDNq4cfK5YzYjFUa3+8CS2wbfHcBg7zUn9mulluP7/5I4Ggmdcxdh
1JrL1jd6Yt3WMS57gP3RDmm+9uPNE1oKkbL2aNJInjL5AaRBl/8NnI8gwTRZuz0J
zoCyC01v0HiQCPwZAWua0zXFq2DNQtR7kdHANzoiZ7ze9+R8sy3IDIFQqLTXx5pm
l6lc0Q7MEhcpGu6hWl+P7gJox0yzOChHxw3EAVrTpn1UJ2qbdBg5Jawn4Sf18uaE
IppHTWtJnt6daPWi93Ix8Xg2tex8/CdFTjZ2hHLWl2aEC++Nr/GobHwUhkGrbzmU
+LuVJJMlydEg7Mlf3BLabZ9BUdcf9ZQdkow/MOCz8XSaajpcociyaSjowfNqvOTH
VFYB7Il4T9/sR9W9XpTnxx96oTfVcbpv0bSSdzzoFVPTeT6ZPNmPo5S2Kqj4Lvzi
bFkPOsiSNjp0sXTG3PAeizHMFzxVGHCiy1T9VP8X9goTXhhuOVq5HRdjXO/1Fq0k
RHL0BNraiKkjXqi7rfLO4Ue2W2d4Br+mGRSjFPLSfk5TnwDdR5kXP4oqe8dhf1nM
aEbXed64awttUIxmFanYagzgbympHX8tK386Oga88VBUS4b0GFk3WNyzyINvlYHJ
5s/EvjwqiWB+OtZoC3KC9GsROs6mVOyN8olvRaYzj72jxaOp9sNAYqFIQRsiDQgQ
0o2ZdzpCdvuLrj9i6vcwEaWzRaKhfEInNCfW1m9mOviw8zMfoTKaXm7vQ1rGOdKu
cVJtm662Ddg5TxTkY6f3qFcI3PR+P8iPq6vpr1WjcPqmwGdZYlMoto2uKM1Arr+/
x+qQ8MOA06He4Zs/o85XW23b6dGh2PK3CdUa7XyB4atmKryubduSFmPzjuIzNB7W
zXTAq8WMOawAZ7NXM6K9lyyteKfVy1sIeCe5OA3l8xEXSW6eB4SriCcLsikSlOnP
WsDJgG1dpZSdtCY+IYci/gZnMmXNc4AMO3Uy2xBSK1hQCAmTMvN9mHAKejjYeuyR
PnJPXT0tnv3UmQMcHEsnjew32KtXlS+s8mLF2UCBSnDLKAj9EsIe+1+bGYfafKy/
E+YHcRFrkg6zTEIPFN0lrotUIHfJEaG3vD490nJoBUFDelsirYUI+QwyzNs6yank
quVFkcxSSDcuUUom56v7QVQ6kTq88sbJOR5j43qokso3qnxRm6RYMg77QJjMNQ6T
se/FLbsLnEg3yGO+mH1WzV5YmgBmE2H2Eu154zeWjF8FOWdWXltaL+J1dgRiXSmD
fae+ucmaJwSuZ0fC0D54mMXr4tIscksI6mzCEEJxb0GbawmmHuFYkoSW/POLjC+n
7V1jxyBcCB18v54qyEhTPfuWhwrtlrI0ElPVEdOoR8qUT2zt2bn8in0svusQe/cY
apVJnjUvtw3vfr4ujr9Xugm0cKW6ulHpePEzYWzLrbspBKhL0DU3bjSLc53Hr75+
gWuNlYzq0miYZf5xm0rW8x6Eh/1mlJ6NsQfcDix9hiEDqFmi5R4iCRx5k14U3wAj
SILZrQ70WvNVLuGujWs9a6/I4vo+90wiRcs7TEO9RAnbWKGi0nihOu0VYTYszwad
5ZYI9uRDC2V4iwzix9V0Z12HQMVki+pVRQJqxmprfggK2fatG6QsUeSgNWG2Z4+R
UgSaPHM0EBLhDNXToL9Lk8fIvbNjqRw5qnkruV9piYyTMtEAuTscIDLEZGrZTves
juQ6b2EJpI5JSI99JWTf76sSvjAJCcOOwduXXmkrYN5GUxOFooXWI0UFsSJTe24I
+Nv4Ie/6h4zUthg9GZXBV4Vdy/af9xRao3IBru6wsJxNApYkiWq1fns00eG97Mt/
xWW0EERphNDk0RdjL0giNLxw+Vi3m2R/nxxDuxG9/+Fg7Zfovh4VqUFkYrzGp6MA
RfPpY5MU9lEqB9PcUG41sQpk44zWRK7ZnHvl4xKXDicsZUwo3uAdC3oxMX6d1K7P
O3b4Yp/jMQVCTdmAqrsJJpxvpfEDfM7KN2cZBC+KxMSuAZJ3uxwy9VDjDsyytgZz
ikET+6aDXkcKP/5Tb9XFCmvHsHAKQbXDW6sSAjINUZqvzGzaxdudRz8mONyffqkI
Q8yFx3tnu1z/2XdE4Z2noOSXc1B5fmGqg2DtKNVnOT9mYW4uqUkbanQAzFNZ19sr
fiMq6VO4IATWCBfTMv4H6eAzB5WI+zPVPU2+/Lh6iUySU+juHOwddBdwkBgiC4th
OyivqRk5p1fPwam1rQIbJlPpIvjTwHneL7Adc68oQ6qwszJXc4tvbqtR+dcB3XR5
xxQ9hh1qVzZVVZ9hibrKgxUWBarPIwDUQDyeqb7L0tV4gI9aUj93q2LYVAYcjX5g
xcfw7pSpR/YKXv4/usyVE/bn8mOYWWXzFE7UI8V27aWQ1wPeyzNKugstt+NpzJB8
VvNO0UBV1D2nM3mPWVqosXKk+jPh+pJT8suWbOe2i6/jHT6cBlvWKce+nqKwNx2e
a3V0wC1MqKLSyq81z0Qt7yC3Qyugx/DxOSmyo7z57j1Abz2ZG70wvpu9VorZOKdO
5qIH0++KR1xUSf87ALv8uDBh29XohyWB9HYWmXzMdyaUCQnVA3ujfPwMbqQw3fv2
QZPnbLaYptLzlvBdNWBR+2O4bafWq4PImHyGDc2IFi4itoVQAX6Tsk02XJzJGxtK
/Ic7fGOD59676D59QiSr5lUsfFdPyhV/+J5CoAPg9GCG9/Y0fxlSCd4Rwvuaoi0M
S68pPsIq7/FCAAb+oqUesqqUBiQKASKc0QUDR7BgpWifkLXz3GVTp9k3ZB2/rU/L
N5cMcGTxvHtyI4jBVS9zoZ66pIpy98lPDrMeH29E7bVYtJ+dMx0As6LlkjAaMGmp
V7rHRhQi/LrtlAEwHBqJxw4wEqrcMJtyPwQL59ibsKsE9EhxhYa209HSl0p5s+P0
/7D1C0NCa8R1ttfX2wcnrvcEqwIlTasIXoBtI2WpQ8YtruWKOsafEB2+qGrx7nuF
hpUFL/7FicvJJoeEWUze2NCLBuompfRyDrM5df2QhaE4D8UzNur4M2rSIDTUChbt
PD9C8Ujq6u9eo1GPBbBmTEfwhgDDG0Wz3NAIfNXlOpkrGHJaTAXMrudMGPPsGyW+
6tjAK9YJecuZjoly88PG6qqgbA1GnPoCe2f24oeq/EmBX5KSym07omcNjNNP5SGG
v46zT74ICvAhP0a/vRBz/yQJ2uTZlsCk3ho+YIhlt8d+jkEnMrQ1EDiCvRtBGnKM
NVinxnP4xvb59E5rvkjw9CwowmwKVpqmh6liwKm+hP1i7uxhps8hb4u6tPSfaAZZ
BrYoz3zA1AUAUM6cAkx54agWFi1FopoaziCkszgq8QlEC7Rqn3ZhlOkGsdFrEXce
zPFTHM3eRkvf458DTi11czEsW4SEHvU6tmBoIM67b/e8iVJdYV70jAk5lRmiIQkQ
00O1sUu570catWankegsDHXvoF4cBZOPNGNzjp1sxScoAL2o3qd5jB/28kmIPjaI
aDtw9mX+8uBqVCv+nn4dRXk+ekOOH0Yj3plIy0zoC+/9AkPC9Ps0te6qF91GmQSG
U/+wO9A6zQpzwzUwymgVEeebkSFxDyTIi3wG/4leeUA7Aw8Jgz3hg0J2fcmiA5H2
ZkGlRJurEAo17o/Q2iOjRyFBIoeFKQISnw6fI9eXND09SlsILi/+Q1LE/AYROqxL
grmpkpFWhbNWybiWn56GJpsbJCCxEv1VPTQL22D7BIyvd+AI24VZHADoPNv8zpDS
vcw18hTCC4DyZDGaKEMdIBidr/uEobIryzg1NT9zLgNYaWIPnoypsa3MemzGj3aX
09WqthH32k31jD2qk7UjkDI8h0URwW8039kwXwooX59BsO87PGrQwLqvWhLunWvc
e9PAJnvaeqyDn4Iggid1cMUxn2ZOhC93JjmbGybqUP8wqrEE3Q/lnN54MjQNc+w6
UkYJqVUAT+kU7ObovgyojtDc+oBLpj5bhrAdNMgRqd72RvPz8NVgqAdd5w7N4TFc
18z6nxWIfDV1v4gdOJIT9pRtsWbU2MHdN9CYdM9WJx005xeX4z5skJRiDrHRt4QR
X+Qx1ftMGHXsp+/s3dMpdx8YApNxHcZoQ2/z7C+7mJ5MyU5Z+MHabKPE4H4V7DSB
Zp2NNgbKRh4hwD9EuE/PKtcGET8oww6KgoS1OFmhD5u3vpzw81lOhLXJxtxYeCyg
kYckdVXNzSzO4FJCjL+WtyTO36Ue5ZLAOr6EMP1GO5p+yTcuhgeTPEBjeLdL6J1J
aSTFgKKkSWWlkadHP5sGJdw6TqkW9XSGyicv3u/SO3MeXOD1wkiaq8NPtGUqHwFc
+tW78/UFVkE0krkwU/fNVjVF8bnEy2psDUuklOca8qdVbo77nbdIBwh90OTnZoGd
XKfApBxza+hCRVIz4BT2o5UJplZbYvoEDk2xLOoC0QLLcPgNhVIHaFAjqk8ha8aw
iiACV4nt/LrTJ9BcZogsvecMzIYfpszkvrMYpcWzXHvH7AiogqJiLGn1VhFJobmU
5jFS+7JmQVVV2dUYRAkQE8ewzfDoiTDmAFng+QNh+8Dg3+u45ilc8K4b4bmB/gvF
Pu9iuU2bv/y4s4gd/z+sRU3Rcf/Su8Z9EWP9DJTaVMr+NVUPSfBFY8mHPxKwrB9X
yA/nVJehqfY6Cj0pVyBzonEcGOLDkkYj7ZQz3zD5aDsgswxvljGTVtpxbSxUWYmN
LWKKYsjGncz7skJRFSoaiKnXUjJGkUhXhN2MUrkTvTpjNEB7ancX18Ao0MEPCPPC
lWM8rJA+mR5EQ/GeBI9znrocnGk4sEsqN8j5UtL/PpYGpeiW1hivdOI1Nz48VZJg
Kp6oqHuPjmUjF+PkGV5DBGxu6yW3UUYULfDOjBJgQEEFwkbJO7uKe7k5dqqUW3KA
0nM6DcRVnpjWipxB5xsX4d0uCfiX2WhbH7PYdp0eGv4NBMj25MJ+PSccRXCSC+xr
PNeqbfLNTo4ZBBY4zDxIChNO0S54n5O59pbIP6/Dwv9faPn22TI4WyUhGAKuBt4+
Sm/qLOhUUeSiJtHUqV0TrKSnPwImI47zW0EDz8ZufVoayrnkRumoY4ih6K/XOnVP
6YBr3JBMTWQeylaJMQ3Hv4JLDYihAP4XGZrR/oxcc8P2aCbF26KWqkGFEaJivq2m
RbKzGYmSKOC1DdUapsSEU/qcgU9nxjSIz28eP7chTvCLmIMXb+7TRKoSKf3yEk4Q
/QrDKrnCZ1kdAGCCEXQncvp34OSuXSBrnxpFMmRkeCWKpRvzPYzy7Uzc+6jl+3XS
iGB95awp16Du5GJ36Uy2faIPT2gw80Qyuye6Oq9GFVb5U6XqxoXBkLLMEQQgLbzW
TrXEAm1aOq7+9KZ++lWhtI/6nTuqky5m8tObampRSw5BINu+Pw+oVAPhGunDJLDs
Mv8spNzMwUnCqCzPJNYkpbQTbUd1wifE/bmCPcPBO/uk0wfID8cWzUV/JqWhrPQO
ULPxD6dQdmdnTh4Zdz6xzAq2drtKaZ5tm79zpSToeSKwkkVFAc5wJdhoe+PfV1/U
suHp2q0XhLNpxWMJ33FZINIq0RaibueNEzBZHuTM5oMeph61zrMXUUBRaCwPxHEC
zcKDOZ3CB1UGGbYr08MMqkWG1EndJNvbxj1GzGept/4SGw6o0gch/V7AjYZngchn
++CSls5QT+1jVTFJNrZSFZzHljTLWEi1nmDfia97RjlSVcJt7iyXV8SlbYdGzENQ
4HfMrCsFPUf3ZQj+AaDBdxjXExJ6reTsXpJoJOtei6Lal+SVvHJoFsx9pkY2BRRe
vsKOgb+b6Idjal0kvr0TCNdua/a5cLJ5A/X4KTK6/4mWSohENpEAs0Qg3V145WL/
V06XXj+k5wi93fS6HG2SV6ma+ZaLYWU1EQ1pgabQRi2L+UJctLnnNXJprsk1QA0Q
Z5RHne0mcBWphUoPuYDe2vItwAYFTPRF0zK0Ja8qjkl/X5OWRVsPSguWXJs4FeN1
aoXvgM5dNau20cHypvp7cL2uPjHpieOQq3tftycrNyAOKTDjFvnlNMvRXgvLYxTU
TUKKNsUibgx7G6FR1AJ5foDCKLrsdqm3tUV4UmHOUx8Iyu8yaqZoq4Xb3fsQ14gG
52YI2NCiYEQKExfjYRhShJz5wtjhbFgUMdPezo7NGRMuNBOgJcbBgcvSxLevoh4a
f9D+mwiq4QHopdR2G/JBx47O917AWpc2YxgkjUyS/9dZ3vacLGgF5ujwNCihfCL1
eZ6cFObHrzbngR40INilNrP8AfEkHAZ5QX/G26sS1stIBG6q8plxpt3SLe80tz24
01ugpQFEfwq0wxmmt0XLPDEQ2zkGUN7rQIQ8cKHFRtvpIV7LyY9MPtolsAQNQe2m
VQix4tSef+K2I6di5TSTKMYfFeHBabtDjlKiCTunmV2/7cnO2IvjGR3Z6D4GK0WB
GdMa8wc8oAyeJKv2S3TYxKFficNjnQ5dZNJOSnadMAyQL34sL/SHli/dAzxgjN+9
nxR63GUYobCGM/CvAx18bqHkJ/1P01tPFNrO4wtdoYz52+QgD0Y2AQRXotbBq/Kw
tN3BQUgv0+vJj8d3u+OIoswZGZPr26sUcRhzos9aILAWM0yTFZwejOopNxNhTlLE
Z2YK4m37/KyZl/N3IqJgcHEvwKl16bEmtrBfam0AXQIe4Wegp8oEwv0Vp3Fzf+CC
2eBio8rHjNEXocm6d/LXSiCHjeJDC4a3gkk6DQJulVuSgGvp/hmg1b9QBlE6XI88
rHe34Jw70tRh9Cfl+hepFqTQygptiTYfpsN7Qla5+9HSG044MWRCACRG/WDSCrd6
fHvVhycb8GSkublOEFvaWDUc+Ufp3vhc26nodtqRLw8wHgrvForVDnJv5lYNpW3A
C0G88bsF5IYRzl91Vv1MVyIjHTsROeGkqC0ckhDbTfRqRAcxHeG9Y/2LLsWdCpku
11Tkze+LGg4YRvTp/4J9FY6EkfXGE6iSyN8vf5EVq23DhUz3emse6d3m4YpGoJLU
5UrZoT7Rw51ocjgogbxMBDSfXVzHOlTcExQ7JKhwQR1ONX3hwnnYb5xuif5GmmWg
ZGg18pJzJ1DbhvHeHHNiKPKdPHIigoSgx2W4FamiTMZ9a0jvgIfjKr0gIfylwkMR
EhLr9CV5ZOJxgT60mgRIkIwCHQAyLdTclfuP4a0Iy/zcHOKf5HUh//EQgIDxxZr9
na0yF0OyuGkZmnTu6aOvPMX3Im6Ghar41k5O2HZWeCChh9vrUL35u6v+A+C/kF7F
rvmFiBwE/+NZHVy9t4+MlIy5r1oCRHI/Cb1YT18kFAdT/FjK2bUGH5kp4FFAUuJ9
VNduLxrp/MXmFayD3nj8POPWrkTdIaXO27B3qtSg6xF82vEoWUjLuKnoIX/zSThI
SRwxKdGPK2xsp0Iy+XHl0BTt2xNbTUiNSMkVrTy3VppzykfKw7aZVYsWEsJU5py8
4EOyTW5M0c4Z3et6qdYt4CJjaDpKA0DtZ62Ls4H+LP9+K2LpB59ELU326rcEV5bs
NJFCA0gt/qdc6JvzpIsyZnicZlRZUGL7Vx+VoFwws0jnfrHSwW9m9GDzqxh9QdlF
oTvUFi6vHx4Ma/yyTtsVgqIGu2qBA2sBJPpOrvO2kT+zm/jK7NudwADgPOFcCT1d
5LyN966jTiLZOJbdLZBBlpNmf3h2W+WbYNAxjTLwPMBwws+pSvspsRVaiBFdAmls
FuKiUd9V+I91qTHxfm0vlNPgVNFi6PGlNaCrTLNhr79LeBOmbh4Ne/DcV+rfzngA
WyLYoO8wzaiNFa6iUV6PJodeY36gDG9Uvtjx7ARPbQSrLaA/zFvzGcBMIFg2JZV1
zrmyyDpV0nFokqtiAHrG9UayUoy+ooBiujjQ3YaC68wUf2TCxiHKHB5ScQpPfGoN
IJoXLwuZTJ+B0rbgivbTbuMtBoajEjD26OHcaxVTob+ins6FS0NWPsAGuHKn4dzP
VD6ioFwo5siS4WTHfoEZBpg7fwUBKgcmskEBr0rpWXyIvOFDuElt7DLgbYZG5QFs
TZa3m5IeqF4E3B3d3o5w6E2lW5KDDwIIR8B2+aXUu+DXfdmAib2sCsk5UfFx7RTO
vOGxTQF9S1xqdq9FwjSzIPBwxoq800HMCH/skhdL3FAlzbUm9T95f531abhwBMJ+
xFU6tusof3lDSkDGvjpU7wukmclVJvMzbOvdoghMqoyoFA0njhO0amuFLFuM9R7m
Ay/uxruY+aqjYebHiJszga4YIlCbTBHR+xTnMhiyLOt4jV0PQ+Rj8XN6BWbKA1QA
2kCF9Hd19s+y0eHFYT8juMGLLFe3T1vJd1pM6M2QKglClmUg9DBryREMZWext8yn
4cx9pjTNO78ljeIWcnQB0mSrSWtEnfAwp74dig4wvJQ2YwUapxhLY3hqSuQS5J53
ar+DDFeEqaMBL9DbBljpqnaUiOdZqoLS+AvBZhrI2L8c2c4lZ/mU2o7xxGiV8Vxj
Q6MyO2Kle2j2DhxYW9Vsx3M6yg5TRxqXHGjiy1mS02ze/X/ABldPuuJiPi4nNdyK
LLR2Wx9idkQA1uoh+s3RSS9qFVRyZmN/m+1E5fqK+qtcD3eXclaZFZLQWD9JpMr1
czQHVmthPEmB4ksdWcHWPZUaemenjfoMLjlGOltHjD1fwK+OwoQAzROB4MEQldZR
Su+Llhs9ZI3HdDHmWNkc/YQSyseVwok7+df7NmbRsSrMVzt+6acElH3cnB7StRVN
KwqDiqM30Am6BqQp4j+DE5v1jC3uUzsQrIyfPKzwydTPxhlhK+x5e/f+qz7ojc3M
Y++3yrtWp1ES6ThHCkqmInHGJfgYiCwqUgWKrnh2J6rOZkLJAU3b5NbY/MDrTFB6
MYRAQFeRoWM5Wiq262KqkENX8TSXxki2ZLdPp6H5yZFvJI7TOdINKBwKizhobjtD
joQzknUxzheC547vVTvU2hDl5OJr0eo02aYVr+8aoh5e2d65PALlSOxUjbbgez2+
74tUMq8+z6PSudV0e7Vat6YmgWrzGxTId4TjUf88kkW/eL/3c9PPvYCPb2oDksKU
8npQpF4NXBYscEAPQnMwG9AkKPaVB0Vzz7CjE5brxjjozUrAmAHrqLVzhKYQs5q/
FHTRoW8fFD69mX+NAeVjUFBJzqE3wi6VlYd63+5UUrEQcO9ZDeUyA3Owg8KOxGRm
7K/j+NR1U+Pa+hvO5Wy1TaqGKqOarpAY77rsy3UvtVnI1wZdOXNr05FWrI+QjYjI
f5V6dZkDnitfC0QmGxFkKu8C6pA0GPXdsn2NWmumrUMaVD0Z5VKWVMe9XCpVRtTq
RgqiCD7Ufa7Y1pW9cA1msTrKWrdh1mPAKt0CrZPYhwgFpQvUyjqW1ZDXZ72emjJz
0hCKZGSNfuj84iFOF1ifr6odWfzpFjtxzrJE1RjUGq/cRuBjbSkV8RqgiXi0tiq9
qMg9q3no+g3X1IRsWkSuqhOlEPHz1JI+JnxWU5jvkWG25MTOK9ZbXg9s9sCCycBm
Prvye963dKwwWbMFDPnncsnppCNstqhZsLrFHoS4bbiLXWQpnA53CjI1Rk/TQExt
X2SsKrR2g5BRQ3Yh+DFkZS4zf0Lfmr9Am4VekPugMbJFlLwP+rOR4t+jYvSUMpjR
uWHwjxVEwGnr9Bm2thr+mWI8J3HSgbHrkhiiw4aj3CCA6mgsodnzN8umgCUug7Ci
suf/9w9GpAmHqMiL9Lps2KynQmp/p5Fst7vvCNUF/ZoZlXGTk3GOLEmsnEYGmmyQ
nM6vZBXGRFaCmcmwjLW4rINnb3ic4gBkI2rpw3OaQo34JS5DnXNeVRr+c1eBMknY
6SJiIKav7a6yKEPDUDigkf6/jxxo28zCteoRgEEM/guFgdYY6jeq+EsHLztMzF63
JSyT+sMUjacq9xfAgOY2DI2y9Pss8yJbaM8SiadS1UEO0W/4VOMhdrsG4Z+LgP4i
rWA0DBIxolmKWbNHujJCta7pdmhy4hOMcuih8eECWOfelKY3ai3vlDxax7Lx0DDC
5zTHApuFkH7fdlyxZ34Um1nqFB3YszFGEuWnqEjI+0wbfg15qJvrpmVfRyqK60vQ
+Rffw10uJvcZAnXa+15WjNeJfLDxXndC7NDFQVssjAPEOwfPwZC7SBzac/7PHyPV
xrceBAepTaEyn9HpQFo4V7dF49HRsgSGRuWbm3IF+AFLuz1G5/wWu9shqVNzFikB
pCGcwFnYuRI2cxjfjoigUAFT5BmO4rjazOiToYCtLbCpajcnw2agAo1e8QGt6+B9
iON3n9QcI2CY9DnuzuPQ3d0NJdHS3vNQDu7cGyxTj+LbxNcAbLGIuUqMAPHDvBdK
lUO1TLMJSnHAEhm6YfURShcOfRb/J3ZawVSz2miKP9l8yBDIUfyx8K2ZaZEdHm2C
Yp6+OuzGZ4UMtUYAObRaUooLpO4t8wC9cDtcHLVic5XfZ/xVC4lXArQuMiMSY6F3
4mvyB3i4BDkLrsJTje2u9jydPIvKN7wRJMBTRv4LkepFA0IH1UXuyA9nIjPu1Vmi
OFuFXs+m+n3s/M1nV93JxPt4tG+d8mh/skyQUx89pI1yTpMmY4zLdVezbLcnT5pK
lIvsleQ9yYMlEthWY65GCqLLOZn7czH7VzuP3Gn0xeUYM9tbnbNjW+1ntf6tNQ33
Pf0V0WM+n2isZ/JVP7zV81fQvhVhTbTz14MZTT6m+OMZbAZ1JSrOlRDEyCbgInKG
rg4tj60qJchDUaohfrUrws1EGGAb581/z4xNmBvArFAnBIE3mgVCBNmdxNV2hHqm
4DmQZHeNGtp1Al6ZuOEaXvk/RW1G/7csOnMCeWOqXiiE+512jPEaHJxaE177er9W
4WwSEY2wVy0IqhZTyQ3hMOrKuBlK74JSRLwhp2PdpMW4mgNThYDINzi2dklZdNju
9j7/ufiIcxiGc66VIieEFXdYbi4TFiMul2YXwgoAeGqL2Fj8QQ7ohUlpp9mzCERY
iNWTTLFLE6JI3OvJlPl2n3RGTeFyWXV2XEZGujO7/MunA05Dg5MosgOyWkgisddC
zcCJxBsViE/M9uYgaXRydRXuW0e4IsKqInQxYihynDqjmSC2U0I4SVbqVZp9CFzj
OvOPdq6AGzcAfxeUt0cQH2mdk+xy3zYCSi0XziX+M8VW7585GbLkHFbcEArILSLN
SNwYeDua8aerGiGzLNPZxvfkoG1vpe7gd06PZTLrY1CEiKeuf7TzZgRG6TErPevD
2ThEmYM3Of10v62t8r4h9jn5xLElcLu0ooRH7/P22hFEXQnimqxdydXK2Y8Gncza
my5nNqTwSmG5macxN7BagQU1lvghNLPtxg44uewnquDseXtl8nnLJutdhOja15g/
AmWScQ6OVdnq6IDqgGmWZDFuNw2pxFcxsEFOYEZSvxhteP2CtkMb2U1m15FiQ8yH
38baru76jAsgKRb8T1pf0j3Dp8U8OX959X+1N3yLSWSaviIU7RY2I84wAQP7Gcxd
hhlS8c7u1/4iGcyenhLZayeJtGcow2SmkQNRLugWGJcm8waFThaSszvjmAx0ygwX
oe46l/5kZR+UgryUwmBtaaiRTxMgQvCU/wANmyADrchxuvkVOnNH2cmGJMcDy3K0
la7T4sKOmF/zuTEZ2iyT/ScBCfk+QsPIDn4TR0YmEh4hc/+xyY0T8/yKyYvyZ7Ja
UKf201UStC0K+VmjFXcVpRC4Vt/ipQwnJsk5ujq0FSaBggNtrjSytWUzAtccGt7w
H7QVqYxDJvouL9eZQhUKkOsEXc2JcH/X9Kg88sf8XeO8UfVCD6H8w0J5Z2/QXGow
zFiaktwXd+gemzJOqqitTPAwgvGnX+CegiVIJuOhnd0TvKLlGiOXIsB5zZJsSsFa
N70Kv7enK1Fnpf3oTgc7rGNAxws0uYtkTkwOSA+/Dmzjvw7e3E4MA7/4HeBLK2ZM
w8lbZErjb/4gqkq1KdEx4Q5Ab60Q7bzTh2iOVZY38GI75EvR/UFe6EqslWJRjahc
SkWEuU56LU1kj6wWZLfmWEGqomkL7i5eUAb+W4Vw8UpINKeH7L9jyVvbTjZnXpCn
e0PeyiXRFZTIsu6DagVkjouVBNfh0Mf6rnHRquKcetyuq8WSe8coMlH4rUc2MUSg
35ZEcDchoV9CWJIeXax4INiZ+jh5BkJT+qn7U6HWcmry+CcpXMdDA3s9tmp0h/uc
ldE9Uws7YkuJ8zHxEZcHdWWwts8PGfQnYPXwCsOdBidFF1V/q2phIwBntLY4YXzm
aOTsO+FnSodfDzUJnm30TSkAqV08VskEI0LioViMkreHUg3N4oduX1DUrr6Qx1KU
mtailfYIdkb9by2iUQsiT5Q9k251Si77+W9pVMfOL27NS05QytCz0DvxUpvSpzJS
h2IBnE5oLOD++TpkgRiT6BfKuWgrszbV/iyGZnMGVRSRuqb/aXbQ1ulIkyk9MDSw
efQTnryalVSGJWfQry3EVP0QYqD4lTPAVubSfQpyMt2CsBx73FSY9qKd6l5d0g99
QGLsZVonCAxmztlRUu4ce5OaJ4fjMdJ3zCGXBlQGH9XAn6hqp9UWtQ99SbsW74o3
eMvmaJfmmzGtcbonXiKQTmBMp2zgvCaNdvweXE59CO3S6t4AYH6A4dtT6UDmbR1g
cxunR0MlKBtFEPfqPvXGH0vdMkT5wXnPm21enDXY8nhL8qS+jUSi68XXjp9kLFFv
LH/rN3SGxQxyH2x1sSxz7ZQsajLJMdEvTTo2OPx9m7ImL/9ROgzV6gTI2rt+WHFx
vwPWVDGvG32sBpWYgPlS+3Ifr6XMPdCaR0BMhqGlhCm9gcKIwhTa0LuxVUk6VawI
osJfseotaRLOVf+UDcBnw1/VRLizAjP8KlDsrhI6qMirJXEFQtvkWzOXQcwO7Hg9
F0wD16/V+xyFqr0T1EytqZkFL3rl9sl8ECxRd3okIK3nczsvVvAcc0LDBq38tzMe
iXwhXXhNCEPawrv4+kIG/Gea3oXyExDPLmVTI+BEJHmy/DBcHWHt80gTktXGYiSS
YieRvp73Fb3AbDugDTbkvUkswhon0n+Mvg8GM9lskJuB5fQOClrWeAIQOBX9pPEn
ScFMwLwqFORwLTrWMlKMXhHJR5UKAjRZakI+L7rWYpq3YV/pJc1sbmVigT9NsJB+
ym9GWNlpicYdpAW2Ec5Wcy6pvn5RLgdRRwo8Wm8hOnweh1HEu0y99V7RbvdMd350
PNrYwwOvTMYY1LIGdNtSu/LTyfku/Sl/GqAsHzeYqoQDL/ow5pkmMnEt6wUX8HVV
OtqBZH8evkx22fmiZcKemsHG/1Bj45v1bDNKUukO2n82SKW7hs+IkOmn+DRBmL1H
4UQU1ubkFR1vqLq50uiddKZ/z682zN67Ia2ZHovurYEytp8zNAat9WvU84NFUzyH
KgXEcAVApvNXO2IU2dn8uLch4iA43KdGnP1s84rnOmJ4acxzBhxJ2Tuafpo+AKPU
dy05azsAgrH51elNt0WXE8kbcqw8VChRKFKke9SlxaaZKIHiYGnrlF1ldVa1hdXa
ivdH9ntzKYLP077cOp/vzVaD8x1zQCFQeb1fCIfVdRxBiRvTd17w56cTRcfHamW5
9eMKQPrvfHGnHoWaai7EUAlE9vjkGPkEyrvBv8m/xGAuhtIcT3f0FQOnz9Apcm//
DCgdWOtll6vcYtfJspbcoNgdaiBTwJSJIcHUF4xmOxoejvd7fWol5YawxRVNrzrf
NZQjxFVxFo7AYWMoH3O945THMlCm23z3Vn3OVcd6iMk7rUtroLpEpwMLNDfNl27A
8LQWKWj1j6lKOy8VeR3Z0MSWgu/MhlSLP5j4PFh1jZJBPkNQsdn6RIbhc373Dq/6
kWuq4aCKqXAmyToGJe0Btpj4U0ntp4+ulyDBv90whSIPpScshUi/UTlir3hpY8mA
gGsR7f9Jr8+2iY9lujr8pwTIxt1DfLfzBsDhRTGz5yCv9WAB4xGRjRvebsUt3gJQ
LAKGV2SKPwx/aivRDX/xs0Cqv4grbVRtX14V8bgALbsemUVtuUWQ43HzhTIJVMey
3uLRAvT6O8Y7IEJQ9ShfTWJ0vSDR92lxf2bBzUGAMaOBwzxokVtZoAl2W1zSrefg
aOUarxJu2hpevZHiZhtlK9pLoHO4znd0UFLTUYjeil0lNJbXrOXAQOHmLnl0JMwC
uk1p8G4/QcW8EUPaSbhj9Cf0PLODy2P2Sk7habNPnocKTCINzJvbpQWqMBf9yuGP
tcFN0eyPzY1h6MJ7nhBLei547/hGnjd4hMcnqtcFdzf2HuwaB4oU+paIfB5Y0tiZ
TxYNcpf/zr/W6kGjL5TtBMcgdblCM8UxsVEjb89Cr5Y69nxLOCqm79QScfWUDx6P
h+gMqCBlh0k758j1pYfrcOi7NFxO9dDAhRc7gf0RKgv0SsQFdrAmXr61i31kBoyp
Mm8ES3qqnfbxkEyW6bDsDnv9ZFkjipjvyZfhy0baAhJsCWRjg67jlovzyLm1o+da
bpdvEPBm2ajssjLLt9YJDEpowAqcL6d6agqKIp5536J39rsUFoNxRNYMlawMKfTC
8gdtAu+pWJ2PGsLSeHpJsaXDhJKkLlYLJKIMe2NS7Eyu/JWqrDXBPBjWRDpg3/mJ
FvTsd2K5o1zIYHRwBl4TgYO91xo9mMyJui5j3q4/3JmsjlU0IjOXiVabbL/awoiP
d9/a6fZPaCKg0+/iRUvjlT38VUPtYZN4IJ3TOLJb0siiVaOgEPKQZmk/6KL+HR36
i0ppEs08J4+2S/DP5a8nqAufISGzdI2h0sS9KEsQgqp1V0rpou36kM8HZ/N6nL27
Q08Etcpw0Xj4W9/b8HBDURd8M4TWMyBOPHZaR/nUenV0OQUc74pCvjINkbhEIzC4
+AHvAcJt330kUQBU5qNPMr9cUp2CXcAK1V51OeCC2g7af+Q88aeLxt7lHHSyUAUZ
VzoBAb/aR7MyUAmxHSLM66J6vE6r+pnGoFknha0Zp+2JwYNb50ojTgyh73k5um1b
HOpBMCax/plH+mhEQ49x+KkNgA7g4tioSK5o4TDJBQjditweXrGJZWnYfcJi8M8Q
roewSvdM9S46EXXPaptejIrNIyjY7YABWkCZvhbj47Rk+QoIbs/knnhZgMAilenm
i5j9fUFazNK4NIBHbqwkPHA4QGPzEkfjwTk5G5cae7eaG2HDhtioElOMfU8Umy09
/9WiGgaIXluI5Qk1JNhJbD3vRlvQ86w4gpDqT23aOORJpEciWQsZwP4/WLSSGxAu
PFxMVeEDeaufEguEg0X04Cs7yHBoKvWSKuG55OZGHZ0/78UpVfaUbela78A4YrYC
XtdnFz1e3Q9Co2HQ/bXHyiDNFW5EVlt3oJqxaXt+ALMJ4MNVhkMYboElJCMPE9Lf
v5Nqld4QBrQOf8BvLKjdarJSOLI3FcvfSBGFIFFv52GoEiqS9RGFTvIzcoHY+Iv3
fMuSf3v7LGCb1EaS1nCJR15idLAzu8xbM/lZ6uDHAA+RTLwoJ/MsMiWWaTeES/KG
/uZBjZWdXtFLgk9sTRcyhBaGpZBvkBVH6XGYJ0vrI361IuqdN13TLbGHkRdXunMP
SISU648TWVfmKXR9y9Cu7BkGrPvPryyzplBgMrFEDwVsBaR5M3fsKinGymyrchFV
n695Xp/uaMGCRm4LK6aW0YalIP7FjDzHqOpXEi6SS8n0pHbcrVDo13V61oohtP2P
OTwpWsnhz5VEI5rQBUy6KF+xxMaRbJoIMjGdzsK4kEaYvK80WjTEY7Z/VId+gBo8
3yQeUZAqW0kFzpMF8IeiXw9gyRxXhnAK772bmwdib4NoikmtpVFUXsT7T+9/sgTe
gPczTEPrsiIik7TWxfSKsMKl4a1OG9wZnB+xBCVgJ2qp2TFdCwGTgv4b9zkj7ina
arjKqZPSXho3D5mVZnCGBRT+MFOsZWEXrCkTpB4DzqT3tIkc97uXguxZGtS1mt1a
Lm9PS8ltug7zi6JTRj14sOzRawQUYVfqfRgRfenmpsbyD2eOHDOEMai3kI7Sn8x6
yOzyEMTqtk/zvlAUAzRmCW5lOpBW/79ZqGKeA7nei/sqAXu80n9w+APPY8p0aGVE
RK6R0lxat5sLvE0yQ4EUQQyBgPLcOUBUXkt/3gLZyMyLX7yf9Q4gWL5Q9fA20NZR
E3UjsvXdiT3zRjVaskdMRw/3Zj31Z29ycBj50CfJrEp8pFjrydi/XIPJfWgIrsXI
MngpOeeYbM+s0laFQUTLMRRL30CkYReGEO01e7fgTmkSdXEXV86UJbUz5ffOMPZG
S+OlWLk4k5q4LPTXEL4rl8cUNvIt+mJMj7OpkC8WjCT4ml9SgNxz9aqA4ukbG5cq
bjzP17axfvxrbEf2G7hXSIbazrcNd2UcxVR3IpnI9h0/4RAM0IgPhbqtVUFg46Vv
E/yF7GWFvQlK6LoKFkUqmOTVmMM4BfzrXhJptm2+paPkEdk/fqRacIHxEg7hCt8e
H8pY8d9FZxOpUWoKiT/8S3CnZxQrMtijC1NGpFHToO7/mQ/S+zwPQlyZ01hhqvo6
24NSjM1t9+bdQ3JtNvJ43gts0QLBjUi3UIGa6O5Un426wKlfz0mHJqrNtFANrrW6
rRdbM60HZsLztRl12t2DZ7FwaIVPlWnpg/aogbUl6tOxeVzVc4CUF6aQRLXEdnW4
qXr/pxksnRyO+y4WldSG7hq8n2hoBWRo1pIYLqY1Kh/MHk6A7iHAXzG6DvgBnoZz
8QDKpN+lN9qNkjLr5BIjMpKrM/39ruKuZx8EG2CsX19ab7XY9g9yUyCDHud8tMMw
BE1bzli1MEIlLjSPesvFgOaCYtaV8Le3rVHwWuyH6KGcbK4rAUvPdGYoZhjM6zPE
yGIxanZil4In6XOOwsPEUKY4r/irqhLwuwDw496ftW5s1UCjnIRvIG08j3/N3F6v
EhL27wyKgGsjGUfyzrxcd12v+BYmlYzQRLiZ7bhFfH22b96WMOz/zUIYaCGuCDiE
S9vH9mf+Ju7ba8ySpK1M3Cx8u2ao4BeBGm8HTGXZlLH4ntvDdwKf9jNloF13XbOV
Ep06FWfmoH2ZirX9U0nYv+sQUPLf4EeqQX2SnYY6WLEE6qM9bFGWB/85F74SOBrj
X25UoTugdoQ15ohjcuxVn1AjJ/kDfJjxxt2UW2NFOFSF/n3ub5CpYagLUDxtXp8K
HvZlgZc+qWXK/jjbxZXzoTH0CkEYnM97S2dEl6WijJGP3eWVziqT1L/49Fcv3KuE
lWDt10iDSHE+dWv4MNF6xeXPUojHA99pihyOxLVjklmv2cyHbP9iUgGecDJCNiwZ
Eo/k3T5TIgVrPezX4llNrFgK2ffXec60GBGLLZo671W5U7f+FMsfsKIiP6ziqDY3
braQPI/sZMOOU7jIxxXlmJlrhiczlepT/mb9/t0fw3BAA9JQsUrmBiJKHgsbvRpl
mtKOi0Am+GJyAsfXvku2Q9oStsw23LTOTKT0Ztxk2HEnc5W9K5EoyxAsWO1OBSw4
Qa+XkitPEGQsSFWU5mLCCxVakkouc/Dqq0/d2qT13gATbxs/8zWMAhgFpaybn8nt
whhFXYXgUrmxneBilJ40OiBDHzTa/UGJ90i6P8dRHnF3pv9JLQlG5yQMiY+MlSnF
myS/CbUBAJ4s+jqG0IEEakud5soNhzzdHggP5L61zedbT9NemJgytV15J1VFoQi6
mBn3goWJVAsV9c4J5NwKTHfabgWzkPYSTCkjJj6V+ZA8LUZsjaftLMRHScoTkpO2
bMXbw2Kb/iDWYKXDpHHIeERoElHf3czC84CTdQt087ShbfbfSh0IFTOKKKty4rmT
rtw5/wdp2jAxK4Is3pSik/kFMvmqrrCRMSMeCyv7xa5JfONmwXUS1jikhqqoEypi
xBiuY228QFEouSqd5LeHYrKBpdtg9xCdfugYQNd9dQ4z7eqvlvJQ8qUNPG5t6+cq
llR06eIrfvu3J0/Z1R3L1oPRJU9ZzXIGIQEF0x0MIPU/OhdPQ6cwfvpEU0jwnEiP
6zb0l9V3SGdmRfbc2zL2Lb0I+svIAx7B9da0D2WeI+gS2iOsDJQqIUZM9PhEzbTU
aXyF69ktIL8wN+MoxCTrGahZxIgiq7rafFU3glQ60ZpWdmLdVaJmJ4crdNAPaLsp
L4nW6jXsKOP++me4Hlwoa2fFtoHhNPTsjfk6xZJ7z8D9uEfVJmaajldmDKkme2Do
KxFhNc79T2ff8yVaO94SqcZXS4Uh44J3/WL6tr/xLob1sRX5sBdNouVnXpZpQUu0
8vJ6ZdFLJJtvR0FyofNZpcnG9QR+04hxJ3NpGMIbnVQp8fzUjAFOOkXvwts9MTq5
5LMJG9vz4rvKfyZtt/SYVN79J/MhUQPr2KFG6L+xkGtHr8RxHA5H82ms+RLx4Iwj
0RHKNa1d3jDoh6Wd+HoInIqr0QX3MUsMQb6oVoH+IvR4fvbh82NVlMHvHVsR1HF9
lXeH55miFPs8fEfJtTT1lkQip2NGHBo39VY3jWIQuqgdJygkwRmg467WLCFe6Q48
1U1uhuCD3C0FYOkjDakcEYNwJQ+HCLs9uonkKzFkZN7X1xzjv2iDi6XJ1ZwZ7Ii3
qOsQ0EeP9WkZPW/nbeur8ToF/D0jNPBmevY6zpDro8+jdCTg1OXNVjmGokjXYNWK
4tyAP9Nl6SOZPhxKv/ytyYsJ+u3vDOhCUwW+gIqQ4FUjiNFnf/g+RDvlidzuSplQ
TFrJ3sv576K+XqGL1ACe9xgRm+9KwODXk5Mzk4vnFjyvLD2vxQGV9bq6CPWPG736
+04RAVb8DIStXmNv9RhZi6U0zQh4Szp7eFud/zS1gB5M1ayX30bS0uOGn/0r3xlK
12fFKatTpHY1CvlLhp1i0LVDcOy0fa2wUzWngQQYbAePSUY3k9yKetOQzAPQpbbh
TOTiJ12vPbRdWii9y7NsPlKrOHHvkXMlhFOaRC4N3CrFessv0fth3y91np5kBl5L
7r0rZMVk2j41qFl4d3tIVu9aVA+najjcDsxn4NT/iinvSxhC/8ihoamI25Xv3POy
oJ+lc43fiW9UMGYqaI7UsJak7V7FM6VW0O8XBRNysmFWx3HptQ4ANwUeoBGeUb5h
m4W3o8pKh0/1CFZlHcO8A5iMuwVGU6dvnxHTVFrklo61iehtjebQY3h6jksBm9/6
HkbiHOZeJXHX5vGDACnRk0Fh8U7LPYv8Rmj2nWROjq05ENJNoLZDEOWq9BKrvN1P
GSg2d9S1yX1E56BkKuJGOJm+0RaaUVuC3+PJzJYiXoGVXiRVTW6PKxosNsFmQXL/
Iqc+/jp851c2WgYqNS9OjmE9I9vrt/YNCr7+eHgRx72bAGcTtoHYb0PSlvNfedyZ
W1LKm8KstI1hH3dyI+trvYBeE/dvLI1s6RMKtnN1A6AVYkSRrDF7rC54f3APaDWo
Q1ApkA0jUEZLbUpBPQqyAIVOyYtneyfcq4hk3v87MYRWCKzlFFmcqnvXYDF2/R0c
JFTYMHfcRqUe7tO3++0+CfKXygBzkKtXVqBpMNNRVFoEoK/ukIEDn6eN3jkYEfOp
il10WNdmuHA4xN5ipkFqrwPaJKZyKKf6MVmvkBONuq6qEWf30Z77XqkEYA/jAdBK
lqQw5d77piVv7gsX1VtbzgFYd++glFIqzOXHsfwWGubrx700tbajfV1quTqNSplS
8/PpQoQepqI9OVPRfBM0kZnSaHOOa2fLBmZA9ZBVR4QhNOxb1YbopxQ86oq8RSot
34Z04bmFBh/vjSFjoJYvnhRTcTIzLPCAj6Iwu8wVNMe6J2jY2Y5KgYQbpzstOAUf
xbvhfmrjmbaV7HeC2wAYvdy4PASb3IkT4vES8hJ5d4/tpAWTGmICRaLvukS8kCvF
dwNiR45DCRTDEaQRPtJRhGzTItzqBnM9jeX2md4pkbodP3DSkRh4Oc+BKp3Z8vph
knH8/fBQ7oZpka6lmw2mQUpWIjwGBIuvTk8eKCqna/Em/mPUdQdmoax+IPeCvsaQ
ed8Q4qfJJDOqYSahmu/ELQTx8/dLp3TRF6DJp6Pgk4DU1SJ5H1NE9Fr+ZXt5wFJN
SkjKmGekVUqXHYy1O+kwZd1N2PY5zDBvoHqkbzaH+MZk3JAd3FnvPDp8BJrFnqwB
wwZR5Pc264K3RXKuXR/iaGX1gMFjuZZAnZ3jtfR7lObOq8LHzbO216/jYiWEZafC
B/HFsufbmRkjArQ7GT1hg9jGDry0nPyyNIXeIIOQhC/BIQ7YcedyNiDL5Om6ZNgp
2b4hquP+ZOcfgN04xN/4SxfmtF3K5nwMhC6YH6gYz0Sg4YBYNEMpI+4WJiqsjANt
eb4M4sHbfq3rZttBtGdtSMLVfMPsrojvTZ7I7+ZCIMvnpO1NkQ1uGSAjnIiCMMpa
Ug7mq5R5xGLsygSISW+Q24BuqfYb29e0DACx3V8AF7L2YGrK5QOyqKJ/MK3YT3kn
qkx1hW2zy6VGd3LJipK05RLrvgjdGcb9MD99NLPmFrfb26ZYN2BHD+f8Fz4TfDLs
AZfNhPgPw9INKFUKGNQy+1KOVmNtOlV48Yi2LPhuy2hHfHrm6WgX0p0/ZgyGjfQA
BZZ5XKIUXzZ+MMpq0sq+5KHl/cLiIWhoB5vNMT8gaSZ+6hyU32sz8fi9EvXYvXNc
qNidIhRRhxJ2Zs2XvK1NpokbfM5GojDkMM6KTxJT5MpxhA8xIUM/tzd8/OtGaTJS
wi7aP5Gzgzjji3SmBngjM0ZLdRNd8TjMZlDgkwuA2OLdVey8UtWKszcr0bpphVdA
/Nhz8sBZL/OHz4xaEjKJd0Rirjhxkikx6xK6jkFAqaUAAchM+FI4HR4J6YwDcfS7
oGz4QvX8LBooXCC32VSJ8UBm0WCNv+cC7YjshZTdBXG0FVZKdp0sFVe8wic9oQYM
Obscf71yysBlCfc/z9goVDylbuYfMYcGyK7f9M3px4LNrYnAy9Df/DI8BF8f7C7r
7LRtKxpw24PdXo0fPieX2X1Zgd3dfGu/GX3zFsCZh/bnXYHqwiS3Yx2Zad1keZ1s
qB7+kC50QuwbPGcUtfXNs+7EV5a+1MpCUOZZSQDorxwA9zpFfqC4Kz0h7c4e68AY
4yEWir2sXNVVnSNpT2SYIouzEfJESd71Go8Um2PI8VvV2uhDsw2EwugQuR/duq6X
NZ3ZSRocsLzmPfGLVq8hM39dgwIj4b7SWDXfMkubiJB0Mrchi1A6xtwCsbIDUr2S
6aCBdEMQwUA+n7DYld/k/gppt1soHArzl4nqtsKrqmI5qT1UzsO7Fwb1+nfx1EBJ
HfFYwZdSc8abK2lCNdUXpqrAJ2hO/EOXJbCtX1p2j87pFnMUfoOPAf/12qq2zr9A
tu+oySWPi3iMyeeyNtwkPskKESq1UI3qse6wvgzl8atLH5DZfqTXeAj85OggaC39
GZoKNSXhpTjSQ+0bYjzx79cbTymF7XiSlqkq5gdeN1B1e1r368YTpqybXdiiWjg6
fnp/I+HuZQ7v1MWjdyKCsbZ/XZMK+N4zTxaFdMWirQ2qmevKMj+hJgb9AZdLNZkJ
wXtYc8QmniREcbVrEpBwpJ554DmGGNCnii1dzyl/2JyMBWqfD/gFdiFN7TO6Ew/A
UOFPvWUKbAVjsthreFWGCZewix1pBYQYeCHag6VoNpZkFJ6rs6wVF7zMJi9bxPU9
knqMpuaPUw5ckPvOiwcgg38Vdf9U7Ili64GRsVWWS/3iglc68AVW5HNgKNH70OD4
5Dg/N+fCOkYcM6gR00hJ7sSrni0BR1LGY1zjhxmfqg635aj4W6wikBDooZtNYcri
FJDFM/az7PDMtbUMYzbcI+uJtjY7Ew2moVQh4cY3pOUxqEpClZPzNvj9cTYE8Xws
FHQnnRpEzujOue5slDOaVcWbFdnTNMGCTIC/u/D2W18++iUhGkLGqFX+MNX+1eMA
pAhWQ7OqU6v6KcqpmdyZNOoK6CE/NraWrUf0klVPywH0JmHa+zv69tkDav9eHdoy
duhFV5WXQEj91kf7cL/OxuauN6vdI5n513CXauZy8tfdUyZvLX5Y29IhCRfMd07o
1Vf/lXCeRY8AN58OleOukTNRyNvZOJNKs1kt/QHwpCOs5oKp4rTrLCx5qLH8/Yz8
wN8pSar20WOnGJBdQUPRKnWkReWRhSyXUiY+MmruVfWSbfx61jmzp92flkFIyYWv
74q/IlGVd6J5Lnlnh/yhvOAAcq/eQ5vPpyFJua+rwFVDrm6fPMnJtUHb+S9ry4sc
SgGL4ZrwPZIlDPFBuoXZVj5QUdERSifNmKWUE8qANRAz0XUzM4LQJYCuRyf2kP4j
A4fKghTfOxSbf5YvsBfFecMZv16eYmVdlXuDRMyZ2CPD/Q2gZmLkqGMjxBFFDP4t
iBMacifjCQxMJF7hZ6aLJ1pKpOg4KbUGpfBL0F6UfYbI/FExCHDvjFrvjQmEsZuO
xsu5WFeXGMjf8iz/mPo+g4WDL0Dkui+C7AVG6mXe9suffnLce2uAAukqCGS/5KLU
lsEoLXEAOhXThTOS7feXcU3fz+WlVNEqTerjXUa/8PVWi3sOObL61u6OCTSCgR7C
JXE2vzdZUsBB6Ogy9gtF7Ucto7VKKY+dtTW8Jozswads+vXrcOO1yrvzR+fKNbpM
07fRR9Ubg+JD3v+57NrUCMAuRJRHS777bnL5V+eYPkAhkWea0+PJoLUBFV/ZGUYR
q8wsI8ftMPGDq8cYTBdHEqXI2Bcuf06i404f33qoGjE/odA1Xx7HW2JgGGJLgqvK
j6LYrpwXnEhiXhrtSJsYc+IH4hkZoixZq7kB6JqLvlfVu08DiQuhQl3ZnY8M8Q7Z
W85IAQy4H2h5duimWt0QFPYL1GdReTwZ+Lw+7HUsKGwstUGgsCQuXeGV0jtaqNpL
PSN/HzhPgzRD69pEfAMVdikNXVXv3/cNBW4sX9rfXkEBHuxV11uDfOpxDRR5LGZU
tz2b7eUBgjZCQv/qqan81u/ysDEabdp/w+SsAw0WwT5/wbk0YPC0OCv3d12FDEhC
Td/73VefCl2nw1iCfoBmv2YbV+M4PE8X0i016/RiLmu3zqVrQgisPa4UqtF+hPcE
vje9G8W1ODDHzR+M8UDrws3itW3KxmHklhlltvFaMtBv39SN3AJh87kK2PA+6kxX
BE9d3kv5IUa6n3KOAW7AYpUuIbE35x94MusU1vpBDKglB1SxMTZdNXjotMIh2MKI
Ol2pJiMlCQ0hYGe1IlBwL/SGU3DFMrB/+vgVfpRHekZD7sn/PTSl4Z0UH/d16ilL
rZeygEXyVK7C34Uj6faWSNezZxM0ndhvv9qL6P/2DWIFeHnq8PG6O17nnxAuGgeq
6Jnvbs/JKL6Cbgw/0WLxJmYKDg6VXQA3cqNqFS/YYQRyGX6kmog725dAGQJ+QTiQ
6jtbsD+HlnfI2yr4YpMzhAvIdFoGKGmhk1AEoKcuOeuXKxZbo1vQZiB68nMoJpdU
EgyQA9Jdq6Z7LfPbpiFgJQ3tBGHwjXtxrOlJheyA0TVpMQq0IiRIBpm5DcsX320O
IofmU6jhPOJqjapzGgwC/c9yB5lHG5Ldd22XqU7bGHL1eRvRwZ4a3AlYRgnJ5rOa
n5kpsdoKHQpHR8MVPPkxzDt7Ec9Pn9ald3nkQU69UaBmPHwbVpNHIHWYQGUUkAoC
vtf9MmGPDM2tSSbye+lUEMvoWSM742Sglz6z8IpZ/Iu5nqJB60DGM7DToblqIhIV
zlS4lGMfu3PmajdJYAxlM+wd8W4u4fml7tzEy7p3NISoEoog4ATUJ9/k1rI2YOnm
snvoeVPGRtR2Uz9jjVDsYnlYvQGSPTUKI4wbPUphYTugObMJ7qlfcagfo3abjjWi
CaKG6na5ErhwAavIXvl/NveVmqvK2GNiypAFGkUYK9kmIZs/mc39k+LLFqZy/eK6
vNtCp4nsRjepE68t72X8A/np8uo5Z8D1m6MPX309GTXrzhFrhDO4qPfAQoWVV6It
5Y1mzIhDMuuskbHXMuCJZuSEwQyI1SDR0Kj9uNvVrF/yl89bIBiZWbZmfWuKarPM
H3DTa3kqAAk2wInDFx3cjfLeI9nDrGTCatGYl7WZqCoLpH8y7QmQOGUqkNaNTXo9
1bPq/4sMQ5zUqOYtQDtiVgPEXz2gi5HHGBu7UzQ3ipWdzWG1vaPs8pGEbILAkgoM
dHV3c49BJezO9n9c4tq6wP+zoMneIWXgpVyp93melkInesXAXkfMGiswCY3vmaVC
UZ6Y0RUbIkefOeCmax6ICJy4ZtvZIv0/f1s/Ok7B/E0nMCzgdfxjzlY08Xrmx9IZ
rNNbmCsSUesuOc+BBpiKdqqvqUneHGYJVbCFaDnnov5iIGy0zqpfh3uKVGF6BSKm
XxRp7mgc5ju3taw9RG1ymmB6MqILQyuFUIr4ANrr2MoVFxLbMR0AsdEUDdOPZHS5
Bmg4k/1hrTvlPEd84BO80DDLkVxlGPVNasKGj08tXS7emyiX1wGC2QGY0FVlYw6y
12tEGLcNSy5uPqteYu7i8nvE2UXWyK5fEHu2Uj5fOUUGubyd0dDY+6RjnaYWLLIC
hx3aC2vw3ZLcE1exxlX+d5p0gPCJSJ9Tqzg85asJQsPtS47z6mgL1f+AfBV5m12u
hob+vXmZA/Mqb4UnmO6fq3alcV/FDvtzrzD8GZ/E8bj2oHOFff4hEPuGWmX7NNO6
6c1UEmPG57dZFj6oc9alMQJLhWM4v1fvpflbesS0eiEJhBjh0K10ceUnOQQOfdBt
S2Edc5YqcnIJv2QxTJWDm7S9PCDwMhw4LOzIRLxB9im2P2dq0YikYfbvzCWkcXQZ
bo9sO7YhHoEy4xvYfT9SfcuBZHzIi/GLVnTeUxLRG5OGKPqV4fe9li9gbMIRCNFS
GD29Kx5RKFEO8pnnKz67W1yRHRJCElphLMRVoOPHs0omhHqhIaUn2XrbNXj3HrTI
+Q20Lb4AY0lcgQ2oVcVMgejZ3eOCVmrhCY0G7FtpncGZVPIKb41wQYYLSFNpe8n6
oV9SEHkCZ6mlmrRoq6rFTUztIsdo4zV/oVfDsrUS39CSItkh7QPsXWkICESXIH1g
RMyK+ZmV2YA7NMnvR1HDQPqiu+0EyTjoq1WqdaoQZhOWmPolZ0cHOT3B7AgDAqk9
TsQ575QZvrS5sDs1dCDo9fj06OIQhvWlx/+CJtHV3JWRJNlZLubPP7DGpM5ITBSy
xqtzeGTrcO/JlbGmsHzroZqo1mfiF+8Jm3WpSSawF5cHFsQzSbHTY741mXdUqHVY
WumzEd53Dy6gsHJVBPq35Oo2NXZ29F97GStJ193v5LOsnp0k8FYefpngYgM44opZ
yOt7fziWZpsZhLfu/npYP/IgdJyiTbvds0Ez9xMqe0f1LExZ4VSY1XwUjF+tM8ue
qN93rbut2aGk8Tj/fouNauioU52g9qyybdRmIlVx/s2nNadLnpr9C2T+4pgwve35
IILVKDQ8/RvYdEHpV9AHYhhXvDj7dMjHG9p++NBu4QbnoIxk+rRCQF6l67kwvvEC
JS0vfrDRvTCOE09+PFWHukACZEmChgzPCFQXouPigu0LYZ13URPEFyDEqX3++k9S
B+Up8IJGO+2TA61QQ/MrewOi/6KH/0/oQG2IYcMV57f9zt4sNurJ88t7fR+EVNQR
0IGIMev00KVqiWVv1e0f6CE0NIR1buWNnNKdVHJBYdRcAN/Ah2z31lJD06Q0oPuY
nv3fJKFLZqYLZ7GJr0y8uTcZTICRruf0bPverf6bwFIzpCP9JWbtAYmzGn3B/QN4
NF28xMD8ViytuZf4nQoe/Do1gKQdU8q5zjZGOO7bpeFB96nBAe9WAj+XOxNOsjb2
TJ4k75PNEv5VTkouAUmp5cREn/Zq2pgDX8IWsbYY55V8at0NVWVzUSP4889olO4+
QnIO7YwA5xFxs4mMv+HSRZNXRtZu4zsssAadp/weajObu+SaCdSau0Xih76ZLVLI
wCY+wgOvla64W2CX7opulWdFonOSeOT7Wqe4fgRGirmFFc6o7SpkTJke+CGVZ2rd
xLo/JMo6n9pn8nTP937wd89LTc2AizdqXoQI3W4+mgvhZN4eWfbrcDYVqWjLQYAM
1FQ3Mf8sGggKke1F1JXYO/FeG18UFw0UQ+pekfTiQfEtDzYoIaWe1gPU8wRljha+
ccw1+KPtDSxIrB41SbHq6ekikpgcRgyVI0O4uAiDW9cwR7F8K/c1EhmKYGhmi5hy
mnFB4sXqd7/sNscZDCuIVOnR7QFH/dCxGBZeNCip2VXfQzYtAHwonXNwpgDoATdN
KqxTqFHdhnKJ5lM50j0HbJlEgjuhCjgJrhQSOlrikigqC8viG5XUQjdrSPI8XkzC
4/tYnyF1iZkF8OwKzaqDtYhEE01wjm7Zj9hpAwgqOuOiQ8W+BdWlzxBEQ20ETIfp
RA8WVXiaVLd2w57Gl6BoOtPuuW6sO/CW1i8jxdhZLpWYtiOMDawkS9hRYei2mWjO
ImCsve99lIk0VEaDMQhEvitOVApTxcEAhb9BxAtyEJd9b+yKXoVt1uIWZoX/agJD
FqWIg4fki8L59oZE5JEQWnZ37W+H7D8HMga/FEMKrUaIvzWTNoMMneOOlV+XEPIp
SHorbgM08KVZa4pY6bmb1sjpqWKMKwwLzhSNhSOS1UjcwlHN6vJashqdWUwK1HRs
FS6LwW6fim4FoK3xQpLH+kaP08T8+y6psFPPQVBF/a7241KGwbQV6av0qjr/ZtOU
nIugGZBFZkW857QzaQHzsu71QtipL0WsNaZr+VmtWJIn/5Ug7eZduHoisTFH7xvQ
2Kkxn4k+8fPBBR3bl5yA6k6HRB5aEZte/48/ogt0cEOyNckpOUHeMiNpAQNNQWHA
Mc7+FgiqI5ntqEdT6DYFrMgpZ7W8FAry+hPjsBaSTjsOyewUjfmBp7sIuxdmuKDj
IvVu0vj13Wt8aKe67N4yiPhSLwlf+TqKrvW6rGxPaBiHRsZ0CA2N3oyrPO1UUsAC
pptom/y44DqhbqdBzApBq0d4gIUHdUy8/q5nydQtMLWS/ysXrkPkjznfse6wF8+G
Sx2K2GREk3DZblxS5jCEC/0xi+G+Egtei3vkGHFJ5pr2fX8+mtizwpUhEB+8yqUM
Y66QjbEsSW01rU/A7qb7gXn6kM3pfeJRuNECHvLse6pCAfujhELBegqUAD8KtRNB
LroZwtP6fipBgBrdAEmDfPbyI4TVlOxm2LgI7heZDRHuicMlrRnYCbPWZVZOjSte
hCS3UMKRCXfnkvxLdNzOSeQxeKsaRE4inSDkuMjICRzPOPzQ6afsXKHFJMIFuK/z
3v99h04DpruwY4WfAijoH4nGooQE1eaDqHD9peVJ3nkCcfO0YdzubUeCa7QhpM/C
CF25erwV1wo8wp74ifzLe7wt/wjLo29m3R3z4L6oBgvoehB/l0mh5mXNaOuk8nnP
VpshzcgB6znUtx8CneKbB1xxbDNla5NNVZlgDTl0J+XW0Rm21E58KRbIeOhcKwC5
yCCWCwi2FXVTJkTyTaXjyVV+Ah9waM5bSr22nt1N1LoC8E4cDhgvCuHEN1VeVxEb
XI7Tb+PYKFmkgTDLV4OwT9yyDA+zx2mMk+ganNSTl1XyvPdjKopGql3ukVY055g6
rxIH+d0XRX3vwICAdSXWCzDjHRnK+0VeymY1bi1gjgyPFql0k56VXF3ld4CIrvEn
v+4sXCyXQpTXNPTuTSboQpwJDeIfQnU9uS8qQ6Iu/v7Qyg2xy8874HQ9dpofVa2M
BdDqKDyz/p4PsZrUlWsny5+JYPgvF6Qjo4j27mohOF/nJyklFCtAjH7o4C4RQ+Fw
9Qw5CdOT2vjYEeQz+DsP2jUFdQKVZVWrHVQJu7YwBWa98XONsDOBIpfyhvsAF3bM
GqiYAKpkp/RQZ3+04buofQDgl3OCrRZLtXe1KugI4ATbLW2Zsa1i36ip/+KU6TAN
CfRzSS2cEOnAGFfEmn60CfwV6pSyYmNDNKtxOI4NIOhv/CP8LMjoMQvL8Vftygce
OKZWjsBSqWyzjQPyStKGpp1SnbLb5kb3yLqTXUs2BuIutcfJQUtt7jghDVDuV11r
7TeZiIuJA7CaztPiOhjHmQhwr4e5ARRlIfYqVlXjlgh4emb8l0LDYSK0HTdjEfKb
Rx9NPav+tKKNfviAwUQSA17dVAn5piapgI5U9ZDwSRvsozaPgM5qM/szMpUR/yrm
Ddmr52Qw9oAtL9RvGvzkTd84Zmo+s4t+XY9Nup9x5O+LwwMs0RrojT0uZMmdlGCo
fPHvZm95qiHLF+7h3QkCSQn9XAFjbUzmSiarqu5S8SgFeXU9L38OB3fDk92Z5K6b
dIjsMgHeoSsNKKwA36x96sGtZUwteccThRXlPY3IhOU0t8QWrrOOuVMwt3S8fxzs
O0xg6xMVRqEkG5wVzv5IIH4HibezIUBa9q4SBzUjGay7Xr69yZNXxoYdhHAJMCPO
IUQH6y+ryhORuPDtGFzr8kkNPcWrs5CS5E7p33BUHOEyxmn+mut/w8eTSOuKsjcS
0EntYj6EL0BrLPMaukgHLTBBOEJZOZQBDBSIPkal1h0jWz+FuxxhijpdXgTmB99r
TDrlT6rIi5YRIIt6vRuWpJgB1EZgcq7GJNUjCH452VrnFOmniTubWIfK9ZTWotxZ
16WFLL9jGBopVO8GEgKCXIyPBqXrCCWvp1EvZd0+bFgK13N2cgiiGTvuC6TQlmZv
W325EmUGlrAALsgkw1DgJP8F50noSfhzNlONIe1Yv1qwoAzuJx5uP8OyVlzrX48v
YA9sy+NKBB2u/i/r+YCIPlfK1a279ds8lrPwmLVXZ9HCKOCwcm8v/ImXleyJFLt8
HE+1g73pm6MtVUhzH8ti/WvafYfjeFusx1hn+rybtY3ZwTzYwaF2Fmq52pg8phXZ
o8vTQvZY51FNFdPgOQV/RpulfD+QMPAyD78Nb8waODMJUoly/SFSkIdsTRPmEIAR
X9DkJGVnKSTfjupRYjVvpvYkpz8vy0GjGKbCRshu/WYZD3vW/d9fHvjVGQSVa/Av
y6b6pVstiYNqxj+ipAUJEodqyfycAT5TNDe1rJqWSe3u6ik/DkbGLAe+gBsnxdrw
TPhyQgU2xiyXxbkd0jTcqqMpw2eNNF8cv1chMUp1LUoA1ZL+qNkhXUcqjcWHi/r4
kPkxc5u3NP7RJesH6HH120hup6TxmyjnQZkT4veSvqLyQWbCeeHqyctiGRcry2+E
TPej8MVDYayoyJFAEVItBJ47f7jBiMSkLJzmpJnU4Hkovts6aynIhmFUafnLtdwV
RJ8bivm4zqCo02Ob3apM6slHdGi7FccbtyfsyXaLa9faYa2daX8V6sYwuWgcsyzO
RwS+inmN9Kn+GVGAIbEHhjYry9GXtEgalB4bFfo+rFizDBhDWtelORvuNxsXyyS5
HUsC4Eg7eW1smx3m3ETBeK5WvG15MbtSwi3cFu+G+a9mGzOaANjIe3Mlv48LNRHL
m3c3qMoQ/L5sVfRbzt68BfF573pg1c+D8zb1W0hHrKmFSkKelOeDKEa8+8CUxnRR
TmTFg/YYKVISZv43w6Q11pBUqGANcjpp8MbMoiknqv0xtUJHkOYM3xjdOcWfn/iU
xf6KX1ecLqgGzdUVHTI1R13eNat8HgRbiFUmvvbtdQYC8E9Ul4rgyJkPjt5DbUvZ
jHhGjlJJfc5H3awcU6yNRSBZhHBga5EPJEayyJIHP4qdiEUGISvzb1kU/3DnpRjm
gCApi9CBsx8AyCZaHz6nTCPzgfMXJVADbN/ZAp/01uHbrDAOFXZbAl98DC5qW1PP
2OjWhAfCYTqqJxJ7PU2GJ8A8O8nuGkwHgXw30tGXLQFwp0g7xxY6ZOhiGP0FS6lV
MyVDNoo8eJdBL1RnyG1ku8Pq69UqRVQwZRBEsTyApQZYtLbQUlaM9q5vPf0V0Vw9
djGeha1+9XamOXcg1flrgIiWpAI965MjH8ncaWmZnWMRM1k8vAkL3IY5amd4T/JS
XqZkQe6yRabOXZYIvn2SUEXYscgpfP84G668o33y8X7/5gE/fkcXa0ln2Ixe6eFy
4PwImb8yU1D+fNkVQZeUGCvKHSobKLV4YTNXofLiQmcrPeVMg+7k9RMxjxdXOksb
CsQBWgDZn0/byaQSLbxBnTn5D3HTsfrK5KAz2YRUpcHrq132Zf3Zfx4PNOCWZr7/
XA+d1duhXipCZNj3eOXfuM+pq6zk41MG+h0VNakT9f+1oXRJZ7FUPBNLa6xNhege
FH/oWEvngzipFHnvz/4z9BIGkC27NY9RYw11SwwQ876yoGNo4nZ/P4ZXlSYAqXA7
PSbDZVakaff6UmVcQMrlXjFn88puUA53HvweHUn5ynAZeGbKsWAFlhrC/5kuRzTh
97Xb1P10Ie/BDq+ZvcHRI4kpJ9+RytE8oD1CFTsH4SJgolYUjrOJga9jyw963wbG
/dIs0CoqOtbWlALHVvkUb5NMUHB9K2/9DtpnZnWRlSiDGi2d4HfwK6lHlZ/r1yPh
UCCpSpz4toXZ1r8UMYNTXY+hPwY61hNwLd1xXOhSbnwm8Yvge/cgbQWASi5rc5JW
BwTj2rtEN1UBXKqo+u72DjBHwRYgTi21xIGQQiEK5jMCkIQSrYPL3ugFCmG0kVNh
VrrtuOs2TL0S1CFU7xS4Nx0WfKXZiD2c7YegEnlFOHPNYsemrkuoZpQEwEiyRGWO
6E0axVo9tzF6svPT39IIStaUBmV4JRtmKW3TPRkxPWEih0eiVw2bVhAr2Fdbt9I+
Ch6O7d6lsFQ53IkdlsgrDLQ45qStifBkaKHwZz8xoxUnBOVRC8egbcKpVTal8kzf
HOzjxrvVXFmldpIKJeAgjjvlacpEgBBWmfVLTH4lb0rJ/43tzkgEdqGrmEHfowsh
9sYej1mEelZCDHZAwBVaeiFxOJy8kgtQwBftbw6RyHJE0iZ1U5/IdRYz2PeLjCOq
AmWKmKcpRL7F5Y0zl2M4oGaXrE9QJylu+gOvy/LXsdluWboWsCFiS0y1b5xthlQg
GPpAVPPdH7mF69crMh2Ehz21xgM8aAVZJJaDO6IzFjhEs+scPqJkM7BNBAEkKYGY
wDVmSd2NVkOYq1tW9D8v8SkR8EHtnmV02a7oE/l70zvcOPwz4jAx3Qi/+WRBaLP3
MZool/8xexr7G8LUTz36b/B97dAK8id/Dn6If5OQQRiGrXBS7CDiRx7RVdQS0egD
u+8fBTTU3VHJ2BxdIMranOXeh92ntotCs+6yOkeRDRUQi2KXZ8nOLMO7+nsmVPS0
0xlkUq9DHK8qmrbWmcMxaEirYnBB8JeiMLbrRuhnI/G1ADqhQ8qjJ3p6MaE2/5r7
0RzSmkjh2sE/ZD8BHGpbGlOKx/S0Lzo8gwLr6T/mVD/Ebe+RZaGVHkFVVJzF+LQO
Bb77JknQSCBdIv6yVNZNSUeqYAE/4UG/heJ2Oh/DPz2OSapGuL6eMSLULV/vCRV7
vVm3TGvqW082AjFsHdTqV4KFOtzVnSaD2lFkxBvkwQhhDH8gvctVBpB6eEzEbl+A
ONV0lqfyCN8UMHWjqlZhW8ApjmxaFPzh39eU5+zr6zCa4WjA/zr4IcKFxN+s+vP0
lkMQTyKlb3D0oBLrtJ7V6A+uNImfhjT9K2dslUHAKip754W4oh6OI7j3lCwzZ8bv
d3MTC/z2tI9CLbOe3v5cuXDA4brBj0a4v3HZYrwCKPBxhZKsL8umSJ6vmAZyM9L9
BQkmSJ3nyPjyuSiq4O04/Gi7iLJSKOL3v6CPmia0B8vclMUlz5haET4VxF6Q1s9R
I+TeeJU2L3e/K6/0vCwMTGCpGSb1JiZZ1lFcj+p4A0jzp6z38CRP7q5Awpc9JYIc
6tK08BICEkZCRSrUrWvlsy8ZYZCQzBKndl+I+aH+nISFIhQWOtccSndyQIGp0bkv
hLYOJRRSLxQcvlzMl2vvwnNYMlj0FoTdjbziUj6e75Tsl/6o/b8Br1sLDnc/z1Ru
6chCVTSD9FxNAfR31nDFc42FfEyFDY1+nsmhkWb5WSzqFybkr3qZ5qeO7RDmiVkM
ZvKJsS+5xHrTadbOAgqcdyryhH1oCP9Wy+wJcxVpDagqU+AylMVbNPhPAra9jrLe
xsQYAfBB9xPgOIl/l+q3jmFQstEG+mcd33lLXk1ghxwbXf59DIcJzbxnARnBG6r7
rAOOafT2gL56dTCMfpd4nCmKJwmeflZU/rfONxJCZyR5XzOMSPvasfXBjMKuRnWc
iaccmMKZuufmc3TtG8tN23THpV+39kFxWQ71O+QCzF3beYgo9++DDR85Teb+Bfh8
EExmzqd0lWEC6NKkvEbK2lq9KRlASevFjRjoMVSG4TdbWYpGMouA+IRgW7lfLEoT
E0NtIRyEm/C6VIWzebmhS39pt7SL+oWrWUs4zGhBXA018h94iaksIO2+qxNMf+Ho
dyRC6xwLTi4uMktJS44GHP8nhEwqam1xtXyE27Ge5+hVgMov6Et/ytM3UtnkcDKD
CyCHZuYR2gFLPCOYfo0djpEh85P9EIImsdWHw/Gw8h7+4JyTspHKdIRIjIFs+VXM
qOzoCifNxTkmGvU7uufNKmDYiPpuxTM295TTFD9cmzvRyuCMEKEw2XZEbYl+xjF5
+NrWywxEHM2OPziyCQA6Ga5xgbmrYC1gvkThUM5r+2t0Xk4mRsmTzxqJ31KqPdzM
60eeh04iZ4dlcVHrucEfLrVWzQmjVvMIy23mR3/uLjJD822t6hRIG4QQMz9jrm9C
FnS2myGXzUlOGWSjUcBMM1gA9F2kDUgCz+zhRf72DsqBWY5ptL9+lD8NSSTymZTM
rI637f/pYqjSqM+Ykc6ydMK2g89a+RMmkjI+O5voZTgA0gKlSCSjoQYSAZSEvTNE
qYeTlJA/MOkgOUX0Ftvegm5ukAlN8yZCRz062FyIg5+YjRLu1ikIRPd7cgmE/KEq
fRNAk1VMIDgZ4fa+yn5/4iMJZRVLAmMPb9faShx9Pr6MgcOgThQ8ZLiwyXTGc6vy
xfCdDTsw6LdupCG3wdaT3JSrCXlUMQWnYrjQBPKU9pwVovbl8Y/fXMvM5SGgAKV8
XrwuiZF2/xLjzYmW4RxNFqz9ptTb2B6g+P3jS4TYEVpc1Y4AnSX/U/tULj7d3Ykp
WFG27xr5FkxuIf0wJCh1flsct53x0BL/iH0RlJw+rT+IOlIk+gYeKDosdPL36lsK
veMhTqF8y4ybZoKwbBctH5J6FekodfFAQtz/jV6glfZWe8CXNRQ2wRq/WaCmVjd+
Cb5wOJPYxHWIIWKYievI9oWRD9KhReMuL2tu5fCMaLbFi3ZlQIwhlyT5kYoDIzOm
p/5VyYpeBAYnfFe5qYPlGvReAB7UXUkCuqFOM89lK4M0Pz6G8tIdvCn8kbddiK5x
btCt3eTyxZsv1w33bximK56B5JzkgPssJMTFRjZpdkXxvwYmwwGY+IS0didy7PUb
QvknY9+6z6tIoLtXgPcKTE8/b1ryxTWPL7W9kiXP6EMC3LR+m8+TOdZr4RuiLXC8
Al5ig8Df6crLuHKtzu9VizxOZg9vlpSx4AdBnp4VUAJyqaqsuDwG/gMSIRQDGCuc
EAn0lrGiDOLv/j3gKqClVT8DKj5Oh7OTLSeLhfylyUSCTpTjs0hyJJCSjvz04FL0
nnPhPL10mrmO30OACKvDvR7Fo2mH7L+lpU9WQAbAyJAAVfWdrkyAWSP5MsmUS1V8
el8lPydzijBGCpc8JsjPdpWyLZg0y/m5ktSknw/veTJR6H4WEqdevBz4K4LNUGfT
8uP3BEJR4MfSREUGWuGv8zxz6moSmGej6TtVbyh5wEDA1B6qOkKauIDI3JGGUq1m
mNZqmP1vjBEnJOu8dGvp9D+wzbVsr8WAvlp3tTps6HAmzVNUaFZrChkmExFNPign
cofntAlNn4pquwlLAEzenIMvMK9x4eCVQxW1PqcN7NBDBVgI6zjjE1HoYLSumEOV
4wL9VwQtkF2PF9DJ2daOV/a9QEmGB2sSO7JeoSIAwTV90P00QxDYEiGOaoL7XS5Y
a0WmPrBeGXtkFCMz9xrMNXjCnLL3qWsmSkZ7SCC6XIqTCJHGwLZUc9/e8gP2As6b
QEWLUHcDmkwUBRVP8NIp4aUMSlvWb/UfRWX0dwvSZh/4MLEx5srZ8wzzIPyeNXYZ
ONiQwae8LxPRylYfSoHKbqKbPfGFQMvcb0JmJn32IyedKUYlIU2F2wtgFk0iJ+zB
nlDtXkvVyqiDhtUCiUJ4Zorheowhw5u5LGgHrzfgPeqN1+2t17uZM+yN5+YEdY5/
vxrvOFT5C9jDt+3I0h6xvKKLbRQWX+5N658eq/df6GJzmG2PimOoOC/qjlXvAn/K
sehTcPW5GfakqCOA9VEDleYjLP2V6n5zaaZgjrgNmwrq4i+XKMTKBGIC/eA/lovg
In9qsPWTAkOw0bAhTkqcPEMybnPpvZG8YeLad2Z6hmS+w3AZJFroPsw7czJovkuP
j8zWtcnJD3iVRVnlZXmYDaWqeJ0AD1hkBlD9s5IOE5covQTLYwQjhyJ8B8/fcfEt
zNFzOtRnPVI0/vrSKiwMaEkhCiuwmujpgk7Amc891SQ28+hDYbXfaV5YwbWqtN4V
WjPhKJjk1dlErhZXn27NaXb5PxvVbI5ZKGHHvSLhkmM9lm8TP54zaELehliA57Aw
73kWeDLrlwo63fg4R6KBLGgU+UrcRDV26GtEPrFpFoL2gbPaj1hk48oMStK1ASG5
dVXfUH1hcxlHGnzIi2f10I6N+4qkJ2hkgxrCYADgnTp8+37NbGvv8Zjc/QZAZz6p
q8/l34+DmRnoN2fBBcZ47NInJLxp5SkmIg/HC4YQTFjTRlbyYnR+VSMsGipmfZ1w
k1pDBeru81/5IS74cldexiTohyNUroyfhyxXymIs8H0jZRwp3J9Yjq9eb5LFltyx
Dkdqcfx7oNW726B+gxYYPCHDlJwVN508xqW2sNxTjRckcJUhybAFZ2ZJNSfvTUAB
TEGYjJTFqZTBcF+wCcKamm3hs0dZjL7B0cb8hqdngI+UVUfBReVpTWLp4GpWCJz7
acKqIX3Ay89bbilN4vQMo+O354+vFKF9s7au1HCJ22c5wX534QwRi0mJnOhjCSNN
r1YvwtgJewwpqZbdtQLhcOi8CJtILYXQe17nroWyYCgJWtNpSZY4O1mLT8Y8kimP
WI3ZThWTHXeO1y7+A/L8L1DWdFAVMjL8FaNwxlDmfq/+Y/fP2Kp22hg09/9+LsDs
YDG4Y9pyfxdCoKxBCNpBRNY0hSOeuw5LKI/oo0/+mEjl7RLrAu2L1hYHjAWk9XXh
tUhfXBgBPXgDqzLAcMugVodPY26PAwvnt99xJyIaEXYHJSK56A4gw+5sxiJgHsEQ
T9u/fwslIcUGWkkrJTwJYbRa/btQgrHzEEeXvc0rjXsk1flondRu5ED8O+hYVXQV
B3OFDi0/BfaqN4eUhiMDX9AIgghT9rydYHXuaX01rkQeMx5GUA8ZH2iBASECoVfi
Mi7XjFXDbM4NkedtzQJAJIcMcdFf7z4/aiCQdsjqOcP1LGVgwYeThy21jJ3N0zVa
cAn584IQNZQ1+KQX6ND91CZcO6Z2nJ41zhwdDvfJcViX2cL/hzHjVz/5ebGr98RT
VBBYBrWkk5xCAveIbHYTxKe5laxSdcacKHSUdx+ypPVzVAygEMuF6Raxp7DcqcMl
JfGppZ5qsHT2ub469ru8cflfskHXVGYVyJOLKBau8HguVq0RcOvo68E/nUi4BqLi
GL16Voqp6HmH47Bs3C4M13++38cN6+0pzTJD78c1/marG3YIsN60xhGiCIU0y/wQ
2v3twzudcd6SO3mf4rspmM/s4mppeY7QVT2zHkbXiXMk5igUVVfGszVcRQEmc4zV
yEgk5vbos5sKkHvkT4BL5QCf54uTmGPJUnKLAdf8fKWGwPbJPhT6NtokWFYfhlt6
iqW47BVrEfSxrYAu6oAvUEjz7BrMp4k2Q1HqnsvfJaJSjupKsvDLz05eY1DA+oCd
QGRAV40klJaa55s40ZJxaqtNZP79gN9YC86Z5jaI5QGXwb7aO6NFdzwVrl5jQ4DJ
cIiSu+OHZHQ5wevn6IiNLphbeav0a+o9GlyQjIYMmyP0n7/6F54ZjtIq/GW2stG8
+t/nEtNS9F8T/WfXjGOY/Tvze6YENaetjjA5LX0Nx35Iw6dPxFMfdyLOwjp1cMh+
5OYMrgZ8gGueWP+khaBt4KkbCgi1aojaIjW3pH1nSdCYy6DroxqZ/jEtLJtTgxHc
x/Upjh/gkS35P2754vxNZiZIqufESM24p1TdnAmLtwY09jufLoGbVSEFArmsYhjx
VDTaP+aIuSTPLZRIuYwxdzyhUc/qIos5AE6Ac+Lg74CnoflPa407pSKkAJCF0qmz
APlQzHskk1dG4X31oj+kLY18V7XJEBWqtxe9InOZcEsYzeCE6yLY71BeBBSTvEDb
WyG4wo/YaN0MZ9LDDuHSel0/QXCN6LnsZyNGcEtELl9tCb0YXe1rrjqMYBNgVr5K
ARAtKGZSpwwmQsayiRTeEXI/DDOHuJ/vFMe+V7WS8zp5VhiX8zH3foy+Vrsg7k7d
DQoraeIDrmhZ86l9LxkmZKc6MWpBrSTpSKlfGdwZoKtGi84TZtyNz8iFojXtzQDK
JihqVKk8IWiyUBqR4PkZ1EP4c5VMJ4+CeHj1g9A5LP66OEiLN/yNBtmxn+PnBBsX
JrsEphAK9DKyhyfchv7eE4oWKIrz/NwpxKilVwFp2cFkNHfZiY4YWIUORGEoQfYX
PgCdFPTJodUzJcq3Is85Mi8tzs3zvboi4Cb7bO+gVJwPmJOopVxConL+8S7NTVmC
6ODSSg3Jsn9bbZytY8gHzPyKAQc3LGAFfCiItFnel3oJmtIGPskAW50wBsB/qe/A
+RlE6RBac1vQva/d2iJE4mISG1HAY9D8CjNKnkd/2JbcFEZfAhoEC9wwXgy6LPkC
naDW0wIqvH+3dh7CyJeQkG0oRdeHDzAYAP9iwQay2pGX7xmuxkau9YGQczuS3VnV
uPmoEaJBbLDa8n+GJcN1CuScw9SubdeDW4U74nioLjZj4LMUc+gRxlrcJZW7Tzm5
LbyWY+BvE/zcbLK+VVa6XiypphqH6E4kuJrwPwhLubopKnR6JVqrL8ToYXgwBl38
24SiNAOjrdBbZ39yyEDwksQ12jhTmErAR80ZvdwfSdDTORYTgrVnNwImBIVFYWaT
NO8L+u+wA/DFrVCWfKirGbwGRMqy1D7PconpoXMo+PmIvd/kzusvGLvLtGm3diMG
ErYI7+HIKpyOq6zBH+lR1Gfd0tmT0UWu1S/LxWuBxOixtE/uaDxutY1kQJdfgozO
4cizgNt0uKwVEu/eY0k8TTxrAAZ7c+52ifcvESVjXTQCGlwxvoSzb/4rK/j5kWWC
9JZduxOqvul5gi46sCUzhQKcjzL9A1btgMVsgMVuibbjZfROmKRsm68haWpT/xzh
RmFasQz1DFYha0qwGCcD/8HmYR+bcWW+CIwu2fhsfTbv9+bH3fvlGPeWxxh4scUt
ICuRj6+STI80f3EcFLw/iCsrq0ZqafRY9XwjNo2Y8hFU5MrXFWyovs1x6Oqehtk1
hcBc3oC9Nss4Vcp5pHwPgGzwalLQyHo2c9Mvz9JJcWTVXvsW9w4RdkntYKu1ie1z
/fEJZAgxCb94EIOVp2eaTx6acFC7jDeXb/wlB8g1LRtSK3cisSvDQmq02dglUwXL
nwIjMpKHq6l0urSROwLySXT4bXYwSorfJ9piffZThMQGcl6KUcf7UcPe3d7UXnsI
lkFX1ah+C/aiegXYdLgm16lYZCn7MnVflMQyMg+daVfxSOIM3u/yqrkWekMTS2U3
/+m1v+Q6FP0lycRWZ+BlQz/gtlY29HavqJj2YXElJjzCpbaODjaXJpOU9Mgbvn3r
ie/QY4+WF0PlzOrQP4kz5cz/KWQfY/jT+FaBvi61pY72Gll97JYUo8EXOdmFLecp
wl77HdQ6Kz7zFofNtKOztcoS9q0WDvc2oDXT+8xNa2TFv2ZWuByWaY1gYzHT5qn9
nnCg0oHQl5ElhApe9KpWOXsdkgZ3ZMJ77Ec2DJSoV7Hd+4phCOFlwZqREOm/rptq
yC/Uh+dwVG/Cujipz64QZjPN2z29k6ieR7oW9qs/7Kl9SJ4nJBOglOO4/EQyvTjn
lAmkO5P5ljxGLDRByII7H7tZLEKNU4CS9h8/nlchgdh86YPIi+XWRyBo8dvUmgdu
1OTrcxOtBjjn39D5hThMM2R5fG8bfm1Jpqf0gwqc2xQ66PhCrw3gBNQ2xUaN3UAh
wUJq6mvbPqC+LHMOhBLn63GyaLbnAjKD54CMJqFRJVlW55rwciXvK1MV/2ogbYQg
ONzYPaat/iPQU68b4cQ8NPtenYKBQutVCIODT6S/+UYRdCX+ZAOny6Usfd9IOtgk
b4Q3FuCCvAFKkSRSzqelb7Mx+IA1EEw2I+LpNnD7tXuUn5ODugg91kyscNEohxDs
W//JwdQGP0Elfk2iTM9wAZPOBIuYNJz/flsP8sDpLs1unadiMSiN7EdH9m5gdd/S
e5Q9oaSdXkkiVb65ZLer8d0K4aqA9sF7WJTjqSOlv8BmPe2gY3+8C91gqy4R6SbC
Q2dMHkw9vuXykpAwaIowvbuJ3yBhWINdsn6SntYUo/yEuHTSA8czGfTEl+N2PUYZ
aDAYhUZpW0rpEAlvAhd5YIiQoNX7iHgn7qIWypBUh3+HtmJNN4DNOglerHGGyh9a
6CMqyVedGB20FnH3L9DjcW2AKUnkmasLyXrPETxcuMWweoBEHLoCu9tmoQEG2gvm
BcpMw93NWqjkByMj7Lh1TJoJGcZ6H4QHnd99DGPhaD0BU9SKGz7GrRgCbC8QgV2f
gQ9V1g5C5vC11mA1NR10KYQ9JvZ+9VcyywvExUsh3mM=
`protect END_PROTECTED
