`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
huFcvWttgtMuzQNivEvC+W/Jk68NkvQmoxvCO/rMUsNXvPu5+Ndku9wJVE/JO1sJ
/ao6qP0xGjdaQFS6mffwzvGDJHCYVXM81Xwiez4GfD5/xIqxBuh2ABVa7JGKzztg
D5CAn2RH6fs/9URT1LMKTTTRFPE8Mg2gGEd3/F5lHbhDz71CZEn1leUs1dcNvAzI
q9u+yo4dqtUrFNlVgQBZRR91rC75YBSkTTDcA3PSPmv68MwUDx/y7OFxmNbEu1jt
ruhZO9Bpw/muizKmSVX8e3dVIGWOrNL3VjcNQBbwNLZtwyuIyDD5z1tHnQ41VSM+
WCQSss5UpfAjMD8UWnR0t36UkxN5j0zRUUcTad8TaOa6jIuUpGkGKjwNz8y1aH/j
TsjJPDllTm+Cg4x3bBIXzVnvkpYzGH7Snr9/VVbxg4Wf7zxZO7qaIoVKWwVSBEz2
3I2IoODSxv75IahoVsOJygww/tYQkzrcOcU3zHnAcw0rvUbw0PCkcOV1ixgZJgxi
scPSsleaRAMDF/zAjlqahOE7jhSHgA7gfz2Rekr7js47QlOVYYDZEwN4095Zivjp
HipNWL0879bvwQtK9xHhHsuWxtriO8gMFYR5Cg5qrtZY7kY2xITHBKddGdkBS3ei
fMdHXk88hNozBjJJkwpam17G4JCSRt8pUm3GoGVbsgecMTDjONo3J/m3SmmXDaXj
8QCwprdKqsfU6YlE4/KPSDXa4151EalA745WhTHgd9G/OhrPy/sTbhu0Z6lUNgQU
nai+VpMZgbq4Mq6rtGqkZ1f+/PP9rtWOtmn46Hu1PgBNkpEnhWAbzp10QQqcAPe5
nE32BXhUOvZjBGNMRcca2jMf6hNI9O2wokIRLtfWqqa4tTljlEqFYwUmtn+PSIv2
vZBH8PegW/mNMldrzfxRJzxVn/NDBWqLDCkv3KU2JHQboUSC6IgICnWzCnDzMIhA
kZaKzBA/tLkM9DyDUbcjhAlkd3SjyuPOPwE+zGtmZUGQDtRMg1KNsa7S0HK+AHRw
fJEHlkqUwXNU0xDLPvtxgH0rDzOzLYFrKmvpmZZxb/64sHJe9MOmX7FT8scwVe/7
+z3LtT3OkppEeiV0BH4P9lULFf6GfYB7Qdi8X1sSg1H1fpbLRgTDSnKahEfM3M0N
xBx3UiSbD07UBY7+OEB8DnOcEKEZ/8dDVFMh9XYDvVy5LrDpj3u+WKIGLQQd6v6v
CijJEwe7xJzgkXch7Q9y1bbaKnTOJltgFwwrsNNYHmFfZWpB2w1y35c2G0sINna3
CrKoTo6f7n9iaWHN3FbUJXWNdXD6u1HEyUIgURoUaJC4yW/zhkcfCEwn3ArmAba4
2dSg2OsXQYVuPraIdFktP9+32QTyVAdIarSZsAZrv0/pPUjjY1kSi901HwZH0wkq
cN1phYrNdn4cx3COk+ubvchNI3xgi0ajRSek9En4TJE/Pq5huRrhIQGhwbVYYc4j
xCna1RFJW65hJvm1Rkuxk7ZW7tHeeC0Ww/WweLDPVd92D7Pnq7ok68GZ9wtKlTVh
Ps5iBUEbxFi7KO8oel8Tjnc7mrywCdOoi2jpBOo3+SD+/NBVxvKBPqgNInjp92wK
y0shuPecnL7199P9bSYnYpS5SXBqlsOnfWixL4yVNlV7dZMq5/yFb9iYlwaJgKxs
P4gu+EQlNKOzac96J3QcEqv0AbGS3gOvjZb7PRHJPptOiNz1snBpw96dv4XtNQNH
P40CUWxKPMf6XizhxM1kqgIODNZVSgFN9PXBJ5C9SaTqrT2ETOwp0Q2kJ/z7pu2A
xh6DdFq6FzCQbIYnr1JkhGZ3CxPtApZKZzWLe8oDOtBHDcJ2OPMGpnw3Fqs6z5lL
A6JMpGs1VYrI3poW7VHyhvKVHaUx8/SXE3gF26gWo73QAAPweJeS3NFKo6YaGHFj
TzuK2GRjB0wSyWErk0BubSR0gK6Jfrh9vZfLcmB2fI9MATtj6HmTDye0VLL2N+Bf
cXTjxAEAU3bKSpjTdY9I8sA92seyxSKz82z1fsu65/ICnAPpHE8VUiQha60Fsr5j
GGypAX1TCtT77PWayakNbawgFdGWHwDxh7Ej79u5OSxYtYg5fpl1QwNLoHcDeN6F
iHkDZtf/58lI9zv63GxuqfgTieJZRYiUa5sdsUAIy+mbZCnJf+Hu6fq+DT22KazY
w9aOFenKMBF5gQlcVl19Fh3eBZ7GTMgdk6VTf1KeRa9+VFSOdovT9BtI0cBxCUCf
wNraBwZjgsGwMDMk6/FqQw13GUu8ZDEsMdLw6cl4At4HshKTDywCA5f+TV/3EjZA
xsocTilA1rCryH0pzZxwcC6kd+Cfoz6UGwlxNOetnK4BUrUF393mp2BPYhoe4OFp
XWxh+wibetkMtvmpAMAq1z+/QQzGu8DRLGOqbBpo2EYizyJiPItNwMn0o7Sb2wQ9
qj20nCR0ObjiKwQ+MQ6psiXBKO4kTWpcBAVX6Icgpb1tvI+BE6hr2TQ4QRG80jJ5
eBTPmLgO3p6rCSXo7RKRN/8jNjr3S1GO/Gnf8JTVEBrwqXhYwe9wO5zT2zyHXkSe
7b6LgGQR3iJ/jv7n1DrZ+1suoFXhoKPm1e02GJG17FnNwtLnnCobk6JQfC2ll8T7
mul/BeykicNu+c/Emz4Q0WrtGiMGg7fT6XEJtntx+sagkxKXycPPYEOT1evoMbnr
m9QPT8e45aRqBQwHUD4B+0veNzSoBupVJ4NCU6my6jypFPXAyTDu+Mbzw7DuZ6Em
FTMLIbGhCbChI3hvDIJsXEuX2GU7y1vaSO5CMCi0kSiswJ0wyGoYgWD//CsCHYQH
WN71SFjyXt4URKskQUm8QjDB8XhlKCf2XwjvxAtTfHc5RZaxozZyV90fOjV55j7k
eH/bJzsd96wKYUdve8nNMN+ZBCPG6r/Ldw42V+DeUBBZRDaxrrBGhs/V4svu/rtJ
YhWABpVETP8Uux+L5PnZVJXpMaOrdq/sTpBl7Q9JsrQhSQPMKOwK8TjH+FAyG6eC
Z8llCzCf+ax1M5PhZppNmdyi128Hwb8iuMCPFUNeRbBz4i73MD0Uq4F5Xl1mwKHb
rx3jyM1DIXaWlnUwP5sdMUSpyZhor+QjJlqPqjf6vwGBbgFXXEFpBL0/H56KTudD
TLo5Yi9W1ybsQv12l1LKA5HjxVndZpFOLELnedR2uvVbSqeM3fe8vMrubxKQpEDv
InYYcdnqYVDrBHS8P9EMlHXNkFHINS+fKWJaM/e3b+yNQWAzmgjmIrcU7DUsAFKi
YR1S+/LgpXNvy2qAMy1zhVtbEzm6keH7u1PRZrrlSYY=
`protect END_PROTECTED
