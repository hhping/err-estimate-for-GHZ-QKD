`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZW5TXpL/IGB1evVQQYQt6okOr+YGRvXx3yGm+umgB6kqqJbX2YorhkMgfLBb1Za
UxDgzzDqtRguVQP5g4+WC9jSiNLTeefelrcwmswXcoT67987L+8Jv6920/MGXxpa
Xhl4bdiaU9mAG3xiECjXA+nxvsHEZFxqQXHR5YLQc/8L8OgpIdD83lcB6m5lnS2F
uH/4c/Fja5ATJ1ZSuuCjUiKsgYdTwuBlBfIgdLZ+dLF90TsGWt/e1U5+VVxS4wuF
ZsZV4vUvqwrIzvOiFeq5FMZ7Os87+1iydM72bTaCcmaWC5fleNZudhSP6hTGYPjc
uZ9UUxuyJouOZSRzKH5y5gQp49bCFQj1tdQwWQ03gt4HmzPCTOj4sYRfT/SlShlj
hj1N9OtUm5Rr2SOjcndPKlyDdwzxKo4nuBywau1AyMjkAL6PnKu89sbURxJfTO+/
gzfZezmHli1HgYIGxM9JssVpWdDqCQUWVvNpcFMRHO/yIBLbKXoJDG4xRSYso/Wg
rZyP3kpWxdcCS8vANx0WHvPU21B2OWhtYWR6ekx+JFElSEAiE5Gpkuf443XFx7ij
mSTdHwYtjHLVtH06Mg1iaIf2Xtv/eOvJPTOwic3nbgaFkBb5nG7AHNGyQvLBa3rU
cFsSLiUoU9tJEM8VgP8uTfydgXgPyuzQlXj2VwqIGrWXyVW68WZH8yr0YSlq1KMQ
RAfJnZ8BKiTRPg2DkNlzUuFYO5m39r/gkN6mJlBMiEmOo45YKT66dVAF0vNY79sn
2hgWLgJDuwyvr3ypuobxQGZDqYt2WkGHwv/oZXrvSuTZ4GN0ysqkHqyFH6I9KRAr
Roz+vqm3JltWeBYzIW6EQIMPCxCFfbrFIFo79slEoN1nnVadI0F8iHcraZLg0DNa
f8TgvIv8Rq2uzesV8eR3dAR16KIiNzX6bZCvmGaDdktuMLHdX8dccyP5x1bmfImN
+l/KJEkyYB0IYfxukWDkJq3Iw30v1PAriDLzhcJY7G/X8dfhS6TEXe1KH8SPhRpX
4R/snvJzHjFRmzHcAUC1OkRfAl9+uNfuapwVPt6AHLKWsXQxLqmcFhROq+8uOHxq
HZ0ni05X2wIejbai9CdHG2QzU6y92Bto8DSmg7fJJKAwK994RnIeJSDBkS/IMNGZ
o+vjOBp0TYt5EeUwvHem7dcLoRky2JP2o0IXVoh6IdIIHzVZAjEF8eqnZ7Jv0V9J
y+H3OgFtkDHD8YktlnzehyADkSmW5LpDowCPNaPSmWoFcfgDcPnPPRQbKog+H1hs
QKZvBTjUEcPbctPgWrnkNjcNJIIsvQ6JtNo48VRhdKJuT6g0xeEZpYKoXZlh3R8Z
FM43gnIzgl0YSFaKoB7zlM1jzsPlUrIRoBT2VbrWvI4V+gyv5BlFL4VArR4CKWWq
I7loYGFqeVMmqLFpl6IWekHJtULNwdhg65RsxMSScCSEGyt5eyCgKM8vanh6O+U3
G+L03LcK9qytXsx/SZZvTcN38urpQqUvLMTvXIBzKwTuKzVp2wkAhFPRa0u3vvkp
QEcH6S9DjuCU04JrwOnyUUYJM6wrrajeLxHHS/fwpWhiljXaUkC0fPqu39xnpZ2L
JxNZzX2+RDAjAt/hw+4+T+Yao0nqgNS6lfsr1e/NQezX4e1qK6buDDT2DV1CgC5U
pUdl6i1cIAAOjrj38hSUl3sXnCgR6sjLHDzF2+HS9giwHzBAhzBCOIxFdqm6Devx
IVszoGYoJc59OEH5IFsA18nda5BbnPlazBObQJDOEXHjaGR2qIAA3bEu6GfzTn1/
TAogP5msOkRgIWzHfiRU5fwr7jyg3sPYkrWomtSOSUkIDts51re+Kv7EpptcUrnp
lcnxM2zxbo7kERhNQxCIzFwSeBteZL48xzFe+z4MCtZwJaGs0lkFgtdrFHw2WfVM
KcBPz/+L90Bh59zrkick+7sbjubkkNdFXiTg2i2p93SdxAuPMzRUL0ir62dUlHWb
0YG/AoN7DnRquSnWZXT9mQg9MdLFjgPnPN/p5FQ1CciOzrqnb6yeVAIPB7srhkOC
10eviDJ6okG3I9fVZh5PaTbMz8WoVAEuTG5qzot1kJtM26fway+SODCdo5Uw8lEi
ei0QF0tdzsINan5qc3kT95bHGiapXUdSg/wkt2vueTNBu8BQJOmsplCA0am2Bkvo
IafjlDsNcGBwyjMaLI09qg6dw3tp5eygfl1WxHkBMbfRuHpU7qUWPakspPfWUUKm
nqHovtnNkNMAUy80NGHCqnpSFW8gonGL5h8F5/HR7L57Oox7hxks3KNVveef7n5J
6qO2RocBLBYGJOC/JJG92z0bhp7iwTRgRU+94o3d8tPc4cJJcRkZqSpb/hEkBEHo
59LDRx4f6ZgDkrTHXwNz3pH3YNfrfy/KTFAWc1aKLfQ63yuu6h0Plw++6hPisXFd
Dy5SsP7q2fzk2Q9/LwgwshFxmDrnf9qjPUisXoi0j0pYCD+ofssowSIH43pgsvC+
8iv12gy55QKevrR/LI9CDYTEdKRt32PqGhgx2XMytgtLHQeNJgENmsQn8APH9B5A
ufjX+DTLfxWg2u2b/iLd4DYQ4REUNNtmR9JvhHmYlrcDqC3MzdC8K5gY1pzYU7ib
jf5AsIMNClIv6ywSPE/z6jdCE/lajLSdE4LZoxnXyGm3R5/qTDOoso5RyWNuVzn6
qxSYaiE5AbXwXalmwB8o9pIeYBaqQserOznn99LrVE1IesiW5a0s7s1uVxucqFQy
LLfhxJkt4cAwpuIzLjXTJfEKZjJcTWKxicjVoMWX/PrcOoAfrQVn6vjSPTV8AKiQ
778YnL6lpDGW6BMJNWtiAa4+9lHNnjn6hVofGXP9WrVaQVexCw9CR5nD/hQOkE0K
uTITfDFUMbQXLXCkYXfPTZa3b71xYOs96uoWDZaz/qU5YJZhdPAOVZ2Ox7Aqi6U7
BcmaCDApCwo60oOIyrxyVcshx4FqFUrAPBxl9cgKPOm0MuJsRw/F9QVD0/Eftaw8
/HZ/oUERw+UBuiWboGefR3IczcfUdh2w7yhvY0MrI8L+AHds2RysJ55QSi9q2H5c
Zcq0dKtZbPQDDkVK7xyFpY3C9nXsBNEAbnpKHGQXsDHJWUUKegVoExmtxfaiVcO3
wWcTv2vXZG8o90W381R62WE7/s1mE3QFD0wtSouBL2DEwPVqrYlB0l+1DMs2CQiT
DYHCYimqgcLmMLxB4l1m7nmT4kpP0LGLycuzVGYU+1Bq8PZmQWC8W0CJyXmsnNvV
VhZBV87FPYio3A6BDVkinj0roxu1YAAhu8SJ2WRQNpo4Dgnuqcy9CLY2AV/NP3sX
VCoae/uS0uTRBaAvbXTJ0SB8TPCMEUMtNAhs7YCjxxt2HlJXwLeq3tkvmIzYyZF+
K56buD0Ovufx/uT7yYeLaFWdl4lePweoQH0jm3gyHliE5slqfGeRJqz1r10zGqba
xMF6oQyl1xXW5AMXK64sd/66kA2JU/E6eZR+hYqfkc95gg1BWL7nH90+FSdAtO2o
0X8KbpUqGiIOE+ZsqtS98zn3sDvSWKMTMcC5ZJ5oCphKwLcybHlei3hS4e037zzG
LK6xKYMVECfuwe3XToyI/CM5tLQupWZ2UAyCVHxeF/wdjF58FEv1IExotzrs6JqX
bsuCokzYaRfGw5nz5wITzXnS/hh0ZdChai7FvNo8HrKf+WeCoOrlKZEkL0t8wjnf
6izM+0J0uwLlb5stnuLPos/onj46sA+iAYaCwQS9bg3CCkFfgnlCj96dXrFbkPvI
hSYuSK7xZY5D+s/mo9s5P313yysqmu2WvIabEQz03schEnV8PvyVW9UM/TlB1elG
ChAytqdbUPe2uFNCMMZ9AM2nHjOpkJLK48DsLQLDGWhI4CEn1DE0UfUrElToKGsT
AZEUgJM3hyPt1sTR5TzwbNE5iUhksfMXTDLVLqo8v+Rr94agUldW4A+FSFhNEefJ
eq9oSUGl4wlP9yp0g7Wxa6R3kpgY25H043HFr0n/1aWJdAtlgAPvyu4KXnIteNWX
QSJjq8SxFPljweE/GNyQIvUJGs7/KNFLjvhuXyKOS1aA58N4lceCFoLT/oTHv9yE
`protect END_PROTECTED
