`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CfriLvtm7j4p+KDlXQMe7oHjlqLoSiJbYM1YY1Rf+JGEVkHvbklgyErrsYzXBmpG
ZYs8TyJW5LbuNgTfj9BuugtpRNlwWPkUoVbbifIMsGMkwSVS+loq5anlcRv5uxIE
Bi6r+rYBPgVi0Kozanb+19fK7fn1jjVkvCkOzRZ4SnN8FEG1E6VtBj4tyrPTZki7
MhImDCYfOJW/ouqTVRcJWxpF54+cNIoZiX+yDJiHRFBjzaz3bdOEm35CC1SaOcmG
x+Ja6majtbJhSZdKpx2RIJu2lCEdiBOKHYBjvZNB/NxmDccHuag0WBu+u/EY35M+
MwnOYcBUG+Tf9TS0+3rQaotuwcw8xYMNxKidYzKo8IRT92rLoEkhgSwsIaMs4MgL
bchmOFF4zEXNrDCyophQ45kbddHXi5It1Pm2NN0/rmM6nFZVd3KKJPE3bt66hNr1
3aDI70bA6JP1MsbpmfQPBQTjz7LWq00RYVy1786S+KjIGgTR0SluwcuZMcH4FN3E
kJYe1YBfz6R1aJfmZvD4TDG9l/6Kv0amR8tPa5/B95+TRHzpJV11eUgV0UgjJair
5op/H1Wfl0/jguLyrOV9dA==
`protect END_PROTECTED
