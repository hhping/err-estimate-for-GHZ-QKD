`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkfpSA/5trVvZy/fmHeN/SLl58pBw2HBQHhRr8MhwN2893012UWvP21aw6s0PwpU
VWvjAOPLTKckVvxgnVuB4AEvfRVKsfoHhyebzyUmGLC5BD/ycYVkyrm8C2BakGHR
eppZBPS+Lr14ncfDJi+PgA6B0Wb5RCdUrhP6Gn2g9kaaqhOy8p3I2b06Z/3o5Wra
r+FiYQHN8BftXQDCzu1duD8elx2uEyDAw+maNrehdIfnrCVQ5dsC94jHOPAXyd01
mvUtXiM3nUmkHfFLXeO4OR2dIbi65hzBPQLVoSZ5hD9wDOlwb5snGhAo19UXjp9V
5B9pPZEqec3O8YGMj7s5m4T0dyjGAKqy/SxSINhJPxrpaatRkSxHVBrOY3MDOAvB
rbG0oQMcu0M02A42ijqRhQ+pyxF0gUC/Dl9k8wFVjcT+436KqRbaKxgTy7wPW1fH
jAF/FYdXaG0Bz9EXIo/Jv0K2rc4dJ9azPADr+SmHWc1X1FdyIHc/6ifnbQwLPK2T
VzGQRLv6Cbbw/XUMNILJaBfLSqSc4GGl8gAiKAi3n7xYiP6JoboXbMtHrIyAgs3A
jHgnxwQFg6zXmo1xE8jRf7uLXdUALhQOnKoB0gu+9e6UPPEiMTZsErKIR62u7dZM
Y+j6OoGOtXGqv+e4on2q49OFK6hcfaZIGOBFEqyG006y01T/qD7z6RAtnakafnh5
GN3Vaqi3q3IMulOJypsuXqOFLWOEUOdVURLlOQ/lN/vXs+mvDn0ZbKo1jL42VryL
7Clnds2heYyNIsIevFbCCVNOC8xwbn7sXlXDMstQFlrK7GgfIWy3UFeWAEeR0ZXG
DN8G0bZVzMkhOxiRwI1XsRyw8VH9ghuTivy8fVaYTfK8u1/6Fbc2iNjjshJCGepl
xfOdXAdbzYeLAyu/q/B4xTXfz4E55dDdWlnTHjjRegOwBCb8oNNpeHV6l1z8FRKA
FhFuOXnTFMJrndas/v11L8GHP+GKpPWonaIa3yvaWX20n1chgMJgebRvriMdobCo
HsCrHOyJg3P6SiYpxw5rzYuNieESjWIa1W4MFzkkJimnZ8ko+dhrDVYuDtP1OlN3
aZ2iJEpt2SEjZ8m3USPDBw9nRnUkaAGeAvioEuF7aVPt0H358cu6NScMprll1VJg
m28q9/ceeb5x6ng5IvWANyiJxE/xSe7AMQrYJ8KBmR/yh6D72Es5XC4kaxUn546V
X1A5U6iXewgHVtahvyiUf/w0KifaQFckoEp/osT5R+MeDkYm98U0gr9Nrv3yseCC
n6yvM8UgsFcaYe2RrYOxQ+9rKBQ3fAExd8S12jS3BPPC916g6KH4wVQ58fRkQuc8
Bgr+Syjr0II9qGt0NxqXdyPELCbDnqhlQhQSNfaKJM5rYVvW8kk1Rxxc34tD4JO7
cMKCfG9mK4EBpCLgrcQ3jzn8xaoPNI1d2rCo0UNPHcpBeiDX/rDZA9F4UQlwCPg9
sSYGlYT5roqMLrR1+ENkU/U3gI2rhsQlWIfM7XI9XxUYrqnj+ZdQDSymBYtJw/L0
gks+kwfMKg4Sj1zdegcXOonwow6/wo3rPhSFv4vlPHmXp8y1FCWTVdY2+cgyGY+f
WXeqMEe7L2Mcc3IW14pfwie7r/Ix06CxEL2WPolZnc37HbX9cfKmx1Rpd2y5Nyk/
2IL68ddO9frejeHfAc1DyMfDV2t9a4Yg89a1QVbHYMWAT3rq++7qbPi7VpyLrE+E
eBjB1m7pxJs5hz13n1Qlq+DJxoRKIrWq2rRVaxLCEOaC+RiZTuFGnH/HmKDNsoF9
/cMG0xcBuO4mtaiohgE0gjWrN8Tm6LquRqmPMg/1AqbSMU+wtkR8tpXbAnAswgRt
FbMVU60Ueqplp9nNmtVl2kQQQBOc1aVlq84r1LtPTes9OXXHvkYPLF9NiPBseQbj
dNGq9eDqo8m5YTMte0cS3S4RCxYd1g0jGmo8Pvkwoush3hGHBr/SQoMiuu+CQbMZ
qRYhvTgY9j0oHBrZYj4dO+dFuouLz7oT8YdykdpaD0/IexVj7Ln2g1lf/BrXYj40
7Uo77dvXWL1TVc31JRBnxdLBBgPnl4oQNjaG/8J176ZVSnZ9VufGS+hMU9A5WNj2
Em2GP9nDWIPi/zlDjOysH2+jdaZzoX0fWIFGdeZboIKMfF//ghCztv4+KoPUA4Pp
ZepPdwGOzhnCliHSJr4V3Tf0Qllu0YGXCF8cb6zRUnPBFi+kuV1gLKuxs0YRyFil
TZkW8JXOh233sLghvFsBkA5G9sPFsRU0UzuHTr5dY1qolFIt9DclIRztRSFkkq0p
rzowmvrIyjBbRW8TdJzAuD8Kl6jDOgkv6cYA9zxDsh7k+uLVELtq80raiDQYp46V
tA8kXrnxf5+w8aVT0LYblkycR59+vc3VLEKAQoaRMLaPDB6gstJ0FJRBB1K57Jmf
SKt4Y1sZFUAyiTLLGmA24GapzaXDOJRRDaeyMGE7YAncZpOPffuReuSZI5n0gBkT
oSBQMrbdzf6i7dqAhPvBwTXQDlXncY7OX6krB8SSnInn/h1AMriz8UKybeHdg4mG
+OguXpAC8eMSRMKtIIWR+gMldxIntOaRB6PMVCqluVKIias16xgHuGciOewCxMrm
LCVZwbalu/gxh2GA6OEtHC5ldDmd4CtY2AKsGapjpBF7Gt+iefj6MuZYhC2DdD3Q
xeCR+7pfevZ7FK+gXxvqJU02QS987eqt+HaPq65k2B27Pq0CZjiZMqZhHecgJ+te
Dl1pPgAHtX7aPqrXzsuxR+gRuYhOh+W0icLmNY0vg/dr389g4LYlRSxkEZwo3aA3
cY11S5o13gv4RTJ2SE+42DPpjKILy4fS2J3bF5goNF8VXdKs1La1L223D6BKEXu5
roSqeRKfPF6ovuaBf8PVKKQRrq89O6r7VmSNmNtqRRECVZ+WnN1BkgzEDrdPkrrT
pnx98zgxxoZfcBPtfNzNiJ4yroKE+TV3E2qLT8QPeOQbjk/AZrERMxD08Wzx3LUp
wmSK9w+2rQ2Aqyj6NLBAOa6rVqZMy/6AbN3PoS64Lx915XHLJ7ohadaJ8HitpbK0
vAQtPz7Ga6MQwdz6VrEXH9d0U3VPJg45WzSUc/FuIX0=
`protect END_PROTECTED
