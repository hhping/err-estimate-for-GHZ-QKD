`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rK7ZUad3pazoUbJ4eNP2fof3yYCvYpuEHdWJKKNXGOTZrBvgG+FTfVIMoUaITm24
IcVpVa5BfMxuJlCAahkQz842Jnb/6IP9jeYaX+7oIZQFWkiWHSMv8AYoIO0W0iKw
NnPsK7PqlTdJqVWL3u4w5h8maIzwaurW1/M8SsMvTCiffCUtt+gvAahCkHLIPQ1I
7jRVomCSlkJkgb1ynbX5ipMnUMTMcrBpc3NChobvHxVVhzpjEK8zqJQ3BYiMVqWp
YOjjQx+4JbdX/Z9IkVryqKlOYYr/VJD7K5nmK3w5GoPOHcSP9y7R+7hh9eXJ2Ecf
odokGaCk3Amn7El0uY24Kx7qElwjTZQ6X5rgXxhox9vCRnIjtVvVGK3r0rtFvSu9
jrhZxrVExif5hXkvsxFQExpxiCVvBFDGtFzSXLr80gznYMN1gEcIfnGjI8f599b6
Z3WJ2N+GJH2SA2TN5tt1xuzq/MYI/V1PF7v/TRyv+/itVFN1GrpwtsZ2hcQZ9ehX
btv+Zbqb3hdSFQdzAJ/gONaUEeR0D7r5Z4y7QrO4mOgBx7nuwuS3dszVXcpw5z8Z
XtRK7YyC5eEE2VfmkTuC92Jx9EUeZ866Ku+l8gWcAu1N+cmFj6a3ZUT3eFes1f9t
Livff2L5EIMpl896Ne+/k4/Byj7sfLLF6M3I19RcoN+KbFWEmCiRPWVvEk19yG6y
SbADphYt43RL2SS1iBiVhu76S9qcDbvt/qhioXMZOO6akaJSrd5xJ4rWlLH+/Lv2
0SRLjdbJXjvN/SiQnrloPHe0fVfi/muok/ds07tqaJ5jdpoTYDLu9xPk7g8rVRTp
NQLIX7nT0bdcUqfUSXoZjLKXXOH7yE//2+olD9BYtlBDdKklgtpE2mBKmLlH2huF
b8hYMyPkQFtikzgu66LsNqQvE4RDmiiHnslTXf/f3herawpbERef6P/whhUHowD5
XjDtRdiw5B1/SJBLORLM/7i37hLKR7ofwqyrvqRQ68Z1u9dD3Y5iLCqeN7RK9D3q
60TTzKMc1x3OMvxPZn96yX33kQ1oHdvQdHZmb/SVAm6GYm7DOiSJLe2jAYUL9DQ5
jJCA0WXkOyjSLcj907AaebXwXe1T8TNigGoOTdmTVcdbx7FykbyKVebZ+zCVMxjI
Z0QcEgEaAi/0F1ahwMMl+gvvHiAiso/UW6yZ1bYo0DREPqh0vRlvkoJaWhcM43QY
XErCKBEzMalfY+nLZ4w7LV2sZe9ybfrCbKyoB0n+YhDj6SOHP3nwt9zC7Hjn507H
NPNiXQDupmyKL7wNuUpNwGl45bOI6f+m+bF2sfLnY9W6B7F/2m/Xw0tiJBmrLgkY
+ZPkSxyYzfRw6kQiLhvgPrm4o3UD6idoJFjo/uiK6QbosjFTtcb6PfVNS+49p3FC
2ITwud5Oz6VMYm9PXNKixXvjXtZsqbGpZESTmhtgxJRnpz6H3Yj1P0preMuwsnEW
agoaYwj1a2z7Bw37GD7rAifmdgWnDs1BC0/TqjdkgmnXA0SdAKdBlGyqld2Enl6i
6N2j4AFJ+4qgMScjCaOncVX8qEBJ3zXHcN9R2KU9h5YG8GzEBymt2KxRd4JKzlGW
+eebg13lrVgabG8qej3l8blvX6T0rp1RW94mGGV9bDlZ9cBg8ZvX5C1SUjlqP64k
fietjBqZAdUPgyrt+6PqY9OEcpo2azbQ1oglqMbKed+pj6HwtvfrrO8J6bYAQ2jY
X90v1/4auO/u++k049Q1ar8kYtCFdMDGNuaoVCPbFM/OjbuBhjZZdcUOElG+B0Zp
HddbSKw7Nfp3NujLKNNaUVF+sWNft0OSnQhF7yHESeURlM2cec/N2OAVaM7y/JZI
kvOeK3HuANNgdiH0hCSs42SgDHS/l9NrE8uiVBNzJ7G5jc2LUTbwJ80ngIg/JGD7
E4VmaphOAMjb19t1gFanZU8eNPkyrwhfIR55CjGxYoxndU5MdxCe8XHiQ4KuwHI4
kYNAEAxsHnum9pmzR29/a2iPftNl6tzopC7C1EVgZvwDfBGrSg6lhWe8IwKDj9IG
IDVfTPvEzRxSIc+cJZ0I+YQiGmMI9SkCsydIEwevTYWX3It/9SDbsHfTQ3n+ZKfg
2ADdFAZCUfQpAuRpy8ubxtHv7y+13lXYTWmDFBuL2gr/p1bYp2TQf0GKvk14gU0B
jEJtdT7Wb5U67+eO0r8AvVCTbFfSKT5hZnBlXcdvgZjdJswlq1soRYOmM5h0GkMN
8RvLt+YwrUxYCkO7Qz/q5GrXHZCcbrG+FWNcbOhneop5knNM8VbCFICfancwzvqb
0wKlQHKTJTcCYTiy34ffkdl9Z7/SMH0LBTluxkMoxcVMVP0IyaenQX27zO3Clb3P
/F9NIFYiN46syt0mv+55cmwUkmuTmaxrC1zMnpSd7l3ntxG7UunDO4NqdBOL710k
/63XsD2ljQLS6R5LUXwJQOsrjgwyTt/j9a5a2x1St8UAPBoKwigWb1fHfJHBryRd
DMr112kBmXFFBvyzNX+qMyQ7pMaVsyltEvs8chqihegvtq5DanbmBHtYPOfYA9/J
zHK2wiy37hd6QisP9jRgalonGg3zGi6fm3Z52B+HWlHj3q4Od3lGk0QbzxD59bFX
Z253d6hR3BXrbFEboZ34rBihyXHrx00ms39YqaOfrbLE1XChNblubEYS0+VLnkJw
ZAewnZKgjjikX+pfgFsmB1QGmlnAUIucwQxSYkkfyS44myKDGbU/y1p05dwIHPj4
FxCUtwnVV5VQpk6JqMGSvo2wN0zsMNZqolvVdf1+vZEbI/z9B1kcZTHef0/LywyG
1QsufMM2pPco6/vNekjCylr66R2Q09+X2BrQrOb8Yu88h2F+rZjYuhzLVYKkcAHf
ErWLHYfMZwX9ogGGxoVqR5xS54aVQbat3hDAbBdW2sMVnKSM5XzsJF5KebgrhrWR
7VjHYyQuc6u55IMSmMf92ESMajDRqN7tOA/YtgyfsP1p1fhFnT74HQf1ekJpkBUu
NZ4BNQ5/WzcOB0hVB836ta7nX5uPcqwnvoV6fMa9Y1gUnQ+4EIyyBXkOZ9SRfSHO
Xdra4H+v1ZoTD+BEoeoBD68n7H/U8nxc1KZwDBb9Nh0r9Np4r7uvBLyGKO5hJaz0
rauVgE/6rpOjWIGPMwqUs+iOdlDUZ3MoX/kdlO4ZXsiKfN7s2oCmqrKTDhq5H0MG
iXxLNiwUZGkgd8I59pEm9sJtQ1FhvhZIzJbWGotHkOzL59TrMFLD2Ev2izDLNqXq
pQG/omSJCRO+buxI/QDuNKMv2W8cfG8Q7IoK6TKGOX+z7BbnVDIWc5ypRwq093Ww
5Th3jEIAnf5YNajncCrO7M9IRu0fVS2UxwA+szujBXyQXTrDSeAfJLOSUUShN16F
BxxTmOAHQV6vmyld7HlSVAoK6wR2ht0kOUUrdWR9+r/fh1l9/t491CJdE/dcsVXR
E2LF/9qkoJffA0mlIjKFoNu/8LOl5qxIjD345yaLv8Ourtk64EWnkhi8iQOqNN+b
Fh/QAqOPguv0lpysqhC/BuSq3jJd18RTeHeroUQcSzbCg8b6zvZMmxyI/BGsf9yM
mFrzb6ohnvHyDZ/IcCfZmZjvCoEWtJ95Eq24eAAXB4ADqgE3UIVA1WDp8KmikbN6
+0ICwGJSuK+uDWX1vGidKJZo5h895G2G/mLFrYNEc8SFPIbdAqQqGZ7aByKVm0mZ
/hP1bIdesjcO6dtCpvreKeGtCD1cg7FpfOR/xE/AEC92lW/KJCm6ou3215c1wguQ
06MgJ65WfuLnOMZlevcWtmi/Jgr6SR4KBeocwMv50NrE6pb/7tL6mLmjqoDOGi1k
ODFZ7yIvoNXLg+N5NFnbnNFZVrrJnuEqA9CT6MwGRUyrY6GLTOd0+W+uz/kRqXjl
ZGWBt7rP+OtfODJwi6tfrX1zZVxKdhgwHD2iSi6OLzAR+nu5k8bEVCAVt9izjOFd
OPhF2wk9H6tWurVDGOojUbsxkj1KdGOC5xllXI2+xAm1DMjBq++fAMS+jGogr704
aLkOAdKksraMKyGnBW0FpGMc8818GwdDNxXiaxFZuh9qV5jkxElkm+6pxiuXmCsG
2kgqMjw3uM0uQhSPv9EjBazcm/Sdhz4/LJPUgrTnB5wjvOex6uwyn5Nyp1NHJE/9
S4WySTCPBClPqOY5RFDxn8eF3KlSHn5BBg7Y82ZFVwBU735pR+eOWs1fOQrrwien
ziZ9Lyy60Ztyhx8M8LhxumH0xXj6vRAIXVm5nQm6ODVlT6+ZSBk6eNGJhnM/kITJ
RGQw3eZEqdjqycm6pKn9YUfIu1U/BpTGNCmigBtjz0fr/84Xsiehjpo5sE+A4vLl
QqpaivrrnA4p2JqZ0MID5HeYAo1GaV2u4PD3jW+K84pZ8n9EneadFAJPZcwsIpio
Ix6e10BkUHpS8bARy5+DU3m8d9NQ+1L5Iety/EInQUDbLEElPOZQOtffD4VlkWW9
bU/NI3rF3KJwqX8NqTP0XtJE1Phjjx85g51l/fyWJKiRwWDmDHJcPr4iXOSqAkR4
bYCNLxBsmrO1Wzu4g/uKvykKZ+PjaUfynS3CePfd2MihYl7ahz8277grjJYGUprL
z/LS+joVKjQIP9jORB+6igpfmFRnNpIKEX53NB3y73si5WnchALlJ6oiV2rS6fak
Cji/Ja9Ii4gTT7zHBgoGTygi0vt4JbbHRO4qYIG+q5JJPOEKZyq5H3gihlvV+Z2g
w5IVlKrubFZ0lr2AYFRKoNEcSIizC4iuZ8XrusnLNKG+9mWiTj3eF0U56OnvnCo1
wAGC0cEW6i4d+DaGX3OYRTAvaVGAcS/BSg8mdJvCEtFcsFb5pj+DICP+5zL0wyjo
gaJNIi5/PNqpGmZQCOZGlH12yixgdh3Wa8BICP/OCrCw9JPi6X3fFTB7t4FVNmjE
/mAcn7fyNrD3oeRl5AGZKTo+4v/YtBVnTXBNa5Z3aNAU58FCKOeZm8H34tXWYSmd
i9uiO0VFTOuCfYQFuCG1EwdlZi46S5F4NO5BG1rd48JyS39LbU1TIwLUNfaysUlA
41c5ekbx2ybilMMeV8kphOd8ek35KVrJteenE2lbIPjo0A1d1ZeUpjuNZZDtm/b7
fP2+2NL7zmqRvnDuMX+3Ebj6Nw6yqYKOoHH5znLBt9bEaJwekZ8zoVNVftF3TGBC
JCK8yd6g+2lWLWe469aQzbd+NdS2TJzDIIdRnxbVeqF8hH29hFXbAvH2awJj7nat
kpDNy5L6NnSYnDB5MSduZ8BbNC670664eeHngjDMQZMwR+pgQJze37K9EFcqZj7X
IAKJ4lV83dz+NPNUHKCHn0HqhxrHRubXsFae3MaWFw6xbqTTor7O8Ybx9bFMQjnQ
Hx09RU+Wu1y0YZLD7qO98HDrbLAVcPQUmehGWOV2wLCE816T5I747Pt0W1cAU0gs
hE9qfPi6AWmBRxZ4FRtud08n5PuAFS24JkBGgEvwBc0WeqTRIRmcm8kcxJMng+lu
EJj8SES2Vl90W/7ac08mNQwpZ19j228fh/PMtHxQCylSnyv39MkDHEfxBt1+RqQa
0CFyhwDqFZHO91uJI/rsmc+abxF4jVfQLtQQXbJ6k8dU3PitoaSZDWJtp35UtGid
MDUc7EL4Ca3B7EOx8hEt8Y5UFZcUoAqF0jipBjhuZ77wUmnpFDEcCwhoUGaiI34h
eHWXp4tSCJkjiIFU5135c8/avgbYIGtBxu/U7hsJLhrV0MCDXPhDZUYY+ywTdSMQ
5EqZZyMkakHnOsVrayLGsCNsh31tLND3lbZpkEFmkPM+lgNk7bjfGJs53LabsP8Q
rTkYzt15RfVX2OZzgAHcUgI0c1zoq3pM6wcFOlLz3soG6rV1/YH2Rlze8uklivl6
85NbIpWB5b6hZZUAJnjHV6fR8IoK32ewLYLnhp/dx8TJmVfubDQj9kZg2nRPaN9B
6wqdmcpmOZc0ycFgKMvfXAvNkD2jOIaJPPtrN1cQhNls7E5wpE9GgR9iyJVCrHdS
0aMYqqNspsjExlLaYdeAUJLCW9Oxzs5yeMZ/ZzITd6v41i34St+epoP1+KnHQY61
b3jojC9zaPMj9JxGWZ02t4wgZrivDznYniGnwaS3GPbRVN0wgnKhsHiEI3pAd3q5
oHG6RHBMB9YbvXB1WiyWpcOlygs4JgzqEh0y+AtzqCXHerL01sZKzy0hu+6IAvkl
fFEARidGlQmo09xlPXOo4MYnDGrscgur/QuLHJtUIoDNCEFl1vstnSkfuVtZ8t1y
ll4qUz+KrXzgWeiabgMz1/iFqghpisd0HxNxuprasFPGcZtTeKUoEKXEDLw9z4Ih
r17GHeYBaSz10pgL/tu1hXcbIYka+7yRrUMeECBFDAKcozmt4lVxyAcsvw2TtJX9
30HJeG1jZYYmUon5lJ5U9lQmr+b0+4R/RIei8eLFdh9fUT4+SXetdpDwJIAzYU83
8BWenOH+OS9dK+87IeTFPdVmwgQqWupM05efGuBsj5p3w13J/j5PgPEtz+nq3+PE
2Z4MYCoVDR9kZJU1yFce8ZsLZoWcziZsa/ef0YXf5GOXgBdj/MN6+1La2ZKSirI8
v/CQeRBCoThOj9Yx/m4BX8zyrZUIuTYLD+xc8ObaGIBggNoZOhBjXbVTSe4C6z/0
QYKn4dx4fgE/+toGiUHnHTwcD7qpuwSPibVudHfB9CnBhfFcl9SYoVmIqzYQLkhR
2ryxFQ0dNyWAmqJXGkDDX5LqXCKwVBY28atfORZzT8UC5uQqx0AyhIPEDOf0IQDD
j8v/l4tsE1oZF1JCFTXMgiYsWxcraUZJTWBp+0yMZ6E8O782d3UCmm/npmctPNTo
9o9neINFQIn68Zghsv6uVy2rPpqNLv3qvk5RLrcJUYoTCh3imkHNzOVC31uMUat+
fDDnamKZBvXn3RLsfobsFl4esa8zedrjfkrHActSMSb0NLbnRz3adKdSfsFm/ej7
dZjmZUCuL08LDcDniEdG2XHmhi7GOlEQhOauI5ueMkvOdFYQdfWxmqizOdU/RmYN
77yjD9ZOlzrHwU5CTuiBqNNcMln/nQ8+TvFwznksBGSp6rahCf2BHvwR+gdCCYRK
ZQrGdCw6UZIa44DiTn5rJEc2lV4oACRhviqqpCxUPwc4h2vUc0S9PmwYaxNh0XMF
EWV99NMZCuNeLaiJzzx4VcUMpoPqBdZtPHAukzvHUPuhGLG9ctiYkJBFkTdUMpBU
yCyOxC1fxtIxoTnP+wg/i9ALih9dFIVEu0Dr7GUU6BBIT4LoOfqfmNHAJdFGV+l+
YtUWUrnNFdORG1moyc5gsF8EgbBDMap0STpgXIvEmj7+2jtUUum51gjT2UuS7xSI
XfVaAPVoUeuYb2Gaip53MA+Mnr+VYxE5uAL2GvTzWoUT3iKRc6y3BQoLcLCr/v8Y
p3mAAZKsLnMPu4ryLNSRpvlBpMcbrBRfXEkIlyiESebbDmdL0kTjzliW5v8Z/z9m
yaAWb3rYELiNGLflm1SbfeR6i4C6eUArYKeSQcEOlBMmpB3g+RZbDMGEHas0bh86
TjGzhbV3tDREsQvg8QaSFpNVV3kIIarq5uhqbdbDLhGVuy0r33pg6wc9VrIAmzok
SpVRCMV2dEmbmcU7CnIKBPeUly5S4LLesWWoEULpbU52eGRZaqs0AZv6vDP7bXr3
p8R0wWqCt+6g03SAGwM3GImwcImnLSMpd4MNxTEIaNxjUVs4T6jWyiSmlIq7kaBb
J47x3YHqHVxkrmcgQYVUnux9Dh9mXiM1l1eWzGP+S5AaHDaPQkI9TDqdZtOQYzHS
S4zKTLfdG1CW0DEEIC4EBg0eabym1IStv3ufOOAMJVxi1zHoBjksrnIXdqKJbXfJ
k+RtVIQDntghtzw9fRhjphIhD6vQVwH7ttQfK6aJHV72jcO7C9BLDJpS83qLYq5t
BQQtWhZoaCMRPkhqExXi+OFFl5PXNjRp2mrGXuuRzV3fHrFADJJsScjyELlXyyrQ
top/pi1c+e7oj8EK9RTM7PAA0zjAzvsGqyrV30Qb6x8USa6QKMD5CH4fJfnNJ1YB
vka5v7jyjI7Y97kJcFcAmn8Hr117n2RQ+RgFBghWrqfRKPf6/ECWlw/sI58AVm4S
eIitMFuK31swGiRmFytUggtpy+vG2209OXMtcqZ5e6IRezEZRKtEta8GTc/MlpkD
J7e4hIpI8ckbWk9gDCi8HUa+jVFuenwVFP1Jj9HD5RBC+77wR2v3lhBZ2GEVkTiM
fzQvs7VdsUxKre0zZO+2DApt0N7D5Z+5XrRXg+TmIYrNjwVtxOai+n4c+2njgWp6
WZ9dEs84+XuSXWzablKH4aOak6yBB7ethJxL8SSANp62e592iGYU6WgfXik7zAq2
IipktsXCqLAVK4JOS0TkjRmu97YvnuuTjeMWGlgnfEHmTzLSnonw/pB93wdsDIkI
GmpErCMwgA9TRpO813trpvPD0StzzAzqwUVM1EP/qGSDpumvNJNJadGJDR6mmWw4
mQUzUTwDc5aTGuNwU1b3TYRZvQV0U14+E3urGW/R3H9B4EI9Ma/a5n/V7IlFNBhG
yMudVzmeU2/iWzCubiT7T3IPpA+4BKSpFJiMP5lbhGjYf8S36lPVoOIoUmfvFDHV
aChQj89ku+qM4ia6Rh+spVY3+D+U/KW5x8KnKY+CGUWH8enSOtxfHoQCHJSvJs4H
FlJ0PoY/l/rZ41o9Uh9JvPr2rep+jWOYwNMSlASRcygPk3zeV+Jv8G2L04vyz16J
uBcsZYYLfSu9gHiapqFCG1SGEvXpUAzkbCPSCq1g4ylfdA3I7zhfvpIZR4xevhc3
K/G3FpSz+J5ttlUeomjfVJ3Tm8OruvbOhmazko5CkYylh8aXvCjl+AK71UMJDeu6
U98VJ/QNWhMGKP9gMiR+PU8IgV4dQXQYML9pVbT5foKGPL/F8KrXdmuCLn4rtcr3
pvmVv0JKKlkUOeO6tbu///zQ5JYClUVIg0szjTkM6ivldaGe8gqwgF5jKzro8fhu
pNKlNGHPnCTMjjNw4lGU6tNjZ7Hf62uJGX/VQNylCNlr6oGqDETvaC4STttmcPW9
YRJsTqwxRKDFEIHBaC+la7NYnhqFxCsVxiJqWiduW5TDyBOzNsM0o7Fm+Km/Wqte
y7Z3HkCcn/OfVCeHolCaMvwALTwxKoxMYjZPvoOauq9fUeFHo9RLtOzz/iWBiF4V
pdQnb+qZud2CB/KDgwb+mtIAXOyqNvyY+wRgWT29aO16E7jZyUy8U2u5QCGFcql+
iDwQxfAJ9lLYz8j8Yp2ZcSQBAgzbmdq92sDi7ge3jhFlg4QEQ0yVUsYnTwL1fsVS
6glJv6FfiBBTGvFmwD9wvlJez+yuMipUmm4GJ1v43xDyUFyWvKSRbG2jQqgyjyeh
5S+FbPCUCEEOnSdvrhaZmQGY+/Tpgb9CLFcZ9sURuyDLy8GLATqnuDv960fj1Q6V
fWYWnT0BTRkpsCTirpYQyYXkoy2Ryy7nsVSyf9nxqtulN253atXAHYtcTDSddksG
Ejk6f1JzNphrNOM5AMpeJNqvhQMhQ2HQZaeTYTTxKtHh9NEHE9mRfOjFokLgJrhr
8MppMumlHvrw6e7xF1gYvTWdnlczdBY9RuEmPJVPHtVd5k13nhtEQfL8QVCv5UOC
ATektjaGWgKprfnr6IsjJ4EwEnwbEvq3w4Vv84NNNIfuXuV75vRSEh71vq3n45bF
SwP4SQyi0AJjkuU4vsouM5WgsFHLuUBhso5dNpQ/9HyKztilBHEkaerBwGcshz+c
zhPxT7Sk1GLwmmrNoqvv/e2hRW0u5WnZYn2luTDVkYSQc/iJmwadmiyLPVxSpGS3
o76Vo2y2zrF9D/utqireWl4EQE/vTkOSyyMZSvVk9wbirJBlR8gYqrf3p3S18uRF
r6rV3vvB7lqj1QdgXy6L/fS93VsEQ9FKbNVIbgEKOWik+NSUvgVaTPbjVG0CzDRh
NYHcqHIIOgEjpe5kTqD2hLevOXImTHknrTtyyLoVQyQRKGLLtSBGU3oOQvSB4LTB
7UpLaqi5xIy2So5KfmCHMc0yAc7v+AdNObGI5E0PqbMnibOWgjc5vMgAoj7gUWlZ
bYbZ/Nz1+UIQ91LY8GwNX5BxGXkMVVF7OMsZaoylQStYMt9oBy9U+oOLieKdX2cj
ZkHZmmPfgfVY8DjRi4Wd5D5+lRZS6lEiHw0OcjUYXz6Yi3Xx3jwZPCPirlSCmPXR
YD4/7nGvxKCu78NB9kpvpnXVreB+4E7p07kpI0v1lEWFyDVirQRiyH+bIfJKDeW/
DnLBDyHQWGpy6tK07IPnA9ECTBlQPcfyrCTK6Y0kBMpBTMC/TtlwQF/P8KypTPn9
nVfVvf8YVoXIumVWEx3CtAMwvLqI5BlUiYzMmTfJW76ZlZp0w0hzRkDA68cNLVyM
wgGI6Cq1ZKtxxNFZu+AFrj/sPyNTBnWEh/gDLAyi8cLa/LC9CV3gqnHMl2WHyxQR
loyLdUxXJGmxttIxWNdKfPcx/Twu//wyA5Pm2cHhjyLKfoAD6wA3BTHX6EelUR0e
+9YuWhDxBHF1fWLrkjuDUieVH18Ap4S8nCVF3UwWjFBekNnx7xuQ8+NeSEpJafj1
3KFoqiPqiewBwd/jkRhm8jx8/iBKM9xj4FpbI8GEpJxL4jSQOUI6FXAwsE0bGiPB
6M8H7f7uN3vNfi6+s+hmhZ6dvEuK3kyGld8ahGXFzobFNLrPWaMRP+K2pyGp7TWb
KgHVzbE3BY1zxDL4paA93eZ621gR9ADlaz6UbBbx9ip+bqGofzut5ftMS9KGwJY5
qfnwpUpqs5e0dg+oqdD+gXq8+U6zQgMOD8sy/yj4dH+52j+keYTZyY31bDrGIIZ4
4B02f7g8VtAPXk6vqawl/3z808mbji6uxvRdQSGWGTI4Zncj9mKrPh3cbWkF7wZ+
xKyV/vL+njjb/d9t3KBjfI6q/o4CGHetgSSeppdYxakPbj5gBl4FEYP/vD1Q9Vsk
gnaoJBe/tRw29HSyl+ABSQqKmGsmJa5CgkqiGJBh66hMTGV61gtO/1f+kUx8dgpU
bgiHSkGBX3n5b1V/RmZtpZKEc2/hWyThUuLmhZp9MS9wvS0GNMCeTWH3DddDyobc
enyxF8K0jl/882Ve29UOByB5CSqcpdkllyTnoANDJmXqAfHYyw0FD7WvTknXb3er
RJkZ+U3zdgQIqa31zPDoov53fTzxS6mdAxG74lnDKPDW7eLQq2lHk6nBZ5qJ8/85
4wa4zIqEvs1C9OFMc63AbgqHc9WVgden8d8jtyJC8K9jkR85NJvCoy/KkzLVI0y3
ZipOQrsPCGTMdx5m/rr3cZu8IrFj4DKzFqW9aBpX0dDaVwRKd6bZ2TTDphvxUyPY
n/ilEL3EkZeIwzgTakRH5B81DZPR99Mb6CNB5hFVY7s7v4rYWcsGKHXIqPNB7AB9
XxsmRtuzA93R007FA2+UIxNg/lk4AJeUdyizhxvKMqZSqQYW9z4YUyBA7xc469Tn
c4i6ujsEkStZ/fGSCvYUeBIf1DA3Pe2s/8xA3vb2zaVZvXj4CRmt/GIvlxuRny4S
GAi9StPXVB/USawOAEzeFMWbBiXjM5svNvQ468jEOd7ktpYc91IJgKzONkovlN9u
wpxpU2555XlGolLAOqyUGDInvdYHwDox1p8mghooWt7yd+wEAyv97BjB6LdLuZ0n
2gikA/U+GsgbX4rAsvpqZo5wyllx7AZeuFYaEvhz7bZ2czyZ/J5J50IPtYrHqF9X
ch2v0bA7BBElG9/J5vuAdDyxKzGUlFYxIpdxNod9EUoLtFL4898tGEIAMONRYwkx
iGKDIG7yeKFOTjXhJwQrHc0f+Gt37/D4f4SkKvLPip6iFJCn7+94IvxyvBplAUSZ
qj1K++vcT0pzv8GiHPkepj3SorHIbfJwPR8M7CmVay8Y+2dHxKTuT0CDjy5fcuDW
yAT8BTxmCd4AJKc2lxskgMDprqmSKdj6HHGTTPlIoW8O1Hw72X8rRhGH4SiGrHRa
S2reh5hrRRlWXtEPy2ffTTnKR0m3BVzbBpDjz+GuHgZr3ChbO2d8g6V0BYr6VV7v
pEkXxCjhe26q3X2vvzfpOVv8AYWStVN9CWwQ8xgXW8ZjGhe2pb4W7K7ijoNRlrjg
WJpkvpYpl47oyClUFGiaMjfBFKw/FWBb9EqOxcc+I10bs/IQ5oNJvKDyBQmcKZO3
5MdwTX51GfsY+VLOnCTVDXM0S9RZRuxv47U778a1N1buvpq/zxbT60miOASB1wNs
z4qPcdP0fa74SR4jUwsK9Tn521cF4sE18fmsHAQ5Hl2+hVKyzzLaPgQmAt+b4sy7
vl0ut4+b3ToIJaHudiqpa2qmqN9AlvRDzDgR5X3fGjmN8ZEpClVBJvubP2fbnOdA
L9t2l7jCs2abtvwIQVayRJ8qom7s+cnZMKHNAKP/go1kfikmdlGouT0RGhALx8R7
g971rZCBlIfOYWk0JKwNvSQIxc1X3GJfmNBR7G4kvAM0cDAWi9j2qJTgjAC3a0Hm
gT8WskzUUvwjqjFzEd9cw7Q/UAmc438A0Ja38aPu1Bhl8tgx+jRnUk0FaCXU+RKw
asA2B0HZidNWQCuVQrfA8cc02VZWbDVB378yMLAqMfg8f58suAdB0jdsuvIaE5eW
gcb8Y7pYRulcUkIEI4hlHLf/HefnOmcWaSYNTUxf5NlEVoEhGqH0I79+ims+Dz2P
TGTS1p2Fm7WKyIg+hhqYfXNLjNnJ8tX4w1lxLdpSRC9tIUxXSjuBxX6+FkX96dKk
1LHLje7ge8v3gjC5qM4jzhk0qXxgb6LDQUeT2AwANCf+xRJ9SA3qhzezjIezSwNd
TbQCNZd9Q+S9kJ2Joq+15O2MisEmTOMOSb2vs4nNPCF/b9Vsm8S79fAsGmHC/aEL
YXLe8hXGgZxR4VHpm/4mRdI43ftf3IhApblAOv5G8xw2J4kUiAZg6eMGzyixcGif
GdJkWN3rMiEp7/WYnpXAVNq5yElDxMw3rqz2Oj2loS4Eus8kc81jmIvC8h72AMvq
L3E+RfvhuIdyVbYmmaAyTcIfUvHspHAZy7hDEGBmB8KPaFAyKxnlgdd/3o1fp5Ls
PEhLMHZ9BrZmXVgyQtqizzTXgCfYvI4twExAr4bFVdG6fuFtlxNs+WXeIqzD88FU
oL495GpmD2sn2aGjtH5JZrITfyJcnS9F2wbTzV6Nyta57HE6g/ofLRhEvsNpG/uZ
qIWnzAfBI5uHFIdk7+Y4SnPL1SwvPO536iB8pI1SmRJouYO9XMNnCt5niNAvvqrP
36pmDT7dejWDdXJ8zgxA4B6hSbUbxHHiHPWdCdSTI0Sah8b20a+PwqJTngReby4A
73UMdgBhLMrGG2OHj1ClTyB4q8QGh3tAWjCGv1GIe043hBqMRavmxPYQOSsxg5AY
V+VqM4orrYACjjPmnH5IaB2k718j0QFZpkDbJ2z0fWnF57vroza+zGVIRrp2foPQ
BxbYOgTnu9tJji7s82oHgV4fn7Pous+t41TnQAFZVo6OzP9JgsUYE3CuzcbLlqhW
qJvMCrDPy7AWWi6qth0qU+C19BQ6MJJoDdOO9O+f7XBRxfb82JdJ+esGhjYWzM99
wQ8n7tSfqBG9DkoobHUihiBxdJ+pt1vuJ5WKsByq879BmNJ70iLMJVkCObleeW5L
MYOb3SP5pDMErAPyLzJGuQprs0Xkd2/Yo+U4jvCFVx8ACouozO5UtatHTCQ07J7+
7ESWY5c+QadC+PwKybS9dxm7SoAgg9UM91uTVzirqT1smKIiWd9ux0BFUHlX+ePo
RhQ7W4Zb3JT6zwB1W+rQsLAevBOc3QflDIqp79BC8I+ErPSxLhOexAIfZeuz0RcN
wknovxPicoOJFXdHsL+Gxq1Xdsn1ixKGPt5YRe/FykGKLOhbzAh8liD8Fq4t/qtK
+0xm9z+qoID10xK73oEI8MGrRMpoTdiQPKi1Ko5xKfN5csFZqd3wO0XoUK7NGAEG
TpppusKt6I2SHF6K0zq8COl4CFnQO48lFR4dYnmYEyduexvHTE4TFuOtMily+uLs
MZEoIS3kIZ4a0c1RxkyE8JsX42Tcy5q54qPTNO8M9GXKxtK2PPITCZIGt93rV29F
xiw1K4u/YLv5uF3o9YSiPk+7lLFIzq3T+BttDo4UCJ/T8rRgIGUa2h3PCKc4bqoq
Cu8F7L6htuuCJWUwWSYUGf41dFByQqHWPJn2tsNL2HNYQVjJNG41Z6MLcQhQU6Hr
ka98OvrdeoZtuCxje/sXKmcnBiy4Kh/84RBMU8ct2oPXYKAP0BvKmZuEDNAiZmrZ
2ASKrI1cSap2WbifxWj4+kcXbzeoEsq6OyDDXQKIJr1Zys7P3tyr+W0ov6ZICq0N
w+noMJNWTUnnGEcC/3Wp6zMRIFshOx/EkXswjarq9iIYTvq1Gmln4cb7RovCNTgQ
1MCbWyT3vyjBlbM9YkFYDNESedBh8gSWoIgjH7HZvNTXIsNGEaxE1TCnU5pREXtF
rhUA1459Vhek9zTmaIkPa1TRsvmDIpngSFNL7ngU5aTEax8Ahxby+6O+dBwYVekL
BUF6HIDqfNi6waccWdqNX8f5rJ1l/xpnGzktQw8DdA8GzKdJ2SglUfZgcP8/sN7X
WzWwpdpTYo47XDqlZgENnwmj/ks6zyp/G4YAuMcHJpaRvOE355puFnKLG7sGt7w6
/gyBbXNCZj/pjIbtoalhefv9uJj0HCuJsgCX8OOMVFK2ls+GtR6FUvATkQkq235+
CFiJn8s/HmOxubd+uMMrMePSR7NW2f48Ih8TXYU6ZfpCks0qObQX5vQZXetty9ny
PJk4T5zbrDhZlG8JJzwp8E8q/c1zlqYEfXYApKXvIPKJwUKGO4cM2FwXtDgp0Utj
5h0l5ky/TjMad/uiLN9pM6ravX+I/OaouS0foAJvM0EITeOfWgo181ZrS2lHD0EU
b4vJLO4o0Llmve/eCzRfi6HVQfhrCGUyoDVhE73Vm+b3E3Jq6Fa4ak4PUeWqDT18
hFwsrg2Jfv1xyDs0h9SiMkjUq87GbBe6PPxzGxuYB8CdgrMCuxhf25b2335k+Fwe
hSfTldO3QT7+26tRiaCsDBqxfUXtgzoDx/+sW/xmCcvnr4RbDu4pXi+IiREY5jIh
BmIIa6CvEVHwvb0SWhDs8F4F1A01wiJ6CMfuId9qmF57D4i8epgG00fe+XG/5Lok
bv3GIDo0CgY4a2oybn7FPdh1qhql1nfCumujEIFo3kCRfZfxAD6qy1CUR8+Xl8VF
SkkyzrqymGLijRTx3hy3JoRATXkFeY9XtHlGlood94dY5ntMJHH4xHAinq2MVMMp
IbUyka57nR8kr/Ak/fMbbtWZm24I3oA2Zz9LsVhnwuMGtHkfMkr/mMc9QYLIR+L7
AFj1t1KOrGGrUTNCRkOh5xHwpT+VnBb3HqFgCWo0nTmrEYnwMHZhbcXcsPi4nXeg
X7zgaXx9VVQMeIN4KkRLzuTcBhOEi7mMygKo6ii4j3+0sZzZMOngsJaYX092SSx1
Es++hyGCTwjwdJNKnAqXhuyulAliWH59IKM9sfhkFrws2rKaDj1JmMujb9yXIJqy
iJ7ydRDeCvA++SMSPrQaayCYUZcPgv74Es21C6qsO9LTTnfAc8GZxXpssgj6angG
J3rk5JpnqqUXPqE82rNHTVJpnX+BgSC/d5Wsuozp2/JTGhwAzsB+ZBcSsGBB7QnJ
oxKV3+wS5ZJJblgYiSXYOKfOSkV6hlygf1lnTP9fqDRr8D4tsJMlcL5WdvEthl+6
m7uDFwZhBeOGNgMBtPvQO3aA/RJgsPeeVmk3mUjspoTFIpuk+SOnA01Bx0IAs6SD
Cvt0fFebNSlT7+Cpu5O4TwNzH9VnWwbm7kBMR8WlpDYlvYTvALvTbN71ym5+chln
EzknO6W34Czdcj7ddNB5CMWVmm2PN+OvDIylkDKmVWIg9EMb87dcEAbhS7teetDF
6KAa18PThdkWxoOnJqq/5M8E0sqPtU1Hoyn2SYRnk9ypF4lyZuYUEoI1tLqPpmLR
HVqe1s2GO8NE5HxH/eTYc7Zl5miq3kOUWD+FPv5rQVeT4N6uflx0jiOH4mmJD8Iq
F1o8V2a5/87NFb4RdqAkWkViVReqK6yedIPkhiYwxAvz2EjKE18NQ3wxCF6bfqBk
J0VBR/HKHY6C4XjcMZ6R2DRPSDAtFgZsNiN/5kMIssBSpVdQsMkhYm/ObaMG3B7K
u/rG3L9Y9ytMbN6K8Geb0GFwJXZcb/UgM7R4Pj8jZQ8lkG1SU9dfMzJrL//ALu17
GUM5rei01zoOwWLdTEd/OiOIS0yo09CzmkoQvMNTKOKpxLLS7vJs+vjY+TUOqb1O
tSLuUVknwObamFP3XCnyLL9yZc905a/FvP5vDAKeGqD/4pH7HI0axRPB5yO28soE
bIJ6xgxnjdiZ4qtW2OLtWeVHcyWpUcsUM4JS6BhWcpJfvKQzEgC3Fa43yViIWmgs
YSLz1BWrYBh4GC7t4CfQ65lnKN+29L8hhTlRw0VN1UOLI4QCnQjsrXeObdObyGrG
c8AYI4CAfBOKAS0j2eAuW35yjoeJ8v/mBM6U4HCn/cV8Ug2NYtfLWUbQBrJ5qW5h
tFyIOIPDyaHpucT+BSoiMgE7a7EhL/H3jzhau3Z8yYbvBxXfwj8DjBLwKV/W0crH
rGOfGv5hqVAtdebrxIkcyuy6YSWA5ceynRvgEvzj6be6mH0ZremDQaFxn4Vpq8eh
qADqbWpx9QOnCdubM2eFh4NyTHbljEEPlQXU+ejl0Lnb3Bi2D2fInNksM5aG2noQ
H0KL4Lsdz1piXsLxaY6ONCr42UJocxD8ZAB/+no7Y/WNfs8csG6eKs1QXkcGZJSV
6YBbDH2Wosy1rYLn/G1hciTe6F46jbg84KpsRHwfD2bdMJouASbTEYHAfAyC9QQX
lV+TGKLxjjhsSnDqPwatxuo1tUWwS5Hm1+IZyP/X71fA5bKT1SVGDfX/Xxd5X2jp
KxpsAlSONrOy/jTOWS9vHxE6hkZvO7SBcMYDb+bKj88uvNxiLl0UZnDNcA65spIS
a8RS7gLPqIqy9mlh/CgJX88fchj3N0m4BkAB51LKVBJ3g2QHHo/jQvaICUH9XGO0
cLXx4OlkOLflwKCcXAvI98lr54ysJYqgT8Z+YLDjwjtg69PQ6M26P3GtgqA9PH+p
8TXYirrwzt0Bx1kdZGeULZLvHyvqmzgPWfnWfXhhOoVjtk5BlKxBNMtbqpGRnqvB
d+yLkuBYfbFcMRnuz1QVyIZefnonY4TWjo38frfJeEAXciK1TrigNcd+9UtexOw3
BvmGhICBe7b/URRButj5AuTW4RXovo6GSa/z2RGhUytZi76F15Y0vSU8sPsYFd+N
+EFJASPZga0UkFyvtQJ9sFhOozaVQF2U5c9qmrdFJ2DVlJlvTvBiDCmavJZZAESK
NU1cb3a/QSJ5wmgy/7BsrAFzCP6MPY2i5l9m/9Bf/KiQRs8CoSwK6T+DnMGcjNoW
ZKArnqsrBPn6mPOHGqFDFTChgkaPoQ/wHjp//lxSVnBUMmcFAGI3i/OSmE7S4hg1
7tNoijXoVuNpEVhOlSVJ/DhrbfF85eL3L5bZSnqDAhAucOplGL+19PBW401eAvND
NcTRAItG6aG09Y+b/VF3i7ESWTYySP24X9+0QcGwljyB1X1/VtCweZgEgHQiuHoX
5XkEmOWKbKjS5i6pqElIap8AZjvz9bT0jQSmKcxSehExoLL1GVgQhn+lFHkPhlX9
ukhJHaiI02b/ivczY9JVgg9D2vBGLsD26B+p5XoeDSrquqsZGflm4MFM8MVOaGzJ
q2UhSrbt0KBctBOlcok972MLjOmx1Jb4prikVg1M5hAoEzvF+eAzAyooMTvGEbGZ
Ov3QTNRUcTGpzdtOdar9PFYvc+T0bvkxnOQhWNTUdRyR60nuU7qxr3Y5LiRLtso6
utv9HNsK6OQvLmce3jpa8lYSI53HiovkQ5YbaY0xudK1lBVwDy8utYFi/nnKqEhN
1/UFzlLMBNE4CJjwOwsSueb5ceaIQDtTudjSMvN8aLFpiSKKfNLSQBCm9L4uhjmo
tYkYkd2vJtKFyqKsOtjzTYqlru7c2ntXxRFVnpdmcWoFzRzNXMMXElgWq7BfaT8t
ax8T97Cg6T45hP5Ir+WLQ0+yfQhNJlomVw14A27QmaaPH2gmyLMNRRBIbvc94o2m
jfrie8FJDhXcX8TXBVf2QpVROF24q+aEhlgiEIyjUsvGswL2VWNV1OAV/FDkgajk
xSdHd1Vj5t5yVZYG9Yp7myTNKkVCiYg7JGtI3reYhHDdXByl9ptAjH+rfrCOVZSX
2bFsD7Gnzf6OeYjFEkv+xf7n6yJDqCIpZfm9VvgZktrSmXWTdFIGlK8CPsy8YuYB
hwKnuWENe5IF33lVawIv0a5tLBObZlvYSmeuXd74dsICIKTxoQazvxQEmzdu+Td1
QQUGj/AUYfHciJAOaotyf1WgGMKNVGNyaWrVMbnQbFB5q66a+lz4lTGbFyRBy4NC
HzbXjV21I+TQfxq4q4uq3AA5ujjHk36IO+xQa2/YJhu8nk3ZAZyxFh4GO0CCXOft
mTHmdlyoUHd4PnRT3hMnz7EOeUPN4ibWqvx1YNw66ICyEpPpLb6cY04NVcyiiwRm
lKjPrnH3bTU+dXfpXfqFfh2CHEoc3i/KFxZR9YIdrs0rmsNdhnRTY19c95EEaO4a
l6OHs2zO9NrK9FkM77Fp7N/WTitURirq9Sd/QBSO5QuDCYemyoK1dCW4eQM5rug0
GeFvoi/s6zNMDN+DBaz/hbch6/mj2RC1ZmNPogjKCI0kkIuHaY+OcfSgLGDPXtt1
TPpZv/J8TZbsETWdIgj3MUv788RPRkg5XU5KJ1IxhC3ib6rmUpxo4eAm1nRLJOBV
OjA8fMMMcj/dw7hSNEthlunLH5rXYXsAde20XWis9iTkl3erAx2Q0453PBmmRs2z
TjaYcGk82uG4KS0RVkfoVjozQ2iZliJoREaucoLpTyhircgECEUpUO7w5YMEVrV+
F8jupPWD5IGjwavOrD3npi1Fmb7qqPEixSix7QMUVg3O5iDArShaI58P6RQ5Hdkd
SPG8GgEsXte0gzfU3YfW7XM5hbK9QJMyQkSpIgyExfD6D58EpgdShR4I9x0fUCzH
tUvlLkyKee14bnvDfYyLEcf97WNTOkYFj7INqyuAoEahPVD0BK5jz+jBf54Od+8k
jYXUyUx2//xKYPWWa7SP+gSm1AvEKBnJFsacD3L/9Tn7ROluFJGE5OfQVLIsgclZ
N/wTxEuUtCnaJFrO3Yq2XsxtJltF7wKSQezW4pNZGCAw1yG1aIOlmrKZxKF7r3Qh
1KrFq7s4swCMKcSkDnuuU4YD+twuFwBCyrLTYg9741TvbAcftGSbv01Njya1hQMF
3byDT8Z+wKmtn0robam6oPHkib3N/C5DgC+De8+F+9lTmcwHTpwd2tt5tu7CkqcA
CzRaiR+JziBmk6xnnZ8/YqIprtDONvEnKE7hGSuklW72y+tpklUT0oIISqtmaxOL
urpFkSFDDLk07GUOVPiisgFJFc2mmpw6ktAsIb/5BHrbyOw8qyWf5hTI0B/bym08
d86YR0AgXqvXthpINPXXleaoOhcOPimRcU+eqTSPxacEweEYfgTnSedy9mrj2Zhi
4m5Yv73ljWUbGQ4UCLGg+R1P4x3Xsxi5gr1h1OYpuRPopWaiR6juZ3eVf9nX2sNl
LApo0vmfk0rZRwujiESJvNmIu20M5pakqWqJkXogoOLfOJAO53JYOrpqjzEhjRYX
6p6/QW+tQCr6gNDRIs/Hphh8o191wFG5/qOQNtVFLEDmsGcJMHjs3ikWo64S2RJ9
ibLA/GTc7NdgT+J007U3+irVXwJjf2NNmD5B72NvfN3CwiskUyNuZttfnP3zBeLN
fSbpPj7CNnIASKryyXtGN53tWjobqKzUEc3KGlaVXRXjCDR0UGLC2j+qVY4kJovX
a/Gvh69l9hj/njjShUt1oADF9UBPywzGg89z8HDlTmPl6sc1Y4LGa0sPIJUJZfbk
0WLR1D4gXYa1VJ62Yqoz8q0JdhsvSJDsEoyE/vDb3TZfypfdEh7dluQquS0mZq1X
5Tkdfp660+xXJqrMm5LCl8BHdepV3ndHMbQQqYPntzvMkY6fpocF6K7qFwczIKaP
lwZ2Hy3F+OhFjPxYcBN26sdrL0w1bVDfpKts7K0TFgsyMPYBRAdfSM1kyzRvF+SB
Quz8dOPqLIHTQY1Xi6KJXRS54ex2uiLR1R1yBzzIxFJqoB4Qm9pe/UUQ8RX0+cV/
6+aPjR6MkC0nHr0w2thp4xWbt1kqoVxeQ7kNesK7/3yOoSuYzoiEOwletEjbGQvO
Mz8YLBnhdjGfUHSWrf1I+xxGXLDPkBUxSpzoP75VpIAdvuEqPEEiTaPL7BTwpt/x
HJ74y8jXKDtck29JAsW9L+cV2ESBGVI8TmcgQbj70d8Jj8YlLJzYrNf0wTGgiQ2Q
RNu9mvAlNH4oHsxNOG5MU2WM2sUtmEoGjbsa1ZHT1yWHBAMYZaPC/vIiaIQt7Opy
lCsoIkLtkiAQtakYjkax/7VW3SsGQihdY/8Di0W9EY6NKReeBQ2KZaasToJqPWb3
6KC5TlPp+bXXjweHLF90NpTlLWxcn8qmwzIuM2QhCDS1s+NEbnjRG4FkXKpBNzfZ
ZBR6i9aMJ4+RAzBg7FH3f2f5B4RgNNcinstxc0SURijKfPeaMYgaepK8fB52Ny95
AnPQIVv7kkklK4+A08jPFNaW4haPcw3x+4vnU1wfULFBzYIrbhXx0KzQ21Sn3Cq8
LQ4gkrt7SGvHZeIpW96a1Kk81cFkvOBvHVoqduGQTRZylkhVtLfNWhaBck2594/q
SjXCIH9TqZPDoilppxI+f/PQzxT5BMTYVHsTknTZCYX/+dzoCzKs6h9uwoB2Xhmf
bw/EXI04Hd7rknf9UabhtEngPwhWhU0GdMpb0yT+SUX7GohYpAqgxvpRzThU94Dq
n3m9NE8Nbekxc8UhzaV1Z4ssb/kN2TWegWODnuomk1k=
`protect END_PROTECTED
