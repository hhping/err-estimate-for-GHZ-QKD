`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NNY9Ds3PFB++zK4i1DNPb299rX5s+llzDZQ0O3Qh8mywLNh6uM4MXEHEKlZX0XTJ
/0Q5g5oJWeIohn88JEwCvLKQxebGk1HjevF9v6Cdd8xj8kNqF0MxC4Rv1x4JyPJA
2asm9t6zFttdPc1QX36O9zNBrDfvYvv7k5eBnKmwTGzLYUiKY09nWv5gn7MZ8BbS
MF/hgBKy5jhOKXD3pw8hOupQSbnRX5uT4OnnuJeJ21xQQ9n+AF5y2fArr/GRvs/b
VUa2tYj/+WTnujyRfoin/kTibfk9gVL/MjjNDOWSTvBslelNC1/tRgBgdiBNJ0Hu
OaMn9b+YWQDrP4D83HzOBOgkIwn0wVxetfmB5DD5qHfyola1GZvSlHcvRb5lCnda
mkaKK+yQzgG0wd+XzgvLZpgeSXmoICVePQUfYnRm6wsSR/1r0xCA3GnIDwx5zBWf
tiolPgxf7uWx2j80/TUP6sZZKH1vKxP9GQsw6GBvHTnfb94qbAkcoiVTp9M2qLuV
xW5dovTvZEdv5lctXaFWRvWqRNm2EJVHtcn3fnSqM9V1edS4fm6+yFiL/UuXuk+x
fK6mHwbjmXtlag/fkO4Z+lGiSWjm1RobfPdRSaNaEpCVaE/YJnUdYTQtK7ZxJ/ap
kTG04VxoGbYzX4WWFnHe1jVVgdrmjRvfpSXMYmhVACnFvxSFtlyKvcm5DZKG3WsY
9POlmG8mrTJCEOrKhLI8jO2aKVaDahdpTek5O0Fo297ufkLiYOyHRCCbrqqjwXE6
OK1E1mGAGhwdiyI8vxah6g4/NXeDvMxuvqFXzIcRQdkqb5yt/pOWZo4URkuNc3/5
VhS+o54KZBEjuJD7dCVyKbE1Ux19gJJ9Ha84pTfRB32/+ueT5e8wWht87YuF+Ib9
10wtsKaJnyh+Uu1DnngYW1M7aqITuMOoA1eJtuv6xg/Ssd1A9N3r7MiZLfPDj3tc
se32o7oe97h5IHNjMzU5Nkwuu2GK46/dN7QhDGXs55dxjvJ4ge+N94iN/ro6V/bf
Td3O0OagECCdWmKOriMlPYSqw9sa6jW0gQLDBqcle5GQxhoTtcI3WNqWm57SOTtS
Cp4tXkvcu1d/mUuMd010Oy3SiCvQr4kxq1ODjl2piB2c1Pe1my8/6i0C9ViH1dfy
6Ajd6xxOTUwWiXUOwT/ZXx6QxYWc9JMlfxBg/yH8AxP9NuUuFTvJH9IGMpHMJyV9
aWETTH+SCVZ6ONi3r/sJHp5EMzQ5158u5gL2NgV0pszb24iboCTDc7RtJwwu0dpk
PRG7lWKZBcjpVKbFb4RzD/Xw3bUtJfdcaAxtgCeO4UcWOfquUEwn265hSXgvekRb
hHmmeOstMZ+DMwBghj0O3yvBJ7NT3YlGDXul3gbiXMxY98Czqoh47fO612MdOU+r
aMXMakzVUP4ymDvshJwRxGz6LFo7q41U5lrGp7wiZWEbEUp3sHsymi0JUYRnu/zk
YIWqUnA2i7eu4IkiEl5U/mvGbxzOafMM4Gr7Ns+SZr2ceXCFRJUx4BBer2XBUIz3
IhslD2XEL0NcXEpPwRewM7kH12+U2t6Y5BA9Z1ehovhxZbwtYqgIwWDl0fdSTaY5
8UgYTD+KPDBHfQHbZhB14cB7/qzRDwCIcFXiD1p8+qFdZQO8wcIqaYXzegE9oGyI
//kegHsvyahmsXbdhDDzfES03EHsxIqGgMZr9qykfqbOaVyBlUs/ZCojFrwOoX+u
cCdGNIdizl7Zsn6jDojvmSnbkke6BYpOVE+Yc7yjdVAvNfAidlCTycA+oh0aREtT
o5+//7OubSBzpqtalfX3I0MHv/dOZ8dfWhw4Cph87HrLdJfAZ8/aT6nIEt62PO9S
h8MNgiBkNCGqjJVzRo7Kg+RpRzF6oHFWtgW/ejS5Xv5q/vTNM3LP216eQHP8MIlj
n5TM/ZtRJScdjAzU6IL7g8DupddulCPCQLuYZaIdSGCuo85yu3KJh3AxyYdPy5vm
truaR4guBvHcEutS3HzYndDtvZETDen4dyc8kzTDr9TqtITwqaqtPqE0OTCg+yXz
sMlWTKdYxoZBsK5DaHVIqrGr1Hz2P/oaMV3ESR+ilt98ZKywWzbewz8pCW9QRHL1
LjWzltL7Ybsd26Eg/VYoeNviJBZinRS1Q6IefBdy3JX8Nw7Hd4ZAJ2L2rH3MJJrJ
9vHsAKzLj+z/SAjUczklQzL/FDANEI9LISCgFiILfo8CB71RhKbahEv0yJQPiOpN
FQLR8JET3qKTH+JqQfb2CNu9MhQLJjAxl3DRecasSzDfAnxqcN2kHW8lrd+hiN3H
fnrqQr/HAhrBwfxOqFmTDVuCjQ7MkWyFSh2rPrs91Nc/20akk+gtDdNV+z/OkYc5
c1FBnLiEM4MuNNeNH0B1CNEe6AISK3/LPfni7R8Tm06vKDSu36V6uFJwDF05JAbp
CDcjDz9/dAGxxuxUU4neZrQL3oD9uaRwzO7e6dlZix11IpBHcA/xoQl2WPpwbIku
4wWbWaiYM9ct1dCcQApUGlTWHUth6upb3nvbDTMMiBsDSSpYVlNV2IoMOLYtTjBq
t6DgQYzPj9+eaGs3bPTJijzwOY0j0anLbOg8mNpvKSC9FzlyWygcipzYlPpkcJ5/
fNTWqP2O5LX0k6i3LBXhBIhVHH2O8G99kLtVPQTjUrNbYPVKHB8hqUuTMr9UVa/K
H4ugGorp58iS58RM494FjeEeN12zWjbmezBc3uyD7gpFeXtvEaKMQipuw+5IxWaX
WVYnpiiBJxGniOQmW/SJK+HVB5TZJx35GhTn0vHgMpYKiYL6r9KQZXA5wGJs2E12
lSwpNrDTSF1PqAGcO7lRIR30fJbC8YXTOEFGPCCXmAQ8EOSkXNEdZ+cVcocTrIJc
Tsa+qZRBHiRO2j8IOBRvv93xHk1526ddkH6NyGr6zmlggzDfdEMyPoGoeIJpP/Xl
3zWMCUw61U2PaedvDCfwK/Liuog78E1NVbvB8QVbQIyAkmYuOWdQvI3cGyqI37O8
WVD170uNbNynECh//9rl/t1c/WuM8ysYf7jpPj99wno/fOGJJaXGTTYTSn0MBkRX
H4n8m9FvO7hq6G6IjDH2WXwvw250KB+xigxxLMMNdUONafjRFWTUx+G5LbdSfVaZ
pMFftuqkwH7n10fViMLAtioc0LcO2ZJ3g8eJpBLvlU6Fvr6g0UH9Ulr6acOIp1RV
eYnUIzWuMTVHBEa8y5sVyeHNDw8BV7x0X6VnJvTl00DU6+iSOYNmWdQ5LBHy4/Ic
CRV4ndufwN9RlqXW7DsInRYjOAucY0rKbEl8xvveTWIeic4jv/wMcEwIqHjR+1Y8
gzM7o6lT0lLCfVCd22f5q9OZGXPdRgtw8ZXAWHiXimXGgJNXK6y+magOz9I0SLVj
gUa+J6VzyGkWSHqBCBcT2FJ4uvwNVsOK1FvSFBELXTL/s2Q4AB06iMHpoHbirJnG
RjtczDG4IAYJcAAcO30v++Sqm6k7HsG/1FWaqOlM4U51PdU6vcV7/fyxaTR6QlQA
sEiwOxm868ytgZoA9N3jrXa38EkssGxBMFYgvSO+aRKCqk+6WTQZub+NhW6ckeE6
P4S2fMjRSwJzMtBbJ6SIbzGT0jOuDup6N8ACqvf+2147uh39w0NjUfhhrieM+apU
TnBpDiNTy7o9bONUFaw/fKwByjforor01R9KyYAYs8+j7nRPTPvWD6YHCjKJqwxR
2F90EGCJf+2xB1+p0A9zUvfbpXGRpmkn1CKC05Uzisnz6JHHpioJGgQw9pUKfXV9
v2UEt+jy07s4+w8ge4bDTW8MYzVCwjVR1RqNjvkhJNi8q3g/CFIgSyW6rGYOIMWI
VnRD6Z7r/wyW/BS+rivLwfFSurHwluBCT9Syh2pKt+tGwfoncrieFLARUCHU4e9V
nmulsxXzzHJvXY2R8aBifDaQ8aFNoy84yUpJQkC8JaBwSUr+8enFdDqLOHazR6gW
au0DDEQF+QVHK1OTsQMJ6C+0w//ZNddR/FPJ83weWH2Qxe4IV7b9PDqu/x3RO+ZA
NSpOO/LHg4nbNO5RCtHMlbMBUeLwp/PNsnTc3mPg6EHYdTuxUW6UUZLxEfO0joDD
KRqnjmw58i6Ti+K6gayLRZ3y1P9ItSmKBs+W4Bei7HZJ9KpSqHx0kwCytVh0imX8
w9zKMTvlEWeuykJIIESehOEok32NCFdT35Ty2+sKIINP3vWseotXgij4Pp1Y9Rap
h6nTFdlk1DVXFrDWr85Qo3gubjgZCPf2ZfVH0Y3DC5Xmj8Yz4lNB8XiCxomVVmB9
xCLbiISzTBJBgVRnZuD3WqWKUBGxfGVwRjolev4QK9Sb92ho4NBQROnz4gXj2yZa
+4BxZeDu0dwHPB2ld1DOSZjXgw18ZGlm2w9Rg5450YH1rw1INXyf10MVH/8Cscy/
SQGVyUIl29ASI4YkGkQoxhMYSPiFKScugEvg8/884gPP9caUrdsU1jmyvpSxDmtR
4CTacz5VhxKkX/b0JDkfxNJAQU7rDfvWZxMfw3VP4zAH1DOChedXKRdV6X0bYH8I
8/A3R7fjSm23JU+uYBJdMiS+H/cTfQTCuZyfKj0oEYou9h7ZuYlWRahZo7KJWOmt
94zVmRr1ap7qQ8+ocMfFhK7F+tKblMmqyCYVPPaYU7GRo9+v3F+AAuhmXJ8w+ha8
jc2+wsvEEfOYSwrx+i8WtZzFiUNojct8K6HhabEUIImSdPUDKlXNW8MnXZT5raSl
b+qvZjWbj/omQo6a3CnDVaWzbryYUj2c3j7yi1c/8bVl2ycH8rATzR+EldqeURvq
9gWxFjW0YDOHB/3HH6/IElJyyhCdOKQwED16ij9/s7hi88BFhHZ+ZuryHT1UySzA
W3SpHLMfBzfpD9vX2IqQm37HqG1p4R68L8kcd+/CP3/nbrX/I09SnxpiZzal5SlT
vIedGVy7eeAaV8mHanxJ6rPxL2M9kSScBKRxS6TzRf2/DmcP6Tr5JoVgspSSzIQp
YHIDUzc2xHGo9uJ8VwaiUBxIydf3mMkY8bjDUlJYU2Y+ZGt7jwQGAJvCiww0aZF9
qfCjjJCZu49ioxHWwcLGB5HdqQv5oWTdD3+qfaxa576VLMn1jqRuqc5m9pwD+Gr4
6EQWdqk7v1zGxijlY5xqe34/I0wkZsEp5MkAENP8qZaHHWGskGBY2sbfcvX3OOmN
F/A6JtXhRysM0gzNkbY6wGlgW7Fhrv1qNWWc7FI+ZU7EMd3CVC/LdMfeMgnHYteM
FY/lLiwiOgK9F6ssry1EsyKmhwSfd6oS5Ybu5OAmGluTnZPhK9AYiCYhHSQpmRCz
FervdzDSm3/zYpYduQSCFL+yIHh+xpb+A13iPcXGw7WzfykohQGGOcxgDMZU5Q69
XBSC0lfjLQjvfEcSmXddkZ7VQxyqC9nAKbR/Rebynu40+EBLsJko4n3XJ0wPzoGy
PBaGOy5JK5yPuBomAHhOfP4Io7lqcX0yPMkJLUHOrdmJriNpAAuEn38+2YNi7q+N
bl1O8FaxcYjcwVw+PsZGcc0k5IZpbvA5A6lgLE7MA97da2DSwSB7fiwhXeeCn+4/
rk4/jpljGeYD5Pcqk6nIEe3kQfMCz9/h37rbcKXJWOiw9Q19COc3vu/0+ImUh1S2
/UzZDkwJMS6EGYHZqLYyGydKN+LM0JvTicLMawEk4ENe4VpBcdOgv0sobS5xWThi
Hhgsy9cnNHhOw+OCEa7FsFY9Gjdy38bzK6NVhmanjG4b/vayxWJiDcI0e5917+dm
xk8H95evZcj2at5HMcJJZQtv9EMgz124lAt0gc0aiIAakrFdcO+ngUV8NmnWpcfR
R7UcCl8+aLbfAJpxzjik+D7r9+skiDQpQIAmqe67QOlYBNzrHTCg0D0BH1ek1FyP
afeuoKxYd/sejdBq2O8Zr/IAlfSFG6fpbjdkjEbvpyAkCScrenUVEojTf2wRxWXl
YPMtO4EnQSAudDf9VFBS6+cA8bgB+KMRLaZm+bXBsLFAeXtRYLJcPVyirPFERzKX
79q5WbzU+slyQjTHRznU4tVm0zOSvy5sah4qZJfx4Srkm5QNZv3Ew71dVEglTxFx
g8SeyC2lIBmD3Fr4WUIoP+gsbOzMKVGCzJASZjk1j06veaiscc0KuDUeoMlLf+z4
CUDy3jw6IRDdvU5jtURr/vIN/x7g7nlsTPhxzYQn397DfmYrHxCcbDIPS7stTEsZ
f8LIcSB2ZHOVSSHkfk44HnwXGMri8S77qJXrk/z7iRp5b3utMpQsD+72/ifDoaUR
OkDwzsHSA+4jM9xf4YQKISGjV0/D+DWFtI4+feu4zXfaUWMWWVKHvQ/YwZufHGkq
zeGL5E1LZd/piLHq4MZ3dtvo3Hbzb5jbObB4p2Lty/yAWBnJ4r4YvdHu0285SwEx
P6aKwuybJGTkpyPzqkzyoraTekVxOAduuKMcrcL5xcEg09cS+dQUTjoLfxYevvUx
cHVDC/PuH3p9R2dfYrVuYoB38wMijrKxhdgaay16DNacmGmWZDRpj4K7JwzqPloV
nZfxGgoM1bW/jBlMDxQasHned1IMqkSsLpjyFRBjeapM5Kz+AnjaJLb8b9649lcj
ZfUWZHBuuMZRLKTmVO0QQ2ciGaUMNBiR6JkIlXA3KF8hWKVrN+FCNjsJmKz9Eq0M
pWPK0o0xVukXwIdGJKqCyTThiZP9vvfxjtxkEDks7/vxMrADzTAmg4gvbAR++ylW
6K2Vh/J6Kg+KZkYsJENj4tVbVHO9YpABAxuNaZx12H9k6RjbIYhw4KLuifHXTJby
890eeEW8HIH+F31fiIYMQp9YZZ9ifY52qKNE+J8VFUVZMj9S26cwr1Mb5CPW8IZy
K3PTfwGv2T9HnfdTlIR9tcEo9rTbCDurnbO0EHhiAG8QKjefvmRIDLmH3kczGdGn
8hlKDp3g1xST/H7uEVGjOPHp+hwmhwcovH091qqGCAFax8u5B1KjEBuFvZKnNXuD
9yLq7+K+3r7m78TEw4Armz3K2WXgHrGoRFeub0wm7AZuy6PMrO55gqZ6lAT3fcA3
FcCriQ3z9YuyMQERXKR1xw29geHjCLp7/pdLROEZ0apMxozm9I4VIvAdvBNcOSBx
WiyvBxYqTCiwULnIT6DTLy59rcb+4vLJtowihfyj9m2tkKQ4ELYlCiCFQ51ZxiV5
G6cO9lCv2Dqb8DmSQexg2VlZCa5LbQPUi31A0csYWeV8dNq3TG1TzXj+4HyUzv3t
czFdtYIiIfdD+50Z8FOgaktS6Kz6xKnPbs+/Xpbkss4pQlbY/3az0m8zLTxu+wrI
HHbch0fQjY+oiR5/cA4+yb0u04b13FBurv/lwIUpBWB7YTk7c4bzYE6vL5OPoRC/
iMCqmBQnEykywzLspnsD8sP4Pa9H6EhJ2e03hoEUvqMV8CCJKibIDiPBGFRmBW0w
QUIJ2HZfZLWZNPwb7lM1/2tDCIBa9KwwqyBcI3nV2DXMDPug1dhK9FJ7Bkci9qvJ
2GXem1WqKM0KPBfoaRhch6SC26a2x4R6cHZtQTWRnpyfXqpjhYCcG2j8WKcc3ZyF
eBvZorQBY6PFiOdIxoBTKI7CTffTGXOwWHpqGdlaMStT32FmDCdqvA5OKxcc77Gy
m7dBAfT7ZlCmehBUG7aTCjboCh6Yp5b/AYN4WBOYJ+jcKnd7vBZOfYCAGcft1M0O
vWl4HotmkUdOg9mSQuixbP+ZxzH6RrxKlmpzUCpwgF3FlcjOCawXL2thZhIUTVYH
K/Xsig3bknyTQsZQQsjmpmcE7n8OIKtgFAbHIDrlRh48KGks6TsqH8kz5dSVdWXi
F9oCga+TdcrIlTZoL5vpmpquiOlGZXJnp0LXdsOYZrFyKnBW1TNezocBq2cGDS9R
r7IRikzZ+8QCy2gR4H2GTK0NjfkEf2j/O6zJRTXr5BxAr/rjs1iniL45OCUJxuRD
P5KDQMTuAZapJduxjtqPAJEfjiHwNkVPnKK3O0SW6txrZoUcm+tZrNysAHn1vIjP
luxx9b8whPbvH64gEP6mXYha5OYH3aXegIi9ozqhqtboZ6eXNat7NP3IkU7sFeCO
TjBAOgwsRIlatZyZFj3gywaVvGPe9d7qi9Tq09dJ+Ok22XcnH+ITY568+PwOXGAM
n1GGFbbYpfklgsBgsFpUpUFgkbKha3j5m11W9iECAzhx50cG3Qfrk09ibi2aIH3/
BPz2/h+u6JPBnCZ4aUmr4Q==
`protect END_PROTECTED
