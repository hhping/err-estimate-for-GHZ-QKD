`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tRE9ImRD+gipAwFRXpR5osjtuvRpOLCVsprsyVy9PvITmjLLl2ofsSROgo0w1vC
QPzTvXTfnolQ4XOPZcaOKjT1DNCR3bpR0FXT6Zmh+aP6oTm5Th6xP0yEjzRwWtHW
N1KI27PipIFTHYCK2xM5eRPsvdxN+3GjaxBNtBU97kOhCTyEM8MDr3yVo5Xa8RzI
N3kC5qA94vqDKV82HPEDe35MUTQ61ktVua+qSpvCAlM0y2kLDbOEMoVtWAfM9dul
kucw/WH/D1GRk5Bm6bq2jn7I81SWRz+qt3UqyaYrvc1hzy/lyWBJVgEk7vwwl4OX
vEONtFc9n6r3HrFdNRfnEjt2kOMOXZtki6vMwR2WglsJaf9EUqaALu0E/2q9i9zR
RIaq1wH8mwjp+X06AUROFyJNjHF3s8zsUPmNUfsTulLJ0cJuMSiAn+fb+uWBBDfG
+1mlSeHCaekZiBcFC5S63yyy0Q3pSSjk6mqZyVDOJP3G/rSPdoIU/W9A/ZM+BumT
jxw94OWamX2Nhw6gOQ+AM4WP5O8ShmvMleQYuAH0n8GnTOXoMVh4hFabd44d41bc
k9vvxSOfaQ6bBYkBiwqDVq0thJ2yiIKXyseDWhYlxtOk5c7Wul72bRo4uRmUxeID
+4NFIl/fRc/3nHYHBgvK9Fj89tg/tCEFogNLqB1iMR0d18FCiCJnNTLsfQmHOoAZ
g8farlezjSj9/7pftKsmXeS5lmC+18XB/B2xtK18OOM=
`protect END_PROTECTED
