library verilog;
use verilog.vl_types.all;
entity TWENTYNM_PRIM_DFFE is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end TWENTYNM_PRIM_DFFE;
