`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D8S5qRxBEEDkV/Uq/GlkJkWrN2Kvpjt+h4AJgR5ME9mwVnq0+34fkFqedH6mL6Zv
efJfKtHOaAeaNITmE3ZjoAOvuP3q0M17UB0oBVOpBN9FsKi5j/ahmNB5GJFx/Tmj
hjz8/vd1cUtdq2IRLN/Zc5cIWYbb6bJmlNQlqE5QZS5J4D1XJB0b2o0FZ7LpT86Z
F2nULurqZzfi8bZq2dFXNIanDl1ADynuZ63/L5JaLKt4uezLG5aSgo8RyxFWmnwY
tFWX3i1FKDnGyeCPv7hxJ+NCHv8XbMkd+mHuFMhHfsEIdiNXzRt118ygcJuiZAGX
gOmZ9LTxI91Escur2211TTLIqVy61Dg+bwSFDe/GJyVTlnUZ/XdHiFroxZBOd1ka
V9ttKlKLVNVwkY3xYTJivQ+tEgnbC7jVK+yPLZSRbgO4jwhqst7rrf6MKw3lwy+j
d4jYCfPvbK+i30pQn4ArGVn5MkCMl0M/Muq2qAdVfSgQU0dPR2gymCcUsFTKHJCY
tNQmKyfTQkYxX/x88fkWudeHYZcoYv/ZMKVgsepVhlm0eCBxOnCgE1bZLZ7h2m+3
W4JikaRIzcH4c17gCrxVLc9JPpSDHIwiPAtDLBE1aI/CJ/fCTQubVpJUaqXqT4M/
uHPcSDkByvgyYDt9OH7/2lab/acAIaURxuMsPJ0AMwsnjnFLnpdMZBYVEZcybp4k
UCuDxhuT5i3dZ1F0kkNmuqcDMVZ+2wnPqvudSvKN+q1+EEp7exMGL9lsvlL2vuZz
CM3jlS1yEtynL5Mkg65zY2pLQuqECv6oTW2rpn0uo92XNU4nQyBz5rpvWMhBbbxS
FrrjI8KxT/qRGKl6er25q4vZw+yboS5PYVA301wvtWyq0GEXF+rrKyhEdajikhFm
FEIB4KXqhfZh7TlB643xxGP6wS6bh95ucQv9f1fslII=
`protect END_PROTECTED
