`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1FrltspOO8S+c2D/VcYT/MwIqRyWaFE5uxkanGunwHwdaI0gZ9246OuvevNA9QU
RnonfgL6LMBgUZjO4eNDQ/e5GSAEO0S/iW+fkKwkWTKGNy95fbA1MVi7/Z6JobP/
xnMnlvNUPviv2NWYTRHGlv/rDV40CIeROiBoXtxB0VIqZDLxfzTmCXhCIklEaIkL
B/HDztEZ03NtA8BRdxWwcVM194M/LY+9C798KA2ZUnHjGQSIvdks2I6gUBwHCyyr
YmCX3FA7LHyiu2MKHB1lRadITE34uIQcZ2wuScjhxgbB6zz74v+4ZVDv5gdQcIZW
EHwU1ASx1DqnVeJVuat6RqD3XQnu7jkeiZedhz6P4GMsKF7Jrfx3bPFwfpabLYRS
0/WMJZPArn2bLVEj+/OtFy469DdaANrT63wmARVhuvrYB7RzcF1jFC5VUPlxQ/Kf
swY9TCc//BDaATDJE9Ay8b0jAKeHXS/EaTx4YqjJp8Gh6P0KYq961NWABpMCggBE
/VXDesHk8A2u1RbJjh9I+D310VD4RglasNvRmFlGfHYZuuLllVgBeWQbkAuI0u1S
b/kgIPVp3T1jRvnkMiLjDC4EZZFPAHHsvdr8yxXEzITkkBV/YAqwHm29smG44IKb
CA4fXbic3LpdHtodJtsHlmvqKGEd5iZ8nR8sVsSVvzVe79QYWowWE7GPq3HyxeQD
BUawbY0yVGuJX/niLCfe1CcIpJgfuvppVNBYcoya9/AZpyOGb9J1AtxRcHjBX1YG
Nd/vB9lxuY6xSwm/3FJTuNIJUHc2Lb9RTUPF1Lw6bxBoG+mukpcX/stoIwu1T9SN
0T3X1fmk0D/zBG3HALdY4vUREaRmvLdvbiuZSdJqcAPqZbYbDMvSB1CSpHrbtwJT
avH8O6LIx5t6mOv3ZBfWEax89Hn5aU2gj/brggKGTgBUC8ac+68a3zkCli7qEet4
JZCYxV1HVO4q875HzfffcMKNOdq9UdSU9y14hOrwn8i/ZSISwquTaZFhop4PMwXQ
HzLHaKSbJq+Gvez8XC6E/BJU3V5gWJvuRPi4NzSGau11rsaW4+8Mp4PG9jVmThdR
MIEnWq7EvkR0KKXjwh6bRER9qY93hJuQFV0D3OdIRp14o2b5mv/Q9sxgDApKri9r
big9OX+S4lF1BOTeiuPBs7hbHPqYXNTC97NAPTN6cAu8TYebkEyRmNqtnOun9SlS
9R5VioryDIA5mv4EGz1vRO1uBDRhkWDAgSmQYWpswtdws012T0AT7d5ztijZ5oMA
RmKNjESy+JMz/R6Q5/OoFlNo08CYUtHj2F+cqBFCd41YppJ3CLvJj2BgYtkRogng
igm7LwsDq4th+hXV6eflvPrSt4Ok8IpU75odR61J9D1idv7Dgbr6IZgHF53eWvef
ZtnRCpFin7upbgnsfbI7EtsJsXofYSpufbG2R/ssSUf3ZmN0txygZBA8xBW+Sh9g
yHGRvueDZJ5VoiD0x5x4EAxDHtTlhmIJ5jno1TFwlk7UEt9BorYc3/C9QBKgufYU
kNwBXOeseLpsM615m2bS+vJj9yfCdwKgtYMVB/Wg4vkkdvSK24/FbwPHxTOwmLif
3JXIyWhXTSBpHmfYmP/OPXfNRyzLHtOZ9LQazjTKkcKlOXbqlVzTmdFLBuxJ4olC
eIYhPmrgkeaBOKb+LpL+vR1HM80iRoWVGPtYYBhRSZq194Fjgei8UBwKl34KSLT9
dtsqwjbRe/EDtbx7BqnXoH4ZzH5g2ccBG8QLPMZlTifgtxVlSvhHttA8kcmKio0s
nS36GIrPvBTl8oEE0V7rL4018zlnMQEcRwmJadO7u7ArReLTXeIu4/vuQZeQhb0q
PANpcvDC4y/3jpUBQJ6HDq2HlkT8l3iu7RO9zq8el2gO/Xmb4Aet/VuT8Vod0ZT3
zAIyOFgkcDMKEHC/3GK6IboFOLv7qnF/ldHMKYD4wkrPzcv2OBrgQSqqilpC5t1K
Q3e1rzofMh05LjgRsMDZn0d3HZBZD237VmQvuHr+akdKRAOlEVxwsHCB0mw4fgc2
JdwTzCXDuteoFRSnIm3qHg9EJvKSTDO+5ksBE+9hRDAlBRM4gpovkt7tCRBIO+Va
R7cwYngbarwsnaYPV6siAm4jVCZ/RGVn3qBGqP3ev1blO9JC5TIEAEFT05idbbtk
pU7VabcPA1U1saSu2AQOgbhWh83u8yNwRRhMCOEBK+CeNnpx99lBlQZoWa8zTlHE
BFRic1YvnsmvU1A99PuJdXtA0/Dgwwupr9LgU0dJTdnoT9BngQUcY326dlemu304
`protect END_PROTECTED
