`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRhe6mtYConmJbQg1/pFzo6WqSwChwowgkrkiR7FHnaESEd+iGSG9U2BLsbgHF62
MuZ2tZBDHM7Yyou/RqJZcVUrk1SnLbNFuKWOLX9aOP4halyMqeTS67bHrMv8ZsQu
uAhly4Y8PqAXqn32FQRq5WvVNnoVzNX5rCezxrluaSUI2GiKHYjuOEwk41nv9ixb
D/OaW6BsKa+TUQpl7TKfgswsmioGBT+c4xJxGSKuqCJm+RZbzABqbwk5xs6PiWu/
1pOLdT8JMdKusSejdGdQMDdgE2vExTVB21EfcZwJm8C9iwcXaJkXEP5WslDgdHCm
2oQFQCUa2uCJu1cQuQw1dmpnsmhRMGhN7OxkHoPzOVVwGZeaDjrYiXbrnYphHKkk
9jwS7NgS7SsNtbqdqxuUzq02QF1j0Y/Bs9lmo+vMyrtYaT/kZV25jlcU9kFmyMXD
Yp2sPXXtxtuh/hLQUYT3vHyfd/LMA1wYEHcXBc0t0Fzcba2xLY0YX0Cj/UpUd9dd
5xQg3Ff456oPmy4BUh9J4JAQqorGvqbPE+k0/NlZlD5wk/F3HaUENzXZBVZ2KTvu
95SYbqkgwy+QUlZuEU2+rTk274x93thATulf518hX1PRE382Bh+eq56h0UXGWPy+
TStgmEDG36+3orJeB9irQ0h13NK7i8OZkTM7GhBh7mffiUnz0Ix2J1Wlo99aT20r
RQCHh13HXEypym4sqzykrfs8UN9bcXwF9Jt3hNWmr4yASqfv6Kd46BTY/BTQLiHa
q69uMSXeua2PcTvoeMq3gaPKgU5g6AqTzACOUvq+PxSABY+3ooZ33lw7QyAA0j3F
5W7KTGGn/6SC+3dmlDjoY+1KnPNUP7T7wyr+m+1R6m/WpDgMpRq+neAJfr3TpI9m
9sFTFQPJoy25kKPw9x8nsx/EC47rK0LOtQ7ecR6/5YZmJCPq2iTNZ2HoVCoy3JMh
OGkVSts5e4aWV3Ao5Fbl+Dt2ev/wGX78YZA9maIuJXTn9f7TwD3gBiJNlWHRMRgb
u8fMIhX+so5dcBO/yKeb6LGnZbgSkjxBoSqDNJmPdHxOWHx4NWWsUEC96oH/+6Md
5b/l7ueVcY6PVZ/KzWfz8aRobDpEWWO1DB64RJOu1XkKPYbedDYuGwsd1PY24m2z
JNynOVrj5Krgp+rf+aXJlWkhavGubTvaPVigX2ZIpMiMT8M41yWzd7cBb9LWVsaf
AP7wDAgvt9CSKsbe/rlpVxWwT7XqUcXa0xRTdxX5irLM9IgNWjMaPT7QIPJFFYBe
WVp0r+wn6LxYVRN2nBypE4R3FOUMynKXVqL2raZKQhlQeIIiv0Wcb7T5193ATsSw
mb1hKeBJLgmHNdcWOPuY7uVdtRVe/nC1uD0CGblW4mbiJ/n6Z5//PkUY6uaaMymb
PnDsoiUcEGeeEypafZNvRRAB5V0/lcuyZU5VjVm5+qLiOj3ZxG4co4i38fRNpHwC
crimd6S0JWDe+xBf0vHd7qMwcx5rigxFttzwT4ab8dQFkgJDiTBLXywA7q00A+om
zMfZS741Z+2V3z71FDor6hZAX13d3bkTsJTnu39xLIrUujf+qZornm1ft1f8cOEa
xTqi/qKd8KfN1LhRvsOtZbq3n4Z3EpzWWugfKBVYL3uaF+A8U3Fn6SYLrwGsp3kT
pf0T/k/CVNJIM/Ej3dnDptEh04D9g/htuHXDRqekcQtGbm22X1iv+WLByTw7ad8d
ScT+VIDpGXEKFj/pHf78fUa/vKy+P62ofhu21q3SMINkCB0KfvLxmoY3L4lwsopX
Lt6LJtZPomik6JQkeYdLpp/ZyqlKIEcK/5uSgi48tvLCJcCl9hLe5zPsrs8yqYec
1Bl5T/ZJ8UMwuRz+dLewIchbHuw6W2VgY6X8FzT71Pu7ClDJrTmo2QudcPAw+l5D
/ozwEcRwg82GJnxdzbVDXVZ8BLfnvpeig3e8mmnD6dPQQC/qm2B0ondwtGV6Or56
v0RL1mrfxS8X9Df2jMgJC0OQ0P6D4DAMTb7Rb0DuOlmAZ0ksjthxO4LMoVvtDieJ
vyPvbEnV+bLUZoWtCr6nMo7QHgj0DZ9HLQVP/rO4L1Ay6v7jVqqZs5G8Jkx/9aWF
Akale2BBQEsR4MlUzovJSkpXqfvimid7gKQtYZSOAyZGCOqUV6KTpG14FCiXV6hl
7tAyc7bqoanbICvpjy/DGUTa3rhnWo9FGqX6bZi21D9V61U7o5ftmXjWZqnvb5fq
gtHuFbl0beL43aSBnEVfK5EXvfcacd6bRxnH0WISW+mB1FUgIwLwnlKDNxPCVwjD
Sq6J2PhPREcsGUNbPWDqrCJFBd0TUnNRazwxfdMTNMjLJ0JpmMuQ8mhSNN9w+doj
AKS3rMoKlS/QGQ+c1jWXcGxB8JNZwhUgDi48R9UF+WJj0YT8/UI+zgY4ijpZ3ESv
4zo4j8NRuu7V6h2xDxZbq5y834zxsTIfJ86nIsGyG3E9MWu5QPUkmMNmpXevPgKa
/mNFUrpERnQ80WT8COAAmKvhfEFyfrvX7SbFBaANaghMBzIR6/qyVtvPrXgQz3zW
KF1ggSaDEClHi85M9r2Miy8bcdk0H3oRaLmafQdRAlq0sGDybKlCHudqwbJ5bsbw
9icW6gm3tHO1Ea3nE2s2/QfiQbD6CJFhX0WIswAHd+RxV272FsTmR8jsxzt5P8n9
E8/PkmVQWev624in2X2upZvwBYuEQ9kL7FR0a78t/l5SkJdDjfsD6oHnRv9Z+Dc5
h2ErmSQ9R0uRZQfklRw2z4piZkljWrzbLRisY5D34IUBfyDvvEJOwmrXti9CFo0C
RTwe8UJPkgVzGxMpRGiDzNDoiHvPa4TclMy5kPH05pYNx7HAh2De4g1EQRfcbenO
Pd2vYNL+URjGco975D5khifux2J1057seJg6bOBM7rIlluB0TmCvoRd9QfQNCjb1
VnldkSdcdgNg4SjIV0dXVYGFq4IvL+XgfQTyXHfT+3C+AU13PnIgc+AzIsDvt4eY
lQB1Ltxi0xEF6siiU6gZ00hCDSjc5Z1Z1AXJo6lqAOFoyCbhXnKN5LCWFg0Ja/qh
/3lymxzGFWcmcvKb5MCy9Q+M8QEPlyY57cciSHqSKhMNlIGruTJgZPuZd0zpX1Z0
/hsljSZ7YysLDzLzmPTylEtGhM4sT8HMAUJefys04nHapUKbRilfDS4BL45yPPjW
JncEOKs0I2zdlgMv19m1XNfuqf/k43tc7Zx/QeKB26ZKgIEswLByN0EkzK3qAwAb
QPtpvEXdgQ2H2LafMkJSnggX1KWwKCQGvAnXRhQ+IsHViCICRSJJJMXB/holjIHv
rl53ehJ5NAuBYDYpyccbW/UNg3N825BfqpKATy/E111O6if1GOxCjPOI6tnRPbLy
XAXpjxM7x/kRJlP53jjOg63dXbwv0pMcDAqyRlvRJXU=
`protect END_PROTECTED
