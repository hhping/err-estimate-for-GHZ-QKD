`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MkLXAP3IjfVAIhjXr71xYq+wy3aLvNqa6x0OR2Xy7EdPagO990wUdHfVs2Gyulej
VtYfNpbR7xHVkxg3e7JDQbkUa70+znWzRw/6EpwgWcA04AG2KZTq8ZaxQwVs7nae
hetstXLUFAW4DMdD6B+avAgV8XpcPAJxp3C6faifXrwv5onCEsy+oQ6CkS/UNlxU
BSKlFGAaShYu9URnhHIZ76qxNPlekaNouQ2a8fKlfJCeIdu7m0at6Air1GjNRnYa
rYa2r9Tps7VZMVHoV3GSHrxHsO6RjOIAS9eUYBVX8GOCluN4B4r0vA+NnlYUXgja
8i1PjYcV2EDvX9OYrm0EVPV9WvJfkNlgmn9Zg67vjRsnP21UFniVi/2gSVPg/gp1
a+jfKwucNbtVlFxDmf/b5PvrOuev3wgQHRkUwQXGWLWrgsB5AAGbCIBoGN714+97
Digc/TgD1H3yolTvrSD//O/q9l5CMczBbfa0LF5q4p/a5c+4BRoxYYnM9yhaGT5w
iNTfvcYIuOMo8gQJtuSzY90fC/sK9Coan0zK1Mm8H+GQIyF7j3c7f4z7ihwSyx2E
5k0WKzdkw/b2x4XdAWr1yLYXy5mVv3MrYMNAijgnGLEIUf17OSAlOouxx2noxQbP
QQx+3QzawhYoTn6LaXzNwVZc5II4e82c7JPtOi8YnLCjldFfuFszuShh6efZwHTk
mv67DrG79aFmQ0TWKEO4UGo4y1CT/vKSWlnk2KK3qkSXk4y3NkTLRfFwbRwx//tY
hG3oZBSNLhcv9qZREazRs0aqcy1xdsi7lJLLy3pBcU4LczBhlokcB2J/CwM/vAY6
adKBzm0uykr/w4WlVdcikbPbTW+J36EPngDTD2FaLvcfphSNKSEqk8J7rAvpCGTn
7AGgDFeGe5Upm1m9dXKhEi+KwcfCIgGfjHcCXnQ68XNIv6NnMnoEY5AiLDNehHkL
RClZ5Z75wAnORv1ZNt6cViroaFKNlhUntc+wvqpAwxCFkah5o86NtCe4FxBD9dR0
s/iWLsycH8WwtRcpSNlTZw4jl/jCiwqkDHPcKCAkZfVNC+/9bjr8yvno4TWCmDOY
e2mYj/Tf3zvcDg+5yh8NTA==
`protect END_PROTECTED
