`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LBxu8UBL2bHvpHAhHZaiv6j0ashx88/SKeIAAsCRPNYChsQqpL20ncrvmXtYsnVq
bV9NAsWpsmSf0mdi9JSoSlw507vU2ungYTGK+BX/cFeByFt+SwApsazhe9PJFeGp
POoXwqiQ7YJIT/KInZExggLUddtbRGJ2tYL3TN5hGHdLAP8rRI9EX/L45gg8xNat
oa1gNIczc1AQNtR7d2q5DMTZXH4IzrcAGsJ5ZSnwrkefDZ0DKTDQH7S+Q4j2t5gr
7G0xbOJBdS/hhY6iP59tWjBxu8IgbE5vwiHVOAl5STKxjHpVBE3GpCPTnwFrtHzG
zT2VOeN8QaBgRj0DKKgePoQZkUSu1inxm8juHGVmbzBhftSqfJJOLabBRlRMxpUN
cfADnmBoOiKM6/6i0LBdDx4JhqMQZa0bpm4Y27f3vAqLaAhomFO/YFFrueo+iDnq
tquKSW65dvbF6P+UO6OaMQ==
`protect END_PROTECTED
