`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QimhsMAzb5n75Tq5mfq0Jts5w3++eI+7UQPIBYH7KIyAebWDtZq6nh3ovwlTioL
lmO9csxQZbqlINNOWbobQHa7zpK3ykhpZB+3Zw6afJgFcaBuSwxqVdhjJeN++4GD
8aAjpw49+9b6jktllN+dZOZdCi1YcgCuHfoLrH80IjDIN68b9IRgQjXUeKLejsqf
SLUpnTzZeUJH0SufcmixEYBahAqC8Cyk3ORoyLDafatydQVqeH4ADqhqfCnA1zgb
3paM4B1xMEq93gy7RQWuIuXs65/2AcWs+e7b+wdZtxXBMqmP8mrM9dEtCY0dIUq7
YEt3nkKpm/yfl7z8LsXX6kuMbqgwN+a8YBGshv+yGSTq4nXPLYXRPYxPIR30RFUV
FqFKN2OQLBf7oXsMoz3VGH1bq3w3IDLsw4Zk2qZFSrvbukII22NZC/PxNfEij3XX
Gjpm7IPfVJjRMgdQFQztVYL5P4D1WTuNeSYaKT6p+MNZX1QBSJ9gJa8rMbTMwJAC
QRBI8FqcMGmuifLRhPgFxQFbrCaOs22tdqqxZSf6426/lUxpyB5NDmz/85v/Fm3R
KjPWYbOlQlS+zGN9V/k+lZ6OP/LT8nXlk5AedIPMj8YxR5oMoDUFtcPk5Q+8V5aF
bPTid/gAUggTCYbdp9KEWIbzcutWtmqt5m3C1QwZ/YdkCm+SylW4BscM5mNnXoCy
Nvrlm7n0XM2jO/+E13H2VLdOwop8O2FaUV0BODl2r+GDPHSubvlBTyZUVRVW5A9B
iZSmdij2XmAr+tFwweNVIqt+778mZfH6KMzcD218mFbSl27TmBRSPDtOrXPIti1A
fTCf9l3v8zm9EjrY5INc6jE//tthluCW08G6evYEq1slC18dmbjYY9gP+1t0OLKA
DNblHlFYzDJRhwDD8H8Zvm8FrwyWAUvGik3KW+Get3frt6cPaL18HlVA/IMr/Ky+
WB/DC9ywpNjsx8VxR5/X+THm5HmVrWew74ZbgE360qjtwshSsoJEJu1NkLjdCqvs
64ofD6ybm1yxiEs5rgn2Z7k00HIwq8T2jdrgvrSofgg=
`protect END_PROTECTED
