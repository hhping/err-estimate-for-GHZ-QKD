`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+PLPMnmU8W25GtO9RuZXSVDxGUUIo8HS4YafWBW3D6Xa+78qsnJkXullK9pUYvbu
3rOcHEqlmPBIBbMSNZvgXhBATdj2eq3Y+gNHM2r6tBpUod6W4vWmGJUNbkVyF+mh
4o26leN8Pc+ubL2fr01+hBRr07KyFj6vEB8OmesS63mCpLpFJkc6dQSvWzw9/lu6
cLbiuVOVLfslHtVoWEVwbwA02Cze0N7aWjJbc0uS8LuqyBatJxl9oumgIBxNiuUW
fE3EyUULDSStdrLsm4/0/4SEh6QWUDfBDngTOR6tjTG+J1/ol38eXK7OIC3o7+OE
Z8PvpDIA/s2DmQkwI7kZtVRc7Rr7r0KONGCXyckh+ZzOXiWdCcsKrBrriPUWQ1ol
WLUB258MjO6yIwlhowSx0G+1XQIyIsICN95FAkxDZJ3gySzTuJ4Y8jO0PRGoAkj4
CM33T0YSYNAnwVr7ngnLe8jkS1v1Xf7FCEk53FKnh4At1xjUjf1L0vw6aA7m6uSo
wAVVyCrNMdWL2ls+2FkNVlB+7FlUePrPXEOFDsm3nDT17on2CTBcDabBpj1IvVaq
c58JMXdpBVomsaFPU6kWj12GFmSdMlXANNCauFWFEgNj5zGIkO0f3RqUR/K87Y+A
Lfqouu0g6n4s23+LnOk0XsNhY+w4nkpiaxvQ1BOqavKv2ybBdkHRoAjPCFD0rBys
zXWY1ABWJVbTapuPCRwNf8NHzDRHH/xvvo8+fhrwFgsM8JpyeVFO5jr+ze81ehKN
SFM+m5FGNF5dsAIRAz7RGars6VMq015GRZ9LZ7+H5EPEphDdSUYThD76pyaeMGcT
GYf6g0Uztpsso7IgizlaHIx3K+t3r+SRTQU45RrrCdFTtAsJbiqE1da4Rx9eA4As
L8fDvRxqePHAM0EAc+DnMuWgBjrvnIhiTXDJpQLkeHhv/2SAbPEtS8WqSCmPOLvL
xxKa1AHCcfXEqunkbdDPjD3oVrO59MVecGG7A9P02p9HCFCKLHAiB9kTXLC805Mz
GBvqhau2nmxoot9HZBSalgwOr+8O3P3VU7lxkq8VSWDnWB55i+MYLsnhb6jruD7M
b+cv8B9lfkSrW25nhX5JbuujpB3eRwA+wkszcGZpuVJgodovEDE2mkfaegEgKZqz
KBFVfGZ5UhHnTka5NAQRzDYCnUh1oZ41fWuTLzheLENN4gMS0BdyvrMl+dSTyeyF
i/P8E9xEK6qs+mQrAY/n81QED3YVeQo12x34FDcl8o/VS5vrPEQ7IAV0K4G67tl8
iUYi5GwWEFssirbRiBEI+oOmiq7BofrlFMtMUeV8M0f5s9Y/s/sP2o84hQGNxo4V
0MV2CJrXljWRBryGHBXPPdkZG2Ekjgk5efrv/xlsidUjbyo67kkGEax4ixo5pzCi
QbyTA7QkiEwkpabYJsYeio/3B35jCiHrbBCSv7tSGS4HViRIKRMudfI1MvTzWWwC
0gfkkhU8uD0O/he7XV09HBiFE1nJ4QXSAJjivCl2lwCY4Pt7NtWVAXvOC32ymwlp
2ZMLL4gUx+EwUFQpbfkXlwB/0hLPdpd9E94y2S0cQrnBSUDsWaBOP92IaWFMJ1uz
3H70ndzbZP0iwC/w+iTgMHq16vmq0VIo1XuJzna1vKZfyFif0B5+wV13UnNUO68l
/b2AwUy7QmeFmCtZRQ7VMj5VkwlukPygEBaKhCynVURjqqkD/qD+XSJHFX2vr/k9
+iFkmMFJkQwEN1iIA+Ej01lpsEBy8u9P9HN7OqRWjQD1XE8LxVwRMkPg6MmoWb3W
cGGPAR9ENyENDpPvNolgvpJGew3okWcaUa7coUR5YkskUOkIqt81VhiEpXlrLRQg
+R47e105CD0O/GeQf5BHbgrCPtmbN3y6XwdfAKEFBEhAnTfDJMM5lqPcspNmqUtD
Gu1W5m4b+FYS6tAamxSsLX2ufAEDS3waI7A3NOMfz4JnMfHuSiXlG07Db7Nyr+GN
GI3iWhOxAZ+7CcRj2wtaNoF6Lm9+B5UGRUPcLQ7IYi58hF2f9LQBvPvD1ugd4zy1
aPSHAKY0PTX44a8wnD95M0di5Mth3t3UFF5seCmkRGKRw6t4GGAjJ7DtXBGnjL49
lKoFYbEqcQsdSxb+fbAGX9yTM3BK3dGPDC2Kk8BvEgRIkNO0DY83ScsENM/Nko0X
/OQP58h10IVX1dlOklnzgUwP4RZ8pNjkxibrd19VeBYjFnuatz4O1ML3wWwn0nii
aE4fJuox9dO0WjuoqpiB3keNWYTOh8O2QiU4qfjGel65OPh3DPufouTTc3i7xZwI
GLKFDm7LFPwAgZNCwAZFXvc/gUs2Hy64FCrt6zelFncB9T0PGNhcgQfCUx5c21SX
T6526+683xAisTUm+FlzI8mqkt8Z1+2kxurU+yg1P9oTTSRVpqynebHrQ4P5K73N
32lneYT/qO6JQCe7vg3OfkSG+3Q6ZikbBxJdCiVd90DyO3y3KKD7/OqbaivKbpK0
qOGFgbC6N4eMjOzayXhiPCQBI1AEsSNbNtgWyI2S0HHSBYsTAQKT8KIRjbzzAXSq
Gs2hhWtWjDeoR3xoeD0RTDeKS2oK8XP0DGXhQWlxcWCYAMxYRaaU2aTW9fWOfp5u
bO+JqqoibtKrsaGJidYRxOM7X/xPjENfPYdVe+m5lq2QnzdtWfPkJNLUhXAd2KkA
UI7vv9gD5hXyG4pi4+IR85F/T6KyfYDREx3q11xdjlA4aq21hC+aSI3Igr69LHDi
9v1ZwU8vTRJWwbO+el1FUGF4MicqBUe9XM/yP5bGVmQZfvW2VGAQj6yXLAp6eZNX
WsJuvE+GOV2L2DguqMw7lwjzTRTWfMOvHWYmHqsmsebkrqHjYqHnoNCfLEbr8cvZ
ADYzgd6pMyCqS8GUUsahoxZvzLzx3g4iarK9R01SDmFDh8u/5iv6GoG9oPFQJJQO
EzwsCYNiUXB2KCf/S9dnTos4asFFs0vT9Uaq4xvej5KBm6S6H0gFmyPUncVWy5lG
PYKVc13T+Um5pH9vuPbnClY2mmaKg8SWHY9S8DLWLMxZm2iVxhCSdZHkYQlQBu+B
u0cgGvUSV6HBpoi7avhBcFhweuz3kxfygx1PMs4YQNLRsDD0Sw94VKggW4zZDJw4
2fIWSU/ewF4cBWrmGS8rj/rg8kvrddw07PoKe+nSLHmjQkQo4w1W4R+NNes/angU
2ZULDb1MhKA3esiVXHKdBc0XZirH5bVEnrWStjDUp8gR23qr7eOZzaF882vq8IhN
IAbfV1EUwAgsyBjRKV2Cn9HsYjB8SRbDH8qZRcbaLjVpmwZ6ZoKkIjWEan9KJjBe
rQQnnAL0vdxgmECAbBEG6LUxZv0zifKvEwOBKz8Z3GBSCeiipXbyVk22PXnFxJZR
K0WtTk6fEjT6MXOnwdwm+gXzxsxLrmnAlNXUmpU8QIC+FxdW/MWZrgYIK+ftYpzW
SPBL6b/xxQ1jcMRL7foWqAT0WQ89F8vPyYNWyhX9FD30KeEGSp5HsXvl+Uet777+
z5Xgtf/Pcj1zZa6irTa9xt1IuCy5db1GG3dL0TsVqtxnPOOqm907tq/xAvqewc9+
OL6AtaaIgglT8DKytVKrCKltQ0/D92lySc8Ipn9Ear8buYM1cbOID0oPqguBnQmE
pCoWiYd5p+hi4z66QnmkYs2x5Hci8iW2mAbRk2r6N5MpjA7wJrmR4s7g0UCBo13f
elZfkYOVuhHA2OQHyNb8JAkFWDMd97NvwVCg/f+XLU1LmKRquG5TxjikD/WDer0Q
fU5bEqWYpJvxv7vJNTTn8BSECFsTWDk/QERmHpl01aJ1bXPlwzgzXJi1AhAfAQXs
SAzfgqJRKwnlRDRHEEFAAgJLduE7ScF0BNtkuXhIaxlDWnIvJfZlVpVoT16ok5C4
zLWhZuN3Dj4qWKk0tuwFkGZlFzYjNEmrJC8FiyJJynqMt5gclRtWhCFTL9r7LACO
1/W6Kz6nnYRQHIrEhbiLyx1UZ01keNBhas3lBicFxHAcX0C8qBj+3kMcztEmXUIR
DSgs4cHTTTdEGRWB1rBC3EjOcnUGU/BttPXpwpgKDe9H3EVLnPFAcZ1kcliJEiyt
pdh+s3fgNQ95SCYmntyNKBP49cJQCnaCAcC27a9NgB6Y1fLW6doMGCIm8TQB/PpM
pBBhtW0pQEfhSNcCC/9dQa//TyE99MJkR3SAQysAO/bTdJHoI7KGL1rN4owvGjFq
Y6mfE810O38thLb7qCc3jAziG+n/piGunx7BOl4qN/i+7PtOMg9bviTszt5GkW9j
EzwgaQFwXUQvRYyHRigU+ICHqmph0KHfZ1RG+IChY1AgZC8hgeiUEZwFjlcbU4BA
UxniMSoR7fP7hwWW3+g71buM3A7XfzxNPbTbgW41NRFrZJjFuKmGHTWe3jsGbcwA
DgSF0EsuI8NX04aG7MUSYnoL99vGrMVLQU0XPFOb8wDsb/MQg7qGaF71qQ7SgQH2
4WQjmxntoI38vT33EYem9I5Pgri/cwdIT/oHo5bnfCBokKLeuu4Ok0I/Qsm/GVM1
xXiIBFEw+zpI0zsPIOsZ2mIHamlL0auyeJy3bHM+0DQ5VGYHEIrFBhJUjpQzjSzK
iDbDZK3xXmxIUL/e3Ihg6K1MtsSEy6q05HcDoZEY/tR5eCLT8eHzAlFdO9GQyT6Q
kzNjTG5ILOWaRXsq0rHzhzl591ZXAwWFzbruAbRT58g6c1X8gjfLtM1qMmFbYiqi
hrJFDxLyvjLpDv7/5VffR3mJK36luGxCsg41eqoGbdA7aqrMPBJCWixAdbDtoJMi
o7R1auDYuJd8oBEYY2nom4pyfPB1Tix+BkEZIuc5/2fo//P4RzSGZYMvAgVPR/T7
AJqeNMncUC/hApcu3QaXJIOG67+hjovJeivysSVaJPvFDZr29e9NDz355T5wPTOs
7j90FsRVzKvOBM0RYo8BKc/7B/Vyp1YEqF3fO4v+0Wcptu9A0t92uRJtzY8fvY0G
1w32s0WgN2DigYw4of24zn7SlJtWYIubd6zHT1jASbC19PnhFL1+DHpJtZvz3E8P
MYuGq1hhALd5sP8wTj1tECkRYMMyUq8va+oepq8hDD3d8XfBRLeBW2DzTuGGrqu+
KudzEOaikPjM3e+APehj+HJ6OSllA/onJFumsjhll2028dV886hI0A+QjerqW7VI
ZHJxqNnXuKradPObumpAE9d4UeQrvONNNJ4xbm/VTuz5G53yRlUwgqiJLG1fWrds
s+VkxzHwu7MJhmbgp3ns16aPr7m2XDlwVwRg1otSC90F2oX8F+IUW9/35rHU1EtB
DCOiwrOYx//rT0d6tBUReBmf8uu7SU2uL+Xvt6YORsi+thae8hVVpVD8EMNGUbWv
MM8P5kyfNnGnA7rB3/W3VWbuxG51iFVRhGFEnESO/k/4P41PsmtwaPBEHcSVtCJ0
S351ve6A7HbilKqIK6Jik8VBCy4/Lj2Lqr3xttp8KaRw9Rz9GodSLKfemuJldnz4
21HVg6kT2LxBbY5Y09c7TaLZZAjHmI/SBw0DQ4SKtniwhaSZmE7bwvblRkAZw1jJ
/QRURmVOMBdssVlehezjkYIuG4c7O8R7wdsozCx7hnT3ChdJZzTcfTN4ith8GKkp
vxsnJgi7elrH6qhpZ0Qt+4GBILaKiGVxyTqPKIbju4TjNUWu+qGoDQ2orWzc0PNG
6yr4g5DjGTDK6ZoI5PU8LvB1byxNal3+sT/NpFtLKz37tY12D0+3vtAVWvKoj9/B
mi1KNwV34LBDZZ+MYdUvuyfejH5OqEC20GBFSnjQ0F1tdGc35IdbL6DTYjxDPQte
X2BCjGDbCckuH6IjrZ83qKoZCvellEyiQs8uSLCy8H0wAvDSu6dfJOFvR0lETVnd
ytLvIlc/9HuZfxuJzOFI4XIujLG1cRh6LbwVxPphxGkhHA4hfhaUYl8JX/bLgv4T
bSJRv9+fhkm6Ak49IGHTc/sUKtVh2DmjFQd5ne7vYGH51JZZYKNbtOTomopSIo4Q
aJu6gnqTpgXVfbgQ1a35D7o0viYtGVyKbyZeeuF9AR3rtDP3MZUAnyanSuSIlo/G
ZUbybLBwAywjhirtTQDVc7YR7sWOkaqRLxmoLdXQ0wr5SatnTcABLw4XgAJ68+HS
vPGZs2Xv9qs5yBTZJRF+xLJ9KiPvvMxJHrDSOQrWwm/IyvnQlWbTx0qb6QhbpWz9
47ZSI9uOSMwhNIm9MufuCS7+vdXJHL6yKQ+OuyylEXIJYvBRl9KG28Ms33921MCo
iTqBJg7Smhi58muV/sxQphqlKtynm3Y6i3Eyoji/h9dm+fb3n0HDMpD5vw9O19Hy
9RXeAdw+R+Gyr351sowhYiyLcc0YYnixNSvpAo8oeNK1kuXKzQWf2smmHNTZdOz3
oV0HfCUzpHiqzI48lOQ5ponqRXYS0prJ7PKH3fQKfSRiax2lGjikrx0uyTeI7ZxC
OzBewScPPJbkriKYQS/mlG8OpzCp9JY/xaEO+J90IpTyCKC3YTrRhfweytbbGMHF
GlCF5UHXHFgfRJ+i891p030QzMIxuamWF+3lbBjJt+ws+E5cPnyEr8pYZpKZCzzZ
dYoz/wkTzD6EoEwWixnVeuTccn2qvMDhjxEcG2HllFsbmtK/Ri1w1/0A8Ua8Pwhh
bIgXb5z8+x/fxny8i+qPbeHjOQxeclQKR2hPYzOTP4kjItiLwrSz7SxIFbFdsQMC
CZXSex2MahD0vJFm9Po7NV0VSCqYpBit5nRJEXrBv87KibPxcbDFF7uvj0dEAo0I
hQhvJYgNE8hvsPHEoRzjkaSeVTTIvikT3EyFJnuBhjQ3adc+fHAaVk3Ww6WL8d5Y
suIzxS5uQmHcevlzcuERdDIHHQ/TYmqK5cMujKRsigtI2s19AiEMUBvn6UkYVheX
ViPdOS+L5xnaSJ4PlGQJwGf+lLprchSaFYXyZ0G9UfzRAUz1w+9V61qbKcnu3qJC
6WWrRGj+UJpY8/PiZUxwPA8yKl+2nTI5q9AT8+Ls3PQTdByC0Y5jfGvr1wmZYcKY
DBsXKBkfDkuiuzowwlLPIbtQ/9QgcKz6w91bFDlA9Nqs7vQEh4BPhRHpuM66dU6w
eAmor6/9uYdXwGRigL3Gmj6NrxX29snqclmHgl1bIEDn/CKTCPckhdzIqVCfPN1X
j9ivC6um5tjSIWIDiCVMCFiYpsxPED7lJHhSrx9K26Oi1It/3w9pUTTFtdTMfeNU
8cfQKz2O3JyIC5frdzkYLfFjipIq2Q5b7UrEXIzVL0RYXJKUlFaocU1avDnneRZm
lqx/7wOFRtiJYHSRh4NZ77O+vA9KwW2vhtEe2Mve+yuliuCGeAhYk8X26/cz1xWp
ooA37HeG7WD4CisIX2Wj0D9lY/4V4KTKDlzAsRjVHK1xTyPABrkGRo3FzPQuJmfO
1j0ZMxFuRlmEtUuVKe9fVKalC+H9paneRYhM4LqQhxh3nGXm6dmf8s4QsdRK0Wg/
5Qz0LI3MmzlEy6yeD9Jl4hRTkUowDspW7aYNdRNrEBQvIsCZGHMPWb0NqTe+IQ7z
68G1RBijeV8IIXH0TKMoVlb/oLCcAe1TorrkHW1eqmpuyIu9Fyyyx73nnc8brron
0fNwflhlNgvyhs+RDkptd1b4h/IJNM8Ifsw7MeUpqtlK+ZXMOnjTLzx+iL3k5Uaa
lu+0R5CjuZls73ZpvgtAgx5xrH6J5Sr28u+7nqAwwo5jxHQVfDwBljfCABEKFSLN
DADeSNWG59hnpyM63bfP4H3QpyDcSIORArpHTgjxKcQ8ZFCNrqnOveAhKiuzdiYY
B/l2RwftErIqwnkBhMdyDkLs0/3y3DD0FgXTqcj/9tDCeCMGS6g0rYDF10A2OO1F
w8uz6h82PlxRBNL7d1Bnw4q9gXmuo1XeCEO+kEbN0ihPb1+nLNAHtwoVREupu7FN
VqWUmlo8/Zpm7HlObylaRFtsomMEiet5IX/MaXpg7BZTiQF/AEvNzpYrkb5UiU/e
aUdTF1tz5gIOOc48Eb2dagSH3/X1+nwBuwM6ZCFxi/aliV+i4hd8YEz6M2vLv10M
K7iyW7q4HwjLkq3D4Vz6649ri69e955sIc+GFz9W4B59nHTm9tqL8Z33/BGl5Gv5
Wlr6KkJ03qRgVcjdG+AB+odFLxfjpF9oIcMgkPUa3IOgFJwHhaN0nrLIBBi1r3Vq
637dRdved9wgXRWN2aCLDnEvvujXpIJ2wQoZst8q8EMQrhL4/TzqBJB/kFE/sh2u
DygQ+436n0ENkfuWbYXlTTlO9m75notJBuINkR5+JXs0rKtblNabUUyzI3sfouSy
Btkui0rujMPGv47hSVI17fvsyVDMNe7S86YkKRyG+2g6wX014wyzll5L/DZ37aue
KY04LM57TFxIYfGnkTwYv5LsO1fE65ZsxiFzINOypoJACj/n7Z1hymo5WRVq0UwI
K1E7/jMo8z8K1zXiq1Ca4gMMuyjjFlLRPsoWSJVnkGBTsHm/BMqdmU8KdaEw/BOg
LIU+KvM7JSbpJM6VkrEyyZH3yv7VI0VOBn0/RyBzpqg3OGtFwHQdw2+ENY2b1wGC
DkOE/paDjRuDJSouAdSmWYvfivM3xxCXBaOjuGfs/Pc373Mi7oSAHjXXLnzEnVa/
yQp/Wo25AKc0mlYth8BQyfiWNACRsKwmzRpSkBYUNGFjwh0Lkzguo9nhbAJWaNMI
ML5B2NO65NRvhygmhdwFZYLoBgR57vhdJVZe4N/e4bF+NkWjN5291a2hX9k7tzo8
x5sXeFzFfVMI2qXZ+YVuwX2QWLFRkuK+d9adZOkGo1yl4s3+TWJzWRCY1+2BAPFu
OkmVc6cSZb3l3Kt2M5kGJALvXOoG8YkcQdy9AQfJeCX66KGJyr90GnaIqKODGaOE
zJwEAvw/rP23f6YL3Mjz2e13HPnwtgJ2gGpPcca9njgR8GxFd1hice9iqqXbtqam
SppMGS7AL63R9an3ysl2ziJyPeD13CsA8yiMR5XiHs0qQI6Bf+l1E7yZCL4a98bP
9Tf4Byr67Bgp6JwDMLf8o2TdhxbS4CiSe9VcVgfIlsfqC/QuOL7eI/lDKXFAIjEj
AOLd5+mDbPaPGXwsGVptHYkgD/BiXtyg+JXSHK+JMj+f3NCUfui0sh8GMKR7OfE8
mm8NNEQNjPiB7GCf7oun9UqDZuPbIQ/uRfA4I45EtJImyq3VXnjDMXfg2sSGlYke
4IUsH5M5xXNjx62u4c87lvLexln1/Cps4Qc713HCs4Q7115dVlBRj7S9jYGCxELT
SIS2eVj4G/QXJjCBqYfAz4f0UN3nBFZBaWsY70bnueODfuuEDHKV7M2hLJRshstl
F5/bwZd4kq54JbvHblPNiS5cLgEY89s+WmQmH7SZqLG9pqN48S+5KMEe8PWS8nlr
K+D2pllfhnj7sKg1LoZ8TKdTbejAh11ELINhs87yauwru82MuO3TrXKUIDi8JVfc
kTmL8J+HIR5QEvssEeLFCaSMkg1Swf/4JUKD69ydCXlwiE8ZJ3hNBr1tj+erYSgr
f7+Zk8bHTNcO34OGy7AVjjYnrWazndJ1vtOB9N7/VIMKWVCmqSLWt8MuaZYTTDY4
7tm4otOTJHtXIg+j8bAm43O9zzvUMl+g7axnf+wWDQbR/cJeHJnTPvZNijaACTA2
5O2BXc0xO8w5bLTvd3KJrHhQ68BI590K7c0vrdU+pWzR1QBJaPhw5V36ajMqFIWG
lpsPdAdUhCx7V59ZiUuUalJeuWCJDBWMnpLjiU+W6NS9MTCkiknA0YOduQ9YT31U
5DBPJ3xZpnWv5RTWiyF94muZOlxHB7/4iFJa24MUfEK1exc/dxvoDl+WrzKZGQy2
asqkmmTqTZ+wV5xFjMW4T3YwZCvuk9YHFx/dczVM0dGeVmODnnPDKSGHYfnodiJs
8hrl4QIBZVB73bMkkN0aiWdDii7QftgCSHnfEs9k1RGIhizNmPRx7UPoyTJDYoLE
6HEEcmfJ/SR4HucaRzlBU+DfV5cH8z7HTSpd74uFgBbEiF73bV2hfpJfCjMTzus6
o/+PunytK+Nf6Z8Z9aHgB8qmWE91vbCYVccOCpCes+c7AthEmZAqGlwBaPfIc0Vu
AkInOZWLk5GjHqZ9FYGUHWKtHqzNfXw8ePag3CkbVAIywyld1lhBMxvLUHmOO5rI
Nxnn9MNtWyOt+VfvlG0NCdGNyQ/w+4cvXfwPetZE2MUCLKngS306g4RU7vGJ2o/7
XgBgkrksfK6uSeTWy7MVFS82w5pC5pMfIMezBHDGWn2cEXRPdm1TbRNe7HZlmvp8
c9J5ju3Y7Hwu49FzJfaFjEG459hR11pBW/RcOowB7r3ADHQooECm+cPgSOK0CKLl
5xZIXaB4YTeYK6r92YgtunI7636GjtMkSysOQpn9K0tDnV37adQNeFmvrHWXQDcQ
+Bj3wBiw3vDPSiU3y2kc2RDVH3QjD2kpVptLLtP3YFr/36tG0s0FqJYbagAXY6gJ
M3QDEyzUBcLvJgp9K/+OA5kcDMfWglRr/sg6Q6TgIIlCrzTe4yxPNscytYeMeXeq
axgCve/BFNaoAE8XsiCFSLkvdO7ggKD2ZBUI6lxzrFiZmBoOUP5tsyvwNyVMtTpP
XBjAJMqytcKQreHe+8VKKlX0iJxYvtIkq/MmBoGMz++ByhNrBrKigMfVEhTQfUjM
ytoTD+ragTrjp8HtIFyjiNLHt6sKuVIKlD/HwxaAGqSuxsYIFP4PhvXZGIgpKFWo
49vVnIKM4jLzkB31awqiZTEloi8y6hRrTb7+iBBTaMesmkVO3jbSDL0ZARoQVKpg
2SI4wPDMqabE7gr7YSOv2gTBZOelgpjvgqtmPrS2QSPnS+TOHmgX1oFo/Jg8vWFB
cO7oDu1mxG6jppixmwORNpofCn5UZ+zwxjymULDorXC8D9kd7QBzQdVdgQTaYsmV
2BEnTr5aj8jocFyG/9ZjK/RSU0b8PMRusmP5iQ9IxdcOUrnaPx5ubKBL06G4BZh4
KvM2SQIDGcUSOjCQ/mLH8Uayof9GzEvOTkl81T57E+itCERwpprJxmIune/NBl3o
zHfDIwfZ2bv3jpKwubH4Z/OCtJdH6pgzPw9OBO9/P34k3l7ph1T26UHKWxA0HGEK
fpDaMS5DieGJ7P/epYVh8E8ivBJdaa2V52ep+6qMuTa5hIqQaIDaKSSVLGelmvVo
7gbFCODwt/yQEd9pEVYlAZxpEzdSADuJNRuO6Htz8J7x8PIjkD6jM3e8zeWCJeAB
FJdGFH9JF1f59PwlzGzSmTnbjEKrb6L4BxlwQ9wqfB26nqZCMALxRVFyHFt6lsrg
OKvF7tfZIny6sf6V3SyujrbI6xmglMPJ1to5crdcXmNHEwgW7q/ZGpViHLkv1vzm
u+cE9ulsXEMozDMNpINha5Mpuzw4aXIBxDRmQfHRE3lEFXrCwj4fhF3ybH/bqPjq
0WAN8H6zTvvVrXIAfOuJWmAPiX9vA3JAAvI3Q6pJlSqIjzbG9chNwpqPCz2wwhzj
boXu16DF1ZQV1MZ9n360cCXMiXNX0qybXWk6gAxPcqD6R9F9GR8Tn1DMle/7Z7lk
SNybw/4usOmgY/U1pNItkU/Oww1E9hSLt0TKxnuQsbWaGsNy8J26toOud+7hPxt4
a3D28lhpaPF8ij0knm7BLJJu+euRf+lch0WyqIYhEngNWGApJA7tFxrQivuYUSvA
KON4PxmDZ0X22Wp3WAwh31qX3DnGsgcQEYGcFfrcmIYwlgoJjIa0GLJSdlYesLD7
Wz1Z6w2jBjq/U739w1l64c1q7/NzesjfBrBN+qD/DEbQuFUCujYJgQ3WtyNcsWjB
zifOQOhotVAFPr3fX+Rj6Z+Ef5WHesorWC1Pjq1MfITIYzR1p2ldbuXBiYhPeD0j
4HS21ANWryZwPH7JCBol9+ALH38Cv3ImKZWhrVWUqPGY9DzWDmmd2jnEVfxO1BUx
qD6+KZO1hcSe1/ZaWww2J2oetVehAJqLscS8MpWB5S5pialdaVv5cBoJs7ra3jqk
Z3vAUi7I+qHo8NQnLpEdiP5mFBKmB2K/vj7/h+/Yv6zXFd26Y63Vfg3Rq6QG00ub
5wjQrwiJgNzb9MnajLroA8p2JdxDEvlw1+nkNW1GMn6E89Dqa3oV5r/IYwRrzBBp
IElitRLf+HDyZPp8Hgw/eF4QjL1Sg+U+GQ0RFDHCgICxZjaOtalvGBuh+9f2cdyw
J/GoGVzVjmzgaLv0CbF5KrbFvd/gjd1RZZHkzhelSLcnTNpj5bm4Ke6XcsGf+V7d
Q+rABnC5LfmOUQF8+2ZQp306DsEpRlp9M4z1YWpWdCaF7RPnnHDBNLd5/Zn5Pa/j
OIemYX8QEE4evVSy46LYGk2ALBznt7ks19HskiBYbFcQVR1O/SIExAIZ+eQiC0dF
+ZxA5tm1cUssk7SJYYJR9VnHjb/OQRHlm9LyVmL6KYWBDYeVis3f1iZz2AsBOQE2
MaVsMYO/UrZ6P9Cevom2XBbVyX+DzQtkf3FoJAhiJ/muv1uCdnR6bgDYoJQT7vu6
SNhrzpCVMDvv3UNgKntia00bPo8QULPCQ5XuWZ3a5Hib2dkR3UMuZiuDlLKUXjGv
kqgmkDuYkxzYhS01F5B2lcf7ocQmcQWqAw3Rrlui4UHWUFJQhMSXMgkUvO9LmFgS
mtFj2Fe3u4edu75Lp+mlqSLghF20OqCgywGTbliumb/4l3na/0CCgHrxbudoLRKG
v9S7vmqbbyu+ThD7ef0tAiQT4raqhVve8e9wxo4msKhoXDdn/sKN7OtLlIulu98n
jAE1YpRFFdm31nmpSF6MdovTFmjdBUNKJYbZRdIQVBlEGtAHCLoleVN9JokktRCt
6a3xnrqipIAFbjiNCjqZouqAiLqyFaD4y7+P42JLFI/HbsvGcgOtuSMdN5MIut7U
AZwGebyZ15vRfH2iP/71sfyRPLlo2gvEezCZqUQv2IvA1Hq5sfFtKF4j1k0ZE1b+
EfD6fXhunES2ym+7xqIgFEMbTNEQPugEXVIGFRp7kOPkcQTyWGvEoSafQXjNZwZr
+AOz1Ltac6cLJ08/mpZqtE7OzANFzGjIKqq1Yvp7Gnb3z/hFtNgq5ChucpvpAd4v
TTHITp/qid3ZxIJcdiJuWqdcEjBaJTXNW2YhkQG1SYyM+7BpWhEW7VXyCl2CXoKV
RAlKFvd6jjMwT62WWxlj2eJzlksDoYIXtKf5Puuk++qRxLxRi4Bc55LeT1SvinO6
ZYTgNW0Ts+a+C93fe1EhFGar1EEJaqvebrMSGj1d61wPVYOewTSdORoKKlaGCJIn
X9nr9rVjEfCGvuYoVlqfx28ktsE6+koX0aCvK2Yhp4mYTpHog2soC7ydT/4FFM4Y
6Ms4yV0aSQv5BDlfPcfe/FaHLAYUt9AXuaRLhsk+Pt0SyqL9RTrmYX2Y0tZwbP5p
SVnh57SIMfocL6dpm/5O6vhNbbyqvPwkznRR8Wvjp5jH8va/cEq39oPAKywz7jhr
kjjJAhlpe7YDZCXFlmuizAPVj/qjxxoeeEjKfa5OkCs7DBrI9Qbkiyc82axUbGnF
6YB1EDjAhZt8JYk/E2afg/U/Sx+ioeUqnQ6+RW0wJTIkiuHa3CRrTStifZpEEwYG
AM1BUpc9GR75RN00bC/w1htGyeDwsQVbL3IC/PuT5Ru/ZTDAt+XXfw7Km72cF1RY
k5bGAXmdDJg5g+EZy9tsjg+NCrYp07XhszF3CYmL2+hDcTcZ3paBN+ytmqrVGcrU
U2J0ZhbM02uUIfSGta7xDcAoA+FAgU8WJppRZr/5vN88AfHL2SG81XxLyDbRkxgn
hk94cIyGy3cM2jegw5FIKqefZkV30dy0OW70DUns6YF4DTZRqvs8z0LWrHFVHYIL
zyrlFltVy9bpu165w7dkM7D7+AdIxEcjf9p4etlIi0J+UC/oHVKVpNDPRd2FOvvH
rEYfhcwEo5jD8UQ3xXWB1wfYZK/1cHFRA7sDK4+cQvxThVhUGNHOnFZqsWSR34j3
kdVj4nMAa8X9Fqoxe/QcbKNOpAWOxfhlnSKXvnDbpQr2KxIgugy8RpCHXoj3VDGE
oPFP6Si11LxWITKRlpZzaUbZivZkXWvAbanUbxxLPrgmvx5MUHPPquAYfm9Daeg6
KnaGgRCPfxR9Db0BeLkNSnwBR/Fh1wqJnBdMD57LqO3C5BVGiICwppv0H/5gwl+H
IKhPBGDaIss3pjqQYhEKnCQ0stOLz6o5ePuZFes7G4uakvsGvzw3h0tNyYPiDAOh
gjKZTH77fmWlKGyu1CysSwavSAIRjr5xQU402KJ2+rFfSBbRECIe8jZ/xgwcVxJG
EHo08VfwaoOPPdgRzYOTSX9sCp1zAWwegTii8drxESAKETytpfLXn+08VgSV9Y7b
VR6HsTE2gJhJacZTYUTebL0DmiDUYbiNhOGwNDSx9nujLmtBzq/BGY80nEooYRcG
iQZ1qG0k42BJu7IUhBs1kygw1ix1O2RJJMZZ9l1HqvozwBkxH8aQnLUfWkibmf3J
ZPMHmtw3RXHqvJ+xTrauKsToARQh6FebhAnn0EuWNeMS9TV6str/et2rFHLNY/k6
Dsxq9MwOkq92zYlSorH2h72/wcglJHpE+X0fQx8WUHoqpGwiZHFrZlpAMtzpFnH8
odHmbSkG7/5ZrlH7nc3dYHlmY8y9u/4YVgzar8YXPuzet2H+VS8hO+CdwNx0Odlk
VfS5CYxS3F71BtacUeUyh0S4NR3989g/jvRYaaKhvXX8RQrAT9mYeV1QlEZU2sPP
jsibzchOruRKICJZ+F/pYPemIOAt7ZfX+p8Ss5G8Cy5hUigdrADGVleODpMCNCLy
msBTt0HK3XeHtG79G3zUTVxJzggpqgntHCF2XIMOLKLYnPz3RqsXgy1vqUk8S7tZ
DMnmp9YielgPecSF7Cok0nVo3/h7EuXNSy2xI6hT7TUehY/Z+lN7uCZzu1aghgsO
PtiNSl/52d8RFWVDTG8l71lisAIg6oKIW0rOGZkSfIftqT5sJ3hW/yXx7BFl0P4z
BxcGRTZJlKEjPWWyGECTRLvjb6y1k5DjkKY6Lr1Z4ihjRFFWyujRy3Fq1FD0nqEY
zYvxn69xsYwzP7Eta8+EivJEawUHWSAuRQ5x2XXKbA6W4sxO8UhcdLHEr5wCl8VZ
ejxpwNgiLKPzFSxd2ymdVOkbz48Md1dmbLF6nqLNUXSnBHtVPwk9/6Bw/hAGr0/q
gJbppyXBQe/5s2eoA1+GQBgQoChIGtCseVJsM7aYrjttgMvjclQYHuArUPgxAr6B
WfKxOS0/GuM4HtmUMoudEm4mEayu1J3GgafjO0cdku9bz0bPZt5XrODOdowIlFfF
TDx9YzF9VbxaxDKGhY9shbeNMxVN0xbofimYje9RqggRUCZl9umXHqhatKTuf8Y2
2W5DqlRkm3qw2Wcq9beamWUR2Pnb+ApRiy/EsC5O0PeV1vw9kYHwVM28YA0cQcWb
1E+BHDpDn0lDeHhv1NP4tmo5Zq93iI2lmy9bAuSCuELjCPoo7Gtmwofij14dAnIk
1jR8v0WTu5jK+puoxtvjFqp3yp/z2jXJbkSJEX4hP6j88AjZIp4HFIPOBC9aA+TE
ezsDvPAor5ySMKkoEf8DWopQnsVMmdPZNg/65NkiBQXWYAcuobFRr2c252FwUu19
G1S6IrFU8HfkL3RShkca6ULRamyyHeoOXkj5Km9jIq7BPstta8I5luRH9uGsNmvX
v3/P5Mb5f3DWxcNAk47dUUPrg86k/8eaCNJdiUClquDpoqItCAM553RmsZl0Vvg3
MLHz74rVdSUnm5xvdkz4rCetdAYLJCksJcztUboaMx/F6TGfUB2YT9Rb9bZu7YY6
W26FI4WmQPM/QJUozJJYCZN8NO0foP1/hJ98RX3UXLmPeo21zcJKl6cEmIUm4lD1
HUILusZGpNfywZyOh96n7kQIBe1g/MzTXK604H9lyz0JaXlAS6Q/r2Yo8FyWMXdy
AQNwFvSn09U/ZBbN08K0zjoWxcATUeU+j/FeTM8D4QkYDrjIcha+otmBi7iQdXpZ
T9C5w9vgyewux6F5kVAOR1yiqlTWwgwRbYtR9c0ue9Xyj1jYLw7RfateQTmsbEhd
ZXJzMatYY280VJ9GQHIsqT5INK+yW4DelOganX9Bcf4d5A3kt5P7Q5qcePFwV8yI
zm6e7CyqsvT1fpOPzVH3xq6rZjcIWYm0n9Jh7PuCvmOjwkq+0BzphGTilJ0TFNOw
9Fv2hEoYPaVwfIq3J2vBuRHKnvxpZmkyAYBboovPvSk2E77yyroeoK/nouAvhuBj
eDVjDnKQ1VICqNH+/90DMzrliV5Fn2lZup3ORoMd82x5ooGRbONsRytWzbimAuo6
t+FZPuudDxJjK9omUrgNxoW+tqS/LCSVT1Fq1sTZwDhOg9ZGsAzYhNuCV3s9nsN3
wpHf/cYCJU1Q5kiRFIykthF6zW0AZ5+iGqMoA7RT7UOvDMm7yZ+gSjBbnfEasaw7
8PaLZbacfIKlXx5DseH3C9yDyaGlyPCWel5nhSjtsoiVyACoz7owEt2T3xG3UNEv
4SJIFSTOPxkDY8cpIr8vRg==
`protect END_PROTECTED
