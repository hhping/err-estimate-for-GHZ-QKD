`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j1EyKNEsDt8oGeUt2CjhC2Fwe03mDnqlx4KSEvjzbxWos0pqxLEPAFPIL7CI4i+Y
ECwlIXfUFXO2cmrE+n7Cx4IR1M+AqcZk8bMCIZWxTvakOQKa21NNq3JcNKd/jBGV
uYNQ9EwIK9hP4ydOx8ZJDlJDWVXGRd5Ev9ipcTXP4G45ZTqTyqPMY6cYJmbRM7nW
o8Hb8WPqkb0ZYw8BNKrEt0V9LLXHDklkhVD+O57lphuxpG3U2n6KJ6CsJtyYvmPr
KXtV4Wc8htqrWCWJVEof2FJ2IDtIKNo/JIoUgwd9RyfSo+zsaqEYpIq7GO8BBqyn
bbduUgwljYfUO3qqM4p5ZDCc6eojavVZe18EEMG+LE5oaSFLFqvagd2yDvvYXnn2
HLwO5qeTQND3u8mo3gq6sgcklDW0yepCbE70x4/tPYym2tQR3Z7XGa5pZXt5IaQh
9CqI3TyoUf9BYmI8YHnl1DnaLC3BfJX9pC35hxIofJhAIxuf8aRSl+TsxHjII0uj
ruIQb+MFpzr2BmRM4uhcXSyvH/1NLPsj/oMbjLY16RPRLjDdsZtzNi8eN1n7DNjV
6dEw/gBlZKcJ88syTGZahXsxcpjymrIeW6sGM0D665W2Oih6X8Eikzzf5hREjtEd
zjKRZuRL/PeFP4QpBcq3kg31i3DqkDTmcly1DxHKdOoNqqOqkNft/DxksIxF8t+X
ctjCEipTNgUj+f7+Keh5cZyd+0mHS8cZqIb3/uSmzYvgY1iKUXP1kPEq3i0KzzLx
jmMy3tXh6Lithm2FdjvQ2iPC4ZvH0B2Qd0xcse9AwpRvmK9DRajCduQnbJg1SOlP
Gm9dcM0Ia7w9O2sfbCDnrz2IlsSzsw1ZoJTdtK0M9jBBgVHyVy77hYsjDSzhSKSQ
sAQpQn77GzgQ4kUFreq2hj0J21il6QiGo12iwqXSHbDy2ujvIATUysWLjhJhqL05
TdnnJAzxFM4LSRRQH+uEcBaFs61EMpu7hEq/jMSQllEcAhVyKRDY0/J9pk5MJSjF
+9qvlYXH44fDe70YM83gP/feOcxH0AzaiVOxr8rjshjUtk6jlfYVIg0i7o2UpVwL
+qwtIeVrAKy6ofKw5NahD3PdhC4MDwb+7AV91y42io854IKa+00Emn5+/2nBD5Qz
cRbQe3hFv4s7SaN/z8L3+2f5tyuwIrEaVOrfyTpI3qM11taOi/3J271h4lEyy7nb
iKWutNr9LFgCP4WeBzbnLXqyyt0Ytfz5dZrYorRbemT1PaigCo4Zu90P/wKmXsbk
aGDZNSXvy2jyXuaKIWaWR/HKqCZuS4vmhyUk6IFo6rEfcUdBVydS8GWoE3U/MZeG
uIVPct6acYhK4JwKv2UanWP7Gi0LG8YNcDxhcLHrt0fgXbUTAWWf9eAIG0JycL/u
DhuEdsxKyrxHGHDgm2qnUdhfzqUcF5mtgBehiTG/MNOSXHKbi9oNK7lBo3RFa48j
WTJp7fYWVCzX2P5M1pVzZQiqqOpMTbRyVgYyzv1QhPK0T10mGI1yDUvTfACEZgxv
bQuFvWrWpaFknefP9YJsen7gNNqF58e+X6KMx6tB2F/Y1/ZY9X9qQNBXmKBPEzIb
VpDf5ZxsdBSWbQzqT72fsQWrwW/KR1UNRN2lBpzWGgdq+0Nf4+H32cYlTnhfkMns
8Jeu1Zsln3DgAgvKvZdlisI2+Got9vAzMYVAEnc8bnfL0bdSSXXMWutAkedXCEcD
wue8CEUe2YglY2LXxgln2kJZk8sbVQkd5EMtOibkE7l6AtO0t09KwDty73AYTkON
t1uVKTrGuG6Xmol9TB0TpF83u4MccRpTo+nzIc6sJcFgKu7i5bBVwaIQ8AmGMkaL
hv1As6uTYFwOORbcjNy4vRpHorvaiIQZZEEbkR455xhKA7hKjRtVfabt8uTlJOpv
5hygq5mBHrQItdqwlElk9AbpdItd+lSxRawChhj6KX8fvlaZSQctKGtXGwUBv07A
W5d73OMt6WlCFDGv0E1dleLQ9at7VvWlCqu8YQd8vSjKKEoGzHBGb5yITcelFkcG
zqwFsdFPt05pZgHRlBpHMUD003pMGCpvZpKXuOLCuv0=
`protect END_PROTECTED
