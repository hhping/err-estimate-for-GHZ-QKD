`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A1QpGP9rVTRUi2tGjNd+bcMvXv83kU8gEArKRAtRjqhidzIuR0zEJ2jRXpx8IquC
xeIcGagkQCbymgGqTIsFb1edCQNMz+8F0t9/gI4nNkVOZS04ggsIk1H1Wcvxeolq
VG4GGOy9S3lSNBHTGgxb3EfHjAutvb8v/La+5KWuMq3hU/yGDcr8LJyfYiz5RpbW
471I8dVJjeM7Z2d2kw4jQ5ZGXVnarWBEJ3Qthw+LSrDFNYdKgbSh7KfDAMtxjHFk
jE3ymgnJ7a1llKuDnCiZ1jOPhC1fHcU3xijMjLUpVwkDV0xpPBecOrZr0BRQ2Js0
5uvkagG6UOZWh4qpsOwXajSHfZHjOHvTiyFhaGHAShyRui2sRb7wa77cHGqD82As
qt66sS+0++sOhB7Y/+MyvMntdRnwxMy8FEs5EXPNi7RmxfVwF50a5I7Ti0oXg7o1
+Use2XDj0Fcfe3/OWcgr6SC0sHvRFt9tLC02vhispIthGhDoka/x8V/fzjtT4tCn
OxSVk2DkHz77CNjVY0xKfU+pQB0lLPPC56kRYK3cStQbdEqYWXzoBZfKmbfYvvuN
famDiiUe0i3Xj4I+kx5zLtunJYDG9XFh0VOhVv4dfbxUpEtImfXN8W+psz/mGTzc
WbCrLgL1uzdPPyIqhdQQQ6hGGjbKNKUZ9o7QXIbx62AmAe7c7QNrX14pNb2KjiSY
1b2Hf1rlNDJYyl4bBlNe/P2WPlxG5QntIhKq4Xli2cL+BcwE3RgpX6ytNBjwPNSr
8u9s+3GzjyLyPtLzPGdktDxIIJnQ/bACnLpYz2Y3yGc6Obj7GrptcRcI2KZUvrFy
Yy3AwTZwBpd8+PmclvWAJ6T66KW4fSzdX2EAciPLOoYnD4q/6xAk+ek6vQ07tXN/
bT6MokVEkSNnzZraPdZGKbJeoF+1hT4M8xb69Y/LYx6o13nGphMRU8fUCdjGA+/a
MzX+5ClEOiQ8XOIIxQnuPBg7EkfL7HTiG7R20tO4wXvJvkelUlrc9BiQzXbQBTKV
Wa3A3SeZvjn2F+gYuFprgNdBhqbUMb0bWNzR8sDFY6Z8/KSlG+VYfd1Ow8mfIIZZ
IknCojeatH2xln2b5ztP6Q==
`protect END_PROTECTED
