`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MamI9irdTZ2BkTogcIFAPRcHHmXAiNBu5faCDHqFkSzAa+WH4AOwB59z0uIEl4o3
+OwPkIF4uMBiVxPxxxHaS4GtizWBt++7+7pxaqpKvHic+TSLCpV5uNrec9UzxRYs
24BlneFiKL8wbCm/nATqXKRPdPnl+Y4kxNMuP8wn06TRfkh3gslnpKsm7RxW3TNK
+67X75ci0g+5FvO0BGNTgR6udjnVLv2bKj7exiY/k9iUqRBOLRIvabJJbtdcLcNK
tcYEkEwsIfzilOY8klPQV+9HzvNJDkeUzD1FcWywfYKoXeQTHNJ0ih8l96B+exLx
3yI/8cStDGyLxtx8Sc/kX46UJwbWody6KHetMy0WNt4YMYLhAiVSiCkYhDhvSi9z
/eFRgU/qqM/7XjD24w8eoOi//GC/30qCYIDbmjg6GxJA6VChZwiUTF5b+9fTa9AC
lodFH2hOp5SvLvj+ZQh4Tn66PgU+5dW8nOQOi2fy3YnYp9cZAlhQN646Y2BwlARu
o60hUu5fcPbwqRKXJfI/CIHo0SOWjbPZOHISBLUiNO6LiUDdmwkDjemdZ9Z2chdN
1PzG+Qm0LeGsnrI9kOnDNZ7ehwQUBvI3Twrb3qNEhRi1+ZU8avLEps4VHzH21/Uz
SieO95T6tMdWqf6oewSVrkqLN40etNBWqsA0NwPe+quHqRhomG1i86XIKyclelEY
KcUqlL9Ygmv2qlsrYpIVKTCujMLaVtc9wrwH/K0wx6/YAK/axclnVa0juCCwJ8Ok
cBty/WAENLIOygG8ObJqWaTDnfu+9qH/XN5Ht6WcTJd+k6bsn+1JfFKAqFav6ELy
45G3YYM5Sl5E8yxuQX3xtJ33bNnE85Kt5g16vjbzGk5nEQPolXErjbo61mdlesbg
3eY/IRAdJA7+ySgQuzDJYuiIwWpFJZUbon9wul2tpLGctdJsxH3eqpTFbEcuKrCM
L4qeMMdGHb18ZlwxhKfjdXQnkhQ2g6eywQcTLwzJIKauCLcyoZfGNn69NIKsypOT
oAYuFe18IFy3cOwniGIyePDKkkXo33FF8xJC5PdmvFxYg/hVBmAlRUWrW9kDgfk7
M/WKLPG9T9BTM4VOXW3cs4Drg82GnE16D+9Himcff5WI4CWRR+dh24yc6NChpkXl
3vby26os1ZQe1etAHIiRWbJ59YyEnKcalr96beTWgVeDQ+3lW+wehtM7N8HCqifF
hKOMW+sGQAKNUyZHRBjT3dEEhvSofUVH0DUwVGMvBzOUsTBr33lmtRpUt4WdE4z7
8zrbwCmS4zAVo9d/rp0xQY71jIATxgyiLSR+A1gYgyAwoCsxJ4JRQKsc9qRHroPd
EOXSwIC7pyLpWtTpw5+0UGaHbnPaJM8OBtL9/DCJXkV98Oecg4qM1Pfn02dLiGAm
XpvegTubo3b85hiST6BV50Teo7gq8abY637nY+GN198vvM5iCpgU+lTr/CgGvL5G
DAvF+kgoPzucnST+dhDsFso+ktEOeQkgd5ifVe3HcYP7rKO/+XoHQwBWCuBPPkfC
PJp4FIqDDDzxQ8dgEyGmRoqimsCP5KcqW+Iil4mco5HjOTSVcB7nq3a8L4K3+JW+
MDs6Qi81VFC5RcOf3YWnXI1yuRp5mLDJAGOJxRJH1FwtUbVIkQW6m7zhAtQ+i+7Y
1gt7qw6LP1wAcJYkjr8oWAbSkvCBeLDbLMJDY2zeCFo/l/wGsux2v6TwuqyZ9kgU
V2s5HSrf/9QByOC+OkrETbaYwm/uULtaJrjBvNU83cqHmFR5hJCyMu5XwkhLWpcM
Nv63KT+vaL5ZVXM7wpfkuZlliJzAFcbD1cftlNq5lctsD9+NH+RSV0McUS7RkQd9
z47169b6xymvWfuvLKgDbikkodRckk4Xx8IAXl/ruIOcl/NA1QEHhYEbLvxqY21A
BZm6w/BRCmjCfEzytwOCCWRsa4zOuUVtjcjQUz/nqGzTj3+/2dAsrZ9DjfPtywbv
17SwivwclOqox7imhv2PlgcCSzzhEpsY9qCINdq39pTSlz2MKlzxu8o0FMlxmS0d
RmpLM/V8tvpttbH6lD7Ed+PmaW2+W6e/eU+Q4ABu3Q+B0EH6/IjowUd8cJtyx3tL
SZcRGVtTA4ovRH68WFMlC3Of2OwEDEvjkLHbEXC4p759mtWj+pJCMvGjxY7ex6uX
w6sJkvlOgtVZ5b/WEdp3PN6+oziv+E6TdIZu4NVe3QJD5FO1tmOxoXSNg0l3PiLZ
dD5QqCMoIMGD4z7DZ8bA/ShpS3aYE0SgaqkNE9hpyMxvInInoOtFS9bfmAT3LP6h
QXJOXfHrciwsJx1iOoswWel+ayRVRDXh6i/03np2R1TJu447blDtqltD6szJ5lL/
w/pVxFsnJzkZM35ZPcs/BuNu5h6frZK57rm9FiGSs0F+8AZr+4hrNk+YrVydJdl4
rdeBiAYk4+sKkfb93wxMrOLunSoIes8EhuuciNK+WO0YZTPjpr/AnRGa9pGhOUUd
FML6ja5gDQwkAvS/Gu7ZzWAwidFOUwhpg823iv//tGo2JL0AoAF4NcQqw8THfWzT
GcV3dsNNOIrSFzH2Iw0yRYDCEYGrWHqUutp2xNk8knEIOBdxs+hgW/Ugv9EW0oeM
Je4j+sjgp6L4ikY4x44JhdGhLCcN6ulFpfU7NKO9tWZwATT03B7bjfwASckfVIBq
9+8qLmTQgoVIEbQ2gUgj+KOgWpO2rsfGpKLl6leAcvFPGzGRLbLWOO4cIT53DP4a
TwaXtcnFov7fBsmcg8SiS5oO+/YwqpihxMu416WJcNjXGimEWl4rAs4cWXceAKka
nRAkUOWIbUoZahkIHppXW45h8HyzwoLN02RMcgx37y4IHkXDYrX6MyixI3Mt6f6h
zCi9oUt/HBQqILG/yU0T8b1N4qNmAWjA+alJvXwE67a4dt9XjBXAR3MHkntvqGFi
TS7dWgNyCODn8VaKL/F0khM/zC1/Y01ueoZoknw4C5kf0UoBl1y8rP4AOBHA5Qff
NwzGUgRWhg1CJWHlCdaxYdjR8AfnJ997gPVGAEN9mGDU+4q9P/W8GqG22fjW5lAt
kE4LAGjfxSkFnFgqGp2bIamYgbkfxNwuAKzS1iIokNBLeTmTzCubmdizapfTe/HK
B63EfaE8JgH4+ErzVKmbIk4rjGfanRTYjXuRf+LHnoMwJMePNxeG6sAY1O0gFJbH
47D1yl/YEZKqDkkX3i7JFQIEqNBCIOCmdhy/7t4fc5QPRhw+HJOppnpYfoX9KHkS
Cq9KUJ+/OBtjpjCZYfpH05fe5BCjU6F9bxYuOv/6ZGRTWkh5fWizPi68TzKCBgD5
TpqUHta+AJow8k9fdLAq18lJ/ncKqgZRdurlO1IDT2H0yUROaMFi1/WLMNMr8wdu
6UklU8ldNth8nj+ojUdpva38snzeO7HLH+Ru+FBm3pzng/xkBvR1AW/GplRmkkUx
x9Px7WduS2DaxFHayffTbxV7kwHvZkHk7cc3N5jnE3bOQx2YVaTH7v97yk/k3VPp
oxu5mkC9D/hiC2jNyUEfczZ86TFo+Vv3MFgLS/OOngp59vYNc7DxZ6TiMYOSqg5E
OlJZ1sRnxSQbF60jNkO1+IvWciGZiqoL9DTk5T1th3JbswNxIOcoavXpzxCAM1nb
G7AAlzCx/Xf/zy77kFyOjfogMeJjS4diruihpdNFKYxfIfSl71H3Bf2f7VZdy/74
xNhhs5sUE0oUk9T5bEIpFsd7IA3TcKPSEtWYSVYRIkC0KQvXowpz0KFLxSbY8A+9
UsPexhXrDNITioTUBWxhSMlBxrLMTf7GwIVGC4CZpGHDZSYeUYQacua724tvg8mv
4rsq5LOBDvkTnGyZDlQuMBm2d7K24GQC1b4fgh+8gvPLdMrzpA/PD33zMahCI5xs
f+8SIupXon3EoE2Aht5dqw==
`protect END_PROTECTED
