`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibCfQzxRI74a3B01FniB34XOeGZUmSivIxRxTNrK/jgdG5cn1kxkDgledie9oo7d
NckueA1jbnIovOaz+laCTGalOVYZLGcQX1iyiWCoHVRLuubDi2mX1KqtS5UX8Qev
rR801GbJ08tdFTlkSq7t9RLLztLDzz+aFr3BC4Zm/tpJMmzIVa5odjn9dyqeT6L4
uVty5luulsf9flPldcxecnWT299HuJOK1QXqh4UTdcPLWI8AptYGBMMskclX7g4s
AExn5L/iXxkaaUEytYV85rbsyCL+HtS4cBS+OWTJwXMrkPjdxvkVBy8crie1xvoy
UPsSJh7KJtwq9ZCdFknsRxpkUcv2xMBPYMi6EUdzRTTfpcp3wdwpCsDqOGvhcoKA
zqLK/JFsqBHk/YRQIAI/KFTHzqHSATMNmWnMLn2QsvN5Ih9cIg9sYMfQFPQ6iA9b
2y6nUZMrogYFYLTS4fsXP55fta90mStwhDku+Yd7k4uPu3ugMKXVELf+ID6OMMJM
aiNBokTk6tw6wuqkQwo46WeZa53H0aSQn30mMXc4aJsYL+Qvb6ItBB12VNt0VkUD
v8bue0l/Izmspafr+kYKEznOVHWXhI9VFDz3xfp8134VA1d24tQ1LnEgcwak5olp
rM4yGcybAO3d2+TdclrVEv/4RIY4hhP3Bm/FE6qFWjbJCs0VEd9SfTpsLQjFehkw
wkWYgwJJd3amZINkAZ+5FwxDnG5KpEYrk8zlauyCWFVkMc3B79DnF3AOynxheErU
bRtkHmJeSNCzBUixGpXODL+tbveINMoeThXR8vHdeOm0nuFXqj0fG3Rkh4vM2Q/G
a+RsU1RZYzdXdRWtWoO39hbLCnuOCazeLZAU6jioy+Nzn7iVKC49XRzZhQ79B+QC
wtw7uJBbMkVcb+URvbaSuL/QCvNEJgmP31Gz2KuX5tb1oM+acveQjyaDncaA+ew0
xTQxmGT2kL4XlX+Ife2q8CoP3EU7o0GHkSz9fYjKFSPi2CX7GTdbU68Sw8A9bUJ3
/QIfkxzndb6XszI5IEtb9wDQHxmJ/w2iycGtn/cbOKojdl7FWyY2odj8NcVXWqHW
WBS2Kc0RXTngZU/k7qToqGj/rYkPguBQ5YOSo2jyBMFDnEDW6BDRmqQNSB9WK4TL
kN5JLWxAO/tfnemEleigH/jnVSCbvahtUVNbzHiy9Vqa+YrMKCRajVezrcbYynVU
H8Z3FOYFxcHAdPixQYfKdJdML4JFOrk+yF+SpiIdtZaGglf2CcYeljYMQVREZaMJ
o1QqyjAtUL6p4RNuTXYXifvu5a0C7j1mDT435klIK3VJbFCSDnpp/2yKfgqIy1Wd
wc3tzIPsx5dDdX7ZCe2jX9fsqpEA4UFAvCqX+X7bqf7FeEdb/IlxSdJ1uZiv+yoq
S3vJkoKTQZVtaw91Wzr4XF3tNeEzvhUTLhodN9Eug6uMLpgd/v5g0+7+eRpbbGUX
`protect END_PROTECTED
