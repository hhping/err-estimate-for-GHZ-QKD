`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lW+k+INEo2diZUSu/y+e+Tp4lk+v77KNBK0uBdXGGfkNuZYoIarnx+gdphhtz3wX
hx8Nwz5chE7Itu7VKQsDaL8L2wIIF3kWL5/+PWtafvWDAFjW37eJ4qkrikY/qUlO
odyU1S/iOBFCyIVBivLhHS5pXzqBMI+6hyVNvOTwtSgzw/ugfR/gqDVs5zj/Sjzm
3vlYimCm4aY8+HWMBkHSe5eQvrlQ38KH2MBAhJIfTs8PqcxXbcbLD+yeewp3Vlcp
n/EMKEYqL9iLp65Vb8x0NZ3QteK1o6fam4EHp3efRlW9jQrLOz3doJGNtdx65z+f
eaiz5WCYtNqhNplhIbctFFmgn4ezfwf2exo5TuyOVnCup3wIWsZSGroVf5xbTndQ
rEJqeJesfMBim7OEGnOcDFdvlQ4/zMfFqLAdobplSTvNaaju3/EGT0MWsRoMcSGs
Me8K/mdDZ4L/jZM32H9fbMdbm6SYPs2O0bh0vF1TT8XXIGXWIrAZKwmZJ4ZlVzbp
3gQC+6YB0Z3HDTBrzjoFL25kBzADrXhiwyMFhw2zZ5vK4tcCNKuxSgoRx3G0lT/o
t4AV5J2p9r+AUSsjUUUkz5WUPgOnTKbG/Ank7eblJJM8+s+cJ3hep1hsqHA1LPdK
qN43wP5ts9UybcRLcA761s8LIyeIGvaja85M6H3MujjjmZTDKrAZf1pRXxKS3jdp
3eHapceJiH8XQYpsj6YyL1PjW9C2sRr1xCJsiVwsCEYmVKy38lM2wkSYXXKFDH+8
CimZ4U90i2sq+X29ukUTu5vEnHfPEOiFHPsI/O2Cw1S1Uk2wcKBxCPsjJzwuQl2Z
kVa4y5S1rg13j2lSVHdyBHPQneV7lV1pKY5+eN3w7RUOVQkZx/9vrJ2MpTvfz7qJ
nP1yH3S4TGrFBdcpVtpi954lCKuei3zSYvHbFXIJGWd3rWWMvkqJy+OEemwKJY/o
03d499QVmt6qsMDNshLYXdf4lC767ZadAeYwx2DaE0eizNNYCu8AGu1ng/2HxAHl
6vC24QcG9TBaVRQAoF24kuatSknEUj5AyYDh5taE1EuBd3NeRojj1Yk4NtBe/yvO
SjWgcQrTwaz08b/vA1krNZmEb5zGKN0SywBP4/kpbgXnsEX7jrXqCwfek55m96Zz
uFX+Jc8drOQSaVXQ1ivl75f6KCS18h4p3thGApzTsOj34vIkS1mSTrSg6jhFITii
d5YKis4AiPGhfRs5qbf/O0tb22snbnGepujtjkKNaTU1JuLvJ1hl0LVbc10wyrkO
AJ0dQivJs7tt883Wd914rL9cisDB0KWDMddVZAQDS+fUQjQG8ksEtAdK5kcF1uRv
I4osWE5iy3oiUgFSP/674bW15RInAmuRUCzSEqxXt3YLu+yW+Ske78lnhjtCpcec
KbTYxAvooCZQF7xD2dojMeAFhu+gfYdmpZdpm8rhO7tStkpIL/XhdViIscEgwQdg
w4aNAyhXMlkfWnZh0No89piH0RuVqesr8cv1iqtwcAIayUNXcCaN1XOddgAvd7te
jScCzeyDO89Eq2hAUK4SsUsYzAqMHlP3HDKuXFtWaVt8DTgGtlWGukPYJRyr1ZeU
UEJitfGOiFg5QHYXDvpq5/wVxvLrYwytJeJBpDDjVI9/SYhGvPWso0cv9+yFhBee
tpfcw93soWHFXBrLHx+HlWr09p40SU0sR1wUB13TMG63WBW9mYKDnBwpxwxgtog9
Tma9hXSihMQtTQy21wdsgczWy5qQbEQXHPqn8Td2Ec15Mvs2lRuMcdvFUKRMO51W
xVotLwb/D4F0fVpILr1UVHDOqqVtBuYSygI5AevLDlXMoYu6eKgTdl0n0S3XVuse
h4SPONLHTyuGXENp9C1bk+wf9GymwL0pHzxXLePpaCs9Te4VXAJBxMZWvTH2e5cL
fUNivaX1y8CkYHAl5EZMjS4ploAW3rQhOSwb504yR1VRiXDP9q660kh0wf1fnBeJ
EVep7gZ6E0Vuzu/uulogAHU5ZX3GSZwonwI316B7iJRwlDrOBrO+kB/kU3snEa/W
+vf0S7DADucYkvCGJi8h3ZAjLqe3trIX7jB3c6Sb0eiR885YW+PaDUHI2TepZnlg
utN7NuErTUDjkXto/UcOb3ulVGZm70QBTIOAgkSQ39PV46m/Ab+zN5Z/22k2JwWl
WMPzlq8jljwuLSvHeOQ0l2yh/FfT4AhVSYsFRSKZHZl7FKR99j+z4QqKTA+CtwM9
QTvbo9L0WEKdLvFemEDEhrwWSSlmyVYI5HQg7o6bWU8yF2Pjz/gy/Baz69Kgm4yY
rCNhIm+M+lbR4JIohu84qf9q2lGl30oPpjVSm9wlBgUZYp5q+0ndyGNLRB/yQUWM
ecdW6qrZdSB/7hoT95K7//NWs4/lYpfGiylfQItmVvEAi+7FEtA1H14D7mCuPQk+
zLbKUm5KBn3+l9eafLhq+hZVwBCgyomSP8FbvRnjcfrWPqIaNif6Tq4zcCrnaFcl
JASjbj8L0+/s7lPXQK3RDcoRXUS0KdiwA7c+UfUlbgHRV3AptzCUSkZdZih5TIyW
K+wkF9XYxJFNjyx25RyxT+ktd9dfEYwCWO03rc80MHSCHmUb5dl5bmhVxFB/A3D+
y3iatq2fJ4FaciPhZdd27jwDYVQnHNd8sqyFNrjMfVOtDDcHW66J9QcWCbYq8wEX
okd9QYUf9J89ADI09CNxNpk/93YrWkv6AoN8e7fASYBfvVtrTn1Fz+4aC4mYCt39
+qo2z3QiR+Zbad3KBEOMNCQ8FEhO2MYOdwPEHUi2/U2UDuwADZOP2mRKvq/DKf9v
qbxpTaGzfhBPWSpnprMxbEbYg1FLgZXWvwIqkApHL1TNfevOTfPnH0lbawzGn5uk
s6uzmQJowNBaVPZBWlf9AQEQMLYlkgnOQ0t6Ft84wjmIOp4nJGh0UDcqc1bnt8M8
QNw6i4KRIlQKAjtwtvJ+wz/KRibu4sYiU8Neg265zBeCm9jXfyNGlqLIdZtRSQSG
SnDDsQ0Bpv05LfOYk733jg==
`protect END_PROTECTED
