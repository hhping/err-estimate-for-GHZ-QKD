`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKKNDxUhyVG2kUMRuXMsqW2vzQ0iOyjAF3XtgeF/ke6RU/cSP4T8GAS7R6A37o0a
ZZB68A0cJBNbwW1n8cgaeA26YdBR9YLYkOkUqCrcKt7vFnGO7C+VkV5QTEC59R9x
E0CG5jIGzso+Nd4RaAIrNvucwO8rDNq2EvrSkW4efBsvzNXtOhCGucAJu6+40UNY
zUjpMu5IFy72QU+Ne0knFWokrX5x/D1xgai6DhKXaqbx7hRW6R33Ogli3oVWIPcX
bm0hFmp33e4x9n1YncWSlGuat5pFowTu6inqig3itCEYpo95r6+WAv2disO6G5az
frwDX3SZmVTlY0ZdEWVlD3fSpSMKQq7g/K2xwPD26ULURAmYA3ZdjOerT3oQHwPr
rn9OeAM3INFyDo3/ewXYEjPTZd3SoTfxAALpIHF5bk1FZ4SKNQ3BePP4G0sC3Q0R
00L9H3hvMVP2g/GUMIqXc95KkYlGmxi0QdA+XUHkyrLOTECasZW0rI+rfw+DjqhE
FtJ6g1UEeB/Gcw0FFISwnYTwmoCjuDP3+zoE2SM8TdU/kzmpbhsmlA1PetaJ7YX9
WBr2Ugq1RyKtFwu1O1t3eMSMk2YDc9r+dPr0L7AtWTLJYiNVHejsUc4qIgPkkX91
`protect END_PROTECTED
