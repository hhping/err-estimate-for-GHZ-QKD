`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdz5zhNU0Sd02lxEQDGHtdaB4Sc77lgd8mHFyVsU1xXCrdmXh+OJZSRh9Md1MUYh
JAf3DRhca1SlUeTOKubFqcMpHq+s5GYpHT1D3ZZHlwhUpKRSiagIfVAfg50KDCx5
oQKQ5iEJtjAXgdE2d9clAOmzDHTTK8yTz27gSuBpxXwLPMpjGrAxjyE9wR1iYwoX
uHlUcVGZ1VAAMEPTSIU/wK8ersMXMPo8gGvDXfJIwX/iBqof0ZpBZ/s06SLMQp6l
QSGq5Jr6wn2YDJlb1HCaFcC+Mxo1fZcm4aR8hg+aI5Ye12Iq7dKnIyox5DsqR+SI
qzf8GJ42qX6Od3ew/JwCbHrf9duQxvDNxSWh8Vch84S8RpSLbFZ99maFFRsY/YfH
qAfaS/6bycCTCsCIXojEKhh4KlB1YGCzllBLKJn6Q9I1Zl82hkxyEuOmYsWyCl4w
5IkMWIPMaNDgDS0qDJ8yel+p5RQRpXFiJHXM9HoAjIZJGHaFKki60xGGywn4m4p9
xDtEeCBYBfjLP4jOP8Tni19Zqu4L7oLLW19HKlQr/tZz/XSkLb81QRRiN32RCzkR
MG1ElkxOTwQ8P7CaVcFHtJOzki/IwPwyFZNpXBLrLnZCGhakSViAbEJhmpufg18B
`protect END_PROTECTED
