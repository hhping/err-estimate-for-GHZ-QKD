`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2668vJddcNQFMWvD5lXmYF3INkp9mhVJNSvYpEhULgWOi4zm46cfsRB45LyAM5J
2KOBHygBRoEzOAPhlm6/l2svqWb/1a6BKW8TXYBVUuU3lp7+847YU6CEXGl7PILF
kfVAmnW9vvt1/XRuSI0aWjv3KKtGP4nmVx6OVMb+i0k6eL1W733zUwUAD93RiNb3
4iU5WJR/tuc9nG0CoQ+yf6l3qc6hGGRSYqgULpoMnyvUyIrKeP+r15G2xAmFFJnO
nKkPv0VmRtmbgsaSqMoItrhFXKo6U9fpkmvwD54ggZejQ2kv7RfNQ98oau+POdLP
5oJ+hhA8/key3UMsd+l+/378XR7IIFpSb8K1wA+/TfYnwpYSHnan7BtZ2krYQf51
4MCQY2qJCVgrvGx9qkT3eTwF4ANg2+io1VNe/lqnCv4Ds+eHSb+dvXjLuQeta7ht
TmpkxWfVJ+HmgGN/u+47zDQSDdl3uKvmlWGV1JybgBj/5jz/ahdsUIUruxR6nKvR
Dn71P+a6QoZL6oGvEOiNlnC/nMqTG5fyS1siJyz+FkDCv+q1DBrvJ+rx7DAg29cr
1RvGCMSYA7DX2kXcIFj5+ZlX3giqk3UF5pP/9tWVBfpyVJPhrsDtJKfsPhnF9ZON
wVXHMd7Zf5WWBgwJbWWb4NW1Fxt4UueljWeGEeVEfEKnwL8ODKB3zsHWx9JsYZq/
hVItuLDPdC3ysjD1mNwPJ88xGY0C7f4R2FtTp5aqf7IFi+O1m6iakHlWuMW4kLrJ
kxHzCyKSEV13ED6/dQaMlWdbEZPiI6F4sJJlMOUVTmq1wW4zcSwxtcwg0japX7Ik
hfrcNRjxLVo+O59a/GzK2w306suhnbf5jRTz/F+WwW+vzwq40rhuIM0W7q4/1GT/
+kE2zMQnekFC0ifMstXfpmboM0vz6FiDhPTgzRR7oir8BbuGGfMpuXzncxtN13Iw
5UwpzPB+a1tzs9qUmA9xIUFWruuuMA7rBM1SvZbJJJMubdIOuK6YxgdhpSVp2jcU
HKtowlFor1cqbEYDqGp64K3rsHb3vLzcF95kRj9jBaqINHR7SIKxpHX1xzInmMF1
KsXdNietFFKKkkqMI9PK9fC1v00HZGJ/x3mWJtNkD9BRTkjFu+5AGTmaY8MHWudZ
aAz9Tm4NMJY1D3WY67RGv/MvJLJp6aAvJaN4uJA/GSm7cYQUGKXcAgFl+GQPzDuN
jDei3Iz2h9mP8IDUF48xzk7selT5n73STDStlI6l+O4Pw7DhXmQ6tJREbzDc8Hxx
CZ0KQNVDWKsFTF2P/+Do3rc0byVpUlMuqemcbYQu/M9zeqwQPf+5nRAz0uT/KNAQ
`protect END_PROTECTED
