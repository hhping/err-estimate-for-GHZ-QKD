`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7C8/XxbxaSdwE6dmTBgVdCWGkjAZFF5nXtDuwX9A6AEWOGghVuXpkfTgsW+v8u+w
fonPIEAOXN93/ulLGmBWjOCSiP10m5DdTQcx5xxssYSsUDBQPrZws43nRJcuiNku
JtHkqxTm8fh0S1+4ljnb6EUGjowIbaWc6oAPbgqz7jWoI9O0H+vXa4cdaiOgcG61
LwGzGBvc0K0OrxhWkWkGOIcJ4Xwwg80Yw0abHlsVxj+jel0KGNv94mOpF+9fxzVd
Ah92X2qg4t09sbcbvmGhmAqfbr1/bLY93ZVz2c5Hm7SXxQdGoUJgMokZjZlC9MmQ
Did+sSFDLMkXq5CxTzX2HUc9v9BzicEpGPXJAnHM8NSrzQrgzDbS5K1pqnuRPzfV
Ovav9b/w1Dxm2JNkezmZ1iOVjqMjcSImBGWHvswVRcrIhMT4YtIBtlD38ooyraEG
Ik5GRZOBQAvmE1MCp2ani8k1qpuOa/L+JGBz36tQDicGtd6+di314rq/BnfKHpgh
WqKhDDrO+bi58FPD92QXxi3p0cCpxSY2/qI9siua+flyKKm7sa/1NK9nseeGtWzh
WX1FK7t+eb6rwSKU8rhz704Uo50dm6rFmj4Uhw6k1HYsIfNdwDlw4hiwhkZ7Pnrm
6d4Ddne6u1O/oK9TEXMkJZsWLYDUGI+XBgR7u+SKFez3DvPAM66k7SmP1oVqz6ny
WxyOOle2t2tPvTJRTQh8wvTeqRe65lRrJjkzHzPjxrhBbL9kL3fR3oqi1uTxwjvE
4H3l6s8g7j3GE+85aS8XGlH3KNqoQ0fX5n+oKumrccZkY5KdiWXYWVMsIuwQ9CWq
Yh0oaRg52YRE7MQIUUW+uFBP1jW0RFLe6ZzssQvXNL7PP2lg2iThFzLZmr3/6Jbb
ahBtY0s42aE+O0xSavg3o+wk+cdhWNjMfGsrMY5+x5+miw80371d8KnnBvUXyX59
IyZmA53XnvIK2S5cC9w9VjoOKsnHMkmFqGEL4XQS2/iolIGlYOOAW689rfJ9/D9f
jPu10QmFEG90Aj92WesHuDAts3q5gjabW3P/r73UaIjYVc7klj6gMQ0+xkjTtnhr
9vE/ocbcFFP6Z5ARwtN8eE3eYfuTzzZOWWdr2+liO4SZgE2fObgxtqI6JOT0YKiS
loDnnrIvjEWaeV0bAZMlTKUgXpDMKTgjUj4OZuFV41ENjuAmdDXFxgQvCQh9ADJM
SWRLGWepycvZLEXuGnH4G4znjCl75hyuLgNVOVymSyPcjQ7zV84DvqLoUEjt0IfH
/gQk4ILeZGgZy+G/sA0BSBkqASwLJ7astCc5MqIMbiUrGNNLZ9AudMRT8DtJWHQY
OZ02lYbWbcwIR2Fz7VCDuA==
`protect END_PROTECTED
