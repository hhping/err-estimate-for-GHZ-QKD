`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k/xTm6Ir6m8J9uStTw80ZrqwgrHtfL3+SjfAZR14RtoTJDvhyzeQKXMW9tv+AcRf
W1qhkRchpiShkNQ8fVumEm+C9bbjzpv0Iq/41STdZDDV8nyhdCNAek1rmEP6xVUY
aYikDkqBg7UNKFtHAOM93ce8l43eEnA/dSwrSefJ0K2h4NRQLCyOU7m43Nwfs0Hc
QOZkwc7f8/b0SIw5OMtwQOP8iIjoZoJwze/pxZj9k7wZwjnDPY/adhtNvPfvLX8K
06g8PQVDy5QlyzdkDUKS5iHrtawVYK6YqfjIxdFCr0okS+5ah5N/15tJLK9gCPb2
KQrRyc196BSZze4XaqJjz3fWehEx6VF7R0adxr/exmr4D2lHd2n1sNCa3CYWBsch
FYH4ibACqliteIZAGdYQIuBIxVgMPWSD9vUE9qDrBeSQCDmUY/w8VFp2K84wbAlO
pKFamMQLGB/AjMDvMl6dgz9TMCZlCTv2D/yNEdCV93oTReTXpPw2Ibtio6mHt/GU
+weRwF9XNdHuTySy0UdztO4KBgoZPeFH3BZiLzaWaFaiIcAUaUwDYCq+oARzWOzN
f4p4KUEo10KzxDoiOMj2+vJb4rI0lv+OsD6cMyR3NHpIGEXFgfJjpWL/ZuBuClwu
0EBILdojyRNNDjhyrWe7Vx6VYEuZkM9wNcxUdsTx+3LQm4PVxKY1friFmDMYCPOX
NST78u9slB0YrU/+gw3Z8SUrO7S7K8VL8RYV/1Ef4+IAEq8S42ifvJyinTu25K0b
tuQSLfZzRLhvu5Df5AH04BfFs4oaeMP8CWnJle3B54xaex0W/4vfvM0aZaNEnA9a
`protect END_PROTECTED
