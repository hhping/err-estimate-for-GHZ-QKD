`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5IEbNixEcaP8S3+V2mv5aDBahmBPbN+tH82f7yVkknHCGEakj2U5yLfaWaoKbBdt
8Z8RowYi8LqE7rP1tiQVmAEWFTdgCSbrO/IVrGG3j9fFI1hgEKpdUD+/+aynZSb2
u2VNWnaxiJElx8LGn6K93+5ulH7sCGn+HcHAJz0PJv7sSBMaJpB4mm+v/ZhGt53q
IX/6pBEWk1n1zQRV+Go7KsmSLOo37QsCfGVmAC2PydhROZqcJQbxh17SE0DUbLLj
ezb5jwUV74YGQQdCjMB1SNgKF489PWBZFRomb43mF82RAze8Zt+CTjYncnnUEXA/
NTRuLIVvm+qlNQICp1h8fQYpGfXhy6o+/rW99oHu9DjduWVNkXz+/Q9/e0u60+os
cqxuf3WHODKHQk3fT74mYAMM/QRAJrJEVxW8ISpS5drC7EyMW1Jya+7bfzrOowPA
rW2If7S6TstVKy3jhfehzgcQ1DVYXXc8qyxME1A6gIMyzZUgR3UNQllW9m5ad14N
fW9YBtzXJSNQn2r99VAy8jc24lGHWjhle9sTc6DjS7Uzuuv5Y6xbBkWeQhgxV6fc
7Eau3mntY8eAMn4y1XjYy5LchHNQRpeopZg+GxYALWxUvpa1G3zdFa0WqhXdPJ6z
MleMLRDVTzUxXp8efchmikR+Fn9Nm955mcwu7+B+6/WuV4XPxdOXBb2h4DEr0O6A
cNKdNEYI2Yr4kU3GlXMHFIFtg8/gPQ/2JtoTXHaFGwn5V4OJ6dwv3serqClN1HhQ
`protect END_PROTECTED
