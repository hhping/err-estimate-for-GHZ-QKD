`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SV8Pi/lL5sX8C28VsdESMkOd0ZBzQQMN+FoJxLVmEMTJ1TwigIiL3w5GXvmWyrCk
0Uvzwtj7hnOrzvxyiEK9RVXc2vIslLrZXQduy6IL3DUXQ4hsDLZhDTwTcs4ttwqG
OmMsfBze41v8m+aoOBdYyr192Ag1G/k1gRTu/MmWB326FQskpvcscgAuer6pzUkK
+Jbdtd/O1JX9kRIYIMM5sP5g/XJg+jeHJLc/mpa2ZVw2vsTg6gBbZOtfjHcRdLHF
b6w8V6pj4721B3z3wrE8sON35nLGtZ2miUX/V/jV8ZPxcrY3ThX5OHva475yO3y8
Y9UyGi0iLFGCqzdNA+VrXaaPCHF60KEu88a6U10lzxYm3DN8lMw1DqpWrrHijuuv
k4yPRoqL3CVgtyU8eYmX2PyQ3iyicZlyzkcH8LIBeNSCAdl0wOY4xnGFg0eHdfSY
1zJ+mShPOGyTsE+DTyT3Iu2qabP6rcG6lobkCyJbBWHuY7jknJQT+hdYoE60fe/j
mVXneeQq5lU5QLoSDwv0axRtQYFlqN5afOZHoeWs5JTdBlgKZ8o5X34Ap+Dbjvm4
eLMQgjA2hg7kDMe0o4Nr+ZwbbUij5ikhwXPO6FZinZGeUEVMVgxkB0hf31t8v/TJ
rlUWSGmAWnhl0CQvCrU742boXu3879Eoa5C6Yv9mUNwJC0hRHAkAH5poiIDXYBU1
8jWCIyRRY/dtGHVMfTHVsmyJIzzSqkp32Tfmu8Mg7LeKX8qAiriQKzedBFQtfb1T
Lq+IIBDzXTuYksRTcCQDnWHTz417w9lrnPQ3N0fJNJY2vgjUZvms+zDXbdEzHP5C
X84ftf/BkL7dZl8JYKV1GP8brl5ePNQNYBVQ2kZUSnMqTvaxYBq5SAHZ1PSMqxaS
yW9Ie5OsXcCcq0N/RAasacjO4yFRamZ0ZgC4WmFojd9mMW8blb3lTEe7I4X9uT9l
xZf8cSQqgwDtkd0+F9MqK3sxkNvD6eX4VZvoxZSsaZKKRdF+KhkyKsWPGaug+Gj1
6eV1x1JENy/cRdAjbiBn1oLepxPsZ6y2uKqIB7GdSw+grfV8qif2HUTPhBIzuVZO
lC6BlsAjDpME1OjWH2k7hakgMxwV7VuifSaJtgGUxoJjkj1lkNWZ5NEHcnQvTtfX
sd8BYGYcIc/ta/ngSlfjsVXxHp2EWzuE9bm4tYWqxFPWySjlqSsC0NiUe9+dKnYx
62EXBs8/ARgNYji6W5ETzPhx+FPFg0H00SbWgJI3+gbKDwtmX993Wg9sTRqepEyN
RTpAcN8lDn4rCZNOOxxPhetaRGtPZNK1o4AW5zatzNpT20c6yBw82qnQHMZzFFUu
LlgiWcOIUX5/laJbrVE9DmTPWVZ4xSObiDD9E1pBkTrOEO/6AJefPrM1KGA7LYkQ
x4ImPy+aSihmEySozY/t365ymJkvC3Yk69L4krAb2oywGJkI1qY4SVyXfO+Z5NJQ
io5rWbgdCQXVRz+3KKaUc6ApYr5y6BLJmHhDJ4C+XTUvceggcoAz3D9BJsxTyMPs
evd5LmVmXg8OSb+3Z0SxuNzDwALLdkGaibaNh0ORUD/KvObU7PYq/2uzArAipBSq
V1beqJ2anPrjxtlkDWGPCRXW0cVcvdI/pQvh2C27IaA3arKFiClFLkoVGUoOi5fg
wJSTOiIFmUny0XB88KylFQ==
`protect END_PROTECTED
