`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUrM6pJGH15miAtIIox6x4reqrJV3ZhJAqRl+ivZnuYdbu9AScQUZgTnW4rdfYKj
0Ra9Wn5YKlGaoo4mM2yDTQgKgIA9tDwjl3jESQTJrIoKyoXaXrXuEFK27MWfRe90
SIXQf4Zw5SpSKeqIF+y53gDBj/2eTGFYltxzoMHipBptXoTxW1FmSYMmij4Lv15Q
X9tMA8NVpsKbllFqCmoreEQ8mktN0IjJUOpVBwkuSVyH9Fn4/K4qpoyIyEGshfnZ
rp/NpCgbrUY5NPizeoEDEKLY/KdcxIkeYvO7Ad+qovSmvPHAIZqmjI6N7K3H12mA
l25jlV4YJOE6lD3us3UHSmFmJlwmtOqqh9oRunBsFxnuib02mtQXFt/b9RGTPTf5
I4y2ufUSstjf7MP7YS6odxDphfSjuwxNWAIqz34y0azZft9wNDbReLSJqt+6OOvw
LkMLLByHAPzk9OQtx9R1Ud1wyXZ47fJAsL2y1XOIXoAou7KxOx72JDa89ZbnmvDc
ybhJiVV6iwx1XCWeJWRrtFmxW9djDwB/bXrZnkaZDwD0Oy4JPMehGGab62y41Z2F
PWeAHAOQUV/UdKGVAvV3rOJRWVaC4Y0R3bdwvDTrNpi2ss0LAhj14SwG7du/Bc0x
k4ZSUSQ78d0Ge+1HIDLwyUMV/mcs+iufjuVy9gVOVNj7Ngmt9eKo3Zo0Ua/DGAsI
k/kFPo88/Q/yqzcNsxJzYICwj2avY39llSh9OGi5ewToFYFbLG/6WjTwiYodcAQI
TianqbcIvhXQVE41vbnoXf6ddQ704eJxA7RSSlk8zAFJPEoB597u7mVUZgJKAH/Q
YIa0gQkauzVGckP3QOTRiSDgFUWR2Fy/QSWkWLE/h4g3VKPnIZd6vTvQeC7g6Lwf
PnoGLDucEKqyXOA0sYH5K+o33MJUnMBbHRoRG9Urk91t/obyb9xKy3Prnx6skTEj
cfk2lwYCOJxoGpVvzkh2CZ0KuftWhbIQgRLO1p8iZu88CF3+Uy+/bO2TqgWXDJ4G
R+ytnWP5Z6sqPslVZLwhbSGzp6yET65U9WLpN6lI6ygKDCANqSO7Ra8LJJG0dl9e
8qqJgSv+X/lxc6zHKJ75op7ghUa3FHcPw7gMhbdZpR5oh63knCzPXhhwO4at8fzr
PUBeou34LzaZig16UKG3GdQgLBu8h8kmcWQk+UaOngXjNh7rvbX24ixtIBS/c6lN
LV0k5cOsTx8QeYdbA6uekiuCFreMH20SZubdZl2hpwqQdmxG5zmEqiCF5C1/OHFu
m4tLhdFhArgW0Dmw7/okl1ZP11tLSBNp07u+ydF6DsHS6IONEbHZr/Iw/5O68BjK
PS7fs92ImA+os3KtcRSS13/J+MTab9cW0O/rndMFYcU0AmJ0EGsD/kDtXXcQjqdA
v3dNfQM6J1Ha1HuT8X8MPEZnyu8QE29iukaiwqOzvTgTK3nMvuKEHUKa6vlbwqXp
XSvGtj9u3C7wP9kW0zK7Rfp//PD+wwVLAFOS6QK3lAPT4ZqOIrQeLhgKbCE0yjxg
ULlWrm8IrqPEdWXLdjqLV1gk1L2tN3vlw3DQ03D5WUI7A7/amQHjABkbswTlTfEN
PuUIyaI9Joo/uRFSsWuXrgpmTR5kw+/h8GCApwIIIYi/mxaN9aW1Vllqi4435PNd
EByvSx8Q6nkZXHEYrYkcYoPoTFhPgNLfHX5IB3PCvyBUGJU1MxcU1h2IWRj4U7V5
SfgJvrkbytbt2wVFtbsL60LZ4C7tHaznffNcAwexYGkTX3gPj0aGLHx4OrioQcn7
KbWYJlahcZDd+Fs5aQWIoK95qYBa9jpHapRp0kwBSXhSPlPF3qe1AMj7vjERUukc
I16nadmO3xnfjrZQD7KFFBCoAkIHSk9+oyVIP8AuWR62B+kWHQfVp4TK+hyj9QaD
0WgQGRC36RKShMPR4GMp1k8IXaaqXtI1YwErYVwGDrIqudZbTPdLlGwQrbwiPgxe
3O5yuYNupPtShw2js7NhjC9UqwTIM+RQH6m+XLOqhd2IjB9RFCB0E7ljeoyo5GxT
iM6JATrorEFOdueM0Q86/mjCPvYjDLTbP0Vi3gNme5acyTyjwkL5qdStYvMRWxOy
E4YlofWjXA483qbhZY4hhbrmHoKRPpE9FvRqH7pAWOwescb+3B3hL5s8YKCo2gj+
qYnxce9VsJLObrhdbh/fWBDzuqN/gXoJZRRsfWwq8/aDeQC9Zw13aZVAdTGqF99D
ul7NI2V4ucZ5Z25sDEzaz4xTEB8R3RSxiGdaK39E0YUtv64LICM8Z55rXxMhZzuO
TDnLQMLsWJKA3fva8It90lzfvU/BPK7EzdayBuRbDJIiUACvKf9xERQ0/Z8N4pMm
E9Tb4L8jit8E+5bcgw1sQTdpPm7No+ydcNMNSWweFMgfRY/1qsR7E6SoUuzwVkVi
mH9X3KT4k5qlcSi7fFInTo2nQrGuLwFAfTIDXpS1gafSe+x8cubL5kl6t20OLrG9
VyKSq0eTsOfpwIS7tnfwb7812aOC7wenBxdN667qhSkofib/yJZ1Dj761j2FHGM2
NKvLhGC2sgc2WfGAoZgSklKjtrzHRvoeiDyuSCrs++7g1mrxarFD4UR/tnTEo7Oj
0Fp/Qk5A9V7xYa3/7EmlhvAXccYPIsY3PmWDClg7jP/wquE3YD3Dwpr5ys2/y5pA
6uObHhYyW19mBrDlaKh1ka841QaFqN/pNt0gC3OCYYq8tCGxVXRIj4LCu4LArOJg
IrH+/MnVfoR4afUHs7wiRldv0o10MDVTrgqsnQXYFcslHnfhRggzrFjXyZ2vqKUP
qpWuNQ5zWrOLvqL5h/n3Eg8vK//1toh2cLwSPYwiAP3a804M+L+SQbqzPX5Llnfi
LdPITwGGbh3vk8VDCQIIHLKqr44uKIG0HZigxFt0d3DwvdKJIcgmOLEv6z6xUy/s
HseOhRe19b/OUbaTkCsEo4U6zubc+1uFEk1JFfOdxHN8saNme+iI8kA3UwK4UVYe
zB9+BSVte/SQCuJarBkZRI17COZXt0Z4Wuqlfy7SG3tS3fRho0uEKpcnnHmMfPIO
Fl/wRkCy40j4m8l+jEQtcN+lC5vdHjp4Qu7VdCSnTV509i4aaeRa03OCHDYvquqX
lgUkt2wiIr8DbTVSY1s7aM8jfZ/l+m4IVxHiYhRF5o5DNWGV6VVSGPdAs9xKmMQR
dYeJoi85d93lhbBXxQT00EL1njTQJ+x9faSecVOABLHAhy/OqgEbWE7mdqin84JB
q3HPAq7yH10j8hByI8KwfLU80anpqIK3BM96r6+4Y5lZbh9IgjVcPH0lqGhbEkj/
8DgAj0IbhrsNH/0j2LPahSNOO/bx8PcsZjTGaA4cTCW7JQuac5It5FqC5n4AT+3n
VJTdxzaRk8xHZPasMYjXYzvReak6/tSjcOFRn3lae4Fdwf3PzLmn39p8TiqFKhrj
ooxhh+fucDvNnpJowBNfwpcvyAD4qTMD+TJSiBwjgykFEbpi0UM1aJEV1+MQvY6d
dkjKy9d2letG4NnfVNpNElZ0w/9vCQzBTyj6HSc9iUMtI7NItiZOlRLvjrs5WTMj
bFohpZBE8jB3NIOWScfMhV1W8zba+UuzE2vfmfqCkkBJfg3nzNHI1qReNJlZhqhS
vdn2KTRxEgyngBGVmOzasYyfHx15aTJRkGMWJmXz/Xbm9/oUzJ/H9v319WsMvv7m
QBy/mgkUhVndkeMj7YX1JAk0LK1a9IJSYLqmEZ2yHB47+kKtdQGy+H4WPRxb0xew
e4oSQYZyx8SJEvpXS5u0ZkgXjm5nipqqtdIGRt38O4n0sQTAZ3DL9wWaTxKFeTop
4SQFD0mNeaiuIhli1aMLntrGpWviXLYXNkOvm37DBujpcn1Y9CPG0t9j3/oicHVY
jaL0okHpbjq/A23LlwugE3JPM5icgwO1RQs+wbhoq5qIqmhM16q6lPBY68MRDLYH
FmFYGrl2iu44Nx+9h8nhR5aGzL5N/MJP6XK6DAWl37UAEzo5y6raeQWUikrMoWFb
om7sXlTso1POCG4etErgzzNew+PzpP6f6/joRsKB5ad+YjOLeItBu3rOaUUbsTwj
`protect END_PROTECTED
