`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
40Lx0zf8Vl5kZJnWVAtPJVxIypvGParBupPu7La6jY7mu5E15HIQYKMFktJ5E7OE
Vfw04iJNLQEy6dLBZ+xGjjdejHciR6v+OAc8JDGROgduCLijVS1Y+g8RU6XYGODB
RxK1ugTQvB5WcU8U0RQV3PwD7CN2wEhhkbtPDAb2eCz7v5NchyWacZcwMCPgJ3SP
d6u+dhxqvXPbGIGVEGe6SHdAx5Aago+nXu2eUDWyxcNs4ORJLIaep06LmvA9PLyO
9XN8L4TE4C9lQ6abMA6YJbZxw3lFrlR0iEVck/5SH8zwhE2pRrPx8szoqGVjlsYt
5zLLLV7Y/O1fq7U6qC0bbMkyLsShS9ivpDOO8eiPzS+qa5GgjEZwjg5ZTp4GXzsW
b02GYoKPq4ng7hUrkhXDudvw0tPWPGP/oKry1CIvVVIDmDjPFwl2tY5WdUuTFyzh
QmMnULBy1+wA/Cr9xxA5lTODcgigk7mjwYHzhWOs7vEkyIjyYgcqJLAQSyLo9OVQ
aHqcR+RMUF61ZFgn7ltRSkOo2mSwjfJM5LzPbQKlXokjnp9CI/uCGdQa/A2RLkgS
m1oP5kUCsT+AJcX8Z3/ExvJNNhBO/2tdmTglIy2hZFvdMTET2ExbZlvRRsAV4is0
k4Hv7vgMyIVtodP+sIMl3YDs5Od6TdDer+usr3dK3AowVB78UE0oiA6azwGM432K
7VfwgjjzqE4ZAlgojI27tQmWb0wYG8hU16izd9GOJMRHTBN4WulXWqHIxBSrH7eZ
c7/F5YvbHYr/FTsjlygkyOWkFqLoVLGiFiz5N4LHlIt1NZHM5Cn3ULvfPtcOl1dM
QTHNMGnnicPKf87JqSKZY2xD5bgYs+7hbFeuBeTOTD78kKnH/cFGgkesoDdU3oRw
sIYr577Lv3WndE2ZDrczqxmJodhjvpUq0uufkbZ8DHZ48NOSz8pAk3E8mGcveBqx
s6y5wtGPAhbtl40vUjlrHLlHI0r+YOL8lIv7MRI4auzKVqk5BT6QLK14ehhAo7JY
zWBPd5UEOVHfpP44HV+9oWac/KsZGpVdpT2/wI9mgxI=
`protect END_PROTECTED
