`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6jPjT4v8KGneuIFf5QK+sNOZ92F6/hDbPCST3K7/YmD+LdU27LG9YScNRvJ+II2
A1Cp0c7u2t+QGu38T3QwH73T+VSldqc/ahHjfpun3OnS24usouGlJPSRW/Vpcu1Q
0WNAcME4wYPeRE+kkFcQZPJj3H/IsqoCZ2xLMbLIcQydo0S85bUHgY27Gv4yykEX
gDI4MM0TwTPIrpIi1/K/tRHNt/sEBCkFltbPyF05UnO99cgBO2j5mu90mi14K5wi
ApvPz9KmZqiuCQjGAs6Cr7AeC/ImbfHc66QlBXdkVlsZXkKErbilBOEZA5pH913h
NLUIAxMpO8Az2e+rqBBkOEF7ldD7UJFtjjkoxmYxSntQXvmxyI3xByc2/ygCOzJB
sm2IVQZIXV+ZCiRzCvA3Jnoch/oZip5PQUy5Baq/rAsl7rKY1Oqy5kQQxyE7gCrP
ujIaPtvyRVuLZCNW1tIyYWCbMqcIeKm0Nzy9vGF9O8xQLfKlHL8Oqe9FHOf7w1uB
BFdf796YuPnUmdnVkmmSC1T7Tw5lPDLuInTSdiSQ2M231r8yLh1QGvx0ASgrKq8F
FgjlxczZwRslFX+HMAH8v3f5BkCPZzbRuJMrD/rIiOsMaW2b28t+0BLFKdzvKhgN
uCt17z5BoAxRnlgC9+Z0TW0c2OIKYxGXYXDYpopQod4=
`protect END_PROTECTED
