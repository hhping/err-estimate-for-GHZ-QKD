`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTyR2qIiuuvNZkwkAOZ7Qa8jduhpnvqX0ViQ5Ch9cdGsqWWoPewvuQ1z3sGxWW4i
D2vqEBMCuXVTGLyjuenBfGJqulQ4PgjnRwoJBI3clsohRDSknrer/c9ey+bmnCu8
pocPtCGcS0ejXxkD2XKuN8f/3vX7mNe8mxEisi82yE0r1Uw/o+o6+5qVA6Tv9VbC
HYcoDVu2nGLgg78xX4eByVvVGiZ9Bp8w1jDEbp5EqjAH1+igzSAJaZrRaAwS2Vu9
PCMHD1H1nJF4+DYHaiqSZBpSzWI5xip2skWCwtw6SNCFEjMF2wy/fxPCm6cTE49J
PwihqZar76rq9ZyoEvyGDxGXuEI13GmYS8LPrDG+xQNc/gEaf/S5mfqgSJMczqm7
fPiRG4v7bQyyY4u21joKLEnTDbOiZ1xwM++yZkdn2G0lPVJ7Pr3yNwcXAlhYw0jW
gSXpc4yCpR3qjzyedfg0O+dMlTiF7SRwHLVUkhZ/Jg2Tw+RVX0BxZl5wTbn9i1uo
jqCUv5FtFu1ZI5SISzplObE7VxidX0a6BpDo4VOzZw6A2L3XlZJeeS6qQYC9oIPs
B0X/Y5iIgX7F3gRvou+uL8jA81s0i6XLgSxEXY+yMlsjdXF9JnFC1/wTC0jvqD+O
ko7/mq3VF7Pg0OXLB0dMXlsjynldUmCClpL0cq1r2o9cICmikg14BS7AdSQ/jD4U
W8Qd3NPjq0Hk0y87CsNfUcm5tzlZ+90+MLH4rjuzkgYs2gfu8xerO6mZAabCAkZe
liikkvYiKuXZ2KuOYjN6qgKHFlZ65KCgx45pm1JGe10i4iIFunLhgDj3+8P+5PMp
nqNWAlOLKeitKmiFS8cuEVXhFoC6xX4UyBQLtE2F8t+iXIsI1t+WNeqFPkyUo2Yk
zjp97x97ZwjyN0U1qH4fLHxnsF/hNM2srT65PrNVkojDomMmAkHDgvpuW28z+WBn
OqrzY8hrfZINGqXCU7hItN87jjwLCQZP9iVZbVk+fhKfadCQlQhge/2oVJZinSeX
61WkYNwt6mi7UOegy+Jg4SKZoFWkFc5ft/LfbleiDbNYDlCo6d/LPEudAzK7t4tA
6/n5UG/hSi3IrQeMuJOb/SI6ZBOzqfQNN+0EWiX3EP90QT1VWwsuvtj0W+omcR/J
Y2+8/FoIXxd5cHR1d2FWgESbk5YketybXPH7/R+eC3zxH24VayHv9kb0mNVTN9Rz
wwxu8ZkXtcR8S70NqI6+VatcJrAkikXiTZSMYy5quUOM7WNK0dGRXpZGsA/BDPcI
la/eioGXVVJGXK80RgQpxj+TGcHr8ORYQnahH3vvviMlqKbiwXlgTLs73paMNUmj
5L1IDcRxZxlU4EDLPiui8HdV+AoPBhUtZ3Bj4pZKrhp2t0gp8E3TJw1HTjRcBH8c
t3QQCRfUrpXSVcSUR7Y+6/zw8HQqRgm5NAitWcppTFhQKwWO3wIZf8xDnak3d39T
etLb5wz4kdz1Cy60rsYVe3myvJZmYHK5i1WVeJFouSt8nZ+Nnpfpo5hEeScGTn/v
mWELbI1APgilqbY7uaM+l+XBFy9hY5bIrw+HBKhJR1ivieSGek4vPK1AEXyvQWxd
PnWnnrdUtBMxvpYh68zw0NB6vHoBHZbXQbe0jHmAdNaR/8tndV5daDp/y7Cw2SwI
04is7wLhBEj3pAzBkXwPqC1vjZF0v5tvj2/1Dt2fXDRakFcaRro4BFkRTryxMWGC
63jY4Lft70ZYPt7+Gu4F2u/J9eWO2PzJXMQzsAPhLPhBw3ntXiHivW31u7GiVm5I
7falWy4mxDG1oHhdfecYj0vwv3NEo5cDTiZBh+sXvW6uuYNHjjCMGv01175gFpKG
jxbsBpIZ9jTTOvrZz2aLfdcbqnB5dotzAN3IFRTKH+olr0wl2kOqBy8r46hfasjN
6aX1S9wT4TJvhVMMHBHytDp/+tC8X8w48rWqS95PJcP4uLaXrGuAsdPJZUvJOsPI
/aB5UOYEmM7lkH2n1SK8SZHgQZ6rIXXsnQqV5QvtKnFqRTTVegGrpx4Ew3V+TNgA
ahXcTmiVLzmvKoMHed5Hg4wpgcXA0pKTrk9MZWJMaCCm38byE4HNI7NdJBv9T3A2
SyDkuEm282QBkNImK8ZiAk9UkL/Kpm3dJuxy5HSwUPhKFi8rih7YvZa1pyg4Nza7
ChrJTvg2gujAxF6sKO/5moENPC06leBTQV6pX8NBe2y1ZSW0Pny/Uhw0RfaaHKMX
NvHSJRPTm6uGSojuhB25ZH3cAaDL5MsR9QmOQszAxZ2pbQOSYfEf9QrTZSJp5X9x
PmRKE260tiwz71zAAgDYWi+aqZL9YxqU++Fd0qnfpPPhKNdVXneDO/3+Bojt7RyI
KfiWbFf9cADU/bkuhNXE2Kq2UivRgAOWGafPRAJC2j73bVF58OjzR8GhKLyjb6E4
3qoBLHvROMNhVaXdXa3LkHRLNJ7n8oWIcuGAPvGRG3pcYFqkmOsfnrQRN3Hbv0f4
7gYGGqMeDt2ezNK6jFeU5g==
`protect END_PROTECTED
