`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GPlf1MxNpCkihpGY5uXmcVL1wwJjWJZGPSHapxZ1xN5pqTaevcAGmPcTOSm6p2OI
KCJUaFCHARVPf3dFmZdCLhSpbYxnvectuFwGraDU1kP4bbI2oiAtp/ALjEo1Xin+
5RWQWAegYpBOZs4Zam0HitqBgWTFwOtbfa5PrktBRE8R2bm1AQRkCDa2wFxEmqK1
j9759u5JVnYb5bumjYJYdtFyWp66Db+nlo+Z8qKzmErKy0DWGvxb5GwrmwSWDZab
lzdsp3ZRqyXFUq0owPk751UN/Q0fE0a7e2Ic7e43BUJt3aHEqyU2IMdNiDo1bkb+
Qzu740V9trRh2dZxsISJGC6n7HuaMOHG/lCxzvldc9YZ1f2L3zYRIanubQNpxMd+
ylZakm1H5og3L3FQBpGa5mxrCNO/R87VkGQxXmqITIl84+0KwujezaX9Ppb/72SK
1hazb0IyBus6WP4qSRa8W8EgYfaymZ2JwDvuRhWbiMnGhMgYeF1Ql45ihvvbE8xT
j9E1NdM8WXEWXSMXeXDSnmM3hNS9ZH7p2tQhmDpKk08vf/4r77SCjg2Dt1p2UZpV
`protect END_PROTECTED
