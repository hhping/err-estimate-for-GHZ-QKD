`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jTuM/VGYGKaaRBgfVGeeJWeJX+0LjeDwYUW5GTJDfjImvVIyZYAUn8wqwTj8rXn
wFQM7tIrs+vlrSCeVkkeSjepFOFeYBeBFT6wNzj2Y3V9EYwcWtUkspjCbJcuY2Mt
2rLmLlHP3yAg/T4rEqe0vTitCltlJ6GrU0Q+1Kru4koM+20UOxVj7sEX53lGC9WY
TFb2ON0bfkYW1kwZV9g/Dsd4Ph48OZ8veqRDPXwl/JjWawWXDQFc3pELd175yZlb
v1hiw+hLM0N439kjpmoqTeR+DRe7ydJs/p40xyhRVCg769EoWSgPjyl3xU1DhV+P
XdIgigqALtTzVvkeNEtl6qMxipPNI5Xw1uA65gcuIsLfn/SGXLGEWW7W4f2MYB2k
a1CA03ZLdAuE251sIfAcnhJzIp2djPNzTMm0+6mgsVPkszb6ele6JYE/eYN4jhqj
ZvIHWLsDsdRuHnxfMAaTNbMGAKl/+2oZObgLtN+R0RAXfudduP7E7gpclOBDvzxD
WRRPRWWDcvbPCh2aHPnNoaC2UyApX0VBXiQ7X1tW0DBYYFBISz830a/KcLYNpbLV
Dz2wFIK0M6dX/9AHnVyvAExNlvG4PUSToxz1XVp9cQnAp7HQNEKwXWni0OxRmk9N
LXprOUhM3IwrO4Hw/dN9UDvy3wHtqvlKhvHv8KWtAo49v4cWkUw8qpxw+AkLrhiF
f2mZc4UjHBCdYi/pqVvBxmEHABgGtxuybaf7U6zk32iVX/ndLzzZjdvkc4pE1pmh
Gbos9uyq8vjWwxw45tchT+1h76B1J/hI/H5sh8oRVotFTik8VzXvdH9ugob506Df
ZO7WUE6mwwNOzIMpxY9vKiEXl0EkIN4skXAYCTml6DaMvuKiocjzVDQ5JhQ0Ydnf
qHN6tpL3M4RNgoaZzhsvY6TdfYxEMdQapTzRfXmGPrcVGQCyoeIve+y4bW+aTAyv
HFwgo1lW184JNKuTi/rCWDUEhwSg6HrU2iu/iHpeRfKb7MUCJUdXDk3j6WgUxRXV
PF+ocL57TWeSgElEu0g1Z3mBzAfaa+SSvUBMFZpYDgRS7AcZB6ZoT5blnNYKLQYL
mqzZUYR9nzb6WlTCrAZKKB7chowtvE0+CpzK4Do6Dt94f2GuxMEHV2Q4o72B12Ze
dOpoVXfdlJQJQ2MZ1NX+tqFUNdV3JH/MAdwNCWsUdKMDYbkwVWd2tFKNFEgz7wmV
XdZ2WMB/UXxhOkz4ie2XkgGiqv5Gw3s3v2Q0M2D89cUI4GYD20HGeej9xzPR87ky
MNvkHGXk8jvImMn7sp8zV707ci6Lf297ZUQ6zxXWV6ESOl1DuHd0A9mPrUs1+rea
oPHhDzJ1tAzjG7OcsRVCIiClqQbgu/lZZPA7fFFyDSbpKXxCBGdezHcASNZ0tNv0
`protect END_PROTECTED
