`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcdpFq1wcSh4kjCgY7oHUIS2Sju8VWmrcx+9zshz+s1D+CJpc/86WZ2VqMtBD7Pl
0ln2djb7iZzRYXy8Lrw/INFG/dIlTWzABEiYBzw5+JfxEDTuoBSIxLUOwWWZjPam
QzEX356wDQkmPTmBE7wkPcTWjuWTSIrNBrxYj/G4S9thD3Fc1bF80cRNLUCB/TmJ
cRX7ORDia42R5tEnk2IkMKH6O9mOOHI31tr67rfiYY7tMZ2eQlakNZ7qgBBluE7w
DX8ulst8r7YQJfK39QBX95Pck/n6rhwCb9/w/3uE/IjIjaBdR62+3395Azy/C+Je
yLo8lPQix8WwbkqeEuQhpF/XyQdOcXdwXMdg4IGqLI6ImBOsJ/OZevEUq3N74HgY
IgVzv2jLAO/t61VHDJc/kotaoW9u391L+nUPBHTSP3OKddD6VLhPpy9pw680JiIa
oJ3N7yX1QZcgFb3Rm4nHREn9HX4RnwRWJMIfWeTsMbHyg9funfMdGab4+0/k6lVS
OYItn4ehuJW4UqISm+ma2lqJofcvTXWHwDt55hNh1irCjtDpk+HP75qcc6tjDBdl
NZeKFd5VN2+vaqBumf4b7CRjjp6YbWTNkIUXNQOl9h3Rdfp5nfbli46CaA6dyNa1
ar4mU+HVBowzPwdOTf7KVi64cUZ2EbQXmQj038geWnwCzCymqTbUJFa1bB+vB/1I
vbfjz9tA36Z+i5QIEt2gPgVc8dcPe3WNggkEdT/nEOhcmJlns9nXr0J3GT2JoKqf
cdiStl1mBdfqv1eo5+1s5ukXGdEwdWJKaHrzH9UYZ0lNR6CeKwtt/ru13TW64bAo
uyQ9iNMyEFSd/AZ5ztyjnsvBnqLykhU+nqI/mLL7JI4gUaxobeYoLllWUTZiMjTj
eAKg6moCwiZFBUi15VDRGSmkilZwXe+Vr25XjW4XHJB1Btf0N6AzfbUGCzKQzOog
RmmHO2ETi/F/JB4qLuT24Dm/Ipv0ahuea4T1sOWCoFS8iXv2D/NqNYLT96rehh05
IWIeRE/g/6JGxM3slhFJTqSrPqTLUzzoaJo7lHr58p6K2B8gehJFANJoylU/YnHj
JADHL9zaCV1lXvS04rV6Ymzn7WAVol2IAFhPeeIDJ/9pDoOCEZjTxQPrPG9QkxyJ
gzanCyG4JRPFOxpv1GqE2xNUmXEebxeQyrQ3rDRq6kXFh5wX1PU8kb9nAa7BXbnu
K9iVFpesvO4BTkUXHrVrzJPuWxjSdSkFgywO3dFWwRKtGng0xPiBheThEkbPCR0e
z/gLcPE9qYhpd5ESQxgmKsBYhT4Q1owk2pf9lSGlmyY7tE3j8ekEBcimelun0kW3
IGU4/9L/rOeI32KLH20F5HMJlSnXrPDnMhX8hBeeAAgSUub7SymuzTjhYLTZLVou
xBpk8UhkHyfXyEFBL0b6ZCiitC/mcW5QL7c1GIo+Youz5WPzFsZbLkM00QOWFMWC
i1AK5wd+7KXfvyLdOSJJ4ORLq5IdNXJ4M0xQyFkH7RBvuZ1JmODVNNZ6QoaQyfwl
y6h3Xpqa5yPQxtPmSaPpnbBREmaXeiHUxf6mU3zEE/15q5h2acHNZQkdJfspIcrX
/yLUI9hUV8rS3u5sp9Ww9iFdoJYYfpKrNpx08j+3mJ/Ed3iDKqGh01ohPFKM8xJG
IKZgD1k+B2CghD7RFyWFRDl6dU1UC1Am2EZroM8aQZACYiF6QXr/Qat880CwuUBF
IZF2xre02S9zfxcDlaj8ap0YQZqnlrOrfBn38TKZwOkx2UqiHzD+zw8FZ2SMeLbi
R8koeTMxFmJyaqaK+M5KfaFLEehdX2IBNAdcYclZW8+g38el6LhOBeja+5o3riEY
1A6PGqn5pQT3e02GN92p2EknqTYYXUOiJAYPgMM3wZ7Uc0/7EN396vsAje88FKoG
5qufTSnzVN8E1q3kVVM4XMr+kS9TG/LlKD8Mh40n06fEM0MIvh3fVyUKp4WsMeTi
/I8Ves66osh03baG74xwt1S4uX6xdFLW6UA1QmT5GXLaUOzE5p6ZAz6whplDSmCV
GAwgx029S9lG+IiboCkPxxalkt+HN1ZopBVDuVyqcUI5G8cHKB0Dd3kJx9LBCaXs
30y+QNdDKGgovmbKyDV4ILANN08z7umtl+Yk0k9E+8nDl/6Fc8t3vCe4AAHCCF41
i9aEiAgIMDwM3b0cW+Oq+vxAAMoqavI/Sjr35UhQ+dzTNtd8bOMZ4ENtkaBd4xCI
Jrir+6aHeFuNUf42JGwIujBEimLdSb7JNQdzdRuqm+/CMV6WNRF0sw7eXpeyVtD6
HMJUVRyDUau3bh+i9rFS8cgwuzggUTIVD0eY1qITBOkdPF7aWnz9QM/TBGf8c7Cl
V1hExn+Wz2IchNTGfH8eV3sbS6lK4r0wUHOce3Xc33f2QEqgJOcPDIDopWXN4tWX
qKBB7FwtMouxei2MuK8TGAzQl4LMo7c97Uyk+0m0eIsJHtFLZ8SCqfLyjxujGKGR
sSpADWjgjDpYiWynKRrhen4zSIQjIoZyYBusVOeFQ+SttmSIP0pO29R950O1MTo1
sd1bf28UMdgk606Mwv4R+FI6F0pW1lfkz3fCTEY6yO+lKY3DiDTtLiqIF6X6qTWk
YgsHzaA6+nwIw7QPP/PFMA/HrSHdqdv+EkKY8V48RnmMbEJQ0/Il+GFkz+2Dsfqo
XtPTc5Mkhmvdmkd+GL3l9le4c6lgdqHJzdnj3CiecxjK462kDOphK9N4py+8hP5Y
0WMvyJD2KEISoiLxuynq6MfMOxJQX8ACAT1a4cvzHmvKbZGj7A04WPJ5ipKBdISK
jVoT7imTdyhKF0ytJfDE+6Od5rkpfZlhhdhEXG8VZwnfiWpJyAKwxpZwVBa3ct86
ACu5b23ycvLxmmkQsHmZB5BW5IsO8pL4z2LyXtVUqhoeO3Rj7GiQXu7mrFXI96/y
5CUDU6aQ8Be4R8iQuzlHHzdmWhx0B3+tc0FCj5MPPMHV2BhLbwZnSe7MCnyzlbnB
1H2VO6ubDZ0rfFk2xdAkBPR6J3pfxnBnaEpX6hw4JT+iligk4aZBxutjin+TNIjX
BtTG5iyvYmWtBwDejOZlKXR76Eh2GMD1ERwzQtmyFZ6z1YPKR1M7MNjDmXFsVBoJ
1k4LVsWN3ardxw6pmPCg75yXPLNbeNKWNTTBqorTOnbcLFE2XbfIjS5TCXq0+mht
HnG4ew23rQ9PymvHF8/omMEhgCGxmkExkpVKXpCnJwjUyIgh+EOUFQFu7lwU2/kd
WXL+qzPOXp3JFLDagfYxmT5Fax+sB+3SYop5fmlQB9oTl7eAeXXT0QHfNEeJ8v+Q
s2Jw9PZ9XKUmfA28VHx2VhjYpRgRKBwoCS7KS/AJvgagvpbwNLdjxHqf0LhPWmXE
JBr4F2VBQDitMW/BvTGm/pn9XHNWHyIptxjaksKLFeXgonMYgdTeWPdz3NemUTcL
FbFFf+Qgu/PANDFvnA/G6DZTXi4OPsoaTb0HWEmiDZSLOQyl4TgZSQQND0nO+9sA
mAYTRimTLHyooK/Y3jWdO58ZSBtWZSJh52kSH994Wh9m5x+cS+6ZMhSj/zJr+QO2
OoqM5mQIJWXfSbEFkkbQzlBDAMluBkiB4SZdHA4kLptr4JrqY6wmPlxgqOTdT/j5
3aH1OUvICUAihVhKhQj8BdB6rICO2h/oKVeW7MEmqlCkCfGGQNfnFhFuuAg4V3KA
7NVrtQm5r5Oyvstgf30kNbPzKrJrQfapQ1M6AtDl+4GUNMCqQ8Q7jDtqVoBK+GDm
mzVS19bXB/hA3pQd7jIjzFe564XDgl1BHTRVReFBOw05qzWJLWDk3Mh8xvwmo9pb
VVuJGgKiEDzkx9BL4a9eweEHXtrLLrD/3WMSvJ73j58keTxcHebFQB5SDgfcCUd/
8nmMx4z4M0QjsR9DdjARPpMbzGRvSjF4OeK39SBGWwziW6VoBvkUPLy6yTEf2Rvh
q4bo1cMb+nKf8QE9dWRovjAL6A48Lp4ZSCn2Zni3OQsbMkiesies7k9ECuGn5Cjz
Nc20DN2TP3yD7MTL6gpOh/DgTECkHmxPYZPxqWdlq8mJM08iPkD75SXJVQInLyFm
ISwl5KcdsfmT25EGT8CzcpXxQOmwFZBOPo8RVD+Ey4QzYYNhphS0ckSB/Jv6Oyjm
B4xkz7LAtuzlGVGHwoyypf9ORgx2Tpmyv+cD/SvITATvu4FWjUdT14YGNGb+n4Jc
BHHMzl4j0zQuZwNJhhAG1mdIIXLdUHnRJvKQZD2b7/ovlmoR3HrpfkMz945Wx2io
mIoshbViOco/Q0zAS/AZTE86SfIGvYVsFjBi3CQ150ubUMdbEejZ1dc2bgbFNJXY
3nKK8w885Y6LusXl3znQoTrOT4EP6VKKowkpGQqQf5BGimi78PoGiWzvDkjdqLGc
BfCuX8Nl1L1bMij15VXua4d2jAHxRpZTZTBOuVKcFAxdY4LIA4Kp5g0hNcTq6j6w
P/JeJAQu31nNVtG1ul5iGk0QLjQelnQ3LnU/q8YoKqu8FO+kOOShyIE1TuDGgbu7
uOLvW8Y/aM9s7RwldBNW3ZJaW1kX5HBCienVnup8Nxy+Kjiuh8fMz+QUaPbOd54S
szm2XQtjMEA+YnH2/JgthrtnKx0/ZNpaYtnekniCgLz+K0bbT4wsDpwvUNVfNpWg
O2l5m7pxSaU1KrUKigKIJSqVr5UTA2bVaUNckDT3TcOhFq903lJSMt8Tqkjt4jtt
1Tkr7QqjW5c1z9DG3MjK6dZtPvx/3Ekyae5Wn/5xHFHhe9+2wI9C75o0JLo0V75F
W2kkLlM4mz9jaSGDxmgWn14I9q9B+Uz7xqW77c9AExxE7+8T991drSW1YanHpI6+
l7HbPLagAzkP91ezNdGrfV+liaXKI5YJL7ee+dxBWUAQJanHbpNeBlR7B2doiQ2P
L/I24TGhmaqHOk1nJVThUA==
`protect END_PROTECTED
