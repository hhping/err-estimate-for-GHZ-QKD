`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rQBHNIDo+9GOdao2Yzp+L82lyBKDxbHwtz3rkn115haBg754slgkVIHlAU/eHrDp
P2NAkLkTDTeWb/xxRyYvQmMkKUqG4joGGuTN90U5hTZfIPVz5ml8jNVd+/9tzY0S
0BH12QSXoMkvT/0DflnpcEAGY+fW05n0LzylsD32ge/rAHlVMAk5NDHoi+Ot8699
P21lfORy1AcJ6nt/DWYWPmnp9dqm+xNh4EcJPlLNC8uzmahs7YKTdgSWer2yiHwC
R9pyPVOpVyNlEk3IDMhNDc7VJ5UT2jyWjEt558v+/IZ9Qu57ebkRkRwBRfAWooTf
qNlJFTrzDXAKEKCDR9lqBB+KDbxCSUd5py2UTl4u9fX47D7X/YeFPKPTLtI1lfq7
/+3pIXbZsVnZ1c2B9848jujMPqPzqyo8ZTCzfdPFCe41J0glmedDOlZOK1vflC6l
JOvaivknpqBXsTOU8JuFywH+Xdaa3cvrt3fXhGUFmUkuAtaW3w0pFPJU+L0/9rEj
1G+fit9QRDh7LEmOp1Uy/g5idOrP8MvcASy6n9jN3d0cGosWFFNbwpcGclQjzGn8
+qJ/sKBgoFthIdqYUzuGwsFYUhyP21kJJEWFmIB1EoRMm/1bB+G40OZ4/2EBj2se
`protect END_PROTECTED
