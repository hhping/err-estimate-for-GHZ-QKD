`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+lLeWzxkXPDzEhAmMlekOTqcC3sRId0TTdU+PxzDcXGXTtrlv5AgTsJ+KLgvrj4
lO8CPxLUgXfdsYU+RQONga4PaqItZ+CC2vEcNuYUjlMXbo+F1GRQFJYBMJi/Gkn4
TpAdwprSOl79UpVJdWKo7DkUQ2GsL+slILhJGF8luvgZYaneeqi2xk69leWKostp
MEIVewGTmD1jmATM6/IX/1ytpL1BQ88W+F4kE7piMSu1+y15VjSoklrbCvbTSFo/
T/eyuGtfhf6DXoIV2l8jOjcUVpYKJFbU78wqzaQ+vdezVJ7cZNctGaFCw6JJ/bL9
QM/eWTdQgZ8DNOZJsJA9htdJOo1T0Ukl2TECML9UEyLKa5PSUyw46+U+keA70J+V
xA0lkYK2m9mMChF6nxTWp9Por6zmAx+Tj/yu/+nEvs+wSjTKobUSbEIN8+s0RZ8b
HQaNbUo5QhlBwBoXQ7dFflc3KqhJ/XCa0TfV1n5SbGhjLrzGRaPYtdy4TkSjo0tl
7/h7q8t6qzCbL4ooKyj9MRj1HUFsRiD1xmWw+fz9D/gdCeO21A2CkQzgEM0MWAd5
cif+ZQth/xGckvB1xkXnvhT3xa/vWloWhpG85gyRNl3SZUTrb2yiyGFzYglTLgJo
PWzHE9wsgdUNXD8fW2bkidOo9GEH5XpgcQL0rmwLZJGV+edevPlj/lnS92ZzgZu9
erJhlLcFybZWsewZLESZuFpB6y8i/bxMAcP9b1L4H0vxtbR079vdWZrPw/K4rGOA
45Hj9EEtl8/ttq5N2Oaiowhd0D2Arg/Nj5IpgZlhtrwiYku49F1ueS+iW6eFPkKY
FLV13USmomgrzOd5kk8dMPjL0joagEOOG+Yg7GD/z0YHT1Dd0Lp+0q4dZ7Lxtm+u
6TayZkBSmH/KjF9AoW+f9HhX2gdAz5Fsi2Id12iZSXXrowhi3O2WYRl7EODS8D1k
48vLmx8HlIe9wjE0cEAklDnSTMtCxr9vCr7kFasP1et4c/DaKQGl+xtdbA/vcwxb
BF7WLIACcJXMAn4+ZCLvGUi9q9b2xGQ94qx6wd8+wkv2tL4bQPPLOiBHocmXf2uD
IZCoPn9p/9l6hpGsE9yFA0d9DzdJe3FrD/ufCWvYM9+3MZY1+GHrY4+NskOJoxr/
Hm6JPy+rsqf7rYz7FTeu8sswseEqp0eMb8xhF+6Ws9fhW4Zn79sbo26eQFGU2JIf
sj9SK7IMAv8SAWhYAPcWfXqsMy69Y6lDZe+lx79eSxG2jPwOnuIC0hivbP8GwbWe
nPDwzdGlPacNMvuNvwd+mv2zHyxgV7fLOyM8OAu7H4tyOwCa4JfJt+DdhC7Ylm0y
st5aScxVEaxaJGpugpI7EXcPWY5hS2js/DX7+/0+DqazPQY4TYKXLAtHNqD96rTs
0eFiKQDRZ6gHXdsoEzQQs8Y0KpS3AxiR+UOzsgDTqz5UAeeKOF0z7UArM7GEPtet
yuSijpq9wK85cRpBfVlafq66ZoLriZNU02RM2WsUaKoA6nPhf1NpjCkMrmYTJusu
2JWXPu8H500AHYFv/Q9nGEDGjNlUipNpDdI7ulvP0Pva5suL5hK0zr71IAwJlwGn
NikhIwcNrEjWTLmOzBVN7SSczPCOb/Z7Mr+FYeMhQV5lGpomE/dP/OJiFU0H3vsL
wNC0SS0h8ZQfHGYE+oKmTVvCXsCxwWQi0yHTobr9iSQbQyL6srK0A1HW63gmE6aq
hNfKFmqrpQcGU1sj5ecwNwngsjRe4wyPFiLCVIkUW8aEBRplGI4bRI4W9mnuJYUd
YNVITRCALDUBTbJMvPuss9gu12z64pcq3whjey/QGYZXLtJTg9HqtEW/QRfTAypZ
U7zIAmYoGDWVdKXbblpyfebf5U6gEW6L5viL8LS5s4K2luxjvXIV++p69WwqZWSW
`protect END_PROTECTED
