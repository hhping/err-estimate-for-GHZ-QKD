`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ceNN01gyolMouSrlrzsHNaiF+LWelsYR74Jtthqd1KC2QESINqHOw70ACeDbkrKv
UYh0Et9LlJQr6bnIKlLckOnX9N7l1nIsuV+pnW+WETnvjArQl6M6yyIMnezi1AFW
6eV4qjB3AbuZMiNsbU+r7xBQN4/fqZxlBBNJl19bk78TeMj/WYdSdSkrZzhc4o5D
QVGf4ifXo2JnDAICzQKM/wdYLizs3BDXlV11ztc1RlzAkj8LIRRkFDmv1Llaq6ww
0rfFMB6CYX7wLutFvkJ620zdGrf2nQyie9iC6Xll+bc1+LN2WetwWq6zRebxs6jf
LKYaLWt2tx+1sjTvJeUUqp8DvGnq4a5gcWzQUDsfeo4ZNdOSIkYnSybeJOsqg0mb
HKyU/O+Bu8vwyR/sp0nb9QTUnaTx6gyDrKjE7SnvN9iB4QIDtfyN106FzZCvYjMH
Ye3NVKy0Y7m2YUWX2jufAGsvXs38IBqSX/8EBkvKO7XvQmnQPHuCO0j1RfJnrcDe
/f5HiHlOSH3R6ak/g54QlV2mN15YapKWgeGZDQK6qP4KYo1aqLvykNtIBBchtwza
Zill0Vu8bmURzUAlmvVr50AhVn6FpOoHPqu8QAuct1b5DP2KaVBWkhwLVxqXmGcA
+EW3sKd0n9837pE5MotaMe46gyZRbDgm06UAtukXENGAGWpveVcC3EsscQRSCNWk
dZBZ0abqutUfLSUchJ32uhcccLnQKHY/VJ7TPsunML8KJAulO66QaiGck9iFxujg
BHLuc8C8E6RNcYEXOSXmEgQfdcQ8m/b+gyZ1QD9X4o9OxxO/7SgO4MmQYM/YsIoA
KHbYnJdSVG999G39So37cBFo/yaEwK7p9A2BIb9RFeYnXjLxQEfuoZbsGrvgBXqY
yRSnogUeKFOYRWVeKMj/tFgtFV8w7pM3ne+IivWAAms4AY52jS7eeCkrhXjWpbWS
T1t4NjtvmRJ7yDg8UAUiZI1eTRgtQQ2l+9GIywk4Totj7Se0p1JI9nEJCfCnHunK
G5MGOlEQY9nULDcP/sZQl8RNdDP9BIcM+fRMoY9snyWGeNKJVfOAHgowt15Jcrve
lBdPfUUXVHoWeyDMA5I/3UqLvJuDoFvceGK/J4HHpcvQoeBkgWrxkd66DHOREBjB
VaX8BFSEqN8VDPqessjigHcLi9V67nUpIpvUIL27cDnj/PmYFG1JXXMlZH2EyN4y
p3f2hJPIY4UrZNlmVurjH1Tfd5Lj/OtxcBr33yn43BgimM0HBpClgVj9McVK2oKo
ogxlaI4GEgv4XzwVLDUgC07Sd8YQjHLXWVFAVFHZFjt+cooEMM4eJeRpfQzXQBoc
5v3SA9SyrQnaMsqIY4Lg8uKc5ZrlBuLwqkk23MODsc+JFK8yPqm4GTb8zRSRUu4l
ZJRgSN9N9ZAi7QClEb/Rj2AHDw7q73WlqhTa3wFk2WKD0+N4v0XJdnuABWyOq/yP
re5czM8wce3hakgEx0lGqRtd01Rx50l58BFpxcDUTaTPcFnGlxD2r1UYNQVACZwZ
G+N1QhPiSf5hEgY9yIXyq144znsfMKjG1WvxQBOmA1ZRqmTB3B4lS0sTaZrhjH8g
M80NEnUyweZNjvo1cl9Orp3HTCGIFrhgfXoeqJ51ke9ZQTjXHUSrFFiEhFDiEWyw
Tfxr0JmX83C0r9CM+t3QKlOptyVCwzcTrJGFOzc3tFR2GbL7D8NyKtOTif1/Qpyn
/0dTXwCJVl1fIcNV0c65qQL1ts30dyXrHVQbCujM9I4EmV87+GxpPRsZsAGjDGfY
w7A0voQIuB0zvmT7RxyUrOH0DI2VwOUEvKEfprsTWJy7dmq6m8tGgSBxAFBrD6ny
MAN52pKylNUDcjUhumtKb3y2jMPBoq38qvifKgP9EPPUtiXqq0E/Ec68krtWr8eS
iUmlddDzO//3UvxCn6PZybWfxH4+l1t3CtXX7Ijjg5+2zdES9rAiqCz+U9Y9DvDT
fG9LgPFIrE80fywgputfEREiy6hFzi4QccJEqmbIfuo7l4ye0TW0BC0gjtc4xKcT
LRDmz5DbcvNQd1HFjiBmM2GRPmyNkQiXR9NDkBUqQA0tlAEH8za0iKc7QA5SCHd5
rtC0VHjymg9X5q7/sdMhWLtA7tZ7wnRjmI+4sFvG2ya6WhjVEDW1TFaZzr8AAMfO
SkHtr/8oyHSAH2KUsblB2RCTdIC+euUMNoPcMOFTJtrdsKL4t73CtfDdx6d1q/zF
zHff2LEwhuGRMC0bJwNdqWln0d2uSOjJpZwyBxrC2Z+m3FK6WkTMjiD9SVsjBfxY
iXBt3XHTiofhRBXNqxcOF3+Ohx62zydFhvX9XGl0rMFc3H0Fx6BpaqiDK5QyQzT2
aCeU+GXbhg3UvXqdDsJk5uW30QLuVaDcMdkQ8C4tvkXFlomR5aCumSDVx1UDbI/o
WL2kKGX6TtMtrA/nYxb3Zi0c5sg7Q2mqjRajm5LHUVMDdus2zVKWZL9YxXgiwU6+
EDI+wc5ZkxdVivDgLXLEvs9kXLAFRB5k6MumT0d16K2cD+cGPkw6egwivCIWQyQy
lt3B7BUxLRVBRtLxVtV4LfXuNg7nulLv6AesYS94/m4a3BrNTb0iQFQx6tYuC5kh
Y/TqK+S2h70p1oOeBZBIcpWS6M8heWz2l+0ZFB9qNhPzmCQcrz5YPLgrupHknMDV
zBTydQeGBmOjSnJZAMFlB04DCWlMjFDs5tEux3nJ117kk5yTipPx4fc30mA9TmLg
UqUILXEOri//dGE1yuOckKkc9ppLNJejF8ssslCDVMs4RmIwSZP/WsYHeD/tK9Ah
NzfiQCVCHVCSttGs3bPqoN9+IdB3TKb5rkhM8d1x1RD0zg3VMmWQOlE67+ypcRu4
cTSBIEXi7s+2xeyjlUDcMIavfKNMraO8vuBs24VZd00RCJPMLLVMws3J5tbgw6ht
dpRWrGBgCBVZE/b0kR0PhfefrHISs3xzpWbRWP3d3JcY4jBiWkH/UZfsI3pVlEG4
jz0E9VPH0v9G3c+9fvNwiwfqcVAeW8/bqOomTFmnWSbYkwlsfm2TXjScyGufn8pc
DNu8dYm2xHoaOXrpc4I0YuhTSoQm5FP5ilU7c2ClSxvr3IFdzgSuDzcX2vz5fZsj
TxyFf/ocTgnivhw+tOt9W09sKRZbsEekkKIF64mpsOLGSCLjEHJtgJjAD10c8kDk
MDIno6CjP75sP7uU4+9hcYfsiuQA5wzubnDOtUFWVh9+DD+i2E0c7O9T/0tSYgtq
fCuOwqxdMaGhl6GIUPQviu30mV0AX+5NDsvO4fL4fhcnRJtVZHN9KwlY+43QYMhI
Moxq9lYoJU8rYl76CIRJAPGsWgTWJuDPODlGAa8ei+AbH1vTO35vTzt8at2rIOIP
Ctxy8+qdirfM+t/UAZvWrUsrK0GlStyQE+SV+Cg4HDvQpPXwaaxsH84b2uSLoquS
RraqdWiEuh8s1XHOZ/64Uo0wUa6SqsEbMeb2KfHQ20+pyXrJ4DAs6T3E/Cf/gorv
Yg9MMvSZIIcSf01h5bxAmZRyIRCy+EOIbNG8IuRLKvG883oRPUBL9KahtkarhQGP
YiycpmwYY6+GS84I2DhUNRZjapSiJV3eEdCsm9a24ppVpqySISdlrnIiwM3eCL6R
1mg5udsSHYp8Bb2XrAcVpowY1mQxyF/rvPQJMCdrZJdpVFCRNBU0YsIecwws0FeJ
`protect END_PROTECTED
