`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXEwYqCCLlUYTe3/5q3nywNN/8BNnA2A2IZFBMecoAhztKObQXmebgP0BTWXWUdE
uLxq3CjmSwAhHTApo7lbG5ePpfDeHEKyuzjzUul2w9DUj0hT2oOyZA3cI1kbZ1SA
7xrrUtEv+CpmOKeLVHGIzONeMtZ7aUOnK6CAr2RpnidugTOOL/JLcCi0nZjN2VDU
5rPE6DoOr4zG8+YTqWWlvcJiK2Oj6QPFO5XTZiO2lN83Dy2Q9poxoIzSg7EERPtN
FTM4X7TL9CFLWZoUQOQTZjA5ojI8Wfb2IC3CM2UzPRvGAYrgF7dRCrVtCiKUmy5L
K1axiun5FM/60jbTSMucgem/p3FgcuraRROzev0dH9OCjIuBkkZdsm541X1oA9xs
x6rsvtDfJh6IKAujE3V3xmKqLu90Yj3eNmFzhqtavAvWdrvD39YTy4HXt1IKR816
L5K/+2ox/3VdZaPQwQxfscE/Po1s0rKpTqFyOTMrB/9hC3To/gAUS2M1KtBQxOww
SFkDa3iRDvwS1A6Meg2j9n79J6fHdb08cXFnw6/vdCDrq8BhgiRiyDOzEo2af9jQ
0GyUWOE7cXTg8NcwJMpxyCpuioRBHSeKsMGF7IYr+k9/RbwXw2BRRzD9R9bq3d2P
Ex+/6xmlItcJXeA8wjaHlKpH1xTKaQwHleH+zbfvh4Q=
`protect END_PROTECTED
