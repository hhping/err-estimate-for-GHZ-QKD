`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XvSj34tq0J7W9+hEFBxetP+T+59y24tNf1IHZAXPuJqJCAV2C1rdIuxS6Qp95onr
ABPaLUwihlQ2rnVvSD4Pn0D5/wAqFbxvPlhUElWlpP4QJv+S51eMaGzwHQEkoiYC
3IQL1Jy2eGZs2Z8Z5D/dfQiT01umIVN9NsTn5oHDDhwy4sWVJ7yR/DDP9cwYWLIA
ohT436R+6fk44SYfBPi7pPQz7r7KMQwMN3CZsadxCeS6SkybflAdqd75mB/6T1ej
Wm+0Qtgf/nchTmYCWSWGaEWsEPnM/tdrbBLemHDxI5zZtojnHUGcVZW5HmBDIaHK
LvuVzsImgDbV4H0KfwjejPYn4ZQ+mwSkKDxdJJOoA38HCAQ9ttDECPWbTogRSnOh
X1t1sAUgYUiEBqaTC36aqrX6aQ84/vxx7RBKZyDsyLzi/iSsoKqTOcmSlG/SZVee
ER24uCpgzvQ7rha4+qOuu2C05JlgBzk13jMvCg34WISGNk37FfOWtTFSAhMIQrKg
FxWUeew3+dZBr8tmThRQ62qXMc6wAs1nfr77YPf7dsTcT5iSdvO3vOhKliaRQQit
nlsuVQgLLp+sHwaJ4gU9a/VqE0GvoU8EqR9WFFsuA/3D7uhaCfjs4OFU28UVqGWa
qJG+3AzfiX/DlyPeDCnwOpVz8xUymKq+h2ZYzZWibI80+iyjhNeS4oxTnzayFNkJ
9wjYZgIjfLYjp7XqjLQp+t+PEXIWXPy2k6X986qvavbJIHVd9UUaKrgoH33gXSbQ
wn1dMZp1T3dH0B0OFEHMQimHhCbwX5av7VLUy2jWVgsSpxtj7aHqoR+SV984Q9qU
oII0zBv24+pxNFCTfrfIQkjORg4dzNE0wQKNfBhX6kUeZSBfgS3bN05mof56R4Op
ShPha7lnSJt+i4Phpp0VuRYWS1frIJgLSXYELC3lqsH1KQJ+AW65oz39e88pVgLn
k9Lv9AxZYUvGe+dKDDkUBDoulImAX2iXGq56SfXtZgVguWRxq60q1ex12YeGtM1e
R8QHbu9RO+047ug8nFhqP95EUqRNhqmIXnqnQHDuj810EPR5jWYIOgs9BRGeoOWE
QlMQshf0LcjjAXXTrg2xrBsQ/zGROX1AQYejqvS2nL2FJfSLXPk0o74x2PoTxCOU
KRbzIp37XHJFJUIMzdR0/9Yb9fSp240iQK7C2H+0eBeDrWSCwmUxZhEHiCb2Tktw
czIg1jzEO2eSe8k+HWNZY3pVQ6f9XL0u1qZDfcpdAFTKMAEm4zNEI2w9d/QgRpYG
BB6QQaSnCNjrmz9IvGncgDJjA676hqn/rtuLn6dsOesVPCeuPIxhMBRU8IOUJevs
Yn2IocHlInNiJbMPw6W7PTzMl511R4DOpk2Y7jTFhZ3LW5fBzU9E5Tmgt8yJbNji
1pR+g5piwEm6z+qdW3V4USGLLN/frwC3nx3zn0HhQtg/XAuGtE73/DyYL97slPxB
OmRKr4/G9Dj65yWdTynpm1bY8BU3WiIAklFvafxiKxxPE08l9AphFURGR5N2tngW
PWhvQURr5VA5ysyyQFvTom6cfLTeRvd5XbwfrqmM/GK2BD+oAVofhqzwoNRebZiL
lGFnlN+N3u0Rr4VOFwfOgAvbsAWgcSmPzowZoTaDXyRANXRpm6CcZpSMxiyF9vmR
oKqHCEhevsZ+jCdi4L/oxOJ8yODi5ZEPnzanuduSuKp8kpR+VZTl89i/XrlxJXWo
ZT4EgjksAkdr05sLfxBHHs7HqqR1ZiNU5UVZaRBIoTULLQSePg9XEdc2VUQC5ZIe
zv9ujWAy+COD94TzidIZBOaZpAmf7t5nb/iRt9MxEgmZEM4o/LEuZrSXjxLkm5PY
MS/lYmlNojfGOC9bw8ID8avIiijdkZfy3IC96AvTnJm/STKQvsTxIG9K75Dp5cf0
uISSloKhGsxRLlKksJuniw3jvx8/NyzgIjEeShYIYoSJDyacX7xsfgEndEf0hxgs
ce/9JVWIF3sbJk3LQ2DFKiWt8poynFDViiuaa2Ud3ghOKzsmzQmqOP0RVG08iDwa
KNmxWxqA/cX3T3uaxneTpt4UtjOb7nvCKCPxsicJELQP0Ja1DXNxmx71j/lpYBlb
LWBZ2VnRV0PsDfVPmfg30oL4dJhcLLVj971/ksovtFoGkq1AjhJJLPw7C/xuPons
WrifpCWdUN0yjYL3w1cCZJX+5NwR0LAb66XoCTXV31eb7bcD4aaPhP5yzxm+f1l0
U+Y5Q9s5sm64JNu0MLWLSVjxOX0TmP1gTB7j8Eu1XftapLKsh9d2zsSgkH77WSeZ
MF9PU4IBcGBs2pkZanSdN1J15E3V8Q8RQvY309SY/O51FYFrTeZz5dxZrZfz4Qxa
SuZ3E2ufIOutmDnMHfEriBSczNFothQG915FzymnCshXEsRJnGQSNrdx6p385pWW
3D0XjiKT3uhMNCRcDyYMh/3ze8VVWxgv+lJngBW/BpARwty3tXeuLKiylSv7yXA+
nObO2pz8oUVG6B2EjQdwhLLX+PbHKW5XMDdD5gVgMgTTgVJnaWDp4eg0neEGBF9l
Re8HmSCOoaRUtZp4QjFQzl5m+PaY0fZb4XB6YZJfyHDDgjLPZRuKEyMznk97U0Sd
rCZLJL7474RvcBMCkSMCDswX0/XCk5YtEMG/lQeSR2ohQoD11gn2onkoeKr8xfHf
AdJSL4P3OBdUSTxD3EvMYiG2GtwZ60UMaPplMKC1/d7EcQYUBY5ps68wmgPvWtJN
Bn9naS4o6RWhiK+mzJ4gwNjNNqWwYiWhePEi5UL/XXEKcKOeCXOGYm9OF11EZag6
SANaeBRcewNApXu1LWk+2BaPKMlFDDdVn3ObQc+Xuk7hTZdAPG0YwP5cFmwPetVJ
ctLPZ8by28VSb+86o55+59uaxFp6jbatXWmL6RHG0mIVFwJwg0vRlD17O0P7o42+
R56bLIr8mpS5kud2ySx/m99WhswirMGB25GGvJYIYHAFrg2baAnzPqGVQwVXAjtv
M0F88vZv1BKkdnEzuV/lhPco9i+pKGH/x+GP26R4FK7JjoVhUcTiAPkntdZt/HrV
mQcfevM/WXbN6KpII7svd0aUE/tBF7oVnUCGkbIH2ar6ukIz+YQT2Tjnd8uEmGOL
fHbj1pf17Aq2R8Sicuy9BzR7A1NAm8P1VNffiOs+gv/33slBWF93SzFTOD4Lbyun
WQlaxtDW1Y/2IyBy0EzZoNCPMz6AuWD1A/8mGuz5SSx8/1MG4My8Nml7AxOcjLiE
hzbYfEIA+2RCTX6giHqQewt++FkODOVf4lWyKXnZEprPf8886UmDxGelbPK10Cag
8i0H6lRo2YQrraX5CKG9rEo3bPcO6qmCDMly0Uc6ZzhrEcNF/W5/NZRmcVqkVWyu
MPUf0VtLgO9UUGRyi/vmgMs4+4x/KAwO8xBsICIKKdrpH4C5cas44+UD/k9TcJV7
mNWmnM5rwaD+kF7AncynugEuUkGUYmPpGuuB2rvsOpNuX0PpaIbFFy807rGU9+80
xeAlVBqk8jo/WixBmxOy0B1GQnAkCEkSKm4CIvWex9+c2fQ+lU0qaYSJCeIOZVMW
kVxMiQ6uCo6eFl+IsQj+v0O96V5QC03nZCL7WpegbgxtZ8vjQn1CkqPGeExNVlWS
0/PY11bTq8RzfvzNSjImMYpBTZPDGApfN9+R9aqexL1mvzoQDErKeLP3PJ6fkrEm
0oGE95p973DsdrQpAY49yjE9X7zbGypFpt6dW8EmYqLHFvKb2qKa2MvryTXek7JD
twk3sLS8WcjzceEMZ3yCzMMie4yWCBalzSyrYWeu10ReaLD/PvAxy6+NAta0PmsD
zzhXtQAmvt+PXXCWXXSfkMANI59EN3jNlnHqIF5w7RQDFNlGembOx9U4HCWR+QCo
kHevfmB1YrIAhXbSxhhkoedEvNUNPUTJ0l9XuY72vCtXSLXsl+4uOcFdL7/V/0b6
fiJ7rITU6vM03JHPHOGoT5etOh2CRUTzX6tfhBDatbV246gMbDQiuFBE9s5D3y09
D9F3ZrrbfYO/3ndFdk3dFmkXa9r2vR6hd0JOQT2uy6Z1j5jlRBxGmU3cf4am5UvJ
xCfo/3kpZkitT9DcCBPIKAZKXdvtiBjJw9YzvIOjvbtzY4pcl6m5hOng6TqyL/68
/EQyJECiUphg942hTyt3EdDShQfJ/m6lJKnVv7tGs7RPr7HDDdzrYy8ej/ysHR0P
i1bVs5+2ZKsLr1lrJ5a/wVaZ0BquPbAscpJ1g5msXmW+PANeA/M2PtgUb5TAALoK
NoN3otmmrpGk9v/qIMCcd0p06lDQY4HQ+GWkwB4i5D28MZ8GOLC+DUxDcmTQn0TI
Gz0hcbUkV6q9DCAqnrX5PQJcvURyC1pyddvD4pTDEIROn2V2hBIV31Gtf/rjguEa
Cw+5azWV1fsDWm7u4KN5DFtFNYw3zcf9/fQEX++oFyN8Kydu8ehM4S34aeE7Mwg6
`protect END_PROTECTED
