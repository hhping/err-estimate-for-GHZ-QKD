`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrXtesTgsYZOpE0UzZd17xLlvq+TuN6UTLMil/k7DdYeFJJcswlCCo0FBvUnnYZB
JD1DlYds88RxGovMx2ZSW+cdNOTDkBS+vP+/z6WLVLz1iq+E2dek33HXvPOeWIOs
3DT9ZuK6kMX8gYyIwShrw94HJlEt51pD3Qlnc+mzcWMaKnhwuwVoKtQWQdEpILTg
f7Qr+gzbD5ztn6v+EVnMB7L5AuSoY1GjJZ+8F58ELYsCw1BAZEqDt/1+qtWZ8DWM
D0TPcxsjX7+z9BGcVodLYANYilwgF6XwhIvhWfPguUEbGAM9oHtlvfzvTfZWp4BH
BcPb144nkJgQJloLk3MQCs7o+P5IREDI3CLtspvpWuA2WFGlsMyYa7BknzyTZ9x2
cvzFXe1xvcdpp45q50YXcpXUrrVLimvx88JE7VCEvHlA1hvydKAfofS9Ue+Vqjfv
AwheTwHsLSHC8C1ro4DQZOH6kkE6DJb6zz1nKul7/CRsdr6sNufo32xcvEdwmsSp
jtfVemvPjAdmsKThIbidJRUBaD0pTh1eUchArN6BefD6vnt9ubpV5xW/zG6pXCg+
bZYmtWc/vrjoV7X56Lfwonh9JhUHwCkv1zrNLhlTpkFi8IH/z9AZoP9k7t67PQVM
XA/6WiCjm6asBYsC1oB/VBmexgRQ+kMo7FWXsxJF6FzTyaIqpZm75NU3kHgbrnIR
NkW13V6l8hp5LEMhELEePpIthT9MpzPDFvD7TnyrAK96hXI3bmsA6+ac+pwv81Ln
IFIw0ZB7WmcIqdw2k++biml5SXg8UhSOOFzwFqzkoSbLgDwQOFOGDjtCwTcuRp02
fKxJbkSjx/l6RIPGLQ4pxdhAdmVgmzQzk5C+/0YeBe/znDKPhZIlz1AT1zSotf3K
6WNwI3vNR/jPvdzIAD27Dq1UKoZhnUAJ1NlLSktDgQTs/UbFkDSszRGedMV4zKXR
K3esy7A8n8TaDmS5SP2bnigewvONbGJwjEsP409RDvWzBMGFXStWI8rZG0hulgNj
szlv1J0paJrbe30P8swoxBhuMGhBTMFm/vW5nlsoGD6Yh/5hICMx5uWBt7sGazqz
jl7z2DoQXIme7wgcBf5od36vjF2zecU5bOgw2XGHF8d55b0Yj0KZ4RddlXXu68Ux
31R+NiIQzdO6hTD96u5vXt/VXbmdusOrmSN1zK0eghGzx8WWzksqy3M1UM4rWxut
Lj+i2rlS9Gfa4dvte2G3pHkfPgf/dINaamCPAZCg49yJ+TeY+newYQub7aVADvwq
RzhgCnXB80wYzu7vJOowh/V427C0nJ0ef5Nsymk8rhgS7fWiqDziPQLQXVfhHwFH
gV1TeUaVinLCePwc8wt1DA==
`protect END_PROTECTED
