`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aao/o4q4ujNa2GwLgr27QzFrGzsAB9zOeAIAO2GpHsZU52CHfljMaJVqhkpHd35O
uTi5jm8xmJM9gQXhJPGy/W7+cLzwQKC8bebUAx0Zjstm5Fb78GsR8di6ZoWk9xR6
YGswA9n5WkkcVwSqQb857EqnYKVGatZn8YmWtw/a4/X0fu6Af8LXah//xgqEDEg6
ikICkadckZCRCF1ApakhSC/0FV5Dcf5f+TCNSlCzEHjZCnFlwBmuOIUv36ChZBdf
iV9N6FHRuqBn3zCiWeymKRzF8Sz+YtcyTEMWUmjNCOucDYrBDNw4BN3W2lYbDw/v
nFxSoDAAm7ycQnwsSRj6WHxoPfYgiNG488nzfbjNj6qit/qAwdAOpeH11i3+ZLAt
sfFBO+XZaA3TqBvPNxuvSfN98PfaDuyE2bYZju5wFuecI3HvLXuorIYSs/kLaJGX
PgEqmPoAKzl3wAUgXTk+dMFgA9H6/jhJeOX/WOGKM1pc8wPtcBhmkO4d6nKlemUI
la7r7KyLji/DMFc82uok78O41tYMHm01oxvNsrhjoGduwfEIUXOrJFc9cQFixz4R
tBoSfR8wwxpL3HwB1ArTFQZckqVz4PNn8p4Cy0HgPREHU3aNiS0AzDYR3QHWw4GQ
rb0oBK1Hn4lrOpPsdMW68CBts4AUPSJOI0Oe6/YjDnRkonR/pohnXoToDyoY+x8b
cHtIr/wTK1YYq9IN8VX8aRIetWRqNFEbvdZcxPvHYlAZgQ/ps1X9Vxcy6wtMXQdE
EdvH7WG2mmclI9lnkbuwGbkO89Lj1dtzuefRFeLkueN0mWFn8/JxN34H7rlOkVKi
8M3lryiHkndmcXRLxJnBgQLL37501TlVa8kZilvCLAJonBQRDJtVbEv9/5woUPSs
ycDTaGtVn5jn8tg8F37viEdxZY8gj3CJ7ulY2qRvITw6Dr43kGCuOKbN5lXGEWFC
0qPnyi6RGKaFEMG/fwh11/hvzh4v3yUviNVABNvmj9HZNcWePCKdyJakK6ltoKAo
1GrNlSF6OBMi1r7dkqGtlQ==
`protect END_PROTECTED
