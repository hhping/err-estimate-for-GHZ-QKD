`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0NJXv3DCpQhsZ/NXL6JIxsb8v7zRu04y7U0g38fPgaAzwKR+9gvyaICEYLSbmkLP
q5rhSJVKF9QVlY27P1uS0ysgLN29VYDzy0YmRH8a67VvNvQ+V3vT3wSB/N9EWTB5
3oNXMihr9BuurakGlLfTJuKjYEnBCDOJniO6qhTEVqD//TwKDHDpIiOs61ilKqS5
nXPFzpF/kE35QI3K+MjqDag2AVjBtk3ENPYO7lapKm8y6Syx19P/lB0q0agfW+Bu
9XSYqG2KNht+ixz9tCzLx9BIEzSB7PhvcJO39aIHo1nsbJ5jDG0DQCIhm9EA/o4k
F/3JNTUfA5kTNTI8TGXHcbtTuHhHuycCm0dwdrCDGL4yqe9GNzo9aUwGZ7iLoTg9
QbmBpBq7en8jbX+K8d7UE/DLXKu/cFI20ZVehxLEXaCXg+KF+7c7sfSHLDnt+tLL
tEFoX7tyJA1ZA3b8874WO1JnCWrHeGcfI4iyghZMvK1UH3tcaD/Ygf1g7up2UVvH
DhagniLIEyLXA9APDAbsL60joqAgyDgApWMyyEHc5J2j56nXussekisW/3KWcCJR
qzKs//CNE3dTg1vhMZ10loyac8owNGx+WYiMnJfEoHhHgRfBNh9K9djIBinPniU9
eMZQNJlF5sv6zFCBoH+X4xMF1ULFNYme+0QFnlMlquisgkQ9AerVHLICYIQ48hNc
4/aTn5xcp2yhJhtaaIQrH5iQ/Lt2/o2j+Hc4sC7JRr55SEKsfHCvEMxcv6OJDrLU
dojPRkRePcylnSeI5LyPoVYUu/WbuOOXgTlukOC84GL94Uto/alc+abW+Uh4NnLu
1fGAMFCkIvq/31zD6U0mfbtVpcOAiqF1jAhAVRgY6BIKZ0lMfGrw6PN8VtBLbkpJ
`protect END_PROTECTED
