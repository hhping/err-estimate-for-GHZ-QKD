`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MQzXth2DEfsJgSi7a7bIhKvh8kBlemtnC/aktwaUkH9/s5puzd50HpwstZKU6MVu
MPfv+24kSu8sOwFqQDA2rsBpq2airHgRRbie5XWCTDO+1vz8ykGf3FFVA3Gx9pBV
fbDWbrUAuCIuYWMPz/yX7ts5N2ZNVx736AO9iukiy82svKmaldzpvbR4ak3GEkHw
GuqW7rkFahfD2N4JhyWjGRRMC8zyYRfyrjRKuyP3ua6GHHpa9ixvGNcUvIX1H1CY
OGOvUoLgMxYOdb52y5pk3Go8eJYui0tEnS8HgpeoSJ7xhCv87N7MXsOgfctd+t2e
P+lqjK9BAPoLfBOlPowpQSxxaDHzHM1JC0xAt7+MyYt2n18HZA2mD/tDPQf0jFEp
yHwZQfwFhdVP0hnJ8knUOk9zSUhGMsB9OcFcNkbERhLYPCT9zs4GpAk9UwHSwRZ7
/eCq2iVWhySlMwG0g/461IpIjZOHiskSaGGROvJPnoCovMD6JDj7RfYBmH/nZ/GY
1U1imEuvyaRX/qu7EsQMr/9AzQUNa6OMyZVaE4h2xp/iHeFHxkNKHPzJNKHB5Sbb
Gd5ua3lHTLvb7teHQuJA45k64Zj/zG+4Vmm0ONRR4DTwjdBQ7WrMiRcUnkOWrM2c
DiH1zYXeMZFJR8eLjbP39jvM8k/fzqi1J0jRiVc+dj7k+f51h6pP+H//5axuc1R3
ZwOLBSmsj+bkNlj3KSZoSkNCV7u7w19YygFQb3FjCc8LzVgZihLglXP99VJAqdlX
6IJ6AZcPa3T/p+myuG/2x5I3U/udvbW9aEQ6QDcIqXvyAM4L01XjeKr0ZqwGYs5u
9U1hpBf3sDKrvl/AQg9z/+O23CfLyqjmrcwRHaGNvi/lR2lCFfyq+ElK+ZRmFdn7
NK1R9k6/lutUIZn5NTvfIQQJke7k1yHNSwEKJRpDELYg7ByAWUQRhUGNVW+I8Mex
HUzuUjIjpVOUMRkes6NroKaFZyNXQIyVcWB0lOAekq30otXat/7DwFyQhCFSO4n6
xtNnkVXRwVFt1cIpwL+XvO73LG6aclgb3WPM5aJlkkh68ZapMHrn28JbXrFpzBSL
MnWjy6c+vR9S1Nnr3Wjx0doAjO9gm//w+pJyanmgD3w2/hGhAoARWsXbykOXOrSX
e/2nR9CMrAhEPRrSSlj3xKetpch7I8f3GAO/Jby+e/ephdqa4CPouAvwR4vtwrV7
z151qz6Jn+wEGVowgKxLpWeqeNVg2beon4jiOOg4h9O/U/+/+jUP6FBqzGKWiRiL
swWfSYNcnhhPjpMwHGBQGuUK3l7Vo3oa2ynmdbJKcn9wAfpzGgBdy8tRBufaKiam
iuGNE2fH/d5dWQEPUvzsP/rNxVrikfNM9pTNcMBIsvy41mOWqlHQFpCAsPYs0aXZ
8eAPAi0LQbUK4ctHyqqAEELmUj86V1nZzJa/1nw9ULQ=
`protect END_PROTECTED
