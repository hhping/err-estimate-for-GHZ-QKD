`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1I4pDbOSFULhHFXu87TB/oz/pb1/Vj9ZZiD+a03vAXaWfWZ4rT/RkTcuqzEGn23H
T3JLwiosumJ4FFq3oAQHNf8NdpyAsmTk+RCsYbQ61+D1JV6c89KsyJpYpqwiJZDz
uCC5VKyZbp9pMUEJed53Ux1B35RBe9GQTP4Ul80oEhWHvkcASFJOPafr/yc2PVr/
3yueajVJwjr83xvxYJQwTCpaqBJN6m4yTU2Jw2WwSexTXrNSZgX2aO6m8sotDP4F
IJaoAlVhAqLzq5T4+0VXFSL6EMgR9/3B9R3+9IgyjJzxRNnZqaGOgl3Ve43OyZhX
1PwDuXtRgfW6qB9MKwZyfYz8o1b91/5goN5oTViDvcAV7/47cJM6JBL4ZQZEjvNv
Gg+Cl51lIajBiMvU8vao611fSoP+ii+86oCAtwpSbOn3ppXgqqPdIb2VvC05zR1b
ye1rRjy4KRhRjCBfFcjcdN2QnzLTVirl6N/nbwSyRaHphEYd6ML1Xv9ZLjneUSoM
2RIRKwhbzHONrNIdweZ9TPMAmnuDcDzsZvNKVUo+WHk3gAThXAEfDxBE1GSq3fdP
ozBZzsNcX9ZiC4Vlagv/fnhvNNQkqTRsEVa9PrAfTzdwzlO9f/P0UR4j50sLgFkJ
jvhRwbqkYu6leMvSG3FQk5+hdcKA8LVUHYdHXldM8pUXNzBxbsJ+l0p051d3WnQg
pMYPr9YF80+9zpE/SMoGJ2bwg2hMGUAAJsIxyYsRWVXfYzfallR+IVShbqVmtfg2
aedZQr8kiCZoauNsVoDdQVvBBLpHZvnswj1/CLvNLNmj01tQLUN856eFUbTuXpwv
a96PxXyg3hCkATvQ0iOhGQHpLEzqCp6ObCMsBm4uq8uqdE3mRQGc/gA6c3rUUoRZ
1vaLFrsnKV4Y8G3G5yUDgLJpPUtRvGh4KLff5vJEkDHlzn8a1N3c+wyDtpGQkCYD
`protect END_PROTECTED
