`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUvJpjI8ve+yPsrE73CeNYd9yDd/F3amo4ctQ1zQhEyCJbtDdjzo5kVxB3JtHMrB
BuA5+zr55hM3ve6WgMq3KN0TZlT+jh0A70dtXLf5BQ/J4/QDMa3qJPrb/3NHr5JW
vXzmDvk8FqrEfKIfMC7VDfGVyoC05G2PKhrcTeqd/hfHKoQ9dPstjr/2Ae8IcAGN
FpkEETb7Sm8riEchChlKxfq72Zia+8J1uSx/Z+LNop3ggVa+CIwybew8/1PpW6vE
M8OInmCyI5lJrbWAWdxN063xg9AbVsSnEiWy1bBEsfc7vesONB4n6ON08+OP8l1j
g96f7CEKi6RHrhn25foM+n5msjWaOW9Ml5Fdd7WHj2dKudFqPeo6qhQvYSZGpyoq
fg3YG/RTUE4rO6kLmYHLlkZ3+pCrFlv10Y1mGpv5f3OA9vQ5mL0JEQs3tEMKyoZH
gIgtTWFKqX98/X16TspWHjbn8wvRFpEatZAzTVkSaLUKNU7HZAsdgPVNOsxvYuS2
wlu8JsgQewic8FkvomymG+ZUnTyj133XxKdmCbUwsu+tSfSnGXY9xJW6Wl+VjedN
tNhuBFcmrHx4jgNjxKiBZCt2E1+oK3+uZZQTIvbLdXYzaIdCGPaWopBBj9gU4nEO
KlB82m4wsqmtF/m7pNasnSxff4gU8MMLPwBU9FWzHw96TkoKHItyY8AmZ7Cg29Yd
LFn0nMbyYlssR0Uk69fjXImJqRqXozkH7v1Ag2nA3ucfkYW5waXNmL50OCa4N5Ix
QL3/0exn48czcLKBw1QJ6rzgQZHdJa1w2btvxI8sGD8w6tbztzRQx5tbKmZKBtcw
9liWAW6WJc/eWwByF8WaUBQ6rYoF2VGOUd8rOk2tpebsWadkhphpElUGQFJ8nywN
lJ8aPvquXNyOGbgMJWyVXVDKWluytMKJx+2DooomK6nWU+5Zw+qijKJOudZSFJQd
x5o48oVmLzxOxRwMfw5aBmGmgVUo06n20Ncqz39DyteLOKu93MSMpALNv9Ukg+a4
G2t4jK97ymuVSX2jKU6eCsQIG7nu38wPciH4NaD4aYRWKHIRelQOf/fxSE0eJRAQ
Xw/gw+Ddc2LLWLs03yqfIVgRYxCgjpxvKRkXTa9aBJ2ogVwY79LTPHhwOvGxfaOQ
pQ4kue2tO4QW+6S/uwptBPoKi1Nld08TrckT2xI1r0+bMRDR4H3AFHR+ZkJABOBm
sLaEIzBVNefhpfjhHB0Z8x0lZnyZnmtNKqN0/w/RgKeBWDBmTTKipShlzPTJRARd
YRolMJgigCL0AL/mYETTWVxV0H+yUzo9g8QaDO0AMCE=
`protect END_PROTECTED
