`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgJLpFpugOQXjYcsWiLwBDil8lK2GF0hfCMnf9S0J98MVSMhROcUmVbAY27B6TAT
Fj6QrBrEXQBkgf3htwpHPuIU+Gq4PPPYkexvas0+vZ0B/ZFSuM4QDshnjdtxAxUw
lmHoSE9OxDSIoqiQEEyVuUQb3qj0aANG1UfYuLcWfi3TSxTdT46lVEkAga/NjZD8
npSwDgke3Y+bHyC3skE3zZ8nePJPJ/LE+zD5YzjBL8clpaJFW5AuoXvivFGbzJYx
Mq11QSHJ1PtnCYbe3xjl7KRX4eMGXQFsaAnc5IAHyLk+LKtoM4FBq8/8pwXASjpT
cWAQFRyI+mo8jZXdHgRBrodLN+TToU6jNDv9Lp6oDFNq4rbYCPU4NM7QF3fwgKeb
6yAF49wPDhc8q2OhVGrq06sAyUgr68UIlCO29/xyBSPExqK+m7iyz7WfHViQ21It
DSADbPfaQ+FeXUl8eEB/AkvhqrCe0Z5IfaamoRFAV1v2MhfsDJg7f/AbQqVvYGxL
K/LpmeZ5tATnStUUsfrHc2pFfNq3c0vVDyEdUUo+WJXfFk6so3k3r0N54IJ3SLLG
9dIQXuytBPdpYxDmdYn6pgeoZyDNKcxtgi3Cg6vS7s4aGHst34xXtIopwOJ5zYIY
IyhjBb6NGG5QuH42Y6MCjcutuD8JelFyxvJ92C2pcg+iWPNB7BwzhtSfpZg++R8R
OgLml5PH2oh6VHzkXeaRyf7it8+tWWvJekxOqER88vMI87l/TI13dj2rqEUmAysP
PBOLlZAi8LeXdRSMQE8PhuG+GAho5nqrejtb7Iixec7O1QfaTKTm+j61xKntqL6w
KZc/QyGH3sbHy/pLSUZo3SC7ZJ4iHA/UVR816XqH7yzj7XFL4AfPWNlGsYiOrkyy
COBjCzg0YGNLoA9w4DV8K4FNDYMcgL/6BL8nFDvbVKqCINTTWWeBHWSC5Zx8M0r1
C8fKdVkiQXI0+dqwZLvmuk9B7BZgzXChkTS42bs0lpI=
`protect END_PROTECTED
