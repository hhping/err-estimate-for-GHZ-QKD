`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WbDrLJwF5f7Vx6aCUkpodVrGkmiEHKqce77EosE8j+E2AMO9SKcvR5EJIsv+Gtn3
IXo80eGwxJYdBMenMxv5BznEHpeku6THzCUuTJRXCw0EG9Wd3DHvGlfymBTP3nv0
NZKp2fQv5Mz57owdXV8/mmUlYXdtqvEo5U4VjVSb3yJgc7HaBP+K3fHiCO4ji3zC
VuI8k5calbpcrZ7VA1OJMN4qPPOSDezJwca7/UHoINSuVmo2Vzfrd1F8DvoIASwu
3RXq5gz+pBY3bYEhzFSGuRy/RkkryYcIPE7gWQdZkAgKved/vTZoRfpSogN7bXPR
Hxoe9MPp+1hka8h16by9zmehbxqhPKyIw0+MibkKv33043Cr5SvhNIuNUU9VHgKI
Aclrvr7bnIIjVZLWBs9TGgZMsn6ZBbLnXG/pzUaNSiku+URjLWuGste05HcOJ/KQ
vefVrdgBdsuCe+8IupnvxDnZik991VgXJ1QIYVPgwUCb6p49TyCHukGY4BGGUBe3
3KkxLN3luXh7VkvSlRrUN7A3XuGBUOCx/M7NDBddRpwH786WOTxR2wzlfCBJGZJK
qrZlplDnicG59tt3U+R4Di96knJMic1Bt6hvdEA5+DaraX7SoquX5V9yaGvCTkmr
c5mJwFwKs5Np1pw0UkG/6PgX8OhtUP2wdydhvd5qzA+0buaB7PONnKahxe8sduNH
sRbXfCLmnPIwV7S2VhkV1SPQ8HA+w2a946pZhjjN169K7bbIjhnOUtIx2BZmgdu8
v0W+G8nCDrYbQeF8DR9MJqgsd+aFeaGhizcXF4MCg5+20ZTWorS2toebnPiZd00s
N7ojB+q9aKh/JXoKEy5ZtsqREvn39xArvqsUXv7eKaGi7ob2tOiUNy+sWGTr+Ly3
MwCZ2ouqN4JfLpQSWnBYd1BZU3D5IV+c5ZqywETC4pExcV6qV04jc5Q8Up09cu6G
6OgL0snIdSLur9ASs67QDXtLOwqS+VsvpFDLNsLpfVo8aPXBJlv7tA+MHk578UyS
ju9tdgSw5c5ACkyOQGDNUvnoE9c3uBniC7SLQq7TIL42QkMvxWnfl6amM2TERWuj
R2R8AU3GXpTUkS82wOGTlDpvSntZ9B5FM7B5CggiPSHybg3yLA7wRdJ3RCFVswKx
jYxLHpKkRvL11XcCo9fsomzekHP2xHPNamEUsveD7rSUWoDEsndrwTBMF96vwk1J
Vti8SOjz2w2mqFEHg16cekH4nVZnzqiG1rfqTuey4gKzUGeK4+dxP1aOIXLLCuU3
/502H2dkrpCdV7mWBOCF66z73xEWBPxyhjbHGZ9xMvx76LZSClFUHFxSvzsAu4IN
shCr1JKPVUjCxOwJuTxP6XxEwTTY+ZYLVQC+QeTpB8nD9rbsdxgojddbNUnbAINL
OyTt8entuPDRHtp4a21IGQ9JGUxIHGx6qQmwK48t03wLAu9USdyRpNMG8lQv1yVo
4Wk/UG/zeo6VWpKD6Ji0/9jWXO85RyIiHwXZ/RhV/uNyGVUOsH2ayTI0d0RidqJI
g5ueI1kLjPaLivES5juBZpMZaqiOdKHmAJysLoG991MJQ3BoV+MX/HsXRkte7EOj
Pmf/0Yytb5Y4NmVTyKSMoxi5t+XNX/g94v9grwj0jgAbPbD53/5008Wj0OKmzAGF
m2VSt67lg3k70/r/uS1uFDZaPG49f2fhqO8EMDEulu4eC+tgOVkGWyI5VldNpZFK
aaIZyAhnhjElOyf3yAo9aHxBBts3w3S8xiR51FMSSOCWqWqUPezXH3h5bBSt/dIJ
OjetPepmWzSj+0sINHy/82KmkNJ2ueXfIcN+hQ/9fg7yOYVPEv4bXAYUz9dX7/wo
yoA704moEJkI0jrJtwiWMj5yNBKcQOaDNtgmSGFjUtv86L0cf7QjNcRb+xJsbbCl
EFsOY4aqcL54IRoRkiYLqQ/i6/7Yo2EPWHOwGJq4ac5EbfR49oYnGKkBjtht0O2z
+naYR+8IHcwmfnlIJms5aVabfTNh0wDn2IY/BA5ZSavzxoG9Hp4rGO2ldMWzWW/5
qS0kn+Ve8cRg1+PE49gayl5DdhkeDNIsUWwEm6sC+Zm2QMSKc28f8WrRP+NdkF7x
kVZUJnLoXbkCzPA3ba/hZRRPVtJ1PCqgvMQ+rZbUqUdlUGtNVr4lExsGeVHthaPR
OC+stRsCeKTwkAMvcOYL8NuLT3iDOWXzyCNL48YUGc9WC08GWTmd3briqMZvB7uy
Ac1owLKqstK6lJFA90N6qEnniroPA5VUE2rkMRhrGEGnFfuA36OnzWoT9hgJxOno
J/BpXLUw0mz8h7NUYGDhHSdMzR7fwZFLCIjay5DKHtC46FlVnLCxNb1zxihfDOIF
hfGn7OzTjySO80+GXF4+4oeHAztXU0STGOVFXRcoCHq7gm5LEGfVk38tNYElGLRl
CkPRvPrY0E6lZFbK2mI2M+iwVhsBw7pf+iGt/9pQMD6Pkx2GuOsitBXEiNNU9v9i
nbfTgj0TZQRkuEhb3V1M2RsPVXk3nwd4C8CacNN3ncNHwy2Map6CzeWYDZ+ugGg5
UZiZl8vEon4TGQu2LNnnXuoxrqp7RnutfexHlhdQxALocmB+pQquDckZwA+IL6Ui
TCc3L2nqsc2ulU4NkJcdt8CYuU98ieUZDs6yDYBnkYi5EYaCU8r2NxXckofL2Oft
tYQJuV80iz7q1AvwPfY0bKyr6B10FnBr+c0+NSAWjS7DF+/Khcg2zQvrPfNcrOts
KBi6pBRHDJE4qAx+TRa6N0q/YLhkV/j2MV/jtO5sHLWwcFYvWma3kaXTpqNIGsUM
DgLQSKXpl6UTTP8hjYWjbz4Jg38wnxEyQzdPD6xzgz7TT0D8+FV+LCLnTkaQo8iZ
2sc18UcIBLWquJ/41CiC6oXTz9hgig6zAuy9okULrTHY/H/ep7PVjXMZ1eOJCUHv
KRyXFnM1XeWvvEhC6/r5I6osLKCywT0z2tt87kba2sFQb0m85MxYwGMVdadTETSc
ep0hMBFVSy6YeEp7R+k/6OPoJibaArDSoKxs71967kUow+5WRHKZ6Lmw7cRLOUfd
+6jNbP+adMHN26c1m8UzRDhohX/Cv9lxrU9k/3BdkKmQFCH5MsruZtmSHL194D22
mHdCGL6tC1Icv8bhI3SiEe7ikYlz/kOaerzWDIN9vijrUedC5HiVAE0nbu6yHz0Y
Q4ywatruftqQaTp2LkDNWNr61nNgCL6OFlNnMT9sBsNc34Ks1O1SgvGQLfSVLRII
XTKm0a9CzhiOk3CheNuvOgcVeNNGaO3Mw6RBPLqxaa2SmAiFqf3XOYsKSzFEY81I
/4V7swGuygiLlAa0zQDfjVH9b4VGggFF0n6gWaIdPBiPQdJLMnsfQNHsWLSRZOLF
lBSakXMa+9pUbprSu6fBGcaHNSWVFgLlW0sYCibpcuYgn1j3Cf6oL8dqwniattJE
YodJSjB1D1TCbH0WMoLfHMXUk3zEBD0cPJF3emBH8og91l+wr/A0LGK7qVyaQLku
itj5m4YhHq6NrLJU0NDtoxqPmPhT6CEaqkuaVaWM3RUp3Hwb9cL44df2ATssIbM0
BLbAwj2EGK745sUDndZqhRtBXR/MsOsC0vFPT2lwAntadbpy+79QJBWSqGa4PEMl
Dpb50ioN6LMKsaHkEPcc61bvN2UXozL6X9S2gTduDCkqjogYx4RWx1L0MNqrNI7d
rjsw7OX10hzzy4Lm1LM30Q==
`protect END_PROTECTED
