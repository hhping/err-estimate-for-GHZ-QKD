`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSw+0l7RBr7Oc+6EV/AnY3qFrIUWcJi1FzhksqbA0LyUsqnfSAf3djvUgEdhU9vB
WGrWNM194mHoGVqUbrhxOOJ2VMjzZGh1zTorrdyzHXnoCe84rzp2mtWM20ku+QWO
K+XwU/LjzE0YogYN3U193pytIxTlCuhDQCQ4kpsG5eAx9Lu7Ma4JyTWfA9g5fR5G
8QlkLuTehAmUTxhomfYAD0qbkzNrtwVE8pLqw5NYIbQOKUbK9xNJDIbofg2b5eTh
FpxIU4+xRunRsjs0jZ62GYdi27OCPvm68zYS1s8jYALfC0JpY436Z2zRzBFp5t0I
DyarnL6SaO4Yur4abmTlbxa+oh8t76DDCZOVZQ+QPR9mqzArWtzBfEWcV9PNkfEx
LuBQ1apAuvcRFDbulzop94UhLgkMSJglecIiRe7vj301gBaENS62Srqs8vt3fnvG
fl77I9uRpXVwwEU45hw+4Mqj9yIa6UOqNdiq1xOHVdG/MKYbu1D4Sb7Xe8k/wAIi
s2baSDLySgo1UpCHVdM739RUl1UZZLmvcdtrriOGyE3wMjRaxMBZOC7symb9dq94
qOaS02aqYdcfte8UeFEGAfPieRhBhtp4bl+CAIkAuE1jbfPDZXK1s/mC4AY+JpHx
JY8lqn+3yqSfyG2usITtv6tLqdTlxbCGA8jJd5VlGz7Nq0j46IQz54uxKG+Nod5v
+w25eFJMVGkCdRiPWxT7KnOATNX8EdGSI3HH2KeufmSkdM5q3QTMlICHhc+cOAFK
nyVAsbgqXHuHcmfmLEdiMT0pYUe/XXbhekXxcXs40HDq6Ae5Ut7u5DxHoeg2SETS
oZdBm5EkGfkjnC+XDYWq4A==
`protect END_PROTECTED
