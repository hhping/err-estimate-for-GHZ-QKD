`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RzD1Av6ARgX8ULc9v4wxWnw8ImCC49zJ7J5308rWqq0w0Fcz+IMSguENYqyI19Zd
gz65eJXCB4Op4IG/aSg2Jjp5cMtvWIu5bs7acOjHMNZevznDrj446QEm7B3/V1Bt
RrDKwEJRO0W+HxiszWJeBATNa8qvNODFbOLlcautP4BmCQWuZclUOxfKbh2ux4zR
S6qgCxkxDP+WNHN4iBI0v71dnkHf/BfbU2ds59iz05GgFtQJWfpBi68uLjLrlll4
Kh4r8zRhs8gjc+sEZ/EfhtFy/AIPR4lYW1OLAe1AhWFKmiVBgWh8G0hO60NSSFbb
keZ9peYvyc1zgmMpt6Pyd/Nq50J654+Ho5Jii/WMa/6QtMElJ4hPMiH4TgNegxTd
zf2fC7j7nKIkoW4O9ZY6JnAqnOahM5RMMzKE3plfOH+kDRl5HPBuyAuid2m+Czkg
2Tv7V7UgLPso0XR7ztvRds6O0tJyQeafYvHTf0hzDDpZJrtI7MwG7UCmrqTj7Gjw
Z8XzAswHGgq/sNU+bpOU0SOBphHlSXjqiJC1izkZSYirqlt8QXZvxAaiH6O1j0fR
lcqNQvU7aO6ilwQiMHLQcFIYGxQLd0C1OEXp4gZdpgkcW5TGlXXfekMsHFElD9r2
Z6vWprfoeeT/x8UqLPolCDYbfKHc6srbA4AFEKQV4PSLBtPllayF61dh7zblurj8
P2SQHGC3P3lsn3ljvZX6ePAd8NxFqxy888NpfKpxyolerI4LA7BeEYjgh91JEy5v
UDXYgiSTWTDqSNhdjJp3z3JGowoV7dKy9sZtTj4It1m3wFeWjB2nsCJFMPQufXzI
w8Zgaxlddu/yAO7WgGJuBS5MZWei2yL3qZD5Wf888hUITMcTS+UM+a0qfAdvxnA3
5G2zdO3FM0bJi7wKHLGH7k+POKoZDbgM9n+WGTOXv5CgAb9J6DGxhRi9na5zmiaZ
TQ6wWmfSCZWNyMow/JsR3FQu91wq2xzgpFD2UhnjtfQz+ZEZAA6QLn5+mO8itOpE
OsF/CAYjs+KjxI/W3S76CLFSH3MZzieWGF94jJw22oxloTEEZ9u+eGvdB1/JOp7e
McWQW8fLeYBF3uJimhoy1MiRBDWXRRq8z13TmAlfgsknFrhZKUxxISuArY5WBLQz
3yFYCsHtKOnUMkgPtoL+opTt4/j2WhzwbEtBLgGfSIPFti2lwO4yZfEymlVQ4euE
XFH8YTsW7CCzNX5zsB4Je/a6dh6N8OXt9FwpvxmZ7M5A8jsI9aEVOWbb90aR8HQX
2ND4joen5ZEoEUpt4vCA2p5rWPkYlxWr2EE39b2d95cN2yFsughMdpK5cuReeIDH
reLjT5AIhUxhpPdYJW92bVpiDvGfVdwsgsjxKLOu6YcOyOOZet0w2aw4xRAfac3h
5J95MTWa/QfBJYVNbAKIsBoiz0yc28MHGkGyttU8K+MsQ8B+Dp8h8YURCo7+LCtS
dhpF+Q5J6k1RX5nYcLor3V9o3VW1BR8a9fCmm8OkD06u+6YLTBxOhFe3Idprk0d8
99S9rEc7/U65zRcKeHKS5A/GUtsiw+TBBoE741DCNX60evsIBKQxaams2dMs7+th
WDG1Y8hUoMTQ8ljQ/1ZcNiaV3xVBKudbcklYQaNTba/Ktowr9FcAB7zTaBvx7Yuc
55Fj0YsU4KAj5rcQHVUmqIgYTQot1vN9yoIykffMnqvjcB5b/OU1cjbM03Dh/bt4
X3iRx3GUFsxtCk+hA4eKwN0tRXi+Dm8R51Su4Y1xTLOA4kPU+tW6bKw1TXYMn+1T
sJXc6dmGXE30nxFjuAc9SyEhXQzhffxZ5YIh76dTPXxTvpQuQcaRN8btJ1+hhdqx
HaQbvDhTpbe+UbUiv4RQVzgK2oiNOJVpbq41I2IgkDBEOi6ckZaIwO7bJjyHATBL
OgKozCGv3IzdQX+bC9FEFYGBF/WAj13G+a0UWjPaKW3mrIDDizfSR9gnc2Zmv+1J
wbCD4NBoA0TRRd8mFvzoiO8Vlkkfm0/Qj2QfuaoZcuTMSVq7Mwv/ujkUkHvUQpv9
rbZUrJl2O7fS5FvLyPfCkniopoV/ry6goqreeThKM95S4qlcTLsRuLcxXWJH4Qda
a2a5cj90+VxLZ8DX+OTZdt97ruzmo0P+ZAdB06JvEBnsjl3xJKaWHjZlYeFyLHHs
U2S9im3WDkXmhXG6feuWVQP14/ODrJfvATuJYE+S1g1yxSIAPRNNgkjHub9hfP/Z
G3mufyhZLtWvq6JRfhxxU2q5erw22byNbhJ+vDiYsTQaAfhN2PECxl93P6I0kT65
Aht+nWUahEkTj3GSPOMzgrMD14hqa3E/7/GAae6qfItW/jlQrlB+j5WD+cQlFbZY
8e6QDR0WPfjEUwPPAg+esuMlWmCntPQPRHHCB2vh3a9bERg9XNo1ycSHA3ShpF4B
WLwLPZfmzDf1R92hpTIsuwM11uF6EKUTvpOZEozmtzEWG6r6Fy3v+8q0psix5aKp
wTO7kapBMGSnOjXSIsKuDmkeaAMV9uKccL7huNL6srV6nM3DXbThz+7dudzCCzSm
xhxSaBLEHiHWwWn4dEZcWsEW10DVbAMZ2O31t2DAo6iZjeE9w1zRsKVjXe9y/I1Z
N2eQjMBZcHehRUl0QliyxulfPVqO/SEFF2K4IvNfN6jWujXVdFaznw9Ji2qlw6or
oOt52BPch7F7i9Hn5nQ45au3OMriAPz7fnebQunvxvfrsFelLgxRrqjkh5dbl7bT
z2PxQC+AT/C7cnEr0e7/YcDhXixPkaUgxV7UBRk7pKqnqZNHghJiijFGaKEG0Ucz
Ys07p5wEQg6/FEuMD4i4Wl4LClJOcUCXT6fYvR0LWIVlTAtRkYgYSb/rrqwZkaT+
J5L+Uc02JTrQAA16sk09RNJsb7d7aB36jBnfw8Qs7R6dqWzFXRoJKYbGQCYa8yl7
cHxs+pyrI1wTZPis1mPuTSuyEUQ99v7JAFes31+pVEnfHliYNFi29tCcv6OgExuw
ptXzX1EIKyqLX3MTNZsNSsadk3tmNlRd+0RLoxBn6h9FqD63ppMWjyVVI6bglz3u
6R5V2yIc1KDj+twxrebfxzOT4XvsQc/cLyvIpfmzqgQUuAdP7qTluuAb1/ZedaKj
18M3BGZXrSa6Ld06xYyFt1XgK00RUrC2lvNsVk4tvTB/gKe94o2HO8y33Xod3lPh
cgUxcfTVTUZFQyPe+ElUQZr5cMKX2u1DkTJyrEK3cOKrW62+qHdPIaIQQMIrYm5H
vr0qC8oEbXNWlSTTSGdeuTO5mjkWvoLjO196WYlrCdKBmU970zxk+iXM2hMy8JlF
ylzMeiXT9CmMCppU5LVMSGX5pbUwCRy5lsp9IXOu+o5U7iQzdGIfJAcRSzkXfZET
jvXThrsAbDXL1KEDz3xXMAXvLznMnB/xUox9P0znIoJTH0DV2xSM2BKYhd0QesDT
8kbYK/OiQXM+7Eb0YtMzyflVcC4q08bzDgnZy3LRkCyCrCXj4sgkHt3YHiR5Itda
gzNHIspkNSseLbbHbJ+I4LkqbyRJxLypqK7Rhe8eM6Gg6M57U/zYKG619o2y+xVE
4icUNWkfvkQ6t3UZXADIHQ6Js+Y8x8YPTNPeOBxDNXio+Cbf/0//rL0Ir/mF0QGM
ju5tG4p7lLr5hUb5/sm0Cr9VrzLbP6Sl7XcqrW9/5ax+6cUGV9cfv8gxP9GyWvnw
Pv+6Tpg0YherO5p29ik2OUVfKQfh2yflaqwCjHElVeJv9n1IQbwKtIeOjpesWCuK
lcNl4sLlwtHFU3/MbL6UDUtlAxg/YTYxWicAvkvnNZidC3niXKWWLj4kRflGabOo
ljQnwMRSqQMfG2TqQ96gFQGtB6vmT9eRSszJRAlfVFEDYuVwsbUJuJPOB8Z2G9jQ
vIt2pauQQoqH05oQtbrxQB6z3wRrcfROzVZ4nhCSYZNRZeCACxq0iIWAIGrb/9KU
k0x3iYvhQg94p/cKA36lXwKL01Xwfa4PvQwdTsyBBdJgul/ikfn1nMyftGX6l+n8
ZvL9dKKqTk4cr6LZAMMnyCKWJGn6CY9r/qx9Fa0zYSETHADSTbA5yUfzaXzib8J2
qbRCFVAkPpZIQNxTV8tdd4Nh06j18RH+PNrQMYCXJfeuOFa9LPHdTjiFWxwDSqKH
EZAn3+iideiKsarL7tFPacFa2h9B6EyX7suTon6Ei/JCdIFLF67thSud2hfnZHFd
KmLf3963Ca6aEyiPrllBlDJB/ARromTFlWgURRWbycCtvFCo8G+m44336jED0t1N
ku8rvofebG/Xk1cW1kli2bP5IktJLFO6Uw1/rlbu99BSpOHchypfiYgfezGygC9U
2BTtvdzh/j/6ZR4n9f9NBgy7q8IeRmGmpMslC7diw43Mdj3udBriAyqwEH/VsGqz
9KOAuMR2BTJ2O6qmQotCJW87t8+kI65FHdvroA6Ddjau2muArHwxNcMK7e+jj8I9
0xIwo9KZx83EZtLFOgbm7KmqX+5Ztij9FA3f2wyrHVTJlA9B9ESAfIz0h5yim7Gh
S1xAdWdrZGJPLyHIDycOquzFix1YoZszGfU9vh7k3R8VWvfotCznB1HhnqzvhJ01
lZoD41ojA+ilZPNYDwO+ghD5zm91/tliIouxFCBhLrNV+P3glH8gICvLN1EBsUEG
yjP6BeqUpRtKw1gaD4IBEblObuR6k89HFZjX8dHAZlvDVpt4CN309zc4Mwd6ze5N
yAqbBhNFBdog+yhShXcz1RdlWZLfA7clLQZ2K0lyuLlxwJcJedc7RFvEdhgpMxm+
nsaRk6U8lmeGhDBCLD8SJNngdviLXACMoVDt4C5dGpat9RQP/mc/YFmCE/IDH+uW
9ZP8eVGMje5B1gBJdG7BMjdc/EmIJvT1RgVh2Gz5YP8ad+gfNt7jECo31heCVxFE
OQhYDkzwgOGMvf5vD/q/Ow4laDyv3+eAzs8ldqFfrQHn5/p9Bg3HSQWvcsyfqIpJ
MkRPJsS8AeSbOe7vTxJu9uGnDCf9jlWqgQ65ELii+8O7NnuI17ojDZYxfFtMYoJN
6tHJgrArNPqic4ap6fve7PoxWmwhIXYNh2xg4Z7UhG+DZr9Pxy6mxBn0mirIf3Kf
5gCb5CbuBhFLlJjUQ5LP8OQKoATW8pIUFMqQSHW4ZO9+e6Mu137fWb/TATavd/2a
hQSjo9JxHHk0TEByiiX3w2AP9S6EVpOjzDkv4ILwRWLjvbkFLgTHXxh/6nT2YNdo
uzLxvCrlQgFA2Bt/ZI1z8lBKG+cNvqpz9zFVewkhk4PeYcZakLnaxsgsvvM7nP6C
vGXHEfYbdJnJjOhijV1pBRteOxIIwcFuE0YAn843h/fNKRi51GOul3O2xo2OMhv6
nqaRxQl4t0O/uJsOIxAG+hthXehpdpNMz62da74Wyzj7DjVMrVbrs5t1uzTiTp5w
Ww4mKWN5F0cYwnv38BRKpyA1umr5o/n6qEUTpWPHPIYC7p7Knf1S1YMERBK7fAIi
EoCUCWtwne3oup6y+JE+Xsb0MM+ehwKe3aRYneM4x/zQ4ojAgaQA3ek1+KyFsCKY
m+NwDj4xlDhtE0Y/mNBquY3YLMpBGBMB9Z0pET4OJYFJ50MsDcx/q+QIqcq5Prsj
JNOG77lqTY/7IjSWJqJGZuYa6k2A/wuVhwab36xwa1s7vBIK4gjNeozdCdlExVMW
yerS5/Fi8DrUPKpaO5e/fbSfU4j2Ikjqs6A1DnblVqgJA8eofYSMn294HPmnrxWc
UphKtQodQmtSiWGkWo6g76XohnIsFLt3YIbsSMowMZCfiQkw1O4f5okYwCQxoWs3
n93PDeFRMSAeRQPqGKSFZPpk0T0vpnUsog2BXqWNil7Xg0wPXbNbKFPX0rBtFpKn
Z8FiDkChQ2domUeg/OJgSjxL59nr6dWSJc2Ha+fjMRfmj8slo33ArYpgHgtDb3at
ZcxNqthWLi1qQ45jTctTnk5BJKqJbwdANmXx7Pb0D2kDCLaEmjmjGMPN2vwP7WJr
qoWTFaOlDSbF8unfQ/GUj1faC2Lu/LQ8sisUmfAIuacpVdoDSId4CUpZ3jLtNFSJ
AlR4CyiIfGRtBviYTdxmieBaNtP5yDaD/YGycFcKuQ6119DiZuIedOVOx0EwElf2
ePIyPXkmoNfVG9cZiEdw9unQBQFlVN7GepQvepayBtRevirCQvXtHwwM0R5W3NVa
caM1lEh5DOf04gnkOohWmCFXYQfJtVxVOWsHM2MqiI5tQvQcnltCBTsu8RpXyWzr
Ic6L4cRgvCQJWz0Ld/fRrjQQ5rCFvkcOrcIRKOD5hZwAFOSHAoARFvUyRFZ4uRdx
Gf9FMRb4TqEgl89MKMipcVkz2P5i6hHHLdnfyrIL3b5urFOKvmrgpJ0YJRICaBFS
2EQoq6lpHVHo8NSm9VCMze1WkP3uTUh+GLO1rWn2fF7d/EZr37FRE3rGcOtR+O0T
YupnIn+x9fhTYysVwcT1KkdfZ6TCtqsoYHGhe5uT7kOiMQLjSqMEUnIvSoXHoSHs
qPVKMHt6pVS/+S1qpptoSi5eh9vs/IkdstXBDoFoaOVrhytr5oCI80TwIwbp/R3Q
iu0EMXXfNx6TQtKMIGBnuY+NuFjk+Gzhh33kyMZWoVRRP5bkQodc9CRLCZ1aAjUg
pzeLqLDh9dWvAy2cWTWfxpatpu9jpF7/dnRInVw48TN6vPWNK4BGQZoNJi2RF1Ka
yrbTc0kMh6/X3/xowhJQoWdo6KinPhvMI0XW3qDZuElqLgu3Rr2PCtIfxzLo3sL1
U5huvjIIp31JNLjVUHZCle68eSHYp6m+mu6fCo/jsaIAyQ/gm8KjW/ln373afLsS
7/gH9jKEGtX7AexCCMH7AAXoAx/uRexHFXkBJsZ5/tLzSkiv0fp+w9wxsJ5FS3V8
mND2McDGoRz8d6DhzW8QnoxLX3sv/KNa4Ifr4vngFMUFSpJvdKJsPE+ZorSpqgIl
VQNtWwtb6/e17Y0OQW5QQQvxo5V0UZFuk1fLeX0lo8ux1n95edzkUHHa4ZalmSxA
dzPLBe78XSypJxThzUAVBceJaSyUPuuMDIWiRxCWZw3Sa2iy8RXWvOcJReXolw4A
ddZBudXVu2YJBIXyV08rpvw5KQxVILUyQayj8FeXvGtNjmBJf8rd5MjiHVoYjCSm
qiNOTNPG9+1rQU5DoyQFIXl3SgikgUaQ42hXJ3b1DyQoabWJ7kk/dpSSYGDv+b/E
U3OeWhgQM1vhT3zm/aCPDZWFQdu7CuRj6D6wATPG9xFArqnAtQBCbjIFYq1+JsLR
IT9uHGhkm1qIGBOJIUfhUV9O6nqEe3MRsWLywOFVJjeTW61BGBRwWGI7IJs5pcpo
jJlic3DBSCzH1Vv12pUF4jSiV7RMpG0mRaXyImqatQKSYYRYcXusIw1z1M+71k9y
llNT/jmOhou+eF8TgdBEfbA+6RZps6995dkhZpXeB9dVjP2sd8Ls2ZhG5cCewFbT
a9g5zyW0coqrjtnnZK1pxgq0GbJ6soLIBry2FAGPD6Vs/b3JZEg+4yOkioz9slOe
HQdkKw0RXGrYAbWsxQUjS2/uVptI0DrTeqLcd1ZyJErq2T3JkyDBDiUZfoZJF3VJ
E2Xri4hqB1lY2ffAx2ygR2L+YsdG1ffkzA+KKQNq/tag1DRmpVs1MW/J/MOcPPDj
klZka82oqtUk7NA4Qba1TSscULi4X+dvmLEv5y0oQHVUTAgIsC8Os00Zrvxw94Uo
+z0/u0kg+jU04/wBVJVA51bT/u1Q1sU+OQwa64BnH15VBVKMPlDX+Ps8eT+OUgPU
BEUCeJQ5ezJaXwF1nsCybDdohCYB5i5AHLvE2scV5C3f3RExVFWT1NRfTeN3dlb4
HrzaVKCiMjpfCHPHQoGFQyMoBoMC668FSJtYMHnzYeDjmIOX05A5AFOcK6Psh34e
Us1Icz6AI7JtQDsu8+YTnJvJqEWE+8y8qnwqv0792rJoRxchG5FcB4ap8AxrKkr5
TQm/pHarAniT53gFgb7FjScvwRDPLskJvYkVLwrtQgeGrKhgJ8lGvjIixyAbyuYu
DWb/TvvnAi/L80Imk27KIja8/7Nk42Zmucasob4lP09PpKF1MMXjyt1q90hGOkSf
iPxk6mE8ufK6McK5JZeMlTMdELNm12EpoVoRjoy/y1oyC8/aCW/oVelNr4mulSog
ESQH7Bx31QNV/dn4tnqzBnn5uKPYK2FFPy83aQ7QOQgOHbbSA7W5SayqTqkmcFTm
WlO8KQNGAZYlnsZKwO5c+oJ//mNEU4mpd0xNmG1LMmuc9oSVWGvUv5kCq73rsta6
Ef+1boXddCSv6IT119WObGiXbCoaItjkngCukjOCCwTTErFevORoZ6TkTnqenjFc
q2hc/qVA/Hex9yytZDBlLGedjcyVNRp4fghJmklP8EtCgrHizlfIpzf1Quh0tz69
/80HW/ePzxvBbMBIz/xeFPxS6ARNWYE0ZIqa3cgly8hOUcohVLpYAxhT/AlEZn9V
se5OfYumNLkYQ84qaGJnPU1TQ6B6ys7+cl52pls1WIaHq+6Hl6AGJZjNrAtzPnKw
7+RAfnSd3y7R80KI8qQ/q7NcBbgyRBkdvUDglJAmxVUmnEyO27/wmFKdP+ruT5Sx
VJlbN5akWleKr74IiBpNqneJPUZx/59FsnHyfYDwbZDE7Q9TAPnrgHQKA+OfJYpk
2+dxDzh7TySi9Lf7M3S9k/9Wd9DdR8qJaQWDWJwMGLFaS9S45CGorb6cc3svF7/b
dW7OZLcbwfswDqtSWskH5xquZpi4FQadqIgu3iZuNcwrWLQzpL0deXbOAUErPYNU
mG41zVAdme5M/Mm07SyA8zF0vXvxHYG1hOsDx5tyOOn8KQFCMCqsHX2K5ggtmFZM
A4i3o4DZt5JMcCcEDacsDckZwCK5S9pGxaqVxW0kI05yI8WBoGw/Wtlg++SO10H0
zuDo9Hb6OJomZUeXK7uQiVJ/xgmAagY/AAcndWTikjVExgLN77nPDrGl9m8NMbIt
op0YiyHKq4SjMciXttDOXebPaMGT+VTWQwgW3H4VNIxfkSqtsArmnY6/4Ddqpj0F
OYqf/JcrYkvGXu3jSJWUh6zsNtlMruNQ/6AkHB/5DHC+86nPGJ7TwMQ/uh6gUZki
WEy9nw9U0A6CbxDHay5h2Ocg69AkefCerYoVVEyKh3gZU7wvpuZ/XTUWJlIXsr/5
YLcpOLYbrGsKstoQ2ArZ/RMi4D7sTTL3qwR7Ani6g3MbXEmZ5IanJF0Cb7s9UW0I
EwNzh3HSnQsg4lyNM+e7e5kWwZkgW03qep+nb0FVidsjVQuCBMYhOqcfP0BMAt9o
JJkCXqoA1YPz6SA/sSOGHm/mx41cGhTQXkOd0rD5OsYnMfUDh0Umf1JO2naHpipA
+SIfBcjNpX6teDPXtt5cXCn8dXE/WJmya+vkQPpH2ihbCdJgwMWkeBdXQAHsY3NL
DqpHVG3LWBBK4m7GGNSfEYYLtr/PwXL6IyUI/S3Dxw/LFwTpgtoKCHRjuyLUikSl
JKR3CHRO4tkjldlnrdlkqNc3SL3hdvJyg6a0qwbA3uVl2fjqMT1naeqgjYLI/o+r
WPvLFuVigqbk5B0UAi78ECbEgBvLcUbDcvyHSYudQLkb0JtKBGt9BGlB8ZxYpesg
QgqVGNcUNK24pV6wsKu+p3JKgirz1Dg4SUjRNeePXCDAbYTio07WOhvzy22xPT8E
Wxgsf/uMeEQHTbydhUP8gvLZU9lH8sBQ/PJYEIMYSW8krqUyfPlE1mKezc2qGeS1
RVKD1entUhicUWFiHetY3LANNUZ+WD8ALESn901PyMDpJq69hrCL7I6TW7unau73
YRrP4vKu2JuzbPavUgT5EKkBc+nyP+I+g9r/HJMrLGRaT6oFYh0SoulvrO7py9Z4
cgnsHllbSTZqER77aK6nM6ikEX7u3iKPGwfkm6XcJXJ804BV6AM9JZHrNQ4F7WTb
dZJV+6zKJBKPj9RwT6K1y2fPtPdKJPGX+wvSjLgdIdLQa5bB5PuQrWJs74Jh4PFI
Z4KqSNk629QCgqMVI8F+bAYoAFi/nKEeLIczc76u9EeTAqwYnfeegnHxqPF3NSKS
YvadnQEL2D7LgmWtT0fhd2/xWuND41/4St1tyf7xaV10hYEOrrzV7LFaUzhauxe8
wVHqH3uGDkB48beko/XX4m1jLyIpJzh6f7BxB7dVSCHsC291C5kUUd+njW3OIFEU
EH0I4IoaNEBIXqciIyJGQ+HIsJRjzvN2Zt8kXfy+cupzy5SPdfP10G9WjoJ88a1c
WmO7L6FO3tvg2mZaivY6T/GZ72APpJnPzZnO9j1YndCeMxJSNGHhlvT3ZazJ+Lag
+HE25jU9ntccmyFqC3hICySQNoRW6xY5X5tBIm4yPX2FbMP/3TbmdG2bNgRy4Iql
CDXC6F/y3lncjKGJEkz5AV08wQXsGUpgIqrnY4Gfa2EroyyNaB/zxRqIhPlDBBxB
kNsrP4NyFcawjRBK3D0NWFtc6DX4ky+TSjFLP5OdvcOMiVgzNYReU4lDYVPlMTNa
a6WdMsg/E8qPRu16Uoo1mwF7UFoXgcqEy9RVIKfycZVQWfMiRkPXbdjmS8Cuonkn
adHpEH82EU+oIQ5cisR97NkbsxROi3rbNS4Hie4PyoBN4NivWYtD0cIw9Ia/bbaJ
3FwBtrenA+pjFxtDVPJDo17F3TmJZF3SKSe5nwP5Uh2YjiMZ+poIsJV1Fqf3hBQM
nCyGSyOZVxYsD0GTOivSAmjDIg9+yXbSODyAczcQG7y+t1jQSgUtfK+nE/Zqa8wx
KlgpJPJoMu7vLIwbV9lLwclUaCbqzEDshD7LNoNcwnSU7s9sxW3e2ytLzVOVC5+C
vQulvbbcjjlhzfQ+3SScguEr5TarkuI8f0Vw3L9DNiiYT68bEKyX9u6IaiBv9But
34A6/tpxhFW7RgjcGixTf9JI3OFYQB0mVRddONRu7A4agsn2ViNg2iIVCr/6mCCb
1TZ7ztL6Izas3jgwmBE2jw+S5NRB5mwgPj9h3ZI2mpxRK/Nn1Isrgp5kcuQrsRzn
sNBn8Xekjz8Pu2y4G5Hbv3AtUt12ycKbLM4XozTKJSKZTGdVNEW0DBElxtyercP4
aIX7LRbxiMWQ/WVuOonGjE2zQPpj+r9GXCoyVtAFVOv1w6DMmNhYN7Zd2G/y6z8F
VkknHF7ACFpHK6kiVWPxiYXQR7Lyi63NInWyiWgkNvuort+f6431NfMTw306Z8fm
fSwo29hFyvSjZpnDyGVGQWv382PkFy6AdbdJg3wKg/fIbwXs7yo1qPz/zw/czUh5
fQ7rWtla/YkY412LQCcnUlI0cTWXDdkBIDPv9C6tctIWUhGLircc3VOM7Xo7g7PE
T/7mEGnQpfAK2deq7ZHec+8rM0HWzGRwAKek7RnHPgWutuXsKUtJ9O1AlRxUIg7H
tpCiauih3MonhX3Cv1l2JjLmaGS+RvVZe3JDOBQXpZ6wNe03eVd/JQb3bdJQCjvY
BMqBNK4PxQhuLFxtyi1N7quagEAQF1ia9w2B9Bf7wfdlvKmUCX9QTdHSRTdWZ8Rq
DxZga00207ZbIsbndrVpQlnjYtv5NvkKo236AgXDJNaDqxHRxnNumRQ2J5akdAN7
u/fkgMg7ahmv5zK1Rs5VM7h/A5sbSpAYqAPh5/22+kJLg+iI3hwRLu06gBvxUnwg
9TelYdod4jr84BfawaecGDQywlTntQnGRiWHh0flxE/88vL6xSQfndWB1sHqIT/q
ZOIau09FiwqyRSj6tT+vmmBbfK/gpkD3IqUPznVxJ9qkkkjoOHN6jws6pgpsTUx5
ciMdOHe/JNYfZZyW3k0bgAre90NPbNdfmj3+c9VH/PTbBNLvBZ2E345E+sLpdP9g
qMOFWVionv11sdPDUEjPFnQj/CafdWSwrjqbz3fG0J5da3TucP1E4stlLKknvbOJ
JS8+1jalQXoSgMdYMo0WsEM2/suiteGuHZhPDhgrEPQWYbV4ULTga20dcEqTdyLS
ZBHhk8avrxPJS/ofZw+N/wvOnpfxa9F8HW7HPNZjZA0JhzASrBCm3Ucv3S/bR3zy
1kcCAu8lrnk7Nf6hW3YHtgwQEXkie81+Y7Gefb9uI0jeHeMfpCPpc3VPbd2ecYU1
4/6MzgkFariqAQ+Ua+UbCCRzI2AgZ2pV85FmemQbVuLXLR6E1LOftP65unirTFe5
DhmW6nf1Qyh0Q53OA2yeu1UyWGkkPZlYVCiD6QAnGeP/CW0akEXCl8V2aKpnUqtW
Mk1/VyCzWpMeX/bJf4Ala/6gXP1pDD2renENToUK68QfKxgVwd3fAthtI60lwoRW
e51dt4QQ+/SmGpkmG6rBw4G0Rgl4AXfLkiVpyU4xHsWIrDBLxlST8cJpZVfm4DPI
gDheEMXUR4Jws7V5AYxvPNbtkLf1FGYGEKMqeQmNBQTE3aWEj3oSLnC1c1oq6t62
KcnkIDeC0X/VfFFiYl8PrOnB/UI03I9lFEjGpBQ01v/tC6P63gYC5isUREpyE6P0
qAo8LetyFim2OA855mhKKYZpeikQJguRs/L62hBX5pcBtL8FoKhc86Y/SEuwW8nE
lmcjrwVV2ZUfTPd8ND/yRIjR5fCj9i9721/XPbKTPjssWLu5RsU0UpP/4PUliKJr
6VxLQIfUd5O3C6vdUJNekH++UK2oOCJ8Bu5o8s1pyCDEk7A7AEuaN8Z5fNuygxX6
L4OrFz+oqN2aCEkaI2vT3hjZwsyQIqmHqVPe+a7meFwufIcHwbl8BrNBnursBwUE
y1xkTd1XKM+Dz6LEnje4HGZegO6DxLN7tp3cUPmUVpSGWzefXZ00d+UUzbaOlrRU
WrhRAOg8OnDfJu3TrkkonpK+/Ysnz/qEjnPwLJGEwnonKtq2aKSNiXiT0WM8f1Wi
e5/HTaoTrz0lPPLjYdApJollnbZi3AhLBTktyn4hNWfy+80BhzfunAs13RuHpMz2
Ga8dQrFV4vCUcOWC/whLpbiEubYUN21PNmZ6ucvBiTmDHRP1ClmiJIu3CNqNKGdJ
GKP2Q3DPirzx5g958IcvcbxqwqWM7MRmbAB/F5g3pLLyvGxIFhMNo2ZFtSLR9pQH
bFEnYobudrjnzxtzoCs2Q8XWlfgpxcMfPdE934xyMdx2albMD/q8VgiuZ9VGnKb5
iywiEipM4IaH9fDrPvw/cVRejS430PGgAFNPSg4GWQpkpJuCqImBnHP0A4Xp9chK
twIEJifFZqwrzP9uVWYMB/fO7tvDxRLwLleWSxOLhe2VGgAx9OkEf8qAfpZI+Lz/
1trD7FrelppJKV9Aaq69fd5lLUtEUMilzRJGkYl6zGUeIFWOkkCFa2XbEEbuDrIM
tEj+JBzj/tuJJArxkvb3xd08ZGCla5igskEbrlLAEeZ+EHWc+2uYnkQqRFPa4K6r
xF31l0E2A9CC2OZDGk5I7f9/qAoVjhdaMxq9VSz6MkfithU0HsyosQU4ZNvPQS7G
cXBhsgzkKVheRfYvRPBiZPzXUhJAnKirpInYf9lyvthIg2kWeOlqzROZia+Yb0Uv
57i+0yNu0otTQfhX58CozOhXALIkntjamdF1JbRP/DmpmyBcxSwx4p2XbbCHzbGX
AgbwsZLxxvEesdZLnDkboRxM466TJX2FiAGMd/97JhytqsFT/JLaPiKHx2jI992D
q2d0GfSd0ZkKAB1v3rglhu8K1S3i+0M03raKNWCmR+nHFEoL0CU+5WGSaNUAhdaN
CmuZ+loc+PSXVWeqo4hmiU6aoBnLZTyfnhTLQ8Sw51n4QDIYQF77Uoj8T8kr9639
hdJcrglki7iXJuA6yQCnr8mC7K4SCGI/oJjMwB9F6O2avquvUIw7einElMWrtwk9
Bi8g0ltRx6/AKhJA+m8PtL9Su7dgBqbyx9J81k549nm0c9rI3WBrxf3AGT31CC4h
w4BmiusVUARp2gUBVDky349yXYk3AkwkWfMU2D6fIHUu9FNAPy3ZS3ucwdDXSO8G
fBX8sQfv0lKpTi1tqoPfHGtAdIGuGkrUSBkVctEE/odDr/pSP5VNJEkN0acpXR8q
8Ig/2GtDPsl0551L1DmRb5M8ZwgvziBA68LzuswSBtOFRs8RmdufEvM2j1J3oVCF
excI2DgXDJ8eKj+WfAz4g5o9gSb4T5jLEAbF56zyU5pv853WAlJn6ZK6ARRnG94C
ww5HbV4t3zUKXouzrPw79xH2jH8ao3yLzTa5f+Yhqj+DpofytHQHnJpmaKv6fmsy
qFq0IaTHreHA+kA54QsTGa648W3fDQBadcEiRulaSr2bisDZUcNlFPXdiydmXT0+
aR4082SnmpfnE3qnFKnZ2V5jodDIkQr71VEuDihjsOAEO/m2FdrCgPCGKIwlzggg
h2vJzJOZr8/Ibw447vMCaRCYUFjYF9TpIx3shbl9lc+U6iIkx8w0f5fSo2oAeKTY
Qsy64qHz/qLqznXBOxo7f9jr68D8FGZw9vE08fiedpJEdIOJGmOGH/k4Bu0DUqk/
nG6LtQfFBt3I1y/qDoKqJ1V77C/wjB73DFyobUAMrpQRTBbFTiWsHJQFUeBJQjk0
EKlUc0kyDL8amfVQXyqZcsnBznsgk+63VzGdLa7CGBx1HTiFPxjPCIcCRntTdn2u
PpzabTLeyRMs4P+fkCvLQYDXWPvK47STS031kbd3T0PGJ7JWSp2Ww+56GHxci85I
525xBMIo/OOTuJLHLJFvLXUKXS1mflER5OlE6x8N0FRWjelFFH3IUsYyjc+x/FZP
AvxhvwGLXVIIllFdzqN9kvCjcbetebg9IjrzV8ElaG3iup8/bWqi+CP8tcdM4ydP
PSm5rOcv2KGdWECa4GmyPG9Fh9KcBF13Qgo219a/MpVOx2b7c9auyiZSrm1La0ks
pUpji6CEOA1pqEwUkgKNsIpw15YLxLgIsO4WrbWSpWTnGx9B96YZlx11ZEnCxsYn
BlMyBydn1dZADFPG0TSs7bjb1z1K6/hS8fA1+uyP4u3HjY/iZVXQIdfQlwm/vp9C
m+3aaIqFPm4S7O8+NmJJ7bggKemK3r358QorvW4h2og5g9Bs+Wqowx7MEF3QPdr2
MLtdXdbuCaO0bD9T3Gh2Dn5nu5CxgPoSiBpudhHXWzIH5oeME1BESN9u2bSHT5IC
OCUadXRf6XCvyn5sbrhu6s7sGvsD8saExbibjwiwCxx2+6BqxUc/LpY0M8dEB8O3
Ew4RRxiH+zGL58xwgFCVWW5621lOYEGFeT1WDh49lDe6U1IG8/UHULbjYz+PGFWy
xDXBZT6D7Ak1w/pBj6bfRBvCesb/7Ie9MJ9AMc042EBNwbMxaGWTAunRBzxF4Rf1
O4Fkdgq/d1W/GSoEsfHvyg5g2jZhTmEp3h8oYK2NNvRSBWFPIV+SeZg79YawSUXe
Qay4MPjlsEmzA2dbDAcjcTfziSoe5/w3qeCyi5jLz/XOFPXTLP76cO+7MjKpFGO2
L3f8UyJnwAfKtL8frrDtY1wKCFhoxrBP/dx3KzICpuyUkJSAAS9lZ1SNuHuFyT7H
uo0nrpfFmxj+m8rrE0CbdJbu8DWoXaKDdM+aIcUc6OZJtM7tAdIGmyxPT/Yi/DJw
zEKb5paNrhdey8XEsA4pykosf67wlmJe7WzGe/q/WodDFKUN4q8w3OYbk9/RGDCc
AKTagmOPL/qJ0pkWxxPblTyeFzJcUJOw+p1FxsQhqmJlTpLz8FJCuOMwjYAtxI+i
+3+FJdLe4ixiVYT3FxMgXJ11coOJfN9Rfau7gBU34R66eGSKqqvJfmeflng6a++g
SvW5AmFtFBREM47NcranQiarDXbl/sQr87sAal8v/uR+y3hcE+nIHJI6y/qO2pN3
RWJ0hj7GQIT2llY7O1uE7ssphEV5+YvHYEVKRlGNCaDU4UMHU9O9gsZImQlduA9+
40auksBAADxK2a3Y11ZeNfN8/UdzforerFLj15RGZyUtZxhFoAJ/z6y1gZD8bvmq
yv6KPevgoxWoE404M+akDcKnOUVoV5a7q2fTtgsU+8PIu8aHig7HpVdhBNqCRjPz
VaPaQGZCiUMRYKmNSx9ZROSmDVWGr+ZNBwCCekMRkNQMJA15XiKlAWBE558ZjgI6
hNLhlgQMBJU9k9AKWEdlhVABFmfS87D8Ibsefzh+Eg6+88C1jezSU3Vg8OxidsZG
0cxDFCzfjsJjGpAglg8huOW56fMRN2dNstH3FwS1TZ0zcMSa6wmSOr1y+8FiqiT0
vA/0jIQQLfbWgxaOMRxI//LQfN1k0X6f/TtUiw01BKd6iWM2oCIsIyOaIybrBq09
gGv4ktJVFcx2e2XbK+8p0Rd1OKuyPA5PLaK5rSGVYAhEBhpZRuP9VQedu8/qEpxP
PFRNA6Quz/Xz+7wjR+8RdFe0IkHO4Q+971FmiyAF4YiviLJzxWY44wZU/eSDhUrT
1zUwA4T9Idkf+05b+6SEmUdsHRth2MpGytxiL4PNQfBUBVx/mHry71r51rkipxAv
jCs2RfxQyPh1EeURUpsukfL4ZMKDivAEaSPWWQyB7LKL8QXgXtiuz8Qz3zNXsse4
ARvbRpltxmk5SgygHQZjuf4RfqW0j/YgclvB7uWwE61zt2nbqiXzqxe689M/zfH6
AoI+zpJ/x11EV654BjkBP8i/qryfu9rN4tYTcSpn1qDe3P+1a/zYYdBQIB/Rh+Xu
rp2OPSLaTZ/luBJDhLOW/SOids/Z5NJh99vxzDvBbPyUPC5MmV1aEjcbLI/yc2sU
jEZ9M1EWuBxyrn1IEIbME4sPS2rewwsHRsCiAKYsv+VyFosLcmChRuFnv/tsOn1i
hAAIB5OO93665ouybUHkLWyWUv6/IZehgETmGwwPHONC34IxGuA4AlaPbwzNA0TN
BYxzWz0sdscqKAIOgrwFR/my/cOFp7icDSiEcOPN3EgQmKQFRCq1czbbb2AtQWC6
o30sIsf2h4X/gebR3ind2qDpEMAfalLHwU/LNa4b1vR2z3K/A+FvHhfVfEwN3QUy
P2hlnRX2Cn7uYnGF/ubQfFzMcN7TYnw4fEHZwWs7r+uMADym14Gvj1M21EPzQ+9q
ra9VWK72kRjPDlGR8/LwMDysrX9lkib+cw6Cc9jtFUg78xrsI1ly1v98M+bhgn/P
Zs4QwfUrlxrT8B4TGkIMlaPp/tLZdeXjk5cyo307tH8ql0IXMwy6CeOcVUpxjaW2
oOIkkd8pvLeZX3KQjly9R2JyC2bNZD7CNt9IxF/HHfBFYgIismBkWjY0JPqtMUP6
XETFRcYvSui7C4uMvJy6DC85WEFhQXWcCq9/T4d2XOakhI92itiVJ6iYBVW0dZlR
KYQ+I3lxdB7B0dmKOIJxIvNkjbbzs0ZeR1Z1CXNqYd5cQbVNLIVz9Y/ulFZBwnIR
1PqXvl4OqX2bg1FL0MFK2qg2SIedgRwXPF6ci7qNvwjnCI6rGiN3iIOxP6B5iKFy
diUsgFpMpCBCRtJGT9ZS/5nVN4j0Ok7Cx1xsWtTf8JHhojLcMbVSykrcktBe/doh
M8Z4LAoRG6Z7BTzKmtrBc4Q1XfDIJimRPMmyq3dW+hoZiWwAmy+NpOoMAJAkgGba
b1NBdmJNoqumCafDfsYuLVLYKLm+b089DpTXq0lTUhrXMcR5AzC3q5pRf/mFSEnB
BPrc693JfGG8tGOMTLTQXz5CeiWLxn5O37HlO4NnhUYqpHuJ3cAnNuafFPrA1oxA
3oSDzJB74TLVbqHuGHs00ZHIDp01IbuL9W9P2RpUyOzXTxdg2+XJW6mV5tfROjJV
tIPgpkqm04kq/TRyVQdpf4+9q7KagyH9gW6RJoMZ28l+ayIwjFJyquAMMOFVKJAZ
GHaknd7+3I6DBd5uDKJKV7Y5868/ZXf4M94TAQ9cY/sAzj3dpp+9/SJOwNSDK7z8
s2LE3n4ogDiVXj8HUPL7CLN+0DKax/1YyyQptZF3TtCLS87mEbNIbyP2vEzny72l
jx8xwO2H15Nr1hEytDR4D1BC2zvSO3sxS+LDfjiSATnJS3GepsqUP3ykc8t49xau
K4ewIiMpq7ywIFfX+iSnbkK4wEfvndWL5CDQc8d9lT7ZbO5ohnd74RbvQ1SJAVcb
NkLe/2PSondQkn7oXbdy3EcUgSu/RoNVna9UBLrwn7nFm7yWWjx8oeKdom9FwDXx
avudJ44l06kLFPATlQcfidiYhp4Q0IN3KvffYjbrJWjqz4N0XoopLrKoUpgsYhf+
SCTRHTG3/DesFOyo138V0rvsWR8jOWsPTAgWSCD91k1u34rTqPKKN6Y8El0B9G2v
Z+6nKMAXv7tPpuuZD5d3ga+NeQ4waMNC+NCkk90bAHOnL1G6u1wqmTclv1oAAXoA
xCaTApysPLQxzzLGkch7QICgJtjcRZ8QlhMcAKsn/NRGvu5QS90FH++NrEDY0VRR
WVb4OPNPwPdo+1pbPTU0wOYVehj780X7VU+UyQxNuUeRhQpgaIwMHC+dLZR0cUPT
Aq/rAoW/fVWAG4vjhTRtoK67H6+Ihu+DbbGONy1OYON+Oc1dLmFVB4X+x3Vcr2Hr
P2teBssVM49ZaX0eOh7GF9UQXNh5zEd5ZVcv7aeMyNOtHOCgC7Jl5YhsEET+l9vz
ddaVMtnrO3PwFJi1RTVIhvdyAduADVilVmXZBj2lJvUuen+/19drP9CwS6lYi0Lo
E2UZWwFAyegU05EGGEIlKLma9UIdQdWzXM/QjhqkDP+mEmfCtq7zAmH2Z7EuljV/
qsyrB7cZrRUsYF5p8FzyvEznR+24Mvw2tXzs5kdVJYW/3/VIzcYJvhCuCJgJIDlq
VYE20t1Jejry8mxI1ybo3y/qXCyKnFbBGFYgApwWxEt6mh+uEdtA6Bn14MP2+kvS
GtjrTLSS+bEr+7fSPdLURdD7mzzirxbFqqbOy3h3EPj2OADwFDCEu0xBbhIelbBF
JY6MuiwaSbUJKeMDf+wpKST5/USeLu2LALZLFTNuE7/NhfOMIM+equUWVVx4Ux/n
XvJCEdV5rZC2LwD3kj4plwo/404pYDnr2vaZkl8rSolZoQATeKWnoKwuVujG9Vvq
9BedPKLh7IhGWAxx9oWo4F5Hvc3BjppMm5tSbQ3OI1stJotvWjfLSD3s0YPZ+C3A
6BHONY5HNSVIELTGaXz79Jf2pmrtDZnZcMwSwlX//xR3CI5qW6VGfy5lV1OWjbZ9
+0KFWQFGeufUfk4LlLr94xUEBtv28wC3zNl4ZkGZXUj35vxkb4qiRdZZFm5EXefA
2aWiCv78tjm0ZeU8RIcsNQOsIPuafxHmNkGwMrXtg84LBvRmNJax9p2/gMpu+jU2
g+KtsTxh5uKIxTKl8bfQpZ7jKzj00DrPqLodIbLxNeTnUDHa3ECxulA13RU9aCwI
S5uQghqnoS8MlQAqxgOo3zhLqk4gYeDbv+IcC5LmHL761mhL+7dHTQa8GJoE8Lt+
ZSBu3eIc3MPCiPxpKTbAlRvNyrICMZ6yjcdPuspW5IfKaBBzIYcsGS9rBlWE6WUl
FkSXONmWS7aIflN8z2tTay1YF0NDmhzbOBacZH60KsI0N+WDG4WDe+/esT1ZAsWk
El3T7bDBGxwK433HXbQigKzOPrn+t8/IOJm1lc0/bdhgjVzuwIz+G0MVq3Lb11xT
J5/J3g0S9ezoSbgvVX3WeN8197fh9ZAiXJz9xCtscLfVtnMUg4JNuHZyTMWpiEJy
rmSppGWJDKyg9LlqlrjryKoUqI6/hRWYoLT9wXxuSPkZc71eOxGM10IlwLwMe301
aUYsDmIdAs8Av7TjetFOX8D8d/cNf4Nw3A1457Wl+erHBLuzZK5vpa9X7nT7u/Ka
EjpXo97wS9w50Sl747DPw/MP1CPNpyiYDAQ3cO7sz7eIaJ9E69vdh627R5qL9cBJ
wZq1r8HfB3Olx+BckbyNAo5KiZ5etHT5bh5Phv+KnbO8nrKspEKstas1s6atopi+
5I7KwFJKbk5dZxU1oOO4yVcIm81Z9k8bSVNCkm8QiCpCB2KrGSWuo/4pnH3IsIDd
f7zgvvOd0oLYrz6qG7sH0bVAJ8i6IUh5+DEnraA3/z85vbUkDcGNq+xE1EkZmbHa
/TpxIDcWVP3AwjoFyKmbwpK+SXgfQFP78jYrU1UHTinWnyb8iZ+zfT/yf11xII1X
wbwKal9aO03f+pAvlvK/cVaAEZDMzoP5WnL5zfSWohI08xliWvQMXQnFTZjpAxMI
jzxODVM4Z0ME8Je25tt+y6UMNQjjkwyLyV/6gay9JSj5dejZkLTZW2OZPfHxekZM
SZRTJgg1Yc1vQQhO8P9p7zzIEfT4xPXHGSpGSvo6o27wwpdw+FhiO0CTEmZcpORe
VBBLKQ4oqzjJlFuaDag+t7shVILkSmO9AxNKxookAhuJgoOSCCPKpDjQQJl8Tt2R
Nn7dklEFNs0N8zUNM0md51h4hU1UwnCNPhdhsS+VNJ4ozbQY7l7xRh8dCWOvj24L
3u7AiqmtwjDzUwDuFayons45DJ+2BkTI7czUdhaNOnMDjc8zDmXAPrfNPJdjgfPq
gG6gNJJc7ySr7emWMCoDiI98R1FkpRVKwM3xv0J0+IGp6U+PzBe+4kxtS9izKREN
fN78+pRuM+6GnxtMr9G84oWwFRYqK2QHXfr2RV+bVCyMj2VoYKyIFgXEq6ZGyIWB
I8xV3FtdzyW6zp+HfH4ETSdoG5dtJxT6XqSwjCuzgltoDxOga3eHeeLwB+p6RL1K
WDJMEM4C7jpHEYeDgBFE6ixF3RwowHMgaLRO9bT3OQdkVd2ggTiv3OVNvLZmS8zL
MauiLEySJIP6KA18LCNzUAX+HUtnFyuUYzMnv5cmzfes0toL1nqqaYIoX54mb0fN
6VZIlsyHD+7h1UZkOTw+627vzea40SnBLK1Py/Q4frP119dNH4FWkdazNrXqCo+r
8p5Yp9RzmU312cTMYzbt2e+uXHPxgxYKTgrWht7076o6ZJ085QFqxHaochk0lGQP
5ejaoq5xRxI4FLUAKSUogToI4euU3XoPqRAuCJzBtMozRXphETHX9fSfHg/DlFoQ
AuSVZM8/yDMYADOdrQdJ8N/YzQ7te9wZ3sdVU+6va0GsTn8489HdoKu4Hjd2xFec
u1XVE5cCaZFyRc0pieMK8VLt9KDuDOgM2p3suPcYFX+7QfAz4FmKHEayrmOK4KDX
x+neR9p4QiS8cC6WDC8YB2z6zrPS9NpUiuQWf7lpnQy9ds3VBaeWA+SsCIj72vq2
w2EGCUZqX0k7BDhx63+mgtt4P3i5tKn6n2204cjq+JJLELw52Awwnpkr3vYCjTFw
jugHQGGdiTsa0w7pOJeWUNm7w6wdgcrmsuivudlvlTagVMuGvp6fRHa2h6taRhjE
2lnTmCWwEKE2y4JKLpQVr6T/oUxcXEL2ZTV5sS9I2Cj/Gl9FgjJOkE50hxuyySnN
v0uU+f7rguAZTlMX4y4xTkvkZIWHePnVy4cShZiRuW+94MuIdMja2brt6A1ZyMHU
De6g4t1UInYqtZKca8Pz7qITWa6tnTNTPDClJ+KzA1uXCabKnODlROKwvu5mrg/K
/qg8G39TTKO0gZuJNhuwXcXI5T8VsOrGmbZBsG9qDswAtZyvnNYqrsIKdxbK8eT6
ruCxHmOn/D5ZVmhekz566cZtpQuRihHxT4uxJ01nW5CwgsuG7LCttort3MzVuAIy
fn9APNL2yLMwWTZkCR7M+PmL8Fbg6MDxAR4hXN5mEO2dW5EHMnGPHJDH4/K0WVdh
gyN0I73R4cRcwEPXFmJm9Y459Z6f2eU51eW6d2YvnsXpG320fHgo+VF+Rie0mc0G
Y9qTWYo7TkLCtpNeh4TflhJNDYvL6wzEa/yQT5PKY+I+MwCEQrCeyprugIniCTn1
0ByTAd+cTeIkRJFKPSZe5dnPJmJQfIHQw3OlKsSwXjAIEAHJ/XRoPqIkdqxsR7Xu
1gOAmFN6IF761FrCiTrw+hMZWDZo4WxsjPga4F6L1iJT1fkxMQZwcMDgyNyjpFkU
2jTfyWNtNUGKMVCmQ3tcAz3cChHCMPN38KrO8MrpVXG/41LH6my3DWLL4n81Vojz
QaG0f9RE1Lm9DnMvsFO8ZdbmgAlcMDqa+rhu3inch6XXy6qjZ7qY+TZa8h+y4NlK
Svl10jKlXDrg1GWVyWo0ZSLSSccnVtcEMvnO91zZWm56v7HBmAkW79YtA/Yz0EhA
h0kCj8UxTxUwkm21ZuMNzNjj8FajhmewYUODfU87dhJAdip72/r+yDTOMYjld4y0
+CcnJ0jxLlRhZrJ5dtEAKIacDNJ4VhecYzuTkrRS9DJ/h7W6kkboB07UgCG5c+kA
XWkI1/NHD/KwGtwkBmQJqeSP1NFrIo9iLQ5bVj+fwXuZFFVu2j8yi7gDfRJB0pN1
qZRU3uDdyyVHit7cMqzvq56ylE4tk5b/pRGLBt+Cqu9hBeZoDPVYtYuBIBuww7C+
XcWsohB6TrVhhcYt1/mCKhsqJ99DIekAWGrB35o8Ofg4QqOdJK1GYzcQU2e1M/5N
obRXKsaiTx7CjyM/RdlMlME6IiW8Vavi3sdlkMGfoDfr9iqmusgKFJI93etk+28Y
YJXbGD3+vIlj0P34gnBuoP5kbSgESTJRjn/seawnH4csUtW885ADsiJRFeEuBgvU
4vd0sZup8X9pEv4urbgDZHDXc0xmF+23WOWKLkFEt9r8CiiL87zisqgyO3A6/c7n
Gs8K/HdYlYANAEz120x5DYikO1NiVUSRKzmos8qOHgg0CbE0+DI7M/ki1tmFNeCf
4xhcJpSss61H4lTxsoBVIR9URM1ougkQuAf/5vDshHsYmcq9+MyYakkT2UxV4azk
VDPN8N4atkkUSQqi9aJ/P6W9PRwQkIFvirY+QYRWHBjJU11bZYdsA3J7LZX7cnqh
zl/pY/pXkPo1kdW6qcO9Wpn+YdfcFSxTX613PZL99he1eFUGXVhwWxJBdNrkkiO2
0syBl/PJ1I+l+64+0QlpbqIETcyj1YHjs9ow/Clc/o7AR1al8RkTPEe/aqMkVx8Y
00oqoISdRJ1hk8kSs2vx/VD+cXMf91/kqZs7Cx1BC1TyFRgncdCgXcUkF1fbw8ol
RoesHEsu3Hm0pb1CP/6Tpn9K71621tPkRYJ5MdXysidSjxLLkYLfyvKIzlTVFvVQ
ayklV33cwkirWk8zDMxUkjdp8xgpxIhJo0BrEDzECzlygdCjFH77AEYAsH1oushK
YqzSRlRqzDMEt2bTax2hABDfTrSjeIRru9CWvrmGKqokGOact+broof/bMB4LYk/
cc16Z82wrbARGQ53dDIh5jOV0028MHsUTI1a/CB8Xs14lPUPkoKQkappTABvu0nL
Mr5A7B/jgIHVrMhD7Gs5cI8mz3cjp2X25N4xEZxdMm6O6EDZw6MRpRvPcVycIoTX
rrUVYwQqU9yycZW1tVqIXDiFXkFOu4EXXTNPSHg3I08jsIaSjdqeKMQgT3gs7adC
LSs0sJsXV2ZzlkH3Rwt2uuiVjOqzTalLx6LkH6W67RPKzKnjLDcWc+6rknodb+N+
Yl/VtN8rB8XDFYf2z7M5CsE1sEimSaPVlUmx32ur4yuMIOzde02cT4+6C7vUn0CE
nySw1d0s0617UgJjaCtggzHT9xWKazvCi24zo7Ehe97xAWJeaQygUlBiLW3KfVki
rvzKH8YW11nZ4xFjV8LTxhZg6BEJ3N2OjPuMIWvO2H7hzyTf8KHwgjF+4TxjJfUy
PIHgsMx7R6P3grdY34qi8sUz+22YxXGQaFH0KD/7ZoER43nhQ/YIbr1my+fS8ZFa
ey26yUswgLzj3REYN7OEY5n0pTpeH72JPKnCd8ZzZ32SKM/94A5TKn0npUN19AlP
cEoB4eWPSEVX6Pdrmr7wH2khgsADpahSCbGljiZbP9WTP9eJTLaMqgWwnN0+6FJx
MYbKq6qhdy+Ke4FpK9g4jzC1syHFvfIr1gLpqWsuqfRa8DE6cHEJuM+UXiInLMSt
lbJFoRYhN4wO5Kq06AXkqsvuXUgD8cRmvaA8FvwHcQdmGssZRzrd0o8EHnKy8M8N
chbTfNh/ic3xcgTRx4sO0GJwVNFb5ipF13DcNM+J4cc2PJZt8Uc6jr0IT1kb0iGu
KZ/qxD7gH344936uou8XkPVvIM+7rDfX9eMy9/D8RNNqS/A9M688SKcRG/ZBKcmp
r8LfcNIx0loEb2hjRCTUDee3EZD1EWh/mG9ftnWnZo5GtHzMd5xipnfBECFzczON
ExyLjUz1o6UVFyQ650wpDRRZf50TH3mzwRa5jSCehad71JCve8k8oy3+0sHJizau
UH4aklQVp16i5JE9awcLsDV0lWwckkfGUoP70kjG/CpOUKCfUJpx98d0U89MYLMz
pbrPEjOsFU6p6PTQbE2oz06RWXA1o2uX7LlsmSLTeGnsiSwosFKy5G2pKWqIdpDG
Vf8sADghWl03aYhAM6khXX9XYcPkpAJ8EBO5I7Mrdu+qeF9JFozYwU3RM8xYjYoX
nkt3MZfyVZs7Fy566PCCfeg3j72ikUl3R28tqZj01Zvx/Zf4hTsI7W785lGQGt1v
YY0It7pyDoeCUvycWXeSWhHa6cLi6Ae2RQI/IQF8h9DxPi2dMEp25OgmBoHHAN9U
A8GD76P6UBYkQQbvUSh00aumR5NeIqNLPgl3zaL6il1f3qLGnTQJFhFD2nA/N9n5
IO3FhW8dXeoUkslx44SgOOhOKGCmCl5efkcvmXkPxig6Ov592fZduzS3yhFHBZ8o
k6GlDFJ2jsIy6pJAzoFFCfG6lC/ClFektf1DZ/CMmr/ZFOXf2K2DGkBZbnoSPaGY
0hhjFAQ+VuBrioRnwI1tQOQ+5D5sU/uN1ZOKcWqYfg9eXAGtwSFv6vdtcqkOPvsZ
z/5fLkFi6CSbD11v69O/HcwTwxOIWhhISXcxC/x0eAb9WUWL7vK7P/Vmfq5JQQUZ
qGPY8qxIZ8wuJHHTdqIkpaliUYdG8Er1UWBWuqe6Dd3BSSJm29+MuJlvWzUyMmCs
Z3jcot4wAv+Diaa9nvLr6u2hHxncMjgXGcfPWRSzYaNlnJLqaFS2ss1+UMuqTQNO
0w265VsN1dMKjT7CbeTKEsz1+MzSqK6XouFrSF5FMSvaoZjGROJhgotv8C8A+prN
TZZH17+nRoeJHTs7wQxb1CWSEMu/jzCd7oZQrF1V0x1fh5IOWGIBQk+ziYdZ/C0I
IyNNbXhkBke6vvrG+lHJPQTorBhntgjw/F5iUmozaP4XAEWfnn5IRYSm9Frc51Hf
UFvqY30rOX9VQTvBfL1Cd7u5K1C0XI4GrnnR7Dvhf+kuBmDxS97ISvDfS1q7i+Q5
PfJf8DsGwUCDEnDamwTjnllgA0I/3DWbS713bCHdqIAFt4hhv2NktUOu3+q02hae
gjiMSAGZm0M/hYbVdG722wcRWQIgZCXbZE+8Ryh7xSX6MeZJLq0vnJdh+bcDH37e
JhKLKqHlyk48VxnmJnzGOhP0NCZEQGLi2irR/iUOpPxwbIFsKEVc+lctEghb0qT+
xtCYioXwrRRJZXbc/FdX+V6a03heRcVL9BUXK+w7LzfeFZUMCetku5QTOtLQd/0k
M+kpaRLS4PdfdIJotbUAgBZOHSTsuSkyQ5iMvNYdSMlN4NLj/7DxgpdjZM9D3KAi
MFrmT3CM1w/umNVKFJa2+n7ETx1Eh/mTIhYrGpPELVWabeSe2IKH8ZxxiXe7AyNP
jjkY7IYem9tiIZ2RWPDUKBX1kXUZf27074IPXApIRrljTW9k2Sf7cVDW5a+su0J9
BjD0aXfjpxglLyO1HLxjMNTVIXVGg02gLP9NsCdDPY7C1cozT9ZSTdJN36pHrP6/
d8iF3xJv3mAWrv/XU4F8IvmitBnj6vIGb+7fEMwI1SaLJCzThHgPZWi2PatOUPE3
WzgAl3nHjH/M7l2rNmD1rJjzSj0FO+Bwis1waTVEP9xaxPfpOAo0x9HRGujefcuK
G5wUcWvquOJckipmveUbeUUdkvPdOlqK6BRNElCLmY8T1nqFn5I38WKF6yMC8ouH
9XTwupfIuEX0pBT8eZomvMPMjJO8yRNNssrAb/o5v6E+1RNEFDCzPrJjwShsQUZo
Do8bDQkXdQAkuH00clWe3RADnbCgD9sqk7Gu7xiyYUTeQMplvBBqHkN6LwUsw4yp
ErVJIkvqae78Jpm+Oyz1Wu8eYsNECPy3Hbp2PeBv/24s1rJFj2lmE/BEl524u7V2
VOh/IRSn2gIw1Vwj1so/91d7HHwH1Zb9ljDJ3Ut2Gijc13Iia59PYk7oMsJMEpTK
btnMTCbouHmQOPzfD3IAhqj4V+dfM1QXu/gh4b8cMAs0BmpzZ0aeIStAJb2hjI/1
c7hZLL435fGzSDyPE0BfNBi3RjpEmhyRzwQ4YMJn6yyV1rXbebgpHBNRju/peWas
Xk09wXI1BpepmmyySGspyPPODboy1LjUpJ12CqXpBq0uioXh/XZKURiqc7Nes61S
rjec318Tc3+/F+XQQAJ7PeKa/Lir/Vp9ef3J1J82HpIhza2k4FCawx0MCuBS+7iQ
4Ht6iF3KCTn3LdNzzPTMp6YBVP85oCzQjwspmvLdncNiHLY0eADdQf3ijQluI1lc
2+Y/5HO+RD1p7csV0kLF9Caz1mNKxu58rtgGsBElUDt8pBFK5FbDAF11GkeGOByn
2dilpY+9mEH3/RVIyjWQSNc64U71LaFzCAcxSWHwwELKRUn5avBum45r8I5jegMg
ZZ5FKCPYBE8JIF5+aTy947UvtfEGeVWC5IuZgWjkTj+SwTKCNPJ2u9DLkw7/d6d5
JgZMMvqKJ+zQuljMceZIXtzel+MNS3iIRwDBTQDTPuuKnbbKCEfpY4vQ1e/DtZIS
rXl4bD076brnneKNTk7J7fhOaSRmHc0xAl4S/kSHczQe1fAR7LxOCzSj1RltxdfF
VRwig2Sc3CCiJiLfoC7Bh/dxV6q96knXVZIQyRqeOVgViWvmXcTyUzlKu/74I2+n
1baG9XhVIaiZFg2FxFg5hWUoUsZGqidZT/J9cm4xVRV0Gv1sC4b208FhMjQzivZj
Ujvq65crNUpMVM6//mhBt9LDSOG1C5f7UDzbWOaPWHsbxufOXgr/s3WFJAyU+BoR
uq6XWNoeTSzJR/EYtErnV/rkYt7BH69IFi/whgp5IRncPX7g+Yf2OruGaTKrbwAR
dKewKlAuzsSFBAxHqSI/R0rffT8sxKQr9NtRjMxJX1BLbrVg7af2b+CPwuojeaFG
3wlhDnZaxmRu1RJr4ORbSHOBl53++wxKsL3atWw+T/GiQGaHsv6BhudahZXXSsoK
QNbszCVttZ9a0Q0FlR9pUUKflabb2IdHzHBx52QmBnZEK3Ol2co+YXxQ2NUENWm9
YIbLGd7s6IYHRaGca7UezmFCh2AxM0IJ/BVBbpcmgYrCDRwxXDwtg8gMkPDC+BEd
91nlvlvDcfMycYjByoI+j8RwXxEN2dybkwU/3GJvDi771yhnhp7yBGg/x5MJ9Gdp
qgj/Zk2D3meVM55H1fjxxDeElTXuRgnK0NR3GzP1x0YkRaF743I7JPMuxjl1tkUa
TSMQO6IdeVVKmO0qV9UVFMWy8EOH0UDibL+plPFZSK3xRqzxqhT4Jn0gvaVR7fc6
u5RNNR4PYgrPVDffODYEBsqsFwUknPArAmF8T/LcAmD7+bPpwb0LQFG3O1HwR3B9
HlmW9PeJ/Sf7zwvScncvDDt5uzCw5Gz45IJKXV2GEnysAeIQbMdP1lKGARzN62BE
e0FKgrZy+Vq5Cjv2EF+FzRmSWn/GPfaMT80vMaRk0WxiXIcI8siTR+0ffm1pfigf
OR3FLCPK0gXJxpItJFh61Zp68OyHsBTV8I/Bc62spc1fCu+GcfHp+yFagA9wQViJ
LX5657EFncf3C8MosScPKQ4Zv5qDOzGLfNPN7I/Or6Px4lBGyoBYq1bDBjkDG/ZD
mZTbaa0bjabo7gZF3rzlDXcTekj+sSg+hg+kupF1SVE5MhslSDO62DSxvfUUPuOS
ovZA8XJtJzjGEgs567GwsK6m7aW+0tJf8QJMkCAvYgrhvwfTHMwA9Qcz/3i7Tgpy
ztMPbtf90GLAEKtzuhsUybUKXgP/joUbLjnXUsnu4SzLoRrYsCYa2thkirEOooJY
mlFrBBXEApSqJ6mMcEbnhN54EPEMl0tLxm7mujQ6B9efzD1ttr2rIxfn4bWvfGIT
ZffAycorqYz1Wi9ER4wdnSscM0Zu7glG/GTVSWIG3yXpFgd/O+FFZuFBNYdvIWcW
2fYHRIk9cevpweutOJ4v/nNgKQsFi6EGSklSKRV3cFJalp714ww9+DlIJurCB4ai
puS8SQGyVdAkkalC2JR7EB2Rir7KOOr95TXgdgbjoTGpd6NpbRM5kWggkewylR6k
6pnirKXTiNsqNVCzQuNfBaRWjTNVKiXTULvDGsZFPP4XsHFTTHwgBgKWkIjfnxCd
reCrSAjXVDQXuK0VHzrXofVtDOuXuW46ciqQYnZzMZw+iqcd2qryyfY/2+Y2vetE
MT7hYT8co6lqa7geUhBQH5XkIJUsY2hbkY0tlZsFy5n4vnVCH7k/D4OvZkNEMvKF
4MiRsKCvcrsZpP7utFBTnMoh2CJSxIgffOwGOyMVE3Yv752Pgblm9Anoyo0bkfCq
G6ZfKDaFqvKxakRCUYCXJMEVoCXa6dX111ChKAezi3ZtoAwOipwyQoPqzYhypdyB
qRNsjKdlt8XD9915sGyD+lVudV5/XyqUDQtrgJP7TTGPlTbNf33rv3lc0gRw69b6
awaYLi7/6TXCoOeP16FBKVgVfjNhatleSvAchu3KFl7Uvg4IzedLBnVUztnW/2oP
685Aa3uD/DioirdqC+Mregtq8pcJax+51VCzt4/Ofv9IdPcCM5+FEHUzfjBdx/fJ
ZjtBd0bhdNgIpkld7M8Cx7XoLLULjWIPXf8hmHmq/viHB8nOXPFaRdsg2GNI0N0c
c1FFEdRBdymnQTK53REHjnww5vFFviJAV1RQhti7piYn/TrZCDdUk4f2e6BRDTI6
Vl6ByEW8VsbsUmuYd/IouC890UMKTvQHR6qGuwIh386o3Lvn7ULGj06dlDUm67VC
39vLx3xOjeIh0R4WONoSTIaCqg15S9YjqciKnZnpHeYQIee/OPH5kPBoI7Q1C9pA
FUrpAzxawWAIbGxA8kqtGT0elKcqavEzwOvSYfm+IH5iaYf1JOhY/gMGWNm7ZAlb
CTH3gbR1xTQTBPpj1EjMmTUGIZSKYcj3ncX+UEv83uw85m0GoTXvknWFqfIt1h3M
hDS50AHnWMiBHSuslwQPtd7g2F63CKxeq7xWQVKVqfj748QNPVsdZpnCpxPsqr/E
U9Q2UMFsJQNgQ/GEbZLTOh2aHQWj27Nd7xIZsjlWsJbvZdj1vwuelxThUJkSgSZZ
Y+SXklGtB3m2SLiEujLPO8SeZFhSqaYEROXJJmVtXiqGCYAlRJfc5Jp3RDMzCocz
PBFk+/3NAAeTHB2zDIJxW1vXi6MGozkurtOQNXVD0hM+wu1PiY/lUdZwRrs0tC6P
f7zJoleZ5GBUQgJ7nGdyds0fPGYFUi1Rf72QZimaSKccHRiXWH5fQwTxCO40cHX3
487vD9n3aYPa5m9aPnbyxL583Tam+BL4P43CV/2mhTGmf/E/xylzD9Gop9UONUks
ptoMkl4Oh0NOkIFc0PDZgPcWzYQGq5m1AAUBmd0kfPzCTQdoyRn1+SVq46eDpAjZ
Oi+UZbdVmlXM29RmYC1lXy3KWTKkQJyDMj2ZBQVJ7WH0RlUzGjKDYUAx93KvNkkC
w4RgCGxFmerOR8WhqjVJcoBaq+y44oeJ4vIJjCoTH+IjpeFIGWrrpjsT/C57S2Bw
vwW9Gsxqd5DgCnE8KV66HoR+8VkHNCW6YeVZHtM3vF0cqeYAIrHnFFpjOBthwQl3
ibYE2bRPT9ThGRhrCPaztpHtsVdrXkiYtCa8GJN/TSeFmdDW6SrdqoFP9+dl3zIl
DtFKFShqURQb/KeaT73n4HWhpHWyZWOlX3Xp1NPl0Tr7OwlM3/bYEO6iQOVL+nz9
INTDeKM8AVEiSopXI84eb9wU2yI3QUaccfX2/FfvocLHGW94Dx+cMpY5JrV2MO+K
meUPYVQydVhReRSvO2vswmIi/PIKkiOsdKqo+bxodKLhLZ7haXOCh8mPTrxAiP3Y
FprMaGsGoMatbj4F887aP/gocewsMuDNKspKBkhqgwrun0LDEMQcv61lG1atZBJ2
HZS61tLh65YzJridmvbiwTPRi1vbtkOgwn++QUtSloDoXWfPao0VCKjdrYugPRtS
ZD8rRzb+AN4Nc8bBZ74U29bcK+Hp1UiMNKwuUYSAxwXbLy1K+D8RAPlnaLhcn0no
J9eo3LST6v4yL7YQC7u9QJ0gVE8lOpezKKgVV+2b5V1QtB5Y1FXBJUMTNvYkZi9w
zQ6XhsblxZJzw0SBSgKVL/5A4iMeUGOpSS/P3v5nzOa0AZkRT3TzzVohnwmA2c2h
jyNwPbdusoSz+BISaQfY261VhHcJnSzbJLKxVwfZH4TTXCCqSYqrOxzXvCJllR1z
pBCmDxUhZRj3xCJtJsY/sBAnPujRGwje1usiZbQHoiULVlPMyQ3LROGO2HsHlwsC
XzYR9CqkxJQAKn5BFPWSPZ1WXWRWQeWKtPq9h+tx8ULYiIN1X/1XCdKJKLZaVgJ5
fRjI/cUXnZp80sp2AipWUwc907tkjgJtpP+wST2XQ8PXyd8Osgx4oZvgaj4vVjpC
8dx+zSZqVJlBfLpvbdpjxVag1pv8JSabSIqfr3TwOEdd/pa3uOJZneRITevVRO3R
Y5O3T1Bwk3iE73GTX7ojZsCnYB8heD2AbIX+7x5LuoROXwztyhxCeUIHARIYtfbi
0jyOmUUz3XngO8ei3FpaPeCneVKJQRJ6o6w3XHo7QSqTwkFMYRzW9MuGKrikW+Ho
RuAuxepGO3XSAuquYZqKSvQPgYtzPfKYqaLTFLEiSldBKOEKXDQoPmONfRUvy56a
a7UsBMO3bcpgaBMONKpj1HvGFJCU6yhT/X5i3l83sIkpcBVIv7MgpV8PLnVp18pf
lVKhIZ+yXY6DpOYUIq5Cd169vXBinvJz1WytFYaOX8aLAB3k89NSSDsis7F9f19e
JW2klqOq7RmWrT4L+nz8qF0BZMSJcY0G5rB8qJsFS2WFYxQLA5klNyTNh76AQIS9
OiKP5ZfzcrrQlz+vGi8c5WT51RF1WfhJKDHpmDUlZooZTWWYZVdhGH4NUK5GfOIM
tCc5aby661jEvmS04yUHFjncF42VzkCld6ZJ9YAAKIBBtXTnQ5h5MQ+IgSzMqHv3
E8QwvSDtX5F30/C9u9IuhEGFaUChwsYRXkDRwxuf5zPP6VefwcvB3iDN618TTIVY
MB/Vmo7gvktaUx6eFhjVFVSHJMhd1lxVB/wb2uVmu+KJAraIAAAEVvtV/ing7+iV
c7ds/D/g7qdX54JrQr7Vv62ne599jMy1u+y+jqKAG25NHcmV+/AEvvCQS4G9eY+P
YsMllxjYVc6HHa9e57Lj0e9SR59uC1CNWdRBmboECsd+KQH0htudQ8efOwapj1Wi
nKxrAJGy7eKTMr+Tagx/XkpBPFB+0A5UiWEIaCuiwTyzdEy0r9Oe77zy6Pk+D94s
Q6MxNIeq2YRaf35Njh/vcQmhEGHSmUzjF3Srvk5ViyYHClThU78qMk2YOJFy73OD
psXh15+6xQivtmm1q6WqgBdDahHAjv3DSQVkxj26B/GUOxKSgSC/syv5OSUAj+mO
H2kJFujiwnEce9l0Qe4AxhKcYDO9aMW25RaY5ViBTWiZ3dxM6Vvh7RQNdbTI92sg
NSjl9nBCpg/LljTlMnTSSrX+oUFCp2/JihucOZKUIbh+zvk8CINsYnZwGtSROZrV
2husA59zJOo7vHSUfLIjeyOh+f6VXhH6rK94aA9zmcq+g3JnTO5Vtd+iXWi0Q1Da
8HnbhWUSbRw9vgRhIsh3DwMQyefkRiRDnsxS2YSnjkqgOWfAncHv5EL9uKUtUNAT
stPdmAxpBiNZKXthDNmU/+t9iRsgrHqFeqGV3Nn+WV5kgxSFzXfFxYGS6zdZsGpr
qp9GTKNRbLro7wPT1p3v2HMEkW4fXPFY3lBUo4dDnS0fgoUbl0cYjYf+xjIgafhH
oHSeSDvGq2De+NOq5fF6XFdpNK5EjOin7+ugDcd69cyOaTqrStro25MH/V6ebDzC
PFloS7Trqta9DXC/98GsjsvyllX9xEYmTPmiAZIXNQHC3eolp4x+NqHmvmV78Fwq
uLU4+XDgdbxVlZJRT7iVUiitvUKM0xggmM4sjZHROxh7Co+uZTMCQpmu5ykGIjtw
lrWMPn/0BHRmyCjX28UGhH7XKyDBqjazNlKt3Ek/n4yYXQie1QEMn0T0QXRU3hcy
D0vTsOIWHrMIvt58YvGWukq7VA5qZm0CupmPiZ1Mr0+xWVA/9TdzP8dD2SUtg/N0
RSmuJO2c6gYo4I7av/iNHwMfN4U3hbVymezBdMtGWrmEYAZqRDbVP0htrJRMmbnl
No4zesAbL2t13jjGubLYz02loZo0A5srIPDowpVcpmDONFjC7LLy24jULcOb2uE2
nDYvSNL6r1PCnBFRQB4tY5RWGi98Oh8nUH4qfSl00ORXncZUNyUC59wsNy7xnELH
fIFNAusn8VodV0DIb12pGJu62da9r8LAzbQmJKWn12zc6X1AIOqQFQay0xz0L1gX
zd+KLw/hqmTfgZxb2L1zjTlql3PdUdHLJp83W5uatFcnlFCZvr1n3uY/HjspGVoY
pHDOZfo0aBPlr1/Fxh60CExxMX1qRrPw95eRCzdH5qv4U19EgU4G3lqxKExWb+Ga
u1NrPMi0k8w8rGLQktFCfg+isTxeh48Csqgx4PPQYdfxas4rZJL4mxW7msBQVBCJ
Mcd47fkTpOnx2XUXSswb/U1Mc8HfsUn2jn59H8lakAMXvXUII+/YDmlhBfhZH++0
1cmi67SQ5sHqekSOW2/m1mzhrE9BCfs80tuJCb/Zv4OmY+tFigslt0jho6mefYMU
OLZtgPwOgELZOgGGJaHIo03i+8tLQzK/dmUoTczDplwsTVFtVk61WoodymhoiECI
YxRCxl6nuFMYgKnE/j3XXHlWrv9OSHyjVtJApDr6PN2GW6Kzf59wXqEWnfGwd5+t
oNPVoEjDZ73VfYWZi6AdXP3it4uwJ0L7eBftjP4NmmS+cTx6nQM1m/sLJDyDhSPh
sQYonOoLgO7CsgAXsv1V+w/FiWf/9bIUBmDH/6eLX1Lkc4murncTO1N1He6zkc6R
zHXomYy5ziHXdqGiila+q95VOzEA7N11PCsqlOlszvAIGdwKl7dNlcLDyuYrJiql
dhmqAuQqS1MdYCY/asmZwANsf37czIUVzYdWJ3ozUZywibOR5dt1fITYHFpazIdU
ETVilkB1jlj15PRQkveV0tNSTGVTZz7cFmHaBhBi0OP1d3KWr0CVXW4c2/jtw7Db
AhB+4EjHHErfes8GF51Q5LFRySLrYaEMUPvft6w11D2OHj82Yaac1+R+nebmXte6
JEHYApGrSrrawdhD6iKINmX6T9w6kHQmGBwdp/zJOroYcFL/FP8EwQ+m1Nzwu/cQ
fBNrCf4R9mUQZXQEwgltN2xJnwYQAhj3tEzVqFmNa8f8LxquP6trpTw3gvShq0LS
V0AtRlKH1b/zn0ABC+tSlKV60rLUA9kx2ZOeyLRwa4ICTw8626J+rZCs2r8hMZyZ
81kmEetTuPY7JGpuIZ2uILMThjOA+EjydLhIcT33OgSLRohAsa/M6NajdjPb5v0g
qxbe+XhfMtYVBGCsaruiDI52zMR1rpI1XXG6JjYZnHZpD3k6mRfTHjQTpHOBnh/x
RfgSTdt2xP9fyXjWr0zb8OYFfPfaEtdlvK7vzShnoYlKQGEiLMn6ltxdiMhmY2ch
qSx8ouAmCMRWo4C0ps4US2NLJRqmYU4B6bAZxHEoyRisGbrhwabSEmIkoMKU3AN1
r1vAaPqtwIJtFTOF+oD3Sz9sq8yUHKlsExgxnzXrSeeptaoH8Qc9kyjqskDojsgd
RpkXdPhI/Buz54MiFX729XDLDXDHktCRth2W5uF2+kZ/fwKaWVgTXjxDROejAREM
1gZeKpJKGuLf4AwI9A/iYy4O9t6qLobnADINhK3NKNV8nr5j2aFbo1DYZRV29ZJn
oLz5knnDUT61fJi0kRXRCui2Vn9wa+mtYHBR13auOSVfMEkZLp4nbYvvV8YzepZ2
GizyG4Fr9yDAmQ0tFp1WqujxUcEpWZ7TNd7vC5wjAfOZvLmysHd0VJh2K22gsKag
7y1Z4+7PTx1wOGA0+NlrPOZlmjCLFGXCIKtBEzE8r29rkZPxg48BCWF6FmCXhGNX
2qqjfY51akwt/7EKUcdKOrayzbHxXU7hzvfeRUiiYLkIJHDSZG+wniAQfcLVN7Da
HJHaNHReHmATPLY6L2iP7n3TVzrG/P+4ojFv3acge3/DZJt1wzAt9sR8mBUo1CHS
8WD57vFk6hjpfVNi5PAfAL/0wjozRiseWt5C26dh7YgaI2w14n7oHzAfx37xRpCR
ZNW1JONL3X+WZAeuMDNV7Dc4ogYmgXMxHqt2SwjlPYD8qvqnkGvQ1ejXK9sJpGum
LRLrOTpzxknLqG7xumjw1MrOPZF4FAUWVHATpXsqhBlgS+vRFJS666JCiwibtt5L
F9PEmZ6YslVleSDxjtAif9x8EUVPX3yUVnh/6Kd4AMTpVQeoFI32RpaWXC1Eg8So
C9jppLqK+dPmCbGmMpZl76szmuO0OqcuWC1rglAsrkz1b7+P2CFOdjNotLFGv+ZY
yKc1sIWYGTdliaxRHtEwe28QfNvXSxRQckd3gJ2LfxvaT9drQeK6/qZY7ASXdZTb
ij4RxqgnJMrc73U/mPOg8yfLm7jnu7AZIf7bVM5OVsSR8OXzphWYNpb15WNEJ3UG
tW8VBUiAs9MAUa1SanT8r43ud0CNXX4HOSKavZyJyS0xY0exgPSJn058ZFsCEX8m
syvJVSBQN80t8q7Su2P1tjcf3JIe8+E3pRjIVUedc5V6QVNAFQJAYYK6zZqunTKb
c/i52KGVooBkLSZelgR2pSr0CeipAGkFWDen8iFUc8PP+ySHxMqdJ58L2Iq1GXEq
h45v94wRW0NT/aQ5D/C7Vcx8oH+QlPChFYSpBb7kq48S8ChhpKRYp/GTD2SvjS3d
XWiNCiLN0NF2zGtqjwNo6tScGasIeEBk4ydVXEtVhzVyEz0Tn45CUjYgG2tR/S8L
QM10T+lWQkBr3IXWdElpM1/rAMKooysn4KLMZl8BH3nxAEMEkbIRjejT0v7PksJM
o+MWkwcinwkLkoln0GjFC3Dl0Lt3vfeMjoMYMgDeXFZ9IbuXBJv2WKpJPCXYQNnc
IfDxEWj7RLnhQ7wS4D6pNFB00Y1dcHqaSjOPValC9/2HZPQYJ6/wRx6AcOcF6/Tc
3zbRHZ/yWX/386V5aX5wQG6RZi8qTDsAtyi/VH6P90rF6ShYOyzAXwWP5DQMm37x
tJK2TUSRGtVvAAOmTmvC3QS2EhnPBK/jzWVUNvRv2H+lDJnU1N7dJ+m4iXgp1IP6
tKhvhvboGtiM4/14blASdvMEnAg4Y78pfBNhxVL/aLGWWgCTdESHGotIEJD3CuyW
uGBs+ntV4zEEp9NoQ/C4phPlbrnGBGqDXBIu/19fmsb9iX5s+JL8VPaAYsdAkGgI
Foe7ycP6J9BJ4/8NnKpVyDIHkcS/LG1ofPnkH92B45kCvawmivRl1pl0fzFuwrDu
gzTl11KtXyX5CCiVrlHfAE8BVWyGGLMgfjooHz8P9o9/clUeRvyiWio8ayhpfeAl
hOn+vNQKH9giW/ifkznThxs5WvfZu/1iVNbMr3H5+qpqlNXBsrjqMWkjKwBcAptX
0+tqkb0DrSmGQ5bKSyYMrBxqRmtNw4lla66uRMN7rdMk3uPDUU007cUdSMYZIeb6
xiuDirkiQ1lhvWLT5bGD340Lt4giHZtZTwR27dORbcDCRGW7Om4+I815d3e4tpu3
91G+qSapdMLvHlOLHdLtGBMR7fWr1d7DrjzaBHpf8K4v7ZwjLXL83DLschRlErw5
wzhYp4UvGzmiaVLZUey55sKYf9nCZkVX1OZIhiz8Zi7ulsHQF2KuEqi7maZVdOfA
DA7o6ThcgrXa8hTLzVAhlwcj3PNiAm31yAc23RsAk1VrbVil142kYSBzI5sBcyN9
PsSp8vUs1jW4pm55zQt9tyfmYLO4oGsN9QZWNgKPsFIPsxHE7OeuTUXyOJfq9n+Z
0KLmjIPCKmEzAKjruMZwKG2qz6k/MHctrGs3L+6Xd97CncNlNI1gSOh93GO4qGCk
ArJ7l4CzNTN6nDAy/+k8/kIuuRyd7+YIpMqVOQufyZAb02csU41RZZN+jU/OwCQL
MPocHAfbpNay817p6bpJEpIR9AvBo8vWr7nVPLwzxPutuIP1shH8cEVOzuaFGWqC
ifW8Jhbt1S49sijGBmKL9SzCsGo8CmQ0kIJ3KWDb6Pobi9VLp/LfkYNr+4VG7HRM
Wi0Eb1XvbF6bA5mh6TjK1EcecJWlqRvyvvRSWiEufqid0lOON4L1ylIkD/n9Bp8R
AjtagFSRp7hPC5CpqORdNFtWC2Y8O5/maGLpLFZUstyhhYaDeO8ZX7/sHK5unLGO
7fk7Ro28sLfOUmrl1gAc244TTyCbsfpDc2XZt0dr2JhWn7TFaYADad2yQ43p+jFL
MEukpUGFionoEuK1N7ymK8Fw9Al+ihx7Qc99//VnwuK8HbJrQK7bCyEqHzEgQ3c7
+jEAkigBrci1H3et4c9tsPvGq4beeVBgmBQbw9U9QtvcYytzdEmhaMth0c12bg00
cFaOIhye4AB5//tf4dM/nzdONowN3utr7SODhPvUfHTcLmRLUWZrgbzrrClWwHLv
9+wYDWK6Yf1Jdxay30HX43zUz0dIh4fOYHmzPOPaz3Yd8DNtk+fgAR0UMbSgW22R
u8tBxw0SjEYu2LzL73BJNItHxgQhAhCUcxfFaIUMkzOMAwCPtYsc2Ix2hx/MKN/8
MB7Zf5uPDeJm576qRv15SKpYVIfFiKamIN8eINzTu5mDumktcjZR3YtqROLvivJZ
qDDJU4JL5AInKOpLJsJMz16rzD0AaN8bZHtrdCIRbY3xb0x202vht5qBv3sXw+3K
e7zmAjJoqQvwbA3704G/EEJkxDF25+//aA5QZu820IKIQRKOA7BigPKTsRZD53lZ
schwqpPTTVT2CzSXQgHzQV0hZgvJjeHsrCSTU312W/9FMQ12FCjB0jMw0iU254lP
O9kILyZlzp2y2syV3rj3Sb1pExANq+ZsEIZqA35iV08+0rvDNtolJymv9yxf5g9C
ZpO/Ag9mY8QKD49zBlYCWkgHJIUS2XWcCKCVym2UfYT3ADSF2uq12Nafb9kLwsAC
pSI3K/6u+d7+fgxk5/d/5uDqwguBjr4bEJTXJJZygxL/DEkpb7897nJYZ+tUAWsm
uzlStgNT9C0wPgE4mbM8noW0MyfqlZxlRobL7BDfO7/dw0WMFwdQz6jvcC8FTwHn
ISOXJEZP6cJuey4Lts8Dd2FjiePqczP3GjsbotyX9wBfozxlp+RCAeqD0sGPlM3E
WtKoscdv/YUpRWBaL0UK6mv9cRgYxdy9QEMzIvXUnz68oA25QgcgBEeoQacZ/Fuc
HeFukJMQgp15otbZIlEm58DIsSj9GkI2o/k5YMoZA/mdcUz84ht0vzMvFtfWYk6z
78Mk/BPqhnEDp5An11N3hrp3uf5Od4chyBpQo4TGkSQYzTN2BA8e1N7ZNuIQXJnV
EIXgZdsrRkyILDi/g/Z3hr0FOk7Nm/v8IqtTAr/6Wq3vK2anY4r+kN6qFi5JMlKM
Mw2KnlDQ/FJGPRfFkKTbjXY7U/U/VhGl/ccSkpkDYTNIiah5Keq3iAl1s1ForIvM
34nplwqIhMOexHKgKPX5TsFLswAVNoz4ZH5ODzwJyVeYc0HewlOszPYba7+XDHCo
c9+D/tvBidlZQeAa3hapAfB5mHAuqPkZbcSajwwFzVaeWIUcVZYybHJt/xtQk4pk
/9ym5KX/ELFC91e2eo6SJcQpRpuVMSoAv8A3qZr8fjFksbaG1T5+Yl4lTbdvMuh5
lRxdRr14fOTwaQSGRWsTfB5Wr24QdNBLIwFb5ZLttGs6O6o0Q2uia8oOVh1IrWc5
Z55xFYBTea7dNVTdSNyGvtG/DAG0jKXr3ugNCF4XxF1JjF6qwnXEEdILhNmAUrmL
giMhy2H6tcinsRfRzeDXSFok6VWMKxjiOJTbLpz/Gk3SLd72++y/2josiQa7DMvp
mvCeYj6EhG6JOZPc42gZcSXKO3g6Yvv0fdNwvkG4CvQr8guG8zJIcR2VpqVZG1aP
C7bx0R4LzUwmEFIvYpwpAipXPzTOPeN3e1//8JITCb/WI1664gvex0yQ0Rut9yuZ
PK0QvA2N4588T5MhQLhSP2u7dKl6ueB7uHY/9EM/1peM/IdvDNgzjPVKt1cltlMa
GANPWQAcNP61wvawsjV+eXKSTTnFDGazmUpzIcwbGbT34PT+xn8vyN++GpHhaWpZ
ekUZ5tT9zixd+HVwMqFt+rCu65PBq1R1f9O6x5VoXVGg1m13aSlpP/tOOhKbLuiQ
2UJEwwdHvFhTXQtl5y0G9wRjHvSol1Zm8uhp3w3dbizZms0aTnK+KwDzkHTDUx/A
nzE51W2It3umNHXHFK5N2aa7PjGAdRfNRwNRQCMC0jdH41uFjRh1zkX/X8kxPCJe
g6eW0lOOrBHY7MFCUgcLB+wJT1mBP9iMEF0a7wDN9Q7vvvkOzJdH/3KktWFG0mcK
FXIED173i0QZU1HE6Hdg6ve647ZFYUWJRqoMuK2y1u78ogZgWJ6RfN8BUtnG7G5v
uDCNxLjyX/XpNjGEi64kJpwKto4I8jOmBIsI/1M/KA1TnXpPjfDQFhKGzPFZhnYc
4LZkOsKpXaKc78r2xwfHNaOIsmgmbzHeKBXLB4Zb2Ln7NY/bMTF1qlILDAqAbwPO
6ehHiAhCDR2efHOPD6nI8nzZZJBU8qyzvNa8nXYnDq9VBlnZ4BpbVnr9cWEq+Dnq
VynSrniD9sZYjGXvfVwC65wTKC+pyMgMPT9NFEPN7Dvzfakv1u+DVfwiDUxk+pGp
IhkemEzRwvBlgneltXEaxkwjb41YLfAu+nER90Pn6pxJFqlEWwuZP0LyOXeNcncv
gCRz5JWFaxfyFVB54OsS1cSPYPze8jLf/ms4s4QnM1vBO9tRNZOohxn3iMin2SZm
35eK7OMHoFyJjfKskbU1Vhe1xqlEeDEKIQqnf+S+UhROqDmt/U2CtKa2ALeTgDDk
umW2udOQCDql7YNCpThd184b0++P5AF+GOr5y23G6oDKyk2JNg3qcYn5A5D0iX1Y
Mquv027XDVzwA+hNaGaD6Ixqn6U5GPlv83Z8y2wwjyuWDdXTWT9ozWKpiCeRXtFM
73RYwU6IKvcnxffkZVXpTGtxsyao/OQApYnTqEiLsy6Hn/jJH8v52W6xDwnfMU69
UAtNA8QIkCrOw3IACFHeRXzhljaOBNXY/85m4OUNATq5suHMh+bKiGvTrcwS9SXM
yGvIxrhRzLXx+rMqR28EdjDO64k16uO2uTy63fHgvb5529HguN/iBN4aQ9pnQvtB
HtRtK3W1hIYdfHVdI6dJd8QwSqR6FQcQjtach7mjgkSjkKUskvn8tt1SkuZbM5W1
gJyXN1CaR9DLN55hAHL7j+5r5RVxUvyr5ADrrhMsb1W8lcDYXAM9IxSLKhe7KtfN
Nf5lFYQmWGiCbY2RvqZ0QasrU8y65CF+YftslGyAnmDDz/1SeUU0JTSM9KD/3iK3
F+6UY0kxos8o0C52Gj0ZU1uiyHwihTd0AH9W7StGsM+5MSfCumSD5kZALkyCGvNs
FDYeFtN2se2hdDxz5OtFXLqcC2z1x/lDBpvck86gfFbfoLvhUjLZPLqeY1p2Iy41
iYdnPC9RJ5aEsHINSydC+2XAKXUW2OTLEgny6XSe1Y2xDVk7o7tyXkCrsOoH3rJY
KC7fOoWHl9ddUtIvsGEGPsmujFCpah9VVy4AkuWVXNfmqnfgSh+7VYyAeEbvhFMM
HaAlhbGv9e/G4oaRqmYPlCy5dMyKGIzIYPuH7JQmPZCtfGI8fgAf4aBPlHS0cJY7
JlpH0PraOR7he4UEIQMVHkGm/XObcB7jhJb11CSgmnFpgLez6Lp5ECAz6JcEAHDz
PkkEC2PDeemaPprvLDJrT09SxzBbTwwOTPpIPNrXS5gv1xOFrHSFUK2o2EuSAyKO
lqhjPl7vX2DPTBd04u1n4/lqSJo/W+mYYBa+Nnc3280ujKXeMz3w18z7G3yf4d4L
MJPVrFQLmLDz9a/IfOLX5togyGGpxv6r9BB2Qu0G0lrkpWq5kGVN2Obpg2SuDNy2
XA429VkQFPvlwDsDgQWFhWJn6zImkO0ueb2zfbWlaGtBZOCeBuXI2s8DVvEoDRt6
y6nUmo2KdL3a4b/StGhGTSM80R+oSfF79zHVGsblIrNeoaW1x15jbhF15iJMPqUf
4dik4xKDsj9zDqFoS6r0v1ouCO21p1WsMwoEExoemv33a2HEK7xY9+rjdrIOEFNd
9n7+NwWl1KVLWdc7v3uJSbX7H48BJYAdyk9bO3UlvwmfDuBO4mpK/GgZV8JdgRGN
2uOUdN5m9T9YIAU6U+S4dw2OgvdaCmyBC2nUlZPIz0nQFmtyG8YUlORcZwy+Fp07
I7CSxyO9QLRkHer6RTeJ22DVevrUggAwJgPDIePtp7DepR+tZEcpjJ2Ll6almtN2
05lmLXcOqHMeortNaJc7q9bcF4/lQ2TrPhvigWef6w40+uTnDOh131uYKDfguRF4
EOOkRGwiXJSf94mQIt7UFxO9+lzEcXEo+VNwQWzS89cR/y4T6GbvafK26jvoGJ1/
htpXjWF+5e+U88Kkz17AuBKO4TehHNZ9wOufXboMt1TZNzR6juCEs9bs7pcXRPdE
f43fxZDnyoUi9bw8STdxc5QUfzgpxSBu+j7FLcpQ7ud1+5GSSZQy9R87pN5nQlx/
51baUpzLOkTVWd8cmiTuhTy7Pn+rSzGXu7yfTxFQBSPsF9hYkU+0jy33HkcJGE5H
7KOsheIS7ucUHEtgRuvTJ0QT0MwU6X3yA3c0Eu1daQoNi9FzS9qRU9PcLNrdaxpl
b8nEUYqg93f7qO+YEyRYgiZILSxrWeRDH0tFBRjVsDxupjQI+7vf3K0npiSw7EUU
8/mpSx3fPjLlxaHpuLfXdldIzCyybJNI2UOI/IZgNXqifctrXGHk6KCVvJX276Tn
hJzuCwoBUbIC2fU4uZ5STnIng83b4fA5h37Ly819bTIX2a/s3LPFcGQUHPV2nOZM
EUn9OaH9pTqEP4wFyD4RxojmioIllTX2fg7pQX9HuOL5Hc8WiA+r44ZF9RjOMITl
IEO+8QMkOEZeVLHizxZyKMOX3NKS4rv9PceItwTpmXRA4xOGMT5xZWyNi7Kt3Zl7
TgMymxJ6eNr7F8bnChDo/yVxZJC0Fj37f8PwPoz4snMp+9Oi058BW9O58lOG9oav
AyODkOmUVpGF3ceXFPhO5X+6Zf0gX4NjpCUyc4PgU57qhhc4NM6ZEwNxyHIl5/bB
TzTYmEz0n6MLrxkqm5cxkKVsbgN0Zcb7eUYFhoh2FhLbLI/s/1M67IdSP1YZW7gW
AalBmUT+s0cvzbMCSbmPGxWh1OepCt7TfGuGIxOzIf04MhVQbCqw0hoggRcI9ys5
nk8krapXYL9PrGvrOrIX4xqMcUe3h+jTvOhvB5F9B9eCxh5s2eTbaDaQrUUJ5SDo
Hq4s9o6TgIE143r0uabDCNa2rg7R95WhQc5IUw1mHz+InXG2CU+AFdVd71R/8Ftf
r8fssTBoj1oWeqFQNPZmM6XFyTV6ktuwCcvQBINiGXkI9i0W6gWc0Q7w8Mav2KHW
k1kXkktnHX7hOsym3ECoDc6pePfQW82R45IVvd6jlyj7+LUlBk0dvP2uBWjRe0L1
HZZ6cs4Shnpp/gLRA1YrwP0iOreS2BhoyWch3a+h1pGLimQDX/6WOsjtnUjXfq5v
W1ibQ0jEvzI22Xcxer4KBNqPixtgCLf2UsUUQWI6GAcNikQWYtE50GDuLpynh9yh
WWjekiBgA/Vn83GSlMeZmYVgGYsKE4tE6kTONXi1rVks68VEv12CFPJf0H5anQpB
rD4R6r8oH47Xx+O/pP72gAjG6CiFaQWcRIaqSxGuvnSOkhAVdv/Jk4O9ELWe/RZs
edMj1iMo6mw21PC7iJW6a8FV0/FBG3b8P1cHrWV5DyGooaZNy/VRhaeqHWI93jlL
pVJbcXG2gFxPlkSwFBOdlLOWqmrk/r4F/P9HxYSsa5NGrYbmcNJvHsQGZo/L+Ibe
k7NDqAfDbMGUTOlt59vAd9dPbXFNVXVd2uAIj7u4A4sQISB2Hwvdvx8Gy49NEyaw
Z/kLkpYAt7t8Te8lvde3lWDhJohHFmnukQwv493bIGtFdKyDmaxQmkrOgnv3mZpI
j7Bzlj782O8NOKolhWVrGLUofPSrde34XkZPiri9l2LE0CqM0XFXOfdJWdWb8AnG
XCGjxsAoN1ra33bXxSFBHrkAxsNfB/3Sya5tMzNrVHHCnixVbjHMt4qv/gQ3UJsB
Hm4s9MlkMTL/xAC0DL7gT8p+nI1iMXc5azWXekIlf4COvbc0+m9WQu1CjC0uFJQj
zZeMjEl4m+3xpCesxkyhChD74PRykGLnCgRGYe+6q96Hk4oqD3ADebb8jamyRpgN
q9lmpyPqxieDj9HnVfU9VQ5GuTILen1cYwoX9nUCJTBVkm/LzyrAZrI0dSQXysvU
4fjYHVBM0i1gIl/4Re+AZJaYHjzR07jKoKqvgvAzZ0zsNTOAZPuph+b5s/EwvC2x
t+ErEeAqYtfYhDoQ3kKTGA0ImQ9x14DTMQXQmFXocbQuHxiHEg+IWTfnUaDt0U+5
yRW/q+mFOGDOCI1fkXxSnVOnHZUHixH5Ft3X1AhxOksGsZCnAHSQQo4Rd4zIiEZv
hIC8ElkEkicTsLmr9hn5tCfp2IZYH9uAIQdaQoAWxeW/gAbfkP4tqhHwt20jPxSa
pqnArQkxdiRNr0402aAz0wWYq9CVytu2Ynf+poFxrmQZaTeefYDUQmLr8onSHP4W
hIVTVgPy5HPaHV6M68Z82JL7yVguUK/CLKyRcfOyFnNwpqniElPDh33kHW0dmgub
jTEdecDoIgsOgZWm50wiD+PXetLjEJ8fNpcMPDQfWM/QNUlwi4YYaubtpccai67H
omjK9Dq3DcvIEKl2xCh81ajlK0IkJuZX1OZcqr2cmxj25rHLcmp89FGu73NzlsfL
uMMKJYfBu8gDRNHOJQfuUUtL0/6AqLisrO3L+KjhpcE83wCsDtpgEBM6tqEUHm/2
j/RCJ7Kmb+NlOuPXMQjRwQb+fB++B61769YmLYisQR2hyy2PoS1kJm0UUDWtSZbo
vvih9s+k3lj33YfVdHktItnAXfLvNBt1wfBfvPH6Qc8C5dgmPoDn6t1685v8XxUq
bguGkp267LKZX/UNUjhMn7a32/3joMyHG+MC0scLSqDscRSrgRHXCu47vKj8I2EP
dANubomxNmAbU8DNCJMHvuDba/6IKOssw8fXUCWbrKUt7WJec7aAOLjtBQZSYf+k
JLkGCCaTk9jOYThoSn1ZS4k5QgYK7AQx74PTqhH3qKp5GgYNG7Z5WnV0M/ogB0Dn
ja7PINiBgseioemkXrNKOMvLogONbodomVux7BwTDcDtMn7j6rddq/qUY8oVN8/2
aEtPLnntwKt4Bdr5X9eaQIq7WIY03j3liCbVsCwwTiNRKF6C9nGL39/jK0fHacZR
uRCnBJWc6FiP5tyy+h+L66mXwW7P/cHsAh3TFmlMJCw/5pwqpOBrYYLVr4JqzorN
saLIn+fPJBUwG5fE3jNQizExDxK9AwC0HGsmOMOTNLZlLl4kmxVXBOGkEwHG1052
9rKei1yCoLEiCCLAXiUVCnP/LvAbl4CNbM0OpF1JjeXJQKFP0X8onRcqXwtcGsej
i3K9oHnV6A6NPv3zlwyD3ji/HHYUqeVwJNiEbhBmSxJDAMB281k/hhdYQ6MYAt5p
BwR7fkMF8G7yv5uAi4gNvhFrwxEAJvdmD3znhLBCMZWEfko7ZwAb+8fZz01kRYxY
am75dJsbdaDLhf87vv8edxbbR9NHb7YNtHYD/eQCESFyrAK/NZVeh7YLOGoVSEiQ
q2LfBXwJpKxs5l58Wh+0srYATaPslsm4IvQhYKLuXXr9eJhTS099CYDk7eQW3rHA
ClTEgsPGC6ww+IAH6lN1TQqp3BVQ7HKChlPiNYem+tb4/5roV+kKAg7rTOS8BZLg
m47wLM4qMDYIBwQDSbv29W4ZyBaHaEeQkS8e73DknVzvTK43F/b4Jr9IJ8dlD4Sj
Bc7UhKLV5C5mdcUslC/nwrZuRj7IIQ9zUWctZGFnS7rW5+Xm/t1HKrVLJoczr95t
+4TrgdxOQmdYBqje645wTwdpdeMdJx1NTq+SMCKXBPozSC74I3Cv5f+MGJb8KDLC
hJukCSU0k3P8Wi+eud8vYhItwUYwxpLFORJr7psm4FFNl7KBclICIjVikA9kiT3r
gC8FmUV/GbgxoUaD8NHcZ6xbWWQjE+DzJ+HVnYsZggwG7LOBR8p6JA0s2gpc8vVN
RhYLzhm1fLJiK8Sg/bwgflOxUSp+UGFTikFuhS+ZqE64jLx54S+nVCmZvXhGgv+H
QEzitD0LD9Ix/7JKfB8SvUKMiBVJGPv7t+VaHrgUszbtuPwA8WgbVZv9W4iXyMLl
vGl3jq3u5BK6BTa8gIyi1N1GltNQr4+lpnBJI0b4BbYpPBVqDHswPZWQVOM5x3T5
K3f4LURcBd+7CTQ96rgOhoKGbMfsC0tJD4wsFPczlMmgiZlqjJgX2DCSEP0pu/Rm
zPOJOnYaWWj5pxaYem+chnsEIcMaonzEEoT+ffuOK8ceiCtWZGS3Q4Ky620hLD9/
Kracly8jApyBQgSr6+fYRAHRy3jiM16LUNbEtOdahe4+JTt1SKij5J+2I7tx6wv2
mN1BYdNgV+2OqjlZhaKrXZAHceyqfceAV607wGh6PhZZthIWjxO+YedoigCTLf6C
/SudwGFvqOgklFopReL27NbIaeRmgKkdRzrbVEbza4/woVlcqNEVViJR2fRfJQuo
JZ2qQCIcToptO4pq8pJ5tZKA7GbqQcATsioqQgo1XCIUsdaLmT4v0FHWok4bWcU8
T31M5uYiw59ucYClcc7Hj4/uvUqrlWN0+xplTCGdLlI540BZpm6c7lFN/Sc1lGBL
pn6C/PhbgOtS46bKAP1hUr2cizItbDOlwkO5eNnAt8zEQU1XgHRurBh3ZgmhNFc4
gMwKKdUufq3DUTfiJaUtr6EN2pf8UHJPLqcX2pc8EJglsEBLK2tE4PSzOYjBgqH6
zxVYLj2o5Ytd2+UehehEGOLAohGeg1GS4LssaOKOhw9QcuekhR8WxRl2VsOztl5s
Uhsqk/ZpCX/yvgbqr4QRJ+IKurWudH6q6To4lIYYYeHZ29MwHiv0BjI+MWMzKWsH
SP/kHIny4dYGwm1w3f0o3026oMZM0KbwV3tM+m+VExInCIBqAMfgbayTsssqXSkN
XAxFve2HMF1MrnVwNgFwonDHPmtHwRBPIilOLBlEGpiCn2dG5Ll6aoeLaBECeYzG
fSf/KX7CSRTi7bRzQKf+hUOoCpzbegU0KGnJ3qV+Vn4lYVLe5XMZE85gfHtg5sqR
U5UK1Slne+RlhxYG11BCgsTueAtfO8YOY6pZpTY3HbLei+dNkBFwh0SAPIRYyF6H
gpNfoT/cvjvtIYb+TnfDBOQEhxQ8MMzYypWLu+VvPbc81v2uRLguR/M7MqXVYSzX
NJTTrmi3xOpDS1KW3Rm5Ipu7OLtgSyG4xpEJIJ9To1tT2h1YAqor/EVa2meDpQUC
UMG2oFNKxJKwO5igmx0PBAoPmegrBCI/ZA/Jxy4fec5L8GVrbxf544nuVvxTOqB0
BpEnL/aK/k91XvkyetTGZt1X8Lfe52qgBOhmXV8N/xBRsQpwb5GyUXx3WgHn2EGB
qjf3xL+yWx/CwiltGQPFW+iIy+o8XTscDpWBxyt0wXkJnVRfjC9Pc3WiIbunEqsB
pIIbpZUcs+fjnfpfoJN/Ehva2VRgtYa+WrBsM8iIrZZMYkG0OTk6QOfUjfjHAEdA
zHvf51Yoo2hKMr+QkNm+EPzLoAQVwKNrxvHvPAyxX2MyMAeKx7pcOnNY286vYNgW
OOJPXobVqFDtj6E26uydQ6W9JYhzfaBja+2DNeRpJ1HbzvmMAuSeuQHZ+poOtY4T
WhMofoF2wLhDi7S3ydftnpGJ1Oj+/Dyb037IVLhig66hD7vTUB1+bQzDmgR8n20X
aDunEoUlDUbw20dq7+21bBB+WeyfhIJH22MAQwmAzHhZ6w7rsf7hemP+gZUA5Hn4
9/EktxW8EtwkypBYmSBEkAIC+fiLckr/9kQ4OUDAkLJdf8Oyb+8dzOt+oQuvdzPS
HM7JUb+kp5AtuHW0ZslFcpeh35RytBA33BDwNyT7QPzJBxwyJJI++RsAV2DQrH1C
4l0Orkob6bNHBfVVYugbrZ891jJOQgMlyvRHlY6CQ8Y8PH0zWccBsGGb/QHp5Ipy
MpljDinGaImKziYKX8vd+4tnUHYu2N/N6wUK81OYWNF2o85mEl5lwrqfkE/wD0Z9
t/bQONo5Sfy9hDJ2lrE+IpbomCl/p8ibjqhtHh6/OGEd9LYfk/JJFXCkpt9YmWv+
Wq4Dkxo3OawU4s7dq1LfrGzUsNrabMyz4gm1BQ/WrBWepwqYUlWkT5opTCK3wQJj
YNiRg/79H7jAAuucSoUPzTFQjWAK09XgozumjRiPfpKvwvCdxmugFTX6ZzfqEIhY
H93k+h5xK04tlfetMTkEEZe7qjK42yKyFf3szrA3E5ikmQ3EvQBFKTgy6/ji2JCh
uaInAdb87ldvXns43nUyh0HMstMb+BygQh2YhqQx3+Z3kWLEhc33h93etDWYwzoV
BHb5x3tngjjAnGfpsUGb1nlQQubZkHDMVCZynqJdh0hliRsn29Y7koc39h75uzPO
VD2teZWw/MkhFTt+t6JFHk+xrettZL4jwRFaU2Hl1hqZRb83MJvfO5OfjgO+QxeU
S/0Kq19IEabrh5+X1CFFnFLMNDWvC3PeTTjhwjAghCv5mfnEi1ydJFlUqM5J00I7
hgh+VcEH7Y7x9TjTbzhHHgsRkNiushz6PC/pwuf6g4IiFDDYlzL4FO9dMM8KrP1K
JPYRyLWA3cPfPmuc6WJ/xboXQBXFserA4+xgxLyv/DB3KP3EYGSJqclTecWmn2k/
JdnyV/f+yowWjeDNsc3qmilzSM83nX865BRcBSW6nn0zHIgXLft0fKIBEcOppaly
8r87ebOVB48jJ53MPmIJKajTpQeqLc1tC2q/zVSj6EBzv+OBQBdCBvnAJ/NfDbE5
DvcMqE28kzrSJt+3q4095t7oKTMg/oMuHdb0A5BMSJ9gAYFFNnoKqzo9fUF1A29g
l2HiPGI3HbjART6nI2Q/gaHQoIrb9ydL81kit0NJNSsaTlLQn8eedFOvCxZSoldw
A2roS6XXNWhCTcNAt5HTb6kvLqmyOBfO7sASY9wSFMxjXqQ2p9oZuj6OdH2NG870
+kQvoT8o/HXreLgLtxgQuaQq8uaJIDyQ5EA9spTsW1T33xS8H41dgja6Nye2OPJ7
QZ06N4Xz2KHPHCF8YUOZ427b3YdDxP3KpPPUYj2HumrMzQSFe4UK8ukrV57azzhk
OFJN0lxd1yEuvIywOsjvxqIP7cOegCJt8iS7Kf82Hh4WeJVMhjIc/p4m+olX9uu2
xsWHEder1qDv+xaX3HAXLWzW851xqTNDIB8vrzqQq3mETCwH6v+fmvr5sRB3BBzq
tROJveWbstGVeYF3Vg9CENCwFwp6NHAYv/i45IGVJwelr+26gqy7RWxTS3+74xyF
jTCZ3yBaVOztyg4+8GXXcLGdtGsMhVCRJno4YHpp2AWmtxU4bF/LZ4WWcgus0+IR
jDOyK3p3ngTSzg1F/+qz5ukwm1dwUrLmatUue6xBC5bHYA0aKhIyjngyVapmJ62C
LVjq7O0d3GZLqkvrABmMuvlOtrzCzVxffkT3gmMSq/hg+h0gkD+sSNXZ21VIwl+D
DkMJmgTLRHWbXrMJOn84sGJyuR+T/TNxcy/hGKrUhnAVNxZUBySroogYp5bUc9Ie
fb7lEvl15GhYedXZC0Eki8hM88/O+HHUP+ehcCWG5t+PPA8dW90HLxXl/UZvcsBg
0eAPzu6KxCDhFocujDldDKKYJUbb8kSYLmygFJ+M+PlQAr/92zJD6mNPdqW5lrmQ
cf2WE1LhiNt/qM6tDwbr6I5OnxlQ5SF4bXBvOSBKVH4jv6UR/JYATyO6enfU5kZ7
gd62v+tS3MkpvRHaia49z/kQzeLjR/fcsOU9dgqUwsQV1Jg9jgJb4lwFGpOxStiJ
ciNPpBNnwmPFGr1lLtqpu40d1SQc+YjZxJqjONr3D1U494c1V1Ai8Y6An1IWgweI
bTMO42MV3pCIPqgv/HjFEeOOu95tNw717E37SCBQPssAl6svLxV0bmhh+kAKj9vj
0XujL6lI5LapTUJMLoEHits+F1hyLaCP+9uGFkeSmUfOfNn9MdrxtGW7T8FJvQHg
t3skkE7X4PLiQJChrzfoVSrdkM3KDI9Aqkhv62YI3x1XHuPgdYaf7kFzd8knpX+d
nervjPN11C9vKOT1QXSeGnTtoesTJJ3rC7+xzWBDdc2fI5rfydGn0/Nl3VQ7y90k
6BPXOb6Sn3ZTqgav3hV0hLClU9cdPVqYF4xrDWcu9UFpWMfL7f4zaNO9cm/vhANy
hUPMLNqSlLfp0FUoAxLsPnT+r+WalkFBmjZH3p7wupUlecfm7ZjiNj4Rm3W8m97E
uXfKLx84bxxVzEeKxLMnXcm1kqocGjN3nImt+Rnqk1w63uU84VqzJo9wmXmgFMv7
ecaOLaglb7gI0P2h1JyGaZ7kCCH6vMGC3p2X7OS5L0n6fuELiGBvGh3/m+bpjiYS
SSuZEOleNHUfMLoDSgmN+w97MwcnrayuBX34SBXSxZCVOF9J1Oybusr0R2pLebt0
9USLb/MHbiR7HNkkqHwK9Vzd2LsbH5d5PNJnLb9eMC7NDHV+yEiwnUOJt28vmecH
5Ulh9rIOldk4cBmwB6VydoTlqKdsVpNwyShNG5OEz2DBmikoinnbdiVo/kPxiFZ4
vU0KaQeofstD9okPix5+BA0jNBPqmmqDKoXuzQ7Y9UXPt1a7C+ia2D8h8LUx6ULq
CcnHy5tnoJw2QLVehjNKzcsXCXt5pB7kyCM6uhj1eg1sChRdFsOpHtNUyyc3Algv
jQYuEMF2LFrt6fKCCmwuHo3O1sF+60zlhFSArmYVtiEdJtAk37jIreEX+3kmoczG
PQA5zUg9EYZGQXTQftt2qoffRyZJsNEwtVW96Tp1ACk0S/IHbI/MSOiaLndAVkEz
tVFhy76EYb7vk1Cv/MfV8acDpdWBGciRVpYv4bQjy1S2UVUPCIqHrC1zrsKkhlJl
xm4m4nB/TPt84UmYouDsuqbXv9HGaqUX7BDnpP1hIpDYIf8n388xCGbEb2JVLFWz
lfgvTZAjxI8Cw8ruiiwjOLyHfpUbvX8At2OyNDdtKdrLTHb5RHO/gb/VVBrJXG7i
2B33xWN9fi/Vbznka1UYk/Wc6DSghzc96KEQCqt10IYtHa0bRkSRhqoTWrg2Rtjr
GtPZpfhehf5qy0sOa27Pfu0s8b1gTJp7PJNxwURyavmLra4fjO7urP7JDzU6HrpI
VAvwqY96hO+fgXxeD1ymtMOVTxGNTUrKTf3Ur/vv8n/U60SC5xSq2GnFrZRPk8RE
urPEPBdlPy5r+/usHFTqfs0o7GJDN31I69NZRk2+9v/RiMm887OsA2RqK8Hk2+DT
dZGPARa04RRrWjnDwp26P8IXa+ECC9OepVk2/ScZ77sBQYB/fbvRkpxK+Rjm0PkO
LGsfn6SR8AhL8IDY/kNT20ycnsIkHNsfMZYtwjINW0VnIIyfFtBY+Ju/7RkRcR75
4wM2tBduMb+JOk3SNwAh0w811Fr1RirqlO8BYwSm3hFvLDp3sKAt2QXSz+P8/1pi
E3VVl9tZe0o6pzxIztMDvFf3U/JhaW8KbRkrVTgUwhDjKL3LXI/+DdHRTMXYIq3N
ma8OhIwUakz5sDScAxCWBJiixuDl7hX+qpPTed7lBk9M/gyCv2lpI8NeRAVM0p2I
CG9DVQIe0cWdDpfc6feYi2z2HbrYC2vx/X1uul0tAK+X9CgeN7cWuhk0Beq5hh4C
OUe4uqmrf1X4PSpm5niE99CC/io4PucCQV+h3ad2S8T4cYvOJWjeYObo/bRww7QH
+6KaN/8UGg9rg2tNkKF6Qi5JyM9vus4Ob24GIVrm+e6m1uL3ESHiOVzkvt/KSUn9
WZodgEsLiE/LqssUFFBviZhMTr56GInsc3cxS7rPlKWttyaL43K62cV3/en1pU/X
90e7yxEE2SRniwDxdPk/+f4fIlEBHcXPpV6fFFogccWQmLBycTBH+yFEGSJTg3sm
lRIxwk7WDVI6oswuhHMFMninM3G6dqDtyRQC4DO2lNO+0325lZCJwDKBMbKrfTi1
VRpwQS4GwOG0d9YrPuezzapWvyy3tLKWhlJVPxsVDP7xFl8cN0U75GMrbHvo8+4u
v8UdD1x7bw50bMPfO2SctSxOepPvl/QE0hJ+JAgDOHlYkRwqU1AkDkq0d54GipCs
6SckZO0umi1H35N8KFOLFVIYf0QRJ/ZxMVi39CzvUhHRHSPmZAum6DUQ4i6pNcLP
Gcggn+5tvGd7Gi+fXKWV9NYncYFhXCGyXB4HeBd50J28OPLkVfgqkSHNauFCfQC0
4688LPu2MJgud+TdAaH0LKBZKG+VpPeZ3fVwI2c+SYSo/OPIOOZJbsAPFMN2LO8B
RAmx7gwR9NjPXtsKhbTaGNmnv2d/3ziE+yZPUPGUySnrIR6x9KqTtmosNMX8EM4h
nM4e0VFBvBSpWqG/qfq8U3lVusEwraIapJ1aVb0c3jmakQE681kBCGJsOgddQ1sc
Xek6zIQFnYV5pa2RUJD/tugstyH91lfVGM568bR6SMmi7uelwHE2bYEz1kihnTVo
EMBYT8YhOBliGOqezd2NunDxK2EoXd6FwDNbGN4KcTKQFy8MyLbifu+szuhX+7JD
0kTJvuMYfoUh8tALTG5q1aJHKZJX2OsC+UvFIAf4SsofFX30zwpubBKtl50O0FOU
H+ex3+2N0xHr9rc1Cp8eODGsNCfanuWLzz4GCl/uVzxj+4kvvejS6A8UpAqdqngX
zc4w439L/S4aGSFz5f2x1tqOPwzB5Kc7NszG+D7Xfu3R3FniOYs6oCoCrT7Lyj1f
E0o3kOu3YP0AG8X1ZWqDEfICXlahJB52qU/LOtzh2StdMlHQiTN8PwZeKDcAYAJ1
xi4vEWQ7HA2BEulZiokwaC55A7eR8OsvgBXqc0rfch2xu8DtV9v2z2733b08A04v
L5OT7J0iRXyFMapef9qzF0M0aNxlb/m6v95niQEoiB5o2TiS8d3OY9hsj1hQWmhA
Sfp1xRabg7jKBbkSxQqccHKO8j7FuznpGXUoyu+p3fCET2eAsBFLWsEJxAzqXxjW
yDvCZmm36eZWTbfjt2cAB4k+cHHGse4NmtpudbZctAMZfmsCzJwdor678ssEuWrg
NHGsDm8IlCOXljaI2jetGyioS4xa76Ph8t+AviCHz2xCG7o/45sWr7SdM7p0+HTK
+1j6NqiNRDIGxWNEJ/eYERft8qJ4jlUc/qkfX9UuiSGg0K+NiUcvuV2xSqukAPS5
crxuJmfAn5pFP+0AIUx03UbFyR8RZKujxAHkorHYt/ULWa4CsNL5VoXvmb7rTju0
MQ/3XxTOkiqvJcOFHjeekAnPpDO7W2cIUWo7ljpZQBbCphaYn4fDF9Lwohqp/yac
HaYngZfNhbcj8/kNlqCL/M3EvxBgGIPyG4IzSNbPU2MGklp9F+Fps0VZwzkhQti7
SCU9DAjooqsiZG7Do6udnZJeZwPh+VxZ2dEw1OdToxMxKZPMG9BJ1xm1Wtga0squ
/9XoM6prfDJhAyw5zBLUllMAg1rMYTPLefwXyx9pPAdkodDip1rR5YQV1tPovKOj
vZ5Yd38WDbB+NTkZVq+MhBKeiAk/2DRHF/3mXu0VqlqUg/S2rT9N4sKdkBhbN4ye
VX1hHpbExosKlcC1QklPuFEbKKHLzfMIOHhOUXooTXmRig+W2Huy/Sx4ECNsMWrj
boouvFWeBwjeEsSF+xuufAA0qaWDE9f+FIGP4GIFB5zCcN8W1+zPOw58SSqdgfMG
fSmlhRwkHQehxIKSydvwDQoTqEoZatSEw6NTk9k3JNph2uCTlSIa2wTeqx7cpVDc
e4jj3U3PivzPqXBENojXq4t/WE75yo0CyQl8yzfr5/MBvn2FgaTC+7U2Av/wNqC/
cSN9wHnYE0mtkXAi6mNyJVfEs6VcjZ5KSo4scYYIMJR+4CIL06pr3/h5/0pud9Mm
fU9ucnOWiDCaqew6pLGHY8hbDcqU5G6nEDbIt1j0PczAkIX1k6fGec/hcZVjQmxV
uJozYUh7DZrX3HcbmAbbglYo7gJpybCPcpG9BD4PEPjlf+4S5BIxJEr7fltkLYFn
ss7l3JZGXbDFkoM3QYPPfyldtfj3YtKyHR38dm8Ib4YzKBUon2ulegh3aanpS3MM
V7GHN87Ovsa9RUCBsIWPjRk1KWEpcqkMPhysZtBHyhBpzMu5Hah0FySi3E9+9o71
4hxWCEQVVjIg8k5gmh0gJ1unkmnjVVnXD4C9FlweiVkeLKI20LvhHY0opJIqch+q
dXu3TX0XRMhylby7t6VBGc1UI/EF7fTO0c8c4uX6Nptqa5a/BCZjkIQc1RYc5ZuN
hqvjf3im9A+GW7cc/wkjFkN9zyeVtkM5a3QZ1O46h2b4C+q4reIHMyZtzhjUqRV3
er3kEvkMzFbMQSjbyPfJgvfUJfXVAbRzJHW6YSG7I5E0qIBXf9cJkkwtngQo45I/
9R+q8fqsXpwSSxqn71F+J4I3+pu+4d8IS9TwvNbRR98PMkMOVNCIvCVzijJs36cd
Y4xAO+maeFLy6rbJaosIa+I5jJlgCUq9CVCi0P3x3xeZFQjv3cbnfWcDLetJSR5q
8xEJkBb0yoL0us3/pscRDKO11SLNe28iuFQcW1Hl8qEzY4Ae5ReXfZSPB3vfMT0k
uSlBegCWi/BvKwEZoKsbYliAteNv8peyx6gXg+7alwsYaLHhOcSUs5+/MLX/FyoR
wWci8svixIByActLpVpsD/jaPYskpQpl9/gWJkoofJL3gO3sLHFGdiS6rSkmbB7H
ghPDJQIsDwNahhHfEjv8D+MVhQvg3QjMZEiDG37S7wZY/KiNUff0zaGcjqd4pCZw
5zazNmHzXZCZPTlVjovZPoY3lLJQ3Y7YiBscYGOgcx9zIXnTYnV7EvUqXlAP9zs+
wuN5W+FF8m+TIKzog47dZw544w5YrjD5+21oFqpFw9fdyaDDL/adeLOvxxmztr8a
zyfxGl8+mSCZG2DRR28taC1RA4q9aE7NgsbJa2E6KclUiXJRAXuO37xw/OXFFhM1
Vfql+/esj1qJQJ+rmuCeJ3Nmr2FdKNdCrre1duDcMxwpJKUdaEiZUvpm+U3WaGeV
yZEk0aFgMcvsvLsgyD7EWkycRDEoJifC5LyVrnbP5EoCvVE+OgoUnQCpsrTbS5nw
p+T9pFpIRp6YgxsZVU1YCXdIuw2i5kMEZR80KErsOvonNS3804JBM3QhdEyU2msS
+ha1AZwdLLWEce49f62unsQZIYPwmIQ06rCT6fupX86kEDIUMpaf5Qg+v3gpZPuI
FLzQO+ta3QAwCinl8XG6bxREackRUtoeQQSPnU29rRvW++5YpvZ96/obFtw9H38j
SGnx9SUtOTvbIZkCNcMkn/H617tW+/e7rUgVUtsofiSTTtG8wegJ+ECoNXgpol6d
JwG0mNPBnC/EXonT5+COGCa/+MXuuGdPxezCbFRd8ee/J2SD1rHXIi+ecQ1y8m/U
1aTQVXrMzrOHEoUzJLm31dwJOgC33qYBEZHI7i8QBp1wkjkeWlHfZ+VCgL1ihMbx
aiNSjLYkesYponyjhF3DuT5dFJdRS1bhw/ySqNAkcZ6BMv58hFBrXyvhrD1UL/7r
576rFwqIg/CP+zqpTkd/fvGgd3/3KUlQxjsfk3eL/w1C2pM7zAWk5lXb73Iw/jHT
CaOGkXonBTIIeR/D9ModwGfh8xOJa+3h29z7W3+3LtQlLbtTslYF/M4brRpNfkH0
+UBp3izaFQIeQQs9PrGbY27yuB/P1aegl2nedha0Lro8kaqxxXrVChnybfJeoazQ
VymhtbYmbCy4uZAhFsbe9vEB+7W8EqBaADmnbhK/Ex/q7rwF3kp/OGc0Jsxs9Ju0
4oDdsavmATbthkRsR6AqHJHODJ0NBy3ioC2EehPjAKsnQKhKwePmB6GsaIUk0+C7
qjEevYEyCXeHiso0VlR4mh+/a1nuXr9ktQJqsIN89Og9ikgG/5JFvwVghtfB4nNb
pN+lcIpeo5oCTdcXAEnPf2RfX68kvLW8Jwi7EakBiXvqcS0iAoSmmYjG8Ox4pgLV
+fOvS0+K6Q2YULKyYD+++IkU+wGmXOo+dT1c0nqJ/DhnVpNb8q7tSvGzCxZhUrTM
2kxsERRozHR1LGJPQOSb0jtdoW7r8mWcfa4PIqkqh/xBBcWm1PHpxFal9c98LXNx
E0DBzAb3gi3vIxwMLpcXBFVJhgzkPnDgsRnbUa7bzArsY2I/k+Wq/sRNA469si6X
6bQYUjtS7ZL0U+O1YRQZnwJgMQOgloRpWwuvivhzqnvRNDNcSgD8CP5InPW2W6Fq
C28cuj3yLidHABWVXpvHgPHLGwzHpo5cMBGd8rqChfc+otZHnp+BDQWc4s4pzsgZ
/K7io6kLo+lazlCEDiHWLlPP9NhbTFcXDo9Xt+bhMtRVHRo9EcVjZUTH1FBZH0wv
eP9hGEqbJqGsd0IGl1H0IJr+KtoOWTIc0N1XeouQZNyBsLhju5BHjOQ1piBPKvPO
lxHVZ27hOxRJGZMnl6w9t7+weZ32lXlMRW6uiqXDjolvcKs7Va/O8aSo/k8esPVr
CutUUCUDDmAmdJyyPkPQAvIvG089s76G88iUSiRe52Ku9HKnoaQ/g8PQx8LyYejB
1VMdJQ8EnIQyOJafhTjT821lwUaC9zvvcL/VsicJW+NQl4v96iRE/48yMBzH/mGl
8Jz1Va9fpSBAyc2uTMW+20sQ4VZorxSxo2ApXjzLv+uiN80kDpg9TqXIzXUDXsmQ
dVOaye1RjmRKhNPgJ5FH1CIyyPut2GAPiQHZvKjl+79x90a2Ta7u8Er2aowcPn2O
5XvnLujdMZ2UQXDIckPNn9FlmxlhpSg3kYgvY3auMYtnZZWAJ19e4NWSa02dXwZQ
AW7JF9pOhAKsmfry25zjDQvHydZZoJimgzrz4fXb6zwtMJA3Kw+wnsFMVRdQvNLI
U9XQdTsaFDwR0qY1i+bbHmCmCPPVy4vKfbuWL0HdcQxLDVdVGwQDLp7gSnwXoP6k
Ogm0LeijixjTb4+uDxsJfoIYnQ/mHShf2neEo1Pej1ZAwADs+rNhFJbt5pNrs2ef
4pGgKj1vxaDr29e5TwLkgvs+TZPpzHuCno4AajkiU2WABgjxXzwTVtu9Rzjv2BSI
rqWxkd/j4j9eQ61ghd4fAX0AUx5mMsjAxZ693E9ip0ZeMNa7a1gcZAc0R7yS1hzi
xaOo0AbWuCv8D+76Kr7oCmMVNCwdRa06UR3V9gh5bIC1xFPV7FrZWIs4VtmgcTNP
1nV38LlIIha7+n/Qg75NW0RSY8CdR/fXQgLVSdBuyiZP9ndEXKfE3L86h4N5bLPE
5JqRLYmeZsUb/ork62HFZcLfX+ne0Y4QNxL7IMohGOhtg71b9U3Zno0n+FQzVLq7
P9pH/8K3UIKlaA0qrxotkX2B8+g8wTlZs75XHO2AtSD1lsju8qTXTD+rPl92X7d5
xAWASi7dybMNxbbILIOPaWr4onSb2C5eGFtOuNNHOemGAigjOEJQ9YYe5B0Lprue
qimXaFOHkr3DgObj7yaEQrxlv/O4FFX0Vux/+i/IVnEtRV2JdZoVTYgauSV6mWiE
mxpjLO/CPzJQOeR3kHbfFW430KRLKSEJyOLcKm6RGXM+S8AjQvE6YfpArJuR9RI0
qJ+mTxdj7MdSWpuAli8P/rgv+xCuJCGFNp+uEvaM9zpLDZ+DWbxdrLm2PNKpXH7u
6ZHHk1KxqK3kP3uthXWAQel9Y+qwiVGmUam8Bf8n8w04fzPjrrGja017KTp1QS/+
HWwY8708wlOpJEMrA9EYeYhUmJvKg7zHTOpYVZC+DTXQHE5JjorN+frUB1z8xZOw
+2veQ/G6DNOaohXTf7qvk6GxiI23MS3D//Q7/oM8gyLaM+qd1YdsqM4d8namD4wR
K0F+HRw3iS39fQ1uVcSSVSSY6XDMQ74KE+g3FchjLDwKo3w6ZG8V9SbfKAO11rhH
WRjy7tEkSn/6YbLWK4Jdtw4d3EVKzZ/jpAHjvAoY0phXBzD/VH7s97TCt05phvgd
b9NcfcT5xrSmS3+fijwgg/z0eAw3AwH2tYjByoykM3IUnuacVIBUNQzoKTp9bxnU
/z12IgSgCDxXeR1ji/E/Ssd70oc2o/VEZd09u1nCDa8mTJlnWArJYuYdmRAjRsBM
MBu/8rULmEzkOqUU00MGis735+AMCGeq6SZEHgZHlVBwWVBRX73AOWg1V3QWk/wo
2EskXxPPJKrGl3axA/E51W3CN9vmailGv8MJSgBWwnwKHFGXuv2E6A8U75f+VdFF
9DaDX0a5tl1RjqFtYBKmJ33LWYlriIvB5m3P3Y9u9bNtI4utyGLKXsBB7EslXmBO
KWq0EumoDrKRlD6Xwm10WsYpIJq2EVkaB+k8jGashVfwSLKIT/XyGXnRN8+9NS0l
2AZ1vv+yeljgCTCJWYbBJ1mZsS4aXM0O7ge+4Ego8jF9ZXmm8la5q6pdgFexdp2g
HFcAkZIW2E4Yjkb9MrzH6iVpBZEMNMjEV5WomgSSdNdpXWWef3Re4mBz1OZztrpl
HteL3es4zqc22RkXQ2SKmN8TJ29WbHUebhwgKZa02T/6r0bpghm9dTjaIKl8koQS
r8K4cTWXVR0W2KcO1y3cz9PcyjQ1a9D2ZkOMFomB7/vppQkqASUyIMwa8dJr9Wsb
`protect END_PROTECTED
