`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMVmekwRBL5P0Dbib/7d2z3vhxD3gPEyx7uGBTRQX1Cml3iTtzmHKI5qQJW/weqo
+fNan3CbDSsCuEcNWggiLE50TtxEUvzjH+1P2tgpYb1oii0j2GhD+CeueCxBNyVI
yquBt4sxUIBjRnLjZMh5rRh/8aVSSexCtkBYUZzRRzQS6/9KobnO3nrqtxBkWDmf
rGHlXzfKoV/Q1PtxFqXAEth1c95pxg7nhVNx7mW5imZKzZ6aAUFifModCjzmMGCy
aqPdc2bHinvT0kjz9R2VN0JiDtKKoGqKcejqiJRWvryAQKaDiGKoVXuVHYWv3nsR
dDBs5EM1FgN9O08LtkANyD46CDHUzf7YQ9bxbMJp/gzVDZB7y20EN/4dksAf52Kr
6cukL/WCvYPgIG+juqxx59BsHEfRVLCJJk4lUwxbCaNDMX6Z0kB4u/vjpt4U7Qbx
bnHOMgqHurjDXNZ3tEeQUseRFmN6GsqPoYEeFB8eQVvy7L3g/Wl50Rk4VqHZtpBp
S1FQhTb6soOUlwn4Hr2vM5OmfEeiTzNgE6QKMfkjAxFuOS76SlZrponFK4OVrd6d
Pt0fvlMhGcmWmZcTJ97VLlNyMOgJ6v9nz+y264S9loFS6gBG+gVbCFNvtFLxWO6o
zH/2rm9IcQ86EfkO45/dpWxKaqnlu/rVz9oepdkKfZko7h95gCcypnBbbxGYHlCi
uYI/v3STPAjJtYTrhkjUMFtqJ9EKPn+N/Pms5xdTZHI4zFZ9U0gnfN4iPrEdKUIu
losr4g9o57t7q3V4WQ/n0Hx/DFvAyiVbxATmSHn3bgCqSB0r9Upu2cxjkxm6xpOS
BOaPbXGo3Ti+0ir6qzQ7+nyk7e7ky3bVzA7w/rvCHv3VdvaZ28mb0mt4n/SqywZq
Y5aCQRte3SP52guJWbg7VrNOANyDqQNoDwuPQllQ8w9fmTM8bQfJ9X9ssya5xhXM
zx5wLmyjDIpV05MTZk3Gj/goWSoz7CsDuq/Dkx7eAXIws4ApylJlp/ZhTVUzW+di
uXZ0UjW3HX2bttw7AIP/8jPz5zs9cVU6tzyhFxw1hucKJQAUotNeUT39LU1FgSQM
/bSWnNTerJi0IV8lBhsxB0ox4tiBkWvobRiRqfJgPeKBskg4apC2VbuEmgyNNPgg
otI7A/w7KweCI8nbeGi8wrIZvwKTWCbbR0geF8YryH1cTaClJ0FLiLi4f+DDNO7L
jpI3tP/TEXghzaBbaWMDXyB+XRZV361kEiAKcZVQP2Nu1mvYLBObOU62/+nbi+1W
Do+U7d0KRH8dooQnHbx8MfDlSHd1fzZqF4psLzme0rvPExVbvkaWVpmMBn7bbmSB
rtM8FJ2EYTcO6ugfnZZeQ8jEhp8z41FuFe732OxoWlmMOVNWTsEbfIK5hJcIGyMc
sCs3aJlXGg0FMVYNcEYwVMSZy3VXMFO/ocWoSVrL9lGnSHauL3nfPnYjWJAkeucI
iZkohqsCcbpfJlpDkR9jG2KxMPQlt6GKlXNPrD3KfK7XMP5a4rUAZnXfnx0c4Ld3
KugCkFgBBEgaWUsWJGOpp4vD/cGA2Vl8ZR0sgenA3l98m/Hb+dkIoMKI+1sPEmfz
8ueRc1MjklwstVcuARo5wzge/NNfgAtfrzUNLw4J1PU96hZTsi9HZQjN4UUpjOZa
T+Db/SLVTX2fM1jj5HkbjYcg3KLn7rGXyUaL0YxnZJoM8HhdEHIyMM1CXPpoQdN6
3+CWkcBStACbVXBSE1cNjk12ZTPq8VVSZltiQ9wTVu72qFkh2VD6SS+ONbdGoNPn
rme/BJ04W84bkbeak4WiiNJnAlcDh896NSjyEPh45wk/8YJfk5Q1RelJYm2HISN1
FcZwvW0pydbmWixXip+i87oEDE7ogRfdUQOhXxXDDkyEqoWuEB0iDCbo/zKJh8wD
RbbQHvYZeqbuSq+9dmcVu17i/4I2kmkbuw2XsyQjL0Ln79CSbX0sRgcftWXHHKbL
7mY2Xd9AFNsP4sn9Cne/e7txwagafXjvhVySdfPz+l2Pmkux4q5GwGxGon/Ygm/K
2i/7Y14fELcb36AKRi7PYuhsreBfSYAog94Go5GFKl6+i4DyzJsfmcjO65P0D0JC
vNytE0NNC6KApB/4gZWP7fiEGwS4s5QuxxYVaaIb78Hol+FEBM8MUJSo/+Cupm2n
uQQoExgaJ1CciDoRGVM8lM/yp96NcT9vyFePjX0Oow7U0NIvG3l+ed1QHRWCFiU8
zRp0IYwXihS5432Tao/QrXYwSAtHUpcfo6/yBiMda29NlxTrbCQ8iBCBzI5jkxT2
`protect END_PROTECTED
