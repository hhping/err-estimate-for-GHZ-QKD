`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/6uYEEzxIGS7v/y/aaLIWSmCNDjCDrXs26clpO4RZf0mcLNnqfLJuwzunbRl0T5
0DdmRpntfAcQhM2YE24wDl9XAWKd4E/OiDBnuID0C7rpXsScZM8LmH7NRDDSNhZC
daQhc6RL0A9HDYMMs3w8wdxYtGucAuB/my74fbbMa3o/xAE/3V8MO+I2NzG6MG8a
QKXS24CGtUJVrggl3XfQl1HxDzVHxj59nOxUB3fBkmEJ2BaSxuMClQCDFYER5pyZ
viCqBNnbe/aMms4VTRQZDylYZybwRNegc7MSL5W9L/WBGeKFjI4MgtSAxOPJnE/P
vYtvjGEFMD5pVXkmib3E53fz5+9Ql6Q+anZk77p0prw7gke+Cy9vxIwzoRqBoEHT
0vSD7A2gWpUBRwkKbmxn9GwSVI+/vQi6X1w/R1R/paBaholZ46PwVcv0xIs7KmrD
YOuh/341WKvA8Sfzx1P9HyOuT/qt/zNzjMfeAqxj+xuGkMoDRbsN2/4r6dgZfyA+
2oBwN6nSyPxiTG/FhhticsLwlAUWCC+FgTOQHt1KHLASZgdGSSOuCIkxwtXcBXvi
RhdbyHMX/uj5gQj6H9UPnAYwgA99sKGWhOnNMDM40K8=
`protect END_PROTECTED
