`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHYX3CyiXkcPMkJJk4NhD6qeWZwgtaXokXLPzIfis3Cs98KnBKNo299c/vOqH5gy
D4NsSpCK6e/8O8MYfKtgsplAjHYGutV0CEqmpXLv/yLAPwYnR4SQbB9dAtxeFAeW
eEUku7XMnwSuRPhyd0Kz2Q/GiQhsX5fpiQGrzkTtj1av/+hKi/AWzUEPREvcSAzY
+PWVwigaYqVa12HXOlKmh8mWtuznUE+kfd3njL3fxDfXPGgO/E93EN/jnY+RQCml
SDpCwhiI2yJUTkh5MTahnUqqsAJXv9VPOStlUrDpAqbmoY5XblEGXNZxazsabSVH
VyXWUDRg0awcmgBwo2tgxodcvd41lPyCzBv1HarWzm44uTFExevhr7GIdEP6j3Od
V2KgHhlwVf8bLr5zAKNRsolCI3sHRCyAHLbBxx1apDmxnhvT2Gn8B4L2v4aN1F24
+YQCmAqaSHplPmkCGUyqb/b1nx6diDaXyVBHKOqGlj2JD/A8waAm9NoS/XKnVVmX
oUHOZ+U2YOKjpMRDtyEaG7l0vNDI7rubGYE4UbNT7ZpXu+E4B9F7E29D4i0g1ZU6
+Q2i31IhfPbla5XyHO875TNqf5V7hzHY0RyGFx/i6huTLA17juxsysZ8UInNin/p
jqQBDlEVd2ZuR8kredU3x/3wqnI9JOaxa+ULHRv/XS8oH6rMVb+KPaU/aLzxBe/F
gyWKLskIx1x3ejuFo9di1TcZKGvvM43TvZKLlKBEsb0nIInghtuMJYv4gsLg80/n
7Jlgoz7o9ENUuSMmWu9LWqXFii0gDdITtj6aMqQOBUkLHxxxOhRbHaImzJbo4MRd
AhIGpQkI1vw0q62QOKhB3Www3QbTF8zT99CV51hKRTe57KsDCmK2G8L1fRIfQ35X
QL4rg5gCVa/Ne7hIgGxWXRyFlEAQ0hwHr3ZxTnPWK2HWA/yia+jHlMAfIG9Gcwx4
HvLEerbC5xpmGMEnwUl3aeZvWnkaof7syzPXMdONK2Y=
`protect END_PROTECTED
