`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DF3wmYygUPx1R1ryG73G4LS7qVRFfsmBNgtrOjqNbhL5U/NailG4Z/gPV0MBP6AY
LTJmCnpRljIhuO9Y+A38/Lag4iQ0eb2Wo/87VCGMDiHE1xsmfR1jMWfwWy8BU6iM
drkWzlfAGfv01AI3eR7K/ewk4HNCH8P/AHmOlGL9mjJOzf8Fpw7JzIWfhio2tHlK
8an1z0K4f8XDllKsgnvqB0fDqwsTyyv4yI04RCK8vRnDuTnWOEXHlJkbijXwY7Mf
TpiS7SsjddNEiLzfGK4m50J/r5n8tyCtpnVJl8h81emc6+3cqvCIBAuceybyuhTw
zy0tVDMowePuJXFdbOrqIPFcsiFf2wPY26OB5qg5KiFsJhb27P3SzAg8/jSpu0jD
DqVvq1jRa2nWNwmC3h5OiusS/lrKvbi3iBp1Dc+uu19fXndCpLY4pTa6DybH3Hnx
G/W6rVWHvrEEbQzQEfVf0KXym7h3Ai281VaHLb1atSGczJArn4ipJrk5xhcF/6B1
S1aVDGh8VU0T/jZDGitMr3w51OpH2Z71qndTWT5iW4wvqBJgxvlHspUSBJG/pl4/
LtXoZlHXhbLgACfwWYH3Dms4MnLikwF6IJtheeQF6nG4Gqct9LZ5zzyHi/cBhHJ0
5e2z5seROI+bUvR87qeQYxHl44k6NM/gQjkz/CZF2slWJG7GYG4ZPkZjWeuCbM09
b6Vz2JZUuNrRIgTUmo/kLVoN4rVggv9Zu7ERN72h3zeybP/hRiMFGfWFjSm67cSK
uMEzMSgfS7Azo2oTQyqedVufBpVE/ttHkDCMN3pO2QtIwoFvVHN/zvjnSwJbzgeC
RQUiDO9FM5cOKPrXulOPD7bqqTBSsREsa+sSoc9UfChYeRiff2aTVZF2rUhIuEIJ
Sa2ksgZaaCdnwcpJlvTPxfT9xfoR5h5qDLQOOQqIYQx9A1rgW1pSsDg78V9W7MIU
w51RRTyGf8J7ZAYPBbctXQ==
`protect END_PROTECTED
