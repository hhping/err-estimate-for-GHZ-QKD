`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/2xrfCDMrgEfXYgvRU6NQTKdfFNISBoUmIlCl1aOyBXnoSw9tRH0s+XwYizOY5N
3F1pXfUXkc+98Gcf3zeNYc0SWBq5/r2mf4SEJSKs4h2wKqzs6597Rtjyrzkwij7n
DnMbv/FFEriq0XpPbgc8zS0LDFY0+eL78/D6H4PNnP/pYLthv/6sUuw5mpesFovk
b7nGhZSV6OYXVw4oJ68JDnCA4O2gzz/A9KhFUUjEo4qHXfuPtqDLZx1i4LugTaLS
VNzJlk9vZmvEa5mFTIqC/oRfeBm0/ViH4M1JG7S+qxy8tl93+4961TfeFZt5yeKE
MVsbF4yEOnRl0rYJlkuLwRSVdB9zsqjaq4uzNgjOVHpy2get/e1dK0/0vJfdh1mk
3Fu5BFu4bc1cgW3oL0gyKXzPquYSlqQn0GILoH9ghr1p0hstGDn+yKMPtUiNSph/
QdPL+d4JXkmcbvT43I+V2Ey1dU+SEi5M8vPTOZAohG9eSsQdOUlADYN1Wytj+vqB
FuAdoHqx9Fi3OBWT9c6MSzwNhMQIgfMmA8p3QYB1yG1K2mOsDM5mXtgLdLVMr6ii
Uo9pyYvWslOgm4AXGVEtHmkJ2QNl04T1KKQl1NALC091a3uRuE5s5rM7r+im0X6K
2lRF/u+T7KHLs9pIzdtAZ1cqAjbdaGgQAKVgyNya5BtZf2plkMdyUgchihhffDNk
FdHGB8jh8EOsyl4uTEZQ48pl/XhTFQOxZPp3829t/T4k7Prm35q4+bu1ueuFud01
athHjzFPMe1fVSKyORPfmgOCGBKdnTCLdJipNOcO6q/5J/0oQwZLA220Ptx90Cyl
VQ4gPl/hqczXDDUDLmKmxx7b7YsvPCa64841jSBVcxX6fWiVCVfHLEgezRXXYY4H
R+VBpYrPSNaGGfkbdreI27jsh8sFwIYYYwcUGuzTPWnHjfY0g75pXcFIxFjmFSnH
omI+52S2Kut9/fnaWdPchnWZVtRTFrpoqx7WyqI8kbCCBlo7f66N/QXQLh7YAuTk
o4oBYe5DCVjw58HXPB9U9m7iluhya+zl46asD3qZXocQkr9mbFJw0DdS6MNy2KJj
HlkvsRRpEpCUrLZ0qtgyfvHW+VbNbHELuJE9qD4ooJr/t0q2QegF1/zk1KksdNt4
QTYNUcOaswMgCGPjS4/GFXUsY5AX0pqj+XVe4RbBuXKRenJ454ZcgHxAqGF0oZn0
/Qw9v+7CBgATBFJNaChWvQk4+318xd4onUwR7o17kV2/TC6GMYrVp8X8T2Yu+4Z9
HqufUKjLNtjs8S/WRkrd0qzhA/VeqNjctokhrZZ2V79wd7WNU5/zXJK19AG/JOPx
L6JsP9ui55xlxAWfed6mNpA1k36oESqxLSpF+Fa4jyLW+gF6PLOfZLLYKHvJCPQn
8FJB1I/f9OsW+usg/JQriVDEkj7xxyngBVD5xnrB2Ych3mJ3BqDnmfXgOedTjsQZ
mEI6tGFfSTu/u9a+YX1o7/Dk+UsgzuB2sIAzm88lVuaVrTU/rTm1R2gmI6VP1axZ
1Ne55HBdt46kKMJ6NfJ3E6sDViOtp/ZGOKIBe20vq23Ia6gRd9RD8jVwmuHY4T6i
dibEvD2TbTlXHakxqV93HU0I39vrWnY7x+Kle7kkXsoL1N+YxgNUnS2cIXNz9XW5
IW3Ajco4FxbLqt8nIY/rYvsUrCYUDPqt76HR63L7ZzGLAmCGGVNRVRhMivG8QdM5
0RWYUGoW1u8TDa8ZvseCSJxiTV7sOHDkxuEhjzI94znhz3Ixr86y/HPG0H0f5OEO
p63S1Odf7nVxeURcat5QQnoMaBOO+Ny5iD5lmK8dkN0rlzZsTgaH6rLdMi55NjUW
55jIoVbuj4193z5K9pWkD+hYGi1N2O9zvqlv79eazAG6t+g3v4QdLhPNqI20O/Kf
tY543k83zzQ0Ab6Dq9jUAyb9A6GrcxjUbNWnfDRSe3TB4y6Q0EF5FEiWJffkFlSb
CTz7Els7MBh5HUpwNda/keziAdPd/TK5/6nbjrExiRKcDl4VNYKpG2AibZU6xTbz
FIucUYhcDPXfTv+NRNAYtfwW58xVfXF06Mk5WYRigFbCAzfFUkjw8LrC0CiJ+A1r
FC62a94mv+1K6TaH1eTWs2iMDWlM+2tUf7WZSfwy9V4hdHfqqp4O+mPCAei0U3jE
OEZHH0pWsdHXW2bMIh8oCFqS80uZOoF6aBUKFp3OJG5XC1b4/3TkeE0eiH89EUwV
mckiUSgRm7cka9bn/wbV7B+jgJ+1b+N8UQdOxCIV8z22go4E7AX7EbReQqX+ThkB
gBhWM4Qlba51+vUe773RyHtT84k40A3Cej0JtNJEHmmbJbmfVbyzLZnewQEB3iMn
uTVoxlvxX5Q4Vo1UF5XNAKy97tHU+GdxLARkNCCDjzCR7YNAKRooE/8bEB1dDrlg
TghI5sLZAda2PP0EhXMWsyraDbc6TsXt1S4XtkWFZX5DYtysXdUMOKzu7W+9TNlY
KO4hR89ZAOFJaZOdKWtehGEyzZb0woKTDQT8kuJ99DQWPaTjy+T9/kNBZpVIMhZE
tY16TJTRpZeOe+qsrNM7uMmyust8wA7GcNs5O6B2s32bHWNH2mJ9F6dqMr7ZmBty
xnRUtXObGpwcEpjjAspv11S4hT66QxfWhbGm8U0LlLtOqLLyIa/9z+TPdm+pDdzF
CiQtC9Kb5cE0Hm8X4+gkG5F560t+FgDWPAKs+cUPDH0HWnNh9NYrzDt2OmT7K9Ye
NceDFWl+Otg8ECpe54iaYHBZIXYCyxGTr7Ac8j3v/w0wRhlTddLaoMnpV/pzStS/
kpGZ9xUB0K8BMrThB0FnU4tkk380gcfne/eDdL1YAYyVpFToeSnhqIW151LFN4c9
VqgS3XNIhvbgoQSbW+gmzfBR25HCO2qInG7LvfzfS4wyV/keDG/qnBzv5SquaG0H
MuY/IzMsCbiDO2wOZwoNj0PtzKMlVBxCsY6dGqFgPeBQ2F7pdePmL8vFIFqe1vWG
FQebO9PTXwuBGA/Jc7FMNawDksBaelFg9FA8oKv9nNcktwt9ZO+5c73NqFAcvKVE
IThtPMM0HstFJD+eWpGLrwjn5F1u/JUFpxP1vED6gNL6CpAuIsSt3hmXc7XPTXkZ
X4TBtcpfo3ncPrFVo1kifUQ+29rZMPsRksrzyjnl355YFcH4RAYeI+oKL1Qs5+Ly
sf2/jKyvtWraW99pj/t7MpOelBQlA9H8UiscxOXcCvg=
`protect END_PROTECTED
