`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyIydSNlrlAs3J0cBZ5LXqRQK92QJYOHWvdsRWz4hjx7z0cHaoLVY91GSwmJEYYl
c+Ze5y2U2Y1VM5M2hB/u1dz47qlqG6JXGRgB7iz5mCQfU7flehAcIPggWySRar/K
1MbXcbrbIl3pFrkNntCCZ8FRu1DHCK3KUoYAmi8nCT1ci7lAEqgQvB0jC1ge+mC7
k5/r7GfLrKlGZHmPPmchhErdYJANcGWObQrONYjcxUkbssuS9d1AHWFUx05MxOnM
P8xClEC0k28wrEbbFXcgZAViTBvIDk+1hzBR/mZHHWB2C/m0B/iBvdMiodxNroEU
8yTZ2xMzUZwnGbwZn7hO07PdGtLBer0EEl9GYDLmsMP/IQ0ffnn+Jisz0buDUMrR
CAYwm00nO2kFmHiUiA1p7ozoHmWtwRlOTqnV1gMGQWTczaiY1r2N1mODGGlwFbA9
FTu30UErvzr2CIFnab6piwGjzUnI1OM0nSiEVxekYeAEJqQY/J5iYuXX2bU/BWj8
UL0Esj6vDlgyXYvUWJjN4POANffSt6lBr2BSNaAvSQPj0nS0LsEwLhOC9fIVca7a
+l2Ow2roOhboxMQsEbQImhwWYgIP8N68JwCHaJCekI4ysgCWy3occoPOl6P0RrI4
eNfdgtcocDsSZ8/ASFSW4T1H7qkfHP0XQhDzvSFGlRd3JmTzFJP88U8I2oWqEPgm
DCCB7enR/76IfRqXPLw/NvjF8bTNGPYaeHJ8Xkooi8hOcd9P3DOr3J6ATBktGX5v
oDE1pLrSMYYJ6So8nvWVa6Y2Y099l259uEQAOhPLH9I0utKDA1Kb7/ld03uYJKeJ
spVhqkl+lMz5CCGZthhABaOeyf2tB55nxVMqrG9E59MXDYxQWSfFbibGNIbTJEte
ulj4fHxVGS/yHnoKMeZSwcuOJDgf1vmp0SDqHaKEdKjQpUXTSnwBv3lJAG+SJnDY
f8TOOYZdV47yr6l0Eu9W3MmCDE3GaqOyX8HxYQK+383gQ+0FXJySI0ULTk10VTQ/
+5yfLUZGdX13U56S+CFQiAkvvCSj9Al/05N2kEbp9fPRGRatSFl+a4jBRcd37UBr
DWatQc5biWP3L+/PeSxaXSm5ULAzbFnZKwn0sp15tkacUjqoupGHdHH9k7Mh0Y8y
4H6zUoOzflfqjCarggENNk4jgbEDFe3tjgPkP6qNNme0b+u4fykq3s8iFK0YWWC2
knZpiR+r8GqyxtZx9utYTy49G0IMIJhfOxetM9rzJnNvPw0epVKLWXwsw0n16DPT
uFPnhIuwYzeZvUTA9R1Cg8DmVwd0SfaaGhbF82W841EYAgZnoGgdqOVr5UL8HrsZ
RJ5/28BYolnQpyp0phfKpO1lcyW15fFmMc5EwxC/YqAVXuHYzSARaoZB+WEvgm2f
AgSfeLYlRv+3W3jUKhlfVU6WdmMniSCLr6qU0jkdzl41np3LVKPP0aU3F/90Hxg7
TMETCa1yzSWXJQ2i28dPbvexRfVdvVUfko0bKEh758he7TEWMq6HBycnmT6j0R3k
39/Yu0GBArV2k3Jq3H9/HS9XXu/nOwj+QZc1SeWLdBSb4pcMvYubdgGZcDkKA976
IilVj5q1CLAlNn4AODEHXMO58WpvggIB3OkOPirExaXwExjcwmHYlUxDvh3JpTB/
yU1jEJ93cXGokywqMBOMjYCq6Dsq1lu4BUlZr5Mxxb9eyAIv3GqgcAKtbY1Bt8xQ
E8ydQVIjdNgxIJZdsmVA2+co1wuwzPLvUkdmGCZ5f+34rpuaENWevcncVS/cnuYJ
5eOyZUQDORhRi2OLJbOf7dlfb5IfZaQGPzUHwvSaQeG/W7qafifErkvhRQCrxDhp
ODTiVw+JXs74w7Z1Mq5Gf4Lk7JU496JVFD0NyLuih9eqNKdJUSaXkSa6/yRazRfW
EYfnZVsgxdWYshK1wXbX8reVQW3OQBiJTUwu7wdTSMfohy0uvrFdFCioVgNC8eoe
1dutSNz4mFZhx2zlO6/Y9vLfdZOKsROb9qGUNK3K6pRyDAgcwMQq5Y8g3A7niPZ1
Ye1S/GwqXf0VQatFoDJ6YyJOLRBpP3o1kYdu6/2VMYc7LPaHLviSa4AlwsNhAoEx
FzGd5+Xet47fTVUtsuPEVoKLVro4r65uJds5dQC8a+1SIJ/mkiphC6rGRz2xP7cP
PGnSv7Vb3pinN4ZMvx2LlsSs/Wcy4y00a6ynMx7byFDdNhdu2koBrcP/XS59Y5+g
sDJLbq8eaYCKmRAN75ZqFheDnSBl055YwCTSyh3nQNrEvYujrFp1joFRTWRHIcgR
/tRqutmsZMLWd5Y2cxbXkyJz0AahpMNcVAzIbfoSAt6DfHFglGky6dKLq6gtFmV7
0RZ8Cptv3zHgz5PCGpxOZLmhOA0kTd6bngAJad1zeCG4dxcZNNNIwW9vS4rxbEh6
wmMplxcuKxeztKfQNRKrXJSpsflKueJK0hNSo/i7sbF/2lYWygFA+LFGOOEjfoF4
87Lv44IzlrtiPGbtmPQc9DOhy1RuCSSj2+NBJbUiATTgy+Wgiy7DlP66lGNCBBct
cCWEVjZXgljuZokdOnHTzoXMnPgKbRhUSMrQO+E8OvQGjK/DbOc1Hs6dvFv7ILnj
Z+jSbE2dUOLRqH03NrS8wFI6sEy+Gb4k7eFEPmJz45fp4oFNlqZLYCOGPxBD6SRD
xhf+FzYfVwDLc4VcnnjLEBPmFtk1joFROImaU9Y6QLG5gFtgFv/DIpoT+5SU7ZgE
5BeQEhJxtMjyf1SG+/DEHseyL8zvUi+8nbYjZKtovl8tfgDsJ2f9m8dSEMtvwAjZ
f7TN724R0aEL5rfd5xTgJN862UJ3JQXgTKL7xHOfEy8u2urPovyOoTf/6CvzZ1vy
sQfDgz9RZe68pZXUJIpuIJUBdMxQvrVyTIohqSbckzTmvsK9YRHVJFQeb9QZ8vFn
lTfbPEMMPD3YuEZwioN6oB6ShqiuN0Qor96SDMQ9/AYFYt/F0W7ehUuRLlegNlRc
Y+yrot1M2lJQR56d9hxcu3MlfI1ziCCy4J9hZltnJAD0U6CoS+/1wmoGHhc/NawM
P+G2mYiy6/4ZhTrHrUNLaVmt3RRDOLvdhZ4wMQV0xpdpwxS2EyoHojowOdVpkDSM
xFe+2gjXQxQn2tlPv88t+D7BWeeICa8ViJJCNB+q+3aUzZOWLA5X3OtSMWuQkp0g
+4cgi7MGTQf+3he/JYF1/idJApOd3ONb6XPWn0HX4AjbcQJ7gUn1VJcD6yqEYv5m
9y8zWqdoNoC7agiUQwAQXnqLkEkZ8tzKRlSmEdrOJMoAUPXbUjkWtcM4UjrmEFrA
oj7s+HY8mIUD2YjnEEOoX0CuDrDTq9Cpr4I5gzGnL3NQTyLfAF5+dJ+7xiN+Gb7T
vtNDMDVj7+oBSoMJfXmb08Q+1q+Y/CSsmNJPLzlOH2IRBCJ9LbY1rvYjIa/e0osJ
88G09ZLOS+pVUfYz014o+Lr9AIf1haHaKE7xFWvdHpOU8Jgolv84KbnTIv8dlLr2
/kEAUxeNY2BTBaNaXm4VGU1CbLxjMO5lypKGPto7sAX3JIEHwCO7bTR6WV+plV7w
he5WDE9ol0FOA4nmr4/QvStJp1srZqtF8ezpEBSjXstuRV4jDNna2J6IE6B4CEgf
zDwetInwThfvEvYGgCsk3GtOmyjWyX3HdqwC9yUDUNZ3XQEx3rrQXbJjyXAmRevM
gE2U4BFvNuE3FfM1Q+ARPtpo8lhMkii6lOaV7fOW1AwwRBgb/l0wwGEADAnpPc/o
d4xE9Ee+RldRwDzEJc6RJtkElSqEuElbYWmonpzBIu5NW44P/dICEDAsXHDT1scY
+hlpdSO/ctPlUzTRhe/zH4rSWG09E7b+lDThy3+/tDzORwhF9dPPxEFK+9ZyzYg1
piQjjP6uzN6XJsUnzJ7lRdB5AgTdwM1186si0T8GmjoKdWORiUm+HZ+OZVBFE9F2
ShimNHt9FKYb4lfvP08TRFj60aMKUVVpnmP6zH1JblXIkMdN4oTyq44Q4QTi3WWI
qo4AggZRf53KruGdIMPWG/kSG+0v8eYwi3aYoNrz8VMzdHwJR6tOm8FCkZNZIx19
CIXFBXfF2RSqbIK2jKRWQGOZNjPX6EgNMn0r+KgI+MiLg1mFO0hupfbJG41w4Uk4
saNBRDem/mJYq6JesovFcjKBRENglZYyMy81g3yxTFCqKRj7zZlaRo/+UUZMAddn
001+xwBiSYmSaOFCwVaIs7oSNfdqrLSUNuN9cdygn5YPFYU0S751CuatN5BoO8nd
fJtY3y5JkHqQv+dZrQXVR7/G340TjQ3P1iiTmvvLqRjffKXhCC+aibs8cnNix+3t
CaYsjx7Z0IONWZd2lRGFQeaNTeTC0JluChc5IRh9DOOZ6t1++XeMKzaLt+kFBNFB
hEeeh8aSYBK8ciuElkjw3J7xGWk2mesLS8JlD0gbBM/vDqA4I5NGtCeW2v/wGqQ/
zHftFphW/wTaTYqx1FZjV7dx5Y8jAH0osm7hSfR28Y7PkrIjs2u5WOTihZLzILI7
ueGRwbm4TL+tG54ZKID3OnQnOMO0QBAX66VteHfDUB22dGe9IeO3tO0oMEumX5Qe
7BTxcB4cFq4FHYXkwNrrieH6LVc0Ug1SKrEuO/n4+DHZ7eXJV5GrIdomNGJx8cpe
IaMbYQr0mx4V99SnntEVGakBzFFt5TiSl23XPCU44UTI7bbYZOQYa9s1eYVTDsCm
CQehSkPcZeqaVLzdzrk3whuKN95B5vnD7uhq6/geKlw0OKSY1niTgBAdE5i2iR5J
QJUdP5x2n2V6H/Xsn4aNuRc0esvv8no3xLN7Xgd5IxG0iNY3HrRMyKqLp5r1jf2z
OAS0Oo8QBiEHelYTla+X4Zt2GCLw6VqXvHEvlHyQUHRyPJv++8n/COHIY7W5NGdK
K7N8gJt+bDQAjHubTfGAywxGczYmf/4DWJ95XdeCugq01OFJzNTeTidsI87/2EwE
f2ILbJldAi7EwPLxk4CksKdbtZSQD7a1N2iu+DM5uifeXKVbX95Pyj4Atb/KIJGX
FhE6DUxk26YMSIZpxOfLwd5pplLudEe1Rkum2pvixmmBxW/3M5PLm8rKYRB3Evxe
8ZtD7JiqcJihaND2WbxqJWgHNFCb1KiZEqwd+W35gVMZv1MGwGie0Df8UE/Obo/u
0HMUvnDTICBttuDK1I8+SockJYrvyWmdgKmkIq8DmMsvsNODYLol35Rd3S2OjtCV
IJMh/3ae1tXkfgrejWzXpUu5/hGqy9xLPKpZtkm6WXI+6BC8ZYQj2uoCgJzjuZIQ
jq6bfh0iG+YL1992/PvYDJIrc82h7Ukm11wkZJYkQpmD76TxqEgHIcEvYJVqhAb2
DQg/+Garij5eQE+EbUynxe+VV6YQFog+bzLIvcFWmlBrNpW8fvl2a81g/hnzqWEn
zaNmTQpYzOfSv7LQQgRU/C5tsWJ1fRiQPxxtMtS8MK2quqpT858H811lq6da2Xy5
Hu8JCPgC/1BJ1lRgCyjoH3yitF9F8Jq/H0Fa5xzYAYBPurCA7tKswjEu+KG6z7E9
Gp3VYZgW1vEEsYRZeavpd6GI3ts59C88MhBwZFVR6nhlYviAjpd4ZK/CLtK0Kary
B7cEPbor0pR+fR3IkMcwsJo9qnalzepRCFh11QNe5wBPxP06k/NTGf9pLuYg4g4m
vdY99T8heQ8DWTih3jot1939+dflUJEHOHXvIdbj1+s1K4BkmXEUnTqRF/1CkpN3
LXpGxxony1TE9koagB8ae+M9tc+BNbEmEkYqFuPyx9Sil001GIski65QP1Dpy/K5
JOtx2T9AOtVZf05ML+Lw4dq8/yqdjFinR9ZCCh+lVulefU25OQSRssU/6RNTickb
+TBw8tOK1sIWqXzVTQvFeojIh4nPNbhnaRhP/nh6K5HFYk3mKZf3s6e5HIHg7Zoy
Z9wU9BCBrC6yW8Y3BsU7PZCegmqipNy//DdQTESzMi90/qjkYNTk7Bb1BIpLF4h/
9Yfxh2IzE/eBbCrED9LR7ZZtYECb1/vamw9Cz7eds4zKKhCJr0yrcJFwQYU5KUCp
6Q2U8ok73veyHmLC7WJeD6Tje+r/2eZmX+47dO83FVAamOnTE6oCtckPALa+0deX
Ggcdad3wKhjtAkOnwkaXfxwUgyE6WxaLdxxn1ogEKEiG3LywSQta9R9eS4tqAzrc
yyHD77keswwQMocT0illyAN+seJ5oPrMug05zn7S6BBEEIjtd3GRfxyPhaSZLbcD
cb8iF4BZARrURQIvrz0bZPW6ZZtXmzL2i2FrxAUI2v5pyaMx8OGhkc9/8Tnxltz/
1ZFooBKRJaAg7AA0fW2vIT5u/45Pn5qim8bTGHEqDugcajCvTxzzXR3HJa2tws8C
y2RUuA+WrZLLmJVBrwMDo2uoD8U24pw8aEoPLEZbLE3/Zzi7tGPeL5aA7MEQjYsu
5MLxyU+QLGU/R36el0oN4mT2iv4Oub+bJJyoszXTOel40V3RKar71K1PzAIv74St
IZGBxoMPuuskIpKpYje3sYBtfIWddpZ9MuVlgPzg3jdAssjHvlXcFMiYRd1wGjqo
9WIx38z0TM4B/hll0h+yk1cCRo1Z9Oe3rNzq8tIXpOpsGk19GUwdMy/7bCbs2CGm
Vb2C1R9d53oZVbbKUm8bXOUramIsEU9BYvoRNuJm437/Ns2YtblnfZaIbXwBGLmq
I/DGqGS+omQyGJg3oknU3ESA2Ch5uWhUxd9YOmi0EfdTT6eLDW7APMp7ipPn6AuA
ADk4ZCGeWYGxMXLTUVTG73QRExrnCEVMTZUsXxYl/w0TOFnzNQEkpVQsiJRHYgIS
bS0FyLZSZ7h8V3MaTI3+Ljr+mzKWpMTBhHkOUWAnlbfdx0ePFq7ikLLOnNhS3ynS
Xqdh6haGPcQwVNm7ku2Po9Vm/A/JDdUkAtoE2TrVYs8PzT4TNqJ9gYNVRQBVF2jm
PVxpGO8ShXXSqy/mQkLCexc5fF1D+R3bwwipF7joC3nYSJTeBV8sSPRXId8YQhRb
/JLQXHfmEVkVMp52oQqj78VT419/NCEsv7AHArxs/uul7zZEHUZjZ9nHE99TsvZp
YsKC55amspD8pw+FAuGFuRAdL0/DEOExhUmfCztSkB/3dUPw++3/A3aoX+hqb/Y8
VMsP7qdJWRkB/Q/KpZb3wdjpEIiwGTacn3dD6eH00tT4MUxSPUCwvjgcED0++S6h
tGBcgctL7ikGslJc1ADVfbEtm6yctQOAuLQp3d1ooZPTSfK0sf0EUIqa64UM/wfW
hKrsr6kEScpM4PtC8iEd4afjsAwYC4jUo85umhIEvRrviT3B9N1hpRxOlsXCzXme
wovU6ZVDSWb/yWVZTDqVDbGHoFTykAuF52j2JhTtHQ+HqaUf7pk8cdl9Aqc6IK//
zLG4qOrYyGtjHPSxX+Nyt0TljSxQLFuUHJ1GRopD6aqWI1mPUQQFr9gfGddLWQ0s
Fdez0KwSm70zlhulkkwO7OkZncZae/YH3UM58kQotA1q4usqS7TbK2MpL73hcnom
kcCI/44cmnd0Jk3MxiQmyJmilsDaWLTRGWmbJA14xEdAtJ+/FZCKIjDed7cLOlQP
ehU1tpi7tcWYMPisFJor6J+j7stLWtU/h9v1M8419ygyCHoM6YrlbR8X/AeuW3vN
M89OyEu7b3sqykc9k78lPYhbsks88afntNjACp/pV0iUbL0iPIkJ9Ov0m/JYmEof
7rwtaTZXPULKrnWOD2BUf6X9Pb263Um/vr8IUv6Nlz788f/+AR6ClQptlt6qThzB
KAXzSXSyDDrcsfllbXU/Lm7nq/0JHXcUnPCYheBr6cbEL86DYODYhEPmmQb+K7Va
z4b6FcGrbS0w9EpzOQ0G6bZ6VIGt7Fe9Heo1plVkFYOTnp3NRjMo9UWu7ieeFI+s
w8jEXExZKlBio6KkpyjXiUOf8XFEdSBuZTstjNHwpU1VL9fJ+Um/zMbjYhUOCWol
9ZNjfj9zZ+0VyshC9SKKSOlADAFetb/fm3UwJnuqorR9ItTKPBFRxB8Pz2L2bLOJ
ftxSEXn4xNVmn1XisZ7e1MDulBkQVEaWCfgUvWJ0rRAFxk3+CmvwFw+uSvc6f+8H
JlLai6lcslfXk3jWt9zquuEnnEcftwC3FdmxbQoenwJNrY5KI5ugVCnkz22Q01c2
CQv9r/Z6wMRxqoGd9akit6YAWlYfViK7gy2KfX3YBvvvJWHopSqNXE4+CTIgSuZg
W8f9VucMOseqplxLcYlLkVIxZBc7sNVefaIjs8FSVZ/owa6X9CE1zBRk6FIcDkfH
`protect END_PROTECTED
