`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4UzFJiWcSLsIcW4w8CU+bAfKLoOU+97q6nIxe0fenskusiHkXT1FDrTJSRkfG76w
WNxd1BfkOLWM3XgN9SffLZYoDIbBoR4k4zsLhj62k49ofOIrkDPr8763B7K8kYPO
dc+AB/wy8ynpwUM9+DsD/KvhJ+vbZ1tfJaS2NL556R1yMmkXN7cNMh+GNTS0FYy0
KpLIkL1Ikappg96AzeE/iNgb6REPkvOVIBYaxm7PEgMdGKHNPBkXNsTXW2dGsuo7
e3v17tKYv/79Z1VrebSQRQOdGHN9/8etakZgpdtHQqIUL4yqvtU1C/ueH+abtr3M
iPzwCIsGqWcLVRJT0iKe0l/jW4d2xBM5liJtbXlfBIqenCO2Tn2FdCutMcpFOhqB
zX17gnYZIYAKnazqVMjgLv8SuegVCizchstD/JfUfIQ9PRlRlj9Oty8IdsojjAxH
szcw+mBN5T8RYP/bYtzV4wfh+rhZPX/bSRglm7r1vRdoDz87d0hc59McgKE0f64H
4IjcILw+cZR7o73aSmQJwP6eUXhNyjAB6UXX0HWh2Mm4mONIRT+h0d7KIlzFxuOX
g4Ya3I3LoN/1chk+2V3YwyqiJJn05QL5pJqMyf+wXamEHXz5uEvprKBAFf9ldxCx
ji67fX9d14BKg9Sr4M5awS1nVlofET+vw50tAOHzLq/zEXDQM88Q45sHN6y3Sgml
J0iPap3CiOt+suxnm513DprvMSuF1KFFagZWVv8QaqL5DRr5vM/mB0xk02Wum8cb
69/BeL147evZZSUQxznKcq6xWSNj0GQsatpXlVHgxQBUdVW+aCO+txlP4wjD9Tue
`protect END_PROTECTED
