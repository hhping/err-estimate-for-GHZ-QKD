`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrElMddIfj5o7tzjTaDtViiIsoUeSZuP+hKlCwWvBlBDfm7FLC4kVRe1vsJ5abbZ
y2lVgAu9qF0u7VrVdQEbPWKAV/AUGRwBMzccN9VfiJ3PGRHB+iZeYIrBaT1u8bCo
KhNk6FNfv+MjLWt9hKuZgj/xSbwOnMdbWot5kB1B8LbeUYwjNbp64AsQu4Q+toKR
bnCl75BVVW6jhalhPOT9Y2949YOEz9fBjoFl8WinSoqBylDc6vuHD/9PlhkD2cZi
+WvDu4SbpWocoVEZ3h7QrzOdQAa0cQ7C4UCYSPZhbB4UfujT3Cb6jq+bWCoSH2xw
pWF1C7QSdHZv4CgmvoAHgETQAQ9E+DLUzS2dVPmMMtGQCF6nXzuTdYw3OeZnAotZ
WSuXJzU7IYgoWJ4y5ABtdHa0O+hmJnSFAK2OydhPMO2WUA1JQecJLvxMK7IyjNQL
MD4mzEMx7xGmwporz6BwU8ElHUwq1TCVRV7+3zBK1uAFufdZ9lexsMiU4XIPHAGd
uKQaQi5oaPxnnT+MzvPw15gqk4PyWoFLeF3TelQ4SAt52SsfEWuXX28laY2ndVmz
TYK1fAodGn9W4gEF6h+RjSOF7CGNkRLv0ELWO3FW1CNmLav/5MG+sk8Hlf8MUA+h
kyHAD7+8uPT88osczkbZOe2IzGa7SHfVUlMV+MMcNUS2XKT+BroQz/jIm0q+mzAX
uWlwPqAUASMRjtz9svdwuFBFbHeB+75V9NOTFjq7MsF/V0addcOxKv3P3tmBdzkw
FLGpOY75hPse6aEM1y/lqfQxSi/PulGGamzCkLT5LXrskOY3aXtmg4AbqTodylj/
/uy19yxmnI6E8nUKnWTCplRotQ34BgqHZllsPvZnm9oarU13SOtfZAA7TgA9MOl/
rQtx1FE6RXUWXeYILMEO/kKf5XZNMcx/raJEZ1Kk6Go=
`protect END_PROTECTED
