`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f3pgezNnvfKSdMYm81JG/llDN6wgwJk5hmM3NvQsmtcZufTrTwJEBhfMLZCyrq6O
VoqKd8ZhkfjKyWGJZ1K7fgCubnpyIqxPnyuXEYyUJq4K1mGkoDObuXHl9aY3ompc
3ExMFWJOXgvLuQ/pVK1FIpMSaC63ja/MnO49W7ClIrGaPw00q+FjFztERWFT91vh
Sc5vXyStRxIPyePVKVT0J+W3stcDBAwZQCm/LsF6JUFH2pz13+h2OldFFW0YOur+
MSd1AmHCghAXPSjk8LVAKyZ3e2B8Z5bdDedPdM6PXDN0wsNINPe8jA5WYFY7FMFL
ZVaJ+oZM7clja30E6cQDT/Hy/lTo11+HdpXr61qSk6XCjcAEhCkfgXWemL7zqil+
E1vTEs7pCSRgQ4i2uwDuLYtNbv/KTfMdxceD3G+//a4GgQuP+GlwGBG8sifG8XeD
Yfv3xYb9wSFKB72LG9W02JB4tCyC8oYJHiSToHRuQdj5gbl01DEmbaFZ14hqoXwG
2s3zoDTSrddmCRv5mtllBIMDmFA2shDReyPJqNuwRB/tzmqr9VCb4wmYmhpaBvPu
k/kGW+MQDZPAOtIbe0idX7Rw9K5j4G0CE2BnJYMnuanaUPsS5/P8LKlyCTI01bVJ
tech+lQhhbvCSO044sClRbUt/PVyhPQBN0YpaldaCnliXFGQq4AAtK2nWUx2tKre
/8X10oBFwy8MUXzkjRQV9EuiCYtL9fpFxPr1kLftZ20jjuACRtXhYAuf4nclaInP
URsOv2OGG84CnzEK19jNmkIB1ofaZYs/UA6taPNK3yqh5JdnuoefeFrXmQgFZDEX
h609JkR8WvDel3GKUmG5kcYxaGv/3/zHNGXopKaJcM71e2p0VYjwhDibZKT+YA/3
q+XBS1OfJlZ4W7DHxpPqESt2vvg+S2acpF6uCNEb6fmPLsGrvduEB3saz5fv7nHr
ivkRdtAWdmQmdRpCSfQiGablRnxe/fxw6AtdGJ8//dp8seSwDqpYU5CChjtPSnG5
q5AXX5c0jcA5oTT3q/cXEDt2hXt0XRi78t8YbEXcbfv4LXdYCDA4BTWniV4uGCd2
b1iyoHpw6kxTf1w69ZQjX+AH1EI7JaykmClASZHboZQEBGf4+qnuTbEkx89BI1bE
Z70/7mqgLpaQ5TDSbcM0PzotkQvpf6PEInAImwGvjOKzpdJ05XO31H0joLUw9Ps+
5HAw8D/cqLjXNGiKIikJQQymEeRkurZYBxXuecYdtWr9m2zYiXhCnw68zBBXKMDP
Qpi25yK7nZCqsc5myJCs6SvWQZTHrRis6pJ/Nx+UyMuLK/FXsC5QmA67Fnc+GCgQ
STgzXmgUw5iActWm9WI82T82Ihb0kQgSXMltz20irznxX7f2aKvwE1Hi76fxdzd/
wVO6MZJN10acxWn6jmqCzJ9eCQzZ4CmAsmnueCjRSE4DVxwPj/CXXGIwB0iA7KCA
5ajjmC9KVPxYbeg0mv33dQ==
`protect END_PROTECTED
