`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1u4mP/P5CABU6kiBFDnjdbgImbr1xIJDaRSOXVXwqBSZevKDOzanWOh7OMHlR9iC
oKBExl2/DEI2cZoi2pWpwUfJQ9nc4wS90s2ug+PF6xrzenH1bh7+y3BUzWX56+Df
sjswXti7lcL/W4QZvXa73BDfl2H4FHa+X9GxW8/c8i4MnpDI1l+s3zd8P+mO63QC
frgnMVOzWs9uauAzKgOPz7eYaLzH/SGi6QYTb8kGZhhYcU+OQ09U9HaHS7HJlW4y
IgeKR8hjkiwBJcp/uXoKkLl9xqP4soKBvE0rk++nnr97KIlyGltgYvk3yN4T4dbQ
VG9jd4wF/2ZiDFoBOHHKxyQ3dBWYJUrvzvtJMr/Qlqp3/FNaCUwChD/iuP9RbXtF
1jkMAZcLS+mB2wnUGipDmvFUVzZvCUgEkYknJ5MQhtqp40jo5RvXx0HbAFxOpBuV
V61SyXvvDk2NuhWk67+Epl2ijdqXri9U9hOsSWlqTuTbsNp90VXV6iq8dNLgMSC3
EthmTV2zhvbGvOrgO5sVK8ORiEmQxlBuUfiH0SiSsRL77Ab4JVh+BDm9oBmgjYDf
yWpyYhl4jHQMRhF9kg2wxILilVKVwvv1Pmb5qaoM7+6fJVlosxAPMDwVAnTqCqFD
kKAqp2qjsH28L6Ie1TtD+/zrkvL2zoZcxy6JjND3vmmkxVUnsLRSymUSdnZYZgjL
ys0LHm9DjuUQr94JcUOQSeW+IXA/xBSOX2DCx4AsB3bmCh8eS+wrvqr4OLTMmNw2
vN66Eghvbr1tnVWF2lHhVNSvV0NlAuaDw6bGdWC5zc2GFxicy3BHnzpuhz6/LOmQ
GfixM+y7mnAfn+e6PniPYhZt2k5JDoIPqAEihyqupqejcBJCknFq+Pnt7011Y+si
ApaStoBVGwNMKTvxxs5fMrr28IMr3nm/GWmnkR54Sl/mE/4pU38K17OjMxNMnutu
xkjaWvnaM9JJi08jB658Q7k5Zvrre/dUgvFElfd1i4haXu2lrAqcGA01rLXNMMZJ
xLFlBFQFGqi2+ApN9AUx7gCm3DSSHOuA4BCqWnpHa+DBVgNaM4Y/IXJDMmJGjq9z
YLLOduJOeYrFUhUhtPg2PtU4GWaykUX+QkjNENTZAhclInrq2qPZm50UGYfktcW0
Ru2UWVwpvOPTgVmXYiGQPpk3CxrQiCr0uKcQ75uLylQ=
`protect END_PROTECTED
