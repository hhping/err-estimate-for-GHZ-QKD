`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bom7KFGPDjZQza2QBN8y7E0xkyXXj936Wb4cpSNh7k9NsUO9mhl7bYRdenuGvdDs
Zkhnzd7YotJgMcKidPVHjP1vvM4YwYOhmbF1HY7DF/Sz1xBbjS5aMjXWSexxAOGM
jQz5iI8SZwvHj+3tOjizIP5mQO3B4s7xBuJZ3zvAyGS0Y3zMY9PuKkggfkQBJORa
BLOcnrx8KE5bN/B2duF0u3+C3dQ8EVud7IKz/uhoXVvZUYeBaYCSE4kcxT2AxlMa
9G28PTtTNETyE9HEpjNGlmZc59wnqzbi+/4tVfPVnZcGBJeCbNdvFyjy3tA79o2i
ymAAFaNNUHLLZEfmOGSDGC3JdeD86gyRDHaJVmaVLc1FQ6M7u6KO6p1oQsd9drEo
U+rS7GZvrbLZufzuw8ZXgB8AkyNTwI/xzQ9F/K3ie7W+n8VcDHGYh+Vp8+emucEA
cZ6v1jEoOjnn5zhlP7b5+vtXYy72MU9a+BAuKV67IqhSs/VRsCCxD3qMfSmHaD4l
gejrQykaFocje0NmbswzDR4n/Ecyx1tMBY9ZXDUau/nPaErCu9ElVwBT8AzlVfDx
m+Fqrr1NRuKIFHxLv2a6owqapjTGy97EBuJG3rt1sFn/rRX1Le2XmlHW1hsznxhh
CYSJdFz1iESQSXinUpmpq/lHZSu2WKFiHk83js6hkElXpRKLaNilWYisYiENYm8x
B3u5IHj66Mt6bLNrP776UFP5vwtdP8KZBu7kowjNwY6RKfrjq8GhNmtd9wItLv3m
TlZd37N3BekSD1dbIL/0dgvK47XAxpQIlw1dieuxrTStHFsk+0gFG+vdwXIZwJTs
CyQuYdUsR2VZD1pXKw4VAEczYF5rkqMx8/DOw7ZE8v76WoU2YnEAccq5jK5Ja3rs
rqs4bNQO2nv2kVLYTTn+Z2oj34VpAKeAZLU6IhgU4P+elvP0rgj47wAP/lyIEEjb
IQQXjyA3LOCmsR/i+jWiE+dcBkXViYDAESNe8V0U9yUl9UW4+eJ+A9rwDo8MCBWx
uFyB3jYIkyVB0IgE3TZHIbCjmjY9yPZmsO374/iGGCs2jLPm6Izk6xxj6s76p26Y
uJZMtBxcOkCMZ8Qu51iaD0Qgs7Lrx3mjV8nhyMGwoaAxv2+1UgQvE10SDUDXqA6C
yd3kc4NoxYIYXaoHcGa9j9lRkreh5HORWGXZ12AFJR3jX1EJeyBvI2T/hlR2C8Q3
Z7UkA0nEhN8bpR2JqQSqaRCsuU02BNUp5jDegjRKlM87HQEsjyIX2uCQGGGEInVD
iu+Ga8YOdRgyrzm/86kgzl4Amn87lt+3gcbtVtQTpaWRD3J0XJTSfB/Qm61IjC3t
3Opi4HMq6k8SzQ6SZqcYhc5NfTCunOxD1++htvLDx/NMIkUKdZaYnIcy+CuDvZnQ
zbu1eKph4zHiCclhr7vU+i6NWvIQ3VidRG9JHzdizxlW2+fC690q5h+aRXTu7X3q
ltSlyWvVUgp6KXEvJbbcR1s4ntUXPqoh2dPxirG5LuhUY8HTyT1/ZoogYFQnvnvD
2QGbrCHyYF2i9ViMgaCF1i0phupnnK/Ub0Lk63HymlM2iwTvXPE3GSoQS7GjPXPe
PMvV7YY/DNNiVq4rFLEDZLr1M/pJOix40j1kK0uuk1gJpOlIBBcaW5mUqA9u6R16
LTrKBwg+L+0cFIWPm8GZqrgJ6ZFphNvq1hy7MZyRw2a8GW8uTL2RTLfdOAKIyGWv
7zFkQNlyLeMQkRxEIfpogdAN+lvYD6FkujZJCfjdJqM7YxXdAvqpNHO5tCGYGfbz
Ew73yRCm9nj3NmClYCLQrT2ISvaDJZNPJl5dqKZnVwBRxzM/PMQnQSZuFuAuCr9v
VXuLpdpIdWpb+hSl0LQKfbplTAHd0usu2qNWTb0HwE/N7ClJnMRDrl8ZBCkjFlPw
pgDTZc9IaR59KCIVu6vrzNd9sbe21C/TJM57N+uW28HfeINLFKqRQf9oD78n46fz
djSVir82JadRaGp5HmPG5kBq0BTdwGwFF6dsXL8WGttrwtCg4Z7lYny59Efkbzn8
UBJCq5tkrc2B3ig+emk6Rz4NKrTx/0Iyu1q/lx8fGgebcBrSCTu83hyAQOGZuPWb
6DhqBhk84hXwSv0QkhuM+pGLPFm0s/ASAwGhC+tAEngunTo09bwuSak2IiF8BlnE
cyynZ0ZhSshTmQ2ky95gxEEy5jHhOFomC3Wv1sJ8KKzJoDUPJDgLtH3TZOfBwLZL
fGBJ8B6bgCtRFNHEBQosTyAdIHxsopmxx8M3jVE0qAxHsTKWZUk6d+SwXfaNV1ZN
BpjyLyMXl95QUX07N5Slc/Iw/XTd6E6m0fH0ERivMS7TOJimciwB6cNkZ+ExRzK9
hp8OVfyIYMGxp25PgdsIYKOj0qQDYCByQnr3ezbBiYbwuO4E+y7xESC3Pqypz/Ya
gP1R2+QK1odCRDG8gSlQsR4EuZELI/NOyZUIoFNBO7M3oXcOiWH/SIfXGYSI+QLg
jQKKeiDlhYgF6La5f/kNylSmpLBC7uMhCaB2nkwnmP9jXomijzh/DQ75HQEfAHuc
yAAysI/PZN01Ta8hINMWMSHtYsssHJ3/RItNcQY6DKkNubaZsuoE3ZI1OINbttTK
5WGzLS2tMB1/5NwkVzRNSQ303I55z2ql1TOv2ueiYR6uFuP44jktObx1LF9PQcvd
oxr2hgLBB4APQxQu9pLIrXaqX/XLt8d5HUkkzUElM3n3i2hv8pH3LvQr990HprtP
7fMkSzM+Rnjo/PU22GWoteTfrlhf8sXtvZA9aPXOSq9dsLLR8W95W2NNEexdIO9T
9cIdzKTVt2XfOIKn/YqRj356c36b00agDupylWZOC5nM4sFuFapbv8a4y4RmAN+U
Aq4odNZS6jFBXcrRCMrBeg==
`protect END_PROTECTED
