`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lfwq+eq9pc9vaG5k4hHIdj04TEeycPNzj4mGcqjRybCXiwBHkw2svLWLUieC+3i6
8bKYzymdVKtFKastkA7pXWhTf23aLjQvG78T4KyOGzmKO479oDhGtfLlo60Ti5sX
zSeKummhoIo0fu+BLRESOyNoO/Kr3LOiCThdliOwn0F9vXaHxjsCSjIQoPhLa8fO
50FL8gnBnBkTNejIpi/uNqAAsdr3dStnJdiTx3onKAl3CZPkjN+h7E0p/qnafkbG
VPf+VGeAk2thKfmyhMI7QfD5gzdDrEgqSf2xC/13owHslBzkdDMWLpM0HtTq4LOS
wk38cjDtyRvx9EmdY+D1FQec+mAvYCUdTptzTS1e1I7Ey5519mqBDK7ZfTALR0gA
V+f3j59Mr5bP6+DCVDdA0cKD4vou+MYA8YsVMGy46I9zXrir0JR46j2C0bOnki5w
ay+M23Cbk+DEaWxne1osL74OnTXVoCxsM5dk0o8lNTihvIrqt4awNlNyyGy+v9fC
Mz7CY0B1Wc5iCRJ9X291dhC8yKXKxk5WcCPOQ+lJJ1OnQbX6tD2PWYgKhcv1ektP
ySfS9Y1/A0uYlTVQBh0XCUX1ocPCp23Ym8o9o90htBFszSxFjXHi+ffVbIkiv4VH
uuI4hjC/ZrbYPrfhchl50jIPEksSBFZJNl7vgQieRZQlqXeqgeh7h+qXm9pv87W7
+Ok7K+7GfSRG/rQ646jl4Rk2lzCGpj/GDiTxAyWW22JiXFWLDAJBmkjUENYPlAcZ
xt6HzyA/5mBNTsorwbSdSK8KIjm1h0vUcVLNfuXckcZ6YTaDWpbNrgRg+jMmU6/Z
FJ5bqxpQnBJ6WPQl5mOUpQ==
`protect END_PROTECTED
