`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkRgd3cI7VOm7fBqpglRvbbiHY8sx3f3QU2jzS+eGKFK13fsWQq2y7xaGpE4zAcm
N5UlP9/4u3RNCSqHpmhjkzmmoeMLu0L87n6nGv76//zwIgBQJC9SQR+gDFi58Wdl
8SZRMRSQOfmjJh8aleq9EkX8TpmGKD+QA9xFztc3i7ErJCsfqqfoN6MsVpkKTd+W
NqJzJAWpMeu0qVY5Xjjh/AFd5NJzL7SSzku+kty69Ng9MP8et6aWqWh2PIu17Y9m
c7T5AQZRpdqTqBUzk5MSJQaO9l7028uPU0MjFMwHQ26zmgefOK0knrbkSrM7XYVD
m3AjTkFtZ6LXYkKfhsNf5Z5foAQR0w37NKA3SEtB5baxgDxJOZUnUDBEss4Gu51r
6qtEsWdvrMySLOa/BDBu2yMjgJqrb1zqeF+gx/rl0AN0jJ/pfutnF+8DMctJGSYK
8b32KepuvaaCHxYUqmpLPXw+cVEUn6sZokw0pwHE6MkhmNdQtM61Gdecz2pYq3TT
AIyCTvJLZB/4EGbU0ifHwgsYAoe50ggw8ytT63PkFVYBv8AvyrVa4d0I1WHpk7tD
AnbhLb7nIVTMHVh9BUwIev0TRc35b1Xp9xouLQk6Nj4FliaBOHEUOt8Z7UBB4T+h
gJPjN9/qLT8nl4A6MQ0gxgDVdk/wni3PLvYNS9yDK8YpOP9yqW3IiXwjABh/m1w7
tbQgj5HbDgvWCZq8Y7bZp6+HKeIcfVSiUQOFe89zR7AvIInN+s+TNi025MJPMDmZ
oq2wCQWDmXOyaD+YJS6Ilt0eXTh0xDtgqk1i5ojA7WHOdr0egF8623mBEEcg6DSt
IA5Qrkqog2JIEb5YwaVxdxNuYJUywvmQIg5tYylZZFEs3ima2paJ9iI9zdmZYLlh
opgi2yvt7coTUWBKD8U+1yMzte9j4QjsevzBjxPhP0adQov+QTbif74urEECurKd
t4aMu+MO5nXDldLWCFEiMfhcAnIpBnyMS5oW6VUfbfRRORPIzfHpDYKwidaqZ809
rZ3jaaF7jTT+v+3PIrU3iBeiu0+ViTJtXMOWzGLEEQQrfscOqkoUcRzW1p9zgvHG
Z/YAyc581KLbkieVjIXHKSD0P7oUvQkW3/qS3vrIIGBRCut2kE7bmbCIeGuXdyNq
d+6HWm9183CtoN43esg1jg0DZF/BZzG2O6Y/RU09UPqhbLSJk29HvuG8itZ4Guya
QfLp3bAUoOegnkK79Ce0hbUxoLa6S3DrR1jkJ4MUe/YGPs2aq33FOsvJNHu+ammF
LSt2oV+60ZT1b7rHQ/1lexPrYV7RoyMku1/2n9aNIIROHhMs7lVb6xItLSB1PRaD
xx4fxSR5TO9cy7p7Mt4gH1MKqARzn2ytmZBzmnehIlVIB/1F/zgz0Nv/n2IPahfu
wpWuFf7PAlmbrl3TQvpwv8Q1Pu+i96YoBOTAKrZHzG7szg7lBy7Z1SeA3D0lWWDy
QviTmna6t4WbEkAoovrKsMrO4S9V2mzfFOpS9sW8iqCiUmM6u+wPo9Woo6UQ9OzN
8bt44BpYZgwOfiQgXHkr3LsMMXZKTd09jumottPtAV6EbmZcjlcYzxwh8Qb6/nKD
mIfvO0J50rTfoeEiXmU1oSSknDNyewLTMzMUSsVbxq1vZKt1QQqpTQOjbzsIJISQ
mtX89z7Z5F86jcjYqGLcpjCdYX/y5v70iiX0Ov1M2Rp3LpTTiJ9GUl4RfXGHVt05
NuogMGQt22ua0sN5NnVtTouZnx/6NG4fSsloZNmEHk4=
`protect END_PROTECTED
