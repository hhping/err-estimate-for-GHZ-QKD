`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0KWjtJqL5SlW2nB4jljyKQtryWbLlV0xk56HT16d1gM8wLKo10XB69a4Vxd8lrU
ni4UNLFx0MuZRG/GGF8mq/fd2o3C42GCaiDzneK9I89d5naAVNENrsuJjgEjahL+
+aAcCsOcfU5de1j2LpsrNBF9U/GtNBhr6LKN/k1l1C9dmgw/XeMQcdC/k6hzElvJ
tYyQJ7nKCxfiFN5QEcdcsEhGnlAAK8oh3R7UAHPJsAs+HETWLXNd1H08z1KBc2Yc
gdj0JWCCMkO4bzlWIUdRBNxQS6+DNrSB/Vv9xadagBp4cw6SbSY9wjXBvAcLWfzi
zANugt1GurhQNKfIF+gr53WIMun/EFrP0sEOe5X4v8PVvfP46eFd1icIwZC6qZhq
sjGtc67b16znWRKOpxIQWlpzCiKd8K64HCog8Ela0/i2shIthEGAsO5LbCEIfbz9
rw9Ut25vd3ZzOkS1YKugW11uvKcoqvGN1w6AUy7Qp9FLhHY8Op69pK4NYVtEYj41
ouFhpR66NOol8zCuB7mThuuUxh+zvOZXN+vJ/8rGZrNUmil9R8FIk6pN177m/2Q4
OCR8MrAXDN+CQJADpfoQoJGCZ2czGCaAFdYFpWKbnimY4XNSFgE1I3izDQ9XOZN2
n1jfg/7LBa5iyCgN7Bk7FQovWJQ7G02DOEykkN5uRE0GAZd3z4YeDjyu2nPeceA1
uTiehioySlO2nWR/JUx3XN3TuN98BhOFdffG/JrxwlN5RcxM89ZeHcJBe5YaKQqe
Aa2d4P1yhiaSrU71XkvlTUNHoakS7c+akKEgMACLtgkWewSfHqy+pffhiQKJydeA
0IrH4vVVY8TQ34KdyYin6LV4WzRKyAPQ8Fw0KzF/50RJZ/OUmhZUovL5nN+BJKVk
xnqFk/qblKB0xO9rd8B5flMXbmy/nfqA244Xd7XhFnpvDvkNJum9T1AYRV7EwPaB
13v+2ZY8Fmdxrt+z3ETIAbN08IhhM2NhC6qyYP0FawZBhmUM8oo5M9EVHgQGS174
0y8c6Q1LWgbltcNU0kYtRa4Qq0ocYxdMIiakwAUHixgumRMS8FyUgAnXQlAAJZKv
z9X8dtpnDvKQXnc8vGJMeL/x85SOhN/RewC6N8rW3Oxa/JHY5NGw3P8+BKNSw1u4
wULc43dVD/3U35tnAujfaSZdfmozEYYqezvIn0AH2Xh0GvrEcp+3t0PiuO1lSEec
ruuf2eKTjjMa3QNl4+kCXtbq7S4+Qs+ZqrOxstRd3040/OOSqygLCbwxcwQmRHKZ
PC3FR1p5nalSq4jJ90BsEAhAmY51ZCUhGPFpuQDzKVEUgacuQ075n8alcqUISOCz
`protect END_PROTECTED
