`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XIrkH3pIuAWi/q6h81HpdexKVoqQXnlA5y+cQptA8XeHoXEOkQd3jsZ0qprCgGAH
6tgNFK6AURCSLPJe6pIdJRwYaZ6sptq2bXrerQqWUimyplFztK4bnJv+RDnw9w8G
rFtILjdIlIS+4T4Qt/gF50NrFmvNOdf//cAavTea6pTq/I5fynMXZOcDGHEJSRca
EIoNKhra7XcSe3tmLu0pE9WPQauJKST3OoroHNw7I2b4eo9H/hiZXKsDGAKaukTT
cQdDjugND8i/NKagfi80qh5u2tL5lxCT+CHX7A2lFj8k3HYg0pggdfXkpTtinSgE
IpF2FxI41bjlthZvjv2iurlymCPIKR7das/qqwuzxf3rncHvcWqhDrhWRn5E/zW1
6W3ApQIASFfaHqIbzcAO9z9ZjBJ40O53uG+XaqVnDrqcdM88pj7sP/I7YkTtMKeo
9YQIrMGMcZu+WOKe4wNEG+kQpSL2iRpa9X2GRqePq6zUILg9WnMijaP0KyVJ90Ct
Krtv2OiGl5XgHwkuZWYEswzdEshpuqCOxuHPO17EORJn/96ZUAnjZ5Cnu8cP7TSa
`protect END_PROTECTED
