`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkjh3B90yqNKHonCnXbgBYzCHaGTPqP1fbFNBDSNbwyHP9wtE5sMueR6UwepChNR
Dw6wCcD80TbbeuRwDi7fKK50mzNpJKMA04FGV2sZcBZaU27VI62mgkqr+vpTHPmb
q9ty3Mtt1bR5KYjxi3vi0O4AKXjyqQFnV7OH1Hqf7w2NUtbSu0TvbScctXGj6Z83
/3Pmnq9kQLwDFMyffpCjz2NJpLh/T+j9+WiE9THrokWqkM7QEqnT31bf4ph3dYi2
LMOjH8F3/OiSV0mk0M78zdrNRZuMwgeDoHerVpBMLgeuzazVTd8RhTm5FJLOTCyt
3MatQs4uN1IG73yAehn+Fp7X64BI5t9I5dak3Uw19h7zYsSW2N13ZpTHqnYiv34v
d1YWRjKHPMj81UUnTD8Wl+DhxEK0FVEJBBK0I8nXXhTrPJlMn5C+bsdjmSAZWNet
VC+UdtGZpdgmwe1LbFlv5qIiV6gttlWK/gNaOpbxRs3/hJ+XxLJoOkhNRRhYaJum
xUKySC6SJeG0CKIKHbrjHOhofkMzBEpol268ErKbQFpBTBfT1LXf3kgxvxaXkFb4
sVeqrbcjl2Ous6ZYqbMhCj1e6BqIBA59sSvD5QHdZe+4Nrmn5c8Q6l5x9E4Eb9/b
rBB8T/9BcJf0Rb2LsSNQahF6gqhVmZnq2Mu5QBseRZTEwSO11Wlr73XjTCFOwUBc
9isN7w/uc6VxeOsnjhREzO6qCmhb+84zH6K9ou/ZfFxWIIB/ht8zYC9/UzYn2cx0
0OrvBCyjjuTWgX84tGUFU9CVehbWRpqERFj3UF19ExgkDcCcarKa/9y0oJU4mf48
n7D9mzI2kLFYHCBvdh2aVrgnjrw6TqBKLQPYk+KwQOp/GsenMUbuE9RHmNSz/Vg8
+expZjdI0bRTgE42CvAOULUZ4+qxW+5eGZF6ds2VcvKTXZdvB/hLU9kSDz822Ifz
q6gqS//XaGg3flUzk2wnl35DqAyo8/B+/kMmEM59V69ggRC2CZ8uoFyVHcdJo9UX
j3SfbSNRCJGoj4CcxFS9BXUS7LrgDFbFPosHjM9lN70C8sXlLxZXnTD3KRovDrlJ
2RA2rcrJD8NuPj8LGOdqexUxkXr9+Ohg4mY55ZUSabd0NRzaqtyBD5gX1AdZvkdO
qfa8rsMy979yKIFx86RKPgvCeNikVsDQ9HmI1aTLyKPmh60ZFv9dKV3OVu38DuR+
lITbw7WKAOEg9Ge/hCWqzD95SACBCurNwOvrenG0Wv9GoV7prciEw+sObBM/x1Fr
Cb5ZPdciIYAwDQeCCOXp4cASIrZcj5SRfohAhkax0c4ZPDqSp+m3d9ivQAME6Spo
YvBfA8gRnMWAMipJM5uThA==
`protect END_PROTECTED
