`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SGg9kuUwLIaIH+4J7WkUhebcsStftBwI/CTqZ7WQuNZgUGDj49eTfnSyejZbaB8X
bHpLQLKu8uRMhLVUNepxxpwpJv/gq2VqGDl5P3g4L9lHHBfAji5/4k3Y8ZyFmE0r
SLmebMLEK0OZm9l+UMiGMZacpHETjuCvQTrxpd+zBlrN2sQQyyPyztGjThcketFi
bE0McD7y15TulY7s3UdQ8Jo0PD3SRp+Oi5TnveVcX7Ittzz9/A/zzJfgvrrI8dyr
5lYAK0e1x6xLmPp3L1GFXUQU2dV9Mku8RxRsSB9Xm02f0/tS3hT7wnPDe5AJcUEY
Vsk5GqmvkJGEpixGtqnDL+cxBP33fguN8uQMKjdeihOf2yLDlSe7ylPE5Gdo94+j
B2vyCtB417QLj+5ukfpTZLLaz0BVyidSvba4r+AoAqbrvW9nUrR6bZ36+o0ykrM5
ngG0H+BvlSFKrOFlcUjD4rm1VBrEDceTy1mP1v7ZxafoDcg82HBBOi+x1UgznZgJ
OT4nOVY4khKoL1ywvxOAwGm+u3sXnuriFdnDnIVJRo4hKS85jWwcFzRPdOTAscWM
LPASWS0iYpY10x159W4MjDmQtrYyyJ7EQ4eq/jw63g6mULNeOsnNq4gJM+JWgRJs
MkLnvy2uWq1b2tCjoUtdgr+MPQj/HrZRT6nHdvdl4CowEmnezTl0DeMMTXMicYHv
zLM3E7yPMdeG9WYeLgenMAwTP3Wx2WLfkS0lvcEI+ALdxD5phJDGpKxYKdaNleyD
bGWbaAnM0qLUyTKs9HmaWHgcVmP95SZg1i+HEWWphK8/dRaY94EIBxEuoJ8dtMmj
efLU/kcW2q2m4cBckA+Vv4zA1e+CEx6ARnb0UV1oJ4rUBV62tdcAKbboUwXCvmrD
56vIcpV2xvgyuafpackSpTLWMonTu6HATphZCu1HSNFmoPItOwP9+yyfDB3bGJa5
VQNT7Ti0u16MuIfQo4df7LpeWyPi1egvVfiXXOS2L93KDM5XybcYwmp37VsTxLYB
yHfwiPYYRad3KjqoFneaDsIbsydG07EZHvs5w+PLYarMnzXvPb2n0QynflC1TPVc
UBE83m1kVgqJOCvQFjYPrPZ/upbgFK0svRClPXeVRF/1mghQJxj4Dj4ht63uVzN5
nrtTRxeesQCjrXtGdVKIUqDrXskOXQmXDdndY0PfGKFT7g8G1DzKUgIh5u4D0W80
3YVCxJ7qRXidrIShd0eXZ93oxplcInkGVj9BzHuSwUXZDy7dprwSg6gNWm1lDWhr
slloNsjhULlRHLGYkhorBRfPj8WNBFpS9kmP6RTNUEI9mmPrGRGeUOIFks4azHIP
7l7H//bfE+Ex5nx7oztsuvUyPFtt1KZ/zHLGRUi979tokqicGY8GlwVnKspZ2Zhh
XXkRugXNT5VF8VMDi97kxg7FJcnpfvXXIewwGkZ0aLY=
`protect END_PROTECTED
