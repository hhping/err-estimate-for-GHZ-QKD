`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VYvnDjUH1NZkew23x+vyPIhAhnNp+Z6gRKINpkjZQDt05I28TAH5v4ZZ0plDON5m
t3cxeVTuqWjGVfLuT80Xq1mbksD/6HYJsQ5OBua2+S84fgLrhgHLhBv294CJfLSA
o21evrXmjeYK3uAJMWkngpUrOARgEo+8S+B/efY62HbXcJ7Lke53P9+/xhRFHkQG
PeKgDcAhHGCrgosq5Y6vqHBnuAnpeo3J9ptUbuc0O7lv/gQfqt64maCEkHCy6lTN
tfbPhDU11gcDP15zrCOaf7zg+1DRiQYvwCxBenofX8QwbU05FPL/LJx+LV7pJhci
hFkvobK/Dq6lZuTgJrPXGeVYY/CR+mSWOAAWAg6TGNYo4VQFXW6iN1Czz4tNXcue
DcQL9UhLhxg4oRrtZNYKT3ze+mJ6h9RVla1Cgn3n9STug74rCFHugCZX9JUH2niF
nSanZ7JSWMdtl9EXr6UAGkLeINtHgxOn76k/1b/ECbyelwGjYMxNLSm9pfv2bVA1
7P/yxuO1AzP4gIB6eVEHKrD9NK5z2NUCgK7XwyiROeYATEVDZwkeczR7M3J0xjcj
KnmJer2NM34Zg96usntHHxXFoYsQ1rtBGO3mWwh7KK09HNhtTiWmCX59J+gAOTgA
Lq4sb3U7vTWDcJ9Ry2QfkMrZsoYrJ66/EyvLqD461YY2ZIVPi026eO3IcN7v9kvO
2/bk/jucsVz7Ka51pvGkDw/U4IHvRJQGB8aO5MBMluyJqWGgsWteYk+hqvfqb7O7
7GYZ1k4PoNs4LBD7HKS/Pokm1mziYokhMl1/O+0V5GQESAb5StLfS9TCIYROlsP5
t2Y9w66J95OudB+wOEZ/mFYtLCjzerwGhMq/V0iLMdQ1nH241GmmdbxP1vl2l57v
rlp87ls7AwVYruSFIlR7y9xmTW5vc2ZQaRxd7aHiSdWe8NkoHl3w5jj2dqcPS78p
rUXiTgct9GwTa7q6mtGhs39vaiXep9s0Tuhd2mZrdDrrSQnQhcFCpSX+df/zfC9S
Ch18yK+dI91Rox497NlrPZ/7bfph94ZCrwvVpqOWJo3raCPpw5ZgsGUpIepaykI0
W/t73cS4ItImRxeTX3idgPWRMToZQvoMmEE0poDeZ3f4F+KVxPhsTMgUn5PMjFjD
EiKKPsKNrwtW2Ms7lFcAL0d+Am8W6ZVVFWdpZGe/pq4jbVHiR8VjeSngv/NMt8ri
RhPmb22qLl1Nwy7TcYs6z/cbIQoikA9Jd/VOOlkTS++hT9tYRjn/rBwSJ8mv+p4Z
vrIIGnoObNNy7Pu4rytd9QZqwRc1S33H1GzS6veGtd1EM0C/+MaGdvGhIkkl32uk
tp1PAhxLSCKBni0cUe4BEzTRj+UCgXBDIItirY+uk7u5iBJGSU/z4AmK+61wlHtp
1gMkspH1rk/sGO3Y/0EfbtHyrrHY56bDhIHWcsNqCPiw/5ws75xBRZVuq8a9e47+
QKQeQv7b4JEXA/NTJphbmoBSwOMKIuKh4KPDn6yhwg8s8vd1JDJWGiP1FF/8ILK8
I2dtVUQsQS3BBe1E/sZe9GNUMs+C/nAVTq+UUfJVcaJu6NrwmNiTJeaGTu0cMaZ2
U5Y2VmCT1f8GAzd5ldBSaJT5AxZ//B/VgLeXHaqkpe3Mt88DQclsZTKx6LiMDmNq
zRHLCguZPuORcw0KAZ4VxZTDpaGw/8tGDDAajk2o6C+6Qu8U2MV2usODNrHKU6AC
8nVgD7BsevhTRN1gVoeKJPzKq37GBdmLWGuZ5rupdS+J7jfxWO2Lbk48DhG0VluO
eqJjRoDpUFAgR5g3U1IXdSv2PGoxIcF1yHy0yuM+O0WLWqg7nON/u5p+KV1mj5lb
Lf31zexw8k6j//8aKS68Ecmr3AizTaLBngSgM90CvBHYUy0NX9xWkiKNoSSWATjM
qNeTuDOr+9AonlXG4KED1tx8jlZ9aUR90WtsGu7me5rFKgx9f0Rup1/yVKTnkJL+
ZuVgqoLrrNcoLQJIlrm3HFpqUfieNDEgDAADxV+w8TD0b8KJihcp13EcMfZBr1MM
ZHub2+yGXYpLqRIfvWOm2P51oMur0fSXNHoB53HOy8//4bgIc7jgLYyPzlPSQn7/
2FI+n1/9sVEe66dPpu6g6GPMFtbAAlcEXqMlkY4pYq9w5hHWncs+UgHK2YNjLIfc
z02g10pgtVe9IPvu6o+aShIIZO1jRilCMfOEI8zYr9M1cqmLuUlSsSsatUGEyWOJ
rLkogRTcUMPdG3dYrKoBuGfwdZ25jWdFuRnI2wFdyqR82vxvv7s94pJof0aEwCZL
XjKElOUqjUWCX/+7ugBir9/gKO5WlAjJcUi2rpyJeh1kDXdeB/NEYxeLcafyTVPn
ZJ1LC2GZSlB0TmhIea5lhsu0hczCfV+Ne7a45X1C9xWzi2CShGTyDRbYqG0B1ncZ
ku8BVYotu8qQW+MTbrOzipqzs22J46VbOlRq7ueGWxOqgy8mPKLVTYxKbsajO6ui
HWyCCmmpxdRVcCAKJIXaq8VZNVXKiS+IPyysCsiVqY74rByc8QaL5dtdnaXea2ez
6pwZVAlBsjq7PXDRimvnDuuHcSI6z2tc3M1bgb0O9TsVm5CpgUjPcDyBye8rMp6x
g6yNWASJ6OoJ8j0K2/CjjlTO8+dWGesXewDYSz9onn5qf4xWI8Y1kNgOE/ufTsaf
cvV/IlgmncKaZV7cZfXJjPIpjpvS3xtMsYCXBhpIMq7gQbR00wINC7T/nrOJaVrh
QV1G9QWjMv4KNIot3a4BJtiIaHWe6nFZRto9EXdCRmF5sxjb8NEtL1OTpHfgN8a9
5T/NAt/JLF7aqIrpnYurB/sDINlNkVMHZ+Am22DXQYM+GHYkVVYCpVAiTlS370Nx
cIwgN3Ov8p5++/otEnlc5PQgSSMVP5CO4qpZ67RHW6M7IK6PN+HwsKVH7T47a21l
MRi6DFlvKy2BfJAbquoIvj5i7880J/6JvSntK/EYlBg1qkhH8ptl2x5pLSmVtuqp
XFrGQkLTCSnki/VkgOPRQcfyysHfaP3Lg5gzpoDL+FxrnEjn6dXwNUr36AtNXZa+
J3RVKma2ltdKv+J+QN6L3GJm9CJUPNeAO94tpgUfY5oIBCDp415iDEsNc/rF5dyr
ex0PKvv7gPG3bBnjqLhjff06BkeIPUHLIY9PrTZHX66VMeFZQW5gu00mFkX0vR5j
S4qK3tiKQtb3MOPtFsrbvu8A9QAeYG5LtC6gLIE++H26Alm5+89Gb+XbSKVuNi7C
xgjESw2lULPFJDs2p99JaQh9vuYiSUbdwN2/ohISej4r+Zvkr7jiC02JcfS/2szD
3OkFoagsSnSgiYN1KHeP7jLE3piDpkbgneZruRcOMmJLUR1hROhYZCN76/tCLKbY
e7MwCk2s7KigBtIDPUsgNgdai6lFUZKme2ZOSvxajmN9ekDMzc/fRB1gks6ZfRKT
bYCeRKhTusZoaoeeTPyqy1dZ0MsHjWfPCyNGHO4/qPYUaqJdpR/T0MPEoIJnOegr
cbOQhTQead5kqvBTuQt0T5hlytUQnxpBKurRl1Odqek+ul36rn5otPcOh5ybJs4u
ObRDxnP051z//C4CbopeZSIEjYC21IS1WT7moBCIs4iat31RAeEtgmUZLCvRJGzy
aIvmL9pqZCvGMsHphZGFok81XYuO88HLvZKGDo4pHKWCbjX26czMdvWIdWx0B7H+
wQSB+mvUySOLxIkLBr+MSpuXCWJDVmj6I3OcOZydnnTdGojVpZOmvH5Z9xFIzfSK
gFdpgFQbAX8Vp4PTR1KmDXSd8RU3cr6AeyL28Q/X/wDQd5xk7QWSAY6nWw29udoq
88YPaqXe1k4B3hVVcApdMjA4/wcA+DOo1IJRq3CQz/eBuah2FYbv0wMkyZSYMeup
pYyFEPthsGN0E7H/Za/XtrTXH4pZysp5iJp3hbJud5rn6+MpPEVz8u8pgwLoKt2v
F4t8kj9T+P4LIJd0Opusck5Li3zP6o//Bz9Ziv3fK8VpxQz+i2rHWM5qvs1nOqcw
Nz0nimziZYlIlkWu33a2GOfSjLW+tGvQtWHNFc5rKPFWg/sWTKkYgy1J397yUOW3
4S6Aj2E/OPFKVX3NBmcrq3+a2xMJrBZYb5jMr92CqJqIYRQ1wnOzvcu/oDh6VCcw
pK/lgncngPP/KQ2TEqT9gClFG++O0B+0krsVH2Wjou74dPuA100q9yTyRUfC6E3N
fb7TxFNwxsEdsZZZCzaqU7FP2NXJFnD0NaM440FWbobwxaUvRBveAruPYTFYpcov
lK8BGGWjFce+nhEl+maF+u69T/KK4H10VTQVZ2wy/w+NPT9DJlK2W6xzMVpdQWOF
RJhp2y0Pko+aqhlvJRUQN8jp+SBgROnX+AfskFLFmAy4DO+RB6YUxkd9le2qz36m
TqqeT6Yj1eW7X7/J5Q2jINTTtG5QaIUYKV3n9MDytp5pkYLMRQ8fWAT4qy8ACvA8
`protect END_PROTECTED
