`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0/rFdemoIqDFV1FlE564aktGB06EzvYQKuKM8jpPbzWmhxZus1rBEucBDkFNKfs
cZQXup9Q1BUV6/MaSI72LqD3b9W1PTmUzZO+2haB3cEzyT49rCxN/DZxScCT19hT
tSh837dMhhywuXFQtFOKhcicBYruJmNE59azVpg+kRgIiihG+ej5XCrzs3ejDzkd
vAWNy67hqXUfzWnAc23dMJoYVNm8Q/QbeucHrxdFpBWDvBPmkh63evhOu7R23q1R
DL8gfcy6NCqQh76GzymfQD4ch5mSXiyy8swNgLwTmCaTbMkcXcQhBLpO5SjHpIlB
21tYe21yFquU/r+qSZMs6AuWVZDEm01VjgHu2/eG1M4opWF7W2xIQKU+RRyi2PrA
eiFfSwVm4Wq0Z0jz/z6dWz3Mvfv+3Lf/uooEBmWTltdpp2iN/mVO6HgAF0Vb0dW1
Ll83Enlsnqh8F6WXb4WTfCyq+MwBTzI7ca8WEOXt9hISpkxTAUYybaqoSwpWNdI2
IXpcEZ/xRYO3+Kr3w9QK47wKTSE/MIOJKGp3+BrAIfM0zHXwsdL18l2CEUDwMQPw
LgPx/autIXAOyq8Fjys8wzp5Vg9cWIcBRdKeTFAp2EUvsatLGyeBQRlFaphPqhEF
eIC3tQzmDaCvrs+a2DyKLkXxmLL+ln2K9LKvKtKjNFnEEWGqf3Wyoudry5F0M3yd
T9ZwdbqwmzsZWT9E7cHX84S5uSJVFUzMODMSAr/PPvW0HcA+dpT3oBvMmqUCbTjU
AjKrzORzcaY6Ds3L7IhLqSBF2fp+8bm+i+OTo0R76Edx44NqQskL1nIbOjV6YULj
k7CoBkKqxrPn0uK1UMBw9XAkvE8D6Y+HU1SJlCBZxZciRHwFY8H7nvxWOM5odBVO
aordFemj5nuoYU/2yMAdDA079KoN/synl50HldxCFcb1vHdt8CqaSP2FWytF6eMw
Bl4uXFQzBt6gihWB6hA7nCi/xR/rXqdIJb83e3EffkjrFZO9+P9WtMwkn0MuzICK
KJyvBhhzfhyhfPwNQuwrxdDXMMY/hqSp7E+UUOdX9JIKE7fJDjXinZ4ll6q9MKRD
6W7GTxwLlAvaIEPmXYopScSt3t2041drsFgwcpeas9jaekRvXIi9RuQbe9Mj7+jr
/pFB5g++7YTEZ+95tBtB6bWS+nYoxu0boxNMo/yR1nY/iCpdOr88nAasXlR9gIwK
86VK5ysQdysld5aU44/2nwlpqocMNR7/cuQ2P0EprvzdW8o76Wtk8kC3U0QzCdR9
Pp/2dWhWmHg8WT4UAIqpYO+mqjDNK0zKKC0ieENEHHcmJGjyIrSCZypMj9E8PCty
O7rjOWd7jZ6xbAEp62rEJnZA/ZAwf9jmx0FC7DemFe+AMh4oi7sLuK/XfPswKHQE
YA0qQHFnrsRKASdAIFReAqLd6ULFbubWOjFCj3l6ArA=
`protect END_PROTECTED
