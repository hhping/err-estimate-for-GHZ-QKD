`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dh+l4u9cGsJYWBLHXJL8862/rEfHM/tqZLZx+zWk5Yw5xc5YWnvOdDWGSjkQUtZ3
9oy/d+52rFcXfcsyYdks5uZK6Wvae8fI10Zwd0JZPqnQUG6l82Ac2zSzdYRCNQMF
25OohH5jIcLr/vFJQ1w2D4KCTI7BDnRNK6sanQdnzhYLBrVnNa34O5kkYJ7hgwC+
3dffY1TwepccD1cu3ZgKd51DRbY4Blc38R0NXhkPCZJb56WY00RdI0BbazY3VDaL
69uJX7e2Rgcfc+eVvbPYTcggiF5/oNvJZIlCmIa1FsiVTKBo7xujEgvnFHopE8Bp
+c6PtiVMInT+NVCNLQqv7CckWYso7MqOpu8fZtop4pEqrD/jc3TLr4iXoIAn5bAt
5UneON7OiCPAaCCWlyb/m/127l/HxA2w5x+t6RnmRXlrX1G2B0WTVmUIT7DDkp44
rVGdsumpIT+ViN3W64rR5EO5Ukt071P5hdDQHadzfs5YYW2IrrTczMuMYU9No6+T
OkSqn1Sho5LfXTp2MvNP0985+LJGzQSLPoD0bZIhI8FqUafQ2OlmpQGLw6TCatoc
NFHh2D+YTwGQ2GA2ZrIxp3XIDBS4OuD4skrmy2JhS9rSic4/WaqLINe0FEqoH2Ct
WV4KUYUzGBOmcUGsTuS6jphRUQJxMO8mE7siHbSHSIh1bmBKmOFmj/K0gmau4ZJW
zeypJboXQK/GIsin4zdDulXlJMVUZHjMxsuM2GIB7qJQ9U5fmoI7rZvV5eFjqi6k
pKro1eF6TNJPAUKfwZCJPA1qNiibCBMUB9baG/lnquSBH1Pi2N7uMegXepoqNt2y
1N3PdeMGhKIc0GBtAQ1lG/gbkrbdNYTivcbP4janacsUBFissAE96V+g2lFg98tT
lxtlxdt2jaU0kRCDE5k859vWqsu0nERnTbV7ykW95BGNh76q+ERKw+6oBXoGZNFA
qF4RvSZ+8mFhRZZg+TxMMU8wRvEoRWW869043z2ydwoC1EvGHuBGTHc1gTmTngqc
2VGDLwTJrmIREiqecloiJ/yMqxpvXcJlXtF6RLzpZsvOsnsdTE0RHFyXozZBqchY
AXEV+uUyrsUaQL+tHvH1E0is8mi/c8DG721H5zOPopEmlaurg1SWA+hirX9judPq
ytpEFIX0ukci9yRTAiXNSD2X4e8KpQ0ZENLmKFdPiILYRWa3y76Kv+TU72XhGqih
dWpKcsUoppicoQicE4jJ9iDYfoKRlvgfVy0dlgN+7xri2shtuYjwG0o8BWKOwslB
A/5uJ94/aj6VAV4CbaMeug+K1yBVdYa1+RzszwXRrAMUxE+qtRv3wOrxwK6q20kS
KmbP0OOrn5wd0xzR5v7vsn6nFCH7C1DxowlNAXUe2zBOvcHaF6PfHY8HnSc8o3e3
BEDl0rjsIR/VprWotxdHRFc1WCtwWXGTL6NRZD7DMZLtq88jyOnK+fgcKfvt39AS
Y60D2JpWJkBQPsd/abJaG/ojVbejO49Gzne0FVRW6lsMNUIk11JQhumVx05jsn7i
w24xR7aQl39ZYu5fO9z2wbsKyEhCs+YoHpoVb7Lqdu6KtuJFAOzeEo4LS8X/2qC1
aApOsOB5dl+SpVLzMRGhCX+sOZ4MPiYkfFDVFup2+CGBeOnhrCEZppt02GGil2xa
5c2mj3XJPm30bFes6hyv/ZL1MNARkvg+iG/qZYW0R8hLQceKmXH+TfCXEPe/PjqQ
lQ1qncTEfH+PTFKaJx6Rj5OTZE0TamyrVeXUJJmbRMPgvWGFFvypuPnLQi/h5Q0u
h4vGMFYORWYz4H0rpWnpzQsZ14wAKLYz3c5oO7hzhj1qQdiy/7nuKV6l2ElSujCP
I5MI0LFqCoGRStqqYv2h9Qn2htMDzPIih9EGkhsnCuUbwKMUcWJoBjH2lRvbOFjj
JDwdO9GXkxN77cIszWEtC2EktYCXnoxskKsXV9fy4OizLK4lUYjFhyJB6EKEroyW
kc5vCdx2flj2Zb8qiHVDKBPFu7nni8UkrNJ6tctK1vig+ED/7eg8PrWkPQoFAIab
NR2hhSsoo3jnCVTYDajpt4MmS4h+0iRG0I5JUEyNwKf5wvn7dGbgvMMH/ZE+i6Ba
b/yw2HqyT0rKtpeBFyGCNMc45Q1eiTzmCMEUG0dXqYT+aIcXSnwpCK0czxC9b2H9
EH7EpwtkblRMGKzwx0+RWkUyPOGFWTQvpVJmnIXP5AbzCCXUVoS+l94mw4D0ioJf
4IgVyLpSBtchjSIIVJVZX3Un6vQs34azNyuh3rZz2syE6y4jFkrTiFhCePiv+y8W
z8F9saXbt12ienzRgJWqmtlFgD1CT08qhjKqp13a5oRCiziRuuQzjckAv/EYtgo5
5+QuTpZTGyUAUQZ6frnoBiA8rgJqWu6qZ1r6Nzvz3OVkTmPYdo4/kOSZFrEsZPj1
R3aho9ok8nBld0uRin8CIW1G57YaobBpfwcFsAtm6/NII3QiCta4LUZI27ILMQpK
F+1XOzQTur+YYVHA0UFRT0vOKlvV1cS2L8oeRYq8D3g6Gjb98Gz8mzgbdFt3/+tP
qnPE6h975aone5KmQcmF4zB0cXu9nYx70A0vMNBZqQg/3+5CIYaQrRZjo3NP41Ik
a2j3k0Gi2Fwy5x5FgVEHasftZ6hQWSrAglJ/A/zFLY2N5KjKhnDAnAugilPPnO7Y
cj2/c6aFdYxYDgA0WG0mxLJimBDRK77eNPJAM4fClGDW9dwLacCFuaNTYrUbF0Bh
hejbeM6W9b0abNf91n8DLADH4QdihEpkLsIkGnhrkIib15a5CVrz23L+VZ5t8zvW
uckNW6kBCcDryS/hPHHNvqG04VPh1e32xcy+jErV6ai/lFN03Lt1gFmiKuRIagwn
fwEQ+ipcNsDcrBAwersaT/5UFkvXRs2SnADAHzSN4YT5WANpL9R3Jofvv3rO8+Im
63wns2ZEgRhVikVhOeFOzpb3rCr+BbEnS9ydO+evJcnbBqR6QpCWDaSu3PlU09GJ
Z5UJoUKZIHfFtjgZDWXlT/KMVcbHEBPQcRBs6DLeSM8N7ENJNO+gnEOr3xQxUQnl
/Y0F+/WFK4gtqh0TSXKmn/tityD8uWSO7jpp7zdXJJIUYfXUPkmid8D5qRyIn02C
xUXmo+O6Ib/wwwOujRzHyh7kYx4D4FSYybbolVMY6mE+UvIXrd9lfZHqHTd0IBDy
gNwVU+7p6s02Qxpb9wDpeJCDcRawNdYt89RfzUDe1XT4pWVnN7Xu2Zxdn/0/pfKR
QZqSR09+BZMZYK3c0RVc3eB8apwD97p96jQfDR7PuhOISXGNwx592P+/SduytjPc
QrFWziob2FrxKqZBhcaU3ekBtyGPCO7MIkAqQMyOR1BkuNJL1gzBQSfRQecY7XVE
84kZtvoax0h73O0sxN4kF/tFMy78GSq89gCNMc9VeS7hBmYkQneyA71rz8JNuC/6
nnHrkSAaxMcyNc7slXrekJ49bz1HkctLLyEhDK89LL3+dTV/2Qp1CGUFk/evTRgO
4Dr3oYD5VlImJCD1QH0w/AMDxYBgq2EsmnHcxIq2/nofAu8G6aFJ6pYyFKG6Zwvb
c3nIg3eGrRoWr+kocSMI66EfgFGWrKBmT2LCxJyCsiyJq7zOQXna6ZK9kFOOqdNG
4h4/gIti9tgATTgpReQv6XutFwJ4CbQDXeNmem8V8nuEb5uXp8lJuyJm6mocUokE
RuFWcyNGKWiemjEN4IB2SUbjNsTPlZQ1Ib9rrKv8BqnhjyuetMOADqJ7fjX6Vmcg
VBCx3fksnfiQrxH+u+6NvhXPDR/LNH8XMhNjU2/vPzwqKmh/HVRkgn2gtycpbuJr
jR1p9VnC1Gb+sgB88qINp1yk3P3dJuXncpAzu4Bw1+w9rEekKO7UQy1mzU78BhN2
Lu0uIkrrhdX8h3xaVnRcG1EjtD1H86GuCuv/4vx/bGfvUt/zRpnhleJRkvq28z3y
Jf0RuPwuhgKg8WW0xTK9qcAb18YUrAiKMe4A9RIfPzoWTmiFymzzSHYHmwB0m9ZR
TAphjOgshpBFFnurCNQVP5hMSbxnd+oLnCf+nxBElLAzJvlK8Naqm7lX+hXDLgYx
U3Ucud0gTj+BnhkvohZof2AfGVijZ+JkmhetpZLJjs8CxA39FGtuu+i7bBWgjCO8
JV8Omz0zeGjbLS9aN9Qh4hiyN4qEkgLqEpWwF20u3/O/QO6odkXRlCI3K0z6MzWY
RMi4G0zWABXLnWZzMrUI1yatev81EfTl3QoPCboXzdhJ0+aiKVXHIpJUJcxyxuKp
LTNlcWsYxHsXJj8uFkLuqq3renrbonQ8rkjCzycNTlNuEgO8GXH15f/PgYQRKU0y
AxX6SIZIFOhnCde67DVnXm/fQHqsDwG0yOVvU47hK87Qa7UYgyadctGqZMTVY8ti
FZrEJpnkVmy1EijDL9kXuzRJCTVwzAVNCiw4H6/KL5gOiw+GOamS3l41yiIZNpiV
RkI71wNkmNSePaCwoOEpugqR5KfPsDmh1s3fw7E3sjkIa96k6hq6jJIUHSe9KlPJ
tecuAey9+opmEcz0S7eG/3b4GRwgJqCD7EGorq93z/vaTqvKfR0qDR0obDHqYqDh
ejzVMRdr/4KqXQsxmqBue6QC2FCD9ONKs8ubVcytxg/PHaAzHmmK24IYCLAPWuo9
Uveqkv4Qfv6Mm8TjpViX2zCaLablafiVGIeALDT4GQlhOj/CkWSJq0uRNAgk7HLV
UbvuXM8G3cj6ETSBeAVVpDD2WQrNruYZMFe9XtSBBoyaeKWA/c1ytDsCI3QTNmpt
VX9DXHDfpHMZSKVpeMrBmP/KV2d+YFwHz1bNovBModnEn2JPw7u0pAE4DRCM19ZM
vM+36ADn22KUXfZe+9XDThB5JDtyY1ewPEjDrGoLS80AOU2iUShVE1J7TJPMjIIW
Ipc7JaLQ5XfrCGLEEeRgBArOhvjqNFyzPOMjIhm1xymKo5LFnJj4TjiPOBUgXDjf
9cRguyoQ7DsiFrrn++TqA6ipl8FUhczup31wBKCxXBEaYcBU/Vn1kZA2xmicNrFe
VGCqHqpvUZyCqP0j34Gr8SV0KoV1rcGbt6c6pMAOuBQVrrqJsmgfpFkJ0WFY1LzR
OWkA8Sceix/F8VWaXfAw5snW+5y9yM8qmsIdY75kDjuksin/gaGDQoOTTyIgre9k
5wvdxP8fr0oMbujDEXiTW1Rz3XlgQWDAnkktlUhxINL+DRZTtPF4vmQuKWKu/Tgc
Uf2HBhelyoZvo47DBSOVrNTH5HcTSxTrJbNNhtIXwJs/do0B38roAjCkYSIno1v1
kxqo/y7Mb+05KA+Z92ywKkUPVMXSxh59AUq119auZqZbO66cAueKrrI31ZaaAP0j
d38iZQjIwLIpyORnc7Z4Iya9YxHTZmeEJWsYaGNfLX0EG6QAwsuhomU7ny+h66Ua
Q/xsQXX0LW361kaaYEgfbsJ9pWYZ/MhJDLz0bQj5aVgSeoWPH/qWdVubZdfzf9FY
NKrCxu5OUnea9+F8gw3KnLKTmSiD8EiABWHJmfmxtSLiUFphMUEwhfubEXaAnXdL
B0UJFg6bWstTczHBQ89xuj+mSBPLDvtRIHP2vJsmDJhDWpIwDd9fwG9PyS67IFE7
nD+9Avg1ol/7SkBNLPhOTayZBnbWu1DxAm3/4sRSTI45aPxLGGhT5j0mwZrENxz3
jbs2HwoxS38JGR7HJAMNfXAo/YOhAbwQPB7hOpzhD3nwsFiyHamp2hqFUomYurK3
ekTn9mFeuP/2eIggAyD3wStiWadVSmZLOY4gpNjLu73BHebNzRy61Gt7f0sqKDP8
xLUQAp3QciRKSdIjZoAFhgLMz5i9GtNftgZLDNTQW3hslFX+ZeVfSUyE1vLB5Ak2
Uxki8AegCwh2fDabs0Q2xB1yn2JsDUpey2JpCjIC205r/BGxfhJH4er7v6yklayG
ZZ9IOrlaWUXch1HBuHE6WnlbRjF0cULqHKwLYCvy0/iA08AXrX7HdLRDvqGDg8Dt
JcLxke667EuGFKWtrqqTmZNll8oqASFGEzswrx7Rc1hbWzvx4SDGXg7h8MNI5z8+
le2xJFN4t/+AW+6dZD4KS7r7/0bCtkrgAJgQAPFoQthqnWQBrnXG15NFVNkZPd5M
b2UH1jPbBy5QQTAYuECkkosAoohz9+zXbOjeSHrTPfx14UU1mLsaHEzchlHUQxxf
obGCQTb8pN++D9k65EvbQqVisbJJoSNcZ19kAcdnXec81+5EnscITbqiTSUHpT2C
Yyg4tUaBbTgtpbzydVo8xK0Yh3O0XUFEZgAp4PxlkjRyQJO5Rt6JOOmM20Y3LqYg
TfHgZIFUa783tjpzCd3ZHoMqsp4k2p8I0UWfz4F7ka+2ENkl2KTS7ecnUQrPnbfO
Q43xtoE31A/N2+BqOh/U1IsxA+ATtsZYE0klfpGODA838gXjz28o/2Zcaewwj7Zb
fdQOqQ5BdEX7jJZq+U6Xfuq7tMp3ho18t2QwhsPpO57oPys+izbI0rs3h2hz+V17
t38YPFae8DXmpA4B9pbMShZJKvciFFX6FKWXbaxGF/XHLKqamw+EXmOSuheCWRHJ
zhsR+QQ+n7lux/Jkt2OWXzB2So09nI2epuiYgcOpyoaSgrHxKAvuOgHycYSe+8aG
W1gWdAadFSPz0skBsVR6pGf9w44/ngbD2lgXV72fxosW9PPw/oyuDAXBuTkUnTDf
iGPRFgV03Ak2H1YLKBbOsw==
`protect END_PROTECTED
