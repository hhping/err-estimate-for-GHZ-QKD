`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dLb3tjwE0E87jhPyZ8Z+GM0MxmEw7EfF3C9hfQI7xcCHVRjRZSLIrMSer2L76Bq
m8iU2D1vegs66C9GKM85FzQi5AVWaIXYKblrbpXaj+Mx5JJ7USQLmYt+F3E207gl
Q8AoH/7+insnYGgyQvgzdGRzn5X27PStJDkSIWN6ecQh0FoYYxqdm0SiSg8Z6wBJ
wU/gEx3xslGiXcklaNTycbqwXSGTbJrBulebU8Hfp0Fk3wHxrEkOxTnm2ayQp7Nh
hArPyaWn1XKiczLnlPFpQOOR5f/DgtA9obFAUNYvIB1dDu9RyQrKzl8CvcjfkI7Z
G9h244F2+qXE5o1926plNJlu4H3jXWKzVejq9WX+yZjhfhGWHaqqm8TqmVNMzAr6
kRUiLL+eI2CdgBaWRGY6xog5dXhOi93vISrkLwVgcw66ZaajwPToLIxPoGSU/S/s
CgyAhBtko3oSWitVXmLrep1tS8L44eftg9uduZX1NhWkp8RDIAQNRUgl/YNhcPal
k1RV3yMbWkFvYHt0DFN+DDfyrBvnqsX6ZWzhzh/KooIfywlUFr/uK0FRhNP1C5oE
yDyVb3PGbwYVLSYnrZ07UUl8uLGC6CpIzOsYB1cU7rxeH9kN9wJMmwy45w0PPYjg
RIE1msmtol/7d4T90BSAJrnEh4Rx16KEWKtjWiQ7+L2AxZpJjm9GZvTrtOc9tgcI
V8Cu1qbyVHfhtkt61H2yeJm+MeViVw1GZvHcxOfbwtz/p6erdfucK627mNwlchaL
oroF27Nhmmw16vmODD0kgCfl7u+OHUQfUX90u/IMBCDUExjxacz/DEXeZ1la8pba
l2D5Qcei12yjPgCP8w/0Q9iesmocjNqDPvxugtABCAnQmkT3Z7BDaZ7//7KUTfQ3
xo93hE5+UFGlqxuDOGcOAQbB6VsSbgSUGKrpD5OVya1Jbd8T4UFmHPLjLLBEcDDi
dExvEEYzuVEm2sPJ3vuz5RPI4oas9P0tv6uZv+E38kDBf0Ju3V/H2E/ghxwjwkz7
L7sdM9y3Dlx4AsdBnJjvqdEWSywTwyXAVa1igTT9VMB5wthiposoBwwgKWE4xxnH
YZkyh5N+xFWq7Dn6NBKLPTF5x7ByUGc+Zg4SahnfrNX6ThFTxXZBjzKLsBXetFU4
rfoFWKr/7+BkvyiB+QZnExO1MeliOJDPMrmF204sH/WcO4gOXml8wOHMEL0nIe0G
PuihGXZ88gABlNWhxtmWns2CRueSEmKshsMM+elxOLBI86k0OTy6RM9g/j0SS3XA
bPdGc5esmzUqCd7wVEJj5UasK3RpBPSvEy1vTb7P4wUCBWhtXifezBAspvaKQyIg
fo7iouuRBLMP+i0o35WcqLNuMt7tCTt3s6yq4LYFSxt0aoQyRwIORvoJQyXuluzA
Qm8Dus43lkuvtF6jX1LPOpFJqumkLSBiBja/cd8RvjHaFZEQs01I4ogSDaWskRjE
NSviyldIx79A78U1NVazfmAdNicTH6U8tVahE4kZIuGubYZ210VD1VSOnhBPxfcJ
yFbEacvoIYMTDrRzrzeBl1woHDiDiLSN+GCKXJmJ9/zR9Kw/19g62hJAa2WpZbAv
b4LZOveH1E9dcJPDiMIP+qdNDPXXsKf6eMB/XuhmQrx3zTm1SHUwig7sczeApD0T
YPSmp+IyBHzGtz1SWfxtxrhUs2pT4R5fDLyeMp0llvCNERal/VE91N5tcCb6viD6
VKtBYA0ya4qbKJ9dHdFoLRJ6uXTA2ogxxnaBNwNH439N8HILwaZjGAavuZord8E/
OrEX9V6fhe1+bjTqw0oQDnlXji39myI5R5o/zTaB57K+ns4NkHWOcg0zlc/PvpJn
/I0KF3F2itn1Ei+HufOBG0Djc/XP85HoabUcQ2REiFSk1JhBPqafR16t4RhomYd7
FcEWyqTWVMKu+nGQMbuIEe3n/5zYdIGloZGF6POngzeNeNUYdEXskHclw1hA1/7Z
yL2sKiYIaGa8eZJX72a/sAPF357zrgSWS9fyyLEtnlRCCTP6yHpWXy0frYMl5fmx
JbkB2qyLTHyqBmYWl8LiMKdJaZDHhsVOFzK55RNYB9QtDEQt+TURPCii6tbUx3XI
+ePBurRUqjDRIZ8v1Kw4VfSZP/ttEgg08Cci5sL2ekU=
`protect END_PROTECTED
