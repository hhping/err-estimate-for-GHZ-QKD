`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/a4nP3xDEj5Rh5WSR8XnVFt1PgnXVVb2S6NcqQ/7Qv5tQPZKzDRs+oM/F0f9AO+
nuCDf9o3W0dN/7QGs4MZRJ8qo8TCTOXh8PnQK6LmXb0plg2pnu64sy8c/TtePdsU
+P1k7LcP3ZNVMT4Y0zCusFddOVgO2Kz8WnKhT8klDv73FXnBUY5wNi5c3ig9YCio
4tO/ZJxkZFRWn7T0JP8feXjSJxuXMGLOJ98vsO3U4Yxgd+5P6jbGALON9jQytciF
KxVzA/+oImU/eua/mRbVcfZRhlkkf8NP0HmfGTN/UJLjR7DD111Xx3LrgkIhDwtU
EnNNrS9C1fwEYr1IyXbyJYd/VE9do89jCkW58IgaxjGRuWKEjCz4Kv7qxURFZbP8
lLrgszjNhu1G4/uuBq/NY2lfXWggciTWz8UC+8Js70gg3/XnAEFAyb92dIiz3Rv8
n+UZYikdseAQeTxZNZU8TUUXTj64Ahlr+rZQT9DDtw+/eR5PD+tPUs51FfGoPHeZ
FTZwK0EmGi5fuwx0a445VjiTi7md/UOorudqfq90dwogM8mqBuH8pc0u4U0aXaC1
RVejwBLYPFHKAuSvstQObh0IQ2c/urg54cp0AbizokB8zHpwwNDVGXYV9zWaR/H3
dmA/rbEWoxYpMBfLvQ5PCXsRqCCBufzE0MKcQPtTq8OmhrtRbTFCQjpGQQ0HwLeg
Mhi0oJizWWipEXLidXP1UhpdVNVxDtU/lfjJnRmxvkDXX8h5R0MbQZkCsMeJBWOK
2Snbi0HJ9yThyBwoXqpfex+78YZrSiR9YKzoOn9RJhF9T6YVzG5KqkrjwgCoYXCy
blZ4bzK9j/+hryawTVHQ8A==
`protect END_PROTECTED
