`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RvWZz2EXD4IwUqftqBcs/r0BGMashNTONVKxabintX9NoP6GxRLQM8+rZ2SkWULX
NcU1BFhAzVamdwOU+2wlaRpKG2uyX//sBASIEK3NjHHx1EyU8E5G495iMT8xuseM
ydc7V8qzNyskBQfkrGwUVNQSiyy8GBM1hMS2EuqiTjaVEYYgFHv/NqbytBQkX2IM
98v2awSycOaij1Cwcsa1jXG8EeY7Bw1+WwRkzRF46aclO2rM10yu7ZC7qdkj/NPF
Z7wL+uPuaPlDHP370Ua34qShTh1Mh1IfTur98mWt9wI5ymyyD6RdTp9mU+UVi/FG
0KOQ3/ECxVjy7sobGWRUjNheqt9EsunMWCSBqbbwtjKqxMqfNGd+xH/FBk3Bdxq5
lMzkamsgC1QYkt8lDhDXyzgxzYgOIzZRZDD7CZdLGvFEWtLEnOhfzRpcNIlkIOul
GqItR43xuW26InxGDDgKbPqdj87MNj8GRaZmi+6I/rEb0EdqwadXC0wLEE1fenrW
TUmGp6I5dfXfr89lhBFPEDJcaRfNQ/e/RjR3mi8EdXwDU5DHETSDWN7kGg9rgShC
uFXOCWYUmeOnTo76z3g0jGx6Od2/oJyY+rfNTbN4qWMMiuMDi3B7MdAc3kIr1SJS
2KrLume3V3fKPF2kClZ0Z/16ALOiMjNqrYMmjELsQH+GrFrHZBJP4vgNCHJiFBWN
VAaoaOMPJcyG90PIAGHxsi3593jE5v9Jkrn/lkPXPQVEFEvHa4SQY1UcmBfeK4cx
NgmB956qsyuUm4lo//XbeJZaV1wOAY9CF4paQv6sImAUBlQTZ/NOQtKxTyCtvB2I
qiTcW6tzZ1WsiaMnwGVYC3awie8KaC1udQ8qM5+2VMIMiunJdlIbFBSa//m0+ttQ
bKDcKJx42V33N/7GRgL1EVG9Cg9W+s1On+U+1BxKkPW4PqQIqj7p2VeXcY1LZJ+x
rPTPfDOyc8kn8QCMkTn5Izkw1BHtDZqrF8RsYKqyKZ2d6nqO9d4Fkcomt4TrPaer
e1nz8wnytdRN7a7jCkFk8PqPyH/aas7cR62swra8DZcIQ/kk3PwOrIwGEQLSuBFc
KuIFxNn7tCN2nLKLLL2LX7jR9G5KAY0d0DcuZZ3EoRFVgREFEC+HESpv5bgd12dC
5SEJhiP0+jwIMH0Hp8m/zqQMU+qp0nBNFE998NRIp5qptOvzcb7r9JN2ULPDZXjS
KRBeoDvmSiFmS740pX41TuO3okJs1k+sC1pBhua4mNcAf3Cjsj+AtuwgIfDTT0zG
4nJEqg+Jt6/pD7xAGY3fO9HS+1/IAiIViLrdXqTvMMCEFYO/or9a5XCQbkHUizmN
WEDo6cEbf44gIeSYNLlBsouz+f5/XvjvqnUvGdOmwzTX6sOrkIBbRFwNjJoInEuO
tT8vWcqj6SAzJcsDU0JmigodPU/ty4MErEbsMSY1g5Xp/uOAjMwMDVnBapB8EGVa
J/mrNIajj6za733OY7V8tWpY6x5FGdb6ySkgeWGtyJR9VyVdAMpHXfSNXS9XacHR
PoUS2IDdYa7n5cPF0R515CraC+7H/dFrkk+Us4X9w6ko36CFiOU0iy9Q2R5hg/Z7
gf5FvRrD8NLqyCNKu2nang6xW0fUqleTDpi6cJFJ7RBDRwvZ/ZuCgVVPR/0mObAM
JNodS+EL1Ppc7VVQTjP9UfcgsonvuL0pEjaHt7e/aOKgz5/9KtiMsAStO85VQX3C
U6P0f4yzhKDdB56dYEw4LB8tG3g7UqpEfK+H5oel0VauL7YKbSKQ1xfeE75Jgq2f
sxSNxnKp/KkcVFjoulOpEp6CLb7kNP6fsSfkTfCKGkg/M/0TOCwJNpzoLkvedSaq
7VpWY0B2aOMacQvx0DKTtJLoM+/hcbt4ZWPSNkttId6zxXj/KAIi4Htzgvf4OqSl
f0YpISAolMSY3Z32YiNnpI8mRWU+rswVfp1rUz+5w/DHUJwHSssaazkGFNFQfTM4
1WdzDDrqSrMtAyyawZV35XBKMFp6og8HXQUAslNpiJRFQWCtODS589jH983oRHiq
Rmgk3cOT88dhsKuvmxbE9Rlg8aXAc2qvmRq83q2HyR+LpZJVOAiLO+1iOk7qmFyZ
GYDHlacYaMXjitEkTOBR7qLfKqoCCcAFVvzU0RN0cjPIwXab7LaAxG/lumjpyIW2
BR6tBHtOIcve39/naTxl36DqaC4UTpgngD9JVwqqVAR2roeUnAJhbwbUhwAYxdOV
3bA3XKkRvtydk2q4NzEu7a/++oo4Zdk7FGl+htg1Ru1pB4aZ1bqXi50q5vGx4Xfd
ajv56HtnEIM9yKJwqEdRhyCJbhC0WT4HjB+AtfI92cUjlc1g4PVCQCVg+APOl0Cd
Iwuj7TDRZId3g8wS3Y7Bfa/vpNL06AgG+pqp++vq2PlsaYdB+rP280fQ80lbcR9N
pWBZbLZJ4/keOoXmfd8ZejDs6AfY24Zh/jiZyF0NM1hy1tFGlfrjDBFwBl+bea69
qAl8r1c3tk1Kl03hQKCPpj/xqh4nJG5OqwJhUcLDWR4o7JGaiHGb1CcvyEY1ciME
LpPu3xEZ8KIExen/Oul0diAmjfvtd89CowsXtibS0bHV6voU1C6iYe0fg4iYm+tm
l5q8YtG9LVJVCLbTY6ngiru9yI6YTnfhfXig1Mof2Rxoz4rgiFNTpPKUqVfBB/T7
2CELAxW327oNhDb/PBa41a+i+Ck7xjkzlBhS/GSggi5pKms0GNW9XmcE4dY4T/10
0hkel8hDQiq2A2wjhPw7uuYg9767URVGC72l+YGRoJ15PDvCah5jOijMJA9s6c7G
voIZU+/YiRsObiMS/Itoxg0sU1JZndsIp5AkFJaifyV2RrGJZGrRXvFaT0C3EoB2
ys21QFedsDBA3yRYdXUZm1gcUfbqcRuJQKlrubqFHktmFfGkC/MW7QT3V/fZwR3z
hGs82J7WuIFR3p3JuCZEX+WXJZRuIzIkexvX0Aq/aX2/pKgiDB2ewbtliq77ua1b
VbHvrWWm7r6ujXMJae2XuQNoESDMqYCorqkJkibMa4NSlrQycBazTWMQg0xuGPc0
YjHAH15T4f7+PYYa97Ewq9hSHLXJ3EOstug3wn7nqkbt8uuBfI2E6MZWLcqCPOyP
e1wjo58BrOuIc1JOCljtMvU8tApc8cJPh/d1baU4HstrESxd9/T7dHMF1oGQiCEj
EMwM296bqXhxagcOOr5HPWVRFGx6C4rGgs0/n6qPv6TVMTB8xv2rbijXXMv0FSTS
KIPir2jVthOYLqeQPAxtHtLY1KT8w4K4Z9n2npQU7k5p4ATl6+HtuVTVilrnFgal
hHcqdy3PxfmyytHwtJCuYTUZKLaDNRfeTid9EDR3tLC/vrXEsSF/TaoTR+tfi5kK
RqWZO6S8zXJtBV1IlwXvPGp8YEvX+9CVgbDDg8Yott8AvK7th97yVXBRNhv0eM1c
Bq5xAoRH+JQ4DKhrmdipQOfy7aVGB8fVb8UCbHQR4QUMW2iGxsprVIJ2h9C7zUs7
FN0bhXfhLrh+9BZhlr4W8p0x6tJPOsTc1z4UnsPzed/aNMAS4rKLULSsZKUHgD6v
0pUC7dHWBPZYeS7UBtixLIBK4jUzkq3hxZeQLOhmXRa3SpKDsYBF8m4UL+rIvF7V
wNXJz6hRem9SDUotEuliEiIOKQk/osRXjlz9h1M5xyC8R2qk7VfhYbg/g0C2QB3y
OHZd92/a2wZWL5PNhUVY3Ngv0WeY2mmji5LVuqf5POu1NQSwTvgNKSKcguzGNR+p
rHPfBQTU230thQrkcexZrp3Xv5zqogkY3/8lZYfxwgor5W8kfIvhqFp38awYTdah
0dELXfAJJwXmdkdm60XHW/McEYw3FwG2Xq4wZUWVrkS6STwnPWAaZRE9cHfg/xnj
39Arve6KnPeSNTs3FGOi1thtITjKg3yjQe7SW3BFoAk=
`protect END_PROTECTED
