`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWTjl0KX9oMnnb/woSqMp/1/tUZWQqlSC1yy3xOKGTZ75i2g6NvqEVO6E2v65B6L
P5p8rrjcRogsZ/z7PPJpKQh/tEhhYvH9IARNEYRpFvwBHe6EZ9WjHCrEXAwswXD7
AlwOuvTSzBolQlR1N97uMiZa1upKZEFiiZD8Tphj3Zi6qzhcsdkW2PPUKan3ywzs
91uew5LgaAfeMkaI0yzO8JpLc59Ht6XHH3ZfLdljvm3cwxX0KZPiKuc0z9zVEMgp
LHWli0QSD4KSuCHedkJg2088ZNUSlpzj3qRnxXQ4+qzHecmvFxUsLLKiuZc6IQw7
Sej6kkK2CUAX9nsZR4CB/Y/r13jvVwxDQcz5ki34sNVjMo4QxpjR4JzMgUdI5qJ2
gkBAXaQVyjRt96HJSNyr9bqa2PX9tGCyvKJX0BA+1LJ94ozAJaVp0NtA+PZbwGXL
idsLmejwxOIVipbq4bxlxrrrlkKC6BFJzYEvHtesddotueKN1OjrM30fqAQf8S5a
HB9Kvta473kgZjixyizQavacnMA1OOQLdTVlwoFvNeIrV0aMTyHhuLhANypjZRX0
ivIHhjhOx7Wg8imzybVIbKQl6oMQ2RdswUFMZ3oc2FjYubDWwpa/B0cFC+LZP2c3
bhxLim1qbBw+an7hMVditVxVwxW1VWZoOd/2UDc8siS4fBhC2ZGAq6dziaY+XrEm
2CwcZLTLDkxfqjP8aRr49g6pEZFCe3E/1KAPBYi2OX6L3hA0yfzFiI+zTYOByVSh
cK+A6LVib+0O+B2xfcKYbij2dEew0V1Gf3lbk7hOzFkJzlz2P66Y8/RQIWRnUz4D
9AKLJ2COWhwXMFH7wc18fkp0ximsWeRmuYpV2fkHMJItDaNvhsxJYQsYbJdri4Nr
TrJyNR6vEtlJncSUz3zZaK81zfItnRSNzRT9uA8UXEe1ejY0LBtcQBlTJDWuyH+S
XfSjpH6zA6q1ApneAlKF7qQY80fX7OlJ/P/gFLz3tcRo836SNBQYMeQV7Xxxalwr
advwP1wAKUtCQRdA9rtdj868J2RacUqWeu66I3H42D9rQX9PFpI6A353ggLmCe08
kVizvcuNRN5tuZTIa0Twp5vKDxoN4/fYJFIOxIlJek9n+FsLshYyraRo/aifWA5n
xAzrfokLsgr94TzVm98JXNsirb2szTgqoQm3LoKY9NGhrESvmccqAHRB1/mU18y0
bFLXCkRSET36lcNr8swaqIoWgTf0Dq8x7OAEktmgOiunIuKgxgVER91W8+kyLiOM
slezMBzKrOnf4RTnJFZadE9iRF28bNzPGQMLrVyOCGOFRdNIczAnpeijGM+jkT3J
cYXt/aBIjtNJDKbNKlmRVlNu2OeajSmznjFV34hbOqRO7/e1dwnGFGlWB67mGlPF
/3ePOd16f4zqWZDOsVSL6GZcXjJnQauwdJqd3oQrPfji0qCBoKHcKFBaOBSPvJqb
Xc+LoA4mtVaoDxNqvO/kN3uU6EgGqGeI93//ZYK1O8SkgE7zybQXqPgP+gKRtAUV
fgwuKudQlPXdndM5K6p/QjIMzdyCUxaSkKDJ3hzszYuipWIISj6Q+L1uBZva3tE0
EmyNRoK4nP/iAib8P99Ie2T9Wec1UX14v80xP06IscCYEuWF225pBc9rk/SGPhg+
F1gIZJjjVRHCCfFRRXovhoj52NKXM8y/Xwy+LuaoMn2DQcAAIdL2QZ0kekr8WghN
zoSyoWb7/Ea7dTOie3ASBb62nd145bBUkb3Yho5y99xis4KP4Dfx4S0SjripP2FT
l5msmkIJ1go+gyEaYvs/OpPiD0debTed5VOWFMMpaBlyIurLOYf7axbgKN2BW4Fa
kiUiobz7VGMsgVk62NpSbA+9+Khi304HypcDQ9uOdsPFQSCiMn6k8KVpPgtQY/yn
VqNWFVJuHgKa3eVicQax4704SNnXVotGOuJZXBV7JoyrXfHv0iKDyqAPWZ9tY7ka
4iYQ8OlGRRy6H70Hs+gaAVrXcPVuXOtIl0OPtXORdTA=
`protect END_PROTECTED
