`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oORVmtPVtZPOUaDWvdZddkAsqggUHFwk3+4f4nUXxGvfN8zSKcCDZO1MW6L22yTV
0I0WCKjVb5VjgJWWBFwQIfTR2oZcMksgDGaqRED9qLOkfrwwxhAzbkKbgDeur/vy
pGridqNa1Fy25kRwk+POQIVmWn8HG6j7Tmap8UlN/SvS4eAigGTj7HUmZaiA/ejL
PIMaH4LXtJv3pV+BspjWdRM5rI6+ui+5w8VFiM7PpSy5oV3pXPdc8D28dPM4QPlS
DTIyL2EkqJvCLAVe2e94RTcMlARfJeEwLJxARGqfSpvkHurrJZeeJlQfTNxDKtF/
zbJqOp29KK+RCpEcigolUXm3Em5LQlL79ETYE9u4sX8iRrsNNd8KGXZzRCN1fINp
E6/q9yvPweqgPCicku9cQtipmkq0RXdoxtQFZR1IN5vSn05PYYUw9kKE9ZyhYfCX
RvBGo0qzV1moYmzMOUAL8dvolhzzOUoyoO8Y7XfblYqLioU+We4DK8OQSxeB3pzO
vyj3euQEZOf4SvO6eIMQ4ET6CGhdh2NRFD6LHrkI6sdtOPJXF7h59Zb1hZCLH6CZ
U0MGwPPYXT6Fmq5Rw1zODvnA9s2Twfuh255pzD7OSaRddNoGCYEcu12LzhMue1oS
kiptlki07LFa7m9LCO8ogg==
`protect END_PROTECTED
