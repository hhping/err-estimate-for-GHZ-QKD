`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9X0K0xjgnHECjVU0t1BZ+syR6huotkm+WXli6EjbBltpEuo9cod+kNeBgp+zNLem
r7c6CnuJTUzV/5vjxsxTYUDp6G0BWURVNAVPO4xifcVJOe1XeFFgVlkRPySOFiFb
PuI2Ea+ogCq5W3DMpvrn5vWtSdsaasd0THN7Dost4Eo+lTW5r9zCWZ7wXThJA1YU
F28ZRX1ENM4nzYxxnYJq7Vjdw+nL5Ta3jdvFl8ZoVzgT72cn8vpH4OID8aVPCf/4
K9E6cpdXzg/zlU20BBNy6Y26qGzRzxcys/7n9euMoOCZEOurAVR+0Xk818t0O5f/
x7MqNq+DpUhYRtMnvJ8lQ47nzaIO5PwSE/mygTXa3mjNLkhApb/a9oczMA5j4ngK
VohwmDMfrr7mR010c/LkOdxREQtrRB3QpT5isnbzEhoFD6Y5Rp6yo87KhIgnVH4h
kZPLmGMboPrd3p2aD5bZUAABsMYJe+VMMEs6O0+s/u7d9NFNS4tHZbE2McGAUPr8
2ytlOPElFxJiQRRMTpS8RsuDjPT6vFjDQclGSecpHYG1mjmqcXU3ImqFLHcv3t81
FJSSw6uyLSYDEqA6aa/CeWpKPEYKhw2JoIgZcqQmqSr3un8ygIhqcfZZf3NN0lUJ
EDlvZTWuB3U9C+4uBeNDZoL7U6Otj7LYnB0vSKOJPar7ZFV/avldp/kxq0WGMXn6
yEil1Ci65yE9npX0syAwMm3nvdsy40oz+fAyee/rFF9T3e9AybXcq9qmVBTzCHKR
wGx+rJiMmrhfLssVecRVP9ldC4J/mo4Kj8gaHwVvhc6fyKA4gkloNAOo65HEOe0q
6D2KURUbea+cn4PcEcmdWeb77W9kbtkuYv953bwq85CW98KorJIMaUgv6BxFQ4x7
geQ3Wj4fM1ZpAjTxO3EUWmDjj8ml/nK8zTsS6Jo3OWwksNgSZByYYDbhtlC7m8Nf
s3S44PtSPkWLF3rwkQpH7Dz59NHI7H6cKylf9c8gpSJojrWMkqoAO1tug9atCtEj
YQqHm72V1PccTpmaJ5UCV3ne94W4Q6NgA4bpuIjPKgRxBzJAx3oq4SQgVsLwky/w
F7WCKJHzErnedKmXB6pnl8pgtWi8+gpKPsD3EwWmYYDjGpGuqeRuhcJe1p+eZ7wr
WmtfIejjoMSbISXsarVNma4GwRnxpwrOTE8oTcgefYTt2pWN2ndiuNvfbyqL+Xwf
p0HNi8c/a6N9iQA+az0TlhsA+Bl+qEN3FcYMKUjBtuu621bbI9diCSWj0Yq4MFXS
RU/9efWR11CsowLEeDsa1XfjauUkmQ8WCF1aXcZPyw1uAJZJYHl1lsuroB/HwYAR
2bi7ZLZAI6y34tNFdnbpxBCEOQeuNp3Y8x6vsUuWjazTJ5/T1XyWZX7kuZgWm/s4
RTehLYjbG+H1WQq5zic5SPJ7tG/HgTp67AcmGYhzUqn1DbOgfTvvisA+ILavkoQ4
f0Bm2UeeG63z6YZSvhdfxdI40M9E6VjVTzG7HtawcjEUFhhzbouXaI43f8eTFKuc
oFxYOSKcaaaHCMqLClhRis0dugL6lBvQr+MIsMPO6A71WtlNSEo8jekBerTB6MWh
7XTMAcWTSKFHyoxJpLq/oZ8pUxMF2V760nHNlTGJ7iWFc+8qaTLVZhnvgnoVs6Tw
ACULQhHw9160R+bAAmH4ITQSR9MuJrAnmMGERJTxaxugJfHW3h9xHeFPJOJnA+Fp
wQW++ogj9fLRdNv8QjRPX+iEqJgp3gsN1afmS/ScwjtNGceh2VuIMigY0/3T8loW
dwFAYeUPUU35PurNMps6H29dOt/SRrp7nHjA8B1lQbrFauAlLocYivFRre25bLw0
efm3Le8d3P6PCZWbqAsi1Ylr2j04Vp19oUuO8oKCdSG8XyuglLQMPy3MJ1CtRj64
ZCvSnVxkLt/si6Z3APqNNJkW9M8rkVrXPhxf3SQkN2wuOF9DIl+gO/wOiArd1Igr
lz+38NAxVScudvryaoT0BytYZCGSy5JYIqHQtfIP6SU53+KKDK47+zf9VBGEax8d
V2PP/Uythw/RdmAWu1z26DNAx5df3me0rCJggjKo9q8eaN+8E3xSUsWzv1RPXNe1
9OnML0WyKpIw+RvovlZ2aE6CtYAFy7JaDpsBhden/fcptbJtYKFe0DyEHv7FqfuX
DmElmMBCXRKA3dNctpnC6Tf0MplfYrpTpJXgeCriibVAEmlX00iJe5dHpVCXhf65
h6Da3h5OMY6edc1PeLg2efUcJEOkJY4Z1C7t+cSN3T8RdswhpRtjNkL6nHQ3IkCe
jD+nowighl7mx07YiYMC43QNXwzm92QLVkITLLiRi2CdEs2dEZqXliiYT4xl5d7Y
ZiujmlGmIt4Bd7WBhWLroGDZP6I71WRYsSITORunqdf3DIrEYxxi+fo9wYZecJnd
Z28tjeITfWvS2vVOgaw5c0DaZ7UJ7EBghLFKNTpTFiJkAD7TJG6ZFKAcDYYVLp5V
pIe7JX2Kw7cjrAYtRFtBqH7KPIh+YEYChNscQE1TpxnYdkKAav7tiIhhRVvay+P6
gTfTNWYjB4c7NOxqEv/uMFhQ7vmKEr4jx5eaqio9K2jKE/ZV6qWS3ej+rAApdeY2
A7YzBY8NAkWeOEwUzKVA8IZr4XYJC126or2otDR1CkIr4Px0LaTDA7a6Q5/+fEkL
DQDuQsvSCjRZCdlMBlbiHE3FfQO2HsPDcr9Gvem1Bs0CMRRBf5AhFhqdkvtMkI+p
H6gnG8OdIoVLizB6vzvxZImF3N57nt2guTlPzF+/hX6TEDPCqzjo31y4WHlHXkMD
xgq2etYRkzCqBmYr06YuaAlqjTG/a02Tapw1Q6Agiis6P3w7xZLZq+cqTrei3/hf
ZL2sAzEZ8S72Q58vwkpA0q4fhHSH+/r2BpLt33TH3NVNaT03U32YfjsPyfdD5M2x
Oknq4wnownfHW+PWDhO/4gbStX5ws0st4k1830OVIFohujTbFtoa0khfqwunPvO0
30DLAwRnfozYtKenguAN6ngcyhDfbXKCBgDjXw9mcZ2/EA9wgGsvefyFQbr43AD+
dNcHktl0hHOXO5ncIL+vBug16XElNMvIvPPwzkrHSVnboKae3Epj/ADWmC9KaL0Z
yQ2E2Tgas/BwSN8yzbizRJQgcdjDMVzmYpo2qb5JYiL7RilLrkTD8/iasU2PX/+3
03r3mtBvGBtZbm4XrT6AIFx1zDgMo2ivYamufModMW9fDJRsFBJtzR38nXSN8Lv3
VhGac2qJEHrqcbp5yzzlY0FwSZ/XTcvwc67aQI65HDrFZlNfkMhOTNwcgOJR4x2T
e0MMrmu+LlYaHCj/tZgIVXx4wmUXP/qZ2tj4upi9jxtNtZ6ysLGaw2OY0UkXiACd
sKezOMOMVA90KzCexVYcQ9x+8Peqm7b80XccvUAZXQrvp+P5rEMKWX0wXxZ9h8L2
8XFqOWny2tmqvmz9zHdblRJRows14sQpfrAdFQMaks49xv7DppCbvdCiAdzbFJc2
yzU251qwvJc6HV85T/rDFd2SQWbT6z/NPxzlHyfv2ANnTzZ5/bzNVM6c2o38AMV/
RPOIKjDgi9DWuV7XNLSWcaUFVjlO/wOvavEIxqjSD3U=
`protect END_PROTECTED
