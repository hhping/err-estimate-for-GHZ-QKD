`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
buW8WyMvcHj1GB6/P2OQ7ktgrIO2JUykIC9HfmSteytQADamKqR0ZC4PWBt21Sfl
6CQ5Or9wVETxz0ALd/NAypSLDiYXON/o2s+6PeOpSuUXbTxA/s8zT4qOJbdaBOJz
qY2GazEfqWMZMZzn+fxar5J9UOBrODvabVCUCj/pzFSDzjOJZB6icXFS18UWwvzs
wHp4p62zLjxJwy78J20EQubZXJTEEvtLhHLPN+yajjQrm0adQrPAxj66iRPS+ZXT
JAevJtnTY9keOWMgc/Qu8NlVgTvpMg7gVF6RurDJzmnfeUo4Cy8oSJ5XxtiXvIBo
6uSJTb/DjRScV3SsI8VhOSEm3gnWNrUVauHWXEygt3hPlx2CyvYyI4uZ9Vnjwtde
mXXQGA4Y8YXBVRBBvgEXbun6diMhC5hi3DaCgqgEenE=
`protect END_PROTECTED
