`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cN2hKt9TdhoPfbRuaF6mAlMQKSJaEYV222PEnad/hN1d8KxeK/NLtYD0WNtjGeFT
optu5bMTwpxj/+rgFBmSDVRTebr9e3dssvIKn1oaiZLgTHXQ0eZ2J2OCFBPlyCYF
g51kTzSl4dG51HQaPEPIYfHk6b9kxWM7dGXAYw4kkDhJxd7vp4JfillTOeOJFsSQ
JtMRujj8zAmXK6Gufjv9Vd+g50uvjOD+OmdWGhlbdPxGg9P0h2wAges+9XeI6qnM
6ZU7f2Ta+BMD8BrbfQ1OxM6dyFQArtDIoal+wMpfEfVWEWjcT1zpJtnjEo+PCjJJ
szIjr6lPoAmr1hFdD9TG9WCfaHGlVb2Ft3CxKop4nh/Jeoob8o86P0KiPsDc/eP3
ZuFrNoOXRrWrJoNIBMG7RWNthUZKRbkyw0NNTKSChZc4YKqxgHLAZ6zGdIPzyGKN
cPgILXX2ZiCdG9LpupMLX1F6B9QNoC2C8oXmDbNz/5TkqZDCvWfPbuyTJzOfCxL/
K8QAHuV/6uhf11nbGuRG+w+yrOdvzfRAI9c+arHGJuztMYHQIqf3RJdapiGqcg+G
6sDnQRXdXLfoIAYXYRs0tauqI/6CHheftnIcOUh7caynuI1bBHqhDpq0IayLjWVX
Vwxu4OU+JlA6SR5n3BVng6hPISOUlk+RrYoOpZ/WMAlWedwAYGqa4vjXOejH76mV
8DVj2KnBM3/YxbZdrGAOPbZOqKaOI8+xFPuyAy92zBi3dvkaSjY8T//wVFgjLrxr
tWbokkh7tleARlmANoPQfg/3PxLAqM6kSLz4XmOYdcKLQvgLOEem1PJTxmI+c0xu
M5tdxbykTMeN9EUf5BlB1JZywv2ULv8R4lb+qEWQoWJ1NU4LTEgiVS00DVtBIsQ0
vqWzX6mBY+u5ocgRa7YM6llsiWjRt40DCl6JEJOCMP9HW6UCavm6JxX0t7/g62RY
skGMbGd+21VRaIkhzV6b93Vmj37SHJcsMMrxlH+ItWOguqCa/Vri0vel6UC9btg3
UieZojjKv1EaLjzHirHTtA==
`protect END_PROTECTED
