`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rUSUlS15BoLtTWeYx1hx3fKci/vQzgir9qj76T17hwKpF9FPUslQ2C5rRCgNTW/
YKZk/GI62wfVpI3XuqUpPvxp3LGYbCF2vVnP/eKlXCoMuQ9KqR7ZMFHarrsMFPXN
gcSJ+0SRpWgGcpIeFYtAiZSBzUEpUXsvOriJ2nkqkBIQQAuK2aUhl9GAdR0Xfkkm
gSsENwmBCWqtJL+hfsfN9nP/A7sJyFZ1zAI4Fk6/uIB6u22B4jjPuzfv1E0ugK32
OzXp2a/Y46E2mBvFoi4o8c5V7u5eKuILQtlJ0Z2liU4oIeWfcJEEE/yS9zCSKhVQ
1RW3SJeZuem1JDO+MvBUE7ZJszZBQTeCGKzPxLzzWcJY2mxUPr/4gwKBwmMpj375
8jvt8BA7Fdz/6k3VuXWD3G0zrzHNT5Y3UvcXjgDnQZ/mEtBiXHKVZUV8SGbHMdr7
TmdjL82ihvKnvbjlK8mCU4SBjYtbehSrIS/DSEA0zSvoZQ03mw+Tr4gNy+D3cL7D
SJcH3IzPbqSzwyAGLYdT38vUMS332kJGf4JpZ4zwlFyHjfn6KqPuXHxlW8bn2VV8
rppNuG24H7cM7vr3HKYz3DpB6gQzm/dXniTzqMZbPx5h4KeyAD1XB3AIGwG12rgx
+fMmNQqz3FLFBTrq4U1kxvHjW3Wxq+wtWizRTNn06SLlEkOZQSnlCzQrTzPNl7cn
CoHGFXjAsq8w3eTYyCKnRVkxjRuTv32CHvm7pWOgBgjaVvzlCkVYjRAuRwk09Msy
gRkamTE3MYSMtP7PAKGPQNwXi2ak/posTrnYvra2tqqnPEH9K4TLUt+YIcWF4jbh
xDS1CcWRuA1HPrG0ULXgOZvC4NFUtAz5pjn2fKsHqMayHz0x3G8o4uY60uNBuq5K
2iAeGvPIP9GlXFslSOWE4EGPeJj3/LB1vpnEfuDMzBKwpftOhIWQ22FFAgaiPuO4
bubVT5Jocg78irHmrfcUTZFjqx6T6vWKLZLmRpZAMWHzPu3eeawMjx7k4u3Wzs/M
3JUPVRu2eXsW5OaaHdGJzmetBLNoMOguTBwtP8gGSfrDw2zFAhZB95QUeCmguLFk
tc7n38RV5+/ddYu6uJlEW8EuHdPPLakc1TJTvwF/dT7b2li0h3JBAO448c0REfVf
RSTaPWYpgiVwg1Ac33E7i3FYxx9NfYKh3gvNWT7uvPo2CLJ7VtDU0M+Q4Svhly9X
EnheiU8DgJKSyS97xDV0IaYaLYstCgKOiEAzlPdBpHrUfD87t1zYwQJyHSFSc6AV
94AbHkiYSwTdSlZ8Ao9AGurA5i9nzSTDaumQr4fdAZWCvao/lbHs1e+VckApvRqr
`protect END_PROTECTED
