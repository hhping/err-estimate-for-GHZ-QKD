`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGfInfodPrC3gn1hG1JRJGKXMl4r7pqXyMvIKEq0oQmgki7RtY63R4sV5BcCqgeo
6ztwPjyyp2dhepmqzTPFBs8QSCq7gW8YaU9PzolLld1gjgZUf/49qv4Jz9cMb4bJ
mlJxCxpl6TWvt50/TOENzPb04uT73Zba8Adee1y6LmGncYOwmTsJYNIQTGuEPJtI
9Ou0PwmTBKDYv9J1ZMPkDtvQp4v2FL1khYVs8ryMbk8x/GEn3OsCNbndkCSa/yBw
ZcbBmVdhAHw50IVGM29Ca+YFt86r//31u9iUMwcEdpyMiHIfORQ9N+HwNtlgsNdw
nuOMWw5AP/qO+1PVKPotEFesa4yqGQl9vZBkskCF8JuLLDuPvdItIWOVG2SDtE4s
fErzuVd7zHFPI4RZaudNbgEW2aFEV4yn6yzpQfMD1PcUCpEe9LBUMB9GaP9io6XC
gOnE2UFnbWPA54whT3/EledWFzAiMoRkdtp/vKEjTxSU5Pb6OyxS52Y38i2hixym
2Xa8kaSIwi//m4NwGlJezxKgX1z1YHWuclBZ0etJe51NFi/gSY/WuRqWJAkvss4f
nTRBqMVj34RWuqQ7Rs1Ag4q/Ga51qydw9X4Z8phuE2x2SFFFCyIveSRUG6CGVDI2
52EPQelVTHA0y+IXhcq3ioyd+wVOAZGXM3swOEsR7ZtMieZkpT69zJPfkoi3NjzS
8vzw9jRb7rH8Fmx3RybgP7+uKT6sI2SEc552RCxABFZ06bnCwfhfrnsiZKT/z3RF
Sfura8QxuPbjD314umLI7KiQYXEUeuw+JH9SXiJeF8I=
`protect END_PROTECTED
