`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gNMq6njV3MXsWNSgO2JYafbOd9eq75NIbQ3SnGv6nTEuM/xgrE0wvZzNqVqE5Ida
/3sgATbJrW43zbUZTryofvMRkQN+TUNvtazYqEp4OYEizwC0fRUG7bjdoqk14vA9
fDrW+mnQX1l3oOOKNvAnyS6Lo2DeuRmGVJP/7szL75CHEErrqvianuzZLJWLCqZn
4WbxKyghYT0RPSB4T94TCIWmjlUfi94KTtSIgYG3W4g1gWFb0AEz9OdZ21BxXobb
DinUJtQWOnzxJfbGA28zJm7eemv3bZbLgOqVxI7Yh2SKB9S2YoguoKd9md88UvZn
IgAgL9rF0iIuuvrfInJfQSDL5FApCH7jpVR9EZwhO2343HWou+RKdxTL/etnV8F6
q91Vqx1a+TOAruQGwUiqODih7NKNXxo+ditNADj81zQhuo/YCpOTIEqH8vqjyng3
OUS/LdPmyTzRh2myBltooHPqS0rocaYMq0DtbC8AzNABZipKhTaSuzH97Wa//Z7W
lX+INM/4zydfiALB3/HKjrjpW81ixD1RnAxliNS/HeUumBIjwljEJvNp3Uo9bzjl
d26QlgCDWCSN6hEFPVVFf9xFhBMhg1ZdhrK1KHdTjjsUH9v/HNAvVvMK+k0Z6rTK
wy3Iy1fWWB1x/z6NZ6sTpiZUjpv+ZSBaJMmitrvbHfKzp4lPYqfPKIVW2JVINGy9
EB/yqBKr2AmnTlZ6tHdVF6vIl145agSq5PT31P6IcAWRNir70PJgBPRHib569DcJ
xqNgtKjfzpM9MY1u7vWNzNzb88UQ9IDK6kGO3ucPHj8Bhx3c2ZxoSj1LPhNxMkxY
+3zFmw2+qAA4RtyVxSNdyBL0BHJKKk6dqZ2oVJk1ceoOrLOR6IG35/bId7M8dYgN
S+OTEj1oOe4WQi/3PvuElMLtwcwx00dupsoBIPFX/T9vUe6vOxP+XzlbD1+DPSgK
AroIByaYQEgEYidELLkXNgX4bIEDJ1M5rCAAc9rKsacetitGefabS3dmSQM+FXZa
r/75Y4oTqD66sjOXg/PJJ5HAcDG8W4B70qXKNxiyAmzCBPa6BBa4xQIBBRVd08Fs
cGLPkt+8hZe67sc7bz2k7p5EuwYq9ZlI6DlnJtpXd8Y4+VVXfREOWZ5zKIzWBFo1
VnQHRJ1r48gxiFGuuOsF27ChNrxR03UrfmeZ6K0Ehxj1mDeEzVe8acymeBypaNCx
0T7lpso8TAHKmCRNisk+fIPn2X10/R0GdXEpYVj7a6liWFuaWdMpcsCWw/qETs5r
M/DKdHk9vP5/UTUaWw202vcFMlCQtq+6HCoY7B1MDWKBPgfQAUnIfeTyXIn3W6RB
7LwtmhxQFzlQ178wMityhFC4CfI8De5rTzUlawUS9r9QKupdZpYjWviXm1GzMrh1
LYPqahR6nmHtgxdI9zwE1FW3hoV3tsegFzykmvLYjSbnZCt/SkZtRuIYrpeC9Zbc
ehltdpO476CEIFYdRuPRP3DLaGWD/V/Ajrn7JxIsm8A/oU4Etd38iWPipaYzwaZ9
Ll5SZu7UEXuxkzaLoNUncgeB6/qlTXnNcUkzEb71tqltVZnvcWbCm82/z+rJt6Dc
4ntcmSkH1fNC430sB7kogEX9HD+Q2E8ndRiFixTHmDqKZLEdkfHaHyej8s9/A38h
e7phe7BFM2+JqxLaH8c4BR2tZJojFK28X5sDH6gKiPcndjv48xMaE9PvaYwQ62zE
Pm4EfVfpCZRIeOJyEzV4Voc5cUis/FeJnChUem4R+adepyfpYg47yH5ihPMKNsWC
IlBfJqNR/ZMAYHgRVEqQGfVVcnUCkm3shbzlTJnH4K231igNGB42bIHsmzXnW471
jPQzFg2ltsAETOhAgr13LHGohD/RTjDkiCKo6/pIozOKlKrEb7tSCs1m44np0LJi
qXqWNgDdr+zUL4Pz5gJrLlbmhWWrLmpPzztMzcPCcK0jGhI7lTt5gAlzS6EKif3s
y5tCX5ObGqxCRP3eOgYygS/O6gHS/W6xlBYPNFShhA4DvVHLF7Zeu4BxTryrkgAJ
Itcecxxv8RHVfgtFwuhLfaj3R5ya1sZpAiPgjk5U/mOQrxB7O05AyUZRatSmENi1
G1QAcQ/3M2UFzGvA459RTjt9OZq9+Ske4P1b5sTj1Y3jAgs/ZGtY3wR+oI3JgBOH
IYjeTZfgHjg9S5/pK41CTmb7a0haVbCSZyhIXl2YIWZ64TBFGfilV3ks0HRd2Det
V1I23EnoeP3MvhCeyrWQhUTz1dT95F4wVdsz/aaR2+EBPBDCIT4sRduhjxyVqSRf
xt1+X9qK5MVJ2xNttJ7hAsC6t4lurylOSvokVKCo6Cjy3s5/4AsH2axWQyuE8Hh3
cemXSiqSECOJtTW+WmXR5dpFlsr3323Dm7xIEfwz/oLvagYSuFb7yvXLTGlSbILH
KAsnLgoyzthy/pDDFZpFMA==
`protect END_PROTECTED
