`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pILTllAqLQQc7VogzpX+SC7V876HLzCLK5C/KD3WxTEpPkcZVHk3pCGC0Ne0NRoM
JCmAFUFgevsAYTxZ6ZEC9sl10ddqzwuPN5wJ9VULGNaDmf/yU8t6YUDVG4NDVu2a
BQZ0vhyhZLB6oWdi2j2PWk/S6iDb2c/oa1UwCntxlFiqS7V7QnPZxIAK2XZGb1Xt
CO24pIbJaiUyJ2FsoSRCadILIYshyCeMBrMiDf0v9qasDDknpyqgl+VgX9lwDClK
IUKnYPltJPgP1eZA3f29F2ub1Ge4wYIPrBDsEH3dI223WSm/j5x3GkATMGwJvx1N
IKlrE5f9o6va6DynXfDkiVqCL04kDK6cj/HkOtdPRshrs6ozc/If2NVdAHuvjP/7
PXglscX+KtelRKKH1un0SoVZw1b6DPMjv/qB/kT5t1bHmpAvB25Kw+5M9Rsahj8t
WXNtUpe/CpeBmLP8GiuqhO6AMdJNIqSmX+brFjwsbhSQCibpsNbbcIJbkzj0PF61
`protect END_PROTECTED
