`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tecxGF6ipzoCe0GKsnXW7kQ/yvkRqABdyzTAIwsgn+530tEt12dlXUsCNLqqjwP0
33T5JaARHhi08Lbo0uXJI5WZIK4nNHQsOp+p0h2G5/QTACdprtMPJereIoHQH4Re
0qOTA3hOtUepJ9QNO+gx8Ri/DqYWnXOLWgZqsMJ5RFezP6PYvZE2QB6t/pXjlc1M
2asD8bJQtVr6eIla1KcnnDWflPLRYY37uV6Opc0YuWNSbSptZ/nKSdXq6GBeVqao
f+OeGrXyBDKZKr/DxXoGopeBKksRa7LPhrLndyZGxSemMXR63NVfWrpY+px49BPr
DDe7VQRt631LYWUgz0f2+M0rfq+GjHKo7Ezi+aRFR3RKFoDCepCXyn7AmIeaBFfd
P4Ad3BAgxqAsxqRl8ZPKPlBONyLQ0RwsFZIAgNur926nUtfgaaoDzn19aiEEyfle
gRb3kzevZcMGpVELFnY6AarhCfJVHkrZS9IzKwsWU6VnQro+7dmcO16+/GoNDVCa
3TFuDyUuaHpDpFYeqt0ZT0yKguNLiaTy9YFY2KVKguGX1bChdwcAXipdX+Tq3/IX
SzsG56vyEDTanMceGjUde4uDvkG+1kJc1CdkXFx3sgpHdzzZzbYYfIye3L5bJERT
fR9tp8GbZztOzsPapV47pWO2JVS6Bu57G6aI1kifBUI=
`protect END_PROTECTED
