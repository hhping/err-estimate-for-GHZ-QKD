`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ync58/mYBAQUIuoR29xuRZwi1dMctEQOTPwDHKoeO02pZ08RbeGGCxHhacHAZ3Et
bZe02mB0o6D+02QmS00VTvhWKUbUw0gJ1UzVXZP7kDj2+7wwz0olA88U6VEWXPWu
ixn/voiooYhHkVnjIFlJM/Lj3UDKmv3U251FkDFkoosjGNutrVsbFa5yB1kNEcsB
AkJR8NvNa7rMPfKPtAVjv+axXsZUEUsewjYJ8Uc+lFYKZSeBrEWmn8YylxL/dtzO
2m5raNG8hM1UySEalLSTsbAm8QbLV2GRCdSiv/LJY6kkZ39Q9OuGKghn51LjJ+gv
LmURFQeRbuOnaLG3lOC7n3LY9B5cBoRqDYv1UNsNNmiAB3gniykeUYeoIr3w3NoS
E19GptuDfTjI5BS8IsXFrS0xVRVAS77eGMkQWtFP2C3VrF3S/TZGELxTkWQWANBB
j6U+HDmCTxDFNXUuuFVPZG1SbtBJXplqgvHsquPALOZ8s496OAr2m4PpVWDfa/29
hoon6O61ae2ese2aHk9343UGzfZDSVrHHnvoh3lz8HulzpUizZYTmpY2kE2kFRZO
WBFaVg/eEqKg9szxDuKdlcTMHUh7X+tgpQhH12XisiHRjcTlpUrq8XDMCddEbjHT
B9MfHEMxD8Uks1gSAbrW68QVCalTz3kfQdXZvt9T0IciNtXJzMwmKLkY5qFHQ7Xe
kEKT1SkUc0fiOgdiCLPqp+CbK8LvtqI+f7Vx+/0cP34vvq90YwVCd2nKO/eb7Uoo
bHZl60wd4a40E38SiBAx/n1WrcO1SPS7xSs+nZasX0aKA8bHhn9KqRatoRL1fHnw
iPyFZoWp5wh6NgDT0+PKFIuqp1dC+fgMAJCzQ7cBdOZawnSaMUJi2eG22I6TAirj
ItfwPz5hHQSbO5qw2I1owIg/K+m6wgb7eUYrpzeXvjlGbKdsqmlPB4xMaSPXSaF3
X8Npm9Seya1MD4pGCU8FvhJg7taY8bFeZG/p2ROQqIqac+uCg+0htLbujo1SjLMs
qVC6y5kR4TViKzA+xBoUG08Hq5Gyr+F0F0ooQVZbWLl8nniWlwKmZAeFyeDjzyDC
WKh1tX4a5FyuO/HKorYQXZt/MSWLhYA6uJal6OPguxAUvv21zwyqMhJskZM0t9x2
/oqCxqa4yozSZGVGoAh8XTYHhoiL1QoESUAlLE+TSzL5857RI6oJjYI4qpq4+pNs
IBjrd5eOebJovF6Uh1TAjGsrRKYD5A1GmlWPKa36mMRNArNn1qeyA5UcunuMNo7z
B40zVbF3Fi4CEFPv2YimEmEJFXyeRm2dqrsyyx6L9COQedMfts6n1uDj/p3kcGnK
`protect END_PROTECTED
