`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Mb3clz3xmqIhadnQSxrErHyfwWNGjx95gS/xP4PL4pn7ClZaFFtcJ/Qlv2ZOz2U
tK+3JeSr00IFek9XyaiDSc2hf2xgS0/Jwrg+IElY0tsgwc6XnH6ssIWHfu3sySAj
HfJ4gjN0LEbGtVUeWe8rcKGImSyZHWncqW1eg7LndJz8oCNNOpEzeCRFjXlnxofM
tsKLVW0GBDGfMuAbGtIPwFpemfq5p8WzILM2VrAL3JzAOTLywAsF/Sr3hWpxByS7
jrxPznG1usmQNglotLgMXdsvnW31vawXKWNP4KeVV7N6Dtv+35c9gBrhAiQaIJxH
rKzR1u02P+Ao3m0vs7Ko7UM8vTGKG+pVUGAUUucTD5VXzKfpwJIjHHSgWB4FdVnJ
j8gCOGUwDQe4THr+zkQgyQxwm9FLZtEouVhpkHzOm6eYQ9RGVDp9azygAfFOxYQ6
u+y3KJb5y6R9pNJYz5WbXWi/vONNYCtkFr99nvboX1jA6ot/dQgyrAj6gF3YW0Z5
aq86cGVnHbz5p7QZ9ma9AbPbJgT8+ROls8OV1bTxCAbOnhCjFE3Gj26ZWBxE8r93
hebt0MJG4TXFCHUMVpcBcarGoNUQSlgxppOGalFLq+Xj0t54lBD742zHJCNStW9+
wHSZsY2dO89f7y/ufvUybevPiB4j2ts3qCPFZHXfiBgkyfScdNa4FFAh6vjjPDC+
iw9RQGN7GyeiqwG5xA3Y6At9n6sxx5ZPBIYNAOV7N1sitRSmzykV8tqqObGgIGtX
L0hu6FIG6dPH1ea2xnhfqhTbVlQviLgtZVZ4GNf+CrCYdfptxQ294vAEnzFgB8AP
L1JZX01sb7zJau613VabQXqk9zDTilAg9/6SMHuOhOPnRq9FDWmvna+Wt4r3Fkia
g8rwAnCBseXa12sbmrUxfvB1k44pjOdDfY6uZy5ThizEE02iC2sLzDyOJSJAj0O7
YhVMBqWeve9+YmB74G7wziNemC7bz+Vlpj9U+B5EJb2sRTTY0pm+74gHVun++hZJ
ZFX+3JDD/s+ueVGR/EdXThKDrOJsU7SC2XXUZ0LJtg6o4uSlzRh6si3hFUHgW1s1
4ClVKtgxQloYg54lfOvMGb3Ba8dx++eYxv2UtQCclwhS+UUhCf28WJ0GuDmyyF1g
cJoyZWaDal5yZ5roKavgWVWmQfCZbfxZhBJR7PBmMS808u/MA9dXLFO2VYzGZoPE
pTX8bRxRAJ8MeOfy2C6Ycn8ac9itgJgOqqKv9yMWo4Knmy9fXzqX7NVGMFVdUbh5
LblBivqDEBfvjWoAco5l3Sxo7jnUt+a0ZzaDZXNiZTJy6FfnRf/GY+Rm0A4Anuqj
ZViLW4E0h2FEyadCEEO7Owrw3yfRsgxOegTBS6gWqgRNWmZzSimLZ4tdqRo1uuyc
gqcnYsUsRAVZhY0gas5krQ==
`protect END_PROTECTED
