`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
piGLyL5EheFW4ft8adpRh5CI9Vu8s3wFASwFLchojQQBWinmuZud3XaEv4POOIHf
V5duyIqVrowUkoUIF4hzYPgGORGL1d3xAfbmSVlI8vAW4AuEmqd4/h5jH/tntq20
c4ckfE0mcajShhfQHUYAgfBsx4i0/TSc7oiiH//xnvECttYvsG3QVYL0IpQbCN70
x33fwDcWQ0lSNTjp5XsXY2llwqhjkqmp+fKs2S+VG/zYDloXW9givCeQ+/w1/myZ
5TQwpLx7F9ClmfZLlU0L/+qgpeqrcfDuRPUKrtcCfKWcAQDg7tKYFG0Y8YlTHyPb
+8Aqtc0fdNU8Z9PtX0Dhq84HTH8UpKHagkn2M8QdO8sCJ+AIkhXsoI4DDqokiOK7
GocgqOFXjj3/nIj1C0ETTLRJEJL13XjD7Efvp8b2qtJ7WBSMeTSnDBa6B7dBKoNF
XnQbCZMPS2WLkURzEKq8cTIgvKVEJx1UT2ehZOVqNefabrBuIclyucgL4C6jws9U
Ad0YbGY67Z7qkC+Q9os8Kej6uxnuoX6IDNHIs/iz0JfnlRBuE49T8v+otjn9QtIc
zFB4BWe9BNe05eYsEiTslISBXXIpUr+lU1t3FaDMLMgyEXsSODFSWuyp0rRBs22B
3nJby4XQruFvcGwtXBLde1LWHz7z50IBKmHg5IOmqy8pckFrOwp/DjL4REfehaqI
zDskKURoCrY3AhDog+cFjmAvir8w8FqhK9pWdkkz/MrmIuGTcBGkSeh15BGEkJ2L
tZHqeEC9JAYXJNx6hvGwwbEV+WHz0kH81xBQucbYUPdsPGhqCBmyHzgOPEVTlq11
l7JTQWbsSIagDf8Opsoh+/pcjb1CM+/4bgWoDf/XDU1U7KE+xWUKy3LUAqlRBRvY
a10VXdMZ77OBYAubUMDjEiMe3uKZb0ZbF1CbyVK6m/+0RofMOoPBqsX2NZWhjGGe
Ak7r1QP1/bus7SGkII03jEjSzQR2JemWTFl9Hi9BtQAhYcj0sHsi8r1hntVmMIDH
9DZr9WRf5KcaInh1owUS/br5pcCeHsoEXKPCyMdseIDu7Kwpo5othyw/D187AZWc
LFp3Szoi/gdP8JRghnZeuVFmMtcbeJYjUt/YE0nmVshbKtyO6wrt01CQbbUr+f+o
LgtDbN7sZ3mlFTtYuYiCiw1UhsCp6B7lp0RvAaOQsI35RQiTeufmzYt7k9COHLjO
Cf17lQhsCLB2zP9HF0sXcv0j1XUTs8SLGLiF5+hCHcLPKe0iWwnStfsYqw8ohOAW
4/dUzN6HWKlUvJ3tCnM+F/PpSSVr12841E+eat+iv0tEExjDpx5SWwysLu+rP5CM
zvb4zrq8Jvu27Aez8umuUqkUUPp36yT1ad8kGlXfrZ86vBOgBlcC38Hz6KVa7X1u
m0kxLhvdwVzeCms9jg8yRMXp0ofOW4S9SmV2DYAohXOyLvbMCxUXDEWoYNgvUzlz
KaVhjvpLR2o9ticCzWT813Cs6+XD54BSMneECOARWLgNQvToF1xNegtmdxZjNu8x
/Lwgh387xmV3F2aN+MldaaCnFARkgCfJXkAPtvsUu3RsBXc+FFsXdprST1TQfL37
LihL6O8QE7oLH2hLG7k8l925wDA/czw1hMOfBjejkXl0czRiuK6oiO0nQOMeHm1I
9BnIe//K9A3dl4wu26r7wOw+gAQ4gx7QjbMMulMG15XX2GDPPdq1+2+XAzPwH5xN
mSmbVpEEzpuLp2EwXyDLVezmk8xSZVx8byI5yDAOusIHvFM38PXlaozAllK0OGx+
pk48j85C4r4uOVPuB5gQ2WXU5ySsw2sV1O2xATP7pnqWD5qPJjMcRY6cEkoSUyTS
C7v14lpDi1BqVLc/7bp4JyJ020DDGposnNt/D1sISu7bGPtra8wjPl0TAm4muL3G
+30TFxjfjQzfuLdHVa0H5rdee+kXLzFjnqkHImf6VQ8ckQMHyg/WvHM/wZ54ND4v
zM3O4iOgz0ObiG9teKGBDV5DwNKecU75/6fmLtcNyuP3ZlbWxEjU6z+uI5Ri0a2S
SIdxE3ZJ6Q5swFvX2t89HDwBoi4E/x37AiWakgwEqpwVKgf2muGJGtz+sdRAA+6P
X3gtgh/FmsMicQjlwCUr/9mvpYXZKRaKJKK5+VzcTqqDxHryFAEFlhTHmCW9xjsZ
xIhxXjmu85ybiak9e16NUw1XixBH/Izerr0CFwG/eHAUZhB4fNYpnJyWCZCU289K
qKyrvwbkZNS7aLDglQCQE3rx3oZ4ei846q3E2q0y1QPJHpQZnlRyXm8ZgxoqzCvb
zpLDPQv0bt5P5Wz385Iuw01GZWmmKH7K1e9N0BmHQqXXShYro7T4OreTL7H67r6+
C+COGNazKe/6oTlqe0fy9FO/jWmgS4FsWMVTFZ1NKUNr9E618kUv4Rq5Xb5g3Ggi
r+CWOrWvkZKCk9dSE/K+bUU2WhhCUGbIkfKLbBCpVqxNAkcIxvUKm4Tat1axeZf7
QzlidiLk19bMBgR4CxZGdOp/yY8CqY2h90uzIvgOX8i4lNcvOczqANVdIwZYM5Wh
YSyK3V7JZGeH3CalJNZksD4cdOtpjbxv0pH25qm664Snig1nWFlhafxhvzQ49XBU
z7E2jwCBxLTJahl5dZd8NXO+A07AKRc9nAM5q89q4O0qn4YQKVEOrRoKDD6rRPYC
WdtNbeFg14N/pCtFCfUzlhIaF0hgDtUDcSWZgu/Bq9wnOkXo/HjJdxkcofnqOh7I
6xxvz2eYhyPHEBGf09OsMl7UHo0VcZXTB/lmGOuyxZReM1/V/miEMSOrhMdv6npt
W6Bb8wwDe58ld9YAQUnHh/EonF/ZUAT9GONNkANMBvIWnhC7zSar+TLC+6YTu241
Dq+iL2VFH6O+kP7MzASRPOqTWBnVB2J6kCYxjLyqJFewKvi9CWMoy/NLdBELPhhB
RJUD6g5B5VEpnI95c/jc0J3H8jfZ+dHUD/a2VqphPQUQLH/UvIqCG09gowbS8S/G
xFtg+Wia+m7qfTIBlzSj+gWuZerK4wNIIJUCi07IfBlSj/uqMIXEh3NnOG6a10B6
PNcKlRXgsJ1EHnXXtThFLIuiVvQxhRyWu2DIxTopxPstjYTLlVVFzrZqozrXfkbW
yP8bj6wSVxfnmVzRmJZQYuk3MEFyAez0LSYgAHqwSJmgHzs5iMXz83OJFcet8Hpn
6kJPxsZ7AIkwfC04vZj/YLW89BzsnifJTCanI8GJmMPHGHs6jmidN5xWB8LOY/2W
uX4wK27UpqIcNgN2PC9erpEoa9XD+TkcV0AaHk18QnKxM+bqLnst9OSBBEjRYDG8
snng9+oP+9nGSUs9toglfB5MFS5d+sDXgOZScVh2Ib2liBqeD5BBm6P+S15EqtcC
jqT3QpT7D3K78CwRrA9wH6OGV6IJsYFXYqIz4A9Zyy1iwT7gPuLFGVj3FtX5JrUE
TQuElcTWDEqMZ1JmElHhw/YXXWwNxr/MipUa3GcH8EnRv6slyMeH7sDj0nTRUYPA
kpHmsJqUqpQNsLeYU5nwTajhbV7fB5qez8nQAnf6nic/veanYD0rMP8/3hZ+iBz0
Pd3h0y4aHe358B37VLukMyC1HLLoPqs1S2t/WnjHKPeRQmgAxZqCu6RauIUVoRUt
wzkpSIQEUYy8b7hcnioDLOTyVcygDfHqe4SKRhAhbt0ebZZTydivAHjFwINRqE8Z
Lm5bB7p9w8nGHEX+WppptW+5ObJYeAa0zW52Pv57tJx23OAKeLjQWDnLowpIMWax
qzw6hLpPqUhRyAOo9YfNHE2xpVau3vAW1IyMoD4G5/A/CnLonCZE4pTeDWr3lZ/b
K99rVuWXbPhH8VhFFqeuV0boP492uoiL6lxn0jq8fTDPMZ9hAEsQS6MwK89cDllT
5nFauFOZtdT3EeY1fXDVxPhILLiaNJ5GUV2AsB0ueEOzDYfyP2sj6V59U8MwFF/P
qQzcF6CYz9t6lDyVQPdN4BAF4aaw3Aqer0dg/5jEQysOwEg6Vp5hged1XIBAaDCN
FETDN1JZmzJNNaFW4SKV/99cdbyBKi9RVC1bBDPVr/jA9w3cWNkHL3oaq/Y+mZq5
BlISS/i0VN71qg4/gIzhYmtFIBLV+cwdaHoaUKlNTXlONRV6SFeiw22mwYXulPbB
Pew/yXzC7ikQI/69ANZDVwNN1UvyT+EyAF6KCm00+WT/q9AzRrr99+u4FuHK2S17
QuCcutJpw/rv0jYJ4inqfq31O6+jbLq/oWm994TZEUuSdhDdihWxntiD2jCPdVlK
Q5vu50ZjS2c1aankozIYIGqqUroDWyNiDfttStbtsIMn89DdR1wC2KI86B00BAqx
ui1MWPwGlTeUtefDiq9HoTa6TGbTtIWSWZsvVNx6MjRNqX+T4KMqoqePb3HqKZ2e
gnuiSp7QSV8p+KO4EDnxnZOH43mLGoUei5kPo/1iSuhfK6Je3kvl1UzB0diUCwQP
eheSEaLQD89s9uAB0uDZPSXpIWkQP0hwX5x/rNXkusORWIVxhdR6MoX2es8ua5A/
gJfBU2ifev4qIId63KAoBRdqcPZQgud5w1DYYOHYpO1vdywcKK9C8SRqIcSswEwk
K7Zkp47mJc9ozX1MS0n6Mowhc+7PpsXHNmzaMBQyxTW4x9X0F8rxTq/hhb3+2aN+
vPFP7AzyxiGUofFGl1in4byMSKGxOREcFKBy0E1fvfr+ppke/mIDbpBK6jrw+6Ry
7oSUgidVPwJIl6arUno75AeUvMZpcA6tvOGDB5mGDst6DnC4XbRDnTB5Onli1sij
9h3FpSzTH08K+F+hfXdI9ugk/E1E27PK6gcV/TOFsdnOQLlN9PyDa/QXrKaWDg/3
aePzkQLuEO31QhxWgo0yxwFkdVuEr5uaoizN+xdm7Dv0yQ/6dNUv96o/B8ZO1yyU
JkmainVTuXx+PwRlou6vTfPJdPRczo9i5K2IJrwpmVxUynOFrwzfYB88Xnv/Sjey
94jO/n16ytyIbJN+UgKDi/pbeNora+MrYhI8Y1k6+NMaOx45szh6AZh5LqiLx8fv
6Wg5Nk2KvjBgi0tn6GtG7Ai69tiQx8IHf+c0lN2l5Ngp936ypGluCy+fW+VEOaAN
BSi9sQy9ZB9uPdTyzpy4llm3mF58wYQa0evdh/ouc/NqCnU6BxgfP72v0iZexVEp
eweOqpOVr/dlRXi4cjppV6432qoE6nH9R78TgPe4UBwj3/DEutd179tjVOAYeJO/
6Jns+Xe+YEOsMF+p2HW03coCojyEE0SGnypkZZDMNj/M/rYDdXTseRbsonB8gdJH
eq3DMstCFJOZ/HGYS17PO71FqchH0PaypxlMYM1AYvfm9DCsF9jqhcEPS2OXiLqi
hyVCaLDfsWxGtkOa7wRyVnbgqvVpSSLBcVyR1+VKMGbwUxo9ZOE61Sh61/p6Y9m6
WVnBzjL/n/LhWOAqJ9RnB3eXhD0jDgchKKijnFA4kI1r8rEqpl+pAKMqhyN6FyzT
xOg4r02VqQHi+vs3zClmWkLw4Xen7V0XVGq3Kgie6tjSpld6txLixZ33seTTmQ4Z
rLrQr+TKL8/Rr1M6cBV7Ui2HF1zrVFRFmfyE+5sunW7BgRkXuUF5ZRlTwYGWOoaW
boBUhEEVXVmzbcna4md23neCBw0ZQJkBf39VZO5gU1y962l09kh5FN6HovYKyCxK
znUQiQzG7XQ08bzDgFTUP6xQ6AR46xtZ05d9GhTRF0eOuNUrQtxTNqDFVrwNg0f2
ipbZrUks5YEyzPz5uyH+tvS2CZ39/Cou5+LgNqH6c6N95kFN4zsIdZg0gxYZMb+F
0GtBEuSNMV54QIc9VPSVkKOdqCD09tEkx46WEnN7g+6VvyZrp5oStuf46r5v94mH
Oq1NrUEHVW9/KAmh6+jlkdBMYd1TbjQNhQP8afZKTJVz3KpKchS9ZYLTU9zjEFPy
msZigUYtU4BZdDvTk2hV2aqMHpRISxBLLFz+SCN75yEudNNXYG+HlU23uDraTgSy
F2NIRb5MfzfyBjD7xioTr/JN7h/Ex4ivpGoFmORbW3OW40axPXHih3FHd57iuofN
Ah+fcTz08RWTYIJs7KEhX21XDuRAIXr9iWsynPvorA195auxRFyQ+AutaI8CGf5D
FtHPpWltC5kBpgCHJ7JqfQy2W7GjSM8s+fCiPXtWqeUISzI//E+7xvBP1ey+szLR
tPPrL3ECRNoTXdwEf+CoeVQAxZXvXsdvdAmp/Nlwkf/9IHt6Afperxu6aeROg0P3
byKj37Dmc/DsC0PgePuMhJ3LQIb0PeJx8/PcrejTiMG2PPhM7TQ1N2rnSaDK0Ew5
wwfn1epRY03BKUvcEONOlk759aTBwj95OvBxGE1pvpm/fJMeBZhDUCTIK+mzuH9C
hYbz/ZZbMm87X1eyezQ0s8MBtVwLrrKKStiIY2YOWINQND53N9Asw+yJmN0WpN22
GwFtSd4uznorymMkwlTjMR/K3rJNkF9LijkNXauI4hd3Sjcih5myP1+sQ8YLXUYZ
DBuZqxhiUTPXFs8Ue0lPhXg8DVD+WnedpYR1T10iE4UH1buAXonkQzZpyVdOwMTq
+IP97b5ZnMI9cOo9Bm2PJd6RGUt3ALBcZsBv1KB071TC8uooPQREWzuT9FFS+uxl
qe+Nk7qk6n0fWkGHu6L53D/Ik/QsevIesCO9qCVJlWKb67KPeDBXIjl+fjO69k9l
D604hhZzU01wf7D/c3rsUEbOxekqzmdyOUzX0W7HpnYlfWhRFqCBStCbt6LgrQ3N
cxwqw8SKCxSU6KqdjqtkRLWbSVYzP/NNwMEfbu2tCX/7kcO9T1jra8jvblMyzRqQ
wzisNj/eEWofJ0terxj4plzWtY1gB7GGMssrey6340nljsZAz+XkhkC46v+LrlTE
JBRZHs2BseQm+zR/4Z+tJO+wH3IlBi0+R+SyDQg3zuwuqwyVzEQTaTsyQuMoim/p
dZSzRBwSGPBOzHLxg6kn4v38GlSRugIN43W6WcCkDh66kiTKMEN5kqhRLRT8u5QW
7hb1bCzQdQl2XyGXJFMhKfRkxW/rEpnGvv9MYEwF0nzccLIAJfcCDSS84mc7HsKe
du+37QZGn/RWT+DEntO1J1oImQ3g9chJ9mxcIXrrbx6S8R/mn2lGwjUtNWGGtukE
IQeAoy0NT7SMIrZLnUDJygvWfxlxuTl6hUMZ4WirqIHeblEPug/RJ51rasEfL8uJ
YhxCoeYN6trQyu1p6SrYKPpuaHAyJsdCTIMsgXX3/6u2RFerbp1wLslrgw8H9y6N
JeGn0xhn5dhmysRks6G8TVXqZJJGgxoImoQeVZDxiUokH7/eshVOKuEr9Sjob7c4
w4qDGC3f/FgGPa7lvt0Q4L1BNTGa2V0G1B7xREoIsIg1a3bvhgGnn9XzfnBYsqVH
PHFKHbnEh30b8zitjplsnPamaqauoCm0y8jWA37cJL54UGCxuRLtT+Jry5fhbkLM
5/TiB+GLkILPAxMozF7DImn2lwX6h2xCEki178Goigu5eAyPK9moxtox+cmJAGgh
eP2tXb2SW4G4DGuoJISGq9j1Z8g7zEGAZmS54ND/n46Y/exvMy+OcgzQqHQ54nRT
0qxL4uBX1ZQtBJlHuEwSH1EY63Nbg6FzPo6B4FolNCUzJW+XNYb7eUr5KLzFzQG4
E6tihpYbNnjUjUtW1g64cZCv8EvK5736bHHt+lZ8NlaGplYxcQ6/2z+82/+uwjNM
37QdFojibF/AAYgtcDSPzfIpIooOmQ/4Mblzcx4/ZCRtJ0X/2llPgWydVnCuw/h1
lyy/BYzBMTKuJIr5efLwIyq62lFn5iMm0dfOWZP5ebMyriNw0hQcSTA/wwB28YQ9
NSqstrhmBjreY2GF4fa/CRpO5NiumALB1on7WbzOvYEcZF+nl7oAEzO3MU4+2Fnd
Bx5Va6jfWfWNu5inj3/ga8DtChGQ+XiHQVBUKxyoHU1URHmTLr7NTaUj6GvsNa1x
/BIGwMKpesLNv8jyIAusuSOlwlPFtKf25jBW1jAjxoYR7lEq1N0m0rfKtzhoLWgZ
UBOQDemdtEKtz2bpirmO5pJNasBCPUxWBVyaaXYbtFNBb4/uWSW+EqqGSyAJ+Hil
h+LkaDA0Maxlmh+VYnXBx1mgq+WwUt4qk8DLsxLbatyj0U7nzjtGtTBiQ6t38jyv
qOEH9jy3h7+UmTAxwaTsbUGurFbVcB+ypeyur+Xx6irA5oR4W0hpC4B51cLPqGnx
cW7kp3MQzRV7k6RWXd/4EOOs7I52swzKrFguedTkjWlpPy8QYa7KT36HmgyfMNYc
ejD0uucXNy/9F02vFQbafu7ofHy0+WTAIKoWBBEiZXGjg90ffLk3EBfb24WNpSVQ
hVutE+dq2h1Gqyqy7Cyb4WLUuf8l+54yhbtm5TbLKGFAGPAbaxqWXmxE8UGpD4hV
Vjv8I4+XH7b8dLZsd2KzIKtmVCS7JN//BO3XYFpb9FdANe4WmIAD3N28TrWKE1dz
TCBehLmYYxCvtRtZSopwjSdxTm+yq/AVa53YVGzSTE/vdFNor2NULb1UZ8JkGKox
kun24aNmMt137ZLfT3c1JJNuEv1Lagiq1EYu0EmgFuS0VqS9U64l1dkrpBQFsEdh
fpw2fDh1Qonh1CTAnCLvRtExKM4jzWT1eMxjM1pz6vgTFIQOrvLqp9EHc9T5gwJ/
nXGXAJbwRWR6WnUJCz+wyqJ46xgZ+RSxibNbL0dmdgG/0i+KBKpqZFG1ZrPNYQlX
8TNkwYRM73EePzdktZHDe4zCnBvUJNbXy0iQAGShp+rwVLM+/wbOLyPylZkrFgbN
U+du662PDkfF+0YJe+xle8G+RyYwA+XfiqvdORWfnrRrOKUl4+gWqBYVGc1peQrP
4Z2NfGKEB9c3AQUF4longubCIp9Ym0YosyxKNXtplHQhBoLfIuxAqc+Hh/GWzwQ/
C5m2BvkV+Yg2axkS99EVMy7t4oEKeX+yexl5ipFftZmStVkD73/pajnl+wU34ENG
pAbB4XsmONY/Sh2qhH0XludAUPooeJvuuddvCatudC3Vr4YJSkEjjeATIG5S+JnP
dWsCK7pQszkh7xWK7qlOWNIP/PR+r8IeIxuaydp1zzOAANpvl9TiV+mqwfJlz2Ir
PAiQ2VvpUIc0o0tZ8MP7/I7XMebWmzkPIHilze7ridqreCb/6SD8KUhm6L7mnJEB
p4DhoZAl3rhyIrjJAV4D/uaaFTSjabAEK5xiKh7+6C/mlFd61paf8PMFRa2/3MK3
tVMHrQfbOl+95JV7mDXUFZiGfpltacQozE26kC0B/34VylayGSTZCs4gTNjgQiop
awSM79mxK8OoaIC6as+zRKI5bRpYcFKa+e46jHOoXj2tAF9EYastYSGtt3O4O/um
v7EUpR0+FDKYs/msWZPD178HO7NL5yeprXfD7SfeIKfhDeUad9rGB16444YGgiis
rdQGBjFjxOAxWVBiH/Sta5Q/58H0CMcgMeUoKFfonjcdJK7h5MWcUBY1iuTobz9u
Ee0nvIJ3lb6XODvVHRbr9HYWJpgb07rn00D3RyxZwiZfSckbdYeqgn03ebs/47GY
ww53+WWdYI9zJWrVxL+X6p+T7O/Zvo9ho08nV1S6lquwpV5x7ZWM3D0IIxnINgpC
OUybWIiRFd3/rpQM6vd1IFUqAfPp9XySId0LD+IzZMCKKzm9vHz9nURHZBn2x7aU
4lBJHvFwEO6mc0PW1WCCEZVa34TtX4N9X8U4zVY1bG6/wF1ZH+YuxdeIUfE2cNJL
Zc9ZwoEFWvh2Y8cJnUd55iGMP/R4YbF18+Ctezax6KcXkIsuRzy2hHJdl1IB8m/f
ekZgM6Qcg4Lzzalrpp81QpnnZobOlb1o2gVgiciOM8tpM79UIDaz3eTJEehhhERb
Von6mGTthax0blZ6Ujjrh2u9q8TAro+I47dq/T4XlrhFcLlTJqH2QsLbtOJBCTuA
zIv0tBVx0Qdt+6un6p+aCwQxCJEu5PwL6Hu/0dlaA11PdbM2/fA62RHb0GbdKZlu
XurQ+HSAQOE3pKTWofDtPamGZ0/tZrB2fbJ6vMYxAlFcb6FxS9PskKcC9XJLSGsZ
uhRaMdthrJgz4JALy4XJyJYTdQiy7uzFgJYMf4s6DvejBBSEuSfMcMwBc42IbB3v
qRq7ARDy564oJfMHIIp399Qv1VHLtIoj+06UDppcLuMsd18nRwPHJZb0tAzC9O+n
pnnGA8M9axPaejKHqlyBUyUatpzkp3DmYqCHcu6cJAHPEvy+gtZe5amFEdUR9VqY
3JFXb2Q0uTY5y7bO7v6P0DDobvvHMJLcY5E41ZnAj3k9esuMYPb9kfIBvZwZ30ze
WQfQ5HqA4dOPH48uj1NaM1eJPRBtIm0gqHY+0NjKnPodTT08zueLxlQAeYSZos6s
Ld37TrfPqZ3NViUnKHmiA/kJeVvkm6qBRWNmO84d0b/VvXrbLE1JcUoadQpbjudB
CeULKreHvjqnW6k+ITzvUodKZDNLOOz6AsXA2R+w57HtgrFra5X0h/v3FPgrqx0U
516VY5kTMiViIL9jcyK9VQ6+DPVGg7IZrqKtn2f6RgOOeXHTcNf5CBwScYDzh5La
FIY9oSn8Esi+ADhHhpVmoK90qi6Zl1hqDSg4sV3Uh+FHwz5OvQ+Tx3jcx8mYMd3y
9P593/l+1Fzia+Gq7buWQhFecddy6wuem1UPKPNJxrcBXqq2+mi1vgHFUhJioOp+
u8g7dq8ODO9aQr98gCLqpa3xJ8RRpTxwNWFzHBytv14TFoeCmMgYNMhnnypEpMol
zvZN/kxMCXzhyC68nxCHQhiqwkuk0TisaiupyNQWLh0jJFECvThEEZpKCdkUF4Pv
+XrXjgosicev47cIfdkZomnIZOpHeBmoMN2gQSLe0zxaWNij+QrHEeNk+sGfl6GB
VPC7nvXa6vkYVQ/hztNhsEikdA1dC+3+V3wcUOXaxIN6XKzuwM6NhocVGXFJsbGS
HQFWPcLP4FYLHC7p1j6QUf/BmC1DmS/F7hA/m1laI5BK+Oceyo19p8qPXsHdG1BW
9pM5j5vKGpddAADTZGvqyVIBAtt5shKByPVBjMgZvKngWh7ZtD3pNFuJSgwuZp2E
ub2RLKkVsNtRUT9dFkI3+jvsnv6HSs4FdI7wHb5c/Xf/ojpYFPOTfkLyKWMRiti7
llJC0815nhA4db3Ez/k0sBj2RkUb+rYoXc9a+enPz2bx4V7FtGt2sasAGke08NQC
mXTMbgh6r3GDEorYje7eodV2lIM1+8M5xVyjCo0H5lYzWxHWAHoaQWzTy8AuGPYy
smU5g3m7rZue/6pkwRmti133qDZrZY8S2j+5YuvuxRwyhfmDy+qMReGFu37UKlcX
+jLlnvZrROr7lkq3NBuuS5rIzGltjTVhkr8t0NZ8EQSTzWhKVunOezzOmaHw7Y34
9oxQyx/PiGFVD6qmnU/FrXAelEY8cOp0JhefxNeI4m0VPwhARWVTBQaYUim7/mT4
qGTBDtdMDuUkIUrTg2LNS3VwZChpJArmtR+szJyIrZzw54bUEbvSqYuXQo0utI+z
ChCOwT5JyS2cvmAFmR36+pPLeRgJ3LoqrEnAJsPiI6633GhPIctG8gN4R500O+QO
XmE6nPX3rbTyup2fVQKnrbT/1xzLitWZkAVHktYAuSgvJirLxML9V6Y+Y5Hpp6No
QS4+/gOO5tlD0GutgZ50Ifh5ajeL0/kDowfQtC6pqGT9DAGcNhfhKzgFOTrh2ZYs
ocPigcwQqfytlRadbooevO8e4QU/WZXCXWrTg+91/5UQH6QP9u9afW+cU1mwQFLq
uXiy6npMJNDOD0u0i9UN2UpeJbcb0ZdGAkQuKpXXyELyPf2YDUb5oqe1bCwErkmy
Z1zngYclep2TmFPVMSBs6OX3QyJO/2LIklw0I0fWjX+hgmh9vRkwX1lLr024VweO
jiA0Y4F7s3C9XARw21K3Ct8gWaKPKe3ffQrNQGBGbxipNSPR7i1qoINCmQTdAkZ9
HSnXR7qBXIAHAp8/7kIb2VmI8LlLgLWrw1oO+QyXbZUsrpdJi6Z2THtqTP/tP34t
L+gOj4X7hGstRiFrziUOIrk0N/Mbr6xCgZimxVBdd29G4kNbAyb8WWEhlP3hxdPm
cySCi4dq1CLKI9TuImZQ0PuI/qEy+3S+bhuj8AGjS0S6pMoq2aHWJQ8vwPvYnkCB
9mmBX9duKbLr31Fia+xMNVYLVn6DvPyxcvCo60oe+MwEXZ25ZGJmj1WsDZK954fh
QdeRMaICZ/X97wuO5csosXGoNSHSILvXBV7gJZnDE1Najb2hvOyKDZmg4kwswrJo
OVebk5slI+1CRLs5tL8MyM6H4I0njZFucUx6yr4PYS03kcpsoTM1yt2HStAJrZTT
itO14i1TQ8loDHtVqokj12DXBTSoQoD/LFB0N3jZAJvYQ9/ZSzIxH5+IpA3ILSxT
gB/l3sYHkWT8Cecpgnl2JwDPwcT+5rkCVNIG8JZro6W2Sq0piWI7fRnTXdqjofJk
r+PPlhOF1XABrQpYcLVb3YSFx7OZqZFVvW7ej1gXAA2U/wBvda1N7t4A3F8axM4r
Wy+QYUjRerqUmDqtv99zc1daxPZuvTxRwG4B3yh6NKUB5ZXvp6EJXLrnbGTtFy74
RIwEMkqWl6dQvesSAKXnxMig+AJh90JkElUCxkALbOnaglVC7R5G+ZLW/+U0PDbG
IT56LYWfazLROmvVA9zkx12FdbDg/Nb2u2DEWVylQ9L5QhwxYGK3/lMUgWz3Kros
qjU7PDFf/HaVZW/nglt4WT4lK6+NrYozv/Jm6HpIJaK6tCg0YYP1+qktaNq5XIZR
jz1b1ukcR7e16e83Yaj0n6vxwBJwNB38rC2sxAiFcAXBRG67SSyRBc3b9Klfi1/4
IuoP0EMxciQi6k2/ZH0jhZuCcECteIjEdgUqXg7hDRFjl2dEXhwSktLJyhAQpYYF
2D73n/xGsxI/uBL/myxgkTd/duVxPRdFbVAYsvatFFT2npZM8dVI/NvCSEplY+u3
3nh90HBm49NIIhnrBoVYyHx3LZ97IFgxZQ9Xb4z/wox4o3N5M2ICAcaxf1F8mKPC
ODpYInueUn82DMZb5dtbG9cRI0b3DMwWsZEhGfS7fEgk7s4aFp/mY8gvZpbjZjap
kcFpgjkR8VS4+9LRHnLdBV0AAxoaFnyjrl82W7AAdxnZjQQwluU0o+AQRUclhD9t
U7bnQcTDd7WLKqDpEeIZMd5y1lDgylCEX7nVf1gQAZ/JhO837Sk9R35eCxh+PQV/
cwVl23X+J2IOVmLXKAnHfnzKgdu6O6Hwv5NX04ppHOwNTJuyNPWPTem6caHRerk8
2tvsSytJq5GOr+FOQCrCHEThJ3ANQWwsGUFc0Eyj8VlgIyxGFd6aOrnJlOmSQ0YW
ZqxkrrhRYNkrQMsffePMsLToA9MXyCZ7NnUYQO4QlU3olU1caQB9FDJkBPJrAhoe
eTPMKUmN6hsDU6EVlpr79/Hhyo5Br2X1t9TVE2XCHhHAdkCRyxFiK4Ts8R4YrYBw
PgnFKtUYj+iueXEa5MbqUrj4RcEtlVD0qiznYq3d3PYSI71/22YzYxeHS+xucjHY
z3ZfLT8wsyiItSaUXnflsdm9DCYhhlFEYGadqSSxDb8zfhz+9se6xNUPEgbl+nqu
rcJdogk9BMRzw30nCl1yKAeyiZ2StvjVGBRCSfk+BgJ5fT6x30Mudmp5towsTaGt
w1sPuqGZHx2ZtIXHQkew8x2Sa4lWQYjRG5AuOZSanXQ90+bOyDKG5L9wyCXEawts
M9YWCUw/zGKVQiSpAmYLYjGWCdW0jpg5VtsAbjxQ4j9jLDJsrUhfgEOdOo/v90uE
5hg/zZgLVDzwt2Zvs1M3lHB6jpNA45OERJ2wEphB3qDOH/dUJ2WDhLzNzqBieYK6
w1PqTTWzoAXtdKWSQ4TlpIpyq5SKkHGFYg1OjJC85UYEvre7Ms+ZNz3krTMnVCp8
HtBXEjZHIOdq7dH6pxLszIZEVlilhQNlNmzEtciJhjQYPeK+MQVh9Z5awdBIRAxM
K/lpBxcMxu1/Ehqp75j/WKoEjlVTd0pLpN8Fw63+Uj2zH2BTDQkrazE7qATJR5MI
cJGSJ/Mf9ekkeDpd9y5rRPlSAhy80do5nC+ZZvwY5BxdHLgqs/8mfliZiP28UMrB
e87LPccTCH+h96jIhRYKbwd39DJFZqOAbsepoOkO07quMk+dAtg90FB/yZiIemyW
8k9jKgedOPpgsfNnii3gventSr7YQ9rAZSZHXSeda0dZqnswySrDM503hLk2dQfQ
GFugadzmKT2LCAUyUaPHam59FsP/jdXUm9hrDJBNmFwSB0wPduDqxHd3jNNVoMSi
LArR2wIZ90g38kosiL4dmf8XHlf0CS6YrMXMV0G4hTloizsI6EVlO379agbUvPYI
wvwOim3CC/AIRQrmUj9Upe7gjiKXWPbdesj8UNPZ7QPOCapla/EdWOsnlv+kUm/6
keNURwV9zX78lfq96QeAJVpBPwM/two9Yj70hm5nk+Rq1ue2+QzZur5RLGfuaqFC
ZU8piGbI+A2BwGrZS9qpDf2NOmY89aUSpeRG4DfP9i2S/yi/Fri1lSmZp9cBgcxn
k6RxJt1bOqnWmJZJ/RGzSXhjDHobIQIkC11uj7twclIW/dQEojQjOn724UidH0/n
UhLl3e9Wljr8/MrGCmSETiqWeOttFwFkpjyEe8k3h31YTT9OT2EFtTwQh4EDMqMs
XfbH1cDI5KKfqifaCXxw4m+olrouoLZ7e4qE1sHD0BD6Z40CziSc+3npKy77yE3A
nAUrTttDj7F78Z1G7Aab3shVrvJEokjENAKyyRKjSQxu4acnLcl7aa8tnI3f1ei+
nlKcHJ7EfCD1QXOBxYF3NsaMN3kSkbs0qA1Ds1NEu/azJo+fHM7APro6ma5Bmbgt
Aji3ES1//5HL3JlkiAultWGcKq5//yT2TN+HNvYkO/EK+o9rYfWZd538sPukcmE6
akQw9uhncoCQ7wKiNHYmfzDpLMOnnmOi+2etvplgywZe3TRdn80KZrrQ+cwRXQTZ
+MO4sfrn68vELFGyz4lg38jx6YQwm+UIyV9e7bBo3h7fi6y21nWYwB3jcRmlphD9
8djBgogYQHWZSNXaW/MJsMNDP058HFSycTpXshTGf8UrBnQfYCBPWZ0AQqF7A7L3
UdLDwTb0S86DN4aOUtw1slEea6QcMZC4mW+j/qlb1YRgqqKwIFaj8UWbooSDcqjm
tDL0P/JnraovXukLfZxenCfZpgU5VDDJlE//V7Lc4hZI8q/009wo2hm4o0VtwjJt
g0XeN/WoiQy/RsVtvPuku0N/lBc79lKRHLuVFeyuyHn/lWoZYejb3piNl3JzEloG
B9Pjb//J1ajJDy0C80kKaYfD+KKaVG+Gbzn8EhuTGGFMHj0ygGAQeac7tGWGFRMB
514A1FWOWFAcmLadXl46jSxprUyWwxHMcz7xKe6cSkgca4zwhW+OeGPQEBVG6Lvl
XxbnUkSa3d2LNj2JpJzl2GOxBOYGkmY10ADY53hN7Q+gHiSrAdGPig4q27UiZsm6
B+LVWBRjWRjwTMENktyUQY+a8DxyH5eN+RHd05mhnPCbuRiA8wv3Ul5xDeCi4XRQ
STIANCkLWQ8CUt7hl8mah3dlv3iJCS5v7joshvVB3reJkNK5VkqMlTbjo1Ez8GWT
WTdtzqPWo39ifKPL6HAaFwH1C09vJXFihe+C7Qo7k78Myqa61w+kYp2kf+RmnnaH
iKFLuhui/5CMQ5neEY1cdQf0QRkWbjsWtqEi4nbsXBE+CRiHRKcYPjpVMax6/IKK
okYZhW9qtcbg+TgybSzh21hn1C1bkGHCTOClyMZbEv+d2BgKfVu7Be8J+vkVrywH
rL5IhnP3yRd9eEFQ4Vq57NpiCOurNkQSblUtIFvhgFzJm+E4ialAWBxBP/sPiQNE
8JbMWqXPupjNT55aB29VQiXtYT6+VjzYuCWrYN1DF9q4ehDIb7/SZEQyRupKh5aC
DeZvBf2JOKGv2ii8r96ydU7fTI+4+zMGIJXu06zVCQaqm64af1YskW9WOmhfivol
LOjO/vdfTMwr5Jsz+TicvJwhj0Nr5uTB0UACQp9BWxx9x88zwVQb3lBzi9wFyhHZ
LgR3S/Atj/3du2HsS1p5K69QlHEXUSfkRT8mxrslHIcAPywHYEZJtVDj3w2rEeR6
0G5KKmpty0r63zjHY5qZW9tblG8NWYuuUT0mJunepluNgVAzumrhZUJRYcQwtfWA
r3rpRPATLFjPC0g7/vstdgIznrblnV6UkOm2+k2WaxQHZIiaQTHrKiBbfPjlUqsY
2TbjrPafWWO95cDmD8fj14Sx64tb8NpAs4hmZMO3a8pfe1mgMg9Rcf6ZVOQgi2aX
9LmI2ga2XUg79jpFg/AXzU1Iz65JDZfl9G3T0ZQNlzCxmGoLPz0YnfhEXB10hiuP
OjKADVGbBCI5TOfl809kb9sPuAaBSd+nAQXa+e15kmyCyNQnuzSShamuuKRwnIhs
crCubIDnZJWts3KcO8RChuHFl2OekTiKh3tiz/EsHcAWqrwdrqO3ILlEHC4ZPcZ1
mZFCP+dCexfcwoEbEdwbmIV8gL0HgSZP9qhQYBp1YB0g8Mq+t5D9LkNMMO/bMGxf
iWT8F12sRswNJyjUtt22rUjafxVT1eGwcFooG6pLEGCyoL6XkzRaLYxrdtkGDyMg
LPxutkuD3VNJHcdEetDuMFo0N8l1WyZp0TkHFj4VvjHrIgVXI68Ib/KSuwVfkNUZ
JSU31L6n1N/8WGVb5M7I5zSQUZwCdHepFOlUe0l5LTFUpM9VEm8P4O8FS7I7+FRz
Se9uSOhlIu0s+KicE7R9qwB0h+BGAF7amSYDa6VHXXCjaK082sqtgJ7oFVQK3VrR
4APvRaLfMXtRX90ACkU0r3ZwEJ8usgZpxDb+BdvckFlWN79znMTGzR4WV9jXFIw1
qGuwDTC0pw7SEy6emel+qVr2x8ChQ9R2gm6Y33DO3MNxKrXjV17C8WXB3DPnXeZb
XcCdCBVSVI3E1e3Oxb5UTU68dusJPbHF2BtBkI79G8hgaz7+/EMeurgrviWGicta
DbSoKvO6Xj2Rv8hgJ4on+62+gkVr25CHE3jB5jUDO3qETmW3LQ9wZedHyeAVW/pu
xLTrAe74ZbpzcIuQiZN1Ct/tf2y77tMlv2uwgp6wcPiX2kJQltOjLikhmTFrN8Ok
fwbgp2oEeIZy3i78RU+FbyepgZ2WmgLcVABLJYuJvuKgdB1T+0LNGHHIhQ1xqVMS
BJjk+lhffBxpvz3miwsQiR+AUhRBOP6sksAhCYSY4wYoEju6wZL1er+V3n3Ep+Se
Loq2ybnscNlmUwIGyKbxKr0sqaqstIYYb9FzBA43XFhsIaIi9DUjHOULPS9ETJNO
F5BcMX8bvVeFRmawXBfkkdUG7iAXmDZU96UUb9NPH6G7MLuHxrZFCAbZplqYVE+e
aHi3cHOwUm7Z+aulwaRr8EataOe0JBgeRz7+PUwK4xiqkeZwAxx0xt6vI/tgokqn
fSyRycc/Pp2YDxEbstrOdx1MXMrrvIl0Cid5JnKQkgyDi1LZ0NHVJyZ9crg5ylEF
z/WC/j/7ydicwli0qRev88EAurTYHWjubgdjRoWu1hC4fAmeIdJkD8B9T+iDyNZg
NZ9ngrnX875qW2p9gO+9PTHC6QaFOd4iFaq7pu3DZtfGtiFYCl+f5BqH2T5nvZ0Z
luIdAyCTk7TsEPwpbxC/z/fuZFO8vKA/RM8b7TG7/ScH13PPL/dKTRWT7SLjpAu0
/fq8XbdL3+fFHq605d9KbvNdelttK2CEuxMIzPp3gOVPToJrLWmlgoS5lElMBz9O
9jyQRnsOdNmDrddUaY+y67Vw/ULg04Hfxotv0f0p9m0V3y0LT3qhXFv69VrUs1U3
GOPSc/T6hXpvNwStaCKvBdPAFk7HNH5SfKcwV76ae/e7z7a19Ty4b+mBjKrD5y2q
oDekUhqDGYSD0KB2VhC2YkOJktdUIM+LLcKxaAvGwAQ9+mPOcAKhRylBbRjQGauS
6GSZVvFbKXzpZOmiysWM97IhH1153CBnQTXqj7E6ESFbxT1ORJcJeZGsIyGNH0zy
jxhXCqqZx4RJuW6UsS+Vbx1tcLJt52CYRzIKAI5oTQH2Z6zw0tUkBekxCq6WYa/C
wpWEMRU58NJdCxcNW0CRdC0HvuGom22vMb1iTRZUiT4gsUcq5SlXbtYKb3+EX0YF
+GIEoLPbFhk6kdIEehJDOJep7JpMMDF4TBeyTxOmvE6XM4SaFvDoFyznG/zXRXLf
a0bu7wsyI7aLHJr9rF8MejqsFBqwDjMm2cxAynJ5dn1MZY7DYnc8SRhQf0vepbgF
oqL7+OoTmGpOR1u1iJoPlI00VWIcnaSJWPRN6mPztW7HwtpxNbB6JeGlBpjxgQuq
ywjt1qIz1e4u3HvnQI2px6vBAwsnEceNizqW75m3ctBpC3l04PrUHLPIzJkbLbRx
0Oeiao2tJm//lNgEueBXn736N1iHEhgpDvOps3YwwxeiKZbmsAj8ekcDYCLh0Kun
LQfuzgrcUXEwJT0Sg93T6ZrN8fG/G4L4SO+je70RwnkkLzpp2jvaD82yVekFLHiZ
jPeXwgTMBTm6zibw0qpx4wsdsQDXOjdNCPXC2BMvTJx+R+rbuwqQtjG35v9xR/Cx
/IC01BV2SxK30h1eTCvjTw2iC99Lx1IePEWz3X+xltfm7YFALzkHODicMo/q5Rj9
1WZhcEcsLiodRV6bz0GxGpxEbnW+xDqx/6oYABvo2HsV6gzO1Blgk4k89At8OHZi
Xi3cLK0A4Tce41KqJzRhASeOlovmLQAhT6jXptQv1zAv4DkIWVBPD2pxqGvPnz3h
6A25iMngnMdXcpqDZU64F4YPymQpGqU5kNn98JtYKFvDmVDdOkH83IoZUqeABz/n
GVUkLg1e3KfM2Oewa4ZmUwe7+g2eH7OmOKHffHmSYWf3Unr0P5/XeIM2J+/iTciF
zVAofE6XQatxvDUhJOdQZW88xn6HtljaJ3mOppLzdJyGNpkBBFCw1Yd7SiGeXjLE
2vXZsOfcOEBlFBShN9LH0DkbBCSAraA+ELdmoPd6VsIyiPaj3WeK9LYsdtKMyLPk
jdE9EF2GKZ3h2xXmiFSrfUVX6JvXlGOarrGFwZ9TrPpKgq2BOwhy1GAy6ZQS1qT8
bvvFECvT0T41TRvBFtESwTsLkQXceX942rH6Yigpg+h8fA0tUpn3v7RnqRp+YcB/
a0eDX0uh4yVeQwaH7/QcxsAI/Ssz66hVOwKVx018KYBpYzHkbpa1cNdwmBurwFsj
27DXmimcH8BhgTymz8P7ADX9PbHhDk00whW9P8iAbnIeY/SxWd4gyEeod3+YTeIb
MWzBCwZlHQKhq5vWB8I2rdDcDHX+SowMX/Ct4wd4T75sniKv7hCBhQQWJIt/tDYy
UZaAdaWxKtALrkR2P8GUsv7Ooi9OxmruYnn+xPWWVE1x0WppYZCTWrjJoDUWFZsZ
xTJo+JNLo4L4Y+OE4eJwBQGcV/0aJLu8HvDG3jzc/+NuirmaTWsUCz0pJKQ6UMd8
qOXqF0LIPFNMg0uYbnKAl+gSEN3P8cyEHNCEnb1G82i0fqIMhobUcVPclQDNQi7T
l9Iqqu/s2+8J5SQMqMUkDCf8v//BIO/VIXemuXO97Z5PN1b/ur5EMPIzC6BNjhef
ayPcNZFXFmIirESCaGagyyHGOXMCQZZS50I5KPKn3onJpzWYxlN5Xlp9WKS3FJwS
taAPZEpXI+eRh4RlOMR9Jl3w1475n8zhpltizXWpzJjD1Exvu+c7yySIPlopY7pv
kDV70vOE0d3oCdx7cwEKsY21asBht2DHtPN9UMdfrGanEwHIR4BlT6/ID+DrAfC+
fhtsPW9dn3ZYyVEugPUjruOGt4cQDYootD5XBkJ32FC/hRyslDSHhsADNnqXSETz
9HY3xML16w5nUMdPgih5LWsUibPE2U8FJi8J0ggh+X4yCLFQh+z2XuZ3NgQZMf0L
7dMqLxbvzlG1LNhGCMZlImvknGc9wxgJENDtskZvGMDz/Lb7KPAnjaosDvfT0Lk6
uvYgawzIJb0ySflCX2Y39sgrNHNCSK8MzqcmixJ0XIiYEILpDkJX6ECTg086dxfb
TF9zPZ5uSjj6HYoQLawFmS6fP2PA53xh552/hRKrI27ECvtfa1f/aGlsZwGZaMPd
5+FNrEl7YKbZhFybXn4YgQAOYqsYw3KDnKhXbrLYqLI21/r50dhG+vjujgXJBQuR
E/AAou1HjQYrMGjcswjRjDxxgKT39ASDNATF+spsPKixZP1J9btAvIzAu++4RlYK
5hygx5mTxMuG9QdSEQwOMa+xUzGmIo50QIKYUNaQwJfD2TxVrCaVrd5BwMz0aq6R
/a1NzMW+hYL5tt2afBMXsRJKhYbZsJmoiw99d9/SL8kTfImkDlq5VFHXZp78bACz
vG1OXWFP4km/ul7szKfTeOvsla3x+XtIDf2mWNMnQ+3KDmNCoqqMP4C7v0BYApZs
RzPKxk1nKALO8zVbmZU3eAM5uMr/a6YQdoVUdcD6XflquE700TovDfnCPgic5kVW
UBeigo+ZCoYNxzm/aivTyz2D4mLSC2khJTeTWFPRwW5uKdRJU+UhNrP6e3k0Mzyb
M/T2XfIPqfwmkN8Xf3fOIw8YqH9qFsl7YUjaWSvaTtODTKwNb3CJGVfK02KYX6NF
lrtPQlocZLRpJZyt4vy2vA/+JDKPwUz6npgzzqMTrTBOP4UYWePvexSbw3b+Bi+l
IhY+G0XTwwJ7PSy/HNeU3mnhFPgAwJiSQZJTvcF3X6fSZ8jIrI5StCYyrNL6LsAf
ad4rw/4qRMZl5rGwOvb1bzWAtUXW2v1+oeli1IDsmj7H6mEmTKPai7F/LdzqC6aV
kLHW/4d14XgocZ/ZED2ItDDDPOdW6LgrAQgz2AvHady4iq0Ae0MgH9r2LuJ090FU
JwYWV6kjMlN29idps35cLQ0/fLiE+29g2/rVwKBAuLrGRheytXRWZgsTZfQphxmE
O6S8LnxZ4uQpKl1L9LPa9wf4Da2nJDKkABg/0IrEmLrdpOR6IHp0ASccaIwSZ4TQ
nIXlRQwpbatozoN19Sul+ongm/tOGRJEl8XID86OcE0Z8n4w2Kjv8QtJfH4fVsMa
l811wYg4CMW0AD5eeVdR4kPzcZJUHmnjhrOJ3zLBUoEGNGihOjOyWCn63ONxpRp8
GF3DCSDyWvj1Uv6QajqfHy+bv4fQBcfX4npmVdiWnhHMpTVILsD3LLwFA5u9w9NW
yvyeg/9+7A5ju1Ca3Om3RbokPSgLZHyer0bTIw+ceWY+TAmyUsF3ANw651UCeKk0
WNqyXlRA1RbvQIDD9w1+e+LcuRaJUcNohbt2BRU4i7nlvJeDbiDmBrbVnCjgopK+
a4cO3MuvC3Xp6VmQrGpatlLzqHpoYliNl/8+bUKLmXfTMEmuWgz6p/Fl949Zf/XO
0J+45tmwUfAZbjSmTiN85Kj/uVj1qzJJktF2fyDGR56hVDehjHV8CHXEM9Kr5jVy
DQ7q8TcPSVu4IR2oFB2X/ElLhD0OX8hDsPZYuexQJA0gcilJ5AgMhCiJGwz6lG8o
LgaTXXdppHXI/G6pTmRbuYM5s3qhH31cx+BTePuT/xwVnF9sbun4Miw+nbDH/NrC
yu3GI7aj6emHldLOC9EEWQyxzONtEIu8903++z3MTETIzO3SiTCNeBqKZIicQA8O
kQ5VKbmeFBF5SSw+85tEC6Kzsx9zGVFnRThtvsYeZhBXFlPKl0bxPWSdMiF9rXo5
PhapLa6EKIvlbsJmTJhi/zvMLr83kaPfPlkvaRNTZw8O2PkuSi7fGX6xveiokXco
W515h9BwBKWvq69Vh5zUyYuOCvB2p1m5NI7leeSphesUuk3LdmEqyViIzzlBSZxD
HR4CKsehziMbeUaWztfdOu+jlHCZvxtWzmoZm4NcWYLJbQsivb0Ojs//M2aKlwGG
4kh8Nag2dOxjzO/9UQAro3CCzMdpTRnWLeZlluHC0aH1XoQVcmkUORKvr6zrdvB0
SVxsXVqs7LNNz3YuZed/FYwWZ8W5QNKwrX60fKuLfFdRi1mE+Lr91F8pvkdsxd5K
u/ybEZP/pksOXCdcq9w3TUMIuzQmn/iBudGvynBKcKYko6TpxUFsgH/AX6IyBlse
YhigGAKfTaQ7h8qGiJRjyvhF3EkHlJ9kzMRMKo68NES6oJC98lr4WM6LRqdpSq5z
2yY0mboUgGtDtgMuYwLv2CKl2wdz4wB5jKKdYNZ0o4KgoPnJn+TB2ksDSVNTpnc4
AmSZOppZhzlXTu4bX5Up2Frb4mSD8dl6HH+VoqyysgAHSNj/h94I6c0ZUU83X05d
oYpkl+F2b1m9V83gapMuCZkalC406UYcEMnZ/ZNd9wr7sSgpTMXEjYXLtDLLTwOg
myEeuuk8guEJsPPxK6mW29FqrTM5uq43cLKK687BiMqqxPZNh6u0xvRHnDcsqKYK
98hBklu7gBI9FAaMijPWKn1x2fkvSpDBv+gFkvJlrsG9RcdwFrz5Zn8fxOm4Etgf
QnfSEbsBwmiJ7csMOOQDeEO42CAQrpmXFIeb4J6pWtudefynWFP4HMWxjgic/0ff
6mnxp26iNFbvoO5C+VtnJqwwxqEyPrVAs97dnol6y9zpnc3b3qLuI5stclJU/Wwi
kyyERmXKJjjJL8uFMGQkFc003RUAe/AqRbZlNSomKsxB2XxjBpFgQESmljiquXNL
Cn590vVWD5e+wZtHBWus/C5KHTJHVnfL8zRi9U+V0x46myYuARD/CGL89mGyO5b6
DIbOpLi+P7iFSj8TPTfvoG6wRAev/RYRNl6c7hhvVlXQiXVzX2MCz3JmdFMEUNi4
qVRllndAMb1pcvWgBZkS9+y4LXCtZXffQGm0YlVqnA4J+gYfp2vG/C1szxCxkZYH
twCn4ICrSinY3YfBe3vnr8FcLHVn+NdqvcRgsg/n8tTZdvyOCiCNXzyec2b09KPa
uk3mL4BdvqHY+M3JoOR6KhKdPYAky+sEEJEwFrlE00WZ7noqhZ0gbry9frbwlbRE
ydz8uttUcIm62rvs4o9rjWckIi07yETQ3EN2brWmFOn2bUDmMZNEk4FComMgBxHS
BXqKQk/j++j2+P3X6OwWtlGcwKO3I6fI3+JGVCeJpkZVjToz1Y+FPvm80hSaqgeX
60IgzOh9kZ5RzFvIy8AA8Li2QnHu3guHcJV346ljGE9tqMSsJGnBpKjfeStro0al
9j8ha6TG3olp0U6DsTcw6eXIwcKvqs5rUPoimzlIaoQPvYov+PovpzorpuDZ5fQ+
3BGum3qbzZjAw5QC5PR8sIIHX4GXNO2zEM1UrqZzJCzplH7q4Irr/knGk8HPu6gi
XsnoRcIx7+PUWNxrpO7Ly+m/454/MYPGhioMT+/N5jH3gcTge/fJGvm3xwTELypZ
Ow3bUYK+MN29R+MAtLdLstZwGTsPWlRYDwJ9qXeCBMHc/r2QuH35TW/VtZ+R9mDr
VdAE86ywvUwJ7ADOt3NkJ/vBdfoM70rqZex6rWuh3cykgwUTJOm5xeIfW+JcMKye
wm1dZ3Wiuv5V6co3Zs9JucpoEmrQSFfAgAiMMQ9Nmm0vEKKVbyeD3+jGGDbkEhMZ
yTycscbCvLUMTUD6NvlFzR1TS+1DMjzcCovVhtMjT89Qs1MrKOLfmtG+gAzoSOmM
LxPmW8v4PVZrb74WrxSEspGU1TMwMf2RnZypbwS1QoOjemJXOfL8nT5ZMVaOXdo3
0OG3BQzWMfV0SGduYHfcwaDWGDe3Z0c+8JWKfyPmDUjWxt5TccqybF2wfLQFEAKP
pUkkPXIDnOR28cxY/iUUP7T9+HTfpAbYPWujQUGPVrYB/SGqtnqmW3aW9Lw2AZ/T
0bFbFjUJczVOKa7R8hRetF7tzb4nIrDBHpng7OM6HZ+F5bS0HTx573H/l1AximY+
7bXp9/nXZpokMzxwzjg92N8MUiUNFad2ztbUymI8tFgBR1Gim8/RC0LW0o6ytc2u
h4hs7HwoJyDZ11Af0FAVlzBKuHM40A8MRTHWnPqhTZUFVMKYiqAILuhabSjoBJbv
MWm/rnq87/g9TSjZmYWGBfGWX5SY6fPlzDj2N9mDaSYFFIB0kyxhpqc9iAiXEBUC
ar4RGudNZxlA9HiNZHr5kI6X9H0Cph41+6y3biWISzuavqUqwixke+FpoH5kFql8
X4xB6ybYGB/RtUePogrpRorS1jPlMtSeD5qFZyVGI6slzD9YWQ0djZYwTnru6iYl
cx9M5UvSfaV6kMnCRmdn0tMDwaiibmoi4gjJamuc8Skzk9qr23vEwjwOIuV9S6S4
ETbNxSy6Iucg6wNLqCO0UVPWv3tMAiWdrEfJA4mSiOloSXYPUnhIRrsIWug9isr0
M+hw4sIOeqHCvJPjcpHcNW0L58fBTqd5Lc/32cUZ5XEX1UDT2N1OvEuC44cbvOy5
a+83jW6igAb1ZFW95fnhLOydm5m7boTe3IAz21FWwJX0lNC3mLbAB66kaRQ88c5P
H4XK0fI5uDT+Mi8xtiupXKWCUJxk5kSPzfKVdPegx1nsiYcNHdlTInFs/SRMfHLe
49+nGP/6DANWMydFIpXT8TlYnHMb0AppybJCsnY8iox0ZUFGMyZ7XTQf2jNL5yNO
Bxop9gtcSrKV74s5cb20jbgNQ73veRD2oGbqKFkQYADm48I9W9CHcjv+ZJeo+6yI
O2RnOicfoB2lwHvLizvofGXa/K/H4Eopw3hOUR1YV8gKyuzMHjsutcVyZpIh6px4
nf8rHJykIjQznBzlhuZspiDlm/tfMQ/olKzoRbWkoFt4xiEB2u8egs/tP32f0whz
Kz62datrrJQkQkVrAj5sh2GlfNyp/NwJUmIWy31LHiNOzrXNfPUil4PWsJFQdT4C
PnPjOE4ev6XITUmXBwixPjAv1DkvqPkfiByJ7uUqlgDrcx374CcxZXG4PeVEaCJx
XupUIJrXWJjht01zcXscX701MQXwF7dR1lTKbhGXefOeN0OvXRmoHRHMBuMH2O+u
IOW8H0j7MMyMsX0xp1uluJovaLYoYdIimFiclNMNej67mIsVflsljpvvnLAq+QLT
MQeHGz4z7y7Vn6+r2NJwFUolHoq6xRx3pICHe1VsvkKmKVsMJZdQb86IwFi7Qsx6
dMhzJ84LrG8tG4dfaVO0hGrNwE4DxnO52OFi/1gKYx+mXCKPa5NyS9L4ex765QcK
OVtuyznWgiOZvfsMyzwTi5hdckj+CD1Fp+zBRSPHZbuf470V5H0TAGu6t7m6SaP8
RGIjJoLCs5v2aXzlqBHUpMmKd1nUiPEOfdNqx+cAfh5bbZakfC4oIrVjvCFDuFrs
5ENlcNaMKpADbeFg9Zxa4FKatAaGNTccm45mxzkrdKs2GibacANTSkS4ZW1jnBdE
/6VR05w6MTc9l4caia2Io/aDbUfFEwpPqLTlAimLPTYT9GjPEx1MOIoN1ZN91drd
yuUwdK+w2zhwHBD3kBw3KdeSyQlm5sLepUK3W3VvFZHdkOyxFv44kZ0SOnnB9BdC
Tvykx+RHhx/4r6NJ8rLBGMkbQ0Gop3YjfAqMWGb6hG0rs55F3uUCY7oQEuiBVeo7
LQdKXEdU9TaoILPoqzCxfSabcDNK3nIKZGIuMpN1zHhH7DEncUQM1NW1oL+DVv4v
AyM4zr5I3lhkitsZlbjP+F6hKczzu7P4I8/nvaVJegRpF6IHRVj00v3H9prE8ISh
1omC3jEwLo5dQVQd/o57TQd+zX/oKLbU2CjeJv1CC3XiRXsdmnZhzQbfkZvh2T9Z
o3RLQEPRbGZD6KGbAXLdSeu8mcJxTJBya3s8WeWLvoKA/tn0kErx/xupA8G878Yb
SYf8wFsDuTI9BvJq8dZ4+58neKtehOwOIGYqFG7C2kYpKgBMaUrA4t6K/Ix57RDO
61VxIDpDMWii10QA6jp/A2IKo9xbL2k/u2/rJscgmJqusuJVNvJUz9n16M6xIwdT
26/1pq9Vft1GZ6jzw4KCn+G8woRK753FnJvn6GZqNePRJSkmPbzkJn3rzQ7pqDKE
GIiAufttg5NagusO0SDtdDcE67lyNgK7S+GhPCqaC6PAvUUXImRkroIOgT/FpOfY
maKR5mmjnxMT4kqVcL4PEaXA+NtMSF6Z264WoH7dFCg1Deaemv/dGLmm4NZxZNQk
CeDfLuqgqBl1pJ4x2him7vH+cFmwI2mxcEQEkN20S84/OL3+C26wIRhFS6I9/tJu
eNhslCbXSquZiCPYH7cZcgLe5RPb7jl61Ms1WfW2Jp5naKkJ+0j27j/wjwVaG4hJ
n39lVmAjmJ6eCYWl1yeb89kb2e4cQUA4bR/v/+JKQyX6oEHqDU2nSjgGLBcHKIBY
pRDaP20mFnSDKmnUlYBMH2lQAmfwInGKtnTzhknqmcUnhvpKmk0U6sBH624fy0vY
g58XEj5DwM4fyq7Dc3QywhkunDakwxU+puZvOyW9tJ3igPwIz39Gj3f2h397i4gJ
uWztMlDwob7D7W8cCGpG+LMq82XVxo4HDWNfOi45aZyfhH/EleECNeEsMosHYBi4
MOj+epcNex050617vXCany3OSy4DshcYWhzQMjX3/kTYTWVIIgPTlCbJvYQCkVdI
QbGEisLIKeCS94U2xIFdQcpcylhAQCrAxSd8QB1W3+vWE3LLNbyTrqbm09hMlgRV
v3LyCBiJdVqUdPUtv/j5OjMCq+/e2Ks2xhl0DyrgNylUow9+4lCgANDNIJqZ+u16
+MJDU7GNhOV3bAFpFcVzmMkCp1V0XtGhKcEfpX4ubfBeIHRj7yVm/2BGFzfdHHpb
ZIPpYxD1JgUOkKtRbYuOhhM2ISldwBfyvHu2zhTGFiAn0XkVFbUvSrklva3xZCqQ
4FfnJYJLCvynPrmyX9kYKaz5jdYlHCFsDKfhivEBCrjUsrzEpclUpn/bCERrQ0/J
g1oLg9rh2PMywCBO+Xo3GSZajGzHC0bEtSuuQVMSAu1lyIzhFRCK3q9TN7par2jU
E8T2htUcby9IIw29bTM4iXsqt8BpuUNSf8YTq3Th/AkFyNspBqCD/7kMbbzlq1QH
JF65LFDKVFxoKGHbPmGvBXhRSwTpIDnJujF2xANODhLizXzqHz9+OEKfrpM4h2rZ
DiQzqXTFbrBIV0bnF9Yp+BEYNVU6NokddfWxlSEJN0PGzpyxOlrcbqwMqTNwkB25
R5IQ4pFoQ1flGUAQ8Bmn/m8jBrN37r3h5r2CdFdEhca6q+r8NWQknBBa7eedqM5c
c+zwjxMihERUZinSjk3RcB/WOGhXZicOGALsQvuU2SCPaCO4Ix9RbMuikXaND6P8
GQl/Z4T+VLm2AWLnbAETMR7m7XrIP5AdTd9xmNZeT9amEI5649qb+9qfKpcvmd5M
BJGmHbotd/Mfy55Ml3Xt5U/QkBRq7Qbjz65jLqXA69Cju4nf8vF1kZWBO/ExLUGP
W1QR/jTyZ92zCF+4sfVG2ERGrHfnrEGjqEoIaFf12lab39iTqcJnDCiAMQwxmAeY
bWMfGThdh4jNGHm0HF8kqZE+YA6wNyjgA3jCzCVMnzydFc4BwIytoy18MYYEm+3a
5m24bDa+e7nDP+LqBb2IHcRYHVL0s0goNbGs/qfuuwq8wh0laxhjBYvf5owXtV8N
yCjGr+zgD1kbRWOprkLtqMu7lcytlvVy/cVkhrN3sQN6Vkf26xB78EbQiT0lfu1b
xzV/zRjusiRH4b0sNiYeEJyVlh61iuvtE73SuVNFMMhd79eTf0RphTPiWuwTr2fe
PQGBuWfEgTaDFNpXb1VZuPs7Ley78cd1olV7lKrzr63WG+tdMWoF8sPEZGyPd+p+
G4AlAm9YaFL/4kzAIjQRDyfn0eZYL1GJVKeJ+eQDgh++s7gwZzFFZYdyh4ACDP4h
M5WahnwlCzyvwwUrn4rwSs+j0H18g9Eoi5iqv5Q31yDJS9Sg047CRE+tSxm9Kat+
kOMx91APlR3/D91Fqhd+zQLoJfw2mxt50dsq3QGRHiQrsZhbzV/BIbb/mk5Zop3V
ODBiiPZSgWYwl5CTk8gO5pGCv6rkwtAEXDl6COdqW4zF0YFQKE9SNHt0N7D7a5g8
GENC3puCUYXSI3upZShVOA==
`protect END_PROTECTED
