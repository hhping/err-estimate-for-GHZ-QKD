`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4SmZ488PtiPEn9gE6AugiycfzC5K6/zsPIIVWlh//SbQ4XEF2GN1FOPFT3xX4VT
9UOsCMB4KRU9b905UfECeQ1fXwRL8Pj1qMuynrtJTWWKyT/HvDGA0f1qvMmYkLnU
PRZKOfJGsA8wsSMPdcSPCUxbYi5njydu3Ryw7DKHzYYW0MAhGhPq6CsXNgbaGcSQ
rqAarhrlvTiBJ1eKnCMf142G47Qw+h6PNlWc+yhzoimy3EoL+i0bgqZiE3OZ9kXi
YqNmknNrFL2Wy3uc5UE7pXzz0/pAol67zsSGU5SkEXpEfwU1qywlLwaQaLrW7Rw0
8g6xK987dE+/1FsJNs2G455jITxa41mPnQxink+899Q2ZGs7MVlJb1daBXjvzw/9
Q3C7REeKC6S3deEqhXEJ/u1xlg+eB2qARYBkqu/Pj2X9dt142MkIdSqRlntyn+y+
mcur84L3WnCbsrnmnB6iRqOypl0uxKE8c9EA9CgfE2CTYyaW8CqMnp8AeKxNrzGR
hM1mJFsT3YBP2MtHOYThcNV79LxEodPBgtzRihWO7izEm6e20ojey8l14+yFgG9N
mbTTUaAimEile4g5rCmEiBksPllnurZtVxNqOKEleciJF7U9Y/iwNx/1YZ9RB/qY
4dRjkRfNSLYsQD5zYr1ftZKcY+r4t8JeWlmlBWGqFFAwQhP7Dk2Ez1ByvyZ1v20i
YSY7lFraLphzp5usmfd61cdMzh447Vt2JVB6zkwEzBxSGeF8aeTBiZYg5BsRd12J
Aj6nhlpSeHvFrj5Fg+H3GcwL6czRwUe/0inseWtdhNPPxuO6LfvPIFFlMetxdU44
uTL0yds5QBFfOCssTWIIRLpqsZnbg8MgBlanv2x8Za92RXJkOR4mVoXZMxUQIsPT
nFS/DnrpTEkxbbKhU+edIiy5jKz6a43gsuUbE30sQM4pVvj/uUQR/mt0vc/Cf7Q7
`protect END_PROTECTED
