`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6AlxHVyyHI1NGTMMxr9v1CQaPD5rWwz0gFAa2rroQhWee06ldpv8qqjfpo5FA4v
YzEL6EEL46LmO6sYVADMphTPAyZcyF4pyWLFLk+FwrYWOzVhrLuAA0UYljJ6uOYH
LITiBV2hOz/jbMYisFxmZKqiCv3vJlYYv36Sl96OXYHHjpBc+DdDaGQ/sd62F+2F
uUnxRATyICH87z1j+Z0OeGQnj4aGTEfFkXXBwgj2zvwh58BjtP3wWpJIGC8P8krK
FCn90UPrpeqpphuOOR1kiFoKzsPJoj/dNZf+zeSo1PQ77m+J6+CGQR6OxtyUfpsb
vbCJelTdj7b5r3KgMIGLOnTkUKLMI9zdB67XGsWNZlaLrSErxL4GwSbR7NFflxu9
RkeuXBpC1SqoXpqiqv4qEVikQGDm1FUyCNUy+OEnJ3d9uxBWdQTdxMc7/1FVrs+D
eKHQu/NKpcm3rLXXLNY0DT5+0JDBDNYMg5z18YQ6+5kGYgOcrxQTMVAQDZlhNSGV
gQZb148REu0SgcFPT6wHPnFBd4pPIl4ol1dXTinVvVI23m1k+5CFJocfwdMA/YP0
n19Z6fzxWTXfH9BYDtrflVjNA8hJA4EwHHCsdIynL1Efxl2Raow0XGHqxgAAHJLD
EFLBQN/yEDG8zsIZoSyfib/RkXF5Y0nxSxAXT5FZrvvz289GNnbThN7jdxFdOGIa
STMrajo+faINsTaVbuDeXRIkEdzxRsQL0cx5brSTJgj9z9tt85MlHgBZUeCe9+I2
sf4HSlPkLeWEefycRpVmT33ZDa7rgdc9PJ51qgqiOP7E8ou/C5RZW7sWnW32oUYA
6Gqk4it82r3lR0n3ibQXLYbDyjZWAuwph8oGiJwzZ0v67XvVsAs2aXawpfhDmh2F
P7B4jjZM91qjhJYz/EtAOOUN4rvlXinM/YXAAEpXLolwXKbO4boWg92Iun4wzUWG
GWKrSFiiwtzSrHM3p2ph79IcCZkLKY49w9fcqcWzj/IubI5Ku/PvP/Jz57xJ/tIg
UFwTokpxuosJCSn9KGlPm0LI66EonjWNF2LzUyBAMKlujy4qlrdo7dDo+vZSAYsc
o/qUvZLIrxnUyux0r2SEHrE6krphNdNqzQZLhY7Cok7uianyOtWgHkVyaw87xcyz
Ump+T9D/X9/uw3KKV3npYQtsgC0ih1nWRnelZsspLyP8f4sfrFlU6HCWmf1a165j
5TIbl/bRX7U6cXUMGMnmSaGmy+oxL8/DxN/YqAkmLqg2md45HqVGlHRvROU9bO/9
UBiSeJRnyhFsGa2isdiQc/o9rczWtfoLhkUulkFN61lRSBpjfMBq0Dp5Dgj5xSTI
nttkBgJ4WIpdMgvXlZtbB8z4ogvYaqd7uoBiErZ5Lj5jSp/JhaveRnJ6PkpWyz8E
JRttdhcdd4/zR0jixzZ2pNYVSsunX+8v4T9MsZVHahAu8s4bhUqikZusK9Sjid53
3g91p64meRusbGP2dUEHskBFVB/eWTgEQi3ChWw9F5L+P85Y3UYyZaW92O7/Fm5t
ruBAgZBA2W+1tzenojp4DxyeGUbdCy8Cn0UTUIKBu7w=
`protect END_PROTECTED
