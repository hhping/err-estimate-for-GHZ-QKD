`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yEg9+v/OAQZYWeKH2+qbC0YMkGj/YciSHct8CUjHNRwlEH4FWkyXKF4rhy9eJrkQ
i9/GuSGDAN9uUxdRo3v80K32HECnS3W2eSVFi93I10cEzpDf8Ms0bqX/h7GDqpaw
+Vo9acRAtze8l5ujiBpiCO3gFnxN3cO9OtLAlu3yTHwRpScRrT5XO5HGCLs9zGXe
89HgaNJBuVmu9TfwElVUX/ZQ8fWrQmdYv4PwwtbJ73csdD2zgIHV4SSL1AFsKZgC
atnxOy1+N6cdXFVkaL/EEpW7REg0bgu6GNPY1Bggcd7TZ0jYQkmQuLKAspE6wSVN
V+Y6U1O+IlQ81Cjpoi1JmJMKOz7wJvph11I6B+gOfmQ97Gqp32RujTuAdlmb/2Jv
QhK+4NCZ7qPodxQwBpC3hxf/k/tlLEFmbiInQ02sMdlp+7QFDcHJGOi7j3ZN2ohM
qiId0HP2h4fqcJGojTCuGyHgdaWFQYLPUtmLjKjy3xLVKXEKGi9BTPHCBOxIE4O7
YZPJaW1UZdLy/Wms/+/gondK13UrcZcCBVlAm2przmSgX7NCCW0iWU9Zsxv7YXvT
/6XN/0AEIPNSBeK4jnlfVJDKpihUNYqx0CQfY547d6ea9g50KwzGvJpLiDa2BgsK
0ZdfH6W/xEf3yEMFJx68RIR+M8bEtOc4iCl/Dzqsro4mqssSUiJJloZS6mhMYOeF
xTFT6saB3R5QVkq4zSgvvE7qU8e4TGkgzWOvvEMuM+H8478JewUukfnJ7JVMkU/R
1so+ZZnWsQvzd6lmr4ZggOoPj0VoSkvP/Si8r/xxKTQXNIYIGJQKhX5uTjZafm/P
d6l6HoGTqiBKV5L0+gRTXpryRklcMh2mqflP3GyxdDKKDT2FogBhsLQsv2ashqU3
vDBvwrn6kQ3pp9aKFRELQTeQwXAnu0miRVE5kQ4U707+l3K/4JOIP7QzrGf11fRt
LTu4zsEp18hA4kEmzm6M7YWpSP3g5fbRaD5DnXfwjwTyc27eKULJuOYEyQwN9e1e
i/J/dkNoQRZtd1/m1b780vmzRMgk4Bb1UBdyI3//yOFNunGdgkKtPaYT8B8IKDQz
HdDHznmGcoxiGx2va9F0c46y+/ZBQccraXmbvTWJjAv0cYmABiHSZ/0lJFbGyXkl
39/QVSlxIIadwiKB5fS0C/cH5l/T6cpIjaUcpqB+2ExDrq8kuMVJeRHnwsyTiNeq
2hr4+HxIeSLQ7gtInQcL9XjJcO9WzhhMg7ZimZGwDr3qXibeqchmbxQvq5aQjVrh
SEniTuW4mLiesjfpDzK58+CwAkJAHsUI32y2t+WbvoinsjYTzrTgFllwoGtaJTyv
SrtSQEbnFQQcvMIjQJ3jXnEbpzFnIbahszl/NyEdz5LQkfmQaJlEvk9N+Zjbe+3Q
UmCjROMMSYwxWOPy2OefleTcV6i/F8U5BYddb2l9MLjeb9gNfi3rJbOI3rUDM2G1
wPoUVbuZ2IRaCh865MGIcHNecE+cIKq/uXVqn71JNm4H/tg7S0gWNQ5p2n7rCT2h
whNyQZvolScprJSHzxVx/vmH/sPsODC38GjWGvfO0JrjRQdKIhASs2uSB9Jsdy/Z
dlU0NL5f/KM27Tw8uW4jCMAg+3ptuPslo7bpIccuKNe+8Poj2Fu2lFooDeHRH9KI
zaprBP/09eFIQpzae8JxJfImdrFR8+hNalBxzNBTylEC3ihdbOCaybaDGdFnDLDA
FcM+tq3KNN0936zfeMWvESx55jo+LHzzEQasi5k10TQrggSVkkrtuNTnVx9SQ0tu
q5Y8TrdyMvYZtlUOAxyqu77JCfzhbhFiJdjx8zIMJlxQCcBjIjaopsmEs1kh6Xjk
hgdrO1+PMMO8eKokLBpV+OgKMRN2xn84AFkqZ4v0Qod0JBA7LvR5mJrN5Zjgqa0u
4lQCkfRtiUhi/7sDov30UShbfdSGmp6sBxXVTRo1Z/KzaW4rmEmwz9WCje5eAI62
o9tuwmT97TVyuOwCEppCx7+ZfJGBSJq+5ceFCmXp/bZPO//jIMC7yyrig4I1Q+RZ
OR7OG65Nyw5HCc49AplmEFMoHA5cprE6vYegNpevlvw8JPKcFQ47kqpj4zyfyXEt
Wg/XOL/PVZPa4bkfhtICFg==
`protect END_PROTECTED
