`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HHRIsHAl3ddNtrXPwB8cAcaBEpk48L3vjP2oLGnwhSeOuPkLgDoOvisX8GD3RTPg
DSGuae9I+qt4mtPvkX2KjZhce5Rh1ImKHn6Pa+s8MpXOp++M8HAFYE+DATli0qUj
D+K2F6WpLYnjLhz/I6nHtFRH2vHAZ/9DfmgRDeDl/QNcmrIh4RoH6udobzMI7z1X
lQnIiyZTklI1Egaz1rwmiQIuf9HssBXgkCjP7tgzwhIyvhpythUnhW6B0qkeypfs
jnXBSdlyP2qm0t6AMlT4LiytInz8/eTo7DcvBnl78V832/K1JWyK/XtQaEKKqKN3
oL5yYW6pRnBUtDqUsgSMTk802VKcE6ieVIvaske3hJh4UApiCZ6oVLFjMA/c+UUl
6P+D7zYsDfabePi1pac4KFCFo569OFQgyxPtbrrx5V/VioIQFEBuo8m0ssHWf4fo
qGakaB0qgNWLv2+TR1QKeBknX4kFr6w1kZZ/+piRdVIfQkj+NTtbpXln0WXtV99d
YUWR7g0sBrNoe/15SrEyCbcPZ0pNYA3VVob3T+k83ALDC0pGAYOIadqeTP8MWw73
tew7sug0TSdG8AOd5BrhSfwkbW0QdqkQz8hv5Q8n1Jn2rUX6JNsYVvmgIDJAamJP
blvr5Kbar3lblWRzhucj4wdIlbVgoQMTCSYp5I32HYsp+gZJDK08C1Hf49lvnqd7
LTrgTqvXZznKkBqHZRQ+7xgWTY5GpEbccjaXzEBJfhwVKCCxeMXMjPdzxlyCE1+o
m/6yDfYxEFNALBENCZ8LeVNCmE1cGEi0oH8y1Xgg9zH0KZk/+SzW98N0zeDHQDUm
PPo9KefoUqh/NzXMaRLus0K5jzR+9y1aAEbSJxh8Uj0uuxxr/dVd8vYgx3eXlfFz
J6DYOT/yVi0JdpxNQDi4T4XwSfPrzn3c4XXNCkBhrwVRx54H6QKNIUjgcFzndV9M
VNXdBPu6z7gSmfMwbLuiYSfKF48g3HJF4Y043MGgWR/9oxEHfeK5lNpjyP65knu9
Owhw3kBGgb7/p/zLVvqUFXYBl2JSX4zVb92pTnhML0fWMUNJ/IXr9YhNeeu13eul
+fZrDF7V6w1dJhkYweTzx6cXZq+vBPaVuzG4hxZbagVjIC5qavckPfR26f37BvvQ
tdcKiXNOBoPIBscktPyAdWuEL2v03hI7Tt0khnB3ROP1MeaK17R+vnHvWGdc/4II
iqM7P98Mo/z3lfVhT4KgPOaEpmLASIwhNHWy/EjKSBHcYvI10KeGb/3TCHRJCBVL
mfVHpzi4UDSe5CD5a2Z1CT+TjAVXIvOmbAIuDferiEQmVoVSt/jZ6dnNJiOT/boh
8qZMKALR0daz1qU5W8ES7fFzxPwob77TVLwt4Zc3KSY7eKBqS6yywD9YBHT22wB8
1BAHnndLEj4boYiWFnIt1G43smxPqGFSNlbYZyZp9aZrZEaMid2Hhn/Sn2vFq/mc
JQaAKhQq8MVboAkQrfzr1G6RvateYUsr3enEhiBrW32L4N5on+ynMfEbjBqZISaQ
GIKIeuserYkhEeDJG/4V3EykQbgQbRNHdT6U9Ee6/Vk8+2j4ojX2VoGpp4/8oeQW
LrUbn48JRHnJEwUJ28fiaF5oNI36j8y/QW4Gy67/NfYHLfxiRWgfpEHLEO76sYI8
1zcsIncpPP6eggfF/kjUanW+dFbkd0xltQAyLrCNSFmcJ/1fYeo6oi4hhBMayUjG
apCE0LELHUI7mHWKiTd55Bs3eq6mGgat9HnZ+AMiQ7cFKmPU0r1zomF3yLjmvyRU
fyVAv0E4ni+lfZgpOQu4zrG/YGassL6FTp4h0PNSShf1a7em6LzY0EF8LM4f2SiK
CEDlyXilUAnK7qQvyBf1//09Q0f2SGPR6sm1tOz+cExGNM3bKoojshh83HkxcdLr
3sl6DG+rQaL06+eOnS6PpMAPADC/1d2rIL5qjFkU21OYMamnEfypdpI1fMqscnDP
UNZ6fdQfzEhJRwnt6PFz2J2ZM3YZIf42DAlMzdE+JuoFabOGsFJDitzrx9UJelCY
ro1FPXoHs55s6wp61KxddgQzcXykKVVJVSjTMidauIQaNrrTaZW9v7j2qndXxtoR
BKhrCk76jRyBcnwYdiaFKR0o61DNCsOlwfvE30O2yUVLDrvaLMscz+0psy6aCLUr
qHSSYNoW4pKZHvca/EDM14XnIMNxhjBbjYODdrnrrdgeOYmXi5NvrH00UHgKxknx
CVTZEWwuKB84r3kWaRFuF1PwBCojrOp5YELdsn+JCrG6AFubXhm5q1HS+v9Hchk1
YYMUxmAjNmpFYKe53gACOrzxS682rjvNDEhG1Om1MHIuNOVe+kIOvQgLyTsvKP/x
xs1PyE66NDj8a6hJ3tJm0mw9I+rnXoPcu2f9/FAgz7fpBm3wb0vFqFGazt2XwRjn
hQ7Y7vsqgkcq7Lj5AFx/sKEEFeIgA7Cwc0Bi6BIUakCWJhBN+FSs73PPH/d0/EYd
wFfKNfjHduoqzxIIHvREVoQccNWYlxQ1c0KwZmy1PQPaAzYSsr68QixI3UoBcv/O
9lnDY834ShRxyl0EYXGduFdbfgEq9EkGCO6rEyVDNMkKqNvYgQEs/Gb3IaU2QPxu
d1+Hv9A7kj7uDKTVP1aypVviIqvUwYQ0fvqIXACFN/UOIt03CM18fWtLAJTr1/ML
ohCvtn62rQeVwI/EzK7mRI/Sa8vMuKExT3OiywmJchLhkn+QTMULbhnw1O5bnPqJ
f4m0yphQTvBbSdtQdRxbSWpes3OMay5tRLumB654efkawAsyDMTjrIi+xYEwjsRr
yBPubpqnJMhIiDAKdjikorSSm08JCt+Kxrch1bo+Appt8/NZAC1cpGnmABIFwkrl
dkBDqDnEM5d2uLj8WdF4HFdEQeMZflq1jozRFMSdTMzK862FcxhMV9i7VdEn/tQt
aU/Q4k8lL107r4hR993glV048LKRmyin6N/s0PqqRdYF4SXGotV0oLNcnvJQ90kI
9z/+K5WaftOotyVCWnQVN7TiAmHD7Tu+9/h73rkr/iDKVwC1k+17edqNv4fjAd19
RPuHrzOYt1ttMfeagkhaNsdikz6O6KnWmhf9wYC6cDw7RWeWjv9WAXoufJ33zhOa
vyT8n8JOAtaU6lz1fssr5XBge0qmUCY5vrNPeLBu/SnTV552C6IlAvksKcwEoQip
YcN4lfcv+7oP9clTM0DIQBD+y6L5eU5b3ss93WxyYZDdsstaPqZQDzoDR4Y1wbVF
EFcVpvGrb081j97C5am5Sx4i2S4248ExhUVC2SuLW9OWlvaZ5HP5jG5naiZYuOw0
a4KV/hd3sqAWVXQzI52IT2JKFzSvmMwpgU4W+7oFWNoOuq9YCH7kD9IqPlmHwTor
NEwQRRuaL7gpEEnNw1n9tfYD2xqgGnkawrlWk0F1j2LO/dZ+MEE1xNE5VT8PYgzX
NXFNuwzsDGVK9oOSqFDsEgtDMB4qgA/9Mj273pcZ2fwy+zXtFve1KTJyO0Wqj9ZD
BwbPKACPsoqmg0HBGjyNdeUREc+4382IvPUA15jxXuisSAbAOXId7CaAYK24g6Kj
9t4pt+MAmwea9HcdkYt4LlMFvcbh3mGXo+GIQYSdlpu/KDgVKrZ6aO01S/Vgpiye
RBlc0QhtcaqBiiDmu1kY+/UNqPLW+YbkJPaLHzSU5OYPwZ19Sz3rZdxHgH1kiRRs
RUg00/ow4rFEFoRCm0XPiJGU+txx2mTge4NPbcvLrnMLcQo+VdFMTnsK5piUmNI2
HN27s03rwq/0PNYTkuwcpOUD1rAxqygF53m9chK+8/QqCvXoh/WIYMB9KJ6cRHOx
2SOBpu/o9mzrScdXyyFjP50n8tTkskXB3CI8OcMYsSs1Rupu+ZPTc0rEC8eZbrB8
tObm6G3NR9ngjeEZzoZ6O9Dj53nVvaWZ7F8I0pOtlPMtbxf6fBhXtYfQvlUcruIM
7A19+osNiTtdf3VxXQRzNPcGWeDdN4mDPjByz/rJetqL1hWPUckxaoPldy0TlYT2
5wtyTjIp+pLGZGzep9WDkN58kBSvMgGJcFIccgF55AMQFvbUjOxtkFxKLuLOA+YK
Z3kvC/wwfWM2DQLZgelVol1kWT2ITFCPfs9tHU0QF81pHQLSMwbiVKT7FhzU5oSv
JFdU3lzH+P1iiHuY3GV3VRoShwIH5CTvglbYqpL/5kdZdIwXqQws1No0M+55/USW
JSfL0c1idUi+13DDTD/ZxQRvmtYq7oXlzVmHAJUXvISgqdod/Mpn9i5FOiQagFzS
NS7cX0zcj5wlJU4TzzBIpdC2x1ytcXfcoEHbWyny1QvWCMa7j1XId1Ylmmeeo4m7
pI/uOVtvVbdXmFByawhs1eF2JVBeTYnI6So7EL0FVKm7AVgWkTY7qr96wCbiFcvR
+wd+Qkr0decW4e540kahJjixzqGKot8HSpo+3hp6LEc6E385nBzdoQgj7T2pW0y5
2cKhMttNXtu0zxTbggezG6CuqsEU8pRrTuDO/1plgBj0XXMQdgOu30a2jcGY1rVK
ZkubtjHThY6NpEPRdWPGo+tMNdmnx6aDHae6v+0VAvTv+0mrsWlmPquWmDZ/BgBx
gYk+OY+0ddj+Hq8rfqsuBK6B/ocvTyeBRkaNbt/p+KusiEMKU0MMLvzqCa4Hs8Si
qR9/dA4s5XZBo8tvA5EaQ/NV27+QfcbviJ15J3Ep3fnZG0MRntMUelGrTSlIhRSX
ZW3D0sn1gkHUYKbQ4tFSFvptiH+3okZYWIteAAPL1aWJy9hhG388h9cJqGHvFni0
KgfFDGpmyypsTsTcsiWcWRLg1B8xOrUM+JUQKQm5cip9ZPLcMWQr17DHud6goHB4
bmgdLNu7sY6SlpnbYFrkGjADCplD14MGpD9Og0JVeazp4KI8n2ZRatxsPxsSh8zH
XZfkLByIsmZOjM35CLijq97EUCUxP/Y4CDgUBhiyAR+JO1Oz8x5WlKhwayY3pWcH
XdYGhcPzPx5S43AVjsBYs9RJnTvXULOge0g3zkMNPRxqHr5/ot9VOSfvmRpYEUCP
UCjwb6LAvldK8cyUZZ/BrmcUu9AbeS/dTyCde/KrS6U7ppAY9kaYKGoOjtgoCvzn
A7ZPRLL4nxF8rvkaTdqbCHpX0Z+gqgXcOKjd2zNlnIeXlkrTSMeq5Y91CR/cFEDe
1oLR2XQsf2Mm+vbZ4R9zhuuKJkPuYv0PtqHq1fkTM30Zo4bqS7/h23ZFfprKaDzL
CJXhYd1/xFQ6w1Hr/VDULEIWlt2vD3xDY6l/HUKjVJbbZ6bwjyTpPngnHc2fTwWz
S7gotKChuz3yNPrQaoHskmVfu1FSoUVSZN3cZUTVBtps69kFov/2KppJqT4ItH4j
Yt5PYeyngPCnTtszvQrdvwwa3LNfEO+yzmylDJUeIFzB/BCgV53WgS0b4EBYjvCB
YuqK/NAfnKwkMWORdM+FtFpsdoPOVAT9eL42yC8NbdssUUbZGtW8Sd7cwV8/mc+7
RJ7mksGN/tCwXngLwi7s0THcJ5yQhJGaO5XDWNFVsN2XUqfkKashM3YTPp8DRVaZ
Q6B4Uq+Pr2bpGYlGmAKgHf8aYNS1l7GLFDm1WBgqHqk+OUVgtcWrDGuCLmPyzBtF
OI+W32MprP7kKtxpxTyiW0xKx0JRtsomzRickqx5agRPnrfA+1K1PkrODFIOlvRN
HD/d14bjzvkyo0LQYMzA75ivEoBm9Zu6PAbLWlbznZOaDCMaOLTks3foemwW2EHp
O3EGLSywAdCJT6Bj372uYrnhFz8E3Px3hXtpMeNyVz3UVDUVqaItV3V1OEFvHs0a
VGc/AP5gWl2I75XwqtezBMOWqOeZCKXqBayeEzl5CunBlFPd76YFARoGHE9vDT/m
suvinMC4+xiGFFSC+Ry6tjuL/n304QJI2UvmsxeuAnbVYcCNc7o6APO654hrsqVi
3pErG0duVLR4ylxAzgE2I/0FmiPDPiBLmfDlQ7///CNxUOJ87OhSFL79Cr8wQKiW
i87/ShdMVBgznFy4JAKcjWKQ3Tj+BVOZtGr3D8tokcV2Q8Y598r2rMM3PardgZm4
wBKH2yDM/eNbTW34flT11FCwOJV4bRzTWtUZQDnsPRxVTvk4POeF+gWadCzHj9Jv
BI7j75AFubN9WPTt92l6H2nIzCKz03GBQ20oT5cR+zhK1LMSjw7Y0N2NxY1eaqkN
Cgodv1kA6oX/TyhjH8mTSyb9raP72zOB371xN/Os/yAVpu1QZyj/YBytFP/JjUC+
uEulqvs1nJ8NxKuy5iOXyMqcQADP1SzKG96dhSX1n5SDp1ruRZ6iBB0yrYyEsaVn
Wl0BE4E2kfidutwRFHmvB/azWHz9YjUt+FivK+TYUGBcsxgkKJXqPl++/L/9Ra5P
8QTrD1+aKbHytppwTFc1+dKFdNaInKm8b4HYelW7mdNokHhFIj9Mzy/LVpRCUP+g
HntPnUVDmAkXeov50UyL4XLf07h2dXpSmhDs6HU2/nsroQzBYPq8nFezwDFkEmTY
+F82QE1IlDmC8hF7FG6AWY0G+rRZzICohdrpaJtZGk9R50Yk4MZBiO2Oh9EQiWyX
rDbfZc+f8u32q2Certnpm9PB6fXs1l6Weh/SWMjaspmavNo9dxsPQPhz/VVRm88N
eRJgAWefGqEFm1BP0fiBpAJvbq4EzdWuPUz/TDKxekAx7d1WLUuB9kSR8Fw873Mr
pMh38b3xikhOzCUVLPXOeQLhINU+O8lFS+VhoxyzvfE2fxYOyoKh7qgvcUCYB81P
xAgg0FWXa6fDxEzJB2WHNrd6dkL2fFXn28dxZKPCRT3jwptKQYAfCZhy4DDxptQI
ofoLYFyXT6ZaET81pqnbvJ5dc4FsM0ksVYhYjOkxBTOETizX85WHiEbHES4Q5HYJ
/XDQG2gmKMGKCyKgRnGfBUdxFRk8P7c49SErMentN/2pY+E08G1lAxGx+wjup/P8
nWOifQP+ymXaT/VEhchtMbW4xzBZ9dSpwQwb17YeheeH4OFrFVxoRQdmzu0Q5cI6
66f2Xrg+ZRhjO0yg9VNEl2H6l15apVpTDsKepV+g4hy2sg8ponEQ/dS39dqJuxlI
mDwC/tCv4yZUja/z6NfwcWzUvc6mpSIgvMTorwL2nNB9nu5nnI9je+9gxsvpZVYU
ukRLLgHsbdH+a1JgM7cHqrfOflbnRjNSCw6V2Jg5rjTKiuZ7wSvnfhHDUM+bMOBs
lrBBwi1ye3znoNKLIyE5R41Tm6HSsMgF0clbFpgn6Ytml0Xv+p99BgvjBMzOWIFJ
VgnPwVmbQfw5l2AZniUgcQrellYDufH2FMXzhcV7+5/iQLzJ4Y69y6ve7as0wzns
yeZWpshZJfEb3v280VraiyGNnMptsF3LjYeeWpJ2UDsNG1YTf4eh87fraqQp7nta
aZZDyf1KchgHgteCiMH27HU3vf06uMWUkGXtf4jHoAi5VimA2vwUro5htSQgw22T
JrbpqEPDu+NFYuL/XUjyPevJgRlYUWQHGIxJivrzJZOtAQC0YUlMXFW8mJjD3Siv
Q7NR6B6Fl/uTGqyIRE8Pd002XufdFrLYeRehSW+p2oX/jnW8jWn33f3vs+LQc4rH
B2RIZJ96yxdipB1Oog/+O9OxTxemgDcLStO14IDwiYvo6UW0iEiHR/eP0wezTJgM
7J3RtP45XEKOdnPA3mwCz6yC5qkW7Ee1YbBkob528Tu6Lzyg1rKAIU4Z/pnZMtG+
PoZi9gYuIKLsPLA9ZwAXru+pKgzYWXiU/dThzLCPTQsFkpKGeX+F9xSSUEk0Ydgb
po3LuMfJU4UzDY3myXxmkkOhouIk42xMRfa0iqsTAaZkD5qmQ8vtDg3XTvHGGPOH
B6lvT/wyIjCLERw3fwM00TxnRD/203JvEucfcYRjA0VZoENilYF4BH7SE6WsHeg4
qrQGC3EWVt9hxAXrigwjiWdDHqe+SoKXVw4yMow7qDv+fzFZMBg0YwLH2Rn8x4VD
l7dkNNv9MTY1HjzaNHa3VyPu/tYwenzcsG06U5BiIGRpidZPF3v1vH0AYQ+sc8wS
d9AjfzEVR0qsAQ585IzgCmqiVRxLSUfKnIorj0BwQ2t2Iesdldt28/lc2bCIGpEw
PtTmWuAZ8YUxOBgG1eXfj93jS+1YkvxAyaLQF/vZbu/ESHUT0KXWXkGD/riOC1FM
yJOJ/x08jDqxoWsrenS5JiQE8RDdLiUTefytrRmREyfpQsyB9abege2BF2JjKwLQ
R3sbVtkq8YpTpr81agcz0xNvXlLdJp5D77k0/z3y1v8ddPz2MP9YXHpMk7k8tf3Q
GDQB4ewRceSgedadgr6YyexsyPklmLhwU3OVDK9OOBwgid7bboQ60H6UwqsUHR2I
7+Ivm03bAOS8zTaEPZy+jBU8cFSS2XhTCPjOJQ9zaJLQ5rNMqt6wn5Zpqc5MWBpL
mxA4ZnOj29/NUeISbcCWGux2wGmGMCsGP8vUkzdM98Mhcw/qM79w/wrGmQ7POKIW
vkijpo/YIvy9QnPzwNlBlNMFMws93Nz2RcBaOQz/TL2i6dG0c48iKRyBG2bmOv7t
cTO7xnkWAwHssYb8pELRGI5KB6PFDnenz2r6H8bMPgiNaB4pBJYvajc+7JHb5Dwr
PrKtGW5ELgwVAlPTwro3ZNdNODgKcxEzltgjH7+RK85h9do/cfRQWUa+5f1IZd8U
6UZaACNjgnGy5t3UVVVYlhAcH3FHrPM8KRo5bYlbQFDIsssFpUNE+Eud5h2n+TIF
8fk/RhUfB/+aE2/IT2MNM/xNzA6vEZ0v7U+Q8+5rCy1ZBOs86AqAsUy+VSVs4Z9E
qtJZ82zwRQJ1o8+ldagDTEUc0p+/iA9mPi6BRim6LN6dQIQ3X7PyuXWbNEwLSmh5
WDMQCRbF8wdj20IbBdnwsx5Ad6KJxtwHjQqHyw9hSS9aPhP3T0ogQ+PThtU44hrm
oQscs0QCxjYn4bGjreG2kTwIDXxqC507F3YhgXdsg1K49wT/7gZMTRqfAPmMwUKH
AAiLhOXWFVQzsxgjiZoEYiZG3r4WkKKt2qFGqRfS5LgSAjWZID92+6Rx4uhth9M/
YEDu8FooIlOvHlPbcoKq3meiMNxf/q21p1kI9YJ8FS+LFv/1H46aHjAxPS1mKeZh
L9HnsCpNYfLl5ROxdj7d4PjncJwW+oD6PGictUpehzvxw3ii/wYDIkQaheawQ0of
HJobnrt33eZumiDJG5XBxeevmGHDsfg3vPj06onfyn23MgBKIDnThtzH3AlfqNrp
Y4d6655esKiZbQtgmHq6IuhFrkltBM0MytrjOc3qZwJseNzCeN8T22hVIQY2crRL
z0K/R/jzn34flNoRuieVfjK2Bx/Obgs2rcwI4k15B9sa0MKGIAm/69GMxE1RiWy+
2ZNqk7QPTEy6x/cNqjE3fw3CUSdpcSG+O+Y2KysZTl1wsT3TduxN6CALXjYOI1st
hv+Us2aa2PtWmmhkslP02FgXFX1qGIR3k44JRPNjFBcgBN+uitgjeCu6v2sJCa7v
vgnMblXlqPrHXexM3zd7fq6sj2r7vRmbAHucO4RjX0ZCfcgIY8nkmrN9caHDI79s
2wJtqy1iobLHElSgpsJMSdrvB60Syn1jXWm0fCac1FwYH8y4OJGYfcmmGJyXZ9ZS
evKWmm3k97qZa/wNWyZ7hg==
`protect END_PROTECTED
