`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SclqFGiJ3ZJKbhwQVDNdD84SBResOzvCPDyGAWPzLac93EEgkXPDOPFSnxZer08O
H3cXBZ8OAf+k8urz+enrVJ9o9gilANfYprigTCEAgALbdFsLEDMK3rKjfs9qMFPs
fiKx3wdED/g1DQDgnZ9vfHcBxcLGyBth+62uq6qEe70solzWgvIMzSKAmTuMEOAQ
rDzQF+hTL+EtWxWjSyD6QtwSBa7PB0vNdyMX/QvNQ1j5zJa5JJZK0VlnOsRWabuJ
Ecb+hZbDtvZuPIzh+hqt2HzBsF6DLqIByPLH8ZmVFoH/v1B495d8QOEWVJQeEsUv
EOf0GISTnjy3SZq23MatHCZyQMfaxjzyaKumZZDwNxd+RtWuDXKxlaXpn4V0prBk
Pbl04/L1rDvjsED0TvKz/7evnuFu5Rkzkg+C2ci6BNrciPCpyjCgEpu0vPyVXU2Y
H85TX/IO5TXB935Jrcid+nZVglFoqGso5dst4MsvMPxvNFMXIio2qdUMasKrqzkX
SrKUPIecZOMDZQ35Nlsa2UAatgyd76VNQZUwkUmpbm1HaCVcYhvx7pFpV2MXRUTQ
ZNr3V2CwEm39C8aN2cjCKt8fAYZwXWrblirmUkhKbxZElb6PlMwmbH3mMRCIGGsR
LwNsx9O9hH8Y5KNdLVAQMA8AONEu9sXUqgf8r+1ydbTsTl5y+jE3fz+nJJhWn14i
uaFIpTR8u7hJdCub7r4imxUMghO20tiRSOMODqIsoC8mBwozMdAUsLGBKbHgF7vq
UH1558S7llozE1f1EmdgKZr7qKtE85v0Vg0Ni33CIiE+XRhD61I/s56RTt6jPNb8
u/w69h8kJ5YxPDR/gTf5c3PCrnElizvGAnDL77p1e+0ZQME52Wiw7uaNzxpes8Uh
R4xG0LtJX5TWN0NLthTJcTnU13Aul4EAPStApixYaDNKpJnh7QDWC0GIgtIGTmcc
CuRRkBVXhTZrv0WhWyJaoktA1YON1mti0vlR+zhW+jGO0dfkjZlDWm6FufiORwPx
Xt/G6i2JJ28TkjDpp4BFrl82cLnuauLF2ziDOcxam1wn+2/awrgiQKvBIToSIH7Q
1BMWgquG/qqI6pJRhtcxBxU+6Xi0xXn/hr2S1d7CqzHIK/xWdn1RbkmTNsEcLU/2
0Tf34QaHLFtaLI/Wz9FJU8AlxfhQMGQ7lpNP3V6NS6jMM+F+IhCJYAB44cyrC/K4
zSPyNKdr6SB+55cdHQIpCpOBTTkl/8zODxqxBeoqAJpqHzQZrjXoGUQHwpDBoKcL
0eIPH0XHbHst+d6lAVtrPz6Kg98Ey2Zp4AKaOGaehoD87S29EGmbYAYAY52+1Pu1
WgrN0xUOoICc1e0f7EEJccFddKiS9Rm1qe8utlaqDrvBepAg3QBbu78bhXNRyu5U
9150CazFvWm1SxpzH0zn2X/SeqcY8wQKeOxGkez1PDqpZ+0lht/PhBSkoObgDckM
7DNEe4RLTptExNA5+bj62HtifQlR/dMCxcuC9INhp7Fi6SgjcC/QrlnREhTbHEE+
SUrBYL0kLupvb0DW/6Hw9cb0ckK7/eFYtJBJw8MlViF9VGccAPmeNJ68chN3pt9Z
epBkEqYG7lLjMB3yxZ4dwdfm7rF7sM8coUN3sJWOMn3XX9vXdXLGTawkHpNusTMz
QXhFsVIwt+VZiuZUEXiDkI1sUiPL9a+32nSQrxOJKFCPbBe8UonfdxsOWDw/UmLG
aiJaSq0VDaASOeFtF2wQtjvCLclw7GQttXvNSxzK6I1/p56AO5HFtuoxFD/wDr/F
KB2qQzl7qrzJnrWea1uIsgnH+u7jrSZX7au4xrwh5JHzvnUeEQ3iFUc/5XT0eZ/M
sQDTzSnEDZQ6OYatLYhnQDJHRCxgb3LBIZUKBuSMRLc1meWj35Nzh8pnLqsP8GGD
Upx1XN/ZofhHCayw2d49EzpwtajYV4zaM/75V0hckwS6L7heZnOleTo1uea7LNCq
ct6p7TaSyY8zgNzSOOU7hEf+sWUlIIoo+Kfr4f4ZO9Xmqy1cOZwShQ6YiTJyCI5E
J9iFD3Sz31HLKaIKFXYRUBEhBBdat6Pc0syw2XdI8h4TLwTbpoRBGg3A3jY5Wr5C
g0AIo4juYlnqBDSw8SU8LrnZAjzII+esw/4pDE9diVK9ojztb9H/PKCADXR1Er2n
WfV+zvTvnZDA6Px0EDWahtF5+j6l6QN7Fwfov66+C/Q=
`protect END_PROTECTED
