`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIZ4PMVzNla0gDUEyG2OEgwt6AXeFi2fo1WogDPWh9Rw3eLT49EWnpGSlZDgUYdt
ejqUIEMnQrOjPy4SDTu67uUkTRPifi0o1HRQ0q0NJs65X4MmvhReTruD7hYb39f6
waqSwhllwmf8MqJRpSKP0KNEUkPbpTDnI6+iKst9Rq39NUxRoTmeIl8NID08oFX4
pvpRIw6k25bbjP7CC3sK4GlEE5JIqBoDdRuybOvdTw/HVpQX8WshvTy4AZLoR7VE
msnFt0oCl9pPqnTbmDtyvLk3Vq9HVLGP73sZb7cPLgOyJD0ebUM8XkWF9mkkpoX7
ayKyO7hJztxvVvYVL/ZkwWApfBFYbZnrx16qCQkph8lRzqyAGiGBAQH80I3MnL6j
B56ZgKaiWEHofScUPLSE787MW3v+FbetKLsYWw6Bv3thDh2gDkqnj1eU5h6kdEt2
SK+Uqc/2ydBdqvpVEed2QnOVAxwNTLHIk51al7zUC5xg2Ky3wMR9c8cuYsBzcWJ2
RbyBvy4sckS5cBeZ/K4WeROUnkcEoE6ttXu20hAwjJVuOhJ925j3ccKWeeEBBvCf
3VtqD3ZRfjJBBTAdAMNKcEC97ymQfve5Dl6Htm4q9u2RcqQl2um2Da/CRpqn9ZJC
WxqTZ0/OXgO5uSJXI3ASmMVPg11JXQybhzBBe061ZS78my2/CfbfxhHW183x+BUA
kk5vMJ2W2acJF9BYqbobCAnY0XsfxodO10sieOX6WHaDajOsqdYlDj3+v5cFPF98
kBwKvw/QDjVi9zs4oHUDcl+yLnR+o+KZ+7bWDpFxkPOpnZZxY8tU4kmLmJ5L4VRT
EBHin7DkrAujBqj/5LtkQk0Clj0QnPdRm+1nR0L+DY7WoxBQZ8zNHr7DztFS5b4H
SrjYSGlyY4EIM/G+TkPxKj8A68yu+RPNMBFaK5SQZjEoWkM7yO8pRIWJUojgzvzE
KQaCUOD09tEMH2UIXSOb6zyhkvG4RxOPJlqSrqq6B/tB+LkFiI5EIsy60ctj4mLV
NYCywgz9nPdCV4UTDzc1ZcR0MGKoIDBSFfOGJqBgu3pQ6y9TVYiVAiImanlKu2AZ
jy3muSbrU8Vj0604fYluOamRszgzSP1RJ5NgCT4a4XW8lgSOd5adD+1r4OmbtYzn
sKDRKxSU/StHO28RNcEsxBG1MLnD4ox7ogJ/EgmJzNWEVdk+6U/CGpR+STFlsvEe
XwzXDPGOi76M+Hsb85Zu0KUMeQ3y2fzxgPWdL4+jy5m13TnD3kZcp+p7qQSZdif2
6124A8r3o/9jWJzZAAGCTLoYeFjKUPrdy7gWxOz3E+KFVBFs+anJXrqaC1/MOJB7
i0CLjuY+AH5Ib81T/s0nE82nxtE2SAFfJKRjUd6mMtXmygYeSQYYaAoD5yn/r6cM
d67R/BBKKl4A93sQbD8B2vD+Yhho6nfYvK5mLtbii+FfYEY9eR5fbwIonLe01mYb
fWxsZR0c4sH8ygUhUp+CZDPNu0j7p+rzudfI0AVRUqgmj8r6Ycg6HOsISM4HUeI9
RvrLM6OgIiPflN4c6/ztLlb8G1SKF7ONaVK7rXanirBor0qAHNVg9J++4kyDLpY9
4Oy4hSZ9vSagqQ4NR1HqyAsrXBt6UmEX4rMy+wovJivyhx3nZU6UaaJh1z8opl8b
sHeCGOqDoq19HAxAcnUhsLYlGunfOqCFj6zyYPNDOFfJUSi44rlYdeMxP+W/K7uB
YUJpuo8ktOdQeXToVvbsmv7aI+VjVr3bbJJNcFJ53gJkvTQ2oObl/ZDQYYcP3emd
9FyV3m24CpPe6qdHI8o/BpS9GBg4qq9FgP+xMuDenZQ7+hzorbpAxiEeKcFk08uR
4+oG9WBmB0OVGE1bi0l+VuDGLbqwdfvVPJCegiZd98QhmFYFM0RT8T2UfmG9qZFC
cQGTysBsy8NN4jvbVe1J744QlplLuUO4YU3LpADvE6ALrOmCB/A8A4tOVzHywFyg
QHWrs8yjqkFDwD46m1vQC8wsjo0aMocW06vmjf2bmUyK2Me8II4G2MEiByY8aBmx
w6mKcu+hcyYhKgQLL+BnSYkKYeyJ+jqoSYEmub5NFsRXRaOH96t2HJEeNA7/Z+J/
4drvRJW1t/PmBuX6Q2iDJCMcFzv8BtVwOSodVBiqsPrginyvDnKhTWgxfKzPJgiG
pWJTGkPMb1FEUZdx9pVSiITz7yIldDDcmBqb2u6vvKXCgU8KUtQ2wWD7xKrv4pod
FX4SIESo32WnqxphLCB9CV/fKZrZa7JLzq1PEZC/V8U3FiiXCKXi2RTV6LrBkR1g
`protect END_PROTECTED
