`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ip/qtpObU3nsPxbrtgrsZTrR5l9EYylikhu5vFB5nwdJF3btrcl4DnMHk/ZYFS/a
1vuWt1589D9KlOeRQQlSMCi2sINRjYcRX0loLvqVHdzzx5PG4tijs5RusIrzNOgG
ESZ7zSBkMvly4QFjmnS0MJ8pgWeO2OlfXHur7iejBkYOVv57WKrz8oV+j09/NxMu
mKF9/prtTQWfuzBnaoTIQ5zpnSjQEtpi8r+wRgHs9P1/v8D1lYYNzvF+BO9ItMq4
+Vy6sYQjUGsjjwLHN3S8SQG34RJt7wYgzTqlPeqpdPvJhbl73wqF6zvGwVsMN8lc
8hyL3PehBvUsTNQbWWgrGTn9GE8NYuZCFuqQf1nS20EZS2/AJkpjmPkOka7l6bt3
82gyzk9N//AGk/BE9yIcLE5n40xzP+r5H+9dLXA6fY7NCgmF3uwO1K7Py9sVWoHE
QrXa59VME3L5gg6XEa+TkRU/5a9rGrpsNRhlRgzwPX2Vp5N9E96RRXo/P+3NLprG
fsBQpTboqvP/GF0cWbV+M9fVF6q4lWqaeJnXT7uo6neOXkW8N6kylCefW8QZEc0l
1blbb4ZKpiVsbn1KZmEWLHF3tDsLiSfJZNodchpfp7xkAzf/ZxkftdFYbcSOsvY5
7h2XNwtwN4OzRGCiblYY8eFJN73+4xnYQ9V4zXdAGOA2bGHpLknpusDHndKyZ+YU
AeKbpFr66cSengRYvqnNRChORbwm5kMreDZv/B401VWEgnb1dzfQ+aEaIxA0TeKa
6TKgt4pBhkYkXmH3FF9oc6CSDy0qjTDWAXavFCxZfSG5KatIqYJJlhatLZGW7uXF
DMERFdFUUERX7HeoZzrS02ZkMZ1Qjm3lnVtox+4vBUfSnVEyN/a26KEzL1NwMVli
P7mTgqTufn2IuBtWQ06xAhailSxZNdDQf2MJBwyMm3XOUeeHQ+86Gee2PCpb8dmT
W5Cq0j+FdC8kVtXlG3xmXLUrLV9DQAhLq31Nud5sV/QOor6Vm7yix65rbASpzsXq
mvQHtjMVVPOkvLBoaNhTNlipN0vL/KghmY8CVewUA3qMl7jSC4uIAHUktz3eiH+V
TiNRqUi9kyAoe/QQyeWp/KuRLSwBj2r8O9A2r0NCy6pOyornrFJkZFbtwQHrpsVf
Lx2Ri8E/iMGftDey+evPkw3lb+sFqkXOccL4n3Qn1l4=
`protect END_PROTECTED
