`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kt1Q+Kqsac0qSVtDHVKor4+VxTENgjSu0Lr0rLvD9iqWWa01n1KgmZPm9lE6JR+K
Vz5Zzf6XXdC/qE3sECsowyBdTfV7+joQ2MD401uj1w1OXuYECvNxKxVCIPXoXlaG
B8Z3Q4wqboxQ36sGCAuHgkiOsXKU2FBHa0tdilVAncYvC+Vya/3lqPbvafO4NnOt
/91AGHxQvw7VDBgjni3b7elEbYDF5dF6bRygWp8+kgjPNy/YL5Z21bui84gdRETI
wSjwJJOqKx2RvHyhP0vkKbYz82Yb9MlqxJHx7eEFUmXsQaemPv7t4OJXLwy3O/fy
6OlTt8X3Ly27y9l/dGh8kp/ZRPSzTcLdcUYQVt9xSWg0QMDzgYuCqU/4YLE9YXZT
fACPIns/b+Zwja8SVKzvoQ1KqywtpB5v0CZcnzLNZiVMOrkQZ8sM2b39bGNToLdg
FrX9kRNWQTNhHOElqGRA1odwx8tZD8JmZFvlGqQElJn2kv45G2GIkneJYHOK0OMp
VUQcBX5MV5D9k/MHgMtgASBMAD6ZwBft/W9rdtKm+LN+wG8bOy1BVzM49JunXHnF
+UwWzpUoOB0w2y07iauVyDNUo32lSBlzpTXP+Qg2HmXaLOba+mg3plsDs2zNopCw
Ihgv2BQVRkhsG3CnZ++q2gUrnoiNeZ12s74Ug+7EHn1cPjj6QPipvj12fYXoYSD8
1ffbnWEiArR+ZUlUdWAkoPBru9dOoGRNgyzafLqQgLAcHZtqK235GgIadM7Ywt1X
8e2SkZv+EIM3LNHWONNJAP/LR8XW+GbQRSN4XLUDu9B0YaacIc1TYuUjfUmgUaR6
Ee1wZh+w5GwUNKbrqdzgGG0NUXvasdr5POtkeLCVttjwXa5mtVzFN8Kux01duKrR
nUSuA9dxw2sfw7MOcMlf4mWCqougO5VIdtqik4KsoMUW5r83EOgXzhDKdN3vmaIG
/sBv+G8eW0DljriCSusv96hypM+ilOtvLKtd/vx4WwzRkxnJPNervYUacbKGc/o6
AjW9hAxFtuW66aQK2nhWrn0fGA6dmSZHlvpnMgFTZRUyEjIhLEEXKJ5T9gdYf+Ac
BQtZBq7YChvVdEQRqU0s87bDco7xlZW8hm0v57UDPk1TQt4JhfzlwzvhPzzP7dRj
by6dHHMFhRxcmPquoaGAtRjPYS7p8+vx7/G2wqK153TKtagFMxfVYrhT6XLkbyPq
SW5dJTRDX1M2u9Te2wvTtDtseGMenpTjyuiUxoMDFPxBqmXZv3EA5ZZiJH+/p7e9
`protect END_PROTECTED
