`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHNrXoW+tceo+abV4fDT4qrdPqAf4IOB7RQVgDnuWNiyiVNBYvkJ5JVMihVIpgLh
5f5gn4rOR5kIMcf6jZvOfmEUKPSE9mKqvSutuuOzYfdKi9RK7nnuJzH6PEn7zJr6
YENeXLIBblVddITfnCXRsduOfFomwsdcziZtcGdq/CFg/w+e6be1TZUZDlHmpVdx
Pp/1NOAMfRPDMYq1ridYoCu8zdCFMrbSpF5M0ytI629PigJMJZo5KBRs/CKEa+cs
4ba8ZptJzyhp6lg4jqS5aIpYUWRT6eHsa6B0uyTK3b4=
`protect END_PROTECTED
