`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MBNa5hDjA9/sDoegfShFnUI0x7TSFW87X5FGv5N8GLruv5nbLavttszNYvzmU6Ww
XtT34szrIHgCyOzukbx0Obu8aUTmmD7qH6J1xToF462Ds/z7HcAihdnCzZCXr8MH
2isjDBxofIfAwKj8rHPeMn3m3OEAk1eVeeToLp3KNQTpi06U6Ph+iAIpqwZLNw43
NEy5O3rSzyXDp1HXnKOEZRvLjDSCYm08w7nD8foo4Ggr8nUQWR8A/SZCu8qPpKE1
XkfcnYMeKHoXWCK62XxM0sw3bmQwFiRJiGfhgdmkCCYBMUl+/vg/DerDTpPB0zKi
Bgb9WXc6J99Zn8hxeppS7jPNzBL3jaJmfbABwr1qtRHDErJCWUz00QLCWOQJzj5b
+4bqJnYhSw5UqDLVgMTo2xV6edcOT/WELDkMW2QEyGE/5Wo6qiUWMB4zkmuZa0P9
O+dJh+wzCvCJLHOjgccuH1SE5YfLedzH4A0x+p09GUEcj26gExX1nfD/p+ZOZRsm
uXn6sCSYhI4izZ3TfabKrhxqpGt8DmgQj+9CYARlK/dKcisqEH4SFcAuwoBRIgFM
/M5YoL5XLBwx3BZxk1GoZKvXYf59b6hgvWP645Ccwcg=
`protect END_PROTECTED
