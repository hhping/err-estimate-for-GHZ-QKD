`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f8q6Lym+bQWmaM/prdrNZHkld8sccN0mIL/zqUvor/viitUcKho2NT16leMNYC0M
VCQUsnX+EsbSq+YS7kezUU37naZXBoLYQjU1lC6hgB6rDJH/ucIKIjfKyR1ZoYv2
9+3e0FtM/KjEa1mdT3XUg268V7p62MFENgX0Db1Ka/ONk9XhxDct51P+3ta5pB5L
3dP2qBTTIni6SDf3kiOTSn9eNLo53WYKdlCbXbUrfYNjJLWAY1QeAjSpl9RINGN1
aCefOGdp0pxYdrXxyYCvoj1b8QWDueHV/75TC+HIx6b+LvvVVY8HNQTEUd6qBIs/
WUHxO4lT8ssbEaImMrv/tb80wcxVyJpZB6w/FT4FoG5tk/B16vO+w1B8iwuAdibM
m39KmChbO23SyCjZ9709HEh64aRepEzA1nB61kbzuqgZZ4YnxZjaIg79kAydGV+/
9dQY+e0dX+AY1DOLFFQNmGZRoJBIeEjZOdpmJ/3XYgoW3+5GCD9vNkkRvOg6x026
lendJwjA5Wmw8c40W24pVDBsnvYN3QLBrsw7ojr9o3jMM7abvoPS8S84MdrFwI8o
PdYqXfgqB3H+7DXh1Y51auSaCgcahYkHHRZx79Ag2+WY3KH2+f+n1uEWPS5f0opl
RHR5SQVRnRUK5nHWu5ecit48fEzO0zcD6jd5dErcBnB4h5rJVGGr7YZkyyBvhQUo
VmQd9UOxhXKQkjmwslSxy3rIoX0W2cHX0LLkRUiIrxR6oZBL2BImcm37IC87GGj0
CCyI0OqI8NFCROzgh5Awzw==
`protect END_PROTECTED
