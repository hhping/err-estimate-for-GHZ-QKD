`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JVDMkTG3TpfUXqDOfvmixWYw1PwupucQ/IJif3NHhDMkHgOpOrt2AbZuYrNpi/E/
jwksxKTuTwiyuWwglgCftd9Jot/ttJFN/YusDFAqrgKzuJnmrnzkEs6pBEyHe28M
rMk9CWqX2nCc2h56AAsuZWqL4ZNsFJL05iGRtiFjpPKvAtL43tvIPWL8qSqItusR
p256/Rt43b2F/WVcm1C9ni9FePMfuGVG+QmV7+YI+krnFQfRoRNVH7yNwJt/fvYV
7OPqdMA5g56JivR5b4k290zKXBN3/asR0NaiMHV0GHVPkpM1p6avk9GDPZI4aeu2
BFaTTiGL8k8e/6H+KiHfd5wuCSNPTwUXxO9kiLNsXII05bqYgDF60p5yZ0JscwPs
R8qx8Fcvh03XK7WcL18pKwwvpxh+Zrz5cIcfBdAliOXiXZ+DzdKFe0NsnmxFC0Ty
T4UyjVTbp+N2cEz8cMmofvj0sKxp1gdYmbAL+hTWBrD/fD2GTzU7i/37WVHMWBoU
va6KhnXhxHS0u1YxeFBSdivl1idqrhRekMTTTRidvdxQirBiB4ew5FByX5y3wfQM
7kBQdh6RTmqXxFz3DETfsBUNA7x/vg6leIhinLGsrSoE0e/MyhjCHJeFpX9u7R14
hxh+/thU95LZnrSY5q35GNUWRzvTsL6XUvqbgfANbBRP0HtxKaKAQthpDh5TBokv
Byqz7HfzKzBkJyU1OR2pLVZO2yS+5GT/A2eTe+RT1VN0qHjit286EJiUY//aKSXE
U2k1WpfcQad2GiK1e8K/CHLcWR2Jiak8S5Z/ai5uLTjkvUO2ju/wuJNJQzucIEQe
zWBelTOtGJ4azXhor4XkBeDU8MgQZ0+LLDOU8gel0Ru0diO/8RAZyXTIYVPC4Ddi
DhDPETkfKAgMr40gIAQSIeMwu3i/CJ681/jIpt83nM1py9g+0Vt6jtm5tNxGCfM/
F5x+XTUBeiqdGokschQD4WrDotqg4FkreIyqUCHq0GdNFCrJ6Mt0bBIxuG59tq55
RHspZhN/tfw6P7BoBaNckwhuPkV9XbxOGozDfkWjL1322A6wCms7yOzERNn2FIiX
9ysC5C0P2+dLVt03y/hdi2EvsYE022kx0vD1Sxcs+E8eHPF7TjPqmHy1vDfWrK7l
9fRk+VtbH1AxUkmELymXuerFULB4ouBuEPzeNg+Wmsb3u3Qx7obybzq8xTwQKPm+
rkF9zTPcqoHuaSoyN6IE/ZfaQaa6RQb1STl1XuIddoFSfGcpSobHMgP5RAztZ3Xa
bnE899tZGr2P6JfXBR4uUIbjIn9Ow5lu9W04VLeQZdI=
`protect END_PROTECTED
