`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JRWYfRC6nyl2uWHlFarCuSPskumWR1Jfzab8zZqURkNRVj8UsMM61VAQ9NQSCfGA
dQ2VzxNaxo+4+8gBPVId8B4jjTAp0emjcGBpFGEGDZYntj5rLJ+6jDu5rzU+tWHQ
MTssSZNJ5sjksPmZQP+3WAWUNQcaCGa/23aBkGvCyusrnW0/hUhCJno3BbSef2Fn
OX0TapC2ARx48ExHsV3pm+o2K2QWKSf+jQAgB0TYSeD8PLj5f2ey9f8kVY5etSxH
+KGr7xSZCgV4l/kyRY9dejWoEHmDjI5QqzqyK2sFPfJQ03ecD9F4N9I2hnQ0lZGd
D/PTlmVnomC8njnDEQnhqSli/uZOVlput3BSwIqDoJDygDx7X0p2VfFvWIYW+DMR
ETQaZbqN5CkQp8rSEPATE6ib7B371bGtvoBNJp79h92gXl2TZH035uoU/2KTrH3F
YyCA0g4SEVPIbAGXF6189PDQV7MwhAl+ycdMOBcBHepvia9PPYRFgIRaVjCue7ty
+ImBUmMNNW2/lPmGLjTjgiKBWfCJwCc/HrMsBJOALhNPgur0AnVA1FCNWB5jd0GN
wD+dXfvYL0mZLgKgUp8rOEooRRvzNURDzFpr3nS4Wor3OWJiefCzo+7u096uSXvj
pQx9c0zHIOjzC5WP/VD0iQ95+9ds/VTdQKONC8Pb8IgZwTu6zGz/bTS1Nra9cvvP
5dQdcRrKZhNRErbtI1DIa0ocJCPvDW3bZWVnsOUEk3F6xSRTxGDuvPvGSfTOtkUX
o8C4EhMaQVwee9lyhG9viL42ygr7Wu+XPejN+DHX6MUpzcRPyDt+vxyGK36yVryu
rrWYwCO4ruS90xlVOwTdRA+xkBsXJn7MOs2j2rcSxL3h7FPvAt6zKZEDBEcL9+z7
eLY4T9DobfC4Ci4qki5G83Lz5GaUZnKz2qAQ7xlA2g/2G1Dr9nNXG6zhZusXtPA/
niPKGuPoYpePYTp4zAhkX+zfByQkgDJdag7ZEuHRO8DheEbGVeEBSA4jxquzapOs
/Ib5Pefy1E0lzQRfdpS8sN1AzHGvEQGuSVrzzXnP2cEQWxQV5R3WA/XHrKKFLaJ4
C1jN//AlLQdta/TSBOKopg==
`protect END_PROTECTED
