`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpTNnjK8b9bXK9h+epb3mGn8EMmRZZ1egnwDsykGlV5yeGZrMKXDYn2GH1SS0XjD
TBbvDoUMuqmT8KWeEJAGrzz5JA802f7mBuIqi89sXJt+IT/i6nkMfBr94T/+omGN
JfW3wgtl0LttPaPhdt16ey604CSplM63nMvmPb59Vfty5qYJeTg4A8BPG6GqYUBF
gKUf/KRDq1eSUhfisjCwkqeyxaKXthtXLPeliu0BKiU4Aq9GSmxfQK8ElDWENNtq
HlzPDsot0Elrs79bgS+hrbrK6KK9YDmCRHbN4lZ7DCi986o7/MG4DnXqit5iEXcj
mDIdup0t5uZv2SZsDv5dq1Doea18d/Ep4Rk3vZdjs2xJh1/t36SUthGTebCLgRIh
BiG3gcd4Q3y9+2kvOpvzx2FusD/VAp9OppZUtyZ4au5Cs8oKDlsEx5f8clz+DkVp
kA4mqa4h3IicnEmwSMZ2JMzYNw8GPzSu34oG9phl42ZJ97Ah/WvAyWNPRQLxapdE
4fB31xjll5UqC5XyEhVoh+ixIkGcBMAzI8rI+MsaB3YHpluArKV43TQuouotsec1
pt4rfyc3qwGaIY/JNXR+0DTnhGv3vMKW3oTKW3cLAG728HHEZWjAxT+7OiYqXbn2
paQ7CjMw0zp5tFNw9L2vqY7bEyYStIbZmHQVVwiv/TizMPEHV3OxYihUpKiFZ3ur
eQNpfeXVyUGrM5dNvjwKFhOlgbyCtRSxwY2R10rBc5m7Wy6cvqU+RXBiGwU49gZa
H/1N/J92Kcw85IRmR6U+dUPAUS5qZA3G+Vzeb9hlWqFZYDtL7N+2/EQ2B5Edkg7t
GVzZwyj3nMrHM2MW9+JRsnqrlec1/9YQRv3IQdxgIWc+UKSh7yb/5+Ked3uFdmYD
FuzKeGZqYisA7lqv5BjnBpIiKnFEyq3JjU25L8JHjIvC9F5WW5esytrUXTalYffU
Ih5soCkUJiUwnpja9dOw2MjLS2ifsEYZTawr2UJ2UsNl0Gy2OVNyOnbz0HJg073y
4RsL9DQPJSBHkQExGf8ncsNwO9WtAq5RKsC6/5+i4EMb/NyQ+GC+rjw5zksPcSWy
CbUANLVj2xVjSOEnCGKmdxyiLWGc4oKGXIL4gFTy+RbqLPIOO8wXCEXPe6eRA4Jb
yBF/w8i92JkGV8hUkUI4lD+6q/LIZkdyzg7FdlIj4PpW76zIyAofQsclX0F59dl3
2Es4U4xP1OFx/3Q3Opf5+KgT2A84WCtK2H4TcQPIlI64GgQGORssly5UaBP1c2e1
Gu5i3gvLIcHfzPfOoFiNyEE7YywjtnYMYPoajY9SGNY=
`protect END_PROTECTED
