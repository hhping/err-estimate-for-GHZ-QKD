`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBbZbu1jirGaHXeYxHcX8B0h8c3QMX2uzBZK9mTwdwt336kDg617QlvEXvZFsppw
3bCA1voX1Zo/Q3hZIfcdcYyHRMpjwn7C7BzzVMDjjegw2ZYu+x9CTaeuMJ6eCakS
npVXVnPfEvtISxznRGRhaIhRPgmItN6pWK8iU6oMzUyuPQVKCbdZut5NTxsNFFEl
LIphxx3Xv/QbhStysAq4WDDsB2ZI5HsMXB89Uz06daijNugw2UKw4jtpS0bdIQWo
85D1U670UOBb+ZlMdTWytP5rP5957iF3otDqGlJRlk6mJ614YHredGE5K4aN37dw
U2hdDYokMEoPkp4c7S0Ms6i97MFjiw0qFoab08zyWnNcczrYO3Aioiz2myyc0WLd
qV7IvX4VfbfMNnQ4kQJvCLPKrmCn6AFjQ2ZCOmx0ja8cAb3lrgPUr+Vfu/QFBuWM
ikSXKRY4HV0ZWB43nldaGRdVLSWd5uT2sli3BvKlvTuY89DYAvCQ1Lx+VPnQTmkt
4mP4V6TqAsFHTQlAJFbBz13mx4kniTTPsL1P7zkpBlI24jsXNFDfDRnJysAmx69E
CYiPe4nWZrKzPx0d0E5VBSeg9sRJlm/LWc6jE5n+dBbRPw9xu0Vn9zq4wnPbYurg
vk/q1DQ+pecHzDrrI0gUufI6hA4GLT1zBBzAgHLSxa4RBXAYmafNUBc+xsGDYVrQ
sjsp6zqLSBkXGowX/sii9NH67K/o6gILZp4fRGMJEBOAHB2UW2yBt88DB0P1PDP/
Q7A2jAwsAzVan2cMrIYsCPXvSndCJr8P3YnAJcnPlx/s7m1d9bYtmmjnX/DmA54j
pJ5YRjjaEhPTeKJfLKTMP5pgN8OehHYDZIlx/pnBArNo1bJw55XXQyVwIewzEywf
uPwbT4OwIY+DvMOYYJLZ2aqy+4EZHJM4ilrSU8813QQFUFRjO803G56NUkVZ2rKx
KW72fd7Q5A/xWpvntiIpqK4CjxZoAhJw4rq5mTaP0khFlIU1SBNR2zUQlEoJk3BC
S8cZjUXIi2xJpfD+eTDSF5TkIrnaPLR7zJ/gKSMKDsLmtx2NPH+vWdrQ7N1Jw8Dy
KG3fut3jNOAJoQwThWh7VrnmCrzg0CAEgYeZUhcrf9HFKBIGaIObwGQ5+pWgM/b6
ajxKwmLSHXz9lBNqHaFRjcXKHf2KpuwMDA/67EoKur1Iw4yaUPWay3vN8g3d+X3V
DEXMLG8MXXzVM+yxjnraSHkZewGVEuBt1yQAal5IIp0tCvbzkK6ARys0qS+tpPq5
mhJlqiv6PXH1IUIgL2sQqHaQSJR0Wp+sF2ZrA/TNV9ni69oiSSqL7WQk4Fx0omQJ
7FEDARy1UigSXzx/JSBxvpFohPczS0N/9WcBmNX7JQ8zVH3MWZhq4A0eHZfb7lg2
9nhvRz8NLQGJRFmxwJmkSD0vkpFMk9Kgnn5QbOjgSyq6uUo9JX+fxlUsEYTEjqrK
mFamdwnOYYk/4PVGfH2xFNAK6OjidbmAXFMgE9fodhOA/a47VTaanTstwZvbjrDG
gZQAhTwFqy/6b8WtjumccJ+RkHH36JckyanPiZA+c+eRgQ/1bPdQyF1ZE6DkUXYZ
pzLyLYbEPj3SPBKI2vY1A9tV9U9k5tjIzkULGKhDwx9onvaSzq4RnDG9Yn0c+5o2
sXyDQLWTDOmjJPLCtjBnoW9GF7MXar53arSt4ECq8T/YxV8uNLywvF8RdiJZYZW1
zl8wig4/nK99/YN7jEWStZcBklatZM3mMjnbH6eKWAGUypp5T0zNxZi6vTuQkraI
Q6TJNBPfY9PCb/K81hLdgMvvglf7B6ZSxThNUfn/vDfGLu6JT3e9eAuxaj1TgyYC
nCu7kday6DHZKC0QuYQp+0/n38/iACBtZhz3D9mEUc2g0oJXUKd0MnpdLpwicvEW
ghVT7pxq+YgDhZK+v4+FEKRjiod8XNJ6GYpbM2T6XPI1ueJPW1/SkjcKj4j7Clmk
zIgD7gUaXiCRxVl0g6lMNeOJNk7r08TosBYhz1yudszFYRhXGVnEb5yMv5MmQmYK
6vndvR78kRTCb2JXSyMPEMLq51+u+7OgboDBt8cuxXng/6KSCGw/P8Xn1WUtwFki
ESv0x4zgPtuEQvux6bKaiPiKH42JSPRllzCWNsSNu0NIbb0/FKjQ36DO9OV1zYC+
17r0xUAVsPrQtM2hDoo4+CpCQogLmqCxtzQ6ih65cTxxUEYmUaoR9fHDxxZ+ntaI
JZfeQzNcF0Yho6WEFkaGEKbxgxKFZdXyp2jSG71AuvrhdLSENz+INums7fxVhdeS
qgWAsHg/uOMbe6tGGEmhL2sXJ+ZN1FThfciIzmNfwG6/0COWURFjLmMwbjMGFJLn
PR00mF3NgtT6mlGt7ogxlbmdUY8ZWUV4j0BqzR+jN663hKne2NrdnG77OOfUzBME
2S5E8Tf7U/f7D9ZczB7V+Qwng73rVvAdUWEQ0yUa+89MeT8Bkz2inixvfmP/vyt/
jgnL6YmRxPBpRBNIYoe1Z2f0Dph82J4v37OFvjDNv4QW4iXfyncDoqzuDM1WMuYi
cEj+9lLRjsvlG0P7sEqhmPBXWgKo1VH1+mwLs73mtnnMFl1zna6orjDIgAQajufY
ofl5TmELIiFEsLSyZOW6vgF+U7AoXh0xrzTb/nTYHNgiaIhXVQdjCVJnEBPe1UBR
EbyjzqxzZA5NoNJ+ZporfCm15AnM+mzFTr0qoNXrfrOqCy4fbNi69tqGDgKeKxXL
Uz1O2v+0AFD1XQ8PtLz+a9OgXgm1aP8Q6eHbXEcWYo6v6lzcJ1J29uyyDvYAcSOt
CDhxjrvPQpBVrtlEQpXqBLWh0ydC+szrWYQeakhFu7wXT3jWG+b1bwJepvaDPAa5
raBbvKXJY8r2OIpnoxUyOgLAVMf0VpFuBYdCaCu7VxquiPeQ7v/cy3E0tdUBCaHc
8qN2Xclisw0joY23QJIirqi7VP2LEeYyqUHuC214RSEtdDP64GT92zfqq7RPaaKC
fFes9CnDMtAZwI8Iit/FxBVqUqddd8aamX0vJDrlwhH3lYjhJ/lUW1kCqcu5bmDt
JQY0WbFtxh8arhdoA4zWWoyKZa0wjPl6i65IlCpb+AA0tY939Cpe54HfCk4jacA5
3KqKd9nc2tTPlP9IHnQPM8JQ6Jbg5qMIMO1u3QMFO8fFDN5oVXtIE3h+S+SFktDd
gw8JqxeOG5+hLHrj2RAYFIoVRrojowlfDgIBVbDnsyjdvdhwdrV6UasfEvPTIj36
m+C+BXeOvGdL0kluLDVE3or468JGPPlFGctYk3Wte4liSHHdQDRMHVKahqUCJEnl
++nHth2BSK+GTwG1arVfyjXwDe+dR8QZtLZiboExUlDNmn62JHTsL9pLhRW3fFoL
tlg++VDr3O/ixtVTDfHlLJmFAGWf/xMs+sxgO5dcdFRGDKa3owBGWuXoY3hSJYX+
GYoeTjNxk4/pNoou0l5YjkoYSPLdrSkvDmz91bvpfw12knu0Y9NTlVXX88s8781n
nYnJSMpdChU7f+t7LcjOYi4u0XfxuQ9Zl/POYQHmseL5Va/6hZ+5sn91r8z5UZkT
LmXUZFtTJBkhQrKkJii9qoR1BXDw+X+cxd38DqFgynmxSEbfyyhq5tm7Wp32ibBv
g51PFSjfNupwghdRME2rznxQ30+0kECvItRKxig7FsyH2ntbAVz4cfedg2mZwjn5
vewmsIjQ+CVGtt58stzIYkYqC+eV+/nl6mGY5mKv3OkxmmumWS2S4uscFKaFXWBl
5teaHukweWgL1P0DlGNMp5aahcGPMDwLNKTjCTKWGvSpYxLqIMItnQRD2bSE/Jfw
Ac5a3VHt+LVoJT5j9EawcvvQsQgoBaoMw28a1J5tTE7B21/gHp0lIdtQafl65HWg
wEfNtkokaB+8Tgn0vf/wUVT8ayGk8pdXqSnpTMLBPc88VL9+xRdcfvLZTTSj/Kql
CQcwl+mp2gc4vHXPl/gK2uD0d1yI59xpipmRK8STfXo3OSiRSW6wBaKObQyDZiWl
Eg5b5mwEfREDzpsb9fcjINQ6gmZ3GDTJGqStjfQCsGlPEN9Xqe3I3JqxEP9NDFYy
DJrUfUf57PhhzmMuAC+AWbYVDOM32K2yixRhOOZF4UAiCTe1qwDzdH1v1jbdzA+p
xzvrNjsLpunwtCjaFJz5PrhBttLuSIhcPwpyfrsALdc4D3FqAGCKRW7eZw5cNO30
fyyNBuS482FMZeMGbi8siYoAaReS3ffYx5QZTbO2nQhrU9O1XSB7sfZUMhvnhUzc
Ni+1I1UrU+UPZSdpTn2CfS+8Skj97hkMB6h5YgWk8W8vAttH2y2msxrmAGwVB3Nx
VG4ZfRZaQj5RSQxKVUh0GHIkE2OOVgjAl433drJAwUm2n5B9sFBZByYu7e4e/aX/
bYfONLPI5MRtkpaiqtI4YPGhnEZICAius15a4Fq5vvkusLBr2+ZK1Ep2NDbU53WI
OG5EmkmOlM+TlwRVvxCKliof23ZlorsKHhXgHsY3YfsXcUbe9FRB7Q1T+B0xRlLN
Tp+wXFkQzedmZB6PDf2yOctYaBQdgbC9TpT9oMDqvE2kVnGYzPPQpag9qgCf3gLq
4n5gK67smXFAMkargag/3yEZ3YYCrUiAR0iCYdSog0bnga4XhQSIVyRzODVSvTT/
FPXEni7e5SQSEYDUdLj5JVdPEa53tDIGHVXKQgNeCI8HuCVvyd22xADwKCc02w3w
6J9yVqyWqHkI1M0bIlVQw/lqq/7N1RoK9X2J2L1L79kYmXp3qrCXWOjBZk9dZnaB
UahkqJExaI1/ailvJ4uOrGVPp7TNB/xW/xwHXIbRowVzpmkjeChHAsqac28Tu/0p
1H+tAkcEVeY0WbjL9Yw1ouDp9G8UR6GpxTrfr/XBwWs2DPSGtGRfe7yt49xx7OAO
k7i6BMEqQeFbOJHWc9qOmbOwsc2F+BtnnJZ9TOhKsoL+fYGvTbsbtX0D1VHFk3Ci
YBMIDizA7oqRx5w8i73vmXQ8ZBwzCv4ZE+4U3QoGRJ5c98tAqQpGXnri6aJ/790i
mV86qGiqZLPKLk9iR9MG/X22bW2B8HbxsYrV1GGe4KmnUANw3zhUUbWFZ3G4kmgK
Z4UJ5RDNzfzJkFkJrRKaVGdDG2Z76p69cBCpFfLzhpBo5kewRGR32oLZkFOROzPv
K2DJOtSbAj8uqvGcWAji4ZthEVFbXCvhVF4Bg1Ft/j9bjcyxzstXShrW0K44Q/da
e6BlY4OHns2e/AJK0hMCzo9UnRtum318PMdsdXiYhijbDyMQbVCQYudxBzMcFeGc
EaFakrcxX8Z7KDrH89NoKPwUMBPivtGkvK2IHtNDfAbJGyZoXDlldIDJ+Eqh99vn
4rcnDBRDXtlTqat0AVG4uRrw9EUDbTiGekFG3mlZg8W2edyQaMUFhh4SEyL3UPR4
B4CACKoc4/qNcUHGq/MCfMTsqwvpXf1M0KnejAxUaEsgzck6YKMEDRINEQ+pjXDb
mAaRuHqMbr+LYuhnKii86fO/bZiNokw+ZT2wHfHMjLeLtNhodwxhm6f95T4iSUnX
DnQ4YHbkTTTRhkZkiSPivnryADOBRJxtWDJN9tgi1jG2sPc1i2YnNyc5Y7VfIs7G
TsLL6MwIIpuC/uIXr4BMlv26Av7SNiqJ6PkM9gHfXW1aJiuoGoDSc8KGwkb7Fbiv
mfTLXgFBH70G1WUeE5e+fQm67Na61QS9C8wbPSySoXi5W/Zf80agLTHF38rd6fJ9
YP84v0PwVf6cKV+M+HvC3sr2NuZosDT3ThTkRfJmtPQclmelmR+cI9nOObiCSrkx
d//sgufOCDGYtlRr/RnBVAaFeChCEz/P+hIgFS/zYiwREst0z0MdSoo27ZPoR59t
E0y9TW0HpWaZem1CdWbdEQvU5oS7g/ChMw5Yx7TqxGmY1BgzyQJoon1WbKGVQbbx
O52J3oIC4cOA4BuJJQBAiS/tPtrX32aK+KcNYB3ErlLtVar6bY5LOYUw7Sq96TJY
QcuHm2NE6U6RmQvWuUkZFd1AKXPgzhUzgqdBXQTCi16bfN1ZC/j7kGL/+VBVDPm4
sJQ/Y3qVAoOuZ/rQt/NQZgEdb6WhqGQsyli0cgs7jQvkx9VgDjV/+hxhL1iByh6H
CxYhC3DSXCAVM2tgzKW1ur20xQeiBbrLy6RycfcaWDIAxi3f7h2a+1tEkOVc2U+s
GRsP+DaOenrhuUnHjJmdbdxcRvQoHxEKUGJaAgJX3msnBZlbGE6O5d34bjfnHfev
qs9p3cxk3OYmRV5H+XVdwLzSGAR4i0a4RNGwpYy5EuLYED3BE8PU3613uKEQAfvY
VMrs5WjbNXUgnL8tBJrPoKyCVuzotZXTsZD4P7IgmD8xOoMgr/a1ldeaVDS/APPh
wtqrWClMatD4hN47c1I5cMwNQ+734sgph18YqpyK8nNATJuVBwxfAL+xnr7HD1EF
1cWWSnovpKdBiyle/hEazD4xHr+7SFl7WGUMfsOEPHCOp6/EgvZWP4Ns3CEKKGi+
ZlttLDWp4fKP0TrbqzC/BPogYqZIvU4wgD9fNHiCEOBilYu9b6SD4AYObwPZ9Zah
5t6mor4lytrQtuGIzMCMYc4XdLloiPPG0AmpXv2dXL/pxVFUKgIcEH/gSD0FthqH
3e6X2e0qoTgkNkP2NGKaW3GsbSLF+9AlDWaGOk5G2OSA9SSsrVMjiAQBV4ss868X
vYQsw0SGJL/kXZw2qwdgU+8zck5QKnHkmZDj1eMAR+SVRc0tVxlfHe8ZuSY4MtGR
UX4+lS5dojaBDRO03NeTiLsbuU+WrIu2qfCwhJwBupNYdAn86BJsMOMbTRxuRPyW
DLheigXVSCKUadtvrL26iEdtrKDCm2ah5LOmxntRy3zE21eXnimvfZcNDRh//PqS
VZMNs4Fg+oLS2h+QivzI+ypZO8nN5ok7vWGEddYwCam65IqdOtyrB0uZhDrrLAS/
8Hj4F/zL3hR7SsfZRtexbPcpUMvFQ5Vwq4+JYirHHQlgU0JgT/wKQFAuzq1IFTWJ
VSAGneXA6fnzIe+SCw7Ljx3ONfSxvLHOT7BqMzPrf3B1FIADM40jQ5WmMT/2b1bq
1vi0XRkelP/6NNdLrpB7izS5md4VuYq501Z8HXM+zs87q8z3ODI4j2ZrgNMSCEM6
jiSCRPJcP3gWzKBiuyzWZqCvHGgqfK7z8EPIVm5BNfee+EjHujO7sTyFAUuEzIvp
S6dgTanSL15cOOBI+f52UU24DvN9toWYXUan9Zg5h7y9Ry6v5YhVKn7WQ1Roa3tz
saUVUzQTSrquNpr8nrSyx0EQwAW9h50Rncs2NqvwxXeTQRZoM/3707Kc1AxUN4U0
ovde7gH7SSXwj5NKo03Um1Sd7FxP0W9IJoUwwDEFlNbZxrb1kb76LpEmtW6PmOO+
UogYXV68NKykNLxqxxjpoqwCDHOIQ6cFFy0VRZCwZ6Bnmrmb613gfR0uFA814oxS
OP0RZE1n+3+lHOnlshnATSu3uwWYX0Mnj7reopV1gqoG6T9JVO7nguPIt6IopSaz
hKBlGKqjMMFnYSvgxaNEVkNycN3htzfFo51E4oiOtTMKTe9SiL1EBjL6DpAWxQ52
L5dj9OhVNay1ThfDuakWJumM56kcV1Fp94xb/SYJhS4ptq89LZ6v7zMjeCt3rvgl
+HJd92pbdi5HRUqpH0iRQHZqGbCgy+z0P+El1oYn50wCE7s+No8nXJKQIIVwwGuK
0ABfz5zvWG5sKwXdokaEcYqu79To0SyinWLc266clN1AETgSCahT6e6AXlSR20y/
3xiGp/IlYZFPvpuzV8Xs01mWr1y8SawukU8XnbiERwPfyEF9Vglh/CEryoRLekHr
UeQf0ggkVV6MJSPjxlPSCh6T7Dft8Cmd59IT2LJxjXbBopUCdIlgp0jBZnKy4alm
1SulUHnOfxD6RkUiGVeOtv7PhbtpeXrIWuAco9DGonSyNT38dwuwHZl53jeE17v5
WxkFs42KMKajePMCuc6t9dTILCmIKB8vgAM6KG4Qb91w8L9D/Su3wqJ3T2Y37GCS
DXpW+CDbzaUb/qbdTSR1Z/E7EnU8CVFWVqllkUOp445SP20k3TC22udKgjF2g5/K
Odf8tZVzjmPPDwYtqeIdIXQMpeiDKcFA2hKBsCNvPdCUN1RMs2hy9AVpBTOui2x8
Aw6vYvLdQn5q6TWIfbuihoAc/uyyI04375uu6qBN+/R3GdvTHV5Uz34g3p0lBS+h
gcLCkkgJ0lxtUJ+8gDeyloc2+2AgjorPFnO1u2XHqpQlzj76SptbY6RcuFqYDjSM
SLFoNUMF2FuI2G7hdFImsQUih0rqMXzBnKzS3hEURFGN9ujbnjt0RrVqu2WY6R92
EM1ZQnN4JxsO1DiG5pJd46DPPv4/JvVmOClSfuXUiJqxbdcXYMGQppHFfyB90ZZZ
IacPFtBAldzxQSDVvZ4HrDXB2/vDXbBsyq9JMqJTow2m/zx+I+4XLQ1A2SMFoicB
iumjX6BJq8qUgNX8jV3CJn5yAv+L1YLvYQvhj14itKcZvqyi92rIAT7Eo8eCmlgy
bZWJPuji1l/JaaPJ3Mpj6nU8hIZj4QMmNPKQYXs9D5nkAjBfV8Tbs+3lMYKGJGxd
j2MUPDd2WjQgotlayjyFghI4tQZLtycuSquIwo0gggEkqo7PGBc22m/CFVXQQHxX
oB94RrX10Tf9lqVXAbcbGdLTEjC5wCIzxP5Q46WyM6Z3De76Txb/Nhs7U9ZY/7JK
dcCSZceWdgJu2kFPnAOI3pXpfP6YlH42tJ/jZ32130Z6CM5l84l51KI6n0m6ZWsX
WH8UGHlP5yM42aeU1D4VJy+376pFoi68ENLYrCgBHg45VwhyZzocxLbxUqkrSmYu
hQWMalr2zKtAhBaRR1vALlqNqwha4mJq604Jg6bGWFYfw1M/haVVN/cfvzN9s9XH
eGiz7iEWaEtDQ5VwgPg+hE60UUNTJqCPQRV0zEJqX9FfEVLzUqmAhPT3dUuba/oc
oUHvVq60itcUv5m5piK0EYI5/ewHt5nFex6V9aG4s1hskxm39nI2r37qhb4Nf/LN
ZseKZZjUqOy+qX2TgVNAMeLq6qaK0+ZBTC/CkaqUuLXyf+Dzgcy0TcIkOB1PSmKI
/IHu9wGrMCcKVY35AkAvER+xNOOTkQpqdWIvz8FLBxZCCv9mKoR/VM8etOJOexg6
byzDed7zNDOl3PlJOdTGt0oIT66zpKubUf/guLe8TrWoijuZFvI9kaS+fFN+Dgke
cKMqpWRByR3A6IJyxH+PFBZs/X4ShvGDIT4xanB4ss0kRxOdtZghpBqCG+ybgTaT
v+Rgkl3gNb3uMeuBVOm9yX843AXgqJWc0xsrhi2jpbYRMCVxJcvJF9E+9c0Zzerg
zP7Vlj1WM/0b5gEH+6sfRvkVlAwccEo9Bw70uEKMJQOJfXAepZLMlMWQ8kQ4cJen
9vRvvnkBB+Uw7Yp/zHObfPzmDVa5wzkpDAowwc8p1cXXTUBJaN/92MKBCcAXxnsz
I3CBybdlV40mSKzGiaRwt/QxdeMTybzmfmwWiEKOKDyHP+QoetCc/Vd/p1Q/LpDi
rBear9xtEsEx4fY6ARQv/0oHapMXXHH2D2rIgQcmRBDNUAsU1eJmt5Gb19Nb2qGp
bfoczE+use+qtzsZGc9jVgeLkiuWlfeu2I3/3dSvAxGXZPU7XSxzEZpuIdi4iOG6
vev9A2Smpzm4yGRkBYy6y4SszbLOo4ZXXpa4Kbytttp5412LXWchTdSHsU08ldYj
+M/nifkazAIqQ/3ncCVeNxGFqz5SK0A3w2FFX7liVs5cEcXELTSAdP/jYT23P7AN
mS7WpkrJGwcRcaEnGCUkHUvyzgAoY5WarhMxPlxXw3RN3QJ1sk6lLnMps1QMM2bL
TWGY+lOyQY1EQKqVq3pETBz75coQvhCEfhxKOLlXILPBbv/pf0rm++oHpwlGYN6r
PtUYPLFMZkYMkdX2esfKqw8+uJtAV7eML32Vw1O9Zb6QfrUnodIcoga/+vxed2g7
KX253suGuXiBEiuT0IyOoPgZp/1V8UDMRctjev5LNRdD2l/LIMylYhSNN3e589rs
JMbfX04PJznbK6I9ax4YCXYxJu+sl18hZpU3mtJXcC/KTDXpdshyX5mQLkMWlY1j
4fdHHvcDUJ6K3v8/GW02SsV7WMaepIq35WHxFwjvnkDgHyJqvQDUSAPqIWXymqH4
nhccBXwJj8ALtF0dhmZOqz3wXWtxC3u1vFrNoDvatQUEyHwUrNt+evidfnykau6a
rpknM9qCEPYj8olek6aCg9jkVbDE2XNJqGGNpeCh/FJBO5CzfhPp4dQrNeFyrTSk
YcZuJyECXgUys4VQ/oKZ+nKwKQrwiFr3UBrgmTuTs1PjjE2NqBS6/1vaIDolmq3S
QyxC+YHVw/RPD6/NR50oT7pHIAJ8IW9FUWICN9oYj/hOOQHWPxntrHYl+Y+VfqjA
CqmNOxsAC0Rn5E8T0UY6p/S0gosp2he6zjvG3jqAF8qJmB+gcPp7+7mtrNlSaAc5
yKGy+AWSA2WQdep1hvYnsHVc7zKj808jmfPWeP9MvTtbR1yLOOJNSuKhNjjAGN5+
3p5xLh+nPN/7W43ye9ye3ocd6DgxMmkR6vVq+S2YQUFqXuFKrIj3NvtxOcqaWQwt
YTC2vfjo0+9ROZA+xM3IFECUkdMI4VUwYkvsjnRQ5aJ73huV3rmWVZD9oIzsytwb
TgToh54VXy7D9Y2DEeaeI1hEPICdH26D26qz0BKL9PVQ5uHvAPuah/3gXZBoY1r/
+8CZYJYPXTEwqe2RP1rNMsB35FDz70FmbQk7aBBpTmorMnO0PC6wS7XNT96Hy2uG
nvKabftzUPQdENzc1EKuINWNpMMmvmO0qkOJMJk0K5GN4BqeCmMU54deqVOr3RZC
aH4WuoHv3rCkPSDtKqFckQzudliUiF87Yp6Jg1kZSW/sTCQYZJwChPKzuaDD6XKq
ZQrQNV+cnnH+/HCSon5nr1RKDptzVGIDvNS+NAx4g56rPYmvjXARwg731VYd9hKg
xg649ulzpm+vwYggHIJpuiP5CBQupvaaaQRDag6uY9M9BusKMSH9c1rIgskiLydR
1ps/ZFrT1t7w9quo64+7p6YJSZ3hMowFCsqohLdu7TLVNKpXMjt8T0Ex8zW2Mf1S
wVUaGj5voGtIcNb8faHiJsh24YH/qAGliAYUIBKIOV11HA4LMdXRGgdbEw/W7HnE
Dw43Ue7GVAp12bp+ZyJZQ4eAR7GltDzQ7S1yMRpPxg+9+83Wj46rh52aLp41wnYb
iXwx2tm1ePUuymU7viXDeQGsgdYt7kmHZ1/469ESwuaimtOn+bIGVR3jYx1LJcOP
jgT/spM6k2CTQpTajk8K8mwcxPeF59rTrzI5G4KDTujC+/Yeqwm65GJ/P6lAoVaQ
RtB905lFUJ/uvjVDwPRImOevZWv2d9LOBuiL2kcDyZpmUz9Xn8WU+GYd/JoZcNIU
2v8CieIpp2/kLuJfBDk6iM+EpkiHyrj6PPNRsPtXh/itFKpa/UXH1NngzUmVqhsB
rI5DXYHA0Fzjt4Iv8/BafVU7SIVETXt402VfkSdqSErobobkAeXWgpg+3IK6nRWg
Cp8OpSbpyaqqM7Td7Iadus4hTdjsEcOkGZj0BamxHg1MWERIZbdmfHB3nv9lE21S
DZVZQanOTWF/zwRyVRlgnKSWssIrmivtVglSH3zlnj8+lLy8ch45W+iVTow59TBm
30U3GMN+xd87Iw9FUV7htp1FJJXu3hEQVSJhwQWmpGZoD7Df8eLCPYmj8xsxFMql
+fLxAI/6wtqD1oTJfyn++Z2gkK2jpv2iHbeSWwfTqBdkNhtrG6D4Xy+prSr7xmHZ
GZCd2j3VXEpfhpqcnLn/Bg/z5A3aEAvKy4fErQhXpxh1veBWkrMSL8pbQ+SY687R
TAP5pGuOX5XRee9S3F3OHTRcxo4Th6H33kWsk52NMcJORMKIeRqI8A96Zh9cs5xX
R42cR+kdHPCzKQq3KNmyHFG32UqWPcouu2EGIMCchYBKpO1vZL5aMBfbiAShHwM3
8WGf51gsDK0oluQ2wIMAyiFFdqGS5ciS3PMRJMyr2e0PV4fjq/2KPLQI3uWU+qfF
JYzvoNXARmeVdft0BUW7HUMiy02dhQEkwBg5dIcE7fHxpGLALricgYFEwxKbXodQ
gTDGc/AIy8reS/iD0y3CokFrra0Xv4lfn30//4N4zx6mOVt6JQ4eyXQZjL5l0a95
k1YeVkmngRblqGqI+gFtrhgEI+ieeA/wjiQoPZWCL7d0VDFQIbUqgj+APPnySXRT
uApn0hfDjz2WOEdHe3hsyXR67/DmdR9A0tNgP/9cBx2trC6OqIW3rgPS9qRc0yqA
spxMXWrZja3eR5k0NbKtQjH4nlkIdDbLiQUvlVFZzcO2h8GpiKTKqPmk3ZQePZXo
NVu6t+HxaOgb2fKd23/MRdv2F4G5KOHxsmFdPr0p8K49LSAt88vsSzMVa1eITuqZ
pktMCT+wQJqeggt7tBvRrslfdOHlpDgA1j7cSl19NBYNKUpKtJhb4vUqzQP9xf/u
Z8YY7xy6nPCVD0lqRZrm4FeQVGcbHCZkPKwmC3d0d+a1RYVjwUoltsGkX17zRvKr
pPNdwQu4dAGt4ni4z1Psx/b4ttXXzTun3J3LZ81LwfpwUyBAJ6Col8sB1REDiRM/
re+KIIyNZTGkYTz1N02xB9TMblME5KwwW7Dq3B++tnykzTUI7YIT/YJkouZiOzQu
gZ0GzYgFrrgwxE0dTJ8lDnTEZe10OJXt++YvufUQBndqXAn2/w8zA9hwvChLVkC1
jYJdGBFc27Kh7zqHS0QPmbq6JtRlHrGnxg/C83GnZ245BUXYhXkI36KcUfdFzE5h
Ia2x3N6EYmX492sn5s4i+1ULEwsJUS1XHSXW2FwuEI7qi0VgeKLO+9MGnH9aLIEj
JlCVSDfBPJnaDjffWhbLnjz02wRfjexxH/tx7kC6yqkJVkScqIzaouCgQWFSrLDr
Lcyv/wb+DKsmt7lmCfNGCtseRcOyFxe1xE3rL7/GjbmSwbb/c+xOENxzZ8PjIU4k
M4QLglxcHTi5Sg0gMiTbB8sjst+X1celJJZDM124Oxmmsve9ogFzingqb2PTAgDa
cQwzfceHESUuvhVR77Z73c2Xs+fVMg1OasFfl2eyTxkEVxFdTGqqmEORkAVfU1UT
bhEGvo8YOS36fxAQqaTHoIaVvS10MZ2KZNLZqNaOOf0L0K5flRXMll7OTZGlpd7z
VBF0A1irzEWTc//TPWaD6F8kKMF/tY35e5foOqtNj8bGnObU6gauhQu0rTPlPqsI
Rrqt94dwuJtwctydupxFCspOa646+tKycpYkIqT12KdTQNUzLlUzY5jW1CwaA5VC
AGcZ2cK63pcHyddjEA3M87lc6wlnYi4BZ0rESdhXChVopjy+RdRbNfzuH6Jp4OkY
xMGGaminfV1nBxrf/SbJX99QRAUYnrlV1R9ojQy1Zxyu+rekpp8vrCZKE5GZS6du
5zEgEYs28i8OxSkzhr8Re3xyq9Y7M/i1lXIlQDqRtgpQZS+UY6sonjSAm5rjTepW
8bSDFvGWOEi1u0vbqTt/hBv4lSAYjzblYXapmcP2wPItGgYztgSNgu4KyHPQKvml
iM7fmGVc+Bv+Crj6T/oTgGO12wwAeL+OgvSF8MNjbhM8cpDdWj3v+KKa27pau5nV
kJRCimU/Q+DiF/IxJWwrss9swO9e/K8Jd6ZMpYZG6Oa8MGqk/KBxSxJGoWT2+iYX
MWWo65RLeyPP0JKAl8OZ0gcDNc9HAnyypoQh/NM4nyMmdyaxMMipLEPqSb+xrP4v
Rz/UINOk5p+LycikP4bmwfsfkiOQAAWLe4kKn7xZ46kNBd3rJmVSN5iCx6L38FXR
TMgsBKWDQRW0eSNKFxSPRVl6dZn1jVIFWhH4QyhWy45VsT3d55q5nTd0vQD26xZx
Bjv3k/PdgGl08YXHs255eB9NGu4YnTTgRGA90EIHR7UKhnnPBMxk7wmTodfJ++hJ
BaeoHc7ReBYE8kTqIXyqZwMx3wGv9MTWiIJc/HjLxpXv+skqsTvkm1QbN2Iw1dBL
wKsmlnlS2EnruzjsVXFOUEYvM/sqtLHAF0nsdsC2swbllhYGtUt/Hkp+UaMX2Ug8
9SKslZBiwNGlWw5eYWshWr5O9GxVzlFjkoD49Zv8KNTOZFD2SsB9PHub6yp2AZed
KQf+yt8Ir2hthgzoso2gdElmJMerh1yUig13xbwu9YKd9oPJWbEgNOMhPRdynrei
o5nqLHzXIW9IAXRGIp4HbHHJFirhLLTM6Rd5IMEbtx4KVr3QqGo1mvi7x41r4ZMd
CQhhMJwnK2NxG7e9PsatX3t/XbDuBDabgRRznY8uQt5U6BNHzjCesLoaiq4pFRBd
oRL83O5NBzTsCpoNkFnHRgQ1OuvYe9peHXI2c/17reHgvL8MlPtOtJ8PpCzG3+pq
im/KqKMIzPJ1un86OQ8YqESjb2vsrpYkdVs0NJE3kb4Ijl+n0TJse5FJF8gYkiIP
O4Tu9591CF/MloyZlR1DMePl5cSbBjmRiRtIFqgIfrZVgwIaBexjM+0RH8X8raps
K7thwhoowDMa9T0J1FME+dvfjc0fjrEbrQ7geOzOdxdH3zf1RkKrYdFix+hnbgVp
dqWE/gh2NBHYRnXaasclwx43fWeZ+jngWjrbpbDzf8bWzGJwkaAGBK5Gdr2ttVrb
wjIR7erN00Iq9pvPHsPwCw9Zc/cJCc2X64keFkeec/dykY8ffuHuebWrLKQNmbp7
NnIAEADdWt9NBLvEPR7fQUsXwlJmtdZVre1omk9oUTMaaQv7dLVTQcYn3XixyNjL
i6oq7eGCld2p0FYkVfJiZejFa0vHLy5b2mBJcvzx01f71cmwDFXESy3JEshxhsZ+
WSiH/BT5lEElVYd9mctTBANYmTeKgfhUk1Kv0M6rCYVuAOWKcPxiQjhQqnie7Osr
NE8LISpvSMt3uipLnZ9/IOhX5c/aruNKq3sb61j3RkHVWNkf2cnrIpF6J8iOUJUe
mSj4gatYm0r2NT3hWWkP4x5fh4oH2igT/b+w3zkR/mVZvDrYoAfwCJEytAH5Xu84
uEsydv3wT4ftKFHT4/UcVg8z02Z7b2pCYpANAGrb+Usy1jkK49nLS7WppUfYyBEL
YIN5wc0nMMVL/xpe2Kpko8yPOGX4itsK24YISFNrOj8C1nl51XTg62PoPDZNoxfc
3K7AdVxBi11P+2DgiMZ7lcp4WazadIRElov0NkFD4lA8qBWJs+fxafZzmibx7mbn
pmRyyfv9hTbv8YMuWmMB/02zC8nYMYZVlf5cQ6o92V2werweT1q6ZrNwirjBlytD
XsHOy+OkqPpZNP3Ys+m0rzD2LGFAV56b953YlCL9y1VAvw6puF+WnHhOUrnGfaCd
9UP6rvtwoeVRo0+Q1ZYQ1RUB51bniTaFyJqSK/U7bHXm1u9zVMptsBouROYOUp67
Y7FDlaau2Yjh7dG1qG7Hw8yPbJiRUz9GXHLcdnaj9emXXFNdPiX5PqKCkSpV4xDi
gaOq+l815HOJ7l369FAu4RMVj0K5yzRETyjG/Uql2rVyDGraSjshb2pKmwK1VHnA
T7lHvg15r5iKrlw5old+DdxKJN6bjfSm9quf7iZO2pSDh/7uQRTU9cn7VTzCAbII
17Kh2brn61TxQwGIs0xGzDhnI9eCVVToJWDhDj8FTg6q16KbmP6ErclRk1HO4GXY
ysyOm0mqc/8b/CTtAbph3JcPqS9TWWm75OKavcXxraytYxu+O4OFnkvGG7xw7d25
I3mDj92MmDSiQJaiTOmVCjLZIiugp0WuhM6xx5T5T+F2EQq7V+QgXXUwJ5G5a/kr
ccU4jjSha5YEzcKuBLBF8/1aeeZe1gZF+ZFJbJ49SW9B200Y3cCZazHUwTsISqRL
bHIifLEAWNVV2LrYJkhKaNiDnbjRs1ILtuMimXVGp6FCojssBBAT3WN5btnx3al5
V2aMiR9ti0rB/BQ+CxOxADLwpUp2tT27DfR+jJuB5yox8Un9kYNhAjhE+OZNM0Hk
dCpzKsDkkkVzN3eI7YA6+M73IFzoUCBdY2aRNJEs48rGvuY6BXdHxwLDxK5nV8BX
RioRhV6RUIshjRTJV5bFMvM1m/bSlFGLgQqXQvR7vIQeqKcfvQnJGoriIFLoQSAm
MM9LaF4FaPtS9U/MoOvqPprS+PubpLbUgR6keeEQVdNd7SKkXvPNuwIlZeGIL+vU
fR5flJHElOFCcRzTLOIguU/Dwn8I/6f1V7XX8JkqqkzhzzwEcccJiQQhDwR6v7Mr
5t+2vflJ35R0y30KPaa7ngMBSpuMAvltbk+1Ia2KzDCXjD2TNZ9nYM2CMBZAVD2x
mpOyQ6fVat6I6u2PxteWO70ICeOfY00oV59YLWVb1+ZvuclcREKyWyFlsKPeIvAg
VxOf5ovNiPW0j3DZDQO1Xg3tZc0uWN4I3vhWK2D6nZaO6RcIWTcWJuB3EMlILIet
QceEcZnwVst9z2vBYIA/DHsa21YbnrCKchb1c+e6+Fja3a/n/WkBT9rXMTQnQrm3
NhMFcVQ5SGausU7UloKrpl01svrXF2FwrpTYt4+lfPDEslJcOT+i0zW/59VQe1d0
YrLFskMccbkGndHedKqJow7Z5a9y7kkkx4SG0ny4rUi54zdAJRwfAWzT2URQzY/8
T3+7tSVX6Fun2TfwAwWy+sDVnIGVtS9Z6NgcMwCFQ/awY8fVx8zVIURm+DziaP1M
hiZum9e64RsiZXt3bl8VRGqyEXkaYPSNCWcxUbi8LWhsTq/eBrQOxPunqxtLZ10k
dsz0eMOCBQRUpD1iB2r1/MwVMsjNEC98vv5nr/e7yALyKno/eE8AEaYQDBslpUI/
nNMWD/eIGeDY0CITPosR2lXyZGPY39823YA20X4W7mZjqWFEoDUgXMokN9f46KDk
LVZywco1LIklG4FWFPV0/CjmYrwPEVs1XfPVkjUzygP9pmrS8Ft5Yos3QQO1FI4H
5DP1m6k7wVW9FFXJ5FOsxIcnXfr2tEz2CqWl9IIzB2jMbIspJuRNbye3WgNneNNk
KfZEly/i+2UHA29YKfv+xKH9CVQhUvt2K5r4BpqKi5jGH3FUI7fZyqh4ADAPZS8S
A7b4AMryD54s02/JopaXDjFeD7S6IF2DkpXEkzv9NZgBVHZQwxaT1lDHzbWbODvB
GLwaOXsfeglZn4oaat92NuzASYBtlAvtHzxE99E4SWYTHSWI+8NVy0YtPUaFF/4/
rQIAKfmxBiRmBdN1t47iYVaDnCZgeUXlBLTJD+bBlWpOMqoIWS4gUogW8nnLM3fU
9pLVolA6PkqYoiojVZSNOuWpUQ0r+kgaIoqPCIAfr5XL55LOzdi1qUTL3mxf9Fys
j3oeqO+hnMOjKFy0Y4xBfMqb4cza7feIKwZBpwO9Yo+rGXNEpR6mnJFMIwnuUxAr
N0ybMQQjpRTZE4LjJh/JFN7X10jz3zHVYL/mdeVyUtbpNfvbJ6lD/s2Ha/wUw3hW
XNQwjADKDLD2a6JQWv/dZspUkBn2trnGhlrUNIQZd/FubL5Y853byZ9VD/rMUwyf
M0Fr0D54RmTXrXUxmT/bp21/FpJHpIwKEyDSEck+HMfigY5uUUU4Rv71HgjlhX19
p8Wmg+ciwrt65EnF0Kp+O/K9o6ca35T5eQjxZ6Iw9hVRNqj1cqhGUovP4cSZnWCH
WM4Dh+YOVTq7G7pMbJREbwr6Wt1qAJleiFCVUNcrMS3MXbuaU4CsUtgQPwGfNLdq
fjGQnzW5Ra90/TXaqh5QTmL/3oBbaZa0kcq00hkjpePzU0u+4sqZk37fRAgrWJrG
tHxq6cxLvW7Ox4e9tY8zWr0ZP6GoUjAg24DMct7UHDRKSoyN+CWt6Md8VdoAoQoI
eiF5zv2LZ08cM5WtDhm1H9t+K0FQm7u8sOdBRBJspHxEqm7A/Vic47ggvVTbAhih
J+sgl9DFPgcfEDcK87uwLpxqav2m/0HcDZssqFaR6Zy51dNSIbJqSD7U3fC6lcZB
f66nusWYKB2Dx34tsFKDpraTeq7MYOelJdJTqfrdL5S17bH2y+lkpkLqmUt6McBn
q+hCPbssDT+eYlk9GU/8wMEtr92yeNQ2DsPwAvBouxMvBs8eUii1WPksl8jWpyKr
pQzQ70Y0yGrnAo57FMAyQ5JJzolWRdvi7nWc/AmxvcII+kJYLBJ7r9LaKKT3fCTi
hRaZvNzAw0w+hMeyC97J0RaFUz9juRN1APxWK/0ksw+eliZ+d2J0X9HcCNF+J86D
o0a6Xs62Zvy0NKS8ULVeCM+vqybyx1bLK3PHJK1dSnLXgMfcyng6LSBf0VgUcW8o
8VxDNbXpWWsDnoqbPE0jg6hU5zHfijuCxWCdAzR26otaTvXAb5NKaBj230Sz/Wg0
QtSgkZNDaOX++dabZ7YRkXVHJBLQOv67Is6fF8BLgw/aFckINyus53/mcEy7+vpq
RhfB4zB8mravxt0/O3ydVsRMszb4LcunZoF5Vm0Jptq/tvbZXQuS5FRgDUKl+xXL
28EFvb8EHg9jxPHEZvUIDHKg/djyjpCuT79C+uJkzAASH02W+ySTYGTKFB1Tbx7P
kpd+fanSfCYfzBc4YY00hbXAhBEBZk/rPWsl0BHumKRSj1PZCWUZr5RLnv4tsewd
/S/IXvWk6JHWzrXDiO+pU5PA0pq3vSzeCNFFUh+hJ08sPReQ9j/TTn0EpHDd1RAq
oUGstXmyW9Pp6UEcLq7Fjlb8zlw23l1A35kaB1lWIe1hJc57HvfpEKbNsCe5DsUx
w5Uy2yI2xTixJ3bz9HwhV39H9/UhS01Ex2zHLxYWexqucZYgroU9Ar1cf9yyfrko
D3iZmCLlmiIh9bNti8vxrs4ZGMz95S0ZNkPXjpe3ZMAsjIx6Ho0ZaTBtQIBaUjrW
7TuvT7kenNUw88uRIgGrVSlJV9aA6ddfVBdwhMS+CgkEqwOJxPuVmSf0OjUlE2Ml
heeXmePzQ0X3YljU0In17nqILSMshCeQavsOOqiZDc86yTitLjzCPiElRmHX7Qu5
YMnwEzDntmAv9aPTBotyT2O1vqy2B7RemrOQH83LNdE49d7ctmneMCBJfHkW30w2
V19KstFoL+xo5gzJtO64aZm80mXEB0VEgSQYmgor2yoWN1DpVEBP0jzU390YSJnb
QZqaxQULpPDtLLpnv5nq/nNpVkTktcEI93f3Vgrc5vZsNkTTz+chwEuvqZ/cf7/u
qH6I8Lwj/ZcVE7APYxBU0DmIi1IDLat3zioA6ARuDeP1xuFaOaF+VO71G5XjSxtR
jMcpRU6uAamzaPzSR47vJ//Arz1WQfjDv2NPKVoxRgNrj/Xo/oNa8iiXVAWLTx9s
kJPTbZFV2D+x5fT37FeyNEq43kO3jGcWfOSc+Fm1FQ4/ClZpxdkHXJ33SEhA1PWX
oCXDksfGayUu3GWL+LLe5jLuU6/nXQ8b3JwzK/W306Sf7gkAPU92ukWzCHpe3cI5
0XDkzOgkMigowK1HR3MnGqzBM2RcD/mNJrb/2Kss+AFBe8S2k4wtFPJD45FbmAv7
4iJG85q0cU69Yg+jZ8408CjutBBNe1KOWUWUruoc/4luyTBVjs+Wr7zUDjXOycPB
tjqv1BsAWyhMOgqIPat0FLzLfwZifSvtKnrUZxjOT3r6DDwTiwQmS0WaiFlx2u18
fRWas+CF/pUlUHjLYlYHBQ3A+G1MWapZzBHM7zopN9vP83Rv7ZZxExIiVpKNAHOA
ssCXxx4nccaneEkyn9DrPYzSI9LhLKOkvY1XRVb7tm6diqKN7VafQjwesBOvTHa+
aatPWnISgouq3btXsnCLXl/Vs7BC9scyictqttpI6IeRNKmHL7pnY3gMiFkFko8G
X6WS9v9ORwKIJs9JFIlvOrpglKDW4rq7REhC7bLx+UfCoLUb8EVV0xiKXwMw+x6p
HJcmmS2J26MrvB+h+T6ijCUbrs6bysD8CPGN8e9FMT3VU2Mur0TMEvSzKYI4Q+Nm
n3TiRKTw/T5oNDzThj79K4TLL4+TH7CqhJp9r4h7c5UJi7W1U6u3/ID02Zee0Hpe
Il+joC3uVhGr5sD1W6Z17bvpyyZiNrevWXBfm16WnkfGv1JoD19M7b0FyCTuE9dz
lt8Cisg5T0RdaCLD3RAU4IL/IKZD4y5+D0aZdJHAidj+qqjM7Sbk9s6SN/hUQwwm
N8/LYbdRb7oHUli323BT8/ZvR+hGUkaaX1o8iEloRyWUNlJ/C9siP9EZvbFdHxe/
sVeN1qEgzUaYwazH5wt6v6Rlqv7G5lsOBwvqUx0F/DE2hvAbKEj9WHn+7cb8jNob
Sp0r5c6+xbfBsHW9z7d+cl/BpbcWQKGYAZNGA/vjo2RmAKZ9D2y5zPzzXAuXX93P
ssTqLAwuAuylyPc+bNJThkHOQORhxMIbhQTQHj9TVHN7m3P7ADS5/RkghGJ9k2n7
GY8OVfFuWBfuDDFFewEWybwaW+yEMdy91LbE51fHsFcwwZsFGs23MAm+miJiAkEB
F2SXHY1xw4ifC4DB3yZcZ2lI8a0ZTRwiq5MqNZDr40TIyV9JwgDmWaTJ1cY4mRMS
3w7Tgp9YA9RjkvbyZbDqTeKjiWzRUU1Bex6350A997jXRIE+ZWDn2tjQe23Rbd3x
Qado+navdhNK7GRgFztMuvkHfmLLCNu9R06taC9G+JtZ7PjLxPsoaSlErzy0zg0R
b4ktCVcYiDE0fMOCjGEAYzqV3mj+/IgNWB4KLOkj1yDnIdTELjJZG323BGbDWmts
7wJ297yLa6SUilR+d9sMknl8UJA3ouB/XitfRn+2oxtQs69yH3YzJ+vCJHv573Rf
RBnh4kvkDofCzwtQvtwGd0aBZ5yJRDSGFhjXliDXFHDJDi/lVU0MHidhg6DEBL6D
pQ03jepajDuC6K+A34piG477m7UdFUdQOC+g6XSmX3D6T7+YnM4vZGacKr284lvx
LH3j/TKRZx7oVNw3RSKl9fcqchK2o/7LvNxE0c8r5jUtksGq5IuhuBqySZ9tSjD9
qGzwkHapxiqXCAEdsoDqmU+tKYAfhnMPl5l6S7tlTU433V21mm+VPsk/WkCdP8RF
h0d3rkPCarXUz7cT/9Jert77HizFWjXXu3CQLdExLthAWW5SFnaba8Rkfk2yf72E
AdQ1GaEpsVyogd7X8zLKpd06P0nxDAW3pjThobKcmFMuEpjlHd3zMSsCMBJYCMW2
czvw12OG3iFr3FvPVCRavy9EuSPzVm43f35mIYF7sVkbsYav7/HfR44YnmAjVNiI
GirdSX+gbMHxmfGIFE8lN0DjumCpy7PifJ+t2uIeREE5zEcibtpL1tP8FzA4CEk/
TnSI7gAgGh1AKhvJo5i77nZsfuUOaF+HSnjSseD2UbptOhDXfFb2XIFFc6BXqQbS
Rd6W33QkbWks8TqpwQ/8jBT1b9yx9dWqNqGWqoCRmUgwXLuk4XIepLOQ9l0GApDG
Rq7b50WJOoztKupiIDp+UaRBRaUxQnTXy64uxGsZXweYzFRaHoIpOUYWlLfStUz5
WghzvLACWYjmvQ8Xvqy5cmbruOg9MnzG6Vc4kTerNgoyF/NGtLqa0aaCRIS/Bisg
D9xYHcYeGVUlpz5/iCkyIRmpHbkjzLiZbQstvL2hLBbKQTSrYbgUgvb2D/emAm9t
zNuKlkul6JNj2n1nUUTeZsy7Pb/6siMJEeIdfT6BZyYDiUvuLnDifhKyq76QsI03
cOXnTrV1UwKF6R1o68IPxhp1rAyRbQilq/cbr3E6xy9QHKV4KClODl7S9LMYNrvJ
QjgVvyZ1W7oAnqSz/cSBPpf6jR3wnBLigENtQnfOtlZCcsKTRK27qPa0ViYtPl3Q
kWENTpfFPy84CNlQseUHtRKSQUOsJ7g6Lc4TYDMdHQlJZfHstU8RF8A9SvRzyx7G
RrBFf5EtzF7UHWMCR8nQFm2g0VOxwk9iiFmip765zh+g5sWsYh8RcDYEVAc0eTo0
M7zRxsz9rW6WCJ7ukhEkvQyqXnWyu1NWz0iMbsd9If2qBfp/liieXBnHBB2xCDxv
QnKhipviLas3wRw9PvDI2TRQOMOKcHjLtjE8//td0fdv+PERf1TvOJDYGgbUAhIs
4sU8JRCoOiPeMlkm8MMz/wbtVQBUNY6mDuO2nvsf1dHYYSivMBSbK6iGltD0ah4T
73827jzwiPRcVNu0DceSRPmgXXsAHFqfu9guvy01mekzBmFA0n/9fUcYLeKZnkQG
e9QfFFah6KGOMlQc2VtI0XHKHnaQaLCzZyF2vCkYRKCIWHZepZlBB8QKExHQY/cV
VtGPt+z1DqkhQVDxdFg+KCyEPWBpbzUUGwrUFYrQVwGgDVwkoFtJDXT+s2oHOhwN
Yo8b/bTppJsBNgCY4i3Nq3NrDjOPeJd0BLDt2vr6W00LwYbdceeCQx1diBeM4rwz
jKwG3F8+kMnhT9YTNjemAEGgqOf0Ma96g5K58OcRRmTj/hfDDTZ9wg5Jq9+MqaWQ
5Fwu/IfLR+0X6Qmh4DTKNFx2vaGpGQYloAT+UQQyJ4HSuyObtJzyfODiaA+ppJK6
bdAJJcgWWHcPUn0+4mkkcWuL+va6XjzIGxUxgLoi99UtK6K/glj6ydABKtYBr3CN
QgXN8XeHNo4Oiil+swmFZ3JWASpxA3zerTDRRGYSU/N+5xvsn5znvEpSTakbyxsk
2njuuKAMWkTLzB98KN9TqoQaOwDPVy1ctDbz+8+d2E/uQdI3rWnW1w88wRUhdgiv
7rO/BnqvGWNBIg042iekjcsai+ZUszlZnXXa8EUCaXvhN2bmIALHlqBSJE1MLlll
8SeV+ANMc3ey4o9NIvAEpVTo/Hivj6U7Y/W3a1S9EyFxdQiASKCNIbOg9jUpVR01
T4ORVm70ciXYyXlK6ksOebAZEOn0kK6NUlyj3kMrdRlYyK+Iy+gdVq4MU1Ciyrtx
x522IVjs83Kse3+J0TFTd6rQRDQiOEhCSaBHDpbzXzMABHA9nQL/o9O3JHpiFm26
D6jqk3cQIfK5Zf1ustFE1kGuV1yWa0cryv0brxUA1sQrWkj5WIJzcWWZas+o2302
u9QZ8NhnkL7L/qL5dnv/bGSjOTIPEAQN59ENSBYSV2uyg7A7UpuD/41qqZ/dWlLv
utxnhZUNa02ZSwHm/4DoZ1QOn8/RuXBTP6dlv9xj2YpRYd+x7Ee2XVH+9s+S0TOR
ue2ANO/FPqAbTIujknt1jP1HI1NsOuqAU84xoP58+Mgn1z9oACZ8njfQ1HorA/YO
dEXz3c4B+Ipv/01JIEQVJ6LJcdlyMH2TwJB/hBD1UPA6cotx2Yfsk83ecOd71WQy
afUTB4kaeJOLXN61bYjHaSVawkWkDEBJxIhIOHkXbZU5zpvHBY+8rKCVu5nWxsGT
1TH2fnRnBSCYHlmCwifNNQRblZDycWcXI9ldCv7dwLxsoUhjc2HzHu/SAKWm9h2D
75yk4PpQSLQWvvEuxqMvu06JSXUB7ZxATS31ZPmkzfddYsnjBTCdj+koFB85yMrd
/fwjgXDsQZF6oJ4K3eo/alnrcFkXL4S22c3w8tGBZ29Ed31GkdeREntqwbgsem/v
2ZddNPkcNFzdwDOTOyi2urnXOWl7Zcv9s3W8Wh4ydrJLMQMCqFyhwfG3JmnsAVWC
oCEC4u4BW5EWCn5mhU5/ekIFO+8ssMmXzccihSwvvldzEr+uKRAsMzKXiwSboC3u
UyTnDSO7Arj5W6nvXUyD6lM97as3LLndlIvgr4yoqGe/IF0jzttM45mntoC4pRIZ
//QvAe/H/G30bMU9jCajTrnzWh6rES0uiJWdEmXZo0dx9Zo1WRy2wxwy1XOSfxPp
GtjomKSxWTJEZzBo+rygNS3oya9NP1mAupFQw9I729dSJPSNXlYxyw+9yeS/7GaI
E+AWZuDVjkp65p6mbdgUYe2O+bxlpgbuRBVLY7kTXKlm+QH97zh9S5qzePE6eSHu
pl16e80IxD11DFcC0UO9Q3jqOblKAkFY5VhPthPg7ejfqhN8GtaH+31lRbDM1yyN
qCxhehQZPNDEVP9Zx+evzRNuzQvK+t5VirCwIIeioywZ7A3nMSWnpP/kdUy0Onb3
LM24q9T4W+D5uglJ6JBi4t9phNH0mGmrsXQxn/P0U3YjDMx7wQ/Ip18IgypL7ekJ
NPGllMP4kZKziN5kaVtbfhv7HHjkZos1sU4wwO+zL+Sz2JtcwXLyB40sHY/8wtUy
hJ8p1ROzZuAWWdHsZI/ywe9aTvmkefwdv7gLZCfNYUsISG8ysn5+rwo2EzlnK8FV
EQV+udJrKHS65J6A2sSJbQ2Z1qTVdVxytD5JXWo9njRN43TT7Sb4clGJDKfUewMT
DBXN4XdjEBrkIz738uQ3Lpg6MqTU/0dCH7ZFaWN03C2n4uv+nHfAIheNcBp0PZPk
uGt1MatYRSGe+mEKIqYxnQEGyYy+LUKGk7HU1ZY3DPrHIy3tBmMYOagcT489SZyW
ARSsO2Ig4K7bqLXunDhFbOLMx6j/p69Sq1QyfKHM8Gk0ueWYBVExjrlbSS8B99Mk
shy5m74WnDVsJHhBvFkP3KGRgS5eNTREY7Bp1dA9TL5O1KJhNiFIPqsifh9KZ4kg
3sPD3QOcdrwzkbsl/5f+qRQqeJwBZ16WjhPJso8rV8gXtfOry9D9PiSxd8kisbOD
vl4u1jxLfUtPiHAw7mrSpWBJ2WzTXtsNhzGulla5w3TifcpmnJ0ZvbqdC76TAmKQ
EZhLraqieq30cZP6lL9gj5tJ4VBptQkQ45fRDecWjbybhncKlBXT1/Lkckq4w8t9
xnVcISCiGZL86YbTMtZ/pFbcvHtkdRMl+O92KUHZtbu0GX1vpOn7OI2fuA9v4mWQ
y0YPY6dpJVxF7+z93DxifraZMqISV6AZuR6qG4tFNaAeXh7b/iqhLdGtI3jX9PNF
0GIyZiljTGIp78kIpBGXHT3OZ6bI6QDFzHep9RXZvkP1V7kQX0MGmpJnkWen7nrG
BMD0HHz8W5+q1aTPzS5sdnbj1aEqTxA2qvWc9rw9ak0pgAvGR2Azw/+R349/iUIF
72R+BfxNfpo+KIEPoZb99s1EtuiseU42zczma8Kb9b7dlSs1nCrSTh3nk1uS6tiK
SdUw26p5onvZwl//vSKrpR4VXrVqRutMH8Zl/7R1GkpEenuCF5dCKgpXHj3Iz2Sr
k4Dm77QkKc++WZJGLHDRZsAB7Eqk29/rVVTE6y4Y3oG6ckAGteWZ3SwS4PqhI/AD
+Ci/HFCj/+qzXFIbfVtztClV0bN6T7m8dGsUAE//dNjNnuZzkHmX/2yOYXTor2UR
gYTyj/amBu0NXgNbHEK2j6V7htW1LIFIcis2Nq9Hy9c+x4c3y7yjThK2ahxAG1J/
VSiZCtt3k3FCG3Bg5WpwZHXOCMfShmg6WFT95E2TLQMc3cC3OiZMpZkeZKNXhif8
Z/mtpsSbgfZ8WUneogpL2qVMYqSQemglGNay0G6RGzkDycgp1knG3RZ2Cc0AJE0K
8o2F25LCe6Vtq8Sz3SEuOXrrpO7F94ZgKZBS+h3QTgBivgFDagaqgnZfwMHbYOmX
lSTI6ZaL+YpJ9WeI6CV70zWkLcVK9AF9wmnvYj4Fhy+rkES4oM60FzU2R8Lb2OAH
wqrxyfngX5zcaCMuRuR9WUSV0CY6Ol3DaLs3vYd55kgqqkoa9bAn8gO9Dn6PN67E
B+cX96OnhGeAIDquPDnqptQ/e0alNKGlQnudZCcSVSeA9jv8yWovKTQfpoCT/SEO
Ltku2mBmTTUpHyAvR5JxyoZJrvtx/5HEdHj5W2S6J9ieSU8ZFeoJSVow/0E0y4GU
8ur5h28WnR3aK22mMTDUQ9xiVL3kHD/aACtDGBSacrjS8gr0mLMKnG/QcZxevNnt
fWINtI2/JUywxTtV+vj9/1GQzk/6ZkgrogdL4OEIaRDZgfQQw008c0xBKGNB6a3A
N9u3J1wi6pPRQ4insssF9LaUtqCmCSJ8apF6Yvg9/kIB2Oeaxd0NoaJRN/PX+kww
QGBPfhRh+KOw5c6le72mcAH1OWHKoigmDk5uvgzUO2d0XK2kJiAvRmoVKUgxOY/I
ciEYg1J0j8A296lMkWK5OraOLJ7Wcfs4njl9a4sC6CZfnZ6m96NKVJXkQE6tNGcO
VKBLGw3zzNErg95FQfwk9RYdnt+br+iB7d7yR2sjOYFWmo22YvW2Q9NjFiCso0O1
FdOTJgSgJkDcuUHnxQBYIV8CzGIEvWl+Z8F6hxvI3XJVaxX42X5KjK/CozxOHUpV
FeO6phG2bNU4VmhnJ20x8Bro90SQnF2noHOF/i/RhJbWp9eeTX5pgxuTZE0tOZCn
NoTWopp2/qEZ3RB9kQDv4qycolw8cuLVfhWRmAmfReQg5tCSg1KO3FjLhoWsITJI
z2blwd+21/mjScd4i/pk6RpwKTrOEVwNMbNroj2KgiyXJEzPOkbPQMKGK6gEGb77
nOwbhFoxF470BEFJ1mo4ARWkxMcYHLMDQk2RZ/kwI9LrfgZ/w+sRN9EWkIOgxpSY
L2ghSFijjHM++dhcvirq0+HNZxXi2+vlNNAHR4eCe7W3VYyPn1sjsg7RZ/mVk6YF
+fJ86COUbwvzy1RFVuh6tuBqlCs9/htL349F1Yfs2Pe6DdVWAmyncZvHFOO9OIlk
EH/MP91SWn2UW3omrrrHzmGiPWoXL7bMNq6ReT+7MyYOWPkvqWCP8sGDgnBf/2F/
MyDFa44fRrmZ84acMijuL5lUqnj8iK/x2hQ6ykP2UxPUCHjBrqKhY4HvfKOkP5sz
p+BkcfnJdaQXEQ5k+JSb7c74snH1iLPZL8nycAj+2WDHGLUVHdOnFZKBf77L46XB
4Nj2GSHNa+HSVrTtzghISyq53NZEhDri9KJEhZYwRBSzLzuhtxx4Eyav/fkcW5A5
4d07E0iePUlLz5FON+nSfyO4bSoRNmZYWEQmrH3NK45Undm7bFxycTw07za7OE4u
ssJKddXHRtenKUhchSk2m09jWjzg9pd9sKgQv+37OYt+Mg4Erx9RhGgoSeHa0RIk
XokTjOHnTpE/aFPqt0CqeLMlllspuNn/47yb4KopnMJc7QA9iyx4h5qXvS6004jN
PPgYvFpsDANQISY7QNZT9VXssfuvuo5RlKtPeg31dcfZB9vPymhtj2AO9oaR6DVK
GU0PSzfrlivez22wToqaeQu1YxUIvAN90AWyLmzdUWFU37V91UqORGWSgRhQdM6X
LZ85V//JWkOVAzdoifRDtDNPCbrTjtjCuAY+bekgwyL27Ud+VD3sKEzMvBReJIeB
IPtnGN5OqL2vDdHRjBi43Sr3YwFBIrNq7FtGaODedGDMbgxqXnqXebDSGFsc0t+1
HdGF7+LE38DRGpLWLX9qs2hZ/5+SiwAI931m5dePD8+0dkbtznGzDUg4O2MZnuYd
CxXt4EM8JysomG4pV9QqEU2lJy8kcTX9AqgVn3dRJ33xCfXGSjmXINaWA/sccudd
gDhu0294MlG8cGguHZVeQNWRtS236HNL+D/DXo9WNgrQ4IaDqw14zS7DDfNnFRc/
iWNNU8AQJhyFGRNNXSSR6fpBNOF+x7axfjMbROL9uKmZ34kMdDt3ZjZKANSbuTcZ
grWikXgonHrw3bLdYJ0D5s1230zckE5oGEqifKJG+hCXk7MStqncQmspqRXvz3OW
ejYfwf+dytQskUDO0v8uGERna1i/PFmhm8J6dQjKTA2x7zQXrz68hpzToSF4+M3H
JodF/RvTp9TZZ49OS927zynXltRyr+KPh30mAqVTxVeyXeRQmVTo2FyrgGDLtfRE
6Ddd+niDX3ZOwCLonEtn1VX+9wpk5q3no8oRR2uW6EQvpEmS+fOJtuT+mF+RoGvX
d+2vpJQqiDzGnMnCPcYu3Gj6VKN83FFZDe07DQrZWp7u1mpmqnRCF6F/VxtX9GJU
ihcE6FgVeeQj5ykIfrNk1+/6m8TJChPCUBHQVkpcXq9up3xI0Ena44q8686cWMey
Ztnrg3+vFUZlRqrSKtCab0o0h1uTEMBq9jx5AkEOpmCGCzC9zRodtBdCIINERa6v
r91n0lqMLjfuHcA4BCH3mJvKnDxfKr8c7+87Bt5XciJvVeU5ltMdmArF5OxeM9Iy
0c9mv9AA5wHxhpNKqm0EMSP5TcgXAKfI/U/vGyqk0kFfALsNnTi7Fu9Eo4qwz0QC
eFPtPzOFcpI6fFtht0X9epE5bMh1ZPPEVYE4NXJEPjzZ9iNyJknlqFDm7sxBNH61
wQIeMqI6zVb7/AHfjDYkp48IWNP/DYaHNDazLSrzi3u85dE7v1MPVSAWukyWeYz9
XiW4OtZOkGnQA/LvvhXxiQWV8cAqkum+OSyDIE3QXzMeeWEOq3BtVnDLsS4EbY6o
piTTQC5rc9xAtBk6PV7z5eSnjtf01m9IubiLtRqBHpMz24JUt6Xa95TczR89Iy36
Fg+x//J6DnYi4mpPqselFbX9635xxZIN7bp0+xhCAXKjS5j78lURc4OQr7lsRMjX
77bS2xIdeBGRYPe1XiB2P3CCWtaWiqHisajcC8SgLAugxjeuAYAZY8Pq7cQV6JK1
kHZs0IiMsLaaMye/zld9M4fUWJ4MnF3VLFB/pu1w9/m2M4Lsht1k3aRI+KjFQr2x
4zTIikrE9RN36XQNdgqd4z9DvLHrD3RUsAnjIrE5zEqjAVyLl9ZMaUO7DK8ICBrp
YBe6+QF+v6ysBU0ume3WM+GW2H0yMR6gtPoaHndtrusJTddoJX3IzzJ8oqdZ6ovf
pQAuMCvI/uzUZZhprnj6h7TpzZcjJbm0+TatdhIALm1kMXI9+gLP4IUR+Zy+tKbr
sLH4v6ifl9tsNS8ze39b6gNdHZvNr+R7B9l7yFqCSW1RFiqnDMtQdMe/bTx3lqO8
GEQU/3eZJKM9khTCsiJ0Fdw797drfYwyzQLVua4H/Rg35tiJ/tcePcf94r8rANsj
6llzmXdq0HM/EX7hHyxxjF7H9HoLcJVHo+CoBGxmz7oZk6ExVPBc1KUnqrms/YKi
eB8jiF1ou9IAWf8AT8qLWKan5CKoVc9QoaMu0Kn8z2iCSWmnEEDqA/wuEJImL6+b
UKcdMQVASMA7gD3Q/J2m3sPy8mNtVKSXEYAl40h//uECUGKhbZYb+Z3iuI5I1GtW
UcsNBkUS2e1O9vBD0u0Nbzm8R1trAfV+Ny6WqYUuXQXxZ6G3nTX2bUq6vfxIAFAi
W9O2PBhSrIV8bPh7AqChbA8on24faSyprk6Uq82xx5Na5DnY8PeObvc53RpGrg2Z
yHHNrNcMndNPXzmQR0B2yvsEtRnEuUyJLi6FiP/omsQ4dEVjR+WDtE1sZejxISOF
dmrgxzeLabxyc+zyImAuTa2C/445l2ZnXVcri9k2mJ5YE1r9BsO+AFSi2hqQZm8e
VaXYMFUGKNP2qK28uctH7ciRgW9d+SsDt2tOmODiG+LgWLcqqH0UQ/dj//Vj0q+N
B+a7nqeYiscPG/lrPyW6iQVK/uVAZ3gAaRXgQC4oDqE2jPg5Lrb2kT4chUkGg6Rg
Em3Ydb5by5PCrb0eYLi28GaR0TzbPWbq0t8P1lSQHw/cF6PZ/CaX7MS3zIClYufn
K08i5mLz0XOErC80e7+GX/LFNgRmS3odo4MT56DEbeFUcarWyDz/U35stjYDFRvg
fpirCmLDLWeCV9Lv5qjNlRxf4RWdP5MMxwek8bKBMlSTZbS/ij0Zo4F1CAVDdG3D
d/ovJ1OkKXLmR+pFmdJW1wMkZD3ZQQpUUTkSKokPwF6oLnfmI/HJyy0WSMou/O0T
DoikcYt+6SmKixH+o1qlHhZUx5M0NvHiY5F1sLrE6ybZdGIhCjCQiFD2Ph//0BYh
OTwTEbXq7nmlmOhHVjTI3qinHK765zdNgqZHoBQcPazneh9cvHMW2tInWnlfqUDW
3c6SW71M6/ZIOyQ58dprlosn3v/7m+wwfkLsGJbOqYl3H+HEXFdagZ2W70cdgVuZ
ZG0MUxlxEEdkXviIB8psYKGp0avHOsyvAZbDRegVs3v17lRD8oZZ/GeFvOZrvKtr
Z2rD6VBxju0GRtHEcEhBiHIgQCw4UEMufJITOqiBjWmqF+7UaVXpmsU6vAGk4UdZ
ZbytSxRaifPLpHeAces0xFSVnLO5BFdASciEt2E8EB3WE18vDu06ZI4uedOyXIUY
2Tv6bkXFJaEBjtP31aQ24acpiSLJv/WOPIN8Nt2xunjh+pQrAy5GOL+hJCUuPHBK
Wzno7wcDqHlOuWbx9gpaTVcoU9TqzeJUWhTiknD8bbdDp0reJaz9FZeEA+b7IzH0
Yg3jfl4sZNjRUmJtcidEmncHOSx/ntpapBp24rwSY0i+6imZw9oNcmYp0hCA1DHf
K8XrN+4FjwXZQUvabMe5Ko8YFHf0StwrCLyQvZS1ekJ6hnI31nDiUs06XcwzfW9G
7gZz2rk2EKsa9BlcQz7SVTFXGwUEfHHneldLc5fM78Yi78v1ikR5YaY6qOlp7SvT
P68u3RVfH6xuzjlxxsY2WHVcJ1kxwXeAChu5n2xZiW8BWrLBtUEQElf3E/je9tJN
mI475EOJ+u+b4Rvam6nr+bTkEJi4jPnt7tsNPcQTrMVQ4YL4cqhPkhsJdPxCeGOE
jojWj0YFu7WZ0hELLCcwW0dngs9h8autSDm/2/yaWU0kDZE3qz/8HixH3rH/KG/I
ab0MUxfFW8u9b5xRgk1zwf/lowZXPVu13QGuIOwV2lqgMcBTiqFf6tX0D6oHwW80
Bf7s2Y/RiUDd8YatXuWeIuxZAjNCshQAvc6gclR8pB/4bfRjJDP8N4aJdql0mGBt
Sf2U8WW0JMqa+jwGr1o5Boq23LalBBnd4pu8WB0/lKCihmkvWLH80u1W6amd5iuF
tOqW4sy1lBYJY3VbOeWzMQcqLBW7GB4fu6rmqST6MR535SjGrfxkp4l278kXZ4PQ
7RqtYPNix2SLcw2cxukEWsGnjzqVyBtEO0eBxbFGCIRXA/TtyyU2SRqtcFeaP917
7SMegX1IFWtZhkOHWx8gqasztNZEC4aPB2nVGnJGE4RL66ipnonT7mxfz1ydNesK
A97cpxrBg3LWgQJSxpdR473wCww3vL4y6BCxvF6Pz5uCqBemvvYwSOmrDiIcz2Ju
ZpDOmH1U6e+kuxZo6Inz4C1ytSzP8y3qllz016xTLliLVhjUxrtYZzAf7FHWmkUf
9iRK0r08NC38Kpq6DBisKvAOyF0VmexBxtiNvs4IOxTM+m6MRplkN+94q1S/AYL0
Rwk8yzhsqhMqZd95cy0qoTtRSmnAc0do9WbBwLO09nvVbM3EsFr7CwT+cDDCEOU/
7x3NBr7Q4BMxZrSOcjkICB0liwWj3S+qX+ZHRi6JqfK5a0R99VfJeDOd7qgXx9nZ
/TUU3jI6k3QMpjA9336mmPEG8VHWjo9bLSH/gnhcG9qNzHMqffPPFO9t7DEOQFMN
EKE6LkZopw6Fm3pJzlhmxfiWcwPRqE8hAJyYMpdaypVGcdCR8UBmRRiueWmwusN2
8Mv/FkkcMz+tyoPaV63b3xzXbHXInEWcPwzliz3jRYnM6S7fduDaR/POBrqqOtTK
5QIhRtuMbPoGUapCT5Wbq3NAV7WJ9iHsqjvsLw8aAyGJVoa96PLqErXNWQsM44py
9nMty2DpRj1IQlzWOfbvXbNsrluTzCWCLlNL048QXXrMRQAes8DAHsKIMWWwBx4G
sVjREbPft0Npw22quca3tMgxGmW59LceQMWaYloPf2SveSzk3AE/AWNmw+tbC03M
njfBP3C6dOg8nbAG2DVUYX0pvuxPGilNyRbUCmcYLk48rEXthXol9DeafoabtmgT
Er5RnIYae6T93gkI5TG0FWtxiMlRFCAS7JY2/2trTeu5Kpx6m7rCWqeoEpG3EjBT
UryRUe8Ap7VJ8laYkQAhlJeAIFAECSeqgy8EAkLgQul6yTdC5bE9ouC72FnrmOd+
l3hkKAJoomlXqDkVyA98vdzu48TVpJjZOPujlIfTI3NqFvVJBPmisrpKnLTiar1P
aLnim95xPN2FHiJxhPlkCU80nSn1ILTdVcPUXvjMti95ziQeT2OBRS5p8kqOCF0I
Fu6AZ54UlPMKjapT6/VnO+ojVgpK0069XpNRaob5i1qY2BHULZQAiU5dCZvefljr
Spuz+7pChG3zk2SmB57vBlFpCRimv9in3KiOh1Jk1A7oQt8tuC6TM1Bc9HiBIcfZ
u1PLybKaWCPvf/h4lp9G6Cw2Q52jVvktFw+H6vdP45pLHC/74P1gjkHrDk+VpVtO
B87L/NEWzICxrdmlYaCKs3QA8cvBNN/Mzr6V364MopDufqurIV6Z5xKyPIUIM2TZ
z5V6gwHoeIl4wwBEmoJI6d5reCnfyLRR9RuJ/cl6ogrFkmb/umssmNhIThxcYoZ4
rngP/gpMrfUUUqLgmNO60tsUDcCm1MsvQICtl4Di4mdPN9lKwr7dC7CDifkT0Dlb
8zPHDWIy9zFgrcBSwkZNdT5dE9VzMFPKYWaTk94VXD1FMz6t60J8QP9dnlcFcHzz
BqFV4t9pNZ83m3Ikpz5lSl/DGuOlopTyBCt9DzLwerDDg2MFMgNMtk9eNGcAzN/j
o3+H9HF7wHa075rrytuTZ8PPWBWSpfz1aHC5MXkPIgx9axYTpsW7LtoUuUeE1vkR
ZwEAa2HOWRyFymKibdzLSyQPXm3fHCLPmqHwCjG7O72ZV9EtQtmuee3sleE+PQKY
jfmIfEh+uB9nmC1dcVtsm6ms1Xs45eRZNlyaOAR8VmR11nQFEuVSnk0WHKKjTAXE
RRqnAOj/+u9YhaLKEQ9LefKMDA9hyRkRkR5hHFFN7occJTNX9zEEjY63lNG5s4T1
Qjk1nTyAsSg0vdHBdWD6u7pWCVUgG7qv1WlO/T19XJBVewaSlckE17TmBTGjL0hD
29TT7KUYLuCdvyXacAQeL+DLOUUZqdSXo5NvvjeZqiORr0lc5xWN82O5kvj5htOW
wubNlE4QrYlJXeR5zQojpU0WjYj8tYbXoshbX9NvsQytUWJim/lABQgICzcyO0ux
GF5e0w8viWbLGnDO7Tpqaeef6ihgX8GnZt8NU/0C1MmIQcto0Q2EVmNzyB9w+wzU
f41iEXOaU40g5x2fPeSiFd9ggclUo3XszvArw9e8hXMr8jqDdMXYOiKZ6WDnHPyw
6Zyird51An3Di2AwxuDAyhOUxRTGs75B4LrG4XwHScJ5qob6uptrMZBmNpam6Mmn
2Y3Wy9aL50BJLVf/mrDO2LMb22GAbd5ORuXPOBLETXg4Dq49w31TeI10TTKnUUTI
Vi6iPjQyPSQGAkgNxAtHWAZNAS2Ye/2HslPzuXbplFViRF7cGp3u0NxqrzvUdv1/
pjKufLfZoB7c+Ul+2i5gl8XOefq8VFz+LSFnInjEr6kJCg9/IQ3y8VFcTa8DGxQO
QzVlwKhzWv9OyVVKpl6AOB1W3ptcPlr6CAkbYWMngsBn4plAUs/MrypUIQNh9Z5B
QKCZVMgcZjaIFunZO/Hz02sy1kJkV+d2qgxpCOVd9VEiFTNPbg+3H8saHXfUhWwH
oBpT/1S15jif9+8pSqEXJo2LzaH+buSdEWlBhhSLFohzZgdjFKDcNxQ3/9ddw46Q
dYKWkgOjmlt7UH0bVn3cMCOiNJY4QxEEl9WWsAxMxO81k5Qyt5R1U1epNCADWbPq
6Vvy+yqIbfu52OIsMjN0sPYAXTRooZZ1UCMBIu0yKblByS2hIfhPEwQ8T9B2VaAm
0LSzFtGh77kXYAzTpPvMvHqO2/KmqAmdYtAG2iO3h67KT//dIijOvZMwhBqq4hVu
Sx6mkGLvpX6snOqmNWp0/TT9tLQVPHsp60C6+CGo0pniO9YO0XE1bTJyOhuvKr59
0aEoQwVr0psV7gy87XdRU22Uy1dioOqlaoQaxcUi/B+QbPc+GKKWsKu9hCPuXd0B
KaL/NhgPFCmZswSPomq4RRPha0FjZ4nt3uwzSSOIixlvvDdURN6e64MtuzJe8QOR
wyiFRCkEA92BLllo0DjZeOItwRBM8vVtJcH4lQpJXeolfNCOWDqOfpcQHVdfUVps
X/1wEuoiCAO75JFcnttPm2WNkR56NSgFQPQ1IIf0iUeVdFcuEMQxQ6wz6QxJucqP
fGIyrJuu9ZfQNWB5dHdAkFKl6CnpgSmo1hBzI5sKfA3U3ES6i4X9JLc9+wmwDFUK
XIVhcsn/nkAHSKbb0hHOWteg435WLdGKDEUIHi/BEM2ztvISPQakkSNQqsoSq5E9
m9N+ZSAcWGNNFonCdbDwW3OS9vr2fPjgGHaQszxLx1rxBKqlZy6VPiKJFhGChiqg
m4lO91gXTIByxYn2Gj5rNtJ+UjhnUN2CBXdcdV1ngUKzq59AY/CZwX3OejDC1Sxh
wIgtLg39iHpkWel607GCRQbs5Ab71yLIJXR6vwTKFvN9B0BmPoOXk4HD3t3v+MTB
MsM+GKxJNQGr5woGcCensK8HzyxjwpS44kNCRaL3ZRMrZ1sFxTO7SC5yVdZSdHdE
RL0MOkkIRd/0vgV/rh/JPQSe2UU8BDwnqprYWAFQfvzAAgqviMkMnv4QGQCKhyO9
Ve59KUIb90bjTAxBXHDlPafCXS1Q/DQoUOx8NJFj+BNkvEyU+8pVihtVPejNiVt0
UbBlNomloYGn8/lpcVFJUb1eRqrfmPLdsfV0OmWFHU7vszQhWEAlkTVluhGJx/oB
efFBlLxBZ/Liwj5VJRCcSotOdrrAVNzLtw9IvhlBznLOQwOhfyBgT4zgiJ1Uhwdf
NIvpwHp/ARQXlI9PJ83gwnZOIYwFOjvbd4Ud65GnVjAVPWSC6pjpwnYIe5HDQVH0
3eqrlY4HZla+Wd2v1ZOIMygTevXVGeDtFhZ6w4r2pfMpiFcsDV/D6b1ldsLnHDKZ
RSJlUJvFXm7a9pg5HbSmz3Z5n/eS4E9GraeCkcPeyTVZA1Iwn+ub+iHfMtO9oTTd
zvfHy9qs6mcISERVB5t2mVzm3irzvZ/ieqM0i1Qzy+TvBxc52N0zjnqJmpy00via
kN/PzEwvA0J19i1FwoJ4/l/g1U2Fen4EswelnAwsPxbPJWuM0lNtYzjkRBUPMaNK
uwpc46EY8HaiYNbAk+PfoqR9+ukqXiiG9xvheiPGBYbZvC9RnyXkbnCpCbtWptXt
r/2KazEewdUNwrllQO+f6OPK6hWlYET/6nBCwPySeqe2s76YsJdMvi4ueDhm7RZJ
o6axBP4jkbNkom+GLtlwFp3Hug1mmE4gHOtNsQRQMYc64h0ncrhKlB1Ky2BZMke8
42ADsvoG4vq9Y8N/U+myxTbZipF2yU+D2R6mjL8vGy7YIyqUXJdrKEQlAXKrLr0x
1CVPCC5EcFzycmc3hY+DggJng+9wRRE0JNZ9TTEbdsUHEUMF+8a82A6OPE8D8vun
htCq2V0yh9Pi1elYd+LFNggMgaxUPiQ+aHbZOzvtpnSi1aX1xxtclF00PcjHPAPw
vbGMF8dJRKkjt2YA0iEi8J5P3814rCPKCy164X+OpMnWK+xZ5txcTMsYRt0cZyb5
UHV7zSIcohzdPetADK9lnR4Am60BR4jtrpPKeOEKw+qGgx9ZovNd6AfGF/dz9Aq3
+sYRW/YwR1l0YhH6UEmYl/55xEKibnqRKTfQ3u8EXJTDOn10cSba7CF4IPLc3Fmf
ZrGGKuPB0l2OpPkSDb5E419Wk0pCCxsPGJorqoJ+pJ3VcNS2+lt910/vyFpAXCKA
VmGpl5Y7CigJr3sE9hJdJxmhnAoabUiJbRV7Wt4FiWLY2EmTHlg1iotwcafUYkfP
5ZL5uWY/np2lcJ3uhdQ4KDr2Uvo2sMt59SfVFp4yik/zGWuofCxP6J3I+ZtqrfG2
DqZvEqnIArtrdDfhapbuo53DcS4cUxWE7bG13JEPn6cNDGzWPbK+y4ZHWP/4GM8Q
4LrHp82YTM/1PTdnvzffO2TwftUxBi3e8fpLJEA0RClys22I4EGMoNGEu07tWJpm
VhYTV+mAxKsXUT840e6iBax5HHDujJT5rHo9QBC4X/WAZB5UHKpOgCCqS9tTLpKc
BVlXEmCD3yXTCHLggtXwt2DFmrqSeK3PiTtEMlDrAFeZ/wr84cDxMQHX9Spxlv+Q
FH/HOK41e4sxgZK/nX9fYBQDApPPzHxpI9HWU/EIqS4xk46Ir699OizKZzLbomBr
Vz85+gkJwXVPRw6G4hY7JDWsZK6gJXgD5xtPzMEDWh9YjEAs9LD96MoG8i/Hl965
p3To0OGipTJXPm4xTPvDM6palzMKpGj9kKJiiwRoz4+2mtFHuUda3yFcustl9QcE
JEBNC9Fm3Bf0FVLNHcj/W7ek15+thEoXKsvMbLkaNH6fWB8YD40YvYUPeP4GqV0H
s3+jPsAttPPlt0KHQweRRgtvvYi41Vv4WE1sWunO+V1VxsVb5Ufo/CCSaPjjzecv
3XllrF3trztSA6wfFKWQ8LZRRtI46D+AltuoPyxLiFDmsh2kTUcuUx3TWtSM0MRk
GkJRaqjwazyMWYOsueWvwZbBhnq31a2jZl5COb2D5MWHSCYAtWQsM5hghQIETHhg
zSP3tCC6auqUjPBKvYnhZy1AQtIrTXAuGce0p8jgQ0KACPJB8qThgf6mY8b08sEZ
03jvKYZ+4FXAFsDi1pkB8RmJLaNuDJ08XChPM+6WHH7Ds6DuH/HDvUE5BqRxBG3M
iQBcZQogyJsONok6B5qx8uBYtoI2uXk+w+G4FhlSsWRng7MZCM1pP+Xwqdb2aBzo
q0WldyF1QtQy+phzZijH1E0VtHU6FsOjw++BojzetsOCUyyZcFAHMzWTNtGZtoM0
GD4FN4X6GX6+PhnDOHXdG8HlEIUfCpHpmdkZnbCBMiwhWDhI3ZkLP+jv/2iIJu36
NeYsB+a9PTga1CkC4tv2TmqQxLP+wNyskJDn4Uvz5e2ooNBf2z1Ou4pXYw7oM0q0
Ncr0KoAbp37bIsQBirLlrO8JeFBESTKLWHI4UkDNBH1W/b88GFWAvLF3za2WklWe
PqbhJsp+nwW6fv2OIM21QvMbK7bQ1/V2rSBxn9F5cTTHEEtsr9O2fwQS+HcFu1h0
ChloSj9nhuErA59EunpN/l/+pcVn82igwj39a1/nMsKrF6vqzLXeQsBqmYy5XDMb
2FfDr9xshuiMkVql1llaAp71DBdPNu9uTPRfkGC+jThUEEUWolLxrZ62Aj1b67PC
7S90POztuBTCUp9fXPF4+tkiBvCRfc7GF+JYh5VpG0UYbcU9Cli1lbpYIWFivfjj
z+6cn2qsyLiao70jJKxdCJcP9kin4EgWp1Pn+nM6nBJrkOatQFLILs4QcWDVaVNP
Ts4KEaOt/oG0rNcYRnOdCYrqoOevSfXS/VVXLV//BPBX6HfxLLKjQIh9RE4SWCvk
IJ9Rw1ULqmEd8P6xo8f1Tx4HnS1UTQ2Y85Ss5KXaTaESYgmWhycfhxyIJfQsMO47
0zDY0cS0HXOSsQHchLpB8Po5mzm3L8kul3p3eGUtAQ3DASqr3Q86tfaUsyvON1Eq
2ZimlFQKcOKaWFSplTwtJ2YjWqymXx8rJkzeTenYflVfo6ojB2JSyF3vYX8aP9k8
FgwI/F/TKARyb+2GllTY33DhR0Ea98qrv5OXESBPG9AZHglXaZDtXFiH5ahLGU6I
Np982/a/3NdJ3QHqySw71M8gCGdnjSMGf/3OAA2fTur2f7LfEWTSNnmflqmP3JPm
ZCzv3L/ZwElYTuIBYaQwdKwpREXJ5GS/7Im2E22OmVpfknGuhK7j11ELZzeRRTww
PGl6dw4JUYF1o5Bt8haiC5mEaY11NayN+F5/8NpS3A2T3J0tzVhwEYfFMKVqsZC9
Gm20Lw7VkvU+js3BaZaA+L7NQV/tyyLNicqYWsP5UyMiH+RlOnGnksyw1s9kBjLJ
0/HvF2U5HsuHMZ0gJeTmYPb6n+wRFKfvyMmN3IEMT+XFlvvPV0OMSr/RaHkLwW6j
1xpodlgTJc4kN0d9sJ5HTtTlp3ezHMimIzZF1/ZnmKhe4jgexZn/tB3Pw2GkRuiT
SiOPpEi4CZJFyOcS1c2mEsF4Tfmy+hqFA9oGiFgFTfaqt2xDOiVOXSYdgFul5gLZ
y6w5gwOYQ61l6cICCJXNAfPuNCtnTOCSSv9vJFQO5Bcpblh1Kt87gF/sLKo1u4v4
cfd3O5VwK376qfUN2Q6djr7uuwH7valBdwhzp25PSV/ikfA/NKVWOEl+/l7nhsAT
zv73EjvMUGwKE/1cPGHlBiOzLvr95sVqNphkY/gdrimsfRRXDjxvMccBrhTUsNFW
i/S8bxqW6xiQtidd+3pKNs3/BaJnhFrtdd4YI+UL33K6Zb0pIBupT2JvDCk9/xu8
YDEMtdfgJSAxXhfsoxHj8uxCkZuZJUUhi96xQ0482SJ80Ugy/ZQ/KktLf/VzXQH6
zduMtGDUeo1vohHpqodY8S3LI2A08XCD7+BMtRWY3TCE6sn4amybAsjLCxmBGqBl
LmQtD4UCCJKi6A13pgsaIfc4HMRdOxMA4MgORO9KNouK/hrY+wv9fIfrXYfDVwke
tPq65tpxGoGlcCBUWI7drG/WLxIJ7B4kTSEE2RnA+Altdoq5Du0sbtJtEMbE3YCe
1SUEEutYwzA7DB/SLlKEXpxriRJn1QSVYwKR26Mn/7B//qBcw3IKDSn+fTaagIwf
nBqk+sgOeeij3ok6hQ5hiCowscCpu113guYL1wpL4nAnt0pTPa9lFecEfPVK8nxK
hZkhcq99S+7l3dyPLsx1m9LixomjTPh+XnxpzQVRRmf8fYxwbJPt20HIfJH/9Nnl
yi1cFXJNhbLuRt9In6nltT4E5riyiBtZTq3sAW2boeFoz4eL686m4yiLz6G9mO6z
eeIkFsQHcu1TTi2ydzlu885nT1p2SNAQcelCrgRuegoHlm+MvLtpZPAYXRR3qeH/
MlLZfw3UIA33zdiUMwGfvub52Jtsfc4KdhqJAXo82cVtk++bu600toSU5TmgQGvQ
zg0FrBtcrzlDoujbgRKDAcR8lq0NbzTaAHU7m3SBEteql2hTCpglJlzFpmriMSs+
jG6XaxsE/p/dnRP32HJG6kcP/XV4kjk8y6JYseF5SFJPH55l4prZ0LziC1VDUUFc
UeL3R6Ms6bP3O+LjxbCXKRPJSmnwxkRboeL+KSjsMHvfSKDTpjvpXGBNtIpAQ97C
BuwaGnzn4oltCkrRbcHlyv+9V09hAiN+1RHrXpeq4RaX6j3wQRZJofotQWbKN/1j
MHT4Er0fuXC3kcauQs7+mL6uvqaASrWPLRn2x0UPUxSBaLR9WJhONCgc5w51feZC
Qssxs/N+D3SMeFadCz3SY1zOnQLxXXKlFYpEKzx9UnUirTD8SnIzHyeFxxUUNZNe
MX7z8rJuvuBtMT6Ke8j872/erjHtonLhgRPCszuqqjcnvy5hT+cCI017rM0Y7drs
0idNKGCBnQKDVU0crOm2hyThE0iqlSDMGw6obS76AbCAPdASzbI2SZ7GSMSK8/Qg
O2umo3HAcXmEfgEKss3nYD0J152Pdp8DfgjW3Q83ntkuGiazP36qwfsBnbKxfZ+4
S03bu7I7C0v9K7wrw12mUwX2I00SnvFQJoKbzPRjtS1KiTpATLEFJLlo1jruGGsH
aStoME5cAcqWO748wOnAa05MwJJWLMQ11GXXV6TeL7SrY080SBsqPyu8FAnmahE1
dBcERMIAnA/P7nRlvuecXmpHRw7ZjUCT/Gq1GItnzlA6pWdNRoybBWDFhj71HW4t
M76UA3e+oP1CdVLBNmnxF8DkEqhz9QeQpxKX2hzN4XOmkhAwGJx66JbitybJMnaU
0PaUdLBpozEvPQdxK8rTBwpayxAHJW2wvCSsk8OOnQaqseF5qEVs01vgF6IU4vTY
kcNUMmM/218EHrzmhN46MPkLWvmjbdHpgLujxJdYRPH0dSYebJlNhbEa0yVlzk4E
FQ25TeVsOcYqI8PEMCrtFhFCGEtOHYICeSDyU+KfBG4s11YWIR5T74APPiAMbHn/
u/pAt3qn1Gperg6bs0Z1n0uMUsUtZkI/RBtBR18r9MtN/HdCVhtMXAwxcMoezZBg
GrGgbdDgenr22qjrko2btv+2bI2CAiZUy048Hn5blQcLwTIQeY0bV6Gj6HSKVGUf
9bJvqXB2Iz/5xol945sbvcLV6nBw3kY+DGctpivB3m5UyDq+03Dv5m/VFv+PB2L2
9U1VV2sgLhwS2g0xA+NkdI5qyfXRtRWULKXPPfhbxrbyfBpUyjdPyC37imFoYE6h
U9YdGajqN7jLxZ2G+eiLsQ6XdsjgKC1I0we4bR+5uUHm46oe8168JVf5zXISPrwo
9KXhMQaEj64tAK1Dd2441bKB5yT3T7V6CvofOv0bBnVvciFaNEa0ZsNBbWDBSjv+
lKmjXbohQyAuj04xnu4xWj0VOCk6gsyZ17FIJbPTGGaDeXSN/lWErtkSqzN2rFkf
rW6ofzRGq1s9QxC5d+/rDubxGl5a2535GOqzenEem9ZvCgwuhvF3wkHlRCzwjtud
mQ6qV1B+8keqBXV32mEqULY2AWUGEC/0O8LJJuL6j5jhN7Uz0OWN+O+vzhsNo/ii
H9fQGtq6RuhsP9r1dxGGu5+lwA8b76T+cDk9pk6eK9A7x/9fGi3ny40B68si04rp
vtbZ8w/kQqizJQRtDFDbeueDy8r3JkLvqlPGWMHhijw3oZOjTTK6/rlt0r/NmR2B
bo4X/kT0ws7pJNMUrzkxUKcVozMOsfdRip4erMUPvp4qmqNl9rqX9TGDWwcXnoML
6Q5aWBYvhIIsg927RXjRql2uGw1KDQGbRQ5Alm1BRhLRpSr/H+wzxo7E4BT5Mgyi
VEQ8+mcUNPDBWkm/8zbbkzt5lCavMGzPMv43gRd6f6mR7JFn0mWYg3Ps36XvvXJw
xJzIYtgI/ATaKDYxwTUvkXmStm9JEhA49eh6rznQ2elYTLqR1W2/nfohIP0xnUux
t0nSdNfYF32vIroS8mci7mIt+yoE1xndJVbS7n3Wqb47X21tlLmHjgZXt4t3gcpj
WhTOciwor7hhhjerNxsaDDOCaMp10Nffo9rjqSRCDu8OTiO+wVp+ZA273yXnKFn+
SVqBIRnCrqdgLguPbrwil3kdvwlrN2TYVW9082ODxezt/RPGD2U92qjMqMDS14Hv
2oCZ94aR8+PIuUELqvWhD4NF3Q7xsB/FWIpalpgrTbF/zMqrzREGk6MOYB39xKGb
v5HJSK2V18Q7sdLnXHpJ7cceyArYyfm1v0kCmW5XWAI7lICpqI8/Cfi5jNSX9WhF
MGFHCgzuIavfzftgWacdBKiYpRovZ5LreczQIhTAJBtdmYEVd4hVajAca3W4/CZH
1fUH6ckVe/d4ixhAbLU0/abkLVCTJu1qy5Lfw9DWq1BS6LBDCoFgaYdSZvIFadNL
n4ZyC7qWq8V58YyAyEqNzHX+OpDStmogjrkFFJh6iy4QcLA4P+gY4F0LVLbAOOYN
G+gr5qeuUT1SdbwZ4SiE7i9QznhF4Y5GSOEzvLr+AtDABtlRsuYwEaG8p/UXTYrm
ln2m2OT662303+mXVj5dlg648me4ceLn6NvfQaA3uAYNXpiAIE15pJE8bwVSaLKA
71NeO0iCuk2BhAwpzY0/sFz0whd0VdO02WOB/QsHRx052JqxHpBEbbAriGJ6eVmO
4CwbRwVzKlDtBEJO2qiZp4L6hprt+R3AAWPXoU9JvBXscoDwMiaw9ky0tP3Ha8lQ
lXtRGKMjOFrttkF5SK3r0gJMYWa51XlEZUejI0SYWy4kG/ZdqaFDmN3P8r0B7Tsl
HX96ScB5JJBQghHyQrM30ujgf2gUVdsRFe7VKQxKORR8Z7dj/Eljg3IhADaMJTee
p0w9jnf+i1A95DjwvvqHxgGjwyeuSHNSRJtd1oT4A0iDUzAT8/DAusP0xhRT5Q3R
eKsgIvrIwjIo0ZtJBDdMv0teIgmTLkIiKrjonktM0K9gOzkzT0QnfZQjcpAXkEiN
l3yPLD95RDVTGWmKf/MgwOEm1x5H19DSBZODgwBH10KgQSyM2gaBPixKD108dnUy
pnvV6o4ojOxWZnWOtydEDszRX9g0MFdGCVC6oYLrbBbn4+kCkpwPWwUPHy7ujDxr
x8f2mPbFF+ec3+3FsBl6Nug/no1mhUAkjCbNab7ZwnjNyTMaRWzSL34Wi1A2c2Kz
GsObpprfbswzYgMPWYQgk6pGCA7MHEolvn5BtaPDf5Hfe7bvOYbd87B1Q2Oyxtt5
u2HNZ9zNjZoelA3pO9jTM5Xz97P4jYZiux0KV92643v7unQbYegAiU8V5r9U1FE3
7bCDzV9zxR7Qu2X8RHajn/GYgjKVxwzB5Spuzl8jFw+mOi+11Mkecz1oJxhwyxAI
p7euisCjdQ/L9IuFFf55aV3MHSjl1jGlLdkg10Qhmt2Mxm7BPppRfNBSr0+avL3/
0GJ91f/JSFC4wULZOr9m1YK0+jHGf4S36+R7XMtso1a6YFlz6qIYmlM6eQLOCVfz
U6E6x1amPoXOcK2llpiPJ+A4F5wSxO04uknZU3g9J1MbpF2C/ifd9gKz8id+wk4T
tUrFME/ccQMRwujJeaOpPA4S7MBP33DC5hj4xlb+/K54XZlq1ZRYJeW8Db+6M8nm
sdu+45n9Q1k3QYcopzzFU03nKR+jOKvcaeDduBEioxjpxkp6BJGdwGaKgZQvcgqd
yUc70gSAqT+2ui8Hjy7DOJGl9NtIRF7BXbMhGO28APkC788YJX1trAoEk6JaAu++
OAOCUyE+U6ohHZE0Zf8gCcjK1HIC/WuXnTzUv/nZZI5CJfUtcR7jMjgsscRVH9Ck
z27j0/qWclooa1G5AaAvZiNF9usTcB5iam2FDi0C5nF+rCEtRmNcFfDbKmbiZo4Q
MMEliNnAtPAlu/by8sMLLr8LmdiJLW3nvYlw53cvpQa3ZsJCYdxp40gmYeGp4kjN
oIeATzjDSzv7OOXhyeVMtM5l+moYeDiFz0Kp7f9wX4eo14bCawldbSpYspURdZ1d
5FXsWSLq0KrOk3odiA4mwUIu3gf34a8Axq0d9ho3ZukTLFuRZXXRPzO02yaY3Ld8
HfSUg1rl+kRTVOHQaVpI6WPUVGSF0VzKqVav4UKUwN4hKvcpYq0gKnzKQZm8i1uy
iI7sAq3v9cSe6KUBV4jOxJW90fvt4Sj9rHqmdLWRI09zh+ltEZC2fePyIubtwa+o
+FuCSKBzGWh9tl/SPjAXw9r3KXH4n+FvOkByn+EgN4QuuEuuEpK7FnVEhLIvfMdf
bllgnoPPGYJ3zAQUde7sKu/9x9wBHvLubV3c4X8GxRQmodq/19N8qgBVy6JwwGZj
nbGoasm7szdctCDUtQ5DNkygQBC1oBvksKJc5NudYRWqHX798xGUMaCZC8XVMmuf
ssAwakps7JMPhhnreATyM0MXpz6aG3hI+MR7jG/bXVzs1Dg6YRlNBK6esPqh5CSs
Vk1uCGsGYoFuYOGFs83NEinSVvR4/upeWqoO+irQuOa+I1I1dLiApSwy+NHpmqI1
to1TasVbxG6BScCYeBniJ38/7Uo2EcTeeePNrsEBiQq9zLF3fUfSQ/sga7EJj9yW
8H+CL6eR9ppEtO+IUOXACwxVTnl7R3tHcsli0s9evSmAsxxQfJsfV1uh72jgkSW4
JrNMZWuxVgMMy3NJhQtvsE4/g72woaJf0UubjEmE6sjaWsDRHw5vTKXxAN7nWGVi
X9K1GHyp4PNMyXyc2ifYtjlUwgPYF37aeOBL5ggX+zSKaGmbJCrPfI3zmArjfacH
kG5bPJNKmY0mx0s2Al3vEEymJHSC8CWl7nCLrsUeiWYQ+9APFBW04b4pc061srKI
YpSyxa1m1OPiVn/Jx7D25cPq2UXNzNZUhHg66bZ2E7nqicXcrHOmhmo3Jc8QpzYZ
1GBO/X/SH1llTJ4ya0vXafsDtM+8+EMuLIb93M0OxjxX51CVJ4Tue3TMpytp8XaW
RWHWvmyQNPtoStDpVV+Lnhwo+H03FnYHyvlsW6Bqhc2tHJEPKf+GgpgTWfsZhcxz
sT1z5LboNatmW+yjb0iIeyAP3kZDYrJ6mpSNZp+2AmKnd9pWPERxfGH0FGfkNbhv
56MCdN9PRx4g5Sy5RmZN6VbZhImjSEmGRGyPf0bXaGs/BVPHpkjZfzPYkKLT8pLK
dJRRK8wCCasmwnXEFU7y+p0IUB3D203BjsmE4xz8nNSulHD3fHSmv4D8783X067s
UUfYimA7X3qy4YE5yyDd4u8YRm91YY3a83C6XaWA0ZkP7WssXLCNKsTcaDcCx3/V
w/w9Zd0pB740bYwat3OPw44WHahxmUwYEEfMOnfnX5qRxQcE1fUmT285lL7rM/rT
VSpxrn/VZIUIq6ESsF6P8kplXi7sr5m0QtwjT4Q0/5QBpviT4hKmE4SCIJ4rQjpJ
KhP/Hon1Xg7F7z6MT70S9OO912MtLq75oev45sEaNTiyesZ38IEdtS2ajkiNs14G
fBN7YlQUbaf7tCVerG0HC7H2/f9EDceCWfAI1qnREnzlXVn6mG1IpbtK2IgX3jM7
95IPSPJYtuihLVzL4nimUksWmJjziBNKwZ5pfXXNKDnqhhgkDwy2brSF1Lmn1xOm
FLRqL/6LHd2XQ0ndgyzzL+uNETTIt0HlCZaU0fD4nVIDQgRbiwuhYplnkWph7pxC
hSXUONZNkCaIpLS6r92vlnYFqfyGzFwTyfN2lcGl+yY8XAGgUlvVoLrvSXQdXBeN
AG/5/yvekxxEIgF5nWHZBtzOoZ+YAoh2dF+t1SBoV1/TLD7Cgr91VHCR+FJwl4pm
GUKEnciUCHZ0ivK+OE/uUyZuLKUBqf/FdDwav7raYW0lLvswuredW+2u348B/wto
S2lkQfgSGsu9S9wMNHD4PcwrvuySFh3bHMgBSZxau/gjmiDaq3/Bw3MjwQx5/MJc
uZajiAwkR4WaLUW71LTC4mIKHYHgHKr1xehBS2cTOwStG/8KNky1maz+qPsj6gtQ
o5nvBdZkCg0exlK07AMYtmM9dJCehobe5kkMMxVI4D5jBaFYGq+nx5YCFQs3tu3p
gSmU/iPgQ8RTWpjTRrL002CSioLL9U/wWMtvI0uIagSpi9E/xWIUJhFg0MoaSjkI
ohN7/qzCfsd8umE7q/b1K/+JZA0/urKXS2v0k/zSvqTRk0VMo6EWfDacnO7f+chp
FToCAZs4mtfmdoZQiavQoGS53QmaxSHzCP0XEEwSJfEG8VQhpGpO7y100B28Yn/0
Ue15jhYtDtdgjC/1ZIMTz9ZFNBLAPTt9BPtq6sSBU0AiaZzp8M0V+BP7VF+bCxZW
KWN4URqd63WSQH70EWy8DyGyELlG6GlEp1ni4OPU4pHIkvfYLkkKgtU7k8R5Gpe0
BJZvotoyWd7iIpNZd6fU6P2vLhZg8pc0CqkpPX97+deuvZPMSp2/pxFwFLYZC8Uz
8jPPlLeP4wviP639TJpx3Zq4k2kbnCDTVW9bJo11rgQW/CJZoqp7issOWZiNUC6v
+0DgtbNo3t1/OVIFjD+yivRGwc+6HCXQzErXaeM0K5OHFXEu4RfvgsasBTsLHeYa
+fy++BSwZ/WYrXSXrEotLJ+kU0Z18x1d5deP0Hhv3p88cxnGR+s8a9/e0w9R9OFQ
yBrf1lA+fXWHpF6z8o1mOKh6l12UCi2l6CmGnIl2+ABmgCXNbDP9uDsR+e4XSuaB
E32FMWB5TMk9EwDb88XxGxor3KQ6c8cxa54wF7CAOc0vw7tCiO8w0kMHPW4GsSOu
Nifnj5vChuBd8kUXay/rTr+pKHrZcKTtJByTZonf0Ffh43UyBv/UjPsxYpX7dcFv
U8ZejAMbtmKdc0FEk31ODt4JIeQlHE2CltvK+NRLLtucBP+AuLT3S+uV0GG0Pgfe
VoYwDTp3Aeo9SC4kjkWkdR5Uo4OqMOvc3BLTXLTkVLo4rGkrj1lAC2k0xbC8qmIx
ll4kEWLVK3yIqjRgROyUuzh0nMTULxf/ed7qh/jcWds/5dqMtHKm9rz60Wb2I+AO
mUBz8f0mmFPNJCmD7EHdNm0LAzPar4QBNvtyjPO5ZA5GuJ2DUnQGa+SzdMVf3lmQ
UqeqSv69jUPg1Rc9WmUWtkFqcM0rZ/pzklLVXngKBNs3gXDJK4TdYnGYjbTzbY2C
EaeR20vif+x+IHOmxhZIi9gdabvFrtIowvRXkPdRUy8ejslZmk/CR72tGIj0Xwi3
bqRxcvE2Pp0zmsGcObv/IM1v/iKgUS0HpomO814OqQlvlLqjFlxUadIO6EozfyR9
whDobQZCt5Cwaljp6hnXd9Izip7wJZK2dsuqR1J+8G4mBPRzz4oDSUD9ybnYKciW
1/ZKAO35skypy1uzzz6Tt8DGa/U2IbCjsOqd1/J9s90RVKeHeon6EGtEQOl2C8rE
IL5/9SIDaqjVSZFopkwtcaznSFD6bpoOFBtSXzfAbSLMEBagxOGN0jxNXjUMw8Ls
rrbMETxadDZ3f5mCGMd+UmmGFOw0n+XgA4P8P03wq+6wo0ONN0UU67KumyUqoh4A
HRVHlfzGuYohyFoS4H6Z0kifMsDPDhgMzENzGC425IC6+TrXgq5Xus7mCi52UEb8
wq9BaXkYEIK7EpQZFZ0h2UvmZrfvUXMVGLASwmcx2qE8igzhJG/rxbnht0ftwTHe
nXybzT24WzuSiaSK0/nYSxBphIk2Mw2IIRXS5F5AqkZxzm+wiWcWGZSaeMtRQX2n
eyo9nLM+pRc/IkFjzzd5wd6Mq2DejcG1xX5wj57PPFiX2dWHmdXlaCD+4a/o85yG
hidiMUiX9w3/Q5ivs6A8cXW59lZsap3gbmcH/gkGDXkvDncTd3FERGwNt3w0QCp7
UTAe+AsLbpnEV5cJRgQB2UFA0zr6X//elB//f5H3XqQP9b10pnIjZHtQBtu/6iza
7DbxmHOjZWWUBWdPQMqTd9rACxkWckhMrqk1Nfo+pD+P1u39tgpZsxtNx6el4xLk
lFYiVMQzP9Clsg3ojtLQdYeMjYF0jFjdk1mLWPskR34cEVaAhaMRDOB4zTZtbRj3
yJGvbl7rHPJIWUes+K1Ww6bQUcBx6pw/ORQ8zDx5mo5CifrcbRJHmQV8Pz/RlSF6
qWt4py4Y8rZXNCMnCJoZhANELzC0bfP6wXHPWfzN6XpjYW2DaSCJKpUU96eRO1M3
iSue8FxmOB83gTfBrK9/OK6Cd2cL5AgMma0QCjha2kdgkSVS36h748nOL6Ws0A7U
tUOV2tfAa0EsEUhW4MeguvF1ERou7kmpKsQyq3z7+/fTp4aMJZC1h2/53nMr5OTt
fqR0quWCcqy8N7Gm+QbwZo0DH5XJ0+GbJQXMxYYvd6ih5LwNYhu4DyNhe5wSbd74
EQrNSjzzTHuhoHihmlkW/QWXbLywG4wvvcPpnJIN4PHULSbpmmOs5W6CEdeCckZS
x2Zo9WAKBTGRe469kk/O21t/SOurd+sxDYUSkTLRoiv8qOlhKiaboK4K1dp2i2Mi
kfRLnK54LJjRjyeH1WmW7rX5sahMSloNGqhKK8sjhAuLK/DhKB48vA0lryHGkQeW
ZdS5c2tbKlr59EqVbxPD6zORrxWQ1Elxiy1cIUDgsSqtL49w7XFy/kdJHHfi1j3P
Gd1FAnbLXoa3i7IHtiH9sFyavvZjn/yBK/RAtMKaUuiQtGCjriPGRv9HsRtC2Obp
T+YSmCzs1C7TkPpznTQvCPdG9GC4q2IFLEo08WJP9JN1OwEh0id3/rXQe90vZ6x9
+P6F4Ryjxu3RBww6LDTyLOxbqVUpJqNkf6W/yM7VozxxWrxTEevCzdEcckmXOF9J
8tHCU53sWqlWcATTptcQgwvOnwyqIM5Ge1p2/A/4QUHUH+EAyeLVs/4dgy/mvTdK
EtgeLyNiZLkgm5dLY7xSbL8UOm3ygSe0KT/K5sti/wo6ouSXCmAaqgRqR/crn93w
OXZpmzAs7DjQKB6AlSexM/UkpoPnuppMYZJkNoNCPQUP3kPF9W3XQmhTJ8itoRDu
U9TijQ4jqKrsvUpzq8Mxkew6uOrCuJGt5symCkUnIacekWnIs/B+rluPzEEFpoeE
1U06iRHtvpyf2epaesEVYHqMtkxMacqDfza4KIW4NqcPD+ZE+vKsUU6FycC/Wb8/
4ngqd9lVvC1XSK+ISVq1gwVq3AG0lryw84hAoYb77+txoCVtDnV1jwQTkrjaPDOD
JpoO9e1LGnNIW5jcckSXf95aGNfy8ndf4fcn9Z1wVhXo4y8Xdicbh1MpsAybJ5iA
DGKU/xaczQubbhN6Vp45A5cucoiMCCyExqnehfyNb0xKAz52zhkGg8vz193oGqJa
4NJrBIgi6Uw2ofHOkJRv8ZumJC332VRW89zHJg91F35HDw8u2rMgWfhV2OIIE5QG
MmVnYZO7DwxjbI7XoZXKFFlq4xAgsmo7mE5eF5DHuOA8IjhN/Vna+424WwRW9s5h
dph5Smlqd/tZBJ8yvXuYvWr03lwqmW9DDDrIXxvvYMbyzgCn8D2GmhYkEuRUn6A2
FAEsjHwQOS2YdR/Mo63utLHQnVVc61IBgnSqb7haamfUoHB3iqAEdPtuDTr9bxNr
ozCnK/tytec+4Sp+ZvtQE9fFuj1b0znqZn89nrP88onogq6rFY75zoUgOKJdtj+l
HXFxvQKgqe2vOFElNIfj1MXa2xsBAaKygGO1nxnbT7dvQbLuaPImnZmvfTkwCxXY
68/NIXie5Fk+zNw1uzhPpnwNIYz6LGpJFwATRNEmGTIaTOxVPQ0JQWUJkqVSlFEr
k4/1Cowg5u5dySAuVJ9uTpov2k4vPrq1Ay7jdXBiNqwJUaI1rwmPg33YfTSq4hZw
DYsuc/pcofjAXviZCVDptiXTioX8w9AWP8995L4V8Xw3wgjA37Lfi0JFHoHCl1AY
/ML+Qy6akbEID1aY+X/ihyo4QqNthFQ45Oq7IubbkrQmZ0qecWONHPQRt1LKpB6S
MMx8JLm4A2faxztJGOBgPSkK1YxS9OCvvTC7OrchDN6/eeWXrZfVwp/sVCIq1uXe
kZZ0CSjSgMPnnssvrR3+gni0EWxPiKUMAek7A0hV0gWE3UofqJRxKZWMu0dMD8Zc
G8IS1WWOCbjFz2slbsuvEICwnU7qmNskiLa6FFFj3Y7QDCejieP822PVtjLmTQBs
Jyu3fvzzW+9IPggS8rUigGbkf4kGcABmK/OhovPCwkEM2OZBBdamgU+hnk/SD1zW
tgp6+Fe7mA4zG7YxZJ5o92VVTDRQCJH2+g3Kj6RKtJmMUE0PHLw7xFEhSnIZzrrb
3YuEujqZajVVBMhb2TgetYRna7umwLQ8B6sxcdWGshpm+tSHO6OMyXRAdq+KtFOX
7c0bIr56vDtNkjBb6lEjxUnz8xLp6Rkp4IedLBF1FzcAwSWuhzR6boSPZugTwn86
zr5lksVNa2EbhPJm1WFRE0R/MWAyQhVeRCsYlOeqyaPVezpkpNqdZGs0wWJv6+f/
4NfPjlrf5C6hV8rQ3EhkpXPdqG2tL1TOXCWWBM0qOqjR+MVz6eCtmf5LbaXKYHrX
gtf+2gnHrP2LEF+1yRyJt0Wd0yZPVxudb8jE3DEvnvEDs01/4dUHEtIgnVGmAwgV
H2HazV7m0iNp011CeWLLSt/hjRUAyL3WsVPo1RvhPVhVnws39nPF2DVzXq94oMTy
lUOLE8vXjPN5u9uL1ugd7RD21lF66tgw5o3h9t8sk/PbY4aSuWuFHRyxHqmW/swx
GjuExAUWAAuQtTPrfuy+UxloVlFlu0qb4HwiaNtJq3S4ktlN5k8lz6lsTyg5rvvy
Sfmf2QVPj0iTMy+24DrIy22OSlYO0KLvYb2FrVo/806WQkRWxHiFhq0KxLJq8Bo6
DkQ3ikvuUR/e+OSMnn9gp6IjNSbGFQrvlnr74JRbNdeJskOq6DvEvX8JIP8QujKF
SiHoemggpHswzTTv6tVS0Pi6DrZ7YA37OvtwIlQ0NRPPCU8jR7iqbHRCVIFGFDY3
j7a/9ZMaGUwhzJXplctFM1APD4S/AiIdSlngINjWphNiXS6Oojd+hGKkaVUeeZWx
aMU2HiNwDJaWsUfYthHLc++rIpYcfClb9O50ZOXeF77dxGsdbiTVDVgqZcH6pOsd
svioZDBI8YiuzifJAvdfSBonMZD5j47e1naboknE22v9yrVu1H4FnpE6a/2XHF7P
0pSvoYkQW634jktxuM3oWHxpbQa/PDvPqgMlkzDAqRe/JWIc2zGVdCCiWCrLEN9E
CbDi6JwpqavKGTVqH+DHYRPapoUZPa7eS3zN3r8dCGwUJq1FlkzLYLeIrN1O7/pc
jOD6nLAj7pKNL9a+pJoQqIKL+5EKeZPEJH0KgbvylZuw7yAhYmcG27+EC2hNdM7x
NvwXmG2xbYGiW7SmQyteBqtGhftJedh8Tu4gx3jOTHB/tDi6+jk/H8CQ09IIoLok
H42jS8K/+31Gw81vUkl1acQq33tlve4diPTABDdbpuWX8knMGbiPRkmA9N+tRnpU
h4HGX9+Wjp3XLyJne2Mjmp6uhFiozW50gQ6ImV2TP+jOAOJ7aut9Q9yC+SdtfTNE
d03xRjyccyTXftbSTClL6KjNKM2un++aW8HhA9y6Xxz+F+TS0jkD/+HGTZUA0/D8
Q+4KEaAAmNF4i62LAyXMW+42B5MYVvEIVdo18/MaCccqf2PfcqKyVTVD7nkIxQxf
QWu/HfhqRFnkOMuTlmnfUxHpqmG8OgpulESfM7KE1bwpZn5RPLB4kZW/2DH83txo
laOxRhaWmjQHKzk7RchNhcO2pIPRghO2/D2QNWrNNPDL3UG35Py6NBAKyS0OCdhK
TumBH2ugVpxyyfbdjngIiOBhqC0NnVztSDXN8mJJcirZP0WOT/pn/clrp+V0cLwL
SwINFWKnEyc8SYwmEYqJnfuBYElcxdd47klawSCxIW3WdutSTS1XHYLXN9IK7h6W
XOJIM3rW/6HxVaZiUcqAtB0xmuK6E6apvyoX0S5qS2OIkk+OUR6GuEGm62GIQ4Ye
7Cheg47QqPMNESXkL+8+laNqXUCDxWrEES94xuq7JIvPcUBGJFuZMHhZMLAF0D/P
w1SRpGK//foLKznFxuLe2T1hEV++5E5pCwvfkpTyV3COl1q7/2uc3Qbmb9pLYQHC
6MgTvK/kzhRiz22yBxv60gVBBS3y/pNxhnYS0IVJ0fnPX3hsafaeuGY5D4UvPWmd
Z7PdhDgpndiN7cX/3lasTjGCNOB+QKhtPT50nskcwtwmzPG12TMjQmwDamrYxySa
Hv/7haGVwtBRQAeLsrgFaow5vdCTBrugcLdu9E0L9tXLlLJvU4FwaG09USB1ekow
BHUofpSO8RYaHRK1LtGVxcA3tRZPLPtiLwOv5EMkafyvXNFBXio+x0sgar/TFi9P
bh0EaASYR8EzPMU9rvJ0RwK1/HfI3pfHwrYnokxasJpCtC4RNuxZOlE1g5gYm//2
zXaxOuIuimETl9MZs8AP7aACdX9C/VBZIQY2w058PzKEfbk+/QEISI03v0hDSW6P
TuXoFSXdIXHVDhm6mRctA7xSy0f1aZ/cIqcwLXauzDpdoIBP3EWzMQpX8FyE727M
613MJzZcdOUI89rS+ktXXIKBW/Q+Nd8tlo0mB6/oEDluNxRpjxa+lQrnj3SY7LWK
evvahhu52jNjZQKnblL0SaWW1cT3Sd+1sZ0aVHm/qHDeK8wcyJwm0AFPmWII5Eyb
4spQvwMI0mtwRYW0XxowxE8WHdNUPTfMxYi350NHkkfdTlJS+hurFfJ+vbVl1Kli
4zZiLrWPpQbuVZQDCg7bIqL+szWRGLhVji+CAcVlY8odOxlDJ3fmwI66SyoDLW+Y
mqtmlIhKCxLfs+DSp2h7PUfsGZgzisnkuzd9xZGXL8zNx2fDmo9o7TDk5I7kjn02
b2KAJ3HBErqydKohBJvTY5Njr/nlduzicJ4Yga70qUdzJ1NMniMn9jq00QsVAB0P
2Yvt07rb5TiD9YQ+Rfp8jEdlfSwyyX0fKtUyS9mCbBzAXgFmKCFqLhwr0Q9D8Nkg
Rs+yJsyCZVBqJIMjeXPRjtoLZv89CtgNiULxiQqVrl6shsn689KCn6UmEXDk+Sfm
NMNFsojrvUXt2IfAlosr0SfjUX6qO5Fal/pcgl/u5HWnqXOyEyGKnVSaBQf4/Rop
ZalhI0s/pImGAWmOBeeDlBd/Spkn7kj6zXnmIzW+OXoS4dpYCxD2Zg1Suq5fHt0d
1H1AUohXyIVMz3hIYd//ZKDXMWlu58jMhhvIz8lHgb9QjuMT2UgcpLbzBHW8+Jdt
LZavDWoTBYQFdkS+1P1iI7lfN/G0B7jdbSnJBh2WZep0leg5l7EPbhZCmPUq/TWe
S280bi4n5PQ6bNOPoEiRXQV4NzuxHIPpKV1RPcvCOkgZ9QKAdzWllVj6isVHORlx
6u0E1T5blFj98+tzfaQL23Dru89GqkmzwktknJLHmv6Urb7QGSknkyu+DKbEWBig
ri0hsz2qK5+2RHqCH+pkCRWrN9IgKdqpgbwRWTQlnj5hyFzu6plO7gIwOTgWsEys
znJnM28F2SVvYY2yUzze1Y5etmesyq8Q/6rjbwnlNpYqM0jnDmzyrOiQ4Uc5F4f0
D87WyHhdwnbt+GwmfXYgaV69f8cVpZWjOxgMoJ8xdCE+RCNNa7ViPfBKmRbGW+Je
eCTFUUbRCLyzJYw2XCdxIPwHZqtIxDs8ZsSA2SAs11LmjEiIBOuEcR3UaS9KX1Nn
enmWx5Jd3zCP7wA2pXd//u6lQnfG0FwdO/r8aEmS1WfiuX9EXR9tJNL+xrHpYH/c
vBF1yndI7cG01L86MDij4XFsmmMxNl0M89s9W1Wb90Xu+8yc0qaG8zLJtJ3nyuKJ
6rsQ7ox0grvzsw1DPoiI9BSN/r127rVER+AE5D1smh/G+xSfpX6QBaErb98iVqkf
lUIGFxd3czSrWdsc9J7UaTvPKd+UJA1+kw+8aqBKg6RbNns8SlAl4i1dVH/8TN+o
BuQtEdgAA4bkhH105CVvdBNYag7Uv2GJIxm2S8UDvA5DltcykaVFx0plmQxacxpx
vEQLJxLrUGmEpyayLs4UyxTbREgWifJHJHkyI2TKAMgkXAQLlWL0ztVJ6EfDZBtz
LKaull2XQ0XnrgQYIwpQhirC1IHxmxjWPKlw7LCOfQBs0gB4HIg3BgRxg7LhqnEv
6zKt/fpHzSFLRlZoATl73OX4En86y1WGmxBlvXyRVlQPBSa8soSgjuBWC9pVrbsE
e8j+cA4l/q8jk+xAkUtOVNEAfWKA/8hIKm2/g/ruTs+Jj4GwgcTldAcD5WAWRH/B
sTTRszMnrjrfmMYjoHEWhXZMKGK0vzfygskydYeeLFpVZAbOSo8dLXluQvylHqJo
eNhCTIzXSZjjBO8lzxzkapzwVTZWhlfMbtp/N63BoA6Wa2mZdbu5KN4lZB0JFFjs
Jvx2qF/JTTli10/0P4hhLAtEAKsKBrIlfoS3jRwxD0edioZXfnvN4veC7YqNj+VL
yU3iKBeiTeBeqQCCqHJ8aN5zZLoB8/YGL16VlVvbQCZ41Fm1NUScdFaAPnQxABtc
lHMnvS+Cn97DRtRz77mSlr1QILg714QXa9cztzWJvD2gsB/KDwEy23F4oHSjDT4n
8GSR6ZG3gh7lsWWqXHttjXMS+QjbdWFmH+RImL4OcfkkPc7iTDsb2JB5494X9w2G
QFTdyi1WWn/UDUUXumqZ91RN0qj29tAuBgGgMqbS80UuYX+WQW3BXDkvHVsjNzfk
ntGpkxTdcy+JbpPkW0p8qY0FDN/i/U+mDL8dyDcW5F8Zb4zsDKvp6tWFKeudFda2
aEUQ+DsJ9etcl6oiiAVQsZlpeHCXBhsn6MC92gDB1Gjh71q5xR3tz9Qxb5nPwbWZ
OOQcmL0QZFWXNHU2uwguC1Cz1kQCn933LNSeWX5RypZJ+dsQvwXuCQBbJi68vCBS
+flHj52cg6hc46rxz2tDcphjyd7CWc6BKJhHWCHB/hrXJUJ4mL1vlfqav43Dvy1j
VXyewo0w7Hv2M9vCixQVlvM9UmGYKp5N2iIxGXWJSVzhNYQYd2G/JyK+7UJ2cX4l
qJ9d64QfQSauvU0TCs2W/27Uiq97Wl7gxPL1mBinRCFuZ0uWrnZwIWBGDFDJfbbL
c+6NE1dIcO7nBfKpUs9H9PHnkBJge4qkelhQl7J54XIy3+m/HGe/UaWzVQth5vEN
EHZV2/EIO1Yhuu1Pd9XnT0FDiHp5S+f825Rlk9EXv0hacuimLee2mwVxnzz55y6/
P6G4LTWbv1ATFV8zzrf58DKVfLtqdsF2eXp4cGerwi1fNynpcwdH22IV+IFkP0gS
S8mVHPcq58KwZmMK+3KXBzDS8ZQpdEUe9gfaHzYiRXDGmQDTLwXH0qChqk+lSrYA
skSycKYvAM/uPFojyAPe0yclWlKzWiqv8X24MWUHnJWm7FUVtHKyExBlCscqxtEo
91U9ovE0H2Y8ri5SKko4EiWCGStJZHrH2WjN14dfOUCbP7zQBvoTySCkzrk8gtH9
x5vdgbVqEAp3AS2B041Aa2lQ3Ur4u/M24cBYNWvX/rXrQMvN9XbTojIUDM8t+GRy
5yC2y8fV/VnKmtmVXwLbKB9X/i/ofPS/opwa6D0d4+dNXWEJ/W31OLa9nfPpb614
ewBWp5G5QyZ0odCqMMw0bCc47oqp6ecZZVvzAMr0NINsOlQqXMdBrJvJV6q8tDZy
uW9W4w2rC5ihFkoSoEwNMzEL3jtfZwGHvAC+lIJ/lH0nHQ06TZ5dzCe0irGoq+tQ
6YgnoMdFewokOgA/A88eAIqpY0Rr2XbcE57GLvHf/wWjV9virGkH4zoFlwTJ5wUK
aPx6fNoDM+HMudyoErujw+ogJrGUd9otgn0NHh+oKxnl0u6gJQP98qcOh7ee28l6
Mk72MD+0RzhTW2bk8DnygV5eouTxicJsbJvol/BA0647AhrSZosfNGsdmIVvtvnG
gy+uOKsdQpnqnPzv+0mqFJTa3KgXDpqMrONqD/5lADAKCY7BEluEKhQrkGUibVQ6
Uz+8RHKBJCjHQ9n95OKXAQLtq+aeIrIdMSpW6AVk4g5TBKqJecwIGFQLkdsIYTNF
LWp4wKgBJnnzsLHjsyUoT8bZutC60OZ9Wdx63t5E+35n0Zb4ks7V4861fkeD0mar
poEKc2c3FDDTslGs8IVkl9EcDkFntMxvr0W0qhA3E55KaUNyxUnXLWXdClpg0EL6
2hTKCI5CDTOwX4wOoXbF5ieHoGigZGBVuD/fPuvq847lHgQQPdN+tj5QgQk3mMz8
MQX8Kjs1pLq+ib/0NthBro0zDY3SXds0WRMkdzQDNTmP4309sb5P6qfLFFIurAHs
dxzHT3ncf9i77S3qnGx5erm1vd2UN6cL29OVOoMiAReBZMohMa5a7wgFreJeu8PB
/hapUzyMuvwUjR/6N4RgaOeOsf6YJrkJLvKEjo2eWGPYJP9q/e0JVOwyZ6rpJfcm
rOy1M/jH9dTltxRrV2eHonMUYpE2ByOL+9z/t1FoooJbA2APXirU/bP/4KNJqW5V
x/gCYeJ3GUkuwNSKvmZYwqBbYDZ3F5E8z6zL25sGFX/JV+teCSeV9uhjgc7PxTEL
+Yv5wkD00Xrt3ZltpXnT3kQsuj/ewjLAoyPHJnhncLQ4EEugO3JdlJq9xqufxoel
ixlKdZNb2tP8Qn9wAAIVwQH9DRWjeOs1aXRTXz0h4D1l1P5oc0BP6DFeRAneLC42
bSvpi4pKNbN5bnXqjhVPpFCuDQlcJGlbxyxXoP5bXCCfjvJ1tp6CBdTXtHK25T3j
z/6K7evusGNRcyNR/huj84u06j2ZPGhHOaWtYcIHLTA9nqhHby2O6OqWZ1S+JdWh
pvaAs/J2dRFD7uJg+Lzhdgu2Rib6BFgODASUFUKIbk868fCRyULiLMOmeyihyMtn
mrVPT6TnYbFh51PCwX/X8xFfaciKPoZfun5rQ0+DX5EkIXl/CP1gs+QtJCMBO4eb
KZvbUWYZwv/QpJJzMAXw4RS5vo8okuwb3cuciYfrBQSgnjADZ7+Hq0UbmgnErXMC
fH9yOY4qQhUPi9OiBr8GeBYa7OtaClV4DfMpWWOnYpg7dJWHjykgTBVBmPFadSAm
g5vVrNrf62vUBdJHdIqPs04GMMcvc9bf/f45aOC3SbQbOnJZcaTgrFp5VwRt1gB7
KNtqFp5KfHtWl+Vvsq9sXQFQPzbL1NF6b3qrhIBgk6K2MCBN/82/ghHvOOYxV9k/
tugdhySBk4gvYexd5wOZug+tzy4GWFtQ9ayOzOeLkjyWRTfduZc5cuglmKI4KLZM
5WjRpmt5PZa6L15UJuGGkFsJaclnu7H85aaPmBI3llD68gDxjJBmad8uApA45mXk
Y7FjBebKM5Z8GfmDtj5eNWInnPrWD2AHc/lE/fCxownBYOmo2xFyrIXraup+yY2b
GL9PyA3PQLPkGp18dWP8XogNKPJJhkJVvTAI0GAvQQyZ2aUG2l0NTIN0iZJ9dlWC
ppi7rCs3feAHILacyv7pW8RTsw4HeZsNvmDwNXfJVxFF8MSDuUGiXPlDHXsTyhlU
73iqjkOAANEplwL8rcEG6uVBTqWvvTkPWqS21HkkGN6GNsOK+0SwD7uUnWYhMofO
mrjw2v8BfIctx5rd8tQxjh0W3L8CyOESVmVZvQ4phaxbwTqnlGEfzaUlrco37qaT
pZtJv8uREBtCyUMH8/Z5l/NyHyCu66jgXgHMSQy+NxMzq1/pHfC9IXKr760N85Zw
cRxEHH8iugmUa4Z43MpkazHRYlNdvo32sybYtQPS0st1Urqjv9L75jU9I43I7qFV
A8M+Trfi/g+sEKxSof7oZD/984ZJD+pLBDDI5F1yayTO/8PGV54exY8HkKwd3vg2
eKC8QwbYCH/omDPvnC+XwC3W6ON3hQub/IjwZIH3wwWmZUoGZwSmIUNccGIY1FrI
E1wZjK9o7hSezyz+t8rIchLUV/jP7FUokPcOtls4CFukgxhtA8TdMkznyLMP04CP
DxAH2CS5MsZMzxcFbCwXfgtvNHiT5nd//AGcjO/D3vjakLpFQKv+oXHOBRCgcwXX
TnuUzKOpgNo4Rz5HSZOxgAcnzNcplzdKHBs8J/1obF6FKoC3yjd6MWdLQKChX5JR
eOL0YlCeaOf4h+9Pi6YMLVC903rNyCvT2ANcQrCQ0B8x5cw4fo9hVP/dXHHICuPN
LPzFXxxObwkpziM5O+6e5ZXxCgoo1vNdcUV2VHPNbyIHM8FqVOPqv9pmCZODFn43
UDtcmaR/5XdmEuX2SLIovGX6YTjTVeS/xDKXaSzmUg3hHTzU804toi8CQx3TCJHw
1MG24/NPYQZ0agQqp3MHIHLZO8soAcmLj8+4h6/SOzphNUvbW1JCjex0u5e42zCI
hhWviI7QA8fvsKzf35p3fV+ncM0XdbflS2kjj2mTBNsKtZ3lV+Q/ZyU22nbU8igs
8XMN+KQHOj0Sni7pcQkooNKU19CtgAsBwUfcL6TKus7GYYOii/N47bAJLeXr1cxa
haZnTmRpqU7f0k8k39EQd72XBb3B1nQuqwVMI4a8VNoNxOGGYmMbjKtkxA54wuTm
QXCyrmuAdm0Q3HlLkkG3rQfCKSG1CURHhr0/JAZ6IF80Kgw5u5b9pA3MvMkyeVeE
JZQxb04LXRESwBnYK+ptbIzaeP9lD6Eo6krkyQ3tJg50EIaYhR7MRQZCGkISzLpE
ZFNyPyc8qM5XI3Ak6wYj/6LZn806fyWA6rieAjr2Lh8arregJrIjPgwgnlQBoXO7
CCuuL0yxbibxGxqyeFq70BH7wW3X79NAJ6ON2A4tKymAn6JZ9Hf8s5TzffoiErj0
D/+45tvl2xrh1jemfGoHpffVZHHFlB6ai9c/faCz4MElFgv9NxjTa3V5SIRKCjdw
WEPds+18Lp/l6BZSuPrw12HREno9rAlA/FMahfZ2C2K44XhUvvs8XvKGNv8KsgQC
N+MCNobuH/JnXe27MLzPZGqzJGb1/n8pUbX5DXtBBpbRIILSevJd6cP2H8MEHaNP
4UrOeP1EQL22SgijpuwcXFBXspIOrAJe2IUqVbrUEGuK9abJC/QF0zTN6Nsf39FX
aVYdITqdb5DENkqeZtwnhvMyJ7Ev4BuiwnEJlmqCQOhgw3LvVchJjNjgLGwiJnIX
ErhpxVzVwOL0IUh+QRY5GS3HSY8YUGm6/V0e1TWOwUq32myNQExW2fql+2BUi8/4
/GI7gUNuL/j9+bRywFgvXKhaAWZeiyh+bZsmvBVr+dWxtwxm7FBj1DaakeK0Wcae
SSBBKPoOecsxjuDTTo9nEG/kvh+44zg35/ttRweIhaMqTQQgQIjyx5UiWFLkqWrA
penUHP8Lk2MssicK2YzzDYe9jnFAwIUdZqGGquJmz/onZD3LM7cADaiLgMQpds6o
CihJFpA6S0c6vTOkQLIt6bPXYwD5FRxXvN/JaQBDYGL2m/hwfWWcLnPnOSuECvPC
zrAxko8KAp06/hIzjbsmHFSRVhtXckiUPABB83dZ+bsDxes6q58vWyIYFylRYrZz
Hm77Fd5c22bzLdTEvQRsb8SC79gSHpkGEiqLnG/v00dV/erb3uYG5+5eQCYx6ukm
XEhzQ7DT5vS4P2DGx4Lweuh3qwWejEfL+KgR2tIEiXEnHeEF8XsUu28vEn5x1V+c
VFlSmijNZxTspWJnziojG8CpAMPbQEVjMr6lEbi8e9LUd0kWx9MmQ3cvi0wUcYUl
EW8pp4W9Bs+mDmDv8u7NfXv8LCUqXiIsUFZy0EMHQCv1+PccWyPxuZVWtdJQxCuX
s9SAnbPk6OoBea7F87Ej/hd9AxT6QsAhgwnewiSciBHCUdgPstl5QTszWj2XrDGb
xNPgmIcZcr7m7JfzSBDFlyafbojw964fVltREO+sGrlom9N3hWyZe38upiUF46BY
h8GdBcBy5/NVU8lYiRCzHAM/TiQDrqi2HR1vEA+/aSr8/vLh4A89ZQyy7SP28IvU
KoEF82ZXQ+Pp/u9IpJX3RtuR3YGqG2iA5cyEfmJ911w06Ov6aM58X81cXJE28Pb1
XMCiTjjH5u7W7YcZWF70QA5PPKSm7MIVt18e7a3gZ6uVmb4GkoO5QqgihsmcEdsK
lGh+z+ET1p38xjgpbT4gon1oTkP60nLSTNOuMkdLH8miE01sZFR8KBoPOMDjTnSK
NNwgfpWP8+ZoM8UruqPpWc40+TWwE9osBMABOgg/hwhwLn8Uhe4Q3dBYuJr+lnTL
nQDWsIlZbfimrkD2faouE28+kE49r/hZMlxhuF0GlCCTaZbRNjBjMgZ7xGWKogGO
ejDkdQJ82EM+jEby8txwtwiUARBrgFz6JGC7Dv/lG2FfFuQ3qy8CBjWIHuPXtzuo
PSwD8ScLuxgLjQTE4wHPDOdxfVb+CgO/E9gRiZ75dYOVKYRv6sfhiXwEe1MFpOh7
hiR+W7ip8CltkRqzPf45IqIGfdekRHJpuDW0Yck6022tyTZGKmwgo5TsWugCyfTX
pbdlfuVOI/raY5e4kne0dp4HZgq1Q1Yd9DJ2AIAMnGtZIDNgRjEe81SLj/VVL0kj
Qw5ZqeaVH0hmmbehS34RmEw5+IlQtou4M8Mq/P4RM3ppfsDx6i4ZeTzJi3azM7HA
i/rWeFoFkrE7n2yHgMENwnfwkjSpPnwqql9yGMLMsm8UgsGLE5NIG7xxEia+ZQ9K
fcIk6hUkkVfhYOWEc3LblItaBS9TIyHRnFAZBE2wqNrvgmZWLjR7oktpUrSSyuPE
jIMitnovsPYLOLynEnXhJBc/av5NlaDuV96uVmrT6w0Omes457wOi0B3kbldEsgV
W72SEehio1mZpO3/LHqxGujTX7zPqNOABdB74lhvWG/ZXi7feExGhdnbYTDl56mv
RRufe2I+T3U13Jcc+0rCT96H4RBVBMzdU54DSCK9fmVfWZ8cduUbwgadb9vFzqv7
8Ux9C7tZxvnUrb3vm5DSjxuerLiY2QYp/8NHC/3yLwArlDEpha9ODnjJLw5nz4T4
j0IPngwuON0A0IS5E8PlHJUU6wUoOe7+7oZZ2UTRh6zgE7ceorJJWzB+OgRe2/sE
J4zKHK/PSo8jLN7TF4VgaoaujRqfvqWcmLZe4l7CxrDy9Fk9BH9S+uKET3jNiTn+
NnOibbK9fb44EVgefhswJfm3fTMeviQlCdwTyJQzbCIzRj9FQdrokrZfT3ZnNfFQ
9S9jsillAEJ+Wl2lb2UTEAZsgwl8GxX5/X4Uw/pCxArIGmW4/p+2BrEE1iIvsw1m
xFQwjZvA4WLO+tqEdK3kFk704JuTSzy/786tbOCwMz/L6KkgXW+4jxu2PgWdIC8m
eg3xFLOlrYnE0bT+QintpYnJfEpdFc5WU+DktEBoYZ4Qr0dO/JF5c8RUrq8F2ipa
3cN8MArnVN1pBecOzP2lphHS/WnRG3wWvPPUCZPx79DoRrJSZil9ENVKw6ooH5KR
HsG7epWN7Ejj64TnQDJ8jFF5CGhQ2R7430EUzl8Fhn23stqqBMdn5uhekHFPQjX/
Frgjd9z9pBZaIW9p8NE2HSiYeY4LU3QQMxTXPQ4oaoz+I+/sT1ZnV5Q3yWbDXM2r
7xTKWFYZWPmDIU5nqkbjeTqu5T3HpRtld4NbX4PwfjMTIGBOx3FcVgwhN/tXewGp
zUINAC7Rd+2hbVoM/ZMvUoqjtHqybUfat1rt7CzrRE15IdUno+kblP55bpM2sDDK
O+diY3FZNVktF2bk+mJnff6XoAWbxJ65k1uZn1HVhQtLvyP8N3Yc7qjD7r1FbNvI
z7JBfelUrlxXeF2sZLtgRvzplDwCNdzfqg2g7XGMLiAseq1qigVXmlpk7JuYq3MF
sPd55BhhCXWO2HqdphvOQRCY6RyytV6m/q3h4HjvpDDb3ZSuTNla9fTaZS4p2uwN
bOSbkzCc88nbIjM1ZMWg6R3/D0jfUwx6R5aAamxdYBl4E2F3570HhEiNP0x9B0YY
k2lPQ3D2sZ9jtKeo/qkeX/kAKCaOaWhkkRHuphzHkidZQJMjSun6v99EYpEYmEwS
WfitPhvd1gpQTMa4vHKJ7K95eo89uekBuirEl7+YIR0D1hwTTKtl0uEIjOb31vUX
aNVZ2eCd3T1cjQSzWSPRj9wvyoKH2kNvvSSuKllxm9PjJ/lL4ZJxPyky1mbuA9fc
xE15eBg8Ex++R7vjUZo3yKPxQ6WDUbtL9c78nWiwpCm7ALL1iYalOr3tu4VKR9+k
loCZBbkC9J0F4Zl1IrZLYWDma3O3RO60cdY1SyadKxOTQkbWRXnWSc+45VbZdru4
gd4rEIhVz/+pWL2kOB06ZFX1H5b/P50vdxdj0DJUjoJYOCtIm5RR4Jrpe0pLrCQG
cLWVZyAfZhO/aILuXv773YzGIV2+zz0E8Z2GPFGKoh7xX5/bJv7O9Vb13GOmU+dQ
GsW2cXH5GOEiuPJVMRuUg4/si2j6zXTGnGBcM0DWe2mM7i11pTcskrRltS8aN9jz
fela3V3hPWLf1bSB3B71K7K68wZX31thAgw6pxGTzTnavMI615WCd79jOn7MXZWY
ReEmvbdSjrH7OFyTwOWusP9TH2+NGjUtG0fgIIRY1dWfLRjtjMGIGw++hwKmmu+d
1O34OH0UuFxfX9Cu3BQmiMijCqVbevlyEhmmxoCuAK9UjaVlAv6mtdK02zPMb4tw
5SQ/WLtvfsTebjJDNWITT/VjJ2xikRyB74YoEeZUNtmLJ8qaKM2c9e90qJ5nPHPK
UVgvSUgCj6c1STXpwOGpIzlpchNHhB+DCjk3z4gnmtaN54cWBWYCW81Fz4IKOdmJ
EnRDTVqeKu/5/xd3f62I8kgxL5s/aeQx64LbwUy/51XlVGjge0ZWUZDGF+TmyscN
qo5biUjBWVYJl3BLDyalSDe3Gq0lr0En5Y9/PBNgiJPujST08BCpNLxjuzoOu+S9
pqdLY/PqztnF+jmLDAepiIdd9j51tzhVgLqmegFn3tFxrRg46rg4baiHUTg+WE9/
CCKws5rNEUDKoabzpEQkr+3zjfjaDXWLTvJCUfJAuZqI/Co8xQHmYnWQAlHyavxa
Z1lDBKzq5HEPHc/9ahQx8IlyA9b3K/MYC/yv4eQBPatufkDkwA4xXRaqN+L8Ibk+
LhDMz5ZV/vunngox6St3tgsYRwxtyBcYF+wR1FxOMu5s5ZJ+JEHJQ4EKDsDhxIEA
1FNVl81xUDwqAUXaOyGJqfSq+MOwEvaXJCEF0t9lDGOZRT1SzHFKnz6+NfXvujBF
BSvPiLCxu4f4GXQWeXKyr935gKiCxkkX20OMPEHMW9uG0b/lgA7nKSyVaQEgexkM
mCBA9lCFopL4fthJ18ivNp49YgmoGXEoj0Pdx8O5Uv+Mi8UHGjzSQB8iaAJG10y9
JQrcuo5yQxiWUi9DTpjKGreo5nldk5WIM1Rp8ijgSd244kATD7Ix4McH18WDo/Qa
UIzJLSWqKZyJEvMG3ZfZVwQM5HEoViz8ufB5Sk3KHpIBtFr+Pzbm+wxuK7oPAm+o
lbG2P7PSkVANnDwn7y6WhMat12SOG0gS1y2e20/ISFMWDypR+L0yYIxcHi1nEec1
r7nQIxmo/djJ5JPUxCvNXWHA9Xv68GLiJVaAh+eiG2KUZKYvS1FUT3lw9owxKltj
tAsLAi3mIqQwv1GFSHFW8dGbi/Z3Q6ZvOmnfgH6Cul7OquvO5l4FVe/WYDIhnE1D
/wO3FG1kFdYgf6W5hgyjIeHSqwlH7MasRSgOT+TUVEpUFG4icVJzlBmDMTCBjS6z
Amyxhuc15z5RFuw8NULpPNb2w6ihX45EB6wRs5b7xAzHjF11L2lvYOmdXRxD+krC
FVceOlyFCAIFK5/UoJf+2wFxlOiVB4hbtyaXxNclvUf/FiE89Aq9bs/LXJaZ4i4A
kDqNeiqr5OX4qipA6V3iSo4SD/VIQr5uHAKXb4T7sWUW0ZwdPuMjQSDDKihogrBG
561F7pQzDNv7Gl8KAjf1ZJ7GzqOwtb/Ikn8uoAo2YPoZlJdPFkU+UTEEUe3UrNAv
jKR2KYJZ47NrdNxdlFDYVTJNjgeYEm+WGCctqrJBSkwinoQRFuwErSx7bmXiyDxM
zMyaP0mRLSmq+/Qj0W0hgsgz20WHzjqtDY0zChbIFioDrnLSUnIBPEAp4P+8vmh2
+bNr8OO0dFJJ9ayfllGugEbxpBYLsetsenNFeyE0ovTYrzyO08Kt5pGvAJ0kSUFh
dDjk6NLMclj6g9xcXIKS7PE+XfOaz63Uj8tlu8LKfybr5B3bsdsYIs+SeDwjJEtr
boHn+M5vdzm4fK/bhxnVI8tOBHYmxTJDC88yE3b5u14eL9UfzmKTDB5+NCz3vV9Z
RLzdqzfKoY1oz5CiZYs9LnbnMJywBSRVVheT8CjL1odj20YTVsTeAlDUaFG+L+dV
D3t3yTEoUfh3LL38SiS9SfPzweFYxats8Wsiag9B5FFg2KsGEuMd3bXAN9H2icPd
roijsLjQr28INhL2mFDHqCI/kRDH2cLa4PkUtmjrz9cLVwvrZguU/mAxkX30j9yM
OIfCBoHqYrNOs5rLOKmtWuzhIL+5v3kZdL9B9ZlyoetAzwuQFEMfkrKTh49yO3wH
AZ+HarWG6aEg1Uf9p/aa7BeQAovRJpzN0LaRTbExBtxKRbEOwpGsenOo5JEJqrTP
fAIQZunTGx8gvS0KDz/2AKdnFx8z7k/73BsbDoA3qJKnPshGvoGix93VDioEewEb
uNFn+L7CYP7UksY+4NFLzusTXb6226KjihjVKR/VqQop//zTcmNQGzeVHwsexfvs
cRFfy3bigThxdIeGbbZEMdwgCYPYuYNusna8NHc9gnnB0lUsP1zeTbu6OfZQcRbX
s/LUhaq6kKxIUK6caCqTKAgPz5TpAlSoxdRXiEhFMyUYcKwzBhwCy+I+rl0rVbmP
IwZgMABbh68qGGQCIh7ZMYZNZGR2TvsD4SlGSru4NcN0R4l9kbeMDDOpg0mIrbnR
MiiWbW4sljVjfoGfLEnRcW7c27w4U+ZDE9ebzBnx8HOYmYJW7K604m36w8Vrn4MG
arsRNXM66BRwCRB6PUj0d5GDTjS5fKlDZ7OYpc8ILWWvOLC8y/p6GazI5Ch1fQ8M
05Kh2fP95pzPFcn3j+pvTjL0Yf+RbvPCSF5zy/IG9tgOV60DebDjsvN131t3cKb8
lwe38Y2Kn5ZNVyJpydJk2I5W1Szn7uW6zYe+E4IAeAGB0uhJhzvnIa4LuDfLm2F2
vguslIc/TAMmy0mDL+C4KOtcWRRhZze6vXg6xn+zDpKsnz+kS53mwQ+OTadHUYSh
v+4+7AxLNhxfT+DtijNMwFKMUw9YTNLldjYECNe4B9SWhlrZLvgHCP5kJobvIKL9
Az5SWvjZvzdSMYMxv1IKTZ9ZoDx0/0ZJhIt6s9Wn5uZ/Bzr+L9MnIvuEp3DcUgLZ
pZ0rLGrYkQ/a5pLp32z4VPIqayHhuSkeojmVBjLzhFsb4zRzavf0lrVkNq/APSz/
IGQc9+znwDmNm/xBVzaTtTQyWl0XV+9M9pIfZ2bKE6grfmdX+ku4vQyBoae5EKTW
nSMiqn+oZ0OOSAbn/bC0zJGkozePNOfL8/uo3vqc/BmVsI5pC9UK/UID+6YrqK4f
DiYNbwJ+siKdg/lQu7mHH5D3wVH0P4GxLHL30qNkzGB3N4Hi6GUmFsIvPhLroWEd
qj4vu9/bKp3shDr9hPv2eFGsM2ieWqPJhE7TQvXhlx33XTEHi3Ul86+vNYSPH+AG
32JnoZFADvk/IpI4cUYcDobX/KltIag6cPmjv6DGDmAiUkzfhXjn72lzb1KDzK2c
v6noqhjkzEjULvBgJ+BS2ZKDLOUMTL/BOE/8kRG08nmROZustFENS91GCfxOwW0u
V30yngE/F6DUP1svulQQEbu9byN1B5NDRSH/+XB2WzPe2suVSSw42QqqRrH/0i8p
0V9i+08Pq678n3yaJvsJ3/bWXjUMB5v/nJRsSPKPkaB7eiqMKz+ud0iuj3lB+3vH
OpjyM7zIaiMsFaZU27gvZtwsm6PigFa+sOz/EMv4zhkjRmvEN20+FdxBW0SXvdkC
pTqvnzoh71PrFClvJsWepBCiBEqU7A2+1KrP+/+4nsI+AaCVpl14kqkJotMUTf1P
Lj4ta9uqrJbmXgolT9bJE+Shg7puLOZUXEftmX+wcZW72aHtlXaxl/l2ZrzZUHH3
+9eXeBBHok5gxajVRHDHHNgD5cR/bGarjRMM4iCq1yxTd8s82GOvsZ7GFDGEbX5e
afktcYLn66YJZAX4t5c9jgItrhqGPS3oU9goXdcmwuO6c3FfK1TKibQKAWaRB/lY
JfPLX62uGrIRTWdKbRH4BHiO/2nW12TdzT6a/0Z19W31P00VzI85QTjS1Q5x1hz3
zR4WJhkNnrN5wdlFFULOA0bisORqp0ywpeC/8x/vEIKA1tt1aYr6TZ9/rOTY4QKq
VsSkl+YJOKnBXhAXyZz9yPuLfbyTanMw19Gac5BWEQNyqV4qEQLZMgckI+Ccj4w6
yoACluIoYQYIijlYxTWP7hMygDf5VyvKkf507H6y9OgIkb4gKl6YGZzth3pHei2a
StKedgrjcG4yoy3ihwHrxrrSZ0wuymkol+YdzU2ODY5VKfPnGRrx4JkUf9Wenbof
LY01V7oeTXPL7shC69S50ZRXA5AFo1U3NTtfNGW7zraTa3qZq8/rKKKnvIrqg9vt
qDOzjHVBBfMJ0eNLonJ8zFcVPni6fCdt2VKE+DpueWF1jHriDsuJGwU8Tbf2jg8H
mL2C5/1a44MEMvkkafG1r47MBE8L3X8VW+oZSsfLAQTBUgqzyX45u7NTpAZFVgye
p1yFFivEG2y1ZTxNcOMqCI9t6hmAn6N4CXzgTfzxFuwyht3qcO1ey67ZBLKD5kEd
ibf7PQjXRp7MxJzqZssD5iFmJZErPR2oFvfs+P3dkJaKvgfg/o92rAggQKmFdl49
9SRsp4P9/uNTs1y5sJ+RMiig7qE1WJkS8mAhOg2uHx7HVfSAH2xZx63SnTPiWi5G
LiSYSj7tuu/HoD+0EJp2pm3tNbD71lAv9MHLExkqZby2an3rO9d0rpLx6UqY7qgp
YCFgPSwpmi9YUjtcZSPgyF38rdxsqgTWkhfKkOEgOqTAgwDQd27vbbw4EtC+kXhH
jeGkbvWHiCttwLB9UgdyuvPK4dLVHKnPpwDy+qFGSucjFa34hkwPKFfRCBKAUhnr
wtDKZByyB9d5TwiGVXZE553ubFc/I536UokoUkt0WIUCl6PFJ9Rfs8ajyOc7bUQ/
cee7OC48GXPNzjYuAxHAlJKId8stvBPvlp8oIssou9mtE7PJ0HFIyuUiyvTSDm+P
1exxWL4Nv4ew7DauppAgUkL/bsyQD2yEJl8UT1uqG/+6MgqPlnInJGPjyxDKcvSY
nt6yC3Q56hm126wQ86+0qwoMzyjEXl17yQCoRIv6h+tso+Uow2EORMOZ1kKISwWe
/2y7X62NShf7j+X01kK6YJrsEljmt6VhM4w03L2TUHfUu9rnsvaJqKFGWu3g+g7x
5OMi0PA3hA46Be+sFWqqJMuG19PFPxvH73sRWehKvuBL/2kC5sGOUhSylV+UmzWJ
wEqsu0BRf43ECGYsphmlAbBM0koA03zQAPa66ZQJ6FQwZsqWtp829W4gUUDtu+Vd
8rtq2jOXV+njp7GYozRyZNpxmAoQmTL8Wt/S1/YqgroHEj756imOdSoFKidTYCTj
zAzSPGri6vYmpHaunQGQC+LG0WDNCouGM0wkIRdLBgLtXdWzzuoiRlD5CBnm+HTi
XwWvl36KdX7lQ55UNcQImB4zvbZnB3pqxL5Zb5Z1XZDILBfoTlqA9oYeLSLxDljr
OLDtZRKyZO1WuhbeIIlFQVsggz2ShS13mpkw3onsMBUuR2cOi3S8BxhS2qwDOe9j
/EWCeFhaSjif6EcOe28t242vusc1w+yW/uHt0+e9KREi2+0hWIfGZ92VceS+SNAg
g98lUJ1+PJFirsVX+rNFxTJIdHvYbBt9UkZCSGokiB7tjJwa+N4To/PkpSz2vtW3
1Q0OEJVIe4rkCRorapvRPxtTFL6zwYLPRB6XK7D4143tzSTiDdXmJ9qho0h8hs2m
88UnH8/A/tKCvDK8pmZS+yuX03HVL0ym0WblTEtmqtYafUhj1e6eNv9ZwAoBYE2I
eWN66zA8KHIKeDhxTicHM1+/fNNxrPWQVw1hqoGFfWIqu7Cck+AKujoJHnJYMERF
szp+wcXeb0ssNNNvWi22QeAIsk0ZF9XrQJGn0fmVk45ocNaK8DzAtBYZ/g21sBZZ
ruXfrg993idvN9472pZgxBnSp2HBwEWYQOHzidzSr7cjKvCBg6RpcImo2w9Ot/yk
uik2GpnMojt6N/o7/Gf3tuH5sIYSrzb+7oEyv1gCpXAa5R3F72JYTLlPVxAMpBAg
GNaBbpG2XrHbH+eTYBQ3GaZ8WFFKh+5TC7SYf2b/tNE=
`protect END_PROTECTED
