`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtKGYzERKgZNijak50WRS6TinicMr2tXEiRPdzSthVUYXlxU/raLxtRs+JpdY8Qy
qsIgDHptxoIvrt02PkZ4EVr58jQdE6faFHCUc5MdObkN9u27Teq+rRf7UzybfD9a
LPQS5vQMfSi4Z5Vsa5TRc39YwXhwsrCA4mji6XgoOkmNddyjaSH3yNCNcjrlF9el
TH2Gb+DjEl3Tll7xsi5yzw/mtRzWjCADijGgvGEgLGG5/ItiIUFS5j7iPp02xV2z
4l5tIojZJoNiaeX5GYi62J9qEIMwhYC3nS3RTu3zOrTx6P3TicCYN4rlT2A5UKub
EhA0zEMz+WnN4hpnUTYYYlHj4cBz6cNEQ6a55aUMyJvuSHKkkRmKZaGxZE93du4l
Y4FNeEoDwl1NoMj3J0ZN5bJTpnP6mgMZICqTDgVSPFIuc7ugRVPs92dLKHUoYsl4
MArsn9/BzcnqsYyRv+n3SayEO/ZB+Z/qdBjWkQjSot34yNwfdIHuq5Q5qpGjMA5J
eyAuM3mg9GjFSgB6g0go7/FOSOi3rQGDwordoYr6ep1Vil55zfJ2fxyAl0jsSBJH
dJiZLzX5b7ORZnPiJafaJLcHL8dxIa+KqRyzv45yUCh4aQytZOWGDL+CPK6IZt97
LZ/u7rQb2ACPALc073wLi7w0TddRXXiAcjJPYq0tsP0TXqrDfReaqk8zaSCNvcSn
xT0yFwY/VJD9B9mGqDBK2RqI5kf/E0M+AhC2iSSqavqZdXQWIy4a7/H+GKwDfJmC
kEhEUdc0VNqum+ZGSFHNK2yeB2TSq2l0JT2f/ot91yIepGxxirEgg6p7qA/ZM7Pn
aovQq66R6fqULPOcH2vkyFxqotzv2homiqmSPmvJQbHHrzyOTcZX2D6ht+0WeZbS
Fsx1t1Zy4fmSnpDoshioNulL/2qwZ3YoL5I8+3EoM/udWiN/0mEbZoHcOhKImoNg
RSTG8/EmZNm+k2fOyz431VpAK+zxo7KP4CGOVxnEXAcdVYcrpnH1AN0/8vQqAORC
piMdD1mXMg8I92Z08MAlQcU9pdyabhdVqaJznjkR40nzHAyAlT+xSGSq5jCf6A/7
q2W2VXvfkH0+ZgVm8BMk1M+6MvIw4SJLLboOGwRkyHwLjMOUHeyzwa6uhMgWaETb
rbFGAUhCQP4fQESyDD0l93TeaB6YUYoh9q+tepFPTG9woaX45p1PuOW3KsXfPHA1
O3eiZVBGsO56dKxrlHGUKGVGL+Ix8ckfhftFuLaNO6qNpzQzp4KCF3b6VGUngrXi
mT2TcijC+h7GBdBi4VaY+y8DCHuC8yzqcj6S9gn7ivVmcKvCQ92JN4OdzeGtd8aZ
k4rv3aDu2IAe8/I7bGEEh/gtEcO76u8tgOt2QUcns8oRTk2aUn0fbvLZA57EGcyE
M68SqNjMGDTk26NfkmvG6zHXcLeGyFT5hDc/YOh9x+9LsrKlORMFNLUyW9jFJrK6
d0NVgcJ9n4ndEDLdy6++DIoxqOwan2y81hjF508Tfgy5/msev6JoeJYeyB1ol/a1
0xIiQDwsKVt24L84nvtMPLEZaBIqKWib5QkiUayPxdoQBCY1JGTAgP3bp1i58lKa
J1+iPrXQ5ohxaIT4fQDd1di/31klbXyIvMvL9G4mEQ7ea6zfhqZ2xA38lZrTTCYi
TdoUfNiRnqO1yVsgJyRJGCIZnLh6vC6NmmGhNTSW2Bs0+k/aqaE0sxdV67TQ1yxU
RmWlU9UBbCZoExjYcTEofA==
`protect END_PROTECTED
