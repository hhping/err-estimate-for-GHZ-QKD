`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3jaAWKwAiP+TOsYDavm58m10dGM7LfVyIB4/x9u4MWJHBLoitfDvExa98S1io23
fbULk1swuazJr70LT9cUOkS3iiAEb+LAVMpiFgRouQAOi1jwx7WGWYxcqcj+3dvt
WCie9rw+VK8P5F9O3tjS2FKgC3TDJ8FrKs+4bAaFCdHyPohz2ZAkHFD/lXeKMHqh
uMMt2LOS1j1F66QRJilZlcSIit5ezE1yIXeyWOrvkQ7GLvcdnejNDSBoY3jpyNi1
TR2OvN0lqaxG1G2MUgzTH0i93gjGTMLjJIMPJCIhaNk6La8wuadeevqbArE0Q/2G
MDgeKcB0NPTKRwjKVdfgfOGJX3RSNEUuLHwggti/qIQeUUe7fdhqKlJnq7XVtLuQ
DGZ67W75fY6jtzQ+q/xoZ6MN7uy/DOPipkmybLUq+ubi6bmwstXeYKG5T/+HGisA
Orn6dDGBZV5k0v+E5eKhSVimfyW7mG79HD7s5cLUhI3XcJFyM2OuenLu2JRZhH4L
jn/Y334bjYilz13/ITyim+oLRrlJ3GFHLExr3Y9AhJ3/psce4k/t1peUwVlb7kpK
40VOu62NfKqqNpIntNki4C/+3Zak2oyt0jS5nDyzVREaysUsnB6Ax4cJLGrV/3XO
ZpZjOSr29b12PnRoYVfdDpSrDZwHAAfAhEKcxvF37qO1spMfseI2r7Z1bJzC5EA5
w5qnA5IJ+U0diuko0v4UYWBPtbmMlRHs1pp7Re9v8017akvFvDJ4ZfJOogIkUaBY
bySCTsR5LdY+YLy3lBi390ms+iNIJr5kE+PlRPe4ev/TZAFOSxKYvjymEbL0Q7io
8tldrKL0tDvRJw4uZEhTNt4FkIMwS161yvPYfD6rKl3Q0Bl7qBBKoegSZAsk+XlI
Sku67OxI1D7UNqrdz/NkkiuGIHauXENtmweWh5SjldPHY1jithqygn+zWaO+dGTv
TfNPgWJjJCVlze7WCxGRZk8WoHueAFQNkWP9Kxi+YQeFY0Cmd4R6t8ZSfwOnhZYQ
9ai+SJLdJwKEFtiS4mUiYMAMi+9NxMZCMX6eavuQrc32TBgac2OxVlVs5FLivWlO
ljZY5PG5gouT9BNNIj0Aa1IbUDERkl6HHZhr3RIcGSEivkVCf2zooBDTQJO6qD44
rbevOVH/D7nYoWlV5uSyiVGEbTzTLVT2Cm/sONEwn+CZWXCgsXqmMY9Ou2wv5/Ar
dmKM2ENu3lOm7REZZGBNaejskEC604Jd0GEhtrcIKlMjF9RADPxRSwoJ8tI1A2RE
FTZR/lZQaeL3N28N8ZHiE5Q+ds88lckrC1EqI9CJOphtxVItHIxQ158TYb0cYEmA
JUCnzufvLUeP/9t2akUDxMiT1Zl8+2VIq06DD/o9Abr7gWDI52hnmW51VDcwU9oz
em3iSY1A2IXWE4Sg+drNE/RFEFzp5hHs3B38WFqPaBfBHmAsresOYksc7m/cP4th
xbFSkhbrpztXsTQoaDdu5RYiGZjd5uepTieJJU3/879KWrIi8ja8dkPIobBNEG5R
eFtUhVaLLuXypTp5aq0Ac7RRHjw2FEHAmZd9XNKqTJdmHCBE/iKPto8KSpZE+gaO
mfp+YScM6WoRu2ofvZCxIdI0DkcQkMJEITYxmpfIpGxew6BYKqmjvR96gIQM/GeV
iMDGpvnI1pDouQW19kbDZzGPMSxF51PIXhToY0+AJheZ3vD/G2n34oT8JUqnMXdg
2LamFtc02OWYIlbPngzJg68/c+7G8b9bqb1J+d3XpIECwtzQfOsDiBsFte44dBTB
5FcsUn/KErbRSbCnF2Lq1LsWt+6R6daweLQjSVf5tYY0uphIEUuH2niuJEurl/8g
mwC1pGzn7SB9SfbHR+yiTKXuQvVUgAETz0dLgZ8iQ5Hcb6eg0CtAjWnDVhstTk1B
W7l/WD+2oS2g41O27kw9P0MHcXKsvyrxI2d7YvQqhuPEfLdAuPqxg7Wbd1Gx2j48
dg2Q9gWUr/w7zpJnoysQmyhQfiyNqHB21pNpRDPXOCdrjdh3xU4WcfTF2xZsiB5k
ZR6y2KHpKx2TAUQ789PYclI4vpcnKDngn5B9oK2IgXERBf00Tcfj9ldxudsvd8LG
C5Kn23l0+v8ciKrkhCo9uFCMtMtvWv9nNpAEX+eUSxgWRlNeAQfgxAWhs9/C3Yw3
qmTDwiqCGIbIJsRdGC03i12njsxJbLhPu3lVPJv6B2LaR2jn4ofE/HDNhiMiLvMF
U/AZLSfRTBjCQvtKRUBAFq4T3kasdrF/NrT1U1ovPhIfVqI4KMXLLe9rPpApJwAo
oqi7PdaUT5Ancj8wsOflgZDh7I7Rp2XdnbXzxv9QZw8VniasmPMBNKgKS0fysE9b
/K/zZzYcCkZwsxvLQE87oN1o3kD+E6PoK3Sb1uh9ZWR/OknvDR6LjK2qX/LgRDE/
N7m9QzlfMRKQjFxJ2HgtgDEPljNFBDuvRFlu5ksIIcDv7ZZ3ohZdLeKcQ/KHwqEB
uHqlCB3CpndPZhu941lbkz8Irk0jOAhrBcKliRoWnFnBKZ7LJVEhmVgz661a26CA
NO6Rgt+BbxKmR3vSu20B841EHY7stKvvpSLYvq8qhpWbW5bQurg8VdQRS/G/nXbH
`protect END_PROTECTED
