`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0uVpS3JjzIlgzRuw+gnCMzjfGXniceGQFbJj8hxRqBU1ZPTGNdpr0CG86z4QcEA
Hf8YCjZOdZ91H8mQpd1HNRTFTi4wZy0Ia/Iovmc3M/UKM/2oXNME/UBUC++wIUh+
niPlNw94z6TnQRmTOO3CdgtJk2eP3l26zKZ4P1ipQJHP29bYAeTKcH8AB8LF+SmE
oO5kXMFagBs3e+xVrDDgBQt652hh619d4kpVN4qzj52a/iFNWqjUUlDnj8sa4fV3
4gh4LEaqu/89JuIOUPA3s8yyTDcvjfyvUuMVRAs6KpX6Wic1NTgROuZkNxOVnneR
kwUOOorcPpkgg745LkeA45WSGLh7jNiHXyxQnQm9WfYkUhezmh05vRKvHbu0srkn
/1dG1M/GWcYExkKFtyzU3uMrRVU1hOQY6xRdTO7rK+4MC3NXZ/IOsY9zZo6xpaYH
i0rwb+6HLc3mK6qncoUnAIfq9ebXwnvji4nKyAe9n6WSiESTEimkq2MGxmQJXmyO
wgDiNocGEJjNCnPg8SZ/gm64GNfbPV5eWCXVSD/dkfrp3OaFPwV3r2H84LiMoU/C
6TrXhSoKAJaLHne9kEHLRl8il4ch1pQWdHM4vRPfUKPSQHBtxdGayTFWa91AzA1N
av8b9yu9YExMgD/3/zWoixb6t2jp0ojJg9RnVgDqIt9lMSv85e3Gknjlt8PTEIDZ
PyRY9XFwfdhtTDkisAYASRtCElw8/UQVUwqDDGjrBuTkvzGb2EtC880K8+dxRdow
0FtLmsMUTpF2PkF8TRArsensRUZgmtx50f4w5ccL3Jjq3feenoA40u3Ugx4JiEcv
0MZKpmsKjIvAhz9XqgNnquLmcsf1sOgYMRllH02mPJA+zc/SxYlzMRECht1irUA2
A+mnncHUrtqi2GKAYL+camHbN8QlJWy70PDUWHQwDDeNeEDc/gsPOBRcLfvRL3ei
r/AEt5xJ9SZpt1C8edzsDeIYHSth63c3ai1RUVNOi6ZDs2dXbQAmOtw7joxJQGEG
4n+/oxuvzuLgm8v0Rlfpb+PwnZQ0nuEd4SWT9yx6ol45teHFZ6WwglOsvbJxYtRG
aNS02aFlkM1XP14VImKhUwz1IkrR5bjp49ADGaJAf0ZDMWh7tALHSa5Q07zPQc5e
dxlX55cqRmWRjvQOmjaol2ygNCzddnkcCGPJNlXkMrZNg5XGnlQDbUB+CRhlu3XV
ybdeZ0Z6Fj/o116S9/n5SH5znpDOghBh55z4RGMA4oLChEMG57qHDyImFr/EDY8s
`protect END_PROTECTED
