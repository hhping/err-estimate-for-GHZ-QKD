`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAxPGmHn1o2S4FjbSQOnq73VdhDaz+xKN4mIcZLGcyx7LEf0R9CF1IVMoD4ZSWtP
I/aMwceYOwvyvpPqSex5UB2NrNpD+2gL+LD5zDX6lEbTJcbLPFdVsbPrdeEQ3ii9
lf3lqt2tgfj58R3YQGVEJbzck1J0DCoI4JC6LcrJzYM6VYUEWp4WlYFChlDn+zyl
Ta0fWnPWQzRA00/rDTX6clTVru9AA4XrF6Gwc5OEhNAdvOq6qUpOJmDoyYO7FaY7
DLfZ/vU8/LTQcYs9meWgGtrIyceQ7gKfQqojfjasMGiLVVxRasATzevYlDIEXTL6
2Iup9lxJgLBviAp/LDJgtvHjSBu9bLhV4oyTjpzc4RaOKc3MZ3jEx245NBN1QpHT
18yaDp7z6xU/FNfd5P7LO5L9DXNet/RHYm3HZh1MwyuOOhat6q1UKITTeISkfGL9
ja3n8p7MUnYJFmieHGOuFdq8PkmzB9x9zrTkaiQ5uH+ViGpkFXL4G7enj7tDWTB+
E1leidCNd8uY5ut2Nz5znkRwvdiH48Z9oGxvTG1z6Xnkd5wdEdPRrqpznb4QNkjV
IT+VqwvRorhhwcbCes4/j8Qvlz8lED6o9vLKJNh/2rp/q5hPhxuvAmqCZ8xWc+O6
D9VW6Sr/rB6/e933gy8C6Br6AUe4bf/Wuxjus1iYlVI0D6WpwvpMk9Xb2fenUMW3
WlvsqqIwKf+iZD5twfUOTa2MEHkA1MtNoDP71u5YVnxYKqd8YfHtpQQmaQmI1paA
+AqJXIyaqavQrESTr/rVO5SRSg11l2ZhzPZWZVYE7GT5ZH1g9eQwnRURzdteDflo
7Es+LMea2alftNyo1q4T8xhoCmHrR3tWGu4TLceGL8DTpMT1v4dxyU0gEZPPiAD7
G7SGCxSiAvjAWyJ84iyG3n7YGJa7rK/kGVPrnrMwKHin5Q8qFQ5Jw5fUo1QZLfbu
u8ttmlpmpX2Kksb/wDspfcCsiFrWf7Y38YjzEw5h402x4e9rT6a7jgdOv0ivriwg
`protect END_PROTECTED
