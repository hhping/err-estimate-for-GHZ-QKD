`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
96ksk9KVrwUbTIpQFjwEFDx4l7VAPrEHuit+eGWM9lwYXPrG/+GGiQKLz1slFQTs
z3Nw6e7ZHfcbSmuQYkLWEdjBex/8fdmm3IVAEbet6qV54S3ZcuX4RBNuAEXdrkDe
emTNuCgcQaX/qc1W7CID6p1EPViR47jeEng6iE7U+ktVyPXpf0GeqKXj+emvvgds
TkaLCTnAaEo/PUdvdNC16PjBqr2aflB0WTpgSuL5ZJHYMXuhXvLqCpAFhHb7+VPr
V7S9TYgHVfnJARO7qpZJc00Z8hHk4Y+Qac9G3HjSgco/hUWYkjVZDGqQUKPK+80C
67WaHxzeA3NJr8GH6FM/mgos30yJ/lmxqvZuRJ3fxmJAroj5rDMQH94LQS8e3HIR
N5WwWmG8ETagEt8QgNzGqRtFsae+jl83pGTHzXz9RpBdu3j+KXM0E0lzqM/2vFnO
dZLQDOGFRb5Co9zKlkoeYqYGW8N3arizxONG4kgTI/DkL731FXuBxnuo2W26ed+/
HuOS7EZvpxSeSd/l/IxBmtyVIK6YwKNMl/zh8yvMbIoYqh/DnBNYPg0YKF1AJIQl
kRLuDwFGehSKo1nplStkDDR77KD0lxTNG5/ggOzTQdyNQqvQQ2WvGZes4aT3WeRL
Cq5ou+4p3w9WhPgoBV8A9Z/HhRTOWLuHtbJhIXYl7sOtzjBP0mEXU7Yas45Xq9LO
wL3m2/fTd2nSxilDhcE8GA/sg0T52QFt0ZQRL+yLzQtJxBVpLetBOxl3HJ8yZqyX
q9eWRbzPA7U+Jw8/+Y2ZXChoDzd29Bfoa1hrWdds4yCTQV/iIE1D6oeLMVbIRYz4
nV62YAcpzb5YjZNx2+bdgwDiBfqa3o0nu0HcTN1nJ++MTdhdid3qHL6CyHBk+X/a
t9W9Zr79dfi+qvaDuPbqPxJW6n9KArvwrnV8XbWKsBnt/YMrNLWTifiZ6A7iYuxz
+L88V3X3pLGNaQ0qOM0zrO0XU31cz1jm28+txmc7yJVtP9CNtZ0+Xvc+pmc8Az3Q
Pl52OOrTXpG7IW01eMk36rkr/wERfLElKwbXC6jz/3tDCAwuD1JYBhPeJwJHrujd
6jRYUO7/F6uhHzY2TTkGPk9ZCwL+K717hUv1s6q7H+NaQNYtYmY+/kfd6eUiP3Yx
DYE1fJgg8Wx8GvrbFLSwKUhVVZokoTN005mMnLOPYTqro/VspnxDfRWa6JRIo/5x
Gk/qxSmX23oeXzvVCiulj+IdFPLOG0fHTn9woir1Ymkxz2doEirLZIF6E7tM57J0
Hfrk+u7AnOZY8pfOKRlYS5EWtJ/B8iwmtO+bTPGglEe57nCz1aCpFMPsvc3fZydP
y8MigoWSBxxaJJk3nC2u6WkvstUMpBY6RQHOmBpHHYbPO8h9AK6fnTcwVzo35xfK
`protect END_PROTECTED
