`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PF5ag5KRTuhbaHw6q85v2x43R56b/KLm/o071pIEiOJBK3JzazHh8gVqo8jTbcII
VmlZwz8/a1qA6GrXj23jFtEITu9WLPoEG68U0LlxlpOs36uYjt94bGEqBnIkgERu
v7K5xuq05IGhf5W1CykV9+1h9XLIcxMOExYQXTufPO1nVHE9npfZH4Bum5VG6iRx
nGcwogWwLUWUUZil0LLNPP04SdMJtXf0Z0zhjvYNGm+Iq2WeVp+2eK59jF+f1tl+
cs2l6Q0wLYQa/C1RBtdZJLBuE4IS8GR2IfoRv8swPAvw8QEnrM7kDFPBv9UXWCVn
1xWkytmmsBoyH5+VpVvF+TZE1lra60kbGtUoNmcrKmU47jQlchs97hohdkGBZivK
oHbOLMjQgHdleZ1wMPV77jjDvdAS1ptucsCooviZaOxMSE3hekkK9gQu80x/DqO3
csPbRMIYVnq6OW5QKA+7VOwYv5OW1F4TvamI9mTsreWE0FPfjvseR96RtVxsWGeT
bIlhSeVJujuY+WyAXluQDShzCTlaQ1gVD1v+qvF0HIJMa5vFiy2wdScYCS5ovXEM
eh80LmG7apspW2mIexmSfdF/37IkIpYgHpZzm5ZqxTeuS407VjGdN1IymhbViWRR
EF20Ll0g94PieyxmvyyoQm7jlh0p7ATp3CbsVb7bhZAq7EGYHcQ9blDcmp9lUIe+
b5K32vUXuloR9w5o3pOiFU6LbOTPmdj0JWbPJNLJroKPTfsIm5/ShRkYYKwGKtR8
mrLAnpUJGMKtuvm2tNkiiQMy3LyGsBWPpoaIFfDcJ4A=
`protect END_PROTECTED
