`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymbHUK/5ijoNTvISsQCR5ApXOjJXCWoCawl6AQOM3+Su3jBJR1dizzTHl2iOhToN
ggKlZsyv2ajt0VDn0Y+IUut5E2EBHgEJkYEI51qcMBXn4mjPSYHE/yWChIMbvj5A
kChETOtjACFDJj/VcpjA0RBc2S9LyA/YfJuivCEImWp+EyszV4QzcpECqXfTdHz2
aRiKjkHZF/vjpvlnlmTe17NeBHOCPROtIcmTi1h63XioIUY4vdEx3GxF5mTndQXh
+2ItwI73qQs9Cv98StubTPeKRLFGW7Y/z3e++e1nnZ/0uKbAIDQ3QwH0Y0+yZ37s
UwjhmztV3eO8FOjzqANs9AU9zao4PS48Ql7DgGk1341kcTbU4d9hdt37jI5I8nfC
MUe9ZCurebgVWRXsvNtSN9BxSOWyJvCVL8V4OLMP2FYPv9daxTY0pygc55M7+d3v
poekiTDyvnKkdxuWtg1I3T4+NYuwAaLYYPsN4Tnz56R7fqO/RtwILrG3uLMxTFd/
e2MR2tgBe74nGsCXWLupd+CpxIxoiYrNgph3VXycQG9TSziWWJAmyN3+gCsMjF+u
a807rUdtCe62TKzQdNbskeQPm46Qr3a36uaHT9FmpJMoDRpV4tpEKkMDSemRxUOL
4UtZ2GFj6dtTGJm0yywU+BrxJI06GYSaPHOYOy0FQwEvRJ0FiGe3Yu1YP3hTTGnf
cyKWKBzwZL+KctIPtSAs7XzjU828Fm0BR7VIbTFan7fk8UyHgtnE/0f65f5o+6Vu
zPfiQzX+xVnJ3KD0e220HzD+mElf59ulISzqRqSv1in0oVp7+1s9BJGe7Zp1EMZr
1H37xxI6mCx7tcDceV3CYAmIknsxhQuaceVE52noEJgsLzve9Ix3cCfg6858HamA
ydH6K+9/g0UOq/6RvqCieV+JZ0+QLktWOCtIqQfX8I15+FPNf8NpwSsR47WJ11Fp
K82Rz8e0zkfbzEPp8gQ4IA==
`protect END_PROTECTED
