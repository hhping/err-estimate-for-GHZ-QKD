`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cs3rx2Uv/7PGFhvdyJEOGnBcFIqn1pA+QpiElvkFgQFiXI0I30xajlF3ShWjK3Gh
ZdqJ5KqTku/kdbqHFJWe6Ro4UNsTm559PDH+Gu4bsKJN1X04l+E7Wl4Q07qzxh1P
IZxO8REnVTHz3BYVB+yBtZFvF9bmzXvIBR0wTJzYYMzvBNPt+vkzJZXS3FS8N285
1WID8IAzmdygDy/sogJKBjh2DvFUYiWALFZb6G+ufcQrMLiKuWWbi31hGXLSzs/K
S+36fFL3rQyzlly3OwUPrGUF3K4MKOA6snZU2PI1AbQucavSo8HYqnH3rV1aJ3tD
kDzqF19W60D09rm3x72zf79NqlqUOPfoA0A72Rde9/LS8q6u2qTVPUi8wy11qq0b
Hpj1cLUgiRxriHOCyBsbCCsa5FuYDlVy7anPJaqA2cBXPE+9+apGflys9n82VXs9
oqMsBK9vRQsI48k0KO4NRZMqiUkKl6WbvKF/Cq4IuQ8DOV4b7prXsCJW9Hi6qBYU
jZjXfrQVIHs8RhKkUS3qjMOyoU6/F3s/WZWjKLc9DCR57CVvbPxkkEqGFhDlU4j0
vi+KXhxRJ2HLOFcHGgPl+IEUfr2ZpIF7HIxUuTaYxuOqX2iieoGli0jrs2OEjGJl
Q0zUti6J5tXzCa/V0uNv3v7CHd8Xw8ApqVZABoAjBluCbZWwVumOH9tyVIHZQYGl
6ALQKmrqvw8U3EJyALe5ABv3yPmTnDomaaVeEvUZVz80mEqxlu9RVLoLldxqnqNR
V74qVqco2Fkjf7s8lT+6JCU4EUO8fsXNgvsLnUzbL6RUt6g9d2BL/M/vzs5IrWhM
K4GxQUBi6pUTXwSNUbAix878fOFbSmQ1/V8E1PrxR6wgORwBNjtTWzxMfTYVTgCr
b6lC2zCxbxX6WANKl8W3dqGQ4KREpDszlxcYmzs/YSGL18oFrzj4psPCc+rdsk+V
r5qhY7zQaQHmINjw8w3ubw==
`protect END_PROTECTED
