`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZltUB7+zXPaSpi3ZnC5Alx3eyC5T9mNthOxZriJn8Ky4HSDlQmW8B2BURPdPZKe
g+ht262RIbRxu3WG0dvhCkcodtDwg16c73nD0JocdCaFgqun1hpsAJLeTNO2CMwZ
3SuEOHOGpwWvq3+mZjN/BArRtP5Vmv0cFSWNEwdrobFQzBIB+HM9YuHSZLgBJ57p
1AAyMBV1IkwGHBvvWtoXyCdf48fYUpUEKoxBN39U8HQALntBIOCAWjFBdNsvgM4S
NUuumFQb8sZfZoPj3oU38rvrAL9WB0pHwfCQd2PnwJyYvuu+Mlv9GTmb9B4vKhqy
uvRtCdrEXYneYdO07hINZVHV54vtE+MtgwXt0vENtkWbxao4+mWrZvN9ZhOCqtw1
6hgyo8Qozxahi4hX9GMce7rVYCF/swJ0HITkUjvzfSuW4d8lsmivFOjdibNQIDUi
hAtqfBNDNp4mruATYiFOGHuEB8ETO8j+8Xy2fFiOvOmExC7x2GJAcbkkI0cUb43t
QaFojI4VCiXD654ykYEALVOk5VLpckRaN0YOih8Zrl/deOSM/e3nPsM7fpYYQx9f
4FOZDej7Lte6zHrVbYf9W3fn2Q4ynY/+Jwe++tJwaTRaYl0J+hyHNLFMQ3CvdzGo
x22TueuFpyPrUAPEnnLXK+t8XuZluv6BL6r1ogeefJlrB2OXHTXOgtf9u5bjYe/h
yjmWmjV9Y0WuYV7DpOLjzSlsxT1477NlQGykhaZo8tjFLIgLqj5McHsV00+14hIg
lxPKQ8oMrhoUpZTFFfsLV8tTQ408r8QzqLtfvgPiJRe5UvwUIjvYSkVYXua5GQ7a
L0PCbXK8v/79lTvLtbrX/dHCxPagyK384NICDOBn/4DbFhnBMjrD9JI6ZxYS1rQc
hGRG8e+2ihBaXkaYcI4WdcEeWJ086NuDVd0uo1zKx6VDMtG8qJ5XvmovPywqs4+Y
9ta2HmB3ueAnRttkNxk8fd4dagPNiWgnZbcEr79ls3++5JOXP9H3r4+OhTk8Pvcs
Ffz7GsnoJDN1noWmiiB3zzt1p3a3k/TLD3q8b9KAwCIrBlNYAojXewlbkvG9pftd
iO5iYRW8KvmT63gYoOrNCkMWxkoPGGq4yQJ9xgA5cDF9uRAt73+TEQ5B+UJRaXVg
tSSCp8AUrek5EqPW9E34J1DCOU6Xpd7L9kd4ICWu4nLMvSfif/z1y0+xnYbmaI0L
CeL4srNWR0pzMc3wUzyImjKfibVxAcZ7mumoDRz5OwyUxyfBMEtOHIMHah5S16Tz
k3P+KDsTK2ax7L7X+tTE9SffPnL3dqLFLZMKrAsOoFQFW9ZszMqnrRVJXy02uPpf
N95fDcbe5Z7Da0ljvd6lQx5rgO66cS96G+wNy6HZYVvsQvQtQOJT7b6OD6HpXsYR
yimtL8fYaRn1GTrRSlEuEJfsMESpqYZWPFUMU5mXV4Z9ZcQsgWog5ZjfSDACHnBq
/dLf3Teu3x4pV5uabSCqsJ8ctzDP4qoHFMs0Bk1fGYpZgHvyyZn6cgwffv3aCnMf
9pfJh7CfGImKNkNmJYENJ9L3qbSM0PDXy/4pbNKn5fachtl3EHzdf97glf7zqAgM
ODmHocv/KYs70fDqNDdBhSzcl6Dq9ReyEE6JYxUWZvBXjGrfnVN2GBzklNgVksTd
fdpUiK7BaPtfWrciKyQ5AugHhBGYtswbLjcUc1WjuZmW+uGWehd99DUzNQ676kk4
v4B5uIG0mGnZbyHjd/EtlkBQ7U4sa/fvscPl8j1c5ZbbSxmdmBqEL4VhIkMbJQwE
529kgHxG/mmhDaDkmEFC2Dz5+EGtXhJ6TpfLeugC3W9TF19kRVzYPC1Og9LuiFuN
WnNLicqzsLmVXV8LvrHGameBqpV6Zx4mFHzfJRF/AOc=
`protect END_PROTECTED
