`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U9jytzC9+nH6MTdmWjqZnV0zRo5YbwS28/ZrFs8TLd/9dv6IEob8qnMmo1nmFYLR
pUfbSl6uNr29TqqXBttEj2C9VzVDgDgaQGhHJB/CCwtRqBvcNO7os1+L6uFsWg+n
tvkjG+ARDJJKyvwz+zi4hTDquxsaBfUqXL2+dlITD4akcr8tjUu6cfCd56lbVDRf
gSqT483IUSy/JmgcsiP6m+1ph6eShwIVnFQvhcbZs2M3crTj3qOFgwujhTOzWKr9
XCj93L2YDQ2JUbODkwR+Pe2iZrkKt6agPPZxUvDADu68bYwF+eQZPPhRe5e9vpli
LGXTrbkvJp1KvAd0+/e80PwojBpA43HOvUUbecEjpsGMN/B/N9eLzdbFdFJXQbfZ
R5BU7/GvRCfaJlmJpvRtgAdcg+QsWVwhczm0DuavradHo9Zrz9pUsN1e43QcOu5h
7/jwZZHrKxB+NfcaZ/F3RTNG76xfzkyZVuFkXRBJQJqdoN2mGxi+HCsP1HmCIaS7
PuvXA+BVqfAWWpDcU1uPxjCoH+IjzEQ7UYDlAHkbP74XOEqodfBri8VCMj/vrfYU
vzq4n4/sGqrFUsJCHMNCUXWdVy/mAeuLuuXM0Ekh2G8OmYBpQl/rLaNZi2CoLLLa
/7/8gOmUmg9oenS2Sjdg+BaUeW4GfDP+aYN+wbvt+JoNf/75+0K6Lu8mb56ZFj9C
ntc6sh31ODVZWOxqa0NLT/7LrcMArm8rLHkHSU5JUweIUVVJnnnxmzZ7Ul0u24te
u7FSkwB8X4WHHxk4jo5rRfVzLjPyv555COdclZ7LWH3FMUk8fwBETzzZOR0/nilC
1G46RgRB5hN57ifY09CZFA/iGn8SdAiJlIt3HX/1zokdS5cJ4Ky8+MW0QHfMsA2x
XwJOC6FKeLC4erB1J0HQFpJRAcQcOw2ZX7PSDsrhjK11OyzgzA32lH4piCqu/9bN
ToUSDXrnIamZYmSll4CF0jzNV1goE4paa5pQDzw9fjVIoOtywaekeGSfRtaUvOCi
iMSLw+kFVuILac0FnNrpZe3KKfJfHpwAwRaHwKRSC+0yzc4o5ce3vA3UR94r/WDP
dc1TFpSvJbd45wfkxOkZ3YzxZgWcyP9MaSEA8wRnNLUaV9cHXeE1dnSDI+aop5GG
rBQ05kPjYDQ3C8eYdMnHHuDrEkUu4brD5PaARRjTiqzWNIsL04HlARSGXTZUiix+
j7j9n8eYyT1MbgVymDRs2eQjOlDhGoSdJ2Ybc056aBTrplgJArdIcOBxdxM/eh8Y
fRShGCyDhtrw3OVzH8RzKlF+YPVC4yfyh4TMvlvRQKdeL3eNCnV9OaB1xH2pVNg/
KLBUIFW60DfQugWJwxe8JcqNT2Mjs2oaS9y6wMlchdUENQvq00k6zMjnOn1sqtuj
+yvRXYvdNTvWCI1Aq8J8N7NW5mPI7CJxpEz6VQTx+ycpM0vkrxZ/ITNN76vecRZR
1YeDNXlpNe3SyDD4voECXbRsmHWqdlA6R64ngdBN1Sh9l6o19qXsUOT4zb95YOEj
lM/Y920RViZp7wpnrWNHXGaWDR8Mj5VVHpSsr3iK7smJO/3O7IRmHlqMVSjwmi3/
VdRvWeB73I0q0/CwmRDMRB4XP0aCT8NIBBLlfJsWn6ZPW6rhigtrLJyL/qiTNNPz
kHEM5GGAFAZ+Ff3CB2xQDdIyhDkjnOWukZLd8Enacu8lXfSXQ74F10o70pdQEz6e
cAhan0yXjETRSAmtLvG06VHLeFvvxVKtZti+7e80CO4UjNHuG5f+DEH+OJkBIl2S
lADUrBx8E3ov+ub+QCAwXjdok1lzvYlLYINIrKLwHI9zpx2YQTEzz00Qx9191j3Y
St46qUXqy5wWMcuJ21g4YbgYl9QhoRfBJAqnzetEV89Is2wyEZs/jwxxmHuyUh1S
C4Fqprnj3NqfapALLT1qSYRcyzvNUvxmyR7PSQ3o+f1K0shZJ2Kvui3CH85O1IyS
Tn1YpBCyOod5TTNL/4kIg0sewDbIbNwK7A/JGrVoVcVwlw7jsEZcxbCwFPPyBBgr
rU8rRWdHTJALs3YJuV+5s3jZZYppdQIkil8b1I2eJoMUJ0T5/OSPkZfld6MOuppq
HniatiE5bbVC2MfFntPkBBa2DBbYJXGTZY+p7DgToFYzaTMotb7Ox7WazqwuytWS
4hG7LAljJMDdnh44QgB3JAGD0Tu4mtWcrMukcQqIDl+RSj9VS67IZA9UQm6Kqp80
Htqq/DIM1i3a+MukEs4SW9NKAY7Ne4p9q+3E9cy4KnjkP+z391zLFUwz5rcxAQZ6
JQfeN8rF1xj1GXLAxsCa/F7mjOZDvD9T3VJ2BiRGsu+H8jhzmDLzSEI4b9LGqZY7
ML/Oeoo6x180j9z7TNfzg5p9+RmAXFnUZIxTJGJrWW7poMUliiUILbU2RSX+CLYO
fWS5ES56HKJYM292Lkkt7/DEO7j9QrlVR71sQtnALx/HAZbwUmmFhPMM3xNJfIEG
gR4iTzl+0NHuvgifNFGjT6MpS91a13kAARa/v8+TRz4vK6EafRj49g85ebHbYHHO
Kgm3dvC/B5PAhxVZI0PO2gx/WBMhYLW2CFsSE0Xxi6YrbZI/Pi3lGtFRfb2YfQXn
z5qM68DN0ENke62Ut2aBbmhduTGrWIwCvYN0wGqNJXo8lVJ84tsGGES1jFc+0KN/
ChrdM6dya09OVmidwPnOeC5vCH/QnoqXMa2iBRGh1Qpu2PAbBuIc26ke6qM1Ibhz
5q02oeq6WoON+JlN/yXMGH6fxfh5PkN9itcJazXGSRRoEUzKtYWt+VEfZ+2czZlr
T+50wj9eKUfhGIdVw/Ej/4WreY5TxaFULIAasP+ApZ4n5FzqgDrM/FlZCKql0haf
opgmHtzb8pn5SPQCcKTc6LOQwcrl304mf3/tpy8NmISJj+UiEXUNM+enUbnIr00m
XRCRBYUxGsgk7C8rGJz6T5MQLzSP6O1WJoBbPHpiA01tH/xN9dUbtQuQ8bW2RK24
L0PINf0i8RBf+SJWsGp5A8H6DaFxBbRRj3eulEx8uDGKboxEM4oaPSKuZuKNVe8m
vv0VlgJOY8rQwBW31/JcU7sB4afzjTLWTtuwfe7eKADh+UXc9jaNsI2JqcUCg+ZH
s5HQ3HWgUDZoRKVxXNN0pM9NgvH4y4vYtrzrNNnZAmzQGVCalrMPs5NUr2TfRq0X
Ag/Dn2OpqrJ9LuXJ8Q8M3FvXr8AXcd7JdP678KL14zY9vPDUP1TLD2jKgsKLMZgU
JmXSkR+RUPJrk+RKIRH357n/+9DpRsdscWNnQs+iw6zhJqV7n5DpDLvRU4xjMuPm
g06X74jdfHzj9pd9gMJWqXI7zTLSaGRR11nFvwxjIWGKyke/ly3KhC3brB6h2bHC
NuOt8aYPXMmVRZPaIz1AChNjrilxBcvDLvb4NQdUC2+yU2ev3tunOVosN896l0Yj
x+JxGYdcps1fh9nt7QHeZfYwlOLuB1jmw0Sk5AO20g77LhCIUmUHAfkxC/vZzmN1
PBq1bWfPz2KydaHX+WL9p+UlNWOKBOpYGU129WIaa5K4hzBXnjPLxDyqEi8L6B1Q
RIONiLx6a9hpeOeEJIxdqic4cG8C2XRg1t+NFvsL1drEw5W02/T3Pl/h3sr+RLg1
SqGOvj4CcoVlDpezz8fimg6yu8PGeM9Y4OmmfSueoSUP4cw7VRfWl3nBMni8/kVk
P0Wfa28iqTZi4gA/RwL1Y4KpmcCqVD+Suzn4Ux6k0BumFhJlmcdmsHvApJpTDG+P
HFAtsroy1pek/uZXuDD37McdV34FK3UUB9Tw4grRB4IW8IdmBYMJ8ZxH9jbrbDIB
0KojD9ibf46KPd9xwjauahRzXiIMNPyhAiftR+iOWRLNQ0YJiBXDkyWX4qfnBAAd
ka1pDtTzL4vIvqUOTu5hAgg9V0y+x4aj0h7IhiXUT19Au5Mm4scY3TiIuua+8wZh
AppuLzoSiucWbsKqNRQXtVE1Vf9ydSDBRby3dMzTvSCotw+L0yhc2S1VIqMUgAg9
/DyAVtsQk1siE60CyuBsncs3MIgldXhHKDecttK23ZciEoajUX+VBIAzfCiTc7TO
voKu3d16quNj+X3FQrw0UvWlcQGJSeRRfFJHZg0w+lBmLvHzDLyWIeyiherf9k0L
mv2YSjdX7pCqCUdTjf7SSactYC7N0igtgQl0QUW8AZo39uqzsDrCZnF+dMqpsIpk
UNj1SmS35A8F7mHIvd6HC+HZfBVMOfb8WcneE6UY+phlC9g1+6jZd36qD7vjHGww
Wo7nKfz/RCQp5glNCx2kqWYHMhgx5lO8AjdGOFl7LouEcro5CmlKhQuUTPXvhLaK
rWTwrp3F8eo1y36y/M1kP9oK18QwoJEA4KEQJkl/IDmAvbeLaaeBlUUA4CMGJ4ZV
2iUmtVgwQgsQxwQtBNdAcxkK3Lv3cClHQrYXeXRKKxJI1SJIwnOnzhP+ymsHHUSG
H4QYJJ1Q+VOxCAYxDb+rBQM/St/cHCLTtfBpAiRGwyzNCRAwzKu94MEXMZJstuLU
RwVC41VCXuoLM1HUh8WlWNiiZoiBOzDgmLCk+TVv2o95FBZw+b5kKnjgL+tVyxSE
ITZ7775tF+0AW/mIdgMGne+04+hIKVF1O61nvbrl9aV+aOwAo/62ruBLvtv0d5D9
zY5JGA4vRkHIveu/tOdqOriMgR7PwgBwcbjmOwstZ7r3+QUQ1/DpXI/a81YbUZtl
wgLXzsPahIapn4EsHYzGyWAB5FyB7G4FPw1x1WTet4uUG4elV7LttG0bK4vUKpuh
pNcEkx6v4FIUjCrmSo4XUxhSMkJz3tySA9J4/o6mqrs2F2nkAttsdmrR1PfUCcQh
MgAd8/PW1ox53hky4TEK5vuDHZ+AKEFWscDQCYNe10mkj8T60eG5RloP/QvCVlS5
t/0nNAVzRywf1drCBsYGdBx92IqstSyreEnOwSP7/3QqVVGhd1QFlMftBRZnx0+q
oWoJ07V+//aVzlHesmzThYIRNaGkI9bTxX/EuXnR05/ier1nmkkk5uZdA610ABIx
Pmx2E0ieGuTI21kuKuOj9zHHoDYRLno0Ytf018sf/IvygNFil2gRrti86rHF8yS5
nudASZ/CO8k9ASzN4VOP/FhPLxyhms3tTEu0qx6hlYcxrOGRh1GrL9Dki+uSXxdC
BhKmnEteOz145OiTwIbwY93Jg+zYAL2y4EWPH7iwYFBRz6cSzCxoBzHIGKXrEEXO
dBo+elsKWi2n116VLJbM+aUiNQHF4fuQOlzGOYtYtpXP/bzXjKjdziW/ZW+JYMVF
F8TMWgKK4vUNt7sl7UBNRCul3oXyucpTmKJ9dNj4R+ig+gbVbGqLumpPP9D/oYtC
RwM+8Q5p9+53cXpgl0zuPGLwxvxbi28UVwI5InAypJH1s81iASeqWo2Tfofrs598
DH9x99QWTvK2TG1i+3s2AhX6MVUQTowO8W+89QcKworedPObD7R7W5H8IkdGa1aK
eoBc+d8JXVvmturf4w3qMGJQmxt0FT/wm/UOcruZW9Ga8oHUvjNoWp0jHAmJfbcX
U7bI2H8OMoKpQ+I8235ME9YKd4uY4qDgzqxvPQ7lpfBYzF6/P6SuxRI9d+jmzKOY
9A7mb4abOwl1QNVeDKRvTK2k+W0LuhkTwLuev1kOVj1BT0AVe/X4JypkAvtxvM/P
R8Kmi3vsJR86WHOz3JSp94KcM7CTvLHvfOj8UZuX/ozMAXalRxQqZ7aEhWXKt6dK
o78//AAyymdbVZZuC2m2oGP+C3vr3gW5i0Zpx78hs/P6x+5k3+Yl93COgKQd2Wuf
4LmtLcuj80UsYbQJSeD9aRRLOLQrxm+jYdEAwwbojWsv2i8xxn2Dnh37uV/Hd/w/
dBQmnwcj4oiJfYlGguLlHa3vw2Am5RegZ9pB1I4D3cFnukonVrizvEnUt6EywCBB
B4saVgOvHAxtoZhz0P7WUpb1d7m+gRKCeuFOmRwOnRbQAuitkTDfb7otL9OPE99H
y4ohHzp3CNkC/m3tu8iQQjPWhAI1OZrQh7kEuryJ35HusEDUr0eYk8QIvhVmvxxJ
lPAOeWfb+tFYSBFf6Jce6Kp747JmjGTeyjbpbCa+5iAegRwE7mPZ5fSq1OeGq2+1
6dqtctOTIv51zGEsCbwh7fMkkVnbUA43i0/C/MSx/HEvAfhQiRkP5zYnwiSRnho6
SfHKgYpq242MrGQMrbK26Vvpq7Z17amXX0v9LJrl/cAzpzr4ILgKULDg/8tXHyuy
7BUxBQjjFQ1FkrxhpN33AixWUcUTFrWcq12Oy02iB44PWUlNcMjVezJ6/rxOB/48
1RBBeueg0X8ubCPGGv1EAj9jqivEPfM+k9aI/+3HLyPFgyGUmtZyauiPfYmH7TZE
ei0OFU28qbq7SkgwdcSXoE/TACSj64sMs21hCwOuE0ircHuRIt9LxzOqDijCsw3b
ZJ5puRs9Ziv+0cyQ/ZYkDrIsw75cqbgROtggq1gl/cUv9QwAnZehlDD8d0qDYZBm
I/iW2Y7D34ZjTTYoNwY94rRwTt3kRKHdZvbGVitcjV0lt+1sPous5gEesYet/Gk8
rekAwjdq5sYHqauBd4vlYxXl3+AEGRBUP4P9mJ6YCTRi7JPLeEdWCJ2f2vWSrCrM
oESf1dYrkipeCj7RHl/leyhi9H9KYMM7IQqN3c8S19G/2JXSP5/djHl5GpBZlUvK
1W8dz2VVAoIFoQPKIncaY67Skc/oaYvS4fChrgMhwTVpKa196OY4Tk0Mjx8MnZvh
TKJ64mB0HvbbYvHhFZovC/0u2SdjqnjH9j9Bfus+k7Eb9i9V74Nut4AzO96q6gVq
5DyH8kW2IHIq1z9PkwjR2qHSgGoe8KUAby39BhuzMOLGpPLUFSJNdbcLp/1FTLzK
+A4ZO1WCroxhxsR25/4+tGIifX33MhHguIzNwXc83E7IHvwMynln9B9bUoDYcVu7
pTBYCQojMcqW2877ZeghedE/O4/vzDSTM4i+iZ3N184m4qfggOv11tqI+kWb9KXh
+4S6pIK8cqeDeLcJWQ1SgI5AyGWDuufMre579V/BeUVtIKqYxmQg57Dm6LgcJNKD
0RJSeofL4s7oJkw6Ak9eQBzZzTFayU76+8xVFgkucTH3pSvXBVd5A70WVMKnlz8L
XSdhcwLweEgDIz6No40CkpSBgzamZSdfOmhDm2RY9M+3ZOznHqRWAnHh8IaXUnhZ
7gbF7Em/DAT0M08pQmhVzA4Uz5WveY3YclMfLRCrIreeuYW9nRVe1TzAJV5WocsR
jA8VqXr2K4BuZrBE8sh8o2BsC4dqSVUs2/kZkJP9slvhDhQ87C3YZ+yHeyvXNKa8
ifO10Bl2jagIuBFNgxmY21tqxPPLI/K+ruBtKoiE28MHrLWe4ihYcWaA1EWFL22a
7EtynoWrncMBUTEYwBHVz9NzUCTIihclzkUJNfbv9G8l56vlkaWso0PHUS2TuwzT
TAJgbpSZaMnL+mTUU5BaWxKZrKEkCGOxXCG76i2g/4z2ugbGYPkr644SwCPRgs44
QHxnqYWxqpDa8ELuzXNRVs0rN4K1xwUSC+A5tFIFJV0j59kWVAJXnjRvKNtfkTPA
c9WDoQnLsKOE4dOb5YC1PJ5aPgSLRSgPacyZhaJoDMAlVAoJ7JEOxAaVTRK9eLOQ
HbmIeeJogerl82m7V8N7INfT6Zio878TUO9ab3ppeD3p0XbZaKQ1TAPAYW7fc6OD
hWmk3Xwpusd2viNkgnHEV0AdTd/yW2OK4/f2oUfj8gzLrpH4+Hjio96CDJ3Y1Q5C
8jQQ8vrNfbATOFAvGpmSbwd/inY7SXwAEE3tnGk1/0XBMwW0G6BhdWbobysf6GHp
BPRjOfsTLROPWXKLtawpe3snIarBhKzcLkITkZMtkKsYVlcJRPpoFWyccJL7FxLX
7OwjWc1dDlvwSWj8knZpJYC14F+Izdz1PobI1ezYDi+t5lYwFsYhdzqjPfSMx5jf
Dqa0NVnVQ7Ell5/fPYAq0tA0E3znbipgr+zl3FmALlCCQbr7CWNdpgsMhiHmPTRm
rN17H5USuKIXfAa+oSBxe3TUiHsyp0riR+eLZkiwn5mYMH0Ndhj/4M90GTkbvN6y
ywV01XiyM0TnOp7qpCoomUBHfdMWjP5fgpQWyiAEF+Hd31+cp7FHoa3RoFJf4a3C
8WdwOhv7Kjsp6D2NGPXH2pbkWzFnu+ZyEBG4PJqMJrIoA6YZ1/ZIU2QOFSx7B6AF
z5OQWlUI3UH7yFlCHDw8+EyUOVqbPEzJnrtZ0odKoIKtRdnzDsLVGeznn0rJr9uh
tUy69myI3ju2Kutb2H2zt1fztanKn9DuHylA+YDjkbhNd4bH6E8PcQYRKez4lPNF
1EtxsdwvKFF3jUPRzY0hajz66bpSmM2FyxrT4z2HJ/P1TWkGL23e1EWhKDyZMIuW
PikgroM+LvXus/nTLrqvARmJhaKeHePABEmypuShX/4x4Mn1DRtwcPm4YPQAR+rc
NQSnw2u01nOxkVpotJ8bXaF4tbcoaEIjgzO44jQ5PObUZDSDl8s4P/cH0Jv83mKP
DLt03iaR5RrIbWNJg+vyViRDN/CqSxmxPjUcHwsQB6kWNVL7M8br41bMfiLTTSBS
Y2RupQmLmEhpZyzAPBeO8ZTONKSO9G9RxRYyRp4+hxAuUZIIACbKQj8G67d7blmG
ZZ0UEPrtugqX7mBd5SrVg0m2m9pzog1jw21N+O0aKJdPH0T+6LcWhogUiUzQvos3
m+DY8MjsVcRLBj29/Rig/AygkZhXY6xK5qIIVXgNTch6HwKa5kOuiqTk27f9PoIR
bPf1XJHjAyT8xcGob8zMho0YfLO8IHekqKvTk3LVSqTxiTpEfp6I/l+0PpSKruCD
JQwb9JbpJaMENIxuy6B9VYLeZDn+wI6ngRX/P22IqWtWmSBdNa9fYMK+8KKibnqU
qpKm6givpiZ3Fbvi+K1UVyk2Zu/WSGOS8zkgIozDuBeSQUiqZVH1nXzn2jCpK9pi
Ezyz1CcC/z6Rz4jEhRULyHTNHKhWR7BnRllahDlXh8+7GjO1/J3xSXvLpX7k5rTt
wZKlyyXq76gOej8Y1qTbXGbW6iesdzn6SF5eRp6EEtFqq916K0ND83pEadkau6A0
PeEPQYi7MA7TiFtaYCGbCXkODKgCvIjgwjVL+bBFYLyEc9fGmM0RGasgUM6XF+5b
dx+TDZ8eDkqua9tl/oG2RnQaT4CiWshB41lsrQZqMGQJTYygRNlAymdC28Wgek1s
uYk+6WM0zJojl4j3d6Dy3mBbuf/NVsBnN52wdqUCFhe1BGFDkkJLxBNGo7DqXylk
TSHEJX16A8818C3N0v7OjTP+HiRFC4tqNkJITUhcab7JJZKKvisJiP3rcv+FD6ap
VPr0qOzbCaT4i89nxPAlj04QfgbariQq2nJcSg94PaxgN30ks+EXw7F83B6C99sJ
c/Z+zkQMgbCTCLfcIpKVVne9WnHpjU3dk9OMlsVoYimbNOmFPGRB9NU9Olyh2vTV
8HSH6SnUR7hTjPEHUDTWInCXdYxaLLlCkbEYeHaPE5FR+xW4Ph+uUtR4+u7n4fhW
jybmTX3V8GFaw78tOmIqrqkmV80PkZyN/wbUcMRQBOF/IgCF7MDNglb8x0lccyED
9wcxtQ/maVGasEQNHjtay/YlFD+d50UFatAXnZjt2Dng6zIwGGo+FSMAej4LgP65
5OZkYm1MzsbHvWi++2a0Gz7PjmEBup6QKJRVYPOlnj2+8hnDHfDarvUHpLnvelgi
XQpbrobop1gWP6iCvvn5Yz99O/xUtzTuagUzQqknVCPhbUx3kGipMAMHzZjGXUYs
pwQ4zbVtMG5BrNb3NZCBvc9NLssvjww6u88Eb94UBF2yIXFsfrSRm8TsCuC1D4uw
r9smoAEJ78/62Gp1A5b6/GHTQXBN4774Qqz+qI3rE7DTM+26uELrRaWIPVM2uidw
OmTMyRnojgLgi6hkoLphRXPZsXcLuv87CMXiplzINSzQSiyFiotUuAVjT0dJqqvd
oUQYXH9lt7jsnGzP4RTYzWMd9PeiMzu1kR2AT/xeyyCtW3Sz4qpVwMf2w/NZKm1u
wofIMACY5/Wl+B3G91CawBveIExKF63CCyuLFirvFJUG/X+4Mxk1PAQxf7/WOw09
dDMr4BRRZlY8gxyCK4ApmX4AQ1smykPufDr7FF7WSsAmkoxKvw+bP0v988Tj5m3i
JmJYPjAiVrZ5BYDKULSmvn9LBMmEGai4sK8GHBa/y+8QBZhfvYZwC1IGgWa5nDBB
oxMNxlPQ0i9zLjTl7S54+PVCvszN5QQRA1f8S+vZwGA4Onm1ideJFVo13dXeLnry
riMLbpsCnkb2YTBBzr9htg6MjqijWZQY3Sg0YpwKbVII9Cl4ukGgXXj5p09a8t2O
gwVAsLzcfAt9kL2LagCu6UEzG3fDsGpZZUgZFihuvI+V0/x3R3lKc7dKt1Ycv0y5
6VwXbDFQc5RP3aaSwjk9ewMywLJPvOGY8RvWBMYVkzceeG1CrLTgsnJA3QLjfRzt
m6Dwhn7C+77fHKSx/iN3HIeVWljb7VukmA8X7Nz6AZepnSlUm4vOLyNJsZ9k+Sya
QsFEhjcoOGBmCQZjA3edCX0ZiAtelPLjMzY6hJwrs1sJbvAkjBYSacMam9FVC0/s
TSXV7ZXV30yRMy/AqYU5K9oREKnOK9LgZhmeyQjp193GWtJYqNRh7AvvZgjnNHP0
j7wVlMVY18IIP7E8xd2FZnuyGwI3ts4TorXZfHATbq5vWkOMSsoCWidz7bGDYdyq
h8/zS/7omy+ON5hzLsPXkjTg309C18J+mol6I9VhLzSYB2QdewXfV/zc+co01BvN
UHxNWtksjc52ZCvS7SfK4dd6bmtFzlZsORfH+UxeRfyxYZb0wYDsMDj8Fs5kM/E8
K7mX3bNxQPl8rToUVPwLSghPTK4GUx1qq3Nx6EdQpvHNzls8yHOydbV00k/dfbsc
FBgBWNqGpvJfHkrA3+ZQCQc5/pqj40Yr0Klplo7wwkga8EFkbIk58pRuS9tc+xlc
ufH++p4CTS+wIJQisGvJf0CZ6gW5CU+m0OzM5lJERkWV0sdfaze5c2nLbJK1g2n1
0CpPdOeBvZ+T6SdWNYh9ABQBRQLmNAmJsfrS1xLzZ7n+hcFYaKCP1+jDY9zJFMTG
QzVSNd4JBewoi1xg9nHAqyiDLSMWO9lz9Kf0Ij9S89CcdjmJP2yxy7wNE63/V5E8
pe+ZMZTgEDQapB7gc/I7oJBZgWhgZBktFTwmzmIXJof52Ek/mbkWKrYg8tED0Ex/
Q2gWf+tBVY1cZBkiErtPk1WWd5H5tqTdpVS7jNcJXxEV6fTAbM20qGf609s/1n52
w6JvK2GFqu6N/61ASQgWt6Jf+kEdk6WF9shfAs5Cg34lxVQi5O9kjtPsbOOI0Gg+
Y9jPStUaVXG0zQVIhKyee9ICV6sQ19sBS67dmKKJ5/CH9cDeHdzDRZgUn3HKvCa9
zR4tTbF2z4fppUOQLmF1teNzWlUzz8Rxj7fkNe8m0wl4sVp28QUavt7dBPioqDRz
kpaFQraycz67BtoAGBCdTYJTby15YNPoMeRBMzpqFmN/9m4ZNOv4eKgK8zLhY8ut
WOJ7v7XgoGMoIAN/UcgoW0cUo1TTol0+ifotJzt0D61dgKwFr6wRKNaKcXOpM4sm
JcwrJX6Uc5KnoVOOBCZbViiWOn2tNUSGgXOwbHbHqRauWY4kNKpAVNGgbzeB70TV
RXXVCw97sEmPXwA9LlSB6eGFzbG5G/YTqxGPsYIoCtVWGb+MIwY1WkMiRDy57e/s
0MMlKFaqRq32BzD+RYGKGN/waxvH65bfi0wky1PUw0CoThVfO/+qyby2gejcbL1Z
iv1IyTEQgcl6EX/n0e0fkScAlEQcV+xjgcgeI6V+o14FjeVv12PEwj+hJ15WVLr4
t/X8anZGiiXfgA//W9NXFZyDSNNfnxTrec1ou4Ykixh4grl+A1mKFutbDb2Fw1uL
RCry3DmxIQXuU0pcAX3dQTiMrvDugYoXGJZqPybWibe+LsEACxdLdvuPW05ybQSo
e9T2saX2ZXdy4m7oPiiW7fMRMS9eyWj5nCnsyUeZv0khyHPRf5mZVh7rRDHip33w
8DECiCgRX0POwJo/WLpJweQLMn9+hdkwWtUhZl7T1TaKCnt4HWcrqiIlhveWxwFY
EaFmoxMNmj6Zyel7IA4A6XlDtoeHdwxmtq9OU5URA6eMdZMHVBlQQIsLTbkSaL9F
yU28pMfI/QJxR7/PdK2B4k8VmsxmMaiyYS3AC8CxQ8TDO2gMgMvNaRQ/9F7Ojk0z
+41GB2X7XruYdPnHf58/Yb+dxyhN8vHaAj3SK5UELEIK3GMjI+dhFG3d01ct2vuD
kF3obcFnxhV2XgTQefwgTe3q00dj5cvBc7NALzPjwVsXlEpuh1aTlYhdr+NlndDD
b7lSkblMdQ/d1J7yLb1rlZtkBT1hqTrNYY6MHkC4hLpuscxVo++tYp+5YUgGr4FG
ko2pDd9bLhz93Hss6fUo/Dx8n4O6xtiSmef9r6hnLkkBTiR5QhRXUKsOP5xEXsvQ
oIaAeH6/DXbFPicHv4VN74AKQpY0jIMQfhChjxEfmh1uRbYGNv9FB64kGPYuDsVA
HqBoSbiXy0iip2y1FObRLFpdoX0YImo3cDXVDOGFYRkRbEBwnLNtvaLhhtYWr95U
Uavr+tVmXkLcP/AnNi9qBB9zngOB0AmELTG/JGxwzUQrzthU760iLUhGLFDt/DUG
bJHr/4m0moUZTt0u7kHFf3xxHdxKEy39UjT48lNSrkXSoh9xKTOa0uY2UNEeDaPk
6rUKuXIlsd/+5c4GHkk3J+4qAhB6O0nak5M/J2tcpIl387W7ybI0JGkVCQQmtXnC
DMQz6hAmcKj9/zJAqzV50n0pftZbdNSTkUyM8yPAgrtPprnTXKqAWIBUn7fRCue0
F7sqzKJzoJcxxRe1SU96sLE5XGRBi34Dlr9MkaP/KnZDB44nQ7WbW4BMH/+RCVXR
43ke7sKVENCNuIppo+FqiN4DuAoeNtT0Pmzu2dE4nNa9lnvDR1n6LGwksRBKRe9h
c8a4w7J1DO01qolL6xkh8ECOf4i0UXf0Ym2f/d/mAUJOTesxSWwxdiYOja4t8gKD
40wl3+tVvBBUWse1bOlF0a8saP+t9h5zWmq/rizBhWEzsgqtgJxFoSy7SWoH7psp
KDrT7EPehq6KqLE90XVU8D2LiIQG0gxGb1Mre3AvC8ztQ1TC31jgut72CYB5vG9b
UNB5AekYCqBJ+Ashegm3VMGWOukvfnWFUPYLHUlSST4oA1qqGZb6gBlu4CEU1laY
+FCLwwUDpANj00CmNeflSBmxULSZ8NWzY79ps7IXYjQhvbk7Sb4vT9anSBfR4YbM
Evcv7v+lXa4Q3dF67+Gjst/VHtlBJl16lAaLE4WIo9jEcZS362CxlknY0VMh4oQc
rSNWEEOao7PRyuW92AVUpfchr08hInds7PxH+2NFQUO9BRMqMZSayDwu8G4SEyOU
FgPXsbc5fjrgFzB7JCsboSdoYtN7WbLdmVrhV2PLhDb1nYFEEhN4Bmc72Eje8qFn
wBx4L00wsMZAky5uByADqndDZRM7PHBoFZB2LzCY80MLYz8VI+2cnUCmQqC3DMzf
KZ6zQsBXxoRR5E2lN4OcZtj8nGVDj6oBX/sexhgLg+GNR9wJd4TV0oIUO7DL1ZfP
T8d+xlDISUrZ5JBS0tme2hkT7EUQpGDJ1M8hELo2h+foiOKMryP90oZNmgepsvXA
rTx1UgWpwzPXVDsqvPwGAnelx6qNX0eKhecaMtyHhZ22oE10k8XDCadHBeF+Cu3U
5Fa2y7PEZUVjxuk6VHjRsQ15q+7FNGXGE/uvEJ031FMqaug1rdxoQeWnkAygosp6
Q3gjqrRb8RJcgd26CdSg/qenegLiPk1qJJ8x/YCThQiiUR9hiH+KRIzUnkFeQQMp
QEkc3EZ2hC5w5FLKIdUmpoIKy5LYjOsKLjT27lAJrqy4xsjRmFAX//GXRMij7jSW
DHXBkl+33ZeKZGGOJJFEGKhMEvwqVanRXiLXLfqe7Ds2yPJqIdQ7PyZwsgralGMD
CtC4qqOQMqhFfm5d0OaX1y72IlQeQconwg4rlei7jAROR7Dt1Nv7wosWAuH0F0Jp
a56qFccfsSc54vXc4+ZzV0MWrVqqRKnhgFk7D+V6Yc6+G3+DDW5dqb2bjcng46zp
/A+mtPFjWS7emROuPQ/D6I7pwGOrHOlVeZlDtUbopkG/8agxecyJoCSJbp2+w2AW
MImVR11Vr0w6IXCJe9WduyKaZanNqjhoBAu0Ur8BMDC7CU5xFZkNUplpFwGPo0L9
oFUrJpDryJ6MBgPuq2syZEm3TSkzurtryNRdLc/FF6wb70Tr17bE66cDEOwzn5KJ
8ZJuEYsPnzaUVVVdB9hebkTssvByM7RjoVx0yUV2yava7FGes/4sCIVfZK93h6n6
1SHDjHf4o9gjCjYrb9iQTUl23tk0B4EZO1fa7k1YVXPQJUZHswzNOK3XPTn+NAs9
dC/HZnFZYyBGAvzQ7dEorClmH8mRH2KJTBY7MjlBceP24ieBOgVtA7FUMqF+IA9r
FOlLPS389QXiGWwWB6rHgSfbe0WqHnCbRtDu9viI/TPvFubqDnSogBus0WEB/wAv
r+FVUlw2Gf+luV+mANfT6HSFw/s6JCqMbRimftUFseuvlGeb7XYxVws+knBX8AHk
IMPVPjtkLicER7kPP6WzZQxz8ry+nGphYWGK+LP6k25a1QGWyjanbb3wWhOR927q
06xNWjgeDgCLM6H58QllCBmZIU4NQkKH7++hO6G7a88tM08LpNOVYLIFj4hzW1/x
AvG2HGSuiaYVejdBkOh19EbKF11fIS2IKslCy2OMaS3G4N6SihB5PRu5qVnkMU+f
YDXxCOBoRR2AcF2ctcLhNDePoLzLAINzlPkbde/MN9WzUA4xDz8FEFBlm/e6eRAH
PCjFTqLgIRiFwbTCfq2MHCb1PoDnNbNeIqjoj5XaZfBt0gCkq4Os/h17gZEefhTl
2I2OBUm00GTuLnZpFWjFueeI//pxR/Sb2pU9uApxFTVHzXOWXz0+/rDNtK4kMUMG
lOlMg29zSD8LXQuXMxeoTIbTqT78ANavA+qr+lZ6QZHnu0IQ2y9TZ49ppHxLaXZX
MnCnjW8jDDhl5/lzsVhEutrTzQRxoq0xmzG36/TZ2qcb6t+N0z+Xs127JxO39iqN
gMPb7t51DmXWp2OJZjOjsmF77/Md7R2x5MGaF6AjzSplvN7Z5ekEPmCZz38Ofo+/
44djr8zakMHm/0rk1niL26ZmNDUkFLYaSlJWjjJyv5INNIRXLGD/CdmqStG7pTXN
m1tOTGHCUNmpXTHneOLOX1ZJB5xmeFh11TlgR+Us+NWYZfW72ThaBUkIrb271PIw
znGNhX37GdFkyQA5fmfauGhGShACFV7PueKfCsVrhFDjnEXlyHbdBqDpF07/tBNg
yGN7RSQRjITLoE5RN23FSNqCCr0bkruUN9OEt6wlRGcUVn3xr+x0IesF6GwY4LLT
e5hIZc6DHg8tAthX2ngRgLK8fhdDAh89wNcnQU9raf+DWKIM2Q5vcWIssifDTca0
IHWbieXCbBh+UMx8nEfVRBJnsxBm1NC9MASEeaYIR2RcqdOVQSFzYjoVWChpGyl0
/tQJhtChSkQJ84vOpaxiIbcNKYtcQyhBZiI2w5dpw8Ou9lWxNsQzNEYGHMkfr8Pk
2YFraSB23W0NrQuC1va9RyRlg1XVDzLXX1nvu9bpL/FsTSpkgnJwCpOng3UMnkRP
DcGt/Qx89IyqtDQvGQnho/eKQHX+SfupshNec6bE50kNkhf3gzpLj0/BHsJp+dE2
PGNBCz3jo/7YWL0QWOpmmS9frq5qgRweTR0hgwoC3ssml+NRAD91tAILYUuKgQBN
Cb5DlRnsmMECs0YwHqdQbcg7HrvPpWs2R0uF3ihAzM6bFpcRlQex+ZFTPqtZ5AtY
5qMBrxrhzBC7X0FhEKQ/esHRSAArXMrAOfVs07/Jh4oaLz9UxUrsfijaXzeSJ78l
0N4KdmcUajF1UQb/8AKQN9wJXnpEySOH/jR5rqk1KjMGXgEZDW/Fzhw0gIxAEY52
EOA8EtVGhryD595GYdynvnRfgzaqUmZkC4ErMZ7u/LtmlSPc4dNXF9JHlrB/d7L1
kGLGHjG/qu64sKctFzw7VJua+uxEjpJDflgGqlxoZSzl0opZ+QOLtbBCBTziiTFw
F8WxtI+lum1Q4M6vW28iYfvkURlSeQRSokz1ArhITO8bzkFgxOtf47sa+5mrY0Aq
z+gAcKGMti3LzBEhseIiEMWc4PPnlktCUEqs5hDyjH5n/N9VP+BPKg1GdGiphg9d
/gRaW6Yhigr9/Yu3GETSQd9ZxCJdaY5lf2KXDedQISRWWcArH1Ft23ckRzCQEOdf
QTi5uEGS6hN8lHVVrre39oM5gLESLDcU8fo6idQPHbYeXUmJtQewywqZ55hdw9lO
+AhwH/HHt+SSDDd2+p9jQ89KlDWNfghxXxvvpfy19c06tcXH9c5ONlbEWj3ybyTl
yv7Hsm07I1KefXvgJ3nM7OLlhiHkFMJTEn2aPwAY7X+N0MyD1jphu8qKB6ummnGJ
eqUX0ZyTtCxmmX+7bNSlVKWRCAdLtwYWLD3rcnwgg8tK8dfOxw/IXhCCV3BUAFvu
r746/iDINDaB/JysB5hAm4qF4hJzXJLAKFsw8Pr2raIWBTqw4tJsZmHNX6UedPdl
XA9PT6mzkp8kyNKkzVaat3A5rHK7cVVzs6Ysw3JFqwvelDXs8Xgz0x6mPSSLqb+9
/nuYJi6J6KxAh/2IC3sQgPg+ekPQoNFeJMal8HCjI1a86iZ+HS299VVcSOtC6mwK
ID7sgHj4DEEQRc3D1yVOl4Njus2aslBCmIyOAAjcam6Zs+JakqJg85f5oLEK7QwA
TjFfVopLMq16UiwCE0WkbkgE39w88GlxJVp4tdCx4SFJZ+uImDC4ZehkjQGYUJrL
IBiHDlVSI2FaAMqm0pHM23d6QQV31uYF73k0fmfTJUHcbfSWU5QKq8qOSzfIfdwt
25cpNe4SgfiWBeaaxCVswaslQ2JwiNhav+TTbQjXQL2iPizdidrv2gEP3Excx1ND
0CVFOOWYYVV0pS8MVL/KLvsRXSlG1qHDN+NVa12r5V7iKMJku3PXMJKgsbG3++50
yMDU0tO30tfm+ot9SAJrLtjLDo28dAMmbayysYc22Cgix1FGWd8FzMbI0IeSq5xo
QYZBojAnYSiAdGQhFgiisJKL5xeiIOj41/ocDI0q3YpsGzDbE0Xz0rtB2Qgtb/PZ
dsz3/wXNafidHOCaP+7dBaCnz8GaHaVQhP/GRLcDCaKD9s2iv/H5kn+9WGuHU/CW
cTj/57EbAjQFb6H9/u8NQSm4k4sdG5bApdR3hq1W/dYFva7fSnfccpIK0zFBiQeJ
rvxHHYPDypLXE+m3WMfATtIOjJr7VQzElCwxzk6kT3aNRn2T/QCCBK+Cpl72OnAE
jL6350SzGu+260nGF+NWmUHbnMWs6KiPomvN1Ox0tegofA3eisIs8NSc+C8ec0Oq
bCR1sy7iAoj/eU6Ay3geFFXeuKis7Y+w3drqrrKckjrhiYNP3aO3627iptEn9XJ5
cBDtzUEUOERQBBVfKyGed5ecNbtVN0h+M3nWljinHbZC8lGx43+TwfCxdAMd/0qW
K9A08+geImQXprQUNobcPgyvG0+kj9xSH0WHusiXkpMdVgdgJoch3o9AmRMt3wal
5lCfSUraOfrxtl7aaLeNoagFUaDFMbuZi34UzCrkbKMoLbT+VfjrRkbxwT8HCmyI
Ta/khDxu/Q80I9xoqUuUa5ex6ww6PPwk5hw6vVRXhl2qPsA/oKIs8fruxMBysKRm
hGpSbDK/poEj4njs7+Qlii1FuByAJKq3WPiHW8L3vB5nKvPNFHcL8hDp8Qq1xLtN
f7rAIeaWKyCRwtTlW3YaB/4oFzGhOCFAkQSdtAD/fwsK0Nk/+PPmiuNSgRa6mH/m
u8rld1nUROL1YujO9jecESonJcwXXNoK+M8kS8k1MnzMAYNnjG6z5gdUI4zoMELp
x/mzTVnE/wdKeiPLsJtxfRwl4yJpTzWeZEZkW5HjznT/OyL8EzP2yustj1u60gLs
3hLzVzsC3w1t+rh5HAiA9x0lFWhwX4q4NTV0WaK1RaAz13vaC5mEeNj7ZWS4yAWx
SXtFk7PpkoyjQx2vcO/7jLEmMyO3QI5fiF371pYu97XnfcY1D/MzIqeLKsbYXI2s
ejRjie45Z48/dhb9LkD7Tq3n6PVy0K2l7hReYukGibm+SAkdkD1sQR6oRgi7+28H
9jinotUsUAfnN5xEYy7v74QGABY7ykxc1FKewrIHPlxlOorUSh7BLjmPjfsFMmGZ
g++RKNJSwNNfxzm3NHQMIWU4kfkWPbKWXhXEyrGyrsXk6j0vDJW77BfSraOkGCSm
AxsXZJQMLQgfFmp0I1QmwjugWMa/MXX1hXFuBVLocCxt5zddFG1kFIVlxf37JHdd
19bWLEJx0cvnMDNiOv2Wnxxqu2iGoDZOSh4Ckfly6Us=
`protect END_PROTECTED
