`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNaD9lxNhP6woFtyLWPWzASEt5sjWxH6WM1nexmDoDylNjocPNZbeF/C/V9dOnS5
flMYbixI5HXFJwXsStmuqnp+6VKAjJTb0dbebrOVojxGcrLyVKcGm0Mwowoesz4R
tJyMUdgQczufH3JAPSfVZcTdMURk0aHiwkNkMXQHvyhkmAX2Y82skT3oQlM9jANU
NVVaxw1O8QBhOmda4z8YzWJA8HZQQ3wjMiQnlR1KHOT9xCvLRT/P+6qScOKE1XMt
sCMUvN0RyzJj/+C4NwmXasxmhp9ZxTQ3YMjX3cn+B32FJP/fqyj7wp2VvLt94FRe
kHQld+oYWsVH01p36mClqgXSq+k0OhkozizEr0mQtvwwrtYT8J9QFYlTC6KCMpH9
W39o8DlY62w76kWthLGezGzgzdO8x7IrEKl9vo3AZGn614yJzwvMENGsR8ZAZYbn
1R5dMoUCZVfQkru7ieXQaP7yRqZ6dcAOBWVYHffws6LCAE1xkm7onl9BiGgaVn9f
iFIeYbF0TEtm4PAnd3CeYIryKk9rFNPSTFW3wvDQonFqjOuHk4DFxsfwszXMW1zp
6khumip9fk8v0B6Eeep73d1+oCjKYP9vMQutzFV83Z7E1Kv8Jx/VoZqlfYJTj+/2
t9CGTB57OuZksbm/GAPgDiwr83IdmUQZVlTxSUwZMZVIufkoi+nU/FQz1c272Kfk
SU8UsH9kJvI3YR9x1fKkMAamT7x39HZCrBsmWF9bfDQA1OJtbKZUfGghHM1fKsj6
zUqUtFx1Cq25yDb+JNEiaWALAaPeWRDffjN2gnhM2q14ppJSGzoBmacV6QC/oSdk
O4CWHk4cP6z0V3Vz6G/oMxMk+k5RIQdHkBp+fF6Ptq4XkQ1jg9JKjRwQGNLoUqmS
0qEltpwhzeahvlgf5Sf6lRM1N9gnTJUYgrlTAKU84Cmx1RyWdkKxENim9ie8xmrX
9WZgjKOUY0L0x59GE9p3xWti/gQsq0gxRic1RdJXsOCIxZDXPR/EJSind/0k/nOC
z86MZsLCyKqZQt8tJl6AtMkCWMZePl0NX8sJKukRb1ledszIIn6yZbgcE+DQdDZp
LUJtOgQ88NBshSjTUJeAU1jBJOiWAKqtd/sLFZ7I1fypqxskZFL2QAd1DUCArY2L
aOz8tbQ7H9g7ErAmsQKEH5mRVP6AQFPnFkC8a9CzrA2yHlx0MiSK7aGlmINeiTSe
wkwj8g4KgC4SV7xl/GQCmrjD+IBRMXJ0fsDPeksnzRE4zPBb45sBn41Etczut2NA
WXmQgb94Hb+TMxtKvsyPweP5ePy2kjbby0YBp/RY7yCfBk9dms/JWj7c9wNJMjj3
qOBBUrAJvAfOZK442bNeXVEf44UvP9QIH5UFdLHwnMWLGbrGxONKMhKTF3VccmoT
mFos4i2Y4fgC2YwnepZE2liXDNaIWBLUawUpUkLC02HNLs0T736VN2oRVDoTofp3
93I9gnOeb+kXKR1GlWbP3VfYqOrnr/5yM3szfaVmk6l6BBxU0LRkEJBL/VBf0BnX
6COF/s5GeX/Ue+tIf8nEZaXA+NAJvk31JRtQX1L5sPfZ4Q/76OJ6s3I7ds2x4YId
RZWnbccNkh865r8F4LsRdSr+J3P7bc6mXeLOYplpW2vCDsuASHqxAG5T7wlpbqS/
pq9FI1K8iqlGaRpwQF0+pSVpKyiA/rxjrfsRWj757KCKQjTx90aNABbfi1Cn9T04
+BpxvtED1PjlOoxCms5KV5GwEcvrgXCh+V/o3L8CAHi0BVloIMct68N6QhjFDlro
7+yM629bXeASSn2vuBtYVyuRSxSmIWUlVf8hR/E+mDTKDf0tzUiJqZHoiwjo1TyY
OhDknmsN2DK/QT43LGr1yIv9abNrMdS22E47Poo8c3bl1viY5zvr3+09y/wKQjHl
CRTEwfug01yjS6uZA5y9+M2hj7mSqfkvtEfBW8x/EoqtXY5Q0laoKpcqdo8vpmAD
eHK0OPYap0jYG7sKL1AaiXi165zOUKN3vY69uvIjwC4DY5A+veYWeYuVQcxlkDa+
/iU5MeEoRwmA8CKlXAto8t/8cJEhuoZqyEcJma1CSAinTtxWt+XsCDtmDXM2nJAE
l3CS3WuDpSlQhDywELTXB0MNCLm7NhUisph0VSGIGMSHz84UpNfWF6cf6Fl8EbCz
UDkgK3Hs+VjoDb5duQkBvtg5XVUn9vjFfCY7TsG1sq8uCuf6oUneKB/JUCVYzLTc
18xdF2FJLDmWRQuXDb3zYjMKAA4UPU3Rw2kNzncZpuGc0W42uKYA/NvwBAc7RUud
R71jdg0Po/x+PcVth+26JDH2bLUijy0JT4+rbCE9oL4xYXFx+h1DH8EsfDUmo5j0
PrfQ8k5vOa5G5C0FfQtBf6bZmSam2mQgVT0K3hvXbZoYK001dfJPWN8K9nFzHBPv
kGblYpUchFSQqd/kpO62HcXb0BkRphj2Xo592eSvfBjDpgO7ovgCfJIPMBhJKlQJ
r/HA3DLCrAHwn58bc1+TMubJ+i34hvnSO9F+uRmz7NNh53s3Q/wZUM3exq2mLKro
PItFEPAVV1UqRgr9mIrlHOwXm9jd7uEWDhMDL5Y98J+w5L74XoBKcxSSKCti4KO4
1K92i8evqqJu+PvgSrPmqqgnsWEb1I3uTS1/RWpW7rwHm9DO6N/xbHNbDsOePrmu
SBvAFLl08rB86yAaQ8BCMuY9krI1BfDbS03RYG8Pc44f4N4Owpx450AXB+hnFkAu
VrHSuNAgCfZSolpDV5d9cRczov8apoqZ1kSWQiSd9U7pKAj5muO3F4FKkphtxSSj
dqfVBenWybJc0B0FlIe4RWP8ZpaBb2MQc7XbgrlWG4lUNZdF7CZ4HP3axKmLmgBM
mDPLk2duQr/o2hyNe8zbRiaJxEJvBA9kXWGvDSw6cKOThKEDTJ4TK9boHI9AsnPL
c0COSdxI2BZ2abeJhfQK/U8BWFIpe8I1uO5KbiLhGKcibYu0ftdunSfLoUobza+z
GJ5jYYbCkMpWda6nNQ0ie5d4Vpec3FqmfBR39X5630E4wKN283H0Q6YAD5qwC6kD
1hGz7HdNeha8cFuSPQ/Z4bfpRKmQRvRIdS1GEfGxIrmi2cxhZCzRmVwqLFP3v4Xw
mvOU9Md0506XBDzey6+3Righx5lC9CH4qRk6Y63kSgqkRTmkDFQBeApuTs+0Yjkv
ez+KEMlZeXncv6ifh0mLFhI9ab572V6m+Cps5GpWjHEV05NcLQ9HJ87rVjdouNVd
wBAuV3fi8jCReTI/rpyIcOvv8vCGCsmbB7tZv5i+4UXKtjCfNrbGfcErg6DFoLo2
2b0eLqt1Va1sKSvpQmYFocQBg920Grw40BRecebAIVFdG+IH6DGNw24HOI2watrL
KSz+4bCbIc5oTNm9miIYBwD7qP9VjRcTElv1hpw06Un2wsGEbOtIP1Ju4xvUGsKw
vgHHdFJZhSeAozi4Go4AND7MeIBsfm7a+nYSxENvtl2nTN/WtqMYsSVaq3mlwpDy
7GOMXK4Il8scVcCUOzvee7+LaRR1HkRvve5NezhJXyBQ+xw2HvZpEyuL8MpT/AjQ
6F9ODSsABCOGqtFtw52TLFn6WrW1iY6cSFAUZoFW90DFZXuFOYXwS5hOAqHLywSn
Dk5tXgcgSoy79lOvU6EtJKnZDyBNmMq/XyJZk8sX0MGsRMzxqwEyVyiDu4eJPRbS
6Ap4uIJOoY/zxfpqkFlafpC9Mbc6Z4qR588dpYstyMYnNaluUzKoUOQNKAihk4GB
RtfOBkI+qir9kiP4hKbwST/KG4sVzsT6eF4o5glwYB/SkP3EOicEK1HIAynV6Pb6
ym7yLCFswt3lwiVAOqolCeQpT3cCL/0oHjrAsXm0HfASDgVKTWBue90z4+qNewIn
2uoll8EIPgyHm+KgEftOVqLyfWr80L1qtB3uhRFEKupNSrS4esHq6S/83mH6PjAI
hbItfTSS9jEfhF87UUH5hFLWhQfuDQwDfIKDsF8tlhP0neDjE3bDXNs8RhPEhQsP
vfHKH05NArIlrqUFHNs2qhgY6dYWb91jAqwBLCEK0mx5gzLNCu1WtOmNwcLztKhz
+1bKcbCckgjJ9acdtfzjmnGFGkN915NvZbpGm9wkgA7JvYm4/veUgYSaGG734bTT
FpNwAvklRnRQwds9Lgh7qqfH8X6Icrhj2AGtdQzhVuWuoDjmWu7tRZXyd06qwOaj
r0aoaGrs5TjObNFrbwr2V+RPD4EXGQa3I6UHK/9q4v02+5uzyvS0rjtorIepxErF
Fq6yYKPykPPLYtb/QPy2UaeKUQxVNhaHLGSBa8A7BWESZu/xw9yw+dBXY3Ux7fU1
wmIi5Ujph7cROwKw0knNQEFoQIZEnf48zS447owP6cR0BEQXLnxciv1tHtT08Sot
yGppel64IC16X9x4ydJP76qXwebi+/sDd8MrpqmTyhaYJriQGJj5TCz0MQgbemOs
tkTSdYTxeHy/eGqBtAXSs1aHv5qLEIZXM+l+4GTouRUu1CDDmYVm4uOJmolqsfix
I34eAA0wJFoZeBMyX3Sk4ODvKkKh9HhIoAx1yy7KAB1DpM8JaOd0ZAuDyxItOIGV
JdBz2T+nihNhKaasU/inJsRJiaDVWMgdbH1f8Ke2s1/+6N4G7lWvi2bg7fiZ8IZu
38WPLX/f6MyAYMrJrESVa5VzwppsboEvjBNL29EstkaN0YURo4W3v/bP2q3IlL0M
XiN5DK3qScHG9jeOfuIPLQkUxDyrrTaVB1lcKR3RJqcDdMoX5G8u0GvO42VNwLPS
DJ23bH0fCuLjqmFBhPwYYe+kzO969rf/2sVs82GpVkgf8ZLl+vzKRnwLaMysEWZ6
bQ80lMLvxUOEidHWB4dlMHTJp0gLtFXrN+NwndCbS6lCRAm5C4TqfZb2VXgHQuaI
/pn8YdbguPBGClkPHpFEJD7bsPPBoSJN/pJBgV25kfupIIbNrB62pEtxrz99+jbi
p7c2ndwr6uytrhtFp0IWyOlPURD8GJk7laFGuE6/KEhw50i7h6UM+IvP4ErDOp2l
Ij9NpPMhwoYHeYxHc30lnq9Lz3eka2kqWgUbiGko4GV7LOb7h42Q60aUH74NOQTt
x5eD76Qtr7bHDOku6RNUhaoI5QTkHThtQLG3UW2edoLHyKl02r14kOX1LnwM4WJ2
+B/jkOFELfSPrZ91v1LXCQ==
`protect END_PROTECTED
