`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xztbLzsPgpaXFVnKVDKspd6HKYETGWohce1G1N1kHAde5+6hqNf9gXQtn3dhKj4Z
1Rl9ZdURwf6+Iubszgx5q/5FeNaRz2TTf5TKRreHJXkGByQyqGbBZYvR4fKoq9jW
oTLFtWmUoaR8h+DBhFVOKeZwX/aZUw/CZlig55weTiPpbVmip3+g4bFPSjNCzCYC
GGMUHtlvulYswT9tt7UW2uGVu1wzY2A3hMWKGcFrfmSXFhRx3ZfKyBY3aDnZpNrL
Uz36DqOiTfE3SjKIo2t5dwj3k9cG1WpPT8JaCfNtzvYB6wSqum7Ix+EbRzOO4Nx8
F9AZLhEjSwRlSCPw9th1prQyjFNla/aP909y6a3l4E4ED8tu7OFfh8EgMoGJamXE
HqXDSmB0JQJ+BJEQ0LR51i1k54JSfDwQtJm36MMNVLvqCLAYalzI6a7woxMESbTD
ibwXk7CUquPqDnKNQnw7oM9AtrNDRwjhtceYkbXVQbGbyRp0sONls/aoLuv3cwfy
BAT607H80rAndTpnj79lmlAlDtjrVwf/0OkHh4eAb1w8TZFqeIBzUlKW/6pGX3pC
p/CMLfRPEZGxf6G0UlwE3+SF2nl1Tsu++6wsUt7ef+DvdoXIQmTwWJzGDXWbZSTi
J2hQJjZKSfyZy2Et2ks/onQVGS+r2PlX+J+dAIhw4gIVSX4i99h3Scxw3cqS3TEi
xNlivN/VtdekpmxMYMpbhEXMp+KdfIV7b1RHTsPu9iyEdhbr4pglznO1iO4XbEwX
q7ZZi1WN0shP9TPLNg2CWm78Tb9jXn/U/Vuzf5XlT8sxURdLLkFzZspKJX+QKGRP
yp9TK99RrwauZ/aqrAnIpeNKtYBrLnMbeL77STtGyf55sxQQqJoVaaLTO+1X/W/f
apeKCho+frEbLuoKLJN6nKTIN8POJjbxJOwG/2Xxle+vikuK4NoNhPb2xmqVsJme
RoBRga8WZxfWAcrZMS8ghoMaL4Z/YSfI3mWvV8tHLS+rjDKUQ53C5QtUXlRRnn3D
nq0c6bWodLgbj/qylIgQFry5BDvMkBRYhgcZjGpC6Z3y4KC2vX/CVO3a0xV5q3nk
8KJ+JTytXvXw9RxkVWvGxX8SYTlA5m1cYb9LGon846BQUNSreFyvElqHrEM+p4cv
CTw6+RgUGmpxnvlm4eyNWflWXDjUhqaJSqoH0OeGmhLYlRgzY6TWCJ7HQeCgA7+4
oNLj7uWnqS2m7hd6o3mihDNQTEo5sIesa7kG7UA5UhAwA5x/rnFdywwgI8uFQArk
f+izHJb69lXgY4EH4bYDDr3yUz4P1ZC89qJ2tvmQaL4=
`protect END_PROTECTED
