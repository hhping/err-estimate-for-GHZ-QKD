`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGeud0yhWoQAqzljX2lyUq+1I8W8JVKTiDcnIVKABXA57SWwC4XFYAFnctVbCYk9
wdArUQJISMsxZq7I28IKvsKK9aAHTFXNDvmIccASpvrGJ29GTgEU0gGy0NGNxP8S
Kgr2jUHfs/GbGiH9qreNqM2rVoh6aQoWrIHi/uP+5Q+QH7xUHBQo0+y4659wQ4wZ
3Voitfbg0YSnJ7dbbqNEF0IR6cklalgPa0zBBdt6nRyYOW5Nfn0nkrhfw83gyymB
4mOz7ckH1q37uXD5o8n2+9VzNk6Lh8D/H4aeuRuFMdxMFYzWZtBzqq8cfKrxz2OT
b2GQj3QKuaVYSmGoLkM1kb0+CgTPjlq39mIf4ATrOT2ZzNH9hZZbk6oVPQ62iOXJ
oiU+aC/1eTA3N1dbFhqFRJ7jEonBx0Y1FawAohZi+vLv8S11tPiS8KbeE8C3YmnW
daIdtc6QS7MY0Zs2ELi/qdPV8C4AhgSA90Vbt0dbDOWIs5etqx3zhZHbAnMUShBB
8j9H3pTO7zbGLJpOPi/4neuZSCNgtfF5ybXeTciB/kEJLVWw7iHTvW1DIv0v8a9P
ee7Jcb1j9kORXnbSI730FCxuvbGSpBRvJSdBbth161jR6l3fiLAtjvPLqiLkNy81
Ufvcp2iNhA7NQ9Rc6ejRHz87HF1WC0kUL8BW7tF6lEOBSdAqsWu2aGopTUeEXODv
1VY54YtnQbxY8W/J2Gbly0HH3M1PmP8EZLOZ9COSNNDzN5L24cyfqG0gQXVYdGBc
6+DWHatKmGjvrh+I3ZGQS7fKxe8rtjO8kSm57SnPSIQnbLeED1cK3ahf/jGYayWa
toD9o5LJzG60rq4yJmJuTLS/hl6CYCUX7c20/9bbqCFlc61r2tqVIZt1EM257RMm
NVbWeZ2ll7MH+iXpe/elUZczjybtVHWXcLhCKx5RAHDBO1MHHDwHDZ9TxQlPOrA4
EMIt4rZXOAHMTAp/LFAegbD2i2+okkllEOH2bap+LnpszLU+zAK2i8rLi9Kw+P0I
BzMnAK0s32uIgNkKda2hQrNO55bJaOtEh06YXxL1nd89ukryLKZlgavEGlyRbWea
ls98OW1J6sNB/+F6Gkx55ZzLlFIgoI0sgLt2N90YDGnTIgDD7+eVqFkGzPU4d87m
coPjhiNu+lrAaa3a4zZ8eSNS2zSHOaGcqzjk/YQpdONv1LlQIudzEapuwlg9+5ek
Fc4y87HTiiP2wD57WIZsLGdTD9suFDJaw2NbD6n4k2n99CIFaaIn0WZUmYN3l6EX
VPQBFtF/cVlPDx7W7YbvKUYQqUnMIXVe6ayFN94l9mhJ3mCcy1UdheWSEUuv+m3t
sEhEqMERXVdxbV6w7M9tWKBxfo0oclHRuZAu/F1s49K0dPmW4CpyWErnyFK4bk/u
+nGffnD3jfeU1CGHfgykDpFeJXXFkB7zHx6H4USwMQPTEHBdPeZ/R78TvQ5SGYhA
bS2QZUrOiXy4w1XfEL+RZs0ReGNDFL0SB4C2CW2FgAIYwmXKqyifHapZo7bh1wxW
r/V38bKVpc0gKOyLgycD5Nf7d6oZDFEG/Ce6oCc1SM+H74NCBv3AlzklrdNVi0T4
kWijsVsWwsv29Cu0q9mEKJ+gkfYDCTgcspcbSF9h6TorQkxucBDh8cK1ycKhxQHa
3qswV3lF4IdNavL9VRjM7eXAGw/xNxUBwJp+dzyJgpjrRnlVi7tJY+1/BbJXZ5Mq
UR/IbM6Rr9ulPXx6XPg5DqhOu9Tbm1MuY6fA2RznaNSaUf0YhHQ6f+NOjdwR8IUL
lXA7VOZ1IeoHxLFjhvH9FeNkP8D1N6i7yoUcCGozG6g2srFRGl8SDdCYlf+REtAk
8Rs7av2dsseXJLEzdOX1jNw2rNKf9lemvQHUyhX26RxGZBo+CvTqaK2bG0tYELq6
DD7HlQIhSYRcLTet8VjjMsHABbFPF7/YyXW92y7bNXNX2d5tPgLCrQklqs/63k4C
TECwfTdp4VkuUOrYpWqCk6Fr78YIAz5ydpALkcMDogddvLENifulHoInkL2+XLCY
J0zgjTrXK7ZFbxLvybeFJ3i9Yvc6R09wgI0+ZPpROr45lHtgAvY6qKGeOXm2Fexv
P2s8vqXOA6pIQ8UJr9wvbWPGzZv1IfdZx7VoXh80dxUFf3SyiRAbvRpGfauwGCYM
yd+8fLWap0l/QBV5EPW26C4KEpd/+q6JG27uq88QQsx7Hw7wt8BtgSqKZxMI2aXN
UKMMLHuvubEukPMoeAImZgPdCjUf7X3WPl3M9kCV4FElYE62Vq7uXVh7zlhNPqiw
EQmed6oNwukwhd4eRD0l1PgxDd3S5QX8kVk3hMQNdHjtPAVh9cfi6Q9l98q7you+
VKsnI2IVfjDNohbQrAYgRfyirxmk0+1yEO64MV5iDJ0wRP7wp+cv6o+zhhTqC2Pk
6rH912LF650dzAqS3FoXMiZ0ZYjYP6GWyMoeZWZSFSOBCXwlkP2wRNU1dW9Rk0ir
ocGmdK8hDufd7MBGsmqEFDhMw0jF7a7tdquay8tstYxwiF5VBY5XfxEmGHBXqVY9
xBcASWTdFuqa7YgR8SidiR9SJbkD5soptY2AHxox8WrrVd0lA0UojnyDj94tI5Tg
tjxXr2F/dVL+Rv4p/zdtbv5zwlYCPguvGfmw32haDSjTVO9191hb+KVwT59ACao6
HMQyHUIE7nqnmEaBONmmljyz8hWUS505yN04Pu7fgluNKYl6BeNs3aCkXs7JxbYi
mAkxey7wtmRqtV/APls00aUZL/ujp7X8Tk8iRoK1TOzf3biRPFwdc2qm3RVlg7Rk
aKFmhSWRsRBptSCzpoODgXBlaA34CbyGUCzmTbEYx71JlwGSyH4R+5E7PLzYiZR3
AlXmjRPpLowR/1KVi632L/w4DspAA/O0cY7AXO+nLWweAK1UypCzsVFCZOshz1xN
cOiXyR1qSPdfsg+qpC5KrNDbfZ71iLvIZBSp1QLeS3QXjL6rxQRaU7FM92cQUAW8
hQKBx7p+oHJPv2/qzPyHgQ6DJ/xn6hfMpdd1k9Ult5sYt9i09lp6TjRaio2icjjG
TBjesHY6x0kY/opD/XV/TQBklpZG4a9hd752MN/T2SM5lcqzuNg1gYnWdafjUAqZ
nMnjp84VdtBNnaUOVJQ2/Nn4C5nyvPijbj9d+GY25NYfQzbqazHGgJNcsDhAnptv
jalWLSjTCiEZ4fHp5ptxQSEGjkmu3OoK/4trYnaWhMUqgnouboquTfesJ60UjIQc
lHhSn9PJUnYt/7ceSpVLu9YLOolBWaMo7lYsIgOZKa3EDHgl1HkSa/+CDBKQjH2D
pYXlKoN5pN9JU4i0WKscJ8vJAeY8GMk3s4m6scYg8VaQWMlpsTM34koFfikz52ZA
3dEfDYs487ds/Ga7STIvmDl76J/HC2pOfLcj03iqTNh3FvuK8umczyVDX+apydM+
sMsLj5sZ1kg8xT354XQsno90QgL3HVgcTiKeavXVvnIvdTMlOUSOi84vTWN92bQo
SpAo+myM4H63aVAsYvwa3A6rwPZrJYnHwTrfSqcAha9a7dlXf3B6nmtdhmHzpDQn
d2W5//aAE15qeO/TzrkYrz5hBm7Ghk1hH6Uc3n6iG+CKNU6MYqyVupxHRUZ3sG7E
ty2CbRvwSImPme0enoUG3qPUXdmbIhC3R6tIWEn7KuY1H5WAykkclfLktNZaG89f
NyiOn8MT5hhA9TbEdpyOQnZ9UtveweTs2CubQTxEr/nHICMFfREOC8LRjibLVcTq
s75b63czarJ2mWcCk+oaQSqwA5eAGpw37ecLmm5WomdOIGdTzi6sPKtQoU8mf5s7
mI2XAGzDMkLAP/3+LUzQmJHxMDdvcNrgbquZtOnYGsMKTSGbM8CxwP+ZXwoPxPwR
D04A0aZj2q/VefYS0OdIgIM27pVWlD8PH22L+t3RDZ5H8V8Bm+hdeuY7kAousGBl
aeNYmMcHuLsedljsteZWQle+u40Jhf1lQK16jlrwKx3z3Hkx6fvO3gkm+wx4iw4A
tfFCes1rdjQ1Cdl58YTwHWmVRf9uHLSYYw2l9Vc/Fea2NEHpff2RDHhqMxRG95jN
NeG7bkskw33Q/YFmsoafmRxNXb/TnosNkrxpW8ipW8VT1t6t96K53N4kywxBWUap
pSva+aNGTPGJaN0t1f3GXIVYobn04nyaJbP9vGKXCAlRTFP2B0Vr2NQ/z/m/WgJF
WYy1PkeaO0RInJlF2sTayy7P+IYbfpOfdgfSK90IDV0k3iUlh18Gn7XvJgXMvUYJ
NvTLnqrM93tb9vz/RXAcgp7NiL+LBozL8MbB9xddXbabK9dAVEaEmQkthY17M4oL
74imyi3CecllaKyIT7ECV+xuCIcg2aAFBsJAx8lvXvOSdI9fTZDiTlG8myaTWPVM
K1CVuONuxALvEICIN+hcURQEvPIkbdwVFeyqtPTDVkIu0obJuXVpLc8fxXefyF60
amISRVdwpM9Tzk3yPKTfQhAhJ+vfH3/fcdKNjfGtQZyJUSrlh+8o6Tm+Yjkf12MW
CdhUBlSDjwuYBu0KNjqE8iijzp2cXfrVuTbeCqImunMcN5qwdJUQKRTh1knkf1R5
sfKPUOmViai3FvgUQT09FRUnCqrRWBW6pcti8n7eyBoT2w2m8hSurgs2BfWawuc3
zvjrEAVsGucuXl7SiHcZsdzOr+FETczNOxcd41rgZZxIIfbJKnCwndrnND3o+WaJ
MD2yCZdrPfpTBwfWZa27ETQyJb9/o2xu1dbxlNiNWOwq4DzyC/ca1IploC7GM3CS
GJ9hovGyO2GHYGYnkycuY2+5IASh/Fi0mCpPY8Ni6K9JNWJ6nJ3v2OddWl1dIX3h
EC1jJmXZ5SHqa1rraEOw7pb5m45IKhtWx4NsAyUc7ffBpuwDOsnWeFVfemhWFaQ+
KwyZPwvWW8U2aHqNQQn6ECx7xnbf9zH7S08ScdmtkQ/oa0+/kyNeaEtqhKA1ohxm
mqT2V9PXx8EVFkzMmwQQD2RHEPlYEgxJYamWpZyQCIltsFHDlivT5qWr5jGaGATb
Zmk97NxAOaBOKM5VIO7Z1rGmjiAmEjJB5xk8XS+kCMbrtyA7RTKGGIvUWq5ry0e/
9a2rSc/eKzUNRtYkRG4h16zm24bSvlOBb/wfZP97/Ix4PU3DOUH9ScjURok/qelb
uAqHWuSRvjmG5ZYBJ2aQRA+7rF48iT41qhLybt9bLzJrFvYfzm9RoBuPcDS7T/tO
YvUk+Jll6DyCbP/Xzp54GDvy3Nuxn6Vkl8RvLA7hiHv3CU9+CTZPdfhMkGK5Fihf
5rrmOVB/e6zo+4WGjH+l4uI87FZymbdHdRa9IeRxY+W0NtxDAVQXrlbxEhgSbbcs
4+WBZIjEsJx7Rs/GV+nOGq6KKtpjaqoiNbjRPQl6N2Pvqxh4asIDiK8ZXzuFKdju
LF7psBxJX3WV28xm8Fx7VnfgBYqo/chozWcsXK2cocTXZy/BH03+OFcTegYEZ+gw
U+D+eGUM2ARClBpkmynEMAxW3zte2d/qLVF06sfbh34ecC+yl+pcWgG1pYHTph7I
14QlHltm9+pipuK6C/n7DR6HpLpVMYG6ygbXZlewBYEEB/5FieBlSKGHhMEVylNV
zn7AX23PPdDMbAF1HLI6V1t+tAQAlD/OugZCuz7+Bj+iN/FCTc3FjH4X4lmBapJN
nglnnklY0okZPgKr5Vx1C3T3OBwvCGgFHDEbf4+Lt5fJKOIqS+2B/Ooa9Tp934qC
pQG3LoIcQdxt9Nk7wIa0f4QDxy8tIMURhhF52wfIUwDu2jBTaob2y0YjB8SJhr8a
XvS57BTPOvVPFHjJVfq4b1VlMlcpZbO4/ia1HtEMYvrKemj7T5pe/yShbXIAq3oq
stwe6jHuFOMQGBBBfN30RSVIgqqNRKazzHBap4bOn4s2zkTGsEvhOqdUDixely91
2ueUyvXeNRJT8UyEg703EhYC8TXVbi4mYo1t9gDfW1o8uEmQhh+kH0fyl6hz1Wf4
EOFfsUjQTQtSyrIhLUjHgonPwrxrnDEo94mSl/+SlprLQXVOv4+Y5vUUvFP6azF5
hDyV7WSVy+uPs/+Y9VNxlCo+poiDnbAEz/owdks/8oUA7EvlB1VowOj1P4XHeIE1
QUvPKSjnpzEt4ypIF6cu+y5fIjuiwOmq3+nHVRlOmseW+AYc9IQmfeR+WU+eUz9F
6hGrWOuKTPubBSP3/GO48wovJ1uI00uIcMkJBwR6bqTBaQZMlS5JY/cEwbccRhdX
RHowBSkhDsQQnb/fmZ1pYFt8cS8QRr6ZP2bp0l5hYwumESRiyxbVt+Uv8uLUciQ8
Uo3P3OnPR6Gttf5gN0WWEEcoJEwbd0qce/4/f1+G4Dec3KMzfKX6m7sJWLCAosx9
MR+hTFyZxbJ1E+g7so7ZHF4K0/At0V+Sgsp72PbiCzPfNNuxUuDEdc6x6DfqWKZP
Lf5hr0d99OqgwzlurlbHCR0aCoHDP4iMwjjyES6KD2iPDQTvYDf2gK1l6/9ShIM3
0zuGn8q49emc/bjzOgW4kTwWrmENDEw3hTh3W6iu0PVAUrLZDT28WxGZG2waRnrd
b/DIMSpw0OD+Wd4irL6fMgwhOQKvYoK2iLBGIPcFSajI1UL7Lnd2bl4fdHDjZZI0
bOC/xYSnCmKi6YXEhR3MBxAeLfpdFgPdj7c0UXh1hi2hi2dxNE5Rli27qoYqfCmG
4Qhi11nfGTCeQVlo0j5uTp93gClkTZ2FESSoNPoc3NxGWgNrJhUEDfAPnd5NOWPI
ykQImjLGIlFaTF1c4QTpz7qn+LXzMgUhtrWFGusbLQGBV8+13h8xfzHeLCl7dX1j
4QAnQZsV/+E10k/aBKdtY/TxZikaMHnd/1Goquqxfop7kwxR9LZkehHI2Ul/pNhz
olV2J7gQ9lvjb3kFp2tHMkjx8UC7U/Ofj2Di8JwftxvOwipmttrOr3pPtvU7P2Zu
+ScV81b59CvtTvbUfoancIkOF8uMXcRo2h5yJE572pNvnpj1XnMJsKUpAb6yCUn9
H6Mr4wXkxHGXQCcpmu1L9aEHoevvgCb8O8a3WHUMIDuaLA23uaK9VHdk65No9U/l
FyiQuI/4+JGAhF+FH2GOqd41b+3TGRAjubOs1ODSR1g9s5e+J8IlFi+sTWn5iCtN
MMZFWmAsafBoJwuUifq0sW7RidB51sS7OIfWGbVukcLr4HDJZJvkr++DmNrJY1n4
X1mj0nEfP1dNr7GEx+HoojdAalfe7k1NdsYNJgRD6vyuXV9OGhqv4ak5ieHqxlXt
s/gnhkOPyzoPPMk5EhnHPzSDQisUa7zTyzbU/FKKhfgWyNWzEArma7TAGkcev5KW
nvGPalwzSastZGmp0hBJjUoWJmCD1/xsdb1AQx0a3VAmNnlkNBxpMOolHnHBTihU
cbPl0quQ4Lm03RItK3zXaiBzOcMreZjqXmAC+98tElN2Zkt4Dag1X0u9tcL0CceD
/C8L82ky4VAjRd0QpcAQx4CYvR1MnYBr4WiY0AHrzepIviWaoMlDV9zJm34y2nMy
Awp1w+gY65ivimWN5+nVUWzmr0YXmQVBQ4dU1KHR1wniCLXs+k/Sf1yHMrG7+ovU
wh7vpj30uaMM4qT5RND6ZUpa1bWZ+aPQuN1SfAKt9JocVs1LKYW4q6voTpbmLAKH
cgTZcaOtsHbE1gSJqFefL55Cq4TGSV1UgAspDgRlSftL7Bkl/W5YP9S5X/3YoidQ
C+vCPEpPpVMR1OUbsxUogKx4DUX5GT4+fgWYXyApOlEOi+hdsJ1qUGk2TeADP6d7
RMWccNTEq8NFFH8oe5WltKsw31CLLKXZ4Gn8G01R5clM38GhLJKQLRyZP9ZEs0At
NzB3vidtJfY/JsWOrjfLHtgqOJSjd3OtntC1J7fJ5Df8Szbglu8xoTKymXg9gQlr
UkXDwKR3mLbHwKyZ9TNgwobYHkk9cgomaLpfqmMkGDZF34J0Sr4br+Yfb6/Nrp13
LlHia1I5Tgs2x3ckHSWS0C0KxEX4BIMbQ1+BmUaz0PfM+12MYfhGauu1cTugQQKH
pZGDQhotmUQhwtJac49DzaoWSnGOYXYdFw5mkr1sDyNSpvzUuOhj0cCmqSslDsRI
trRb2ThuIfC7rVvLQVIbKui+CPIJWw5f4OeeZE1LEaZHoWXo/vmjqO16b6UNzqSA
y/OnMM/KWACY4MVdsPsV5YJrOBvD/ntLSIMcq+shcyeqV39WKRZy9CTIFE1evzd4
3MdwlqiC6KXOTEWIkPH2lcg2NR53o+VlDJ7RDDcFcJTMWHnBr7mFFSPPSAxWtEnt
GPvXmySVv6AlVwgELjZihinPLyqS7HLB2D94vNKKMj9FNyE/d75jb6VFbo0PG/F1
RBOe022XwwJL+XkVmoCP41YM5y2UihtpJl1Uc+I1XDP0PpNqACLbeywrPx6m4W0v
NbVN9bL+KW3SP7KpAvXybIbTlYzWUp7cJ8WT6mWP4sAku9MGaDgyg5xioGrTP4T7
axmgXpmcDAG+JZUM7fGaU0MvZDlpqlBFqDIXpka/vypNi6DaPvkXmqMhsXFqU2cN
e3yDYkDJrfw2RCcGgbny9KrjF3tjEpqz+ae1pTlTuPfrf0oC8afoe17hE6vPKx+s
zObH6UY4fJS7E0+hjx4QFrAUVL4WrnUziRFlEIMEpB9E2ob+QXXva8HgmSqz98W7
3iIeswq74m819xj/kgRRqOoueDorhzc71ZroVOslAd73ZkmN9+YOn0VEShWTVNxL
5/bs+lXb6MZUlQoaVnaO/rCuu604V/btfC0ulFkS3IHXkLl+JsK6NQ6vE1ijE3M5
c7Uxx2hgtAf1WxIqLdrwlVRYGArfJDA+9hFOeoTH03//qegfqYOcYaeAjBfQ4MCL
cUJ3Xjopv7kplNdlKSr+b8GgM+9J/scVNBQWQacD9/Yafahz1OsqUEE79CaI3ti9
jxlFGEcYk7r46YY1m4HXpJtey9e71DQQ9hiraHByMH1PWKDqw04ecPhmDhfv8lmI
y1hYN3/hvpnlIL3Vsa3KX/WSgQodYlm2TTdlvFud1HZ1cBsQ98wzkDedZ11VQN0U
zxv+OLBicai8DE7QCYe70BZCTcWOkX6Q+GBMt4SM+3GksfuJt62MzTM+LdH9qCvZ
ThoCtL8MMSSEKf57315j1TVmLrF9PisaWhAoSm0sbBVi+26xjOj6E1iREBPqHzk+
C2BzegjHDIZH9emLyb+wHOBG5r3KRHBeMLivrOyyybvWgYRbRxMdJs80iEHig7s7
5G7CuZBT2ZG0M+XCAWzjORzRNkvD02ONGrEV1c+0Wbjqr1b0VbcTvCV4zU+yCsoK
iG3Rf+XRQew+pzuwEd7L3VPP48SamNhhTyzWgN8V4FGy/MdOrCvWqmrv1cNeRh4u
PGvRZoOM/WRhFONEb+CpcmU6JwV36eFvPpum7W/vOzMmwNY85QVd8gbGTCKZGpn4
Nv6IUDrgepuStPddBwW1oUlnUCm+eOJt0DYnaA1gWunWCxvsQ8Z0L2+OSmEzRq92
UdMyneKCbZaWQUZ9uuydsdpz+0j4BcRrmCLeJGkwQxvzBAECgO8f0tbb5+Fnebsn
//KqHEfYs/GK8hs6RAOWaSNEr1MudEfCl5Lhi6E6t45ESUmEtvUDoJsC1VtY6BhW
QHzIJB5VK7XOY+Ir/gHaPKx+VhNKLofOjBlPNIxn6kIGxsZ/yNiGNBeS9vzSi86A
kfP8OM2pItSYn/h9SwWI5cFiB2GwSN1/qn6zQsb3oENwtqfobO53ac6HvpjqrkUd
kuqCu5HyHcDAbihGS0awU6KE2mcR6op/xP1PdoFc0KRL43MGe/zJgVSWZawDqSsM
75/+S3kk5mj/EXxEGjpAE1qfz192TQpfMNkzDKagcL3Gd4QDrWRg0CmQBrbnKflB
Ga1nklbertUU//yAE/i8bZwiVqSBiCpBJPGCIJ1lacGnmfyFd1XhS+MDBSdxRMov
NUIDA+0wdSXln3u29AWREfXXGYwZU7z0VeSY3Epti7zc+mOdQXAnIo/ZI4cEB5lP
gW6WoU26WyuzunpcIfufrMz/e0QKx5akPFjsfKtIVjkNpLCNa77fms6fphQ9nwSE
WlnIqKb2QA/vc5qVLw/twowMEqwNvkfIyoZOuSwWyJ3xR0CVGyzFyvuwFYHCB8qc
QUBYwLLnnE0MG7KvIqjq0UEYAtJWQrcEZ6DkQ27ukJfw0qR6ziUc1kZf6IkC9Fmg
ZshchygraVTwC1IMgMEb9ZL5WlitB56YLMmp/dBqUppfdsmybmkE1RO/pav3Pf8Z
iUAcwrXTr04m1kPPuCSjVUBIO6JLivkiBz3cFewH4phPSWA9e8TpixIMB5lwvCu8
mhrkBYsgBO0x6VKBO2VwMXrqCZRoUHgl1aPcPj+esX2vKLd9bepPJ2mPgT67spED
yIBCBSksI8g52x1tfzlU/F8GjGHZghecXEtRV7ppsmwqyLL4h/JgDTOI5xlJ4CXQ
9O+k7TX79dqsf5gDjDW/6BrOmJTkLw9iG+B8aPzcMgU5snmtEpeb8PktD80Ob82J
f4L6QLyuszW6N0qVErhY85FGW29UK5wSEVnQVUlOnqZbS3ysKpALZdo6vY+h2xxf
mLXPoIxnT4l5PSrOfWbon47IBVbi5KQA2cPr5jhTCPHnQ7RiqTIWN6FWfKtEpXMK
wVrPXhSSIBBjDrtXgePczUEJrCJuqWWNuZw7x1lKerDQjLJSmw5UxWJrQENq8CwB
tG6nDIDlpNKAgMTu4RPUZafvuNK817AQouqm+m68cbnO08jf/89BLLkwF6x/SKrw
rlIdH1xLV6nS2iZdTtrPiQE+1aWbk/enmmzjsiF7MmtIqzFGZVkHENKnpMqc0Ryh
kixqQINaglZ0c3z7jjpL5dP4RXp1ePRWm/7U6gcjHWOWN5ER1dJMnqwuUE4tAhzl
krQK57AeUVVJAedcCzbWYT2OqT9/DDqnuaKybCUUnonrHgaeChkeMKpLyC2ySAHa
ZmSnpOvGZ/3r0YmKyFxIxfoT1TUvxLC6wk2ZHZOYoGD9U75ml5eSOT+g5oEKoygH
WsF+mW8aeYGCNrNAchXD8FnE54R9b7wT9pdtG1zBHgJycSD8SODgG9ryNm5VkfpI
zf55zwUG4Ju29+XRil8lmXyXQ+pO5hTHzR1idbhbxHLNMfpLahTRzip8jcI+sF3m
0sNtVEifAmRJDFzOJRfwTlM55ANy5yRGWHFWJbNfwk/1mjMQapyzmafV6Puli4gl
Ny38fI+l2cZLwwZJ75/7en6+wdugA6uedjsLhadVBKmG1IaivL0rTKZTyTxpbzlO
7sFq0g/6kfgYjqd6YSYIjvlvnTqboAjX2cxxvqYyJRwtK+Eh2SkpoVO1VG2K1RHx
sB+j22ALES3LkmxF+Z5JNoVhPS67zrdDb2kR5vrpUNCQjw9C5luVbENCss/cSLvV
jkb0AL/hN9Fto3Hy+T2fEdH0RGU+68Uvy2Q1c5I4xKU8KfExZhAWFIlyB8DpwVVb
0UWBB0AvUTN64BjcLC/llTkNBqhjSK5b/Whb6k5JKzyXu5plJbAFpPxl04C+VXoT
cFWzPGcYkXG1Mq/1/um3sl9Y8taU5/Ejb11zd8vpv6IXw6g9MGEi45w+hed80i0I
YXyw+rjoPc31HXPDKhyoZnXvGbB5SW8mpsujm7pAL1pNyBYXtZq/HG/ouCL0lgWR
Q5MLnC/Q+Efc964g7RO9F6Qyuoual3tyUZtGdl2Rsy12Bl/YZMLkYLNFBPRpuoR4
unWePTK/dDLLuXJB6y2KoFednHfImxUWuFcqITUrSneidRZX/apQvRSuL+mGLb6y
p7GZfDEk4xmide89VjXUWTDXn+IXFTsnxEdFxXxEixjfdYUOGfQKNbD4pPwAEs6T
C6IYUwlcgBM06rhIb8F4Zv2VlhgO+XoymjchgtzAAADYtmfD5V26L8GcxHNooIF4
n3KUpnJfSBIUUoonz8iU6L6JOdhxmB+xdADr39qnbl6t00JjVDV9wVvBk+d63J0Z
CO6KkIkCjIljTxMwXi0k2pcx1HwbHg2UDTkNY5wVimCmpzKCQhwMegVnUMZAFd+l
ex7CW8iXZdc/uSObYdC67IvpDPEu9LnDrBQVTqSjjMA4TfqqdJWAKdeOLifeFnOI
e/o3QVRCC7owK7ijyeG5gh4M84ZxI1NA3JlPdtIz23l/ZCX+oL3bo4Kh3N18Qvqv
DopUdo8v5onIeY/xeTP3NYopAy78IgFUdJxdM+qtglhCNIAbiaKsc+VON0czS1oP
zItSOd0e4147LI/UQOPoM6K3EzQzfXRrS5kE8BaAWk7EomcG1/mrruyzGwmgHjBL
IDCOIZOmVuHI9Xb4yogy1VEc0knYye4hgCWvug/K8+RmKEH8hgX3zKy0bWTFOGEt
f2xZWZWjEwRLwoc65PGSnKRiRs968xtJud826Ab/EgZg9sYONDkcvWcgs6WT1eP9
uw3VlXy4edi6liziU0S3F+gp0o7xkvYbl/idM1T/+gUjZBLD6bMpSD/5tDBtqWkK
NOtnZHWkh/cvoPnH+cERSwZUwc48jupoVqWqZ4dF3xN3GJwuD3xk0RBBnHC6dWgy
mQNNA8ICuaBCRGiYpDqZrsFJg88omPj0NRadoTRIWx7fUWFvl7VXnmfTTQHXAaZf
Rmy/us/Db2fbkOC9feWrN9TFSCNW6Oj0Zj8ogTvnBUBQhccQTRafP1VzvlZHaSEy
w7jNb2Igv28ZNBLNEVJct3gPAKkfSWAsiePdHQgGZsr7HfgNWOc3liDurG35y5ew
DrnihdeRr+esMzz0HWD1pNvXubfyMvOAZKVvQ5aLbnYApelKjHrhCLAgV27LCwyI
boR5Wz9FCbtWw1eMC74Z7GZphDV/y0tQonpShiT03YauqBxbiVCEDfN2BvKh5HOG
DWlUkiCYMMDoqpL1O9KHGA2/fwZ+0aQ+NTNXHZamiu0ej4Z6wfAwEq6H0Kroq/p0
GwEJjlEkHZn+rd6B4gS+uLuOWZjPVXZpDUR0XORWOPaRIu4ARNN+uLNaft5MTALi
V/09itpmGentkwh0kh5I7rpQ2Pka31CDX5YUNiq/ku2BSnsWwp6UFc6246DWpQMC
kT2jrt8LaWjEVMyLWcGMYobRZ3uyp0lPkB4gKaeaBuE+AwBnQMHnDY5rR760NXzf
oUvmKJPClZcTkVwOuXx+C8AnzAMbaT1SQGyckwGt9qAYeBD1vI39pMK0+LAr0dpC
ZqbvZ38ZXrYv+dqZ5MuiNWiKCLZWuSHqD8brU+5l+iZthua6heFGj7SPXc1z/SI3
K3e7MuuGzCBwQ7jPtymBeaVXazVzfkq4M5757OXhyhyWaRZexV92DSBCw5Q1d47K
Xd93OHRQ8oAOo+AAEb9tw13eSQQigXueNQEf+lfHG5wioEVSZqNOob9WApX6sbTp
`protect END_PROTECTED
