`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjz8VjzrZYmXC98lW2IBSIxpkLYAAOuaaUUTk/TNuKcxh/ppCpnp41t2f9Z7uwRA
dwnl9aRH+VKprnb8PPnlaogey12M3OqLmNq8S7F4r45wgabQkoKhfXtK/ZKG1vKO
6YVcWg3693Xy46DiZyDTxVcHjRdLfZj7y2109V+HORxCZoDcrRt4qEBES/uKmigK
zt6OwZG1oqEf2/vdCIg2sSUo5W3m6BgeQXFQm6eLMsGCTOrU7y/m/SiQaFzQRKog
nKwAeartYGFlY4XMh+O15siPtpg5ZPspvLlbKoEwdHySHAEWRywg+ntxC9SOy3aQ
g6apaQFSaEyTe2gvH1skCcKf6y1UvvS8UHSVxMCh2E5iF6wa++CcYelEUq2pxgrA
nOdF/9g/+ZzO7z1v62PcAsn/dIA3hTYtHjceEqgM1nlAMBEjAieHT8UtHqhaeMlf
uGhZ3XsNe8VB7aKTltDVyA==
`protect END_PROTECTED
