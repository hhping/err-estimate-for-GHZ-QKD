`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Em7hLTV5SqVFkJc7N8RSvk7tFes9JU9zwl/t1I+JAFdR96r2zHE3IF8opjNoUpQ
bWyHsBJL6lGvLV22kjX1L2V6PGCFgHNgds3z9zpJr1FIopCa5CGvX/+o5FuT8BLJ
42OfobXQPYaRiviruH78z56QdnEuiCQphe0s4CdbGlPLWKNDe48QlqbPiy9tnR5B
LnczkxuCAcyRVphCVt+7o6kI8ASPYTTUJrHDhN9wKxpcyQcQGuailn7u+uBj6QCk
lLa9Nbs9yACijX3ZSx8MmjENwBh9Ul9jr8xC7Zqj3fw3LCs0upC3k0p3HjIExHm9
ZRdbwvvj2cdxz8k2uNamDS3L29qHfXSRY+wQF3bb+qhEwgv8l4MYJXix4Dbeiurl
llogUM0Nya+iFyJj808/mjDESAYOkU1iibWG1KnU+OXCTv0IYYAz4ZG79Jqw3dNb
aQF8b0A+NDAxMwZJdRwxnw9avWEvbJEe5RWMwR/qHM/iSXajyyMYnF37hJyTpmW6
YKay3Ei3MASvAij5vz+Rcf3ArUDYjCN7ZEHWFj0xMWcIJeG/BQu12gCPv7Rd0Myg
aL+SDLBwgv2HI9mmX5Cm8vYIdWlp/6ZyRziYaT1YPSSLk8gY8vFbIIbDHyrGUez6
Cvf4L8P7csp4TMsU5oxy/eePqn1HlPYTezr4dEG18wd42IpkRd+afS/dpSjXI8Qb
83SoLJeMM+uTdApg1Iu/4AdaLLatfJIohwnXehAmSZxxdG54kUixrM5+3AIf4+rj
CaaNkc8sZyThQfmDDo1yUQrL7E5ACD+64KzNTVEFgtFQya/cJsB3O3cBgoGtnUBP
zLplPoLzFiT70YQss1WA/5D3r4E+JL0ReseS7yzr86aByzaaOfGtDN2XTcEDv4S8
IeMY0oZl/+YVkWn9dWmsEgB3zBmtzLbe3vrl2wGETNCuui5/h6Iq7hkA3zvGglBc
TLy3JtvgpKWeH9OIAAx1ipXvsi6FjyhU+XQEaMx1fIBOvoN3EMMQkC3R25evH7qb
pAxy6YrzWlH/I385wEAE+8ebGss9NpIRtJiTP0DqrBNSphGlk0a/0xBA/DqM4i1H
4di4TSydQuzURyuYT9LU3r/SRfDxFX6rlkXA8XK0fOS0zoYqEOY8bIh1qYBlMROq
Zth6DB4/SDRrVuQYHr3vWt4b2OxmuCk2m8dIBapjn43fxRyZk5Z/3EA3VOGpycGM
xmjW/Z+nKajE7k4Pu9MfqlVGMFZ3dvIwa0PnkXB1yWas6ZksnwI64GpkWiXUN1vH
s0t+6w+OHofhhb1MduSvmfv4it7PWt4WweQsqHwpBuHxba3rp4Fhl/sCMH3g5bmx
pa22Mt2EyLTf/VjGyI8MQKdYARIfhJiVA3HpVXipC8w1DrGQpXwhcBslNx6QBEY5
Gy+/QAPtFcfue+n4vbvIsggLOWan7NsZ6jJRT4pXxB7bGLwtAMBot2f94Inxka7N
UOrXaFhtEQQrxCl4ymsS7d2zUi5Czzd9K9Pday9gABSsQYjy6g0Ka3/MMBLRhsTe
74bgc61tOLGXHNNApRnADlJubDrCesZ2tvgfSmh028YDC89SZItoNX02ZXqO8f3O
2CIRGMBFqQRaF9RFCtoc3eGZXPK49xGHkTAwmZOdljWi41lmo3+sNiKHM2LgJqh2
2zfN4CN64yUw5FgaaSCoEIVHazvnzESk09B//+UQLKnoQQ62Szu4/mIZMH1FE2uL
RH26AQUc1HYGjpICVLib31iZb3hz70hYQiZGW9AtlrndMfHXW6/q9VMYkxOciKaH
4QLXF/ejo8v7mN3zm6QdMKYZ1ZRAqrAg6w5pwqn3DoYxV7tfhFBtSrBvhTCw/BsI
QR8emS5gC+HCcOJSMMuukr628s6pYSsLrrkabNNUeTbR/bN1QnDBGvADzlmoUpNP
jT2l7O2mItJlbo/vPOo6N0FPhUtsxIt8KuKb824YwGG/B6sncQTEA9m4/PThbG54
8NzF/yecqtGBxlnMXdXCz0AWlWTSH5PzxSXkBKlbBQN8U/qgUD5zI1wYOdPsH5uT
mM+MH+LwiXjTfTohypATpjyo5G/RHA5ppyDTkovRH9CoLp/OMOplDoqvSw6KG5mu
EfpV7s9eJW0ewkEQwB+/k5MSnjZjP8V0jPrUGel1LP8XrWcf/so46W+e1a1W8zji
dRngBrZbjOQH+Kucyz+H3CZf772JGKu9WLzVg4oJPSqP24EBNW4RLxzYFI0tORwE
8Y1Esx1uB9wZ2o9VjoBSU1DJ4Fg3CKogGUf/kec+U3VssQq0O5qVBR10P45mA2FL
eClkK6LsIUvUk9mgiTm45II84ezNwX6x/Ci7nFK7BKPxnhZ3Oz+rUiOGFt77kyR+
A8ubRNNnMf6IRckWShrVM0/Xtzh1LSQwSDqm1jzCOTu0TEGvWr04DmaCsa+s96Dq
vh6bfxb1cgvZzHTk4Tmk/bcZf+eOV89WB3cmWlVE3RQf2JNKnDunvSlRZTGaCWJL
rVVoqU+Tr+RzeJpbd4QYgoutXz49MEze8rxDhnJIjIhiCZhEraGIrCvxIGME9E9K
usyz6GbLvjeRHI1Fk7Oh5n+vS71GsYio5XUntmpY//fkATpUC4nXrek8J9RbwMSk
GQMw/aOpgPam/C+Hhsj0sU6TItbpX2JoiqmjHgv5GDeCz6obkASN+GmkFnedGczZ
I9kOYeLMXkvdLeIFpqK59Ff2B8AiVVEJrQy2gm6U5ULNzUQPihwDY1RNsO0QKRJP
g5e+vtmjyGo4GRZ0MeT0A7MEU8BB3EL1O2RLcjdT3TiKLPqFPRAm46L9GnlB+wsf
nAEbXaJk/g+6T6HzF1r+VzOyfsmWks9l/gaOIWwexl7TNcuyzICKDIevF58Pcalh
R4hnrpOy4IfMPFZPvWGH8lmBQp6yKu816vgs/4NhmDWc4wS0npMe9g7aqZPVHIsD
jAVOVwxbhGoqLmEvdJKX5+8iZCzpE8iH9zsm63glrPrFlUWZIm+7zwak8TnWH02E
xcwrIVIfHWLAlAURWwkcxIx0Pn+S0ngQnYBdg5s4MImzm4DtN5tCjf7EXtzHHenf
Skx1c1AQG7uhc+nM9h43GkDft6xWcGMJVEpPAsDwu6xds5KZYByKLMvPWGE8mh2y
LEP8x9uoAWxTbiEqVMnhnftLvP69AVarZPb2sXD1fLHvsPU6q99ACtHbi5O4qEDW
P6Y7zpcC8iuxe4Rz96CRSDBOgrR9rhwuNdZX2yw3KaYe97DPyZO5Z2nummSTu2R9
KgjewvF5xZ5WEsagjztNeQuhSxanP1S9aY3+FN5mC/PHPo82OWS2tfX5+1pMwyBs
T9wNYpTIXkdBUBNWD0ezKHUOzW4N27ZVh+Y8nx8kIoAqK9FwZfHbzhqow3D7UWWJ
x+WgM0hQr1T1fiWPOTnKdOy3CmB990VehQz2IG5E3D13B2XDs648yIzBRQWtfsDx
Foxhii0Fww2Brl9HiV997g8li43idgqim6tm6U5P29LeYdGBDDoTq4OhTVbLEbgG
QbV1O1Vv/mYkVIjrYvW/sOwz0NL2GL5aApjRw4RmhSJMfj8oK6XruhEV9H3QDAQ/
eZpXhDyjmRpKMjtLwm/uTVwRToQVUOu/+KDFZLbFGBREjwDzVtj70Vo7jJKDEi93
0McDPD1M7GmZqYaQxTodVOom3tlDK/J/9eyLxHijRm8ePIvzrkAP78PgOG9FqdVA
sGrZ93KLOsc6/0qm+iM2h4YcHpI6Ah5JtkCoCdcIXTpCfY82KbHii9YqVYv2WJjD
QVETsWKsLAjZhaaZ/s5M3XSVwY1QARlF7jmBYvcxiB2tFQ1lcx/L4rV9VtjI1c7v
eoIKMXguE6QGJlMEB2/5jzcNoNO0pjAzHyy7BdYxsCEF/CkSvfMbZvw1yfw9ojTg
FUjULodSYPqb2l2GtIl+onzuAAUD4cSBe+5/5mwLL7QEH94NPXYrq124rG94saHD
1aBXOqGJtWmeD0tHJef+gDHGXUfzVogStm9zKzbNjoxjnuUQIqZrIgkMP8hSZMeA
z/p/Nj1Eza+NlBKDodz51Ffgg1nLv0EJ7gBNcdH2z5KBbJZp/PbMTeGKgfghNeJi
CXKBRs3KEdprotsWM1z75Qv8ncvLFb3O63O35mgKSBU4tsRmMAtZSvkF2rYbXpI/
JtGovgM7RJWoPI4I7LfDvjyYIxv0hbKyNH9NZSdv0DOuN/Nu4A123abkRy1s/eDC
2nYKu4J7UB/smbZZsIL4t4/U6TVTKgnEq3rYzKVmnLNBd4nk9HiLNKg7P8EkMr1v
kokzD5V5mE7/vwFEaI3BosuUP3SwQdkSCS/c71OYdFVYU+auX4snX6ZWbHAhN6gv
QKDa/y9Z+Ll67zp+qNpgBFQMNssQG2XtsxTLyFG9GMX3XV5iWV1IUkdyBHPlVOXw
Z6QORZ31fZ7m8QSKC5Pv6BsYcmrvmKdG6x8P4dDQMBO4k/4v82X7pQNhjn8WDHVY
92dpok5Sz5OChMgKDJUrUJKvzDeZvjVIBaWMcIHKz+2oQH9M5pvzKeSA5pD23Knf
7GGAclDiUTRo0uKLUkDEAVgZr6hBWT8bhCKGbvo6l0gP2ZuiRJy9CoepVHbAu717
ZFMRQgPaJDtZUoQHkQq/qfw9N1GTMOP4OVJ73Ehjk/16JLl+ntbbTu4wIcG+z9Z3
lG9HExRWmhiV6oO4uR/85/+n4ICDSf/Yj7PdUMv2RCSRaqH+Ed5yQqTqUW0zO3Yj
TZdJLXYXwQnlr9jXVaGXvoQSZQdFpPCysl22hXnkpVG5oZMk8P82/iUiG9J0ozWA
9Ft/N4mbNTWQ7A5/Wn1ZhiWpjmT1Tx9XP/UQsDyAS2nx65ou1bi5aMmWFnovbSt9
DKhCCeVRX1Zt2pL3xIZycN3GeYEcWv2Hg3BeJhsJYV6vWuSQzoUaZxPYBfE2M/DX
6KUDviM2xbyrDBOWyZ1Pe40eD2U6R22Tx4UNIfdmKgaTtIw07xmThKhBfzjPbxHm
QAq/iROyKxYOD/s/FUBWnFthKB+8mCXB/NygViJGKjPw3cRVhyDAIZbIKrlwuuPm
OgZyxxqLYj085FtW+uwKCiLxP3HipsJw8/HfXr72OO55AucK8IfnNCwSSTff0t9a
0f+rpMuIAG5xJ30TnjSjgg3axD5rorW/YNPRCAFsoiKvEOOOvrhhEIPJhLs8CALZ
1U7hMOj8nut0PQqkL52usVaHtBOF3lN62wEQkKb594IIihs4iwL8/LAOKMnLY7YX
+7LgJArTmKFGEbCFPTLcttRYTOX7czeN2CUUfjPNSLJo45PTLFXnZcrz5TbkAqyC
c+RAL4ZIuOWmTjf8yp3of43+xgLJXywi8/iHNG0fqoZXlfUV8BCGXWM69B3ol48i
oNEwI9c3Y30QbKS/jRtJ1VSCCKBF647jtBw9tgj+sNvoIta981wF1deCtLQ4174Q
QrDFbC2qum6ShHJVt+qw7xw8SudIMheZu7YG0lPhJotI/gIxGoUOvhBiaXqP9+8d
TEzZo/Xmg57Qj9OtjrnWBDgM1gCpaJwgGSNi17zK57GoKYv9Gk8ETOs79X8rrbiM
tKKhIuXCuDgGk4lguSwLxd3vndXV5wyuk5OCFRsshEoHH84VKXOrxvD6ga8IVxzq
EiB3FYCKK/P0LPlCqxDBMGT/mDl7RrDHuh9jDSYOvPGGLZNWnpvvAebQoqkuwmAY
5NU1Rh+mPnf3DKEOUFWW8KC+WiIjimTKDEwbJevuAoYuFYebcy9hGBmvlUBwtS6f
Aj/kygjG/Um1M1KoYT2o+jBOZ6KuyLj0Q6FRKTrcmdKAZw6EPPcZPpTG0YwVcyTy
hgQ0qm50Pyc735a3GhxBk7qnKYzvvQVpxQrKZBwl5ysCR4U2RY7YEQewKctAW4Hb
h1h7RFobld+DuzwqwDtOy3B2QlTbNDuDCxveKcbccLcFudDsasx1zCIJKCNiXEiq
wp4V0kUCIZIZdjOYojvnwXvukEL+ZGJsMBlWUpgscaMLHRiqqWTWPgqFCaIZkpjR
`protect END_PROTECTED
