`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efOM5cQy9SI2Ns1NkWlo5vzfwidxe63qinbsRLNsnq7ZrpViRt9vTPWVDNuNeIGL
PE4DDLeRQGyLhOQfgGvna6pv74agp09V7ztl+ezm9+QY/SIjcooQUqbP2HCnAdyl
ilkhl8TjvObVe3VGNHmWlAXbfnZefjRFWBachMKrfH9UQu5qEtE3YgIhn+/S+gJW
UJYds6C+Kc5vemL4Br2uj3NNZnXy9hPUt1PUHRY2bK+XnN8pqCEHkwUJhz7t4Upu
QRE5VIwH/6bYnImAnqkDp2JzXaOfI7yhHgg3Fa2nspbbGeIOYlzHyqry/6Twcb3Z
tN3pBRzpXEIf6x5L/1tgUkwXtJjtg9hXFls9+vWATHOMD2Z0YzwBxQE8P/oCwATZ
N53rS9wZyBRilRIbaRr+QhoE75TH5JooffJ3wxQAKSYPWt8Cz2b6HjlPRfgrqH8P
SZ9VWAZuAUQAqN5wO1aOWZCGJj3C2ejmBH1p+C9TXuEetYrdSG6phe0vDHjO0Evl
QJN6d4UQ/UUBTDCCPKpCaGW0LFylpxI+LYBs6TeydcyqIE+8aPGYljZTfv0AaGCi
79ZI+zZZ0Sk/NZOR8soNSOObr8eLpdY+75HMRwdu1RBfeCPhiPPYVFmi4RCf0jjx
yyVHz3bwLlakkSnKZI5TDQQx+5tsyprSmvTalxt0O4oH+IoyGjrtqvn0M+5DobGr
z91sEaVRpXRImrbilKsFl2+6Sr34t94A5XrpddokYAfFaYsI1Li53OFBcgzdHRVK
/VGnhCJcTr/7Gd3mZR+Cbv1ciP/UDP8grpdpXylrACi98UpohXOzs6p0kHAGiJBg
s4LUVGh6lFKdtuwJ+YFIxWwm8xovLWjd0UrE62G1wMt2uPy6Y7JDbQj12/ndWerT
9mV9iZipR5rJasP1SpoWgUE3jgUXafQcjoClaCjEhkVNFLYEqhKoiZD5YayEcFtJ
KmE+JMPy1/szXiv4mkDLSK2+DdSr+aNrgsd0unXsj85rg/pppTIbTY7aqKNJCpNL
SrubKeGtVxonmScA+Tug+hrJFVp7jJOij3BaMA7xAnHt4c9BGL/kSerhPoRVQCKw
cAABP4Ath5t1euexPseg+TsMwVGcANnveY2sFNP+AbkuVKqs3MBBU6UVEORSMN5R
XUvdnsTT+P9SJ6l0yzvN+xotKFmYwF7B5FvzJCZnKXoXGFPVGHSsfNFzHjSwC4uz
b/KwY78sBPHTTp3p9vPfYulIGEyO3QrAzLX4aTWXG0VJu0Ootfpo5ZSJbzFJzHuj
FkmxFcb1FbVt41nBCmXSe9qGJ6e1xyG4whp3+80HUzoZc1ZkAz3QyZHmF3zHbFp/
RmtuQttr7O4RqMG5wHkx1LayL2bTIDB5WssxSVDC/FESSofRtreAHKLsm2ZxUSFl
LdlakIEAcpmO2Lg5d4g4Ol2aNM8GDfDESwgFQKoJV0g=
`protect END_PROTECTED
