`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I80nJWsWsBk4abjRfEKpvmeaJskh/KnULqeuDlr+yJhJXuDyDz1EMjWrayWhi0Ph
EFwdRoQupPxXnO+oenAiUHR23qqrrCoqXCMVQyW8LolIuemvf0CSErb1Q0BtfoRZ
C2nNfpJXv0e46qQ/Sx+O/f9SS9xAaNGeuvQRRpyeEtG6B+kZ+FdpooUu+v3O+Ly1
eI+55hmUNZyGELqI2SZg1DUGSUOHJbzn813f0Sn8RB4tnVuKI40fq/V1RX7bUSXj
TnVgj1zhd8+VqAAnequIqPGSHoth/f/OAJ3ahmozMw1ksWd8cgBdaOgG4yy+hgCg
KCkecesoTuQerv5P44iBJEZkCEGuz0G72YPqeuHz7zIQ9fAKxPrdolRVi1EzCoK5
D5BBIg+bln04Ruqufv/k9VMxrF7GsChvKIRXYrbQ8Q6rlUblFqIr8JdbciMAj+pL
yOPjEBIhKHcfJr/CQ8ZNHGZvEDsycJVuMu/XR7ufbKcLY773tHKSGnEPPAbiWpZY
gj0g7uezshZ4J+997Kx62Lky2FGcYRf+Y+8NHRmIy8cgyIxU/t6FnUT7g7Rd0WmY
dg/dWfILW3tl2Qb21u83oyjSLejWggGuz29OJFs58o3kzXoAHqUTVD+R1T5nCq3E
G0mMGc2WBl0iDb5YP1ByZtxgyycNQmC/e1Cq/k8h9t9wx0MbC84nk9Fa13HJeeZw
MUUpTp/xA3xM6tIt8Umes2zQxjNiq1tkNaFQghnoWO+hyKHyIHpsu6IadI7CGL6S
uxkhZYTWuMhSzEl770igzRZbWGwSli9uFQc6vfEhFmbGpCnY+NMVPqc8yAlDcML1
2KzqBuCrG57WR1B8RpNOwfwfuiyBKi4zFP9ihxvrnd47ZNLEJ6RKduKa/i3n3dEd
PiZLfpIAl/bAX2H8k4QJ+plIQ09E0a83UoXAhyZmu32k9aMM2neat+8B9tAtOCEr
LNVhENp5ljITJqalbgpplIAEmXys5uk8/+SIuR87LHTORR8/+GsKrZpEysoUIeDN
gJGQQYkUHVgy1F2SMR8klnnjrFMnrggk4PGIV4y/3ZbS9wBvKQApo4gUqd1CXV+h
yiEfUa0sv7e8XVOs7D45qRAaLZa7W94VnBWPyI0g1WjMAjzL0ZJGHAfzOw68Lm8y
G2GyZfVdYPyIF1BXd/+DwZB8WT9C5GJIUJG28XfdW2QSE68TTQgKg9FkGUX6Ulkx
asdlNa8Sj9PKzXuN2BVSDNIOpQM5B2SkGyYmioqJOpsgXfn+tBnrHqRdpMClSdpg
hSnO4w2ZUiDuyf/TaKDEMRG1PFlC3PtgRxObpNANbZHLx2Ml8zI8tbNCXkfhAKU3
ZucHFbW4pASLjYxNOnt1BJ3IhTH2rlHewUz9JDaEyI827UES9sDDRmtmT6uJpbrH
LJCabMX0v/yqOG2/BAnJBBPuWaRvpfudKPUZDHbb0J6ckECNYHslZ43oDgQWlho1
aFTcJHW10091yWYbjG6Jj/5KyWWbanHw8CH7fHolRNt5BMW7CfsQPmKe9pRmVts1
cS6DCHbbvc8n0mtBpQQZ2coc14vYFpwQDDVU7c7meArUnDntD4wsDr3qr8fJex6l
P4fBf9VR2r42U/HFu75r0K2TQ2KRpHpgy11oW3gJjlk7kdteJpH0fwGhzYNyQ+AJ
MuIZcp1tG79i8qlAbKFcAg4rxdVo9dvzVL8ymVgO9OGg/F5F7hEaTzdMfaXpGAt4
okV9xKjUurRmGddP/y6/kT2z/Ptac1evkF4pu6ZW/lFt0OWJaNyFYTAFdvW+37Az
ob8VtI1LNSNs3OhehuO3vhN3TKd+K7f+BPvSm8MpLI59a0OUrRogOwc808N1x78H
9Ekgaq2nWgcdS2CfVYWQRg==
`protect END_PROTECTED
