`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
orySkNGcNYP3/0vLEYH1ylkPFSV+0fLY4qDunQ9iuuTE6Tv0qv2FeJXC8wh0fDle
CK9aoyvqW5SF0Q6YJUnPa1uB3Xoegy0V5VZaIyK9PeTORC3zqh72+SzAlZ9rR5dT
EzzNMCsN/sFbzC2hUwgFQP80ip8/gFp9iIlqkxIXhhBBESwbrkyUTjE+Nib7TLXV
c1z5DHl//x9JKK+HUucSlLBxuzFfwbJZ8yWvm8lbHayvG/DkKKyBZkH1BUwl1+PB
XxOBGsQbj1YDGk4GEAAKctXPJfQ7AbbAhxjnGaEzLayzIvunyrzP9ZySvUw6Qvqi
q/XbJc6KbwrzJbRcxOj1SvEL+FKHBxmRkwR2cQf3ZiY7Hr6qhxkpiflTazoFDM/D
nowwnoQLW07jmvTeQMfYSBsg0AkeU273xZ8k/BSxWvu+vhem+e34+94dWE5OVpNf
wXFz8MeWO8YJ0OZ7KiuE601J2mzUGQuw1GL3+3EOsyjt8yzCN09u+RzFvOx2vVr7
p8/THtwb80BSEJEQILv6GuOwI2yvRX/sJCUsB0Sm5uT/lgL0/3QbGsDREkydVzoP
pZgWFWxlIO44t5A0WWPqm0eCOHWlFWclcHnK586VnNA6iyXysDrOqM8pBnijWRVZ
m9P3VTXgA0ekm5VjhM8Yw5AjXsYYf1Qqck3f+ez2n8FoKfQqyn6lZ5h5d95cvtdh
KLZRg+C7fm1T5RUlPrGlxblziR/G+QqUBLZNo8NI8TUTXBwnd/EsZSKRTutqGj6V
sVy+7y7HbuQo38+cSHesZ3LWpa+lFCQstMu/XIKnicTIR0NCcgcr+894BIi3kO2l
F3fSt23R1XAAVhQFdjBIflS5+ypwDd5UXDv323gccSemWI7XqhW/LcgoUcYFNFLh
36c3IbIq90O0HbWAh/b3++nhCbMZTA1Ci6RS0fjNjUCmBL3rllH/lbsyRTZzXY6Y
pFIw69b/pjC9ChvpgFojGFWQMcyAosghaZGnuJlnX6bKSx+hG8DTCtjBmZ+6H+3J
Pk7BcOw0NloHy8fnplK5i5rzAge/6flYdTqgDBeAe6mMPS68ezjdTifG9twbdAK1
hbqNuUFzGQ9itcj9HQcD6Ef1ezl8VCsFJ0VhuX2F6DzewNWdniyYJ+CwoCUTqdGH
lcCpdeS0c2P7wGy1dFEmqSJF6EINlkXFDq8YdgZ6XTRdLH21HHHmVwZDUSD0Jc87
m2C1odK9z+ksiKPT84J8B85S07j5WnRv/5leHzvGboUJFLlQj/BHawZIwNseZwU3
G8wHFu3p9RoQZ1TS3nV8pgOMtu1LyfTiPrsHq6mwivzEfYmp4nRMCZF4agHr0iPC
bMG+hj+Mtp8cikIaIu3kT+I7taxZi1eJ7cor7cmqp8JvGLpRS7s/R13BmTBpakhq
Lon+MPMJL15DYO3Duux6Hooky98dBDkGX3q0X6+I2j9gFPCQK1zcywBpWTY9Zgyp
dyoPeW6IL2d9ySjYHz0YGKyQLANTlbFUR+ijuWVEtidSre2BDne013HnXZJ+ZAIj
`protect END_PROTECTED
