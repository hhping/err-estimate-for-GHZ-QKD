`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y26FRbYJlQXPnjd6PcfAOmplldOo7v+HeIunU6+XdF1zGR0QZq44o/iLBcgJgnDH
YDxfJjQvvGDAtyzJ252+6zozJKkXH8YjCeRoZ83ORUbVIwc+4cRlZeZ7BjhSQJH0
9ozwLgWmPQA9hffxIO50CzNYME/4yqh4jdP9TAdFoSGzxWzk4U0ImmzO3l9tGRa0
d6IK+weUkjqX/X9g8+h1aA6WGkXPLy0oJ+plT/kNnI/SR6vo4p9RicTapXkfarnU
BVKAekyU+DSaORcj01oIn0qcGBFL8UgM28HxyqvhqZqPRXF9Q31iWPrCWkFn7NJU
3Neeos2/1OaF/PM6wBhq2edHfJEz/+eSXGwHpqmONvsg3pfs8eqS0pRPNhqnxHNS
HqsTUW9TVCO91sx9KXHjn+b6yD5zAW4R5/5r88UV/l1Nwn6GCXjksJcXFX9TC9Lj
LtYwi7yydTxv09WYn2Eq2UHgW1+u0WpY4XXvSJ+NNg0P24usrWxBgTQKffiClxB8
m5aNA7ScotVslgcS21M7INhNFjRdIcPAgpSX3ueH8toeCyJuVsfLfC+mtepcErk6
FhywnPWaKdn9c2c2YbvO0hZd6/rQa8327tTpmbqJCj1HRkIiRxhp+KPZwvazniHv
TPubAPemqrxYk6/agCk2/MSDSdpHWGHK4OvNhyNypsXbjKaIp7U825vFN5AKI/Vd
1aSKokxMNNXa+x42hVpyDArs+q73HEJgFCkMWe2jaGpTLbN9SKmAFt2+sfiRl/Jn
Qzg0E35ASd64Iv5k3WVff5ixFVvXbjUZ3AHZe18ow5e3xUFg12x1L8Jq9f4M1LTW
ABpxuyepjyIMibOkdkW4/+6kVJfqrQ9XGlH3mdi+f7J5KKff57keXAFFWykgZYVO
kfJOTj+gUDMl/403SEmRAhaB9FiQ9ng3inZtjM1AiGqBrRM99Hw767xNubkoUa2A
jAYM7J+aH+h5ZZRe4YMU/WCDLqnw/u9mqXyX9e2KFbIqUbBjhLsNeM1YkApSpI19
Lf6eG1JGI2SLD6bSG+nw034HDQn7ljg9/oCIVy03A71VQzOASJIATtN31j2GdIxJ
XqA/yu+gdxHmxcCx7UWCYA6eExDeXUaGSiOwntwtA4nkMw1V9U9Yc9dZorYLmJpQ
yV/dBFN5ND6Q58vyoRzK2w==
`protect END_PROTECTED
