`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fp4nf7UK6002Mhtz3gQEk4iGN42dZgX68ZPdSoa5zKmruJHnGDa33Z5DnfkM5DQ
Lg+/brKSRexlRLTwi+LDfBZKBqbheeFVl9Zui3UX9t0NWmMRgPNyz7iSJY5kPawo
Vah9v+JPD1fGAbj6xqkkmVH3votmQVHvFt3TNV0KZkSn3hrRnlc2k3MozYYfBLb7
mN5frM2YjsBxgtKpNnu5zjF+Zxjalw3tYNaxHft1Oi1w0Q4/gCZ17eZxfHV42A56
w3N9uGNFArwKYUMAqfuPwqgZTkTcLEoRl2gwiKzauCYoD4IsQKVnuKKD19gdWRKo
OWdZ4oVgex+Xp/MvRDbWiHzZa4GdN6ROrNBxh/qcwr3EXjIEczPKvNaJK9xWtLjt
uSLvr1kXeG8afc72QiA2WDLyh+uK+CYs1ndfHuVNRtKCoa1qAKYgu1jXHiUm4Fvx
Q2BXSkrH+L/rjCjcVvOaZDcZiqtZncFwjIRcnq0H2TJ+mQ2enPR80GpVtwhwp791
Hv9pLbu11mNIhACIpPXRMQQ9ObS6EJLSU8/U/hZALpmGjkrtpVwTIEleh+l+G2wo
NqMQETYMzm1UPXMJcotdtC1qaHERSEco1ysZzM7aCuw2o0py/oQ3mZMvbDfFr0oy
Q2wxezf/SJunShRp4HJ5w1Ew1HPqjGvY7moFZaVMPBPLQJLTBzWPEsoAGk1I9cAc
UPna3ix4eZ4F3QSJ+OaWwV7MY9mg0jl27PPtjDjaSZrIddvM9/67lpX1sXsbqLhG
tOotKF7RrsbtnCseLuL9qa8uZHthC6CMLHgcMRgDn1HzsB7jOi5AlhTn/qhaXg+4
1sKT14mBQj2j2FAknrYwqGc5pQNKVy4JOuL/RrjkyDalo7Mnfr6/kSQe6qW1lJms
lkrfD/jVuruJXZXLr5dKT/RDstcZhC5AjWaLK2FAFUP0L89bNELohcBZPRasBZHi
kHfMK+wwE94GLqwRu9lay7SJR5M85/ReAv9RfwOVMdy/JcRRJ+AFEKaw15lgYv36
X42BIYdLayKUBDLhDTJStGwBo6BVL3/s/PaYEcCFzS8fJJRTaspLpIutkcKB5R9r
bIo+uUf545gyh+tUYvfsMQyHvY2OgqEVL8ZM5JQLUBp8NhUUO9oa94FhKXoTLT6B
ZD9WGGS8q+jUwKSutqjBQqpQRo6xDsgaSRmp78U/gpQwjrTmvgV9mDvtyIqa6OnP
`protect END_PROTECTED
