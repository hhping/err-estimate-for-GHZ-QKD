`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67UUeHKXZB+B2kXJJxpqvAWAP0fYIEpTJz7MeycY6FU9sT9Nkc50DThUEet3Gxu8
Fx0ftqgA5MORj5VmjgU8b0UIWoxAmX8voUFuSaGbE1MARReSGGn3C9KtxUv3IkIA
V1k226wFdQVpM8IlB6TS45cq6Jku4VNz8HmbOmpQbpfejMTa15iTvrZsexiv7Lqk
FCgE9JzunToWMPJpi05R1d03IAH1MKYKPI71R+LF6yu+TWGbSnQpOKBtd9VJV9jo
AQdtYU5Fj6meQxDB0qqrEGY6ge/3CucuGbGKDqYLD1W9AO2sb+tD9Zx2mJlkiBhG
ltzucoS+DvY76Oo26c7hHNE3yc/aD5uxTEhPyydk5/JzOgP8rd+u+llhvTjYso4f
vwf8webhi/NeQab4hWeAmAu5gqfPEfnu8CGVShfW2cgKd6bwAEo3zlFWK3S4L0P2
pNmPzJoIa0omiXrewYs9d7QlpWqJjf4g9i3GAhrQH7KaX5q1oNMMxH1A1QGS0sZh
onJDFEQICRJ6+uU1t18ctFu1nbDJ8P/GFLsAJUjzIOF2niuYNxIDYtzz4Zw4todE
K4EiWyZ9vY7w0m7784Sk5+hsQjM2+C7CZLMEdastQfY5023FMHmfqhcRL7ONcszz
QymbZbWxsE+vyYd+WzBhQPBrqHRDJ1eJeYBRkYLyh/Q7+nBjIgbdZTsq0KZ3/Ure
9eqfM+h5xgpiqnR5qxazc+blf8SswM4gtH8hPpwbmHrLGDn4+DaehRxNZyemhhvK
L6uolfLc0p/qd4oJKelHOKan/1wW98voQemV77y9DxUSM9L3OMURBCbAoZ+Tcotm
F43HYF0Bk5R/fdIhOSji7AWb9ry370HUyVe5WVRdXtp9i1mFUTm+xcLGvhI7h7aS
tV5ZL1HKGkoDKgIZ2sS1/hvFTgK599jDf9K7A43OrhTa4kH/tOCNURmrhQbdAreV
xam85cgYclMf1/6XzgAWuRt4bHNGtB+MTOvgy8TQ+mY4AD2ru15ICm0lFO9zmpYI
`protect END_PROTECTED
