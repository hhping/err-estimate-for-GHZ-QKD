`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXAraJPO4eyP5As8vwT3dyYzuuCrx2td1ilz/f/JUopdc5HacW2fElFXChPFHKGi
ThIsopvLq2/Lv5aSQMmjjY4rwHxYx5jwCLncRqdclTA6N3w6WshDLTIQATdFFGNU
00+Srt8p67T+JSye/gs+xqN5ptKy9GGhrOGOLog9Iw0gxhiJs8s7G+1D1QUW06rm
EVVWy+ZFSkQWU0h0pvXkdFt9J5+CfITbTWdkbTXU2Gd98ogzu9Da/c9hkvRr8PAe
QZgHGJ2b2ld5ToRG4/gt+ddl6EB4yeGS9TTgbb+EcgQcB/rXzSZZrUcyypG2NgPd
HeX+PvuSujyJK/iitAf+FZO9+TqgHhAeFjOC2qXh1xQ96xQ0i8LDTWXizspbyPyB
/iiQxie5j1K65W/7zAPlQdkEdWx3M+0fBzl7dhNTL5bJvg/Jtde7wM1cdPAYxXch
9UpHeqgfd8QKVcKAYXVUQ/BZJo/Dl0zl7x1kGL9C/p3xt6bmFRBe/882R1f2/D6L
B4BT0GLjfUxLQC4KyaTV0Ob1rbmteNaf2a9Hz2sPye1LOvmxzo6nzUKCSloj5ugs
iix7SJ/Ama1No6z2XyMOU9u5Pi9CPIRkd7bdr0KZFMxvGpN1CtL7E792SAer/1hU
QzbsYoi0E39LyeP6Rn3fhoFBbtq9rF7XbRRXzIEKyeUlmw301yIdeWyvLoqZQqpp
iMDllXv4mV+qOZx9DireiZFeZAP4jrj5GixyqMTiJaouqhNLvs6pIq8sWrxL1u9y
vhu6chmBDCqdZbj7QXuOHeD0/qdi+U0r0wzS+SkiWvhSryzmZgQkf9dpKDeYUqos
qqSsC7tR6+gZmVqyyOl/wjRP7G+7CyK/H/c7CI9XkUfCChuGxmSeWIE5E/QF1UC3
k+NXOZfp7/pqNc51drlKp2EYy+7RFmNn88KrdQMlRhgPEcLQXQvw/LRKP6Jimpti
maAV31bHYOBRCnUhF+1+axyHQ6ewts0GrPucfIKsR509aTwF8NpXsXDsKGjZjutR
ZpsN1x91Se/tNJ0n5Fu/K9ZlrQZoIEErQBoRuq8RZ1dfZrHt9frR6Mlem8Bmlf6v
`protect END_PROTECTED
