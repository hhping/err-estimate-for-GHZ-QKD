`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
en0KfoaJ3Cg3IMrnzm4bbDJ93vlW4drxOEjRGTI73nQCDglvCer/rX8A5I2+tdyg
+MJr+npLSUq9SKJgB19dVETW4GZtex45+kwKtlaczwkMP6A9FaOfiMeN/JQDTlaj
E2vaVXGVe784rXp6RZgMUPflFRRcaFruhhc0Nvz4ifTqTxFKFwtEcjZCjMB5+By6
41+EAhw3WHwf6LOGgvwA+zm4BeuMW+nYby+yf0+FO5vvz486sSHs6iYVt8eSJNtI
K9XqdYZ2J3rKPLawD7le1KNl0FJHPN1OGUJSFD8GDW3ZakoxjrJVH6LjnK9yKfvG
PHWji2vF4NHXAHMP4ZMLTgII/TWl0RBR1fzeiSt/BDs5JA+ZyUdjRC/K6uNxPLpQ
Z6T+Nh9k48RnZzLzFQxt3W4/XeZNKYJjEYNI1PYQ7Pd+aRISx6//0hHHpKTEVPZF
hy1YXMYaD9ArXZ9i6IR6NTlYxj8GE+2VItCvXMKBW1DODe2nbA7f6s1nLBtzEZ3z
MrVYYJeu/X8m8RHvtddtcAufmKFCYI1RjhUDd5OWh4cA0oso7snhWlda47jxJtGQ
7k/rR7f1DLKR0DaH9m+nI05n4moq/syMwCClDkMVrCTDkGp8L23Bmuihmnh0h7Dz
XTkKr5lSd9Scg5X8akI+ySYTbZG109PPo+0rQ2FaxzUfKupBQ0FBZvYyD/7imBGP
Ld2DooP0lwpTRskKlQrmDdSX32PBLcA6+BeTb1ESH1L9Vxjkvl/HyyX1TBa8LEqH
Z6VauivXTTCOhfvNWCmaH+8KGH8LmX91Sxx7Tz59YDNG5FanvyQIpsIXQbIpLZS+
71a2XcPOH2HZXFqnTDUz8+jklr35QJxDKLA0ACHt+2weSMHUg4v3Wg39cJAkIeQV
SDU0MI5VDBLecJ+Rtr4tT1FkxQSKD17kss0Q7b0m2lD22Is97FM5js29DiMBY0wh
SU2raEKsOQzamQvp5EwlR92O9Ap0vF2NCNaWLLu5CgEf4jDcIkUtAMhFXkqrewWn
waH4toyA0mjo/fhr9znV+crA6v+yg8SHrTc7NfcawHjnPS1yyA9lfoLPPsJhhSr5
hHFzwjgXQtuIIpt8xbUhceaoK+qcns0kYbDto1pq7ADLFT/Ukcuza3bBGoL9XUyy
4yqQEo8dfTErajqXABLRz/bt/FaHorcx3kvEyIDpDJLDnUc3hEpjZ+TOo+Brpqsj
VYYNtbNVk+qX/2ktxe1lqMHfpbCoZv7eJiJjP+5T0uxXeYEVYsH2ykv88UWl+8z2
xVMVGkxpaUdLmXHzbEXk6/j5bztREu5oAJEMEDlC6XJQ2BCzFIr4tqg+L1eWBrMg
3cS2DZtxEBjVOkhsJqPme9IjaE8+hk4ZzBhWO3iJgvmjDF/3fFd0lb4MlnhmWsl9
7UwwPZCxD7ulxW8IXz+S6yiS0zFS5G8Z13DTj7wRTVO8XIiYAkM6vp7ZxDN45l6U
awJ7pkUa6uWwkrLX1rTRP9MvtAhDTdkEfanS5ycV2eKlN21KsEY/zMYAGnLJCQz7
jt2B0Ht1PWW02k+ipeGZUkSigKIfMmuvOVEPWe5DrfzfIPQ5ZfWjeZdFWaZbr+5/
DBF+8awseSBbENBE4wKz6iYm6jM64A1q+QB9SHWJP+mUYuVwmDyJY6tl+BhzkQSz
MtKqk4Qt2wvURmD0UMqjwe5tsMTQwJ5JXaaeEPnr98km8kUZ9BfnNSvrI5F9dyWY
julIspJvezafXoOJTaaCk0Bs0fP2lIUFR+aqwq/m/OYupXQcfbjRgKpOpYaNM7nE
HyabcwyGkLxtYvwFiPga2anllk/8XPYiwOV1eagUupK/bhgOSnPcYbtYZEdjH849
De8fRkX2jPabi9XwGWWiy7QpnecYGkTQY3qDoqQvwNF6kQq9H8VR3dhf90CjZ1tm
8LHQ3ZGij734fGqJGoMI1xrVkh4vJM0oEtu9oId2iLpEaCYjZrBvZ+NQ2GYB1xA9
NK4aF5kddLNZDLTqv5+JPNeFPDbciKJmpGRXOLk1V2tR0GZhW96CMW2qGgaSIbXC
OyGpItTzTl92fOu0nDYUfoK6AysOluOwUyJT2x5BVIKc+mqWMGoWluoYgaJuLfOj
`protect END_PROTECTED
