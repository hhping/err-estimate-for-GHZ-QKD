`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vL1Kk5mnbPGCq1efn1b7P/K6iqVFKOz78yQ1xtq8HqtFRHrpxDuM9dqreEwQ2p0O
AnAL/wPqKDF34ESBi/EHExRN0ZaOyPw9NlWOhVow9iFO6B4pvL040lrnryI9NYQQ
kxgt767BIe5MW/cIRPu5rXu2QH7hqFxm6QsxUdqgN9GZlVzpDwsFZNHRSyMq/J3h
muhLAH5RKW1OlKEsBrhkyer4MxQh6p5Y0rUc0/COF3i14vvbDWS7zYJV/7CtdQCd
ygmWqSnfBYIOLcTB2i1lYjd+4y7jYFXB7WGEIO5QQm1xVnMGkOBdW8Ja+U7iGsHk
mSDaw/wn+ry2evQIOQfM0HDxxyWUGJbkcUQCgh+SiBfV4n4p2wEN5u8KnTYkFkqT
Cb+c+H6PRqSSE1ES0E6XyOg9v5OBuhLjuMkKIdYX4jMVMdvqFojCqqABb8vLXJQZ
ZPi/tu4dgajP7ztRSZZKuQUvBxTkFTC8RW/Ds67GUa7iKLj1LfX067TSjPT3qXmb
v1JMfbJ/gnEq0NI440UXR027KGgPV/45AkDOfyQoLv0PV2C0k5Uq3UuD5XVFtdUD
0GVw+dNwAgwGmjll6s8Esg==
`protect END_PROTECTED
