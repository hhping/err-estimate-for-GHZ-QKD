`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8kGPHV1MuVTEpfWR230ZepMT01L6KwgsfGLImFQmbndxI+5u/a+Z+/LBpwSsJWo
5nYQyMAUcxEBh3gsnLHMk1bGTDqtWvtXPWIksipHhzA+oL7dczc+U5xjeFV9iJHI
qhUyK4HH2rWlf4BVMr1SF75GzPrsw/Y/VwKpWxGCfCjXJ0Olltq+F1LyAk98UC2L
itacGaXEle9COxpbXGV+WN6jemM95V2zHNTvCjGooI6zMWbVO6b10SwHisAu70Kt
DRPN5CkqevhRGeM8Okz5fWb+OnBXLhx8DsVneOSQcc6WO34ckfSikozuRW7kiGmb
E6U2R1z3cX8SP5H4UV3IxTnibKTfQxgwWzJt4DebEZ4Z2Oc5vAVoSP8IL9oWzAjq
bwFAWwau12ls1p6jNwaUy8phBtS9kok5Y2tAh74J7pwAucpKvYb1Xx8x7IdOmYO4
7Yfd3v5H6wojLMGrU7W/KakY8oKGpB8/r0amPUCD9O3wXrxwB7TRbDVYJHlHOMap
++6SthIlsgv6u6mKSwrVbYxSedqNFsCuIFeW3Y7jzuIBQ0aONFGi5yrmvgLTZpi3
tZvC5qqf4FK9owdeRvAZT1gD1uJFqwY/GsxjwWRpGI8AstGST7x5DY/8ydKOsERA
DfwYl9BGkHowtOf4gsYCBflQ3uSca/QmPtMzaGmlBDvDaGHf5A46kFmTVLyOFmSV
o0E+iObgDE3tHrNiEXJ27HrvRQlaWf9ronOS6s+7DFJVJfx+o3jUKbXH4DQZliT8
Aekg9QQkhTaGXwULLxIaXYl06pYkIaH6CB3P1i+gR4YG4q6RsmubPSEWuY7DFDv4
MQpTMYSWu++uW9dspKZ6dMR5G1lrfdQW6udsP2hdGD7tk6nAFgaIoSWlR0zU/cb2
0HRurIn74NtelRc6XhJO6tStcQOqwxKeposhCqJv9uTd9vT4Bk51ZBSU/IrueUU8
kc9TWB1ysj+WNxcLcd0Rs7BBwIMq4624rH6pwKq53tkp3yRcEIZ/vN3ZaiXb/1Jk
G3NI2Ccf7R1924Sm+xtfpTRYdgg+1AEZXo8qCbQOjFHUlv6Hq2AKDwZ1azdVY4cC
o/Nds3lpuogMLvp+we0mGkAdMq9Xw4nqT8MOObBwz5OCtH2M0tJtqgwb7OAEYXEc
JyQ25v+3CmvG1Ah4wSAJNllw1XVpcDzoQCJLhvMjcTeCrzP38epnpysUkSX4Nce9
50tq21Lig3y/n88hlB5OuSFE9bt0CNxj+3N5RtS76TMcw/j0wH6SvdU1/0wEjUFD
zWd8KkgX2b2l1JI675J3G8qHP0h006TGB9cJTCOhaSX8tEoZtq25JQpyZOy2XCRQ
MmRMQas+jXV3BNgQ6wvjxj2nLHZ2/1hEwRXwD6Sfg/JA4b+XstkwVPC0y4d1rFor
4mhDTyuGwdwPUMo1fcexT8pDyIMfPTUYcGCY83zTiDAESEqguKO9VqBhXhWflVGM
3iPfFC8LLcA3R0y3mN7SZTzfcluPE7tYujeKeY8+hPqAIcrfBjroiTQkXO8hVwMG
cgjJXnV3jrtHCO8dWgtEe7dr0AsMFPQhdJ7xpQk4tbdGw9YsEA7VXzjT7C+5tIY4
2YoxY4bnD0fKVmJIEJUeU1+y3b61hcbi68CAsn7JsFJrAr0UxvU1KK5GHntsYvpP
mTI2gGDq7VkZ/lcyni1muwzMfQBpxoJmZUWzCkmcFL08NpEuVL9EoqEjp2g7yIDS
FmOJyyoTMzOHFxsoKA4Qkg==
`protect END_PROTECTED
