`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hfxZXLoxzrH38KCeyCxc3V2irzAWoY2m1j+EsJ8sAhwR8A94dcdvbw9lYwxuZGIt
ZVX1osTUYujePaPfcKP7oZGMcidFDoZWlFqabzUcxrFjrxgjUvnXhSiY9ZD72oGx
MRyrCP9zlP6m5fqL+wcFzVw258tTyGUt/5td67r8u0i9+2Qr8BsKoxki+vDhbbPy
gSQbzEUQZCy7CmD1PV/daeufZ26f4aVjaYrR+t8aZn2InXoY4tVM9dBU/TGnpq6n
PySsW9UDwryg20jtB9jK4Y1eEL1JZcvhtfN/52GbTXGAMIpvNf1ZaD3O99GQuuX3
NjLLFvpFatKUKgrabts9jyVXapI8mNJLddoPu6CuDWOxjIyDHp8zgIr7w3afpx3X
Ar9qZlosu9pNrqF5ZwtbvVPtIHZN1qPoMxiim6ruih9H9hvl1q9u6ArCU/DRZ61q
4tpt2lGyb5tRjHqOTEeRadqFWiR5natIl2l5NqWBA7pqwsPFr+iltE+DsId73kxT
D9mgluj60/2gfo1Ej6xjKdpWMZ1rBbUz149idcKSlXlWWh1/I7JBUlQvy8eRrEMI
bE7xaFc6kLazDPg+ZWozPEMy/c6cN2Aq5cAnTTKtsrHWKBJt+UIW7E49AFViIeQw
LOSVYN2pTqjW0iKUJugDgd1pQfF0duoSuAdmD+GJk9vIIaEq35VirOqaVrhpf6kk
S6rUQ5A+H2tCm6LS9znvfSYAQ0XhoFssrAWXBmijA+oRkdXg+hepTQpkDPin9IQo
/54nHkeCnhabhZkoX0q+Yi4Y24dXBrDGarPpl56SNNvN83sPzRjcwGB3Wj8eXZCg
NVzxI17C+MdaKq+kxiOI3xRirESLg5cVcaH6v5lMtf+CMTHG4wLalJmyTuHLUo27
KZBemOXFb0Lqkbo9YDIkge4JwZ3UJfue2lERGok4MGWhXn7KabCwLBtoetjM6149
weejAnPYAhtsOw2/6xkhm5InY/nRN572gaGH9evmW8vaaLWaRjvpVdHvVar20mtL
KkCj7mURBIjnavAnmmPVeFSpXHu5bz7i02m6SXj1vVhJwcbEgRmW59SgeNyIN24Q
3ZM4DTeNdG9noL2jvosfB1enHxGH1J56vYqtTTofYWDv6kL/lCljJJALpJG0HvIa
+c0JnCN3D050kBsB4OmA9KO43g2AnYAGhcqdOkMoQaONHiurMmh2DYequymyh3TV
jqONLrRL+5eoy3KWZm9ri9118L+a4BQHKCDbTD/zq8kuCpTBDsbHA5QIg5wbK3y0
6nqG06retqb69qLm56SkLH25EmO5tLMnJzjNLjB/UMtxRxJtrm5fC73Tq1p0rmiC
a4lwcwdMpHyDIcbdSD66kl08lUx1pcFF7ftJomeZilCVjtKhpHxLlsGdqDKdCQKT
yx4Xzen4BCYkJMdIGaMUPfQnaYRltceGGAs05DncA77lENakw+PoCzj/aTjXHHQS
CXzqdYb8h/bh1Xh0OlK4ew==
`protect END_PROTECTED
