`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jB322nZ+QTMuSCliHOxilpPeBoGvFxshXtZ/nLMku46jWSWuz/QyiQoLkGiz7Kvf
VeCze3X8hgy2971kAygJvwsBFRWxZKx/MLs89w9SXOuuhfDUOQnORu9bioUUpIjZ
3r+uvGu86J9cHybeDgJ54Jr+7sO4PPzDtVR59Nl3kiYeHo1cGYL/FhX1jV296xLI
rlI4z0aM8/Uga8WMddm/7acP5Rt1cshIkLLAb531AotR3Zj/Ul8mtu5mTswf0Z5j
Q1w9wEDNYgaROd6HRZcSGKFdUSICxC7s955cDOzSbPzSGcEZpWBbpJNBhMbTdLZi
NCTsidwLDOTYqf0KsCJRhA2GtMIRt7kaZK2uib4T+n298b6DwRnJe7PkF5YPPAuA
dx/XwE0OEn4Z09odnyj3U5R0P4f2s7SxkcQOAHVQBS2lAh5YFjqA4/pOQq1gvwsx
tw3gTtvPnPhaeOEnC6YS8RoHbqw+3nGJvk+mu16MZUChVXtpjyz3l+lJEO2L0+bw
ZHUuxCOGPgC7jpu990DQX72737H/V4IkXnG2TfdilJfCt5MODh4LOIc7ApGTA3e0
lGoiZAJVVLpUEnobWTTNrlhL3LeZj0ESdmswaYfVNYwj4jsYqFki2zQBorSoAAsk
hjVYlEU57CoH8IBte+n7npkfNXSMIYt4mN1fNLrgEvC8VkA6CaqpkivgGVabjGEz
Chi35kHchGBoBIccAPWVvDu0FjOtu2Zn4qognB9WbDZTRIP7WH+oOLN/snyjdBzB
bziEyn2nakA/uIRH45HR8BqZ6N99j/adCLNjuV4FiDNgm/IyQUX9zSTNSUmsJMcY
btDLHxK2kxLNKhhXhYJ1z3WiGtFe0G1NI3FQ7kN24eQ87o3Isf6I3pSTfpMSr6BA
LRA06H6RIq8+8qR9eXGVy6ksExV0aa94i0zGp+bfOGpkzqT84Pf5qHNcwygwSQsC
oE+zIDE+Wgs7T/7jgLZOa7Nd9QvP5G+V0NNQffVLNjkCCyOjG6CwFM6w2ZkVJtD4
TaRsTlfp3MimDbM+AzZS4HnihMn8WWd2TWbBWgsT18Xywzj+hw4beATApnS7C9HV
JLAVaLP8+5TCxnYeGl3euUZHkbhGsstaLNqlWyaZQbZV81OOGfohxpLZ5Fa7Oe6k
gG62/+7Z9A26UxQdgE3cUBSpPr0h+onbz9zgSOMIxlmhJ9GNjlqh6HUtkm/5LDfr
x5vbiLYCWQ4Qjobg+bVnbaRxIsD7CDfx4XYDmPQ3iDoV1RH+v6vK8YvNjiTLij+G
bNIHbtmWpQ1RG5MgYDoEgEDHZIsLcvXPziDchRRSivKT4FptDF+dT/TY2uFd1itb
lFKmdph61S9FedC/dPJj7N1QQHAPvhSJKyeoEIdOhT0VsxdF0gLzmX8iq6svEoSX
U31glzOl4g+4VY3JZ3E1Iw==
`protect END_PROTECTED
