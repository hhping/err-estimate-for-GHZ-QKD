`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
12hGbHQq27ZzCP2W+PAKjc0uphyEJdjjk0WNQTyLZhnEV3ALDXbc44uatFX5xvJh
6fk/Y4ty8Rwh52899PE6rVFY7ObsfS0QSbWBgJudfehhRQKtW+/Hr3S9/NTffRJU
sQARL1I001BWceGEbes1/ONa5x99d5rpKKNH/IMNJtFJeuRXfJPV6joSgpkj6Y3e
DfrdXBwiDNVFrr+WFZdA7CrBF8hpTIJcLf82p1D72Lx1Gk1ZjT4zUk0LyrmtYhem
92kF2oERoykebPGgbj4OL3mRy3uRE8cMTA4odvfs3ZRn2kRIHApInQwuMeoofjOb
3E8e0T8aC/jHlIe0XEDVkRQtNv9zXEep3sytHsV+m6wk2PW6top3B5jpsDV1BAIY
zYEuwhY/WXP9OagTazNXv8d7kzy8dp7XRVCUiqsUct/bUqNPJNPvN6A2HtmY1Lpv
fSKIaSV1c9WvzXYks1pJLom/8b8ydvALQ4SMJzUll+FGK300XFCxOKEb9xf1Gt26
vgTaBihcMB5/VQe6TMv3L7PvBSAkcnV0rbkwMjXHjLrErdXNOpoEZnV3nsydcwLh
pZpXAtJAEzcYcBT8JMoMUl0KsOJJDeIXfy3budcktKneKVLVzdUkggkxQzgYPyWP
kkDCQ29rRL/coG2fG151dGi5yUtF7Wm0gvmWAJRF91CVl2llYYZZKh9wMUrZ+qqX
RMZJcljLrU6A34hPABNqS9ZKOZvJVTu8iIE9Bd0OqTHv584ufbUuuqAos+MRoV1P
Mz4rQIWw1DsyYFNBkWJ3Fr11CtZ3LMwVUKwShd5SMQ6cGGX/X3/wCcrl8U+E3M6V
7Xq1enqffrogExZaL8aOeCIHBk7nRx732bRMC6Q2cHku3YFck+DQua4sSW4xUmIJ
5aYCcUlKYUYzIAaw98Y/d2N7if4w2YyvFRp4XFSmBMcurAiVbkzvXHJLEfbi1wHP
xG0RpocY2JXq+vlWdrYQnwvfZyzFbcxaEAGuW/rExYV+pCIEJYCtrndSi5j5/GrY
n6kBqe61DNX8TaIYc3xZILlzyJ1PS/7MkO1erlox272h8LXTKRXXj460c4o26FJv
cq2/LQmrSFHIeuYmy97L9D9KK0+A5DmB5RXHqxySdzFHV0y4zuVSBMmIm961lWHw
grJq1ikgkpL+Ev9K1e+pXwneuQDepAFQa41/y5r4u9d7HVzEkV0ID94dN9VmxCOP
iyHigxLsZN+Q7NuP+qzkfNB21ljRo7UfCKzAkHZZ8tPBMHZiAJ+As9jWEkoyl/+K
MKAOnRi9YRJIv+VjGBUYFYP0JPDCMNSdZ+1Ax0lA6qBkmL8tJCbqntYBl4+6sgOR
FdNIuYt8O7HdDEYKXRvRJo9Nrp0k4Gu+mSFdpEhgHBeHAGCmzGhq2piZqv9VuQ6I
mQvO06oaebJArGA/dlenZw31HtCYEzpA1I+v1C8rQt2fNAVjy2Q+RBTZ6QM+SSfH
xEDJGdsr6uGBgiyovGrTvP2HcXMFTx8Y3sdReTPlfP1H8MY8wtieCrZ/1ao7NvgN
OyAwg7Qv5xVPs5bAMQGh1G6vjL3v4xGWRTLXp3FJaWQrQkMOTyL0adr/SyurIwXO
oAGR2COTH15xQdwmKGuE8XVXtOuTTvbPrNnowZHRItgTtCRWdAHaNFRMCcyT/vaO
4XR7CcHkBD3+n9ngYiOCVqKxxd0cLmsp9zoBT8rL3weOfbYg+1IO22Xfd4KBV7SI
3OUew3ACJLasnILMwdYNSMglhqz4Hnr6y335iCmsW1Bem725Qsx3CUr923tRLxu5
PBNcHgc4TyDlLYX7+GIm8uzuEbUkltwH2Q905DB90SZ6rwNMj2TRZJs+XHdIo6e2
fW2WA0evmEc1UNOudb3YjQqh+lJ3IJxLRV558l9czb9xTaKvEqoZRl41O8Nou6gk
PfQEO0zlc7ootI/SxVHDksMGmkbRwFRAE8UcdOt5uMNEkrNg+uE4tsczTZlKy4xe
C/JHwVEaGrUA8DPA9WXZqLREAllg8u2neIN5bDO8EghHrKpBkeoKifCyRP6Brf1d
uVsujA3uNW5qj+iKYo+aJyvLCKVQu4SryyShbsuHa9Z/R/xpw8KthMMOPsHfxXjY
CD0pPwF69U1vjw90EBpq0xXr0l5j1xMJdkcsc2/7WwSr+HiycWlPJfve7fh1uT11
haAtgdhD/yCyDqZqRA9UlfRzy+pAx9eNiB5AoKC0DzznFTMccZGiEshTpq1PgRs5
8O+t17H9L1DVspf0mVw7AgMyUsVZDgMsVIEk4V6kHedGqb5xTzTdwxhj4z/p2Iik
hoCg8dfuxOOpYSxzfAmo6CS/JQz/C6E8Fdhowgm7uXglEX8ti33rqYjCPlUScPOt
abh68VJ3PCM9SpQOfmthwMpHP/pmtP7JcQpx720mRthQ/bGB8axPkuKmmr28t8MV
+snxtDgV5X7PYXdM5UENtPcB2/Q3XJMtbDgQP2w8MqZm9IIpyy/O+OrpJhh/GIh5
ZobMACZ6yP45KPGjJ51HXYUC0JXxgI930bOtdK2GyJvLB4sa5XwKdScU4ZF1kfes
Umukgxmru24lCjNWbQ8ZY6Vb+tfr4IKuzpCHb7yb17bshxDJ2Mwn5lOiWTz4Bkl3
mYq2UQ6r5PHXKxXoBaQNxjsnU8f2FqQv4aZNMbiNfmaKrjjVecfmIqRMhQ6hrVUc
LijgNbhMJ/8gcwfEUrltRuamT2m3FIYYpqQv3q1hvBhBT+yuGj1p/sFdB5MFvdYT
HvCB+wyOa9dM1ULHsFfKRmySQ7BFTmwpUwjn0ES9oqGowxJsloaGOnbmqFTlA5Ie
2hzAj4P7z2pjk285cXzAwyzfrm1RFvav++7R879Kcr/BTckiAH4C7kbPEFKmuVfY
m+A5j/HSuZwFqSaN5qX8j8Isp2R1I6rhaKwP+h8DJLC2eTuCA6mEmaaTwklEQCdd
Vs2xWe0CocQT3X30nrtwZmc0lB35ZjePitSjnpZF57DCFPFBpmLSVxpHvYg3cjY9
sSVWMXpt3HAp50bBz3fsocbvTDn/FQ7aTaqWogv5VkGz9DykWsBMsz/2hPNDTnn4
EHbvOiLiYww5vBKn7l2k3kt1Xhf85q0AjOJcn9AvxJQTRvcYQwaURG4aCtTFOqza
SWEtv/R+kOBmNHMdTV+9/8naUDV39dFjIfxXSTwwzlsUsVj+QlVKGkqbm9Aicc71
QSo5ECyiMvgZLL3r7p0w6i+wUEYagetrmeJm3p9airyYFbatnPEkJn63z9gIKFDx
1lXvHss91myjm+tNtqQAXBePg8poWbalj9lMN/sSiwdSDflqwMwLrDmMs1eg6D1t
ZJ7biATczPuUdEW8KGJJmeiMRcHF+Nkc/72mzYboB7YaEu9mb24KnlImdQj2q1Eq
Q3bW/fdV6CJEZRirNdCAIfSsqrV6j9tQhKqWcgKxA9HFFV0mPY4chXsNfa0EFLMk
gmz83Ix3sc6zS28ltXDp50VcCpVb03N4yUNnonwh7M6KGm0rjpGz5kHJlNUm9avE
/veI//NUivuMfDhXxaNj7RjiAf9uajWhlkELjYrRCK/fxM+QGE1rL4qVgKjG5sCC
4kEYGH8jz35o5f9c0JUeOvNe0BpzBnOvIZBeb1IGP4/FRL93PfmHCfMCF0wXGYW8
/omfOBWXDxHbB9bqMxBlLDnIjmnxvXDQYRVO7/ZZHdtBgRZTw1Xn1rgXfAATPwlo
/KysMkzqs/FkWS/gDnBUepcKkPQYFhpkqDEDvjW5ZIB5uOD+uh3xv5GdlWYJIUkp
E6HHgqAPpHfS9pBXFVn5qD3QkqIizMCjwmioOIMYx+B/SMUabkAB94PA6uMz5Xsb
0BbPRja2yOue82JMp0mrIFoLkr0FmtAqxZzYyhbNXvqpF8QS9XmG6N+BkN6b03zk
WOnvw6/EUjjkEf80tZKJPPTTYe8yrfVcLihpXC+J/u8N4Yto9Mqqwp0nLEoE11YG
MlzBEWZe0xgg/jNc0mnI1ljzBN+33h9DtQ9sx5zXI+uLiRA5uvzkBsVQCRy4Pmqb
Ipc9AxXE5mSbTShhXawH6vKytmnODPtWx2UZqJoJjxizomJBQLSmyqd+BLKtw0Tk
/6jPMwLpmWs4ItvR5AvPsie8nrhVxbuOV3vxmHzc9cR0jQRFe5yurmgHpYPC8Lhv
izuNeCcMsB/OFz+OoXvkoh/6wvwQNHVokldjkUznVfH1N2CLwzLZmK6TaxxqYPjP
5oaE/YS0OqmqdFcsPhHIv4j87MjzDUtIFTbfByJ80QFjSxqgvzKI9HjhR7Vjelb+
LZK3LExDMAf4eFVwbsr0FT9ad44P/upWC+vljrf44IlFM0D3MiRd6qt/AREHCHq+
BuNHPdZ5wLQLqlmlHEIR0IHExZE9eEIMJ6rie573uoOGCz9e4o/qkhuJn9LqKWMg
GIUfO0CgCHkDMJbYBJy1XDDcF9ci3b8ILmKIxhJ30j8hXPEfcEJSfW5fNC/L43zI
h+8X3OiDxH2KxIPGHrjvaNUIt9PQQQra1wnApNxiXtslmoCZs1oJ77zP/pzQe9oe
i2j/YEKeNY9NGL5XGs1DktmMModM6Le0Fj1Y8Uv+Rxq0PorsF0b1HZs8RJB2IP9F
Q3l7RC3rezGXQVyVtTtaqT+yr4hyMxTJh74B78+S+CXhHMIpOq+ZmVp0IDb2fUd8
vgueLXcn3Vemb5IAgMOv7AmwNL2YlR0/f4MwvTC/7B/zA+k4kpoYiu9iY96i9WYm
74TNWqP7E77ek5p68oFsPuMAvpUVHqdnWsijQm7DZjthjCUjx+t7Wx0fBueCcSGt
bQw70VN15/A9r14RFvpfNNzKgCsze+OnCf2B3FbTA84iiB5dIRiIQdjnLlvQoQVP
dd5XFmd+j3OrwFQQZ9jU2Ks2X9vukcXR/wtLdFVZdmFeylPbTP7GC5KkU0sKh8Mt
g/gKYklpR4uwqXT0IYwvilEpLDYIdULJwH7+6kBzvHexOaKbbXeVWwWy2NE9sB0m
rywYU3ca5BSa4ja+c8atRFfLJSq3s7xXuuoUzoAqDsdiuhBqNu9lUYqLDpL1Srvh
r21DqA7ICljN/YjftDD3SsgA1HD44zMI65rY99G9khRKGGjMvUB5y/3cCQ3a05Rl
gT4xJyPNZk8Wb51HrX6JJHz+zU1iaWBe4ewCAimpOe0=
`protect END_PROTECTED
