`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yc5bQEyKxSeuEW9ofXzvFsItFvaqKObHEm1+bphza5a2TYR1iMsQcIstKIBPmDo
B45FgX+tJZIpz/3dgcESo7iBO8YNaTYnOizRcYbm6lgeWxQfUWeVlNST+jrB8pbR
8dhMuEfOpC78TmgnJbAmDy6s+2mVz3IUVWvnH9yaTNqTMHC4nBWr5aPzUOykO+C9
kIqoF2w/FFJE0Vp/UZ/LsVxuHWxXEEfcfS09vncx3ZiTW4RahgzCr2aDP33UecPu
Xz6CKoaVX+/xrDsaitNzztEkzJtMEbHZ9nvOK4I5JKRJkwZVl3JB9at+RkgnDH7H
/65emnKGhmVvP7T1jTzkw2MMcNd2yu8qdIAd/Oj89X5HzLdvzyvzhhBh6mX0TB62
1UfOTTSFDuDSiiNE7kum5f2Suzgk7phKQc6E/2r8olUd6Jcwns/UZ5sBxD/y58yk
VzsJm6QxNg6x0mrj4VjDxTqp1Ldf3KmQQwz6USLtabqS/L9E4azFbYZyWTzs9DrK
GvoPM8iMs4MSPcrPmOVJdPJA7dh6V+L/KDEBs1SK5ofR7eH0JHU+Gml+RCwzQ30l
QzlO82T3+SCYQVjWo3Vnn4wgKarGtpDBKASIb95kN9NDxJE72IX1rZtPWk6nDC9E
OY75VsbN7Kz6M+47FnWPpBIEkOjcwRGO7O96X+808cngAlD8qJX//Wf1saIeIJyq
33q8PTVvspnmnOXdyaQA4uvNCaQOGvm9HUozegHI5A6TyaBYF1OpLndjsXFxje4K
HJXVrFDv8S3pqWDF/GKZjgcJ6M57fevDWdqAEuYgHxCbJSxoIdT/+h6USK6/OyJ8
KueCCRYA2V1UjyBUJDY0OXRr0JcCEXFQGxMFRg+KfbOQ00IeLRNh1Kkcba7w1fFy
s/0Jri3s75esheMEMoPQ1n8w156eai1ijrA6tF/h0cmdvazgKif82YfOC7p0flz5
vPuq1W5AXHFdnHvMp+Cen3TDdAh0/q73oKWHNUsGfxTzJT5yWbGitea44Sf9+AYw
0ndt8QpjoQxa6rroML2349LKTmHG2bL+M87tI/K9Jwk=
`protect END_PROTECTED
