`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKTk4oYVdVfJ4qGbSdY8RasqnoBShwdmip5kbGBcoNZSUWYlTzD9OWOS8wOcYzK+
CjjXepp2IRM/uW4osAFVAx6GUrzNwN0Gs8dJFmyIY+wWpSNalVi7R23UN+JotGSl
nGmnRNZzH9cCsRyfVAs8xRWk0NBBc0QKXspY1Wur9DtNtA/mR8TkPl/Rf7I9UHtv
MSnwiFDt6+GXM7fq5hLjp+RyD9swrM+AZYA6WyYSHB1PkDv/jhctyCn8+kHdlybi
9g/NttpTunNXDaGAKHKSrOcQbRngkL2KVeIhyCP/+AFiIz5r6lvkk9I+X7Odxfk1
Bg3s7xJI9pTs7O30gQwl0aB7LBYKuCC1knXLLt7ShOAChUoU6843OpTv7zpmhPPp
v2U1ZsarKFsWlW7ajAErsFCg9d7aQhcYE8RiRP8yQlOm5X+d+qkX+bouIchx5AWH
klWkPcd38DNquq1M7gCthsIc3tV7ZtW5z+ca6V+Dfx0X4U6M7pq3nTEW6ZNLMu+p
e34621FXuPOflrjOWMQs6OGLLRNDemt1VQ/fooxIgqit17UyBOxXu3iFitj7CQT3
185iTnOZMoonmWVCxGsQH+rgwIzxxnuTwp8YRnzbU9E2y4TrFmt16I/YX+QMGFFI
nwvm/yIeFauK1WTedyb8KDKGzcs7zvh1cloDkk1YLbouUTUcPh10GY42KLkoS3n8
maQ+CCPouClghmODYKdyxZiNjpC/dAc36gvyn3g4nPSmPVChjMZtnvV0XD8R4ECB
3yLCsh7k0aDF6oUuFUt8+HVPPaEnsGVBlvmcyfk1d1muFWSd1708fJXd2QkE0IRu
nIhHCyqDMU5vVdYSbm3Dkm+M6V7QhUnhJMKrLOAg2DIKn4Voty9mUTPqvcJuWcTC
bHNPbOXkUBgUTpzW+4QZSlFN4wI48V52V4ZRABVZO6OX16BrzvrFVN+cxAF0l6pJ
Rye6g1RpFLoqCKjNX0WL0QMIUjIUQF+/ZZgaqrmpp3Vl80A9Iu5b6wd/jEfi3opZ
lNAuoz5BnYETNRp9OIOmh5fCBp8gSYwnK4wMUf2alJmOSxBKTR2CCpyvzgmP9alf
rtmp7K4tnboP06Ge5w105byRXClhw1esB9Fe0OQ7Eg3l9FTayI6Lb5e38qUO2ySl
nO5IoH7W+AezImvRRStb/75FodH1rumW4+9vUsj6maPk5X7HaATkp1iqRMgOUApq
d5PuvX99eERYTIbRo8DHVEdSMg4RFDOrIv2bvyvZtK1HX2ZEuFiijPa2IHuFK/kY
hPHreV1exCPdEZpLs0tzR4D2kMHmW9dj59Wp6xZPhvxyf2USXp3GSLqK6rs8r5lS
wl1NucnbsrsIM/pdGANoIgyUYw7SEx0TuCk+cKYLcrM8B7k5jYHJ1Iy9hd72UjEE
tYboEZGQRpifwW6oi7Zji2BlJBV9ufqStOlYfNwubieDPcbFfIaIfCc6/6pA1hja
sN1Y3L4fEWu5Gyi1Spzd/y7pnRSfcO8uJcbb0kF9S9t2FOyTgRmBtAnOrDUxGMWh
1Bd7LQfOxFZHSWfB6LDS+EF+4ZQz7hPHN+ShN0LMkxKPfLS56QFfwxCldpfiqv99
CnsysbaajzujNX7sYcAG9ILGO1MhMDZRfMdtteEhibCTIOTQdqYW5ESLZR409kp6
3s9JRB/UwkrjqGUf5TWazzbr1i+ZER9hO73Di8bJTLD19nQsJWbW+tafk38/Co4x
DgihhJQnvJwaxBpF+fHFMS8XQnC98BURJhHZtFVyZAPUkW7x1+7jOkOcMOhcoTu5
sgqh+r00wU7Ql8+cCVnRxiJBy7mFDAoc7qfNuOcVV8Dz1eduK4jg+cWzCqVFNX44
4s9FvTuJ3bw86f9FrgA4IzKpqg2675UKZks69B9mQq9s+GYL9jGKMmKVg98ce9vF
yZ7pY7c1eZ1MYuFirjeKm2aoE5vvca7vIvYjOe6eeY4=
`protect END_PROTECTED
