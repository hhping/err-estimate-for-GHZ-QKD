`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYWxW6px/xwWgDt3PW8ZlIakNxUrBtWAE3+40pNKZ2FAVTh/cXdcS2mRb5+v+owd
2AfMxf0LULzLIbSoWldFKONpZT+JPpC+h3HyR8U+kMKgWAKPyen2YqB9AKSeTUxu
LrDQUJVOCs8gxL8oYJBRj0t++a1BmiEAsbe/7sJz/DpZfSNoRnmnDoOT4rs9xXjj
U7WehIC+cZh1/NOinkafRuwmxSLyk3/V2Aoh8VGnTMZeXFeLz087qRGcmzY9S8pQ
dEv+u1Da45tIqqCK6SolPDikjoc/L3Z9aGsjgvsQSdNtq9dVUivyp6haPY/iHw+w
7kMESyFES79v4tbx6Xl1zYyYsxtHM1032eZsLn4DTMaywo5+JioF/wha9Amd6QqT
EQ5jiuFJJ4I+MDTTKUcgFCNIX5GOBWgpIXe3hWSI78ckgG17tdmaKq5F1GCkqrfJ
rzG9jztna9A/S2kY38TQ4P/bFeaSwyFtPirmU7oBCUOo0hu5o5sLtuWGJbko4fCU
yS7A5nb78+1TUwsk/gCHcQhTidZX/KxSiKriro4qTiFn82fo8CoRPaSKQL6zvjnJ
MErbEDVUpG2WywccFDbHviqcIoWCA2IFIh22BwK/w9r5zTIXk4ZT/y+y0HMm4nbs
FGNNTSvOHu8AiIw8P1Oj7JypzQJBVgQEwCJVP7yTaXI4LWY1bO8MtdpakrAbNDbC
nNWL+6R0xqGq5A+E+jI4i6sIDgJAJpq5LBPw9AbaCJbl9NjfmgA13x3HFIxPh7Ua
CrgVcBMMA9s7DRXDXQjadzFA1w6glyFq4atQeq5KzzqHTIYh2EOkYYg4eE3jBQwq
CR8DVdJ+qPJQv4xTg5ikcQ1JNp+Zd0oi35oN+PHaplw1ct/ps71W+qkSad3m44Hj
3f/TCbnn8LX1kxgFkIOGT8ZkJWtUTSn44clom6DLpn5BbRJKhGvrbluE5FZFu9o3
Jpf4oKBTLf+XoRAbK95KCwI9F5OkWC+TCD8kFa2l6m6a8rDuN7CBROTjZk5r0TV0
5gfyPnIBYGbo2ZSBkv71vKinbczUV8/wApipLs5pEbp2AGkUbh7EB/TujAG3obcs
T9ZQUdZwelaoCms5dYLybStl1FkJI4hlP1j6r1inJysEnCUxBpKip0aQeFIJ35fD
nn95ldAQVqiKQ1zSlpgd0YZgartgy0RAtV9Mwqd6/a0c7Wwc+70uDxirgWCvXnwR
fAkYfUFKFdSYjcIW/t/AFYWJoVxrC3+Hka2yPPrxlUX5QlhKfJjBhECBHgoYsvKB
wr6GNZL05SUiU4WXRtSraQrndc7McGzXJ13NAtSGI4YaI4V5hULdeAluBRKubQUG
IggNNxWmXdlORE4npCCX0W75ePmGCiNkxRhNR/DfgRpWAKIH+8mUi69LJD0g/Fai
wmmMqkuy1DSMRqyPkBkmppJWsFyCVtngbBMgvU8fSMd6g8shEAhGJk1fSODP/zZx
aP/FHAUJxyiCH5tG2EbaZx2pBmkgqORHFs6k+TZ3KhbU7gIQMs1sdrCLnhAr9xJa
hR2Dt+4Lhf8oHKAwinzH7jMYrG49zF+k/Rg1axczRB73R1DSMNnrWERpYw6b+aTo
XF3tLuiFFEjORGu3qsH/hs9j2lxKyX6pBXhS1tWcv3oeh18EQHpRP85hfiUZ2mco
Y8qX6CZgzz1Oa1f2HMzFlSEY96OrrgRcfjgD6y00rnRaO/RXmEfvzL7bje5MwU7W
N9tiZxp+OdYRzuSLnaOlYn18B83mJzKE1SF+kwrbLGA7WxTrG0SchbDF8p+dBh7z
viNsYHIXqCindgUYzn+NhADjaI+MkPyeu9btl8slis75YDAbHtlyssT6dTzFIg5p
FmBw4spMYbrgAyrUdVf2AEChpLbnOMklO+60VuuKbGOCOx8UhLq1lzaeC+RZDIfx
S1QMZ7FDgMKZb1VwN/fxrqGafqDtPUeCVuJcSIBgKT2UGys+DqP7/bZb0n6Y22Ze
e/65kdw6osieGdOAxJST1DJKQ+qNr6gYZ0M7/eDSWn7ypmWaFtYQRxnGsi6Dcolk
9qKUBMgpIJ0yQoSOk4QkSRTFJxFV4AVsCUxs5A1IPJTOsi1Pl1t5CCvZZgFI7733
m/Sr9/U+yAxBXMjyz+VhffuJ2Iwn2BdHUTvui+IIjmo3lCtwizt+E5X5lLnjGEhq
1yVR0QCf+CN7ZhAtt3c+3fwhut8HHf7comY7kVBgUQFDx36e25IO7G0yye3f41UJ
uXgoXnHwjKZSDUV0EPpQKpp8wpqfh/saGr1qW7jX3LgI0A2TZEiY/QpP3eDGAc9G
kVaUrXm9W3WZDoMj7otjpjUqoBdw75QMnpQ0czLNMItE8AnVWKFwItEz2l+oWCxd
ARFrA7C4NymO1CBm9Fvk7IQyGdz6NfGsDClARWv+GoL4BFY5tpzGT5VRoCtQI1Ob
cHR22uA58pumsd/sVcizVN4rdpca7D+pQS2ksEpPj/POYOdMAtV/Mb5th0YgQL6v
tkxfc6kYfAAeFSrc6u1r5FBawybkYo2cPKibLmFNrBfgFvGZSd2uWLoQA//mZVJX
lUDcRlIJ0bqopqY82YqHoXI65DwCUUkFo47gop5tEKYk7CAshU2SLzGnP4YIX0Yt
xBCv6LfmEzXOo4UoAat9sEKjVfTOzzGSHWoeXQtMCQUviJQrWWct07KO39VA/UPn
VkSXMgS3MMYqL+y0uFD2TrJ/48JfcCHxGMXaB+b3gdgV+HaABC5cxViKKKNGDI5i
wF9yytN5BGKmuo3DAqXhwE9OtGLZ8XRPBhxnmko9xV3eeYCZNBE7XYrGWOczBEQA
hT0WYsv2Z1cUr9n3wy6aoG+kjZgmk73vHAeqEweUA5AxgjK7dVbSQhEmdw2wbvFO
QHIEh/uSJ7T50YXyDO44Y8gyWyzmInYgAbAsz7xeV94SzTXyJpACkvITK3l3sjUB
DNtcm/SWwCUodBgXsEKP66cPEne9Y/dnyLc/JGxoFKweZItwmFStqVfXlBkNIZAz
Hs7J9U2+yEp6K2qZxN3p44iN3G5syW0HU/7VwZfmmG6rzLvc47f24PSSmfzcnDir
l8pp7DxclT/u7GMP7bFQzstIY8JbvQxfCGgVtm4DRfQfOKT6TEO1efBECjv5Xfyf
ztVanUjORwQNyUziLdlvWFzt/UN2HT3oyFFTAxeCKSyNAQXaoiLmk2OWn9w73UFI
/LbfyRqj85eBuDyAzbK8SYVrGVqwyRx73Z25wr3qq+naog4rFGESAcy0rr0H0GLj
Bn0jcjuoEm2YQ86Neg554Hk8qVPaZiwTUDZj1zTh+AXWCR2wtZ6ehSYDZRrDSAse
B3knPCHMR/ncZbt928hXoGNYnhIY18x0lUlMIjOntZ0PoM2yFgbTcuu6o17sZTzQ
B+y7Gfd7b9WrtSaaZhOKCwH+pYy57ECWzFQxBw7LZVBIT4E2/Y3Rhj7pK98Q4KGf
FWc8zFKNbZJr+4O//VmPFYuqg8WCKu4dLoJ/4vuKgDSKcmyQIR0wByNImwrc+/ZB
2sxyRCn1r2cEbc/iKCuSdG+rFkdXr6dscrTSUSshRKuQBGQ1Ja7DZU8VChkenD3w
40ItS20EkAovoztMVkBWCmm2BU6QBSV3wP8mkW6QHm+twrUybS9mhpyvEChek8Us
ZySnFBg9oINV+sa7UXsTwENHWipOzn0+l5kmmaS9XIvocTFK2vnGS/JlRg+/6YDB
FrSCBySnMDhbmIVoa1tqbZPqPJDvJujsNtu6kIjyJSy6sH78kplluoJUtwQYP8JU
IftzZ7QRbATxth1v6AJVRAs1aPF/IpGk6bYJNiEYRHXYuke+bsxwSpHpAr9aXY63
ZsAAeJAELWqErwHJB/cD4qqbS0tPJG7pVOD6M2td0xe1y2nAFFkfORxYK+t6yI6V
CeBnTreJJMqlt7FlGZEr07oKS33g2owIjE5+GhkmRcc/Dy83+3eeW1hiMP/LX36w
79t9Uq15I+Dl7w/rSHmzY5f/l9A43c1DAgG5b4X2mhKL48h1ANvsiSd+qXEtfpa1
LpyaNmkHzWXWA2OGfsw/9qVragCwagqWeKZiYrOWyeblssnP8Drgk+6hmO+t8NpM
1VWaXKIgTFlB4PT5Kqxddbdsvljz1BoKSBW36ojhPuOF9VCEn4ZN6uHlTQhKaDC0
5D+a6GNW6Ldlw4oprbEM9HJpDvxHszsKhE6MpV9QAIblu0QPQlrvSFl3uO5hshKx
1A+87wHaQME/yRdeKwtq3NjofkosjoxDGhZi1Bwmo0yu3RtelSp7rNCTKaQLI3pZ
K8+QYqSYB6y++gR5mFDG9k1wEi0LsYX5VmolWndhLVDH6xaf7hE2fhXHlS3Lmo8x
6vGhHuzaSIFh1E/IPxy4GrE7DIRT7kFkMew0C68qQxJ6M0Aeo1TSD2slavzD7Qx5
uDAYe4YE1ZbFrZFGl7pv6Hf4ztU1GWm0nEAdyhaWxvZLdZJUpxOcSgPNo/zRKlLZ
WdrHO/9GhzGp+I1M0S0kyHrd4D69OO84JhvVnapwRDauCXr0hd2+hyf9D9dBpf2J
EyUvOEWcp+EOL1xAmp3ZYB5tNRN0SMBw2NW4zp5PKeseR9kxsY1m1V1um7Kcykax
+MG4hXzhtU4XM3B0rX8ORX5zd0zuYcnVpRbF3jG5YNNG0WV35DX2bUx2LlXO+Jh7
A6QkdMluZscOZq6wc1xp7BwtnGKkRWs4oRXx7qFUsgV28f0Ksr/iN2uZMhWymwtu
oufVEp/vf8Ab9fJQfpbVM7kxXrzvk3mmIGHUhh8mINnCQh+KEzdg2VvueX8OSYbd
pV6dZt2GRo4Lmr4QJ6/CEDQuwmMG3bEbtMX/S9EgZtW1lCMbp5pwk5IA+Pq5uOL0
bk/QSwTmAessCdXXKCbuFsfjULlEyeozGTuDkGdop9c1TAnhwk0QmyHwR4j7fP9x
Mvz/D4onyKTRoT/MfyrweJhwh1wqFwQve8zXPvB9/+DRPFOryyxaC5eIAqJJJ5Rc
ijY9gRGw8rDDAAQL0j07djLcxH+8iSuy81GPV25lexO2Fe00rawZKIBoASedl/vw
fyMHPVsahyXWwDkp8zEgaULZZFX4nDkUbh/b1VRAeDzdpCMzoEaDuseJpRxW5mab
pQz3HFkTPAaWls5kRModq7iinZaas4d3MYbEFRiS5rsFvhzIBBFJeBVwx+4eTD4x
cfnNJWq4H9BS7tIuDRj2xHdjWqC+B++c+XMDhh74O6Is/AvQjzyM5xett/xlrnqx
HYw3s8o4ggMpgNCSpxySNhxE2MOmModEPw5W/1JnbvZ1ey99N6n6g2e0lvLFtma2
f/ggMt+O5yMRmNJcmBp4WqdkBGD/81kFy5mY/CGZs4eKLN8QD+/muNAWqAyK8XJU
sH5eJbHERzjsjen1AHTovcSA5tnkDTZgVEITOVALjXVvThMTJ3izOCVYXMGmD+Io
50+L/vGIPJNYr/xqASF32rUNN27F84eGGU6f2WZGUXdRuV6r43bcKp4Yoqouz/g3
IDXHsUN+Jc/fe/AgnklzrYiiUfA43BSwl7F2bVJ/M56NRzxjPnMmVo06Fu2xqg8/
6Yt60mxt3aeU65FNjWjYPF7QeBL/vR77nvRDzJMOk/wxNhtnw1Kq/atxxbHgMQ7p
QrSt0FfqtA54i6BPJQfC78peh7Mzc/tO13pwnCemmPVzYSFotenlMR0IJknL60cS
tfE9EUlyE5JpoDtiG/JiHY2OsfN5NwPpGp43CbM5CwHJEIoCVU+F8muetwxs0jgO
lH6dg2ARFviLhy+V8NSM4je4sH1rgMVP08vAIiVaEj8w36k8yucGeEk+RuGD+JE8
GWnNkLsjRg1/E2U9ZkzYBz7rJ836/ceIW86w4bDkmn1m+JKuZV/D4HUkuOflK2yE
vBjDrmMhfKmmO9C4ERps+SjPHE6IQyEGSKxkDxeO//z59ESCIWWa6f8fmY8j0MRS
xvlvfX/Zfz2nxOUPKVc6I9WDxQ6ZYvZ2LfUiAZZCY7pWnaDpy9zrD7I1te1d/UA0
NB0GhwuaMC9iFusOtPMjE30vL7T1q9HXccGE6b5pGYkqI414uqnn0CrjjOYgN2X+
oQPf8zvRdI5yNmaxcsjASkX2szsjq8e4w0nKeBeFz+n6A+j7APr/s0JR6m+PS+5m
Yamx6EoqRGDDdz6xZtx/hQRdzJVpOkjtaiSE4O+DKvhEhL1hNEEsaQ6z50keKxH/
De7u6NtCCYllmDx8eNsC9HH2/Io4jAf9iLmisGuxXuw6pzte4B7GBOJFQ6hF3/G1
M/lZo3bLjKj3S2kQFiB1mUn4TlcXIdFx+c4Rd+yIxxEABE9raKwEjo1TORXgechG
7ZUWw+mcdjtrlqYEuqJl3/OBE42IFhhl6zQqs+ZU0BztVo4bs1Y2JT5nf8AJG0yw
RmiK8IO70Hs+yTVKT5kiiOIWVwXrj2Ra1JGTbrR0WiOk3XK1EadRFpB8WEZPpjTZ
ZH6+f14K4fgOL+CJ0BmdnXqC9ZJuPyA2iOWhU3DjxqiooY8TAQ+7m7hmLqoTu39P
98BwbPWaoTWKqASDd2KYjMuVhcvNeA1G8GGjC0Xoxrp2WRgW6MngOJfQPB2LvGoA
V7jzCFWJo9+cyv4rQf3q3JvWxwgqa3oS4RFKjUyRygkgQgACB92UnvDUbHRoj2Zb
5EgA4GKdgf+/EA5DV8dbcrFFuN/rooC9WzxRVahxdY/pPpxPnEFX/ZX8irqWpedr
xEMqjc8SVQ9/TfmY9QohtDicoRMl6B2sA/kjB6h6D67kOoHSqHHHZeVE/nryPy2X
c3y4PgB3h+2n8twRlMzmpyrJavXWJd9PFlpOc2rOId5c1NvT6MCIn+NB42LMzONF
BXWIeSOBs6GEvXboDD3BC7lm8MvZhsSbm2p0pbKMRMlBZnx+08Whno6D6bVC0M9c
UGypHGjH8jeDn+oHuARhWDKnr/R2fhhNPgrUkpHYSDb/fHtST/kSM8nt2f8OIyS1
RjHV1y5ERr0gFsM6vZ1wv/TZzmOivYyCFson8sV7nFqqOG2eMgL2lX9k2Nnkadm1
fCCEmMjCMp/Q5JfsA9mZlrbuC5TqvhMexzYpgh1f5T+qUxoOOTlAc2Y0uuo1xxfE
TqPTWul3HLZzKSJcxlKWvFKMuZ5Ygbgtnm5qKiWsb49UGf/8gQuS0cYKtIDEwZLU
0B7HDyBlToLxaMnukLP0+wz8Op8oEI4gQD7ILOtoBmgpXK7U6wtuYFK3RgQ/fV2P
568xKyzeV3AmBbUk2l+Eza5/A6ey+cYi4xQXWolU7mLRjm9SCDfQRLGfzZEIADDS
lpNGAKpZYWieyh+RO0CKXlLATn6QLzMTF/NQz4KCzFia1yreAAmKQAuwUrOx1Hsh
kgbXe5vKBpVo1N05qCCzXRscpQxVlSoqDJDS1Ya3a15/mYTawyoVIvp4se7GynPW
dn9He2zXYrf714vVpO7xGyvEw7InrPPjed7Javs7Vac55VvL2IVJMQ9EPzCzOV6F
1v5Vo0jngvTds/BdKLhmayqWRtX1nz3rv4CWyaQeVgTJ1SoKQECzImMJjRVdRaBV
CqfTOsilQgWUUyp8fN/C6AnbasBJa3L9aLNofNd3t56EOEjcUuPRuXPr8HVrLOys
MoiWnaJHlDDvQj7cFc8sQmNGQQSW7sS3wMKAtU5kWZfWer8WdaKzJK0FlC1i9K5n
fcURYgbJwUdCZoPc5nP4pT/xC9fIZ6D/pBOrb4BUnsW3GtAvoBfXEu/cQH5c/wEN
sGS9A46zAUELZrGLLp49tcUIEIGE99n1NU1eKU5JWyCqC6mAzAwq57T51Uq0HdJv
Lk9hEpsNL19gZqKYlQ2n2gWajMZ0lRUMnHUnXJoCRj8uHEYNqvldC0yi8eVhWSKU
0o/GRSAnloM8TDt1CQELz4ku033h9pjUW1SFAA2ZjV/4MmYHzYsnOaad03rqTreJ
NvYoo4Z39R3GRClAdF1+tjcCeTIAyJlP1qynWwozvhiGR12Lv1B5eHA2BWNFTF7P
8e3l07ddg6LkATi3JCI4AScxn8gVl6yAhyK32/ZUJ+BuXt1A5CmsM48xfc727lOe
Wql3aQduLjiBYcGKqP0cSJcG3++iFyY6Wqm+CrtxhxygYcyKuqMRQEMHd+xJW4Bx
ZK92ileYsPqCsTExU8LkNYvQ/zWWYTKbU6D32AqpChlhZlqgx6dIVOn9Bug5K/C0
WuC6J0P+nXdpj9nCfab2CV5ypNzjg85f7vvqRD1FxJfcs371gkTsfj00far3JLBB
s38pfy4yYDmuoMwCGSRiB8nt4YyGr6ec5FXEPYJ/YkSAMAyVKh91fl9M0kO22j6H
2+uKiWnss3SSNEPZmpQN/u8wLYd7NM5OmGd3lrq9NzOOk106WagR8cn7Y3wLXf7/
1rGPWaDI9d5ukez3pNjYru8XIZQV1dIzxuApHTpGZ+YCMWq3iuM6x6gJS/jhTN9Z
Fh0y4XD+4lRGkzgCVmM9gVcm1Z81qSFANauu+WREr2SThmz8TmZXqO27Gwkah9Y5
2d3be270bNUabPh6Z10CflzP4oS/AMwB3u9zxq+FqG39hXyHvJnLwaEQwHUbrht2
yOWzxlUcV9GEAYDZRRqb4kx4O9b1+1tFsUYc49/V+Fy9Bcan9U/V8l7sqCzSfS1U
N4MrrqCnkjpEQMpo1LLxkBDeNdAyNVgyUZge/VPmzKlbt9APYX0B2FLidS+7+uVZ
GJV3g9HYWwT82fWrDtCnDluGE6EM4hQ63sOa85RDFy+NiTgDdmjhyjsO0BYjNG7o
gBkfUJ8nxk6m2cXaEQEUO+TVGdWIE6NtGOK7VmQs17wcjZcla/MsQiK+diPIBh2Q
nj966VQQqc3ig6orwhRd8nHcPyHdryIoze9ll0DWLuA3XdizpKjrmIQpEABAOZ/J
NeUJaMo9BY7qDdjyDGEir9hle10cEkThC+MWv7fhTAulRrNsrvpMDEuDRYarWQAr
KGVXHSkVKj2zILTeuMoATNr4l1tSW4SnbkbfVTocIWZig4GHW9ZGXOAP72iw5tGn
wPoatmBXSC3BcMDQ6J4PyJ2abOtzCa76hISIsbTEV6eh8Q8JwpgXUR1drUy2hjtl
UCxqsXJ8h0W5kefzMgAiGLduqJNOERHwOM+4XfzzZqUJsZe0f4w4g2F3XiOADPQO
oiM+Wfibor+lvtSxCSzZubj/AwMZn6cWjZhBP1RMmNlN3+Z/1e8Nz8nB7mI7kg6F
fG8HRxQ/l8i1bD6JZ+XXjq1FSX6UHAR8NGD9azmbhezU36a9o3rNN1X1pftb5zRw
UJmfKBi5mwRRBMk2PrmlyttL00KxIqYj89+Z6XR+BcgchPJCWbuQQmyWGVj1t1cB
J8Yf/i+pw62jHY2FQ09O/F81BSVwM8Beed/pNjao49qPTa0qp3QwFUBFMvQMrZeI
lHxU6eztyrhy4SPxC03wqOHIhNEfekMU1l6ksmQWgOJvktpZcnifux/Au7ZJ6EMB
Rb/k6pwuF0IcC3qMHCHfhV+DCnIA/aYLxrNfrJ1pdgJT+nkLSJfsr+Go0oSRR5RK
/5QR/GBNk3aIcaxDD6hdJWj79DOMxCvr9vP02IMqzflcyPBQiik9Q5kQ50gdy9FY
s10RzRu6838iVTOLrLGjopQX6TS1/G41pyFrPgaqGdJjQ/XlKv+TZxZ/3ezLIBtc
594HF4xKgGN3RJLZYPNXCX5R4HoB5PgJFzS/40ptedYb/ICwj7umw7VaW1ZPPH8E
mTAq3IAiHrWhUSnMFVcXUJw99AB8dsrBx8LAm2IggAmM1YEToLaHuQ8X5MF6Fa0I
SapiTU7HIjv2pcvkvvthEnfGzn6PeUnYCbnHpT6vqY4FMzdcrPlyJmDFpNqPEkZD
I00XGuf9M24f+65EipylsZ+1bHZfgh64mW4xhe2iobYkpVvK+7xuFwj6kcfNztrw
NdC5tcUcv6zMleksmq3RTN8xBZ9qUnBY2ZQs7l0xaue3pfyA9/BfnVyHwYjgux8g
eO+1OkgM67PMEyCndwZdDlBYxWKXsHayd3mEOoCpqRQGtNFkcVzUNJ3YWADFXq7G
/ZsG54XaTf8JwNefJAFqpt3VscitK0heAU2mfbNdRaT/STNvB4nETphYzkEsHcT8
PaoJiJ37s4E0Zw0n5oGg2voxWGLVQfN7yROgBwNwK2ZTeHNao6srvVyUhi+9J2F8
gLHGqyARWzh1xC8cYLxpd7mEnsL8IjwX/ajVYaixB+ooWgUJzNiBHEOPoTVzT3mU
Eqpt4ynpilIdwKe3c7dU/Ef343pROL3PKln2fJ1XPQBovp9RBBxzT0ti+cPvXYuU
tyWcbJ2SVwTvpu7n9aJHWijbxuGuJd4ehBNsPBwFLZsUU+r61vm18QAQSzCY2CwI
qNMgdC/ZbWMAeO1on2CwO0ka9IuucprUtkBITibyujQ2fdpbT+BngaKe7fAmH32w
IJ3BE9UYYtGR64JRLTSFoxY+tGwotVqCbswKF6Iw9dl6NhIls8w1nIUA6kRJHk+T
UFheaIfNxDwhbAJFoScxdq68/jAU7TWPh01LqOzNWh5lp5npKpD2DVusEJ+52AhH
IzzfY6/eof6uyepij/cO2e6tVFT2rFsso1eKT21wpJNZn2w+OUIocEmcMYJuO4Fl
vUVvHPefqCFcCF0yu4FUUG5/+ttAV+yNoHBhb8ukYSWZvwxsiL9jMKOHbHjTDovg
mxQCjmTAJFBF0pRpliHYGQuBlZEPElUyjvnM7qJ5dw8gipE1uTk487jGvvSqYJNj
6StvtAwot81wko5LkCMnIp1/OUSHlO6aoduKkDvgNdU2k+TovFHAuzDDZgSi0/m0
uzhrBVcFFwIDPjOxVLGNIuh4c5OmWpfXowcR8hpChbCCQ07cqWkS7iE/4vOSl5Zw
ij+wudxNJuNuqno/fNkc7qFg/v0XeTGmoNH4QeJAf3fcs8dKEG27mriQn24BbrdS
JNssyvdpgsFfltzSPJhqCgmGTiLOkfHehsh22H9EMsA/LpkLqI36zyrQbynpje6U
EwiBRSEXia5uU4BCpwTPjIcVksBSrvP2C7EhvoFf4Yb5ltOWr0WCkBAeDrpVm4a3
p+TgnEn50nJT0W1oMUlQ9v8eeTMQ2TGQiuYEcFL+Oa0cpXtU/4IXT+tTrAI7QkGv
QdCvOSq4EUL54L8yBHd8c/NpYSrna84DhRExxCFOttlZDnI5i9BC/jzzGa4FDdrP
gG+xVAQqG2SyeZ13gSW7BxTTbLxdZ67EE0Q8BdDSdg7gD2H864XmcN4pFA7+33wA
qOmhQvyV95Z5BGrMqSIyz7NAlDxyLYNgfOS9hclpSxDfQTuYrz5lHIDZnSTR0+la
B7mSGuVvXJGJQbN+d0bGayJfe8WUBrHl38rgoPmQJ9+o5dXqXntn6E5d6+fMLM/K
IXzsZ3Ha7Ylm0GgZ8n6eKBA/gdO0wC6r0QyswWjoTxl3i5N/9QfQ6zw043D3Qpm/
TReluuw96huoDuceIyH4qxQ12ivmse1xlr6UCFI7fRj4Ba9BTAg/iQ1suAyEc8jT
yGmzpkgQ4VWIlXZmJ05J99r2Plc9u9359vOcFAAhCyQ1YpQ50Xqhsc6Q0ZEo04vZ
RIowbiC/UAO4bTTIPzSbP2MtgoCXv/MUupS5bBE5gqzPPmByQKcuWwl4HivagwqV
NJ/ZWrgW4CeFfY/5sCoIzptRAFq/sAnu+gYMqUjCxHvz3xMkkANr09MRhuqN8rmo
mMHqB82X9AOmCcQ7qW5YHg76fm8pe+mGwteYlI6SUCeXP2SpEcJuN8zND0b7xuhO
4jNxUbkx/Rxm0/8Rl+WAB9d+onk/75Wx2B7/JYT4bk3kCizBKKclACmc7BtsR9JD
CigLA0KGpJyPve/jgxxKsjKdOKtHRu6nSoPN64RCwIo55yDXGx5TaLdwYuw+gu1J
rW36/NwhXPwbRrilWhV5nSNPOCKiJ+1pZs5qsbZ3qFDSA8Pmwp1MlGon2+NiS0hW
zYJdvWTI7Rd8X+XLPn2nIz/zmGK0nTlMG5ncij/wljbeyHsWFa4xB3Pt6FejZAmY
h+Oae3XQU3zva2wdLx4/S4T7QUH9M3AsCNl9JBN49NbdhlMbiC88m/ToT0hqWnRF
YPqOAprzwIPUo8zoFdyU4bU/euUOxPjOTR3o+845LqRtBH16UhzD9NrSHCM/1DVB
wyksQ4kZ0gOmClMXq3gr+T5WtufhalkxZtV0+8vL3z/MPL/oVJmKJYrlRt0775uW
odXPvC5wiKzDKooGgBpUCEnSFEQDWLLfUgQHU50CXdSsg2OBIxL+XUWmUUw9kmyS
yB6UfwJ3E7OW/tcDw3eC451Er4uhy2V+Vq6RK7Ktjj99Gs8xupqKCZCNVSgHKJki
HX9X9bKkNPDfGZ2sW3btwp4pUE49ZdTdgHmCQnQ1gUY1A4Vj2rZDwD37Vg/7xDP6
Ebiyqi+nVKJ3ahRDO3Nyy1zY8hj3dYh48xOEFFBNCOMWitFR1LtywrfaGiVxvKyX
+a0IqLQ4avP4ojIT9YspMLMLWw4nrPx13hAmcNxhsHDXAYthWNEPiaUir6fwu9qx
HaBglxb7FrW9naWaRLC7F0ZUqD8WfiW78uUWUWldsRxFhQJNMraVCS5iCxE3LZVt
7+L4ozqwYGWWxfHoPzXDeDIVIduONd6XOeT2pCM4X+GRDUmNAf5/OfkPNrl8ls7j
a+bTK2IC+gG/rqM8ElC/gZHd1Q66aUMTOq9KebuWaBkMPo7+udmDGXjHJbsVig8g
X9hOdUHdGrRgeSSTwEgswQNv1OebNKG44qxt1SEVg39gOcqZrgCN1G5PnYqfFKZb
tlZDERsWqzGLyVZ1QWwQ4LIOjaHMNjXMqwktKuggLhApQIajnKLDDvkOpVrg8zF4
puO/A5wsxpULQoGcBIIy4hD5sDujP1Jf9VivsVXI1Af0YcyGbx0S9de5OdzmBlrb
+IeOGaoT9PP8E3Rm01xW1UfoC26P9bpCzWKFpghPgt6PXHrUrvd8QSkud531emFr
v/U1Wsqe3KgCq0MjUv7MfRUs3WGThXN7IX6xKGWOVSvgg8Kk6spAv+6lSiU/FcLm
L30wMMZWbpXGuOVJwAKcNMIM0WZwVhZfK2H0nnNQL9cFzkkW/YY94O7P82YmVcM4
ORM9kEAVj1LT0X7V/IuxTOYIHaI1PaYaQJiv58NEY6vHLq17uD4AWGxxHQmUk4f7
Kda03FZQWDjoWIUWAVvjXb0g4ZoIyi1b0IiTNhqUPGCvmwk8USIJvYHOY4DmTnX6
eUg/wzbtrCClERK3dsc42Tst6kQk+DtvR3CiDGtXsWUd4DtX9nbmsIhz2ISJdE/n
tkTQYGmvYqarJ7wet2ZGolS6cZ0ObSCYo0y6zLY+OqzRgfOK3EcmBGfseeXomIvm
7Klwk9t1JMV38yqUFK0vyLVc1FU8bsRIWqbyr97mPqmTPA9T3ismxD6zMWhmpRiy
jmp+gCkkLOYenEy9jhRRS/plTccAk8BdUj/aIRxuUtxgSlcIt7lLA67zcpJLFLJb
SW8qpHwwiut0zSPBmSM/MXJSGDVQbLBkr2oTcDgvD+2HTK4gYjjg9/jelUfPwlpb
Uhm7LDJ1tls0SF5robVEpCdVrEd+rtdDQu7bEv5Kh84EdVkNFxMMf4nw1jXSiEOU
VvZEYwBcLUrqn1Moq3V6PPlqSx9KNdC1U0ls5yCg2VAE0Ta6+K47quxYf2DMp7uu
zdo+1UxlcxwyRBNgU8i8FGAwHRQl5Gmb2xn79I9bRC01cuER1pXFtMvRx3c8LnNA
JVWCpIlSmGE7L2O1l+18YisSkvTOmvmi+GTcKj0yg9TY+qyAXwQrmnqnWsqmEfWU
pPkNiSiHtzgunnV+csulO+xh3EjkbLluAw/xgm3doERuwAs1AJeGIvGWzQAC8d+K
I8CGAtvGum+RVkzY3QRCiV/YUjkQB0A4lyZlHTUPOr+tf0ifbcB+OZYXspAdBu6d
VHuf26Jl4bPf74hB/ixDCnzPNLUytj6u4PPDkQ8lflHo5m3vzMNJAdu6VwqyuIcU
Cbt2i3tagq4zm0lps3MYdz1YH8MKYIhbVdEa618f+UA2o1wiZxtbP1bTfqZg/X3r
thuvR3d3ZeHanbNXcb/zQ0V1VmKJCSV3PYebI7e/Vf9a3Wa9Xzaog51TitBc0DBG
UsPxhKQxmOBfn70iKu01REmvqghRGvS2kfsHvcGaoqoARJqZ3TPEHx1H1PzVDCjE
cFKHjzVQfI++YChZe+WAGJEFMaxbCzWw90wBmwyztizQmpjucN5RjMcmrI8rXm8V
EQZY6YEp249wPFu546GnC8n9OfNRixc2V87YTbKD9jR2k3MGiyHs9S2qZAuodecN
R8t30dW9B/Rb+sbtfa2UfVCa3EMre0Cia0wFPpOK5axid0ZhIiU8GpOnqD5iIDpo
HeisMWAb8q+LLOY7208zk0CGRZUbt8GiTtCArVETdOl6NAjjHP8Ah/nD2V2uEt4N
sSdxPzxy9vKqyJAbIQ1N2LX6cK3tyvRaue8NvLvQBMv2sN+UeLLU9oH7Fur3JP9g
35T2CJXA6FlDsXnpENCEa5Qy4KdMSixOtzdMJjZEgLHkOXKHzgcwJYEsy5BYYtUc
IjY9lsfrBTaxndTyKsGybtifIWuXEobANBH0JUQrSf94kMIUSriQMMoIkQtYsUsc
by07cu/uWCCME2DfPu4bcy+O1vduDZKPwmfwt0SPb3rmeKMfHWp79vGlkCI40eM7
kI68oc8iClrDtvHwOr1XeeKouWfjHj37k2K5RqDT8fWxDIQxRBJTl7uU8BlTZWlO
yTVTTBLmnDAJq6mmd5Aoc3IL8eHqIYRzNOMrP1wlv2h53HAhJbDamzP6bxlEBAts
NSzaWbdOvGZ6/fpVJMYJ7t3g/veWQhw5PNQ1mTSsA9/52DaVLnnbERRe4VPLkvag
XKEirokHcj+Wgu7/XLQdOFLlqDxsRcl75ZoJa9pqbF4eYlbWFOuQ2Pfn2oKTr6+M
qgyS0mDeXE3l9PZ5r66oJcJo1PitZJj/kgyEFaUUPMGT9kpuqEFKQ8dpQV3grBwt
4oyDhYp38+jM8psl09Jt6mzitJr5znkufokpRZXVxMfwia82UXxtLh8QnYZ9pY6J
xCmVRNcln2Pvmhz6X1pzzEVqZ9zrLdJPS3aLcnyZ4/qcKXnJJ2IgO/gsPfdJPUkD
gY5j5Lfx0rUaHpIv15AH7xaRuN5PocbD3VP0Aifuj/wkF+r86u/+dv27KXCMMDtN
MzsSnvOoTkP7ADfdu7Fk7vCcW+95yzbwDmZ4zHFk3uCMhFPKziqC9dsQrRcfWzYK
Zc2Dy+8Znsn+Wq7IrEja/fwal710eC9derOTdTQwWQZrX4RuwvR66JAWTx5UM0Qu
m3KjEVU5ne8zKQBF9ekNUdRx9BGhXE2qUQFVyWqe4zmUZFN7lko4RNUTzHEp+3S5
sml8YDcQFmabdg+HgbsrPBpJZY3HR0uf5KbUv8qEfrzZ7y75DMy4OhdphL1cThNK
XTGn5+CZAAu1fFgTW4XjRQpS5IqD0iuYeB84BRIbVqddG2B3pTKD+wg3JYz0iehJ
BpLBqGRv0EjhZe1mlPIzFIn8dAD+1jR315etc3vtV7mdkqOm5m4CZG0hg4LfGCzV
oRvAN3xTZoVeQnjgJOpqfioe+uzrl03pRQEVTMEmaxhasJXMbyRQ+kaMqycSpVlA
ngBqgD7xifAVuN1vMft0wACcTNcByy6jl5UFiKD2k4lVuSwXzVIeD5Gy0asaNaJc
HioIQvxNCNxEICcqYIV6RW4IXaMQaenmrflu5jEmaS764du0GVJiqoRWIuuwRW+p
EyXEXWZ63sBBXI8m+3ydVdVdIlNrLtFcsUCosvJWTOGBvy7HxbTTBnVFLVtN1bB0
DSBmVv5r7gsTufiI3O9ovDuotV3YtchkBpwkZZBH5EVzOGe1GxjGccuoCptiDj/A
mCx45K9vqsLeW2eUDcErUxUhvRet3HQqhPhXVgLvE4oBu/0V4cbi0SYaEtWkhDII
krCqLbWCE5QfovwyR69Jh9ProeckFlZ6bxR9yVx4s+q39OwHzAhGa58Qs43EBAuQ
t/nXXp2D+N++J/a25QBIJdMyEYdxVx53BHbEwUg/WiTj1S0pIjO0BEFZCvGEWN6m
La7caDy5eogs5SYo7J78vePDtwms7OeL2XBSy2VDntVY7F+YTensJfgrtmmTytG0
XDoMS84VGX/TJO4ZG3Z+vgAVJcFwZzB/TtxNq5IodLnvrIN7mYA4o2EgGWItInPy
COBf10L/QniNcH/2GuwFDD8b+auLxlJKGlg1YhPYm7t6Chtai2PFlxRG8iGdPHYP
yZHmKwZk8Pw4inkfplKzI5YWL9LtZiw1WHsfrhtOcRuN730AhErz5YZkNL0xx7yO
BNH7viroE8UzorSTUUKQWxOy6bBRDbJ79ETGZc8PcYE6sIWgdMz9CUvHCavT70UA
//1f8bXF7x5q86oCSX3hJ6vYFH85H9HEMDBE8mDgxncNE8dl0ukYEDLoquFB0/1K
tlk6Fps4H2kwhO9DbeeANdK2BhUsK4jrlG2SoCM8vuWmjHchyEVKH6ypc+bAriSv
IVP0ncFkctPyT30ykK9+NF5QiV4hgtPeheTvFczmzRwHZD0doRMS7PYGZUjvMzdI
ZUtnFn7MZPTyAc8oqpxPV1xYoqQPrGBNJQmJl5P605iXKxqeHWBooYPji4dpySnH
4JWR01btYc60JXk/mg0iHzf/VEHlXzDiurTpG9R/CESTxuMuYCFWSEZiabWn9eaX
AvwZOOm+aOyvO3O7pZgxFgcCBYOJo7fQ0uQs38w0l4OgOH9TIB1q7GvYs+KNcs9g
fZ/JmQF372NmnJYWFybOK7YktWItrUOh1pouJMNhfabKOlhucFXKioBT9FGrq9QQ
0BIAKo+HZZiRtDPRLoUfxRtAhzObrHZoYzAUB0JdyxwucB/exHUKq4kMrhCXA5RU
SaRMtwwvEI5+2KfvYLXLq4koyejU/CJY7R/MZY9XZFpQjiu6CE1t5WnyXFbGhiuO
4CCq5OyOgDbm8SgREGOl0c8O7lvzXiv8EPk43+N4c3Hnk9oNUNmOGkihX84v6E4f
vjHMIeMLbVGm2xWsEgtN1NkAI5gr/JyISzOZDSypwJ+y+avstOkP6SeH7lIHYeyb
LsRJTlWortOvAzw5tia0hK5r2gUgOfY367Llqkq+XDBLfkAzz60HxtL3O8WAxlv3
svWXrFEbBXbWvCe4iRzfhBR5tedPHOx1V26TeuTafRi7xgoc/VUOzAsUMVendfsj
xCTXmQPMsG9w3drvHWcH1LQV+en5Zz4+wW3ehTvzY8b+qzTpsqofrDK6/+wMOHch
/BiKnoRmOS6j6UF80z1Fz6vsO6FNHyqJSa7v3hk0yYyVB7figCjAHbYawwm7vlri
C6iPj4fSlXau/H/PQPTVaMgZXNYqKk2j+ZIhwT3r0oZ0+o4WRy46A6bWeMMTXpbA
hDEWFhehxZWnRGAym5j9RUwMonKmV0Dypr/3CiGxc61fkaSOeo3lz9M82HIaHpb+
Ixln5CacJB5Ajzhw1GG8dJ1ZuuhCSK5DitMePDE9dyvE5Q90UbJQhMWe12RmEf6c
S9PwejB5U0m+waOzsBDkn4CZf6DMMyp/E/Rq89khohNjgQ7FuxviZEVU7QAu7fLN
aaKJ1vQ8cb2TyQuErV3/Cyl2+MrOq97eKtsAsxHZuJxiRNqlTDqNbYXnMSAWtGt7
Xz/aG9LIaOV4isp7Sdh0BEyc8o6GCkWNPYzjZAV1aXzjjmXqID5nqek6/XfQ8X3D
NjN6hbiiTqjnzuH7ePeH/y/hjQYquQSMlL5g5xcrp4ST1j2fJGkYJ3sf5ygq7NEp
BSQbf7qRW/k/amBivEdIUjMsYiwoQAGKt2VBdbZxLNBqPDJDbWWcWOx+R9g5ot0Q
5LyeBmYSnKN+5wdcC1qpbUV/05UDyzJyxYLSOEdm+M5mCBq5zhh6xvERxnsZIHE3
/K249hT5neYrMqsNZNRJ3YOkT2RAsGG4BgamwFp6V/JeMuoLMeLRt5SLd5dguqEX
Ov9ObgOkPNw5VKq0Bwi7iphSl6IanHGdESQKpsVBpff9TOCW9KNSZ9yFlMf14MsC
4YJhW7CV+kukLSHET+JfE46b8ASp3TJFNC6vJ4wxb70QTUWCNWeecAqrE4MFHkwC
e4qEj6WInPx5dVCGDITRkfIyzTZbDkEG1dv0FouoTMoviDs4jauL1TMN5iMiWuJi
wSwF75uD+7emLIYe2+g4uCqv6uyY4JdE2+QrzS+yA/jsi1vnLWL0q3i+kmeHrgW5
RvfieP+hFeTth5v9SRmjbCgNdXzXEG7i2gxXTf/iIFPB5OBYioaIVpgS1sx25S4f
cC+asAd5j8PjXHqrLk2XTMOuOYuFbnvS9RxCUGzRTCuCKng+7/FXSjvQyOsM2DyO
QDx9RRkvTrt16sclZUWUrYOvE10YSzo9uPPzemodISbO+CsRaXnCGMoXMRNDlOnz
DGsIX2xveOfhpLxPfJ9ob4Y1kTsjiiD//SUecsdYcBDf7TMEF4SREsUKfyOzH39P
SRzLJOJPqhkOFgt0eEplRg+dEJMSJzVy58vE6jjoQG3OHLy2EOcVViZjEI2Lpbas
K8IT5uVtv9G3C7/Lm65LTMbFo09kJCtetudOLctuMLAt2CZwXXXwjc/pb8s9fYkb
mTJBny95pIs67gMDdJCGQhAxsOYFdqtS5lRGTyR3xR7hr8BngfuoJtAF/DlGg/tS
QRYtAQZbHVh76gZ82vVe5vRNGf7636i4FjMFV1+xKuZJwYYTCpSwsdpzzpmOY34A
rz5Ce2PQukm+M4XQ0Put5Ijm27+O31QpYrJz5iCgSaGnBPvbrbeyaF+HXOyCDYQs
EYwBGKsh2Hq4bvG5xcFKHt84daQvgDDXI8Z0ulRG/uNdiwrDs4Pf5Oh6+/sb15j5
/1e+2OkWTvUe5iBbMqznWT0iBIo3KgeJOakD2e6wICMfAdmqHQ2xnK/N7UKvAx8B
ddLWtX8ZwZx+HKr68vdNpQ5akYZUYGmyYS0ZL6yFvgV0oIw+0vTCsXCebEgIVu08
IfqRWFf9e2tJw1A0FJRonVKrpMmzJVhQeAbDorF1Hzxg/fMlT+dfbgU0vPBtsj/e
S2mH1xe3SVMMYA9MRg6pnIjRtWbyuSnjI93nwTKkrFLXWBDqUC8wjtsnf5vNy5Yy
2Z5+VvO9xO/N1rHUwsCEkmkjo3LM7tXfmDLuLUPB9LzOXyHIUU+l/yEWJ9UkhVHK
4vfcHMHXeF1TmuDSD2aduiMogp2eDzjruqoiB9eLPxfYuH1IzTYhwEXTypA5Jkrl
uHnVTK3nXgciZHs1DvROtgGvDx6J7Puwx+tK3a4D5c1qHFe9l7RbbhWBX8+9oMIF
soOLnhnft+lD2q2bL8pi+EpL76x5+/kTuwIkcQ9tTpKkfuiX+UvDqZBmXhUHttAs
TlRzfGET+wBwq+sdUIle/tyDe2GBd0j9U5YHi0K1+NIYofv0pfR9fYHmvdkLlCs8
NKPlxb1HKTH89FZ5KyODpLO8B53KImJbnajGrO/zj7b+P+gYwSvOT2rjlJakv6Nv
OB4FqJSLoAQCa5xB+6M5/QrPdSOivPkYCdhbEDxy4xfRJHbeL0oyXCeaUR3EuQbh
8+Fbaj2Wd7NlFs1Svy431oybrxfnhpKO+dT7JFNdb2cnQHvbnCkB5EvdGborRTDF
ejRv3RF3ma5MyZGojtri1+rkLIrudbwXZIVQVYOgDG10a8Uo8Q1z1RaI5zRcRkwB
Linuq9v9zchzb+Jqe+N+LimK+EmgyflW3SGHrb83EeHLjsYYidGXN0IxM/lCJjOm
xf2rrV1g0bcEIv+N/6+51BPXbpIe+NrQT33M92beSHyTqQKD9tkBIjHL4d08THnG
VoHi82oJnUo0ZJMixAySWufOG3BHp3R6RlIFOI9Y5jDuxMt3qf28ksonpKZlGWd3
HJ4l0E9t/uflEDYh4jOhJeO7e8D+Ewo0GEhwPczHXOyqjtdVBn4FCFL0o4ZWFjdX
D3axjtYiQEUEUJ1bfKOhoqnRmeVAAQ6ChbbWXOEWmzqvEIe69jBYRh81V1aGDfZF
qdZxU6HqReOg5Lx6YDr1nhCSSA3ln1RcZU3/m3vMuVci89if0Es4ZuZKbPRIPp39
zDB+Cv9VfsS2ewz5SZnIbHRVJkU8YpjMLGyEqUd3X6uDuMzrGun9CLb9q7QuBnMl
2sNZOIbRYvv8Kr4Mm+OOKH8L7l177XpxcupjhvmwOvg1PGvKwFHK99usjnA5WqPy
ivqU9gfRzj0D+KqTSYwuGPYbNF0lAIPIKnVw46msTstv6Ydjthzpr9fDY9p0zpL/
jVvqS4yJDXvGxxGZwJM4cGfXz6yqMAAkF0+g4SXHmadIEsHzhnW59Djw/1ChpzB7
XBcPMspSlTxQm3iKd6xQMJtMl6YYxsWsMNt7MDkGMvD/O2/KdWSQZzSzEa949rBT
DjdOQy8uB1ndUiS7mXXwx38MBIofa4+HVvBmEuxa+oSR0k4sBelEjKLFT+ku9Z+0
doEKHvgEmjrXMC9zOgPDoWt/kvK12eKtXT8rOS6ilTfxldejB7eUUErphkl68A/1
D58yMHVZaS5N8MCSScdTwVgeiG51343uBKnldp43gM79VP/tg9iOH3Ay7b+Ajjm8
`protect END_PROTECTED
