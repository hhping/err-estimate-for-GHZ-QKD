`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7Nxj4aYizDTmLQ7tEqV02i31DEZAKdtzyEtEkf/PvTCoGu6Jpf5Wn4XYvyDDOs3
2GHTyRLoVMyN2ysnrPojL3+I7fk5iqxiGbrtVEUi5istxaHQHmEEgb+DtC6c/W9T
ox4Q2FRTVSL0cAygbNlJoShyL/kpafdiA1MlBnANp2ulTX5Yip1VU4NaJZQYAOr/
Z/5OQkNTDKvdSUGZPf7LCCnGJiq5K11dcJlABK9gmbp1FriNZe9Lbl6MsR42Wof4
lHI6IAk8yf2tO6/3RIhenPFpUA4GQjw5LDoT+5Dhl+uSD+eMa31suwlnyOZWbEHJ
g6042L3m1PyJ2Evxi30EekApXNdaTYc60DfGDHxB5N9fIMiEL9nUCc0JkTHwE0F2
KYSW8XK45aFuHk+H/D/W6dk/smKRknbCu1fBJgEi/oy7LLj9kRW9QdPbu6np7Qgh
mofy/cB0Iak2idelwEHIcF1LaSvyKUSstXCgDRuhmM64cCPpVo6uk5Uqlw/Wbd1z
7McGYHoZQ26Q0/RD4S18ruEFRrp5wrJEyWzQpmWk09MEiJmpc4HtoenAc4ntL3ov
iGo2VxsSIJQqsSJWBAfrlspE6cF1/vX66+5hx3Mky6nrlT/e9Daxc3nf4bUwkfIW
TLAwOzLVpFTncmRZS8ugofNXx77W2jj/FTctIlpLgXrdKOEJE3wBI3uCAf+VG5wz
10cTEUhRU8RmQsHQIZrMPhksfuLcb2kxCqwaPp3yeiQjMm3IeIyMsAPLegIKpsMP
CWjs4QbaG8B3sYrq65NN7vmAwEM2aBqw6tHC2sWkO0SRb09/MhBg+ht7+uFn0MdR
ErPfsA7GYl9l7gI+NKcYvkVexZVl/j4GMAF+CYxsCKPbzAy0WEIKL/uQ2c0QMYwP
ddnk2Yv4rjTzLfcKd68DVPvnJRrP9fKSSe3vxNkYbtW0UWy2rjEUqMDIn7ATIb5e
KszfVXtivs6Zm5QjOQRVT+QjhVIB8knt9ZSH7GLvFrN6klyPOVpvncPHdycSjWRi
5ATyJzDQ0HuXVprB1FoJXmVfKKUShbaTXS5zrn2TlJQ=
`protect END_PROTECTED
