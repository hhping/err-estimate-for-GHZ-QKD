`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gm+GkZ/SctrEOjC9rH8gtFGYo99dAjIKBbDls+rSh4W6W1PaBU/iBUxOS1BpEL6D
qfMAZhVe7UR4Vxkpn3YIZXNQeYcGzNeZEukXKJu40iuTO0Qch4MqNFzR/7rUyFov
B4HKQUdvc4mYO/4O5hxeOmDhL3XReOjkGkp+Oj7USCWQk30e5zw9Jlx37MN/6IQo
k+cyNwtMZEtb3EAaXsvok5y5WvGu/9dHFT84bWFrtfjdqcJZd93iHKMtH+rH19Wy
NaM2s5SRFozI0WNUqSaKOU29NhlnhE9FKGQ2I3Z5EJBZGb/CQMSNgE+TahrBGm7j
6OM64RnMUI2ZyTgm6j0fF9pJF1dhBiwxF8Z4odiPcYxhAQFBn/iSibU4+ZX6u/9K
GMgnE7PbWzA5PeCl+6GEbxgemPAgHGiLZAxK9Me08iIkO+SSUYHupgSuPIqsC6Z3
5QOue93ZV+FFRH1SHXaWGBH4yjDvOT44ZUGbm8tUqH7To0JDWIpNmfLuwAcrC2VQ
8Sa3zh8bApnKzVtTzzuoPUHW5ONmEVUmQZPLQsJ2g6p5W3/usDnLW4Ij13RoYU7i
PtHsfJXX8MZpLR2mYZFYurl1UTx8l3tI70YfAuS3YO6Dz5OE6ePJor47Vm5SYQEs
VctYXuTINftdRCM4Ednme7l9FmecsxSdiFZxu+8GHODgZA/aYXhTfRcYDaAlUMuv
Lvcmpq5cbITOHfIta0kPOp6VGd/y9DNjRvjtynCwyhiTB2q23t+z872Mur+rhoFO
EW3Ye5R3xXu/owJ56NO/4rsxD9N+YSEvzdpE7xqvJMZr31GtnLUfeVN5FGLJawr5
atLJkQuu+K8kz7cWMKYp5GiCngsb/y2BlB7g7EBJUWjzzQ/6xcBsnHZKgSjTkWLV
ISt+XXU0jccLbr3xxp+R0EXqGI2Hy2pLrVFOvsAxgmoY3nQ+EEldNeo8mtcEaZLB
TAvEMkEL169qrMgs55JGU0ORdPqezjbF0dgtVHQYg0QSdhivlCZudXCct5TzQsrl
VbJjesRlY1X3uJe6mWaNeqAi35K+luvxbbUqXpXv7unB9wWE3j8dM3F+ln1BBZfK
4yReA8jdo81xUJ8Wog+Q7TonPtdfdEzmoUacVgrroSLm0VQAPutxDBNS3Ys4s7EJ
qMtuiLVp4Jrgxt19xJfKcHkkmdTE2OyB8QydDawY4N8u5rP45KiCTuuhccfqdwrw
2A8/3FXHx31ckVr/USCiH/XlS2IrGPoJ1hyFSM6O012yicHPInn7GoyjD5ShLdSr
sbnjnM9OSRxtIi4ZhfyPyzWBQjdGi0Cb+JGW4NbxlykHpw1H+8NJ5tgrFiF0/pXl
`protect END_PROTECTED
