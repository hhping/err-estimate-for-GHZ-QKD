`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rrYG2f+X+JbZl79JDbW26iSC2RuOMTKYK6QZAl/F+QlmIjc5tGISKE48/DbwMaYX
aasfLaqH5cUE0fJjTFKv31AVhZxANYB8xxzqcvHVL5mL++GXIgje3CP8oWq2Yu44
hH1A1xS9LksQIbWeaL3y0We08nCHMDLH7MN873aOthoUEnJHqXkBQvwbNOP3JlF8
XsCxnkuAnV+AyaUBpI7ojnQMavLTAqW4Q9vg+RcuS0NvRLcMOo8SOO2dmgRdrGSw
A3yTzIxsetoRSrdh2yLdUumGxOjNqGgrZvdEW0/SRwYTT5OdUnnKOMgDtcEvHV93
fSS/ZAVcl5lwWkFxa06qPf7damok3XPSBkl1t4oFXCH4tauNu2iwlvjRUH/Hja+3
wm1xPs+/OhPrcNCUy+fpgPLb90oXb9rjr4BES/lrU7tVIZQYFRwTbW5fsga2McKm
jiRwORlA0tDf1isklI0iUFUc1e9zv75bmfSBzNB4QOAdDy80KrScPvK7wKTbFKCY
nGWvLE4mrrfC2awnaM1URq9NCtpKDyE34o+2dsYzWGVDnZjtOkcgP0V/Z5whdsG2
FQCZ7GkFSkwOmASoSzlogRsrqy7oRBgP01cRZpt1irVxk3LVrKRu5NIdeqfPjpza
vyyDldezEhIYsqdMcmw8S7J2GCUN5d8m/NBKX+zw2+WTYpeNZM2NYVjzN8fOeU/4
/PUPM4/7btXU0/JblwEHQlL4dIMvJiU70stFW+i2S8x2xEhOiK7fgCAs4jdaD6Th
vI6utr2GBtgVJAFDRNyl3Q8BwHuuieLaGnE5oKX4IfdIIGE2gw3TeV+UlQj5vAOc
LD7nK2/90FbzOaWa5c30UipDLX+pnEykbVWjOeUiXISrCZJMYdWOJO+eX4SGnVs+
eWQld6LHZAvUi3jADJJ37Quu2QkQK0zPzZzm/udd0zWtMOv8Xaxqmal5nNcYCrj3
j967tIKZSb/JEQNd+w+zTdG1EqdUK+fONdL426GCR6l+tyEufoUntLj6uKWcvfZR
TR2v3DgL3FLDkc9YTJHEA7Y+IKYA2dyYKbFBRPGfDfatwrKjfrNwFt1YeNs+7Kc0
T4Jkz8UahiHaCSoHjQ0vAn0cfTtdBGNuxOMGaQmLaN/WgVkDFlVZi/E6X/esEvds
7/uXA2OPVDjdS6x+wmcLUCucUUB6PPN2Jx1f4J06bQrd47MSLL6BF2YA940N5O1H
YLaOV+OtiZ99ObMSep2lhAKzw7KRWSAXxwpxtMOMwi8rspQ8QxFG/KMuE0TQ7TI4
clU0qgS4ORiCdncK2vBzHXGy4F9G/PCj9Oi3rQLJrOGPV5jg0oQzcTrn9DFrwCmY
1Eyyw7HRiJa4YA3U4xiGLuwRFeuTaHmnJDxb/lFlv46bb76zlI7mwKxI1gVyZLoV
HlGcxkXS4MzXgtiR3BMlRRSfu9/oFQ7SvUqTth3R4PE/ufEoVxG7HM4cFz8WSz56
+huIdYj9G1X/UPWpe9cUiX8U7IDfajyQlq80Lj7WYnhqy/QDRrKI6/vNi4ljwixW
cxlP3y67dsVw2tXDUcX4E3fl8gdj0CgdwqkaX55yd/qkTQsOs0kFWoWBHdqIBSWc
fEaYgq3VMpo3kDQonjw0HgHDCnK2MvGFHOpKUFvGPZBm8fjfVQrNQy5jSgMdQgQa
qKnIKBHo96C2LnAXBvASDH54B/34H07hwEAfgg7N/WC7QHwlTkuHnzHYaRT1l5nt
JyoRLNcKQqAkWpNQhNeV/rieU7jF9pHhRlSyS6gQShnXWyUGAdY2Q36otCZdWRls
/MW2kUb0Jhk1WcsYmoM9itEhSD6TS/MC7JprEwUaSSH3VOfpxtm+0rIgQwQ+Y1gS
BJjYChy6xiqx1KCvNsNsztrKBuNbvtL0XwnBja6yTAioZaNXetM6rfJrrhRywDcc
EM6GDxeOhxAP3Pl1rkhZMasYVVxJHlYkVAviByvBCyNCnXIlhveVEJkpPASP/JHw
RyhN6cUaHDTLlSts6BZDVOQZARwgKGDwiPZNysL2OOhVkPh3hXCLCiTS4T+qc20J
R/zdler4XirCGuwZjCNwbHNUlzJrl8cODkrWrX5GfbIVrp31SqOAYuVYJH8/OsoW
ue/tXy3JT0rYucExToOPAn0E7g6olTYfntL04kRlZV80QRrZ4bTyRT9fLibPgc82
eWAp7evsJ9QD/jNBE5ElbDX/pRbpp9l0r6CtUKTIXOcVxqa/wYNM0xgCuQBN0+lY
6vUNzXaJ95TT2q28rzpqBPgqVFk7V9gNZTU3ZORjHN0FDpaDF+3r6k75NQEv8EmL
AqW0djmcsR20aXoRfQY6VYwaA0HT/SGjp+MOJZQ1X59crwP5TsToAIRhGfmuC9BB
xY+UoBcdvfxHHKtq+pEKnd8Swd/8gfLsF7jmS4vjzPUVrLpXZoAeRxwi2TogUyIY
zypkY0eOe7vlF1anioVU1JYdmtklkcPaMnoURZV2/UJRDQHbkmgN/1lmWpj+3qoH
QxeLthgGdq2Wbf4ap4Tl7BF3liB3Fu+OZHrgVSm83kXWHE+RIBiK5rcA1EwBsdh8
aAWpWhiXN11iawQA2kRjnNI1qIDThQX7SBuy8nRBJzzefdlrljl1kO5C4VtgdllH
sDjNFNo3zPbOoGNnszuA86bLwYYYLDI03b6BdmayvHkNMuE0l7n9XGsnf8n8DZKv
r3cg7CHkWX6O8APzCe7pS0VPvDBI+Wkk3ruzwTV2VN/fTHLP/e35odhpB92Iz7Bg
hC6ou5Og+y14EqMGLR0VI7som60dtBTeq//ez6/11wF1VsDNvBbMlhblhVWiMvBH
t82pc2OacHK+IF+ffhBuIFYM1G5vayEmMytK8jEuZfqgwohXz5Zh+OAjXVBcPtUy
OnqTdeyjr31tbcDQEuQTVSvFlmRVtA8ReVA+Q7TufU70fQ6yal8NzWeHSaO8qu0/
tsa7GUD+9obVBFlYtksY4PqjOSfUhIe0Kzr8AX0ys7QODr1eG7FpejW0hOXb7zqn
Ymkg2Zl7zkwyUCn+1JNsTzi42gAma9K3qDWo/AMYC9bBFJgTUeN/u9LAlzqZDOqd
PJH41hcVZAg6kPtAPuc33RYGtqvJvH88hEsdE5RIq9xWYsizqlVCgi7sDiDP2cZ4
FXF4Ht84jrze/i9LxwF8r+3iPDli/Gq+/FKZg8Ta+ux15ip2516mCgtto4Y+RrJg
3pS8KwgwKqhQRxd1daM9x5jqxvPI+FbFQQr7n+pkf7+mshfmf1Dtt+SRgwjIG4Pw
InKdme3fhlC7YL1QY6MxgO4WDoXbRPdr854XE2MEq4RNCEon5k1+LKmnahxxTwzO
zMG7brqmB5galHQQHfNy/dssrdBI7tpejFSBa+pPooq07h+Yb2BHR10LQRYVF7Rk
/IiOcWc3tHl22Iwcxf6r1UO1znpDD0AuUGZJeLZ2uOtOHWGgIAb5TGC7Cp4a+ZoN
ltjODkScTg/n+hYtjuiAOAhNFfTRlyPKwR0Eg9/U1g4KH8De8CrXj+6rUiqv4ryq
oLQUaV7VC+s3LFLYlFQneXCPmJZzAdDQVntvscYpcQ7vo6GzAU06XM2J9Ki01+pw
XO2q5bmaCwGvVGZgpHn4OzOiu5bRw30TftUROMd4Ip2sJzNH9NrGab+5WE2tA4Cm
UWpJDhElgRe08N6B1OaYNMZf12f08UG9qKNZAFIHf8aXRjL03+D45QqJ1nSDxJ/l
qIYX7Pf9wqelKOjOss8xo7u1VxoMsK6qgkSafIeuMb4ZyGojAGYmRa1ek53/AK2V
VspiDKdSZJXh4Od/+QiyPDreLTILrTE+R7bu0K7PngaAXVbjz6pJbyaFBsU8FeG7
iOUtAlfcSkp0oQlqXir/4mXgTfcTnPRH3cAVagVpW/ro01SAT8PMIqzN4JcCqauQ
Cuhp6KFcaxNvXD6BKTugJO+CEWNSOZt3jedGrmq9+YDvIQf4FFrA4isLUwjAlnFY
j/hjmapE6EUvNV7WgIObW/KQcaJrgr2hKhy+Su8nzNuTLS2LH1BePsjyOKwGk7Ws
aXRxofWUOTiI3Z8f80MIRqBJWsi2ElWvVhMGr6ConjyVRrNQ9sNuCNypUhY+/OB5
gaQTlZvHP/zjGn79T+u2hF+xiBYW7UjODkGn/jegIsc+uEINab85Dm7aTjeHYo5q
3c6239Xq9Wyq4lYIWV3CP3W138MIbzX2o41LpCEBqU5SpBKyBf5Z/IaVsnm4BEej
1rXWkeULNkUsfJW7VlvlharKaiPcm49A74UbQ4433AxpaFaHlvzJmfeWj8dqFs3R
GV9rm3HF27LCBVhDHOhatyd2g+AkM9pyZs3YF8QvOsw=
`protect END_PROTECTED
