`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ym4VSmbdcAnuZd6DTxtC4UJw6BcqPCC/wtwR14KWlIgnS/PZ6g34rNtcUTcIqQxQ
zyNl2ZyfRJzJrCbWoMD7FkRU3bB+K7h0lWkasuH0bNaOGflxurpT7d9IbysV6IcG
mxTUDpXWiedY7Wh0A6L82rk9yBSL/catqhbIgb/DEypCSJquJpVIG8B5Ga5oHMVi
S19bRS6TzZnuKyz9U4eL5ASA8hT97qDg1qEBv7bQbq9jLXnkcTmAwAlTA1NF3SiV
FpqxIK5VFcTCIHXHQXmPtAbTzFQ8q3kc3OjcZ+JAUVwTjNDwgMOu5T+eHpcqXAsu
3WE6/VrzoM1y0/rOTUF+Upl7TmqAd0vMtR1yQrPzzf+Loe/NIZfN4xwye1+dH2gC
n+p1avf1qksPFi/ptb9QzvLTYgyJRvpUGsT/1/wzQ1UFM6uvhZ0ARexwNcjXGfc+
v/9EXzc+a2rMNHJP0GRsTNiKa5vaUMElDsuoKGnXh5SDfVbwILbZjnMp/lWGmDCr
BjO2OUvj8ZC8Q4zr89BXKph1cq/xXoPRFQOm7hqJYbtBAFIENWFVcxSqanCxRmWi
K8bvZhFdJeFkD7lPxSy8GvTafeQ9j85q6mRYTl1SzZeUzSTnFKHq59WXjJWaoBKJ
RAiKFPxdUNLREhtApPITdPHcZpEkTfA+K4tnd+Z2dGqE0xLbMleMFX1mIsruqjtf
UlqhdJLekaKs/49LgAZBWzaQcjCyiba+ZXeBZ+g0dgnswG+tF4R/JIRSvSmOspyf
oa8lAChl9IruGQ0BbLptsLaBk/RbbjakHFl+FJNhWL3UiNmQwmd/pnkhzDclEU7M
1ZclNGFY3kMoNdDBz5e9cK/BfqxdI5/fYv3mvmv/qrBOb+zK6Keetw/dOoRyDwis
uLqbVKfI5/QT34Hz3eOvng5UJkxiNMDE0NebDyIjbDEZkelE19V2ecnZDlDy/CfY
JuxoeDF8pegJmNIuIIbrB352VWQ7f+PhZRoHilOnqizQ5iwCDowZap2sh/dRDnqq
DHbvLjQ5BHlMBRfEqh1SQYIdUB5rHkIBwIG3VV8u1Q/+48cQGP4xiHtj7reIz9Gm
GsZcHlozUaz+qVeAcZtG6CluQGQdcLORrmOBdlWPPvGr+vybk643wVyPqYtPppH9
`protect END_PROTECTED
