`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/SFIMAhqCkGAiS3OB4C7fWnCHHsqtIPkLvTndGP8SVIcoxTk7zi5d7NJNGvhUe4r
sGPaprq0D8uuS4u4KtXKTEhdno0l3XJG/ZskSjyFq3X60LIsmuntVMh5zVzkOOgb
tNZ1Y1OkU+WVnvIBbvGQF7fH207QUz2dBbSrUSRryPoFJ2D+Fei7hS1CxtRQSOkG
5q8mSOhOT7WlnigLjod3MnxSG1uml+DSwamC9C65H9OqwW5dJ/ME+4uzFPubfV7F
YAQ3pBpgmKmy2f2NClrDzLcEsZihUazQtM/9mKyNK4JyPck8Ky/nFiF/FJ1jMMsS
+wmlDnpmtITVmJZRf4B1iU+8Z+rzjJjZty5o1jdeNv4A0yjSH/exq72LM/D4Ro/Q
gKIFO3m76BwuIpnCqMvcX3/ikVVJ1eshWzgCAlo048AkYcMe2CIfzwebaSJdMWbQ
OwGxKGZdtQYp91foBQ5eQjwij6O0mmNxR28INWuLixb2lvCGnCTZ7/vmIDaWQckh
Dh5mAtmssztcyidrJ7iD8z774eZd8La8eZP59T091Wp1YLTi8m/H9iqGunf286mW
/BNKhzz0ceVXzhZpZADtWyke6ezo3UAgmKOZzdzyP6ta9Omb9U+0eBmO0Y66uJ3Z
vwfg1MvSJxAs17a1u2ipXZdCBsZkgUldXzB+1YXRepbTiOW7GG14glC0I2Whke9c
gr5s83qhPrgLO4avLUXtT92/W9gteV4Sps4VubEdZdEt/DUiTFXsF0cWtYRLIOJ4
faKJNn1yCRSkteiSN3a+68WBqELo82JXfuxb0wjj3Uk8kOrywrsyOA0OrXes6STF
hr1ZcFOvYsgyPrG7KOIObML8+S5Z9F1yIKW0Q/bVsatfGpQi4dAt6JkXkJ93X8Uv
QIT1KLRmvFaU1klucbFstcPOEXUdkS12hLeY5d9ofeX+JmXwNW+XjsjOqMpPGyDt
VNKwxq+wsDMFnAUPhbVObKNREvisy+KW3a7JOMTfIQLUFWIHAR15ua7xJs6fQl1P
7t4l0uwflHhbL/0rJdw/x6X97IFzZ+G+jSh0uRySDwAfrXf/hyjftgOWdUi8vLow
BCnjHzVYA76Bq+AR4Fs15iYjnrFG7SobIWgzav3c63FVLZcGhPZ8fkkRhLPF5PqC
Y4kkHAlTpm8QLaD0ieI/gpJ/o0XTY0SqqdFrW4Zi44WAjAnpekaXbcXwh7vpgis3
jAG9lF5vE28Kule1y6aPaQ==
`protect END_PROTECTED
