`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AaFlv1jox9I7ptHrgLDgnU2qI22RgvaafviVRD1dZy+gVFy7AdPSSmOI+J/z85R8
NPiV1xeqk4E4A7/yYqSWcobq43iMtZtMd4NtS4l3yaQdSKMffrJzu1KdR5nXI9GU
8LbiAh0N3/LpLIFVy5sTcSZzl0GT19MScyZeeEuRVlyhLI4GgRGdF7X34+vk2Iev
asfH7G07dAKWEfrQ1O0kYaCrdyv9EoLKPx2HYJ34Z8KzNZBQ66KXv0qhdrkOJJBz
95EKoQf+X0q0jRNugXnwSVdFaZaQunFlgzDr1kJj2ExbWpC8qirrgvklP6umgPNC
L8yxwhMYpxgFgsKJVEwJ1m840DiVY8k/cqiQ38dCP5+ZD6o+F/xpLNP/4hOkpgA5
tu69kTYXOH74BCdOtj/ay8kEAfOQVS11ZVeLXn7pK+Biug5nSck5pfKsYuDV0gIj
EsXRCN1BJ/3fnkkRZy9CWAHvkIFvsQUgdUTU+4kSnJmKkPd8G9zLZqwvuLGFVvfc
Wq5kco6zFi/Q6cIX2gpb6rilJs3apgGQVNSdL4yyqovVnjT1xQTusQ7IewAbMtDS
4Imw8tRvGcsbpbb/ugOrawlgPIKW0vB59NMSoKhWFOHHFQFeTt0tBU+dyk2OWaXw
z1+pc5/hEOZLL+19uc8cctLWcHlAJIupoTQTQV4LRnEVAvcI2PQeGsXuLNuSSoAC
EPTv1PSQ2fXhMxonqDIagfWj7tYQ+n9/aTDcg4k73oZOd2A54cgsUkMiLQ38fRd/
rhsoy4AQm9UKy8hrs44I14mFLOWshrjBpKM0H09+oeH4i5+F0hivC38wN0CKvXMM
O2+fM/BGvyu9J23g7lnI/iwTCGB7shKuVOUHla4dSZl22SU+tpkFJTC33gyvVzfP
Afg3gugu3lqd8QiewOd4fFjYHrYG3p5Ow68JIvgwCoA9EctOp2uXW1aCAJGzdneH
osgGiyCDwHnL82SDPPmdCpsoPG0hsH2vXG7mQEv3dOGTNKJ+RELW3SX/geWZJTYj
axoa1wrmmbPiUMaArLNAOGXbKwUoTzBshnbZTKvlqLqyWn0qzKoKUtwKv6vq3iOG
3Uys6wPdFCyPP/DENtrdbMWPWWvIzf85OVdy5HUKt9SwMuWY2r1uoIHBeMszwTli
xxWYhxkCVOZIhItIuN3Mp06H7Jfev99PTv9wTlJI6GVBM21bLG3Wx12wGish3jLZ
I5Uqxpkayz9DTbgZzj2TCRDtjYU7IyRCmMxqv/kBiZCXmjfjJK/dlIqkcr+VhHvL
5HyWzA601aDZ6io4yWXCCb9dl+g5oc6gYkVz498zXQFNKNR4uGJXSGfRZU81CD8A
z+SRiR9L8qLFyo2tQNnDy97CUUCbkBMhBLdbPVuncrppox1s/aIUwv1ZH+lqAAmO
hseAWBw+3AZPid+QQKWkq1rTAackQ5oiTbq+/fkANcHJLev+oaNsuECtmbiXur6p
eDCCR4+x28KQmnp0RJey9OJjXOcgFYGiyxG3dB92KwFrVSE0rfOXnfdh1rSHOsXa
ZW7uch9suyqCOZPmqYcfYLxGXbU4KSM8EgpblkRlDtDVFW408ZgF74JovdPjh7mX
PN8UG6bcEk/BVaOxSsG/vcyr8Vxldsp+AcmQaXq8KpPB7OnI9raOVcDPhHqB9vf3
Wum4kImcVRkaxilvJelhScZv537cqmVNrbsn+aTrjqdHEldf0nDu2WMET4c0qpqH
w5v3OE/Wc6YCYg4srIel3dzCvXIn+L8TXl91ggEQnEsLcuBzjUV7cCPqbVQYB9jr
SRX/HRSJ2u/o37Q4eMY3HqYxyPSP4gjeQ+W4bi5BkATiHxzUbk2A4dAtHcR065O2
lCAx3yfWivJkWkDY2zkOHnLgTVb1H4KP1GuNsoAvS/rW0IsLl42wQO4JVpZzsBBy
BlBLxqb0XW/7Eoz/hfWXy03iXFGj4xBF6gMk4zUl7vg8HSVsZ5ZJL9R1DCSVyEwD
e2W/idInhI61UgO9+meKTzaPkk+yPGmhYPst91j63Zrmkx24nLANETPBsA0/OOf/
GnnJKMmigm/fbm9ISlaUMor1LKyvNl8MY4vzkjah4om0YqUq6KvYgdrr7G6a3C/k
Ir67/5vOdNYC6lP+FGhT+W7Hg4+EF8eVa5wkz1FgIZCTykL5FUlHiFxuApLVZaEY
zETGF8bmvNhYB86xpgBRtdpsvZdTRZvI+7Pqmi96lep05UQx/ZVw1GddasxXPlzf
x9M4wGgB/nC/88TnTNU9eDB3m3dCfrlMWXh4VTpGf0zAJHUzhVoBeWxF3V9k4s3n
Z+3CLPKDJquW27z4I6DfsQnc11PbLXyWpKEkVbKi37VUW3kMiQ1sScM1cZBHtUbU
f9wzZ/22JogVz4PRIaTSNZ7TLRt9TKNmBg6vSCcAmzmLGLCDvrMi806fj1YV+wUr
0Gb5X4sWfkXjmGl/OCtMPd96gdkp9Pb6rlAbp3EH0JxDZaItZYX6IlTaKM2c0Gbx
GoTVCk8vgHYSeENIVZx86w7YnQ48TetYhQhxX/Rzem32S7FmcD/ZBZvxeq9tTOk8
Vj/wEhWsXTa5P8LZq3/3d0nz7seQJG7O7cVkI4H+H2Bpza5XOjVfyLMdgrUjE6B1
cdE90FV9QnzBUfcbMllqhZxhz6wb4puKJejQcyyrziTeJmdMJrDM01piA6QEHUjO
FvxFjkxqeLINTV3v02jlU85ODV/bVkeE7yIiTK2ITECBAyIJdgkx6Jc2XliWDDLm
nTnduTweiBYGCH1nnkdMYDLLf8IrrLGQw1LnJHOHY0QKDt9X8+RtiG/ta53VCfix
4hzk5FPX3/7bVvXMmpziPbrIuwqoVg12TC45PZDcRai/mnjk3W2fqaZyKLdAjaJf
Hmk0tgcR/neAU1KHwZHFMkwyEwDGMwA+WrEpDAv7L+I9e1331Mc8Eo4/gTeC4WSO
P46Vnp1cNJ3Y8CiRSJJdJ4fDtVG/Wq2Uhk9NDYrX89w5JUsZnQTfExN/Jv7LLTZs
vhF5TStVMkr42tqoHsRmdvFCmaicSkFvXFI+TWv7yYW5NgsvU3Mgxmx544XCAUjl
sDTCOFB7JFGIfX7sGT1WZd9uBdirX5nGYqrmdfD8BOeyD+rGgYWmEUG685rlgMzW
38q7uQzfcKP2Q6FFY52ekG55J5tpCJRfcf01vPwN9+kXgHxQGfNOGQmoe51MaTU4
p4UXt+F9yrKIrNd9+Q6HO3/IXRak4TuBTBEiLNRuh09B1PpobKoMZfPlSO9X8oNH
PYTxj8y8SGC6G1US1qhu7+qbHbYJzHoZVD2mmOjjS2EAM2R1iffO4h1mK9MnJBlz
kuJ6lAHVvZSUW2m9CoLtjcJF2ASdE9NlKFThFtyfsSfJGR8YR/NENkMbBifhUMwg
3tZLGJB5w7vET8tjCXTJHUO80XiNdD0Tcj8do43dSfAOnpfWfQBZPCM/X/nr5URp
7F2W5lS1zPWOMlLVSaSduFP9z+7E1vhEXM6Cm/VMqjtO1j7PkzEawHUfUcYjex3v
09w3eAKrbouVUeo4YoE/Begps3PQhu3a5ucNMFZ6A35DuJ7H1il3afz59EdE97HQ
MyqLs8oZ2UqrhwHPAx6F/CDNF//KuqcIoH2GR7w2HG/cJX/VPbY9ybxi2NS9jgKl
DCXBSINbMjNTIvHuZj8lhkeHOczCIJDsXh5VDOAXV7LhDpHQMZ3oCFx08YgCdk0o
DhhzIdRiSm+yZucxcT/iCi6c9gQ6n+u7iuC81zBusvJg6qr3hUkjfWfHwSJMJt8m
99NiNPzyTso/I+Rou21orjUI4ZtHPoR7U3ss84P6a2wpPzsc5L9s9UegF1zxYnyn
TR3hEdONcvtOi3b+k3/TGk2iKGDvuOmrCuDCHlh988qfpjZP52LG769KSouV9Ue6
YotR5WONKU043auikpkA3ECeda0ZxO7sxSyF4Qbar3/J6PJ0hjMND9SV+0NHzQTb
RhOEJ0O/LHjimbavDMmC5D9efMzDTd9kP0op21FUYCWdr71cFXPV57iTnYmBxknC
LDmVOJajJ8onSCZRtnzDXv/Jyf4TKEPZFJOiX5CITDuyhsE7VvfRkjYNIJ4StDGR
asp9vUZUANbWmBGTQ1lskWWLElsg7rVMyUXbEM9Qo/OoSzMw0bQSeEJBybCZlpic
lU82hTH/I7DKmzEF1CzrZrEu3zN7q6aYJyDRTSlR9XH0x25KkrwdrDmIdtRdFZfm
uKGtXXWzFBfakUIP3JpjZpwOGYM1Rel0/DnXcakm8jBAYfx9l9crA5oW3Qy/xYyD
TdVkMgmkiG4fbOG/td9cMweKfMK5RoEKorjrHdMMtlnrE+HpjSmhVGbmWQelbUx+
URAMMQdrjhvXYmvhWmubI4box1OtI+OwF5lVO0pPupcZ8qAOYeZLTSG0MX1oGDFI
tZoh0+jpFVoQr27zsHBphgbiTtRcE0q8DC4YWAqpiIJA0os1k1LlzWDEidhMTrjK
gbmJxXzzD0Ru7W4mkL5NpiCwg+9o0gBLKJmLMKZ+J3cpBCoJSaDrg3hKPpSrOgHi
nwNwosKZgtXQOXwsZziDykgD6aHNXZmha1WycFXrvaMRlx2m1hhgcjRyFoQf3KGt
JmIn3b8o54s+erDV8s8TL2n9TDuY9Rg1XK6FjTLeHhe6TSSIoo2OuCWuknn0RsDc
vFE19nErlIQ21DuSRUgrmAemCl9epJisl87/2DiVU7if79kYG9OBJboaXrM6F2lE
BHJGSYmj+XVx/gqkRswWDgbNlnvP/KO1K66n2Ij2Z3LQiDfQOJ0lj7wKDLdb4Z2v
gXotMc1LpTSc+pakKZkeYch388UMebYyPI1ZVvZmiCvZ1fwxAzM/T0MtBuoqte5j
UwfxhoOIFyeB4GhQcTCXTmUgvTYf6jFJr1DTWpRIE2Xpbo9bzx3vCq9Fj8pXLzf1
DBRUgBNMd9hiPGhDRYBMXKY7iOoYux8Cnr+FrLn+VkUV+U759t62di3B2hnCgdgJ
izrpLotscvesBGU6pu5QLB50dB+xVrNFVoXW6NeIHZ3bcIgcEUn6U8Uh3yq0Shto
FYltBtt4u1wcDc/T8retIghqKOljEdOf01oGZxSp0Xf7LO6xGSfXEfb6xKFncOys
VQQ5z6/I4X3qXZSnpHWOqxxs5eZaFx/+x+oF23qUkRxk1VZWsLamEfg5lCntUQu8
5/z/WH46xefhGJz9qFSZcELz3s8xcO64TWE498SLY9tgQKJEL3llJimFXNaLjIo4
fke5te8/44paOWiu6oRHcuBjDI4uGqLVGmx4glKvkoZz5Sb2EW6ZdigUf/2BHpzz
UNFYOqmCeKIy85fXg696QxqZKA1ZPtHyG0QGpNtKh0snnW+eisdni1o89osKTySN
csR7PQyodbIX+d8lHRMd/Q8xHlI+lIpkvKO18/CQ/ESriNHsrELD/PlbS8ePW+Ao
dgAoe2RtKxqw8t+oL4QUIet19rGRH+kSniXoYahs1/2fQCjAqkABFJbBP2RaL2Oj
Im+1N5zoUgYe9ckxwQpWYFt9AKeuyzGXf23TQiyzOddgQIwR/WBWwLtN/xGKnzr3
2dfn7hnuW0X+sSx1WL+gpctlCznWAWe/SHLncM9l4NsCaKwyj/dQw3OD8EhQhL/9
a5A0Y/YoWmhZf4G4I6ct0nOqzPWpUlmkjg/ody3lfafAE9iyglopUo/PWjNJ463N
bTlrBTtSMeyazpFywHonpmsBIVTCEcHCtv0R67KXVqjqkxslDO1KW11u/1no3SSd
roMrsWKoWYp5j1UveUIBDqoraTOrpPnxf+HzEi2bc0YyvfbH+mkHM9AQdvrJu0id
V2LO+tv3bhw/hHD/2VuaK2SgKkjPY1wmPpnWBleSGw0T4Xb6kVvy3Zo5bGd+BvXA
2RRZDI9ZODPDU/GRhsaswF+64p+vHFFUYu3y8N+WTKE1HCcaTW2jJNOjBR0DhQmf
TUdlPozu40xUUYDjKBlzQwKsZA5i8feC1kCKpuiFvp90XWQH1Rg5hVLT0F0WHPfw
IgZqVrhOxX8iOtGdDYhIeHR+7LpoVBQ9ySg1oB753d9IFBiQ5nvBLuiiyVBqFoQx
`protect END_PROTECTED
