`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LhTj0HIxqjJYeZTth9rhJ8IRWbmbhqeoPeR1AG8xhRFMCMLaVkvxMExABDYj+x8R
IjA+JjIeywkBv66vs94tmRrP8IzBqZPf4K5yeDwx/8IrwPZdiMCrldodES7H82TM
aXiOxAww06TfxznQ3pBNp+yYyuMV98tjPGMeyjjSZ54FYfWr27TGTSsmldtM7G9b
AL2axaic7/2NYhsgorsWYlz2wfN4DGWJm6C8QgmC6F9XhzOSFr2bzneW7OXOthfD
lyo1PDoTFMa1YrYQk2aV1cxOlHzH2OHjeDqE3XfwXfYlBsNxn1+Wm/oHp/1Ai6VI
1VnU5m8ptjZb46AKFQcno7QgK8LXMbZsyrAm0EgW3WFF1aYtJcgNQI2Kq6MMXXaX
t+4iOex2xWlKaw+2jvl8Y+ZOudmD1pREmzp0ybFt/9xAigRgfJI5g9FhCzT+3por
2f+xuWax6oGPwFK2xjMnq22WgyzYy+vbfr5fm550tl/KVbT+vY7V0WOMrOP5rv5g
SQDNGuLvdA6qRNjJKx/7wP9hVWOOQuaZD0o4pYqs8pG5rTuQzOKItHLnpvM7yTsA
rWzgskyPADoV7Fy/OckCXatZJaKJJyR4CVhe2IXbEEHLcOd/AjB/1ZFBC3ugutLB
tYTMH2YWFfsdUymI7nhmrWqKqLGPuuIDk/AkjMrLBP/H0tYdpk2H5zxTOBvfgbrm
sVxwwt5MFIKHASe421b+L33JarPGg9ogJBnUBk4KEdfHHmgUiXQGt/LA25mWJgFi
Z+6ZTz0nWAO65C2ddgSzAhktI/ujIHr+tvGaP3PmrQsI7W7xAZA2vZZEfeo+Oubb
tauY0kr7kdbVwEBWOzKZW9YP40jCAJNUjMjJpMWYo6UKIpkd/MR4WjJOHGJfTzKw
4po//gG9KQDsfyBj9RJPgwQxolySZK5UTNoeINKjwXALv+s6TLm7b5BQPLVjCxRT
f9In9hEChSJfVlunQlrqTcxI2m8JojkPAEYA1lkVeCagyyq0RyJ7Wnv2cFCqMOjg
J0ODbkpDOT/q6pfR51l6t1j2y87hs1IrtQ4ce9mEXonk2hYw1f2ZWK06mWi4t60V
80zxQ6zzDcirNKRa1FRsWlPAm5yoqQ1EWV/QlLCZrGH2MD6AyyRyYSaMdF9pNHQj
EDYKyRQ3D1lCWD3nhA+VgUzWdmDVmOPTV3AIBKCyYi9ZfYOEv6aAhQqcsEqu4ccf
Xo+/WTPDS0Hxm0Q7DBznFOuryUYrWr4pkwuGFUb8O63kNW8Dlz8rR/O8n3Dbz7ql
PErS6CTYCQMq9ctbW8n6420JLU3l/9cQLKxql4jCIKBzKMMaLo+KRi7jRhdubIKe
nj284lt1e4ok2eXWg9mnqFm+PKaRaGN1pA8HcAKXl4ygP6l9MKrGTFrDqL1cSALv
htm07WZKWKO8A1cuQ3rweMhedZi0eG32a2vOGyYnHWPvszxaG3Gum4z8iejSf34b
oVtsoLZ7HcDghmgfk9FxvXkWHOh5quV4nJIKdbtL9uQMuAJ1kMV0oJiSGnC4cbov
7peZ4SfJ3XjHy5mRAJm3if8ohSxmt80XM43Of+1p7Cg8rbLRogybGJszpX3LHcv0
F2SeXLN1Q9XMq88+HRmos6m3VVqdZkuoCcAH/ajbPr086s3WtLwuvg8na+a2PNLw
NOv5IrqarUjBgb2cx6N72tDpvM1FLWm3qrKEDEMlrzGH3RMdlVEdoPloTEUSOrhh
8qnf+sY8tfqq5STR7JxqXPiKKHzOKIoCH7PiMROXRrg2SGbMsn0zGz7w+4Lnsbn9
OShDP/Xfxwhs9KM5QZ09YHShPPCeiEdW4qkZMG/LGGwX6ReRrOw/nrvjN0dyuKuh
n/V3B/oMkYZj2PW92xV9deKZ107TOJ7WN9jwI8RG4oVVrw5rXgl8KL32rxpMC3At
MEZXHKMPplVR3Uz39Fr7sx6tNR9kmNdqqKarqO2dSl12ANUuOFb3zk0dyJ8d6GVX
zlIGvDcsBSjOTjVfL5QswCzG2PD3C6kCs2cXXzPa/yfBEGkUR/WtkIZjhm24ndTV
r1lVFpWXzcoeN+cMCOmseyRBvAbsy/17ROUVKcu5v548R1G0T9dcWBtuFUJ6OSPJ
e4nVMyC81k9km0TxYGOqXtsZWpnhEMGvA5hMnbn/6ZEUbgNpVtnZVzw8ELDai9vh
KLjJpWJgdikdsb/wy6gUp2n3gTl8popxDrVrLzgtMq7jt1b1O5eNjV1iFPdfQTRC
iQTQHNMeRdETenyw7153K8WtnoN7pfqhL02LdU2SVziiJL+PwzQGGj1qoTwLOAof
686Ekg6ZXhTWc43wS3E+8pqA1pWPm+e/aXjd/DF+gu4egbBp+aeBA7FPIEDA10ct
ofVjSwj0tUIBEjY7hkpd0MLK+WG6zIm0OUG5/M/Zdf+sm6ToxlOyGneYC4+gKOml
TFHMvNL4H6aVdtnxHbH9HtHTfKrftk2Sy1LsG/nVxArRW/Sr/BqmNtGc893UKvDI
VPT5gVS/T6K39/R4etXbeaHg4O7/wm4nLHhhrbxBNTWAcE6VEc2OzhLZXOve+5MC
yCIC8YtNPCf0IFPGstiUIGlt0qrYWQJGQRtwRlcqHjFBaNUCNFvc0yjUfposnqTn
FJFZj2nfKoVkL2UgTvB0hjXz+gZW4wGZAw9GHOU75SkkQvVVpIZnUKta1KssK7mv
dU5rs265/l7GrmeujGX4dTnvcmiGMui7nJMtSxL+dMQnUfJ29oFHqmoj69cJvFfd
F/S5ujySarLBHbbyBHyuwnz6dy8x5Sd7zLQx7n1UT+i2IHtNcDwORV3aQ1kCvMSI
BdUeBQXMMlLs4XOGBkD3GLDlkdZMgUjtVXibKgqwpFy3VVgXJXubgKBbbfbxwzOx
Ui+mEwJYJvtOPXBy5M0S+zOVkAwNb3/Ww62/ZBwo9CWh+SehWTwWzvCvs18KcJZZ
`protect END_PROTECTED
