`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdwlZd8zUQoc35iMRzrRKo4yNJwYarxFzrTNJatcFFJFj+a+KfDe8RVyWuMFFHhq
/Z+QTEoDtRalDsROg3t6dmEhx/dV4UZ9KJ3McXNHk8wzfK7sIOyq8H1BspdYhzNm
lFXqT5WUmKL1FVmI8xlOkBy8i/zM2npwpiCFwmYzQPjYkXKm0Vyaui3GSGRuHu7F
oZmcO1qn0MduBJ0bMjl4T046qfltSOqxbJJGfSymvnSbDBz0mCd/xKv2ZZ9aLwof
SnL4hnjYkduh8jmllJOdEaDlPo8Cr+X4GpfgGJOgTr4Qh2bLY6H+3Vp4W28XqO8Q
82tVDN6ei8jSSGrazmc39HWGIVBuUKZbAsG3YsIF5IjqW4q7SQFvEPkuPnShmsCY
Q99Cej4/MlABY07yEmC8ukizfp4ha566LYpagzmVR7YR6RSF1PHvGruNsK4cltSb
3K45ppTeHzJY5MUiBKPR+Mhhrwj39rq/9XYWfw7CyzrbEd7KjUyJxFN1qYh4trTb
e7Mwndpke88wlb7hT9Xg72bLKJWae4uB4Rk45vQqz5xsieXcssQa+iL4RzYrC6AO
K4Xvv0x6ijcnKMoZEJJ1wSYutjsSnZaUvY/TfBpHZZVgFjnotM+qpA1zO/shGnyB
t0YNvYRFrQLoxjOjGY8ay0BLu6jvsVPBE5iUf7hJIMkmeiSNvZ24YMndv+1wIgVr
ByVqPIHuUOSN9ZbmUTyLokgrtxwPzCInWqgIcjmAmrIYDG18+zqE0YvoEGwkpacS
vOJbX0mvESxGpQauY1wSow==
`protect END_PROTECTED
