`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tjn27WhzHSLzMC1WXimuZKoITSsm8lwnmEEJVbUVxjkg20Eatjs4lL/brr5NqBpl
pYQECcGUfS/wDyu0fYMS6VllKrX0Aax788o9MOqlorC386CqoOb63KLLYW6OYce2
j76O6BXIDUDNjKyIAV6/xVLq8ZvoBad09hwYhtBa1Q7TNu0Uwi21d+aF+nu734V3
F4oBiRP0qPDuD6nJnVdfZ5YL5ppNbu2Y6082mtydTGkOfv2lsMjPmmnszH58sofd
ehTEIlGICtN2Ink3IhaPtJD3/a4S8yyw0J1I7YcjDzG8iIes5PwisKR8gIlYHNC3
6mCrLf+r27mLDPdrYmxqKwYfi7r74iRe4hcikXsC2y36pDCXVIYuJbp290IOWxkN
GayuewTu1AvOC7JY3JAkCveHV1mRMfN1KyI9bK1g6DeK45G4u5MJoS/jJTAdNGdc
K4STTnIV1Xa8B9yeqCbWbicL347RxO7ekgQFK4OQ2JGIzyQiDm4VVhO/vH0afo5d
ETyIm+u2priEGwZGupkGOOm38cf4pFoktH76RT3khVV438PFB+8a758sj+rHyEmm
I4sG8Wv4cQlcUljYw/4CTp5xSLYzbBlz34sxKEk6HGONIYVyX9Mh43efX6dKaW4J
bj0zUj8gIFRtlCz4wWt1hkWQE1GJNdoRaM+hJctfRUM3L0ohuZme9VRq7UVesHb4
UX3xBcqMBIFHGFGOo3CKoX6jEkM7MRIsCha8tPSPUUuxPa2GIwIyk6L/4EuMpFJQ
R+1gy5UYoeZK2uB6efpd7wfgE9n+FrMrFm3AqBI9+TXfF8SZBbMSGtsU2ll0OMH0
uiPF//Xib4ykUZ0SSYzz/yiHxFjFIMfgbP57MlVtdWcJ0Ewm3z3QhrFlXv5rKqb0
84aRpaFUMzLJDUejApnqrft2mmgttUwky6zMc76AMPgaDzaCY31PQ4iNx5OJ3OtR
xDEKGexxi/ejzF6000kfb0R3TdJz21A5hfvgXlEEXNbdpzJHJOcpTEi5XtMycME6
yzZpvCFaH6dMAqpwe121Vg8Wm1hZB+Ab5zUNMzRJFOB9gm+4HXaS0LR7CTw/pguD
HNoAroO0Lhh81j6iUMOlcvvZntktuv1x50ER4CEtGfibgM4ZCWz8UStUpu64Httk
XZjnz07mkKuZYAyoloCWVPD9JuCu7NqXY+LbVvhF/z3pcmD/JBgXuPdnNgDKk6Py
knC3VZSZebLPi9nAjrVXJPO1kCnLUp4dC0jKwdJwvhJEVxLNwHJLk8sJ0MB27Ddm
w/Wfh5gUWJ3d0GEo7Zemqn5Tth6b9gWvOqHsOiycrobY+BMdpMnP8X7sonhsk/m7
U2dJhdNIFDzviGe9c7NhWHuNoSut6zMUzssn1EaB2e6LTxu50iYQByXtv82KJ3fc
xSzDoiDfdXIb8DmuhHU6MNQcb+t2gtPVtyMjDu09EK6vhtXd7vCgaeHg0NYh/1us
DtTcry3qpDJfiVDnmyfqrOPNgA3k38VksGw5mXd4X7MzRHrBsu7Pc+I8lUtMUS9o
Qb9NJt1qrfTOsAZOJK8uA8yrjIt4EOv2pfuQ3qtayXOJr1QxWLBP4/mH7GrTMk2W
ieZ2fJc1h9dHwJ3pgwqKsY1706Zg02imCUvgX2JpVB/aMgEOiI20rFy9AtR8/WXF
3HkPa8u2l5+6B/HC7AnC/6ftIf1Tb2wBjaRuA8rx+ShtCPbAWkaCAywtXIn7NtvD
rsXBL8ZEEGd0WJYNQ9/CVglBk+Uu8dl/scKL33vjx2BvRFldLMbvBv4pPOJY0OmU
/ybJCKBH70l2viDmQc6x4o5KBtrfqce3nBDDRLCj2xCumntIEN9C5y155UDgeCqd
UDGTaEGYY2HhIlg+ONUhwH+ERQY4aKujB+eYCBMyRo8oQYkAWntTgCjH69/Y/C7P
irsFEOPURKbK93BN2cf3vPj6VBMJ7m2XeQolFi993yvhkhZi8QF3TyxhII2rZ2Lt
s9KegpjzKq0xW5foAlAgJBpOaOSmEm8fBM77eM0NYUofW4IPdFF93aeHAXDKepZe
xTqpmlwq2QYIez45M2vyxLtzHh4gLsPdTZ/av+AyfggpxVEE8pdS/sf6IF/MWY4L
V+toV8Ozm7kv9cE4NmcdJzbRo4KbdM8ANkxrRSGxBnf3Pjp+49I3qEtgv9nw0ZUx
URSAmpBKt60+v9WtrUDlPMluvcQSBh3dEQNI4U/9IejqAJ+wXJLOgxScd9hhlpiE
jgNYtK6R9NfUEQW7Fia48PrLoZ6/FDDtjm6zpeV1Kkx2oqwsF9Hie2jBG5f4s/tv
il9xh8mxEs6nUh766qW/Hd+gqetWMcAxmF20B0/hIrFC6Hz6242e986c/0ZJOE8a
AkZVUMDZZXCeNAxKcAHgTRvsXil35j4/MlGM3Qf30G+8GUTDTlx54busa5amMEPs
rp9nWFNnGROzzk6vZJUF2N2posXSLf9HX9D6+SOvk/cSl6vTXUAZeRprlx57PHG0
p8v8qHdGo6csqWXc8IlhMsLvZPYUFLtvRm8zurT+WjsIsKVTfT5LTlarjU8eijBb
av/x7LgN/arUp6Pbka44DCY+wwVVFmRLwxEJBcy+HbNIeB3pbh1s3FJppLaxRUW8
deDklJBGO2kxDVdpK/YkUyfqg2NZys31JZZL9peINUVZkXUMEJlr8Fl6hx6wUD/7
fAMpMkSu2nAx170EJ/STHmMJBSQjmhXqLzCwP5G8kZnTXLcXSUUNiICtnoO2+wWO
pGjitucARbAYKbdfHeJ/mWgPYmmTVuLBXjGZj34KGY9BHHHap3+KRT1oU6VvoJ5g
07HKZuYHvv3HTqxK4Y6u9Dqx2Fexu94Du6CLRwWXzWAg6w1J4tuKaEuAmnjZm1y7
oQh7txk4XqZSo7ELIYkZw0EC97Efwo3hvIivFIjMRvaxr7DDwcMlh3YKxIEjTXfX
DGxIiNCcCYEDXIcrSCYP/NIvQlRZIF/Y5eK2XY+ApWGTDnjNx4ZscKAhRf1OUHQI
vF312yAlV7DV/8vKKhebegtwNdJokwSO612PEJNMz4he/3YCP5ubN1KIqQGmuFy7
OdZaFNcNwNTgU2tUOi+Yfxq1ETPlZAZxALNJ54Wph3Ge48CtoLb6cF+5g3co2uNZ
wMQexzv9T2EFpjIGwS8YWM5XlAtObZM1wHn3H6vy7Q9uwZCubg//EfFNYiJvY8hj
whCRjI0BRwXAAjoF1EDkrwDyOWXQTpWSMnlkPNdIATw=
`protect END_PROTECTED
