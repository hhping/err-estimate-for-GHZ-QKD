`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+W7XNAFMMF8bm75p9DXvOptUj1+kYathT1cdj/imMg2g95xxysujUtohFWU9P3fu
iGrwImzEeqZ1AW6F6eaqRmHbZOVfnunPreL5DZ5oFmV4VB8nkQC29sbghYyxzlvD
B5z6tdmhwrYGNJhyv1tUdcoOq0//7qUweNgKJwrNwiKvbNymMiEhu+FGgl4L8IHi
26qv7I2pHQ9SFNGjEynKcG+j3tDhgy/R//lmgSlrZz2Ti58x5TAXFwB8A2fyRJmd
qRYaSn4Nuba7lPffZ6orNUf2iFIcRvLRiSSsmWbjob+TwnPaBKnGVqbsT6wJTiTy
RjFckmmUyMstjmsFTXLzY/uYancTSJVHNq478Hw2vSJ5ZxiZTiICaieamEXc0LNd
NVg9W2wxftlxjbUs7bGBJvUboFZoIl84XiwCVjM1Z107l5LmoVOPWLqYNlrImsq+
ecRhDUMFJiQXUwiGbTr0Ji5oaDchU9LMayY4R3KPStRidlfXTsctSUiZl7hv4T5E
`protect END_PROTECTED
