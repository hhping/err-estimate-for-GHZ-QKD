`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jw45Xj4URCY0gZnpUJjXnuvup32bYm44Pcgaegevy/UFuDsC8F6+z/XBMhD4x4kr
6cSREPbJPBdx9dit3yd4MtWrsyz5wZY6N8N2UvYMT7NkE1GqbzrqunfXyudaSvYL
wOHtdRn/7QlM6hLfoH/0aLBJZhDx2WHe03mFlYNWTpFG1b8WC4Rc8dLPJUaHo7RY
cJ6DxwacTQcefZ9VJmQR3O8UaURtkSgo7O3Bk0bZHN2+y+sXTdIgwPuwIdZwnpyf
EmmS0DG19Ih4dNeDP17m7Do+onEHY1eyt4WjO6ZijALEUpvanYH61KQH+EPI7YFz
BmC3POER9hjYyKBhFG+h00AKfS9qki40OWRqVI5Yotd2WRyJPqZiHQbD+UR46Q6o
vWbeFx03jmwtYsWMWC5O2XNHzEUgvNW4jVoCii06qE3/txlro3hx5AkZUzF4gg50
AUcZjop24xtZVrH349UljWUIL4g8KPZ91nRJ29QaEE51j2TF5QDgiwWrFViroDn7
YEvgwcvJFOZnFjG0XW28cWxbNmeOwuZOXKE7C/59AURt8ru/k0PaXkgbivUL0SGR
xfMcWYCfCuCdTWbcBmbIpr0bIcexxisxeSqMt10vKvdQSp6/QI/KiNvUEHMDbLFt
j8CIM6eEM7AxuylFZeY5KaQORCkXIcPCY4Q1bnlmXgGv6OQKzv7TFiTGWGh2csWq
gMrSTXALy43suRHCUipeQpJO0pyJI48AwnxPc7nhGPDSEC96ZV5B9PTBslNCVr9g
wqufwlXvjdqCV0EzeU0wKJj28nz+6JLdG4uDIRqq+j4LyNHu+yPnvQ5BWRgFgSMw
IVk1mHLj2yPOFHCGHs3Jk9lpS6E5LBdUTINHd6pu0/8ePwlDvwpayZR6oi7Ge+ET
YAyhDm/x1Mggy0HuIwJIKVn4Vk6UY8kvgzN4d6gKMKXo7K4TltQbbcQxdSlsqBka
c0QKoQY1lkTo9HSs4NO4EgcHBoLRyfIPOVsca/2NGDmzrp0sjWBiUybnjfqWtZUg
w10cQiPHv9yCCPX6RowhOs9/dfwjnsKeOtgQFd25qfD4kkTWWx5Yjh8/Zf1mNuDq
5gpun6tDaEEDStj1N4fmA3fhADPsSWUYavgVeoC/J9xwAD79ZpZjWrZpBdrSzdWx
A8YcCCfHVNcTgFixCMy9NvWBkzQZGEZ8mFhppHDXToP+yA5JWJsR9MgnIdjmbqbg
NsVmdbeH0v9TSdrL6ICRtRzJCcFbo8orLL1jJmaYH/afridZcHcol8NFqAkm4yK+
Y8wazwCzXskDk+zuDCJa2yABoHEHoRySXQJf2JtR7vIpyywTSmoOo1GIRY6Z+hxA
ZGpvTAb2j5Sj2Xht8fCbUDpOfGMF+wOEN1/PgrCVgFMYrXgKScRJ1FhxaANeaBIE
wla7uOyTHmc6uFaDQ2mLq/8jzqfCoMXsbWH9Nitp9zFJp0kNsJOLRn44Nk+jop94
8mQK+MQCNgKklLLodYostRB6sXN/YlZjXDP9wq4sdMLtyr6mNEbFEg5/PhEjEQeP
KaoirIbdaxjF5K90zi/VTuNgi2Vh66eXUbE5Crkh3/OxqLZBVjcGlHiXC8dSxeZi
f4z3P199FyWNoSXrcAYTTX/urbaJbGN3ELJjs0iTtqQfzy5ohZmMxlKJAApdxQn8
YoJMQnbYm9qyZAxU2exKpVIne4OfbhSQjs9nM33igmR1vmfEQap2n7wGkRE9AUD7
qzvm8gt4Jp5TDkYrpFDedA==
`protect END_PROTECTED
