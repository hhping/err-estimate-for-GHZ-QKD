`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YtdvvRHi2AQAgjky9S5lxshnDXvd6MJTQ7zF7lhNW/b4eSgBjeB61cH5FyGhYNI4
4nSkXzRIJ6SE0K2IuCxSy2lwn8T3Qd+mdn4T8npIx4S69PSkkNlXRK4l2wsJLQsi
lXO/EvfJ6l7bcg85EHhcBI9ky1aRvHUUcpOn/SKzCoUEKAYbZ4GufZBiS8Km/oJE
lZ2RLOvwTtyg5j0R0XoTkoh5sNKqdxN1++9n6Sri69uqWREXWTsmBMPDZyoxjAM2
j/o7a6MOSIz99v+Ux2nf0MQ0kFUwdbwhvceEVq8jT17iRFJCrDDQynt066SgTXe8
FS4/IJMjdN/EuGN4ziId0rHFKEvCE1SzUd7wmFBvwajo+zJipLCHSMGOnvEjmIP7
y4CcZVDgJHsRTa2L3zSB2IYpjzWqdyzWdcPJpERj7hyGqGJN7933KFnZNOWJL9+9
LZaKkjIz+kVNj24Nxtx2Ky3NrX1MQDZIgMY+WZGKkmZdt/JMNWhZ9fmVlvs62qg4
`protect END_PROTECTED
