`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uvohm9dVysMCVMUW0RI22F+9qwyR7YGsBrjm6h6rcqYGk9T9aBsI0hNiIrh+SBEG
704I2vaEXzrpCQk3wvpYrvBh8vLzG2iLzARjSVmtsBaEhyE2i6LORfJfH8jjdXK/
VMGr+91Krb8fKXmWUpO/qL/TfRdkBQBiJ9omEbG66JeFogyX+Xl4QiZMNrbgGmU3
kItySsYzpWW3YhfpHIURA+dWcOERklIUxQjMWmXLmlMjAWePJo2Q+BXXAGhxYGaN
IH5bjahaFNYFZjp/hlxX8ppGllWmXXf0almXwxFlDVV7xTm5slFvBHj3C3pNIgQT
oHusJx1Nlwt60Jm6/VROg59kO4/5pq8H/WBRVJiVoz36HgaGO6KGX17Dx95Mb1qD
p5IaRpwSM3atUycxCvTADnQ/OtEXu1KJC5UY2e0l+sdk1RuYDEMhjCrEnGzXrjZp
33SvpUfQsoafBJybWT+vDKAQSdIgXi8HRAqKwyS9Pj2CdZOqDqu/wrBY+ojPgd+j
qBtMVeYiOODvA0ehcTZCIPHcrdAd8SI21l+0KY+vxL9aI/Faxr29BnpyVFx7WIrx
BjlbqMIwI7ndc7XKe7fohbVx/wLiaGq8ziyJWPPYADxh7ggliPl1QahNND//qAey
Y2bmZdOv+rA+KXGCiQ3I0Sb0jJPUx1FHuBXbA3fPJuO8FIEnrhmO97tVJVP0Tnrf
DBACOZbGobGZpXHrqBE/GGBLWwBCLvgdGcT5pOvVD3X/EzqGCT/8Gbt25egzWTJ7
SxCHbEp8U+l7KY9+bvBfSPqC5q9Iw0A/rfV39nVxk0TG9d7UtpdoYqVe6z9QLO0C
cUBIUjqAVKJiAwSB1z0tCzkURGKgjMQACq3adESU9otMzx8WsUtvA1r7/Mc8g6rq
JrIMZghsCu4lh/gazHX7slkF5ZQGzlcI4DtQis6kTth/ykoxXuhYYPhUq5Qa0k90
0wM1fJVitQdJLS8n4Srj+dAvw+D8vUFwzAkzRPZcFc0czkXWTaaPV3Y82ZWDP+zz
8XG8IYbvIXfTs/Det2ZjIq3hfHEJPPFWhFEspwsFqQTk/vnx5xvLXIb9HsSxHfXZ
Jgay9TDxTbtlWF0QjHi3xXkhrt8CQEJYHci1ociqZwhj5n38dFmwSGcGKE5d5aDY
QIppOpNjNQA7iStPuT4F+SlXWH9qk23jve8XrodF3UWDaaHXVZ2MCbNvBbBB88Lx
yqkvfXELOjWR0l0H/QgD8go+G+lEUvDjiHLL1PdImAMPTKz5Mrk/mYLBpqx7sgzF
lsB2OgBtx6AHcX6EkFwveq/f2kbpRs0vk9CaSf3X0Og3YITpefUi/6bbw6wmNYIy
ZBmlZIQfkCD4NNYQ/wqUipn75/dopVc8YcdYmVG2TC0fnEKfDYUdQOEVEIXix3FE
yTaN4n21X+7y6L3Fqv/JbL2zCS8BTK54frE3pkMuxKh68Y7ddvxyJ8W9NZdyg4ql
qQANJGixQ+WAnwhRfe6yZERchY07S8RpQD0o1KLoxM8/TTF0Zz+Fe+EX4UVKcRWy
M74Qu6lVYeBNWu+rsFvuBWw6NASmPg8JdwfQjDPvUZ1UG4bKi7W+v8ut+7OUMNSg
00KnN0M+vYf5b57sxhpgLNSEz13EhEgXnvVhaDGpOrrKtPX/vJ7aCDJxef42ECy3
TB0nsfOsQx2UB7GEN5A3SRgTOzcul1Th+Pp7Z+JAOxsX/MwVnJ1xOk/oC6l0YXsr
CUQ+cTqcTID0Ydg07jxIeRYEwV2XU0UZFg3v347Eu583/P+FnKTwIowD+0682x0Y
zsHqmPljArixQdpzZULOxAxZxesFTD/sCQYs43LRqX9frExEKl6LaIseiR1QCf4s
KSQY0HC1YiaUGVhAL+qHRUJKpcp+ktr/8DU3R+Oh+B/3QUSZAGDEowDJuAyApjKO
l6HxeEIxx89TUhoeyIRMzpXwMdDG2zYBNMmYPz0uPQe6OCaZrBNw5OSFJEkgVlIs
7zPw+zSgOtiAbm0aZI8/rmY3OMgYGHEXQKOt+ye5NROF6oWswHqX+fD4gT0PUE1U
ZojItWBOsRBRO0GWkZ0FwN90GTXr6AtkozqwdI8Xg7+aJeH0WeiJ5YYSuAHSmCQP
ADCDvHdO05mz6xFABsrx2AcKvP8BHQduL1DBnPXPGTi7sQkh6fz6qHYl+Ai2vpo7
ZRRJ901egAmWkfLf8CoXUQAocislle6QOAs4HklgXjt+TbCCSDCDlt0Wd/sLQUpl
d62TXSqX/q/uLJOc3sh9d1LLMcWiDA2rzPjpLLuVKT7IVlmxygVRUokVH37s3B+r
r0aciy/wsWrDIFcwH5Hsk5fhl6TN7rx5Oj8cIh7VGLGdFpBMILTl10xoCEgTQm8I
ADx0s96UL5pqj2HSzMaiAHrB+dt6TYxcIZwXBNi0M8Nnh/qu9fb9aOoZ8iJH1Gw7
I30bzRLRdWoF9QZGa6MZV4IImPoWzojVIWXmooBrQx1nfSz2YNAnKqjLJhwvfJMt
1UAoq5SpZDiH/RDcy9sy64kDRYOpIx6aBEfBlKevOVD7DORLipk/5dN/9B2uUAat
vIdrgJZ1UZ5p1MHSSwVJTlUDrwOegWjzd9UScdMANqUvADTVO3Sf+jr7xVSz98UI
1kNHInwn/zdUTPValDzVMLoaaMMoXp1quVViRe3eNIgpQTNVwDL7TB8UXMfezMJf
PYmwkWYvvawc6FLayO/w6JlZwZzAWVMOIbWqnVrioT1RKju9WpAo40YEg6BTawem
eL/6f13E9N+3Nf08Y37anErtSarxiH8iVfJBpaurL5RMVIckjLIqJaCINnQI8Xkv
jdmRWrj/gLSUnNjpRYsmG9i94xIQpC6PwaA4AZxxE3tAvjf6hYXYhnWwzfBeXHWf
YJraRyp5X4hjJ48uvrgoPgXX1cOd4AgeEdvKWVxUe2/pIu00BY/uxXz2CC/yOQan
OPMNaZHRy9SRAXmyZw/0kLrrYG7J5E/ru//xxe+ROT1X/KvqYVRu7XdBPNDqSWoF
SqVZVQMVxoBgxPaO7JBsdIewKEKrHwAklOGJ+rya9Qj5Lte5bihZ5mP2xNcXe7iH
XkBlJHLw/A6qmzBjkga9u3p68UzMTdrUhg/Tmywu/Y6tUh5bfS4pEryBQwW4HjGl
bkNSQkiaVlogDQa8YB7NlIvcRdl13m6NlvI8D1YlNZrjAZDqAh63CLZrlaq1Wb8l
BkBiG2xFn+LQxHUeOBn2JsD+pAI24Yf6kCclpRxpe5RZ2WOJAoDcpW07tHLb6vRl
16GlKtNQlhdkNMdDx4/CrA7LzXq+bAo1m9yXZDxvqUGTTzvovcCxYKc/PG+7OFdk
Ce/zkg8vhe4nAvTi7fxbJY0FYEB6RxQwgEexbdrhSGTipeLd2OZ4B/UZvKarVbgt
jAm/KOXXsu0cOCWtY4VWcBqDP3CftPmH9FTTK7HdqZ6AtIhjP1CHZfs6b3dGSv9z
bi9WbqAR/07c3whxG2ASMpf5cVi/zmXQYlx70jV2zHhO7dxkiIdoD99resdrF0HR
hy1XUe8WWAjVg6f1nK91NocwDk59KVljKStnWteNa2NwRem8xD2QEJTCF0PdiCDL
0egpgXwZPWXZvYCWw17bun4xea1SJIrnDPsixBuX6LytpikGyI+RReTKjZ6sqirt
vtS3eXN0hNLoz2Bh00cc1yZZ5vEq5BFoU+LVFUBng2LWV7IqJ7sjxMCcxxD7loSO
k2kNoGOtr+cbCciiPhedZfo/SS2dUQ7+mUtgiCa8deooLJ/F5smThBktOvK8+Yy4
vNPX5jM0uHJ7MXlFzCg38R7B9dRBB9obH4hpCmN9UcDW2vgfQRspFMHqc4tgE/+S
nduOFRxkBmFOEIUR5XG9ZV26TZ9GBsVzom26L5AuErtAuuvvM1zKkCvv+xu7dhCT
1dZAdS3Y/FxVdBlMMhs5MFfW3z2K8PJC1QPAVn8xVsVXZtv8ZNsSbT3nmiBUEmme
xRh6kyMm/SedC9pDhZnC7vwh631s8WEVLtob35Ciz2JmCKbTQPA6Bsg1nHnNzBal
DZ92vsj0hHiaH731e4PD6S9Pcgcie5I+XNbA02PeI5a9FBBSni8lHjx1quKC+ONg
STBGEwP4BlOm0PlW/1jYz9/25Jd5DFKIPnDp80uYr6si5aTihgO/T5ZUHn1kaZ+c
jBDNjeYQGz2Z93bDVM3+boI5IFdSk/ED6FXtonCH+nVxt8EdC1rcFlCFg4OB7eTp
nkRcvinePYN3czw3E+s2hAKAOhz12ravUslkBLhQgProwfmlfU/9xq4mzS56ZK2s
83TjglPa1+VRj2r2zb3qtwvXo7YTdudp7pqpxbxRiD88r/5jaNcwBS/Hwls3jR9b
4hLowO2MaI3tyyo/bLLtRGti1rJIIHFLzEY6vwxKld9+ieeC7DAyOFvxvfHhn9Do
nofLjfwPq3ydYZKlrXgtslF0JdfB3wAm1yGWiiWPtd/vV+rmDZBiFXFLf3Id4RBJ
6Xrb/W5GjXftHjmI01Dwvvw6uca1/jb/neozcRnCI4Jz1KfV9okpM81CQj+yM3p8
3mVKtaBatAgjJtEIMYuIuGZb032g3tsRVcgI4EVSnIHfiYD539GbZGYgST2LQgVw
ZAGx6CsJpkfL3bBvF+Ajl09IB8jVeecBcx1D7s8jzBqhLV9AXAdWTYQMVP7ChQTc
o6mo/kkhRPqe8sbWc27U4hPuajfLyd8GAaWs/iM0s1vyclbg1AqcfaKu0y7GVzd5
TQFiXbw54eictKtFWfPHq9Dt76OYb2+9hveTDi9yx/LlZmxLRltYmK+gCNBFEznI
Z0TvyyzIZYNeEKkXVaAulGNiTV0a0mJP1Qs84vvLoetu+0mNlJvx5TuBBaXNocFf
HY/XM1inSrjdZgTZ/488SDi5PiIiY35S6igjtxsxTZH4rK3oUOtjM9az0FnBvF4G
LUFS3pVvxYDAbJc55zQUKeyOkilLlQEx651looSuXipoEYNQ0iW6spskB/XxuKoF
hyjZJG6I5OXOzGKq6ukKOF+1nepyjeLGf43cMyDV6Zgb/aC+X3VfkQtAwc+VVjgF
qZIM8m2SkDd1kY3Mhegasq5UEvHBtOg5ynaNPvpz4eb6hzJNGb8ZvNRyV41knTIs
JMTHckb/tnGdvNsqR/IQFYvG5i+20Xsy5FqkAm27IjCelLCDOWQjUXBO5X9SESdY
tsJIhzwzf/OJy/WrM51RO5qscRrOu4RlvsLfBtc+KHsS9lJ7lzdsKQwOVx1vs3KU
90H6dbgC3Og0BT6ZC48O7rMFhS9gF9JQoX3fgIVeQonrhBc7UF5HaD3UjFdvR+77
/EpAVi5YKE8PZWtHECH+a/YRVl/gKQtiEO0wnDi91gDpdJNdSqmxyZBKhiz22gaP
L3RbHEuHgZcte3czHU8prZmogdcK8/X1TYNbp6CuqdE6rcg6MPzpK39R5vl60b6T
s6ldgt/FJgX471GJ/gEuIMagIA0I3Ag10A4lvhzyiJgUhgyIMcqBzQOTC/KKQ5Ki
bgiApLTxZA/0qIN+vl7Ef+hGMOo7+xriIAJ/s6BggTKJb4intWdKUWHJPqGuJSXE
bywOXAyol2AAkMCWMPYbINNAn6ac2NDPbhSmStWJWdjzvoVUYmagIjPNP51JARSa
DjuBsFA65azqaUmxN7uBVnm3uXxJ51cwgEPMWgICeE3XFB/9CQo1q2SsOe37Hbdy
Evq4mE2Wz5iJrOFuRutUqu5bWoA0NHAag4YnrFX29ceq0L70sLo20QAJ6Ots7rGr
1dBUPsLn7Co/zUI7fGMXmmuYDmIgfWVEhsh7/4P5uvFPtIjsbYxTJoz30iXdQX97
pZCdPHkXL7Ulg0jzKt74u85LCTPhuYdyPPLX784EsrxD55s54Ucm755qxh1tfZ+R
o3iT0+NIvYsvLrWpNB40LNuwn9GUk5x32DptV2Rb7iYCtWWnCrOmbpNQvDNOdSjB
YMExzs4Fz5m83Wf8Fc6gGVMTUmgNVlgonioysmC12BfbuLjPZog/njnmCUUedeLk
lQoXyN+AyUuRNFuP1bekMIdVgmwOdU4s1dTvYqZAVTucvdjOYq83VhQnmLDJSry6
ZqlKVLf01Q6PqFfsQhpaMx+xgYVgaBIgzRrsVamSAMlh+082O/cF0jYRNLECLFYh
VE7SD/SpGg6a/wDbP4DB8hCaD7lNcjnFI2TRUDjwnHsp79uOH98u3mgl8qc9Bpjf
esCEXT3erIvYFm034BvjfwandQVQZH6hsPSuGK0qNfSD2+cQAt4E/NTEbbaF/V1j
JyiCEModVDKLrrO4WlIO5vNv6DVCOunvOUs4nq0baEiESvn/3I/cXEPfTTSpgd5y
PAs6/DnWdQwztA2qgaQ71T4kENaWX5NlPZWBz190ZIdNh8MuGi5g8MjA6xT1iJVr
KMjijs3aE05iqfSvTFHEe+SQG3LVUjysiwo2xmNmY9fv9ChM89/gaeTkTWuhuqqa
LK9o08/5t/u/ghRCIizL4Zdxy97XBCFh/fzT6B8TpWycYcRVpaGdRefZsvRhHTlH
GHUQhpwUOUqzOTBOcuR3B4mtYZZU96FyabUi/4YVc7mgET1Rc4YWvFcdHX/B4Cbu
VZHL14ITo7ve3sor/9vRVFqa/CIRz35YjqIQJ8kJLRT8ZEoRcz3kBGovh9qTDG0C
A14S0l62Us/US6Ct0LOPHXUtDOmg3KiKvd/eiScl3YReVdb045W9srYS8CCe0qy9
WEVKYJfh24QhWLvfFPBCZ/8LCjLJuAtfb2bxPqBXdD8GYAvWwwvtxyUl3HVBvf7u
GLMvkPzntFv6TjYusovtuMYs9xkNdEwVtEQaxC/aGP6klWVKB2drhZZ5bym/hm9V
QVzOql0WI5zpMtyvnlt9A7MqSmq5VjAmEQbm/Tsh9HKI2ud6hzcwTzpQFSSaVljP
YWVTEjXO7kiy5CZQAfFBp+kamKAVMh4LM6hojsc1ul2u5cTYUXiVMR8tr0AUKgMF
406DOrnBPfb7mDpNEdhB4yHGibMhD6+L4Av5AoxKaM2D91IcGC/Zngv3HqOuMCXG
EkMyLvnKu4oW2a0feil3ynCt2tYMl6G45boAgv4kObULXQEm/AEnNsZW89MH/cA3
ctepiKGPohbxdCrG18Ddfh5dZ989FJT83SLABcAAzwQFnJX4ubs1VRUn9WGywCO9
NH7ReGq9LeNqGY9qd1IKjuh2s34IsAnzvJY1BvMMlpVVX2cL5mupF5NcWIX7O5hS
g8zjNVX0TUgelcf3foQYLGmXBITPfdWDZlLShO3kpiyr1gp0CkljLfWGKkOHB36q
KY8m+iKaoZM0c253/xrhUN9qSUPnC7870fs8HcDpkCfrTqbkq8lfhxMtXZmS3/gX
npSEs35ykX50oyyy7mc/dkE25D4nn3VCBJnBeJfLngApl0rhSdILdo0u37YP7yPh
gsem4uWBvkWsnT2zZ2ww8cwSWOWj5+L6Wwp5UEBAcciLKi37seaT1okwbQBuPwCQ
GhJwfRSUebGCFGFAMwSz1pQTrLv2869CQ5kjvWpmY9qBivFMQXmA8XaRqv3g5n3U
GLuDeb+KkH4yYwpg49o4Fz1zl6BSlOJGLSKbcLxTTO1ZjrqAUrZojCGCEfa9EnTv
KtovdgogqQWtUkz4arw3mSJnnn9Mb3YKyyXTvU0xluoxLP4nvx9tbVj+FfC2+pU0
6zAoCV0+PH0BVE0r/SGLpJoLDo8dl8ge54ZI3RGpF+/qcTlZLAOTCpjsOWYBw9JJ
8VRPTPYPwljLU2icLAF+KAHlOSfLNkKaNZbDbzI8PQG9vqAX5Tp+4Irfzx2Qsa95
oTtv4ZS6UL5X9bANdG7Bij6aRWrg+JHbnxG1W0RyUVJfkgNrMZ6XrxO69F7iG/rc
KMOzb7UecYTokZHT5cGUq7p4q/Er2gxfZoUPktT3yfJ/cHBGSTJB+2eN+w6hWnRG
tu0dg4PinKYG/3/jEiagUr06NraSk6w7qrdMkxZMxpvtSH60Jce8S+bqVrJb3N5h
mISa9kD/KEJxGZUm0eNpdtFQzNbFH6AKZrBDRpWDGVsTDoleolbhBEj246PeICW/
A+VqEUWgnLesdhHNY1dtnmfBuCyQFigxEB3n2FmpJGGh7L6XcwqzzgwYMwpPeieq
ujT/gN2GEXanITXAlw+13JaRYCRhRFRtutvAioberBqoWaTTZ3qQzQclJTcENeWs
lTiTTKVACDbhEjU55fECIr8XvanQaspxrBAJr+ci814DMlANAIvEH8lnrp0Gip4+
YAQaGPKSPY2ukG3/2Jw0oj+NQBevm6ZvHZCat3yZSDYISk5Y/+EasTFvefrL360b
jkA82qhAna0xpL6uTfZejwuJ9Fhn9IJvS/O6incaOm3dLzkmu1SHDMBaC6YVy/CV
8zMRj8f+r7TC/hnnaV2rYV/w18DR20W6xAxuBSfv37cqGHNiOCOonYTxI1AdVdeB
pQ0WSQdM1MDqVeFt1Cw9fN9wSyMOFPO6v8MXGNtcZfIGmMF68fRORRUlGcPaSogU
45nBmhxWH/PEzC+PvGpzFXK0i657QgMdY3bN2ED+YIM5/qkb9KE08+acyKcopObn
JTTeCjycUrUIZ7swd+IrSd32gh+MuWrASdirq82cRdDOq5O90M0Sa6egeUbsEB9v
oNlrk47ZKarsu/CHxqBJ+W4wNDjXE4AGnXcDMfAvWW4Xxds7ZAcXQyuFPQ2GL051
LIzNUULGGcC21mZfgCjKr6EpSG4N3k5deC8XFvKbPTxEtauMZeTNB74ldtHf1oSV
u5omNxujwClszW+6/BfonK51IwWlTQBMCYZKjemLgWSsb9R/wfWzVJ46WDEASd4E
5zpBziC0b5AaHBqjUW9+1U+ms6gNN7+e2Sb5MOGRjZT1Pqb74B1bnzo2NxJ9wt+i
IHZS3j0qGWePWtkMeMjEHpNQf4trrZ+oGAQ7F+LNI8Fa7XmD7byv9KWsvgErm8bq
bfxngxtJ4qFDFYBVe6GhqkjPa4Nv+iAJH839nT5ayPnhWWfqM/vFwTaBDMJugXo8
enqsJvhU9EPJXfcoC2YnuVewbLu8pOBPmHl0wPveMSrulAlyJxYkHhJOTamVzhvx
7QzfHbN0vaA/wPPxsWUlc0p46UcK5qSBe1+ZcQEUYBNiVgSGdrT6tTpTz7MctBUP
cIvRAveFfeo+b3gwhXVNHfjnZ+59usRD/SY6hjTUdZSyMhKvJc7JE78mhKFbSbyJ
VvHThKWAMfSIOorN3AXk0brK7ljbiT5fbm482G8EPqnaT8XoHNpL1hyue6A0hUkp
CY+rJAN8As5e9QnJvUCrAFjJKDob83dN0+BjMJT+SHB1yQMkpX7vWrOkPquo66Mf
yMd1PSyxlS11K1u0LSNRkr/Yi5X6br6nn3Iucjc7rpHFDrFXj7UmpQuqx0U8L5j/
x3HMeIg53kMpoCLH41XVmIDRS1y91yuSMNG9LzjZo/GP4QjRS6hMsfwV+8627Io3
t+1cO/jzw7E1V/yh7Lyo2qUn88JV3rFDE9VQ3IMDpop0iGdFqdqbVPKhkyMGt//e
3H96hYsP2RcGFltmPlT1GtSh8ecT4p+OBjKFmF/LVW98TNfgrIvuz4e76sJ7mCmj
IIr7sjXjTfkvQaX2R58rOLmbq0RMCvx6MQN7nh3Usvn+8f8iamQL7iIqt+2rwDVI
D9aiiUsvRZ3qNiiJb90b4ZxD8yzLJSXSJB0C9Tnb5Fit6+wH49l+z9CnbK2Gdadr
FCjHBVgBoiO3BYLK1nnMD/YW9uzELhe74zAOG/yvWnWKh7u27CMco00jfG0aH9pR
R2seP/5p0L9XkL7rCRvLe3MDIOeArhkOGOs9qT3Kn2ops/0j2jOWkJ6hlr6pxveV
v0GsQ6d4kyBTueoj5opnp1lGL+Guv9V1SAlM6tIKSwlhlSxvRnkB0LU6hRkTALmn
l7O9y7Kq+bYmAcNjzKatyC6qZjtK7BrunQKGPw/kwi+i2K5eH4EwfL/zCTDlbicg
9bziUbcD7mJ5LH7sgOZMXkIRduCmIW79+D8EZy1dPK+qCeSeezz+7ElrQWBiQ6Yr
Ypbb8NW1tgVVjFxAwlxT1mb+4jSjqe+mhV4qD2LE2tNO0TGbESZ/E0OQpAnMKvkI
woZPaRdJekAD+Js6fUajvcQLMn2Q+N/KANyA0G0wJcrE+r+o9qLhxxtnwu41UJS6
YhZGw1roGFez7FxCR1+DgBavWWQ7fEGVA1rlH685OV5IgT2WkXiERxDAu3SsGUmu
Qv/dqw4vzUcPSs3dsmsQOhYIzID35le4TydewRd9ed8=
`protect END_PROTECTED
