`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJSrt9DHmk/T1RXxl1dh5/+BvTrKS70MVoKL9Erc5iY1EaPKID2zErxQvkEts2Ow
xnJJ8xHVlMDNTeD8Uw621nSza3Zo41HsgFj+Nq46BpVZWrxXEik8dt5MGNiCEKuP
dfdY2rIg+wuxYsxdKsKa149Z4zTawA/k2f3JvTVUOg1qj7XZZ7qaOZv5eDUt8LXz
ZHbXn2TQX3hqu8EBG/d4kIV/uDwy2zkmqgST9WixCVt/Zl90P31eojuMIPvCXXwr
KO/+8YBvdTdjtOwAkdiHYci4APksrSLgQ/cPz++OIKMwTEVVyAPw3WukCpvANBq3
H4WLFpFtG2RhvaJO0wU3FU1dsLYAAgf5L+9QVIG3kGmP43v7oWd4asekk0+LQBT9
bUhr+HzvF+0bmAtga+Qb556EMHOL4VjoVvd/yHc/o8p8aszqxTkKbEhJqyqXRqdG
jEElqkLu5uDOyfP1/0DeD5iPMXXPg4ZCVoBgkz0QNL+Ri9ANWerqTju426SGcdNr
zfDAIIyNLCCKfAONMuUy8Zh0UEtFGyS1HGqls/QBn0pP12CoBH7xKa9m20NHeAMd
eqVrCwKCfgUkU7fNvjq2bQ/eks2U95HNC0En4zC4ohpBtfAPxOCZxiDDBy1zlqcg
vQ1iqQHSeM1+VQ3qqqAIIbYvDEvGtl2KzvBtqdQx7hqc40vWgXtKmJtk4PIXRTQ3
38ARQzr0nWc24qomG0n+R33WFOiJrtKQXGu9eWiHBh1cS6BXDeOnVfIXnt4A6Fqt
PH6HcNCzJuUs4Gg6vZxMoXce8A74qm6tjMyr5KQ/S5cBN7gU/H7Ntr7lHkykyanG
`protect END_PROTECTED
