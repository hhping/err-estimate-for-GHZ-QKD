`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFNSfx1TYYRGzISw4YuTyGHl77yLzUqtv5HlHHiLCYBlmcWR5jMp3fbDrwwrPadQ
NDT792H0IlFfs5UZwVdDi0rBzbn5EA2UYYdRcAHVNtYHSsseUObWbBCG5FcQq8rJ
d6A1vIHXbac3S+vyqgGDqxHTo+ozxCYgchMKpP7QEw0ZI1jJj8muBR4EeedkgVnm
HqpcH2tAln1ENOZmrq+IkPwsbGr/sj3vE0jbBIRnVQLFE0XewE4vK96yWobpuoun
wV37SNQS4v8JE3Tt4d04AQE7nxkqAe7+zyYcuwB5d/TUsDVrwzmvq3CdYLQa25lV
/qucau3WAF8/pnHV3pGWVtSimQ3GjFKTB8kXnMdRpHvfYd3rx1oxvO/M27CmWR62
JSK4fHMOokODGVhTHgYXht4DmCmsBfhkab7wmaEZGpQS9xiedFB4Uh3ZP2b+kVOw
Ov0Kr7lGRGqIIaNaP89LKJN8CyW1VaLkuyXLBvBmfsyLStxlM05tFUzkZ2M+zF1F
OvNwW8tjPjpqQVeG4+HotvkducGp8lSTjxBkkSzX4kkE5hhNfscivs4Hh3rAPZmI
2amXyJWX0vWPYcqfOA1PL3+lvC7sEmaLBHzMwhC/UxYxCiB12GZ1Maek/xzeVv9U
HhnF+9cGZUvo8mEF7WcOjaoWFO18Zvd2hJNbutHXVENg2jvkxlgQY1nFs5a+4DL4
zms8yQWu10HICncwgNLs+pTvym3f/Ok8WiM9IdmZaKuz/mwBDWPyRMQQoon30nbZ
U7KRYD8yh0fWZXUXZhN0Zb07yA/AFZqqJP290R9IaoJMCfwYxzv5dSU0oT0WHrzO
GqEDCovmdP/I4Q8KiVVtag==
`protect END_PROTECTED
