`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHLDw39lPTRo340C4z+r2ArJvmHDsv3BGhplqmQKthbOkxhANyihD3hd7yIm2MPl
G77wQpXSlltTMR+v68A6OpqyjLmDWLiM5UvyvZaoPoFlIIGojzZs1UTAyn3YH6vg
0kmGUarYFMw2ciWIec3ltKUoTcZ4SkkQHdfrh6mTY9OQON5CqvhhcFBGTJnW9L+y
WQ/jty0xs+QunltaPGL26eDImwULuv9C9Y9TEyaWqN+9xIDtGrGoPguusPy7AJQ4
24rF7g+qS7yEsc6lXiCrO3dJ4Al74Pr5jjq/abdfKzWSbZE3r7mDrm0AKbi1jjhX
Oy1rm3NdrlqZodsOFRSDTmke0RVkYL2wIdUwgTH/peBfrMNCMPgx6jEIOW0fEk4V
k3ImgsccD9MJdDJOHgnbNHrbjqDWX2Vk2LVmCdHtXpRb11AecLVq1getDUY3cenz
SGB+A7WV4gAUDyvESf6cKqbM0bKfHJ3JOwmhbmP4BJOFbNVI0IWO2UHCvQegkNYh
P3wXPIemmpf5FVQ/jEIlA0Iqf5dw1rRCKkB4Q32S9fV6c/xw0wy7WG0yVTTsN8Nr
J16kwnXCFZLU3nS5nZnM0QY3IvHHBzvJnOv+f8/pX1+sWjcu2s2qpPmmrqoEp948
Nw4kuImXLGDsswA7fgJAQzpb7ptOmQfRHQ57Aw2rr1H0ClxHZbXj7nmh2NMMD7Sl
TrMZjrVXYf8DvdMCi65SPIllLECqyze1nRLY8Y7HRX5RQzN53KLbF51Iz47MY8Bd
IrFm5zfDcQt+Hj0RYYGy6Q==
`protect END_PROTECTED
