`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jUVM25z1XBlxu/3p35VSJSaf51NL+wEuEZ65TwkFf1Nll7Q/qtODFa9PIu0oaIf2
UutpGhXNLFjMWBdIWohbiVOY8E9BNeewTvJxZlweStYvow9gUKgXmvj596oO010I
k+4J/2VkKAHICsctdhZ7aPZpjY3cxX8TdVTjsBXSNIFzeZFiaNNr7POhoJi5J1Yq
vjcpZvDgx++wl//jJ7fda2+K4F7ROxx26LfWjaAIHD/YZtQKPn7SXJDge2LNZUoA
oviE/JLYQwfYR6USO6rq30OFclr3H08joLgtODfHJ8yqnBI+Wy2DxlvEUGXqC5W4
4wOHfWj8pK2X5pHMhyJuRimC3+zgF+bcHyorrDinBn5G/MqQgWzTb277syw8QyHw
yhficYzFO0YbN3PowsSr9+arLrcbjI7k+1d2wb1IaUgfm6PEKDGr5vob3Ll6hGcT
5iXZI7QKbRlEfRpiKV8vQjUHRT6SA7pi54xwOmrhAU495i2TpnUBHIul0RD2CpwK
i31GzlF1XdrS+7oZT/EKT7gPDwtojUrbykf2vivDgwwt3+dIE6mdXpuLEOtTSupE
XkMT17hitx2q4mHg0lvKCZ0OQkbwT0sGpiF7tEkCcs/rJlbt5gCLiRD6f7cOSDqg
5vL5+BQqdsZVqcaJ9Z+5ismZPIhLJiHyTIMyGvlN5kW3a+Z0ZwZeG1holt7Mz7d7
08Lu2ULmvao4iJeyBHlr9ATozdEWuSz7c3OFFiMqQPc5oZ0sZltwVKKzjS/7IR8P
mujoPL/hJUC2YQvkQrWhLMsCU3nTkqUCGY+ZE4lCdsJRw079phDeS5/59ObJcH6T
zZm2NTGCTJAeSbG7uAuMsXSj7Nppo2GihpsvKSQhdI1MPsYdKwIfR9tHrfkHE+k8
9x1G6vIx/+xfBXaSefS+x8QrhBuot/a5RJKTMZI7p/s=
`protect END_PROTECTED
