`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYomSkO64o0sCZjea0Dwo2m4kAfrk9YpCfBoYfxkZC1YzEPO8zxaCjQ73SE54zFD
KXo9kcjquwkOlOY5cMuzYXGsAAwyqjZwFMC8xq8IR1spw0EWF4xljAD2ZcUNpmFz
Iz4sP3cVHzD9SAosK9KdLg2jv5vCW3Gc9frTf/OQGWbcCJF6Hb7TKN8EpL4MuD6G
HV3GQ0Jpjtw4l011axS95rjEFrvphsmY/GjFYQL2a5kG8f4+6HzcDMUJ9HcFpJIm
p8S7897IIRjGeiHhKMpHnbyNX1qjdbFx7siYXsHnaeq2AYwi/94X0qjB5Uk//5SZ
uj0FsfX11JMuAZ/2IYTSGhD3/LOZSzd1r9ujhwGfvPi0x+IngLzaFfZ7xmO/nmpD
SfFyUlyjXVMNT//zW9iWN/g71GXkkKmN3Ggpd3INzTtDcJd6L+Q/vGV16/cFxaaS
qGDV/urj/ECJN8NVJZz8jbUkK9wtvtM4WiRZPSCA80rbINiGqGarLPtPAsj5Q3w/
fm6rrBDd1UDCd4NOhGNt0y7XH26fA0x/tu8fOL0/9dbK/U59uYZmum/WeUbucOvs
KpIM5cjwRXfb/C1votF5H/qaOAPpzBXiKn9My3j9BlxhDduJUw5j5qquXy80dddo
85oNmpuEz3GB5C/1FK+Wjz/YzJZymSYzqqql8PafFXcr2CS2NOgQEt9j/4ULmQS3
/CNwtHZobm6yXXVkUNyK64EImlky7LuNexGws3GSOqJTAjdvpvRl2eMGJXFDy9xU
3fNtnHag0FkBE72vN8I4br1yVrAjMiBItkgGCFwJq2GG0PPYt28OzgiUkNnjxg4U
op2ZZU5P1Axn0ZmTpOaJqiU7MVAnF+cISjqXMJHQlhzdUx4+RqBQZM6rrUKgDtvv
9pI8nGsuJ0NkPUX69wLtJ5FhdP7yc1cKq/e/mBlH9AKHzDVmghmQrNE7D9MgZQ/V
nasc0OjdVOS6PrBWNKlHDwchQt0Ryz0MU7Q6f5xROlceSI2CD8oZJs9jvBUHGWAo
KY202fJGImvkvi9EZIOS4E7N40lXPvxjJP93cpZYdG1QgXX1kNYf81CqjvHmtZLM
uoZ9rl32KgIhrX9lz1hs5h2SquFmJrLUgb80ggmlzLZXjaOLwkciqzIZ7okJyDp3
5xEe76iZLyh9ND1x05dBQLHg+4r4Nt4BQmWM0BVl7XOaCONzbJyxLVHWiT9cUDxH
NqReSMYCmpIacrkQN6O+JkIek8aXehvzvJ5yoga8piP7TM5riZyDyPen52d95wgq
DKLjGqjDSI58Eu0fXTG377JAB9xz+FP89ID5aeLCLgxQgYA8JpipgNjwffXWw6xM
Z6aNMSN+238TuNTe/S3+NrAOZfQihJPsUHAUMlraFdSsM0hJBnEL3I0aTifwrtXc
kxXNNYZN63papXJ5fB7rTCAAOabgjenFt5qRGjLsr/VPYC/+yKvDg88ECyQkVoKI
JKSq0bWY2qtILQYk0F8Rcfvrttq/bpUNfamrOIoZ1tt6fZwQciIiTZPLARqC8k66
vK83ZU2T4xgLfeXBGt/YhoqnBgINTSSfzfh7ziIFp+PM65OmnzAdSy3+ZgkxkoW/
zA6/sEpUUOIpK2WlU6n5BaBWJwFSRMvkq5Vg05W5n0ETFNoevBKPFNZmuyYNGXBA
9PdMRVN7a8oPyyQmZcXg9vbFSYG7W8ycy7cjp8ASO2BSGntkXeSUyEt3jgeStqqf
Q2wg8V7HKr5Z3YVxjMk6vat6dnzr/TXDsLEPAgpE/oza0TjvSCplVtj+stShjOIo
O11iGpSFsCSOM2x265ylUXOoiUkK5Y1M5Q1ptkY53/OYKEr3fwV5zDZGvKyX3mit
cRb7HS28gyHxkRrDEyQlul2nvnnvZa2DJvzg5oCh5U/VF0jFoelULHBIHy1rA6JV
zOThCLo870XNKQ68OSDVgwYIBXD6FeHETDXMeelQ/5fHQcKgsfQHZy3aUi+X07HO
AOPGqBihy7IcL1qZJZRuOA+WPoxAym0kK0EXxngwZTPykmXJWMAiC4BemU4ORWf4
YE7ZDT3Yvx/gU5M8AUG1P3HpBl9NXipsAiEeCQT8mQ31ek/KBMY3l3N1PJgfkgFw
nlWCghz/XR8xjA8+cS+wqSuXEmiSMqGTXeOXB5Ry4A7TIxJIPF9tzt9Goh/1u8Hu
sXFKmDk7VPCwzchSLUetZ3z2SNKUGL/KekupwnILs8vWfWv9HXLoXMtCujjRdzM/
eiqwHxce2M678MEz/bkDJhdAmeYKALpaFf8qD+0iLRxAzi+BS2EKIZR5wGOJSOGp
PfWQZm+BrNZluT269av05Hdjh77QAZmLZaRe8lCgmSOh7RAEYOVrxZ8tXv+7+KSF
QNskxx03wPX5HGnjSPtAg5He1ZBq+YfPd6sTCrNgo/9W9IyQxh/ZAhqYaqYFhyut
QNrbo/Cw04Vo6dDbRarQOB+zp90c/eLhT8V+1MtfsMTFPk11+sDv+u3GuWw1NXNv
gmM3pWY9i6HPl+ggkIemBb9VCGLd262mEFB16ysW/VM3nXTJM35xlIfDUuacL7NV
pfcjaCyNyQ1DGinzwJAnsERl/F0owQFOTi86o8ZAdYFjJM1k3QD6Cv6DIC1WaCaY
kQ+JlkbNhSDOaOySNvx6RAUOnebyMU/dJSBTLjH6tFL2qx6mFQ1bjip/7dg1QzAU
+lhYsLuy3c4Ygu/nljrpePD7/XIQVQ2HrzaNGXLjjL8HTDf9d5z9UZPxjBMsBg/u
rAPn+sBsVhr/LPNyOJ6dxO39pIBheip2TF3JmCFwbLxRqTMnB871CpX4RX6difjt
cH/zyPEU2/3j67m2QcjhfPLneLC6Xz1wk2HbJrhYxV+1SVqqNax4opsJc+IsRTmU
/WlpywCBpmPtNAKpWYHjiewMIu39gaNx2+WKKLwPv8UKU9qvw8tAyCLkBNF9oGWT
WtUb3uA/4A29RgWkYLzKp22K+5h+ozAwMmVo/tv/yil+P839RW+lRn3c+zWd43rF
xhdjpnuHsfsxjabOlWOvsyxoWwIdvFJYvooJznK7LQlYGzI3pH/qxhaDrd/tIAFv
d9CiCk8nMLNmFUOYwJNXkIRO1m3f269hPs14lDy0KhtpNcH2z+4TPko0EsSf5vni
ZwPDpqG36o/oFV9ok5X3V9Gy2PRWKWTQZPwyRyzEeslOdyqar/vL/jMBoJc5/11i
Nv4CZ1Bwg0uN+5gUrHFh2xfJ/zSuJIFTBHxDxYrOUWjfX4tjkm6P5jt4D2+LyqpB
DkCR+Bhm+HhhHoaHgk64vuGsjYdn/6HQyWAgbXtfgVBO9NRmJB82i5CkbVn7ce9i
AT3lgEdUlOF7TuX/4dn6PORqq894NNGWlbo1gNRm3K3QJR5cPxTsHrj+274O0B3G
5AwNGXOLIHQnsB74eAEYoZHXG7hnIhIxaEh8YYxmlKqydg/9aJMDgxAreWjtcLLL
xky7FMcG9U+Y6HyEzvn7zZlMry29ilZQEBdcDEEf6oAoR1FqF5mRhCZpMFOuQ5k+
HjhA2UC+j+PrDHkf0tjfjFYktEq0AXl/JaaeIDc2eMCyAlGxRkSsgf3aUw55SlL5
G9cNvns+/eTrNS3A5VC0JDXg6HsPmDKnE/CLlPkzgG/RE/dtTip3DkLdQ60/NJjd
9gQ9/RUvy3Y9hR/pUjlZQsdlU4cyjxJSu+4kO29A/jm2Im7RWgAHW1OBm9FMPxAj
/7Mv6ai2G6OX2v1JNAX1mLKcoXNyG6OhhWedMhTtP+mUrNWYj0CjIKE9HoNJhejs
WKhgSjC+PrDR8RTZg4fw6SK+afnRLzPvUJkuZGZbeZW7E/A6MWnGEI19ZaixdRgl
m0MZ+7vVwceQJ6LdZbOwHad1GhvLeoM00QZQ/H8nBc1mQBERIzVdxktg8hOO26FR
AQL+iCFtUgjgmYIogUAxAV3NUDsETHGOP03Bo5WWLam5rqTSr5viUEhWjrnJbYAw
0uTMZ9oj+9CmUVXVkdptR1mfZdNno4Kga+MLe83PiidfV6ZpJPFGcnUjHOvGHojz
ZfAnc2b3HcWrPOGswDGOhJXo1SpFlzc8fxiwm+dSaGrH4I1jDDr+93BahzFKWwYx
YqGfOFmMvyrIGaRWT6+/UpQWD51FgAry0DDFPzwU0l9dbfN7Phlqz8GXq5zaVOxV
EIGHRJtTESy9a2zMA0F0jgVsxxmLyZ2x5s76Q/FfB7qTgoGx90jOS8RvhZneU5+C
an8ZHyxa66eF5iVFy4n/cKy1WT0MUedbg6tzMQNt6BAO//v3gTtKKBN9fsTAs49j
NszcXMkvns5YQncNRTFGJ83huhvx+EK4bNeCpbV3APBWP3phCCrFBD3IDWH1CQPX
BuQKjm24XPamRJ+Id5Q5GgqJx2UYZfIuehb+/qG7i4qzmEaqlrLaHwu4yT+g0zO+
BzmTM0+p5IQUKPL0DBQ2EbhpNcgb+rIeHbr484y1/OPVZfkNe5BtmcKzfP7taRU8
K/9ivgf+avcZLNFOZp/nJ6dT4cpyDaBdnfc9DZaXZipVYgkAlWyryNdIK54WrgTs
46d6mJ2OsDhPA47tFoUSbu5M0cUX05UYuTFqLsWy7nVdVIVsqeHx+dGDXMWvHdXy
M0YIhEVtHZm15OewCM09JakM+jm46qaozwy/jOe+kX+aq7nkyLuZsN0/0nP1yhTZ
AK9wRSpiEcNwCE/AhyQKmga8sn6EC71Sb9OBsoSKOg4YnKKzZIX0syeWwQZIKQaD
BxNIF99ZQ9oPUVmpw09Fk8od/dwU/m8uk+JdnE9c9fXm3aTq1jA4i5a0K+KW6kb8
+DAw+PtpnzGsZCpSkyp7C5M7WTOjYW++kmlxH0FEtoQFb34Tjer1FLFP4BgsVbGE
GG65DgSeNDLh4HvJi631lsD1T0Om3HQQx6ubLGuckmI=
`protect END_PROTECTED
