`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8McWQt1yMHlNJxLDoDBfxfpqQRL+3Zqxq99BgxI+r9GQsaSmq03O4cihDsQPEMN
eSZbTMFCST5mNMvGQrkb5GfSswWtxZBy4WEd1FgNzEKipZSnmlI21uHzmMjBQRjh
639gkJiBkfv7LpxDyUz1L8DrbuOgeERW7OB5laMmIdDCiU/msKypjh/6yVUI2YdW
zaARXnea41MB5usyhq34iihJGqxB4VGk6UyffXtIRXKcsr/vaUx607J36eNJxO+w
okJHYRNRIKvUUhiN1dTmSyzNsuJHf8sMAVbq9hnTFfLhhaAZq8jH/Mn+ghfnwSGg
oIcbYp3KSFckJr8ds0NePDr3OMI+zR3GzGQr7NyNMWMN54MObC2fRDAF4kytMYjm
ynwbhX5RFmoKBrmrnq6ZEBHw+GFL7cO66Bq3FBaIfGsjpeWGHS6R6uGOT90XXL79
BQw1ldCQprLQhznv3G1EB/KCBCmRVvZ0BGVzviH2IZ7tapG78E3e4CdrXzK/KZ+l
pvuqEn+/NpcS6bOBXVxv6yqjzg9fkNZZbuaLbhnjOV2Z8CX0hhcj9bT7pNPEg9zf
kwZt6LppFubr2E6J689NLnrSnndal7s0jRpxLiMXlVyMkRsh+C+DxSDzsEt/Jqyx
vfwGmIPYhLwBWY1zGPBGSw6cqqrm63EXLfUVCfxuQYqMKG1otjXH6183WrDLYTwy
ZweBmb8ta4lRZfoc2pAyVFd4ynut2RQ6j3gUi9RzEv6lngJxT1/tc0k6qIrCkP9L
9Tzu8iWKVI3QNTX0DPkwmskLdXGVoWCIgU+Wri6m2bdNeB/bHEKnvcubRh0DD878
KXfofpZ+DKpM3qfBCcwGjBbmaApnZHuZBSgScUuYmSSkQBS7nzB6cYnFX4NKksvC
GpYyY9n4eN95eIMvUEfYw4cRIm2ysVlslkxBhs4+n1o=
`protect END_PROTECTED
