`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJfl89WXEHwxRIxlNcp2uHXljodfuqaZIHU8YWqgn2Rn/9NfcW7hwI1xhxRkdwlD
A7H91JPkw6oYCOelMZl1iZ1KHIuQqicBomVDfbmUKQqQ+uNU2kWFrbCh3+Lc6LSl
iV1CGeKw1reQiLXoqYIuoVyJdcHL4YtQMhf8T4FkiLVwpIMyHq8tmokO1kZ5Xi/k
3POe26K+8uBfEEH08xoRAY6vEgqbCN1TgFQhCrJT4kde9b3qvwims+Rq8MnYDNy8
WNpQL16/Gbemqhp/T6mKk34Kt+Ds868vh64qckXZyAOy/VvATuTavHKMrLrUCf20
S/qHqZWWIlBPv7lfzMlIhIim/5X8a0BCJygP0L8jyDreDc7DuTzq5X6hw+XlMm6F
EsWyXly/8LGs2jAPaofeOHgSq0ds8rd1ZOZBvtN2DQwQyPXlkbtbi57N8wALQhcQ
4WDJE3H1K7ukDSzj+/583g==
`protect END_PROTECTED
