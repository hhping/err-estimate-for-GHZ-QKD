`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iBGczwc7VsHhSGr6zquxbLjppcPjjxzt6/mVQeiJVUOEvqsNKTN0Ue7lHQZ0zt54
kkrHEGSD/MKZK3lMKpWUyO9nji6+rbyokZVZPWY6OZr+DmeOioaqXBZBF35LmcmQ
3ON8l1M9QTEOoA9a6ZtasKpWCPHDosGRnGYJ6WEfkFuGKHUP92bCMa9ROIHbmwMU
OimlyMqZVcgjlmpL/13qkfYGjQwPnLk2OMsNl/jInqoWqfD1oqGVsUmOTExci1r4
6eJuyNg3QEDwENOaisIZam7VH5WBovCfR704nqe1fQsorHKLovS7LajCSryB1anT
VzB6tJfdUrGOZgp8lcnariWEpnLoQUALEpACED7jWNN4z6ByJECscxT+bFdJ6k1g
Q9mlz62PRgybUsiZLsCHFjgpmJG4ToHND/XqqKmZJT4IcXtFh0RQ1JLHHF9CMJhl
7Ozw1ajZk3wljneuNA0SjEFtWSeGzgTwSM1GSSdtDvlEi3VxyUYfetujrPoFkQ3h
qKrJSr+x9YOiY70ls+prBDKJPzrNEWSUX82d4nufpyRDTgXK7wsIxpP1+rMMlOQn
a808sjO+A+fG9pZCABqvj61/74/NFo5QqkQWXz2GQD0/7vD3Dil3kibhRXbu/JWh
QjBWbg3E28K8k59amB9WZxp0TgqGpqtM6tc7uVaRpF1y0Djgg+DFpmb3friedBA9
YqSz1vv3f2wM3Wu1b0QmVb3YMlb6aSexq/iRIm8qPiTzHYjKrmGtlfAcbSEam19U
PPQSAxmTv4OZigG7sLUe7fUAGNxfAlIlRiiR8xG4ws0=
`protect END_PROTECTED
