`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ye1uag1AkH14f3HGXYh4mXT1EhkvxhIKXhEX4+cADfs+GsuU+lMK0R/LT6YhJpN0
2DrLfx8RSJAcI/Kc/a7plRgbvkzoOeOzByBFbFZs9RVruqixvM+t+G59mDld9VAL
fIbzSbfhd5RE6trOdjx33/rHHPiZ6IRLFitS2e/GKy/+e8mg+uKTipXzfFJ9n+UG
`protect END_PROTECTED
