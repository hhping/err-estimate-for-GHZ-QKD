`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EV7vMkxqDBsSKDAq4xX57T/i38ZdR1+jjv/l1tyiXYvn/+8pk+IgwAC1koyJmQqJ
9X1C7nN6XvvUPK9Fs2fmth8JH0hGHB8jW1WLK/amlvgxSGIW/e/oCaVy5uoPM7Sn
6ozsFRoTeOr7vH6l3X1pAzKK6TYPqryDHw/ACXyN52XTbDZvpgv91a8kC4SRNins
grPUfhFBuwe+9t8fj/xyo3afM5H9/f6KkFDK2HwNqch1gih93TSvk05dz+gh0aaU
hJ1Dnd8r002CiCJabDe4O+/v2vm4f1A8kPYA5v1dRLBvBrv45lpCjIDZndsE2n2o
ZZ/5OU6eP8XjkZagAj+40dlmvzunWfIntshFwep3ItxTAzBmVFMADcNBllql0sSe
2t3+H6LobVHgEDvXHKyM1Adb1k2GtfJeKuO09nI7Ztn2RVDRYmXlVBpNujjRkPAX
aS5vO4HLkhsmAFXd7G54LZKu8z+NS8q1YKbbN2IDlsaS8bhEycku6vNPmw7s2GLs
JWoqHCNTNnnf9sJdyx8VzAUl0uWrEs+xd8hC5ajiUtNv/YOFDvgK9/U4f6fvVCrP
MNdXr8zwj4KtBZeEg8IQi9P014H/YKGJGy/DXbrYZVcRa1OcFpJ82cLGKbTk8p1p
0I5INaJoYIYoewPjRwVzOAAxMTpvOWLdEjsPFPOI9Dj98aqBqRO0cUyxce4Eggt6
jVltxK+gmIjndCfWlJyurwcSHUkKC4ST8GwXXOUMATE15FNYpMW2tdKz3PoVdkS6
GupaKTBYU/WC27EfmG4oya4MuQrrtvkNy5fnIJwAbpE=
`protect END_PROTECTED
