`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aooOOApxudXqf8B+7S3pex5rZ0/m1nbG7cNsqnbQqoSJRNZsTwPD9QQsnWdWMov
qMsNRngXfXphhjirL50V0BTZCq7D05mCoVPZX/sskG53w7J2qji76D9Lg8s7x4+m
gyNeSxd6STmh/D6odfNsIyQXvRxygdqvJAxFMxAIAqof1HIVXkbTBTxpyY8jrF5m
y2JSDcSjmqaEIUlyRZoDNfuF1sUsWqiKV1N6/wTftvJ1byucmAWtl8K+pICL6VbH
0NW70Mg00pNzMavFYXinZceG2itSHcdqHTj7LpICNamcVsRE0uSwoVu1Oe2DLcCk
3Z3bSK/qCmJ7L9i56jI8Fx0bQkn0ems5pUoskD6cCRwGxVnGtZjA02TtRpGKx+1H
6+Ct9ep7ykoHd9DO9k4oOKsqt04zfzFLcXMJuxjKgmPN6zmkL1vSpAUx+h7gKazn
ua66dzvDmZVwArNvkIYII/fXoLyeYA18fZ7WnoN8oK1bZ7qEhnNCJabDnvJWAjUv
niMP1FF/JYJ+3pYewEwLQWJPcHeUYv67FbT1Rw5QUz6qKNDB1Vr38LlOoE8MJX9W
BOC2vfBf8SBagGpGZcx9T+DbV7etGEMsXHPS9+uut/oN0ctvM2ch3qBhuNfo2smr
oEyRzzJCY96iB1YrviCbUosxy+j3BAYAjjLfutn/6OPXkRTYPJ4PfMXru1asmLgY
55y5LGL3HpsirFgM5cXqyJ/RBcPygJJgSMI5TYO27Iwaa9mcwip41lmWrcF002qm
7tSILM16H4VLlgF/BBZNqQKh0KwE3S6C/m3COtaurYqfSftrBGHmQ0YhR7W4Gg2v
v3XOPhe+FNJG4nlqO4QYyE0FkSb4TfKatmuvphT8gDmICYnFo4cC/v2VjbaWVY6L
TdDC4rPxNkSMyrHF/gK6Ssnp3W6AE/HArCFg6M9CQtpdK9lSd6p1+bnE6eHRl/Qh
P0MiatI2FTZsfQJaz8B3wJNX0pwiQLYHQoiNrMYFS8DxHrr/TAiDO6XmlQtos9So
dSj0gi9JpH6lsdSqVPuk6ZnLIxcXGv/AqW5GmAgEgRwZweGMPWop07PO/FMhfoYO
WV+DvOXD22GuXdRnrV2z9/gkna1O7TOJAdr+gOngq63dJBowk2uHuvtnumsU1r0A
/LDoQwB9TnP5lxood7cc6PhIjwTT7D/yAOSZPd2nh32DhipF6W3F2y/Xod7S/Ckm
uRhysL5QzAEikbtMH3xYr6uS9JV1k2yZlntZRu8heCAlX8P9GjdbFACnaFUs50Wl
Lb5I44gY0x9XwJXTBrSZZDS92sQ6NpDwSwbwJKviCkTgi3msDEEzeGp+Lygh3A8b
4CIonv6WuoWXVbz6UBSD0/xSDgH6+u/4UGlD7/oe6m1pGc+LW/aPyKZEcFQd7ZlD
ZLaKPsb2UafSBakw3u7MkIWUp6yMpM6laiWrL8HlwZGvfiz9Py5PmIDkqUp9vBn6
QdhBxsyvWGLBl6zxMcfwdewb59kXVt7/wmSVdx/CRCh6Ub+ysySONnmniB+QghJ0
btfZ96JpkSz9bBlUOBohP4WIV840ZYeVHPsIXRV/pM4N3hlvCG3q2NuE8ZpkSX61
ySWo/JfULemE3pPSdclVqPEC7XZjnV4ZI4h0RGPJ500GD9EHwCNENQceCo9CytmR
vkC6fzi0g3ItKMeAgHDlw0f+K+PwEa7X5zYhOjIwWKaSBWWpH6xcTSLt4rbyQJCF
mG3QVRBmDLtMNTvTQ2Bj/fgTdHz6Hdp8R8MqePIt1hqdJePECG7wNjk7+ryamDAz
cfNyaWx6KaG84kuKO+8+NVSRruWTo4NfW2i7EJ2Dwqq+v11N0vJ9g21vwnZ+/QUH
jDlIJ9/gy0um1XbNQiRoUGIYwUfbjQITW57BCzYE2R0NKqqdSt5LmfTwY3PtK/LR
WZ1iehKn20q9dP/wK/PUJ944FK+v1cAde/1VOb3SbcfSY4ZYC84TMUAWWyZLjl/j
qZV/Cpg8B/RkckgQzfTP0Xd08FOp/5kUAJehefYhWwpDUHDRpLFP8ZtkGzJNyVb8
teWzw6LJC3OzkBQ/+QyjucLI02e5eSnSI9eesLHgQCtV8ns+3nOIfJ05DV5zzL79
IaKjxznMoAIgXfCSrXc9ZD2rdxz7AhqeZut3vgudpjk8RwnSE4FRLgga3cZvXBQY
t3/8cZyPYsXtnGI792QaV23oveuCiSdsAvvPfN+YVjsksnWE7ysFRHVREsCB/3Cv
RolCeFpYpciUlbBF7lpOWhAYM++TlxONZ16zesgUj183hoZorMc9/Q3yg2rb9EFe
KyFAk8WC2S4l1UkYv2w8eqcbV5cqaIOCt24O5he46DEzVFoxGevri9v/Fl2lWGSW
hBgutQ3PbUUHPeUN5eK70Hemy3kppVnPrABVJpxDOFYOMHLsj8E9Ycac025675Pn
a4Wzu78gPOue97MIIRPQArh/OeRapKC4ngMNnjRi/S3nifuWgclWU7TPLXg6VJ3A
9LX6aJzEd7UImSwh4XaWsz1olj0UYw/meELCi2ao55ta0nqnjDdUWe3P3Cgb3tZW
w9Ugv2rKw7xB9WbWpQ5G7yUGuFq2xnA15wD4l5EVab6E5sX0C5MK2b+LIjakdIjN
0LiyYs0Dh9I/cOG8cMwtNBcDEl1prMC8xvQZshjZrApZqnvBscg5n7YgOtw2D4C9
dDcN/gN841vCHk6Cz4rw+FGp2xGLpaQpwqtFmqp2FWNKRL6DzCEymhH9T1ecXYEg
lVPlPNQbPRYn4pWKZf8oW69T8KjBsH8BJPooAX9G0cGZzSCIlVpLRJCdbHZCs323
Axm0Yt9CH144Wni8UPJBCGVA0ZdLH9UTVhifQZpQqLiWenevXNk7ZzCxDtovmqy3
rhsaIk7nFGJO1uQYJDFN/52Qdehhnc1Yg7hvwrljpwzldOk2Hb7uUF3MlhC1etpI
g+rac8CyI0OaKeRiCprlxjumohEZ6DhTFU9QtxUzeGT/G1jmand2mhb/il6ZlXmV
2JqtRvyCA7MArRd7FmFCTEVdbP2mJbsoLEbnSUdfRCqeSh9C1yWGUJaz4sN7ygDi
/8ClUjKa8JNKko7cYIF5HreeDCMD95iaCHfEYNsY5zaf/ZjD3S2uIXAtECqXS/vb
oaATgr7TivY7IrKwtUGPrfXh7Q18f3fY5BRP4QlegLMoOH002NqsbGOSr2rjp/Bk
wN41jyWtBQwsWPlK+YHdHWIaYw4c6cHw3LfRh0eI/kdB36KjEB8t+5B/id0cB1Bd
j2WeH7/ZUnO7Oy8nSj33LtUjVujuf+pqTgFSlkMvgjJNXkvVDMaWpuOlRtqB5on4
TfmfLR9sJ88bEStmBopLKFGt9xxwcNSEft5llu6Odq6aej86KzKbRb50v7FkEYjN
pxLCcfpsnUVrUbmtRKvE2bNudoQ0AL1aL8xd+OmSqbjvXnW8d3qBIQV5K2bCNPb0
8qzpIffeYIfFTVJvFChIAsjRXMToUM7j/xsegdW6fFrwyA3O1AwFyLlKiviGdKTM
tVWx1BK42jwdLwKD9FnHi9xSx8k/t8wvVvc6P5ue8xSnJn8purF8IKFMMap8V+w4
wVJ1H+njW4eBx+IGlzRBUGzOcc+m7/ppYyIquA2SSbbHR3idAhWfcUTKyqwIBzQS
RencSKhJDNXcsyb3+kb29THvhzCe1XHaX9uBjDlwmH5gEft8cWG2xn2hum8dhoPR
Mn/fq9nk1tEC5Xq98yCEw5kTr3PPkXKXA3YBbcF9/oGGcsCfr7EvY1gPfSO3M83b
N7gSVMprLcub6p1HACq/mnXOZHyungwhArOgUkAVymwNT3yYRet7naRX/uHwe7Of
b5+MFv6E/1FEbJwWa9b53WXC8ipyB8YSqRXTOrmz2DBD+cG8fEpzFxKgnIkE01rB
8UPMraNB4xnoF8w+aeo+99iI5kfoGnpVtYd6oK5s70cQj082d5/BCo9lo8RJrb51
GMIv3pnbIq3ZeUDeA3GMHlctmOoIrWBIZuWCgm+z7LvvaM99VLeQDdSF8NxfspqA
Z5zEGeFR8wwxij8ckJw5GKQiS/1EGnhMAbJitgIxMLGBK9NMUkFOA53JRVx8q1G4
L7XGSun87IdKuTGAzqDdwUCobdoqrjzQZX6pycweDCtMmfJhRokTifose7WzJ9wf
WKYTuIJxs67d36rYSKfMcYFAOwHqW9ce6af2U9eU260A6L/LmYe5xgM0WNhN7OJ+
VNqNwqHxbpkjiN1Cxdi0V9MGa6mTUwaCfE2GWmNiVfwYwfcGP92faPJL+FW3a3/1
kvyLkSHTpFP/ZUuquejG/oINOtpCs8OfVwmWPFlxvPwI3jIKm/W0IuUoXznMCqeA
A0K9YiOKqt475v5c/WPUU6WC5FlYDNPsXOrwzFlYr5jkMfzSJglsoCdz7My1PZPp
6XmRfclsWdaulkzl2ZSAAxGqlBpw+RlGd9sUF/NQ78Osex0Mstw0er3fx9VTt2Yd
Qc3qS1Iy8k4EK7n/yZxNgmo1YfiWl/g7ZiP49W+wDxJeb2WhwUa/4m87vlWyPeix
9hOe+wdw4VITawQeubJchWK3WMMpTnu1ZMUEpmofDNK7xhf/fjzIxbpcaadcTvxw
kJ+ZwEcMKDC+K/QxUeObuGTQ4bn4vOgmHPnfCsHtXq5XkhmtaiXnq5m2WP+/qhcr
ONwqHwety905WN7Njuy0Bq2y+RGDTwJIuiB/ZX6TAw85dWCO+/56BLgCI7TsJRyd
ldaDuNDrDKicLeGIy6uSO/DNmN7/9HpH8UrJk3RS6EJ3dYJDZR3sqb/UNUfRMWIT
i1CJx6qAuqGHdjv0VJHb2NwSc4MTiPn1grfYUchk1sFuSsfFJGMVucB6sZkmvAnB
8CeeXkNo4YiUr/C5z3ygaSAR16iQSCP5nVPiWphHKhL2FrzCzn/97GLEjymyQxzW
b7DQxVtf5o/4nzjVOMQInNnRAtSU7pyUTLg7XRHPe293uwz+luxf9314hV5Klf9H
Jm8HdyLuVf0rp5WfL5H+EbqjVmu+fI2WminzfdZQaERX3QfvbVO9d6D3HY+pMylg
HlFhGYdCy7gTfDsnv5/SAVTrPSSKSa42PrQYXTZ3wfV5c3x3GdOZWBBhyJ6sM6KF
28K/WrkqsmB8S/1EOaZxhMeOYjOGcsrztxWsLD0N6AQXndrHdFrv6k8fa7VsBUXM
LKHJRc0/JTrMMqi1wESWTbj1Q/F+bAh++AWDsuKbGoPoJCqPnTg3z2V5arSQhoEC
VxBSVX2IvJHik6zSCCjiCsRQmCkHpk1qgqyHG73uIQljlEB2vABk4TeaMuUD60fd
oQd2oyCUtkhXwNCAHSy5G0foiSn3JOZv7OBa3LDn6Rk5TiNAsGvStHue6cX9Nkxj
0i+pCkDUPIeiRqINsmnfX7SCGCnks5N0FMfBC5O+4AUYfy7nbNg/l3hZa2Xx2i/7
hv2LHXSa3sp0BzryoeQx3BJSvo0C9YsjMWnjNsh2DVrpOm4S4irDf3MFtGorBAc0
1AZqvN61gpmo2Rubm4pFGriJilbtUsVSbQ2IcisRilSyTbLJwY42xDfjG5L1/v3q
k7GAUyb0epx8mCB7YC5QKPMobq036aF6fKQB+o5nBt33udEBb3LgQfwMuGnt6n8J
s6ggQgd3p+zzjbxAWxqCQijYeU+127NbGelSXZ55YRSOvotIj+pq4g+dsCDtDF/q
8Og1nUl7dZLx0YwP+e3FaVBrDSNZAg4AjUT5dXHFkZaZh7wNWJXS6NxhRA6geomD
gS0b+Kl8YKfmS2SEhzoJD/ThUgTQ7TbAeH9y2edRAQoO7vWsld6du+rZxLJohKyC
OoSoKoCBDnwPRZIehUddcLVPgukGVgc0wEBPbwFNn1QJeEesCP605O7U8+VxVZjc
pT3n8xKr1OKZ+zbVyrfwdZ5kOiv5pbzoSh7+LQRABgPzsFoipA9xt85sWHQras4g
e5crAwMUNLOEbIahV6oV10vLZpdGmg3Qlhh7VVSSstvNCljXtKfL2g7At6ekvxhE
5DHMf/JGnuRjHC/3E1E+nryEATP81ByHq9mhKsdH2ESHaekglSbDsdlblZYWKuzP
bbt7am1RHSjX1syv8qIK/z9V0U75L4nv1gKg58VKzoKGnLDyZK6bPNlFYBvZ+Zkh
mNDQ6+F5kgD1I5x7HY/AtRh/q8aaiesRQ6Jvloj5hAncez+2RSJ1PBUvcRC++k9O
PpL4Rmmova9111A9I2snU/Klku0wvIohI5v7rswCSFrWGvrfrvnOkTFElaDMgqRR
bXAZVFmLF+Dh2NejBTL+OS8AYnyYMi2snWZkcvb/w5pzb0P7sE1/pGpeB/NxLcmO
RMrC0MmDQDkOy1okWvPQY9QRnZeofIWfcWI20U3SeR4hYbDwTtSLdOnM6GiznXko
FH6kJj/Vlx+Ja2I+b3n7c1c4D7uSEq9MRfsFk3iuoSHNEO2ayip4X1SOOmaSQryh
wDlhfWsE9l4UlR8EX3F4JlQnlo3DA96luMsjB3LWLuV6r8g8PZiyYMrIt4lIa/PA
+8c+r9AO1nsW4Au0O61G3GRDZ4cEb0HTOqrEvh+TGr2nPSbO8PxsIqmueZ7IGzQN
irln2icPpRaMFmUiLPt8UKl5Z/bMl5qxi1XmspOAw1cy5VdiWrrIZpzqock1YIRf
e5u8p0fuMNpmXeghPhnp46uoGV6fRHFp81kAZT8LXGTjfCb5+PGDIOdW4OV6euVO
SFxYWEb+KgP9grPoFaZyOjXNQt8IRy4RDNt/f/NnBlcGjGSTcO0djWlfvU3XqwrF
tnUiFiuyo42bi6xhibHVPm69MYKGUwUvUFAf8kp5drI=
`protect END_PROTECTED
