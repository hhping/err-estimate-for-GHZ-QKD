`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uty/Wa8wIDGUvRkhzPXXKkpt7ZFmc6uDaUN65uLGmBhvBL7awAk929c+vfbHhoOR
5bIrePV/tclLm20DEawPVtkGtTNkEN4s+B80VRAzoAuQE5dbC1uwEcX1qJN0drPV
tYfXoBd4whRTo9w3nvmgYDF58I8q3+8Pizzu/0/WfuB7Mc2f72tZNLrVCAbNiEKg
o/8tooKcp47ctjB0oM98cEXvNl11zGcAsy4b6boC7lIbr94YAyapX6vzVnGG6Wem
cj2GO2FRKGPLTbLmt6xAIPcxFZ+sJO1lGylY8kU7YJtaxge3EM1HIxPH3Yi3wwlX
M9oKWmjoGLQAGxykMhASM9F4s4+QWp5v+S0O/WGIF+atfl9mWQOszZhDtWkEcqjy
v1NVc4A2xFdvFViH9SsHPepRZk4hNAGCE138YB3+44eBHV02hhom/S58nKBUge8n
leo6+DFmy7xrAaMgywXyfHG9aGqEddU/1oZMTvstyfhFllQnIHHrZlcj4sRwkG8B
PGBhw99ngUM6mPs31OyrBryeoPywD7ednwltINc3RLWjwnVdW2dIR35sl62iEUb5
GplvlXMxtk1nZmbWotnC1ki6V+H4bYhBu315aKLQ+FyHh2JJMWff2HGQgVi/GVuE
9BbirMdwGlJ1ntxBSj6bFVq0B1e9vSS/HsYL74+6c/E=
`protect END_PROTECTED
