`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eHsTCf1iOSBnP/1Nkp3W1T3WjPRF3RpPp+x7i0EmYaDNn80UAZr6KGIPuB2kBpr9
1d7azfX4lJTjkT7ALAIoagnlojHy9pqdUhvs2vB98bQUPcPeu260XtQzbhyaFrmt
mlLSodAdrXKNZk7KqhQZ18lmO2b2FLNWkuHRcF4u0PHKlBbjKsOdPg/SOG7tJAK+
KjhYdkUMpNT7e4LxRYkiFaWaBO36gCCrc8RovfdgEuIErdFGO7XhJNx3AddXiYRS
qTl7p28U/Ypwch79obtghx/N34MyPb0o1XyvUcvV/wykVmuCrlolPOS1RsX2Ad6/
wDzNjh1+J4jmv+FR9F5ZLu2shWFJ6RLiB4nj8Whe3ir19Dio7IcrkPJ09RsoNCvI
rjXNwFW3+u/gf5rkYRBH4w5zxqumSsU+3Frnv/dwgc6gAofa+rQBbCbZMnYOauWs
z1cQ4j+dINXhdXuCNmfA9gSUqLrWxNDvqyoJEWqiNczK9RO8qmOEUxFxteC+jS3P
UU1ZWzTJxxffTvWIEk3o8tR8tPjyv7Z1i96K9AufKmLSoYCpl2/L8CObwwgqinvQ
BGJs13PZewkyo7EUw78+vZrQihXUR3PriF1p3XXpfJ9pwVi95hxoBvSnYnFO9vcz
dhnbP0DlCidKIVUcS6EYTmGb5kWmGfh74LEdO4NBXmcHA5bIs3R1UJSMHubu8eQU
g71cFp5hbMAty+8fl2ziGskms9+/bl6n44tKor+pzDg9tHqUm2GKq50CfJH+UVRk
W71E2qE5XYebJAYnNgDuKA==
`protect END_PROTECTED
