`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YyBcrPxeHVQ8SZE7M/ZYJBwMEvI8r5suWRx5SwzYzfkl3P3EP19UZwAujdkq2w27
wAYc87mnnjhJts7egivEJcueL6tMh5dOvtJ3dDWtCTPy7k7UXBzqY92/2gA6YDF4
fiRvM8i5+Fbx/MP9HhjFAv8ZC1qHpThRdpw7j8+oXmHtgIk+Vke+5EWB+9ar5+z2
dh7Iy8rl0lTyDeIWt8dMOeREms3+smxcYQdTMEzWLlildZLHU69RA+MikQkqKiP4
RWU4ogllbDJA8bzTDSyRqkFLOd4cm8wBvOxe9CRhWUtslxrPLvhehNFoxOeqlMCI
v/V9o7mglWsw+Osh6zI/7bk7RHg2bz00oGQzu5un9Eo7rQGY9W14y9AffOELjIdc
AlDKZXjK33lreuejuws/ZVOV4TUPAe808tJsDX8M6Tuz3K0aLGJCtw0QfATG58mU
DrgZx7gH4X/5RqqJN5ld/Do928vY9eQsDqz6gzUgeTy+IcYahKXONfLxckuK+Nnh
Xrvv6P4nf3yV8iducw/Hz1Tcc8z70CWr4NE5pWiovR9CR2N2Tsbm+Y88DozQKOsd
QC7jnH7PkDwdiHWxXIWe9I7Rpkg0me5zCmDFrYo2IRHuHenbr6uoOiBjAc2neyrz
`protect END_PROTECTED
