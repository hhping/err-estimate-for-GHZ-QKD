`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n70ayD8Tc+b+d6yYxJtiaGYX+JMFKdQyjN6T8TQAX3dwo7MM8pofurUR+ITzMf9N
2snHXdbV9oygvzBlx+rD4hOYqtaGoI6sfdUAlZ0Y0bYFnjiSH0CleXuHrbV62X96
4Fr2EMTBAqtBiOgSAXizm8vu5A87vYTH21gnU49jffS2RNoS0KiSUOo70HtR+Vf0
KhvMTKnYcsv2zo8ik7wkrN8lUcIZCMElrMnUUPu2Yqd4y77vcehJmE8g6QSvCzga
NHrkhHIUINgE1RjH+I/x4C8vzg8UCASm4vab8AgIl7CKOnZ3CHS6nvF1BQ42AaLi
KkEnqody4k1qz+wcslz9HZHkHk2EeXZ8sau7KV/K78Py3Y4L9joDsTf9fnV2v58Y
WPEhst5hZO8mIotRUb31ptr0C7gvZsDlwzDd4mIrIEyM8BJB4LzaNdVKZ5QGP2uL
PwoIVbIwsY1D4UCBSNcn1vrZUxOv1ToLhs/+ZyiGTQiT7jzZ2LKzBQlaI3UXvWyp
G51H3FXrv1tpxn1HeGq8kgisXeAyg78TJtq55jMB+/lKFjIskl2OionzPmYUi63q
x9JdKq7t4QXASvtWpmQ9ns6RY1Tcj5TL5ZuDkaf7IDcOPGV2hEJitl9mOeW5ueOV
M5Lx+7QTHifPXgGSwgr67ifR2JTqLgiIcGRoH3UBoYZFALD7yup1F7mfGdC0aba0
SNPjONsam+tLM8mZ1CAgnT/Nyb5L1L/zractDE5d5fdWvfL22TOf9OZ/XW1PSZtF
KhzbQHpjjf5O0V59W2DUUJuhGRPDmOf5XHo2VZk/t0RcKhBjsxPPeeSubal+X33W
wDM8UWFlN060f8nupbRBW9H8cCKTnyrRESO/FMy0gXW7+y0DsCLelGonlF6n5lq2
/tqZmWI0hgi1OQyHlPU1i7hr9ytpaBikkRQ4o0fX3LDBp3iLbBNPwq0xJ7aWqRfz
jJPxYn2Z/B2SWYApkIFg6qdhbZhjS/ThjGVIaCt/tur/dcmGiBYeZfd6AM9gi+jP
mwJPIYlePs0r+gri/syXdMD842YfBw8VaTzKLM/doeFpr7UN7Y5EbxmyC6/sV0jJ
4k4DJI6jFc6raMznZ6CVl/zDdMOwek6Vjs7MERFV11Rb+G6rEaV4ES0zYJq961Tq
rr+UVZ11AZFKBJUk4IGteyIuCCnW5nYKbwbuGr9s9/McuKFnsOh95t7thI1+Nq+B
kyNTRdO8SRA1IB0j9bc7Pw20/YkPt13zHHnANFlHRsWglanRQnNfLqJGE5Pv2nRO
heJws9WoKL5KlHECP0iFUXyAqLVXj1gzIJ1Jnmbk3VpEHofiEuOdLCm5/bu3oaW0
`protect END_PROTECTED
