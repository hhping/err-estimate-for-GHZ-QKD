`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ja9vOTiY85g+lwblE4RohhZh33q+5mh66bfenBhhNXu53EuqdHjpdbvi/SQamWjo
mGTbI8lT4FJ2tJDthPknh8qJfJO4GU4QofNncQ5HBLMpsfzhYjYfJtZESQC/omjW
TGZQF7LNaEbyz2G4RGg+TrMPlFvmu6cAUPgIQR8LUkMo+mUDtHnslb1caUZ6QF/d
md0dSUdbQqq9J0iGl2VBbB038yw69Ao16ZbxyphY7sTDbOgOhvc380NdszthtU23
KnTXodUhHM5LVsnClr8Mkmru3Cyamle5Ahf7cnFqwBvJEhSVBr/SZR+ErYD7Tkm4
FMMaMDo2xEPspvZYwq8pQ7E+VE57Ph5U/Lfj2gYkCSoTbTkeFaPn/Hf0YIuoepFO
7LUL3F0Bgq8Okpcgta+loEr0rxXinbtkLOCN8QodSuXwoz5gBuWsi15poSjsbtJU
5lEZM8Zq7HnvzVdLClsQjms4HxQOoOyIwHcsRdreSu44AD9rIi1lrAHS2H7RDGZf
UKxTdPwMQcfMI/D2g3QT/JgvFRMrgqJR1zIfEad97xdagjpStRHVC5I2UY/xWbLo
qwBi4JR8mr7VOtMeCBTOP6tXyC+Y/4LDm8iVhrNh7oG1nxdcH7qZG5at4NtZI0zh
yUYbMo6IIshYWJW+8l1FEZ1cV0129FViSzWJoTRLPpnIfMwkq33eiLB6JB7us4Pi
9AIKCyX8fgYr6a9KZfzYIxVOJeG4D+pWf8cDiv5TKM6aqDY1DxS93z/4z1Qgt76Y
IptpZaUjQvSfMCtqKTafwuwKCDJ8TW5CnhzQf+h3d2c=
`protect END_PROTECTED
