`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j05PZj45Ck+097Ss1DPdnZvSr/Vb2ZndijpDWsg9X5yIYAovO7n0XSwzr9DuXmZH
CrKkD1QH4pWNfYDbMyRB4JGPxwjDSZiBvkD8/mEUn0tUObU7Rq06pwx14sclvvl+
3T1jQsdLYsKzaw1Npm3id9buiADNfOilCt0f5DBW4mqkGWDz/eFRS9k8p5ItK6QT
CDg/HwraycwoDvonFBNMoiH1ajU7AkIE6CLFRupdJhMbizgoFhXcajMcOfxoHWH9
tqCswNbKVAszUiVr7oAPfZcEsabiFYOmT/ElZcXTVDFBYcAt5YEAr9zS9cQU5zJN
3dK3k5Ri/eoK5haE94FVxtal2svw663Dwq92XB7kVmSXOqInpMXcZltIwZATHoFT
z+zxoQIUci8+FT8cF5wqr4enq53sFk8S9Q+0PqDlcQpXde6yOf5ZJxkPUj86xAS/
Cqpfjh48JRc45+ampICIAeEMbl7hF5LdQ2qRXN/GMMBpG2ThDpJYd+iay+4KJh47
x67RdHg1EQ17kgRcaxIRoTQoVsk1gc6ENpm89X6e7hVTgNszvcOicb09kwmIagj4
pR/CRQPpNvKgSMutpeM/OKxq/ico3MknBdNF42oIXt+il4B6wJq2/SpXBAjdOHY9
9vlCYt3Jb0K6nHOO8jzFoArj8gGM8aAHCer2hrDEbqs0ZPApGt+2fetVvhfvvJUS
D2FmADf56uf8ybN9gun4xs3uz9yTNNl+bGRssL/vUpENzw3r+qwjtAiZIjpGKe4P
jygCAXGD/q9BwG4OESnxE1COd/a8pIGyjRkZcjQXuN8=
`protect END_PROTECTED
