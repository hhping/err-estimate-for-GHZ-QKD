`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QoB4zb5zgxu76CL+RFGdXrmiG/3zNKHiIdlxR2zptLfkpbV10RNS2ftXV0/h9Wxs
hiRygVuOSiHguvzzRGjmTEN+YRlgE7bqY6LRpNWe8wWywez2R02nTB/TNXNRNgfs
G1S7V4ET5k2gyB1ZAJsVb5y+S4a9kRqdxquTmK2HVfyFEXnpopyFxI596OLTdPAN
AmYJQjLMEDUZiI+viM0t+4OWP+yuHYYuOoNTawZWmUyou5hl6yJSLRY6brfkyzsq
k5SLqxiLYj5fHshQRRTagpiJEFgITLWLL6lzIKes1AiV00OLS1nLU0k0WT0vrO4e
DF9Wyu75esismBRxRA04nUFjblEArVuL8o8sBlTNtyGK+JG1FqvJMsCDFU44hOll
GOQ+5XsXvrrx8m+JUpPc1Oa+PfYY8c/JwhQWmyyRX6S4MdOgD73MddqLtOWcainy
WcjE6qkVaMabY4qZKRLpaLbgwvn5bQG9fDszvRTEom1uKUYo4dyfOROCzWnlvwJ0
ZIZmlsb2C5cJe8fE1PzuNwf+haLjM7jHmf85H/rNDiWtTLMP6MvJrhClvfE73kK5
NLzs6ry71cTWxrDT/A6XNe7PG/Hs68a/qmFDCDedB2Rf6mLFElBcUD4doF9X05VP
C+J9s4Z24HUb4eveHrzwto+bqoekkuw1GR3mVDQOrovmF6EU4l0XUn7wYnl0Z6St
3VO8HN+wV7V30JuL87ApHLfLmFF6Nb9jJK1CLb6IsaGYswMcYsKldCcUFaDw+yOp
TlKwp3zyzF+WDaSmqfzjFMkltWSWbCwSyfnHs+PTldtsczfSNKTMkfeQhB3XSiVb
oqB08/UmsK23WfPosPAR7JmFrf2jETK6AoWtq7aEYNztdsJKcx0Mz7OfEX0q9rnL
tOBvFES68G7uucjy9PCELDLeSX/cp28dUT4t6xKdvN/wpMlYKCbhTwgz657KOV1m
NuUz/Fjq9IZpFQTjFuGJ+eRp9satCqyTn08uxIneenWmAujT3MPo8dqIhAwnFhgY
XAY+rOTVa7qHMB5FuulGCQT70a0Qcj2s3oOWMmlBKtwHFFq4uc/hoywJ7pNHOTsv
/rT+/tsY+46lgJGpD1ISUnhoG0E6mqmqqIQoUf89VqVLz3lz0HvUV7hl2lfcjBgg
R0MSoNTAAqcBTqNM+PbIxDRMsaXcrIzlU2ZulSWK+1avk/yz7eLwHiUS3H4Cbk7D
gnH6VCTOQ7c2r4kig4SGCDiFrRwwAtf6NYhbZFjo93S/0/M3JOnbK/QZplxjq3cW
dvWWNLIn7klObfeIfK5+x8liMMB/V/2cRpdmeGBESQz2zVSC3PBdCGzOZzNrWyDq
E1NBy3F9mfbo6Cao9fV/+bTY7WcQNUD1+5IuXq7edC1PJtYsRkcOo/jT/5B24+xv
TSIi9WgxQjfxCN1OAc4BiQtkWnHI5KMU2WqZfF9PNRw3hG/5idN64mAL2h+Bls1X
lJZ/UG3eZ+3MtKD9ryt5pCzGCBPoBSSHKFZM0fUmC2Yy3ojyLztHBqdJN0sNcHi3
TSDSHSYn88zZW9Jx62WlaTNf2Zp5eR+uXrIbAASZ0fc30VqpWim09l4uZKhb5I0V
/5xFKH5lssDePme4fiFpy1N59H2T6UXxRjhvGvOU3TGfKl3p3Xn5/fdheTohAZ5A
3ONB9mwfUvUcbZBIsOSc/k/p7m5k2wLYk7ExEXUSEUlq2Q0e9GF+weLSZCMx+cx5
gpXxcYyT9mDmAt+D/70ip1yg8YL+GtnuSOg4Nd5M0sNUwxGwMlJRF4EvL8W/lECj
cspsFIVw4G8yhUZ98VZFOZ3+12yDDjCmN5ooLaZTnmp/2V6z+yFO7LmcgasBMjAg
/lGSISb4QGNyZqv08lYf6osS8kIOn/bQJgsWWMfbPHKqq5QelMgzrziDeUlIEgEc
fVvAF7MoXRRmWdGOHcxfXD6IJxvCsazqviuwGMB2h/uckulAsKcrTGxEITHo6UiB
RpmRjnHauEO3tlx/4O2EGwYA6ujAIUYPyyfovWUB1Th0T3KTgAHUnk2TC32SCJ8K
uKlq1l/hwBM67dfzoZ4hQyr1ILbHsx95lfFL9o4hxS1ncvZbMVaOdUCjbSxcxxls
Vwj8dTDg1Ng3fe1e3DFFUEuIinANT1hD6A3W6yb7fB3Jni/PpiIx1vCbA+T529D+
Uu7TMlvjklsMsKT6ATHUUi6P8OIKzlYthwbTtCgyI2AzCLuPbtkS2m3nD1E65brG
fq52QDe0/oQKy44rJroNpU2570hEDCBL+RamSaHfPrRsdo+dW+OylwZktmcPaMA8
1oJsSFxi3XwnAYBCflqXrWsN7Li5IJwSzKWyHAz7dZ9rcfPUxCjqCLAWjAzr+WYM
N0U3/FDPUZFqqdnIWXPhcQ==
`protect END_PROTECTED
