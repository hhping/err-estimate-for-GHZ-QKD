`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3obruMgQLU74dudFFQc4WBQy1HjLt4rQ9SO2wXOJSrJDzg6bwvYmeh1XnJzMxyN9
7n9a8J8cBGjqTPmXCa3uUyliwQZttMaSvbmzJtKKBZ6sf1rGlQ3qkgw7L5C+cJG5
Gsqw7YLZTAPPSz0d7ZROxLP9b1E48KP3OIweYo3m6nb1ma+hOO3vKAUgLH1OYC2M
4pDSFQbYxgNMfSllm4/68TKcBLmeWwA/ObwXHj+FSHUFC8BItuYynDAVJUBEB1+c
FBdAOM5U99nJpySFh1KEAoGIfmoyVtW2Vl/hB6/MWIda4trUaz926LBN2pBBis4+
p7cyu2KRMe8BSqeJ9CiKNCo0KFxEnPUEYKsBiIUOpI8zINdKdn1cUj006iWU1z2V
nOPBxiEjN/J2WP5c1hmPQ2s1cgQDhfBpwxKvQdRubyZ52HoPVSaA4CJadudf5cY2
5mW3421O1qB2dTXdDAIsIPu+Ao4AfsBDB+4sDs9fSQsbEuY3B8eh4z2j+Ui7aKTO
fdOdptehrCFmx9sKa5KhB3O5TpZG1ARQc0MRLH6Qp5NyMImtqEYThBzSM3rEffz0
jtxMpjV4jiVMzk7YZmrfj+fgbZFGo0O9ILf7updTu8hqpcrKdpBFrZbAP7PxcZE3
wIZxv5VKtSy9uORvegFxEZFIaYxkEYUVgFHDwRZwjJzskVY7qUTLA3ZrvugLxfCq
oQ6XVZcJRW5iSwIt9SNRX/H3R1UiRTpEE0rphMPPl+Kqtq6zKyc8FjlMDOS4lVpe
HhxZU5Ebn84dTcIU/wIsxRh8/pTC1YFSS+AHXWSKLFjJy2hAJbMw+7OIFwVkLGnE
RB7HzGHkjaIP2T74vqphRJWryPAA4atyknnRZNjg/t2/NMCMtTwSc1wBI/MXR9Df
AkgUlHxLlW/zx3oDBqTUEQ/d31pVFWlB1np0gVU3ZNt7p88/4hF4P9Dk8sqSk40K
qd64RZz+yDW6XSYLb+dxKzzfuI+6TuhCIfDS0xZVE2Rhwk+C13wAr7Qv5MhgZAPH
f8I0cjOxlGjfuSBLs67M8/CLakeAhrDEvkQ9Uh6Bv7FX69wg1KvyU9idfzDSDnIM
sdBR/OoBhUfrVydEiv1Qcyr4vtFrTqLz0xVAArDMnuk=
`protect END_PROTECTED
