`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ph+GGAq9a1OKJ+PGNB3CnP96WfKoicU40TNjDUAzBcazz91m6G9nczSESNGbCoum
+nPgukxG6/mmr9scF4NVbYOH4pNP0FtPTEnOu+FaIgqqzzcW972YkDJZU0yjVuEc
zrGmAnAXry3aJ/TeKF4WuT61EsK/r7oZ6UgwlBpq4KSV3ns5b8zzJbOlJxhbXvDH
lDfGRzRAjkSM2rpcU2RLuvgYJpKmRWj6AhUg/B6vr8LBpJAD7RBgj/dvLDo5Kjq5
rjUCRnvVgCfL/NRdWxg2G49RdfQ42yCplAXmUbusbVcT5ZfgxevQD/ZnhmxtMQgc
aBq2HOZRB9pQwlsDCB5iAYQAPOnOf2NaZwx1AlijIagTQNFcp4+cjlbaNVv6bZE6
n2z9LOAvNcXHS2rdy8eXhLBRUK8z3PBCYNEraHGmOIPgSATgmZ6Jd1qvvdxY2BtI
+kZuOyUcVn4QDVOX5yZzgy3jTouORQe6KJszgtnm8Frf9LGNr0p8SQHRPiJlelCH
o+F+WGFgbG5KySqWx8/WFg6ymQZgr+bnaWNpzgauoxtYsRQxJ9ZcNV0+lWhQ22Sk
S4muyCNTy1H9eW8BLhT9IR6srr101EfeOx4Og/AAXcd3Ss0UzKgsgg9/ZopFsSoP
YNo/AoexvzheOGgGV3oqn/asnaFdA1GvX33qJdjIgchgE3pCBvnSznxGjxc6sm4K
0oGARpwvUj0zL2XVtS3awOD5gs23MQzpmXEpWlgT/xpjWrfMt6TH1KGXW93WNS7f
7g1PQkf4MlDBrsZCiUlaDQ==
`protect END_PROTECTED
