`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOmLLDqzFw94VGlDEQ/7QuiclwlgjZIXOe2BfTpLIqOsZBQIuKZHwMrVkXVHCKCG
obiAuJ0iaJWYOYN+Oti0mKiAHqPYPzjDJ22/Cgk2c3FW1Dmik2/zgMg5mFbcJMDv
pqBEqpUbWqi4Gn9UVb4FzvHdFaBheIMIlTVdpwfsKHW0egvsehEhqoCeDDpA41o9
74ylal50/G/Lnzya1kiLUEMxyqcGY/GQW8o/QBADS7+8uMzZOvBWiQYjDjyetioD
rJAyIbrOLF2JRd3o4ttctOOeqZPhX0Pj6cM4VQlK1kT5XfMe5gTkbOYLSf8FP27h
GcxKzrtq5DzUt0y6jh2oUWRnRhlb8Rih2hXN+2P4WSTu40q8AzSp0idlyA2DxU+k
QHlEL7BTapAzvFvk6WeP6YSPKKc/mSXc1fk3pr+o/GAve5xWwBSNn0vyqr/zHsji
L94FzfO4d76Np7T4tIQaOsXqc4OnD9jIIUeifdVrPXE70v1P5MCvZEfuRP6kk81z
L/rcPf8S1OAjb5fE/Y0rczrud7JFYz21Stt8kfaqm1WQ93WWv5n77Sd33dILWbA3
8k6RIVhIgdJpQpb+nM7IFu45j5SltNOKl/YMoW5K4mQ7uE/0XxRxKdcbru7+WEpv
E5vU23vGuemSVTglK01CKCTbr54Gf5hseHV9c4jQJi7FVykjMTVvceY+bTPoqkoD
RBygHnpfUm1Pjr5COI6twfVsDVRX9Io/ztFGTBXQfZartb+ZUujvl3tqzMxNq5RY
fFXR6fNajPwf1QlzmySBCVsqwjJMV4kq9tyXh/uq6grE2fozy66VwdDI3vdVh2N0
5pV+ZsKn1nAhd+B29giCZS4CRsdW3Vaq1PKi9Atd+uhHv+vgVHAKFoJ8F2wWSI9h
EIDztxLBkHN8RWVWF5IlElr+7218xymreaWQ8V8u70wX/RSUe0BFBqP0VB0k1gVB
OAL5bfITU8OSOpHL2zWIbBwFbwXSIcDLw/hXatfGlRKLjBP1g+Dr8y4ZNACPXWho
9MVlwmp8VtyWHhrZqOeuN73xTu3B8lSbzB8RLVGS71BIl9fI1xjJ3jcC5xjLFbc2
SzZ2KRhU7yeyQawmhG/y4pelHh/2N/tGWoyHps+LkO8sX4vDnfZM8MMpRBh3f1KR
wWkkGTVKiS0EE/3MxC4bzGAoNtqM0SMMSDGWsLDCPNlQ62cUr2azEUBo+1dJBwYn
cg+2lNaAllLZ13FZYgjMpztvyeVhTjBAS73z/kZ3qm8sEHwOiKnmky1QXmZu23kj
Co28gWTobv6IlEtUz5SNDhki1ykbx/8GAF+Fk6ft9IGb56jJ8ZI9MvzmtcoGI/Kt
210JaFYnuv+MIbs/tUG2+7ICAtJhOObGrkNj2WpVjclw6H2MquznwNx+gDcRZixQ
gCtpOZAsMLyKKYYCp1lV7QeYFnmZBlWUGIAUssgpuht62ja3dVx1PTJChvdf7kVy
sw1jUM60813tIVpaN5z+KRpHdEPFZXoaglsCuPdhchfq4v3yt9SCdyxHZu/2V6XW
I04/zznCarnQxUklJp5vikHVlLCj6Yi3EyQtXCB3wycKd8z07jd+eIwr+DGy2Z9x
NJ/LF8zqseS25yyfFTBLY7SqsZ6SFOsxxCkZjD8oCUiTSsAkEqJah6QCAcnLuRDb
MrWORReESrQdf+OOPsKKAEUo0rZUFaxNYkgLgNP1AVMsIT4Vy6tcE0l5ydiygjgb
YEoLqmAZwhT1qYtTfCLM0PA9bkBorzaKB64+G/QP1O+jb6jIP6IXKdSLCWIZOzWK
iw7oZsziCWhjBlgBXkFagcugX3fEy/tUcOskXZKWd+BtRZS/oYa+/qbVGuF/FHex
8LpO7WdpARTx/9ICd7VcvpE+HmV+69CJ+yyTbPtGAxoSFroqxzOCrgO9JHP7PVcA
YxpbNhewRo7eDsibxftMsvRm3iMCAlLXVzDnsr+kYmqZYDNrw5L7YwFaL6X3lBzS
cjvStyLXEbBCxCb4Bu6xzqkb+lBh4ZgEpP4bE+2Nz/CPI6ClzZUv7mdYLIhyznXd
yMuAoTy6UCEWiZNNpFftsGp9yUUeOtY/rzTFi5PIza4wf7d0MHjXyT0u3t4bUBW6
JS9CSPolnjAV+PdX2agZ+MZWmgwTyC2Q7m70BuHLnpJryR1+sLpSfeiCu2iADeIm
5nWe2mWOegcl6CTaexyCDwhlAQMQV3k0wNheUJqoriV3ia4aAEW7kgaKbqbK1ocO
uIkpS9tvQgklwBB8O6Z1V75MU40WpyC3qEX8hdGQD6dZl3XsgtT/5oUfzJ2fsg9G
ZnZ0HyPK7uooZ5CrWQHgfp+cFC4FN58xLGatQqSa5Tvw6sSG0lBfGV2Hdm4ruYGu
ePHS6WRIkO0/9dUMyDvOyQIYjqgcS0wQIRcDwsF4UqxbzQEg6R5DSVh9NHcHHuXm
q0IG+mrxUMu5xVptaOY20FO0suOpudsLGy2mlm7Nxpcz3wUXE2UaCnKuL70HIrnw
fSWC+kZGwwbIKMCEB7i2UQ==
`protect END_PROTECTED
