`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGO1fbZNOUxjI03GeZMCfwJeLVnUi8kNpJlZVw8DiM218MUyMc0BxQ5bpoU5onV1
Vhj0xD3VJmpjGCMpqE67c1wj2Ppk1v3hKejn9vzdu/nWEjcBTAi36h0XUVNwDsim
jsCw9duqI7nDXUbayAU7l4JycEwJ5yzU5gzFJdDY/Wo1GEE85qiqjbWfICmqyCWy
QUHCb6fkTIxfs6SvskMwq35hAsd8k9gAHwz57Ap+4Vl9OfNT54EwkdNukiUGQ4eq
IGLDbSHwwgcMxsvyM6j3lxnsVKbOttTGdeqMgB/2Dv9stUY+YAPGPM/KszRrxbIC
Ybju6KeE4l18w5ETUxcXjoAqXbhZM0jbmqE87HMH8Epvmamvk8EOzHGtcH9wGBWC
UQgfZAoFpy0U4HAmiY5S7sB0U+duvP7QQZvWR0N2zr4LWEB4lECun5BFkMCH8v0m
mu9dDAXeWGM9u5I3YxAMi0SbFWhrDzKtv1G1cWwTnxL6Ava8vjEPPQco+F8HYnTw
13EvmFTRClFaO85gibBRNi4unUq89J8SkwyseFVFBApKVqBmjVop4pGAzYJg5h8Y
PV/92NIhnAuXDmRUILfxQRLa+sH+7kckY5mASKnP8R64gyxYNa1jD1TpzXt8GGgJ
RQ/iBlmA455GRAwbqAFCwOG5IIuHpkJSunLQ3LIaRAni+SDivUyIIGCcmvs1qR/I
TtV2QW3FgQtGJjIVDjwCnkpfrp8GGdHGCGpdRO+NocuVW3nNcnYpSEoXdwzQLUV4
4+tAx14h357qmDSIkbzWz/f7Jaxc8Q8JWR+Cal7zEy/gfKETusr857ZEqO9kue0o
rJDkHnjXyJUy+FvOv154SXy89F+Pe1IiCt7uuQgcOPmA4GchH32bsY8SZKh0pZpH
FP5Rg2Zpl/HxTYQtbn5pSv5yIv9iLZDDop6EgBv74KVzwKjEen9usK3pBwJ/LT4H
eHKCxXukc1bb9m5+JOmpFE5uDvcKgaR7WmcQRMolyaKkb1e4ewU1QrnzNaZn1Zqp
`protect END_PROTECTED
