`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gLWeaqkXCF9NaZOjPoqXlYbdTBxYo4+7aWojK5IRI5/uWEOTvhcM9FPdscLdmq+h
8ahJUXxzfy24OHwa3gjxqPAzySzm+8UaQThkZOxAmbEdbpe+oSoRCsTeHg/9FTFr
EqPOPZIHQd/r9cyOFK+AAjVhOtdBEgDQFpBLegs0dp4jykEj16rt9YNy5XRBQWlM
xYR6jvkIMQvpdQYzx7ucDkLX9eNsDZj/oF6mmKcg/vwt0SVt7pqukbKo+6YqykSB
ubp7+kloynIZ7AoIBDoWIiZl6aGpnGJEkp3smXtjsvPVZGFD4+KQPXmvXtaaxO4k
2UOCYRm3N7fEJgZ8cuKbQRH5H7YA+JtORNXkXw91zB12OwBDT2FtIzFmSAA5APkE
nl04FVdeQT3SYAAHDBXL/U5/A0AFXSSNNT0TmdpW7F3XBtWqO7zjI4PXfFYOXBOa
hKuCxOwKDUJmrJpfEC7ddI3Waz/+QYpuqKC8I39W89CIHlBnCYI8tkH08QwutzF2
KbCIVyWTCZFi5NCBuerqK6CbDSDPufqcWPA8f6+Ge44ip9vrX4LO9r3o4mVIwCem
X7OaH3pTE98/6UOZWEpaM9uWHpq5asFa2mRs5YfFk6VVhOSDswnZmhgt4PJck35g
e5ewMO6h27VpctUWvEPdtdu5esH7/zTvXgTbKfuLOgFIrmyhbJX1ZTAF3BWtYhNc
1I+oy7hQOx9xAApd3riB4X96QLA591bwtdrLGNT5czYf9WM3EEjO4cxiEjy9/4ZM
EHcQS9eELLRnqg4NMXwt0S81VfCyLWQT1xzG9hO/+mgnjNufxCgB/wilUkljfmy7
91hkfgiPg7my0IRkVA5dTDrIIJJ0+RICHV0Uao6ATk+OL2z7gfJfhbH6ykYwHtKc
doWCm7ufMvIbh1tmE/TR1233G5WXcwD8rbgYMUcK7bS2eNQEDW0Vli4KFsTQ6xSF
El+119TZ5YKGIMX1B+Z/3owHBwbR90teMOv8CRN74bX+39gXTJaqB2KLN/lAkhhG
dTIyKoOCeWLAEY2YGYxun8EJsqq6zSRDytxamcTY9CKUCUUJle41VZ/70gFQVTbz
UQVA8MMen93nVatT0kYi9I4JQ4FnEXYspQ94v2sbARRx9tmF1lpNaN7zM6sIlXj5
rQzr1MH5FZyf+2142H930bWtAZ9YZ4iPMejCuVqbC/ZyM5ADiETu2+m4GbTAaiOB
9bHzpAnFQnAULyhjFBK4/BWDE5kDMwwX7MlXdX2dlhebTJvvUUUa48CfUD/a3LDC
0qcUt5WANwHsWwOGwtJfubSHEoM86Iqu9cKMA1oTgEpFeahBlYbkqotOEWv+GiiW
w21Fs3ntGIAKZgA3/XbXR+WVIh6sfDz91YD5s9Wh9sUTohdiO0OGacy+iNkhF2Cv
DxTvklkj/hlPL9TQD1LGK1SZrIkChUUkWm/QBvJ12b1cPrr/jFq4eROknSF7w7OK
G43vFfJ4fMgPXhrk75K+U+rhHZWfnxlrNtbRy8++wNIbRjL/KtRe+pyQuohYX+ot
TvP+MDfY36arDV5FDvPijY/uv+8ZYjLQ0Cy9tSM0BzHVkydi/6QdU3C94OzElILK
3H8LnMX2YzK+4OrKE7ByXAg883IDe2ShRfOz5o5Yc2imzLEZwclVCIGTzDOSXuS7
u5nq3Kuvbgedla1mI2/QeE7HZNmi5bquo2OrVoucomNhIMliu6MX5TUC8rjMnfvb
lbB6wj3y7YJxpMTOQbkOv9yrB4nCNrFOf3CqoV3aXiimN8fJ5eXcjeYOjqUaYCBv
Im054xDqTUizDvrcfJaVSEgoCT2TA6bq0qef9NJtXywiLtat72WbVaKr41FTdJlb
c6ACZtW+zW5R6OiMmaIXgdQBArC1CrVqrxIwpYq4M9PaZKN1BYZVc5Tvicyc1aco
g0fMQ4KpYsIXVwg4rL6Fdiw+rLBbwZUofrnGCstOLMBFJKhxF96fMT3qKgnbUw/S
xaPSGhO1rOaydh9c1hS+uSrkDs21usNCZxwMmFlaLou3+5q8ZYv5Pkr6Qbnj0Jqy
H/E3+OXQqS7UYC1YDAgvNtNA4qsNipBpyaTjqIrOlNupJYATVixtL3aub1uaqMtJ
muksvV1xqg1M32lJEZ09RiPVNiSTzi0IQl4vRTUqNx/eUCnLXWHm0ZsNLcehBVXF
WAcjSsCtRhHNNssCJrhSrWHYzU26fTO3UF9fPQhkXpgNi7M//6QMLpMTu1yFb13P
aLHUPcKklsi69rIXNO4d7F8HJsT+dHRnBz9a/z6o4VwRu+uXz/mks3jblD/UIrcP
4PMHwqmwVCIirQW/G85TZF7acEb7rtEj2GFoNP7vlt99V35CkSyl68NC+DZLdzfe
MTEevJi9SzmIrhX9536CdeZDzB+7/Szwdzo1o0gnC9wE8qlesyU3C+DrAx7wLHFm
Yh9Ote6007duUETE2TVDwFm3RpWMLQcrr3qRHGQxh8XDBUeuFePGdiFFdxxxvEKl
6i78LV1CZ2Wm9hcb0IFEZNg+fR3TM6hRb9p8vpLLICdpTCsYU7E/nauXKG5KZBo2
G2OqFZ9ObvHBCwmDDHlS6wyiUf9sWJL0xTxDfKLwnT6C8EbTWt5iuCSIwpXYXY2T
73UOzNKPbTR+JSh5TBSP0Eu0oX3jI+U8FHep/sZYLlL15IWvtRzsZ4G3oFCOr5ed
joU8CgCIDB3Uu4s03KV/IVuigIOjWUCbUVDXGspq/TlcT/cKongY7UJGgeP18F0E
yC1Wa2in5oHX2mnvk2NI1Y3KC0trsJP+m3UYmnprwDnKTxaHv8E02mAyj//RLcAQ
WUOmrGqUh+7pDRILL1lgCW14f72JEbbH009qiMPWw2hwbe7Sy47EDOZ1yq1aw31K
WpgbEXB+dYmmrIrzaXlsYHtd9VlTVinnt43s+E7ctPX8DgpAUwoNHxe1iOWB2/Od
dNkkcVN8FRl96EVy1AMpilBvAIDbjYUL7NhTTJy/CPJcNy3v6nSJZ95XsxyZWN5D
4HFzbCYnRC3q03Fo0vQh7aYVSwSaSh/BDBEDyH2lGCOh3eIa7ktudKm7LjZd3rfb
RvEsR5pcgqO91q9xD9mXyxxj4J+PvkylX9UihdVoZV9fMu3HNGKFVdOdf/Xc85fm
i+VS2EKobUf+fd1hZAyIJNkh5Q1bvmvkIkbZi/r5cSOjzyGzNE7xLmiMtxOSlps9
i5jb1riPNM4AVrAEwyD6XSjmDnTLbR6xQ+770y0HXrFyuSXrwCC1lO/Dfr6BYs6q
Dq/uF9IIhJ9HA2jbkelYZojoNzzOWEqoIHwaq7IJ8ynrXr9cMZZEWcr1SgBRIDOJ
7HJwUKwz0L76TQa+HrJf5MkbnNSDvaEPqq+NFlch2C651MzVSKSsVBc9w60U3HQx
eH7OPJm5diD8DjcJKfRO0MgR7ya8NAfoM6o98z/sdcSP59HtrUcspsvg6Ikv8iA8
wRUC5d1D0Vn4NBFCr+LU7j2zCU+A1Q97SqtL2HZC1jfcOJw+YhKEUoFTsv3KsLAb
R2aDqQFOiqwmV19hzsByMOtT6VFMsfYwYFT9dXQqgLXfop3g8pYTcVGMXMo0+3Gr
v++6yPyFu343mSqf4ay0LOWFnsIw1MOU/qFkZe1ISG5SvWEwPUgANr6Z6usfcGMG
CPqwNEAGJ18z+nBvtGgHx+SmRcIF7lhNagrW7CXAcouDWbHaeNPQDAZJLj+//mkd
lnBQkR1HlVWEwJyJBOeePFh5I5bFNcM4xVJJdbABuKBHOzxjI4hhj78X97EXFmNZ
6yBTNjfVLi+YJMwuw4xZvlASj26PM7+nhk9Gfa+pzu506NnuegiA6gpPHMgAH9A3
h7lNoNos4i7So9k4u7T4hcpxEpqsddaOWOak4ATTRxOzVVVbk1+wyutuI0JK6XDd
Ndtf3Uw8/rGGWjshlDTldVRhsZtLDEPz4XV/s0DiApEbYtW+Gsg5BWW/NTpHAUvH
n0QY6v312yvIW9AJgR9RA7GOm7Spkd4VMrfKbbkij4bU5vZgffmln3TDxEJNgBDT
e4ULz6ca1OdY50FRk4qUwbOcjQowcsCZnEATuXTbqUfRJJKBTJXltiwuwaMy61uU
6JftHTJUKfcF6EM87fFzds4m83SrghV32imRzV20bEaqv7X0I4GpTL8D5ySzeCLo
sCmirUFNfVIvKQIBllIlZzHfzgeLA1yi3aqiQL+OiInH+uiGDsj3LUoF18Jz5wNz
j0YyvmZ9NZNbQ/rZgYoYSXR+cMMsWbvB0HCDn/ZJf8IqHSu5sLw0WFdiwm/cvOE1
rzZXCBp/d8iS3EE60vy5Ku5icDVhJv0uMSfQJ2o2xUihXjiadbVrsCCU2bjqVY6V
kkVcqNz0dgT8pIvnbrtZrtmYnNT6uAOY4iTP6aWAj8YP9dKPo+WwdJGezzoui9eX
G8bdldrj3cUmMJxXnzUbyuxeaZv4EEM6Bf/dykEIXC1f+TXe5khYMep2lzIlA/jt
iGuYyFfPE4ISD22ZFnquUDtVYxbXpqMllH6Lh8XBPNKtNM7uBReDG0gU9XMgalOU
b17haQHyepjXLq8JUvEW4fDnwKgUEI+prAoUzNCuX9Ic3K+x2RNzHSpvTqxMGznH
+RTsiWkJLVruuJqo/NgJofqd/n93MPKJS+G8dLCgmdHHRGQrfzUe0wThpHgpLQ9u
v24qqh0KMyqk2DmE/z24bqCx6NWzTv71fQrq9B5uarxH/xxaCtw4DcXFD1IsChrB
wc5mS8iCS4TuFXAf2S/z//BU5BAN3dmvTVC2/QaD2+FlDIgeT0faDdVwTlSFYvnj
sJGYMNMqvnqqK7p7O0KUt4bNPMUOhEeL2EjrnGXVPlQDB9bnMqRT2rMj0DkFLHWF
IEc65P/paY2y0HR7ZiStV0lrGueOzHhHqfpAIidJxgTV6WveHHosrf13RFX363HB
uMvvCWFt+oZ6Z4+ws6c7htq/7DQmDTZzLyMBlXCADd6PDc2ig74oSHHWxjxAGQLN
V/e3ISXgQ3VLM6J7ZdzbtVH0zhn7YhdzPpOlbdMEfEhysAoRwWFUe2dj3SLsO+Ub
BSqmUtG5x2rRPrQuKH1jW44tyGKHadALyEi04YcXIoaYtvCamKQGXxCZgzfWoN8J
r0O+uEXdD00dK038wZRQuaq7u47mx6dKrghleOvOu4KTU7ux+grdaWTKK+HPHf5A
dJZuBElRT0x/sTlan4kMZVmPsh9/EhTkeT3AeJ1ttPjGt3DBVqYfWauGits3I7NQ
ujAApUAXWILcWZQdPbftEcDG1wdSOji+1zZ56oRiYfl22elUdR9aIXg0RQuBNj+1
T6ObqlQxuU3bOXjjkaaaqqAYcmnzkoBn3vbJujGpmZ2hf1dFUbS/5hZsT6+Zlo+k
QZc3NKexRHoipk7gaEOpqVzsZ0gKFsLwo3m7Vw1Es0+/oaOrnEV2Wyy36BFUXqk6
RG5MF6J3fLZdJuqYKoM4LJXvp2Yk8oD1Jn/lZJp6fgGSOso8tfCaw2uaB0HUlqP9
oE2um5Lb+e6o7W98zBk7XPBQE7IrGytlRCqiO2SMxgpXfSacleZhONjRao7bZw7c
bh51Nk7UDNkGxKqQ289LfOfEXQafOn1XfbBXwC/byDxFa2dSkiy+nBzbGxI97m2B
QuFt8DZaD1cpvxII+kUccOvKfopCVhK8QUCZWOWN+I6Q5RcyHORrrclsoTlioTNx
WhSFe8MhCnGEJqlmYGgum9+oXnfud7QvmanAYTwITZVZvOAjluWIrC+MHNdAA8re
sdOGHS+QuxYbqpH5hs4BGmJu4Vz8vBIFo26f0EX+tv8LVUUQdvZvIsv8URrSgAX7
tSzLzbQ/F13OMs5W/z2vdfVHuXNhSUx3lShez5lGL3q83ZAOEt3ivwkx4Ssn3yzg
Rrlg6OSo2lr3B+5yL01dt/UH+B/pS7QeUYh1g/KUC2NIjcNfHNQwgwbVQRUc2cfW
C/mjxBc7yWOf0whzEBpPaoQH/k+kwjotkjUPNPRPjB/0VVr+SKDndEaORxSzeQYV
TSBsGlAEDMthoKM6amaqBHSvq+Z496GK0+LDw8xdtCQbgtBcQ4980exFEvuRr3L7
a3xHHGJ0TvROLuHNetvFJRWI/I6PpVb+/W0uy6AlxmDky3pxeIutY3lxdeL0biQR
RDLq6CrwaiqXiuLtbt6+Ek8s37k3xac4lVchQlgEVxQfK2Ib16AlYGtYW//EVhuy
TOsCyWvFlnnFDCxCucsQS7w+4Ep3QYAu+CKjjnHIk0r9ZjQ6HV1zrNFT87Xw9uth
k+iYs2swANCZ+UtDRKxUpTe8+5oea1fdJvGiyuB8FInJeJDwWpc+9qBCRcHdTXwE
8Y6amaqR0FpkBiSvh7rihV0rDLinVnxv4l0tONktpCX+MKM+jH2HDQEhhhPuwV0X
WI6OTIRNWfABiERKxZqZlIw30HCGIakxmKOmbh6quNng74lZSjpdcgHV6fhLbePO
hP/Bimk2T8ApZbZ/iLW1AoidIanBPn0y8Q6TC6Rgf9oVwCI/FGbMuUGIMRDIlRr4
O+DclidjGs2lpz2DeSYttw9OJGLi/POZ340RYpTnmIcw+yyG0K7/Ll/de563lX47
JpYmdT5XigCFvJKN4lZ2Pv/vorjj8O8ggq3hy8hfnvmLpmVQwYQigta7aTG33sQS
Yl289DhQ9mVfSjc9ksR7jaOZFcrssiuVeQuAcf5mqJTNOeYQJ2nktYDz3LDEigDz
rcBW0wRHcZmb68npD7NQOhghQsEcyhFvmvcyaP4Hn2lmwaJZee0COMFt++xkq0GW
EeqgU4BF96+RqQf0pbm37iTeFHuWBkBY7yfO9/XnrCMbAvwuIlCuTmAAr0fUkYvs
oxgbco6JjIkjPJQPgWSqR9R1nIUdjJeeKQCBvM5gzZ1Q4oeaARITAwQbjz0j8O6P
ZTDER+1l/mjN86oF1sdFlL4mDudNnzQiT//TW3STtYnfzfxcQfFCJKCYk35kiZk6
DyP1MI+I9wyF32UpGSWQX6YGh255BSRX5QoWgmmyh59FqTYBWErtLDoGZATVDcLG
P0Jn220jTHzWhCpDEEGd1SRZJXD5KFwY3WisUvtaUANCKg9fvr/VhVdqjxAXekcU
kGbmk4IXAIzYNGcQ34y1O9KpPKoPPXm20sftFi57vwRoa8tFW9gkddXtv6WRKuYU
UERppds1FTmEubwt4nwYY/D1f0y7RLeSM4Mm7U5JeRmXE1A2UErFBbLYc6BL+ORO
1TzEX3wUtDxCsoR6vH91VHewHzJwrnnidYA1rZEaFDcg1lpPLFHg4BeAimH22LbY
vMhvviRz9zVZKOyc9h+6hTIxgtcX7+BNXEEmgSVtNpaP5berciYl7KfMVzfNfx2K
bTa4UGdMemeUckKum8zIyy9rEqVvX0rbb5evrOBwfWsDBYlGfMNDvqmtjDVUbjmH
emP8vp17lMlGdt3rrvT+xLZs4Czdy6En9uVq3zJeccrlCzfUaQhP7mraVqKQYEWK
UQpayTimG5n9PcKblkqgNnivGXd+144aML+EoHaUGRz+VzETnM7hTzwV3Wldpd7G
ngoCiQJAmCoLVYqEeDAu0w/PVqp8FRZpoMFE4s44zEr39xLgjui95BEHZ91X1TSI
Y2rgK7zqWgBaNFkt5nIKA/0Yev5gqpXN6Lh5dvO8c1pxTZQqFXs4CYmeHcqYA145
9gUiSxZ4tjHKhKR8XjHQ1sqldtj1elUGqpfyaRtQYB+1SSiqzzRUWY6eOO2470Lj
bGShrnGG+34QHCUiDCDUjMlepwi7Rse3qxiXG4hMD4gnapdblNvSvaKqObMaXr+E
d1y61snHDeFO+GI3/djstsqjySWU6nJVWxehIfvc9sOCNFM4ioLasb1N0+YjilIQ
QNiqAzrX2odydEBV5ukszjN/DPAcyjkMK78E76CIRSSgdZ2477l3bGUxP5/2b4k9
+sTtVAjhPiBoBGeu+JOCU/QsE7VIkJuKM5im2/gQD2eDa/UHl2oM0Rnn/0AYBT1o
4HEJZN6UbBIjZNDiALWUNiU8mT629z/JD9D9UsKz3keKAdF6fkTJRNJ9Y0lbNiNF
qOxiLvn+7oe0vmanV1Cat+MbSeEKQ7+aeBcTPKLrTZ7T7S0aMbA4nPPcF4PxJIKY
w+cxvDMyTVL2xHrE5UkyVhZOqJmhJgvyq4tMTV13ZvGJD4DDob/aS1HoDMPlgygB
VrUP1Lha3RJYlXOdt8YU4aBWojGCFm9p7gXpzUibfpGgjg45XRrEkcVVdkM0htZL
jkKe4Hd1uEQpWOvyMD9ha5k/GMQ7Oow4CJY2wKOMCvMxaNMU16S5yIusGtb0nVS+
2mYmLIWKfTedTu4hQwA7NO33Ib7Bhjgs+1N2lqPVSaCgWDUymM6LVPihHsGexSRG
lOLKuvcbTYDCCU7F5Poavus8y4/0qDmdcqjppc1Tj420Ro0/uzPv86rd0ZaC7ZuO
N7XuoTKejOXPSAvhvI9ZYOWOnaaEdyHUMtlAaD7/s4R4bWVBEmF7wDP3hzfhbA28
QhcAjRhFpVjGNNgJRYiHoJqSukgBUhMAe2rjDEqgqnMCkeo/yBQqUIfs6NLUC9IU
ANVt7XBeU3RfviQD4SGq2+xriOg1ti5lrnfugp8rDuKvn8py4diUCtdpt4kKt/H2
JW6yrGKNR0VAeAAOvBAAwlEht2dKBDKsqf42zCPrCDjqqVWxCM6MwlCm5y8Dw0kJ
xAgUiR2khOPqu/1SRdiWmMdppJB9iDL1S3uOOQB8HNRIoxfK3+hGonte+gCrlrVA
laQ9Y/dpyXai6uISS2NzyVNI0vXXn0JDxU9EDWQxjzN7Cwb8w5KFs3+zc04r0+80
p6C3XqaUKnRoT7Tj04U7o2ZQBW4E2vKXi7GFtyCM5yHMwLuV2g2Be3kR13l9NK/D
XFQ4bYK/L++/Qn8B9Iuer+qgqVQ4hwJKND2zK66yFc2B3ADVtkg/RPefsq+rzPz4
+mng/LE4wni6M7UkmAChWFwqqBBQHx7aY6Y2FL2IYO/YUvczC5QhQwBN9/c2ttUl
z0QKvdDWxljZlmmK++pw5n3bC4x+k1if8/YnE+5ZbuSuSLZLJDH3N6bnQ+aMcakg
lXWdGK7D5HJUe14rr3e0sdn07NQAWcDZnLPSVAT0wiUwX/uRx95UM1SCM+1v+rV2
nt4pP5gkBRCbPt8XLSEqdXRyB4Ujx9lTaqCA2WTAKdchNpCrRaenngzCuO0ZKvZv
lhpLGcGfH06ixqJ1KbJXZOzfws0yPjfpqpDrgzLQwe3qV96ssn6A3uUpKP6w5afE
rFhvd/dF+kIUCgPmJjxdur5VvRcWbp0KJ+e+Rsh5itTk+oBPY8ulGf1zxVMdU35Z
9OUCjxOH3+H0IrVAlGwfVlrI2eLnWnLQ1DrNurACmDytOYjNl0+A444cIdbkThNf
Iw3x+gB/peWVlnm6zHZY3odolM3ZA1G4xlNAsjSvUtgf5QV8UyQKosozMroqNTmD
Yc8XtUTTpTMUokdqPsxm6F8AkWCq+xb2XHQeMdrVMBn0GOODpldSA6xUgSr7p7+8
4ayWxjQs5fY42XrabH4p6UtKnyYztd8uu08M7jzfr84dnbzzkdbIUxAt3ytGt1on
WfB1IVtQUjoPZhNjFLwhOfJBVMM6OQ52+/5MZDleOkw8tI5y/odEgx+gjKT8zn+b
vfyy9DVjjdAqaSNSVfK2akphSQIfthAFZnUOk0yHeYv/QuiW31axrLRhrFHCMF1n
nS29AUkfKwgA36+1I5FS0z4pgBnSQ+8zilyQiWM+1FyQlmgyNRcuh6KbMxUCwO/C
uU+x6a89CQimuYcytJxIFos1Lf68noVIQ8CagBOoUpZDWER8zmfDw5dIMuVKWGZ9
cNSYDfvCGDlKBqfnI3LwLHAyC7OVtu3KA+07QI5RPL7J0bJsFsMA7FbDctXkp9j/
xtbvr5icuVECcdel/gLcqpX7czvzipkg+da8xz+8HrdWJ2voQLI4yn9lNOjD8fVs
2IMQNhFD2a0Fl44T6hRJIJkNmjl7zOm+UP6ZEoYesO+nFVDsm1M9EVERgs3Oj13E
ZX9QQSFQorzDv0WkqbJEWT2EXthFICo8nYgUK8zlvMqhUds7ltQPZKhuw9YDKy06
JrbPGTJsE6MIKZ/joxDUgiTEtxziitlMDeuWYucgfAhFoF6l527ovQastqsCTukI
sUfpWRposuT3SWUToD3hvXFdu79PTXdKn394/H6BsBgKLM+i/siJ0NnfmhPc08WO
lueWjiRSC3PpeT5UxthtkHBVU7N8uy7QJl/Aj4jAmQBTNVBzOWK4yOFXaQh2W5j8
1VZyn6I0Wcm9o1Jh3d3ZltJH6lMQ1Q//2HFe0vR1BjsBbgjNcuiLTMe19EmakekH
EPdQ56ZrEFSJDyQLlU53lvHbKoEwCfPckvYWTMOQT3BpCE4Iw4U0jdDHiMcGc6u2
LXjl0QTlUkVOMwx1XynJ8lqrEUOSqt9kjLcrDzcyCnquA+yoG4MDCwElKPN1h1qm
llZWgoD4RFJbhZQCqXV5JRwDushww7FMldYyi+tJE5Xe79K9PGP/zD238mV9wXkF
yMWn7hSU+Z5s2YEFsnBocZ6+UjZ2b1hhv/3RWM+XpF450K34yNH7jjaYcxT+gQLn
sBNz5smi76XSpjMLV2HlqKuZM8b+iQu2JbvutiQOUQQbIiml8qkOgezUeq4anqmt
HyV6KzydU5aov+t/gIj+ewpHwyDALC8FYXgR8OS2i0shOs/lY4hrWHqBuJKGVI7e
sB7e4tLuky0dz1pAjcgm4/vL2iXZs+EpEGbAvQ4l1dC/nhOHIgfZJizR6zSzXprN
xqWIKwZTf4YaiR69GR9HLImOFHQhYSxixzaV+XMYA6BwZ8GUfdso8vaJ4chFHkn0
NkmnmyfL/WBm49FY+g6QyqltfQOJgY22REEhqpsbeIMmqivnAoQ0NALaUUuOufza
ymNl6f2f+W5ZQ3mMK1HjJeynXI57hzBvnJdwsJjCwM6KIWVIlDBr/1CaBvbW7G60
Dbx+uL0V23nuaMNuevM+/XgX0QgNhnLoyPi74BDSVl+FIzwu6Z0nWsSYGFADudaj
9fipo50RQMxavKuq9cYNl/3rapFJWv4w0pZeUiZvhM/FJET8Qvi0xkCYA1VuEBP+
okU/bQa+LSWcCG83kjZ5rPar3wArefBNCEnQTMMLRdr02/zot4Cjz18WGOCZpywR
T5LQ9x0rX+q8N7FL/u454dbWXek2vLsiVaCwUqNGLLC/rzpgYDYsUeJ62I2rWrVo
RW/UDpIH+jM/jph1eFi1YhSCILeaetvhLpqepxZ4VakSzVOLMOLtBYgxWsAcVwXs
4oqjMPE2qXzy4cQ4uAoPL+HHIY8rvXyD7GuxcMFMSpMqUwdeH7roK2LDWeUvpFYT
XCynHNT/CHhOVy2oNzqAhwvdpOJiNCPz5/j/94dQVzAYsINqIJTvK0QhH68TNRDH
1ngqQup1MI6iST+sl/L07Pgv4LAwA7I4Wg3BlbBpgk/xx8ttNK1vNhEaqYirWKRS
b9rLLpA1mx1p6mHtg7iOVO5RL1n5vuxaJbSaB0toj2isDr3rDbIKZ8gw9P1z4WlB
iMqgXNQYQi0AMBdcitlsulwnP1NSXvoRJcPRUb1JJ8n4bmZqj6dJui7gIAL7ggaV
AZa7mMvndrgIlxHi4XgZX0hYZkCPCwj/lSO/2kvTgz+QuFgL+u6Dfoar4mpsk6wP
1UqAjnIaISlLtfvhb3J+aFiUlY+kHd7UIFlhUz+MQBBmEgG+YpmNJCuHI+AK44W6
KJBLsGSzKpMw1COeFIiT/AEZi7HwJ/le9KDzsF5Vwexj6sLfTMaJ/UEgv34t2I0J
YRJAMHRrplYPS9zFR05WZLSMkXqPQKYCqxZyJN+tWstDiQlxy5UZkl4u52FlHDuD
XB5jEzlnfr80TeBtj/4su21pq8ONKyFk9z/KALflGI0LaoPNJcKQL79yK6SC7EYT
lwfDWQ6vZqjyvAl8fEYwCqajvr9z0wqIJe1swhwa31u/TDCu/H4sxug5DA7Om14l
9MHt/N441QeIOUcnQA0AtbKjtx9/BMrAaBLtQqzkIZ3gqmcomlfm8rzOSMVMqsQY
LoUcfve4zeZ/oOmOHRWTvaMAPnOzErUDu7lkTsiLcCtJkTlFwPdxqFSg8LiJjZd+
3nsqunHE2G9d7iX1rKWnKcncGdCZeEO8SteRm43D2qIzTngeA/XuYkzd2BCwFjGc
XLRw3O22xPsRB2V0d5HjElInM1Cl1AQbmQbV6G7PqhziHM3hQcvwYvHSIdyZarGO
qfD9347uJZf/DiBZTt0/x9JfI0E9TwS61FUzZGlj8UsBuUNBGMdNZaTqtZklkAZs
4uLYa7DwCheu6hfE5KWVJQ19jZojeJVDDg98U/Az96CAVOPX0BTNh4R6EmbgYe4c
t07sn9U+z6tCMRn37Cd248cYcQ7oCPUdyItfq2WGWFRNXAL1MGWi04C9ckSiuQJ8
+KIX2Gc2DbwtC1q/k3xFDDGaHl+YwQc1R7IkuwyUA8PMxiF6lvoGowkDFpAWhbXW
9LhvFqzFQCvsDL5rs1m0QWLCG2iA9pyopv4Sqkdvmxs2GxEl4QWflF00U6goAx/D
2U9NYgPOiroSLCYmHnu8Ev2n5gIzQNUw6Z7ohiAB4u/AUSOkLq7xnO9sew0wTo+N
zKZiNCimgeHBiOuiY9bo5FsS5GXPva0MbdKlb0zBx301TYIuScYEt8GxFEidfrtA
5fv2la81YotDMHMvT60r2YEYh/t0znC5CdVc/gZVapklD42O4OrdNrIxgQBHYlF3
eSjszBGlzYU2aLGE0YTnTC9EgTthdGv31mWgSgvMMqamQKmC4g2ChlL9qfzqMnBb
igVDAP9jWWg16xtoCx6P+2bp7AlpicBwRWUR53OoAHAt15+NpYuEEkDYZGJC/Bk1
2IEDjdqHAOOk+t0K9aiXEL9/CA8LLtHxiDFEdYmsPLq2fA5NeMGyI6yiR3mkTQVg
ScsDNdpAK98+LFO+ek5FBKQ8SaEBjf4IXVKvnGKD6FrmVu2JbcY9R4OTo+VX88ER
8W5f3/Jd4rD9havvh/SIvi7xzz/lg3zujjfiJ/dGQw2MJ/lDAN5tvTtthtNHPGqF
9jQKJu5UN1pQGP15xYwCnhMPqVyOJBmRzR6QvDhvVAGo1qkNx7mN8qRo/uw7msNL
RncagyAYrWiVdjJhB4WmoJOV+5N6VZ6hlQES3mdWn/FMWUaMOHtHObs7w3gjHNw9
iADSSmK4b2eKn4xm1V4eA+ML08nv3VaclfPZJrE/H2/vsyre+JDpFI5sDKT8nx/a
BMMaOgZzVJ9odZQy8d7kITCZnjOOXLd6Fz5RXuN0TCo7IRQQeXUCkBinA5/KaqE8
E15TjYZILcrIgGua0a0ydr8g2S5lUns00rroK88rFrS6/Lrrp1PkocEgeC2+HjSn
eONvZnj1cg13BA8Rb21WseWe0bITn5jDoRQjHh8n28kPA9JKDshpq6e7c3GZGkXB
fGduvYFSO0ELxBsfDcsa0LAuTbDI0ZyWOwIkmIwlw5jgPoU7s3pwwm88E6MmkEPN
KK8Bxrpwp5KS/zWa/W43TLp8eZZWOgQAVB7vsIZqZPd7LuvjT0pk5fNrT+yXK/N5
18QFslhILXs0bJYjrnFgTVuJoMso/agGhZmtHlT+KtARLFR2y5tpr3VvBkDeRcDK
I8bklFi/O0hdKoE5BVC8uQltXMIsxq9rdkfRqd+Javg3oWFatlnBq0W5TW6MxR76
nVS5WArRjN5Jb7al3N+KGN+otaPLtU12ss1dEzLif8EtXMr5bUK6oIC1QxOt153f
KZ3zYsPv5LzYT9jBYAG3L+cDMCgYcgpFPiMOuHZW2fcc4xIebgQxyD9S8mQhFhCz
jf+Cec6RdvTWOffwqRchyyuqRyf/ndt7k/rxf+M9GlMiMmivFkwH1mKy3WjDl3To
ngqrplhx2Z0cVihyMP6IdPympjUxodqJ7pgoxZOUyBlhrZVwfyQE4HZZkEJc2IYF
lnvZpgNvu3rnpDqPoB1QSCXR8VopPCQ+WFZh9t8whEA+77P4yA4Xl6p6OHAMBNvO
CFwFgxMurczyPlpuPahzaLZ9peabNxr1akhn0XkE/FO+KgEfWdS+UFi3sZWJH+K4
wGqxXnRv48c0xLMOdY7QDsKYIXe0rZwmpq6yVsxEyLiD8BXHNOTs7lHgZJyn5Eo8
VUm1mVEGa2ez2lf9G9qdmThVcdJuVQSr+x7lKy2QFhbcjlboANvhBScZHrkzkuv/
Juqsfw00fv304kjDW9+GB9m1DqBD8VTLRsOpLpXRTRv/pJJ9ymnPSRXdGmbf+bpw
amEaGfc2GFVAsXxeNXCb3ee7Uz3eAXYivOn/gUWpY33WTsLmKP13BQCNEgcJwW/x
6VWFHZmRw0Xq8COXZaI/fCBB5dFGYkHD0tAlX0SqPlT9nAVkr03cd4Kv19o/3533
OH+QMjRnuOWo9eUMDfRYWQI25ff42r8/TsZBZVfOJ2fC5ecc65ztcRo6f7FbZ5Sp
gNRyoWY86PsW3LlinTomjHbZtFR3DBYDG4L2xcZCW9nmv4w/wurDRGxylHuVXKvO
fgyzOTJxgET2rRQLyBAlS5DxC6CuCHNRqP7rjvn+W219kFzp7+8FW2Dlxx8DrO+F
+2ltn/Ael59WNmuappZgZiubTqNtTudPfr9XX47FiH+2tk5VtguMtTut8mx+ZXqS
KB73wCw1e1xpInhEXjVYjF5Vn3xq3EbBMbWA4tlABJayHzUu7AcapRf81GrgmjsC
K5y7FuVH+YsM0Zq1CaL9sFvWy/zvROlAekBHv6aXthl8Sxxmclu0Ybi0FpRT8t5V
3sB3JjGIaHfG3W6XSv9PNDXDzk/NkNRLQs16ab11bm0+pAj0gI7GdEOhmMW3tkBE
+0i5J+zRWkomv70PBUV9ZMmih87KTfn+mNLmlkIjySaT+6tz2yv9pLYz8m0oLYxE
nelxRISZQEuuGvhuSdzbw4pPhh2fTfQcfFXI0W2MH3ibL152/HNSkpAG3yOqT9lZ
UgO1ZO1eqfF0BnQzP8o6BIWjZgYNrv4cehyZWCkVUwhj4ZdYOjS7F+tDgPIaDECB
l9FmYkdOGT+xCRe3+2N6HJbQoME0LB/m8MXtyHsnTxvhrgTEGAoUqfKNH5WscIII
Hn7xymr1YJc8stxFKeV4Sg2P5UARpAnVSv1cCDX9L1MsZrqRVL5HjGV08IAQW3AY
W/LzXabwZEmNC21qed4ddw+a03laPil674y/DixyOh/vhXS2S1N1vXz398wOa0PL
i1ywdaVq6iyxr1reKrpCOaXV0EYZG8pUoawCee9lHmv93kufORfm8G8d4gKQ7R8z
eglYAcmrf8J3kdzz5uXDM1cne1b70aoyqpKld/hPf+O6Syzng2PQstK2IZWxgI4d
7gkiE8qKDdtXlvlXjxaz3aQXL2NGqS4WjfPXvcqgD0zDU2NXqKamhLhvGSj7HBVk
7JQnHS93aUgE4RPvO9PAcYUwtNBcd1jOfWaCA7fpBvV3XJl52rDltpZ8gYY00eCa
P0CPObu5JaMTHJkYsyZfrTajVauZMZmBKXL1UR4ykwrkkNlsW81p6RWUrgSX1pK2
xjV2rQxQjXCXhIevnaigxcCDscdnt1W/WGYY0AHDqzIoTx/XR8TDk2AEH3P/eOjn
n5PX3n6ni/c38fciWE1qX998yqlrRGx1WHwIK9i+gk7YtF0EGy/Vn7fBP7n2IW3w
c/BIV80TvkE9IdjckdS+W4HgZy1pdKdbZwjiGCbTffdmj7z36+3PYi8shcO8SFF4
Oaa0GaPQhuzCkXB04oWoPtaWtoudB4cESJgGX8JX0Xx19i7dJIkrvX4RlEPpo9Wk
HgvfErgscddineLd0AndbdVTWrUwKBge4HtgVCRxxvmeZdCSEqL9YGJlHUxTjG+p
s1k88UD7tDxskObdwcWvIYHCPzf1rHmSCSfsJc+NoempikPa6glZgyM9LfrckDhI
3V9JO5/HiFHt6RqBHIIc49a4D5TBCXbmG7ZErdIPU1h1KhLPL23e7ic9PV3sJBfj
wSfXZkD2wLaxfVJ2prtY17bhA0lmYvPhuwOu3ZyDH9yXkTIF1nCtxu4HopJuXxP/
B2hYcyUz9OyCZUBIXPr6xr0tvBeD0HqxAmRTBhdJJ/V/a4+KYsUt3Sbj+wBKIn6e
Xhp8zUDGJ6oqSo9J8FHvHufEF5364REPtPOe0JyVfHiIKOpNK3swU8KlUGXZgraY
AdD5U4YaskLXFkhGRlXxidMY9XokLHD/NPttqgl1eMXec+//ytb6feoEYnCWxig5
3HXX5BPLysk+SB6mq8FZg0m+ghp5G5D4rXLk8EMF0gO0dRpRgt3YU1GtcboyIUkv
d2AbuLMF5KhMqWii96sQXvsHxjQHNKxcWMhKxQuNdb81axIhcFWtGWwz+MVvhIgt
NFx+9fUqZnTwlXfY/B24qn0BeJoFk4WHysfA0DpN2p5FOlM3lbD/zLCySdpsOqhf
fdp3mmvZst891u1I8C2ynceefxMXmjHah2gLJx5QojjEMQv9MqhTWpP9JcYZK6ED
w8G9WDqEaredUJl6oo0cNGmP7qhpOI+eA7sdHKbKakwjwSpA4Iv0uiVLhRUZXi6O
gcpvkHFNuiQjdObjTbA/c8h9oaMwmMMsG8oXYijtsNZsZ2n47ifL/3cAznrhedHa
l5sVDVkQ+v4PLe61IF/mqXgyXoaTFLldUrGd/oxiKDGKdD02p/Hm/gHFuddGXzRy
d2+IXCSg7pUCsSUJSYqO/k7r+Mou7riIe8BRKP1HELaHsFE680B2KcX+VAJM2LV6
UthMHc5jdU8SY29MN0C73Z5ksJ2qg24xYPZK4rPURoyLXY29v81fyiMtCk1aEeFh
30YLAMRQ0O5m+uWbwslJ/MxO6E4eymSWSQpYBFTVrTKgn+aPHF9xGvdw40m5hVRk
PApV3dXKpNZ07xr1fp6C4tDEZmn4UliAYWPaSjSO09ZM347R5fqENdsbQwuZqhTp
q8jLnobV1B2/MXh4yUNvtrl12R0z1GW52SD63S+unXTI7YOWkh0UZNvsZ+W1XP4m
5/+4iBbGqZs8RRogjV5ALHsuwW8agmea5oznKlWWSHYkBDPf2eA7AE7BCm7E7dHC
/V9S4C2txzlBe2MoumRunuDU6uVbmzT8pp+4WYbl/APBu+elYkkrIbd++NbYNDaD
u2YPLAkm84VZRiIgcbAwkNh2roHXa6lfK4b81lukt19Y53ILt9mTlG3KSOFI4iaC
39GX9pcuwCBiJXjDfpEuLbkoZyJ2rGD89Z8WG8FLNY3YpZhRYtGcn8AeYaJIop/U
/DxPcXDvbziu7g8sfSemA94Z8kKn5/rnppqsZsk5SP1HXVCswvWjwjBw/Z/LwxkL
vwg67h3W8unZ9jHrSAEvJvdM1bPgJ4SBv2/6//IwKaACfZrwy2Z+9MvqV2yC7tsB
sRq6l6Jl7pXftzcTh/8tcqZ2ZNtePACaKVhsnk/vjbtkuLULNDf3Zzsk1vLSiO7O
d9eZmSeJHTGAp4bb4Uhrt5uN3QqvWya6CA+lHP9RgnFtqnaUAk6XHq2H6rR5Ddn+
lrQQmDo4zdM8SnYNgceNFlV+PGLL6RQ83P1S9oxc0DGv9Jk3b08/zq25Flm9VYRV
wQrVWCtJ6YqYTRNv91AEOkmKWQimzDxE6riHfXfAPQFpwKj37sVXh5nkFNAOZAER
D54sepz13+ui1lL5LKi88v23lG89MtR2OzB14IGm4Df3qWE78P73io+/l7I9lfSD
yoWwQxALz14dgrvvbwFy/UpCvRisWIbg7h1nWtHabPGmg9XvtzieV4xLu+MkIkjc
AxIG/ye5eZ4HeqxRM5Hl8IvSwy0+eWzPZ9AjhjaF7z2AsWUphQbvzGacUyHsCgZq
RuCLHnOw/PmHpMthhyl3/lWrz1GbFAecLtrSRfMBayNMWDZEMvFL2NVxN64RokKU
8igEHWjfHREGTu3HzbuXVSqyTNrXB/zrIr0DkaLrAO8V8AwwU/k/uk1xqky4MmTn
7wbjmOzGheK58kWIb480+T/K5zhL2rp6M5kyDWJuVU8+ITcYIzznLae9NDqd2MpB
8Uvnj0g5YLx/jY+D0YNXv7YnBMCPD6PROExwETSSRmbfvvo8RuNrWpGJBp3QJdsP
u93Ivnoh+Wk8Qk0+1ACHSrfFEmr0YI7BgPZJcj8j6Nuvzja6mkCKjLYdtdflqJu9
xtZcsdgd7IScOKp260zKcWkDK7nL70DoY4182GoZJbIcHxcHFXMp7mqB7SNF1tEb
eN9AflrmMy1ShAPsaqz4rwj2s8CvTwCK+APkSpr1ozFLBODEpm2oTJ/xvuHWVjPd
Y1MjqplzBOp2a4vm/SAAijgYKNcN2SuhVfkLKDME0+fUhXDLTSBzadWwWsFrvzh/
s+rOMucJ6pv2qucCCqqpDE3L0YQ4r76Es604RpPgvNqIbn04ZRr4qhm2EI81B0sk
Ys0ulLBM7dQUCoKQEzhIAmcsuCiCmtiyl+/diJCKExCS6y8Ncb9thHHUWCkKsSCV
T69mm7hJUTwe+LajBSQmFXuYL4i8xyzGOyojl3adfpDZgNKg0/cV5npZnubXRZ1U
fCEX71vuJ8kc9dpj99M/6Ugg8IMSLxhadaZnzzpZkmwPbgcHaUoHxA+BU/ZZU42u
AERc981pVr/Yb9oXlKBkeo1ArGKsw6lwfFa/gqL/ZJfqdyFvCws6wRA8j6sFITqI
Ux3CEBdVbK7iyQmSJ3oZ6NV3d4EdUfthQkA307E3RRfM2HRjgw+zZxS4FONPId1q
EhTbljBLbiyewyhSwI5uHUvBNprAesoT85aQIoVcU7QPi2WZDrqKQZVtWZLK2yHc
MlM5NEHVltCDgN2wWPMwPxs4dvFotQWxyUW6XBKTjen6mx3URXUrrmGlJSnpn+hv
i0Ho3GHLKBRWPtr2e4cP2/lStZaHJ28aYUkYTMhgMoUjG6qHdnuiUTyMiGKJt5Wo
oDMPTmylNChQH3IuuNrRi+xZPcfStFj0NToLu/s99sxGi9u8dPInycRCdGVnsnuo
/xfz382uV8kauiUqPyCBhoRWETXO5kMwcG7eiub6HGo87ALrvMzAoLKCgRodHKM0
kGVpRuY+5cWTEe+q5jilSYylND9sXDLwdeVkjLky3I3uCer0b/4dPBpsmUVlB3FA
VLZ4qXPxydtThGYzEGX6UnWqRqLRFfdls2lUhhZ7+pzLUyKielUf99Foer/3XWvC
1HMNE0bMa4Ja1/4VzgE5krDf7BiwuKhw0x6fsS1sYBpWIdPZl3U91FpSRX7Ct9Kj
tWp38m6sF8hAm9SoycLqSem6yoUDHoIgGDcsguPldOHePsTHeDehgMVm+puEDUft
hbaDV9f6LiwBR/XfiSq6cZptZ/wg80nQhzM8pXl8xDpwtC1WNwJjoUwhxJpq776B
QJG2U+fLoll8IM+QJNKAg8E95x784zucBHxSYoSI3BzGxGiwZ1Svz0XuGhDOGa1l
YbRfoTzoQZVT1yLidNmc4j6nO3ASCM6ShfJEe55pyinfTa8t/loZim7N5K14eZcq
7ozxoGIFsNxXgIYzlBP/YkOm1s/MKfklFEarEmpvPZTP3SebV1uoFzmnav+3SHR+
qzXhJjzDn1uFHTLwXo1Nj/TLX1JiMN75/Ty8r37kPLIJeAaq3t2LMnFgMs3Lk3Cg
BAB2xDtef7q1rGphFlXkWZhJdRpXT/Fq2cXEU48ynPnLk0auaD8H60zmHenTw16C
MbQH7cFx0HvRwCF3UMPFLZNfbLrC6Wu1KIn1qDnxy0503L4hSJFv8w3W7L6a4brS
lq0MDkBs9V8Bw2CKqHkknjEzqjEtSETNfwy+sOxAYUSl3pZZHClm6nS8l/lccN0A
2BOymJnjcNwN408OaqOnJyLjNKRugzjmCNng5Vfh40sKHVtzAcGUrJHtXOc4sCZj
h1fgpT2jfrUEI2XHDUUNOKqhTO55rnABjxt3t194G2ytNoytT4+pxxDZlGRq0Jgi
IYlcDyj6vNZj1ScDA4wBj8dsuYjqVNMGLfENeI8iFNRVdlTPwu4GxTLNJxWeyyR+
GQGAfccV4w6cezYmEQZoAxUPXA8/phLWnTzK26exewg8abioGpsZkgCMVsRb8fZL
05Kp3Zl3SDVhn9/EjqHKVddihJO3dIhM13OtLVNEG0C0YAX+rnNNsnJlA9AuGHss
E2NWP1ckTwrHARY8MmP4EqCFs/OKBA506LJdwhPMq7GPbk3CZrJa+s7H8UxbH7Tl
uEzf90JYGuPmUByScHicrr4w9qMw41dKQKm2mCyDG88wDdAZ4klQJzG/LU3gmTp6
6PVdEkOID+0cxFi1+YHvfb+IrxLZ6YByCosIRsP3oBFspJ9K+TfjSE6MhgOIKspl
s7rUYmqnaNeIxJMc012LhqyWa3wSsqJJXe7ZJXIuxOaeZoY8+p9f7Qas6HEsQzIy
9mdlTx7tloCJrhfhCBlDbE3LQqBj1WYJk34SeaWFNUWHr/TmqU8DQ/Iple8QJOXJ
wmEM5PJIjij9zmGXVO9PDfv8SPA7HwgQX14cOSdg2mlut/g8m0UDOWiGVIBALHCl
fUKWWyleb6Vn98AZ3tZri7yYRfJxxuBo655u+B7q0X/A1lA9plE/Osu2xZPSPnf8
5cvmN5KSTxQXP8UOzR8Mt2/PeI/pB4AamoMCIEVr80E2GbuD8sdiMNp1ktpt+iyz
uGwgsCPSJeQUU3YSKQWcnfCV/3rHslZWstzVa3hhCXQSpSLMl82xhJUMJnNwKCNA
L6BVsfhge50dE0hJB0I27eyz5BqBX4LZW1CZETTj3N/XWBBN9dy9XwSUZlk8ssyY
7v2sShwnt93X1eha0AV/XJcMvkzSWjai7VbRxLWmVyq+bq+E3ZyOeWvgTH13usl+
dDdtYNdxLyNHJp3rxvMOlbDzb7Yxw+jz0BfqwcBppGce221og+rHZFW+f7cSkXgu
EJKNqOKw4goKmLJ0Njx9GwHd6zfdUD5GUVVqU1+GOnR6NSfNo92X5NVlPgJQ0HHh
yd4MmtZ2Yw+zLBGBChdRkfKuiXBhGG2rYprgodL/nmmKDOl7if0bmLHI/tAftAb3
VD+3IP7H/48mwaxyGAYJpfCjMbYv0OjKDWlcNnSLbDjMvN+Ctua2lSSYxfAB5biP
d1jX4+Ix0Pc6J7I8gQKJj0461oilD7A9kKwODWXooJCFEou3xF+LPe+w4qYRT5/p
x60RKEcxFk+AbJHH6WM17Haj/mZp9kn2nQil8SDyoRhmnI2GuF0cispPo3YQCgwM
BzzXvq1iRaDMe9hTeYweORXHb4q5l4ETQoefZkhX8qJMoPpW0SwjgsHrehNN0p1V
kj4mRFbfPY6iZAJVmsTlqRmsmrvyMrkxQGZWvIXGvsoHZXafnFUrIEVg+bPA2N/N
jKvmPKlHY7I++i9Ie5ICbhQoDGN90nrSQjyGVBhrLoE8u4ROLC7SNCi5r1XpAPC4
IXRCVqmN6LRu/Knqa22IzuPoaMsMdFUbSgUuId20F0Hlrxsm1XcWxzlZZPdZO0WX
H2GwHwRj1vHmlKoDQFBW0V6h3TsSV34NRUuwQhkYkMITybd/vzKAO4Mi60XqfjsR
P5Eu8Zc0Kw4hxUN6KrdYN0n2gRe1pkGst7BcA4ilYFlKEBE+5eHg06NDYFuciMU2
3aRPBgwo+xTycS85kIB2eZXWA2hBAQCsNfJ09wCEtYChInKDMt7EEFRsFNmXm/iP
P3dtebGA/6wg8HddB9nBxbtgQJwW0PVf9l+K+YqBCU54rC4qVDvWljD0412f7j5/
8H5K3KAUZCXcNRcKbYNwsgWOy5PwhkW7Ph/zwFecnIqKt4JN2Ob5rVfBXPXaPN0t
RLsOf8AxvpBbM+ixLW11ybNwMb3jXIUWzuc/FqDVcyYLMj1XNkCsH+G8bStmSalK
/fuCFpKGQWrbk0XG83a3KcyYisL9hvyo0d2D94eB+MGzARKRxRHjY2NV/QHbcJxN
yrQ4B7t6B85YNTkhsKbTULcTRUIR+svz8BoNO+8jO3KizeKd23Sk17T+CuTJg0bb
FppmQ5XdvPDKaK3aE4IOZdC0Me5SNGQjg+cupTatSZKL7HCX/nLlIxm3qOS2M6rp
gXheGM0zo+nBa9FdxEc6c1o/2IReN2OaJQ8e0YnRKni4YHCD4dHB6/vbs2f+Jg3z
f+3FSHeCoofLILnDJf3puXguGIatnFNwy2comEe++yf0fRdUQhZxY3dKuIARHwYH
/ACX/xo8a6eHjz7nodQEYi9bDPNJT+zNYKNLeQe13KY81Gf0lnXTpXpwAOxRoJ5X
EHW05oBAn8HPn9DbK8fu5Bb05myZZwzGvL675taq2VH2XM9rCXMZLkAjKWyYIbcj
IN8ypglB7mqRaGxV+0FIkMSaR5iM1nh+9+2rknpdHyZCHSU2hRb6Yny28gvm5dQi
45FIE5Z1hgx3loL/XsVlM839TcpzuF+abULA8pK5n8k9t0Tr97+cfPC0KRaNDsWx
vgrLB8/tXmvZs9JS9ScMFMQ024zahGWwxHAAaOfmaEXoStmTMdDYmy6U1qrgaNbR
ErVZH8ZjSiA7aNeFrCXrnuT/1lNm9vrIyRA7zIX5mEF5SiT1FMStMC6ddOCmIRW4
6wlnfqC4uPu98jhsDjz8LRFaNNiQdDqiT0YKiRxXlFfOSnDpyAhT0pYNJpTs3C4f
9YtlE1PiOyz3u38giRma1ITKEzJXFQRAkU5u4DxL2t1bJ9p8gYbzV659Je1RP+Hi
+K1Cb/39h0GuOv35m7KpBhsBIePxXGe3BiVTxt0495mRAL4Dn3YxzFOz5Ej6IFCe
qzQNELhBpAXLsyFwRtqsJG89XKsNfnFMU5v+uXCiRS9lBj3JyP7aNOe0HZ7usuwa
M57ciL0Mu2KJd/qpmaIvQEbQRlD+NQQahRDDFpmKZHHYjrHL4fLLnYMXbFs1Ezc0
UMaFlvgWDG0Rg44grAT6xT1DWSfW+IRNg6eUfmeDMh0FMqSxzG1RyCg9Yq6zFbKZ
Mj7ID+dDu81m2UZcZTnlUW4EsjgWQ5R47iOkwAF5JIobEz0SbkQm94CMba3Cpd5x
5kgoL0WAo6tq/rhTlxdqrD5RyJsGZKp7s/R7dfwq1R9N3VwTqhUAwotER2sPjPwr
ylytlx97cHEbQmJp5IHzMcQ72qcBDu6dLeoayMaX7/NneTfR//iaonWV+cg+GW9+
t2dHMye1/NDOZe0qmkff+wZB/R0wqpNrAJrQDY7uIG8h/ReLEV84z3cIxrygfVV2
PcEhBBS3b+kCB7NJ8TCSaJwGsFGQyFc2P2FWrMgiMxi/ZRA6pX5T07OlWCmmB51R
mS18YikeSKCJd6hqqb6w1dOIETKPP+6qUEaTVZcbUSKVBJrT4r0vn7ORZheyleOq
p1xvouKYw6VdPkzl9AcIvUvJrZ21hgQlh4CEJ+C+1qvc/Nw2Sh16uTX+9HPnfilv
NEYCe4E32s6LrHx87hp4M77Q9OHnHkDHGJDMaODPhD9e9wV5c17aIWg5YCKwe+Pv
UQ+F7HVqJyO3w5AVolosKPhGP5kEaPWMeznGrY8pHdhRUNLVVOY76izQCnBIiM+d
6WBHaKFwnA9vOFbDpkr7POuR8K1Md7vo54gMs7dOwrUhZ5wGBlyHiGhOBrXDVfpS
miiUPPFZvS+BfthnwgdQTP+1u0k0QGEskPV4EmJW5lRRjLllOxfMUiJ4GVtGrlf5
ZXaekLPTr04InNgUD3Tinc0xRSJwE0d5k1lOKRiZg7gdIKieVe1U+MbsD4l+YjHo
bmC4Th49UjmNpUNSxKk0dqEVjhgxeSZgb3bGfZGzSY2wVgrIW9FN2kHuSZSfaB7g
y8qoQoVgJEX5HAq1VefDcvwSw2Hz2U3WYLZS0VplFlFxWlc/s9ERfFgx4sTLAgBy
UkBFQOdT61uoZ85InCFRFtySSALWkXoDRFZt37gESJrUHgAvQrIdjHrxK8NWDTSq
6gkJIHMJP7J9SOfVi1YuSR22P4majapEJm0a2ZgP33UGMCsaT40pVCFGPNYbhBjp
Xv7J3u/1kAk6FsVnPohw2vLSlOc+5s0C40T6CMnbIWDzLJIhycBnah2YUMsPAQ3Z
ghpOTzqpi+q/+2F4vo6lww1QYkbgm5MnX5bKHmiTxc8cyELoLmmiY6aD5x1P40Pw
53+/kg1yZ1e1L2StcjeHmYU5/LE7xcHoN1mpgB23qsTzBQ07EC254kpXao6zZe14
G2NPta4q+5+odEuW82ykcV4xsuOVytAFZRcBriHOb3pNPP3TiDqyyH6LrITurvEH
QHcSZkQAosRfTBpkciMp6lfZN07m2ajBTm5N0ytsGOFVY9LHyIU9rl2viEHds6KM
dtdnXsTFdvfNUuxq+8zXqaa0uGYhPjFRvjCrTSmQERlUmL6LDYNYY9xjnORr4tdK
bp6l+R+28keOEa2Rui7Jk0zxD5RSk8MFojL8vludH9gf3W8yz9vtF41jAo875Gz1
0JytRxyvv/e9bYeVwTydFqXfQ8hw7JtBBAjP7srsewdNQy4hXB3SM9/+lddOV30V
2Ob5qVKoSL6GhHCKbm98gn0l4BJB9KfTpiI9LMozzFuFkfJ8ftClb+OcVBP63g69
RhzOyaW0XII6SOCBz/ibpgtYF/YQrOoZmzPc3ErLCE2xWOUcYTRcy5jScAda+Fxm
4o6uiZuOEF3P+n1nNEtaPPGjid4fsG3S/Lu7Rmw0fsBMegL7P5dLjmqiB33j2xSN
E0Oas6F6W5uValzGDQwMm5qO41vOy4dtPmD40CgVG5P2tvLgtlZUD3fHyNPJlTri
lTB3K3CTcDSkk3i+bj0IKvEfHlyojY/NI3tISl5Z8mS0SV5mpIf/PXAZw+suyHto
JnxrCWr3K/jXJMox+mPTSIfuRUPu3jWRymE6K5pmA6xeHRYo8nOWJnJ+j1ZjE4qa
i9GIlA8srhdY01ESqpxMt1cYudOb0oEGn5FWqBnHi1VoWb9NnOTtyL/ZD4CE0SPV
PuTGKYHIcA2nwBQSPFNltOd+l8mzKwNXUy0RcP78D5vLjVNsoHfCsdFSwmX0gS8P
Bj8irRqdrnljhyRdiGNm+ET9Y20sjk/wtnka6i67e841g2JKRHSwwJza8EUWTNmR
XszYmWgLnCC4wcAxd7CPVEMrk64fVJE5mnUip9pUoxMFQ1/9QyY8oboqd0NuseC9
LRRAUSdDrKCnH69XvDMXgXD6oTWAKVe5pjNcdrWCqtSXRJhfZhTadF1gNUDlEQBZ
ztklvu1OWRtQYjiRjM7iYmVU2s36bH2H0m8zWmTNTl91wefkfaJXTpnMwnjTAb1h
kSCOPwW7fG/em4SRojjG/osbFYOsSegbBjV2NuYo+K6L+Eh7PMrjKd0uAuWq9NaQ
bSOgzfw/EePPfKyY2YnQqTTumSt93DHNg5cAOd8HYHCuGo8EeSHhi/HvN5AUNObP
Sjp6yT6UHFAeeM5vvHLB71jHZAl3g+EV/yoWHH4S5YxJWwr9l2iv9wAtp1p3oRMy
iCajdPu49CGs7i4Ky3SnCxP/Rp7xmqJndtQGj956ccJ6P8VmIDFRRVLAvqgItk/U
EukufPJKaqApjSMJmHGDUbst5erUIbhFoAnBaQw8SJUMIwJmdLQQKmsXU5l6Lw35
4buc2SwW1gJYF++Uj12dXbgKQXdZt1TNJ7grvyt7fATVtRBYQ8cnjBqjRBPLxM7z
9PB9mxETHZCdLjXzXJNNIuVvgPr85Kvje+Jqn3bXiqeXmbM6jAXKzOc+litxpKgp
sGXMn7Q8x7Uxrg4ytuvxlCjGxgQmyoF0FuoRSyg0M5FJnDi95s/PPgKg/pBzCohF
1BENy+GljeYSA9/E6Zz4k4kEVezItO02A1VSxycoEjRRpBi77T8EDZdJ2v6KHQKP
HRrMgYRkxAUzmtTtr35CKooRs/t0EgWi0tsOMg2Y0KA434Sdzk73LBfZGU2g9m5V
5qEXw2EPNXG27lMGfdb+thrTS1yeaiEi+Thqjg0D2CIFJp+8uFKD/Oqb03lI9BTD
m2SN7Fp35hLLKqaJWsmDoJUx0qlKY4pqF8xTtU7UayiCJxWjSQZ1k+gUXxTxhIj4
IZtz48hpVRsb/U162RtxbAkfe9rdtEA0t3rzsB9kBcWxbfKPYY5Sq3LGW11q2F40
0dQIbCNgt70Dmi5iGRExATKUGGW7OlaTmuS+sNprjJSWx6lIk/0XHSlXAaGg972u
2py5U9rzWax3A+8bCCelfHX84k5IkTMds/PTzSTqO51MS/TJuHtyPCzSiHE+PFac
v8U2yuAbAo7vvdpl3TBrXnoPGPXGPi3YXItcSUE+f8iai6hMgcAFQLFUOBNwOA8u
h4M41VyGDq7oJPdwdnd3qYLpqWbk657dZ5m9O05eVHpRwrkFJcLsjwmvxv0XgnLA
hjZS/XSr5GveJ4H2NahnBhpIJofbQpzZpA1sMqTwZialz+RtHv6U1bMm3KufHQK2
w10pG3MIv+oaqpZr6amHiz8FkguQnKM+JvRLPoLv6h6bP7LwUqbHtM9hROIUOkdc
Psnbl2WmK4D2yMUSWcDWcrTbJGjgQi725OW1jYVSyh836k7KLPKEKt9ntdMgNdKo
6BXld/Dem6kOif0f3pEXjf+kNX7+vZcHFkXfRY2SW+RMWvkPxtrCZn1qwx2Nqz0S
QsJhLb9Gu25tx+dohjyADP6689BWeKMh2LfN8pYdaHnG9rRpQa+k6fbEdEMX2Mtz
AzkEJLqg4cVqcBJbDVdu4ChJK9kZFsAK2U7FyzgnLDk2o6I1cQvumwCsUNwnDHiy
o+3WyiUmOlr60cGvWpmpt19stuTKhpVymNwbdKAR8yIGmaaokYiXa+ZiOVi4Qzfx
2F31Jr/rjsz4lKOWDiCGD31cpu9JW0V4NIA8+2etaPynZ7VQkPQ4WUKYBg37dZfY
wePCnxbqHjs65HCGmVf4C4oClTV1CwG/ssJAfyQpYoaP2I6NqhD4jMiIjz+lgiAj
igPCZS53bncwiwBSgP1NLyo2B46TmrET/PFoP3NkOet8Rp9g66Q5yLA6uEBgHh8J
btLihaAfpa/eoWk82DSVbbXhhhNYsTPtPkSD6a8lkAdM5NyOTU2sZ0W0ZeDXiiQ1
CXqHxccL73KYqZSuhFtFkwGERrjAmIo0ozccjlzOFximpOYRCaoggg+GzVlNcQsB
AvjXt7cAhnXCSlWQ6OGm5PuPM7dKuBTEgdGp7X8LmT1cFTs4UvZrwHGengDk1qke
zGQ1CCIGu1EpC7i1B0DJ3tKVgtreeLpYBTBagFWZnRfrh2r4m7EKnwYMIq+RDC47
mZeC3Y6pryxyCIy0EjtXvCZDufTqEGSjBdRp/kZlAfKKKop5pjK+FQslEq281jPV
Th+IZQF4sSueKPw26CIfvtQP95fIoVfd/yQTfI5lWQAE1Bt1axoskSUnvLLNdgT4
sIZx4tQEiGD6/m/MZhaKcDEXYgfdOxkxsx/Ko98UblBV2u2JjNCs/qivf2zynL7u
OZcFuO4jilRndSZLmIBM+qxMXRimmZVlZ0i9odV4WAcnApdC0RkhkNtSOAVQUpPn
inH0s7rEYNSo8BFgDbIqIyyXRzqc4VTA1uoSg9phTZPcaG6JpZaeYlmcsOyKL/Ye
mtJD/KnRaNy249EyZyKdaqTz/PyNTyz4adCpv3xvXvaMYv0Fsv1u9XPdXwgn/4nf
Lve5eWf8tk725oCHipQ6t0LkqfLW/OyTswq4PKf0L3Af4LWaHOohpck5gDIFYoEe
+A4o4PibOyIQ3s4tTMesj8FIlx4uEK2VzsQZs2kRqGQnbP38vk4jyBNrT6LLrcRy
ZrvD3gYQsLQVmzNjDXsqOQmcvYbQ1nA/XcDp7OFqf4yIKdkhCE7O7ejPXk/Q2NDh
9eYMZETPDbx0+VEwEgmg5LHAdNQX9zNXsH/irwFaDev5/inJPHl9PsAKXglpY2AW
lkCMg9MQDcbRsvRxDvk1YjCbQ0Fn9y4a3kOnHCZFUvc3ArI7uyAYvMCJEPJtLjpv
m081YvBlJdJ38EFurx1z7BFx5FgVAk+93cfeDCx4c0qzDSffvAv6YDTEql+qX0qd
TgpVd2T+oYOp7DyTSn2k644JGWyfYlkDReaBY3/1agQrvblYYTaXw5YvJkhN4YCI
FyKHggtHncnQOiZIIfWpsD7f43G8TyeqkltJrD4BE0zSuyauEBhVEwt2+VaH+gCS
5Vz9tThTG+szzcuNWHwpNBsDkwZBwS3lUKDFPQrOnvy17P0Bok7NdoIZrtfueC0n
YT9LZc/YO3eGXCA6pNg6FMIWmIVCLD27H9t387r5mRfs+I85mkLoJwl7ZZHkVhBb
a0Ae2I933Gy6//pbqHM5VFE2tYKqqRvB5FEgWYqX/XMKli53nbt/roTfiUBzL+eL
9oHIctmgCs6A05zI4Gyf0BaUhZJ31npJ2QIh7oegZ/cS7vxQXR3AQP12vToI0xLw
SApiROk9HCmgeXJNryoXMaSNRwFjQdO+sZ/XdiXi7iNTnmsWaJRoBgZpOTcYXJU1
j63KyEHuQoebK93par3hYf3SlVhTeiIGXCihVtbC5++rbe1GZX0XqZHIO5S19Wql
cSRV9veE1zr/+RihBSq0OGdJaCcHLVradHKwGbPRVpn0tEpGi0hT8r3M51vuVANd
8+tW899EfoEjO1qceJowBO7qNW2vQaIxTJUrdmbnuM0BYbSPgSR734OsvMkbx8pN
95yJSaHRBVaUdv+ejcrpeDzvFkkYkOecbKLiB6c4lmEXHKdxBrwzVFMDuktC/DSZ
NlaVWawq/X2HaSBobjQkqm1X8tnnY4nC5FE39Dthos5psjVXjj7nvNNaQyACwYRg
h50E1uMBVvti8ofqW0v+4BAYaFlWRHCwbTRrwVThUHpBNIKmt3WWwWa71MVV/WVR
NgdI6Ayz0AW+lzc04AArszsKk5XHGXLgPk+wr4YrUDZjz7bZ4RAvfccG7+LFBJhW
rQYz/XEskLIlgbyaaZwRNiwmmY4kOPUiT2sH2R9IKdK+++xHye9aRYB6/EcfBJXN
/u+LDdRnuEbLt4FuIUBmu6tsnaMn5qwmRCklkSXAx3/veidKs7EBYDWM8c9VKJv5
V+ezXWEpCcsMKRsMnHUINzqZtWnmKqX5hBBxh++GuFFL5Bm0rMyP1chUI5hEOjXt
nHC+S1DFtRmwqVgE6KhAfrjy/Zxr1urepk1WWmzexOvmlxPo6HJ7ubI73/uAWYrB
5zAnojKWgPr8nNbPhn2m9ABie7lctlBYeZG09xv7gme+gAnBftodnh9AeH7WBYpr
7z2DMdVfN9U+O6EL7rH8Oag18UPtr5UwytZMLWOjT2mZWs+Oy+REEVObGZlEXpso
5dafHXMqBk/eid4gBFIkIu571+DvvAcgX6aB+yaC1KjnzjqbAfbzX9j3dVXsr4hD
b1xc42BUhmv4xmBkV/TZ4bjqI4rxqVLbjr7x1fU6iKyqDUupSUg+Ag4oh2K06L0u
3SNBUkOELkPcJczxUqwLS6Qhv2noKU2Q8l3EPNS4L4snCdDndDA79KauoyngBnbF
2GcZOB0Uq6XsJDSWHp0lQ1a6w/EmUzN2TlfaxOWneVhziUBoeaVLW/7o/vrgZUrF
3TqwEa4x5CGvuxkcLtz1n/3xq7Vsxo/XfT0tNlM/00Hrmfvs/ThjYEnOKZKTMqUW
FrfGWAkhnK7ZY+LWR5muXSfRAMh9FiFImaJ5WHFLzamagt5uJ9Ti/nUhDivgFP8+
zjV6vIEg8Bj0ABNFNT1awvMpISliNPlVoemfT28n0H8FONFA/kTcB0Cwj2ZBoTPg
q5CKVD69lrFZMS8t4R068de4RdRu46QE6p8Ki8rkLSsbMU+uKmuu5EeJKeXifrCb
AB0fFJBP9FIVedG2UMPrxoOyQzbqoZJEl0/tav719m0l4q95YgOcX55bvRJ7N9m/
rr83oQXm7uB4ZbM8xnzTyCPQcroeACpxJcQBYBPQzYFlpTv+iy9HPyOJp9q2M1oD
bMVZQC4EkvG2DK5yrtvWIrXwPBxSGvZfAARwUavibdABGcohKgXrnzY4Nzdg/jHU
Am9Oml9zx+d4SMgZ+UqOfRktbYJS3FPbxr07sM+XaR056YSGZq0yjKqCwFzldZ/p
vHgDf0/qXvcjtJuR2q4nUZdTJ+E0BH+QbtP745V9s8Hz9JJPsop6gXFMBzeF+92P
d9wQYP+Xkfhrabj39R1kdCXsAX8vQ9r8MSV0UcPMNspIVbTOBC10wp9Ej+yWnkDg
ScDt6jjREIFgIWDgv1jPt6fXfyDI7ZUPWf+9+q0mwf9jYD7DVo8LvPeORUyuOO5o
IfTWdCvhUYf49oLh/RczNxP9vozgK7m9fU5rShKzuA2KbtiwV1dI4CbCfYBXqPrg
tFeidx7rN19rIuJtTUFiNTCRPFsUIJWT1gZFrwqZwhF6H0pZXy6AGFqsZ4GSIOS1
1hZngOkJ7qOjujfKnAG7sHatwjW0745whcGepJEPonhSgr5hlBQoh/KjTtotjNsr
PSKAGREaQQtHzg0CdNNXAE8B8kqWLjV4Scg9NpvROOAIJQlnjohSFU6LG45UEwhT
bqE5LiL8za5Me8fkKI5YYd3s6AK/cGihFTc4CsUqHKvaYRZYVfb2TNVoSh7Hjcxy
vuFxsTWjuK3u+C2yEwfwpKG2DqvZgsVom6piCuMJpQqW20Bl60/IE/B4LZGaTOi3
fcu2s7CpuCvDWcCTdVouQ+dVXXZN51TyQoC8qbcFhuZjDo4JGs34cR2BbYkuvJv7
8QLO3xnEyxN/LINW/aFnvi7Ju1nN6hXxu4GlmqoaAGFWB+1hl6aLyO5w4oomLbxM
wu2egEbwoijPvS4TRlrl9UuDYEmA733Bq9gcaCd76H/hEYylPGHIlLNk+O/ir05R
VyDG3aZpQ5tjxcRpW4wd9WTdFSolEdB4xSgavPrZBptKm7j60oXRoa5SAEIlnmSw
nj6vZYzdZVcDbxrR2dOB2iMfNRqoPE6Z23aIZ8B5fappdBK+MYuheWUewq9QAlok
HpfpDX8f2TaxkYt18y7TdshRVHLJTlcwM3/aNLtGFVUZ67PoM8w7jcIcKBamlGrZ
pShtpmLzVqPBkP9Wu2r/zu3kgpm0Tit4Nk6dHnnpVN0X5fklw8kXjlnt1oayivEL
Tk/XMH1TNPvYD0Byuycb8jmNFXHCPMcI4gdw9Xo6Y/wU7OG+1XwyjoLeBdS/js3Q
5K+LNZiuC5FuW1apUT30ml8JdKrMzCQKtTT0fULT3obtTHka9vh9hHMDeHu7ArE/
/ikAwRaprN+J5H3rU81zJhN90l0z13RbmdHL+zcAJfVpdMgkIBcE4TNODyMYnXub
2ESqpR8iEGegl4//0a8v244KePlmseetAYtXZfpWlI0B6GkVQrzDf1Cr4iI9gp8K
/khrPOWLOJHlmVlXmshAu8FDGimcnAmmLaHqVAwQRBjZoLyOUJ7utPEBZpJvCv35
JNNjRg4s71kxh0E9sTDp4fLHyBI2Vy12kzuRDJ3f7CnpGeQYorhVRllK+3D4qM2l
OndKJoS+g1LYf4BCL+Qf80ggptN+XcPUVLHJkDh2cYGGuI2IF/S+VR7XWcQKUmIh
t7KvsOHE9rChhC60oanpqjed2FTc+WFLXzcrNXobYUiH++QGCinjLaiBBQIpNdPm
nq2KTWQzNJwgqEzaKw3KAv//IQuex4jUn6RLMn3UgFOwoE/nUX7JMAiKkW1IbV6n
FxK+3ba9vRDmInSaMk3YzbUGRBEcl6bwc8xDCwswhs9324J53D6BsxqXtI3YiPqZ
Ve11jgEjlpjSGgni05jqxW+RQWPVRxjqTySbzC6LdpRr22av2AxF8taAxDdXlSbL
J9UqFZQwDynJNqH8xkOWsiMR0e8TH+siw6w/NAX+W8cm6UrK1VGj3jFebsQF/tJF
nJ6RnKCRMw2ksYx8dNupCtE227j52Hrc/FanCccLJ9Bs2E8IjRWt6e1S6MP/vbx5
IIwruyrABkD/wlsfaKvSnYl2WswCQ1cBGFNKyzrNPMGM1siYzRyyxmwIG86j8mtX
tvDIkgIpqBSjTe4h2hqXxCa70AKfao+TDB5BfexLWDZ7K5pZTU3ySo6Q/SGBisxp
m+eRju4lRVbX06oGQiThc1ceXvwQSasseKUd9lmdhzJmEMgiiBGzFHtL8X5n1Cb+
MGG0cvGKAYA/Z9pZBYcT1BoEr/NchFgMy+tE13wdJSOS+om4tlmWdx9KuLrb0ihb
IehLX5/Gr2v2MbwMVQgh9bEl92NF3Fixcvyy0gyw9wf4pNHYDteXEveO5JsdD1Ju
EEXKsbkMSuNvWAdyvcJf2fjkdnRGNpGmstRttTXhZiKQoO8IIdsrdzsmaNUOcywB
ci/E/lgIURn+Tqy0SVcQUCwZ+YDVkJT/eHZCYS29t3CEHeDtbM1Uph7Yg3/O1zNd
nqTYXqndLH8tijjdwh/8EucYE6EAIJrpWdS5SPnaQ8LWbrkRAbspaSLtFSoc1uup
HWx/anVynirMQL75VjB2MU7HEQtJ5XWFk3x2yB8DufBmNCD53kmocWeRWT+NLCCG
BMGlMeronaKfUmuJnz1up4BPDshqz8yxWdvfXG26zt1YW/+1Gc63W6GYExJjY31B
PrV/yCmwdF/f55i813zuvHBcEuJxdtPeo1fsvAz44b3hks7TUCBONSK5JB37qg/Z
a+9X9JxRuEosAA9X3m9KRNEjthGTltIp+PcNDbiPuWx0I5SUjMIY+ioIxsZXggbd
YAeEVjSLiDoDYVSBQdqJn64bB8YOiSeWYUcNXtvzN1NbyCE4kabWBdN4nbK9ljmx
S/uANTF2J/Xi7TtwlI2FwZBtip/V4zRPRQEqL62Keone5D0RMGojm0NwysJxQ2dr
P8opgGzaGfWr+qt/OVEOaG6HVGP5o8JRGZpRaAnpBxhbCRlgSvCGJY7SXdnx3Qhg
9LU0m9A9T+dbBcvjJ0K/HsfRjhpAN6b0o/4mqwVybqqaxIVOJSfhov9i/hRV1Kar
VQIWIFSr1GTqepvzEQn6U+9+84/dYFNpTuZprEEaL9P0JEbn4ym3H+pJntXtHTIV
hz8ybi3QbkH/RbfSnZkrovzm1/ftlFnGmDgSqvDpAevEaS/8RnjfAXDPBULxVn/o
veVqKoTctMi6i1m6mvsUqThyGTdZMBVXm9c6odZwNlvag7SwgLofqBnQCDcLpdi5
8PzfUbgIqpKRM3SpgGu8ldhA3YIcpWbkf2HoIUV2cVsg7RXIY+WeTACCXEuRr2i+
/Ojaik+eNHIgrzad1Hl38ISzl44FywHEyPxAgnxb6o7JRCaAUDxR2me3P7aHk7CC
wRLIms4QL2tyB+rLxV83Po+hwoBqH+YBC3VFYvwNawSFD7W6JZK8hxhFUVhMC7tt
8LvQbXClOflUECRtvBe1zu0cna+Hvswjep9LmgzE3r2dzCSW0WRIBZgY393/Hluf
8pwt3EY0NAkpOi6iAMQC5lsKtlio/G13Fc72Zs60kkdtGQfEBTyMu7mlA7wVxQ1I
voTGTqa+rhaoWQrDIDBFeO7VP1ETv9oVDAwNiUkiThMANFY9i6YR2uhNrNpvvXUE
0s1FpX036jjAnE/FQ+YAdVNFBxEiCWh4GNrbcPmWy7nV4e459b6c7OYOXxeS5ahD
VRyibk1BW4FJY9WTEAy76hVYvQJwW9WzkgIY62hrcKDGlKuTc/3tuVvnMCUTdOSG
npBbFPoHyHt2m8gVR/UVWEh4ljMsuZK9/xkww6utYHuYzdJsAI+RyJ2MK9uzRJ0K
KUs0qCEWBQHmfTeVhQBAYlYzU2H24lOszbfBfubHfHulsxa3FCyFsZ4jI6tJ3wcn
84Xbt/OxGdRWPM/y/TDoqQOdrgSYl7jZCBHE4g1j+B42JEkyO64ZcjEWMMK7JVCw
sWaF+f+u5GGyUXGq/ZgWg8NRpxLUUqHGAy5GIKchN/sGP0e//NvwMTBNwr2yu073
/zM0Vm5Kcqo3uiUD7tuy7tewwW5Lytj7CDeWi70BpZzRP1epxnkM/fopI6AY2j6O
JBSE5WaH16/2wD+veRDuwEkggVEiUSZszDuoV0z1iUih6QyKsTi4x14wydeGp8/m
g4jbRk4NCmCSs/U1INhNI/aTmrksg/5Icbujwxx8MJyULQgN2q5kxysyYzcF5KHL
YUhs4B05AWiNPg//LQSWPutEtQmb3DdR1sC6JHFnqLrzpIIo6Ecjjfzysvngtk71
F1xgXx1XifyAkMQOh2AbetcPLDPq/H64GmcuS3c5yt4uDdoU8hRNmnjHrJSwtq6r
c0z5udc23ZTe7GicgRQPRtCJK3Q2IcfhD9VwVpel9g3zhCqqtHq7VYkJbgWGImXw
+YwWDYdF+u87O14UjkePyYuC1Y0dr/OnvROV8nUcUk62YGDEqaeQxqxnbyUCukZC
Mh1k8EILcD2o5P7ZaK7yakmAeY7RkJCOuWLe7VPIY5HmJ6s0Lchomv8sfGyNaEZp
aVqNELuzbP2aITn/vBi50h9zjetceqUj3m+yOfsFThhGJlw5qbQB24dmRKmn1CBr
arSRE3WHeBlaK3OYYnu+7ecsCrKUzBe5Ykzs90fGi5u0q2jETjgL04lDjGgwB4AX
qKadrVFPIiY32oSGc7gqLEuRNgQd3PB7xWvFzolaKicIZLhESwH41pHYt0tI2lMC
FnC3J8hVHqv+skRh3Oi3Arhjs1LOEUOBHdV+FofKNzSu0uh+D+fcv7S2NMQoNXHg
xTRPzhDCWrB+Dx9KJeZKAeNmSSvCgPFxLc9N66W6jx4icdTT9+w4N5IBc7Jmuw9W
E20t2X75WruHB74UGGAnLS8O1VVpMft9mMGS22vBcqYxuuB0ycGKZ2QoITLHiwF9
0o3ecDrLcLRQds/cHV0F60gE5XX8ibEuZR1TolqlrEaN7k6anIv1a20EyBafFjPI
xn9BpyYQhiesUp6Bq63mj0lmTJSZxK7/mWHGq/tfKah3pyg3j5KghDVS+YKTSUnP
FKN24eHiLMoJvdDMrVKiIUnNnF85bp4b4njphkIlxDuZbYK4QfGa4qK6JPOFRowe
L9z1dGS0WTJucnkpItIxcUX1Y1hMDOqHVNfH3+FQTJwGlXoXiMTCSrGsEWbf07qg
xP12H8e5AYekcoDrtnjY63OxLhGXtQPwygHJ9q86uJbeO3DlswSviMAaDt5vX+Sc
dr/6QG+qo6gE8vn4Ji8KySB6EHgQ/hLf2NJFcxieNnizkotzPBuflE7wOgsICI8+
4H54715WoUCi6MmICQk4yvylUC5DYVUnhKEanoBj42OWzKTqCtGp96XxF6ahs2e+
ueqmty/7SyVM/J99ZBZJqfv5KElSgZ7eQEdJE3yVNiQ6/IlghDwlIfKvS+e/q/fV
8a+R/tOEAth0PLdEldqy35CsV5DnO2X2s1yhb4yBJeDsq945nkCzLsyAIIkQKal6
RO9e+1/PW92t132Z0LG/p9q81K8OTlBRdOeamrZufKJG5a+uYhY150Rl+I6gx2Y7
WkYDS7PymNSV1pkDDEKiwAbS5n1I2RCS0D6lECtLfgCnW4+fpuu6x0NzH+OEDLDw
GLaS0BmjOKZ0hrvAfev9AYAiymWOrWCOe2KBetBJ0hMUaVC9VMCTmVa6H4Gczfst
ZfvDr7Fm6O94Bh/xLX8VB76Pz0nEFgGe6steaGKO+WN63cVcLLD+ICG/MrO9hOO3
/A6Jl+K8oxpoPBXZDVvdfN81FNlAUdHKFdXAPbCNwPzdq0kchwqNA1ho+ub+/pNr
92gdsd5xUsGFVAGYAgAFtRzRIaQxWw4r7bXvqAS/ghC+JKch7kf54lc5+vlmT1Mg
Ecdc9eaLoro8sIjnU72DquAmLXhKQdMBdp0/061hOfZsU+H+XA3E/bsvOZ+D+izS
P7YZugup43YzlXBB/xpQXsdD5vIkz3nNcqrbptthYPpea53ugve6+c3GW528Em22
EDa7Muj6/syk6ENqXipF3AyegJvKImonsbKSFVQ/ENYUhvCSHObFqNEgSk1m5OYx
5Cm4IUFbMqLB0Oa6uSvdpZ37f8niVmiydlQ10lXFP+PmpXY9qK9ytDlri8dDFh4O
NQFJLovwfS9rkAZJ4pjilrxYOAxbV99H1SnzSHeVCmrHTMiZiyfUaLhMSVLsBbyj
frpc4xk/wQHJnKvvTMqL0yOS74A2Lp2E0WQoTYx1Bm9qyTop2yuJq3gmRFa0Vpn5
5cO0sJjBV0HcT/bi/N9iMQUK/BrdndI7cNuzmGOK0hsQ0tRBRgxN/O7omDGs2VSr
kN5LKjDSDvUe8D8ino2AN3LSSmNA2/EQhvS8/8rNyNKjZoXsuRc24UDXMrxnH0QN
1kMYrragBck5EiOyH8/73apz98Rgkqtl5C4x8pKh22es5Up/0KyZO/TBspI6Uu/1
zzGDz1r2vlP9gwPw2QZziBSu6AUvvRLKviU57be4mqna2RbzMHFHK/eDq7v1CUKz
PfdaNKzdqs/pS1nIH5ym0DYAQmKgz/mT/E6+vZBR8z06WuNTNAhxKiz1h8x/vugD
sYi55shyKRl0H7hULHB7lwduz8UOSRrxKlpIdiYqPyeHbNAH9ysI0sRUrtZ399uf
xQtYwZ/a5akAV+3slvm/GCfekuspgnKuwW44pYm4BkOHFQ0nJ0zYrt9OuUZf1/q7
OmDAd0RyBrYOIL6MsHaBmZr9NUcK/u9Lksgx9QkBo2lYYNvPGc2oCa+sDk/+4TLM
rOBVYJoDbnkeLRWuUpjru74hYtJOHyj0DBlBqvf23S+LqFwx5z+I+w8eMSQ08s/I
YyWwyBWMIMvWp9sQWLLug9SHZ3V9E/EKg9/dAarK8+nzX0TyNr5oA+R9aQ+QWj+n
OAc0GIg4JP+kPWNEEAopYOefCPPFft7DnJHhZMJfhOMoEJ4ZINF9HR68lcy7qrOB
9qagWBahxgrQnNqHhxfNIDfpTKLoxUbbYBiKkbbmk4cGM7mu3WUD8f/RCpe21ISF
yjtgnmJKWCARpMc8bX3z36ez/UnZKXmux1z7SAn5oQmFIZzpNeLEmpKekpXm0dqU
3C2V7ycKt2+kfWPpDMFjiJmD+t4nSEeCtO72khclQ0WckDS3Ed7kFScKMcoAJ95m
adBCVkvtuCjk5Nbxk7ZNF1ZnOwAfA5OLZilspZvUXxhqhz2lEmkTgUh1Aylqq3MT
pzwMPLjVHShIazD5zij66fw0qg3cBG+SKcaFZZ7OWwTpB7DtaRyKDlIU7NdKgfAg
GEVNREnVorjrIOrwetp5NtWQvlcO0A4TAYOgE5ueW337R6IR0xkpSNjEZuX+G0oR
IJrio4T3NssQ1++nSA64y1/LOsbvIAObNvxijsRvvEkV1tnU9V3lBnwqLApurdUI
nR4q8V22fhoAeQj0Fsb/E+Od3zx/w99EEkWy2CUG+qtF5otcT3Nk3kNzzattIQbJ
4YiBN4xRAsU9cQBEz16XgCRy+6xVBF+jbcr0/yomVnDfaXAm7ghqBX78fVO81Yzb
ZGVx5Wd5DXhwSkZ4mxjnrblhWs/1Zs3FSm82jhIuJ2gLqWp4Plpnh8O4ElV8pEXB
8TgTzJG5skee4uJcvJPOmINoeBkSFq31YFLxmDOKr7+4FrkRuzddGnJOXFsjzxqa
X0IzTRO0DJl8ZpuC/gN4ykCghxJ3UHSnIx8cUttF4ry6OlU2EvAk2NF6BWpwayde
WrVe+V6M90fQKXXhbhRzLGm2K3iLDQkEii90u878Vc5gBygmckqU4W+9ycErD38o
39XDXTSSncVpPTGyP0VN/zQKmx9nzKxapjtUEhnReYCnIcLO36TysBPGHysdokeC
4PWaMIJWZr+6I4I38/0Mk5u28yWxpCFlWEXJrjr7niDbxB9y7GKb8WvlFgHCEo0V
F6o2L6SL/Tpjx+wpN6Q74RU8mjKIGQEy2aqtn7Mwb43cxAH5bFtRtffj+rmu4NlD
yUugO8dqTe0hWeUQHzf227j8n0lgKFPjWOm+cx1R9pOS4aC1f/wKqolVqgHF9PCp
mvgpt7ebD6zaiooKV4Pshes2hah58lKVKdjaV5TCIX61FlRu/MqKDmsOC37M9fXF
dKwSctO5cOfBR3+UCFTnghTSNSzZoHfYpJjupGxVeSLDkygQ3wwl4sc36mPh5uMa
kXM2/zp57hDgtVZ9YhaR1eN55khzs7QGFxz0shWcPJXfjcKdqQp9G1c17k/3lPOq
dG2iyOMX2FpXkZ8BfDl6IGgMRunTOEfdmqo6Ma0Vd6IXouj6zqQj2JVHyM4u1TQA
o0lZumJDjrJ1zp+XRDd1oAA88DP11ndzrmcEs2QMoQSHZk28rqFZJrPiE8a787Jn
x5dUKaynFSeBBgIy6j/Xu49XSESMeLll5vXmhkXqwdgruNzTYYtL67/4mwdraxL8
+0CrNu2d4+oXxydlvcg6XnwtX570RYDBhXXoDIsLgtCBko8iWo1SymDU/3T649tO
QF+fXOQQKAAIksxto7YVVYYoAPp1NHXSC2E0lDV1mqXBXMnKwkAzvD8LaF8wgJ/1
FLsdzCF+YfCNlgkcSgxR/N4mjEEsEDSt5p7ea8OCqvo9UmeOebEuzNZj3oJ8q67p
zH9wnTnDse4leKWr0Mnn9UfZZI1ajYlMXKHYu09rQ2w4sGfM0Z8800l30d6l0fOb
j1IvhcCeSUTuegCg3HSGiXWZq1SAdJAg13uaAC4MWq+bOofz6Ytt/fiW0qsHxweg
xr5mz8KLDK5uhCFNTxmNgEwA/ACWzOxhUsVhWnZekWBRhdurKz4BPCtqClWeIoAV
jmWjRCw46FTW0YHpwdIuU3S1pFPVgXNl9MOMRNa1NZOrumRNkM6qJkSZmYJubKxL
bHpJtpq+JrVXxMxr2+Um9jJx0OP3hlCSOU8tnclup8+Vueuz8GnSQ0LaA/8M2aCq
4ITJ6gv1ulrpELptWm/JHp+N6aqDNuvSD5qJcw04/UIkjujX1GW1SXufiZ6igP02
mcmkjE5e66Yt3fvrojC8/IjIfUktf2J3ZAglW3WLa0BHsQy7mshhwsUVT5FCe7Ra
501FyhsJDCU831pC4KmTZ/NQrzSf/LP9rJrVfCi2FMSN1788I1uTEWxs57KFm1WO
XcfruVKdeNnoVNUI34+rCTZ/D6inUceBeSwrD+PXIKMxDL6Gk9JQlZgPyoJ39VSq
oGmj9k0ntYXcepxu2v4nVEOOBH09rvSYtIC+8k+CoIzBre6/dcziU3fcuQ6ATO+C
h28/Wu4w546C6G+GuO+93tmYXRKaWER/ajQ0/Niuj+t4gZUxQQq6gqku6WYRzgze
/A3kL8iMUp+/dQSY1e7BwWggUUyyp0Lum/S5Y5mAJ0a9mbY7Mc0M+CtO344xpESu
T77q5aVuj9SsIQfyEm58/5ZLJYWuPVVLDkQabn1HPBIqtszl+cxFI3dmFsYkjhyb
DQNs+Xc5+yZTcZu9G7bPbku1GlsA0jWVR/6izjjZdYP02N8NOOkEgDNFzGAubgx+
92R6xpkcpUYw2YyPFgRjrRU5c7UtBSkVViNz3SBOIv/k3yl1oIsbq8dKh7NPJhPn
2XNawSR5KcjBdGlPEWv5G3tC8rhHsoP26pLZTYst8ZyVvXNHEU8dxjCeT5MLbo3p
f76yrr0ultud0/lx3uLEfexzt5Cz/rnrY6gfC+BokfqYV0xOP5Ora3HWfMmnsjNx
dOWwYtL5wp51bjcunLhikL7JBl2VueebANV6qNkjgtHdXfr3dZCxsx2S80CaAM/U
leidy+bY1HaToxJAim3sXhmDoSvkfstlhdTLeemVMHXcFIdhlFpIWR4TCl4TpHOh
54OFV5+1bWYeSzdyimIM8+w/p+tTd/esafpYaRTFFhpx41O2OBwJL+xxnM09GCjM
WwofCFoBNww2S79fdiG+s8Ayhv7vDbruvx7Lds8Olg4pnk+rtRvl2ywRu/QOzHiX
CpgUV3M981DoxgzwANoqxTtpm4GiiJ74qdK9Nr5g8SPYpHZqgRKV6ayZqKhgsHdx
nYxxTOTForcSW3ZrkUOv2FBt6Vt5dI634Sq/+sh7vksxtkLoP2d0ZrWJ8Ma1oOpo
pWn387Vpp29jz0vbn4EnYo9WTViB1Pd005fU3707Ifs22GtJIFWlsO7z/YmJyTus
T8CW3NXCMkyq/fXtp5WJu0+9NdrOREYim6NuCfpSvC+vb9Pzrp0uwqcjxzKNHx8r
R3L+X+YPy414AOOnrl3K5fBPzHubpLGUVtMziaN/UpjLmZUET2dO1TWcohrs/LSo
bkxwGleW7LVYEPX5snp6EXBEXourPFCjCLJQ83Qv5WalqyifTFnoYDb8RgQ1zXFL
j/DXZinGJMmy00NFf2O1m0LjxDexYqKV+SuZC42x48YVgH+Vvc5ExrURwIgphvzh
/gx8g5nf3ufP6XuLUQzms897i4Q9+Rnam7B5zBc34NSrLEBp0bCiMGj9gyiBIiNK
cOIObZKeyyHukN5S0n3olKzE5++2aZWlvFCcsMl2aQsLKA1PmfHDqE8pW1ertu9F
nl3OGNKKxgSMO1B9uKVk/ZKf/f9FZ2Rd9W7JROqW/NAsAy/7ysksu6gJy3PwuGAi
+HPF1sTVrnAkU6+hjWD9GdrmqXfMVsUB+XN9OBPSxx6/OS8saQ0A07UfdNabII7W
ks+fSj7KZZd7bBAvZcNM6SOoTK49ZkumkIxRDM+ZTh3ZBAj0s/xKKtDOWuHuuUbm
9Xz1t2wFE4vaLuQe9mSTJRi+oBftGllig0GOkiaTy1mRUTP1OlMg1T7qV54RbPed
IhSY4D3akUkUSsN87EX25tkbkPp8FgiQxFN7AYStWvg5QeL+k50rYkRUYuEcgKVh
9XT/mqlmn6rouzxdl1hqKhCwk60nnaq5hBzAgMSIaCHXCAm8Krv2vKQU8f6Mu3wO
2ofVZi4ePig6SJhLhSYNGsFr1CSAY0fT9qNC1hS18AFhkalX7U8yh08coPaUOuUk
XHPs5j9zdYSoWFAUirxYJJuVGveuuWP3VzZougt3wcVurMonXkOMOwf0+hjctlv4
tR3nQK47CBa+/d/e405QMTjI9Wac8wwHdjHKFj0sv3MhxebAetwjkirPURwJEnx4
xrvlR17uwdq7ByzeKKKa2ZzfHbJoR3084/8Qq3wjC0ORQNnyIx0LmrKm9epkThzy
3ju8QMAp8r8Ed4PttY1O+FY7i98EojL3dhPmt91ugV3Jc41YMaVOZh0vlAtMJ/wF
MEWk1qQv4vofNvNSAjh7EZNxxPXLKXzVOLzr2jh6QQG6y14ljvZR+YHND0fv43d8
/yWfobMCWq9IWX25upaXGhCyV4P3DT/ttYQjkgnuDiABtUTGGKiddhTl9oXfLNHc
p7Q8aGSINywpH3Vxx7S4s6hgOhSwB70E9D3cGdt694ibHWCyuZQ9zQR4nSeMhr+E
JNcsQ/f1txBGA43kqUWUARAbQaLYDbIxlfWiA2PUXgN1PDOEVFQZ8LouvZLsX2m3
G8URqMU9YwMHTriqLfmu8tOlWkHJki8qXIE8DRvrRCXHO1BkwV/Gj7PLGjWWS+2q
OVVfWw/6xP/bpGYY4ASqW+5brvum82lLRH7oBozJ/0aZVeJpw70TvB4WKyH3FGAk
r7mbOSfJUB2EaNRcme+ieGpa34szvb+nBBkIhEfP9O0iHDHpZFUC37lOUgSkInI0
SmARmyxm4ImjEEgeNeNrHZRE1cLn2Zhzck44qDU2yjTpLHQpJ2PQHtfwSI51fDYU
FURxFJaZPip6YcUwfkIBitRNFgOpUurhLoB4BHaBdGCM6cyVVGQP/uc7pjiVJmR5
f2qEiENMmPoRGXFZY71CNKJHLxBl/69dSWF52Q5nqAtaO5+XLzLrY25mKTMhooe1
9C4BZceOSOE88kVhdAxtCHF9NgXkpN4+JZLXx4Tw5MYmXsa5LsolExg0xpYjJK0l
L3VTBCmE1KiNwB8LeR8S9bdFWRKZYA04Tcd0/F7dtlW0dwIB8AjQH0wtwux/3way
Y0m6/v9AhYrSvh6Mlucby4FP94JA9eUggrcXutEfr3yunn7tx3E0r/2PPJ/osvUO
vCZHAZBlLBFvbjQVBd7zgBrfTodqVZS9uBHbjVedkyCAHt/DtSVlp2BcQPNihgGd
jons3H0yNVl0mgr2oTBvAmOTVTCYRC5fCa77fC767O3nkCk9G9UuMookOz7Q+pTB
WMDJcHyD0d+YSJKZzdWy7VGM6z2cZAMjHvP3hBPEeTXkW1bfgoS2D8Hkca+bczjD
1CmQLq672UiCyw0bobkF2QeqROqaoPwH+jGuupew9kaNsF2bil2VKtDU3a02SDh+
iPNHPyUpDjkbwIklOm0L6jt+46Q+vx+v+fYmk0u4rLuIiLMdSZsppsrXZebgNw+Q
FGyd45ZQbq8lL9FOig+BoH6F0sxZ76w6SWZAunA6GjVRHHY/2JKC7u3crDiTnplv
r3Vb5IGzjGV7ZQVnvqWmFIb0WF0srxVxL02h2Vk6bg2SRGtRsjs3rwgUGqytNzoH
C2yh49w1kARqRL/9se8fAqCzoEKKHpa378ojtp+V/L1xTp6zmFhLrfABgLtdWZFJ
aE/z219NRZgeulcDWWbUlev55MGn24W96GbnJI6YePMOXd1M+d4BslbhXJh8ieZ5
KhxQ+Ie9V1bdU5GiFfvTWnLQ2HLJMD9VyX7SneXuWW/WBetuuv4Rd9AyiK93hp1u
WXQ4ZEPtvZTXRv4fF8CsOSzM5JD/nNgj3zRpW8+bJT+oTxfEVuDq0/Deuq35C+wd
diOUNkm9akFoofDEXBCfmff5O10HBbur1SqlBPSwTZ3XQINFGRz50b1EKbIIwiHl
3lMGYK2WsRuURqpQ9nUcr68fpy8pdhVixd8jdMgf6Q7hNsckkTqd3d2blIPcTD1b
ndzCBe4f6acpHD5CMWULfVscLhg0SQqd7dMRQwjKznfhcqtAwjFsq2C5KfJC8YYe
15nP8y5Ezh9CgwNUV+BAlb4WRc+2LyBdHzj2E6feumiRR96xGxlAzdQEdqdxkBUv
MjLOZY/XrC66F5UTv3cP61I90dzLVk0NiPaHLoDlS5ykB1MfvcTPY4Gibas5LMhf
/fHQgExxpBJk2Ryx0ZDy+Ntpk5JuAEE6WkEfDnjnpO639u1+1sZ3twUDs2WJzuEL
vxa6qJQ1jtZMeRDKEz0i71d3lYDP4aJy48nFl+h9qlu+AWDTTQyRFBJlPcHdXHgT
nncG66eXBWfxe8CrU/xvsjaxRzOF6yMk4S0lMPgue6LqpxxnDBjIIlZRjqjABB8G
u6Qm27EZRHAGr8IWA9WQIKQ0JGLCQ6oIQEVdT0T7zvDJJ6CcG5rUuB7V84qhNBaO
CUJlQRAh7749C/Nhrl7Oan/UytNP2X5UMn2fXRBp3nt1xwsCMfZ35To4WcXbb+oq
9pTUxZsgjiuKZU2jMJQybbIHhIHbFRCf0vKp9XIgwyYGYt08IlUW/Q06iSP4ZwBt
5BC0KaOnTgBbM+MPEgWL2TLIyaA/mb9lrsbLqW74LXt6iCXlMcxAK6pQEBC0Vp3r
2CMlw/6jFNfzWOmoK7mWDTTvvxtq1PIHYPF0lrAkS34DJYMP32XwIdOI0HNedXfG
QiNmm4RXeESrnsL/Sipmf6n35vbcf7Q9CtFU6VhLrwg51mQbGDaC9igWa1g7Etkr
mtNRDA2mh3j2i+3d6DT3IGbUDg4LNfz2hERWWAggxyjLhjiHyU4IBO0KsdkLh7eC
ErWVvO6KoawVGJJoVLQ2C7VwASP35N89SAJDfxZg+r/zWL/RdbYteMDOEEbgf/Oc
PEIn70G7S0+JeI30WR0F5EXpbONPybSxqN7FCGOjAhKxsDPuVYz5Br4sylpzk4yA
UknJegntv4cVT1eV/8EAIKycbqjbwQnNa72uteQPDV20ERBeYPuP5VmlENVXbXim
xe4c9hXG9R2n86WwvjCQtbOBnGM2F+qtFtI4JYTw3E+SiDae4eGFnuYG6PyIt/Il
TZMZM/1GzOftuPPeHWG3OXQyzDLl5dqvsTp374raAlCW/lXULJAY9S8hgk8Or7Tn
oNX4StTZL0GluTrVBXxfr7VjmUeeRvVLipa7lW4pAo1eXLrDl5Kc4lhB8KyBRgCz
dItE7NdXd8+MekP6EeK9rlVfQbI31BY94i3+aTKuIpuLR01bFzEBPuknzgVifB/N
oOVm5elSrgCFUB1LQ7I93Q0mwL8rWGBBA9DLfAPQq2YJPcXLJeKZq1bKdYUZzuZd
0s2ZqZW4l3tjA8VbXDAb6FQXlH3ym2QSpcq+hMZTMXtDZhqiQbV6th7OhvXUDPyp
avv6Aszpw9NYGcLIV9nfOHuNU7Zfrk+S31I5m2h1ubw6nIbW0ZvQlckP2UXzgfFi
j2i/cDhz8yZ0lBdMfEOh+zBLjMUI8axvQbgWlln0DWDCiNcoYNRdzBu2I3EM8k4I
P1MONSs0KvjpbFgoCpxUn/+6teMERZa4uMBG1t5KxMFv2i4q+OtfEQm8AMEQhJAA
HEd5crDXyhagCMkOTf6yFeL2s8sgw+0qbMSWSpDOq/mmpqj4TnJBdhsDn27XmkQt
01vTlY889C/iVpWyDt7/bLV/2i2wjJHPP71ZkrJH7d+D/3kCdtW+4Z86liCQxiAA
vCkjtuRpVTyCu8z1EeAD7rc+jG5qXJR8zqfs8BoNm390qbZGaygtYW++P1sNYJlP
9g2aicMghP0R3eNr/bE5koSROBmgYxoPV5+PqbHkhWXzUzxvSpcXnMhqYE3FS9Ij
Hyk2lgJ+U0idsozewPORKh6Q/mI4XJvcadlMwyV5Egr8pfd1ZrTzltoA5KWQ7TGv
3uiGCf3z4IpIRUY5Zs6en7I4vYa5AtB6zkZjkc/4Nf7jOLIQyQucnIHtyJDehDrJ
96i2nhG1y35yat2hqROuTAUNX/FtP+4Ht6fb1fmjTR1+Vu+eStkXFelKhl2G5pAm
CXESS3Y1Ho7mJ/Bx1n90emmSZvuRxAC8vWATHUaqSKldVFYt3sUe4cLVrXNyyyoN
vRfo1HUW6rQsLatY5pMSGuntuXnqp66Rqs79nOHcHVfis4D3UTiOa3MupOeq9oVj
fyWwVw/n6BTaYcxUIeWpnd9Et/qyGpAEq654ipy7WdsoWKlu6/fSvn9qf5cS90WD
y/v4W3cuVqUFhR4mbRCfD21+oYKuWerB3XJp2f4++Q0l5mVlXVnmVjHDWc0SYvxr
j1dlG58xNbeKdia97jDaP/AKmuPK3uMfcbAqWNGacRkb/VWXW2a7r/BjRtjyCBu7
E62FAGg5PZwQ8hFXXvD1zp8nK/01nomZvuMuEbW1eN6BCfDFcckU2elT6cblmPRu
EyYkd9190D/ZmVrjAukR03j0QvElGThPD5xoM0XbLiASJQ8eEAYXP11bTNFwt7ps
L583TTUa5nFkFNlZa4ko2qGINNcDSGb2+jLJ/uNz7I9Fd/kFA9VCDYSXm8rMwxtm
IUu6xNj69vwZ/IpUUk9HWYyA+KdytBDxnm3uBgAZRdCKXk2bl/E52NQAzy5Tqgeq
doOs8BZrZ64XJ6I7XMzJRGlRKzOrVWTa+Uch3aZDvk0wXMCIxqzRmcIVoAynsWtR
qXYQflZ96ujzNlU3SQK7OKsWSRGXuY/Oznu/QRe/5031VerJmuAqfUzVLulzH7NN
CmNdS4x1Ux4LtZ/jh8bkWav8QLsrWXEPCXPERQrhXg6sCDYIl7hvlFLPCOXi5zbA
Mzy2MbsxkG8f+MitHo94pPzS1Nl8yYqoNIxKKnh/iEvU6yqjRK1VIx5K+RHKgzr+
wF6RgSbWU/qLtjJ8a61AiYY2U8Fh0zs8CTNuEn1tI6voiEQgJIkDOAZRDd3MnGKG
+r5q0A4SBCoN49GKmlonoHtVY8c36iwcMJam/nNqpIGXBPQZYrFdQoKOnR7B3+nP
zW7xFR9O8WpFdZKjlZLDwkEcspaQqsbOq1ehFEZthWcbHic08GjR/QemUkvfMIiT
Om+0URd7NwXPIULvga0YHkkd1iMAhlhzW5fduwPyXjuSoGqWrVJisWhTuo4vmfZt
J5IDEzyVasZLGSLsxhhhw06yCylPAdNhykDIWPCtEgmw7Fb3/jZnEID1UmkTVE34
WYwq6FJayiL7pNDdkweUCq6ISCqXFtI/eQW2JnQ+kII4mqYhH/eIv5Cd+73/4ksI
Wi1tAHAiEhxsvJnc/7Ag5pQ0Jf2mHIavjO22dR+qSV+8IzRXrgrWNbvPi+u2gY8u
SFq8TiQC1NCyrLyK8/EsVDYmEMBmmdWhDmIFiAGHrOQjh1qISH3csmR/KfYxjZG/
KTAn2MHDMsTdXAWZcyZj5a3NmybxoQRuHr0lw0mTqhBYA4zVgYRfrsaF3ttzhvF8
UquuE89Gu0fgu8CobKBSYI+idII/vprZTPVnGT5jW7ny02NOpigvxGpjxw3WUiKm
RdF7HYlP3OsDCpDFi5MECLS+wY9e7u0tGo1QNLZZhTyoxDZDU0cGIXVaxe36KvK9
e4SBY5MYFRspRq8ikeLma0OrR9hPIHRQiB7b0/KhLAN6zcPwXcTa5NlhK7LB25FW
DVJ815m+L7AqRAvC6iCxq1RneoqOnCuXIVBS1E6haKF3gaCykJTQPibrHKZ72IFv
LXNUzcrwYpW+pgOfEkFynMA47IPc/MthBljh6a+v+R61FeaIzl3dDdvSHBUNFyEE
w36KkZlzfy4USOSyNcnDOT2nJ4stMiBh10NRxvc3+QsoN6KsYjwjbJGaGv49KhJp
G+scl6udjVBPAtwC3KWbIQDmTn1sLh9VvJLIAjPbZCQQKZGUnLqrOR4adQ5TOU1X
dvryAHlLpJZPBOQk8wTnj+DCy26pLdscavfqE19TzJHchMlsd/19UrIla90uepbV
YwvFR09KrrIviL5L+yDYp56dkBWs28ICoayoglBA60g4cQ2mmKfSt7SxlWujHDnK
a/UdarcAlX3y3vJqXTuHgywvrjiOFdgaEugM6DJTdL1gr+Q4LKAwrdy5/6naKaUV
0tBK1vwGuDaBECdVOrJLrUxGvhz7gu7KcciM26G235YIHoEHPq9LpO05f0FEX/3J
Akc3YFN+RbmvDBnurUI2KNmNB7DYizYhypaf7owbW2HTSSyUi2ALBZy67Fy2gwzO
N1c5HZ+pvFvJlJkLvtlm/ERDCFYMM222gutWjmajGplAnB3B2imZBMNoEMND1Qnn
qmlNhXgt6/Y1OT1viw3RQk0Na72czbZhdKZy7gADiBBo8MJu/pYqfAcg4rexglty
SCIDy3Vjpx8qxRgYuuCO1z9//WFvfrGiSGl5azpJycK5Nr2gaNC6fKeoBr0oCBVu
bWlTGJoiYGRKzpYQm5OKF0urIH/WKA0j3APRXWTvt6RiCBramA2/rzwGCrm3fl6X
13mf+Qkr6OMDD1pOJCEH71D0YDSOv1CVqDhY2FfALfV4BxfCRQSWf/ozFuBiBf/V
+6HDfFM1dWoThhYLMfGlo+bBxqbhK5RQ/IqcvrNK5BLESpfvE+2Ynwc4EdHEcdKA
SbU/OinwGlCSLBM/VvlpR3VEdaiRFf7YioBwYPmUgyknixKpYQD8uhf2V8vAMutm
hnw7R/AFfWQ4oPQPeMwRlJSj+nSf0tCTS4EJza105e2aq/bSrr9GoE2xBdl/g+HS
hupvOYvXhWfe6D4UTLu8Uv53efMbZHvAQAuKKtcRhtrSfJMq4v3sgVpXNy2fWrLI
J9+DbLDGPJ3IrdVA9jDMbaXe65Gbom6XB52zE4v3N47hzCe6W3jKJYLm/GBLkJaz
uogzzQnGx1afUk1QdHg655loZ6AizE0SzxtqnLst5UKB3xzUCM9T8Xp3y7h1miVY
u02zpeIcq9eNiPvAWDZknF/JpCoeOBbHRSQB6FTZsBsNH8Cg5rsL1wV8PwENVjId
kW7O/VIZKu9ajKiTLmHhhvOw0ACDcbSr2TwxzjQ0Cny7QA5jSh+7BQUYrlYZzf0B
GyG6rRLG8XOU2YoIK2DGYOaLPqWXQg9C8LeKMAmWxsI2Yt9RvzAE5Oz3t7Qw3LRy
NyWYnrcJ6J/TJlo0Wm7stc7LZx0qTe59Yoha53sBl4L+wz5wdmgS/YD2XusycIsa
QgzzfLA+muDyT8JGkN4UuQ3R65u2fTsuUH3GJs6lWR43Q1pXDY4PXSBgKKmFC3yE
y4XveoRuzFy2l/YCzaalK1zBx5yBHo6CMBvBR6QZ71v4jdiJwzqF3w/FevoeuSKR
Nsw1l4X5yW9YOXsLBmNrxADdNsAXlLU1rVUfXpgY+roB2uAzIIEvhfcc1AEfuAGa
xHzkypiwZl6Jf20jhik++pQzelBw2iQHgGF9D3PwA+u+k1YS77tj3wTciWl3twmO
DGMJrXZdPYgsLR4x3W+cp6kj0zg/9rjbcStJqxA2Gje/BJ/XDKF8EMycqWydC0bu
kVq48kr7t6cGh9fGw5juCuzRJQTlrODWB7CzLDXCytR3b8kBWDPtVT4SuR+InoaQ
KK6tzMdbVBvNoPj2U4n+6zx0HLBlN0mhBlQSZW4UL9oZvfcyZfr0jlhYFCyK9ufv
8lkaIFozjxV7z57u6gQomk8PFdJrWuCOnVrNkvrd4F64ETFlgICIc/qoZeDO/TXP
l8y1RoPn2AJZc3RGKxmdiOQ3Ks+XMMr3ACYzSQ2x+1eXF6XWL5xMySbfcFnpFlrU
DP32abl0cSKxq512YohloWpdCYEn+ajQwfbMDiXOOkekRD1bE0qUFumbTKr0SwiW
tcTfYAXAYzGNlYR8+tAaLLWtfG8awzsdWpKp2z4Z9g0M+qefHHp5bDU3XVogER7p
vDHKSDaQnSIC12STPCSV8gEhJMqpxPZdtKNkQkFRVY0xW5A4w/6gKM6XGy2krKmB
DFFxqH55yCpL0K33khJDIvKU7DIcOj3pZau6dM/veCQoWGncIzh4YnQTIiLPtrLk
FyNSsEF72Gn206heh6pYMOVMATtIfuGC0vWbdalsuyahbR/ZPmm5Tc308vAmvSkm
Q4jE6KcZYi34xlo5sU+nz1CA2cTFvsqSQjQkYYum7ihC9R+oubN0GK2htbDHHRs4
IiMwj7fxMkvqPM3N+slN/NSWbyY0iUxQyrO7Rp2Ip+6ysjACFSbJf54OL+s8qayA
Ad9RVzzULwxqUEqvhqKpgdjM4dzP0LTmiqYOtbs0ejsRWCgnUK6a6mr02Jmv8ESf
NlU7ThKE77bN5ckbFGN8veuU+Zt6yqsVQaHj8RO9FqiP+9WZ3HO9F2/NVIlq6x3y
z2W6hpnp3Umqu6Bn4gYmgvKoyDjWn/jfx5qXG/ZbY5EMnznjGLDrOGbCp8oAGZBS
4g53Mynm7l8gB+fUC7NXKP6ru2HcpP36oDjA+mIZMMN1SGzmXYDcpa60O3OQiK/a
0UST5aNY5pJqAina5U+0vLWoJR5R4sF+VktV/SF/yL4eJdFWHnItkGMDfBu5u/MU
RsKNUbpR6SjpbXbyFVwgUjU+VaV7qkTO/kia9/Im3kUE0MutE0vMsdyvLVZVUHf3
VD9Z0IINTsZXoV+pOgimkt09937U8cE0BJ3FeWu/DCBBB1DSaSaxxJZnEGQPkgF1
sjYO82Nn3ViTlh5OLyA0EHo7PsnU57f7FQjt1FU+C3hpEXwPbfoJuCsDhFXLBaw+
/XzKHdzRBEAf/KzLTOrLIiYwG8MRw4ZE14OcuRsC+OxvB/7pvdB32oueyOpqkiL+
ga4+gNMzX0rexy84pfj5YZ4ljiH8F+P2ZPvKCsXKJ8cLEjwROo637prqm3dZ9Jbd
8pwHOkEAgy9soK4UA1lqPDKkuLsVygOHgrcfLQPbL9WJrBo64ozZRjbYRZk3uexL
z8N/Wq8n+u885TnQrsNIoC3E4amKx/BE+cyisBNVnQY6iCaC9vK2qSXZI8MWpvP9
9lvLeE2auOmycQ1vJdDZRyJJoe3B72DWUTA5WUpyFO9/58ah7oisSKDLarFC+VTf
TUZN2x6uiuvQZaZ7UBa133ksFUfjMcIwjxCHUZLCRWh5TcictCy8g85wQL+n2bN8
oq+nL18873zt8j5Yv8zHVKF/ZKSL0Mscd9UC70lJDNjlwz2aKw21HzBaQ0ycTYpw
FhGj20zEJonPfeW5vlxDyapJa792nw5BEf0MTduo8pvKv1H6H7zTaeP1ncKYSaqI
8A+RxDzO4h78VzrAWr15e1iQnuUqRwlQqAjMqv3x9LXMToGnqMP8Fmt/DbwgjCpn
1XMqu271AtJ/PC3yZPWY8yjtnGCL8pm9DIx8hhz5LMgrUuB0LBN+L2xXjRfzlhhF
XhjMou9b/XHBqKrZdO7sVSSglpxDm+QvBVknpjoLwSlTpO6OE7+lV6XXcFVJoVSh
8E8WiB1u+BfV9Yu9JuGmY8oJrvWjQllHuIaZA9xTTlgnoZHJxggwpcS0AcIrwIMs
vC+6mwl3PFHgCXk3VU2SYcCO3LvOc6lRvCWIKWR/Rsnn3pekWaRk3iAeSEPWny9x
FZfIc9OC1wVFqz8Rmj0AOXavyWznU3VpanSn9ydgYHVYkRHJfFc29Bo6whfKYKIl
t8vEvhn0Ug0E/fG47uFLzKa1vKCGyS9PjG2pcmGhOYWxhW8383txGSXUQhcR0R5N
5wr60LuqYts/buLTD3iyZWrswWfRxTGjRqEM+hDTiKN+9IDBMnKfoBigrNHYG7MM
ynYyfFPjdfA7RIRIyrG5tfOgzJJ2/KXDMGlhaD9VkGVyLLfD6JEiDQMIygvGNgsY
UvEwrbTKGquz87RBNGkl5PL+kN4u1B+FDadDCkRjNENlQKvvb3RT0IOe9En1yTL0
3TInK8djoIhQ+GDiAzo9C+seW0BBzLVejzb76cG8rq0Etxo3fghFnKTLvuLzn0ev
qQjXislGC5nks9zKlk/l55IBXkRJo39J7RNRzADGwgpF4KPVNdP6vEKhepSNXdX/
cYxiUhNzuOhPI/jlZcttQBA+cWSJXwVdsztJpGlVCojHHttRpaIAhyZ1LGp5/4oa
4QZe3MMctXjI90SZAoSD2RgVuPM1+w8+8SNbpkSqgsLGz0dZLYG6tknunN1kElOx
aGBqpuOul434lgAEpj3aoWWeOG+FNd0C42kN4OBdJnMk4wbg8WDJ+iLT66xivjjU
vJm4cJMAkvrRszFlHrjxnz4aRoWtUzlum2OQK5m6VhOCPL01trIeILapKc5E8xpE
mr+wUiH05ODghlCyj3ODI7UeE6gwI/n95AoMtZy0awHerbdCCRHU+SvbZi0G7Mpx
sNtjW/GTMeLRV+Rzbgoh6WwhBvhBQs9nAROudRIvz3eW6P1De/fFFYENsW/g/f44
X2krvQRjBrEI4OdfMLo/yJ2MkQfYrDmg7fAR4I2V5Xf057hOVvIHZjH5GyltsA/X
atd5+4KFCPCPLv9T96WV7ybYnvwp3LeCYBoO2UXRKm9xHUA0R1CNbdq9Y/3oFnuO
mBq/OLSGW4zPHeoS8sWiVNRDvEa3n3G6PMnRIhskl2tS0NfrLMZoRF4jdBi98j8q
3r0cXvQE1Y6OjKIMUYpKYOrSaN3ODSbbqnp9PZZQtsNtpDPxWUSMQ/+FxIUwv268
BImituJdRynTER2dn2+5STZGipQ/Dean+Ah5Rakzy3BjEURdHtBTM116gm0Wdh87
A2TlabNw9t0tfVlg+LnXDpU9IG0XWmeZBw2WHGkKc39nMfyWQDPK2/OmcBvxcsBF
sYSuXw93oMNLaicm9gLfjkGUth6FE456Lb+iYQtXdEfn3k7K0iGjYOL+w6thrIaM
AMIaHfXWjZEkCoz1wg8W5amH3f/selACk0TFNP7i0SwZeuJA/FvDjiS3/VfQ/D5P
OjewRGvswLBbHvGW+/z6pjPqKW6wcUVYiMbc6u9URSpsxGOp/bwYuQk1iApCdktR
EiWIPnoq0UmUQOI7WZ91BanatLc/elfqhT5CGd0xD8/XvGjW8RvIz2NGB/YiYlnB
droexgTowYTJfQScMEI1SH3V2+Dg9w3lwpsumyMGRNXFcAPo+sZgE8nd7ks8zr0w
niAdGY68yQWmDXuBkXG36aznA09ueRvoofDRiZjKLoF07Y1tIINgo+FzPs8NDOU5
3jnVkQFM5KqovC+PLtmLFELKXdRnpI9dkrHMhvqSYyDdDR2qRdlVA2BFP3Id/eKZ
vlEn2/9IQ+6qAG6k2FMAevwVYefXh9qhKm0JSx3/H8H61Hxn0SY+OAPhbSXTnZg5
PUZVmSFaA+wbuZL4xfQ1oLhtrHp51iKfzh0Uu7WreP5V1V2mVX/5YEA1UGHvzcZ5
0cdY2z988vcbglmLIXZQGUemxp4IFZyPYvehCoEjNSRynjRyavearnbGPwkdfZrU
MXYYukUhnj5GHI5DaZ+DQRsP/vBl0677bhfjC0JlBEbkLDXJ0zUtZbkKOGo0IyXZ
Kk2SnETE8iBsOnRnYaoNjUUVyirZtF6yV5A1W6iDn6NYeMyVn2/dC7HcGTEMDI/P
pOkhbFPsISgT2yL1IaT+OiCYXtscPGisN4Al6YRKuF73f9BrFgUlNB7Ej0qvuXSc
dddWMYrVqEJtmbX9ZVMJlYk5Ep7oQimb+qKKzz2LJDZZd1XbDPYld5BKUtYAcQeZ
vHax6+FPSG7Pz2/olyGFP9HG84FKEi3VufkD4W7BwlrirR75o3YcEkVFAdRbX/mK
sHLBEygfYafjILzxIOFR70F7i5FRvlaEYljNPNTHX6K2MneSTGCvqt56bP51oqQP
UanKwP95naQhc35hhdJecD1947ygDqXvCr9RJeR/DD1YG2e2W4PqL7tE9w0cfpVh
V5wJ0DH3q4dlUmVGrMseZ+XBeY7b95JcU/7B1O/apkrN96DQpoXJI0zek9YF6fag
MbODL2kJ9YqqQlI9mIepODhm072E/XNrnY6igTaaWFVE4oJY+AxZN04OpApIbbBu
2uPBJ2B60pqaxvcoLRvwfQX4QJwah4hNA6uLBeqG8BhAdgWX2xxGbgQh6orCM/Vn
+X02sVk6ig6TvU/TaCpeUFfCljh2RESjO9odFfr7voiDVVyeNyd/CfZ0Gi2bj+uU
TgFC+uvBMxAglqZMoR9gWhGNL1o6NF33gGvH0tHyQGZrcOPxCzqXAeMHsSmFZVV6
5XTd6uWfNlFf9arC1K9tuROP35mNHZiioyJDAbMEJAHS4mkxZk0YKD9bCcPoPybt
pYuA/eyMgnGdJd9mAOeBoTH1ThI/NNDbB0wOo4kKU2mWR2TrfDtwaHi7K6EcuBPx
6B/+EItqXI72gDBrnjVmv4I8rn1PynqZHYvRDkFnqiD1AHofh34k429yDN+T0A/w
SCsDO5buxZ6idW76Yre3CcR2sy4Yhy8co8fBIGd/AoUW/zIq79WCE+kEYfOXHQ4c
t/S5RotGYkX3gB462rkpv72ugMQSYoglQjhp4MG5YnTa+bRvnZsRf5jbiPjvsJ+G
qv203dytfnZyKJdPhP0x/m3BwhDAXcaXEBvUOCU88JSqPNJ8h9IKZdjn2DfxCh4e
Wm97smWd3BnHsVjkTPX+fVSb5biGx5uThzSNk6V9muqVVjNxHU6o5wIjXcy5wnuh
DA1ckq7zCj9N1qDc1rHQzUpDl90xqJ76U+oysyzHIXlGUUhhHC6gn3Zi9okYx1NS
WlsnxIV4u1i6V8JoP8zHmkixDpkeJiGNh+GJn4VBmFoYq333c7226wftIej44P0d
UzsrRz1KVjVmmExYB1EQASYf22TDPvSUgmRp34butS7bdcTqZaKkq8uSLJidXqgn
ocrAZHDVrGotTi3RNUdO4EwIYj7UrOD+g9tWuO8tUa7WyV7DMmojIL4U4s4XSZGQ
N05YDcjhWGkxO52TKAX31DbOC4cWfgLnMTPH87JCkG0cAVeeOo6GGWHmD0ifqiVm
hbjpdw07RMMOYCkX7i2PfXjD3BDs3szxqaYua5cRmlBkJM5xxN+j3HmgGL2+xEun
y2/aEnNyIH3u4b+f8eAPvq+3uvKOX5c6F6RvBqANxpb4NMOAQkfN8//S53O6Gm3C
Msbje0Z2E/EdA5iUV7ldQLIarSHHuEFkFqfr32UdYDKt/rWk5U4mcTwQUhQ1kUXA
mmVMhzPzTlGbVXZKI7+F68L/qYK1g/JjlSCwyHPGTqkl5kvgyv0wtkVjEw3fL3t4
9ou0fxSP8Eu8hFhssxG4wfMd9hRhdiGtJdqIYWofRsmYP8KxlGQX94bqT2EpAvp2
9LDA31rgusQ6Xi+HfblQ27qZE6XveONai0zGWS9B1d65hOCw721d/Qsh+Yn4IZ4Q
dhMyjsV+57zgtCWEa4ALv7GdUQT4JXIw5eXiSoWplDCXWPtA+iztss2fMa/QyTLd
6Pf4UpiUv1BrJMhBAwky9EeYHzR/c+VyS+08crMjppiT2OK/gaqR+n8zu02UCX7e
RGCEbbuS55u6mDf9E/5/qcKZ518qrhErEil8wgLLQCSQgkGR6PgGT0xGQVvzOyGU
uLgUjBvK57TGi0byYOqKVPD3vpMq41U08ED4+KLbg7vn8u8Bp5m+TJ9afr1bumcv
J4EyaxZEdcRT4CsQ+WDFndZqF4PkkVPh0UEaF64AerdFldzPCc/26L+2nZnJIz7H
uNr5QnUhol2nWCSdTx/XATfCWRQz7Y9eEHqLcNkDYi6XLFT5cY3HRFUGzgvXL8PW
XQbF8EiPAPMHcMM+YXrQxZHuX4fOmqrkmDU/GC0Pfe3hpEOzZk0RlthsniqkM4/i
H3iuXQxcp5nsFeY73vwQ2ZgPxCDcFPmteSIi2aX5KK8MuiN0rXDzhCogUQGXsgPC
VJ0AaDKkddGtJm8LRcNYlo8c10NnhLWqwGimP8M9tjSWuyx9ddOpFxqiG2WWnz7l
EQ8PRLkDgZKosGdaoV+Y13baNemuAQXDNntitZ9EGqDjlZcCpeAjxYWfDxijZ32w
eexOn+QSWhGfdVW1x++f6DM2Uon36pzJosmxU+SG6JfEyw/up5R7ZXGuTP++jF3a
HB8n6n5Q89yS2Tlx3FgI4/8hV2AZNu2Vdp0mL9LEkp7XMk5d0/G1o0e1rRjSJYny
91EXGsuqH0M+4NwDFpmICpcMBppPaC2tj7C7NlKD3dYQnbPaSuCgTJRYOXFaE+vA
vTkhuElMYcKAX33YbWtU/C/P3WWclJRyYG87SbY1ec7xIg/QUYC4DEF7T8WuVwjr
b1+OwgAQ686ZZ8Q0xFmvP3rNdb8TeX/gG8Lkn/t02mbfD7KrFxdbjdeaO5HhrU+2
173nEvloucMyFQjw11UbkmSFRpScGSoXPgl+ddbzF3dfLO+nWcpu/JNVhFjQ/tY9
jnGydBFD9ZfeRl6B3gqXoxVWml80GNb5dZET1XzUTvbc77w3tbNcpDg8YhNku6dT
7H/MWP12+W93wKqahlXwuDtjEl1PAzi+yxNHSFkd2uXiAtl8H+NfegOoGWUTWCcs
Zbkxdf472nVxBUg2hRsL+cX0BC05Wc0LRvukz202Jw9fgBOiNcAel6W8VjQaWIe2
xektMStegGeU1zNj2GFLAqw0afUKh6FwS4yjehRTB4CuvCRpvOfLLJIshg2GbYRY
DOCGLinIM4Pa1IcUGnQoOqCGH4w8qoAD86adO8Cj3nsTIWUKyHcrHux9TGhiQqOu
1p0Pd7w7iIo1EWzTiEsz8LTnKuxc6RXK/Zh1Q3OFbt5vt358CRc5RgiawvhOBZmR
hkffs75zjxeMN6Aaj64dFza6U3XTz2v10gxYypp4KH4Kykmf2etVI3S8KAzDTuur
kWtTldIUFhVnFbDZk0KDp4kEWTEzuvStKBj2geYiDGCfEeZavnoeGT7RDdgq7BT9
DTANRhWHpkf3Xl1gS2ECOEej0L60eTxfVO913p7mBz63UXlA2QrT5ET/EoQNLv6r
uCqfOpCHM9kxHn/j88JIQI/P1tRBZoJu1jAxFADH5Im1is+uU7nCQbu/y/HqnpXr
sa8b4rcM5bbJldUnxm6XVgUISWRvIx8Of5+84wvEQ9qtMX4MCM2YkJT0f2K7EtWB
/Cl71fbEyVQtDAXbQvtDJDMIJKCMvCodVT9wrXZc4F83KjvRVoh6G+l4YK28m3Gb
V6a1EuDtnui6jsoLLHpKaBay2cafOSM+lFAoobyXpReDg4Y/hrskW28GmXuJtISJ
ilogJ2mvN3mL06l77a9F2JPUWMgzQixdTgTWuSfQq9H78f+wJISRZfwsmxLDKr1c
gzMSgc5ZqZUWnc6qkF84iIb5RjOJdVNhVc31pNk+l8dxcbe3Al7WqsO6p3jpKzkX
/DHvhNngfGGat/segRyb22BK2xRdjKj8F8VIEgr+9K1ZWJXecrJ9CYtQDSPW+CuB
Y8ZcyP1/msv6uPWhI2vsYaEiA4sP7+rXlOubKPTrLti7ljDB39naFlqPj7QODclo
qgdB+NAtlYcu5qRtje6Z9HrzvFi9RiatzesldpAkTIyccylCysPBpxUP2U6pdXBQ
EaavORlg7ZEYsYcblwFy+af6A5Eoaia5dxyPf5aYNm1tsKnroYj164sAh060Ov9l
KENw0jMILdAIchFRjYVPpnRGHFCLUtRz4IwzPGl1f2pSOd7auFHCCd2KK+f37ClG
Q15Xo/w3l+ZquvpMpbu/7zBLNcGz60BNskqtbAjmqpsf7nKefZnfSAUCCJYphWib
qovJVrgiDeBBbTlGCtOvYzWXD/WSh516ij8oQrNG4nUrhyPmNlygXVzWEDiQrvbG
q8iL3VmpPaBQia2dZYiekGfhgasqTRuoljx8vt+ncFzdOU+A1LBt+0/JvM7o/DEe
SETd7hosjTSBhkj6j82PcgTBT2UzGhtfzg5xg1OLS8NQosJA+mpA2SWk0bBt8phW
FEzPTs+2mQtZyRWxQ33BctY7lzhvzXhb1oyN6D9oYv7NJvdHNntlgwk3iuhQHSTB
kaQLaAgeImVe0lSvI1obmSmIBFTQEYNZUnVWazY5XjxPxNk01mN98JGLmBkyeput
f56IBVTnfM6Oy/vsq/5o8h0jCSWlcn2htoreTA/rsPLEEVCVsJWzdtE9NvipOxhJ
L+nkyQ4/GjbM/PhK/z/EQA6XQFWZoHLi2mClH+VaA2IpXKjuxtBNX4toewDWy+uf
rDrMuH+QqEsz1K2yoj6OZnM9fKzulQPRBsuSZlQleRPMwWJ4oznGtbJcPwcZpnk2
uXCzC2gAPgTyAIFUT6k2vRr0WorSnSx2saN0AJ5BYwFRWxluP7WP52B4avl7hbFM
oDTOQymoOA5TCshnADwX2KLsA0klgmhl6bEMlJYf0BGflqLs9FOZLoKnEyar3Kdc
Y6mkfYHnRiFK42jh7aI+/g3OQpR/JWEik66iGSOGqqFUQyf3T26imlgtz/Bn2vh/
gCSvxx2SVFGLfoDO5IWZyKKvZQlLRhDhtI5nDssRb3cLSaIasqq+PkqNQEyI+GsB
0k+kovBYOsP4Ehsw9NALVumsQJ1ry8K3TF4vT/sQgT1wMTDF/SRgbbmYHGkgSsmk
VYCf0jsbQU6Wy/UhMDPfFAkIK2L2OD+4NVpEqq4oekZUimWCT0UMCHZftWx9LSoK
ZPhkVMtITqjBUunkb3QMwocuW608jUT4U8luz8/9aPyKFm/BnfcgNoe8Ao2+P7xR
T55rbrjTOF+fXzydRIj54OFkdYZQz6aXLe/tGexHlYiS0h9nipBcmo6UffV7/dPE
qzLDE5TgRjXuRE5XzVr/8mX+eru6Io1z4UTZJeuWZadXAAZ6hidaDHr9O6AnkuCa
ZKAnkfElJi9Ey82v6JKhXmB5bCtoUXgj5cxmcd5oQwSRqeQVvu2TWd2EkACdeFsT
dA+oQOx04ISN9+UzOOXdvjDp04G7hhN3DIsQBX3NJSMco/xXZqIz/pLJ1O7psK48
WN8I3Cxa0LbGLxFCWnZR6y2pEjZW7zq8+WALvYlcNd8EfZ7G1fY9f4uR1o91Pphb
wO2+r2XaR1I/VwIFJrsX9CNrHUNEcH1KzgF6zXXXLPwz+lUJOKtUFSgg+GMpewG8
b/T2GIH3xGqPXXGICVm6fRFkHlM9DkNpOwb1b3lXYLflez1rQDikhd1ykC9jysti
tjtKDlIHZcpVt/bW6WAhC2YFdBM7VHNPol6AE3KZQbSVYfE4au/m1CT3JI2Hglhu
rjR2SyopM0SYrXDAJ9opew6mNRgJKlHlAzUm0Tgb9U2h4+FPIYSYDwMjgUO+8Tom
3I5hI8qmAaqJmjZJhqYSx1J9Oxe5GGTToS6/oofKLUwuLF6XedEc2uFXE4ndATmO
uhZjAxVRfJ/DgMP3SVhqyD/0gVHXRf+m2HnnN/8E+ChsIZyI56Z/Krtwe78gCijp
fUofS14s9pYE1TI0JU8wGIw1nlN5cCjI+ir6boftgqHuDbEmaj8oLvmiPdWNnxjc
ajJkr4uL69MMGEz6Bu4GJJnU7uC25vcJkzwet6/8HiVkunEEAohNIs1UGPZ9FvQl
2M/zxvI54WcZ8ErIDm7BpGe+rBgf8Omvg5DkovI3Zb+wOtQS6X2Vzi7nzkuUDWni
U2K6mn5a9Dw5NSsVBYhUdeHdmAQt3tW+Wk6yLfK+S88x1vAD427RO/YKt2pYM6r1
WzO1STulBGmxAN7o7QP6WnX6sYk9UPYthE6v1fJ8y64myr7S9fQ68v0wwWCaJSMi
NP0/h8Kx/NPoIT3stcyAGIkdNeIiffNBjjzXpQHjXUm+YDkn1gFI5rq31FThhoAl
M8+c71rFURPM4Pa4pg/CZv9KLlj6BlMwzx0Nza/A0jafW/rgauGM69rXTrGM80dB
DXvGNyo5R8YyRbNKCCoVopT003Hmlq81VJUId15GYQqas+5iRDthgBFnb0NmU2kG
9xUc0axONotIEdzrSfze0l35+HIX6ZuepxUw3j52dIBOIC3YXpPk9WDf0gEWAk1+
I9CgnDSGRcZxX4+VuheWta+L5DGBUgQDnwPD633Vx+bPMpgGRPwJGXlFmgnCdVat
bHo1BJ6RMgWd58PXvpaLKw2RKqusFgK3Q4gAWlo+k1XV16pBzhcZ9KBIrlZccgSB
jYZ+/9q7G6O7Hd7Ml3vkmivWFe+kfEp3IxxiDpM1sP+scyGaKm3CadUKrMKD/1vx
T5/msftfqRqBea9UNVRM/2eDAeMVU00vHlUo4U5XMW4rfOCNSLTQDISf0SphoBvO
0HUNwYjOagPdflstxVUtLnB9CplqzheFuLqwLVch2uUh+TwLo+D2XXpN1t39iWIM
WH1AUQlTMvBVhHct/LSJayqalgNTLo4oL99BQbePi+HXKIF1eiwBdebrbFg0ZWs9
`protect END_PROTECTED
