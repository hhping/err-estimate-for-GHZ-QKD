`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/5xHfB8lIPcAw3s4R4OnagssPR4cyjTqn1GOP4ApZF1Q5RnrBXtMAlMkNB7pfyL
yHGBB1KkAfV8xGzFAREIsbVj2f11umv/o9HFC85QJPvuncPe2LT6wJNhu/A/Xt6G
SRL5fUToKQ/+WIhAF3XL/f/aAdYHwI3vqyoQDbxGlkjX0x9mf6JxxMtl8QKevcqN
fXXrqjw5ImVU9mQ+1IwwkG8N/0ACbvmWqq2w/cwx1OucHFYMI/KdO+v/C2KnRNLA
2M9unWWTJw22OraQ5RFZ3LQWWXzAYXvheshnoLkoqJHtILr6/JNR5BbM+HTXy7yP
9RIv9O7FELi1S0m/aXFtqdIHd79iRLeui++fL8AGGh0g1yxTY1CvnkLnTvVFdb0T
xLwRVjDeHCEZF/qS4mH9rKqMT3dG3DUHtU3a5UBIDp9O3uFmVbIM7hBQjMuLLOqw
LCeNx4E1noTcOInfGPAhcAanLBMRPLzKvPJr0F2D3Z29vxeaD5lKQ7X/u1ggi+28
xVq967YqNjOC3gJ2l3wXcLq3vVIJpC93rfgQnaa27GSmnsamYuLQEY6mZvHIw4cX
bKLA+JROl5NMy374Jogyxu9yp/OXWqnzecbwfYumGFg=
`protect END_PROTECTED
