`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OzsHkKEF+zy6kuQWSoQ2gYfv5KbFv4A9PgXVA8/N4rjJLIo658yM6EyhO63CRQuJ
jcDSwZxHVk6/txUjk0ftFca5J9VMRr7rlXv9qJcFPrIq38w82VbYnex4ZmNfEYww
84juR7KJY8Zr8SeeSnUNkVJXrMuDPW9mKF6c5fH/iWG2fSuk4u0JRBbfA/cxyd6F
O/vAb+vZJ1mMcKQCAJ++hngLiQVJHsJtdiy8Fm0GRC9BUt+VbKzav05rH9YLSubV
OPO742PQLdc0+q3WMsm3XVtzLq9QkwH1ccKxEpFg7uv7/pZmlyfnfSW5lqJJzsAd
8DWSaloTSEhAfzGPbEFKp25fQYwX9icQt6iWZ7iYSLoIeRiAo6ddycqCySwjHmew
O8d8qK16TuVDcmDYX78iBREGRTnw6V9aHIi3R4CLSK2K/eC6C6tCS9HfgNBIvjCI
0xv9PblR1OdjvgW+iTKnTtm+ZS34JWQQM3L8xVKw1HrH94O5Zi1CGWEv/9UrIBq2
XyjYwA38xAK8FAxWLP2gqD4HZn3hop4hz4po14SyHpjolJ3sdprUiJZFyOYdd6Aq
PEW8ZzSQ9UGBFo8KJ8UcH0n2u4Qo46FY4v8yoydiaR9rOqvXxh1ARMIXNluHNSaE
cpBK7RfbZCBfM/bDYRFhklEzSkILbidFZ/8w9LowPZ0IAd8VvsJpKk66uqXmpJPr
`protect END_PROTECTED
