`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qhTc9R7v/xfw6xB8u3JQxWaEaqAFoiIRpOsZ016IqLyGiolnxNS8+KggWUSqQO/r
pK5FFp/GxBOFarc3Il6yaWq/CIRVWDpx/Llivst2u2DL5ny8O/TPWU+roNHIZ8nw
smqOZfPx3wuRn85S4BHVESqWglVnSpJTLah5eCeVv3dtphH5LJLYVQF7sMrw6xpo
X6KfydzFfvE5DaDzvMee5KW330Wrn7oGIQRnZv9ANSsEWXBPMEBBZdsTwwIWAXNC
zHc43QdXDbA9Cw3BKgUg+/8Vo/7GyLT5Y3wFSt1dQ4DQ3PkDCGDBykXmVjjvAer8
9/kAHHFa8k3rQDIngnj6OiNtBzZBoRjIik/k374zMPIqE+nFJry23NO7iYDYrNKx
KyDP0E5jCioxAKAH55rYdsqldp67NkOU530Mb3FCZbeGYYSqgRuwLQ+QcpLNenvJ
sDrTnw8w8mTN7AB5rc8q4xuY5WMAadLgNXp1FDSAjCV/AN5RmpE6lOvichxhVnlA
rGvNcZyH3iuwlxKbHm2pkXqX/B3ga/IZxnc4lU2hq+wk/gvmv5MdYFP+gIhlQ5FZ
0noxkzzv+5+f2zjI59/FJ6m9hFFMU31JIoSPKNm4XO1OuNA2FbaHLwtsfNW/I71H
h+W2bzx5SG+JW1AeKIN7BmsW+91jlf/v4/LSvvl6ZM/peaAUVKR72i5e7dT0z42S
xs+6+gYm964khlTrdKpA0A4Lnjf8RjjnUHvjxGzxjcyN3KvjgMVksNNJGrHQtFQS
u2Xm5cSzT9w1xV/l2p1B6Tq3WAicb/jKfs6TKQ8LCWg6qkwwJWHKGTkpYnR+fzna
zes5RhlJ9PmEFf7w0MXntZIz1ySiMsDQMEAZbS52qgQTUk2gtY2Tk8Je3bjFdYwn
y1yyOJPjTgzBJePxl8S3pEGG1Ni97WZyXDYwFUA6lR+zuwO+PqLz3C//YgjaK3RL
aLeGdg9j+hBfTlS+ssxr+aiN1PyEt94jXKk6WM3ys52Ty76O0NHneRj3zb4Hgf/w
2B6e2sRWXNfaR/FzdS4ag7Xw2JK8NkpTnfPIVkL1e+UT51AsI3nnhouNKG/y7W00
mK0GTMp4NvPOpiZ72mTrFmj9k5c4gX1r7iSXgHJ9Yxp1Qip/UTl8lczifvOtfoPu
J5XySADZIDaHo3s/JfNvoizgIBPNGFCvPWPo9nX/jbh/xjSiaUOUz4pDL8v6vOUq
vs084aGPg8t1hAjXHDt4Hhw9tujyfj0db7GoxK+z9FHJVSr4LXhZEUUG4whLMk/g
TMmlulFkUOk2Jyg7Q0otGR8z1gaJIxpbLaIbaNn3w/ehMUBqPHNcvi1Skgk/LtUA
S69Wu5h/XV83gC5PopCfSO54SMtaV5td3bv8FWk06h+0ahkClHXmyvithTqojcjM
dPmHRnwEzbEkBspTp6Ra8XoNDqfgPbY28nSzPWXoPRsVZG+q4otR/LMi3GoO4E3k
Vkw8Ozih1amn2joluu/AQ0tOuEWaW+1IDh6MBrgueFkzqth/MscVZQkPzfdenYV5
efBkELzr7oqhcujuHviZcAq3BHr6N8eLwbko1L3onOYvBmVLBKHcK3lsWQGjhvQF
/SFU1VuUHbWu/ofJjgko7cUA25lTqkWU12i99iEtPfSHtowPS3InQi+Sd9/GHaR5
6BK5vShihzJxDxygov5YbNuLvYgIU3nTIOukXHWyF7L/zKgdsB5CrzPA78HxuCxu
3JUiUsNHbtQ0hCDDMBZYCQHMbnvad4NTmFQ49xezWeUeQ665dtuwiiWITJeb2VcI
kBK8XtLscMxgfq9VRk+7IJW9fgZpeCbl1GPrZBT28sbQ0ND+gEeKWhkUp2sV6cao
vDve/10vRHrwo9NOnqMKe670ZjYhJC/KDNU6ZPfx6zUk6BNbSPNZQZmMIRXXWvDp
KFg9nLF0FSPmHeDlAMAc0c7x85LSR7Fs25y3p08qDPeNHYvzvs918sp39K8V/eFH
83H8V/WMzlT3Ro24+9fiCmmGSqeYYmceeiGKVbrcUj6RV2QyRbcMHm4bTRxkKxp+
kFB5RJDrvPS6Etg/RlrcJmgWtwrNJfwDPSR+l70UWRPjFGvTv+JW5kraEsqmYuPO
9cNeD6IRPbRxccay/+CB3VlGTmKwzeC0XUsKmP+A4Pp0gD4z4+a94PSVugClM3p3
e0b3kbbdF6haIfzdPQ/QrClyxRw3RfRmViTbZUO1S3QVpNyBEdduCmYsajVz9Aiz
w8yjW3pXomG8mTd1zd6m5pQB6cDAnRyCveBB6sKYa51hsVeVS/Y+7qSKFQrWhwXo
Mv55GPu36PCZUDjW4islA92dHx16Xt6u71zbBi+7YbND6sgxNVswADZJC5b8XeIN
p0jgyBw+UHZkisH+2rgV61DvONm/QNOIhtMlrxDZTBBmTuo6J2C7s3i1WtvwDrAd
HozLC1TpUuP9kQSCJt4xqMPg+rWry+TVzNdIY5yzrurg3+GDsS/jAtC3SK3o3pMR
iMQyT5s42CAgdJULDIDgNSyua0X6unJKmEIhC2+7gnmw0lyN9ynXJvLT8nGnOAWR
PlrKQoiK+C5+c3PQTmJFU26FcFtSmRwEwYJW4YlQcKvfrEg8zyePb4WgFRPJDpHY
ERsvvjmUQXSSLkcFN1XTtdvBdDWxuQHE7aUsJWDK+zU8V+PaXE/vFsKvSZ3CKC4S
KcU3jKfm0SaKESR+Z2psVo0YYNYIc9KQSvXGull2D1PWmiGnqrNE+MbMDLvIh/rX
dY07ifEjtNbdFAg0b627gV/tZ2KPIZB0tCqcXzw6FmGILOLq5Aew5a3M1kl+reTb
iGbTNPFTcBMxmaJLwJ/Ca6kq9XyoHqh9nDWoJmtIcL2eq3/AZQ9cIuGaaC7CeH66
iCoie3iYb1gCUJogdn7pVHTesPQ8SLC5BhZGiVHwQBpByvq8rTeJxPhPbSGdpdva
dtGWD6UcrlX+V2Fqr/JtZPfpB5/dxw9tzf+NUBAz08lBIjdqTBL45UdcWvoaLVWS
CYD8yNX/lTJU2iYCLBJA+W27wRWvcFsblbexRIKETA69hJQD2R+94yq+psPjl3av
zbTdJ3RXxcRakAZb2WAtw8Bau1dAxIGsU2nMVd0ouCom2H09Ca6Ls72foT6WvF/S
igPTwNctDidsTy50Kwo+RHR4cyzMlWOZTVL8o0JsUfLQNgE5A/qk6XpvY+ojpLc4
SUXNptS2AqQLo8GS5SMCeFVdQ5wKqt3URsSDUYpt8sBi/Lk7xWv9TJ4DPVG6uHOI
ep6vSO++NtKeeozO4HiJPSPdKHAJf2CITyR0hPPj6UsDPVXDWbTzm1rwjXyi2jfT
UhrL2mG9WM9h/MEE27Z0e4IP2ZAr0SsXqFAUJIWoKJAwq7BErwDLMrNpbf0tJdNx
snj/+Fno4GNBCIdQNDr6oy6ABiCxRBCHNnbVCRcvjTn8Eje0rNrmDpUFeUNLclnG
jLxh5QSkKartJNTQBs0iV/P7UakA47y6nQOFiux/rzwelc/9KCK5C0nER1juSgjA
kFbRbPc3ARagCS9576D0EoxdkTEbB62Zce6dXT3zdPkLJ6BSwucLudmGE8MQwpDA
xLMfUgvLjg1gs8/X2n/R2IHUH+NKkN3Qw0z3WhKMyG62fX8m9m2TcTaIcHMDtpt4
RgTy4sFA0ZqsOLjdiKr7Lemh6YXl2x17uqs851tH6tAj/ZfSI190U6Kw2W7gseKm
9qhvXBRpz40XiweOaxOPcEhqXhl+TvzYitqPMXXLc9QnSREGBOF48kdgi3XVYP5m
Zy5lCtSlYWPZhshTtOrzaNAleqFqjM4/lAQzDi3/LDFvBw10AepasQ4JBr8/IlpU
fc+Yztw/G5ZwO0mZeNjFAlmuJwSYgo2w0J2SCHnDOlp8Jn9xPoi4fkxo+/j8f0I/
pO+oj9phGB+LfAqOYd1TZDpnqGVWYgDBp1QBiGaU+/LlCEDipZgP0g6u+hpn9BHd
bH3VYVA5zv8GEEIi3stLGf5D0OfrYluQ2k6XIHxgFyaLwpcw9GlnT+dcS2eRCo9F
bexp42vuATFHNdSrZEIn7hcKxsGBZe8F0zr9/8KDP7MBLrfITOCyOEDN3l39j0MF
x3Oq3MOVGiMu729VNPe1OmqG7AewDpp1asroWBG86RojNd3RMPGp+hnYsPQzzNK1
+icZedCTbNYjTN7kpNNidlzzaJIETDYjxCD1OFBdmDmU6ehc0H+GeAsRz+cWpVTq
hBLT4o1XL0zcT9t92+ZUlY+ZEoK12a6tKOb8k/NFsZR4yWIVGgxojNYh0MLgPirM
C0/Ar/DoDQuJySHWLJaEIUkf/FqjNlCGV7Bcs5iU5dIwmY9kHhtREtdTiQrPZQkG
YXx/C/ExnUJN9LzW3r/zNpocdM6jXrsE7ZqzMLQ1ShRuvWkm3A3lQqlcvk+T1U2Z
XA3ZNRkqlAroylom9y5yxHmHNc9D6IlF0TjvjCWbYcL1USg/gX/WYMuSugQS9il3
6y7R5kFhlJAIJhEMMZKOtjsKbJS85zSeL6SVm59D5VLc2D/i9jqfBy9dEDJ/8QFB
mz/8/wfFMePEriSuMgaIHrkRU6VK9eOg/+PM4OhAfJ4Eur+I4Mro4j3Rr1pBvV0U
6avuCbpSDg0aIEB8R/4r3ECxdtoelv0El3zxJok+pCIZWvK6uVMRe8uy1O/dmyLi
vrRaotG11D7U6YsGFd82zJ4sgmiIZCBUexWc8h6XZgZMFP15IK7OzeYnkEl/KhR9
I2JmqZ0NCknqv01zcOrD27DxhqRIUIAoMjPwBNQCrXYocNXwGVHXQlQra6JPqiJ6
5KUgbGAFwqY7Z3hUqCg09313XLqmo/ZKU2Zz5rbhJiQDegp9NSRgEJQ6upbEPtav
YNuKzyEnVzZscnhkdJE1/keXJlmwyEmxHQmeyRY9udO/7TM30xdvYwZ1bpXAcSKZ
zTFrCFDWqw0TYq5ATiC/CYZlg5r6auidUCL8oXp8Nsqmp2RaknP498XFB8AXvHt7
jyaZkEZnJuUhUCS9xOY5R8SG3yxSX/IkMp5c6XN7Mx/38ZL7wO+PxwGPObA4UdIw
oxvslVChILunBvOlZapXuoIqvH5DIgJ78hqE1Jd2xg/6Djnq4w8+LvXiK8sowQFg
m0Rfi1k7fwmP2fB5deF4KkzRBdXsR+WqlaXkJUzpyQxt8vFqqK8TS2fR0ozdj8YH
IE1vfx7ONm31+KJ+wQzVKR76xfz9iFwVMVJXNoUmsvi5yDZny2Q6/CoUhC2UwI+V
y2IKxLT5KUudKuGZ8n6YzrfIqVzbkz30XifmyQZvNmIsKnPd7fwdK/8Qap9RYBZu
eTlM6X/eNY+UVRIbz6IUqwKKbGGKj2k127fOxNFq7/kKBunAR1gsSuoW7QwvKhif
6IJPHgdjoz7eavcZe8lWvdkorn6muFraKZHwW9eckxmvdsb7qNYWEoZfSpVEmeSM
H/SDgA69BdXYZ0yv3mJ0qaMUlexCZv88G+I8Jy2WMVzDM88NrQ9JNEszA8WGqsS7
MLDc/ZoeE4tWzSS2z1yCROV2lABHs96KERvtXUsZ+xMnPgf7f/eI01e7ya4hx6Nn
7YpXbaRoKAjRyMi1cY2KffEUMqdLJkUNzDhVhtq4Kbf2ahYp1v/wGdl/YdqkZ1+B
pCYSlpe0Ma7O7s0Shg2Y+zblQVIiLF+F53Xp49wQZX5W2sKVRZNoNg5gA38U5z86
JpcGXJVAiVS4Z0SlLZjaGAykI/FMyutqGN94aQS7LSbVch7LED/T8Cop2ZSWygmJ
cfurwbJBM7KrFdCwCGz0Ffgnkf4974lRJDycxWulCzoDQLYJU0SkDyYzilHJUBnx
HoBH6SlqwP/XVABS9w2GCcwDFRT/72KQk3VfTAxgrCLBQH+29VPud6EuoSQ5BbLn
fjLwjuO1OEEArVMAAh9VYhLQuqBoTiNiosUCb3VKcxjUi7tuY4gFr51KDjFq2XZN
bfG7j1Ia3m6uByQ2b0uiu/NhDUCshvH/FYrdIloYhpPGV2C0VWLwKsFduxCkz2Mi
F4EacdGyjBC8GW8LsiNN1Vz1HYfNOAmkRehAhvk5a93LS5y5DA1igx+RSFzmLPmO
o7hyGCdL2ttb60yR8T+wqZb43Ze0PfRbv71rlK4HAX4SA4o3N7rhZqIk5mPZ69rH
SlndIXR6Z4X0gTdb/50i6SYnhGXFPYy0KGicndBjkhf8b8xtjrJO6CrTWA44tjh9
yZ/ObzQqTWolVNNTYFgLuTYL0jb3r4yUczc0No/noj0Evjc61I5RvBiq93xuM4Rn
YIOSZGqWxIkMIYkyvW6A7bg90IWNR3NiRWEQQMtuWgsBZKrQWd2+WacGcBB6hMBG
sKV+qdk/MMGv8hU0+FKvfmN8+5TWbdwunxEz0xBTfgrQV3JcORKeHBLRFkAe3+4E
qtSuI+C4wIRiy9eEIK98Ba5posByetZdC61AbD2D6CQzk6EJl1eGKMorQr4UCCCP
x0aEpG7Hzd88JPSLA8t9EG831oflwTLG8NWKZNDl0HMZPEQroQuysZWlpsijmSi5
IiQrk5D9AuMOeuHXmFFEdLlTCA1fE5v2+j/elUP87NiVtDQiie0aRj7eRuNJr0Tr
fD30D5B9fuTH5O6i0Ecb0IDWSbCreRfry+WFWi98Nfl8qguCDbHW5vtmT99YqQMg
OlCMloMb/tYhpn1IHlIt8M49nfi924D8WIDIq8YFZO51o+l/wX8qfOV9j2bcsfnP
TqBsu3ZwxruSwPwV6DbMN4EkX86XxKUFkGVR+qtNSftqOIFags5QZDJSG+EIZG6R
WaIh5TXmBI5bde8B1QeRVL/FHDBta9/IdWC5AmHAH//kFwL+wFTIEh+8TnqubRBS
dd2ZqHTonuGY9BpkazxnFHorrJ41AUTksOlNyuUdoz0Xrn81nrDNG4/mPY3rSDiJ
DctNNVL7ApY8ErDlsLqD+aNjMmLt9C2FfLjvaaf5nePY1EvbrBhMMZlQyvcXzBpG
r0IvSQikJKah+sTHCp8q4Y48JalaYcBTVQyypr24MsjKP2Wkn9Dl5DVadotvGy6r
dTbth6sCm7NriyioSvP6UuoYBlDJl3b3bI5UoDGjlT4xsC+qWiC9Fto5/qL/PX3b
cm5GcVDLMSRl+g9XgCJ20hBYnqTC3tATc0hIgdbrJVtwonmusHWUElispqBx1X/K
U1mEVZgKZTDqmNxosZfePWzFqOcS6UJSx1C8aj9IPnBt0LLJ7eTbBwffEZgjbjJV
bQ7HLL12yMJmOtm/tzOCZpyLQi5NzIyBkDjpmYiKa8dESp5pqhIRo61HhrV5QYnO
BkMdmB53QzX8c5Co48KT6C2PiWON5t1WZtTRdgWeg1kc41/L8HkhNeWhl9P3qf2k
iC4AIhsLy91r+4aQdpmdnzrMH7r81TD1JXpThuACigEcDB8sZQDrcX3k4kdMOOfc
JHURT02TIAECfQnDNsRveVGciOE9/m2kh3Zo7u+9n+KZk97g2PM0i3m7Cd2p+Zjp
7nPJC45uxywE3zgvooHTxgxPWTWNeCjSVFVuPxO5LbmGOUH/tgbHMrxdowyDzbhx
YO1FGoa8VTKvar4hFD7OZMIQmT0nUrr09niHS3L5Gui4snkatr3A3+QeGMuiq9fW
UCVgUMuBfCF+EOE35iJsFPGxeXGU0da7k8hIE1qO6b8zn65gXJuxXK4dJun9llkP
0T99pRmFYfcgJFMpDqW+4KGESoMSqw1dboL0MeX86h3Db/hfy/ZqO57m/kHaMwHl
dBwMI37482fHowtATYZldyR4Se3QqKL/fIbsSRJUO0tx6NB2aSV3OEWYy4Anprwp
LILvculJ2o7BNvLBE5IGRmtVBdP2sJ9H3+CSkpb7CSlPBRzT8b0e9ernJgZN2CNj
Ot2suRyM7ZjaJBP89Ot6o/u8Rl3P07pIp6ElFWpjs79XjPCqrZhnQOen7fK5Tcfm
YjP+TA0j6qpXISI2XrX7Y0AbJ7YD7gJ0BOzvG68zTYQtwtREoFPWsuCrTd3y56iv
NDMFSipVTewAB75OlZubPzjyM2wonAB1WK1LNc9ArLAxz1x+6XSB0WHeS7m2xIIC
61uBWF2VUTIW6l5OpilIhB5/VGAHzBBSZZ1yNwdzgMngRa5VGQ/ePvMNBCW1Lowv
Ydso1uFr3pwX1LjhypKAQAhPUKzw+tf44Vzjt8kYPLVSUCsSpnLwWWYl3SK43huG
aqsV0mnNyefUPcAh8o35ZxNhYkggCXYIpjCYUJzDIuWDMfbMxyL7TLF30ubGh6v5
v3XlyuK3qg2SDADxTsQXPXi4lGgPfvE8bP2ZudcG1o/nMMmUKBI5lgel5ju8NMIU
Hj6hP+bhbM9h2nYoaXf6PIDq4gaprAQRwFJrLtbv3tCPlnR/AD6LFGU8SO/euUjv
tcuqydk5QpvS4Ih1VPEziZaDk5MAbv/OcBy3d8GJIX2eCQ4lIVS8L9y3QubOiOmv
ED26EfUiN1+NDx+u9xnDc2AUk5jbl37qVCfOJppoRduOyQhLQBjI70ppy4qfNJ5s
28J+eXLcS/3os5pLPQHOC9/pVpUN2IzPQaGGzhJ1J4sJUy1YNtUpeewrHWTtXvB8
0DhezuVVHqa+e28XiE8tC+t8uwsLkF5CgCpnOyQHFflrOutzAIXLdKr1Z+Iw70H2
VqnT0RBpxyWFlUKlMoUClUKhLMXs+gPxmnrA50UAh4aKi/2YHsO6NC1u8Sx7u7za
99kToCTJlXHd0dlxh+fHFoWy7YIHLK6doDHFmB2GuaHMGh+Zsea5tttawzQFKNuO
aeFtsQ3s44GG0wND4MJwoumox2eHkoTgGykPsZt6XNL4FPNn7xW6N2jdPDULkOTE
pJMKQ6juqAR8VqKJGLP2xsHcDeNSWExhso83SrkGX2oWLUTRv89S4qe4xtw2uEAn
FQFZlu/FqKyf9BI+y8dVqVcDvLrpqf4CS9S6kDuiUsVkv/9IEzCB6Ov2xpEWFmNS
Y8u8KxG7FhhfkexBtyR4n7LWjdqScTy/7yYOxf63lIX/ToOoV/y7gw7HZiNrkQvi
ysvMqlpTEXtuGBsOkppN8K4/B5lAOHw6d7QTQpbvaPbaPM8x8yFAfJo/hJvI/eqY
yqj+V5avitHeaEMUnyQ1wRy+ZJRHinUd7WeCVDb+mYOYjuNGetLUaPIZw6waTwsj
30iITJyAcUcJTKlQnTAzXs+bLkgEbueli8X4C7cpGiTcIk7lmFruvrW2kKPBmuKg
d54ZsIsSVk9UtckMRQ4UcmuhkBL+gxrRaMx5vZ/RxsTe7fJ8aM9P5eIA9e76984Q
tcSpn2TbxPsnM9RpHnFL/SpQqIV3lKvye38ahwalYGdGqeFH3CZR4RS+FUU7YERd
MNbVzi2/yRO2zY/SG4C5zTyyvauWSfIlmDbDByft3JO+Nff85iu2XcNeK00D4n+E
GrQE3fBZijmqE3QGPBIdvbe9FBniE9P6+0X/CueqtBsJq3IxDyqYbeJppYXFj9rb
A/8sPDFmxxo9JwuwGLvJWfxM9GREQoZmFBNRfFVvBoaDfZ9QUYnW7o87u5uAWpeq
YMOc1WWW2EpjnYg+oL4kCXyre8Uan3PJcffA3AHPJ8l7dSgl9S4f6nUkpABBpfRZ
YpEt1LUl/J6DvMu25OdcSLr12mId+y85z+5c7wLWigbxV83V6PdQVWGHETbb2RSI
6dWDeCNGIvKEh6PEKLDozs5sBdiMR9LCZagJ5dMNGHPVGyypjh39r+Sxbm7jygRh
rC1V91ymkLqgbRrNy/SdRwzAuBYujVgXyYU+GbvOzC/vx2eCZUqqmyTJ66LCJQGz
Q8Hv6T7qSG+gsUEBBnRJkTXtlWSLuGuEhoxo+wRb+L0ARWOjSQZvBsgZwr068DGl
aEcvU+rIGOBIYbJKkqHF+6Fmpi/MQOfJlJ2DY5FH6bqeWhsr8MdTbKL7f5ewlm9b
uiIzI6RD65Ailuuoe2USkrClc7NvX484l7F+P1hIKMN4gWrT6cZHi41YmkIUk/A+
Nh3btRPvRkrHy2ovGBkfQeLPhE0qnKbQKX439ceMi5Kr8TKGTGOj0XUfjlAAnbHv
9KgF+TCLUHZphxhH92bCMsIECaTQrcwbFFL5L2Bbj4HPt4OTj8YaMg41ny1DOL5a
AI+zlMjcT4MeGw67qMaBfkTEx/DvVIHiMqxlDn4SpZJQJ9eDv748bRRYhHTaVxn9
q772UgFUN+ATWtJtOzXTvfeT8Ox/LkdEvxRzMtPLNSNlrq9E9MG7DDP6sD+E+i5n
AC2Jj3j5dWZpOwrAUueUYaEVwUIUaFdnSbTV3dEH0b+87pAxOVWPevVc/PbFyuth
rbw+LkyX9CeFAuuCL1+9HINeMjVqnKcdG8Vs7jBbXXIGSWvVUmBbNodbWirz8kac
qzxTeGib3Zbswp3an5a5NFPpbcE+/8COw0KCucjYwEt7N/XayspstuKN9NR1T6+8
IFLZsuPWb1OQJGzFU/CrGjSJd39v/MxCi7Ntts4llTEfUxYKAOu5wJtv+TcVUIyV
j/pKq9l/LvhKyC00hCslNPGzPLInXyZf2zUQI6EhO0KXV898Rvh5yZnKqy3NKBTA
YQJkxdIn/2UhdUUX0kl9kZ3ipXqaYliSIP8jyBX6yVzKQ9WnQvjFC7nBX9xzsBaU
hPwjeRCBCl3iWez4Ag7XIe8Ypm+x0MraV06ktBLTdnbaKrc/79zB6Cm89MbKdvBo
LC99r2nkOLWn/VU7IOjKQotBUeBqGDsZHyf5/oiqi69O659C7HG9pLrYQe4RPxAc
mp7I8RvdxSoKOI9A+tPiInuZZZspxUKplepLwHS/RgvuF4H7Im0olOm04TeRfUNk
ci0BB25TNbwi+W/eulMcrL9qOuOypOepWxBT0W5kIob+6hXjf63tzL1s2Ekb+DZe
bfox7OvX07e9pEHIm3WeItrVTyisK7nr7VuT9ttTnIv3zV4+Llrtx7xI4Km0NLxH
rf12PMET3CqixUEHAmjinat61j/MqcknOArJ0w1EwT45toJNBUI1vgsy8KSLH+Km
X1D04ZD3Br1uZZu3Cy11V/sw62btXnmktTqXBxLW8mINZOueNR8h7hTLC2NMIiXX
ovkiuA9C/wNfM+lb0FyP6bjH2MVoOCx+zYSZiYTYKnfbv3pKzU/MCLUxAqePBJCi
zExjMTdJVf6lqoAaqme0ELtysYVTxoe0w/Gc7Emh7p40moSANVHvqR/a6ybwj4mQ
tjHKgk0XCldGwZZAi7bU8Vz9YcAcAq1MoaU9qNFvvN+kfi8gosHkoV84acneh/Ak
M0kSC2SW2ik9qvXuxy7Sogy6gxRpW8Kii+sYjvfz5Z0JuQ9PSAOoSpMtrcDgiQT8
QYGSdxvaRrtUM/i1sUGmAavaGMjlm7MYJv26Krf4otQJk29fgqxDZgMrK4LG1FfR
4aADJpsyN3M6RLNLYEMZEaxIae2NKXeIGD+pcwZagJcCyLxcOK4mgdHm1xiwhqGQ
oROnn2UP+YaD4IBy+dsjYrKValboedYI8uh1G6di7Rkyiqgddb5iHcneZ5LX6J/Y
b0O7WiIif+gVtJfJP6T5Zp00b5Slx3wpWp8jQ2dsNvlr4d8mIEci/ojcrBhBQAIP
DUpYXsCSadqRGA/5WI5xV+tSoUcZjZQGooU0vh1/TZ0010kWSUjqt0cPIqNBshSU
XVH3kBzyjBKs4NZfrRi+t52EbaSQmfOQBoEWaDMvPLCZC6atTRzHz/254/UXP8dS
sjJXaHvZcoy58wF9TE8l2lEIe4wjqlwUcTMrlvQAzKYezkwDhKYGNZACeSKoP3VC
TixwEiOOEGshbWtunsz6w9HHv4xNUg2ZY5yurpIzgAn3wcRmaU+VJ6RRt9lBW2+o
wpU6nXrhAKq8qe10kIn1g2tLpBy8moLbhmEKkggvXBje6iMcPKjUPSCv6vdbRQCv
cgkHbS9o+mFC9/Dw5J9k0T7KBk1zlOLDj6i8a3FicaTNZjmuvb05lbg0Vu1Bx+Yp
ZY2RLqRSz0bolkr+RWwHu7cWD34t4ZbYwlFz5QzbsYevk2c7gNG7OAs1isR6/7OZ
rA4oD7hE3EnFoYzu3whmfM6xmq8Xk/mXn53C6rV23onx6YlLfyG+rJUpgvrCT2N2
XmYGPVs3LKiEC52nDFmoRZo/G1QZ6dFNqc/N2Q4ITzCrn9PD8oJzI68rft47TAe4
8oSPuLNOX2x/lNrX/l8/o66BUnXHa95PzwvFUTALCVnMb9y3b/mBInc3tf8hBsqH
uu4UgL7/Kn3Tv/jXi24u+2nBKz2X8ROHKPQbZMyLk9Sofijlrr6GyEhXIJtql9ds
j3CrTcL2gurY9ivMui8YQptoAm5d5+/OgrMbAAzE+aOaDIAx/0mMQL9y+KiSXG2W
fNKpZFij+Yd5ZHsuB2C/O1gR7zRPrhO+4CsUGNCYksE7cyIW5xFHrdwjGdX/38Rv
dzydIaA/16ZzC/BG7dCfWAAUQVaV98J9T1T4Qh+OquXfbHcMK17dgXL1p1uz8NZu
Mc1bzRFJSPdVl+PNR70cF/jIpI8StNTqITG0JJ6e0IBrkKe40W5t1mIetUkyUijh
HxqRmN2+/lO+Q5OOlruRcVJ3UZv9PVmemyxqRT31iOa5BJqyH/+zWSjQo0lArMLN
aQEIF8EPLz7i9tJTQw81WK8oYxc65y9XqmnPtl/uD/4CyWIWggthHNbCijSnIl97
QRIJcj38UtiLmdSwuvyu+t374E73jwBacCOpSz2GJBQi5BQQRKd6hzDvEnhc0jsE
O4KYMwxo8N/cgt0ZtE5LsD3pBTwHHrK+Xv5dD+27A333QnH7GZhTzKpxdt/g96sJ
eYxJ/TvRUSay+dC3uEpbGZQf+tOMT4CJO7JHkoywApkN9mKmt++/L4nXslju5e25
3d3UXIDdHKDuzxvLqXtv4b4+0z6Qb/ay8Ue9vvRijTNjWCJwOq3rpfreErFs0rB3
q3wSZNBXK3Ipr9nL04xICSsjosB7BQmmsSLMgwdiBzx2WA7InRTaf9zTvIkhBu85
2OlClw/0f0u/UNkipGFz3vMx1HRrTB46VluKil/CabX8QDivpQYuwoX85X+FYaHe
H10do/etKtTK9SJxklWDKYATAO79wxQ5Ck2K/kpdYSPJnELnx2zy+7Lw1imUoRx2
Tihx3AOTpBCTTrHib/K0aVVseM0mAVmAK7PdVJEEwjIIvpvfbMLEJT9nrorOoNUd
vHTMJdSjRdy6UxMxBFhDZEUsh5hNrB7JTpqiwoVuu/oudiAD9ZwvBqaNzpEEK7JX
SSsuMtlhJBN/3u2neSy3V5r67Fjy9MsshFog9VjSqsGfqtMrgqzh+TCM4w6VUQrz
tWMpvBleM4iW3DaG1uUnGPo7H7UHpFh95qudEumaes3YyzLU5RV9aqk2GZ9tlJko
EpUG4bkG41YX1kIBO98ZzrzciNm8dEbm1mrpfx7IyhF7/YMLPUO093BZE6gIoLQi
1FcTCTkCnbfGXi2hOzMXfAzT0Sajo21aiS2vYEnfGxzpvBRNCuRwL6gqsquFI+th
sY8QbCs0bByvDUz/uFcIxWejCBSH8WAR3EYTmfvxKJRgTbCqHfkZNsROYnqiGWBe
R1jcIn3VACZOQZkWD0XgdRSxtn5wOQYukv4PqmG5hx+ybi0jitlzxDfg1qftK6ck
N9GfTJeE1qzntJ1NOI+NY7QkmwN9V98s+cRi17pKEPPGi3Yuo2T4jJT2IoyN/JOe
015gw+XbZ7jvLlWoPU9FOoH8poz8Sm3e2PUVQ0E42D17DpkWyAE+ThnXPuPyRqTs
jxJs5/sYrvLOmG4Y8xQ3SnBcYMlENjWDCl9ZCu6DlYtuiSrHxwy6EVGJRnprpkTb
VOBpeHXyCAxQ59pK5cBet4oI+P3idffewFStEBDbicnoAwgKNLrnF7L/yW+jQSpg
C31sFHuOlzG3rOCPvERxpvdbi466eEn/85G3/tL9qBFOSClYIOqZw8NYWpBAw1Lp
kJFwM9nFnsZroVnT36S+1IMCW1qiK/wXibqugSi6MoNdLcDuIbKYLWW13LqK5Rd4
aCRYqpM8plJxlfj1ZngQKFgqJW9l1AS4nRx6QjLI8c73RN0T2fHka4G7Qzf7D70C
QM2rHMcmOkZ9P7wTxCZsyT4j1+G9qUkNewr0XmUdAlrAedIPJ6MZttxIUyWRtiZ6
7MszPafJj5QFSdohUk0/UsVjVOQCRbZOZuRKQbHPpEGyEzM6BNrHNO66dAtF/b03
Gsc6nCrBZczx4i8OrkJX8PsBldzA5uYPvQ9cCLRLY3HoL0sBed4eXaN3Wd5YX9S8
o+XSIkpFv7xTyCGfX0JCl3IR2XGG9U1hRb6Yn/DPWQsdadCOIY49EWlOGsxgAVcM
aointzca4JSlMi/YDA+g93l2A+1TmduuW8cETtJo8gCJ3Z8IlmqczMH5oX3dxx80
KRJvZoU7WANpyNnyCi3Fnrf/w56hsYNt91sTXGGFrn7/DPM4no8dDrPpuGNbwx6f
dWtwGukoFiDMmHNbzGIyP0Gk0e0xJulgbIF/lBAa1LV/aKLUad10pS0JQpj/7lv3
M99zpPnj2yZsjyhw5cTrBdH/jV5Q6ixkwYIrpgBNic1PBr9Ag7mt77IzIwFvC/Ko
kjP9FzIniZ4dcxfOm3OHNJHeC+oEWA6G9dDyhv3VPTDzXSoZYcCj4gNQ6b5QV3XM
mH7Qo5i5t8g4+kLlZDpfOUoECNMGW+CSqV9UmNXzYfanfoz4wbUh6HJ4K+ayT0ez
AIN4soTrAGxCULijh+I/vewCaWmRtNNiUURtHlkJ9E/tFvepk+lrQKhPppeubk6W
l51eSXltf3AQBJAEt8ypSdIo++7Oyw5PS0gStBYHQ+03DzALTmgyWur+FAEX5kIN
fzz1mBJMF6Jynf0uAxq46H1t1v5dCZR14X0VcvEnjFE9Uny1K4d9iba8eoSdQe21
mHM/vXJ484FxG/CRPDVQlNovq76k85JrM2VGOq2N8p2QbCN443Bazpcw3DgBMEI+
hpj470dqJgzgLZBL86G+VB+nkpJHBTee6k9i7taYfc/8gZMV+Y2Je193QZNd00G8
m3pFQoWyg4Kanu2Rulsb4VhnkZTUD/THx16UkEj7xzJEknYQMuYz2zEGjazMXl4n
r/mox0Q+fVBC6vVydeUeOTrMpRYRwGoA+JrjrbPq0+7T0vq3FkNtPHSg32eMvFWc
h/DJbIWH/Ilcw0OmdrTeVhs9n1fzgU+AxMqf3G6hUVBgBjwlOldmz2FKRIkjVLoA
1PDGQgn9sc4Wx5ByLGeQPlkI9qQU/iroVZe6T9RGqH2STYUk/VcMRVjmWkvmWgDw
AzFVA32wP+023bsmroD8z3VVvV+IcTboWlarzNRREPYioPx8Er9JJFZum6bMcd7W
I3XAURZJSUXRu2C67HS1EPp5ghAnzYA6nCTndPT4FmGdWSzzAkRzyUg0sW4PYJP4
2gKu/ThNDf4IbONmvlq9ziCh77neF2VUSE1oFUN2uv3xu4ixjzV+rzT2bzvWjYV/
yplOtOqyUrSaJOgaQSGNdqEBMqb34rPEhyHQSuw5XkGwo9juLgf5+hn22jCbjAm4
L1XNvvNZVbc2Sm9rOIZVgUDDdpxYfGCa+Nn5J4sOagtGB3IhG7KlF7581YZupGfd
h21+3hEv/fcT7+563JI97JT2guI28Fr6zNQvJ+eWbFtnN3gPiRGOYCTBZVaYvN0z
kfipasBp/dThFZT3lW1yKN2Rk06wz8xpG0698wy2tnHHW9JIOCQOXUBjuXFqvVvl
rCBCvo+GSr7njQzmopaN1Y88lCkW5EH+6n2aLWetDAcLnSZ4lkR7XGc8IrR3Rr/n
nNCV8Qg6K5WDGTs73GbjOgVW3+/5mwMdoJaTtxdohHnRuhvdUbegkchxuXNF5xCV
vU3VsYJcrIMhpvshEbJj0nwh58TPnvz0u0yQMGnnJaW/3UIsth2AohuQb4xO4H8O
i7xbkQQ8vScRmUQbkKuYKOpMid7DDdd9hHtghSx6/n3GePv5UK8uGmZqjz9Zvkqz
bBQ2091/ERL+E7DQ3VaRzvLC7aZY6m8FGXJNql7aeI5w8Cd9B/z8DhVbrmlSm+sG
xEQjgPpwDPZr5Pl4IVdP5ybFsjOPw353DhyDZokmm5OgUMWEiHuuYqSDPXC97RMq
279BkfyzwzNUi6Aja1+uNNakgCFeKeIBLq8iXxl3atHFkuqITB0vcO0v4ZHFFqVq
0D9C9WzKopZXW/QHcnWcEv1ImEYgnDNd4yVA2GVlvZzqKl7YCJVERA/wz1MpiH55
gmxRsjq5UWbn6dn3Ax7BVMaiuWaNY0W9eHExfRe12DpOiJxHcT7mbsIeKsDltE4e
CXGWsb0aOsKXueozLzhvKQ5OAiC8GyxKiepvRLgur30JCpFWEJU8+VhqZa6q6tnR
EeNc1N7bBS878Misu59iPDKQsbVnubgI0c1ek67bS6/fI6uxkPjOodHKLTiLqhW9
d/NfGWEi+4cXgBtSkAudY5GcqFiq4RKzkmU8q/v1yOEbjqZHJKNg/iUi5IebgfQ0
Dv3hB5s01kzG0Q35MuIsVoCqkaj1KIBtRKrfltGwPOdJh+etB8iX6nAU5TJonshV
7N2GDyt4/2EuUVDUWK77M/8fM35MJwXfGkkLzqhqjOj+dZNYyDbPGFIS3mIx/8h4
FPiGv88tslUSDn2GMUKL6p+uJP9b4p9kw2E1WYp5+eF9eqvwMtP+C0ntoEFmczk8
XAb1a6888lnYZfB3Z4JNU/CxLe8CJBoxCaLKQ66WfbFl9cyDp/cAHJN+T7GjSVka
HdzHbpdoFfP0LBZUOf88TJwcZnv2EX/TdUa5EDDJS+hfU4OiJB+VEClUqkaI4aWt
lTHsYDV5iv4UpWlo68O/n1sSQoDWoyToXjcBb7o2JJ2GQbD8eiXLjwvaMmIGP/+7
UVRfLWMafKbIStvR/6Mg8tSYzK9Fx4GAIME/l1tt8NJA7rtL62bLWvd3hio8gkyL
uW+wybRUpH6/h2JuC+VQE/oqz6/J/H1wnEwaH3MsWmM7UXdMNjZ+LF7r523xSwpm
NnhXw+UPjV+FOu3T3VYtYRw5og037XaMEuglYtZ1RL9DrfcwZlKP1OlQjhwWaNRw
AAXLtRO1NTeCSusGCH/Y6yjwTsJgdFCs5sGdouEfnpTHqnF/BlBoSfmUbYGdIPZN
iI8q/FhdFwp8NXiFtrTz7sk5l1WItQrQcmzqTwgNCU95epAVVd9Su49xAP0Jfmly
z9iw0NbHgNZ7I/IrMN04zWRErGmZb+YwrXY+I7EoF+hrpLPezyKkayI8EWkOgufW
T9Ya70uRptWB8O6BoHoYhxGB16909H8LA3sVe9Zlku2mcF+VLmPUzu+tE4pIBfMx
dyWoMa2PYi7niFvILbPTi/vXEToUqKNyfUFQ0/rMQ/JzNFaPywh+OM+YWfvXU9Jl
L73E1Uyx9pMRPZgLtJHiODWDeSOwAhmfZylfqiIprBNo3GgMXrJtk5xC7m7gJwIq
cM7NWxO7eWAc5bgeCob6Y7etQoSym0GvYYuGHi/o6d2tV9RYOx98upjMgfdZqNne
Ty5Bkf9hFnUzL4UJ/wZ+J5+CO658q9eVujigQbclBz/P1dBbah5YBd4ZnEbTrhqb
FW016WZrWizgWuTbbiHUcaa1I0SKM4XIUL96Kl2EExujczDT67f8GOE9ziwViBYR
/r0C5c+sPAF1tErkJJU2QvaxwBD8YuhUh0NOJr12mBgSU8fP1x4/wf1GUuKCR8RQ
Jb32o17g9dfgX3VhINLzXX5UFCp1oUXLYw9lPnqOkuzPWkiO8IthD0+jG+nssKlG
iNXV9zQUVq5MAFeHMgHH5xrDed+Rl0znlZg/3Otxig0nJeO5gsWR3QvQJ97WVVHW
Vc0cm3psDAPPurJmipXnBtkSrDgNKlz3Qx/IV0MtcJPRIbTtcw7HzaYP8QoFu/TL
YJeZ+SvhotLyMaEsecbc2mglSyzJBnW7juDaVV0CH62Ko3dDZPx9eyy2NhNOrWFD
mt1S97F659nTgMDAU1uQoAx11oKoC6ESGmyNtvWbYcVg2EJAG71GCKgAZP5go3Uj
73nKSu25C6vupej2MZsrskrsNCR3jf22RuLxus9zdB/J2C2LhtTwuXsb1t2XwxH1
NRuNlNnAeklZvHHVuUGaolkZ92fnyaAGk0pXWdgVMWsuEQkbllDjeRc8W0NpQ6lk
AZzk8HfhcM8+0ulLZSduJW9l3yNJg2lXa4Iuk40iP0+gPKnJn5DG3SAd0QPPIn/J
bimsT2wHzUGY8luRrA0iZmDKvGziYeRWwTaN+954j9GkoW/u0HzQ0f9GI7njRuYj
bSLE2Qj4DWT4IdRLuWBP8woeE0A7eshpVn4gjQhhDrjs7MWO/p+j8txl4H7eb72b
+lo+XWaDMB1Etr2UkF47edXEOmFBJ81h3PQfuCh5dM+eCAvN+EuNr9YulLG1n0Uy
4GA/1A50oUJoRRLo+uYqtyj20DlRnFI+lxDw1F12cAjDBcwhiK//qUWus3AHfU/k
khywdpqJqIkhkXqXbobSSmvnN2cMSwOZ+mUphlykvy0r36Bsni2B3qzEv7UQ4y+w
/DQfWm8IREj6yP3Zkh/fuxMPMCVqpBv2Ez8jV7vbtNXFs7HsjxMYsEJyl46aoycf
lHjYtxfXo/yZ+AweZLuzMBfWN6o0NLbVU7geiR0AIq1/cULUeS2Bf1eZtbNpikap
QIPstMDhLoEeh6UByG8oZWpemPw1V00RD5Nj+/tIT9ZAd5S25Vvbo0HfMCFA1uqm
ze85YgMlDt1BlqcHRzvUHkNjGRLKHCFlMu+QIlC+fckeLyyjZ5J6BLTKVYkWFD6V
iMZec+Gui6AXYrOpa1Bvfi7A1CLjR0dGiygnt8Jr97hAviJIPST7r1FHZx5A3v4Y
3UWN+5pZpjbkIQT6BbO4yiF+foW7Ctbnkbd1fCHwZ4qkUgUytjGK5INFAM5yZQru
yUdMlXVHXFgz+ZCIQMn21uSRG9qhuNpowMrUyxqdmkH6CxB5A8lAGVTP+roISppp
gmw1zC+SNHw/alPf7v5S289ROEQj4q+Ta0a5mgoZmwrUGBdAwANagq/I980jWIb8
JgeheVB48ZM+1lKPePLuENaTW5ghAPhqkUBGcCrkOFvETfHurqaH6p+n6hNRej5P
KKbJ+zyO6/hWEhNrvnmBDUZ2iopIVATxgFCHSOB+W2Q+r6G4hOL3PVtUEy3Bc1Zw
xJGIP9sZVyf3ThXjLIjO+TUmJ7t4gNgGAXo+6Ei3u23l8gn2yUWgAaXPaaYPNGhX
7GTaFMk4u0B2W8jy/NnpZx/4XzCq91/mi36NVpSHjp9XRYv8HNL7ACaJL3AhJJH/
UB+/KLRSewcqzQNX4reWX2/z2EwxUufS2MlhY0SbyHFGa90U0PMsOBeBEFooMwJg
6qdypOdttb2RUUKA1O5OsdXdO9bBpspwJp+xJwR8TihJaCv6eKLwUWqcOTX0rXpF
V/jvRS5+X9QuZEFSm65gHnt03ldN+0vjwnDrU92g6E2dDlme2hR3noC6LdZU0lOC
dG7WQ6QoBJcHmUUycq+Ir7QdE4cMNtGcmvMGvTr9zlpb9cDC5M6GRVzuPeOvCZOo
PM77g9hP4kccztEvr1wxRAjzrcMUrExa0QUDTx/ogzHTe+C0akkYEv1zYQe3iuSl
+j3+2aikyrmwLgRLCmG/ZF+BkbAEcfN19zU+JvHiYrKb3dupRCqriZGnhcWXtXih
8B+tGpviKk3BhOym3UtFoYiga+sSGwjv1MRcYdzuab0jwMmM38UWZhQnQ0gYY0CM
wXUdmddV9ZMzFvBoKLCuOLNgAYtiUsitB7rNvm49VgiSwUjs6pdXZ5M19bHtI76+
IQSDftmaPpRqGgP6Yl/eCMXDk+t7zQnjQ1SpMdja93ogo7cx7jwFEB/hRTRCEmtY
2Jol4BA973WrNw7agizf7AmH8iReDA5fn8dbspV4EG988QiwpIwhdKdnliQNs0Nq
1wNZK03VZdNVnGz2Qxv51IKjtUmvo0lih/n9GFEkM8ddtgilkHjepa+9MHfZAniz
VImydX+FOuDILgCosANqfqCFbs8nfR/WgxPTJEqDalkrBHEJQTtGqu4V3fah08IX
6vyZkdSIXxdzHw5SZidB9Ou+NTYt387LdTXDu8v1ibJ17pPb2oe74lIh4KIvi0f6
8fUfC9UYha8GB8xAf0L9m495hbCJW8FAA4s5ngJBruG0u8/Kep8a7edJS99N2fqU
CBAmZrv2Vmg4Tf2GoZKeqviwUs5OaHvhd8VgW4ZBxOYj334XUpV7Ws1gLPV8UelZ
/GcICwFmAmedwHF7m8pGtXQwhXvnuElyUJZvtpMUvyJUBzSzuRMsIIFN2kenDKhi
vySZBm6Xe9W5DHTWTeDQjoPBULcMw9fRfrwSqtBcpnqThBjUMyvxAnruU76cR3be
E6QPUAPPowQNiIO6+A1tb3TlxsvyaopVP5iy+dIKuA+3rZb8STHj/JwdLmDFSqkV
ZQ1CzJymcqtzjCjKha+gw5/SRAYrLsrlL9agTiKVydnIf1dwq2SEtOXZe5mL5dxA
hHmvT5xQMWqjs6jEOPSJzjGopRypJt9cv10OOoLa/C7dBnS+yWHPOw86JLJDQx8o
fS/kbx6Zx+cd21LqXV18figuGuO1Faf4wHz4cCeiQXN7TNGHshquQ4lRdRewv66/
RxsbBmEb3xP6meA0QYg+rb6veUjqoZqarBM1JQk5qvQJ8uHCfTJyWNP/21TOSw5E
vUXU00tG2NrdFgZR+9MenoTXX8F6f/3zbF3nt0rcYgWP8lxH/49S7Tk2E12jumu3
ajEcBsam+vypfJeF8QY5NPCG6wq1Eb33ld2hwex4weloDHJpNDNeKedYgztF5+Ln
qAxD2lKeclxmqVLSFNx9h/dKd/T9ntVnpz9/gIpuLThfZgEmnbLVhCbZKYmxk3sD
Q/KtHu0jqrrjbq+Tfbn9IkYSDpgQADjYbQxUiJejWgJQKLxbX3slWKyo5yJzls/N
INu80ygRrmnFxwSYmHeVN6R8xXXSplR/eMwX0fAt1SzNQMGS6qjibDM+U81DICoz
guq5pvFlIPFwLXXrtTGKEcRpTnpmN+lD00bGMKYwp4Hbv4RDkWKnPP639CkdSOQl
YOqk3+z/UX6GWweCn1SuKbHK4G301TA2L27t4rklkvCdljkO5DjJVwsgWGuEGVXM
Dc4BROGLebTlnvkM7yvzLpHPRJBRmWqjtYP13sJ3xe7gQ6wDX/R05HVAuKzVnGIT
VH9FLfiP3v9TUjlYBYwLHjb9enst0B9OoXXtx0lScz96QTs57XFECQlS5JTN8ZCT
T3T6ntzFoRwInaBd9w9VVSvPaOH5gI8aIQrXQNfHgEtQFvaa26PX/zuU8NSbYF5V
mwm4WuqTjcQA+wkB5Q6VjwXRUaOIOKkHGie8yUyDm75qU8+GahN3lGq/xYInq/u8
zQhLuZOe0qWDzddamuOx7lHKcz2KN4SEe476efH0wXVqgzsQKxVmIbQJjhVu8tnw
a5bb3yA0gDZYTBdzxjXIZl9VHslm1wEXO34APupkP9YO6cD/7p32/hVOhw7E5/+W
SNFGdZ1mXl9ONlZA85nHidLJ7Ks8uVOsGBH/r8CzX43ULVpqmfcEgxmJ8jZ6/MQe
iSLN6CjM48+kUbGXdRrWI1hebOyfR1d2Yam4rXaBOCgFg5uqKPyYAiTm1YcR+Uno
HV8f4/KlS0+Nfc2CXDFZ6mdK4UwOsV1leujZQT9xNLy3Sn5GGg377iW5AmvQCuVf
HN5B3zcdaExLAnXV/UP9G5eoyYjBGw2f+9RiWdlHdwCfrdoH4WOBgNV8umC0o4Pm
5tX/K09kKGTys2FT5VtdUHsPbUY4wI+v3yPSAUaydU7Zb0eIRVYudAvGINFWOwzQ
VOMwj3BuERF4CdHHjrYmbTe66eFLFpbXB/nihluAOQbHot8EFuHyniyw1WXaRfr/
F09hwgMaAJrO5Lh1N16xqbmPck9Yz/nf1RI+GFFZGbRohgy6IJabRPta48qgayuR
Kw3x2ZDQiosbTXsmgfJC1yA998FrQPya4WGdlw18ttiV/XftZUsQOvf4byJMWoXT
q0v3XY2HCf9t9b1lhNb+iOJKkNKZQidxafdYBhVZZyD/4wdC6M91766q2GQ83ccJ
Wdrh2VvLCVrowCVJEVLJou0veHABA1h0Mf9qVp6gIWGmBcRkU9QvXnJwmllTiywI
Hr2mnTyu9ZzagsXSpiOwHa+Vlpzg0YMbPhjsAqr8viIVvLhHTckEJv2BDBWJSMgj
DVhCoY61uLTnN6UtpawAjEnVsIHiedThBN8yU9ed3V+Rw8YExUghI1p3LBmQ6hxS
8AEcPTF3CutcRHACxo1GwdyRWRApOPb8dErwqHEsT4x/F/GCOxkl4dOkx79TTIdb
agpasGdNDGTycUo+G7ojAneNrOLxrFg94DnOzm1CP9POw07c06x3iKBtkOUH9Hia
iTMlGrjd3p/FgrmlczQPOgYZ/EVufgjvyJuVvUZK2PSaEF5PGCZDoJ6VzHZHwcYY
EEya+jBkb6IymUf8ujdmGBklC5dnz01oI76n9qxhUmoAmtPi9GqfU458yj9YsRHD
RAN35bk0c1Xu+vfHoAPZZH8MCgY/A+mlco9cK6YIpNVXyfuguqD6PMNyRP5Sb/QM
y21B/MTtKOike3EqnQ4iyDFQ+E44HM9+tY7YA6kW8BKGsx03FXOOU9w9wEXi26xl
HeCtjPfGpZ830hcIOqUmd2Wt9kL1ElRYQOCPmS+0RHDxWQmcNjLJUR1PILnYQrcv
UihU5SJ3/XnhKLmQFvSvjM52F2mkDPUVXn+DW0Rgf956D1MDn5tSA8LEC7YOp8Tj
VZgzYQ/6cQS4NuQYBv89e1HsSN7XI7As5D38ogirnfEcj7UFuN19GKEdnRnlTtQh
1xyBqtTsfdmOAVwxYIyqdNCgi7CJ2clVMb3HsuUCk3Jw4YnVPV19YexaaQhmsVwG
H4IELiD2uYVVtnNRG2ZKDq1CDCtv3ynkBmFDB7gz2P34pLvwecPMQDfzlQwtnAZH
Xi02oL07awkjnYZMbDO3Z1UPvljNN5LWJhhQ0JQd+M48Jp+3QWNL8K6l5BIT8XgY
aA9aGUWhAInRCjWC5mjhZAMJZnTc15VNXCWY9tFuGPK3M+vGXM3wOpGoQUwRge0G
q8jTq0S06/pmqM9ltyhT5E/M8pBd2KIZq5NiCTizghzRXjKPj3R7HH1Ghi1mQgLw
Ua3uYAet815g1W2b9RA8Ha9JI8tQ9cHlwoeuUmh0Hq+rOjEJcfzThjrSeDW+oVNb
iPn8nOtPBN5TX7IpK6zvM4toWf+l6jrMI6qjbwv31Q18PUeu+2pcwUwT0LSW5yBb
vJq2L3iy7zCniTKayIho8fM17Y+I/k7HcPoUYtAhTmF9OpS3QMhlJaFPxjhXof+4
Brlu4jtFKSo3OoyA4IcKqkhyfasl8hv5DUyQlAz/g5AYYhTfEuUU9Or91VbfmK+D
wQK4rHkchOG8yqWaquw3iB0Sx/UyNQj9+IIlXD7cmla12EOPYbQQD+I+01nlYgsP
To6rAFPoOxLkh3TbXCy0xlkfE+5BFXiVhyl9KWxDw2ssAaU8zePT/DmuEmSw9RBk
RPv+mH09DW3fUM4kmC+fbQhSG6lz9hNzy0H9fHIC9s5OsGpg99W4R4UVEwvpyuQQ
8isZO/gUDj8kN0JxggAJkYzUxo1od7kdFJn+B6tZRDEfaWVjDUbeDxbvlCusAlYS
Q5Ao7CvsZwgEOuryyaEilfZzO280jYboOOYmcbOTJXiIbCTs4ls9GGJa1laXCs3z
ThKWvDCRbzl5ChbSfQh2YSsCRo5KnUj3rrLF16BI9xtOLiZLFMfjJDPzTmjlznA4
Zaq76BKjG3V5Vu/xbaq0Hc2nE8/w8YyrWyZbjrx1DYDOUmAmgApPb7SVfdf/CbPU
63TpGjuI4h5CDFFDfQ6qOcLoFylQ/CtCF20PlNuXeiHQ3iC9/3LsYPs6O9axwZcG
BSc1KhHvSMwvs4+WkGWzwrrhy//v4Ht9JSKSxSWvU2Jv2yRIiOuvNUs2hP+UPBdF
so21b0MLbD0hPLHMkAQdpLBPF/5bbd1XHiXHEGM8TOyJT0qu/s2JbEc6pyAD8Zar
OojX7tHKiOJ8YbofnkHjMQ1p0u6dsIiqSgJIPGJe0U36G5egtt/05fpzFhQy5B7i
a0BEG+GJXn62Eusn+8uzuXiFp5QgpWDs/AlXKC3mmiBwIwocEyCodN1/Bh9ks+im
wuV252rh6Ox7qbfZT8cVyJ+zls3Cao7/DQLpBMxY1cAunGqTqomqLVVFQKvLe7ED
FIieSCADZdWO+yzfcE7P+03kecGgViUGKd6/NWd42r8BrLlDw/DNx6tYxpBNMf0N
iauLKbX6/mLf45ThwK6QDHMXRP7nwzSIEZvthythAibTHqBdUpyiixQEPMQfy8Y6
aSkJ2LvpQ6+NDJ4Lr9O6nFvkx5nG73buNReDmWjPfA6cW4R+zq23LXcUw8Docdfv
B0k4dFl+JsjAr2vRWJ3kr3yLv8FnMzDFi0eLo85GHH5cEjZfM6EqyfMsaX0UHpK1
pfh+bc0jd97k78udQuwbY4SGuNrNdLT2YvpSa69L7dkYC/0ezFfDhlTc3HnajEUS
+FBXrzbklw/zEc+tv0y2dU+NodyC4HxB7qBXU6tUYA/GKUrSxLCyoX9AM8dbqXpA
uYjXpGnU0uECm+FBmgIcCMHV/nnCD//uQTz1vSkNy2IxQhBHjkprRKUb8WSHWnwO
jN1X4qDv9BKmkgIlHcgdAprnakTYrqb+L+U62Dz0NVl3nTgz5nXbZayb4/TSHcNW
+mM2ZCVuUq8xEkiUR81CIb5n16bFmjkyCStRNqfH4Aa3Gyf2YOsP5vbO1uNUp2Vi
UJHhZmMAYHXNBqxad3wjtaJbbztLt5ql1nk1HeLCkASg3Yt9ojKE0myOjufIf0Lp
+Jo9Al+1k7/HM50x+7kWhxCbh7RrrUHVNTmqFgEfp4bsyigKvbQYJEbacvm7lB8u
b82jQUHBl5i84PQbjKos9FjEdV1q9HQc5RRr8Ic1a78XKYfqdsv5xTqP9yhFy7f+
dYIwr7I5Ij0jMm6jzph7KsbrMN43v3tcBnl5HU1krit9xFta8oTFk7D0ICLIgfzt
Ar3CTJM8rqVyFsQJFrUEhNnvIyAtKksJx0NWo5YHJXQO0aTk9vrWv3K4DOoKTvYl
MZpYFXmVqPbT9Rk2i/js8LVkM4JDyJdJ3OBQr3oQ2ahzy2B2UlFMt+NewviHHeW/
wRifS/BB+NVf3zUAYmTSIw3M5kZdTqc7BvoVxwRDkvS4/AiD3XPlVuNndLz2bkYf
oYgMHonRSXqNicTwHYs++LBxUGfQ04OQ+RNKhpGxzCAfATDD/3GtCApa1I5mE2Tk
UYOSjupTtsJjaKHHXPqnLpT9ZTxEE5NGESEy+3aPCRijqi+oO/sVg9nRwRK9SHqe
XWj6FRXxb7kBU06r2QzidEDTf7ka73bddVdWVhFneprc3Tn+3HLTieagRSPc6+6I
UqLtBIt481Cr+KNVkJJIBLmHsFCDdIk2q+gIkys8Fxyym9N25LtRofNUIodo3ihD
/PEwhyy0mgMwdt+mWJ5qgu//+sINU6m55PXCVv8WlP8taqD2FVlW8RHdFn7qA8Ba
WEnC02msX1VNiK8wvhpUyo75bSXB96O3N1nDmHsSjS1A5nK9MpR/0vRDn+Ldgbww
5L+l24jvWf4HIfLSADqSNhEfoIUZ7o7qGn5cYjua5y8+v1QsFiBiG+e6TccAOewz
dyEa60e1tAfJl8qnUlZkjljNG4o1eonPaxFLx/XBLZAHxCYLr9TR13N54ES7RNNR
zYFmz8B9ahrbZkxl3L4HNyWDVJE6RtpYJmXiDPc6WOaOuNd/jiL9U7ON10KvKwa8
nDseEugkqnPuJ3UzYGk1y4djYXJHgeMBrwbVLY4laKPktTjORItSX48Gx16EYJYN
HuuTVQw/0kUpI3zVhv0Fk9RViCHyfnpvUWEmVIEsMldPwzZicd5HBNJnlb0J6jgw
N7sYuUFCh6rx/Yl7//C5VAhawOYp5nvWQM9+eJIW5c/bpeOCxoZVArxS5YnQTh1M
Ws4ZuMRg+2NztO6Y5dNw7zXvth6Uabu5BZPr5nhJpaHiekYf1beAqm8Hzh8nbwd/
M/KyD2tzmC/toT2WkSD9V1lcegiE+ZSvKPDnwQuxDDLRbmzsX21AjZqV0oO9VBdC
FAWaYo6Q9KsBgSU9q0A7NAjg9U6Aw38e3CwoqnPfj3yqXwd74SpJDgIiMx50Ea+5
d0oc/kxGWl5z+suIjiRaBOXd7Bu0UiYVWv4M1MXeW3/SCFv47MLlkcowt8Dcnt10
z3JRsWeBW5tN53qjZ2CUG9OsbrGkkGJ06pJtVLs/CNZaAvpDKmWfPeLNM5X9KBq2
RXCzFL5miekYaBPnyMUbx1c9ZejSTQe5mpSujQWhh11J0s/Z+IV2W/qGUullr+Xz
4CxizZ8VQ8SsreastmyG0T7szZOPOthIuR3lVsbOXLG5SC3bswIZkmHpZn2d8w5V
yNdHsqBj0ZcoI2IcJbNA6V23uwhchtjM1XBn4a8nVdVbX7sChwQIWDq2477G58GY
LTeD1cJ5a7+iR32jHJ6xYsu4BnmG/WFmQDdL+egMdI7XTvsk1cFE30H3gJeypt2a
cD1jdBCBbXgky0OzKV6knTGvWFbVARrTr3EfJnqgzAviLcNk88JZHXx/yaf24WS2
nFbLeVkw5bgpqEUcCW2WHGTVst+GsywWzZZY4lBqI4h5FP2pR/PQazpYi4Xg3FrQ
nPhNzxrnAZCzJHy3NgIu9AexCK/aK2S3rXsYOH0LOXc5PN3ZpKHcSzPk2zVLusZI
OHXkJoc0kCOo5OiGcsvc2Q6Tc3t+lN/Hp2Wog9GnSXsWeeGui+Y2T+Nw+mqmqC+b
19gVbxlMA6uQWagw76JfOBdo/3je/CE6Rp53MBxbR0INg5Mlp0GUz/4q4uvz6fR8
+2WM7xkEK3GuhLUyAaE9p7+iz2BzbxHDm0WufI+5YaG8XuYf96aVqqE+f8UJxNCW
Zcov3wFr7cLa+JmeyPL9i7h7jCzpR+ZLvj3OZDTuHLIEJPluo4FkVrVNT3vCjtRL
JlA+EJaC70tSmrqyEdrhBMB+rxbGwQRaKZQu5GQc6I/OwBbofUNXv4ug9QhI44a3
OX2UxuusWvNIEPtfvrJ6EJCwnwGq9mGLl8cEgDBdFgvD/j7NTQUv3FUP6kbv6wNR
0+wl6d2Zz9baUjrqFBGxj9//dlx4UegyrMCkxC1I0j/IaD9gz24nsFMvz09NBoe9
rYqnejEHFrL12nGu6RAfqO1bY3eyaaoBCUSU16czxmigkLnSXYIv7fd4KEr/tf2X
PrnHrq8ziugMNtl0SQPVrgkHXGhZCIQgxQeuAqJxFsyV0gQXwfr7E+nisfE69QNe
qc0h2cd//bXM9BTavBvDF0PbLePvFv7/5jex8/u28Wc4jpWqOCWmz6cXZJ7FeOGx
9hgl45uaS3somTvHOalE1kKTbjLYlb1SozuSbHcvE62v+FcRU3c6GaFcVorGkOSM
BP78Zpvfkka2jQVUGjUXup+6eEWLCUjYezl8dPuVgia/s09D1YvviJ5rV1xgZid/
P07LwiI1ifFnPvpSKqNB+vm8K2300TEvZVPOTi2cuMwN4ZHwwPJ2yXzhYVEU5xBa
CJsxW5HieA2RJEl+u3VUFKrzqbbCOGNQjDQsFk4ryuwKsdAuj03ZpM1BjP1fkzFV
/zpdYVlKdN9ra8TQ5lHnwQ0FokIywUhKlh4xy7rj2dYD8Xmv/G5aXyPMPUZDHbWI
U+QyaHmDSuswQ9JLv74huKD8dxc5kNIX/4D6JNpO9fEbZPfRjpZLrqc86DNoEhNt
By6WpT2EWItjdfrau0XS0IZG0mIjn8FOlWhNIJCEAJVLvEBEEd6KB6kICUELfCql
fJcbakFUMMgh/GEldbNqVqAz6RA9P4c8qU9hnH4XO8OfAQ+rCKZve6YIfgROuo7x
iw8kTBFYx0FJL875MWBC+hZBjJCHE4XVu9VbVLSkudXStP5pjFH58/apPBkZ49KJ
wuSaEgmrAYb4mTng35cxTnEyW6BoUP0gdqaKs1eQfRvgdYBlSywAgE46RbLrLHgR
LSl0iB4TAwWdvLZO+1wQBJ5RvowkmLLDHWPAUM2LTbec2e0hg2tHs8RkPodbinfH
DHqwjYjhKyTaC7VR1stOtoaxaQeBb271QUkPrT8TqgGnJ7mJ4TmPiuMEPVdprGfW
pUmHk8d7dzE4Rhq/0NdvNjd66gOuC1pbg9Cp6gz+f0tvZYgEzndC+K9GNaEUfCWO
yQFuMt1HWPyKnIRiJnx+ZTSJk3Hsa1c5tQFla2r0nW1yYxqibqb/CANCoM/THUjt
TC+N47jxdp4kL/gFrzlvcw0Tn5KgVJ4euvqPrVM0+cMWd2GyVmqP3Cl4uPF1zbPq
3IieUwoLC4V8jnZbpJRd4wbHnsvQdiA0yi59JGfDPgBpIsWcdqW7M1LntX9wTone
1zzizRFuOkapp1nkW3PppdzCLvuv1e3E4dlJq85Ojwx89DJRBMg0V8dzgn1FDUdA
G81QA3gDmtZQK1LLoWw5rCbrWD4VNWLATCT/ZqsM46PyKtLdUMRabQ3AyrC0PAdc
KsDEGC7K+MrwOkqe4yZYOd3gO+/dJlDDSsJdiIpRUDPFW+127q6v9sY1SRHvJZ1r
5FilRBV3OjjIV4VrnhT5wHJp2kHx4qAxFr8V3kxKQ93LPOghczutiqXxIOCmxVnI
aCnSkFizpZoHMbiw7JNtyGuMVUFE4kXpLsl7qfGARc6alZLJ1AVZ9mp3AmQCQnT0
n8zCgt55QNF06UaGskykTYlRWFjtviL9iWoV7smn2YOnuF0EF2NII8E5U6yyIhu9
QCYICIwLszIc9jeAETx7PsNf7ZQe/aWIWs5r8lkF18wuaznJyi+hgXmplTYh3Emy
EeiT1ykcg3s8GTfwKoFwteb4FyAc3v+LCmy8iNXM/P26HsHLx1n5X9PX6jB19Ym6
6lyLACRXIFJE5wBctKdvns/wu0KhobIJHjU21e9IZ1bAkYEsQejihv5AQds0aYOT
SVltnNdPIRea1Vwt8vVqS9IDLyqpn9I5VQlaR5F7y5+eJizKTjGdVGIqbecrkq+H
GpxLu+GbzquO3qyRAQp+mFUZgjR53mmd+4Y8vGUqFQvdJSjdzX0waFVVMeiM9dtW
p0yyxjKeRYc7eWBWKxGWxOdE2aOKpHGmdYbsNiio3VNihaoXLbGJfs8z9YEvKA/i
2v3ZHtHyojsyAfkFqbSKyub1DO0586qnndgcvyjljETqPGdXH2PRWcIeJ5n+tjqB
y2206fBb5WlQlKk30XlnnbwfqHTqoIvrHoT+4Hn8CHDuIestw/YVEjbReRmF6r95
kv9DdHC6HucgSvbcx1yr8pxxjVFg0QdFf2YZVsKvTHed0KjZlBTlMH1KNb82hPns
oDSkm1NnPwBvHuPYEpwNWKab3jB0CaztsYwcFARbQpz3eB6NtorOpQ6DTF5hJULX
6fTxcyTVMl9NLpZhxHBv63G1I1tzP5Cy+7pMKKF7C4rnxL4Hporod+4vejoOzA6G
JZ2MSTye/xejOVJ6fdaYyML9SHVXr6GOQovrPc++R8Tjmd1lVEfjoZESY89KruPp
7vG9nLhE97mZQj6SkkjgcAn8s0hmIutN4687CwMAVTGNtqvkPSLYYZB/UktJ6NKA
BHSeyBJHWwkLYN/ltEx3Ilxico5TwX7/PApY4jkyoPTjQ3b6zC0aLAPYfm3mbwim
B+ZB2CpAkfNeZKDupD/x82P2DE62QHljjKOMxHMRRKmiYsaUEIf5pjY/g4hvgU6j
jh560pNw+nMjIdLHx3VAs3gwvGwhRs5CbG7Hc2BKlBb5UOR3vS1ITyj7Gv9N/eGR
GBTizkRn3PpiB7ym+EID8yCXlLoudu0qPtQ5/c5Gu+cPu30SKP++pBHb43taXpkj
kwOWBP56KOFE0M+yp4bFGF/X3tGqfgHsDATqGIL5NL6RIMdHZxua5CY3l+t4sLiS
eNC2I1Ouwl+njumVcUulnpFpZoZnPVcr21NjfFyj5mGdIa1PLKx6DLcYgvpzSA93
EGztNNriJZ+5/GEOBJ5sF1WLC0Ywc2+49yttFqXt//7ECY754tW688LyagAyVfTE
7uTqYEGWC+8GkiE+aOrdS3FXtrDAYo9cq2T7CnX94TqbcrVxwwXDyfFRqKurMDkO
Vwv5UPWgLKO75AORrkIdbE/Tig8njrDbqTSZgWZshr4wB2zmmR29qEayFXivPxcm
HzxQWLefb1Thr/G1BVe0Bifdq/n8grZoXFneMUMP4ozYCwYuy5MAb5Uc2JGbeagQ
Jnnxj/0DAOutePqtRe7SxZ5D8D4tHswKpGekS5quRmrvyQJwCfpPBJ3WgdTx3+12
JQLnDiYzX+XGkkyuytCXYKWp0O9TJpw+ETknkkmbN2Dy7oGwv9P5W6Lqs98McIS6
VwX+gKyK7EfSl6tcuZapfin7IOB1jl29u5S73dhj4PTTOIt6Qlc5+AAdrDYVn4Gr
bcbVDeCUivaZatqSisDoloAOr4UitTfQPHaZdPPAc0XnkzFJdDDItjd92TZdhDi0
60+Yz/K/o29NkkVun3juVmIe7CY3+DigeqouX2s2GWb0MmiiLQ0MzOZqj40Z9ejC
bm5wHKmbEOgBwNrNaY3GMMYWBckYAN+4B5RSRGpsJj4oE51cbNLjxHd3vuitbLGQ
715hr9tpGX6B3xliIiajPIhfUhfAxHsdo3RtqgAJKw8ckCT4YEAcRosYt3TEQtzK
eIMqSanHHGUn5nP5ztxW+hzT+AMPvMA+SDUALlKYzCe/gIPQpggc4/6DYDmqgUsc
l3OV2ybLhIA6LU6hh+/GfYIFrNbyhzCvdCkCj0LkkZJrf1NeQrDuvumJ1oUOKIeR
JKi0Z+wdN1imzsBCcQFfL7nG5Ja7+gEJqTNR4cElJOMjrWyjUOysj3Div34OHGQH
nxNHk5NJQxoHw+0r9I8IOHrkDBl5EvFJ+GmUpmQ/aUEqmdQQpvN4xYhI9LfZpzRV
4H1LVLNmU1tutzUPoYymB0GPgdyZgsrqNRzDWO+oobkswuZgF4wokFtZE5xdRLWN
/uMIjCsezUVebT1hb4X/0/p7ADLDB7tkGneAkpfJY9BFr03oijWldxabhf3LDkiK
JQVYqtImdcsLkgOuxJFUVOzdrSL7a9F5TxpWyIREEocLjmnOeGrPAnvQVQ7YCNQU
bpck2SPRNNVY5SDGKunTtnl7mNKSrGnB7sIQYHaCuqVEX0Rl5jtv6TqitSApW0X2
wHD5ELd0NXnt/k0X1eKt5QSa/w1m345kBdYbc5u23ZCKA819OeRP3fmBbLqded/A
CP49xztXXdIl31CzMO5Xv6Ddz9UfuPmIerRHJT8xSH0i4u5V+KQx2kxOu0dE3zR+
jqRbl7ivl5EveKbcylMS/qjCRjPwt8/obTFSU0pEyWjKRZaiTX2QOas/0DMmdwwo
Gs/SSMQIcP4mdo5tkRzPE3a4g1bDmM+6Y6X/oEheBq2ls+r7YAT6A+c5+QMIjqhG
vX4+CreJElvO5QOq6lFa1JtKedoDDjwNmp7jDJg28N3Rfe/UuZdPuADe2MvFs4J7
K8j3zE5e+qF5z+Ha6iPeo3Krr+KMOlnHnxDAfcIIzu3IjHzo1bGGeuQOqE8HJ9sq
+YwxSo3ir5kh4xch43DxheMYDRje48rl4jP/tldkt1WitZfMIqdUpErfxQTVsKUB
LPGnrAhLrpk5Pw/ZvcMYcZMRSqW8NwzVB0hWguzXCtiTuP4HeCDQdBajwsGJTqH6
9AI/QfoELlFxR9Jm1VWKUwr6hN/En9m8off5ACTVLfpEQ5m9St5jNbI60FA9Ei+I
6/Vq0eICacvuy9ZIlwNyotoiHOWUj0BC0W35l5bJOriQMWkuiQ8ID32dagAkAi0k
WEpsjM2wcBVZweNLlKz46idY2wlIE6qyUIwpEgG528drIASlratpti1NyCoEAzFG
GBdYMiaE5q1VuPbUUcuF9GEFlNYBm97XG/xicRG+Kb3RZZGQxlyQ/G1B2J1IJJQI
FYEdvEqw++KShSAVu4YZvreY7fM9EnRTDUnwNVPlGENV8eMNLZyvxC7V1uZvckKB
PNjd37hxHKY56vvOOmv38mVVIYFwWlay7UouBT1SYQWRjq8G0RveH7Wz41O03K5S
pb9K2r8BdPq9XSoizuLKA/CXu6CjuDEqrGZofHrDyKBje9kcjqY8JqEj8gr4Zb50
2pdpYNeh0NzaNY70/c0sdlAYmet657QdrCy+JtqRRikzMcAB4Eqw+bxJE8Yq7fZW
ZQ5BwuRXjyuT7AoxucGowvWDABR3TE1YEI34bW6mXMRNYzGbyO0DUbhQYgivzIcg
ZLThXG9VRzavgFyTwBF6G5Tw2lmiE31An+XPnproQf7Ryyjj6gbkfg8ZmfedDz4v
kfUheWd0lxebxrxOIAScFDCj/j1YLkW+N4aISkoISIlWFnfxg20emWxKB04rehIe
IJc3mFd2cZPznpkHWQegMb1S4VJgsglG+xxjf/Y1Qvv3AjE0E1mjf8IyrbugRDUp
ZsptRM35XFxo8L1aABGw11+bdoA+i6fKzUzhMuihnVNp7aUdX1qMo1Rb0sFJ0NUt
Jf1d5lRHbp/YrvBLJL9Czf+yhAYGLouIV9YKqor1Q+4XwDzglJoq/mLck1qrF/Rm
071vbrvBrZp1/Ge2MrCo4+0Qv0YNQipunwqIIsskGTtMv4Ie+zjHLOx2+r2shJdy
V5RwtMdCJLNyULyHz1or94tqmVO12aH9Xn/nVVVy5zCdiu/oK4o6lRs5ZpwnHpX2
2Zx8EUKMd+apQRtNwBDdPo7KkDijKSapyY5r+VtIqCOYlRUJEpU31R+xej6H4hUr
GCDyzwctnvovOZV7+v6iY7Yn1bziVihuUKjL+gCTAP3CiE3QhBn3DMWmou6s8kNk
rV4kfxfq/VIf+MuNc/6okpwphchckoWmDtWctrJyz98frNhQd/YcIT8b3oi7b8ks
U1jRu+zKoEQoV5oi8Bi4NBbtcZy0BPLD5UMV5F8uip6My37giNVgNtL/AgXPUPm5
vUsQ7LdPkkGSBVXzt6Zt7SlXJu13gHq9Heqn9AsVaGcismgp08j66pDQBonlbINX
ICiFkrP2ZOe/GuS1Ha3Z3+MNzFy4OPQpmXJnyngEpGfV6Pfh6PE9xETCmx2h09rJ
bpsN/+jp9DoKWd73XLE1Y9W+iexmvGRidIc2Bg2DK7p4T/5kfCOU6lYF0dUXgPAU
zJuAQV/nVVmGNyP9xH5y/rvrBKHd4+HoS2o4Wm+MwxVqrY5zXYNzyrfm1XBcg85Y
6eq+jyTKS1Kuge2oq4nG4sxhzpJ0eXrTuXMT/ZdR2k+1utIasoOuSVl+bjG3Fmgr
AciCN/Qs6efgzeGBBivYL2P4GKn4xaaa66CmT4qK/h3YtNRTU2Ul/TAn0jOS3IY3
7osAB4yhHYIOmY0Eqv5XI8tiHV79TNclWtjpfZQxpWa3xQJx4rTqeqADZI3RgqoI
XNG/iMF8n2MDMAOts493oawaXjnZEKpWHNd7vJouOBpYh7Ls/eJ2elK+J+cTPkd2
+5XzYbM+P6YK0tY0Sd8CZAr9piuoiK5R8DarV1a7fnWdjmeJeY7Is2OTn7xvUyUJ
KgaKv6xpArcPPW6JaTFHV3WrSeCnpg4BVQAfViNai+Rxvvq0MiuvHyf/EwFOgoAy
iZjmJO/rQH9xyFOnsZqTJBAhT359IJGhU8LlYZihvjQnm120yeZ7bmNE5C970aY7
fhBZsVetAiWqoUTfiE3bldoGV8fGcst7CKgq1nsbTBndF1tsVW5eOdVTGE67rZ0T
0d7h+M6cz2HUL/NyaiJDRno2YJCx/YF9o0xK6iufUv3GycXpzS1r+YedWJD6BIjZ
FYYeHWAR1LCIcMGy9cZyEkGgxgG4gRty6KB7A6pcQDDGqbYWsgVPASSOONnKMwYe
dm6/fjCkjpvgbGVbXSJYXOR1m9d/FWLDwFTW0AHb0DQEHnJe16zcuoTIO1846fEa
Y08kj3dytJj8ZHldPSpj2VndX1uhpHfkLmYo6YS74EM1iUy2Sy4bJuu/yiWFNPyd
YHsQnVXLcMgwO8/nbsY2uUCjkrZY1N2S54UA+kEpsA/Zz6f7iDVX5IQq7ZwYhUd6
0+MxgBWDi177gY5cPa3T25p7y8/a44S4HbSPC1dvDKtD9NN9iekdxTayKtVh44C2
DHgNN8Y9ooyuywR/gnsuuF4ozvDdUyzN/QK3c94Qtm2e0tSGR7MdPHzSzokp013A
1fzfW612Nc2Sog+/TFFJq3Kr/lDFrN/hHShNiEL56gdHFR4/Kt479r5ZAfiqRbbU
mVwftx24w6mc01bxxspdz7IEbhTXmSkrvEuHajw2PNy697VCXWqQtTS4jdx/koXI
3eIAC6d7LmE5s0XFFDaqhFU/ZYHNrTd0x11aFWTbsTsuT+hNgorMZYJYyY9AUOrB
YcFkSvO/p8Ex7rh+5PogbXzTMowKtGjpkBVDd9Tcna0KwUmIZfMlRblF7TgZNKGM
QJVnmMbnxlEJH6VDGmrrDtpyxHkwRANgBH9O+T1e9WY6NguD38+lDr8LCzKZETf6
7Z5trB8JoIB7Fa2iBW8nT9AdvPJlfKXehGKZopLUCnzzBY/cX2kTe7dN2uIKN/2d
PukJT1EsfbgWR+Eo2zoW4Brif833YwsDdoT71Inmx0aPz6hO4DefDLnQpC42PKKT
54OhQGNHd+1y7qbQM7n0aFFU21DG6fzGZCSlj5WJDfqWPvhY8n5XVXQW1KFNAfy1
H3dL7TubPYyMRxNdhcBpHIuxf+O4LnEPcYvIrYVy18CCihdBirT4X9/t0X6W1jGI
NyC6ixPUW0MxlxPT96cwRSXjbQ6w1wtcnikRq6FOa9n8g50OTasXtodbmJPxdTrS
+jAPl2kaBXlleRv42TUzgUXCyhAe1rNyI3oYfspw7QmJN0pdlnXexeRxyLiYeJjE
+JBk8Gu4KqG72YruhKL5ldHtMTlILyRUKZz6Y6gImgVDEzoY/noVKo7uB2JIWugb
KobUjjODwpPOK+2HCe5G7XyFhN7P+wDwXFqCKBsvwURdF3mRUBT9OUZzlyH7YlrC
7gqFsinRiNG8F7khi29ACnvmp76HzTqC4llHnm4GFU+iPRffutQB99waZlcDbtrg
gLD+v8BBV6NvJCU7RFLGaXhYvsVlERByRD9dqKTSuhM4bGIOEZLpWwRZjMWWhjze
wE+lzx/N5w1CwBQMcsH7YN6ogjiRWkqQl8Bf1cxL/C2jmeQ4fOu+Ys+hb5yTxyzq
386Ml0PG+GL92VtO7KOPHo9+eBfAH/y73E/mm2Vk+IcUQB/3oThxEUQt7rCYxouH
H6AgNPeMvfaqM89YOnaHsZ2JVNcqCo9Wow7f+LZ4HpwSUts9C9i63LdJNyXzisIb
rqKEq3qQPLwQwXalX8yU6M436BNOOt2Io83S/bNB54lXJ3vMMXBdmZSgjWSFbhwe
BF3UKXPdm4zw1GVa8le7iLHW4hWvVMQlJ5+1slubTOdy2nwqkNXgbdTQ2vx+CkA9
hec6P8BMT5UWcUafSu1OPbdSciXouO/FdH0OVylmmCr242lYB4hhPU4USDSI2VPz
3SMQ1z2t84EjV8aZzialI1kbOscZXaGgushdsb36xWspz165v0s3rvM3nEcgfD0I
S0Q7mTkybtg9aw51bM9F46HeJec2s1qPzW0ZIdTRRx/nK+/ilU8lt1t0AXgeCLOp
XpZIc+8hbi6G8kgLQWtZOXismUSvTxVFXTLiNZ/vAaWrL0cWIkMIaUGMBqBBppjG
Wi7u4YRGonhA9bCMa231N4y0fkPiuRylBcVG/crO3LIgvjHUZtkjuUW6ZfoddUoO
8EONylTgKdocArWc/+yC4QZHieYx8v1N1LmMCuiFc29QPTO+kEhhSCIRX7FPRYSo
sMfkiDbkl0Irky/9NXdrMn2YdpZivqAEft9kslQiQZAIpacd8pVgEcVQV1ErJLwX
WAsIY91fw9waIbhH69sFALGF0OH7odcJB8/B90uUp686T6RoBDQddMjgeJkAoOrW
EkzcwJO/uWcKEZknOqcXDBbthLd5pc+khYa2pmcyl4DrxZm5YPpBGiUZaqXDRhJp
BSuaKRssvfM+2dJ7RhRohZVur/NNbL2kG/DpEHC1QKaJnjAa7M2OhyXX3Qz2+xZg
I+5lgXg8lf6zNr3jRj8D87GywrGa7SKKp08sFKq2TFXgHvClNB/5OxRDtdvsaVdT
LTHUmB9LjWheFzUerEch3DRWquzZq13X7ML3DhWruC1hDglsEI5DhWgHh+uMh4lN
OFEtY2/ttbJYuJpva3Qv/fHygYGc/TeM/vrCAHUklWhGay6Tl5Lrm7BAeoPi9bs+
0SIvPJ4yZHO4okLdpkRVu3x/7dkxyDyIeyw3fg8TXUW1ZJNFfzPLyYxnHpdsbUE/
Zva5VPEgRYSzijdVrrJl6irY9hhKok0LXEHs3SoGl+d65V0YJlYeqhkqPSO0zKD/
hMqhzdgUvA44dPvIUkm8Xi51sxb26Pl7n/EcL0Fr4eXUGTVLDP64jrfowVyF8cD4
xLIyzQCm3SwcEcgNHdQeyBNaJlePiSNCsUGTYXdnM8s0bweN4eO5zX1PCsx3SkZj
9GCLyKiIIw/iixdCiycZBaZjvlNZBejJj0ZN3JCO9EEVYGAeZyyPiCFJ3aXR6Gh8
Uj2YExdc6v5QPZzkXB9WLWAM2+UBO4pn3m6oZ/0dnxm3LmyTCKs9fcjc6zySOx8+
G0hJjkBB2pdXsLyvEYjtgkPe0X8jwXo20EGyreUjwWtYz53sivIdasplAIAGCIrm
a+hdg/2tBSmL0I3JIEGpB4r7jAf8iWo2oazb7auAWj0R4IsPbz3lqolwhJYjgwtV
3KABZtawmfr8BPeHreuM8irvDBFhX8Q43ED/u1J91WM7eWseerVBJaEeO0uMO/sc
VfWC2SI5d1Sp4o7Zux0lAAk2rPa9JjsUlp0LC9feiUbAXqmrefcaqCGrVCFs2UAS
b7m5QDqkp78upzlLW1OP6jlirSHihaA4tdgQuLH6g3SLWEHjeX2mkXRDWW/EvKDQ
Oc6+yKRM6xxiNiOvMyt8jFSTyfLElS7M4xeC4fyU48QzbhAGRKKgroANvJlC5CMX
anRzDZ3sSFEl3dh/eLoZXks0R8a+0y5lMbkJY4IGeUD1DALKe1A8ZTjcZpT2LxWu
0FEFKeZZr6bLjLwK5pspE7e++GJ3d2LGHTdYktpHiAwlZRm402f/OYhbOlv2Dx78
K6GvVLi1gnHCkpf07SRvX3/37cScCUfVLJC3qnTda+cLUwRQZnrN8xcKsT4kb659
7fxBzIzsZsDESdDeBgJqOzDIkJ87BNxrkHsVTc1p5L72KAN0EXxK/AFDpQP6dgoK
M+ha7ernf6uc/VfPt4tboOrQZFAnunn5UT2KbpIzi1p0cEzSob14m+IEbwY8Susg
HB5eQGLDGJ6F57snYuoNQuN24LStfPDPnFdyTRirW143oiRDA91NcgHG+Y/zPe7H
aP0mDZ85pl73QMo3oAtIrmtcqN44LBnwjCoQ8BXPdUE66XWtRnWVcGRjZPwSxeMF
BuhBA0WFug0dS40HmSsAu69ABTpMezP0h4eq4oDzbeRR5JotymNWgbxLm6IxzdSI
BT4RHB1GCCNHP3z5dh+46vEhYRvpsEZdarLx9RGz/e8GaQI/nxzBx58jUVAQ4hti
5QkX+7vDpZ2C0dAfLSZe5b4dB913XaLiTVYByuVmYA9Y8YSxGVA5QzEhf4r87gfw
7mSSuWZkUXnYSDKqcvXRszV8SncDYQHFrE7OrRb8DjDaFqKktFy9dldkRWFDZ8OO
WlEDFZpcl73xOA/ivYsPTWoD+JdmKqXARWpvVJThBv5EKJWnjtu/dtdrZuCNcCVk
ehZ27Vscn4hcEQM4pfvdxJmxYN2QLl4BV2VMX7LxHDgsMSmzxbOVydIoY5KFthBD
/hswGzbneRG9xSVMFH4GMhgfkwQcZXONWMzx+NyKy8kDePDwu/Ii0ZCRGe71ZYMM
vO5GUhP0urZ1J/qwMJ5NPsU4yLCrFebEaxjn/4Y7ILpf6xgDm/Zd+QH483ClcKWs
LdSEgJqEq53Dy3poTB3imaPHTc34W4kimTNRStPsgKZ26Gl3Xx+ulH57/Y4o3RIv
r5pfjezKqSQ1Mo4AqKCCiqxbeEbpifi0PiHhX5rQLq57Xha/sGdjRQBFFP5rbZnn
x8g/heGKpFRKVPqMg1lMcgu8WDnmR8Vb02GPTdu/FfCixS/XNKKdyxHxWc0JTIBj
ZZoXuAXHqbzM/SnuhHFZxfUnIq4+Q6kZqQW3imWlWxCPw5Z6YETtzETHJ7q8wec0
5GFe1+BXZEgSJQsRcKoWVg9n3Qd2i2qJl/bblAocvdBO6na5W9yPYmyi4ok/17ZZ
wXUnvZjS+xJGRXOgSpZ0zvoNx9jWm97XiVNcx81fMzLvsflH88Z59CrbsO+vGFId
GOOwkOxpig1UrXbZFa48km38IAEmX3Q7MIIxFz6LwfMqLaIlGBQNNOWUU2TBVGtW
Nu1JlSpcNj3eiFqKDvIQj59TXys+R/tJ/v2UpMsFkCl/+1v+uQFHpRNJz59xmd7l
g07Ki57NPL3ZGEkaVdl7YhSUR4/Y1uZZ1nLy/J0S6Ois4C5Fzldkb1Gf5u2/K56n
SGyY4nYKTIATVC8/c7gHjOXhe4WBZGBTX9XAg9Dm34Mf4Uqa+eU7w2CvscRmmcH7
80WaRV0lMPOBBy/yL2dtWAYkAxB7/D+bIanV5exHlCFTIIsdK6xwTAtA1z3vmYa7
Ux1lcJ7hVrOcCSU2BmAh3kgIxbC3Z3lLoRC/PFPOC8hXCo903h1s+RCxyvGV+iUr
vyVgVpEPBbbOHAOYtxxd+K8ECM2OqIQXEwugC7Ex5CQeTjK2rpsEp1PI/qytLoNM
xHr2SLYTokg566JXkosq2UAHJeLIy+Mwoiy8Ve0dJ+UOfhxR5RsbT2nmeNjedO/U
UNHIgGgbIgyBwASK6v3aJsfpA+7XXtSP1xbNfcHR0fgZQH1S17ft5oIFdewW8lfZ
LXCsux6tkNkahxiLLV2jCZOYdpzCDct7xnZl5wXgEZD/Iw291uToU4AEbnWhW76H
dsEgRhI9BK//hdlcWWT+xFRwnq01s2ccpRRAQaSRT6q2XKFZho040gR95gNBLUHc
jjz5yDwLcLfTXyt3/mwKH2zXRb0aupq7oShe5WE+HJSuTZ7amdVuatntr0eRzfb9
S4MZgnMM1xogBVIBwl/4KxvLIcF3GKcjARdFzTPPORxJ5s+0OYbqDZ2nDZP7E5xS
w3/YBOoOMRrYum+qHHiK7010cq+fNV4Ha2z8+J60tNGRw6W+/x7JL3CuE+Nv5h79
lyWH47UwJAF/I7IRk2eP3XQ8QOh+BdTHA3sLHWvrNejxsq8dey9hWYFIOrJOalty
jL5eqtZwUK2n4HoB4oz+MwJ48/+WZlMkzV2rgbhEHZ0AQDBjsk/8iTLNCdgr3uXv
1UMddlTRvDQ1DSBi7SzAKpV7t2Sjt532IgD/OuQEx0bRD5RYDW9R0oDj1/CwmcM5
f+Ta1+5O2E0siFf0wHNvfxkxXqrXPlCRpC6YH2+d+qddtcfwb+XYrHav5PPqKTjk
mxmXUYsIi2XLARCG+rWcwoe4CxLR+qKWA5i64XU3/KoDgFT1nwv2ZEufeh7zCdUw
EL8JNBpxUwZ7EIM615kl2RhPYdSmFJSlWhcWvHaavp5TKjNRAH2zyOug3rDpUjJS
aRa/szfwfML2fqG2wy3485eGa0tvJm6Kbjpc44HvmDOrpupD2MTK18i8vioh73+Q
LcvzgUepHsttfCCZWJUdqJZb8wxwLOnA85JEDhkPXoJfAmzQsWn23/Rl6C1r8o6z
E8ecYmEPEoo3PNR7Sq7jG9aeDdFk+eVCVA9BNBSkkP1fWXNWnlD1J/S33rx8rQxj
Zo+GGuXWZPWKi6LfjUQqC5AuNyS2Arfn34/Hfi0KCTTupxUWQx0h67onVICGyA9H
IpSmhcTKtps4Mlez5828AYVDw5Pd6WXn3t02HXDTMnBfZ1TxUVG0jrA+L9KVLJi2
TLi6yflDxmGSAOqUhL5ClH8qeExRhJbp43gPjuTGyyNA1LUJoxrElYhyXZmyuz+Q
cUEdo5GCPp6yopVykHKCWP7QPWyINnpMYvQyvRiMiFHCbdcN3Rfb2XiQ+7jr05V2
Yot7mHkLY6ARmsPdVjx5bISSSJ6bgmtJRRw7kzNLcebqaJDqc2MV0gNPHtskn7gL
7UwVFeCJfkQIqT0vF+yvjrTHif8i7gKcCwRw7yT8kxYUVYbOM7MbNK/r3mNq5mvp
elDH960U3Zi/iNwiYC2AnPE2BQ6KExK+b17y9WYz9v6w6kzomaWDhn2Q53Cdjj3G
m5rhD5bEP/CBtBH4PWqku7wb0Jpc1jt6VT0tmSMUUlKqrPSvNaKmi3DZMiX3rjOe
H+U0MPLpw83ypEq12i5iI6YbGEsmSwgXiv8GKojYeShJQOkWBg/Zrw/j0/7Dquz0
v0sR/OozNdVKoc9XRCfiWOM4sNhNiAojtO6z1FhOtttIklKK4CoWwlNVfGVeSNuK
xT1QONfPDn6mpv+JnptLLtWduWQ/GDKU6pQykZBb/bmsGudlsf6uV3mXkV/1GJL4
63/thvjHFJWGYLTVrJuSFvGibEivt6Smql3KHlASLKYzFB6JaAAEKHf9u20vZUJb
sIsG8hPuzoSoeZD7/OngIvEnPI31tvZwQrHus92xpRJ38PFcBdKIHXRkLvhpG/YX
TY8EERI2ciQXR5TYm9tyxL/MccjTu486e0aSUAlphyQiczmyEFfNTt0xouIfxWns
1c1WXyI445xEKPThVf9CaMs//brxgNg28omGjK3kveIA7ozEsYLSqTeB3FM0y52q
VmvJoipnMixoI0QZIwHaCOkBPvh/x3hvC9QOdZjfhCKWBPZm3rkYZEUXfO4goUpa
6PdDoi30D/TxXOSr02TV7ZmH0Dg083TZ+qogz0SaTjRgDZMclEgfsyL4SQFN7pRZ
OqPyOpFfR9JrpsFf9jO2SFejpzzZTs23JPHUeJXhCkrXP3/V2P48H4UIvanru/xD
//hUaI8SG1O0izSJiM6/NkqjBihIkUWpcJZXRWyDap7Uq04CrRVTmfaR78x9mpYU
TAdvr31fFrvEmrlfE0AgJ5LZB66d2v+WZsGeO3an9yQQLcVzbRJ/OwNUF5eOIsUk
7U5BZB/5RxGMdKKZ4o58damsWQC/pJYzzD12mB1NV6MDR1SLvsxbjhyEjhQZULnV
UKBJwyAaJi6iNJxwTEyabRNCM+gg9dxDDKkLR80/V8jIHA2BF/pbBsitGpX9+geG
znnUhxnLBdEXHjTi2pP8biLllfBog/Yob2PTPKSHPeuA+4TDmv6bCd36Lyehfqmb
3SMPTGi6NbG3puv11xn1PBvGwTeS6KnYu0gkXmg1a2Y2ZQdCxR7soB1+LJhbiQV9
YlxGiC6houZSTg0KIrSkiciFELbXNaenR3YmoFMr2Ta+wo8iVqcPeNSOOIgpZcud
+tIYevbJT9nnozE7OkfHX40rL9B4Dz2Vuti1jjihWkIdvnbiDk7J41CzM5Nq68Cu
ksIO/8QsFr+g9vMxTS3Whb+QgHR960LUL2B02B3rdPcE4KHbikDQI4W6/SGIasbp
LgMeZUJS9a26BGuDceoqQz+prxNGBRPuMqhwQdG4EDy3JN9LCWaVMkUBUf1mREKB
CrUqSlGBgmAncygqS9BjHaKxpso3DzCRCCT30N0okRmYaoSRAFXK9+BxGdHVVf07
525zO98p+mNXVse8qzWDs8+UdkDPOu4Et074Qp4pGAKYJvoTUoB7ssFb5oCRitiT
d9XxjAKj1Bmc4+XSKLJ0f8o6Oyd6nsJ0X8+N9fONgAmvmF8u7OONnUAKz6FdrmX1
hh6kwF9elc8/HIireKCOEQnLwOf0I/Q6Ts4deFm+cGAb+ABSNmRLkWFMXyDeTtnh
60KLh85ReWbKqeqgImSLBPBkRgVOJGSPyickPjWHCyDoQm0t2xuPxobnpnwkLTkS
8DVLmkrDrDg1iD+JCsdKtE0WqXY/lywsjMIZ4l2OF5VSROzOGBuSo9JhmwBwNJu7
BuGLiSglsqviTT2IrUwmkredGowkheoF65yiD7YaT/8ZFmsXIV+411IvoWmJE3rd
r8bC931Gq78LDRv0kuFBKXON8MObNwwv7Xn1DlZrMcw6RLXwwsnrjegDEAcWr04J
81ISL6APrtMJanC7789m9pP7j8XVAyHlImi8HO5ES/mMezEyzTD/THJ+kj4AGbSm
qzan/nkSvzTYmmNtoSewnE4IJnq7wKvNeSPtSXRGfBOde6FA+X3KeDvkL8/pJgoH
fE0SgAj2khvVOlz6LudXMcK7mvwkb192IoiW8PzHyp5oZ2alWaHDS3YmzHKk3kkY
vOfoWR9kaD088ACc60ThMNlsTkQslQB6cAcQg3zmwZXFcHAb7E7z0k6Me2pd6WbE
XtioRK3fTvQNbPeyFgKALl6gcvOuE/zupRoBzkOLIzYTDJeCD0z6pnDOt4S48TEV
bMUWsM8T5SGxMrYv9rKPQIThQT1XZ7+FNuAYVNTWcBi8qR69EAxkfwAtsY0VI+2S
3nVYq9lHOkX3qZHTszyHMz3Ru7wtAs3ktJMYFur1Wi+JqLhzkxG1Jin0iFuNrn99
B6zunG3xGq5nMb/OqOlZNW/JCviWyPCrij+OGA4Z633UxOZodjKhqHGLOL/Yqlc6
Oa0gfoTPRY4wtTgNLItpXtiviDV5aO3vEzdd4QG12NMG0K5r0NIJCpJurMeSBsbi
qPeG664s8XCA6F9Wvk7YAI+icPWo+pnCLHLtKMM6/aKQX3ALEFpfWTkEBDjWgrUx
dLZDAp4H6+zI6wnStcWKdBBosua7Z8L42wuEKeukIZEsZthM2Cw166oFU/84APTN
J29zH1RTovO9tIUTcMwJ2xcvZWIU7d4sHML8Q3dIBD5k52/i0CjvdCj7pmADRQYN
w1L2nxSgApFeZAo8bZigiBEWxNnSKET4sBuJY4FJah1yBQeqUtm5yp07xKjzarSV
FXXmrzua2Kw1DC54/SgvuXpd037x09iGXIbsI8hE0buXic7J/rm7lMe0jXlhslAd
/DfBhItOM6XtdxVQbsbQpMwvtTeVKElWVFyf5VYB8/fW1cWwGFruZIWp1wTFwrF9
QV3vN2k1dB6FK6rUUcaKI7KrqZ6P6NtYdw2xBw32YSEUcvfHhrcL4MkIbVs4fGQ9
1SQVfKkqECxAHBUwZk8D/88qSdLC++8QQtUZM9GH3t8cqwE3OX+lDA6sOzU53ai3
eDDkDMBwAm11r9Od/6uR3EyJo4G4pihB5utyyMCvklqvlBuaBXexBvoCv8/KL1iV
Fe9ni/1dzH9Ka7Ya4g764OkWePwCntfA0H1XNOLD+Vxlsm5NZcFtey9eH/cSKsGM
el7yZ1f0Vj9+KEpM5dEhfQbNpgY6xs9cH7aGR/x3NeOtZ0pH7FXMWa/tHjjS1euT
4xWcTtdruzjp2wK0p5SeSxQduYV9/DuBaEP7pwQmvfapJjaj2Eyg1AwWulmNbwRA
N5aNOSraP9upZbfbuSsBHjxcdioNw3WZapQxt0FDZ4tXhCWYQ9FWZDOiZeU4GbfE
CNGxlLo58RQOBz2obbvkzTYDl6tB7eE6MPA2C8nTyVTusvzRDxcN+Gg7doVOKDOz
9nmHlOJPTrtR6GXkYDucK4R8Yl8t1eIBVu4xs7mxlIguyVDijJ1MP0krceTY/ktZ
zy4xUWrlktZ8PR7+EufgW+E5PjXWPo2J+9lC3GSL2kqg7ZGv5pygFdqmTY48FqiT
lRl4elyYfHwVCGt7wySTDjRUZwAozLiYb1NnamNCZijhsOM8lSzYs7uYlfFJScuZ
6mwJSi/RDRFpzhVxK1vmHxhiRjBd73NXD716teru9wSPMdPzNdzo9/1SjHaxFAaN
Evmc6EXh54dYQmyJO8vLJ4FNksteVoS/dTvIWjB0F6exYftFgxY+HsdH98M8hRcc
oMT4W1lirsYMO+sohVS34qp1t2JJao9oOBlq9xjkYWvuuqXcDjfNoPqM3NgQle9i
AKbCdtyaf/ACZSmUTDWFgxaDkBccOYTaes7Xr+XONkRRjvnQTeZjjIKqt3ulKs3F
+TxwnpNy9AQyHw1QmM07KiNc3FeDTq6rN00bMkGoQptUwx0AcWcmh44T3y0WsS9p
WrlwYNFTTJDaOKhcE8uuYOToponJg9SI8lEoT5VoXBjQzpgaAFQ+ZqNt/vgOzCS8
AiEikeE1MjP33s7YDbfFA7dvSV5kUsSt4oHdBhYKcpjA8fgqf13kdDrb46RRdteb
cV/MA6RMPpeHgZEY4hyI/yvgS79kG8s20xWjYGCe0VqhvYF/ffZbucqyAXPJOUkg
MXAS3NN/epsQGCkjK9TOVP3tcfw4ML72CMZ2iZvVyXyWRAubfHgsfijqz9ZbFsXL
ERpRXBbsw8+uQIFULDOihzAkWzURnanD2CL0ucKjZZ0GIkEGxNF0GDHrR8VJLsF8
n9iesxOKtd9IqFGigNLV+RnXToAGiWmU4iuC1XumU/qe6IkwrmPzVLgKue3sh7IY
8NZlcGSok7uiuwGWAFo3KYfcdxH7p/s6DMNFOOHO7rHDKisw+ZtA4khELWDAAlVE
85ay8R7zmJE66GHYiw1anQTt8v7VuBrqyi+eZnAKUNqfXnhizi+KVLfUsOZ6j9e0
82vQQ23+Hp21TQ5KioMBRaorcjPkbRjd5wmfckk7fS8jQ2YLZDT8Ob6ixvJpTlWe
qLoNrL6su1pXGQvq3QalOZj/LjVXl5btburF/vHLEr0zJgRE2HgVw7j/Df24DuHm
zbBWFJX7icFCSc/Uc86NjbvoxYq1xpeQyNhk09JM/3gh2e51PZpHHRUs5HNmbMzm
znDaYmQSghqSoapKKUjb+8gDxvH+6dGAKfveFLygkhLEy/1/iXFxJo+P6eL5kI/k
ELkQ4FkJHAbzNmj7UvKr8mtGYbDhbERvMOUznpMi5Y6YNNPBXly4KweiKNv4tVhP
3IyHdly74qLvooVnrgP3ka8ni2fOcpgZzE6LDUxY8J8b+XxBvSzdgURixZC9DSnL
AyjI0K5nPYfImM4vzodOM0KJY3t19mfPLtiN/WPhAxG4QuEZUef2pBpKTTT5JJf5
K5T6FMQGDoT89xIoECjZiU+MNbxU9cjtiZgtCq/PlU8th8BKRgcKV+CAR2n3gn4H
JXK7ir3WMSNziR7JL/u8fQG9WFyBrmePibOvjZ9i4V3MSE/LTLKiUAtT8DmFWVfX
hEawR3UCTup7n/3JjflQzPoOMT7ECyuAxZh+RgOQx+IP4RJfl9+NowXb8Uw93ljU
Fy4lDLhbbhag72G2yNnG0+gA6lFBsLdEpTkiJODyafT+Er3X3bdV/MKo8ex7kO9e
m2z0KCZo4AZNBn0FpUOHiDYbw6e3pQXHeGMUkK/UifLxd8ycnHwJ4XtY0pKKkKa3
sYtLX9z/+XYlDLEWcmZ9V9M8dblzx2UAUNOwmbLzq441D1K7OcFWDh0UrL1I793A
JFGPnO0oWZU+0DLM7dgEuRvPr7IUInK5IrV88LLht0wbUeoNb+xPX76BHmQs4jra
a2UEJNo++DFyzouujoKRblRVfxn48xuKsUuHw3JbS50pAzpwTPeQWJZCf0BX/1hN
b2qsy131IeuzF8qz6MsTdGzExurB9SYrtcSAY/QHzdCWCBUsrFG9rRM913j1so0R
k4OGDmY7njS4u9jMANIkTRADW5VCUX5Uq7NpKNmnMQC4u4+N91cTYO/1paQ8NnzA
OjHIMiQ9bWdHneNdaBH8ZrZXtol3+ZgfBcCRBJ7VA8p7jFLGjxmTN9KRQN9Y9MGL
7OkK5Zi4FN30DURRz/R4hKRpzrux9z8NlNgOIGuDC2AnnS2AfX4VwbcAv7LSnwb8
x7yWYuKTVo2H0NJMoIH5FJoGjTYvGRFKnsoCn7jpLJl/myvpthoj3l3xP5BpPFtL
RMd1YVsFzwPacCnBTsUQBlNKz6j1BGkoPR+FIwy0zTGmpTZ1/v7IELAKGC1xaYnC
+f5bs87jkHmb2OiUHyXHrejpQnYgDXZw5UAtB2u8RPL9ZI9+a6Ws7N8h3JRnLtrV
hKodVajxhgwQ9wZJLCGUgZPyRS6dgtInTWXfsF3ICOk/PLXw7CEMKSjWO+LXdnfU
VQ5/XS2Zh1zI7V0OrsjQW1gXoRC4mcmwFJ3EBTFRjd6hYW54b7h875xsOgT1Y+2Z
CsWEzTy2DC7bXSgITtfq2TO0GytMU0pUAyUT6000VQ1QaPWfjh9seN0PPhB7AKST
Uly2aVH99+TbcCI43KvQkGbp/e6aTMytg/gVerI5/9USHhw3ZZNXXRNNRvCHgdyC
1KGVhfww1tKRNLk50bMuALM0KikvECaCNoi+MfgGqh53evA8CH3uMmNukJZnm+sN
G01Iz52lSbgAMHKQ90xLWudVpuZvXW+gWr4erIfYmMRl3SNqvZ5HoRftob+UzG8d
WlzWmVMoxgkiobcDy59+zL/a4a7BBODOZbsoLzDwA6/qpTrTAIZcXAmhvThbCfXI
SsXFYcz4FSg4OdcqMetXIFLWmLRaOaQnc2DyQngc8tReQNgzb84dh7YW/yJbFFXZ
SbB4xyvYSjPbNowXiCSLhtnxRe+I1xS0egTsT2xOM2CIGNe5kCkSxhXjq77Gw4Fh
FaWH4I3YnXorCXOrzgnjqDaSSbKtAslqtLHuyx3UtjbUPqqTvG0jY3BCoja3ko8B
kEfY4hc6FZ03X/nzHso5q9CL+oLQ846ywh6tINOL5DKQ0JVXNdTTWscdYEyrPkj/
IaJVByfyPgcrBPdDwuKiureegYMpFVoD7X6g2rl3sC6wNUYfE+wCvKI+P6mmfA7m
JuZ+giNsZ9qx5wO69U6ey8Rge7XqNR2TxUWM4gXM81DM9xsR7JIxMjOTq0mNfzJI
INTaSaDkbrqIyknRuOMTDtbIgL3MpB3BRQDzuRPpkbqtrkQ5OX4G78PIC64Q0Dpf
f9dwg5msEgP7xFLBe2/Tm/i41foGIm0XffGUjg7WTgE2vV79TpZJbZsi+hq9Wcva
puHh5T6xCQgXJQBA2nYv2YLUv8FNDliiUkr2EHrRQ5op6NMkF67HVzHzixhtwNXg
2oK8NSF+1GkVPxgkTEfViH/9SAz8VEg1EWFm+Iun9PkxkQbF4YuEaO3clpj7G0x/
YXiIn9xjVor8YdFN5TuFqtqEiJdVwwVx6Bcju7Kx/yV6tZLs0eviNdhFvFAqVH4B
6YTGMdQPEm9IQbYtY0WxX4P7vzIwhfrLMEMHEO1AgBkg5t2hWkFUInIxLWGc329q
wzGQ/K9PGOUbAkphEVZfUeDmxlwlC8Rv5+42dmz5MGlDNtMEnnaW1Hjlpej4VNb5
rbValxN8B9h51oFn8E//IMiKtlWytihp3EAKrPu4fFtZPoBCLvA0CM/BxMSd5tdb
cC9U3OwNyjI6cSK6B07Nk3Wo4Kj3nPe7XwSJq7LAMlhZzuQMs84Vz2aNMKmursX5
EgbgsDCNWxBChA0gl2VbsHsPhoUl8w72ipspEsZf1YZWmN/gz2x1Gkjq3848jAdI
tvByaIKFZrIm0XiyvZOpWmZ2c5I8+T706aB6nx2V2W+yjA24EIk6/T4RZLfa4Deq
q6Z32wqui1I9SKUtn7Nu2UhuScs8eIK/ifp+eoG76Ie0gktMtNpNQXvE8BQlGlq9
ralJ7i5q/8qsqswDqzlgBJi9H8fmzmOmCdOG/Xx6TYLbmMItS49XvtymYdwqU9Nm
LWJTWD/2NdabFY/zWoZ8qyXhbPbuQS/60JeFFoKSDQ9vdzeFdJdMiNBVbsDoTLzM
z2wb3r9cE2fY41ujJnc1pMQo8Q5R05x68Ky596c0JjCHAdlTJa+b3z4IRUzTAUFv
n6E8D6GC1dOaprvX43wmMfxN6Ne5pusN9aQYSbDW189L4GiNSNw8Bunz58NEsb+9
dMf2HgW/Mibyflwgog5gU4qJJtceMMbumPctI47ZGxo2zfYZx2/28T2mRzK22M/g
mFGfVKUvAN39TYBiqK21wOaLqpV/BKAjQ+fp7ZEyKemZXNZhzDOVNzQI/7UfSfdV
8zSu9Vi7apl97FK8dKWm18muTaAj8pR5nCvfGXMO0xomko4ZS0DUkoobAEM3i95/
tKRXMjy/NpDVTgLUJlW62c9QPLbfOswVs71kQ1CUV3SvDKncotJ9Ga9v61UCisJI
wPyPyQENJMvTFyqBa/laoHHSRnkBzFcK7i4r+pFEAIqrr9vbqY55/Xao5jzoScqR
Kwv4HDalpWqeb0cVb//y4kHygI+p5jTki3UPIeUXP+WacCFddLvBStkL5a2yE9dm
5uqjjPHYQBtgRn3yqAH3bZN8tRep21lJJm2WpiUZUkbxFcIdqVQPkvFthLYERvxe
r9CABGfc9F16nLYFl2JYGQ0OwGei7fMdHfOSAb0M1U+ucayCO40wPMAhmuIBDX1u
XAgld/UHoS53obyLFx2nF6/IG+NgibcwzB8itJSQe+/I94gQIBAtQSozuaLeN+0I
SPPdKPCpTH+wzDaaaFgxORRm5Def3dNWskgjImrjuVuKiEpFm+DEZgYGU1vxhal9
4zpGfO1M5mN9NT5i9yGkBA7RhX7S13hooyRtUG9JHnvI2pWMUfB/8ZjqPDUdcM2/
Et/kobZ0NUYPPlBIBmWYrbP1dBJCykTRxAdFgUHF+R23NVWafHDKAN2Q4aZn0j+i
iETtduAf4HnQ0mCamsmEPCCtEpdop1mLp5ukHCyDoMQKQwSYV5d+EsYODkvKx6SI
FmTZo6Z48fBW70ekQI0nEppEhHz3FEw+mfbInN9jvsK28rfRt1pH5zB3zifMuhIH
LcDflWNH/LNuZivcB7cA3biKMw9TQqNzraOqnGX57aK5zTn/N4ydn4V6an9o0fZp
dPxSgYk00jbxE6gn4Cu8owGZyk8qLhJfi8cuhmH1qRljQ8YXcaQwLvGR+eUKAVPd
FIbx3Ty24pFIiptv35r6FYa5OxLr3dNR59TxZeiu3B8T3THuQacJunB8Rn9gKP5X
wc/QqJ/XPD/PzjDJK5QLmpr4o/ip36f8blEbZ0vBUJlhw3qhhMmIqUC1Obeo8Ql9
3/sv5l/1f0mJIr0/3dvvR4/xSvhRPhx3rvWdNdJNCCfoaVQrHmvLGcpWcUzJMhmW
hAXU2XtZXcPnRx16Hv6PdABSQ0COFpXIzm8s6+zg1cnJT3aogrHQI9w2P+yVmkPd
ooE2A+u6YOztGPrB3koQ/22sVgXLd5S+QvMykq7tqaCI5VC8qkKNSZt5Xz9bbG1V
HQZiUesqufcScDB2aIQ1UncxY9/h/ssdCpl7jp3aYikGYUtpldaoeX3S6Bx3iTXI
xcdnTew2Sqgbzez67AW9SMLkfOzEBGg8J5QRHMDTxLmy4mJSZSuwSwojrsKMN7rh
GYwn4ahO3/pzv/Q+HXQM/igVcoYDZ74BSlFy8PMJI/tLckZIVhul5MHMDgko5gEX
5kubh10r9cCv1/ixov4z6WJYoscUF3BOm8Ffv/2awMg3m6/oO/Q64pzk2a85P79O
potp2zbZn73SivQSiwH5StJOD7OfARrKto2OqY261/ydAQmp/pAxq0AjzYWkerEu
J7kbvoVcFRX8RO0apRyUL3cKPE8BZ0DahkxNTruwgDuEdVUNZ1PvmVtiyMzubI6j
L3mgZ7v9ovgLdgvp+wMg+IM0U3/g+MOw7XmMAlMt2JA8mgvVAkbv70BXphHzaJ0/
6mk/Iy+5v0XlDek9mtHNfBK4ejgv38Ihzbuehzo4mZhvpPwSEFsXk9o4unWyfTaA
g4eTJMSFr3m6Mm39MJ+oI61t6qjc0ccQeJwhwIa1WVxZm0anU466TahQ1jbS3+Qx
+kB3Fhj2KoMWWDCWIvo0S2u+PBtdkrPLTjffBSv8/ce6nR1bSXVI5QIWnpeJUtei
iEjUk42o8fXfQ6YQmi78/KMB7SmhXYY4QAIrH4VkVvEjMJT95HQG3bo6eVkzC+1k
P3e4sbxuaFLtH/BVcS86ykgIBCdFOmJTfxpIx+0kFIZfPl72np/XJWceCRM/My7K
oPwA4ABTfSPlJ4PfgKI2XFl8bf2+yf8AjN5dkI9cAXuSuvGrlPdrmgFrk5tvBzm9
da0wYZh0sOGzwsmOU3MqkungymM4Nbix5xuVLSVBZE4zuDCfHjnhq2HCy9W9qgi4
Zbs4uHvMhjZTBkghsBBafR9ZoosV09oL14uMeA1bMIrFKZFmK7WWQA1u2LOzRQWR
cvMzLUvfpootu32DbhbeQt8UBgm4/8ObuCCj+yR0siawxlPh0+hVBjlJu11HhRBa
IPPQMLuuRusqSXe3Dy9/NQ4/3jfidbjnkea9u76Pjm3O857sp0HjSQ4urqtFXiOp
IxH1WOlKaQwF6yiewi4jAUCSqn6aJ/0XbBXeVhfLzrqOvA8Biy/5yPir+nq9eWSq
NkTkLKpwoTWRmLDKv3JzIVA/d0P7DWiV3bCKqPaxCCUhW2MPnCfZKnieaYEpXpqc
+Tw/2/P2vhip1AxOxTIWWLMEHthsyX/uFj/6YdI2ZeVKiq7R5JXcSvlxYo/wMikG
DTqBhOb5tjJun5RedLtRe0UugVRJ+LpyNIY+6Y4xeqjXRVlRlmcgNZj5NUb3CSxp
pO133HkZs8oICh3XZwStCMm6C6gdResfVtDy1SMSwBgrQfhhnc9Jl3CiQScRBIep
dgDaUsKd9V6C+DKIAS2TnyUn7GASAJTmjr6CiGw05RJ3ScfZxa6vpDa/16e7uZw3
PY+DKi8mTCmVZDO2/N4IMj50dgSfgxAfGr+i+KHVRDuBP8eLilTvI2BGu3WZDnAP
1D6AFPcmJOIYTVmL2CRcmaZxcvvPBe5AurQNb3otPELXiDH4W5EWFurofglVcY3w
EYeLIkq3d82sOztsoxw5LgmpU5N3hDU5lk3Pm7XQBnM1Qi/12s0NX11fMEb+4dDX
gcS/fzuh1ldKhmBu6K1HhaA5BjWhAtTdBMs1b57qCMP4s+exEu3LnoLO/L+9xigA
jjVZgpimsqbaZXqgWjhfHFrecB7oJmwyGTEWtENDnjoAOesCrZaaiUkpQAwKz62q
FXwqeYYMgzuIZNeSuP2VeZYc5s8i9XJrhK2RbN7HMDeQP31fbr7Z9gCjsOOWXdvR
JY6mAAmPW0G6tiVU6428W6Xc9wr20vmDJCguJGARJrYYEZ8OT5GySkmdSpowaoPV
ZvHQf0tTrmSafQEJ3o4zNOaKly0KGES5kA0MYHgAg7/J8jTMJvUz/uzYuWfT40BR
T6aytlOyZsTQD3lR6iP4XNp6+vztj+7XjZflJeWORou92jjADB87EW8OciwM+1K7
xlnDOZqLvxpdITMc8vZTgUhjVqidlXLaUmMr1GySLEil/bmAUh2hvtDCJo6DoleP
3IlRDDvCxXT+pfNcPzduyH9brxKBP0J/16UcIxktCc2pirhgv6qOhoCW7YKiHyad
DxvnupU6BfBFhceDQOysydsEoZ+FHArqDdakoaG6DMZ+wtvAgrTeCbzCULthCX/l
PVlULTB+CAdi+Igpe9Uex1TgDV6t9Hky4CKheKw11kXGp0wyoleLMguqKVU3Yjoc
g6LD5BUuMPIsNjwHrTpALoZVvxcxwwcWJKBC5LptVwb4NPqRfB73Wr8YQdtxJiR1
YH3ds/TLpbgV1JLSiq/GuzzfN3o04oYCs8cD45clMpLPiYRvz8sEB6Ri9EAQ4Xgm
124K28owXCOOacj+kFg6AbKnEUG54PKNq4HWiBdtdQD69S/+wkaG0dYOvBl1qTzq
7oEvLDE6jymS0ZxdtZmNX6PU3O1WzXB4ayY0kRuTJtHKH2S20DyUi3SfWnrImrax
SSPfCq8F39GujMswZAa7/cSKn1EpA+n2Vj5pYpQNlVgMyUrnzyu8697LxkYZyVvV
ZQyZql2mLtIQ7pRhjagPPSKqT+/cbtHIeTpxyAi/HIX2MHZKjJxWn0B44VX+wRxW
nvTCxjJsZCQYdlxx/5tz4NevRiRmB4zQ4+wN+55MXOQW24eDgz9MMx4vseSrMToa
OfoAqDxOV/j0KmghCKmuWjo7b+07uqCKF4vovDMGz8az3y1bVWqII6ZfHYWz8gNu
6iUJiwda498KD3b7enYAvTC2dp1xEftoor8TP74jEHF6izu8UDutHsQ9RM243K82
p/IysSU2zWt0q23HoZkGlQvaloxWILrNqrKQCsaNE3n5SnvmmxLLpeXJ/15tvjzp
sMrdwKP7ljOyoyeYbBkvMHaufQS4XUc2T3rSZ/L5IxlZSN6zjQXzpzCI++BeRJgS
DDByFQD2on/ht8vK69SiIDaPLJ0O85h67dM2KABQoXP6PpfWe+jexuLs/ZPC11UX
1gPR/xr4FBf5O+comTysV7NOHqPAR0VdiohNYxzdHe+eHmuwrMlp7hb3ecirdXOQ
y3Twam4rotqX7Zy3OZsJBZWOXn3be7vekCKKEtnrPS1g5OYr+TB1zqq+L0Eo4hO7
bOKSgNLnKwR+Qj0IPDEL+iGzvnEh/sUKvBqliEJjiWKNlR8mRI+4ttHoj3k3uF51
h8RpeXvuEykA9AkQ5i26RZUhCHpG9a5e962+Ym378zI6C1HjQovDwTKB+4VnWLXN
5Ih5nlGq0Biwf3RHUN4ecPEO6OU4hQfX0msrtUz+4lIY1iTFkRtp/IQ42dSD8uzM
HjLchsIGPYbQwx04CEcE95gxjFRzYAIIRqmen8oHi0DNLFeMfuCnj32APuYMZEl3
2ZE8jJz0oCxlEDFihgmxLStMg2+8EGYBGj6AG3rL0GHQ4BPYkskIdnvNNuccj6BZ
ag5uHWUQYANO2xxJQBs8h88xQwovZq0t17zoZukK8d6cOgkV9KHYpGbTdOzZe6fJ
Xpni/n4Pji1SdTGbDX5AD8AaYtbY6fe7uYNg4tCzTwZL36gwGt5ehUVyfcrPHVWE
dSAK0PD52AWDcO+EbF6CO2x9Nv1ML6YKW6dBhRQRsH6pFhJmQHI+2qw9Mc5sXsso
gxitFmenopzBe9lTJG/4h7vT0OeQPH1ymDsGhNppL3yY2hZLpUYJbyvhheIIyzuX
zIGSK7088evxaOTZ/8fi6Pbv8YlhjDJFDAKxtu8w7RiuWSKejbUk0WNulemyvoZR
4JTVIJI2tkAB7d2PkZfysZ70aQZakQU1/EXYFVm04nPrv4ajn5uebl5Z8styJn6t
WYxJ2F/u+tWasQay2yd0ypEHzP2dhK+Qa/kgcXQPfKz9+lLkg8lSYj/tEnwbJc8Z
3SUHyDJ8osDORV7GLXF1aTSIeZljnzi7OMomEne+xDq7PGJWKh69whXUn4xf2OWT
ee58AGpmINGftaiVajCXKees1dZWh1f5lY1y5g0ZTOROYIl6AXrC1p1bsn5H7iot
mukwfskdc3EHHJSAw7KjssobxKkje9pErTjGf1vAdr6X9HQ2JdR13jwoFQNIqIaT
dG17tN9bS6kXKxN9Tv1sEoTMc3mMSSYBvQPykeRA6vgx6eXu+gppSA5I7eEDVGKX
knGiin2N5uFtMXYrKR3atNCJHx+m2aJX2x52zudgVczkOhtzhshjCs7r8x3T32KT
2bLDvrjjsKndHZIQPJ1f9AvG0cLyapo7Z6eKVqNzqMzgjbulzVIpamvantgEE+Mt
X7mnrxbx51CbC7KeekWyeJFC+LqCtXMLj/G7jZQuhjJhyHF7ai6LxUmnsOXVsQnK
rD1OeYJOOrU7l0KEwmTdtrdbjuWwa0VLI1IcASwPfu17Nba9A062vAtlasTOkaWa
BXgbphMKydytNswIB2vy9x7R4ziXaUi+79RqQ91ktpRYxlgOb+09PwhbB4VYjAyc
/h2yyHkg1ke2t8SbZK/PcuNC3DMYF4a+ZvksWXvFV+9u4u6JZrHZGe2oWrxqxzWk
MdFoDW3gIxbTAZxYxUAUBZ2dYV21y2JnG1pEKco3YGIb24BPWvzMTHd6LZ2ArGhi
tJRVh0jHTtWbyrJtomNFGDz9TpOcPiSkysfcipwWawcUnqy3OY7RYTctMpcwVxgb
6St6VpfqFbJU+Osb6doHu6JENZMi/EAtFcwCAu4lVPopl9TiGkFiAVgBhuUlxVm0
2k6YUPWxlRrpa0OItYl0mxK+roofb1LnOUYku0sBa1joFRYeoE3tlgDx1Gk5RntT
GC8qpKv2ZD77kIspowX51tvFQn+HLeloxhtKZaDsTVuAayNreLgCkIjvLNzViQYW
JOCPQZXTS15uRpsVy1u7dH8kDu3Ypb5EAhm5jvMw2JuTVvcrCULUu5Hgf3t8Y1Im
oEmCv/ewaUE9OVzCpprSuokWgcEI3IADqo31+4NfgYrSyJeHI7zCuVb9w3Hh7L3v
8PJ8w/+NlcSMUfaUBeEOkVcZHJt4rVdM7FJ6TpddJytFCI280pqtOYmIAMccpVLY
4nlBHKKbCFxayOOYIDSLvbpsoCQDgrE2IZSR9yypYSGC8afHqTuk7DA0VMQnjDi0
B5C+tpriN164cpePd6Ta03GS3JEN1XbMiilaGeQPqfnKFJ2Khp0HgPzb6aOl8gCw
OeC9FKxTQxVvpEAGKgXEQMWijhN5tFzUVu5AhnOFno0KRQ/dhIZN/25/auh5+8YX
zja7SKyBrPpPBnx4dpifz9TvOfnDo/CXKYBKO/Mybe8Lz5LxgXOI0GD3J2xMcuD7
ZxZ1svPuVpP5emFPFTWLlOlVyBAaDnxhhfLw8U48gh0dIlRIZjfJ3mXlFZDV18It
YNWuwTP0FGxAgEpQ41G99DWddgj3dvezhAuW/qtwKIz3aGasYhvqd95A1lFC8a0K
hSo3W7nXaAxZSlCIcEnNW8gTeKOAvgN7/x5KY/IWRpCgjEaYo5lR9cfKYhvsU02t
0+Gj1ML1Ho7UtQlid0udXa2eKy2GjS5wbSXPxMhbliLzLmvMhxR6uWsBp7vaeQrK
GiZYaDYb/SYZb2l718wlv5KqJwON2r/2RdYnV/pEfDpDenRNuzhrn2TdGZrSaxBc
Ol75T6C5jaA6m9ervSXK50Cbfq+L1MSLlsQ+kCCyxQ0/l6vZx6zx04GAJHaNQQBM
0DhXSSj3vRfyTWKFwmvzALKNH2te7uBqXTw4MzbEfsnANa8xllkTKgiyMJsMq3Nk
m+FTjEqbj0qOrD/mUfnrqHIMMlwcUNhNCtF8Ij1Q9jcw2PUuHGK5ZQ/gR7tuXDzI
+4x6X/eNmqlBmKWhi8yeJL5VgzXWOyV8ax7oxn28+gbsK7QZBbJqUTX5Ovz7Milb
5ivRCgiz4OKoL7yNbm/QPWKO/iE8/GBMwBqeI4fzvBzKImEPL5qih1u/sc22kTe7
aB6TQSOd3cJ03uSABNe4TwER7mbPkpH7OqeKEaOZZixw92sucBU5JFyyI3N54Iy3
79P8tpu0qdfSeC2wE9Ouswt+r/x2VOAaztrEnFfx5ngYQo7Tab76GkF2Mhm4oKu+
mSGp+UCuTqiv6Ehs+krQEIJY3HunzL3Xa0YH+3vXj8EPTyopRESkCttUqPl/sL7Y
CJUYTpOIOyJKDAlfBt0EljSanElt9E6A2v0Vr0TJ7UiI6b6JhCld69I8bPcYeJVa
D9ZKkun0soYg1FKvfx4LMrI6hSRJDlmpEX6Gt6bwpz+MrlQnSRBCTXvdo2LShbnT
HHTUQsREURuatQHLSk80KW+4wQhiHe2ORThse2F+wtk3n01As9kdEB/hriFFAk8j
4nC2RW/SMAAGXLm08TgrjGPq3GeDEAfECoS0aCuVzz7VBzHU10DIa2EQ4RTKlCOg
bWRD7LGNLAxn8FRsdBvDcC6Z+ThMFlCfsbx+tsReK7B4ZI9a/uW5NBfFUkWrnj3l
PeabLjqi/rndCFsD5jSy/yNzdgSp8c9CELVY6N8sR9UFXaTvkPBfsgeWKsXtVCAK
ecMI9JP3BekB6larTUBN2HlDX2j5VzepSahbgrlRE0ZwuKSR1Vs83LNET4/My1WL
TcNiiyN7vgEW0gLyT9Dyx/HOFvgLR/lPJiNIELaGMmUKT6rrgscTIPu46/yLpJiG
k+TshPNG5Iyqznsr3rfjk8WkZ5Uy2VR+49DE6p1kY7fOdSud8V6GDKrixR0IwPBZ
r6qoMbU2bg50Zoma2EiEPQgyVvzbPK1Um7bZHhtLeWZEA4cGnhJ1oxhn8Gjckg4c
l1y+Cq3ysEWD6NmO/aQaxVzWkXMjqNL1LNKrVgGadVy1uZ5/bVZOsRJwXkdcXv34
LNKNYOk55AeNMVsfeJ23ePLC+MbUHZx/8vN4kvFvx3lfbcvjkj5am0SISRrcnTJE
esjm26TjncH3OXzpZrTCy1rXWrJkWVRxlKi/TU4qtBUpEt16/UP5gfpM8qx0PPjt
2YLgZ0nQVgBtlH2LaejSd+OKPFXVahL/5u3s2nU8mYjZQ5kAv8SicgF0yDas2Mc4
44CgsHL+WqZBFgte0VMbA38G+Ltq8X8d5NWB8areeojTqx4P/rZmqCKMbcrQ+2bW
fdLjI9iJIEQePBpTr9OPMyT/gPIntbQ8EMoQjqj2jPtcvpV7cKPJvnm1uTZj1wpd
kUdVYiry/MGwUXS1DeTd+3f8Y9+gcebi3MTVKC/0mbloknmkhFJZSqSuzYirggNC
6kayx4Udr2m+J37PRElC415bjiuRRlkuN0k8YXbAx9VV7wWv0dB9NYE1wM/RlPlt
vy8z7kE40QA7pQA+QfBuswjJuyHbvRmNlSj0Xnlh1r3JfPA1q/TZK/MiiICUjK8S
wECmcxZdv0pBS37mvB3Q4uHUnlQ3HpK1gknuShGC1aGny9UdZkmZCg8F6Nl091Fe
DQjPa+EWrG1H5U6QcGUwUUhCSbwkSm3L0aCurSFvWdAWvEbQcqPlrotPQWavORpm
JFLFk5ftMkii4vb8rqdw+nZPF+iWKwuUy7XIp1pnE+iX7ZtBaIqJ3IV/uowdzjGL
7rRafo8Oz0zZKjsBuJ3viV3THXtFeRkqHjzxCDxjAXvL6KgGFliIh8wQvt2QwT2C
yseS2iL9ytOemGQRq/6JPh8p+AWS9cN3i7eFViq3HP0/iRJlFxtB+f/X60jyR5NT
SVmrmH4Dv06Zhx/733dsye4HHoK3Xh9off7ZDi6L1j5QRpE1xI9M8fn8BrfqeLn7
aGN9nXiBhyjNXK0NKbXE7L6FVDGykcwjULFSTTioBo+OM/S2pcyTo8gvyJsFeALL
4xrkDi4fCPjULjOL3/6TLGzegpWBxBneCYQdEN38rUsLxsIQ4oi53AGQ/kBRrCUb
6v6m6Q51VTEpbGbm3mwouLNhA19LOOshb6el0ml5TSbxQSlQspjHU3zi1i6gyfa3
n8r4f90taulg/I3Qt9YMj/2JLWXt+DS8Lv/EAk+Nc626CuCzOZpH7QxaRzXOrb92
ixUTVTAUmpFv9CVWUlX86tWxNfBF7PjUyUPu2a612VIlzpt/OZinETpfQLtGcoNW
1xRsDCN1mXXeqOs9TRqYo2fVhC4dIXpUmgk3M4w74dj7OfiqOTuO4hgJg6mwVNgg
qJhovJRGQn8PDCiXkGW24R+pdM4jRCkPZd4yed0EhUwf7w3ziCp03DdWvqhqfrCr
gkPTDNpkYV/vU4TWsz2DLAcNxPbYj+IcE/IQq9m0bLQscdh6oXyEp3LITkRf5SbS
eJYg1zR7297DXm09JmNwtv/NCY1QlAyKWgE6zGLiUetT+Kyz8ut2ylUtg0JQmsaF
IzT64DU3fQXlkEtPf3Zp/1q024FrhrxnWw21JYFa0wZ0jXrMaJyvTn2Yhgju1r0e
dNJmoP3+bnbiegplt7PbVSjUHHscQyBjx7i5xQtlv6Sz6kpzO1vCYYKWddzskNsw
7ftcs+/jJZNFT9rnNvqBP5vkUzsXhR1WfcHAo9GMtJoFzc3FsLIthsu506Ub7HGr
MUN+wNYYQh5CMax+IQzo8LocTN/y1ZUuj67iN8LQS6DBU/GwUEb7fzWRIQD8T1JN
r9RYt+rK4aqvA8TAHqvqy2KyHpTBCvUhMAebAPXBLmxG8WH9Q6WJN6tLO9YyCeTk
icK3TfnRupzxQFwQ/8J7kr6vAgXFk9+WAvIyvr/5qcKEJClcJ26y2zaxQNvI71Eu
idU/IdSmMaAM85WoIjWDehf0gctwm4UbteChpR7yA/n7liPSFk9IWF+X2SSVzWX5
1rAkNSlY0ftO/4nSaWCgxzXVP0zIHzzJVKIZ3ez9bKu4ISQh6du1cXiUsRJoHHg/
9+cRyDyeCjTq4Uddw79BTfF1JokzSoVWW94daaYvZvKNvFH9vzxsCV+uTF1n139F
teU/tvYVqNK2lKdMbqfR7Cn6klk2bu6mJ/nIFD5LWwU=
`protect END_PROTECTED
