`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Brkc2vnCvSCSkp4CY2ewETteTUD2+xu7B6HTJx6XhhOPBlr16Bno2CmpUe6FMM6v
8IGpiuqZKHY5jAF6KR2ifmOCpTkvlZSFB6u2dG2DgcD93u7bwwBAL/zGbP+WXBXP
KYqCulLFH86kTq9Hh636XjmnByLC8HV7YFMuMq9lrC08cE6GyN9b0Afflv+iRd6s
SS/zTU95HF7ThQkkFGpWacvmyxXFRv/WIgO7zgHauQ88s40SA0KqaDPlQCgI04y3
Wm50cbGNIBdOTVNcvfX2670TaCgCvpbzxLZSdtHUaM8ribHB5/X8t8mTHskwmlaO
O01TKLFybQZjHYqhGoR9MvSpZOJeBSLHel1uHmSS4Dsm1D61zIG+XEVxxq4m2Nxy
ZXTyvakBgOmOCKo8n81Cnn6F3dpb8Sb4Uf8QeFGZcLHZbLVHi3R73WWY42Pu6hO1
EymuvD6kVpRA4n4C1dFOJ9jf0cZ0uMSiIIdYxla97WnfozczI3QesY9nPBwMXrC/
OFgCP3PnpCJEZpWGyIb6wfdh6tZS1V0cUL+TclM+EPV7Dwkc0OgPIgnW1mvdGibe
pU2n/ZtTYQRzysrZBjPdJ8FlBMTuy88/IQkmBERZ6mQNc4HCZ791mrcEJdU3B2R5
Nqyv2FewOyl5YiO46q8yQqdMxFaBm15XJzHC+pyMcASbXItDWqygykQlpQFlzmzW
oY7YmQYpZEDI8W1r+po+HsSQu30reFJzX1ahrLOnggMkC4HZus8NDw9G3eN8qutk
JvD4uJul9GjYyvPtRi3Vr32vT/D+LHAWjMX5dwwPshyA22aTR5aHh8LAQSBH/ulF
HAFuA+HM7gce0ouMJCmBtcoro9ODeVbUlv0GjAzD20jJzrI5e5JE8pe5+L5e4O6h
S7KG1bDkzClNfQyMWZ9o8WUE8MDWgrvb8bR7vFjYESK1X4YtInlpE/6ImjZlPtiD
B9ZqdZ3ZZiJp7Q2dQGQcGaW2jCv0ggr4WO1KMnv5QSSnEP6QwdYQXTo8w0K4npra
/AYXi6U6u9fQpwAKm4oAU8Psvf+qwrTs4vWWpnRNB5pF4kc0qGCBdJ59e/WMx+H2
vNDYwg/RXfU+4QN2CfoffNwSI+nACLSNeV39HIMwbvGmgbq0MeKkoJHlAV0zDPvc
nVAYqg/hzCKsDOAs1Jw3YBr+lGDcY9QkpgfXuQNFFdW8j2pqNUDls7sbqnQqIgdg
l0o3WB03ER5CI32glgflS5MuT204eB4oc+hw5Xx9MGgQwgZiiZVAAHS+kPudCOuj
x8ybHO4bkdoloPqalQtJEYr5GDSzND2T8Xx2UYnZU4jyHTLoVuG1Psz1qbxNNQbe
`protect END_PROTECTED
