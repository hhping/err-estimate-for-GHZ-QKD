`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YAYgugyd78EhwHEbdt4+Aqb76hz03po/Fa6MHN6sFAlgZpWHss6LM22z54ydJEUj
7nCxKR9PUVj+ABA/pszw+XN5IJSn2U1YbK7bQgJlkr//3CzKoKzY9lEU3EG9+7b4
kmmtytP/+Drnj7GyBvkQvf72dmAQkq6NCWMlPHgBv6TAAUcrNsX2NMmct4yHky8Q
P0X82C7rVl6cHk+yej74LHAZ6itpJ0+U14pwGws5S9yZytXsXweTzO3Bojxg/PtY
GMyN6p5Ok8ySZmyFhKTeMAI4jevZVhlVV7zVdoJp9zVwUUulAsnz0zWngE/tm8wI
Q3MCaT9VOen9shbsxOfqkMeGFE6SE6osRSe/8N9NmoUHXV4RxW885EXpkHkC0SGo
v3+1cTb//zHdoMwHiljiY6Utg7FEFUGg1XGITebFWYjgUWqD5dLpc29zDqfx/Mza
k4cq1Xr44TF+mrc0zlrYwqkutKuMN5vNrHINdOWbIeSBcpPqiuCRQ6sGsq+4PViX
QKCEJxYVWc9OXzsx2inEMXODOJDUXoyzjZy+g42jeoFCZhWY362dKzEOlA3Doy/c
35qk4KiSuvENJX89+I7T7/MIfipI+bmyFhgo7WeuZDsTb92q2bqk3jvXhN3Z5tpp
2Cj3D4DRahtUU9hoa1v/uWxCMTac/lO43erllz2bxbAy0iZ3Dg6SDUTrk+ytdhLg
CisRh0D1yOOaFq1rEA5dNcSvGRPRFOy81eeA8HaR74j/v1MRMg6pfQNtlyio6QL7
Xm6CDXg5/uLR1eVqdsrNfPtaGKeTO6MNaDexK09PS48T1KI+/2uiMgsbQ21AdItN
`protect END_PROTECTED
