`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jK2TlFtyWVUKVX4ZzBPSpwR8GnyOAn+K5u4QUXWfTzL4dm0AGMSp11XZIt96l1iw
QIR/uNNRC4THQF/Q1ZISFvK2R5RR+3uSZdYbISJDvwxtsbEycMgIDYa4A8hxjINW
CdNrEZOgdPui6OfHhhUvwBdJwJc0lzTS/ImNy5ybo/g0ce+q6+HLclaZTPL8hAry
Kq2zo6nH+CBGDnyTwzPot/+Nu8tBrovKw/zfdrMn3/vS9lz95FdmiKuklvkwZd/h
2WRBJtPRgT6anfj3MvFVtS8m9c4TBqGGuo6vYLRfDLKoJvo0qvYolcXtIyr8Eu04
lrvssyXjKxH9wsldmowfdMGBTbR9w2YWjMhnCszu+Uu2zGiI/y+rZSox3EcsKrrQ
MHwOocrzYMf+eqVDxAjeDpddrl4BVHbyeVvE8BR2n6EYR+9tcULvFUwN1616PfoE
bQpvnI2JJSUa4Hari+8YikvRbDRtbzbFRVG93zzrzSfknMS3Ud4NsnSz4tAZb3rz
8Gk2DO3rxpMoDiaWXNg6lOrfyY/lfSEswfrjYfjpyFmKAse4xec1BctxhIZ5i6Pn
9fgau1cfhAfAyP03uPZxzGjtCM67Kq+jgT4V0BOU+wZVyNJc3UkjRJbDevp08CEb
1oxwWgDj35uGdGbqrmw0CQ==
`protect END_PROTECTED
