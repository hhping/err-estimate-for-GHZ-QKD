`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrJ1SpKY9IgqWBcuTEBI98ZolhhaCs4WhDc9PIbn1w9OPicSfS0gCBDbFAnOg9eE
N0NsptipuUoYIEcHvfaKAMENR+d28EiCeyOvFR70VkxGjJFMCO7fEMkUWifssu30
liRNEkt3FAikjboTRl0zQGZdv3RgnY+XIhJ1BuIzujW9B17cISuI0GIW2lT49Cwj
x88XnIgU7m32J7JoA31J9n8KSUG5M5irLUdyBO6xj4+n7rZ/GSeqkIW6oeXXk2oD
PvuuaOBNwXgO02uYcIFaSrsIMO2X9/QBuYfkB1T0tT+3AjMGopHZznJHxvdZbPE/
VWw/FYoOvCAZ+eidvH/R576JrsYLWhWj16Sy4MLJJC2xElaoI6TPne5fBYg/kfbr
eljptc+f9V2sjJA2LK8duo6Bf/VlNghJqH8lX+hJZ06FRVLEqqklxtiwiLOdAWs5
RQqZnE/VbITfWPNRqFlmrw==
`protect END_PROTECTED
