`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZVcr8/nfAcuIKUGBRd7l4JQjhE63pvF6zrV7xQFrE2Z7UN9e4TU+iMZWDeLlUMj
0uOqp1JEOfvmMtquYjUwYygZ1ogKEqLb/OSy4ZFBXovJMlfdZT8ZSw+5x75mxLep
DOOvj3C6Sc9NQgUHt4nluva/97jKmNTsrvAcxMi0uHl4hvLneMeFjNEfn/RjYwDU
FgQ+1T60OrU6obzIDL8F4pmpAhmDsrdv3TqRn4a6kbuuGzWjlN3+Nk24bT8TVhNq
lG2YN1jdyjr3EfrL0zKSMVCZrwSEVSb/vq1oAc+dMDPZXsVryl6Qb2bS7pDTw7XK
+/wy0LE+CWokHNFjuX4LrKsXtw/bsKL8sUUz+DqoM9x2aeqGvf0TddzmRg6XGck+
YsFeFn0dzHzQJQR+qTWOfF6lfvz71mHLuFSOvGMIZPwOstEv0hUisC2yAivFPoiA
bvwW3Qbp5N/XxA8SkcDeAD1iTnh/c4NEawjkIaKZIFV4Lo2IQ+AhA77R8cXG5EQu
045SxqdoLhUj5rSqBF/jzO8goljQl4sZmTixgUhbLx+HpBTNwJPuMO5nfybEXe00
MxG4uiFG3iYB57SwFtVUwM7yRF2+0qjx+HgeXkafbBWkXcDGQSM7FWyy+QHwGsSe
8BVjjR/3/34LeaLI/5bYRu01sTjE3sxJIdgRuLSsZEw=
`protect END_PROTECTED
