`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PvJlKpzXLgcQbDzAPsKgVpf1uSUNcUEYHfJ8yw6bsByHT70ufHe/0I3UYR6NL6zF
g4NygevTLiyLBewQX91lKI96KEsoaEJP4g3AtS96vFwsJFkU/yCvNagvHxhR3TgD
9rOY4Q/qrbhqoldwy4qTHabNLCLZZcJycJrKZH4TtqSeL9dE11LBMLB2+9daqPPZ
Qh//Y6UDSqhj9u4oi6qKA16NGXgi88FrmQDCltuSUJL6ZPW338DNGOchBWrZI8DP
brtBgKb7C/ZNZCXubyUzbXR1S2r98uwP+1Pru31IEatSlbO9qSzh7LySz2wK7u/d
RZztigoODaSUTkvUR6OyadxPvtKIVGsk+Z9UaO2SJN3jYz5x+BFpK2F91aoiSiSo
Ddf94D6XzfzARqw2Chn+pfndmM/VI3pCyXUR9uwIhBncnusTZUITDyymgn7X2RA2
odTYAYn6JbeDtKljgQ/Y2rmupC+KXGb6NLwG4Jq/XX6lCjxHelQp3ysGBy+TywQJ
Y//2kx0Niad4Fs/NBH3kt8TdAXXcJ1V9dJTPQLa2vE3O+NbNsrl3g9sPRjX93Feh
gc9HJ35SB6DVG6nuzkeEmtWJHWzoaTjw42+UMAiaVZFRYIN352TZyNu+cpdmAH5L
kMqhTn2i5Qjzs7x6inFU6N2iTlur2n4bqBjwvwJDzSFyoVZCiaGq7ME5iGw7DOEW
DZp8zcGQKgqk5InO58a8B0LMWZHqEyjDfjt6DSAInggymEyObgBgQcSrvN6YwS6N
hEh+0PqMby1/foWs+mvzS3GF9Ca5dBhY1tFmKg1RcR7gZ5BbyJ2S1MNlzBnLf5wg
dWBhgYAIJKGdbKNr74pdngd7+3SAdx4am+NvoaN1kaxGi8U5EHZgBFzvDTJUNZTS
wcPvm4Y5GiAbkaacN+/6zv3gjqHyGvUCd0f/Lmp8ZZzLT+9WEVHA5w/O0BhYshiL
Gvi3mDsPc5TAFcd4tZjLQQpbxXWLgjgW/3KaCnK10lVhAJ6dul2smu+XMs7GFEUT
a2GL+ZSLUUd7LQV808ZP/68XCl5eN68n0dnW0KHqzGZU+yl8hnUez76PXaSAw9T8
qXYMpaHWIvhTFhn+miqNHtVfrNH0Fl1xbdpJRS31gJeV2mAG86/a3t0YIGTCTkqA
nAWxuisBiIH+yQZu/vF/SrB16p7kRwD7+EmXxO9ndUmr95Dcc4dsBX04EZWuSR0/
ta3voTOhS55m6wf0D04XSOw9bRZBzwJMcb8WlLmTlAOXg5VjONFabeIIi5tsZQAq
+gxfIojrc3pHe9fUN5WDUe6jAvl+O3jKdO8yBXGBHDx5gNLPebG3cc/VSaTtRD4o
VPB9/78DW9tPIenUA8mslVEX6LrtcyCw5ZY+8d8eSoMqrhD6kVVTpzEasaUgHXQr
pFlXW7MOLaiBzlxnjx6eQkLGqQI5cXBQHToqqGTkGHAT5b04zuk9M1fQfTjGpvWV
4N5uhfa7SKCKNU/Jje06iM2ayA6IUtzGzwlb16gMjnDb8wS8HALDeMZoi3KDkGIQ
dVzVVdE+6wBfljHFLtBvC5/x+AR/Hz0qWvyJ9XEm+cX+1Z+/MzKamDs/jsxEp5uu
YgSHc2SojlmGzBZEKZ66xLB5V8npzVfTPTI6qCVG58TCKpShkEvFbT3ewUQ8vFcf
y6KbmRRXqw2OBx7n4AQk9HwNqrnth1vtWgnFKqFh7clvqdidAcmpL2yNVfvMVOCT
tdBoNJiyIVYkMLDaROKIujZIHvJpE9VfaVEFEX+Mw4fv0ve829+KCiWUYkbKYT7g
69CUifBFuPMzjL8wM9Hy7y2RXavWgHF9WkNBiywmUoaP93+6QJQEPinHacsRLPPd
EGVZ0wAgtRNH3fOnxXiIIobr2QaTbqB3RW79AVX+tX84KFI0JuUiYDmiOl0uoo+V
nNzktjv4NiolfJv1DRtg0h7vN1ZHFYYZygICpQw8pSl7wUsxAAivGtyvTaICWe2w
x/s3hBo/itiH5QpoGyYq1y+7KTZThT14n4v/Vu27qMyE67Z3yoDN2QY2wkbYwbzS
WFEu1ufOeiaoLqxv06A/OVCXZDJOQD63PpAhMGanTzTALUYbJsgBrGXKIcX5I358
75ROWs511j7o6JHd/uV09JRYRKCUDgD+Hd9o7SdaBu0A1JKmP/d8dAsUxIXg0JwO
r7EWEtQP6NiNmyLnSbDw+41OrrbP4VsOcdEprVB6+gCludzYDITKAwgZRJBPH70r
drc19wz03Dp1SWojxB/0NVxUrCP27B1BDsVc2vwJ+/Hzk5v6D0sgjV+9k8mRBNTj
xVEfuqqAiEjqT+72NiW3ZVvEDjZRvdqnCegYQh9Uz734FtWDLs6Qt3f6TLtplLVN
uKqkKPaVX/Ov0ZL1sgreige0dLrE9yxWbT8pnHUpzWmtTNNU+6lEViNcDqvAnFuu
GldIlE0+YY0mAQ0HfCxM4azGY+k6Baw1fp4pJj1Vn0hVkQ05fwypTNe10pFlOLCN
QK0tGVHRDP0BLVjnP0DHB2G6gWssMCGy62RkjsTbaC5iiBttCppNPUEk9a470gLR
ifZwEz7DhdYrTIUY4ZcoGx0yby2L0uBpusuWmhKVlHgmhHfUe9E7LYw2H72e7kpk
UA0ZwDv64+jYqhJqovIFwont959Ot77lxHmfZ820Sv/rAmnCCclYWK/Rc8TYCC0N
nZZ1uApcXnYJ9VjUaUCy9DZ/3WNEvhgmOY0k+zIB+pASyGd7sa8ivFbRWNORuL2Z
LziQfKnv8quj2lXGfL7ZvNzjDlIScnFAGkmrSH09xpS7sT6q630qwS1GPKsA3HUB
nvAEtzhcEnbV3Qy1C5TA0bPUNptinRVzaRdH4/n0n9RWsBR8H83gm2ssg/XV9kjO
Rq9c+ly1lEnlRwkPVgh1YMmIdekTzE2bF3NyobAMvMMcTFMartqRyhHD6CeFAyIp
JRLdYhLZKTokYvISRAJO8FKqLYrPah6JUW+s1LSySCPqJqz2ND7YHF1/VOhl/4P7
DG3bT2dRjIBelqsfGM66GIrjFEy/CHkxnwA6ksih5IcdSCuAXHi9mrw1Sf1+981H
vR8N03K25XjMUpyeGVrRuEyMyw5jdnsL+F5vZAczKmkRI1airSd+tiUi0f91s44Z
KC6PYL1pwL5rowqgque2qz2RInFWZ3/o4pMKhG4358cq8AdvNkJbbuSYm88qu95A
/aGMm9Ly+C+FQrcWgZyc4MpR3Ey2JDBRRYbV2MeGyxRytmsmPtVMrV//Lbm34KbV
vdjZ5v4tqHVTqna4GCgoulQdewkE26ru097/aJWXGUSkP6RLyLB9ipRsAHfVesQW
62qa6BLT5D1S2urklcaThqYR5M1JsNB82WLla7+Nx+lpShfvjWqGEQIPgcfT31tV
s8b/++gbJTW/yYW0A3AE4+w3yTuW9GO44Cjyzn9eeYAdFX1Nl5d+fVIEA700v0DO
ykxzOnVXWQQ6pXcFbT7/YvnIqjnZ1SJCo2vLihqQVSAmVNkNJFHzgr7MC0sbstLs
GzoYb3IHwuJcFNwH3MAyolDHPnQqq50Wz5skS4LYiilO8kjI0wd/ulVSjTvgDH5K
MXhnd01Pds2wXHU1Xit7hwi0BNYhvPzEiQqSIE+cMQPo1JPIr2x0Zcl4U1iwKPlD
o2w02rkvC9XmwqYe2M4HnKIR/Te/FSfPUpksAu3t0fL8mmo+WX1K8yuxKNO7JnfV
jLgBryHoAenk5pMdQWPYmAVeNeNfKQKXWGMwU0leL9OWYJGmOInAzFVlmX6wgEdp
CM+W6kxr1oGJh23I93kYpMz1qT3RkeZFGxp6Q5P8ehlSLQsX7NQKYpyFprA5/RO6
g2IxC4VEKbGHYOL6k0XnN0umR5JUlqH2wRoiMNf2rjiA2QVK45RbYnSP1o8nQk7L
NWv/4yde0jNsQLRr8DUvdtaSVro5a8FpeJO4N8sdVQPuIG/P6Mt6pe1758gNmbuY
S78khtCk8qC105poY01C8/MMrd/ByRZVli8L8EkKPbAnaRMetmXNqs0Fbg3phYmJ
E9FjpATJHKUIcRIQA8VZplZmZNLjcB8VH0ZHyDHBEDc9woO6GZzwtGDxwHnUagIy
/fNXCib9GRL6v7QWixTdPXmATmwxox9N00n8Md2xTwvHnofBqW29ef5L43Numg/j
9D/UXwBQiEafC7KUAaMA9Uo7BNu5gfMLq5YU12ex3l0K6ovmvgw4pamCbDFOJzfb
2DmSWoCj03Gpk+bYJfW/rE8yRB0eHTT1UZKMmB5S5EMueXxdEstmwObL2L4h9nhJ
4qwaybR1FfsjhkXxbbHDea4t5BeR8/esWwsZhO0ZFstvajvjH1HotcNUNoWdE+NK
2fLMBo0JKysh6fFoAlwFkj14Uoa7p+iWiQmxrv4BmA5erh/R/WTgqAqvUSZtcNNS
jXe48956jWvAhtnFZbgKQwss2B1p2z/XK8gPWCruXpE8hTDzhmpdWaKLJ1DKOtz5
gjsWAxKy0rqtR90b3sLwTy0ytQZFDZZAo0Ymn1qcG5ThEekWwT5Y61jkXel0UJ0p
ro4LCFRJipC2e9qRB4Nle2JsCLCOxDG4Hvfzp2SfO9O1JmQtssm87oFbrFVqOtH6
6wo05gOPAIjy0tGr8J+vHI4/SSsQUGUzB7Y0zkPQL2C8GnFb2bCMXktDZa0qYtrT
xrSqcjfFPptxtEC9TxYuzc1SFY6itmyhAQ5a/K+sh5Zj5iYyqcGI4BUBTkzqjaod
5eEXOHHNwBpzg0esbAJigxJthkWs7cTzQcBotLIA6Kg2ZgBNJ+/le2upI+z/ba47
a9U9xFJgi4+ZkTB+AkA/1PWEIViQfhOrnhLVUaOtnH/dRlKVr3rUt42hx5Z8gQuY
Krqn0PL+sMOEbabdGaemYBFlWtE0XYdsuVmdTIsVyIcRSqJ7VAa09zX7fmm/dR6b
FkGepD1PKCedze5566gDPYZCQiNgUibYJC2JahkX8cSF9kAJysxlPD4ITgmLubpK
eQK1z4sVJ8gAQvvYzBCQumT4DMvntTVIgiB6k3NjjQxf7OVb7gRPlix0wy+OfQYI
lMYjkesBT9WAElepM/HTTbbLYifc9VP8EPqqi4lxbg1GCk2q4toPIwx/+ZO5myju
UVg62v/II57liFN5VmnbZN4m6mq2Rfqy7IaisQwrJjFrjlFdcKd6IOLcS2M3sQX/
AoRhvfqHpzJ2GzQ/bWp7i7jw/hmgcjKTFTZWCjIG7xt4/Nck6XDtAiW52+Qv854u
EwSRJe3HEsHcjyTgDSm7nAAzkUXkAxQLZQMWXul+XSM9YF0dSTOC5QKyuh+xAOD0
LGrcr2F56Qgkmoy4Gzb+7lKbxZ7Q1XnuEJc2uJSJQzYCGwktHcbQT/eaEB6zp8mE
kgRcHdi1NwqlPI+x5Ig065Z5fxKoYj/uTdXdfMBZFacJn51W5+3Ovo/by2hbeDVg
yNjHT+PgS5EAeUEce++eowr0LS7VApPyalt8vjW2E38IelYzKvNZ7RXIOzoPyzHp
u1R1QgJvDV9dFt802+4K4v7XKPmPGFKy72vGMFiydXSKB2f+rAj540aPckiy4v9t
igxDis+tQb4pwyR3TUzdnjAoqG1PQ6Pg/K4zIXYi/rOCiiqTiVjrHr1lCN4cn332
HYN/q0Rez0CYzK+PdfKpFr8xuzFFcRSFVVztL5ntfzUzFamaz88nZwtKbZ0dO+6S
eRTcfQNbWDzPfsOUcCb7P8gXczZAzWJQY7hEKo4a/e8zkcIyRDPTt+2k9FFJZ5pF
qEuORpb1fnCSsRcPcXejHyf0rdYEh7N6o6PO4NikHHqeAGBsfsSDlBZ5ThLUywXX
Am/WjYdfv5XN7fidnzL90oOcmIiY9z6Am3EFc7kly3292a4/9g7lyXRdRurPwlMa
EZiuKk5TFRmByGQqX5eeoMhsBlzkAzzx9a9+xDtOjlv4KSFnh86sGcuefXqPPGDA
MN3efIKx64NgnUID4YxbaLQXCdgskIn5R9iqV3nD5Zw+ADRpLjnyDRYofIzkGgTk
iaoPRsX29EYRnvRsv+jQqQcWq7ZTBewqWeGc1nYhgrud2eqoUJcthAZvujhMEYJA
IBTIl57ySddv3Nj7Md1U82XiCR+b4gAejtfLqw152dxIb0plKjYNAQhJry4To89W
TZI8DEXfc4ps0rdDL4BtZ2O2CmK+iPUq6H0HC67WVSbq/5O8ZuFfwAPB7fVeNZ/W
mt8hrMR/74UYHtxK/dYu/fRsQQheyuSsrLNo8wMYiatPzGJ1rUoPMl/3TB37Ih04
vLX5DPPnuyKsM3ZxskBtpVCTWknWtjqajVAiTAmwAdf7S9xVMAFjKm0lfgwpbh2k
PyAssuTikiQwFzIZTVXhjQfMpWYdyg5kRQz3cp/NTrG+hwcjnVMZxqqmiRoccFih
085bSe2Yg+NLOMBES1qh9rslhm9jWiYlSmqOWpxX33hz4FHLHkQwmpHZou3SZBHB
XIM+9xNpNrYPsRzROrdW/EFpOpN1V05s5Q9sVbkATEImQKRoKA3aedV9pReWaaDK
4BObVLVygQLHHd0SPbo7aPPnQ+hxjwY4bMDF2QcKv1QS7hwqYtc++huXDw9cN94h
3CJYdT+5XgUSyqqY5nYWx8vZIGrPtsthrJC9VFf6Z9ybduW6VeOny8hm9ZbNVHxo
Ohyn69SezFJMEtlLYCYqs0+xMl2ecN0kFH+YGNeg7vK1t8thF7QchU9FY1VjMsQt
otX1lQZVJC1EtXeEVWrqwjp2cmQpYi6bh1yRQzHtBj8FBH2Is8V1ZuR90ymVL2lR
iprxcyLRYxekhIm+YLTeC/8d7Wkfs175ItgA6jD7XR2780dN9jsShvXvKzhDoe0q
QVrJE14v/EK2h6YGCZ+d7ao9VWpC7wVqfq3+CNUbqFn3QPzL5xLFIaDmvjjn5X9b
tam3c5vtvAV08dsVmHG33g+xKTrgxggaE5ns2HWwLuKBjeCr66Xqtsi9NtjBZK/f
MVyrGczCBmNIHyA7NUPClFklYyw1WH2vbh11o5eY4msa7AeEzk7RNT6P3PSxgjpZ
6WJW1gc0JbaLLQraOLYtiks1WKPUjTQ7mLaANtgyTGcOL2nTeKVYxNUFT+z9IDEN
PemH6Xj9JQJ2c/E1RhxxsYruT+QVe85iUqhk17HprhLK4ERED3TmGQFH1SwO0WA7
vnicySYb8rJzUQL1SPjI7PzBZM/GmtJEDem6OOJKMEj3BUMNZJMWSveYTfJYKydd
euRo9R62O7wu8FW3c2bh6fpZtG8M8HoZMABBckCLBoy4RUVufMkySpumHISy3qRk
YV6Vcs5dkim+FUR6t6z66/s/tDtLRVGahlt5bnv5qltk7zb0RdJrxFdL+NXDywUR
vzMpH/k/lymqnHVfRDbgm+FPfvXRkudBJLuk/CqlnGgFlu2cSsmPijo2OFXgUcSU
itTRsqddbY76msVXN7AfVZA27ArJHY3Ohg+VHUZl4k4WqYNVcn8IuCeT+2ID4mZ9
DaXjHMMAdi6ddmLuXjOXavqe00voGMGcudQ5ZdZHl1Y66R6NW/bSslQtSb9oJt8g
ZFBRgEj7uPHe2bwbXGzCIL0s3DRZd4CPeIcccujbZ3qRAEFieVZGS17L3ZjS/xdP
h0/98bcPUUENnRa32/lgo1ZH/ltYHvvPrj+QfHJhYZ4eh8h1+xIS8CEqLYrlID8r
nD8Yt8XmMFZKRqE0u5DNA6qVoTBX8kMOO5zxiAlfAs1QPc2dJS6t3NHMuotpVSmr
+i3pfWEm7wr++yzYnRZn7c652lu9/AbfnmE/IToh2xs5pSu5lHSID2xkZUDK2O+T
SkEAXKeQbXvIzbUnqT7DBZWTLLoBxG5bF47NUkFVfGO5NTm+rZpE1qOyjL9IslAU
gScs2GcW8H/uJ7XuT2MfK+2PVrzZt6LgZNJnh5iipBzhjFVFN4bGn7UynqgZqwE4
LkgGUB4zA5Tk12q3rsvF3PW/2yZfJK4FuW2BPgGzpfkHFaHYReLCW9rHGhFMDk3V
K/IqRI6jLn15Dg4NKtXyvX5WgyU94aHVW8KvvnOWAAsmUq6uyuRpAzXgE262xnjr
wSWo48KoDJWFXB/ESuVqDnnfPMmn0pXoHpDmjlJfajTzKJGbXIy4eNV+L6tlr9Mo
+CnkcRMkWidm3gKvO02yzuMhJPCmhPTrb3OOK750nAfllAk6RXFBL0jKHyqRyXAA
MJcSQnmp3vv2FZ8KzrJXLbGU5YmgMaNvW0a5TAudwPc8ve+DyjszQ/G4C7y+FkE2
bw8t41p8Ay54JNqLJSDQnrjjqI5IIOrQ4i4uA0xJ0h4DdbHsuDkIiXjsfnVla91k
iAcYBp7ShNh7tXDjIdSBxdoCYUMz1l3LPnPmlCvMNYNxQvS074ftxuCkUa0dcfin
IGltBXKvZBdbFChgsM/43jsZSXAuHyRMj59bJecwkB3tjyG6MSejo3N4if760ObE
70eaIs6tHp2vKjGynbx1gTJ/BNAcQc/krvQzTreI5Zj7VGTQVhchg6o90IH7CnEt
0cw3v+1yM+uY7BUb2+P+r+kt9EkIQvnD/S3f+kWgaFM9N1TNnr4o5EGOfgv6v6W0
d1WUvuGhVmn/jxkQ1Pd8u80tAKsGBKjLwmP75bVFMRCyZLhwya0P6NPCVh18eOR5
Gh/XKqAOXgzk5D+2V5+cxTdQk4uZtJoWkh+kMPXGfeoEqMdTqPSCynyHCxvohSFI
B6oRZOkJXXC51bXme7foL8Xt6weVsX5wRTA9iS9cCrx88PMGScCHJwaCh3d5KNbt
6deTRUkls7mSpNDYvfIGABSSaMOYUhESoTA6BAcP9ryiDOY9GehoMakNCcwnOBWr
xxRHnuJ90T4FFXqnMTcw68Atlp384QLbuFFE4cePrpEq9IcrbGiTHfwyoKjoHveZ
/b8dZwUqEdUQnPZDTYL6nJSpefwI8cgHpT/l6OFPzjfoqrLaEya3agY5mYaBSi3p
20FhcvxupJOI3le5dF0klYzQj5cAZ4MvITyOIaw5untjkQPxqnc6KMFGjuNvphLh
`protect END_PROTECTED
