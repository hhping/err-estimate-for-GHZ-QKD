`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZIS/POUdV7MjbKkjR+255gIBIx83II5Iu1FGTHRjibCy/UXh6nPWZ5LTP0HAygI
rcB2KsiAEYHtYxNrtx5Eaaj4Q7J2hw+ZeBwSg+PqNK9q1HHgZmaD6t7A4alovOH/
iEdbxt3QI7l4QX33ZhBDFF/kC/SOBEvTn28bNCFa3NCSolAMRXAtgG2IbyVOybqY
w53Y6hGmpNJ2UCRevxcO/miQkW29srarQQxqR2Kwz5+2qKgmBXCWzID0ONVmEiYi
OkJdkUsoypnNN3FO5+FCdVadY2qGKjUpXcSo9GpvysRP90UmlIf65z0Y/d9K+3lB
X8rZ+TgIAOwaREm8Mc8weOeGwtMLDFDD5rqVy/07y5R6V1i4dfUtX526YvCXA3e8
2bnNOKck3Bmu225LbQZPmUQfLBUyTrkyOugAI0khMB9saicbdSm2KOSyK/2bZ2Cz
r6bLn6IzDYTD4as45HlGLQ2ST9Ys745hXQBvCPk4AxLxInHiPTGty8MChboM4QCw
mnFSmeigv4NGLwnfHQUD/BgC75v+GSffsEoR+uTj+x05FXeP2gAxO4Hx6xJ76WV2
k2a7E/pOzM4a0/UzNFH0j2Pn98kR9F2dzqW7TAZ7XqKiZio9nnI+BlY57a0As7wB
ZItuiPqrRWlgWD6ZJ4LWSnXFDd1aH/BzZorJGZrXwweTWsMyG2wWzUwS2JMQP8N4
l94TZ5JvUjbuXALyW2T7EUtnj86gkHWX67B0w6w/RG1/TqvtaWcJgbKr5gjbCMG7
Iz/jvTVEB3/Q7d3gHVcjf2XcliWsKTk/i3aT/Sup8srpf9j2H6M9CjYwIRgUJL+v
IzuKIbX14oKFk2Leyva+1nHId9CYQOI24x0Lg8QhgCPuUzsF7HU1RdfoX2siK2un
HcnFP6Nl4JZdeUOIvCzsvTFvdVTTjUQ6ir3Ev8Mrw5m6EQytE69i97gnuywxUckG
hv54QwhaTpeH7NZDFvtjzEd8xDugErhhUbVfd41OvqvhKNV5CujzMQk2ax6BEtX1
PMp7X9U6Ko7gDVSPyWfehOhO8X84eO4cQX76klJCmp3ac9324tpuPjchNzaJg8Kb
nI/YCwteH8OQJ1sxknPbzkuEpqFH0Dlu7KNyXHyyHI9v2fCJMez/kf467kjwm3Yk
CXVVyiq2L7K322c3mQeXibpBumKbG9H8J/O11lIXoHZmKrSaBLu0xAbfbVE2aOZH
+e+D4XKs+CTkznYM2/uGgKTZ5cEhYw0+eaUF2Qgu3sXIKiwiyznHW8oBVBJ3CXux
O5WD0AB5MYAaPoMxFd6oyAuX8wXfCQAHpg6v46A7KdT98vi18e20+BMACEeZYAiD
b5wSjoWFolYoFExwwe/4xIEPRVYMT/NfKuK1JRPwXfJ1Cg4NLb59RIDb3Gbrjc3m
JwGK333x1EWlP2lgI2YCUreE3h+5vkcfyeJsSJmS26oFHSO6hzdQItATZ9xiFMmn
RB8/58+zDH7N99aw+/sREVLmD5oUc1Z+QS/axe7mq/YLdCpmupwCQ4h0e38s3AIY
TVK4TNBAcz3zQDs2BMCv/IqNdXeHSUknfdzv+zKCEhGypS+XvCGM+JQ70mN4wxbf
Q7OUKUxGu3B2My6VrQPd3nmK0w/PeMIRQsA3K2AGx1KTeDrOmGhuIRFlFPQTIXtV
IQHt+x5gomsPVPnWdRQYTXFX+ld39W+Z8tHpsahd9lULVSPSkS1kLM8NODCydfqh
lPw9ufeQ5CV/48+gMxRV6hoosOfLhd1qtLs6UpIckOgbTr5eNdvY165dVJDVY+FZ
JVZziNm4zjUA8qIkpMfufaslQC2uxiHgZFGuuiUHeSWfezIJWOubtC5OBWQaIate
GF3p1NY8amcRQeggKGx9zxYCyxLLczNbPTruX7FblvwbdS8DWf3mSO7Fhn+YqtzX
PhJTuU85AbJAj2kL7dlW1hAj22FmfdbrOcBfcHj7Cr9hiLp4qi0HScOiK2Kfkep2
ZXze381dLSxsRuiblNHDLg0uBAwcolbAdm3nBdeqQAnfj1iooK/pTFx1L3F8EzQN
5tJ5bzG7ZsNxrgHZH4J7bVpVYFLLETadIz1zBM0E2k+okcL8Cnh4q1jbbRdE9nVE
GB59LpLmOVgjvcq8t4CHEy9vt+IOf7Nc+IFsADWqCYP1096sk63sgV89cZ6Xs7VZ
tI6lUmclpVZAPyAIUYQCsWWjaCUbWS4OTsUl06Ppc3K3dpsWwzrA21PepyU4ZKdP
5MLErjKpIWQZniJPrwVptcBpXL0+IimP0lqRnvySFZhPj4ExAW0UrbJv57BWF00V
4b0QkQG2TKSZHuKyVUWW2fKJ5OaL49pt4PV5nb+kTV4Z3M0h1NiEcfqXo81/DW3d
E+S7tkXKlpeaWpT3GeGIY96Hr5XOZ/rLKwwHZz2l1Vmce/IZz0CjcQUn2ya5T0+Y
QuqzfZ96c4vchdKsbGYq1swr6qHmG1W6cSflK7za6Fjl1VJ6AwdPHOTustkZFEHt
VKpXlKND32xLCR+iXItDUAF/rg9MbINCs1KLMhxaT9/o4N/cXAH8nqipsVWcuj5g
D07rkGp01aUkYVQSa/mb0hicFtKEVK4f6sztOiBTnQwZTZ0RMrhEiehJqngvkSas
vXyYFKk8LTNb+RDlSgwurgGDr9v01rCODaJP9X6JQZRUJ4ae0jfUC6EQ7jaa5tEO
5VWGM0p9mYvmRLko4HGJtFKoszjR5R2RFQqSdWKaw3tkBi7L+CVjGUFkecdfH8vf
iTWQiw2Olht1OqirspHR7pcwPZGFqUkHNhPr5KBa+KPe+C2kXUsVe+4bsV8E3EZ3
nnhZFpjgMm3jb9ko0tG4/xAei+dGkeY6qqbDqh4ycdk=
`protect END_PROTECTED
