`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUHU/rZeRKdlHv8/HcFlru4jF6g+tyiv+1snbhClTeBDOddplQlV0SqtwpyraDfT
iAT3Tlr41/KILryn2zeZc7rZzBi6oYwNJy9wz4Pial5zI723TYK5qJa5mShY8zBh
J6Z1AYj5Lz21MgSZly2ySjm1JYumZTFWGgbxFyBoy9Em/3SiQQi+EdeVszYOYiHL
pFYuAnFBt5+fNJBotITL/Ytn9znk2Lgk61U0ySzcxijNTeDcIhyh4nERjzOF3hRP
8wcqOShHvMiVuBtOjOLct7EAlBvfzo27oyIwO8dxvRxfc+GrfIv8M3quME+BoPjp
W9hJuZ1ZfHUqRn3VnUZByXVntLc7Cjk/hmP7Mtbasjpy+BSbUg5U07CSjgJCQeHu
+Vprr4Aoud7rmABsAqKhAcSSWQtXPQ7SoiFotZK7n1w=
`protect END_PROTECTED
