`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZq+ouuQtgYSZmem+lDw2UNg0/AG3FZmg1GOVUC2LCOGZOArRfl+EE6bX5obK0+k
2vPC2N7boo680Qn40F8mjprmrUoj4riTmpI3owdi2KBZjiKvhKYzdpyknJ38+EN+
woOWlJUQYCxvehNsUeDM5TvxBcKc1dIp1JFAlSV+nJLYDwnarcdu0FwiRiohlWNC
sZFUixzFd26xP0qA3omu8nGw0B3qI6VAyZ6mXWz8TFBP9krHH8iA+RCGobpi3iTc
C+m57vyiaI6g9garL4Ox7EIeKdd7EHM2JR+cwvbkhQMNwhcgAP24/RGoPfTtulcH
LwImaJPGv0OeyOFAO7pIBZiWF95lF6t027+IDawdgFNyy5soGC6StLlydm5DljXO
xRo9Ix+W7RCr0mCoBUBB6kx80DDufuOUINsrKnCHwftvRJZovtEKtHEZnittbVAe
XoFk6V5dq+vFLbxnuEEWCsD7XpWpk56Ex+GU/VYEnp1vYSOciKTBw9IpMuZMiPx/
XjPzRGuufeMxh83c1vU7yVL9DUiY/dp+Q39gTavEkL/qAVSOG9AP0h0WPiRKhZ2c
Fzkgjjcu+aZmDuBUSjTkP7IvUrmexrIIIYisUmKJFwTCP15mUy9aIpQSgZeKpAYT
TXcuvQEFnD6cvkZHLz/XgmkccEXemt5RrOkHOPJKPUsN9raA9s+ccHe3ispTGMS4
L4qr8IQc9G5Cq6a/g5wKkPcOBSgYRrFs9fdqvhcZFKtf49SpV38+I95Yx8gNF8A0
qibvaS49UxFZxmNMpb35qB1+JHLN7ZfR/ayuJwwT6Obj7F5RX2nz3sxxkWPPUUDZ
tYjlNLgUbtNlN0SHgXekNxIBeGqZQorbRGKUPUZxba8lk5PJ41AFYDfZdEz91vca
kfps85WXKiENx0WOuwgeqxw5aMcMIoX3Im1hvt4byTKVcff0izI1o6il2nXoqYAe
rBdua7u3fclPrBfDJWPCYyreBNmyvwESlivcho5hG5bHEbTUS58LvDeDTIq36zh9
BpJNnocyrIWnsZ/UMFbmG0LGqvUjThJwJo6xCE3fYk0Li6WaMabPQh8obbgx6D4w
seZPwrmTjXVqiC/mI79YJYwsJkDbP0RfGenSDpXdyGOZwojdE3GyNtXaNJTdeP0d
pcPGkGGNYulr3XFzNNwIV9+Aa/cnGUfO8Bx71cAlGZcKvTimuoikBhYNmwdBAJHU
1B57ID03QsTBGYNv9qMsdMgGXMQcZ5wYv9w/cTI8fUKYmORw/1Lf31BTvS5wSMNj
qGG0unjQMsHtDs+nOgTe2NzzwTcSjRtXCXpJKPWnGDxYnGXkSQTwR5Z9VX63lvnk
7m/N0T3fAC7I9oJ1RJPwAWBYpl40hKI7Synd3V4S/39F547O++9T0797Cs2TSt9e
mOwA+Exe1F97E1Qb/wrbl/u2KLo6YM9mQ+IF+2BtTp/cgZGtwyRBR30ZeTwVzGii
+95sUX5OoSnckLDl6Hw+8UZFJXY7EGljuEYqLiqgiynyfqbQXDPUwkAU/jugU9ki
EzWVlhNF+FGQ/NiJNc+/ulf3pigVJAy6TYBwHC/t/bxxTvlXFX5xP1YD0TOO1ZC4
v5pioUFFQ1GlGaY6IjQ72Tk1X3sgUR4PJlPVW/ThluGo3vc9deFvvblC6rtwGtsZ
clU71GO7TVqdZhP0wbW8xCGrabGh6C+z3VENJwUYNIRHBjMMFFbA0qYXwhtUqEOC
JlRU6J5YwwM3znOo63S/avdTQa00jmW4JKaPK2H8k3U1YE9TLUnHYBpSWGbbqdZw
3KljJnRVMlDKAgcWNYLU3Djz94Jglntcuf5MjClbm0weliVVJklVFsjHp0LRQmdd
gqBn+jMz/1HPF77unAav7bhaqw6MX6I4Bdx5M1mf95tqw95yw/33nJkn30KMq5+w
1vrNqb9FZ3vVEHAy5X8Z25w8SKFTPt+dmDui/FwrgSYdTNeh3bO8vCNZytR2cHQZ
JqxZjRiDVh8F9kOjw2WeSUaMddUjeZa9RC2+dTu4Dp37VHWtdV2Oq5G7tVMMFQxJ
7s4iRLsyqWaYMQ1PalnSQtkoyhepti5tn/wARkL1r4REhDlLEyq/0AKX/dFUqK/P
iemA0Vblf8hOTWoUsbiBS5YplSnPSU2oHw16c/cbt6/PpvAoKjylUnK4KNrUloMz
PtilMsWPKYT19z6wn9UX0Z1dXjLLDLs7Qd3q1jDaZ1r4VY38hyLzCtul+xRP87e3
jGasW2RG8G9VlbE93N4qaeSkQpUcwsLVuei7ff1DiIgNMz3az/qvyKCO+dQhuaUx
KbPslWIST1Nx1tqJMQ8KUzNzgeT5wvPAx8Dec0TO6vlzODUazfW8+i7oq+Qxof8R
G7koABTtUSz5ydN0JGiE8V8Ebos/FnhtgCp7/vwMNY5QFUcM/uUtukle1dzI2ChR
q+OWm3GxV39eEffjUAwIsK9TFeenCd/Ad9gQhPmBLhPzouAJFduMqb1GxBJiyIJl
ak5Wr8LrpBA3D2tvWscqETBoGpnuuyEhAEOA7xUaIfk+ASWR9xzOznMpujHYvk2r
eH52FYVGouO/7yKRMetws7jnOM0wsf29ahnGg/CaZY0oB8g2MGFRcTeLRTjHeb0Y
ibGwMTpknPqRg+LasJv9DzY6BJNBSR+No5kNA9bMs/jsx3WMZzQdERBVtYlB2oB2
aWjHUpgHfGbTofC2460heWRLYKEhr8lKO9j+yz6dzn9ou+0abolBCBEJQV+MoSU0
iEa+uORJhnWVrwmjF2m6+/8D6DwyzNFlwRFYdWgkXoJzRgiD3dXd9bVJm3U732Pq
+f5Vz+WFd1RFoPMW6c8sZekAlufmw3svVezw4orM/3jO3QGN6PrM7+tEnZSGObPH
Kzy0aN4nRCAbvpcUrUFIR3jAhD9+kpmfvwWYVuDT29EO5c4FIY2eF8pM3pzhfPwV
ULy0ljo1QXJ2d9s6zxHBSCjmN1UkkqKonTsfiAAN9cv/emCbt6mMOKk4OS3kKy5V
cXVEMN5gS23nRHVYX8DJgZm7eAC00+TnxvZwnt0ZsQ53kdMVzfU+u2s5rSdng8CE
4q0snyMb/8kdCzIyLEUce6qTXSomxUu591/CQ8a/noQnotvm4VdnIxUl4rqt0FfG
CeQJ9mSNyV/TVxwvzYCk6mBk8RUmfKlSxk3+HgassS3P3VOKJoknfvy/3zY5N6gQ
yLji1odxXWdQkQuslblAdCN44Jv+LFO0KJQQTlYmj28XTbEfv0i3UZnBrsMB1j4U
HDH4QIvcZxjnzJxRPRrbQsKnhi8NZqA2hP3IIagF8HcaaE0yVKKT6ORt4SKFTYm3
oCe3o/ZdIz/RTRFZB8gGBOu1ISoBVLEQmz/5CCsr45uXYVGlynPVF4I7EPC9l9JR
UVJlyVmZXUBh7ZYK3O4wwRWo7fQWphyPw1UEUCbLVgqNDAb4ObsXFJEzrR+RxZ12
w+pBaHOTgx0VYg6qu3uygT+y0kL3TbkODTGYxTaIYhBQ+VjRZIWja+gRx+4k65U/
WayhVdkI+zV0Uj16Tp6QBL74LKg/rSbJYdq+qepSndE=
`protect END_PROTECTED
