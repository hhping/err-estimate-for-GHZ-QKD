`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYngj1lhvleqljnICXo/XHgSRe46Pv1cBVy6Xc7hpPV6AYVqF9rqIRf9xD2xl96V
LI+Zz4nsmycpzHHJylPZEvsQz9lX2/XSGtjNm8Yeh/NstEzy0C7TSKh80CleLm5s
YKdjbCBkTBf/r81uhm5cg5Sog++7eqToLFhzVAmBGIseKVWqGsgfk4GaPsmVTCZI
/K0hlPtxmLR2iD2mDlOXOTK+Kq8EXeAU8IiBKMAdF1KAi/g7DMS2QKxQhaToNDqq
DU8XpknsJ6sD3E8r23VWdUvTpDTZxJ2964vBLOeNDA7LkAN7C0/ilPd1JSOsVAX6
NnAKDes/o3GoQgkpwffZCkD476mL6Jp77bLTrcsdmF6F9rLe2jz7VMA3CYQMBgxh
UFgY/OvtO8b9kXnnSETiv9CElti//Oc/OiHtHQke5Q+IpxP+kFAUj89i95AzlD0T
ZT02HRtqNoJ/2ZquwRJ9CCYXm/0ofA+MduLICjLkccR+hWX0XFZRaWHhOf29PX3g
2+4q0PSaqOnDOMZPx1f87wJRpYqwzjlBwj6yn88tWmbY2kk4Dzm50uuzz0zXwUP/
Q9l1SHj+HLdolYf6Kfoi1mQcvG+dcshC2iJRbDrSsCHv2YGXaZBC9JjcztvLhNbz
GM+eXgpOokFAixlYgCPQ9QxD9pu+aMisqGSx14l7iqnk/s/v4NP8HQRRx9jAI70x
3zQtsOSLM0O9eRCfDiyHpHXlM3PODdNtl56bY9Ae56OP3zCvdtzBoPZGAqrqwX5O
LNbYeV+SeBL5Ej+zH6kfINN9egWoEaXQici/eYDwJxBqEVUVXb9gMpatSNBAejRW
Cqn1+zjAesLaSE+ueTbcidB/e7+k4P/IcS1LrPgBsuzwvk+4NiZs715bfcJLm5o2
T6HMtbrubgySfNfB7AYRuEFUY1mkE3LNGTbtAwG5I04SUsLJkGNX/nTFEeWw2jb/
Bh7/N7USqGoMB7oUMmnLA9NvN93H8iy8wYlI3Z3WB4OcHbTzoB6qQmXxj+axSGAm
ghLsrDWOXquu5AkauUq/rm2oqDVvrss1mnnzMe0Ji7QkUYghZAirB6o8NK8N0T4+
SdQMble3QZx/FLkyCjPEkibyA/sSs5GR5YaEq74Yo61k5LGWEPFtUEJ94hmeR/AA
nhSRwV7GzBHPcvdaABcjyCrBkIYFlja80JV9MM8Pge03NOADceluQkypWTCEl6G9
XRC0HpJgr+DDg0K9rLaSoAmF1ZW8mbXIWXiDCokQFg2cGKeg6+r2rZaplRblnEr0
TKe6JcuNXPDr5zZr+ZLxZErrVLRKdtxFcvxGdVDsOcKkNhce5x1rw/sppobl2KBp
k5dfzq2fXOXqlsviOfzcs9YLMOqrCtl6o/NR76EJ2C2t2OLbt4IMAwyfc9kWZ6ZM
Zeut4FKjkRGzjuD3hPgG6hIuVKiuO5lNpM9VS+JvtVzX7q1q183YHgx5OV3J7wC3
/vI5Z/2/eisZQJEfFibALqgCzzUGhXPAC1UHG3ip8T+4GOCksFQrHp25A2WbNJXd
KzMio/wSWWnLlGXBBEzrM9f93rFt1DVwapb0lZza3l/QxhbOz5fytgTN8FxwLa9t
R3JVMhKu/ZaSoPad8FeULE8b1mgWom270pEkLJKPtiCQGdQXtSVAzB915Y2SmwKI
uicNHbqp53Ewgo3VeUJTr/lQlE5ObqI/0rp9gqGKXWHCU0UkAwjh57uuQPpUKvX4
DuOY3DrYdUqcPzQI5sBYnU5x9TmMfrbA/Ku3D5L1KoBmHgJczyjD3ECt9YVsV6eD
v5fpKa7mdQS4P8WrCOt38QLEjEjecCNiTafJLWhm3I8KYOtsiABktSKx8DRoTM3I
BER/wDJvCX8bKAbjDp4e4VKUC4YWpiz7sXgjH2+kveFGCiZCibrVLABYInlTzaog
2XHHNSR/m1nUepv7tgBFxMkzvEgMljo9ULm/lVJGlbguwhlWc3/ZVG6RAG+4s01P
pPpKA8ACuK7ztWE3Lq/K1J71+eq9wTC1BppCb8TLg1N3IIRIwzjQKtrZB+sOuLIR
+quq6HQGE8kYycf9zLd1Cna/UnaXJTXgdcfYzFS+ECHyjJSErcMGZ1hwKGf5S7XV
QLmscEqMlHe/EBcC31aaIBa8z/Vv0cD6VhUDhCVl4Emp3LdRd2TcyFVnB1dqNNgq
jzR+/jpDQAQTbUcWCwnOsjYgUZDLOO05He5M0UQ47lQDcKoX804cg4xVlxfe0oqY
kpi0XzAUN2xTcQlBzPrB0FP1rjYMLV3NPj/n+XW0rrjIQDbddrpbjLcRLTHTPO47
3o900jo1NiT7PVc6Rc2KpUesJS9YW3FMKE1VwUtImzLGN/hiqKQZXz23wOpp9S4k
PATddLJGQbIZ4ldScPDbEbhr1Lb9XMejA6YkaGW/hNrkTAOO0wzHFYDBgzeB+dM7
Pm8gIAF8dSEoNX7sTZApQra1feOza6UbmO2L2LwzqdUVJCKPwKVIfOAha7ZfLwVS
AeeHunkgMG0o3iTID+qf13HlP3Vjp6qe4FdOjohqZ/MIQKwtYAfFrlPzgrggr3oz
TN5IbYOoMXDWgAXy86ZQOXhQgpN3ytgVOWhWptrQTsQB4Zelf4pomWKhKDCKf+3A
Nv0CcfRY5plIHNkfVUUxnWrn0f7+I4qkmwU+qzLIAZaalDo//n3Tri0eu+jBTPP+
3kJ98Uj99z1w2ZKeYf3vh5aeVsF2+vcHRScC5RiZR+E/ncxWF4jeI+gRXx5BIDQp
dL+EGELxvSOVc19beY/pbg1y9GFHpeUgiuS4gnM/ydFhx1KZ839pCgkxpePexYoj
XI5TsP/k+EATqhpCqJ9lW0GR+fNbrCi0r5umr1kMmBh1NrC5X6XwsQn3ypoMVl4s
H5yV3Fn6/RVjotEtljCiHuH3wg72woQQ0UAkH7rMQeeXbheBTpc8uL0CAlau8QRR
iwT99wRI6LTm/UsLJSzef/jhqNTDQwIMG469ZNrB7vL6rH1GJ6W/N9CmHNLK+ghx
TUmVcHXCiXdBpez0vPhB08ke3X5o3iifG7fDeqWl0oB67pYnebodd+MYrJPO1aWA
TTLlNrJ7vgqtpGu69+d92prTvNh4ee0l8m6pXgvRWN4DxWMF64r6l0I0qqKI8/iJ
LXqLW539wtWr966DeH/tPU2BNamvJ1A1okjehqXGpXTliK/cvIn9kIcv6YukjAlr
b+R7rOrP0fcQPSi7ATvKcJTWXNzT3IM80yDBeHWsvz9AjSwpIEA2O/KiGMdWAmGr
Ek/ln0NfATxsqCoT/nvSON4rob7ybC/WyGAmCU+JYT0cUlVEcu/vL0Mpfe6dgFth
I8pb32Gsree3PA7KmlZd5X0SxoDyLTYmjGR46C5Th6JAv5w6T33vgYw5NbibKSih
48GH/gkBrPt9QElczagIjfv6cKha8sYgH54C+CKRK8o3t79M/ZJOsA291Xlwvd1D
wBAv3pT39TOWWp+c+Z/GKA5dpo7VZJDNd3H0gYPIYpSN4/7KRB04qik+4kXPWZnE
97b6TzkjCrmvRLFOA3soYo0sWapU58hqhYV107fgcjGujepqAD9G0Hv8c+wenyIc
Wlc+anm0RAZwgy3arGFjibZbafVV5M0APAnZIKl93FMgg84bvwNG9UT3DQFhap76
QdBN31I/yicR/JwrCrshWvAg7oAm5FzWLLW3H3oxd7uj6t0zi5TCjWDwBG4qxJDi
vPr+SKN4ss/a79mg4+cVPFv5NkYwIteNP4EfsOsfgDvLUhmtP61kKrujmBGmHka1
XF3797R4VNnR7rFIl8oVzOKDlt1zyhOOVOGcLmFa/gL1ImtlD095Q42GajT2VBUM
DL20eEG1XNKotgHmhU4x401eJDwJIACYFt4YBtY6AZCT3Vj3L/kVkm/rKM6hHKts
hULlSoZ8/rWtp591JlIIQ5+jGP5S0/MS8bwoXLYFQL1+3F37xigzzXFpP3ATSfJw
oiNw40gFWbWn1SbwyZ6UEfe9j3LMsunCt+g1ztWbLjCqIE2RXUvDkw334S/E+A7R
IdVcRFyf4pGka5wbOV7ydZkXuhE1W0eZZwrv+Zry/+OEiZXFURwbH3tp5lxtqaJC
8HXMNXJUzKNWbB6isBkdAWQdiqVf0U5uuPmoaqJhjzxgAhhHtj1d7Olwd4txTSdA
XcMO1Xac2YfPj/3cnOZuYIfY7Dv1pQi4A89ToqLtRWEa3sq5U1PYKJlAdLwn2zZl
MiGDPutS40erwnVJ6ztmZBt1eoAfrgNaJUJgYMAN6D8lL/4MM8vWMYZ4qiLY1ggy
DTpurzKKrM8MTl1c88M1PilP3wdYqlXw+PmQxqDCSYeCwPZHopkeGJu01E2CbHGT
GgyzU+jQpShiNQTZAW0I7NXJJquQLB2DGWBTPDDhKukKKsg4xWvCYV6atxKDu8vZ
Uv18Cw4py5e76QKZ3O9hbQjb5a/VKmlpnOyASeI26Qc=
`protect END_PROTECTED
