`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gH0Xa4cy9FenhK7cY3mR//E1IMcw45S6CBtgEY5MsKqxE7FrwVbqAv7dt3hEwhoM
cqVQqSrOXu51QUq0A9/uxGFHR24+1F06DYDBPdHSriW2wFPKUr60FGGmq5823DH0
6KO2nxfb+mOfD4Fq1fucAGkBCRssCyZSyYnaqyB++Rr9Mjst//pVNMQP2V0tUyx7
yICqFJCntQgcO/kQzfl35/Jm73/GX6PCTdS97Vs7TgCYITSm8aI7DyveerLP19su
gyPb5yAZd2tgWIfXevaxU/U6vFhmVIsbhKbyAeZBATphOsh6wolttxqDV4Kxv7db
89d+uj1oOzFUVmEN52n8fXnJplLEdN4SruZ+vu/f9SUI3PnkFS2sYPVNjdyepS+o
sxg5uA96lE1mJut8ITCwLx2WNk5u1y+CKRpIVDk7Ck8L2Ehsn2AZQcmtRmhXhrfs
0Fe/Ho0vDyVKEs7Xf3psDb//dosKQYPHU9/BnZBpp/lMo34u254n7xL62SwuW18T
HCY10yDe/K9WxrxqKwvIqhMAfxi9WDlbn6n6k3leJqLZbIh8EAMYy52/UAQ5o/Vb
j71Sm5flRKRiSfIpEcrfTz7ISvLzrmUiwEWjoCipix8KnFotmXXasSFyQIZbo4AK
td8ZuZ3w+sSw9+Cxg39PSJ2NkdFnPxN90DVNg61GfYHmmfsSZNkkaGNWx3yzme7c
xu3VeHKHPYc8GHu9FQ3K4BfBQzop3PInFObhvDNXbszHDSm50El/PMwJPCwhaZHT
jN99ljkjmkaaNUxQ9/8D8VTZ1h/4S06kwEUL44VVNcTPWJsewrbQdSqluEy0YSvn
w+QcuDAK6ggB/6ejya8WjKADUmz424VlkoZhEx89TQobk0kgNKcTrkIw0dXOw6Vy
M9zwK9hVo7Tv3d1UbN7ugH3bHzAfsdfdMSc8gAFnT1qXxHVvlZ+ZCDcD9FenptDG
XoG1hR0LfnfGYFOcg1Ez/ckc3GkTHI7YYkVkxPFrI4pn24GbS6L5Nr9zBIW5EzX2
E/pD7VldX5dLY7mRr2e6+64K2awYsjdHVqU3rfrO5SsgXLsywB3YoL7cNqtOcnZW
FockzbU60qHk8qUniZmImaE4JJt6p2nF6+ZwdLyIsWs3VVpHOTgzR0hn/Ahc/BWg
5DPiwtrxQIw++pBzCtDYthFT5BxS3MdvWmoTg589oYRGZrYmHCmEPLvUfNEQJauq
JNAmx5T7a7d3ioKQii94c9j59xZqoaeVhgeOpSBHP6g3R8ObDvj9G2mPp3ROPctz
FvomyNFl+iiejGXQkOFIWo8hoF49rqEOug/+3gUQvmXhBUmLpPgOyUtv59+DqRTh
Q+oWGvnA+d3PaRJekZKgAUgg9RnYlKq/AJu0bQJ12Otjmuk0WMl7rhojVcAYGCB+
xqX9ldt4MS6wTNu1o7meSjNCn4ehawerOQXa+1Bpg2BZI2+Somz17ZFrjLHua0hp
7AdiwxwGkarvsjD2HIJx2jzg5YoMgoLfs6cz1NpecFeU88r2oW+pjD/Of30bIVIA
BI8M1fjE3iZjfAlVCxZribr9QgNZO4jYWUIs/j5sWuMNGH4KCfCfckygJjr/8go2
V8BqUTK+K47VG1J9ditJQLJm1+xE+9VE5NAwvGbfkqjbTOBPJhn+6YwTPYxThJqm
QyKK2Smj3Y/UVB88G2wbkxy6MctIQVQHbr0M4KLDVus=
`protect END_PROTECTED
