`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulXJOmG8SFdrsSBzfuAeuare0kWlqeptLS02lm04yQKGdGx7wM6GXp1m32Poig7A
BD/JWsLFeMc1wVcJ/YZ0z+AXfYzDjmMoPIVf6sEltkBi1p42X2rNx+Y51oOhhI1F
eVMntKz9eEqFxgGJmjNrMuAh2BPyyR22CwzV65Nq5zNCjUoV9mbKhDNHVHok3mO9
HYAZfAtRsEoFFSZPQ/6GwiC6PcWIssH8lBpXupq96xiOG2YcUi7K4IW8O/ROdcem
FOt048SAQOytKvJroxckmTL69y8i3uJyHYwLQBPrHTUu1QsocSYhREOKStq5ASq3
ELU7rb3yDKLVlLwu3Bncx4Tb/h9uzRzQ3k4Nl5GHzJgD3euJuH7ayqzjn0scK9cJ
QXCIiJmGJ1yA7EMSRKNQGBrsrDb7DGe8kz1AEgLsWK8Kc0DtZNwCFd0qtrqwZvl9
N6kb+XI7Yh4SNJHHXyrnD9tkczcCfTrxEFp3G5iTlHHgH6q+XpE9Wis/R3FXGTMC
evnIXBm6GR6IkKExwfZ6xNVbtiwuZy4bGvPa/Ao2j1lqTJK6K92xgmA0X8lwB3CE
OwOQW6Dajmfpz60jjhzx9OsHy/2jAy5biziaLkX93YZxsT99/1wwLDu4YafgZWDR
x1FVcDNm8mcj/IvlmnmwtwU/Rv4D2DiR8olHci6j/eteRor4C6zamz4uvlIiQcQP
Zk/uWjq9vkTXMS90Gz/c5lnq/DRgZ8CzTn7zREqEVeQhhND1dIgDikJ26of9XBng
7T8HvyJkEnhnM641Vuzj0lIUt+mSnRdPsMIdrB5DXqOXSb/F8Rx41TEAF6mKwYcg
NHHA2xfMYp6YYDLEWJgI4enI7VLYWt7pTKO9ptM6/3y6xq47EGEnDiem5ctVArQC
g5cOcUgHJI69MVhoKSQ9t1t98kxDPD6VnQtr3IpHPUoQ3ke4Qo2WSa1GwBkxSdMi
MTKYPyDzfowDKKW/8gRSTqTlnA5q8ZbXvRWL4nFxZ3pcljv8gmqtnrZ+ayTv1rCC
TTl+Nw3E2aUVknqhs4FTB6gal/cLF8o3IRbSL8qby7LwjKXw09lrmpNArrhFd0hC
+4Uq0nwFX8rr4NtVsBBYvBfpYdoaSlo0uigolIzczMeZgxYl7w4k+Fqb6+BstZ7I
Fs2DHkSX7qwmr8YVAM6/NK7+3T1byZDRryQvm6dNy624oWkFJjm+9RcZOS1Ak316
z0/T8QqIPSGXuLEmWh3e05wKYi96azYUepCCLNNlLwiHlES8zf+EI0H0FvEZaxy8
di8DJNVhLiNC1WsdFqHMT9feCFpBkEQECjXn9eZtp6UhtECo8LRDvQ1GXrxKeOmb
BQXdQKDMpIl9g893HFzEh4xc89JRdjq4QxXhApwGJK49/EVBMeERpWoFUTvWRb+4
QxbNyPduIjjpWlFuKrKYk54LhmA57/hxv3SF47QURwWcAoRE1aVCBwrxZaG9mIOu
O6Mobo4WZtxNW3W7boRetdOWIA/bQT8bfSg6T+DzZsH5IustkcYqg9EZfuGhlSMh
pAG4vsyFnGv2Dgp8QY1PaOBSOpVrtSv4JlcIxfV82pbIh+ZxQq0o3a5P4Ajij4ie
9CluTymeZOsEx02EdJCmiRyjQ7B73iNlrdUYAwGGCsw4t/z0TF+nQh6/zGdrZiiG
V3BXgCk4uADzjI+b941iJg/zjP8zaezANviJGSIIb/xGe04WxrBjbPbOHG9VUFKj
x5WwUM7durfFxtK103sFxeR4y2p/NS69va7baROmTIXAZLn0h7fvudDpx1t6Vsrs
Fi2QzlsH8Wg1gSwYZEujNdE/FILbIt3C9hmxQwmI0/CiRIlro8+ylLiAuJRzu7x1
wnHVr5VRrGTzwN3H3A/pn+2yBYVqp6a8JwufnG4BZIyS6tO4WymIU5g1R30zEoRU
+HZNrl3nO5sQUl8ZiJfotBDsHjJ4e91M9a6GfJTL88hSMjIx3bIUL54mgiyoqRsC
X8QN0pO8RSwdIs9AWKXEtgnrAM1oxokEfxY6w89qOgrr86oWRFBy7NZ7sgDohrQ1
/uo53HOCGj+XEEewhnhMH9tRZThFH3BrAVCmrV2l0dEyTl+gmosvbNL8wT5cTaIV
GS8bHfuURHKRitQ6JjOn3nOHKi28laN99dymMKVfEUoTc4gOl+10QRfUKzoblSl/
R1yh+qZmLXUVhvaeo67YEwrpZUEWWemf1T3Nbu82S/e+RmLPB2VKjMlk8SESgb3b
Z6q+5+/J6bkTfu3q6rLr6IollKO46p0FEMaoghZzIrVHD2vMozAflHPfRylKIAfL
qlv7by//4x/x+pRy9C4FALDDf30tYq/mGV8DXSUEmi8=
`protect END_PROTECTED
