`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NdXb/cZ8GptSXnAlVs7dzgb9VsW3X8dF9sDZL4JC8TNMyy3x8ujvHX+5fLjh/Bue
yTyZ1xu2zcAcbxYm7lCMwz+UZeBLo25xpHTzWaHlJcGNwlzK/TIY3X+1ghpTxCCK
W3OImEf9Bt3eTHrI5gS/RKHfgLBwJudHaFlSHxyRNvfR5/JL89P3/6OilhEjH2xW
5FrMpc1T0/8exfsZxRurmf9Nfb+/ZTgBdwMkVcR46ly4+GxBCzwJJkr1dgKbzB4S
u8q+/9n/QMWORMt5TdOHL042Lz8w+0yUh6yKWO4t64oicLstHkzL0l6Cz+1CHdKF
L6Rkp2JLKrkr+QWMa7G8voc0BfWJt8aQqqmMtkiMcLeDfmSN2W9R8SGMi8Hyxbn9
NLcR4mn3iKB2ApgCzvf1+O5XoLTn6tnGVoYh/I/2bHbLxik3kf0zdIJ4fc6du3Le
aFZCdrQbNn/oSW5G4TYplA7PoaFFgP7NPDCfnQ7IZvewiBPoHQDd/b60CdyrmMjT
xmioAENUkOQxEuCfWfWST3bOFWT0Rp9Dt54BzYsTFO51nQ+ZtdZmbIuZFn69F/E7
y9rLf70c60j/z1YAy5bgJvqWp55YflAX9oyJsDeTVsvUpbIbKpwHK/06/a3XhJlI
SVrggw4PicYM5/grnsRq2mXZi4IkWNjv54SxR8/9q0djAlnXtWgkjooKULABOw7/
Kk7nkKcRX5sa2qOztMbUWxglLmzC7Ew8srJI+f74UwHbJe3LlfLAnZOgeDDccaYc
BZz7a3LUK48IiB0+it2+8f1N5cDpHDtpS68FoK7S1mm/0RFJlBfrcCdW/CLAZJ05
0+mcuyei/sfn7J29Rwes1PdfkC3LFcPBCRFN9ymtpWbX2rqSASzhebugv/5YZVN6
Lex7DWvcu3O93ByqVkOOlEdXjJy3LVDR4ZuuOPHhMzPUEehqDfYY5PJBuadVd2Wt
Nqah98kRcAzsxyIpriQ5sFa3f7HKBCiUE0vw39ZyzMGNa4H6UHftwzhOtWkfrPrt
vejLtBR/HoYbEochdo6mB/BsWVqhaWK8wg7YO9GZepVRpUNpHPwT3QllE7YYs732
0p30H9zyIjl4xwEk1meJwFjwFz4LM8HbGR4dy6Y2IXEk3CDS4++Xz8jR1rv42OKu
rI5yBrfZLa8u/mKkEfePmK4Q45GNOM+bqF3dBI/JA6vGKe6gX4T4KaT4/8gun8Xc
Y5I/wi3ApPB+6vg+Vic1BJHM0DCrHpJEJr5vwQZlGfBBXUCR5Zcrjpy5/AMvjyWj
mepsCmAg34g9YVxN/8WEfmee+fluGKdAkkglxU6oM7o01vEa1cRdg4TF35ECxsYM
FzkjqPup3xXsXAPOa5iVmtslKbZOUeJHbYNCjJRC9pMER+GDy2BZuPz3qhP7QKNE
BEk8AI3V+jlftW8OYD9VO+SuNH376zztg1aFOlVF9ZYmHxHaCGE/oK/ALuznDKjA
qODG//r9RvamcYBbC/1UjsBYSrVO1KnFUF4AYQRUdaocff0sCA9Syzzk5As0Gkn8
Vsva1g0FhUBRTuQUlRvv17nZ2iv1YA3SECyl6pQgxRQkmdtao1ObVOCCu62o/lro
ibW/8j0BkA+coU1pI+H8ky7FDHr1+4MO+5Vys2QHZWz9XtsmAGXFs9Y1gaGRH9V5
cAQzTTtSyzWqg513so+VmhRutmAh1WHOXOQzNL6WWCAF86qAnwoRa+jS9pwTHbKF
f8Q0LlQF8KEkexjSMiS73VZqbXgvj1zOruDKtb4rAsBkke2NSSUS/vOLK26Ggoj0
gBC+kTVNpBlxLd79jkCwnbYEKJ2HW3D2uJ5MTRa1kWqd9jKbG0lN9cOlowMYaeDf
5DGDmbMR7o5q5PdeA9j5yCSNoAK7F0K41qqGXss7gAvcsOzNQ+KQkEuhhyGS9o3Z
g2IIB90m9nzZ+CZpTXCRzjVK6d4L4lbIqU/N/aMGG3+Px7U54YO65uOJm2OxYxUE
elahIS28iIQts2q0wdOOk2VgJcOI80zitbvIABsEBlnRgolQT0eVO2V9yRTSMh0y
Yi7iKan6np9/baNN5NV9qhV1qCmJibyVb84Zv7v8gxpNCuilOT53nDF0QPTGc0Jf
O55rnbY4o5jSyYI0bsSHFEoxMblpDW9R9SiYBsLg7pdMmbnGY2ys0No4wXDGRo2H
xbhiM57MC31A1WnOcq2LIQiv+vL6UvhsXqvDae9O7xj9xbiFsfimU5PetK82P1qg
cIfVgc+KE24SatRDszXoPdo4dEHhrx4zD1MdyKps/ya6eIs+yLszws1P7dfEQs/L
PbmFct2b1pWNWtWD+mbUhYgRN5gtPiW7g71tBdWGouk7fGH+72O2+TLyTuIrAn6c
2l1hWTUtAfes8o5AUc0V05rsZbPUAKnYaj/M4SylqreShDfRlQkZna0ilxFzJulp
BF7itWZRwDBkYYQWPe31N0LB01zaOQhgUXLh6jRy3FQPe3DEwJRNriigNzvzhEn5
Y9paaO/A8mn89ju9NUb8P1rj5+EXzUSSvGw5TGBW1MGG4svmccLRMG71nge6l93i
t9gjn4/vwwufaBcHUjGT+kTV4x3x+t0mPgbVDZ/hRFPrXJDDBZdcmuSHQo0cZ1Ds
bx4T/6MMMIUFLKFameWo3YAu+ntxrMmXrGZkaA1yv09GElk+dFxhwgUmMglVMS8/
`protect END_PROTECTED
