`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Shd6Z1ETeIDva9l6oCJFNXlAYmtSoWgaYNNbnk3QHU7nwZpOx11YDZQvBM6TB4Fc
r3kNc6yPe1kKAcqxy3N9V7q86x+16rwW1NAj1/fw4DCX4wfQ3qClhEK2s5dUagJ9
qaHjRipyYSy1J0RuR3g9weJU1cRbEEQOX8AoBpY3vGo+e1oPenfCkDfEtfU9MLAG
mdkk5Lpw+VqWMWCvQLqCsaHogSQ7BT11gY07BdJOmRztghFeUqkNUPy9fEBL5KqJ
KffCFo4w4qBZRPFhY1bMcqsmhXOiTTd4zBBbWXKUu4beM8CLbrPlIqWEBWa72aLa
fXmp7nGoB4P9e1wqQcaFWQ9rmb/x4A7XAgfetMt/bj75mvPQvderNfXOafgyuRkN
8+u/IJQmrQleEwVxS2YrYw==
`protect END_PROTECTED
