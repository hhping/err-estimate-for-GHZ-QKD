`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXISpuCp2FR7bzRLbhJCo6R3R6D2N3a4flmJmoTf2tl3ya7tYgGHbenJrFk7BKr7
dIyTeeF1DtJuGc3F5iBdnCPN0RnQqoWZY16TLDr3id2ztHFEFGEJ1Hwz2Pz+KAwG
1aUHni6mH6fdErMFao+BD6xrLKWxajlq0R5AZ4l4UdYE31JljR6UaZLkR4H0qamk
G57znqg6klV10QLfDDUJtbHeie4eY9VVwyAsEXeHRyOpfM2M0Xb3kK3qycoK3BxO
EVetaKj4/TJgQdX5VDw0dOEx4txpM8Xh5biGRikSxoq83dcmCmvHVRMgNRwjpq2I
OCxevDI/NHR6qTYLNNosUVVmdQpYFXUZl0glfT+34nhM1hb9MLB2dnobir1kjGOJ
gR6z/Ql8pCBDYopbDPGD0NWdkcchAW4HdQ8j/Cp8KQL2bTrVBTSpfWdBN3wMUiiK
cRjgDqb2TG1ASFbhpgfQDB9NJHmggIAH4r1D24GUJK6S76hf3W4HwA83hvuzKFFG
O06iAomKGOxCMNegwxW3Uocsn/D38TwOMFKE21DDiEai/vCG3JDaB9yJrqmjCbKF
VC+p7/b4FI6MT9jYW8yGjAq/PjX4fjRWAlf9QIhGlhcgFMWhWtB23w9TtXT4Fndk
LfYV+tLSxyK2OoslKXJIl9w+pxWmLGcUr4twEXjLH0Sst6brwC1wZGbbR3GBUzKu
fkLTKRL3x6DWAkfp0JeW5MhRiFW8Ny8AWgySPbONukMB4xJAGEJ05NJfY3TU3Gw9
TcNNQzmSmZqw0nG9GpI47uhUv8qCW1d40ACAztoll27QXCzRgQ8WIyP5HmZR1L4Y
0/VPtJP7KlKz3RJSGtOsqibVtl50vVW6KfRf/Z1kbpenfgpTWNtnagx3fYoKku0+
YJ2gZtKBdvNmAqS84djRERjX6xZ5vh/mjK6D4hN/TjY=
`protect END_PROTECTED
