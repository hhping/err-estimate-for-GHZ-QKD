`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wpLcLXX2FQP6Vky5yBiGEo/Ybi1uoehomSUuozMnjdJfOM7PZn1CgRPQzAESqNPL
pUNQy9XyHWmDAm2XhawGH9+o2qRovPzz+rCN3azyjTN2E7k4tOOQeagTHc/4Annr
FidfpfXsUnogL3egwR4dcOqDXO4Hx0L1Id88QlyH+MXxcSnp/2pmsZ5J/lQNSED0
9KqeOL15vqc0UWpIy5q3HRUDOOOGHhOk7O7Xk4Yton4si3kh5CY707ncZ9JKwdOq
+vUQnBAC2roaYOcibglMum+/aXb6KXj1HkORqOi6W8EiCJVrttHNIMALIhHiqCzh
ozIPPlTg0oqvJoRxHgOyJf9PtbPEwiN/1aoqrFO1f15nBzpFPJsKTD/WH/w8Eybd
5Z6KJxIWSCrMBnzfaA9R6idmQ9/wTP9ESI5x/buUDIsMDJqkcMdadhhy2Gf2LYtg
Et4jk2wyX9R2AiGTD3BI1WiEUpp5C9Qn1ubOVFWhfqUU6r9bUtq4SLM2goH7r7Gx
ssgRb45bgAkZvLgQfKLNQQKz8cWEqz277BGgfcCc3vesrghXl9a9CMrfFEu3ioaN
SEw8sfYJoaJKSulRABCrI0g2GpZoEjvfu1ovbMv2iLTqRrtypTibLIDnMx0RV1Nr
pHeHIqTIcT2mUtKl7tuqdBrPlejNYrHINhCmwuM1X8VPw5x6+AFqk8gDoGDpcIqy
vOxXkETZTV7EJc0lfbyXLbuT62qF9EdT92vf89wm6HRH+RYZNoKghZiY9kTeg0K9
2kKjsDVleG1XLVpNr5vuYKGUAq+CKtIdkzMO/IKQ1OCOkc1QVBP0LEXhijujjJrg
gHM3I4k9g3X4CHVuIsxsy9RHRVpeH9avWJHwOW2dcwEDyQjlRC8RLqgprTYny+kz
T4QoNQP8MhrOjR1WCncSVvsr5yerdV4I6KKLxlFqqURwqFNw8iQjRMbwkT+mEMMC
MN7HaVw+wqp2y/RIeZhJQ3F2n0t9Z73+CZfjTBcvq6rRDXvp1xrCDL1KrvZh9Hgu
q2ZgiFYv4M8uuNgsCa8Nexa7REBQij26zDmKuXDYg8/7kztVvwBhj2E6BNG7LYW1
UXLfM4tw3spBeOdYmtVpBCP8kRjX0HjdJaDlnhbVxQPb45y1vqVlncI9gy36g+km
my150L220ScYbyJF6ObWZmyNMd/jrqW6TNDUCHD2k/wh31eCon/fn9Vh5QJZhlf9
zBHWSnjlt3bghYFJjEucsg40t0ehTMlDs1REMHkIYWPB/YvzsMO3aC6rKIQOF+ny
RA0ZakcP+7o9Nj+uZ7MXiA==
`protect END_PROTECTED
