`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ScPAY12gK8etz37Zlr14G6v9NM+MVK1y51+WQPmOxTFhBn8aZknHCZ3AmQsQgRy
gxdK6nJqa5LWNVd3/PQTzZL8fFGINq0l/BRgSTRQ4JN/TaW5MbTtvq+NgxKQdgHl
7yi7r/5j+m5gYngwVTvZjuzWJeQKkw6eSt7SwmnB6R3KnOswTzAdNwW+MA0ko+bQ
oV4YqBmleDdKcXgAoQdBthdrf7PRYUmafrjUq11vhKhEBrIEt9Lb/uV7Q4NSKH1+
LudnbP1luyI9iSYyG3FGM5GiOCnItr+toluwO8ZiGQxXE68HmpPdKkzRfguyLsaF
KMJh19yZ55fhKkRJT+Rip3m/4UPkkeUTmt+ltdjCRGhurjz9PIm/ShYsQWue51tE
QVYBbPXXjbfIFfBHdML+QmdDJDwLr4tOpWDzr7ZSzs5F6ZIOcNamtAqCzw1D4CYV
HKWki6LBOU1ZCf+6lQLo3Uxg1BFs4acrTJSF2E6cXl/PSf5HiBQvy8nK4mMhDrvT
JPkfDZsiyDJ/pjux41/a/PJHcac3rC+IhbKQ7TkbThKrbnJdcLK67KfaBCEnBed7
c5ImRIl/EDPvEh6rVcqJx1p/yfZWRR+V4yuXqkO64z/3Jpavis30lFX5oXaW399p
P7zNu5aICukBnodSFN7453Bd/wG4I8SZ6TKrIVsi/uDmYV8OsZgpnU1vbEgOAwdE
ST1zC7odd9fts6lAt2vEQ0/YqE7eDd2k1E87Gwjan8Yx9Oc80wq+ctztkWv5ep15
aqZUVSwOSRB0oM8A+mJ7yAMlydDfPndPQvdDU1NTtWuTe2FZ9yWnABVX+s+P1FdK
+uLeCV9lStXKHEowhy3B60UG4DgbCRgo5tvweATRuU2pVVnV/EEBFhl/cx/qgKa6
66YsDC+DS7rvPljen+fJAH8HDV/G18ACWuOTsNLmkdboFsTEBzUHLXDKzeKEmb9U
7wTi42eDUVkms6L46Ckq5NASKQBpx249qwKhKrE7HZ2TyjVOuElIxDmyvcW1KwiE
WK+YpE3Q75z7ppTJr1gdPogqr11cYrTxjXIxiUAbKIzbncHZNR7vo0tWe/plnq4E
g5048tAgOWKseYcZId4sTYlA73KqHkC8eh5dnB8DC8jlbQL2pPhvB5eiN/4NcpRa
jxDPSCyBS7aVJAMzmFRLwf9cFVR26ldUwUTzsCOLDrjaEklDxqgfjzFM6T5r+2YL
Pnh/Ugv1v5CcG2jdNa8Nl8DbymWWQWr+T5SixeiCuCaiJLEGeU78iQNhMs+yF7xM
AXZcZWpBn5CC6HUD93lLjLv32vMTYFq1AeFfn1/4qmNpKUGVR8E2CFynIiH1OMKd
NZWBOHoWMPoVPUl9ekyPdHnWTtBdU6E3G+80C6xsnZlgz+pqDcGsiuGFHAEg0oNh
wCVJzVcqqxJqclDioace5Ha/2uviA7oARj9CTFpCo6yDvmTvrMVzEldY7zXRb1cs
R9rxp9Q606VHPDnj1MLj6ZGcJcEOPD61yz5i3WIRWGPvUVMHwRq8KdV1LfilaRqR
h2jfMAUfNq3deDlFYKjUrh1oElAyxDXMWI+YJCWL9qudTzteoLNqCqwwkILEPaTH
3HnufGinXQ8grWbRG86bEXbHppwSqJpfs43d5n4eXvkwdFP42HfELHydsOXL5++u
JCMhWtFiUq1OA34y6baL733XP9K28/bIrwekMFaud5imlsNqMbsZVlN+4fgEg/vN
UwZsEq3RLs3g5yghWHAiV4/OerSoilqYGmLh56p9z07Wfi4A0osSTnTwakIezUc5
wXIHnJEM5KlF3SJRtJtoNlGw11ebMDcLz5h3suVdxJaVI79oTUC9iYI/FN7MyfRf
g2WLuiOO6MbQVvSsjtoybhUazuXUITEDTCLgG9n3xgIU4I+vC1X6OzKO/xWfPmUA
oyiIeSRoaUajzNpNtBXFRw971NWHBnz82Z8U50+En1K6VSeGeyrVd/7r+cXEQrZr
9avUfRCYEmGhkIhISmpjFE03+OpWLoslkfWlAjHM+DtmB7oIbBmszDeRMe2d1ZTY
M+HGepYV0J3sGS9w9OzEhYqfdUaFkOV4E0gCgaivNDN+e+mt3+u9yT3lL6R3tmrZ
X6rxEj32gS/CsLc5UsfnUTe0Rbmce5c+EvtnsxRwRzqYSDumLSQcHSVdxbTDOiXR
yC10uu3a0R7NG2wVtvq/p5JJL/SsQW4WpIcqAOzot8IGMH7j7hV7YScU0+n02Qbg
2p/bKz6JvggYPrc+sHK0gMGezH9WcVtbHph78dObnCSx894Tj1qPq5Mn6r3GQHtx
hUxjsMGpudJhQnSSUBkMOq4EjzYhukmGvPc5prTt1xOA9BAd6aZyx5n3OkbtYKbp
eyhMyIS+wYZnfg0rsbvx2vT6i8enrggvRdQBBcC8wsTzxaHxeCPZKEmhzPxEhZlq
oOOGN/h/fZTw+5jrjcdZoiiF4sM5eOLx73pqC0Ho0pDXKla8jg6VIhQWh5xF/UDP
xtHmKjrhjtF+kslfI3nMXt8rCitVcfdglGBzgCOPsuAQ9q+nL1fL/cd875t87WGa
DlFRex4CiRss0BfRyO/oBYnM6y2z7emjKg+Tm9txeCavXS5HXQs5BSCVWsE9P57A
eH+vsWVjomrt54R0pUJnVaCphRNSf/k1GRZXm3qdf9zcUncJLtopcz6jkHthO+Ot
bismzjqIK0Pu12tQXX+wlt3t6KtVO1Ntyg//k/MS3Gkaz3DoGJ1CF4DS6zigdj3t
AnvnQsXFYe5L9ZGaz+OKcRKnyoDgkdWuIFBw6SEbhgNTxldnoVar7yljes+uD9qQ
nClm0RZMAxpcs+351/HGXrgUblCQDWVw2CXCZJL35SpwelxHjCkdnhitSqcqG4dj
PNuDDfgp5HOe/8zKGhbY2LuUlK1RICaFymRmnb3lvbRyDSh15a6kL+znplZA0StY
JVU73eJfU6YZ2IzD9rWXleWadyy14iHhI7bzaSCnxnt31Ts/aaq0ktIDEL7umQV9
cf1o6T/tN3OfS/aTpFaC6VWveD5EjqJdbSdqRm2KiehLTyiV0i8Oshqa9FNWVoaH
AO6iiQ6V7thwtiea0kBgTX0xigM6SHNfzEOnu+hbk1nukP/k2hDO9ZYatIYRy/67
HqgEY9lnqHy5EjcEQS/JUNyUrmZvOomYJN+w9t36Bs8XY/aRCc6v995t6XMW3zJd
bRbOkY3Dr3q/aFXvC3QCoMJ5lvRSC61Sl3pnzel7MqiDP7TfYkb3q0JmyMuH951v
8ziVIs4zoSaGIkqdTPjHfSknSn4ezQ0fnx7GTF5jRIwADWFNXoXrjf8DJIklfws/
pfsZ5GLNq0ZPvY8JpRq3NWL6NBCxaWxSmPWIRTuGKcWPtqOrhC2MdX994muRDSk1
ndOOaNELj/iB+PHkqaf6+e1/OC5dAwQULLO7PReSkCuueBe0Ujaz7iUgyfeXvaHm
d/xJQfWrVs5GGjayihthn5Xkaw+bkhiRiqoUmZV5WR5StN/9A8fOX9uDk5v68Jtz
BZGpMpD52MMRrps6HWknlxk4IdLAlrm4HsN6JjyCVXMjfBRbSV5QWSI3XzIVkRoE
DOq31cKThpoS6bUQCwWk0kvIA7tX/yJQ/G6QN65vGJBS8fzV2ieEkJqjMqG0VhuJ
gyeiDBT1Mb8Sjzye+jkBeMh7JFXg1z3tyBHoxORVGj1enbCC6YpWfDsrYO1GAjm9
02etcB522dCwE94qwxsP/jLbwO7pWX/Kaaxb3xqlF2UKrHHIwqzwjUvNYbW+H6uj
8bvIdr3JKXptGpajVIIEKahUQVzL5vd3+BwaohOcq+QfGr5qHJPki1NV134Qy9Qh
T0U+XVkueRkyaqaP2B3/NGLTrlhqAQioaTAe+ebRlR32+uCcXMpeAeaoiOyRRUvS
OS4N2wvw2AP59+U/YiPsiBYuWA4v6t1apBNFVnsKNgiR+EtJ1KnjJ9P8E5YL1nwp
6EfkhT5TwTN5kPeh9vTyKlMVIfGv3/ituJkpBfsc/mL4fvH1AFHlR3re4FtjCGM2
v46zqtGzkXrbDKzSsWJ03danODTixiz+igtBOWQnaTf3vq70v/n1aEqcoIHAjcKq
WFF2BBXKOtqbuVy2eRjaKUMpWXmfGeo0ziMrkTheOntXvZ3M9ttRdNIpZKQkAnsc
U0UGOk93jmdxOVy8pWSvqtdRQmN0hneIKcmBAqjbN/fC4LBHWor7+hgqZOL2/JDU
/khIj26geDkLMP5gU6n4eO2cQ1zPzddUNQ2ndpx6kFI6Nns3ZpQMDN11WnB4uMYa
r9zA/XWQa0u4x+MlVn+BqtqVhExBQ2ngQz7kV19DlA84O7bDEJrMzU7V7adGwJtc
3xPPyqtpz8JT3XwAPbLETd7OKpDf3gvxln8twwA4Uu+4wUgv7DY/7Bw8dFydYz8M
yDGQJaHO9EocsZcueGfoRQOUDVntz27TTQ3V2noPPI2xbv9fl0G0tAXPMuwuSpzw
1r/ql5VIUK4Z1y0oaYeLsSIUP8TFHcVAXjWDfHrcN19x4d0pfPYpf+mYxDe7xnHG
+1X572zXoSLIjmRMwS+hRDkQu/Vedweb29fU0/BTG4mpAvpkjw6YnwF4LphVvVGt
beiWFnOBq2GTAByZGnqfjhJuUbZcGkZudekFNgF1TQkkVs4hwitPhSshiHbPLR32
NnUKT7ajbVT0vBOFi6f0X2KQcYRWiO1yeOi3bx7MqZzXso/zHRRSxJDKQYI/iCYs
pDnJubHrvuHMj+As8cUQlUBZtO5wEihYqgR90ReULTifjwIJ4Ldc9tqdFM4QLIHQ
2tQIcRnd8XwwsKNXdggUkkiEdrj0HLpEE18+7octCIL/Fo5nWx3Wqhm9L56Llrgq
Sr6I2Af5iCIa1Rw9YQv+LKhGjuuJLppPWGN4o/F6vTUGbOzH/fhGtPPG7rnOggsz
aIizKsiOt/cn18oj1mXY520uHg5CTX1DsH1C5eNz9n0xaSkSM9UFwIyT6DA91wIi
gYBqx7DJ/mJyXa0JQztEgM2/A2NB6ap+Iygz4DExpJLqZ+slBOrZi7vjOKZPKHiO
Fgsw+bqZaWuSrdjM3OgHio9/nYiuM8eAU7FBkLrE1QTaT+Y59icZTt0nX9SO+W0H
l/9+ab1lavbdrolC7WU+YxVvhsU3cH/c8z/j0IqCuieTt0LZUMMrqP2ltcIHFyDt
YhCVwxyO/YqXzRCQhu1ThfBovst/1k+DlaVczuitSjzuRV0SZbmmrPCsP4nQZq/o
rS0Qgh0GFEAWIUBYPJZWyv2/otDuoNf/eAEZM11Qf/t8Cqm0lSgYEO6V2fm34L36
F3RZCQ10PajAt6MTnDEI6KGO3EblR06fsaHwUIQo/cvqhWGDZ4pybNX0NdVltO2o
21g8piAvm1G3CBZ+SCoHFoKdToYrmtHgGqQaBtzXJns32E/3CO8Eth/nkxE8TU9p
A6CaDhkL40Ii1uLKFnybz/sQ+6jsiBugOfu4ZA0qC7uklaH6Y7Tf1VRHCE44sgkh
78yzp8l6UMGqrY44jsAJ77bgdhPbcroRJ3/hyPTsgxWIviFrM84t9XDPW320b3mG
mDSuzYvVSg22zb5D4KN2enAee1EgeoNfoffgKHNGhpBOHjPkoIW954GnT6KpDzVH
S/5cf94S3F6sCOor0I/KA0KsJddf/ZpIuFFwyfC6R8Nw3351y0eCdzvdoAYEqOvw
74vhycV32vDv6BgeOwWhcDM/VzNg8z4oHRgfqLhbyliSZQjo9AZGXFhlguH6F9Fw
vPVmT3axTgMoZjtR0dTpBv1sTf2tGXcA2nj1qx0mqzzLpzVeJMk/08lbK1/i1SeS
8t+5uIwFuXGe9R5WTvoxJJxQpwckOseQFqXMUIDtYWAjImT7UH0W6ByisaTyhLMl
8vfYkEgAQprHc+ZGGgyt/1dzVDYIMcDCWtRwm3kLQXyXwC2aLjmsv+HsfeyCf5ke
+Hu3Itxwq3qXfcg1OUSX6i3ziNZ7XeQtCwBkoma/ihM11NFZiqxX1aHy40hE0ynv
svRAfOijsPlXcASRtdAONnX75QWj5hsniEXPH+hDjdX3g45OeA6JeJcPCZDS0yTl
u1qmKzsQ7PnPyqgMOGwjOMsSISJiq4FUzWutbDXm+2GwogHjTKJDJzt5pdlRDl2S
IB7XZvbx7y0KkDP+p0qPPD7C/4DJum1DtHzMuH0y+OqReKLHbUrfbxEs0V267BJe
8/MtjXRf2svELP4DlJsWhCB3r/tzXCPOJylTgQpfIaZAO0h3eeznLTHzp8iHb/+9
PaESqpDBJvQK9eoU6zEGaDdr1REWL7zIH0htQyRlDodH3pm+zzFu5c4kbt8MJHZ3
8mvBVj+INUme+thVn6Dr9w4UmDJ0eDI/H56mD1W1Hpjzk967xSSn8Rwxfcr9gJOI
ubhmcTXLHgN3mZUxdep65qtEFkbYoX6xUCJkgFAkEWyCTYb/JcEhDf7o5tkYGib8
B9IQbJPWxj2ErMr0cAoJgYFuUz7zN9FRLFI6yFGft4BANoBF8cV+aN4xSdYD7n9m
nxNaRzgROIQsxOLFugkXevtb7VkOXkQR4TzKldZtE9NKbL59w1cw2jA4IKO92dfa
rMH1qgfCt9ETNmk5nW273+3gTfpeo044kXrTHsh5o8wGU7DpBODV1Vy8nSwnzjKL
RcuTrWzYyoG/N2BomShzlVtzorl5uTP/Me0RR8+s5R0s9sx+hhnDb2ZJo4A3nvWx
jE0RTyFv8sPdo79GrYuBicZ3AsXVy93Qogn3m6tggRMRRaB27Vw0h+ZRXg5gGlZL
m1f9OmpQLKxrDuz/3uJohA6PPJ64941Fp8Sohy+iQ7PRD7FgG+EYVbemntlnLnkW
vGiMAKBgwwowzfkpBPuM1dNvuATRWtY2C+P1QIny5nOSfZ1k9KyYi3NMbw6KXEeX
lw1llTwDLDw4eiJ8/jddOu/zwgbshXyxEoJjnOpZtMtzgrSOeY7R0KRzbgCHiHI+
ktYdkwbCNuMtPlM9S41+85h+7NLMaZnRSqk7SkvNDDLpyT8Ed+of3qrlqo/b/5Ok
gD8rdpKtumghv0soBKnhb/WVKg9Ib2wiVRRV4RJh7SAZH6toXYixXvFKwUAdPYSE
APt6g4noRDRiicx1hq9P6rQ3Ty29Z4yrInQIKuUbhsIS3syfduRg5zeW2xMOf/oX
rYh9Tu/sl/7SRc+hGfXS8Z6WGOx7U7MnxFMXC5mSZR1ri8EnXiQ/HKPQtHkQLYRc
Fv6oeqzYO8SHjMBxpzlqu0CUVhFM6kXOA7WLDd4/pce+Qa/WpTEvOC69dVarVRnp
kr4cMNa3ld/OICgwHDXIzTLzqSho2LP5gem/ntpxhDKjK4V5gXjv6VXmJTQz/WWl
ygmvK6OFiyzD/Di3vtIT/PRv96AVkCHnbRWUb0Q+A/2JQimJ8Qgr8/5AVqRVCOfI
Y/zcm8QjJ/mpBrKHEGNjBPOvq9ILLp84wB2KhWTY1z0DUaMvT342f/qvWhCLfp0T
XCUVSZifh6grfAVtdhdCIx7VgVd8lPS9Lg9XK3+q83nx2HAJpXMZPKzYUvqezJjO
KgtmRnoALE33LWkC2TEi5QBynS8MYaSlWDRpyuxOQF11rR50eNo7qR/8AN5XVE/g
yjqKA7raygpE50rxBwxh9p/H4Qvs5evuqCJwFi4R4A0NBpNqAL7nweswVKxghG5/
k63EpJ4AiG/byf2wVmVfPbDp7W8sqXBZvnAn6H2QoKCi4GyNKPpNJMWdTAC+lSDl
H60YwCUh4Sy44FADGTYc1UKyLZyGHRtuhITLpo2iabDSsMoANsg5q643GhbZB5H/
WC48+pxlFvzjBlejxOa2ZcsyOJ6GPjVKMkz1EBwJKnyq/qjezOIZHX6Z3h/PGD/s
w11C0DlABulraDhRKByvuDEsgLSqJ1G9CtcGdUoQCdIGoWZyLkKrXdd/kML3K9dL
Z5j75XrRLv16tXCS9sL+xRHhxDowr5bN47A+DPcgKN5uH9TjI3xItPl5nvfKzA4c
GZNuA2rJFB/UG57cFO4nZGyp6xfEJyaeZ8icqgoy2U/hBlez4OjkmIRp9PTevbnG
/gqg5GGd0YbSXDmtGb58pEWsHZzzVnOsghSM94sgldeLEBy9K1IRWSFeAi2vdo0O
08vu5olYtRlmRKcL3On6xbmsAuH5Lkzv/0+XZy+DiAv2l/ntETWs8NZbcEhpHERL
8n7fdwDybaVIdWSM1wI2JiwnabcaTlH57pQGHf68wcPap9zgtckL/0iIm/U8umWq
mKjTjiHJo+0X0g8dzwsRVS62pJdQWO8bcTA6ppeU8UEm5Y6ZxXDOcHtskRJUakpU
soEp5bEAAGO9lG/E3bI0SzG7Sjx/pUMklujFl+aNa1F/QgAiADdELtrkdOaAC7UV
vpYkx9kXFsDxS7k5IP4q8JOI+D2oDTI4VzGdSoY6qp9X25QQ5/RItCLSxsvmKC3o
f0QurNvAq5Dt37eugI3MmqHITRr34Tzk75M177kuGcE4dtfo6YiucI50+B0l8kSU
nl4NboQZ6xtb4FFCvnja8evi1+QFhG0Y4Ij4XC0IqwG51AIMenRY6aiZ8mebOAHz
5xZEyPZHEEMt27sueDpULX0GLNm0+ftY63sAGnJTCe3BPniatq4B9+VxooVB5wOA
EpI/A5eeyY0C0UDXowS95zPxUvS7c1Sof2cMSvQBi//egQdXNgj0uXxyDimPQNs/
5QCMnYoBq18y5GZoj82u+pjZ9ul0LF6L+T+PcqogIogics5fDqoakBOf/030rtoj
jiy//rX7kMbkjuWD/joV/Of4Hq+eW/3qENqlxDyqcfDe+RKIOkm2LMZYezQxREF0
iyPb5/w4pAn1cO7bZxJh4a5ccXL+dX9/3ssY08rXX7Jnxn1QxexbyO2ont0YleOw
1SoS8n4WICH9PZ39N5eXWhNkKq/t86j7CEpT1J5N47tQCKZl74k3aGRQv7D913QB
sxjU7Yuy18a1YzN04ix1kbfrxrsUbisPcMhQHiAp2NIM/AXmP8IwryN61Mz3Ppfz
TfBSHy7ygBCQ5eLWh2ftq4fpmmlppqdAvRhqwRNIO3p55qPRTKIorpPMFEyWR5m+
ndJe0s2y+Shzxjd5FCaPDPSJrwr5cFKrQgExI8An0pu1Kyp0T82KN02sJiJ1KE6u
TA05dll8KyK6TZC5YnvTC5lEdH8DrcQ45ksXf29kzhoISj38EOVn17TETFtAMqgm
Yp6cUy2epVAINk6GGE26QTLMh2Yn1sXZ74IgYxZzUpuHCN0Mrp3xNgrhGcL8D9Oq
ChJtZ98DTD5QvIkFel5xSBEZrolX/1JsIdbHgDE0IOYBRidqroYgIjdborrtKVPa
c2aCBT5pelh604M9XdVcCuTI34jGOV2wGETg6sW8/kmJe8o0JUuw2ECCcLOOl4QM
wCH2n1V27FrFSZcfy/qveiJnmvqE4k94K2bEERcC7xf0pibMiIYgMj3E2YDFSaiq
cuyHWwkU38Ooj0MiNrUEi51vufDv/VamnjNlWBmgo/iOtJb5beBxbckJgynPsj46
SL/Ntr0m4jth2aLfTXIuu5y8e9fcLc2uFyxrw1imOvXe1qp/fTomKiY5lwbzDGcf
skBjwqFZS2jvODV99183WFl23ItK+bHyqBGqGvROiI7IiGHvnHaTj7EdC9u3hcNL
/GXd9t9jY94sWES07R+CNiw9PPW7vU2Vfn71fpe0CpNsbmIssWrXWpK4/Uv2Essb
nGa25ph0bXVHy1vsepHfbHgsHKxKF3fQwtYApVBE6476k6d/VqC7hmaL+B99sGts
iuoBuXzviHJaVmuTQ5seOvEMdch04gc/SJadQDxoTAzRcOoAjvcipuOwU5Jqut0P
hZfmNa+HmNGtO9qwe28XUDLZYEAF4mGX+BVJkzGW91SMPdrg5PavlmeZsjAmhLlt
11vQUfhkQAQJn2WrZdaJeMIvN1aWg0eKjXUhyzZatUbs0WEbcThfPta9kqjCF13L
W9VkT8kw8r7TuV30bq917pMWJy0gR3Wnq5ZWkPYoQbn7JVVjds+cxMFx9wjRZkqW
kOyEl6UkJgVpXDBGo+2kVw+PpdJeB8Y9qPQA7pNnMRtvYKb+/nHHcaHhwj9zmMX4
PUVQ7mzP87VGTcHRYET3jUk5ljogMdhXsPYYkhUuTt84IX0sMSFPpYbQZF4VTkrS
LmfWkeRdC5O4tBlkpYmKdCzJVq77MMCbFgWANOf5FK/iaQ5alsWS6L1jPRt6ECap
LFCx5vir1jdNDNPQulPNmx4WqlCysFqyGIA4zkdtS3IsPU+AYeHkngPWo9BFB/Nh
5QiIbThgKMHJWfMkwo2CGlHj7ywCUynl92kPvGbWSENtCiZoM2qZHuucUT3B09i+
xZmUd1LBFFaHefOmjlFgg1u65U4VB7B6y3D90bAHP6E6zVPOr1T2Y1fmOApOLryR
blOIOoYZu7BxGY062Zo/o4wvKa//UnB6F/APlBObwDb+DegtulvmQrsNcqPezC5Z
eZ/FmAdupFXMWPzjjXkx+Pk+W94Lrt/Jyx8P0VQZ6vVuaIsb08ktWl2P3E41kIHv
G6mhCQ5TEz3FVdC8XMMDkWiJLcpP2Lqv5rsUNJeF7+gGrER2/DKVtsR9jlkSZ7C5
Y3FO5JbW2ELJdDNJ7MYd7ylzJ6rvcvTf1rKN2TD2BAIC4TtH2EV4i/3CNYq+ckc1
IAoLBneTiZDVnkf/v9w2mTKXtg0VRUYYzCxD89JBmZMnvZcoRwT/6Ryd2ptOjXNT
X1XfvyapTTOtdmUJWt8IC4X3mwFsjELn0dPMdQ/AnaM6YAaunGlcMs5enCSkJMn2
FWHE0AFMixeYS2dEIQaZU5YrXj8TODlffUgdxc0k6zTwgtyBmYxAfAFMwp7BATBM
yOz1b2SyqWKoi0fJk5dfvc+7fttPAyDVP7/W3fHWW5zOO40rzIJC9Szleg86ju/x
ls64xFAWdfKOlEwCpDm+dif6AFQlhQUmV3NesbRkQPksT3hygXuXN7Vi+Y55FWy2
wRtcvPyMX8lePI0RHSVnJvQoO98ylhwjhIKjhRyOmG35fqASDg0Pshwl2FQ+uANl
kdrCFmLVDeKlI6f72w/NWokLVKRqL40G86kNKQsLKpxs1FnOE8qRqJsK8/If/3Zr
3qQLr2Oz0M+z8ng+W63cQD9MZIP0dh2HchgIiLERmpMTpEjNAgTRQcH1zu6mZTSZ
afxfIkbQmlFMvGnRyzi7+cRn2B7CNevW9nAZ1HN3yV4anGQ+tlCtYwY1FYasmMC6
m0KdDFJGpYgFEXvK+4s/cy6Ck5KWm5XroLYNagJq5Mu+F4ZVrLZ1+HLbZuiCGCfd
KlOoc+wgjTjtSnEwLhQ5CrHv+mwweYXm6nYcRdJRpqsj2OJAuR6Zv08ySqGbdKXj
/QC43W136hrzshyWtD4lwtofe2dNcaHlNg1/aeJcRIdNtK9lYgLmXB9lzhqQw2U6
xdsyGIbLPraxcympu6sGX5UZX86a63P0U/ArPPfqF6Xn/OyUyO3UTmlDuh8CsS4T
32hWjI3Ar7sKzAAFkBhvW0LNEFFiZ5gwH3uYAPuw9i1yV8AR/92fsddo3pXwvaW6
xzqgVVtcuQSCXy0KigPP1LurioVWV+MNrcCuF/+vHpAQnEm6NtvHdcwGglmxhttw
0VFoaWJjQL+4FRAr8eYTBHH2c1m9Xq4hex3DTNs8zUIXap6pImdcUOhlHzgLXLP9
JwYMgSM9rayd7ns+ScbZ1B2NgB5Lcaz8aEMD193dNqpVyrtFn1blQL2E9Pcc4xY7
nnCLNB0IIFJEcITiOzTHYG+BosTKJipxfCmQb/4xRE7j8tCL+KRd0Eqndh5F4/ry
N5KGRbBTpePnl+fWHQ5/sS3c57O24QzxZHow3zjgKr7AjaUJiXW12ZKXNz95bbxR
Yfok2MKuRKqDjt1TI1iFcV3eG20LlZS34RJezsIe7uv+KtmHWNgxpzmUUQG0354B
A0FIM92aLE0lFAXxUyx4kxVQKd0xNRjXoJgeDhXhdcE71Chi39tL3v0jfLY3Sg15
Rbs3tws7sRlWC2aDjUfEauWAfKAOOisQSoVEyyI8Sntvw64QMTkLr95gAOnpMcFZ
HStfgT9oItkTy5IH2Qowu0qGBBDpAcRDOTnaSr3Tm+HcHy6bucQUHIg/WPrcNSoN
m2sYp05H1P/ZRLUnk20TRzAsSPwW7jAmI8Iirl0YEyJkxWzVKptfXiYCxrUE916/
bRSIjG98fEqI1cvTPN0acy9PzMZ+ZRY3KuATFpe84gqdjy28pKCc3qAcvGp2Jj8s
fYxA9BqpcCerhWL8atdYz4WZ9MAmKdNtQBPpLHlJTrYcgFmlae6L5y+E3wVI+Iee
CcmaVKy0Mm3NoG0042MHr5UJUZYCqmzldei0z6xgDYDnGQ2o23c4VcoiL3l6gOZn
9n950YC64PqUgMGUrTOd1euQtcZ6usXgkTgUrxuqzAgQKWJrvj7gURAwWwEgUk4g
onde81OPI1HmmqaktDHh4fPIBLX5/w+jUKJqwLIl6cjVGhLmPaBnuhk43X318umn
KLKo4qS1M7zig0pqNDMRfBJJjs07ih+nLzdLFBAZnruy6o7ctnZ6DjWT1/AqrgGL
uEal8GTWfRbPMCaG1e7b/w6Pywq7bB9Y90HENJ0UEyCdevuMEz7JEgA9HS35ImtO
3fPPgz2QcevjekyZbtDfRUjP9HonrSMsd0JC6DAYYqqk7VD27XEWnqYgCCik/RMy
jANstMP35B8lYk552S24vLRC7YliOYs14dfbcQUZ0yFtcugQvVmi9lxuFyWAESal
k/Q1CdxRCgAzln/zrMjv18LiO7KM56mrK3ydB+4ivjBvql5wrpdHixQIAw/jM0kx
WSNvsVq2jkKctZO7BdYeHDnKnI9nIwEGJc8vSA2W9UyMRDefLm6SYb3PqFkYngVa
FODiMfZWHktKxM4zYk/oY5EBFrYL/pOZA+NtZLeuX7MGPDHCwq20p1vbsZSMQ/Cx
PkxOTHrjmPfGpG18XWh7gH8jh4QvDfjXBprZ2veJBBnj9LGlS0YBlJX8OYkOZTvo
UyQb6HlM9eM/U3tK7C0zFycNa1RnLzOciCAJCZhYj7QT7sgQJHi1smiDdlk+RMgv
41WEKXjodKq/25qI9ivvGVZU15gtFTsDan3j7g5IEL5JVEZp4gsiUlRlzYoOzecw
OsdUh4P0RPooF4Mcf7wvo8ahee6ZWz25QzEzkohOnYKFGpM2YEiCoXL83EXSwN6r
H98k8J4WRGEiLKnP33OP6lYQ92jLAK1i8jcFu6DFkNK25VET4RuiN3lYk0YIJUJy
tB5vqscJvrHmPn2nIHh3jr47D39bkzwXZsUxvdDL5JBn+8I06NnJOgJwy3Q4Wmja
eILhswKxdcNISAroUT7PrSLLac9gTqjVboRcGgWnHweOSJCwlV3Dy7MkNZc7s2kS
kSKnZz5Yr4GYnP8E1lqm/sPcnPSNVjbcPaL+7IDlHmRCtVQeN8CafFk5txnwMzol
k53CyUljOGJ5zY42rwJwDSiBmQ91gqzgD21Xxt11TdDIFpH3DmrlngCqmyXTS79n
sNkbp2hYlMpPpQRk81WldWBsXnGGrbFe9kcBWS8H50Cx8V0GGYrGPS+OFFdaP19W
q6Z+XzWxaO52wTdtAwAZY6MDCXPHOWWistQhto9kqZDByBPGQS0+h6YuVot5tiAy
ME+DXCL3sKaQqg49sVotwlBSSPFzvqZGjSRauBicdABpkTCXTsS/1noZCDFstJFm
m803rvquxKSeZHyMOk4Z6tTDBbaufyKQMBNpr53En9AL1/h4ODUA9e4jsI1F6cpC
q/kIwCN04MAxEvmrOl467B+nhoC9+uLMsGwaVUA+MENgIJY/SZHi5CQD/lIecBLn
Gt9/iPrqr/dCyBKSethrUDxNzwQcIAE+dzzRnOULlgTNnphfnzaQgkAZamPPhK8l
1o83t0Fz7Wafqbn5bxqJdn4KGSvN3kK1vIDf5nt0aAMtwy686II7WL4EzpAu2tip
m0lfgNt+J+l6QHeUbI0x44VA78ics0oOxTgOzfkPeVcGhiAIoZDzUycYngvkuPUx
DgOaHgVtIrMjwFR9zgx2KtYI0ltsJ43PMgR6PKM5/gntHzUcJTeOLafXhlBZJQq6
1g3PStkS8hxnQT2kyxoZTJBj6fUNFnIAb382iAXD+UQYCPFk12Kw90qJs9aqnS/v
gzYcEQzkSWkR2Iq8NtItI/Yhlno0OTvCa9+gejQbnegZ63nCPebJaFxbSPjAlbpd
nBgDpLfSCM2XHjruVON6An4qWrxPYi3I5pXVeei7cb5w2soYy589zvDT4jsOB2W0
mINcapNuwu/JdvkR//Olv2zVlD2UWkY+NAIbrWa+m1IIIExcKYgIj9jo83oJRPJo
eE18VXkGks8hL5PjprhgDyuF5GPG3nZgIhRKK/iG4QbLXz1A1vnAPG+N8d9nnaVo
FNlQDgGTMxLOF3Pkt5RXbpIGUQOR6MJARdovz3evREeJi6eN8zpcY0WKAKOzrIUz
AKfLiuQ/sW+jph2vXmfW+d2zA5Q8Pgx7jyWgmq0JzLwPqOJjtwBJ9W5rz83JJzFy
ID+BzefivmVjgjSeTPF0uqiq0BiLQgNIHIFQtuYYd0otWPizuigYplVw3EjSuyRc
KT+xeC906c4rfmwQt+ehj4UBO+iSIpf+4rXZRaiZlBCKpFKtISDPlbOpRxqUIPFF
eGzdO3DSEahpQfOvJiO/mLPCi95FhPbser1jFo2Bdn82ZR42U8368BzhD37TcUc8
YB1IKi7obTkVm/cv2MxTkf1LF0LIHxjSyMTdMGsdS6fqYslcZDO2yPhBRzHc+CH6
+xZMvHA+uWca6/tk3+Vz3qwz6g+ScEtfQnRsyUtaEFyOZhPBXMovzpdDSdaJoR7w
riyMzt8XGclBewxOACJKdTnuLawxlgywQALN7e69LmmbJLJ7YGsICyt/IOTjMFyG
g+J3VGkXg0Hkabp+2KMkUXDbkAu7iF8zh8hTU5A1GdpQFayiBixOclXM2qjhmovS
znoPQG1HGMI+AvFNgN3j677ZVTxFOtFSYvCkwNBeM+hmYm3YiNRCxyWOBRuGULf2
iN21K3skKsrFaq1OARq+KcqBX3A24L8ZJLbI8SQAcAVGU0oC83SGm0IEZwb2fcEF
CyG4WM16v9rhegBhLX1dN/6r6Iwvdv8+af2uzuFC9rz9rPYVj+Uuzf6oPph1d7lE
DMeQBYUa+zUj6W3Pe4moPTMLaMFchs7ShXckls4XZGkwwt3wVREgxSYOE2qMQo/7
aSGkRZy+PPXou2Z+m8XQbv/koz1ESsDqiQkEYEuq+5/yUBvapDLexAIomzi+4TC8
x0VqCF0zPEfDncJ+vX9O29SZ8yhwjQ2hl4bgzywQDTJdzvT7jo6vlZIblqGdn8Dn
Fy1Q3xjWquwV1Zd43FYavZgWJAKiUSRP9gUx0kc03K40FeqMBTZy1KFRD6lSX4ol
hExCKyoPXGkXoC2rbkKH5+FPl3Px/JFYOxIwy9qiGWs5ulhIPDGu8P9ClIbalKoK
Lw9+m/9WHAC9N1qvGd6Bytoa1HsfOtRVObNSkbXbq6yhViKMQPFvXy53zWw+ULqe
JVtgbIp5Y270h8T+JUFz1wiV9KEfcc+X256T/4eVxshjXTNI9ZkM2zoUf2dM77QD
f3Og3MUXYPtjdePfOlpV5lE0w5ABEqXdUMu/ZfIDBiaFFSpezxCHC5un/fxPE4hk
9IFJXgzv77zn1ZuvSGz7Lr5Zrkjwid3wfb8fuAy+/wi7G0MibUIENk5HWk1KSNtX
elvwU4kPuFJr1QedFWELHsJaNpHiMAiXs/DO5XTRyda6nSw+9mtD26VqnhVpFlGw
UmHUkf06aquyCxOTLX1d1CMmjC9IQQrEFdFKuX3YOLH+Swz7OxT3+cH9SO9DoMXI
OeROXLi9Y70J8fc2ml1Hp3GuDNi/ptd8hUKrBgoin06YbvV97uC6hrC831hSLWgh
rN6FQxz2WOuCoI4tVn4xGxLewTA1ldG2A04oYrG9phcPR9vOAWDFo/vfbiGTwiKx
QZx3V2AeKJn9KZID8XMFt2fampnRhyFRYIFEblGdhqZIM256GbmPBeN7SYucwo1F
dTOq1+V2Ca4dNMpD/7gQZOvqzBTvbQsR/KEN3Fz3vzHJw1KW+p8J6Slks4K8Pv/y
6yzr28e80buFSyuQeF77lCoCLuPhOWh8PJJ0p+B+9sf3v50kdzjKmcmbzzjJAen9
9TOKloL/WDwC4RVrH4iYhZ5JpDOlR9mF5+cHq4cMXcUryIr2pBxQGnB6Wa4utHwK
Dy5x42GFirl9S66iaUihHXe1/rF5u1vvoJLys+2CLV+aThiDlM82urvV7ocSmRC3
ZP+it8FVcg2kDxRdQ7yDbta4ZTp7+6lbiGzgkEiAysDPoZT4StfzkJxeemVd6ztn
Jg78mPt74++x4/uKA9c61RK4LAcdT6jc/W3G0eKPPGAkmpoMoS4iKkd7uGS4Fj9X
VHHv071kFbpBfCpy2NTnilQmWomIStJeFgYtmury55CFpdqQWa+BEWqgc9Gg6T4x
bPuLA8hF+IEXyrrTsct0yu60gMdZdM2uuCwgpLIn7yKlRv4i4STLYpg4x7BoHXsB
hTJ0k7p1qnYwMMm2q4O6wOoi/3rLy47fgvU1SDlw2jDpFo14tTOtn2Qj4qCepo5h
bCcD06PPAMgzUPoM+CNVLoDtbhxrAY5vmtJuQb1CtYyYUrkJ9IKLJQ4u2STxQZsT
trZoAkIsidP4TC4skKZpAnzSJatZPyBXrqJvXh60YIKaMBpauD+osE3mto8oAyKL
DdygUcSltILa7/77XT2JHOLqcH05YWfp6tPprsA49gsixHujeli4wdPIacx86svY
gjdL+leGRa1JPhsiJAnBMlCqczH7f2SYVEqVfDsUuRO4u4sd3tkBhkkc18SNoILx
36sUYh5pL4kRISyR5DNYPcJPN3Y+nYovxNqy3uv3EHwwS0aXXG9xclX1m+7CF8QG
z9I++G0qEK3RBhFB62DtAKq2M8Nl0hk0x3e32pXBRgwut4IngHxvszRnQAICEPDQ
6bvqwvEOGsff08/t5/FY+tkTPV/hjBZjsyzRu++6ErZLA5MwPFw8PWNA9MREpAhU
V/mIyOdhxvlt6C9ASIVqC1sKnjpWldkR/0Tb1SM0kw1ufxaoj+sD/gOyIKD1DMCc
C/nbLdUbS8/acTpiXaSTdkXa4iKTyGc7aYoc9ap35hzcvqr5NR4lWXeFHpT0eWAn
pwv3WYhBQ7KnnIi8+VGe2HQ/yWALjjviqROWvdpry/zkpffDgzfvbYqQqC6It5qU
J/uaXkL5mxibNODYVbRvRzSNZMb/wpGqYz528EXR4L5J8ZfsvPFrjBbJI31G1T2y
tY9d2EM8BvB1AP1TmMZukmQjhL+wKQM7oSZNV+jsFh3ZtX/rfsgMofFDfAyfpcNW
CTzA49cWhlS0G28BDD7jix5O23glc6OZhXgSKTFgQkNBMgLFVymmYyQUCQzAe5X6
VaXnj+AlP9J3mWr7sjDqCMjZrG5DTe4+iXuOPzgW6R1nHFHGfA53cifUGk2EsZ5L
4Xh++gqsaQz02F3/48d8q6eppJBXpTRig2mwCM6IUQJr5bi2m8q5LQuTCeOOs9OJ
Jyd5Iq0wnPga615sZ+sJeIwC6TqOUBAvN7p76M6WBlhfcY+Fw5HUvZMn8rekPakv
L4bz7amXJ6VCpenPg/gnYDNhypQTA/Zwj1houWsiPrgZWeL9HWMdzl3j//+mBCWQ
T564adpQEwbmDAgG7UU0pg2BStI9mdm4VB4T4GaqatL293oQpwTnEBaifT2+IaEj
P7xWdz5mr8ha6FRdScXMfj4VxUVWmVSz+g22nefTs7KmdnydSS7rW+cyKoG0R5Jg
JH8k/PAUKpGU5PFl4o4pBCe+8hFKcaWFEqXdDFp4q/CEHFwdo6TPYPY6q3P7/vNH
bIJmUKg+8mPQvhJQAg0P4+V+iGwh1MIDE1axUIgsEqW7SZvONpbcxChqV2yg2Em5
RQGNmEMyQ/UOUJ5T8NmOLAaXZvbzVPDv5r2Xi5AkrM1ZTE9rsfruY78iCKal3PAO
t06LFhXSTIqdJpFNYXYHU22281dio+HH/8J6cn2z+5yIbWqGHCAHpuhTj/V5j3XS
Kt0krva+WXqe9Nm5/BBDc7C0hB6yclp+vcKs4Ych6t4Uz05oNsdk/9X/fUQ9T4A1
lQ5CM14zAR6amIbjYlNcl+qN8ua9eO1mN6dpz72GDKJBi2OKUlBCvC97dVT4JfeV
jVKjMdP/VsTCzd6bvjsrsdEbLr6Ebw/Uv0/Ga8tOU6BPk0OvADvX+Mqkuc4eHdYX
w0oNxPinxrRK8IFCLWT5BoXKqVHFhbnlq4MHh9+EfThj0Tn8CR2nJZK0stQwsm6M
Qw6MUTGBMuBbb3+MRxtDhl2uuB0ucNjbrcZ7bW0pCFg5XQljq1p4MkbPKcQ72qVF
+iM1cBlS+749TxiURpvqhshSm2ogdOwexhAyAa+UnxHSQU8VCgobVtjAmARD3MFc
CYjlQS7QqMA5aw9u9eoto9XO9nmYCWcQAKaXO9NlrzUEOvzKWZcIPcDYa+RR/2Wn
/ytIUXHPptCu+sgwQ65wmGQ+3vrnvFgSl3AT3dLG4GpXjWeYqI3jdpcm311xZcZU
82iyXs4UmE410KVm1uMmpza5rK7GQn02tvpw7SbINuRWKJKTtbIlSAF644Xy2YFE
frixt+KvpM3Lq0dUDB2RCcEhbZ7pZfRediKGtBQh5VKFjzIsAe0U30AYjRH+0jY1
HHRXiTE5hZIdH6UMcdcfDdYoZF+dwUKaieX19l7oHPUuB4Nk8fhgAtB/syupYO8f
NOXAKUyzm3VtvkBnRIKCj0zXBeH/xPIZI1F9huXcn2hLdUpSV0DQdyEAPZiMc3Kt
kT/oOwlEXku+BVJ2IAR5JovP8rF1r41jdbclZ1995wSdZ5uu43jZve91QnybLyNK
qaQx61jXDRKzC7ViVaPYea0iSQmyapVRtbcbaxd9Xo/kD7lxBJBhAvxUnrriGvDN
BxdnNHjhW+s6K5zwcGi80mTUNTrif0wfwlQ5hCrdo++pwFlFs43K6PgA9YgS+TV1
X1U0mhVOSclTJRA1ba2p0soll+m1lIsSuuSTTE4PX03Fd0aSWGqkxUa4TezWdk7N
JVTyK+YgTGCI6PQMYq0kAnqzPk0AaoXWvzGwE1nd5RVS7pIHaUirV/yLDcBTRfnc
VLcUP/bgsrQN7nKoclUN0anGS3ON5Gva4nXLhrIWzTArQO+unUdtWretYabF3ypf
fCm1Baf+jxtMyHFWy3KuiYrL+MLcqt6ux/Ty7pxMHh2X5BPQBGtVROdgygcsZDoa
s7yZvu4JKH/An1k1qCD5yhzIoafgs0WxjGsqExwo4WHFzCul0WbRNnn8VYktIPoC
HXanqsvew/0N11sC+WfjvIBaYRO12GHj0Hbx8MNEg9N096J9WlGhgJca+N9QsH+B
xvhChf0BHlmY865eM97jRShpNjI98qJyIPMbhbRYTtEG/2L1iqEm8NzYmqdGeZB5
cGSZTfE57v+zJidEy+GmTWjnGSxLMkuo229WhDZzDNK1vAw3hD5QHOzfxriCP+57
lExDzAeoEFI3edzFd6qyBPoKlGAkOvAOj8TLB1wrYAGcqX8xXdba9dvB3Q+VamXg
/nrElvUcWxU7L8Q+GRIzxIppzxpGy1rhb8vdM5BeA1T/yukljhkRngvznCGy24Uo
TdQunP0LUzxDww/MNslQx0I/op3+9qPc4wzlMcw32KH2JIDr7Tp0Kp59XgcC9WTy
YLJY1ATuLWxvCnAnq3VWzmZus8X5Iz9r+mls1LhahEX0qAq2EoLoSHYUNKsbTv+K
goMepw1DN80TC86LHfnXDTjm1aJXeVSznPkKS5CoDk3jPt0EdO62wXcVLo3bmtZk
b3uiPVahDPlbllk7c8JSAZZwT+GbkwM1uxUHzQwRUmR/oxPbqKQ1WPbFmet9sFdr
cbVC+3O0fFRZ544qzjfGp8jbkeusJUOKLCmkYEBzlPTPvuWtGTUzslJDWvstgiPP
AGA7/XHkTgPAccE3rTojE80Mt42OdHhtUr66GocTliQmWPPxNKfgCn/gW5lIlqUg
j+lRkzc1hIrLGdH1/IhuwlZRxzbo4XU8R1HLBLVR4/w6gO9gRsDij4FQ9vbBTvBy
qOTFNCyzM/zLxZSWVF6kCJdQYJsCKJhV52WgIH2uzQ11o6Q5J/xP/Iwbyh4FZ3iQ
6ypkd68LcCH2qGii1PRsKA+Nd/vCpZxEmtl9QQBjQg6elDO+Ra0NLChVlEPxe46x
dqKz74ajMgv82wB2bzEPA6uMp1L34jOy6zGLi0ZakUBBaZFSwxjfXluO5gGbdj6+
LQGvv6k/BLOKrVvzIJKT8V2R1lJzUurr+koRAhNbfWNgRnZbmJ3EA8ZnPeuC/ef4
hTiUmK2vqZecsQfh+GyQ+/4Zwcj5f4Q/0OVaA2NNRpTX5EMEwqI44pcRCQZ5yLvf
82zbvlt5xE7+38t2bpYVIlBRcub4DdZ0lu7kzWWRpX8sR4xBx/hqwkb21OAochrN
LqkEf+EakLuM3NtgJFtTyb6jNdT8NbNDCu73lJgwuPk0on28envp7IZPON1vs7B3
UexXo55+dijUpj9LrURIxWYonVG36M+m6kAaXzq5jFUBmDJuD4kQZn4EdUWm6/of
HO0dZeSIZ7LDr7zA+CmJV+vllDTLgbSceTiCgTBr+JJ75eqGBBfFwT6YjwViCE+j
fWn7n1qewfcLUylw8fevGSlRnAnQd9JcHwvKMtCsUVjy0Xt7qo1oekJBWZSgv4B7
9FciPkQfuzbOPdfhbSMRST44H/s77xFIfcY7NoYwk2B3eGBBAAly/plv+WjQMvEu
z8n/NpEvhks5C+T44uoEC0jj4BDFGHfaY1hstrZ1w83NyWAO3yiv2TeMjEcoWO3d
7vfrnCOp7qwWxp3KoQ3AD/q6br3sKbF+TXMV257yXTR25+vpeQfYx3eh9WlkXqCi
MfGmxsNKWAs7IzWuDH9Bfl9Xwrn9XP9j+PVRZKkiukn1JxGlSbtUwcLLRYXoZ9YG
xXIOJpEl7z2KrJiqIHYe8b9FgYiWsxyzAlT+an8cCVvLpa1UY1r9fKbb+GE8OqFh
D2ASngdiQw4v8f7/YQ5FDe8UmFK+aDoq6baEStNnkjiQmyKjKFtLJOIoBIyLXupr
SGFRXQLehtkycYUJwRyjsyEcKa3pWbegb+zGxN92iNNF+9zH+69RISLwPZom1m8B
/lGwp47lfR6o2LPjG1evSp4sy6kS6AKQzbDb5V3b8wneuM/ColssqNtDNF2nny6G
5Fl52OB6Nlzb/OZhIHkAtchuP2G9EliGOcYLv/3VKP27TDPyaVGL79AasF1QMSHG
yHn/vn/mKrdVyFztgTw3AC6IuwzBouQpaWKLiGjfufbeb6oUoI7J1GKxvN4cSFNX
aM/t78lpXOn0GUZE2zbiFABFIBqh3KlAS3LLb21paOfiQSjRYdHEJiIVxg9iPT/J
o5YbpGYLzwFsDMQiI3VMtmnIsqMPWmCTN0N1VbZLu9KNFfe19ptBUqbOnQJ36idS
6CyoVR2WILr0Fx5J3UVSu87Toz3NcGEdr6YLBZ2PNBcmxyqDUysORkS+lN+01hkj
2aLwnV4rKuYVzLFbU2G6axfisS3uGn2epwCJZajvwo9lB9PuZ8TTObU3cYTeCP29
iXmK0b9l6VKAux97WvyrqBwD3f2vcZJ15bTePTgY4lAgORUuQRSjzi2+LE7a0sV8
oHwZKnO7u8uHYhF3geYE5rkW8Rc3j6cBEKIaEfnwRXyjGHfcmobNYPFikVWCl04V
6UnixMV4+QWe5iD7IEMIPoRIA2M6XMPfd292PjQRhFmCyoj27A+HzW4PSdImWZ/L
1aQ06oS9dpzPIlpkQuDRwgaHkMr+n1o5oK/vEK/kqKmQ7mUppz7SBiz6Jx2ebhAN
OrSR936uGVJajY3i9hYtLiP0ZwqN20CMRfP/q8mVS3n3/QVGdfdYxVeLYfGr3dN6
GQvWAwJ6lraRIhwP51Mhd3/SDoiijtLggGHeK6/Z59tWsoM7eAIE+P8gBdM0pBZu
urR7440gAW0dolEQTSGP+0ITGUGs1ov6hiyP6V7YL30xZNSxIlQqhfizR1DkP+9Z
S8G/FUDkm2mFCT0MZCkMzoNgpKxlxAkzRtVjCH2/0KRATLAj421jDNgJ/2lma0Ii
oW4ok8Ams5cYlhy0qFJx+cl3l30TMqTh6ri2Cdy1RKRrlhpU3bSAgy8SzTH4XU3N
yPpmmVuhnT296gjuf5Dvx5j4RN2iM3EA+S0gMBrRS5iwBc7NyLnUnkEZwZ46eQA7
BdJQX35hlELpmI3693MA6iWgzdUoAMOjV6UwFCw0t3lKA8j6skMmy93lObxK+i0l
Jks/koSo0w6HmK/gYsnX2g5jqqLPq1+dlggB3XYkdCc2CDMlc+Es7eSU4Nx36WPn
eShdseEFv+2Re51GHgw9MIePKXeUs8IM4AlgnQpx2zSJsarOBjUlTe7HOJ3msvQw
S+RIi6ERWoWRyMezyKyelTHkptUy+35vC6qLPFYzBN5pUu1q2VSi5Z2S1Nnc7N/J
3Q3u6YXuzcYNks2lUiJRnmxVlqnKtdJu1QPsayEpup7zo+7M6QEb5jJdeILTXp/p
rRFUKqpu9ZCSySYGJ63aJDhy+7zzhqcmNsSotHUYnpoLAKRi/bfFMnbCKsT34Z9q
jh/DdPrp58L6y4WqVf8crt65Vy9T773C495ym72hruQg7bm2ZgezGGNo8fZ4UdyB
02Eqk6r4j6rMdBwnfRHyD6DuuY5ZgjGw4cQR7cGZ2azwhVNupk/sF3isVVwAoZkj
j+WMSVJSPioPqqx2vnHaoFCUYmc0piPk5nb/fnokPUecBS2F8RHL52PAGWVU6v6H
c6Mjr//yrNMApus969Rdj+bFPwaX1S9RAaD3DdawjOoZ/gVi3syTyfEE5uhoXcWz
de5FYeu2SdH95totFhbarFnK6jc/zgbETyptXPY47YfxCI44f3GpcVrXlVBRrSHg
xjNhlRbWiLtdRpi1hng/1EvEI8ZYwJ4OkU9mPuTMpHYVtbfT5emLmgj1RomHYwi7
64k/veF229Szjh23eZclvoTlNPsyBsdPq8hvTn8O/ei2HTXTg606b25xEtAOpu5J
1u6W7o1l4KSq3TEVuJu747NBDgKvVIk2/AJB/vum14Bu+x/iOjU8W97TKVpm0UCJ
WSW5nTSJEUtMiG1kTojgb6sFXzv9Rxwt5wmIB28rU6R45te8BH6uAlGg35iV7B9J
Q1PuwVaxVSu4oO/oiwUrBYEQZ55FhQY9NsMR9T946z/d/1T8bHllUd4XuxCnJm6w
UEkjGpNZH88NZVGOYyHAwFoFrHerCpM1Vot1nqy3fJbC1XUXOVFmZk73JOk2O6ZT
Vfa4wBKNKdttIz75+VgqKvZETh4aQNLY/49ROVvBAr7IyNBcphYMpYo3FRKGUF+p
sBuUT1buLqMqboKEEoCgnHqI/l28XCZ6Sgrs9cv96zkAbM8Cf3Ub3g4Wvge3gl9R
5vscUerC6vD9J3ITgFhf/vVUk8R6Hs9nkdA8MuHU19YKqycEu4k+7cPXcavlJVh8
a99fnf8eEaBNqi/gG5JPN3tpvVhsNq3k61MfT7Jropbvft1nHlLlW1xXQgvKtA+q
piocP5fgjEEO9wvWxUfQGF6L8HyAzUCue7lTVCtgAXzbmJuTmba2DTroNADK98y1
2LIePYR9jA0Pp/BbjQLMC6R+/j1kLmrHiWJ4iCO2DpOfbGLKAxx1ynD0MPHs1pbI
hlY1qK0YytKisUhdAnnvLatbINmxuISehOhCOW6pFuJlPtCkHuw3QqI/tiTqCuJq
cjdDx0J0vNWyHCIM5nh01msv94qTNQMXlWkG1AoRgHXEpqPEwSSh+KBm2bVG4QzZ
FhJe/4IHME5rGyld6Ayj4srwgAMZymt5YCSFSHGsPJeqqOxXX+XUbunc7aXqZs+7
Ij6BWHjCzyuljoDfXEuqFMEiCbLJPUWZE+i3hqibI5cb8wmHE5oGqCqWqih7AqyZ
9100hSE5/1/yRz7DIylIlFNgoukjQcfkATv5pHmFaf9Ik/nnzsuu33wrNT0g/KIE
0fqsrC5X/HS+DOLNyj1KAvzOT653bY0llKLRNpU3zyp3m/OJiBlCW1eIrb2WT0qH
585oYNuguJv3WxX3GxnNKOIkH2nLHMQqvA4lzCyobOAoOX/6L1hf0VxeljST6q0X
5vkiMPhNucyPmHeC6o/31c/KuVKroPblZ+rkGD9a4AnGFkpsNOAsg3RZmNlvDkEr
J+UOLj8/9YGeVKeCuHNkVEnb9wcuAHoEJsEAZswnpTKVGBB72+UWcBVdmWXJOoiS
09sCKUDpplk/1ohet5KBjjkjqyaJ7Qpl1tVIND5hyv5YMHl1u9gR63QKHFDXYEI6
htUSjuP8g30q7cFBchzWLSVq71vBme96TUl2jXEMbV0863peL37+IgUw/lRbtuZm
RjwBXLwnFFa1gSibFtmSauTchnKvTDpvofb2npmg3+UQWpaRv4eX42mtFaJNmAyr
H5cO8hJjdWqr5gjofT6xzv3tuNwAb8Qu0lZxyOq4mK3tLoy39UkTC+GuFqrFaFg1
bnpFFCB0RnK2PF8lXqn0GtqXjiJrwkpmAvhI9ZQxNoz3JEzLWCnnT/PFwm5WVXsY
QbnUDMHM1BFmzlVJASHkTQyk78RLbl/VxNdPoAfOcrK0atIxM3S8idpbhkWQuO0M
h7bs9YLwV3Ajfq9EjY9jfWV5OR8t0RyazmiCHLCtXqKeJKpxQX1J4s7l1RufSNQZ
BMgcrGcM8ZTqhm6qc1V/h0zXSvHkrhCBFn/wn2OSsZqtveTBpsMG8GQaAi9Ick78
V9H4YFMW4cZZp6FRGeudX2j2o96PRlyGjss+1La+vLnAT80Z+BQv5zxWKXbaZmds
YFkeG2oohtf+obArdoRXsOUqF/2v+TfbJzBj/ks/3MPoD+jLRFYEtS5gP1CE8IZG
TS2jjA2FdrHZbOrHKjVP7R8uZEra2vlNHn6LokAUa1WPpAKH3CtchVU9RI5y+pVw
zqXOy5JJUlTw8awU2EVw3Q3N8UXp2lAnX7FCcM7lLM976Xrf1KgZ0oq/ocnJC5nZ
ouFTF1bcq8RhXjCcM0dWCXalWthZiB4hyjH7ABlieVdovoDvBOYag20oYi/yR9F5
XM2fcdyvG3kaN+pso2HrnMRF6bo/Irl9H+C2GL9XX7YjoSaT3JpXpYkrFUCdkJ3e
LWJGoZhmfKg2hJqoZk9/jFYYhaCJFYv6sE2iZgUMB1FtdHVOTMqCCO/0MkcmLp47
WX1Bp9xqeFW4L+OBv06SymFeJj7pOzGXczHsMqnON2A63jt/UT+2L5vF+4igoNA4
UgbmclZHuuCE2Z6/OgQFKneAVz8OUbzCVS1LBeECSx74IetyL9+iMQ/ey6vWKOC9
xMS2+C1KcRZoKSupBXylIKreL2hJgwGkVua36U1weAeEi6R2IpWQriAccKDN72An
LauQCLO7Bu20C9XwigTRpEaNlWnUWTZIihKSmk9yPsiE9gaLdb9lVXwBpa7ohQp8
XlbEimefGXtsnLRrmjiv1ujuUpkidjVxMY6VHqIb4iKsDTIgzJ00+mPCkqIO6Oci
eww2ew0b+TI4+QRq3xhZ0Do5nWxd74AOh/Rqux6ZneZX2eEqaGc1nGq0fZLHkEoe
yUJzqksC+AalitGxynpu4DinCY7LCSySaXlzc6bCgPS1CcAYnHk9NfUosaNuf9eD
ACrzS04KqSYEeXpmAoof3jMZp4aLr6Dcjc7gXyHT4NBW42VJe0WJJ8IlTWyu/yRv
+Sg9YmkSzdzd9NHI8dMktw5EDDfkcbYHhK68viWWvH6raX2160b7HcEKAi0uG3s3
lhAuXyszZS6y/A4l2C+2Vpmr3s5u8+Nq4tDw4/bYCcAcyiZEsk7yvmqpYNJRPzRf
UGczrRZ+F+mz6EsO+1INtxXKtpHOUdJp8Yd/fA/qUGK4cnWD+YbxdUv93UoxUVMe
bqjJYsRFiiM2udzYB6HzWteP0u13KY1aLM9JrQIfJOQDN5TNXxsj8UCz+4aQu6Ml
CU+ugBhIsW4INEtQ44NAJuH5L6W6gs4Mp56rf399USlIU+7CR3PDojZLiFLnLBGQ
XvFrw04z+u/Mz93ZqdaN4DBUluXURBTp3wG7lCrXMZBQNR6++Dr+hJpxjjuKdhHw
MjLoMC/vFzfXQw03yV5phBxW7JUOWGCMq/lq5I02N3GoTbGz5362HhTPvt/kqspa
Nflc2/Y/x24Q2HO8rMUTDQmR1dXxZqjtYlNTT4O6LbLjNZwkTC8gMiIy91SAuPqs
Y+9jl5zNLyNwKHOV/5eCreqXTZuCjcgeHwcaQCjzBTOfpWPEYK623JQu7xRbMV9s
tK0/vpk215vK2cbEY/VCoHXgDfBUJv2zslzFARCGc49YOY2mTdzEdXNXGMq1nLNS
o8VfDRBpGbnKSZe88et0Cv6BO3heJVYpq601IpoIt6KBaVC4YUfNXkF3UVek4WEG
dp81+dWwxRcgUzR3SeT8yefNBSiwNJ3bkodnWYwnqynwbaNcaykK5swKAUCT5cLe
IM3ZOStn8arCFb02oM3JOfzQaXu0JRC+c8FR59DlJWPxvsFRyOLrd4sbbTjdb3dh
W67kyNsW1kll2oGw6aTdSJveuoNkWN+E/9E+VhQnWmVdd0NB4fwQb4r2gZZNWNJg
sIXryMo27PzVI9hKqGu/6P2jKx8n0UgaLGPkQsJeDETIaB8nHcTfvsEIWgsi0FDl
amRyTiO0BrkQrGNf++C0bnkp1/2NbLWpVag5d6P3gEM3wxI56xInQmbJ4Nc3gzFk
H+Rr7leoCaJX1aIKEAnu9QUHDE3mQDZ6m1DVO+1RPtHiZ2rj7mpATqjtRkInd5vv
2xNGPaFT8/8xYdSCvGr9USyBt1J7mnPivY0Bsdh1m48l2K0dwpHhLOe0ByL4v4Yt
/zsP1d64Yv9eVD/UKqg+xNl0aJ0F92OwXCClQKZQQOEFVFOENwfEJqlQVOm5aukT
5KyDM7itblsijsqMLjxjc0BoH213AR1sdsYQ6pQx3Hpl8UTL7/rNmgkh8D07KKk+
6TCSu6xbE19ohYCORyBS1slUvKgcvBFxLOrElKdLedfItRY36maMpl1Vj01H85N7
2jVD+ZCjB7YS/BsMcpltNDdGJtn8J5aODA80ITAmKM+9hn+YXpJTbXdFmk09Rptn
g5YkfpwrO5U+679is3cBZCLFYAFpnS/DxQpbRJJu+6ihJaKGq7mVmVouG4fSitPt
2b5oXr0aIH/t1YnTfQ/lO+F5psuL74FYZOaEsJRfmgFRIneZp0U3/onoPpIAmTM3
CqFdhQbBFAUs1zh5Kn/UCcfkgUkfugceNqAJc6YDPUYbiGLDngJuf4p8TFpTgYzV
FCVzdMjrUTuu2hfmC7adZXHXfI8lsFxUT9B6cz5sf600rubhLD6pO4wXJKf2vrRG
sjEC8qTd5/60ZGCjeroh94U72fmiVIrjgsPs7NPPL1b4KR9qkeqLyA8Q4omnEYQn
ZRJdbI9pyZSt487TJticeTBWPcO5GNoOwDHrZ6ykQmcMb2X4DFigwvr/aYEq01Pw
WSYf1C6zHZ24d3XUtRSqigOpbfaFtUcDWtZ1EWIm6y5LBEvR9WUv4s6ARG9tOf8e
xkAxyWJkxSQTni953yynVzvJ058sNPWJq5zlPIBMStNQI3s2z5AYSLRknPzivbUn
xcaWHWH36dluZoVk3nvIm4JC86O2W0GkupWxEoTmQUQ1163BWEAls5nmwPSUBeXA
H04m4ChkDmfNoF1cE82ZSrQh4QuMZ+lMF36dsVlOCBW1rWJRVPzYFi6jfeSeZAlT
HVr4YSDeOi4t6LDa7+vKRW6kjnbWg22Sc59aYatUw8Mu8CemhgJdxO7AFaIcoM4l
pNnhMWnjio4iH1SBvrG/zq0vIYsaJ44uM5jQuxZMyhqvxr8Rfrv371sAZMB6pLD/
8Nl0bu4lbDeKmSFUy18LseoCT1sw1QO7lxuQc6PCvYVw2qgrYuZ4kNF1vx6R0/yP
FSHSA+e7HPSMpKEJvNjzUIzFoN06o7g+Yom47/NQhK2xbycED2/YUnldaTY54QgQ
QJDY/j3m+uzXbDT72yofkwZ79yfnsbsb1ZnQ6BoRbbGqzl3Vy7oMWLj6yEydf4oT
sC0LCzqvLgauOY5Z0akz5OY7JR01s75R5S+xTN+fn0DAhEhYC8Cf3a86KDMBRShD
B1s4TtmM+w8i24xC7e4AhzT6ffOQV/ef6PJy1d/Y9CbwtlPgxZJp95hYu5mP+lf/
ZhlAQySSr65FezDMdgSYHzc/SIVInQ2DVYh0ayUgFgmp3F5no2HNi1W+QIe6eQS6
Qelz2d3HQ1pW22qqbtlkdUUCJWiu6awD3ZKRRNVamHbUVtQf79pVDaDqqF3R7PRC
y/ylIPLbtMBUdOwNRfrMG4azXYVcC4HuOb6MGDui1dkjt0Au1ZVTjNzV2cX3mYQl
Vy29QZP6fCUa/cCOR2IDG7VFG2Qg3MT7Qj/y6Mxxcynoh1Wx60nQwIxh+3Lo3mhh
E3VpYSI1/w+N1Qqf/06TmND9KZkGIEiLL5wkEA7kIAxogn9Q9XPKdMHuPrgBycHG
FDIzknLXAGqifY8ahFTmzYM1ayGxWd1sUYuaKyPtLk1cPaCCuUupZWO51A0MpFk2
AxzYrXw4NSiUF8hn46YqRVLz9sUYGcBaLPe62tdu1UyGRozWgR318a9KF4GRMc0b
O4Wf7wjSB4HekhqT8Aq7V7UOGpGYKqDURiCAvlYPb+WS5rb9RuJwnfdt1kID4BXW
qKdBS4/qrTTXb0hEn2KlaZumeCGoKyvd09GjWShYrTjkI43RIQas4Pk+37dMdyOG
PxKLqxRn+y7D88MgEprGh44X+OZLkTz/FvndQShTqGVYrA5nb5UX0X7NNYTCbSUl
2ek0p3Jx7cSQiYolNVG43FwFET+PCWQZu/EOOkr6q6fSuyh4lZDtJy+CDiVGgK0v
xlpoAdgC2ec1UeZMTXRCu27igq1G3EWJ+mCoZHv5nV3cvmOp963dS9rBQYJuOfCt
8v4sRBvHUk6DmY0AYD+UxKTlhj04MfJJmH+Fe2WJZ20HSmzxaytLXwKY8IGU1I3q
jZuD1h45lz7KBasPKaaikcJWTWy7aVt2yUaCsmu8ARwYM7m2TKE5fspnczeqdUMV
XTXAvSUYq0ZsyLNYEiiwsnNWp8KoMEvKPxWuIEn7k2+UPzUzLp0qqvvJYIzP0h5z
aPj3WlUyUCSvlT2O1aqJTlHQTdZTUFLMJT2MWzGf8mp0D0l8kmpzrqUvZ4vPiROS
PjTcPENP1/5iuSCmMqEB5ChSc4Qq44hCDA0KLoLlE1Rrjz6xNvzuxWnaeCvjmeJt
wW3K/GfbvQ2HQF2WIkHCaUK84opnioed1t1N28zGzkMiDVHQr2UwXk5KVgEo7cwX
5S+GGxoPtG31y0vc4VIlb7whu6cZbwOxfEOJwj6ManKtLj2s5bqDxGanNTvjIvIw
yHltrAo1Seu+ynAr3ed7Rtqd9d9GLYDAcQluQZ6I3GLLnKUQytK8Yi0PtZaSLJeV
0iku5VfCXg0W/pkuGi+NM8eBaZkTBtPIcP6rpBaY68E3EMScgz1UAoOxFd/1KibB
qyQ/m2jbUQB3bn8mi9GZB8PSDyAXc2ZONy6kiaS/aMd4tDvtlbxoqK1TQEah7/B0
TpXmdoeX74LdQkE+RGDJFbTRrjfpdPUvqdM9Sn0b3WTobiZrm+8S4Nw6OjOJfFRY
ouLO7hJJfgyS1tArfWl6IrTh7pU9csTjzTfuQ57Y5Z15wd0Xx3kn46SeJkhDdkQF
zgVV0U9M4ATDMn5P4zrOWhzKCEEqUfDOxmXSgX0gowUQUyE5/o4NQPiCfALFn/8r
F6kqbdwvlxovL1dC3CSkavuGYEM8t8lQ65UPtakBaJoiGxnDJTos2zA/Iqo9q7BV
UGxRdlpuyvv/pTIqXXqnTlB4z604yuge7N8kTemhGfg+QOp5PgH+3h8huM9IfiTg
wxGIUV1nxgVmF6SIKUM91oj+N1w4P3sIeSSE+S16TvUsoFV8gwikbJ5UfHDopwcz
e8wy5+L33LGCOEiwuoP4Bv7nG06Kal+CIZQ0Sn25haB8xNxqnLjPmyrSWRebtwae
d+WuzdG2oPFsemos2de9Ot6t7TyVYVCB6e4U+sSkCQf3Q7nAVNDGcmBMSIMWi7Pv
q8pbZ2jpkaCyIhajbJQ9twK5UfFLXDm7p3kNCvVaxg2qnM/JkytwS9tPiFzIzEYm
t4RcfVvdyRudPSclg4/yoYgxAG5oUtO8RYU89KpgiAXU/BrCiXkpOmfWr5X6RSX6
wLRkWssscs2f1lPRDaOQ4Uv5N8OPbqjV6rwR9SnlNjzhjGqjqhpViSEC/cu6jpzP
vTejhBSCTc4V4QOpnnT4Hhce7wjpMqGExIGR1F6ER+B9XIcWKbt/rZ2cMxxDDd6K
jMMX43zjDLJOV8h3AyLrjGlGHL8b9lfIlUiXmatBemd0I5/CguuPFkpYEd7thNgZ
/BYzB6iHulI7jDooc4Gh+4w0YpJJolvKnebehM4UzIvUOcF4Xoo5CwR7Qt+0Yicz
wgIasiM/7ptgOJgHWVF1IQH3dfxZmVLDw++hD3roTJLhXnY1wZJdHl7tHUXB5Lot
nBAP7k35JzDvLIAr6pCI2mNHAyZFRUsYmbpc44mwDGsF3nxJbTIbnogbtW6Q+e+L
fRJvs6Ebxk5giYagSKSnccaHNw6Zy/pcT2MAftOncUV96Mw4Hmu61hbV+GS1dHBS
3oVZIfIOt2RMhYXPw06Q0pFCbomQQ7zGipQic2jLrUJ2HlK5cYIAKGiyAecZjtxN
kXN54myDCBT3Epi7uhaYk2eoZT3CLTilpec+yZ9/B6D+WSe3hOnD0MGEBRgB7AO4
bRojRBzPy3BrnNHpv4Lq1XUXtzowg3Dn+kEy8+0XAzbVd+niVYqWOlmwU4mX6wOg
w3t/Jn7iPgMfsSL2Q50Q9bj9szjVKxLOP3ujNbUCaunXrhLjKJVbiRbANoYumLV5
YTOkcxYnIGA1G52Fd2zeRoQjgf0sQRllvYiYNLO42EOMf37dwoUzFaTcG9xAcdOA
/o2l32r3UoNGLNqddHAsSaj/hN25DdNwht9W1zjjWZElhouRW5tGMCvUI9EqSWHY
iIF7Qu0YNLde80DKWznPL37r/hhk2pQkrDtccIAmRUfatgxaezYcVbkXO+XEYhfK
ZOZmUailngtkPwI/wwlG5y6zDJogjbSp0hc2xFmN1tJYzEKmMustWOxpB8ndFUxx
iFBk5WhGABWmE9DjGj4pyTtlFwETefc41uS8xlkN3XpNbKRX48n6CJjm+CCRgLZm
LG1jdZik88XGGYgVVlI7Cl0bVIjo+A/4kaTzpUN5txVOa0m0oa+XsqeZuJ2x+F+r
cERfzMi2sQIP0QYtCoeTQ+gTb+4e+JC4NWlg2+fEMHVnjSgzrCefAD3kyZ8VP3SO
xkE991vcVElNZ0ZAHLpzAD7N6W6TMcpYgEgqv/iJ0/erDxSVVLHcEVKNOrGp3F7k
Q6TkYIIKizlri2AgYgn55v64H5iiTyGI7Knw4BOlk6hOhpNUiuQHz6dneIvyG7+E
coKtBWjhhJEwIYXbQ3QUCHf5JBqxyvKUZ5ZQFCWth1pfw0Mblh0q6LrG6x+npM4H
J7U77gyK5kPB/rxrxVmTSV2qmAdkPXGUqOdLfbJaYjwqUy0gO8PtNXweoJWdtnmc
HahHYC7uA3IgIYTSSAnikvPJeZgbX/1cH+VQU4cSZb6W7GSdKHrpNZcjYp0pOAf8
cI/O7RqOgqKmdTHXgQNIZBJO2mtmf71BexDJV6KdEoPnUzC4XfgiBheJClwxSgeB
soiRqWEGkFYSplztmM4cJirmNoVFXnBec7yrL7L2qDwcP8HSHKYl+Y4gk/ONsmXo
FTAurKljiKR9U9hkv/H3haZWb6S84N0LsMQgW4IWdLDTth3PDmrEsdZMg0uGV7IM
nnqj9gnupIWKvNsAniEyjX43l9tLvmNKdmmPW6egekT+LGMtgABvqvw3jT99Ld9Q
SgVoj+ilssSAzjduRYSssv12QzCP7YU45qbuhDjw95inxs4xxYONx/EvpFvwbalj
NiegM/kd/SiOoJlYE4tDrozDD002GR94PgbPNot0WGzkYpcOR+i4666qy+84jmqD
ldLU0LLYlRq/qr6FoejQm3/kGwGopN5bOcimJvaHIyY3oN3I6ZY8Fu3zlq4a5/8e
Eb5W8cvwcphV0Sava9c6xEWsLOn07o9oip/21EZubkyLIuPe8GHaPYBTDzvvjl5X
txJYbXHZSn3Ayf6fNAH6aSfbXZcUC0VayL4XzeXMwSo1hRYU1dBrM5y4En9PMoDg
rv3/rjWqPu6UC8XBhS3EVB949MoZUrre3AjlGOUvQi2WNWxjwRZjkv+eMcFAGBpZ
dY075w6VL6SsPEHHZKmtjjMkihhWm7tivUUxURquwxl1/i3sEVS3MiVJQ5Cpiq6m
KhPTcU66bwi9vQoPV84ww4+JWnrrKSEU1ASzF5p45JAdvd2nvNhB/PL1bB7KOdnU
KETfN9oqM2/QyHc5VYUmT3OkQ+EqbzyAVDYtlgfBAanZauSbmq4x9AvR/8JrnHQ1
13i2AT+4oHLomVvANRXZIE2iIUW+b3KgwGcR6+pufn+8nxLe0b1IXEgi+rhL5pV/
RCFOs3q9Z11/a3AbKTTz4YS8ZbuSsR45lYfOM01arh54FWB6P05ELjfLlGrl0Zj7
ErGi8Sm36M7Eqisk1UKAkgiF4lw3eAqHLOFfetujDgowRRtwe0okJwhurqZVlbij
EagDFNIvVVOGuV8IvJxr/BbjnBQTi3FHafnKCbzFZusSrEN48WEBnPSD7mxah/zQ
JMuIddtInuc22sphpFUTfAi6KlPJ+FsBisD1lJ03nXvkk+hF0o2a14/KIh1X/CAY
kyiWk+Ws+58fYtD87agY929FnD8mBECTdDBJYO4UFDVTevKhQC44qSgwN1/syBO+
0coPHpkMe4XlT0AiQDoQ1GQ6iQuRo174fp1witbEXIiBe9AnxKVfJbvb2raKQMrW
0WsaD8eHva6DemecBUHojRrsv9Zol6QKsgrr0qH72oRN6m1Fd0E+r9nP15yMscAO
UIuLVDhTuz9GqRjJHen92TNx12yQ63vXOTjTxg1IAy+5rUkwhlbPYDIA/HyJvGKo
HA6KgQs7LIW4VZaGCNNnZH/dLrZblARfpXgsoB71nYw21sqKAs8dolJVYfjzjmdy
y//d6f3i2vRveisdq00Bnf/MZQsbD105Q2WYxd9861dOZi8cA6omYzRgnK/2Nasy
hanE3T3lVGLnNNYTvIjFh7Zon2K1tuKevQNxY4s4263q1sWjr1tQ9ekb6qep4QDN
Fkq8IIzyt4twjmRLlKzd0MqiaNyAkD6NF0QRawUWhdwUIx0/XZfkyOd7DMBN6WZd
6wemky6In4sSov0ZjE/4jQNt5j7gh8o1MlRtbuzjCoujTOAyKQwUYZqQH+6L1/my
quqcKHuisYdN+fYgKRiVWjWDkcmETADHSThRq/pMjKUKCeXuSFcbZO58aqsPLVnM
Fm0nCRBvxdEhzV2yiW73v66GINWMMUPRBumgguhnWxOvQeBFW1n8qmW6ptyovE72
h3G4SbDjm78d55QrypKuZY9r9uMPq7DrNIns3KTGgDHki0jjakmdqiOaVLUtFQ2n
XoFLXDOHhqkuQLt1Z7TFGNy916zKenRx9QaEtZjbaYdS2CF+0iPxz2bXhpp7KKAA
+60inC8+fZK4TXQZALxAwenPDsdqDTwwGCvW0km8qkAGcFL+faXNC8uGJgXTLNTs
iZH1sFRydRha7Yf8W01HXp+X57nw2IHwmxC/PfTdfaY6OAheNLUfFz4NWEjBzN8m
Cw7uq3afPL5pd6cTY/zZP3G3BxVb+R8vrbOfd2jWrM57biWPFvVywXZsKNO+WI83
BCVkR8leSV614mJb/EMuOON6CfqaLn1l/609JDILn/CkTp80mfPKKR37UsXzs8bw
a8zZTL5MDSF9QITfuPPoJbMyF2kXIa+ovsG5Z+1zY8DkW9NJmbbJksUIkHt7voUh
RlV9sR4ZbbZbZtyt9C0wl2aH5FInzrKVFK+3kTvHzDyyTTMrXAS8Sle4rxHyJlfq
M5flQAIyZ97LPYGlhEAMnhMx5BouNrI2VhOB+x6d18zwtxGO/WPoIXqo0aUZWaqy
87ZjqqTeu117A4TIyRSIu2+1fANn5cibeI5gM6+XbpNDiqf/m2rtzPu6qGTq8DGd
oVfb/Src7N45jve1uROvECvl8C3j266OOD71tIjt5dqhJ3Rgi0fIwiHk9lb+wvEM
MFv2a2bbiZaMDEpvn1lZrzBGbVJ+JLNsLuYlKHErEXpM33WBi2/2veUOL9kmFhXG
r5D3KAI98RHw3XrJ22r8kvSi+XAE+uEv0MfFzxke2f4SjWnmGS0gZvSVy8M+yIEV
O8zyxa+tWQ2NxgUl05s2l8LM54Ea7I5MrMe0emoOtjAfKs4tLzm0vU+gxYQhObch
E5QisZGMX8bS0xaIqhufZkocZygMieoiWOF0cN16VG2uats5TS2C56qmvthnnwys
6mxj9bt2jD5V4SQJOBh6GperHrSUeDxvQ0FQ1MJyfhOcQO9td+mAEE/pvcp8IefF
RGQIjA5/0ZUPH9A4jd3baBy47/66tbXKtGAY0BvPrrpM38PqZ44Bu2vWUHzD/Op1
EAopw3RpggJ6nNMBnjK6IMCZIaKaaN0ZIADTcRlHg8PsCTJEFyt4Io7eUBR+4lby
TIBfgMWUhA49xecgBjLX2Xn8yQLgtQr35aDQoFdYjb8Gd6htxPQucS4uzv/G5Lh8
VtOHC+V//aW5h94JEZCka3m0nBnHvg/GZ1ieaPkoFK4bga7zNRLt/kJISo7ECSan
fGsatFF+ykTd9jArxF33VAhIebdeO84SdoViu9yAwWRV2iY8DlgmxicTDYXoF7vA
w7tBn0xYwF19KCBS9oX+KHX2KrSLY8UdiWcxKO3EXC+yOJ02Yj36j0r3TTF+hN6D
1QYn4CZpZV2y85RZor4s58fgxMX1TDvBX8lUdweX0d4jVOqDdEcC81OFHgXPgO9m
o1MJlIMGbjoJFKXD+jtFsxt1auwmg7EHV867fmoROF2TRnstTtbdk/AI7QmxhAhf
pre1fmd6F6+MzhE0rWFwW9frKKIsd9Gd9epq3GxOCAShhUEc59FaWN+3JQ707s2F
Z31kpJ8DdP+QDyylsL1IJ3TAa8o/85qkfhCRW1gbL++YnUmwJXiUx3jDbA7iuyxJ
04Rwmbklil2L2OeK5kgzmsAYm8dZpl4WwYSHRreycs63xgHqRkY2G14QJK0W6Uig
LopU1taRU0Gb8GVQ2mTrKHvsg1LKnbBr0d/iokBUwHLzUtl/R/ecaJmES7BCNsi1
3xSst0YBelrXxsQO2QHbMdToqyrr9QeVOuLQM9wiuVmBKFh5uxjAwoaLu40k5/UJ
mphs5ZI4J+gDjRLUnMw2dN/2C2q0a6SVcIC4FDjZocvGSHibhYvGH8T8FOQEw0Dd
d8vMbyRZ6A26saGAUEUTbOzDffw7kHohz60I7j3rqWHb/yuOQZ7v2+Edx57KNUNt
0COnjUmBsa53wtvntUxj8Z9R1XwkTaQeWQVEg5sKT1eldhSUdsvDz4ky5W0/L4em
3DO6MDa1Qxpw4d7X/u6GEUnToA+Kkh9UqO0KuFIftZnFBkRGmtupfpwN5ccfXBuB
P1LUa8y/JWJbv42i50Abvh15FGwtOG5FGhRa3TGhbvs0+bBFB8JztFWViJ1oYX9Q
pvLNgKH721aeQWaVQREQ/G/Qwg1UsnpiNIEIjbVKkSpRg6wtheskEn4XbwRj8485
Tii90A/+aNJCJcw2tKDvywiUJVP/2/wDDEfcXsjhNNLEJghseMUM5kOTOpyTTzWl
VjhVcsspoSSFCkfg+2mKGhOgDha4Xki/lmxsmqoEcX0ty2FCOrZuqMVE2HvK7TsY
D29VcbUDF3DzW7fbais2FtHXK5ca4b0fJwZ7wZ4zIULUq/WKT1RIwl8YjsNjnkAD
qgBVbifIg9fAVR7nIyeF2gIlmhUm6DzY282AiYCCfknhs8Lj0FqgLoeGt2F2niEu
Qdx4SYiuxmQRnNLr66Gc6Z/RdhcBPdETCXWqAZxcWOL7g0NvB04+jGkGbgDMJ2SC
0oCTwdmMjZht8EAP78Agd3Ur62napM4DNgwAb0w1vifbdaZJsRQbfalOk9b4+3Zg
iOKElgEIx7ORoZ9N9AljiB7TaL3WxrmqbWZzAoq97cOGRPgD28EOK2KGK8JKPeDL
cpp2dhhTOR+rDV3b+eE4+xCnHyc512aZzieJdnfUEGfeFN7vU0jmgZzp2odxwpLs
J7z7IwhHQhO6nqGNWyaMtHct8UqNJmwuUwQyVM+/pRO9hP/06EWIx7Ubn5I2ouVj
fI+TA725XZvxFHJNUw1koV7744B/hreMA7FAAGkXU511+jk8l1aPefyLxwfuGG23
ZjfcJSD5lJ4gLTz6dI00/jGchb6RrlWhckPTwnx5NOLGt5xa1667Bz9xEACkTx8T
ZUCI0sjiG9HYE+xf/B45OcNoebFtYPhWvz2uGj4e20uc/lK8feTV/s4GCsaZOTth
XTorsp3ZxYAK5bOvqCV+71aQjJtIzYym9HqafVBBF8Baf/gseeUZXLPxHAolkfo7
LFkHSd/DaKH9cq+1YcHjW6CvBiM+sIstNJSrd2J/1/gTUnpqgNpXHXWB1fyf/uVI
VD4eSczxRguG4SzkHYq6jTBc7vPsyWLhuwr6/Ojx5Pc9MW0H7eziica3Bs6kTHqn
kP1VvLgUaJOtEYBeUK8EOJ4/510RUlvKN/Jx8v+zBa5ZoKMYbYzH/6I068v/b76t
Xa5C2GPbsZHzgrcUCatL5A+yXAGO4WYXuuHxvJAP7tvI8LhUqKWPh6haLFJSspYS
yVmk5Y77nWxehK3ioZtgNXDvTH2Rgvf4RE4tg9vROQRckfOWi4Qa3XClFpQ/e0Q2
JMDjYEnJBl2rgDYrZ6Gwm1/bfkmEbzZBbu8khDFLOsIZnYvOGJV6Lne3+PI5zNUc
yz6ks/ZEDB1i6DmomLUmO04eoqou+Gqk0n2LWRMKZ7qW4aO+RwbNIdb9bafM52p2
uyR90p4rKnsxsWHzRuWxiOlJcKM0RXvriWJoyvwGR8+ybIo4DBgbyrGMJRm+oLoh
8rKLEw9pfaZh9JVtG/ofgsYOLWhFsAiitLHzncJkxWZlLdq1vaezREgQkK5K0PMw
CyYsJ3TpL1V41+MONwVn4KBbBwq1F8U1hR/3nkmRQ/d0A1OtUasKvFJZaGxtNYeV
/fwhfG45SdejSAgBw5tjqp7Otm25Q9DW3eBdqBzdrUvujR5AqLnHB7CdLAkve9m7
tp6iGDxSgducGdCZzWTWH0kvpQzRJ6fUYWVU/WvlyyKf3jz2Npbbt3cc2yqYSiUw
WwwHzoaUK+baaVpn07wBuQzH7fzMx6HldJFw/kBTle6y6eZysNGA5SLV7Kpy65xp
y3iqeZnpun9CnV7r+r5DdanV/OF3saUeBGUp17bD3YWJleZEjsen3WGXvWhg6MhA
nYEK78zHll1JoF3OieAZUNajGzh+5wuIHjJ87MzV5fzAnZAeQuRl3alff/W1PKyS
SdksNYW+MavsJYGeIGsWvkAKLhtwi7o4eAVWeDtt3lv/+z2P4OEU3a5LOc+DfZ7T
wiC1Qw0WE9vjcWj/lxoJtpjso11UhC/uMLNJP4QADNqE4KL9oTDLMzdUOEh9XPQk
czl8p6hn5zA3xfX8IeIutZ/3tFmDnyzPTDocP1f2FoXTqv/ImMKJvWddd1pUjdt5
LwGtO7wxnD58/HEegSN7P5iN/rmNgM2/HMgZAwjeaBVrklAg8jPHpAFbXlc+Wst3
jrC0ObtHN/AbsLBbQtkEcgy/sEXI2lLA1CzT9JHKFfIIHjnzn7eGSbW8FTLD+/aw
TlbcgMvEWN8AyCys9DCxR3mKomxZYOoNWRX183j2icmFBDlB1ddsR86d3szZozTr
yiz+uJBGgq6BUFI+AS2H8l6pgrI2ozqdd4YV+FMG/9toXfuvnQoclDMrC7gFxWNT
OEi7uJV0E2ZixEgQ/YKjh6JGmWbLeJ+Wpbu9SM8uHrfqAmnsgEt20ZDjdhp64mO3
x0QTVUSI/i6mNyYeuMncl1/lLBI+Rd31xE320+9+P8iTA2k8XPO0iXC/4XJRpBhR
6gOmmQG+R4j5skentZEO94LHdCVmDObCT2VVihedCA3iCaiitKkcMyoa4jsIOGnA
K8OvCpKEhkSnv2yAUnTw1EHyNYksD+35Dk1jKxod3qIb9siONxICZgYVCJYtZHhZ
K2dcXOoNn02mYFWy7uyQtFvSS1MKCF3JTwGUyv7V2p3yU+8e2gtZH5DCD8/572nQ
fSCp7Drj8LVCksTNTabmsytBpQRwq0V+7PiQVH3I73TYmon6PsqLC9QNVqr1l1MH
BHdaY5OJxiBG4TvQTDqYWliIvSsp5bgxd1FKTxEGmUCHY/x7SypHVSC/glHt3/vf
QqwekIF7/FkuD916/Upv+Gp4rPENY+mK8Hxsiou2r2NfIKuORFa7ne3sOI28eToq
SoJSGtY1KdBizckPZe6GSojrPYmP/MOU85QvipU+GCJZ8oZIjpVr/nEUieO0AlZM
9IS7V/3jBkrgt+G82WL184U89dm3Q2L+LmtbaJwLXQ7ZsdsVDYQA1OPyO8rPL7cp
jrO8pZOnLCYOTj+QeTS6+DefeaCN3VlTXR2PgkSB0zL1ldi0CXA8Qf0qruZKEoCw
FKdNzCY46i6pqKGGNnwd9sxZK/69GUZBPR/f6fC0iutJDMMil6ZirJv5z2JgwwCt
6WTsWT3N27Hs5e0FhM0CceYvKgobQkNcS/lGSZKsFGUQHt+O9TC5eisHiz0/v4tI
FN9lbeujAt4gpQ8tJk681aDb/f1OGtWLOqRgyezSh5wvVUkQoQdQPqhl7NU0dcBu
61OEDgKD39LZkXT5Ukn6kGWnkBWf++vgWKAk0IxdcTwgddHmmlwdlYAvAez6foWy
SMgKSrQYxo3EPbuir6R4kNYO9dcveW9Y9ihgagB1HWex2uMtxOMB7ymbAKyYfDwr
BsrOQKe+UDv278LSNK6kdQeTyKCFYM2UJhGWj4IhNzy9I9ESHY88Cd4BcL7UL0iD
gnWpWrlR8aZwDw7VGbqyz98eS+WrCbIixQvLEdNkN4K3wfROiAZzPzpV4OcnC3jB
KM9nk8zePaZkK0LEi4JI/WL3OJFFjDGPnrNJFt5EdwDFawuXiOIuw3xAJ0ZoCmPA
cf4I7Cd0Sg/x/ttUH6Q2pEcIMC9+3oClvhrTQcGkX1A7YjtZUrOVs4u+fbwOM9Lv
7XnJQq6JA1I5dt2sBJ/LTfpttXOM+s1xwbNDDRTZpbrcFqoyuESgzZXEvRiSdHtt
s/sZqGhyVaWw4ks9365QaK/Ooq18TuiLWceC+S1jmPM5VMnBpOHaP311Hv1gWxA7
ySVjkLjWXGJ+F/Rc/BYk4NLB6NLkV6YrMp51hpLU1O+ZSre+HL8UI8hna4Wzw2Ll
OxkpxlTb/lmFlwVxxUUGYmchdSIpZxuuA2EdfZfwfRBfQFzvTkMJ+4LyvsgniZY9
EX3E6f7O11E3uHRHlbl3AjGTHdFXaGOJyWAz8PMebLBmYSxe+WE5bP8Dib797GJV
rOxZIJGHnKzhE5LsLuSJwTTrnfAdmt7G6TGfb+dwZIktx02jPo1O54Giqoek1DFS
yr0csZmqGSTdkW9VjVxyXXzbn43O/NmMejtb64G2253DFM6BddRtKOuzjtJwwsqg
2IMt/DSKU8bxJAx+c/9iia4CAWlgB8vqgxDVEvAT8mnk/0tMEdfaWmNdzMp6Y7jR
Dt2mek2bYsRpw8ZXG87C/r2YYVJXsfSC712w3EStkXQxalO297AMDgDKx6EDkZp8
409A9KXQgU5Pu5K4MeIzn49wOsavzUvxeRyTOEi6j+rECuDYvlpqR7sXSmXwWcrZ
rkl4UgaatHwZznBJYevwY1bs09GjUEBz9GmXm0dJl2OSnsivplhlzy1nV/VT3Ri2
O1Viqh/1jeWezpKIQ8UDtPsKMNNmtotZFRbmTziAdgZJUjsWUkiaCYa8Gm/9djzH
tLXyOcPaZkW4c+3dBsNGA4Cpm0asl9KrAr2wLD97CpZ5jI59w/GlrWaqOJYPt2MV
lw7fulfArD3FZI1LwQKrTZRHpkqHrOki7u94VCCKx7FaSN3wLxq6AYT1kv4tQOAZ
V8dmcmdL6EJ4FN4IhYLJhMN9U4iHi3VhJ56+XYPolISHizL+m8LP1pNk0QWFBPWd
UorzDCxENzZTcr3oBP/eV9GqQse6wRE5vrFB9HTx1+EBAWgi4VMeyJOkjzQdcUJX
ql2txYjAw8H29wMSbHyAH/pksjtkGK3s5Bp6gh2v4ZLjKh+FaNcBxL6T/xUPlpYS
Gqj6IMfAvIZr85gl0GmC9rR0agwWQpd3dhnxJR4CYUWFf9JLBxXXUVhCfYYww3Nq
VyP7z6pAwy6qbbMbnivX136L8qewjfSNszjnxUsQyGU989ZTwr5V6daNP4ny4/VX
84kNSkCXvsjGC0gcGLOyd3gXeiRi3DxzJNUXmkQsmKipS9ikqImnxVZ3rqSa3GdF
svd7bljFloqK8sBahG1MBjxKCM4XqZEa0gor+Py/a5mw+LrZZiGagUpeZ2RC0wqP
S2YZFRtIakumuFHOsLo1nRuppZvaiE1Xbril68B3rb/AVddHGwOKXgzoz4O2vtdr
mBlvQbtdtAw5jvK41g2dTf88+QcRqp9dQJ5QmQ/GZ65ltU5BpeEYDWgAw6lv0nDO
RoDFLC/N9RM2Q88PdX/LiZqz+FleYJ0ns7HOVdOqdIjcvFSsZWasCngpCDBItPab
0305XS0lBI6N5F/+MHH615M29EeNLGSfOmJ3miZjcXQ9H32dpm36snypU0QFYR0S
ZjZw603NcuKzxfjH0Eng6G+cWcLLCRJZc0VL5Ezpe0bZkBLJvWBN1ginikxGN920
2CVcC9D0RXgb/FiIYcycIFxU4QoIhBPo7J5YKVa4qBi3ZQDVQmrPQnoQtrYh76Ki
Zy9jLdkZqdrOGZ2as03+6Yo/t0o82hFP1ISGZ4P/KoeafVFH9jeSC0AKzVvYz2mh
dXwcpD8LrUsPK70+qZPD+z937Vp5t0E7B7k6yR5313uB8paYYr+VZUOnWhmRSmT4
hWHt1F3y2acTiogC2g8aQGRWinaZRahOItUBynxf3YK9L2pk1gDyzQmcXV8NOCSn
QgYkqi3u27cSCYb7gUoVBvsPi57coC00/22jHDQLcgJNrOp1nYMFF0vXCLoZbjkI
hd4eHMKhLJ9RLw3KlMIb3wol+XkPJlWni1WucmT/I8KX4ekdh83V+4Is4ixGMm6D
pp9KXFdeie1dyLaLeFbq5XK/pYFKqiQhtMa6UGYi3BTQxAQPACY+FwVG/8i07vM8
uOKSWCHfDGKc4WwK/MT2GUrj0FvQKHUtwSeQFctfz6RH4kpPMbQMVystzM/+UW62
U6aXgUN5I8LUKrLgQjfyeZEqG/ISCiBj0tuIVZMiksPcGsIRz8Dm2E6tInGGMJJe
+F3Qv3U+qGR9ZahFqkFZ0jpYQsh3rR+y33qqDuqt/8rtvjh9riS3Cz8n6BFoPrH0
VxKq6b0R/2UEWUGPwPIqB7aNJ1M1jEuZVt4XDQGBmf48sBrLNRWypl0w2Sn18Nl3
YhmQL+eW33qRmPhmZ27JQATECV++sSs0O/d6KLajmwD9be8r5gSaEeAPOsvx50r1
M1Ju7917ui/DqrVq3ID3p7txiCKQQ4xW2GReS6eNy/5J89BOBEi/VqQL8p+Jkfs5
E5A3X/2sYInpzgL4JtD0/gsfmozBjiL2nQH3lva4D/BLG05kjggb7N5PSf3dc0P3
fAm+jlEGk594sXq2UcEQD7Q1sjzS6viIa1Ld38X5j+KpiTTSEXGmql9biSdbrvqs
4+HBZ8pr+GMU665YBUtIUc8O2Ya+eBtFzs4xDXuB6sSj5yNiPzEb2meK39yOWb9C
khzFNUvdACuBgeo+ETl/WnGh/I/D6NAAoCjS+dWU/wrkZoEa5on6kcggUzFGYFjW
0La/VdutLn/33/OhvDnpHwDi3ssvb4L61fvIfjUza/H3hKudftK5gfUTfor2MaWC
yIK3rFN4MGPyIPJzvoM9uzE5yeQHG9nHwKFoGfh71K/ldQIvnb2XhuHu6qu65fuN
Ipd1TLCxbI8dath65+lOZaBZCoPxIRUfBUvJVst8YnyYpcaNKeNoHdWGubAqL1z5
9mkmaHng2kMH7k14rQXWwfOpKKhOCfjP+lsNMVHL2uaYQIeqraaHyWOEO+NIhY6o
p70HzeUiQnZMpKssxpMlL0IFykZzrLCHshG3aswjMc1LGmlmAvLlgeUoFsC5sLVK
bqWQkwnocqxNd7zXJQ1hbJxkPeMJ1VzlhbStrFr/sFUL3fIywL+WxVuE1sCaomwx
Sni3wTptS5GZQOtFmXoSD7ORy9C0fRsmk21uXvcMNtSmUEt8yS/3ezKSKBDAvqQ4
xeelZRDpmC7AcH1JVybKxNj6glT5alrvZu/luymw7WIyh5s6eLydQKqGV9auS3N8
mgJct0rqbJcsAdIpI/C2dOBzNfe/r3J4DCbGPIlNKvAmh99gUkwMl5whjrkgdLst
xTzvbut+htmMlLl4Kq59CLp/BctHaND86NaqC/wDsfDBqja+IjM76QrBQVYqhqC/
PN1xcM0msRwA8ZU6RS2eWxa04vW+JqZfrJlhS8nGbPiP+GLzwOCkfZ+fYLhCCIxx
oGNC0oPIsR2axbK0TAH/iC/IGT59mu6kTXf6kFjdmS3WigPCI4m6YHjIsECKDFL+
wiJrEWoeJOBRXYF7ZUiskYAuaJeMO8ow8rEyXsvkTCyCZpeWwMIxGqDhPfDHeI/+
Ok4l5gp9frxUWS+CP70kIa8FufGTDVpDWWaO7ZfbcEURKTkzRYtwbJ8u8kouPePz
i8YY/fb4Maie8heRN0zb7YXbkseOz1iz5+dT01+zMtgq4VcLniois8vbYrY+fgee
42pLtM+2pSylpfgmo2MsnD3n1xkt5K5bqoQzeGxu2XJBULLvFpQMIygKnsEQuWfI
tw3ch4RGjcI/3UMZJKXdhjiwefMIkCQ5KER4e8ECCH/IN7/p6cYnVH0cj4Slalad
Cv70qk0T7XdjOMwK2I4W1HrbN+epakVyy8zhuOefcPe9fPKgTLZyocdCwnIybH25
+vhC1AR7a7yZFwAn7WJ2O88fI0za2gCeUtI0OThD3grkTpPXEZ99e4OGLICxD4XR
aXi59ScrxjvOpc+7ZUrtAGET4PIbG9ZsyLS3jhIrlnR/wqYNVfUInM2gw/avh44U
o5KhDC+Y8hbWiEf/QK9xqhxwnE2DDnH+zrlPDABoMMh3/C5sFv6F4Qpd6N1FTINC
sqj5XhSeiNhpeWRR6cW7z9ja4YXLPx8Xi/qQWWzGWaRXC84AWYfllRZXvJpxR+Jz
m3GNu/Pqc2kGbYNlfgvdsEvBpHUkwZnJ+O1dkycwk8GgOUfSuqFO9TpoIaEpLOSk
FOh8GFCOz5eIe9OcsEmHeq75PkmCcBbHij5uSpC1j8R5x3DJU+hq4BGpm46Y/UhO
HM+TivTnMLRTL5oAGJGxJMvrjCDQznwb76X1Ll1XcxCGgzJTFRqGkT2NAMyvpV0/
S+HLXgYd22j0qI5fi7spCHeSNjMEC8ws1dmk1M1+ec71wRIuHWfltd1elN5mfgVL
boo8QiXWAPoL8EIC6v6fAC4iqZqRlOyNhX3myNzjzS7xlBxymzzyOs+izbYUbi/d
OnzvMXtnEteDVc9Ylm3z+rhPTob3bcDsIKLCGX1yNwSaLdJ4yZRxxllyWR1ehP52
HYzMzffte5uA9zaH5U4dAumsMTZjoyvaZZv0fveu/VSAttJcQHGy9b9YgTsklVVo
esT/2Dddr/Zfins0C+qVRPn0YUEDbaqycOEnspa4tB1YGUrIGfw6uBofhJPiF4pT
3m5tka4X7Z+6Y/5Otm0HQYCwAm+g2EBjt3t3K6fl/IBmh87EWAnXaXKRDeETrevS
+T6fCDX2eaA3S2Wh9oh56UoBBWbkFRLMCZEJs6zwHPdpowmU0rMBAuvHb8ZzAlSC
gjWbkNhe5KymoeMlVqttBmpZgUJmVP4dR8Fmu5FqzOF/aILUOhpEn//ggx+3ZXzZ
8KKkW1qzwsy+572YiTRPz9MSnchzrKm2PGEQHKpNKO2tsY7+OwTQscmAJmwmi5+5
zYiescbILL6H6uzq9ndfzl8+UMqNK6SBjLf0g1x0hCUAdPOkaAWkpMKPvKQH2/Wp
LJt+7jIMahZ8zCNMSVlCcwJ1M+5h0mVdyXEFQUGBnj74LMAl3ayUSysDooU5SudP
7r3vqryDc1YeiMxW+/c6JHo67ZEMuv3NYdRvHqGs4OtlCXUrR+pHsjG6/2pH50v8
Welg3XRNxidB2l7+HESsmuQhHIgqGvUWCSnAeR39+YxQAF3bvxfEeKSy3v+gMGAH
qxB3WCfquT7kp/bd79QN2v15+SPj+GIIJkd79382ubW4TCZQo33rfS8PG9vkhKue
Z4LkW+QTPWLBl+YC6Qp3Pazbq1FXB9XYy/JUssh75kC8puoMYi37i/SeC8ZQZBcQ
pJEfZ6W8yXZ4ZeQVwnCdRbcf+ohK8C22VpBRQCLnGMQx5zfbSEPZvdmG+B4oyDhi
rTUBCR6gdmvLlqISO4L4dZcqiHUcZ3vOObX3lsbYoY8xRjyxxH+O2+05COxM/YVv
u/DtDhYmGfW0HGn6czROERgdCj5xC9janp4Yn7pTdKTOfFY0yts3Ig1E98k+AG64
vgaMGQfW6NQKBeFaEeAU7V2x5MjFE7ip8ioIEUXHDs7Xib2a8bnzIlXMEYQIX3g6
OMFiIcpcMByMvFxnQ1SpiM091IMyS1nUuQjW5n55dHSDZzlvAHMwZFkBEyYsKWwt
lBL+tuqqtQNEim1umE7Juu6PDjCQwQkU3Ow/ov5Qtj+y8sxvjpe+/f0eKZo4PRib
TLnG3WN9yvPJZx8OMhgSGz/463JwNbmaN4EvZ49bWF+t7OncQYK/iqbEg3N6A+h+
+hqM/4dkYE57EUS2/jNJciFD7yEP05SzNIJfsDc2HN8vd63kqwoCs+IF8BBnpdQL
qSA3bH/jlJdbfp+ZkEfv0VVYoVjkne6864e6kAtqKEfXkKtDvxrxwSDR1LaJUNBM
lQ1iG8gUVIUNE2/AbArfqx6bGX6WpmoOSWln4YeQ+vVvYWRdfREfGlBajgTDrQAX
hzDAkplkR5RWajCyeLZf3Jco7OsqZFex4twBmz2flC53e6NCDO7h8sbwKarIFhqm
YcGbjwrKgwkglzJGzGC1QFc+j+ujnh+kgCgne3KJZ2PPSFm94j/FHUXdSsUOX/xh
6AJZa4mLqMKWiz19WggOu3RTJ5D3XE2Ykhrp3z9MwAf/TB9oPVA4YCoADlyPz+WK
NwmJh6vW9dkZqj5cBIb07QnEX29nFh09mJbWckoMkadHFEGCbnyagjZF1+9wtMBn
6MTYTBnBKUMq3QB0bjI+QMJ04mEejHiD5Mg7YcpTYRGEYUmpcK64kASV5CZGDxxs
r4NpL4rsNIaQbN+TSweongasnok7MRfNvcFucWcguEAqTqAytteVg6dd2TYh6Nyq
VDBmUpeARK9XTVXT5d8KYusmxB8+ItUQ1lfojTfeJDkm38h08qHngzgWoqyjl9Jc
6RD60Wo9c/Nk0Cgw3+d4PzRKkc7UG96MgmQoLhnLKrQzn2CobFAQ0IxhCLQrS4d4
F6QG0fiQie18kYzPPOj/PpAaJQv/opf7ZVGckQfMsYT5391K74HPzuNjPvWKWCVm
UCaGDVHTHKKt2kwY+tMW0euz91cN0LjChn4plToO0wEFW0l63XwKEaWjwPU/VjGf
vZ8gkjq0HdGGEeSbHvnMNq5aPDHTzyfimPJ5ULZDSb1A0Y6cYmvMegh76Qn0On9y
2/oi+99kSWI//3QKJMBPPKIgGe+UtHL29v3oYtFrEF2yvzlSSDy3VI+MvBrAEkSL
BBZ4qpne1GCFOQE1uwOPoR/SrAOlFQVYLAx745pFwsOJjJadLMgwSszk8Q0n7fxs
QcgSxnQ5enw6ZsXMEID88J0y0OlaDE4//I5E5D3Kf3DzR8tbr6tHS+XVk1M5xmnA
DrVqFXrPGjkq4gmpjq7agfp+L1qstI/7nFE6nxd6MBRFAZcb5f0RaOj7AjAzE0AA
NFJO7jRqtcMTEXHoFVxDOI2Lz0fdhzMG1wYbLFKdKGSUSA+zraRnBgHUUuMFqvgV
W8Vz92KHI8VXzRggosW3Ot3SCzf/JNplSht+VdFBEk5YXur2de+khr6viyJhII5R
NnnB/stSuyYsrFzluPhPjgrNVkfam1rQgFJw6idAZvKzwybcSJmksbyiU0m8msPk
wYilut7a0IEz/4zmA4gbDPGk8v7J6pyJ/eq/HK4OHX9ZfMZWsaJZCEzlSwz3+0O9
djv+inJZXrt8M4aQ0sWOyqycPAs945KAwyVCBj4DLHYEKaYOkNA6ZaiMX/MbTJr+
uQEd3FzUKp4jzu9Mv/0w1pAHnVTaFqwLqktc3QFm785ecCBCUlBQlBeMlbJ2DxeL
5IH8/fhFkOnnjmum2LenMmwMV/L/B4sJUOLqOLiB6wndP6bOVi32pF6XQ2KXy7rI
8cyRQjEzLO2Vb94si7zsBsDIbhgumtsKs+rWLDxrwMxqCfnL/sdvmZn/FkicSGp8
PPIumvAUtJ7LP41O4ismZs2mDYJ8IZ5u5zuPs4+sibZdNA0VLjh6U8wQIayQAFdg
lDb8zf2dqDMRD3GipnfaSz2kCo52DD1dOGjQIiKM1qcQUWy45zAbCwgiC2W8ByFd
BJsPlOepCfacMaS4Hdq8NcggiUQWR6LAd/tzHqD4zmSKnFSwy5of0af27k9vHxKB
Fw2SUUm9+KWYgdrYvdMXM1U0JBysM599VghnDRTw6wpV4nIjAGytdTyBF4m7AJtv
IccofXC2BeoiCuCLZf63nkIcP7QoI6n5DIKJwxGphjjZqN7CPn1yfVg9NdyLzNLH
gX4l8scfM1sdXYgt70W7QO6Aeis9v21ENa6L6neywf3IXw4lbqh3fUIMfJKkdaFf
P15N3wurP+P7DLixWKNNMAeXsgSS21AN0DJ4cPoORz534ncAD/4FHO7cTYM7KSwT
b+8tdGRGMDxirGJcOkxOSbKlRLIs8mkRHgYHOMUrquwOWJzs5o2l5zYdFh0wUaY9
PThY99MQtcBpJE0z3RvuxBJ9hNs2hAvlEciW9u6pSX+sf7NAmQSePxSRkHmLSsmZ
Z4yM06mleM1m/nYTIfBwztuHTe5WoJdW4L/KYteweVaZAa1K+uPj0OVL+vIlaIZY
HCIq1oDlEZ1o1R8KXChrwifP9ZAG59WJGse635jn5GEbqETZDQPYRA7SLxZ9a2kx
Fn5KsgS2QLvyuArHs5MeAvkGJfmifdSfDjdgn3IYmCaxknF/uHuQ5EBftnOC1pbo
6TDZOmLBOv2VSBj3Xz7EQSuf3qZafKvzMr00zP+7xnZbSw13+vfi0TP4tUevDRR6
9peb+sLIi+JhKjlklVXmT8Zi8RBOvFZlk9kSvP/6MTVF/OsjvlUWLaSg4isVWje2
z8tM4LyVWz9bwwd6iunLUnpxDUuMPGCpnDITGZe4hQ2fxmvEWOugg/6kCBRzVBFX
GOUtyr7C3yg1vrIlvO+fz3GUQKSYuPYPiKi/mOhlDvW35vPSdb6EuyjrwEzo6CUV
koYsqRS91nRY5ztIM1xaZpBjLvpHqXcYLJx+oMQ9p3mvNJ9Bac8ffeJLs4dLXmEZ
cadxNv+a7oY9dqXimvkw3mnsvI2hxD+OPkFDd9ozLMdg9Qd2agMR02RAB9gPqobQ
43AxnJ2yC/ybcQCDUdyDlyaIrS+x/UqAKNi2pHHtx1A6FYjiwp8i9TaP1ZXvC5TH
2XSXzPjFuf/qJSfX+zRTQgiS4xUJok2Z5vG8gPAuAt90aOk43MEGSRyaTW8ryBrs
f6+16Hk+lnGI2lf72iWf1IyulLtWdn8vAABKrgizl3tRZJFuclPLqAMkdFxOVur2
8/1ewikEuqEOBvEZP3OlAC2+IyUqihgYhD0CJq8Hcxv/pPC+mKOYczlyS42CbigZ
zJ9WXRc1ZJRXdnPlTKIpbccZ/8EmLelQyRY9ltzzogJZ4dTh1cpZZEUHzHQ3PEXK
oc7z+rZ4RWsDwp3bjjZq867JAONCZ0TzhAbX2vszu+V3BTViOK+BxlVw1qqmChDe
JqsM7pWCV80sAgk0LbQ/7YrVEkt5+24ftJADcb8qCHa4zd8M5h3olmR+Tw/suLoQ
3Yz3fgV3fpiHuITZalh0dAlN3EYpqcqmThlQrX/n57qwwp1Hjr0S07BFV0gRqaI8
u+iMb+k2jYbI595XSD4FMYUOG/z/8E2MOgrymJ0LABmqWbMPW/rrOZX1l/7mlUrq
x3rBJ0TsQUNygu6BJrAjYl8tC6+uY92kXrfepZrS7OwAn0TwnxC5c4/Ff7F+qvx+
7n9wWM5w74PiUQH8GoSjQnFUkJLASwlCOKTf6mDx66XOMd5I1cslmBdQBeBm8ogA
u9gi8oA5piU3n91UBIxTyYgK/6e5u0qjQ8nABiWLXX5bCOgcXeEchHq33hB18mj7
KLVQbR0vDLXuVHjnBJfxQKX2xa2pzMI5dlKvQ9kPqN89Iu72suYcKGoWMFOR+JrG
G5bnEgbOIZJtu8n5dN/tp2RRqlBY99GxWSpXghtDqqyVxwekiIi+G52FgcF5/gQ9
IXK276WHeP9RKFlZzUIQxgm0jZ6/MFi4kG7VYhFNV1fgyyeLiJvyGY5P82ZjY5J1
9Ty1spn1hr40ccbBeAsxr3cb9YOeHItBrRXpBXSz5suSLJUXnVcuc32KNarrIoqF
iI0N9PWCIB1Ap0ByJcfyQu9C7BFff8juoIT3C9Zs7TRdmEjuDF3U30AXyXNm/47E
uKtsEGxlQsEnXaOB5ZbPUaJ5zI8Q5UzeSreUeUwqZZy/PlA8rtNYmjozWOze/NYJ
yLWzeuc/8xc1hDKdiUr1g7syHzI+97ka9/WYzlq0NCEmIjL5cpPjMPHXp+jEg429
iRmUTPyasKnDnuxn955FF3TE013K2wNYeZClT4uPu8nY08HFNpA+YRLRmilAFVJh
cZv2UX4GFkHcNGYh/EXqlfflXSvpQaZu1wIfY4nDFbMQ6iABSYPSvEl4uDBExj2y
BXZNFsaQIox+TO1nGxlfGMI9qPn75FVk+bT1n8rbdEbipAO8fP9Z+1pp9yaRXa1j
N2UZmODyhs3IMh69gwPlNBmjAaz971h8P7PtSbl7tmjLFRjHihMoDlW1ZdsHgNuU
PqvlZEesZ8D+8KoDjGue+za3fQwcszJwFiRSsgxp8HujmLpSHzs4pj7hF65b7Gnj
1eaOcXh1lttCHcn/iHm0JCw60dSN8e0A+SbTvlqHkzUBb7a2NSrK29JaUyC9p7Ay
8l8Fqvj6eWuU8Ko6C2e0DiJhIFeYzC5GYq9dNHbS/cnjnIEiOHyftmd5YXgcf2K4
P5AM17sIaHQ/Rdu5miWlnYVFuJSE8svLy1TCk1GYHrdfOHf8BTsiV6jfVhr/v7W9
vvgSSCqRTJFGA9t0dRmJjmDqh1KqkhqKSbH2C3kd0JRPVqrnD/dGmRgnACgIErPK
sAzCOS3p1m+YLLFrtvE5ZZxWHQ3PtlDzUxypQQyyoSDmHNFTbnm6BU+iY14st5MW
ulxlFF150UQB6JiXSYUnlpKPMDanSGuf5EpP/bSqBtMWVF/qGDlwidqKqzdSiYsK
xz5iSHIuGPmvNNr98dkZymQn3JqzakpNnyk464yWHzPZSrid7akkoup9Dw2TXuBK
NPUsrkYP7dd/FY2r5Qe+sZr7ves7T8cta09n4BGNBkL8HC44XFT18Qpn475jhiy/
uO9+kLUNsUSQFfgS3DnxieyiMKiyAX+su/z8Ubpa9ptTqEGu9+bn/3LRf2qxcdri
OYaCfSKwgfkm4XCC6zc5iF6YS4Y/LgvXlaUXNizE1EqJg4tncceUM9KNxvG2Keoc
U5Ho43QSgFEMQEjDV6U7UtFi0UQwotVIKZnkzfGigPiQXaKQffqBFW6VvUstOpe8
xIL9nhLlHWx6kRL6DcwkKXsON3bGPtbUSwdUpc/zvXWfnbJWFFZUX/zg2AwKSdVl
084Y4y+e2vrqfgcuvU7gszcx+RdqClAjikrKcOs/Ge+64thfozXPXPQI97xeYnIf
NN0D3ZCLT96a5PCN309m6PFnBXzfzxu3ZF5UzVmlayHdwWMfEIFCmhKVdsi8t8XL
PqM5Zdnt0zIbm9iqjXi8Ks1Ww4xUijER4bpcod2krBPwMstDGEB1vjhSyrd6L8PN
nBhb9/gZsL1Ywe6iU3RIodQnpFsV/PY23/Uu/94nLHdRlfKQhxxuJyVcgjq+OO5i
gtvvlqSjEUo1OsY3kwckXLghHxrFHQ9rXHzYrI4OVc3KEBOeuTz5i8BWxcwEpWqL
eHXaPt1zTDWpwfB1DOCQ1SeL8kscus61RyUH5Wz7mf25UoWrFI9Ins0uBBOVoKOR
GxHkZ+NF5Q55la0BaZOB5K2NTbBoHsZreIJZcIXRy937nRs+1XbRwUugNZFH9EcO
Vkv3/Bp0TdftuHq5jomnPdHVHzDFZYoNmYtVhYwDmPNqdSgXvEx0Te7vLRAE1cVR
Z4Cq/8ron//cB5P8x9xNRZZjKTr30wiispnE8VR5CWV7HbjIdqwH9r7HlOQ9AM9N
SIfZ8vPTNlQmLSX197cfQXEd1PL93KzU07RWI/yCEQA3D5X4ca9YiQ7I0oPQk4vh
px9XypBEpK7vrTH25ggOWyu8535c0ygRISzZydPN0i5rUHc8LfmPar+Rdn+95u6a
l604x5k4uxvjb2e97piRO8n91VI2Cd4C4ot0geWJIK2Zz4f2OLHbNZY0djRolBur
DHDvEc0JcZ5XICgV+u2XWESolrvVUzMWIViat0Qs/yXDs6Amkp20LkEoQLdOxKhu
1u+H7toF3bXtTYPf5hq8K09CfQRCmR9MSpJiOlOBNJUZoe0puL6yb1teFMiFO/7V
4i59+4KlWkGvKQ0AB/XDu4y5QCDkHOnvp5TJKadz45hYkOnHQybTGdxliPtVasSW
BU7aLJdcBKY+5X2SGZIyXdEpzqqZqrHVMzO8Z8HS9RdaUL4uIlMg6IZhYc5Pm7xp
S4lvkElZUvnCd92pqVtLso1E/WE328ODADKTSsvzuWNWpBjR5FuD7USy/0neS3IH
c4J1Ql3dvFUGyJVobD5QIO++/XQb4x0C4w3LJH5uoy69SvvARRrNzAJmEbpuZVXT
8H9w3q4/G79ht4yUTxfGHiDqxKIk8dekIR8zZ3BZwr7fyaaDV5oBaSH7FVWGNX3W
xbQ0pNPAr5AIK/5MjE4fpPA9EsVK4I8vXS1iFaq5mBBiu1JqP/pzsRd3P/4mnP9K
wi+nWRIIzgNRt+9qbeXDMFVWX0W98rZTD09bGluF6n5ghopdzFKzMJa+A38Bfmzd
o4q9owY4LGCQUoWitlvRZ1WE+qbAAmGfBnaEDCzQBeX28a7CPl+ZtjJSFIXY6zRZ
rrvXxSDljwhWuc4XyXPFZr9Ja2qSRSx7NrpZ0VDv/G7DSrqnwv6BsSS2gsT/HPAP
cTIdlq6nZquW5zJG3eivakdSbiOZPTnciJBFk5l3825V3dU6WFrSA6YF6CN/1LoI
2bjxltKcZMUkmfIvyNPmlatCK370NyOEl/Le9YxQi35cUAvXK4Fx0MQ8Z7bzzWKu
3NFa3ce0C10yw5VSCFimMp5pRqO5BnZig3UT8+QN2H+Zhys4rv4AEUnWPHb3Ud3Z
VpS9mXk9KAuFm/gN/fwo8LRNpaNEOHhswAdwpmoehRAAuSh0MqcJI2Wj0klPl6Bk
RmKK2Rouk3hnqFeWak42oXonn+0p3Y8wCyHKBix5Kc/1Wk1iBzllQ2bVFbMAOTdL
2NG30go15LAMuZvTzRt11nCdmfe1J/3iwkRiOopIUoI2iWV21Y9so27m9DLmhoMJ
AUmTs6zrO8manpr8E6OrfTyQDHg8Sw/9ECXqjM7YhwuSyupFIaaWqia4fc9G5lDh
EN0rXrsioRztkfd+73Jeg0OvD7X0yy/KXdW7oRTWtnahAbLnWK+aLeO3SRwniFLT
4lbcHN7hYDbyJ4a26uzf+odnbTYGGE/wMcyYEXhG75qc1h1TiYWZ/kBaXQm75slk
6Jl9Cpl23X7wX9Gb/P6U4tc1h0Vb10bhfqFdRRPRjXAKQ6RC7ejxy6bsDqm06ULG
cy8093ZF0I8GYM/CposfcB7N4b6A98AQ1wZYacbto2oaUFg+xDGAj1fp+PXMlJIn
0in+ESAuQajFq9hJQWDEdAXtUS43bbX+R3vVC2M8ZX0ZNDXy+u4IHHdbDT/RJCE1
Lt7hDOm5ym/2ZRAAcswadclDnAduP+md8MgU4fKHAFK8PL2wZTchLoJTBcYncb71
OSGEsdDOUkDr5wVsYhdBNxXsAC2JYaTjpmD/GIFpF2rzgrKDkqXHuV07KN0yPlVt
yqnx6iBnnHhGwqXT7p2mjvzt8RGwH2LN6/Y4XSgynhi1tjTjX7f5DJLjtaQZlDw8
+PzWSDFDoI7sXPwZHP6JJ0eqTXarR3u5HfEa7SrjukXPeeODz6/EEhDOLBXU9Sne
jOMRpXuHx/JBhv+jagmzT3kCLk5x6gGv8IIswxxh3V+u4IUamtXmG0EnjClp9LgT
9FfBrfGocp3+Ip718O4GVOdRZ5JW30QpWZaNl4wcf4zZv9oGdMbcfTVmyjqYK3jT
/jUQcHKxkZYb6JwmQqEExckG4lI+Y3GH1XITdTWAfj2h7VjnPUgz4AZ9CRve9PnN
MON3iT8ISmjDUFOU6OlNcDPy46/yKbcIf6ZIq+bwCTxkOGIKLzhuukcHO0I8wlZp
GmSzIuOtGx5tmDMGpPHGVp+U/8nJTNWXE48J9ZWEmT1fhA1tMPlxGTTtm+YJvfBJ
6/Fss4qyIlcmoClrBPIQ3usoAEK9KWhplmNAiKabJLiX20js+ljl5kt4dJAcr6Wv
xDEFkXbdQPA2NX/sxpICFev0xBJkJjkX4gKsV712Yyhb6wxyX4zpEnnmpK3Wd9xb
C8qcMuBsBQ9ypI5NPx2M3e3PFqZqU/AwOGXECryRmUGv9vl93qf0C0g4Uhu1Z9f1
kZ4ImcIMYCoXBVyEqgsoXvTba7tjnGqPbgQQC6QTXWC4e1+P4IRRHtAT94Efbx8b
5XZE+h5rnO8GSk6fBGWBKDjr3t7nfcWngyAUiFExITrLFiPgD8LwfBkamvC/T+84
Ljia9/43czX4FAxDoCGUVX3fNOvcPMoZOgZNU1S1+oDm8WFAoNXGTbl6/lDiBC34
Jd9MOc1iCTGepGqYbpt6hjS7gpbUSwX0DCKgQJ2UOgL8912QAdBFSUW2n347RqPj
k4nRsFH7XoIdEO+dwDrNTfJpiGF0/FLMogXcL02zHo80aZAO4zkf2JRfZ2sGxtzb
0BfGZA27q/A6678JK1YJUzhSYgA/Mff832ZrR36rlFiGwxSQk6bdwjCjWbcb7Npz
wRfScn2YCQOh6mCrPKJCf1ncgg9TWXb6V+1P/S1UtIZQ28fG1QdjJIROQi74ZIgx
hvD5XqTvCAihMeQfUKtR6IAE6RK2m+s4WrSVX3OICFmmi3e7MoT30dWBmFAuLBY2
V2KOvNTUfZT3B4GSzmQOxXzfvLhYPA3m9cRrFx2QxsHcBLRRbT7mBMbhG2pqBG8o
YGsgq0/pmWjBpq+nrYocQpswGhr7NlVjdWxpw4om5hdrgi9TN4QulTQOJUiSpY6Q
U6x6lXqsD8saOZd9d4Vd/o/Dkf112QK3TUF0jyXf76Ywz/i1p62Ij8c1cPjd/rev
FopbSuBcgvG2P9SZywlUcomdILdXl+KHnm22bncIYDnAQ2WzErC5Q0i4n8L6Jg0u
DoDM1WhLMWMw0sk9ulhjg2LsGdmPVTOznS1tDjRcgZJ4oB5KyzrQmOQ7quBy/CiB
G8vZGByaaN/WaAMYQHNLdMg3KbTfwieiY85g3MlaOdCFODA5c3Vz+KI93rdwWGAz
4OVm0aCidshp5HyFRdSCpC6YtfrE9emKZjUPbyMU4SEYvwI0fQUwbLkE1Ps37Y8H
iiZpyPGu5FdluDNHR0KLL3ZtQzzfjL+UzNo2faPBqEmJGW6HcQT08sxvAO3XE1fL
YurDQSO6pktLNx8iNjZpg6/6HMjxxsjBHwHVj1oGedIBDz1bh2XnRl+jsOt11RZ3
/jy96jKTcNEn/Ue7WATlc7CT0bMXi1oZzA/nRV2ei2I2TOa7z6TgyhA/Or0FcXRO
24HGU6pc18MfeCo2oUNfYTyk/2hntHelLeDatLct8zw9wqOE8wZsBirn/NGgFPxv
ENDFFBFtR+qBUXXhjQIVTT9rNEQdVn7203pzLN2ffXmEYdyaFDT8/JCDBzY7bHz4
Tuyuhy0TJdyw8f9QqSicH8pSG+sKa9z6ineaBndIpKtHEond2nCe1mbkzYQsW6yj
xFpxgkvlYcDaDXOcB7xLNb/aqb/4/+OWaVFoUrAhyTEehThAsJBipzJ9CGIrc7Bi
Ymb94Z7pB7cFks/8k+Jcl0RlqWs6MiQopzaO7AFyD+ZwfOKhgIp+tprztgzq7M2d
Sf78gepW1rKkHMT0+3vmOZQdoPkm/DF74H+f1HdeeLYgU13a2k7/4UGLyoYAuNqK
dA0LI/q27dxT0ZJkbCfIpKR+MIqEWZEW525iGTTwXK/makeEeMCJSTWKFLS14Ys2
tREE8Snbu8Wx1dgsZpDV+NWGE68X2TEXy/qDEuYlad6a/Fif6rFocmKbTznAAwvp
i7zbclvB0yPu8MJ4CR2Wux/4t94DScM7rmr5bhVowafJKdJLeS7KU1tBMNkCRNhn
Gfmr9xFDvuTnhSmnai2QZmDoMTxnvYUTxNOeaSYch/akM6IBuG9rrldj47ETWkeS
kJEKIbOACPkFTq922omuJDV+MSW7aUaxZHItynqsL/YzDtsAFUxSOKQ9FioH/xUu
d65DH9tjzhmdTRt3vlg6GBsZsnFzfAaW1pEHJUbTeG/daKAriGh+45X7vBk02hTr
pV5Jy/8lpISFXpRxh7qfeOduWcpDg0+0dNTemNRJwSpAPMTJW64l9xtQ5EIT6SQY
h8i5J/cNOyytfY10P60E8aqef2zDKB36SKb4UYmow229KikkeQYLIvv7/XiYyjcQ
R9PJuAONyHPdN309Pprhybjh5qcO/1qrI41qev9bKw1TygqnD/3gbwTvkOmNY9pj
IVBA3ZFz65vgJ4MeYwu6hwy6dYtUpLofuysdOspUCdfuhk+vrrm3Am4tbkI8iruS
sflEWGdNHbKommhGjPQ1IUg1pruGWubQ7+qEXwOMeOvsodU8hKJbuZW131sz/IKC
EBRZ/165YuXD3nAJR9MMBZG60ynuNi6M71s9uQJW58pyFG+LPfa+7ZuETtJVncZr
UmW1zNu8p++86cvCffIb8TbbJUA2OpWCxBHV5U8isqq90RLrPuhnbIrWcQCq653M
r0MW7qrOuMXZdQ5Z4RTecRGXoo6aq9MLlHHF9HWFoLV1Z9Bq3aSn3fWLTEyzgn+p
RUoSJWebZVudtevAqLPZgiseHn17lHnM52FZpa8yn/ZP3c8v+s9gRLedVrAGz6RJ
o6BJX6DMb4kCGJJCfmKCkkkYMKoGFMp/T7kzg1zITvT6s02fsykpEWxsq1hhpTBD
9g4JCeOAK/v9qDYQbCa2VkWyp2fN+shNXeamt6scLNJCG/Rh3Y/s0xBClwNo5MwW
O0U1U/UgFeiTKURLJMSQplgVkeTXLIu7+QZCjse0TA22yBMD9vCkk946WFYKscVk
aLojJ+aZSHbtCa98ucekFAiOjgWCaLaoRO8SmJh0kNKwLUGecAHPRh8sQKYWA/CZ
jxX2XnZiB/FDZ9ofjlYEztFONCGL+IIw900+EhFWkZPTKbzCOqt9xp8d9XT4SG3Z
QbEQlkkU0dQoA766LPwiToHsEDaiuSQdFrO9rnIB6dY2uwJcX+M2DusIpHTODGwU
7GEKxhl5y803hLXnecx8xIzcJrJ1xDJ4RQjxzPHVIYdlA3GhNxLD24Esj7+qjMpj
NAjKoEdX+dl67bZkWQOLZgyK/Bp/Vc58MxbH5CQ398RtXI54+159r4scH8dcyejM
emLk8FHzrJXvCLgbbK6c+K2TJPdZAiBOT5yWclQS04q67EwtSIA62SAnVzxDMj4J
zPgSnijNxmpM0aSXsISdUTRyqqH+Gla3wXrnaDkkyWCOkwUD4yvI060b7Eo+Q7JC
miSv45ka+1OegBLiGqvbMCVf9mR/0BncOg0u874E0uvBuJWsTfAqoJNwwadVyFdt
UIROfreqNPymDJojXBza/Dn3gdeqlhOcExJ5Van0Yh3f/hHmtROXncWLDiLoxedU
XbYm/p/k4SI3zeAkfQyLoIK7zPWB+OfSXe/xAht5UvI8PlGAYJ8NAkPnk65QT6HU
drhbB4cdBKY+9LgnVUwzjSmOD4fpUl8pcMxXzbRR8KJzEzoSeIFXsX6WulKgJLaJ
8kr02wKQWW+HyBkMqyX2VU/qeqKcExPJMUEPm2ZVF7u9rNpBITRUD4hHVvueUEaR
jKdnpgNz1Fllm5i05LCLe5ZF8VkYo25i5Gf5RALiX95iK2ewZsSnkfttZmMbmhit
xKv9kGGw3B0VIW6bDGuTT58VTTWKS2ZRUTJ6Q2ywjcUh0yDD0NXcBcThIY27OO3X
ScnL9hRkAQvaPPYGAPWizpOEZsb0iZPp89O2Q2mY010V/6JuyTU1KEb8i+gqEwjK
pk8JlhjMnzLKIztyEINRCV5WGxCZF75vzKidspBj6GmKQaeOutQ7eezLxzCu/BWd
lzy2lY2g14uR8msaXjcylVkVtNJVrC6DDEyyuTYc3ShuHyAjMkOde4GhozgR96MS
oDR7VNdZAH+CtzmFmZI3EyLlGv/0BZ6LPFSr6azHlmE2OEcWSblvbr7jNqjePYDN
UP9fWWWLr4Fgfl8eUQqhbtseI0A99aSC8d15f9VSJNHqmVsUk3/5+hB9pmIGMvn7
np205fEMrt1QcPjWpOGzy6cFh/Bmkr5se7hkqfRzZHfXa6TQ6jxZEJRGqW0uM/A0
1NT8RqLPyVFCGAK9qdtcg5OP/yjZR+qPkmOPFEcO6UbXF4U3x4ziEhYjc3bBbwG1
oEudhfeFLOlKnk7gjBJaseagxEjuAvM3dJAbAdckzufBR2VYP0oIG5gKLYMn2mjd
jHhub8L3+Vp2tSxfAfWszKmg87HziatbqsobKcf/w3Trp/6yQ+1F0SCcxI66xKgC
OtSLUV5ILba9bcdtUWx1D+ex2W2VKHnYtTAYgRgJdZBNX8e7M8b/PunO8oygWf1r
Gelwi0mDYoktGbcCOOiDMI7HNn9QKxSTsrtG7ifw2mROED2oZNdONmi7kw3mj48r
IwB2/+9J2wZrEVEIbfMO759QBkDpjQcBM8TKxtEmuF/lVz8hSnHo4F5dprRAwxoU
AUnBFWAKfPNBpUUFjx9q1BXqf1L7CTWRVJlb+5Vj7AXMieJibAAFWFh1145WbTqj
XspSVHzHGuKL37xuPHxXZHRed4wH++ADDdbwM3vRu9rXb/vbl0v/iiiBFL4kg6Xl
tkheYpJDvj756OKoL7vi88jEazwO38e/IGyK90C7pKxS0oDwpKJHjfggF52/Ve2Q
+pDFe6j/jEETdYBgiMGHkcFX6euDSex3+Hu25aGwPYXeFb1kA7kR0+MkZK9XfmHp
GnZwZ62NZjymCw92QA+H7//YKlSBZhWIQy6PJn37I1hS0IH/uY0czDyMVxXA2Vi3
VKKO1ZPr6HDOvX8OQrDZcpR3+dwydUG9AoNtgNX/yX7Xa/RMHcNStcWbAnYqCLpM
cDZhaBjVaKuQ35jjZ/mDaaNdtPzaFx3i1BUzpHo1R2a4EkMjaeWwKK8dA9dulAEK
6hib2t+KfgyVAuW61oMDHFctYXe+d57dt9ppsVmSTXYZTdpfiagzFbFFv1uXzrnm
VCfekFNEd3HVMiA4HwgwbdFTQOBhXNYxlxZTEgeVfr7ohCWhXKdJFdZnwgtxob+N
2rsglkDj60y878bj1QlPjiQZUwUTrqvXnyPN00LzejN3afFA1fcyY0fS8SdGjOHv
l4u1QoXgHR/ixabyyZfMr8nbaxs1HAfIC7CHktA9ke0WkSj7m2yTWgRBjI84nmy8
jAEqhwYk0lCcxWRi9o9BCg==
`protect END_PROTECTED
