`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wh0Fi6pt4P5HbNcON1jI1Yy0meCvl4ImnxYO2NU0Fk8h/RnjxDqdSufOO5t6uMdm
Z900f2d25BpehjWtqUQBL3Jy1zYSoL+fwZ/A6SWzptWI2JKWWY0bkEfbvK9Nb9pp
q/Jz4mL7qlzKZIG65uJIgCM2Jni572Fu+RutlJhKayLd7Os/3KdiSUZZ2A34Ee2F
ppa3juOXxWe/XcD4LQVer4F0OM6YqTKc1+95QOeiCk3s2Bmtnh8RhZO3Zj1yWnIt
6MUF/G82mNbkdac2PjEUEFMcBeTXIH7zCEp3p8JoAc9pGgNJcQcrJyIL74ezCn8T
TPSw1cc+35+tmxpJ8jK6UcztQ+g6D4GmDArwq9FkXCtpKoLo04MA32IQ4+9fm/Rc
9MPmYUVPE8SHEySpDVLzCUEP1CGVExxP2umUBqFe78mKhtealp4OkycOriImx6UO
U+hRpnM+pq3ZWrR2fax3vNksfDJ22LR/220Mzh3tqcMAmjY+UAXYP+hV8gV8vkMR
FEW6VYSTycWUiu0ajgcLkXZqsnP2KfDCSjJnPFydzeL2dekv3hkkSshutnRFa4Dn
lAn4SPs4a6GFcRwwTE23GbB4omJqKtZkvYJCJyQGXmH+a/EUysfmZxb4iPdiim7S
ZOfu+TVSlRynTXwGIiTs0oZpR67LYtEUOW7ERYAADzI=
`protect END_PROTECTED
