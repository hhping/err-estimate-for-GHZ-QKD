`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0UGN7ZvMPFapWsyIOPJ27+EjBl4y5bis47kzg8Efth9etSLFKypMKBbf6DTOTG5o
PIGVjpm1t78regJrPwPvXUiVijKvey6OAOVFarHvm3hjk6TK2/6yZWlviZUxAwiE
RXXRiQw04ln8MorNO9MqlcHOZI0VndUxwmxXTDKOHr34hZ9WsZqVZhL4TH7wpTyv
4yElyvBQRM6Vvd1udD4SGSDtfzInTydbSln0ReQesFalAl9vb+5JT1ZX+lTKFiCK
s0baSvJkr1yStcaODAVILFu2pPU/rvx6jc/J2WOHRqKkiK7Zn3Y8Uh0smzzfGEOk
hM/dKisXeZeB670+6K5EKdj2ftytcivw9XX5EpL7WJ8FOf9YfZ5y/ob+TMZyl1hN
5c/deZE5idTk0yWZ9mcbAw+4rp9NKhUyAcpxlLgZ7o+hJvOTfVlGyddivmpQqeMF
aQ3HemTSOagjHcTyrirxL5sQ0sfexPYYhCNdyu+fXa38uEYJz/etH6aV+Xsq+hX6
H4wZZP1NbvjYNNo3WezhSd/NiatSSnoDXEfp6Y1Lb0X9QuMNtzdqNISdql08iF33
kVyW4ohLRQmbNIsodkERKeDaimDTSLte1JdENm1nImmP2+6AVG9fyCAeznGcOVqg
SVXGQXbi3wQmaJZw3AMCIxmhpGxcJygsxNR3JvZgiCVI60E6Uw7d1RIQqzF37HTc
u47gwXZY2StVNKLLwNO1elELsgsfSxAxjAIJ846Wdq72+y1cu68ZZxajjc8doThN
BzEYwT02onlG0Klck3HO5z+pKGgsBgMdKh3aiKZTqFVMNhFnNVJISBduxVaFRJOk
n5O3Mhfw+lJPq/tF8+xaNFI5dsaiQ8JQ6YqyNWvagDl8kGrJQcF/BKT4xq3+QWxn
xdVTogsuDeBdFuMpbL/MwPtgAWITwBQMnv5wi2uszGssJrJI2IUALSuGx01ANEx5
gQX987CfO3WNQ7z9VjQOerSsXRXZmT/zDS2FX69JQ47+BZ3hdBQDXakbtCKab9Iu
JPSmJf+5dG00+lLpmWCLVhS8Ixzrb9/D32LSg/KjT4RCaur8L9t5rMmhlnJLCIZF
qMM7ASeo4U+rIOuJg+J+bbUHDrya70kiap59cBwEb8aQY9/Y1uFFBU6KDyEUIjzb
ePwEL62G47NaAvFPKZd+Z3EnymuXK4ORRInhs0y7qAPjjtn+B5tA/1Fd/aiAEDvP
+p7r/W8Tk9qzU9M1Nc0KnH868+5x1jZQXMlq+G7pIvw=
`protect END_PROTECTED
