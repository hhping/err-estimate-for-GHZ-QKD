`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kKnCHyLsgybs7Cx+im0bpCIaKFrozfNSOIB+kwDzAZQ0nNqnNeBgjYVaQPSzWQXz
fWCIWfiJqyDpfu/NGid5iXGOsjVLxoI7gs9nqORojsMvyjIYTBUTGBl7Gxxy95ds
IV+nGvdv7sWwohFoP6GQ3jFg/+QQcf0i6ITTtr/vXOSS8qifOkxpO+UmAdiKk1CI
GUqmJFGw7Plk90Zovo4VyMEcIekqfRCnsS6AYZ5NYk1ymyLWaXURcNxd3SPxVN5E
6DlqQiJnqKQ6Xp8cBRbrk0BDKILfIq4kZH6Q49OdvbBmZGU80gTEOQTJefe6OlGC
KF8j0onyPX7OZfW9YJ00OifKdF44xhwIGjZB3K8lNC5JpNhlWyFct7kJsnNFICZy
B4hGf6xDj00GosOiiVWrazdmr2dMUzBrKBgujl5QwnvSHE2CkM2Pj4Woq8vBRuoq
C+q4FttTnvJzNF4ZV/W0OIpQH4+FubRrDpGHuh8yBcIvHlce+79Zyl9+qt2x7r7y
sowbiA5N25GRKiuONhBlAapfnSFZkWlXrP9487TWAix3/aWBzk7PBrdaLJDF3zpe
x0VcwXyR76ccMt/89KJywvtQNH2C41vlRECw6u4GOcVB/QFej4ihUsiwZcQ3HSr0
KfLNG5PSSt2ndcQMoB8c2gaGlduWan0ABoRcmZPy8pc4iVsA0IfsQD3kanCOu54R
4/hq/A7fMHvctZ3md7mLJ7/6eBWBXTOTqbCP6xzuVid7NEY83tH0/vl9X5WsycQv
aEjSGQ+6X9Z5CgCOk1HSvxUA3S95Y88Xn9KBPeXNYP5c9rpTlj3OSmNLAJypW6Qq
8AasjoRFcUQpP4qAv+rPs7cL+FaZAgBMpiiwmGXb9vsZyEr3MkCcXK+tE78bdNDC
4fdE4eXer+catB2/EMHX9f001VJv8oMQA5lYtcCII8gbB5WMGicSQiVkr636rN8E
Gqyuzfyr3pH1sVeI2f/3MRtCnobTV6YVJrIFWGseCRhjFcppc9+lo8HN7AWNxt2V
LJ8TDVsrwnAlKwbkjJ9pcu3LgTFZbRwKNIiQTop52o5rsdeBFh8zSDMrYtk0wTfQ
2vWrfhqJj9d1uCstkk21g38JumuqRcuFvoWsXPMXyNpL6nQoUK0MAA4KARVeFokS
iz0DtBKMT6TQ0m24de3mTFnW4dao24LDRjLQKxv9Z7/4v/U+eLNDBMU9QzAgNd38
JRe45GRfiW088R9B9IKG7ppW3rM0jZaJ5ztV+IqYdirfAF3TL2iP1TKuY/KrVVhF
YGEmBekElZRrQz6bk9p3qqqws26nEJourQ8pDhvsox3JaAIhQYoo+0DDcjQiCXrW
i8ygCeeWKJ3051GoUQxgjuRaxJLVdIjrwjKZFzfIFzso0ICfrgqFuHy1y5BHIVzW
`protect END_PROTECTED
