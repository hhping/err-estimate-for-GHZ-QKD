`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ECQMeonMzEXcJOBaQmajV+tcTHVipGoI6RsULcJJvtAcTACwt0RG3usNjMmGNaS2
tquX8dwnd1N7JMObunHWrxl43yfNKA944QwSrCpFEvdyJUHDBrk9MHlTpeJ+1BoV
Hn81518aazpqG6duNoclYzs6D8t38+fz6IlF1j4nsij6Pp1rgd7SHI6D7BX1bwdD
Oxh4I6nIQGUjwd9gnEFr2F+/RNTi3pgjF3RYIKlNsjefQpBCqRlaIPmGGwmHTIDx
`protect END_PROTECTED
