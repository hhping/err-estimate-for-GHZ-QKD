`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qh58T6mNR+VstA13k7j0jSdgQYohfXK3x4QUWCVyPjaoFH47ZIT8cTyX9eT5UcEH
9zRILGDbYY0zG7oK7QRL8OltbEXSk23UiN97hAyG/IoBeNrskcTVk+OgKceioX1V
XKebfDPryUgyceoe+mz5vTk/5Tk6PF38DyeEFT3pZPIXydB4CmZmk5jy0Tn7Oxe3
aleKWJ/DeDIaICWVXNqmrM/U7s0fdteeW/3c6vCQGxfoAqpZXBlJxP+JfUWg44H2
hWwh2F2HL1rvch6+F70c2gPKaytqWz6q99H1B1h/U8sRTKgTG3hpV1iK4hodgyqS
dXqfwvZVGIiHjza3coGS1eZQZh0vIXTRQYXJ+exiLBc351d0OLmm5FwTstMUrtqf
7jsZvnPVWz0z+9UbTdzanh3XULK996r7N1Sx1rDqsRK6mY3uE50/WGV8Oz4Ole1V
wV9D5U8vqn3yLzSeUTSyFr2TZBc4S1zoLF1l8HnljR3lH46WDcLbxTJaa0bPMiQY
51PGVtsCTw1XKSMdtn/h6Mv2FQlOcL37E6Kann5dE3KrNSw4s7tWhQnF3q7sGc76
Ebk8XG4FcYY2pdiCyaLeU8RWhVkH2cCqb5FiuuA5R7I8GuziGfx6yeZEKHJhBakC
81XvXfO4X8ssef3sj9iaRQ==
`protect END_PROTECTED
