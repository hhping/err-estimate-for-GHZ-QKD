`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xXsEttoYH132NOW9P/4jD+yF/7bNdtBJCJd8PzY4RZTyP6TmtphBQOrjKvisQuKg
/8Ma6y8cjDCN7DjhwlFwLBN/sIy660AKGrdmjTgNngqPsS0TmY3fFwHmvL/uuH9L
PdhPQCSkiZD1ofLUuPKjoLsBM5mnQmP1Xjx9o23X6IodK3ZZtZOYm9a6pk0k8PM+
9nYPA2Agxg+D4LZRFkf18lzR14blmBE2e1a+a3ZDdjmDevrPvWZI7voRuNs11kL0
MOx9UE3hxmI+qCQhRp9e67l9KvWqUsh8WLcU0Evthrsh1mFQNtwwNQI5IOTvlHay
Gb2boevoZdULFzlkUWT9H+IcJdtbN3Nyo+azURXg7Lg1QefwJSG1KXdy+TXLS0Ch
6IkSTRtpc49vwXytA4kPYl0nN+Ie6zmTYln8xA5VCK0QW6buTsMwYeaGeGdPWHMG
vXwvpN314Rves3ypSRGW4Hys0C5xzJXnlmDinO5tVICzSdCkMuT4fzCh2V3p0xSA
TIMt8MhgKTJaIRaePyhmMibXUrfu0Z+ET5j1M6a5TMldfcV3wx02YJpD82HV/48y
P7KtYcCAguut+KQiroZWhn0gLt6+LAlhw+f6G4dhdGt+tMHN3fGIdlN2q+uo0N6F
soZod1nj4r/OtFFFz3W7Nmy2nupKMTW8rNTQUtK/eseK8Sw71w5w6yiiHxer+ltr
QF4yyMI7JWEPHlcmSAQwSbXsA3WgDcMgyNO3N0XSN46/qyqhvG4+5TMyb0KjR2Sp
+Ou4Ji8gZVYlXtFrlODudIyPVUzb9ryCZE62lVvb1wfgkLspPb15bNcKK3RAVKOK
qrCnPv1WWSLRZdEFNjmk75ZR4X8gR3xo3NpgzClCAIAHUIKDqmbEQTo3OSj+F468
Vb+B7CAI8fnZiHOd2zlJAoir/OVwlH7QLjEzehR4vZpWujLo3qa/pYrIhNPDMxke
QW69hqP8PMkaUdfpdkGEVzz4PiORBbxv1AwkfNS/WwwzGUdeP9FqGAxGSSYQEvYD
eLNUoMSE22TrpR8pIjTw1AK4sNkPtuQ3qI64M6DjuEO+5D9CbZN8WR32//3X3ctf
hxGET7c4TnxQQM1N4/UxssWVAJhC9xAErbkR4vMTctWG0ZewHnf8WVq+fAiYibfP
gOsqphk9wcL6By24QHLiaEQO5xKhRpGV0KkSE4h06WFSyDop8QWsBeuuuQHf14PO
A7bGeLvfTQplRxVWGg0QZR97vNAuh1PFaRC0wyqGpYAhnood8l+EGsU8BEA6z9Hk
jBmqrjjoWmdSVnJoks4E2wzGDpYcvivPjEDcAM/OWfxTuVgcd3mBQAOoymfWSI04
dgcZWhMIW30TPhu7r4Sd0SUEd+8masvjJRT4el3ln+Tbfv2xHd+2boHr0T557CK3
mtni3gLO7KYk/j9hL/6BdPUJoIbdL9AEPegySefZqJK9Txz/SIiTN527RQCkPBPe
nqLJT4/yky6fXAPo7TCvs9qJFmL/HcmEHzYH0Fyr/X8nb+jW9JFt6VR1eqXJ4nQa
cCpszBq80pgqGRzS/IBOwkOEzygA0FHuhlckQQsJjxZS/S2furUA1pXwuf3K8wss
DTYDCrnAh7fdLFUr+qIbC03sM7PRhrF4SLNLKhTtP0iPZIqwgl9GUGQHpuw//nME
N7nOM0FSLotmRvDxsF+gUX/DDBCkeMidhA82kJ54ul1yc+RsMxepE0lWfO9jNP83
B2xebu5Eg2z8j/NsxLkpLgGxqP3CD7VWoL/R3Si1G+RpiGfIwWFuUcsvMZ0O0nLU
+ggo1dIf5/GwYOQf5id+9AQNBKAQYhrNnDXJBEFEVwvvbCrbG96StlLi7zcXDGxY
2ybNQIK6Esv1AxErbnXH4sbQQvJ1tpyBnauPcnSq1I3hT8gX1Z43SJgX04JrCrmd
u37MoTbi+9iEwJJrHI/2WuFgVP3nf+v9z3lpkvA6Bce35F93+39mrw0qcDOTVXhn
VYL6V8tm/scVyzEdXVye3AtmqJy3qddjUSnN1wYxqIchclhNJADzzo/vbBaergM1
lRznX32qmYOZ+ynjymRIbZ5q69I8133GKn6y1K+VL6U4maGgNyKN1j38CMSPHqHC
VhFOjDTwf0RSVyYug8JnHQ+MLwO1+qhPcp6vsH9RSoiWZDvhASPhWZntjhwH7xlx
H+XL7PV7fALXX3k1k0HBKYg+ulZtyGFwhLN6KkWeRJCb5hHv9q/aiOOyxKcLQsd0
2DD690DTyR2bdECK7yy7w1bsd19KMZJpdoRErsVd5iS61PgzUpG3GICi6iGo2zRf
`protect END_PROTECTED
