`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kIaYXIjT6EJMycHHvGKlOoGgAEIodjbQMWyTOukW9CQtUfci5qa2aVTiGBq7C8Y+
LZzHVp09/0NBlvzpmVFcaRwiGHpDreLgewUdE6nmVXeW5q2do/eRlB4NBI5lVw9V
9fG/FlYAsZJooZGlS41OK+YkUZj4KfRJam8hCjCTcU581U6XGgZB6oGan803vZD2
0Z6sj2w04f6EC0nVWKgxer/eC3CmBgJprfDsQ8Kyma8ods9LoD3ysm05fYpE3Dep
71DNtiUpzXq1xO/RDdXOfAjpCnAEc5YKcIEU4xVMippuZzm6puLDmaC50sjxUZsH
PxGkgjJe9RNVi1eL2LaE/pAe+SEbT5kgIZwIhF04fjVawk9GrBqDo+i3Maa1yysg
FN5Q/1zIQgETAV+FeuWiJAT4nb3DsL5RhrPIaMxUmyj5TQHC8FNbMY04TYkMxgL9
uHY6xAtz8MG8N0lxnGbBqIIfMZ4F9cYDv/STup4vqo9FIw7MCTaUtc/NEMXx28QS
MoUarxe8JNmdDDgtFXdQHqi1+5dqr/Vh8OzAWoN1uYDn8QukvVDHlkExudp9yg1R
6iI02j15wM+ttCDjcLpVpke3mxfNfIBl9qTNylEhHcppzOf2b4hjS1XiCkPsVped
mCPScSs08tWll9oxqYs993EkrGmKOAlm/ZnmDCQrylesL5+J6nn64EX19ZX59t1K
/2iFmhZctCmmLJ6SZCrevMTrlNnJz5gcw8zKHsFEccmMj6Vj/IcbC1CJxN5t2y+4
uyCrUFLXxA1M0ZZqTXrIOi/bC+tuJSShud+ENW8kbk/Hr/pvt3O82wf4Ds01OWuv
VRkCIEap9RL7liG3P9j7DP/E1/oiG8bTrlKthqrdV2WwHe4zAZkpXdyb1nOG0dtf
wZWNCdYkgEb5u7ZDASIOGXvGZVVcVw7NZhtzMB6b6md6FXNlqUBbJWRoWAYubHZk
A3gjspcaoTFInh2gJedLn8XAyoN7oEQldLuGCPwMyCY5fLs5sl6r0wnNL2LDXAB5
VL3V7ux+ivwBayHC6F7V1dPMuHZZjYcSacDEuq6MG8iGxoYKagZZJ8PEICOgRO3T
7968+nNVnkEy3GUGFWJrGiLXw4wDZ8PwuvJVCVQWVm4kD4E4Cp9fPIc12Kuon1mD
2D5F53zzBjBRfU62qbGrSuIort2eqUu2oQV4v65ifiZVfuXsMeXSDD/RccQxwH5r
rY64290Xf4PRUXQSdDEeakP0YARdAUNrUCJ9aCm++e44PGGv1J59gpHk8YVruhUL
0Nrkvk03EG5FnEcOLkyjt1B6lj1pZem0QqGmvtkMT1OsYXiX5MV72rVBR2QQT7NT
+IuprcbSw4TMAEbAJp1MRXxdVCYiQWj/EjaKFdUPW8jne11WZH6dWrSmQXDeVBH3
2qSvWFvJPSA/FP163mUaQC6byEI6rDTAFzNeUh7PFboEoLFDPvntL1OrZNRr7+1m
j+zBBw8CCZ2gJNmT3gGnkItprrKkVyiDUa77Q31k2wAgSTD2ubDIHY6prTNvl/CR
gTcpWgIdByd4zh+AEYBNXkkRjG4MqhfwdAE71s+nNP4EOjyaZ4IGfcb7Jg6YUrmV
SExDJZj7wZDhxnx3LcnaNweyziCHMbiGG1psehgeJFeSk/ruvRlJpF0YRHLH/9Wk
wiDsqUGtxxjieGEcI6cmwOF4z5wk1m2P2BBcq6ne9GOt7J6DMHUXOT5gt0NQchYH
fJE8ZpYuHEPTWmuucNHAWqcAHPKhs4onga86fCgsg+rXkKb7YsWEZVNoqBZSuJqG
WH0cyixtfLX1zdh0JyOvwejFqRH5G+3HCqpqTBdJuual+/M2HDRkKoSN1lUEL57K
oY29Clj23X0cXArM8hP1vjyKxrIx1ZQgiujOhuU1di1kZjX9Z0y3Bho51RPydINA
RpbkwRwwHfRSdeoT8D8GeA3EjpbJ87TSWzvhgOYUKUI=
`protect END_PROTECTED
