`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GcYWM4GLM9F7u9ytfY1X/LA2QaoArbjyYaR9IxaiHvssKgMwXdDt5XZ+4xAn5BAH
nmKAatOw7ILMGeyM2y9PfYKVRIIgKa0dUmJ2+VIPjI9XOCYENG5URvbduYrgx3CC
nUciDmZOEQwVKC3GxerBhkknAMIf2Z3ZywLLaWgtVtmxKRDbQk5m5pemWXaU/rPg
yNkiaJ64EfcDfdCZBXe33Vkzlfvv+SUIKnqK7FGUHe16Vt+xKbpCvVPDyjj2iK8/
OsbQ0J67wwezbwv7evAXF/fEzCO+IdFnzVlOFzUaG/FVRGt7sIiWyjjXMraTxk1v
UaxROHZDWBQO+lirJmqQn74qSmm7QmoCtVMlGT11nsB02Fv/LqmQcYVQdSY1GP4h
KBxI3s/xvgprmJI3aTzaAYkhJjppazQaPx9iLS6nncF6F4j1oZIfpSQ6WZa72nqT
oboIwWEcUqoL8ih9FeK28FfFuRB+aQk9+B49gsGww5SbZT0YfJSMZ9T/y0bSBMqe
fsURSJ8gumCN89L3GDXJ28s790bAL2qklqWNm0VA08PwORh/oo6z7/KzbaxF/O92
+PHxcN7OdBJPkyzimLAcfRUEauCGsB2VJGzDZfUSBGxs0SvQ0UZ+GKhQsDX87cX6
NemE+5qBdY/CDMmIUSzZDy+Ckm4D3in3ohk1CQYQ4Vm2Bmf7ePijmvu0gz2fStJz
+1SbJdJdhoGWnn9NJVRk7hA9BnNIku7In2IasflqEiLwLjxHdPAFFpjehNq7M3EN
cLZdpV26LkbuSTM8KfqubEUWFFOt3NyQklNLp0ZfvYuY5msVLfWE39rbVG2BV6RO
X1fJH02iBsFDqIfG2LmET/1CD/bgfVudDVIugcbAa4zPSmH/m+tt2oAR3D+539CR
y6maAyO3154l5kkIgSIAzYghO+HTZ7KJxqFrzVVHPFPB6S/9+3T0oo3bkvVgwRsT
mH5FQuvRSwfxGklyxiAkP31zb/p+yU0FYpBz15gyfBtGRh2JV4V4FnDGXfHmmctR
4EFYGbOZ3JRpjI10S8m6PuWPlEhyTzfDszfO+ipoFztZmO+aIhoctdku1ylupZs8
LNvKn7fVh2LCl0QN52ELhUJ2ZGZW7OEgs6D1K5GatajAxmCh7fBLoRa6QpUjcRTH
b3MyzcWYQYCrJD1WiDcMujuLn5mE+dSMc5vsMxf8nV/ag6augCmfRS5X4gLIRhuB
OH19t/mtcfIwPYzUgJhK5GHDNRLwtMSxpnKH9jDAnlyACwoPYZISeRQrBCxk4dIi
Ucb7dAFT/qMEz2PafedhtjbhToCkiMNyp6MJn69s7ARP8M75WUzvqEbkHF/sRpvS
Os54hL1TP+vyC13kjvdZm67XKTJoWjiuDrvCZ/xyoSmEIJ1F6SZco8eA3sgxJkuB
HV9HVHTWdxkR4LpoLpP1P4iKs9EociKbdT5Zn9CSMZUptqnq4F+5ToVbNSgLQyym
ng40+os2sA4uWL3tLXV9iaSGSJDQCLpq07LckoID9hK6OJ/ZzpsguamgRY+7Tc0Q
GlVew7hvhtr6QvmwdUMkQB1y0NvfD7OMNCDr4kD3LeEpbonu3csIOZ4240thYwVX
c9zLKMHRWqEiazoNL+I3N4ipZxfKdpVwugmhX4NQ23B+XWRipbLNjGgHLJgg+1Iw
XK+80dyXg0fbaQbbjKPOmRSUlmD2+p8wsm0FrbDXbsxOyJf+JGs16jyfQsKXzFk0
j1Dpwm0hrA5WhEal3pSRcsv2S9PH5nUchrQzAFHhBgJ66tlGUSWOzugrGRgPo4n0
h0rJ3gUXbItaZ7Cdmdm+wP6mt9Ps4RGLxC6abelq7QeRq0cWa+MRfVLvxMK8EsVm
FeSd22a/g1qeOeC6Wnp/gg/u+KRQsD5eYdPzpwefm8QTPT5/1W7qqS25+MPqI/aP
PQ8+n9MWaQcWLsMTNlHjAeUWF9frVNDUpDongyVRa5EcuvDsvbYsVnGR4aaS2qE4
iv/hovTxN2VqOveosBHH3Ul3c4qDMBf/vHnAOxaiXAF0ts/eu4s3y/UzuhdSpCre
x1KwItK8FXtd0QnOJRJ20xSLlZS5+ZCc9fez6ozCKmTGPfBDUPsDznVf9kFR/vaa
sSRjKdh1tjufT5gBhl9dfcQXyX/zWSRLDS+5Y7IrI8fe+jteLXrxx7UAfqMGs32T
qMMvFDob4om9pDDVklbbRZLjgIoMQDSI7xyxfDCweK6jPZ2IznkjbFr2WKAY2PIV
qhdE7bUk86ikeYnClYVnZBf3CSAF/ObQlAuRbkKPM0pgajtgmmvy+7W5jEYTwFNy
x69MdFzmQnTLndpaRfIagzRG9nM48q8DXYlBB+rpAbVDoLhNJfA1JL/tLwbcYBGi
`protect END_PROTECTED
