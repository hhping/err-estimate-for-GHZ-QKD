`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+/7s8nF1NQuBh0oImUxosuHfnjTC722MaxBU/+mi78Yltm5xXVxLnIqviKyFLInt
ApzvVME8t++r3viIEZM6zSg/z8vvLwoIF6r41tyzZmAocWKfW1ZVkT6oFDMGn04Q
FVQ+EShKpKS/hPcZ5WLRpn0j4sBsOsMUCf1EfJtnMtsw5SV2MI3lVNvhACTQ/0Ke
mII7SOurfLEoH7fnqU8wG+numxLSETNy3/YeMPMxkut8wIDGGZwrVRNFqyHExMwa
niGVgLyHJbMMJkTViuvd3yEAXAOSKMNOgsqjEey9yRxFpa83VAeYhC34x7Jg067n
QbiQszkI3BvP7rXUOCQcfhKOd93VEEiKvhPXj9n3Y01oMBRlMbuycWgpVydp/bPx
uFeJwBrZh8IES8jpVf76PPpkPNc2ctAh5pvG3iUZfpLCfmroIDk5IA6yE2UOKX/U
HGxK827ScUuTWj4EHidHCZzbol0Thai4wW9C6vU0VMK1hrGhY7HtoSlAEcGnIB8b
zF2nbS91cuk03suvcNUR3y+KpEZRQqLD4+oGeVEmKIHaTP43k/TQCS15BFGLWwNH
BtFTQYUYbZZF/3e0lrokAUwktzh/AUSO7VldegASZwseb2SZHNxF7Sa/qZds0ZDT
YssFXoSkHqN8M6UTLpdMyG9receQWIMfg0MKw1mx1lYGmYzfMgXQ1VMQQh/pZMeH
1D465IetfeIPeJEej78u/F2a8iLCnsdsl2WMraGlV6dyqRPPm030abRLDP+pmsDs
ylLYxlDq808q9hlpMnrk9pqPqXGMFnsi8RqkxxHhsKEWEd6y2Fgz4dUZ7R2IATiM
fzioHQg5q6y/ioUznKkwbS56pdqzeWlrY/DMQvqObn8320rFFM0AHAWxYfimNV0V
dUshTe3kZa5z8iJuXbVh6ZIgCLlNSRvEIo5zd5zfPqZJGbhA+NuymDBfogCEDn3H
7ZfVtcXlnv9WvAfwjiIuG6a1qp4EAf7RGmP/NKinPPtFm+GFsMtxWYPjs41U4/y9
itJ1GBJY7s+R9/3gcO0tdHrIu9qZcTviDSKB3whVdaBUEnzgGa3LrzMF+F6Nt0OO
wjWNrqr6bsYUMJbKIrqrv8/hXn54tC3RDQwkA1gNM+hwfC0Mt0WS5cSchvLdIvmL
b0lkweb1G4cwdLrR+LglhhsHve+s1oPxqj16t81Ul1kwJlB2JWp8lhYdb7gHNPU+
iqImXME8GrSh9vJj9BNku1gx7FEn9zXuIuBwaLfYpOAd4CRyrGRWofxeJHRNgUfg
2n41s+cN7d9O4EGYyl/iGx5NVjOUG9hEk7ziSBZsPrZ2wXnWAg0gkdqedaOVlfbg
4WEJfGSeMUzwGLidL3CwP31jF+IVw3nZxswFW1PS3ryS7LRDUXrgAY3LZkWRcwRu
e3DF9TX1QKoaM7psXvtWe3yMStQ8LU0UySuq6zu7gTgibJBPydHa7049ydiNSbd8
0EZl1fcYhPqc3cIrmDoOqiIpReqYjbnAAlVL/uYsvS6/Cob2wpdmMaNa7zbm+uZL
9Vm8q3GSinUbESBZZExDxMc/Wgnl1GYew6XuI9uV2tohjsiyO2svJmUDXy6/PaKk
RZGLP3MRDOQrsfXfqjc3oZa/jD4LhPqX37P9hss2PVtCzqm8sHnJa+Zm/d8cWS/s
qsL+QYRpgChCqc84QAqkAsN5rYqM3hSTPbZ1yOTqx7ZS1I16Pc4qhMUKh9WueTGV
pkuf0Ny3wMcA39B1nW1t+eS7TvEDH0eSy9INEkTeLAQUfT642RLzc0vYhxrRYr9X
t06tJh2WuIPJo4bexH4QeCv8EX+6i2P6/n3xUoMii82w9H97U8leR1Rb2/P5F/R0
R9rY/oH5BgHizYgUjuKH4+m5z5g1XQKVlYPh93FLw2Eci+pbtFYVZUkKwpGR36n/
xjRjPNSXoa4pwVr0hy1pPNvcrFHj5PV81/8zra7voT/UJ6vgatxlK/ig3vu751Xb
aXt0NSToIXmzZrvTnoqn9ROaiWpHmC7O4eeHBfbthmC4vpJXb0FFP7cGixrEJiHO
5U/UUAS28BsJ+jd7aju0wc4nmgvMn0Czg464OIIB/wzUNMkRLX/BJx2OrLg5IyL5
MHdOUuXupA/MuDrqUZr1ctidCpYMHlMtDKNaAmnhZBlztZTyR+y8v1Oq1KVyBYz2
/BlmjAIaVHhRWHZ2J/5HNVgwlv9y2wqgwms/KU9Cq65cipOWRDP7t7MLAMLymWyg
XNNf5tajJb+2ZkHnC1BSOLy3LZtEBHeubdGHHmSy7fZaCcUOmHtx2AU3ZOJGnUCD
qP+baxUYFbbaPMBEL4Ew9Q40wgdDNldFWKcy7QWJuczyYH7i4ieqjsLgSBMC/mye
lkgysnmBB5vB4S/+jPBY7w+4hqIYOoVU08jHCpEsKVvE3DlAvUso0uLLWs1rYLK9
0/8+iuVLZYQt2eAE5YgnqEuq4RPgBvukh0O5KtptGGw0ajbMdcKlgz9MeAxiCVd8
fonL8FZ+DbLk4/WXP0vgeKMPK7jkFG6yOqERpQ9zAgCWhBUOZnccPkjdQV1HHJNw
Q67JuuthPOUg3iezycmZiPXH7LR9iBWZFqDqzYfGdnnS5fnU3ssQAh69F7iUkzK4
GH2BhT28vy5yiXXAAv1rsUS+c3G2wBbeNRJM9dXDK91tUsA7niAT/JWShG3pAf19
uwAPuwgmg4758/8nteJWdPKx076cJNy+SPzuPsCH3dSHyZF+OtZ05ciqXHh4BrUF
qRlT3/HUH76YXktTC5zOielZrxlPcMfabGoovJsSYVfzbie1gKl/KZGI1KU2wNe9
lAn7vVVC0l/sUk5if0Q/EqrdQr4Hg5yrWQAuNYP0N+a5Q9u08wcY+DYmNWfYF8va
K1YmWiKUq8FJ3vend0FdYL9AQtYDWDAKnRtzdWkNMMt1VGHK1L6owuynx8j5p4Y+
teShF1Ntxfh9UfBM+CUDNVJoQLiKXmaHken6cgqJyCHRVXmaacWnZ3nrzxgNXaGU
3kqViMTFllG0LqK5OoLtNQBVEFqL0foOSzdSip07zhTYbcPRWNtHQxH9NT0lZHxr
LrPzQGSFVaB1QvZFuh1U6hRxy6uqKSEl4SnUXESJI38XeLRHxJ977jUmmZOG0DcC
EIFGmXYhBOULGVVGE4/LCAghX6eknUdk4QeJ9bcDu6TQ3Lc9r9tAIFQGc1P1BN+5
`protect END_PROTECTED
