`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6y8tklwbHVdqvhSJTo/vB446mqhzstTCB38s9bfQ5YNFwtGsjpOGH3djQnKbDL05
fbGmzZ2/8Ru+8G684r8grcbFiGy89nBZPUSIomkqWS/N88a2GOrbGvP+Cd4rV+BL
GTfxnro/xWt+0tApV8qo9GHEfVu41dCiRO5YNjqEH/8/UjE0lXRosTZDbld9xfaE
ri3frSgQqxcHZhnKfkp9RlvBLpwvzbsF+7zLvp32wruZkj/kQMzb3PX46xUQ3K4c
KiJJviyAsswDf2Et0w3+b2ZHV2X3ARRK5zxuLOHM9umnS439fSX7QxF1HxfELcwA
8TneTX8FXbi51nxgDa3jGdIkfzaPNxqiRixqefeOJ5L1vgEhVB6Zj+HeI6w9ZaLi
uRkI9FFnTewFahhkcDxwoWd+y5cov9mmrpx9ZvxQU1qoWCPccG/e7L2HsnGTg/Jn
vKf/XwULf+aAr/Rkn5G/oO1AFbJYSyEylDK80WGJUSo1ju90zllKzllNi7lfftfR
uXc34e38sqm80JFr7IDDSeqattTKpx4DdZuLaeZ7kUk/DRoaVn6PiByDC/y3xfg2
seIjxIJdDCWpKTjoK2trsb71HuqKzcM7KSKisoXbxS2lhVVxM0vgEJ5ciA1z5xxK
dkGONWvzuTqMD11LcoBlmw==
`protect END_PROTECTED
