`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+WcVsLNf6Aksh4+oc8euWyNAd9zRzCP8+DEcnlLZHzEgmz+2ZAi/M4JiLdu+d8XP
2H/XdTgZvNhANuROp6Ra5iBExbNzzrMr+4vL6WMnkoI1KuQqOMlQAutu1ioMcoh/
nrmrehRd+3W2BPCT2Rd7OwyoA2Hjw01DuJpXVFFeET76fabMKkBlV9DACMjomOyv
EH1tuYlU1O11MOyc9aLAmE4WCUiOYI1BSRmXvt0iLjEi4ZAuWgn70+ou/8PW5pvB
Y5ZiBF2a08hoO/hD4rUM0DgzYNmot+OTVXwAN979rFfG2YI6jn2ejBn1St2D1ey4
FDdzcugMvjfkNnyxyHdYqnfNP4ZJ+Ekg8eFxlYmiwg3r+BHAbT74khq5nKl0UY3Q
040vaJM/FrrLDzTJthOY0jjEWuZaFGn8JaigDWGn233ioULiZyMgxdQHW1QLGFV6
4nqhLWjF9p+AwEl/TWMKwfBxLzzp5Pl0hQkBO9Ale02XWxkGmzzJ0L9rp0xAmZWa
fjJQfESCqscxL5VsdsmWXzmzArDe2cPl/U58LTGFWnfBXCTGy6D7glvvPJnOhxOc
4JzuyXF7V7NiJy3egGHTzVuNx5eaEh1oTMiWwAq3nkdfYXkz2rMb5pXMVLVeyIDm
fDWrNBFYozXnS94gHw84pp/liHR+UEcStHzeH2ItFbmFH7bnwou0EhEHdVKia5AU
ui8iPBNphr4kqfZs0xIBfAslz2m5BF9rInr3VCxEvgyAuF0oPKVyWMebflWwWvoy
sNd28UFqerkcLrTo8R/w9mIIPqGzPTh9N7n9LlYdz7/UupocJHH8HSZtu+zpKGRF
58HZP4sw9KDp8xcVOE91MrlDXEn86fR47K1uwWG5SpiNERhGLRVxwDQMW0aWDYNI
HiGunWX38l+ZXsB8gIKXED8Lpoak5qZhOzfF1z+XuQh0BJJNHhou6Q1QBmgTPdyw
jhkPuNAgBUwAjaaAWvCgUfeA3kLC8PDdk/yX0lj8KwvrwmOn7b5/4XoOjrnoC1ob
GE+S5Afx8GrYdBGj+wDJchWQqLlVeRvG2s2Jg3Ratee1/YlMbbi1li1knnTnv/MB
A9ZUrHvLHRWdc9CNqOhstFQ2jVt7ZpjBqludtUG2ioE1eJ9VfKGJHz/S3kIVsewK
fJAHiUz8Z82OGdFyTAHdNzJh4qjddc6eOn4HtJGgXJSFR3h19xmbLqGkEaWPBu8n
V3w5tkauOpNOLT6DYA6xgGJYjS6q/WARlu2t9xMhYut6awfL/8DGPPNNunhjy9hz
4ou0pe4gDIycA6Yg/O7ClyyrP8Kjm5CteFfyBSCiGbJ4pYmz+cRa/lE0pUUHvMt9
L49MEhCtWofC0ZhZemHvx5oAFe24Le8Wm4XqOY7EkCT6RcZT/5sj++faUp1Qnbqc
vCsecXoIeRsu1wxKzTdOFritWu9F+G+rxK2hCadb1A6Gv/VmHXdo2NAwLw7OlZWn
VVdiETO6c9/xz5yedpX5zpxfB1bzhep/Tf2/8EaQ4N0=
`protect END_PROTECTED
