`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYJHld4xsCy8PX1p7aNbBPN0RP7Y5hg2JutG+G8oVL0OFiscOpF8MTYfvrsAPB7H
/uYBvQZTHYM6KzmqDtRlkOuuZuAGm19wg7t9CW4subtkA+jYzm23a5cq3QLfTWTe
HKzmtHHtRzbv2BZOQtFxovDxNuxhtErA1XQCCfOLa2jvdSJsz+Bp+UfLxtNiLQs3
sZwR0ru+7LUw1xbm8aBD6dwou4emkiwJ97HhaKQ3Z8ejCCGnllfLKgN+Pn/s084Q
Dhj23GDrpFzmsesvTbJHtwM0rNS6JjeaMmYlhhzoHGFtAA02jwbuigdE9t8u5G7d
zMbez4CnG9HQGCZMh9TW/FnzyZXbjZHFg6vPOhJNWjTJkSXBtl1UdGGXisVjXYqe
GCxsNPYD2oP0SWi9yYHjKTQFOX6Ztdg3Ff2SurB24XnTS/89CacZZwsCIV/X9X3J
mOc3bWz4wqBVjNQUxvxhwQ2oY/n2reh8GTYYzjUDWwo=
`protect END_PROTECTED
