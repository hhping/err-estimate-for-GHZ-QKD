`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+EIwjb2YCPdBtLFmbH/ZFRTIFgDRcTGYjxiXj4dtf/kWjDbF+0XZ3dAoHVkHFvhX
fZib6FJRa4fxwO3o4tVFnLlFGHVBeNDXPidcsjv8U5/HMM8zjExw4Oeb6wGnCTHE
1PhF52U4TvvExey7MHYpx8fDx4tUeCN225KHXPTJZqHlyOAEW6Y9yy1MotSTUWmU
R/0oHlfaeIzund+q58wOmMXTqaS5qqaNZSqKnAc8Vq8/9l4ioNWm7QnK+Jap2kI8
gHJ9bf2nhS7+ZOGALo9S50Tx2tzM0i03NQiRvGlifQnvwpHgBWD1NAt1nUmoGomu
iC8j/891aA3zLrFqe6gTyPBxj0w4p4zi1SqvtC5/J5Y27nTawaRBdS2nbBzVjn5Q
f2Jg5mDyyme/Xl+jV/0/mKai49wQY7U0ai0NVcSytuE5IxhOCBHlAzGgOEV8TAqk
0woYda3BSBdlKzfABKr7UqrhsVpRDHOJQcVkgNHIJotSrP1emD7gLqawSz1DuhMg
OuDiVh++v/BYMZPhiSq7l/HMSpijRHD9cSv12Or2I/DYCQwA4ZTw2txTd9Zlxz+r
RcLMfD8KiQL8irwgKsPFFB6TKNt6rYRpvihD3K0d2DeX19QsaJ+dQHSfQdT0kPEu
Df2tUb6/GV9oddFemlHKs8OPvbt4yZKbz2UXYnfCZs+4fPqBP1cjfQUoxhZccvWi
f+WxUpv+DuNU+0Wp58OnEQ1//Pz1yffkCWx5ZLczTN+mrZXEUnfeN/qH4KLB7V6u
OdzbsRh0bEVTIRheEbpE5DAW5zMPVD5VmezSkdPLWd36Xcd0qijdQjKwSiLOvewx
mYSuaUcCxItR/gByDjnJCHDmQV7FyBZvmpW5fWvtVAlGlQB9I04nkzSfKIgtHK6J
gA5tGkxgK2+12AyAr7D8QFIYmLPuCgRKALRtkCgPjZNf2s4lO75bYxD6Q+OTB+ft
9hIng+vnGqxEGwg/vegx9MdcUBI8SYyWs5NCAJk4fPOsXW+r2b+RGPAvuOrX/nt/
BN2bMJuNf/vNZAELsCTTuYZdodLZDKkiKEi3ej/jr0WskeG5O0bHWi4GI5v2KtwF
lSiKbT5wREQntlj1F8MZyLKb/3WksewpLhBY5BDy9sSmdwid54N9I6n26yR4NK9O
fN3oMUsutu5ngCntozn7H+lGZ4wpCQSg+9eh0Bc71tqaqUfsofpi4VoDzlr/k978
9IGG5RzVtcWTCdgTUfRvaXA/NpabhD4POzqBiY6zDCilY3npjqAfCd5dXL+dV/6W
dKf7C9R8bM0y70YidKjeMYlhPsM2Qad0zO/WNXT6asXq+yY4JLd7DPXkrdHnNZPA
Hi9FfZByYcV/FQ90tgTyGsfMJn+1LKs9Wz/ex5C4yXIRfh0FzGyMTU6U8/jGiVM/
SJd1hsf2q0nh7VHJF0XR+vwypNxZ0uU5C8ns6KvmIUl4A13akvEeE214hYG/oaLQ
3T1Gx8QuUB2497VQAQuuLRRXZuRV6TSk9FSp+YEluh5pw2k2HQUAM3pLeyfQjs+w
u+IgTvfPE4TmornnfTQmMEh++kJGaGGa3Q5neaK9uKGz/grtPBOKsUGgx5CxY5nb
h1jMgzoknBEA5ZGAglNBiGLUptA2bZha05t69WfYVHSYNWCKvFhYmal/0pN4ZB0z
f6oaAeiAf31HnAL6BUBnQW14ncPJ5PA1fBhhsLTUcrvr9DUhdTJi2644kquqAmoP
1yy02zQ14icbnYMfLpP4u5RM7KA5tm5D0ANzQG+0M5QlndMcAYvSKKjYpQzAG7SN
oGJ1vgygUdAgfhrwxSLrwxZDTT1y9ZcXVSWLlXtGYYNhh+aJ1g6JPTxs4iyvtBQ/
zHlXuxbaIkP4Sv52XFVkyKvQAOh5gVVT2aDfOVzHVYm6tYJZzZ18WRNeDQWAoeDX
sTH4FmmdiS4n227IBFkEbTZruncahWNNHLRfzh7ybIDo3NuTAlw+FBMxYe8EILMh
9ocXKL1Y9PnGvEwD6A3hj5wmQ0NqIJGNqDU9bbkBT/lIKAMxBfRxPHZyBfQ+TvPx
Y2sLPo57FhvwYGnssiKB7A==
`protect END_PROTECTED
