`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHyRaDdMBq2bWx+AeKoTyaupED35eTSgqiDEdnKxQGANCXBNv0f7ujr5SNJjex5q
KUUV8sBS91PYKtn43N/eC/OJL7dwj9M5IwnjLeDsNenodS6fI5InKFunrtpo5Vbb
dAdyTo7mUZTAgVF7bOtv+NcpnPZtdbSLe5bFevgtHAWy8XwdLbE6WGNkpHr03aL/
Qq0snaaAm4RHcM17KAwZ4f+XzWF2HYX2nh/CqBcmiir3UeCLUXCElK2pUSB2gcxS
nfKjuwnvepzaB4N+y7auJLP+snxrKvKyMORX1gaC5/Uv7nyLNgQbBUk6tNfrmoB4
rywxG/bq4njnJn7wOF8Bpn9mixQGVMFe9QJb9vXHr5B4Fn1bbitF/eij2W2M5pFU
vyEAqAesGQ4yqwW66eZu3kck/ajTlkROGX6JdtMqjMtNBhsc8/4t/z5AefCO/amC
IGIQOabZMVyfvdggmVMO2GS0t7omsliTgR51cRpFW0YNExvIrqL2q+GjIkxTA3t1
RKjGcjTKoyqG1hPuiX2bvchDUzHXRjyId2kbQs4xCaagj5zXXbHE3+d+R0+mmS4O
/bBaLI9FN1vpOM+w0jOoOx7tFPNqrtbsIkXwr1xs8YrI5NLW1d8BePlmqC3FF86t
WhWZhmkH6AcOYyp5tbeqdNurK8baCpTqExY8p/RHd5r4Qpz9ZoBRYG8m+W/xUIQk
QFsvfP3GKowWEXvVsO3ZED+SCytZqLX2So4wrFAnI93sdqQCqn7vSUwwF+NfSRG8
xPGuSc6U9a8a3R4bPJPzvn1+LXLwSuPv0/BooFflvCJcmBv7obDAkkxmy6q09bv9
V/CENdCdVAAm1Nx8LLuRGTmGKAbM9wHDE93rBs4NM+QguXi56ADDbObcHW0I78zb
rIKuMH2NUBBUXrwxGwHhsKGYe80z8hGT8x74lHJcWg5+PrFiaoFcx4JpgI0VFZbd
uaCUwZlhZIq23bu6nuXZrh0DN0alh6oFbpmwzNYHqzoKauTs5mwcwTLoG3i6W6Q/
`protect END_PROTECTED
