`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gI0pY5kszlUpkPCdIsFrz10CT1oJV+CR1EDKDlzy+dvtu2hnal+7lahjpsFv+FvK
lndCUhvfmmZzV+hINYP+vZMBgnE3OpTSPv0oA3EshtKiujSVJwe7glR0/+T7vnTq
aKpWbbwtZH5GxGV+2NzCtLo0uIsIYxmrJEnKMn5T1tJ6XmD6oLH8QHTeZzq9IFVv
RAIqtAJkRuQxY+IAysvesgnnTuyYdT6HNB4jcOja3N0M7hh1DoO0GdsJj0UM+X7E
vHF/ncIuzSgcaWYeR1AAh7uyLYhe/TzVLus/pGNmtzMhhGWAJOwglxB3IO+qmkoS
8CfzmuwC5y4u6j6zaU4Zd6By5H2cyHk6BKHwHe9XRRlQcT31k6TnGuFoVHIGoujX
4xljZBsSXSnZjf0cpbR8DaDIXc3JJ/9gyH+O7/jiBGl5IrqioCK2ln3ERcRObLtA
jzQR89OVmYsHPCzSlk7EANI3MtWAHGNJc6WIZji3w5QX4TO1dqwo9MsnHqvGU5h7
MRrIzH0MQ0KmUtS1VBhS2qMUdGYPo9JUmz+bsWmBAxuxg1R5PAjjPny5OVY4h7Xe
9DYIjgkVzJWXo6VaJ5RmI4FcTzjvGC9vmE//UUEh4P8BMz0fUOXZAsQxdWzZBM60
weHsjHxr02Tl4CWvFC2ulS9LaKdmijUkQ48VLnzO1FkC78GfwxAcwlY/mXMxiy80
M/GVrke2+Jgx8rm+AcvuaY6qyTuK/O/8IAviFMIHh7CPbpLpIa0L4Wy/PZDLYnyP
4PYrLyzM1PUivQizY+Tnp3t8qPXKwzI2vB81Kpvm2roVeuNE418j7bo2m2JHR4IW
ghCgnpHxmr8DJGyAC7h8c4wJgYnVJ2XHxOqVuKLQu5yXkivq73jRWTrqS3j/SUcw
6NnX2kHyIaI44uwCLfx0HaKMGntukThf9WqQaT6CX+O/hTchLU5nTDUREnA2QLJ0
IOL19qS0AIjtDJyvbiL1MZeBJF2eDyYrC9QlzBPvM+6nWOSp2/jpGt4ZEIXRhPcw
L4OSlO7Ofx+zHlOBtwhHG7N46IoRQSGrHUpteQjE5X/J54R4vz6y5nKxxS4WVDsd
6lgi4H47nxe2lDGevcyWcxSC0NBb+RA9zCM1oumY++Xhu3x7iAzxg7hYw48mpiDG
tz0vE/Yd7meN31bpqv5uRCZ1w8b4UA0oO9PrnBlosLIuHT5rAB1VqF268C9ZHY0h
1OARTLTa/7RaFSWJOqrayVia6fLZoR4DoMGDiucRCrQq6ekJb+h6NljPW4X8je/W
i7jtKf1FYIVcRmaqjWS8os56h27VPYAsIBvcJy0zr1xubp5oZMsPwuaV7d+FgTw/
apSFwN40la4tdfMvbEWJjbRBbaW7SMrFkJeUKiCbSt/k9U9R51q2497sXvMpXLRB
cloFNBmYQW5wEXMA06A4KlUlMYMk+SjVcssh5tJDJCkAnrjfxoCU08ZVN3wCLxks
OOs6z7TaxJqRTzbWXFZxjtvrQF3NOp3wGEBhprP+DjDQ0iqMptq8JQw61EJVsnaM
77EiET8+L/O+/ZRSAj6h6abnFhVXyT8ZimFwik5r+Bcpm/8OMjikRUz8v14gvSZb
wqIKbJioTQGKxL6xIsNn0kl/8eGHsQAhv+bf9FpyJtlnGCMSl20oEe7cih/RR7HQ
yVxmeJ1Up7Xrptigao8hagWf8U1dU55bBZ/ZGMHqe8mwA+usygz/8KRw3ixh3Gew
aIcbEr4zR+hDGlnNcwiZw1vvClXagdLFnpu/GoX+iaOufKVGbnFQSDFHU7aJNRcx
0uhus94Jo4FagEL2Idv0UocCUhmSF2UlIHzgGSEsG1/IGHfrrkX7iFtqmqEt0NJd
ZcVKqgGQXhIPd3YTk6yoElVoRpDL2z+4/23qNVJd788gt83gEZSUGbOVXyn0ui7Z
9j2yHFCq6z80Uq/Qcvv1klh5Xk8DrGQbQC2yj2owEU7n30bfqFKJRZXvha3zeIeR
3AVzNhIiMUKJOgrE+lnYIm7Jv4MN6CiOx1YIK/2kSbdiF4wOm55GqEpH+WDy6o17
1wn0r0Fn6q+4rjHwKOsLPEgA4WrAEjyewn6EOm7IFyljphbHF6fWNYnsV4V3JNHQ
Vmi3jaYGF7sncpJ4MIhaBvA8Lvl8QppB9d/pSK73E0ydkfH8VUERfOwn2K8iuZ8w
Ob0i9T4hm2prknQux15YWpwbkdzCAuiebZGAM46w83uYMolG11FO4Od6seMbb+C8
ZjNpeaNCxC/YDhJbocwi42GB5rYqAnDtr93CsQbgpZe28r57ImqU2LDeCe4ppmeX
ady61zLbvU+E+swHHKHk5xNw9hq+lpXhA8h/4iTnq+SmM32saQKKfo5p9X0SzgnN
t91UAyuSNW/jacS4YZrqTNflsPQqwD904LeR+9hE5FisDrXjuHkdJMQKtzqjSZZf
li6mAtYOSpmTvcCHwn47S1EDXEGUjRiKS5DbXbrs/qqPeX4Y226QkzUg21Frjkgz
WCWbajLtcJrCBzNig5jmXUmwC0dk2t+8U00iuDxA4LivCkn8/QkAoeQGR1h6X48L
peLYLrTjlWtjoCrsXtrBLztHZBHgHsUNDPXTyK74chg8L8C4s440GdO76MzXn03m
D1LAfjPlEEQU32Hq3Qj5PB2nTdZZCZarfJJ3FRtGsqS4aYFSDS39+7dvuEkFZONy
GPQYifH//K9I4WXocpNUh4IG+w2o+4wBGlTugkqgyD9KI1j97R1LbiUHK3UWS3qa
hS1twrNeTm4AMgBIrJu5Lw08nJPzEZU6nc1oaSa0CvfKVapc52j2FRZlTLXh452U
lh7ovD5pK56fk6XL805Kahl+41FtsQvSWWVOSwCcj5UY/oERhuvDqG9vgY14bMf8
kBwRMDK/34aeRoRFsDM7wYagMEiPhlWtz4XSJxdGek0KFNPF/fTFk3LjLFl6hTj5
TOz8Y8LUSX5LflVtwfaS5fjKt4oFzVUUvnp1X3rNTx3cdm0yZg6F4zbOSGW+Ww4v
mYK5cS2X/B4SNouJarIJ/A2j2gOnsPlHnB2Una2vzBizbGoneB7uCVX0vNBeTEv3
ZdE1zIrwuttnFboCoWJmPu+4kxJJoEGOM4GBCvSz1C3CdywQCpmQatacWtNRXdUq
zgHUQN9JkyN1LT6u0iabg3GY74EMfe4nlM9X6/DhUVr7japMNpwuFn0/h40iIH3L
l7CYHqplpbuexx7gv87N8sIUWJ139pcIrWVFiOhkcwMClFHyG8QnEeV3vN1yE1fa
cCF65uqRKa3ZoNocpDrgB+E3++qBp+nS/wxsq7HgURUJ0HRIIXVOoA/gSQpSf3NR
Xav6mszWhEqWEZQ9zanLjd0Hj+wHBXLm0oDkw6MU4eusXgrSYrQLTCrAWh0soPdb
WH5tACpVry6+U/lTVYZjiciFxu6kdi/Kwoe+jioJcNGzDvxLDUq5Qm5Fne4fFoEq
Qut8Z3wOwzQkIWNZwuy/Qg4t60rtiebWSvEBCGPlTMU31LGWv7nxkivZ2XUstIU7
6783q0rRv2GVsqnI71QXFVqWzeJt3VlZcoRhxoU5uEE1TideD0XhAWV4AEuWU6dy
4gR1FMGwTdXVWLXz0MCdXgiZoqUE9Caps7eVaK/KvZD8u6+fjzEPxAeb71QfgseJ
mNEJkMH4Zp78hdmPM/coyy4PyUVoNQRXTBP2I/OAqcR0fJY4ZUkbtxM03NqFc3bB
5IEnDQO1l6cXoQTP98QEyhDNl7wukLkFEG8lQDoqGXbclyEnSZamG7fxYVm/MYVs
QonbNenTS27z+x0k1wILTPl4NoTyibvz4VoLCcoFL9XyU5KEqC4HB6l3yw/RY4KZ
0hZ1LmDWtOZ7wmOsnkKrINFeCy2h1JVF2rZFokwwkbAkEDPyVTOLK8haxaNrm1yd
Uv2PPl/EGGmAkw8YakMcCXUEyeDr2UtZksiSWWrjdMF348AdJeSW26ouBbOKqMUP
VE6X4+naOZKSTFyPW773doJdcQk+0OHWM6NPtv+9jFeSN5Cy7FOHiXXduRUM4bZs
RWpqoTaPgJ5zADxsVnMTXwVDOpx3Ali/mV+9uLKhH3vVU1/8mY2wBVM1MTRdTGCE
6x1CYLtpM1ULboQNFTGhy8gCzrgrvvpQnEN05rqVLZBsCzP7MPHs5mb9XHH3Q+xG
4iIkC3f6LvsKN4nm8qZqa3Vy5IRDm6jXJ2npxsMQzdvAMJn2C35BiIOZ7OQBwlGR
OwrvvDb0I0sVJSlUbrbZ78cWcc163+612msSFDa3yGwA8D3pNksDIW03nRqfy22S
7qVgVn30wRoUyJWDrMUqRX4ViK9BY7yABnUjkNUbQSXTcv8/qcnmtVtPl0dsIDrt
JmGKknmqs56j6DWlwQXpV+5TjdwDWkA4zPIToImzZhYRZ9mZBNdRsc19eXfNttXR
fP91WkdX9YhcH4DTVF7Fq1Z2fEV+6Z538tOUyoOrSPA1lz95WPAGoGJ8TD7ac4+F
fGryl2g3OqVc8m/NKyfZ0LgoMfgFgHbmTUM7rufzA/pUv8SM3xgtm91E0Da2nB2o
R/ZdCnPc3TjV9PjIFoieQzT4jSE/QaQXrIBsSphRTvLR4jyI8z7uQhrrqYjUCCiF
KRDaOhgV8Z+KilK+YXDxSVAMp0AI3ujNCmi0cJfCssJkstrlv37DHEOo8uypMS+y
c5t+PRDRfyDG5WSYv9zo2C/i2pg6LsX07Aw8vdw2CTUwbubsxYsBMzsVKOXlj89F
3PeHChntZeUDwpPL/P7Uvl3o3UbQMRriCwQO8AKz6vyvUFaOBp+P4lueojLL7LXd
oB38oq4dX41WFdHpz1zpaqLSYJoir5hw7DKvw/TIAiD/w8+qZs0C0/f3/9MnU7Lg
iTR9OVGWegOx+9x0AuQ0pE7Z5kZDrSOvjg64OiA07al27HILF80SeUvv/JUgfcUj
K9aG3uLqJOc1bPrTkgZ35tsEoRFcR2xuA0itFrGDr5AnobSc1qamN0ovf3gTbv+Z
A4xj/gPL0EJAWAo41IhXWAlkmjLyg0z0conaSf/2qCzHw4qWiEsWK8Fs0flgeqXz
VZrNWlGkkqaL7a37n1zbi2xo7fkQgs/jRoZjKKSmUYF3SRhNmzsA3dai6+dxq7Ww
vhZ0zVKzNfrJyXRMfzj/C5FIWKizp8ekwLWe78usPy3pkypgzwAEjPxmKOQJbLEK
2PuILdQ7CBKLOBr1F/hy2l0TJGZw7BiIwJgG7pPdtvRt9DkgOVFgpSM8F/YJ1ygP
P0t8agq8+eqgPL+k6wBny7/2Qz1cCT6gF8aTPZvzhAbZr6mxeVNr5X2KHcMvvgFW
heLvBl9/0sASiR2sl+X7Em1SxdUpBei0QA7dhMK0tH7K7yizXJbKYEk4nbJOeQiX
RA5zeIG8hbJ/XP6wEmNJpWn+xLEYYjGHqTnBvpBa75bm/clJoWjPwbq2TNxNTWUu
HzEEpynDufohxr4Wlt1KgrG9bE6fPhER6Sc8d12/nXv9tDyB3Ty0oOU0QDeK7qsm
XFUxBmjowwVM+/9FPFsvw8WLGfABBIQcxaw7vm3PXK2R2Nl6fvJrchb4dTmheLsA
1GJj7ehEWfCVhaic44Gwu4PhHVLBuGzNmrasMYiLKZc+5BYfFTSlICCHgtL6aieT
dwI8sJr16BX7utTnjivYx8NOYfCO24x1osfsMXMvrfSIQSuoJdXh4mG1r4dthExC
EUeZoYwH0QW6rIK+JDeVgsatIHTowcRqy6JBNZ4jMIwVWzvJuvuRBVhYVlfHamDl
Y+1u3fS6LBwK+hke/lT843qWnGbSMjO1R/AeLt6T6GdPu3zVKpGzjaKQXViBOCPA
KjEqI/AdbNfO2V5DuIFQnJxE97pEvOJjeZIdU2hnfMkfDNKI6WYyblXkIzCrq4VB
ooowCPpO01Tw9wxo7WmkM009/82wCZ8CRu2XRp0tgHLHrdGHwtP4TIxBJfnTVyjp
oFJCrFwDsdwtgQ9StYcpZVpiwFj1884PhG2EbaxBGeUo7/dvPf6m61Quko3Nj+I7
5a1mK80njXFwbQKVvLrtX1MpPEBDEvCe7OUx+Oyz57xql2S1ppW+Rt+4vVh6DiYJ
Q2TDvOEXDxUNE/qADCX8sn9+2SYDvDKPG/IRViLSXkj3iahhJqGasXGZBZIYm+hk
b/aA0grKrL0ojIL6NYEjmjjAdoJ+b6DsNC21nU1ZCtO/gmmUA5jIiqfPn8EKZ4Oi
SlTfTj090q3Se12EBETCmlbpJ8z8T9nxw+fKFF3tsunwoHrdowJGfyu7AucIS32d
lW/X8JH2M1MGqdoEUT7iD1rogdXs7DODgzUG1PWlDA0D6mAMEe24HyducZ6YAH0o
vxw59bXyceEKQo8bp9CI30RAjzyi0cdNuLc9qu6ySSoi4rdfAZv73bMqiLYSJ+91
29aqZi+F8mesg5bhGEFB9VHmxA2PFKFZO6nVwZInHQcsOp1seKopL79g8Kb+jFsT
q0NsM8YL3z37kY7UtaQp9bmRO7yNGxHxyDCR/tp0NkkrHaxZB23HMgnK5huTVOJk
QFQBDm7X+5Y7Nc0pdJN1in2qNzwWKCdOwX36cj/vt72BvNDAjD/BdwpFyJWx81Mi
OnScZPt/t2E2hcsFRDE1Tlzu8BFfo6erKqN4kPkr2a7BrMOZzBPCWeOWbtdMHg3I
04QNGwMyFaMBphom5OsQabHCbQmgdffOV2GzZvggJbPzjfGdsKueOwaex2uIdoln
BYVtpbbM236tlW7suOQleIK6jn4qTeHuFR1zwto53+zhV+iEJuOQm89+swhR0Qhi
1EjhjMJM9G4EX+QLJbNO8n9MPoKPqZfve9QXIv0JcNezU70qf2Pj9qWgrIIMegnw
7nzpzRca1ZNJ2VXf7NF4ElROgiC3a6nmG9bZgE7LWdIJFrDOkH6i83c52jooCWu9
Xl1E48npc6HBA69i7JfRtvekj6yJn9tmLm0dq4kgo++xNaaVD5nB3iVTZ+KoFFdD
IjJwduM+d5r6KJmrRUDZK4idsVcCr1iaQ3iwRzaj/fT7NZd0hyUw5Z/S7GEQLKI6
8JU40vOiY2rnBpiZlrKaArSdvMQ4FPkUc6MNeQHhc4tUrXB1+oWdLnvkrfz8Cr1B
n3w3ZWsO6BwTvZpbdxIdK9nfxh7+TXY2i4nPUSGpo8HbGn7sKg1NTxe4wItfaESk
sOAnuENf4XJWYDBzEB9lyxZbSe61TMdcDWTtNZan3hxWQSkYm/m2BE1aT8ZGFdET
N+MBxFP8MsjIMIgoZHbcV4gviGNVtkXWqawMyo9fB463NGc4XxBVOgMT7F6cOEEw
uX/XMNK/6osbaoqbNnwtzy7t+7dnD4K+LWnb/nO3vXp0GEcHk37YQi0OkvxqS/q4
Gqnc0xwokp2GCc/yIzs5U1ZrVmIIf1V+PhDdk7dBQZjzRpoBtBNmOrYX/zwGOUp4
TyXWS/hLyeKES1M27z8rywygQXWB38cliHgwMESIL/nNYLeERqraz8sAlIyRb7DB
X3ddUidiwvim5r96wRVBtJDiY4tpuwZVZEf6gQ1ZN5Pp6Ynkxjd7P2WOBguINGHK
29yuzpkDkjVPUZQC6K5cYVWaBPvPCXgqYo+0Jl/3bexMG7ALeDPBuk/nIOPc8shl
GFQ6LIV1vnxhMG1PDNNLTJcLpv+bS8PlGs4qr9ihkzR2Iu5sO9SnVkJDtE6T2iI4
sFBDgXgW5Bog84aYWZDA8alrK6C435vqvCsC1786Sw+FcV8qVpzEvmZRgd7YhgWk
gbCVD11WBuJGP+5i99cAZmOOaHDb64Ntm68kHP8H98crh2C0X5GJhElGpGEkdNe0
oSHmqoWAFsio0llsGcoQuifp9wHEiP8xcpkfobMC+gxHm9QkU19YDuaKjyj+Zhzu
l7A7MRE2hBm6v4LtBxX8pELkRByFkjMtuHhylahDFa3gBcFjpRxE4gb1PhDgThaX
rgZduZcJC3bd/1VReNV4Lj6bwU8P6zHg5Pmkc0tKeWtRjE3XYRmqj/fy6TwX66f7
NbnqJM9MfF+tzCPIj7jhSSPW0ZXJbRwD6DD1OI+uC7sB4PFo49dDNZSYETZpHxkX
Nfpm+lZfF+f3e50c8jRBSK8zVZCMMzCfz5JiH/CEZSiQGboPfR+Rs42Z3MT2olvb
VcBqZJY8IykwQkYBZe9afD0fGZX6d/cWtZzGfHg7tLhc64YCzjsT/ldE62GSawYW
fkTqo3QbAJlbvZg4HVVjRqeZqnF2e+Yr2cNtVgLj9dxHmd4Xl3K39up3H869toCT
NEe+Zpoj4DD7OLY+okc4pezuJRBwgqVZLcNQJ+D/fkbnvM5FO3JWMYi7UZTXClK1
a8Dhyng82DHbXB89Z8IPITbrEy5y5DKVvnzptPipR6ilzgw0zyQWOeXZBKdmvOpx
2eDnOQ1/f915x72f5xbeBMO3RaoDreUqTov72uAYor01+a7hBns7fEugpUaE5juI
y+ALOM2jSpegYzzYCY9iPGP9Ss2ng5m1+TGnwQletpC/gPq1Uij6BSAdtXpE0b9+
Xk3yLpLyUidxIbIVm7R3C1t6wVWx9806F9eUnUGE+txw3kwiJhBfM734yj62KWat
kOe9M36HDq6zNHv7e+OwqTsiuNF0l2rAj6gq1qXZpH+kwxYr/bMf/XxWq/0It45w
RqvN8FR1xKsxpwQE8lN3OEC82xXii9MW1+4rvBe7aQHmwnqGDbM8qiVjA9fmN76+
VrYMca1SIWeS4XKTFVAENbH7l+cwWSf++Yfiv1Wz/JCy3LHo9ddXzRwrujdKrdPQ
/HpMs/xS0CdNn4vXfetMh7Afve7gVT6Ht6tXOo5BK8654H1g0hyNK+/w93hQAHYL
m8THRb8cVsoR9p7prO8O7U8NL87lhptKfulbg01PXYrkwenb4Hg+gTz64qo0ZExG
+xSQiCu0Agg9FYQ6H6X+r3eJx9aVJCs38Z4AFHe5sWpP8TpMkBA3oYBL6lk6N0Jq
fGeAycaKYIt30MA5CQEsJpFSjsGAlZEIZTrDUJemP3iUSay2AG4p+d7k+I27hOJr
3QK14PSMw9DweovypXEnjHgrdzjKqc/Qlls2QNzpNNOi1RyKCHwYzUUsdVC9c5Mz
mrXL2ga/NjPgvu7E8XUMRh5kK70xknklqwm50x0klPIi3BzOipFKHfb9RHBWEY6Y
1+gle6IX3vIQs0oS4HGIc5LKpZ+aIp9okGl0vL0XQOnU7C3lTuGwVslEE6xA9zqY
E8kTuA48z+2/+PYMWb4CrxW39PLA+3NWyOW3y9aqSD5hPR80raJ6eCyA+dr8UbO/
8WKOobridVcyx/cxtVLDWptkBZLEaNUounRGg/DvRuceqe0IrqS37cQ246eYptkU
UVJFfbnmo8wXIyfhy+3VB2J431OVS4gTNEYio4xiC6dc+XGK0e6gvRxEoLUQCJWZ
cHVIu0mD9XgL6KKlTng2SZix1ElmIf6K2wM/5UDsiV5uj86k09qyHx1hz/Xxa6kp
bOnzskNtiU3QmVDQ5IVo5/tdhZfC4aisPBvbouKirx2p5P7ijEFCva+iNUynfm6I
p7z4MkVoPXuxLC7y526oxpSjH4vX/PPTzQ6pS1JbLt9nNuX+0MLaTkJWV46+pQFJ
2M+b+p/5mwX658+TzxOXDd5r5ZsGEJ2MUS/USAPWsDM0WO2i5llWUttfFOcm9rcu
ZNMI7SrID338cYBUzIWRtHOopsrxXT4QcjXkhcQCTcdgSHxOzY3GASB8fZw579hY
cxfkOuPbo9o2wrQKm/fndr93iA1GeOJLOqwBaJxhpUT4PPFZ9L8vrm+gCbmJFfWf
OEFxwOFxpEqowoauiYwVoiHbB0Uo8Brm22XDnZspDJ9PIKMJNztItys8bGfOZu4J
IvPCBYxnYGLuU7f97ludwQRb6Rh34SboFvwdl79V1Fm/Gm14nJGtoyuH8hx9hEYv
32BfF1l37gg9dpLZDljeq8PlMrgyAWJANGkvvgfwObjiDqLvFJ6PVxfTm98qTUJU
pz5uPio6S8Jm3NIDEvouVEGW1UAajlHWKR2LLikwMb530XQayiPTB2mK1Bqo1z2T
jsGDN9Dsw/pbnWqr6PM9H/yVWCyePvRIESFZC2kHgrBSobOCqjZrE2kPXGA0k1UE
1bK1sEUkLpLlVTcD3zaGOIZExdTPJi24B9IQwaV3eaJ80IwysisIEIaw9QKl17E1
1tg366vfdHNL/uwkJ6oLpRdels/hntjoARUxVxsC3reO8SxX7LPxPpP2e8yHWtha
y6zv/TucfAWGc8O390kYYcKHgC68+DdbnZJ7JJH2zjEQKovrbdXjHQdEYYtZ0Hq6
cjHh5QBmk/gaQkGWXKeJR/3uKSVt2V+uwFqEx83BnURtqGuayFTEIbA4KqrWObDE
X0FN8wTutu2hupjyp8Ej9Wktbi/zLMrYlkartN5/aJ/Khm8pM/GGPgGD/BORGC2X
7taSwg52rT7AFavmNHV++Qw/WyjwQBZPvVXnjWgr20+o3OFIBO2e1vO9T3n+XLMy
T6OHpQyqNCN3WlO9qloe1O5yG4AdYGPnMRAr24FMkIWGgtSndkDiDAr+A/jW9zHN
H6zTX3R7bxbKUTaoBz4fjPAGIpf9r4n+HadIiUGgI1EBksZd4ELBDDs+IdH73gXm
RqQIzjTCqXnN5EfxuwXs6dh/7FqEQ+nWwT4jzcKrm3U1WI6rJjwBZIdXvk7lYkLY
cguO8x2NwZILmRyGQX1bMejB9Nbt3OMWqPN8SZM0fcN/qKSQFn99GFSvTmDDzy87
2BzG+B/OHc7AGDBz96rjA9I6ao9jeHEsciXtSYOyNuIYAdcqAB2rjdiX/dH02G3Z
TZ1AvBxJJ33ATkPbc7IEHs+c7jci4p/bThMDFUidX5b0eFGjuwAMS0MrGKt44q/t
dNWf/SlWxwPKFqD5638OPznlGKfM9nAApM5kK2cTdE3TELo7MXkgS2hmR7SQWEo7
xPRy8VTVc+txrCWuiC2wLG+i3zJC4OvRIUlDtipbFqq2XOYOZv+nuDrDDk/PhELa
iQDYSKCs8a+x0/12xSd1gj+yXiMJF71w8CrjxxsfSPozqpNA+oBbULzHhhtqlZ8x
9xFzfXJCd9L87E66Jx6r5/xwrmdZ3aGPGwrB6y9sP+yDw3pj8UI12fvn8zGLdTI5
nOaTieXvyj7ATwpKoNNEXl2+bboHmWX8Ppeo8lV036PiK00JAuVV5GVOxXtQyGMW
oAy0eeotYpEZqdZ9CcFsZzgzDSFbjZO6aiVCz4Uf63qWNudgS8DOnlWGQrVW6ECO
oqQhcaST5ZS2Qb3R4mcol5n/vbgVeDaqNxevazUhkTGCTCgudwauLQ3QHrflc78L
SDqc5nrkl49DYeZIkTGW5c3KwBgS+wpCXfvVsb0j0bGCN9kbWHdsxTNF5vQ270+Y
3uwSDodW135sCKvKKKtLhS7Ffm62L+T0Zx17YyHbFzeg2E5b3Yy+XRnLOqK74vw0
6Y3j8XOV1x1qFRHYR2awt7sK4NiYRtmbXVH1azYMNVQTz4++jhuxS0tX9VvntcbN
NTrjLKMLOEQQ4xqclwn94/kXWuh6OtnsKmGcaGOFV7HoQFTgdwa+6AVfLECwdZEL
z4cZ+DZFhvz0MvjIdbJ+qArATK/F8OlTq9BXl1zWrZRVv9x29RFgaztlKruFjunM
AgTxckt6SoVS1ji0HLIZEHyGdY3JpJNUaIrla+vnpQjSoQWG0YP+U2pJH3WjcA5G
fl272fYq/XhsmDT0btEm1NXqkfImaG57yoyJbQBXpk3RaPcPmny8bn7KU3GNdh+a
KFle0EhLsgqQ9TMW2tVGdYrnWdECwxR834cTYna3964pwDjwrIqwsAM772+vIWLx
wbfxjUQi2tRJyFAMtRGcc7+JLwAS/G2bTDrlAekPaBpH8zRiwpB3IvivK00Ee6s7
bONzB9BthzmcFgF2O5D5NCwag34ma2bFBEzorWtww41UFI62P4lbHK+xsP2M97Mx
BluO1zpq9n2YEz5J+eFGUcR5tou/P9AVzuoHQwLFLs2/KV7M3bn+TAR40jrJhL33
oETY7/N/RmaTS7c3zaj0In11T0xmfunBqlKzAmEPugZ4VuB4UWThiZYhcC9Dcwvj
+anL1mBjpa+XetBAbYa5yCcOLPetBNae5HDtJOCra/ROYWipeQ3bvhz0qO9ymqqR
RxVa6ZmSqaLTILsECgqUF3uAv/IMd3W1kopmDrNZ1cwBeV5UkNwIjE0KirYL1Y6r
jnjcMNJHyX0KKR3KjWT5oKs75vGLvMEa7FSDwlUVVY30/u7E84lUwmVvKhUx0fbA
9hgj0AtNIIzaK+cxYOrG0+Ji8RdJNemSOcXz2esDzuOkRsj5+aDevaA+Z4jm+bBE
+xnrGQ7Gvu5orjnM0OF1nQveKi8wEtQDIX+i5BTkziQ4YE7LEmn1NsiSk0+Sjx8J
zrNevvU1NCjRGJid5gn19LFeaZ+76knzDnbhlpf2COEJ4kWTpSfGrOJk1so9lZQt
49+ZwKG0nMvVyRjMx+Z3UBb6W07mSEHOqg95Vc7IxHOzBpFSrb/DdcR2ZXBHB8+j
5jdd4yINFXjfCuTRpvuD/AMiXqwOTJsItDM5aDogckVJHWc1DFcO1JApf3as051I
mO65wuZID+46pBDIkr2apxRA6oTsRkdCPuD6kvlF5eLBqXFqmkjpmJcTBlKTrXWV
H627t5qyfRhyVIrv39V8gBU1tp3RBqZKcoLF+0SKo/GMoyeRQPMXXEp1lIIUxSYk
DDn9WAJ8l1KChPYmVhI6T6Ip5ta2jZ/SLgJe+2po6IsJXkcNZLvDzh0KvEDvjLcd
c1CWBngTN7xDCSO6JFXnFlFun/Bf8Yx7k1w4giDS37Vwbh0F5CvhlXXl3JxGdKQm
sipJDkYN0IRX6d2k4E2KnBBf0kTaYRktjhc+T8T6q/nuDmVXBF1JmNeO2MKoLU/K
9i648rGBYv0Z1UV32lvvDtIm+FnDk+xtmAzGEtm1cpK5LM5DQ7Xdrl/ZfF6evAP0
+MTYhJP3vuDyGh29h+AAwhuK/OhkX7MYmOuURVCO2SyCaOUeby4nG9sZR62f1dQ0
KpCaQHducELqMUJW9dG2UmR0c8wti6V2YMx6v/gEIShPe4tHfhVDK/MSj/cHQ4hE
uDX++9DLoUJGZFlNAX2WDFJl3DuFVKIfqNu8vjbqOPiNdJa33dLW0olkt+2+MgLl
TAfbiPaD2Hh2cKi+Uho3DiH1BssepilszwAWrslrW4pmq3Xdr58DZ95jqjBIyY1v
KSkJO0Pnr+rqVFu2VIP7DXuMD41uz1peOca8egrXkX4KCGbQMWBV7ERWkx9/+WNl
AvwW2Ne/dgBkf4XClclAhLj5SIZJn8quARGfthmuGuu26wZf1szA8FkgHlv79OD+
szN3rN9tyAjq571VgpCM337q25/lC13lqgoqdjdn8twyGs0H+rW7mIMWxJcQuINU
yaN5V62gAPrlWmNLVDyQU5ffdQeIpIg4Jel8AVuDcpuq0CdTFaweuIESZv7KugXH
2KK+PopDSgY3W1cdDRMfTnenPzF4jzuGm82e+1ykjL3XHCPlI4tYLVZmZ+SvBmwu
txMcXyD2LzGQNXp0TmRea0sJK2x2ZWEKTZYFse0rz0IKe14+K9/MLOxFN7KjsX2t
LjzCweSygKznDVcauHv0s5Gtfv9Y11I4pjgakE41HMwcADkEhlfPX9YWOFoo/6be
w+tZmAR+GfkXw0yUP+K8/VxJYdw8t5lOEc62hfWMVII/hxpOgBtz1qJzrb4hGsjI
kJgLAJldA14jKzQc0p564LVjOeQat+8e58JhAdf/CH+Q8DyOTTZMNmgCLYO+afG3
j3pTzlWh7GFzSmAjkGQg5SZLMGa7dZ8TyvuXDr38u6nE19aW8tCXYTzN4IAHupOa
Uy4sDBm+nKqNVg4mi3mnvWBFA8Xz2nd8nFMdMTDYLYtoFHHjUBrFz8iVg2vuiBW3
6sfSb89hOuxHLaB78UMoZSlNqa/o+/Xqz+OTAu/dF1GrbwYdl1sfn6xjuDBo0ugp
3ewI9YCKebJtfrxkwSRXHHuekwLUgYzeMor0Nnfpzkx+ZMkPiuJjgk/E+Jx+q8MS
IMG2rKxYenZN89C4u3p8S3lY/mX8tzCz8Hk/7R6Lx2k1697YcdbBOpgRs8BIttZL
de8DR5/+JifU6c+9o9SCoIvo8Cg6noKhItNhfnNyJf06Pend6Y7lpYTMA6P5EgNj
n36hMBnokXNuzQZQutmWKqNdttYW+S90bTtGNK/IxWBqHG21WSlyyy1ArvpWviTr
yMH6gQSa5BDdfh0GShWBMQ3Hiihbl8SNd7mm+OCF9VBAnWLopp9YgjmiHFwPX8mE
mlqWl2CnF17wm2rDUcBXLAu14CkuA6bVp0G540XYMSCwx+lBO2YanthbJADX2QQv
7B4rky8eiH11eJoUFOw8a+jL2EBNFEDKk8vj0rH/GmsNOkiBb/GE5GEQOmIkATpS
UQ9b1rqAUGPFOfXEG6wTncJIZNUhCimY2N/Rmf2Zcok3zaCv/aHYZxSHpIMJ9jhd
D7veI8gvcapSYaizI5ZuYxYHlEi7Dpx6z404ihNjIOKueeLaqpmxioxv6So9METV
cDq6vKdwuUN0npfd0zRrnDFOmukNVV9pdVdi1Xk2UkM9uKUpOicnYuu7UGq3qlWi
GyKLpjco0Hyl6vlTevhevsHgTtfNIxwdgy7+7it39r8d65zwaa8d68dPxiRxvJ2h
FPP6rzHhOyVHEJFfRvwpWcuYbbhaMps8dAh0CMQJ+j1VfiOlnVAjXYnUIiPvD7ZC
5fcs9fZ1JGNttzJ3oc534NwfM+5OoDpGOPGe8iLXVoiUQ/5lNqiAlZNDb0EVYoGP
KJJsB6PV43Jhg0QmdWILd3PQ75MyKX609D7K/46J35PisuoEyGK6y/Z244LQPUJX
Ep6t0JS5vsTR68YoUVBvVYzSpDKp6N6evarEdTS3BD2xgfpA09WcAShF2bB+yvE/
4JKSCtWKTj2+r9//Q8QKazbkgXyXeAai7re7VWm54RCEZbpR/SidDG/fdcu89s+u
68vglP9KAffwBWVnJ5l7wjLXRCrpzmggwKGxfs3AcWRfb3psh871Hdanhd56LSi2
wbgSKGpvvtEjcmBi+Fge3e2gK65lOvKr6MlSd3L02dtnV4TO7SeVNtk2lJDSH2w6
co+gX7DBXNoagRhS/O3mjRokPChUQyKrQxnuS2HNPzTxNoNaIGpuBWCkiLvC0GBl
2/woK3o2XZX1+6O1nAmOsgzsouzEkI0SYtTz3mxbgAiFa06sYgtMiBAuTSflJMsj
AMlIinSbfHICoj8pFXgy5nchhkiT23PNMdUJZIP+3VAIra5PjmVe3wwbI8gXP08F
wVH4MTeozEq3wjrNYF9KIM4HDerJGcoZBmS4sHV9e79dARXprbW4A5jaiYyISySn
i4GAZU73+F8rfwHLGxnmz6ZxNgXztXUDRsBgolDsKZ1kbp6YkD8Y8Ip8olqAyDvm
PMmXHekaNzzBYb1gh7xpO+Ou+ahDBulpA1smTwzjW/mbIzQklULV34AgKu5rVlad
62PEfeqpLB0YQo+GIqXgme19mL+RaBnE2pEUJTzwHTSopR0Ny3qq1CR3GxsWHRaL
0Vzrj90ve5a/Lvr9FuJv6AaUiXzBK8ZDUDT1QSvwddMqs/4MSerJTDu5WCLiqFMG
45oY2Z5GGZLJG+cblh8Fy6GIbUHRcdmaT0mItjUJCzRBBcvlcMAO43mNRCZlCyrL
8M5bXUX7DkEePptO6X7tFD6u/gtpm5ZzhpkMfCVpj3v1gLf+uJWsiQ3GJJQup7LL
2LjSKqshZfPyrox3E4yWvyJUGcPxv6y5IU4bmwrUIp2vcn2urDopoXikGY5WtNCc
fr0sfsjBACCJn/Gx4jklSk//h9AAICaooG2ZheKctzvJQtgQuhNnWhQ8yyjAe2Ue
azMPhlaOR8Pqt+SQ7+biiftdRcmEM6LwxtZfTC9mijv2TFZKGcxJVs1Mmlg5sGfI
666j8WXCRV2hUlwH0I84Xn6lHXDyie4AySB7t4qIohZmOz80oxDuIRk3YQBazAd5
jDkoY0EiHBnrcltnrVU2JFCtYFyTWZv3PtPOb5DNJpCFiM4YmXtxHruyanT62NOr
OSCYLUywakZhJE9u0jdyfIbAsSEvKjVB3NNvHoKInGcYyQYhV855+gcJ8VOjRICC
FpPoC3x42ni891K5GnIguZovGzV23CQZAhXbRoYYnWuJvDORBHM3ECoR0ZnGNd2O
NBL2z96an4/pew+CFs/UNeVJ3XwftwImqkqrdG9Bez7L73KQedp/yp+XbRrxPWDL
QPcRqyGuu+EHQOhoMvrX77J9WKswqPuw+tA9j4llG6fSCIlyFmOXkRgaHiR4A/pw
Vj8bdu1F84z70r1LQkBv7hkN3wCkbeJwWpZcWir7MHfO4AFbaCG7Hl6qu+M0Z/iq
dgjpVhqXbISKsRmWa62WAIGvC1tTca6skxQpKTo7D4pi+k8HkOZb95wyDh4ysm/B
aeYQkNdoQNVKRcv2a99MFTJLcgqwz99z1EW12lCV4dABg+SM7ZqUlUYDNbjfOlFx
zp8atUMAjpvxmoOZsbOQWSq8E7wUy4/TOl6gG4qujxK/IIExQ+9l3pt6l7DsIfta
hEqJCFzJPosC59pMYzVoVnIpCSF83cvzEL/29UkiBarhm80IBlF1r9FxDxrVTmx8
J+RleVAhIa6iqpbmtblhsSU2S7fMNuyB5moVBD0LkTlVlX8cc/a3/Ft/5wrw13A2
8C/y5XDO8TLwkPgYyI3Tb0gdKSREbJcDYVtM61mXVJE2KCd2YXlHhZkB3laIHwoV
azG+NIrqULwhSyUSo/Q7czgonTZJ+oI9qJk5baG4T421ryQ7DiOSTPj394fY6PGH
bIwwJYF05PO1MO4oibBTpkcpPQAoUJgQPY+4KZKTJ4LZgkXgFGofUWdN0rK9xIss
zV9CxNANgUoajy8eayghvfCkINC+iI1uSjmp1u3T0i7+gtC9vAZu5GqNl4CwXHvz
0i0Gz5SoSooiwAG5ivXn0PmEh1bXWjAI/DNQ7GDBNpqz4KUISw1VICZR8FC3+nXR
jMR3bF5U+cNSu6q4CF7EaMM9Tb8GHQlpp84qAAawv8w/pskIeeAGKFdY/qBJOgIC
nwE3e7xBrw3M90e7oFCHpGXzhm2fs5dt8QG9PBxbQA93rjs8ExVchnwlnBzBeULd
RhyD/AcUgcqvqIC2Fu0onmhmbrppmFCmx1Rd9dH2fGKCmWeM/d6nJ59zHBCBr93W
+ZApDbppXXlM6s6zLBh5k9b97UP+ibI3llnmOTeHqQupgcKFnXud8qGTgrhJbsMs
QhMslOCehxQCQ0wp5f/g9oqAQSnWkNHYnOAzqvLHWIt4tzD1TEMwGe7d+EAeaKE4
jeR8V1q8ud1QtZ82iy7lMNWr6wrym9+fxEWzxygpVSak3y/17h3puAGNg1ceD3kY
sxvOJp1tRk8BJQgkt4BxHbDPWTWltx9yIo3RZV4DWA4heKT+wkNkgIh5CJvx2lOG
VCo6/jjmyXuAOTKU/LOcaYMYO+wS2Cpy14iZ2nSXbvNUypRw/oPOfvFCyMn6wSCg
OVcnF5CqfOsZBGAVWf/fCrLrhaP8RlFIHkd95dWPn6k9KzakNySW4udOfq4PUxYb
HSyAV9k9AnL12I5P14DlnIRKFfmQJ7nRBQTlvBJfJ/td1TmIEkPJmD3yC3tHnH7l
hBj4DvyywBQisC2k8Okw0GzT7tZOecMKR7C1v07NqVmK65quCB0H9K9zESPTj9+x
zGs2zdc8dg0sEiOtebHePGWIhVr0QtrgMJi1p6DE7HWL2vfsb7+yrFCUKSlNX6Uu
fml6MAJ7TeUbSZcsjUHX6Fgyaz/sJ9ZIK/rixDZmWadhEfP/3FQ9Xd9jGzEzbp5d
elA+HeeN+b+o0pwW6zEGB91v5s8a353gm6VM4JykX9pihd6ITWRp5wAEPvSabjZ1
N96ytsNT83u9coPClN/GZO2xq780LRRW7h8IlrEYqTpglqlcCnNghn6sQfzlw/an
IMBA3GcZRHz29d09Ael05wdDfwJuAwJAH524r8kU/5UPqzyAOQPmR3dC8GOiix6I
7lyKVmXzDnHAFgc4s/+JGY0xmXWg2zQp7JPe4l/km2i4JDY1xH3bBCaXjom5yBJS
b1r/p4zFpfDYPrKWWsTJISuCRZWu8rSmO2JC4YaQYeZkxXmOvbkLw4ZD2YJlsnPj
gGeulPHBEdntSaC4oCuTSZSIx1vr/+MXhNLIX6nmInFhQeyG1YOh7R+h8u0IdLmz
YF6y1fLbdwPxtJSsp0m4ZWvHgmYXBIDFjjZSs1Ipxu2/kZBSRkkRAE+K5bUks8Bi
LxIs6QeJAnR3FG+yO1q+Up1qmf1/shLchuPjkPSsZJi/+YaYtqaN/RK+BSEWdbBo
YQZ0IQhwUS6Qe8gEzuOUMHmDneiztwkJ+RJjOal8ylDtrEqzA89VtQ5NJBda3/04
pHyGb0X1rzk1aM4cJiFaG0V5yICWFR0alrHYDF1+w+Rd3PCGFwmcZWG+XMdx13Cu
vzvK0Aiftr3DB75IMgBzBGiYpwKrPARoxuwjx3aVA85SUR6uudBpgS3xpAxbRDNu
XMGPA53h7vyy7akoXkARGmSwSJe+zLZXwX71JWIOcCHhQqLAyg+00+wmy2NQUzB+
zmOcnOLEwmYAqRN/Z+QB4JWIMOaFRaJ4f/FOmIJHgXVvVmeoUY/ejBpvszmIiz05
Vib6AAkdRxDjusOxSO5TGZCByQ4TC7aykQ3Rn2L6gh4/pq57AMp+cU+/C2BEKpPR
yu3tsyDtK2p5+BCYPBGBCYOToJhZASFc+aY2kpbtirmeFHsuZODgxjyX5Drn//x+
MGjmJjEs27XUt95iGq0vKomXclfOUQVvYU5oXvQeS2vR5hydJcrXzPxW++5VVt4P
/DoaMQO0n5eLs7/6Asje+VTPH/h4CIu3P3oySh3iJxyPKu/5E9T/ZO/dDduBQW8W
VfREymDAAvGB8MaWV0QrnjygOoKrXFli9yUYy5xIY3HiT0fHNkZHE8/nN7Xl4gwP
M6/gvsO0PBarflBzUGzbVayatS4ZUUndDDa4bLJCN9hFeolYuh3Yui4ihSy2mz0r
a86hFdoW/GqX6J88jhi+v61PmySl2AzScsI/vP5hhZGB/2EU1/g9H5IA0aHjRxqF
6cJ6/dDaSBr4dQIqmy0JCYEK9CTjsnBcgRQub3fCa6piyRdCwe9r2wnhQbqXHPna
4REPgfwuWSJ9EYle+sxMX4zfE6lLMsCR29sVBf09m5SakuDSv0aduYHau+7U4VRy
bkQi/q8HyLUiNK/pFnyF/MA3UN3c/8Fml7a6/SLHZLHNHrGpApWsFXsRo2PX7OBK
ROu/MlAaFuCSrae3AmbwBbcUvnrkSJCZlofF9PKSH34lQNQZ8EpvU32yKjBGDRua
ztRNXkSKG6t3+diZJpqq8kFjTPqTLOvVOKSBW0X8Tkn9Jr87JSDIFF4iX0kf5+VX
8RepJlJ6bXTfcLdZLzO6phhi3suqXPpTEcgW2gXLS6er0IrC2wjXVbY1fSU9JUWZ
no0BNPM+Ny9zQTb4mE7Tm3xWWucB21HFncGnqff3FzqDfQKSvVM6kdISTcgkkaNJ
onV18dRgnH8WppaWwmQDN9IhOIBSYDAXK2KSTZWUQXXL9XcNIFNDNxrNtblxCVBX
woSwyiujzTH/jtDtzpJHw4v/+Gzwc2zm4RTWF+WLSqM/7kwbDeRepSF45a3iIZLu
jm0OOhXKlsT8xlkqOOhgcAdvtlqKl7/Tq2iOkLiWFvnyejp/wPJyzP0NO6Heti2F
6u/C01r/R860FwnbPsKMKl7RZvDMoYGTtk9sKQAUOgBEGh03Y1oycoy7MmOC1OkI
TEVAa1/X4BQ16IfgR8LHczfpKfqOlhti1yPj+pe2f2bHKtc9ZM5KaISIyRPqqPb0
w1SBXZw5vD3ZcG/pnZPIlpPZ22ESXwFYa85BxJ9kWyD8mlIqO34g3HsAl8sRxf/O
k/RpzmL3+YRLVknh1OWYC7F6W9/bYXL011PJ5zepKnUp8X9FzAP9kSR0baQZX2Ir
jQfxdGTkH42mISj2cEDT6wp7f/4XVDLYaf7JT8Usst9ZAFFYixITbuHvYT6D+mQU
bti88+FXUiD93Of1NxQMTTxBi7/Z5NxeMTdjMz7NxYxpKHBZ9o4FLrbfY+iVNqd1
AEMNqNSXZ2brwKzMf5TVIdL19wAgR3Dwui/Wp8LtT0rXe7XkdGm0Id7umNM791Xo
jCaUoHXULtNK/cMXjPDDUWk/egssuvDjJFmsRoiaIao5Kg+SdIiQKEJTPLOkqzra
CGsbwrPd4PKf3OrwSTeezJ750oM0f9pyZVQ6hTTqr88XlyWBtnTqgGr7nISyrBBk
aQsXVP5yI3kejiAw94MgjQ/vEtvri/gqWCqaylRUVRNlZW4CVnVfnQ4dQQZrodBd
xC/BF43gjCFNQ0ERRB9X7QwezwRR3PrdNsM0eFatGpTlpxU3RZz9VzEkmULmAD35
tnLFVP7sQih0w5qMx9pnxrsiGUblAYWRuHndIxl1dgLFIGEntLeZ3zVmHo/TQosZ
oIxUtcJFLnKWuhvo5nuL19MLr+AM7QLthSwIpXONbazNsPa4nv29WEOKU/jWlfGD
inv5pUrMeTu5bZLo3U4tvgnYxYhJwZwyzfRQ//LKmZ6r8diBvwFCx5lArjTeVfCm
qN22IARfpX0d62WdfBwf4Hbm7KXI+Yg2vZsWgPrILA61+b3jitp6pvHZQnhTeNVo
u0FPYmJq5EOSQgcnHkSXuvgmUGWqKImR+UW0tN92r36TOQD/ElzlaBEIJFCOduMO
Rt+cKoQyBPT+8dzIdaQPNCiL0GVo/HQ+/k0erIV+qHFu5nGnnfL3H8r2Htt3rZW6
Ipi62XGvJL6EDRu/e4dmXPY1fWi19Ejugay5yF5QdUWthcqDN8lzZyWCrgnnj6L8
dSxViFcnYwA9Mv7A2BpHxspBbbDVPjMQT6WSeRYIc1t3CrwUBmECzRP+wYPBunEP
cYtD1emxc6cJayLiFiIAsiyVrQbEkkfiLyY+UUQhdVabAV5WlB+JhtORd7xxL10d
7cOoyD2dAmW5WqBIaA9XqoGTl1REI1ZqN3o39ttg33aSDAd3VW2omV41q9JKft3t
+VbYhJzXNbSN0fd1yLaeBovKToDN2rKlIsUwhKmaFd90AasRWtDXPyEnTIUYnvLI
WvxOcc8dPSEc5uZ9LNOY47KdSEL5k1tXWcFUA6YDrw3tCFqQZ/1cEd3VVEoP8Qxv
/PJ0Mmgy2abUSM26ZZrN0thjN3EwpWATqexmcdC+xfLCWCMUIR1B8g1eKxr3dSR8
RrFEOhxik9eJMVJG8QrmlPFrEeczQmcg8WkbiWBHX0fsGi4XYKpJrLBQTPjdSMQC
GUO3rJuZuMuSJ9eTtJtBtWgjAdRDHCxlW4WG4wz7tf/7HcsvWiEi0X4N4C+AEITk
WR/q8OTNyLCbNROsvH39bZej/LnZgsS+JLIkp4tu+dU+5jRKo5nnS7UNpvhpGnWk
XV7S8sxexfXAjJwCoP0k03NNlYxPL+b4wef3ttbYy8PauNWTk4ikspW1nlIOPoCL
OeRqoTKV7BtCD6Zgbeo5ZEpAlG0aGdNqETBsuw4cHTXjxritauxOKM/e/f2odZgb
hiddHcqVVLIZJpdywl7Gaz//rqn+52g5xTodNkUjwEjheRlpB52MUtJIn23/kE9K
FQLNMY5YXb7aRmOKeWOy1CuZdZLQzW95rehti2Q0rJtYQbZ9CqFilzBpHuJJUq9o
Lf1gj8aK2o2mCljYipYbBEpvgDAaD2UYQTX+h2IOAOmR1GgB1/Qk4nC5fR2GriTB
hr9TyjHznwZlakW5zFM4fhjzacxCXhxszpcJhbvJ0btNMTKKOzqpqCImhOsqYa3Q
s7KF+1zNKCbF1lnYjGRW0ZePCa0MMx0U+3IVGbKrax3hgdWkSeRZNrVmYb1bqZCw
a0Jr+xGG/YxZ+eXt3k8fFP+ujNRt/M/jZNHBybLTC/V497OgNqYQ+HWeUTizKswA
OhDKO7rNFItFjlW5cjngBfv15nh7vg/LKfUGWUUjms5ChzgesHbYnm0lrqj+csk2
D7XVWCV1FsUQk2jQ5/qs9t2M+59avbjVOMJ/+7CdurSOH+gwzMg8xRkDboQq5VRi
s5VQBXAtxuoNVclfz+uLaoL7OFSjC+fyk/TN3hN8fkBIGyxW2wNof8A8Kzsej214
liVx+ExcsXSdw4Ws8UyNmbQTYbuKycFLNRVWavxG3TjbtZgdY/0tg7Iypt/TuP0W
JUcJiCu+dXO02+EfzvdpCgh/fvbYsKMwv/GCasM+2ASAcZNKXdTIO1pd6tKVJVuU
lVO/mW1/3D03SYuuKPwQWX8LTn9ylztES5bHHU4WaYkZylSbTmIb5A+53Fwb0Wmm
2jEHpKB6KxyMMHFwuSlPCfQnHWzuwTar5rUGQ5vEPbwjfu0w5riGaiglhRg4QJad
3hNCaLDyeT6WpHBZUw38eQqYCCbhyPOlglepvibmey1lV49JD/lWLCnnI5b2BGvW
0YPNpix0oJiqp0c7jNuN9B0iDUqLX9fmiWg/7vFhUKRJD/q8fv16vZFoqU91FjTT
NjbDPVo6S5nxIiV4l3982LDSH3g35Hnz63OaJOSrOvel+ol6Jcq223Oyjbudj4Pa
IxQ45TjcB203YkroqLjSwOQ6aL3ZskXLdzC8AfbTtJfOoi6yWgS8yEaMsCeFPScu
1NPjunfxV2ySsQqtnv1F9QBmoVJ1oU/u3Pw26TO4Iw01nYEOsmPijyCGscYY+k70
H5x2uuadZE0vP5YPpiM1i2M4EttQzCNhg/wXGYRBw4rkB/vPsnnGfpBz4/kO608m
KZFD9z2hHbnjT3CJSwCrzVbCdbbGaiUX+apD9BiXoQVV889J4d7KDZMixeWSQDt2
T+JbOPC8EaRJZhFXktiywyUfxfWExQi/xodL+KdWfw/dIwf16fZw+YZVOtvsaney
rb7SVHSLp81XsAvxnqVObkmPT3FzH0VgXPyHgAB7CN+D5C/sVJz3eurt+4S20TBP
0HByK7qMhvSZoIuAcOVL1jR06IWxvL27cLcNnHDNLrVo/0b+cbJ35g8kZ8OcoaON
SBHmIuKWvZYMW2q0IsRIOOJfXIzPx+WRHEpOJlCNPEfNiFaZrUmpJMnKddQAFWtC
EjIrO9RTxUP7f/riYzgw3u60XelHXn8n95H2Lhgyf+M/lkd6pF0/UoJdQshWPeQQ
Hn84b4pVSQ0AEhMgU3PoIvnAtzpaVzeeuqwDjWPTWGMShQdg5M9OmFd5Xue3ZfL1
gc+dDpa5ngl9Q/nuDWpI6wGMb9P8KzfTbPtO9W8cnGVTiG99QfiT7tUbpFZZXz+H
wmKroKpMdMUqkr8E+v+Cw1jyqYSBi846aIFXV/2Jdk/lxPu3yRXYLoDVj+VkMygD
31WWSmxK+jcyCF8NKqzNs9gmgfaRfmlBBfomh5XB2Pclmg25NrmxRen6+1jddzJl
IDEW9VeXpTK9s+eva5XvKbAu1g3mTNKIgPFtxqpe8zc9+6WBKE+o9Nth2wv6cep2
PmifNk5ZzpkCWtNSUp+s9xwNfWUcJIuzONZH9O1igVomOpFD5+lmFl0pb1EQHSId
560/nyQWJ/HU7a2qI96OUcYPdJ25P5bCEQxqnFX4binq5mEYmQiJCoXyBTiS9C8s
3685vaNavdwZKZY7W08CTAwelJKhaQlw0ajNQ9pYJ2S+PRZdmQWgz+GjG6lKz9be
zcgOkfSWGuPqN1f0k+xdwHVkZVN9xeJ9SwTKMI7geRhzO2xMxY9rzapDQikUFmc3
n6wtJmlGc1OUodJoYb7slOBs0vDKM+sNojJnp82dhjixkN+Xfh6FFoqpHRd+BqnZ
he++MHBcV9R1ejA1Z1rh8TZ82RQyCngIBKZ3eN0t7ATa9/Vl3KPnjVRIoMGZeRP2
dXAjUz0s89CQJsw3Hw/heFMaSqFqFivaFQ0eqTwx/bihG2JNiiPyh7P61Y4O2kcE
SjUQgeW5cqp/j9NWMyQ27lMH8nHI5sU+dbprATdBdpHqPNCNhZRaEPoEP369FrW/
v5YF5K+14oyhZl5266VPhpVrh679cWmeaPrj79RgjCDsRy836yZh1658kLwLG0VO
Mwvvmbh68k9vZd4wsfs964yUC16k6x+33jCkF7i/CE5W1uZKSNloIdsVZNo2PsUL
bQ/NXULuOxGiYC3Ysc/mw4ynbftAp5HldXkxuVOMSY15uKtncjY4JtrqOjvIJSFN
Z5CjIrf2Cus610E7M6MIOLtWLfZBL+of9lDuAzeJUPy3YDkNfwbmlyU+BKSFIIFD
krCWSODYQDCZrttWcyfMxPYdqdN1J+0YOzaNzRJlvihxDvXulrQ2oXImWMW8LZrO
8sF20EZvtXDGsMn/UrF9tzH4My3n99tfg6AM4QpBrx6fQfGWatxFALIlGu9kZOP5
Nb59nlKVAWq6rIdZeOSbjgsucWfo3R9dX0b2+Dg4c3qhFdMHmTVnzF8H+8gEHL73
dWEnDLhFO3trbfmVuM4q4JXzOOeXVsLdxmangiVVQgjjmAH2TIU2X7W2IHMmjg1W
JZ9zdVDRFQs3GYoT1kmrh0AUScyG5hO1r9WHY4jCQiIU91VB/alEVzdEjW9k1Pfu
qyfFpdoSuu1NcLRjbVpetXXz/2DXn3Y6c69pON2v6sliJMhQ7ZZRZflQfy3Ya+5P
WGr0WJwaBnXvGnoFnH0ejzrblcLBDIqt4H8rfYgyVqi/H/d968Iz7pkeXZBdg76Z
Krks2G6qw+nAiP45q+5yWxCas01aJJqcuWt59vQEA1LOjF7UGefDPz98SRQI43q2
EoNf6wgxU8YDPOZe/5/8f9K+Vo7/eWqGMiFi3P1fmzY0HHWWO8xZNV/XYFsjSw3k
zHjQ+A6EmSvedqSpGL6vdlJDzVQWxC3MXhkcHt5im+TmOQxztK0SKLpgSt3rY3s+
7y6HD/2rk9OoyaeSgHUC+YqSCyTAT7Df/0Y56mQLqpnaPJq+00JMOHve4f33uniF
me6T7De52fv6FOFZsFXXQjF40XcBdQFyQKWOlse/hIj8iBKSPndI0GKDZCpT+ZRy
8cLaptSdQRp6vKeAJT4DPDxK/Avgn6oZXtzl3tEKPu/LK3uy113ZATsxqHrYyeV8
84OP0M6fYaNFmCVfqS8HszO9VhMWIWjV/+x+C8N6/jLHi6o6X/+BlbanLsk3p7wc
1tV+fjKqXQRL2PVqWLdjWQOFgzZvVnpLolgBasHS0Y4L4FE09OGTVyKNMCMCxKre
kLXF9c0fvpEDiMldT9BPqENrxQrU8ML5e1BWWiarGwYu5Az7w4hQa/mmAw1eahLX
7nTag2PTIUCGu2RhNQwqnIFTdTaKIw9Gqfb8+NXhH6eEXApAuiKdkV9+IZeG+yDX
GM7oIXrfJDdcuOhmyELRh5nd6RGTEFM20WwaG6vLssFfWrSIt8RoIqme/seNPzpR
qDE9HomI5UVXQFni6JXB0cyVExd6glidC/IQ7B8FHNeWFcz8n2ShY+zWIp4Cijga
UYHJGRPu2zUNvla0d3EmFFjDtwE3+065D6TtJcVVG8JHZ7UrDjJ4ll4wehDwCQP3
NhVVWEfPg00YdGwpHM7Aww5Ip3WoKl2QnJ76oL41gpINTgX157URvA00PDatyygq
m73Jas0eel21CPR/reqWSOdnpY6xtSwwqFBwZlFoSbq04j7wZnuBZYeGY33DPip+
dY4JumWeAXhKv4L4f8kACoIOMk7VIvAX3FmkFZXCxeX73zVaweJEEdoW1ZuWsE7E
SJSppTNBWCX/Q83wrxpvwl6Zrjf2YmECB8eGAdqvKBgW0MLY/9QeI/dex0kQfnic
jYhz+vd4SiOMxmoyX/fFtH1t0sDGwcr8/gmJPoq8y04MMj5cyUptLZwNdmK/a5jT
t0YdxQ8kVjcq/qzJ9xnVrFoVqS7l3MFd1eI2xZWTjnW55Zt93U/aHIg9lTexCUAI
m+FGDSqZ6aZUXzdaHpRXy/sha+dif6c+BkSVTZlXt6eGpf3GYMzpgcXKldL9e0V5
SIkJKjbOHZQ0+KS2dhaBRVyWaOApN9SZX+BTgIbDACHJbzncfPaKG3qsEwpDnYlJ
ftZ9rXzEA8RGyJsaH9/hJLXI7tPcEncFEHO5WTSm4MJRKn7Mzwzg0BVejLHNN4yP
b9omrcCmBmjEUJ3INYLKbQPuV8O+Xgpeqpa6Xs4syY1ZRJLNvBEeoQQLV91xpYgm
+qphtn6Ho/PuNGdgspSJECpizYhv8NVqWuQXBVWFs1Ialjquww/1LlGWM1sopMaW
XwzPHucvZbK97mrHl9jOnB3MDX+grqogSkObajMeREBG0S3yfJzFqkY4hssFbsA7
I8fJXstiUretUZe6PDdNcdXXRxYV4woMDie62hAQeGaxjHjuFTE/DnVxS7owRfX0
fkKLtpSR5NEsdG9RYwDXnGeWeP1ky4f/Xxm+Uc+bQpkpS7TsyR2gWKFvx4wvuWw4
Q2sZaAh7MhxUbxiiNW4+og2zgVUtq0hp6uSHUHV0whIdguEoZcbm+FY08DAGuiNn
mqeEGUlERQhxvvd3e0Z9LwqFiA0XFQbJguLPhWWwP7VzjlSJeS6jGq9YDYg6W/aa
lPMdY3iL3SG5RkKtjtXpwSwAp5vuY4PqRBxxqPUXwYOhp9VTtu/3WG0jomZ3spg7
e5dHwRs0ky9ue5rgbIlClRGd8RK3T3LR8gPw6/9asthcfIQfCKuZEAe0uS/wqaQt
udt8Vkq93Y4+xyhGQsLKSACKhPTOS1gZThIFpkERlH3v/7JeCDjwpUysvp4YDMnC
Jb9KGlnq17/sRTWC0PFKkrWc0D0ElvsGlDyGayeogxE8nA9MqSm5Lm1ofposrUAW
RVX0ToeUU2eCE24b/l3+IzsfNdlkWi5Z+BmDWzqXbfemjcKpbUrotIWTNUxBR17W
j31Tn2tl54haPIUnne2LLN0Yl5W2nEYRYgQuzEA/+vakVkxgBG5XQaIUpb2fKQ9V
Z/fY4halCk7/F4Gwhd0Y0qRWukjXPNzV4U8e6Ojt433q3Rm5riohAt02dXqHBM1g
wYIcpu92QmRoGHTmVLA0fcwAJWHxkXg7TCLqaHlRQhRMg4uPG93z9BkQpzZqbzHv
0isra2WxHV8l3+UenuFM2/hLML4unoV8C9QlAYFfy61mbXJOHV7x9Bx6MI95pxLI
vtpOZXJDZPLmRlBbT+95FV6YYAj38bIqhpqnPQLqaXRrsNn6+RBXOIH5LZS7VUhm
y0cruuueMoq0g2IbGOCtnfa02Y931GN+hC949FtwodwQvpTJ3aSJSYxFoZmF3ORu
myFA2LqSWyiLAqcL/LPKZYHwCbXW/jJfaH/DWs5eJq6p7X1s8sBWmKjwj8UpElea
XiTpNonQZXU2uHXCIlSKWAkauWDoJKybqXqGNZYdWlXZe5SQml1FLgcq/84jhWdZ
BYZcr5BeTo5PXFsGRTxe09S532yiD/AgRVGsPwS6TCH3ZiruU5lOoHNBecdW1rhE
pFOrnPL+JjRDxcjI31IMDBar0nNqIMgpaJWHIL6LbImfgLBgdEeCC6JxcZUgVMcM
K2h/Dqzd+ogTxIhtFOp6bJn7K5SwH96PAhnK3IeIgfqnZfTjBngZ3XA4+HskAIOK
IB1QQ/4KtrUoedu/0MnouTD5/xCzoKByT/QRbPz/7S1+QKAUsYWyZy0FzlDBZvaM
X0ZRRFI75dd8dY85iKj7+WTKgz1Vc2cJmZ4IdAtZO4wjej38iNn7e7PhT21zsK51
VhhuwtuZUb4g2iFkAye5VPcl3XDNWKxE2x4cFxYAwYkNpkprHvWJ7W1SShxyLYee
FPnbvyCrwnwRAuCUIoS/GKoTm9WenkRjI8A2/PuYSFe8WB/tAYmELJL9gj3xIO5H
EQZUn6Je8HMbP+tVFgS8P1nEhsCa+FPqzaEwwCv8YZ5Fky4sx7PLyDJyz9ROZ8Gz
poCMEeb34jNzT0ia0AS0Z60IZqhJ3jBU0yzYu9A3LcLL3e9sjER+TVEU+ddVfdKG
Ij9I9WBRvz/maW7G9P/ZdWSOaN21TvJyK8CZ5K8uaNU4/DOGL8vksb14tPtDTVK5
3+YTEIgCqoFvcgS0CsawwYKElHfKMPM78XzaKCMu6pruHs4s9H2j50t3JGsX1BVp
w5BSMJOGJNKIeZMA9ZPEE5iZQNUSz/HIxeaDOL+646V3Fh/l/Zt8KU23extWdsFW
xv2cJYgd0AtZNmSswoHi0SRG6p2Xc6o9h72c4XQy4FxZSzO0V066rW8ITRVgHrCH
x/itSAxT+8+N3/L94P13lTa5vqaXoRqvmks7Bbf8sGCaphXDGRZ3asvhA3vXNyjr
PixnKsTKQzTszIO5K971rNquwlK8kMrO3maieMzYHndSQOqhbvIBvCkfnXCLBL/M
LXIjxhJ+buwwBYfPVHWevnk+KwXPj5yeIsDE8Aj12skuiU/ZRfuZsojOoT6mX6pL
XyUKaNRYHeJUgk9URAu2xjCA1mKPxir7YkAeWL/7SzLaiBbtApSC2kDmvJ4gi+7B
NLSRRcN29s0Ydwf03qhglGATqvrg1jxmLfmCypMUGN4JflpDKiWa8B5P2y/hDsZ/
MKkDAa4/jn+3zCGIApduYlOLXbDkiyECHSQMWFsqVIDuUBAnPvYWM44fjK0e6HPk
RCeOOgcA8gMDRdE4aRkG+fglxv5wskcmJVeOHSd7Csx36QGXb+lJeqVJ1hX8kLer
LaByCCmUOxMnFposTrdNvxzbbB7BSDFybf/2ZoHIEIa/MZY7M3hsED3ngry4dRTY
/6Ob1e1gAnuECy7tmBp1RGuCEZ8A4/zk10zL8lq65z3W3aiwgzsGr9U8gKpRIN9q
uYLvsup9PVrIs2SBegeTBDU9M/H4GFKR4Qb2KxiYgpxubRhb3vyTF0XiWeOo8lKF
Z+sxiWeNR5LlY0pdsaiS78eIuzUW3JK6G89p06cjxOhQDbEh/hAV3hXDpZgE3JuL
Hv1x6j91ka02n786PRRYRg5FJn8rJzdZyxr0mZB0qYIBkXdUcgB9T5P0e0Ypxpsp
DkAT2YOLt12nj1hksTHPc8tX5YmKxZNFUA73LJFV4Ss1/u1UO4VGtrvGPch7a6UL
SFJNs2wZ+Oe4Pwrtw7SgXMGt3lNgOpT2agHCwPmkVoJuUK3i2nI7kWWvz21roR8A
HcIz7OnqjOHbP1BVEssyHl3aerjKZxQfEvEGxd9R4/9UKM4zLSEkOOaTLtyWFdCz
szJPI/PzGrw2hw31SpTizfwgALxf3E8b1vJDd3a/4GZZQ/Y/VluLhRzxeXSIhBVY
+Tv7vIou5c3V8YeRe400sZS5e7OqwWwrqmOXc04DEIAFLSXEK739dlmdPDsMq6lx
usDp2VA7TsH/44JgCQIB3I7M4QZExxGF3WEKmd9FhnKuPoWNyZIseI6+HWuaWoOe
H35GAe+BHrpCqqhbIbyR6mrDQQf/NnXWK/ivL3uhBdLXdCKesHEBQ0xmlFv7H55a
WzxtQrGjwzJQdEOX987YgU9CdksGuR6/YLJIk3rYt4JrMHReCEIPdcZFRyofOknG
/9wCat3AFeheDpGR4M0jYMilWfOIQq/sjPJ9kLjWKyo2Qy5HDHowBRpnW2btISaz
UD9j0z5FqFBHIrF8sNWOU337z7qovzSpna6qI8uxHvQq9KC16GBH2QnjNyDdxQEQ
OhQjSPZmByFLcvE3evJE0jTIJqKV8kv5XQk/PZyg/twuwfzzFlpewSBbcNLlUgCN
QnDPFQxwNgKbQgKq6sUKE5NOZfKwQegG+ilzySV/iknjEkg0Tlk0EZrgQrsbSeep
I5UY7mktNJrsQcBqHT6PRMrPW88zvf5SvVPXYCVTnl1jBRKqACP3VkKJQ8Dd/FPa
ZVfvoVRqLZ32kFE8FfYNlUnHxGyiQJQtaQIGYseC6gddvF5SzUCPtkTd81wP+u/6
S/Nv5GjAtPu1anoLOzGfh9s4a+NjV2NTC1Dxfm4FidPd2J235kU6uccBRc46S77g
IdtpLyTeO7pVl8oAABa2rqlRefSFN3medHKTYv6YnCxPzzeJhmuggOfd5nSsQLkX
fitKLF29cTFet+JqrE/VMyGWkeog4D9iXK8HH5EAMBsNyjVHHO057VrA374rFPIX
rwpkmOk8M7yATitNgwkb6959vOjc5zecLW4BJVrx3zQ+thrUkbaDYu755JGiDgnc
f/jAaGoef3+SMndTZS/6k0XSbkRl2h+JgLnO59LGv1iJbO2qPbl8zTuSp99ph3xA
zuuwvgjmEn1SM5y3ZndXBOrRE/goHsSkQFcHIcPVLfbeT3a1G+rkLteFikPqVekf
FNEMejYa34m70JF3U37F/3K5Y5uy0LUigBji/lR+hg3tZA8wr9yi2d10qJxYWJsM
JcE4O5opfB+pQq3upEFWeeXNqfG+4lVEU0WeAl5bpw35xegwB3xI1vGx382U3ugQ
d3FabcfYBEGWP7ijc6HBf/O3GQ6L72O7e5E+9W/RJvnQNdOAPARxWQl1WCY4jOsf
6qJGBTy0Q4I5EvYOiFhGrPduEaRvUc+brLsvmrF6Jx+V7Y+2aZy7ogcPN2F4G3QW
0st+aqEbI+8Ll5Zv1zq5wezC0pG50AJ66ZfIqAphd5IOpnUgp6jco1olSovctgrC
WMQtEcWFFrEA5dQSFmfLCuYmv2a921hzivp7sXDEnBuYhB2W1K4n4mIO2k5z35VA
okNlZQxXBE2duJYSemOo22JltTbuqP3/JBL8xvMPgKvtuH/IeGbF7bNg25dS0Qit
Z1CrU8AHY4IvTK0VY1UnKo6OUVyg3D+dUZ6XiMGoyxRIn/4FJgmQESZWqjfY+2dx
xeJp79u/SUUCh+QQZFbBgCOpeMpc9lYbwEBwsgrV8qCPSncPke+YKEztN4fAlVtO
MO4QbFTJkmtT8IOvoee6Q+bG4+ncXz9yHHQZbHD1+9D8RTkabQttUo0LR5JYe4GM
/gi471K02dB1YIs2xCp73UN7msZfPhDsafMCBVvu62WkNBRVGl+wfIho7ag77C7S
1qw9os1jv8weCd/k3hYIRw01fIvDeuDnEIkXF6Uq6mDHxhJjIZFAKYAuoE0xy8O8
WYMxs4vnwb7XVlb9iQp5av8UabXcFKmlwcG75qA09TncgpIQZEWcguoqMEVTJebA
madhn8owe+Ofpdo90U4iDqLjgzEgu3RfuHo2bqBtr4Id4NVZ8UeIFkZ1zh8QWDe0
qn+9ABTjo0CRT4k0JydAbVCi9br4JJSUXyI1yZcMGybMTSraOgG75DBMGoTT/vQz
GYehLfgOfRRzGc9nezTdghiLqcCBxIq0IhViGHCjCOL5KteLckc7LiIj8fNFypc3
ZpkR7jo0gX5F99G8UJa26MBw76LqcmpyO2MbSOfkGKvZFypsGC6ClsvH26qGZj1h
1Yedy/tLILcMI4XsVRuPei2/ks62gLysE64DqquSX5ZMkPa1lihVX8Rrm2FvqFO6
fsf/4gGiMfVYTI3zJZgInoLrhBF5upM4KsXYUnHZQyY8CCxfv27IRGCNBSpSU1ZN
dAkM0WPY23Lo/YVu2ae8MTkNztBh7gG4XnZkyPQ9c5AhKAShJlUcdFy2+xcXj9Li
cudEZJZGRW+gqVxLF0cYTBGjaHawnRCFmXQEsZCe/DtOkFZ8E48MQuVNHLRrRL+J
f74vGek1btyAxu4x8XHKOEIZLBUXmyKPqT27x246aRCM44zRD0ObqXNpaznqM6Hl
mOQLp7qfltgjwqt4ERKFYwcFOn8QaOgBlZC2XECOcXFmyqwAwUN13Gc49tS0F/1E
q9Au2dbtjngTd2RCBlwAhOCsF9f4k7EHmnno5Ce8C14JuKm7TKLKec+A50XMXrNC
24ZQ3X8Tcx8nWjTTwT0SQe2zKbeYmIngfEXFnCORrPzf0adzjM74E6CYuj1mluaI
u/gyLDbGY6W76gd0HBS2dsApFYX+zTj3tEI60+fD8wR4QbAJuqtQTZCILnomtHwu
3E/oWkW7AsiQ2vWvRv93PcDHhPuZPWOZcKW4DC1XIayiDT2jRt+KNjYp2C4LeRJm
2lmD50Fjo46fIhzpTH3av9ekTRckCBI3OfE65usCyezRKp97A3DGKyXxNQ9fgRR+
21b7bIuII4UejhWz4MLRXEeO6wua+UKn2LE8B73T80DCXd0cJM4uNh6BYdhHA/jd
GcROYozPYXWJt56jpRzUdcRLR2/2IEu3KRzcMubJagr5uUFtYb2dAtt2W3cOo7MG
me9RUKyayqCqWcZMYm2m6NghujOR4nTyg5VixcVmci7CxW7L+4uIc00yJQzRzNCR
vlM2+Jvqb9AfW00ZIj9qFqfUS6LdBW9j/En8KEuIEu3IKBM7ANGJNJDnBDCJVdH3
m14qVobT5g9iZSiGJTFh1kNhcef0Ccjw9t30Sdj3KXPksI1MxSTKh6HqUx/WD95m
ANsJfU2VTIDW+Dp7rZLSMJ3XRi1E5+FoJXsEifSe5CMzwGjvR0Xj4nNFoJCbAePe
Zbtf/ATZMWctqBu9FbZn6jJMxqQrC8+ok41ozDAlnIEL6NT3GLXYedR+Wm831Jeg
zj7T1qHxKpaRVFvs1ZDDs0zBPTM7kVWCJXDiRnxsSxdYwBm2JFhsbLDzPdTpIXn1
caTaYbTancf2Och3BIYeVVDh8uVNeKMsdVnrTdyR/jRY7P7ek4+yKgdKiqcVhSum
8loJPyy4NwLKfklNmWpwRN9e40dSOnyV0kU1LbO+wjoDvWNWo83gfsEtf9j/uemL
ZWJqNkzb6llmhN+svxtyGofpa7aAnesQTB7bYNfCNpBgjARx2SW0cbrHfAq8Fj7S
0W6Vk6Scov97yYcSdND9JHMWGG/O36PFQCTFVJD2sB60mV+Emu1rW8IVFyBwGQ65
hF7lqgtuezuwAKGqMTEhz5N/bWtEQfS1zORTgEJaSaWFLx5PUjjthCTaYVBCBZhD
/bSoph1GhHpP3Po2/tIyAQPRCgsadSgw7zkbgA78jfmzyT1P9OOWlXx1L/uo2K+D
VH9O5rda4PrIYoo4CbxncbI6lwccaa9ZuGeNbz6hPD4caVShkekcChi5PvngAHV6
TuWnjgpuT1tE1FbSVS0fcAaYiHhmifMyAP7pmpbUHpgd47DVtrzNTXG0/sI/h1oN
GwKGUFzQ7oqYgHUt+PcJ/0hutPbFxJP7D3TMB9+SnIzkWPyrn/y7HqBhXe+cmZxF
zmG97ABvbteCNmyedBSH90PkWg3Br+x2R/naMO2HdqwQRw/l4tLEOSQNPoJbJIyK
EjcD1vKYlqTjV8cQnYdPCdVXiZQwOqjQABFSDYlbLOY/6J9fYkp+gctCNTglNhkE
jOTvXdrik+S3dOazd8r2hJO2XLMBJ07pp20J+fupskch5b0L/DFMurVwaGd5XmY5
9hz6M/rC85GY7qJLdsDA/gSZV5dXxwMzWYw1EygMVis3UmyGyiJybOsvwKrlkF/1
5XtK1IAndKyfzkSpMA8lYjpTjk2Sy0EebOC7lolUBvWRH5aKGuj33SKrAAWtLIyt
gNRAMfbybcnJe6rYbRwVrCJgZ42zPyfb62E7VTkdctiby/zblOjUeYoe/N2gEgrA
jgPVJM/qrEjbcqVOhhlr0xOErFd9IYbbl0GpAXYT8x8ixAdxA8NSkjj34qSilmUm
f39a9P6vVvN0qCMS+R0Npz7nY0x6Ct3quYHk3Q/lcPThfrw4uG6P+jxB/w4U1jxL
MEjjvHayLisTp+6+9cT6y/F8t7z4iTBclZyQoIPyZ4fBrnaOJ9MrXou0riAs1rHD
oKL7uMkfDIMURQr3OF7gmQ/XZ5iT3AnJqlD5zShr/hRrqYY6xKsQ0m5h+t4Fd0Bl
SphxzJ5wwzDtXWaCqBPpBfwwRI0sZBKR+8LpdmTYwBrAc3nazFDsICyLqGXpW0+j
SW8vokSRC3WpkKVSNz6eLyz0bkwq+iPmHenBSKUimg+qVKyDpXSvc7pbV1EjfA6b
czFwIV21jEHrMuh+vrMs4zhFAvJL9T8ICXKASGyldGxYbZUEtqm400XV+4fLwHzV
0dLDL8cO/fgXpC6d+pLyt46zF6QMJ0JFMq9J4gSEkRISmkxM6rtJ67Zj2HIKq3y8
ofWN/5ve5ONpayls9FhrpblfW0/71HZwTatr/xNvlNkNYcEFguRPFwi65wTo3Ak4
U2GrE6ARONucMwwUSSuHDJGJIkxdtpvJQSPEltLtV96/xYVCZYwdxblVLpS2K6Ns
vxpRPxitpPZga+gWcHKELde2BMmRhC0cwEW4yEoeMpOdWNAdbPyfY5ZYOJTvx1uO
lYoibaKFMpAToktUTVXbmk18E/TcaDS1BAAMEe9BpsBHCGQ2+jXtevkLRv/pjQ3Y
vunn2o4aQtb85pt2pbiYOA9X3s8cSXMbSkeHl3bvmN04tyZ3ImzlB7zKC+vTujEU
Vw9AUyce7CKXy7357KOIHpnXttSI/VP+oAJnGzHWizAbLv/T5pz2CX7wrUB1djSt
Q4HW3k1LTLvWZdr2l7Tq8sOEsmneBh7HfiG6knYfCdqQZDpszvxKTufCEXaSiSFY
1RSJPbQaabBSXMkdRNNfHUNpWDexB7MGR8XlDvp7REPJ3FmRvm4lPvV/lFXvtkBC
W7nZhGzcK8tduvJQwgvlIqfOgRm04M1s9VLu8YolcMwjEcoYYPosgKtb1rHb9Hx5
5iOy3Mp9HVbUOgQfOZbqKTq6oLVirY1GweerF+r3Ls6NQQkLS9ZNkuADRZVMVr/f
2Vhk90hkuHkANeAjzW1UYBmPoJpBXxuf+XY8GXYPkC/ANthrH2Sp+i/cmAwTIdKX
7glMdpjzzOWmwcRPcPzQOfMdCqvHHS4t/++z1alazJdK2mSubdUs6ulxnHN95qZi
o2hy0ZWhQM/sOpQH2riN8PFEcFBDEvyPNWikXAH+vSmg1hjF1R4sRyJVid574h8x
jm4QhTHHtyZLzae0S8jauaREA1S6dkbbnZYZSa3nZj+tJUXRYUZTpBRSfJpogKoe
EdZ0JnRCRnawrLr3iNoUINlF4F29iJnnPRXHVFa/2wUW+sDfWvr+zEO04v6soeC6
cQo84vUnKk9drUEZ0mPpnr+4WKpySRnOhV/M4590sJ+7nkA+meWjNj5mbS3Yc3KZ
oYqfnbqJO6D/ZjZHeX96RMjI7u8jqOdnRUH/9mWv0MEvVL+gNbztpQ4TDy1V1T55
7snW7WUS98/DtQ18OCsC6REQoqQPt5QYU6e/WUYGt4VMCQdRWimFuYfQgo8bi54b
2hbcNnYJxxPxXZGHsmRLAYOoAuZ0u2/aM+cD5q8qcKWnMj4eTfIP6bSJZjwfASA/
dL9B2GJclyMu6Z0xSWbgok5ieR/dU6AdZVR7iN1LGvf7NmZyQ2D5aBiYWJtcZeZ6
4cjHeY1jIyqySIeaLpTiDSqjMu1+SoKTidpm+R+pP1Vm7pKqnvzvigCUoQPilUtp
nKAhJE+J9y51FdiowhgGQExM9oiU/+CI4iQCSL3ZMPBko39y+SdYhN/PfcZkkzm4
AQKSlCFK0EqSQqX3bwaIr0YyVCeqIWWJeruaaaeGABkzn24GBkJB2TWuxcpWb+V8
KXsBh32ZLvwvKsPwriJ904+7RQwU+pVsxu97AKKQlZmM0gLaR0VYnaN+0xd57ORb
Ou9gy40K2cQPit3dpgBATPuoBoODLjElvPOlpMiOa0OiphFDoIrqAxYv1lq+Apu6
sSxw68BDB0cGIY+DF/b1Zzxtm6fDm+t2yh6tg1W2bdo9bL0SboYPbrx8r5JxWMq9
R3IzRmhis18Crkrwy9pYbKlbF/MxgHbJUEpXNfq1BcSDkhN3QiIUQgX1qn482E4b
la50sh5ULGLhLULYXujoxpTgr6HjEBEr//uD+YrqDyA+wsiGm+Mml+6oAA8k1v5l
6Z7eUOBOEIBVfEe2PUPT2J8X9bkytsTa8hvZfqNYxWTEwXbIb9bqzl2fWKnQkoBQ
+kgFcc2hdb/YO5SBNFUjmM/jdqCBdXiZcCpn+BJ9Viw1zgYROXbIKco04ozKyUrV
+pr9llobIQ0Se15ewvK80wSm7LwlnJXB+rWA1aCXpv4OtI2dJiHvSsGi7W3IKAX6
ZEJ3lU1c2fHQCwcctbX+z3xpfeRnphxPVx6YZZxX5TUlYPXsDXpFfXVOQoT7Gp34
Q5FtAdF7OOoLVsx3Nr7epXFLUPaxdklvE5ba3p5oA6jA/evhvfQcsBI3YpY3kRRG
7NkUm7ff41XjSvjgEwaVLtJB7JxMv0uVu8OaXdxxJK7MaIIsbQ++CT95hokGraUp
ky6nJEoLDzT7szyun6FwNaRwyms67Dcx6hobBcKNBWpOvG3ttg7YzL+eDy/NrWAf
L3X2MsHZiObndQ6GLj3jlugFDfFdl9L/BuAcqA6g1UIWjfoFVW9+gwLRDxZ/AFO6
iuOdo4ZKxP6wN+q+3LU3b80znX7y6tSF7nqT1kmgW7jX0PYPmKCktebY3iRtRFyr
t4JZPiPEg3JXr8nMUhNPw1I8cHbtfGNnjsnE43Ib91GmsXINrl2hUCaebbb1XNLy
w6ugB2fSri3Ln7IOdwsN7WZOzJrItgHtQFibNrAq7JCQ/458uEJYPPDI9KG896VD
gapvPpg3R7eK2+oagnKglpbjQLGkZBv9DPDHABo5XRIW8BFNs4dZx7c44vOI923A
XNlNXUj2+C3+ZA71HGn+TuyjMe4eO5Xm4wnVIU/vZ8jXpD/IIKpkIFj5Smv/KHO/
PRv00/2H5wQyB7bl3g7ZSvCGI48LWgN1N5BBunie2zjevylxUz1al0Ji533Svtb/
9cNV8DWwcBlTTMokH66tzMTgQNPtY9rO9nDi7IQHUNPtMX+cK5MaglpcMHmy7Ctd
RpEEc2XnFmpWLCU2RmGguCuSH2jwV5SI+T1LajJB+1q6dGLPTPLMr4d6hSyI4xZw
2VprUQWemijniTYCm0jw/TKMji2S4VO+m3TPFceShnVokdI1yXwjXGjnZ426JS/t
CQpC/4R3L1DlpDtv4GZKwMvz8QVzg//foGygIC+5R8cCebXxrj8vqB/vZNPvnefU
H4kE6c7Qg5Znw8lbXvRlHsoxI4DOD6Qv5dWsaju1So58u8i4lY+bzH0ENDKa1zIH
QaRcPrJEYk1YVBxeMrKXwVY911GhsVwc9rCfdkeeMHZkZa3NnKmw7ZXalU4tar9V
82d8SixzB0IgM2/Lvikc+MGhshvKp2bh/lL1TjhbtmIHI8/h0XkqQJoRLyoRcI9F
cxak6eXrMtSGz26KzAgpobrSYMlNcEGXnHDjQ2gEflcFeDuSEka/f+vuyNyzlxkJ
QdHcDN7dhyy2zzj7y/o7u2X8Oos4tMq1uAsvBg/Jm6qF6FsftOZx13S9gXClc4er
zTnhLJB4YBQ9dqxc5pkpr0zOpVR/sRBUykpURLEAxco2pqjuBueDGABPATrXvygw
XPtvFSSPA9CUcR0Vf6IHcf4QxarOZKyWHNPOpwrzzdy0MynDtvFR9V695SLrrwCj
Bdm19WV6k4uGRnTWpGQ0EyJ4I4ODvx+FM5qE7eyMb9Ob8peNb6P9969qgH/6xs4T
kunjqPNBTtrzoVQyBOuoIRWm1/xJHtL0ZMKKF4C+/27Xlotq1Y/vZTwQ4fi4gHOz
UE348RFjlei9MzgR9IQKo1F5jU2016rlNOF+yOt+kIkuqDsDih6XgcDsczVMcJpy
i95XRPAWWK0CzqCsuFAW+1N+m/2B9nss644nbHXLH7ZAOyztvl1jaTKbT22fJdOY
UUxrm8LikwBOlMZgjj3R5kiykjSIIZDeNG2ckacQIVjg8hfJQzdyJdk4tcyUFngh
hUjx/MVWBT10JsyE5iYbc4CLrI1LS+gei+1C4KY3Xaeqz5gnp6VLI2JHgBOmqkBa
tiBqPdD4DT36C3STwZYL91H2yI9XJo6lVSOGq9aLaLH+xpX7rXQvqokp9RznlorP
+RO07taCxKMs9VZ+aGYbY0EG8+toumRjyLPmFX+kixhmypHOslI66CjFekkhRtM3
65GwPz1U4N/79SQhwSCIXhVtox4E4NxJbPSkCD/uxoGKeDvEb6G5ey8AbqmJO7Oq
xvTImoLldu6xjSZofpdDSh4F8P6IbdHdG5H2wJEFrpour53OQo1kqvVa3WAPa/HL
i+Ht5IPAedpqhV9THK9fTBATxKSGy0M8o15OUBAXXseaffy7QtZoBG/KVaY/K4uP
SHXxCF4nLjVCn0WFMrIBp07ZFtnLF/PCLBgbzBSsKNjEPItA5DuMHeQIihBcTVss
7sqBEQ1z9qdjEFONESyyEl7YkNQC3GeYupwgkzUt26lPmjN7w+0dIck/ZSuVXFD3
POK2Sv6SLrx1LcqQVyScTR9QW3n24AH9s5LR0kKf2KgcB6RBwq0qYZa8LNtO6S07
PcOcSXXIJiwhYjYXrfhX5DV6uqPutGXKQf0qNtrEf0e5aodn092SYtjA2CmZgxb2
8F1ByMDvF4Ue0ADySxn2WWfdcmmJosvT1+JirBDYc3el9IWX1UcpyaeMYhTSzhIt
xONuFaQfl2eQL0q1M3DNQW9NDhV3KxpIN0f14BCj+X/EsmyrwIaSVaQgCMWNFncK
QqsxHMJLTHH4hSgRGBufiDsqtdpG5c6wEDmkK/H4PSDfZcKrj1osTCS12lUFm/au
DQIYR7JELrHlUybRiwR0nrr/HbU9/wl4hx78eSo48rODY0EmSXwwJw4f6brRMEaL
K0cDWCxYum3bzNGfX8onypcq5ddSAiU0nSAJCHCsE7Eu/BNHo/ByIjJH7okOB5EV
Fy1PqGZZEjvTMcr9oETDCGJzKdoVzlqdeEo0Vnd8zx8FDkN+5XMtT+yZR34pKGX7
4v3h843nvxcGHjfaJl9L4ea+VTAf4hMHnJCqvgD50T5jz+95a8Iiyb/lGf4ptMO2
uYFe69SinY33Q5wEwNiXVZSMA6QlJT4RJFe+/4d5m/Wj8KKaMYdC8zCtO50BYnqR
TrVLzaezEl5HnhWb4lPl84LHBFKrYVI9Mr4YI9FwC/IlwE1rGEhc9/s1/+gz7/nm
5WdytUnY+LDoforVH2xQE47W58iY+cyEEc5xbRxaKzRQPpT753aNlXac2xC+19n/
6+8Pmb93E8NxbC//ycKzO+UZ5Wxx/B02Xyp6bueTZkbca8XgYJqf2rluYBisz9oZ
VdtXbZgTZtgNB01jGiunCNHoQcnF6EKOAnvwbo/gibI7TSFQNL1urfkFPo1XZNkt
O6FAj8R4bpAFHpLQrNS2uGGebZQkEbyLVZSuxFDvPh5YWxxXIPJeMspzwYrAK+eg
9wFHr8aHEoI+jtAwbv7E21wimzDMINKHi9WSi3ZU9LklJrW5dvhOyGHB7rfgwKvk
g22S7JqaIMfAcbsfwktK5ZCs778/ZnfryFTSNNw9jvkGEoOFDcSMANWGpTNduWJV
hYzLQL+E1TTKmqf9fcNGViCwl1lj8pj15gVA6f7SR5lzqfiJUh85DXMsgoHpstuv
EX6UwIxpB2tC+Lb39JA3qfWWsjk11jso5uaq1d+8mJXm4hjM+2UVZvamzpAF/TCg
IRKZQzEBux1aA5Sp8gdsvQi11kCdtBX/ype5+j1V6JVfAHzyeF75YiHcwoQtvXeB
g6Fp8bysBN8kitMi2To7yDEDXrGpV287+nNv2Rq+mQOJH8Ja3D+Z3XfBQFVanj57
8xcuYsJ7wj0QvLg9lP3bhw1xLdYagmo8mS9VnBYiEJFSYXoaUzr0ErKvvzo1wnC+
0gPVkDwreF2cv4m20tfA6Y2lZGzS7tzOExx5CIrydSdkuD5L5cO6SbbIm5+2Ub6S
CO7LPiOmRMbAZunTvB0o6vFfDLCbQzqxDNCXNGjwWjwIe8E8yLOPTds1CWRv1Ave
HmFI6FdtBHEBCky/Y1/vx4Bo9rmXxlF2+lH7xlb5yRzc05ZwonhJ33ggMnJIEVDL
LgxwUuU+F4sGFfNQTypI6xm6ojy7tjAdqmGP1AkmL7JxSuDrHmMGf0uX4k1tAE34
zWb1MK5aRvglM8H5nL7JPQL+2LgaYUk/BJMFcwpFJ92BWzYHQlnJ3IJAyVDaPRS+
u0sHr+IRW0qXtNNG6hU7oM0tlOpdgCPDNo7YlmLKRS1knzoTfLY9xPuTW3Ts6BGx
JR1XnfPgHyrMxyZC4jyGQQV6FwEGaQula+KcunZUgH6zQaiF9zufb7YTnOI9MqiQ
VBiUVpSDdfViw0RXcy7AbOI1CH8ijmMEpIcr88QFXcUl+fKgTmpz/C/fpYd4XUW1
V7qeJOIA5cSkWrYmbQwezPDKMk6tp5hv/b3j90gqx8BTSX7DnJ6lJ6TcIHronhwV
WIYgOjVlDQFeVkAs9CA9nOHcHD0ClYabY1zebbSGmb1WLNYdNm6WmN8jxN5YMPBJ
6JvNPkeq2ZjBF5Fnfg2dkbCO9aleLnoB4ZKt4JAT8lTnJtwrXO9w0h6eMJHk+kgj
AL0xGIBOmLji+UoS5ep7VTwyCZv8ccJk0pIf4vnLJ8/156I8doxjRUgvX3IL5GXj
JKW81Q3lgOalegv5AN0HfI39+fu4sV5WodLmSYIVoggEpxXcv7XEP3oNHQ3SV7JJ
Z44tMZTDRXLbUD0Jq4MiRU8nPgah3HniUrGNigQZahWLl6Co+I+hWhDdGr+zUi8b
tznbZ9fBOrGoEVTo0cx6ISVulIDq+duDjhUwHQfybj/A/OuTiOq5s9Y+2jdpSa2I
lRqxc40z0uJ/BleAA838smfD+QcDPm2uYEDuBTVImawJmO59ygt74E1vQvZcQmKs
DyzfIorUJ/MaDT6uNPvpoeix2R2/eYRdQhltrMeSTCoQ3m5X+uMn5+j9MStogMiX
sbWL5nKLBW3xCFRzQqcI53YvIOBw6FNQCT97db9/d4eJlwMJCz+7DUM17dY8lsb8
UarrEAmyn7wWRosCiHAzvi9EiedW6MrFgfJiMXcD5pj5Dj6EeJu9SkeW1+wV4YB9
dsPpIUcpiA75SKtacKMXEmbxCU8jw/FJiOPmw6ErkkRS+VJeZ7eJHCIXaeIv7DYm
Ak7xsrr/TJOUMkWJV8i33xrxEW30xg4HDYKOTiIJnp3IZ5p0Cr3x9RNB4lx308Pa
A+HBhAxvVwLLkVAs/FJ/hIzO9dfe/hrK8s72gxHThqADYDXDWKErhQaftyda6opv
OcH4juMa3gSS//+sAr3ZV3GtRHY3bnov95xbluPvFyuntNA04kqmXPqqMRIRRuvv
cnxANWKlWs5oaa425CezJ6G13Y20DallJ/Hkqmo21Si+PqwE/63sWx6Hm6UVdmp8
C/RdJBH0KZQVDp1bEVfuVzCXWN21m0ZbTqgOhdjO3dmtUGM4CHadh3K9AbqgmP29
yzhHFe2hn/Sjc46SKnD7T7yU2rs6fdT30zXvKqDWBu2HihB0gv+hzOh5ZGHcXAlp
/P8UnDsG/+Nuf+esOvIHaWQQ8Cvz481FE53lIzQzaJLLpiFoBxtibPNuqi+kRRac
OD33pBFDxbNUMNUUXzb0myg+LL9JoeajQxj+v+6kXUvJza7VYshJ5kYviCXKqS8q
L6VKgcGI3yHP+w93UzK5449/KavpCfsqgNeRyB67RixB6BIjkng0Y9n7SOb70j6W
KPciQQfh+CAOXb/orL6IPFkSzusFK5tW8n2Zb4mbmiQ/Vmuu2QmhFF5rBZi3SWJK
lK+mXoWdDDMbJ1F8efrrJVx8EwP3YI0LI7y5nZKILp2iAxZWOR4UcJO+yYB+idpK
9A8dj8lRDA0kQovBbqa7e1aRsYAVESJiPGIOpetnp/9V0uZzJl4hYtQCOf06GgOz
eEllkXYCSujPJ54PJqiITdbLKGoQL9Z+8v+zSHt2NhmvcmzQe7WQQQyF/bLpCho/
DKJnTrKVHOqT0zPP3WnPpqxfaFNTtXu0t4YhXOFa8VdBnX2ZTYEgIuir8AIEMtxZ
WVNwVtdwmm3bs/oaR6pjNGT1j/hR/CJWo7WX55LqdGyS+yzy38Y6iZeQkrio+qq/
iarmdq8fUlW96FgZAcvG3savwgi2feNS1GlG6adUpzYU2Nwwp4Se/5RBah2vDA6b
OdbxGynMduo5I9ZUYZ3Akpxq7Rzh7m2FT/699raXrX2OlMTWM5vLQtQZWwPfbbVY
Glb3W89VMREIbzEl4DEaqRTf6QCJsNfhtmHUhUn9OKd0e2Khqgj5EgIpWrLWlJzm
8mqMynihREyhJWHPWTWVcHrORwGloJc4Qv5JXmWp6Mg9QUCm0Osa9NUHFchWs0l1
+P7EknbzMM1G2W3pe7Kv5+XIZwMo+u6AAMtavPb3m3I2LiAEI+nUGHxa+NqVeFho
g8BJcZb7WuoDEYcRk66Acs5vfZDyc6/sITExxIHOVI9diso+4Il/obzN60o/vaW8
zflNofNUBgg4S3isAbVXGXH8Zap3RX3B4i/SxvISvx/Rw3YQAmbhLOTavMJKMayF
Xqg8S6N6sihKp5SC0WnaT1MbTWw2M86OaoPV12LyPi8bb5eGkH6iFrhwQ2i9cbIc
3NgXPm4Zmfmmja42h4VY0vjXYe/Cql2uA1SC8Fq+DqS9QwAUOVDgoAmCY3MqOQKw
9UpqCcZf3uTY1WXaWhgum3ZLxbbBJuLoWVhqv9dUbM0X81qBkpM6D6RKMyBwyD/n
F6vWxPZXqfvMJR3ehrCiAgMNrTHMr6hmF/F8IPnwz0w0+u6AxpBNCzJZbc9ODcFg
pytwlhTl0/kGkbOfVA+pXf+DjI+XtLEdwKNgD+m/ZMV/aBAejbKjvDHNrDyrfmaz
0fJLj1Q7UCZ1UbdWn1FadlOoCQlxnXLwXAKSZdLwRHAxurFxd27wiYgu/3e+jMFR
NMmUJuZ1I2oT4D9TZlnvvwPrCW+WWrFVb6FZUzwJ0qgWu1xkpr3fju/BEDrX9Lpl
mk0rpeunemDwEixMq4ZZyxlKpJtQWuyBwilfoPqMC8sJles0MHN8jHIztAOb72Th
YXkP5bGJw2+eHtaCPXZxtDNX6Im+yIW0rvyacUMigSfE1miSxxnH12n/HTt/X3LS
20UHqPwfiweBNSHOx3Nn0WPxVUHDbHuC6A7AlBORPl0C7nOitgWajPQrgA43wonw
HyBQKtixq1a/Fu8pY3JJZIcsCDVUAU8TmCGZ/ML2L//zi4ZlDlK8bcFgZ5K/3UJH
qEtAed8kw+rEDv9T6OI4VlLjV9gd3PkT5ova8R+DSps+yBAKtD6rfqOrHyJT1weG
cdOqUXHwCav5T172E8+31G0Ne46IlmtxBJ9YF5vAnWhGz5bS20p1m+DfOhqNMIM/
mv83kEt4+LUE7n2M4Mbx89rQstN5FrK20ZrQZIFunQrY6741TNOIPEbz+nH2zPxS
0mWe/u08cOQelVphQepC5baTD3p+ADUKTmY9XosUU3PbDjZdz2X32ck+pdxC+lvK
okokycyE+48ChtaJxa5S2x4/nRs0jCIjyBycG0sS/tjd5IRO3xsZIllRCOKiOPP3
rD7W1zoa51KxTo0VmSFZ/RSy/n1lmkHinuEjSWgbG5PeGixaRqOhQBkpJC2f0iY2
cGJ5DdyMROq9KNBJGmamXmy8F93B1WEmjsuAmCympk7o32lAdRyZqnn6xLgocssW
65rSIQTCGuqK1EMUOvrMmyoIbwDRwGWI3/d/mEfTkVDftrVKUEZmHkol9Xx1K1S+
tnd980iFQiKpV4l2km3HEuWARQSZCUigGtmp/qGPfbeeez6cInIulH9eJJ1hy8vo
OCjicJ0GQVkaclqc+umPKQbQ0mSu9qQ0P8rlCjGQnzeQRe9mL1rJY8+MhLLZcqzv
yjGCFDM933Vk+8HZwZqjnHH7qioBtpSyDUxEjt/6VR0KxkAtcueaIvzcBqJgdx9k
HQrQ98FOvJM9cxRyM1mO3eYcI27v7n4B3YRTPJhN0ZaTJSGdWkZ4z+qo1TX1ywUf
gzKVzgOdxt0cxba1hkPST8JbfVpLfMd05sb8BHyNkYNSz/Lmktrq5THipoWLI+aL
+egMzMmJ5q7KdfRYoD1H0CFEw2rcbodwf2R4/q4VfYKd/Q//lZfe80h0gTgKVSQs
4kXWFP6XTZQn8gfNjdV3ZVOWbe29RyIUTsT+txkWZTyemFOhc1tCyqFgufo9YnLq
FAjSpAM337F61rBSB+hFojc+eWt3J6sUIEqThZALM495PXV0HDy/rqiuizVgHsNy
G8mw1NOJ7prhEc20sqyLQ3ySvK+XqcR2qu1Qd4FPZZSVK9lzkMrbX5AX56BhQxBL
/ypAh9chnaUyCa0HFwOUrHZfIwDImwIl6tPNKNjnbad/0LUXS0heftRIzmPrTbpi
ABjkmQ71yEjZ3MG1t9QfVI5oOcdyFXoFOQ7DPeegwG4YORsZFT8SqrpfE4Fn/vBG
uPJ026YH0ocRAfGUesXZdOMmUukjIFxLYKzvyvRdV/eqr/+38AdCiyzJWX9dbWHd
1nupPROAQzi4HQ9mZratuAr+0kntfAeNG+XcmwC1xzvCI1Y3GHMQgPgxx0YJepfp
epgEsdbRhfYs7+aGR+o5Vzyu6QpRWE6CIF95yNSP2dHxoCZ89xM9aUWqWDYLdJZz
wNucM5NJJHuVVyrwcavOILNMXh2wZT+plE0SX96cq87pMM3hPcFInlEDWBqWLO56
nZ2MOoBx5eRCPXukpkAtm+Dgs3IhfDvMyzWKlXP/dd9kElx2nbF1/0xQCUtLl8fl
7uIA35DsjzAbfEvUB6FGx1bf0eWVDkZFCgHMoTj5J1+aSMAryNeLqB1q51afVt3T
d0NMAZZahClvtQMO42eWcJZBEZ1fzvBdy/z+iU40mtsf0wPX5Uh5MJj0lMswaxWr
0GqI0tfVdQpzE/Cuc4JAQhbCmJ8UrvmRtVvJrGNWVdFBWcMyfAb2677oRx0TzA1z
ScYfIZmDz+5bk1qeY2jDqIDognp8JCetE+vWaTwZ9ueXIRgNE7SrFtRrMzuVc/K2
SXkDVJvk0CrnIkay/q8dIHLe5bf8v5c3pMxX/INCjwfpKU/t3oypUXCrT3gEQgF6
0e5Td7mUc++SWrgOcOjrJWD/MVJz2CA6A1YOM3OM1mHbpj272p+/mGtkVCVxAdvA
s9wGKgbcolCZMxtJQA1qQezJcmFwKPq5voZF5Wij6NaaUw51fLk1kjSQu4b4atKN
in8dNt/qcKi2fMqmpb6jZ6S0tyIaaV/XHExU5Pvu/oAuW2Wa4iD7CqF01b7hxZ+f
T9Dd3VTXB0xKKYVAwS95sNtYhukBdTKwK+Q9s9ssuOZVF6oHTkgTitMMJCDNSaXT
kTU3+aqz+EzbZvI3ij4vcwQR+3V0uw0qLe1rEpXKVVhV7hDuVwooUC8bbOtfC34U
xMT/+Gs+UIqpLXVmr/mLxuKRSp78HkaKTYXEm6/Yc4jTTO8RRdzoeB2Y6AngH9pr
UyT/aFN+/4ee5BzY1qRsNV03OT2PYQ4VoTb8+kbxlHx1t7NX8d6Xa4+2NECDGnU1
oQ9GgKQwWcaoGYmcujQdaCdNjWKPAAARqOplQ55gMxracMHILsko+t/+eDoYH62k
IaDPJPUSN/4oqtL6RmcOS9DdhGAkaWkrp7+k/DTY2yWiehNWeOnVBti4Z0j7S/s7
f0rsbVqEk6FJEy8wPOuItYOjAXtQN63lI6P8SSsz7OAMy74+oDY1QFa/FzP5H2x7
ItyoFs6eFFpsjwWDadTXwUkVAunZGakwjuKoWtW+7TCjzobNn1/5SZuyV1kJvnZs
Jbeyi9HCs6uZ3l3InamHiQbN63BQDWgjcidQX7zocLJz5QX6BsrjuX7zxMWa9yDi
/BA1lxjR6uD9NID7uW1QSCSch7/gwn5mItvIqTR4besS816K8hu5EieT5NA52ch7
EkFJr+fYQBR7M9aGLFrRl75FocNmqOnX3wAz6B9/Oizkq9y4Xu6I2OXuhTuJqaK8
2i+p3mb2kEep/g/qXjvskE93F5ejVp5+xqrgTKD8vNCBMoF/M2VH8WWfzBi4QfPd
PnwF3i3Js+ghzfs1cmDrpe8CeksUSb2ukGZBBdWF1rpM1/FQqzAa7pTKDvqUb3/o
brX9VXhKgA8wfI99QBrbuqpHShYIY42oMj8UuMmbATBbczju6XLyzw9cElPxiWRN
4OUfBG+S5HcFQ2t8ean461fay/h9BcOHtb3eqAukOxgxi1bBbHtqdj0yBAtiMJDq
FJ866O0JyYsmFkCYRGlShGngfsE5FYVjF2DK533v796dTDfLxQFd1GwiagkDGTvf
PVpODjW7eoMwXYEG3sKY2qgaCRf5xn3FnJ4AwNy81E/3kPPIphuGwHKLbFz6ORUa
GJqMOFxDwJgonUuyRpWZV48L6cdZ4ohEwxUmEhhOnHdRkki14cw4iByUhDYTQh6D
NyuRkmLY6OIU/BCEX274NRBxL8iUDz5BDXdXFfnbkZ2Kc0LwSLxH5o16t2U8UGNz
WWBOEF7LhGQccmp6ZsyH96d97I/5/fISiAMAN9CFumStLF14mHymzXgkAzKtiCr9
nBc11977aK4BmLHFRLuFSHq0YvYZ6MFwV4m9keCHA05T+JfvuCHndSxKVYpjHQ38
IuXxx76QOnkFfb555/AahXa4fZN9ur/yuB/E2tcnyv8WKmmkZO4+zVkXvqjs8t+m
pRELJg+ALtZ7jhMDk2QDc9GwF25JIN65YTzpBfe/lQtYkKKvXuF4YvhhjIXYOf+g
qUTqV3PwQXdmmyLuYMWLt1KBCqjKhIvkddiYsw9zTqZJnof6WGOeqp+8A52ZHa0o
2rPufQ8Y7HcBiXudrRWWzhixmwlgWVbuSoPoyAuRSH7D1q9w1eTtWA8bYWg+4Mvt
6DTW2MnFB2HMExcEDbEKX6o0Xsj6btibKQUzwd23Vsmso6rJs+1i7sj7DqdMrmEa
EhfaPkzRU7hjfHVyPLzk45D5041URPRTwVNAktadezdWQTqXE6y8peO740sJOIQd
TJ/4zB7XPZM/hYpcD5ntOHJknjq3Ii/He5bn2M0X3HZNWKIv5U8u7XM4acbzFT5L
PLm+BG3anERqKHpD9pmWOJyRs36bo7565aqkSyPNRikFnQ3BGSttCal0krmiJtwd
PLbP+YVXeM0rmR/4h9YYXuP8kC7BjkIoqtT96KrXTjpZOE4xHF/cugpe5U33y6oJ
A1xWmgupepGL3OOcwJ8kqAcVQlbkT0qaSf/B4yIdbXy5wM+gZWnSZY53Bj/rLrOs
/6EfUhT+OFKdToyrM52qImw+Hlqxld0W4hDF2SoY0m+PgUrtnTVOSUfG4cGWuA1I
iGM+zjuM7RG9EpTTDS7m8z3SU4TVXpKcNeVOCs/y4uoGO8Qk02o7O1aL7eIGkbcE
+3qh3n1VDILsSdRY4DvgI0QHF7t+TnvnsMx6CL4I6M/vtzFrZrllVQOfK0HqWSHU
k+2flcdGjWksl68FbW71tJszrCHYH0h6k6g7zGjZvtSO/c9gYygnptDvxFlW/2si
RNXRZoQffPOHtLLmT0mG9XnwPBMSYkbJcT8BN9Zra3H5nRymkRZlCyXyZHCcaRBA
XrLvJlA8svPOkkK61T/GxCNDrkPSk2dbnMAsz0uqLXPUHU53d5GdYMZVjTJ2v4pI
/uX/I/108i3TLKkbQ33/W0h0kkJ76LSjcGeBGLjBiC0hUIGFNwR/8N26Q2Wjh1Xl
CNxmB2NxgTBSgFK27Hnyqy3B9r3xLAPbSSNdQhz1/o0bwsFqYzmiyt4z+Pi6ufUP
eABDmYk+yNWLW3+EI48dg4TYbUs4GzTS1eawPD0MP0lbX5uTO0yNCaQ04z7h9E9y
x6o1Hs0o0BsY+JKzTV7TtVOV6/6vpgNWgvuP/u1jjYybbOe3LF5Fd2Ly1U6ft83o
UXBXGw+1MlxrOZxfj50w8pRkilG43Gki0EyF4s8N8IGGwcgFiTuBe8+mzb2VBAL5
FvG5DBDK0sFYXBxeqZv+cAAvcwhdofj2byeEdBC9InBqt3FVMOXUEMEG8zSU5C4s
R2zzJi0ru89ZJPMqbyylaj9LQw0wJ+hXqgedfVDU7zpqdc7IkRBdoG5zMVXeB1Iv
P/IG80yEzsVtYLD/gSx0ojOjfEhDNt05vPwtBJmG1ah9GC2SuPmn6dpjZWTIfw8x
UpriWPPHEEFybzJD7J4fmtaqETMI6LeZeIgKBQgevc+wqai8j5iJf1QYOhuQdmWI
Iu5lue+/bqnYOOn0mYJgx42dxn2ZuCpQvwK5ltz5H4M289Zyo57gp5tfNw7TuNmu
XJAgMxV3yhhzzQHCFDqolspWGKxe4et6S1XLIS9RXlY4VCjtNy6SRopruNxL5HOI
fgn9FQEgNafiCqIbJel2dIuKRzzdmY6FIgboJesmsH9kPqLKf+nVvugxu57iHmu6
GL4WwKU91JjhV/+fPPl4WLQ53yC3DN0V+yobv1KsaI0fniJwQ0qqLX4FVgfatrw3
sQJ/z/E4uuXBuBLjT0vtC0iMKwv5lvf+b2gC/sMd7DDaxjsYH/Fbqb+Y6+PMSsWI
Toeut0bHQ00gF0HEa4ExzR0ptQ5Sg1uUycilsVQC6jT1FpNCkJthyyBlKIFqinae
IWlt/mlFKnsEwKrG7JdPS8DnKi1O+oyZawb/CGV4NYuvW2ObSCQ+HuPljUnUWXUm
pcE9ZtBJBlGbk3xkQiL9aJxREmTd9oLJLlSSaUz0wGJBAoUulCfv+RPc8WWjKT7V
O5yzfc75urHQvAlep84UiV9OVeMz+yOKS3jPZHw43bZl/p5yomovzwG2XTbXrPFk
i5Lh+N7s6SRcZA2YrFvdVHR07CiSs160oCCWZMl0TUVxCTFYf46WNdzW52OOXYym
DB0xhTu2X3lV3WW+PirsqnwRPsM6KKSV2On11T+vkud3qxYWAnBnFOA77Th2HdwK
jW45o8F3QFuVXgy8bGmbT3TkO3Z8+QOTYGPB2JLKLSEtV3JbjBrnQfeMaqQhlk6a
9dFYxr5Duuo2d1+h82QTYoyAv7klQEFc1uIiZS50ZF9gJwuulPJ1RrKxnqK3PDtk
ihISWf9Mpjr20I62XmOhKAv1ejlReGsPnqzh+YqUQhsBekjhJiWa6eaO1scjWClU
1fFA/z6Y9w9a0XlsDhZymmD5cOe70BlHiCFg2aNUzTXuTKfU4WQGHYic2I/dvIfm
SJRABVsiqPSzIUh37qqRL7uTkdCnMXp57c43Ec1PmtgAATHchSEjVBnAY1mJQLEd
diL6SmKfBEXArJTDWn8Ot0whHBkmtqWj50iG6bfHB70vPlTI1sl5caXYEJnJ8jLi
VZYPiHA2clk9dJkxIrQ+uGctsyAS62wudPNHyOlzBhRxs+NaxjwiHWjbyRt6sBSw
YPAJZ/7YVHpp+TFYlZuWgsro64l7J+hc6n0HIkF3VgCAAIwvK74jbxoVQiTbCuju
NPeVPf7YD8Cq6y47gWzdJ+dwmm6u/3wjqdH1n7VxNV4iVzUBDewHQJhDf1Jdf6iU
3XuuOJ3f1dzZmvNsZVLIsDkWzjt7Q0pV7a1+vXybTnwhZMbsakintpmIJJwUkU49
qfM8mWZKsLLMlbzZ8BHNbjPm9nOpmgW/kZHmYJ9PB/f9jkV74GwqAJOqnSqzgX2L
txvpg+NLR/3pCwAutDVscEkQyScGrz5Jn9YoIYwNtDyYaptUoslb11acbY9GEyFy
ZQ+pEOlEM0gTu4OH/2V5YtGPkHl8Qml11ivv8YhSoX1wcOu9kH6PunRfr3/s4DSu
zkoQ/RsdgxyJKEldVQSsJ7+pS6JvqHW0KFxaCPs0JcfdvrdXd8aUKgl90lpsGPKd
iBoVFmAF2SDaDboabF96syRiv0d93cTn7Z0uMFTyv2hN5c6iVF0pwfgeC5iHAdKP
B2MyhQ4O4ZDsh5XtLO23SOtettNglw7ffsamxiO0v5i4b9CA30/6hgOum+872Va5
ds0GXtEapLms+6icnJ30L6W4tKezLtvKS9DwyBcppJ9RKH9eHw0BMbl33kyPWBsy
DzIwpmhcGXlyPURE9Wzsl9Pr2xe8W1wQyUCEEDJ0MFJwlKA+bk8I3x2+66valYh/
pwa0HbKk+0v1DuVDAH6p9BnbhR5h+Nv43twkIV5HpbZzUtAkGlHymlt1FL1jmPoX
+pM+brZfzGkUgX6SwUgc5o2cgsy73j1NbrMG0tG5vDulqEo+oEiPZ5AboK0r3v3W
wb6b14h40TFITFseoBcb1ieacUuAmjSfYtoO8o2Qp+h8mIcPEaM4PAxK9ktFXm2c
JNeoasoLRwHOGrAnJg4AxeVweHUO4CNWTGHRVH55Dd/SVKyxPGnQl51Mt4GXyOFO
k2ZbC0A03recxH2cEBBYOdFSekd8Y6q+M5o5wu/TanuPbNrz+QBs8/UPR9Kh8vlY
6kaCZ8qrh+OPPD8wLQ8CtHiMl7mUip5fOJyxF4NR2ZiXWnBrCNCnEAZsx2dXrGtr
fjBmp+6FuIhj68zBrqsHHtKaGeuZC6kGgQcB+mba3wpTcoklpJm73AnIc8P6/IpB
R3ZgWI+WN93YjRtPemhf4u/7sOawcKApMUkXls59MuzvCsvkjUh+jMEDx1T5npxs
l4DJ8sWWpSOcXzybUSyKQ4SbWYQQndRP5lVd7c2bYl88H8P2P6EtK1/OLStd4dkr
hGGigmu6/LTtDzZLEU14tB4RpIl5mvnOaxjJ4G6FEHIVsrJyBqFOEnySsv27vxuh
GptxOvdqUzo2DF1NKdd7RLnmB9rxM15kccUwf+oYOG5rBsMAH0tQshd1aCPKEAZf
DLVtQqgDb7BqUjgZh1pHeM7Ru37omTqjJ6Wm/0shotyqNh4UuEOllULo6ki8O+gw
UR8Qrd2QZpI+7roJbk8Hw1YDQTwQ7fd5h7QwsTl4YeoieiIveOhEUokbzlGtv7H5
WpgZ+XyHiKjTLuLlZ6CW1m2gbpL0yjXx8xEnb0jQ/OqDmkjKaxb9uj+qBZNCHf9w
AlWlFeQHxzHBTVduFcV1jLZ6TLIXoQmCp1XdgesqjG7sor0SXRAQxXVo4sn6OUo3
j8Prv5Sq9TlPhfxy4aj1IMGrFvgHSbf9mi2Bp/C93EInkCb2LK8/VzRtcaCAS44Y
5D2sGXb9sOd4bKVgs1n5bTtTAV/Se/86BWSrG7i8iEcKXPgyvbKg012w8zAwE6Gp
0BDuZ69N9CH6bUNF/TsZAGjhpXUcwIG3BPbTGx3u7eMgD2SiuyH1F2IKWhu58gIW
MOYoRdijY4t6SGPengZsXTpTQCjfdlqFDsi1ZIeb2Yy3TDOa1Gc77YGhP4oz5bJ4
mU/brd0GXb8A/IJXgiE49k3/K3teAxkd+cY71N8lL0Fz1s5LeIQdy3vK5gpUTbkU
MvqIHGF2oFVf+OD2sO4tSpVfug677h0zsfUWTtd+GeANUIYa9upxVSpjxndKWi0p
UC7gK76iqVWjAjHKQuiytliZME+k7JVtrcsAc016dx0qKHs3YwuweJbRysCFAnr5
9fUmweIQ6X3N3vxJIelCIeEL4Trh1MFoG/tkz2dsONbaTvlOKCFhqQJvUtUo7T9l
0D2RcZNn/Zr7Syr2fQFY6dgJy5I+0ES6ZT+lp9pKAsHByfUoYOSTOhJOtCusjs/Q
ekcORe+mL3jaKrBQu95zFbE0yyJP8NTqH8FKrpBO6PI1pC8L1mbuFVMeW56TNSQU
g/Jy50UgqJQXnyslPkIoGF7quJVHFposEump8XLMS0JqmeNPNYJ26xtQ0LS5VQOY
qD+ssT9uk0FBXcgJDBZFgH20GS99MmT2JxWOb+nVu6dQvvfeFz/rr+3CkPUyKZN2
3y3YIb5wCOKHw88IG0fXOdclcIvZFaZ4XWEP83qqGSzzY9Nc99iS7zBakQKC+zXj
nsEELbn9Svodc+2DM4X1WXJf6SyoeFAVj8UqrGj2HtQNWoB7od+VCI5P+4Hmbcif
dXrB2dUQCTEk5bBGMTUNczQYFc3Ie6hpHdkHk4yUvDvn7MXIGiqvdLp/AiaG4/Ve
Hhaj81SHXIN+QIAQzWNwj6hPiv7+9l4B1FgVXaQ1HoKtFtCe9CCuqvLEjBge+KhL
eiyLDR0Lzy2cP1RVl+ahZu/Hw/mkbOT44/TNHTfuI3eMarZXwD6o++tDtT7tPG9n
0wPQSitjUPiTU9d3hBTCwZwvKjkCIoAtt84pyh/W5OdD2AxSvtOyuzGRvbU5cZi5
2x3n5BmPC9F2DkQ2HAtsh7Miw4A1qkM/Kv+uZJmq/RUu0E5GNME2WiGAgOs8Nh7V
72qssqqRjI57tREsiL9o3H0wJ6JoILR/+RIij7Nd2wU1KIy82W/SSGQ73NU1pcnQ
qzchulwfxiw//ASMwK2UbP4zqz8cULG64XN7vZyxBTRGfFQF/K71J2GOT12Q6Izw
mZ+ZqofPBTwWj/36vjXMbhqZQn27UFaZYCiJdi9Fx6oi0B1CgGvEZXwXogmZsd1P
Ncry4mfdDipNc2KTBMVCsGjUZm7u817a0bOt5EgxddJfeAMTnCXhlMwbKRBAv6KU
OCTOCxq7MbGKlth8l9Pc0I7ZLOMdadkcVBGMygAsEajO47nY6DwGZL203wrjo3gE
Q9vfW+vXUDWaRIWxHiIEZ9oaM84k2tilNiiieJoDhKPbbitxky/yGnrCQ7ZHFj5/
bCMJ7Nsi2/t6E0l10cl6BQclh5Sz3vfL9xk21OoXiEql0BUT1trAhJP/yhddQOzJ
jCZ2d1iAH0MRwK1MtopWMvPHr3LXtFZGrjAGG0rHk2ThDpVNqTzp/a/lQroLoIdM
uN+v54mz7njqW1pWjMrUK5QvJymy4VrRRyKgv8hsk4iYcLSBTIAXKuhh1Eh10ra3
mBKYYpWa6kV3vtFgIhB9B0pvujz87vh2MZGTD7Ct3oUGLes3Mf6GVzBfDsrmTmT/
dMndyFigahvXr2Eea9C5PCbto0wvzZpXqWet9yE/qNy2a1UNkgiwE348an2mpyLR
pGzZoYepQ07wzGTvKDi3yauV5SiM5q4p5Qs3sRffKI8PyWOTG8Rj+Nt1ohF9VciJ
hXcTbD5mh9wqA7JF960jT75s9N+oSIV3PLfXZWnO2Sth7n1uZ1kRjC08Lfu8GpNU
ucdQ33Zm5Y7lt8CiE5QgEaVDppUOcyBW6ewnoAIoSg3jJBfqMbB2xESaALmxHdoe
lkiRvji3UGevf1TYK3U/ZINdhPvteQV0l62LUYBs+C+bEhgnh7WZ4Mpl57JNoRgc
SRxZtn+l2CB4iUolj5lY4oAHxJvgopjSGDgzqNA/EQhO1Tfxeym5Ao1xauReQMAz
5+afRGz6uCsjJOmrqaA0ghNCLWkcqLoxqR7dvwDD6kjOW3IMRJPBjqeIopHT8B4M
lcnfXfPuvqaqAJGndCx8/BWDJrV+6nZ/4k19G6ZIl6tOw0U+Se2jDlRxkJbSrxyk
Rm8kHpylBZ4oxd5uZhnKFbUnhc3jHJxM/OtJQVdFctONeC+1aK+aCSGHAuVbXFnj
qybalqNrAfMRuWCXTgMyTZo1rm1yctQJI1NJXwM6UGaqNZPzJMkTKCBjYl1pQA1I
2EPapZ/u45vNidSMi7x87iTz9ZlywYAo/46nWop8LTqfXxzk9b9Y6UdE6xu1HQIW
OQsoKPzwow4NeeUJpD/tCDnWo+77ysSd+cWQ2B8eB0J0sKmv+N7UPLF/m98KR4uZ
+vNKocc0jHQ/Vmtd9gyinRW2GU+XhEXiZZyHJbBlNBjm7IS3AWjxDSR6xaN/ZCm5
ho8phn5sd/ck01snChGfY/KP3ZgqbUdpDdD3lpsRbGrxyGREnB60FuazTnPbGhp0
f/FRcRXA3ZHw19paJfMOMtBvUh6Hsd3OTXNjLhrvI53mtNIsPQyo9ZR6v18o/edT
4FX9uyzk7OVvKJXc9fX2AG9Iq8YieKgOLUX0nF1cxLRokVX5ZJ/5mITkNpHozper
tU5HJad7EjlDqCFPwMJPrymSpz0PbQqj/0l3afBvlFHTycTzfs6lp/bwISDFbhu1
C0sBeG20klRxYTnzU+EIiZkZfn37AXSV4uUIQw5Ne3gwBoClgrKSEXhtDXkJmXfs
399CVSkdAuGltzjuD3+ZOXAxCrsLqfdqlxkq3hoEL4s5dXKwpTUGGQef+lgo02yb
gPblB/wSS1SeT2+OS9yb3cNkw8b3QITYU+H1jnVRjZ91bhmrU/Qbv5W8Gab+mzSi
Ek7Dg8kKxz9awQu731WdHg7zHiSPNlJnkbVxAJl3o4T2mAAIoFiL9qPft7AYOnRz
CzhjlYMlCobuMpIRHe4cu5okHzZiYIThhgVpjiOYdwdJrjOLutPgajufvbOd7zMu
W2Wvyj7B4z1p5WjagOlbSpL4yc1O41+iUxVMdYUEPPFFIVOw8htV7gVei3CjM7IO
sSyCdPO1CF5bZTCoq18TwGgNgMBIUPSZaGVfYOLMS3Hr0AvU5nYg2zGo2tuQFqgZ
ocIKJWZzJ5l+OhBGs8c+rZkvmg5lGukktlG7Xh7lgOAHhuE6L8xpCLedihpXgPfj
R3saitsh8huajBlGZNXx7c8ekpOv+PRdG8IZRBoKDhoc8iDtrLPon4QDSYtD+VLF
ReH//U4+eCwLy7NvTkCPciaFR9QXXJSBbnKVb3cGFDLbRdld/diimSWo60Bdl3DL
KCPOSctTzcwmpt/A9BnMmScP+aGoUgRZLxPIosAIujYRp9un4nGkPPvszRE+I7Vo
DWf3p/0S2eQgOu/vrDZyJfJ5VFH+YOzDbbHhi36n9uTtYLI2/KCYkMw+3/DXAdqA
riC0JwrFRRQETLbmrW0besFtc5HJCr4GmoSi2q20DLzDqE0Uj44U06mYXQQ/v/0H
zDCS8UUCO5Vya8IuMoQXWgB5J55xXiWKkuSV798ciIKDgb/P6waLRL32aYEkxpGz
UrQr3MetoRpQGcidBCgQSRy+IjWCxuVtK9lTizrOB0Nx/K1jDXADS6v6wwrFABHU
qTwttTv4q7BGvFKZmZJ5HT9vr6ZCB/vuqcF2vUfkP3lZSq9epUrzxC0Qezb/xFyF
fRrZuJmc8gvivCKIOXGgg94mQuqZssj9ffJC8Ol1ZZP+Sim331IIgjBI6fKblRoX
Nk5IHIkyBfQ/LZ6jMJhJQAjqs+V1xdCHIJNNsIOXzBkZyxwxO0O1qBf/0jfAXX58
b/Ut7lxhDmGfjoadvx578Xrbe6a75QR76sIDWYquQbOI/6ddQNzPK5a6mD5hmJ9E
X7tjpPWb/chOULskWmn+zaD+ebbyCk0/pp1ZDSTJ0iJezH4/CsxQTW1FvAHoOKuS
4uQI7DKSfgFLEQS1HU1IiIFc9wEm+v352sD3uUQSJD75zEu73/x41dbYYoJnE+8x
sk7wSNFEEFo8AaCFQMUeYKy4ikntwPoxKj30wOzSOKCZfIcV9lZ2vmz6wRSAp3QE
4tUAyna/dny2jYt9X92YkBJqLF2+JtgyIEJf2FnsjqzktC9/t8EU0zAJLreMWcsl
G4hldljxzo9LuICCSF0Ky/blZNpqq9AGhstnhhIj3D/t2EqlRMvosyayXtzNQMGT
qyJvSbYwJyfpQzunkB7phEPLCc41WsTg+l3/8+sPf9Y1v77cKBJhE1j1ua3Rc2Au
7R+a/pmHRwDE+5URZD5S7PW3XrCnQPX0ZulPc9WRQcp5rDtBFv0xVnibzaldrUtt
REzBbZC12dZFJUbY7s9v7ABnENzyu7qs86XiX+t5NIOJqswsuuw2sUAwRJbWhCU4
wtzBNaioOO7mbQH/b2HnFZzKXlJNsljWJxl5oBHgPSswC0YXLDHIPR+L+7e70Ai4
gxg0w2D+MjTxyJBo5FG/8OKEqg2UIY3zRFBrtTmbtD55mHw0s1taCZhuMo0mPYnR
hV/Kv+sugUPCKzPCwnmi2xT4GHMVXU3QhtFKJ7nGgDjy7r4/zscu9ar83J4VFJqF
vWGRba1C5IJvp3LCgS4shgI3YOvroOOgnVuImdT8Cy/HhJbKoc38JMMa4s85fW4C
gVnUYfvHlvjJVwMlBIuMiwqMDOR60WM/LxFC9+VSUdcOkoyYZvos9Su4fTz+KNyj
8sitmE+VkLuFYTb0/iAkC0F3KD11pFSXpY8ir6JD6C3lgdCO7vAEbWZGsXhRij3Q
AmdTx419QkoRwUPMp3gm68ZNHnyRy95ZY45IRSwNkpf/psEbqYHruC9dS7/Sam3i
CSBrHh1c0WEgP5jtAv0bPi8SjhSz2D9qQXqwd0uSx9RdLVUVntuCoEiwF7Cny1FN
IrjI63ekqjrxZyHD0Bw+Jadah2/UVsmlrE36PxPjQFlgWmU7ahlXLcd7IR1oAuJ3
Rn5toqrTB78bK2Yi8Dzfz1OMmWoUxKw3bOQjnkXfwp89AY17zmcL5P9ELR/pb5js
vsOmxi7FAkKThdXNX1tIGoN6bSlgeZ22QZ7+1TGQM8hnjiiteQGQ5cxhxtwB2fq1
fywnmLFJQYSFPSs5INvtARAGfj6C3b6awp5c752aJ3Mla/5+9cUHfoRhW9KRSPis
CaYjRxPKUYNayWFZ0vlRRwAaOBTlIX08aDK0lNdK/OAoIbDfju4vxYDXugFPa030
R9z6NeNW8hkUZ8RLn+F929xGeOVtGm+Eun6jdfyaIwtJjpuIF28sg07KKGj35gjO
A7OFl2YxvdSiPJp2GcgAim2XN3Ms+QSiR2HyNgUKAOVXajbDgqn7bdzOlZTKVWeo
HFaAsx8V13sRuEuAoa1BqmS1CjpyA16YqglFQNodNL3XpegTl013zLvx9oo8PZXK
bDpHiIjiIFgTOvFrJdBsFFqGqaVPpSm9rop+tcl61jo+mPhoFIDlALfvFAEnK2CE
sCOyMb7IRl11haKI1fnlT4cPVzFdAUJx330oFYVz3RfRI8NBTs4fWltMwvcTBYoV
Ry53J+eaYpfe4BREZ8ZD54mWF4TAv+nB8ulGlQF1D9RFCz1hv78LxWEO3vQp0qn8
6B8+tluZWcBXj7nWtXwQGd2MlTsgR00qz489GiZEsZg=
`protect END_PROTECTED
