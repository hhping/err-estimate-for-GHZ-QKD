`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQIyg95w418slVp2q7+bn5IT/+hBXgpWjs2HKHc/E6H63lJCqOO2lTYs+PMMmbZY
niDwMmoOVKlGnzldX3c3Lyqp6ypTAvIzaJsIg8LwDH0WEsvMdJVaqZj7VL6UVkM6
QvsE7zQnDNskp/l4h0kxG5BM5Rw84JQbkwiJ7ldFe2PCBPrM6O1sf0txgWcyXMag
TpIujVta1ANtJuTK8PMJ5/IcIOFJXLhDQhXd5fw+vkIUlnqnmmtfOe9RF/ym0dV3
bvIo6E73h7NkGcMQIkxBFB79Pw3JQXQrCQ9MOaXlTjpJDXW3kTpIMaBq0sLWutnq
ST7xETIMBhKEXJCdCHVT7NZmfaqJO38G7OHAEEhfqyDPfIc/ONqVkJz+x2LGP2h7
4U02MFM+ugLE9eFqNNmx66RBIXUv8e5cYwl1M1AcD8NkxflckYeMqlbk77yop/hu
Ch+q9PH9gX36a9cJIrauyGLsXeytNQmVoQQSfANH2fRuph4wQNqr6FAxPrOOwDSL
gH8l5wqQLlX3hbY5V20sV1Ib/8yNNI+zs3BqV7Qz6gkZ4OQ1IqQWOa4HrjEWCWce
IrXsnEqd2KygsBGlJPIo+Bw63+F5wgW622FdWnaUdCLW4gVkaqu+OoFERPpQMLM8
CFBIJvR9zyNb17lPWXWB8pSEfPR+/mccARztzb+WA52L/UB1R6vNDt06eUQ3PREz
6AhIMIjPcqo5VudXvdKjxAr23ptkD1pKbFIyOUJ+idWHesV4R9UPRGfi6jn5fGqk
2LRPZvgeiyHNu11Z7kV4AN/j7j0j3yzhSvmzgGoQBYwyJNFTWVzKl47LtETuPUtk
+hyOXNiLtrIepRp3Z35TmKYquCg6DdCowqsVh1y9HXI1mvPIoLD+z70KjbA7zmDV
KsEZQRhY/oReZ6oJxeKIdVXqQjBhCqHJxZoA0MJNEy9HIMgF8bXgw6IAzxGukcH7
erQkbXxSr9SBWIebum9t8Kg/tE9D25RNtpBnWcR+t3xwUIj6h0+KikqLieAA/T4L
7KhIQzV2Sqn8JMD9sEWVe/amYhsFne8jaI4zK43zJt3J86Mb7ueTvkgiVwlT4T+8
BZKcY5p0uXsLMP70Mc/ADTfKJ9+Avs/tCi13+TXxMIlkfyhk8BKeBgMiZiVG9dSB
CfKzeuYH6v3kq5a1M7uAf+N7pA/pCmKIX3OoMJOuQX4vWE28O6iTw/3jfxTt1f56
O0fjRipnS1ukByTYhEACeriQiX9Oqg8OkKKtizv6+yW6IyH8gFl7jJplxIUmr83S
+EBbgAgvrMqe4ThChOuODpI5lmWKIGO2KwXlWzuTorzcKTmT1UZ1etz/vegcc206
NIZ6JrHkO4+uPOzsl8AtGNQwBY19Y8N2YhBBQLQimgiNqX5Fhg4MdzhgIYG1NweF
g2i/nyJ18vm3tF1A6mnSuxxotNOb6/SNadloDyAWGy216s356owzqOXxHzzjVL2B
qmWmabmLf55K+KPgd7U9HJvpromwUqr+CvLX1gIRB8xYitEuZSuR2wWXXmn/AED/
VvFJ6ebeldd/IHuNYllW8DUxBxkHx3E3fTNSGvs3/quFEF6X+ndHk93jEo1lCZ65
b+aU1W6jHp8mIQL03T0YaEfXaY0rOaxBaFO+HyB8THSSGsrcSAExCLiMiZR/mslN
a75v1bs8uyTeD5IrFGu7yR3Wd4RVX05zuVmG03lvVM2ZNPziK+4gxE5nVHizqzTW
yBBILJ2TSC8kDMral23nZ7wqSwft9LUO/dmpoLSHS4JxuJyo6OHof9bhGVATrbBY
/9SzII8rbCRKqeISJBk5P1nIBZevKQSLYJH+4YuL+WKxcNg5MUcposAZMZ9GvOsD
X8j3I4IVmXnAJIHU7lqSBgEtLQ4xinxy9ec2UxBTOtpgISRWwN5nJthDyZ86Oy2w
VHvEvxoS8wfa+YXZ+nbSbz9S9lLkcTURb9DSK7/oOnx8/xOKP/WW6ha+xSr1RB4J
Oif7TtMWdIs3iPkhxW/yQsZXkJcEF/v8Z5d+raGUdsM8GbBOrOnBk0wPNDv91jMA
LpwlxE2LlPqxYRmTQSJVhGvqv59qftDbiF6gfKiN058ycgJr+CcNRQPtHFpAxeGV
d7SClHl39kSrfn8wRmdVdg==
`protect END_PROTECTED
