`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2HVaU4n0Cxjk5dzS5NCvICH6mu1ACNbY6T/GoWf5wfqfI6np2FwOr2cVD1mL0u9t
WGrCZhH+bm048ebKF3c22ihrW9aBpZRGYhmFcDth2D8IC1UcwJp1A/+c4w5E0gdx
K6Ki2rWMlpZg9hQE46okirvpfcVb2g/r7I83RcA1nQ7q75M4pQLcm9G1vQNv4a45
RiSScPEx7Ar896C/ySdKBSCpMLb3e6HffeidP7MX3/nV9330+BMw8Gfhqpp/P9aH
F5Qz9Gy1gXwv2hMjmBVkigpcm2hh1ZlaceHT+AZ8gcW7kM0xg1CrHTy2WYDS3y5x
PiWLFfC4CTvSH4LjO8Mgegnmeos02AGTQB14adhiHaDY9SjONT+qeVjNpXQITUkY
kZaCDxxbrFPfTfxb/bwH+ouniS3uMWsW+tBVCGz1FgRsEdwUtTu61iY487Hvs7RL
xitSsNQPb7DhWpSgi6OSQzpp3bNlW8ZrUFDOepozHfo32ps4eo0xHfJ4xf2+LR4r
61YsAtgJgyRQ06GW+Y6fwTGxqxuKhtmQQSMAx2BC7vXnvgl3WvPgH0mhwwpPrzRc
FycFWuJracwo8ngMnPFtZ+AHIZmF3V0sD8U5w2yGSfHlKX1VUQzZid5P3byoJmt7
pum6ZSL/bq/iy8rkQMzDv9mdc2OFdpPLLp77Dn0uhFuN0I7Vgd4eYJ0x/qiIDVpE
b97/WPpWozRPZto90gUCtENIKrbDO56njoSWyqBBlDRB77T2l3QtSi/N6DKc1w75
rRItsbWkOSiarEvyYQz75NygGUABHUCF6UirM6K9xdjPu6o46oQpXHXE1s8dbpXA
RcjMXD+3ajKKg3E2mHXbTZflmbE4DacuRBF53fB8pKwpPiumj3ilu7BC8TqndpZ4
ck3Kvu1myxgwoCaKaBlLgOHcI0MKCXPaJehO80W9wzv6Yc/SpCONjOqdJt1F7Bkg
V8nEGTivoelJr+JvbVg/bwBre67EPwHy9qPIS8PPX6F2LhsUlHov44JuwSsNQYey
KSWOrrJrcHvr+uG+k5u+6UaIqzkzsRuA/EXW5DVdc8ZMrbdVUb1wuMkBEESdnxa5
IxohW5fuP6+8viCK94pg0Xbs5qreyKo0Waje4MXlZuTNeOLXGT/etC443nfx6fby
d7Eu1ELVfafUhGmFnmQCNuYQNdo4rSvGARi/8akPXIrY47+WVu8BbVElAqZ5oRg9
3LtURHUCHkb68KspqKu1NDveiKo9/RBRQJuH2YiP7pS6AIZaMm5pYZ3vZWUyp7OL
7dWhFAlEQ03rB1EYgKZZfTDE5WZMeeQbt6dbpUsTL1yAWwTJxMgaVdkKtw1aTrmH
BX//lJi9BPIE3LfZ0jLxEFadpeeIlJYJBsB09YsyRkVXKWh67i89lG0ueZkzTFbC
2fSTySj1fFoLuRQfL2S3GFuFJ6yQX3nefGBcoNtOVZbFPqZ4htnkFyQv7lFfoBK6
cGqV4ODk+GlzJwkn9XTNQ9u8dWv+vBEUdA44aMfuZs67QaNXMi56EQ/rhTO8RiOj
forOQMiB/fadSqWU7oY+GAFa8mZNSbOqde8B48ZdwJL+nQmlO+JJm8QPK1pq1M6Z
fUXY1ckNocfWBFHjbtE1Q3NHZGhyNKsjDBu1HDOwEH82ha31jrCfYdZ02R4QIe2l
RsbQs1jQ2uwqQbyQl5RdLpdzbAmVbu53pHmzrXywC9G5RjoM+EZgFQON3N4czXqW
RSIPBB3o2hALH5VX/qGRDImPv4iE6qiUQdNMpjx1MGw+EwFuO5BhFoZoLKl6WDJL
goF74qcCcpugMGarvZxbi4O5AUhNEYapCHtkUcioLlbeIlD3I4XtAmNCG78wk96k
+117VThl99015/Ar37IOpELS44WxxwnhW4A4xGahhBHx0EUEhLgAFMAwqZqoZIw9
iM+gvNRd+edpwytsZ60sNLrPLq1FvNcRqGi6cEaEf8ca0EzEwv/tm949XBJxCYAQ
tWbxKufC7H2tmZbPBhSTohdk3N75M45LtIlGsP+zJEUiWIJ8rQ9kF+Wh+xfr+TBK
HxpbTKb1+6ASNs472zjGOaLUtzb0T5iNtD3tERa9aiL+aoukDBdGZVXHk0dS8dTQ
CXtg1d+pLKUa+0xpQGVAUfW67F3Bcp1zP8EyZPUNWdBi0/nb4wXepyjE0E8gx7LP
HQp3lI1yOBIis448hguTNpFvIJTYlgvJnP5YusGabPRBMpRAzdPbKJPgX07ykf3r
nQ9svnzatrSyTS5CLTEVwCv+F3xsow7qfsT19GFdeoqhxvkCNEWCFWrWWgFHy3mP
ENOGX8oJk2kuCiBrHgb+qPWgQ0NUz3umT/fLXIorU6pFwCL2eqZXcSM1TZKpwhC0
x5iLS8xwOTykNtMO5jJtxb+hVk6I+vYcZ1i7M+ex06tTYNMzal3rAbZbUlotcgYK
pvuIyojy/fjdBUGpJ9g+cPy2vHTw0CExtVb6LIxoYLOGtY47pHibml/m/NiCUfWZ
DFfIceIY29cVwC4Iq12TTb6VbW7OmeswzqZoMweWNOeRlIprSJwscGn2anF8ukIa
U/RpffaUfgH/5nI5/r7lok3VzAZIxQvkr/5C+4wfZLXsw3Z2nYAKkKAag7/Fq4HS
BKBUy19YpVX+n0Ut9cWd43DY+4ohDeeS5b+P9HKrlO7ly8p48AmgwpiZz5getziR
nuBL9gmI7EMmzCfPpLpc27GVJE9Nlwe95fC9l4qQF6oUFClnrjuqxmujPu5tz4bH
YMQ7Zy3t0UNc8GFezryOhMA3N2KsMSIESF292F5lqcskWhYGXE+gE7UWgU7/hOAA
bztIYwzthSgYvm72Tq1E/284sXWPPYd/HiPansyVPK7cRYxb6k1Ii5qogqpV4KPv
/U7meiI39k/k4MsBWlr16fYAZZTMosU2HE0R3AdHhUqvUgiKv+voyfDlq7cdhI3Z
Mpgk5zw4BsILq3k/XEITmomI8Sbru360Zaem/7A8psw9Fn+n6MEWGVsZyhn1qZDd
zKcMVTnInHEZ2S4kJo7+wltMShdE/g7oggBZRxddoESdD4FVnTbbHv1uxOxhoKEV
PgTUVcx5uB4YcUwnjwrS8H2yGLio3LuPnb6OAd3eKrHWS9kXtgGl7vivNOg3lztJ
deOmqAma4uB3BcNoRMcSz5pTbr5mr4hO+GPFMfiyF9ID8LSMS/o8+u6BvPLAAv5N
AUFCuyABR9I/Jl536M8E/J8dJTZaeyBplruEEHLEYtVNJlY4O5YxMKyGpW2AQIG+
yuYLpEqhp5EUYlE4JMPBM4eL3pUEmsmIDSI+H0T6I9BDQ2y3Arou0zBVHFtxa8gP
UhSUjC/8rzbze7E1rOf2CCsx2P3dSJzgD+66MLF9vKaQunH+PZR8NkvvzhoSPkYl
a6+nhl81G1jItr+SdIzEKjBE6dupr/14p66ySMy3RD3M2taAmIWb6Njo55ZIBSFk
GT1rRu9xd7bZIrlnYWPvUgH3qitTT0vmNQSM9lHq2zEgWx72DqgwGIhNAZvKDQp4
RU7iBCfKJW0XZKI+1Xc3XPnG9DGGu62GwHXBNFx/+SH/T1jQ5Pl7akmVBuD1u2WH
OnXQTwzAERrRxcC70j8OMn6IXWc/3z3QOMXPvH17ygfZ2lPD3jLKIsFsN8ToRX1U
xGe5Hmds0s7NFE+U+bc7TS8DX6wMKLneDh4/DnkmAKU/09nsXsKjUQAd9sfdx1ds
cgDIepaAW3itiahC0i6XzSOizEYx3HEN+t6gFh5YdDMCqHFnR2GXsBLjOlyqw3Qm
pIPLugtthuXT643Y1jXZ4TikGkOpmDHusuPbA2DAAhrMF1uKRe/zPbtunGOqeT3p
+++kgPSlAe2mNd5w6K99a+BjBjvTJNVmhM9DhMsjt7jz+7Z9mqpp4b2xKoIfaRAu
X2wBYB6XvoO8CNtX73WsBJco93SPIkNoIURjyL8scww7WjStpxK2mQUy8rMDAT/C
1UOYcAh6TvVCDgziUJCeiQc7NlIbSW2tnLfBxArS7Y5EAIpRuW1GsBTRUYYyoEeB
APYYtX4/LEZaOCDKNvB+ew36Gq5k4EhO8/ZjtMchBCAmR+qemI+0ur12tDDDvnqW
+ZtXJXVGbHDeaKCXEstHKO20d7MYLAdl6LMXNZMxVboiYX+UwoiwVKNPtv4+sWBx
fE8fC7obyXFcH33IqtyC0o1jdGBUcrCZMTLEgY45NwR4Ew0W+9kPs95hS5+X99DW
BbQUph1LXuUSK9L2Ov3pOr56BYh57+/Mc6mV4Qln6ny72RJJrSeTNIYgPMEhjBn/
13aZfMvDJqb8Vm3GypcnIivy09ikxX9l6inHX/yOOBnkhzSAGSfBKSlQNGAuffDv
N7Ue/iOV+HNHOHsVUQ65EfIH+qTSKSzaR0rGMxXvtGMFLVfrXSzpd0QAt1ipugKU
CY6sdk3jYxblqsBJC+mzExkJaZzMgjDszkkdsUW18zO2MXcpNkPplAvnRHVAIt9q
8Wsr/PN3Pre38p+1kqaJ5ZAPIPQqhN8T0Ooeu5ANnff9Xq3pEowy2/NdR8Iz8gRg
5HYJkOOh9ilQc3RP/3HXSgLe3iJgwe2oQ/eJBFz5y0yrinB6FVoPOTvcfXnGQRp5
Xj6CrU+Ln9bEuovEGSSOkw71WxCnc7yQ0XCWo0JsQoIYyBV50l7W2marG1Z36wQU
03DkXITGAzEOdEKqPIpdPm2Q1zMd5mLVHNAgEF3CiOzYEcOt74n3xM7xctzKj+Wm
MqGINUBXnAAlPO4tnzb+TLmjA+0TAcjN7fTtDldDCWaS61VqaVkGfLvr2mfA8WK8
+RWd46ZA2SwLfRXnkKD7v9heLkgfIj6Rr6P6BxYmjFCLtUP+25oLeXJthYQKqWeY
YoY4RdVZWaVu/g5RTfofly3OFzb5UkzCLmZGVN0nm9WuwEZeA+klwWii0omA3GKW
24OSF0hVvhapPBxWZoVTxT46odqf9vIZ2xcxZE8NRLBr2Z8kSznMRC898COO5bQV
wzMfybsSRBqFD8bPpO0yQWuo6UQukjzQYDs94fHc1VLhfOpDA9EIqbzipqXKNLbf
aghmbmIX/1leX3XYUN9063qhmQVNCtyQpxwQzZt8RcTb8Gp6OrjBwOxLx8SYznUF
HOpM1/sWork6wVN4dVswiXln0cliRNu2bkXKmSU7NY496p/mdlgpqy4Pz9DSo29O
7XjoqSxz/f3EHsSSoDqkBQPGp+G1G8U2b0hwWl8hqoG92iJltDQlXYKVmMKLXKBU
ryZT5B/8HcuK2GYOp6/udVwPkq0sS4qYZFvyZxMlDPMA0X87QercoFP2iyp2uJE7
DX1MfL332+XN0NzuLEDdR2H+0/Z4Zti0c35hBg+EwAUDCcW1/slyHUHkWyvcGKOY
MOxCFF5Cpd/7KODuMTOFm8uyZdm2bjT81gZnchK6uLh3dWH6CCs/eLxvwy7U5CbM
MaCAxfrKURNmvgP9J2STT8iwRIEIGh1NORHCqTGf37qgnRRXfvgdtg5F0C2zerUY
rWo3TS0rJRBgZtbv8EPjaEWcjMXMrzD5bQKDgj6zCRe3Bba+bvh3xTNR47jE0NWT
3RvjeOm2hdfrvFtkx4DS0cA2iiavN3kteia6P6bVJ4ngAZ6rMiIV1TmpCWWo/m0O
j5Bcaya5jIi9UIejDiva7+/Qtw+IVhulJB2MSzwIwesQ9yi7gq0jrD9aqYFsoXVV
NZlN+65hByQaHutmxeViBe4Z/tzCCCiAghr4uiEMdEO/TAcU7JDBbREqGhAkKLZg
`protect END_PROTECTED
