`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xY9OK/FUDNIkx1+ci79NuIV7FZXAgdebx9CpGnYnpqJNpMZgUbtNGmgoe/XeABbV
ffVvrhGOENUj3YKWt2HIKI95xFcbDyC3jPdPVcb3vS71rqLfHkEAFR4rqnTtixaD
sikbDlloGk7cxVwnRbxIO37ZY37/2+6QJPn11Pi5oZ01UT7W+nDWjlLXb6lbHyHf
N1weIpSMosWISWLbYH6tFfiCNHDtSTLrbJcK+F4sNTC7Q4b51Fyz73O7iOrFbcap
VyrrkS0d7VU5pLRMeW0lBCXsaK61xRR9v/t05P41gDONbo8pYuoa1E8nAM3w61QS
/RrNgmZfAKIQKCZ34npu6whp+giB2DRsoslxJ9tN4nJZqelU0HpDvJrqgAoCtwxe
CTNECTuphBAI2q7CFnDuHMxDKW9fllTfNSeHVw+3z68NACbqU1pDKedrEAVx3jbl
Asq0KrjWBoqi+mvugakwkiGPfhr+Zxp0L9Azd6qUjpdu34TEB9t537M1vN37XT9t
znmtuGZ/foFCruvhbBQC04HfRBZtumBgcqZ+9KNQIRmm/zkVmWpujE+LdoVwsXNw
xiL5laVMk1ghggYkLnBWYcp62GvIBkqQf5xwtHgD8RUFav9L4in0f48mo6juzIh2
FshcUGag+HiIhdIGafcEhYpcY3C70ZibbwdT+G1gRJ0XphUmq/eoJL5+fNmmMclP
bkid4HmeXJQsMw7Rmmqg9G0DeqnCgBknsIa439A6WjtK1dhF1gkF+7RjwLJ4Y47Y
3VqK135f3vYRpeF/iAQ3dhUPDbZPoykBfVclNHGXNut+PdxMQHadCkBbxtqgcnz5
F27MlM8cVCNsadL5Lpe86lJ3UJTN1cq5QGTxv8tXrhtMObyHQNX5lwKdqwmM3v5G
PAfwYBTWupZKdzalWwt+IwrUWHz5lE7PoL7A2w3O7jxy0tm9TMIF1ptkFL5NR+hM
KtGTsyUFVE8DKVW7B4bj5TA7FYCzEQhKbrGW1Dc0KLltdTAI+/15xM15FCtHHjZ8
rsDWy7RIsi0/hBwYJuOz9m0BgCUyuGP/Sw0X4CqowHTx/JNqVX4SNkYf4blQuFBP
/gj6sHarHTR2N/zISFsvhNSMPSlFuwPXN5PvJ8EafSGfTKmqcNnGdW7LD/gyQb9N
CADfkNzjJLISGMg5TukPnmBEq08msHWVslvXUBWT6tgmJymZo6wjr3f8vRuXPCBR
d2ORSdJQXvJJ4F9hGDs3Pxvwveg7cGm1SM02oFFGOjEVKvvI9MwJEPH4XKr6oMU0
9VlyPo2qmnFfiKu6njEc8baRd6yMk8xQZWEnRB1PCm5IQlk3T1A4VcqKdOC0qljh
BGb+qOmKmThXXnSrL2zZyaoGY0ZO4ARlWpLgkcBLyK6hXh5grRFwJOsl0Cgntz2E
yqFBWgvQWzrypWS5IqxEaCUisQePtbHdDuCVcfnGhu58SeRzPKXRM/yob70HKFuI
Xfsnfmoq0EHlhSEM0DjIPDPTyyewKYdY7fKoaiRFc0P/JOoUCEy959D63MXguRuS
lKmfOe7J+5wsBIH3FqDQOD+FLUlxroPJLl4unXRF2MxJD9NyIBAOwX5qOU5l4tV8
8Ln94BHJPl3+npoqlr+x4Eehd1xMkcviwInq/a4ZcfbhdkOc4h4FOY9wBd4WlASv
aCgsVb9UuPKGXYhTMFRvyQ6SeBwuwVpndjCN8OUcy/JHetfOirmDV/JQ/NstC8fY
MYyH9NBv4ZMbFfKMwRI3w3n2SQHBJ/ebk0lnmsXtEekiicZL5dhFz5POQen11QWM
zRqSEjNQDoVFVpbsvsJR7TU9bUmZgzKEz9NAE2Ylex0gkP2gVNuLE2xs8Wnw4qMu
aBe++ZWhnhGXHbu8RKw3O5wnZGCWRzJk56l4aLOP4lOzA2kTWHPRK0Hpcn3nmVBs
Ljrf0AWLIsJl1oYR7NwxjuhB9m223Qxcwop+g0mJklxE8oJOuqNq/EfpqjNABUkT
AL9msE9g5HGQOOfa+/Q85SjK4j770AM2qWOe2Su/ydaFpkAaTnpjsy7aMrPYIzp5
ZePJspaKTrfILYSu3nubkiPEl+0F7PWjjrfTP/C2SAV0ZtyVWNbYkeOCxgq5MXZM
Q26XPNiQX5r5e2IFDQg2ft+YK9oBFsMzmBX3PlV3GQqHU3HbC6Pij/29V3k4Kppe
ckJIRIiJGnl0xqHOZ+n80PKLOMa0Ch8v29qdUTg44SjNZB+en+3bvE52jQViP4+f
lrw/ISquJXmwH+CDZscbG6uyVwmeLuis523mTMcY1R9LuAM4RtsBJmmBc0LBo7pp
UCPeUHGF6g8BGeJROwUlgECv/WpjE8P+Mxde0AflIa8A5sNIKyiKQq2+Hq0lBh6x
WvLmSIKSamDAPmup2WnpMeiwKLxdHJ0jKilDgzMbWcAHPBk/zx0g91BLg7OZC3K2
UMRizEFWOE2XfzPtWrkSH52qRU6EQsRDE4J2C1Oyot20UeP4OJk6n6zCYXr6YJzS
zI5SVqp1fWdXyjKSIZZbkNd8vZXPoASW/OFYyEUQEElnyLVS+m8teJjCwr3IflSK
MxXQD24OcdTZeHpx/h0mYe3CxRrK8Fiada7ct5lD+CedA1N6WUIXKziAxZbou17b
zMNjjTp9wnxtrK1NRsSh3veYVGyA6j9/VKWAdXnqdEfLnXrpSyrP9BQQpGSzR0vn
4lm2EnYcOiu0S6Kt38ewjRAlFsFVy3TwhS6g+d/QoY7nvfkvoFUUgBVtwcES3Qm1
AmDh4GRsejR2u2gwxI37uedJnzxGDHF6qODtytIlIKvvd/kgpbTJ6BdrsNQhsCeQ
h/8y+iORKw5xXg+llpFLsecUuJk5JJFt/C4I8GnP2arW9wiikoeTllsXNPi1EuF0
4dhHjHVhGCkkJffzlS8zfI0eBS/9USmi6facRiHkAeEx6nJOxpUNLDD4okoDOaXe
DAuae2P4i7FtMLII03DvQYtVADM3VEy5vOO3BzeDL1n/EnijRKbZJOl5SRRyE3uo
9uYh9ROGmZQNkGDDZcf7owJJG9dHf3snXykH7CmGsUBSHVIwIwAq1tkklfr9NRSY
HVqWhsVgRKn7QI+GHNN71hvSvmTrMKDRj551JUE1bj+Wdw9ev7AreTxmujwvT99B
9KZ00uE0C9MI6wmVYgAYkFuQtTAOrhAYzzxKU9Tcl+084CVJnZ+tYjcZXbOIomSX
zU+B6J5mmVZ8YN82ajyZQ/s3FhZJiSbqFqmVPWZMLHzeuJL7GMSHERBX9/7Nvt+P
i+Y3hX5QIOSFWMXioLjjdEXYpnBbHXRcAlESOHIee4afhrTJCkb1I+p1hofyY22Q
NwKOgvWp6cDUnJH1ZOLnUm28LYtZ2V21by9mQbZtKNUvRfr9EHlZa7IB205Up5fF
K7lPM97+Eqq2MY+ureJlU+IvsCdJIZLo5fmRoba/wFvAswGrUeAvYgxAcJRIyuc+
kjTBtal7PA+XSrRCIE1X2bcGyV8eju5Ky1xBGcovLJTQAL/G4zGhEmCnvXaGymaC
qrg/UQGCv6EsGw8fRV3pSwMUODbiDPZ7Ja27n4RE4Bpdt3oi3E7JAUYsiwpQjQrY
obpHP3LM5jKHzNfNY+uqEIDJOe/HxjISM42H6583B60uZ/ln3x5XmrZOCWRW5n5W
9H7XLRgYgc0GKQzr+FkR+Lxghged1b02PhTTohmxtdXgFaa0wdBP7hdBGS3WDjak
JH2r7JUfZMYtpJwNU6UVAyDZGqpP8lgpXtO7n6bDEP4sFqYOQ6yVvV8xC71tmJz/
b/Z9iutka17Qapy0OyLpb6W/H1ycSsjsKv9NTXDAHzLEvCDz849pFe+JonPLg3/n
tLMd+FiVU2OfGg0LrRIHS11lWWpWRAMprTweMtVBTkUNFK47H0C7K3gB8KFArNv1
VVqce0LGuJaBV/Mo6QLvTOWhoyrKFK4iUbTeHRQJ6mHhJGI8EeN7YzccOTF2iPsk
`protect END_PROTECTED
