`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6OWDCvypcOT+RrZ5oOz5j6xwUtkuhiSCvMXZ+c7dTYrVX3WcS9m1yJ/lDWEgslJ
AiO0rqZTj+cCcOzdAnRR1XLGUKLPVS1UxxD0j7adzBqJQ7fKMQVysLUZL+3jdBED
+C2KeTm+aOM4T9SyZLevj3SStAeSmqD07S+QejfvrqLoGBCpFDZpODyIZkscefKe
CcsgbKrx3gm03VvzRQWfKoUgM6afrTleFk0U+p4qYxmBT2eP0DduakwY7FpYLxgd
UQUAFzFpfkfe40ddqRug15H7LaB+LwoI9IblG9OM3vjjmHiWTrcz4l+LRBiLcGfy
oIztrqamL7LvtqlEM7+qURjsPdIWxGKhpOVCfv9QaAIqF/LzZ1Ahkwd4//tCk2CR
jM14WQuYVl7gzgY3evbBb2BhXhZ2GOYRGBDZl0MqzddTn7/hT9EKq8MM1JUs9lt6
7efiq1OZvaq5nU69FkjnjRucT9IP9myjRrrzvvqOI6S7o+uYMnJSLbg9V4IurSX4
NVzM9pslyHsw0WW0N3sHbsf2ixCADxUfZyrUM+ztSnhuxBvHGaVTBaO/lEGM0eSg
`protect END_PROTECTED
