`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POVM/td1sIl/d+gDvoXQqlBH13DBVXxfu7Oc8SZtWKWpr41jrzo1862bsqXUJwgn
tVs6vWq78Pi7AhmAtjOFtvlftrF0PgZ4+SVaJNywrpe5gpR6AdxUZtP5+0sr9OH9
Ly7thNh3W/xJYBMOId+fZZsIkaBsdO4Yr6H6pR+OLK1/dBrBF2fV9rwyyF4QFbvZ
z9b9RkhHsBOaKhlQ2ESkHDSz8wkQH0VcrCoQLC3jbRmrC/K5PJTBYn+8FpD5yIBA
xiQ2j6CH2y0Nf2ReAWSjauNTnGdc0LvvK9Ba8XYWiWDDQgrL8vimcJQY0sxNJfHn
qnNOPS3THVr/LPwIZcYbavVRePuv4boQKzxh3jpLAXiPPl41lToe20p1B5/jr5kJ
`protect END_PROTECTED
