`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72zw5qmgcrVl+uHHoG76F4KhqFPQkaTQmgDzzL0iWP/wszqbJOgthIKeOM9l64mw
E7gDyIxHMqiiC+C+mZDf7rz271jDfUcUclBlvrLfFTTxEuYE/k7k9BmwyUoq0EUQ
EOLv0l30AiW7UFsXLw8kDrmP/DVb0FOsMaFgXgoowPQ46VfvJzKdiGMhC2TG0Pwi
hzzagWCJ3sVHSv3eCvD17WsBc/5jCCC/eQlSSMAops8dg2ORbM14Hmrh5eLEt7J5
il6M6nYjqvTzjMdZMUqwx4DvYTVUW71Fpfh3Lci3z6lwB1aIYsSURRghmbvXmQKd
Gp45K+b8vQYXEANIXkmr0+0kEPgXapHQ9SMxHidpJbUTaJNqPqCk9myjHtPc8vN7
mdYa5mq0Vy9zbpVjeALuTdyUvO7glsZ07MsQF6cXfMtMUI26eGLhjASey+G49VrM
I0hYn1LAeRg7DjRpv3Pdk+XkH08Jw7tWs0qAIgvHeR8VKkzp9gY/GHro6/kRR0Gd
YJSPnBBucy9bzp6w/lZtQGg134/5Hbg5DVvdMbPbaCa8kNzU6Gl/Nr6Z1gRH6hXK
HqZIYMIuutdBQi00B21Plc9w2EqHKlQy/r3dVQv0VTxVusV6rUAfGICdkGjt4U8d
LVl+Zirm4MNOAeKoHqjknfxfGnJG8wKmPTLereIezwJ3xx8WjKWdai1eZOWPKIVG
iJ3Gqsv5qsfUu6IhYdhhqPSNcDiCVJtwBMpEjDHYSwiPa0Ubtsq7FiC0/R90J/+v
zNxJICIs6nK7nGCakrvG4Vlipk0BeXHG806fh1txqqMLUB+1zDB338RGtqAkim3f
CCxiUiu3i6y2L0QhgItPpg4DAoiKM0kYsTuU1RCWMDB2PNS+i/ZJF6EF6uSFG1sI
ibrR+n9FibRSVhRjJpG+ND13zyjBjDCmZSdpM2rCdL8JHySOU7cpPMYbYsGpndO5
nY8sUxxhmIXFuqTete6ttk79NpFL7HHKW93F1gqWlqduWKjjSEC31eAzg89sSaA2
pIywRDeMO3rd4iaCXJuNgzZUerv/fNryWUvRg2yWLiR3/PA7OrfT5KFLCVJfp0zI
6PEUUIIWhh5+WUQ4f6VOnQJw84jeYl6q7Qv0iqQFjwDTpOoX6alSci3QnaNEvy8B
p/V58BFWrBjKnA2tk7B9e7jhVPsNNxKf0WYJf7L+KyCW7F5EPkHHpsEzyX0TSWLE
7rbhhkIpeIC7iyvlALUUDUckdEla2vIagN6z5T6BDuAX1QnW7GcjrqH8jMfc/xuh
rjitlMOxLnS1n8+afPJi63TSqrZP2mrkqQebWcCfN57ieLpPC1tB0wYBo6pgVTQ3
XGle2cknVLqJuPWbgCWxJKQ0pBIsHBf5EN/5JqAQ8QrmAOERjVgLxgFYKd8tSmVz
QiSkQTnpA2N/sBkWy+c++6ZCRrZSutFljlBHRy/zJewx8OFRWDLChNPNipRP9k74
ZwB7jw3sZ900ur8xxmotqZ0N7mg8SxBpvVQVfj2LB6CCX22JGap0/EBDrSX5l6vI
+bIiFZLwrLEd4is4N2G3cNMQCKTJh/vOiZQ9MBQ1Weoj4XgCmNRnSXW4MrSmPbW3
ZVapd6Zs438Bv9ADHUrT4OOWeaM8WvkVTIsNDNbhraYIrhae0TDU7mAEstS0HR4F
nDufZOxe7fDctmrLUxEVylkuON18QPwuN+XBIHz2aByUsH9Efr3U8A/qCDh+jmUN
0gSxmcfiRPZoWzl2LedfGoD/X1TtZtAreF/isCEYIpwfHbwNHp3J/0CKR1jeRdrP
Mz/I4HK8AwL5TBXX9y60t9kDqgyfMioqtE8e2e5mA1dcMeOkPzmUYgeKBwgvKpfl
uQvxFpI0w/mgI6sWWnxLC6adXeDSRDBOImpL9Kr8Gqk2Gk/O7apCHmo6HcXXnuWi
c/miD0slkk1KYWbVW1dXF+W/0moI49KnP4ACMHfbIEPEC4qQ1yU34fiWJcpnExmA
UElaJSC/S2jLy0cYZh4rSI4zYqubgSVYqzVhvk8ap6Mn/pRgIAPznu4MPJLoYRA6
kg8i/pSccF0Z1O2PIhD5XQ0A8mQcRDKlb2doDPo2JGqmmo68E0ErX2fSj38D+K9P
bPK8biEtvSSeN5QUqPaao+01BefTZJ6tcwcgDDAuOZRo58BnM+XgVXGte1RNw56D
3G2jRmrjMB3DGCPWPT46dhq9mmAV7JpcArDH87ftQ40RSdycpbna088v+34/3U3g
OZ8yz7WngcS3vghzzegbBemadhKuD9UhSLNyo/izAi9UNxJV3PsRlvljWvOPppFs
Jirl0RpsfMf0If6OmMvl/hckSs+RxbWRDnVIuc9KnP0ex1AgLo7tkdHL6I3+ooMh
yYHi6dLM0Be8zW6/ILqTLkprCcaQzOTMg5ueMZSh4sPtT2AvzRmXRXMRnF6i4OB1
zag94zwpt2HaQj5CAq1IeSYQtuEBG2mxn33pXy0aoX+9oC4W8stZTR9riX4vdCtN
5k/t6iE82vycJoeaF+Ho/48WVbgZBl7XRTqXFgO6ZEMr+Y21iJ7WbSgW6CSX80bB
z7K8xI7hQVJIhyxSFyWqCisSZYtaVDL6ovq1Y3KWshLn0D8edciG0XghSVLDnOPV
RiOiyp+jx/qx1V+1Ca0DsR4bgYV6AwBHiK4vPbDNh5nbopzPhacbMRLtcEzvAMzE
mHUWtOAkv13Q7OYj3oOMNkgO6eMOF5tmMVM6D75HmjdQjmBoAtGc8iXSkZNp740i
hPf0RjGg2HtyIXt8aan3HWZ8xOULj9z79ngWW2gk1GmmTjEEC4E45/VPLl8G8df9
8euFpUL1jQYxul3cyTEtrMTcpoKglhKBQGsn8mnze+idkvJn9EwYf6GuD2XJ7NON
1orEKYMkv6xOD0h9/1TYZKqx2B5jda0yxdsjvslFoQC7j8LUKrYBzAO8MmnvOCef
OLRohgK2eOK279S4zAdQlQ1EAHjN/P4X5o9uB38gcBmS1/Bom+WDUqUBElOo0Ck9
Yff1Ee0HR0W7VCdbFlQ68il37LJKYn7xeNGkBEmRFPEBzyM2sHn+QU1x2vS8YdgV
aNjlepWatU5dOCN/0Opfa/r3qPs4e53KMuShOqGCZ2Mh3LM5xHf73+FUcUrfWV+3
smgYMj2DHlZHWY2DFfbQkL7b5njf23U5Kj2MMgIuJpqO6a+MdqjNSBFEj+SYxbxp
G8gPMBEZZb9OyWkDZceSAvQ1PVelNGcBrSHOtPpU0xZgLRaokROW8cz8DgjLvLxJ
XljvwV8g4mK0xkJXiA/e5VIW8iLQ8m50qS+QtSM6jq/CuWs63pW3MTdweAlsOxnC
sSJhkbTL+b+Vd5YsucKpnij/4pteYwWVVZVNLJr6g3yDC2OQxfLsYUfKas5mK2q7
Av0cjowXkNRNYpR1gmJjIchUpAnoKpiP9iKS/rLvLW/pz6v+WcS+BdPk+Not8J4M
oReIGreu3cOjXbwFhSVxwg==
`protect END_PROTECTED
