`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbsA0osxMPAyvA36OhIBP1wSWiwy8A4wHJvSiyZ8j8Dc+e54VuCQ5rSaPDr4rQaH
lgr3iVQTMtDnWc40SY6McMGPk3wJsfK+OkXQpygYj+dru9uyx4Zym7w/NBrpeO8I
osIXGNARGIVjhDCCaEzL3GmqDxWwqFVtpIMhKbqUA14M0+/XZY20KlmBUB94SV6x
PJrgRBaubAwFZcxXcq7pfIF10Vc9Sw6RVxuWxmFSkxwkCq6g9AynCbnS9lLov8l7
l5b8SDSlNhYq/QXqnJtO2iAjxO/WxbabkL0AzATVAADX5u6FTOSz9wrMlMNjqkZ9
TMCTIqhtx+5H7p0jwKFPnQA3d4ZZjiS6Xneperiov0ixduDhJkIdF2gyHgHqtu1T
bdIvAmn2REZvXR5H2prYZz2tWPmcon9FrMVjY0gGxzNtDn7MdDogOkR3O6CJrSoI
3ke62uTims2UL8V/x2PkhPRwsBOiUopKeCWeOgH0nYpDYqE937Qk/64Mtmbtm8UP
LAHQ2b3K7erPNzIZnL3uVYh6nzgN6vKhiTyaYgjAyN1BRqd2QvLtfoI4VDiWwon+
vvwUr1sHbF/WiZB8WxVQ+Km2euILg2sXLV3Ilbp8IeATnhOdSz2NSaXAtxSbhlQH
FeKqypKrv/tdyAIaax9T1R7hrwfSJq6EUHNv8948SqJ9Z10brfN1zpt+eI6niIPn
ZkMUoYcK6nW5efKMH5++e4BXpWgvRgtXkGEArEkvH2C9lQJQzw51uWx/CEkQMOx5
9t6naSeu6gJO91fK46IMtY02okUqBkDzdpep6yR73i6Pj+yECzS34PAyx3pjXqEJ
Nxv8QSacujVx23uOPcvZHkT5CEb3HZaQfBy01G0LMXyG4ugXJ3rPc6OYkbJeNlvK
0K6r8odEGCiF7sa7C+14waIJ5vh5Vdb/K9EgX2SMQH7LRr2ylxhfuqHqU/IRos3g
op50qN1q3WyMnuwJutZ12Q9w0uswh0uHqtbnpDnQ/0AOHBbu5m5xLIyOP5l6xq9e
0z0HmE27xTJ8pFLRxnEwrubJis+bM9Tk9Hc5HNDNlZTDh6qTX94LjrvsO9CysNMF
n2MA7hLpS6EM7d+yU2RXBC+SPSvUj4f1D597N05GUxmCNXfonMfrE+zgisaqA3sQ
7m6F8B4yLj0GY82Wt6VMKcOMcB7qTC58h/6TDSUM6ixtg4WEkwrsXDOf0UqLb2s6
NmdPHrocKuoDbXaZeajuJCSvS3cFlnogCeeME1uMplqGmz0X0g/6QN+OznzUaknV
fORjSpRMTgWda/1lKl/bjeDQZ3+zp+89267xbcHmuaiHCfc/IxL+1WZp4moPz+jX
eoDqlkMz51UaT9HnRn636uaLj+ehTOVqZqG4SZIsqTFZPYW0HFWe/IWoLF9LfO9A
d+bxQeZ8XLq1DvSrL3bQO5fyzg7KIh4Qoa8HizcNuoKS+QofZpPsQejiVFULUu/G
UpRix9093ymLBOAU5L9dTN/pHWP7ZAqeKoiaSqrSHyl0qW2qPbj0KkCzrO2O3bnF
QnO4qoHcTp1gq5nkvKer+fHsjZ60kThG7UUGyzxZEBSTJHHL4Sg4UAMjtKB/M/GS
dMWIdGr+mAsRzFN7yvT4pSSS01fL9h50S4NZBH+1w2eVXcTZZdX7xfW8Pvhvb0O+
GgNywPbbGQSEu2kmsSwmu68e5yM9Fe57QS+fXCZ/31X7CxZHjlgo3//0iGMxEzXy
dpdCCnyMbfMZejAE/njzOsvwlaGDAnY0bZStocVKachvjGV3zKWax3VmwxlL6uh3
rLUineajy6+nizAwwUkRddk+d6gqk8fuogDLFAb3BFs=
`protect END_PROTECTED
