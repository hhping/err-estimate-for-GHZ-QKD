`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdLMYPNXD/wYn8KDBFI95P6pnBKCuo/YxNQ+fQ8qFimMGNEUjdV4juY4yvDHDd9z
zb03WLrYKescJjURhtKyk2V2s4neOYxExvRPDHwf1a9CnZwMcpLNjo3n+zHPH0sL
LJSZ84EMWDOaFgK3pKJSZxwIkEYFDPPmhfNvGBKY6EzYf10htGtaY41kRyCPeGfq
j/ORJyqHtqYvOAI/N6tr8htCGvv3HW6aORuCN2sVFb6VWE0yR6gDyCJPvCr3/AEs
vgkh6as5v8mOwS+J5nzG8fydVr2RbSlFdpCh/AISQGh326+T9hDEifZozZfiGgt/
W9PZt3GInWByeIbRUQLT/8H6bOBiXoQMDvPM0VWUlYdzgF5vjGLPRQZX8GqwMi+P
hl2zJKrCUWYsGt/kECVq080ztE5hcLrD/D0QtLDD2wwKGBrOHogi54SKZYQUwZcF
X9aEjn8S+96mSW3UNrjfaaNXD+lr9nPxy5CuZv1PlraSS42pF7RV5EgzX/GdRbBE
tjKHFEKU8vfxPM8POG1l8CfOUSXYNnEDQFXmGN2/Ko0nRh7MYXctkObv7XX+5dLr
BhHWQ/N64QMm2SsY8rdD6k8cGfhOFmhJX39EyN3VoiCjvq790v8UG9xT5Q/gR1e7
MWdHydgqncq4mQLl1+ViDV1ustZ3dWcVlzLHhEFiCjlhJy2y9BTrpnKFIhrVosR9
F43Q2Njd9j2pzoGaZ7Lfdv2abGasv2U7JxaEuHkjV3MePNJeawRKBU24Yusu5M7V
/yszC7A3BdBcE81iMav2L5TCFUkaelDS3UY1eOGNilhYC/mHp/h8WP7WR80GDnq1
RbMZQOqxeYPtKJcK33g/o2Nbni/+YwIEQ7AVmXrEx6sFfB7BxVcCeEAaBwKyq9jg
1WYWdBQwklKDIP2EUwFK0jkDOi3rvXDpjF7P8jcPASji0leSZroxnARRuzU/wWaW
tITTb7qYpOczSLFf74vKZAr9op3Fw2JvFbRvbirz1J9mYnO8pks0bG4Gdnd8eLWp
MamzhfNxxXEipLiptoH+SRWGOQBrKbgQvI6edSA+TILwwR++zaoDN5ZB5LuB1U30
tChJ9GYi51dLFQtLYyUcFwcRVZrz1p+BUEPDAENiJYIGZH8zV2j0RH3svux2OpyD
lb0eCCj3tQ4q1wbrtKmcJqyyBkMJVNzGOf9AVdrsCOM+7yTsyC7CITMOTryWvjUQ
P/f29yiReQUYwGTjaWN+iEiSiT2vx1nLazUPxgwZz7lgTAnqeYOyaYrL2eZGFERj
vFu3jHC5ZRsyuW720vrIHQrsYUk6LLM5iSuHRubWIKM7U50FJYBGJqz6VLVzU1aq
1O8Cex+Zfx6/Yfv9Fc1nWEhW9D6+wjtXpeefyzf9psHm81KB+AIguAC5vzoZGZXE
nL8MyuvQRxTjEF4qGRgMHO9WRX35bOz5otpJGZOoiAJjiI6npEgZz5aokukZT53E
jWzJ9UD1R7tHaODsfhOibPIkm8r/T4wNTDCiehWljOlFCz4e7DCWRvkMRhtW2ujC
evklayxMwGbI+arG5yJDb5C/BxcyxTWrm0qrDAawggp/kElpe/GNxFpI2BztgKvB
F68o0CNh1lXlwrD3WjwRkzT/P1AtBW+KdhBygiy6oDyimftdha/OzMAnEoDye9sU
4r+Ia3HwetiBIOeKjyAmt6KfnmCaXJqJtqlkWVm27utoyMt8snbLbZ+eO5nAL7bh
wswgU4p5eExy8fXmzpS+foLifqLHLueCX7saYlGM2gIDORia/A3depo8t6k+GywE
9u6TifBHu8foAlOaQDrJAWafIXGx4JtMVYG8m1Wd4Asf7YWZHfvpIrE9vY3jiaJE
ACzEMSVKQskKdpqoIYmhykVP0Ap0Po0GeBBK3envA+voDSk8ojZqzS9fm7NrjKy7
iuB5vOYZWcjw1PKg5UpRCPHt3Xq6vq2bJx+BcW/9wktldO36LhVeDLFf7qEaeDcP
8VXQGcJ+5owkH4Sd2zcplfNJLXWpYglqqTeGLAXuT7HfHY6qlNKo8AzXtL80TIPR
YM87c25R/P0DOAcqpTKnyWUTHOubTyf0jiDw4xtTEKkZzLNslTSekks8FMGH9fm2
iI/Cybg19SPkIN95SRMXBtANam27dS9hVlF2HWwnIW5xpsxKT7ifgzFYNe00WIBN
WCcTnQt3a7rppUsrVhVVcXxB+52mkQ2edsg5JokAcORClMtlPrbb1IE6zDvd9BDo
RO4XSuqohRXkWvMyhqip/sCbP+UeUeJ8asE3+DkPKPY/VfMHtG8Ij34mc2rGqj2V
tiqgGpVEECQC3oa/nd8xfC0eieTuDC6+9FKkxj4n35Z0P0fIX2KIPJlaQ2LAs/ZN
Z3UgXhCc50v3ZcFthcE+hQY04pZv+I+84KE+8xCxFkSgMY5fBmlcjLUyO77AKMb5
biAHXPiCzH6OL/21DYWGyl8KMBe1gdAYevFUApNRMEiJWUUxTkUu+6sinWwJ4LQe
eNHVnDTlkyU5x6Msbg1546JVHvHLpVLU0w2hcld5zIfFyxXwhb5xf919KdHnuDGL
lXAYD9UesTN/yw/pfYVAjQ==
`protect END_PROTECTED
