`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLE+xY9O2Yrhej2nTcSMdCRsOtgLPLpYcIgMKZncIfj373ETjoU5QE9O9z0UZkTI
FPl5w4SYBtcZAkE3c0TzXt7bW2buBYyvEKLbeFwYHr2+G0AkgplJr1EAiLYPnyTh
WMPvmL1z7ZaGArJ75UCftMKde6nuH6HJkbQAQKPbQ7GSnfw87mnoTGryF5MyHkex
n4M6fErvAiBi7a6tIgtyjGUGjzqtXGHSWNwk7Jy0NkMM/TQ7NQEpvOQNGa16cOPb
L398xZbbKdEt56EkoOdHRluOjYdila7HYQpmite7PMhLt4uDtdcIHLksdgBL5D6+
+YNY8Wtjx0ia9fXQbJGwOHNXRcbiHCyq2bZfcT7N/JbqCgzHyvTbK5Crd0PnXxFz
R1ZZcCQQy55oEonm2GJx8ZyqDkpsipkiqnXOyhLtZ7jr+wAEaOReFl4O5Z62WnSD
Ox9USVbvdiGzm6XTJiI2ZXISHDTdhOxsIJpE7+xTd3/PY9ezJnOfHsMsS4WeFv9q
izsFjE0r6A/AyEsxajJXVw==
`protect END_PROTECTED
