`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UdrunPIthDf8HRN4CAImDzYPSfLu9g2MI6MgZU52Ki/mUfLHpVPyxs6uC95z3cr
vopotVnmUOmQ+eHcuwKSlKrJAd2MkOrI1Y69xu5zFEz65lyvvrhF5T1I/QSyV4aQ
TELDXQ/V696l7gu2xxtWl/EfhJ+18KmsKJ7c/Cm4gmd4k7fx78t16ZWMi2NGA5vK
s8kjJwJPZf9QJIERKmpgogX0SOCV8Meg7c5zD5kBUza42Cf61sWMeWCGlcE3ZKpF
P57RDSpS/4qaROgsKwiehC+KlFEBGqUSVS11S0vZsd5WA82F7yOwmRD5IhTEKSzo
oK5br3V8TlargPXBxfaNQPDCXCAlEKblLMOQG68DoXwbthCjHX/cE4STqOFvX2Z2
fgyG9wHNJJywLM1KUiNRsEFf9JUfnnzV3K4R2dg9uDnfCGSS9WT4mVBwF9kk1ZWa
PBBJ8QkOgewqYrXQ3MMvIXTQI5U5kVIZhKyji89GRTJsScaLa25417TYiSnhhwKR
x7DpT8RHH6i8TutEjrfs2YpFlFQr7SeooI9Bo/xevkYuWM+pPGNonCp2OUIdHlFp
0583KbI/M3EIEfvjdlsEWw5uTwbsWs5z+X4SS5jVsdtifMwkUcP2ozwSpzsFuxr8
0Nhe6Ij6l5UxRyjgUzNDuQV5mXTt19WWT/eZ3Hlrk8yYL2wvDjOX8Vt3sqNcbXUS
al2jxMoYPMaJrYZ9/yIvog==
`protect END_PROTECTED
