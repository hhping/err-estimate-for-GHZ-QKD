`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+CUL4PfNGqASpdmgI7nBkYnkbR+/VDva3SZU3EJCFLe016vTud8/YXQKfCC9HNHE
ZjwhjYrq6BVUX7ufxkM26I1XcL9w1nHwKWequRspx/XTNj6T0ztNjdkC11fxWwt+
bAOshXe7kfFNGpg01UJUR/tpGn6Fw6KyM4De5TuldCA/eRnqwXY/9CEqa0YSQSy7
LMcZkZEvEhIvFnjOG20vZxszO/80dg29IFBg+6UH9KnDKtGt9wt7vJ2foeNKoEBt
RkkpdDol7WvqcobRW+EV7lsqgp3P5mV6G+1cn3lAQrbXwryjsfXddPmJzlg5HxMV
64MRpnciKTTjUlGRGEGSt/TS6I0PBlVphHrnqpIfqiYZhBfCtT09AojUsB2IWnMY
cbsFJTrMgAq7+tcNqw8o+gYqepYykesu6sD2oXcgLY6bDG1o5hkVna14mMxgC2Be
A9kKj6AeYgqajipqpubKZkAt+NQHL3xIdm78gJdP2MLAmBrfa+ysKGeUtMZx+l9M
FqFiFP2J/2QWrG2uFC9MtkkRsoPYuwgVwI/uuJL9r9Q+j1y3bgwSat7EafHs6DNG
XphvkjpBZaEjXMj7vPrQYiJtQzrnLeBQnEU28Kvk/8NMwcnD6FCoLJKiFKWLexSH
/y/1kGHtu4uIaxxO10TmkDr3OSUI9/kj/JnqKpygXmPQuPxyhbbRAbRLP+G8PuuO
BoxMBZEQRhsTYm2T2IK//2RgtWwgDxZaaqbh8Pajzi7YqSb8IPBLomZuLvVO6D/O
9J1HAtUgC+yJ+iCJruUwAElmG2WBGacvj+vbEJrcJh8zYDTO7BE7o5Znf2/8jcl4
FSd2dA5cld2MmGvZI6OvdRYPg/zq58B7LUCQK+kNDo6ia/xhRq6qDmGqnEYYLnxp
4jjyBWzbvrTtSACoGdCr5d4wCMIf1iL/i9od7tfxkEzZDGobHSTdxtRAnBZ7j9os
zieQxyOt2Xh2g/7WYjhLkD/zsbYESRaUUInWAgaR61Ht6kJCyh5mtnioab4aj8N1
gZl9UKeiqDmGy5Tj4sCv7rMSFWb7dVnyIJS8VZMXZOzWO0+++R6L3tV9pr3o/Ygj
QZI8YTMFf8UP9jI/Lmjoc3XFoexHBRneGB2iM7XOazBZAhrtKCzauOcItM+zIS+i
r1dno8AcsHD9HQAmf8oU/Ttxn98nhXTyj9Js+1IQIkkG09aG2bQ+R43jvBXiZW7k
a5owu0vY5vVERFl5YaOCPvXRZj+V31lUW2HIwc/Zr58XQmsaLhujp+7vaW9dKuwG
8hcD91VILbKvoESsKQYD+8V3c+KsCM87tE5h6T2my5MaTs8ukdjU6U9H3XWISwb6
qar98WTZlWAiJPZed0rKS9g8gAceKeIg58gtLaK1rSKpZR2N55VeHEd04FDXwvoa
AS7g8FqmMlGrGBtUfkV784amRk35m9GHrZ5PGMF52qZZ3tSF4ERuvGYVb76u+m4L
`protect END_PROTECTED
