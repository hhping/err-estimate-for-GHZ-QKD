`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TthqYGVzMikalwX2xzHBL93cMD/iHOFm1YVcJLEY7WFSpyc40OgmlplpcLP0Nv/u
/90xIGF+Tln2TGg0mzqDvSIS6bq2cbM0+6CxTsIzuiPzuKZScP8Aw6s/ZPKSuGuG
fgbJSkuRU0WmWfUWL7FTTXJ5j64qUWe8/WJ3EKe72pXRHNKGq/1abm/RRq9M6fVo
/D9pG/ofN12+Cpoz9d+UKdWNQEzH/IaGfYJe6P/LccIfD6XdDpSr5gl1x6kswbm9
7uaOPliMlr9C7g29puK25XxHedTLBQx967z+0HulCHv1ZI69ysjGdKIoKIND5ZHg
40q6L0cVOSWfg7jKHJwG12bzTMEKlvDUU7RVBb4IJGThV+cM52aPKsVnLu7G7VWl
HNrOsDwzEIk/vaQpxbvkLNlDwxuiZ0WOyNu2ZeSAZAoDkofJLp6Cl8XixI0WH016
F8MojNciutdzufzmQuv3NSAwPRaJYXV4v2HHPEbq5GfeKih62Lpg2pIBHu9nJPyf
MJYHn5fD0wabq9p2/gRtWuyGb2sgsp2kw9zPIbL2+ntgmjMRiBvXw4Mc7nNszWns
oCU/5xjQabv96DdDiZDSmneuXOdAw45m1QMvaIhrcNATtRrG3vC8Y/T5Kd8eoFyo
AwHM5bcOJgPfn+iSLa6OvoriPml9kK4SFTUC9cDNPCoKt9XVq8zCeb8IrKZUYQo8
vC988Db89ONjeKX8emZ6r/p0Ff9h8Nr00itV4fuw/GUX2jWg1EJ7lPowBYXcmgQ/
l2wknf2mZMjAD0nlhIArRFolJhY9oSEzX3bAZayvR7T13B3oKiTu1livK3uCZmfk
1DKoP/9fVQyoO0oopq+cISfaJX3KnDEHDqh/nbEIWiB3a5tegEupSPJYygoEtyyB
olws93cYw9qkNchfkj0ms6NL56YvM9HODNsVGc4OZ47Bp+KfuEmi9WCr8GaJNucZ
H1bGdYXnv+HWKxYAdYm0bCpE36zQuHexb8Hkj5ekNxGZafodcCkc4WuChl0mX02E
4+kKpRnBLNEF+A14uvKixm9CCEKHB16WvtR5MWdhsiNbcJ5YvPq0oMbr8/0nR+/7
w0CmVK05hZ3yKzDqUIvXRw==
`protect END_PROTECTED
