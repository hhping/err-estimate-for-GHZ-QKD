`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hc7EhkVd29qPKCtCkOVmp6bMY7O0LyGJfAGAuHoVNgXiAoApBrNaqgyWoIhFlsos
JnW9MefQv3fD1faSITgxoC5Ylk3TIc/Q81oDgxdV7cojkzlXtB1M2Tqlg/uZFayB
ZQVaAl/MfeClqQinivtXY8zXcDRNxliKGCeGysoCZluLY5ZvXHg6HoJCS+ZNkcy6
JpI65AJ5eA7wIpDHXXYyDtvyxqkx4+xjSSFeydcC7WhIMVx19RqU7ZvE/45fyAc8
ewCk+YHb5TAakJmb8fFMlnDFsiy5icfALi3HaSvTBO80vaLujjpGgfF5MiYlkWpx
4m+e/KGbPaesUM2RVAuovBPsvsIdyaY2Q8ZJAVaGDqM=
`protect END_PROTECTED
