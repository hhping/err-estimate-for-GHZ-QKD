`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1aVs/lSXMU9Gs8/ogIv1iU13YiMg4knwfnTNrcPPFpqydLk6fpwlber9t7uha+K
bwmJUaTpHAsF+E9sgOMIeDrhicwly0tU3H8LZWuqHLpS33exx4RUYFt0e28LRLJM
JeyNNt2Yq02ntHKme6Q0eseO6NMBwDzND6K3JEoVJfuPdVyGBPl6NDHSnInnCgv/
TEpm0RFBkj+cBHQ0/cwUeWv3XcXrwqaeu66UwX/07Awf661pPTdMcyrAwc9lm/0G
Dv1Kww/UlWtsz6WBlQI07C6tnjTtaEfASY59XP9LTykXqygrix8yRpOKkgsfEmZ2
cIWsZ025INvULrm96JmD8Vh3DiVVW0sc5gXSGuAkJO1K0bXgj4brMtC9rXW/Lm3s
DQM6MwOSkUmzt1cMJI2vb1GGyqaOJCzvDY08KaRzu3K4p6aatKq6rlzAWvzEUqb/
pKBb+jzLwX1a3vE6g5SqSH+Z2XgjWwFnk2FKJpoBjNxuPArm5NMGaNKOHMMzwoRy
OnpvGytFBUMYennGgO3tUK1vYp6ouIs5gtGPIc2ngycyD9jwkQcPvNmlFXz2srW1
YOWLFTIAIm+f/4wRqOZHGCQWZrC8+ieXraaq4FOu7zAVli8MvOQc+NW175Yinuf7
B+gsgHQvPy5ucpIIYM6DqBAmmwDCJOJchjNaRZBOb/Shr1HMLdqCmGgvUXzRDqfG
lOw8IU9rNmslApL2T87kaAlqeyWg1K++zMwLmLpWlsrQtcbZUjyxauIOS3/HWKYi
lgP7wbFqsZND+fMoJQUXkm9MY+UHrl9L990mY7729ZfxREu8NdOgDc5H7J2hYHCp
jqkRR3hSG9KWenAmjrPDPzXSV7HjdK+cjtMkj3zZ3HKATBAdyo58/IPmbtthf1US
vdCKD6uwutTbj/+DinlGQw==
`protect END_PROTECTED
