`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fx6zZsPW9L1C5jXHSgA7NpwuuOXnGVUkKjkh5Sm1F3Pc/yvfLDD+6IHqPPc6GiY/
FdJyIZGym+tb2yT8V4ld8rH2VkCj2ioPgEvK59M2mR2zGQRpCBM9Nx037GFMb3h5
H7wxvOyRK2D1RQpTgegSvnKdsjcZNmwpYsXGfyG6ohxAJmVhxrFal082dMVxW9lT
12EkHaf+3Tcnl/MnkcMcVA2GrTuKxfxIbZqgvxYmyljyejDRvoL06EM5pZqMHT14
0A6blSFZAtSuDQgAkLG/XLaZfNxXHnfX3JMfrNQNeoOPV4/H8tIWunOSMq2S6hnB
DhP1VklxfX+VVTAESJkFwu9ZaustgPNzPi6NZSjQdBjXlTIk5N09AxdLhJ61uXww
0jrRjuNCJ26ebU7/KmaRp8/6Du/810uKktoQ0uQQc/S003VlvUwvP0y9JrDbOcwm
1CWDaK2ZO/ASFJ/ng1z6VkQ8NrS3biP/E75rCyl+qVflirNVV2tp2QJNZQQ2UKdK
YmnJrLvzv+fKW8W0FGgfLtzytCXU7tYgFzMaKGbX9zam++5ydpTlaEoIlAJcAU+t
awT5bovUwrY9px7rpYTBq5cNGqUTpzoKtMm502wNV+3Hz67S56lAD2YBfqqta2BW
+AaQ1obCVTJdyMSs86v+8yVpoHcnUNhCC5GCaUKVkoYhc0D9uqgbjeFHQbbGEv9N
tXwRa04SZ2lz8xkm0vpLXfcO9LVAg+oTEFzZwoEBkVzYbQ6SPNeEYF+T4VhqqFO3
tqR9ElgMDT7g6/0cEaFER4A8SE/tvNBPU5fJx3rnt2Fxavn+Og4+JOHLYqsxOOfz
iODWWmSQ8OOsb4vgE4NQ/OD3bqFiGc0HiosVOiRBML9EDzW5tBPaG950ocVEXwiQ
CrgXiGqUFM8DqJq56QCKXl14oaia2da+BbE4j5qM5ew5LJcC6IStekJKfp/naV/E
RfB3MIL+vszHp+3dOc5dpr2cQlgsMteCjCpInFpXtcS2lM4HwKPM+udtyWTunO0h
NOkT9c3yybOGtT1NZQKeb5dDNLCbKd3TcctGdGEKnRE=
`protect END_PROTECTED
