`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HY9FYCK2qA0TLuD4XF3gbnV8Lbc/ofmNGM6bxx37rUAIK9q2OXVougFcGvJazyO
xsHHuM+8DLHycujzlX0AgAvOfOMSqLnfhmPG6gp0d7w8Wa5DCjdNZiaXzhLViohv
XdSrXjGwBiDGMjfwzAws7/U+9u1jS8KI7y0AP2nW2apzQpHlBXrBayXEoPKxKyKW
t7JZt/5WkZIzzxjlsOthzYAAqN7USSWpuY39tcmGh7+vp48Q4E4A2KQgsUynAW2y
fP/U4+MBhNnXC2m1hIgG9g4Agj/T2JREt3SrO03rGKAj1BcF8eufXuvPY2iEOqHy
vBJprBh7gyHGHL4NqgaG1SkP2cU6dY5bdKZ7lMsrJ6iGdYHLApgYTufAi6QTXtid
VjDMql13Ase8gKiay1noELk9RvyLrpGJDd096YKfmy8deXNsGp4DFXLYEn8xZvcc
V0F68R+SPm65sLb5zLK39c6bH4SQqu3TRTT4GG67OIQLK1Kqfl2vAUE+XIBYXBhz
a+q+uZNzn98EL3z1ixQpWpclCsVhlz1Y1x7Zm2IHsVGzV7l7zVByWDebp3hQUawy
iNcSFiu8uD1QfOFa178x9X3TGSv3JnK8m8iqSuWlKZTHKvvTX7Vn2sDbffVKEFDz
BF6KLGCiORUp291+4LGqrE3VyQDJFu/Qgp7dvYKhhgoDeGUmAV8IJUVGdvUV1BNX
dJ6qHTxTZgYlW+qD9raEwxj48MGzLVEohd73xtCtlb8=
`protect END_PROTECTED
