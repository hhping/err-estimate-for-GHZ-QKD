`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hroV/hJVzFyR+CvwwII7fDrmJMGLMoHsrNwodrdPLX9tsD22t7wyOj7O1YUVaQPE
BfmquVhiznXHue4NZFSzpUwv5maNx9FzYmnPMZv6CCmOZvW439YmjNJcSzbpH9Io
jdY74yLjYY8+ypZ1QKnVdjDZ00/CQNY6Xdly2On44nm24UykmBKzYDtdgNUAxlAX
NEQ/Q1NUTanBnXd05rHyIJIcNckaKSqrs7LR3EaRZL5smXLJHnCw0Z7oo9HGnX49
/TH9+TgIC9J3gNliFIhAalyW4AnBbGSiUhqLt9W9yzAUWPUawwKOKm5Dj+RlofSf
VOO4Op5EFxjz7HpUsOqYI8qvjiSfLT6SisqKMO/Koe88yYcih5GGSmL6a/rqSpnx
u03ZgarAZSku98yxiWfMbzuEzj+zDQdItUJLSyogA+7zU+Nm30o6ugnRYyPKwFgm
eX0qycOMsvu9d/d7Lcaj0LeRk80kF80Qaf2R1kuWFDqI21mWSZiciTmg2vAau01E
VN8ZAZAPswtgS6tzLuq74qhylZz39OaeNi3A7vrCGe8SlAi4lbL0+Pw9rL2Hqbqc
K3Pm/0SSwsiyRVBh70X+fGMHzX78nTWqMLvutWFdJCSl34ix+nJF6tCfPRjpuCUQ
YvEfxpfTEFckKQnfuqt5ou6RFdtXSvz47UaJLsh5fwBIxRfila3uj3noGX6WMfQ4
l4Sel4oRdptAWd59CnYIhbqSj4DotHmtoynf7f0g+EJJFmzgic+hBTC8lPPcvXSG
2LEk2SGj/V4IW/ND+bod1+/E3gHP4SAjCOGC+YOv4x0Ed9clMUbks8c64YWKSMVK
uYwcU+dA4ywHfffdCTvK3odx+q4xei1xFqk3mf0K9+jAREjRHKoLwRWNfqzYiYPW
YKTJ2hUMrs8NSGcZQQsuSbcdi2e7tfWYPOy+5CYH5yg1ebI8ZhvkcrdNPYB7SWCI
gdExOoPtMSN5KeyjLTWCdA==
`protect END_PROTECTED
