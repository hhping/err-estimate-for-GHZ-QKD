`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzlRoXKJy/NFGHHSQf8OG++eA3sBpdHsjDMJOVxypYKLwqwhyB6U9Hg2rW6qrQ4X
fIL4qa8lBV8cS5Q/b6wIcTSx4UbO9o8nGZn2aFvQoLQXYc5LHqcuDWSPQPPd7BOE
dldam5n2dFQq+J+0RaoXX+4ossKK/WKB3L+Q33+A1MSYcgqrWjY3pgrOxCYXKszd
IncLt5F6qYvQqe9DWDy7M71fy3XX9pUy/++Qg7x+aod5QFsbAiiZNpCLfaVW9F79
nfHLXPLsnn9H4+CUMHfVmHY8xs4XBJWF+HYQ1fVHk9AM6H51/FwAL0jI8M3eMZ4c
Wme6qT+z0fJPf/weC7D0XGYKCyMiaOJHYfbpq4ba+I6t9AiPMxgoipukjOb0weIt
ysswM+MrT0ijzd2CCMgXCpQjncqc+azScBHInzdVPPSlaoHPK+Cz6l1y7VHLF2+z
liiVFbXFpur7JUYLxydYzkD0CKEkcTUVLXU9iUBQEbmKkflLDLZIwL9PuemwvWRD
1gJPGeFe0bwVW5EQuxWFpdVM7Gv7wQaF/ikt+P8/gbfTwEBOjh8dvAbN0EOp0yX5
Z3FXei3AMVdXl+B5QqK3PzxUiyihDbrZutDWs9agqQg0f1qGkVhDv8nUjHZD3uDD
WySaNQhp094zcZ2UdWXyjzD0K1m9pX8OHNyn6TTlOsfpX2H23p4hrI/KEx4r4pAE
KqoyySzh7L0bioKIQIzVEN1ZDzZsc1tb50UxE/2jp4VchhBHslUqG7IvRMMVCfac
IJA1LpH4VKJ0fVA9OoWhAZhTUC+IpFy22blm2vRntUOBZLEb1sz8vYpBBskqiOWr
TJP/R5nHizZSBSgR5L9YNFqNcGozp6X0+fnb5tHQYFgwV/8akxUH2WoxPoDK9Wh7
BiX+DI+1PGF2D2LDTQmEMJEIIsx0lcE4CR2W+Zv4RQ/U+tLXPjuA0Gfm6qUEvH87
w3KC20sS+OKLtuOQIW4HVsi6HJZ71db6PkVx5IoWXYiZ9ffrIxntZT6ldNLZHEDP
wnc03w65YFeAV0zUgAH/OMebyilNXTJQzSvt6c57PaQjWQECI+Y0wr3V1SlsiGX/
ZOfZApNc792MsrpwWaYDz/PuxvFSQKqAHiaqG0dJ842XF6yK4AWifDEMaPZfTtsZ
ZiVBLQyx0Ggos1rr7cJMGEO8PZ/4SBH4O85B1Y8oGFP6DJjkBKVG6Bej43vpWlQI
9WV9CRXatLQ3OtLT3mkbLbYeZpAU+CccxuuWM2ep6L+m489jDJRz/gu5vJLCTeMQ
LrPB4+mef/uWgC61ve8kCOsJSb5gi3caWVxXduuhKfyptYBmkr+gqE9xVNmfyxKg
Xc8YYufUG2jOXd4i63GNsgddvaMKx/PCDIP6K6HtToVj0tUvj34636+QAxMNK1BL
Skfi4Wk1GZmV3mmjmtoDmM9XK1RYk/ITWRJhBj4PcyKWFkDVq/YCFcMQ0CJjQkFX
tg1zIg2S2ajN+N7P6Q0Yf6/OOrIY+pXwu+C/s8ga+ozE08ITX6Or/RSgwJAC7llO
Vzl0QMTl9vfqlnmQCJhjiiMjHXiBTK89FF/295Qee87pxYmQoVwEhateTgNr4X//
okVIjHnew3Ft03XDfLBLyjsKRLeBO2jCyXdGaN6LG1CwayZ7ezY1RdzUZhdo7iFl
LMRVJnZA2NWeDHcKCPcbk4gTIVU1/auQ3kFEsfM7f7Q+PiYBJ+yd73g0OtoDGT+E
rdaVHXmuzZjlUoOjH9+3X4Gx+A48R4exouywxx6Htp1tXivH1gvjACW+h40I3xx3
ayW2ky4dwivPv2CovjJ2EnEFulSta+80ndn62QI4NS0EZ06vkhTkjSRv+aLxBzbK
4PZ6b3yA+gLUAUSBJ+HA+CJhWEPop8+93DqPw0uMXPYDe3xzoScFtM6f+2MMwNZC
e90Ktsjs7qOz7lL0qXyXE99U0U6gtOgTxxdqlim7Rp5h8m+ZOReq6VEBm5xOns9W
1S9ASFtWxg1dOYm6fVFR3mrKs1u31AsKP7UGlncUfBFFVUP6gxAyVeZ+Pdp+LUDZ
rfnPxDyJtWXyKkVvjxyY2aoojD9KC4XqWdbt676/vhaKKE3mby1H6KMuFo12wUTY
baFQaU/Yhwrp8W0oY8YVKjq0ak325bf6hXoSxbvGYyJcHxh1Ek8Abwz1xroAVLLC
PbgplY6+4FdM/FcTRumFKDMQDoX+xutsXJqcpViMyJTsXjEPDdMhUd4sGS1mQE8y
VZko9J4HkR3xiwxbKQrXI1NBwRuSPT4nsrXImz3g0KIGFv6b0afk1DWk57/l8LgY
hmk+rdbC8onAgh3XyJA3Vn+Fc+nrRSR4R8mGqBJLV4eziE4iF56zIFVOVKn3DlTW
4ArHsxujPuU7laaEpzbciW+iPMhCabEVznMN7Dh6owfeWvtJJJJVAxEdD/JvH8v3
w11WGSvfFBSR9W9Fvze7zqIWX/fROmTqmlwmHl+1q6GCTTLF1J8bFKJEv2dV0uPI
WSjcZFJUWbFF/VMXX5P8usRDLa234cIsU+2e5MYlI70mWPHaRgw5gwaytPedXPNf
nwhEoOGA/rzItMpEJPuvGOGLNRIftsMLiwKa6RqxcXirCjRiIHGPnpkn+PSRUn1z
VK97Kh93bnB3rxbioQ22vZdkg9X5SngLH1PTd/y6fomYh3EFc5l14zDhxiJXwMGP
cLCi6MNSVJCVc0N0vbfP93R1OkYfDEHCorZgtFDY6hNn1Y7+tszwZHR/hA55+P/t
pXD0EjHHf/CT07E9oGY2pG6t80MMRe5hH2rRkk9+QyEZcX+m5O0iAPPObb/XibKE
6sIoQ+F+kXTjz95l+8X5gClk7dUahdwkrqHUR5HUumwrQ3nI1mPfPrzP3R2xQQjl
YJRr2uCVld1tReP60YSilECR3OEOUTTj/p7fTjvBv1S/ek9JxsJM/RXGdPdTf8xV
a8HXOw1u+3O7FjOARK2UTokW5AzuiNMAsmWjx0mgz1kwGHgTXK/uZMeblO5bcmYX
IPvDTFcl0P6cO0L2HeHBxilMPJmE+WNGIFxSEzc8Vu2fn/462t1JEuxSe/bZzfWb
a6BcmhEN++ybYb7U7x0vLf3C/gUCIX10+1Zsm5JaAy6PkOvq/cNntyqatRQs/LiI
PSFBLyaqEoLFryMk4dFXQgnL3fCPM7glQuYO8lN6+8/xXmKJEMqQY09oZeDinin6
C3H8WnNMnybcqK/c/YDD2M8Jdiz+IQ+1GrkC2wz0smbzTtNocda0ADmk0d68db6E
1eKSmkHGUKZtuBLOpxXpcTo3MSs7/HTlsMApVQIgoAl4N5476LrzNOWW/0PhW20K
jklXFkBgV/lPWnqP0iorirs4MiXZ6yiIa+wG/SalCE9RKVzk4HFWWjBcWEruYXCS
QkqlaCD56bsEt5pZ9n5/6bJ5otAXaqc1cOAxG3dl5OGlHQEyfBkaZArfRXsX01OM
OmUWRFPWgyGgB5LMvnHP1REYSC/YRz/q9ThFIOlRrLRDhLMXweSRTllmgo/CrInd
NQJz9xXSncRmim9Emu4Q+8+v+XsGlFTnIf8U1c3DQ2Xp68vYhxlghZMdY1dodmlM
vjAAI6vH5HinjMbO+9Zgm5R34YItBQh9m4UNkGKg/fK3xWG7O43AdmV3duoYCsc6
dW4bx4s5dtxBgwTEPK0OxSns3FmeLXPfPC/NxZJJB29ml+cKA8AJ74WDra17WzrS
eBSognbO6R8y0EvQ3BvSIyAbuBtsKZGoLpZ6IhEwEiWzeoW7g8j/Vi7G+fwfplpu
lfwjN8dbsQpnQIvqw/0R4KLGOX8Uo5WOSvtSPBvfeHNgubHCNJLXgKq1lggSYzlS
8Klxe0SCKX/k1sfIL/XDtOW7e9C2B+2InoSIR5U3B0iC87uV4ej6nxOpXAmR37Ub
okEPQ1ZLZ0nBaGdy05f9BVcSUyOm5Wc3pSn+rS/3Rtt0DxLvzyPQNdX9pFlTc163
Z9lQhbRHyXVkWoYaLrzXlVyERetm/bXv977k33xL3POdH8Q2wwAHFDcyk/+dksq0
uH9nPzu1VfaA2altdrz3RoY0hjpTym5GalfjgQw+CwBmVOoh2Et5oc49w+7UTEo/
0cxX49jeM8s1okHhDOsWYYaOH7u0xjg0oRxZRWoKHaPyQj3SOuGf5O9XnjxZHsZ4
o6Lhwpm8jX2BHXGjKjWHzD/EQHnsOZYgg0gD4SdzjTDZcpPjtsRkTcj/uCOzckI/
zI9QdkbSEIZ+6lJmbilz+gDRsZCR7XFcHqZmbByrzMqFWJlVjP+DGFkJxR9qw887
CS9ueIxdpfWP98IXSow7qVVhvN96pez0mwy5cOdPwnv207CzQihJKSlAGuTVqBHR
AhJSRYXzcGZiW5IoL4hFEiDe/Vkp26dJxhTDACYUsG/GSTTo3TQWPB8umoiGgLR7
D1h1EGfqkQ9cWgsZAS51rbpEz8GhPKvOlCbDtUiEYfJet5i5X1l7qTU7YAxEKS2+
42MG4TPSnt5spm+MyhYqOLSZl9cbpnPICUYgno+Dt2s04sFiIYizZfI3kQ6dSV4x
XTSQ5xuZcPq/OkVCbBftGNSVHxquEbR03++gN23bqCwNyMUWxVcwuxx2CqEkH6zl
qEaLLSFx6akLYqK7fdctzMnLPiJm3BoSwq9QhRT5x9FniV5UC8doH+lR/YpwzL2s
Pxw7jtMy0M8mR2gY9ddo7tbFRaqa861OoBHiTNqvCWhG1dAYxshdNh28YlBxlwxn
QRSildM+EWXXySRfe5raL5h/ZXqg1o8qIoxQw8FZelPQc/iNCsX8y8p6av1sZe7O
WTMXOE7iSOgjxLYtTkxmK838uoDfqbi9P6XvO6SkfmjkQVxfTBaylncjkVl/stRq
fZXofAzNG+pY3UOgm2z8dOoiieqJYZ5e81oPFZkdu/v1BYwxEDCEU4rwsCzR7BRo
IohVEKrI4LOU67zcYs3KKy9+S7vIVGzkfu2cCbTCv5gOgo1YqF3KnLsP71l52QDV
H4VZjf8WML+6ThnIGNPDhkZyhrspr+oOpWu1fP+M/v3Z7kgFRLEdnwuI7Mo6fnCX
di0Xx7L2wyunY6+uGftpIzRJvhqky7TzYNiqZjvLu1yM+sySSDe1rtV2+kG6GOXY
qmrfGE19GWRkVblKYHZsM5meaSex3FiuVfozlE3wroVX5PhFOZvv1COMp3rHa8p9
QO1SNgOvUK/GuhESlZINB3ej+8R4uUChHOLTQdAJTXQIxQOXWRbyNsBpWkJDEmBZ
t+DTV3fHsfD1dcPcjrvV01OwcDJn90Z3XIj36XEdvdPXfcq3wQ6tBADGCLiuO6T6
GTt30rYh0TiJ7DEEB8DTWrGfyXl6auHPjmd+OMpH7+XQlz9UY1FkgIorrFratysC
FDyambsDTAUVsDSkJI0eoImuzz/pnMPAcRHPf9Dn6uW3nMa7pPVLzZnTp3njbd8e
JDf2db4tEROaLGvFusHnI8i3Wv1zwmD/3TPLEAJ1Tj4m3kkrSKEh5Vtfhoj4jbH3
lno36gQZitkSJFZfw+9+th34GnuRr6FUrhKnXXzspbHNUgdDMXxh5JkdrwoDsq9B
LPtUWlrokx+MVX6mm9lIsKe1/I1iMmpvSKFA4UAwn1RhNHWG7GPPqbQdZyvQPLmV
2Uuk7oSvQr53bFJuhx0m3GlsaAf++xQs8eDTCC9grmCtKI2BEOrfoFF9YEuWjd9x
l1m4tHRqVTJawW+Uevt0Z/itZF0nhphIKlVINSqTzjCxrqtkU+5tEPCZl4hZwrCP
T98SEBLMCJUXBwJwFKKDWqEIRFAKVjLu1L0uRmrRlE89N3/Mmme2nFkyaeyRbcFu
rAVnHA/Nrya56pl0UTeo8zK6+AGgMT7LaDKx5k/ZN0e7YIeEm5jnJ0nvUbqqw5Ru
VZB8oDIM+XWCtQ6phpdflJY0WtszeeJxWx5FAlk5FHmwEPjyFtztfjAlqpCKf+eq
5E6zVEP49dbU2eHWjsgNqQkGcoPw5wkkZV2OtUi4MMMYtVjw6PDbN4MsMjWqRIPc
lkTbTNLBgsSDx468pLTxTd6o3W3un6PxdGt8jHOHSAwoGn8s00nTrPIWtTP1Sd1l
0Md8207Nb3n6HFNx4f07BLNu+bV0bSFOtR7gBwxdUD3R1wij8QF0YqSVabQMWgdl
ZJKc38s3ZVRlfv8aAKqHKPr3T55/B65GrtZlzmoPAHESPs/qfy9R+ivMPcmEIqCF
AwwdHzzsyFDTjXMEuDXJDbUkdkaaSxCtgLwqvFzIefhGPfS8bu2uEzXig8DHQO2Z
OR6xMAJSspW6zoqiXFOmWAiKDVLOndNOOLGyTsed4NftemtydpFEZ+zFYEebzFt8
na5enazbncw528+AYtp/l358f9xerWER2gLzWXZGDfcVyKQRevCfD4e649a1PAZr
5gwKkSOKUZUTi4wAWzgqMXicvMravxIEnJDXjr9tvCqoTmQKYKyxBji5qbAqOaae
I3dLn+OURFVO3x1RmCgOswOFIh3B5Z2LE7S4HT8KE+/fmxSB1DBOp7itopZ26vDw
lMOhxkjQ3pUxXiBWmgVLUSJGDTArG1l0hQwxRC7WF2lJDFKhj7Jy2UhcuiiT0d49
+4Ca2xpQZ1mHNosBh7Dw7vm71hpBVq8ww8lGVc7yUquG+Guz8MecFStCo6t1x9WQ
e3YgBPX+sWZ0mdTAmi0/kAmr0a5jhMQEHyMGUgdh2M1QNh9mb7d4PJh+31zJAiEx
m0JtMrNTrHqyVGn9ReozZcqLh/Hg65GjQFaCDrLirQar6HwXUy40K32TkMiRAvjb
5k8hYp7W+aPb2MgVA1W4mH7h3gWkMWM0grgL79MHQP4BJq5/Waet1Y7q7JcLAG4l
grPUOg8dqrrjokgaqohwnS2avMg7x3+DKzszuUuiAcgbA8yqQO8N81cBfHqiq0i+
JFDPwRP3MiI0gbxKfU68T42t/K+hw3Qr7bv3afrvpwJv0b4o86PI/TWZ0+mDV2db
KDrHDG9lVpP8P0QFOtISZxNE58nG89G/Kbkr3VVgF6q73d17B0goVEKXapUw5yI8
7cXeLk3Qr41BYBY6VPNYmdahqkjwhiY1OHwk0h8QkgXFTSO4tboyNsHGyKEgyG1l
u0ZtGGZ9WYGw0OnR0VSnAchUD5x1cgOVDRC6JuTsV7eTgQULyNgxUsRIsz/fk5Pt
u2ZdN8v1B641BdNqGeiVz/1iH5kNXyew0Ok44ppHQOxkvYzYEb68PKcxt9L9mLxf
Jjtx/OFRTeL5614/p2IKCtflrsm5doOuZjgtxXH1LM2BhoLrP/nnKUAXUPa+2kxv
g1O7yNzySggadaJS7NAI6CCOJik96rEvG//tuQ3sqfMiryoE2OdojCAft3Drylkx
Au7shpBRRainBeJPKD3hsYvmvcBPGf0Ias933fchi+1JzNWumOFXMS3LhasrHtKD
xBvlVv8clufhnwc69FGXCjMIyFo/L3iOF0EZeSZQMmZH/H/WB5K10PSpVIqhzhKR
m4COQODXLs3rI74/S2WDf58fDORKslxJ86dpz7mSXMKqdJK2ltFUDe4yirwx7Vgb
GsbD5mmIa+3jLMPRACJmKDDQVxFt0IQGZ7WP9agxQKFxd06ZRNkiDmVwHaC8J0Ql
zTgVJqXW7j9XdCywsyyOVgpQ37DmugZvMegEZONIL9O0lQhxe9qYj+CZS36wASOO
n1aUWJrtYInMKr54B7OsrTsnlq6rzR60yBXySlfoEp+Nj4tbHUj4Xb2YQPQcMfwJ
O1/BrJ/mOHp5bdzRK0YVxPkc3zKscfqV8q8nbbZnFI0lcakSdfefGWeXMJb+CUDw
N9+OfsvOPGtDvRI12o5eeCYW5NDbxMr3BF8eLMbsTm7tET9T6GqQPRrJQEWWQvv2
kKhsT2IgwyNoDa632aHvwaFu25Ji2k+DZopk0cUiwUt/zFp7ZN0zvMZw8wxTL1KR
lXUXAotDYoytdP149PKBPR1KtQaP4eCNQL8hEGb/ow6VsoVNjLlchLkt2kMFs/bC
a7hvtEvKzqKXAnkoUNt613MKaM/EOEXOWsfnrp/1KNuo27S1vrsqezfa37klNpJE
ndAfPidEQPq0WtVL7hoIqwlGGCBxlcte9jLyJ69gj3nNNZcvCaBJLT6PjcWuyOXz
5DrJAn8IOhu8XHAemrU6gvayqUtSktdZHYxK9CdV16cUl8H+Em8mLrFWAqVmh/c4
JwF+ktVe8ARe7mwp7YphwZUPBf/Dtuct3RzZCxvylBNiNV0p8kGdmGdcCMeT4G4l
80eLEkgOCa4i3PvkNmlPdITmbGmMsDmq1CWnEi0/xVbMT7RiJhUYJxe3ErpjuCJ4
xsA21TnTmO31p+C9FoK1pfjzv8c+Tny9hBvjgrtcVFbl0E2+MPon7itAyOqVtB0B
KSFBPPmbu3reISjMSe/6fcTEcXxPEGCWsRKeuxhQybRJNbDw7spZO7PycJS7/B4+
iNgCc/d/gfmN7dCPPlBROaei0zMgAn2udknlyup9K/44dX4WbbZTKmTdTVJ5PT8F
WRQhbbYiUSk/bG3P+PHy7xfUUe704HUUXD5NTB0eK6czQQ8N/GIL5CCeLK5fAJaU
O0CDSbSbgnh0yeA9FA3g/qDU+ju9su+er697nxl++fk6AD7pomY0EG/gBs2PeTL2
chCHo6LVHjo+xyNnx78QPQtstRALGtqQLbWYTDKjsoPtsd34UDOdzGyi5pAn/Y/x
CO9NtIfnTNOof766ZGrIzuiYJI8toXm0oXgmiDSPixOPnpefcwKhjM7jzIBA7/b7
XwoD4PaDDiC36D3us9ezis5HYAhq3twEDmJ8f02FXy4i1K4a1Mfv8JclsH5PpjJO
n3RMPfp+Q5/4wlC0oHerNe0RxsmEg+DRca41GClThptKULkjR/teppDyzoZh7pv8
u/CpHAWT5rmelDwdz6GdPzU4soXyG4pBb9CeJm5BPwoHCYTZAqbVojWZGtHhaYxA
yB7ftIJ0MJiXsIJE44MDJjIEf0cgovkT85Wdr3rTK2E0K8gIhsAYAwW5csF7ruQ9
RAprLkvZd5moYLnwEENc35q17Yo8/2jwQG7VLZEofcyQVVjMQ/HvpazvM7dcxPwR
aizDFedTTI6pM7UUUNVBxOAH47M9z2V4ymX6RIsE33a6raOIBNxJmecZGmqxOJv1
qxoCMnBpxfdaBXeDenpVpsVSD15PnGaX/NFP3xokFiiz37Ch7gMzbqimUdzjCFzA
IEtOxRQPFkSNWifkP7DpSv+5sArhHa4jQxWeruuOCTgh8jJOY4tkQl+Oo7KTNf3b
TlN2DPVbWE21uNic/iZ4DjZ+w0USMqW6rsaehmL+I0xHaotVY/uGVpf6b0EqSYpK
nfstLWXI3yeprM/SX7CW8fwP8clyjP5F8K/0d52zhrAnkz9G6s6bRRJwNzmZJBkc
lfvI53JYU1027qZWgxS3I8NX6QwKuzeS4AdyzhAfFTqujZIPMXeikaEOEP157MHj
ex7lqTv456vt71anqVqaW8HKV6AZvPYA3ExXKY/TGsYp9GY9GWx+ixy4o5AG5QM/
05oYMflfHI7VitZV8/qFo2BgVpSSt5mwSuftoRmF6vuus7em9kxR1YROvEy1CsVK
Dn6n7u2XNrlYLcmWUj9WdUFja0vKrEfmHe4c/CXlWwWPc0WIiz7+JHA1B/BsA9nx
wct1/5EoTZTMRwYJl/PNz8jlXUNIf9zEY3eRI0cTWLQBN8e7/w6qj/9o0IxPZ2CY
HfLARYbiM7Pk/sOAnwSSSstYHzZ67IAFJhk+SZdvcFL7gVUokMQTedQI4s8Ws+jk
d/vhG0lKtJqJ9Vtjn6MMKEW62XEzrn1rOvjyWro7ELnK6Nng6YWg+Mpxgcjq60qn
ObSQhHsHTTb3XAF5f3Pg9CxSC05qe/6I7mpuuQ11HG9P/UrUstBeT0/cks7oWisH
rCAQD9Vsy7eOlb7CjPyppW7gIODIMdCvOwQoEYtqPD1/2cBVYrmPYOfifnGUY2Vb
Qh0DiWHmL4aqao8PZDweWstBn5WVx9t0P1RPFvLncwSx0770O4InlwnThNCKrgy0
QFzbALGRzqzVdKcrDs6XkMO2vvVji3qx+LYmMyLvjUiuCqHkkWi4kAPNIs1VpaCe
RM9s9xt5En40qlOoZ6WEV/dUia+VSedCL1qqnOvwd/NE96xoLEGhhfG0l6xb86Wj
Dwj3ROqSusDb0HxUJ9kktLPGwfwAnRefazNQwvv5knAHlpGqnhmlqUHo47g1Mwgm
r1KRJwAlTiK6lqBJj6/9yazFuLG7Tf1wr8GyKmnEq/pALbBa/DdPuFsEaqO9VP8n
onhgWDm3sOhAQGYwUkMsbf+OSzdBtkY5TX50+QgGfsj1HpDji2QaxU2KmWTQ41YY
DVibA919kw1iOl6An//lgb0Da9wlhO7rIfeGnBBBqedohv0qIQQufez6YoEPP+Zh
D/MOgjVpk0Ay7mHOqFCpQSmAcAu2OGuRA1FTl7B7Lgj6Bq3Cd50W8BsAhMh0mvMj
MgQNRj7jBfymGk0ftH/hOGuNxitmS/e0957EI3yFQSHMLt61oVSy3OmSw6U3FG/s
zhvOKw8Rhe3U5czS2dgAHroXZ2sYOdgx6Vq8mhx/qnvpVI4JZTJ819dOJW049F2D
tCoSmlOZzE3Or4NEYwFGQiHTlGKOLOoDBRCSrf2FprU7xN8MJGDxQMNxNv0GfjvV
foKP0izqO/I1J1XTbHeGeSp/4AxzzIcQzMcpKr0pMKLYlaxSXexh6CBJTuoqvmvp
Y2vVezIf37aoBCdzUBDcIGGIPpA9330ymYn7EU599Vp0m1mVyGGq4iH/fj8EWg6s
lvPm2jkPQJnhA942mZlD9NkPW3fXPM/UdyFAJ9GW/sswyr6cTlB9+pwAyA47oyjO
MgBozt4eLYsgcEbmEXAWk6OAzWhV4nSXFMmL7BXn9QdR1cTfXdkJEgPreFFVA1to
HDXzCKzhb/BJbIAVnZsRpKvbgv/i2ZTdzjWWQsJndn36PYv+AymB9rdwGU/3ZMBU
Kh5CgVBW9FGwMOZN5pN45SBoovlPoxifAM0kY40o8Wnl1F29ZkQ71vcJi88D9hub
+vC3OzjF6J3uVVuQENa3Zav99WsJR4ZehW1QFaIr1q6LjnFPg6kmo2dyUONUUMOQ
bnmDp4PlWjikxTt52yrjgcR7SEDB4dXJ4GnX7347i9p0azPETrhIZ1uvYKVqJcdG
ih9wBoqMT1WnBOQz5Vt4qN9lcE0EItkci+KvYr9IE9UO1nGq5Ti5iXUIpHelAS+y
JePijDqZCEWnXKxRB7+B2wwHGkvHSuQInG8crehfZVca73/1eRHMR7wxPUeeN1Wm
FcLmh2CEQtxkE4tV33w6Pbon/8AyNSc8NosdhtLuCUNqudhgrwAjKmhHNwKwIuj3
yag9FAg8eewAId5tzosjs4e+gV6YgcsI3Rru4GAdyXf4UGdfVu2/KK5sNI1CN+VR
z80lpYwIXRWkZfjaqB/H2yT7OTWEa6qRB2aY3dQmdbsLhY6iClyEE8HHnLRZJmdQ
ju8ePEaWxSvRnDQ/k/768/40XclOVJDgWfDg2rwvp5Oq24Pddr+dDvrbI8dtd1in
5cH7xSV2Ao/6sjo6HGYgrPthlIug7Z+UuzPfVUXM+J8ErHma7FJQpVWPz9YGOZ4G
RGrur/lrSgKRJ7Neoy5dMFE4Aco28SCMq41/P8jK+KyLByeNkJd7DTtXzmxIJMkC
NvesQzPpuOgRiuDrSmB/cXMFvDUpk4laeyOlyBbzh0Ncxk26HFl8xzRjHNrdbqod
GWGsvk21f0OApeS4PkjgiYHL45hSydJUsJzfnMy7Qr1TgPOGjNQ9I8LOzgXecrNE
1mdlzH51qXrgjmmapHmDqIG2j/SRsCz3ZhxQVql6D0IaEVcHIPB/In6/CIk+41di
7GrJyDcyL0X27mFbTu87iTmXqtW2ZjV4K48mfhl7PS+GCzfqeOKqVT5pd5seRyma
K7Bwz0CMXtMw+H5z/NTgtjqQSFGrEnOG2TUP5SJVuwbJWZCTMzL1EiA9ZCzCdwNT
WSUTxewPdtBdr9ON41fbU8ZAMXxNbK1MLu4tm2Zc0ZSSX9vGJtQvcUglAMFybIDZ
Fbl31EEV/wGHUp90W4/CVl++JIiprXiCHnveZrxELKMgf290tsA2svaMwTTMnoDl
iwy/RWM6BW/i/ZMb9IgXyZ5mJrYmflFNVw7Bnd2yOxDe+Uxtllkb4mEuehm3ooF5
H+IWGzCpm61yr+M1LRncT9pdV/jw+QKjbTl2IZv3AJJ8sM3+CHDWsqxHMfVSJFwx
WBaaTSW7XIBVI5lfzWpTiCUie08XV5xCxEo4T+/zpNTj59nBzVEmxRZxKl4iqNBI
05pfsocFe/CBZTE8qpM8PH7vqGBrFa1VGS67xK89eQms8Z9sLNdPVzGUcJ/q7uXD
56zduQglXIhrFXm4TuTs1GOrcN8pXVsmJHkBBQzAV9f8ihTW2gkN2abI5CEwM6hv
WYeIVOaoxMd67PFDA24J/t3BhQlItHjcMb3RfTK4qH5ByAEVXtikW5wgwuye75oN
w3XL6zq9kr6pnMltzaqoWHkWBvBqbb02cKbpvfZ50zDHAKnZBfoRSmOVAhmbNcOs
JXNaaYi87fSegB8iwbIjpoWz6BiOQXwdczbaFVuDuxxMlUd2Bq67p4ONLtCoqAHy
QZfeyMUpOKDboSPkoa1fcYcPNpqJ6EF63ONHB8XOy91MRauZ+lQuIgMGu7fD9XUr
6VRO5joL+0iWWFvaqh5CToVK1Vq7EMI27jcEB+ACEFtxUZ3xF5NvaXv2a9depNgs
Wdi3muw4C7B+FOESYtCeCBK9IgO/z+69Sadq9FwkAohDhjWAs91KpPUHQqvdAQE0
R6cNiHVe6sdlV5IAVnCRBRQdW1nupcyjgTZTBETbuojL0g3b0oJ+ovaczg2m6t7S
NRqlhGdYIG1BKhkEaknc6L23YXtiruIl9Kvdjl1NsyAR5ySY0Gbsfi2hQRb6rGyy
CcFBUCuRSy4EGQkiAzIncUgzatlQVVzyphbv7JzJDmCZqfxTpQfcnjXn7utUpQAS
ZGjJXCHwl6T6lyI7NqSXysq+mLqD2ffWVRohhr0OXSIRQAavMl43NBrxawVd6o4R
rZY1HpiBv2j1qMtxZAyxThT3JKojl8mkuVkK3THEex0yjg5HuHpJgkwUgkh1c5MG
CDKHhsVkHPswXx0ZB18G3QWSagMrhZGjcTDKZdtkAfYDAXDO6e7DCSzRGxvTy5fu
lBw3XofmvM+oxdxbLmtsjVg7nM2+5QLaVXELO2hH5ObL/qdsJTc6qIFo3lQwcnWP
HvH9v9nWuYYe2M95mYU6mhr2Euu1WDN8cKUxPMrfqtOPAPgfjnfwBJrlIR6QUVjM
GUGHgieEhbPsdtc1BjqigNMc2+DlPNFWNsrH5JwtbiahFo6PCAzEBazDDKKNcPxl
YyTx6qn6QhYmejRNQasKWUtzbRax1NxKM/y56pk8P6+vZVwaSDom8CY0tHVhRtSV
1PFQEFTsZE9gBNpJFXd0fDJ6bIaLsWsptfyuLPfcRRXDxf92beS27v4eC2M3swUL
1UkNnnAVjep4e3AQ75ONjQvAF6ji8MnDVpWT2REEWcpyhMo0RAeOgAundjvkZTeQ
YMYsf2ntBgLyOVXffi/kVPh5v7fUsekT8QQpqmp5qchDP7CLD3G4uAU5QVDItMWS
smSqDPXUqCwKq0gm8LiqG5NK8JJ7HWj/IXoKl6xbfiPNCapZgBD5g/272XNQ5r5i
oV/kK5zvtmyIZn7hyDCBcwoH2MPPEeWTyOsspAKe1MDy/IkiwTZG5ye3hWFnlnot
y0m0IC98TeSTSvVU7uwrjMN1RoTa7TxQS4EJ8y0n6iXHpQtCFb4yu8PLSscvl5B1
EARWNDS7tSUUbByH21KNTs2qDyRamVNgxeEWrl8coOHXYAlya+TbX9EDbqbrk4bR
UaGE9h9fDi8wGW7AtVIDUuElpGHqlWPDKjAdOSrriqlmyMaWci0hvLeUkme6LiO0
xbBxjlBS2qR4wGvU+Jo1LFxWzFrxWdPENFc0tEUgcMkghNxP1BXgwOaroBmgwcyP
LVaKegad9O3piMpgtbpLtiEOyPT3P85IDxpMZHpJifJzDJ3D/lqEuq6PCtOV090t
TLVlYnArrkJ+fgCGFXK9Bsdp0K0tWUUfJAUWQgVlQbKJoKm9jJQdjASuNbPiwxQr
TOxSXGulTWlCpgBcEdbwUH6A3pP4eg5KkQWbY21pKDIVdalWMdf1ORXemojakQf4
brrwQD806km6Qf3WaHJTg+scIRtB9UajelUNFPJ8+7JmdS/Yaxcy0d46IdnQuQEN
oIK5U0KSf/TQde7sb+Vq4cTY+Z8NLXQ80UyR3TapzyncGtWeK+vqu5Rt14dVIgdN
r9v++DXWUgBp14Y4Me/MbqVjs9ift9/IzTARv5B3JEBVRH1hec3rfknNre5VGCMh
SJYvq/IarCmqq5mYaiqg1/A9w07QkuTBiGJ79ML4wSJjfWaD5aHhuUtvevxnmsf1
Igm9lmOLbmMVZK2NIVPJ+RiiQfO6J5yC84M2zQN4vvreXPSsuyezj/kEb/ZyfwOu
QahDePviwlbhk4vZA46nybqukpHuk8IGcRc7tYnF9AiHrq4c9OmplPgKLaIpJv1N
uHEj5VAhp3UAU0Ac7n4Cz6B5WYgR9oR/cORWKuZ8bxXPdzaKEQmgnKnR0SJQtl+n
Fq68/NAwsxqyeaSR2KKAWsjyL9hHFxbJtoSbtpKE5zCeqqInTNY79PImELc+3/4P
D0btaT/GLByto3Hn/vga+eJ+uRHaDOTwQp6zyH9oZMRxu0W6/8PemoxPnrCIr0G5
vI5WgYfbAdzsSmMJhCLh2iyMXg1HPdoTgA6pmJJT6zdYSgWBdLdyiE6MPfqriyPF
/4ClFcDtcm/eG/OHRngsq0uRWJVgT89qrpV/3eNqwBgMpkNXBWzfqruXyyWzdcdK
4RfnTByqwYC2RhDhU05OuUYQ170SxYS8UPFoUN1rLtbr0WVJvgNwEAaJy+Z/qf5y
fn2htN6esGDUttQIjeJP9poiV90NU9aeGsRccVkUiQ4zMz/IG89fDaOqg59PeHdw
Q69fApdbiCOpIe/2LW5vnodK+QeVgK0EY2YFQhzXUWdiYzRr42YlWy5ZzDk4ySw8
aWhEdt0hQqm0hHcOgbP8KRyTkCn25w2yxNbquOGgogoTir+L2MONCgoAI5/jHwjA
cbGTJ9frNu9WtpCEfm7leU7mt/Abht6JAfRB0Iddl06BtQN1wyupirzOKAc3c4Xh
PpSGAZ7dz1C+Jmapaf2LQcWBeduYH5cSZXYvS4WEJdUXnJg7A3zYmcS/bZUF+k0n
koy5QGUETT86nfXJkTFGNNshwlKwN1CXmRN962JlxloYmGD28GRTNmHUTTsNERMN
yvl5AoImwDWmfb6ZgAFsMBydDDWXGne3BubZgkXOt6DbYCXPQeNiBkMeyZJFs8mr
OvlT4kfHxcaCbqqhhvosLFmzk3X4mkpSDFHmPODwxo92ceq6m2xsaMTE/3rRgfhI
6oWtWoLafdCNY57BckcR6B6BgoCWYzLxk/gV2vDoFwYEgOBG2a8+Nq8+mROsv4+M
0fh67TQibKH0vB+llFA4BwxRoIGxRs/TdTmylT5Q9e5iypJK9YVfvsJ9KHrVwibD
37C6MhvHYJFaSbw0gvRH3C840sX7pczin8bbbF4ChLpY8Wr3paFrS4FD7rKWcUhj
BeSNM9K1H/sAzbNCAMf2/48mR6H+vIihakoPnm9OTBDmSNQnUSfDxVs8VLBly/u2
gh4Fw2qhbwrhPwtALeu8I0Hek8nPQGUcqDX3bb9kmV+gQYvqqPO/yP1sWCQVPY8j
FhNkYM+IusNOuPMsotEqXSzjRBDVAdxvKkKhCkq73gcrfEVo42hgpojBhcvCnP3F
J+pROJuxyOs8zORqqAgtC2TlCzFno7ETRdj3vyArGgCUNs0swcTE7e0pqCclMvdl
ihN+vsnhKFVqMJrrQYTyZLPhXucy7O1IqPsDoROhqFFxjvff92R69gqzJOEf6AX9
q+LSRpCRfrdm3Jjqq9gy0dMFTHu9ZnHm3rQfIFQa+cbAwNxUAekDC5t0T5D+IA0i
Gt7WyWC45HNnABnwJmGhfCSwI//ODR/yYHby34SHmO0aw8la1RrPaArZ7kqpnkor
vnVilTdvC01syTE72b5J2oKWDb7vcGAp3RKDTl10mKKfQFzx3I+A9vj3YISUYiul
K13aY0CdhSqJQtriUyQmkxi7/vabipaIWOG1VqUj4dsSJRbglv+etbwyLtFhrOmW
8DhSbM/GwQFYbuS1GAiCn7ZoVOO4Ks1wTLTnwVz5u8AG1E5NDcmim119JkPEKQCM
dZhXdTH3nIkPz9imFG1cYG4yAgOiw/DZjtYibZn6Ulv2iyK47WuQcksZHuMgS3mY
mWNPQ1FBkDYh5A+lO2TITeB7lRu+AmuiKM3RpPLeob92Lxp240j5YaKYSqdXrlJW
+rLkPo8RVhTpm7jGe0ZWhWyT+1gFm5YVnuwSlduYiNFDL0+xmJYHXrVbxwSUQiJL
O1Tn1dmC1a/0ljhocdvxJpEhZsTUOnzkTexplKCVzhCrLoiWJtnL92UGoFATe5jg
JFtjysiEVPhyG0y4Rzitmdj9Ba2o3MHdGZc4Fkr4BttGEILRbxY6US0E1eQ9v1zP
izC/+EwR2anUoXdwIjXpbiuA/IE9XGOnjouQWaaR3c1jAzVoj0ypL7jG/HK0ouVs
5iVvznmZxhIJgqS1jJA3sOtkEWmh1xDiadE2Ozk7/b4caV7nD57mnnQBcSRusHAb
TX3MJaiKPT2VEgDRF26QJqwDptPHFoodTkalAwZSgMm6Xex+Fgxf5xmpNTg3omnL
WNkDvK2KmemdEfZS7AfuV4DPZQOIN4IV/+/5GGffutHLoXPigKOzHRN1BrsHc3R9
c93yVD9cmJSONjIUJefes8K4uljzf1JmODWesIDqCUI0Ue8yeg8GwgPKu2AHz3X4
u5koTFiPK5jjEXe5CfEIvD+dpBVOrMepPmJscZ30yrX+nTZqY+rfceNe0hLgELDm
Bp+FB/L/3NRYXH83gT06M9qtJpU72INNvnrELKKwIYLz4pGvLmMobRL7Yg3us0sf
x4KpFJ+MAoQYyzvn6yks3fDCh9tojfzmKlXzYXPyrA+FuQebYksLYkT3Qgwa/P04
H9X/497doRJf50ivlZWAyNzqTslwjbdydOgxtvo8KJrwFU+4lwXh7qnO+loGu4id
Ap5kZb4YtZ60kfqKVUqhG88D9MakoAhn5bJgDO4kqlm/1B+8X6xUZZ0fzv90j8Mu
Gn1FW0y6AP0+HIOYiZ7tbnY67hKnURayd0M8sQhYhpNmzpQ4PCeoiqlqkx2cNFvh
yEgmhAtjEMwRoOwJCdtiZec9w4LBhKwdiNW0zvoHWWwOynFcwZ8z02eVR3YuLwM2
7S6PplQun0ZNTSftWEnY4jjm2erZMK1Wr/Dt5sJtg6gyCDcR5dV5fOTwvLJT/2mq
yR9zbXFFwZLZHFUJmeml3+CvgyjD1HilDwq7VyyNKczpgNAKuSc0EtK1+8PHKZ6S
TrUBCqP7bZrWZsxeXaKRdP2qH8NETfNUCThtnKCvqs5t0+3gNF8JEZy2/VW6geNs
KZUCHJi9qL4B5yM+ZIQwqSOmgdWFO6+uTMXVLEJcWFJ7Rt0C6HRmuLwbT2MAqYEI
WLYANvxvD7J0HHj4kT2vq6NuBtvwy3dmnGClSjL4a9uwYXssi5RU1ze/nPvKm73q
SbicY+3ZvnM5fzrFiS9Whe1afxF0YYWmm0O7UFTkbGTvRkdmkSlymKj6ktCw4Hiz
qyZMOgKn82XNR+hHlSQ5KHuVNgWCFpBa+FzXHY42PgBIudFb2BiV7xf+4l5V6coB
TGggjcW8eGQnamDJuEirbVXjxbml4phEChyLQyGJjrfFBl2wuJjX+uG/nJs/Gvmg
ue2qUbhlTN4VDUP4b4i0iqg7THyt6CW32M7AXkcezPJ5xBoI0b0OXRrjl4DvZiEG
2MtxDZSJ2NBNxRngrlBiOxs/u/XEKhEU2lSLyw15rvIEjWKDWe0X4/rRax7c3r4m
hUtcc6m25EZet8pP+Mt5LPoVoLNduMHWfwze9+CO6n3DmcmIT+PSmSnulEPYl1Ab
6uHc3wv248MSMOX5O/xvHGb0WC6UkxDetSXqCgoUciKd9twDsVZLoE+X+PN9CE1A
Bl7HA/BVSlX59Rqx001Zw2U5W18VQySce5HrUL9glzfoDhqPbRMjvrCgnae1+oeX
fBhKd7MzNUAuiI8sDrWMtiKA7w6tQHls3I2pDj0eyIY8i36vjQtkO4UzdCTYptvl
xm8gtspGP/E3C4xl8zpEXnEspc/lKjmWeYAuf9IaMOQoTdKXKQGIbUs0Ostaly7l
HiuLO2wFCb3WI/qhD9klVoyJJ1ru4WnB1vyV2S8BtZ8+qwECdK7LjzrkYT/cjRH7
eevVwqJUTXDi+uNIyBtMYQVfnSmYur0F5h2f4U3bkl9m6YED2MphkJSp3bQ/qRW9
FElhqRyQoz+Xc42GIxpcstPDNDrAV1O2TCUH7zxwHGoWFgGSMgZ2NOPHftdutj1h
dw4tBQ7UvEqK20iN0eYu9pxJmbhrrabxi+98dCaETAc46vZs4JxqzmgPdXsL2qMi
wkX1Whyk1HOjvlMDqX8WIf0FW56nRmR9zr/NFEXDYfg3f2ifmr2U9RguduDeqvdH
Zdv2zBupspo6x0ge9o/kSx0nMBCRQmyLSzHeaCLOKDODq/5qGUmNx9HBDDFLCk1J
HgKkbVU0dOlhu1DEEkaKKTZobXaJy1ll3MRceGRtlv0Si/lSQFJvFNzpY+tKZZBM
/6u33YedTDyBVqk/uDp1vVxK40Rq+UV+gjc2GasikJmttVRKuyfcFZB2JS5IKiUx
7qqUT0JT/zzkMLp/Fmrh30JLzyl6S4Eaq7KhYv0+RFxM6bbU2t8Gih+9yfZjtLZz
MnMGLOaWvEZCkkowrqbiSxXh5LqS35OvszH8p6dOu7fWJuab7Wkm/SM55RYaQI+F
d3WJ1zEEHoVExVtce/PufvHcwUDwJUPswDq5vEU/rToQx/cL7Mpa0hy2HWVaFjPM
1PJDqWzrmGN5QVn3NIEvjT6PC6HhCLg1n0cOZ/PQzFCSb/mysxh0X16UaUx+K9Hv
8chNWJLqQubTtrj7+yUaA2Mvs3L00+PZtURZzEaY+6cBb66b0HvZb8nnncGdmz52
XUC2YFu9QS6swS247GvM1C42A8vy28OyZ2K8NDEpaynb2F+k2z0yPSRLZwqK8Gpc
M8HnyRqdY1tNxmqEwYpCxNyeORv8Hz677qVQhh0FuQsmLg5mVbJIVP7wRHHdcj1H
fM05G0WP+0ftgFcVjg70H17TG4tPmc6FqhVGy/sniRyKMEyPyCrEpuR2NlWnEdd9
MuHev9ciLXpSYnvLOLm4JHGZsj6Dl8ETM058FegCzVwPnZ1aRPIUMQqm1Hp7EXpa
f+ZSKywNe6Ex3d1WKBZk+XPsw2ndnR13cbNP8Y2ZBIn/RN9b8zP1iTwymWQZuRpN
FNVj/WgesQUH1t7twItwnbo1t5Yqhel+Jmlyn4/2Ht76rmv106FZ09N+rCI/TN1D
5bbkrOMhgxweU/TekPFGjPHg/B7eTUe11mXLKjMTrwSkdI9ImzhQwd0EATjZCOwE
8Fa3QQEhACIi7FZJHHoDiLIGhfaHfHLgkG8DvFNGvMkqT0Hb2oUnrOTyOwoJf7yR
rMOFQuaoXmD6ZgHKc7JGLQOXWAuryw2iT5FRAJ0u5ClcTe1AuqmrT0Sv0Dr9Sxwz
S653ryh+XSSGASAKPP4ZSRXOr36EXKLGXu+B4KNHK/os/nh0JdoYwYrNcSBtmu5c
zkZv336K4VVFizMCGyfoJw9qNmTeI3704ppLOHUVf4kugIntXQSxA1ZYs1RHwPMm
zYas1uBXXSQVq7ukEzyETaD9C55S3ux6Hne5cCguOEb2JPpgrg4ZsgWbQWcq6qRb
+ZACuuk5ixkDeJ73EOUKr84Z5x+iWONdWuJU2sxk6iT31trYxemvPZcovE+FQADK
g9I5sktJUkQDiL0lBIyJpsV/sNzh0CVvpF/fstEYhuXPWLCwp3y3L4xYbdHaNLyQ
4z/Kg9vrmsIB132LuockUlm3AhGuQcp8b4J0CR3kzUquXj3r6BkgX3QrWxKMnLD2
edqGwVP/Ejp/UThNuZZkKKOq5WEpK3eJMxDM2GmFi4Nso9LJbax6FBvqnJTphDht
Zfvnhb6xCf1HbH+pWWBTqNfGDm9FRdHi68EU7tZbGXNfCojx3t+nz5pEfQnYdKmf
jq8lkkFx3UrKhVhljoHnt4SfR4kF3TxdleqR9rRI2IphlylojuXHhUTXblEQfsZC
KnaedVQluEULrO0DyF69mSZ8ZgrQIwcGxwegfffVNX+PNXbPlfUQYmBKtJLIzxMO
iNIirWNj5y7E4Jf1QrAHPq3F6DurV8kr7x1hV5lzozbXzJK1TRK6SSqlaso4eQNp
jZrTEUXykI+FuocT1D6AXsWu+zjyemCmGRaZuoGN8Doa4cIkbkWP20xctBYwDYQf
HLfOPSIwkh6iX2Epbih2AqfPvl82ENDwlm1lGYun9viApmooIl/2ByVlFriB5Ei3
Ksh3Kq7SArbCv+a+5T/Rs6X1UVvADZx4XYBw2P5qkaYFKzL43fzoeIrNOB/eVMJF
nmyfxErw0PhOACxbAYBVje+FGfbVjBJBECPfgq7rZt3mTKsWi5pV1VRuO9kscmoT
s3tUI9fBM9q5O819B03ibKytHyk/cpyTHJ0Tx7HNo5Q3BGx1wMb6pkN0aJoWkze5
Et+96bJbaSVw4yErHyhyvhoQ1AqYDbEm8SJ29h/JJ3/HVTzW7UuhigcSqpa9nitZ
kyThafpHc/ugrM09vO8E94ZnnmHCBjTcO69lYP6k1Aks/T41R1uRYZaM0JsUUPF1
fGQNcSha4z2taxAaMe81y8c1b3ElXN8riAQc+nPwvOiZo3HMjvUabihq5f5XaaQt
q3mD5LdHIKXkI31F0RotPhOYIO64pbRELf+cEh9B1bytzWc4hHbjLYZrlzbe2Qp2
Q6hiGizS+ZP9J+OeEC/FbOsrsfwgKBWnF5jrJfVNFSbtgfwZa6AVYcIHroCt+QpM
P17xTSEHpNErvw+R2hw6G8H4MbrI/9oFXrtJLEAtTcPeO8baReI8W2gyq1zGYTsX
cpnqUnMuFLx2A6TFZUZPU0mKEL21Kvf5yGC0OLRQUoJL1C6RwOrvwBGRaSmXk1hA
bCwNra6mcbnStHkV6PVCmtifw6ZuncKsp+3Xldsx5W0lWFwMWgjgWYgLVD3KfEck
IHLGk0lT7AJpoVZXgAaSDN9ttz0kHQFu8Fg15Nc8QCwhgZSKQ3NNRSxWqi2UWcw+
sBmVCgGnIkHKWM8aESsrNccyo7oplt1jwMY/B2HvNVOFcx4WieA4hpZW/qpEquLL
kFjFqwfUDCXXYdbah/83uua8XQQF6I1beFsOloL8nWgDpt+2pgAQBsRU+k+2DEZt
5XRkopOqop9CqyHfjifogx8KYUf1EFCPqgCv1u1GhUjQA+VA+ixWnoNKG9LC2o93
/ulXKeObURR7jjLUzoY/RRxC486H+EVUDCgSQJYPLsinOcuBztSAcVHq6Q4rzeNd
7QcTeEkHqRR6DdTlXE3JMF64uTH66+0rgGtqdYHZNFwd6W8HhAajEUKmaNG9pw2s
CszXiaQm0CHVb/qGRfC6pdjATAyzGoLF9K82mdCFa0PjfuD0EiA4h8tn6CXOPvr9
lXfKiIP2ziCB/cTU0GF93/sDTy9eqfgcBoS4ucI1GGRKBOTxA8qn2xjioFzyJJXy
628DNms+E5F9Lxpf9UsRimCrbx9/bt64veNDVR3HLmJ8CCXGHbHGtAVAZ1gfGq31
yzuajGgAp2OGASJFwHneir/5ZXY1IqHJr9Yut1MlTMcsfKVPNb0KqJ4WZOtEEvng
Jgm2CDyKAJCIdp0O9+1bD59r5sdsoEsgOUpu+g1B+3lhGAqc7mniobL1BCdT5ZN0
kaFYEMTY9Jvur4gk8PUa67YtwEfkuF4a5wcOcyGjm97IG/QZ6s9/DnSVt5gETuiq
23Oad+BBrTPKTj7T7S2a8K1NVV1TGhN2Y3KOOELWMCutlkOrTQZmvdWFWtFmabmw
u6HQjTuW+kXp24XBbyuSA7Rrf7sN+6EVFQVTRs8qn5NRxyeHrTX6ZKvIpyXUXODn
NGIAEFIYcWaHIyfLKLeGvXjpuhqg24huwVbNlIDQ35z/9b+MFsv2vtPzxymToHg0
q1b4BZn4+TrOmHxvDshhgfGN9MUBV494AO6G+kYtadK0Q6g+gfShJS/pCs73IOIX
A7FoM6f6+SEossnMUBVrxrcYhMbQJJnW+O9nHu+QVkcYlPS6nQIcqsnNM1waxhAe
GMm/psPd9un8gEPH92xK1dHE15G2Xq2UW4xQWJawHPQzA/vOjGKob4CSrGFxnoPf
MAaSrR8iYsJAn88386I5WwMwdh+pdid1D8wye7XfB1/NLMDAYDGN7cNur2GHsk5Y
h1FMVhWGAc3QXA6DVWlPUEBp4esq3Cb2n3LWUX8cW615r9W4Hp8EYYHelNwEjWHF
0auAiF2pFmgPxYze3Ukpqd2tUrausFvmIs01/Bjvh47/QsaNy27muvE4MnOFY4Gv
DOZH3dPiUZmXitB4gJg44+TXmjkX32wVN3WQLI0naAl9lJD4crhsJ9O7iKmd7WOd
CiUrvCYMkGgE8yy6Z2jONmiYcCUFzvCJA5BmuJElXQSUO2P+h6qAdFbfo0Ptpr2d
EZhytDW3vh3m6eZttexbNtI4+UFyBLqruKEOiiwLLjqXTD+kN8DuIpcHzg46Kk1v
GxuXYLLjjMuX9CbVEoMTWD2EHPNtZQ3ZV8pM1bqLKC9lgHJWhzeVAbPR/ivE1Ws0
oQvSN8Ae1MSTgl4hRbvOighn9bKiIkpNCmXKBgTj+0k=
`protect END_PROTECTED
