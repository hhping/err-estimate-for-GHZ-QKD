`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdsxABv723f+41o/fzW4eCnC0vMrpwKXEubIwjygtWvY2zmGKBUd5Kdxm0DuU5v5
kQIPBBrtxoJAEc+jq8sv0k5aB9BVUWwHtzLha9syFcmj65WD+U7xDEeu9hdyCJfF
Z+7hioNjtYcFb3lqGJOSbm7857W3/bR69K/PTFoGGjs8GgbDJEhigwY+kz/W1lQp
uQEs7V+qnphHiNewPB4fyKYDajSKM6PPani1ft1a2wPuiOmABpmoobxzyJCD1SUN
LW3PJWxe6oJY0IXHOV4sh/IJ2S9k4EvnevJpLJKjTnpcrfrX9bV2r1aiZBRooR/p
qkfVxHAgKjryN3d4jY3UEPgQ9Lj+CrLFVv/6taQgGgHHvxSSGIAKlEE3QT35OciP
x7goV2rW782GWrBotKLd1Ae6BB8TzQzeDCH/7CxMhpKPwNYhJomFkjbBayLh7NMK
ef/3k1nuk3dGJJp2mkP0x755la1rAVGQH5qs7N70dyh8BkWTnQfdP6siC3b2THIb
JVbgeaZFUSIiUFsQFvVbjK6LgXkRp4fHPNr/onE0hME/3aSjdwQzKSwUp6d1X27V
oXySyJy6rrTLzbv7jm0vkFmeLjNEkYJV/WfNMj0PQOA81dsGAob25X/PLHuFQSmX
tAu5ukXDirAE2EAP0JNOETB0c4qD8txMdr4jG9mcJs7k3wGl64/gHeWiaoAR9So0
1MYcQP+EBYN20Y4tGmtCB3N4DsOXL/dUbXr3w1Ivkhk9pquITcRZWq72V2ZQAOD4
umf9mCop2mb+6uI+4Oxq2ZAZEzvoeHkrhQ8UEO89yjsmKOdfABdYO57Xwlda2ZB3
TQhWD4hg6+KUOgl3ph3ugBSXiyt4JgXRHVkhvSxANqymOI4tdgxJTwLMs+Yjk3If
jbjBKCEHvnrLy1ZoYZ4NeZjVhPPeMQzKOGElxI7EiyNTPBskrKVOdj5LKrFJhA5c
V6x0lfZFwVFSbAVB6xmZoo59OReKC2M29F5UuQQOvvJViALD3B1cCB/GsiQXNLYU
SepqDTAI4mBb41VtsWXyJ0iBng8Ao58rlGnHQqIvjok8FHwsk1LjTExMG7q1Sx5N
B7ZwyF5mnTARG2+Ly90Dc9yAbO4cl54zuL/5vl2TSispR3YcuM8za/Zlqr5jIfxl
m8bIf9k575tVk2DI38Hp/vxWvOhq4o+9PRMshwGT2P3VBu/Zq/XHqUnvyzhaD65l
6uR3enbewupmN3uvSpC26M85uA3Ce7gECWv5umdIjwEb8BX6Nd7ZlN6hoGatZO5N
/kCwzm0AfeoZzJFKYik358oMQJint5M4aPYIcdV8pRSgcClyyDe1Q7YwyhJwLfpJ
NCBeZ+qoVL5T2f0Ta5IGBQ==
`protect END_PROTECTED
