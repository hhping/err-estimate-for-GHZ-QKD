`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3gGpCzV0dqxDyZOWRfMiaRydKjhTxBLjcoHZjCAnd9/5K3cIQr5qwxj9uCUJAJWn
4qDW0pKXc0j/ClFCk29jhDpz0IHKR/wvZZAvlQzU7o0+6vwE05+WKTMawNszq+d7
nRpWYvKVp5cRajlCXur8pjwRjtv5t1FVKRIEfwmrFeZDE8WQk65dIvq45742AsDq
PiGUF+cYsAbu7KQlaLIISWWVLDXmz+iuJs2vkfH7k9S0mhWnsN2qW11PkNiBcE0G
NtSSRAVhBPCKaXP0xy4Xsv0aIQ/fp/yacrFQzdLK30sqvdiZg/0Qle8rdp53Ehme
Kz893J4ci73ksXV+6UOWlx3xIj1Q16M2G2lgHGw2F5qVkQfESggf/03US+p6J4rH
sNa41fgjYxfvGSkNUuxDdkanKMjmFwUipIelatySJv77M/8ni6b5f8C05Owe0psL
PUocIgkR6cQuRVFF+Fh4afczcjsyagHAMxfL1otGx2fO8Avd93rkpLeb5a30nl2H
orPYXwF312MiTBpTieCfRM7P34ejnlkQv8pqtiagAjk/Wz+9t8ya0c/dUL4TXUKS
zBQ3C3PahEQb1OGSshdIooKupdT1/jxEoTWrK9NOUt0s+Ribh646u5ZOWxsizF+Z
`protect END_PROTECTED
