`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcnoX3qy1EIZ6yukqZtx12QaJhSetddFCw8hDN9cU3FQYPZr5PVBbc1Nh1P8JpT9
B4mDcDzQBheFFuSuoEZai7snYnqQ8xITl783K4RZhfqGB0gtozXI3uugHeivgvLR
YTdaZywLuZa/UEGtqCyR7kWPrgRJQshBmEox4kHrFh9cj5puZ8J3b1HWm1Zq/trn
HnKxxhyWMrh88ewAHjmq0PiBAA2CoffdCTnjp5bV/VCA7xajVw1i1aV803maMF6y
fNuB09xLoFUR1j3nepREJaG0rQ/emaJyR6BvPvwl2AsPbXW5mzOKTBtVZEI9Wdwz
Qb9wZ3nrEPlD9qHV68tqvJ6ejZxzuBwUOM3AngkgymhMnbZ3GpppocCO2FevVwO5
kTPHAd04FgNEmIY1Qh5ENGDb0rz5ZaXBJuWhYlkICxYO+8tsKbN1tG8xKSOWhauj
bEE7qdyhdq3z0Xt6lzSFKK8m9xjS5kiXD0u+kB33OlXd5MNKNxF79FmFnHDXWLxR
97PrbJMMR5XUA+BVKaD5LIDWZwEWAKfylpyD7YDaFxeosVB/7tDuocKFEurNO/x4
zQd0wdRgj0kCMYjO7QdiqZafmAL8wl9Ynmt03yGcpeeTD1L4FiT5I3JiWsbNzupo
5M1NAryu8AjuYqaGhS1O5eBiTmxT+nwjRwJO9vOtKsA5t9Un35juFMtsFqPZ2ebl
wLW1huDWh0PciljCo16/Pg==
`protect END_PROTECTED
