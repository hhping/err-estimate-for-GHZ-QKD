`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wiTUiBluGePxIfT0APgnVDXgLVQJCSQ+mL0NFEKpdtUy2aU2LdSs6JO0WhLKGSAT
CNWC7dAVQQlg3VErxr1pC0C0ob9lgnDpzqpLdepOGIRN/UNgD2NUVaBGJGf3vNoZ
cr2rBCWjN1KG377C92CptLjfaYL7bswJ11OP/M2jllVqDXcuW8uPukx6U9d58Ebm
Qe4ico7MO7I9SbXeibfpmKZ0pYjlb8i6N+FvNczmbiECr7ETQM6leWKWd2setRhB
zKD04igmd22su/IqZfBI7zAS+jz18U6lbEoTffO3ErVmwu5j4N/rzMRF2Xc9WBOO
gNJ9d6fdT9wEZnLFAPfHsFZbbxUEyYEemmmRZ+vuHJDUBFEhuBqCLyK/8nW5czEE
ou8NNZg+y/kskW9Mot5W9UmglQYQEpcgtqMqR1BqR1JDa3WMFp35ATIGnQvolm/U
93TmyQEVcV7marimKlwQs5WiLRo7F2kA6Gw0++tKCS3IyGi6G2F/OJ6Jd/R75E0f
TWJnLTYY26plbMLxL8gywNoU1lkpUwlFSPqKJQ80z/08XvuX5ws/Ezow/NgAYZDg
O3WRih3OUBaTiqe4iLRFdkeypX5u15+WN816i5hyqVMo94gPS8vTdSyiC2DHuCVN
bjMZOWKNLUdk+yVXqyZTyg==
`protect END_PROTECTED
