`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0NYp9mqEfXkZsuSTyGvz1FxYX5l+cDhJwYptSfn7d9AsQbRM9jCF27e+HtkC0Vc
eg/p4/2sDXc9GM7WEGwbKJZxaNkMuhS91SL8m/9I9f2edhzDXjA07lkW9GkqTf/9
qGS9lGXZ4+cIusz5Tmplr31n4fliywjXXRe6bUDkQjucaDP8lrouksmb5U2+AfhP
N53zcgNr3NBokPrT/B16h9Ig1hyAMbJ8YkQNbqdEu42deN1XrXot/yFVe+eZbnaE
oWgdodtfxo55l0EkNMMvs6VcagHsDBCqvnYnmzCzusVGyI9NT35pfwz9ZK5p8xwk
8hru+hFkWVyysuaAKI/z9DonxsFzx5P2fbcAlatz9yQ+1AvOCsnxtdyd1d/b5Ong
vuGn1AsEb5b+szWDVGilwLk418Qozp0k3IGKioyr+UBbg2dgEkN6KIQWrm201M5B
SORO+UMAKUDLzZLsk6/ev3xgMQ79NZsAL9EIoxQGEuitV2aCYx64poKvY9JRocpi
nG1KkC/7hAwSq4ljUk3sv1zK0SfKhFURC3+Y19leJn9/o+4lVd+Ar3rJOTt8B4On
xHsWFZoGMVB3xkd0JETOq8DfLtphpsAd+LzgVKsZqH+wzDR5WXqBhUo67cso4YjD
IdRZNoSGX6fnZRknnCNxjcIM5sLOEXbrRAwzp7PPd9D385YnCtHELTIojNILoRIQ
yo8pLEa5+OHO2WXc3UtLHwMdKz0Ox0QoLQgFx7Thhes=
`protect END_PROTECTED
