`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Od59Hpl/w4iEWZ6oY232LgDz/BK9Hd8/GGltTvNf62wHs4LCUCQeHvm0d5p1oGKV
huhXNKaOvyWCIkqQIIhKn5O6JFqQ++n//YhOlov5T/G/wcMECkFoE42N/axFc4Ew
Qu41c+VrBZH4TPRnf6L1F46TsHd5p501Rt5Yp+lDHT8qzIMe2yQK1WmjcuxufWHQ
E5bu5hWjFLRMYv/VXDsvlNkwVgAaPsc4gZBYOehKwwqJu8KJgWmEZMgmcPxh+7jm
y4jFlDtix1SmVnujSM0yd+YuHZvpcC4lHKuoXf7AaZ+btlyp/kBsRNepc+BASHOk
dA1NeYOyNbVWTFxBNMBijzsJVm5+YHb1mEIpwZdbUNMLfFWX4pI808rlgBhx6Bc0
l7fnt8JEDvG5FnhjUE+TKWv4jV5jVZH/xEgP46bOGEoixgqf627OiAyRmovhPW3Q
/vguZ3Ctn9BA/oquSSjUpo90CRmemVB2tW4wu1CpYsmVnbVliW05fFk0i6zRt4pN
n61PJwT/qeEn/eVbQHWGJJUXuSPd6hKfWFK31j/FDT95FOV9CwlQi8675h+cYkV3
4ebcRY3UkBjTsDJy/EOYgjKtwSksE3DfcJALJR2qdNq+zLK9nQzptXd+f421W8Ha
XNb5Z4WuNONT30hxapLaH19Cs7TKE3ZPOG80UNs4V8Ge8WCHPUbF2AyOa+RECzv7
Yc5LmiQWu/ockU3DTgJlsmyV9OvCwSlDIDy6gGtrfau9NEKZJHeCNkwiMRHxxk0z
6WGDkMdzTnn579eV0EuTWGjb5ktatcV9LBPZuH+xeOowmNM/Gz1GcI6p/LI/8fN1
0RzWAFIeSBSlGgD2XD8MkWPACvmwpicXhaQKBqRZyjFnLUoEbdxDS/m6vYbJQXfW
14c3ymqzyRJEWaOlrVKTj/P76+zOYVl8ynY1jqBPXD2PUQh0+IWOgJKUOl8q6ca1
Cwh6tT4D5DX7TPu/I4e7Hw==
`protect END_PROTECTED
