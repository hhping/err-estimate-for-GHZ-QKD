`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88g/ff3Kp9HCKFcPEYfSbEG2Mft8Ai63CvUnis1nuN7wNI4PNT5UKF6gqQCgG4jJ
i+5YJpvXHLNoTR9tTh/yYfzlPjNrkNzXKowWSsVXpNNTA30vFH+J5aLaNWAZ/nxI
7qFeay9StdK1c5ql0bTcyyOsqp+Q+KG7FD42KCtUG43mUGv26Fp+EQ+onqPn605O
By49xNJ434ufxjQaZKkkLE1JJUDOo4uOZB55e5I2oDR921fiyj1Sq1i0oM1ew9Hr
TUu2dGaWj6BcnPuqRxqxiTpsCMoU0HcfffJiEhEAKv31xINOqzMflTj3Tq8SQbR4
PBCh9ua/e+C144OfT+qRrDIkfPdJ38bUrVQFtuUtgZWtFEtNMyMrGxdzOsdlGPqz
z59nzlQuCf8JoWv5Pa5PotxXBOnAIu1zJOFFHB/RbQaeOgPh2pb6aN5p4yQHBrV0
J5ahoaTHJ+jE/kpMVIw1nbsC0+2rjomIKUaw1jrWGjkYeedgKwnFJJjoiM6i2Bbt
bIHb5rquR9XbYgiNl3STxAxLsFYOwTyPxqXOEVOR+yBKpwb3XD4YvkbtP9m9b6WU
WDiQb81MkcvJgmCYhBmcHsitMiNieeRkqQj+GJkGDXsGLmvui84EYD5F9fqX7QsJ
iNfSoGPUbRAXilS+FFT3QKyzB52Ssnc9KMbQXvfQLpJMUCmsx5xBAiPsM5pKuq9Q
NK5Gd8nR0VJodRNKvLZUPfsu8uqF06hVpdfUMmOeQnbhNhGtCWlHUt333wS1RWma
RQXoU7y7i1BCsEaEKkahAJxyDeSbsXtB/GcgRKopZ6pyQc/lqiac5Wg45mCEWeoR
nCMj+E7FsNUf5NKnGwY2jym4MvgKXRjH/QSfqRgDbyhzS9V5zr1fV/rcJiDUq5Ob
dVCJcMiDqoyvwEJ/IGjz1hSvU12v3hzH3vo21E1wEEe1jYDIBQgtg+hsCC0OvIoY
juePBUzBVkiiIEFKaO2St6N8gybz6x8rMwCa1OOKi/OmxG1IhoHSB54/bmDXmhhO
c2NrzUMk+bhJaxK+YnYeAsCXVGbudDiXMbKGApUkfJSkcTJZ9VJE06NMw3unUGrD
miVJVv/0R4oKz/3eBQpGVuydf4Z3wuJinF0LQbhoKuayl4ZgswAEApEkdMFwerg7
hU5IN0n+yDzFzi6/UN20RVxYwe+HeESVB80ok5bKF/5dRDZLnkP/qgGD/NTZgPSi
vV9LBbytcHA49NPczMVnFTERMhQ7STo35vF/2Y2f1FJDohXNj7ruCeg9+57HGy6j
5jEH1wF1g9fp4u6Jn6JARWAlT1dIALzJRBqsC8m3urKb5kt09xn7LHufhh65Df98
O7NWqWSeFagI5Ol+WHgY2LZPnioWLdfyXYbhr/HCcKtCLd3Ou/QjZgh+TCjeEk60
zfADOPAMDCA8oOuk0vWYpBFOjz1voOMNZidlfsU4uC0wPVwm8ZCGptXIrMxtcmbM
7wKyWjPshXntTTy+TlO0AcWRWbl7D7cmsq7be4w5HRTg0e9139WXoDcQpzBINGEl
Ll5oOT0Q7hNq7SFtgCmfa4xAFPMEEcZbTlp+CVa6jg3BGFLtyhJT4/tNv8a8EMnF
jde9feh/tMulbfAHIxBfvmYbpa/ELoHZQ0/lYEw6itm8gEAHqhXXOfy/oOR8dBax
cZxbh9S8aV2UJ3LWlvsud81T8FGef+FLuxbRBTB9H6ptykaQap/zXSakCptr5dV6
VmLIpxxAdlgwDrxsK4ZmkJ/jDQFKx+ZBvOQoO5emkOmfv1g6awn6h8KnmJf7eUoo
7y0bMb+dX6qsv/o7+50lGC4NsodfzYRNqB2RSILGvhrdl+zAgjkDtxMBXNo4wzo2
E/qpT8zvuVrT77IaUYJDrpSxtnufh/Wjs0sUlbNgM7YSyVKRbZpSKCnJegsF3HQK
R1xnH8ziOCraK8vb8Ua04Y/T8IgTDg9vq0BAAyiVJg/zonQVXEwonvjpIe2DSm/y
153t5Lmlv8AW4KHuFmaz2JbxQRcDTuQMlnG7jKUCT/7EFKnJIQq3yoqFGmNZrh4W
90zb8GJE6sCNPZZ71UPtnKLr8YS7hxsxFrZD1Ezz6wXWntfae88waOe6cJeFCNEE
q+YaLMZGVZ1Ot+rVUHiSUPtw0DM4/uRbku5ijTkYtKHhpIJ131QbfXKED1LgCRsQ
Y+pLjN6yXztM6mbKKXeQfl1e3XqyaajuBGEgjb7avNCmbevS3EshVp09V6lryOWh
uMbyptBFyCEvsxVO92HRipdPDDdz6IUg87r7u6kVdiX/2pNI77PoSxwbqcKZcgoa
rJqYQ9PJ2l/XVV5oXQQGW6XfUqcv+h88/H6M1ZfjiqHyxFaRCxXNmJG80f1B3fVr
g+Y//4CeU5J6eUpn8dfhIlFjLvcgQgxiZ3j1Dk9arTWXNosjJ7hokCo22iIgRBqR
w2U3ppoQixkZrIlK6gtXu2bb9BtOcnuD9EFcuAMdGHLoIaxMm2c7MnwFtYi1g0Er
JD8fZHEJRGcoJoVoHkTCmqjU0angA3MkLiTj3EIGcAJgaUROjYmUcF0PH0XzvXdf
FUW49t53SSVn41Klg0kykXQ9eEokHP+/TtKExqEmEK4fiC1Wlfz0JaZ8z2nwb2O9
IIWySwEJ9EHZF0oCiRlKy59oiNpq3VIoXsuuPonwThTYzo+bmxDsHNvm5uns1tEa
CQOe2hfW7RGY3Mm3Xlvqsb+W9+C2PvnTb5fIlIxlSPkZiTBvVKXX5rhu9L6wgY9g
lpBpRvl6DRobN3TpBpQHCbd1qR9ybQZgeTAUGRvGJaFFutWc9SLzYxsfZutIXRX+
r05WO53tP8tY7OQiuWfM4n1X0at49Ca3jxjBMC2Bd45iBP889ger4S3Nj9GyEu/n
queq6K2tkr4rESsrJBAk0cnR7Pu+J0Hyl24SIIytTt1AcL0DDY7ATHbvCaPXey96
WXHIOVZqpEXzmJGf4Iuwa8qDalFlhXe58m/8HHMFrpTFxFxgAaVEsxOHut6/jeVA
SEBnGRqMcWnq+OhPO0e+1sBsClqVXKWdBCNSF6To7RLsHYlHxJfSUyJOFMKd6dwx
GkjTjrjCkRKr08PsemiUhOZFcMckvut71R/remMZvy6I0+OG60zTmXtIxCsqdMBE
Rxw8jDmBaCzkeB3QFDEwdCvtAefE2uw9DPqE3VmOv3wiVgF4QMnzV4bywEsY2iW6
51Z9SItIQNF/FkvoV83ZsgiXdSRyuRPh7SxBMVV8EKXCVf0HqhI8Rb+RmNB85Pyb
2kY/9Oh10NYtoE7fetAdG9msu+Bg4GxjDpD5af/wQ6YG603ZqrHID0TmH5UP/vS5
I9Isd/Ft3msPnsUbn6kKkBb64rIRW+UFJpquinq7+DqdGEp0G/37i8p4alp1hssr
OKj0DS6LUaXlof6RFPJseazbWtTGUXZiLxVWGdEJuXJfHS4WtPagey43kZ3az+5M
FF6nkTimOgBIKyF/rOHA/8pIyYaRahpz0EYEeF2ie0UmbYTDJ9oD+aDShvVTQnPJ
MbPVT1ij5looKH1gKsaRuTOXS6arwMzr5JrUiJFEkCr02IquuXdo9HBWZo70q1OB
qz03rn+jBHaTZ5e4lZWJpcmKvYIK9SAeyBsVCgYpis7AZABGJq7FYWDXZM7XL6sz
Et7lR0+jth8X/JkXKOSSDxhWq3eeAuMM8SrGK3zC0lFEWAnjP/hHE2R/vgEEWY+d
hGZwvYpPkklLzaYKfcZjRGNivtnKYHu8Lug3FCoiA6xElfk58hg//t/sqXK/p2xx
Rps+V79XpcCADS9M6q9o22CLCbLJh+RP8Quy9yWtqUnJNJY1iogghGlO6xahMrPg
b/iY6T7mX6x/8w3NfFnibzK49bZ7dDzq0iF4pjI/xWnb5ktvNRThv3VwI0Y9OosZ
A70LkHbJK4zhrhQ3cztOWFKCofStbR83pAcCx5LGdCMhZJNHw3OypihAd4+YEApK
6XS4mqHXVUwiRpISVZ58MKLjPQrXjBGRk3lTkX2+/9s76zf/xfIg8Yvi0eZgJnm5
nMvRyRpI+b76KsyxdkHFLw==
`protect END_PROTECTED
