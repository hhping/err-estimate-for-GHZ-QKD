`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppQenOrvPN0oHKxXgrVC+WwizlTjTl9/fw9W1dT/Ro9hn/iHqXP64CYhs0gpQ2sl
BZSogOab3urMLsthOAi8Ngh0yqB2/diM9QRCxtuDwmoYOkEPjxkB6SlpFl3S0Es7
Kyc5iX6rc1XxSFssMGp55ZTCnRVKn9gsEtbDvgasX8kcBr0fZZuJkm1dhOkEHLNp
FmJlcWz4ZvrmnVFGHWUPvKZ8WaQqpO3R6iWmpGUWATK7Fu4cGdm7TUUPDPBy3HUU
F7vI4nX5bfqwgyb+zddKGsrFDzfAq2fOoD6k8dEIjBJmIUx0UaZElBdJWez8+hA3
tFsxziBLAfW19qCM0L1zdSWPgZY9mjdDpDtYAucVPJU82Hka72aAsrreTF/X567x
R38i/oP/fSvIr50vXovpbiiWpT3ESSVcK5adgVeE4JTOQIDKawVEydxpmX+th+SQ
nQtloBj8QW9ptG5AkkFncp/NrJe9zoCk/1Ev9jQXG84Dch1fnxkFOex1BFzkMWnv
aG6FbwLhR2eSukiMIFrX0t2BYlzJfAKZLeWOVPJOnX9nJobLz/njuyOxmVCd2UY5
QbDbTZEdQsqYYJcMX1mVmCYy5XDj8JC2e0I86IiB3OzpyqEySGvx5c+JaO6tu1I9
a2rS7zFKRxnwci66xVy/BlNFFnFMdKiDRp3A377QkU1Jt/7Rc3rKeyAaeeSnx18x
mtITCxufgDsUlMMdBuNKp+1GBpSk8OjYZxbjI1XsZmLmoJmnQJHvzgBC8PQwjXnv
UnCfZCI72W69rjtVHTsHor6BRU3bgPSXTYhQkrXChwA=
`protect END_PROTECTED
