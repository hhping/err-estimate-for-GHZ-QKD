`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwbCXp9WlXUpQIONqe+6HV4JtMXKOC7jge55RcBQOZhFE5hqpr4V4yjgthlV0P3a
7DvVArFq3ID6iWFYA7jau1SLqvza8r6s55Ga+4j34TH7QsANZYCcHLjJHQZ7wV5M
+AhgdeHtx15aDzbVTe+oTDTsKbdH7AzEJF637PJ9ZNjsFqMfwQsYyFg4Z+7yDT7D
OnFCDe+1wlut6W/ueHuB4Kj9HrFuFyF6pNq1URZ8JwPq8YG6Je4TvPftm3q5uDBh
PvBEADjQmRFUqwdGoxNxpkcPxKLwU2mMELi9z+MFgYKr52DLet0WTcPebLDMY9NR
EeKf9+kynoNym/iRiLEI9xthje5SrdBmdMIT2tUEIm1JHtq4oQ3SYLklRPLG+i+u
W0WMmnSS5SfdDW6eEGZrHaQL7RxSngYrZOikPe/DVigbM9UfgBlOtaNeOS33SGrj
QqNiHYVgsu6HzXhIiZqZnapM8HiNjGSWeAxukGpvphQHipuN4AHbzOFlKauAri47
YLMaPSADleW3pOa8iWdHdl8dT+/I/MmZbDA6lrIC2JS3ODNhCdNsseJBXLZPvazQ
QKD5x+ug1O2tyZYFtJesrRVlooAUA7Z5O/jdyg18xpYZATV2zPS0NhMhC1Q8LCUy
5pkh4DF8s8EkDNRINedA8wU3ldoT6NYfvxmA0ieHPqscUsd+Hyb5nNMvvc9RbOtz
E4JppbGMnevhlezGiHaH+wQrMJmTa2svUXfx7n3COpyIf3VePyUgcwtFRn2yL8R1
CbVvuzffN1FD2jMSR1Sa26X0RZl0YjtBMNErZ/Za44Kt74qRBNBAKK6al4g9ODC6
OqfSNkanVyGDs9hC9FZWqmjySSWrYX0MADXG9cqCk1n50A3CnNVvIqVnDln6Q9U9
1U7h2TlZJUcnJfV4Xx+2kWg5a9+IJYB5C1VyZPrVg+GACPbpU1fLAcPapm03VnDq
2HivM/AYKjZVGi9DqwysBj7sccWzM4mQEvYP71H7cOJGw0dIn0h6MaIGTOBZLyka
Sc4/ln2nrYxbvCaVcC78DeZiZeSHN4iikYs1JlWmywVMqVzUDZLeXoWUUvP1T0eF
PIDc3bl4LBvhboZXGAc9ItI17hc2gxnS25eS9PVeC6VuPPF2SM+u9iovxmn4fgpu
YHyzXT5p80cUDF7AEPRRn8O5yNSDy9wjyl8ReSSKbNgCGpLGXWF1ISsM7rDULRKI
jEFBI99hcMSfDoqJLEFU4xTcoV1R6J+fY3gy/0Znp7wSwYub3IsebRDjTKXLH4mu
6C1yjUt87GZ+hBf8RcV/TMs6W7S/VJMapBvUZqr3f+K5WZKMYDS7gMIFlZGNmmMj
he/kXUw1fBzDA01eexTJvVWsw6ZHVfJ6yhLB3msPSyZZhzUpnkNeYZjFSJeqlwYg
vNT0OZT0kve3VmwYgrKf2A==
`protect END_PROTECTED
