`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WimOT6upgJNwxB2ZjEY7d7AcZFJ3x1fehclx9scxyd9FvMAGVbiuPYqJHdZwJ+Ky
ppajFfcyLJN1qWsRvvxq+CN43uFUt28LkkdB5TQN3IMWrYbw1a8n/NlPHcPLrVck
We5Oku1Ld8E/J7EdJgPFqQS6xiUyXN5p0VubtdczOlqAha9WNHfSvEKdBe3wikY4
4hpAOOO0xGmggyqa/zxMH/qif7qPY7nb5Dqg/IePz6EO4FjsDOuKiqa5vTvGiUL1
Y7m7QbzkWeMWba82jJ7CgJrD1HckMNVgG39j5SYZdUkrvdwImOSStCs5GH0ZJhBt
YJV867oM0EW+WvZoStYXS8B7Uxrco7w+0vsYl0oOGxk4KEYTU7JKtgrZhnn209pJ
BcNN9kTtAx+aTDEnCu38kkHNh3kiW22ndSb74Rxwa4QqUQYAoQXZStfgW2GwAi9E
tTez46ZRIycwKonDYSKByC5xAfL0TL2JT/oD9XZ1a1183WQ7ao/fl+QKr7zN9WJC
jHg0A/FeBgAW8lf7pPc+K3EfITDOHHZ8COKyvi+mZqDPjhopLktcnUhj9P0RD4Mw
ei03SWlcwaSgjVzRPeKJp3kuNV3OE0sgwj9rx1IskjV21OUFhF1uNSsTf3ljvEze
SX8kfbCXb+iKeMsv/WB2Kc3N1tuMI9kx2nnbI7Q2/Uh+LNMSJ1+25a3dlvCS9FhY
kviQHJ4IygqnNuvm8qsLfXUGG5MAr49F1MKMDmv2DjgiIHuEyYI61WhlNjAfDIWi
zzHD+aar1KKGx+LeBbUMI4USO/hyn3dN3HtTuo7tUkv7RlCR+ImkDPRvOJYbkGXC
vVx1KTIYy8JA0oXwizmAQlZ5GcPfhLrsCCLdTygO+cUbDgOvyf3Ih8g7eu1edeoe
72RouCAyzAsh8MTj2AGHgUvF4z/d++/KiSBZTdjDVyDmtEmevyA83vqGaET0l3uH
CFsi4xKNt3WepwmT7/9Pg7KNzHbMRY6zmX3Kny44Pt2B53dCquUxcJo1v5eWwIev
vEMUPYCfC85TJoacaAPEuyLr5Fkk5XH+eUmgIEry2pnoR3YHOWUhB2NAikJ33Xhj
/OkmbRhMFR4Gym6K8TIMAw8MNApeCNRws1wFKA6Fx6gqMM6pFMp3J/w+ySd3RN85
FGwsR72YJOGlds41itt4OrYGNzqAocIaK/E3lhNw3tWKZlD1jNordJHBdQushMpE
LOHKk7cNgDgxNd+v4YCl2Pz+QRrr4NZHqC0PdoEuxe3u/zz2Uwhq8cTN1+tGLL/Y
D7m75361ycXqED6BYbUnC8YIHArqBGza0peFtvWQyLaEQ+VwjycLYk70rqwJqvZ/
we4u4ahW1W6SA3OyqjZxJs5FTpRBZGCG778pv+ii1xbHOvalF7BpMsMY3nqyO4NN
hTPwhjbv+rfB0N+wfjwktCv3EPcZhjdJ0Hrf1N1wOJ8fUq+w0BJajhJIO/qNzE+I
8KUBmM3bDYczHVTrI15o2Ryyv9YhqpJxC5LmYIhvajL/TmpJq1RzteCam3682pr7
wem4JQH/E2tCKCgzBBAwVYdDS3UQpoT8O7aTl5+hhnukrIeCuE/XAHqitO3ZiRN+
9FUZkiHlKw3ioukJx++HgXE1KY5gz26W5+A61oX8MRMyTE5lu1i3UMwz9s/oqmeT
GiseOVa68dY4ngwww32H84Bcx3S/wm6jU5amzZjwwZsFmuoxTKn8A1P4jZouOfS2
jZJkh6PjcxK3Nw2u0e+t+kcMxQ7cbgqACWXFB5ay+HLDu1pDfY6SUVpm+Qz07Ara
oaLVMH961WVeqedprUpgqnsEvTzrWfXrkvud1E+jSAqu6aN6BS6ptTLn9jM1uGrI
RBOsKlBV2V9Z8FeNjNToR6g6qB7nGxVJT379YcAX4rrs0cMVWgpjGtx+gIXGXxhM
6ri42UwO8PaxXCIgMlIPlwPFgDlU8ZJng1Gu/x8KfhWKnXsDnRFFAmQLPIg23ty0
wC711hcVK0qrGAe4YyF+Etkv80m4/waR2aypHZK1XF2kBK6ADVnPOodjmIVEUMXt
j27otEfDcO/VQbL39A2rZ1s8I1dK8A9VQti0nHmcfKcZQwF5wX9eP464LJjH3cQi
yMU49u/00G2aT/i38/LWKDZiZTpXeGpp5IO6E3Is97hVcursotjWvYmMKgRsAznK
RJt09BGVyewoeAIT5jTBuagbWgdUTd17s8mTaKHNFhoELcXPpogmDIC8VGvjYCx4
8bQ41bLZRU79+HeOImFJSDmMDRoJGmBZ53IywwLkaYwW99bDCPAVOx3H7R2PTM9i
OHE0IJeEWfCCIqRSgkguKaaR5ugOKE4FYSnb5m9IJHyvh9AKa4HmmSfxDZrrf9SC
0Ancwa6nslc2VN+vqxMBXCiT4fw1ANsy5AOG0YxD/V9Mfx3RM8NSN3ShiCfJKTp0
ZuPQzwKsQmtBUbibKst0SgMbeKl9EePqFNCuACBXnCEYl97jP+fQplsFRaQj7jjT
w+/jWnmrGiYpZ6vcylLBQK/i5EnAC2DJi8FLYtet7S52YuTELBm7YurQ5tOh1Iwb
I5pPYvox8b62B8rky/M4Ng5h2LC6jH+nlpIMrUc5WuMHtjM2bL+kSyvtXbIuD8qe
634r9s8aTUuwiKtDFqf98H5X/NkrNcUnxsDJqqrdB1cOPiF4BuAbOPoer4vMmwSk
nfLiwutuo13I1Meq9ai4zzWO1CCGmzTYuWwE4X4YJq54nPP2cvE34ZwrMBh7rNJq
74ouYYwNVuK6LBPT2T5NoAsDG5zWnXSKsb7v/r4u9SOEr3IBXQKW9hqErWAkVJ0H
YEFPa4iV6nOkDXg4A8w5f6B8ltcBfiWxzM9ZU7vxFZyqYFyPP3RDnN1jZ3WGuBfW
0cv6g/3YC3gknTbPv+2pF8Qjzwgl1SC0TF/S1Pf7UQwN8ixgMDTvoezXzPrzjEfE
pIQ0XF5eyJlQwvu1odXsd+wyku7BchmfpzG8X8QUFSrT7wQIXfgExN3r1XSRfMSO
UA35auwl2zhbuUAsLtRGlOn/KoS6JjYIAemLStvVC5MLRn65lXzCp/N4At4rRaBb
L0Kq7CQPd4LLyF7kewx0gg3xdDu3qobBh6fSYnkjQekbCSfkAp/9BJ56NR879zuM
JhhOf++CfkPsWfP6GMRLK34ve73is8pTtcXkQoA2yg4g8J3cr8p1T0IROmCaVnt2
rd5+YwSATPyoNUCO196Iphasgo4SGSp+Zk2ocj5/w3BTslEtELKDI40WpuObn/+g
lUCUL/zyoiSkUdnljQMxwkLCKBPKiuJZH+ijPkUZ0l+hLCd0kODq7fzXr1hMsFjC
c0x2HO+4CY2pooAmrPVgdvS36ZwlW0sEsbWQeLbj3gLO4CElkPk+H8DcXb6pDsQ+
zxkTFUfxpJ+5IrTvUdY7O33linskz7SQf8ss3UrusShEhh+A+NQBYFMvn1DGj++1
GTiL7Lrm4s5A1gGIgbUEQo4nzIiLLnIiGje0g4ykSstaaGNNvVap2e2IV8UJMNvx
Em409J11mIH5XZH9uhBophZ+MrlUYeUP8OH95bqKvJnfCA5deC+ZouN4nFp2g148
1Hq7lMS8awAjixohsSU3Ywguzw2DV3IsxCi1DiHTFhDwPclr/2kffR2d3Bd8KUH9
7TFeYSOrqjhj8YFgqUcTGPlR2TaWOV4WqCboNOSr5g1x718d1u/PMugS1s+yIgOF
uAQSDYmBhs30LWb7lgOTqArFLdwWpVbmw5ngLfpMXGX8xcdea4ZfpzKLAbuAVl1k
NFrM8ruyWDLt/8FAiM+p6nyX54wGaRlxxjTvEPF+VUvKv85Mie0i4l7+qgLW7llA
U6Pp/CVR71z3t+b1UrQTVXb7nw3Z9siI4rJak7MJW9aK+nvjTyAAPk95Trb2hqHF
L7gxW7QYWjXQziupWhI4LlNV15Ehvqq/pBOsv3AuqEkEWKU9Lv39qF0d+hzUShLg
ZkkwfNHT9xk1qtiK2Vyq+98ZPq4hvAvchyB4gBOY9XGqUPNZFw6yBtUPSE+VtT+Q
zzMjgldEZ8woN1XSrPf5p2SRRoKmox7w6xZG/VWnlzkrmQ2VQ1Lq6IidAc0SekVL
6hqM3rp9mlNvT/wY0OsPAuU4HbSJ9XIIS5fn2lJkZF4M9495cAyn8x/87iDD9zLk
cyjtaM3K4swMwAGc194S7f+kZ/zas2gRrKz/EEqox7IB/09gZdFwPh6yeUbGIiwD
/EVgoyNdD/2fb7cIhwlgDiSuatnVo69dQsXH9KT5N7c8//fteNImRLzm4JWavEqT
ixq3kQLY1oKffhyV16iFa+crHTiS12/t+k9GoloUofVOZGzSLld1+7uVa+gUxAhX
FJaksb7MGBR1117LqOvIhgvQRZXQMgTZ9kCoqieVapYDRZZsCTTHGpKkmVeGEsT3
SN9ZkNN7PnwTzccy5Lx5c95fwe2iFbFLVOEL49CX7PBqAqsSTISQRvzGuwX5zAjR
IreB/oHGBd+kapPsqy5c0RXq09eI4zMzYKpTAbYvaBNCl7d1UjtHc4uhiQyU2V9w
4EsvPsd1oXzP5tB1na9VtwfVn/0IxfvamWG29qnUvekLZusXkYxguWF5Q7TeMzwG
61AisiDSDPa+YaaMk3axGVxBenWs7XlaiqNcOBDVUKHScltUNsZluJsZJ9Ehazu0
ZGDgq15PXeLdBbVtvW3B5IP6y7ieB0oOd6GaU9M0wTUjCc0MRcxmnBmhOD0p8Std
uc12ADPFN2tPusqGVlxUpxi73l5E96AaBplfFq67izvviT/M6Sol5GCNkShk6+pr
+khntkI4hOoJYXz5vbofcaTTnH65W1bUcy+XipGDAsD+u2NgwGnBgZOFzXhJviGA
AZlqk8jKrcaFh1cqEIJ8z8mN3fdIOu08Yr+rhryfnp8+z/tm0LkncYlfep+9+FJL
LmxQvSbpnvqP7f5yx3AchOBCMn72wI86v9h5+J+A+sGuZNiP4RBf3B2N/WeZQRAE
2XLfPq+6UG7EzNpVWlVTr3tn7q6XoFyYRORIq5SF1J2DS+A/oDcS5CrPw3MuRAAy
hkiXwygZl4LsLh2qqPJTpbF1V+w+qMYpWw2rUnxixLjCAYw6jJjMwvabe2FOnaG9
b5VSagRI7eRqwiUbj2mYGMTOAG6g6yV8/BeSpUPB4xk/TuOsYlN7b/Sn3sTktryx
d4YAAmwUWYYA18q2+hE2e8T+u/OgJZlQbarKvvAfVPfYCr38OMbZREo/flkvAspo
ipKP8E0UNMLvmSCpRvmoV/Tl9GSSe1QF1AOhvEjQ7zj7oUsd5ScDp9zRoDjO2T3s
1vItzWuFbCNJiMzqGK2Ed2k3rGRuKNGmrF6xOFNSYV6yYZi/s+usK+ickZZs51P7
VdC6FqZl9zyTO6HLYlklbvQm/GjeYvMMJvJF2fT2ZrL0GZi3guYbyQQu1377sbFw
AdmVdlP2K2jGW2VNznLPsQ9mMPk/PvYti6pbVJtt3Iy1YSgD/1vIC4KA6dvMQvaK
5Mt5vMvvrTRMQRYbqwxkIXtNhCovuJHUakY3dAAiLesXkMVcKMSDgy356eI3Z7P2
vATOdrr+EH66Iwczqrx1dDQFRDSPDuWzjFPrFG7qUJqWKMAXmaJPsMi50gE9K0E+
omRScodZk5zlUEStkDTyOKrlxEimpSi/s+iEYWAjkF7BhznrNQbVW3ri6YhtBZSd
pKyp9gi/bZF41ZTLV2Y1nkG/04b3hd/fLYct/H0J/c1GNvY5tYi0Y/oSJ1/TC7xy
JwDuRCLeOYGxhNMDAVY+AjvoCP76tE4ez7Pyx08FojUFWHyVRO5QfmiTWpgF17V6
rGtH+wi7pazW+GpqbV6EtidEiTpQhjT/W2BJpMDZMTnpe47KWIAkxikpWUy9qp4O
y9MZyn/6r9LGh0mVzqwsol1Ng7VHimRwQpU98TlhwSna8xvGvwuEsVWxx9Ze2Uv9
Jtx9HjXVBl1nKRPWny5KZRrRTkQxu2F8E0BA3TmMEc8/R73FDVHyHpVmNn5xZd4O
0BEdJpB4d2InqLigRtKCiMcI1207unyD+JhUiqy0iTzVFv/kTXeC7JVTC2USEXCw
wtsw+zPZFIXBuuCZQFhSsQgosEjZCel4ur1PbBDM/+Leh9HfkWleQbN8pabe1wTW
eIXgqY5Uth0ZHJKe+ycj2tCBXeGzBuF4xI5EIcThle4/9/kGNR9QrHIBsU46UAOM
0IgvSpOU82rj+2N7LoqvmXof7wzDBbCXEY5gAZYCgG8pfM1Qs3e6E01+iYPeRSm+
CmgVsI8TpfOUQq3Uj0QJQ6ckqdheW12DZlZDdDXKCP0+vBssE+Fdug6HSBTt+MZG
+JpT4GUA571C1ug0Jtgsm9Mrf8GuLwHJn4u5ogosGofUwI+S8E6d35snarug67h5
kcpr8yop/cA3yMExa6Av9QmavlwNK4gS+ef0dmpWfK/4bEGOSivGDRfNGayYcwXW
0kEsu9IagLxgoFrmdNVAV8CuPluwa9sUylVQS6WcnWTAttc7u/nDXcJTdY8MJsj/
NS6VLDxVknnh7kUES4YMfE4HaRmnNMRVBT5gIES431fg4lc1+g13x5QorWR1tLrH
ouk/tD4+/dSvWDCiZ/HAiAhkKvUC8U1Jm4A4+KiXbENpI8V31b+0ykanQbPEq4Lp
8tHxE/38nfk9Wf12NL/me5pt9Mm0c6yYyzTLv+TCvm32OcTNA0dxZzBEWmDRevSN
+yE9GCFPzVqHTvTxh/jG5SVu/69MkBAMVfVHnd4PlMdg3b/tIoQlV3NreXEoowx9
TaPZ37LDYwtAdo3LMF/oGaChlzwAYDfiSlD5u1R/DHgsDqxpuyzl0C8RC8lyiFmC
8heRE8JwQi3sJYIFUMCptg1wq3qef9ou9So0eAChhz9Dhb3lILgMeZBrqoxKVRH3
gBKPtIAYZJZTVu80Uoqwi7e6KzuPF3hH6SUkcRtcCanJJykNIjrhNSuWcD0bwiCz
X/vI5FH2R3+lKUIxkK8IMFB+KJBkk0Dfirtqkt9RvKoVLn2lCiuouCRYFXBHb2YP
5pR8P1wXySgNSDZEXkUE0e88egmoqTRYVg5wt2qcpSesxItrGJ3x8GdjrbatY1Q6
2VDjOAD+DqfzWMpC/eoeh3VpA7eKgKgfD8u9DJ3OALjL9wgmKrjMetwCymDUI2dw
ts5ifjbDQYXBa+u5fSwY1rReNyYJW6ctG3IziuFw/JbsnKigXItNeI9+o5xWCL6Q
9NZcfyRyLjYCC63U212n1mHbdt/cXRewxMOvuvt+djRlVUiHdfwLVug7iSJI4RJ3
GBSaHimKiDcTtQRWT1QDyFXnvmXJ/yKPTEZwymRlpo0j1c+R68KS+/WSVvMSRJ8r
LZsimPBBNrLuKwLSjvIfeT1vuFPJxg1Hh4jC8VIl4xRC0tCs1vrUWNF7XiFDRCqg
vPc/KI3PlIvJWoe1oW32afrrGUBDowk7w20DYpJAVr9ED5hp8toq7bwKqtLtwS3z
jZ5McQQZp40OuWMX3Fsxbz7F/CYXqB981p6We/DKWvXgFdZFXfqR3a2qX54pI/fR
U7IXjmYppto2eNJGYaDEKt2f71GFoiEv+TQMKx5Bwe7E2x5vO8dc5qVksASysZVT
277e5Tm7tbXCKGpmyCE9lw2pmtwd5QUigtsTI1RVx24gAPKI74etHdRZMXrdhodj
ZBY/aMUH6o180PrOW8YkW0EA5UghefVPsCaRKC3IkX1D5pTCoym6lA0Q9Cj6+x9G
2+wZ7upV6Jczh5pVlrVK5Z1Ge3hByizzdaGPO+1gDeXJYb+GkbbMaDYKDwCsjEhw
lNGGmdf3MCEFJOVokeDaYXcTgJRxIU7L4Ttpg1GM9fSBrF8OYUug/WADRS2KVEgQ
tsUbYK0quSJJNSRGOvE+rvNcAfJXKYfPT453IcW9turNlVdi4PNeCjRsXwYzx7nz
7/QgZo5YYVDNdo7yDk2l1qUExEl3gxfla5SliUtA65VvNLK9w3wUhC9JGSq/4XsW
ANu/BQw/VUf16IlOHnNJ9Kjphshv/FVtakqtNyRFrX6gAYzxtS6lVbK96/79cvRb
4WGf3sc2deR62AIbTael5LAVjHCk/my62jhY6QT5KDmnTwTjJfi9bsri8BnplEkw
1ziYFUjzwo8SS30B6na/IFKJt+rylOPoUJU3TULyqWPLpwAmZGOZXuYQP29/aayv
AwcioQag/j+PJ0icW/PjYmITO1s7s9zITU+IwC2eZk7WKU2+C9SSSxqhIw4u47UQ
+O4onsznQTVCy328/YwDbRVA+m78o6Dr8KVgYdZAcD1Ly9h4XEvNnDNW9HnakZgs
obQsuGvjn3/wk1R+R5b4MVxAUrJR4rcTfMHXCREpmegBAhxUhPPde+tu0x84OJVx
uM+PXxf7WorNgMr5GE4h5ka4hKAHPsGY34R0FZyoaFeIaZ4mDVXwu5VAPcXC31lf
b2uhUXe/acUdEhWFuS5lmHxEv+B8c+tDpJ+LgWdqnbHtooqph4qw9s3FWWRaL1VB
zB1B9zEHY54SMt142Cz1dPgJKs+fwi7igcAfBp+1FfBF7NDW2N6e2L1NFsjNHf3P
w7e4DiZ1O/lU75FT4QxrS4nl8fkJDWxfNCDd5fNacaT1zDJ8xILZRjoNIHZgiT7x
`protect END_PROTECTED
