`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5et4wDeUo1hngkDHl8krv9igtnOA4Bse2ghDSm6FEsik7aLjB7PXymaMmWJ1iWWB
2FFWw+V78S9PeQY1rv352duf59pq7FjrVKSCF3dUXoBsG0yLjidjED1UfozCRJXF
P1G6zWl+7mJo54K+3vJcXOHyrQPMJF3LHeM3MVeK8lCuoqVYOVFUcK2yXxuuXWe1
2FiGqlFOD7R8SXBVjgnO1XJriW0ldX49E3nb2oLnn3KpAkFJEZCy0wUXcsY0PrVX
pNfc59SdWxSER9vrEf4PbC4vbTvFdsNqbK4ZwNj+FYd4MzoAC6k6N/nBkbG5ULFc
QUXVVEykjevRoM0ilT+gHPfZSaN8b2olaaFhB6i0bqzBz/jz37PtJx244kiv49Pd
WVAkEiSsFgzz7HLaNHpZZXO+ERLuBwK70siIT0pd4OoPSQrWn9tPnAhreG9pir6B
cXgOiyVmK1dyTTFVSnx94foBBAseaZrDMzBs7a/SRjcWSOV9L3SW30s4jLmjkjSA
4aakPMUgR9Ac3Gxw+GIPZI7IkfOGjY2p6sOhkFf6UL244sy/sYUJKOzaxCgL5w3m
UqygDe+eJCwPW+BX1z5EnYJZSyzHSijCyst7VzU9/BkpepUVZWRGlgGmjFM/N/Fh
nKrmdxOx6EhKJAT+3ne5Q1mR5dB620WhDVjT9K838RTWJVXVutrvEnQU7xQku84t
kNkP9/aRxVK1fWVYizsCyvrXsIiG5flzZu4b2Q1+stGuUqVsycNGgYJ+Kzz7tt67
uZcfqhOhqsMvR6spx5SxYgwhSxcjhuhCUF7+kIgNjwXW7JPPdHhBMcVCdKw1j0tD
eREFrsoMIGmAyKFo3XVkmT6xHnG0Egg/YDlBaOp69OQ4cKnSrViTT3YVZYcXjfRT
nrs/F8K7nBXd+r8qwIYpkPtM7OF4uYkFW1BQebwW3CRhcapUu8XfKGKC65qSwIMD
8BftX68NFvwB3rrFb1fr3b8ipsEsYhE96EdTVZ8I1nlUJtEHjp+goF2/qALYBx+8
1lpdkcDOpxi/2yy8jmuWjR26ZKOuWKUoZw/UQMxfpyU8JhP5J1mDRQpqdAiNxReD
TzRfixR77NSGWSJjVnxPBM21CTfirydweSM9Mq4ABBiv8ouM5vRf3upFaf4/YWGq
Lbz3t/Fqg/ohsJdaFCQgPtCvBxiKULvamNFYhmXgMoH2JrTkFmX3hUDKGvzeC2Tm
4+SaSxUxfmjhX9a4PGxKD7TI7Ytqs0Q5rBwAI8ixds1jfN3M2EqqowLU+s5tmYLI
rNGsPhpo12WJq+NeBJeD6AHEqMXrbuCS+Y5Pi7X+kzpWkWqtcjml1Y+XdF9Q72mJ
eByXbPDocV/R1M8XcG5XH0D7xmLlECM19Jlwn0MH9+o8yTCD9hM78V0W2OLyPtrm
y6ELqUjT/2cZFpaUSMjNhDPaSUUhdJs5nKGRNsM7cxY4soxmfDqCuBlK/+/8jMga
vWburkKYeuZzOsd0edQNXNxXHw/g4c8tNs8fWab1rlskZLlKEUYA9JwcrtlUzTgX
khOJ9UbbNyPbQdtcdQnt7H4CbBIVlMDE6xotoWS2gqXDkjYF/7pW7ZmlNy5HM3ls
xdVx+Vqn1kQphwXqVEX7yXGPTle5I+BQN8DYy2WSj1lnAczBe+2EFbyzW464OtDj
hRf4QzahS/Xd21W1ibBaDqjnEOG0njqFC3bhPbxWhIk4dQ0UbqkQzmzSzNWQ7/yV
lsB1BJW4hkMhE/sgXg7uI2ro5V0ciPuZfMojT/xZ93AhvIMPUIUq/so/Wwnf8mpR
9rPcGdM/AWIYonfi9U2Z4OFRGtQsk1yxXNe939qyT+otc/BGWkZCh9m1NTNRuERF
DWLiBz9fzCmHI4Jn3Skudn97AJZBI3yd2tQj4Dvv+KKlKVs1SAOhAQdff+bxToAs
0CXMizCZcRV9iz6O68pIG+fcm71qwlUJJveN99o5PTjMNz4v6J0A7PFEhNE+ILVM
`protect END_PROTECTED
