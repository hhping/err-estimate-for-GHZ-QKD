library verilog;
use verilog.vl_types.all;
entity twentynm_tile_ctrl is
    generic(
        silicon_rev     : string  := "20nm5es";
        mode            : string  := "tile_ddr";
        pa_filter_code  : integer := 1600;
        pa_phase_offset_0: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pa_phase_offset_1: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pa_exponent_0   : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        pa_exponent_1   : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        pa_mantissa_0   : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        pa_mantissa_1   : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        pa_sync_control : string  := "no_sync";
        pa_sync_latency : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        pa_track_speed  : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        pa_feedback_mux_sel_0: string  := "fb0_p_clk_0";
        pa_feedback_mux_sel_1: string  := "fb0_p_clk_1";
        pa_feedback_divider_p0: string  := "div_by_1_p0";
        pa_feedback_divider_p1: string  := "div_by_1_p1";
        pa_feedback_divider_c0: string  := "div_by_1_c0";
        pa_feedback_divider_c1: string  := "div_by_1_c1";
        pa_freq_track_speed: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_wdata_driver_sel: string  := "core_w";
        hmc_cfg_prbs_ctrl_sel: string  := "hmc";
        hmc_cfg_mmr_driver_sel: string  := "core_m";
        hmc_cfg_loopback_en: string  := "disable";
        hmc_cfg_cmd_driver_sel: string  := "core_c";
        hmc_cfg_dbg_mode: string  := "function";
        hmc_cfg_dbg_ctrl: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_bist_cmd0_u: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_bist_cmd0_l: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_bist_cmd1_u: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_bist_cmd1_l: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_dbg_out_sel: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_ctrl_mem_type: string  := "ddr3";
        hmc_ctrl_dimm_type: string  := "component";
        hmc_ctrl_ac_pos : string  := "use_0_1_2_lane";
        hmc_ctrl_burst_length: string  := "bl_8_ctrl";
        hmc_dbc0_burst_length: string  := "bl_8_dbc0";
        hmc_dbc1_burst_length: string  := "bl_8_dbc1";
        hmc_dbc2_burst_length: string  := "bl_8_dbc2";
        hmc_dbc3_burst_length: string  := "bl_8_dbc3";
        hmc_addr_order  : string  := "chip_bank_row_col";
        hmc_ctrl_enable_ecc: string  := "disable";
        hmc_dbc0_enable_ecc: string  := "disable";
        hmc_dbc1_enable_ecc: string  := "disable";
        hmc_dbc2_enable_ecc: string  := "disable";
        hmc_dbc3_enable_ecc: string  := "disable";
        hmc_reorder_data: string  := "disable";
        hmc_ctrl_reorder_rdata: string  := "disable";
        hmc_dbc0_reorder_rdata: string  := "disable";
        hmc_dbc1_reorder_rdata: string  := "disable";
        hmc_dbc2_reorder_rdata: string  := "disable";
        hmc_dbc3_reorder_rdata: string  := "disable";
        hmc_reorder_read: string  := "disable";
        hmc_starve_limit: vl_logic_vector(5 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        hmc_enable_dqs_tracking: string  := "enable";
        hmc_ctrl_enable_dm: string  := "enable";
        hmc_dbc0_enable_dm: string  := "enable";
        hmc_dbc1_enable_dm: string  := "enable";
        hmc_dbc2_enable_dm: string  := "enable";
        hmc_dbc3_enable_dm: string  := "enable";
        hmc_ctrl_output_regd: string  := "disable";
        hmc_dbc0_output_regd: string  := "disable";
        hmc_dbc1_output_regd: string  := "disable";
        hmc_dbc2_output_regd: string  := "disable";
        hmc_dbc3_output_regd: string  := "disable";
        hmc_ctrl2dbc_switch0: string  := "local_tile_dbc0";
        hmc_ctrl2dbc_switch1: string  := "local_tile_dbc1";
        hmc_dbc0_ctrl_sel: string  := "upper_mux_dbc0";
        hmc_dbc1_ctrl_sel: string  := "upper_mux_dbc1";
        hmc_dbc2_ctrl_sel: string  := "upper_mux_dbc2";
        hmc_dbc3_ctrl_sel: string  := "upper_mux_dbc3";
        hmc_dbc2ctrl_sel: string  := "dbc0_to_local";
        hmc_dbc0_pipe_lat: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        hmc_dbc1_pipe_lat: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        hmc_dbc2_pipe_lat: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        hmc_dbc3_pipe_lat: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        hmc_ctrl_cmd_rate: string  := "half_rate";
        hmc_dbc0_cmd_rate: string  := "half_rate_dbc0";
        hmc_dbc1_cmd_rate: string  := "half_rate_dbc1";
        hmc_dbc2_cmd_rate: string  := "half_rate_dbc2";
        hmc_dbc3_cmd_rate: string  := "half_rate_dbc3";
        hmc_ctrl_in_protocol: string  := "ast_in";
        hmc_dbc0_in_protocol: string  := "ast_dbc0";
        hmc_dbc1_in_protocol: string  := "ast_dbc1";
        hmc_dbc2_in_protocol: string  := "ast_dbc2";
        hmc_dbc3_in_protocol: string  := "ast_dbc3";
        hmc_ctrl_dualport_en: string  := "disable";
        hmc_dbc0_dualport_en: string  := "disable";
        hmc_dbc1_dualport_en: string  := "disable";
        hmc_dbc2_dualport_en: string  := "disable";
        hmc_dbc3_dualport_en: string  := "disable";
        hmc_arbiter_type: string  := "twot";
        hmc_open_page_en: string  := "disable";
        hmc_geardn_en   : string  := "disable";
        hmc_rld3_multibank_mode: string  := "singlebank";
        hmc_tile_id     : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_pinpong_mode: string  := "pingpong_off";
        hmc_ctrl_slot_rotate_en: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc0_slot_rotate_en: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc1_slot_rotate_en: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc2_slot_rotate_en: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc3_slot_rotate_en: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_ctrl_slot_offset: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc0_slot_offset: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc1_slot_offset: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc2_slot_offset: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_dbc3_slot_offset: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        hmc_col_cmd_slot: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        hmc_row_cmd_slot: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        hmc_ctrl_rc_en  : string  := "disable";
        hmc_dbc0_rc_en  : string  := "disable";
        hmc_dbc1_rc_en  : string  := "disable";
        hmc_dbc2_rc_en  : string  := "disable";
        hmc_dbc3_rc_en  : string  := "disable";
        hmc_cs_chip     : vl_logic_vector(15 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        hmc_clkgating_en: string  := "disable";
        hmc_rb_reserved_entry: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wb_reserved_entry: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_cfg_3ds_en  : string  := "disable";
        hmc_ck_inv      : string  := "disable";
        hmc_addr_mplx_en: string  := "disable";
        hmc_tcl         : vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        hmc_power_saving_exit_cycles: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        hmc_mem_clk_disable_entry_cycles: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        hmc_write_odt_chip: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_read_odt_chip: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_odt_on   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_odt_on   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_odt_period: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_odt_period: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rld3_refresh_seq0: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rld3_refresh_seq1: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rld3_refresh_seq2: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rld3_refresh_seq3: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_srf_zqcal_disable: string  := "disable";
        hmc_mps_zqcal_disable: string  := "disable";
        hmc_mps_dqstrk_disable: string  := "disable";
        hmc_sb_cg_disable: string  := "disable";
        hmc_user_rfsh_en: string  := "disable";
        hmc_srf_autoexit_en: string  := "disable";
        hmc_srf_entry_exit_block: string  := "presrfenter";
        hmc_sb_ddr4_mr3 : vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_sb_ddr4_mr4 : vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_short_dqstrk_ctrl_en: string  := "disable";
        hmc_period_dqstrk_ctrl_en: string  := "disable";
        hmc_period_dqstrk_interval: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_dqstrk_to_valid_last: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_dqstrk_to_valid: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rfsh_warn_threshold: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_act_to_rdwr : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_act_to_pch  : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_act_to_act  : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_act_to_act_diff_bank: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_act_to_act_diff_bg: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_to_rd    : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_to_rd_diff_chip: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_to_rd_diff_bg: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_to_wr    : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_to_wr_diff_chip: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_to_wr_diff_bg: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_to_pch   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_rd_ap_to_valid: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_to_wr    : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_to_wr_diff_chip: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_to_wr_diff_bg: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_to_rd    : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_to_rd_diff_chip: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_to_rd_diff_bg: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_to_pch   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_wr_ap_to_valid: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_pch_to_valid: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_pch_all_to_valid: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_arf_to_valid: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_pdn_to_valid: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_srf_to_valid: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_srf_to_zq_cal: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_arf_period  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_pdn_period  : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_zqcl_to_valid: vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_zqcs_to_valid: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_mrs_to_valid: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        hmc_mps_to_valid: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_mrr_to_valid: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        hmc_mpr_to_valid: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_mps_exit_cs_to_cke: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        hmc_mps_exit_cke_to_cs: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        hmc_rld3_multibank_ref_delay: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        hmc_mmr_cmd_to_valid: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_4_act_to_act: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_16_act_to_act: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_mem_if_coladdr_width: string  := "col_width_12";
        hmc_mem_if_rowaddr_width: string  := "row_width_16";
        hmc_mem_if_bankaddr_width: string  := "bank_width_3";
        hmc_mem_if_bgaddr_width: string  := "bg_width_0";
        hmc_local_if_cs_width: string  := "cs_width_2";
        physeq_tile_id  : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        physeq_bc_id_ena: string  := "bc_disable";
        physeq_avl_ena  : string  := "avl_disable";
        physeq_hmc_or_core: string  := "core";
        physeq_trk_mgr_mrnk_mode: string  := "one_rank";
        physeq_trk_mgr_read_monitor_ena: string  := "disable";
        physeq_hmc_id   : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        physeq_reset_auto_release: string  := "auto";
        physeq_rwlat_mode: string  := "csr_vlu";
        physeq_afi_rlat_vlu: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        physeq_afi_wlat_vlu: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_second_clk_src: string  := "clk1";
        physeq_seq_feature: vl_logic_vector(20 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_sb_ddr4_mr5 : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hmc_ddr4_mps_addr_mirror: vl_logic_vector(0 downto 0) := (others => Hi0);
        hps_ctrl_en     : string  := "false";
        ioaux_info      : string  := "";
        ioaux_info_valid: string  := "false";
        ioaux_param_table: string  := "";
        rewired         : string  := "false"
    );
    port(
        pa_core_in      : in     vl_logic_vector(11 downto 0);
        pa_core_clk_in  : in     vl_logic_vector(1 downto 0);
        pa_fbclk_in     : in     vl_logic;
        pa_sync_data_bot_in: in     vl_logic;
        pa_sync_data_top_in: in     vl_logic;
        pa_sync_clk_bot_in: in     vl_logic;
        pa_sync_clk_top_in: in     vl_logic;
        pa_reset_n      : in     vl_logic;
        pll_vco_in      : in     vl_logic_vector(7 downto 0);
        phy_clk_in      : in     vl_logic_vector(1 downto 0);
        dll_clk_in      : in     vl_logic;
        dqs_in_x4_a_0   : in     vl_logic_vector(0 downto 0);
        dqs_in_x4_a_1   : in     vl_logic_vector(0 downto 0);
        dqs_in_x4_a_2   : in     vl_logic_vector(0 downto 0);
        dqs_in_x4_a_3   : in     vl_logic_vector(0 downto 0);
        dqs_in_x4_b_0   : in     vl_logic_vector(0 downto 0);
        dqs_in_x4_b_1   : in     vl_logic_vector(0 downto 0);
        dqs_in_x4_b_2   : in     vl_logic_vector(0 downto 0);
        dqs_in_x4_b_3   : in     vl_logic_vector(0 downto 0);
        dqs_in_x8_0     : in     vl_logic_vector(1 downto 0);
        dqs_in_x8_1     : in     vl_logic_vector(1 downto 0);
        dqs_in_x8_2     : in     vl_logic_vector(1 downto 0);
        dqs_in_x8_3     : in     vl_logic_vector(1 downto 0);
        dqs_in_x18_0    : in     vl_logic_vector(1 downto 0);
        dqs_in_x18_1    : in     vl_logic_vector(1 downto 0);
        dqs_in_x36      : in     vl_logic_vector(1 downto 0);
        ctl2dbc_in_up   : in     vl_logic_vector(50 downto 0);
        ctl2dbc_in_down : in     vl_logic_vector(50 downto 0);
        dbc2ctl0        : in     vl_logic_vector(22 downto 0);
        dbc2ctl1        : in     vl_logic_vector(22 downto 0);
        dbc2ctl2        : in     vl_logic_vector(22 downto 0);
        dbc2ctl3        : in     vl_logic_vector(22 downto 0);
        dbc2core_wr_data_rdy0: in     vl_logic;
        dbc2core_wr_data_rdy1: in     vl_logic;
        dbc2core_wr_data_rdy2: in     vl_logic;
        dbc2core_wr_data_rdy3: in     vl_logic;
        ping_pong_in    : in     vl_logic_vector(47 downto 0);
        core2ctl_avl0   : in     vl_logic_vector(59 downto 0);
        core2ctl_avl1   : in     vl_logic_vector(59 downto 0);
        core2ctl_avl_rd_data_ready: in     vl_logic;
        core2ctl_sideband: in     vl_logic_vector(41 downto 0);
        mmr_in          : in     vl_logic_vector(50 downto 0);
        cal_avl_in      : in     vl_logic_vector(54 downto 0);
        cal_avl_rdata_in: in     vl_logic_vector(31 downto 0);
        afi_core2ctl    : in     vl_logic_vector(16 downto 0);
        afi_lane0_to_ctl: in     vl_logic_vector(15 downto 0);
        afi_lane1_to_ctl: in     vl_logic_vector(15 downto 0);
        afi_lane2_to_ctl: in     vl_logic_vector(15 downto 0);
        afi_lane3_to_ctl: in     vl_logic_vector(15 downto 0);
        pll_locked_in   : in     vl_logic;
        global_reset_n  : in     vl_logic;
        rdata_en_full_core: in     vl_logic_vector(3 downto 0);
        mrnk_read_core  : in     vl_logic_vector(15 downto 0);
        pa_core_clk_out : out    vl_logic_vector(1 downto 0);
        pa_locked       : out    vl_logic_vector(1 downto 0);
        pa_sync_data_bot_out: out    vl_logic;
        pa_sync_data_top_out: out    vl_logic;
        pa_sync_clk_top_out: out    vl_logic;
        pa_sync_clk_bot_out: out    vl_logic;
        dll_clk_out0    : out    vl_logic;
        dll_clk_out1    : out    vl_logic;
        dll_clk_out2    : out    vl_logic;
        dll_clk_out3    : out    vl_logic;
        phy_clk_out0    : out    vl_logic_vector(9 downto 0);
        phy_clk_out1    : out    vl_logic_vector(9 downto 0);
        phy_clk_out2    : out    vl_logic_vector(9 downto 0);
        phy_clk_out3    : out    vl_logic_vector(9 downto 0);
        dqs_out_x4_a_lane0: out    vl_logic_vector(0 downto 0);
        dqs_out_x4_b_lane0: out    vl_logic_vector(0 downto 0);
        dqs_out_x4_a_lane1: out    vl_logic_vector(0 downto 0);
        dqs_out_x4_b_lane1: out    vl_logic_vector(0 downto 0);
        dqs_out_x4_a_lane2: out    vl_logic_vector(0 downto 0);
        dqs_out_x4_b_lane2: out    vl_logic_vector(0 downto 0);
        dqs_out_x4_a_lane3: out    vl_logic_vector(0 downto 0);
        dqs_out_x4_b_lane3: out    vl_logic_vector(0 downto 0);
        dqs_out_x8_lane0: out    vl_logic_vector(1 downto 0);
        dqs_out_x18_lane0: out    vl_logic_vector(1 downto 0);
        dqs_out_x36_lane0: out    vl_logic_vector(1 downto 0);
        dqs_out_x8_lane1: out    vl_logic_vector(1 downto 0);
        dqs_out_x18_lane1: out    vl_logic_vector(1 downto 0);
        dqs_out_x36_lane1: out    vl_logic_vector(1 downto 0);
        dqs_out_x8_lane2: out    vl_logic_vector(1 downto 0);
        dqs_out_x18_lane2: out    vl_logic_vector(1 downto 0);
        dqs_out_x36_lane2: out    vl_logic_vector(1 downto 0);
        dqs_out_x8_lane3: out    vl_logic_vector(1 downto 0);
        dqs_out_x18_lane3: out    vl_logic_vector(1 downto 0);
        dqs_out_x36_lane3: out    vl_logic_vector(1 downto 0);
        ctl2dbc0        : out    vl_logic_vector(50 downto 0);
        ctl2dbc1        : out    vl_logic_vector(50 downto 0);
        cfg_dbc0        : out    vl_logic_vector(16 downto 0);
        cfg_dbc1        : out    vl_logic_vector(16 downto 0);
        cfg_dbc2        : out    vl_logic_vector(16 downto 0);
        cfg_dbc3        : out    vl_logic_vector(16 downto 0);
        ping_pong_out   : out    vl_logic_vector(47 downto 0);
        ctl2core_avl_rdata_id: out    vl_logic_vector(12 downto 0);
        ctl2core_avl_cmd_ready: out    vl_logic;
        ctl2core_sideband: out    vl_logic_vector(13 downto 0);
        mmr_out         : out    vl_logic_vector(33 downto 0);
        cal_avl_out     : out    vl_logic_vector(54 downto 0);
        cal_avl_rdata_out: out    vl_logic_vector(31 downto 0);
        afi_ctl2core    : out    vl_logic_vector(25 downto 0);
        afi_cmd_bus     : out    vl_logic_vector(383 downto 0);
        seq2core_reset_n: out    vl_logic;
        ctl_mem_clk_disable: out    vl_logic_vector(1 downto 0);
        phy_fbclk_out   : out    vl_logic;
        test_dbg_in     : in     vl_logic_vector(47 downto 0);
        test_dbg_out    : out    vl_logic_vector(47 downto 0);
        pa_dprio_clk    : in     vl_logic;
        pa_dprio_read   : in     vl_logic;
        pa_dprio_reg_addr: in     vl_logic_vector(8 downto 0);
        pa_dprio_rst_n  : in     vl_logic;
        pa_dprio_write  : in     vl_logic;
        pa_dprio_writedata: in     vl_logic_vector(7 downto 0);
        pa_dprio_block_select: out    vl_logic;
        pa_dprio_readdata: out    vl_logic_vector(7 downto 0);
        dft_scan_clk    : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of mode : constant is 1;
    attribute mti_svvh_generic_type of pa_filter_code : constant is 1;
    attribute mti_svvh_generic_type of pa_phase_offset_0 : constant is 2;
    attribute mti_svvh_generic_type of pa_phase_offset_1 : constant is 2;
    attribute mti_svvh_generic_type of pa_exponent_0 : constant is 2;
    attribute mti_svvh_generic_type of pa_exponent_1 : constant is 2;
    attribute mti_svvh_generic_type of pa_mantissa_0 : constant is 2;
    attribute mti_svvh_generic_type of pa_mantissa_1 : constant is 2;
    attribute mti_svvh_generic_type of pa_sync_control : constant is 1;
    attribute mti_svvh_generic_type of pa_sync_latency : constant is 2;
    attribute mti_svvh_generic_type of pa_track_speed : constant is 2;
    attribute mti_svvh_generic_type of pa_feedback_mux_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of pa_feedback_mux_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of pa_feedback_divider_p0 : constant is 1;
    attribute mti_svvh_generic_type of pa_feedback_divider_p1 : constant is 1;
    attribute mti_svvh_generic_type of pa_feedback_divider_c0 : constant is 1;
    attribute mti_svvh_generic_type of pa_feedback_divider_c1 : constant is 1;
    attribute mti_svvh_generic_type of pa_freq_track_speed : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_wdata_driver_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_cfg_prbs_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_cfg_mmr_driver_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_cfg_loopback_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_cfg_cmd_driver_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_cfg_dbg_mode : constant is 1;
    attribute mti_svvh_generic_type of hmc_cfg_dbg_ctrl : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_bist_cmd0_u : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_bist_cmd0_l : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_bist_cmd1_u : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_bist_cmd1_l : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_dbg_out_sel : constant is 2;
    attribute mti_svvh_generic_type of hmc_ctrl_mem_type : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_dimm_type : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_ac_pos : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_burst_length : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_burst_length : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_burst_length : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_burst_length : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_burst_length : constant is 1;
    attribute mti_svvh_generic_type of hmc_addr_order : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of hmc_reorder_data : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_reorder_rdata : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_reorder_rdata : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_reorder_rdata : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_reorder_rdata : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_reorder_rdata : constant is 1;
    attribute mti_svvh_generic_type of hmc_reorder_read : constant is 1;
    attribute mti_svvh_generic_type of hmc_starve_limit : constant is 2;
    attribute mti_svvh_generic_type of hmc_enable_dqs_tracking : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_enable_dm : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_enable_dm : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_enable_dm : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_enable_dm : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_enable_dm : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_output_regd : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_output_regd : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_output_regd : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_output_regd : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_output_regd : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl2dbc_switch0 : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl2dbc_switch1 : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_pipe_lat : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc1_pipe_lat : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc2_pipe_lat : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc3_pipe_lat : constant is 2;
    attribute mti_svvh_generic_type of hmc_ctrl_cmd_rate : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_cmd_rate : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_cmd_rate : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_cmd_rate : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_cmd_rate : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_in_protocol : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_in_protocol : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_in_protocol : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_in_protocol : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_in_protocol : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_dualport_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_dualport_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_dualport_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_dualport_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_dualport_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_arbiter_type : constant is 1;
    attribute mti_svvh_generic_type of hmc_open_page_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_geardn_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_rld3_multibank_mode : constant is 1;
    attribute mti_svvh_generic_type of hmc_tile_id : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_pinpong_mode : constant is 1;
    attribute mti_svvh_generic_type of hmc_ctrl_slot_rotate_en : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc0_slot_rotate_en : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc1_slot_rotate_en : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc2_slot_rotate_en : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc3_slot_rotate_en : constant is 2;
    attribute mti_svvh_generic_type of hmc_ctrl_slot_offset : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc0_slot_offset : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc1_slot_offset : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc2_slot_offset : constant is 2;
    attribute mti_svvh_generic_type of hmc_dbc3_slot_offset : constant is 2;
    attribute mti_svvh_generic_type of hmc_col_cmd_slot : constant is 2;
    attribute mti_svvh_generic_type of hmc_row_cmd_slot : constant is 2;
    attribute mti_svvh_generic_type of hmc_ctrl_rc_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc0_rc_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc1_rc_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc2_rc_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_dbc3_rc_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_cs_chip : constant is 2;
    attribute mti_svvh_generic_type of hmc_clkgating_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_rb_reserved_entry : constant is 2;
    attribute mti_svvh_generic_type of hmc_wb_reserved_entry : constant is 2;
    attribute mti_svvh_generic_type of hmc_cfg_3ds_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_ck_inv : constant is 1;
    attribute mti_svvh_generic_type of hmc_addr_mplx_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_tcl : constant is 2;
    attribute mti_svvh_generic_type of hmc_power_saving_exit_cycles : constant is 2;
    attribute mti_svvh_generic_type of hmc_mem_clk_disable_entry_cycles : constant is 2;
    attribute mti_svvh_generic_type of hmc_write_odt_chip : constant is 2;
    attribute mti_svvh_generic_type of hmc_read_odt_chip : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_odt_on : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_odt_on : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_odt_period : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_odt_period : constant is 2;
    attribute mti_svvh_generic_type of hmc_rld3_refresh_seq0 : constant is 2;
    attribute mti_svvh_generic_type of hmc_rld3_refresh_seq1 : constant is 2;
    attribute mti_svvh_generic_type of hmc_rld3_refresh_seq2 : constant is 2;
    attribute mti_svvh_generic_type of hmc_rld3_refresh_seq3 : constant is 2;
    attribute mti_svvh_generic_type of hmc_srf_zqcal_disable : constant is 1;
    attribute mti_svvh_generic_type of hmc_mps_zqcal_disable : constant is 1;
    attribute mti_svvh_generic_type of hmc_mps_dqstrk_disable : constant is 1;
    attribute mti_svvh_generic_type of hmc_sb_cg_disable : constant is 1;
    attribute mti_svvh_generic_type of hmc_user_rfsh_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_srf_autoexit_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_srf_entry_exit_block : constant is 1;
    attribute mti_svvh_generic_type of hmc_sb_ddr4_mr3 : constant is 2;
    attribute mti_svvh_generic_type of hmc_sb_ddr4_mr4 : constant is 2;
    attribute mti_svvh_generic_type of hmc_short_dqstrk_ctrl_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_period_dqstrk_ctrl_en : constant is 1;
    attribute mti_svvh_generic_type of hmc_period_dqstrk_interval : constant is 2;
    attribute mti_svvh_generic_type of hmc_dqstrk_to_valid_last : constant is 2;
    attribute mti_svvh_generic_type of hmc_dqstrk_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_rfsh_warn_threshold : constant is 2;
    attribute mti_svvh_generic_type of hmc_act_to_rdwr : constant is 2;
    attribute mti_svvh_generic_type of hmc_act_to_pch : constant is 2;
    attribute mti_svvh_generic_type of hmc_act_to_act : constant is 2;
    attribute mti_svvh_generic_type of hmc_act_to_act_diff_bank : constant is 2;
    attribute mti_svvh_generic_type of hmc_act_to_act_diff_bg : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_to_rd : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_to_rd_diff_chip : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_to_rd_diff_bg : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_to_wr : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_to_wr_diff_chip : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_to_wr_diff_bg : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_to_pch : constant is 2;
    attribute mti_svvh_generic_type of hmc_rd_ap_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_to_wr : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_to_wr_diff_chip : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_to_wr_diff_bg : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_to_rd : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_to_rd_diff_chip : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_to_rd_diff_bg : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_to_pch : constant is 2;
    attribute mti_svvh_generic_type of hmc_wr_ap_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_pch_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_pch_all_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_arf_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_pdn_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_srf_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_srf_to_zq_cal : constant is 2;
    attribute mti_svvh_generic_type of hmc_arf_period : constant is 2;
    attribute mti_svvh_generic_type of hmc_pdn_period : constant is 2;
    attribute mti_svvh_generic_type of hmc_zqcl_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_zqcs_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_mrs_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_mps_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_mrr_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_mpr_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_mps_exit_cs_to_cke : constant is 2;
    attribute mti_svvh_generic_type of hmc_mps_exit_cke_to_cs : constant is 2;
    attribute mti_svvh_generic_type of hmc_rld3_multibank_ref_delay : constant is 2;
    attribute mti_svvh_generic_type of hmc_mmr_cmd_to_valid : constant is 2;
    attribute mti_svvh_generic_type of hmc_4_act_to_act : constant is 2;
    attribute mti_svvh_generic_type of hmc_16_act_to_act : constant is 2;
    attribute mti_svvh_generic_type of hmc_mem_if_coladdr_width : constant is 1;
    attribute mti_svvh_generic_type of hmc_mem_if_rowaddr_width : constant is 1;
    attribute mti_svvh_generic_type of hmc_mem_if_bankaddr_width : constant is 1;
    attribute mti_svvh_generic_type of hmc_mem_if_bgaddr_width : constant is 1;
    attribute mti_svvh_generic_type of hmc_local_if_cs_width : constant is 1;
    attribute mti_svvh_generic_type of physeq_tile_id : constant is 2;
    attribute mti_svvh_generic_type of physeq_bc_id_ena : constant is 1;
    attribute mti_svvh_generic_type of physeq_avl_ena : constant is 1;
    attribute mti_svvh_generic_type of physeq_hmc_or_core : constant is 1;
    attribute mti_svvh_generic_type of physeq_trk_mgr_mrnk_mode : constant is 1;
    attribute mti_svvh_generic_type of physeq_trk_mgr_read_monitor_ena : constant is 1;
    attribute mti_svvh_generic_type of physeq_hmc_id : constant is 2;
    attribute mti_svvh_generic_type of physeq_reset_auto_release : constant is 1;
    attribute mti_svvh_generic_type of physeq_rwlat_mode : constant is 1;
    attribute mti_svvh_generic_type of physeq_afi_rlat_vlu : constant is 2;
    attribute mti_svvh_generic_type of physeq_afi_wlat_vlu : constant is 2;
    attribute mti_svvh_generic_type of hmc_second_clk_src : constant is 1;
    attribute mti_svvh_generic_type of physeq_seq_feature : constant is 2;
    attribute mti_svvh_generic_type of hmc_sb_ddr4_mr5 : constant is 2;
    attribute mti_svvh_generic_type of hmc_ddr4_mps_addr_mirror : constant is 2;
    attribute mti_svvh_generic_type of hps_ctrl_en : constant is 1;
    attribute mti_svvh_generic_type of ioaux_info : constant is 1;
    attribute mti_svvh_generic_type of ioaux_info_valid : constant is 1;
    attribute mti_svvh_generic_type of ioaux_param_table : constant is 1;
    attribute mti_svvh_generic_type of rewired : constant is 1;
end twentynm_tile_ctrl;
