`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82Sv/w88Emh1XvKUL8hBJQSIc8gzlywfpMXapSTEyY04zw7vH3mgMVF0iyyIcUlK
LMZ06H/FMZ5euM7E6OrGxx9N9RzvlgYd+L7OeO3YBt2GLFh+4jvKv6lw8519ivZp
iiciaUE3kwQfz34D+dU7fnhiDTydjjCi/QWCyENDxlj/qA941sJE8TwmfQJdxzU8
d+gae8qNA6DNgSMeW5YzxlcD7yY9r/3WM43jZzfkhvdY0v9WIzZMsSFNIK6jPNzJ
wCjJ6OlIUq4m92DhS2ol/0yjaf94fEBevmvfobRb/iBnu1eOYAerWruxHC569UwP
ONosKpv7vQ+EEoL+3bsHGSwMOq041PbVkdaK0XbryxE8xo6SXkRdauw6jUmH9VUU
0AvGBjz1RmnmQc2R7AZaqiRWBv9Ln9DtsIRDdLY3nR7k0TWv/Mh2u/rb4q2yTbpi
rDk60wqjbZWDzTbeKhPpyOm2rJf1nj19Sg/Xyhv9gASWkfK10oXg4JmchcTrEG8X
RUo8ofV3nfnGXfShl5s3hOCTFyHlxwGmQez5ThM+UL1qvM2yHNFJ3d0mldt9DSsL
9LBenpK78x3K4dqmMKj2AGfYlnRieLoel376YPTodTUDlF5tzSJ59IxhknSh9FvG
WxGUOGk5s0xrp/PZ2Ta+TJRSVtEa1FPGQ2gYjuMfR5usHaIw+zsaJVhEG2w1AiHA
YPRDr4RV8e2pgD19AakVS95+Ejc4rAWto55F6FIPPEHgsiDJ5I9yIPhFFdmLU9/x
qv6m2Cn7ewSXmlEd7yfsxiKp78q3xYXlrNN8MQoCjhWGxX4OvwhsQK/xhuCRK6GE
K5Y+NlQL/rpEYkgQ3ECU8ohDXSdyEE1EdWnIHtMluqvGCKaGh8bn7yr9luZMAzNL
7xrJQd80Vw8lpGW1PaBOV/LApHeIvZYcGuFFEAKLBS7KuCzkor72UAM2O6OWChts
x03V0nzkIITum3IYj1IuIk5JhH5DXTTGkzFySL5MaMC/2JbkQ5o7KKV2XMhIg+YP
z7KLT9rW3suarbI8525ZXxACoxMkHkJ1PJZ3iSzLlRMBveJJPSZCtwmypCBWpURG
MWojXAST1Y0WzqtS4w7ClHfsB5pTdwFHFqrlhrTwD5p6tnN8Bx7+dW0aWk43so0i
e72/AUeLSG1B+0xTYzNEpyFn+brxPZqpvoErO1bpNQUAFHCbAkor2IHZgxDxMtxS
taA7VRv60n6+1J7OTEa06r3Al6vpuNoaNgOwwjx90htWeeUA6koKQTnSoxz/vADT
gVVSs67ZuwsXQPT5qgMlFAFkcEX2tLEOll0s6oCOwWKrvwA0wlpKyN8Z7MsgVWUt
Xef8zwIk/cOCrq6cg7Kk3gePXudp+B/nFF+hpKMVE0tRTmACCBkoIl4adkna4ula
G4PBscnMIhwylPxmk9w7sQAJ3JqpD6uAFoOqJWmraz4TY4B99mOJj2qjeNYhl4p/
2o4SuYe0+POglqdTYkfqAgP8MJv/EgpOvkEy74ok1E8k0iaGvp1kOJUpOH5z6jha
oDddzkVUatlRcuTt0AIyJZPSshKVjdSsrpxJEvvpGPfo71hN7WOMRHUFT21sPJBi
rZFuslZPI4XTlcHt5frMMLgGPnpDdwsOnKkj4rpu7qaZI/+8fMUm88nc08aip2SQ
cMjBMYdgBc6LnvfAByCWQKLxaoaUziFjqtr6fm4hYTLOLvRU8fmqWfrLxm9p7rjU
YSc/+rKmW+dTpnGM1gTrnjuKDwADqp+xlYzjOLa88Nchj3Z/3QxF9WOmxvzybAM/
/ppzrro8WwN2MJhyANiJR3zNZ4NuT3NoqB6edw18Qb9CAKIHVEPa51bq5uegYAdw
h6ht4Gq34JXgfr6BrFs4Cr0kLfZ57RBvfdyDm97dw+AdwDjXFqlvP45BBu0wXw5F
ozsRPcDV60bY7IU+zjChBCKmQKpUt3lmmTBTiOGCdKzuuBRtSOLcDf41tSNm9dSQ
cKZSaaRe++fiRI9Eg6Fql4ssbe46exhpvOLaQMAhSPVuEA2W7GjCpe1eftDGbnF9
3ll4HKu7JfNFeQVq523342yb06OT4UD6M8BYE4u515xt1ou+gMXJniISPRIZaeM8
b18dbVbjOMpv1uqWZ0aNp/p2lb2EBkq02UKz+eBVKscMQtA3zW6mlJtyq704UGz+
38tFuazUfxrLzHj8NzjUw/uA4sjNlqHjIZeJgxKE5PZfuvcFViCRnjFleqDelkpA
k871j0400yJTYHoR5R0whjK4IS7Pcvmps3GHyagY7QbY9yESlATPrAaKaxVyZoKa
+MWnIV+nWwIOy3sP1HPvAJZ4wP10ndVeaYjNnMXERoixH+YftCmnmNtBLYrYSROS
L4Kg+aMwPB9U+MI69dmIWWOMC9DbEcYF52JjAUo8LXTvVYaBod5XTCp4rj+ea9He
GkiY6gMzfAtCJvMbmnInMeA1mx2CAs64O9Hn86/VvIKneDtc59gBA8ylgRO/id13
r+nzAMhNPAdXXRMVFYcdfdF5AELVdRR65AwT81F7r4PcE+RGfAkVinswSysv2bzk
nG20OJhDWqVGPOr2dK8rZDSMEt6HVhcDKJpyjkglhufcM3ePl+mLwkSull9mTJHB
oSAeRN1PZ5ON93hWPFYfvO10BA+qh8Ofxz2fWbKihj6+iOlIyqtBh/BG3Bp+dWVi
Hq4OCKzf8xFB6zJvN94fjAlKfhyMBNiqt6SR5rci2J0zKm2Uf7X9w2a2zoFclSUt
WwFnSFCC9feM/Zh4lxx6KHIaOM3NkRMrrMYeXAT78RGq2NCSSGTy/CndbBYkg35l
Vya4YqygLYNTGDN3kpQZ7btHiu+AaqfK6kPHpVmmKJrvq606z3YLWtNUf4y5j9Ft
+xgHcufXYCmwVJCdRkrDjKYa6SgC8yY1hVlYQppzl3Q+Lm8+H5kPSxHW+7n4NGRL
p3sRK8W3jVM+p7IPEN/QrbGDQ30tCBtR81zL2pp8yPLZbk/lAi8q+WCXUUJeB8cL
`protect END_PROTECTED
