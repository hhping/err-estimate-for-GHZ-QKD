`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
076gFnDdt6VAOviqcVZqLhueO1A77MPFy4g5UfR2ioSC2bouj5+TMkci0T+V0Q1p
QCWGwnOYbihLU4qmwWS8CIHuA6e6jD27Hkq02TZqmgw0oiWTAkFHCGYaZtLs8Cs5
SsRZ7sMUGLLPNxyn4uQFiEmTQbMacBausikRWKiFLKTv+KJyLu2gTUFwxjQhMLmY
qjjyU/UuaE7Vu7xF/PDo997/btH6xiXyc4DJs0J4qlJdI+r0GQv5dgVCwT5pm0Iv
Elnl71vKVam2uFiFE9uHO1K524xDfpeLZnSFQSzKdNXNmgXRZc6L1wTYao0p59Cx
P3JWxpcHJh19qBen86IJxyOMKG7jsJgV3crm1ilBjL74aSbendhe+wwOU3jhgUJb
iwThB+GbEQ/ylZIlPb+5SRN2J5qQBiQgjvYYyfrNLP6KNEFRIz8z6fC+UxHolK9a
0apemOERZDYsQzvpxaQjpgqNaILohHItn3O2H2iaxXmWcdI+pIG4uiHmNI/NbJ0h
t1wpFcgB5Br3tXDl0+/7kJ6Zv5wEavNzLePvdSttAJk=
`protect END_PROTECTED
