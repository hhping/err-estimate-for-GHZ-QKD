`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fU8ICHl2EgISTwpFk8biauKgfKiVt4RIJBFMzEbNKDbQuOwcE5R++vNdgu7YfqZY
yclPfu+uggmZyq6mY83IhmC6kmz79rAIUoNnHPlbzYF65CEKqwlwCbABN01W6CUb
SdeWDueEVKb7a5eqP+stdTsCLIsdkJpPu+QWOe8CaxRReXnue2NU4Dh7fOn50mZj
6d3mEKSYrpMXTcpX5PtdxBb5TFZyRNmfCk9eCzDaU6U8vqWHNOJA9mfe8Z+A0QKG
kWAN2BsmIep6BWEWvB95Rw42QnaEl6qAtIfsrchO4nW8/KpXkKtmiaqQM382KGaf
mgVX7gS0anJpDJTFDB1KP3sEMMps1HF4aV1y5MCt7AX8TUjyecm2tKuo4X6+SN07
POeUY2OIMzo44ah3GKo6C4+h2AA92/jDd6pxG0gzddLjXMBBQ1EBlO1fXRl+bF1o
uGVuLGe7Htc7mpPTfRv3yXq7sPa4Guk6U936LdJ7QGxW3iDB8yrfg5HipS2A8itQ
iSq0CaOp36W26v/a0OFrNH3fI/FOU4TbesIa9/nJV21/aiDzTiqvVDnX+By8u3ef
xuKPJZsBSG1cnHl8UdLyzuu3RxkuoqrF4bkGWu5HBGuG14uQd+oP6vwOhyEQc0BB
BYhjgB4IAPsGfUlk60vG9V7C/CLm31qS45WPeW0ovvSWhaWi95eDVSaO2d50Sxdd
+nPSpQAyoVvuisgvAntu1QGLogPY8pc+sbik8WkbKoGvKNnHWvU74/8xaO+kOWLC
LjhKNz4fhFuJosqvp2G/vioqlxzM99yYlPPTTycxTmiBy03ENbkiguHULtiJ8PWR
RhFgbWbuNe/KjRKx5z0UI53riKAO8H1ukxR0Mn7G+uBz7sFn8m7QWxonS0nKVocS
Fyyn0uAw1sBNsyZSnX5gRf1GhU4hyscASBKB/wMNdzSeQdvRrnoNdIRPwWMZKuHs
79UcLGxeKlHjGMdoiSxtXh/5K7FCYCZKHwFb1582rNQ44QOtfgC7u2+Cy4S4yhmW
F3I3nXF1JSSAmRsVawrZ35pFAbbJswCLky6IM+j4vtCbR1tc1PJCkTWE3sU6feYV
SsIQrHlakATgRS/gIvXrMbuAeiHUpyoaupFXtxYmy+Xwo0dyAhlwRCtm0cC7T0I+
Lv4k+HTS8ht4/nCd7/i/kmCM8eV7osj8nrRTL660K7PL+m5VDcfO/R/meva5AB/N
SFZ/R+rbf8tAFkdFeWFxatfRMlIIVTZj5bwOcYGaurREVfo2ZZlx07IjI1JU412C
4l5jAF+TAriywtOHSWH0g3tLQH/aYoN+qyg1xYUMZA0ewzTvlQ+vuw09siCeCfAo
VvyY0oYDLyEnDhhBxvYF9A==
`protect END_PROTECTED
