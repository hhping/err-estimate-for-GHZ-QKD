`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUZAeCwNa7xVmzLyMJi5sXZrYANy+BbLlQm/TyH6R9fDa3e22gw0RfoNE+JT6VJM
W5LDhDPieQ7YK5sYXg5ggBYEZPpXyWbYQeEzXzQVgpuWOXCrZMXgw5ItUuAlThdi
jxyl9JdLOwWkq7aSFgKVj4eqmK5RcRdgHHNlURyaYrxT1bAFb3+Y6elr6KTcS9WR
9EOcML58n0BdRZ66Qfq90uEoZKD/35PvUR+3SqFX4sIk7YKkILa1eHGRT9krfhjU
aEiVS/xuYQVgSpifDgg0IA4uUKOIpb6JTaWmf76hicioA/8Qr5zufMULgn8I4+XN
4uB8phnf3bAKF2rilVDRk2wYBASvoppcbFn+vNEqYY7xGJWjprUFNfoiANbpdQFM
CruROlKfc2Cv5E4wJ0qRSLGYlh7YbCX/1z/VlRY/64Cop5BWXS6V1BEZAFWMnyjf
5WiKKHtIOkAKWYyEe137/eF9odo25Ws2RInYoDUGxLjwX5gLXB2sVowA525eLAeP
UdZb1zKJ0Yg32Mxk9OoEOHIIcniq6kd65cEvXL8bhM8vluAdy6Ev3K0BdunlWTQH
EST6mhhd8VqB7EwGefuiiqI4ddMofNqF+PE8sQEH8wE8Em+eOJANjmBkubMY1PTy
RlgShoH4aDWLbG4YmbOsISDpxasTw/LkWaeoNQnnKzfHHRCj6GYYXxhTdOyxlNe2
wXFTd6OkE3KskbOLr3KhIM6hx5q9sJmqwfIc+fKnMNHrt4MGv8E6mLmaKWZjmrvz
Skma9xXwTmOoko/J2GXVFOIsgpzoP/xoA0Dehw0PGmuPbCxP7ayPd9tTpJQUsxJq
+WtCnRiTyybchO1PwfFB7xId9vJm8NZuYCbqOx4oafV6Y0ukYFF0yLIoj2dgkKI7
ZxTFBoYsDW9oF4TXLyL7B5Cy/o1pMcn4CpQgKlFa1xN2o7DscnpjvQ8VgK3/15/K
lYJ/oEAgS/I5M9BR2p8sYJVlownZAYx2TrTfbGjkF0uMq/lf3EzcR/X3PGm/2TyG
hzRyBJORb/rY3mH808DrrpiHPYdqOvLG8fw9/9D2e0Z6eUsiUFz+bUdnwkY7kv4o
q7BV0hqSoHS0crqFosC6q8q2Kntmea0lnG2mdO2LJG/uGl1g8JQmjfF5robc427k
a4qCCIKxRPxWtsGVVhl9MxooFXXiotAGS2K/1Rv4H86FyReQIKFS/U/TetYRN5W8
5/20xK7EnF5XP6EFZq4tPM94Z46qqfiubJY9BPM2BbDtsur68wfqfwtwEvaxDXJl
eNIPYfnTYYvtjLkCs/e91qQNM8MI8p4BLvNI95NpItQDpIScw7aECghPFvluhGRP
vk3gqXWLML1B9lF/uJqojxaefMutibv9m7pckPzcoavGI89H40bbN93nvuKWVKp8
Nmw+DLmwJ1SpDnmYQjsG4LY9oHvCEhZaBmM4YFIuXTLP+syQh60QzHZdZq2HUxcb
iulmCOF/kcXVm+Is0spSeDtu4BYwSMqc9ZjlC/Tsap2Rp+f+FY8/0x1t3EJksFFM
s4LyjoKsIAz7S9yFAIIZTYoICExcPRXu49hbhDt59BmOmG3Ejk+p6QNLUHBq+1Nd
8/99pkGpaBSFyvAhagvT4TaevQpteZ8W0TH4b2ZnZ5TTC3EzVZVsQn0Qd3AyYTIB
jvGDpQP3LO51q4vMFsspAjaGhx7W5rxvxxcXjKcsXJ8diKce7dMxrzUmhVuHabS2
edmVPomySQH+aVhU+ane9OvwdJHVW03goEzFJNZZbYOJKGC7Zq+ipdvuG1nFCm0b
pHA3ASuCx0ZY0HXT9tzfOYlId3PrDtgHYHAE5pyyqDZV95o44puDk8jHfT0e5ZDZ
G35p1sJDRSkhDdoSS77PX/Nk9MxkeTlhO31R/v9SUVHy8RhCHXoOCiZSO7es3Lck
/JeG47f367sGr+nNwcnHOK7jg3E+rnQz71ICq75bE4t0YwVumPyUbUYfhoeSZSqt
5C+13oPlSyLhE6NZ1vjNIkZ2/4gJfgMBiOuh0GpN56Q6lXsV3Sa9uO75k8FYYgfM
MJDEqMGyy3F7R2AbB0KFgye8C7xDt8zQRgY2P0tiZU8Vcb6to9/sMlwOmoadxYD3
/Do2t6hOEn3V3trYQbvLV95AIfBIwQfnJuRCf3R48da3Kn6Nnx4J4hQ0Ex33dCgw
`protect END_PROTECTED
