`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Sg0tkfw1eOGWZIQtpiWZyVumjvLov/6av/zkGbTeD9BSMzqWqXo5W4IYFmHRZcA
rYI3LVlv8cKeg6oLhzv8gHZHQtBOqkbmkvGS2Gq9FyW8A4O1aHFo7KH1F+/Ssl/X
Oxr/eJLvuz6vOs/ant1q9QLmKoBMKUmjX5Jk1fuKp8y6QpOFQWkqeXRcdZvJbyzq
OJRWGi2ucdxLGDyIO/CD2V5aIBCj574wIPc60gK8Pgd2zuMK6z2c7NuXzMZjBzuy
vu0hB3LLpmorliAo85AB8h9JUJaxpHmSFxaO+bgavwKQUVKaf2ftDR9BSxEv58HK
1Hz2c8YFZmeFjttFSQV6g7LUpZB4LfdvFrawI2ImkZ2bpDLmdYBZykGdpmuP26hm
mel4mZDew35o9LD8Pponu/xdlwCBVNeEeWUBJHcNwg7jm37pYlXyAAbzww1j+dpj
yH2YJIEcgUJdNNFg1RAl/VSJhQeoxkoERcDypG9SHWvT6/F8sB9ZgiR5obQFpXQp
783cuFy5IvZMPN6hx7ALq/9hb9H0XNjjw7jtkDOviBQRX4+GiqQa/duJ+pNLWym8
8hVLbDhRTKScefKKhRtaMA37tmtLk2+MixlzfJ/F1CWji1Dl3j4GU1iBlHxsmJ7J
knjH2UaEvHRV36v9Y/zhyR5YJbfCptD2A/QYFWE3YF/b/YMh9eU6/Hc+rZo//aU+
P57z+BRj/xsturdDzQyU+1zCt5PW6ncrQHLK67DbI1bNblPRjAqlr9eNEtfDNPsM
OZ+9nkbbiny8n3cTL+O4YoEcdGfZ8agT781LkkdawV/M9pLyCBwI2N4N4MLasZbq
GqXOsJrewj03Lvr1JWUy7VBeScqqFGqWdu23Ax0pYd7P0Wq0Nt2IJ1EAV7hfZRBA
7IhLPuH6csJSM3a98EU5nV0BLFmyy/vnsqbqQSHmZppDKFg91v04qYX+QZ1Ni2Vx
h/moWYdZPVSa/LMhIwRWl74c7M2VHIGpXtC3JsOMdx4sh8Ei2SdxKtEJmUUoB2Yj
Dau8tqpptlqgNDtZoeK3N0gzq/k98uDO1L5qymJebtCGAErQQg6GP1OAVlcE8S9s
xru7gtvHqFgkSGVqvk4+AGUhHfqmbn97Zxnyt6IYUdS76jHvwNWbQ56m4l4OWi4q
AMjCmHeziimn9kSZAPKksNkhH1gy1JDzSgvT/r9+xe4oFyEWh2KF5sTvep2tmL6o
XpBm5L+1c3UupMiv+E5Pm/octGjARmSVlW2FAnidi8jNb0Q4ZCbBr0WRLmrNdnp3
VkoIMCAhTcj6pVKITy7vuhqc0w7Rm6CfvBCLRQ+c/Nl4oBGm024Eouo0P80DfXdX
Qlv4rYP1ie+Ica8rH3z6GuD7Q1i4Xl/rYkwT/Zogwk27XWFTiRqcw5fn2BvjKERv
3Jr2ISW2yvhVnKdis21bNKD6X76WxCr5Ft5C3xVTe/gBPTqizNVfKWzJTtRl+swC
AxWJuoK92LtJDXPpupbNtbijsaVFLiAh9RnaL7o6PTKxWP/3X7MH/PEy+Dz6elDb
GOGfLgDv/GUM5MUUZ+h8zU2/RiOk8WBAGOESVLahEhLHXACNr8c7YcWqBAjQwPuK
EWB73nl1EeJaevNz6RrLw3RhFs22puJgtVsMUBeVCYcyQjKtAeLBbZqxKh5UapL2
x9zO/7Tv84aiL5KoYrOiH1rIQPG6V5zRWdhbUssTusgAvI+eMWA5bcpFS4j509UC
Wktj+2xnpIWfwGzpRUXVSNqzX7B9lmGaDGVeHeRhoEroAJJT0fYl+ConCorgW8kF
YJLSKO3AZZFPMp4oZ+br20F3UpgdEfwBL7aMbIcc9BKd5fQxAoELg43jcdNNxJOZ
9bqwcTzYPQKbD/KJOn4q1DFyYoo7qqhI5DtacO3/N74ioVZlCjax0C+sg6CBNo7B
U00lhMGFGHAiIOwKO5sd8LpNFe6NETUV+CKs2KFAQaJJOArAzHWaRfSTAcntEiOr
5dxXyWW54ICV4RN1ip4wjX031UWle3fczs/Mh0NtjNSCB2VQfve2OYLuET8P2jYU
Tiyi6COT4xFlUEVShNV2bb9gypAqunlyysBe5K+LlSu2Ao1+3A6JqX37pnAC863d
crtekupZpwbZaifHZAhcPxxdQOt/6UEXmX3iXXKE1NYs5co69ay/nYxGjw7XKiK7
UTKM47fo6ZJnKTZyS10VPubDIuYu21Gl7bvyDOjAM+5skU9b57h2ed9fvZ3y70Sq
0++IJ+NsbtjLERdNF2bxR1iEGoPiAWqYHIIx/F7mAWGIIh/hhhzdQrTt6ZcH/Szx
hLGLdXlzUTpd+fP3Pe7/Uu0KDHo6FkRP7GQrbx1A1Zx3Fh7/GwwbeTbp1I36jMxn
Nnscs+MbH0aKQFSUz9gEoeEZiIoeMGM7bvfLCZg63Sq3acpOeb+5MvKC1G4J1Rqx
1AIUZQbvqjIzrZZpHVSVgfWqP1e3F5+/niXoMhKOGg7zvoHvbU72CLgyJAGqXSXJ
CwUNXr/XWIxc+7bduo6hgzj1JmeZtM2QeGLlTU+/RLJ6KyDzgsj7JUPh9vJikYmL
1MTHH6lhSBpocS+TQjeKbWATAWmXEE0Be9DCu5uqmZNSs/I8/m3tD9k0Czs3y07H
F6yIWDlT+++blaSUehlWXSXIQYqgSJ1oVPeh2bq8wjG03UEnv5E1sXPY5EbilZ5e
7WWvi6c0p2+DfNOnKxYrx+7cJN2DqrpfA827afLoLIjhaTQ8b3ri9jGURlYrgr/K
VecB0+s8I7SeW2pp7JAQwOzyIzUmDeuVCDXMfZAGS71/mnMrxcYiK3QEB8x1whX6
m8paTEFnrYBG6r4OxdNl6DSTqGYMJYZDYOri9ql+PfFIN0xLvHzqwKDOf4Fq9/75
vj1Be72vkS6F64XGBCeqo8HikWnU6bDQEet2GkOHLfXi1D6J7QDEbv+UPOzw+0+k
fNeEHtPw7YJ7MqZgiTgNxSOR9MZlUwRjYFAprCGqVIG5I+AWYvATWnfnf9i3Zihz
N/pMjhDge5EIiY7XuplCbrrfkONcwtYiO1no0HxqCp/B2P0NOGG4AEHj/e6gMsLj
4K/p+RJO6qLZw6er/1wLSkmG113qEvAljx5sIn9YXtCPwv4WuTMHIixCmewEeXqE
lTodJd4dGrADflqBzYcFVkxoG1fe5jDlXgJnmDRdqaT4frdSi61vF9nfq0MAK9Nd
dkLprWoWcEiHFYwRdXDpuI2vwGrVcVQnKX6pUknE4uCAGss4nPM5825Ju1/29m41
Ac1v9/daqAfjxoapNRu/E9pcgY7tutTT9BAFO45kEt0ZE2r5s5xBPBS3QQlKWyTt
iKMPUzBHJS0udzY6R2nPeGCHfSoBYfp6bJ1UwvH3fTr0XzrgWA+Axsy8oNRQeuQp
3tQ/yZADC2qiMiOS0vDCaWxzTuqehd/3CxEPlxFjYaa4jKm9wL3gjpLJvTlz+tyL
SJ/e+r4lXBjtLV7Oibf8PjynJ8OQrF7aJJzHv4Vw2qXCfM0q9ieyOyzyYAztBYSp
ByCnRZnK8aEkUDLmSuSrZzQSeGjY45SjsHdEhwGxP4Be1q6mlKseJRIVZn1oNkeO
QoDImg6cKc5tQIcgd5CQ400setbTB7nlfmNO40np2RdAAW/6503SaZ2fopMQvHWG
MTascGAcwLxnLTWqxyhXy6fvlQxFnHxwsQ4MaS3u4w30o405Bo/1wztQNyKwtRBo
/MzDYzCR4faWD+uq+RLtU4DmxMjnU7q4P9eXfX6B2bOrJJC84jYi6g5YXIr6ajzY
iu/Zo8eO1tUJiam2myfGWGTbbF6z2/HvYuhsHqskTkCCl43nnpIkQk+1TAWQQz0H
sApiqXQ+X4ommsL+Jt6LUGuWgK5/TVulJ2QCp0Wy9GerPoN7xUoZezF82TXLZO3e
MGFU3XY1MHn+QEG8Q8SPUmIL7qn8QZdd00nBu5N3gwpzidY5z16qIetIQuUrj6m4
/SnkICEUBcUs6b8+fhcPwXvywA2TTAKERVB/cnSyjmNWFuwd20oVWhcT70FCU1ys
k+EDLB+VxQWlicSf1ntKz0iL3E/kRTgAneZ6NLwh0VBGztnzm49Tn2b1kVw/LUwm
qb/DfqHS4mZEyoZtprXINfi8VayDPyfI/iWfECKB7t/W1jyYHXczAAkGX9db95h7
/7dprz3uMPhjZAu+DYmb6utfGlB9J9rnJLHNq0RM5BkTCzPZAc2ZTDI7UXwIJKop
e1t0SrjNdNYFseJ/8VAhFat9bMqPE4Yknd3mQcMNUv1wgRJpN3P8HPItHXWpADUz
KKV/0drngP+16EtP3j3b9J5KzKF0OOvP3bJtzkl+tMa73xkTDQ8yImIV+6vXCoFI
icr5JdjsmjHjjlK9IAuLwgzBpbOwYE0V/i9y9rsZRQe9LCcCh+ydlfPrvDVzjmMi
D256Rfj5j0b85SqcnoX7zoU6ELDcsscft81NbCgB5OoLIGrJdz3X8N9VR+HZwXjM
ZH8Xsi2MXBkpohMnbSzzJIrBHADUQmh2Zs+bqRqFFt9dBvkUGHfc9ruIxB621iSq
bsjNFmzfQfH+pzSCPC5/eN1oQrtOEkcwMxrsN02Ge5seHwix7BgogOMLSSyTlIRJ
ByA7zcBeKiryf+UiORd1bEoLMZwZJaxT+NKwMzKqg5MV9f6VvEYgbUxLZOeSK1MG
SzC+Oh2P3Y5ydE3b9nsOIrbRrT1Ux6XlqB8ux4TPEmIbvpfcOAAgdTZcP960N73R
D7tOQxe71rheT2lbDhdOo03jav3iBrBqmOBZQ5/vbr714LnG/S2HUeBrdSWC09xd
lepTbl5+WdkMl9KhGEfmdOnhdc4IHC/vO8DeiwKhMDenr8QbR5aeu0AzFcdhwFw9
phrmHD5uw7koQLa+086VSSmBJ6sRhLoonZ9uu2ekQJa47Pb7k3fbIm9hY8dSDbah
cO7IVBAJHCumyCjwHvrKx4k0z5kgcnDpgGxAXSy93dQeTavdjnTLIgs+GxJ0/mkK
iLgEemWyuIDvtmqBoD3YD+V1ET6z+IR2PeWuVYCQ4707iUdEnR3lemNsEDH+yrdo
YfKAwH1wvT+3q7Z+5Ut9LRZ5CfDGpC55SJbWbdNQ5mNcMbyQOy14DlUbhj103AWo
22fEk4GQd9CyrGQadrIrwdvHO8CERhHupSwr4NkIXZ8OouTODcoOIjyEglxYaDaC
72TU16HCJaeru2ctovgfKNPQwi9Vg99KHt0+ES68jCPbyoHzeH8+0R8aD4hvwRhk
VRtm2TXuhXRIONAqaBspYy1OEMkuSJfh7swQR0/gu9Hy3KilKz4wuMo3mwRWAXbr
A9qwqKqHzNXNGdJqJ8HmVokUZgZ1sZQyTv+QT+UT97D/n+78Y8V/6HaZ5MKp3wRl
UQpswRyqw6AtMyTOuu5MVCA6uY0B+lc7irggYbv2Q3IZrjZeCkldpnqd/cekFO+5
PQ7XhbtrONPWKLqRl4aY++WhQtxtg6Cx4cRtgarPmmbkImvKyslzQKjG1ytD9n+C
oVLUu4KcYCFoVX0fYK5OuCQKR/6s8YcrjDB/apEEG3LUTcHe931eOhItHDDaalIS
dZClsTbiufTWN5Ts0Si0W6k6pINoOdf/7+4y5+2QzFFhe5EJ45SdR0SqEhayI/a6
fAjGASEETMviGz5shz8Rje7rrOhR1Xd8/GEFAL9S/NLWmmNuiBG+dltswyZTtPsk
/ocODCsx6JXg/L/bbPFie/VsPMu+VnRBDEvnOoTYqW6ya8hMXGDomIwFBUTtXjKo
oz8pLJ8DyST9odn5FHZ2GTIfkybM5tNt6GD4lECZanPU+nC0tgOC/LaGx93VfHXl
qNLkYfoxDup/dpcqY1IO+J4hHLxKfsDDWckEO68rNac18hw1GxECd6UfRD0FxL5t
nsALymUwICWaPd8zgmvBSSAcL/h3Sn97jgJ9LA8tZL+Cwfr15a6aSutulmhhtYyx
K9dQiafcJcpEU1/ElY+FyPYNxhz/zDrDpO+SCTUuVWUYd226xrj5MYlvWkELa3KJ
92qFDHKu0POW3Ef7muHpkFIAOH4WQCxliXhpczfYZ4gG5v4E2Q9+2+D0Uy8l2xdo
S/9FWsIEFlLQJbj1qFQpUrG3rakYV0hNAsjnKO1Pcgoho8FcQOIs23EJbmXARTKH
9we4TqeKGp41DsqNkvce5dARM/YqVF0+X35ApbQ4exwiToPzWx1Lnxz4dWocTIH9
XiSX7AplTrDitukc7wNnRm8pRqXBruCI2bgv6nkaTy8NpgCImKNootl8wSRrdo4l
g7iqINN8dbJyqAYcDGlpmfVgTJP5j0pmDF8a9Wwk2PPEUD5KKrxfGOWsu7Pz+lrS
kn92Cp+75d8p2JwoXtYfOGV3N3aU7pjINoJrX6+NBmQGx4JkwqwFH7GrBhnN78jZ
rqFG1ajfixkgbZwegEt7GlHJEEfWJOBNe9oeRiuJipl/99f6S6bT8dt47HNtNs43
kQIMwHMXnQw4eXQyq6YAnggewmZ2qF5Yt/ZQgLFHkTiGDHnF7EyvD+69A0Iv1Kf0
kf1Vd/jIU2gV9+BcIcJZiTmDNV26sA7l6ZFP2GAnez387xWWUMOvvVaMXEGqNv99
DK8/l16p+3NiHuxXNad0c02FPuaISuLgK1C6Bn4wt3rWHp4y2H8eDEnWG0oZdrua
9yctkYJvad/0dmDqWk03hFbDhsWIbOAGj/JgehSDqb8TT3arD8/QAfgA77vFyLxA
opESK2kzIPtEzrwtvnAfYdhgv70q4jZMf1fYnhFtvyRKR6fL3VBYBWQGYwKTiH51
FmDrI8gwVmleTt1IBHHnXg8TOnFNYzweTSHV8ja4sPDZS/2tyjgrbheQVpQyjadx
jUE4/vea2Qq80sbYGkSpjM1DYbHJBoFb3/+ytyo0Kp7TasyQK5yB7gExbsgeBUeY
KooXm3WzXFfc6kXDwjlATnso2cV+BGFD3cEZajOCuJvgAKYNo/iFYY5KGDrrKe2g
ZjXVkrG/x7rRIwAUFTBUEj82K9l2wqOMgUYv93QEhsREZpL1Wqva6mek4J5zC3sO
F6wMbI+5S13D+FETac/UelBJyCuK8mMOS6mmEui2s6VtHAUJMJMNE8ZoJbFb3NsL
4Vne+sZOSO25SeiZ/NIx7SHWWu497E/zyAB9fKsBSge6FfINxQ4GETbTaLl4hu1i
J1vYUV5r3AwvJHTwAh/agWRpVplWnHMWnPM2ZbgmcVrG5HeFODuUtl8ieB0UPk9r
UdeCSosUxjLDSFp1UJgsEWG1yNYFiuwuVVYfDxVUSbIBW8b/RNp5m9cHjB03Y0sH
Mg1Euve1fn5JS0k3DFFOzHezDuZXEMU2CtYjlfI1XU6n/R1DEdnH4FFlv21Ksi7p
mGX02J7rDuF9LqcWXFtEuVnGbFWDFcE17+EBLR993HJqU5ycLtBo94ao5HPtWLHz
H1Edpr/Tvo/u+YhRRn3n/ikovXvyGz79PEq7G55BM0qs3+CEltRjugZaVQufUDAS
MgYx43F5pTZFjlu3M0jClNhJ+jC7TH5b59lgAJNsYLy/LVOc5m/Y3pSvG6z3o/no
MaQCekUbgc5P3XJZ6TsNkpDn9UC3HM6vmNjhEyTbivygGNJF8xAtkbrLyWBuo0tB
XsfYSbO9UTTsP5zOBB2uBvxcm31cU2cbfL7ANUlguYHLqvUv9JCRt/wqBPdUeWsQ
l94VtqlzioS6ntkYC/JWHzquA/t17or0egrwy2scAllTIjsdB7laBy0GnTnzD1Q3
CWdAH5EMI7xegDdiV8RqmP3PnznD3+VXId9dJ2pvBlpmCu3/y1PptOJKnSoG5S8l
ms5gxaw6gxifLlM4ApWO3wED/5LBv+awgYpl+066up+NMrzx3Jpglqls5emg1hqG
2gR9D5eUYEvEQ9FTk/TMrps81D3Kphop/UTDH9ou3Q2KqZY1KNTkSE3TP0/oniWN
Po1teoTn2whUU9DsP4a4LJtdhYBs7RGYS5GhScdHKvuapXKsul2IxNtmiVSwNMdG
ymXsm2LC+rcSYRACfjtOVwrt9E8H2FABv9Y+65r7lErqKyFeLNIUKqNj1j7lPzwb
qqZjdoargv3gmjjF8OsW+dXdBI/VttxLOThB4DtBx2+Yj5FD/ihwxjK4X8Ul9YAp
O8dPfNvTgm+jFe9X1gyCxUxajTjQq/R1jU59IcmlMCCytB+XRDwGcp2Oz85dIrUw
7WEWdhwSFygSd5AyMh9zvhpi+60Ag/6fFEx2sD5CrW1LrSwawLDJFb/wP6Big6a+
Iz+4w9EBmPTGhyBUxvJCJrmKYbdXeY3q+9FlvK5rUTHnx2AlaN7UBXAXBM4xNz9j
0Q291vJxoRRV1/U9WneflFDc5ZBYamoAAWx7LrsM2tXPxQ6OAkosyoH1D9uRLlA4
V/ut5AexshxHFweI04M02gxxJCRSNsuTlCRJDo8WcbxDHPnvfpiJ5uTAN6ptFG0K
W3suY0YUyEjD3sc0Sa6OV2Cu3VJbwsA96HrNd+d7o4B4aR3r9kN5PdK3WAYOjcNk
Jv7H561D6+sTyla2BieTY/claCue8tBQjOYuLVURc9Ka6MZEfXgZRSGi8yU4kmcc
b4KCQ8LgNyZBiQ7R0H0A9E+vGkn1W/xOfce8OL+ENMgH+rnr+dbU+3uwRDtGNeXk
ZpC4VLaot9X0OkU1bzM3SeFWRvWy3cpDz27gz7YQuZRtaVDtKMtWpzr2tLEws4ud
Mh653+/IjSye/ksmCt6LeJ/pHnjcy3krNbktzq++4EYTG7sIMTyEqs/kpNKXpnBh
/j4Df468LTPq9ofQI4/WjogStwLgi+NMUkK6y46bT48rfXznzwwzsGA1aQZau0qI
mQc9+7z9c+n13dmyfzdJLisNbghf/b+Cew69EiE3M/aAsMkWGuQT87WEGd5Ci/bm
4RwnmsTRu6bT8g5ewygCjxhauOTyXDa+k+RGt5dFw5xSo8VXIF3qicz9NeIVE3/A
HfiLtPgc41KziZHcrQITtWPkRhSGhHdbUd108/Wca0x5E2WXnotskxTGd/WfBuVo
uGYf5/MY5eF2DyEIUsZ293B1ftcxDME6/s4sOOKaW3x+5sD/m2+hOuWVSujzmisR
LsoWu5eCi/VIM6+O36zSRxIXiT0M4t1NZYPNn4KirKj5hPFMvoUzXRB1/3y/GjQX
0ZQZOMJhr7GmgynckT/naW6DeJzwMmTSUGZ8e6CeOLI5i4ENCbaBGSGzgG+WgXVu
ouApsxZzcCZuJZ00Y4tqOdvMv18Ifd5KwmE3hdbhDlwHlB8qUp8GJ4LcijluGg9U
BNlhq2KFAQfEO7WaQq2+zDbovvNupfxPFLuAxAcl7cNzEgAv8/iaW3bl2/WcZ7Ka
ZMbqhLa8wtIDydpsniT8JnoQp6aWjDWUXWMQxDTyUOxuFHWC8IQ0QAZ5V4Cnfah1
EsDXoefhXXh1t++Y6A4rIuDmxn96twDA7xP7Gb6x3jnyVZSp3DGaxgqDz0K+mEzh
nV5ZgypgJLP3FbXgO3WqKt5xZMliLFWoSFIUMnxUDHWca4wpXfdyVnQaVqON3Ukz
V3kEQR4sXm4D7ojWsNOpmCq/nbs5ebWtM5Aeza94zkMKFkfJVA0RyJ8FL32fHAGf
qBstyme56qI4Pdm8Gv21KHjny8kT2g/cQAh5/Ssn4Gr2tIgo4Hyc7uJGeH4OAvsj
7aSsEROiY45DpCRrTkT8gOh1tYA7ZpSzwO1wtV9XPYN2H6NHwQK3xbAx9AH7aDQu
YUhnnZb8yNOSpFlmgeqrCX6FzdKZXCW90GZt5w9Hq+xcIpEEk7U8SK7u2fI99m8g
hwEhEtx2DBBAJ71ddSu/bDSouDjj6d7+NfbqvtW9vIqEWHnGTAJrcfiyksHtnIk9
bK+/HirWXURaEaJ1nS0SQk5fVCPIlykDxjVV/26z27tbubEsJFaYKLSBAP4SKEAo
p+J3UsEJuckzCgAfK7N9RARUaYJebCKxOU6KFTZUb1s1xBVxaelceczVh0tm7CqL
EArnzLYA3nVPrjjB1LRPdu0lvXZ9RpjaVb48/dyTAtp5TKTlasFruu+xpWPN4oya
vygThqGswswS469RKBUEx26FVn3hiy/fJTk41bLTAVd3bZoQk5ytsHZmqzliqGdD
zs4gUQdk+TVAZxmEqzc6liUpCdgitQ3byh1tB6iG+bFNf1Z7/QvQE9PjHq2L8MFb
fBwUDzC5JADvrqx1ekG/k7I5z9+VblpdhqX6xscbQQt2Fuu0Y8hK8jRU6mxxGLP1
jihvXrIjxEw+zxR6bzbEby1YOIQRCKx8uYl78AHH9nM2soZ88wh/Zr9yDuEjZfbF
grKsW6Nt1TakivCw/r4FH9CvN+J94aIsHVPsuOLkHbly5eKbuBxbLP7TfuVZebOu
/cYwvX+1wAMhCVjcGVv2YDYez4HCuGCjO5UUubB9fiJ2z7LwPfHjOITkqqKqALT5
wal2nnqQzwRTJTtJgDXHoD16rQaNPq8ZyIhlf5nnMaHvH58Edc33DuArc27I0Gp1
9UmeYLHC54A7hby7fm6hfUsH4hozc919AdOIMMzXnWOXavEEZLDEngLJ9nJKkd+H
8oTFEcymcTtcX59ilNpdrSX8Bb28PchIIKszLsfx+9E=
`protect END_PROTECTED
