`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSJlDHEy2xI741uUl1ZrXpWWgjfh8Bd3R6TjXRiet5i4L1eA7NfPdGeCR+gpMLeX
ibMTOslKLrkeL36MBO/ziLcZMIGuUJaflgxk50E+QIhYOjScpGSGwn8WS2LIgdPI
53Z5vPC0A1vyuaXIJ1qNxUWY2VQGSyqamWriTn3xKMpVr9rfkD8PBERTk7Yq0tip
3AD0qQp6BTzHbO5GrxRORSJZF4d7Ukz1CngW/eak27mzELd1hh+QWmP2EGmCjH8W
ADsd5JPHgrqMZU+Baq0wQZ10pj4R0HvPrPJtxtc8ButV/psBngXAE6Vm19WCf83H
7xYeutTdbg6BO/qebgLGYQimAuWt3v8SKXzwGgqfEUo8DOc+H4C3AyiNcr/+3rBd
Ng1UoP95UwUd7DZGsFfr/ec6ce9Ggl1wwtv+I9TeXQepVCIAork+LIRb8sExNttL
O/ovOcfzGpGMFxHG+Gt9ZrEAyZT6TjfF81GosqL2a5ZwawNivp2jzrkVZa8h1fKC
JzLeo7lLkckmSL9ZutBP03bID3LPx4aSkKrtmjAOKlLrtSYXqi+dbw4aZ3RyUaYz
Hq3L4RGDE1dQMqowM33JtPjdYG8vvvFcOASCL8qD6+lx/oAfEJotJVeNdjxbdR5r
rbmiK9CB8Z9TzeFNDa9AtQ0xVgA0qZCQeCSL+uDSj335UKVl6dso0Q/qQ3zVG7uN
2aHLxcsm4LePrOI7JdsCokSWqbvgRWw0/OAp10bUtpmsEaGJoo3whcs3qosU5zh7
TYHETIh3mdRXoTOxaxqaiGU/yduzmBL65T0shUhm/xU=
`protect END_PROTECTED
