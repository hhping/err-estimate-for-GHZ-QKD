`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BM4rmMlG9Bf0hWuH6eGurLBF+gUERjrlr2C9YoYF34l4PrQ9y0Z5SYcUv5zNAYiw
3LiQ/unxrbnrCh57jL/yplRyXi/B+VHdYcc8g8aS08MOVeBqUd9/S0+YGCibWSsL
w/vGQ6BwI6SqZHxo1wSlbLDyZJhKsdQkAcw6ECrxgSVvCG8DEVNaqp/mTrQX/VhP
HTmHKHdr9YTmbB88DxGFNF20Ysn6/irLVsrxmRP4Nr5iZliOwwLFQJPB88J5OIiC
NfAQZF4y95BUQnZcSv749GtQ6D+bsdnV8B0XRCWOKt9/YVRoC7hDpc/WW/mQ+kTp
CtIYOMoRmBspfLAyHRdiRy7KG2rbtK0V5TkZZjVnNpR75kYJZLuxMQddhEO3ZTHs
GFGYTG0huu9+mVsT1p4qbY4nApuMSjW9mE9mkvP9R5Xq5kO/VJi+qOVo0HvF8mgj
ASM6NqE+Ev3mYYg+UFWrFhZf/ZH37yx2aE2s46+oCmbnA0EQ35bOE0zzNbMog11a
PXBAO9o5ERvZ36FrGulct6rliIX0fzMnbksZ2wnBHBTm2gDhQ5+WBpvoqLwSnaSe
ND2lNS863m3QhUCvVPoqbMlIpyE1MpJ9ZSees8yCELEoudJGh4HJebZ36ZeaCquq
a557SFm/tUOWRlGmXb1kqcAYxp6Hi7Nw2+lykh/nMlPL8u04nR4vXWdmbPKY98GN
3adH9xej0dy9UdVsvubErbv2hKCSmnzdkj4uu/IYIoVePfiIGnB+F8wP9MGuFxqx
41yGb4sUx3q23LGHS77aph6yKxub1VOjmIc85vuSvZ5/iNbHsaK+PMe6sNESl4az
y06dCi2l9OtHKsNKZfYRksx9kVbeHiG+QxFlmJ7LrsM1tCI1y9eKtLvMYjZQaUry
hHu+FxJemt2RX2RoB2Z3xL6PGxnVBrUULHrGaZj3cevoQxkAmT3V511BLe/JQYa6
N0Q2M5u+Mmu6xGTLCStIX/oai67scKpsTQVY357IeqUxydjXAiaSKnRBorro2iwE
T/CnbHE4pjStVEXBVd9a0jfZWMqYBAEn2Tocuwu6mSz6+O4ids4R9WOIa0ELVK/t
40TsJ5IUMEoqbWEaqw10DZaQpWDV1vl43KY0lIvYL9D7YB+8BqA/JftVySxhed/r
bep7MAGeS7hP/hKPAVZeFpdG4Z99f8WlD9IsjkwLqHg=
`protect END_PROTECTED
