`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5kZHdilOgOYp/i6O2byr1SgurX8HaWwCkuLsYwicHWvFdR1aATcMch2voPlj7hX2
F6hTS7B1/y2yPNiV5zLDz8bHi4xQbTxldvVbzUfnvzvOmOgovE3kwdrMscfKxAIN
XipmeWNjpVlU55wHA49g/M+kQf9YoW2vmwBaWGsoY2adL14lKwry6hKukCZWZLIV
sccIhYHCOHXE78kaMAVabRQPbnZajCD2IoybtP8iy4hzaHhUIzVvh/vFp6VBxPEU
F/SBgALBlmbzvnIv03UlnJzZr57I4x1Arsq3JpZ5vFv6Cb4igjDsl2qv0V8YvXcF
8TUmoW7dkE2ZESwvmZeKlSYFt3dJeDMsPAS/93cz3J793VC22KjwuHuVmJYDeqcK
3UOehyjFJpGJUPC7Ci/I1UB/8+gzDWSQMyRVjS5IeS6dxVO3ZBE4M4r6I1t5lxFc
oGqpji5v39A/RJLAxf+TVpSs3SUf1VCkShHoz4W9/36+VlUDBa+ogOnbQC5SPGKH
UFyoWB0BfBcIneJ8XcccJAAD6y18AADAZxXxJLrDdk2XVCqOJqF7WpZMcX4fkT6D
DtCKC4+TxFo3bS3hdi4TEdjHBXDO2V27GQaNBj5oY9OCVdU/mCEYXJ+eSsY2sCbC
cbpeLATc5Q+7jdajMpvm5RZmsafCyaYIND73buMFICHBSyhvE8L/gS/gSmEQiNEi
Vj+9Cfsv0pgx9bksEyemYSh8BtM8AdyNilV2xDUlKWAj9YhQ7hLRbISk/1Mrd0gJ
1xN3euSsRP+7eKFXYhhxy+J8SpzcETwASdGbbOBr4iwtH1hM9h0JJd0FpPC4c45O
zZlxXfsqz430b2vkbsOfP5aD3hJVe1LzgGSrarRHDVSPs1MZIuhd8GT395JiE0hU
tEPB3gH/klYOkM24ZOJMRWnW8e4WGhqp3wOX5/TOPFs=
`protect END_PROTECTED
