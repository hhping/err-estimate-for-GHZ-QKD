`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hg96WuQl0ZbqSAvifeE/4A4X/+TotP/nbhTJFhsZuCxiVRu5K1phgcMgLtNV9atN
1B+DOOOiSS2z/+Rh0bPDoxCCzELWhoMwf+MRb2QhB6X+P02ILScFWboypdf+VS4n
kncUBGAT1cmPjWZ/qBDXGf3sPLgN7HF2PJPbv/fn3CdKbOz2xL9PKfmC0MZdkNRV
Vqq2twH7idSFBfsehmlIIzl5IE7ZarIfRaVo/l1AbMDWgTJxCfIfjLwWBEcJEGkM
7hBkxu0fZEwC/6FikE3RoSckVPwcLgW1ncczWUMMUMnyVPLDOxPGjKu94r4BE2Nu
JC+x5/URxBpJXX7q3Toowlt8/+2/1lG9voNHIxzJ+jPk1Tu/lSs3D2u+LdfuhTrZ
duoG0ZsuhhlnHm5285aIh55Kyy72ixUTYU0ci1cB/1bf+EKi/RYU4XgjL071Zfrf
Kab84RsCOdk2rRHJjTsjZcUP2vnaNNVIqLZlas8eW2sPA6aL49Lxxs0m4vWLShGD
Mxh5ObHBxQ7TliQ+ZXuHnOasBIi09mkTo5VzoVqs8hpPeiIWRcuR5AAlO97l0lFJ
lpwaIsltAA4H+HS3490yUoiaVnO45jZRF2FdAcJhx+a7PdQH04WHRw0exHsXosi9
d3UtoKvFRYlq+E2Jo23U90dlOhDOVfyDG+4A5DEb9u0a4OvgwQ2zi3rI6G6H60DB
oAIJU6N431ZVdfJHAEIReMJ0JW2LG4jzIrHeeP1DnfPivJoBpPC2ey60BIugrKii
LVV3OzOWoqL86flzLPLIE3jWw8qQXuv1J56vwrPianor0cAb5U2Qi5G6dSg1pIfp
xaa4CTMcjB+YZr9z27Jsjqi6XQGCblWil/sAwAhuc/99Z5lqlihIvp2xjmvyD6l+
K7f2xMPAqX85rR3hCSObscOzcUvD2bV4c4JUQk8LDcntwn7IQ7nI0MI28EQ6JuPR
Nb7WH8GAjX152zwkKAXR4j+VjPRAAnSpwJ8UEjfA+i9UPeP/WbP3fAVkJjhNzo2q
VJW8Er8pATo2gozPVKbUel/2vQXuRI8Dj4ox6e4pk4Fmbly/vk9cdSVNenYx/UzF
SNfTt6MjqAbO8G+2vLuDd68dVUS/lFKLK+qoz++oeyKPgqyXV+oPSRMKQkNiS9t/
cDhLVpEHD0k8VlS7nOELDavaBEcYIrERQYaPvI4eBSbur1XPiCIHsddW7YO88JM1
m03iJJqCCK9Jo2+RgpU3bMstqBklrnfCyyHx3iYnPWJjgpQhHpXQ3GNoTNrG4Wju
p3SbLv5RmV4aujgwBV7dOHniKdrVTPCTO5YdzYsZ0pKakapKZndBFTKEYzFNt4xb
Kxgf0mFN1LEsGvKZbKjPYodRJHT7G0ooSEaufgPkFFicRqsEAMSV3nNwTCAZmGAD
At1JGzdhoLd0uo8VZ0lyprkGu9gKBQ25gnA0rY0DxkM61SYB8gxjA9pi/lHfrirS
3eCz3+oP3zdmfmzEQ5dFZ3wJDUG8S3bem9bvIUrnWPnTKeOoTTjL5OYqAv3RnH32
QpcESorVB0mdxtXbxf21WGubSqarg3ya3J8gQziKsGDV84NEUhzUY7VVWkq/SYEP
02In+oZWdTcpWXnz4RJKMPF4E0icrlVEoRSmy1OPqwR6ykxsDOGwvb+kHrpN3hbh
hOBU3U+9EVhAFugS4TmZastJsCnEWkT878asRTt8TUwgQKTG1MXR+LzpIB2UpCk4
mdhTbKkA87XFQj1WSm0lBJPKzCqRVGj01Q1oSXt23lJJSgwTogfs/08OYrCA45QF
wxckowm+0cytYfQVOa7grMxdBN6iYKJG8XDbKIlf6NH2chWPGtHgoEBUDWu36OJv
xXIPJVYhmuSMFzcsvuwIrJuDBARQ+V9gS6yjVN03AZxgvzAwYoP+UKVoSpgVZpQU
TFsBIjbe8JaK2rsAWcNW/earjbdT8K0oYxSq9UATqSjWItW4J+mO2+j245f8McFf
5fHgG35IXLamg2zGFI+HZHcEyymnLiUSJ3Xm52i7lBXigcgL1GGF8y1VnlWJ/wpg
O7bHsSPkS+pCw97pRrpjcyqz+vWw7L9yI3gg0yzG+0qdWb2rJTclVE8FtOTJXir1
r0YHfkXeF2VoIh3aycggo0924E7b30gTCUJXY8wpw8YeNmfsCtND7KjJ4vhm75ST
Z34Yc7fsXxpPPliY7QU6nw4lJ+AnKtp43uy6k+po5BysLNvpK/4DFoEIB1F1n0Um
vqTHi0oNVoViK0zdy+GF6qwpYwI+ry0ODm9cG5BBmXpwYbN2hUvXbFrqGqnN504g
kw7RsAppg8KavGIamoaLjF2r/udA8PG0531l0fp7Y/sAylVBmvEbL8sExiJVFeZ0
56JIT+iH1i9UzEUBHW0I6DvSa8ltCtZvJXjo5eNGjGNxp+zgXyT+G35OgKPdEayd
fSUBQRpU76sMHaovL+dN4JjTaCnmqJ6CChhm3B6b4p6knU/pZcjP3byicCF7XV7E
2epmI5HyK+rFxKlReLZfXJfHlrhisunxR68Evr0qeDIbVrjl9LdSlTfnvzo6zOUH
cuk5diNobbgu/2JuBAmwC9Disr1xdxSsPGfFjDjJhmSObQ77bs9bVVZmKoykYhZx
I3FENYpjGRUTHRPOkZ5xn4mQUrzkj3u0FLYRhbQWRMqBVSYYc0/zWCP71SQcgxyI
D8aNsdI3zXrbka645DyZ/NXJpe/mgTe/gaWG0SnX1B+lhWL8mXLkjs1sD8YvTV0W
6ECb1uZdCVvX/hh/d256cdZISfeMtwiRNu+Fxj+ou+G6Nticse6IyDUWsTrRqMrs
TGqCzrhGGUIXW74emuAHLvf7cIrIX+tN457mZxYyi0j2S0zIdobqWUEeyAUUyqAg
RynPsSxtBs4mOke8bkdNQz927ly882E+KkdDokFZ91vabjKOwbjoSFLP0TDtMjXc
ePzKkadXwMwYWLA1U3Eu3E+IX8odOPe/WUPR3y8enX6bohLluTd+Mn8BYisTG3Xx
ebooquxyiYoR06XcFICj7JAVDjtZAtUnnMq6QVMPnzIahzzb7XvtbmKyFneF5NH5
ShBMhhByR9fsaD6qVq3B4ljqbLT8AInUCU4YyufGDiz0NBr/2jnAi993P/ozulov
JnqfD3Atd+DJtHvBkr/GlEowa49G4RaoNeCJbj9UOBWhzUgNLau+Gj2HkUjSNGAC
yNyt0MD8CBSpe3K5g7J/c0TTMRJSlAO6ZYO3l/MBBzjIWX0p7j5q1x7zVrxBsX+4
ot1nEbL82afeyvEzblHVgn39S3lHL3XEAGpuIJgTN8iMC5IOcuozwBnd2jxoAbDX
mQj3AOvsr1d/2FHZSGnxyd6nokXPwQxr0decJ11PSHgGpH0kYD0U/jf49Ow7PEb1
QBnAjRuYX6p4ZUySuX7/uwebU/TestdkoKuXIhErgcaSivolKv/Y/xQzisYf4lql
AHxjN9jv29AUk8i694ec7p2j2Y8Cth+O6k9elaXwFQ6LRFrQCJDTzJ9rO9wr3idh
zXvSbHTPLShINO309F6LolcE4iVSqbG6xcJ19l4hjQHrdyaxwOVMzI+M2l/Tf3s0
Swbid1nUhI74V7TJrxSAnJcZazYVFZ/exK4e7ZXVHgJs62XpUwYMcEdf2r+WUXa3
cqsFghd7hn7BKPsVh+RQ0M7PI2PAdjyTJHPP8xFOBDZCxahy8qYBYFX2Hd5Kxv4s
COsID9aGdy1JeFBIHUs9k/yJGHFy8Uat9uemhVWGZ0bnfXVcFzIhwKYEDVpjx3Xl
Zlm5Pht0HBGUPK8zJZn2O4zzdBf4sO/t8FPuIhUxC5SPZIVRjFCVwNzoPygAgfpi
0gCq8IZOQefuSXaM8nj9eOd18vorLeDGPHHq6U/uIw3M+P+euPpidEp7mu8Kc3CA
YIXj7jjPTjJqpfkxt9ODSeSTTfvI+a2C93nGDLOo0xFGhW4lVolYh2i8QWwsFzRZ
Mu7VkkORqxeIgTXkoTeNWjk5SMHhYCNVeZMXxuYs6F2bVQS1/u9IJur4qmaUgieJ
WQTgzHKp1JkgYdNoQcIk0j1z5/F1A5EfREhb60ms1IsJ7hrzndRwLcPfWysbfTwh
A1mF0CqrYqnPX+WmfSoWY9sR/T7+I8mQdKRSskABptSb6B9hQI1BcCtyvMFqD5Wj
b1pgt2RyTsfsAgRTh1DSrCeAX+zVvWfGWxRs7BK/mwPV7TN/d5WsXso37J5+BuRl
+7+n8OJ1aIU8Ff+GlB1ALK7P57tRYat/pxXOEnJXPti4hVmsVVQom1absZ5FMUZ1
8YgQ4pA0YhrImO2qnnuDcFBs7IzA+jv6kBAQv9VIxWjDsZuxo/Id9Qtgx7Fc8Z4z
2N3CUUKq0q/53NG0Nb0xTFNoj4cffA3ex1TTplQuaI3vb/94F5BGf9NuELhoFSIY
BD+fzP2L3p6+Hud7t44J1ccAB1y2doceOhMF2z65YJkx1FE32NL74FsUEfc+vKG1
QX9eVsXAQmacZFoaP5L9LkPIeF0DPGcsuYh4FFyJcmEOCU4SPkeRDuxzc75H1fOX
sWp/4cecmwYcSMEpdS3mnyv5IWNSn9URNiTwF5Ut8JnBWBy8yhsa4LUDTEpunLKt
gkuahG7iqbayO2Iq6QMili3hm0F7Pd+3XvLSD3AOfmJopded7qnYpYKKd9sgtAct
3K5JjQagocOo+xN9U8QpWRvk25UptOxRxvT3AcWY8eQ2oSXqmEFoGP1xGmHB0kRE
MnQ9lf6dAvS//TBksyakqCbOPPs9T+6MY74vVPNhAzsEus5AKOeSxHrFBO8jTq1H
DVgiTw9NFIk0Hjf6c/2NVGqQahtHFGkSC0D86YvwGwr86YwA5sCEW12ZbDHU0KgW
TxphVzSez3kJ3/6WDDsQJC/ZmX4Jkhpyubkapp9BOyzTjcCagDtQ/q3xzOnEQ2Rx
jvV7fkUNO+YzTCmR57xSg01o0mSqFQHlyvtgMhw5/2kkbQ/RpjNYhDlqoEXIW9Ir
+07bcXCqknZikQ8dZ26RDsIqeqy5WTsid2EAq6LXnoj3FbXRNMSVxPKtWwhRJj8E
1FP3kHzbMMmSTxcWnhphJSa7Hxry5W/8HzOYvYx3IHO0McHr9+8TpHopXES+Vynb
Ybuar/juazRFKihn1uVv4T0Ta2s28Wg8tU1+ZB9xh2Vz749H3Qq21g1oCu9XeLlN
Cq0+61EdwEWhYud+wyp91T4ecVWzu6yo+WKU8eU704j+MtFDiloEXGn9Utz8/xqG
Ie4TErm/OkwVHv/SmmQtPTvQbjbg8VczBnSspEPZSW861YxezJgHE02Igjb6YqVL
8pZdffdSgOWLlK0xSjQx64/4/Oy/3thk05I6SY/kG8Ny0hCsbl9h+6tMyev0xN1E
2QoIpcTstXeapFkTQPuTFApdYYFs5mPVPyUf9W/lvmzj2KbhGbbXfTxWeaRTQsEJ
OSjo89QaO92M/lB1hmdzEs6irSDpPT5dE02/T78xHq64TC9e/nyjDR1m+m57WqDc
mIk6/cIC8j18pw9gCXqJz7vjOtTP+ZqvFqTDVlqHYsxkWKy2sTaWdJM3QONG1ccA
H7cHtarZ1szLZFwxYbwRQBa4CDcZ1B12+LQNwcy7g1fg9035BRaYCa3fkmamelJj
QxzJVmyj43Q7k2GsUDeVOePfayYJbtXXTxaE2sXPv6ufM6+S3f0XATp4QEpxO1Kh
Rzb6uZXFVfil+3VQAmlOA9Ul/q/cgQ0/CUL2ucxriPk57EQbEb/mijJamaGhwoLS
f0TcAYuwSGErb9pxAjApZFbo+by1OoSDSpePrcexQ0mhcNwTNZBJhchBXCNIPgS2
BI1gG2kptZehrZlgwCksfr5dkSWrwLdLVA5dUd7g1KmSS9CyDvM2ipm9Wc6kDZ5o
jE/hT+h6B4ybdxcO4eFhcIDn0SShCgsRQnN53hSLSx/8DmdCEmU5pvs1WeilvuC6
m83msVBz3BkAq0lEHdf3Td0WhG8o8CN9Ezc3SegS8mUrp3qnOuCNM9eqUxepPclO
MRZ4D9NzP5dYsUqGgt3GdewxN0IGL1AiyvkC2FAilFdqjUJixNooxMN0YyGh7BeT
3lTpKwtVA3l7jm7Jvm0tdadC1nNoimsrx5czI0ksZ69OQpROFyCsqsxrI1EbUlIi
93kqGUICICZcIrTQ+YUHkxYdQ8ysy0+lruCLzlRca+gQh2MNVObhALxSMLJripry
5Ds2EwvdROBTNsRshuLB1cxkMYxp/den3ftyblKRsN8NCgkVDHtzDLEW9FzhNpP5
WI5B1A2dJzy5FZmsEzcWPGxAQYFVvgeiBeZxA3g/zN8uAKO4kYyI8TJWhrqVA7yA
qzzKu4ikHgyFGukO0tY6PRTxvaxqHUdGpwOns51V1fJe5y7Rxbo4SZh6/vXKzsSx
I/jrbHKiy5dR6x8QIWzcMiVNEzL02E/6EvV2KyXW6Byc37Dp3Xib0Dyx7aCT6gvJ
F5vuT7XGtMuoaxonGUWbFqYv3hWA0Q1W5uCCfXLYrNNPSGioBCXHvlIq+epNgxYZ
PSGHXEoQy0eiTWoFD/ZrPiFLQqEFPoHKM//mJkZl5yLLHcEy3/D6WU8d8ZAZsVyD
Bxst6aOc+tUvPP8nzXtzwHZR+sp78b/RYEspoeDnSy0dZFCBh5G3f2q52DdZCEs5
wPbosXtMm8jOHcytRs+vjdAjUzGDvDsLxpdDJJhIRZA7/proek8KUYdfthGkYiMT
jPpXTdT96AlmCm3Q0zFDI8YVi8VkearU79hoMzvQyLvV9gd1AxmCKV+JNToUpFiG
3gGzv3O2jxcuHCR9kJ2D4OKZ6rcN2XIdm9lWVmAkc5qKaLNYfyjrYV2ixslsUKzX
/X7JubxRMQ2L4SMXp7rk+xIRTMHbGkrGfR5yg/sVz63uBaH/jJKaazzrDMevp+v2
OX2wP//dv17hNxLQx/bZur+0yuinY3B0/0kD7M6qLzNxwu50tTCqniTN5bTIp+As
0UFz+pUo8d0GVEmzEhhcM20vk02o0RIzELX22FvjupIDQaEWVyZKbmLdk6/VW+Qy
exhyNDone81EuE/12FyrnsTkQcyYXIrDbqAxxO6j8oI77mA0Pasqx55cTv6Veugx
lxUMzWUpVCV5zgElpkURMzF4Z6XBd3Y1Dp/uVXp//KRqgkobbYa3+cSdN7j9J6hV
5tuUAVOu/+JXnWNY7WwDNNoWjvw3zyFYpfUQCI6CZOGMc2q9a9S24Tt4qJPNwk60
uTaSJU+QAyGawFfWyv7BZe5KE9O3f95wM/WWQCSzHvxo0G5MRUyCM1XNEybLv38q
ikZ2bHchBpxcYU2Ob6+YJe/LPkYBPZCrbOPlo577JybCccZZsacE5zTkXwHCkNb+
KsSnQesSFkzKQy3jIMFK6BmIuKcpL8CKGpWW5hOcwnpcyeuYwrzOPGSlt0BFl9Va
03Goa1+HsUYmhYnpliPKHKaTehbRjuHVIeloysc8d/K1g8ejlbT6iwDgIi/OB3pC
OxpdKxAA4Sc6CdWNSLPw0x53YmlHGM7c+zrbnEyqq1NbsGR5DCE7NNDtkDLwDNih
xoFuuoVrjpRuZKEC0dlsMi8qt6QUyQfmr7CCpWpnVWvGwp/PmekZDcXBuN2nVORv
YW2iDpkJLPqQ1DDysmsURZHt9k4qwUJZD3wEJZzvbAK49w4PnQZ3cF3C78zomv4a
KFrwkfL04AOea1hJRQY7zZckQQrW6iKSvC6RthuT5jH56988gvGpH6XlEIouHBxH
NCjvMgN0lJ8EYsCPwZTaMnbBRrfBxu+GbqJr7hh36K/6Gnfo60WRnHgkXGBaiG3X
q3bSwEfSyBKQXcSrzoooYS/qqz1DXWN15/muTdK2AGRjf2EbR+ByU/ruE6fkyrX4
xzUmQym3budC37vf4t+/eJFzB/9VlCMRLMqJmMasWoLcDZwhE1pcK5+x7fjGusr2
Tq7/NLV54bxCwIxdT8Fnoik4Z+OG/OHLKZx9H1fmoa+Lk7ZGPeipwOEmlPlPfKg2
hqS3jbyqrgk1mMcvzi4yNCI+zhCqTr0AcZpDb3eKg/vVZenfB2r2bPQY4V/EUiYa
OlP1pHQ/5iSwqJdFkEUmoe7ZZzsnycT+8qKVOeB2ZEbfMhAdK+WtNrHpQ3ygh1WY
LGmJOEfT5Qf/gkNjze7xRGHW1Z9/sC2tm3fsp/1ltdSecskBz53Wkwj87OxYkVe6
haqtFpQU50v/ZIWkc80Xjeke7/rjA3s4MJdVg+3i0mRiJejLboJiViRT7voosETR
kDv8SDfkvGPBh3xbbuwNTD26mfwhTZrLZ+QirPig2XahXQ7X+EMVRPOBlpnHXKjP
CQFaiEY2gbTmNMV2GCYDXhUEE0pCIaeRWuwmXeZmY1yg/5qFbUyvCpczfukwGWjE
JNBXEmqrLwnJ4dbIgSuFqIrZLC1JXVhQldqoeWcnJmwhQCK9Ek3s8y6mZsLIu52x
DAN4kDxJZUjiHM5Ro6ySE5vYYNTBnCgSqvUBNlhSzqGUxbhEpVyg/9/Bp3WvqSpw
6ZL4M19jBalhWq385jl6UB+2uCA9/OBGNGfQjEeiLylDKP0fJQ5IRTldEjQTUtVR
OyDISN6wpzq3nqDNPW5wmo1LGMSYmu/mXfgCxUh9lFLoLvVef/CXZQ5F2c7yGTPl
pc8Pn3KLDrHnF/TQwemBib0imyGyJJdIubcpbkLV0CZIrzkyTSD1zxYgzpuk2PsG
7hYT6ZAXCBTig1N8EfDtqhnoPzYQQgcn/yVM9DLyCtrvQqJhaM2oA85cGbm6DMJ6
LdTFgOrq5MxFu4riqF5Q3LYsGerfWm764wPinQmX/9A6PFAgJomH+6HuoFtCvvAG
NT3Nk07HJEVaOmJt9jTvcKxtDr36Vw+ePfGM81PGZK9cZuyrhBc9DB2pPhRhKMll
KxDBaEu5AEZeXc1XFDE1aRjEs4BCuqosG42m3tZRQtnEorjnHlPIA9gk7NKFeKi0
cYv8lx2cEOojWda7OoHvUKdU3FFGQpFO4vvxpo+f9QSuNvZxIHJJjnErMedsIjcr
oCb5/uRlvnKrpZ04EvXzd2f9enc2G/7BYZERKzq+NOBuySH+1GuQmZUsnLodiKla
1voJHZmMfEUABUUpHolYBLpUzP9++uSf3+SOo7I+fOedZ8zqKvjDtLuOwx8zVYGQ
YNPu0TJVLmGrvFRZjReAkuR7xRMHG5r2ktLY7GZ2HEj12vuhonSqSggzZEQu9l0p
I7TwXibpX8f5o1T70ok8lB4Un19hvCN2wLEbbV2QrDVEnzS4NH6gxlZyY0uwQs+B
8tqUzWCcQjnUZxk04g0XQkb0XtWbwofvkjChrRoZTCLpJj5XrhquHwRphjrprmX7
vOBQXoX39itFz6N1T+To78j1Gy6pNXiLBOZLwVhJgU980BOhwqbWdGGZ8rXuwdA5
DBUgEks+UaBKct+bIWvc7tQV1tbPUcawz2M/3M/07lU6lDoZTbaPPeKAs0loBuzn
b6VyqczrVG0w1781UuujIfPtvdvSe3IsnY8tZICiQLau/izfLjfByaA7Iaflth9a
qOPoiFAFp+xf3pVzhvqPQtoGbKotkuB++HPs3e0XGCO3nuhfkbrNwWuiVzyrmPCt
/Wq9mdlnDOAHWa7sIJmlq7EJgLOPAjj1DqNm4nuE8IuJYRO008u38qImm6A8hOl4
Z/Di7z4bNyKBMMapDOAl9OhhJMFmwRICu5U2w/nJjnsrxnsHnWINVVfKb0rZWmEa
8m6N9aRH//rx2UG7KvEW99aGTOJNfdE9pwPL80QY+5Vj4MpjC0fACqbeYQOGiRyn
2E8+ccRP+xPET4pjrpLc0RcP50JWcLoqhhiivgMOnUovA/3KYT7gL6mBmch1I7R4
yAOT1AwKQv5vPUI0hBLx+uDjBHBocyhHi4ZtaFUqN6dO9zZpE35KWeKaZyqTigCt
ZmD71h5szfDXzn0AADZO2MnNd68C0WTSL572491ENovmZyzlqTGt+MPs4gNezzKP
7V78D788XkCI+3086eVwdYwksv2Qmsu9titi9QlC3PgXZxCiiPcVDcEAw5wVQUL8
x4OqSYGhH1h4ZfM9sbkUYcT6Aawgwk8AA18uCQ8MbNXQVhK3Ck3AWvXivFUe7WQD
8OZ7TghdRS4EcKWHG4Jv5VfypWKEQkJbGM+EQasemJJPKFQTBWvtcfd4FMU2q/5Y
xgv2pY5xYB9aTW4CJiTvDZ71qIWFWKivYHdj7m9OfcqOrlnRhf1Eyi9O+/UlxzCM
nOQJCpT2mUliiu/7mBQ5hphHISoSGGyXBVrIyqLOHsh296LnxrizZcqIhOWfxbE7
FVVb9edAQrhb0Z+yAPOpFg0JiSVdHmalzkJ0F/C5a+e1GCpSSxdfNS1sQS7u3W8J
D2MYYVdzlSimupYrFCSWZpjEPyk65RPEVjQjewn1XHviTVm4kzE7Ryzd3izey3qi
Jkmv3ds+736sS+30pEjPIjEB1K/8Kk90U2WoUxMQCfsbQzrcJ47n5ZgprUDEn7t9
bsY+tMv/I54mKjFvFAKwT4zyk7fD1iNq3UabAlcbTB6OoJtxOTSxffVuZ/Z64783
ywqQme0qoWZXkTLQ+tkKwdPfr7FUbIvXe7VDUn5c8OSVt0NCf7pnXC4+DCXpzZOL
cdPRnO8pWj52sRkmv8iIjw8G2vKNy9/iJTZWqD1oCo6xy2ZNVc1yYDKqRSXzUINB
khyzt/G9YTrZXWKWfiDS8x1uGet9QVsaYO76hanvLOOrgh1Pa4vDuwUtBtPHxBVp
KZunj57bQRH0t3HI/HOyWhu40iXiT6S8yoakVlCd7p5lc4G/v9mwdAd36rXsVrfn
MMOgvgNNI/IhZLZbwaJj7fBFD8Df5DuqTw2XU0xWYz4RCc2xZqoeCJuoy1YpNg4k
9darYboYnC8HJnsmThGQcxK4f7hn3raKBRWDAftPCXbMPgILL5AH4IVCihUkO/UL
SOumKVBQCQc15/oNqWPhR9KubLQZj1oKlOJ+xGxjxiqnq+Cdprk/HRL3aASFzP6z
8HAUu/mjHTSNvpHIJtuydn7vyucBtTn3b3XxN81Rs2oS4NmXFNlKHjV8e1PsbG82
gmbwv0seQr+sXJ64Rl5wrpO807GYmnx4L485Gnb43r+uN4QR6pwtOKi4xY2Hskyr
P9E31J/JGOj1ERjZDkTyx+OPgtGy/zy+3xcP6bK1K4sJ2erEmkSS9HJPXsiaKvep
m2tUJ0rx3AVHqRGmZVffU/kSRXtYkCjBUts1gBH1Vkw6dq9Ttl/ucuPoXu/Y0/Et
dafL6QuTZZ9JwuT+AZ7+URn0TANuz0X0u9IiG6OOrGUToSdPXAKLI05BhS0iAJba
PgNA5eHP1K9ven8bwtm3OeNLQJuanWkgusYkyK/0PnmP5KwlZr930mn4/FYNqBfR
cu7uyA7vaQ4LwMiKzFe27OppNv9eqLd18Bu05wwRRSDVbRm0qPeEFWpOZYWrK9W9
/3RTDvKL0fgkVRBmF0TjTls3hUZ473HicE3WXSwYCAo6bGOLHs/YAbixG7oT+DoM
hrBLYdCLPt7mhmsI48Bu/ERC0NUgX7py6MQehvAZXACQjdY4BK49k1Taq0DgtcJG
FiU5p0YOJOABjx+zqFNum9+39jma4OxvW9TJd/YsVAm7ZAXolCiudotQmVhxQFqJ
+ylY+Sl8alu5J88ARHZ7ZR3TvGB5u1QZe5x54dKbVzblWj/9UmNRRZ6v0Vw3Rxn7
VtCUPUnA00P8Wi135gBnEhrt3bQxFS/RoGOuUi9e+UVedH/yza+l5y+H9bCCLpqy
Hv/XaG+hW/u50Xt/ONiey0RnxA0fEAwkxneXWbVCGMoMVpJy0HYXLiSBK+rdUnXB
P3G842yxwSwxE2ttZfb0xV5Eeu8VYoi8bLoSG1CSukeiS5fpOGLSeeQ3YDMJymOQ
F7NqvWW04kJEILDY9P0I1uvo0+pv806UiQ6j/qtCt7GUoepjk/DaLkvGoYoKySsD
CA+wdX3ngsFPocM3tWB+Nr3tsiXOc134QfNFLc0p4hazEylW536L3ldx7s37fU0l
Yo7VnDLpXx2Z4DzJLrXIGbHl+nMURNcrDmJ18NuRcCuNwHHXxQ68U2s+XRVZifXi
58o2sADxRKjn9NZJ8GKg6QRS83zIfuymoniwfufNGcdA7TjUomy7bVg9M5BEmzJG
qJIWL1Q7tVIZmKDiiNJf4Mp35PERDGclR5Y3PbCWM017Rs4fL4X+sS3c+A0fKUDo
CwRysdDwIEp2mJX1lFphRjV9TnqpwD/zHfu2OU/NVo/WO/8uO7Qqnmj/5ZPe50un
EPFQpGc63fBReuFQ0rzsY6FnMA3z153/KhrMPmiBly04sT/gXnvW9k/njxlH8Eq8
e4Gk09YqaRodRYKK/qgefO95iHeEuFeUHkyuFLlXuODo81lf4ky4BzF3afRTX3RF
PAs4KdQhKiEMJSx/vDK/shnj85L6dRCwFrRTi5Ed3TbSpLudBaqr2e0f8c4qy3U+
xLKvhRoVXIq5M8XgkEyOfe1LcaAjgk2+OTWvlR61FlqZF+K+CHkapJaMG584CB4P
bQeNSGjAfRRxAPc2FWoXR6ZGieR0MetgVD/91/fnSgnlf1reFuw+L02Dj2DI4/DO
eVosL6OnUxLCPIom+liuK8/Z/BP21YQG9o/cn8OA47UEwkgxFAwjPxCErbcYeZ4z
cmfQTQpbNDxm4myNk0Oe7pTwVJgiO5CZnh5rE7Hl06Lx01r2GGezkKVa+COcb3Q5
G4fNdr6qtdzIQ46ZjyYBCfUiEhQF+jO+U3v1XG6eFkMuX1pUlVtpRKf99PMdu79D
XNBX3QBKG3hu3ASbI7mvGFkb4lCm1ZtUrQWxivtqHlc/EoaPuKFKn2Z1OkNaWKNc
BXJ3TcMgU2H3KzZB1V8mgVI6kRE579lHYuh7VV1BiE2Iec4ATlAM16mKTiPt9Amw
y0vxinc9DrVIV0fZVlhNWIR5hdHj1TJNzy6RbteUxdIeLGna5hNV37uaWLfHnziA
5s0Y+1C3pA061ar9SVyBYAwt9Iwbp3TgNEDS678c9K6NG5RbrLzQhdjghgmsaoNx
pbRJaYmL3z3sDo8BoByU2cwhoBi+EZf0imf9cn8cpt/6T+AYEXn+6qC9r8PY3DsG
r5gQLrkOzjUpeqI5h3PkDGU3X2fApg0ofH+Tahiq7fq00Za9eXkNxO7bGlRwZsiy
OQ11F6KvmjVk2JQdOB9vKJdICgslmKpVxIcW8lANvqluvL2BIclHg9Ur7ATtLFdN
3d5vi99bYnfAUYGYak7l8/hrmudEhCCilxFTJZrEsqKR4YbhaYKeBUWlGU1AP82U
1nWF+5iYyqNN3MFmzZEvKbzoJjjwCDJayEQ6MhtJQLGRm9DRhHj4nRnTQCRi7sEQ
wHx8SjSVcMtCHh52WDAMK6MMw5e30vZMTmwQVuinblpkc3lYf1NG2sSgKLoxIaTs
ss2ulx2PtqBMMhEHmMgkzeWmOZxcLj/QwW3l5IKZFuSI4eXED6kR6pEkmXS+DFYY
0kZZXuNDiSkm5sUecMcvnwScJUEWgcG96GWsFGpoghxUU50+OXN2stDtdGRVYlaE
xjHX5mjg1krK/0ItT3B7qgHbdxeXaA+egAFASnqdcTkLahwVL5IslDQKuQg8Rsdk
Fi6W6W33e1i5jYZt1BjF6nHTAqYyaGX0sL7WH5uyWvGVy6xxT4Cfe6TqsKrfyePl
N2OC0DJK8X3J3G+R37ElhZT9GJaLIa8McnE3wFUvxOosLZlVpERf4ZkhDiZtQGoV
rh8pkZCajfH1ayIP4ePKOsxBZRjWrmZLXAq5oN8Y/TtZ95y5gxTLnBDURmEXzrNJ
7j9CaPf06GT4FP1UsAkKaRDV69se2Z1MQ2cGiToX5oSM92E7SgWARFT1YjXTebh2
yhcp9lFpcynKIWIlHh280mznpJq9b2tE0G0/pDgUhpGZ8ssKiy5S6PUCXc9U487f
d6ZwSdWNZZw2bDCv3zPUMocU3XAepEmWI2dKGe3tccihjpTPyx6pCZyE8Sh4biNl
qzZWkW6equJSQo/d/xiWR6JV4IbnvfYCpxbtM9rKwaQFCifo2njjfKu0peUVEoov
RHg8wrAhtlmH8DqahQYkyv34kuEg235zFUTMliIB6ds4ranmUdU0miPH8Ji/gQp7
JSDcyPokm6QpNm4WnSfOXEFi9ndV9Ox95JEt2eB0IMmK5UzWyGlszSLru+zR0AHg
AlQfiz7Tgu7nD4UhanqWM7CgmSSt1QDMghvUzdwwCrZJKHp4jzFaJ6yT5NathiA9
uGijK5BeddHLHuL4aPRt8y1ffrOYVIwg7Ost34TtMWO30wxmVyZ0YgMPqwlg9uUS
6gqJPEnFycKOHEN4EXOxi8Fo505fEYZ9YjcSUekEVYGm30iR8i1ZLOY50fUsNdI7
AQWI7lBJiHA3WKRRzKcuav6f9ZK+iGExb2yUd0bSsOVOlfg7UWPvDjkAX2XmHmGQ
axP2M9N3mn8CjolZoVxZv4MGWbE4n70WdDk5CuK2ZW2ZVYDMj0daL3TlNXd/H3SK
SJwTDZDH6TMIKGdQSmZI1mcxKSo5XYUogGqTjIuBXSycdGBsHeaBM+y7BvtvuHch
sm1wWwxdmFHLVjWcJ590V19bM+h9/p9PxjSWz7pL5pcBA2KGeSPV6H5QT8Pn8GQi
8kjBM4RT/XQvucVqpu2uDykOMru9VB6GnErbd79ZZJgcy3fRSYbuBDQ49V2ULj5Q
i8vE7u1emp1kE2bgSVIhqfwk2P25eGVnWevIyJdZeZDMXXHufHGsAtnwrcn9KEDp
sQiUxh7J6aKdZEnSwuM85R3li++DQNh4EGiPzEbP5QJ3Mc0EqhVj5aLFNJhHQ7LA
xix1BYrfcIR1+APSajyToEQCBuC/4gBLR7MtsRXAnQPgvwNdiqS+EkZmMLMuIEs8
+S6ECVA9o2k8RRb54uQg+3JwGBEdmpzAHym+Wx2PSoYAcUKjSMuWia8owNsr8dLt
/p6bAdu+K+slotLOCivc316X7hdssG6/n7upN6V0s4KJBNCfSwIPka60kMvHIlIa
DOszldHe8PMiycZmFjsR+mJoytumVR2fCuQOb/wN9v0amXFw1HPuNXop9bmpXoEO
tLG5wM0UCx5Xy9tFauZa26qqPMnk9m96SuDPM1C9XigQUzw58kWET+IKvO98YVVy
1JBh9JK+U57xslPS3FBjQ5B3khQNLukAMi2gdtupzeuATDB/LbqVQHv+UzTpRbEw
uBPBbQwsrRV1yN6X8hLkkdgnieEZIreojsEeTbnUxyN8lF0E+4aaJjeVXWAn/sWG
HUIaku6VruTgNUQPyLNrT7JAgEMu434L93qmJSJBS3jTd68Dqs/QApsiRaymsBzg
MGL+jahzv5bc0nEddE+vbRoQxA64WETimRdnWV3HPtVfLw5AIPu466CPu9Ovf7OB
76PpRRtXWgStWRIpzx3OAZPlFZVgsNRl3OqLy0ymdcuIoX+IZtqR9Hn4/a7tCE0z
b43V3vTfvMNlTn74YgqOO7PVlcZIOqkUQuVaUHS593YuGsCS5m43FQ6Bfm54A+Ur
1Mg1aFkzSCbJvnrk89/b3zZseNuDrUL+kWJR1BLWAjD9J4zJGprXwtMiekSGB9+3
6uz1py2gr803pTK9usG0n61MYxOD6tsI8jPqgR+yO1V7syPoNu/MxTwnPL0N6vNU
DAtn+xkAFG8puqh4vxuFq8deU8ukRLQpqRBstwSrT5ZTuMQUbgXSlZrte/rO2OLc
DT4FCFDzyyWV5P7aRrqz4yJaYsRKTmsTINLLdlBl0ak1iUIGJspRwUvHvntikuff
rGPtckaYgO3k14NoVomo9QjX8M6wfxn9zOgab78V1NUb9WR27BqeCM9DwYbbd+we
VOxDc9PKiESgoZNkyfc/VY6G7Sjg7wi2gXDCdn/Oa62NniZjj1bY/1OS5u+2Z9Na
tlovY26K3DNVW0tPkZSSF8y92WIDW2CbaOC1JpmjNXvYQDrCYs/bwr3bLSU45r4S
i2td2lgu8M+giIyd12lZRfGn4+5SOJnEQonGF6KMT/yWJLJtzQnxyGvcpp1mp0kF
artBz+FS5UnNDoULnjJmFtRlmqJ3bK4+DrC8Qhf4SXwkNWCd2HngXRJ6vhtkqiTv
ITanNyFgY6nZR0sp0tPV0DqFz7cDtIXhO3zuHeVIBDGcDx81TEwfqCGS4F9f0VTy
e+MNfxVQsvEBNh0aUOP9ZvFR6n7t6oQcERVKEPddDU5J+z0TOaOpllN8JsAS+HtP
5LAOEvsnlQxbh4bJrEJ1+dUkHut2IsAVFt9dP9Uk4ys9UsRWuMfNHu4nNcGv2MWx
ViHL0JrUdiwr+vvXPpTjslSXKCB3S6g09qiDztzlFDAnpXewpspyD2r/PFr4gvOJ
zW2AoKV5WpYBsmq9KeNg9eF4Mwt6JiEeBx5kMI3hDCdLY4KtDIT/tdgzquz3+Kvm
j2QuTuKgLV9xYWS+MphbILwn4WbQbP+qIrNLGV6WBuNINcGPaGiFx6S5raoliQUr
ty/VCfH6ZroJIT+OMmGM4TvvCy4M2YSb4BBhOM44fAB1S8DVVu0gimi3KF+RmDb4
ivVIBgbcRLS61PWeIvtY4w==
`protect END_PROTECTED
