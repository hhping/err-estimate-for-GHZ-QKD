`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gTbfMpmYnYC8F5aDB6AvCNWMi0P+LWoBF70jsPaSFADU6/ZSDG5oFtl4/38Q9NOy
c8hpnV5SOHMxb0Ptyb677GQA4Vr2yq8eA7Ldbo9uLs3gxnt3wRB0Ajmseysr5f0l
oT8TIInyS37IK6eiPxHowhxqAJacmnSx6giChJ06Msea9TWy1iugWqEvySGZ85iN
/rfSXR/QwJ3XIlpHgXNXXdZAmOSROntPL6elDFQtfN+tYHN0f7FRPVCorKL696UG
gMTGbXW8cHqkXe6n3Xr8/zmXESjAwoDeTju+Y7G0Ay+qEyLQumYMvtHwkw9W9WSw
Xkmky6H8PKSUprL5GPYsfH8cfSVqqxbjBV3th4WnC2gwbbTxOXQ+B2yZAytUKi+0
PwlChsyo91bIerGBi53xi7OddOqoM7BuP1KyMYQLFIdPQ7RorUI6Q7oOVEeBWXIe
M1bpa+V4OWyktyPjCt4qUtYQxb0Dy7Dsbx3/+JfDKBfETNL14itToJiVToJyAw5Y
OxCLu+7zlmdtfYs211Olt1oN8pKKU5VDKjD5WY5u1zGah+v5Y+UoMPHfvw7PlIdH
3ky0t/k4en+7IlmvqA7x0IJsPD1qdE4lAv8vU2nueF51D5Hb+/RY1j7pUFfEsFpQ
jgOwvoFw3GLf1cjveeOBCP+Fmt33aMX0055+KfNTCunTnr4Uw57mbmUTIzhBtCbn
TDDE6ETK3qTuWsTXZ3NhlaEnxYogE8rbQZAkbbqwvgXZ2W2EOFUk63ul4k4vh24w
LvRELcukfbeuU8DqyCruPmZW8lt6ACJNn//qV4HtYcRf76Jqx6L1XqTyaKpv4BlJ
wScJT8CHMhkLqLEdB5vzAajnj8eHVIMLY6u1ERQlo2HZKIIHX9j8D4F5TNx+bBMV
MKb8p8pwSPz9k8E7odWlWULLVdhnm7BI6Yfg1cBE2CGsn4cSgXIAbUuwW3JwpwlS
2n/cSXI/0SMKl9MasCugzOppE33vDFDf2oCebBaddfYgyd21VwRHnhPUa881nqLf
k4ugWkiuR2jcobxDGQ/F3aoVPGQUmpSJ7GIvSAsT+3cS09nyymLIAZHXQjQhOpu5
5gwm9gmSWxqZda5z5X0qcHmSziJkwSaENCTVedwJbvWXT/6QpFLqBr1mm3/OU/FX
NQz1SdAYi2zKszEGvyAHQQTyCkBDVTH8LAkzKh6KLsak2h7I5Sj5ciWuhtHAAe0C
AWTanV7dStQwJLSaQN/Kq8H2/PQwliYpj3Jjkb8Ymhve8YhnjadoJjKwcR5FWn/k
7lP+jybuPI/yMcgph5Yo5We1rRiumxZt7H3SfNj2/MdVkVztk+T5g7e6/PIDTIM+
vI13vAiwDx+msBV+L5TI/YRaNgqn/wG6TG5Cs2v4Ad2O8o4ERtUBLxGild49oANC
VvN10qyn63sqA6qDxxcKBNuJ8K70CBJLgf4zn02KzLlfohUmGxHvWEDyCHkznpIQ
saOp90TK4Ilqe4IkLnYJEA==
`protect END_PROTECTED
