`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y1xyNYp7wpzp23Ru6O7RCwhjFkZ8QJgcjrfl2AHqj16+ER7Tv0g5M9l94fYRWG84
jF929b1a+9q+7r2xV7GM0/BoiqesC1fAmONtUX+eIJA+GYoxfcNwiwGCA8uBf4gP
gI4C85Ev3/5V105e7uB3Not5zLB5Z9YEbJS/iymSPhtitn66lDIf+g4pCsrHy2o1
NgcpYcQq3ZG7BejXiPhOFm5M5xnRT9dUQpLqohz7dlpURr+JpOFbz9tPkVsrE34r
JwsECwB7sxtVEWff3GL59krj4zqei+Z6+G/ljtXJFReg1OB5RCvpxrBvTlBbmAVe
eOYz6fEhB5/vRh0+PhCzJQ5niYV7eIsFz3VMBUWsh6sFV5UHSUx5ULKHTiuakuO+
Udby3dEdX/zxPiwVgdrYs0O4zRwn1B1IESAe+Hr/8fa//4wFpFFsohweSnfAlvcb
AIFTmFRw9icOCbJ8ClPaFbN4pNT0UHELSQOG4YOe7A0JKASY4JW+/g+N7jguyRSY
bmzMTyjaBIZ/n7ywHBfKuA3oFwekiFFr4eX8GlQaJgAHmQleZOZ/eTQ/pFAokFaY
ZLMojBQhfE5l4d/uTZLjlrzYD9QG9kunPVldXoYxscPlTmBpkNENIMPGRroIl5CV
AV485HBlaZf6BCaY1ruvDKGB0ty8906Zira7GOegB3w=
`protect END_PROTECTED
