`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KV2e3zVfF+C5kIriyHOkxAHT1Y/GMoGJJ2uky3Zq4AZJ4NTWI8ja8RfNaiYQB0f3
J4y2FlLgrFw/gW1stHVT3GRkoeBUoR0UHL8h4QDpC70/oo6yZ4JMcjuQFDMGr5SM
eertR/y8m3PA48p6Stz+hpuCP/ZKGlt6ZMl0LAXsMYp8TcQSXxWKnDEOVARgkSon
PSEwFMM+z7Ygdefrhywec7/xVjQn2oBuIDogXuIbzC7KL89vXQEUrY+xFw0bAgNH
muboWGleee/GdfS4I01mS689CSBOBK4hxu2Zco8ObbPab5HwsH4KdJJ38xZ1gofc
5qX7iIHpdI2Y8mlUIGkpAV6WD4C8kZrhuhyCZKCVyL6rni8IHp+zV1Sk13csVMOk
RCAnYEp/bv7DCM/LaH9teWT/jALUq8VYD5V1kDiXGCGeFKggf1t7qIvlTDQvI4bm
pczTIc1orK5SHIXBSpKP1QEEAal6whJWtR0ZWpNimNk=
`protect END_PROTECTED
