`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5u5c3zS93Hae4QsQ6pOFcrFzDhqBSAcGo+Bx8NpyCcjI8u1RxrYHADfEkjM6GCuh
B6/HhBvVL9B1Y8zXASnWzh+pfmPG6EZADcdSYfCePkIkCJ9ZRL3hIGk3F8LCFBo1
sqR7IbtWGcXwesBpWFMBNa1cBMgmBqY4d/+hw4aJRK6tvioNtogKenLSpQOFAGIi
VVa6eEg3zzsLAhUD6clJXwMJoP1fwDRJB+mo14JXjmEaf01Y+IIp3JQPWxkUCx5D
jfxH+Z8ABhQNGTw7qMEwd6ncIXlmVMJ4aZk69ExzQUHsvU7btF7vFN2vnEp8vMyb
xR6bZFg2vv/kVIAMqUXB25JUaBekfyk0JlR9WM+0zUkilUb9FqmGMv13+EWTqV2n
kLSP19By3ITNlSNpJca//w==
`protect END_PROTECTED
