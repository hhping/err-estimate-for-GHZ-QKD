`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IqZeDxi04CQyZyUXA0Dh4PQ8AFMkgYZt/c07XPVtXboKym4FPtFEIltWdtKJTWv
ABvCvlxn+hoW3iJPOqMpmWVI5xtwxcSQkOzVryCE0PGymDjgP84Mbc76JdUBHqU6
vwmOm57AqBuxh1Yyap/k80ecLe+GYyEfXbltTmNV8YfWhfkD8zFinxwKqHY/F9ye
6+JF0984eBlm+R/PLVVj4rvwn2YOfiOofWhSGvOfHC2TiIwnp6RuEbNTsCUHNs7k
b8GekkSF8XHB3kx/AnpX1zRvd0FgBDrE/bOOuCE3/Tfgs7lRB60Aw4sXG1pLBVd3
0O8OAbGVqLpZWmaIASQ2Z9QxKYus234sZ/avi7AaE8NvyKL6LNJcGJtIQafSyY41
oZqBt/aleCkl0iN0VmjkXlXsRqdgjCIWYsj0glhvYKtvaffap/Jpwp2Jk5qIC/IO
WflsoLy4RPJxpqq6yBnzc/cd/SylyPnkXEEdRnO3rorm/wWi2vlJcgHuu9anpZW1
N/62JSYq2vp6BllIl7wAxQSX5Dmhl7UmDO9odCWYWfchn3AsJFA9gBRPdpxrY/X6
wkU80SjtN9pZNNrmucCLnM7/QWmCcdIV++UA97cMNYlMsxch8b3Qzc6NZ27/5JA6
FhD62xqAoFQnJo/o+km/N1X4VfM74LTucfZc6nPHd7CPNWSwlUhBs9l6C8asVaDw
c+yMhyjQjDnc27eWcI13fq69U8LnIvO6WkAjGCo1zkVjhpulcWfogIRKa6asDvs2
yx8hauyOcVPe03bhGVbgfGITbxaAmUjRzFjVO0RY/bU4yifSqHnGB6fbo+y/Lcgg
rqStTL4Cs9Wz2rYONoOPNQhmI0haPwyevsM47VPugsevneQltvGoP+0TEwAkyAB0
yiVMJrKBWnbLQBLGjPxdkJYIvrRm/S28Bc23Tn+anzI9QDRMlOFc/m9MsC4tfLIm
iUKjl+RFr+ci0T3MSoxIs6jbXZu9QhR5n0EPeytp1NVuO6JDnkLe0QIFoXkSGc7I
ybHmRpGyA/+R8tIWquHM68yXhZngHLffUn4q/4PWUURXHP/bg2URBosmZ5XAeVf0
C59Cc5VqQjYVv6X3WxKjY9WdyPIAmC77UD9T0cLbVIPF3Txono0vRygkDu4ZtpEb
pAUxaSV9snINuwujDNYVJU4de61RGnRqL2ve1rkSbpH1K0Sl6tNe41IbzpgkWPy5
ksiFYzUbqJzWKI+hJsMNDexwNCIAWLpNw+IU8oCqTNDYP8d+YsPINtJqTMaQasQ4
5tK6Ru6BAPxG/sSzrfsg+0aj/ZK9wg5deqbOmWCeZXt0TA2fhTOhs8RC2BjOwCIi
iueDJvq+CTuBXcZ4MEpg9CfaZgV34TXTDNOhfKGv1pZJsSeoRcb3tevzW6C8K90C
0JRSNUWj6tNSSiOVHfw1asg1aRJWhvm2kjcPe2j1W9orDc9I0XtnShhK9Dqe6GjF
RBWEe/2UAuCzk1XSOIKOWHpcgl9PVk3VHrokcMtn8grmD/IswDIvrfmzltFZUHH8
kSCiWx8mWe0Vl73hGRWgd+79e3m3vXGeug00dHCUJkFLzp3LlijLT/xvHsCixgv2
yC4wfSxNu2p2NNcaQ/VEV8gslnAcs90fcgsBM+FC7gP6psMLZMx3yqvfT7Qrzl+L
qHtGiMeovCF3Zi1gOiPb/GlI3byoxTUDOGESvG3eQEMQmGDIF1EGypunHOoXwHQo
cA44+BXnUBvX08giSdJyC8yKwcX5oAtDAGUqJC8DSPsCdz9d+9AimZ3Mb5Yvq5i8
bonsuI1IMojNNdck39lmv6Wn/6fHvE1XOI/Bh+IheycIbfabnB4tDfQHEfc0wvuH
3lfoQOBJ5iT0SIl8TgVpXA==
`protect END_PROTECTED
