`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/ljhj/nWAx2+jL2CG4hU42Wt0M5eSttV2DjcZAH9p4YbAs2RO2v9bKcq8JbzUUJ
1sWvTxpQTFVxNlxSd35ExjS/NDX/qE0MzcA1xtRK6ors7HJ+sNY5PWa5EajuKjbr
68ynH0wAONNM+b9Fj57e9V3FDlq+Qoq6c8cTAw22+BnxfVt8zyhfou2c5yky+Xay
1M1KbN1trlHbsEKk9Dicd6aBNK/JFa+DVIAhhJXxteGzb4riliBIO5xP9LL03gZT
/TCpVQSNCzwku+dVGT+8Fvzky/TjOBfVhHN5KENYsm8Q8HSv7p0VLJljg/f0gj8s
BcptazlWHB//iNfqmXmv+GpZtCz9rw9X33yDE7ejZKhk6JX+h61W2jIpRQDQzufo
lW1q/KlhHy6WvdtKeGoM1nBStrihyTHCJwdRUcDuK+sZkakRNVSv2Or7nGXXWOho
JPpCC6nn0WXqsqwpd+VtXun3m1MlTnGVsU+PjEyST7DqlNAe5AtelkvzaBOGdPqH
2i91/L0GWmIKIf0dBrHsMoDEXspq2mTPO+s6hDcHNuq0evcSFwS1+yJBPQL06bw0
ExPT3MWhQZUiveo4Qb1F7l0NDVV6N+OOOdEO3ozN5alGUox2Xhc74Lhw+K4wLA0T
yx+R74ALlyvyPQB+n3PV0Wx/3kMdtlGK4c+hDkPvIqwzkw3NHkTD62Fgfs8X59o6
FSkfmYt4M+gkcWU1y+BZhhKU/zyGzsypnFG+o0aXDFHRW3HpghmKtPp34eiWj5bh
N0TcCngjMEq1g7BHCPn4kkLcmHdOTYz99Qas6pv9JT69s9WwBvAeV9/XqDMFSORn
5UcxGel7gMdKQ2Y/gWaKCNV2+8L+JJdeyKaKOOKZBEWFSq3tBzYxKTf5u3dfz5tz
cUuEQAFpw3YkhNbWnGBR1jTckU5/mHkkXVE7g27tRnPOljwQP2sfYdXqY4+ZnaRY
t59ltdC/L7xZqCVn9L8HYDH9ebT/CBCmpuV8KPT8Uhu7HAe4oCQc8lCW0dtaRG6z
vaguoZY4lDi17qFiW5t5lZD2mm1PVWUma3+sfYG4Q1aFuLAoRDiVWylz3K/NVgA6
qTOfWZs4W3ASAxxqPlZg7Vj9DWfB26wL8akELpp53VfB2GnNNwPGq/Rlk01jpt7i
aTU4d6HJ8BhJXozlnc2HmJLe8erWstM9KFjUkIUhmW3CSfckrlLiT+6vLi4gThgz
0//65J7Xsu1AF8sF2cTeveOG89r6kfGgvOSlvfJRhTYEi5RXZJkJcJ6p+ZziWiDb
x4Jo35wXTx2eSj3e7l4KzUbT2i2ZasauPDBVwfu7G17PKffaLFjvCmnWz0C4cWST
q/qRxi+VB5iTaMAxWBpxTBEW6K6atpSxprXpdeSpVnJ46D5VMI9p4jTxv/czyAqR
CUS1GUffjcf9N8ogpmYGnByT8mdVuK9VyUgYA0LTi9PsaVQFahjRbLgC4H12fPSj
`protect END_PROTECTED
