`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XdznUmBRdlPLP7W5zPWVvzuwvDgRHHvuo2P/hJ8eDIeSyXKX/HsxaQp0eDpCH5xT
pfHuv0w25B4OTZZKWzidx+GcsSfKTwvXWpL9PJqE1TtCLX9U+qZC1KKUJo3cGhF5
a5ryfBx4w3jaOadHJ72lgHNf16p+kJ61CYFV2uQMgj3nztLwXyErFXte8L5G5jGF
GeSPnY7wKmw75mGPXdqEBkXvTPH8msJ7iOr3ys3DVY0v7NkYflrNCfg+R81aju67
9NK3giuasj0mwuYKRgkZIITSFlgm/kLEsyw01ZLQGL+cRYd+a872Z0mI5c/qg6g4
RMd5vUseaoicqKQgxGrxImDwg599hCmX93lWMz2vKbUDgcZ0hJwYbpxFmgGUmcpz
xCYva4sBwyJHao1484KA0DY5cFnVAXQLn9SbJNJmIMoEspz/XzAM3/uX93fuCtgD
//+PaX3owQapa2PlTZqZ8UbB/9btbJw+rWRc5bxfHoAy35k4MfZVlX1nk/VhkEl0
bM74TROZYXxBpj7GXtAKNdYXQ85MZK6Kmg01ytZk52L78V8WV8GKQjedVtZBzKd1
MRBcoAB66LOUhqf6WsIGbP/wHObrIZbzQAvNvGeNG1NHLx7sCAXVKlvxnim9BWQ5
Uhr/11xyTpyLYQTeDE3cQT/8XsvREO8G8axsoUAoxyzMKIfp33eEfq4jQjmbNiKk
0H2vz0Vqs0+ZLkR9Kj78P9zH6fOPCVA7lGl5/tULZGnvU5hrFfn4/0G+B47T1EPG
VGcIGXz6NB1yLXLUXVArIDyPc/YgjuU3df9eLHLijtF/2bkqtOSPERw5Yi0nG3Z0
HsnMx1a0Kz17DRweVD/Ty/Ke2TtfaB1sOjqnOvPmWojddKTB8HwJULq5wEKESdft
FdcVIr2BTmE80tkk+rWRATNuR22PaDBQD+8YVB2tpwEQGM77HKnaoZOsgqsptjl/
RGLmZuS3/66QcDGk5V04WpTPdOYzF3N7jJJNhefWgv+SuIHro8Wg+bAOctVobEvV
eyLteFXboOaUZUno7xn+d0Pq951MRt17GnSe1I/4Elm56QaWvKVM4Qt/9duxTFSp
RNCxHtTJKx4gpjfdDiQ+HzJY+khSM/FqiAqFxfOJ6h6FHz5qKJ+2kO57FleOHk35
gPi14S9hIWJ8vHplWxoTehs4obWD+uAaTm/RPhTzM79T7kTc2olc8bJdRLDuwBLn
QRzJc1otwBWPfY+Cu7CNd1+TT1VdJ1Dgj1j6niriLs+S6OgsSWXgWg7J+7f0CDiA
1TshjCW7Tq+smpUz3A22tgDAWamINU4ZVTHpjiaqFbaXj1+qV1xxlNXnRUe87jox
RwDq9TucKcRqGFlDN1BAP8rw3Wi9E8evbdHsm/fIXXHYJWJyt2WnLL0borxS4pFM
VGgCBdnnNS1NRYit5rV3ESLZRvGtJRgllcK+VelczzT9Q/0z9/whZJb/Qg5pw+lZ
maN61aJBqf6Hyys8ryh/piu0ANkglRGwpljCJJzzG5iNdkhXYBNoFb0+icu3sBL+
vkGZ8ss+cWyjDDpBBBfRIrdaDAkiYmIYEXtOz7jXjCk7G1itLrZe3mOzkzwBQ+In
ZE7/BVeVJA1PGtRKARXW884Olz1ClnVYsP+4Cfj9ZipERPqrzGtS73uYiW4Bppom
5fQSxFlQPBQqhrQNerNpcNGjErmiso36fd7vUzINzWExzqfAb2yiRrcvpdlRCaS3
2gCwGIaMpfgc3eqK+rjwkzZFaylcAp83r9bhBryxkh8DFtme3zqSBwkCWVzjV8bO
3qYyvVGh5oawsQXRe+xSeZ6n3U580R9AZawWC/lz5ZYozWJ1aN4XbMecxBfReZrt
qN9fgHKNOrJVjMRP2e1auF1NCG7NuecZfIPv05qpYICdnGARIMdN+dPVN8IM11J9
Ob8eeeva29+5xC2BF2DrZzaxOmtcPhXbeKruST//MiWwfUpOW6vGDgyWnN9cvFLB
jmOkGKs+uAshesS75xH/Sf3VWEoYR/US2c49OHqqfwIDej3J8qZL9WH8y0eiO2xA
A45jNm7ff0Vg4QrQK7jGmrgYXLuzQSsI3QOn13tRVFJnQTB9fgoCGGvGJBM8yiDb
l2lr/+Gbc58HWmBUUeCxZnkwOW8BNhPGFUg6ya1YMHR4gYLSvcxjm34AbMT6XUWF
7Tven+SgkAFbHys3w7REeKiqRvzn0D1ClsZ95QWe8+vUaKfF+VRM52bclS4qZpOz
+N7BBxID0bie6YWt/QW20lwiz8Qi6155Cejyru2l2MDWC4kNAgrv3SWBad6Eivsd
LiGyl0HH601iH6bQbOF+zij44t1PEK/OGK+NgLZJiWXF4FgEnZDs9CbG+upFABJ0
6OS8sTSZFw7sasmDZWjDiOD87abfcRJrXUTO6JJUOBUN92LWnT5HcDIIB/7ngUJD
V3cJcKOPyZFw5i0CDNVCnsg4ss5B1YqAilwpws3s492Nq37ThFd91b7cyDhIRP72
t8nXEzvln/4VYXD6ybUKSZgf0BJ+i6Fo/KCYf/ifrY/Sy/jcZ5I+3x2+5bIoe541
cptmjKE4b6hROshHlNHIa/+UzGdPcEQOkQNU7/j2mnBgYmlsGXmldHA/Mjy0lfx7
GEUa/fcstufrZxbzy6uFvOHM0HccMOp2lJovflemMO2kawQVZzn2lpBEP2wGXbgp
UsjC8VHtHUFcheueUNK0mmUDp9ZNhxMVdfIsaj9efa0tW6K2uvLdd1Fm6TLxXTSK
C0q4MW1yVDCALuAlTEfdPNQqqds4wLxkFSBINDYhqg+C96BKQ46uyctwJSKCEmFT
Pf8jKtg/OhvNYCh+RLXZoZCwLV/LC3W23kJ1CjnpjvdFRAKdH3eIIZQwmzs1ydYv
se4hSFz0Y/CnQYXVrkxNEGMWRlmYakMJpOZDDzBXon1fXCSTSZ6vI9unWBW1TQ7K
/B+ptVDDdCQ+JwtWTjaQPAp63hVgHf7hXbVa58FhgEYobIedJPkXSqhqiM8+B/ZR
jeD7iDuUv/1+i9oHcY3sXyWpndVEKux7AN6QejMLz4aV0ggUgi5bmu1qyhF9r4s8
4lcFS2VB5gyg5onvrn6arC/99g02QUzSiPW9U3Xz4bu1Q0ThXiF0P8h4UxSnzWn/
w8GbFFNp2zWmmKdQB7h8zCOIMFv6tv6G72hqIxKbQVUkkCtdvUykJ2MZdFbRsDUY
0iwOpTVo5ft8d/nxUlli50jCJ6odAnTsEXg68bnOMirB2RTlLfXwiqzUkjSrOy+G
OL1C5dFXKUuULgNy4Ta2iJBx3YMAfGPu9+konW9McivHI7dE2lp6HBzlJ1irrRVG
OKCoZJUAKxu73lr2G0v3KPhIjFV79yEV7Ap9qldS+ZNBOVepkLBG8/IVgZpe1uWX
a65DJPNJTZiAVXX+leBUK7EoiJ+WWZSD3299scQzVim9jOxYYMrHTVhCY0YMTSdO
EkAoBSOzqHrNofjlWd5GdsXj2Nq3oHWXaSdgQd5JI998LpYPFfBfVDFEvyg69FOu
XfYtctY7CoayWawq/R5P8nW3pH1ErbLOZ0B4EU2iYrCRL4XBOlXnkgaVMl1Csvhk
SMgtxTEcQw1s6p/RbZFolfW7D/QpYf2YYanL3BQaBDqKQ1yS1IvTGixO/duaDGS0
anpw98BOuiq8wfwpfdxRVe1fJB+rU8/UQaSuqm3Cl88YTWuhy/8Bx1w+PpBQtx1Y
3t5xQX1ZLlsuFqQigV+kRX5QC427+vT3UFIGoAYcezCU6TH4WPB7DuMmuz2sSHP2
JfnOYqaKp84hsSS1dxpYwaXh4gaDPXEI+zGiH9/Sd3UPWScreHCIl7WZ7yRYOQZU
qAuNmqGR67ZywEiseCBz3WrCC49Mlej0gw30PACGiyHb6pQ55KaNAbsJm000Vs/Y
KVqV/OXh/qMjZCK+ZcLXUiZKWBlss8cxd0dTghewFqifnUUh2Kn3Zk1JUKRxBauz
E0jHqrMluvq3LqcrvSkG40lIvWnNokHzG9VpJsisiTcT3C1/RGWZ97CRcklwotf3
X81PuXee8TR74VnzJCnTQUd4xmetdBpSpn5deTfIfwa3R2eIUEt6dcaG9MmSaNyh
vUCgH//3EamT9HcWi9msOw3bmeDyMtkDKJhA/+a0Sr8p1qAxcnYwv1Ab+4zPGzsp
T8eqzV2jbQ6AR/7dI7PvdxgrT8Jm9mDU9VYIBWu/QwsArKx5/mnoxoY5sIFd3QK9
sknQfUe4NZEGbTDPjNWEZqHS/AN28DrsEviRR70Ik4+07LbtdAf+pqMXNMqsZvzJ
ewTtjAE/6XwEeuCbliASN/uYDbSJqIc7DKpZY2xIK/44oHPKKxlM1rK1FDzGm0zS
K9QGbRhzAYqkRim8AWzeM6U5FjxcaI1JOvkm3CG3FGgQjwq5a+2DmqWhGvPjz259
cl3Q/Ae1UYKc+pLPCSwxEJ+dkiDyaKYiDQSqxWWMLPB6Hqwf0wovfwaYJTBiEklW
Zo3ay3I02f04DfLr1D6rvNWLQRQtzrfksHvjNf1wQipzr+wbc/XbzKmvRyM065gq
GE7QUD4VMiJyboC4ZC48WsOfG1tIpVG8SrqmoWJHQ340K++mY3SBB9LcOp22YSN9
TrLwfUg8vpYlfrHGflLVmxZ87YIjgN8V6dfxYzZ3pn2iXtaEVnkQ+zdSIAv4gw2C
UmbZRrSh7hNFKg0NE/gGBRagEfe3HaV99xBjlTpzy8mmXaQu1Jt8OtBfNKDTZ4y7
rjU7qS7IkmAsUaworMcgAm0h6Tt3gbclGzELXrRWbU8m6KSN+TTvdJPMp/VfJ/1w
M35rtmFis3SicWX4V8k8WbDQ7sScokSDILIeNg+U+snT8L48SSPpKS9rjfOBAylz
VLHWZTQuKdeCgK5u74JZkuzs0nOio97faRv3mReFff3M4R0EdCjestGvq0HQuCZm
ZXTJDM7yS1jr16Li1iu+Y+w1IlgMh4gCx2RQ1lshx41RcQR/RZyuRRC7gvWxAD6Y
XmNIXMNf7hFHpdKhD4mHN4+ZvNgEWDs3pEsqztJI+zmhKJTU/3+t5r65HOz784Hq
9YbDyMD/u63v7rY7RN7C8gbuZhreACoqTM1MM9nzWG73/mOAdsd74fFtymiti3tT
PSgrx00Tm77czewnzRaO4DVtXwcY6KTdxsz9dkhWdKuWo201WSuQfwtKEKGPXtdR
ZyGDr2dg2mdS+RNpStLPGMuOBWXZu+NuewBSNJmqdDYVziA27Vls4Q4N8AlEO/MC
PRHjv0yXVdoO8bPoMMZRpvWh6plOYLDM5ZB6l4vEAJ4xHfDaj5ovWbutVgCRh/us
CjN4s+vF+1/1pxj2ClygBvJeO6CrQLeRl0fUrjl6lLpdn6wfAWkqywFQaH7LHP+1
Q65MwvEYtBYAqFXcgpC4jssqlxUBdkuTQkUkgYtPUgMrju9gNx2ecpIkU9FjiyF0
LaXuizvLTep4Zvzf1s2xGjz6Wz9XMf6hJ+T7hmIUq79mOPsOaMAyPNTtjox5UTXh
FnC1srw1VAC4VTHsM14YCMDz8NkS+Q3QuN3qf0fIrHChlRIU5IInOJRbxPajaBMm
HjC94LzZ0qNlDcr8g8mccygKpjHR/M9ccJ6SKkqwfo0ns+V4jiCrLwKAKN9eMYhe
VELYhqahEe8GqDbFW4/jrzHLyrZkRu+3caY+ArIoTV9hkYZx6z1xd5UNjf8NXqhS
IIC4kRKxUIwEl3nr9on/D/BydRb2VuO2xZqC3WL7d5Ebur6kUTdut7EfSgfPnvoA
ZKtN+S421zJXD2nwXTfb354a//0TK/lJVRkBZwTkQj9NMdC+xgtMV05jzUOvyCBP
60s67e5tHxP77MFvJ1kUE5kO6XgOe14xRe1zJ3h+dzAfo+6Zrp5OTg3kG9dqgZfj
xO2DI1bzB0qQCw4K3Nbry2bHR5J5dVHkmEtetEKIiVdWcTjFQgNQsphY20VwZwBI
T5LsWAZpFYR/fzcSH86E8eNQbIeB6lCEsYe/LU92KnD4UTZfVKVskraXUAg98KsF
fdDh33I9AslfI+SMQ467gr5eHFZ9wYu8tPdvk8bBUsyzmfK7PM900gWEDhUziEMI
UoGePPiMGxG10eWMgVX9r2JZqGNI7T8eS0ZE5EgugGxxB9KlKiJrUAiPr4PvdsKk
P+Du9n9swMkUq6fMD9B36ZwyE+VxgROjxopOtpl7m6Xw4EQtMb9DeplBbf+aoKx6
CP0+2ycx8OGatDF3Q6LHUXlwphiIZHQ3hWZwfbwlzACYeiQum2/2cW3Nrm7zFfPD
mJglA6i+QxCkbJ2JA9b+hqz9UPRzqLkwkYS3Z66DldRHGReeWhopyNdsZZ+jcMp6
luh7PvajyX1gfPThkhSjE9eaNJGuoQq7qOIYcKbX5xWdOXDgAw8vI4+bs1mtmgny
av5rKCnO29i3rVXOShYRiblmE4D27ECFXv3iPpQUYxQGfymwQJqJaF1lD6MvxfYO
VCcc7+uvrtcmJ1He+cbzM/b40WZ2OLhaCf6tO3HVbE4/rDJ44DwTsEmcq8dKdd4H
z3ud5A+xVvrhgGe7DLfniL3SoBS4jh08/3yjxf7AVy8ROwtzd7On8bSA0xUTSh84
CBVed6INHC/vub9MtA2KDF5ZE7lZtul4OEb7iqg60ezXUid2+ZH8VQI2qa/hZvPK
uD0NwZect/UO77k6f1Y1ihsEy8vqU+LrcVpqkvwtRJ9HA/pu8Ed8zrx+y+1o3Z+o
nV2X0otj518755xxKb0oXP0VkDgOz2YOT10QtlaeKIEJONGslQZaJm9QqF0DAuhx
m7GbSX7ZjzD/ZrTf0zzVxtAmtfS4q8VveCqhtfz3gEU=
`protect END_PROTECTED
