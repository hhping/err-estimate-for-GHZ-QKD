`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Th9sUxS6z/1Ea3cGeY0EgQdL+X8fOi/700yIw0/ZxKGk8SX//Zh5Mm9x3t7d6DKJ
1AAgJ4Vahf9n9TFAoU3QvA5HaSS//pBvXiWsg3Sc6gV9wEJjwnvYFaDXrJFA3+xw
n5R99rkOGrv5IL01/6aPi2JXpyJH9iYJwXhcIlWrl3wAqzQz7ZtU4uP5sgsWGl8c
/uVk8Cp0pYJG7nSt3gBJ3wtdqtc2Ltmw38PavNZAnq6zu74MVJULhMCCMCjcbMyT
EwvIW3L8TEu9QnLWYlzF3TmJ6EnVz/3vuyAo/38vptiTy8ObTEMKh8H1fJh0FeIn
JpH+EL8GWVffrUiHi6GAIqSwiHqwEKPUBg9a62tGQh8LxYS0/7lUxnjLcWYBjAU+
vzW/ReptuVDyPJQnW0W373ENhtDTa1OrMKlz1wN4o80MnaNjcmLcFqKe1xDfrXQQ
17AB5ll7S5x1edw5Rf4z+nWsO4w3yLKCHxHl21Y2L0ljsMA01HpKLUgkzWzMhHQz
gt2J+9lm/Y6ahutxYv8KfdXLKcK+fbT5JvIa3+1fBKNXexmztPXmigpLFA2+Ffa0
rjzvwTpU3pU4GPQ5r7LrKFwAFIYJcL/gOw8pRpn429pc8/MsENvFwnMz86RaNgCC
keyOBNlnh0sVhYniyG5UEkrYDFXuQxRPUY8SoMjgMi3FD/MZNyOkubNQDPF10/3O
g/SAUGb2kpUnlJJZeS1rInC9uV447sopLLirLVRmOa4tpMlVZSED8kCoCOtdhOAa
yWXSD6uU37nPM/pilMguijtWKG9oTUgXgcDBnYiuUd0aT2ZRz5GdqxeiNfMNgrk5
4SwTpFACSy1LzuYxw0dIniDAV9pwVoKakvNIFB4vWsPt7qWCv0hp1ExAHi0NOA6X
US/ZGdXPNGtnRrWsuRDDkearTjj/KgHEQajpV2dnq8AdBuZIdyKHkKq37EtrfGqj
vPYMHMp55FPCUpI/G8BeaqAG5qnU6VhmdBjzMjKMBqj90imtXzeTVKifli1aT/KJ
3WCi7atDNjyxl8OFHTgOjqDGI7KvR8hQP22cT3/bm6EZfDGxetnqpUMVRwmAP8Mv
zQ5+QRLWYSzKmUO0FJMUuEm4vOntx+aTOWFpziCcxZhOkq0jdRQnI3i2IbtOLofP
QYuVu9b8eMF6qYapnyymzYq8ClrWgXHonCi7zPN+iZRolyD/xV5ghmX7qsnlWGD7
+8URuncHq0lR28Mj0pPf84Isvw1pN6h5BmRLIds6RcnKsEKCPEsSW5+XwuSwLBhk
65VbAihzohfj4odsVAiNWoosg/YU/Vni/MTdS8I0uibmK/i6WSRHhxJrkS4n5cto
ht6ax55GMUah3lOPp8fq36Z/FJAGU03QyIJ+LLt1tVm2cnqx1TnTp/2ZfGnzD9Zm
FuQks/5JvTMpCOglX9A7WCihNy39NFa24Ztl1KSKppHL7SOjhQ2tsosdPYkAQbo0
NtriFISsQrz4B6ZBMZocbMF12lkYQRxn4UOneD2R7gzuhd23XMUEIOzYeOh26981
Mlq7y6LN8vgw6roRciMOSMSFSjKkj0EK0DP0Lrlhf2kceo2f1q/ZiumbkHVyBNx+
CJpQUuXvE8U/CZjK70qyL3ZGyOPXvTlZBLvVTYHny59nTdRspKrj2x4E6a2loYTh
c0BcwtaaqsLtVDjHPLNQ9CEk4uH2dkDb34O0dwYXwdtRS+PHhYuM4+Plzv4FvV25
jtzfWLMbChBNvgWtxhuo8FwOun6oQ/INlzroV2o7n8QkYmih6TlbwxTgtDTsydlZ
SsfR7Bkzjz0NhJe2dWGfdEs69ruCMNPWlM3cBiCA9vND5fsM+QX4rohQd9RJG4EQ
dHyBWuyFSwJqrVs/yi8i5+QvKmRxznX8X5K0v5WBKM6oegmEo7do+8uHe/giV9kI
GFZBBColGET8vFhENRKJ9yhbzpRTz6RswxS247USMG/uvBHjT+P5vLs7GT9cWroZ
nXtIoq9YwYC/+eKhTmhuAcfIsyzdgeTNiL9X3W3QfC74GB5o6rAszyTZzHLQByZK
XMCUJn685VrvhqM3i/ABihH+MRYTemlZGzoEzBpMvgg2gfR5xrqHNJHU+rP41a+s
poer6Q2ZP1gNXsRdYved73h4YVA/3ZC1ZgUhuCsH+qPDZBfVPRoLMM3z0woWObca
5HcjNneo65yp0GouJTHSmCXi/cLiUxB4saJ233+hHplxDj4NU67VYRkMwIEXIeU0
IdIQbUtAd43BtEYb4qedBKTXxKGxTZsHTD1I6JiGUumX0CaZaBErZiQbQfTIaXTg
1aDfDBpohAwgSpoV6mcCt/2QKmjZ03eYNtnEZx075wAzLu+yWBqE6V3+mOpWGPQx
IdLhB6qt8TJ5JRYpFGgD7RrIar3nAWZqXToY1p+PTHLC78cIBMAfaPvlGiSOVzOa
rbW3YUKhFQpHtzKHkK1PgIQY2LoF1Ex+Xr707x2VnPYxDUgGg1UCA5Plw3WRB1F+
zf01a9ZmHEKF2mqYiZAIBcsB6Yx3htV9Wn4IdWDygLAFHsMRE6MPdhnkVVaQ2fj4
z9tGnvx8KRtoHQwIG6KQxNIefan+jwY7dOPBtBSVjW7UXTaX1Ia5hR6m5il6Egvz
jsgtfdz4pRsXHG6rwtUDHaljg/D6xM34Lp/LmBeyLuPK3kLwVpr96oR1FDHwZdPM
FOLz1PRforp2Zs8zrICeC75Fbp224DAlsP200DxXHxJiIJPQzbPpHRkmNXfJCDdH
069MuwkAc6cIgtCH+Om7hIBYR+1ZE1An1S6w1QKZdfPdf0lGBu8QXUcLj3K4H1xY
utm9tWFNa/1mj0QJh2qL2/zjcaKYRSqGKi09f6zUB+6xl+ViMcFdEH7pDgVaObeq
tml0G5JbY3AxTpCGsRoN+3vW7T9jN/s8PHJbJCLRhzTNLeW/1J+6KACpCtrvzir/
tV9izzsx7pFAsivTclPCZ73lFdZz5JxP1B96vlUYwjro5loSxjxQFht9M2uGJ2Vz
wXobRNZCnJy8GRD4wdhHtKg9SCp3FoolQVCnYT9UtucBQBNbFtKQQbdUXT7CWZsG
0C/f7xVPSReaDXy5pyVHR/l5xVp2qH53xfx5h6RvbiNoi6mO2Io1iiS8An8fXti3
8RSLcCi2+rWZKx1m4eVl4QR1hXk/aJR+AKcCHJ2MbScLcREMfCXm9dKobHRDUY7u
Yiqe5i/b/kuoeQSKuovEb3MMvHWLyQpW4Z1hQ3+KbQUHusXXMY5GSB3ulcdBKFsN
NE9aDQC4kludeEpTshKNuFF1rJFCVOip6x68Z0GS30uYWoFYIXzfGFnSAf8kFHRt
Bmr/EOuttahLigxWi4ZPXE8m8ORhL9GAvDXCWKlBCUtCZNxW2fYCV1znxiJuynUk
zYeFAnV7FAOAZT9Ustg+LjOM5LrkFRrsJL6xuW16utg5SnzxAGFC0fREH4pxsb1K
1qXtRWSajtfvFq8acsJ+YQogz4fHRlQNOkuWngkBSx833ekutVHUDDUmwd9Uh6Ne
WwhvnyySuwKDC6JtI2FhbW53R9BxB/BTckAz5Ch65JkkplLjBqog60TAo7p3eZg9
zKVhVYHYiPu4FwWWqs1zlemSzRRz/X+FcS8JQwNuFTJYnz7GDQ1qksmfqPnwzwD7
0eT8SmVuncPjWVyIXE3QrkKme3teBPQ0yHXaslJQ7HXuQR4bL7cGf32mnqtP/vbO
WgzpdSsH2vNKEiKkOPwBkOL1fLqKNdysyHzXaP1vSeNAY6+sQnEcZIPVFSUcBSQq
7DoJqQS0Bxu8iI9Bkou4ou3Z6RzsKsMvCKLvvUZeE57T+2Kowrhsh4rE8mSWoH63
P9hrupoaRjEdzF5Z7+lCxiwDXaBxitw3P99xFCS51TLITGXuZnProlSFGn5N58n1
buiBnhyU/102aJFDmbqh297AWkssSq4dtMtSqHTN72rpXxt+YjtrT9dbH4LU/6z3
72qTtjwF9Fnhy21JKgqZKEVEnwZ+UtKvrd3yyRkJeeAKW1yeI0/5JuHm2WbRBWKF
PCuOs/CYJYxJIqvM4ohAcBlMGkiufMMugv4wULzZh9UERP2DY/c12GSGB0Z5Zq8B
3acDZLQMmj7wZ2zsfC7MGqZVW/sRLOuOdF430XULLyrYDfJgA6mmZru0DXy/gINR
j+9V03BHlbpeuTq5/UA1kWFOqdCUvhB6Va+I7j43kDkqcx5wXIbTzcty2kdpMf4H
QZMIaeiNy0gFg7qfhqwlBpP48tsyC9wCRmkhwS2N38PmuUkoCG70mXMO+kIcQHmH
ysuKoh5kspC6pNckH7ZPVOsQsUUVN6kV9jxlOs0Y3j4z9ciIo5w9cHvYJoUll/VN
tHhzzTEDR6jh1Oe/ALXC3vZ+WFTq7tRaXcmxWnAqlKfZgZ2Wk1r1l+wKczngz3rl
DcrNRsVo7WtGr03t1oOD96r/LWW/u37U+CbEtb9BrhkqhyGgbtgBW7DsmxwxIC6G
UjrNNwUm4UcKvXnFihSX484LG/tMcvVqd33fO7SdbIU0GEiVxa2F99U3VlteEBBt
M8eBHoqqBySugSVICKRZh9xSaE+IH+FIe75GDMZSIqMopMXIzYC/Rn4YbV3vnYDB
zK5nmJTwpzxrm8cOAmdkTjuKM0PZcXaZFs2njOdzZeoMN6VDkQe2SguFuwwtWfvB
oT/VEHc1Ytat0LFDYJfMC00RxlYy61lK7TLwEVHEOD253XjX7NkADIq13S2m+ADR
dR5UwhxshtXGpkPNsXuys+H3CgRqqvzg/FWT7EgRf/+HbO61bu32VJ/JkUcYyyD+
Z2roELIZXwANB8anpCjlMIELDF9J5ajuDAWut2lw+IVD1RiladH71hX/4odZh0Z0
0cFI/nubdnsz17CnZ17KoexW/v8SfhUvWgxl21RcIrP5b/cy31kihxYDCcEe7r1M
u8z+1gsObH8lpJ6dBggrO3UppQpjPKyF/On0lrYdMemBP03bAW4UkHIgN7RRwYsz
y3toZFilRE0/jiC69zott9wYOueBPdIFbRjlGgmicYalxlEFI5kzbEnn7oWkFD/R
y20uwnM4jjUANtytVT0FmEMUTdixwjmsyZW+G/3+1FU3G44Ochn/nzZC2wIFisRn
3c+w85pB5Y/MWTw2lIJPrIuZHdnWB2FxlmDVKCQW9SdCGU22Kl/+ZrURRd5Ql05F
fN+Fc2ZhBccjtJymwlMw0fDQObQFW4/Gfam6exhiyt4ZP7ritSJCEcLBfU/uOftW
raIcXD/4qQnYCzUAaZfGnvitQ5gK2YoQqnhhU5r6DyringQIK0vyKoHkpqEaQh3g
XqbBVUavuJfTUGx77TMJXBWhnBGGs3wg5q+75DpNynUSKQQxNSy5SF/xYJi1JRWa
tlrFvVc75JzUS65zNK/L1HhDFaMnpgvspzSkuW+i6LeAPhBa3seiPehVHgLQOTlq
VkuMeBox/iQa5A6mHh+Qybl+Nm6VjXphBSyy2q3zZYNp2OkLQ2It2EtHKDegVwSR
wU+gyH4z3FO5SkKXBlNeDT3Fq6O20fuKXGvnDGe2j5XzSii4CSxMb38XUWTjvZhR
uFSnT0GqPeQysDvDhE8iq7SpaiOBBiuWn3NJEj7j4beQ92UuC8qsvWfzDZLCZ6wU
0dSiLgOsQMPGJoj/ZEoJt9j9oPFD8kNNk7vj5Q082TgsLrqV3qXj5XTeeMsXqq4X
fLBAzT5pI1uyjLpO2W4QKaZ+u/DoKiz2vKzuWaOIcp7HnfVM6yR/ERgmvuW3stE1
XqQOLIWWp06lJQBenimpP7L8DBBIDW6ANIqJupmKLgBJ4h98CIIaJ6PABiLTYqR6
ius07OpER/6W0mHcIIZ8pyCH2OlcWt5RUQk7LkrKMClBtv5Wc64fsg4yQXWtNC3o
dXPpaX/OGb7eiH76iO5ORkuCsCjgxzZTucfKqUimzZpqGxDy8UZa3AjnOMM7Kdm6
yDnajH2+b7idjZjm+WiUfmNFYeWwcOG5BbyLcsNv7IFGy/13ZKquBFzhPni7Gzmc
IJdIq/Mr9lam0LX5+QuGDw/0LyuLkhcd49WXkWrLOSP7+ybF+bGe6CUoFT2aSiwD
wIPUjEaPeycS/gkTLf0P0hS0E+W49Qp+XLKSXIscJVGzox3issMynFXsPOvEWVF1
ocLvYidg14IxLfs4VWc3oyCnneOqCVR8lrA0NOG2LzaXy6DjxgCYHEIug4/7Bscp
QuR60xkuu7NEXtRy6WwvOUzOAf7MJOwU3CuIygQ5PPIoEcGsxcjHIeLGF/zzWGmR
ut50BNs3Buf6Lj8x6aSEA+ZI99Ws9oxhQ+Ghgqp3M5E4l1q8lN5S331Via1scIRL
jmnclTWupfOK6wWzsiXfZP78vCxwIkYAwi8UcqKG1L3ne2fKfydKntt5Uf203DAw
8yXRx6M9DbNHM+khPijiJE0LJmIc+AUSdc2Hj1VgjKcmc9gfK5g/dlKCok/DMmF2
9hfJZ4HyqsbDvfwAlIiNf460n5/QWcHA9oZu9+ctB8jai5AOnDjbEn6J7sQH096w
qSELwoO9d0qJOks3BobDZDDcVUEodAbF3jEJS/YE4bQnSJJ6USC+L4NVpFvEkMk0
Dky27IsSN3Kt2XYWOdN0b6YgkIx/xf5n8K4OseKsrCHtgpqRJX/jeTXtlkKlHs1V
5bsdEiu2RAWYYP9Z9mfS4Z4PWjdba4qPFmhhZphQ3HWN3Qps9lnjX7niPPPCAoUu
z/u9WKrkiIL3ENc8LGoRKCfGCGZkhQV4P1d9ZemPxv1YbbRAo6XcyRo2LChRFvdo
KIWXOFWKeaHmKRyePFBFP5fE66E+oDnYjL09K3zQkUQplEsH+3kuJ2bT76l8KGD3
cUlFPx+RDgz5BldLxlZmHqhMurEjdsW3UnJv1CVo470SUrcGzmCJHMq7pvkXJ4hW
0hSr27zvyxd+sEokmhTn/b56PKRtQWMk/MMvOxXtzw386ct1BywfSNkr8GltxYUC
z4gYZJiDGmy47a+oMkhWimqirBeIZYJOnu3JlbdlEUrBHROG2P3LA0CCVJMAjyAx
xtIhAf8kMiOVLWaGkih/bfRcTQpcQIc+HVxbCzktWSvUNoM6f8fXzu0H/4Z2gfT1
6mALs8DzmddJB2XvnucitY8PQni7WlbcEyG30Nuv/5hR2f5zqi2gQZEESIfhlByo
V9g/ekSRWsZpuoU3TueVtJQVZjKa/cQmlkZvk8oA9HuvOYoARw0zTcB/HCQ1UXEm
UkmAtbXBQEMwa2GWpcAWsinEbLdtIvkihyu75iunRHr+M2KmnDwDbmSpLnFQu1Af
aJMIseoH0BAtz0tcMCV74JVok6DeCm8/oCbeYtRWD4T/AKV93u4GiuAhzGk6MBGp
vTwhDf6W/It8v3q8Zx2JyEZ6y6vVmESxy0JPkaJq+PUuy6ILcp8CgsphNXiGi7lf
ODZ+HhHOtNdIABc03biV1yDx6j9xZhpIzbgAt4vC4vAPzPAAF+l3/FgGa4cDrm+R
9gjtdZxzOceYcHD5hW+JmKzzMbLiGTlRsxhaqfkTSrliMZVjtv4jdv9XR2Xw1PVD
taulZ/0+K0toKTRWG4fK1KPYCWvFoKV09srhHJZvh3+ZQ854mdWDONpp0LRfQ1mj
vvqlEwm4mmoOVHIzZswMzc4x8HFWF3Rj4eF09SAvyigElm/W2FQniYceIAgJQ/Q5
CQ7klWY8g67pLwDnhLzY31mHW0Rj0haC2dwyobRmvqWeWSmWZeHnAoIZFzLK6Bb9
v6tIWOjfg1y0E0K154dVo7WIkdLc+kdaEMNMo8njwgLL6nHcx4BXvc06gF9FUh+k
GSJWllZtnob4wIs1O+/T3CBZD6p7ZLC/dv/2z8+ZSuq4XXdr+mTAYAFbOcLKf09Z
0PQrHzk9qQXxmAuHeGPAQn2bqoLQvcGlBSXcwCDvxtbh9K8NO1vkdr5IFUIlld1M
ALfZ8FjZQBE4aK1WfYIrs919or4LmTGTssjeS+vj9RJeH9hEAVQSqtbYwTSlrMDa
3BO/dagDclnZ1QUNhlz3re3j182j+L+kLvpMROcI60D7d97JDuTQQ/rGnMIesQ8U
HiNTw5LFJOSDcDvEjFt6tPfGpPbmbrE/y5xpvNCB9xq2ePazKTQzSty2FRTegJ/S
ywqdD5Y2n73rKUipD6f+ljV3iLezBaGqYaZNUzVbY7IgzqBSjaW9ogjxQChkGnOd
kwDMn51UWGGwCHXISXKwSwubY0gKvoC4RinlNFa0ElMa7gxdjfIdljKSt184qE0M
RNFOIGmfcQ58HYNDKB20g1KParF9t/fpQta70Z5h3VoFx4slmiJatxrEwILyhQhm
cvm2x3fTjbosYzb+rpZZXgql9PKWFmGsg3QI03RQaKmnIQq3OREfRxlbos2kqD98
Slk/Tp+7hZUEX02iB62SAArVg3lm2OtsnxrqWH+q0crQU25JH92TuEgQ+Mb0cjZQ
YKvHgKO9FSfHugzF06uthaivydHV6NbLw0wBzU4ju7pf442NuzhTuRRgTv+BFrGs
Q08ea52BxhGAd2wV3YtuTkJlUb1eiuy3eitOFeXsE4ae93N8jIlB62tWqi3P6JTT
pnZwLQwneT8BKThqIk/FrfeB2SSEEupGuxpWWobHtQx/oVYgQRzPHwPW4DyNijEW
vi5YRkEUwi7bqcgBLffHadTDkwVaPXt+1a99wz0bPOFdq7Q+nN1te56TPQPrqYME
OJHdRSnLFCwEAGnBA9uPDjdjFAvBIvrora0bym+/OgEFErzNvSTu+VBSFNUapDqS
wPM0jkvFTp8PRoxDdzOVvtz07f8QepwZa5wcVMz5afPG14z8XEy4EpOiHoL3p7ha
i7QHZYsPO/10cgelCD5EVj1pZrBSOnlPLFUCxkufAtA8PTKz+e4xbn19/eGrbUop
cdzHaFfHy3mkW76Xqu41Xz/Kh7RbzzIMlbUxF3q1LnrSfbMb05rzOPJFEAINPLRu
WtRz6uLz91l5gfq2He5gUxFV03opgAKbXfZgQVGuZHw3pJJ5X52fzy36I434BsIa
`protect END_PROTECTED
