`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SFSejQbaVq9Sm3NAAythMgzHJkVBQPgbUd5ZeBCPX2PZTIVyx334ENobjlvHak+W
mBOqdmq4z6ugPijLKOQ70F7ettoMpiB0BHSIy72KgsQgvdck0L5RZa6iogJlUZSx
YLqQiNO5hh0vnapMUSmVQ2iSFMQ9oIhTfQJ0za7T3isiBAUcVJM+WuPXZ8q/B/Yr
Z5dKO4Diz9UpMkURWAqp6XAbnQnfdUzzmmOdEKyE2IKnLGX98K3tc96yK6wauL7O
z8bV6B3ZLHqB0nnCCOPUeJBbOxsE2N2eQLS4NdhzDr/U8HQb60lrhB/8ZTc2eFnC
UHCnHO4J3id/arHuaMDHfCEbOD3y3ffV3KvDvZIbifXV0BYkG+sEwFMHIZQWEY8f
2PKgB/Cl+b8Cjqr5XiGEJbj0QllF6TnPf5T3Rus/URlBSA9wWjX/chLEXuMHeghy
TiXlmMg+yGgyXEzPTu4ZR/kwdtNcQfuurp2+WJLa051DbxP3KbAT+zK2s/6K7TiU
JtGqgROiD1hAjvbkjPBlCs8uOAdXP6tHkEi+YWNgXgAK8SVEynq7dTMrHmpDZMQv
1N87E4Bbn2cEKrav/bOjqBUOB5XUHJGCcVriMLHM7lCRnAkWTl6V4KhpmjNRhx1s
v4ezLcIN95NZnHGktNFUg5qFVW77DafbfHneHVlj11vs4j8YrkkHrwVPxt+Qr586
t2JdIV69bHpPLK3462eAsJI/2ZRy2+MU0oeyJ+WLfoDI/0WN6dOD4gvyk22dZWrf
csJD6YfaRk+tAEovYr7COK2coRkWFmEGSxzkypKHspY=
`protect END_PROTECTED
