`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QDa3iHsACJVpoQkSB1CbNormsGsMxSVnOyKUpXqtGXswh+spv30kEHxwqoIReUhg
nni7TalZQu7yX/8hn1RWR2aUDxWbsz3vRylCD9RfiloLQZcJRcoZ7B1jRqHAFRTx
yPE8QjrsGfWTX0HDcH7KDZq9r+Rl6S+k6m0hkKGDGY11FwmBrZpuLP8Ft5phwyug
+aiHxILiHLHlIZFoJPNJEpoUPVvEhW4VFJi9VWU5KglsKYB3yZisM2CTa2MMN0Z9
xxZiD11pFq4TXY8UKK/Dy0GSmF0dGJE6jeWMkOs/PYWB+5I/L3TIB2TtPbGFjuyz
fzvZdg+PDtFhVGAqwcBkkCFWid2zab/xFQKjvgzjfnaDTjvZ9LAFj767xLsvHuLb
Z1V7H7ZgOChTX3sTY2T+RJXLsG+kJkIU1ydakWijQCxzE2BBQDnuvtO8OW3UlE1A
ag+S+Q+n8RMYGJ9jxPYNu5qiEM4duJ12g+mJftOFcuPWJ0XnsGYy0sKocm80k6di
9v1v0BLB4M+ACigIdSKIYPECwBGx8XlOidnD+UPi2YwUx/uJ13vNhIPrAE87AZ/H
cc31IKLCQErXk0mzKb8cbIkEF2dkBFBqwxLoJGlw2NtFRaU9At5AYDE5TiKmopdR
eQpdluVeDIzNZLgA8CwX2m9C9bC5N8vICX6QJG4NtCuMH9mkIiTefb4FPUBS27ES
7PujilpFLE3Z19qNGzIkvL/Cu6ubqVxgla1Y+7Purq4wSMslwfl6/Jm8m5Ma8+3x
XoNFG1yp5YB6FhGA0dUDqo1/Hd+2V+TmoB3xkneOHqIdo8L32yUVEIai5OzR/L8d
0iFVxDqZnoKOvQNlCCfI+AbLgzKSoiExbTpJ+nGhUNHy6z8ZdoZ1Zj5/Nif1iJju
Qy6vj+I7g4GV7FWB/R04wNHYshgXNb2TkGXdGAvDk4ANC40x+QxLAPsxYWNhPR/4
cWLLDzW0XndzB41mG1Y1nTWKhDbKoTLVVjrbyI7RLho3KegHb4fE12vbjXIv4DCE
g2SfqJSI0PoxVfY2yEHMZNKvJOZ2qqc4KcvMAmch9Poeq9butSAZK+IdoOZL7dcu
ltaqFU1O27L+a8Cti0uYs3/0+17mdUC01uRhDpJnGYPhHBT6t6PxbWsNBg6IXHBG
9WIT2+MnLQGrhpIpAl7A+zp27M0yqzR307X+GxiEzQK1hG7HgGMW+JbtDnqEvemG
ZmhcSlB/ghtBJGOKHvHzao3R/5Onc/qL42kdPuJYy7gQQ8RGnZjWYvmco81EuUXa
CsmJaPnzA/6qilLGa4qxDE5xlHV7cjKFczYioRn+P3HN1v4C9IVUlxgK48yXAxCK
DQMWysnHjVNflNbDQA2MSK45zi6e3Yk2oQKGj/Gzk0GUyS3wRW69C+yXESiTPRlz
PxqvcfYtrD9cthpMh4/oqMygecp/f3CgSmE3k+NttGn2PVb/xwglIqa74IoCeIHf
gff86buynEvx+XKnYsQVqk/MS+6BMR5xqSM6OIncruu2KfLG+87ruph9SdXUCEGr
ko4HGsBdP7VELgiZt29pA4005opLV9XozW0hqIFRX+ZqCAg0Sq6szQs6jXF3aCbk
NmcvMFJhVZanK5HH1jAvu6wLtUg5E8JOMimRb5uiKnRVfGtmZiXFHWn8ujTcAqcz
J6D0riuQ4tQWXHpuQ08ysUCZecqZ205jkZpUTK7HNrgGHj6YZZN0BdF+dQIF79IK
Vaoc3M76BtS2XkGF/g/Ha24V9vHb8lB6p2DxpVo92gFmKf0MHm2c6cM2+sN5P7MW
t4dNkf3I5ENawpplKIdCu8rd6kcrpKpBTiWvVOGQfbOBL9G8W371eA5uc5ZhG+yJ
sCop+2eWHwAIuht3JoJT8SajhR0Hmg8hd3wA6wS0VSKdTuRSvW6oWRI5JTRaHCob
OFAR5Vpg9EwCzrjX9/feT+yxI3xy54ffAVPaPPnhFrCSbgRTIGs7fgEyS8xupKEa
iQVeIUFg9dXgEMG9ZFeiNdOyEgEQMy5DiTOCGA2O6D9rOkZyJcl9wx1sKl366wPI
0AvOMIqkcqsGg5YTaVL5SNxpnXUAcqSb28pdg+kIvmvDi6iukx3z66GrGE8LHVPh
9u3ReRleDt1nk6U1HWSDAl3wCK6dKe7jfPgE7BLSFMMOhU5RR73yBUI0BdiGArKw
P4VjxSowPGRVi3bD0a3Go/b3FpbjaNgwBd+OhCmAw5cvqfkeE0e7YsF0Pl2HXWtF
8eNwHLET+c2pD0L4N3E6iwZrqa6BPL+gbonDON/90H1Grb2kjDUAPWQfA0AvvAeI
hI+2CBCiMvWW00gOMDm7p54eR1od1ka2DiX51VKLxMfCpsNauN4NwdBAxC7JV4yR
4WnC19/9Gm92Jr8assWRCG/v0U9F0I5QE1raklBuI5DOsLVNQW7gFhddBM5yPOTv
gzcPuHR9qNtrmCy4fi6dPrIUwhva3aVluPdp7r/UW3Ju4zHoRNy7JukLn7DNqywL
I5gq6reU3Bz4YSz3TMcdINRbHVqKu/6qcbAtsgd1HSD/bUkh6z4htzDDTnSlgxZj
MXD8hAXgRnJOlEWMscP8mDkNH+g8NDxG5KyZiLOoHJ2PFh4M6HiTHhWQDfN5SWZw
CznMKRXq7idPH+D5F4TVLw==
`protect END_PROTECTED
