`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59ufCGoDOVDD+jDbKKl4fpjCK+dnjIhN8H3kezOsPw2pF6eDLLFrv6WvR9GfezvD
0q42Monn7c5KgGf5QoX4G9Wi1fCaEqtcPXMaAipIyIBOvebHw4JO55YqJngMpeXL
7lJu4n2A7Yq7MKkcpe3Cq0qOK3PGj1sXzpAO8eZ0cLTRQ3cp0exaEDMmd2tiT5wk
RaAlXV3Mh8O7FGTScD8ecXy4FjG+jeIij2Fk0r0TwJs8nGrDuOpc1B6LY2sI+Kkd
Y2rHUK8vlcSLIcTp6ZCWQc68sY+7cmlTjpqMJV+OTcSm9V2y2dDE1b8TituGDFvY
BupqeE6mFv+byksT5HK53GQbILqoY7IHf8oFbP5nRox2w6xTBNGR8HywVKzoO3ER
l6qXvP16tNfAGRBrhrUQIm02hYL8k355xyN9jOnYl6Q8wOfqpe/Ab/Ql5FsQxFa5
1/wG+62eQZC1uWhhL7Mj6W8qLH8yUwoD/DxOLpOCVlkvTspuFwjbLrQAeRJVx+Ss
/cb0rxezFmPIrw2alVSaqw+VNzJ7ex2LBELP+ab0qf9yvlnea03Ve6PPHa6fZmKf
k1rHJzVItw95DnUZ883Q2T8rHr7dvFb604M3jsbSGVz9cFVmHaEz+K+uG9M9oWHQ
7OIQ6pPRvfNYFpDWJn0vx2FsnKHzTxTtr8G0iVroolE2jmvAneH7TUMO3ZaZ0OCJ
d+g36432k2RxabSU7Xm1poce3vdCFKHYkQTzPlxTDQhkBqHfzWS8j1M2Z/RZtFQW
7oj/Lo0pdW2BpJgLRvQG+sf6t8ZQlw177Ie7bfPcisBuafyLCvSBsS1ctN4PgD/D
9R8LJFmMpVqYt9vaV+ayqjvhWMdCsll67JA3RVzo/a2ewXCZinfh+PbtoOXVzPIr
VwtonYJ+iPbpkH9uhmy+Ruwa0342t/aARhrFA9lcBM5N4kC/omj3mPLX78bOTBL6
rGtTVROO+bDY/qrlEWAN4s735tvBMDwYrt6mwiukz6K6omoItvUNgfENydFZ2KN0
qYrFl/DXlv8no3iuvDj8EC3tzMgrhTVTTEd29aFHREyIbFnKO6Qw0uEuk7IYOSTO
6ZJmosED3Sgdvm0C0sh1zsz0S2NKkZQLeKt6043/iIZQdvpOoFXC8RTskGxv+4GQ
E+fuL38gp1fElOyXBhKjF2xlVEmk3DUutSgK++7olkT2fWjuBKkLv9WcJg2SFoPZ
TkDaaPVlsJd/5m/BeHePMZ2r0fVZJ6X0nxdJgo7mulidvWBaxogEt6eC3gOV6MOr
jLHym4GIgq0YtFqXkY+gjG8viDDncW8lEKlpnhf6aEifGgPKlwWDedYcQCg6XzAd
f+Xo3DJkyKVCicIDeHsfVKkjL3UglCzVRW9Ft+V2hOm8oL+h1tuwFgfsF55zSemG
8xLpuyPjQCIwsrApfCABz1sSR5vb4x+cLSysAmKs/RyiPP362mcT2GPDv/mKp2Jr
u+J9HvAJlfCa5LD38ep/kwWAfbUQWuoEAfJGfAVwiC7mOjA8KLIwu5UinqcUHkZd
9ZMl7XQ9gSw0f5UVP+e5jFz7AB3MxDV5UvE654Rh8zfYIV3sb3Tz/2BeylIHrE8l
VMYXxKs8BCeAYKD7Of2RyTx/JABSdF4SKppplv0Y62haxXuVnJxbtTOFF7fg2FRJ
U488gAxzxT6EpuFhaKrZ3SApcVpZG8FEU8RfSXhHRuBvqAMXG1TP93zRjqHAiQmV
XR2O1lkJAxymc9kYQcuLzJ8u/h0HgwKNlHkYh2PK8VKD7Tkyht1WlXKR2GnX+lwA
ngSoPR8t5iRU5y0BXMp+eRlslyyLZ9I3C436b4Jmvqql+JT4qS+LUlAuSmlOx8Oh
3g754QvWwWmOX+zvVBJaUyFZ+sGGjhhyEVZe4a82st8EIhQzFs/Vrtj79Y/rqdV1
HuoxuRlZ+RpMy5FKuX1WwVPD/K7BAF8MbkuZD3g0vEqEP3hsFZzLnOOcBj2WIAvc
E0vGU9LL9ThfAd6YP5MR5GhBdE54KvKM2giyGlN70VkgIkvIDrTrDweWygPRbu/V
P/2fA0l0ypKudw1SODJQ4SCVwioMTGkD3sMbxu1KdDoHt4bjHse6WeqrL2i9jkCp
lLiJHO03ET2A+FeT2bwqBVt1S4ZVEABR4L2Y3MKQH3zQfdSL2c0ppblRyY/vwlPj
VIQmQOqlhBodjxHcPMKdyesISAri/xdxD/KkPYXi4vH1pM3MdnpJ/Rt+I2R5Yfae
zm5DG987qFypCt5zWLQPcWY0u5n71gYricBG4Jx34qmLHgyNRwy0A+kIrR24d1Ib
AvNbBXpIjvI2drHweVgELSoVdQG7c8xhox5G2DwrSmOpoWecWf8FduId3GB2wGfA
MuwC8MZlBjqzharFFqmquOplEdvMKaK/9SueOfyHd6OiA34wwlD/iE6g8HBAYaJW
bLcO/PuNuvcIeGmMVIsCGwHRrkc2JkyEtabztNjbScKzhn4WHkRKt9g2ycvZVMaw
rPoOk8GLcFIWCleAsZp9yOH495kbVozp/1ibXmDeAdRhfTElgOHTQb2ZfK5fL7nu
KRjfbt9Tvwqz071mApcqJZ2p0Ng1HQ3jHQFeWLsiviM/dQj5L0yVvwBBHiN6xDTa
mKT6WzNsXTbPXYWu5x67rqX1r0Hs14wQKapiyWwBaz5cLTjZnFrPESNLyeDctqXe
LZwUrvRVFLhWQkMrt18DgTh8iNTbwZ5FBH0kGy0aTHA/iaJWLWA4/8s1qp8EtlB4
ddrS2sMsrHxaQ57Zzye6oYxAsZ/+D+ijqZzMkbdMFyDj4KTRYkeyHNzm8Lr5vyud
71koMwafcMV/+k70HRLITHakCFV0+vtseJ1nBipsNlbqlEgGp0aM/w7s4HB8xXzn
Fox2TsfloTBhGXhox9o0zZqz8BIoplOpISSmh+chHXsaFM9drHbm76lw3NtddBwQ
lVajIzjMb7WmkB+ItvGMY+9xD0QehWuEZ9IMlR2+HIAxs2AyY/iQiwkJCtmj9Jl6
SXBaNnRzX9e6jmsDS5zr6UrBehGbz2VI0y3x3mDhKv9PpgUiwXWs9Fei6Ay6Gerg
yziOKTceaTePDm22s+2y5TcT0qJF2blS/MTldnxNQyluyGQmwiwDrP2qErfCbxlz
rNnv4uKD0VKjW0kmBZziwyaw9P4KelQ8GoO/8JlIQ/lOOsmW0WcAy+VAo8J/xN+9
nMxSFYf82rDawOdnnwDad5ZFq7m1+UJWfEX+C8H3BzH1Kn2jIjHS1gEvMBa65Phu
MDvbve+2pBj9hFGnR+nhnx0W0ltzOjZYlzNfEC8xpE0J1vwrudgZ2z2mRvi99cVo
UTom9/RHdFJzuQXkERqpk/cmzApKdmUk8tQ+ODueHGSgVqSkCRKrRPa4Fqs+fb7L
3Tc+dF3xUN85OeQwP0ExlvmTXPINsrWKJmHBOtscSkaKBpvmrYHQH78tvJ7sQRMV
gpWsmWOcXOGz1TPKZgacSQHMWGimoiJ5vkQ9QMdCEqpIoydMkiWUVhm1CiqJjytH
uSIx18ed1dOf+Z5GnY/fiJNsnALb/Gac7JGBdLgMfLi7qNOz1ULPP7V5YO9q5jkm
u72P519ilSX0k1dNr1Vi50dfiaT6C/ciHWBMQpRYKahZDHweRarWPv69KItFv/ug
exGLB4lYqFI3Qy7pdW2RPH7VWPHv+GOok4eqBretX9vKBfY0AgL6xqAMXjo5bVit
ovgktZwrMAM3sZPEu77cQp+9hQ26HQmsVBh6DsLWGd2UWHKRGwU5oYCH5iT4wDxZ
h8MnF4gSE74k7jiced6hZFcV4gGwQT4kou41WQZT1YaUWSV2B4vuXz1EHpFMFG+E
XK3XW+35Kcp9jnXvXex7aIHgRolTD2f9GUXfAhtMZmmpNyEvfQ2FbOCnHX9IGypi
+n9GFn2z9phtLIoHbzb6ZUpmX345qybQckhuxF+VsD1zcS303UHOJauJRE8rWZYj
cDafStKwUrcDDRHLlFKF6D4LtNXx3VdFpweAICo1gRKPoifegzxarc6q9PDnU8jq
+mP4ib8ptQOc+pmFxIWefWR3Z27BssZPJ0G+ykvgzhSn7YdpLWZTKpOJYr7YVdgM
mUJ4gqfUbmY1WDn5Mrn/6Mp4lLC+EAU0S/+BnLZRK5Yw8XAoR/Ilb/bJYWQNsKTN
2VJTs3oa+rlJnuTKfJC8yvn15Ip+VPqNVOKgTUO74faZptvVNUsPeYZ9kYmPmvgX
+Kl2oc34aWqsadp23ufdFr1xC3GUuZQ6VS7EXGscPFDczfksbfHqlf1Vzb/BoMGG
cbCHouWkR3jfEehm6cwUC8D6q19hjBpwsCD7Z8EU5C+N3Ka6X0zn4mLjb+ZaFhEr
OD08jfPy5pdDNO1QHekxT13wLwqdtixG34oNh/mQlKz53hcXAsEwEP9Yrytn4f2b
JPVmJlJkWsPGrJqFcwqh3SuSnKjJqiuMw0xRzfZ9XvRTMIFJkW5d28y6pM+YqSZl
+aPVabo+lIUZPi7BZijHHpUcpYSCXxWNvtJ+eKF13I8iiLMIXa5fBmD2Hp0PmNbU
5t6L/f363ai540Xh4X41OLSKXDVgngvM88/0kFWRM6rSIJyprQpjp2IgAtImKTfK
DezZVq0Jo/BLA9ho5Z9EiIaCmQGzENV5KPqDeFBeb8hoABZGcNWnnyTWA+4qLeDl
1Pr/Eww9GxonJ/TNr+FZ/bPIcR2qIK2n0k/JxNWkFChrdgEoriwOENPPOCpvzRZf
wzhffqY07jWLQZk1iOmFfj1SIWteyaP9dwPcShKZv5i0qN+ITWrMHkJlkY6qcNze
mPTujEuTHA9VwlGgewzBXVUCl/L1jHUR/iTWdzzCB9be4MZdWWDlDlZ20bvPu5ft
+hT8d0kIV2qlwH36zJCT6v5mXEdbkzMbjhorCkzbZeNhfAfIVYiH0O1A4yhKPsxN
Ld3jGEsYB6mI+Durhu/6WQaRHjcZwIOAOUQUKCZPFlTzqfMBQDwrRSYBc7UFcKez
34cMDFYOWxEthmmVTLb9uemoA71nFtLFBaetHlfTyaa9H54MOrqSUMum0qG2WIrZ
ARPrzTc9uHfELLBsxQ3ftKDYkJ/Vy/KliFo8d2W3SoyxDe+ZFlq8Y/5yxutPwbqz
dIfb3X8EC3NfXNVUWujz9srnPBioe6SgbsoLDGCdrmQUqFomyNVOUQvDrhDxvWX4
0LeTny+zf1n2cudNq1XA3pnrp4Lbpz9U48zk+B0CnrWKFGAZhNWDf0JFbjPBmkSN
LQymS0F+b/jI9kS0MlLWB4sBdpd4WkRAx8j1Bl0fL0wa04v24aiMITl1PB+JtPVi
eWJW9P+8/fca7vaiPZS8gToy0dfHDdOdw8aOOHMyPk2PeYlT9LnsYHCoYfeNcH/S
ev4qQiFnDONHOJFjFtnA9GDmydWZONuIugeQ01YbZn4XhM5T2bz/GbNKrHQCfKPe
9ouSMgoSthOGy+u5zgLWa0j/jSkrp0LIMJPd5cTbXt0hcNz7Ne0g5yk0dN709s6x
w4jxoxPCGboDqiZh6WSgVnQzd+mzTVIMsaHj2poaQKsscbjVRGZKD0UthcXTW8/D
DufoFFoLmCy/rAivH+swAhOlZWbfUd7b1Yqwud1sNaAiAAl55gquOhhfSWLxBIh1
Grx5ZzMZB9cO9XxIlWg5mkTPWpk/dSs38lsTKBKILzbHqEPg8oMyw3SDYMJbT9Ty
UAfPlE19xXX08epRju6YQc/sbJ56s8z80+AkVc9PS+miu8URbVEVh6mG/I4XWdJL
J5n7DMjKVW79OAkPMDnRT8Yu5ae6auStXd0DX/dv0yJzjkNXlonuvABh+XAfSdNI
yNjKdCAbpeZJR+bW4pdS41tXdQMR4qOITs57qrLRh6++fREXvqOf1lbovJOJXytz
8IkCoYqirUZIP3GAyiK4VOdAujC3yNeyX4fMjrKwLhTHwcXEJwtggWfsPbVedYkK
RQHhx90O4uGg7dJuuXossRX+gsmFc0UOpSF13cXBkaqXk7R5Pprnj3bQc+Qm82h4
Jy4M2WlBrVWuIO8IoSTnLBxBlCCtDCNBH0kiicK126JqItbNIZKlQhZxkUPBhl6a
dq6MPrc95c2LGyJpXafhQ0sFxhKON1YvRr5fIcMz0kJ6c39/fk02YcKuwR6cK8Hu
XZIpi52cItTS1ev/wMhrfUah5iJr9LlLC5vtade9YiHLYfR/KL9M0MX3dXbSqvhv
z+925fRheQ3nJFgG8DdFSG/apNCc4eer9VH72SIb0JkeXOZyGxpMwrDTvpSdp7oP
/nHbmsQx8IeJaVwpDTKdcNj15r1BYEabZ1CP7RLGvx4CJysKyQSy/RbgWwtKn/t1
asaYQxd5NSWjXAJLCIGJz24gf00UPUEdsnfmydPomL3JYl3URAwAXUfkZsqxKkBA
f1dPDzPqpYhf/N5cuiZZYkw89TEV7SnXgjEG7wDeVcjWloSnCHMTYmLBesmsGRG6
0J973msf8Z3YagZ1ceS5oO1wskonRNJoZCrLpj6AgSg16SVMfjujf59KWbDal+PG
wwxQdP6tJeF+8USB/cyR+lLnkUTEqnpBnbfcp2xI7BTXbvfqfhreWu/pYYATNwby
P+/w8sfHfurduv48+wWsmL0n8nj7HfArWypTMEcYJZfh8Vz4HkKFeVI2NHq0GYF3
wcGY1xJUc0LsFY+yNYdvsyedrpLvbkiq31YdY2pxQ89aE6ie/LDkxNGex+3sYqbk
cBkJl7tM99WDtc9NHKm2PMG9jl1ZczE39X8Nn95P4o9653P+LwfMmX5frlZ6RLhS
mHZ7FkaUs8sVUsSFwA09llg3qrGasGhn0/lpuNvwUQE90Agm/Pyn68ttwO5sIuvj
97W/t0VVF//HeG4tr5t8GNqR3urB6N/p0sf+KC+3rGdJiBfe6W1+H0NC4RR5RxoX
2ph0FbSWwEaYnHeWgTK6sPph0dD9SHJYGeTSnL2HpoDQ/2K1H2TNSaTmyoj/o9rt
V5O7lcDDWnmwdhv2S8jwbZh5Imy9YqHYneLP+KJKibhMd84i7LbEsgnxdF6MwQxw
gCnFXBp95Xdpwqk2kftTNpxkqyVu4DmwiAFr+YS9XDIX7LWb0H7ZIdY8J+1ODR70
IqW9vdTArk9lYcIv7eiy7uw5XxM2bccADxSffQ2VzyhvLbS5oFJcOxPttR6Oj/Oc
MukbFtwS3i8SypouTZ2Wf2fSUNJYm/4zykqJTbBvu37p9p791W0PRIkryaZOa5N7
aG8LnM435GLWc4CzsRcfhmaVkKg3pz//CZ/Ol43ZCwmCdItT8mtIsgn+g8E1Q+HH
K9AoS0tH9iqDe8PG/2kj0s0utWdlcqcDbJzRfIqVNDWzDaxoyrMCB2bfzRln94NU
xnT6L5YJY2nL0h8m6bmJw45LAIExI9VMKEkHIol45U9dgYHroqlHIGnNlej9veaF
W8ku1Av5KZUi18Th4HErB41Mn+5e2DAjE3kMdlfm4zzWIkfnc3DuvaM3cdkaddoJ
tXmA+GXzrSRnfZVCsgb9vQATywfmTsMWR+XEfjkiy0/53GBlxzsOu3LdZy+2wFdD
xpJgpihPSc4jSgPEb+7Y/g5ADUADfGoQVleXNA1eCUV3rF5oNwKrLbtBsYsVlsPo
LYUo65UIh4xhdAeKh/CxW08LAfxoi2nUOQGCj8emhkESVSo8RHN43KUGhNCI7E0D
623wvnYTHoS4fFEVo+l+j/ejYHoRSUCgkjDgBMVJKPrYOiF+f2iM7xwbWzOJrFQ4
KNRHcVBmbtun8gq7BF6bNlDCBOtY3HIMVt9EVJUPgtiPa0jasKXDaWZbmsDhh09H
2mTJW+AiA48g3D1HEa+mi8vN4aD5L4wLrKcbU4aSOg1MYkXnw+bGTPJfT1NuI/y2
ScDLki4DVi6HEoxaI9fuG1V0fT3mopmNTk70fC5pETHJB5/+nDHTUKE7MsY4F8Gf
VJIV9VWqWPlrNgzJNz2zKeUDz1o9Lr5NfnTu82XFUVZC0D5J5tRwwpHEl6gUoq05
lAhrB2NAKyEuxUlyt4el2GdMzxQSuL+HefWwNbvo5YhLpfCQQTiowk7SDklmYKWx
VCDjVf1AgEMHhq0Ah/kZkWH5/yrhJQ4ZUU7On7G4vR2wVR32kuHarETWjwgjpIPf
JXeXZIixUXthJIC4DUCiGWYjB2Hk2ZLdDWdTnQw9UsTjRF9pIu2bjionqIfeurCS
zB3BUcWTIGkRvL5fCrDr8LplRUv01ytGCFx1RNVCVb8Kte1h5mO6tTunZ5LaumkH
yR3YRAVoFhjmyI26MnqMNiFb8ti8CwXb9UM4Z6FbsNYfEdH9F/RfNj6kDBDuedTv
47ZFaOBC5dw2DCri7anivL4cFrdiGA5eaL/334MHJ4BC5vIJKmrhiEaJTO3myQfK
Tk5w4EnesObPzWE2yv8i7+0SBWD3PtU+1J3IJlwhq+L5WcAJPps0LlUimFEBpYYN
kf475R3392FHt7zGMA23A9TJ+Zup+pWHcEQJoIhCqLt41o9BIPdInXB1PfjpTHlK
xH6CZ4hz16QCGyiLmgEBnSTQxjkhbaAK4Xy+Lg5A+8PYM38A5Xr3y+3SjHq48uae
RwziL4WVtqthYt5j5EGxMM3doRTAOetuEch4laoIIzLsaDosYdF22fkIzJnucxUv
9yy0KVAf+MQJ2FRog+RNUBwDomxysrCoIbGVj5uW20zP9obp7YWUtLoynmCLJ7Fe
3NjIe2eSEsLM/d6DaCY81tSvnd8lA/hb0zaZwt9rLaPZjihpxwpOih5uPGP0ap0z
EVQQ1kaQwLdqLOV4XGVH0Aqg2t7sNIY1+0r8bD4p0quSpR4uB1epgaoaIcvrsl2a
zFjWDnmm/FMuXDmUXcoSMBE5GyeQEZMzGGTHLG50R86qWaahzZS2KwzG1jZmfd1q
C8Urj+TDGkqY92j4KSZClYqluUqMKBUmn+NW9f8/CsWnJxqY9tY7kl9+u4F/xQ35
WXLdmY/JTExjTR/3/Vt+9KFd6aLr/ALMV392kFStK+X6G54TDvUPjcFtWtF1LlSZ
1lLWxmn7lNBmPLqCF3/Kunji5U41Q/loNyJzIRU4HqE=
`protect END_PROTECTED
