`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSbC8x4ZWcci6woPMWeVBcjmNVoucjbIm79Xs2dQeEtPv5cBa3/gMSKfQDp5w9CO
/0VXhEIikpCw7PP6TQ1tGwdjNtj8qHSRgUOUY58uuJSsy3NT5hdaX5uoQ4cqPe+/
XziC0SExiCANreTMf5lMoLHmQ3Ex6tpJ9yW3U1viJV9t/jNIb/Zl+xUJFGaM5N5E
ctv3wGeF61BcslYvs1zcJG+SGIibBGiAAWYSuDUGIZk4kKGV5YayVjuVPCWwpgYf
P0Xad1AbR7a6vMXhjgJKPNyPBnj6QnyQ2iR4B9lvWIV5XeFo1LXqJkU/7+oal1po
tEdicRKwt9F0HGthcwYtrjsp1QEiAec07NiN1OhR+EXlygY0S3mKZ6qIxeTI8Xmo
i01koSLt23LUeWQxLI9gqncUgkewLIALs5kfVpZMNT6exsK8VTuXPudVdaoiVN5X
6w8i2Mnl8+MfgZUhq9C1JF+FGzCYGZUjFl7h4EZjTvsDDCAfWwsk4yxFOfQ/ynrt
plkBr+XZCvOM+qc+FLbSquU1tBDqAWa87hsqYf30gpvBeVscRjoQczQCGVg3kyZ4
UJXEG8WBahpa2Q453xsdgOC/67DdrgfSGU3b4LM0rQ9yXj6T0/0gsbhhGrBEiUJ9
63OoGavzzAebvHKqt18H480azdtVtBSSkq5shj6SFIua55UXZIGAWrp/m6q3Vqem
uURbjAFtEGn0pC1YvDjP2sqXWpByqnb4rOX148W2OyH6nbNTVmIKhhH/JgxKY0H/
ypfP8vgqPd96nEOQVUTZGA==
`protect END_PROTECTED
