`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jdA1ebGmd5/Hxqmr+z+kSGl4Kib52rKKBuJrYmXFKlrXpJC56VQMFwXKIrRsDIhv
DcyUq7ypSCGNKS4IjxpADp6bIOWvT10LqG5LFsagvy4SwrYNa51F0CWwm3JfYqnK
eP6UeaVhNEI0cIJiKAJ4piKppQssHqQuggQwEobS31BbUgUsdn2z5MgQdC16qHtu
iJQLuFIbl16ZVBVI0IUbREegia4wcOhrcr8PJdxnBIovm0K8RZSSG81WgnwOphuT
82Sc/yCjzbxG6335HL5ocGINLzySC/AZM/Z4QLn+B6qRwBkuRAVtjIGn2Yzi2zzp
4VggID/3gFwUnMX1fad3Acv1nfHdMoxdlkcfPOhdVpt9z50pgx3YOX+zGY9nS3Mw
9+iimFKiIlVRnU5YDgvjzuAUxsE+GizFMT1TjXjrVd/gzN3Fb/S4dCqfsXAf6kSu
kylYW/MPVPPG+zckjyZ/WGgVg872jqHF+ByB4kQe+rZjKPgsRlPYggNWelzT+5yV
9+o+tzQxu8uVBXDQeIrSHYPf5lNfKlUUUWeX0TXVRvi49/SoTwFTZAjm86XmDGXI
xWucRWvErCTzl0hAX5iakX25fqbEa2N6LXGkTAlvdq88SdCLNqz9enahz9EFeNCv
1LjK5BEjO+RcaA36kgqZ5BD2iHgvxVjWxenL5/vZ+gp1RufWnXx+5NqmUyFGd08A
PuV35F4AeVb1cX81HBzvjnsnzBjf6pUU+FdXGms3oQrmFgMue5Pg7tRz8voL65L5
9HTTdyx/GTnSHBJroVMOgpWL2yuBdHvKHCT48EoDjuQga1NHClX2DjlVPQTfCu/c
S2aenuL/sPMygzK9uBaBQsiVeoyHodP6CY3iOaTqLLyjmyIBi8zHdN9P1fxLfh9R
u/bTJZnZ2iAOnaRjJh2hHG6H/a5oucLFf169XNp5AzQeUHLuW0HKTZaQmgMSYfkj
Z4JDmrV0ZooWqfcg633l7m9EDFJL1QckMNNbIIPP7BWxhFDdBmrL4sNnMfs480Hl
rcZCRtdHJPPs03uAVul2YIMw6t4Vio5Sc5R5sTPQvz093UPB1N9QDR2NOQGG0pLf
7cCeq18vNbSE2wrjYJ/ynhmzoDE9rS+K0VyleONXaRi+a9zD4SUEecyzteK3vDIN
m8oB7jCIW92NWRnDd/wG5h/FA+WeCf6fYzOiCfLUjUy+cbYaXFqqZicZPt+eedJy
MzsrQWCeB29P8+MzqIkuUfY9UvA4BzE4o/wWKyPEkiZ1nM2Cie3kjFXhfYuY4JhH
5U8mXMYzQtGgoY7QdKDRdIAKksmFeYC2mt06UQ2AS4BYugB7j7xY+ZhP4p9CKNGV
lJIwVsTf4fRO/HX5RNAFh3FQcj0/GL7J0BV6xLUn0wx1oFQRbqQXh6XeSK7uMI3M
e36ndE7zrU6mZJEFRQnhaW3wZ4P6ZmnbP2YODqP/6LgPVqhwQxloz1zA1AKTzMI7
y7ANFcTEDK3W9iPtqy7EFlMywZO1xRNzgw5+Ct3eKhrF4aYT0UCHuXrrrSUi4m6R
Fe3iKSXuIRO8rwewvFESZ3Ipo/lD5t2nWpQH6gOtA1JBWcjSSwKAD0kOrqNd9wlN
XvcgucK/reRNq3avHvsyZdtFjkDQzUv2ul3bOgde3Z2z2KIokxj94181/ExlJU06
Kxkjy4TriT/v68JBUpvLQ8Gvss97umWN5l9EbX7zq/WQcaYcoc0tHPHmNyVuJnxo
oSP8XhHjpIr84ZvVuAQxDpBZaCw21m4HhHcO1DvfqeRPtLyykExogy8I5crJYh24
kw0lTV2UvRsx8xvvtoy0vi7P5A51qxiu5CMKIqXL0BS3VBYGjyahaH/t6Xsph5VZ
nwbMSd/JI4CyzEixjM+SJnnZLDv1/M6/QHC2Owe3wJ5WlChgwVoY81FjFN1yAm/H
tAtRQNCbRT8vqaCvndSRjVfkKEIFdWrZPqtovkMgqqw5/YTXlMtprYJSL9c2ACBr
fcC0N3/mPQi21vbHthzfcqHD950uO9DPTW6X2Mo64ci6BkgS9twuTI8ohGIcD7nK
53bBRzaLVNJGd3lA+ojlsfqUwOLc0DlzFe0kin4QxO9TjVy2Z1zCtCDA54PgvL5g
51WxRF4ognKOHwGJV+9CF4jO0hlnhIIFPKDD8ewVfLfwuNrplQfPCxDMetQuo9rw
kXoSV3J6AIxkrcocoF9pHH68Lr/9CUh/xxJ1wiHgfrE4j6520oEmO4EprsWErXFL
wBM7fGOlukdEbKBWjzgNNVvrigjpsAVTUEa4xm0kLy3V2BQDhVcuq9WoW2s2BEmm
d+DGvzo50cYrCzdmTWg0rZ7an9GXAFSzXtYMD7xYNiQosyydmhY1wSxhH31/t+UN
OiYBSU5FkRaUvpCb87sGdREbQG233L/p5DgdfrigFQsOG354lusc1Ilc+V1HR/dJ
rXlX8fEQfV8p4J6slq/e6LWYx34RZ/AabuLhYXrrA+PZxRICGOzIVT4sn2f/ILEX
4M9tGxNS0ScIyYFNmg0s2iimqeD9AfIMsi3RqfE1FLyK7XnzIGqtUpnrHD8O+9Pq
/GJUie2HFqRQkDhpZVLpwVFYCaLVKYJKsn3g9Wp6GwIOsBeHcD+tTMbV68tusVf9
ptaf63bewIrHPxaJIc3Gxrar12wDg14v6PgLjv2JD0EreUu/jLVGrC4soBTllVdX
tqZhwJbBSD9Y53Ugm+yCMGMJHq0V1DmfP4WvQkkkwP6rc/FuTF80vMwOuD6TPVGj
09Tpf8xk5xzovOaWu4lgnxTLXvANkfyK9whY5IqxiNZPWkyU76Rh5YzkNdSRjJoX
yUGV7uomOxODr/Bsx2YSa4FKUewkx2d+WjuGFZAr2MTnqyLGLl8U4Rw/RaSw1D8t
wao2AFerary/2JOlNIwjIFo140hQRR0buN1RK0AEaajtJA3C6cCIx9gDUkhy1K/A
ZW/D0WS3BrKIyYJtGZDeVtCaI1TIzFwNsFj8rfx3UuuMBuFaG6EoPIp4FmrcqDFM
c0ERyXY10b1S3aoSpKvKfONfr7D6++m6Minww6ohGLy/4sljTPbXzIv5zCO71fkN
F2pvB/q5nOPsInp5v9HaM9dxinwkrc9KBgV4iH8ewCMt6/YqClJeBpEN0dEHFcbA
TgMv5Nvn0tziRIeqZ+t70G1lhrJhJfItf9UY+AJWxEgV4Z8BfRJcWe4Auiez4CyW
MkshBwDRtf5ecH/pqtSxEYoS4ResitXaASyP1gxzLXqBi4npsCCnn+jJvXz5Kr5b
noBmKlv5N6Z4Zf6WwGAi0HGwKqyxDGI4Ot/DUsh3jZ5EXSnYOeRGWI48TNcPViWQ
7y+y5TiG5jM2zhUCujfHL88yz84kT6Q55AdU/rzZQDPCbLj+n7FVyrhX1QEGKZQ5
DUCPCtrBa0hlRobaKuEqj9vTiJlsoeVDF3rQOgYk4Mx6B8GVAzph1DPjnRzGpPVk
xZAvSh1bvZ3e78x9lMAOiQEeAepn+I8+DIfBAMfVJ4vlO2jrihUJJCFb2uIBtz3v
y4Ne3Ir8a28DF3S4tojN5b1Gm9rpZAC3RDNFrz1fteW16aznsiK10VWoMyyTJbIc
PKkMXXg71LwVZq3AWOO3bAFMV8W4cKmgF8nVKYscXzwxN3DoSU2A9G0bou6hrqai
7lUTo8QG6r208F5KE1DrAOiC8sk8z/i1dSuQXlD92PtM+mcIzZ2dNOkEo1DZUlmE
t8VhNCY9fXEcjWPRf/dGnWH3Mq7y2DYZYga7SdYcPEVqaWKuo9xNnudTjAFOLJFx
sTdGeX31sJfzUiqochYhsJYurQv9vhiGmur/DcSnsR9/k8JZyZlBsIqYqz0hFm53
6spsIHN1I+RLRnjWVZ/kLqw7NS+BzROSqcBMEfSDPjYK8Pdq/VtGGs55NF66tfdW
qrVzdD9HD7S0YeAfu1RGEo2PINIbh9KHUSv9nLGZTMrpFtMGtE76+CvXhH6+XH8C
MxG617yFRtOcsXen52/akGtAilPluI5xQayc+vjtNPKAh4xgT8WH9WRf2HXJ39dt
d2VqTv7ChW1VHFH2FbI8Oz4V/1epou+/Scnv5xogrIO9WhMbCrfRwExAp5L3WGoF
DFmXHxyezHSx5dyFcttcb3IkRKOgHn1pB/OYc9p37nKBuygmkLO4Lsa1YOU16Njh
ntM1UuChjeyQ7aAk0DmVRv0JMR+KRngmQs8zoKZbbbnDAU9XJ5ih4/S+eUx5lruH
OX2iC2osFtwjbW6Fj0Cdoa8KnO5Cr4ruJprjX6tCQP4+dRsw2cutXL0XD0RjC/nJ
/M5SBp4kJb+ooWbGC6QuAXG+kphNA7yenthkQbPajoPl3tMK7RgvTYK7whxgeKxA
BDNci46HH/LAJPKL5CFv8Lt74l6vqQugb+/wZguO5UjpOXivuaxbG3gmZyrMg/Rd
Iy2rdQA1hYMwIWAaThQTvBgTK2dP3bcw/zdw7SNpqvQ4lEHrsJapT30bNEZAPgQk
l6FOFSLXlJWqkjYt9YTfV1KGBW3u1QyAA3Kseb7mfX6Gn8KOK9qszArzkz2qCHYp
4CEKDK872HWkq5GPfZe/KrFgkPxNolBECN5DgSarpmeNf+eey+Q+DtpniAAagx++
uy1nSJfPU0BK5Fr5e/rY3IZLtGTFVLQxqt2ttMdhXJox2v9Mm3Y2jpH0kWyKciRB
cFKfDzbgilmTMP2qIVa1XyHyZjnNn5b6Oo9Y6Na+7+8ndw3nz9SoF9OHdCxocfDn
PisZATgYRttMdr/cg2L/LfZOI2DX4WG/5NdHYmoKggD7Q6q/PH+smZDY6GIWYVEU
DL5BN11ruqirNUTQunVcNRcmkMG4gYGpUUYQdQQIXWxa+NIAfHCoMB6ufWleHyZx
i1JZrRXVWHuuzKnHGboqfIfVF0rxZ0RSnPMifwdzoHEh1+jEHORoX0TFxqPUVoEH
qhZmY4178R2L6Je6jgwBmupGPsTqZJXdk4LiW9WvqGEOYarLOl0UbtC4xLYxNCDE
FZBivXbpuViJ+IG9yeFAWttf9aULBzmU0th/lVnpn81kvHoRBiGxnvUe2FBevJ6H
gMhUU4PJvcSsQBsKfEDCKig8OMqDLuOiWIFwJPJlW38u6Ji2d+23IZEtAF4m2lwx
RnF3lH2cZd9sYwjJyLchqDB0xhTv54AQfQztsBd9Mv8No34qWJ3+k3E/jl2UIZhM
oEZGbwMHycKQwVHr/4c9DxynJbhC/9OeWmwBGqPyaX2UwcFO93ETPJms1RJobruC
Uw8Z+3emStc+kdDwHYPDZ27SLHebsUH3CRpBNy7BypK3EM4sV9eJIiuYrZV01FOm
x5fNUjJzRvHMdr6/RAzmndYTmkcHH8JdbKlNp4VT8bNOw5JqEhpRdDBaInAFK/oC
8g4widC5oaaHQ1uTEow0dmkkQ+ath8v3PwlYB5pHqJ1+QZgd3NEn61CW2tAuZA3r
WcV2L8qiZDAuzQnpU+Q2qgEJtDdSCq8F40gpCvULW6Xc/c99shlixcWLRy63knLp
/rrPuFWd321n64XmLoBeagHqdROZ3gQoQMTWfbmVXXaCsDGtaQKVtwbsYIALaTP5
qsw4iO/Ss/Qxx6Xtf5CGX4f2a8ZLKIxAWs5ka2J4TnlPiiDpjy3vTHrWpUsTgu7r
xLSaty9BIK3SqXrqGg3MnuqlAnsY0LOHXJSAwHPITFZ+7rmhB0vK/vDf3E8j+lUE
HCY9DjpzpyTM2fpX5KHrc4WIvk1FWfGscA4iJLwZz4mxk9Aoq93zL8OJmY49/9x+
xJ4DtdKgEcST+hOKZnXdoH6xyj1tcvq3qtLU3zdWdfikixttYN4LZYHSERuQTYh3
mWwfgRjvqY6wvxTBve7Wtv1UtX3iEy+nRikYdwV4onKG6q/xxR471hUcm2c4jd2N
UVzXbx4VL2+cVEOptXd8N6nf2C46UKQxQ9esh77SqFZAoAC4p9a23Pz6SMCcHqQj
aw3IsrRj6jpuINeS4erNX5MX3JgLH0Hn6i7mAoH+mEyWMfuf7oLp9+W243/IAJuy
wEgxKotWJeieBtmOp1m6P7q3TXjE854MVMZaZAgVKLpiFwW0rQs2doKzymchMJS/
kaBcnOra/BRSNhfmI7KArbuQesJKauLH+YJ5jzsFmBH0RtqKdWY8UcpplDo6JJpB
AErPm4GPZoH0mblxh+7uYOQjfCqAbGvPxKzlPjFVxTN29XGg/Npt/wloG9urs0xL
Ey+/7YlMMDvFyrjouwVt+FIDw6hEiscaLpEFIzcZ+hQ4ElNTy7bnGMuTBAzeZ6Uo
mYm8TzS0FHG4YVhqdhyKaEoPmrpPtW7Mx01Z2NH7m3hcxApJZcIOqlldfC5Ty2Mb
dLifwTmU5/25Fb07aHPWm5mV6c6uATeifEb5A4tJllmhUaR1s95YoOhzzO2saduJ
2GQuxzUWDb0Y/9sF52ORyYgmELmXaLdfNm89xOzm93oEiIQMMZp2cxnkj9zNrqrv
cgbTz5wPcAAx/3RexGpT8Cz2atbpDDKSSkOfx/0qyQzROtWRs/eHt6xcSRktmCnF
QFVzS8Nw0+1xq3SakuOL0nfRKe33Zkncc8Tn50Te22RUoGpL18RmwLANJm/7KXRj
gV1JxDnIKAls8KMOz8zT4jNvHHjDsiIRvZogswc2amr6nb1B5iX+eT7KJNvqLcwo
9re0Vk2qbgF7Y403LeHHvsCrqoKXm/vOLH/h/EvjlmTZ0C9JfyMXkuA7a99EvRvk
LThZSDfKU5bv4Kj8sm42kNp5XjPduAvq9UoqC/v0Lj/OaeEFnxRVTWvXlEdisYab
mZ/DJxGCYT/k5F565rXB6fGOELdTFjDYlmUkAx3wHHbcT74AvenqSiIkbBYuRuD2
mL32BXF1bKD+DnZAGtRa5Y0riKQwVnuX+MObEC4PC59nuZiIcky1J/qWkvi//l6T
xsIRmFeb8ryZGFOwikFCz+pqSGOuAdjAOH/J4N+/G0j+2jPwz7j80sJPlxvGMagH
YmPg99hJUn1UdXCYlV1m/n7h7FjRT7uiA50GHIEp107Xx6M/ezs7hE6inGgDJYgo
KHJrogGHsVPxOlN1qyBjL+7fOc0zHoldgbC1ZRMRsfqKW9cqbUvW+W9HWxZFtxf8
e2N4ge637mwkzZwqQ4odEDlyik7rNc/SoxcUF85kSwXtJWCpQ9Xy7QxSQ8wENAyb
xENqUQspQ0OxxsSnyNO2cILOJrVloSdqimWVcDtSkUozKyGzoMzZrRtwvQOf+P1B
qIAt2KgvwUvUUXSj3SVt9Ji7Sz0/uMRpAb0JzPCtJnNGWL7MMVuKVQDXwwYrGBH1
VK+ubG3rlJO3pld9wXnnC8ceI5rOiAE0yAPsvn8yZj58/mnZURSjLYSAmStYAzqm
DJD7YeMsPmpMIQKWAzwtQ4xC4eYp+u3KgN7SIdyoOGn5Fh6v24VV34Y0BwJC1aWj
84JlsvZ5xklWcKlv0S+QKBIVGTJZoQX8pIMs+RV2eUyatoG7elg6hqIu5vuxnooJ
nMwxVmz3rnlZs6/DEqRPFLS78ATA4ttAa0dYe5Ct1PXhjOvKoiFTq1xzfzK07JWh
2uMUbtM0ofYrmuJIue/8Bm4umGEnrJMNoctTvEWcfRiBXBc97xjW+cjdrYBjB5Ch
YNwqriPPGJ9T5mcQsLrA03cJqSJg4foMTh1of9+Xv/dQPlelppFQapfsW2MzxmKj
AwbhE+jJg7ToXaMTto3pGnOGqeyjd8kVj5Mvs1UXyLmf2Dztsvdx3o4m49YxE4aK
FDccCA4xDK4HJLiywqFqZvXSUPrm/WsJmuCURMLcn59MNPYe68kJZY1HBSJK3MvJ
HDXKcK72plui3dJX88gEVlY8Tli4CtZY7yoWiszj8F/6i8gl55VGZibK4NRCmPbZ
Ju/cchNa/yBqVn7O+Zxqcbx0CJ8mY4JmJZac3TA5BcTxXPuFpnvWxcFlSZRB+aWU
wgg6avc+HX96vhSem3UiO+StyrliJt7FhuGhp/dCGbSme2rUzzVeZ8k/KA8IZv5J
B3osY6L39FIMTZKEz4sRB9tUq4k4UhJXh8bP6KysKgTDFtxBSyejyQSbF+Lu/f2f
K3zp3G9j7lbYbw7AuX/s9P7XrW9Khed14lZER32QYsxXSIUxBolYIIBo+AsQzitq
V1LeAWnCGN45tUdGQOWvy6zMLpf0YK4aon8NN9z6nEV2XEG/eF0iVXBi9c4/QWkj
Jf/6yFB71I5/oidtnL3lH3EM73X7WFiOzGotVMbPcu7iqOFz/o02in7hjk4ScoRI
GvsOUoTzExSulIdrNBPRc1D7sCGPucojy79CsSL/YZlyurzBlNkVZZBUJEtrNGaA
oxkumibNPcts9cNVr8P3CWu3pbcpJUQR51nWUVl5C8Qhw4HZpe8qgsMMd78+qfhG
UAnWtoAV1rpoeyVZ/hEqzmAMKK8qf6DRWJ+vF0vJ3XrvUd1q07EbMV7m5p+l3bxu
PrkW7zrk8LpvPTDgu5X6gAfPeTAtnzLnXkHuR6j+yHkU3NUxcH4Wb377Bb0CAVlH
Dgb5db7QjVFO4bkBuY6yCya03/XTKOGgUaJmAA6KYupDFt4jnUyzXXZPDbN0fbBo
Yc++AGs3lA1liAn1wvKD+IOJbtXuSggZYXD9RcX8nFA5V3yAYqbCWcisCCWBzMsA
8lpHn6ApYwYlHiwBcWj9ONEg2MVZ4AJrUATxgYMbas3yV/23hBVxtiv04A971UTU
pcTgpRlxEnAhUsP8PEIDbHFsWMPlnw3WK5/gZJRLXGuempEX2sCXmG2OrMGDkSPY
2FdXgyRSMTsI1e4k5d+fENTytFHuRWPnQamyorZjoppj4VkxIuAdNNnlfodNQPtK
+GAGhYXZi2kROrKCRBoE4TX/9WOiXYbpifXWLKm9MZErecXeckizXmWG0xPX9C3f
2jSUSf0MNwLjFCD2INDHed+5mBnr3ntTj3anB6WmgRIcqzydh+jh0SjlzU8NSK/O
jvoqy/uHBKK+OrAIaQ9HdaHlNvj5PxbeWoOuNiYbOO5xuGJa56CYxS1uvKo9Rm2J
Cufv8+faOsSBXPtZvRx6BJMJ7hnpnKuEtz9MCUPhnvPNZsSq+Reiho3JbgU0MsnC
jb34QrkUdKO/xId9DDAawiW/DqBSyMMhkFTofHNTNq1Reh5i0/f6Ir7Ism6SI1wj
50jRfFkGb8GvgQHCQayVFouPLgfJkJE3EZa2T5Xl8/AwSSpHG1e+8/PlmGz1lkLx
1dC1wTnYYipfVpqtYZPPGsD5thBlc4R9FkK4JY4FNAHl44wiWXNWBnddc1/K/hmT
So9D1vpN/0Ec3+0OvI1eWubvK6bnxxhFS/prZp1vE8TFnzZQO1EM0mKFL/Oa6R9h
9mipdCU/yvVVJ/TUP70XAH9XdHN7EYMD9gBwZBtsYfK6PIyVPf+M+KxH52l60A7l
6m72L31OnqFH83QQY8Xe8uN7YF2ZseWcXmBjbT6kIzBnKgLbFmC+Nj/ErzK3f+jh
w/QotI/cotj9yAWoc36bSTZNGqcIk/UxZXKhUmwheC2IZWxwynlqILnS6LL9mOhv
mT/TsIYL0b5vO9xTJj4rxwHYe0/IHzC8GMsDY3pJpCdRQsqwq0xPse0bE53batlA
IkYb8fUMjfeTXTZiZgfp0oMQhBgam6GJCl9o1aYP5QtJajIVw/s3UCAP0PsX88lC
ZPFnrsCBff34ML7NtJzG38nH6Y+zh3P0TErl4QzzeKKLRkIWKe1ZrlIZLCZaUZCg
hpBa+WLFXw7btlrjkovfAuad1Zjxicte6iajOYp+LOhyR555021MhcRp/Hf23z5Q
+ktMAkTuZkO2S/yVrMeT3AZe8GsxXQBRCPAtmId/D88V14SeGcYukD2ncnWyxJYU
nMEf3GAVov69XX9engJbXxRPgTUw1SAsLlaqBr3sVQOc/mVn3K06NMq0ZyZNYArb
7YPZR74VGgxHxrArYfvPH5mWNagjYQ0NlA3SfGgSbe/AvKDnIkpWcrgdScGtjJeS
AhjisrBSUwV7YFZPE6xcR+tMkVdMnqpP0KvDyoOQ5sVC7YJvjKB1EHAzLTETLMk8
GsVHqGo53BB1WXenFoNflHsx3tas1Dkd8NN8kpNTVMDWBWIpLsVcsd2JNlhAf6QW
5Q3T8H9CBcQXSv5y1qnVG/BuE5HsHZhOi9M+D58kvA0EcqnQCZBArP6vruIEfdHD
t9pfWmMxzu03SnwlbxwmdtTFFdzchUgEF74Llz3Wt8MFB/X7FfPR0IrENswFz3a3
m/xv5Nd6JtsIWfvOCDlz/wp/6JZypmfHpz5DvZIBb9t+/v37UJVaD7RwgpP/le2c
WsXybmxVenINzV0cRvgWiMdQkH/x9l4PWbZEgBxVgSlrOZH/56C76jiQ+ZaxeYYl
MHFZi/8YqJsg/y9LYNzAiIG5Qi9EPObfr8OzRdbtal87AEb1nXGcqfNWB4VmNKC0
x3UhumvlxmPwrWq/9DaqFL6+UJFHOVtnaQX4OuK8UkB+6EdIW668xwz16RcFxPb+
9De5JvGg3zncX2F+514HiImtFHVvUDXX8Nl3tQa2Qe5LkldHSr2xElgxBT3iKVQF
iQ578GZNK9+HX1Lb/oT4wdDrty5f2Yigf6i49j0ST4mjCRynSibymNNUEG7hxt9T
Wb/bzT0Y++rMKEIEdNA39Hfa+UTboZ4bPa25MUDXeWwQFAULFuU8mh4ABYHAtyaz
BezZurjyk6/IJOHGEVU81UyYIf4yjyIM2pVQM9O6X+zFv+0T87/UPswaZks8KjhE
fxW3osCYaqNxBe6d4/f9+Bu7DG/GaVTYTgIQYfeUBiN0DkpTuFyEDC2qSnCGOGFP
XTiUNgd+Vxbm9ffERVcrSBwQU4uE+j/J9ISDQCIgqk3OcKmMkenAze+nNuPs1Lmk
2zmlzg6Ux0K7eVlrElkNmrO0lxkYG7JhsO1kPgdbPXrjFVj8XbFH8N/m3qmWplh2
uGDuXQuMONaZ18oO7TrJyd47UtdEPsk+pXTQo/pX/NrTuNXQmYueWtZGm9BQeUyu
2VAqtzWCbEJa6jlidsPbhhpoVY7a5if92K1kMjeXC3Y2gSsGwJRCONsIOXwru84s
YS8rGs7sYXQkgzXnAgekD+cnKpowRg+7Y5V2Clh1dtclze5RJO+N7wG9D2hBrfxM
odXjM/J2uZBBFhci+0xVsQc8IdvTLO+KBNM1Gn2ZM3NHX+dHdo7ZZ9tQ1IG/pLiu
vmYx7Co3ET+C/cn4XdoRLN+nocoOewArBVodY9w0NFrrfbmDGItOJvjE35rh/QYC
533usCoIQYHvp8Y0zjUK4dbJULc1kEa3teAUf0+dTomhoQW/Jf/LLWfwIr+LHeIY
BlpR6ZaV9SgFcBKgYc0deFM+uSJB42nLJY9FkMDlCCN70yxpYI9uJIo5wjK3WUxY
sD20n/i/BG70F5BXLwOmUAxMqJt39c5L7aWQvu2Z5yt59QKFGcw3f6lro8VOjIFJ
Px8ERlP++nKUGm9Kph5wF7LHjHkVIbQxXvycLTL/9jhkKI1BgXPlBdhMpYgBjmuu
UbtS4m9oyzkaGLyGEZf21IaXBZO+HhbsSYfHvoXTtLemctGwKIsQNWtOMt/7gn36
gW35XxzSbiGDatiwZDYMZwS0fytPDzTDqIMBYCeE7RT0g5Ljfo5QYjOjTdCm4fcN
oia/E6C89M9xnz4JU2llIrW7W0iL7X+Nnv4bJhEA3pTd0cuif+9TUPMzMwfiAzvV
SuqfKS5AaZh2pgDPNj3/64LtAeF1PueymM6DmDR++oNWMmypHZe31kPxXQr+Iyj0
hUNqkyBlYptMvz5gm1RWfEIzbYvJMeyMMUtZGzRFIO8VUcsKlfibn8nP1/oLdZ3T
iyjP3Nv8xBP3xsN4IQdkf9vJYyKNJhJfoMW79qlfBbaYIUKhybgVnCfdGYvGzbcV
36FHGlU4DkGasNCYDPlVuI6zgVzjiQQwiTB1/8Sz79R2wDR9uSID2WQrVLR7oQDx
kFHfO9MavOdYDh4Z7aeNljCG6d4S5fWWn5H+wsn5PHA/j4EaDq9OKZZfiq8OGFJs
IoODTOyD3zHYOIPYhmdFmxvNrBBgx5ZvPKRx7PVlVdnCF54S4uuIvDuBOoqOKub4
qPE1wens4/1/D3z/jqpZeewgQnNiiNbJ1AMiOJNqc4GHGWg0X4kPPteI5E+ljC1j
3QXw8lgvwmYAkTXqGlhJa2QsNI0XUs1yfgVuNFjqAtt0712bfcmJklrBhkVIg3Xr
wPAFk3Vbsp8RvYdS0lRQjmTvViuNVMfqgE27QgedyiEtYa372P6tDHYlweDhg3b7
duedfeASi43xIyoLoHoeJKaDpKHICH8Sk6jd8/dAZ+mzEEvAylVhJtCmyg5IFI4H
6lGNe+A56nPJClh5f3khsNiy05cNuAjfCE6026QHG/k08i4ZwV3DCqtaiFH2neTT
uhYJ7KFCiL4QmjuR+SVkERTYDi3ya6J8I4pJkQXe4xU1FsUnt345rrURWiHY4H8j
+PzZOibxCMQb/AnEREi65d+RoN7AafNIQmcyLOz0MoIQrvEBmRLsur1edBq7dHhF
8PYlLwc0bUOb/YiFFY65p2pzMP1aCd+nKKn4K274CmjBNMxxE/xxTSeDZdlCczpd
7o0VaJ+Tm017sw9qE0cfaiEElEdu9Cd9RuxcR2xYt7Ji1Fs7W+KJet2DBhc2syef
zdQlsyHzMlk2CYN4/0ck6kmai4RrAuFAkNL2Qt5/3LTwr4rnQP5jWo7/wmzlhmlf
i/512I09w5m4oAPvSHiZMbg5X8V7jM2D8amidI8xY4deESJROsDHfdkHOGeigJl5
Bdj49HzvnPbeUpb3ajSNCmzCqbrFJlLRt/Dhj72BkRZfM7mVNIXzMplAJ9uoWvCj
D4RYggrkszMelo6gstz7lbjJ5PUqU16Xqyh7F4X6Nw+TdYwWBVITZBsXjcojyj1E
0A1014+nmWbBOI41uIl+ZpsswoOyQjoDqAKLIwWMqzu/ceICZBCrOrkiiXTp1Fvg
Q9jmDNasPtfh/ZGZJIHLAAHRa+p48ijAdkh7HffQS/TCj6gU302bYDZc2jDL6mSY
rkn3un1JKTDLdubQwU/XH5OGFnBIrVN9GGolTYMXPCUeUxksjH9XFO3ykfTD1vOW
i2jk50HCwOnAN5LhiJ344MS+XpsfEbOQqzO3VarV0b5zo9bSUdIZkXloDJfn8MGK
zHcHnG5akAsMIWCF6GIJTcZQnkU3tqxSI5fAI57akhJ/SYSTeEjnpsPVnymGgFH4
KLRL0UKwRa9wVllCFpJL/fCXzVf7LYr+Hbn8mYFkKn21ITtULA5Unx8z2OGLRpzH
r7zCgY8+NUbvYz1hzC6VplUc7lFsBydNV81bHLE7RsChpTeN8JF19xcov8ULDVf/
2M+dUU8a4W7uSwaXQFzl6nekWY4oK0VM07N/MhLNc7OFccM47mlxm91flvM7G33X
r4VcGf/u06Vl5hlFnJI1pCSzgbKABEP5Pch0BUBOzU4nuouoHH3Ldinf4GJ5fFvc
uUv/+baT/cQvY3DR7UfgtCqwoJhuJHawziybCQ6JhClKd3qCsPQAYSCVyyKDwQ3l
KWAUzYD9Kf+S4kL+14b3JuB+7XVhMgAqCIaFPw/kr9PF00r3ASn65aRQ4nxaM8Yi
3ZEuA4bJm0gnTGsL+2B9ZJal05hMtJgV3rirm/jqcJg+mrdQbMtUVTUFRsmDnOw+
3CnHYpfiJT5Zxf8o/5qgpjI6SWdmpm8xCBTceURhtvar3qdGASBDxVyy5N6I2qrA
sVa7WX6nr4c5yeZq9QIrMUt62KC3Uhw6t3uH9W4CuMEyRX+x9JJprfJuxEfaQ78Z
OkWHCZxIaiy/+A8PBGHah/or9Vb+hOD1hqKCeLwMbNE96ZRd04HJ01RbLDsykCcJ
C7khQCJxTaLMhT5GXRVZ01RILFh1NVweRYBO/eppgujEIZljO1f84xvbG5e1XDJ8
eqagGi4sF5Qh918MFdZjU069cR+RsOJl6aK55I3Sy+8naNgDcdrg/gfVM/4GDaex
uczN2tjdjg4FPvZP9hU+9gWCuacX1HaTTNYU+3Nui+OO8cxJrOTXzbRh40MB9tez
O/FnsFwGBPjBT+DLEnjI4I3OzJlQq+QCLdD7p8gyuPHOqgkUiq1j36DarBbjoP2d
Bq6VhDucMgSa1rMjVmgyEme5kgTzM+tkVDa5PuLk0bB+L2tg/naRe9X9Ib3W1Cqi
De/6ZdtDYB8m5I0Y3fLHxOAyylbonovDL9T8hPM5BiRFcJBu6uPsg1V9xRx9LMrS
r9wSbof5KgH2e2br6XnRBA+yrFrIXdpBpQVmJ1c3SvIbZbVNMTWescO83UA6GREs
RWFgeqlGXopb/i4cY7YHUKCn6g+3IMX3rUKPsuaj5C/Y4T9D8tprPTWT9Yj+D4nt
TQu885IfMoY7Rneti3RIegS1agKYXm3RaM2z1rtjyrAcEUsKAPAzVya8Yj33+H8X
2V7iLLHy8QQ8gByys3O7W9pMRWxdov2x7P2bj3Aya/bBRryOd2NcwVuy7aQO3FKb
po99nE23KBeKbRQajbu8QSelBeCjv1dRS3fdSTEbvCUuCQbvZRNTUl8fTT42f8tP
PrKyGA/mtBpuW3ldgJgd7nsZl/nZ7Xb7HrozO0Di838SAbrFNS/eBYAf22fUhbAM
O/5gJUQa8ujI24ZmyBvqjrZb9cP8zgVoKorpIdhvYIHIdxt/ib/qdLe8t2DAtYdO
3Af4BEnqep7bT0cuFCvilOcvPN5YZ/uMK9n7jvQGRPLW1o03RlrJq4XDCq+hA6r/
qL7LbORpMf/6geJtlfDv/Y2yXNauxQZ6JC+VXwWJiW4z7vH9xIEg+w8U2AQ4oPwY
kOiFo4750rkMyZlj0rn5BXiRusfEwBJEQQxJ6LG+9Yj+0ViyaJaT8QmbMuwA0b1E
ncDY25zpvvY5jorIOribRjAT8OwrOO5OVK/YKjo5pqIzjtNZVtXOxqJyz/NgBm8P
rgZEUuv6OUo2C01cTurT0OPckLtdBk5kY3TGUwnNk9nqwYeFAdL/CdCajFzcOBx0
xTJdkWy9awxk/E+5pYJUUwkF0jAI017uIlQzOJwepnB08LazThMlwNWyE+dDR1a7
pvbEVHY4iKoq8sf4KrQSgHfMr17wFZ4Gk21h9hV2x/tE7e1EOBUMzYhOUWhVnHtO
Vwg5NpSuVoxBu/xLofjJDsGjmY+P5ZDA9HdUMinxMJZzm667Ma/UPyz4yStKSbNV
H3IHnMv7wwPlh4zLZrmJxojU8/4b1rO+2+7N5XkxG1UPGZBxiZ7wugfds6zl5qzD
HqpQ33Z4pZJ0CgZu306/dMVwlx5QV2DnGpU7ifqEJNsBhoWb18dj+H5pQwN08UzO
XIQSB4xt+PCi9fXKUmFDVXGGj1l7ve5bn1UdS11weGkPvh/pp8buJxYelmmr9tlz
Ta6LoEsQlSy30yX6FF2igrDIdjFU/b6gX4oQRWyHabvht2zXu1+NQlJhb/s4K/I/
pd2t+7PxhC7uqyXppvMdHTD2Mjql4BSIAwbV19GC4Y5R0aW34mCKUFbOEgGYVQYx
Amp4srkY6Io69kGxbOS/Pyaje81TfoNxF2f1Gu8qr1I9x+ex+4HdPeqyMwYXQcTD
J3aW9V+DQn3YPZYa6BEoV8orUYSOmHDm3aAqKwdbtFbMKYM15Xvh02ga4ZVOmoT7
oLv1jZ98uWN2vEKKvNRa8LmozBVEKuL24xa2/xT02memb7dywd/0gg5dbPSBjis0
hMunHytXvKLd1oc6FZdEUtbIDXP/UP0nzZ2wlCOH2/xVlu8RgxYTaG8ylXMj4nS4
PK13Wue9P07Vd7UH4g6ZPaZYO1u2ORZUZpSzNhGolbumkqGSLU1K9pnEOY3GVdYr
YDEuoFtZbOmWGfF0cUmM3HiEVpBDVnwmibx2ZGyO9naxoPbopa7zc7Lz8sPorfzR
WmsvccZhak2Wkv2Xlb1WsOTch/bKG9Bz24gPIFnVdPurOqV77fKbwKlLeEt98UZ1
P09vVfdQslWkMjcMHcIOgikACbP8OcaSxm+Y3sLBgldvMPGbIhvz1Po7LQ9zPoTu
Rlp5QJAhgBemcLxXW9z5JD0pGj59a9flMd9rpZVuquYs3oNr1CPYL8JEqWZNGGVf
0yTW0Q7EO8fl8gTQwHtf0Vx2XNhjQPHCOig0wDReMa5V8O9rxJqnqOAO3VpzOSgW
0b3lBrcf/6cO4ya+zZWEgFlKQ09VWt7wcjpb5MJRaBwipVWpXdZ4+efKQo6UcarW
UWKpl4x+QqE4evE+NRcF9VcRQ5AbsSyIVnjh31KRg6eZpWvaL8ieD4pnmsI7sCk+
A8PKvuI4QO5NPmlSCstD9KzJikl8n+GsZXq0vRhUzzNfxacGOcfLiCkbbWilNoWO
lAgY8NvjtdA97/vmRtYb93hUMwv21PJq/IOkZx/CySF6s2NeA3ONQs3UXK54jx+Q
sMQWZGYbVHzs+J6Z/DALvBuGE1Vq0OwlSz13syX6M+hRyYP3YciKfpkAPVWMn4ap
lUDaYAVmV4I9nGk2ixYgRR3GphRv+/1LozODoKVMoOgex8BbFXONRUousqw2Trk7
6SFByct3GlJwrLpWdisHhNaLqFUwy5F6VahJ/hnT3LpLCky1kcEierwFp23vWd51
f4DmTeAb+lOo65fRvzx/4h76yLlkPykuMMwC4OWk0EV8nuiuN/3WA15YM3TOc0nK
5vgxv82yksUJ11fbHAWWaXeU94qolLc4Mmng4qG+7aTAh4dFIwJWxKVdVoKzWKOd
78TKa0AKVvHrtAzrOCQba0V7zyAvVW540XwvFWQIG2smvrwDLAw+PGet3xnEnTpB
N2X68KACR5NRnHmQYhZ1ATvQGzAon2r1QITcJlCjrEsxdP5Vh+nlUi581SPg1ppH
FsUeZvLK3M3Odsep1BWOBLXdYq2xnSnvzbF0FHJ1I5anIIe653JTNuHu2QGeNu7R
WFFbcDjM8EUOqrpcjKMp3xP2MndfRzVyhvSDfPuwCD+8nwOcmBhi599W+3lhhkby
zloDP9y3mR8VR4Wyrn9N5F1FE3q49Bw4ROshjoleL48Z1Gsw+WdHPj4pw0KaguZo
C8AUoPx8Wp3FILFr9ORpyG7Xd4M80uXl+WCIGLMuUwg/Bey6yw6iI0sSO17nP1Dq
mV2odVWu/lxoGQtVJpmahuQBWI4vc3c++8AA7bMGmvEETHUBeAcS4xWvTFo4P1K1
cCCgOPZ9uyYJuhZaogmBRvQT8uGK8HYe2Fcsivi74NqlTDVkBwkGuOHkPj3YMAPX
SWBeG/KjT7xAAZr312pS58S3egUCe+MqE0Q8pAioK1/pIdgwm5IKheVtscXpSbKh
XSn9D/Q3vXcnPADzTKblGVLftRMlYYaQ/IUJppE8yGHxZJSpPkiMW5KKAOclFmzk
3PShmkSIM8qaXBt68UQBzGK9rGL62LWDQXc0u9Kq+zV+HL4+BmO17sihAxD3icVn
LJOKRP0wr9DTBVKjL9GoeRABpozF4dGqR9e/BSGncoNSljIsCt2ieWKMitZqxG8w
a/nrCb0KQu+S9rpb6mqxTPYqdv3ezIEMUqi6c1kWM+YJjgYAAjUhti1rYHRWMo1v
xjijKv31kYJltQH3mSb5UCgVKClL00Cbjg7gpl0b7EkekctmetwV7987b/OmRBJH
4xI1C4ghBG3iuXIZDOaMkRU79l2nubxnI2WUXuIBR0Lpn1G8sXMAHjDO6B+mHJP1
LojS2Ot0Vt+pcdzc6JJgHLpOwxl7jnnKoLmh+wwQQ/RS12YCe1HMD0P7EpClcEDA
wszndIQkVwiaXd6z76v8Wxs2vyHdwTpm883HMZ9hyVNIaVlJJ1/uYnqY3kRed1wC
YW0tQId39yI8jos/7Vq3k1zAX3dsKpCntgCXxEhgvnfghHZniKG61yYSLoB29Lag
A/EPQHXOu+SroEP1asRJ9TQHyyti3xgmBnE4Rn7CV6vtqlQc6gz5ane8GrpUY8Zc
2zE/QrJiszwr413u42YAJLzmL7ywX7JRZiSmEj8qmmCzEe4IKRRC9XFLcrgiO0eU
e68Tmh8VPUV85+hWuC8o/sL+ATQ3UXWPJILmngYjK6URl4httu9OfGSb4FCmMlM8
ZVvWvx3p+8LVEkoEijbaFbKqi8z0TTPeM++TISlvfLUvp7iYZE7ZodWa5+cXg3nh
BQnPC9A/Ln4DpJSA2qPwlSCQop1LFVLM80Pv5PFlAlRuEtTMIClNNysi0znIgQoD
eM+z62XxOAJdb2JzA33UvxOsQRAJTb1F+CZ1Q254n1PQDtLZxkDC9FR36MlavrXX
fxvqHbGhxFVz2QnDMSbYY9BbcV0A7IRCxeEaWqOKOAtI5/iAXRuuqw+lYvOf+GHE
kJcgZid6zwvTqPufizkucfLLLmo77E5N4SqmWmTuzyBu02yJ3YcKlCiT5mY9rLRT
paoKAX1T0/cnzoU7M+sjpe1kX1LYkBSe2glogtvqvo66T+EvOASCLhGs1y6N515h
i+1X6j0D4CCM+JSwdmyuSbhRGpINmGkQCAR0NgS0P0nMo2512az/KbepTzFTZkfa
tJsHZBfOUbmmL1rqJdPp/ZFcDoj/iGNIKz2tZ8qCl1njRtO/Xlo2h23C3/Ya8YId
VbRyFIi7AltoyBYRiWThePIqywuuYvOlHmNy+CcOt0bUSGlyZ15hNs1+brTUv2i2
lsGCNFXVtSuE1bnNhRQCbphLKfu/MOIozUa2rLF5uegi+gbtdkN89Qn4Fu3P+PFu
5QGwDGPHgoUWB+4icpw+HJVOi5OknqsKhjD9WQgfMN4ZZW2v9u00f9vfefhEvg5A
Kcy2yzvYgRWNmuKk1DJWM4zha2mkAajb43JUs+/+S+MUAIl+eqO6zNb7lTMziu5M
9TPVo1P8FIuv27TEojaSN7MpK5wRSIfy7S9GrcrP1l7kUw2Iii5gMP/QdI7wuCHi
AckRSULg0f7gyaIZa5KGzwEU+5sqq7gna8WZU2BjPl1HOZJMw9TWRCpVBURbZ0dN
iwVHTTqHtjLLD/agmShF0T+T/jW0YecqZGkCVszQurwo+hj20ufiIMjD8aJJQZP3
yjez32zDv97ZAoVwFbFx+cTfaONGEj/htvCTF4UgSn4l7DK0Zx83zoEJQtQ0Kc3W
tp/qUVfD4qvVhGzcygh6u2OkxtSnpiTn7+MHEs1x7pu36Qu8F4dC8+Yba1dM+5WY
tzzbqfcWz03XKAEscBSXpFCFgF4paqdLnwBTwcQDr3Ppr5mzhSHdqTb8XwI9EIAV
uWmBu2qkBUjb4uxuniPUxj5vc1JHE3a0tSX4V1Y8QAq8vUyekDWRDd8TUxrT4Epi
KAIVflpmrFbKXHZWn9rqs++bQMoyPSls3fkHt+0ONleFOYzJ2sXbL77wU0AloaQR
94cQ0fxMs2K1llgHhSeL8wdcdgilKv+HaZsuLziENirOOjZkB+BCkdn0FGFsk/TQ
d53v4lTBL62Tnmpr9O8ybS0m68B5aQ4swwO+wD1Iukz686Z/bI2Ptu3/xOCAdGRZ
Y++R4AcP12tCHtBz1nU3v0cCG4E/UzAvDYoTWjQXIHJCevppkgdoKpYGgLve8JJv
WasHQmxiuZShrPyMlPQv+ZkwL8tiX4T8ZSU0pHL6mVw+zk7kgWGdxJc1dgQaWCbH
g5IK7B0SPzHmgI9YLpD2VUtO5FTIqHDla7tBF/GphJhmfFOzihdch8KNSYryvaeH
i/xhA00c9mhJKtUEWHxvYTD0FFniQMSpGjyb9GgKIAfF6zDKw/isGoPYs2UKLViK
XZa/VqT5Ec1voAh1Y4BDo3GV4tsNu+zW9hxYsvDtScQzH7F4M+RS+mNh7ugli1cj
WlYnd5QCOW6EBRsjMJjtH+F/XCHkzGP7ZiZayVa0lccVl3v7MCJJT20JH5FcE8vQ
MZXT49nh3SHvhBYYQhzzvQwVk4QKMdvgjSydBW1iAZvTDlmXq2geE3W1MdWvAZ4c
GlJRkYTZNhbPcLo85OXk05VDTpbQlOaKT9yPCStwr5Jv1w/Et3qtgDQ6HdUFT8Mq
52N8MfN+MmXlbupWSoArVibQNB/bP8FkmKesB7yjlKotlkHmTa2R4m7USDB6oGgz
v7fEl50CEV0YFvGvycHaX8NA8c2fThU5iPkFcQJFesccZXdey9/j7jn/MtS9MN5t
ZUi1KK9mX6Cz0pVJCUZ0lpgSDStCIGqJFAlAjRfMfVe+MpOKSpR36BqzCtJFVIby
4AvvYB9FgFzZBCN8kS1bwqcGzHg8/2x8R+pvvlXpIczq1RhT0k8PsgGEEevysVSq
S89kFlnhM1ueKDR+o9//2hsIlW8J6QUEGXd0RmeGvqyBAT++8fS6mQOxkCREJ1z8
b/Q5+R96I/vQdNtVUaib55YXKF2S6ZOIa44+VnUBJJ3aT2iCRkmTDbe3veZ9sI+O
0z4MgKrrz8+pn0b0J5SJz4IDu/fX4Do/bc+hyrw+gbQG8LxnP0Ru+oafz6XLxYvP
igUSca+AWnz+BivRq6nEUZUqT/tTnacVZgZwCl7tiM4qi0/L9W8TD+Ep1TU28y2v
rm8I6mVoDxskoDbkKNV3jB4Q2ZHUguyv7aAhA7/uLfcppVpzYQ1i+vNxxc70VWQs
ydUGNL4jEIhdj35UAniWMP/xWqo3H+KMNUZ0M36hSt7nrU01qppn1vcfOKTXg35+
+9ArFgeUm6m6WNpCyZ67AJFDv5vZUqPMHCUllE6oeJks5+Wgf/KTwzhvZdikeH1M
MDqSAVyYMX2JctyE7096DZaDfPZu5uPIiKdzU+ALt1tkzz/MOnVYoDNFRY6XSh3b
qz0vNF+i1XEMR9EF3cMNQDgdpCZZ/Y0scmqRocmA0jtSLm6N3KLEPk738+mVyk4H
tQeAsyCFzB071oSs5dCf/syVmmJHSg4ioiCdNUPWlrdmzLriK8u8yLe5/nDoYV76
P3E6GoMEnQ3OqooqOvZOpKC/y/eQqOpb9s5N9XhyOXwwkcOJ2Dfz/3l/DNmJdRry
lrXvKS4D6yEanTugjp8GUIDK64FiYpZkcAz5URn8mfot1HBPQX9ZfmCXMSnJuZn9
eKhQwE1bTVjdsh0eMFHyl2jiSe+k1eweI9hP6UgLI9wLhaXoazKn98Ri4PKJRNCt
VpfUB0h795ESA/Phh/AqOPe5P00L0rfdd7cO/lWtwhkOCcKunno10RysbNg/v1Ke
RzaNpE63hnfHi30kEzsJRLi98rZUQehpEDaTaMa8B2FFS9zS41JcjmqwrL0zc24V
E+EkDMgH78mlXWv+ylL7hJy/2w0T42vGWT2uNEtaHGjz0cNx4U9k1Oitm1cYgeE/
cwP3mTza1Y9tgNXUBsudIttVKgqgnUbqGQfK1ILA8OFgA85zfiNue5bQuooR7vnF
NONsXAfZW8LGg3XT9YnQyRIadq1XNKhx9gsYr3c8R88n+xwR3tvNqURUdkzMZAPR
yMNhS/POdAKOD8gk2zu00XLpds6sBkOkIwfaTGgE21PEAgMSfPW2tenfGe6IvZSI
ijbTb86WKerF4XXTxQZD5AQPnNoaRFQwmbjW/p9ultl07qghEDNQS60LyGi+iefH
CSPsNbXyGK14vCqRVnI0bseBpPgQNIIGKXSO5lg+mhApHbYlO/p5mzzFQQ4cUUj8
OXVKVU50EoMYWzDLivKFtnFGErbo7f4PebU6LFW80qKinUdDjrauKTqo8SM48s/G
dGeayzZgcAfLtDydIUqY4RhWdQ/BuVzO/aEiFyjt8rbWN55KWQP1TxUO0ZUL9Aye
sJCs7x+PqeVl/GjIbBz773iWZXzxBRjHet9dHTGVJ9DUoR8N2E/1jRWLstfGPqqJ
mBztTStKrND+D3bUCeyULsFtiShs8KBA+SYdOGeU/qbTMnKM29sRbELogQOjg3uk
lPSKl5nunNPaZ67EYOonDZZQ17ywGWj74h//jjiejzqzZHVKqRGE6b0cmQ12eMRC
Piq3+MIcY55SlrjSC2w1oixnd+42ZiK9yS8ZD+z74Gib5BYzbt0oRqEMWURlL7Jw
vQEY+GOrFoRMZq85SKLa0RFZuaJc57ulJfUOxo6/R88bJmZYJ2iozYdvDKJeLWx2
wyh0jZG2oe3LFObP31kpd5xODEhY5XPqljU/tJEKgC4iMxgrjg9j4BAtEixDTQjC
bbSftWbNxkXtnL2iaTe5yxskx8lfrBxcVJchWIU5ucZiG4aGNMInY0T3c9lGmG2R
R9Y05XzP/d5KnzYAjPV+SNQxwoYNs7le6vyr9w6QyTGgGn/XGqxF/QgWB8caJ8Zy
JNcFhjmFoO9xzxzTgW0z1fzRMxXEdbIQdK5xdxc6nl7dx4rmxoao7ilOZMbTmt9k
dtdaDQr75VeXbDrdli2FWsg0BYov/Ty7AJVYHVMYGZRCMovVVqPCDHduTgcrdI2F
hlyBJ95tH+fhkhqmmvuc6bm/envgT73a2amYbr0gtCVMJiFAlCfrXNzGzuqCbD/f
sZrO8dcUS6awljjcC/xNneEVPyqi2438GHsSh96isugR/cyWqGVP4MnI7JsLFgqq
HPZrtEYHqthxUK6xr2TL6unRtCCqdFe676wjMD/FV5euCC8aiO51QPwnX3n4AVPw
wMq1lhqPN7DSJ5e9FU2ZZxHWWRZj5VHBbkn6X04UXI5XEejK9eGKRh8fTwvlij4y
OrKtcCfPW1vuXPDq5T0K/u9Ja/EkSgPyl/sLhz7nTpXJqVxEuPM1ieFgxd0s1WOG
wtn0muCQEqV0e7qsv1jW21iCPKhfwX5ntY9SOgbRTW0JG+5jvvcOitUM5xSaOxsQ
uArz4wA0kUkASfoUGwjW5wIzXhZT2sMCQ4uonLP8Vurt7Hd0EiNNaSXB2OX/a22u
dDvjXiPWYf2XVjd2fzi0TmYGLtaUEuYFuAsqPI7aenwznGeHXd2ox9Hf0FG2XcRj
o2dYmBZVfmUhvIbK49VtdecinlFv0nD+SXmP4FNMzTIw7pgbCJuGNM01GBfNIfqK
Hj/d7wwyhRMcecBqHHfzgmUVD8G7stvuxDvpm06+eFIR3L6Yl+vARDFxi71S0EZw
2+Csynl0D7hoImab4MPocfiD9aQr9yXirvij7cJ9ISTKdu0BLZJfCw86oaEfzvPj
BuHs+vFIXzUnelJGvWnuvficqM+Rs7KfwPAP3nQTe6MhRqecIT+Rh1U6FqI9MEOi
35SyVoA9DQJOJJFEy2ptOMleTWOxWo0knwcP2D5bNTmQyI3v2b7HXSdSNtPOc9fb
Vd5vRDbs6NNUqcLa+u77k1ihxFOmg4G4BvHrRQcrbTsn7EnZn7PjVUyzBI9fgnR3
vsUte2ChbHCljQNJoGA9u6JIXVJ2jQ+lC5jIoX+ZDzcrkRcEBSr8hK8h1sb6HwVu
Z+kC/K0tlRXKb220WgOc596/N1UIpEX9SgW/KVe1Q1flDy7wJIynTV+ra6fiE3zl
ldxD/i6tc2GK+XsniNukOFPJfRWfKFDun8wshyNjiwjCbEHhwLAUCwW/xENQ9+6x
9WKBzpn1Qdehe0ikp8A4kC/+/ihgpcVj27Qo+/gfeOtuI4MZzTfN7fHLYgggzINp
zhc0+ExTsLVk1kNBJHb6c4H+XRkByFv9099gOGwtENXEvjwlPYfZLUSnXNq0fKwS
kdJNbnPQCEzaqb+Wl2HrvaaD4xtynV2eLlm38tqYIX62Ay4xQ9agjPsJADss/f+M
UMJk6BiRrjG7BBagkJNPP9CZJ6qkE1noJFyQvA1CIIG2QYTsLLdvKsVs8icTsAFl
amO8PGDd5LdCRYueFIaf/kZgSeuMPdiMx/0//BPKhDzicYWHRQhyFiyu3MtEJdQS
zlXtGdpEHwHonOnXGJqejsFs4fle2q4nbvIQ7yF/dHYUTU06uC7cbWvnkjXVlYYF
nkOPHP0TthJOUY6TMS85ifTjqwvMbX2GdHYlZ/L46IyqDKvvlv9Kf1YSOSCQ+lJ1
NuhtiXaoR0VeDpChD1YfQHy230ScXZKPryR0ptxxiSwLDz/IS3NjYB9JlrkmHuJr
C2jgJwuH4jjjuOvsZUMtQIM/KjhFR9aLWXDFrEZ1tze9ee6naZd75G5TtKnGuYFH
FdReUle+84ulcfkFd8pf2hKQJ8EnRd4HvoLctHKqTiV+ipbFf27Vxcc2HTdiCH99
42uOLAuYI1SygdPJFEHFwU0wPvIFKNxTYIsRRgw0/Lph2LAyg4xPXy4pyqM+hRKe
H8iqC3bZWfxLrxG5/s+tpppF3gbu4qnCMyPu/gvogZD3Xdd0RnVOEs2iu4JC9n4V
DMNNhewGj/4xZPeaJlvUh9d/P9xTMfiIuEE2yCOQSXgQyn/fMFw0cJMAgqs+oLLs
4e7NwqVxA9ytg1zl1M+USRljyc5zibIUd9b7RQwtYKJVn1h8K7YGt/IxrotLMglR
Pm1OPTQJ+GqeiF0ctdp8/hlKhAStM8lDJlNPQhj8jLwrTSf7fV5o+6Ertm3YclIm
FnxRH3ALwVR9iTyxzRj45K98GjpA8Sd1vyVKwxrXaJdj8G1DHW6CshyQ62UUSeUF
2YJfW6Or7ZOPNSijv4zUmEo9rVu4QxeLHteTaWwPH4IwC1TsWNbxNdPiOcEII4NX
k+tZVqUf2VWtVOBbOPR8T/IMN/7wXE1bDwCzY+/AOaNwyDXktaUCpuridTn2b6PI
GiR1yLsjtRYryQBMPV7bQKbvR4ewU/BWr8nYF+0361YzDktN97Bdq7mzZHHyr4Yl
2OKbsCxFJZ8lotSeY5X3VHPJQHFCg+Tk1mKd3HzrgtyTSkacrl+2FreecwFO3bat
EhXLaMDeZuya7wqFuLw1WsuVZ7p7KjodW7Eg0hLpn7aL/3IkCo7chGdWJvyIrzxj
e2AJNPUOWEFGo4EzAen0RDOKljoCT7BAxDFEW0ucZ1SQ6QM2juSsbTCv2dPCgVmZ
KRA010DKZoaSewxIiYITkrHV/mtEfuhltMgSmO4naiOu2bx5BqgW6F83qMNuzqJ+
MZEPrZ8bOwnaKyCjDY32bTSbod7DQMSZCay2kwmJF5YrIYBE18lGs8KZpmMxxLD1
FYOrMMQo8lZBeN5jYEO2oCH/JzSWTTT+TuxeULAh0hJKKpPU4ZPXTc0ao6PYtdY5
HJ/zDYQ6Nl85/mJ72QmxUszjmxSWy5CzfN/hHvjoIgW8KqtQHAIK4gO7CLUPMjcq
PEHGYiLlFwGs9lVGfBADJYqo25VlQ0/f9bMsZwMU5SGtUzwxSVz2/Ii3QSJR4MWu
BucH/RneFuIBfOGQbdOS1v5DcLDPuiGWkNhbX18QJg9TJSVTgEKGzo4ZhnTLUm0X
iq0C7bp3CFjO8qp95fm9XmjBYSXlVdTsXEsEYwKJAE6mA1Dn3Pd/xIlbGiFEJfxo
C8jGF8r/ns2oL8c6HfSzFTzgMKX8s98oaaffkUbPZJ0SfT38nc3rXqbkW89vFcMw
0kJpKgRvVV94pLL5bChtel2Jx5GvH3DfpDPtX+8bC95y17FM58gjOavNtfK7rUU6
PH7YZYn+7pWUkPcNOKKbmIKEMn8OMhW4VjlOtCN8Td20AnArMlO8MWzEbT2+LXoi
9vKu7WU5YlmIxpBXURFNd7g/qLlWUw+4cqCwru4vr1lj1ddtP9ML34LZQ3+sxNiD
+s5p8fl80sQP7UBPv4i5BmVsfwUpXJJKoPwfqyEJFq2TnV0gxWkXKm9X87yxI4Oi
iLEMaE1QDwrwhHDgXbqA1h7S9vNed7mBJdTehSbGUOAF5DdMRfqF16m1ebHmDoM3
77ID/SyMRn76VHuL6VGE+jjlTaklo0AnYZh4o0w+5xY+wZUzEZPl82DabM2c2kZ/
BrtdZESU2n8fBxG2GC66NEXraEI8A3FeU9v2amC+gN6XL/9TW+k6B8kacv9zaSh+
om9jfsmDixuaDH5R0QJkX/BOUf1ngT3d1NJSHJ/hEUlSz7JNnxPS2VBDMp0YD/QX
rZ7ze716v8acIUdp8AGy+B7nVs1Ww0F4RRnr55mbN9hCi87lXiR9ClJd3NrdJn6D
bRG5RA2pgAFh3gfP1ELVAF7oAS5A1ryLqJbvXtF+OqaZpwiOewoOh4fxiEuXyPVI
pl8ze5KOH3MxjIouWFnwMdeVzR/Cl/hzz1feaHQzJfRCGA9tRAERsuqHKmt6oWHn
A6zbeotNISBJEViYdaFw3qmrfGIj9CckvYa+Dfmqg/yYCMe94GjrZ6klDk0uhKNa
4dfpABVsPnT29nwSglsek+BcHYKUabLzXji1Tq2Lt7n3ZrlEgIJWNZc5BVsQ62nr
eSZZlVr4MkF08ZGsdtRziSnNreh5NtfejPTgZ7qAAOEUDukjKOAWV3GAJuBSzK63
v+601UgRdXCjB6+R/XtF7s7oGCUr73JIdAzhUYAE9st7Ki1TGzdub18SXVzdMDrJ
oFOcGPmksT03c2u/QT+gxh+FzfltynRa0lzYm+qojCLkmu+lhOxiFFStxKlkrkgx
KSaj1hzmKBOOdi2p2g5wr6PRSOD7eYHNSE6mj5HyVvOAUFpI2thgL6/9+a6miWNt
98I69/raZC0Z0muxCGt1cKMzK+y31imKnC3HVZOmx+wcvhTktLJKYSq1b8IyYJp/
2GCvyLhJQVge9cNvw9nSEZFQ1M8nQA7nsrHb27WuSpuUg4vV0Q/keZimcEIBobGW
EhQVidMLb2X6Pc0YkTfxH8UsPz/53a2GqX9u9UO3TTaKG3jJk07lAAdt65ZZyfsR
PQjMtUMe2WVmt/4MrvadvUyB5Lkv1s1W1bOnzI9Be/Hk8i2MapxoR6vRLCJADEsx
H1vU2afq9sGRrfgi9jPWam1E2DVRFwgziqEKG7Ma42ZKoT3V6YSiZ4gbLE9VBUAK
MeQoFTST0Y/6FCdlO6Ku4Z/LCUF6f19irb6NT851ACGKBIALf35lObb78gZXffaR
cpX2lDOiVBhuUR25D02HVyjiISJOvmRp06mFIjXiACVpAcADlGGdSYFDQiNSakw0
6O3ploNIFb2CD5wOoH1DkenxjCBUAb2VmnROTQhJKWM6C5zUDEq8Bk60xxA2PEFX
y3Z8BqaMIAq8VLbpCeD1gf4r7x+vQqnBgXdCAYKmdqa5W3wmdqF5lSMxb9isB7Dc
wVPOaSszZH+CKF8rGje/3jk/Kv1Q0Hp5F00IUMFyE5kdq3/W/12z2bsDQPzMZGYP
5ocFAmytBAuCT7il6GJMFVy+eLlGty4P4vLnW9aALSkuLExAs/VyYixw+Rwe8Ii4
dUreGfY6DYZxzKxgPfRDTcjk93YSuZs+Up4d5F/OXGv1VMUemLb3BWxq5QUPMSjH
GJhDlLIydTjWZGBjdHiW2cGnSs15GhOhMefOvpsBhQui+wYmX7wxyx1Z3qamED8W
LXh4iRw7AcOZTK98eyT0EhlxUYzcZrO1PZVMAr5LGNjy6UaZlVJF24r5CHTI1RD/
BKgaA42PJ9Nm51wwcx317ucQMfDPIOCJKs5y7JPrFooDzNt+Bmr+TSv1aKVfoirh
0CFrClxmfEb5V5HxdUQfmr9gxqp6JW4IcfaMoc6Rc6XUpnomgSQRVAx/ReRcRen0
CzGY3GjUvvurHbjjUf1pMSFRYPIIuynN1xWKLMKwiytgfAhG91Fk8QRDQS+96i7p
/iIff85hMCtlDqNEAuzk+IuGHOYR/rbJ+YL/ntt9uGVzHgbmobJT5MQVhlP2dxZf
qmVGhCR/FcQCjKdi6bFtfogX+XfuTCHAB5wwDKyPUv5LnfOa8bzqR3k7OLRZ8j27
dpGOP0cXrqd85Dh6j+6x05ydD5G7xI9KfQfUghNuJQmu2vr9DWDuBTAKcic3yhgU
bNXbetRCn95WlKFrKt5lnNR20BdSUuEi48w2GFxlllD+o91EByj6Emx9uELklO2t
a5k0qdtOEYJk7jhSsALNxaDggTCgjB/kcPyykDZDJ+ovsAHJN6gYtETYUde3ISni
nGlv3ep8mufketw7o8R0qRwuAacoxhYK8wym95VaXiGzm9qXKIpYL0Us63kNJ7dk
gVB88Qhbf2aGWPqKhGl/GlBsxMmqIj4nY2plHxb98iaaJShFB6W8ZXPyY6+wCg61
uL/qNiwWyw8OIFPiTTkXEn8/KYBew5yRTn1W7LAtBouA1DQIBkTv7Y0MW6co8rf3
01K5ENBWLoPHUqQvdlWvOJyXM0Q3aIIDlJ9YAQ+PL4xgm1LLvfMHVkHm2/uHobCO
3rZe4D9fc9nijOiOXj8dxfUSjOEWyXAiDP13b67F2yiLTxdNGcQlTW/9iOc/5RuB
VJFIr7TI1qV8O4S1q5BbIyGw43UM3NAtszG5QX2M75Eml+TtZdk6UtgfI64xYPEu
ytoIQ16lAcxxrudWZxHqX2ZKHt7a91929+fqCPyX+vj7eF8SD3m09eHMg6i+EYe/
hn/wThHw5ziVMQsDMLyUmtZJL9F8kvHHiMheVE0II66omwuxq2uMujdwt3mZ1Tnd
FtPHLovwuPi8Tvbt91GMTN1cGiu633K7krakRSnGR1skLi2JmEWhPNRGlaWIGiz9
RoOH7ElAA4q5rB1fvsLsMhdcTPP/HoBqybxnwSBwYhRdPLN4uL4yznqu9+gJIAdG
EC4FYL6xaETU/cZglvm1QhNhdmokEM4etKcDd4wSKVj/GstMU03lWi01XvRccfSj
QD1cs8qhe0xvezMOQBEeqEralB9dvka9DsFeIYK8CeU12eGRhf/JxML/WjOAwLaA
Ilu2A7HuLspMbBp49AFxqIxrWJIiL0ovfVhlFGqBcziBRSaL8LHS27mHCBvtt/GE
J8FoROaKQi+BJI/ADS2aVyvJ34CwyfDQNgtrWOnuHwSfnBYh/tMSO6k4BaPu2Aqg
z67Mtdl+Hd6wzDf3pdBDsHWAByn2WsnSGBlNgUiVkjZfUDqN6ur647u4b4HHn2tv
ffkiTPiQv1xBLN+tX1Xd83WEioko56jh5TyczzP+1kloggtD/xMD1jMPYMXAOVTW
IDZZrdnMG60peUpY6+nOXjbQBO1KtWlVUAzkstlffW8xVpnp9DI9PjHRgiZtqMgh
O13+Kbs7UnTLb4yjsq+v8ngiLYN3M4I2ASjnO85a55AuiHPaDmRCkgaqm1hI//jZ
votqYWfc1MDVhP9+GFKzZ4sOOCU61Ga1iDuvpBrpesxYIJ2mhZXIhUyBcU6hWTHi
4WFxkXevMDGIJvRwhKi8iqp7wcoZc8UVV+KaHlgYckDhvftZerNG/0Na2JXGpyNt
8nOh61eKZw4qzEWGgcO4Zu3h3lnEhLq/vjpupAakAH3b84CoRp6rdkgCufWTMRuZ
SxXn5TYRXR6PwM91Lkkgr3eoWj9j+o2vOeAG7uvQFqaNBJibvD5qNDQD9FuLkjtM
3xuzMO6ctR0pQMzm/sXNkiJgu+gUvHrxqUQx3llZpJZHV4Ssf6cVRmTS467kimWQ
SEQN9xiUD7P6gYGTZLyT/GT4ULHQidLcM1zQY6QmRNUn35ppx1jPTv/M2fU+k2yN
jsgrQmQdM/kASzoZpwn8zcKAXXAbZupr6ijSSaZmbkTJXCAT2xmHncOXUocT71fj
mn+spK6IsJ7dn9JtaR8k8y+jSZIa+07bybCPymAR6u1PVOtgc6TlLQWuVe5oC3YB
e8a3M+SgCuc39TC2NA7ubNtQGBDPzyEIKXCZ7oYy2E/b+9oOhQ7FLrj8FqGzdwLP
mXWQF08eq2ak+RHFYOK5UHvkGRF938a3CX2ioc9IOdoG9ldFM++jSavA1JpjT69T
stcf7zfI9qVuHwNRvwxIkCPyPs13Ix6Xtwjuhek0RDcawOtZe9vC8+X24XgLr0f3
TD9QWjct3JeV0E7BP7JVP+yuR1xnG/4+3drEcVx0YIirVPcwG6LGCzUTEdhctD83
IasJmnPb6Gm3do7Syi1uoJGf8OgO11pyo/tkKei6if80HCXT5pTXvS8l6Uhxdirj
Jg9MdipMXOg/jKvcoHQ+E1HLYzTs4Bt5oDyjebTdiEYKnDXxBym7Yr4sES3Bxc8+
20dPjPv6tM5SF3m2PvNSQ27aszn3gRKMEiB0WUslQlxCWFbN1zjdqahsaAZ+N/Ja
czkFAx2+Fr0kiFk6YtuhmIRDJJIRi113nQPcnrOTJI2Q2cFg9PyxLKNS/uc9VNrP
W9jVY1IhMojUUoCxuAjHTNrP8FDU3UdsUKpGjEfDCaEb91vphDN1aDIL6UmOKNgu
WBZPH7I5Nd0m700NztvykP6Q1F91pgzaf9SPdvsEyx2rJpFRmqf44btZYqaLhPsm
LSgVmtfBQ4LM1vzLAVzxUw65H/sfG59QtMQn/19eGd0GHEFlvPdcXmsDHbZEsZ3Y
s3NUgq/9n/TSxnl6h3meHJjC1GNC5pcF7T7zEEcWFXkY+woaxJmV31bZeQFL9SVU
pvLo1yNOe/YY8SXYD5fo5VLhwiQ2WlNSyfBWTGRj2ytgeLcYXC2RjaazCKDboqvt
8V8xU+lPNizFiOuU6cJ7buHsDKWpsGytGCrldBzE2QV5KOe+SdBBeptHvwUqsdQe
6LnvhUBgYxPIUJ9xvPcFzfl4MDW1XmGpJHxYK2TjTt9hMqIOBnu8G4GzvfFGo2Z1
GOic04PHmf3t/UGQYHpxIC9bXbSZ4qGC7mhEamZlf/NRipcR4wUeFfa7ZvA5ftpo
9aZgnXYUFAirS9hwEXyKWZmR0kXR9bK5WZiSMTYopljwUlJNgSWPwm50i9Ty8OoU
ieOx/sNZbeDaN7VLB20ukU7UyarGHgwfhO4QIJkbWoZlRjud0WwYH4DLG32j6LrD
bZZHUAHURgU4M3kP3VM2B97HpdgYaeg5aot6GyQ5OYHd2X5cJrGEomcUm9wvMpUZ
DgkWXOr6F7mS1NRauPo00yHUy2ccOxntxXbHzYjNPt+ATDZOmiNeZw2cPAag6JTi
pUX1vYMzWcY4NBEZq53jqVhOByd9YnadDzV7USIMaM5pnw6qynKh4/3T9EibPVYr
rpzuNuXJJxt/kjOl2LjFA6YRANuU4/nGtiKQG7i9oFgAYpkpNxNjUc7TWAKK3Zef
rOKOxUxMvF6Z9t8AjjqrWAUytQheE0OgNFKYEbTccUEBGUqoGDCkPWM9CRm2f3RQ
KJ8qU1wInzdG5rJT72sFuHeB0VL1M7Ex0E9Cl17x3ifqGz1xqOXblbIG3o4ENXZQ
hWWn5Kdea8ApS0kfZWJH5KMwSXbwOUo9ohytr8een/O6vyz/v5Nfh0rsVj+4h5Qd
CcfhRYrum8cgd1xf+deguDEvsbO/65Xmmv77XAs/zoofjNwvBMKpkaiwE6B45EmL
ocSAiPPfBYQTuIi8zPxJipfUN5b1+bYV6/lTo0WFmDIsnGP/6caY7+Mwoulnxxxw
0OY3Buihi51u1JplH/6VlDYZYPAiFSJoQEW9iUPlfLHnVpBGJ5CWjw48FMy41n51
Scd5+3409cHYlcW+Pr8wC5LBVja8xf4UA47gOE/8opWRVJ0HPT+LTPQ7W9aUAZkK
3n7JM6F7KhcYzVAwU6iGGOiZuKXNBpWBufbgLZsJucUtG3ospUDuCGXjPyVuiL7/
rVGN5yQceE8uDH+eb8nVEA5a+Io3BIo4YwFYXPvhy3wm5kS+IcDV+bb4C+i4kwhs
wJnGMEMKkgsJpl4+ra/qdLlaHkknWecCVVkCbw8n0mr6e/Vobw9MBBh8+tHBr0z2
Bm4aFzR9lojxQ21MOmsduZEbAqLXw8hFFoiiSTgKTqM3tc7+sA728E/G+jYzmPOt
69xFvIOIQQblpFNzWzU1TYzrtKiyuo85pMbb87lBDWikMicj04tf5rXHDbmEckFH
zRd85yWzn9bqKS2E0i/vhUIcTj2tUi+bzfdBEbdw+tGSHfGY1GSUMKBtjI28MH5T
5dvBsFXwoikrIIxbZLTpy105CT6oGJ5BJp0W5r+6J9Seu0SjVtTl8I214MHMfvRS
f4Zo5CuDq81Lp9WgsyJKh4Kuco4kFLAFnPGnS7KdVIxVax9ttlMe4Z6P5T4vDkUc
BwUb5OiMYhXyrrcQ2qjpf2KGHy1saAoUN8PvsopxUsmuGdf/wqBvCddVH0NldM/8
danYhkDf8tTtynNb2/OyDfOmqgvpLYBnwqigiCasNeqOUkqHNXhI849f9sB5UqjC
rb8rMsOfzj/WGZo+XG7qG4+Rhcltd6ZgNDOcBEv4/8SZocVhnZFbu7nk1CChfHqx
Fch/ZV26dd5C2QFt+tosS3/uliMRF/vLH9y+8GmyeupsV7uBSj8mX2hdp4rG2acz
u5pu34cD118f0m+5lPocMl3c8Im5vH0/k8c6LCfaty70yMM7zgasHD8QWqg7IIIV
oazsIeK5ww511gOzdyTvAMrjma52JvJLga06Dtb1LSmsuZCpSfIx5GgBnXWO7nZ+
ldnm+2v13eOLre9NK/EpEH14hQBog/fJQqpkNl8OWDw5QBwOQQQlABet1LxSTeTA
4J8Gc+cxpD9+Sy5sR6hgtLQO17F1dtIpp63q8GqJIF/sfdx7gJMaRnXRbZE8CYAU
0M9PRbTpZ0m7JdTwxAOYVyYmsHHQKqvXEKKAx3ZhbzCZdZdW/blq15CYxsdeKrPG
8hnYOsLVIRF1N87h0FcMM3RNq9FjksjBKCX+CKz0fYLzVkUHlLte90sRTWsQlUE1
9OiX0U0wuuv7HA89gGXDxEUmGxSmikOWdQ1PEDhr3IjEYP3J2MDfE5J3zw6uOAUJ
wxYMNnKmwACg4bm3NCwglEVzHMLm5MqYfVV5a/XhKlAaTWSijFKant5Y3dL2QaYL
yUydCvxgtvTbDtJX91XCvqU3V7tPOzgkO2sOyHoq7onO/OyqzJ1fawe1hZOH4kPO
TPSlHa88N34eoxjtS3LJ1NT7jODNTFgs6RN1wGt+2FYACnTD3lY38BzypfyhGzTI
q/T1qbPSKT5vS4ObJMzyHxssE8p5M1kdI9wD1iT2RDaedTuCJdKAKGCGS+4N8FNm
17OOLr0Ie+Lm2qcTeY0lQCT1fqBh1JhwM2iWzqw6TCbifjDy/LXFvzyfWyvs1dEp
iwDN2bpE1hsa/MRzcSzEIQ9/NfAYjEF38Wmp+NVbbZKJjAuxC64BcCGHgQoxEkG4
H9fCt1KQ4Rhbe5IM2V+C6BIfUQNHWNlpjvT50vqfSGTLfJIrQeFPQrp1BLdVfvcV
tUoh/UWF+k/haKnLdnSIWgEp96PlxYc7/Qsq/1vftl+rdt3Weg/9FurB9dDYe5ab
OTax8xbTMlo2Fh0X0oVM23H1lGR2U/8+fD1KsQani1CNcpzd7eDrDPo+c1tM6vo3
VPsJSyMou+X99eDoOsX0be+88v0YMmUDGtWIDphwtyzb5Pn/xA4HZbTyo1LfHmyv
ADMJ312HQGSWNQOF/5ftfVd/FzkpvameC6XL4xlocQywoqmrXMOcEfxAP47ETUBj
ofLsREF7vZsYTQk4JIzRxftKnCJe6XGWNk7hiJ9dQesIkocNIlFBVrI64cE6/Qf1
63C0U1JGdO3jyHPKHKhJMyYwTqnwpaGaUXSi0NfLGPpECEhSgXyjG4pBvHqjCNBO
atRM12MdtLxm8rzFugHb2ekuXENED9pMzwHcDZ9HqXxwRhdzug5gsbO+zJf3G6zg
N9hRlk85yhKt10XVxUJ1Fq7P6ErBcObAJZz3KubX8Ntb+qys+ONXPZqlMTi9ftgJ
TKl9h6GRrFoL+gMYN5hoDcYDKYKIPKCYzFfRA5LUbUlgBshoTGer3jyIWr4losQP
1RX0DqfMVe8WprjpSu0p27CXmsSd93Iu1tlaQH+s5Oki9SSiEvw/3PHcZpNvHmE7
ahbRyD8u4EJuq8KFnSGtKKxTawu1qqcPtamq/JYXZCgvUzSf/JocjygNtcyaFq8W
lP3sHCo5wP/Y7/+TXJlnP0RN4oC5nuHw6WLl77wKXwYPWWdsnGG1CEYecKWZ/lHi
oDJHvKWwtWJ1UaI7doBE+9njhjOigTu9CBG/IXaVVHSz7fqUsLgblXa5cMHLClNy
6OnoRkf6Qu/0lM0g+7bdN05nYwG6ByT1JJGVUIbv6UmusEOf0Q2ayFW8xRwGKUfY
ZtRpCsSyfAms12IIPbjFCjqHmDJ7IakdxwwjJddt6wl2GKn8fDS39lMIgnPTeHce
T3bg8WEUhrJBd72/tnC31+BbkeoiGY0v+Q5SBg983Fh0yT/NG4umrTA6gxBNICSw
GtgHwuUCTwUK78wcO/eoAqcDIX6mS2ROTAv+PWfwoWiF+834V+cr1GfnjY/F4sYY
2pgjM41nVaMpl2UcgZOj5YNKPDRmRM+TuXilHp7tPSq+jpUY0slOGHiD56bsV9pG
y0U9XeAReyBpaM6ZP8FLLASVnYQkPqRe8JLtpI/AZxVQ91yx/eZ+jx8b8T8fmldK
a7GhDG/d149pw+oIM0kILev0cD4qdgQsIZkxYyO5L4+tPsPR7uYi1oFCLshfGnIo
Dcox2ouXeYl6P+BSuMVDAJIFXDMi3pzpzFS831Qwu04Pgc3hxtk2LnmuBoH+0Cqk
aPrPnWF5G0ipCGLUhuTEM5D0SlBmo0MPErnr561RL1actid3LMvlxHTddiHk4aNZ
6KKeI4XgYwjoElVvrJLy2Opp1FWueZlLjIAN9tYuxHp/+ZlHBACm/1xDwzH3AzqN
IANlC/iZArvJ1U6tqIbGaTq8cv+eR1QORwgfy55vkjdkz/6uLXFfhalQZdja2MN/
d73ICOcBTPu36IrS34sckAjxPoDKaTVk4yqweCOxpluDKrBFr96ivfbfG83nvtaD
WkrahkUfwTlFaMREHVGHdT0AUKYltmQgYGO4UfFSa41aATkgH0PPyvZKEgUIHnMp
OrS2qgDUjcTblVoWeSSZsfwBjlFZRPImHea9U3NbP7HflB2HUORTemh9ndmn6XNA
pbE7qx8SsjHaoqe4NdATJFmRp7/EB1ishXTVNfpUFayLdBrBUC+b9LPjGINKrzo8
jzu+jAU5mYE5rMLPQKFhL5n0xr/gD2oI9x77DG/xARnsGF7Q3xuQY0C8IdZs4cMv
n+4XDymP8JkzFqM8NHCeZVSqfBC/1ExtnPknn5lcAAwIPY/IvKAReD8GPdIKKLkN
o+xUkE87F+ovQq8DknaLry+mo2mA5uGbzFqim7mlHb7T8D/eCc/pEX5FmNeyPrDO
/Z+TyhPxQkshk7iznHBDb+AR8PaXnv1ERAyh2J/K85u/mf2/VOrIZysy3oSUkcqR
RPAruVB9pfIClYsTjL09N1GXH4DfziAlXPI2cTZOvK2lAUf2GIZp685XLDKrhxIF
RQ5txIeElam/7yR3RHEs8wbbvqdqT4yi3UgP327pqDK6z//chFlcHPkcakYyfua4
BWGOy24iGgnenH96z+CY65gfYHAAEJSFLGhQWmMB0TSBpZCvWO8pLVE852yk+yjM
zZIM3eDQqyLA5n0+VCQCgRd7xSpH/+982UsPG/jVP7ZB9Ik3KM2ZbFL78rviCOxB
QW45I3/i+tfXCCPm+QqRA+pTJmJQdIvekgEg5hCyX8NCwWdFGOZrEC+x2tEhiTul
wutlSWEB8j/bRQRlQUs+9jkji8tF8YqEHBJ4p8VTZ3DQ5K5XAcvt7FIPpZUpmgPp
9jGE7pfPBiTDgDpKY6D2y/7vzmZ99oC+rsARw8XLCI9HpOPx24MCSS0zVWVqO13+
durnn9L+n67K7diPEV5H9eqosaXMYCD/RzAa1nQ6jkxeFPkCekUWX/9PTR8MJWNP
fUO9TUxe5vh9akVr9T6AFF8tOLRRV5MfAPk1JHufkt8Kv/AWnxKjsKs4+dabQBA7
VtWwBLT1yCZyIDbXcoV72bfd+hpFh24UKy24AcZoQggOI+Uv7laryx284BwxdoDs
+s3nz80TMV8RjjadrOwRePDHHcqrAMb4XM9K6IIRNe3uBYpt0g3pwztQCTnPNueX
rQ4eYpX2FeGzygGrl/VvtvfHaIRNvy45Mhew+6ixoUyxdP0IciXxkYI05iFsGmoY
s2Wz3ITfEMJ9x37KYOy/WPgj2pah/9tk6uF1sovmMdnkLZqoFWN8QwfED5FJeb2q
2/BlC3JHT7FMVnbZqIArQOTRJEATLvreYnrAY/YOdPuB+hSq4kBfwQeRCoWX/ZP1
+pTbIS8lD+5DmVSYq29NldY72Vw3f/lRC12YZVfyMD9Mh5PYZIP/+Ot+4gdn+bew
vdPG1jeqLNSvYl+yTzvuMYhjKiW4z4muhq6peS71TTXPLYGtFSl/TA0Q68SQFCBM
YuiUM/6qOOhrKLkdHQPfEmwai2bnFEj+Qo4DsVE4ajkyAVbwIGM9M7rYuIn/Xn4W
YfZp8MgjPOR/NsukwejpA4LtyoP4uQb4Ecd+VSs93Fk0dmIKT9hmq/tDli20TOad
pgshodxtejq9up9GPhR5Z+lAJO+0UFSr5c1ra2kbJNkV/qOsMctJHIg4iVhO0dBK
DxWFJKp2rW0m2bPdhFv6kAYs+vvkNU5/wv48KQyJmR1sMBpkmd8kPMxThgR61km/
Ax2UrelhYtFThabZ4eRZyPv0B/d9BTC4dZkR8z6vfIYVSCiwcPdnhHcz3H5B1PuY
pVAF57tP2hV1ylZkL3pGHyCbyRxznXKP57COhqROuN+8z8V35pBXf6shVg+R6I4q
HyqdT9wkbFmH3Kxv9Gz5Df9nnLK9oX8CXw3wTkaboGRk2ShjTeEoXO9Ha5gBtnxo
Up2xm5WLbBruPXK0VT6My8msX8gM7YtN1XqNEUONstT5t+//+GWoltqd+lagiWvC
YWcsPy+g7t1de5SC3eI/OqxQHnJL8NZ4rNKAcCk86I8t5jQHFt4KLwa2RtjI5G1a
Sbbm7K7T4vkMjFIcYhJJh0ei+BncT6R27KQaYerw4IzeF6o/wlYS0N0Wl1zHlbVK
8D79Jq6mKPemeL7KEzVA5K6fV/9wB0mu7KXy5X4xppyqcvN+Ro7OV5azF3EN8lxs
ZA3q8IjBFzlyqHUd1/rDvMCDidhgUCj7I3FQ9nfPmRewYp2tfFWkIRmz2SQjwqWR
Mu1+3vbPI9xKu2LOYtGsbxmw2aAlz3wkZBZKcccCsePA/xNdSO+y1gum+bly+8sQ
640T0bFA9HYzYPCynlAa3emxhXpcx88G1PiBiDqxn5snVpC8D+SyzNr2BPtOmKbw
1zBe9J1/2h0NcdfIxLtBmQJp/2bVcdOWW/CVIh0V5D1xaeYyv7aZa2uHs0Sb31Fz
vxvSZ+sqRFwfl8MRV6/kf8sAsh1G3juYj7RZkMSG/02CaJdhfJwVuZOs8RM/d97d
vvBlr0oBqa1IkQv81wspKmRbDVXqo5MBgGUHJ0Pebc1KWFVzDQurnvy6tgud/qnC
eopDxbp3pqSq1rXAiCzDi+XTvof+uRyrZk9tGUfWMrqgRN3lSsGlyyCIC3yyqz0U
tnpp4aUphvgU9yIZDnb95TAyk29J+mBr13evci/z03WzyJWRbRfJmZ7161uT+x7F
EsutrLZfAx1ByCPV7MkNVRSZHEKlPg+wPj88WBPgBZ/0JQckzIOVanD8eyx0YwnZ
RI+IQLe6nhdy5yPCUaEHiD84suogVAw8bbJLMn1fiuNT2W2J/n1RtoGc9r6FZj7n
oMsK6aqBXgu3RASjpS3jSFhKkZdTc8qHgi+2m6N3MaKD/lSYPCQ49WKvCxO9eZE8
lpvbE7SVqIE39vc30n+5YzCnAsUtmnmGopk9ohREBTBX1Aag57vtky8hWN/Xlf6u
fnH8FRJ4w0wLDNcZTT9urRvDKB5MzEfvEr8C3xw/Oy6FlKBlb7k8uN0UBlar9Fsl
A/08l65RnquqofsqJHBq6RbbfWxsaWWAOt2sWq6n2BpB4iu3HsENZibUBlnNa3oS
tmtUSmMEI5N+Yi5+ZMpcAZTobCNzUsylL4BPP//pQy+GTs5XwQ6jmItRenGM2pHa
YlqjYZzxCw9GCE1TizeQ/0b3LneqZfH/pVYRRfTWzjqiJwb41sqmBXey+uw2w6SI
tg7s9bwPBbdZV5Iz1qOQLP1XFsf+EWfxDcjR7tsn6bjd7XAEwhIiZsuzUgagRFHn
3y0I5c+0rO0Wiw8hK7d+KsMCWDZ4untp0U1LjaKOSNtE8nYlVBLu14DRi20gO6dn
MBD5fxudWTsw4RMK21jnrCrnhC1vgbp+hTF/KTjN2L6sKCjHLBa4YbxX/gKgH6Ne
HMctPnh53/e9ew33aSY5qdZSGL0FwDzkLRByBaJpRSXyos/kw7WGZMC1VmJTP8JL
af9jHLUFjrYm8oLmg6PuWqqYa1xzVog0kB8BVH9bZt5tcw0mre1Gxse4thvvEKb0
12Pyy3e4CelwWL48yn6MSvueOA3AVGMaB+mQWFzye3tpuQLTvR7DZ5oNIvIEfBdU
ScY1RPOjOHEuD9BmyzcHWd6KoKAReRJnkk8T5BsZuuY8UFFZPzyfPaEUmf2AuiSN
nyruFakeS9rhHj+lIEPD8VOHqYNrlP//owU/y9YRISDoU1xBLnmn/2kcVkMz7Xc5
ujAg+O7bmU2ArK04y1Mbr4yzy8Xw420k/z2JNFQzbBoeTlsLqbwDG4T1NiK4vlp8
Pmv6FcGLa7RAkC6hABkaeBc4X61yZVhsdQOLspSriPu55LpIWAGwvQpnA0EdrIeT
1YOPDPCK6uDamh1kb0jfIljbi9PTdp0qGe2PlUQ6NPGtO7XT8xViLHMGUzxuKnuc
Dqjy6zafK2x2umYQ8CiPzf7YHR35sDlzuk1A7sx2gF61k/2UM37+BuMRuS6E36B1
wAWwfa36UGc739TEuT1g7VelutOXiYXugwKB+z3clRDSIP5KX0fF+9qUaLqaJxDt
0WY3IsQG7c8CRt4GRj1qYA/ocByekvEARo2ISRl/KAGBzauWzYqnR4QiZM2f+rNt
3IdgGOzz4T1Vttz6VDu3CAsECpxDznONflthQNux63OHgnnYXrQkFajUObeTC3O3
dmcNGmTIBIlX0/O6tdow4udeS8YQoABRGs/zY7rkquQK1depgfwlV8fKHvgV/OJh
SMyqa0tu1L8h8wQ/rrpS7Ungsfzg96Fz+b5eRFZe17E8c08ptlR3X8neziAiazoY
VzVpq2xEl2wqx1o8iLx7nenOhJ778zvqIuDs7Nx0fZZd8HQagjxFiTMf/72AEYUj
NBXP2oRfMzOnTddwEWJ33uoL/dRxcUx3inIrAtD5ZcIUmANA94mMlPfJPmYdtOai
G1yjqcEKk06bVj4zSCYg2w6CDClc/rKFk9beCcRAAkZdngyEZYlsPPxZ9TJf4c0Y
cTaGwuRlZ34JYr25j+RaJcaCaa5GdoYYYrIxZQ7l8ULqDA+5Oaa8/HSKQ3QaNuDt
fSalTXKS5D6PxhwbxH0z4R2kCp819tbDHl3LHunbnGkVby+M5JIGiP59n60SQ5w2
t8cTWsr6PMVlZfJdnPrQWI5Xkd4R0ZWEiiTChWTQKXg2esIudK/M2A/+bgJwMWvI
idUJXCmR3XLa3rCPLN+ffePT2s9FG+GweJolNx7O7uR1jlcMbYVk6gNxFsE7K04e
XgI7nvCxEpLRJdECnjor2QQuVw/8rDnSt813GHazf9K2zTiKPkyqUDmQE3TjPuRn
/5DDhksxYaJN4+9/o89moCwmt4h5qrNc8kRkbyrgykj7UawqICiBiy89c4mW3piJ
K4V5hDKt6ErkaF78ATnExjwyK1HI3zwQAcO4i86xBTvgBiHg16r6f/6L+iYjFWg3
R3b4e9qGN563ON63Cbe8J556HcuAr9TT3ZijYfQOLSHUdXkLJT/PaAFYyAj3sFTl
WDmRGSE8XZDi6ztK2AAzt0jqbHqOPWrkHY1Z1KWLvEEePF25dg8cymtlhR9BqNTV
barKCh7/Z1elbFn1Ji1hLS7raurxJbTrv/301XUa6TFhb1UFhqUMBC7WVVIQ5TFv
y8Q14leJ+TZFPhGzWkQIK0pI96FWbtrggC7m3dSN1muxX3Q5BXBl42XjLCWKzBn3
d4yKNymQ/PxdQSOeZTF1bnWwZVAruBdMfbNdCVJrwgmUSOYOVV5vXZSyMRLLtBIV
3EJGe2+Skn4gdFwrfv1W2vEaaBu/P5Ux3CflXHg5Wdaf/v8vHO5Udkr8VjvfGoNk
8Gz3weu2m9OcdT2IE0cHduVCaoqQ0uJflIpiHUn0LuDsRhZfHbv892dX99FRha6m
eUBvzxjBUIhVZ6PsoPZ2rCShsh7gqlmACD/tm6eeBJeCE/gJPTUMs3ILCSH6bDA7
Vr+838gJEjVw1IhMwGc0KnpVlm66dpnHdOQt4FsTjpZ3AgsKU/5qPU/wpcNOkrYD
+Fp2ugUustn3ZRI+VdMYSGp/G48IzBm57k+o7553ZUBTYU2ruwCN/NAZjifO9bQ4
qa48B2Vqja+Ka/S9M0Nc7FdnUYXxI7bBvA+2eU49wRlCgl5zJk49yU/NLTorkXNL
l7WX7JtKniO3lQTO28yI0kum5nHGc6bDwksFd78/cFazcgkud01zH5s+BJPvY+UM
CCWMtWqR0OAeaeJWbYUbfaB40bPnRkuHyxEsyIz1GA2o8bQdPIOTcPLRas9rxzCz
YiFX9yBRpjo+Wt5hHus4N0yjUX12++Opc9lS1L+uc8EQ3JY+m1TxmzeYz67uqkf0
LA13BApgFRcxJDkJ5dfVA+KFCkBCA63wJpkJk/yWowC+f4jb0X8E21HL0c/D3ZrG
pRgDEb8PUQvIdwb38b+lPE8JlstWyrj+iPAGm2GriHQr/gIr5DQ/3zQC2gOkp9rS
A9GJfAyXmurJwYmS5M21ak/hSYoeinRqsDChwAZ8sHR1uX3pSvrj0T1WK+s/E2yo
hDW8xUjNqcOy+fz8k4ZFazf+pV3t6Xa0g8QFMviF6HVinMviw2Ra5tkP1VjgwLTT
ocIyQtu0IyLEB4LGLF6Ny3a+9kC9wP9fov9ApMSGtcBTZEUsNoxp9Xjbh3bseeXs
fDkL0km8U0C5m4d9NWsUM80WRw/j1l/YJiNRqXW3KFqH0OXNDoGyV5VzejC+vbWV
XfDJYWsxYfU9DAcn6hMmQ/A/UcB8IFhiIb5ts+vsuT+r3qHOoVzqexUYGowPK/lr
YwmRtVyrMQMEFINxWMyK+ZGoXKNdVKhy1PJCBfHGdDcWyHjLE+ffM8hFtxo+GEuS
pWKhaGoT/5ms6+njPoFJUv6dsgBbi7Bc5Z6c806V7EQPtGS1HynIA5jjdc/i1Dn1
ed0zKB8zbv1z8i0eXHQuztI602FL7yPORa7YANVF9Je1QfJKPEoS9w4PDMUAuF4Q
FSY9UOUW0JGxH9wdGqJ0MxXJv9ywFC5axaPLMWmj0OPxVeV0a/APJ6A5tvbrxtDd
YSBZmpOSg7eWi4ZSNPHV92Rvdo39gw83TlxTAMmx1nGfLfeE6R0pFzhxluY7WoJB
HMGTevIaa4ktHkrihYMu+7e1e+3EFYkvm7+NJiAzHtQtBHdFJkL4lxI2TPxmzDfT
WL2yCV5naTyQLktCVRbRM3CNtzVMXu6hzHAdHaj9fz3/uz+ftYlBacF3yILzq0QR
zcoFJ6Ld25St09+lcVbhG5ohgKBYhYVNyCGWKlD+dVbzLpxPYdlbuZxgwDRxwbnb
UhWYLQZ5QQ5oDIxrmTorio1kxQQ5czSz67sT3ouZVtXJE62h39XszwPTt5OjJ+WS
Vny/boTtPM0F7R5mNC754c5FgpjKlMuCLSrCIj7YoSN83eDFzdNJM6VSNwLFG5Xz
CfMHfB70MzlMLMxwzft1PhhVVUTgF0J9R1Wl0LS+skB27LBkuKq2rhFUAA9zE3pR
OZ9sqlCkcGZvDkF/+dk4GHAU6fccuDYnCHBptH+iQ7rAr9463nI5hRS/IdTm1R/h
r0lUtIF5o5Hda6HG5ptPvrREnzGxTEsCy+JRrUeRurGiW5D8YT1YpzV0mxkIXsX5
ypzu4j8cjUldG8SPMyGF4qE+01RlY9Jh8ns9wjR1z91CDQSdyVjs+xPYDDZ/+xYg
4g0NGpGvSu4uHtaGBxbl0MuE2O/19beLM5+CE5Pon2eCUuNcirTNsB9mVh4zsUW/
DiMYOTilMByW2UM1RMsNzFjdHIDhsHE+iU1YAP5KIXH7oTVWciYWcd5EEDET8jA5
fVJfe+Ywr85LYSuptpLaJJEAzyNbUc8qfuYyivu2mml/LtgSGjcw+eRWJA1K/VkJ
Hw/eXqHcE8jnBHZoPTKNOUvKV+1cAZl4TLtXJ7P5rArHz7OtX4oFViZXmhW/kdSO
53+fODwKxT77l8AcRpiGmx8btXCuj/ogqoFCwVbtlIjYpYIPfJxEtFlI4Lb2ID/G
dMlSitDQa5F5se7kqBTr3X3JW48sN1cIiBN2UMC1U1SJhhxa2Vdg8KIMxedrSN/b
GfbkfJH87zVHMno0weuA1Pmkef9V42brspJpL0JyP1NYRlxw5MESbLn0+jnvykBa
1MVOPRPfa1UF8fJeyzko+HFta1DoBbOo01FGJsmetCrIDEg3XMqhYw6BUrmtAt91
s3oGjGpzmpbZTbIlDd/hnLQZ9pSq/1kkPE8pJVTVOEx/VHLC15h+KnXmw55d82sy
ZMJL0/oWDrktcwD4Vy8gNdS0/Xk/Gu+H49S8zVu0z0wvAZOJ1QO80tEM5R3+y1sc
1u52xp7kjjuW8+mpv/TCB7Na8LbkZWccsQCmYwgnedgbTvtQlWx/pQGF9v5FyjRM
hwftFS6pXbfSg9uE9Lcpitw0ExYCYE4QNCXwDQDGqeFS/e8MJVqUNQB4jSbadvFL
M289PRU4zU6NvIXR5/44rXEo2nbCVjBIYwV7knK+mEh2BliEEMZY/nURLaYF7s3r
OYlsWDM9Ag7n9BMukPeQXAaV0cKPSc4fUPgYcmvWQIsK/PdgTDZHo8jTZVFQJWRw
ELg75YeTkl1Lzcznrjcjbqp7/BOS4MvYCvIVTJO7vUwieSf98xwj9bIwepbMt+H7
WzY38Om0N5QfWnkrIu/hrFdhhGI5ox4Chnujkan1h2p7488g3uTdxIEDPKeM/5ZV
JCfDi6lW99Hvef6HJ9QHSJw8oMEu/6IMRoq77TIf2Eq4CBwsbwqm/qCdP161Ihzu
lKlodGNeju9IpNpW8zi770YbcfhUM2OOWK/SRw8vvFZJ96PHm9aQqvtQ34qLifOX
go/mqVZgoZ8w/L0ZhEOxqAEpRGSXl1DQk3dnjQhFqfuI5a2mwsfXicn/19kZBKtw
DAAd/9T8ISJPKV0gobvd+XkN7tnZgcddGq2doHm9+LLv5H6AhPlGOOZn34InPq1F
OZRzJw70cGLZ0ZxH3qJ+s+6GQfpoMxBnd/xcXWGYDq7YXy7rH++SyWItCIqnOJDf
O7euqw977I8o2w32EvgyxezS64Xnp8A4K58bWahUol+fSmkeK8B5CKuAHtaGNDCX
9tVb8LJBJ6jtoOygIA2FJ2i+54M63ubehbdcVU5txvKyYFdYAFB9XwIBqvyvDmm3
oQbziLXUvlvwiC/QEiFOOidhKXrzx6Dk24v1iU6lRJWbNj0anRlMzd/mnpL6mJvO
R3jj3TXLblNSqDN7/ZkcKrWWeGHfJNUb+SQUNfLDZ8O6lHdrDSTcBdOthHl1D7JO
nLyEzXH0fh9GpwlvIa2n4m/+s7EZUMXJzEDuUAPfIab+7Xnz6XNS3TxBepxoU1f+
sL64pJwoI4iEAKYclp7VNI5CbMxg+J9SsVNmfSIfKF3CcZa6KiFGZBpEcesWSs4r
rhWuDjkf2lS7LiiS7517V8+u3IEAqJscIfL4+tcWN/RY8MzQ84CzKvFnFryU5Rza
GoCzOzU++Gh6Nmnl/87zDtxoAUHFXxNjfvQFw/xdanKSwQ324VqF4OieMfLehxEY
adH/f3MNI20D7koagBoUjx4AUivwbYTin7QMug1CN4vXkO0PVw63JeatTVPEylfJ
6fuLEruKqIzUSkNHSS+ksLMJP4SrF7mRWoR0qp/yFV9B2MDMoVWHaNW20dCRpCIQ
uuJWShXX1yGtBakCuxeEaDZlUAdDilrLBF2fROsR1pa8hL9A1G89/NFYoQlAJ2ox
ZYgOl1IgF+9wdieZr37zo6papzorl938WQY+TBHlK5nKW48mZr/Djkjv2+YqgkDd
hbnVsKzpo5F1jSmkWnw0dKjshyf2gRGHbUdKql+5jQGSflZKjHaPC3FawG02jM3X
xYswkliKeBg89VMU4G8QVYfJD4ZT+zcgvY42aXeToQmO59+zZCg7Dgm8rPzb/Vgr
kSh4skaLuFfGrovfcluQ0Mv9rrhnpBlY3HJ9Y2UhjKxzRCnEFxd2XUTVNeYkFnOa
sqKk+RqX49c342C1gyhBkCGz74ZR3M3sbkc+HjVM0fCbjKOE4rphCUnyVb4spCJJ
JOvg5cQQAKqoYihWJsFeVEmnlNk1KwXKWDjH8BQcIIo5RVh5Duz/IUHg1pByLhtx
ozMgk93ika0KDfeFTqd+DxQBWFFkjb2axiiGY/2DA4vDr2CQd45QSrnj2MoHgtRK
iRmUP0WcsqSTUIOOGY+4rPuPVKVAzQ80ic0axIG2G4RNMTBk+9paqJTPHQkgyjmM
NkgFYKeiqnUVjy0vdBhVwNZYF8yOdRKlkaOLzV56j2x8O+YdQCju1/iDAfBdBphn
N94X7kISdTxlLgvetQOkG2pEp4eEqT0YX4d9U2KdTChJTIZ2YiOMUfff/qJcyeZB
iQqBNsvQRzAZzFu9IhORIe+HSNUONtMgT8QXXkO2IZqGKkr40OWT8TAfHjFXgo0S
C1ljToJHheFy3dMsVGeTiG5d9xjH6S3PdddpeSPh2WVCHheBAjaGCDZlgKLKwOhp
sli4Df2vab2Hlw9xm5s70IzafxGghSTPTQ6boO4hCViMAplE+ZEM4POiTUXZs5d1
kprzPdDeYFuwpSdrcdMN+eXrPowgrVYFZU/LU67+bMfYapa17OavFUcCFmnt0wI9
4jQvgSgHGabxJ3yhKtXVvE45hOo6vfl6N04WzXv5H5xYkowb1EhDg2ktQ4cCQx9d
nzI/hJrao78hHbhnCvs+45es0HWhrtdsqZKa2u2LRdImiiHwettyVatLwl7ZmjjS
2PACuXI/dQ9OPi/rm8nHYPdJL18CodkYvVZWuCHexTCPrM3nlSZLoLv1ogZ9nSul
Xj8khCX9XV3vzdV+Cw6JdbIC3Wy6Co7n1Gn6bDE+Y5UtoGOUwBQbjktn6NZ3ACkw
P8j3+Vf7evhCpLNLfRKojcpxKoO4qyUIi7XD2EOfwXXjhkhBKa7tXAMe011K2itB
N8H0rZ7kk0h3qbDfXEdxtQvnIabNK+K8vBLlhhN4ew/q8vF/nUmyqkDgw2ymkRIw
2SaqzOwvjLLebrlCyPzaOnbfxD7CC6c5Sb6feomwN+LsiS85uKFo9SUzNCsdbLAT
A2p3KA+o4Byw396MAItkNKWU0B4Eat3/QiadDPFBJ9phLOTRcF0n82qdCKrJLvR/
EwPGc9TvX+cSQmgCJSgR2jQAvIaqTbbanhnWjUWXEKHbcDm53EhfDyVXZ62JHlnZ
ssbIiCFE7Ynxeb8EJlq7PuqIIzSzwEDTQCcwfn1wj1f/DbJZKbFQZGcYoPTm8D1G
o6miq7d+yEj9Du15xAdO8Ate9AhAyitsVLz2IN+argi9GpMLQIXVQc5dK3ySExSk
rJZI5KKnqV4uvObTzi9PAq9NA1KZrxiRUUUEQe2GZmV81+Gy8Kz8+jycVIIjNtwg
83J8dv3iqNXIxyj7BP/UHYyOWKbCGcmdEAmg0WghGbo7vZVr253KbyCDlP3xH1Kp
YBO6iHT/7LJoGDEjn0wrhfvmtQT/1i9VgkV6EzT80zgKcZuiHfzA151o47KgLShe
ys6JW/1HqXj8GVbJVXmMs0uU0x3JOr6EmERPYZFNdeH9A4SbmWVJUrnN6xBK/MDc
NqK6BWVIZPGgTrHymx5EVUAtkDdyoEjgOxRCjbNFGKVl1Gda+x+V/Z2v8iHojRao
JmFxQGx9xQJEey42eLr1+yGlUpRQHc7pJ5l99MrpzA0LG7yawlHDm77HB9l3cAPt
fO4pnv9WrJwGZDnL5/uWgXgY6a9vHoDafkr075ZY9tfbyKM+5wV7KiWteHTSzWei
FJL+7c0/8+e7I4guIAp5Ilv8WYKdBWlHGhkTPlYFE8wh0OX3AmokQ2dyeB4T8c/M
0m9nigUUWGLyi6DLxA2Xi3EwN0EtdPnpt7fu5GYshejCCIuCX/2xUWXLHFgPp3gg
EH0Znn2B4ayEwegW2P5TTWgQqObYHdaeiUpKlf+2Si9S9kuCkvmbo8NZe7KftPbW
UpEo8RAkCmv9f0HzEhVRFE/kS9a7Tfth767qYcIYfygR7hcnn/sjw7cuPRYkp4Ai
GHuhbPmkYWe8M5JhcLG6e2oaTdBkQ9s9Xh5/RJhGy7QfqWQhUoT6JB3MzrbKZ2Ed
e/tV/TR+0+duuffzMZ0opLVeC2ZT7FgCmmv8/S9nDVA/kDWvEKSkP1/2EutHEB4R
sppqdGW89Lit+RgE4hdkRwD36dd+vab31q53RxWcnzz9D5LdZHgL1Wh84gf3GYPL
+dCClEWY5D7C3N+2STqexxtsQVk6g/PodJB78VuI9MnGrECz04GV3awiOBPMPwV7
8jBvWHjUEMi5VWOSCwH3laVusm+30xn6DhlpchlLQuWc3zvB+JJ8wNWM9DpoY6ne
crbMz6G6rvk/wJ2AKWsJZyE5p61Cv7dTa5IV/l6VbA399XSr8/YjaURqYw3f2KDG
OFsWFLUtTqczxwEjqu/gBBP+t21mIAixLgKYqS8+cPGlWpGYvi8bNdUdcLtxkwvm
MHvZZ3o5CBG+OXUVMK2NRRpn6B/SQswa5Z8PI1r4CIyRQ6WH3ZtbGBcx6spfbePy
9zu/u46d4rZLemSYZyHtmf1iGMt4XeG73Hp/IRiifkb53MI+yKQL/JTqPBy2c2Mn
c32KxEULzAD0W2hd09WGTJpgniOx3Ir2iscNDMcuaFR+eDv9JQqjXpuh2UJoIEJ3
6ZxokaP+qi8YG9cUTev3SZi34I81uLcHSj3YNeOL73D6rdeLAMX+nVGxhzmnP/Gp
+5tPpUMh2t8zHKQlJ+G9eo5V9fvBgig0mutHO4LT/CynQvliqT2nLC3aAdQguRQi
UM78j/eMwfM9r/syZtbENiuEVA+onbkOWTlkm62cm4SI4looe3MPxHqZicpdY4a4
SjFkX7ip43fLCxNYxVDCX+pSRsh7gTvI72jWgB5AUXabTIBZCWDlQR9iDWQE96NY
oi+K0gwmVV+ndlY79QABTIHtUoKBS01rNUJDuLP7q6GOLPmsiyrfg3ezLACXXcqX
wA2B71EYVyPVjoXAuuvJ75Qcvdj5UNT7awi8CTn1H6bc4kzOALt0EaXNsn+f4Jm3
NTEpEbYaf1v317JrbUHQ660oxr32okoGzofFHXwa4WTI9nTS3d7NneUjGkQ4o0xS
DSzpRxOTqfhhbixlVhhtXiVChhnnIpBE7YvTbBvmYyQyQYZFnZPTaApBnzNVXOoO
xD66rWNTx4Y9ctvC9lzDCNpCaC99kCPV9mISSgNn2+ghxO915eEPEuD3n+kGxuXy
aB3pvzmcuhyDk/BaGnIs6b+kzMQThNqbEzP7mRF+avlakTO+dS97CHeAohqMuiy/
EyOAsoKwDEciUPH/Wxn0z6g6RGJ+9kxja9sCZCyfJnfLVdBHWwUJQi2+qGsGpXGy
L8VK3xGT0BQK6rt8pUNl8S1UvyKigTBW8Dqerzj2pHwTEjzRWwYPJl7Z/SlVM8sJ
bM4OfPWjfFgXKlOQr0y/WTy1nKXUde/cjEY7C2ZrgTaBIMoFyXooqCBstU10ul8+
naky/9GamaGSJ51A6Q5F26dCQHGFxmiKeb8Av3pgIi8zLeJ3fGbwrFpPMid6W2CW
83rkIlThK8vVCv+fnE03xZhig0nHcuvtSPaCvzFrI+Qu8WY5orLCV+SadEaZAic4
hOd6poQOeRYKyt3pZK2H+5hStNLoLfDdxr0C9gvA4KHK8Nw0ke9NHGI6Kae+Gnuv
SQxItMX7MsvB1tkS6eIwWKGikja1U0gYlnLS129GQ1aHT389U+jCDg2SEYxvu8fM
feqA9fwp2Ppl2i2B0f/5MffT3G7wV119eUIW37XkCTCqVMY82e/Bhy5tRUfZbm+X
gET0v5V4LZLP0JCvcjWD2g/zLwtBDvXS3ACsdsicbD+mNJnynYnhoh7qTSjwqxSN
TAYXutjwoRCvspKlyeBgc1bnZ5YV+cY93nWSw0C2Hk2Eo4AZFhzqXJx5FmJkc38B
6os1ToUSxGbrVYK47x6E43Cez8JflwecEpsk+ZRCYEwLdfxc8hIdh4lOOVN2A502
mCx/IurFsdo7ufcSYyUAb9SCHOemMC2O73z+cDUAPnNjmOoXy6DhKkrQkAzzEA/p
j10UCJtWmrFPItuKhodiA1hb93TAJAOIXdmqQoDNA6eSuJSy++gk+aXcoYL5rKcX
MwBWoagoQUWYAMEzlWkR6A2+o+iqzficBjQttOdZQl7Wck09w3gyCCJY/n8CELBs
BFPR825aPuCXHMoxm36pc/yhhPAsQYQXugJzf//Za4kSuuD8KQZY4EN8zoA1Xyv0
es3I5EpMaX0QfQAYR8qFmyaGmrFSiQske/KTNzufTNnMiUSadB6hc0rBmnLVY30W
Neczm0NwxIdFun9OkbMS7jeqZh+TCjX/iV2v4r2YhKVnhsOX5xwlyph2Q3ilcoAB
8CeoFr4r6p/PxccUDJzvN+/rbQTSiNrWELJziNAA+g5HhAIn6Of96tZY78+yxA7E
QXI4zsbqSBo6tgviTYq8QcqRpO3Gum35Fhm7Qz2uVCCxxWuYpq7mPzpsbJtHFDp6
LyzXnnMEWeApwWKLhoski1Q7H58XJjrTR3WwePulBnitvzVVNKfAzr/V+abNWr0Z
jyFqTFZ9b3xsKM4vWVhxggha8ZKJLNFdPcGnG4tl3qpDoNJ8t0oGpmQjWO7Si28e
CAMK0NgZOLZk94DbXGbpw6WZxMuWSFAinnkLvqtXaWCM8rfV/BingHkrF4LZvOq0
rSf3hiLjVsMbyQUkVxuG6yhG1iQNZ/kcF7s0cL1Nb28XmPDtRqaUS/9NRD8R3dSx
g7dkZ4XqiYhqavmzqj6tsYMOWMByJKKOq++LRIovq1CYVMpYip7PQsZB1477r8hD
OHQz2I1Vu1sPTZ1UN9fedRFHwvcvm1baQGShmpoeNpOAsUHi/nQEH0g5JeBUxWi+
6gwqwRMvAjffjFSZwD+hzttLxBuK58b/8e3/l6aiWFE4W4kMVarDFGR/qSdKAXtM
hJ3b5MiTnWDTDS/26tWhcainI6OrCusmjBdUZiP/kgYSlEgOuNdjjrt42IEINvd5
nJ8+CumDpYluaKfjwKXOMHMaxIt/GTA77pNiywsaxm4DTH++iQ2lAS2/4sapvUf7
QLLFoZ2I6tqnsos6k1Tn7icE/E2vEBETBnkV2zawQpksKn/T5u+dML5sF7vcSXrO
0iqr0C68E5S1FPH1GBdI3TOGX3EmPx/6pUk6IE496G8XMta2bkcUsCNPEyZCdK3x
jJrkRWLUAAyazV502ZqJjB0upy6qKE1Mn+tg6VyLEiYl9FXkb46QjhYiCtGQui9M
cE7jPVBH8vOKHXxwSqcmscrXJ6Q/IejmRX6Wh52ixbgmYTg5sz0TS2KDK37KtVrn
2GWcUx+Wk7wK1+RbWwOR0/W6u1RbxhsOUmFJsG+Vs9DJjDHw2N5UkHtRYZMF8gFJ
SoNGyqt+m3H+Sd87seAGzEWiBF4awPAJ19KR6OzaMtJm3pebKiK+JEpvl12FjsWa
+ZtWYSQRwqLdiVEKHv5rda74PvUEbAwiROcycoxOCedBjRwQ2liwHGqv6dcyYZ+2
TqwZWvOcmXWGRhWTsv/eQ3oPS+vzgNe9Ym6Ty9DbfqQ46YwjI/KtW7nD7+KtL9Du
49HVKLNOwwKIzK2B0agQx7na26EqphhBA+nDs7suotOU2H8ZljQHg5h3qIDx/iQO
qUCOKoJFB5Rt7LR8Uc3ez0xigDuxor2DBNdNAelpizUbzN+eU5OUStKNR/QfdoUa
rCaLx4faxWUBItEChDwAT+TFVpzNGTF5MRxcxQrqn84xoapdcxN4Cm+5v9wmpuGG
bwG09k4+Xvtule0FS0IG6LvprGJWsDSShev4td6PM4AinDu5pMqUVyOFdpL878M8
PPbULc8kmrzlbYpnz/o3DNzPMJk+dGww1vZlCKF2E7vRr/+eS+K23cyCdNU3oYPx
Rwc/aoph9I02g1Q4VXE6sqm9mskBWVrOA/OCcztad2EsnKx6rCfb5SU0hKod9VQv
+Wat6f9TK4NNEouUAHDETmTnVcSbXPEfm9ryh1B34BVY4L8Td3ozLajwuUBhtMPb
yxdrmwcPFExQYyeGeVftt8T8qC/rOXnu7x4iZ81uPeLo8l447riB9yPrAXJ/iezn
LO7sG/P6CAP6/Elabqse9oRIQP2i0MH46QepAKNmKNeSROHw01lJIBcnAhk1jeY1
3lwYf3kuy0oV9MB39TGowO0vl9V9CFg1I5dpmZ670c4ub9P7bVIWQIJ+IQaL0QPn
0VZ1imcIKLQjgWaY9R03uq93znG3tCpJ/DIq/Qm7fL3hFZHfPOxqfZfaPbWc20Cs
bcVA9lkKO4S3XVVFtrAZ20yXd8Qx0p+dh7q3iSK+AY2KDPAVyKzyEeitLxWf4Xqr
UDWyNQqhL44j1myDhjSH/804J3LFgzMyyH+7avsBasCmAyTor1sN//S3vyOog9Yi
uj09YKSFnK/TRXSrAY2Hu/ypnSycy+jPdriulk6RCUs3H18W22f/ygW97CNeYMZj
ALTmD2ID82tp+outy3s7RZ2bgooG54mi1DGCSCDLxDqnlLnBm0J8HECj8pavvQzS
/p94JYEPZIb7abKSNPFxZABf+WJ8UnKJeKuDFzssZIivQm6CDb1fAZkUbb2ltQcp
hwuN9arprEGmDFHoiDGvD0jXlNWjzbsdF7shLcSw7vVH2Q3+A3WwaZ209CxE4kUk
kqohlmiWzyf9K7fD2OYnZyc6D2AEoba4vERbylgXe4jzrqKaSdaopqPyqDJJtwpA
L/FkZO9ysaNWD8LfUzr3MUjA0gBZ+p1ATCBJQ6K+dYH06ibSMbjb4qtsbfGEtKxn
43ajp9tEcQm4n5ri8CxL0uyULybMpnfGzg02DvcRrTOBo0z3lbtNg6gc6bd1POqA
JpvuZ72cG8f8s6kepxrA0o0vKZKx+m+4B/YtUQ6uT5peLiSWZuLU9gYHysL8xRZR
joAa7ah3F7paIOhRaQFUOqDstdEUWXMg1vvAjXRraAi3XSlJalqAjrh7i/+YWvhh
qNaYo6b8OIWkgViVHghzRWy2ouS0MGNA/Gl1GdnThlAcJohSk+xiU36p6D0qI+tr
sxuQCP6OU/XobVNnO3z6wJrlDqEiO9953NERiHIr/QOppTvKbpXFcqBr6yW9Cd+d
KQghyDB+QnPlzmbwPYwGh+JkU9qwih8ansl4J1gPgbYthHeLETMT/DNGbn00A5wM
6gF41DBPqx0FdnGnCjnm7ZUU6mwQbef8wod+eTNY/E7tuIB5gUJjlx4wD/84LQsR
8oDZOiHFwnVXs3yVg3DCwgXgTR90fEPe1fDEip8c0T9JVPCyFiFuZ66fdQ/HF4L+
1x+7N2b+CIVxDV0A5nYpy0chg+wv2wPyoJ6fyUWZ0QrLWFmRI81whB7uaEwyXa3E
N0sAUcNAAhUzHHXkwQvVXTCAm3Yk9muRzrPIrjc0M2NtM4cprpFopzlQZtC0lKjJ
/BGyzXVseWKRKWmcHW097scFnTcTPAAo0LV5tGaNODiQV5v1E0/drJQPAmKDwzI1
6608d4pF1u7Es4TVqhQa03a6NI2SI13ljb6iaruNZXaGH6VxYAXd85JGU+Fv0knA
gD3nrMf0VB35c7zXaAc34PT7NNmv4HqfsnMNcipWLjePwDNs0/LR2XUrJTcu8+xs
d4l/QviP/g4BayMeErXgZwiyV74VPG/kWufFgiU3Y1E8H4UTjynpBC1iNYeK7Aby
niUfT/o6pKuagIQCuF/17BvRdEiKwS5TGU1Ex8VrzFhFQGQAzV/EWTL3vfgIYJs5
NBjw0rQIhHXs8dvhILjKKfvuza5/RGQ1mEuX/ztbt+rnHhta5jx/fBn9Ki4fjquG
IjOMbncsZ4nNqjmLrqZj6ZevHtUYdIRXBFBOwvzQ2GuniKw7I8oT5mj48O0Moo77
RLYrADD1RCr//jgGb7Lperb4sEEMuelFFO67d9sTlQTmpVE9okjXw4vYViFslKd3
wjPXa8Wjaos1I1tu0ilpFJz7ElyBhYljBBOC1HcLB2appf3w5iOP0xFdZctIjpmK
FXudBI8xzTjYhlUwirNm/0aEhkECQCH3Yc4O8wi83ROHnSdHmZxMcyRvMLFmnSte
agD11RcbMAmIue/c88qszZsHwcOWo0tHwDle1XUe1MmvrotlEzrqvO9zeepUpvLt
ZTKIxOkBwp3lteix9rlvMkQemBmoWs28TqWFG/9gGwDyrL4V+m/uaWmjKEMXpSIS
IArh1tB6CXW4cOwJoI4Abs7bwAjKTMLtr945YqF80R7EPpI0JpTv8tThq9xy7kFG
BOmiZEikN3GXd6ZtweACsa7eLKkMJXzG5Yw0kDFqXKf0sjPURGRyeYwOtbnsxFpJ
pCJN981KQ/ld2e+WxEoq38iNvnzhztSFwpjcrcxwG212P88bZp0kNaSEudjpwrKN
S8uzqh6evVvJF0zPzJNolPfoJZPLWlUvK+gOjamb78FKgUFEkcTZLRsYs/9xzOTO
n9/kM9BHe2MNosHNlQ+QGyZOwze0FXvF3k28hjN5m2E0Nz5+t2LmN1LP2JVV6jZo
e9VdU8ZV4cxptcg85ODruz54mSwOundscqXC+9dZOU4SN7opLGnRIa+EGesxAkOY
sVtaEoPlBz5dzM+WRSUj+rAs7/uDZ6DVp7hxxAHxVZXtLiePq1P2wp1dF9D99dAX
iX4I6R5gXzeKsSrqsSSi9LDFnC1sr9NgWBZWMU6elngO3PWY26L8bpGLgXZE9Fdn
elE+aYEViHN69nAMVwkBZ4aQAjsSvXjvu23OFnIUs7ApHcSg/UONrgsFYg8Sxpby
sTKHJFuv2sQVro2hpwu/9xgiGZu+r95jD5K1VeR25hZskogssL2WV/dW8/smK+LK
b3fkmW2lNduIySTXzEDB6H3+iamS8uJrmvqEfkUhEGsu1/fPMTtQwNwuGqHZebQT
3McL/kavsX4xXWe8Jf9mQU2ea8ILj70wopnlxC8WoaSd7hQcZM1k5K6Ea+bHA/cr
zQu4qWXiMBxGfybjico+ZGJuK+MhOYjLNoLHH65owP6COU1JjMQY3wkQ1QDo40Rk
sk33p2ZPLMUoXChoyUugrKZ9/WQN/nc+F7kUV0EiFt1RshTU9qmyhi3wHuXhLeGM
EWgdPTYbwM6oC1fxKI4uttMn4X/j2ZRDcMzXKU1eZEFEzhXzSuYPwbgIKL22NiaL
AR6BMYmTfobtg1eT13Zl60r718oXRhXYilIbCm6xBROghIzme4W7uVYOqpMWp0q7
dtpnX+r+hEl8iG4gCO4XJGcqh0OIK5SCpvUDNGniNGRCiW3unkGN5fN2Lo0Klu/U
JNiPTQcdcf26ejBgY4lDCS0KAvX/GL0gtUrBs9TWUlHFu8QYcg2oby++SOqhi1db
mXjBRFNatgx7aabOuoy0ich2VRAw/G2/UVneLPjOQvy2H8KOXMXIpb4ktkzOHXUx
dVjij49mCW9nZk/UpbfQhVMMCn3cV71OnIbihB59dLbRA5hx3eLsHLsIuikdBEkK
qf9M9noa0P39S6ZDJzkGG+IZy6wq2SeyxYdKl0uovp4W4fAWc5lL1xXNNySIvocI
cU6zQicTeHpxQVwLx7vBTdEYo83nvtI1NXI8uJymOGjesuhqZ9HjyD7QlzSz9q2C
33hSy174Y5jT+wGgri6KnRdxbagZidHu66UFbLwqUzAA5Hh9Lx6XXXZSiKDu+ydl
Ddg7RbZTX0pqMRZ1yN81/yln8MWaQ59H2mbZvYN2kVXxanw1/d7OZJOMc2DtZq/1
BhfYRsujhUx3BSBsSHkEQMHCk/fGJcF0TZ7SswMdgD/D0gNH4GZh1utiZR5sYCxZ
I+k/l/Dyldq4mJug80BgtQwym735pbaiASLF4fHPytGVaPKXZYQo+44X/JKjlsw0
5ImsecFxc1n5otsSth1iletCXpzajyIKnPxyJXVJ+5ukBrjDICYt0ejMOLwXJJ81
XhoeyOoQyURsK1f3i4VvYIpSicUKA9f9pq6mBK8Yg8QGQrJfaSn/ey5KrLQLm49J
ttSHctE43vtcvGvom4nMRI4D0tPOsdfL0BY7HuuQzQiWXIBSgv0mDTadnGza1cmQ
LWsdfLiMPrKQlBLMqJWyzqV+Az0w732IQhjFxs5sm/uI16JsoVviKG7Tye0SleIq
7VRzF8o7AKX6RnhXiSLrHHjwdNcQduMYWEYdJt9WLeyd7b/J93VHdcpgxnevMk2E
/2JQLcjIoLPbB9uc8Kx09wbWqMMn2Xl09a6VM+jyYp7L2liCFmP7TCk4sLsHdje0
JZG8zUIsiODrd2ylYYADk94s27DDYiMwYj93ZPg4gBAcSYAn08KAAE3TExhdT3bv
OhADIJpCFPUeuJCzuhZnRrid3gbqJW7gL1/6xc3KKmQk9LQUCdt6Ukw45iSM3QV1
2uT8X/GYnv5mywsN5ccAi6Bw9DIXYPIpl4YsA8naapdOk5WXBwbUvC6CIW3AvOQ3
RofjKoVoVV8Ec19k+To246tjzL34zDdLu9rN3FCEZNpz4t/FFZ6z5xA+vTGT7kc1
q0LP/2Jm7M/Kxb3wZSakx/8CijhQb/FytCcn15jyqBpDYtC250SeEZFP77W8YaoR
9pX+M9wuF1igDrc01jiZ10j+vhiGsp8SQVutC9m7oN0tkhGMwGaYbAMQFqp48vp9
U22mltpUZWcftddbhKRw1fLIhzejfOUNuSfMvEhvRQgvH1a4c0FWqR82rpYrtHcm
d+K60lybjbGqJkUpjgrKeOQgwyhQCB3X45rt2L4adu40dolX9gP40Ajaz4wH/qpR
VatQF7qddScSaS1OkOL7Hd6VllqT0f1W55g/RjkDWMdBjJHusrFGSbGWpsIR4THx
fka6PT8W1Z4j5OOecgJvdO/rZexix6XJUFq0PI8B2HZkjlUFZgcZMRpRLA7bQYjT
jKqsWhcn8WwU5bBzH7E3ydwOkHMYuWwqTDS+NSPHtzXf9Xnxp4XHmxZtfEde5w5w
sKQP3MJpSU8XoSkhyTkB09W1klc6qul5orewcrfcagPZ48qfnSncSuZGf8/GD/0K
9LAb1ZgTcRu0qK23AlFKP0CO+TqKorwTM4M6hggbJdj0SRc3ke8b1HADi3nSDKtY
lrZPQA2OM0fDHQSynTD1Pu6F9yrzfrRUfar1yyHdjdmByw1eWrv8Tk+UjCHxJBzV
RIFyfS1OYfk48jpkyGtBIWTaK1TkrU2osPr1G0m+sXAcstgevZWTRfK1wXgEoIjE
azdW/K/qShw1J192W7XlScap8YZ3IQd0cCL80KEy0RCZBdngE1OqbyRxd1BSqzIm
MxEe5SOc1CFjitVDMOGekn/kEs9/In+zCvn/5Vv5nduuBmj3PZqzy3uKtKuAUz+7
GORueo65LBD2hz8ujtWbM7J8oiunOEuwxL6fn0xHLMOdWud0HBW2sD9g7OmxmSoH
PWW2IKlhluDy/FYjU3kNEfKJRxb8c2EqDmvVYRaC+kWGxXrUkPiogMcXtjaA+4Uy
Lgm93p/SE+BuXXNVUzlj1SECQJFSGNOjQeuGfABPU6hL+7ujCgga1SBKXnXEvfFb
GgubNmNqZGuXbVV9TpCy7bRypusKwGTSrlw0U0h46tL8Jt0YaM6V2FJji87XU1RW
3qc1pqv92smJ80v1Kb5vENlEwRPuLTzr3M0UMH6RNFneyrcI3nBQO+0Qckn1RuWm
RTumkUEbarMbVKka6PiXpTFv1xT1DFfP8TEgCgdL3PyG6oEfgQYi/BW822FM1i4+
rzQYGZyEdpSXvAFfP/5e5BuEeev5VCmsh6qNOfWfjNnyhMvZXM5UPESNteWCYy1D
sAVvJzm/hpFyOyKpfL3uOxwPqoBVvs+PHySGtPRl6PhFuRW/ckJmKlaPXaXPtW8z
z4du4GV2K8FGLRrNVt2F/t1FVrgNGwTEaPIFCl64wiuwofOUF0r0LEGgwjyQwgex
ENANoBp/3a5hG2hc/gvwlVXUae0OgXU431G6lJJ0IlQaGfzSuckyzrYtwQSdr4qP
1Fv0gFzgg0yD5YKq8/q+mO57pneLlnz/ARqH6Lc6gURD3qA0JZq5b6sb5ZNAcjEi
PmSyltXyEOuWLdlfFdFfQSzsjKyhdHvU0nd+kwerM9KjTImfU6y2u9tmyc29nHkc
ioV4v9Vfcfd80A+u4hiUQLl47RFki6lCpvcYuEokgKRadsC1K1FpANyl72ywFbCU
UuCjcnAVl/wpKV3vpWKtyK+Ev8zTsCPpht6YG/vvLl/UVPGgEzCbMGVwmd9UqV1o
nSMzfwckEuFno19mGsQpEJmCwi9HXjEzSL7g5UKLJJDBBoDPjtGfMjAiY5d9HLPY
/d55YK36iCq4N4OsTqTPjuoHkC4pbFlfVSD1mYwiej1nsXpvd88FsyPQGOE6QeMW
/58Hsnhnblh5EzsmIAlVr321gfxjG1b9oqexLMxdL25lmj1Mrxe69oO0wNDEBUdv
VHaiBoty3CQ3akJMv4gk2BMIDuvHy758J71jV8vzMvo+zVgiTCZeJsnhx7nrWQ2h
en7ihZFOpv/HLwPPhFSgiOnC8sZpqpGWiPDJfAfQ6c5AqGw4H63XdTBVw+FL3qdj
BgmG5LWTF8JmojHxxiH1esXpWLfuv1I5YstQyKvrBmvXSL4Vb1rqwDaHmN0vRhFr
ILa+GK7cVR9/L/a7YgW5UyznsjZJYXxQIa4yMTJfSCRcFvl207/pjRCYXz6ZcHip
jtUBzPH1URZr5IqtHAQvavDIa2cL+vth2A5f0mCWPU8wDxhLH4stSjYpIgrElOxb
n3o2fHfvNZqdxThUBk+OqhNoYPzWS5h2EP9k3t3i++Z2SKWJYaVYmauQKEG3UuXj
ReEyoaQJv3K73D1+/mjCy175xwN2RhxLWo1y6oERiSWeyzvsoiT6EVNHNYQ9KQhF
up135EVh7wpdmec29Y5TK9Ul+vtfb3gjQVPYhcbammb2ky/q+WtpEfxvdBjs7DjV
8Td9QAIt/cQ92fwt1D4xXZiWJLcwlFvoNwg+nGrYgo9YNy4lDFcj5UEn5T1nHq+L
Mo3ZwON/ZfSrSSsHWkLr+n32OkKcfKSIrUECytSDE1QHlGi7eQiGjuxUTJ73BYJ8
66LhGyVC0cysiBv401e7Pzfw3n2QEp2WC+Vi5+wubJVQn/D653/BbTqP1j6GLm6q
/bngD1Dn7CUYowsJN3i23wqCGcmb/VuZht/cOQhdsR/MmE6J3IXHgjLSC833E4SU
Una5bxxH9OM5c8THTzoYjZ9PqlazvE6o/d668MyWKMMJO22CQ2YPqyvNoblUzklL
OOaAfrg++iOcTF6iMZbWbTklJNk0g1W4GFdPE9cTMMQskZSjPWebApdqMBuQABkf
TNN6TOHdto3wAf18RKRatMWIxPvzpoXt3Dt6WHSLWu7ZYKxtMpxtuu3Ul0b5qNpC
DoJBjfcE4Rkdiz0gjx19zUdDZLmV7RQGgvT/phAq9i1LczDzEScjW/Z9ZbXl0Ee0
ioZaXKoZqYm2iwKRtd0iJRHlFyz5++QVcwtXYbRoS4M=
`protect END_PROTECTED
