`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGOKiY4X/ndhXtngG2MB6r7BJfVQrxnyQ3knmv3JU1o29baeMwyD7kWFTC4ERezL
yQ2OjUVANFX2L9jXRa/rAGaIKPE1n+acIclF5FqugiXLGmnB8i7AimzRTDR/5X4I
CG/rv7H87WKXsHvA35qa3yUyhuy0pdpNmYDWubNtRg43XUEGaRpvToNBhei4WEX9
wYnIKmrFCI9h4vhLbG0SQS4HCfBCUG3DWH4qHlpu55ZIB+YlwPFHIqdLimMk2JQQ
YDLcM2BJrbw6o5nc69iA8EjLXe6U0UUCGmagvuNHYlpZ8KqqelTEBajEPY5WoB28
El6LtAaMVRq5WeT0Mc7HuYZhyo10UK9UIA8IjKfAtRHXSio8LouzKHvf25hk7oqI
WS0GU2lV5fFfHqLSUNJL3vX0rFfidT5LIfAlr0qdq6uPi856JyUpa6SL9TruWWou
KfBv0pBBE+ZrExlnfYPIZBW2xW0/NfU2PSdZYs0N+ezw6aPUj+SWJqUvkygCz8tn
Om5o++fd29/VO4pcfsKYeUqECkXQGVacOrKkOjRbqIQlBRpiMTuDO7V3zYqWva3y
YafJXD3skslLrMvTrSN+fK9bmP64g7OqRKGpOt8BOi5Rus87MTcfs45UCam79UMV
Gk+sRDaHBqbSWpPSDrKn7dVadRkFU2/rwQs5+CKuqIlOxJTgM84kTGr4OZIe4erL
Tt1Ky7LJj9H1zV8qMfzWwFTbyOkRrIyb8DJE5zgbbjdqmUFm7nYGOZ72SS+WHk0c
giKcNLA2oQCO2RWLW8HuTcCmQscyZa5ceQnM6IuIJfXXByp7SUyHVvzADTpUVZGJ
dkZFMBrpOKVkjcEIyWN49PZ7M5koi49z7nex5tFRUun3YK//Y+6X7anyZTJYemRc
lMOiMLC+iXGvqKmXKq5+cDs0IW8zCbpWmcUBwt0RUtXWXUObLwo+2TqEnIEmmlYC
td7pYxZKNuyK4CxCjd/4o1yQo39Z6SEpn+cZKLdM8O9WfDJljr26zglE2qzlViWV
kqgcMpLDfYsCPCqy2GWRcXMxMQVzfyhyrX+V+IGNkXwf4zKocnVlIUlJSCJTt+1h
SBk/MaXISF1q5qxyt7SrEK/pwDvf7pDDgILk/S7sq5NpBl+KUxdkkXZzotEO8wqK
1DVLWC4ZkWZMZ8ghkPPtEeT8kXf+QchGlP/EAYCMD8ZYH3AAvTNwy5IofTCJeJBR
S+oEuhqWmjBw6CIqvdXdDr4AEdluWhYpQE7jrkO9u8YgfuEE3stNjJaTX6/9qGdD
7pLpCt4kCcWgfXOGY3kOP5B+Fu55fpROWL+7fvGQmhtXxI/Auyg1378pc1h+wHCd
uTlfTUruNE8B0f/9xIodq3apqTgKQMTYaZTXysHxCpXg+RWZmr5Yp0S2oMHU5bBK
/CVO8crpgT9P+0yeF+EkOfE6M4KyEfVgBnDzoZGAw7OR326Vk0mfO/MZus4OvwuP
Qw3ozzu3s/EOLKsq/rukIvccKjnh31FOegQVuHME9dEFtXL7SXlvRch+3A6vV/Ih
fK8wJSojxOgyL0lTAUpNfUh6xTtP1C9VEhy+MmzFYKDFu+Wz8mOodgCjQF9ldYgF
bpIpNV5fCqefpUM+rUi5Ip0vczcw6ObOHW92BE854eXbRaHhHHc54C6QrYwptnCV
iVJdbOQHCH5PVFHmwdKUXkZwJlPxrFyy2ZqR8jJmFVv6I7tiolQYw97J9dslaPT3
PbiW8s2WW60lqmOZA/CS4buFJnw/Mm6Ajl1joy1e3L+c+a8rLHKh2XzLo++b35of
Ilyorsq3c/7cHPSlJekB4eE2UGxX8qy2LLaTsl+aOGAGVRzAXn3DbQepVzx7wn18
EI8XyJIZL/SyFuiuRqJN+rn0jP6pRVWmiTRTmFZ14jZcdTT/+aV6EeoZxUKHu/p7
xmMTWhCubHFP+dB3w0RX96Z2MuieB/JqrlLKErWuUFE76xcIDROoYYDRsxFxQMwW
eSTHbsKYTq81XqxHMksCYeBC0dciSIaA0O/gOeU9u8L35AZROPrQVClIDh2AySlj
8nTpXZy7l8euz4YO4+Z6faHkMm7u6Fv4tZcQPnmJ+6SIkdXVX/un39dvBwHySo7o
sA5b7vwjbBI3KowKkh36uFbylvXswtqnjtToEeVy7CUlYWmo56QTIKzzj7BsqeE3
DvzOfp4NOzep6qeZHyIJsaL5/J9MHOiVXYK5kEmTp+aC2BhsaITmmZpMWtEtqpFH
GVtpN9lGrCUSmbrUvLr/yka3iaBg7x2aOyIq6pAcachCbQgNbRls/zD/pZi1WYld
mpQixfiRnAmx/LV9W2C4NvY8Lz4fbXp0k2DK+0HRApUq69IpnqZ1OUnXmrofgbVq
+qk6NHP51rcXFtm/LStwIMkIKVa9TzlbE+KLHWykSK68greWZGYN4QsdX4oTlFfa
8HYlL2MmXTEHGTgm5fWxDqs4djJGpITJcgT+XFqRCMgTI4cY/6mfMcqPJcJe0GZI
NBnJG3RgL0YtEFu4acSfvyxrEQGTPysiIhf3xhCMfnlGLQjnVAzaD1vsaazGyN6W
wIcYuPH1bT6jrIlhGeYi1Q==
`protect END_PROTECTED
