`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aGl47fJWh1W1q8Lwim8zC3uJIUEK5b6i1Ql4DRiys0wWtr8uu9p3ayn8fqEKG7av
Sp2Vvl1xknzTzONCYfwEjLDKRvxCh4vR7L9OmsFYmdQJ/nIfQk28Jh3jYTaXqtU0
/a0KKLl8wREHjYqg4+Gqe1hlA/wulAktq01aWLN0+TOsTq5C8+GYpsK+7ZRCaB8v
tymqh+YShRSlsQSmpbQWy1k3Lcmw+9/KpH4YBG+PtXlKPPibyZYvg354OF4kQ2+4
Kje0xl3JQTe094pJ0VJCnOKBJverknC++mhmIKpXm0CmZglAF+fEuZ9rik4an1mg
iDxF4vL/knik4vrXahZW6aaWA8a0ZcalUmxd9wa1FD1ZXmJpCn8nwZ6gN9SzXQ+A
ts7xDihzgSq1LzGhOWtG14pw2hOl8LioZnfxwehI3vWZ2k3zKDtVQmMstMKdvdT3
p7XdOXmqqWWDAwf9lAeKWQ==
`protect END_PROTECTED
