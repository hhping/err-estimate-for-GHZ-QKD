`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NchLhcbsPaOdaAdLWRKl3pF9Vktje+32E4mir6/7WoC6dhT2hOWiLz9RIz6kZA3r
2dosbvY4izNrpVGiyNfcbcR6IsCgN2v5Hss6uWyTqGC6rmHJeRehlymgSA8qzAdn
2WMMbqDes+pO/Aen31U41JC64c79IU5n3TIBKyqXiWWW73IzfE+3fNtVIjdY5YBN
E6PeKIbab6bG0CjXtwiUF9pOKr+Yn9vKjzTDXNp5eOXecUBmg4v5ENp+ube5E61y
VgKB1yG8t/fUHGaLj6wYjm8el4gxMXEe2L9c2JYkM3toseZnZmVnzTrtWPIMk3nI
ftAzxOQ42vZ/Yb44QqbYutP+FIMU496KjQI63NV69VoaxUTbkLgfgFc7/AxWeHl9
6qjU/lH8U/Snsah4/EsIkLa4uvr+lqwOnQqqNssAjjHvBS69t/joWqgvjW/H39V2
ktA2EE8jv103MXdJFzM4ZWNbx4NOlOWwPiFs4/k/gRhvtAYY/okJzas0faEJ/WxL
4/sJGiKNccTwEsSaJTPHunA2SDFRMd3Oga5zZh5GheNYkI50fzuEzUbX7rNb7Rte
KLGqXCrWSQPJundSg8QXB49VnGSo3yfwUF7WCYyYqt+uUz15yG6UjyfY5ofV6NNo
VNcU3gBq8vmpSOPxc9ofsMzKGHGCj39A7zxVFzORDDZFsTBZUcwa39qLA99BrKyY
Kj4rc88jJfjlJgUQTwx36zLDZenJuucD1K88aUNl7/JlfWwj7pw/KqXmMpQnV00H
PU42y66kiPm/o0FuTD2W/D1pW+PAMbho7ddE9Pokw63KPKu/2asLuqcNTMJP+/Z4
4rTD9AxOsCsexYM3k21W9k63p7GwXoQX9fhA2v+SRsKl4Tm9bti7zrfsgTTFSgWw
F/DYpMTXHItgL7gQ6se1M2z2XTDlVhuqkMfu21P4w6k5/u0uajRBBDEvBeaMEZCt
kmsaqLbXSUj3JTJMEwYD92c4GjvlilzR1aMZKX6fW837z0e84bxBHbnHBuJYTV8I
cYfRa8aChHxNl2+krSya/Hp4wPaT7CNowZ7azhTKBPxokCpgR+ifqGmPaGnws03o
JEewI4Ij4+8DDSwLjC++JSGgVG7bmsrjslUs3OCjSVYnLk31NonsOOItGptT6+xB
MnVbNby6rk567DzGz2Wr5aG50GUPYXtaRYUCwBkHO+w=
`protect END_PROTECTED
