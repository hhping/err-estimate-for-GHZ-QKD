`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98a4EkJUBbsOEFjAhp4m4xg6v7ht4NXd/pCAZbW25ShY6tT7O0d83HH6Gt+uLFy3
NcNh1lkDXrgEQzSZNOFo8JwKNNODa9YYHRTEZtzeZfLSuc7W1x/qZgmF6wW19gFa
XL/miNwP9ZLFrMpXWBNZHvW0Bh4JXq5EhqrW/wGqnIYhqmuSq7Ofq8hv0yYXMNZP
2/6IM51Bu9dsLKD1jXg6L+qJIe5Liw0TuLzx8HLyHM3E7LSq6Zi7ZMC+cMt6pls9
uKzhwQcLTSe49P92cv++9vmX92k1AGZgswgEBByhPTmJoJ9/GKNmkcL2toYIYIni
dJq2QBc2tlV7zf4KrqgPe2j/ZCt1NFKZ2bmnQhGQipk7bJFT0hgHm/QGj9tqlphT
l3fTJ7yq30iplr6wynQqZgXAPXT5uKxgRQ/onBz0IZhMvwjKDBv6qoUuBhH0H3Eu
4IjyOqm/vC8hiiWvakP0SMFv4W9jQ/3l6Aa6zFFomSPA8vphd6EW0pF9L2XYuVF1
oEVVC/aJRkTv/NNM326Uh18AqA6bAGtPr/+8HLQWV7kmtxySTxjpEwqQkK9poI/e
jiRpQPpkiTC9XBgt5TC4d721CNVuzbYfic1o1jQgKapKXt3Tcz/xLJc5kydELzTF
i4+Ls0DqMi/8gaZatu1Oc1bgIe+CK/hHMstJEsHhSlGwwSIwlVBG9xxAFB+w8jeN
HACVYzm+K4pw3JB2YLY1CBT3i9kpFvl2qQMimfB70OjDtZ2M/9ck9QpFW+YGYrww
S1lfV2cM+MVOi6XA+2NPUzUptLjOKi605E+cJ7u9e4Hd6OxVhOz+uWxU2ET6TgH7
jx8BwEGe122FUBz83hOPAFKWlNVzqC/i5BID6aUc+XLyIpr/wb9fyQAFJW1atnBg
T9jRevcceHvgreCWduYJOc3wCaVTYH1o77Q/KoCQ/SpRZSFJ+kZPR1nrNbx8P9X1
4FbL8qt5sNej6wI3Q213ZvDkHoF9kIMh8xEYcHaEqcBXlyH8keHhv5GLcAoPzdot
ukZ48lwYfyivZhcmdF91+/XzB33gJ63XUC0ONEJZnHBdvN5OOgNY/gKIKMLYYI/f
6JiodlY83/Gxd2ZDk/PS67D8Ba2qxrazupZ9VMLg8nhXH/tCd6767ML/aRxiuGAC
H75I4F/f8uDIhdepuuQ9r3LQm50GBA/i+83FRGXrt3nriOCEyPFdrt0zrIa91+m3
zUizB1VF7n47/pDkf1EFzwgpBSwO89xix4a2RazrEX19EycljkZ0PCir8ukvnOl7
eQxX3uf2yq/VXe9hrXGTSDwi5Tz0lBeNZCtHX00WdL0X/6b45Aaoh0RGOzXi63t5
S36QW8silmd2D65bTWZJFAr9SjrutEc0VNlQVih2j7PSVfitJoBdEXyOxh5Y61l9
TkHLYaIaAUC3asHH1aRx3n6AB+jNzhGH6JyM9kowU+c=
`protect END_PROTECTED
