`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gE7FcAfJi3YGCOCyxV8XADnPJuwv3L8CY/Lb06syvj/pRIjcezPdjcqNLVedn8tl
ZqtRmAg4ZcXDxj7CjVxRG0irzXo609qYLijylGJEF4YQi0rJc1p+s7GA+VRv7z6H
vsfFXo4+TCsscX4g9WfViONuVNx9CsQ7Qy0hhG3T2o2jSZnzNoYabGonL8ZoG3WW
8yiYwfHX3mqS8/oKL21RVwUCWr1/b4ULfgZlo/1cPl7dbkVXY3XE+638ox5SZjRq
1EtERepeKX/p50zRLGv2aZq2vYlLikIfNkh0ERaW2yGjwr+gB/HhwHy0MEyaCN49
E4HSiOs3OzeeOJ8AUBpO9cjYdZcGprux0Ir4f1gJJJ6o+Dcs1WowzmQKOGmDtE2k
16KaZ1IxNHLOwY1ZqgpPWA9WHnfLWv3bZP/uum6nUS0Bj+4EIi6WoSmUD6haTzKP
2Q+zCD3RkxFKjIO0FLPNZvzj8tBzIYD66GaRBF4o2Xg7YSuM1ls2ckk8GYRa9xVd
dXAsr8A3KQtubISZAGZUkDandrkLLyx51atmIybnVaYbGcMtC913ECZKIZBkzH8T
M2cLK2+ZA8uhzi0FLL/mJ+0SsTMrICKOuBGKUt1x56tRlZOyTRZc2jK+LrwCgyYo
/qHuzfztkm15TcojyJCCvhxh4MjSwFublGFeisVBprloR6ENiJqpyNJqOWV1UuYY
3K52Lr2peO4PZo9uOdRW5XwCqtHb5QHZ9gua5Lyh7Askv+AjXCJQN0ahLwDUTIrU
05Z4wHjWMT+AhZ1DKILXY/Tesp0g4hsoZRWHyCcx+TALIIO9IezmJ41SqFD68RTJ
0eb0beK6/03E6DvE3kPvpvB12qa+gCbxnEucjpqWNQLav1PXDJo3ItIR/a2CbZXX
0pMbyqHeAbAjUxB3DOearY0bn6y/qjHD09CjqeJuYZ/PSnBIdsFAmRiSmQxiG7s+
NiAwLrZXgnIPyv5lONQKtWbfLsoIzoKXfpEQMLGXtgTRTZsxQmZnj9R/rNyTl17C
`protect END_PROTECTED
