`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUYs6EJRRNy64hRaE70kvyQNtRlKvmK51bZh9Bi5Bb+KWMvqf7n/VtOfiRcw/EC+
wf4aipTn5MlIHv6mmzTFh8bFVjxDo6jtkKE7xOM1x/gQ6DLRdkshI7ftm9d06HKl
UN1+3B6FIFGzKPomgtlCthYfGYO6v7u6+UfjGOYnYncUKZdsQTfBQnYPHIA0OajN
rFOxV194QOTmb++VX7iXlziAP3DumROBuFx5xhUl8RxPurb7yvzfewDBNusgLqIl
6e0C4/CFZDJDANkgRtCONz3VNiBe0ku3nylcWuOiKhRsC986D3gjrDNqXG90vH9h
n4KPDayeawzj6NVymPh7GNWWM18A8a8CeREenYIIT5T31gdP65LEa9dUqtpI0bOw
AfwF/hs3dsz3y3WJan1JQr2qf/elzCrKtNzoUQRwDBo/Yg27ujtxEhW1ngtLVHgI
TrS9gKr8SGHX0kIxFZdDfdCkJDUlR7nHjKFJ1dLvWdTlae5V/JtnbQDgA2fNomnd
CDfwGUmnETbjU1U3ixWqE/KszEOQRBEBEoUWwXBVUs+i1Hd5Bf/5EwuBQFAjECqS
/w7DlrVnjjI/k1hAvAqBsT+2ZvWrVFttSa69LcqUpp7nmjVvGcfNkL5Xq8hSgCYv
n5vsF1qcpnsz8xnh0S0ISryqoNktIPTJh5e/wf8XJrJsVbHeRiC26Mc879DeepFF
jMoaoTTr7RfYl53asXvCLUAhzKe6Y+cBH6TsVbbeC5tKRAD088cNraQvWvdU2LlZ
zGz0gR4tw8xWqsnRS7OiTN1xF0tN5sHN0x+DvwxnNjkpj9cj3cHcXCzX6kWovW23
UB/vLBXaALeG/ceAJmnuE+Sur04pOIcuXGuQ/J1SWKoxsz58pMFRv2j38OMf4tyU
tzLlRjdtFwCASPyw6oynEVAYMzqJ1VxO8kXgufbbgzwsg2El+b83/UQq7HW9euSL
mUwatnwb5IjyVKSU4W8MJSGq57pL/Q8Ta1E2cUaRxR3qJq9nTJ4ImOkBUfsCyHV9
u8dbTVjx58OvXl+rd1FuhKrkWkhL5VBE+ZlrWhsILwX/Ubg7IGap65CTyshbdCC3
od6BAZSUuPvFPPWjY9UvUq/nUXGtjkHZkg5zO0/DiSf/07qd9pc3WPaKwSMMLXFv
l8wd3LRbYv+XrHCeCySSMbTIa7CjMwyRMBpH4LUZza4xwgr0ZJTVHHFA6VMuxunu
23ZkyP7rTr/GvqZ/xPgpCiAEXJiJ3kYcaqzwFwkltog0KmHV/7rSnNp72f29ArdN
qbvRI+eelL8Sx4ntOWo7d6Qx0Ql8mP/4PZtl8wPnmTX6/PyUk0XtoDSIjyZL4nV8
7LbEbdEN2/4gtOtm/jBktfl86raT3NIib8HohWL2wTg8uS99tXQxBT4dJOjEfmGZ
xH/Qkk/JrwWuCxUkLFsyV5k9PoIfS4FbmHvPz9IVwtcDQJyIHiVjAfPj+zDAChdN
5m25m/Qmbo9NCvKlHDOSrGaaweJepQhZ/L8c1fLvApgAhwmtejAwqMDBn1HOxUul
yrMvGMYslRHlrR5Fi+RngPvKOJ3+a2DCChrECtZFRplA1uDrFG+vw+HO+rn2MJ/S
8i0QT3JqGnhbo+9Fy4mOV6jIQvntJH+KTSy3GtrgGLp4uF7iPTiFk3dMDC6r1pGE
bVb0Ii4hFT8jCKKk4HmvWIIjS6JmYuMIqmkDuVW/xr8tNfq5kHVW+ajN943ztad7
no2yxOVLetHEoorlXdWhtNq0SPl+6A2Lu5oGCNaOtu5MVgy0/DUUAxAtwxvJHqUB
KDS0g76w/LBjXmPIRqDfe8dpTV3sTeKq8GDu6N/tNff8D1VDa14wmCrtmTI+k2EY
NjHSYoE2CA3uLg1l7oqRQKWrdzLeotcL2CPhXKRQwVjiCqnZXmBpcQrDafHMdfI+
cutdzBz4j/GBMEbEiAxyCA==
`protect END_PROTECTED
