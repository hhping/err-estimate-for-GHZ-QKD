`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PV9mNhEMSNrZR4q8B08OWLUiyZIom0XacQ97ZIp2I1rMvovp1C+XGogXoBICxufN
oWGJU+jjrgdZGBCTAEObNaNlDmEmyUaxiidoGVC987E4+RxU5aZUhN/AaPv4Tby9
X5FgAaJx/ha7+1J29y/Tup4zY1BU403quf7qEqdWl8EdiOFlfIy9F1kCu8NVhhOP
FLG3M13Qm3oMq5zGD9ZXFE+p3Ebb563nvjlv3TZkrQ0HIEFbL2XxDF7t8Swgn5ic
uUiGpOHHlIAZtPTEgb/PH2LoyGcGXEx7BiIuSLh/OQUYADHXT/NkVnxs1VZDuFLx
iPUxpPM+nYQXG6NvmCV5iCMoblZIZBB/RnYF9Bq6TJfBKKFHYRmhMK+QMEveCgsj
fh5qi0gCGOKkZSRA0NXQbstkLaVpjj/jIHvMb7YZKav1sFNfiGzZteD/fkFTmJZT
UWwxd3q50X5w1TwMn0JO1+swWcFxehwrXMbVfD7ZJa3OKhLaQ0VAmDEFvtzBEvw0
wsmF+0NawAPRNaVBXUrLnhxz+6cJ7/kGfzF/n+zVP4XgrZnZPQOorN0gnpoW55Zt
LaLkq/rjgKul3UHQQxMGLQ+kyPpiaVkCt/xPYRDN+dspgUvkJBY8d+T/AYS0iazr
ywu4d0TTS/AotK/0sdu4oFKmY2B66dXI6smWzYT+uprCMR46UI4PPkkHxFEE0fYe
SVrDNGtdXrkfgyUY2qPK+SvCSkA8Pnw1WESzp7Mxrxxv1pMq1B0QEEE7aLARqgO2
VZ239CSmsPUVg2+3aHI8MEHfnCj155Kp0PId2iEf2Q/YWpAEodUBaLG7Lbn7aBOp
p8EtzPai+dplqSQ2d2NMq/FtFG3pEZQG3EcJD1uHJ4jS5ZFDPNPull2uoaQYNwc9
Av7CRNmHaaiJbLQoTIhaO5hKDXtrCP9qgPIJiHQQkiUfX8gvikC2NbpGqcczduzW
5jbfrrKxGM4Iu82J7h9cZWCGUnnPesFS9M82VoEf9qFNvTsdFT81htTxawdcDtdM
P7aKMZYZ2thMpxgh6JLqkAnf2JhFAMQnMvagx7/Q1MQ=
`protect END_PROTECTED
