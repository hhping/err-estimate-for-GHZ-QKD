`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sgq+V21UulkA0F11pntASL1AuyVMOEiBT0XegIo0nF6mwqGPzAK7MrFh58D4BaKo
HaVEsmaZsAGwl6Ers7CByvV/o+no722+ig0ypLVA5B5rqKapziVMqJvzhnZnIeMo
Tu/lHsmq8+bDdSm+o1tIT5F5yEWZb6Afr8QeQJViDtFCE/cG522Nl4Oydo1+zWZq
GEjiWZrYbcNVdvwcaIuwVFxL4f1gCE3xI2T3YsXLtsKTs/cgQaEjs/05ZiSkD1gf
jNyslh0C2xWp7NVDWAIPtRXq4PGxrgRtz6caxYTCdMpbA3TPX620ocyRLlch49Pu
csvY8ymAzlm0+TnSz9lKio52IQ6RC79oB4X0i2AxDuYQdGBPyMErvt0HqvEtRw5M
EPXnUe3PkHKzpA5PPAekav444u+eRbSerjNWLf4BHd0rvhQbuSRs+aGBpAFvFuXI
wvl/x07jhRW8+XzPHWVPrg6q80JmS3SkoAr9m1jpHbrBlyF8jTRsgMp5F3M0URDQ
itfHsgpFON7bGRK9lkhv+ho7/5Sqj+QPrgBzHGJugsXLo+FQMaY3Hb/TvjrpI6MP
LE/ytGfcd2KPOM/w7PO3W1DNjKKh/yYdwvQEIpn6rEzFZ3O9PFF6DfdCrFs7wt+7
O52MbJjm2M3skw/qo5AeIDU5Fhj8kMpQ8MIwyjFo0+yyDxvZObi8iMKMuyroVVii
YcQg35Eg//ejAyxHvKEOD50xSPH194EF5A/XP9l5H/Tn9L/XZY1ETKyP/uQzrEJJ
q/ZqW6aceKxq9TXhaTGd6MtujXcWxT/OBZl4H+fYrWe7Z6B1l9SG2G5s+NWo+KUJ
Y8NFz2kIcQmtg5dhujEXkaSG7eRRl74d8tn9AxVJHmmM0RqtXhdVjWX+hWTGxU2s
AXtRGC+2chmf922wcKpG6o/1VeGUYUH+TGyF5XhB8P3bP2cqTZgWr8RGpTW3Z6aP
jh2JJosYfq62S+EzMYNLlAZZ/6Mf/e+qjRqKCpDcK67f2A72J/ceB94H3DdOn1Q3
JUiSJnBKHO630wJQYdNOcluXSboPOIl9B9us0G9yjJlcavLeyNIcco0/9iZEEjPn
3ztMhJfbXgV6LgqHJ0o/1jNNXnuWWpNuhiaYa3zAkWO57m72/s3jh6r9M1Bey3Nq
TbaStoT6OS5suZW5Ed6PJGBZTWPxJZNDHaxf0E9F4rmqtqBPOS3S6FqVKQWxK5qi
NnGfdCQjcfDmU19eSNLG16A4nQ7xLxhpzG5puhnkCmflTwYAmBIRGW7woMBGVTX1
Lg5t1v/n4+x4tyXlsp0i+w==
`protect END_PROTECTED
