`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qkAp5StOux3D+QGiwjkye7i6AUEPJ0NSPzdEua3t4uuAtCjw/o1Ddw0PVUUJ1Lsp
B9iOY2bz9AAlj5uE9yYO+Z8GCBe3/R6ce5RvKd9AjNh58RdQgSuzA8x1DGjNj2AL
D7CfLZovmweuD9to1Ob5mInJP/28C0APbgFUh9rf7BnPNcwMWmky9ZqpDTt6mMtk
HqJxaXFPZGnP8nH3jOe/iJVD5mr+7tKN49eLkVDukwSBgupxqnK5NLQVY0tcGCuU
QDUffbbLhJOMqFS87XutI/uoVfvvBc76A0W4hEb9YQei1Kx/C7XjB5BvkL16PZLk
o2799Hd7UZ5kbpKwPvGO/ZbmP20AN8D+wVaMNuhPT4t8OawfQVzsnLkQpCJW31mJ
l7QGksO3dbh4ylgGVGFoTi3h8BF7jNRHimuCQ0hFoVgBuMOyf0Hhh6zJd7nwed6c
RFYzZKbR5rFGF7SIPrr++xKZvUkJMSVyhhgrWZ8gLzOPDy3EekjXzqBI5sSBKr25
aZQymvhD1S+YJ5H0Wsg27vRzYNi4chmLYBiNgasUTOajEtE+U4hbHLgIyOVxyiTB
9FGVt30jg8dFG9UUu1OsP46UnMFkygxlPzjUDBCSsFaAsiemh0E3UXxTpECqP9tT
SeNHn85MYpMRN51pCJgKUfH/5iVNKWOvocwa3wWdyi+KqtFij1OfgAiY97dJ2o57
4btdoEIndfkTUUWM52MFGuuRlO4OzOef3vMwpU10zlPRv9CdvZjOGHKXZVya8BWt
4wKffhHXghtNV8YTC/tuU9USvE0FccE2zJTfESyYKyt1bo0eWiJzBFuN9jDzLE8Z
0jljQGkJoUzjxXON15oKPUzx9/paWqu2pXm8+7cFBPV1EI6hFZdoOsjTIagvkDMC
2xQDoR2Zi+aZErsdf4IwxQ3yauHnRioaPnnRwaW6iVKmr1+itaDKqspm32mmyDl6
re31ZvM+eXpDtpwqMXpZ94dRHMjlTDomQuhzuXbQKs0/NFhmWmC64+VoXcuiJmrS
HB7TPR1uSb+aXryQ0ayVq6Q6+2R8jFPfPuj3J6ui/n8=
`protect END_PROTECTED
