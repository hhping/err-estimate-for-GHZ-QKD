`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tk1G5uo+CXL8EfGd4+98mXywKYA24u9ng4MvXBXyjhXLW5GEJEqXKB3vCNQjz/yV
JY8DRhryMoYZcZdtl/uW+effWu/oRDzeEGBf+MKZpz+zC+n3uTA3eoCH8Twy0UQS
AvIHBE31czwC6xe0w229LQGxM53+arYqLDBmWqw/6QW6S6UUgbo4QtOknrhurTKl
p5sgWP+6iHVUU12YcbSABC8JR6G71OpN6iFzqe4R3S88OxERfcGFHE8UIFyIDT6z
b2U/BGgdJgbC/v5kWsthhw21B4xfMv3Gh8DQoG2KvhNrXWxSX5XCtNBjKS5BveNq
zNYcrlZCpw3TwC7wwxCzsVQJ5SvlPxT4pD+9k+j5tuQWXwxgV/jVp6tOLXqgDKtN
i+t5tgQrmVWDX3Erbxntn+1CXmZfMLcakcWR2tvaCLcdMGdW1v75p8g3VVla8nVc
snT1sYblQtul3p7cfPP0lvDgLsgFUfY+lVjEYoEeOlB27GY39iQ53y+OUJrtWovo
R3qVZXrrZA4cyRCqAF+7/xeXuNQTPCO7ppMU0urFxSIB9YM/WZu4JGjrmLC0erDA
bdJfZCxnwaaQRu646py+qeKQnmVxjJuscFtw67oSy1l4sN9SKHV1Qmhirmy45q9S
qWjIz17qTAyKRRadT1HFQjCNaws73TQDFnCM9CgVTgQYP9Obq281xCnvJ54gD0Nq
+KxggBnsSVWTufx0Q4Sfa1XpKSFm3RCxrSC3NXDYL3ryCZFJODgEAeAuhYIDil+z
XR5qEhUCcS3RjKStFggJR5odOLtlJZ+CigYPiFLI2E0WCs48fw5YhoI5IW3OvQnE
`protect END_PROTECTED
