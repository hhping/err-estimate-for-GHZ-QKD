`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tIIugQsD64hJA71nNoRju4R9LJVTku/onC7GQ1Bl5C6Rkor/kJkoBoSNQmO6FysZ
i0FzrH7aeLUVNLGe0zMT1JUbqkwDxJRSuse+a6va581B8RcJY3suUqfURDcppzFh
516n632ri3Asr7imv5WnNvXW6CZc4rdI+m7tlJzaUGg2oPKhAaiAf8xq24OHr3H/
ATVNPO2iIXRh5xRJmj/wlxlzl0sQ0KbnnNALkg2ikzAkrYqUFw98k4uVgnywDiCS
GLhgKgEXWdqdk/MNqlVT98YtP+1T7lx/797daC3bgZyyAdSK5WnFTjY3jo3f5kYF
lmnZ5GnwYF9g7dB1E21NoKu8ZjlkQ8gAVCHTRBbvRJ0HrkKg+8v6RxxBpiYDnQQ2
1YL74bXuTEPTvwkPqyAWcQbe82aTrt6+WZ7dJ3A6cNHk6i80zGAaU5GNnv3VkXy/
mB3MENTsyJwiEO9BmUVgpQom7euBwU8ImKZBRVd1ILAME/0G7eVq5IRndQ96rsjN
0myJycGhX4pbhrK1bWl8f1gJ+shyJdoDXfKfSIhp4qPiMxR4+iSuWxfbIRCS4ANQ
wUg4LHDM+oUAu5o/TUFu7v7itf1ghzAVwHTzIq1/W6KZP+sriS0mxlgG2aBBotHH
5D1Rqd1D3FYFY6TiHm46+rsqVN0Oh847nLglTiTv5Lzmmxj+/ONTb+gWqcqh09Q/
iXp1YUNnzf76jUBhBWNMMY+LkmtBL+TKRYG7dhZ8RRD5A03HmD/CmkZvOTPvW/iE
0jpRn+doPd1jCiGAg5LRIwX3LtgnyG/W4jVxaWMtZBuSuuRtzwsokzWXXk2F3FVL
g2Gds7ObnJPc7S5Pd5O1oGd1xek731sXKraI4qv3dthECqSak2uOUz0RPwaz34lc
ZSifw7bQAdzBpIJPz+TfV8xGwxQ/uEBjRt3m6yAwPAxnPaRYiUfAx4rTJBJKkBUV
H0icun+K0DTO4t92pRUtXc0/PpNARQ7Xpq4ex4zhcEFzHyujvFiabts9zydSV+HP
yTw8ONeQB1lJExie8GPaaPBCKmfr3OnGYI0yg1KvFJgnqlA6FY/RL9z7tBLVGZDf
+3kDlqpR2JsmWJhKt3obLeJBg8pM0zrXNcgW816ocutxEW48QBipK7z+uOXQDBzt
45UU2uXD9ho9/1gfv9wQDy//Qqv26Zr1Ln+kpOE8J0zC56zER0gkxAaJxYbQvooy
dLKggose3rUVgWOqYn/ev5W/Beh4dh656purDrR4TMYnLWABqDj4eOhEddtTLGgR
/iWSEeFFf0oAiCw6q2GJbr5VseaaC9dm6G/K5LV46ilc2FgeAcepCwWFRhhkb5b5
a2jPO5myGO6vCfypOtBua4z9KThCiAUR/FfK3OP4xvM3KxGU/lfOac7vKMSa1xW5
jt+KGkEdE3alpxY8yoaAslm2F0/OQART2jT4e/0SEet/4ABjy8Z19UlubqywbURd
98TfV7BX3dZ84aV3c7ovLuwRgDn909cAv5kYyd9gzHrQ837dtrYuT4zcLUe1Xr1Z
PpC5pvR7XyinlGFhiyyxI5yRBGi0DSx3zeIB5cy3jr0eEVdeig0pFsgScSP4FjPd
VImIkDOlKQuWSdcbhliZLa5EyziNFfrWUbkUMAfE4SWnixY67OV/oYVUz4oI5Dx3
udeVlkwyQbKrP8Dv0G52Pg6VMJ5ZM+8ElVO/T4+bJAKMnPXoYflCB/4+U9I0FHGU
2zWELcl3n7pkhMUdx75FeN4T7iEdcRycQNdZ3oIoTSQd599RK+JdHysIybkcnApW
g4fSVSyClpT2QL/s2jMaPRTfOAl7jvm982HMXknffWaDYbgIOsLjiWlidZ5imB/1
e2jZdWa56yjGLRPEL4O/qUu+pt0VTptQDh0immdZaxrFfMMrcqKqlDLMpl3eRsS2
gTaLqj3IDNcj5R3u1PJ4ygM215VhiDhiMKHn1C69Pg8MnSJD/X2EYZaSlW6Xr2k0
thHQuAY9Y0Ud1vrJC42eMp3dASoEWZCjWZuJNgGvaquAsgmlsbd/X52f84gpqg1S
S5h8BUmuPJRgVM07u2DU2om5PUmPsf/fzXN+hKmlWWOurn1n6YXwJQcdFzq4KaIX
KHvL7ZOFjQkTM9Mxfcb04mpYaFMGK8CJUjC4xVQSvjAzRbDU8ajGxZmjmcQx6ueH
J4G7EH79aw+oDnvMTtPXsZa2bVWcGf8ULH0IVqx4fW4XrvalcbCpUso/w45CMjdx
I2Td8AK00a9B1CE3DpMAtvjK2jgpKTVsTfR+tELg3g469IQ9QoBayP8BA1p+uxn6
`protect END_PROTECTED
