`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pltcsZLRqvBso5rXi8N1l2+XZDICk+hkEMArEMvBNpIUlZQnqbUdj9/nzIWdej6
rnJ6LqAOg2eIPQXRdUYNSJzSj1OQzxo6WhyXyp43M0Eba6AllixyWS//85OIRvnb
w2MvWGzjAsUFCgmxgEhxwlLYHu9/1Dh6ifZ4tdlbu13zmEKwj6Xk82pJ4+bggxpW
CrIKCFyG+t9pq3A/MHO2d2HVB86R2KDy1bPQ2C3yg/wE0hRaFROIbrKqWpBj8Pge
wOmzszXRWcWv96uQKK1cAUlUnHAdXjhbgmH8LmhOjSCntG44EnRpMxIpEmen64x/
+47zK/pONr2kg+kYGeh7n70ZLtEJae82TyO/XTdUBmUdxl7xKm7QyArWf1RB5v7w
0IsLFgWaLks5cDFQzihkl3/MWgQ9E4a6aWviVSKnnPnaUggJ6wTY04Qd1ek/17kQ
118tUOB4YJ25E3oH4KYYBlZbCVvTuroi3Kx8pfVWzMjAEzoB5wVSyf0ZZTxT5+Lj
LdtTcN8JGDEfpmICe2w2ucarBPFOPYghMVnVBg5RUp4jJ5yOA1B/BhvOdtffq65c
0ACnG8E1IA+18Ea7P5QKbDhhZx77AVPRuV8JUTUTR7wqQXuTmY0F543K8CPsOx7m
Q7sQaHF6sCCnV7ax3iCgwYIeVfoyvJEBoHlkUDV/E8ywyczHwJQLHjG90a3NAvbP
HaS+2oqLHwPBoZrDGPAA/HsTECxP6v4JjV4o8Tz0t5o=
`protect END_PROTECTED
