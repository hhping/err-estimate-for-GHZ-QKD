`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCUTCUUvrX3QtDS+sAmPxUkyACSHzA0BhmQXqyLWsyzWFdyxWLrfEVVcD0IXbx3n
IA4OP5QzsDVMgRMlox5Sz8dFxm1/szKZncxPwxm4l1Wsty+rGCR8qcUucvdIeFlK
05dnxsepwDbTbth6XGJ8968y93VwrY6jWzO1ehyXZyy5wj46U2d0BLZn6BP11dOy
L6VQRQxrfjQTdkZ7OlfMxmX7LSithH6V3CVIHmOU/O/BBNUGyFv9cfJLSflmVQi3
PnQBeNj4ZTHGTMugVf/OEkitTskmMk0WO6Fhd3/OF0dfNEORUHEwdESPL55OUJDg
saMAEkpHTL9/G5dXETXETFq7RpaYo9/sPUzpvkGxJ5m+vzw1XF3ThjiEF5iXYRB2
nyLV6/NMFSxyW4KH6RfIU6ihgV5OGycOh5wKZmLzz9e/Milp/4Vay6biyLGuv3FO
dJzXhi1WcQvhZbyVs40ctBj2iBTBbzKGuThfcnDXuCf6VM1oIAWaqILCbuOMb1+v
1hLL7Xq9zNfBlsLN0akvKm186Ka92ybuMKIMowTdiQLAPaJ54i7IJE5tPLZgr1dz
fFFBy0NdbvFg8NlyRumPm69DnxG/FUsMO9fao6F8smbYXUTSsQyrHzKsRoLN5l7l
TbJzsKDendALHDf9vsSvrDobPy0VKZlGSNWcD0BgQwukTRlIyQKnaT/W9FAbZx80
e/Z4NU7T7Nrh42bL0dOSBvSbXSJ7XUhHjuAljyL9gvmx0vHNTFLTf8P/CNC/uQLJ
of6j621cDFS+fBgZNp7odt/m82KyCNp4gaNmvB0MRqie2uCY+lGv6sCiS6tGapmQ
wPQIuLjJDSAXpMlTgF7c6NDpq7qEeFHJZD+2avWhKB00kc4ZwrvWQt0psOnU7e/M
zrxb5lyySRmeEzAuwyi0UC1JYSrUwkkcRKuJ3BexSNcyMon8pYkD7vTbx4L5TzTM
+SPBJs+IPG5rPbjPXlXmQxxr4WZRJBGu9nPpdzb8TkZvi9sI+ulxeZIfb0S7CClI
SjaAg8DV5ZW2oBd0TgojoC1YZ7WMIQLdlNF4vZrzTJEDSRLi/8vG9yWSEQAmSGhK
WnQIO0YZK8K0cm94IGThangVjG7w6T+nodrQX07Apt9ct9VhM2ns5ERH1NnLD3k6
EiLImnV3iXJtpx0Y5UqnvO2uS1e7QwYNaSialNPWC/XrOD5Spl8o0sRsm0kvwORu
2ZmkS8rfdwe5WVVJ1/6yDvUMqEurcC813w6X+grAqztytW/yQnQc+xTopgRzXt5N
cFeF5Zhe003sRa3sRhYy2LmilTcE5B1F70YDu/odMpSbJY9+JMOcU9RuH8NcLGpt
WRt2Y0y7OABw4GtHx2Pcj4lqgbCVmDrIeJcCb0U/+eT3IRxYaFUJmVFhJA7ZdLbr
SW7rCgh0Fh2Fu6WXKCz2okQz3u8EtgVX3DnBchauFqR8dYViqrMHzHk7OUV/TS2S
TcDXdzk/F0z1QQsranyH5zFmAElKEKu449fUVlUs4SJl/3I7oIFE5o8sT41RQeqD
8rBheqpXvTXXsT4xhQ7k2Ak2fbsipkFu3pjvQI0TleytH+wUN64bPT/GOmwAienZ
a6DGv4c26Xj+40Xx0ud0oT6eIOwS1feDBYuP8upp2/Osu/D/303LQMhzMVqKLCOG
MTTYcfwV7t5mRxkkknaEuiaN3EWsbZGtsJGrBn/z/wABI6nXUqrDoe1rbrogrNTl
15D//IK6zrfhXQ/9ghzZy8/+ffTzTjEK+1NeLRJFNV5hy8hh1ZZbSZmJ52HWvpan
5qgbUvhz506cFLPsKIk4GUJ6XnF/xbWK2WZvwA01aSh05S2jWecQD3f0uCaBrcvj
vB3Lll4uphEo7uCQBWFYtan3Jtvn9S62jO7nunvF0vKXlOpB6y7/bLSNP1Pt3RT7
QWYbbB6a5TPdwogE1TfiL77mvSagzqtu6PjnRA0MN6zK/kKmVgP1l2x+mN4mAe9f
D3yhAUrDC5h9CZQodKRVfdCGoWGfLtBiKvjI59p/vzAziMoTKwtDCWUzoUsQ93qH
lzUxwrxh7+iWFRhnzvV2/r6+04y8Oa6kc2dBYhxPKiUhaKqFqh82GR8ZFtWJ4yJU
lzIOlLhgN8XCaKIZalZTrPXbug0wnlbinfcAUt+JHpXHUGd5K/PX07a3RTElH3La
SMyNHyhI7iEGEaDKIJykDWw4HjM5/EgZ2+2SkyVt6fEUpEIxBrLo740Er3yXtMl7
n6G+1dh148htUaHQHGPavfWl5aNl3JV9RrLtePb8NjkYWG43pkTv0P6Ct2Sux7PJ
38Pa/syXP86h6EL/imF9I9Ymh0symdiyskOBx4SULSGJ6UlwOML9CV7LQ+y4ijpt
ksuDAEc52Hwi3CVB1wwBSa0aih00m5s0W7oVUxKDhlyF+JNKkyKIq/UQrfGoV4al
fsDVvouzOgRWA3E3T/LIWtnhTrEaebDS66nv+AwVbdBi5Jxz/pvQGJlZG4/OQW5l
Iry4WjhkAGwzIODVTi9wzDaqBLTmAC8cYH5d98AAX/81+yPw3Ei3QhJ6N1sPRtaz
B8XDWXth4Hto/h4Bx8oxoQYvqFY3zTCI5bUhkLAzOC22Amps7jYXhCCt08Sj02qM
8cixe9W7AzzpXjD+Brv6d+SIPqFFZiY23V4oLPAYtEdETg2jrzd2IddympwnbNXb
d1Tu97R6DfhKoezEd8Wmo1KMh+51A9tZoR16zZ8vTBRhl13Yb9i/fIWjbR13z5VL
NzyD56iIPulf25bf+8dgKfjj+MB9zmay/b4ASNF3ghTJ/GgbIkcG7zghbv3JnNwz
4f211Ylojkt8AJgpXj9xij1xdTyRmp9KvWsobNC4t79CY7SlhvWxmkQrbeFPqA+B
UaLeOx4NWGIahFp1T4cs5yigFAjM0DfAnlE7wsZjGsCMr7sSHEAQuuBjnvz1zCPD
omVNJFXe4Z3qwDPLDhfuDDIPd2KjjzKRDbN3JC3Deb9BfkuBTZWTDbXf/sdb79wt
GZe3OrBydTvcSQyUY6VawDQI8pLPCdTCkba6tlZYDpWKyZ9cqQUIv38McaQ2Htse
m5Dzqq7Hwmrq9wMyDbXycjIoS72v41KJc33OzkYyP7YmrD6trAVFhRgu+kt04QbH
NLQkkFXjOX1+7qLaHs2rqAR1pk2zI6EKwkz8uFVeLwn5B9tm9mWM1btDqpzhRWkR
Qeqt77LTYgwsoR9aVmxdNKJx/ZjDPnUBspr15sq+i/wEPpTv8Vq3tKXnT+1VTDdN
0PGB3jr/WzSX71wUh0M6kQl2Ck94guEiClf2cKHv6rHW99YQIwIIqOayhSXJpiEN
vJPLlDNf7o/qyjrOVr3/of58Js5Bd+JY3TBAkWI/ZViKilp2nHEn80skv2fJy+B5
HEP/9BLFJfZM4tMwrRf85lS1WB0HEbBARgOa0SI62hS/L9YLtJYzh1d8Q7BGdHUS
xALF99c3PL8XLiJnWNX4HoCTmdn3EvUtqqjX5tNNAaFJxpc+hKbOY8cxhO+VzoPn
nqFn3xhNf0pJ6zHkpliTLxS91sKiiY24jgreDd8zXiKTaJPzHMHyWJ7wuXOJ3eCj
EMhSfJeeqzJNPZasK8tshcstzHt8FXSY3FcU8DXEUWn+Mg1b8gQPBbN1SUofBPpM
NnfbceiExSNoQh2VFuMNhzYUFji6Sq6IquIeOMvLzHKY/sF8Mb+dEue29BpGRU0f
eJH4R+Odsc4UJVIO1oYjwfy2mWvBmSWLmKcYTmngfONE1weH8uROhY7kMGzapq1B
fk01bCUNVvuWgwlQRKBoOJB6cwIjclz9RULNL0rIsQTOhJMcBosw4+2jQLj1WKWA
wSj1ejuXpKNKaduUS7lHe43EfVDcRxgB9dlPFE0s21QLuzDr5MEkcBHGgxSyayAR
ZAGczZh6KY8EgifdqAIRKXfol1jwuZ2OT6e4NySiF4MSBz5tPv/K6R2FBd0P5Jk3
78xSAED8iVyKpWitDzKu7OxYyk2bNoHnveqyToz+cDY4bGxuD93R5n9LgemS0uJC
mvHnBcMxytBBNen4RtQuffnVllDe+XgGgSCYCY1j5otlYhUEUGKTiTCr4OMvB+La
P9J1DozuAmgE0LZ4tbUVLsbKP0YJxID44cY1DPMx07hUJwMCkoTB7Gi7gyJM7h/J
E4NXQzsWwScNTMQyjawveXY6NLy+6qQ2I6rxZ1rmekS5087mNvV81AsNOGcc0ADJ
djtECKc4fW/OPrJYlkfF8BKaj8wp6wpkQiEOv9hgrMvjpSbIfcT+Bi5p5CSwrvHR
9FeWQU9uG8P2i1eZxz8DKO48ufnJ1lsvtDFtDNkt/uh+PEDeHt7WLYoVixtZ22X8
/S1SCT+39Ug/ldrOzMhoRnIksALIt2QLSZ9O/2t4YIpdHZ7nuZbiR+qa8ctRc/JZ
riDwxOUF8yeZtEiW7wvr0Dkwx8q9MjilAp3h/NpKbYADol6QAQoVk6TB+GwemOft
K7IJCjPk351NxmgBk7wJ1BQSa91/c+5KMI0QbL/poHQPVJWnLFrhyEuF/YpBT+px
g1AONrw/Z1SpX5xrigv0KBIzKj+WsngcEhaF5cmwA9cLkMTntulPhaA1Llt4jsLK
xGI3lHNlMiid4V7KJBPG/wJMaKcvuN5Dpj72Ik/YhCzPVZcF/jyC7OH5LkhVVrYf
MXI0Aqe/ChjZwQPxiFQpmS4abHwzbuoosd6IwHtJExLBr1WM4pgxWoxLS7gAtdfu
u8ibdsvFmFySlBi2ewbPsH2zGBVrLN5PUZDc84KpZC9HoUAtPI16E3yDDtTN54Sp
m+CzEr/QXVsXTY+tTuENM2WhgwSw5Lgyak1UbhyRVdNCktlOPqiatpVe8W6opWRk
uWOoyBMZ3xOgHlTDowIz6Yvd9ZQrBrndkvrLLOv5zpdXuN2aX3gu70itwxP41TbV
ALwYUNQIxF5UkV4jZ6A1tN9vYH7zDIAHC6QWmgH9L5HzHBc7YvcvZMHzhF4abJSq
xF58CjQNqjhZxRelzzah+KKXCYJ3cTDlKZKDgiS+C5SvaPInEt0w4ffMmGTJy0ED
6TGSQD1hruZueAp2moJKiKEMdRdDX1NKSJBC4lrSgGyiok669K+1T1WzQPOQyNko
Ep6fJtWv6gSbNToWiv/zSk9/QGuMHWeBr5ynE5y+N/sTvCEYc3o9rFIAmV9ymNuN
8zCtir0qpHshI3T8lpt4XCffXjSmQRqjXBgQASvBNrIW5xmn3IhmttYubbQFNwAv
Lp8tyWA0i4CK6O0IxOYaiY4q0rdeHF31cb7sNMKhazC3cytgNiFMN7/tXBtfj0hf
o13OZ8f9hqvioKYnKgbbDBjwixvjbqU0fCD6fHioKKE52SpHfAl33u+HfdDPtFnU
Z9BkmqalUSNRAHpYORkbMlro4WO1YzxwgPuM8Rc8oGBJXhcDr5lw1ibA2tA0kM8j
fFpW6NGE3Mm4b4pJ3sjNTOfJTz+JzdaDgHzjCXvE+cs=
`protect END_PROTECTED
