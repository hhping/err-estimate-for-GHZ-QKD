`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2e6+1/NAU2VSKckTkZ2xhtTOppH3GAFP+uy6cWVq8cwI4Zv2OWo9VO7Hh+V7H6vt
/tru1+KWZl854d58JDzWqysHThjnzaV60XLhnfyc4D23WfQhCmET+Ygk+I0Rfo8Y
rctSDyIXNJ33inhEeZ62JLa92iTbm3MBLhx5wSeo2wIsWEv+W86qGymFiwGB1bcA
kBTT+gr98HnXPdR0797GGL4P/gO3VpEuLLBDEhyFgfZIWTiPEmcamapVFA2TbWk9
CIBdFilcpL1767eo0MUbYh5yZlqf7i9/yY2pqYQsHbYhZWNBw8str70diqDgR3PU
ccMD/FCOEFFHGICDcpWE5a6oDWJKVssYd4iuyZH4mqze7TjFmu8QuVO4EOQawBEP
rrhWXGymGeImDToYLcohHpmfVvZ8anphw6vwvInHBYcB0oXSM+jrpKmjJrmf5lOb
R86+W9RA7nO+OIBsLsYQK5bKJ1Jatkh3ENCBGzBI8s+ZbwOjJImsSs1lrV9WIEUP
YrJaGH26w1h74ggp/QppAzUXXJ97t3Lj1FJLC+aGicpppauR58wnnJIX4MYY1v/F
QlSBmabS9MArB8WZN7a3Y5jFvGsEbGHqWz794Q6GSv9MkblPClS8UJAiUWcS2JeX
/vOgXXAG4M2yV+QjkOlJmKZUAH/51Z8UVfdbq93tv+5bRX7xGJLLbTkj+AT2Pok3
XokJU2aSNXQmrjQ42+Mro6Qx13vzjV9EYim5L7SgTWM+UO4h7+pd0wiABd5qSKZ4
/N61BpDj9yKIcZvlscPkJbP0XtCkUMycIceHKKy0o40irkD7mjhE/mh01VrWFaKT
jT1XKukUszOKYOdtAehwABNx5ZdBNWVo10WKyVjcmPOVKJyDd8w3eqEbJ8GiKdYE
ACz2ZyOha2Vff+em7h5a2OkTaZbiqYaFMI+MDELLTU010YZQtLjYsJs1te90e7mA
G8cnZW7HUkA+2zacLSHhO4aRkBCBtobX9YDDI880rFQTfEuH4V8KOYAp62CkxEAm
lsHh78YrnfBNIKG7VymsoM/r0UkhFCk3LYKahGeRbP8Ad9RWCe22DhW2EmBM8E+r
bTKKDuuiqbHpzY/TQKP6p2V9zYENAoLbtG9wdJvcJxJqO3vhl0In9MhPfNUnQcV4
XJF22iu9Wpjs7i1mc4yuoNzoG0zvJaeSpC7WVtMoUsLKOckAu0zNrYrmnAqVhIqB
xSVf/pripmxPCfxnMTzjOVhGK7HooK+rmLGz2cWr00VJZC24nx6+xI+CZw8aASeZ
ZlqWUZWRM9Nwd4zhtlLyR8jlA3ekEKHqLoe1P75H9grc9DveNh+QO+Z3rSKsTIGs
U0DDQ8cyMcYtk6tE+vWIIPJ1IxtMvENt/eX1JULDdoOGrAmHugt2KBtzwxihM/OC
x/znJ9xMKnJLl3uZmbMDL4fVqD9LBKAfweufnorRrax7SGL53dTD4DUFvfvRb0Jk
ezDhONFXGXEuUZ8wVl0wkjQeIsdBix34IR3JajkNYkKJfMFQ0COiA7enoeppZAZm
8zoJKPhmdlH7kqRxrLDanmDC6LDoZWBKzm3yMSFUTcfDuNpTP++43wLES2FC8+Pw
Jv9vaMrNnyPPmp85GW78S/Fj2z7kj+5CP8iIqP9hJTGJcu6QLaPwr12F70fBznnL
JKBUPTvFRQ0vNy1Q+PqqFgKDR5VWeNjSE2ELua958X4=
`protect END_PROTECTED
