`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yv9v/IAP2jI4HWET3eyD4agLOyksi/63CuDVxso6HSWyqSHYjSAczXEfkwHe/Hbo
kDt/wndxXvSz9nB4eKP2KloeUn5dbXYVNfiLvVDJfRtcq+W7oQZ5k3TmrInA5kY1
xlgWLO9JoaF9+C/ike/9VI40tWdvoxs+ezCm852SOdV3GEmF8j6/1uxCbyC99g0V
Nt+p8H6vGT8Aeudh7QY3SerYBnLSOkt1aygIQgCixjC9Ao2X/GMHhtIhcJTgaVrk
YL54KvudnK9c40exorNi4WGIYd2BymNQz6LWNmdPuBNmwmH6wbAUOJU260vD2JMf
9tXUpqp2KJONosWYUXDtcTC3Y05BpydT3DctJPJ0ysaQzPqhnxVo57tu9YSqz6Rg
/azFYbB5Ilmp5zh6iHlXVjg2y85WeK9yB8vNuFfBstuxFF622++kAzvb9tUaT/jY
MdtfDxzkdR9p4wdLwW5o/hKBzvSY3ipsredAz6bZu0dbntlmd02f/P3bk2wJsV2f
7wxinqOXQ1MyKZ8rsJVXJMreAWm0ZXkQUmRoPIQl7ETcAMtLiozzMp/8gVuq410X
NSMtyaBnMDHi8X9sXKHd6Z1hU2znmE1IviRIAhKvYMwQVrS1bZh97uhLArlWovyH
`protect END_PROTECTED
