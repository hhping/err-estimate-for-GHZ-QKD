`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vG+9q3En+iWLb5xCXT9FEmqBkUZeEEaq8dAYUkDaAzYW3MYFO0rtN5L8w7+rauO7
sOTA/Q8LtRt4FMb9KLyM8VOa65wdeZEw5Yg3oyHwfKv086ivHR71UUYwJ2wsBME4
OH1OTW2/BkdEnNXnq4mNilb2JrsDslu1WFRQlF4ssAMRw9dYbeBns7AVmxRJ/A3o
PkD2uhGmsg9X8nS6nY3JG38FN2BZtD5zPodVMdzoX/yMiqaFbmoaFfxwusPsYkOr
1INMCHL3xcGvcGZBpkZPq30nAuv/fqV8KIuqYv6/FQBCHp57D7p4Z8O+BzA8jOzU
qjXdnOm+Ie5nOL/F/n8zuRt9WgMnkwBLh/lZSULv0uJ8d/6Z7iPSiuAuJc1ZhNpu
F4B/mDdHRe61jTs04u3eov7oS6zNxnAQ6pSneQ3AreqMnIjoqFvPLQZ/oO5IS140
/kGFZHU60Vyq/IwA8ortPj/pmA2ufkGTRkwdHwkBO2bJI0kkodX7e9d/0goOx9VY
zLSbPzDSs/PxenaN4aR2MCxU6uIik5YrLFyBvFsBKkZhtSaX00H1B0eTjXDcSxH6
hKD57JwD+ZInuEO0bPyDxVRi3zIfdxhF+SRYvUW7jwqzI+ZgAykG0wEq4TLLXbTo
BOgj2r1SUEk2V8H7anlsE91csyIPE4huZXznmVssguXDX1VGcQY0UZMj8kj9EyeG
w/KECp60e33o4+2bmE4K0II7r1rOFAwmmj3OGawS0DJA8pmSHLxY8OxpDXgdlQxU
6nU3Ev3NaDF4dmeimaRn1TXGZu2jY4KcAOVgOIA59joQrpclHp3CV6mf0A77XpLZ
XgDsMoCzxxAfBi3xIkz8UXvsKxwWs+aBUWYhiUcDOF1RlD7PJh+YXVS9UEsnkMkF
ESiRoRkBaeWA0wIhATjLVUh01TD5/0uYgGpzhw6Ns4twsmfr+YDMS5hCahsAd1va
dG6/+t76enTwF9TyCHzkMa4RanOaZ6efX7AnCa/Xsj//AF2KC7EAPCwETXjKoDrp
4hMsQkVK+ayjqd8zrBxtMUTCWe+3zQE44rVEAxNfTWoEW1Bko9QLFcxZFJPe7KYP
qN+UVO76t206oOM4v/WbRDiqy5Z/p1pvXEOgdLveYL4K3yVbq3PLryqUhU8OCqlF
a18T/N2/CIuzmr3506P933UtmEXxICDOwXJaJSagJyAJfZM4T6YiIN2Z5YvvbcHT
hN5yffr/rUMGMt484/2/1SZoEVeDoNOXTBG8j00TLVn9Wqd57MXJpxgOY1yVBqUx
WyUaruDXkdz4Txu6OxisNglYG9tJO+NPsZasXkpOV6G+DgyjF3t1/S0z5pPVhN8g
nysSV9+mjHHrvULoTJggWuXSpuFv/EUShRb3rSwLAx8h6ATvc5mkyLhnpjkbxMV1
G/PgTgM/iqJ6KLXuYSLZPP/uhv/U8lBiBDwTPbE0ugCi3wJOAcjzbgDDO6URDOWL
qlXRQ38mogNS/E9xK9gYRC910tMJofcN+35TW7poJRQNzcFwd+YumRJuPqSe9Ghf
pWYSN7OhKs3ewjnI75tXfGnZwQlrFISzUxP2sC8ee5fzInhh23nnjngL7YuNzr4o
ImQTIkmf5i2ZP9liTUxfG5AH6PFg6FNOj9MyIeXVkFQYsXrDrKV/zZxeR8ZkSRPv
8hpnXSo8UGUNvmhqCiUq+1/Edi7i1gyL+sKAgZ+ebQ9MsJ7DG40tOGZQVCmqWIX6
rJxRxNI8FU0r/LAtmbnqLQIlWyRGd5oOx2HhXfsIe9p2idpFdYgqde5HcIq8A3tK
PhQ3/7N0f/9J5xa9JGPnqYIgrgjcPSj5jJ5nr4eexXSDoRzmSHflShsUb7C1y5w/
2m+NUwriFVNPD11ojTOO4MCBn9zlHbQmiAPgGuz+g4+jJ5SChO9DkLu2a9DQhh2j
KQS0MvuwtVcGJ1y+X4USpApE/ClUvW47p4ESwR7bnS184H7t48ZM4y9U0uwh8iZ2
rhK/X2J0MM/mrLsifBowhrWCspuLdl6V9p0QReUQQYBD7BTFCQtjPXUMlcVsm6pJ
KlcjeS2VQ/88Bg661ejtCJV0Y6AG3XEEq7IEz+AU04eRyknUm/bX3zoj/Y7HAJ7k
P57hQRFt/pkzWdcc1z+UmmCs5AJS1uhL3FnjC+EE9qh8P/oamXM1Joqhngw7EPCE
62fe9h48hA/q+QGth9LaAEVuPYnZBpr4CWqbtrt01T2/LDx+cmbDs/cS1a0UIVXw
XkVN7MUfhRgo4i/90omTp6KUu6CZnu8IaE90u5jxQloN1Z22ibB5GD/iTmT9smGy
yd/H8U14rV4HJIe8rH8E6Ehnm9pGAG6Me5cew5HTiF5a3JuCPlJV2DriST+PqHcQ
PKe+IRnnmc4MZbN7YWzebW1SdoUpa8a2zuCoHFGRHoJFPx5y7XOwd3Ek4SPsziTD
ASUWWEpQMhXJ9y3oesMnoupbTqP4wQRzD4xGiocOPGYFGojLKikvUIEBoC4WL9Gd
2AEP3FHqNW0VicPjbeqsoy1pxxZa9tWcL9CbsDQi065bNCsUJXJAKeBmywaL8Wto
ROG+8lTyKWXBnvH8JgqBkZNimHHdchOXe5JFFG2DgbciDm7w1vxzyA6CfBxISolC
lUo6ltgo3ccrYWJGnJSbf8a62ybvWVq21Aq5c0XVveAfymUqCgC6Lyl3OUro8Ylf
tPuD1/UyiLszQlzncfpmtPPKitD3jK4oziVs7bN+andR/hJfT5uulYga74iDkZYc
NlrpjWPstkO+/BN0E2UA7cWF/6RRA5q3T34hIhp1b4+W6nNtzg3i0Yx7NgRgBFA+
GOdU0OarDvY+9jsxCcb4k1RIkeOGUu2QyOlbXm2pRP/44V+9pFXcA1Iihg6EzT4B
DiOjOaMnjw4ylppjTuvlxVsqFgPQTcdinym9DiEkCXRsvg3KP+dLFDJmpcYRjkIK
0s+M0qjvShZSv25gr1djVL1m7R7gL8RLFa7gqw6ZVMA=
`protect END_PROTECTED
