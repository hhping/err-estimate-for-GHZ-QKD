`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAkTWrsS6tokiTQjJXqzfI76v+4KG0/PD6XEqb3uxEzrxRBmOEbO+oyK3wJBHiWs
r3bgMXWN3a0BjspWXIcqJZwF/RFMAhQ+ivhlI5wTa2kIYBKreHOXh9QNNrFfvWIC
YFmq829pyWgofkxcfoBpUlFt5GFfgiQk3JuQ/DJj75ugXbr6HYeP0omv3gZ8d6iZ
l0VGO19bOXmVuYWup9f1vI34nlmgaWNic9/M+umhHsHtJlk6rkyAnRBBT0KZtZBd
naZaAPxSdJ4vZuhgbuK0xeiqPjZBzXS+4ocJ7N/H8g0heZf9d0PA2EmkETTELeis
lgeTtSuKEtyBar8gWLp0xAAoQrz6nAoiW9LO/QzZniLXzMEAm6dFMdUBIHAbvCfG
AvQNcJamTecKCe2Lj/Zn0aN+CYGUoJe50UPmPjZhJNZDtPMXs5rQUqpLI6DVitfJ
InT4lUJ8Zi9RQzU4H0Ip7qobXLDkCrINj5SiqWbjWSZtRNrA0OZ3Tc1y05WlSl+3
Ib7kpAkHJqnqxTRBimCXhBlrLxrAu8jsSSlAsRDwSjQTVgRUExwl/8SoZPQVtjvL
7vfAtFhJ2qMQ2jLgN+N+cvfYZTMZXzjLtWPYUmb9bj91YfqRSPfgD+r1FzOBMwcI
AB/Jc+BfZgyduEY9gbA4stAiQED3KIvC+uuRumoChdu6GJAoNICj+JEF2geeVnSb
i7Bpr6azs7hdfJprxl7OZbG5eyI7pZjUhnybk2+YESfIbQ4vLLfuHye6dLPr/BP3
4yrtMDa9YI7h0TZ569xM29p6/ks1K4u8IqspvlJF373dcK4Y+QOdVOy2jGBJaF1q
Z/mtNV48lavM2ajWvNMEVQ==
`protect END_PROTECTED
