`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRyYSRySYrkLdSS9G4Exzp67v1gz/njCQrhMLmCA/2XsczKDwP3SQx+BiTtGoh9Y
hmQaKRdIMM6VIZHvUFoW+uErcZ1wMZt6pZWk+WpInNL3IBw4vJ2sfGcrKQvbOgCO
GJMbiJ9l6vvGGmnjpp9LMAbPk7tmnjZmVZjfTP4ohUjK8wuWibrmt5fwg/6c3eZz
Ki9UDS8708wMyNANX+eDUqKNt7dCdvT5PKxneALPtu0e2RnkTIf/Ytjt9v7VIae2
xm1/KL6s4gxx26Y6dw0WCVbHyOShMPPnsZskyqQFNYr7FVVGNtI+UKEymlbj07Uh
wo8bwfAZgGJOBjJybS3f2wkV2rdDzWy3JjZFG4R3gdGG3CLW1hw6ds6JoXdPr8cs
3EJ40EASJPAudrSVLEQP6In6b6GbmG4mazPK0W8yOczp0pO14lDxntkz4oVSUvS8
ZWnhQ4956DvFfBmSjn6Rrf374voXMmWTQE8gSzAisu8OL1d8oR/wklD+TnZP7VBu
y1bTdyceEtbVGZVeq8MO8ylMFYYKG3xY02TPPzcpDIa/RrurD5XpE9GPpM98KMY4
5CSfZ6Jcz9Vnvf4qJuIt/nZNxZtv7pAFQ/udlJ1znaL1xNf/Rcj0SEtQkLSktcjG
EXFi4Wltnh3JU+O6mZvaYebDjUpM1OfpmTQXWIHlFtWu61bKrSvcttqEmZcyH/HJ
fwQyNkO6ELMyg++GBn7eSd3qch0PrZA9WRrVctbGVyhdXpdHTWwXUjK+SyUUj1HI
JtDWOhWK5c6g3b+3K6wSnFByUikbTuqfB0qDzCJRcE7SMLUNCeqz6h0ZyWvz4U5q
EZVIjssCSUi0A25kg7C6FibF+esaMFTrUZK97ZoFRpN4pvLGH8MZ8c3Acmvrxv+M
F2p1hV9XXcbfUwWcjp8VKKsKxSZGFJNnBlRZNJlYQBoIT13N8dyyxO0gOklD4pCg
cIa49X+CxD7xaJNPvfODqyIDwDUxoItTsHvJ6J04xRBanXnGqg6cZHtkKG+xxzNF
3mXWAvWE4/ijMDn0JTZNYNoqdI88HltEUZe6nxpoIKjG2GBMX5DBqoyfCf/fxeBW
CGmYxoYXZhjaLbvbNf6ZkaX2hgaV3la9hTFw3G8wky2J613ujBRbSINH1FszvFuK
Bxjx5s10celvrUDvFE/Z2jgQEndUG350wg1e8qV8y39ngdH79XLZB79vx3xveyk2
pfgS7eQSPkmFB6sfyaFrAY7q43nCjlZI9Y3u5wmds9sOztxz6EvcNH0hkKnk1kgU
nLhFOJrlpK3iA3sXN7Xg7HlNlLir/+qdj2awhbOtGMpR0KcXLQli0PtSYJbpnwjt
Y7SkQrUVyHrgDfAtxf5JLiOslj80gpmCPcHb45Eq8QPS5Wgjj8pkdzbdkpU3SkEA
lXQza5fxr9LG3mzc5JAUd6sr2W8sgarjch51js4CLmTxoeOuVG8e4O2iKQB7PSmb
4mSCTDJPpuhurOdWyRViYpxy/Ho3Sr6hxkwdSwcPdzx4ozZn3BT/B7OC7ZDNvhZh
Mm5SwhZyTwF8DI2quK5N+lcgJ3yL5XwgpswKDPrXNFY1b6vQL7NUY8vDCJg8PNEO
U77LElHfCmhHdE2o0lmL85WYVlp7HVK72PDE0OpmRITIEXBc2J9jbR9N5yPNSvs3
fwM8QhR+UquE0es/lxI79Mu4vZ7OqxIyWAhZWZhL748YBnc412zlCyRHOxJyIdlP
+x77d3qMOfVoCyGSH58UjipXnB2qe8ebohMzTYIlHSOCjOmEXRM0/ulQz4zRN5FD
01z4aAc4CDMe6qmWPXFcsGptEgSP4OL8NyqSs3a+nU1D+7lwKlRaRWei/q5TMNw3
crrK2JB52HcIDiMuVZNH5davEpOJkUO26xrri/WD2O2AMBkHl3t5Qjqc25gIH5dQ
OXzxKTkgFuUBZxJ3sVu9zO1BtBu3sykgi8MNr4S2fqn4Im6P+z8Mve/qMDq/Fe5G
tnRwOhNcxcEUpbt1Tn/GXwwjp/lBXAx6UFH1pd91qsjxOTraluLp7XbceD9erc/x
ukdpWoR6r/nzhSgBlxsPwoZ3JT5eqxh6AJJdCWMOp7U8t3+9tSZZsruTwhmYgxGl
EW2vMXKPcMaLg+39p+00E3yYzzqUSGycswsxvUGoSofhLvpDYc3JGa/ybJjncBaf
RhNob+qdJhS7/gNg5GTvdZtFoNyde8Ab3wM26sXBxV9TM6n5rQh6AFL5Wvgy5K9t
aAj+mBKRbiOgT1LbhPJQ736nddyCYCqBhF7UthsHFe/FFSrC+0QqXWuu0dUTr8xo
Qj8HWS4O/XzlV2CBd5K10mTsF9vkFdLKNMIucggBROMELdptsnFPArdHBhJqny3q
W9eP6A2Z1RavIdHXDXx6u3rrOZ6p0DOw0eXC1QMzoMA7V4lmbGExG96Wy0Wq/olz
C+EeArbfrMsLGlmgFvFQIc4HgoIu1IM9/+XkAmVsW3+XzfOO1XCx3I/iyKGpbBV1
QJtctAuKJaL47S/2YXhJ6Qi77Yy2a08pPTkl8yeAxHYuLw+yMg1mPU7RDbufg7HY
1u89v/P/Dq5K/6qxZWHvekMjoFIYtnGyDspsf1XRyx+J5I1w0VWUGOvlUtg3hX6F
gplNCi3SNOyZUBurohaIaSTLvnA8G9jZn/fcB3qwtuoeKB04ykNOlWj5vt+Ap3UZ
qJV7TGMZYIJDQAkLgBtjaRcb628bke2anbtmULCVwIZ/nmOOorasyZeYiuLROgif
NZ7nMN22rBDh9hSpKL5Xb0rCa9Qw1wpw3oaYAx4roYOjjpa2UTrq5X6p9KUrWEOq
jHXnBdvJ7OYopuP/HbiZ14Ht0Po3aE16U9HQKSDWBt8K1jGD6zeKMvxJOJdSuFs1
M/6d7SaEmCde3JuUp38Q24zcd74xVrUaM6lPwUDxyEXr1hNqdm9JOVPZG1MN3Om4
6ArlgSnPN5GA0sNrkFQUPGToCzJmG1LF3vqm5NI1iXyLlSojpytK8vM98ugBv544
6uNyui8FG7uulI1gqpBg4+AJHIINFxiBId3NDnq2908/mrDF8UFR7P4uq5YARio8
/HFXN5qYCfda0zeFVRvsO+HeRT7ygpstC6RDPQrgW3SWMfv/NaOvH+MWF9JUYyEZ
`protect END_PROTECTED
