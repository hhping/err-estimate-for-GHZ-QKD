`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jewqsOfMMwaLF/9pEoWxtXF7uMfzzb1H+zof768m/8XUxFrWo9xrgwwmNzN2ptkh
/cQbLoAbY+BMzmwT0niam93ZyAR3RcbLwFPjjwfrJcCgke4FSGS5M2q2tvPWgrU2
NPhBFBEjfwpFoccuMByDDMd1bzPiOlXGwnB2pjmXt1w77sbdcX4JLrAvUpqtuo5w
AsmeuuY2/uRhWPm1JMR9vL5wQcY4bKpOe8tqYenPpvpQFKFVYNSEQ3bKHCtPRrFE
EKen1j3NPQBrkXSWy/GA7DBmps4eVpXIOidQ1UiPaRqt8VDUQAsbNf4K18Eu8RTj
5mviFUWJCIl9ytdvCdAYwbJTdwUTVQr8sDmUJnvhQzcvv/keM4oYferEUPgVRJnM
9Yg7B70pczG42FS2LVfjOPwXlSSMAc7J/FnVG/RFlIf0y1N7eK7i/TuKc6vUsWq3
nyhKe3ZA1ytwAemKtskqj9nmu78v+Qz7fLrIyC9nDMDgyMl4WoDKmPZtoR3CRVyO
u5GECVXcbtzrT4JMJkxXgLumPkQsRrCTc0mLCtGw/vAyGwnHVucFxPR571zjU8L6
dKZD7SKhpyrGbJxRXebozwMkArpcGCd2KcSqBfRYyyyvnlYv17vl3cqj0Ay4LcZg
0pQn40sB460ZgL3RPNMEOQEeFg31HU1x7J1VU1XDoeXJ88BmPI+1qMJdkBtDnzvg
s+ZWenh9P3eLrODP5yFoAGfwFWGeAaJjYt7BMjp5knWl6mYBT3MoczKZ9rizk2LT
4sN7x89ydKAebctxfgm+1srGScTpstLffzRw4G7I3qXqSjUMSvfTQJOh5oJeQLkr
GD0+eYBhhE59YOnaQp9Ap+TQsPO/d7lUv2ke/afOyw7tn6WHrVwcK26//Tzfc6zv
EwY1qujTdGC0d16r228J2XfqoTsijOTyzRuLJujsU26PmiiygaWg3q0wg2bTBHhr
oK8Zg4d2vz8QMJKWJnlWm8xF9qf/9OazC6u3V/s0HcxJB1i4rASlvp+kaqoLdcjb
`protect END_PROTECTED
