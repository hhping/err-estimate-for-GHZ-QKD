`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2mpgIryJa+/8ZYX35Ii6CwZDLpbpYAUxQc1LSumADjnNxDhrE09QoB9z9+4z54Q
RJWiTba2gHxRcahFHrkHiZqQYQfqXo0e2i3IQMpfXP8saytno1MSUdRLDqgAeif4
FXDLJNssSEkCalia3fsbOMlpCpB9x6/dNwokE76Wl3TvSXBCi5jgi/XMZ+bw/F9S
W0DiR7IFdNYw+7XRF71e7oDyvdkUwSmkT22c6YnEWi9qgGBUObtBaHpzkcx+N2Wp
lgeybHrmeHxkfCi/jQgc3Agnlp+9RwRWXVAlwrGwiFqIJTEPhQaLdRUc4GA2HeVO
yLvZsIDxGhJNVjHtbtuFS/0YAWGkcgps9I6yBZBnHbJyjSjJepNdnvMU+N/tbOYH
MaPHl6xWQYnBIy+BvcdEcAj22oB/t4s7q5A+oaHfsYema0vTTtRON1R+hF1nqkyd
LOSCmBzW/7xQlZ7z4aVRxvw0pduidyZlXfR0uzPD8TYRPSHbo143wHB+6cY3weL4
Om/PrlqXn0fz1sKHxBs+Wa0Ee1d8TlZM4OwHn/0Xf8xypmnlMXNwtj1m3tzklTrF
nHkD9XCv91lLZaoZfkAKxyV4QlkfrJnTiRWJO3aluRA3IwPsmHyMhAFkoc3G6cvm
Q511QUZJNxWo/sT10sNBmOBs1S2N4DgUaoWgf8U6So5Z2oSCzVJD+dQ3Nz0Y/sBQ
EV5Vgaoi63aAmPJqvFlxqY+M2TbxvPLmaYmYoh+zjqwVXFRBIODV7jjZfQ2CYv+6
L/7h6Z213IB0tpCmwAqU/yUdKqWFokF9D6xkzBy+7QQXmsSewYjvI2SKvdqUMy7+
Lu0Hr/6srhz8R55ckuc15tDUoNGNp1LcrCdYXJ6HZAGkcaUsFvz0s+xLxvSnH6Nn
BgK6dsUZ8ib6XGyvyTBmdft0hx3rZ2hoN8hAw3VGb3ipkED4ZeYshYC8zLwivKWT
hZS+LsRzNkUUbZAuIt9MnbQpCtOgqfySj9lM+3cVFc7YGI9TuFDhuiA7+0M9aox/
e04KPjDCIPbRXeeoXNzYkCcLK9aj6wLWTTT5IJUzYArElOcTj2XIhetVrsjZhy8v
KlGde/1smly8jvlRqBGvbQeCXo3B4jMhjFm5xZXx+dIAc6nena246Z1JYMywQohW
Zo15alXZl9uovE3QcUp1lnqzg5aEKj+URo8M0eyilzU+5evnGYVnmpoDYZErcQjX
6QC9nNjeicP6God4mgT29x/fV04lEpzJbTDO9zWUSHpPINUIqCOvRV00KFUSBJMs
+ywdd1K6M/vFobqtkgUYUJ85wQmDCKdU9cvTZFx26T1S2dbsYc0HGxVYPmeQxL7z
fesX1NTtSPTcU0SLI9b0oQs6nTHONKKTztrQXVFbWl67sw/iUYlbL3WZA4Xy+6kt
h//oP5WgYaPVTqXKpKWxrzbfW6NrHhsgg/wOx4MKwthdHy/D5Qln6itqr6bAVzy3
0P9kwGiVOLqASpyGDb+3wd/N6RaUwdSX3kEGqHdUcVAiQkwa+odaNHK0GVV2/Mtz
I4OsxCqhOPUO9lBYLEy1h8m8ABbczyOz2q5ISWPBYnhPws62ksfOSec77uTveztR
lggseYrsW1S401pFEun8GqI/Dzjx3E6aXWkz5kNV7Jb/wPWaPm41E5tlD0fabXrQ
1k9MrA2ascukJwdqy6eWsDX4yqnUjap/Xw2l0PZ1vmYDRdFSIU4tFxlThdlFh5Pr
RPPoASvZsJ3wG19tZEs0tu8a8UNXDO2s+h99NGIfCYqas+NV1C0ZqY+Av6sEQOYk
WB44KdWvTO6j0f/4AUqp1k03gJicnhpKyvEtRciUkpaKfTpwXUgHISCrDBx4eBqT
5XWIYikSHRYONpxTPDZJFNGD+noPK3fSafH168VED831ZgV8cQiBxC179X8OItpQ
hOgD8+OnfLtOSlpL5e7iL63B25nmz+AMZMaCdWeDq1B5nMbjJMCNUETeXBmfuW9Y
EjGfsfznL7JPe7br6uxZWMkw7BJnXm3hiRAb1BUaOsnWdoW9OcWu40f65UqrC+Ow
CvqpAuRb4P5wlYZC+mF59H8X5VPD8nBW/84ZcStWwME9V8PyReeqr5EXy2rhtFzG
AxTgs/ko5rLc52WAga2Qar65CCEMvrT+XYlP54GerTrp39cMJ/oSGXoUPJUwwWjb
MYOQf6ck8meD51yo3lPnx7o1JfpgaWhQsaLdYYdEcGzPvoB6z+vRlLseokjmmpw9
Dz56A29bQTPkMcBtkRBFJ9rKH7sUjrDZjI8Xq2UySrB/37cmKiDraQaRWJV2k/8o
fqm5f/n0H6pAkP7IjyCuTPubV8E9JKexB+RTFk5D+/kKRC9VOkqFIa5n1PBbd4zU
rCAIzXdiuFWmjCv6GYeN/zFdxIR6BhONy+XUFpnpQPH9JlyGIIOkgv0AXBvL+LaP
3RDeBTeixcQdFP96DEXznbk4xarvDOQPLsmk2jvcGTUAEK9dbZxsVKDCbXcTVwUT
O2VHFMWxX+JkubO1ELBaYo0ANpNch3NhMWKnzzMqhUHM0x7UV1QFhwyNAoykfsLj
Q4X6Tn4WxbCHCU48K5gb5qc7Yjv/BePf0dLdyE9qQ6HjgHEylLv93+z7GSbFxzD6
Ih+GQVKHSCbCLNXHklzUaHegwhMdpR9HrqPFAbFkAPxnpYuNG3My0Mp+m94l+Iru
XRHltgXcOtpiBXiwSK1bMP4/aXYinHFBXZvKOK9Wm36zmwa2akFMikAliSG9lmoq
/DGFxcQ/TqLLwujqsi0dr3FjYzwoBY10qIu/tpOJ1u+5ylPgOLazW+KSXhDknMot
ap0mkCvoGDBlqk+YTUtw7kVpnXAsI4HiLGFLU+skDrSfIF2NZU6dvTnaB6euURRB
DM5wAfcwZMFNyviecMHHkrk+3OihY1XcNCN5Gf6SUyxZRilZtO/Uhf1YYB9ykkaB
bsNkKRYGV2PYLpckBS5ZRoPE9Rob28vvPl93hyqCfctEBVYMR3mmoqbKdJCvez8L
uksmg7FzEdS3YUGRJDvgfzhjHK2iCR+jioY4HJ+K+/Rau17jdUJ4jTaXsMpLZ9io
I5APHcV7hAd9aoIXDPdC4iZHBFfE1G7i+Z7DdfIgs1Q0nmNTvBSskHsqGv3x8Pr7
lqrxXua/XeQIgmhupvbjBmjM8hIfc+tJmJMbesOau7IheuvT7R7QNAmDmLK2Fowc
BdheKT9HMKt9mJRSDfLlT5gALVJo0L+0TN6ywdS6IN7RGogVUO1GbY6caqWc66B/
rOJvGxaBe8l1uWXneyE3AJ9VhvM2epDABp7HZQAplumlcoHNJrNkYT+F8b8SI0aH
GTvqklkpzSBGUdPCVXjvOnkxDmKLG5ZPt+oNC8vo+aoc4brBzGwPzqhBo+wPLUhr
PUXw4Wkll8sUk8WhCNlFk2QDUXj7S8nZ8w7CZzkbakQ0SFVBZA/Ku+B+cf1fvawk
1TqKvkDyRv515SgPo/CNMwkPKOg9EK+E7XAScv+nXFy3yp/dsjYMLAQ1FHbe5akk
o3E33E6XHSzRt9mJcgekkiDMb7+fce2+MykzUUfF92AKklPbpiBOXSQvWkLp8ToH
PkESpPGdjez5dLDpufI/YSZvdyWBaCBDbOPJrSO+7ZjY+Dm5/Y3A1WD6v+iBpXop
o/6Dd/VJ9Tc007Sn3yQEbmSP+/SS++ATXOB2zZ+R+P8=
`protect END_PROTECTED
