`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
orNcd1EjhlXNSDEFsuT77Gns480b0SoIl6WAD60nNhjuISLRQIgBbj0suk2o1cSd
qQCcNdK89TMiLFIkioZ6BKnhx7G1/8+/SVMkqdRFiH2K3LOn1R57r+RU41H9er5G
A1WFnrkt/iPpS2dsyu/Yjaad5aDFy2RACdnyHzf8ZIJE8LUB0qbVQGJ/QBLP+5q5
zHqvmhRJEXsAiDxglaP45Q722NERdR+vpM/TvrZ6xXICs343bNx/UZQntoRgbbr0
WEJQ8KQHZ6hP4GCkQjBLN1D/2m8PG309+uGw7UNK6Ut0jlXELNkcWSLZaLoX7Fqx
dvm6prHgFe4oPL9qBEuclmsQ1KAZo+9hSZeQCBKUDAJbbc0RMcwhIefwlM5pwmpO
0h6WBb7xp52BGvzDq1YCwHpggPXn8fgYphVuK/6VJ1ww1FoPA6VlOPV2285w81Qw
WXkgzVhL2+6lMB+OxAA7ykBMWSIhvBKpRbCo31CP/EXsHw+O7h0WxqZ1XCf0JK/2
Hre5d5cYmuQhPacxdZBk4Os2nm06micS1aMsP8iP2DHAgEsHy22uKzQUizICIqMf
zpl9tGRWQM5NTuj3RzexrT67R6AlVCk+mrvaTLYtDTUpMm3mee1xTDR80HY+IYYw
ON0jGC40aG0GJygEBzD8+haUr5qZsR5S7u5tDu2Oi80WiogrpEFRwfPjXHEWtL25
/cwreuGuyYtCEo31OwviLANpgHlbraiuWKGElllch+9kAUEZp5QYGRhXUtvnqhJO
bRVYbQPMOsC8Ab7fFetclx6guaW+AFWgk6Jm6UfvGVDXFefIfZaaL80+R8URU4bz
d09ihH1bB31TnyrfaB4uprHFaVivLCqdw6Ztp3+lvSKrK0mNlND+pXxKyRKXKOmn
HxOrlcPIPcFKYS7Phf/qZNvJZEputhySd+yHdaGvA0cMkHn3K5oX+IgwvzwqHOId
mY0PkTsuh1QDPnnWq6lG381DLSNbELktSZnyoFXRVeUjKRLRMwjxt2MELtdLGhbE
`protect END_PROTECTED
