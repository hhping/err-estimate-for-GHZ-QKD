`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
erjJtqtS+2OajHd0DfLNmNiwoMz8jmii7aVU8XzbXUtV73CbG+5HEB69iAysrg2E
E8rYvK8jxNRZ41Wqgjh5C42y7+2njqOTPw+DLi3Ilff0XUooKbC6m0MBmv/3CDZm
rnyGVOab2yL+o6ZCcesl22ln2vmrXUlN2O3ZEGNZjua+BkiIIq+iGebz7OwyPUs7
T3PsRwWtbPS31pMUH4rTm91tNpN9GvQbq81j9k+zf3yxxCRgZfH/Skt7BeUzxBae
BbA77uN59yQbTJEq/813SwvwdiipSmH17jXHvlNT8vzaqjkCVoDOt97WNztHiLvx
ARwUDVopImGYT0kd1LcxWPMoOrxrKCHByN8JNQ2B8LwZqrRTkdXJuz7VHFE7qOTy
LUhFyaC+vZw/3IDIZ1hWoyc4vxnvka8AuLCUvXhdy/qOhDnYMgnHn8Qf0mr4R+Sr
P/iZ8Sd788q+K8vwxKUvPow+RaiMX2NxTn8aQFArNEhDrql2evqtWHYmdWo04Ef1
WdChyWjxuaLPsQMld1wduDnqrTWlPw38OskiQPHBDSiebe0VuLxaNxcPMl+bQ/dL
K8hNORf7s02f3PvAZhh3EFQZR87ewD/LgWxeV4+30R/hzttlaPO/l+/DDA5k1BrO
YIjTGYk/L/w1E5iL1An3lYW8wJbMCrjbgnHTPGSTd/g=
`protect END_PROTECTED
