`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+agIVoIXHs81So83QDZWXKpwpcZApKOQMcMHc2IpCrwmNWptC9MRA0xRqLJUuJK
tISIgKzjCQqQYPGY5aWZGM3lviZ6h6KFl/uMAkksrvVas363dC+JlkXHQ29QOQFI
re17AR+IYWnJgudqwgvEJ2olU8Ko5AxWNtpSyWoEbndFFidrzhMqJIN8mM1pfNVu
mwIlR7UJgEG4wChD1xFR7RynrxJfywD9Qu3Uzi2WrZZLkh9x96KZD7TNCtPXeZ12
twzFztfBZS4uUktRUzfwfIahqku14Me7QR7QNFBaJ0yeE9hi2+56JiyeKntxeTkL
rVNMqC+ULt0re+l6E5tEQfJnmtsXVkRu5ohzDRDdw9aWX68/7NbLuAyq/C1+pGKC
fcu7RAs/3pl89EJI/mAXHB5Kq/QvXhbNavWafkfrixtQM3ntrYrzpP4Q34JsUl6b
4OG1shRhj1uvwwCmalY9LYmzt1VWUa1oqn+yhFlZQVoqSKxOCQ6omKNk7lh+62lY
9zIPzxMhnxrofLxN4Uo8OVj8UQmf3NC6V7e9KChtGCrKSgqNqc7gvMr90PkZokR7
q0zlT6bIU1wNZ0dBjOaZmoubpiVyl2uZA6CBBrQMadZ14hzlbDpGYZpyGsFqKPgS
aY6oG7MTuP741tLTmf2E1KtPuQqxwQyZpNbWhJczgXTGlXHIwh/PDGmO9ISzFeN/
KsiRauqfkF4K2NjSJZxGUYOFnbWOh9NZSXMLTufyNIrt+CRry4DoeGCGJW2SyjqI
wQGo0+Wg2vPzMiG93XF6X6z8w1hAFyYuUrgsW6s2fN1CK8C5xNKC0AiBbB2mz0LA
tqIgsJQrLKX34s5AQCMbbdlnDeqaGXW8zv/StwxAtdCCdAtwHKXQ2kLAVqvqDCRA
U4F1YAK5eukkiLqdwfx63iAvV5Iq4wlv5tPd+JFVupp4rR+z8lAkxFxxOMXEW57e
AacD0+cGQ94UObUa1JUV/MZsXv/vL9k2p4KLNGcYJA0W5/atDQ3olbiqdZkKyfXG
nzptPSAIwcz7fcPEJxa2XNHVda49v44s3fU+AEmIzTm2yMpBlO5YaSYdXHCyZ6hZ
KcSlOlkmOkkW8K0I0YL4h4ovwGwjj0tFNQAeaHQ9zFblZeT2rq95Hq00pKpWdZ5I
1r2OqJgf9kELCcmMkRaPh7lEln6Q53CB23VOl/VvrY8sE78Q7jivfNiEo59/6b2z
oATturqE88uk0CPAm2azk7arePzeafobAPgXCOc6koQMjhRXTLpPdsXUgMZgeext
PVi2CmrVTv9s5SnQ84lhQyupJemuZo1onrYkyvseyYQ7dZb16HEZuqjS0cvA9QMF
VGYzPN26ze+M0Ay7KebFTHs5mvFqzPTkSAzIi7RAuDwny+d6npbg7PIndwoQvDju
D9ro1mIE5qWyAkXtB7WeLY0l5U6c+ct2ceGkOU4cA1Xkp417GO+6DspOGrLPBLmN
oGepzjT+eLlBUh5SmLjyG80w+jWDxo8Kurtc1skrAkvK4YCTY1ezIk9G0Wibc8+i
Kxm7OgYT8szCoV4wC5gO/hz3TTYVCLbM1ie+l7N7fvY=
`protect END_PROTECTED
