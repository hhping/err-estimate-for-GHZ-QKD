`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6244NSSwkhXwqMEZWssEfjUCja7fGXZEvE0gDOTtkQcIbc/tQlbyjbBlz9ar6Qf
4KY/unxfss6o4ssPQLhPRZGgNIGMrBzFTOK9mnDDDN/QpPQfH9dq+UGwbc5uMM4D
CP+NRN0OpaE6d/+meVaRcIKwwspkRnPmrEB58pNFF8+EUaqePNE4MUTqFOqBmgDC
XWbPrVcUN227owF1NzmIfoMx75vcKA3WXzjpNZI7a3WHIE8NFhydYbT0V0gQU2WC
Q6N8TnoVbhP8u+U53VxpIL1mlD0TNHTWFNoSd8WyzpDZ5brXCHak8H9POD0HqoFd
AVGNatmQNIOxphRqPIX3T4r4jyy2bUe8yX1iXX6LkysKOfP/nDVIvdtpvrtVAp84
NHfxolZfYRlsPPWNgvgPTrXAYd2T7znyE8O19jQGYiOo79H2pO3wCrg5Bm8NqjXI
h+cUYWXnOcKoRbFuHEI8LTLp54EaqGA9F6BMABIvnBtz5+7gPgnjXeasHdIv0pLW
mURkrRXEKjTEDem1Pj/92bWsxociGGQ5u2tFTIwZw+KK9Vbox+/E0K9v18UxnK/9
/looOX1mZFaleCgNJuQxKP/KjcmfXTk53awisqUOsWkH56aNkY+I73aMj3/d/oPZ
9gVwfqnQlh5WGKf7iiaM4iIRRQpsvYJFooJREDHBXNArBENbMUCNablSuBnt8RXe
TxliL6fNupWr69Z/lcUklTbnfjPSmCSI/zFLhYPFdor4lqLuvHlhpVszj48UR57l
LQGC7rrAPym4cYqyOq+zQhqM1HUYUajqNAWd88AEbogJLRZe7H1dCysTmcKwN1gb
OIoEipbPSYAnYHErGluLkdB6zDh2EkBWbWKw3gQ4WUBP9Qq1goTNpgZT7GAjy4FM
J/bMlsOjvkzY+wRXgmjNw01HkxClv6Rl+pKQLy4zJ+OKOi8fixcRyWcXiWsGofHn
i/En5YLIsif0ixY2hehwFvTy1eRXxtz+yxNQzfa7SLVOsIujFyvZfO1QJ/FwJ3TL
VXb5kBrbp7AZ5vk41xzjy+JuuMNyMcQgjdC6a6EbVFM8Q/SCNxFHKWMPekhqYAlg
4MpQrp75u+/CVRdURNDgKbwgW2X6a6WpGwu+P/aov2fAG1lZZYCEmibUQCwvLolh
11G5k0WHmlcXIB/Y6MMpUNg/vhrx861Hbp8KKveimWT2PVp2DV6Zux50Giqjkz9d
miUsl72QQgqXz/yZugsq1rZJWC//kAeWHLJhthvkUFgJ2IkI+ZHQpzMn338Rs93V
IzZiVXDL5DVrDSFxxRIz9KDqKiYFSV7tPUPCm1d+m5e8Dka36SSrm0AWojIa9uAA
/vosyHFTrchbz6aUDtbT7Q==
`protect END_PROTECTED
