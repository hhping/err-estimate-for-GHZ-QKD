`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jmKCShUru2S4atgQmt+BtQU6tlaQPU8+GlgHpkNWYQ4n0h1Ypmn40tGtRx0engZ
iElpXkQ6mZyLY1W+86rzbVyMLOg3PHJj32rwQOIOqD3bZ9EzTih4JDygsrzeyIlQ
dXak7rmcML+D3tfjji/Ao7ovSN3S7+yirKwPIIvOaMay87/E4qNKTHg5xGuT/s4a
6SL8nrmBx+7AvdXKEpHMVSlZ9x8gr7LlYy+DC4e7FvYRRvhtyLD/+X8ZDU8+8bb6
rkzFZUzJ2N5gx2A3dGI+EW5lKusMNdjsTsLkHaBpj5SVPEY+KNjhx39djjHWXOYC
TCzfSRGu0ij1cfwya5yK2Eom0pHGGIDQqLQiKSrDqL+J4MZuPVSvmYIh2CGR7NJU
emDe9ucnEzQC5lQuuJVCJwcRb8hTHOQosNUyBMs1tnsqP7006KhidwD1QNzKkQBT
B8oevnMuF2Vh1/J4WUWNHW3O7tmReXdKq8CjZ9QNBOL9FYkIpKIaaF0EjFGrePdE
WcEZIfZfYgsBufKf4h3iC/YHX/6qkOQ0RvzDP6fH0MPHCWUY4DTzsU11SOuzmWLy
r0yLR3pjddXBszykklii0H+SrRg1m8H4czdr6aVkLnH/QO2mF2SQkWHMSyMiYNEk
sJ96hsHkQAxAe4qAnNn6KXXaGwKDQo4+8Z67fPWqNmpwhWW1LQrpYHY40VoMtjs3
8tGLR6b+h6pJadYQRitC2iGfC0A1nsybhXK8z+hksegHZQUvadqRWlhUZ0d8996n
Deo5/Cw+cIo+NGCIw47iByDXWHBsCktgANBOzuOL9WHUzp8I+tGfPxjY58oD8lZr
A0ayNDicaXt9zQfcCTDQBA==
`protect END_PROTECTED
