`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aR4VbZowPlAb8lkjosVpMv+dAd/Ivzdu6R5EcIoZQLpSymTaKdomgYiJpcvkBucS
Gs6Oc8hoZh+ifijnz7JZXttTHEpwJrP7r0uFG1jwKmY0TuGu9/C4kWj9OZ2JUzcF
dr3DYiYnBXwXy7CP/cDDdI2cmIULpZ6ipbD+AXcn2k1YbODdL83AAjjD0hK16bhH
reuZayA5C/lu8zuUX/Q17gE+W2b1bayG9ZZbeqfeTbeNrYlPlFhcHt1nAxqXWaSC
PWmxqwiRWg/m2dzU9GgWzQPaQ4gt200tQ5TQOA8m46BmAgBLz8E8C2ips8fwlZaM
xxopOSow9vklW76VqIytbN0PzE1U5qs6mawGtKgsBEB4crE9T3jnBuT/4gy2D7cf
SL6sepRxqwsg9bdEQ0RDuZBqDc7kyb5YnTFgVjeYMkTR8JZxKNLAcoZOIfnM53Jz
NSy3vrlLm/Om67EuKuvrnyE+sA3FxDqAYU21HVrLNZEbEgY49+SLt+O6Llnyky9T
E4gBMldMyJTDeec7YDFB+yV0kLOfn5TNUsjfb5KoHmbNZL0pAJ9SakBKeawYaod3
zpNC96qZ+R2Q39Jp0/UQ3QKIgYJZpd1ggqnEQIUOKE4Ny5o+XoWp9R4XuFRru5mN
aLrN0rH4t3wuy4vMlVuJDDvK0IqhoqyjNXEmH73seqUWlLLi3X6VBJ3bBvnKiEMK
29XABrPPfLmlPgxCDF0MQcCvXhVQOZnGPIZc3yIEuzzlF/o5abXFSAIPA8pR2thq
8rQirq7YYO9WjkYlJyJ0sYcwP2Rm+XIM92hjAQJx1nGfPyZuk6LzbBVWPcS5esLv
EIVyIwKVmNuG6mWqroVVQnJy89a07t48v42wmPC2wfqw/jAdkk6rnezhWtrxQLj8
j3HgZWmmwub2UP7ZC4ldttxMMYHMqCB6pHjPQz0GbG9myUJwxQ9ngpse1ojGWz0z
DiVga/qmDJPkmqHn00kcc0ko/Ej4bzbhd7Q8s1P4Aiyh3zpoXIq7CJXoa3Bkow2f
z6k9xZh2+edLXnS/hcLz+TSPm2xcYK+RPtrLuv+2nFUJOcTt2AekyYgToDbaMC7Y
ciq9pNHgVbLybht+rr5gs5Pjp3cFvvyxiFPbx6LmxHCXd5Fwfvt17X/c3tMB511V
QYiMoeiMvFPoqmxEMhepyLF7wIoNdK3AmQ05ViDWE4nH5HO8Mp5Wu6cBPK+dXeIF
E59xfUbRqoqeLPave8aZ/cYDTGOMkhNhlf3GKiK+0XGnPXkXnQU7hruZEfEIr6bT
VZRFSZzUJ0/EUYHkL73GvzuG3ZPtEs6X5bmVE38LuZg3ObNTusoBfDtJrgnUdEqp
s2HmWLk0ohppXPc4FRoua/mGxTN4lTjoDrrsdzjC7M+lrXwRZbqLN92rohTmIDCL
PBrhroCLTJeVoOOGAwL0c2zF2he1sZ4T91I9GV8Jza7HK7a2lX4oue9VCrMGIOk6
gQFfafhip2GRtauDrottWAUTHJOwoKvatd7SqoaB3yUhEL7NBRz6JZbjGXWvuoU5
446b6P6iJf1ojVBwnM+UJbdzfOWZ7DQRgIfooXmnHdoaH2gvohF/7+o/6UW/LVAf
HHOVr55D73aZq9+O2LJvpIjMpLi+aNIHayhBf98eae56l/y5bnCvCIPj1lTDtV1P
e6YZA4pXopVxCaN+HWFEys2IIDwShBPqFgKI4nQ0Oc+676bg/d/bRucu9G2b/HQg
4R0F7QgtAv7Z3v+YddWHPLkPkoUJNwG8Bek5Yc8m++rAwwVvyD7TViEj3j9pI0tL
lrIC77IyznLmFeGamSsJlkni6KUvilZtUJlfGGxi1CiSRh7VpZ/zw1pTa7NZV/yj
`protect END_PROTECTED
