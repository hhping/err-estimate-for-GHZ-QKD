`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLTNigcYSUGIb+/XOmI/LaKbqlQ+AKNgqUVDH7BV5CpyO1x/DOzFZrw4pfad8FVd
YJXrjpHX9NWZ8Izhsiuj+ItxcWr2cXI9vYqXc5Ks7ankJECR6rRi7dCBgpaHXIBb
2sflXAZ7CSRK2Prjc/Ds3UlFzHgu3rwbFqWMEWSFBACPdvK4wNc0zjVntn2ZMQYe
a0nSh32b7hbOPNLVUE79526c5P+fprItftzyHOMIvBU/k95gjwiRtmkYl6NA9nTS
EXO6EFUyrKrrIPsvQH5zkygFink1s5NktBmFPlwmnhYExDFDzBbbkfbrrMLaW3OI
TnIdZsEKxIhY4+aI/xJTGh4J40WafgHFvkpZl+zKCmMiRQfJeFyh1xT/7AOIxdLW
E4s4J/VqIxFcDkfuuUeSgP6ePsC24SojthKZkXMUO96HJ518qhVB0FHvHpor3g5k
yOPXEFCCbjJypI2Q1e2o8ZyywGlMSvs+jaWVU5KM0+Eeb640eUdFY935YeHhbjRL
L/y4KoMSlsEdGz3WJ5U86s9In2+fguQHkC7b9NU77pxwlOAkQLgVpY9g8Yf4yaEi
ayIhfSydUvW3AsZ+a4Nk+bUHXiwPlYtf7Aen+lKGDPEWu9gg1Xg02DSwsukaKNoK
v3zYqLsyZM7Qk/6mH8OJitCtttsD1Kl53OPVj2EBcuPbSAfsRQwews5bJtXPsrL5
Xszf8/ZuTN0BLOXQkt5cWH7JWhb8YuFo9L0mJ9NvJr4aQNM/03Bm930lRez652pg
/OcSk1oPMGAfsugOl6sd9zl9R++hCNK9AOk1UuzFgoQ6A/MJ9xxU6bsXobtxrNGk
W1mjFtTZpqhuH+H2WbJp+di6REtLmiksgm2swW6TgkQS89mRaeFAX+dIpIdctLS9
c/BF8WQId6plg9VnfufARiATBRnKkhj8E+3oabs7JMEF358gX2CuG/UWAT3NO4mU
EWbSNoaoIjaeF6q0HDmJXRNfEbpsQEQmizt/bEzWq4Lm7KwIc8SGfDUR6k1nvN9Z
`protect END_PROTECTED
