`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7U/XaGs4ylkWFGqqzS90x2R2HGgAunULqSo65BCjNKp9awH0ZHLCVBJFOCH/0c7
jgjBEX+O/m0pM9VoRUqsekDVmgP3i8Hc3KHuNuT8yayexs1HgABIPzIv/li56ny4
3iR2nG0BRzAf0ZKKDf5uQN6SDn7CLdhdNmI3FCp3/vk1c/e+7ulG7e4TkjCfdzVY
362Wh5AXacXc9zZeglU97lycAAtlUjy40vz5t/vlric3SwuYOjgbXqH5ydQF4253
kG4kBcaXK//qDBUBMcQ3XglHXYFK94MPLRYgrCacPCvtF/MXryqxdfrdBWy+sqpL
s29PJ7KxTCvekXACYWPHmn80PJEU+ttQoESN59TnLs8srleJ9h80T041r+RZbIJy
9DhLa63rEmqNt3A92Q6JSbCFOJ27WlSMRCuYUiUZ1nAHKu79i0WZmWKHbcPj+x1Y
SuJRtSyRGms0zzKGYVY5LIQWTHKp0Oh3OuwviuGpiW5c9/m+jTnS4tjlYhHGl5/K
NDZSTWqOLqWuXfj4TwsUnlr7dcGYDy4NRJ0uMwVnu62LvthPKRn4UJ32eJWZNePY
G/yGaiQswazSBtQ9gVQcV2MdPacotBu/IFGT4Q/Uz97+CQFOYWh1c+CRW08/InXL
Bhk/xdeSESxSJAdOkXZDceSeTQmcWciWvWw/Zp9zID7uDvv3gZZtMBUgw7MscHZ1
X1i8Gug8nyE56dm1N+e5stAvARSbtWWpRpB54085cH0MmjecE/Dt/DbRJC1bUndB
rqGCTBSfyuo9PepQhNM6HwW8JZW5NLbDFgiTg6lqfhQWr5I5HGfRWYSaqq5V15dm
RCgYA6+sO1qWiI69XgDDSCpzgGgeymjCjD947SqGWJy8yOLc6zjq/vFbUNXy2emP
Nzq/rboxdvTn6e5RU05Lbo0dc+ICr7MKeyHKX6lLDatgJGn1IN8hJEgHZkmE2S4M
MCh8mboRqH+KuY7qZMcQYohz8FGi+6UeJMudH3tC9oJrLjk38ICPbHxg/cQx0gzy
YDR4MPtSVOOCzeHfOLiI7k66FFbelJH6u7/6Gkr0xm8qVqHso6fPxZkuZi9irecT
NN3Yl7QoBx0Bg6BrC/9nGiD+CTHjztLKXpfLbrWumEy+fL4LYLSMq28tHEZ2KZoE
ex4ntEX3kcvNT/mTUD0mLLxzFoDZGCJYYEJLRJ6dUmeQaniaAn4+waBEtO7arwhX
v9kqXpy0+ztrQffU4BdiqGTUA8xwfvV9YEy6fSEsnlwSOzls9Lz3tkwdrBpT8HNM
yX5UPaKd8s2i4onXvZNYPEUUMQBu8KkU0THuXf9uvzvJO/SQeyhkT41eY616qUl1
wU2SoiJZcBBFJPpz6Gefv9dluPvTHVPoia/Vx96WLeA6v+wKNyhRyDYZbrZ1Jjc4
LCmPIzWHG2cg9YKkafuyYsO6XzDlPMbBVFHVQFBrs0PwRQUdvznrTblfYKw2zo+P
rcAm6yIsfC0MKH8k2kZ7qalJIHiv0NbL3LAm4IbFg6/ifT02i/FAeYsRhBvh1imx
8mqYJOn8rUrfV/0Kl2IBhuALRuHWDOk5+24TH2txEyNsn1TwfcZQpcjEggnrEvmZ
Zuv3KpsXD+8/5VIQhPvBZFPtT7vvGINL2ewR9ntZn7yoOt13fretKDHLu9eqtS+U
jfAgNfRnLYou4yaeg+l9HPl7v8XOWDRE7Mu22z1AI9u+0BnjwP9ascVbL+3tKjiI
Ab+wg4yNap2DIC2UosmM51RLiozxndEDI9VDCH9uLuaCuKik23ki7Gbx7aYdl2lf
F0uxs/WPgKXa5eKdR+dPEO4S6oVz+KeZCS8EdU39fPh8FwToiBKF12VaVtYlgitI
SaxF5bPV8tVktMTIEgncviuVBpgXt1v0IIQh6xr5ACv+bKks4qQWgSUTutfaHBKz
dF6thKZSBjAsCw1Q0clmMKC988s6wP/FyaVlurd1IueMUmftNoRUen2lraIWuHHr
362CogTpp7d12MGMsRrvbw==
`protect END_PROTECTED
