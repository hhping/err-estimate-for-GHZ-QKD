`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3tPmrC1WEUe8B0kOjkwq31xBYSx3KMGBcA2FeIxh4dxgMyQAEhgEULslpM0VdRq0
snFeKFSRxpUeiytqB++WWG2PJdA5G//7aZ9g1C0RX6XpUtRrtPwit57+JP5hHVPV
IqavbWLy5qM6Qm8l0uacsHbwCcDCb7MIUgxhJf4aupRgXtDDof9IgHRGmyRg2KVx
gfk9i6IEnhcvbyAP17zMUDx56fwTIjvulK6k6VWV0/cXPvY4K2xFv4DkesKwITcK
KSp3HArS03LApWSim0TDisBlMyFiG0saZudQRwchSBtP2mt48+aULx44hL2v4Bia
qX4JCfiW3DFuDgL9oFwcwgIm7KXrBU68gffdj5ArKL8aZxNwAYGT9BgUnNc3RiT8
DO3EplaO/KRl1Rcnwlt39alr/S6RX8TyJu+IEnfY5FPvWjjCM0cdN8dZCwIqYJUC
C7DfQne0J8ryf51I7oLO7AXnFvDfjtE0o+JWn4rPhYCGNmjYbrQ8Z0i+HDiHPL9y
ANOXC0s9acuDIZVKfv3/Lk2NA9JOw9sbCjKCCS6sZ3WB164Cky1s3Q8jovFfx8pF
elO8ojFEUI/Dlnxc/8U07yE3/sbvpaDaPP3ll0iC6zqe9/R2xUEX2wOwaV06rJYc
K3fZYJzZM9hBE2oqGlqbbP2ma/s53wfaBRvhd7DKsLQgADQaUI4yR8EtH2lp7Oo7
WAuQaKVvUzzIpK1L/OEij3UU3vBQ4YulNIHrC2aGN7ID8dowY+L4vIGHxEioo+hT
hRy6eErWwE48LUB9hhK6nSL/GdwVu2zCtB/Trgj027delbi+0E0Cf7kFxn68JWXy
gokBpi5YaxhOsWkt75e5GATpS9N2rouPwYX3kbaVJ5ukINdJN2pjX3OHqUD1+7Ug
0go+8btL31WAtwzqda4jOicadr+pIkauLi/tAheNroIlNUI3Ozo+K0TsqKLstCNy
qoeV1nqIeAA5QqPy9DFQUjBDA8FT1EQeYGvRszp9MqIOGYYDK3dF+AuEHLM8snYf
j/pW0zvZE5XvrnaKaP/oF0sZAPuzI/d7gO86lwucAtYhBdmiASzSO1YMN9p6CExn
ETiJZpD6dmyNo34x1TzjyqT4Gk/Pnr5Mo0OHJ/LMEDmQH7oHI0yljFbBdzihUZg4
Prfb8rOZRsemqxDhj4seLBo/iACKpYJn6kO+kISXIuPSBNbeNkIly4otJ/j+o9zV
5OUDUCwSUHRWNv8BUlGbZJSGDqn20VUvBlCi4c1WWc9guzSxDSplK2aPWtMqsExU
GEfL0tUywQgtV/jh5v5G80y5TseX6K8niHS0++NyWMctKfx5NdLiX3BNB4DPeXc6
GpuNww7aJvvoeRvtCwjJEfb32i4Ljz2bm17kZ5b9T1KGf4mjNlE3sEUA7UKFDneU
BthIZBfoImGjv/621+mg80DxrybrL4jq3oRY8Z6eAmPI2GCf6voDCl7LYUBA5Btj
4FVTBs9WknFBK7wVbUthIFoKRPOV/KsVzI+C1NOjxiyMWN5tRd4nX1m7ODjCJgA/
ERVk01NyWgMSs7fky0NCQbtV1m9mosrHPjheiDXUTEj7t8uHoo9XGnZyL5Mq4Yqk
QAGo61JSaHNisG53ZHivfeL+gFRaSKzntgFx1BdzS+FFlIV2ZHD6CusvwUN053DF
bRlvv0uL+c83PmkgmEZdjudG4zteaycVv7Ks0MjQf3+6cye67B/nkMZ5WLOVBRkM
K1Kwej4fxJpgf8aivr4O6UQq5n15d2Zg6MolodGJ2/PCExhrPETImh+NXtYdJJAW
Zha5cuXRKOt92YhUIWqFJnssu52hv20zqPHx6v3F5JSA78omOPdZ8IPl5lmBrpOF
pJA+3wkHbSCxUT1QYcrIC923aKifhIg6eSm9LQ9jKH2BF8gxU2kb+TaH0OAWyfRJ
`protect END_PROTECTED
