`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSj9NZjrBHJr+DMlZNcM7gBoTh2jf2nvtpJzC+AIrok2b/TQL+Jtuu7najXEmegG
qFDoolyMbc6ayhtVTI7FF4eZ+5wKHXjY9cYfF+FHcysQgvmOYpIkUE0pzmmPEr7l
c+MBibtJLgmCjR7qfYxovDisKOzLtziQbe87JNDIzQBBozCw4y5A5DAceeXeWCrA
lxgJRHGi+AfpAYf03f8UBNslmgH1cQCI1VJv2XdeODPNWGk6TRkDIuAruzCV+6uj
H9IE8SCWNxj6/B7mfqDWkGodE8FLG0tBOZ7OQc0T+9ojYV7hWlsKrMO1lBSmcTRp
XILe+SrS+9nihgihpB9cN6S1QkKZbvflRS5VGfjDbLi9eVRz2s6y+JaK7QHIV5Ic
b6LAIKZG10E9Ul7YJm+I0P1DJri3fDCjAyDIvqJYdi7eUbiOOPqN5wdO3C2Pp7GY
ECogXXE/y8GlX5QI304KxQprelyEnDQGlhii78zbdSnsnRSuUusgmmE47csMofKv
k2xhc7ac9yibn+iqag1Mz5/vo/z913jHr06g5+MfrU2RAv0YSWBXGVv0bvvP11Y1
EC75WHjJ5XYOIX7x4CH/YHQ8/WibsiI+1DZz/NmIGbB0YUsJdDodPdXas8fkFAua
F2PcBFmdcINAW1zKMjsJFbqtMXwsmhY+DYm6Gzlz6gc2o8JzUvH0cpNqVlO6XPpA
rwyHm9d7dq/sIPDMZFoPsCqMf/c5KYsflYOTFNuUf85pu8DMugYUE1CPt3GwbtZm
sSOppyJJXpMQieqQH06NNMt/U+j1sbi/0ccZGpOWtGqovOGiB8ESKZW6QuWf1tpG
2Y9Nxu6GUIhPQB4TZ7QNLRpBqwhwlzWsq3M2915R33DfyUGTjRmfGratfKaryJP5
gmj0SN6GROKP+owvLtP/fXD/uyPUZ2G2bBWkyBHPKlLF1T6M+u0BGjtcp3rBYWC4
FLK/GGOSzEY4qYPEBAS8k5lTxCEJ5Ywfmez6+q3BLE4dSuuu55iEcAlnsDIo6lK/
/cKjSDq5ya1lKu6scxnkRis0PnF9w8Ygsd3gdSOSS54lohz8HFJH31np2ifRjH9V
yY6ejnCP+hcvbVAZ6SccvewJihkxIhmUSXR7vYsZxG5VKJMzDqesNNzG82a+yrUX
k89K/ma8ks+3rPkYLMtWQP0esdBgmbYvjv0k6+TB6Gm6VvoUKV24MzcZ5pUGTGRg
h/jccTo4u/XT9VgkmpLmSbkoRmKeEnhtyj64kA2R6+3v3ySbWk15owFK8E+uEyLb
CO7ET0/GbQnjU220IvSJAiLRkpsu7vCBZZzfcgqpdp0C4pgBHFmUIghRdN9mR3EK
w9XOn6oaqf6kvqFn6KpewIFG+mDX39c9cUZv4flMpvfvQHBEtKlQpLbc/n+pi/51
k6VVLJ6GCmee86FDdphJfuzp3mSD7UUHBhSU+uxn4uyLy5+7rA//9gswSSBNfSCj
czigEF4zPJilGTDU20Y7vTW2vkfXD/w+KUsI/qu/tbmL14Q1ZmJB1FESiudeLP0i
uEGpk86a6VJsWAcFbMH7Zbzd14LQrBUNoP9lEc1Bm7xa94/p/PyK4iT5bzYHlili
Mh+ODvRLWwGMgREvcBJzH+jAYo98cPYTG+sxuOh2lEn9hbO451qjp6NqAg/8KcfZ
+IHPGfZnuSQNvlf1WiZccdoU1AwfqrHuaimkAKbxkqGw6+fHxfgFKqzUKip146S4
G6O5h4CZeq+AJoQkCGWn2YFPpX3hLBtCj7OQLS2dUhqd+7vrVeR2n8JK2lEiDtto
5jfdZEVaoi4o3GdmM/oDFgGF2vJmVFT/ZRvpASmJ90wAqmvKQ+3Wo8+fcUvTR6/M
k1gQrY4CNtq0onHk5H16BOm7OSxxpbys/sOKYyURVUEAP+Yfx8OGAbAW9hstuUKR
/NTG3KVPGW35AECZYvEvTshQxPZM5LeS/IiBdwZTTVdyOQ20mb43CuUPR3RNxr7v
rVXCsu3lr18eZ3dDChhk+6LU9pskMB7D5ROF/kI7sSxS7OR8MTUQwXrNejn5e1h6
fGd6vchdbi1+O3l25Y2sSJcul328OuOpIF2iKkmys8eddNd0JMn5vJg43s2rzleS
DNIMDbwUyEREFQDl2R/DxBkjqkXRa/JFpoL6ugMrywQOEgNGB7P8x1PqByLvQ5Rx
x/tzveb9/Yd3as9PY6/jL8dK3CVYFkuq+3zbgginlWT97bnougcVdG6aIjQWsrH+
YgMW5Oq6cQa9rDpzdB7YK/yMVxvQiNkd30YzrP0hrr1XJkaj9fOnbKVAQhh762cH
b/weHH/EnwPbDGJdq2DnwoawJR9bPEVnfvo/ZBNIflEB6muWiHX2FA50c19AuwzA
UdyaQBjWyQne/IVrQUZXIuUXwDrKPJtuc1NOWCOYOd+QFk9m5FfaTGbMHyz3oAD1
jfucPr1C3ugHkkxAOOPcza2hvbNC/yF2REHYiLQ9C++MQSl9L6KcxglsgbIWJ6Zh
jxfUduqmaXCGVDFLeXpCqOc4VptpoFGSaBAG+c2/zXiAZIYGsWWKyIC2Jj1oHAAh
npncM7IIF+2U1sFsB1mThtsNG84qy2fPjtZrAdk7X5myOENoqUaxzU4bSf+eJdZ8
Mzpyrq0LBGWSow5iRGKlXtGRKhH+kCBs86QEmPIKqRwqXOh7O9nck9crRbA41fv4
v6mqLuHbY3UmCoVB4oCwk26b6EFH3sMkwQmDr7PWkHVZT0ZIyEKjljxGNE0p8onM
UNvg+mUafK/03P52tKYaixddktTGK5uYckDGbFk93/c6g5SQ3h2ITR4//P0KiMdB
7n+3l4/0cA0/OQRbZ5wOO5mPaO7FUbReS7MOY6qeKuqc15BQ6JVRzc/fzaQkFdNQ
l0ucpY6vNtjyM5tDJ4Sk1nIP57wtr7W2L0u1WTdoy+4Wp49fh7cg0M2bLS5hBkUl
eIwCLmudBk3iHYH32iWxg7KqWpN+B4pWYz/CLbqv2bgYKNPUkwXgbMfbvmUgLAoo
zsix49E+dSS1O21RMZ+Y1aYLeaWDh14LP3NduuC2oJDoAUSRwC4Dco3Hx3tbeuLj
6micuQPwOoUsNzHQ7JyOOc/V7z4Q+gNIhhloTR6OfumkfUMsG7FdK7dpT+S/ARhJ
omd5zXnhahWfHKB2iYc6trY3YDrIfVFg3PSHFkgnd1cQXb0mYcC4IH5tUlZ3ZFFD
G5s5eLPFmI5yvANR5GEbiYf7KHJH25wc5C132mS8aaitLhfv9AsbA522rNkFbCYT
tceZKclsUzpBx7mce08sjyo5cGajREB3arui8ouqU2LxftjQHvLfJZexGkMkBFMZ
AuuGc++IOsYM7YuGirzuYHjqFeqjtsqG7Std2O24xnzBLwxhjiGp9vrsieJV0yhH
f/NPPp/iqllCPll4lUAY8lZAamt1Igch3Fn/q+vGdhuqcHqgF/ijxnrnANhiu2PT
5deWC7M/gqAK00MyZ5GaTnhxooanez0RrUThu0AMiGtykL+pGBozx1ZAiFI2V/01
xMl6zi1I88YdrxYU49j/pyLRNY8PT0DnXkXLyTiVs5HFocN4jxKk1QpcbF75c4vy
NpMRsKMRZzEZiu2QFwrDB30suHFzvJS+6N+opRUHETFz2LxxTRD/ug/pvkkp+iaQ
G2OlybiJKlitQU4hldoMc4GFkX3WGRk5mZmc2m9Rbob/GNlIMy3ALqDISST9ke8K
k0I5xI+XRwcvRQlkGhJO29kc7sS4ogOM9Vo2EFCZONBZjCgFbvJSGqKlE48Uq9Lr
mJxz1RqGxwvWHOg9l1+kFNIjRAMY0yx8S/+XsjLbnubC6/E/yksukUupGvRs7Tsd
+JRz79XahJAweaizy262LVY4aseqIRmTbMeEH+sZaCZA3k4cdvdxVjnsnuTmbsMI
1KsMckqUEqj+cv3txna4YeXtRoyFi7q5O7FHwO6Oi6+bBvDMb8MqXWX4/07h+aCj
ja1vDvavDn3Dc7F2EVsHAbl8kU2siCfpKv8NSf6cKIc2ET7S0NQIyfI9jl8HO2+v
nKGEmqBQQOThz1skYj5LqpEktn5XNCpi7r77ddf/Swy+LN/KzVYQzab9bwsvy94C
Dm0Younbc/jzBMBGvXQGsmfhcUFHmmb77StFAalf67eHfdORcDcSc0zkpZPZjl6D
fzoWHqf7atnnfQJDH7lxl9Mrb+XjN/66VSPfIzS+xab4suLE/cHcHjGz8zclZhJl
cZew9qnkYyJgOXgwWBV4KROH/Ip0IQXigm8i14HiXaqEy8nj5/sVjFGgutXGdgE0
gZO2HoTW6tPAQbvtIMnbNLs87UNS8kudFUVjUhZMX6nkjcBfuv3udAiiXiobpBhI
jvLWmVRA+XTZKbhCilokORhz6hPLghcaXIPFcecmUQM7eZ61yhU6TJvrqjqqzPdB
Hqf8RdFBiZGSzd6bZUgj6Vw1z2Y4Pkavp8ala+pOHV8=
`protect END_PROTECTED
