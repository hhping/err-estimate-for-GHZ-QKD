`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxxC6+W2zkGCFehADJkeqCRCpYfo1YPH7/vEuN8eCGkcw8YFkJuouHil6tcjJ7bB
SY96OZg9LgCszsLxKyzOmL17jVNtYf9EwpN7MQM3Ow/xYjBZRe2hBBrXuSOu8kuz
2u6AIe5ZerCuVJ16PyNigZZddOnNU9v4PAJCVn3a9yvq4K5J9pNtdAtYg8RGjGdw
cWrJxmApYwRDQIp9zTmhnUib/6R8/tq5Mo6Duhm1Zb74ZyxMRkU/KBD1flgBz04p
cMS4M9cJCnewlQxT9rzcM4IvcQyS/SdlHVPgvEcfeNWcDt3qnhBdXdC6lebCIVny
Q3aofefkRvjxOIfb2bmr01MAnYUUprnnW6pvk3BFC5kc0qiiPtny1eF8sMFFES6n
gLsQNPf7azqdbUzBdpUAXYyC6Kjxddek5rv/FTVUJ5HHYxbCesFSiRnv6Cc/7se1
chhyUDUTzcK4YAc+qfVcfH3ic4laltcp+jkHiRlseqxTDZXaZR0L/XOoOES+0WRt
P0C+P9asay6pGYqaEBFa/lzWbbM1UWx5iyqCAzORwefBLSMotnBZ7YahqWyncOY6
7cFXuG+nHXBFx5OD9Tz/PLTDEKQbwpLjyiVI0xZ0R8ELmUNsa6gMPKTTC6BQEOWi
`protect END_PROTECTED
