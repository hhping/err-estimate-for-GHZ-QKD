`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xyNjUevTpg2ALPHJ6DmOrl+ZLmMEDarP63jSuo8v4JqBaZ50Bq+j6G4vDw+gciiK
cwCxY8FWk1VaDenTr4NQ4TJfhSnl2AOGrfOPlaRz+K4Lt4qIBvNCow+VlYTJVku9
+5D2kElxAcyqMTzD4iQuHMN+vEoyZkqzLIJZmHRFrOu8E5zQGQLHdTAnVOpvfEY1
nhFxJ5y6vIVA7Vy1yIhu8xChVURDOAnlG3qlDJUZaXfCLxZ7bQiYKigpUs21YB3g
kZ2vhJoYrZWs4PUkGvo6cVMl5FdfNebstw7+ImOXAPEjr8DayK/k1Rf3RM1lgMHW
uhl6/vUhgCRqWrHGbrHZjk8ynytAdUd5EpcSQSd2djTUZb7NsDa0SE7M2WsPsi/Y
Uv4HiyDa0RuwsF6Hb0HLWicD7HaSoVer6CBFesDczUdfkmxeXKGRcqim975Oxdxs
1HHlrSZoO99+kxBPJKMCu1mUApymHGtarXY6IeRORQ+nVIHmSbnVeb7WUNJT66qe
qF3dciD4GEsgwPHFmL9M0Qx4rjiVOu/OAqPyOAzJTiAH8apIEQkTm77yzzv/7qw5
lszK+yee9Q3VASUXmD8KS8QFif+cFpP1wHrj7L15Rft1QNI+dg/RMxzzE4z8shsB
vve/3vZPwu3H+HfjNwkOUdYZHAj8XTmJAvzZ8ofJksrE5sbGnNaeWVTYoxv7+cmK
DkjMXVCxLkJoEflWa6JKh7AFCMDC1b7CONay6K1ih+5whXr1ZDLzHXW+pPugTwzS
+7U+TEknK/FXVc3VUrgefWjteiaV+MqW4PEY4XsFZ3Bl+hQqmrQijhmFVSCiyPo6
Io5n7WxqHCzdNBN8cnevOrTq3EYdQ+jfUcMzjp/lb57kVf4ClphbQMCgO1zYJQPg
hw7GvTS05F0yIX/KSMKJ3MxnW+/yjxF2mF7pGeAgSLboFCze+YqEX211JOEpkxAX
L1ZPK+b5Njj7q1t9kWm1+Gct+CZD2WlhddAD5qe0yLOs8qAsWH/1Bg1Z21v0b23A
C9w7pApXbBCTZ/7Uz2Pdo4JDxqFclbnv6QyJRPJsswViLIBBHnMGmrBlrqiVMh7t
QZ27IaU7gUdFnXTdZIwvVE1LfUgf/3pQeYuIdE+scRQdYEphS0NmFcgYEjT6nDtN
5g/oIU70ZWoKxSMwRyrfzOcRbfZ7Ag/qUByh2gHNmI8kAb50bkEMWxLV9ixERsKe
MmghRJphYhbu3rCH7nHcG7sg/2eqYxTuzZ3UxHU1EszWJo7zumRoqGYqJYLMUyq8
qoZjehPUYOhMc9zvpSxzzSBv6AJ2FBRwk7FELOxAK7mpq155+hRBGrHhh5G57jI9
EiO1IRBDpm519z6f7uxHOgGVJQYSekEHY4FfZa1SIPSwmVzGMQhvJDuYbX7wfemt
+LLUbiZ70TgIXJjdVywKf4kw+YDRMm3pjev1LY/JCIBv1U8PZvi9cZXSqOPZb1mR
31k14s2z/wOfzGV6Sr1vvTViN5vKOvJhKAR4e0TkSDdLxZp0z2uid9IwAQwBKOjI
mr7ObVHYG8/UrLiO8rSpl6gH5+n7IHsVWShloMOTcrv9rOVXz1vpwlM/BoIiKaAu
LPYmS1fI5/uKsHR/rna63ZYm/bQjPV2zQN4v3NEtOEqfKr8M/NSpa9eeYLApG/yF
pHXw5ntAt4I9J8NozM5kq0DHhudqmKQ8vOuD4bxZ0gXwFBiZgddcy2bO9D/8VoVU
knShr8pcgv76FaGde7uIzOts0jvxN5CdDrKjVdS61SEpwei//+4hXBv8bEJahf4Z
9yMCBUzrU1bZMVamvwhYYX0minqqzb2XbuA4iShx+ELe3moaLS8NvKAiYk+RRXFf
xJxDjIsqfZjqJWi14Yq5dzpuBDFb7nvATU/NgJWk5rrpRgkosWNqJKZSdb91JEVd
GYV28RL23QRvV//G5lIHTOKMolOpQCTIfklGhCC3RFGlhe1qArRMdJbuhYEbiyWY
63/WEEZR3IZI5aoqAhLTbZVg0L4Lx1s0NWmgsdyODyyTlYTD16ekykIkErvzPTnC
Ov7rFI0Sgl+5uka1eKjUFpobO3qymnVR4+bPoS+hHZ9NxPsObmCfpWDA06oxmU1m
gGDee61y6u0OdG8rFJNVwodncNAFX6Jc2YRkZ3hqsEjQMEW2T489Ac/KPoI8q9Gs
/g3vhJNrInKkWaRCFtpGdkGsGBBn8/0DlPdviwekhjLJD0HsxEDs9ieMI7v4bGRK
FB9mGJj4POMtFYDcthG6OmRaLraAq95t0S7pBwClpX82caaiSgn++YNTsIjSWpXS
jUlG0e7aMMjfclk9w3bdxCVBElfKEd8YdiO6wddzwRX49n0KSMpXvbcfYD+5vtNO
qtSPzy+dg+ecg4/pT/5WUeN7t+AbhD1GqifKYdTeem8JFtewrocq7+DkhfHJvqfN
2t7nf2ilK3dcqyxFM2FIY5Q/BdlbjZMicNQsX35pnVkWJ3nutMM7mM6U1J/YJ0Dx
9HTtDgjB2fPWObHGnQ+kCeLrwTh0TTw/K3nb1+5uMcNBlxHoIiDHOuv5Bl2UqYtC
4zo1PqyV0JIGkYk3cFJ/jcIHrCs0EeCVoLoZiHCeQsjwBae1uDRl9gV5KclhZ8cq
Oi3zej9i9Sx4J2qbyDSWvnufHxrT8JaCXju3k9o0mxKEDlTFh2XUmAB+xtd2HPSp
0Rn/DgHrbQFrLApemnNC3SYxN71AwN1pPtNTd0jZ1+fOqzvmSl9hNxnPYI/ul9t+
hxLrJ2ymOjuVJ7+V7ztW5fZorvPru1gEK1ACT2uWqEEt3vJDNwz4A9NHr2u0KCrb
+FLxdas7Sx3jLA3/PNATvaXzEH6qq0/z9/6R7qeGcypRHGP2/euNRQZZaDiNklfb
H+AIz8wsBnoGfbl1x646hTLPtNXIfUSw+LrZepxNUP9F/UK7faeUx/XVloPAabud
W5V05Ttj0cAr8FnxboAXXNLfafER9+L5mlxJhViFnC7VhXKhXFwFHbu3Sz6q92r6
xFtcuoDj3TsWMS155SCZrNsQRsMpkqPHZYQz84XXkjyPspdoTk3cXprTTJkotle2
AZ4joLsSWGiFGVenXwZ0wjTjEGMKMnG9tso5omOiZs2LLROu18AIj0tqqlZE7rw3
nwGjPD/t3goFFIzcLkaZ5utIgTDn2qD/D6RMIk8UOXykTx403po7fjn8acSuUHtb
sjX/JC8sMXkVl50S8IquKvxfgn+DyWeSCjTf1Sha1apHtWs5+vta9+bj/m80aqe6
vH5RWAdGzlbEvoJvxHzs7pzIzy6c3TVy3jf73uK820KkvEMUhK+hIrZrx5f9PSV1
baKcKg4O6pI2vk1OSqo3ojAmhV+mtAqxEGDmDrOnw7LC0vu+8zY6R4yUNGm3vwAv
ivPJomW8frExe26WeB2JbeM74NRw2xozWEH4ezpvY1ICrmS1n75nHD0K/Qnefv0o
IJjgokUAeTyrEFJaQhnopaQoS28gi3SB4ZgevQ4y0A3Vw/R4XWvIjYSIsUiUX0a7
p2ZJVPZAwU5s0AbjQ8KHbHx20QPuqutYiGqk5iiirrEDLgF/wfPeHMpcYF57J/A1
aPBqwqiWc8a2tlGmWOkXPZra3NAaGZn7Z8Tb/g88n7aEiFZC2v8yaJffvysbNHyX
/6v6H7vCM2sNDTev0DgJiCcpdMuRjiVdnyQoovq8yZS1ZTfPFE+EqnNzLdtYo+B1
XrtqEL9W99Ai7IDRq/MNGYnJn1jEPOsAwUvh+8Oz6OrJUrCWQDn/DX8sK3MYGZN9
dbMgDpg1EoZp+yJA7mahUkmQHKMA+npwX/LgSGfomNq3/1KxfnDNEPA/ORPXuaSO
nix5RpF7pXauQDCSeEr5zj1QrfjrpaNooUHDDZM0Bn8sk/KWTEPgrPU6Ac6FHds8
2dnxAqUVDoOmOmErnSO+yoYU2TebJTZxuAla/mvJIrtHD8GYSC4sKgDY1T/a5XuM
WOg8qc8cMvsM3emoz8fgBw==
`protect END_PROTECTED
