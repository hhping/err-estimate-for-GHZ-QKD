`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nsn2JZV+z8Ce/2oLNhN3w4dn6LlcXBpV6emKVNoRnwOdO3dGhmhr/pr8dlzALLGX
UIgnH0Zwc77KT3j9L+w6G+8G8jQ4bJkkiLdjm4/HuWuLetBOnZgXZZnMIOGviKRC
QhuHMPhOXS+zk+mPjMYXZU+8NQEcOycl2cl8xN9KrUPtcVilsLekKYx+vWBYmcGh
S+AU4ny7ebBqTEMow6i4rIOrUuWTTeYCR8Rxg1tps0vpH6t7qP2c+vnA52wdz+85
xn8gfGoEjWbHJQpI5vmiSRASw6SYNCGKEB5m0KFK6pgtZlKi/iQ6gPiP1v0G3vLO
KgX3V1sUri3cAbWYdHYUjPxtULuWlNGJlaUP0SdDUAsDJ1u5hBgc+NTs20pREdIs
/N+KQgfIHkeBV/ti5t4QEa0oXplmjg/gGrsbwgXR3UvcWEnr10pOI+XgixgitflI
qiklcEX+naUvjx0O5zeI5tkYnQDBsQTVOZfVXpXyI/r9MAhSWaPpR2lVES8gBwXB
dlGrJ8HahZ6I9ndYUuhWVSaokVAxb3DNYfiPNWMeOd2miIMtYsf2B3lzrw8qTbDw
drKHceUMbyuiCViUfxIYBL8DwlftQW3MDKI+Y7QY8KhDnVPogibEqgNsOend6Iqh
6+QqjtSLeXiMFkR+VJjCvTlHRw+Tc/gXGi/Env2K2spB+LVl/LOC1EsYXTpSmrxP
vgmxwy6o1ViosiVUk9mVDXs8sL3d+1ZIC4sgj1AWhx7PVTV5GyJmK6By6fH/f7fX
BiX9dXK1Z6xtINpNw7KHVRDPBH/ymbHL4dKEftOsvytQKGrBWi0yGcH4HUuGP3p+
mZEbjpLHyO7VZkMCDGa00bok5VTa35Mj4ulhn3QW1qnkZLOr/uQmfUj7rkw5waZy
ZBj5Kz09fCVwIbzvjsZGsfS8aJMilBm/mP/kezVhYRFB/UdbM2RsFhiKGpgaBLU7
2UmcpPiQoTVeWrq4nIDqYnrlaosKHt0AUrGsxdF9sP5luB/+VtBLUhRa/sV2FVjG
Ywk7Si1Mx0Pt/ijBUXadOUF8+oWEvC4+BZJbEm6BvahyM1rsSxrC3DTjbh80M8rt
H63unVUpFiEE1vLPqC+z2DAUYMWFLdyzKV0OuIvwvvagQ0qoScpOAv3v0X5YlAC+
yQGUULpBR5rZCmVb6SnVMEGb19N6gCBXYfT5wyVtXFPzckbgqaOhflThP0NyvNOr
bPE3ZFPy8HQKsdD9x4EJAKubehektpld82W++mldgrQgnegT5dOQbAoYL3Mf/aKv
gtINIOXRi7lRtOyZpafh6Ly/qighEZpT8QFg0+BTQou2jIE5uqErSx6x1R0Pg3Yu
9TbizIMLIu/WqGSqmtFNVfEuNuCTStQgZ7/iYSkwvYHbqvq+7S5QHAaME9s/Ci+m
S7zgb95zmT+oP5pJ23ZS3xxJW3oZQhux1ZIFEAoI6YXXZL1TnuaynIbpmQdVQuFg
YQW5MEF9U31BfkoIyeo9yuItb0g+bOzi1kTn0yyPJ/lj3vlN3Oe3MkIdml22TpYD
bUCEEFmv/F9B1CTa1wOGmoKwvymkYHw1/mxrHTfsijzJPsunQdv8Am/kMwOP3u1Z
fNPJkMsqRSEu620xvGY1g1z9tJVmR6yTKa5SRoto8Zca2JXFTwGe1rZQ4OxvTSb+
wOJ3iJPRtN0baorV7055YF4qXlXuc7TJeDW9rX2GE2FY2b+cNoWyNFUEfvGIuFNJ
YTFhlHWYkUJliOb885axjJbuC6eYgmjKPoSDrU+PQmX+YyE6Y0pOsadS6v/WsrEj
HzPuxBht8cHYp+doN2Zrz46258SetEYBLjGPQU7AEB2OFKuJ4MazxWo+GPcZLKmu
dxxX6PMtcgMw8vHRhCmHh3rd+4qK5hzBWYZ41IwBwpbLJ84O6JfXHNm4/M9Zri/V
vGUve87iTZ3Z3i24IzLtbx2NQ0OsDejYC12bDs+SUUlMVJ2NL2bJjIoKrLtCAMtT
Eg4o6mdFYS3pTb5tSarB9jNpeXKFEdfWu2YqB0y4Hv/hQQy+bjGl9IeBqcaDBcq0
Pbn7ECVqRClSVXDxoI3B73WKXiZwbzyqGSo2MuUGvw7kPVdYs6JvFhDPee5625pE
zphQNPnpUSz628mC3JVbt1sDUAHLA9Ei4CFAQM4ipyLBybv29jqvdGchqkv4wRjt
V7OucfvGeu3+A+jwuR3raZdaLMZ9eeAS7oZuFQtATRaO/UPWQjjgoK8t1Jq7+dkO
td47mkE167noWQd2SnT2P2mNXLK4PX1HwpR7RWB42lm0wIICHAe6u8vf2nClmgVA
xUsGLZNXjZxqW7qNe5jLDo+IlmEQQUucB2rF5yrK5UCAIvYpFijyH7iAf+DcmJwt
uTsT2kVCOvP0MviztPOC5DxldvT4W22kPL9FlFuH/ACaJr9h3oNrFFkhDwACmGbf
OVnQ1/Hfu4JJioDT2u6E2PTNPXPrz7noGX6BxcSE41YH7/aF62P3UZv5Hby64l4S
9AkyHDw0fzn6BTO6EFGWfs3Kt8RlVq0IWpweD77Ubx+sWvyaDmPSJjv9fIzI9lZk
`protect END_PROTECTED
