`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htfFhYBUdduxg64TPkpM+RI4gymYNiHT3tZSt9O1zs3Z5qiSAwtvce6c6486ET8I
z6dqRp+SHEyiRlRyWFsjMv9t+RiZxslVsCJLVkdoM0TZnxFV32vEtDiDLbOtU4jX
yqeqevmgEbV/dtsfhIyDS624t4HThWBwHgTLoNttsURZFwdnUXOcuHy1mgBqduhc
2+DxXQMXM6Ll0AyV+CAAGTqrQzakl5J/qhktHyIPWClpJaMnc9oNsvnztTQYrFke
b0AFhBLlsVVEgpQVSlS9PHR6kLBXOLqbGfsxefxbo9koD/Gcx0CxE+qoPkgxoOUD
E0AXIqxXVSuu24SKww+KKmVkEZRicrV9L6UQvZUVPsBaAcUtmI4C/SxhkLAvWQQD
VKgw1CtIDRVkneWLniZhhoq0KJLTZoTcO/xhNG5egUT4AUlnyU3MiCd7waciaU2D
v0WA/yAVacy5tXCXVX5SspLvZFDZGMpYUU5QKIkSYZnNmCanKjoMRX2eQQ8UIban
uHQyE/qKbnjgHvSzKUQjumCWA1hZTtHHL4lIfoMuZYR8vlSEsN0sJouFyw8va3Gg
iHejEe7gzxBdylsu7CSG1DbxjuUQRVJhIqh8C8PD+HIxuG5v5wJ9IqDJFw8rfaNH
E4cBG+g6GstJvRoEDsiXbg+gapVVzDilCCBoE7NJXNyFT8+Od1N1HBHRBD261h8H
CtGk+cPULYbbEcCBoTFdVoy7JLhL9Q6K4vRb30R/GsLsSkPXJPAqFOPSbKGubjao
nZtOlSVMvmFPI8fVl5B+bbA/KU3p4yFUsM4v27Nq3knveTu214NCGdLZhiISVU1M
NZ54XZ02OzFgOP80JoFi6w==
`protect END_PROTECTED
