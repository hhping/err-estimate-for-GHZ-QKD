`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMvqYc68nsj3c0JzJDx31cLUsLfA2Oj3GwGtNZ+IyfIG8i1DpOPmvvWCiV84zFdh
Sz57EQaHPvFdcotj/Xr+b5n5ndms5e+coBRLYvtWtJZ2Ml4GJVRkWwtwAw0WTYYh
EkySp5L0xPzRnTPAljas7r+3a8H/9IofJ9u9bi+1sMnijqOkEzAMc6v2Gvf4wH5Q
Xh6hd6Rnumw7ZKbwUbABGYDGqkVI/Q3yS+8e1HgDBaNQn92b2wMcht7ToKxpuvWf
waefTQPbDOtlqkolgYP1+HCzczFa0uMI4BSV08voHXTvUfyV7aloDZe4RDN2N5Wd
B1Ue/TTjseWJMsxAYhTv64Sacqb5G+3sUyPKPA4y8w8Uk0nAJZqpmWYwmXplxsYD
th+EPIBw0zQj5cy1v6HyXm58LyQb5Q/QatpXLY/r5CibN6/71Z6erawjABYqVWhA
aHO5w8i64sedqVdxOjhAE6jJNlW18hTmSyUvwvodFMG0u4xEUM9Pz/ic5bdgIwlv
STnGB8tJkUqSnwK5i9d5Igip7XtC4PArL2YrE/idvEtk6a0wtVweOkQXFyZmb7Me
/d9fL9SZ+89CnOX9kRMWnedZAqvJorRujF7nmJiIKHQgcsqaupDmgxrmksXJKCCZ
uyTNTbAQnh+Y4MBLU7iZqi+8ffq1KGA9m9zPQ3eIOHXVHb8bF30cuweKN8jjI0YD
WfPbEdAdFaxV+SXBdzrUPqwYwkujWYoyy5RnT0Jjsx23Th1GxZgJtuLx4zfvAuAo
BeWZTIfHbgAkGgp7ymEW5GF7yIwoeCjdxs0wcVvhW6wO9uwIRlD+nobohgpBtNHw
jcsz7xEkFxOgE6Lulz3iRw==
`protect END_PROTECTED
