`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxSy82avQ5KXuNTf9CJxdJXjLTjCsAKx1jlJSeETeBzO89FJ7alwCXxHKmLaA/BO
G+ff631kYYoEpATDIzEVFiHStpPDp1ODOW5ytfEYt0mS7ZO+b4RfacwbAYdhYhSx
trjyYP0eu68XQcOIkqShUn2SxA46OLvphOf69p+eTek8RD5FgnWjt1/4tieWOflu
7ouDS6nkFvn+VaSWwwAMW0T6Dx13ud+qppcLDh1jb3ucq6/JJMdrcq1DHhTvZie+
5wtroN5xvZqT7Ubr+sSUr0rT2AzL1DF4cinB/OGsq/gRKns5z5RTDS4Sb+I0kI6r
JzBSi7+0f5a4BMECdy8bkLB6Ua6YWV66QWF0RWFjbQC1teGdfo8sqDaNwFrsenL7
Kg7HUUDCjRqmJLyy2vOwECa7SHbAc7t4d93TllLCVGHbgokggV7u0Vx9MiWYlA/R
AUG+V5ejyXKraUvkGn7N0+fNKtE8g0GL+2EjQ9HO3NrmNUaRtsv2m2KnCcHTnSwb
W+8d0h7juoLbeQprVXYcpVFK0SGJvYc3BdsDGPPHD9OXc2l+Qb7hWl/B9vfjQ2TJ
l+vXNJ9M4IMgnkrSF2gaWPSWGEQ5M16XNGjqatuR6mWTW1VPfIbvTZK2KcZdPNa9
0FgDCDL3eJO4vb8WNXxQ3vxOiB/IRwHNT18pBQUOtYQ5zyrzpB/Uj/2VWsui2GzD
cEBgMrpxIucRV3VoRvRcU6Z6x9GXHCtC6u/44vPLt5TvY0/iM36GjrAxkUH6J9zD
RI8Oxu30VlJWtN+HnKHLAnMOS70/FI/OP3adiRXMIMjv7KZ4EX7xD+UmLaSn4JfA
6VN0zjuLVGA+8D0M24E46wS3J2SHEvp5Hwo4Zn6zJ1mKtjUzIRhDWg0R0q+2ow0f
k7Km4VcEEWFLWcaa5+KZWF+jVt6xJrXYouegXmr+JkdbJTlDTLyvumUT8aHl846d
JLTtED023vTv3e6lvjvtJbdfGv3lGNxS7aNuQ7aaq2HB/xkSzPjBiK4kW+0SvkgK
KpLUQmWtxRPRYnmELd2Zuf74DkF6CqyDEQ1RZXbUEYPb2RVDMlqJEDAlVoaMyV/p
4ofDtjOFnimkDKJU1Miibnh4UStw59R30Uuv85cl7gK2PYAeqbe5MWtkhWg5sqJp
sR+1p8V5LmUqxU867TeJKDruNcY96Pvf2gaWmQm4xEI=
`protect END_PROTECTED
