`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zm5236b1+OgU5Kj2GoqC9dbwp9Dy/m9lmIqWA4ZzKzKl2TnoC9SJnJRRDb3uk/01
agctMVm54b7OgE63td8eQbA58t/Rt+uOzMBFBUkrlOJ2Bm/g4dMxy5hmbho8XZdT
3YcU3mNsVL+DebX7/eU9D1PQkOcl6FmQiTT9UHYTagsSRRviLg7TwAPs4zufxSEx
oq2OdzMBisLu4t9N45uzI5UaARpekIzKTUdw6S7ow/v3/NP5T02xB4vTjvYHB7LB
g9NK12g8W41JuCZ64pl/wZtGKs0hzByabnolyxlxgnkvL/F8zpMCMlqbKVXRbMxI
u8LCD3PdiufywCRZ2RPcKSmma504gaNsIpOUs756/cs6rcct6vEMbZYHZlJWPbk0
KAmV90Audy6dtsTkCA7HNZW5Q5lTaYbWCY8KKm/wCdyra4S8Ip4OAXdsM1U5ifWf
6bDTsxxNvYj6dmaQcX6HyfSwR7hqNLt8r7BPOogU6suJaDok3Ob9PDnhMgnfJ3om
e9Ybdr9kThGzwEls6j6e2N4Ots0RGNa/E4/vCMQkpQnuEaVvhU4kP7xgzEAOk7FX
QWaU3uHodp3qPuxk/ytGVUAs2dAqV9mt/eCysUQ37t5u2ymi/+bAuFIottECtEjM
CL3KJHYCePLiDaGTMUBMAfX750gOqCyg+8gq24ZZfmWaHTepxT9ZIyEz9wUG1v5i
KTaTKOyy0ct06inAL6GC8GZBSWSlc4sPFkstLjtbW0V3BxdAsYWKJR/gHjgQ9rcJ
EdHGfv7ke6iZEkUdndUDJG0LG/JiTAAow5qLMaQyYo8XdvtHnk/fkdVsuVeS965f
56GmTKD8P22fWMBkNn4zLSnYiXyx7yLujHtQxMBX2uBBMOS2Th+X//pc81xI23Qv
ZZMmwx5cYExjHtaqVKHNw6PIvwzels0UA6BN3FUrDguoiPmz9Vd4OitrS4Ac1fth
0tAxKrjdaC8FCzGA9ryftDBw0i34KPNvIeeFTga8nCDqsfiyY8ERC6+T6JUT6zjG
BPTZLwUPR067dPIEtdRqENoaapBNhRoyJfifA2SmUes1HcZfpwEfSCm1+i165ITx
mmpvJKpi6xvF7qfe1QxPs82+WCoLMo7833tsfC735qfuEO1TLYby49UAoZtR6zqL
54c1VPlsy4qRXb9rld00dyLrV8z1C6WizLTb5rBjMLkAofpbY6QMss9rQzvHZu1E
m4z9oGDE3nZVzq8A82ZSE3bnp8ANsNGTWvSMc94+L8PhdX8RAJi1WPZWKbNH/PIP
doOVubhDgh8OFCf5z6Gy6bbbpK2ZIVEkwFG+ixZPCLjIEQUN5uaWUD8WonKT5g4V
XPwCOsbdPLWvYgsp5XIwRCfEYpQF/nWMUr8KY7X2kre3GDbqjkVqI9zaFtjseAFA
7DHnMYNYcPNGHiFLLIzCsQ/mQl4qPb98dRAqSanZxzjULGOufRFEeRmWCF8Rlb1I
9Ye9JGVFmnTsTjmQzV0WSc6ypdZ5j0RgZ4aaI7Mv4PqnqPJogfByubZvXKSpzlj5
rBKBPuaOowtnjo0tQozjMxJrX6CmPdlk4Af93NYNXgzgFN1jmxszHsixEYS/Vwmt
7A/nmeYLycStVy1XgwWdgO7VhfHcSoF54eZZO4gDwCMUaKHaQQZZM1cCK/CDQhzF
Wq4Api7I4Nn2BeO4rwR+heV0ISXR3E8OewnhJQMq+a8q2uMePD0RhBtspsFK9iRP
LEu9q1fdKbRXkKzpA5RnnNmoo37zMAV/dIJF+Dt+V43S6O4oxsbV5BTNCmoJ03PE
ynkj3RWU+UoaeFcVM6kVZ2Gcbn+XJW0URhVcMvt4IarElsgYTa9IEePSO22U7gNZ
GyjWcMG0oocrxianyHQ3Se3TfZiLzFRyCHMQEu5ilrQ3fIjQEL4PWkeJTHIyPt7L
xONe6hNBj/ly9w134/O8t45pCl9HekH3W14d/c0sCeU4OzRJa2G+6NKJX2Wzhg+7
Z/7HANxT5hN3vySrvRwg4WRM3qTLvto77si10X+glsOtF2fcjbyQxTZKxXPU6BHn
d318eXQiHn/MYv48p+/TpRb6budCZfOQd46XdFwHn7n0ZRBIfnkzZGGpB23JduI+
y+huk7f+b2Kp8aPyha3afKXTzmP0ivz79kaw2HTRudWhnObR0MqWb544mRGu+zld
KCW5PJX05bbbbOjCqyhTgMFXkYEsIunrmTVZRd80KOT2QJHjjx/RA4muKoLwRc4G
ouXEp6FWi5+5d3UTZeWTevSofh8LE+3/aozT5wJ253KK8auHJwrDym5/bg3SOlhU
leCM7IvOyCUBkyFRiJ+dOe1YP8yyKUIqdr5kNQrBjjh3H62NUSwN0OHw5RSnXqPj
tI/Yaq3fCOvYAgafLZ9v9fPeWzdW7S0OL4IPVH+opExCi7b+fIgYWU/jPe7lYd4r
V/hUpBtAsH1plcHjYUdkSxmKhggLcOoaSTFWhgeapyO6ETI57GAHIvB7/jIKVIli
QLxLYD7wMNyjFKkiy2jVljPVD+wPym73aJxx8cW3hgW8pZmluzk1na82CLkWcf0E
GkkAHJyPQbl9hmmma7zlWtr9QF9CukwWuqW1mTeU7mcc8zr/plLt+FM04YMUUFlK
4smQ/WVwW3l900UumIU4pPSbV4+QTNYI/gPVk5HXo5AAvcYqBjb85qMCpsMKApWY
cRCOD5nlYMLfrIJjJyaodODs/I9vwbDKB2r/xkaKQzurtH339vCMq7H1uZ43MVb4
PpwHtAmKwMo2L6SF37ABRDxQk6wk6BfOZntyVLYTd5GOab/TPyiZDjAGoPpfj9lN
cn9jF6ohzeMxnBmpK1jUVEtyqKEZ0B+M0Szbixg3wnguoIOT/0sOWsTz4RdjV4C/
SardfPjOrdfSdm6V0ijuI/LpIFQI40OWlnb5Lbes/ps1WCV0lNBI1AKgl6OOfqqS
kgjpHsoRAvefc1mag/AhYFEXbyOqO7htxMs+8xwXNt7++nz0oaAayc80NWa7Ew9X
cD876rJlSYY4EslSnv2rOAmg44qyvDlplNfr0mCGmpn1wGQkOGQJxO2lEWlKJWfA
po07jp4+e2XWRyIJ7Ur2l/iw6Y55/cJIFiXIUT8nQoKdaKtiPqyMDWO/VrleEelz
PuqgjtQqt5kDLK6Mc1dEVoB3MblY6MqjeqE3fwLtT9pwd3FbThnop0DLjJHAismc
LqTew2Bsa7oVhD4+SzGh/2g248zkDpRsr3HchxigpG80Y6ezZFJvDKx0jfvcFOu/
4KIx3gcV3g8Kkh5jYF88BKi1xQEE4pKjLpFFjXbbFqO9oxEoeM39PsPz1RTUuTXo
2M+FDO9knUHUMFYEyWxHdQ==
`protect END_PROTECTED
