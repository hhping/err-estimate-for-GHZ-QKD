`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0orevju2JuyOLrKohYchcRtBDApl8c/cOqLDvAYIjo0rpv3dBpsTpkeaHNeiSZt
I6f05uomYyK8g7bv2BTHWarUy+oCR+tGM8eSUpeKMH9pO+r+G5va1PQvmSbj76s1
olK7dCcZ5JD3lXTsASk9rzws1D4KZiirNPR3PM3vUXPQyUo/VRJLmAo8HgeQlufU
PQkif5OtRRwoK5KRe+v1cE3ipbp8aq0EGQgN3YIEqO9yTPQEI0OKwxCRTe/cOicr
HB3PmWyTuygYyYyEQfVfuEuC0maOIv/5dtT/aRMBH+be5K0fsL0tSBQyGb6plWSe
3pWo8sydb+8X92yCw7y8KZVkI6qGAdCK03sDGyPUU5L9zasqENVwaPWFso/KdGAu
fp5T0V9vnwu0naNDWPdhuJWVOhQu208sKiBKFIwh/7jcgPeVp21SCSTWi3OROD9L
WIFC78/tVWTol1J018vl0LT02jeZTVCjoYLE+1hi/xJwycTW4OuD96hjeweeopNk
p6eOSWJDuwqyIXau9Eq0/BGYZaQ72wvS0/PMMwu1B7vmV11GITBdpfVV2IKQpyX9
JCydjGBQ1q01c7iRj4OfcxTakytIbrn3wZ+wWq887xH9ydMCwDaV5zJgVcGZ5Yta
WbalnA9fdzIGO7eFfLE9I3CXGcVF+zHiumSYqEV7q3gmNZadKDjHnDDPP/IECbj6
M3PtXaTQ56epmXvcwdvEN7dWujMPQFOoZeDq0gHwj5RPpnubcm2jxhH6iJzMtn7d
eFqhbBSfR/QWp5bQsIa/fRTxoTDisKDmqY9/t9eQixS6Pg4xSyTCUP/hye40KKDk
6CuHhYHb745LLJmW2KeTdje/CVUir47bmmuKKggJZBCAGRqz3yohscHxWDdgVjT9
bjhAUV0bOaI2thMOZv+CMpWeXHcXnBeuoXArBJldMcY0WQGFE7XwZ0ggeZTpu8w2
QoxBwOwhUfo+u6Zk4mozYDPmve+rDe++izbq1/OoX35MNCcwXJ10JhqaKcoApuvn
Dk8bxb1EYtLInPl/qKLNZ+T1G9li9tA7zwmiZouxkr0j6o4jXiQUJFYTqzHztke5
r2lC6sRoe2k9mRSONS5K1c5KMm6Eu4Z5QSyhUjZM3y3x8R4bucOfwIjmd+FKySzf
qI//q/BaTlHCLqLZLQPT2MukR+HPJ82e3UwjZgye2Ye6CQ0IqNExTNXXo1puj46F
FRRepF/FH1BRFM4E7tZ6oexq3ojia3huKOOrMR5vLihlW3P4N6gx6+qsjU031hLB
krL3i4eabKegz3KYljunYD2de88e8v7CNFiUJtTZY629dAb5YoaxZBnu2n3uBXz1
C7yolmF9ePclLG0wERQob+9WJAjEc+n9Z9TCcB6NMddtkyugPzSznxPj1ceWy8Ig
1DhdHmFZrbCTKAJG4sl4zNHOeUTpBRbXxwoK6VbwbdGJqgqGT/ECtDe6mZchlR8a
X04QZXfOlTZki3plrAt1f7G9lpgpdj+15etDH7D6nG0oWTo7EGsR8QQtETGDF+La
wxrZkhBu/cJPrnLmxjk3Bm84kVyaaittJpshfxNkZnqmqoZ4emMm/fDVazsA96H8
bF/93b3j9PytrqGpYfK7QTjWZAUafeUHia1X1PktTPDptoPJkkcaCYAOBMKqyNaB
7gnCUgFVZOkQ5q5gLCm6YcemvIdD4zUVMSlACEwm3rbLA+q6Z0DS0zjXP9pkyejp
8ZbAncEVb0P2X2aIs/Q8PvfMSfc3Cl0UYjPNSynYDhgjluGGyDkR2Zxm/nnJqFMu
2l4u8W6ED+iqjvptdAcX8gWgSQwQRv/3SYUrm9Chjvbe0UYjkldveLpryZIUN9Gr
1HnScxVjaXP0pTuyliX68+wxeCmrIWGgeSC3kQcq9+8nfLWzwmx4dopq6TXmeUrj
dcNpgckqK9JhwBdFUY+MWxtc4PbRTmi32VZv8frTrX2aI9Q/ddMHM+dvqMjgzMgp
MpskBziVccgYUvCJB25VC6LrdYnrWfIlLttevwCpu7I0f+vMrcUlwHWx1GaBSWVV
NwFBZyQZkGxeeqgfLhvCbmXF5K/8xIOr2ZeWpCzWvE/yuoRROH0tdL99+wmWNyUz
WlLK1C2nRXZ/8Slxp4wOmTyAkavw04mzQuLt6pFMtR6ySxRVeFaSFzGNFMtRR7a+
b3N+M24GicrCmKIKe5dTnNAjFXdGU/udZYwHgjdzcLczFtqMSL4NYJdyBMd6su37
t2lmG86eZU49Vtr+ZTuk9rsigmEHyhc6Vi1WiB1jpRLc1IY4K8iJJDlEr+QePJby
GxlEHUetmHt/Nrt70Yp6HFLpChiKjECVF9x8DNMAiXLJlBu0sZbcpxAYzkcSaXhN
+KE0tQXAM+7hZI7VcYb1kVMUIFyYiSsPVyFPS3zuM19tU4XE1mLsmXKXUieilwt9
c9QlrOeKdgIAWRx/5TlSIOeHE9nkvjo9y6oZYN+n9mZ3W5o85479wVHjwzJF+Pgq
811AlkfVEUxvLhIimaO3YQ1MMF4lP8Jkrg8T+WwuHN6pf2DAE65JBpONTB1ae6Ro
pqsT/ap+XsuyhzqDBITFaEbKFEqSBKDk3miCQOsd3r9PRcM3b9+7QNWcd2849c4M
C4J2sdPXUAE40xXl4vVsj39ruB8aJW7PA/IZ/ZrbrfP18TPPPXxuGssQo27fGDdx
DgdsDPyuXNkiJDKMFnLrLTd0X8dKH+/IbpXxYtPXZMTn2Hgt/D2jSvMRANhgIgAi
/fPGgquAihYOv1OMv8pthoyM46tSCoUtg3EUY/4xeNzwXLsfWOfVoZcTfgIdWU0y
UG1MT+Y9DU5TRfZ25+z70zuDUgN+ouRjSu+iWSSPzjyTwwFb5s+23ppKoshj1/Jv
y7Ujfxmaz2MMcczjklhxQb/Wx0a8Qdrl9eN5swOpIk1YA4/EvAHi8TwQ4SNMXF2k
vkOGRVIIgbvSJrUsNtLqo/LWAiSgYTiBwWQENQdfe+8sPWG8EcYT5B/E20wTC5Vv
bhW+zMt+lnu1Cist87ccjHWmMQr0oI/gcMrHmYcKdLS9zKS9d5cjPAghGpexAazH
h6750taWHwHHVNV4z6UdqBx4601rjq3Je/xkQwXnofzbWYVEa7aIhljTl44akQry
CBcwoLuFQqsrBSFMMreVVdh6YXlapO6YmaqkPbjEos5YCka8jw2u+8RVflzTkdxK
3S4AUbVIceJ0789aEHcQ0qmd+rvXvyRIy7GGsRxJWcrlZjFGwKXofjIg0eor36s1
PmwUHNiohcv+IBDxs8rHpjOQSpXunawW0z9T9LUP1PhdWkx2B9aRG3Ikn7O4AE9m
Jl/hYgbrefnQADnLNCt6+weHLw0mGSsOcNFaMPVG9t9Xx1YzaBA+9SanD+iG1WS5
q88Sg+81dn4k3n5WmjLiiAgG1U2GCMXRHsM3zgfhnosTJ2c2KvTqpM/Q8fH8VF/B
q/v2FrVJPxsR1S6BGMQpdBspWBpOWDRuIANAIgOBCvsnWcGG/wYU9AvDar2SblJn
0HmY039OQZSfLAVT/jg0TTwDTBWsuDwDAO5dLW+Snzim7/bnOasuI21AWvt9IfPC
Tu+X584TofZSHm2nxJeMrmJqMOQWF81k5yJkKEk11TImu5EIx1XpMa8os3UW70yW
prwAH5WcJeZ7jh+eohDcBpnExTBK/VI5ZqkQbH7jYmruTisOXNGohfTtONcM1t2V
lAmLaumjVOgCJjOUpBDZ3fu5NpmVGhlP+S6KbqMjK8xVC+t0ZVqBXs/AILiXHCNr
JsZGsCKPb0OEewQsmSWobRzJHmP3emHq+csJ4iYBGtYByJMAnMV8fexYp5tGBNWC
Zqo1g6OkjzBGfy2xEsG9DXaMl8COBlccxpee0MdDtGsUX9AGz1aTIQoXZZq5OVQS
1xvXqXwkSNmjQ6DO4u+MdS6m+CvIC3XTIlsL+ODyNTxZiy+UZe06aw1wzaFCL33D
meygTusncNl7K71Xals7OMkqqAdClhFHCjGoeWuguEglW56FZhnKkabcIelJO0/9
uhBczyTxopmqonCKg+yO8pplYpPxqv6dyZSKMtVd0GzZ7C/+smlMm3Xs+qJU7BZ2
C9IjA64+3aCurxQTUyg+9EqogT4G6chuCZDGa+oN1gpI1ZQ1qCNt+IFe9rVyJrMh
Ph+DGY4RGk3ZbsUyyytTgs6wMyciiwkvyuicHscR68nEH/efawIHPd8mB1Gufwig
k7ar1zoehzwn9F2gHzdgeDhXOoNesY6J+sBGdJ7RJHL20pS0hJMRszveICJVikHb
JKZW3eZNeG4MbWytt2DeC8Nqmp7v5npaRvozM4+8qDz6jc80kjSv7EQVVFTjX4t+
zejnpSwJC6D2qE6dF3v8/w8HSdi0bnowjqOfBXhHTRlKZWuoal6rOLo6tTydT5R9
mmbIYzwVuhlbmy87YrofiCmQl2GD2lrUVuWRAmTbfE7PsIKHmVTGRty47fBuAAKg
F7oJpVJqV+h9pc/uWjhH//KYTEnnz/ts7fw1OCVcVfG6nM+3NMkVNFVzG4pmnYYr
qUENIN9Xxm7DwmFslPWgo7ImtOAdbqdPgN88sQs8fz7wjFZP5pZFMWnaZaUXoPYL
DkMqg5wlsMwKL96md2fnpUOOb/uj43us89I4zKM1m2fhGzKHi1Y5/C0yloslq0I/
iE22zsiS60FeWRie6wVUAfdpq8JimoMX8WpIbsf0riVaP3eE9vhLdNlPThDY/eR8
MWtistAjqYeP8p3lypwBGwFosdmSAFozt/cLHvot32K8AnV6WHHjUMtmXf5ew1DK
EGpRSGOTAZeQ9JNp9iY6wYfEPBR8Ug/l9lfKmo6NxPMBAA8HBP9+LMHK6mr8+xIe
gpDcKh4mxxCmJbDJT78c+CwOhDYUvHbwg6sI9t78gjUTxHEUMfuPoe/JQqL++kon
7h94YvIe0qDYh+ouBHdcd9Je21Ec4ppZQynR6AtLDFhpQ19l83+r1/AjN/o2IUav
j0mqj9g6OwU0aBGmJk0vlUFt9S+X5OR1R1r1WwJ0l1dlPk7tk/8kQbj+ddRjroM1
1e97+hxANsyMvpZISUGtDvS1CpwHJe9f/AiSrP9S7+OrUTRt0B+L5b8migcanSxg
dJMjyGDLomjSnYsmpBDg+cHgllUfBq6dPYZoePrReUMovMTU5gJgMo8Uom2nQwDC
DIRzt+SMz6ZMhbG/Z5ke0O+LvznYYu5n3DcSFgLWIz9DEm1N8QKsSjNu6tQBR3LS
BaJiV2qRYAh939f+V43mVkisquUVUmCEhWt0ITtMqm8LKHH2+AaFyKvUOYrDTdVk
l4jnaD13SeWK+09vD3ueGzYp3dY2+GCaRdhzmoCsrQYTUetHO2yC5hrivxfySjRh
Jxkv7oV6EqILpOa4Q4Eh1oYlF1v+02dSiHclswoln9DPFVNapDwsXGGdW+wDqw5F
C8hyZZkm7byKKFZzVJokr4MrLjuqDChbcFdGZADJKasMUYEF3HV4aQPTwm94WyAZ
f1D2Egf7ocIoiDuqaVwtuSNn7TpZkiJPIa3c/+ZCa62txBham1JTY87AqEfC4165
3nny/cRKO2Acz6Scsvl/qu1evZXYFbhdgVMU7eqjQ8rKKuKH4M8R0Kw5yWn2purY
vWr7aogg0axnipiz/qJCLkr2EpajojxOvMj21tcLlHmMojQTm1FaSPL5CfAZsbwt
0lVIJXjlsoEzce9VhfHPpnTlkWFJyimwcohcSic/IUmOB9UUTljQ26k/9MHsgMQp
zNeNJkt05A8M6XCe5a0OCGEQa42BP32jiDMLKd+BZ6KBaRZTAEIW28p3bxyuoHH+
QDfyUgKuiO3F+xSB9qXwMy7xBiQAWCEE7ahG4Vvz9ry/GPOFBQf6wZnUscXkF/CT
KyUSGtVh5rq4l2pe+lT9dMceurzzx18C43I6vBfVdjxgRSIskvymGx/DrUN1mqid
MWMAH+F/bqTFjVZ5e7hx5nIZbt6rLsofE7oB5ic7zmZ7IOLfSldjE635dv+DmVqq
JGNGpUv4o1lSilSnKQ25Bd+FgSarNisPWkQrQw2iFN1D0K32ZRxizR8ASAr3uXqB
jEEUxPRBj9FYYHnCp8WEaBEDv8RCH67Uugwj1jY8BtmzuPDEL0QfcKgMScc2vH0U
jmaO8A+6z9UFPzDzU57EC9tGrW0EiA02tg0j/Z6VY09w9+VCzevJj5Ra8zF16NUE
Cvm8khwgu21ns44amZK8RYwMOyS9r+WB0b/FORE/Az1zfZyTpKXLCt4/rZIBz67e
QAcCQ6MDVYMcnPeVkaYYsnv+dalytGjClBA7QV9ZV7tNdaa7UQJnHPOewLnmotEj
+27HHqSXJN5dFrWQkBNp/kdv9m2eljvt9Y0x5tveM++1yJz8IFdstcwjuHwlIOFJ
/c5ZcZTnbaRV9Zr5EBOFGgs0jYa0iD2WJUhghqiE8nCP5VhRe892XN4zkdQAYgWY
ThpwJHKfI25szlOyMaMBdk3EYRHuHziWrVp10MIEGM+os/YnyvjaEgIvx+rCDEvI
NHWJxkXW1WLPeoctB+GahhBBDVpBa83weZdznFtw8ssKHVljFYjHJNQrHmMfUVl7
9qeSe3yXyLZ8XfVWhLI9dMJtyYrEVXU/4j+sqHGUD0v+zF7nber7mreI2o98NRLJ
6pYLiqXzh3OGgPaS4Jf15Me049KxNd+yW8DnNbjV5kxTXPs5ATJNf+oV0ZoZnYc3
7hqHuewz0LLiijAtD7k2xZjtbcEfWJRxpHxNOkdQ6hiNeTj1ZllnPMPIB9XbfqE6
3vrxR6gIQnyCpfNHUp6+oPKWEknrWoJF4PDCZJKjxui4B6aPXBy3iGymYi2EOnQ8
cUbps6IZB69ULirDFErq/RcaZ5mqoJvH211LJPLbVn9uQj6TMtYHCLrHJwgCMaa0
VZI2ZegBm0e98PuqnvK+AExZvDd7C1HWzQiUBRidgOXkkRPXejT3UhY9VE8LC4BY
LnoI/SIDS1DVYQZwTdnaKjp+vxEzwkIFgqQfyeeYs27Q5LdM0/GhIDO+gbyRMTnf
9djz4kXchoWja3CuUc5Wg6lqA5tVqncgg0V9JdOOaBSlJrgVRxK1zsPW73P8hDcE
8Uyzevi9O5nX1tz19CxDub1z9JCN8zok9eJSczDcTkeeqE/lovlFfA+NtY9/B+5y
+5Zk+l2ciBr/79tE7fhbOXkRg2Vb7p1u1oImCeqkYU5AudZApCWOTQLnOQW3Sjxd
K+zrOM/9+l0knZpjA4qyqDHZ7oe9BrHUhOe3iJxRrYyW7SuE62SZmdxBjw1AcM8B
Crxoqb1daMuLrWvRGuN98rdaxTBxtIA0oIZOxjS9aQGzTBzRm3dBe8TaV0Ky66XT
zBgHmcjieti45aenLHHIZKwbXxTn4Iv/vt0vj3/lKAG/1cXcnPxdx+xSdH1oFEoB
4N88z5DVKGN/0RwkCDoQ7Oc8Bu3i7CK1W4esmuQodTsMy37CwgeIdMGIqKZMensk
5SAy+mioXFKEqlarOzoGdqIEMxADFqHwMeE3KauYSKplUFl0LfaaXgRD1FFtwrtn
oCjuJ6Ngbdm4IgQ1khNyBkkZo9i6jnsz+sMGp0VeA7MTFc8yD+53c/pQF3qzn295
S6GfP6Htek4T8eaE0pxXkFLchHp85njCqauMumTwPaQiisMw1OQQ2d06x3aRLTzw
9qx72uMOH43KZ411R+Iv1kQolpYrmsSTF9Z6jsHotLP6R7LpFNzCnzbkvVa+8uu8
umvhv+2lPUiiQOuYYOtLIgIHUkZ2RPquRBeGyg4bhY12mggxQpV9Z1Iyq4zW7aRL
id39lTZ1Ahh9B4/DER3qeL36qpHnf4RcVqFdD/6HfwBYLWuvudtnFRCFKQ41qxPB
weRhLyQGVtLFTaMWoWdPTp6vGpZbIENKaoNZhEWMNRmmwyKUlF/cElX0RLhPJ/mS
evrL7ZOwO77xvnSeQmB4k0m//9y0RnVO451GFMxJkOjL4pWXY4GQdrItzcgb47bh
lWNKg9lnKG9bAAXdV//RRsnzEsezzf/I95G2iUpEgruyMbBOtj3svsFm/T52gcHo
6/43cUYf1oX9BHwMkMFopqWyjFjea0xG3dCL4ERZDC47xfelGsMIv/Y9OeqhJB4p
vtfDtINn42fq/kGumu2Z0/I1zzwsjhOhZcJ5wGcclCgNgnsC2brfObksCJ6chteX
8wc+56Ci6pGrQsyY+3w3Owh2slUQaIjEI1njq8WroSwZCgEXOHaQ9LuzcDfDb87n
V3HzoIEx3htUhfkQoxewiVLEWqmrpcrgohfxuOpY7KEOXv1edabD4gHvlquKt4qS
T5rtQsFwnxxcORwr4hV/vcsJD4kTojFVftYd5dn9pD/ZE3ObKvrjIRz1BkMp4/hV
Pd9K30/1BgPTHDY/KZeyDrjk+GX1LQfgHIg+xUyRQ9F7dfkJhLfV6s/phaeWN3gS
Y72gcxhVGB3etqAEiRrjvB8FX+NEQqRvHcEFZBCszt+WA6EN03g59kEESXFSgM7t
tdrYV7xujDrJ1nSHrXhPGPzsiUjyB3b7UsQAPBN+DZs+46DdpNyP3nPQAaYg5ECX
a9xDvUMiex3RpPNsbrbmsYnPFnysVT7D08STHVXBlpxQoNC727xt9PisC+Ow2mFg
TUSGvxGbtD/3Xu5ahLB0BwHHAWP7i5wcJxjPjt693M7cfq/y4Q8B04rsE9N0yzC6
saI/nt6wzh+fBsRJc8JXcG/dS85YIwozmnkO2QjssTtUiX3/hhayErwVWsLyZp1r
2ryi/lBizpPUpph1SNnTmMuxgJ4KUR0G9HWz2MOyErwcetkFAQ7JLQYIKAzG5Sfa
yCUuSaji8em2B05LMm4DP8113ciF81JTBmr+GbqXJxNefD+1vkic2Z5SRn4hzMpC
u1FbujreWNurV0yLekX/ZCKCLgAo9J290J4ypzhOfwTxiL5eGIDFJo98zO/Ud60r
iLoRaIsefLahfz+YxYnQSSx3EVZaF/etqW6BSbpt6QMcoSLOWgci+Us7/SElfiDD
u2JmkzJUIXO0WkaXwzaDIhQvT21P7i/Cw8C3TQ4HQeWjpgYAIjFL8y2ZmhONSEnW
E1I7VSG2+4JbeIOnfT9p9GvogOkIdC2ozrvlf0U2WsDXB/OlSXqG9pJyuYByzU8f
ebDjU60apH2VEZ+BBGSMeAO9QdJ983oKAsnjhkoeJz4MP+jU9EsSy/TkiDIKad+8
GW8IEmv9vtAAYMob1RNaJk2vxgLD7pbnS+0+x7saRiX/0U7Y4/Xzj66ijFoxayNZ
P1YifOYMCgxupSfXanV7rNCp+0HsXphgq6Lzqbiqj2m15DeTlW1lvqaZs+d5vn5t
wQWlmw7EWhZg50NsiRM6S5XQy5FeQWB1oKlZzTtatDQO5pzz3Fv+qPddZ2NdYi56
gT+rwTmB6JQQ4rKV6599Txesn54s8Y2UiCnlDW7VNhoVGj026QRpvXLle3R/EY9+
/Jq9L4k3sbcFlEw30CoVizxEI2uMtQcV9fKM+0WBN/I6CUhBUIITbF3cjoupZgxD
12m13z4p0wLiqx/mvUopR38RYwJpK597b0Yw3UQex4owoIbhMQoHvUQMvWHJRZrj
c6eDu5goZ0XKyc3FIDz53hoUEpQBvCYf9ej2zz79/blm7Fe/Q1xGxya85tmbCLtI
5UsDIKLCFz6FyiC1bB53IrXD4Q5PjHPMT5yJ0ev+iktADOKOyKjGduE7BrC7mRjS
GFd6T6r0cbozM0ALioAk6w4N8tTV7eCEGMHePlZvlDLwNd194ibKtSGDjXcFDdHS
wK6xN0pS/Yp2rO13CFSgvehHZ3QHNAoiF+pufZIj6ocKUuIB8NjfQd+WszdajdSY
npLeesk9zkMPJPrISuu2MomHhGgS+sU3kvAJNfMqsm4dskcW8gnno86jjsD4D0eE
YbXy29aUM9JK0V4PXroIC0nChbrcaWZUehktqJU0Q8nePerLMy8ZyFoINXumabEG
6VeghxZrml5kheSBfzbU97MY98rBCdpvbdXSurXtwuz8B+7g1xbfnjtu1VfqlG8p
hWmb5jCRVqX30r9a7CDRsCq8h/l41O4sGEcjO8I45PiD8lY7mQZ3YTMFTE1q9gZ2
O8H+M49PSUErLD/7sEMnclhTjierzdrBuapHCNPFKjHb94anUOAMbtp0be1YL/Zh
NwegsY5xmZLYMw4Gh237dvrtF0ELBLq41YpT1CFbJ2xiGx8y9Rny1UDlTb4+y3wW
+o8NLmTCPnAH9zelfsxXpNUo/7qTEmvnZ7AsV+SFLxEMsSw/Zsz2nUp0LHuxn920
Q/d5zejdooPvt8JyMpdi7dzIw7vi0ZVmptZCewtMQoCjddVgP/gCVfY4ZAUyBdKx
q7RjWsXpi2sA2XecALfbdIdPSQBJGCAa/HzK/WQ6VzH7/JqcMQD6PEeNnKWPgJj2
lA/NtUxH6e9d3L+14DMP+qZeVfPOQqEa9C/ha5AF1bhcPgfCpIGEcjcl3m8WQNqK
mCc7uJyzAVcumxMy4IbC0PPnrdDP5uRaHa7LIj+ylSa9j2MALVIv4w7RNRCuJoGN
9x/acIf7MXmUVGpkH85b0f0DE5CoYOlW2CYBLOLEArWRXBu+x8Kvugj3zRcdGhap
JwE4+gqr3TSDPpQAifvH7s/Wv38y1UinTS3sHvHSXxxta72t/L3mXNOwny4RpZFg
UbHLfVXhILkSOjllCBbXWTWuqUX/D4g4vGUSO8Bxc8rvE4EdslNtpMc1xDCVqXSi
kVew4ocC4BhcUJqCOSgnrSmXlmQ/lmzIUTNY+4osxG9Dn75qvqY3n0anCRIubiva
uk6Oe1GJ9igISyHAO6CY+HFl8iTBIwWMUsqEGI07oOf+DAZ6irIhFqld12BXMCY0
/3sEYVa13gHf2zfdipraSbsASJS5+1vbG8d7b5nHffo6qhAi+t++51ES0Ld7O1Ol
57FS7rzuMXMtXCWSiSsTYSnNdnUdfkqpcl/otFHJbbhng2Ycr3+rsOm8g9616GkZ
FtQSLU/QM4TUQuwhzXlWz+E8lbBqey0RrqWyow/e2ldZbk9KnHaM+hITz0Ex+lau
QBZP67e7HIQmhwTN7BqaQahUIeZEdh1XNV1CZ0HpTmAISMXTC3/Ewd4g3E6AwkMp
cMHPomuVlIjYFbzHcsU/5SzQ1hBO6ls20anysma3I4BMGTP9ma3lHca3CF8AsATy
dzp8rVv0wgZLbj6bQbX6GfnbMq+eYX1c3q69MLYfaEN6/Ou3OcNaBUvm2E57L5sS
aybzKDZi/getLqkf3bUJhdk5DLb0Gwyb1ZIr065v/nVPyuc3IVVjJGsWM18+/I/w
0ZEGuPd99nzln6GQJ9pmvvr6pfO1rm2RJVo601DXHqPouVXj/KDN37FAtjQwMuUs
5wly7IsVPFqphMEvyz3KfTi5UZQUn6A2t5VgiRtmwfrFxd0rBRuPKlWluI0H9E4I
ZalySdGFcGVniYPxeU+6riMpcDsf5ZOH3ZmW5COWh1neToobpcjx8MZCKWwDmEU7
rLkMwO3V7mUGJsCxU+8PZJfeWoyPSyyjVzOjamOT97F2eJdHtwnzhiEhfrZz/mfN
w8Wok/ZlXtQwEkOOuSW/rtMwrKWmQPkUx6bwGZUXMuWOtfSaEB6IlDhStxNsGAsb
df3lXwA5j9pedh+1SU7U0+vZGat73TyKcw5mSwr/O5xNWpBtPjzvlesu7o1IeO8F
ceIDaVE7/gcK2wX8Pd9rKUUCKnzc3p57u/0PZAf9TrNhXz6dX936DRIpgHGOILY8
CdaSQQq6w8McDLT46xOLXXQm9ck42cvXyIyyuWfO5WzmGOuy4ZTIdbY7gOid9FTP
YVeEKjwfA3Ge0SaFRUUVhR9yETjxydru7pVFI+5rEfXXixN4KvqgMCCdp66fZbao
SuE0EF9XoDVQaLfsEANe4SbJs7TzbM48P/ZL33ODnRLdRleUd21RjXOSZrJAge91
oaGU5jC+66jg6R+jgJ/MJpdv6Hwstkr0ET6KA/JXlZ9k8foVh31Yx725WWnw7Q7g
BmKxFO9ffw2pHj0tdURTZwmQZPzwSoVMTToBuIqE+NT6fF4zYTfY8sz60njU8vMr
EWyJUm7JpZnAJ2RLjlGaE0VWqqWXnK4WnD+q4p4kXJLxiVzT09nYk2x32wyrZ178
dcwIOotnJZHMiWi82Z0m73nmJo0I2/ESur+l+RtFm2DFSgTIBjnrpxxkyJsIKfhE
+pV8i/2yDQNLwgcHdqxEfZq+Stth5CXrop49jFcPkl5R55pZa+OoF+FY3ZPkt2cU
ReaHXjzik58Qksnu7EqpMCEmjrK5YZvCpc5NLJuq0BQUAFiGqWJkj3QdspN99fok
2dV7gbmQIVEw6TyAwmqR6bc7wd1uP3cPXHENzYb2LmGwxvIhQyHODVlR2wkSzpWo
NLoQm6e242hwMpVXZpglgUojDCj8a956axIcLjNMnM6ruT/Z7W0KeXB9k9i2dZYA
PD0S9d84lqib89mFNnafSVD4LIJJpCQm/AVs1WI3kRCDOAiaC0KmO89b38nVHLtM
Usq6uIeJZ1oJf46hZNXvgrxTbOdkSU1OEdqO6CEgwxzjp4CWdw+JCOnjKjboIsWk
p+SF9qtz8ksoqcEoFEY3wdWedb95BerixD2rU13lqAaZWH3aOmyXJcbIj6vmhMP0
vYXAK5T8pnpl7uIt3cqg44qYhfsUwrPercCt/O0nznYEEGyP62hVPRy+f6tQhvD6
y8LjEwOUHlRuEJLcq87YeHuV2WBT9rPtYsjy2sP5lx6No9+MP+F9jVA/ydYeu0ml
WF1oNbP5BDSDjYcneriw5mNAiiV6JOWINmt3yzHOBiHD/gAOXjN4aQwuxpzAxL+1
/uPqREbt1JVNhrDVJxCDt4DqZAQQ53q/hjllF/T6Fuo6tcjGVu9MoBoUiGb0en5t
Y8VqBJVgSh+njgVO6S1kQpsV2zkQodbf6nx8cJ+8xarEvmZbZMcWwB+nKlj0lvea
rw7l/8dT5IpDVb8NnbDdBEfOzgzKA3RDjLrGEs3+u5pWLKmQdvTBapCMb3CISdwb
OKw/xotiVJyXx3cQdQcGsNccRhB4S+07eKiZN7yB73z26EL2kCAEpqMkVXfsFGFn
9T9m+94d4kLmdemgoLVWX6JVxf9GdtgcSmJrEBvS+FFI1SE0nXMNQzwZBDwSzH4q
SQvy87qOe1W2nLaAHc2CJuKd3xgyxhqdNrX3kz3I1/6WusNIF/EAPvNwnxN3qM1m
BDf9UZ0DbCMRZzd6w/mnIAgMtIRwypH0ie8oWzB6oNlOKnNSEix3TgIW3XbizeXv
Dqsrl2IW0QbMZIOUauaJ4pw7UsNWe8HC5GcqnbbxzYkmybW9ZMfnZEYDUF8pnouf
YF+n8zJRITLp1DD68Dtulm+56F24WyoQ7fJXRd62fSlwPKupO7LaePoFrSCORXJ7
VqX9aTsoHNPgPLxrUhRa7fZIexNatLFzr3VIsvpIjENCsSg0gK4IyNIqT85nIp4Q
SFYZ3uZUeicpQk3eaEeKiY28EWvxqgHKewMyndEHcu8q7KGsrD6plaHCdlxNxycv
mZIBs+jzp6rytwNzkdiRtzzGb4iYbOHlJOtCZKJVuGovSGM7TXmouZxv/dImUMYt
LfB4E2tCIPY7XREof2Tz6qEx0/IZJwzmi6vkpaeLqG8XQK8SgdXd1DqX+ludgyy2
oMKiiU6OF2ErmUqZ+AT4wQRFdQGCTNR3bWp9nSPRaHqHO3Rpj1bO80Fw5+/eSs1f
mhQKttgDwtn5AhMVgOh0PnyvJqO1Cx+t1N4sh5NQGaJJ92RYgit75vlndaJz5eEi
gURnJBWEq1InlTwoqAZl0YQxObzmPinjSeucvnm2t/2Vn++BF7EyjU4FmWEpWMlP
OvzvbJn+Rcoa+eDnK1RN5DhtwTwYvq8jzspPa+EOK8g9pKcCmsR1oAqFA5R8BQQg
WKUr1Qj4jeudbsk5NgBUHRiD7IvVq2l+yamYcX0jIYiEyD3mbq0yCxasYRlyzPwX
TnaorNP7QHwkgWvyzQTvwNOLr0e7CViewfdjxL91oCKNDvfE4G04SHXawVym1yTk
vWr8S7XKdO+qXksaIyIe0V+thR0bi7nrgnCjy5R5ORCCYMop05VF8/rc1mYYHkv+
eF/MiZ5tq6h6xLuUkzkBiFnFVqVtXcX10eB0z+n6taUE92UX9bNjI41KUk3ZXtkN
b0+mcDcLmLDiID4whO9Us3xvYU4eFje9evzfstPU2xIeRRficNuNFKJcXJXz3bxJ
0dphC3HIJhsGCkx/Ra2FVrAzgNDjf2NX5500lChedOFdiGcg20KBMsHu+BVLyqiB
BA7QH42tFHSGPgLz/ay2zS2deUqfgCQrpldDrFUa4VZptEW4WSHDaLcxdc4M4PeO
jsLGO/i0Sg0FgvzGg3bAudybruFUIgJB456gevWSCs9XJFtb82qnkkdOAVDb1vIk
/OnLTpKil6WZlO/ROeCyTZ8qfxCizQHPDqewATsW8OfFKUZTfO/etOps0LrZE/iT
pfgiwx/UYgXRFXQVL5BwWi0HAd9rVwXy3lIVrSB8yNkNCV7TrBO+mfP72hnmvAO/
miYcrwmsdXD92Wy8WFCMUNaDCTAOBWXPDU6Y/fQhDgFFF+iDcqY4q9XG+excj4YT
yf7gCAyUmMeRXZvA/2I76d8z13TE2ICqYz7q0L3adEqe85giPjcPk33hRhLN84YX
ERsEUN1nLxrqMwsJwTAhmjD7VpwRjCuiyafCCu0e+AKlRALGf7VRBUpCZR2Ww9zP
8J3n9lGHxWhnMx2Ld5BdRnAF626t/DmdN89RgeoElc9snJQhaQROBuvqO+1bc/FU
+hKh+2P+eOzzO6kbUzTMRle1xGviApiOtrUGX5R+cwSHCX2Y4ob68GM/h/wYnKPY
SraYr0/wd6gXc2fmesK1aja9Z3VzmPwsRpohSwgiKtnRXYThF5P0IsUvaSUWMZWH
VkHlC94nPFn1K+dAXmFnO346LnC0zkFeGUrZcxErDQSfWY/CndDL2dzU9iuViVCG
TXwCvFH+zDPc5ftmqt/zj8qN0Mf0Z+gHAy517K3JnTWgWQEqST+RIlD36rMM1uuR
h7j+RMz+NSyzTLFHz8z+UWY9J3ceeUm8ZISalmDiMZ3bK/b9x+qyspRg6jGs7vpA
/TwnLmf4Tv76fqv/PzabpiCekJ7XZTXOXa681oHZJnZhEpIIjbqsxLHFQpwNFl+X
7HHqmjyVoz1erSyylGRQiaJQzQIzdHcmZdyqwmyQ8yfBuO6HdsPj+iC16K/e1S2x
VL5kw2xQY0SdLERic2D+HhZyPPGD+p3gmGdqagWkwH8N+Ew3qkGkjRohzIVuNOkV
y/mXa+dGtkj1zLfgC/3ail4gbeg8dGAu0QMBnYB1KZ5rZdadcxzOEhkebQL4T2Ga
RJyzTqwsh0uzcv+pO7OKAc6kAkvOHwSXpBwRZfk+P/PqW6Q6XO3SGxKKkW7GTckq
7KNthClJMqU7o7/K1BH2BcmLzDWVOoxsmRmoSBg0yCjmIj/LOR0Nc8sMYDJ9p+7F
464t8bWtuDPUt42EjCLfAy6UsxJ1aTgMZX68SdVlFYi2MzUo//pESuQIgjn+hguU
Vu6Jk68i/5X+RJihEZQn6TsBT01iBWiqLb25hpfHCsFEyEPfTRAMlqukvlq3NIol
+QvltFzc7hg3Dd9/S5oSfpEf6CFNp74kd64cQBhG2set7BXVCNs95OLp73hmHdjy
hDxA5kgSOHMHKb+bAEOgYGA5XfivIlhNnqCmGExqP5gINAVQfzTfL7XePOqxITVx
bOzquiktEmMsAv+J1HhysyKhB5/gaIQf+5M/G4vLLWJQmYkyrEpMhMYeVpU/psYV
iF+JIYGNUO3edrTW9dU0AyoiIvJRTLEraqv8hilrM3irqy3bquLxK8puBkl0uzyN
Hcs3UCyRtvwVTxBaqCOiQ1JI8mPsLcePJzc+5SuR5HsczczU5nQE+XFPpIwh3GVE
TOO7KbQVaJJMILplymbNG46P9tuTedackDpps74LYWj/ThjzGd6rNss0I8o/Dcs+
jJDQyY+SENnt3cOlm5Huz6AKO82cbum9IBmP5uVAu9a71rQxKcqEcjcunz4Rk7x7
QMl4cU/qbxx1pz/8hwRcCyjUlsK3pefODsvayDyWE2nLdLqOu9ux3pkcZ9LBsyja
j1RJ0J+9/hsV8D0hIpu3fyejeqvnmTAxBY6QSQOlMHyHoiI6MWZ14dxwRGKGSbi5
S25XuBDFIp3YnvsWkNvYG/P/PlH3mQHDOtBEpmBjHy90b5OmmcgeVP9cgpxKOv+E
qVJKS6ipLMe2cT4hy8qx/OGAvymkw73cEkUhvRiUlNg0OaPdmu3WfSq21YsvS0ZP
QPRbcDn7wWsU7CLojTrEyb+H3MSSa62sZEv0UyhQ4lh9tdF2Wg40lBmB8fBgQV4b
dYAafif9P3hJ8NOGb0PxmzLf8UBuuWxAKk2VtbVrRbG/8gYi5WT3CcW9XmCRRC0W
ElWBZQRrNp5A/Trf4f/d6zKFQi3XRBfYlzsAyRrP8i7Q/zjbm4je3FAKqmZzZnJu
2ngUXcek5o1G9y/6hXkYEzKcrGjaafPc7uFM0lzznN+qIf6baS2QSqVNb/v9h/FL
mjPNq0KTYk6WVfSYwNaMUmeB67QCZlhDi2uVtQNCCxselMmjYoJIdII0yNdhV0U3
CgYNTeUoWZjAmmYJboqyxbfuMGYllMbxTkyLfdufc5zixdq6OKbRyzOEx88bAsSs
WsT1gJVsuI/QitD+Kjq+bX62VwCgcUhuOjx46ItPjfpJYU69iGamTPZ5OWbCOysW
Liiu8BjNR1QGJzcD0yUMGD96S0tew0j6K6/9E54UxfBG1/JtcY8uHEiT9miXokDn
L3Y1gWcuXVYdIDr5rdyNisw1Uyp4A0PYaJGraYy+/22O6PLbCXZ3lWChF0vzDjAb
PX5pJXIdoruIr0mftrdamJpIOssi/A0IgE4jclNu01Io31fM13hSdI3pkl3cZ7Jg
cC/QKJYbWRx3dLKdCBZJtUceUzFSHH0P1ZFuE+BSIzz3RUpMrXagz/osvCkfEzy/
XmcH0DjNXB1CrbIKCNsdkZHenW0SQeSGAhqvfFkBv0NqeRMDVTowDuhRFmqwCmff
qd46Bx/5jVIXzee8Mf+dosdqKkFatX3kkPMMLZPy1f3hn7QcD4zM8Fz3Ayz7bffo
w4zLfF+Ks3nXCBu0UJV0A5Imk1BQcAeCZRDD7XnxN41TjRTkpPvaZVodQdI/tOXd
45NtDvW3MEx5eCN7o5K2rItonLRX6ELNpE/DcZL3/4GjOWjB5JDxdu7h9stgz3bJ
LaoylCUIHgYpbXpQfPw9GzH+vIZljT5dBD827C0mwX/cSa8ziH7LxaxSVhxrOmPZ
D0DxXee8VsL/Nx0vMJrXyhdhC6nmP6ngnnZzT4l2q/tXkJyk14BhPoqUTmmR7TKz
37HISstAuq/A0ftInkGkXH7tWTFAgyR1Lw4WnDaopMxS2+EGvmks0ZVKTGSJISCe
eO/l7xLJ0PRzG82t3SxB4dEX6NUFwrWzS7Yd17BPYo+VCK3VeXY2rUhfdUgiiHYF
X8c/Pz8FJkfe4qQ3aBLSW7z2JAhE1YoSvmU2zqsHRc8kTZ8r522C2h2aVBQwhKIr
8pkdJagEG3V/jpDbEshEXJu2r0YZGJBTefCj4lmsTy6FpIsY/YQvPo6z67MQvF7i
UhOrSBV2xmBZ2MHJ1Q+L1VRLHnnXs+k3kTyVpaDyGgL3S0GyedR11XKMkW57FawL
r204C+1UGj20PfFvduW0rlmjCmu4autYVgsRGhWuKjrBBNkml67IymrAaTvwRo4b
Xu4PgSk9Sq7kGndURr7DsiRn2qL8ZHz0wluK/Bbw+3q448U4II2XDgEJ9ACyImze
SafvvnmoI6nHlvF/QhgWdBff1BVk+JFWKgHJ6oxJnC+bXaEqPSqnkn/U433J4SCU
/sqYkSNeXcI7b52e3sXsDodHwQG7cJ1TiSl+1pAHzckJAyngNsNyfnyACbHsMh/x
1oI/B59HNemmnGsOPaEqvTHGt2h82ApkdOn8961X2gjSaYPFduyUPTsf0J8YF9eS
V9Ga2JATKq5TF6GG/EfptskdjjiQOmrKz1Lz0+/soKu3ArYAuMya4G3pSAkouB9s
LUJO/fV9RUarh/MsvsjiejnsstVW9EJ1ZujCc9VVG0ypkK/W/br96ei0fKYxtJlc
mQeDOa7Xh1ItxZYSRc3i89w3GtBnARiJ2zK1sNViSSDLuD5vsu8Fp23FGAftu8cj
1KyTmSa/rJZNfa6QNnuJH4c9UqYyZkNFQANuOx6HGqnA3LD+dUA8nSP0CIFmC0I2
6BK1q2QTn2CdFKgX3tS0eea1y5+OjxVQNRJPlCtYjW9llzFPOydlRtZ5EuxZjYKE
Zm+x/TIF1NKolIA4R9259WqGR77Sb0eL+E/vW7XPV8HeaToYnFkDovtHI9WK48Zs
xRcQMuykop5tpMfzR/pEsv/OLle1z27vMUpjIszSsgez4iWS92f1uWopSKRKRA6e
hA029eAAncMLc+LJTq70SdjizqbdTMhP1fzT+yR5WFSaE/fREh1TXXqO6N1GBOkK
Umg1MgBfpv/0D6CrGNrALnDr2m/u0I7CCTvrc+K0B9q+4/mWei+S9Cw+VaW+IrlA
7cnUBK9aqqBMMX33z3w7Dn0SE5LQ3HpKQvIOP2yjKrjMC+QB9D6ifcc3EwoAaSuP
+0INquCSn8sE3Awlqx4cmbYvr33ReUmx++J6WlfQ2CTtGeE+rQIgmPzEz2DhJNU0
zlgJ6YbVqWx2tDz9LTZgmUqWUn2uGYo/7tVKDINxpickftOiEd4OGqtKjRm0Z5Lv
aH/RbZBABRqmQ4Zuy8+XQ7q4Azf9E8puk1if3BB0IneWf1kXdnLckiUVaMsGYWf1
MOucwvFQ/Az7rMnthy4FuJc7zFCk0fmGkjZRlxg3PWCbnU+hWbITH3brrlK/8egW
wBzPdFoRx0AXUKH/vgioIHjZPUnN6Qx/FK83egH/av7lIlWbVh0FJmWTohTJkTtG
Ow3ZhI0l/Gt8FX37l/yRY/3KhHMFPKhFri9jy49KrpDvksf8aWzzQoZQNQjK9R/Y
rVTv+rr2siPz8FEKFXrwPH0MVpIrHkNgPZcAgKlq/2V1BFI6aAJAlSP0yMwruOoM
z9bwGUdQwWISqsSh1tQEvi7mh6sd2mIWxWh0C/5vvGSi4rQmf9dFKTXgyxR1INpd
xoizOOiZEL+dcbHYuMIlzDmzreI7tUiFZemiqxB7Vm3Fb2ydolfka/rgcK5OYwOn
MPV6W3DeOZQsqcnUqafxCdN7sxytY7zASSW8fG20f9c0lMMiKh8nYPKm1aP3UM3/
9inJLLe8r8VSYg/gVBdQ9CbOO26ViJvz3vBTndhNTOTtFAt5zuGbBuIRZeKd9wQw
oNL47MgIWJ/QgFmGEkHsDJjPg+ArZJqLGUiq+lYaiGvij1MiitRCnHVCHmLxd/M6
s6VFF+XLMhwav5SM1HCbpKqspOTewtQxNDix27L1bFSOEBZyv7DqcPRlUCJNtB3o
dXV7wuggY0sHLTA524ElcnNDN9Nk5bDql6J69cPhYCXqXvmyFvwYFP95D3zlEgYA
xQpIAmBtVyIg0iWGARoKJg9FwNxeUsU2J7imYaPjxWRVI4Z/J+2Jlj+UpW+mrndw
9xPmizUdZi8prWLNQCLdNkQZCGkp13feTvJH7Kegc1piilTssw8hFi2acu+trJdE
Rme8oW8mMk1uZCeB05WFdbhRwoYkzsRb73z0g1mOQ7VkOg/wyovnv64FouCKTjqP
bNzj3Xow22KPm1FgzFVO1BiIfEcvrIzi/6qSIZQG0zVCCzQsjiJfdFfBptLksBbJ
KqbMc404cZbUQ/K6elbHEiSXte3UAtIpg4Pimma/VORg7xKpuUO8dk3uO81G38ey
Enrx4X03LqTS0sVUSClzb4qIDUOmDdGZgfrSwTt9t6S/KuS37zyu/xdHggGxtmvZ
SfjitfHgcgS591BxAnlsnKQ44uYpBBBRuGYIj5G3n13cAULLviwY/MQ8VFGy0z8N
aKCevtqS6DvykR8yXbMSG4lb6Er+HdBkgbl1lxunqcIHRyrMHFZ4yDE6XDdvC6Ft
iwopfKChJDQgXRPu3IER/GaYUxdHbm/D/XTEmnTPjtJkXTPLeJyaviN8LBVLOIC7
GkCJHDbNFjpE9JNxYfq3nSdlZZK/YPGFFeb7AC9L768ZHq0BZTLH4Wt0YTQOlBxL
MEhoSDs33YDkZ7zpOonLvGYlVOOcjclKE/duyyqncD04h4wHh2sZjK/d0WB86whg
Vv3+dSLyOSm82iMST9MLFpG8C0tYxcvEPVEjirOFVwHR6UgZX0gJfoxAy1CBDL5G
MycFVomTH+mVLDBfm534m2mE0FEFltprkjbGruQsI2YeoAr4nEDES7o489ChZ3XO
xuqgHEfQe8MUdJz5vfFjJaV/sXsYJxv6VYOk52A9fQWWbrwn5gcDBd+TfH4JbzTB
1yLb6kmxJQeAmgW4mn6SL/h8+ScAjN4XI3ho2ZhRmyHgJcLcHYAcdV77VO9mgQPD
ZL8zAXHrUUU1gv3tKhgH5nErfBEeO6HXNkQpdj3wKdnxedO3Yi0Iz5lhS2Su+pvI
05+zONHr0ftwHVXUiIIvU6Sf7Ru0OvVd6QO1fKHs4TyFXG4BdwK9NWXgwfmmLKJl
cZ6vDqnW9nHUgexxhFQKwGQu/giOBR30nJ8YCzUz2ukyTWG0vvXj9n/3a7ahvbGR
gNrcr0+04CEXRC0UrazKX7D3HwBx2/ZQcffkq+CpVyjHAqYAKfiAziBgVjveF00a
QBOKASA4ynV3q3BABoj1/2qBcFrO8i5V6oNwjoM92ZAejKniir+4ah3p2iSGoz5I
Lw7sHJ9ylBTMKiNika0/J62kBMJAfHB9s/k9nr3DNtIKOOTlNYNB9+c8sJCWouII
jJaw9Hk8jLZ5QPPFXLItw2Qu9fIB8chMLeh+jFQBCFPJsKZ8bzDRrcZwHDuELDpU
K7mlrLSGkCuto3i4gPlFbiDj2sIbkQc5J3AdPFCOkAG47IQRAtbrS5OjCwOiX74n
uNxm+nyCtSGdz1BIkaGHogs8/X5wV/NRvQHHIDmC6+xLxX4EJwSd5lhF2kmbCOZB
TOUKke3x0ZFWqqHO6O4/9ujmE5ZLPrHpgVZoga4zkyeu/3aciurIp2soKjCfNY9V
ExUuW/6ycKWylHtAfBtUd0rfLX8J39u0Y5YvrD6u1waIVrBZfqKV4ifzn9MdhUt9
CReeP2UxaYCudz2WTcTapX2191RMfB30DeVYBa2yGBErMvK/hchzhfe+jR3hffdW
EiJCv3pFEEWn15wJlyFeQt3/Tg4davykw7ymUPkWRWkRPQiDHGLH/6fL4LWvBhHP
J54dFbQsh+HbN3D+boa9kpfJmMAbp7NijOhPDR2EF3R6AbrHRicvUzmqlyFyHgJn
b1Qlxtk/L5OT0m2kNwcmEW+S6hl2s1zXfLatUmjJDWL2Qj161AJjWMdUHs03w1fw
DiN0UxXfgEsnJ0J2XVZ+JBNBlmX7cfsb71OQBJ26UvPC9ZKKJ5U9sgWGzUSjUeT5
FX1M/E1D612eisbAoOkYxxvYdNuPVcs1aKBom93uONVSq5e/9d+34l99488US9t3
snU96zrFotIdFmF++F/r+J4qnLMfZ2Xr25S7QAUfjGUUQOUaB1uQeINnl3yeReCZ
HeB3C03ddsJStJhxlUlZmsj6QwJ3vqavh8clch9t5oXneCjHPL8gzo8Pvfr2uQYC
1fNdiDM87eE9HdW8Gi8204/YuI4tzH3vD4wRMuHWrEFnTTvjalV/YuDm88Z6N6T0
zCqYbewCxEBB8PBTW+ueFhH8ZstOsARGJbhZJjhMyLbX6x91ElvGkXC3D9iWIU26
B3kOKJFyoxm6ONI9JPn9qwR4z4casqsTcKEEy9iXnLBy/+HSiFYYcDfZGiKeeUGt
bMhBaDwuv0Az17K7R9YpQx9214U+N6256ljWECRZZxNJyqPBwFql+P/VgPjqG0vI
RemnkK3XARX9YmP5GdrIHUF9bo1/RIxzD5EmLEJBiwDdb93l0+TaOwdnCmyHci1u
VqLAKIvx/3jDm3JCdbx7hdIm/a7KSUH7d6ppjoFMQM+tOMJ//J/LykgX4++B57je
qvAlIVhyvt2gN3sI5Fuc5JZLEh/ShTTmcX7s7FPcHFzFCgwn9ZUYqDDzs/uKZeae
nnfN83Mx2dFVQ05iUlO1Qk/eIJWOriTT3FvopOifH4Q5803Oh+wukG90n6lCLeYS
aD+eEfcTSxdQU1P3iVYu3kjGsd57olqRJU3KrojDfXqmsYEp0Dg26ZYAxTrVDvqs
jS8lRX+5ji7tIMXe1jW5FyYCFg8MAK9ng5ZnQ+MWXKv1N3PmWp8PvR8vtFn3aSkY
hhzH3MY5+SxLn2vPb9QyomTq/bF1+PCl73rR2FXaNHf9OT8DrzRKp/PHcGK7Zi9u
/3ev/v91+pHh9kE7WV2hooz7jgJmx+eb9988/idCVQv7ZmmeaLhdRCiln+qeOOa7
7dIaALbmGD3FWkxbXbMu6Pz+LbQFDRY9zS1Varz0gqS9PMpjvAjjZjVj+pcX6JdB
jvc5ooWQmznD1BK7B7JvtSxaNclqZnSqPeM2ZwszoslTu6cRU07ox86UQ11RgquK
K9goNFC0LL/QnvD9998tcEmBYt2Zwvn1Fa8LwSFm9Kz04vDSMbQwcPknde/y5g8a
D7zLQm0Sz+quGU2FvJ3Q8RBGoblQyDvCdWxs0kkGvWy/SDSaN2QD+B+ey/4nbWsS
0TK4dmTqJvLEV1PQuSp3g5XEPLYF6cUpx8r5+WavSm5bPxkbsHf5PgtOvqz3JD6E
02d8OMOph2GpprSyzOOcMeKsyxjPkRlXsN+EkoeVnY1+g2VGt8fffrOHJRRaQ4J1
BlN5m8bHF4x70/6Y2Sn+dy1ov1eixiN8Q5fSgoQMu3pnXCr/76kaCx2IHqD1LBjg
W6jibDzqlzGj9lBrKUevWPvXUcO6UVtM7N3eDt3tFcDKlSxY8dyueScO/ZTe8nmZ
8B5UFXGi/mIi1CbqIf9r2uoH2IyaBXl05cprmXOFiVRxyU1NjkCY6FRlJF2T3kmj
XwTD31ynd9Ko9ry85DuK7YP7sugGt7pzSIsjnmOTLpAfHnYA+UH1FNVe0dVoMNg0
5vJISiwUfFE1pLNiFw1i8ahMZxAbZu1DwM5LxwFbdE68F5vAfSHgdm74uw+Ib+aP
cVbwmeO3YGbPTI7qexZisRphjQ0GsHfh/aSgeLRyN1vchzTNePEyGtJDBCdneUNl
j0nQHhuWr/R4h3qTjv1R2iZnTPjCYAntfuQ8O5aJHHLBJiBoNqOaO6Rsz0OhDoXl
uI9ieb1tlGJqjStbWYDhR4EdbgNamv94udNQswQEyDU/CxX63epqU2N9MRKop4eQ
jfjCQKfmTLdi09WYD44NBeor8LBpQsb6Xkic/ITX8yglcm55E3wJ//avp5fjEkLZ
ULBclyyEXIlywiydWHT/tJv8mbUT/kLXSyFKMnXHbN45vNtaAJ3UUTkjA3/txVzK
iWtb1Rp2YfT9ZXEuGwvI5uG4zO59WBASwbHSAC14/aTmZTQYBqV1T9cEphS+R2o5
1vsKusC+EKYN6Z1/laNQ/yBMFp1FD9VAYDjRKBv3cd1rkvgD4eWIuVpn1pqzeF/Z
aG7Q12OtU6w5WRFWMl92hvx6TN54RRhTuOCHikLWfhPBSzeOOyaPxtSXAya1JKdf
pKoQfHyjvulLCD3cnmj5zjQ6vnry7BTjyM7bLikvgbs4S92CNe4qGieZzoaIvyf6
JTYiTuMgRCP8QAmAqib/r4yA/Pigz3PARktKn/lWfvxUpXNvAQZpBIJeHPft3QbT
qMn7MrQe3QOZYpMql5vSgDN144xN5PmwmvCmPDxZkP1ZzVIOQNdneXpoNNzYfZY9
nhM2TgoG53rcdFHaFBPjR6ZQRrNO0sbXOMhaC51pdRGU9Gy/UshTSYp0KM6ABjoY
QYZZ3VNEeR2xyByN8plMnkxpxTNn7uJNfesDtHD7eZeTDnoecP3onoF+RGTpNWF9
k2ZRT23bKe32SnVYowWn6eOKilGDXP45gsJjwG+8J0xZnueWo4ln3PwUCSvtAZBQ
XQW5fSfRvClvyU8dcaVpCisF5G7N3o7p85gj7qWmv8z7AmjjeYKQmAI+W+9Jme25
UlgqwOUipQdqfLt98BC8OhRtdSH8qG5LO5+Jb9yTnfeXCc2xjJmbxnJb4Xl/g0N2
CxBJrj/qNNYzwhovteh/YgwnbCA/Fva8loStUYJQQEIdHCwGq4/+zYSpWcnz/YCY
FsZAJtEYaMyeBcubfG+KhqJsKhTaMV7MvdUULcDLZksCvPDi4al3PC8jbzHNs66Q
PCaJY5BC9QfKdPQER3DhajTcxjfAZ9/l6fUMF7DdSYCCCAvaWtCrEio7ZGfakKOA
hQqQ39vic5ms/BdYajqOc2K88MfsW5AOvGWL6+E8r42l3BBmpENia1bDFBqFhV0b
yeiEx6CxmLLx8zjS+xOAO5jaGjjQ1HmWazVOlaZugMRe5xiIv7lU4I21hQ88FRVo
b7xKykXPItmjhOfaIoOEuVmjaW4Hbsy7Y15Pa8K1VL9K7atidbEQZPZdGgcJpIoW
pmeZ+CALChjyzO4ZtsPTJsRBeLoHewhfkxhSPYN4BjqGF/fkcCoIRgLobBTrZ9Lk
3qYpX6QqtJRX0Ir+CeneE/yGXLHfmGC79rxlsnsr7kuyjBz/Zv/I1+9JscfGZPz1
xFMQ9m9yXQGnB/XiOuemOtQiPUdwNwbgofNU8AF0LISo0SKNA6/rD5IT5GRjRyiO
tVA9AF94bis3dfep0WXi/04ES+h+GmqTRyL9GNl3A0UIuRWG1wVkixYgHI/7SEZ3
rJulf5jncwEAxAuxDR8jkxkoMna04Q7gWsiW/bWtk+a4dC8/mxD85Vig1XlDiwAO
SdAcRQh08TilQ/SCD5NLjwZm2mHad9mW5gOrF6BJEsZr8e18ORA7z8vnu7uuka8U
6csNhEtA5tkSiJtDZljwELqjlNCGFAEKkkzGgMoweSWWF+gZr3wK6uQ/muEfiYKb
bcEj01SX7Lyu9SuHkmnXYbUtnvnlBik98cgiQXcujHx8vRDjpzNc3JCBAdgzYq3F
Mx5MCFBlogPmzRPkticL7rPYGKUBO5fZaFcu1TwVnTHOb7+QgxBUs43o0NacC4Gj
7e0CD6wDqzAj4T1MJw3PTugzjilASozrAA2RVzUkgt8V96ov9CRnYUiV3JhJH9cc
8yb7mBm3sPuQXZwamiUz9WI9ztjUFgTFb0Nzvu5Nj7i3EzEnqSAYOuXXXQgMOPTt
f9DzAzMlDOv0POoZEY8qHsJiaSiTKgLp2Y2Zm7r/Bh4M0gUIQ+YtrkxcKx1Q9MJB
OyzhdapS5cHZpGyNcY01BDaQIG3524ZcNQC9wavzuDGtnp6YHqsiukDCuQ28WmdA
QJNWLugNumn+X2ZYYnOzJ5RsocXrnwxzRH0uzYULs814o6Dxnnw6T8OgqSgdyv5v
7WbRb9ue7+bKL3N/OjACTHHWiVXSojsPGyG9ZJu+r/X1irNLRsI+8mVEdFNQ4USq
FGCFgtXyBm9gfIkeHGi3BV+Xw6h+aHVgkPcl2tB0yHPRgKbMV6VzPGEGYkO4Ut9A
+M8F+n5jlTleh4gojXeuPJEe4D82b74Qxya5q4BEeomeBMDkGEQ8H3nknpSo2TCc
dERAaByWIxeywjFobxC5clQF7nMSzjSyqmpcVUDuPARlhXAhsPBmfo5odHb1WVAm
ckIcmM6tdJnvyXugvdVK0aNjSA9BFIXIl9XklL+kDIqVER8ocy1F2EgSwE60tgIg
MUzCWK25cTLH+5QksAOyk/Enl72+duocO/ru2RufH6A4cCldo1TQPmmoTx58Ofns
3MyQQK7Yr2J4fcgwQrw5A6ld1eKI0+4nVM0xLR31XZfywMi7+ZaAmuaERkV6A3Q3
zQBmjrwZdIHFHc7X/qBKLBt8CzAUULTyhAxXnpqciVw6ZJNH2XMIurox70Jtvtax
gb95Uh3TGPELFw9unKdbD7vI2BGw05TVapRNhnzbkxozZ94r1FVQ5K5Lic7v7O5X
u7LRs7EjakOX3/OicEZKfTI/Cvfe+lGIoEOEuzy4tS4kPxR4Ym2A8gXjYb2qQiW1
04k8OipbSbszbJ/lSc407+HlDr4lvD47CdQV1lPcvEVgqsPSCiXlkIHCETrfP/QQ
YQfWi5l9XJGRjMZw865B2D3eU+u5Dw1eQUN5LV/8we5voCwRWpEtGhGaZaIvd/NL
H8SUsIIB+6+NUYd3ucDlALNUi3r1PfG4H0XKpfTjBsmDQbXtBekYNjIOEdYEdrhE
v6l+W+Ti8l9EaP1PvwFMwMwHCgU7937aa/GgWddQR2rMH1KrlX2pChGUjyHqpEa/
IgD1ajp0oPstA/AhNFchTeUSDhXRluQdQPD6p8GbA24ltxK+LTI91VMwXv5nHWGk
RBqIE+vG9spjBHwIwRnAxKIdr6zUmT2UvN3sdeF/nLc/PS75TXOGI00dsXGQq9Ol
kBazo1vNpF08VJxHlOwghRxsE91kdTSZaBRvMKBdQZaBwqSMCkN+b5Dbm3BL79kW
E7BmhBE9FdF5bxQrqNAgk8oqhHL6Di726kSS5daA08Cng2mFONwMR1z0dw+rMR8F
KnSzrinpmzGwgAzISqFGRStyMxcqenYghgS4pqyb0cFwaMG7P4im3HEobjqAUHun
yKbqJo0NZGkIAKFmcL2Dk7iaTB77AXgXJHr1fagBKHD17wSmW1T5Iw8rFB3nNZyI
6kGuq6eCx7ZcXxBJWCzhQdb64Von4vSy+KQFyyNtZeFj0L2uduh4Nb+L2q8OkBY+
wdVG+qcfql36z1wVT5j5SeYfrQ5qJX2CD7lKMa6sbpPWHsQiJQt2vFAV/Jgh6gEE
d/j9zmW63I03rQcrwHTXBRnNTxmwQT0uwX1pb1MTiLpOaOuOxrIe76ZffVhzG4lk
oIsnk276djZjxIQNDk+MmIg5YJlL1wRqIwLENFmI9hy4BykgX/nQuRMl/e3L4MuG
4hxP1Qu5zlvt7uosJTiA9lhXhJ7nmes0mc6XaphfzY8wsD7eaMnpdQw6QneudANG
fp2ULJfU2hUYvyuS+AXxPUGo7uVGdBs0OhUpoNx+LE/f4zYIDb8q5BGIZJVLqywS
7iXGE7xEsz2f7ecxwhpXfb8IqtqKjttAD+XUgdc5rkx0LZaqT4PDgYd83QT+aS1S
LK447cthFD3vUvSDiMSvM1GkO4zU8DoL3GwTh1Qf96xIVrMVtkxd/14AEtKeDxBa
igpdsMySx5N2htueLiLg7lbR4ADQr69wl0/mkm/w0EtZQHdEOTINAIvuaFox6pwm
Ex9v0kjPg2cVWGASo3q8i3sVElEZh9lYZVb2Gu4fWXBS/iCRjL0280XdEj5ZeB7j
r2rkPKpTh0vqCWjtsObfho2uW5UeWa6E3y/5fruPQpFA2VKUbeZUBAEbYn4M72V0
n9FwLjlnXs66kVY+IqdbLzsjhj6ncKZGXteWPs+hj+13kWBX0wzF6V9s7TX9wEjm
5gfdMsxj37TLXf4RvZ6AnpHhUdu3TR3oXjn+mQdjH4+A3ZSG+y3Z5SyiRIpg4lFN
qR68wwIoPMlnKyq/0Nj4dRtAhXRu+3s5iBwvlwAaLN5O2iC/9UzTR4C0IG9X1s8M
THZIQyeUd47d44aIgT+RNHWAfpI+57cOjR4wnw8I/btxkHXo4jd/tlT1YETOdTOB
/hOW6V9PGtU3xcbGbZreT1ftmMAuMlTH4bwrADKQtL3aXNRCVpjC5IZthhECfrXA
eM0VAlFv7ap8jCU/Ie1gdRZnm/FY6CKdZUt1seXYwvV31F/+Ia1Ithgsr796Lxna
whaUFfkjCTK4+rnOwNBcQB7LFxojBQ1WGSwDW20lv53zjnnYaHCgSjBUoxfVMUjG
Wv7WcyKa1Ne+vKdxoAZPMC5LjCZPbHUOyiaB2bY3wUIOsyXQ/3YnjNTVeVFIBsKy
fj5fVgPtYmcqXsJRk3oTUsf0z8sH+ia3BrG6T1q8rwK8ay+rYWTXr6kq+JjUWCd8
uu/mD7dpPHMsME66TkG2kCJmyeXIVVUriPsb4ELiI9S7vMhGHRLwIJt/Il2s/QHf
4MIEROrfEd5fpdgBr756NcXj3zahWsYwTmze7J1jMjbarK/zXATckkIDN02wHMTP
VfKQ/67knSzgecQNS0t0s/guB4zsVo7meoe+jfnk0JGryBIykYRkkhAeM7Wp6r2s
UKWDqls+9C5pEfYvuWghlsyIhvbIsRMNoeHWc1U5kYq0n97+1VyxUOSLrGAxJlvX
hUDzbkLeD7zL1L6h//Ks0ODarUxHnrsZ9/TmD78nNqpM80QJhc9k/AW3m8Fc/8+5
BUEFCOPnIPvETSMOgsbF16xeBpF46t2ZvdLw5GRUktXdbtGhRLN2ZI7wcgE6mV/+
rfZQPxDPJAKEhoXjtNzvMBFPyAhtOouBkK8QWd0yAGRd/R8gYmNMb0b+uGgqrp2I
EWgmavQjWDneM89Bq/iEJfeLmhzz04edAU0ZZtrj6Wr2fecC4qysuazRmRtD/3ae
ZnS+m/j7ETl5mnxhdgZ/vp80bbDHEYoSvbL/Xdfh2UDnrPH61CAXSLEbM9TTke35
QNspu7cSqrhwRO6m4GWUs3qcpMsZ9Fq4IeFuV3LmTXfjgJ+PbqAuwaDIB5hL/A20
EGGpZWX5bHqzdzyckeAayf4yRpbRTTIN1rPRvXhkZ59C4rnTgVTbBhNOQP39yy52
E8gK32LL5rz88ka/Ly6gD1S0bRCEtwlxfZCSGOPIPkbyY3Sh79K5wtndH8o6P7B6
7QR9SG+tPnivUHmJgJ0sdLmHg/oMSLiDxC9Q9qIH4ThjoO8WyEPXZj1AiIqrS3j9
8stWj2TGD6qlSdtJ/FpaTBvSaC2+O3oON57wm9KJEZIQ7bC0R0XPO6p/UoKAmHVy
S9F61BoQevDrGhmXmNPMYUEyHTW3L3zIYZtoBgBndlZosEpObHVHgN11lM+y5Oaj
f3sSJTJGYPmIAfhrsl8Ueku4J/qBa1+pv8Ydr1sF/RrHS3lYszSC0DfwuUqBGoTu
KeQhd5DuZK01mhL0gE2ISZhofNKAc5vAvT6Z4x2e9pubjPB/uV0LrNSpnrL1fH9H
CLTtUU3V0hYu2swRUPiawwEVNfrL2iJoM76E87wew0XX7zrKNB4zJD8lJ5T6TdBh
8cbfvUFiGjwUYoN7B1FWNtZ1VPSHHaXxy5ujXSE82H/hhAJX4Bs3kqQ7VdwSR2bI
nY9ZovtUoIUzrjA70Ocxi6ko15AOnYs79fPRvnuKZ+ylVE+B+WX4dhMBhjStBhv7
gz1YWXZuVeXsj0HSVaDtcfg8xlQqzOs2LyVOEUU68cwPwLtpuvuiOVE7axnIXExA
XLfaWnYrbCQcvQSdMUTHgP/ceJ5u8mmac9uMNuPy1KrQBZGyD0alXht5jZd5xG03
0Lu64dFLCRpqpQaGkXE09MfAFy+XMkdDu6D3Hy6IdNzYomiViNnLNjuIbUEzypwq
uh/B+HDYkmS8u2CpZHEHiXoRZLhBugEA1WJKL5tlvnsbEJ1pAFHroCj5CgIl1BLI
lb+wY9b5VaJkvzUeiz+td9owSpBM+H1ssN8mJW0LUyPxj5luYuu23s3o8vzlly4a
2Zku5uEFPpXJ/oe/yfer40I5XOPBRxeJVryYsIIhzi3D5Eb442QkTtKQWc+3/rHe
sbCGfjSkf3EkbpUNEw27+/oQMD7QqC4TtSa1XNnYQvXYyLv1XaS1oAonR0HjUdCH
WLXi3Qbui2osgX5Wm2RSbXhboJ9ASy3NKVoaZYFkOJan+F7fvDsk74L5YB3ZuFyu
Q4FfTD1g1vI4Faj7SKi6Lly4CywQ7YaAN/RwGJmGnzJJa4/MjH+TpZJIjUhO0py8
f0+v5yZdR5aL5g4WQYMC8cRSNMyyIVEIy7FOieqMJKqW3MHuFHuKpsHZq9xWOtgl
CMp85p8j0f1y/AqwwwChLGIHEWAykG6BLCgilQ3hpso1tlyNb5Hpprua/IK0TUbN
+bmgfiud21s838Gm0oh30JBLGc6v3sK04NzMCeLOeyiU2khPhjw8ML+46v5Cgcqq
oaGrftuwcqIWvpFugE3t3U7Gf6SF+2X9gjAqwhes2hiP3+3OYHQDDKAnqQIP+B1r
EjOEz9+iBmEZw/crId64J3LnZp2WVCIBELd9jDl2xLPoY24P66uEGRxysumfNGqM
AS5cgLFlYq6XDRIYth+Kv/OvDm0S0cn//3OIsdx6EITNkGmgH4o3LnpxIko6iBmE
UAk2mMrAye1A2kCWRx3IZs/WQ0JkK3ZRrWabBoBizxOudlGI7YhMBAkQML1gxpLn
2U+EkYuNvnL0jBa0n9Mk7tX1OGLWgw/Qc9o61T99IOtDqJe6zUcXmxV1SB1iMdyh
o4bsQ0hlTP2tfXck8MAQytKqt+FZo8jJQYVtYbyJwPRbVEHAAN7FllXPnKTOzAiy
SkOKtfwjXTiczvJNBLjV5/0Ire3sjrXy8HxaoZh3LZlTd24ha3opwd8b6O9/09uJ
a8m9bc+/mITm4LD7yh77U44vgxtMHxTu/VMCB8wYEL5zbL2C3TMzGwoNwWN/TWEc
8/EDGE2t9Jxhxr3C2xmQN35/iBmOCBNf/604FZ6to84HnnDl50NcdccLNEYRQ8vX
8H/iaNWoGeC9VTNlhwKGRQFTYB6u5ZodmHOU5d7kIBP+x5GfD53JVhrXEwGBhfES
WPEwcLBHLY6C2zr+wpGMCyNSDRc60rNfxvLUOgAjSAjDeM6Mltr7gPk9cG28Mmql
wtew8ARGcti8SDVkTOFqQP8aSyYjVEO2kh3FiX7gApqPSNc+ZBgfihOrrNe1MJXs
NaGZmfnYQh6vX2hlkMyUzKlDmaSrZ5MA57Sjd/Q+Hcr375rqsqKmz1OHgxpQiokT
JsGfh/8npB9VFCWL/d3Jxv+ZvO4DlXuF17Fce7pPKn4HCK/HlayuEQVrrGk9YOIU
eP6JHJvCkQ0toU/zor1Z1xeka6WmaMwPbFAtIU+lt8s29kKcqlUcQYwtaF5B2Vol
OsfvljJlzZkC6UUUZWwrBr5slNMPVCIBxf2q0sVGvof/HlKns44w13OklXAsH+XS
OkOZ3qYQKxcEBxt7gJgC6EX7846Sul9s4YnRAuzfb+o/cqPgACGu640X9qgl3V5t
sHgfldYoXBZWeevn7XyMUGHvJztlDFIPAvOrtBZRWIRUWg1nZ2m2KGtzny4hZ9Iu
iSXxF2d0c0eISXpNOqq3bPbykzivZ1CTsd6QqxuMbNQ43JVdPNLHMUwS5RQMT38P
772a04TNmnW5jXR35G0y4eKEiUMTT7vdkklG1/nnNqOfopIaVJrlm1Wl78E8I5eZ
pTfGX8ium0FsqDzmo8qVAX8EHXYR4hfMU6rWtOgiA3Lrxi5+xVqkP+G81IIWrbBY
/AWbBmi7h8CiiRp8kLGyoJI1MvXjW+nfkgj5AbnPhRa0ilVwjiESXMMb/GhBj7eB
850b6SVfArI2La1buWaxeOmNFsVANCAqSml7PegaKMmO7Lga258oJ29MJ355WNur
Fw1eUxAnIOdkY5gekAGbkp3mm5YKQ3wMw6YNYNC/X9Y8sIwf3nj9Edi65Maj7CFp
axyR78xrcweyyYKVQiPYiErWFcDl48USW1Zm3Usraagu4w7aHF1/jS4dqx1XMCp7
2tm+cnGU6GlUgcgJZJlLZoIJgwLB8A2kS3vSi8aEvsmK0LAwfdxO5cBObzmr44su
JWvzz3KSViJp0mKkC6aMASDfnW4TnDVdiGZTlcRaut3ddneLouMXpW9ugjQ2xu9e
+TzwDZEIH26/U3WYDnWzL1x/RKRbWSMahrc/I2ZF1Cm+49kJ/RLJrg7Zye2P7hEM
L0o8utmhLbpLtaTnvYmkgEZfvsvILO9L1Lz4SeWXT7yjxcp55BpXTUsiyukclyhP
f68ehUDCHLvQJGBRhK4IUQrSY035MzPS3YzeoUfGqi3/LVvE7qc42DKas8xd08GH
fLzjJAIoX4BpLs05oT9tVM50yfW5F4Jwe2GyB6vmF28gwU3I0wzEaz/DUidaC8kQ
mripMWSC6I1O7vBySGULi9IJva8wR0qsNH0qbrY1FDThsOrpmjZo6zOOAUElEjb0
5EdgBVdTRj5muTi19ePWC2lXNUzOqdNX3FlKuLzp5IeZh26BJRka3e91ZNzIZXHy
6g5xgXJ1ozMV5dZXvwlXx44dDPcJCFvUIflX+Lr3V2118v9XtlQOl8R9av2WGkXO
T/lRSinwAbnVJ7sE8AwwJY0BIykOIcpIGvNWtvSCo4vY0w1uDFI5pIwuPfzh0oGZ
V2GbiXykiKCwe8TboAilxWyhZFkyy6hofwQkB+/b06BVIlev0PVHoBO1/mZTo2Ub
LQM2ZYNgTtGvch2YhOplfFHi+IbsJZm3qOfTMvNmZWiQOyjdlKAxB5k9CMV1cxZZ
C7jm1eJaR+tswtfIIg7GTI12rxht8sR08AmhrmLayR6ujtBFu4Z0C7mvWaWSo437
LB7aqNess2n7vqi/Zb32BP+GCzjVaeIerjHylFfS5sUAsZEnh5P4HdJnQMKuBcfP
8B/gjuUMB8yIWq9i3Y7JrrX0SReczfNRAZzyi/Ye0rdsT4DKn/0SQi46nq5z3nOj
Ipzvlz86QDuS2uzH3KvbNawJwjHbeYW/hRQ7ADBad/7XYrhz/ifVDJVxlAExvvHO
n1r0rxv876L7W6cbvNJhqPSmQdaOS5HPB47YY692NRG6baonxeR+2cBlNOLXd+PZ
qi4L7rHtRUgCtPFmGBwDOmRJC3xD8dJii6bRLTaBD884IzXdDvdfo8HqEUML+a+z
43H2wnx0i+9yZZtYGPKJvAa9LvF7T+Vnzp7Q2q7E4RTmTglFLmEIN8iY/U9hCpRh
+GAF20BNZMR1gvFuLBIbJrCxi+4DjiS6Vk8LUHCt3JFQj+GSft5fgEY4eXYLtkiD
AtqAwlnqaj3LmW7PU+htFlBGCC3B8JjQu9G5kP4mV1YuoLoThaNME2VA2Nezs0Tw
QU5dub/9V5n3jD8EDLiWlIC7XJ15IzmRlnD6evAvcwLMXzsVfuhoUG3D0BLdhAs+
403ZQksCUer6Bdu6DJgNSV9bi1LIpBzfj7qhimxXJbH1vsjquh4M5BUxGDsQQLkq
L78vExOkk1fOKJayM1O7ma+mC0jdmznW/WuptidtpbJAVZS3BEdMGi4MZ3fVTyOw
kr080xJ4dRGr6p+4hv3NsJ0Ml1AA59o/pcYIM30Oicu6xAlZxofplKojvVT1S1ch
ni5LRngE352s5cwL0DRPSp0Y92qc47Qw5Qf4d5DueU3YwJHPhu3eOAgiaPo0VdT2
Aeohcvivvpil3TCuiFSxQGb/MA9F9a6pyxAj3cMwx185g5gCK47N4Uo9JbgwcQz2
PKooVwEaKyPRjvv3KyysHP2eZy93LpFyY7QnCs3cKkrLIpw11mtDNnaosIx4OIgN
SQO4BoUYlttF3TJSyN2WzK3+2aSr2/6OPpMZnUqlhRdlWVt4HsIEcsq2L0z1HjT9
QSYsp5tXNStpV6DaCDWK4KsofrELO5RtjlAPYY2dxxtzPQ+jISZ1cHlhpJoNhwuD
zmYo+w+SOCocp9eAtHxf9/bzX5xBoJGw5RlYrW9loBuWVix/JBp6Bod8X0mmE3Fu
E4NcINkqoir9r+HKwCwrYGBsDbh7fKBCzu00B1HlUSSvLxLx33nGx7Q/X22rsQWN
Uj+OzDfnCp9oWchv7gebjlDDJeRWHfqg9GAfBWtP8tjz8CDOlDha2e3IQxTefCxS
sDAhcwATh0VfX6CWKmZqiAFWbzzGZcoLcdzg7QJd9E+shq+TkvLVzS4qvYC3zf7L
BCZGBWHBXJWtF2pqknZdvBs3GSI/J5kHPnmDVSalyqz/DjBBA4oDNy+EJboDtiLa
QJ2/q/RkOoFEjUp6wjQ1iv27JueJSNWhTYqe+eENiaNuww/WfVOB0brtJ+02nnGA
r3WcfixdNeLb8IcWh++XoKAZdnUMKesOp0cfOUSObn3bJGvEBHDd4JsuANZAo2qn
Cmdfv0VzPbkSqPjX1JzNhC3wv95CftGEi0xvcp6b8zdz7qrH9Wp8KYqIgDY+4WT5
wC0ss0PeUReKAT7Y8B7VGqxlLVuvVIuuiIbSfNLYiGEvyU+kcpEhJ0uNf79ecyxz
2mNC1ogh4//drU0or62oimYwmu40GTsnc5sBWQsUHJalgZTWUNFx3SwXXgYMRYlA
4Po4lkK1Epr2mLIQzXHhrjIrzDOZv5s9GkMVgmSC5KwjdpOBsxRiVe+2riI24CU9
9QB+fcTdlEjZ9MdgpguiFxB6fN10vskqMYX/xWXwFg0ha/CKhXycrL7gJIr67P58
v5PBLK3KAL3qrx5PoEIIxgz9oeirXFcoTHU1mCoib7mrRCjhXCoiWr2hdjxX0Qik
IvImQKRubX2ri7hh8XumVP/xdPo1h53TKyarN67JG2Oqrapa/7jDOBE5Q0rvoIuv
sXxSl1+pFx8cd0T3GBaybuCybo4KkxC7UrEOP5M7aL1WRnMf+qAOCpQo5U8saWXT
Nu8O/Mxgq/1XqzSOPzBc6EOhowb9Z7sCz9ei6y5Wxnks54d4VDw2JMC0CEk813Ao
z1hKEbb11sFGhiHhgTgnUYtnldatu1zw5Ed2pdZUagTnzYgkiamX/wxQYhdMsneo
XyIpilXp7PUL/wu1bTXJArwwnmguZWBDDDuKJu3Ixko/R8RYz3GzQ/3Mro+vXGEm
AFj8SEGVzS/hzXal8uSIqSYUXJEbvh/GBHqE1Ylxg/jCqRwPOgpAMy4P/8o96U+/
3RM5r1TkmEmz6vd1oQ3HL3ddZ0X1+WhU/BcCOxDr4bpdzc7//s2LLgYejZCxaah4
v8xwV9VXaQT1GX/vHZd0pNyHY+IKFWsjsg4+nb8dmq7f2kog3MEAWqedIQf4yk+7
p2UIbz/5jWSyxUEoILLunDMbEdYwK8+5ubDjJS6792DuD/F4wn0QkCQAeiQRqbH0
gBuHhk8yUHPcHqpBaFF/vqb7x8iIf02cBsS/rqzKAG5e04rOqkM7MJ6TnH2eS0wW
iBCVIx0WUMYzI61wvwLhgHwIst+Uyk8cuEC2FyA9Ndgkc0nyZpKz2uGkGjZz9AbZ
L4so1pNgEvJgthuT4hAwgY115aRdCWH1DYQEd7l0ryAFL+1CJ+oV6+1pAcFDWFyn
ujrKtbGRUIURu24jfZKpRyaffqJC/bhKDC7yE+6UCYexsRg1BoKxlydvUaw5Vwob
huOwOKg+noIoO/6wMirSZqfG2hw/dGHwSsdtEUQGq9myMHN11xERHPeuH43ct4lK
JzBAJ+I+FW019x/8LYcyjWN/hp+Kus7QxBycUu4L7K4M+1M2N8jtbjdPFUGYplC+
wp+ZjorAsbTE4kBEPUpSNCI4b0Ll/MCUdDILYth0RoupuXtFy5kdhMHGerIm33iW
ldmJxf8GS8oV7EZnhoUoBJ90HE5rf6/QN1mIzqrvhQxkvkJ035FWZBIJAF+s7UFp
XQhrxcPLHXeMz6tGlm/MvDL3BVIbX+80dmo/ZSouxeuhLxSDzRt2fZ2CP+WbCKfh
H3fs7hLwNQFz0EE3KU21z80HV0ern+PhYL7mcUHJlYOLgvlKfmX69SENW5oAbn4F
O5RVX2CEitrDOZbH/rc5ZkRqUJdWmr0utWevm37CVh+6K3htJZDbCsjld9kDxu2N
EnT/5frms3TLoo7DY5jp0l71CI62tyHExI4zAgKoZgm6gytRjO/cSUdPKQr0Kt5Y
J8KrhX5wWoxS9tZoHqTKs90iQgJ/88Y46nFBkOMkb0jTp7qmkFl8udjMwLu0hnbN
/lXF38Ts2+NZD0Og8RZK/dclp3PAAALN9Orq28OlxTCNj+1+dPljTOtoyZTZswJ8
T0CN2xKz4k1b5ymFuILkt/aslTjwtRoXm4edUM/Fu7INfzC5EJz/L+RikXyjMVVO
XIXfOxpZP3o9dmSZISiXThEbChyokjzQWNkgbCU5XB0WG8NCZlmwGji77qA3rR0P
OAsbrMEK83cpJrXhULOvgEkXf5P6LOng0HflXBUMahoVQzKCtt1MUgMie/VODnJ/
6WRxDl3txThOmWVUw8uLxoHRhHXrS5eyNtyk9gvUWrYwZ2Teq452Z3+RIzcm05jw
ug6ZpUxlKT0bxbE2iYTvhJah4wRoiBaMirkob8TytkSPkIGKiVz7K1u0CfdPuD8H
FEA+MGa7qsu1VdGPx4N9IDE8XdHiNYuitRqAxof23Wpxzoiqo9AuJQhbIF2bE2Yk
xIMqnGHltSxpvjFRouVjuzT20ly2292p2GCF63GXBLhbJqux4CoRM2asj56ok5az
qXd6GTVBL8kIFj1Q2e/+1+Ndr+IfvvQH4pW85oNkxYGmaDNL45ujNjEnqPi2InQN
73WiC68A3pD9knxfMGW6I450Eqy6zcKlIbfQhGgehxYH84cA4r3bG2V2qwqcJl1p
uhwDaaV8E0cIp+M6tBVpsSBwQcDERXYnMNL60iOtXN9A5fg546y9uzIjG8RfB10b
18zT1VQz2wX6P8s/IeT1C7bdhRy1ONH7rTqzFpC+7MwwUh/MxgvMhHMIH6+Wnq4f
P5VD/INdu2xCs2DGbfZx6CLvT0xYdhhjE95rpSzix08cy0PsiPnIYdcL2J7mZiXL
4aJ5XZ6vJF01pj7Eth+4uxtJf5W47H7wix8huXSKbUD/oRF8Bo2ylqjd2lIRL1uE
W4qJrNt1aC7TS+XoiU+NQikhfEhHSfSb2OUVWNwBl5dAYQMeEJLW9o/ctBDo9bmg
ia0jdEMV69Xj6hX2kAIcZVgmznNAeFeMsJrpsSRtpxvQpZXRNm9gYD88WLp0Gs2S
OigmfqWKeQBi7Sw0b+ni3pjHWcZUO56lPWMzi/+EWodjZZNlHEMI7Ozw/+8UdIyp
79vjUIWM4fTXTAZQt9jJ075+H7lBc0CnhZqVK59A+OOaMETWqL3TCwkwQWc+X8xN
m/c7Zg+dIxWLHs2hnZaGWcBPXayk8IdgSwOZBxXnSqOCfw7tQ+10O4w8A6qKjuWs
+/bTpmZFMi+eoaKbgpXn3yFlRBysPlSbg/X02V4qcysnJcOGTcdA3bNONNtiCvSX
Yr320NFZ3uBkbEgvTxNCABpA7tgSA0ODwWVT5l0kLPVwviXy+YnV86UHaAln4Y6e
kzud0nnepi0G/jeCpeScZLBosOoFNzNsqSuYzb8v6NogAlp2FswAsV+0jY+ZX5xW
e2CdTRM+DRMBSsC9MLyYayQuwFyr0g51dBcxzLPZIUnZkqyIjrRaiHKz80ZWlyoM
4NhjeFjdY4K5QiHXDAn3aDmo7qwWul7Hqsu5Z9+YaR5Az3FRVzb66YTkEZdJgsVW
LVq40mmN9exgd1Wl/o/HnxyYEKg0Aifw1RVXnbFLUGJwqIdgnTsaiyfrljr7Z26H
HKFfuhxVel3zM6k4hxShU7++MZkTA0kNkSBZmOw7NHY6h7zoBfZ1z74RcbocvTY0
gUDczPJjtOJLHnX75BzzL3BaTGQzi/GcROgeDqFnrHgfkLImJXOszGM60x4XO86w
JIBE+xst16msVD2iGP6tptLAJy88hJ5IftD06QWPQXb8M9TYcm7MW6H5uHO7l4Kp
2yBcezLL1Zzn9WL3E4vXMuSiI6LncyhBlnlgHecEXKKNtgCLzwSKcNRgJAk6YDot
Ha8+vXx/Q/5/alilLCp8ojb45J3bXZXVw/i/bxyuKVZlh0LMZGTvpaXtZQ50v+1l
XQavE5KHtXneoRLqsEWI6U4oliCavsydX3z30pVowyoycrgYN7JZbK1QldHiDAlM
dthY1GvCT3J2y+ux4k6UKyKzNx28NxaHh9xJrRKuBhsinOIvPCeZeouZt2JMDQRO
1Vj5wB9j8T5RqXztsTz9oWaBf8q+KFFUSv/DSbJT0KtB0YYv5UTLs35q9CFEi2R2
aWoW4GPB2/6z1NjQoaU1TzBwMXMkR7aURn0qFkyAZVUjGkFJVUuWhBsNM8LLYyp+
jiXFcsurZ+myuIa7s3tbRi3NWby8Pv5xg5ogshzUEIF3n37tNeJN/Q2uegv2JDyN
f7UDJI1mC6T7R3eHfJWdwqyKdd/f4CL9go6onOS+rog9vll8WaPvB3fDY468Jxqj
Lp3cFXrllotGWunu2zz/o51FayPDO4esjsgNFGWMG3iLdc3hQWdAZRAAH8L55lsN
ekB2qlqiP4Xb1LK7tosOiS4a3iupBCxPF1xZ1TCfLeIvjaWnivZf4WExG9SzL2ev
605yFGmz+XMbwS79+Uq/b4S1q92B7K2U5832eT5sXrwMexKgEzjTnAYNgtdhvfh9
ZlWnLZRHJbfb7nXHPn39SkYUJr1zODe/zWTsSMM7knp/6wPYVJmTPqUDUVrRcREF
d9RvTomfUt8kzz7QiNBjpNWAQqZZOIEue8PiHTC2+IvoYxJDXYKQ33SdfitZSYF/
3XJq0vswfnq5oeNifE0510aGt7+7njOlY/V6rwchmL7nyzVDqWX8t2+WXSvBkDFw
9oVJgQk7NTGHbkofkvRxhAUV6Cefxfren6xL4K5zne2o3IlDuzia8mhGHw5bN1Qa
f17swC/uwn1yngf9zW/V5WLIgTq2FIwtfORWhlS0G7jwysiwPtyiJo8Hfgl/Y9v2
QX+nVSyvhRnXY5RxR4hV7kRQ5LkjWvcJTpJnuXK9MaKFZ+v4VrOFgHVDqmPDYqkV
56K9smCvYXBEpHV0XNeUtkjeFP5pdpEfC1rquofeYJTa4eItAhnocmVurPANl9mz
H+bdYpek6hRI0eN0GHIwnajp6EWkp/iTU+gCbDg6YXEngLMN7iYMNjuZVbf/wrqk
n4sHNVCKc+Kp8d0Nw8x+co+50L/p7i/ZRm19aS1YP4e27bPz8s1KpFaKlvbWH19N
mdb4YKebtwutNSuImJm7yxDQlnCQpIqEAJbDOWU+q/oWt4k+XnnJVYIGv/kcXWeO
oLVGf/OaFG/nCHcD+lB6J/+ewUBG90ORRYrP8N3vUvjsFMHM5HQxjQ3KRYMVOBb+
aTTYwgYC8LOxIR2m7kx1C893u3kAb/naFYCISs5e70+8r8lTthwuhaHvVFxisNm5
BAOVGKMWhM1uZStLOIFf3/uLgQy4Cq9RykZLNqFWSZa3hf1h6LtGmooFoMyJPzfH
MpaJZAB8ljserm775tA38qpgJeqn/YjRNUs0w31aSBzzHhChUnnWu2SxGeGsu9AT
jyXzWLi2m4g2Z28XC8uhZliPOihN6szH7AjoVPGZ/jz6omzcYKccPOTJyGNdBwnU
besP/SW0hlDGObUhAGpbyU0p0QafYKQPCS3LVsi1uqvtunJMXPJXwQiV4qgxWQVH
VUtM1a49fPkfMhKrZZgXoZsJUczXf8YQNunYllLg6AFDTyqTynMd41oJjy3mJo9e
ZodLj8J/qJjyxigttCZw7ToNMrrjeRqWUSqqshECIB4cmukUv3USoONkeI7NgEyZ
Ygko1Vx87m1ZCeHSC/AJgZ5GhdScB5+M8eSQZZNHlcseB4TP44/cbBLki38YssAT
GcIiNMJwIDlGrQ0UPoAaHpcob5KtH4NUptDc0s5ViGVhnYdVDo/gh+fYceCKr4xj
YUQ0tu0qWkl2CR4rEAkD8XFgHN2Kpx4hyUSlnsnnjVRLMoAdG/BTGvrLjPQ848YA
7JhV726NXDGft3PeVji36Tw8bFYRnMtFdkO8hk8Kydg/J2QXe2MUuk+hD9nJOsNZ
jeIYpBkmnGV11v9LSYdFQdfzZSA1/4fonDlhxg7srO9wu6ez737ijzQd/HdNzWRi
cdcHCF4fZoz3rhTxL/0h5xcA9/0Wlxp8mJaLiigs71tbeBa6hd/7LOSDg7EW4ENd
OOMRRO63wlSggCjxxaRCjBJrbit7FOqpwYH7/Cs0G96ZW+8q0fsUIVVUqtaunciW
0XWRD8UgCBBeYXzQe2wm/JcXThFC3Djn9ty9KILpjVUqHKQ7t8harm72kEW8kFjy
wzFWp7YNLSZTgzPSJTxFwxW/tOQNwGxcRdHvxRixqUzv4LB0GTBOwXrfP1vIKTlL
GJCBU5zeIEvVbsKkD5uwvLErPtMtSJ/8D2mHHyGu9VScWg37ZPD4FHPabPoXqc73
7zsuSmmIanFYx6HUzDxH95c79ujhkoji9HCG2JOnC+S9Il6972eYy0pBiKirQ9nW
QW1QefW8iz7n2lSKII5Es4lgerSwuLwLBdapeOy0FUVJVismu6sMn4BroTUu63yi
FjV7WDhdGwl64ocEaHTY/oq1XlOPkjPES3lzCxifBXRbh4XEo3zRsLAMajovyj5z
OUtr3UKrNcjOGWxSUVoWN3cmzfqaMxUAytvRhWUtZqbUM67G6dp0zen1lxfzhvUg
g/4qN3QT55mHOdRWwefWtdJHP8Lm45CIHJMGztzQWEH3Gbu5RNXvWEOAOVgyEkMn
IPFfNEwp+c9e/ceZQMUrOYe92MLZqlmouezrnfzyd9vgrsypaOVfgPU6PuPsEln+
oaAsU+HaIqYb8jxsedvMcyQtEgL44LFEcCRnwjYRr6QLajuL8/srrTqzZ0XPdezj
KCojokPWYyl52lf/BEJCKpfCx3II1HyKUDnn+h0rwBa4ogqQqnN7bswWwJHQpSxi
Kow5sao/aL0UPjgkJ0elrgxJFVXZn2GEZzMmaCFTKX+5XO2yT0dVwVkH7/i/psV4
Iqo0dRkMLq/tgsxQmDxzzxEat469M6WAHFWyysV36DUv5MqAGKhwj4WAj928CU4d
8N+1/u5bLkVcPjN65KLewNF8BFuohokE/Hy0vEngNgmv56/bW5YjVfk6Cdrv8vYJ
W38HlA9waZ5Cq/KJwSL3wVWqZt8v5CEmPfS8rn5b3RWYdWkfNuVCoh66Ix5ojH4Y
7P2vvx7vzeTADvtGoiXt4OVb6NChnZshlVDGWPueenNUHu9QAWs9dDff13mOkvEM
xYEoRpLQAdRBn5FbW3Ug2bLdy1p/ISifq17c8qaChpYA7M1xRqvP1phqBcvTPOY9
7rjOJsh0RfRyzIPrKRcZQN4J3kxTSWKrnIbQZUZj40+IGpQUvd7RAjWm1eMRUoUS
+6C8DRCQmfIh3HKHgnF9PZYjWlOoi7gHprKU4zU06wjKCA7yE3d59ftlpHAV4Cmr
W/ev7wQoWYw65YJf+e/j7r+xfL8BBWYRc53dhl8v4HE8a1G/uh7LmMSFpcghZrGQ
ecHMqJ/L2Ps8vguKZDVfT/1uK8HtoWnKA9cZqgi8DXFu1F5LE1AXO8iaThnDl/H5
v2vViZAduG3T3Q/+jk9uEyBuvOi+0lJf+HngaBFHgr1t6o6L5U9X1wArFtydSWvI
Hp0CzHGERahSPyDq5quYIM0PuJdZb6ozz9KiYihkQxC8E7NU3wM4AM0L6uzfatsz
zoWLhtqI9QXbWLLZzP1RjycQ8g/lRM0m8CN8QThR9PC+cCthtH38QXxl0K3NdTOj
vH/bisl9OLxIxIFbbcsGuEUatgE+ifGS/qdtf00DD13R2EGis2b7P4hQa0PoHmXp
yT3mpMjjEzwxaCNZhBhhnIyNCjPSRv/cC4n3me6zYr3EIdY2qphcZlEmm+PMfa+p
rEtfG2++dePGteDBh/TW+fws1kjgCHPW4Qw2X8knLfNkq1pmy0GkMUUoGroFlBfJ
Wdwl3bj9NmTgXow6OEOo6hnZQxdlwW+8kV/vQu1O17YZpGaEXY9h0xaqWu8w+IZM
5Nbbm9G92veemn2IeoJONXsepg+96dQ2un4kDckyeFul0Rs5l20lauYH5AvuFNRe
krV8G1TGsjm5KzbM2NmhYENuqN6hYC3EA8ua1wBCzE3nnW6ajuYgKAOkycsl393L
GvG+ULfnDK7VNr4F/5veX8H4V6idqCijqWM5CA0Zh/nS8W10BJDA0Z3x2rZLGD0R
YOdXydnuI6v9l6yMdxiRlTS3FaHa+Ny2wX6qRret4meYBfbKKAmu6ZbYhGRn9O7v
5Fx8c+sz7Z3rfyclPWps4SES8qj9H0OzcIzGIr9Z5IefNPo+vEpjRXc7SFvyDjIX
ZJk2esFVexuw/5HjqAHefiit8pxLJyekYgPQ6gSe96UlCv6RRFLvzkfaBcD4Qkwm
0ifJs/nznxmNt7P5QfhzRTALNS6Rfp0x8JD8IMgpGJoH72Lb1zY6Ou3AS/nQOrfH
VvJCZ85U9QFXjGcCNCILUTbF2VFLHG2cDNMP+P5j42lVa9RFgfUScf6cS7b5PB6/
H3E67cH3eX6CerXD18flup2emvdnwBNAMZIFPecxojKWKJQALORqn/CoAX51vkrE
2Husw1S6uHEkxsSKQrzwZC+OHOo9iYvrQ61Klb8mmiz0YhlM2fD1OzxlhF3qGCVR
Wu3j5ZWsbbm9c7DwCKZCJylut1YmSbGxKwOAb9+8BmaFxiqepZLmDLIH8ONzwy8H
7IyZAnKeDpqGAKyKce9W1NNRd//9pSXCk9vVWQSAzf21a8Zg2jR87vYDiCqrDqj3
mmmZG4+5qvuz+XzgINhlhY+x+WV19Efh8AH7E9fopfmjmNh8r8JaEHzEO61UOhpn
ie9wksPkijFYq7d0Vn8r+JyRKDaQVvKglj8zq1JtK/cUkVkXZooGY5pusazW8t4N
c1S/aQrZO6yD0oVlsWHttRi0Vc6qYFEzXspH+bBJjUA9WVrG3o48ZMybqc8Gg2Zz
DarU+qwtZgjj0Xb27mORgcw0cscDE/D9Ua79EQw++YcOtEWdXAu1lWDtXH8hx0j6
B8ImkflG/16+3h9ZTHBG7INc1yy2YrpY0tZptOyLCpn3WICRkFDvks3SMXXKcJGP
sq8FQSTen6duwp9pi6SlXAw/BHoftlu7sZ45rYtEgnoKzmjx27KNuYXUno+B0Xll
7Ae2zowlXPJdpUHObJzYeD2qH3f4NMDa1mPTSVQhPO8fI0cvgOEp0UIOZAgnMC+H
D7AGCgHr7cNA+ygVm52cOFqvakdB6IKuxzNpRRbYd82myiG6OeucVNjq14PRcI5F
0dEOiBVZ+U5Hf5nufaCEo6j785lgYcBFmnQ952yve7OU5d4/jOUVoT7T3BcsrQ1R
+oXE8Fzeot33c1AxJzzkX9WR6Y7Kpqukn70fjhrHae+Iz9r+Rm/v6+Fi+yTqtzdA
8rl3soz0TRzfh6E7marpMdXIdHO0X3+WYqy+LJpeugFjb48cmxM/CJM5BbyBAqBn
cz9GfgpLRXEyBLTtGOkHTDe+MuSeFevKpPIMVwd6+Snnki2FRuu8GLxYeSAQxKfg
Kp69/FKz0Yr8HgBNkU9WVET3ej8/gZz9UwwAkA1jUQORshYBpRjjMZCvp9Osxk4t
eIjIDf5N+/wvla6N+hHfWhRb+wAlC8fE18knF3XmsZHxBX2aNpFUyJOnCAilYb0N
YBN2zLYNhcloiHzzBuNvnrzBe+53IqzRq4Qrdu78d88vxnzLAMf38vnWZXjGECEW
i4l5ABYpu5XGnpdw+wIwskzECX7gbeUz9gz9d4WQMXO6tbNvdk1rSUrq4xyGps7B
vlD7H92sVNnU1ZHDfw1awdTE81rLSg7uT+Cmsa6607kIzGfnkNwZbTpTqMCMn6tC
JncYkv4EkS6EJgRf9U/TP6tuo4Ee/pBgEmPw3sfDDkJhCM2eaHa/0YhUCiUiuIzL
KBrvMCbJyQJO2wWVfNGUGUQQVI5zmXjjan+NVrv5ieK3iGDk2GKpfzI9hi7e14Mf
G/bSqkcNruMD2s6j0+IkSEC7wcoSVegjCV0BTwCfuMWSaeB8x8z1akWxCgfV/vV+
8DZoCtqJsiC6WpNNpVTDMKPaIZabnnUJKiEQrtCJ3PrOV0QXsyv9HqOfSdnfA62S
ytuI4mtv5RGkja6l4Th3JXo3mVjCNTvCizILCmVqW6nG2NggcwNLivjplIUEx5rV
jLOZ4VcROyuUb/YQsqWqgtTN7OIS1hwTdTCwSQ4LkcQp81K627D3CmtPgJhifSzw
fDccGHM9S/CztHBg2dAP3d/Q4M2gNXZtqrTb42aJSZasg7Hv4AZKewtWyNXERe2o
csJ39VnnJqiL+cInUILywgq9SASfGkjAvUwVkAlVjOSsROJnwBORy+uKIK9RTfSm
2+4Q7B2mAIvmDpU0LeCARHICYEqVhHZ4XQiOp3bn4Su5fpMom+0E4QsBSbHhuZBA
9lCrNSAwQTdC8Q2gz6LPW24kTE5tzpVoZxldkwnclBYO1ZA1vtx5i6tG+9eGbYds
dBDBoYxEfhUr2RM4tCP9VNr1Nq/POrOsHGXPiJQU6fplTmXsC8SyjdjQc0elCFBY
IL3DFIyv8pCVnOpKHvAGen5ycJLk7/sZQdj1NxNGHYAvSW7OxTu/5SB4A9z83Jn3
xmGnpEulF05y1EXM89MrMxyd0EMj5SLtC6E7+PkJNGZxaUKmtP4zWTh3JEVPmnDu
fmiYIDiAOyJjZzi/R3Qjpxk8jnS+XcmwMU7sGtZh8a/Rq4A5n762qTKbc0QD7gM7
kla8bbRziZ8lmv99ZEZg+fD+i9ZIZzKuYMJ7NiHvQjh91BW/sdVPyfjBqKQj5Nwd
K2MOS4cf3OsPIV335wduPFoga6/nkPuvMwE/LSbZZuVbf2tP6Hh/mXTcK7WEaQqk
vHjlk0A+FXwX77TfQXVv4RyMlvzWWsGxbTRANhV7DwEar3XnEPKE1Aq2o6fnqgUq
0TrxlvmbEXkYflvMYdqGOyPxC8U3Bk6z5/1qhFX/rL2XJtCavYvS8qozKM6hps5C
rtzT3P+A97HujKXvIQpYE8zVlWNoSV4lF90xYBV5ysE7lvLvvJpsRl0OpcHVFKqv
ahoWj7Dp5HhYbW53NEiC5qLqduIm1E7asflqnmTybE020wWf2BrHfnrTI2ysE0of
wqwVrYADzX7tQAEP0DYxcaGQIJ3a8ElC0ihKKNoQW1mHUQeVrgbB60EDffsbNWR0
zsFUF61DUaz+9qWncEEIYXUiWAhlLlZmix0NfpVqPjizpEqL7uEIekSqLhRPEHBH
lbOKEBXmGi46LZMTgCZKZeokYcvnJXrdk6EcBEHbiV+B7sYZEijyOD8eJ7MUkWAs
KlEkDsrbPVKJssAphndXNAYTH7HppVdxaBUQWUAKW5cdzPLwrI4VXIWWrCMrqSZT
ZA22ncFZg9JnwI2DOKEkUTt4ij8vEf4UDZMrWpp8bzyzSVVepquEJ/M4sNT4FzYe
UAf7lY0JYdqd76si6cdM+IRlmeneTpth9mSAzUtOsTP/499Bctur24EgzgRSIwU8
RQd9/lbs/OM4fiK4VK0L+FfAAVhAXIH6bnHxwuPTtTtwgUKeJPs2hwFzgIndev7Q
uMeyPrxaQJ/5uDvmQk2qLmtl87ODwV7iuc3l0j4HBiVapOSpgDdLoa+aS5wzxSYA
+lf53mPkDZd2JAD5xwvwj4jSzQPOwxI/LtrAQYorUjSk7g2s5ai5DZv62twQPUho
TihuXqqs16ppbWH2TQwXru8i63nxuQS/SieuqCs/sU6wGtJOJB4szXOQA5nnyw47
TywpmQAOVp+y2WZRJanjfEo318Pz8h0QqKvGJM2wvmtX2r55EPlBO4kLSs4H9wYh
I2hTU/VQp1IY6MhRPkYv7HVkDXaBAa6O/D5dc0P8eSQx9+wzLLWNB1q1HkGkAaIC
XeCRseuA411wMRUQFFwJidnrjihkVbPOESLnjKX19hERSvN11EzI0ydrSNcpZLXt
BfnR8yFAK9E1JimmRAtmbFXPWHnvfsMqj7r2ap62USyxSMn2JSb3+aGnD0EjWtAt
2OOK5GWY7oEZYr/oi5TX643ty2YtZotkmG2AZMYmVgOuke/QkxKT4z2oF04NWTNr
EY/a0LbO48X0IxdB1R058ZiaA854LIny0O0hurQABZUbvpZaEEKcB9uWtgZZ2dq9
u/MuNaDTgUSM/63kqHy/5ECkUhjHUQfllPj3ZzAnwiBtu/UR/unhvwvt7cmE0OEQ
Ai7NUa08NmiGOqb3y6VdrJ5hC+jYDaF5z+RgfLl8IxvNkEcQYOH200fJJ/Lf5Hgu
ALzyyDicqC0rmHIw3L2uGKSb31VQpalTYIhrsfWzuOOFI8vI6Ri/YqJV3knlkTGZ
AdCqzVmYevIhWlGnpaKtGU0DTx8RQYwsu0jaPdTR917/Co70a/HhBEpec8SK2hKN
XUD+INx2O2RjUGrMeFUWytblMgkR7U7FGAW2qfkSv8EDjxDgY5sh8Gc+rfck9V+X
0euAYqvmDT/LDbpNj8iGWPgLtOGJ+cn5chKsIr0ygo8CgLcDbuLijzxuohVw9f0I
wQ8ZxosVZjM13fQXcYIUOQS/5j5PPHwA2J40OjvLnOzPXnoOeji6LSyuCPPaTuGE
9pzzzwu1JjlqKWOmfx1ezxn6hCG/74P4kCDUA3rYzb70BlE5zlL4rsHzWiuAZgEv
80gx3byOzAuKz7PMCbnxy9QdrRKPbE0IRz6a3+SblrO1vr6t8y1YWq8KJ88Oiqsl
XQiy0BG/5pduPerxzet3BBEvasOUZ02Y6Ejwzd288XyLoxEeGMqRfazu/wE5d8Gu
XgSu5E43EQNid5DksClshUiNggJlU57AUViehwnOpFuDSavBmIBVL4p0MGfetmGa
ILuDhfReo8u4EtqyVaqzTQdMQTjsCvH87oM2UMny/vW7vYnt0Dh+KzljdK0H1i+u
ZQQiLcxUZBVnaWgVsFZEKheyQ03OMIps19o5zczYwNlHf+L0igbSHkwkbDO3ima3
MB3/Go1wRUwB8pqvFO8F6Mw3HQ7ULjSeXiNfQ/tJelidPgbYJG7lSNuWDQW5e+xv
KFwhej0/Wc6K4EJdx4p+hBGoACzzue5ZasCQHF/3Wy/WWgBar3rpBdZovm7frwvN
I6VocYKYsbzkr7xsp2KWk/1H1Wde+5DAKMCwlaWrnaupAeL096d3ks3dHTt6hZ1F
5biSd5zWLT79x5iiKLG10NK/zX87tqnbN7QGqo7Vh6cgkUqshMKNRnaI41tTWKGq
QZfC+XzoeQQr5WC9uHU025l7QuVtnMO8e7dF01LCouUI3HTgAJo03vmKobO8GWEI
FSyXmTkeiMEKdjjy9v43Y+HwPLGoKTqLtnM9pOuA9aGotzklh0i3MdoJZ5agpFqd
A63y8g3MdR6WJiRYj2Ct16D8oHBqR85CS8jEQFW1eHZVjm0OsGC4cVJbCUL6iDE8
Rvx1VfEGtcfDliTC70o4MNlaMKimBQnvRUqK6lVIZrPKCO+Mi98zNNU0MRpHYQEf
QG3I5NLhZfIJt66nvexH7kzWYRqApLSAhV6fPdjGX/rd/X7FzDNf0XPpzW1vA50n
Wi2Oeslh0FzQDFDNqQBUn5pt9YEAmyJtGh+P5exwbhVrKUp+Rkwr2L2k3E8LtlhN
wDY9hExI8rRhPTjvPx46hlj5TfvEK+jollnHE4c2hIvsyXrLIkI5bupjQ6Mtlm/M
I9t5IZKgE7C7HPUsAzSPDAqA3R5cW7bcXC6ANxHM9S8DJIG2eU+EynJ/GhOqN+5c
rf2uLUz9v7zDkOOhQoY7HxsHLkiyJqbS6BpMdJaEOwK+5I+s5ps/IbNdG85hr7jE
2WFc9i+sb+t8kjVUz3vQQi24x0Qg+CIP7Q9AosLL28QIxpzdRPKCr8nGatosDog8
tsYfXAJBq+k+NnXw2fQzPR5+q9nnd9oc0XLEZ9kzN8XNuoVCNZqkQy6WMkOJoVM+
QSOGR+gJ8Cfos6sj+0MtSQY8M5/o3P6sJxba/incdmHTePvcPbJT5dRix+hTVhWi
u7iVjXL3UYW6EuETxqTWFa86ePSulrMHy25mMQhiiix+t95Q3DjnJq30KDvG9WqH
H7AkyHqGYGkIsxGgfS2dLAE7aUaEctxZ2nfE51FQPMg4NJ1e4qqO86IqOG4ZG2kp
Sme929z+D64JUbph78MGjeCZ+ziOhZtEdcHq1659olfedJ2Tdf2XR+crEcXrKyoT
H3IqWiaMttuiej7pwuQJnrB4zY5axT4knjyptm5Pmo0J1dh90ocU/FdgySt+DPX9
4+HWxT4pR2QSIKYyNCfV0090tQza/XzkGsbsd0MP23e68/1m/d4nltcyChAU8o4/
L7waUc6B/iKFrh24Qrn0FiBYtOLIByQVFUPXpO+XFt/7jlmHcczOLZ+Y8Nj5Xaf9
cjU8Fut+YcYTiXErF67Nc6fFrI6+4TmlmMtSCtJK5II/sDRkSsyIR0DUtQ8vlhyN
zYNxXJKX71shbGkoBOz9GFrT0dBl9Vf0cMixH7poDPfYpyp6be8hj9S3xABU8aEw
dO8RWgsV9Sc11D1hA4wGkulHGTNFsonVDjcwrmULzdSpo1anUqWLtxiKa0dRLJfu
97fETXA8UqbmouhbwPxhVSTIlGyv/JwTW53UEiKHYa3aH/gNYLP+W+X8Prmy8Mlw
zJt/6r4mw8D/NXmQ0HFDcRfgTdDvtR2qoWGt7sGXyk5SUHlgyhxG9vgqcWaOadJI
YbS8YOdr+iCDITQbJw/b3vcR8hH4Cu3uVH4l6X8R4S/SPpa+3JuOhIAOwxEK0NDD
GXiU449HEKMrlh53743+wrL/ggFgvFDwtkPiLUuRcitfYjuOLKsI0lqXywxNfQZv
13+AWxWeo+GRFY7T/LgxXqW6CZrhtiujpcVvPAliq2DTTmkt8okxt13Y/QbFLQ8O
uVc2a1r6Mc2Nn59PdFBYG3DBbGEfySqNWZ5bc4soRZHTCY+3T6lfhmBlpgZGbECp
VUxRhkPySKxIrtzxNgjyfvJ1xOQ4VKVIJghH89nYaZ895fpZzd0/oNWrw47vf/cg
CXLVjDrvcZuCuM2GQRLKshIJl1VzaxlvGTvShV4MhnzRI8Xauqpo5UysV668mIYN
UgCVMl5AU2BsopDufBlEixyx3eTbNTAyX3hC6nhxFHpidOlvOAFqYx0hgB7F/k22
tMXwo3vbmxUmF/LD7zcDFA0yo2B5k1fNgO/BELrxVSJ4bqmXCaY0Yha9Y4u9uxpj
rKWbMmVAW7+a7Kf34PqU5yT+75K4TfMgwqoMPh17SXcGTpmJOXnarV0wkyrJsxVB
LW6xrkGSN7H9pKt2VWhEbcLRGIe5qberoAzoqTXifBrb/KZyv41lRqMCHiFALlzo
ugWmKm17ldtqLcHp8iKmBxlEp9hBV8SnGxvtuy0WULv5kOdQg8+rQB9PabDqYNso
f4yZTEsLcAUSp30bYqpOmtcODX3rRz2fk4dqUgqquYCW66/hEPoIao3Ls5dZ9rNU
R6Lut3l31gRCV4ZNtnwcs9r2k42ZaGz5rT1L9aqPa+RXTZ4FmujUJkcsBU3L5TSM
2vcJLO6oh4frQiRmxerYI+jHy3OB5fuTFzbRcOVHpEI7EbOtXESoVuDOviBo3sBF
Kf4/amfmdITLWJYRmzvz1fwcez/rfWsJ+hc799gxGEp1gP352uNcjgqo9faqHfZa
Y90bJqXOLpfb9URWWPNqBiryE4HDc6jkqOP8XWO4t0YciObyZi8xr/fRRCZNJogj
B97I2w7S4KcLPEA3oPizcZlzep9shBsRXLzu2YRnQ8k0xJO4b3AlYLvD6hwg/ZRF
5Wg8nJykVkwOeTVWs/Rr+qG0+EKc6mVUMeDYmSOKMSQpK41rzyTxPlpLwwg06It3
pdaOax9lIK3C0ChSHpUoeQYgpBCTUeUjt7Hcz57tmCVJS19+epdygYDPWv4q59oX
lRBMsEuB+waxN+2qGC8faMmKB0x+dImHa+ShVsPgHkEb7Qtw+Ewfsj1UHp4sN4Sk
WpPnRRP1e0F7FO+jdyFFzkjE4dIR9DV6sGiKM+fGr5oeeFqq7NkzyRaDe5KK0lSC
XcusYIyDhdNboAh73atWbsMnv8tr+dB3Ax7Up+x4jbgyuGb2MRIx1jRilh/Q/yyX
Dzw2xg850tZ/p1Aakr421NTN11jOM/5bOSnmCS1KbGqewA0GkSPMXJz6V3S5aN9M
awZ5FxjPQDZ/eJwmscAaECl2zVjdBuzZkShP9NFsNtTo0aGg2uOTSSz/XCdPng4O
6a4Lk8/dZPNHJ+4cbec/x5MS9hDK/E1D3q0v+0Grd2Bsl5a/lUkDxzENEBT0Y8TE
oqFT0hsKpnCIjJXcBBc53R3vK8nUkW01hlL4omFsvx63yJSWx5pLf5mGgFRAk6wT
CvCdbchyw4km6NT9Mp8jBVmo9qBeRGOCVpXccxBtOe+9wVGuobvQtkF5gRltfszK
Ye8u3zcKPnwF3I6JZBf5qFc/ohOvzAMOxicWS00zKXUqA6DmIzbd1uiHj0C0G07I
bQXsuAoHySrf/uzXkk0LafCrc3uJqmSQOsRgOucDpy0/rM/SRMlHpb7aiLbHzfEa
26Ofc7l+NTZrylZqNKQ820E7u0XGYjs9IbCWBD+KZ4DghKgPGSvk+yy2kQH0sYwz
sJHSAYl4dJYaaH8hpSOYqV1X347v7wRry64SZT/sHKxXp2PXb1Ya1fHZXIPYqIoU
lYu3ACP5nBzQwu4PhD43rzJfMi/CKTLJZik+8V92nsnJjCS6mApBJuWxsZesrCa+
Z/la3qUeCHIBupbjsOr6Jzm4q2CP4vSVMvZ51KLumt1eIav1aGYORevdQuXm1+WR
YfCjm8nJvwTtHkcakvzTLz04OqgyTsCnF/EReYcTP+HQm3t647hENQEpnblC6pZ7
pQf0CPbtq83ZwFKOv8udzOEmcdDCzJ5KrsXlbJHrJbgnS1phOhQ08sf5ds6X64oN
hQ/vescQvTDAd8a90FtpE76Szc3Qb/+0Waj5+gVR1P84KLBKiYPZWlYNvwhh5nrB
De2cL+aDp9qyqWSwziGHUlPC6T0NRNGNDvDWUSGdq0/BnfARenSavMlLWmRIqZD2
yrRx/OgdCQoQBhABe7EFQIS8nikZ3h5px8tYVT8yyaPcI3XmxGCzi4aIdDcTWutC
HCzmhxprAZV0A1nl3KL21Njj3aoMYhkEpQvLFMhPltCCZ2vXZP4/wfqy15mf95WJ
NFnJsuREkXm7GiFIXgVLOHgUMPSFJ2D3wUxgRH+ZVw7w6PCOuOp2pMNPcjpS2hMZ
LEeP8C9/nEtVGVB64m1hTj6+ktVXnhDbn/s36xSiCvNm4rCQ4FJ+HayHZF42NCew
biU1LDch0bfEEwaeGphWLVeddz7L25/GX0OdIYpSGPcakNyKoDUokVno9Mno8RTV
vmb6wna8SX4ecVst5nGw4ZbreHe5SNr7HEi7Px7UaGFQu+pLTuEMNLEZcflLT2R/
70pwNGgylm0TvRN4D74+lyMvCR+2HPzD9VTcdg9glKqvrtOnTwp2G4ktUkmqOvzy
eP4q4JavIzL+pzXt9rB1YrHwTTeVVUrCXkeGux7kCjgw2jIUH8TiSbvgCNkdcJFw
vw4jlPzNWGLj4iVjbO1qMoRiP+1QIlV+8RempQHMNGHdEvnhVtNjLO7T6hySDUOg
rsUppGvFGWbCbBlvr5xDX8WtKlQ/aGPtV3P3TMgF/xUtcvsCLKe74cCHNkLjjUk7
+PCPIMN3CFOpjd0PuonxG+5Z8lvn1ZwaBDJagmhuWNkwEb26buAREcQi6wbQp2or
mQoFpNHste/ElnDyY27YKcYsHYTDmIKAHHjNjkTuaE5hkGy2Hhi3KH2aBv2AdYcT
99t5Et+nEVx2/frrdFWXQHX3DgvqopbHx4d3FS6ejY1k+Q2jR/62Wji3Xtvj7cVq
E663eOTe6Skhgj0jLQi9qlGs0/69usysWnnDWjKHUuNw0kfKJhFPucKzJYF/9j/o
jveTAbGNmeWtKj0JuT5YlLjdIh5nFMMP7AJ7Ps46ng28YxCAWauLfDuPlANVEYtm
CSyATSYDdWYdlPH+afooYy7UI/fFgGOyljDdVc+aS4G3bFCRZCcVFtVH5an9hHuQ
2QXfliDMSWpyY1Fb+4FUuzOUEM750p7in7/BtC3C1jkv9xAGG5yLK2lnKQeZtSap
J+YxjZCsANnNn9Xj8yzlb6pBnmW1sAy1q1mv545ESV672HeLKjQUbNzOZl95yaBP
SCwwRQ6IkgCBhY7rb4ANYKUE2RaT69xLQwhuR/1bdXEa0/k9UELvpjc+VUNClPvH
yHOTD4aO7vVOaxiLXR748hTlLvaokqkHRC64fSh7nMp3j071ziEOfQGQOHEZxGMy
/hrhfrlbYTAjLNcgCjYzr6WTwLZwVkV2mqQo6FVcfYAQZBIAZk3lK9MHgJqpm7nb
HohjR4WNU848b+rxZwdN5RxA41eSp7FZEXMUrwJUb+2o2KtsiyPyQW07f8rrMdkb
k3SFB9+TACzhqIbzKNGZhdpnYZUUvyzrDZ1j36NEssimSEfHFgR0+zWmExuUOcZ5
T146rVfEETAw7M7b0ABGNUpZXiB19A597+fY5r7heorY6yHCxgTm1OTYUYob5V6f
WthWOlMtzh4VBOp92jYWGA74Gx/XfbOVSo9FLjM3d1xL/X4vBk6Pr4nN6eD82tg8
i/mDm1NXwkjNpjEfRFuzr4p8/SHHihBgf3oL8U4M5wEHthPOvSUysI5qBTg1+4GU
l8hZMxZCkGwh+QtQX98IJPi5P/8gm71AMKd1O7CKl0d/zbR3LiPp3nsLkYvCkhU/
MSyeZ/l63MR783z1SV1fHMD+pUujx96jL51QV9xbE+kONqD06gd4x1gFQhcg6zpk
nBBj6Sigj9Y23hglM6D+dP/LEObZT08dO8gKQ5e/awCjGNMErGB5j2P7qS1T95Gt
aNYJliHTXiOTtaRvTRjM1x2P8pb/R9P9BHz/WGyC2Lqd8jjdiLMCv3pvslfhsMQh
r6ORv7+nJ47V16ClL7OUscwY/v0s85UYzgLVk2tRrLJTGvBt7z6AbVfHigDSkCKk
kgVr7gZytSTvaxDmCuyayZxd4zK2XVDO9ytMlNzibOTy//6A1KsKZrxutQEHbDvz
LU3ddRuUAwADRr9qSIrErO5oljasR9fvx5Px5hAkKkRbaFamgTzX5qsGAofsos7F
Ep0JqhjkL6jNpOoXP/am/9jscM4PmBtztQG9IpuEPbg1RKV/3fwO/y53scuhUHzV
ng2277mS4dvrS3w1j1PSuPK2izM5B+wTsp61iY91PlCxdbPVIi4sBorAjpxfGkd1
8bmLXalUlQ9XUxJL8AUu7E1MatJDry3Ak6LPvWfqTTtBhN7KZ9mj7tFLx8YZd2Qh
ZbwQr7eqY5cct+mlFwVfAIatT+zn0LGInomlu9nOpL+ydAgF2XUhI0LuMSd+R85m
7c+w9GTvmEQUN4bq4fwLYoDumKAbbQa/SK+0Isv0vVq9XOumw2VFRSPW1Z5VFX0A
BuhU8YrrA9jRZOkFwZmKstoVljJidkgLzyhqRXrZLX5agaZokb+wHk8jXGsEvBLm
52ps05SZt2fvFzjUbmwpe1drjWHTZ2GeJn+5+UuDzFsJ3imBc1BlmzEfSxDBkpbY
gFzhRbnV6sIaRNbEbLB0G/OeeoMFjQkOgY8ng1EMWSDicDN/YMz8TUSlZ7+zatbI
NHrzfh5Qk3dqyOHDOi72hLRGkP0iq8LXOrFPoTi8/OAXtF2tZLT4YH+zXY6bQwFj
j0PR7GosSFdoqkmrClR+AivGjY2yAXAXcAPKlsV5mqYcV7ibv6Z1giCJZAnEeWlK
hiw7D5osE7Mvl8dD1GtTeI22+Pei3v1Kx/R6jEoifc+fgccc1cLR1eKyAlRZPTTH
ZgiGtjhZEgmQBFGVJJjT4V6eYM8eB91sN+CZI89eQzU4o3ktKXucq8jHuQGgqCzh
TCxhrEowIXglBqWdlkPrzA4/HMEeRzBCTMGMoy9Fwbas8xHPulCoz4gPIsPJdf6X
yUWj/mgiPOENOYX58Lei6IJ7jswa02fkxfRLDprPGjqq7+tUoqs3MPLNgcsYr8t/
bhPDWpNLodAp8NP3fce20+IKZppMfQOTBC1+a/ZmrU3STYOwaraCndRgQsbdtY8C
1/nmcFTlzDoPJkAxXPb+Lo2nPgQzpbPIwsQK80w2XPd2wnpokZU2iIaXqlEl7mML
Q/QmKkx9pcXswqvlx73mIGLi96QNO5vqYGoNon977M6AApl2YUmh/QzfXZeMr9Ly
d1gILCw6r1rNwUp0J7yvKnbr2GFIQDlNwM1azODh2wvtKKhVUoKlMr73DxTFTl7O
53EBRI0UgsKcjb4PdRwUTf6qnzORra1ZNU7mcdhqCJSisBR0UK5euKKf4fFq9tBD
0F3rvcGEUWmQ/6nOUcXsAK3asvMufzPAt251B90bKAi9m0DR5bJlBnF7ro4ddgO/
NxX/rSY07CHUwloBM7F8c9IE6e4xZyo8EWRKPD+5AfGU1dfvuOreX+akBFsDLa6y
Ulea10t4MGKaUn0hZnN8e0kcWnd01HNFU3fH+Ngag+ocsP84LJdSkOmyLItKhXve
WSg3SYq4AKRuvkxSraNPc+0IrkUl5SBQe9Asl0s3EFf9bJmwLchzUi+KtrivjPkj
G+YHUujCjhLvoCh8psu9t6DfkVq7bmIE505h7i+6assIyPlpCuRoexV7Rk1RS7Nf
8G0XsG4GVzV2q9Cp4DIOR0F9U//eCuo1PbIWVCVwA4wHZ7qkQsJP3L3MWWSHEHyw
Fkso9Kl7IN0H3wsh1qviZ/Qv2Vc8KOZvquEUtqTMDoJ9DOdSOHBQGEO1Ur16v5QH
7zddn8pWFhQ7aYlGwR8uUgcw1lyqR25p06K0FEFq4e1xgPy0BxnenseHOSl3TGRr
x3ZQP3rrvxD1IR2KNMF7XSywM3InYwUjX9lzLSxM7+N7Kyle6KDCXudOCDUVXZg9
K1NPAPxz/JDyjBWLBXJFH3Z6w/I5KHIWvXVa1gUJIXFOci7L/bTPSn0e8TnEzyjR
11VEPQU7vtUBbML1ZI4o8E+/dHL80B63GCUHDQolP8pUg49yUuLL7yUo09PuAn5w
juA5WyYMtu/XZR/3Bp0WVX2T0D6nO7GgEOEj8YzY0caeThSBZu4qbRYWvOHMkRbH
UH0hM0Vp8uNbta3jc8OjCcIa8sBwyhONR3GL5pUIE737ekWYNzF3T+aQn9LznWDK
HM3FUC6nXmgSw/suFuXWPyhrPZ5UA05sXuCu3LSl2SsnINKNMX+wQrTCTCLvSG+Y
0EgW73H8oMCNyAqFtSHIdR5doQBsuVWsHBD7Q+RZ0LaNY0G0xNtocL7sMTRYa3gW
l6mBfFzMDtOUSmSd01KCPlvuJYQ8KNeH/bfpE7RmYQwypocV3/eZJPnvzcYvEgmB
Xq2yhr+xH8wPBTJ4nJeaTZ1BFqWwf1L76q5U5VQTj4ffdrn9V3enkb4got7xF3Yv
Ks30SDt1wz1iG1OkTCZr6EvISSgAsCYBthqfzP0ovhw1p1tvv+6mi3NSZ1AQMNmb
EAAF61Lh2lSTm+CUUqxsF3lLipqX04/qNDjhtV7hoKPUCCpn2QUQP3R9PRlgJj7I
paFBXzx5hGeTiFVK4pSGwijD9O3TSKR7ajzpPNrsMgmxLIygIh3P3KAw5Pz4ZySl
6QT1pK49+P+6zut8ul9GyS9Ig4YbLG0QIYdzw0g8dut2b3Q9FXwaeEFKwx1kjGsE
6lSfCAf7xjl3cyZ2Db1mhpkycWVIrpTmgCBTEI5K9Oq8LblKzXHOG9Xz60E9Tp5D
NW+b7vLA80P3InQFfP2V+RfVZQU4/gWlB+J+HoQs3dKoOt/17dyKap5UT+4lASri
HRse5wHWvaoaW0/xrxR9fzSP6tOInsQynVjJ44AZ6FAn6O0z0f9HGBPYn0N9GSAy
jfgQi9cBt3Ud2o3k9oduBZokoxG3qkhxJYORACy7cJr9TRdMGHIxlEO0EmT1rCyV
NI3o0plHEFsB34VMXyMVkRzDpP09bLIVwjsFNUDJTRjWOwLghevqsj56xlF1s5FT
hRh4XRLyFU5TQ89cw6GAEt9/Kvj1CUicAFxGWTy4fG7Ltl2sobKqHIVxJPCPFPaM
Cbk5qPvIuWVqdn14fZWuFDHyab7jLQDVNwI5BUxAXbv1dFlx6UtU6YIlRYta5ac8
ecXiutYcd9dpuJOWcBSa3e4jm58q/KPG+99me9QOO/Q/YJ24am20VqIt8CmVa0h5
DKAfw8wvuuv6IKXOsgWlPolL+lhAdnE4B6FI1xBGd/0dnVyq2ttiLS7A8szDD51z
ksOokJvDak9txMeSRd0fhtuC98PxBZNofb3RljTUU9RNCdZuhywWn+Gtvpqaj4Rq
ZXAMZbSaO0BB3CbEn8qnjN+RFo7K1WceT0i3sQ0aEXqM+e2ZQL4SZ6/pIxZ+bLNk
`protect END_PROTECTED
