`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FysoPsZK8udBGc1MmaKXyhgeK4o3DUV+pFuaFTd8YXU0q05sM1fLpDunHsqyHmsi
BZ6iUxFQ0V4uqH++gpAJc2lvs4yhWF1Sx0+umRdcUymdN1dE4pFdlY+/eO2BCRR9
RUSP3tHngqmh/0ZNUfPLFn88qHi3SC+Ca5Uptjg+5f7oAfeVQs9BNvKsgxNJc6Cx
pcAtx5pOVKbd9lMGEHMQv12hXE+xSY9MWG+uNzHa9PIqO4cihuS+5P9rqkZRIYAT
gKnJBB7HYcqOlSCVaep9XjCMdH8rF1ujP/9Rquh77P5GgU7GJHEeUSAreKQuALHu
ou+0wXJ82HLKZ4SMAOXffWaYgXwsmbyPqNlbBs9xCJ3drSp3WK0lXD/IKvtU1loa
SKQlWGWch1xN5NAEGvwUO2nWhqg5MU2T2q4xJWNybs6EfEd0sqz3mfUJbavpCY73
zsuVX4zv4iv+VM8TLPfnE+oYBn/hFRsYr0tzJPDMFrmiYr8c7gitg5apy6ttZpMh
+XpNLf8BnPXuwL/5VoAwiyET7+5QCTeZPSqJSivajQ5DIIeL/y0P0x0Kccb9hmvN
3LdrS3qmmeX5GCFGlmz6tU3GVcVCnqzY4dLKuCPHro+tzvk5vcb/ZZjnAVe3BBcm
bI6eE3Ymr3Ta9i5/0E+zz5SKd7AVaAjOsfAlC9u2Ygo/tSKJW23iNvM37cb3xgtR
`protect END_PROTECTED
