`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1e3JYk6Hw3nh3NnMG9tQnJH+5sVdkhp86JaflVjEi3c/mvsNhp2EsZMoKktbKQ+W
0VCTZFEC7G8PAeR6NuDCpRj1db3rv5PTIRBzCFZFZqDUGOdIjbbdvxt4VNqbVa6J
LrVBq0YEcSdhEs/LWazxDdjcAq68k6k+EEZIiVzVPjACfVM3mmfFtej9kJjPbr+M
wAyxORst2dwk644JRHM85niblVEPOi2KD4sJfotSJ9WKaiRGPcxJufbNySRk3iQ/
sWxqiasEczmXts2BUBMAI3OJSJ0D+fTLOZp1JMdJxiClOQaeEAgawdC+UHf7uLp2
/a9/m2GKuKUzOitWVUQYoyATKDjIHhGNyGbTjFrC4XtgxtcZkrUv0hQFNQZnpfz2
p46nj+/1tSsMcfEqPEvnb0LX1iPJ8Xu8QXJSqIotiE+I1Tx7Yyydy9voljcDqAM7
BSkq+KagEx096dT37j2WHLOVGQajDhQg1FoV0+8widmPCClnt74tTq2y1YhTMWMG
tqWIp6vCN692gl56pbHfjsLiHGQEvrBR9A27QIaIR9ykKi5eVoBqYOo9CB0W5ALx
rPb6LNkkLWii8uDnaEzneaBTxQakOLn20oZsprA72v5Lrx6U8zwTm51cmJiHHULS
bDDPjzzcap91oVCRE15QMGe7Tv51NEXCf8AYMwFVEdNOhY/8giICsr1ITyoK/Qgh
8B/h2Fa9wy05FKU1b8TOErFjDtpTZ7bRiMY2lN3egl+IBXmkR1O3fQVoUXwoymZr
JJw82If+0JG+BFG8aurExKpee4k67BN4Rydv7lm539fQlpMyhqDoJWnWsawG5e+U
3RyRPff9cDw4Lzm9ZbJMKtlWUK1QXN4OseaMSdUk2sVXs8LvW7dKAFcNJqXxBJFk
emy7/GsIYyojgHahC514BhhOmi8lj92oQHnLfsQUWqMEsALEqgBBqcCMqPgUP8vw
tW1ZLH6slYXbVSi/u+IZqxI8ekP4GMAJklEPNHNCqcGrdeL59iBAYsbKFmou2M0W
GUr+RDuOHCZVgJ2efJoQ+lulPo5Guxjc9KyHZdOQtxV5+/yfgn4lCfpaBm5ZbAsx
1dH6yvonIimt0+U7qF2cQTaPWhkSZchTNFto9RMr4+F6MwzGHrtxBcHMhWBCYcv0
5oBaHyXpbGxfqCw9K3/bnuXQRNJ5P1CcxKRDTU/CvA6eZAleHwUkuWT7Xg5QHrUK
Azyhv6AOp7iB0iLRObfckHOj1PfbMEeAGu+tCX11D7SfhF6GNIAwmLn/KMtSWv2n
JYQGifJwXT7B06rYBUXllT+MS5npBJMdedOx+OPpjdnCtVM+rAz4CYSpcLUihYtf
CVcgGZQUofGKogb7x/oOnJYHNGuaCI7PXyCrNiqeUCBBWF/ooB+8BRYPZqOc172Y
fN3ttnP8YgOkJ70hQ2HSFC34Lz13KDmMSSKRIOECCqF1zwQltvqkCtHdY8S3fs1c
cOhZA2b+Hvd56ZLykSNywltIkQvo3S4unnTkGdbcBT7xmKxpzoJnoebrBxXglkmw
OHfS+LuhXb2cT/R08APfE8D2WOm3QOUNU5YQW8FSdYsfX+w1QfCL4NoP+5lQ4opm
D1+Awlwmla9pCjbMtb7SfUhKnPNy74/AwjOBfPYMyXXatYjoEHxyB9paSYknXMgA
9SlLcGy2bbk0yuWnpmz0bk+N0D0ByK/oz5zekPBvBjeFvZdPgk+YBNC46Jq3slKV
phJIIgHuEYzef9rIReuR/hBPtdY4/+4EZn9iAsfUzGs0qplLl8GMsVnAvF1m/aAF
LgGohhMid2ah4qJf0gXBxwdOS67uy9FcZr3HBLsEy7W23LTuUoQlz810kENSVVw1
JcO40E9hsIcZvdDnLO+ja8dl/c7NOBiYfSagt49Et9rFoErUPcuIUV6ztjxqvhcn
Rb6/IcsfbRY+cOyksKKFHWZWKCKxsSld1vpOIf1bN5l41sSu106jQ8KbdMuN2b05
TCbRqcsIrrEF7va3C7cT3Ml/n8spUmF/uhfWJBDFqFwyR7HwR+UJsC6gHq+6KIw6
UvNlFx8nZpe7ZGPaMiQ3EcGzqhzO/aDFK0Inw8eyufe8qarzXpKbvXgHaTZM0K0Y
bQe7pfWpjtoBWu4YIBYwqLJfqJltXtOpPHL/wDkEchWPJT2BfJpgaFmo5Z1kgFV1
Ab8iQaJ6PbmX7OQ0c0Y/sZqa2g8sMtzvdRbwTOcJWX1WfjG6N8FCw/9w/LUJVYKO
cZgujoc8EujQn3Enad95/2+qmauY9/ug7GpPH9DTBVamI+8ueFIZS7TWttg+01/p
NKtvR6GoFeKDo1abE4z9EpsmuIcNihQpFoXLx6yG1AyUYQwRFwj6BLDLcatX0qxZ
gX3aEQHvhqA2KeOpOucyNxHqDFD2JFAjL9xsKgEvKmbWYaOvBHBD3D5u4dBIN+Mt
EWnJQAmDC/jSfpgsD8gK7hzycEs4E2934czkUrbZ7zfH4GCNd19x8SkoX618P1Lr
4VhuJcwEZ2XKhpgvtb99QCv95fVoXW9X1QVUKQg5zQdht5AOvwZ2W8jM/Bc3EAoi
mEnqqJ0mJePGr+PHXAxVpjBiqLEytPz7LJzCumyanGOVivXsCU+WTcguz6JTbzbL
aiwnC+sdvNJDnF/r4EeGTNAXOL7m/n23xU4abOfpbADWxvGzPpxfg7G8wulRVViJ
Lrkxl8x1lP1/BfObuMfiJ2KT59Wf6/5ZyFeCeOUMpI4U+xPoZo5yWcCv07jancpB
NWsqZe9WFaRgKzrX27eaZSc9Oam6WP/LPl7hyJtwAYIxM3CQMla1Nbnl5/3X7U2T
1dLYwslksCNpjqCaW9Xk6Xtf2fi9Q9lpuHGEQETurdw2uQ5r5cYl2N61/rGMiCu3
4mfVScgt9XDNfK7qly77sBqvfWAWgiPj2AsHewB9sgL1I9y8UQYHy6v2Km6IfFLU
vGI5oeJSRzx3jliGLYXpfhKHg6uDON/GIUPeWdniNSaqxZ1n+uE5GYrstZMtk0Km
QlAU6+/v3X7i8jg0AzfL1dqnFDK1wIlGstpTGehiVegChXIQRE70DM0JiBz28/1p
oA59aGzH1SmzG3wv0D8lEZOs6jAllOsYOhjt7ZVpG6k=
`protect END_PROTECTED
