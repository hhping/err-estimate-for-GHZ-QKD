`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YkROS8BogFg5+UMhgDE2iR3tSGFvQUGTJThkuN3p/AvLESpNhBC8c2ouT/ZHBhO7
DO9LN82uAjjhOvHNxyrruEpsCioA25oKKQtZ8aLu/SE9pLNOvLtW5M/eAhfhSsGx
MbBFzoSmShy7WlPsy74fQ7cWo7sygbjkxYyb123W5IY=
`protect END_PROTECTED
