`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q0Dl8oABis/ZInEEsOptXZvl0rFeNiy/fb3BUZXwPEMOdsiFbtSuxQf7Na3BPrCY
ihbcRJikZi2PWdhs9MxiIjFQnTAEw1Q3/nhh19Ig6SIS/bWQjjBj9teGVA67P3ea
nZvJ/ZZ9l/R66HpItapqljg5MA1EKpikx5tI+I9ckFLJQuHyVSe9gxQFpO/31UgM
vcBcsZKrhkbQqmHfeLt7ozso9CYMmBR6nR18N8kuZIuD5gIZ4E1EkxDSi6eK0QlI
BwxHaJzZzP+1zaAgTQQj9vLAZiHTnfCrtxxaBHd/W3PcDrwy4ujt9N9j68Rr7zDN
BuVG0SGy1FUlTIA1+YpIjskl4Pp0CmwoUW0XPIWh6Zc52zHQdHqxgBJ1mEvWrVw2
potU1gNwIsNPEoK/TKhT8dWeYmZux0Eue1DVJR46vLQPy8eCgjcHWgUhsxj1HngE
hIBfgHSgZq2lsYh7HhOCfOx0FSofFjxosqjrB2xhVtLPZfonr3DZJOLDOuTFkSK/
cfhbxvwZjuDz1T0ITRx8dDChvolQwZ/klGu3W12FHJ0tB2RNJ6/riUnsy0N+gSOY
K7K8rdl7WxFzwe2Fz0es3ih+z5WNp9HP7RKYUTRWvZnl3dJ5X68KKQCMRAZwoHuJ
iO4xb/OEu/cwGoHFkpy7oml172O8uYCZi1spECb7JiBFqcTw/EoKYG5JSC6pI7vA
0ceZDLzKCc8xbYBF5pVu0r20UIJH4tVNIWaZyVFfVL9PbLODNC6HzE53nygKl31k
GOjzY2oG59Q9eW0EZDZqjfTRBSWqh3QxgrEcz1R1V6VYGOiIK8jvcwuc8QXbdb98
1hUeYbP/D4HOc6ArRpXSynNMr9HmADW3L2QRBY/F1gu1aL/N3yuYFyFetdV6Amsy
gDUScBkmzUOnHThLipbJg2j6mAF2uSiaQZAZsw7AsoY=
`protect END_PROTECTED
