`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S0xLNjkED6DqcrYAKnq1mBXxWufS2GEcrNMkxn4kToCMQqMcPqmFamU5Te9rG45t
YKO2q9VXJfo0Msyl03NHSe0/Mu7od4Fk3cRWZxumZLuVdc9iEZzgRdBtvb/zI8YH
gzawPpFdwutn7g7mAOe0DOl0o/u3lIIB9Fr7H7LasiHQPYw7fuYkNbcvI+L9D+/H
pzaR+bUdLLSupHrPvoMFfr5OjTPZdc92LZASI9AoWaTvrXZd6y7dBCEgMvatvuc3
6Q/7WLnVyCHSPZ1ALNQh3UNgVTFHFQ4zrnvDWPWWST1U6SsRoFLgWAX0uFueqhG2
9Xs3Gokfn7isXtzEJPLlOpA8aB8koh3yXs/bKICmk7UUgU8Hd3wYZx/GXeyjXAbJ
`protect END_PROTECTED
