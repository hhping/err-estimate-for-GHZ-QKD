`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXdsHMh+wF4zI/k1hNZhXALy2ftpT2uPoVcctuSPZo3U1C/7vFpsL+MGUVFrjrMA
9mu8PbBLkcR1gI+ABznsl8KL00IqmFEkZysxAvLJgosbTJOQ3hnMbDHSqIvzOqZC
wPMgRpDl1MPAy+dJD33ueVBrkMRY2lsEozVHb7dadib1LQ+/2ebxci+Wj8XPKU/P
N7cvvNzOO7aqRKVJnjTepArIT5e1aFzYuMOlZqSfmO99AnxiJc2Lz1u4H6uAji5w
/291uRh3H0B4jAI0729biHq/uYm479Se8frryPSa8BR6M8MJV0MQxpArCP+pxNoH
6s96nxE5+SnF/PcnsBKNbfFgyAY8ZzIPTBqwHIEIdIFg3L0XcdoSJ+4a0eZYHGnI
okcrsagoAbCtn+on8IS9fT4UUDptVPVrhC4kePK+3ENzAp8YnRRZpfgcxmK8XRzT
khxjVx0J86Uob7RmP/56Ffgi+A699zAqhDupceskqvh/TkseJiH2OKNcVCE2/mO5
NUrNfDZkeraCjggeTNNz945/BZTh58Z8RovXKgvZHx7A5idtr9jmuMBJ05RwQgq5
f9dFxT20voNLjlZIpmzj6aaLN9J5IJ2hwnFFuT3EZ/uz+GPPDNkZNyZJyhIZolw5
kNUAjEetIWcspjz9lQw+NC0SUCpnGmSfcJmAznl1aBLWzmNI1pOH4oANVS8KP7la
D61OOxI62fNF8FDTsm2rafmC6+eZCt5b3/mWdXYauOfHADsMg2zyaJtYjMMk0tRY
47+nsN+nN7zwtxaloE3ElOAlhWsxwZ1Uwdb6AG//cHRC7TjrRfZQxabT6A72jfKA
7uc+L++prftdDwOia5ymLbnJVaqC0NbDpTFViNFZpRXiSFkPL2lBGp9Y8WV0d6q5
UY0lyAulcvIWmvMmROnSC2hgoq33K41zr+1g2CD/oqsWrnJDqbNhVwicquaow7rg
Psgzc7csIzrNzCENEacJrQqf/2bD4zofBSH5jbw2s/Dwx5+oLIlbghZZhgrM0xW3
/d6DRvMuD2ZuqnVeoZzYYOQCbZH3bWQyzkQylFigV0PvD0bo694Rg1HtgIbYjY3x
jYw6KJ9OJVX/jtKH0lOEgljl6YjTy38mgdkpmtIBGIbJx5ZlLn93+ZuZKCWO7P3Y
PjyOMUYP21TUz5ECaheebgs04J9THTHxgmLFTelGE7vWr0YYuX4noNCF0OCP9CEI
H0xZta5b/clq9z2a32Xot1QdO5D1iRbejlYxJxcVyrG3UyEFc8/mXP9PX/ePA2JQ
HNP+ZMlSazlCLumUnfkIgsYnJfuNo537n35zvtb8qgirJ/ziEAttkIHTi2BNOL1I
AzQ+It37DSC1upt7aM6A1llRZki+FDqo1JlmRFxhM8O8W1WmqM3Y5PdXy4S2CEUI
63uRQKP2KwFuqNfDHLCAcy5Ah/PsIjFtg/8UvTxjDLKQuX1Ter87hC53U65fB5Wk
iPQilZeZiqG+BiTOJrDYd4kukeyE3RGTmGPS00ZV7t5FzTrlQwl8TPCWku0dk/zq
Bj9xPjma5+QQ433LVYNOzRuH8mawFKaIXtg4IM5jpZax2Jx5wDHvOIqyptT5IXRD
rfudrbdIWuZJDnV+Aqb4Gtp2fqqXZdsCb96fKWtGDA6wcT4bXtpkJOOAgnSjZTw5
kDkuk4WctFFJRaiCo6oLwfyPi5td/Q8PyOAJFtluP3HlUs8b72I/5o/jbIw1+TIP
su9/6WneLwrA6uteXKII1nccnZOlsDqm45eKsAOuYyE/Ye0/jlH+EQQa368Tmgou
bVjTzWmSGOkl1WVCEEyuzEWJ0cKKAqVs1abfZ660QTGM68ytu7oyxb6/iAZRcJZs
oMMJxqpMeSM9ACcKBDivTUhMI+CzkgfJ73D4oWAqhtB1s7v6FUDvXvNdHql5Rf64
8kKIwp4CoocfURg0KsbzBZEGY8K390EmEQuPB+rOdbmvFCwl+D9OEolkgIyc8d9O
Ppt1Ig8rmonYXNF477z3qzWHtwAv2NcIcY3FJr7LcGx5zv0erVAJ27naA9AJ+URE
Z+mw1+mRFtJYlziZ4eaDoHVf7hBcsepGBE6Wrhf77CTIfotijGCo+g60FCe7++vK
K/EYJ4HKZKVrKrvqLr1g5rfsXepXmJ2Cq49jxlv3SjwVbegBEOELwd9U0KbSOhLv
dAxVi7arTXB33EMfjt1UYRuTxwmbgLm2wLcBOgIQKODQnrbuZYovF1YhyGps3cOs
NNoH7wVa+T9aHVuy92mVAzdqkaXHjHnCZ3qnpczlD7UJZ+q7FxoG321cmMLZEJdV
tkqpCcDU1DtFwxVHL4zpfI7IUKyYYqnhQyR82DclSZB26UkfB/5vvKL6zejT4ApX
X+e6tqzmEuZ2q8AoK/X1lpEqW5PhYb39N6iDZpeEOKOVQavnDu9HRs06c5vOsS3F
XroKbILxVOyMnGlQf1GglyrvrvcFA/lB7XOBXtguSxyDllQv56ww1jiJyhIpkyZM
zzHKdy7ZdF1RkQv4GTs3pahikJ88ZBWigTcFLRW11XzlGjjhmhQZuMNXWecAZeFL
s7L8UMw6dyDng+Pa7dRZVWjrc5nayBojS4gdVJG2fuQNd9xFzRXPqwepyU1SusTB
7wJoyFi/3kLXxhewLa1tzA1otaZW1FXZKj2WcyJOexucBHs8CrafKAfuNmu4ibbS
OU6iwCxTNziGscSLjrXr2Rv9TWMQOzZn6MlFkuzxjbGrL+hZ9Ln2yzAEbyhLG6K1
+1POfqmZk0lOZbIjnpmkazPLLcMTtkmPqtXUgtdePk6zgR8lh6ueZsA4WFiOhr6M
d3mGfymUAU+JVPHEWFQhx2AElT+MwSuII9Alcyy1KlelCeQOQEJ7NVnSw8PYDS8O
6x6URYGDs/Tl6aXLH2ZntHtS2U1DGxrIJvEJSDwlg9+DUNj/mnOOZwuMusOBSo3o
7vHwiFjx2F200e+iLcYEs3k1Wr0eKd3fQwnw2ybFzUNJso/eWGAMkJjezB/5hCZd
bz8xZ+1SrbxEqVrsrCD5wtbLiGLfaSN5rmtnjFSvCwnqtFv6FO+l8Suv0Op/Yjb5
Roo2mskNEXwls7muQ+Ga7LAHWWv7su7hL5YjVgb/PVh8X2k3Gdq3eJVg1niEM8Ja
KYIAwTyQAwsA42Di+HB7w6cmpOAdJhn8xdEXwLkhN6xIJrjr2wzYqxZ8axFvz4lJ
fFHzTzmxGHlXebo2NOteZaFy9coDnrdAQ/LGkhUcokRaU3zpBJ1lw1Px2jXwbkDr
LC7/wKE+1OAv8cSo2y2Yhqz5Eq/xZDyb/p74SIS9asKcIMwwvMZnA4sY9fZVoWUj
kh5yyVGsYhSdvmNNqG+/PcKL1VZDhK4jhpazk05sTbO/cZwMR9Pd6A76rdAmYerI
R/JeidMgay9Rbi2PfG9jvNNdPuSWE8ExainDkp8YaMe0Zpf7zUWkNJ65s498cnMJ
uoH/aKGMxj5uf6jDnNEO48JOLTPvqXmaczGteeRD0HEjs5O+Ir2k6YyF7d4fgf51
iwgi/Z6FlNdAy3hEDLC7g5Ax7DPVcxdJPmVxkmq2l478lBs7NK24J2/Z5GN70RQg
ZvZaJETdpCG6S2OFb/bG3D+0sEkxsxNxRbjauNLbght2/vWHhBV4P/gZhkYhV5JV
iQo0C1uuT0/iZgvl/PMHRjLArOpuymIAEYlJMATNYoyxaFzx7U4x3LYE5f4EPT0v
pWow5vKvtFldx+ozpfLZS3KtU4KotN//e/sqTTozBD7masT1zLFZ3grNot6/GRfl
km1yCJOZ0ZxTh+e5mgzAUxeD2zp3z7Om0SOlETS2dgwh5dnuRjrEnFbEsDeCruSn
ua248t8gPoqzizGTYABLGsHL2ypv7xxMJJgN3m3D+fyLy5niUchCj1HqZSj6lD4e
iiOmnt5HpBX4YROSd7QqmZPnNHj2YxAnQtmET+b13XqdqpM5nsN9DQV+ZySb6bJj
JZJVIcCSJDVQJ+BGHhMyb460sQ6lXIQXfU+ejzdWLyGN79fKS8vohTjKNYcqaESs
OZHD6f1/Ngixvj6WBe093206MnQipaSHzXVIc+jEaGO1rQeFJZ7hwMXBMK/Ovf+K
uvqexweemC2uCPWbw5n7v5M/Q7Xsg1r+LktqQ9pfVDajTeEYLWzPx6qaS5cT0JZR
FdHS+Fb8IXg5VRGy2dOR7UQhu97nMxS5G6Ox3V+CE0cTP0azHEQNsplh6oPHdXZA
Cw8nQZs/KWoC0UUttT+yfe9/pko63FL1ySRC40d2hZFDgVcWc2eItYkmmZ0A/qw8
ofh+xVlhzPTESE+5nMxp8D8bm+SqfoIT6TGeEfiRqAC5IYIIcBijcDALOrVHYHHk
elrZX7cwgkuEW9UsiZFF6oiByr8o7GVCbQ3tEjGFpvHTtg6jBqomjqbu9g7zG1bh
VmlNlpR51dM5BDuzJXsHD2ArhxLxjUXqorCPQWsCgfTzX1hKNRFtQtnFOKgRGKLZ
JK4sYaqgJtR2bVWJ8ruhqt9oWQue2VM9n4gKUy9or8IikPZqDE7iIOLRXgzpRL9X
DDak4n5YsDoIYSV2ZxTj2SRbaxeA420Zvri+WDoBT0Gunjnsi3hqy1AJm+xVrQRT
ZuVK3Inje9jPJJOqGoNemtgJHkruoyUywGRTywAPZcsG8Rt8606aupYGQcKdon9E
kCBY0RdoW51clU9VU06BGEuxDrm+O4ZbbFTfobOaCtLtsZjGQRbyYosgKVbL3bJ6
r/uRdmCwRdeWqbsN405azaVKsAbAErk37wH5GUIm+z5HiOcgFkLAJgx7/4ZrBtZQ
NhMJ9FO/Jl54M2fUKtGvRLXmXT4+hOS0V0FU/2xQHFK3pOYeIWXgVSTTxNs4m2Av
pva07bJRq7WPUkY4JfDQV0SjbfW8bazjWl7kE39PUFfeZkhflu25DqxUqXXJMdWa
th+S3cMYx9neJ1fLX5h3/eyh7Kd5ChN78AjaXsJUCCnhK95zojDZBSnRSAXkJTnu
dNEUf7QXrcXC93+IExGj1mxvXc/XLqv/NN4dv/yEVPJA+vP7S02lUTle/VkuG4aO
hfMtE2RdeO5E4QpmMo4aA2y3DYI4GgZ9yvYhoz70SYp5U8Y5aqK9a+6+MazE6Bcj
ZhfU4Dxclu0CZJRxw5kjVpcDjJPDbGu/ueO1+f+Hme/79bInX0Z7rzmRsPbWIMdb
LtdlYxqDf7cU7wQ1Qd9httfcrM3sT8RFP7YB4yPReXsiH5XRDkCs8hCg2xeDdKzL
t452S2YfkAGxmIPS3zg8KB0cafuPA+w1DlQIvBFGqo5VnhDI86tbe2ihrdHCY1f3
bqJOaYX/G5tmEdqFfIrL+i+Lhgwc+YL114EurVCUP4kajngWEZ9y69aXW6ww7UL9
mvSLbD6Vzx72vfNXG01NHXXvao6U2rAkVoFUg4l0CNteCgsV8qsDMK91RG92ubVx
eF5znYXkRqwGqZBTlOVN1OBfEqqVX3naeWWMshrmDil7y1LIF0Rwps7Wsx7d+fMQ
QfC+nB1U0VdE/pG/mteXw7AuN7ExFA+VfO4k9k1z8XKj0cFKTSM4DIOnMM3+G5tg
1WeLyZ84vAR/60oOaJwa6LHfvjV1zy6iU/hLAK4RCQ7mbSPCaPe2JQ+ZN81GjY/y
auTWmSrgx1RyaGCaZZOvy8hHq+49QFy17mMvxeyB9ZZtYJIiz13kOafy2t5iBt9j
CKy+kcSZEP2bkNNO+a5b76NflAvYQkKPxMfpGxqyZKaL/6OqvDzo3BEr0bceV7XE
SAQR+M/7o6VIgYZrkjDs8pLEYVlhyI9jyUZkysTraDhniuo4gGnPk9YlN7y9hQ1a
6uL+N31K0jt8Ty7mXCBLHSFENDehMeaOr/vLWQvTsGDarXTpYGLY/AdRWQ4aahSv
xag/Z49UBGxCHtGC3Qsyy39mpskw9sq8ZTuRBZKzJApTFCjDycMPAyCcvJxUN5Sk
SZ/lPvYHB7bvSx1su+4uizglYqTACJzjEFCc/GEKwIHpJnm1Z21+b9uoXM1ANJQQ
w/RmAatIY4E8NCr+PivL5jR6GDQFZY5vFjkHpN8h36Ndy8Nrm4BXiEVmeaw5nMPF
I4V6SfIRLdIjEvhRT5kYDfHMkgdcDkcxvHUMsJRyGrXRW+hWwqFUyfMIs7IqaFwk
drsKSeL62px0++eTTj5xfJA/y8rbPppao3Wq09jJRoeP1Blh/996as6sKdny0GDR
S0rykQkYYYezwmt7JMCzQjtkOxIECRvYxKrUdhluMirnFGg1DZL1fnzkg7+U0ZI2
cJBFhJRsf8LT+eMIRyeKvi1fh2R/Kra22HC0r72fzdr46rgNLZIh8h9HiApObC/P
19p36Xgf7oe1JltLAEYNfDQHHbF67UZKTg5NpzAPhZ87saXe46uQVkWeZeRvd3nD
8wlFOMLhGDCOObsoOujyBZTZ5+gaglDlnQGiAIVnzZ51hr1rBDL+Wj01PNfznRuV
zFDRDWLxb7L/MCOiWRFEQ98S6MppsWHmJXOzcPu8SPQgecrSA3SVL2Tn3O2v0GLo
HAxl8xbPXoiVr4rrQGopJ+mhUBDy/iX0VGFiUmZbVn3T++kuREtJFkFraW7KNh5m
YRMddFEs3pTTv3pa3gBRgPFii3iIUVgEGhTIAbp7DhE7e1n27r+KOomnYowRy5kk
Qa6gz+yHZpNk+bzj5TG1pJxQH78UQUn9cKme6837b0MNXUDUokE/D+uYXS2GxUFH
56KxTSsk+qZiDECWgSrnIbwa2Docj+TaWt/9NRtOyK4C+KC4hliGieQfI2DwqOcj
XHnkkGIc1/JDN48JUqoA5Y0rX5tA3RpE47g1SNSWHAyK4DAFcJfZ9z/F6V934fnL
TV/WVpx4t0pNasCntuswgv2dXpmcumBNCppOasH/GDQCtSewZh5iIuMTFmWeg8jp
dnHpPz359Wb4RdhzyPv+kUwjl3bwDJiwPIhBwttcuMVB4+yD5+pLIrsTR9Fo/UOk
ICJfPt62tgq7EWfIwb9NgbFTE27IWUQgxlUu6L+SUVoAwygqKPfxgWcumktfPtXV
qWGOXvbqwWS6u+aq1huBc1AJkkxvHDVJWqNMVzlYcnuVfUYmE6BR41QnuaejSq7a
9n1VCYE0f18pxPRXwx1Au1m1cE1pDoRWuR0mNAudKGggrGOL8jxyR0ypR7hJnBs6
2EHTQij85/3gxp+qoBP4VwGWeqhUX+FrO/PTfnEQcLyrLRWB4ACav9Vg+8pWXegC
HFXn0kPXCj27qdy//9aMypa2C9nPfbaLWDWcvegUcupGnZOq8gTZrI/+6Cx7tptu
62cTCL/KJoKES+APxmjMksTXF9FtVY1b+XfmasJKqx5Q8FbTDRJk/xcauL3HYr5C
I8019Nbf3le+/bcf3tCdmLXOvkudlwhj0xUKA+Cjlh4h7ouJgf2VSMIs6poR2ZhX
p/IbxjdqHJJvHMtKU8hD7Ivi/+naVH2LpTH64wNDWCLF31dxGXzh+eUMQxe37NrN
eBG5qmb3mb1Vq9hZF1thLQhVEYeqr/24N0q+tl53TdCuDbUf+xShEdKZlIYrt5Mk
+N3ZPT7lx/jtl/YyStRe22nY/my6dRZ/H/zyNIgfXzIdW5i37POvvMtHT8bzvaBc
6fQ6uq8+L+7OUoZYoVis16s22hKhEWVsJ5yTBNqZlFXRlcdVYGBuES2VK7/iXtmn
M8HfMap+m3EUnuqgAhMRXHuzsBqcTImFPMZfAuCSwtp+i7QGwjBkDT3SXPcJt5a8
OKB1lh3xCj8TzBRCutjmNovwGtHDbPN0g/14vJ76YnPFsx1gqoRAmVxRWFfbmh4C
gEKB0Ne4WWaLzIdMKjsiVcEDh1pq5M33QF4OqOqwVO7/w/3bLB+eTU9AYNKu/UUb
P8Qlq6Izbc3AAjM4bfbj4mIAB2oT2977a+o1h8a8fcL5ooBusu5zW/8T+pWJ7yyB
yL1IQFiTZIkLNWNxClMvRadAv5H1L/9R4zh126cd/qeW2Y8GO6IgeE2ioe2+X/eS
4SVaQXk/NYi5/il3dLf0v2GkGGtPx9CRDxmq/+1ZSaV0NEmyJimPKI/9mNOHvCrS
l7u3EslLxwMEijgO1xk2fUm/0FP9PmvByHhXq8u6Bg5Y59icfN4qkrSf38MPvHnQ
n1CUP4ytSJBDQKBp3F8TW5MuLN8g+AtUjCYxtyRnQgdN/g+Q6AleHpj/ZSO3k8Rm
H75tuTh5KuSnWn23wzcYDZtfp3nWoD0jMiDC25IQQtU9bkQ8FF5EJ6FxkPjSeMnY
SjvYXiqR0RXVpWVIrGuBuENfP0Uptb6R2vqKLV6Ptnkzf9C34/20k1V11N2QUetn
SBXZ6WKSB+kNIBOJMkr0WaQO4aktPNvbC645eWkIdqOuJ4i6hMQ4DahW5ZlyD0Jr
fgo6DzOj6Ybv3/3zMJQsvSrCCt/7EBeWJoT8EjqJLiZJszn4RFCNog5Q0VlZ+Osa
7trjpjR9OpXqjbWPPmcr1aSH7ftbsUitRS6PqRMmN2sx+IhLvrCYuomOiPalz+Hb
/0z/0/d4ZpFiNNmk/ypstHaMCvFeWCNWaJdb9ce6jOuMQYovGQGsnXi4JfsogzAh
Wzn96J9PSn7PeSiDuhh3ImWtzKnqLY5Wl8vSPCH935uAOmdTpwj/0tWRpC6Y8bw5
6Ujq5gUdgnP3AAthrkypAK3PDf0dF4sjvKa3D/XEkcxJ7mF6WbMllqE1fWPfmUTQ
efEXUa6B6JsVsrya+PO+AFdyfEkMmBEJ7fS708AqMgjBreRnOINJWZID5M4lsSG9
fHIAYuY5Lp+nCg7W3OnrQZVVVkEL6kd6I64N+t13kHyUNJSxAaThoSKHItvsKwJx
39RZ/94+iBA5pVeRM2S35WMNPCZm3CJMYGDRPC09aaMmiWvdZ6MZCWUw23VK/bN+
DNpeNRvM22QRMs3i2GqRbjQD6SoVsVpj7S4G8khtFs/FScCls/vd0aL89RMddsWO
vwRGYWIk2zkHhKGKFMR08UlLXx65xTXoVwzqZDICQ/+zvgONdjb9aLPVoIJnRQ9F
gzkEQ97zw/Hc3OF2aa/2xGb0SnBL6SfY1MC6SKMt7P1ihxhUD1X3Z0Cr4YePI3DA
JoosyGWT1qx+SUYgHwXiHRlFf5Uz8HVnD4rEKEgIETuyPsRXCufl++z+X5HDmOem
R6mRCFOVgrtLY9QyJgKIF0W/fNQWlrDRd/AuiLd3M5PlGLFuW4hOfyIgPJPpp/xY
HMUmgOOxRf3MM8FZ0aG0GfpQnuTpRmRJvyFrzOMyOT8Tvspwusc60+A4stKe0wSb
G++L+4V93jPwy/RywZjgJHtofVpTShu/X8FaM29Q9i+loTuJdeCqMvvPEHV7+tKY
l0QNZfxYvu3ZLJ613aLYZJ4BKgNjP7bi3HHzNXURE+N+PSOJRs85lxu4hVSqOMLQ
/BbrVdsXH+kHA3hW8CnEXQ3Yb7B3JEhJN8MjAxKYRBYeMUkpNFS3dc6H4/KHI7n+
V0IObgbRxpp24qMbQMdLBHrb0OjLgZfVn/uEMKyNkmzeKQeXS26Pw3Y4s/GkadFa
ds5+mljjKbX/iyFl0ExV13GKrtwysZRFbEAD/jvqDj2vPBv5R9FXFOF3L0xoxzSz
7jHmTmxxclPu0aXCPOF2j77Dl+mME2enHkkcQkp9vjXXggItMneBOtqgiN7H1KBF
8Hal9leDrxRs9O0YH1CKqoYlghHngcxMoRBp6MAB4R1mS6utnSyQbFt/4JBuD2Rm
P4SgaXOG5jw0gSA+vPnBN/+3uSwbpWE4UFHwsql0WAoEMGIgdXBrqEEC/kptUfod
vlZtQIAJjHHhaPPdcn1P9mvveQ+vqpn+rIKI8GG+E/DNRFIq6hWZz3z42NU63Uhk
CKbuDdEuxreawgKGfK6SGZq9Csy5IJpWktZ8wXfNV/ilSRjMm6fuuB/Th5GnUKMz
trmT+K0v+fnrkmi+tvZnKDY5Su/l189USO5CsAKFrt3MWvrA0bt2mVwplkJhn54u
5QqAb2RjeJTauZ0Wp6CT8cCreP53hyUkGjJWQ295r0yB9VlR/aH/W91dAZ+SlSno
QScwNrSDgXH34wtTk06u/8pzveIQqElVVoqLZlxVcMioqHK0f7k6929m6hkKmKu1
+/LtuW/vBOKcGixQARvuWVJ+s1Y2tXJKokI+hS2RgL4FwIspsKR4ZLLF3eJCPYjh
8X0eQXc0Sz1W90AaZ0G10cviI23k57g1cXuKhdZTPhspuTHNtvlnino2IjSALnE7
wokIQ6BM1FVqUIRrXsj8E3dfABqH5rag6XlYLgJo7g0eYQOzY9+vLysYaRE1zLZw
Uq8QeefgpDbYpV29qYNf2+4gxH66Bj8+DM+gVwLn+Lha75lf8W9IQvqwpqxvBSFo
L4r16ZoGVplgmtV1X4JTGIb4mpZavlGs+E4wW5JqqSZcuoj1rXQ2dRbvYWsdAaaT
xrlmm3YNFUXPaPbsZwfJxOZHMpfT8ZM/Snaya+3iRie3swhEQ+a1Pp9aEH4Fo81n
DHxZGLOoNUohpb/bpg92TLwHFGkPWEvgtO7tTDzq7eVymOvBo0YNuxq2pU+KyXt3
0VYdeNIzXy86sFhCQ2pVPPnCa5C64uAbgiKcZ0IkcrhUxErVqCCi40NEi++6ufS6
PVwMwtRSw80fnMPPs6sz3T7Jpn0atwfrnSi0Qb4HIRQYUE8e8R+l0JBgsnYWPdeQ
lqT85jC/qEvimfo0yCChR8yW5XTqeVLFZCTYRA7LJIyAd6ChY/hoFGFffPbNa2Nb
WC2SpkuObpglz9/dz4hsBmAclszrdCDaAJP29qlGQo5RicuV7AymVfX7+TmbLrFS
bfwZJYJmFekC61dtSMKyFBsQ1mjp57L+sEqKT9XAZfp3CldfA+9ZJJTnIZszprwz
Ojvor/h+QvbxSg91X6zLAdAgLvoh0kwCOl5kVIeYNmW+nBPZtN/tWWhWJDEHBzyP
X+3WTs7FG5tyr5S7TmU4rps0GPSrr4rvHd25YbLY6m1NGO2eGFAG2yGH1nyGexHa
opiiw8jfeXSleOscXJJYT3WEuBYzlh1KC5ZNl7zL4V/fo4fIXkj8Uk5/5zQ+0jYF
j8gfScc0fvG8H/mKAyi1j79SzCmFu4lR3ZZ8YGAwUDFJQNUy+snq2Hkj+UxQVfL8
zrEEUEo6ZvPI18thpV+PwUCXdceqdrXH8oiw0GeZOfYwU8nggaUEUUg1vxcZ2Qzk
EVPVzU1NpuChIxmne56e349oLr6t6pQhRVQvD+4+sb7aONNkNKAGvKjXOa/ls30D
fkCruOUtPlD5rS6El+XwWrpOxgV5CeHAxcgCN7mYbzIq5CNV2IRZnJeqt9hUriW4
tz4YIEhozc24cfBSu4ZXlxIBtuypeN7IsJOD7oNucqLHNU0wN7B5z5UEkaSNMxMU
p4em0tzQXr9JYqdHUSSK4XvW/cYNxFLpJzJgk7ZB/bfBIRNpZbmFNyfC5K9UpOP6
f/VfYtLMu9yKwkRT/urs++82Amy/E9KwnDw4F0n2spM9HjRXHUT2qB0yR0N6wZQa
Tfq5Eb3XxEpEqUM8gL2awg5sYJT2lXeRYliQC/DPAH0L8C4BG1uqUqcXYKgyp4eF
NPdY6QYECIO3urJqrr5Y0DHiTbywjDo8XFzrpm8CLbQlV1171fOMCm/nQOa5YrfM
wli/B1Bgbu9GPE5UJyxoLK+lDLKmCAa44N0A5ifMQYYBoVknExKiGj5LbqJLCCnm
cirOB+gfvivf4oqgDOoQdryPR+d+U8NGF6yCLx1FzyGjhF4OdHlQjrz7f9bhoDUG
ZtwLKSiZ2pjIl2m2GJQUM8d3E10FcE15bdl9qzHaWwe6IUr03SDoz/E1/H7Syj7O
bcP3bFPNLVuwvJSBwhado5nKs0hO/v5EE5jJ1Plo/QlFE7cZDdN6LsyBFFScdhq7
NfYBQDNKUZ4V7RX63lgsObzSenyB7tsjTGB3DwKOgXRTcYNncdALkLHUAZjvbrfn
nnhy0ZqbbJktGYTkIQUkByuW62JFhj8hFxLLMVuznLF/2o96/R6PJ/zatyK7QwyQ
KIlIYmFnjeHpV5a06CPXIAWCkDOFOL9x+pFfBrZBoZ9uDcgKX4ms8bGU36r3bUwk
ODgKCFpaOGhOUGzgQO2knSNNBOH4N4108LWsAGMdg0w9wAW2LNngx7xE9eVZykRE
NQhSzBHJ/4mGynaEZqgkiVyZoc8UuTKs0vXVj6MElgPKNMZZLSKnCS16wTj7hxNC
fG6R8bP70sX2iCI/e4y1WwSz2MXrgppxoJUa8iXaWDxsl7GaYKVvzMYZNtRKM1nB
i2GgT9x0PFvJPEf1+4VomMJjXZfBnQXWeQGj+daT+9xVA4rRJbOo6NRws+U2dhCF
nIgn1FT0vJddbpeNsGTQ0ZAMvyOwtfne8fIAUcWaD+msQlbVoK3wPX7vtDMo+7xU
HTSpZMt6KT95HA4xE6wA6Zs63TrqwiuvKGzG3hnjpSAEQ8EvWcvx8q6b63zKZxSq
IW4iCVlFeUXPuyF+gxJ+YYpuNYGIG94+x+u88xwVRDu19h4FC7HZ7G4lvtZDaQ7X
9bsqZKY21DtV9yqJUlyTKe8U6KR8pOKQtTN1zLmBTmXcbFL92Mj+tQTRXHtVEcXt
bcMP1zQRHn3i266hdjg4NPCgGMGko7hlAQ5O4ZsPeGU5WHaT/HtDiybCsXM+0B/m
wMksSs1JhgtsfeeoLfaPOg==
`protect END_PROTECTED
