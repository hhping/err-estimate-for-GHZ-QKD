`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+UxVPbg2DKmxY6bkUoYmTSSwx7Ps+5Eyvqt2QjV/emShDznW2oT172RjSrwE/h8A
T3qdeI6hkIkA4wLqL5Azz6/RmhwTJdCjNX/TPW34reQq2fXJ94fLhGxTpjamMB1g
J4I6ULLlzBWxCGzum8sVzb506P7GftyfEumrpH9P4O3zC/HM/MK8duHruj3Uy68S
iEnFUpPpw28y512p3XgQiQJKwSGjtryOh7MPHx4hYl2FxzIQ5zgOCy6Tnl0VcsNn
hUEfb+hsd91gSPO1XL8Ls1muaPDgofKHWxg+JTWzTq/1QYDm2PFR+Fx/E0GNjL2J
ymBLheSpsITWD1QuC7RAkNLUu/fUD4+UJ3ugfe1Qn1c3yl+odxvkUlJDE7Sf0DXH
Yq0Ll3/YaCLgfpN+gptnkUGzSvCee8EPUPOmZZYFlewuqOxOMHA6lr2dzjEQ03wp
Cpv3jQDw1iMd9TX5YC3M/23EjtrEPQ254KbHhzvahU45tFrxUmNzMyB/Dr4D8SUA
J8IwKPbIYf4kzXbzaOdugToHhrf4jvdpue/ys5ebVkMJyyHqw1cNnjZl5RXmbGXv
0j2sLuKRqFD2Z77UOmf64vOvFazzK4/K/Y1Hg2TK5/iub6eEGZuQNi54O3C1WEP7
iXnvPWRQcOrLNUiI7TTTpCLb9nefNYEvx109mxjIpwqd4nGOj8kSVzviN9whh+m9
hzq6kdmeXGLK2WDAmcFXuxToc1vmeWxjud5rvJTQQGU+sMEGZN6ESKCZEzHNsZ9/
bZX5jkyd19mdWwSfs7UpHlQ5jip3fp09QwCk89wFAtDBeIHwGFjPgP27kygmUu60
45y+qNhO1GnZgfgcHj/O+Z+aoJOjFpRwEvouK9ailPyyljWp4KqQOuR2S2ajgtCY
Rdjnsv9Z/xKJlmEU1UlSSBbHgOVmN7AhxnUVZtbaykm0A4+n+mvigBSc/u4B8+II
bOaWl4lqNFUloxtCEZo/TKaKH6C6vuJz4XsUxlaOlX2V7rSDy1yo/XKYCbRAvNA6
WeElT9HOGZp0Nt+3scEZkpX8RvUdAPHIEPO6Qmbf4UFVEFciQ6hKh/kpPY35U7sp
Byd/iX+oVXYP0mHr186PrFZME+dQJI6Z84PLJUf7bUKXWi8HSyc0I6PMBB0SlZAd
fS9kjXjgsLEfVDE5zt+2kwOc1wY9ybY1toMh/SWZy9A/b3e8rjZ2dBppDLgOaZdl
UymKtl0rckNonXvk/2tMsKc8kxi8xE4dg9T8hCZydWB7HdXfvttpGJvAscbtXrn6
YUSwf55tPVpOLwKc6VB/L4LDqRLyffbDHn/ttNACgQQjmyl5IC58MQULczbaYpr4
u7BKhTOJF4uXoOn67wnGQAzkwxvAEjWR5X3wMAQGsD09VbP9eaxgbC8nVnoqCE7z
gGxjZdbqfbhSRNsJiEhUBm1+okLX0qEM9F71iZYaQqKn0yVFiK9wKt13TWgtlwiE
NLS5ru4Cb2pKHL7MD4b1o6+lsgyz6O0aa0oKE64dbPgfK0SQ9ibpfO5paSzr2cTz
iDTTzU2Zo6i0XaOwDulvappBq7bTR6Eo9Ir1Wll9M9O8lePH+U2fCIaF4oRV2MVx
eMzsQejHvJUJOSgNEmheY7lWFbkJloncA5gU8e/jorekyDSGDMpBR1vI+W1xjr5G
BrMI9t1SXJz9nhcveMFEc8aNBQWyOa+DeAnQno/J53OTaJFmlVA4aQwqjcaHp10z
tAeK8FbQ0gcNdMiU1n/OptPSeODJp5k2UBZ9kXSuqI3zinnXhlbeckMG2E2SDi/2
aWqli8ZleER7JBr9szCx3NvRoqrPgDhszZDYgPxpXXt1jVhFPekt9bNcqrR3Vq+d
w6DBcVcBpi80hva/9Km7nActmjQJVhGkZOr+ldHJvr0nZ8ffjbxRvCGAp7hWvRj5
xrG9FS8XaCB/eTPgP34s5OgQsB4iRd3jM0J4TZVbiZeN7NJ/2tg7HZy9+TtQGtBd
fdK9x9VyBE5YuxWta7zKEDpHEs6P9sFw9HJ8qN6M+o/LCLHi5Yu8HGQK/YA4J+fQ
Z3T1YoxVAT76H22KPgFwOzysD3rOgkPSoUw/xjxkxtPZM4mU3kdDm8uGF1S3UvQ7
yz/KIKfjWyDnVf5VrDPAUv2e9k/8FVhG+RTaY2NGe/XmQzJbtX3NYms1fNnntOxg
7GSnZXvrPP/5xMCu8CfNY9uSOT+rkVoeuI/6bs6mtA8XSM+hVZC3qSUg48qn2qAB
RFQM7dG7EOXDEfdoXxzi5qtw0DNbXCXPNDm0ECsipImO0swaKhcOOCgi/cujDaay
HiiFOV5T1wTTj2ZiehifrWpeigLawWQdh4JXNDBuioUK9VYAvZ9o/TNMDMSxmj5x
1l01+z6KlX6esyxpGDtE2kn4nuSc6LgtIGPrMp8+7wqT29Jimm2PQQjN4ztXeXW2
ExdOqwSYt8aZ3AtNeTyRjjrACO2PrsRLGlvQD4KQWP9qJhnRPs479B4WCYy5w4ag
8rOgTA9FoRLu6H0rBKSuVFb5rx5nUWJtjpPtC6+cArIBULN/jkA8/dg2f6I7Yh/g
FR9jGGLUaeqefxF52kIogKuEU03VHBpkE/wOdQ5XywkD6AL46OWQ8CpWkjegipQX
srlRzRsVWArA7n8cwXFNk1sLnIC/mayIBJJvZ/mz6QrMmOx/W6R5eWMvZ/yav99Q
mNfLi2RnoBMVVd8XPhWDc4SFjvuq1PUfTk728bm+dSTzq/T7HWwN1zpartfIocOl
u2uHpCeL/85tzGgzU3dmC5VNZxI6ZfuQ0f1zEnMudBZTNXCnYNiEhfcxmoGFOSa9
6Se+qJ7nGN3iRr/TkoIULTuzRTdwGXN3OVrPZOrdXBjfzN5zeslfDmGcx1XHpnmS
9MyqMs9CtqBsALp/5yW4kHFsrrJevVHX4DnmHtGRwBT26Us4xIjv018+5VKF5JKq
yfHde0fG9AcXqyEHvPRGPomPyXbCrK9Gnd2kT0nQ19enm3oe7B1FndLdnEJqxL67
CQ0lWr+RcZJRXlYfAPDpdekEjf1/oRu1cAp4woVXSi3kEF7iCj3SgyodqOJJBQJm
DM42YBMpFqLJ/Op/o0riVgEltQPRZtPkrTxN7Zt6/Bcoedcux+FqU/Hfn2b8Hdss
oAVBOVdcBoU9C6AxuZ+5PxpBaueadAIi1G5311e/osBCW6a+ZFx05zGIyoFLg3xk
QZiTdkUg0VlXmfIuYzSXdnm1AijlUUgMQueJ8ODzMDXPzC6s/fRB2NKVfsfcJfLh
IzrY9FAlJ/j0vvNtN1lCkaRJRXgJ3PcAC2rw4fJ1E6kgVkHlTgyf3WyCVq2BbCtO
0niJvrV0rhKTi5x0skBw/j28eeD2qH2DxT1qkRChJxV64LzBWPGArgDHfpatchiA
+fiy3wXafSqA57MM1Cp1yoYjSlc0wyWGJKfoqcFtUTdatciHKnSEn8aKqRyVzFcO
OXXJ7omB+FiLfSnjVr40QG2P4wI+z6YNFhO8quDulC2bRTYippuF+UUF6YI4c8Lp
1NjOInjHvFun8pLtN4ln6MLaCb7KjNFmhMilKcaA6iQJcfbJTqZR/Yq58+362xVa
67Od09trc8devaEzbAGwPcCkCOeWGbZqrblv0Jsn+4TPIqY7QiqS4M/4ffds16D4
tC3TcpTpkXGP579S1rfkFPZ6S/vFn0v6JYb3Ke9BfvbUWr5MQKX3u67RBmPp+Kyc
g33N6PSGuZOuj9ARs5yVF0EwL8cDofxLAh2ClFNE1dsep1acMeD/fOECnxRCOPTL
sL316gfDxckH07va/S5nBTvrZj2KnNapBT+ghvNfROHnUoO3NpH7peUlUPHBjnJV
2skh/XIFwNGO96UnBD7eTA8qkZd0NGHuGzT0T3tjDr+vjpZUO+aqGXlB79i+/cHQ
aTuDbGTadr+j2QJWTGVgbIa1OVXX6HzLpF74daiBs9kSNqnqGfReDztBaG5S787v
iaB/Ve1XYco9yNm9T5HlhYdDYts7uKSVKt+Gf5AokZjAm114iqjaTEgeZXVGcsCZ
XpCEbTLvkx7z4vBkSDDTglWbNiFJyX+vRbpJrI/PeludFVAG3wZ85pVL0w4a32f6
AzRcrGiGN65o1NhZf/wrQtJVOox414Ev0D2vEDo44kDBKzo/bIO4OdXue2Jgh9QN
0XrABsPkeQZ6jqMJkNhXhZbelLnJS0q1hGAY1sKUJ0DvYXhB8E0T1ukmp444yFsq
3iXJ5ZEVnmIHNiXyfTtqwxFePDGuofoB5kudJm8ZWGJf3AxTaw0py4BC99+RzNGk
ScPlnrZYklJmFGiFXe75JNagzG9Niga99PysiCQDnDc3+dcIJegZotXeNdYvPwA+
6LVngbLpsEjASt5GKrVqR4upRxOBuY6tnL4x/zioayUjvqepMiegaFufww3/QNMg
wfPqzmRuKQiqmASEbjpWPhnR9zJIdU7+Z6ZV2ZxOF1/qkssUly7OLu3G3j3CepGu
hLr6031/92w6U8S+rKjNzkuOdwQafCNlBpwU+k9SUCms0PnHQ4U5cML30RcNdJ83
cGL/RrBOy7eEyTyxfYSsNoHjT4IFALlAYalHBCCYyKPsrdBGkUKwQi8yN6jo7Idh
OXbrAYwOc3CdwGuQPAeL9MO8C6ykwkgIWFjN0WrWrP72tPFgisCNcL/glYUtFeoK
70irzl2lcymJfpnXTtNBv1nOpyiyBqmyfBrfWZLVkD7v1Lrvk6XV0PdfAdoqyxGn
vU/NhZC/hozcDuZ5OzSt5AUdFeIJNOKBRwo9ZWO5a/bibmD0Pb8tUuHMIO3zjwIv
LaoxTcNhH5oTSj4VOl6+TkCl9FZwwluFS6rPzQceKyo2a07WpXpan/34aQxHYX/6
Jp1MXWmV8CaXF6EXpY8wMUKBri/Y8e+OAXQHPfOU2eYhi/Yp2+hA9DVkQw2Wj5Hy
NBNvFcZ8ZihhL0tIuaSOasjxAOeuDxS2zN2vJ3efEbiZRgTyujHsjpR23f1BJrDQ
0X+//6o0x2GOE/e/3UiMAzzox52SSbQmZPlfTAYLHuDm6CW9OdKXaWULxOPmpHaR
v8zqNl6wI+OQl5ipnqXXQXvr3Iyvs+R7xh8DJbHoCFIvq4BRKxWkyMUlPCGDrJhw
vz/yGP5mpTCd0XI7rmocHY8utSrStYlGjGceTR7pgjlEo0HYJfNYuBa3N/WWcAla
KXTsxobwfyNQlFxlzPr+DG+TvV7Tlm0FrIEVGrKKEb8PMNP28ZtA7xDz9Q6J+EwI
dF54ESKSspeDh0HFDfsXp6ILF7PQ9jcA1uPH36b/9uD/HnZmjFqBLQiENRWngtaH
PIk8WktQ+Pd5OGfoxMIyY+BDvhmmZ3OtvcMznLFpPc45FSvWQoRM6kn5jOCZ9/eG
zO2iYDxeHl/xPuBZJJwNWWVE3EWVybmKz3+q9BWbOxINR8m3Yc7J4uc56PUdoAu8
2lArfsiDq6a7KUygCN7Qfto1iuZoFpdUPf5kKAb2Lycqqu7erumzmjQeen0kXhJh
YfxXxMX4c7f7h3jTfespGKtH0e8xYvmieGzj/IgGKkCtaeWiQSIESAX4DUVorN54
Bma3WGqwt+3gKVGSnM5mMhS6Saahj7Hl7ZKzksfUl4emfZvsEc+iZuczkPOYmGTO
1DElADaQjJcBriPsnA3uVCnsEfJInSpIuAmrWnAIMZpyGyDPe3NOhT6SfkmzQF81
RmBfwDIwJoSfaRFig56h4hAU2eWlNnkxjVLwgYZOoGnodr95e4x0JHPmhN/2fR4x
I5msuBTda2fgyzizK1PEi/iYQjjphkqilG0dXka3h503XfwG8205bsLgWZVUem4I
ynfHz6SMrbLn/vYXcZBd+yvSkTy/7gInLD2KiUspYPxX7v5gCh3YawtklPaY/zJT
MMnFYvl3T+cRitT0IjGdCuyUpT+dNeuNu6OEL+EpxretWJa+DxyLobU245zqJrDj
MEdei0h9prfXPb0IIprWT1SBKlPGSc7t3S2pApllio7WDOhK9xQmV530PdAlNSKN
IrKwdC0QAQ0Uoc8BlTFlxrSFdLbSwsBR8w9VixaIpcuywx7YlL96mRFgK7PXFS1p
QkGLiXWtozO79oxppps85OMpF37mzYBcvxxn3NpSKgoJm2Hq73tiZ1cZkGoJq0Gh
JDvyz4W13n50Ny8rv92PH+JmihGC1n9Dvwufj95s3E5s7LUnALvQ1cIREYL7e+I0
hna9czoEf5h8K7CSAPNTSIfHJVLYOigAmc51dOzvmqvh0E5u/X3xVzM/rYPyD08L
iMKQf2iNjEavc3tg9/OWxTNsVMjlXDxB8okIkn1o7yvDSsRs1wKy9Gsylcv9Zb9K
16wMXzIFPY0OtnI6Pkf2fZStM+GHe6c4R2xnRoBZ1tGLadL3OWaMt25/bY69fKPZ
fJxtZjnSyRG+LWnfzV44BvBMZ6RoDqma9+nB5FourD0On1GINfH8Vid0Njh9PBQh
fmEIAMbuxgkvDpgQXu3DorNb2Tw97t5TP//eJmBLMBHITDEGAhbgWFmcqH+r8UNd
01vdRFpySMtc4zHUZakSbMDARj0axoQzesJUpSlSrFyXH1sTdCqWd039LO+sqvb2
4w7k29Xr1asexlFyuedDUTFSk9Qi/+H+m3yzqoBu0GDyi/HFD/C38vWpulfDFIkL
TAwoUvYmr0+KhDt7cPsv8iaAgHXW7RFMKPSYvJKBBU2RLeD4PWhe1/HZEpk+vsTG
SPjWH93m8XsTVvu2C7fY81Loi/aGa1IV2SXxuPZdoMA60dJ42l/yGwq5VnSBO+H/
8r/RDR8xJPlI1FhVq4Tz8LEuJg1Ica+xWG3gA6w+Ss8fNrmWkhwzW3wxKLykP2cR
Y366iUsYtxdKEX0hWWVPB/YGe/5WN7hLfzr2cLVcdu4MNPH0h/kcNgKn+llI4sjP
RLNm1VQzKIGWqUvcT1W4256jckzwTAs+hnO4AKue0ng=
`protect END_PROTECTED
