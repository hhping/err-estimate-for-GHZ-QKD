`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kbCxkqWHlmeqSVtj6SM6jCn9ClDBXQ5RxJCR1zYj1E5UZZmqnA7tL6hoRj+zbZIM
dRECCustbFZ3CWMpxXMAAkLJrd9EroxBPDRWVMqxC+KpZ8gzlD2mCrnMxovog0zA
6/ORbxYP3n5rWmMue1xXZgaZzBsZ91mKt9PTAck/B2gkYsgoISmMb4CZ75pyEY2B
itv45OLHWPAiv9bEaE2BSYU5XLJVyoW5zcAoPRzyPb41Rg1VSs6yNHQE6fJu2jeY
z8JwB4/FEfkaM2TwKofW8Xg5ZvFjHKfmUi54/FREXfBKHb50dvVURPRMlOATSwWs
RVf0YOSdumHr5ZU9uvggtI015RUHWKbIzqffx8OERVqFS11Av6LIeGmSYcWIEv/H
NPiGbV+XlpU+cHnhZGZD962L2gXKGUtHjjYt1Ygrg1vD/r4OGpy10NytLgGD2JOI
oKUdJOmVnkGeXmXAFWnlN60qVG8lObtyXo4WBUT3yoPKWZPFR+fgz9kiSmsJThyv
2l1E1dq5EnbF5C7coiVFDNYVdDlcSMUcJbj9LL/n8ANFW8aAI4DufyxnnCfGr/7f
RYgta+dWcLCondQRfaenVDw3VPIWDGBZ3Qw6NOa1zeLznMBbOgWUNkDdyaHfeLN8
ko/ERYpAFg2i4qDErGsb8aya35ddWC3mzp3lTcVR+yq0ExrNI7l/l9LuxiTl9aeX
64tnTktNn9D0HXN0fE64a9q60gwxaVLwkPSoBiQDAz+lVRjEgyAr2OWVwgaLLevX
Jswj5kP5CTkoVaTL5dpIG6DMgTsrzHBvYvv6Cr8gmB8DGAJncnUTfvoi/pMNzkme
WdG7ylCgv6iy2GO6IpXA1PVKEUUE1Q6laTxUBp8lA+cya0jLb2I1+utJnukjn+Ma
4ButWFM9lQemyx9R0J4erSoyfyJPmvXk+junRm29G0VBCaUdWFxpgK5akJY4RaVX
mJ8Gjf/wwcSFW4MnZWM7UFbAesvI7IOuTBGDF25agWxkXy4i2Cqq23CgWosBJ2H4
r2M0lkm1m7yZtoi4qIs8YHvWBcU9DDu7zRvgbR5FWougT/7kKg5gpmkuU/OazR39
nUkt8kNVOC6LrNVCsfyysrJGDGtnOtred7TVYFclvaqo7tyFupZQ7P1Dooiubads
rrpOm/alhqF1ygwWeKuSTRgIOa+LCfsc9VamJnR0E8GsYb1zAZUpWlMiRy4I76fB
kAN0+GdL0Usjbp83Q7mvwl9+nHJU7i8n6YWadpi1GqfAOasHncjWKGBgQad1dp1H
GzNyT1BIsS4sAnbOG0EH3CT2W/f2H0w6oaEgu4dljPhDTxBUH8MSGvv4g4zXjVJJ
39dmNuauZB75pmjHDyq+oelEQhryVs5MoRBBxMAjlROylRA0Fq3jDRRi8xkdqx3W
cHzYFNTZSTaAmORAAnj3CwhLSSUPH3otz7Y0/9lY1CsCW9mjNHfj5DXDkEuIyvPG
pO5MOP2Ga2f9LtBlWdIvBT4sDk1RL46TAPDTam+GvMxK3O+fvOimTxuEXvL5a1EN
RaenIHPZpzYZVM0q1GDq/14pCHQ48VsnEAQB9fF6LTT7gMMWfYxaH3dxsSrPlCxI
TNYdFhIMXxXpDlfBf931EUXOjwtrf4riHShz+NC5W1/sbPV4vUnlR53PxcRkckV6
bgRRndCk8OJxDWXuKndRvnghjQ/BQYfqfdkcVDipwrMkb3rz3dWqBqtw+h3XgA/D
MlsKNzRrGVLRwVhmyEHrbxmT9a7MOcz7v0s99NRHSw6Yt2doOmwTdZPvZGoWqEXR
YcNeze93DvhybVkZtTrzAPebuTtCEaXqbtYX8wzT/ahtAR1x7E8EgP0gxb0hG65i
A7b9uNauXv+Ex+DN3uZIcmoFV7l2Iff7mwXSgltKJlKENeS2Llw/IpUPV09ZsFyk
TrVSZKTDawaf5+Q1JxTMPUEqyvk4Anopz9jkZpPBZET39A+kv7mfsVofnVhbUTke
qF5iydEgu9IqSlWVBF9+b19zLoHPt9H16laxw+Cfa0KJbUKxu4Lj+tchQ9SLPhha
F9w4Ao41Ahp4ZZdbwN6T+sTDZIhokL2M+SMqM8Z7mypNubM59sehilI00L9dHipe
CIiKiZxrvFVCEyFIn6ihYqO3AbzUgfDZiKhYpdaWc/eyJ+LyJSrSByQGhtUQywv2
y2yU+oEn2RMsygCcaWy4pjfs/Ch7NNYUP+Su1yOQMQmkmDbz9ARrDATfeEHtsIgq
5oJu3BFkYKMh0MntDkwn+75W7j+OcxZ24EyBFMtAFysLaIstHGGmXIsXFUg9glK2
oizkEsmRJJ70FzumZtlYKb41hwlkUKAdKXwF5PPWPHs=
`protect END_PROTECTED
