`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSy3M6de4/D0XayOzxevq+A+uMtRuvpf90RTlYoZOmFtvDhOhzYNfctHRFoMRN6L
ZUUcOcLbq4JfSUGdia8CO1Ok5X4oOn0XQVT7stjXmEQsy49IL9dneJ2j7Rv6roPY
Wf9VIVRiw38+xod0RUdSsY4qlofb2EdNo75JDXHyXxnmMQz60AEmZjifVOdxW2kt
YJUAz9r63r/On1Stw2b81OeHHeT2R5FWHyPqZzNrfdYwXphl3SKXf+8rwCSXDRD4
mnkjAAGJYGAqPMPFt+Nc0XQhziVZrmnjBkNfrP4OXKLyF+aPMnKyNJmKMFLWe0yB
KeOZFaeQ5kTsroSakL6jXEShGriJpBPEOFmy6bD9LnJ8LP7YUZhj8YN2KOZVxaRy
1yh3J7dGVywQ+ZAwvS9FbnfJqyH/AYVMsqQFbo5f13DIwxxhRF8jXqz+/g0PpUGh
CI6YtvkGH+QAgOYj+X9kwIanta7dSen48met/v/qQUaJ4/HkqxrRXabh56mPIPmM
opdfA4tU/1W+XOPWSL0Gpg==
`protect END_PROTECTED
