`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPXnCBwXmFEP3o5+bMXZVkSkCJJHA7JjD1kHgRndxJF0yRgM4CCRWhSYrpNqUM4T
uSHCxAIW1LfArNnPHjnquWei09LGsuF47NI+bt07URlhU8EQs5Qv4gY/U13dwE9S
KJKIwv+LnHai22i4UqEVbtF8Hv2QUkALBXtdS/3CZEEv+6HwHYvC3cKjnh/FlLYV
hy+meDAqpEa9nyKGHixwSPvOLuZgNt82EZ9htZQYEeccrDhR1GxiV7iCZwt6CWP9
b3QDhsDRkxyFkEuewABI0MvfUe2xgyhrj4TN0TGjS3+ClmhRl/zQ4HlhXy0pEJqS
c82FkewJOzsojacFOoGcLhekuE4inFQiu7R2oR6srdt8iL4qkr0GrqBuiWmBJbTH
gdxQqRacMwKB+qXm6ws28pNbq34ieIlZJ6CT5Grs5hjMtLfyYPa/qCXfaLCJmYRh
cXRrw2cZQJEX5N/BE3MyY/NPYN4UTVFMyMJmZVMDt4fyutJYRMGu0XyWX/nw5qsx
z4osSPmtWCMY86s3H9CUkyO27NfXrOOCIr09dcM+0rd2M/CiwZp8ncv187+gX5td
UPPS5XezKaPARI/Ube4cHXfGORsApd5RUrrCVQXcL/Y6ArlbBTwAIby0dc0FVBvJ
GLPIrKpq6Cz+Tokr/oA3FJvtwy8p638NgLy5wkII+Pinbqkstg09Yy4zEMZtXeQx
`protect END_PROTECTED
