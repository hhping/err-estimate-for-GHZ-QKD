`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHd0uuWgu7AJVX540rp6CdCp/DuxSf0MCsmU/nL269OaERAZpAYxr4tbeo5mo12/
20JjpTX4UQrUjLHtft/s81ZTK440vG20nBVMcvtYIbtW99QVxUIH7Ya3JfrSm0uy
CahYkr2pBeeFp1kMAAEAB+h/CmFU1UZM6c0+BcHP0Dk48CSwhkzuHxo8KB4mkJDF
EjZ91nNuFV6fWgcX3mi4uWgJmlfq+ROUFWqMS1DO5K+FNGS773Lc8CBm7BspZpyL
st9NanQ18G1lquWZWJlIQYYNpeBs1i1EEuYX9WNLJnAsv7POwFRfKwHKcaMboTDk
m7xalyf+7h8/CPNnUqfvVfEXHs0nhm36SyVzaHmsMTTpv0hSD6t4a6Xxc4BMzVsz
FZ2R1gnsQy9NbUjM5KaC6it0geVxU9S+/mUIhq5tE8JGLKEkSS+5tO7wT5VO/KCs
CH1Z9uyWYf16aFZMx6Ma6rbz0zYU63KnmmeQKLgSyW/LN6j7bwXOYS1oKK1MhGYT
ZwcjprCDZ5k6Ms/MOEQafOCgCRDZoUMRxFve+P0jE6TAQpweFtUSki1L1QXS3p6G
HSAEyY23WyDSVCeRhtOQ6YN0gBsIpRC/E6ONM6Mx2PU8EoOimfxs4ZV8smmVbinK
Kn1667+2ezByJiqq+5fkt8Nx5uWqlOrTJFai/Tmr2iRXGK70svpqhOzsmVvEodNv
AaLxM3CN1rOKUNFQXqzlqrd9Wzp/UrXGvnkiIMVKcfMKmou7fOe7Lpd3XlDbCxJl
TRx72y9MHUq8alVx+KlXunzlw1KM4EiQgW34SPvWEOUlZM5rpRExOl0+RSv8aZBp
cN9hNmv4kd6twXAnMODhhNfhwbPkSfK3erf34GMJsF2yxim5nrNTIbzdL43sAX6o
9JmHiYV7w2LKiKdzLTkByThpniQumquysnH331Czo2ESMFZuqo7a/PFprHihJN5V
ByVAPY6z9tIgUiDUbyaB7ojpZ93dDPtXxoPoh0tHh0tK4P3Ylz53g63mX3JP2SvV
Wl2yzu+dW6lY26d1QJyBECW50xrYRwbTudE9vE6qzY5Ssn7GRoQdEB0+s5sBjFjN
/uB1WkZ/TL6oTg93FtJrZUQULzhjpLFYjmd2DcAoCpzpYoS7wP74TVF1dccHRjJ6
Xn+i6IOFSTXHdmplY9KU50TXtQ25iATndLN7UHDN5eIWfYWePJDcr3PXYTeEuRZI
71+qIXTqY4VxJK756vIjmGiatfhkj1rKhXHY5FHLt39hS4iT+fmpXdmeuXk7KgL5
GQoUdLOo2TmotuZ4uX+bJeUrDFrqXSjI/cxGtX5+IxcE6vGXgdNi9MEAR/cxTURt
g/pFiZZxCOPfS88zodYsczUYJjeLxjmduY29PA0o1un/1MmLqNXZir+NANkAQ+Hc
fM3PE+U00BRy3ISdDja7V3KhsV5Uy0JtO9a850PFhFK9Z2Blj8P35B3Hz1TRXJZ6
urpjijC8UGXDFcjpK2deK4SmkcajZ+MeG42zREicNgvgXY97N7t98L5Aw7fz+rR4
rh7dDpH90DVU1ooBjO0M3eKyAzPOAxWLcAMS+8wUcPzrbdD3P5Ewba+l0+WJglgt
Gsr8A115cRYxJ+6rZqZB2a/NnYBFbbCorzlczRr4O856IcMWHffTxDppSz7ijPwr
kWDPwk3NGYqtLr0ILGVtcO9e7T3GqMCCNgjwDxSpcOD5hHGFjogE9QGcE/Fy/WJ5
n08FaiaTJ3I1KmYjv8xOjiWxftZIYZk6MAe3aVrUnekRdBABgF+uHu+VSfb12QON
qS/LxYttP7HzYv4TanNZo/pUPH0iOKBNwVV0Zc3vd7XZ7F0nzetB9J82OxXUm50y
wBBJ0l3kbGEvAbObX62SjTW+5y4ksZYR4N+ETFSzSI2zBKwgEv23beBzWcmYDprf
BZAlfKTpIHF5dykWLt+P35OZkRJ3h5n7A9hpslVRnSiQ/3Q3lDg/6cY/mMdWLuSP
TawX3i8FM35A86EuxMGkleTWZkazYXswhcLjQCTRWrNYGQloF18jTQ3NJ0v8tug9
DdzudE/EjZmQjd8hmv1rbOF701bPXucAgygG78fJCfEUbKsIHmjl/u3bw3RFNlQ+
T24KRFIUaeMA+iVhKg4mvqoNnHJioSm8wiw8Z/g05cD17mCDAhG2jj3dXhZyx8cF
5YGzN8r1ggHAhqRr7GaA6A==
`protect END_PROTECTED
