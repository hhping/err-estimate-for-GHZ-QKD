`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ObioFSLfWR5ogAr17jJG3/NGeWAuiZoENsd8+1PO4/xnzdIbuUoWxcLMwK1n94pm
RQy5EVQZXEtdUKEXB+SSpYM+6+DiK7pxiu94xUR4rS8IhBWnHX2fj/DMHgwP0UrH
WsT5XQTd1Q3ZcWrV9Jq+nVxCcsGQtDqhmRyJQyWYnrJ+qCZyTYCx7+eYkd7ELudr
zXkCbrIHoIiDzGYPQx+GBStb78fCh9brSLWxO6+vXnJX9Hk52x7R+J/MKVRZ2IxK
ql8QV4/R1GFm+jJEO664T9VeLxR34E3fFsIq44HibXZ4hf9NkJ5Nif9dQ2fNFkAh
pgXF3Jwv8pMmxoB9otN3T+kmDEoPl9Kdr3avg+tK1zjSb7ZLhfXkWFU1HuvpwKJH
rWEIVenYyyrZJlReEbeaY4HCd8JgpbJSxCl//6bxelZ5BBHXe7pcu7CYiURSHnhi
P861NIsnxa/f8Jn5IZOzfg==
`protect END_PROTECTED
