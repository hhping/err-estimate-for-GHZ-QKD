`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LdJ+FuO+9rWVP0mYdycOMhDO5EiTkuCl3HDpKx1zPsvhjHIdfAwP6FGfz8NI/Pu0
7Cwkd4gX35ugjK46isXK1bN1kfE6T2SeFRk64KDcuJnKc8b39JTGkKL1YzwLpYRu
mhQJdGLTk1X/V09VyOqouKJwXJFCSJzBmdWakYiv7sP0cjwe2U2czsuwkD3KgCQs
fH/r74J6Bw/RPJ/5zRF3Jb/61DJrB2ev1f7kuD80nDaFoqZEWCWmtsazdhgM+sDZ
mLixWIyhHu+8AuothHHgSCGHAtobXS7rUsvSws3eLwUQiFwWHfZPZJ+nsGaKnZgE
EUwRlaKG/iqlHaMVuuq6mJyx3BpoMaEmbEyo0e1myO2FMorBSoqUK0eVmuTZ4e/t
9rc1DV10mL4jDsXspdu15ZzDiyTXZDKLr3u23yhJVwEfFcPycYZkk9Q9UZ4G9wTw
8s9SqLcC9CyIMwYNTzxmBLyjlxcOEoNMSGD8REahkSjh4pinbK8OJnn2gNq9XkUt
5rkfgkC2hNYFhIGXSiL740uL2LQHfK5p7WCZwQlCzx/QzYp1Ew81/BMC5sjtFkvj
R0dkqA1WBg2DL8h+7d2iUhUbmEmL3B2G0wKznJLr30WODJpx5RlsUFDrgIEKwh36
6n50bYnJexX3a7rS7rftQQlXDwxpCEvcKbS4zlPoLbuOKAYyWrzp1QIROafQ1aSL
MTetoBOLk7SgJ/SAp6e6rHrol+1FfxJelfZs2c+IQ06RnQDvbjysKw4ccliI2CCk
43YtxftPoT+wl/WM/Ed/LTFXicK3A8ejHYPg/7K0BX7j/VCPRT8eoRmlAkZBKvaS
aZ/Saxs40zho4TBBgH1lq0feLskfYufi++M9GyvI2wYXdER4XDaiJKG9h5DvjMkM
h2JM+xkLrVTbwOZ3Ic0whR+2CqqjXlL0lY0txHffdoXiOJuJVNTmSCtjds94/TjB
4mHQFmyj3dnDEQ6lcJ3rGufd6jusQRno8h1t9rgZ1vrYX8RAvAc+j6rQ57iV1LOQ
l9zgJLXrICUgJUa8qJWq1tyRyghbJ7tQDa22EpQ2JQuLllcRhSUVWkMLA5d4mE8G
98fCnfNa1Bv2B1yrP/3EjUx68m3fGTdP5n7Q7VLsw5bttHWDZHxJRzUKbLuLlm3W
Z5b5B/iTC627TqdJO+3odJxDi4qjKWd2cqZ/HdcrUJLbqKp/nOJmP4b6woPLGP8E
iRBzhY/Xa3N718L+zayEzIsryB/J4N/epxwYMQXLSdRZsNpkiWZhZ8v5Xwmp6hRb
ME+0jKVkna2OwSNUhYVqjuwu7+Y2CnjSdEQk2rhX2+fPE98MgwrsIy6Aar/IhhqZ
UTqGEqdvgMbRdyGvf6S9PDSk52/PsfcZ0aY+3/yj9DZJqxllQ5jIfyYkxBnSdzcM
3Y47unEtbYzCN1JdUV8FaM8fPViLnfGstXXcarEVrpdjMDKt7ANRHJJG2rEghfbh
YAo5sSMx+BU4VYI6xBwRuYIMTBhAMgQVpNdBwIxxxn1NPhpKOydRsLOs0W0JhYlb
XAAmrJWUVuTOIppa03RyxIfi1SABCNetljMNro7qVIImiSCl2Xo5/D2Z69cQtjip
axmtP3lgWs/wqrl9/Nq5maXHmburJk/RwFHJKn+wSHZmSmeuSg8L2uldVjqwjCWu
QSyB0aGb5ULOz9X15UNIcVoWecYXvmFZD6bOgULllT3VoX9W8asr3lY6aJDRT/D9
mStYONODhODfB4Z3f7C+MSETM/HmS0CsHGB/Z3v1RrCTBVWSa2zt4NHY6fBElBCi
2i0Ga0HR19AZsnB0sXL++3rchLn7xPKfKndF1gphELXpI0bceIUqibG30Ic+W2CU
KpTVB7/i8jZ+wcg+P6n8dTgD4qFE85+5CMM9PsKo7m6woacaHs3ITsKvp56xZB1v
oGS/pJndLIBMUkpa2PmRkpBz26r5/mSyQPCt5MnLbMK6RuP6tghvqScMxB9L0qW0
8XWBLY1vsS7f5k3aP5D88OTpBnT/7rLgHQY3kZVTcX0N8dIex4PHyY1GyzZ0CdNt
D7+K8h2/UcAU1cqXgl6XNGHSn23Dba83FjRjDlM3ZmIkJi4x0Qz3/AaYcaA0ijO6
qyWCrB6QoZYDc0rUy7WAHCJZsRRq0W6ikmsecGPOjQdHz2Vvm9tgEqeKpyMTALjE
Mk5NzWO4vFbDte0MMxFReK9zrkHq6RdYFjFQcYx0Z0Hhl5iLcBFquKOgFk7TtPoG
RfD7wfNH+juwZ+g9qxasegoqe55LwsHRvDvSqsyB5JIh+ygUKxz1chY0q/CFO02t
ImBeGmwK2NvBr2qFS4wzTI99nkNxE7Yh1beTxyzF5mRj/I/qC/or+ljHmxx8b8Rb
5ZdIhZioDLliiCGP/me97wXE03XSbclIMNbeSGHfjn+Jip0Xsi2acJAZLG2zzk1Q
XpUFJPhTDIChLEwvXsY6LT+5yp7mnQmZvv4YAddNsHEYMT0Wi+NPmdNF8qXKqOsD
fP5lO6qDbYRQofoigUvps6NXnjC47m4Kvd2ib3xrBHL+hoa4DyPb+dEJ8981t1Jh
BlvpPewuUJj75UdcEy/EV/XC9y2+FSsM6PMoJwrzThTYA3vcD36l3V3DjoaYSQXZ
RVoGYoLRQmmC0KyLQUV6YvN/kUxwWE5CmMbIB0CR368TD3KwxzmST608tLNe8uS+
Ax4My0qEOg7ufU6bofLDl5v7yoS418HsXAY7ULQQQFDjKKq4evygq5BrmtsY+Bo0
asHi9ytC8mVSNc2YyTVTm7UwZtStSM5KSnRn4hOooH6fWmZQnfz6AjCyf9N/Wbsr
EMoAL009L9lrYsnbqbATpdMEJ+4u3qj+tQSKp0i066CuiTXQObEunEh3FzEtwloA
Lowfqivv7qA0pXFe/7R9p9pykldPDz61IvAeyo8uMaWKDLzdXRzZqlS344xrho4j
Q2ySJviqzxIP8HRj1DzNaGTQTc7cwHL+gVC1rV9r+gkoWYZNUNt1q35hUc5Lm9Xq
rCwnVMtRm4xe6qw6PY5BDiFkQnnwtEvnFVHgluU4ObmWl5h7yM87Vhrrgahnal4D
ltS7ZiN/1IUdsVKfxSJKDdQaVr4Rk9E042UhgPSASWEen4ei6zPrm4tupX6PVHqq
rBXEngJRs8xYX0Q2Gj7QhNh37dj9DuDkMZuTsBB29Ytps4iwBmGkn/Ubl2UZkrrj
hcxihOoh/Xi3DMsGPDiMw+nKYL1Y2Ql3W5xHZDS783/Q/6woJ8oWaNYIZozTFvKy
Dmj462ZsW3G8EiHfBy2kUnI00FEw6pwRCjZbOuumlw+2rsQ3IyA9B1wnDB7j4CzV
KtkNNjwGADHz5xhn42FK94TU7ys3GnHYVE+fDWD4MaAbGXpMvmE28us+5b6kgGrt
0d4H7TKmYbemh4TSHHIDjDSLc2QYuP6dDR8Pd6UrMY7dRymLKl9Ance8iE9rmGsI
9Hm775swrMYq+m+FPkVpA72KGNcHJaGd1EsgmHnh6b4zPkX1WKBFjjGpvmccwjJZ
ANHcfwMnkbP9moNUw1PUwjlfo91+fq8gdm7VXqPu5ZFKRygFPlHpN75Zx1rndIjY
uRs5kJjhhCDjQCg1oSetAmssdh5l9dUm5uZg7Rc13ZyydemiY1acR6OC07FhX33g
3geDU8DAWAn56jzdZ7/RAEPfZBHFm03Rj7A7jeDlhPOsN5WEWoYbHZd3VcAoK9zk
dDze5+OlUTSEHINTDmMSNb6Aw78ZsSb9M0urCGAa0fWa3TdvMIU6mkn36sHvXDCF
0E6nwjIFaUJj0N/KbsRLJA==
`protect END_PROTECTED
