`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHvFjwb4+FTcGmvB11V+zm4FiPLEpkC7oO0t2G8TVjN9uNPwfZHZk/AMU5Rk2zpo
qpxJUNOqkh4TTiRkOhmFBoccIhbPpMY+GUsq+yeSNqfELTq0clcrw8tk6Pj9rtg6
2mrSb/TJ73NqI/XLcLMRB+07915Sp3T8mKLSBos3OarCHIi3U7JX5SQaOLKymMQy
aoqAKF3oF/ekNCCS7DAqm6l6XxHiuDrg5odxuTvduw8C1ud+4R0svauWhBx8Xe/x
qRTyAPw/3h5aRm+9e3SWoo3Ie+Callimt1gJhbV59o3Rwx9DUMEGAhvM/U0vBvxG
iYhflpO6tqLy9SSlBlsjbYSZqU4hMGbZTEmhEtCyrInJnVUYv32wsLTYXBdsvMCm
oxr3EEzVLvMk4EDBAtpF6o+1sJGuhXzripf2DPxhxcD4NUWwQXpqr74mwNDbQ1f7
xHId+nj/d+yvB9rgbRdwfXj6v7DEPX9G0hJLFJnWdlOHi/EWWrvKhG3EhCCMKfBV
i4f3lGYZ8kNTvxM0nz0w1RjwFNrVtjlJB0VE6ttCww1lBpi5tDZGMuj5IUO56ptO
Lr5ou7tQepHHYslqZSosMUHLZKFoWlwLX5ZuNFp+584kdg/KntzjLZUc1LP7C+7b
5KuHrP5RHDfEhgvTbKuIqcDHDFhOXJTy69JB/2SVwX/xqqL1PDmYH0bAmLxqaa5y
GG4DgIyk42ASDB/mqATsqWzzBzvQLZSy6mCpdP8s3rjdkAqaxjBaN2xjXW+2JQZG
vAlmUoqfdi/Y9Ne3SEaMOUoNunjJ6f8fmejCjgfHCIsg3h7RoN+9NxFYcl+UNsOf
l3lHnDOG1yXrMcfCLpzEGXQxl2Jps6MRSdEcFgbCERliRdI4MUED+2Uiq4yrSp09
WVNPUDGLy1defnwXTK9BlK/eOo/LxB2tjfBFfrkhmQnMf7ULrJoVsgyZXlq8QFBu
PRfyto32Jocs1jo0TkxXueIXre6rAJp3w308jRsDDkRL3CE1m6fRjw0oOoqq6Hmx
sqgea2IDCSumVJuR3prw1dqA0Kkiz4/lacm4+OTYzMkXpIl/Qvfj5OPO4XN9xnOM
4+ae4S5vfpDd0RJnmVuvicQLcKJ4vJPAzEoef5BlZXSxmIT9SbBUJe6i9u2VVsF2
1gFHhWTLYOnhEfzvPiTkrlNUHgWIqgXDNixTzq140o5PvPzv0Kf+gsqbQpxsGQHK
cY+ITHq96zCqO4wf7ufD4q9lbM0rSN3tGioyM0NjZVj+jU2tW6JhgeSKkRChZHRA
jBUPFoZKoYcZ0lpWBqP0Re4ijg0zpLWRTTGi/e8ktuDio1CzV3HO+jD1egjHLSum
JzEWh4MA1fdKbRZQt7K5qXvgxvXvqoVwqlotCKZAgrMdtzQxniMbPHvxJXke1ITv
82Ig0zNwJy2yB762qmp9vw==
`protect END_PROTECTED
