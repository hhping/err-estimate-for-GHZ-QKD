`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HR4JjSh50VB0A1xIFDgxsqv7bVoBJ+t8+aas95SM2QtTHdnF275ZmtLfzs7oxJjC
vvT0+VDK4fQlM3vYff3xloNWVbLJhkZnbsBbQfKDzSp8cr1lYquBAKqWodG7LC+M
mj62L4utPtjTyZe7xIE7W2JMk3uioGW/kHOAWIZjGCr+zAbBqWAQ2uVFrxBMzLnx
TVqZIBRAiCnBiGR/arJAs5xl/z/JjOUN29sRoivLZ8jQBFhNV+6S0ZoV+bKrx9cu
4Dfnp8Z3Jz4Wg1ldWxuJIz826zxL/YOtnVXV8Lf71A9nTJak8Lg4/lHLZL8LdMRj
XomYBksUWvz8ieRf/bwV57fkmDGmEP9efvQNT4qWg1tBAtSmYwje0aHy/TXDo5IK
stj6PHyasfT7p4V3pBfWJNPsCdHKiDEzf6dzqsoECSOElhDIXUlHWJqgC24IXPbl
e9kampwokeMUp03+zYXiOQewsB8H1BesNHr69V2FMsLVcZxYnY8XE0MunmDgZymE
PctZsqYCo/gi5H8wjZ7cpYeqt0zKwzgwuqrRGI/YJhFqcd6l1qatnT/jYPlsRIIb
bRqqBuupEt1lNfuCrATWGm7Q1rnz6BHs4TreSAkabv/tOOBI2oehrjh4fsWqlev/
L64B26NuM55islv80xln9YjdWBQuu/htXW0Xd31ComuFyEzLtk4tGbmyTClw7BkL
EtGQmVHdg1BlxQBGm+tV6SSMi+22B80jDPT6FVvnNmu5V5o5BGeJIszi464er2j8
8jLd1y794yIFuXAfpELFkTqN6M9XbxrHZf4TfuW410/NIYpctN+mCZjUWjX/5a47
BjAl5TnB0leFrXwpoYJJw+vqTycpjuKRrDuyBKR/6cRKmnXAtn72/ohmF12Y7wdK
jEShtpOdxbUEZ71hPFzEd2hMYPxlJwve2sJz/q2/FqUnUlMD8LWhgRXZjoqSra+P
GuldnhzVsDF2Iyxa1+zvXLF8d9JGiNjoRGy6egNDDJviT75O7obM9ysMSPKtRfTP
hK30dhIjE90QnV6goO9FjyesuKM/YVlmHWTyiNIccSPKluHdYXAKU67DgmbqiM5T
Ehzob9+q4bYu/m0Ldn9TQmictu9Pgn4AaI1NV+TKQAVRqkICredrwgiH3pnpdazS
WAqd/VoAE3FKW93U2UeaGVS+3MxvjCniuJLOIQsIzZoTaAbm9taMUunpmI7hpFDW
Q27pBdDWCY7cdARQWuNp+daHw8eXJnldQgncL12We4gzORkMXAzCOHIrsmUuWCS2
cATLUVcrq8wzUM4zrICbj9riMVJg59JG8SdQVOsiiHcBm29rR7ux4T4+7R72pQCu
sew7YGhknruOdIGz+cMlF5F6qfIhFjsEqU9s4A7kZ+ZBaQqIuBXl4cF5IBn5UrH9
5f5My7bzm5bIAEmP9jjcSvps0UxbcOlv/zIsuSesSNNoj7lJrbLFY1LolnpfuNz+
hwQZVjmyrSUs9Y8gmFUtM6In2IwB18WOh/A4IIiotCRo73nDMECowYP7GQhrzJt/
mblSZDSIsBwet23qYc2LRY/Rp0XGFdTraOKdMC9GorskmUIbWIvxgsR4lUth8JXX
3v8SfArwHisD/IYa5L4jI6ZZmeW138ZmrfacBPUDvQ5G/0NFVSRK3kD2/r1imMd8
Dm7YfDlCkX3KCoJHWVIomIblf0P/bnNdOc5XBjdF0EVIgLIcRXpLUlJgN1kctKGQ
Nd8RuaBSQGKWDSkXC3pjUYl7ecwdt1nkmIOzzpqQl/3v9aGW9DogHQWydrytvgDh
ecXabasP5UjAtxEmklyy27rwnUuYLTItlsmK6whC7XteYXCyReFOkbng8zlQBpah
iMeJ2C7tM2lwkFQrcl2V/8raZRSOlRc76V9atw2nbe4U8sTS9COY4MUyC1U59PLI
dbEnH7NUwxlQ+4ivk0fAgQ9Or4MpePXAwvL+6c4CSxzoX+br9LxdRQXYJp9Z2qXX
fh31tYRGveNzIoFVXMYQ7kJzlvVFdq1Acd3nYN/e9OjQQs9/dDqIO3Hws1cNVHG3
WRG2aWyYUu6R14kFnO0J4NaxgctRcfecl0n1GXRvOQfPa4PkpkBQxo3qTHcLIr5j
KH75do97/0KvFQKGGqcaiA6ENRhSaLOktgN+8RtaN8xrkg/fGBMpSYULblDE75Lq
gZM8XaR7JkuIHTZEa8UT1MkR7nRdsOvh6eRKcS+WR6fUzGCDhqaetEi5ZYRRnGfR
e2TYsyQ9rKmkOscjO6cUcxifdo4mOlQE4/BbNUOCxFYzEvXp4Dp3169N6EXkb3gY
Kz1GXBfVHvBYG9LfKL9xU7s0UpZFlOVBfTne+jGrnwkDM9yeFZWyqpyw18pf0y0d
KLs7MX4aouTjFiAQpJL3DQq5MKtFAotH5nPHw0DG66iHOV5SycK0JfQBodNBl7/1
UDsn0HjCbg65tPCnCxTkPkpJU+svMCSBE5I3f3J+i1a5S2FPFv6hP69R/ch1e+ol
gJHgfYLwKFW2YmfKM6HlUvZOmrRMeljj7I6ERrd4TZ5PDJpHm1gW9DXF34Mg2q6c
3bssw0q9+9XMw0hjySvlXqxA1XKmrpj7HEgJGDH+216vbtZGe4l76YzILMbFjK2g
SE+JeZIXAAMNhiWzCGQ6ysRUyc/huN3StezHJh17UTt7ZdFUphUfsapK/HSzMIlz
/Uk7byrv7ivN8GDaiUu72yvtEfG1aIigLmRtquuzyI9G6AYpM5KMoE2D5IfodMRL
Z8M5WQUIiLaytvF8xofdXWZo9sC0/dvCDZBRjdXr/DEmxnFTarYonON1ggbEXnGg
xOzMvrSss9rLksTW06ztCly8RjB9cSqOK4mURfYj1ypR6LDF2uOhsGxSrQTIGX0D
ntq6K02NzrPKoVQ6vLhtSfP8+ePdooRHP8FjYlCVO+0aIPXEVuF6O8P0ufWFCrH1
fZxumqMm5gMl3sbIK98nWuhXNJlmYP991WYoZZd7vhxIdrbyM49qqU7p8Bjk3P+r
D8C2QAkg7XQx5HXnzAMruv2CNPwxrcXZ6L/3j2mORKFgJyL41kAmjCVcqTTnUd/1
bQDS831aFCUltAyZcT1iCjqwW1T/6+pwDCt4s/zPCCZyh08TxjbWkloS1WYl5vqH
Wbs417zx+yU/MvQGb4h2oYdN8DEJrrSrsn3mfB2IE+qaozNj7qAWiqQz99+h/X+c
JawrzItrIpnGDDGTB/t9BSMbxzJVcwj0/d6THf7mFensSQ94GRh9tHkYMVOnxodg
we6dP6iEU73yIQCaUlH0KpftR5J/FbJyjnCFk3axDvQK+s/BRT8GZJ55ZIlRFfVt
KzajWjB2eBqcOjEWInJ/I0ep7XEKvsRUeMAhC0AUpXl8dUUMxVz2dBSlNgvfelph
u4fZP2zkj2/j17JOViErjxt7BYagts39qvXaDiIz9XukiF4agPCG666hB2tvY25a
JQ7sTeoAmAo/slL0ubnBp0R8mgy6NchD/CDNGjeKm+qPyXYJlwlNWLFWBFwDMPuc
a/K7VvAHQMiSSTD1zv9PBpanG8ZGJMM7iE2F1E64QOKbNbMru1PWWGDBkEljSyhO
SmLFYdDBphk/4NhtVXvcngNI9Y9lAq1c2/iMqHm2RiIOVsooot1JIlX0t6I9oH61
HdOCOv1RfOTRbO1sTKjy1W1bKY2oSto/keQC0V/jFQXqPYQY4kxlCekPZGm6kMCF
zcTy2qv3aeW4sKcAceQMKwPQQNyZQOPtWJkWuvViUoWq4li/HjsbP3qUF5hDtnxw
bpN7tUPK2HnTZBBkHkPdWfP4ROWtiR+KXUhm6drXb7cdChD+B/gp3olDd5Uc6ISw
GEKKl9zDBslfyA7jQFntF0UpIbP0+/941MR9migzjNR0E8CCyXXWBzl8VpTaBOeB
QnQ3/t8izwZ+ihBsmjTqslL3c3IWPbsQptYOoApcU9+4cOvtPrCcNbiJz9JbK9cb
cANQ6VW4d3s1mKZnGOcaqPbwihitjIQ8YlPsNznKpmb9+miV7uL63Zq3jtUMltXF
EwEC0fR5u2nsmZewPwiabb9GuIUqUlmJHryN5j7RhCaHNp7cB7cj+8Y0G1ibsEBp
zb/eu3CjB3czzgaT8cmNPbGvRtiVUYh+nEwb9woHqOoLTE9AN2cyXpjmBKz160r+
ikUZbvAFNTJFgzDO8b2uB67pjT327XtPcr14UgThHDF1BvgmP6SaKeL4KWX17BWg
Nerd/J26GygBJB/OroCdcP68LHZhc+321ZocUZoUeP8H9K0CELjPMyCSoHgRYYfF
fglHXRnP/VQlZjak2YeCpgCH/xSQh+RDWNZFiYB9LQwWxV6QFxuKPf9q3ZPH2tzn
iO55FUI5yng05x/Ii1ggbQlL8wDkZbh52dS/W9GcVdK2s6p7AUc0zzCJLhT1PrX0
FGGs9VKGb8nkoVjPf672R4POdFJbJZS+yI+rH0VRvjVhory8wR2gms3hOtPrxebR
s8/dJR4z5It1d+AmxcpJ4W7d/6O46gNnkbHY91NJQqp4dau3ZeEMHhSOdJcJalyo
`protect END_PROTECTED
