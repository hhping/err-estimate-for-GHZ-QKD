`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDlKOndGxB8fihsO48MCzp0ATfQhXscNUxqcTmYA0ZRYz604gJczYxmUckVrb6Qs
lUrTLmzy2b6dVPczyGZbhdHSM6Fx8ozRKwesJqlcfo5FJIY3JMlkmycVwyJJPiZd
P8QShFNzwyZ4H3KerctnTcVOz8UmuIHjJy0xKOCW3KZ4MaXHT7j30I3h6LgDtQyT
OSYTQdYw7Wy3KSZn77WL+hgxoxLpAwpHXZ4TwksqFR4pvz9zVekprHaOQezpV/Oc
UI0ZI18rZIyHSKoH1SDGAvG8oUYOsb8OY0s13KxA1+hjXrpr+hjjgy23uEJEJZ0d
LlxOoPgdxHafVQ0aO5p7DD6Fx4hJbtvdPXqZpvd1gZ6dUElcyuI9aKCr+XbxXbCO
9jwMjJJ5MfFS9Vn3m9jWGV3qngLhePH62oSsYK3nPX6YsIWwXLfRpGVGTMSmysXu
7JOHVEzOLE6n1nwDCIZgOULlfPGozR2stcewHcZwju3NpSNcn9ed+dA1e5cn4zQt
Lsr/ycsek0nzCG3hnysOd9CS50SITwsdsiSpM63YnZjSjU1ifJ0no/bf9VBYMxnn
5SGTnlx3N2FxlkdOHt5jv2tK8Ck921aJjEbxWd5+MqzSkuzkuH/dG4P/Oh6TaBkX
`protect END_PROTECTED
