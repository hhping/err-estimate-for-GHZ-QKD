`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mXc4fGDqltClynD6YuLzqPxMSfktzqlguPxPoTcgAyFff7FcZVicgJxBsr8x7sU/
1NvmT9LSzQucV+QbQgYideGHKqs/3t7qIiMbmlCLFXPzcYzvL4EHBnPmcAFEZGBd
zj5zxvDX3DCoVosnzODHq/IVq3A7l4dY0PIoXRpgutnzOHBk/goBIzJzI9dNdAQF
DY0dmmBTIprVS+5CFhbzzmVMCcA5fUeBUUJ+jg+vORpAJN+At7NXlBRN8FUSldO0
X9Bt6GCdn6IPM4oGoWvmi/Bwbmj44uXzPVJlkwOQ9vh78D0qyOW+jF1fC7wF0J8+
IZack+L1VhpQmeJyb8mzdR2WfTfsj+nyqMDCJA2aO4QRLR4Pms+oJfpKnchgHpva
omlCgf+bBeSg5ggVGltZwQulBMYKzfXE33RZG5ysbnYtkAElH7eX0M0ISdeP4ouM
5ztIjv7k2A9G7ux9+QaHkkUGvsHZHGxilQiP1MfzAWkI/uduzmSwoSBrr6LK9r1s
uLeh2I/VQ08LgHgklES/UmEdQvFPllmiioanrmNfHZ11+1gIO/Q9KphsUXjGcZwt
4QRT1ErKeK4kZQVGY7sau/3hSEVF7YWeKlXGxBobJcE/Pia1XZmcwDWYK3QBEM4/
dMBhQK5QaypV5SYgHQga9e4i6ZFkyJnGgvrPTzXjPWmdhiBObEWC4nAkIFJRU0dO
2IEkI70NKGdDhq8gWJY9WeB8MmZYmaid3aLdDpcucJKSkx/1wtGesoow0Hno6hgf
L858bFehJBARK4DNdCcvJdtijYgHsHSNnrqDkfcRDw1zT5/9wR18h/+V84RVC5J+
k6+YUbtPaT/XOgv61jYTCPuD6uasjpG/FkX5aToDTMxuxTutXKLL4j/yUdcvmG1/
3wR0EOpELqk4WsbK2Y8F6+yAMzSscFM+ZKGQJMXg22w7RBI3zRHzNC85sRwGdusB
RV2MuzBu6jpQY7Ja1Xq9bCzDPsSEJqKhbz1YwMwFdsZ2p51KtG+mzvBQOlX59KV1
XoWLVcv/C9jeu9tyM5w5aEBsAS6dLw5vnTby+Qa2gY22tKj2ivm4/jdl/QU26xFk
KoEEUwG0eMHqnQvsGxbsvcLIc3Eseo2ZTBNZxlIiHy5AybCW808enrPtZIEYMMEs
Kkw0qC5dYqSd/jpNUZViujrEh+GFPfRQlmmFIdxx1D3YbFoSZvbl6P4eaiePg+8k
WYl6pQoGMl1zeYuynmLSKsq9hgEYwZT4EK/2hPCHAffTCDa6v1eQGyamNhFT1oYP
uFcajKD8EW6HpZdMsIPA+/R2NQ58YWhD0wG3T68S0/ZTwk4ZIZm4CX1PkxOGu7Eg
njBCgBUrveImaVcsJoV9wLMIHp5CJ38s8Pes0rmZfFEAZrcYORq30da3QmoouVKS
tk7AMvAnQv6Pp3pGMw/8Xudd7zEhUWFUgHhYEf/zvOAPDbbDPUlBGYDEI2y0bW03
1c+trC2uDUOYnML9xlHOjvf5IjvdKcIZeDBcmxsWaEotD0mOqweemtsuAoZoP2OY
q+u05hZdPYF1Po2Wqp3dHSBiKy+jseA18Qk6FEpbH8Vbhi7yRF+YQUWB7bATSyCb
91Gj1FXEt2stoaSJStm8YAjL2pLZFtudnVdWUVqlddEH1q9G9GnlGLbANs3JI+Ol
06oROT4bwEggp61Rvxsv/0h631sssmOzTIuSMw/6vlAkIFz3al6PI2a2dsYmHfgK
4fA6v+SXbe+FX0qL4yNISpwo8o2eS4dsGYV/BY7Fx9ebWleLp3HYkglOQV7Zj2ZA
Wl+J+OfcVkIEG2VD02JhB54ADrI4H/Qm9wrgyJ5VLQfIb81UJgJIG3io5WK2K66Y
QDt/lI78mKWZR0iENqmvbgKXdu9pp+6kNXrIHh+LI9sxcQOc4CIq3ZHYXEQg2A2x
tkqP0XFSnFrZM2fCeejOOusoadRabjWKmtNz9ucOslGPxb/Myc5hFoG/IsLTA6bZ
NWQMF79za6At7Z8BdYBMCw3yR5GvXAj8afFOtGbN3fp7/w5UpFPOdp0RWa/4lvMS
ApuZNDQZxSbYJcLEejxIxKIU0y9wzXZuw3D33N0y0Mk/8q4oDVVwk2BTQ1ey3Dbt
kwRy77hUyTIA+r7epuhEoeHmiMxt59s9old0D1Py54ODZiv5tONR0oxTOUCFqa7U
XMpw43jTf+JEPXpK/Hjleluauy8OTTHLpY7t0Y1ntapuDMrFqOsifJ0cuGxuqqCx
O0EsLuN7T+EZvakhmWaSHHno4yNetCQjstSGBrz2uwhctymu79BUU0uU6ocdrnA/
sPwVrVDOT1cQCh5doNIw5ZNy1r9IAVWhGE51oCEPdkC921jrKl8bX11hET326kr5
lq1xEeQ+YaFvAGd7WLr+YarvhYmOJzGwLTh/8t2IzxNSC+ATQK7WiKuLma83uBBK
i+Cgk34y1mCGpIJapIGjTLZUwgnQEjyoX5xZS/paWmAylDAgatifczI3U6g6YWA2
jPhSbB9lQVcsAZ+8zwLgjQgGIJOEPMv4Wm76q2IBbygCXFXTUe803jMOzli1gGKq
IdDf8G911zvH1CG+pr7JUqGVjYvSQwne3h/gzqOCWR5zW8IfMRtXCvUP1wk3rjP/
4oguLAZTTEcDWImU0BiEynMBaDb7RiVkE/l0XLq28jQtVxKp9YoYm93+tGEyB2O5
CSyTiABhiA6p/MExoSBcXSvH+QYAyCg5tal2QDyhp1uXN24Bi3JRzaE3al1EOPL/
xTD6VB6UONYRhtUZiGfcBjIivTLzRA20FH/lupxYT8ZpFPSxB3tj49h8Y7qrSqnS
r4IrqicWi/JM9T9p8MubXs/B9U6ZUT/zReFXxqlQ6MA1BBegmjCbYIBoRixuZmQR
MAavzDXZz9lRWjVtW2/fqRuV4Elzr/THk3YnK8uWpDkUngApNS4lsSOQxYI+DbZY
5GdCq+cXgPNuoq4rvJ7Q2akOhnuwbsUrV/++qmCRPxc9irCr2ZjvCcUqk1U5QEYK
qMZfNFIDaO5qqjUP45bt9B0KqsXNq4Ok2g6jKWbZbvX8tnRJERLu2leSuQkkPnkj
yEJL8D/RmIqF7BqLMJ183YVn00ufVv0tMUQvn46cd1hZY9nUe6lSzHI3ya95vafP
vMSiul07LkZx/0xdOCjLbuT3m56TULEVVkWTKp9QmapZ8L+CyhMCzM1q7uJ2FBJG
MXfz5twbnYbZpaDcAJVss0SrQ4eDmpsMT8Zo2yvgcmHDB33TlyVgu2xjjHqPnV78
0B31+EQtRCkI1ysHeT20sFGc9R9RjE1z3i3VHPKUASMoqdHOdrYZBMSdW4t8R/Fv
W3B5zI7KY7efvpb57h4y0qkC8Eev7uxZIOXs8bD0c6qS+drB8kg+zL2Q2m2+u/WE
UWf+wd6HQo+nY5ENaq5aFbu+s1RAYq0Ypir2aHoC1Lb5RVSkseqjyydiLrQ4Lwij
w/8RnIbkT/x1UTpsz68LVlBK1TQ28I5721LnKBkFRkQUtYxleGxUOB4o7sPr/RrQ
m1lKsIQBdw8wDQpZ2LRhq31fcKlXxxYsjTX5YRy5eBaP2dyDx5zaGgPCEEVqm4Jk
IaAfd6dxWujJo64DU4bEQrnCPEk1VBtWJCXMyASB1uoi7qLcl/SJ0Ks15TwZb7O4
E0EIz4tcirNLXBDKXTvdrERyT8gAG+UDBf8NMH7Bo0PXmCndAkfXWxbgbApciRFq
pho3XTK3TPCPXpK5iijS1SlrF63ymIilixwLhFdKdcAHfHciIwG2Zc33tVnu4c9H
CxxkpUmlNnx6IQ6PPoK2C3aUy3KmSAqBSyQxO1x0tutMbV0L/ejdpdYaiayRnoPT
+rgin+2eSXxmzX+nfNsvwglGvyS8y5Hp7kxUbZxvYzylLU8tZsi77Cd2ei9rWBUu
s+NlZXvi0q7PLNhdrBTZUSypEkixgp5tkug+xY4p1b05VGrQDFN3vLqz0WwoDIgn
Om9lyEL5FZNsyYtYhvfOPbAk60oCdkF4YP0SApzIAMWchUiDDniu4bLwkMixO7F4
0vMVsmWI4Tca4b+1QuqGcdRXKtR+j/b7Sqmv+UgCA0R4w6I9L2V6n13JafBLPMp5
cSrPkKXctV8xfDF6aM9jAkk/Z6Hy3F2qU8rKOFNlnwEs/BlAIlmvqm/LxjI5nFqR
y333ugxU8p57S5/Du7SmveKu6zFvYZtgvAcqvedC0pyGYBQfe0EkONrjOVtvM1ky
jtDNnhYoyVTdiczwx88m8Kku6WHobeuyp4wxcggFt4smN5LQvbpXghN7E5iYrJUy
3eqhaiAfrl7KecpayMjJXqIMWS52LzoSE4CatUTp0tn9vdvzIPfXPUfbsbDVRcy7
G9RRefsmeIpiecV26crD+YWPY8qUH4Y7PN5NjUHS0DY5GAFNZg503BNk+1agOtJy
gF/CMqbU7Eg1M9IoGh5FtnIDlGp/6MhHkv2dAfoeX8y4IG8vuY4xgW8rfm1IFrtX
EUDJX9zolkZ48Lq9BXuK7gvE2oRspR+qJaKEMztH7Y+TeUjiZ3SCi9Zaualru+ng
Ut5OIfBWtn+muD3bCq+lWs1XPWiTFWKwe/UY9euxVFHigTpWWlmyTOe5L44siLmW
VDiLreUSvl/zVna1wF/hK4Hke7qHzM7tmRsDwFADRVAGPnzARQZsSxZdZHHy9QLV
6Eiw/8FgRisHAfzbeH/knoN4pengrXu+22S9SAsVzUnPsugfHNtN8wKjR9Ug1Xj9
foDmVI/kKliadYrVmllMs0mqkd6hopEmbUanZejwg1HbCNGNbW+rsYjRMJqokjLK
TO+1UaFyMknev6DItROJTGHpEBJM1gc2fjA6lgodjU1/TxWQPATp05CI5+N6m5l6
yyHDJkh0acy89oSn8ayF9D2bkk9ljSMkDOITcZydIAr4q6bEY66M3O9wnFf+49RW
ErtL2hNP4I7ZILmPF2yPlwxOCljgDRH2sMVY27jtDL4/0gkcJGgt5vGRMFUdPr3u
YxWed/FSvvZDfa5J1qJ5ZwQFU58UNd1kkw7RjqCmNFI3/NnkPd8a1iCeI4/ZEFQT
yyOttPQixZfANl8xUGjHAZrawdoakSBZg++KvI02fO+Tzf6SY0eUp8LXD8YQs5Sr
l8TM7TPgQOsK+SNCDGsnAEOmI51jt+wL+rA4BsLEpJq+1jJG/augxD/zxuk6r7gZ
MvQv1hrCVnWi59g1rk0iJooD+G4H8nVwT+AEthwdEdPzsvV2O58ansJeQ2NI1z2K
96vhpSWTTdhrUofXuusjJEtDy4k94Tyg1Nmd4gBshgNS2ARIPi9lQC5plNKx4b+s
FhdZSHFjf9ryQzCZ9AIJP154/QnEi1X19CFV9RpH04rkiAxskdmG9PWIMxsrZTVk
/hDZSQOx3avApkiQLHRBuCTApFVICvbpr9N0gdqOj5KImMomrvJ+Yf2EdNS6b4gW
XmLgZnKaZB4oTtz0c2azqwKAdkgfe6mgCptqLsUlyp+//Eg9Ri1AYRLq7GNODpOL
JEkeIdIorjWLYhq8wEEgQ3JppsruTd4ChVjp0hpV754TLhTFQRUcB90rbceJ0PmO
vp0eBwOMDIKhdWZof1jG4Rks6+3WKQJuwHKwhz1aX5aJv+oKQKC4V9ytIeWy5w/Y
eFOzSnBpvZxbH5Sx/G6D0g==
`protect END_PROTECTED
