`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lRY35WMaTeDJN4ZDeA2w8FF0rptJiR9fYUGx/iGpqed0qukA7+ysHD8A1yPGJuXM
eQWOXB0BYpvPcO+/6qpTDhSSjIiU1Xv17jxkh3uU+8zmApFToofB/om1isGZlnjp
f32jp3pWqCxgs4Aajmbpwc+ox6ZmuOTSq60wCef0hoaqXxsmFRa1WtOc7bcFnSEk
GvfyLQDK+fmLPIovq9D8MToZkwsgzORxpnykM0h5Pcd4IeJjqM9U1wIEAfNPpxUJ
PtiPyVgdKThl+XtkGm2cixUR4QknQUH5gLfOuAc62q4MBYtBVD2xLFHlrR0fO4u/
6Z9MuY3AuW4UQHoXgaZ7rrjntkI9HdWrp9DWFXo6eLwP0ru0W3qNA2TWKeEg9kod
kIgq+OuhfNHqQnCRK8aeFecn8qOOSHlEPQsfpl6k6DxeggPVN0uXM2ttacPxJSrs
m0tutuw44NsCsJL7Lvs+NSYiLgGjv9YJNvBkTKKbBDexN0N1NZp3j5rFGQDmw8pQ
Mbf4Bm0xcwBRk4jmv2FthXS+S56groBE7gqDhPhKSSpIDcxPuJG2M8XbN0gtNfgV
sc/cF/TZ0IUyUYGrqF38n2ijhCBMRTQdCzY0lT0eFagMWJcynzjPgHGf6fQVOgNT
yDuhl52x4LE2JXOtS84vqrXAV2LJCuCaa0ynvKPKWYCLf3JRvSY3vM9dXvgPpHY9
HKzbPrh/Fy/7NdHedOSungjkWjhXzIaQMjHkNwtYR8eaQE6kE9xW8cZ1I2PjJ3cK
SV3UHxNROY5BhAkl68dBP+JuUmamuVOZ6ycIejgKAYD3+QjSCjDXOPyNu3D2QKnW
WvzU30FaAK5vtA7n9jllcFar66gll59wmTjnSyoERkIamZTd7cNzW3LJAHy0dy6l
VHkk08sAspTzb8btdv17RNcS61FQZYuiRQAc4Eq2sWzqa3TyFm0qGTAYB8wcbQgS
PFvKPDEWMIWFEqqbZEXwZDBHXon/Xprstvv7ssOY4fVpfRZi0UPlG3lmV5MkXiCt
NOrOH2m6cseccLgNKi6oi70am8IgbA5IBp4iY4q3nQGidtObNmP7MMLMvoCTMmQl
D/u2F8iK0J+W49SZphoSBk63hTDwZMBK42DvE/frPyfy4Tp7YBOo6p9GApx7lcik
YgxBh0ci7IgjPtYBPAwb/NLrIno2LMPmR/Tg1reLjWSl3fvKGwZzbjxVujAE0zcW
t+rvs6fZd9WNBL1NA04+akubF1CD+istE0RLACDM/k/1ZChQGGMATpkc6iX1fY5Q
0RBhbSD+iJ6tftuI+9kcpN/KojxmmwkWF+MV0IBjE596eXtEVGli6XqK8IvUxIcR
lVPwe782+DKPcLuiCBWJ9jMZYz9V0rrvTYGhp7iLNSeE0/cpSvOit/j0SHc60XMF
xNNbJPEJH+5dKBNxJr3UjkCRUo7PrCu0plD6f4HeMmqsP+IjMhzUems3Vh0pMSHE
eoIqBK8cn72WyiSpBkYpRKln5WwWjzMxtR1M1eivpoZjWYHns+K/j+LblGgn9M0t
+dVqYmtVYpgsdQ/8Uv5D2pnSXM+pJsxAr1OEKewkhtAqBxnqMANVV81VRIAoOflk
cB66JaYyGq0Oh00e+pUMbfSRZ/JU0EJk5dXtN/nZLGp2xH92/kHOmjfwPxVNYBhg
95g/qzKYKyWroWs2khjOpnQvMDalr85hZdSz5kHJF0P0wPwlhh575H5qYpXC8OEH
p25WOMr/qVrq+gjU9ZLK8UbUT6K740dxXgCgpepF/8M4p7ZF4EPXBDxh2cIzmHFO
7WUdcL6GaVkQHOOsnvCQCmjjsewhaRtAoNwBw1PJuaIHBzmepO0lKk3kZN5nNsU2
tfldMR6ETSyeTV3Urk8dl3boQdSfQk4OXonbKZ+AId5iC0rIbKpFP+pfS0Z1iyxF
RYv2J1ykewm57u+4Gam5W7XH1vPNFcnbrWDgYq8RG0EHjnOzQbD8+bdrJ/ZTteEf
l8MjXob6IXdrUqP/Ii+YpF95FqDCPZtIuUKr8pScM499/QT0uy0asf+zvi/dpmII
KFZ9XrvNFOb6/9kyGfjzmPGncjHx5UtFseFklxPHed2xmzZJPIO+q06+23XlOcQn
8EyK5Z9tyqmB621TNMuXb7WAQwU1fCDwjbjFlC3Ncn5L2tLN4uVHBbtnoPAjfjOe
`protect END_PROTECTED
