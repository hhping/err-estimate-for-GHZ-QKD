`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4TdkQynQlVu3aNelSh7RI5ubkRA2ia1VpO4BdvE2VF1UBBUBkUgCm1unmp9tgOdf
RNaS+EBU/VU8QEYCyjzkpmhFBHzvfZae3mauZGPLzei4QEV96Lh0+PaM8BFrIX7X
Lsxi27dxaOpz5zmWdDharRibhrjg1TCYXTfHnI9r/Y7zxzOt/Fp1eDiCao0xlmje
4tVnyMi7MofCqtDzQB/Ch/eECNaOwVNrXgxfYOvwF0RuvQAqs16JsuXtfBo0iJl2
KHo1i1aALNsE7n42e+r5/gHWFdliGyvwL5BBQngH3WeV1o6QQVXHIwSxW868NDTx
7DuvSugMbrFFbuEQMXJbQBoR/QVV7f7bXCa8unhYznJnD606Ev9U+UNubrEK14cX
eRX6pXPJ8VOTfJnr0DizNq6BTsHcHYVQ3FO43SXULXXyga/Lp/OZs3l6Wb440Wtk
emmWgD8heBUeHzi7qO8Uw84c6GQgBnJ1/U6uIX0QliM+wzBnc4qbbDYGibNohaeQ
j/09aSDYgv5jtkp8NrbSNeHRjACjxjo7yvxA9fb8n3pyGcbzaDZOheKQ8przKWd7
9l9usOm+DyCR05DzlUoogZoF5x7VUEqYEZsVusXVyPn/2AR7xtrqmAHF9v6o+lZK
6FHJDQaokgY2LaJj6+TDnds5mLoSkS9E5vr7+Itaqr8n7dl/Sonde5QWjBnNlGYp
JK6wyTW/fNW2QzW5enqNm9CVji3AjEFVyXtmcAqXbJqJ4V+MDJWr7MKBla/BZnDD
63mDlnghjld/hyJ0GluKiE71WAImaefnNG3I0VOWtHLPdxJg/alj8phWnQPFzbA3
tiyu+jAZDHFzCehpc5/IVPV8cOMDirlnrMFY0t+m61e96lkgS+3qh0AgUSjapayY
Ujc4QXqpEDLDIIbSjg9joYUA2NWzP40r4c8+QkPOgKTG2yiVc8zNRah+lF3dCfcM
wHvqktUXz2NjQ+xA0x66dOLZ1mBnvoIQJ17CUdH8CGirR7XJxOB5vIrEfnVq7GAU
NLPIwh94cCWTvYD9T/0bUEuy2GJ1OA+7yKds4Bku9XKFH9WmcuPNSYRJEyxg7Gen
xz9iHgTPUt28Nj7gOU3Q0E2+bz+KtsQ7Yp/u5WVfbTwiEe3g9ZnFXa4+2PzXrjCN
BpWGRFReScjgAd9MOj9e6fMsnbE7fEZldC1cS0nm9md1l2NudUoiiHJ8So29H+g6
A+8q1Blohpv9ztwoZlLGdwy7GYx1wc17UsMVVXDbu3lE+qPmVaRAtg2QN4irih1A
s38KJRGQs+WloOL9IHkI0hDSlsAhz6OCNMvwpofQKNkLXkNP65k/uGrgxmKP1cQG
xLT87mmjLpoMPSEFemnHtj2+QT6v6JZVTUVpoOroicB2wGbBGjnjaZH9h6rvQacj
dlqyiISrj4v9rH7nFKe8KQr1JQPiUyjkCs/44kNvdCAc0aH78JnwNY/QbsW2k+0V
bC/IA5dSdTkrMBOmtK9xaC9sFK2BMOoo9qhud3m0cac34BsaUWlBjNmuomjKlZce
gd8/9sEEu+H2ra6ELLFk9wAh9owBCkG8X0pALlym1pL8WEyEh+uQhb2j5k5m7hft
BTUkyfQ9IkLwxLUYsh0dnQ==
`protect END_PROTECTED
