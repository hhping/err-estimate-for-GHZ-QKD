`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Y3oKcbIwVdnqoEyTysUX5fde+TdDpYGhwScca262akWHREf7QSQhjBGN8MS4sAY
pJOzmxMQLkHC4eKYUvWd1ECCxPdvIkt3LrNM1h6g4kon5B/BiqIni3AGIs5XFjCH
Rj3O7XxW+HEfWobBcNrDnmpbRJPG4H4Nq2KFuL2D9aYhtvCRIX7m8p6SUlxY8V0P
syEVqshikRRZlwatmCbGoQWJ1Isi5SezYQIUwiBHP92cLqUCNcOCU6XRrtl3ejXr
zllUsby9iwsFaMMZfjWpibGA+yHoj9ioOnHhyH9pWWIm9xamICEhgJU9jl3Pu1rS
LtnqE10gJ8vfKHwG7pRtusLtjF6van9OucOF2LFAh2KDMa5s9PjygVf8OVgrMOyp
Gvgo0ZIgWcjRr1AgIji8u10srMJujTfQVrRyEOZ5SzoSTKYXcQj5B3R5ESz0tZYo
WFoDGu7HiaMDkN5C7rniT2dFyoWiPrBpvL/bfqfX9MTT3jKXXRAQvBP16R+WKL0a
fk/zERMonTLY1NqMJd16p8HAvg/SlTa3M6XDfEIIB8GITgzf5rcB//PVnuGGjJl2
2/DU6xOgAc0ID24Pc8Wl7PsArt6ppWvnDwfsoNxEyCW37EXRSNLbZlvHhZOcjBd3
OhgK3zWiCXND1qw3dcDQRBE2jz6SyMp/baJzdqLEHqAgSR7t8/1RLKeaya4dkWga
`protect END_PROTECTED
