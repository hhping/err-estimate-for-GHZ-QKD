`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lu5Q9+G5obOYw+7TQ4zObtzoKmbOGKGhYXih7lB80AmeodzVQoaNkZVGDj8RJDxz
jFaUIQTmHIjEbOSXHr3crUxtm3jpPPbtQMqdVkMPQDjNZhsU+xa14Y6GrfDSRCoJ
a4nOWyLaU9B3eQk1RgfW0UzexJTbwROOmLDNzm2rKIYVMO03Tgf45tKo9IwI8svY
gP1nGVgfvwJfR+/ntnuYdQCY7El9XwJLuIq92henrjD/css7cb8Tq9o/hIDX+PNd
1dqS+OmGFAnjDLijuVE1OsxS5oM5O/VSyYhVAU39/ttd6vtinDKVNw9rKgTwZjK8
ZQtd9S/rtKZJETmmh0VmhSmI05B33bKwTyfGHA60u6iiuef/ZhbC4KOBI4uppZBz
xMvP7g2C1pUKtSaSA+Mh8dMG3OCsyyulz30jnU0RtzBhmfFUA2UA1TiT5leDr7K8
Cilk3s+3tHy1B5Tp0dwqvKfKkjj+c7nlGQ3jk8TERSyt1d4BA+/HDj+Y+j5K6iDr
ORQlkFFHMxrBOqNqgYtuodG16MEj30bcGMzZjcRS+T/FD+quRJIIY6c2Gy8hiv5n
+vMNYjf6E54qehyIn4oLVCSG+hrs5SGyc2v41tSeL2AsH6u5FHYmTMLz7lAsZL4D
+2MQ04uT4nipMTqC9nWezFxZ9Fj15glKiDy60OlyRS8Tj33PXqOlsby1pNZW/1KY
5KAB094hLsvZq6vNYoL66THQlUS11D8Ma8LohNSX/NJDpkpkE63Gk+uUEYF3r+nX
6JL3bsVgX/3Zzi09yZTGbegg8BCTbs8hqcOfLxwyvQy2uRzd3ImTApNKFfCeQTsS
FEkUrXmCgouLBsGDSTfZNje0SBHVmR3yceEwAJgoq2rlJf6qfEE35HnvjQR8aCsY
yGGXHxdNofWwHFZsYOhKCld0cC3zVIQki7Hn4cN8CZQC3KF4QS7+U2JC1xXe8AZU
5x8zxRYhEZ71PyjYC48c4TjIFlNMVIbk2hW9MOVC8ix3sj04co0pn5ZnHFKUTZuw
9e+rwXu5C3hbBpplCSYly+TXCydWF2rNDe5D3P3r3pqaHaS3SnaQTNPSAzzavbS+
a8//esDcAucIdtLHxgRqGFmVxR4F74I3GGniTa5z7jklGZAgB4SErIotG82vxaPM
0E8bMq2LvQq79KKNBlCJuioivWoWL6T7ITYlV2ilhiC+z2kPCeqCbdVa+HOdPtJQ
5SO8tr2azFoEJdjDkf7RO8JSezs88d63RC4dmatFxMfRwfpLGDbB8SOZPbrrIHv3
p2S7717QsRcYrNV9ekNoFA==
`protect END_PROTECTED
