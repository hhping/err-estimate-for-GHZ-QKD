`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rK2YORLbNfwAR2//cf9qVs3NJnDrtHBGddFYD6tZLTD30dVvn2dpwhqJ6S3pMf/
Iu3a5euUcysJXeeHvlK6Lu41cysRrzZlrzjM6z3CK29QSEyjpr2ExAlkaH8XB2UK
KDrrK2uOV4HpD5mnR79dEJSVNi1BgID4iZ6wOmDx4eWOGPcwM44FGlSGFKUipMzX
DHGHgA0RfoWLb6HsD0CcK7OSs++jWpuI6O+bxYLmil0kMLNFqYEU1rK4GdlzdwOA
Ai0XjTCtDsxBYf/qxHFnCO3Gvj9CdzOXjfWiNtKeMlBz3/vxc6srStnkwEXT3l8t
9xOSDRVla6wwg+DqSPS+DM2ZaSJUZvQrWAx75zKxOWBA9l/Rrf2sqJ+wYzM+OKhw
WuJCh+7/Ee1xm/azN3cVQLqdY6Xe6prodjxxa+23QNQ4y3b2WLWcONU2ipZl0I3k
mXDyFw1EU3LHLorY0lF9UaLqxGnPPdwl0g28FCsJ+HxaKc/X7/r56Ayrkn8uPXM0
OXi06O5NKvP0cOteqcBPlD9iryOVZVvGLcD+8jg1/PVDU0hCVGOhCIhHJAcbW50z
WjU3COUh4GoIA080zd3YMCsi7Qg9csCGB3bvzHAqTU+9XDaSe/yp2hCHwsxFCiCp
SeYAFtcUYFl2hti77J5pueWc+1m8A5iOhKUjvOqIlmsr5u5Rh0VJPG/q+MMmlZ5R
64iEMMUA05mDHr9xqp42UBvVkzFGN75eyQFYvPXhzQg71MP6K4p99KL2I5E2uoYx
7YDjs+WeXXqs7dZw219dSYlbsQCdHTGYjpvwHyEqPv/NeX5yrhRy6xamhTwg8/+1
Byxh82NQOwzpEp2gq0INC5Fjix/hVT+mrN5vgRNiYoGna+EmeCsVB47u8BOGyf/Q
dHdFa8AXnuey8aYY6vTpl9n2DlRPkIw0ZPqlMHSXkv0=
`protect END_PROTECTED
