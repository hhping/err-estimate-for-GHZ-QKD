`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5AWQ+pFhZ+ZoEPkP+59LoCl+/LPQndRgjKMZF762Nhqmlv9PrV1lWbs+DpknR1Y
U/ojsko8tN3g09moxXaNIMrhTxlqqNVLrLXGhb6lbfMGtqS4bSD+P+eqIVhqHlf8
xOzCRzT6+y1kHaLDBaLocWzRotRbkD5L2D7xfeQIwSJtsf1bIUjIY6c0wWzjYDmw
3MbBOh6a9gP64o2U+oc2OwIVg5rglLTnlgqOVrC0JbQMqtME7lyaS+Nobj2MWp2N
UgHofwjefZIwP+DiIUWnnfB4wrqc0Q6VuWw7s+YYdHbfvdXT69JsYoX9tFqaPffZ
sgVpwKOHC7SyKTOT7Zxs4ZUCOYOMk1c6w64UvYMEpy6suthDm3Sc0/j0T7Nte9E1
4bLUAI/QsRzUzFotUmYI07mXa/HyMRydimN1vQQReoStE1r5ncktGwUocXWtBvo6
odZxLYGnSrDeRmc1kUXwWyOjjY/4VkEgSmep1Cb4JYT33clESePPFa/6irXtBPuR
DQljcgjDJifwOMNQAJKC98kQTWgaJ849/8W6y9lP5miNt1pdXlDdT3lTcsad4i2N
U6LNhcMliNOtNQH1XyRVSaE2lc7wwUCsLlNBLdDW1cQ2dv1DlPQmajb9TxAKpc70
rCAFoUks/TzP17bE6esZx4uSS3AGnagGwFw795qDg0g3ovaD2vjDwHYJcI00ByPW
uO38wow8v9nGDAzG2iA6zy0d0FPgXCh+Tc7p20FQh/ZYJ69JFym3qla9QjabHpD3
ISDQGeTGySFmyPL4Qz7i97ZSRZxdxMeI2Pp28COtJPLDHczGZ3xifMdoKcR8vNP0
NZS80AgOU/7fmEHxxe6Kwb+b0SLFO+XYDytjMO0tV9hKJjUU3ZvOhqBAMXjNXlkZ
iv4M3125Ycv12v2IU+4XcrNC50Kmv0qX0ud32jU8PbRNJVyZX4TbYZJTpiYe+Bld
n10gB82rv7EwpbxjzpLMKOdNKedr0WebpYlkk08oa7sVYr5Kr5NHXFMAZGa75Fsg
2AL+fPUQ9ah9ZtRMh5UZDy+ZsNMLO85XuTmEEQLmHc4Niux3ngcG6XyoPS89jhWO
MhCOxk8sBUKn7cwU6ibTe9Ox4hkCvHY1MaMkpBHweRRkVTTP5S6sB8X3AsMNzNeG
o7xvpR6wEfKmClLie9vjQfBa7fGhKIFwifLALsdYPQcKBUhAgpXBuwMgVEnxTsnO
lTLnJhn5XkstdPaD2SqCewvmWR8qUoMrdhLkC1sOOwpRHuuG/W9gO8X5KMventnI
io6c3sp44CPuHiJTEOGQhat3kuIjq/W2U7vis2oZtH+iAQGsSOGfIg5z0Km6jgLi
NrHfLKPnM9lib4CfySGzUkXI1MdTDIBCRXcML2LZAYOlFRyVCcdeJtULx+9SxGW+
gsRMQ0XMkWD1FKKRSi1KQplMalIig7Vy0PmIba/whcVs+Mb1WcyonzwWnIDbL9sD
yWcd3fHmTFs6wDj9ydCQ3i/U2wq0GJ7nnXzKSLM5spiLkEEAKz0uNbvXH9NhAMpe
qQRVfueHdFG4f4FPe02LcW+G0kqjXM7NBcIcMOEsc1mpZUglcuxlrUU9wNK72py2
Gsz/6dCik95eC45qf8jEpVDeERKPCZuGRoqGvjIJ1WK6pzno9ERCE7K9AFx/+iW0
MVSzrp1pdBEfv+taL2YL/n8St1bzRit5nVSxDqwOTowPYrDODhuv6EXUA4X9sIIz
i4lN3XvAPRKImaiFSk/cJmqGTE3W/Tx8+zfcenh9DFPqVh6vqpH9sc09eFpniWZ3
BfFzVehNNpsn/zwQIJMluXspAqJEhqXJqbdoKj7QFne4K61OQdllfYZd6woJavRE
ybyXJBvNmZFEBhhfoQCVykGsXIjtjvSBRCbh8m2XhUEpHTBFsr2moUXBthjP8cMc
c5gV4BuNcU/X9ehB1GEvT9JHQ4nGI6+9KJ0YP+BKjoq0ctZmzfR+4rcvYe+2cQZu
VOTDfSyaBlkYsQtPlIuMoDdB28JEbuwQ6yLFtO6S9OYzMtv31GRLJ13Drj3/iIg8
jhiwrhsO/4Be/c6fXwnYl+W7ql4KC0v+fb32LD/MrPvi2RVMfoCIO+eScDtXGRwL
ckX2HFZZ8C2EMEcMinoz8LHXEoApqV9aL6zCUT64TkU5HaWW1AuVTbN9bDU2AuIw
r05aQP0nQN0GPSgFr76orvCEBfraNFEOpdkqP4G6KJnl3eofi84FhNsGO5hW9jQ1
N1XrdnNdlyJYkrw3ZWJ9QQXmgzV9HaKuDPB2tHTK0EjlN9D6j61S6tK3grZBFROd
llHXjLy8u4BcCC4/FyL8EEm+T+kWtVfUSVo8GMO3g/dXy8I1SHgVXiG1raBIW4mB
WnyTnwC8poKKxhhcS6sMNOSOQEdrigEyhWKbsxnx36H5VYqlWIdRqr6O/Nki55Z9
lT9Iuee/LeEdS0pV2QCg+KuqjUKdY4xfK6WGEVQtDiv1IRdFpmT6wPlCJL5C7BE5
WB3KTtZz8nyo2Iq2zvxMzxuWLp06AvCG3MhYdgrFf72pvLkcEBK2b4NsZR8fJdXJ
Vru6Y1TQBCXWsNP7a90lVT4XnLoh91wp9DgCxBOMMWrCrDDb8MamHDU3mOn6Zo3e
R5EG+SA0YaoWapQd3DeYcA9h/jKpJQsJJx/GbMRjLUe3CWi6tFwHKNahipWDeSDR
bd19BeI/Z+xLpo0hGtWAVPNetbQkKrPbVM0WkQbKjsUSSs1X67rZlojtR5DYx8Lz
jcTibcBHz6+4INQNVrSWsmLYWw+3oQutiX9HtFYmTrcuPst6Mo+J5z5bhEPMp/9T
aEcYnTPc4wi1us130VHopEVNf3cenxXJSdMlnTVQiEWVWfjITfhZ3k11MVZLWpOS
Noi7RzRc7yNO4YUmESsLxPjH3XCYQ9QNVUKHZvbARPLw6KiCDnhwQ8Xto6xbxak1
`protect END_PROTECTED
