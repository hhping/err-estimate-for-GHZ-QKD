`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9gC5QCdKO5XHe+w4dzxUuWR9Gmona3FJYIxqnejCY+p7fBMZSQmP+x1NTbwMOm3Q
osItQ6QPUFKs5JhhFjI7JeL8DC/RxDifZHwzKT2CmUyfyqUkb7U0WrWONDjiDsYw
INxpTUO6iPYBdtXAEuDJVb4O16a6NEOpAHsZQWVr+dAcQw6uLvghnfCf1yaRamdq
uJdEsWEtpzhAY+cJWxGLMSGB0P43hvpy0UwJSdMvdRgGEaJ+/8l6GscE0k5DzfVt
VvzmgYLF7ooyMviD0OktNTNhckmcA+9gPOYKIV0ZDOp+frvt1PDSKKgHAGwJAvyo
oC8q+RAwdZf+B4NEk42r2Pbzpuurl4IMmwJ5ilTzBdooiG7Kf303Z5W7uc+CKTaI
kjzpQBdWq8fp2AoLRQ+edkjRVWmAHh1TTyMOLlOZmw16otUfQ/MeiK8kyIozKELA
KmBZlAFUklCxqxBiIvgoYyRjC9mvejXFMQ+01H4Xzf2KY+RFL2rGkKyRJ5h4vmnj
VvVLzAxGbQm0u1yJtqabelhCMrpdn3iARrpvvjXeDij2KAZp3j5XRKExyTGBV+T0
WpoEwtxK+nPK/dTwHKCg7OA95iqZBY9qFE9jb4PlB047KfTfu8C039cR2pg+WeDf
S1hlZzJrERjsihoVqkOQ4R6NpgEw/QQSu1e6GoqJHfRFeP6MBJbgjX4L4q0y0q/I
DtfO03+w9brjgHRYXxh2TPZWuIH3vSrWpWYFtLqQhvWQKSU12Spax0Cd7m/pDg6I
QsiSHdPiu0PX1R3uXfaviFmZHPg4t9e/bvGgGgYMyLkqkyM70g5JalQrRbqZrBAr
ekDIyWap5ToIjBAA/Y2Sb2UvsmsqnjMkBAYPDfVJ4bmbMqMmIk1KB1U8yxwq6jao
P6ffj+Mrnwdi3eeRFXSJZM4M5gHAY4i8DaHKcECjzUkJGqzpmjRG3SLk6seDRDzK
swzNN+n5i3iYYTJ8GL6OxKnxtMe6NhN6RjOGT3IZIFzPW4+23WLQITeBwtJQzvXB
O3mrVIWV2h3JUgZvCk1QiRGMoeuF1vhHnvrZRkb0zePvCGjlR4S4jEtYEM0DEpBw
wfvYBuvoGtariXogaxaEWefirwXZ/XfoMuUwolmqDUvaKYc1CXVNizQMJ9H3qTjv
7TlTPHOnfUw+QdXu3JxuBLGQ0AVU5x4Yv1VST8muRe/CUhH/8HsbgDYz8U0mQWW2
zB/BdTICKe3hg0vu1NOYoPbSOOUCsRhK65UP//v2WRW6Or9DYJMt790z7YGPZ7jI
7opUD0rV/oDGPzpsV6TqT0BPqRRtp8UwjWiuA3Ocnw2geHTHr3YFxj2aRjRutreT
ueZOkLfeX/hnzRsjZOjm8EaMWdHsggYZSOgnA4m98dCrhGtgGXirHrKS7Gc6meis
Kzb6OeLAGlYVgQf4hou1kzOr+Kwty3DDqGomwAQjX88gf8nrYK8Xo9h4vlLPrVDj
NkRbyCGiZP6zxDkGjT5dBBr6zFVlxl+HaVg7SGzYJHOew43iXaZbwSlRi9pZRGSZ
T+eOXkTyrPaKeah5DeEVIMONdbV875kwC1Ekz39gDFXWwgN3FA6IqFzFP1s3TUxj
rLH6GF+xdIAMQYZZHPesoP8Z3lZAUROcbXq2yOGSTYJfss7X6TgrG0x5iePsaO/T
DlSN0yuPcSjtXRuy131P3LSoyU2PXuI0yDJORIuRkXZoXFmdmn+qPejkOlmO0UzT
iiN2zASCxDB5qqaCwgSM0ASHy/P1IHaRrF+CWMT4X6sjLOP3+M/Fe61p0m8LmxkR
EiFCrGfD6ooGuac3LU4UQtgwIP3tqRhgjYpeBn6gnwBkjpsOku7tb/PvN2VLeowz
IvkwEGWJ2RBzjh1F1XhsRbBWI3ilHpEUBOtZ87FCrxrYTPpHGXtwfe59eWxwInFQ
CP44mRUpbNDCD4j8qQG1FYuSo/N8WGsxCdPW1FaLUmr5Hui+FFCPjqkoiy6OInFU
Z5j16Fcf4PpVYL3QdFNbMGgpUYoWSLnxKOZR5lzx0VsOfbSkPYAayAGscIuMREiE
0hVJVDlptqTGMJjNPWXVoLAJwzVjL9jbwcG9FOiaUaQuqekVMw9SoFEhOxQsdLAn
gPtlDnelCKNFqQV/bjWzBcSygzYkKIiLbVzyAAfWRkyw2seM9xXFk2UX/itfSl7T
yxEu738SOPXcyuF9q6K69MQz7nmBA1W5bNP4b43GeUz+Gkbj/mmWCHGkV3UVT677
JjaBku/OVs+3qm0wmay+W+0XYiWDoFGC9nCbD2DW209jqrn8I6rRBNnRWO09WJNW
69J4ZCKtrCAWgNxA+q/nVvPJoyVK7NwTnwKah0IGO0ho5dsFfy7QMPxWd36ZgWC4
6jHmwFeKyznE0YY82FsbN+uaRh9w9k19MqWfEbQY2Gv8prpLsCvvqw7/aec8yrOJ
IK8P7xLlX1mnoFn69AjgjDKADg/Uk2NRhqDjheHySOAZEFiGJZPePThEXl3e6Gl/
BCMOclImEjEMdK1BzPZOQRhKeYZXMH+dgO6lUFd5I7MPJVeQpOjpz+41WPbBkvzH
f/E0WWURUWjfDEU4/Rk/NuvJptzJ+Pev3gj1Yel/TPulRGq4DpueNvshDxfDsmRy
GvWBF0RmnRRFnp+tSoUGQJL85/1LXbQoY338lANi+dESluoPgaObsHNOJfjkA+9W
UB3jE1ER/dxwpQCMk0boDmKZES6HyicxrL09KwmbGlV7MNWF9VUknMmIcSk59qwD
FSG0BDyHwlnUZOGIzu/B1dNVJtI8yhExvhLQ+yp2ib7CEqf9vQgtluFbe/Rrmu7o
BdPu4KNMjj+rL4CTvJGaw/ny6rjcPibP3yfCxN8W9hPEBI0sTEOj3flikAN+IOp9
vXq+09b6PKy2Gwei2h0ZUr1HUdZPLp0tCeNVF3JqYI+M2mhl0WH/iLbY0ks4mDdB
HyGwergohq3C6pgOU7erfHLZsxhyTDJT5GeQRWUe4IxFLD5jtGh2XhlNqKGZIiz8
uWt5JavoZ6EdSNqdAZRZcjVrxpX/hT6vQUK7gmBxjBZfa/4Dd3W73+GGb97HcuZC
Nvzuib9P4p4p2MaX42K6WgcAWc4YnzksHFplDWTrSKOjH+sroaXukitWK+4lF/is
`protect END_PROTECTED
