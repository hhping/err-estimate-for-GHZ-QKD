`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmqKcHo0HOxwuI3abDeJSb8in6iRhIIDmY4gUttvpf+oNQmGA1Q+dd6Cu9sudBdf
o0a0FVp1BVlkGs70SdXeNCg1MJHnZ7DdIsOzYT4sa8CA4OyzrX5JOZxdBATd+uoQ
fqq2Uy+vfZdZXbjbR5lZu3LshEtp8ERRBJIVwsZCROuE+je74zkAVI9LcOfVUK9z
SE9y+m0aLA2NRjcKSwwNZLSczAAAwzMwrKsbWOMX4c5yYhh9hYxxLfbtb4mfztcg
wYuMjAzACd3QX70z1hSqwsnGlP16B4bmh3BH+Lot9bzMeTQmr+IA1fJxQINXgpzG
5pXvPuYcSxZLJUfI3szO//6ra7Ch+RQy5DJrbtOJ4VWhO9EE974AyzlNsm6n4X6V
JysH98tqfb6btH0+QXbk5U/kSxolJPlBtonUEJ5BRm5cld+u7nEWS1iWDPUZ8Q4j
HFTl1BBAasIKnWgzM7DOBp47gQ62X+NyICmt/34Vs3RR43hJym9itBIi5zZXIS7v
rBw9Uk+Nq00YCN9EJrhWWgrq2U2tNkBJIOi9+krV7hDahdrEKTJkaKLouI2DwokR
Gl35E/NKMhpf5eu5R6IeSoxpUIyYP3wyKvTzgcKij5E3x0CksCRoI8WH8navMarQ
yWOf38y6074YA8qr9iGeaanLUHkZXcSPOFK1Ppcs9H09+REhxdvD/kyjDuAvZgTY
FNpUdsam+L3QHfJS/Il0Ew==
`protect END_PROTECTED
