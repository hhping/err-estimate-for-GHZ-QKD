`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhodz0qVBao/0ydEh8ner/ZGjwTW3+GDeyPnKnz4LKB9cwV6ybK97tNFhmQO9xJ2
NgygJbyheWaFUSleixhfeHK/gpOdBGjk9KdSh2RzFRQoo4fnd81FtDo0wAq70g+d
J4gFVKT6kX/RW3WbsnPlmXopA4Xj1nCrJFjBO7eE4IuG+FX2Nq9cHNK7rky59mqM
POlDf4KPs3Ca++9i0+mPdoZ8uDJe4pm377VlgaLD5+6ZJnzfejN5gp+x3QNHfvKg
2iX4i0fp1ZhxqWmgZZCWyxl0rECf31ZZf5MTUrF9iAL7BmMNW7BbB0TYKX7jr786
kWl+LdHl+lc2fB91oCsq93/AsaHotUfbYRXpDreqcfLPj8lPX9k7cFE1YgI2LPpS
vVLQCXB3RhicdD43tPa1HX2PONlE9jT465h7ekXtusIC7a5wAD0jywsfUAv4uAyu
rN8/EmLpGSZsjpqxV8IoKy539XIyz7YZKyU4jf+OJnMoyt3ZqZvdHQs2okkAyQaA
jC3wNoUMBk/Sn24/1YKPvSRc6NyJpRP7xLrnhRy6/cnAGnUosv/73P2OTq0+n3rJ
aajpP8bycIvJYMXnCv+gJz220kaRAS2Dbg4yNY83vA871QKp+XYZuEE28FZaIXgh
zoGzb5DKCWmMN26+18enyZBns04wtkbL7bGSv98D4UrqVeuuOh62WTqZXuA7I/r9
UDZy0kL0IjDxORBLydp6wd0+z7wpjU2YjyBAXpj2XqzbaFSU3nlu10ZvEFP8DMI8
IZb/KKBNPuhAOdCrb1p1XKc/kTa33IU3WmzeGPlosX68wgxKlKzdtUB9oT7dyD8f
2RdU1QZTFeZfvU6ytNhOW7r1TGpeZ3rWEtHAxQyYwcJzntsxvl4PWQPtTSAkDVvO
mU+LjH0vYI1VryzR+sNcvGJBjodEeiPUWvevX+LiWTssYRQyp8OHMN4tprBohUGy
4Us7xbJgdUa+NALDnLFickKRUwwV5hT2jp5eXwbMVFqwBHcr5ItdpBGUpBlsXA6H
4lsbj/tC3ZJ2d1Mg237T5yw2L6GaOklh+oB/X25BqGl72oucW6mzZTdb6UwGqChJ
LfNycnoLBra1+6Ks/tDUI0611IUYItQh5dYTjZTWk1ITxzRaTbz6HL6fzACGMS+S
XIjVFGTg62GOuHSinbzAwfufUBCGJz5fbVCRJzDmG4dAkXjYrOiEF4FF43v15zMJ
cjcQBlpKlZRxoOOlpzr7DCYilhMjN8XvAqR7r9VdaZgad7i0HFmIhYkdu6p/pU7v
wSU3mrjD1M7YZE+/K3fy8Drd0cyDlaHrSpAd4HS0L2IzYYGnRM7/6tPVpiBIJ6IZ
wR7FVQ97svl++ylnRyRsn3QE3I4Ni4YRrZSqOmOsEKrhTG3he+XIexir3oNdqPLi
Teh5et8uLsiWYqq9NU5gcJM/EJmgfGJbGgttrYFOFPkRBKUv3FlBInNvipGsge2T
/S3777oFpvTWdyq/qpRTcQ==
`protect END_PROTECTED
