`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5nSR8xCnEgO3koiTtmfGQ6wxy0xF8/vSzdRkVYogiPFIWERQB+YlWZL0jzRVVk6Z
hib3eaNQZW5y33uhkJSJdzyFp+TVthezWmvgYdOjq4CwxR1JFWV/zOOzrAqFOyQk
w8WHSYJ7nfoz+V50abQ0qc6PCq4r0DX1h8qRF7CO4ZaGY+FnqNxcW0rOs4e63Nf+
munCB5emr4gmPAFAmH0rX5v62teoQLZL4P3xtShH+5asRI+TIDiu0/CHLNCWvZI3
KIsshWD/H7GGb1oTl8VXF70Wp8MGAv34IdhIkkX6K+3BucxyFCGUKo63TWlF6Edz
2REy344nPKJFtchkRZ+bXOqSh+7OGJ/0zrlMOnpTncOw7CneOgH0OGWqS9VJk8NK
IHe5+7IThBopRHNQrthWqC3nevc7VS4kLzWPvl8lIlxYMjPY87p2X2sWjPRODV4M
Vw41IuVvILDvhppwHEArYtPQLlZoDo3kZkc+rH9ZYB/ydZweD0S12lRlhSclAhJM
kg77MNgcjm8cNdi4do25zZ2TviRAX563kvpIzbyzJc91qihIFXDGtO9ueeFAdeUI
3peXEzTQLaKkLoAogPBiJnm3tdeTr0ZOPkyDeBDWojocr1hvZcQSmY9qXMDKAYIV
ijgx82bw4tRxW6EJuHZUd++6MQDfKW7eSdaz35+DtfsZr6FTfsFmZK60+OsmosWH
BJ/445OM3Bww8m2niYSRL3w+D5gRTw1IbDYchs4DfxrH5VAdjUHh8Hnc2m7iT9EK
BlJLRbpKcz32G3lfHG8PQFlTaIXKN7qc1tLJD6w2Z+choJ0LTRQIT6rlKH3E2twW
BeMC802Z6ajR1JPxw8rOxa4JntYAFfAb4f/1tp71Zt/Y12JLYi1nm/hMLwO6oLVi
IEdNwFrF0+GpTJJCUJ7ITJMwyyUQ0EwWTNhJ3ZJ1yQwUhty+/guS7ZY44MUfJCuA
1q4Ds6IqB8dteCfFm2KPf4wI3wZaRsuK2MZfx2aujwylIMcgtFPWl1v0KymqR0Eh
gxSpYuK6MLV1FTgExh3z7hEkS/nL8Ggw7DCVwy93612DkhydpCUs3kfWGKlXLhpt
cgpKqz7Tciyx54yHmOg8vbLcCM56ZqRJmJMAj9eFrzGq+4Aa1GzsVO9XYoqLo8Ol
iGjVOm/b98IbtOE0hEbzjyPilOkwUBldPzzcd+E/xiN8xRqIErPwHMLamBH1RqnM
PSi7YwVbkAt5fvoTfc1HMir7UWM++KPQidSHRRCUHK8U/L01NGu1rYV7kheUoT43
kVpHVYb1O09DEdCuonNJ1nU8/+vb1ZnH6P05qMsPZX1iwL4nCrcC3D07TElryE2m
KlBf5V/ujG3OPWPDMUDTcON9bm4gCR2xVbcwZ90WBAlplr84wEfztVKLAo+1WppO
QZ/A9Jrz6k76S6Z0DzXpV8smyEgojiH84QyGxBmpSdqfXYJXIzspyplbEc6dzl/2
xSAnpNjxAUjTdD1xjSWOvjtNc1hgjy6kpwo85i1d0t5qKiLzVMt/Y2Awplib5mP6
lKty1RPsjH0hap60m7a1JX8/fluANPZiyY1mx0JRo4Ji0EAxGj9kgxI2Ntb4bQfJ
REFI6t3kMMXfoyZVULIhqTa76Vn8psZFzHCyjD5b2EP9us7T2vO0XCO5yRZy6WU1
kLMLY5kveK8EwbYCEoMzVVLuGuR367DM5iGW02vL4dZuN4rz3krPpVPwIx5uI9X2
m/ijmzjo/LduMumgUZ3QppNOC9mrIxkyV8xAMxopF9vCLe6to7Bj/lJBKIJ4xEOh
S7ZqcNtSKsl4JjKOnw/NBGkOwRyUtV0cTGZc589upjw0xm1PtC0AvJU+OAPdTshY
sNQnoaxPOOqcklFV++gOdhVYsxLEbkoB45tcz2iNbbuD5ixeVhPocpfM8H2szbtF
Aur5LHDG1k5g02OF+SxkmMtgOwIQlECKSgSVfXDf0vJu5LvIOHITslNyLdpbZ1yp
YH4JiC4rNLbeQMSnjH4ODCi8/14sMkUMBN4kg1r4TZBD6HnRbIh5QGyx9RU34gsV
RyljdsjshEJ0u0cdYxI2t/0MQvvvj2ue3wxAUG69wQAlPp5k+jpqDfzgnvEjG9WD
JXX+1pYToHK3UQWSn7iPS/Ob3d4Sc3CFowFWwQW2Zcm3IiBhTidcHN09Oxa4ig7r
z7EzWrJ8zb4g9ev4CGxLjzowV9XCy2IxtCq+CQ/5r01eOivYWRd9C3LhBoH4QVPG
BROFDbN0mPuc0TiMrQ4d8/zQanDl6FKXZtoluEI/ZfURuApHbOOZ5j4KujiiyFRc
PVOWa3XhwmhlbQwqZLr8ipBxAsSD8wvTJxnrKyDFkvDZKTpkwJPbEN/Pnl0I+SIv
wBYWJ12AdBGdW/lAIfVAxsAkhry0EemqZ1pjVZr78LmuQXBRW/HeoFfC3fjVG5FE
bdKUMjJMQ3YmIVpAnBdM5Hvi9z3jeXkCJAo5GV8D+XTRuiVCbaiNfogUZvKegGzK
/DxyC6eJpqdhWqqJqLw8Fsb56wTdHRmiavrbZMDAKgiy+kUmuzRtIcaa3eeZ867r
LI0IqHRf2ycHAhBIXcre7KDiahYWkt/OtjJJqMJ9etr7Z4qQQ0Z1RHuImIjcDRIm
eHPDMSsiE3tVQxAHwj7EFolCzT2q0rcHTa5S7eDg9qNe+KGN+ExR+7i9SDztaH/I
EYxM8L9YZuu4auFwa8oiAVWWcj27RTy3Ih0w+bnKJhSJ19Vl8Z5EVXq9hg57BbTc
sqI1FIXngT5AzFL1iKh8iXhuG6zQUA4copxoCmFDstYpjUuuokRy5AdHA1e65Dug
MroAZBTuW1ak2HlgZH45v7CkZKTo6i5OH2CaeXk+EzkzyjQUybWygdmxtg+AqOSE
EOb7STB9B2oQpMh+uZp5+GN1lka4hd0E+rPYfByxKznAWctIS0kLdHHfFUbZGNyC
NrHCoMU8fOQ6rFuvJCnvFCniIyot3YGXy16jVtF578HT9oVdPuyfyJzuJ+mohRPR
Vo1UcSvZ7c0sf8NHUIYN8D0NQumuS964sELRD52MrPY+h/SHDrMtqYszFWn9Ye2H
BFzoAfmMuQT79/om4RqGZuhqax5NXQJknH7oK7oLj4y25R7HB1BaeZ3bijIrnNuA
l62P7wiH18y/1BBFWJ5Cahg4BWosneXjM3IT8ZU0Eb/bvPwGQoLW7RDhBzvc/upY
gNzrQ3oIc6jXcpLIzACpGUK/wh+b4YrLBGTiIQCPk0xivIcm/FnXxm8elmqHv1RY
ISLNvFAp46/h/vO8e8qbaYfu/gudGvkSnhfHXl1/PznBbDdwJ0m+gS9ljQeEvWf1
XxOt7PX6WoCtPx9DgDf+TomV/sDuCYD3IqfAgfVww+4sglvgPSGHu8DUn23l8FPt
519jCQL/dRVvZPBlj8h79IqoYN3yJin7DXDH0EXk5tDhITQvWYzjsbj11U+0YSH7
Fros18pQaxFD65aQTzfM3Nhj8xItA+drMtkCVPpCvAyTTaHqnrCuLHW26KdCFHSM
Qe70O558fBoeQg47338Ztm+a5QGWH0Iz7ihmjIPJKqkOe6yYcPMJ9PmTVs8Y5Eh+
0/G/LMeDTcT/DTA3L+Z/GC7cBXBcdVnUtL/J5mEF4PysfM9Q4Jp+/hvUl+a5zZ5K
aZbSDFAvjS/x7yFmg4hhXVLLNcX2508vXeK832FrTq7QWIqhIqgo9vZ6w6Zczg+P
o33B+ODkkXgYpCxPzPvlgaIpF2ui2n5bYVGSUB4eqBI4Aq3zmadRtCoDXB3DDpRw
Goszc9v81IY6TteH0Nrjn3CFCo3hjPP1IcCiGc8mkf3557a7Z87NYL4gfg4trcaI
gTd3H7XM3u/6VB/HX/p0pC3pp9fhs4y0wXNuvL3Bv4zQtXOmek2OeffBtqdLwaQK
i4J49wh3vIIiLIlOzYgi3czLlptF8lHUy29dFi5CoEkiVgLDf8QeyrbO4SXqrEJz
C55PglnflbbmkWu1O6j6ijFZ9dSqrOSsxGLGOIQigLoyeg5ajwAqi2o3zikJ4Qy6
51OCmG4WI2yKIjWrbKvkSPnU4KNHgcKkIrPwzR9IBjwvShXqqSuXR7dEDia52VeT
pPBAVgwHJVUzusLWzHEtTDnSaG6P8GnhIrccl929lXqCvFph5vJY1VG41gQDFWOq
ZyK/LescXgbZozNc41c4tC0lSEaHNhdJCZLpzboGTv16xG6Z0zjbrFs0z4zavmid
drg6JHwQb40n2BRLFZ4rxvEUnCGsecbfzVMxjgmAE4PTTCkLoM1+DJpHgjL8vYkh
m461NJnKQpplekuU/eCahUvjUK4WcP4djbS1RGsm6YJvooRIHDzpxdXySmy/9IiE
GrB4qYNb9237+x69ojtTeUQKr9aivcTwve8aXMSqDYA0wmcOx3pBL5uelkfZWb0v
qDqs4T0RyVtOH3pFmlY2Yh/ZqrYGYoGBMM90R6VBN8ZmIcLM9ZUOMs4yy3sYLVEv
VPJyjEoD6qUg6331xoo5OBSTqAzdxJ1GvG80PQEYMzsRvYYfH9GuNs1T5aJg3unH
0XAJ6yjl+t7fC3NJuddBhLCtlBlmE72KPAp66lcIViaYc/IvOfkiYFl6KJlRFcBD
hfJ7fbUrbnH7E5YPmjpj5rxMUi+qgvuyfTTHE9Ogxuu4tTAVIueVLnMHdqMmcY6H
OofVEiHpEJ1EeR3dnuy+d4zftXTPv6IB5tLhX/vid1wN7da8DvK9R/2gl2QtNI/r
vWSlodczPnxVgGXF7J8QSUYOffAjKYdhMG+4AIAdnXmaLuxCRDecWkzOegZxhzFV
pPdmq0s2TA2wC6tu9l5RdFL1lrY5hMQLFkdXpyYvXm24EHGTG3zJXSM4NIw5UriS
p74lBovn07Q93LhF/7cucpOPKbZLsvEmJaH4hY7mN+a3h9zIYfMmeqeACC/O5Xfb
dFhLqgMGd8qqFmmOeMCiw7lMLzAjTQHXrT03VOZP3m0tInqHYau4kuiFtIyesMpV
ZSLD6WNh7LVMsV2VqElEv9CcbRnLmM3RPGv2Q0tbYCLJiWi3kZgkxohtFFpX7M47
E1XN8btj107fXIo6zPTbRC2i48Vi3kzSMCmTPF5HwmrzwIeOAUjAoNzpBqv5s4+n
xgV0U2Qv1P89LnUrXXiDbY3SObXJgpsYwrANElN5FLfkBC1iKICEBAyoDKUsWOF2
4w5jTuDQTINcLlP2lf/H/ZyHtWb6eZNMTgw/ul+cVaHkNlJoWcbWgJuonHYhw+uQ
60pRu8rMWdfyfK4pV7tKVgasHIlu21GZlX65OPR016y21jKdYRwTxhPKIGIJIdyY
E3VJHZ15k34SZwi8gENB2x2jJod1RB5FIQsM2Y+Cs80EQC6YhmuGgK6glp8ieKj4
AsZm3tMBaDmYXrnaupc6ZPRwyCbuKy3gU3Lz+QLI/PA09IUYAFH/kQ1GTjv5/IzD
hA/9wheLdkAVSbM9yNX6zjvheeEzB2mLHBw2L4902FJEqHMxeyG0s3oJJ7dgTvFS
xZkM2RSj8QGKEvgTo25ITPMkr+ffqaLqcDHcSTZ4GAO/yjNmC62GdZ+PtUYM7W9u
SxRi5dKon6AbE4rYFSOggDtir7ulH8kCTxsLIITnFDX9wyXS5W4QIwzNVbLCqAoi
kDlYKsO7QwS/e7RAnL1th2fjbzdr+EezewEDMFZrNutpe4IA7tXGF4d8mRLuVBPX
2Ga3f6nVYiwSkzGdoUQRVA6LSqFXgb3TDTGQCQYGqNc=
`protect END_PROTECTED
