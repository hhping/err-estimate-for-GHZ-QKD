`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RESqzz3qCl5YE0ZIBupgRsKM6WniUPMYIu6939vFE7s2D+3t8iCC58eb96dg5dNn
ZF5pT+/yZt/NFGjyT4DX/n1zYfyJqBa4L8xDtHrK8WhINLkyztKcC6nmbIlqQQ/2
C0Vv+YNBRBI+xlD0Em8WmMBCanxehoLEdgFX/ac835zhP/dc+/3+u3rx3w0kcKfU
Pnvwxj5rqZi3+RjtPgrQ67K0y+RdwIf1FqL0GhXGfMmY7xKZxPAuoYwe+rKew8tO
iZ+7iftvC1ue5Q+4vEzL4kEwwIFzu/6Rg60B+UkKesRBwer24iik7r08wkf6tmsU
BuOqm347TxFAE7DC0jtqdXiKgxasm5jfTUWLs6kn5hA+xfJ29Zqc1U+YEj9Lpto0
AKcpOjRODo1ZWOIc5M+4295itUCGnO7mhiJChkrt+Gj1vwW78F5C3txxDnOenbDH
o39ngEHBLTb40ZlofopXtg305Va5+c83MpShvYfUU5gLB6YoixilFmNuaTa9V1We
5sqB+zfwdNSgKchzyV7we127AsAoJa8oTbhLrlQ6UINo/Ggte/Mh+wwagts9lyAh
4cDQFA1HM0lyqQsNM7BM5apm8DakjbQQPSaW+oMJR/er+VfGMGj5d7zTU3bJwEYm
GiWbrmlCWJJ5bbGkhg2bGVglz8pu28cPCzf1X+TAQHHMkdgL56tFHNMVNV6cn1DK
uZbH0ZgAJrzGCrDqVcJPXHadNrmReoXunz8wRB7C6sqEapmsuG1fdNvfUBIxagl+
k4r4xxoZx30IeBQ8kEF+uvb0zBrVN+6wyBHH1gm9THQ8jmbciCwL3m9VnzZ24I2Q
8A8cBgbJqVOvEc6YnThy9mEELtlL2mCxpnRPRiwHMAt17e5AQvfm6qzF+DCT4is+
YkugA3KA7o3OpY43eyul/gPaODc+uZLaN4CGqVEx5T+CtTpWad3KEBcJIJaOo2TF
5jbK19+a0yoQZ10XHCzWnSpM3ScyYB7KlXX56YM7cB+MJKmVapgylVaUxvqP9xO3
Oh+hqfDXxEAQ0Xs5VpT3I/FQ+RxSirNbWtkv699kurhZUi8xzEpMyXBFQ+yEtPcp
vz9KtCBJ5U38l5IIhW5BCt6n7gj8meNjpP2EG0k9Nel6l8vyDr6vxmpbyQe4IPi5
mqj41xZXAKvu21dBCNc2CcNOpHEW7G3ZIc3HjHfX/JMcU11u4Vl36gHEtcbryZ2R
WzvFiMYf7r8LD8vIv9HJo0eqg2lV/kcQiESyWbEOBfjiUjVUqEDq+ENgibvrOstG
vaKuShqauwEonSrtqjpzdvKNo61ff1MZZUAhx1WbOtVBzDsU7j1M8Vaew/bkwFqh
GPdQzLUnXO48jHQBSDJaUMlNSIpIB5jzWSyReEpiEBxYA2z+tqlD6XtVzHV9GhPL
0sZYgQrHT7nTAEkyRFcI27qda6O+HFkEtn5H2UUoFcXwHOUKyu1EpcNWIaHy/oQl
`protect END_PROTECTED
