`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IIgi3l6AI9ksgUgiMluC5YfTSJWA2/5Xp46URY1P8/QzMMVePnV8tavcsOTdZeYM
ZVPMsHOks/zgNxNoN0wgjzz/acuE3Jtfv9JqLwhBM3TjqFImCgcr3wqk66Ku/y9O
gZPPXEFqYZHLi5C4B7ae1+hTNsTs9sRnL6DMJm4WwxlAoncRC7NpMGhgvRX3OFAp
CQKmK6eMdfLHaPgrXTdg45pELiP7Sw1oRGtFAuSZwz1kkQrX3Rud6eqrYs4g1alG
eA5+vRq9HmhAy1UWGjFKZ++oUOt7bLCisvnKUm5relTcoiYxumZAoBBhGy59DWZA
U0zpl/AuUy/+iUgcwhnuEdqxsFmRkmnkL/vMtjRYT6yv3Fw9BAQ/ICCtnW3VPfuS
3soXwq9AV7LQvwzZ0RBdAu80Q31ePva5z4FS81iHqdUotqybRpKil0y6Phv00aNY
ZokETS4Njm4W5FCYnS3SYosHlzJWPreCVFIjhW1qZ4LEYejif2HTDzYdmcKWShuT
6X2K8WWgRn6D2wiiszI4wH+1Vjayjs6/oF9xibRqVz38ZxB2Vx9CV5PPTdc/QgDu
7J8PYkBY4tjgnvkpOJFZ/jnkOz0HIiIOxWk7R2iBaAp33GxQXFD8X8Ckd5cgdYp7
WaNkiNcMKglcIOuMt2vy4xad3ZISxT0Md6dxsD1nCjum4bPJ1B5c7+QUfn8r50zp
dpcPUQpM2wuZUXL5kSIKmeS/3Pgd49m6SKx4NFmXabU8NFE/jkwPyP1OftZ/VkmN
KZO+aV4Gbq4SBdGW425xUTcgwJQyFw8OdJ3YfPSAqnMwLqsjcgPYDy+MWt/2q2iS
E85jYXR128nIQGUSOnixAM4jXCgRkAc2ovCp4CatRyji1S9i0MqMgYZ2+Jh3OZX5
gXixdLIivlO22/v8wwTPCw7SZsK99Wsm3AIETVb1WVW4qZRnnxP7vLqCwr7Wf35c
3I8lJdbyq1RgCYmNtGGHWY03lBWPnUUCZEu+Px+sX8+FQIVDmihWqU+PVoPRjO1P
tXITdgVRdL8SHqKmqQPi0vU93TeJGRLpwT7bHerO2DErSb7zntrdqemxpBhBkRym
tRaPFK+Rl/WQqsUVNgXxq2N6lJf7TpbEmfBDzle6qJVIs51H3TSQ23AyiHSA29U5
KLluq/gJMXbv3cflV+9/YnvzW3qqXM5xR2Jug8nlTq4S5XiHRtuzJjSJmeBGu4JJ
dpD2N2EybG5PcUEiZuzhBxE6hhbHlqgrkT2sj7VuZ1PmdvWsj48c+3iqjhd2WRby
2+bLIUgaI9nqfaStyHebMqEv0JGe74wH01/kENOkshMzr4cRonRUOYwkRqVxUFKv
nKn4nGEunrDnx16hVFHjQyKaYNxK6khKJKujdRwHzasENR7Uyr79QEC8qFfndGmj
vAAazpXI0/CBzM50H9viORgx32VhgCXkJmsjhH8zTSV7asveWIqoO1nARA74n+yQ
aQm6cHqcEiQ5CXAojrHIHZXTe3nMU1ORxf6lhHFP5Xdv3O247VQ6gB32QBHT8wN0
1x5eurguwDSBw3aoIkk7m1FRGhrAQg8aXKMSgKnTe4qJkSrQs+1Ymgw9Fy1k9UCC
hS2WyxOT3kON6wdeii+H/sETIhbbgeejZYHbK9qKDIZMy0CtWfv+C+/IDjoETT6t
BJ0+1aUN24FgSxYChmiL4pTQ2ORho/UKHd4NUqOWZGERlb72b3LnMbUWewtBXhkA
oYKZeGQ5JStSpqH14mXnoHKGyCxojf91E9pLHvoh+1JJRl51YZU5e4Y1NOPiQebG
ar0XS/m2EY8qbPNKCAYdt6c5SKoQJVFNO1SDmvskqC27Avlcjn3E7HatUpJivkVW
jwvmnyv6skfIAbhSHn7bPpNFobK3Nf9NrzJja4lqMhJsNO2M5tyUrGtMGxGM484a
qd5JbYIQgg7gNaWBegCP3nzHRssoCKc5FISpnDhhC+LGXE5zu1NkmBQ3UjsxyC3q
CbQB1DqIt9uMiRWLlpkx4Iy0eYHAS2IYl3YrRmKje9y8tE1nTzkJXUizDey5QVZ5
ENKpXa5koxj90lsUkbL5Mj1FxPWp2v0itjT0HZ2dDyk9b0PVOIV5P7GBWLIx4tGU
DNwbbdNNzUkRzecKnUm6e9tcdcZMKHCNc41C9Pi8NBNw4h3HU1NZYZxbrvGoXvsb
HZhjLJEUfehh9eJ0vjwZlRWOuq8EI95b09OV8Kx5SYKo5RSFrKysiNAgovpv5vrv
DsBslCfEYLj1Cz7LdN0mL0PGREwzZBK0iO0SScwBLH/wrBeU6NLdsc8U2MgcxStf
AYJfajc8EzU2aGBohMylNHp4Y/XOWtQGy6MtM1rtjED7rp/+MGJUHbMKBlZFNrVz
QF8c7bBHFt/cWsW+odDI88krKQoqLDNqCEqYln/SHuShtO4kgFXD9YqHb00uat8w
TEjIguVMQVf1dm/p8YRLrcSQANXoxYVaFGzgr6ZEhA4DqotE2oSzvuEbAYiDj8Zr
gCjOKUDu6CGWmZgVt1tYV6sMx9q0OwRNwrc9i69kmvA=
`protect END_PROTECTED
