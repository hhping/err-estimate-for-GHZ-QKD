`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MowqKR17oApq9TK9L+dEIPt6p6r4Hk3zYmn0mulP4DbRX1frN5ogZzGDXFkRHNbo
bxibIY9omRKYFNgJX+aQr6CEhIg3OhszN1oOvxvd4QR472XIh7IhrFEZYy/1ODtP
zzIXDFvh5DzHjTq8MDlxK/Re2r4F/LZpFGndaEHyFAER6hD9AzY6ZZ8AK0EoqmmI
F22PBkG9JZi26khzrjh42P02SC6fUqdmCuqb4hQIeSSbwBpJL7x8L5wkNgt1aa8z
SXx4F64BpXgUQuIQq5ltsSvv8RPhSX+F88KIWH7AK6Al7UM3ww9FCZ834kjiqOTe
HbpnZ3tNs2JVxJ1P32Ku5rYk5BqezhTTbWxvoublSQRiwo/KzccOsGlgeb8ZG3jm
THFIBOeHvIOvXuee1aRhtweBMiSUyH2EjssUKU1iT4c4t+IlLC93ob6pR1Bmr+pZ
3tzjD0+kXxNGS8vCsDvh4r5WF2/TIA9kE/TPG/rZ1IodC+GIB4VwSkaw+WUSxtY5
rSayAyqBNSb1z1c5L0XQdM/N5U3qEgsWgdng1umFmSTkS/1e3duplDtLilT25C3K
38qdptnfV8HIQmntxbABmAy8K0TWcxwHu+2pOztr8FMYzItToEMLKPtUUGZHeccM
x98Wgt1pcuv7oEGWYxt3rjYEl7qQ7gioTS8n+RKGlLP7IcgGbu4oN7E+TboVnwXD
3AJUTxYm0aSSfWuhLhSa5TtyHLn8uAnmLlbapUl3uVwP2+yNgXpiQZWsaiEEOert
43ODxVtL1rVAmst/HnJaBKOR0agZ7gYOlVa0xjW8irBDN4Dv0NZ7dAY8Y+e8COKh
NKOd7QcIALBBz6BfyJAvH6+vWRc+QCaPdOIRyuuwApkxYVIZV+u7Leo62qV3srcm
eoB91E+F+gtmEBDztYdMdZL83E2PepUsN1Oh8b4FxKI8SlfOXeZB3BO82XFpniaZ
GLFTcKD+qmsvqdAahD6ndoPrrU/whfSBxNIcPcTi/pb3xpl23A4tTM+j0krO/cPz
EMXS+idYBF99/p5gxYbjIqKcS9yUza7TM9YFXawyWLX+/FLw9xwD9uLPZUBGnI2W
oQvURaBEVJ/aPyPbS6f+cQHpAQPuVbiOia5AJ46AEXIDfF+WffO+liD0K9/GD2/7
4ah3p4P/mjlGRqxj6pLiXD0Q8rQUT/LAxcAO+M+XV4xlS3xyLsdmRXfGK/QIINvU
UevFiBYu0xTqtInW9XcFAyx4kJSHjec2P8fwJuir174Cv8rZyZVntZpeK50jUkWL
QwsZ3a4V1sVzbcOMFLS+1/QQ6oyzbwy5NlYJK1OtvUzmx3r/l5BdUfEk/IJXI+m4
S8655hlLctxDXeLs3h5QP1pDGc3Fr1KLUZsMBx44YDxUGYmleq0sFgNHMpVEfPFD
Vr2oZAZFBRfC9FfHx1gIE0gyKHPG6Td0T5uHrjYjhum571tGTW9kveNHHi3OjbOS
eDl4hY8w8sZgkbflj30xu0p36p/B+AA0Y2q8NLj0OTnvcyPlTK1gVkewH+zlI7co
MSRqj0nNagiJS0ELiZQhe5aC4aIE+AjNyWBnv6MWa2m/b8ITzg4bwuE96sygPq8m
yMMWyOahGjU6LBSO1hXif+qg+yX4bbL10LVblFU4X7mcYs1lM9p4BMJMDUzu8skH
8vkZK0DUcAF1bMCv07HPTVZR+0m5uDkGGTwAiOJiaiFbpW55zz4aHrpCtBMIMyum
AgcwQw76Ad7tfPQqv899Jxcl5Gbsm3xBPeCXMwYh9BcRZ+HFu/Tb2lKOd/Ym4hxL
VsMZzo6qaFIvU6/zqZcrQIGUnYrpZ+kBEbNQGKKamfJ90/KBTA3otQrU99b97tOt
ckV4t8ghMNpqzBxETv2oKmi02lZjiBXtdl73haGinDMdN3FUjlqWNyNw6sJZ/hMQ
MPzzb8G4WI1cpEohlW7KVVhlNwr9UNUnobblWzUaJgj9+3ixb8KTJhUjVIqBUx2d
t2zBwGruHNn9p/8vECQQTDTw3mnL7gTwDjNg/UPv6ydp6vmONLsuoeAuhmjNtpMB
ln7ADzq1LFYOXoWMP7ofzq4ws2TCk61S4tPseeRFQ5O54y23ga1qZQ5z5jHcdmB5
0/WysOalQxzmrEDCo60G0cOF4zCH7VLxt9SHVyTXCgNwlS2L8VSgNm/b0s+Y4tl5
ATilvtcMuePXOHcnPHtSnzO4bJ7KVPSZ0cqLAf4ys2p2y6hejSOvR/TdVb0nwdaI
XOJcMymrtztCrXCIFIrXYBTB/NsDXtH9NqKnvgiWBGmi/h+aZ+kgH9vO0l5J3/+T
M8rEncvlnq3jaPKAcD8HM/w1NRcUKLTzIbrHjxLEMfxVlIxNVCbQNmKbdVdkVfjH
f1MayBL9f0lw8apTbjtwMx0HB1BXxks7R4grFIFA4MC8nMRs2fMkLq3I/qBwYlcm
3eFQDtTFM3/F6WOcUTVcZgCgXc1zWVKBxwj+36BR1U7QB1/Gi8HLoBtDordgIP5C
m0A73pZFeydE7wYKk9rZADoZz9ZbFUUKgom5lm1Xc74BgjkeTpMGvyx7NNVodTlB
EU/Sp1kr+NqIIz3eOXqYBQOCItYfJ5FwdRZrNCQmVgIDzUCtVcj7Ts095PbT1oxq
ZElQEOdBLmHor5UKMgzjReMS5BZY1zRTsYFMn1TqyZQbYNPMua5ZGOLP9bc/x1EI
MEy8cVZIjYrsAzSvc63a2dD8LCMc2V7R0gedrnRpvt/LHKBckaJzvmoTqPUH0/aa
8s13MQisMkElOSt9ovUwUXzDAugrcAo/E0gd2GYtXdSN9T9/bjJREH4OYzvR/yUi
X2ezYGx7kOKiMasSX1McaqLWl1nlxkixQwXYHDJtVf8b39qb+9a5epGFHCxqeXea
gwjW/0/lN9+2LAVjbS6fbZbkb9whN0v3bIZXYhPniUCx//+lhVNcAt/HcwBG3IMQ
r+8dY3xv/v7vc7wg6Rsca/3UP7CoEJptpzbmcLPu7P5CRHp3/gEaQYS/54tQdYE5
Kto9p9/0WQ3sxWdYX/nH/huNxd9NWleERedpAEmGzCWFqzq4xLgpK1xuhoor8uD8
GGctdKl58dHfo6Gh3XECL+iDvmmbqEYG5m2aAVYY6ThFlzv0ngkxdewsIVPfQlDf
NbaJBXvNBjgplulf4E6UkF44wcyhDLG9E4IXYTqibnMkmOSaB1dwDlNl9jpR5JHi
FpuPEzYXJN1LGOh17kkKE34T9gDgf5req28hK63AuJhYMrZtJ53GNkvL8i10WFNq
GANaXY5yHuzKVfAmmO4FHFTLUxbR6yRkGVG9/7vFdbgi8PpAjXhZle4nw+40Aw6N
caPtJEJgl4kPKfhF0diz8KkGZfdFARo+O9xYv5aTSTIOJ+n4OKonBqVaWMXp2WOF
zIvocEyq1yhoAUBYRI0jw1F9TQiVEoya6HIV43kqXFy216uBv37krc5dLOnCv30O
Dff3Cw3dlcx+NUvxfNUq4CXfPQYDAT34/TktD8CHUtgpK6rTHAwCkLhJYxZChx3x
DXzEdVRPmE0rqvcO/o1OgSLpE2z7Vytm5kNdNwbEEzEgViXm8rRgAyDXxQMUcMzG
pJwmyJY8FPxpSRwn4WDmKt6bVRCNa4KyQHPehIEKQyCDC5RYPd4bX8JLyuhfHD1q
8y04EDD9hKXiGhyRYbgBeeCxWuGWajyJxH4sE/jHYzwhJQyPKLSXInDOMGbxvqKy
uIbRwmPt+gaZuoyT48VRvb/z6liqddR9sN9Bt48vuLrAq7nFoaHMx36YDXXcVjsH
VQuzxOh6eBhh2qGOpb5AK6smYk8ryzfcON7l7NRWo9WdMh5vkwKj0oQ3mtBX3ACY
HjumPa3P8hDvA2h9ikEE9XJzmUmIRFyDxHcF+HbxCQH+CeX5E9lsL+O0KW4tqf94
x3iuFiwCEYasqm12M9/jp/vjgnfZ8Pv6K/7WJgF7MoUeM1GGBv6lRw+bpJoK7536
kpNVFV+8YMBQgIG5or2R3IujfZSlDiS4VnPZfa8toCapyv4CCdsxXXbiEkautoJ1
xwABKa5p3vQTO7sS+OtgjslFMCaDIwoz21TtysS27XpK1puKHkJIEo/CiOvGYkdD
2CmuM9xm7cYlZ2B9qHFQas2uGf4j+gv77FsieNj2+h7MQ8GAmb0c5PHmfsubm6my
0weakOYm8+CYn5Y7bQvNQrvDbhfnn6/TSTGI06fPjABsOv7L8BOz0tUJT17v6b/f
EE38QkbNmLVJHqmtpvBpCOnfcRTNy+1Wp9qcBu3EOuiRdOJMXr2WMJAtKOp5hy/D
HJLgY7vgqM/u+3fEmdCFxJk4Ue8S4fzM5epV+Z61CdCYVktn6weLK2Rc4S/jbNc1
Oe2Vw9uKKwJYt1GHha5YOWoS7ZaX7T2JhJgXel4hMXH72TcaExjmaefFl5hb7AW0
3sHT/vXJOoGklnVUEV1hylqwGRGYVebPvI1xLMlBL/EnO3lmBvQSFQBRvHDZ0x7w
k4VrlKGtM6kj+EGby5jjOT3XgsiLV8Cu34rm/zMRCOvB4D0t0rUheyiaBLX5PwuF
3r/IcJXEyrNoZ2uGWicBdjs5qbkZVeFjXX0kI4/L1+5yJfzXWtJAq53PCWoPUnhA
SHQeu6ZzZcd5Xfo/tDfqs6Z4Dnfk3TlrnlJ+8Oxwc+enqC/Hb/yvQnL5zeofudZg
KvPi8u31MFFwtyUvkim+XdfNt/aq9V8k5Wvogg6xVUrFtltWxLgi0kyncCWiPAtj
88c8VQSGqYvWT4B2mcrItdMxtPEAGqEWDKHVoVhNxRlNco6zh0yvgmS+zi3D9FyL
ti5BPldNOFcaBg1grhZmGQgUQr4Rebm26VVkS9NoYiEZ+wHGGAiEOR52hth2Xz5j
Mxbc25XRWVrZQGaBqH9iNXZZWnNKF0FOYrAo86HdgmdFrlbUceCfBpuvo3skuCEW
uwZFP8m9Jj6vLzh7qSB/mmk3C16fSM/Sj/6o/ST2dLR22PNT3EiHZ7mdDtluhVIM
NFb2dvVs4sHFFB7v/ak2j4GArUYJQp9Sd4XXUt8rWlGmOPEC5XntqvRuHE0tCBPN
ayjTsjqtXXflFhCI5ecx67FXhwzaoYA2rOphznQPbSTYJzvfX7+2C+DhQOblUe3e
NauiHx/xFRC2gkaTRFt+ErPWCrt3asEVOaoY4fofeI6ttOkKZTyDVy52OzJN2zRw
orPoIMJHF1g3I/sO/36kPEYAfHGlHSjljBUsU4UtSzqv/k5yhJOUhdngBUvtysHG
0mrYgv7ZjVkFsuIJTfMEqnaFA1PuwbnZCM9iG+CSEiqRjNYmQuOnTSvUlWocZF5g
N/K3V3Ts8HtA6m+102XB2NmOD1ptfUPBfwXdm0bpTahorMaSHmSqdw8daP7QTnSg
jTmM3hzjU3pueSBCKD17LVwQOwabGA4DUIz2ZiY1o8kiHpHFTmDAxywm1Rz27PiL
YGLZJH7x4UFZ6gVpDb4q2alEjGsYod2Y4UqQ8JN+DjUbS0QgEXeW8ffMDrNokTST
+H4qXmGaM+UZY5QJRFL0R/ZKwIMJt5ewDoBxCE7dM4eiGg0pSJiONKRMdyTN8558
5Q6kYqzNlyFob7iANF0DpqRFxp6/1uXaNwA4SFQKRJPcUUJ8QmOjgf9L5F7pfLMN
oTLr+FDdkJtWBjFxiJmERyUdxPsPJ7xe1OmylkDdoLqTA4Z/prmF6vxK2EQtw/Z1
pHdXEF6AU9o1nrBfRY1uTFvoiTprR+sFPHfAGI641OYZun8geDbs9JE3OBqE/TpZ
x9PUhe3fksILqLk5U/3TUMErR3tTdW7FycgD6w3QSqIFPj97ItLghycTFm4f1kP8
URkiFd/gj+KLHahS2LvQGVjPHZEpHWxPtzLaaefiDNiZgW1vdhyXZABqxKpfOuiw
8LUQTNUq0RD1jq2Rsqvj7GdvMEWfmI3Daa9M14L8CVmyTZw3sJg0IgUBoW61A25R
edt6S8ZrP8V259h9X30oO4XPiPK2eRxZ7f1x0NMZtsS7v33Zmsrd58lDy3PtGnL9
C69Xrnw4YdtX/yERm+21o6m+y91AtumIavGAn1PTBJukd3pwUloVLZb2oSPeOV94
TEY2kAH3ZUOUrUIfnYtLPag9xoLWBGwXSiux9tGBNPdFnQc48X92IkC9WSPu2sgy
NZ1PK5aSep0Xm50rlBaqHFnT1S1kbF9L4XT5g1qUhqZAnyBCaiRmGfii6tnpU4kP
0kagpSsZFrSvMru9FeZS/ihlDOcp6SJvE4AAiHGWpV8904rZpcU1T4VRUkhpO1TP
ddMK88A/faYH/0CKf271eFFV+LWqLh79Uj/8weQngYnDM0iP0uMUrD8EhE9PhODY
sqKoaHeBrdJGeMYCw+lh9vFT3Amv6+9eP1QmYaMMb4Edec5j6Izm5VinbCnQowFT
tReEow7bBtGBxQBRhQXk7mD3A3NRIBlYloerHA0+kU+avPXMuBZz9wXA/V1J8RE8
/bLh7Jifu1upfIFKI2CsJgfWOGVFCP0/HkFkrFrCi2sMe3jB7F0c6ngBH4z6fUIz
kLImcVIbas5+Hl5bABYe7jZKUxNTI1vvsc4yyzRUd/f8oQUx5q47YSjAIYqmkBMu
1+HeaXnXzQCFYMkDAm8BpYQh2UMKJ+RkVr7UdBJ7csjEdAvpIYqekuZk+SxSHrT+
vlHLWxVYm1m8up0aKVUqQckWiXwwmIDrFGE7wZiGyXR/TiSuUoHcR+Z5i9yXOU+D
TOhI6VUXLF4cyCehMqpcRxAsRdwp2SJCmb8NvO3hcc3zH65Yj1n8YJcZsP33ly6g
meIV9GXczMhf+tGnjolZS86EEUm2GGykSycB1mUbYN2MF6xslzQe05bvKvaeOD6k
gCAp8EFOfDYKig49Bky7fhznrsUrHM5xNy4UeyBf0qTqq0JYpnRd0jIAfVLUeQLO
n3v5sBv9KxM4IxcNs/cX40bssnYmXSZooG4S7qOZYH9KKJR1jLgZQaFhKIdS+pDx
BTCrnCtp3aeycyThSJncl8nHySpqHsOAr6WHltV7Izs57eeAcrfU/7Ba5TnaKm4Z
1EGbAGxCOo0RrnJjviaZdbEd0Y0IjwHTV1Td93xS+8pQfGrNVi7ZSo4z6MiUkR2+
YhwqEQy3aN5POsJWICtSiahqtiIwsvU9VqsBUUPPlipKNr9uuIOYlngZ39zMf58K
EfErMD8B/BQ2e0NkrvlkHwECPXNGLynMRwCZK02b1b7dAVjloONJJ2ZjtCDbPNjJ
0cJOe1OPrAsMkjYDMHHxZZemQKNAoHj/5N3/AIJXawAcnuPBbvr+sCkYF4Idnqne
OBs4hG8WZBR+aINkU5T5nsXx/xC31JJqvMJPUZtIfEz082H3nZwz57ahjQNFzDUr
uTQHWqiix0nPorrTt3ZC1OZujc5+ek9hEsX+l+pXzuuO2rYKni/3p4GQEiPMHrlu
ji/X+hsLGPVj/OA2EkFJBQM8+vPlssdrYmtaA+0Fuvz+Cww07198ts2CnE5tI/e3
24Eq50vVkL6g6G3Q2A4iTM6Kh6jkvg+4b1O6P6mtBJubUTI6d7XDWmdk7sFlnkWA
rLKvGOaPeLT9bb/xZnMSs8T8hjyc+MOfHgJsXzLE/N518qNVbgdB8QGjXwORrYI0
HLCIXTwmcALPDk5vdqRu1qqmy05Wrabe7eLfnR78y/oP18TKntWd3gtoYiywTL/u
zPj+u7dsYGKFu+p58h2KJ4+luv6yMp+/AwR79PWmDEzjuCmG15HYZ9WEe9h3fwlb
2QYB+v7OnlG7Jex8VgKMN3OFLMTGjFbCqgaBmjKRe6BvxGFf3gzeekjerlzYMg+K
VbwC9wnv8CAST837ekdtdXuPoLHuopMrlRea0q3Q0AE7nHYMVqtPmpydRCJUtD+t
fnoHhBbUGqNEFpMl6r6EyuyKQF4ZLvweFtgcj03uX6liBnEjr9FiUSLMKupgRpvr
wYTuXRI5yX8Y7pZz/GKtFh+LX3Ck2I2YlvtbTXpFzHBv+kY6EhR5TyWVfRtODIhs
OQDjcWDEDfLwUsrZSwsZxZHVFW2Lx0VsaZJ1+F4QvLS39CD70W+RScwsLB8WKvha
AzmdtPkDaOHic1UhrNMaxJkvh6S8MJR8KTKqi2eaCtWwDbA6UdfsRXf1zh3D/w+V
4ro8P981ALHdwukQacsgHeTkEngDWvqTLDKGONDSms0khMmrefumxlXOSnbsEizv
7QQZlOMlGnbZ4ySQKMlqXhTdt5eN/crojCgFoSzGzcN2HvwMXj7KbObaItNNyDwO
+AKTxN4KEgVTpCpAQUCsVb3e56uhr6kTuzf9/AC/mmMUW2g5/uH0XKPkEWwHN2ax
tDDZQc3ByHaTj20LDeuibyQT581AXA/XWgAQfZyjQZBAoEcOA6mjT6Y4LdcEDUCA
S2c6E8Fv0+XYM9DwNNtmbdVjUpEL80k0hojTmY3nYarvtT2QOqwp3aXkU16IeS0/
sDx4rZR6nM+svZ6xhnMsSIeOjYDDFGlJTUrSMwsF4x+dV3qWauJm8zchdgqOuSkK
lbp+ZGOzdYtMJRSY52MJOU325JY8RWPdbbVDTG1CR/gzaAYJwTq3PopPsfhZOKM4
pG0rXVSQ8pk9qReXuJxrOX1ui6V74/c/sxPjNzhJvb9wJop8JBlglMTgUQSg4pUX
5QVoid67xtnHI16yK5oKCa+xrA7zS1Hh7lOZzYzb9CLh71cDVm4WavQn5sxlHwBl
1apnrlVAB1D96Fm0oM6RnBI6N8n/U0b9ghrYDtLeGmZkU8jJuEt3qHclrh8BPKdG
E0zIWPi+nbTMEXhJCqL4Ga2ORM5nDvtli4M717WtYhe8WGU/G8CSSPs2V8MQk2a9
fsldYwboTQ8AykF07ZVD3aTWSYkYg/bmgyLyRnfgnwu9q8SprQ3aCUS6W10fRVht
lJYY1dno7w1qVGkjiw3Arceb1k/KmzMDamstxJdoyrCKoE/CAHnAeJNg4ZJhuzAg
AWnknxbe/2D82j6RXtm+05kloGl7YKBDDZuacaU6E9meZLfaLNWVK/zXncZmDnIT
H4yNJDHGkK8FjazU7yvEd4pghYoi7LwrBhtgPdtk8+GZaAF8/HK18PigN4gqaqEU
vpA9LmmXyNeKG059jN2SGRwl2CLSr+5ZomSLDaQYq5CX190mlx8XGBy8xl06gSl/
JlI3FVX1vzd+v5tOEoFY6cFrpD5/secfTxx3QWJZvCNVAQQPo5vMYuE5JfieUns4
slTVDKzmLUWG7I7vscmtYzlXQOqZtC/f4ayjcmKEHMkjgYXzDiNMsUKBRmzCW3iV
eVEJpFHaow2UCxRZBFNPaq1huudGrWeLmldAWmF02ZhOmNszFK8vfZxQzlgysHWx
7r4BWGHTZ7YMRmxUymTTyyG9LUmSRLDqRTe+D53C+nsS4vekvUx6uc67uAYBb0uY
BSpfGZIAPwFoRD24xJTjRyzeTfbo2VItRgELNBa5epaXzFL8bF++lVi1v6nGGVh2
TfK2XY7SkA2GE46o22FTX+aEJYMoDcmGiC/20L01bbUrMXAGj+LVMXok8ej47QPT
BNJGlMBe0k3pGPX3fLIcUJfvvzsZyZDHLYpNtywlFg8NVb9WNA1KKcVdxb7OWf3b
rIE3+5HuhXcjAbTINkZkoIzgiZW8KyZLGorX4HRl6GcXj8hoF3mhcngZekhuvI6F
ZJnMCmYoj2Fw61n3CZzEZE9+qAcjuYbMFRlos0MtlfYU/zkiw3mECIu6dNdP5dgZ
Z8I+x/5OdZB+kj4Xj1ERoFt3ntXaTcYQHUg1uVcwTt3IxdVe2lsl8orOB3SXD0T0
/FVBXd7XEnyLKUjDV4KvC40Lo5CO+kb8nx5FVU/rwJzaBnKKEhBd+3wVCogAQ5NN
TPlrwgkZkA4YbKrhwcrptvV7k27D3gUu/36nmlMdnrFtpF4G3h5/DJNBwOpSfjRz
S/TackfMiGEnA2R7D+0QNx209+2NWODMbnk/YmXR6yFizxLmKs8sfu+2YVEX4aZx
QHpyQwMUjLmni8RYYkX0bIIRL2/LOWiubd5P2rrEP/lrA82z7j1fU/PWtnuDrBna
hTdqBTn5YGB/pJ+aDAO6IGUJpk43CrYEQzuYZvWNnkwte5j9F6Iwya91+5xx0hY4
eoah7CaHgNGfZVu0YTH33f6fJDob5lZhAN2II/wnL6uzjcYs7kL6c0wAaeZuojKl
l1+eH68B8mZWbJQ+rBvDB5mRY2FQ1PWHyj3C/F+jWyC9Dsj3zDz/zIl5M9x8GU8r
X3Z/jJWjMa9Myw9938/YCFZ6tQzIy0TCZYt5FjRaC+jSdDMZob26WHhvpU+SELHX
fkL83pF6Tgztb4cWoWMvfzFiiTaZ6LQPEaNPkASU4xAefTQqheR5sO924hu8Qcyl
b+NHL2KJEf3Ds3syuF+CCRmghYEYY8aMi0beYHKWJzjOjtYuQ4McYHlm+lmvgD/3
6yM5cuqLl9P3KMmK4Uf1X4m+IIQK6GhWCgGExKoSIVUsiuPR4KXEPmPS4RLz1xFU
IXIziWwcZMXf1wdcn9Mxffr1oeXGjr91sBtmfNvq1SRRw9VvH2kHz2onHlaHSnww
GS/8KtHzg4Qny9rN6P5oZRGuEe2LHwMqToTIrKRsDLbz8BFTlSx/xfXD7/SFl1om
pLZZ98rsU9lkibCTrzJLge6iABV0u6gUhgCssZ/fWEKEzWZxN56ZKf2E+mE8VrTY
zafqDh9Hze8tHpytobNv+cGAXRwhYXQY+4JRjoUIWXt3jQPBAj+7awp6X9phk7Tr
1Hl7bK6YnBzm1Shgrd37Qj/YdQ55Jk+praSGYttegxOUo0Ghb6F1QBYCXBhpLMlK
972LUwYgzf8+yuAkRfax1FUdCUewDmNIGomSYhEfqM7Qv2OlCRkSNKHnRPWXBibU
JaoKVIOeFc3CLhxh8OsJZ0RfvnPU0yZwgD+4k0bnF9SQe6eP0b+gcDyhaCFPZKk4
GiKjV5W6ccAhgnINxBoSS1cYBaFghSuPGMefjSLwX12sLS3C2wbVG8Rp9tV0Vyqj
t5g7I6BzZbIHWW2RoDhbfijeygCUe0/9OwgpEnvTeYB62+7lQOG2fZh9sBg9P/RN
wleZeIHMe0bnjTAxbcUoFdQu91uq3Ic2iFQsRAJI3jpUyNdB7JoUoUqt5URRC8cn
dcsoumyf6wF5xfcDmBH/aX10JBVBN6EwFUXCkBnPWoCXzMv2EkbkvNmeJZj1JB+K
74u2ZDJQik4cQRhxy7m+samydT0Qo208jwY/SnwqamwhvLqG1K8JhAd1TVDn9lrp
GylMeYuziuioUvxSsdV+UyyuU4N7tRYtVwyjahR/U8JN35IBwqXRNnn9OmnwKW8L
ezwvzZPoOBIjn3VAhNSlAe/n+9dskxgmDLGkesqrfIHPlQ4eOQVbmYCYOwj6hxHB
g5gJwKgKYqQxTBTNdZBhe1h93QdUxcMvaHHebRyuD8v25QDeHB4br/VVu6oC+yCw
pvSI7ZxK7cIMJQC1urVYqTsvzvo07Mj13WSCmVpKj18bkMKsvUVIeb/F7oI7d0h1
7Eqo3wS2QwmC9kP03PE5/IR1hWwgop657My+pc+0+6YZzRjfPcRhHLlRkzPHv+oi
vI3JyEebaTO6Cv3JqNtniz3qAluF3Hl4LK5gp4zdq9U08R54Jm3ANwF27dxcbxTb
DYFDUgLSDBO+Jr20mbDW1bnCAO+oiFSCbbQ90drhClX1TWxoXpJTfAeZHxe3bPIY
LYdOuofpBgAhEGpOldGoO1bezSQNpQAI3c9IZkr/9mIWLamSkJdONTe7BapWThlM
x9Y2bmyr/YcRncA3kwIm14Uwy4AGKPMVJjzVG5eT5hSF63upHYaWzzV27KfIldls
ryp0RL3AD8xymzwFEAAnK3QV2rmyPw/g4cYQgt1RELEgeuc8FA8QNjauMdRPqu2m
cey3rvmCaQac5mzRo5SX6kfYrMAz0UY3c+WTFQnE3wC7A5Z2+kevPIExslkpeYKA
jtCW6s24qwRYgijPczAsyh/2XhsNRcFgXwDLhi35VcDh/ESNpyl9maksnl5e+69J
YotfLCkbnoCRqzOs3mDhdtmP3zkYI5a68WLvdDUoFTe/znhAid9sn7fJtFcjNtks
yWsEBALSaZntMAtnhBqtH6GUpQosQHzmJRd2frP288vIeaoEWk3kVFnTa3jbR63x
yJk3w1aBZSUOgDhu+PxnMkAp5XJtk1+p7xd88jdcVH71r67Ad7Y6McsQZKnE1qfn
Xm30Rauf4mcFpGLBlvz7J7IjI++tY63I/nMxFxfeeBdFPm72kHzqFVWEsCbn0XC3
Tdpld0Fluyfbmi51epL+B4s0Zpg8+CqVF7V6K2h+IZo+Jm82BEnbosymj/eQ1JK4
zg87/uuGGDbfHJdsmpoJ3OR2yx8blqfoBBQCuGE9vQ2/73qpzLMvQfgPxdYWNbFK
aozO4OAv8MktYgwVQq1SC68Y9IqRmSv4jnstAFJRPGkCAUj09LkQbCnz4Z9Vq4qh
gz4HKEEMx4xvJablyMJLtt9F3/fIeYvThIhr54s1Vb3oPwHzmrGDWHTTmwzzErSL
60gesI92Po/dfp1gS/aE50EQ3ix7dEt+3UMtRKH+5lPhhrkc05ZM8Ff6Zn72WAlh
9NI+HT9mgoja27lqmZE0UKTFpcpbuBQ0xgZ/sl1ID+R05NHPqh5xRI3udDFzRhkW
ExKvPJ5wLPdTPE8HeHqeMkAjAAcIN+eG5OtFvnYmKunzvaXri+rzqjoRc2k0lFbN
ebFwPpolaEEitulMVD46RS2rGayfTEE4JK6mCVppdv4ynRH/sDMA8KxfZSowUMRi
PlIJMHI4YaaRxIvzuIgCr/h6aNrGmYJ4nxpPcE8K0HlGaLYEzz6Ib9tKxcaQIHs5
AWIMUBlsCmveTAJGRD+XuTaaXSd1JxtJ3RRooOsBJZl5knh9ZFBecrZYnb1pxdoB
k7dqeAElTqMRcBGUfJ7MspEkLF/Npw0/9XdzLoLw3QL76/Rsj8+5EBLpUTpz3NjN
GF0KU8UH/r27SGWUkoKkw2/yU/pZKjuGe+h9CJDfgZozl3VjfASvqNemQCTLgFla
l9XD//zXLKSKf44NzcmNM1PUK2mVumR2UxV6y8Ig9/j7ZRzyhQcVSIMtv2CW4/+Q
TbksbvurJXOpakGqnriNuHE7+7uePdR6jgJAWh7ZAUda6WeGhaDayV/TooqGHkUh
5ZrsG8EUyVFMyuuCWRXJUEp9wfsGZaKmNOn0wzFfK6pRi/Slc5+I9ZONXq/avhA7
jAPBxe+p/KmRlHGt8SBfbMECBgTplJCJXeBVCE6hFUu7OcmNyGyrL8kQUzJpob4D
y+qanuNqjDxVB08gPFpftr3A6Zg9EALffH1uupH8oK5ZJL0iHXL5BsKTAn7BoZ08
G29dI1MyRaH3ZtbhKmYsH4K6+7Ag9fUwDQCwClE8G6gQpfH5OoZjzEWxhMbk6ybg
/FkSdOuwQmzywLXz2R6XyaBuuRt9OZS1QH0DBGifT7xlOQ6yBWGcvHE17HLpnqeU
euFxZjEavjoCj0t4YM0YIWQYJCKWt+aE4XkBNfvsZIuaD3WVUJpg8apqSJND0A0q
MVZfqdcDbVgWIJ10o6oYzWYVBsj/swvGUCLnvAJtiBUx5Ah0teKbvPzIgrqQNuUH
IjGh5EMPR07AVlVIljR2QmhQtJP3czkiQyiod9V3f+Z6KzTi9tod5BOTGZDOF6Iu
J1ertOQ6YnNlKDuoUUe3czuVRlti3vyqIvGLANSsbvcxjDBoRXgbUSjscBHBjNSX
Sp4BJVt+axQHj8VDSvrcHg4nIi2KVC2Do3UWA5Rsh8PUzLasUiqCwCxeisNN4VsK
OIMxGNw3BXqsoTo9OS94exg3JerP4VtYBiDmx1dUULUsti99TPrNuwRULOVWW1SC
4IynsUVi0LjMjpXJ1DEeUm0/WuOyyR9mPJuUqBQZbpFNF2LW9EM7kP/rDfBqKhvw
mUNkcBb2uB9UcMR5ciPZfFuAQK6IGk2udzzWeDX+Yzx7wtDLwKXihdI4rOM/TZoQ
HnDaIMqPhZt2tVhIOOOL83nN9wFp08IDoMmk85kE5qeX0e+R0MXnQEBPUg1vfXLB
CfYBXG3YuBiRo36ha3CBPo5GqMfjxdk1jFdlxtmy/ifWHbc6aZetFNkXVPaHGIMZ
pcUHuv70SwkyySACxFwIp68G35we9bqXLDk1L+SLRPm1fRlCw5tjLRSfME32OySE
NXJLyHyOIE+Hq5pPPiOMIPKgL0A8M47/6ESE2L34WNgL47E4CZPr9pl328YC1oh7
b9dxc6R3WaxSJoiS3ABiJc5tTnoVnZ+b4hUqWB6wVqBqljdBaW8sgA+rhxN/o9+F
rvfMmQCJDjqM/MsIIYkHaTBE7Aj/avIIiFf29BlSYkKYF9TCh2MlR6PyYoZtF14l
zufiJuAMiLiNg3xeBy+eUpgvbn/H81Tx1rbsUpd6wKlgEuaidoaU1fam+DjbJzap
EI3NpG6uW4VKnQAtbshdIdkm0W1uUHBDGtwUYDI1dMK89md9BfLnGMg1q0lszXzt
4YRqnmCRcKCsQbeJSk0VaImsBCvvh3qp6c+CdhPoxeVsynUkdkhtwzQUXNqmP9hH
w3sbo4w8WKJ+GuyLsU+x3ZWgKlUfzHV860ROaojCDCOQUJ9QsrllgaN0BXJbFP2N
2fTXFEsWkUVnn4dL3uXu3X3EOIKf25FESW0UwVkIgu+U/f+z9I2r61kVk3CTrNx+
whmtH/7Hg8nJ4/cm6UTNNY0KGcLplvfc7UywXnwMaf3JhoHuF1Eg3pppUeaZUV11
bJ43UO9+zeCo5Gm1rqRwBAw1rTnbdxHUFAO+bBgG6N4bHs1A+IQrNEx9OHhcWTiE
Z89cXtD1SK1F0QeGIWPNtpnBecz3lcURKHfsKXINiIpmpWHUivrEI0UxOvqEAcq5
xrGAYubrTr3OfPJOBCWJpogI8ck7T0KLMtilI/wOtqtTSdgqq+ak2PDftwk/WbdX
0dAf6Y885Rt805oEnEtjsvftxk7pF1phu06xtgejLqvqHRHHBFQZCVKU7RQLObS+
7sFehJe8cm/NoMxjxI9A5n0VrvUs90xnsJLknyjIYDwLzyBjzLY93H3aKnSMrd8Q
8qJ2g8r6fx3e7tvT14tmauYSQYxb4NP46XrEN27RSTVEQohRWpLykNGAzCfT2zz7
qaifOK3HXAgRj+UF93726p1vnXSj1tKjIuZjIhEvh8ymvjgg5X7qn48/Yx+wqe2H
Aseo5efBC+b/loU6Z63/Ca08kgJ/v17Tq4W1ceIjEUpFZ5S/EULARc9ORwtGe/U7
fBFvdKXOwn3q4C8IVRCfoR6nXMHCYyTOYwJJhhQYYN74IDiqusjxk+j0d3ZbO+Cc
0UQXjQQ2r+05qZtL3Jjsp1It70yPiTvCERnLK4Cyak7CoWmOiapM5sQIuSO9ThSm
WKci1REkfgvfkigV2d1NIeG1PB4ZiGaIn3UXNwRBFgnl5eOw0OYPek/roGdNGDON
Ye//TaRgf1KtJ9u3BzXQ48K3n3gyUzvSrwMJ419qhAjerFTJSYsa/tazbkv53MXW
W0kYz0VV0/eb/vB0jKRvEYDDZ8K8fzgAGabHIasGjJvMERxUMq0p55a9LWOEzc9M
0A4zsxps1+0iXGzsgvdUDyF+Uj4Fn8VY6zJK4LgyuG5aRne/zfAeQOg52ThQ24np
ocdqYZPKyx35UpP1/pzIEYtcG2k00/edpBfukRFjH4mmWbeFuRb1Uxi4D2hyUExb
aPIynAt1/S57aoZUpHVcRyiEUPojS/hlyfiUoxQLBq9otTC/Q9ffRHXOzWq+lQVU
Ho5J51df6kH52/2VXtZpQeeNv1tl/rfExGL1KT2cV7r3k6SGrz4GFd9s3K4EiPdY
osoHuiszB7elT2sA7jfIGU46yg4tsTpCfYLF1a14vDI5VOLGcU9EdEvqwBThUyuZ
8Jaml3GWwjeU+1yYVwZLxbI7XTvpxbVCjM2PPyANJXNi6QT/YBpANlCwjddcUFWg
FgtHmBNK/+xLyaDB9rvO/qWSZkq3RYkAv/H7ot0TeD0zQfXWuuih42QBmbbMQrFx
4YP/y5+0vUOBgFEmebizg91HPs1RvxyF8p6lF+q2NETtGT9/VEVOLwa+noxIeZJV
Y6e+QnWVh6zEoom6fy12MY2offCIbvvx4yE0hcGQGwh49M77B77uZ8Fpvbhdlm/9
AAdqCr5PV/fcL9+j8Nbqc/gJvZeeJosIwVQqD7li78PHl/8kZEZwzSAb2XsXE4u9
1/YZX51sniHzL5xJWYZykLimcGaJwQ11/QWXgz6eBQ+Pg7E5jJZz1QeO0Vzt+5mF
aQEINN7mXwq7ymCG3qgi9T8v9ilFI7lDobrU8/ZyUwfcBfg4C6wk77Eb+cS7HWfJ
lmctiKrZ0pNzwso6fzfNzWQJxRDu6ua8moobg1CSUa/lP4g1d+8P4x3dI3cTziNA
GLL84eLrjp6btql1DC+vEEbd2ZfaSwgC4YOc+GRY8xZ9QDrYYjv+CyY+6sNz1/hp
hhLiLxTN5XYFHPeV2XO6HXyCD8CvWsHUm3jbQ/7BKSOoEmpv+IyWP0DHjcbyKtoM
FqqkjNyRx/c4Pwpue4REogzdUoerg6as2U0R3L+BIj8JJFHTAm9Z+4GOAVQDoQ+I
HJoBA2vrnYXfZQ/EAGz2WH4gs7LShg3TL2ZIaTyWXuGz4LpJSVGi9pStYVg94MZS
51389LpFce2JjQS20Cxqnw1x3gdy8twE+8QPGeSq1/ZwHC7x6viyFcq3Kumd5JDM
7t4rRF2Nx4vV3EgabNMUOf0eeUCTLd0U1HXZ2tFdn5O7ZjOTptV8/mJlQlZIGxiA
ELBrjD0Ue++M3O1nH5gP5qsbXzvrtTAEUua24WDCaiEaFvorw+i23jIIPyD7lF+a
fg+bpXYbxY2MJAInAWWjiyKx1igQtIaZv2rD1aElU98jmEuMUbqvyuwItlf2ohfP
Ad+xo9qvglqpydyAjsVYwaDhRGc6zfwJNZaICH7dqzorOhZBMCHeF3FWRf2iC4FF
9cQjYlYKtlnoA7WvYoXYm3XGH7TW2C18/aM55za3eSi1dqIUOnPvw0rR1FCgslKT
6494s36gHhuv65TrQzuowug5Dxg/TbLSMAKqSavGKS+cRzctdm+qx9aj1PbRZpPe
R/hYTYYBnBV9Py4b2IXOtB4B4Uf0N5297bULoFnUQaOTcgY4sI4kIa7l2ypV8vor
j5i6wY39MV9UvchwlcOXHY3Czl3LeTQxcR27ci9utfIMA+o3O9qWR1E8p3D5GP+z
4zxZmscU6otkEDryOgwbEArjmYsxyVr/XE9AagP/DVUvVxRHVjAnuZxfOx0mW5uu
7KVwZI7Vrv13mA4+d6EwzOSET7rG41qNn3QS+wytWqQzlCWJkFd6kt5iVwP02LrE
J41Oe9kKqwyZlgjeo3RJBoDdC2PmOFQSGwTJh8DX6p9GVpMPxgqFZDRnE7pusaWt
KgSDWHYzXK8+ckkmqMW+ErJroVap+IKlL3dACxqYrB+CL9ACy6qYvPg16v7/jNbJ
KOkOAyp9jFGWQygIkurYorhHbX+e+3bra2oBNDknvt7LDyjDAC6/FBlkAcrkhzXr
3o9GNigq34lCF8Suy/REKX6gCPfD6DbOdmfj17EvKljHDqy89oLM9kTlCbk3lEX1
j0X5OJyb/NVlurO5lkuItQSeL8TtNylP0cm7ZojE7jq3t+isn/SPbtoxU7xaIZqr
d7g3ObR4/hKyFQYX4it6KxzKIWNml/tW8s8U239Vlu84GYpzZB+1yeCgndGys4Bd
0y0PGRpsOBqvbc0DhysiepHKRLHS2zB/hFNxuSgQAe89/JyPyZPdF5XmM+SnhSGb
bm1whLE3NKROG+6M80mst0i7fDA5laVFJVSuMwPHSsbH10r1uXyteRdC3m/jteTd
hnDasU0iHj39K/p953D7Lfi5gimBl+0VSJcDts2xFDx53M22zKQCUrLoBJHR01K4
6aAW9KwEIgLMTU7GEe5k5fDw121qpm6bDguigN6nb4W4HJscoMj0CfnidhavQOPG
lLcitl96MLTELamyufi8crD7axCvJd3Y/gVdOvjKzsfsfGrDwCoMWjngGWwuMk/x
Yk+nGw9h6lpfHO+KHAz7zwljA+SrbfUy/VCpdrE3vokQk6ALHiGHxP6cVRh8dBC9
5XUpn9jk2LAUW9a5a1KYaPA2LDtjW2ZJCkUYUI9mBawJmRuV0wYF2OBrEQGRerg4
mwbXkYUCMa/6ZBc3KKQQdP2JMwrMAoE00HKOjUP39Oy6HOC17nv8MR06UO8XFQJp
qBVu2RyAFp2/cAtNgJdMF0i4NnKxpfiBtFhwUMtOminVesu0qPTtVe23KCC/Ttpx
fYwWw+Jj+voFbWLDDHG38fYlRFEBhPVdaBHH74J8u/23x8BdV2I+XJHAk1gSMjNR
6ddr/MixKsztwF3DexBI6FqKPNstpXpMEooNjSJ+YEgE+7AUaYOUxTD45EaZ+BH4
8jlgmOlqW1A1A5V807ARj+Am2jXpSnXMB0Mn6LPgkarSOybUtGIooYHMkjgekqxy
ZN0C3W+S9+8NN7WOka7hCdCt0C36pm8q21GcRrY2W1aQ3IKTowRHY2XaTdOy+EHe
VI6S2SejThHXP6cITWnjEcyQrzjDPbMRHSh8bZqyTxn1YZHccowdsHOgCpulg99u
hfkamMBjJCwZbzK9tOQHKwsJ8NIK2mfyjAeg+hxLk/VeBRNnhBZoVNvpUGTdXV2F
kf2YFnhpwmjLM1dBDTLz+S+VjJ/j8oEdrVgLjHwGKjmhgUwuOcvMHCWQkdOIT/ik
Yh7UeHZAG7FxKZqyJzSaBUiW87nzbHUyIqofzuI8OAgflR93GLpnjBjKVyBuGXS9
hVE5/a4fP+BZ7aQsV2JOd5N4xMkaSGP0yWTAt/58+KxwhCQAdjrAphiXBSZMuWqR
agYn1BaOfdRVQiXjdHlZkap65XcQYFzBoj1W1bSIkpcPlMXCsvXv7c6Jb7PCwG1c
33BiiGbvBRRbcdYzjVtRAm9erHLUofedBGR/7kEqnRdEENsIaPnEvWyXm0MjGXeU
iGXCIeN362ag15040Z1AxD9LOIZBqKLqszU17N9tGqK6C7ZqVC8RLkPAtpoLn4e2
4azluf7Z2/KEI2Chf7b88ElsWqhUpH0m+ybc/mFb+auCBm3SY78RM6l38xjL5Wmv
BaGLgmcR3ngFOOQdJZbYYvkDoqEQazMYKw/ypeKJ90NtYbun2xUykO67I+qW/lwy
xB2ePFPl+WXAW1uo6BWQSMcVtHUk86LHeTy0th2o5Cwrq8eCKf+lH7n0r1bkBPgc
VPZCgAuhPut4Y9g/RdlIIKP73Ea2bNI8JDpnojuUuMaxun1WMERAKeGv+CXCU2Sk
WAnNt2M/RQEUNm2iYQXs3rZY+x78ORncjLHY+5zd10Am7X/eJm8UDWV/WvnVjoQ6
3lTipJ7CFsrRSGSFXbJtECC/bMwJVi0+2ew7xb9esmfBYMwwEkEthYXD6mR60LXl
surkIUvpAgvLNVLMU0+CIWnUfgQkeSSUFlXZsMRa6jTkDPdZywsrJFMc0aOk6QWn
hAEk9M+ysTbxYJWrvcbL/dp9zypvuMnKnyPtrhmqg+6H6CpzH143uxN8gjQg/6av
y5eaD/m8t0yP2n0S7bfsinblHjk2o1YbseaRuPxPFYpTHCRmvsdixHegp9JkbjHc
YaWMAOSDO1G4wnUBK8nEMK8h5sXJLb5ZoWkyHT5QiDyv/c+bECN3xUxxhfSDQaB2
kLnSO9/GLw9kKLUWv+JQzs7YEhRFOjb8h6lmaTHo/4edB/YYW6wm+VLZErpu/Uav
KroTvFiMFo1AJk5Z1LRGx1GQSO1JhDrOiBnQNVntybpUGiAujCNom4YlHy/l5JDE
0ycwVBxvyisSF+l/70ck2kjXeqU8J8zyhdnVhVGODYYMsSWkg8d/1vjSsPXm7kHm
qe3RuPmh09UDH69mt9/iONLYE/niTmvaeTsmH+ofw2MHkWXIhzgyZggDAK1Cg++D
nXjOiJuXUE4NY1BV2vTpjxCT+PGtHkOBOHtKteURT0oSZw5jybDAEwAB2ZA2Avcg
cHRKLB7YgqsuoEBmlK9kP3ZRp6kcdLkRFUyr/j7VWJ3wMicHCpV3Bmfj3oOdFG1W
9PdDNVVYwkVze1nJZzWfdBnVYw7eV9strdeKKaYWXYwbEgpJR15UmJ7orjoYZM4s
hLxd8m+YGK/4Ui6926czTN15yJq+CijoKm+q+oRJ14LH2TEL/DFQifXwfuaYe9K/
ocZR+pI+YBlSlHqyHNJoi8Yn8wYYMCVffjc92nMe4Exy+VEIHnKJnWyqmfPuSPcC
SrAScB9RRKWwvDpDQAxJg7ychtALbkYUh2WXewplX/oigujOTx4qc8mZanERhduB
wNKQI7D90TzHgqaS8OXcTPaWtQtNkBWIhZgDXY+liHNdjOmKSWpkrSskBnjxrrhO
OqR6tCDj/eiUzTBqrYohAr6PswE+cj8JfACjKCfKDabMwJsxMI2uhCMo/GLQYnYR
X0m+D7OJxdyqSjdi8Wf5e4V7SRvxWpda4Zl9dHO6YZVa9YGvsvC4k40ctkcWAXht
+HNQRcJiY3UmO/tzStU48YQsKGrsNbRisCQ6PKvM9fQDozFTtskp+VV8ukA2M55k
savnJSYamDrOyAz94xsUVqJ12MlH4jVqDgHIQTgJ/mqs1XR6scxs1zT79flSJzT6
+kK40R2+hkDPJQCsfnjbH8MA4afms3Pl433AWz8FgnOGKQpqrOPs9xZuCoDbUkWF
UHITACFDPoWkG9lOaAW/pPr1D4aRok6Ghg9dZpBSyzAsyWSMrPT6CxZxv0xW2lot
YkKGVA76gn7ons6IL/xV8pIWYi7BYuI+NQehFYa4dYB2hR1c77FgSJFVvIujHP9y
rg7i2Sc5MtvwZ/nzjKChW42VfboXMXadsLZ3qbTY56lQviDr9hqCk0YOZhmcu2AC
HIMmfYjivsd4KsucFvX/BNtpnc9naSPWYNyX9WcDFQttv7SS5LZ/ECawCSdqyz8T
7tQUWgiNE/IqfHnxC4NuXqJnsjHmiD+CzqSIUOZh+kefQV5131Q6v1dAe1PGWFrH
3XYzRgNOpjWEjKzWaQkBwhGc9CGQgb05VUyz/FnRcJdgIsI3BggSF5yddvzwGHUO
sPoZxOWOE9ypgNuT9qxecYj8SIByoxtmoC4w+gG19x8NjosElQ3mMkvtAIkswebT
VAR3QnyL5Ucr6rzxtX5imPkxpnYj4j+tfB6jYHbGHYU5ZN9efI8tywXo/iBYawX+
Y56CZG/+h9J51U0vpMJ3Gc/IgLIWn/laisW56myGyq57GYKcN6r1vhXrk/Dmoo/P
GunzeGWw1NrAPaH4Yl1TgW+kPTC6pfKnzXKS9mUTvogqr6H0pBKtULHV7ixjC+K+
ni3vV4FwjJLGhIzVBDJC30/iai5Z8E7XzIlopNepj8mFfhvOPteCKs4bLmJrMCT9
1MAJn17grscgV5Oc9IKpZ+6VjPFshZyOJOgfdNcE/SNQ9xKXygNtoLN6XpUjp1lJ
7nTuNXT8K8MPOA0D4dfejFr8nHwzc3BNQ6oLMPXZYfsuuA9V86B8WcroVw5kATNK
mWwKw86EXTmGuiFKj+KSjEwZHr32kv/nfMCvektAmlp6yRSMAgtLLMTKcd8k/ftj
9i4lHpbE6wd+pyOTPgtF2kTd3hHWjcW8ZnKtPgGW/dx/mWhn2zrfUgu2Oh/8sD6H
uMfIzgBdYlV4fDQOxHyM1AF0mF5LJCVN1jzA+NGVQ4RFEb0NzsBjokyEfq2wdNqE
AFTHKAp3y3Zqh92Q0gPcypA6C0RUbuUELg2QSWtW3YoFihjCffjgQUeSHLMXfKaN
m1bNG4dgzqQpDMhIzTHg/L9fp2/+KEk6kY3Jq5UlbCBXBKA3WTakufmeBcnv/J4A
yto8RjqOt7lURF1oZduQS1E6a0NjAnSVbIJ/uiBFd2y0ynS+gWvNMXgWi63VpLe3
nPd/4xxFpXWG19I7lhU7TQjDrvNLeLac/2vdzOj/v/tL7g/j/Pziyd/YIW4BuvRt
mP41/Q6CwDwlQfW+a/lT3D7qKgTK6Bbfp5krPdt/yGmcdD2RUEXVvor3YpSdQtNd
ixonMSbZFUEI5LsjqsJx2Ti6OJjPfx756I7mtiN0UXnEK1n5WwFyf+gv2VGRIWXU
BAVFGmYK7T5+GUASVTudPuZZ+HLNnoUkOqN8WWg+gfJtdr2NjIB8tYzQPFU5OAQ6
aiGcNwfq8kGvo/Na1YvGLoJUz4GWOrt4wAqFkPUiO7f1+/F57I4MBBTiiC0u+ZdG
e3mhpZmdXl+jpuZU190JG/UwIPOW8xfTUGXjfZ+ePCxp0dHm9YXdf5CNIbEvihrU
Djw5N3grDjxbyk9ooFfSEwbjAF9a4Zh51NxSVN5YEfRl1PXZ1h+1e8erDgKe9GRk
5VAUbDfq/48Wqsw8eSpnXDGn1Rfz7ZeHgZj1wlnPtU81ohcix0CXf5892fPwIcGf
kIYOdgkBrVrhg8MjM8AnPyM8DoejPmRwec6b6gjmoUbX0WoyBKIW6PnKqaXNM1gn
bTiC6DBEd6QnouvhbOfSj6Gf9sY18jMqapjDLLnlCO8Ad7cAHFWCi2XVa/0OROo4
DNU+3u7xKecfjKFf9EhQPIbp9kSZnx+oy9HjEj4RaIMb3LVqtJYtIIWJsspXHxfO
tvEFMuM8M07n8Cv/DgR3sd75EE0OdirfNHJsK/Q9bE3reRuLVeo5HACgpW95NCVe
eN+vjLElxI+WSnGbH5Prxh8FhMaZMtsJLP6PZB124Cz91Ea7IcWcdb+zHLOfHlwQ
luaD6TG1MCO28DYxwGwejBJpLQgD717IF86BZBrJLdvSfKUR3qnhCLQKuoMHb9xr
vuwf/DNlmO8pKGuiyUYEdmEJ5oQJ11fvrMjZ1wZRZNcoXIBAhPpfsd5dqtmCogPc
u2HxvHDhj2TemeUw0GoxjLMk7MHwMXwKDRAhVTKSRzlJ6sfS6eswvZIgIuw+clrK
zNCpMfRpVhkMARleIKwPc38gFhDO8aUMsA/i233+xyrHSRMzooNO8T3rWXditKXc
ENGmivnTsAF7VraOsB/kkMsKS01QX4og5KZ1pBAxbdWYb8M4nYTux6CU8j3GCQuZ
H6qMz1TQ8LR5UdhYyEocehdm4cPdyelPq7ch/uOj0wAzxu+zJxWwY75fPpUWKagC
3PozMsk4WmmcaAhmrWiMdGS698bP1NPb0q3Vpl6KIgRSy5uLRK3lLdOZ6t8nFv72
yuN49o2LIDJHaXa6M+DNbJhXTat2oO0relaUIxUTi3u8fHGBft+HaycjoPQC0o/V
Ue6C90oZBOXzUewx2SiGCtlIrqq4SWCbfaHN3gZeSOKIWFNjVlMm7hJ75UujJE3T
5C6m/ng2KvoG+z5+3CqUSQVuJK+s6cuHI9Ic8D18OjVR9L7JIP4vYCBcx/o4iS0u
RltkxP/B+rdfLUMTnM9/yDPSOIctUrhWwOwjXUvi3E+Yl4YvSJ69Cx9qInJJE/Tp
J23NiDCJTJ89P1rPtnfI4PyKtq4/KJiNCKv+lYGsc1IlDHFYf418S1gke5H6hwZ8
az/+KsT+8tdqUpk4gu/BIpczVzA4/zMXOj1Vu59SJmK09lSdSXc2Fw+02zWX6kPp
8q2GQpvzdnwqYNeV9R7gOjY2z+fXw6FrlJg3DIGZllW89w3ICQ71HfXaqRCe43iH
JU9t5xl4Z/0RhxnCZSsGddRrLKlMcmOvIq1zIXJSdpxU4SGqfiw2rbUSTvjw3xrP
qlDQhc6B8CwxLa1a+HjJ+xaVru/3h7zdjEwubhTkf36M6qbdW5rukASkNPPBl/1w
lGE+OxkSc4VcXQZ3bNs8mkwWE/VXTyOGFGGn1k1wBpziIkOtQOj4WYurYQQcb+2j
iJbtJtHT6f5h4EXjyJZfaQFqaI1cphH9jsxq3FjZVsj8265JqHA4t+Ux/PIK9wpg
jXhLJahnO394H1bLmwAhKdxyyiP08HH1QALgKezqaZdPcqzEUK5MGAEpYLceLWlT
ynYuWR6walFNl9pdsx6XIMhs9F400vywdVHVNkVTmlxQyeGVjfmAmZi+ReSviCKm
+hMEl1f8JG6ipeLXptLWx1+8E2p7C41JQEp12VGvcQ2ThmDM/F3Ys/iuK7Jrj35W
mo0+K6wATy4UvlTBbm5XkMQ5B7OcVJJYhqizBlkkTb1A9p9ghq7zc+mFpmAVpB0g
KOeVy+Tvd6EzCODQ57/NdS9/uzb0k53I7aK37/35qIbjlk32zktNORnuZb6X2qeM
BMs97/lsBa9E/uK3aEKwZPwMm8ToCTi8XQ67gpnJ3cwan85YNytd5lubyqLXCnlT
CO/zFUyMQu2wNRyFlt2znN1GnzNHaweleJFCHoN3WO4r/XxV9HGfL9KC52owzgN0
1JgsqgnIsyJiVgNaOSZ2xHLnciCk4VoWQeztD1OazKgTZaI2O4xCg3hdviNDuQQ9
U+EbHalV6hQ3dZ3uBIltPA3LWrXhLwY6WVov9zArr+8lg4iu/LewyHYhURl2V6hf
X93MrEnO500fl/oQQjMwTOrB+ooEPcKMiJ9xXjbDMZcn7Niiu0dWbQHaceQDy3bZ
c4luBmLq15F0Q7E71GAkD4KM0E6MpBxCTJbChBr4+Mqmpy+SWCKtREhcnII4wF13
wTeimHI+0907b9kPe/F0ZQkoZ8wQeKHXZ3yC8z1eIBxK7Q56WgLOApfoLHwhW+Jp
+ucV6hePDciE+xgdgGqJP3TbWVJL9bK5+vmzw9Bb7GEFslLI3kCGMexAHtVSD6RS
PRSAqQZmyRBzxEP1+zxFiQ/vUocKqC06DfW+B8uiQwSxoC8f2eApnJ71kwqlFEZ5
+y/TatBGpLWUypcayTvKytTdkZ3gkWcJ8zPaOcCYyAb/h6tS9oL5MqyO+eyxttSG
8oMo/kWf3z5UH+h5ulk+UupUrlJyfEtp0KjRU0IA2EYAIa7IiT/ICcqAFVGvyg0L
7ZQPbOxXYPuuwLKuXZAB1gi90HOVOW1sTwrsEMPZRcedFTp4aoxxbTnH8rK6AXj9
cgxxm2ssJXsvS0lYoAjAUOyFyFPFabAfENSrx3FM+0/4+s46XJVXxr0bCoj8Nc49
pGTNu0epDArBeqjkseLnXmEbZiRIewt5+meuHZpzxA+uJ85WjLaq9B3L8ayCjzI/
PbRNcjiAGZCEV596/4VKGdkqqNpIzJwogjCZSY54kEWROa0kl+x3k8fTJWZH/Yfq
tihCX/pKcR/jQQNarjrdrO5B7NjG9wKHWHNvo5eFcF9w08hF4tPN2EPlrjLomqT6
PcXdpspY7z5hybDnklG35DuaFyN23dLo0K/a4Qw2+KbOiR/96AgvjkIFlOnhiSgo
kMOp6tvTBhecXRVl7SKyJNdQa3h9mFM7ec95LvmQz7GBYpPQFFf6sMvQmvsqO/Z1
oFg9Gi48Bq3CDxgXQlJDMKXgwEbpOVF3Tfq6GGIWuiZ9XMOTJqKxBg24EI7ZOkF0
I2GIhIOorG4jmj361IZD4ypnELhFchX/1NNgIAdkF6y/FcTXQ3L6nOlXX7L2aXI2
1/bLYIQcuMOSHLxy43PMYWDhOK9cDxqk5q9VDP4g2oyfa3Gp+YSPNVQBjfGQPLZu
ym2tB3vh6BUAnau9I9BnyWyOKhBiGo2aYiiTOZH0VuRE6FWtfufX4vK6DRPnDpCP
XphgUBrE4/9w0/pwnc5gfXgfGPj4+zDUG7nGK4RU3cgU/ir0E2/BvxoysrDX8SFO
tk3JGPZcbuMkKGkHjGV0Ax7GRt/BPESddK6JzCecQftIs2kHiHPu2uNT85DPCu2r
GKDJuXbJagiEKStD/4KcrbA7Jerkt36ZhofWSvXQjMnjVbOmmnUIZ6ETqg8WGQc4
3mXfx4Nj51XRusBKTVBN4QZ/zjVpfbl7uAF16gPFJkEAAAS9U7INaDolpCDUVbGf
r2D4uJrVwenkNw1hcr5awMUe0ebuvuQii4sZfeooAEAOcTc6t8x7GGObFt3wV6Oj
ajFFkrw+qDLycxSuIK7XSZES78fA0uVFAGRsV9JEtJ7M1SywCGL1cWTBakDC9v5H
PWZuTvYj8wTeRv/RbiBZv91pZXjaEk7UpXMAZvkHrLjI/6j5ZXx4MYa6qIR8MChP
6Cj6+OydNrY6A97N6rslfKY6YUQ+5twxa/Qh1dCtib2EO20laEoEIgqMItjGb4BF
8G7mPZhhk/uZvhCSQ1mc3ELrcZKpBCJ3/gFIomELkH71R4KoM83XrrFG3prGxsGq
R5qqG+KIfltQBxkl5IVb+DfuFcFNuKavPtpmzgS4ZpoFjlmTkdoIBpJyZtdCH3ZV
UF4gBD8XuFiGuvAHm4XMuHhIb0xWvfD1X2jHafUtHp7aRu9dDVOeVm3d+ldE1o83
O6n0LL97/L8EFNJIA9W9Br6fG7xvzB/sBkhdKPFQoo7SNyga/m4r8z1dnfu7cxQe
k9EdEBwkNNJ7trIASuWC0ZYcsSOXMSXl2Py1S60Au3NuAw2Bmwn7ZTT5QkZcill6
7RkXgHttEViilbMP0WFW9usOdUMNRkDfI8ik7xShD6poPPQQwJFl6T+f4fph/pxq
7DK/9HXaLVqqjPQe0zBYj3dLsB5qHC/+RSsSEca9g04qpuDkrFvSUkzFX2IlhZZb
etymFYKaKLNIJgaK8DfIPognOfjjXxnoOQHK1vrCVyPFEUyc5RM85KdiO0d/0qbZ
Bzuox3CCyrZjaFBOHnaald9yG4VIrO4SlMZu7UhHJ0mwb0AhHy3MkJ86kpv2UVft
91m37pXIm97NAYlGo36SiU7lS3dlKRfo0o+yxV57Bk0BNAd4TRBsiMN9ctkUO/QG
P9Ozj67LQtEk/DLIop3tP5mzjDfjD5tPTnEPwsFA7Ob1sypF6NBghoRiz91s8Eyw
SydsztSVWYu4Spb7TJ3zYDwqH91cZP+b9v/FSXM0Jkb6mPOyjeYQmHdNL3pBRbAm
pKWX6RQh2Icm60s8+CIVapu26/MSH5/w+h7rq2xCCJ0vv1Jkejs4tSUBJmxlX8qe
BExl2FOPBbpHmr1Kv4nwUDrZXPpB3k0Ln9I9zs0QilECFJsh6iYFiJAekJw1YuM8
DcODLGt6ZaqGCcUNJq4lsVnvTlL9JbcAqHMaRa4kaq5Jlhz0mRO99W/dkNIi7la6
SXi5kmfKPMogLMYLrjEYNdh7AoCuufmQNcLJr9c7PNgY3ciuWHXOXtu/tHs9oHwi
iAmxXH5B+0XceNxZN/ocLq3Mw3G6o4DDynOWTNAYorIkkJ7kSnF1p6Ka/5OcVI9A
6PdsJBJbc1huTt+63QBBlFNZDVu0ZrwUwnqh3SaG+tl2ovhCb9ka854wrYYBqX/Z
+Ap3SkrYf9ohnqO2ivfk3faECVvj0NeHYiTb8PgnpcwodyLAETiYD9QmKPHWGzw7
UVkgbTnHAvE3l4mNmZpgyLGeDLOAtSUTX4+9JZvcCfoYIMhYq7u2g3hphqwFkFqe
QjjotjFU1RRHpgGI7N0XZAHdt+IpU5iolDQdGfB3pkzRUVY00jgvId0rSMOUUWFN
t2sbWLZvR8Pfb3rOQYXGHul/sReoSnHXW1s+4Uc+okBStOwEBbPdeDel7gQLyGXy
6mrmfSS23c3/UFr1/VpBp8LvC/m3ntF85szf++kEJMFEy85gEeTr8iU4V4YhT3Dd
BWIq3QCkYA+qtC3bnmAspuzPi2ehDaknviNK+m9tT42Bop+C/H3mBLAFesPzD5z4
5iDQivrRGX9g08Ey8vAdBrQfKG21ThnadwL+ykndOd7h4ij9R4+fYjES8b8yJuXH
m9drLiYqV3Q6vsZhzE3yUgYwLSEMGgh1h0iRCT5qiEmJlMW4B7kNc9wD4H/qnRsy
oXpFdiQFt27GFGgIWxrsWZcbX08Oh1839hr40V1dV+7J+wbY+Yqd1KA11UneSD4X
mJzpBvzrGHIcT9pLIfKsO+doELk/y741QUjqH05PMvqrnWSDkAu92Don4KilFEm4
NcuHWsFqdbEnZeFENRs7oZUxmDnn2RUcx3etl12QqoYys3ysGQFgRXd8Ojj6g1RI
Ej2sX+oM/LIKaIF5+bJGnCKX5NniVhONxKFyf/I9sxL4hCSpyLOiZsV2ToDHq2Qe
Gx4mOSy00yqkLc4Scz8m0fdmH6vVe39SerYxr3Lf+5+SmREg5tkpp+qqGPMFZHcr
qVPCk/TefGdiHEUkxLDz5xp244hDxioJo3QrdzO51Hx7TgGvMUtBG52mfVdj4jRb
0zS2iUzyKqiCku6y7uoQEOwdysy9NBPi2YShTfVM2yrXx0hSURbli2Rh7Xk+rvTM
DcplV3pP4oi2+FztJnsVo1l2PZSoYgP5ImouxTgMLbZokdC2yQQzf850En59WVUB
0MsY4n7XnwaU4MeKSQkWn8JX6WegzxYoLKyZBCJcqCF1n/21acw7Y2xXMthwWr4d
o8AZBQIqLRHfh5uwQLuLhfK+Y8AUecuIDK0MyFdHmC+zDz1tVCEjTOSUuGkK6hfi
Y/q86qCGqnLb9LHIrSM5erH3P9WD7MYDhZSJBnLcsyP++FMQWkhCMglibbDHJbn/
Qi+nrLdmAy1SlszAvjOgLKUElcSjfNvSFiAcCGw3Rn8NMd2xgV6Ew52HiyDIe4wk
KGOjgjxnP1sYggk3QTD655L83oyl0tbkkFojug7jgS5TUI4GmUWaiJIZ/p12E1Gq
6ZXul58XSGg1YLl06JErEpRKw45NvyoiZ7KkD4zqGiMhzrPln8GEmea15mh56unP
LVhdNYRIMrywZc+U77FaLQCn6nyZWE0sPGdK2MQGETOKQZPqtUS2IMBcUTEx6kQT
OBMngC0gn7nFkxBFCPYVWoKCBg+LcuIQrYkY12kVmKr3DhCnxMwKGoY1Dq7fj9u1
Uo21nUPdWzlFh5HIdGmMdPjYtAC8Wcy0h5QfKH5nlNiZbtqq41PbHnesylbIuU/f
WlqHHH0rhfZtrGUlPFsmFcnGk8ZmblFE8qECGKH8RLChPfzF4IPf33z2LO8ppeFs
1XICeuvO/NXRMX6SyeOCXRl31I/sGKm2IVhdqMuf7o9o+jj6S/gqZIK2OCHqw2+T
H8wglcmLMEnoKMg+rBrUPfEOR9Ck+EFmUXkZBT5zM8e4GC6kUVY7WCmJ4649C/8X
larINcYiV01YrXd0MvjlmdpmNYdrVoxo4QnzFGFTjAHRSuIvqH7zw/kbfju4bJeD
/c7T5AFLm4g59sybUmg7kWpPqWLbhqUBlgNnQ9LNM2a2BnFJU9Pz5OfaCyaPCvUd
6mzxZtzA+Um55DPIFESf6t9mv92qqb1lC8dI1xPJVOx4rCwIVkyWQ5rfVfpVhQ53
3cPoQvcyv4EE8jC5//Cvy2I2jw6JYKoeG3URJ2kOcMiyscz8/xJHj/FFxBRKcVmj
8SE48yBfMmZbxxUfCsQ/xa/H30VIaKNMSWrFP2wg8JcgIIH2AVrfi3O8qM96OTQE
Q6Xzpi9zay/6Ijb7m+9G4dyaGIeIqKKnomnzVbuHSNXWLXF6+WRTJ8myIckOap7b
qU8HRiJJDoBCubTOxTRh1McnPrBNcVDFdUiEMzLEJVbhTzrrVwHpdjIX6d0VevlU
tk9Qjo3FqS8HmjeisAB/TCrR4w+ilO0YvhfaNJMpyZ12cheG9rEWcM/GPmcfKcr6
zMspJ+Uo6RZxF5t8/YnJPzlV/2pqVLYqvS/F8llzXTg5+l/lAVAG4AfkfHY9yq1d
JwccEjcUn6SCD9ewBaEHEG6WqNsiN6vUPB/PGPWMCDYDbdH5BmU80LGacgQyOKOl
alQ132pDWPpwXjmqHpu5KryY6qXZmN1KaMJushhBN7iZSVypsnHSTGVGBXFcEBSH
2B+RD8eQKo6AfCe748V5HvAvuBkW4x/34dcDZ/NMLSP27h3YdAldValIJOUGvmxd
PVLf64nxZrd92mOwB3EoKtvUGK2HIV32Lhq/hFEafg1riKp9LWDUdQ+LPRCa+tZL
1Y6AudSOYnwNjoEuBep35qzVzas6nZcWRVDY3vm8UE6X03J1QlADVCoVL1RwqJuR
ViqXhafU8radAd9Wl+d93A+TTIi0FGOY0Duo8DrZFbezOozWcT4XfgpsHXpCshaj
+uhqrUYpCLi/+pGlp/uz++lH4JDHrfomaR2AimYDOc36lfl7lhUcT8ZdPBZil/u8
S9qU7mtOHXEbX3bNVRcaw/0MmpbRaRmGKOHsOsMQvnUqYl+vZHHNS92GttzZScru
sJkF2xXyqhxW3lm8x3mBXnbsVkBRZoCoxFMhNk3PLLag4cgOvW1MVWTjAxc7iT2K
WJcm9NcNBSWlTENWQIoerjF88il+IZD9XNul6AeokaxhZ94+9ylnR6McDUCHkoD3
Z0De7pbtPjaF4BFKYBmxViSNilEjtZiFaBRnZUqXv+J7g9my8WZPeJnPKLZ6lHLH
3/gbNQuoRlKJsNqAbMe/XHtO1D0Tt6LWtCMJu6sPACONGQ65D+57NQggOcdwBVv2
Zz8y9cghfMiIq/0iZoJE1tjfZ2m4e+Sdn+SGMegqhcJnrJxMETFbir+PRpLu88oy
zRHyRN6+1eeDKUi8IrnoRYOA9BVqolwY06y/d8C8QxYjjf68ogDVbDtOf7HZPzwB
+o34tW4FtP4Vc9qfHCGSqrCrnK8pld+/IVqHMoLtyCca/GL5UYzIIlOByp3zUoIc
MOGpvjvZI/A738ZLegfO/7uQ6vpaeYrmu1/k/Wn/LcKo9lVwi4zTeodqZ1K2wYLM
R8DqkeW6fyt5iW0gCxWkHJBmnxPCl9k6i+Rg0yFLpTqWm0ZW1BRlm54FlhxnDafB
UFJ6sUS6y6EVPJLpEV00Ytj5LzR4aTwgeRvll8uqMf8o/eVDP0uiBAJp7BuIb+ct
j6uHeaBe/pNnKEcxYsuUhHal8XC5WxIfmDj0L0s5ByR6W5NUSnbRHVQHEwH+OIT4
0AY+g7GMH8+lCFdHRUetAzjD5750aIVZuqalktxn3L6vqpsI5VX9H5tP8QuIvVZy
82y8fJcxl5VICUWm37UHUrbJ/0Z6paIeaEDuP1e7Fi+jEfAoa+iQaboD3pmkglro
bgiuypCX2uNhl4Heivh3zg5AqE0qexsobiSD+8WcEPCqNOdXQX5NVDpWOlhH2ym4
ywlRHw7mfY0o/Nh/J6il303BxZJ8KnVEsoyCyTTf1GzNyKPT+d5WI7kUYTf651Xd
xePkTaLUqEbTyif901kxas23ggERMr0NQ+SRJ4zQlnUFTbsQb/WuGO6UEn+hlSmy
JeBcrmF0uUM4VchUS3hkDwKWb8k0wmfnGPSnrDJFgpox/e80qbcmaQiL/hAKqyQa
1jhMH12bcjDa5X4pdv0+eCQTmZ2JuxtSntBBRb78vcsHtfC6uISQekgKO6PxSyn1
8FdHFSDUTNjtUqu+2b5FLsECvRWaCNAoYhX6Xl8JoESZONA8JJvZ6w+EWnolmIsd
MjtUwRSovvV0FO7CL/1omwpsfqxy4w7yS3bWfbJrgKJMW/wkqMkxjEt2CJMZVLx4
/3sym33rHOzCBeiUoTBvl9NjiQh5dTZk6kka4vFk7/VwAIIhU1OivrFwDE4pjs8l
GtMAXnBKQwyIpT0to7VvDEvJBy7mp5QBRkpCTZrkZGW0KCvivcsV2OpWdNLcGi+e
DofR////X7jnUftOV3gqo9mu6UIqX2r7h43GJB3YVLTkFR2FoDDyc1BMXEDt8YGn
XTv7PHtP0lxfGpEVsiZ0OVqxSySfO7qs1pCo2NqZXkWLF5AEHGctj94IrfuKoiS/
Qpwnriedy4FaEcfjoglEgiHJ06iVuxPLQwxJPek7OrijUV7DFocNMvG4bM68nrOI
MgoAh+20A2GytCCElzF0jX/l4XO3dMjlUjAfpOL9IrI6wx138PM+G8NFsBvoH15m
DTdRDkbYfbXv8QY2LBdTbpPw1YosU+ehodTj9gwHy1SI5U9u74VUznLYBnIVYuWa
ldy5ieAfvnK/FReO3S+smuk3o5yvoh54uIpH9d4P5q3LEc/QAqjIhzB56EpKRu7w
0zxLYOc3AkH54kfEchUVbskVg70YEnQZPb4KCUtCjTPWNJictvTJyTj9396HeWRy
qNy+KWwywjLBjkAa0lImAZVU7dGjRCWVOPV6zff3/xtw6xqbzX41GZm07zmBnW4c
wiZWl0bA99uz66ZpY0ux/28YA8c/7tQ+pqyfI+Xh2Z4ZpzRBwpnKMRLgeLzDt5UR
gyBBHqtpW6mWA55iehQQdfCDL/MeY5rEpkl6qXODOTdpfCV+IZjr0WBgcq6Bjg2q
BTw+QDRmQxyRuc/M4MWTafijooj2hYHico5s+nra8/4f0A3Q6TKK7wt2xrPBp66H
hNPIluCJjxsUKDU2DAw+ktQmfsM2qLZ0/9ZhQYPMF9XbJupRdP4aRA+ZWfaE1ZTm
IiA11qeJTJz5ZcpAiFRGBMTDF1EQb4TmlJ0zJawGZlkxLBsdzdiI0YvFI2ES97Ua
KOzxBXPw6BybsbkiwAu5rTfGDuxI5xr7RxxbcjS93PYzUxtWBZusk3SvVdbJNEXX
42zQcPpBnmC/gyfgbllVO9R4zEa9/hpuFHMOr4up6ioy/8PCUI38klSiFqpaSTvV
haXT/5/HKosHGZnpns0NzK1BCCNg09QIE6o3bGXu9oNayxFLFY2IazlzFUd6wOR5
I7F59d6pMZPaGjkhh95UY19TJdJ0tqzKUSU1qSvJsykmLy/zo4ZtGbVS4Tjuqzoe
Q9+Iv9W7Ap7N67k0hJPi7wOoJ7W2OiSiijglCY+Q1WzrM2Q13HpjJLUY2xPCwt9M
UZNpg+dlaTjF7uVOheSNng/VT94rxkLkWYQldOQpHTa7sTjdrh9fiHA3LAHsJmT2
N+UacOtrMlAgC6+HrUDP7aFNU1HHlPkdP2cHn57A4Px0HS/2xeqBhmWOnFVeMJku
Pdq58fvxtpGo7J/fL46yFQE5mhccjhvNf6nb9dufid/qRivXa7On1Og6t62pCtN0
U5Bybo1GcB1KIovUTmcx6GI/3khiv852ZOCabWNo3recdYX7fbBGzWKbp3qJTBwa
hs0jzgv04p8L7kCTo8iRmmTrx6+ggOCTnfl4nkknTdhk/n6SKZD2Sh9PifNcQWZM
Dz6nXggrEWg/NG/l8+j7PrdffwNe9dL1sS/veLdhv3bkEDuZuhlduMEUmXpvv0KP
s1Ne0y/2bGVJClI6UVyU6tuwJqfyMeM09EszfLP4r+9jSHwX4Xwdg19mpcH/4w7F
8zycBJ9Lwci+kyFoudjnmCoGsGxMFsEDPDg2q7ImbsRwosZufMvMFN8Y0qOluDDL
o2VijhnWeg/ZmfsqIRKQTJbbnGogd9Rx91YGYEY1VkebsH9KMFBeprzp/1j22pcI
VAR+G67T6zc0Q9J+Vvp/H5+FteM4/SAW4I5wveutVQPf51q0KQG4RYf/DzhYH+WX
2pJQKmhsGRC0fq/6Pq8kdPm5Me2WYtelGD43YliabWEgMoMjT8+ncn/zkQsPnQJU
PKETZ7aRFv6B0S3JYyu8R+ZqGBIgA9N/fDfqDvUwYgiHDQJOOXzeevy04VHdoS8p
eh2yU0/z87F5EM2T6TQJa40krBd91+qkJ9HgIwk44Oaj0T8C/b+BTpKgY+jqVrUv
3DLDHgYBfs9Z307bpnYJGkM4xLZxV890nBc1z+vMGmcydI/ln50FKyzbLlDZqX17
nR40Av7dVh+v3ycYyyG9M+fwsI5kAv28j54RoWvWA1XFnz/lp2X8wh/kN+kMzxjq
aJVL74Kz4IwGMtcrluSXJevbWdFEeafk7NOD9bLAR0WtmwH632sbCX/UUBqS/gzJ
12oFFGiT1z9pEnJT7SMubOSgd7JrEFbAPjitXkq9e9s9/mn2AbRKl8JmKNjBxlfn
3PUZHeCWrTo9ri5kjgnVBeqoJIReKFmW85bd5RuKM2T7kSF1HE9LdIXx9fq9/LnB
3bcofbod4BsfXy4jnAXC0qHpX0hmlNWO0WWrYoKmeaw+vqbvxdd7uVdxSHEcPLuO
Bxu6cOnmEb/C9HxO7uUrNrHbOUxfbtADsWmiv1BK07hxH4huaZUpoI+1hOjmR88c
laKXzLE3E2p7mMSdQBJaoYbq4r++iJPpblss9uV5qJ7w1+ZCtzp1MZu66jzev1LT
9twhm+dsV4da6Gl4861vbzPZppoMuwjQxveyZbAkMQ5lgs2SV0yfgLD0pdKPi8CP
TR+PZloy/Xy+LEeTCl2q9FPGdtjq4D9y/n+wEvyGIf1NyiRK4Hrt4PhqOFBSqIgO
lnXPy8F2eUuPUrHuy3WQ1aqD3Ey9EBb8jPfzbbPUhHhaNsjGulTl+fjsv/gCJIiX
7fYYEqh76NYMTgbKm28PePpI/2dvTdaoklNPfw+5KVUUD/HOXuOEKW9KTOrbDc4o
fJVPf+xAnT9I8+yUv/mw9y1qJ2+WXijrUSWrBj3WShuEvBP90rpYuRezi0w8S4bE
ZAd6ICNyisvAh91WeJ0xK3TioE3cmnR03vhL4ipP7djdSdNtQUSDjbee2ILzlymh
efcqP1YMaynGTdx0YyylCWn79yIZONnFeuDsufDIhbX0oK4MeYSkGfsCumn0RLpS
13zJcHqMUFfzxTR4ZA45MZBxrcrGi25V3l4zMLPv5j5Bg5mCUe6N75aq1BKFqP39
6YTkiArM9CpToyP/t7zJuz7pgTWlISiL83oZuVrCBWLx24On3ncCmz579ZMZ6Tkf
/c1nmC3zRAImH1kXUrX1TXWVdE/ouBEjC/NTfpDJJleOu8UcFkTYutqfNnjURbq7
KPNH1A6HuIf837HbH6UmZSVPWjawcqd2+SWRdaQIsTvETfhtnRbCvLQU4VfvWwno
zkB7LcvorrrRc3s0oB/+Jcv4ae732yi9YgDe3iGywqTEPaMu2rA3Klxi99FppIc6
px7EabuZm9LBcjUjh1cnywY+1Z7Q0k3iF1Rj2d+RFCNEVXy9UUDUBqtOQwYC88Bt
pFzrqY5IhjRrlB6lUmNQyONfteIj82KzoqlKerMjHiQPndsoQOxkWOvfO0ewkTo4
MZmJ/pTxtLgxrPij6CNKYWH8AUgFy4KMTNCr1HyzGzHgpJq1Y21alBXXpWFYSBs1
I4dbqImCXGcK60RDgLXMVZ032c3T0d+J1KqNOyu6jQ2C6sORlzBpPlevWNO217Fj
hIJV+jBkAhvgzfSQ+4PK7B8OaZOploJ++dWwca06eIHu36gktn30fJTloB5LZ2WE
pZQ/zMMETymX+lQL+QMHbBdJHuXKr9aU/O/GjzYl+AzHKsfLvz3KB0Yi2FDKbSTo
VRlb4CzlNOkbHdqfAc/7BbXCBP0HWd0NtIjrnRpCwDLhHm85K9rN8eKxgdSBzZZ6
8PGAmNsyW/NEVmLaTeNwBYlzCoehpArSdzd3vGlH9Lv7jLVsjRgtsQzJ1R+rn5Fd
zeY4LtGdVNoDCTCCG6pFK/kZyTJXlX2iHd8zkIGMgsy6MiE5VCcY2tzYH0ZaQXW1
vV/4vdvBNQBG2O5oilo4zh5VskKNzVxAvwk/yd+r26laxPCUpppKlQV2ObdaieVV
QwQf9WVA1rQIxURE+9LYPq9WeudbsQljUzqSPfPziP8vepnzwdFuwojqEuR/sxhz
oyHzTA7u30PlYwBi5xOYq2S+noN5RZejolE679S1gY0Llb4fGzhL7cHlLzDYwLPt
PKqSmy9X2Rv6VKAZEyqI6T/A384Phrlv9Ocs/vVIETqHNZvaxOnsoFHxQtAod15q
hZy7wUDdHf+14g3MxYoCvLqOBo8V6srVmMrCPFFOR1f50tF1HvmAoaTGdzKSluLO
kkCmE32wPX8MEErIPfEmyyZi7o1kDvdbJgnzTVtFB46J1U1yUcRQnIF9ONXG3WzQ
kNPSTAnmgD9JlpyvtEK6i/rAAkjbzoK2Racsc7GVxqDSfYhCATempe0WqVUD1D5t
qbmx/iS4kMQD60zBg8pY1SgzYvXSz4xdzmfi4/9Ts3h1YFbTqe1PD/G8qnxqUYN+
zByjN3srLWLeu+McWMwebxNeHoxCp9GF4zUfsuyaGe5B555Q8VPr2hpoN3SL9BDY
JD8zGZat6oPvbKKOm4OYlKISHzHgyv6ya6BYa0a5/M3BTqQ+XvjBG4FhL5JcVpUe
1EMd9mT63fAZw+P/Ig6CKIdij4DgI38XbE0hvMaycQHueVN+C/ASaTgIea5rzzhL
StuncoEBCkt2zQlNwqEzV3ExiP8wvgD588aJqUPmwpYLjPcETZVt5HNDn9u+8mXt
1+P6/9BA+MCbzT3t1tHaVCmm02UNOaIZpe6L5fvWo6DF9+UsD6iPTGMOWi0pb73E
rwW9EzwnoXORBp7Ga4xFYCqy/LXscmXAiky8CJcfai9/DHPse/NYhayD7VuDqPRC
UMq3wIFWW3wvchkX0li7HvIWWRdc3ekHv4cP/F1EQW6Z50zb4wTwiSEf9txiE4Un
XPTwTvjzq8vgEnFFulVoP+yZ6wfZLzHtiyp6P5g/wkE8RL/RbA73Mb3B4aX7OyF+
5cHWtsPl4Ism6Bx0115FIymdub5EjYwvX2XYto8Fj0Wv2kA2V1iRg3J8FNFbkjWE
nBhkvKarZaL0U9WVBw7CyZQtt8Wuewj7DfpbVkQJrOEp5wzQywjSMaEVgIA5eB2i
hrS5anc0AG/j+b6atghA58AlGsdbp4aYKpy69kdF3jqi8um1bImd0CTUgByjIW6T
UwO/VSv0OWZmmPuvBAWe3s+kPBY63IoL/9uvlcs+Xm6drTkuyfybtiVzsi/kR2dO
78qBWQVSsydxcsyXeWjktM0irw3/jZjHWgqCeICNxlf9w/bsivylab8+9sloJ4iA
/v/J9FvL691F3fQloM2p4U7iHOKYfFcKZmlGgv4lfj1ZzY7MuUvQ39MkanAhw8Xv
mVDzeBJGJcA+y6fYz4rIFUAynNSEb0shANhkGanyPQTKQflEGFnw/0+hMpfur0FU
DDCBvEYGQ3MysxhjakUJ1PU/5ZvKV48DkT0W5KGrClLJXtL4qu68w6QmiORpGTjA
CLFuNtmf93EUsFu+b14gZK/i8K6cbMeKfIPObTVQ997GMJaFqsoQkxg2QYut9P/z
0IjtsQwPMpw/knp4VLR5jh4AgxeN7bSYnIYibyL1b/R5vhum7+oVpLMqhFpP+q4N
30fTbltUnEzWKEuwbcqgjXHG/sOqk6xsq38HxyThmeMS7MnL7GofVqkcJhm4TVcD
gJCoXpO284SyyQZV4bMXZpnj/fV+u+mLkegvnH04laSgHcmhyaUeCHhOjB14oTNf
ocsdF9Jw43Qwe8jzf1EqeTysgJFf+3ipZn4h+2k1Q4OIPmh9WAgkvICBHdiNHaX5
VdTNq3CCH2//YD6v7/aIbR3pXsKRUOU0BeBxndD0sb1c2mOXBn94RKV99MqHRCEE
H5E0lQfhppTSvQxqU7pPm2Q8LiAGhODEKtpFBlvrwUSJuOsjCIVuNOXjYHspiYNn
qw6hiafslb9QPAtLNSVwOxrNjz7025CjtX99vwvmkc0F0agBq2swkcqtamDdQm45
Ak2+oVz81sIUm7US+niihoUqsEdGjGtsItcpdMZeq30SQmTnASsqnt5jSrMSlRZ5
ZMkCsPhTIGm6vH9YIfrR/nV/JQ0jQduDLJ6js3A828ulkC8s7UtUqPHvKqx1i8jb
s536VQu+Uh5LfiMcLym1D82UKWUN8CIxwHKRW/ua0j4rBRvASiraAIIQfpBani34
ZRLiHSd3WpEjv/A8/1DJkzByBf8ebU1ERV8Fsqru2G4mumgBx5h8xxFKICOOJkSu
ekcCU/Mp8aDgU+bdJBioG8QBGMOLwysG8/jDKekFAQ+R3cnaDQbSeL8EwGUpyDez
WQJEI/J9eeJJdnCvi/7yoE/4UNb3QTajdoqDvkBGYe7kldSb7ljJ1WT99Ian2P24
zXIOu3nxVqgqgp3cym6s/m5VCONVVIv/ABaRyJARoVbCCeV4SraECxl/iFrNWAST
pUhcwCCE8OSIlUoKg9Io8+XxgmFzbHqJXcVKADVxziPc3/Da0TnmOPVPfUIjKyEQ
o9gNxZJpbYSyblODNVjgC4Lb4DYA3aZExBG0X088ZcMkLxpILYmAYPqmnOrNBGII
DqXbCfUEK5fn440dVARkLmTWdfaLuFqkW8ReVRPOKkVjY/sf2HjTHCPnQOgVdt0v
a6BudOS8uwo9b16NmkeSiO3Iws+ZOslPMxD52m5lCc2AS7Y8rKqjmZeT8CoJNK0/
NLESC2K6hSprHt7Z12Wm0eidsHLHIsmVlwxRzci/foitFIpBO6PNUw5Py94Pe3MN
ZwvMcf38NueHNSHO1ZWC8qOFBM5YSGUzZpNpm/9iUI9JIgTMbAhthazrA4l2TMDm
F19GTIJ/25Cui2kXJmtFrfmYCFl0pcwFhLhrUsbgyozxh+PC+24SSJJUUsmttGla
DLw07Jix/uMCGUD6OvewO9CYZgOG7VVc1kbMwj7xPiECeulAMZzAnfOQ6Yihso/j
d/hyd2fW0S4Xl60YExpZjcBVFKc/Uc/ugvQI0X/qrzIfZLTZg/UnISuM9pvw90Qw
T2wagUyVqxde8ULTmsrgnDs7MoWK5zbA9ba+FKVt4RT/F93klcqcyIstby0o+uCj
A26y+xfu77tWH6gIC1vwQ0r4rqkrx9DW2+PRb40rftoQ+l7BjEY72M6PZ1ifdfFF
9MQZU2yVGahOSxS9PmHw+TJV9a9aut7gZsBTnS7uQqC4BMKbzqja3q3YDuXSSc6I
KFcTYOqkz+trHhROvmj8k95wXQPWGNB0yOni2pAzi3j6/6R+1wFWo+j6HcS+Qcx0
y3L/LQCljC3hZ5iTSgTzExgxmUYxLxcSSMkl9aYqhgKP3FFPepLpIoftqmI1Pv11
xtEuO3RDyLFu01SQeGYYXbSwCMsPgz53c6WO6khI5DIjs6EyTrAp11emGpoOWiR9
WrWvDUiBOaJRd+ODK0mpO8Pmf4gzb1UHtIu9wQgJeunxFZFVzuw5tKYn1ckJJa1p
hPI3MmmFPeMren8S/C2HSX85sho8l/2pNkqWMTmixk6ThdkH+S+bspXt6fzEFpj4
lhB0vq2bXFvQSIbacrNHm3OXSt3YogoxvxjQ7LzPWSRxzRH97RBt5cq9SaKOymLB
Dcf9hOmXygNOHAdzxMQI9x8tJ2imMlhk8mX5Ppe2f8VUqhG5jXBT7usyzJwU8Kx/
Vgd9w05IaTWaWDmMf+CNjr/pkF4XgmE8890OPyqUwII8yhHPKDjyPiVIZ2HwOlgf
RHUvM9KK+n8Q/Vf+T8F8AtV9epXU8qFZblC57qwXflC3CChVJhQ9vdUoaPkHCL6B
dJRqu4mgId9TOZIBQ4ZWYZ+Ft4tjYkE/hFZh5R1EMi4stMES6aWMHIDPs3hcHNw5
jb5IgdvhS+IP6csknuLkipLseC70nH2r3nq1IBa3zTK+nZpUgLi78+RyjTaj2mL9
NF4OoOflxqkvW1z69+7cEGlMIZBfU//qpNo2kB9aUb42ZS8/BF4nZylO0jQpxEaM
EggE57KF6f+YIA9f3NuiLY/EUux59dTyPcpDVQiLnRxGs/hB77kXNuTuZNIwoMOp
aKZRxGNki11u12RWD8kCbLfY6Gb6lsXHrbUuRveHQnwvIwLe7ExJvRmTO4es4Lhs
BdSJisCeMxRjp0qUzij6HA1nZNDhbKaC08q332LmiDEmGk0E6kv749F8STC1RPxg
S2FSAW/73W94A4UsNb6jhwfatjuL26hixCJk+x8o8TX87VMNUDhnn21hRgszttOG
uASb69Cgdo+wos5CcREnDcFXVNxncAlSKMSFnejQSZdXL3S+IMxvHhBDexQ+Gaj5
G2bJ7zIi89+z6rRyK0uWw4SMJq8tWZNaUnreZKw/RyL27ra5SKCYaqYhiObvhEii
LEwbefqlE9nOGjZ23R5e2yfWXdR0PwA5393ZoBN+i03no8R8qiw5bu/MujO7p5/W
Dz8Egi5d7aGq03OsZ/pMUrTsOiKacCRfQ0xJ8Cad0niKmRfwaYmghm3Jv/tSr1Dd
RXJHuFJRmW8+02jnWGX15jQwSNqw0oIgfJ6l//3gfTs0yMfIx+WiZKO55BRqBdm8
VNb+J59GyQCc5zieH+UNyrCO+bgT67H47R4pRcMJU9+jZ3rtWwbhGfLKfUW6cyEW
V53vHGgUicnQW8b8Mwd7M+qHWibjvyCntHML+DtNc3mFu7+JPdeDspEYa+IQoqNO
qWvZN6hG2U95OXxLqPnGLcsgVWtXTHSLH9/g86nos/fI1KE3UeuEfWKF096M94RJ
Sn/E4IRqomQ1HgVEzquchX3vd20yBs1UNE6d5SDtDbSJgJ6zatAGmVB+AhN3G0wV
zIzxRSByjz5Z5VzhzCseby1Zn5J6V1PAkpubNKR+yLfWK/ZQyInZtJwBprJR/Q4D
fpR0mH2odlY6IwqSwucCoUXnSuympZBDRNlQfQsqm+VsSkmwl9mN+2fC0XAOBMPx
EQaBEKyhtRSS2CV84v8rthkpdAIrmk/nSWa9xv0pmiWimVwKOt5fBv/t5kL9bO2t
+3R3ElekyRQPHLkqn7uvEzqsPtc7eBcOcRVunYytgYC7qA9cwyNc7/z8+xrDsvf3
AUR2yDfygRZAJysB+VRb8dXgoQz/zY31x0wruwPnjOE4NoRBolmevNn+PsxJBEAR
FSUQU9FlpWsC0ahQKN+hYoLth+1S5gOZ8F+0iScn2febUcajCA7HtPraMjXfGd6s
DAuJEmY+h3zf4/WzNgkAqQAYWrLYS1f5GSs+8rqNAUYuIya3BQ99ok6xBsfdEtKM
HVFpBhxXnuaE2dgqVipV3QW8OFcVdh+1C9ui5hVGc9JbxllNwIE4rQgaOPluPq94
CRlOaIqZ65lMWsYkP5ubBNTCFdxt38c34sqKIg9F7m7Er3HMoPPTB0fAK/PQ1R95
uV4JGmKpt+FcKjWHz4iAfhd8nYYjCaosdoqB+h1pEeK/WF2tit17B7sEUSFn1CBX
yhi8dXUf4fwOCZrJAwNjhabeUtn4Oz2aa0+Cpw5tp5EawP/7MGwZxFGEgSn9B2JZ
20GqjhQD+fzcYJHghrp1i69zDwvP1mh/F5OBQL7kjYKgS5AuE+qDSFQ/gJYXlsku
Dkb2KwAzWa1b936SL+9KYzClDk3YhkueykslMLhan18APP14Bew8oWDuSsgXPnPw
iXGjo/kzD2Q1s5Sax3w0ubHbB6OAcGaa4eF4YcpDCZ8Oxy8tiE2k3IKG19ZVkS8b
fa6J+X1tn8R1HKjP7KK7YQH80osrvBWtb98rdn6DZrmsqqSFPM4R4VlCifBZc+P+
Pe//KC2dWRM8+lDqAa/eoxkUwvxlXa5BNkMEy9RKoiakM6eKWvhK1es3Asq2oHux
vmxuNIRQDWo05ia7l9XJ1gxYEJIV1AKT4QXiZY/Ypj9HDZEQIflde7QDmp2bdAUc
wlKRVaF/zyyKoBfJnJPemdr0VYIAeON98+Zf0/0u5t9bQA9vIzXX4pebzHTZofoV
+bNnKr2BijnS9/k6pSsFlX/GjGRuS6latFjRR4aLpWOVAY6ntwUGrKZR1ldIvJbq
WMcnQKaFQt/YlVz7hNrGbkUC+GO8ClI8DyLQVukxF1IulptDntQ47VVdNAUd9Zf1
t/hgBgT0UKLOumvPNzhwjWqxJ/zqldyXXVBO/2xeRqM3RI1zeDiozCxbNphC0SyH
CquZ7q7qHgZ+hyqXqMPfQ2tUGQB/hHe+tMgFjfi7QVfZrpyaNxNMPE1RpDzleVGf
61PbPT9jNjbctAestxZUq9vSKJyczUyOIuHZI/aMFFHrqPIhQOrrEPUk8rcXuyvn
R7u9s/neuwVOrxCJ8Wn01RW2ma38QI1BuhJo6ALWxMAv5a9oR8oMvwkhslMHDusp
Ec6iJnR9euLV4yftnOLVk2/51iVkEtueAhXdFiOUUgUpJknOREDFM7TeDd+QT3wV
nlP5TwL80OUJnvDZ3zSLlNzJydXFhGZSQaPns8Kohzi9xcV7O9EgzcWUnUmHu1HV
rCHLFlEr3+Kr3hVtPVUBOBaqGu2GFsDzZ3nHCozyjvcXPzKTbN814qwzfcAZ6moq
dGrKUedEXg0o6IcsVjHGJ5My+wBwE70M4w1I+Vhh7u/8/wAQ07Pleso2zhRQbWA9
WjhnKStPMDsMTPAUg3j00FqWijmVFjDZZLWR0gpdwsddftQOsMkjzm3CcM5S3CV5
73IbArGIAph+xS8q3sd2UKGXDPSQN9D7cpB6B3JTgvltVuXggFGIP/a129mMT/Og
+C7FWn/HWJOSYgm4tq5p6lAraqInGAs3rirlvMDxx0fBjhdg7ayJwpZCH8rNTa0u
z7QYhqguNyyZrT8Rtrsj2Q4DvqNGyaMEFK/7VTX35jZv2zwziJ9g8ddMd0SyjLlm
ljHzPFcqyLuMZIP65APaT4xw4CerNKmbqPW0eLd/fWzWkyD7LQFf2P/2PfMrQ5y5
XDZw++S2ZfJ3GXBlvfvV5iV0/mxBz4VsTcy0KDmLsLfJhXLOy8+airYZU7LkHvsF
qb2gGhoemWURTu3Ag77TfL1KnfHEVRxObOVVOEADjX6IYqmGOaCHApwinURtE2Qh
cZ+Oz5Vizp0PNwrWDzXg8YPpYUDAaVR0lFalxgWqjLSLmv/xlpPLcO8wfzH8IKHi
l6MYIZz+eslzhe6KA4q/ZyCYc+9Q6i97hEg1+J5/pwtnXBCXKBXkuR4+3oNmnol0
GVGVFsCgG5fU5DY94mjdGakWET/XAfRQJVFIM3EfyP00717RA+tudnRApXADyFBK
uelizEa5a9nmMZ/1do0FHsvnoIWUrs0jylWGSdeMB2yTefmRDLC/m1RYmoC41Os6
rA+4IZ93RJIEeJo7mgbh7HnJuI7F/yD0ylMYTPZ9RFDc+uIJTqc7DLjPIizKVTSU
Z45Du5drkYWTyZfx6ILb4tZldFgZ4oF9VEUx255w5aJoDbMgeO19SmOifCQi6SAG
QApSjW4Ob5XBJmW9LZ5raNvm8bgIy3eBUDOf9ByggO0rGfBWf9KqO1vWJdNsgZMt
vRR7TwdYCslq+LLxcRrCPZAfi2JAfV80xzOAToKF40eiIbcspV/NAZzHbAfj3cD3
o+eyL/4o8ksbIiRKAaVadCZ7en6wJsXC8bRnsMr4epEOglVNEzhh++LLGYt0U8PR
HYwZFt32k8z6zv2Zbt7QPQgdoj++ey6W/IGifaOTYTGGfz+zQXfh8cADz6SGIZ1g
171dE4Fs8s4N8UFmvSwqExtJwz6234R+EqlXhlXhsKn8fm/DurmXR44BU4JhHN8S
fb0Jm+ZiYr+1ZY/1wwMyIhWvzJ1oZ7uG7rqp5r5y768nFPfwzoaBtCCA/0ExgvNb
nDmWuVm9erhvegUwzdEwCSrzKPs5Npn55EfESi/PyW2YEGaPtx40FGZVy9+LOXTA
ClWN/0zSDgivSgrK22bTQfyxP1/lwNdfibf5nLRg/hdHUtDsgrlSCUqvPIXgomUC
eY+OTvMpXJyHJ6jEdYvlz8k+5U+8Ria9drVu0IM9ULkihE0lUV5earXt8j16acEO
WHCS0t5InCsp6NXD6BzOr4ro8PmUWFybdG++qscxcYuZIa0TG5tUX9rUU0UWh/ct
MBw6+5CIyNzw0qw7BB4Pj1Bwl2lE2WF3QuV4+sTCcD+WW+4H4cVCl3UhIdjPXRKP
/cy5JMDtHq34Sov4zYTUMyrg9TgmjkLVeUVoGlLEb0/Ekku3POWS0nhmBXrmHdzB
FJal0Q3sWBuDUNxHpeabm8uXkNAgGQlmIO5pGQo5p9PT66K7h7qP4BumYMfjGtaX
B9YlztleLaDboY80WkgM+3POUbpekOSls9MTd3PCej+7/KQ3+q7b6We0EZevZpk3
zxVhDhiYuIWjprL7fILnb+1B3NFOO4mYfPZg3qmmMeMoyX8QHvVHDPh+UlNi+79L
cKDbscIfRnI1v4as9PQjbhZmXGWmkj7CO99k5LJEJTET1jqfTLIyrYiXyJPSnMfP
ThOddFui4r789Xtax5F9VLWVbIUfp41puKldT2OGnSFrMJ7ljtRukZk0PL5kbawt
smh8zTklWvjM8SW/ZNhn92PifWP5uu3tv5aC48YH/LSiEzBcEDvihBLnz1MLxxU9
0INXQmk9se8O8cmAiqs8v583rBJISuLEQUqZGu+T32d0WPXgMPMdk2eiadgETffS
THtJMc66Ye/J3XhuWxdv2o41N92vzN9JORpkauC5gAY3d7FPM8rxU2w/hILr6aR5
21iggbTJo6ebXFoDoW4yiO58McBuvPvAcu6281rITcOHBs4eSKVgQy965ioyKXSI
V5ycar26oO0PsqKDwgW+m1lOxURpgikL3nYPJ78LrQ07F7DBqvoPySPCdLXtLmXE
jSP4oC1TprdqOW14SRkGEri5PNcryh/v7wMlrdSnjyAUX1G+5YR36aWEiVK/rWBf
dDQDxHRed+IRdaXHvcoj9muVtfMSLuEdrQXbl+Tci0KS9ehh44RuBaLKkYmsWIB/
ya5yj71ish64KuKoA4eEQwnoTfQtz/y5swdqrABzz/YmouaUdsFyiOGas3qpEVHh
w9TWrGVrncs8eEE/RnxwVDNwf7Fghnmt08wefhVYXNg2wTtrr3bHlftOtVy7yote
XsANUKsELK+l+piGe50JhcTq7kbGtd+lX0TXZ21KBXzNQ6Nlh9RPalPfxI3LYdn2
7t+a7uwkpJM2c/hL3cdhr5LpAgqtEm3bKMCA2vyJIhBsJVuWjLis6D9+vEGmG5F/
SYPFZddZjjiTdDCiO0XFKHzD1XK4HaznVwWdvFisqBsbGzjiyBxHGBJpZvrAIDcj
i5/9VTFSGr9bAMMPDxtT8QAY3XKTee1Qe0tyAUsgThGr7kEpaJzISUiRKYKzn1Ju
Otof9GxVsLHlbFbUkn3LnvdNPinM/WrpFQy9NVRGEHuB662GOu3+2PE8rS/3wUfC
OLeNbQFpX8uGCEda52mkU+jSeANWYCdB0/dqySEVVGy9s6z9c4Px1MHbSyFfM9zj
QGBEMT2qlyHX+nO+JhP8h24MoPm13/nY68voUWwEaLnD/Xv/BDzD0t5EXp/sXY6d
DB8O5J9NjUVzbK3betVDypwz+VOolJFQQZGhS8bLLzh0bGxRxsbieNK+bgxdEqhZ
k3osAEEkq8wQaAqDJRH2y/vMw6rU+zVWHIFIa9TAzmy46E/ViBA/isc4mtzK2TP7
1SZ9PXz634SlOS6FniheLll/XqzXyYyNChRkULwkQ77ebf8PKQJUD5LUcQX7gxWf
atQhGdIujgzJ5FUPlly7u7q8C2AHqdx83s/lJz6oJrViHD39/E516HgQQakiSwAX
1NbedJXg+hQSuT/IEAkV84UYU9GtPiZ+9546J/Dp455Fikz/9xuuac/yqRmWKztM
peGjI/4+8SM7W7nwLOQsY9Ew3zDkjvkdN4G7K14QQ4Rd6g7ZzfDeXQniDLL69z1S
zY0CtfpINCWDZwih65qGpcAxAXBseS5/UZtwqmWoCiwT4MFyDaMiBedgo5iDjkio
vsf7BmwTV3R1MYz0/4sYRAmI+CN1/Nl4yWZyAZMUCikCWkgUJ5h+optjg0OS86cp
SldoITNXuVgIB/BxmiV10LE8mr9phwWfsf0Bejz/mLM7Noz67seAxmXFMhvb+OYY
8hLYQPKYY3Axz7d+S7P2/qBhbhE4GQ8A1JyxiD7e/S+kEzFrNBU7u+t1SLJ/eFgr
RPtWB9eMt43hfD4RJ+iHJOHHZf2vlPFBpksTz+AOoflQcUm773ahoDrE/SKFVAu0
Zr+/glme77XIRf2oXxErwz1vaqaGAxPmyG9lUXh0TozMu8VpKWw+3o2gz2Bgysx2
UxkfvSfbF2lvt5+W0BVPzZeyH6EEecMzluadOQERAtBKPuVvLn+hmJgXHLtrDxnI
wZQC2vniT7Gi/o4eYVhQEs10ZqahDioKCLAsRduLBfpA7WVGBbg94iX7XB7Jtwrf
+Sjvl+yvJwxMFwktwVnEH269jtTE2s76srNZrEw4CR6qcv03MFvgvdx2g2UzkT43
upi6+Y3hHlVeArD65wnysNWo+qff0vQA+C1FaSt/SCgs2/tS2l9fitAWN0w/4Kna
bT98eAKAajT7/O9d5Y8UV1sY4gUlcx7qlwW4DiD8wxIJ2sCpqXNsITe3PtJznGc0
1QRmfST+Z3MgKjYNtx2ngqBE92FeJqiFeB8FhhLDtW0OLEczk+d8asa1FuqIYQJ8
o23GH+pcxguwu/BK5YvpZEErbQnZAO0cxM1p3s8DX71IItsec5Pk0EXIqw6RZTDv
61rR9neO0dKiTO0q4sGNQ4L9uOQMk2SltOkIrbbG1sXm3BdzrQwZj7agjrgKPvmw
Q4s1yQQq4fjHObR6P81i7sq+KBMl4iPLvW6srYY4Gp2l3QqhcD6W71Gf7DrM1biT
vKsjlGFS95QucyuX7D0veOsLKclZ+qJmgsme0D9tDPNwAKM7Z6AzUjhVq9sGWvzv
IjPEudVuJQaAZfaYFkXyGqQWkccEf1wO5jvMc2PDtY496Cpn6ZP8xFb0YfuIc9VF
iZ8ZBn6JGlFxIKRsIXjntLmyQxUMc86P0+Yz28tY6MfsBP8MzPQjVD1wZoTrY6is
faURX6oty3f2pywPg2NPdYAeIFvWDd16qUkOVtSn4HdIYdAn0Lo3nbcSeKsXWVfk
1WPZxH3ZJdDVMj7cts9+BIg9RwfukjrrCz9Msz6EmkOPP22o0pcLyJJwn8VVOkYk
hATfEhgib+4PA1+hEgHc/t/+llRk1II7+8+6LGSbpocqk8TWcMaIBwlvbgnn3NXU
x7EGxSuPwx8b4GU0qAIqmz/GXKMBxOhw31H2x+adkcj0s3YsfPy0bg1zSx6yCTgL
ekK76QveC0h2mFyakiqMhCjpSn5BC/PNgPWQENvQJKr5YZPYjgHVanSN8fwZeVOf
2WD2urJQX6d3tRhyT+09k427ZyDJohbn4zUdKlxbDAJL71pwzzU1HH8zILSnNm8V
AoCQBAEKj5064smzSxmtyD1p/LcJjWB/HjMbtkDovZFerG/npYNUgHB0ibfszCne
IPILayrqylRCQopoLkxgUgzqLPxQF0kaAdS901q1vMyjtipTSM8K/BYjXYB87m08
Rhpcy1044T2US7ZVaNiUnWCUpTMSF2Dc9UfKF6X18SbiCMS+zAiLUZidsWZE59Dj
v2K4YOmg/eThOzCeEvl0ctMRdYI+SXCvMHW3HgU/32RRCHVZy4h94vED/XC13a05
88ELnKBeTlz1p+4rsw3fH8zCXNgaheNrAttsY2QR6PN2MR1Bt/GXzscT2FtTi8Vw
NI8KEbhUp6io0M4Tu2nGg6RITfA6cbF4g8QSutx+80QE+2nWve8MAIXZQznQ73I5
wYNcor2msBx7XRhjZjwVsRm9aLn7aNfPcCy/mq+tVCIo/EkFtJ2HJndSstovVSf4
Vl7fPftmVfPpBCGkPUfzqCix2omovD/1dVNVSKSIw7CGYOE1ij5YRbEJdDUwwcJE
5jWXp8w0ROXVtZfHDpR0I4uoAOU7p0eUd4EYFkysCIT3/13rxF8zsQQmRSfv6bKX
CoM9ZbdK4yZK8aLxg0JNFRhvubOLy6shIojyvk2hTKhVz+TmmhYRJAJxHQVSU7V4
cjMrynRGF7ZYpPQz3MmPmIMaf+Fh8+LM0uq+nMCQjZH53vy1THABi11PCDugszi6
HO1RFbPtxVdgBDDZ3qaHateolx8BQsbuDgV43v2rYzndjcUN9Bqs1TYggYph5eSM
E8QJ0SfbOlKnYritgFVshoyFLlSCg/JCaPgIdtuBu9shVyefBGtmVpANTy/3CVlS
RXP45xaZQdp+m5YNIwq/HIeRCKwkX332xx7jEOktxNV66eciCM2S+iPjsWYyL/dK
Cgjc+hXK7RpUh1NwkJOkP0C8wd58pWGtrWxScCOOyEjrlYnrSi77EMzzVN+QuUZl
t/okZnTEJ1qVawXkmSRiZ9FpFfmLENLhWFwybIk7nzc0FujseOqImCh4EZ46GDFh
FKfGlmCYv+5GJ0DPHCDDIukPqMiuc8ddAIy4/YDYJ9MCUDMTVTZQ72UAUn6yJXiw
IqUxaWde4+6q29AkeoUPZjWwy/TjbOh50sVkGp7G+HIsJSwIVe8rPR1lP+1uu1fp
5SewPSjgPx6/zZNGZNTygt9Pu1Qg8EZVBQcfAqq7mJhjr0goo8OAKlt0NTboIlgO
sKBK+VPEylArucqlhCB1IV2SOCtNdX4wrFcEpYWZqkjnwhvBubFLq4guTaNDj5No
H/XfDr2I8fkoDbtchhvObQ3gGe6Rp5Ki7u+oEIMua3rkkaEktKoaSmIn+BBaETvi
LAEV6/xAz6JrcpyICF5ePaijBzQuHETbHztwqmuKILIA6RPpWXLO1oBQ2VPncHuK
M9jel2tEGaoC7erSnLhxf9hI37qbK0gHYpSiJKtSj9/3WQ5YZqykUX4HMcO0HTGi
y9UqbfhbW1qBG5LH+4minucDJ4z/nW1pAmLy6ByuKA8KMb/dDhb8EDdlzyJAnx2R
FRNDK4u5+MRNZGyuxsNuUpdul6N6wuY5BNBP8GrnB8jMoKPAeYfE17/scaC7ygZP
kLFkowa+7sSqKBbwZuDO6q7e9D6QWnRBJUXqOsHDZh7S7N7BPTSOomxaIt/jinFQ
qkSc4exhiC4Jsk6jqjXcZjiy6eLH212A32BK9uZnh8g53/OqxzqmI1Er4VURSJie
yqzvVtqu7YxbIwzbiwGZkaJHRCu4X5V0Get6JpypTl2uMaTJCZoMCeFCyE7AvV53
r3svGxlV5UXodzqeMAZovqdzITnT+ajS7eRem1cjyxkr9EkgIipXPfJQd7xJmlSM
ARD0Rx68ajv3dPHqloNfKzW9dPFv6VzK/zDf641qcOtbpZfPYksNQ/rbTASINmr3
zbe0FpvqV6R49zFSRt8EybACaplXYABfpr/aMyfjnhyvvNkqnp2+4tUwA1SNqMC+
l5hJphKM2jMFyeCOVLz+AXjOpYpJXtrix5VIwF5nVTzAFpFBWPss4KOXzlBV3OP6
Sb0kqC6+FrN+KrD5jv15NY+95Njzcvl+I/Su09gA6T4LhC4Oj2jJIrF4QGeJlPA+
pO7ikXOjSzXmnqCWptN4QhVJutYDp0Yd2UztYIDQfqFrLubVB36Ap5HUcosIaTw2
7LsNzo1Kwp8hEve3O+U93ItYUUdKbD8wpCWM7R/EegDWCEoljbki7vVJGOHg7EJB
yqHHrDEk8ubaxoF3JNe9H9HIT2LuoaEIttygyfPyUEvbcHtflqmLD5xpQezZXDkW
Pmu+806PQCRHdWK8dK9fglQXZKvGypzSRI6taJ1KX7M3wCUlltrFfu3vbagNhoWz
YdgAdkn8Hi/+Puc0+czHPyEZh5gn7/SUqT2MKOk78B+hVowmQzlNSpbnKhsKnuQp
/QJ+J2t0iffMkkvImPC8pFHzWNYVflbY6ua72NFSOY94IffeUcTNRtppqCnFiyeb
PeIb78mCIzeYJWNW/dakHTIcQ4NAk7s8xlz3sP61JqSJGe3nJf5TPTHxMAshqP2y
5Wi2QT3cmxNuUppBo04l6yiVzSsxSYjBDXJg/+8j2aDy/PuF65SPMWTfeJ+Kg//T
KRc+oYwP6pbE3SNv1vuY4hhC9tx59lJBhPutCuw1+1T4MaZeeCzLV7o/knHt2GSb
g1B8e/eJvkdXKgOvFWY4A6F5ZPMpfOZjuwAlIigL04XKz/PmQP8vHpPUNERN/93h
k1cmszCEVr/od/2rd9dfs9lzzsQlQGB/EfZa2CLm+RgKyoC/njG4FUup0fp5KEfV
+4QpbYhfrGrZWqEQDuwlvkooEOKRNoUs187EmSG9XtO+c2qe3T/tCUbP2aQtpY8N
3PU7zFMegXAhUXbreEjczR6lSv4iYsyjV6vg75+3XqpKKvKM5lufJ0hnj4PcQ7pY
sp6uf0EQMdG3mReHebaJKLvixfnGRx1/Ki1wKAn0K5oDdy37iJJoLQWwzqOeNk4A
MLSfP+fPndB+jfAkekZBopZLRKSKKWXzW95JDFGA4ifMrys0ihr7C8DZkWJd5KP7
9DWE/8GlNziKQLs/MYVpKhI5JZxeuCJn3vvuu8X6XW6IMIK0L9to0dQgVKVcQeZK
nBf7/Gkb1A0C+P37gyJU0sSZf/iYH7AgjHNtEcm/rOF5Z43tO1Rm5NzMlr7MXyOM
kwCERQQ0/n0GPsHNm2sNVWTp3ygSiHlOReAO0EkRHNZyEiIifU4B53UG27iEUMkS
DB0ggr0VWk+Mth5Iu5mYoGHaqTpjwK+1c610fhEqt+hcP3EJbUq0K3S1wirZ/SL3
njD+gmuElGRPO7SWN5SH+pV4I/tji/aGw6odAo71PsmWrqdqBX3sxSdgvrJmPFY6
Hno6z7vZuNHeVLnaz1t5uOGCLvk+x0ageF8mC1JkYGfL8w1FuC+plMBZs6ZX2OnH
8n04t6TrocsQf0U1d5pPz2gjchqy65208CQeJFh9mu9yh2rnMRE4Duiig+mkNBwb
ag2GhhoJ4O3C8ojcI/XJLPSqFPzDcMXm05JJZItwp2QZl3lAg72SdxsjznwxqSbI
Fnr95ooMM4rFYU3qjiYy/uL9267VhIaCEGdz7OYR+BCcx45ECUVtPn8fUG5cIm22
56BdSFOmhua6YDkBL40OSIqJ3jgqMCBSRSUn+XCW2vDmg+LdJTm1g1qgf/hGX8/s
aH1Lo3NS5ZAuyKpbO75ECUqIa/OKUyrYMVPBk+vGB806AeosQEmgGRNX7Ne7VOlP
gOGXv0a8bslTU2xBleUcNqZwNA2NCL7pBg4l2/GfdMpsUfSBCzdLuonoDj0gcP7P
N+FbMkEUYWFRWmrCB/BjGbTz0+ohrqPxcNUslJ7Dm46kD3FcbATMA4h+d0oBuuvT
Zs3qn3KaNisx3LoxwFY956khiZcy0Op2TxAFwetm5kUkBlqAoCiUwBhm4dV1qWRb
w5QvvRr56FiIO7jXjc0/TjDu5hvg9VLzfcLD0a1cnQX/GLSR7foDlRMers1EzJHd
EQ/iWiYEZmQYmtZNzOpu4X2r5iv47JLwRIWyCyOT2Swl+O010hB02xotIUIbyshu
DKkp7o5uZXct2JzdCi1UBV2CdxdWjHRa1FF3DFryFFwAZOzPqbC0p4qvr/huQ53X
h1NZDskivhdlxCYFjbfTx3fgMQvQzrsEm0pGzIGLrHBz646+/T2FjxMiI+5KGduu
BGdpo5nK3gkUZp828GXSReWoD+2lsuyoptN1FUMBx8uSTT+RrGpoKla573qmidE6
+76rsJwgS4/h9NC0VT1vR+qD11EyMPpNgkkhWDykYnfM6hoHe4wEXDG0pg2yFHxf
ux1at8lkw2mp6IkYVIlknag9LoQ8wxSvjzskkl+W7922gAiiSouOSP3Seg0pck9q
+Q4Ddpfky3YkmySo7zYvZtO2hiJXzY3Ns2GH9C9IZ68BSGVWt3TohXN06lkUuDul
99BNXVYRLhok8MhYS2RgXqw1OKebDXqBWxW9iz//ftyuuzQAvqQhBfQzVwiYxB/E
+2GC23g7nvdpijIuydtVzxKHTtOIJ1gFPU1EFnliNhdLSU8tIyxiJ+Yp4oeM7JDF
It6PGLwxgL80+TnNgpzAQ3wTi+7mN6ffRTCehuctyiKIUTNhfKkSyJQVonMBqPQI
VfI8gKyXJpgPqmkR5bWlyvUqxMeb/vhOOy5MYQTzNKMj+4gtsuCYLgvjA8k+RqG1
xTPHEQ0gd5JV+au5xd2O5r8Yd8jiPi1V53PgdCh6kHl6pih94TNKQRGjwKHQJNb7
MyrMESPxWwGppyJ6z21QoE//d956ktL0bettgULk31G/DaHSOoDIPVIqKvg3tjzl
pXnDGLYHP48I7Fd0F0iZRdYCqrKkuyEIDC5Au9IJT9oW90UEVYDlFrlP8R/MYd6S
mciqJYJ15uEiVLZIJcjKtiTBvlv5yCLWz3/R37YXA6d4YaWKvnJR7KvKJCDDaFW0
L66O9vmBfHKfrm0NpjTz+4SbkMAfO5DvM0VCyRXe1pfUb5XLjh2rLSrl+PFpDrev
lJD+ofYR4lr4V+a23Hj2SZYSSYo+jAxVTFiToKiD3fD5p4Vbh/fKLQQehNp1Solf
70gqdg5jkjY8/koA2ubDUG+1SuVuUL/l7STj9A/tSZYPANPTU9LhskGWnmJP+kFi
znCs1lkf1gsgDzZ5V0vhyygIe993O/kj/2hziEz8lkCjOc2+7aBpGZ5sO2WpBYsK
+5Lb+P+jSyxalhg2/JWrLhpgIiCtoW+uVt98SvAKB6TZejddP2uZ6Cc6d/+amEJ6
YLmDyc2F4hiZ6NSguzX0Eo9Gu67KgHKYOIYT2NgMVuNmPwDkC7wGUTbYC3kCYjzI
AmOr9gx8ggAHsCMCk1matnxnP2urP3Yk/PixBxXH4ZtNKjQT3TBVGuKktBDLT13Y
BupAJxRgpOFCkUnf6d2ZClOCJBbEsHp5u9+INNRaLJXXBUjR01durwgy1CTWhpAS
oKrJyExEanib6/3rrhboNAB0VEkKBl4FVlpR7m2vZ3MMKwi0PJiDXAJng0VTNHT6
+LByUCOeEjskGxZHmjobsi8NSeDQAjWcDU/JGBiecUuphZX09SzzB4E0U5sOiUiK
HOTdJNtQRrc40mcbPsV9naw6B4AFBelctZdYl3UynOZqi1KYcE0uHBc3OxawinQQ
OxCMi5vNB8SnQGnMVxxEI6D155Qa9sNOBZlmZGV+vDb31KceGTsFaK137QzBUALk
N+4kor3Lf/3t6ACV9qBZhp1KocYo80/hf6N7TZRcvdyX5P6XBzCokkUtVFjW7WgN
T0Sgq7E9RnxHaMhhELRlLBAPY45Az9PcRAe10kEmVn8ipX8p1nJlCt08I/+WuImq
VUpLmVy5z/E3sRBjula+BFqeBrrN2msqNEqAr76thJ8qDN08coCmHqqKn+EganvA
QCIz/KuAzFgeFDucSi7zpNxTd/SewX7H0rFsweCljAPIlYfe3x7rOowf9UXLHyBK
uQSIDAONIeUqtt4nH2w6MpGubSHZRFdxsSu720Y7Wq6L+nYx8Q2GDs9legpnGezQ
G+1w3DqZfrUa2ctFSgUJGFW/4KyvBmpIYiBtF60piquMHAIDVGKqqoIeuZ06/fiJ
Z19CejN+zJHG4MwSdkt1X8NUSDeQobryzX0Z+uty871cVzFzxEX3v3haHEBP66SB
wx8/utwL6qXSed1RM15CcuUwoLZE8gbPORiglF9g8LVd4duEgu01xYnYRrziOjeL
wOnKCPVqium0K9kErju4+So9Rk19+dNtDP31iyOWipk6Q9Mdzdj/ebDCj6h4+iC6
SinA44X6WCpCY7koD6DnxGTsUgnqtdZfEi3BXmT2zYn1JgbbjYeAj8OrsltmUvvA
hnrYyjCF6j2AaFZUL4gEMlAKCuRACh+vJKrR9lcC94RWgQMv5ceCdw6zH2htOjEY
Jo+Euy70PUHtSy17Jcd9A3lP1wUxGXpI1iGosm7RZ27nEYrq56k8hWCUmtHBizgc
nZbP2LnmKChX8I6V7991+T13Fp03Rn4c5KDsoRqtkVNfplaoWquiGTS9CnlrN2H1
fEnnll1yQqSwgueNzP7/ekrBXAYEnB7IA5I0RriA7x4LSykh9+lBTa/09mom3sB7
cI9CngrzxnCG2YZLW2vlinqno9W4D09tNy7cAQvC/Ai2Lq24Ruq50Tm/mxMgh+n5
wPbZyxMpMfmNV477PGEgeetKHF+r2eQqvtxkHZs+c/LBPXnOZUkX00Tn5D8BmfHH
1xQjJ2Az/6r78SWhgap7fZR0ltELWk5O18Yw4I5gvyn4QpHR8rjQ43+tQcWW/wgS
MNqVmUvy2TteLxio/44eobmOLNIRuMbWbYRtCM6mI44GFWkKK0OoO4ItLtTc1DSK
YSNQF6xcgQJ0rK0ieQjs2IfCcRISU4VMRJ7nC1mrJaks/rzZ+In5X4Lc0QrW92hI
UoE0pfq/nD6WdtuQAkPB/vyc4vZ1lpM37c8bY7N/qtd6tUXLu6ZsUi7iMcGTiL3T
uG2gRUm8L0mJt+E2PvKQ+lsHmEE/EMTA8viXNL+njKhsl1W6gfUZnGibMXcN1g6r
uxXchQc7jRSyLXHiQN7MNQVe2/s3aMdaGefc44WaUwrgq7XgU+3r5uUOlaxuZaTf
tdP/4gDdX7bq+r7RGMxO09okTvYhPIlfaNGJPIhJpoozfPVGn0u3GhJuunS6y3kH
g/GXAcAfSgNxhX6kc/zO7p2YacnIIXlmrR/mzAeI4wtXEBsv73WxJTCwBEYP0IN4
woNCkNU2trn3FAXtDNpbgyFexAjdKw5ujTgKtCo/yTxEQPMkuZnW22kz4VIQZF4G
vwFOm0A5t1ZRJwy1SShmUOvrZPYX8xSWgxNiGzM2eGtWaqChoeGS2ebTyD/9kUpp
I1197G9KxwddueyueN4kNwDee4ZUuKoXaY6+wjugGqUUz6gyiZwaBtxQTpamNYjk
DMUa5+4j7E5+9zPYQU0XO2y5JYnfktVMdmrQwIYZ8Pa5gC/7Br/1QaCiWQaGhDDa
nvcRlMhQOy2A8vhGqNfBrYcBS75SI6o5XMNqVX8oOjRwqMiKXsnFl0KLlKDc2xMd
cEDr1nCdSGhbnSehV+ZiiIv3G4zgtkYQDVkk7wHPTBz5FY2WK53FwCbQchLOlTLB
NBGZyn9AUNhkCoPaSOfeVjarfAozLkwHZqVX297w0M2q41UWKuBI9fxhbZF6IIWD
67M1z0BdC3MHGrX6E3SgqTZmQkAT1iVYibxKpkHG8rhEfc2Mqn0buEP7VoDf3QuT
5/D7tO24ga4iFNiZP2OCwentsFgG50SeU+lr2VelGDaymK0O39+jpjgmNovIQtNW
G2ogBcIZxnJ/68TTYKAhkQeOZ8HT0lx62r4+m31H/t+N7JXNzf4iqyDiHoBnFDaE
Rmtlu18vtcH8XrxPdvBOXa0iBVkSiX3rT/dMHnhW6JoXmlaZM+4e6T7IP/eYosp+
WoC7fj7XDyu/GL+ua3Ps1yISQpw5heuzh2Zg87hwW9a6dDOfJzG8uB++90hDJVjJ
woEWn4+yiqqFVRXMp/K/x3EZgOawRJoAumMghe3fd06KB0wSpMn04+gyFVifzyRk
sxN2R41Vbp7qIKtSnwtUF/wJwCZP9AHdMQY43qXvO8xmsuSCzHsF+HrrAozZh8SS
uLNkJkI4RUNBERuuflZu2p8LlFPgi7PAYcAMeMBROWmZzFep5qE/szF2uyNrv/ns
DlbEcPiLUaVdjY6apG45//3p/cXjE1gNT9xeS175M5/BcFFk16inEHXlPdtowsJ5
8eGD9KK72yIQHXo5LuabXd1+jtG9SftnQ//+SSSxuIjG3315JtMuAfPYg6lYf6oJ
RRth2HOy46UOsnZ2aH8bxrgPwX7h4PvQrkPIHhUWli02UgT7UvhNo8tb627Q1duy
dwKyMn7dwksIuqEaG4F+8al4yRT43j6R76F3KO7KrjekABrsd5w4OhWCAaFn4So9
kBSiEmf7Dc025Na9ztvL4v65gMOGAJJ9ZV0Bj6cYIuhKc+MmjEn3bWvA30DunV3U
esWUAYUAk63AGlGZhGNzMaaNh3tS5jJ9tCK/0dyTnveNMNuzKbCMQS0Mupe+NBaQ
c2lSeuPZpcTUib1aELdVKDekWSRBGhpmAVGNBquVQ46QKfrfIKQTCvaHyDiYGyKY
ZD8sJNb4yn7wVBjXibQ+2s0IUGq4Zc8bBhdw7+v2HykSj8uzFyoJXXpoRE1Ob2M6
NrZwWExeiWMAm2xfE0SNMMuZxMkHciBc+1psYKX95xKB63sirFJ9/haOXOMUNXZS
NocjoyyahDXfOCNojXACRzKSxchUIEDXdZ0p2PK+JHPR2BDXIEeZhqXhflHJXdO1
yLUN6zVFMfG+QjSH1/aXgvHzt6Md0FVefRiHj5DGRViCQya2nMuNzQHcT8luLP2p
SySvIa9yUa7sgSiwLWXKVY3wkeqOoSeih9TTBmAHGdW1yW5Yjjo8BfJDhF7xQWGl
csnwB92hjZov64Kna9KdYQWR8aRHCHIRUBDnUDeMh9w1FitGslvmDngH6Zyklf/Q
bFTezx4Wmygi93ElZxb7Ft2FW70SiisSn8G0Vy6js+SN2nI1eHaapxp+q4du92PW
krYYFFSPJbD4IbfwlLr8BvhDjJuFld6sgN0CyGVdITaOSWdMmo/6FSJ4ANW6LuV1
bCEoewxFvmofF/VxLljGp4SIwh4IDdsoGtX9A2BmWVfpwBq//msx9TN51n8AawR1
ufQ0L+KEjjcgEs5YynF8x7Rt4X692dQ7KHVeUp8U/vOjYvYIO0AcUxTamQV4CN7H
bF07ig9KKyIT2yibQJ8w/HCwcZwiMlCVXGpIhYBlnx5dKpxnonmRuAOk+9a0yLsx
Nn3kclSMbyiL8ADeXZLdzjvFWmM5jBR5YqlvEZdIOs29gKs7Rppu3Sye1BFjcMeB
3j5JsHCRY+piIUnpuq/MqD/RXr/TdmXXRSxgxItlyuWrIFv6tnjrWqoOMdh7RDK8
eU3zWiE/TAtNFNOZpDSsQ5bxFY4ry8xXgNPOv8gDzgwdT04JTx8cLKMnT90g4Kj7
DE2z+u1FB/2fQenugLxJaDNAsl0ZsNXFCIGXIFiBfrvVS+hVlFarVqB1fV7UyIbP
DJb9qxvP/0tdZPWvyL8Xb/bowfsP6EEOCp+dA7Z2NXcSMT8MTXB4LEzsMEcFyCIo
+bnxUGRXfuveUq9FbtTaP0IkewkEcmvGU+CfiI21x+hqvWdFRy6104+pWW0jkseQ
vLajxHnUYgk0iJtesrHenKpoKQ1MyLT2GWLtuSM/kJZu59D2NA3mAv1QYOmeFuKe
r7Sg86vwP+fmFZU0F2mZDfs0DW6UBu3yY3JgCzN97f1/yjc67r6w6lvainYeaWA9
9yOV/qXzrDUnHOKRkyOW7Qjud4PcXIqYzZ46j5w4l4fj8P3RHyXy7+V26o0nWBz9
4qeIrzzs/ixgN2+c9z4uq0FkPMU53m8nEQoW8QxNhI54drtrnZhUv2iG8aMVMfQ8
6iKMSRx0q4Jqh0aypUkNtLG4RG+K6wwXebejhJ1s1y6jlgln6jzsCErV+A8N3cvb
2tHBc6isYdZcvFIczimGne7WD0k3vp9GideWdZblIWPL0a9R6DZkZdeFA5fG/Nia
Jtgjp8GH1qRUHQ1INMNrkD54RLPBub+VlLeJL+Hfe3du6fh3enNmvCYp/1X83BLF
34NuJ5obfftloTon7mPufwMO5dTBdzJgFm2chXcS9r+Gkb8HccIYY1wbTBm/LMJf
ZAMlWSlZP7fg9lsAAP0n+oi6SJ034OE+s6AXe+PhE18aWQzEzSUBTeBOB3ZNBvyZ
U6C3T9vN4j2Nb+KkZ5mpneByXJKW36PNB4oG9V2yPaQFUsxpgymSJi9pTR7ykBNn
kyjZGB1FgrqQnk39tW/AWxRYrVnn50AkUC0oZoCPo+vRwkuwE+G/soMrGmBiOi/v
6C7QkoiTPAINrA7HD+TZ/sFoA011eqlrlDHNZPfrVw8V1We7Gw2qeIKedcwMdtzI
ja28J389dKkPxVNQ5g2kkuAZGSW8mBxpI2YOaGZCU3tUqrvZMG8a6KxD7O6bnTca
ClRne251B455kSpwK64mQCD1ObFUMeiqe/p7h8vCroDHbKytn5A9A7IJMwEx+Ipx
cse2kvC8WvYq0D87efEdJOK6tHYeaS0st0uPb3pZtFxzW8zceAweJ3aKjf+gkakD
Da7UPLERtZNHCfC9DvNURt8FZZ6mGpWmZZikK9RH9vXDvgdqZ8CGFoUoeYYgDTiy
3ISKffYvEpDyRvEr2I/ssp+aZAPdM8N1SE+FIJBs+JkunRGzJXgF9ZbJWXTSRAuG
gZdTYpM4bIkiNYI+H4XXcGm+xT1VXiq0FCSYDDKrH4NgcfMyTkXvhEhp04qbw0Rw
FA7cRRTrbKvdGS03Al/pcuVvPNB/iU1qv6f9QuMxJIwg6w/IcIwQJ7O5ge2HQetR
8Z12oYZI1KwRQCljlz9/W2haGY70CQjl/I7hIzjGUYRHFtCLaB3FDxR+x2IQ38J/
p94g4qqiy2eiFYBQ/cG4v5FjJ/sgOzS6HrCND6qXgo5p9Do58oWSbzANKADLb2gV
/E3tV3cz/7HXh9gcp3MiDK9SsoJy50CVvX3wkl8jPk2GTg8wW7LpYlxsZ3gcWJVF
JveZg8OpikdMzdoDgsouDpKVtcAfdG4JADo4zptNDDll8LmGasz5h2cjekvIVnF2
+9jCAWUOHQoZAd85T5nOngiPrafaKImE3VbLqcOmuJjywP8yMlKeK+d8c382pGed
FpOlorfg/2oKwUtph9cOabYr/gfxMGxdfBWy+3fQhW15zfq6sCjOdWudsav4XL2G
qvV5W6kGRxjKsScYIqxzc9G2uQ4p4ea3yE7/xfywdvAnnfAA+wDJja1u9HZ4340S
mTNIsYbgqCZYbnFLTcnQxc+DO/L2r1rCm8iq9vkjztIuzpU+L68fyyDgtfzVXtAt
EBdjExQ0miwasMnxiOVA+tbqnob7ZYS21//1s0Yf3Uwp/DXvu6lBh2jC42EmXuAg
NFGYdG14UISNpqGBgH/fvzUP390X40Uphg3qPoegvwP/LucRV5qH0EqToM5xofvg
Ne8OI3xe7CLF+CyvH1X0CJtDL2MVQuBRBTvRmRE99L1XWEPYqg5VQbHnDC7aopE0
VMJDo10X2ZXlTIIsDlqidftVP71auadDliORbPxv0YslIse5aktriZsec7uwSQAG
42d+QJu7Lgqfq7xyJ5XvmSNI+/U6qwSniirw/Xe3NNpQL3VYdA5j6TNJix7Tlyop
xcyN7VS9nPJ74bdISBi/SGj83Cc6A6CfCQDD+fC/DMl5GZSevVSQBlmAzMw64vR0
M6H4Fzjo1DwEk4aFZ+FIUBK3doYX2Hu069SR2bCck5UxUh5Ky08ETz3JRpyopXiA
NMNqj3C+4XCUtj+ksbA52a9f42/X2xKFQvrYbv1H+NJgZ9s+n5E7/DQU7TEyXuoZ
jV1JD3CLYBZiXbEYaUd/QCpTg51yJEd23d/Ly9eZHNfPF3mIsgBi1o3gUVgDpPFX
0J4OCPe8nVsIbDG72np1uUReECL13RqTftObZtKHhYAybf7iN64Ged3dKbz0sDE6
X59kBWBVIgjdRuH6a+1a2hKZT3qHQ6rU33edguvkEvrCOCBAH+kbOYk8wMwgjhZF
DCKXKZCrl3TOHnut33IVmsNC803jap9eV6vwXyOVHhupiBBLXiNhPsGPSyWnRhSH
J2loBjbHz8jWnhmidyjNECJp+g3o3IXkfvHsWgA73T/SmCNUaoEdOlQqb2pMLKPs
QT2Uzp6VBJGgShFcE6IGeiHiPynjtWdKG4DEmAgCG0FZKisshYgcrouYYr9tdB99
pxQYXIt2cmapdD2jrsxo4CDuU5Che7wAlHHQbm1JdkptM4Wzg7z6cvWPHKrKePxH
ehStYefyTJhE65oushQ7aIbngyE4M3VRQjuyey7BpMlLIfv3O8sOKiuP8dae0HXj
CmnC/PkAEq4nAd86LjyStkkHUTSRTOizJVT52gHfBMuM77jKNVBYgQUFIoobikj8
2Jyo2nlmHtY568k0elL7U/bpuuS/Pok7O28NHiZFmHXTNaBOxFPSzQiobp3/sSv4
HqDqjFBGhWlDf3e2ruKLlo5JtkhZmkxage1XgeF8he7N2QX87WV0z0KiubDuhl4b
dkZKqN7dCAFghA4NePR1nYkzTiQR7KQMJD8u9Vww7UK5kTu9SikaGZbtMRTnbewo
vMs12CyquqtyL7cpfAB5PaGtqi9pxAy8eZkWrsb36POa/g+oKxUyRXfwyVd17G9R
Xt7FuHcQg+1F3bxsHCSP6huOo7einZ008ILcO82a3Tb16QSmVSHoys8YWm+wvRPI
h5y409iGaNJVXWewWBcepYsVDawiH9bBZOqt60vbVy42qvAOMudGAQLL8enx1QZT
GoSZY1+gSh4vjYSDMbUpivuQdfmPCMqkUmh4819YmCAxXUS4I6pe8aOn/l6+KJu3
CEZYLslqwo/d84iuWVCxnJmi6bBNgeHxtiD4RPFhBex1C6Klajn2e5i66ViV+27x
XvQM2M1gwmh3RhzDWyzqYg8GNn0raMLo0wqJRtIYv4duM2yKCNiJGXQVx7WZoNyZ
83ckltt6iP+Y7K7gaul+WEM6XA1Qu9UdB9VfqoG3R3TSwE8ipasXo1Wrsd4Rv8Us
HX+rXfAZlUHg3MhUz9iOmUI842CuYBd+9Z/NpSYLjSCJr6vawW5omc6mk/MjsCIO
wUDQwyNl8uSb/axQDQcyOMH/lnzJXDnlbIQNQ/9xRzDDJTzTZP164H3G2pPYwDVj
mcQ73N1wqAE5zzj52HNtkj5JwL5jzugoWVpllQX3kOdktig34s0K613ufVF7ZR3+
Ju4rUW3kOdHaNtzBENbZI6DSsm2CE2pkvJaCGQ64keIbfvWQ1HYGXxLChjtaql2n
oOlrosK9OXZFNPA3NCS8DnyKV++upTsOm0mcINxbGZTKi3wCDV811reoVzsJDMe7
YTnuwksqp4y3fdAplUTxG88K5uVcJwDlzWycE+kAq913c2VAjajFiV1L09gMh6eU
uojf5FxTp3SYM/b4XC61n0ZarMU+sE8IDzYZciCJFzlw0CK0rErEH7dG+TwXAoVF
5SbnOZtjePpkrg89nwH+xVbtvXyFiVFA98hUwFBOYkOgbTFLcDo5M5oTCutxG7+X
8fo448ysOGDjNjW72018SOMpCd36kBotj635wFyK+Dv9kAMutvwi1OV4xdAKa7rm
Q324m40q684PENrXeR2dXjKDGYwiYY4o/DffInA5uTpCDTSwbsYPiokcsyxAYJ4T
/5gtt+ceTvLiXHIFTpyW86bqDbGIdIWTDPCXC/xtLcjxl52pKbL6B9jC8Np8duw+
VOxUqsm0yqTsbz9e9FDJcrZP15Icct09GpKuUiiEvZ1RNGbV/0XdvVntkJ8uk31Y
mb/m9HJWqBJn+eyIU/SEbQBI9rZPljMPCa0gdFEvCYD/AAEQZlZwVm2Ls6EZMrXN
P8jFpRfyVIbDdkOmWgW4xSUErz4kP7Meix4TD6xnhv5JUVPlZ8AqLZlqwNte4Q5i
fmm5pmgA+/cHaTA4QR1u/uwtKQBzOwU+ReVB2r3e+0tr9A27aeAiFEq4/XvUmH9Q
qJaT6vv4FONfM5GEEV1zZAv+VUv+Ckm+GxU5ZRhT7xb4Alb9Y8tn57SS2fu7bdRw
IZvWqAAiQXBpRU0CvI3zXPdSSERRiFH3O3OBgvCztjMvdNDRpBn81GQQhU3kjzi8
O6+HGNRgK/peYFxonvB/IXKBXU/tENwcxp87tmpyFDgBnBa1zcdqmbqyppCzZSsO
p8ZA03a6vHQTxzluWDc1NYPQmt4QZesudKYNpd+DkQH62iNm+O5COZ+C+ga8Onfx
pj0O/N3AzduJjq1UeAE2/ZsMRsT9yMO7H6plYkgFZW7XkNRfnjLyIfDw3RRdodYL
P9Py7PcVC1gorsyYvMRY8XX4d8ZNdJRdAUcP1/SCOtv+qLjCa4Xl3s+qhYkv4oZA
RS3s9XZNU8ap9mYC1vXUDnBita79x+6qW7DOmdMKxXYRgSIo21ELwxTk/MpujVdC
zdA/2UDNC2VMPVTco3vX/isZyxVeE0FlhcGUHqnJuwrgnmvZ0/moDjOzgGE22VDt
5VxWOvmvku5SgThaHpei0GvDI7FJ5zqbJUc4Hs2w54K1YShGq0GHC6dYYtPJO9Il
UAln/F5Gd3eL9uPOFFUGzYT2tx6bVLauUrAQt8cAO/7iLMoGxnrIUmC+NCZhJn3e
KemJDQk+mQN+shvpyl7fYdsBQ25q2kmGOrwY9ar1GeI16wQyTsh5goDJLxNH9/jl
P5Ok7mW/a9JH+PUAUdp+QcA0go1m/plIWsvuHTbwltXt553fZxqtWwZTdhUoxKS4
9filZIevMD7dO0LulTMADFuoiv92/0v4D4o+KVo5y3unrKbxMub6pQ4JM3VQMoFj
safvvnlF3wCzJbMbtEtvtadcOi+ul8qkHGEu/N4aG5RJjg9v8w2po7VBYFGvorm5
X7KkBRIvmXRul8RMNvnsI1+WODtqUm1EkenxUMV5k//oRjBH0dVrrHNI2fmF/euL
4kQdSo9w4EVeZn0Xsb3LmuiXE0AjjKFT08AboO+d3SAXTvWnlFTha0Ar9K2z6xbp
Qs43suW+ZPzjhZmCcMjmqo4IyJrhcLvqQk1Q8k6soCgGsb4HvlC+m5HtyQ+33eWp
jSA1Owxcnta3iegLjmLtQ2/jSDtuLOfpx9Y4Qn6mkmRj55DpF+WHI1/AosIp6XqH
D/anLn1O2dDr7wlfn2ZcJ6uGTp3fm40ESOcDYp6EsAGqHNRMXljmGkIXG/rdMv6J
9o98M9dDtUsgKBhol0lgrBh8HrbCJ938zrERRKVFSN/pvhalbNxWGdJuUSagLyVz
nTpfBAikrm+SUYregHBU4jAOkNGT2/MgqBfCP96WN6XRPzEvPYDQRfN04oie3jYE
svt2zhXUvS7GpX56+fFPKotNjqkj7AF4rB9nL+zKMP+MmbM6ylum6rmNL36mAAvk
FrklVXJ6mk31UtF5FcXA/DVlXy/DE1DKEC2dAxs/FRI8ZrecXFLwRsEuGPs0Y4rQ
F6KxmFjMVZ1QBaYuT8HUuCXYwy1VqbCanfJ6FwjuL3MOgQx4jImrsVnAmbKNHufr
ljMzaPCdBrqg+IXUmloS5/9TqiusdlIXn86xii4O9ag3qdfZJVYs7G3gwdlp+Yis
AuWdyoJpFdC323ufKh8c1CVBu5GHsKd2sDY6gu/GKzf2dTIOH+6t56dxJJGMdlpJ
rov3+YJB0arphdTq7JuKmk8lrxDaVfQjjfFjl2ClRR8/2KOBcoaetG9jG6L98omK
MH8GuEWalCcSBeQZynISAHSxyk37HwEWlzYADJsM5jJKWu5853V6Uye51+ddlU7a
EBlhKFj/G1VYM1TYu/vC2eH2sDSkVGm45s19q+i/LNSHLcJxR8CmPfQJBDpJsWpJ
sup+M2iGwRpZ3jCfAZSGalFJAPPwsufVu2xj95gPYbiggKA+QMczViKt36CJuU69
acVx4eaIzd1DlRHAxZ7oaYMFpH6hZAK9wQWeIrctBQxsXVhkf8GCDRZL57cprtq4
0agayLspzqqrmoXz0S58C5KGlSIKnwcXFoHcLNcGVsPjAtke02/36k4MNaTBtxrm
fDKTuiqCg1KaKuZFtgpVZas4t9sOfaTOx8NCRegpa7GPx12w7x4r7g55WChjY+Gn
Ydp7YZ19gbYpBLqsaFpw2OleBz/p9UT+Tr3WbjylOOGq4wmIH9b+8IJjO/gnuJlK
ghCEaiGehOoJQ1lKvd0YQz4G83zFlS5cyw5hXUwHnmelHaJ5b9nKVj5vJX7A1yGR
1oR5+G7GQBF9o3fYvNi0se8EAzblk8wFbekUOUMkRfNkvER/O+F1nK/kmm4RBDEF
gpec0rV4F7FqxN05eHqyOQ/9KlQvO0iRB3avTNdus7PAgDCXbLE0+PPqdBjthMgf
QvwKn2t31H/9d9xdItiJ+HKwC/qyg9wocwuxEdtGU2wNKG7O1HtK+yryYUUkH9pS
TDw4X8tcQr2hzPnZc+sO9sVHolTkPlIiK+nLuzdvWIREtttXyB5PutpM/kUbT6Fa
14Ys7mN0QmY5cxH3MhXeaLV2qHxkDiW0bncfnVhZmkZEM3VLI2oj8bk7CemZ85De
4mmNqzaAqTLtjRxpitMAV/vMx84CG59Gy84rzN/ljDFKZQeSmoS1cUu24ZDSpOJd
pOYDlY+dwPPzrJRHlSAasLdc4MogGK7i6QBNyWl95pPxgnnZ9q58y+BGedEzTOpa
y+eDp51FO8boy8k2wKLVBgt7wpVIqDfcWfTRhdyYYlIwnuoYTYf77traZ0tquwQT
2YVsFJah43A0wbtmfZcwGLBZqOdwPISCB8MkoY6to02dywcMAvPDuU7P6gMrgZ9z
+Q5iKt0XAvim1mtdqWtG+NL50Hb9lFumLyFsBgn/7OdkgaXNS1QJai0tEVy0/L0g
xaa4e3VNsEgdgz1mZKyjemznPtYe3xHDDyudW3CH0lO0O8pSznZHkkk6ZqA8PYfX
HW0EQB827McK33qpFQXBtDy/I+8qypiYsRU2J8DxnsgubEVH/7z9wxVsJb0wZDxT
bJdx3YpBVJXv1nM6DftAHFs7ADPh+67+31IU8W1jpUOqICzysr/3xe+rixq1uS07
tgws9Ig2vBa97StjtmVBsBGSf/yczWOVW2vUCjqFeFqGI7KlxSUMkzImTGAyIWnx
cN+fLbvlzidC+Uvb6rz67//gioH9R77LouH8a1usQVD53hf3Rvapx7GfBDisluXL
MOlT5LDLTPa14imvIjM7U8fMEHq2Rrm1AmfBqA+ncBceR8goo21mJJRHRkIhZxod
886nRu9ksrQmw2L0mzJRvl9Lwzw5m+YeJ7fvth9ZNvdt8OdK3hRBtI6K4LXuQoi4
FZZPe2cIDj4GAMACRaiS+t32Fu5wfmXrUXm/z/Squ103QAyctpDdcfn3O2c6eUTI
PQ5yPayfGGllAXrlPhnhqXVTW0qn889GpOEa63VsxGoWzt8eqXOfHVWg51CLj60z
rOOqSCCtu4mcl7vC2ec0GRCUzwFjMu/+aRAGJdtyUn42VzA6/59UwdDG+7NhjI9J
6nboAmvLXC7CSyGh4zZzsbg4uAT4CiLNdWgsG1Nqh9vfObGCIMA9t3ugnp/Sln2a
d94t+dcU7VZ1Xszc6q7jp49wKQ2yTnsoK/A2/0os8V8oQ41DwVdUMcPb6ELiiy9O
Stt5RKlsn9LlaC1fs2rFbYR9+aYUYsuia0DYc+1m+s9227FqD2BvF/lK8YJeglvs
Z4gOejJcRgGPD/r78kYKaiNb4ftym0yZZieIFI+RkiHRvbT51sZQRHjInCVjFRt/
2TvCMbGNUX6K9goVVE4e/uxOadoSe8i0JHRM60+I8rI5jS71PTVVbOtH5bfWZ2Qu
pKWm/Kg/HFxE7v+nxraUqFIzjgWtFDyyKeojSpmXnwdwvEajWDcfrEyp5a9Yt0/8
LiEDb7FZ8r4076hirEZobktBWfuOkUeHvgM1g5Z2HQxQZCm8FyNc1e/0HfkMZz+S
IvwbAYtitRYzim04ntdLyrDsB7nrQQpnxmSMfXyukZ6p6YPWbkakCWq0x8pYRe4K
/7sqOxRZ2DXF7cplFc7RbVyobuPPCMTrvoqO+LAP+ScvoiMhGBDBiDqEQny36Gm9
`protect END_PROTECTED
