`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KdXZbPGS1taifuI7dAnhooL8zvcD03M9RVHJ2BRaJAjTUZZoobe/f3+NDeTF2hzT
n/7EEHgiCK9eYYUs6lNMjmq286jAwD3zN+i+Bc9ut1ZHObeyZ8b+C29H8ESgUcwb
Js32waxkQ6IAAPBOv8yVQ66VTyLPVvLk3MPNerwDpkJaUwvoEeMyvZ/atsJ/pQgZ
QxY7sniR/MzAuifS4naRgVkqXdTgkwQ2JWVu1+Siy4Cph7evUzwuGfIYuTZIJZOY
lizE24w053UHBa4KAJGnvuF3uIZRuAy6MfUC4iSUb4KSU0MOAzlnQpeMQ6RDLSLw
JjkwcObO/Opb9x21VPqIhLysuiObq4GdfnO7f3XNVydE7EV1wwyBXC5n0+QZk9+B
Iloah7kczBFaBoDF8rKT31ATBott08OgYFZqT+32i6jT6BvgRnQLS12W/XagI7RI
eJjdm9hnRTqepQwai3nFDmVCrlCUyQ6shLqvfvP5GQnruEWrlURJB1E8g5C9VZhw
OpG2qDi6JCe1yKffUB3B8NBj4ExaMXb6PNVFqd50cniCIgHLxux7cveJmE1baJXj
0vpk/DiObZPHJ4730MX+Wy7peh+/6t5AtyMJaxhoiPrnArbTMcJXhl4okJiKt2B1
4kF58NEkJdtokqlQ6UmFeOF4la1bbK/NnFZj3/H9V0lEs0V77OzfhnmZjx4FPTkM
jGIhB59i/nJZX8n84AQsN7NTTL+OGMBtjWnTmyHz5vGLwq3CfSj/1CzZqcRlaSDd
79fbh5hhpjcMTkFMCxJO3FJJ1xjlDamWQEPJYm89UVH19m6Qs0W5qMwwH7vk6/Dz
Oe4dUOifUB20SSvnStSMTcInsBEmkBfs3nCneENWdD6V8g9ZiNuxhcJVG7hu7wbL
gdXw2yz8BTV7PMiSSCsOoT81OFGIBrK6SvUwKFUHi35QxkQrVXj9N93SZY2JLaPb
Ty94EqvUTm8NiyAmc4AJaNG3iIg7N9YGiW2s+jssar9Uea8oF5o+j59Yt/vG/+Ku
EbQBxseB1auAb/dEmPltfsBa0PsMYR402sMacOQwBTNr/FXvxVRfH7fMa8HZoS+O
5IwhmNmaxYFZ4wHEYwsH/EcBYOHUX62qF+IP90ZbvolshmdMsgNRVSNfBvlPchIQ
0Et+6UaZaT6+EP41ziIKU6CLlCMRBpIsM2S0OtwMdkC+vwhRoONDdZ4pbf9pVXZa
Ws+vApQr71dmNUcjwemFSg7AK3WaAFggj2vukJ+M1UJLm0HfdISalP/5daMw636X
WQUzl+anQgbN5VluJlDdid+vSjTVR6N/kleE5iR18xYBxqzcYlAPxv09//9ejxb2
vTne1C4+ok68FogHjnXkyxDlurjWN4gEfzk6obgCRVsMGXYK0f/ijx2f2clHGVKQ
NcOcPDYN5sLNDnysrR6XrhTIZmwqIR731K23rTOCR/FDDQcy7YTWJClAjbS1xRqs
Wk8AF1v4WyD3NdUy5pUcA+rgoggcfMJJ0U1ccLzK6H1UDrxdFvhTo75YDLBdn0aZ
mDR3EHM4YUXU3L1qlSOhVwJusyEOry3kpFoHeZ3RqupUSJHDS+HBfjhvhEnuaAN2
kxzgqXnS3aOspPnDklw5vTzjrSzypT/JJ8MSJdvDqxY6+KJ4raZYnR3eoUPE75m6
07kF8Ne2krW249B+2BY1mC3of+hraxLexIWk+npkYgQq/VwBjY/aVDlvVWmj6HCI
XvDhflbBWjh+KnopUZn+J5mOrwPLm92ZN+l7aCHQpnHH86R2002/dKYgvyrtgczc
ZGAfc7+JqbciwEN59tpIESWZim85AQc+OeTayzp74iwJ0gsHOWjmrGQ0VoIjEAmG
ZP2ULsKtvLEa8QW/gVdT/OSHROJ670OG/9COhL3lQQRRbVRcSCD3ItIVpuR0fWnd
pSNhNxVyBsaRIgNSK52I9OuO3rvPr5XqiYPGyTJsnrqy53rkcALyVVLwE1rdfL8L
thjnXmXO/XCaOVLHiNPoq0txc4vzXIJh1tCXs34ZlnHW2kzyfiwwcU+4l+9rh8pU
B/PuQOMZliekv+Sal2Ge1+SNBrzs4e8te+zQyt/4y2eWOX3vcARX4gNH7LY3RZZG
zCGBeyKjKGJEGu0D2CgA8e4OOwYAAMrtzUeLBch99gc1OaWSM3lEvlO6qTjguv32
a1eLWyFor5Qi161zjtDy3dsKaUvV9kFDqpAM7Ymaiow6o+GqyVq1xJNT4MBCxHpR
VUBVOgZY0dS268spbc99Z9rQX64d3ymzV+JiF2VuGVPmnWgcUg/2cNB8dEvelOoQ
zj1xTv0N8dRiUsXsMMPhRoPBcl1YT0VF+1v18v5UOxsCUPzIc7rDvI1PQobjvcan
b0Zjwl/QzlXfg9/hynae4ePhUSaAXOFVl2jZEXPR2EEH1DSyYM/WAlMsLq1THqSC
kvqtEoWoNNhLTFU8298xd8hN476M6k6ufyk3KSSv/hRoCdBBoAO4lta0nLCht/Be
38EREZOhRhAUvWonlcoUd1ysWrUUICi7b/YV9mAFHdpuzBK3hLut2tuy/X3avFug
g0ZqSNi9fhvnKy7vrgqTFwxdwCwunAUEDPK/BBia2fkSxX3QckUlWjD86lgZkoXR
v47yxiivrvENNWCt7nVjEZ/x/s1g5mcvSAgW1LIXCX0=
`protect END_PROTECTED
