`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFqrv+dh9GN6tn0UW9FZvCW6m8S73dDGtUaPTco/f5Jrn5QVysRR/e87Gpk/5aqw
c/TidY8MPEI6qoSBrA/Xo/Z1VXa08aTfqmXm6eNvNoWKC1abIcrSQ5W4lE1Skt8K
l+91M28vx7TOkGsNS02c123nZwdSpgGJAD6KTyOY3uq1SIvxSqt1FhayrxZEw6pq
FFr+2MVVbhDirG4IHxo6W5G0jVPYAu9tIiBnCu/cz1RfMihzO2tWpBro18B+f1wn
Jh2iR0Pz9dI/IDAK+HyQgEUdaPqRhlnEyyghmDWlyDe7OEuF1QQJR8wQwnIdliR2
lj/3dG1+jD3E3YZ14xOJ5dRGaPvqEiyTfZhhTBwRF4L2erQ41iAesUMie9P5UF+D
tHNgcUKrU7imWZmKdxYR95nYXrqofjwZHLn6lLRh+Jx302EfDlz0OHAV6BAfUSrI
YXFpqMqd+abb1cYg86DAvYcvD0HHmZ7LezUPzuPcKPG07/JonCoQ7IFJqru/Xkvt
D8dVMHPNSIvfCogFKU9WPIGDwqMs2/r0/nRYvMxsLeh9vkpjpmqGx5jDpaJS7dki
1SwSyvJi/9M42I4X6tdrOSHtd1v6UUQgPb6AHBwKl1QCLkvTDJJO+kN0BpzpqewP
Q6NqrN9yH7/FNrRcKyv5I0720Issea8tDSzdyCBX5L9At7/oRoEJ6kDERjxmIP6r
0xAMr+a7bCkjfcUBKWQK4cCaFig6Qa8JrI0/lLUZVuh7FnMSOVvkavlWZedgRZYi
AYA1Zz+M19rl4G2ZC7LdVgQLGCd6sxfulb1hP6STHTmSqacL84AhMWdfEYo5kKYy
R/2DHfFKqWabdlUaIfhS+XtkpPG90n4nUVqHo2C0+ViR13OjJRspd8w91fS9YUfw
fNUSLYquJGqnI9tfUi8q5X+Lhvq1fxHIumVWwfRNmzLRLNNVs9YR60vPJzsKGitq
Xxn7kdpjvC1ibXJavUiwL1K7e3xJ7cKvfvYtCs9hpE8046o2/a500EREN4CBRuKI
/lG4S5EgzdUwwfg5vF3uRhnbCAW71ctCjxoqX3HnvJ6ptvTwpBKrHvDXMSF0F0sl
`protect END_PROTECTED
