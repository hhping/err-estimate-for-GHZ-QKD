`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NyCScsjun9uPkesfXK3q+MkvSsWB1N0IU++Tlcr1xz2Yl43obsgnBd0oI/POKaKO
uey7iYkQmJ1fvr7ZJO796Or1EazcdgiXKeHtNkiPQTJU0c+fTxnZC6Ak0ncY2ThJ
xcnDfLtKUDzEjLaljieggIwWT3qmShuem9JzF6J8LFP2SlWrpvAk5buKdFFYVDLN
cmYIUSCoEGvu2EvXLewQwPDq/Z8T8T0x1w3AIu6vMtMQ5rmCFc3RtswtnxW+k4Rl
HqMpghNDyNPQFlY0Ao5CChGy21kCTAi46PCMclWcGM/dVE0Dp4LhCIKZVrLkIr/2
19h1IwotJUMZgomwXCPKGJl8xe+no7fbdTR4jl7mOCBY9HQ4BAqEoKuLaLe3NBua
J2VSrSsLZxsAHFG3WrJDUCRXScADNJrbTKkM2evrZg/Ln7MLmNbVmsghkeQT6Vwr
0nXH4m7JPHFLl6rTLbMDyn19z+0hoAXJVBe4yo8XOU4F6GRAQW8pnuWf/jJ+NQnu
mAIpmqmne/xa5f7Dmiq25P7NKwaBSs7rk0Kq0EbTsorAWDmQP1lBSUM7bQhEBLgf
8SqZoX3Ba9mzRQoW64pHNHh6mU4rqftnFsPrks4aeDHdHsLqo54EnvdkD0mRnHAS
ddii2mYiCI7qUI/mjFPlRgnQGSKxk3RZ6mlPLlKtQ1GdLuwzj/wNlpnH2Vghh2vv
FrCqZrwKU7+XtinguQSQ9Nce4nFA0TGBBYuxnCLhwq2lwbvctkpNqJ410R2zscXX
Yzp84QdioEXWAVFTzFWxdQowWJPbkf1SzYbrn+0awvYj12t03NJW1QcBi43iD/8e
FDow5m9ksrrOQpIW4X+ILUodCxCMLBPz55dSsShoG+Ff+Dzm/pL4VMq7vX29u/Nl
G+UaG4lxgeaTsiLTu3HIyv381sIE6SoAYd145xqyixWuyVkobHa20JMQ5banmeNi
oOG1i6C2IqdX0uTL+dRK/Cy8EpXCeqGa11MD703ecWRwtDdAEfjdNB6yyHkLjvQf
NiSrVG+m60a2+u2tcuQOTt/z6+OD4dbq0dO4vWpfjTggDzJrqNrOiS2fjJ8M4K4+
Q6KsnhmPQnB6ceP8G7r2ix7x3uOsCP3B6FUFc3hc8zaRtec9bfBL5O7Lsimc6Upb
ICm++yDiQv1AaE+bnqxbFUvq2h9Zmu+xrl0xqqh08NUSwo+rHbyUAvt6zZgt2c8V
+xXYorWUh8TTGMr7PBRIvPQbC1jOsAePw6imJHwfPhTkOHkS6wW+PwwQjNGqmJHC
DzpHXL7Hzuc2tfHHn7c65jRRyFC65gwD5X0wZ1al6vguMNynZFbVNbpmpwWum+jj
UWkTSVtokwWdKZjFR55f4T2w2uIV5aofkCvBKiqRLAhc0lqxn19ezRW77DrCFXWX
UMgZDfcqNugt/296jnAfpfBwn/vYKQ1pXCpHU6i8olB+1TOyUCqkV4SHwfNL9nSg
pbd+6WFYF6r8nQlzkN/82A6pajNdiyAWSWV9xx6DUq4XjZb/B7PeEwSNIyellGl0
27jpmhUwNL20SVeNQuanr3+b/ueVneZJg1KoDVYzhwnCWWxOo9PiD+97Isb23XVl
at2uERSqxEdjQmUm7DpQ+yIP3Ue0Puc8MJYSav2vQedzQfGA7VqY5o2eAo5a538P
8BIi+0aZIdLaIia9NJzJGDnz78j67j9p0LzrK2Jna/yMhqIPf9CByiBpMS+1fal4
lVFLpgkcsdOPKsk6VE+0pc/Ciiw+ofEpaaxqFNrxa6Ctc7KcHR5mwMzsFmzjqyJw
pCtqrGBEdwW0u4RusRBcIQqXiXzrqN4+F5epwQuNvP1TgwzMCiqAiyn7dcA46mDE
WKnSvBjbpmR8XKB06pIT1AR3su/3s5Hsg5xRX74Mi2R9zzHBJJQtq8rFC7/Uto6P
8Gz33pbsG16B6kKxq98p1umWtVD1qfNJeG4aTMT9IVUKOlV9lk2jzm5cdL0D//aT
jWdLUWQev3VRxm2fz3d9Y9XtlawGKV7TAGeiRsUidhWTifvbBiN5ExX91skCMUrm
zWtPvM5RUUbM+lhYlR6RnT9GOhu8oRZ96elfQFrRpokZVtxbbTf7Cl9VkPVopUqJ
swqXnCAOkYRMavCuiL9bwNH/UZhOI6qaQOeN1L1lqPX7atio0buWhC/rvoyVhWcK
h/b+cvrWKHKJ/XR3H09WigbRvlkh+yrLcqswZdQKD82Qgtwr4xSDgXl5pMRWPZaW
Ot7/hBat09RXK1Ht0GFNQE62fI7CD97Df4hjNKLllOeP+6KZAEASd/9cR/JAE6mq
`protect END_PROTECTED
