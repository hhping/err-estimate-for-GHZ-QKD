`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ncjgR2N3JT7nhPiBKCrbBggXpqXMRUuIlybcAkDd37Yd4FZdddLaFXjA2jDe9gF
/op0B8pKc4lwok+TOTdJYeyBry7AUMXZHPyHppyVkB8ZDWgPV4ZZdZXYVzsJlHou
8obVXlyvAhmmkZ5dVA/m07nlRDDVba4PQqrSwhSYLlQs9iIK22WBOKX/ukBxiNQ5
8PXwkC4cA1JkntmwKPP/WU6FrgWhdw2rdiHrTb3Vua0eulgoZjGhSFHuJ95Yo6c8
NxWP9F8/WgaBmTIjuHsDCg0op1zUrweNoOQEtEeZcq3VB/UUQTurDHyMD5Kw0YM3
ixcL6I/pCSiFmDHgxYbZJSf7zXnpHbplVMrYF0pwyVmUL6mE8iL1v8aq9So21qAh
FaX3jNCfwTy0on4y9MTECJwuEOqRiIsVQ7S2vc5p2hlSm0P/+UvfNn6aEauFk9K5
7Bl9VN8xKibPEJdQloGFFoD9BdewA3t0gDNu/9CHm6xBgKosMl/GoWHj6+NR/5pC
AWRWiYMjpT3lwKVwC/OJhKBD/xFJ9KKyxBPnVu+WonQkPhMYZuITh0wdV0GkDKoC
IawEAKoXMi8f6CmbYb0Y3vdXJEM/Jdv5P9Iw8crZvD1RqedOznF9pW0Imvq0PoI+
ydGuz5TLBYADD0bYIGsStVIfPem2989JSKjYvYEoFtrJ0LQcDx15jDnXmIW5xVPv
hVKqZ8Py1LoOn88iRuRe5PrVaWlL496chQeOnht3jOi+NIp3ukpwHigB/YzC31l5
czOaT0GSvQSXSimrLt1kSRUcUK91+wocxsslSReeVCmfQr/XQ/yP0xpwGvoe4peJ
ZzDBAQrxNSUl3Co9J+x07FgOPm6Tky4ExA8ZlVWGr0YnWk6icTLI3B1NoFK5Av9U
6//ItKT4blvrEBOfZohNt0NheBg98+1pfp9/+lwhrqc/2PosHVdwqv8bUHCPif5/
QFo7Jq628/JL04KawyVMwwRa9MVw7LXHSGBKjLv3/A8PAyb/LC5JmlT27cXKTRhr
r9yUSoMPx4555zWxBgCgafjEip5jgBuBmo9sskWqDVWUruvueC2dJNa7STKl2AXv
+3R1sF1Vlyb2fs7ZR7qYMqqd7te9rj48MOEQnvUHNKyoWNSYlYQqkJxJp6CmZczk
F+LT0rQP3/iKApCgbBKtBNCZkQ6Fi+RciINdAJcCbiUHDQ+/mM2DCNUldSMhDk7p
lLEbjR/MEnLNhF/cpdzsDrg14ZTz+wevdhMq++s8OPaTd0GHHpPl+i+QHsGfQQbW
xYJelpkKf4e61u6XHNQKhT0BV8GWsqTO5kKPnL53sNa9urWt+JXAjyGf1aO2lv+M
qh5xlIjF4vf0BYV3XyUJ7Ge5fvhDVFuAjt2p580romdGUtgHE7noBnxejUnUh2a+
YqacJYfXO9eXw0Whd/kYpF1D9EuSSwyKtK1uBEh/Hzkce/90hgmDGK2KRYnDwWP8
`protect END_PROTECTED
