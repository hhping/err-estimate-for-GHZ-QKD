`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVZd1jBOG+GI64kx8Ci6/riN/I3hN05AetgDP2SZt6Y13TbeVYWWOjlBcP+JNpdQ
fKjriO71yHZqgRg2drSE8rCDfHMhBLnR/DE8bQoqOnzYd3E7OOerUIMZHk9FJ/Pu
tEpHkea2J5CI3XkoKvAnJcJAWYxHtbLOQMHhNSh7x7Tfh89/3vYzFeCUldDOkFhf
nw2j5NCpY7OIm/6zgx8uYk13q1dBXpNsjVKPmxix5K0nMP/nBIEH9T1az/4s6T3g
J0ysFrm91yZwpZp0p6mwVg7GpSvTvEPUBhp54VmYS4Sb85UnGP3BbMXG/4HdJ5Xe
Y0eSQShl6fMtLeV+GqERqEJcp2GvjHqS9TTM5coSsdAFvlOJBqYZ/CYVhueNSQ90
mAt9ysg/jLbxkp7qb9w6Lm5b60NrWcgrsiQFRHD+vBQ7biJwRJoPo+Q5FzZwrQK+
uq9AZ+cA6Az1AR03+CxochB+BWDZTnkfGaGb964NYk0FiKqYcSaoHNRotmOqhvAu
dqzxbpuzxWh2LJpYfTz/5HKczbubMpJGOs4qG0o/zBcoDR9WlxKJdAardckcJJ4S
YqPAuemaSZ2nknJIJiz/rNYMGhv7wiXvZp/Y+540YaAKgDcOgC9isfaO1ZVj/hgI
NKTIMTxX4j6GEb/hfn3ZDpYJ87aSQcLH6bm8OsunN5eaCUCPKb7urX4yrWz0MpLB
90L5/T4KsSudSn3e7VjhL519i5gPZdb8nJR48fylu2U6U3xdglDVRrOwc/cMUImL
YMXb+wfxZx02nEaybpkPaemvqeZzpmvfGO43+hndqTL1qMDHMqssyijgX7jeGfzJ
kBgXhPuU1kio3+PAiJoPXxgbI1pLng8gyDMtQo6V9yvDN/RJ0Jo0uYCrFBhhDxcw
i/ahA/PaYycxIjb7VHEcI4LmUjeenjuC+zrJzZLhFR4=
`protect END_PROTECTED
