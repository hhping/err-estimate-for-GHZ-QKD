`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ioPHA6CU7UQ6F8ZzZF1eUcDyXZolx5gNblhmQWPaeH0bxMW20jX1FS8UyCEzxuJa
tUBEhmIkiz4cC+NHh5c7xgDct431D0JPVfQrVdC0Zp1kJAmKbmY5xujBGWYeqGVD
QPe9euX3mxoGOShuzW0N8LmbjPKmZGS6FFSUT581eIO2mHR8NGrGH9jqutbkI0IC
1XTw9SC2OeYGVbcgG3ochXhDv5NGTr9mjNM1MJxP76syqH8brGsSRLypFinatRrS
ux/TGGR09lTzkOUHRTNtyx3HyAxNo6zuR1Yi1r96W/5eLhb5ZiQEs7CAOHlb5oLn
UXigsCfpy+ZP8/AtL4y+6e9JKEye4Eo1k6gZMlUdUEQ8J5eOZNJAkq4eQjTVFzJq
AwfDp46j7h6O/7mzQCZ1RJO9Vk6HgFMR/0jW9YKFemDKv4cvQETVojjcheEmX4TG
elrYOG23/JeSh1p8/5ifbP5m3f5iSvPMD4pn3EIYJ9W0eV4HZux3hu1bx04+VVNP
fV5FJY/VslRvUoXLUeyJMunQmju0zQ9QnIb7FCmiIBCcPb9Yg5ED3auq6syXFRTy
PY82h4L77Dbv61JNw6MXoHZv6nwG7/kEZMWW8aRUwzb86duITgviMqL6iC+tu7yi
ksbq1B7HmqkwgW4FtFWmqiPb7+f/y1r6a6rnDSiXP/KeXqxyL7rssRICGpaBZP0L
4UeLFJMb2NsN6rzJGizLiqXBMjHV4gEIix29hgoP6iAjucAAezk3LNYc4PzlIxrz
xu/TbcIjOdOolGwCoSiZVMArfG7kXHMVpIY1KrSMK7pSRveAOS0tUTSHBxUPxtBv
S4u+FhYA8H+nHo/h4Yih51NOS8A+8HLyWwVpUVIs8RsEzBGTovW3fSGbujRYEqxH
0/VM379++Pw2/g9brtKtFw9B6ktZhQFB9QDBqo/oWio0Fpht2ecFmigvnpcP16/w
HtaGx3j0+b2JSeSK8TRRWKjcxmXubs9fScS+qOAUu1axBVfxV6TldQ2eIbDT9Vsr
FC2xC1+1y8vD6sMQkqTARrLFEDfd4qkBHbgXGT0+TQEBohg8yJYT2U/6D67P5Yl+
9uvkjGI6wdk2E6BkYtID7HFlVKrVrCE0V8LX+1aClRX/9Euv5E6MyMo4KGRF+6qX
eA2LTtxJ0X9XvyPvmHzAxXpRke580KbLdjJcPtY8m+mjxKMzEw+rislEayHts1FH
+dng/IgGIflsivnFXRUFjCCE4vWTdcZAqUkzZb6H0DC41qDpi7YEGF7fxG7LIHUc
WIXYnrNFiDxyzJMlY9q7Lc9WH2dq4+BrGFHsMuODGZU=
`protect END_PROTECTED
