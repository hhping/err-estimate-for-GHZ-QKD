`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxyPKnKZkGt0niZgiGmcuZK+2abllQw+3fMjZGXQAdl/BnLTyr7pK1DPdrXmoow8
NRAloA9JL7iDC4KWzw8XLcPVYuIyAmY0vQKV0e+SBKX7eVhKsUwaqHDgjnSY86Wu
sIRV9X4+VciUq79Jm8d4lY87EPGFf9L9oEkGBzl8jawjN3ZJBfZo2WMpIdhPacwH
B+YqVKI2mcdI3EpIfLc7Kg6DpVlXK0/h8RBEBMG5bdqt3dqlU+UGl2ahohyPqjEI
uF6gSLNFZM5e1DU+tt/S7qanfps/ePTERh7koIV079vmlMp7DZGavg/INGXDMTv1
l6qsJ4Og8od32R5r3Kxot823eJqohCJJ2uYT8jH/UiWXP7kvlTT0/FcYfQoMok1a
c2dbA1TraHl0bVVzK0QRMSw92nFdVPhEFHp7OdlBz4AiNBnh31XCa2rgY1OZjEBD
2AF9TWHX4LzVNmMgLFET2xvsx/cYCSbUlqJXwTMFewbeS8xdoNLJaHS4OI5r0OIP
8nepQkHaoK8vnT2PDJGHKPeV7+MwDmd5yy4I2iBHK4pnTrysDjB5XtRgIJaLVcDd
XW+PemAd2T+KZLToq5RT199s31+oiTY68MMGIiGkvT3HX+c3VkIFdFkLMO2FslZV
IDDB91jkCNbrbMhn/q3agiJ4hx6g2+//51Urx552Q1eoT24qHgXBQ09ZrdX92vK7
OcUQrceyDFQPnoXrlPFKNhWpLsWxk6jLjhv0T8Xi8G6XYZsbYu6CHdtdM7UtpXG9
C5xPz17KLmurIuo87LjlVLagVb6W5CoBt6KTzTWFw2oyeusbgqk8ImGnOIdO58+w
NMVi4GEuj/bhpzE44ouSea/VFiY+BmekkYd9DppTBHRjr3RUsNzq3zIZYw1wzoDY
Izo5z1ES+anBZkgI+O/ohB73md29hLiKOyP1EhTITcDdIgDU3xLtggWtDWGwA0zL
Q6S6RqHFxDc/o58tvadyhz5CGcO/wBrgRWrZzb05uVqD0z0OdNYzPxqUs3YfgyD4
dooSh08kqcQ6YGjXb0NTZYkZ9rObF+6I6qjE2v8HtZc0oVTgRtzUzIG8CtdKjpIn
E0CVH5oiSediCm/h/9mYbNqaFQEBIS7mF5GGifQpQWEJfCAUodS4SwKXVtCzf+yk
nmGQ93W5yzsxm0uPLqiIInB2E9thRkYWegzI+BZatsqxXwwmKjN/DwddW+jEm0op
C0c+HTrMPECRUNwGIJ9n3nd5KN48x//H0idHP3RFk3S+upxqp0dq5KqwYonphQiF
5i7Qy3SGoPERNHThy24/JICe0toBHW6qsfcNZEVJhmFwzKxNxfZD4gY5PLA7LpQN
9G/P9qQxqEaAVGVSp3j4nnKTtlNfd5DNlbAltZZuVxZDC2gZga/hGNUcJSsslQxt
D0UU9OQnig9OFJyoO7sN5HyuOrx/jTcxfp3uVUcK8joxAkNzSYKrJbBgGF3rZlF4
ilHbp/aXsxWIV7Fwf85tiDBM/NKmdnOvJ6Un2bkQspfCj5yVvMZnVc/1AmVLTg4S
dru97wyp/zP7To9nN7Cpa5bm3eSy4oLaBCNAnz4NOmGIve6SMBMHPN5tInaFPcjP
Kqo3US7jxZoKq3rMjIC7qjpTKGX1DEg7afH2V0NinypYq7gBwbcMzdUy3DnAX0+Y
zYKfzjB2LOxuaJmq5HrYK4e2mi0a1p5N2Y20VjVeolB+SxnOJKHR1q06Ywvl/CCN
FSO5yayyXAsqkNLFF70thFE5YcG/2ZMaRamo9e7HuGcQLyh6Et8rFseDe5Epa9ce
IdT3nVRf81VJVYn+2VSeDVqeXsoDBWYcKjiVB1l/0w7lNZnnMX39AjC+lz//xsCQ
JS/hsJkFmS+no15Jj1m66asBqyYAvCYCemXiYWvRY1Mnex3hgwJ1sOSd4tmyejLE
hb2pXTU+OwwPAT1DLgFNo0eQr32F4rYjKrmN7/XxaVoUtZ5LyMEpk7hN0jnpk90t
Omjvslm85wFkLRU97dtk4LEhR/zMoqWLqPtAxuTvY2/S6mvw4VsHCvibtArE5CjL
xVy9Rbd9MtMklG4neYLnRx7E2MO7bAnCkIW6SLxs70/KOmrMkFK/n/kFg6urRwCV
30jRKPXHcFHojcHpyRmPACCXe2kDQ0x3R9opgPa1ZsJi9mXQsoDGk0xSjcTo/A3b
R/2PXIKLilRzoMmuOIWIVkpWUNEbTBEs0KAkImBD64NacZfnFR3WpSPtXcRsKMYQ
3++OvVfyOvJsKTROm44b+FLq4eBNeapd8VU6EgKcSIb9yDmxEkfRBsKHhB2mWt+g
NJvytXy62aUVvli8lIcu5rEUplvu9MVDc5RhRmIOhVxrSpJCrf48CSDdfpi9LA71
s6tRpXhcRJRpwd/EAsvyzSF0w2g0i6ykKuXu8ym/rXSNBQWMNPEFGwwer1+cuVMX
niccntVvQqqlRx3buzlTVvzol09/N8eUvr6C4Cph17lBYsZd+b/eFL2xfFhJaYOR
ySx0+ymRFbW4fVkweXPhQnylMh28WfQ9IAv15Wn7ZiGCDuwM4tK8AQUXlkYLFS+u
nJ3siE/egJ7WEwTV4+ljShVaN4Z0tl/jBkz/hDw06X9Zyj14TRAGQ3WWIonaGr8/
R4hH1T6X5tqxd/uF7wZg6N1eKPnu6JbBY+sFyqrocQWzw6SrTejmcRkSgyuVDZky
BQSwvF64Zi0yCUmAqaNCEvENSoqYKiQgEmtEAHhStXg8oBIm4X19KTO8rWtzUHKQ
wYRDsGRuVNEt1RWqf8D6+gTmjoWDrBmrtoruhYuXaMZNw0i8tYo5bN+XyeoEFaqI
CUhwdCebcdPfOflwjn44Mhfvm28rypf+GgB6HcGFJUuj0WDWBjjd1tlgyUTkuuJe
1Kx5ElhXGCFOHyxsDDmTV++JUMBeDxd2j8hhy7sBBLShXFlNrNkXoGiGjbO/NQOG
wCxu9B+sKlqOlJ2ebsYDdcu6oE/rkV9VLM+9ty4EAo6RnjtkQj27WV52cAxwHoZq
9J221I00c+JwlW+ifWgrvyJPKSgbuBhlkzhzoWGCsjgFK0bDt7QOS5wZdc2oKp68
98sG4l349yvK9CKsak4GZ1iqWPtyoj4hNaZ2TiJBYA4UAI0jN2CfL31lpYRTAV0u
MmqXMbMDZDpzbr+riAD3FbYzg4RdPO3tCC/VAho1RvuspaYODJMDj7+jkS2Zo+t3
dFXZUEnNAifQ8ekmQlkvOe8k7Gb/wREZogc1M/7oJzCh3yfatapn46HbOFCpkUGc
pIMcAuOX6xkAZt9lj3h8FAaOfcsXW+d6D5ZpziS1XznHQZvGr8Jv2IMfFMhn2Gdb
bznEzX6jz4mlzQGAbqvq8gq2zUKV7jI8rliqhm41K7iLqxgI/8Z1opZlbU1EhAeE
voWWRueHlG7uW+5+nytLdwdlNcrsY1wz10aNQRaH7kV7izfJiyrxFmgYLZepYpGN
PRVM3WAuF7GHxWf5DbQ2lBBSYcdFubr6WsS/ufuPvudbqSiAcT3kBFtxLTBWPMp3
qPi3S0MOk/LoZSApaUqCyQ==
`protect END_PROTECTED
