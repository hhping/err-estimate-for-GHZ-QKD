library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_rx_dfe is
    generic(
        enable_debug_info: string  := "true";
        atb_select      : string  := "atb_disable";
        datarate        : string  := "0 bps";
        dft_en          : string  := "dft_disable";
        initial_settings: string  := "true";
        oc_sa_adp1      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_adp2      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_c270      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_c90       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_d0c0      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_d0c180    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_d1c0      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_d1c180    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        optimal         : string  := "true";
        pdb             : string  := "dfe_enable";
        pdb_fixedtap    : string  := "fixtap_dfe_powerdown";
        pdb_floattap    : string  := "floattap_dfe_powerdown";
        pdb_fxtap4t7    : string  := "fxtap4t7_powerdown";
        power_mode      : string  := "low_power";
        prot_mode       : string  := "basic_rx";
        sel_fltapstep_dec: string  := "fltap_step_no_dec";
        sel_fltapstep_inc: string  := "fltap_step_no_inc";
        sel_fxtapstep_dec: string  := "fxtap_step_no_dec";
        sel_fxtapstep_inc: string  := "fxtap_step_no_inc";
        sel_oc_en       : string  := "off_canc_disable";
        sel_probe_tstmx : string  := "probe_tstmx_none";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        uc_rx_dfe_cal   : string  := "uc_rx_dfe_cal_off";
        uc_rx_dfe_cal_status: string  := "uc_rx_dfe_cal_notdone"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        adapt_en        : in     vl_logic;
        adp_clk         : in     vl_logic;
        clk0            : in     vl_logic;
        clk180          : in     vl_logic;
        clk270          : in     vl_logic;
        clk90           : in     vl_logic;
        dfe_fltap1_coeff: in     vl_logic_vector(5 downto 0);
        dfe_fltap1_sgn  : in     vl_logic;
        dfe_fltap2_coeff: in     vl_logic_vector(5 downto 0);
        dfe_fltap2_sgn  : in     vl_logic;
        dfe_fltap3_coeff: in     vl_logic_vector(5 downto 0);
        dfe_fltap3_sgn  : in     vl_logic;
        dfe_fltap4_coeff: in     vl_logic_vector(5 downto 0);
        dfe_fltap4_sgn  : in     vl_logic;
        dfe_fltap_bypdeser: in     vl_logic;
        dfe_fltap_position: in     vl_logic_vector(5 downto 0);
        dfe_fxtap1_coeff: in     vl_logic_vector(6 downto 0);
        dfe_fxtap2_coeff: in     vl_logic_vector(6 downto 0);
        dfe_fxtap2_sgn  : in     vl_logic;
        dfe_fxtap3_coeff: in     vl_logic_vector(6 downto 0);
        dfe_fxtap3_sgn  : in     vl_logic;
        dfe_fxtap4_coeff: in     vl_logic_vector(5 downto 0);
        dfe_fxtap4_sgn  : in     vl_logic;
        dfe_fxtap5_coeff: in     vl_logic_vector(5 downto 0);
        dfe_fxtap5_sgn  : in     vl_logic;
        dfe_fxtap6_coeff: in     vl_logic_vector(4 downto 0);
        dfe_fxtap6_sgn  : in     vl_logic;
        dfe_fxtap7_coeff: in     vl_logic_vector(4 downto 0);
        dfe_fxtap7_sgn  : in     vl_logic;
        dfe_rstn        : in     vl_logic;
        dfe_spec_disable: in     vl_logic;
        dfe_spec_sgn_sel: in     vl_logic;
        dfe_vref_sgn_sel: in     vl_logic;
        rxn             : in     vl_logic;
        rxp             : in     vl_logic;
        vga_vcm         : in     vl_logic;
        vref_level_coeff: in     vl_logic_vector(4 downto 0);
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        clk0_bbpd       : out    vl_logic;
        clk180_bbpd     : out    vl_logic;
        clk270_bbpd     : out    vl_logic;
        clk90_bbpd      : out    vl_logic;
        deven           : out    vl_logic;
        devenb          : out    vl_logic;
        dfe_oc_tstmx    : out    vl_logic_vector(7 downto 0);
        dodd            : out    vl_logic;
        doddb           : out    vl_logic;
        edge270         : out    vl_logic;
        edge270b        : out    vl_logic;
        edge90          : out    vl_logic;
        edge90b         : out    vl_logic;
        err_ev          : out    vl_logic;
        err_evb         : out    vl_logic;
        err_od          : out    vl_logic;
        err_odb         : out    vl_logic;
        spec_vrefh      : out    vl_logic;
        spec_vrefl      : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of atb_select : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of dft_en : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_adp1 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_adp2 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_c270 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_c90 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_d0c0 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_d0c180 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_d1c0 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_d1c180 : constant is 1;
    attribute mti_svvh_generic_type of optimal : constant is 1;
    attribute mti_svvh_generic_type of pdb : constant is 1;
    attribute mti_svvh_generic_type of pdb_fixedtap : constant is 1;
    attribute mti_svvh_generic_type of pdb_floattap : constant is 1;
    attribute mti_svvh_generic_type of pdb_fxtap4t7 : constant is 1;
    attribute mti_svvh_generic_type of power_mode : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of sel_fltapstep_dec : constant is 1;
    attribute mti_svvh_generic_type of sel_fltapstep_inc : constant is 1;
    attribute mti_svvh_generic_type of sel_fxtapstep_dec : constant is 1;
    attribute mti_svvh_generic_type of sel_fxtapstep_inc : constant is 1;
    attribute mti_svvh_generic_type of sel_oc_en : constant is 1;
    attribute mti_svvh_generic_type of sel_probe_tstmx : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of uc_rx_dfe_cal : constant is 1;
    attribute mti_svvh_generic_type of uc_rx_dfe_cal_status : constant is 1;
end twentynm_hssi_pma_rx_dfe;
