`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EUF0YFeh36RMZ++TM5ZbpW7F6j8/RZ2+Dl4Rf4u13U/rNoq+BdqdagSar6aLpK9R
dFdr4Ady+wNztnHEwOfbeNv3j6ui4Dm8mJOx4BzWEgo8ZT6JPjVJvw40HFLUhYxN
U3411Gg/WaIILJqWt47/hSiQQgg2KKCMtu/4ZTGzQBghOExC+jXhd3Yt4aXlbVKV
7nzJvW/3cvvVromd77Zw7hx2CUQudKBBhcVEEiJ8WNXnn99F/vqA4U0vg9rmPmsP
uLXhNd9wJQYvwXz3YoD1CMrvLND+azDNso/+J0/97xz3LolZ1VbL2C5u/KeTK+VS
roxCN4M2yFiDdBdu/RXr3IS/NU1nuPPXrWVsQX5Ey/ZditugTZcTEG/3sxjwy4Kc
r0lTCm/6hl1KdT7M4MlWFIlz5vX3ZG+n/Ll05zCXZjgZV6PJiGyNwTr3qpAjqRIw
oVyxdf8FnjldKRdFhD5nHp3n2LlMF0/NgU/daNP8FtkMj3A4zVcDPZ3wFA680xY1
FaRmvahZYPwHtJg7cySFLW6z/n3oFLNTDCsKZvSqsTsOisDJw9MCo0qnWER3aIpC
YEYHswZMv11BF+wO6TYQqQ/vmVwkfZ62Q72FH4ddugIuSwuMeXwQ3bo8NzTh3eYA
OY/7HYsU9hnWdBe8xw5J2fJXozSa/OsWxJZPmauaXaojmrDeDkV7i6KhsUqPwxXr
kC6GMZbBzrhu7asQ5FmG2FnYqvK49SQX2721EGMdkSs89WWPiHgWpAh4Y3BX8pWr
HF9cFNsNvgEbm8Oi++rgW2o3LqDHHw8SbvdMjlOn82Us0QgNGH5Ch3rSMsveSlyv
NNOBFgo4g8m+cJTmqI0T2qmAQUJKwVJsh6uXGjdgDxWbq+VdtbqFexQEpjqhwCf3
LK7y9rb8BoG3g98sJJvH6Zfo+0kHXKT80OIXJwObt6rPjg9EJL4QoFpHUqHAySOT
rGgsg5Z0epuXnmM+fntttdEnOKbqGVG+nWWMHxgQrNAcErr5N8ts5VqG8KZkesOy
LshB8R92fof3wC6fsN+Qp6A8LoyS7M2iG829awBBjiKaEIdiJmqVCA17EmJrQ07p
rrvtSsy0+VjlzHXB4PYFS2doNwLGJ8i3gjkzyqkVfsbryZsHxZFH/TfxHF1tFFdt
vegMJo1qJep4oLehfu06i4tu7gZcDMbjAM6rQQuIfLw+Nx78znTXNhdKa6buNUBH
01++hho9W0AK2t0ZDesMamH++4XZ876E20QGpuwMVqyjfHfRCNE5xWWrUg5gVphn
HcJ+vzor6LOwj4LhU3tTQNK9KR4UarxAzLwNe/ijhaYbkH/eoZ4qZkLvVvHacmFu
ldbNAZKi17NvGhPSggxll8trE8ZJjvDApLDdnJk1ytlijGxizkra+HCnkWVxA1Of
JcfpqY05OZyhRs5YRXtcZ12ihldVjgnTS2qWwF0YMl7LbpfWPfHprj8d4FSBWA2s
cBwmEkphpbxygPNS7UbfPgPb/SYauwROeLbfV13mC7riC/cAo5ZkY3Z3e2VKoG8B
ktenhcMPzzAtPqj5LQDMFB2NOzWHfxHSq2lyCZJ6jtI=
`protect END_PROTECTED
