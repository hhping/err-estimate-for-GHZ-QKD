`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EB7NTPJSBqTwaIkZ3NTzU3Wc9ZtvKK+BMCPVRDowM0LB4dTYzh+N5859BiZLo9bG
pR6DHvJiLkkeE02xaEacnI/Jc9JBVDm7Bbqcob240oG9L2GiNOUXOJL/DJmzQVUN
uL22jP7kQNcHCeTx+8PbMkqu89zcy3pZ/wYxzYQmAj3TGRJkf/OxJWRsQw9LgD53
gKi/PyZuVlV2Xxw88f/JbL5krXGK/9JHglq0DrPy+ZSo/qTXQJzd61RpCZNYRnM6
XvcrIwHSgK6EC/5ge9p2Qr21gt7t/N9+rMqtmRhgzHGy/KVUMNNBKR4PJYRMgwMd
Qe+jT7Hz2rD2HH09UMoNa7GvXrMz9zo8e4583+yed1on/2HSABh8OQhxgkNzVsEa
TMw2HGxY6h9gJAO0T84MZRZclWLK7QhJhs+q2d+pwKPnL9hZhJmmQIlYOq98Qerx
22lPe9twYdUAbmeTFuEWbyXQolqhqameS6taFsQiISSnyN8CTXoXweAaOU2+qNTQ
DkBw1lSZps6UlSo6k9VBCWh1PZGtNMvaE9AGXEIBXBU642i3hDpFPOmD65prM/Ki
tf7cGmTv8SDgtwS7aussUjk/ZVoe56Rz2XSQDJlEqKKZxJITJm9DV9T6xU3lA8XY
ViYcf3Le5x6jlokITevtwztmdettEGft753QZFh9YCQjsAbj6Razqcr9HSbwshDs
k4q9mJd5VZCGCoBg5zlu6E31bv7UM62IelHTDZd8xt68OLT+/sXt0y3ibApoZXcQ
k+x6KpmPh46NFczpITiQX6oTP7qzO2NKs8MpCGEH+zDxHBcEM0a7TH9KcgbIYLeT
7vFgRSUbuaCIANMHlG/6YQiYVYA5hwTD5lDZjFnzgUZyWtJ1Yq68cFkGaMy5VPSr
m6Hn5ywEYDBGkBaCUJlPHmGtw8lIS6HzEAo0/FIQKSfJHb0hw8sMwcbiBxIfXxHn
rBFhaT6MXJWTBQFaqnnZtvHRBDwPyqlL77buaWh/+H+hiYjybteOHEiRd79xhRk2
kn6wZ/V+EQ09QqTUR0GwidhAPRQvzrIJqUfYATpI3CTM0pK4cqTfQk+PWA3kWgXp
A+lmNBDEg9waNGbvF1d3Gg==
`protect END_PROTECTED
