`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+I8GwB/aK4ErESiXFIbGgfZCw+AiXoMDNUYoZsLng/fwiBfenGaFkNa2KE8xNvC
ockVWUVwWB0r/6joI92SMV9vZiYvQ9OiUZboSQPaSOH6K7ns0EJPs01xK3DZ3Heh
TgHEfsl2Xy41Nf6zBJAqPBltvZ6i1jwI9ra/BpYjb0n29bkuXPmeflL425Ypu3y9
Gl/dPG26jvvfnAuhKZYauCYqEhEisFu8iYs7NO6n+anCDETIZmUBLcN+bbUNuxcm
ZouhYXNlXhTCPMZk3H+ol91/rmbUGbmD1ZyVdRIe7fLsPj3vMzr/y3ZTaykv1RAU
YTI4E+58+b0Uj+aJLJ1ADJ/ivFykW4DfjmVuEnauRqUz393k1mROCGfCBoIJ3j1l
GdG56HL4S8tvWQ1DPI8kgPX6bX6C7bPxGGC6s9/2wZ5Eyc9owu2ByOXccUrE6Ula
A1KhBrqeXIspg92sUn6KYSfjLhM20+CrEmSts6kdM9+xy/v/AeDMIFH8phQcIEod
QtsbsfSgVBaanT3rI6tSDbNN2vOWAdHxzu7Y6pM4lGsXcp+yH0zc4X97M2lXwPvK
pSI1ZyJV1whVFsVa6Zj13vmpkZyhJvyqblrQg+vttUZ3TLlk7kPzVUAKU8fU4j1Z
l1l+jxmS0kbJG1o0TUjBXduoZJsk4dN/cj7/+L67WLg0fS93mScbX9+ZBRj1NZa1
GRdQu/ml3TGCTHRrtgQ3GeXr+TgnwukPQd3oh6Y+h9EyXTPz/XUOhN9o8INFSbg1
2A6zJoyNzSkfUwwI+txZcxOU+EgNEqeaeJ4JYES9KO5Dgc8qLnulCBAqWvoJVpKn
rWNseSyo2iUcUY8ejn0D7rHZLSLju+oIvSPkkgr3LwPA42/CGQ6oqo7bYJLbrMGa
ZyNrRhjoAmmaD3UBCSkPkTPj0klu8HBVYbE2JjIxjHt6AMXLTZbfZ1CEEFkFWpBz
+8sWd7DuT7OcM8P1obM0ZGVWcIyOSMkKbaMx/nV5WSEUlgxjjuG/aro2phyyLaTi
T0PQOb+9yFNYKohQt5qcz1YZ93XD1pvYfAdPXiHaKR35ZN4pzC3ylY7eP4NpJ43o
1seLjtUTgb97EUbNrza1mZRjVKNYgTFa/TbvubwW8gIqIkEvAZonLTL1d4F67u/e
gg8DZbSLkT2cSY1UMrujiMV1R+RKu5MPVa0oBnWkjJWdsKFhncjJqYW1m3xQEmY1
hZWwXFyEnrG4rSP1O6gke++XP425xnxZYmEKSknFPwEDer34coR2FmiqElcREdCr
nWxCCpdrCFcROd48/EMIey1aj9iHnoXCYZR1IUJAngyfLBoPIySILVvce3rOdopT
ToinVfSjgEk7SJ8/DNbKapaejPKB/w6IyK5LpKuOzPX4P0m4I1jeFaA8FRSWJlnF
bouXcdjS8lSZBboH5L6RGClCBwkx9ELhDuZmCZnw56ZPTgYpVNdkePcKiKULaKpu
BNK1aGKJgdOwXgYfDbddy6wojHiSmXzkkojBaDHDopn9uIPHGTf6npN90S2W2x6I
FgVO3uGZui7SgjmtUuh+24ghwy1FxqNJUXNy23fclYzSQg5Ggsv7d7VCg4M7c7Su
qUx9JBgBUrE1nJ2kCokMT3qDkAGAFpJAo2oAT/A2WDIyuPylX3EEbwjojEf58gbi
USXT9/ygdy+8lIm7EK7INS+Bs2adzX2CMRIZeNwecT+Q6KxJSIwNj0iMa1dDklWn
5OGQKGxECiNFWGwRKBlBsa+3L8FjBF8mu6ngoNFzUvHRGzt6zouJrU4V7VSh2zLt
2e+QJ213ZP1TLpZlfAAxMn2VGxzwHwIX6hBu45gaHtb3jXXUueNMxRRO64cDJU64
EEJC8m6avb4z9Fd/5xq4xEB5HVl4dUXAwnO0u0y1r5VebNKhMchHX75C2dJ//lE1
0AMErxAAkYnzV2JsjLAIhemJaXA0V4WSvuKc79NuifmChWSsPKQvPhDHJmYFQqx8
0ieY2KpUw6sQcSfOoLimn5KO8YdD14c87dOqko81yK+QiVB3CZc4YwBM6NbOgzS0
VzLcezq0bXwy5uh7i0PYqSORWwpAqFowzpnCcC/9GJIdIjwvNbncpJh+6Q72OTRt
llm1uNsKZh2FGIDoVkBxgQ0AfkJeX2JYVGNK8X1d7GPV5x2jtRIu+h3rSTFbTNZT
kvbkE3EFHJMaZrc5V1d67GgBwHmAHntsyr63zxfjuli+cgSBryhaHvwz9Lab/a7v
9knSLHdQMXfgVZ4J8bc4/32fWXrgE4Va06p3/mABKX3v212wkfEMYLlbczyQTOuK
KxhBbEFE3riJznWruGw6FWWWamej/4Kji9iAvpUh3bwo63t/yANbtQgXzcdJz+Sn
3teG8aG1JglEktpvoNRMayWcBW8HRr1EnwuA+10L1DdHSsqwkmC8AGFJOFRN93/g
t1DqO4aAPOLmWCsG0nOLu2+z8Xr03fvtUFMlCHc8XyB4TnD0ajVnFmbr709y2EYR
5OwqvPrhQbtnUG5Zq61Bqsuqt3XUn1+nNoswxWdRmHaSdBY0zD/lj9q67t1xPUow
eGVA2iSf2fnDH7AG8YcwUG2isWL0ax94FgYYg1YSCZr5Ewkwg4Ltwhqa7eqj/Fa4
SJ2fFf38rfadgUBYWHfvrGpYaqPXNa96yl+5Bif9Gkx4udOI14+Pt88daxSPjH8R
ehY5qyBlJBlxHa9wNPv/XCuuNL7aaQiUQqeugxUA0qjExTuj103tUrcXzLQmP+wn
2mGIy+0cJZwUE9YogUrY0CwpEsKtfVpVDKNCA8thLIPSK0m53Akh8wkLC74thhqp
WZHkPdQxK+pTiiqZJraBT4ISJHrrf8qP1naLvSmDrCi2jEkUKDbP6y910WeBOrjJ
uRuZe6uOaUkzFC8+zV1vGOz7V/gJL2OT3U39u7jtcZ/za+JFLugNorNBv6aRTHEk
+eCAPlBFIBcIqXdJ2tSD+aV6KqpnUaEjXhRY7lZrIjapYQUCsXmZYt7mUgxMj58F
R1wY8iwRArCFE+h9BM6LugNCx/hiqkN4tpRSRW//ScnSxhN5gujhiphwAOkKc0NA
RDLWDY7jw4cKy91Vys5f9QXRpK7MNuGEFxgdmI7xLXA=
`protect END_PROTECTED
