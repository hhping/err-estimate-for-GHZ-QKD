`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eX6p5vsuBwwtffEj4zzzk/Co7alhpIz/3SJ4JkakWKxpgs6ZQflBGSkujkX+LH0Z
49mzdqhIarFrJwaXopR/Zprha6LM5Xxe/5cMg3fYMWeY2s68HPxnk+sXjKw3wsPo
Nt9ApXNirA7/P/qBnBktcCCfBMWlXUlqLwgxn+ipBHekqkCBJ8yM7neBXIK4GSGM
FjZ1FQIYEg6M3riDppvMCJ+V0PYFj3njb+Gj6TygXWaWrF7YEnO3oo5MXK5Ak2/Y
le09ngWw3TPUoIXa3kuJIdZ6+9SGGauY/4Q7IKMYrylU9DBNLXrgfB91JdwBtTnd
kK5gKFsIKmEWCbsXqswtGIK17fvM3NDogz5VW1kCXzQsy2kjOCnEJGB0yJaeVOeN
HLvg2DN3iUJCKHqgUQ/tMw==
`protect END_PROTECTED
