`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dw9ws2e7Sl1f0sFPZMPi1zBvFNe/kETePLhhSIWjbR7/Q4X0hjMzp09bIutSfccX
Epg6AA5Go++BuPOSGYBP+Ug5lyK6d8TbDJyEmko5gZWtSR27X7tWwofK1TNHhIa/
QLpSHDLniHVovc2JIInUkqQMvb4JDOvmvlhJQVmwR0umG2F10f5WA09i/7DsjsRX
/1Nn86VWGkQA0bBwmcDgTNzSkG4oEg1JQrD0zyu33DAZcfSTGvEuvcjCp8aE0TK/
X6kVyVPPyh2AcU+L8FWpiZwhn3FJ+vtm1WMkZRG6J2Bwd7bTLDkTC59XDz/bGXyT
cw2LPq4+PonHZ0g7d5S65TP3ZmxXPfrg772xyPNwApnJjzw3Gjw563/xV4b5uf4+
W+yg15yow2XhLksDV61kR5t/WCEvVY+yMGagMfFA5NQlvkGvHuGH8tyj8v0P8mVc
b/uG/Fv8ewwLoqMwIJNDx9G4XP5OobVhng3VbC90voyk5R/+OeHkXsgbfOPfSvP9
DiZ22hdn0TKeTHgTONcs7JCgtwW86un6ZrLP7byx0X70XO4+WNOaN6uhwx4zJu68
UX6fn8DOuznniWjoSqHSbW4EI/I6U32JGPoAwA3edcJeHejuYKfXjNTeVVf6TD4Y
QyKVNTfXGbYsLSK+ytazpcw/VVbTlvsPxkYM2ljT/rRQhird0bavUzEaJ0JvVtAY
j/kHOb2y8D4MoWf5wsTy/zriV7dH7/Yh7pBIvAfyrSHFySt+ta9M4zKJpvZCeCEI
LJUDP0GQvXC9z73mFKFopLPwiTc/orQKVlZgN9z0fJLCLvU/G+KC0MuaSmtkOmwb
slC6QZQwpXlXEWI6O7eSA6RtmlrlKuFH3ZC8a/w6dO0iy59CiPBVZVCim+ZwIcBp
nN+blZAC4pOE3fOMsQw7Jv28SnT+cjwti+5QeHlhEl5J9xQx8CMb6A1QcBW5K3CO
sjqhEpPRCAUfA1YqmXtbLJ5yMKb+y9CNfS1fAv8g6SOIJTw/u+HxSn6ePLqUrYO4
ZWHM5eyiYpb/0DdL5/lAIMRZ/pHO5uEaapI2SwUEE2c8gOEm+N6LyYFBH2Mm7y+W
`protect END_PROTECTED
