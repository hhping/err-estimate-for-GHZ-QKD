`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
927oIzHXosNlyPcnvdaF6xfE0ANTosmtUpvP8eettn+17V/VbyG4e5ulVeha/Z/5
h0W1XsIKgr4FTUtdy4/BA5vDGIAfrsMY9Wq0Cjx2kFiKlPcl6bwSa1OCeNPtqR1J
NcspCIc1jrhQDVNcrDZnlVSGKZnd7QjYq8CZKkuKpyuJR1l1Mz2s29P1HM5Le+aY
Lca7amKu+wiWJw0XfiigktmkzmuQ79CeEt2kw/5xLs+UPjeO36oqjAFL0Fff/PLy
NO8cVK5dO7HirFiYSW0eerfUHywVJsZWmwzbPhL16OPMxLPgpqPSJGQNTuI77vZ6
rZfmk5Wqbly1Z/W+XOLGmhjyxcGtm3Nc4z3069oOka0i/aYosqTKX6v9Co1xh1nh
IxEKzqupoduCMuSfB85WdQ6uVaFATDISmhZs8nQX2g40fDo/whsfUyjP46iD2C2i
ohVuDm4nsnKpAdAZgDd+Vn39vJPv4OeaDkjC/M8RxztcLNcjQaUHtEZ2mgwhkZYz
oA9BCdQqhIcEUBZcYNkeY4hPbIeK6G9dz9Zu2SIOslYhQxWFjP8Fu1ifUeYDbGOV
WqT+Ek1LwI6xiB06uylzOOd6HslAEdRDy8Vxv+LaPGklM+tZkJTrsSGRfSv6l21m
lgrewU1uO3Oq3z29Ea03LMT6EqJJRN28rEMBJIUcw2639tQC2We6QMkBtyEPZTVP
gi20Wmamt0ENMpVFkkGFipaeonwiY/OuRLLkcPaMOUutfdIUw709abNdamMZg4LI
wFDDoiQk1vQ7wyEo+QgV/dZ/emQ0Gs7Yd/5f4KM5zQd1svN5fkAs87PPqvgL8bk8
OhJdqbzrg4pIwRFdRqrOSV4euop8wa26UQ0LTbGA/wL1nozy1UNjIDOEwe8t2goT
ylzBS6WhXKMQmvWv4byoL/H7+ISTpT4wX2PVZMij4aDgU9qeQcnYpJpbUUPx92va
kLEwLpHi8O5WauyY9a07ufUNVr/wXLBLLDried0ec/LXthrLlMTAF2RWyS2T149J
OjAqW/3XKrPO6s/k9KIpqEW+GviGzDSD4BWOIDhdkZI=
`protect END_PROTECTED
