`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKV8UMLmk5aRK3kAYiv8EYuAo7ld2pLpq/XIcK4rCZbbCofYVpovvsHvrRwXKbC5
dejdiCiSVyMw7AT1qc3eF8AVwngC4cRSmqUy3x8+8Wcqo8KaAkktzpaRF9KejCl9
XNdIHItidPrGmScy4+aui1hw7NUbYaZKFNkvbDfS3CWk7JBwPyLzmr2mfr+yT6vz
KD67gQSLLVQsW2anK0dkKafP9hzz3MsP20DotcQgvrxGLEgRL+h4nh+xWbCVFELc
7Rx3LtfysZeTmj9wgJ0kyKz7Pn6vrmx0tnzjUXkRxa5GQ42umdoxUrkuLSjO6I5t
9iQkzpCE5o604H/pWoogGMF2ccIJnn0X8W5a/mWuCRMpAkv9K2jMGHVZMJ2fcdcR
Ilv0V1BgEfdE9NA3yMQQ17EujnQmGgInnc7u5RLpywTJ9HM5+gYDsLn5PCKRohvU
+3mGu0wu9jkf0xDZW91lK/I3gBLvJeHQBVsD2G49SEoTsJL5NF6gxWx+pMVjbBGn
`protect END_PROTECTED
