`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DA9DMfNpDJ0GsqVw/s51mw88m09QhjTTyVsM/m4ill/JEWJRAqSy+JDEcKx9WQv
6jL9/kskkTuzkBtitLQl/OvaUsYd/dBnzq4nTuxqvxZAd72xNMwR0D43Z+Y59eY1
hxQ+kNnjG3W0oth8MBmq9q5cGcYsi6bI5Ub1gEMJhHhnCYhaOxdAKkHlAWksA0I6
i6cMS9nf94YsK6haEu5kNYW7YsmI1vFcEYCC18JK7v3GZeUV2XjBVChGZ9elc2+V
93t9yo/v8RPeNTCgbvKVdoje9jyE3yeXOLSBwMpJ42YU9XSPY3awufXbjU08Ae6x
cur4bSr5LaxfruUbWlSBB456TWokZ/Zf6C8siz/WFWUcTfo+b609y0rOr9M6Hb8F
ATLwXGJvBlSFtP3JvMxBwdgWf3TRV0dW66PKVqIZvlr9VGR60GPWeY9Za/rR6ask
401wX4hqd1orsTSX8XjqFMN7vYsOYHfE1uKrOBy/Yatz2xfKsTk9kigJL+mS7LVL
15rRpiwjRINRDT1vrRyZj56SdjVQU4ndX53zONPU8oCDbm1w1qRAFJRUWwouh+7W
jqlfm1J+INS2nedPhi8xvTqE8fKvAuOkvzAHLzWap9F8X+VRRlhQWYDAnXU2JQ8p
8ICv8REglVMbCSvR5S8NuwTnSNSBN/U25MvLili2LVwkWqYGUaqo75IASGIL3hHN
CHxuGlinSa+wFsb47yKwXyyIgofFNvr9yRQSic/4eGgXRGO/RQ35Z00SU/PzxSWS
MyI1h6JqftE8q3JdSwkG+ozsRDga5eX9QAUduvQHRbdrA+6rI8rFgRxbllcqyeN7
MqAYZc1mqe+T2X3+G/qImNfu4zfMFYWxTTBvrcW0IcqqY6BwNUB925pLS/ZisG6o
a+8e/22gP0NwQ7xFEL7LhROUPbCxrfdce9ezefCH3osjVjzIBpFQgt96s8CQD9kS
YXA6WuVNdjuMCo47eXcdcoTDwrPNugt3pLA7ee8bhgnGiVgwro2UmWa6hr0+8ba2
xGKauEzOMPdKyB4W0L+pWq+P/ZOrBtclPbkisgMfc7rZP01y0bN1gnQFDbCdaOcI
nwtnoA2aSekKfrvGLl3XUlzER6fBxkOkrkyI7/ThbmhqwuwbslFD5EM86z42bY/v
JrCH6OPaoFZ/PhzNVR1FOqKcEv6WtSJF8AeF/mxSDel9/mf5EkoTrtc9e8O8tZ6u
c3+luEEn0IKs+7TktA8wOr/iqwVJ1TRQ+IjuntkhLwuf4qy1NJjnbeKgDCVnFvwO
1ccDX9j1AxAzGbMks9axQEkto/+qwjGzoW2To5X651ShX+tuB0iO4nU3GBDVM6Vz
fYjoyaSOt/1N3GBDjrMK0VGPLsnoSskMT8TX5AKUsNlVCPkaNBFavgn2egbt7EHc
bgp24jUewJ4nfOPLhVy6B1GngSYE1UB+SuMOwVvdXsU5v6Jhbdkz89oCLglWglVo
gKFWRcvTf1NzICVqW92sbAU2RN+z/vwt0wKswh+TjB0SdBx+4fuslUq28Li6zDOi
QI+28PeStysDPHf4kHCeAAkCarK/VFVRjBoVqtDrYWwlnidg5uq0mWTfWLJ/IqdV
RmxyCgyAYT1oBlHwFmmEk46U8cxcppm19Lw4/ZqyZOTfhX20z0Dy5ihj8VzqNCJz
4zGUiY4DUzAkMZWZUzH1DMRjcf6iyP6eOysRX+9VgkarX02iAtFRUwy0T+FjrN1A
gDg7aErDhiYNLGAh7PRDrjTMcGrzNEqpaYtGIyHnS9im8v2V00N1OIa5uGBy2eUf
Iqi6lsVeeIu7iyFCeCRo8jy6WrsaRMA2V2/2rdfmTf3q9A+zYzpkV/ev8Qm2wnML
CiXIyHqExmuhzmZbu0odV3zGhQY4+nKNlyNl83ue9NBpG2lMWZWWmJQZX8U+ysrs
qxi8NKlStcn63xrf50qe/GCAQeNdHThJUQxt8j2AtVvMi27b0mgIDN3MuCuutv3r
0Ib7h5+DcGV+NAQdYcRlx3HsmpTetEF6bt7rejFyT8vomhh+PUzXq8Ryec9fP7XT
KjFxly97U2xjl/ZvuSYOrl2br4T37q55kfKx+fczyrbW0wMu/y3X6V2LEXAQNPa+
diI/HmQyW0MiBQmA31PSFmQw2Z5ZmTGFRFSftq/UM10MEdxxFnRfFKCGEAKTNfxE
KhKD4TA9TjQlECCOQmsffCMMetDN9iqbsS9YwPlrs70zluR9Zs0jbYsY9WOHuSvG
jZhNU2rX78A+41ALYm3Hh0pmEypi35NXoRUUt8PQz1X05/RLwy1oel7o4MtvnOXl
KcWbSIl1f9MPcCBbJrclvpyIDodPNiSOGOn6OJq0bc87QdMretuZgOHbhnXYys/1
vjslmSvhfn83CG6fVqytT9qPtrC+1gFacXZHDl8ohVvYkSMs3ghbv8ai0Oyj4tTR
pMWMFBrlLJIHwq1v4MGqvM49geXWHP4k9wpaAxsUyN9alGXCubmHZwsCyiS59F6R
5vvfp+mlqa6LMuVFx4k4e130GLHUaBiIp4d+NjBo2nznwtrz69UwJKNO0ybPnybm
ZPLkVwl2qVoP4hMfU7CjCJmSvk1AwUNUoGFmLLEsfTnB+KvlhHdO9Ypu1eXr/q7s
8WlSyWChCELwngfloZ8N8GkvTLbdOHt9Igm+jrvDZTlkj2cVGGiz4AX++xV2lZU/
6AL7P4KYfP7VUHZDFuQy/ZKkVy+NKDUfmQVg4ieiCvKdGkZJC9wCwZ3iOtDBXsY6
gK8tPwoFK1itTodEP3g8dZhwCjfuOI8bnjIWQlt90U9jw7TGUNcW1lgaplQ26B/D
WkLWKPjse/OtjWnDiovK//XYsIfizGu/jN7ut5ypwCY=
`protect END_PROTECTED
