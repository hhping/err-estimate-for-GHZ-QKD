`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJ7wecg9sSdnfsDoYsZf6z4MCjJZWzU7nmuu9onHtykP15afz4QhoNdfD9ShHXF8
h8EsBwjirrWp9Dvu/81I7StVnQtMu+nicXdXEnc5LE5FHxYuBxozDxOH+AOnuZJq
JRXBSiTWlzLy4XKLMCrFp5hxR/izWmGmR2/KzuEchGGAMWIWar9av/Uvmshu2siE
qna54hWFugjsIQrQncBXbvlHonQJcNeoOjph3fJwxSFRKoaWwiycxH+HWt0xGRfY
byyIKfB4+zk98Oulx1ETz4cS0y4IaRczsBMwivj1BiyYS2BaRfTEcTL9GCLuqdZd
J7cU67ICT02m8YBGinfKIH8aqMSyRNlCzL9BoAzw0WWFGGfxMwEeknja50iWIL7Q
Hm+Z4rnCAqrHNeSE0crCIlfblMxkROwqoVoH36pyKvkBhHjPXCaZ4L9m8lj5vu04
VJs5FJKeGEwAqWSJDpuOo7yA/W/QEWo//Wvv3Z0p//miLOTQECIv5Xm+mtm4Fwhj
G5+nU3ZsSz3mWqtEVraG9K79wFc+8VeEW57Qp9hQDnUXGEEVjyhwzDLl6BOCYUZT
gZMyKEjQwo6mSw8nmoR5UA3o4i5KJVg0Win2dvkTNsoC6ngbpRaYGrQyny2gaZ4i
58UbWeFQ7nlNfBSPx/PvJnh2eO1twfntXAA5Mdj7lG7nTw7wxpAK/rHTL3zV/u1R
4VTgHa5VFvRXxOd5Jdsj6Y64Dz9CaawwavISnphjUzWvNQsgIJjZUHcDgcD42V3X
fl4nx4E8eVbOD6GKXCN/nti6JogfiTaBjBAE5F9EJuXdLrW5cs6AhTLZQl0UEuDi
clDieJ81DSUIhNvSJvmVxVY3+dw3jqb8t+fGVIogYfVs3DDyf/IVq1E1lS5YF755
8MuyIiEMuyH7dLTkrmjkRwed7+/44lvPFgtPWynldIu6h0j1nmRt33QwmnonXdoI
dM6w1By/PAHDJQmU1CgrG/usYyza3HIamMkjW/6RkFQL8wxoFpEAcyZeBko2d0p1
QZt28SH8U45btY2bhjwetJBZCYrw6JF8nPfCa1qcT+/Cn7zgx7gMNg8subeIydZs
ao/78AmSvhstMiqvpCpsTJgzNDUiai0AwoyZtKKcXSgnOI5pNk8OtD8uSmOgLDZX
4fZHSbMp6vCasK+g8Ij/YEwi87BwmSQElvpUJiBF+TK44JKltrAeSR7vy1krDG7b
rT/f6NgQJWoD8yYLIUzGT21kn9ohrK//3AZTIqsjDJutawytiIVi2OeHwVd8w3ft
6ErMJNswY1/S2DlgS6A74KPuzjnt/noPHMYmniixUWqFkm3hvheSsxaGV71IpAqr
T07mAXAcpTLFdQGLAbNJ9B5pd/VTyDRLxvvUQlD5FHpuGrLIook7WxSO8ftwisK3
n6nIB8azNLLY/sGTjII+WUT/AQ476Ewc0ZjeS+Igncn4y+N0Y8dXm2TwvyUm4awq
bWPYbSIfItcpSJCH14AfTQtV+XY+veSGVc4i7gNe2AGFvYOc9yzyadVXKiNTzx5V
l+AqbA0aYKtmXbAKJFLw8VN8FPTyEAl8oE7vWXtoHshuw5xrurR8Dskx8xMNQiZM
241VVlGVcxmZ8XSntEz9ERmIeez/k3n5kgYEq2AGXttnQVv4V4p4kEdP9BFR7Cr+
pTTK6sXwjaCrYDEwkf02tJwisEX5fQ7ZDZX2EI6v2+RrX8rvLUrYJHjG1AbEZ21N
FXNHGY59nUJIrLymcnfQAPp7nWibOWifA7dE33nlUqOV29z41jg0m7npvl+FC3EK
fO4L7M3AvfjWuejoDp8wRPH+7wE8bP9CDV9mr5Jr14wTcQIGI/3QsSK97SDjBrnT
ivkFQ7v9Igg7wGa7hFGb9/iBEsrW6hZ0hjgIzYrkYTlpoe5uiH19u2S3qrPvd91r
d58rpYG3N/zZcZTdZhPlip6yD0HugJmAd33kTQ1/HDEX8xrJYXynDxkD1G/+l36S
nXrlcVuhqN2MBtasnE4DUYKx8MUgaedFs7FP8yCE0JmdCrYIvwke8PBX3/mRolge
etN2i/F6YMznCozeDyVKI2DX04/LN0ARupG1KLzHsk7tWXXuy2gRD4Gc3vzUUSlF
4EdXHgXLjTO+aFEeT0v25NIgG8YQdUhUWzKXBI9rKWMe+ExbZNi9WFs/ZslMSVzI
UWXuyWYjbXiK9qMNhT7IQ3LVmXdoLj8z/yVSqH8Dp8pytYkngsRN5tamPxElEe0z
HSqRs55HuzJszpvMoNSMDUC0iXDtytBsVGufZUrdek4jbZ82n3AqCuFCf05FGLaQ
Fj7E3HDz1o9/wY3OAnfd4w0+T4wq23XlW5DQcVr6dr5fDg9SbxCChXs7x8W9QAER
QH5BfIjidI7PvA6XX4r6VxZarylWW2JWwStPBm5Qpi1uabWLWNl2KcJkY96xmx5M
QpuBoWCGybKTotKrKaHY34HEDDS6dTIpo2GwTI/EyhMwV2YaI+6lE6bwS6TFiVXB
ma3pU4Ytn+DTs1TQjl/8+CHl34hYTch9wTc/Jf3XbXasWfGVmkNPvSZfZBVfmKwC
i/g1rMHXBoVRjzTRc03JWUi62R1J0T3qmeX3sk++FpJAFt+l5nrOgx1DNOKHqtSC
UhsOhHVrtblvy04ADUOd9uh7t5WARLOlAwGAGjSPRISahljN3rzbhjDovEgAPL5/
Qj1PZMbDFZlFMDMxW62KptQA7rOhgTGysWQN39NKrXPFkiAWSy5FdVGG+01lADAP
czU5VNYsFlh9bUMMLuEGWNn5Y1hXM33SSvM9Ds3h1ibVBkSznA3LOllwe+UA10df
L5gPzlJkA/GwKkUlNU1oJAnlBGRdc8AsZFEjV/Wc1RQq4RvDXG7Q9JuUyDp3IK4K
ya8SjsRvvf//qzcw96IRRyMy5OOc+Si/reIdEPeTkzIZ95itgr3zaa4tJjv5uh5I
XpcgJ8mzU1YM0BeIQx6xTWTJzb62GbuiW7KWZKU9jum5Jn6ngR3wx5jKSSxYnBWg
Prfs7hcxqVW3h6oS0YrtfFByVnifzo1sjnBOpMUO6eewrp5FkerDlyi9r9F9eEdw
fr51wWXY2HoZdkkhO7st6pelDlaMNyszNmWJDsvRPDWZFAA83SZ/gAO3gMkAFXRb
6X8BaE4YgD5/8hLFUxuv+3nkeNdK/NDshrGIYyEfWf1bxzg0Sbo0lkUal9nvTWnf
adT8xtD3iVbVWIvZiqROivdoS7ImMY77K3S0sN6NpwApQLzvrDhbNvZFEBVjLs1x
v/Da7HZKMCFG5CzqDDO6PRirxxFR2NuXTzRskeFXVvg=
`protect END_PROTECTED
