`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fMzjsDhBcPbrsKlRtzNrMNlVB7NcWBReGb0RRPemx7sYkk18i8YVJLDTdF/SQx7b
Ea5uMFO5nEeLPVmarG9Rv2KAK1EyWvv3blWOiEz1zeJegSKbDqNNKGSgV8Ti1D7E
plQ2n5/oeynSdGgWpROWbRwVSoBEzFn8eQzXwxHNEuWYltn4YmBltow/fjyRpm69
K7PQe7q3/+RDL6W57zwopVeYSzpm5Y0Y3rZr/rtRBr9ikVRju8DJA2/E8cGeY2S/
79b1j0kuRQGXgqU6pGOXmce2D27fbV9nzTOaD71Nfcn0ZEEC/u8uRyufpXsOf4gD
jdhxQRBbcVZypg/r90fzRBqJbr/brmIbUnL3aciBVX8Gsa2w+roj4HcCwc2WUGom
W36ZPUxTI2UZ1hR16oLD0uduVBS0D/jD1gY64RY01SgNXj0xVlFiLPhl7boRwdHF
pfL627dqAxAWgvI/8GUvelTUxspPcv3o2OIhuFXyaAhcZC1XlgYB1UWatuk1i6dV
ytfz1EAtxoUuBHvRCG7hVI1CWVcFwrbuk9x+qMdWcoIfgv3Op2QU0IJbYAKID4E2
RbAV3ORWpri8S3HUoo2DxaBebWlz35tiMrY3gkAWp34QaQVNGRBiHruDTmK/UBpU
stpGuQcn8BddGYLDsu5jTRV9U1QLRPKA+YZ+TCPmKCBA/tHL1YOZ/ZmIo9CZxlS+
KB9SLBuxd7glQRi4APqjlRQj5Dk/7ptcvG6fZeSN4aROVzlgF7SHsSnGnVvhqqaw
C9d1bH3WfHwZ/W/VyOYY1BzxFiOuis642JC4b+B/4BK2Vi2hA+1GIN1E1XLRXRJP
q8/T2giw5z8p5ek3QXDQQOWaJ15ZxGblH/7sJkpZQ0g1TnOIzwLSqoXV4+I7eokl
oX+csICOJAhsmec5r2xjN/Cpwe0RgSTi9elHZCPr7t8fJJBkL2Q66ZA7g3LZ7krf
2DZB/Qw0ShNgoZ1sGePLIzwBXCBCYRMJ4gRX8I7qQ1RmEsmv9P+hAFHtDF2LlDGT
RmUl7CoKtSgMVSVmE6JAlPtWJBdc95CiHnjydNqgVlUfiktiNn1yhsV07KP4J/kP
PBKAYm83ARB6AVmjUo/5OkwEi3LR2O4b/Me3us267TKZkuPP2Rg4Q4mgIEjnfIdH
YXEn87ckQB27lXDlp8EwLqtYIYL4qBmer/Zmi58BmO4H+NWnhFV1gI45Tbi7HWjG
mrErgH74Hzsr16Gs1Nix1z8wBlUF8+UTPZZ7fhojudy/MRRr8WP6omguo8uothQJ
NMeyJmmGWJotegJ3iE5vy/2Ec9Y7SiTFNVEwfLa+GnF+xFjXAtjeywKbxCjuRKtT
wGZ7kEc87R1ObPll3yGtO//5cFtbc2yTb5ojdWmmDyYJ1UcRjaRGcE3pdEX+A/FE
/rgcnYkTYxsR65GVtbpy4ySAIrpMPqrQq3+SGOzlFokL/Q3j/Y91T74V99QW8j0f
5ydCFnOohw7S499u9NT9kBsbmWduMCr2qeinbHYsuuOKNwjz3RtAwn+BEWNugvjb
zV33TVgrs2ZWwsLHtvKBhG1O86JDC3gRAPlYVAqJzz8X3ll6kyV7f4CsMllKnIlm
jblK6/1RXeXXdQiZpKak3hAdZCxFausJAXdwp9weW69lKIdVhelbieAL/1YuagC/
03xWBxEi0uZqlJg1peU/aGcg61vBcQMDPGXcBLFwPtleBjareYoyeDKcTMph/mhv
B39uH5oAk/9LSR56aFNKN1YY3XWlxjcozrG8ln5pfvU0AWdpcHSaOGR/+/bDFSdx
uKDZkSXA3GleN/4GPFf7Wq++wP0wkOpaDAbDOB8T0E4RxpazELBxcdUPSGnt4FwF
rtcIWNwg3W4IdBZgBj12lYamPYJ4u/7RRgxx9lDQT5ErCG0P7VcDj41RF8lpx0EG
pL2E8Y1s0Xob79KnHM5cYVyN1ZZ24XpfKijTHxw+dUqRU5tba9Xs7QQEjGimF5AQ
tGJ60j5rd6w9NjVOyOKbAr+hNt78QkfN4EBOAuCiHU64wg3tY+O0PmlG+2GW72t3
tXLKhjYMa1+qZ8LLNjO5pZaTQZmVlhn4I5t1p/wck75LZOEXQN00zdY/zI+AAblY
cWbU1zOPiBiKb32J0xhwS3uCs6q0FfeYUDsff41R3ArdQBhK5H/PzWBK+SHZz5iC
ENW58Rj+IvnJwzP161WDzC5MW3cJYkAtRXOV/I2qtSTyvYW25PVa27Dj2it7BHgy
bM9LogUGio6JXZF+drdEo4dcAe9OvH0kEfVT5UJSycDSQo7cnfepmDZAxvPLwk9K
Wcx1WHK4ONzbioom4PRlenxoiUHn0kfr25r0UuJmjKwXmYEwbABT3Z9Rok6nNTMT
jYqZN1XZmqOwtiGG5233UZMXQ3e70zwS28+4PWWaowpvVQLqS5nbpflLGJAWnA/q
rob9xGDDykjUrscMOln+CmK54jtbMSOyWtxHr5wkpgnSgHOiGTlSHk4GgnVpaud5
DhwnwSn2wuF9dw+nXUfrBZF+zoTrSvnaduZlLcb9TaC4vcirkuIooa+8M0TqL9tp
5GrgXNvEFI1HADQT9vOsENqwQsu2kURVQ4xeiqCQgmNolnc/dwcxvnuPcgknWAM9
rnNUso2n3bQCA9L8GhV02T6LT0bsH2cRg0UdEQ/EconShblmJnq8HrBRqw7LytMo
TLgNZJAMomFeg9CpiRdmepGDh7arghDRpVVuiSPxvQ5UIZYOYxz2ij+bMRa8xp8/
FSe4SvyUGmydqt2jnzRSk4M0bjyJ7IlrOskAJQiOFNix0aLO29hl22DALSpm9b2o
UfJshjb8v/vOWwsIQcvJcugTTCu4H6eowIR6nQPsC/BS8nD6a7MQPHHKT2vxAgFf
8F1ECnpV39ZN9zIKPq4Gf8UUEEOYw8x37tirWlK9j0dwPV5A/UTU3vl3mSRYKnSB
wiGHsczBBlqdxznIkD5cCzpOE5f24fOMokOYlEYtUrAlB4554HlXXRFb6xm116xu
K0UMAvCiS/LRfcFXmRlX4eY+dOFSi5bVBnJ3lZIp2/BmdGE81BbW6r8BB4dWDPqd
4CSnLfG0idpUutFxoTT1Zd3Np2KN7FF9GQLjJFUSBW6yWuxvgJGeUNU6BJVAxyWz
n/QvQSqMa0L/Gxe+h10t9bO9G3hAdRiUdTtf8JNBr3wR9ELSsppboe0pHTdvxupe
vdph/DYsBAMyoCFEbdAYKEiLDEN8g6paPAILEacnZkX2LRTJaSkKa5ZJmneZrzco
CXbdRkxsQxWVfmQxhESUK6+uF//iV/qhVfWGwEk9tIfpizwq2Hn7+k4hsO9SKKYv
mIWOFtcW+VxMXqE1uV+nL3z7vPXKfy7vrGd9Stw49kjKfJutw6RMLwZWmCYL/Kx+
`protect END_PROTECTED
