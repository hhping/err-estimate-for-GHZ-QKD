`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpKUn0BW91pjHZYzU3UZOPdYP8x+/d1Zsvbh4sYdNRjEdkE0KcZYOQXHB6st7v7K
LEazQrKDY+wQ4pzpXgR1UGF/jvxChYIeGeCD/+1teHAZdtCcsCo0Q+/BvYjbA8mJ
N1ngFacjrnJ8gxeLxBhYKz/JdNLlcBMhINJKOr/BhfwIgRi5dQGVBRGvSmftrUAV
YOed+um1Ai2Q87tS3uUF0Wig9XKhTZ5j8iK0j6ZcTpTJoyphYr+wXN7N+fcT7RJH
q+UY8s+mrOGjIKVZ6oXG8gU40jJeDnp6KfBmmBMdJjVeVwHOnC8d8RmVBKNiHL5b
tiUBtuPsDr7MrwZoA0cKiPqwwd4jzPLvt92Z0p8Ur0TAFURrWoN5zT+v6jV/+tR5
KauCJsfPXyW0YNpnwNxejpT/Jjg+fW2+azXCTtbcA529Bh6EgawhI2oTXw/uhO/j
PDPhkPncYisW7SUoCHnjB42kvLEmbygRxaaPn/JpJi0dLYXux2sSR96jihPKuuKp
ZVMTAGWWAey5Mbtnj6W81MZVgWTvYbPf6a8P7tZKh+XIryLba5xmocq1NThCY/Cy
XfWkETGg5ZMGvur2/zc2MFnIQsLCKbX+91dzt1KJk2dCGjEtAw/YIdl4Jf8ytX8h
1nfOYBzHoeHArJVql0xvhb5N8+uUevg2xnLmu9VVtKkpPbAW2xO80ED9AKZgn3Ji
y7q/RiGJzAyyTF87K9q7sckihhw9qUSWiRCaT4DupNlsKvirefyVfyeDh7kLmAq2
khM6MpDrqUAGJL/yVNYkuqCNCURJIXgHg5Rg7f+SvxFsEFLGt0ZvFw9x8RDkvrUI
GscDfEOu4nj3r2Lte2EFuup7t3bRm0TFgSn3LkZhALU6z4DO5pZNOOfN8EAw5lWe
WGqUQxQ0r+Bw2BaExusASUHoboCwl2ofNSxy4lyjpjMjdWQs/Ti881WlIbrxQzLd
lL3EAkml4Z3lYfVGt4gpUyxBHOvR0kAECi2InIPAzLkO+P+DVY+ki9D9qYQdBZcm
p9g3oWWs8PUjosODIK8kFZDoL3Cb+xuQg5yBzp9HBu7tTxzzT9O/SI7aAwOBkuzT
grgJxZfz+EQwTKKUr7LUJeBIkoYRrnc4SvrtxLvtwsjyBbFufzQinBPZIvMHrPQ5
Cf9GwYcZdRb3PAX6c1V4BQEfSIDHjGwKlAp/zXNf1xfHyfk+2Ac0xsZeoqr5TDrC
Jn6K2bgltASFSm81bJawU7tmaP2+wIU849t8qqOZpastaA4KjY6Cnyyb9TBd88QD
J4lUeTI9W6LSYXvWEv0qWYSlN6ZblcY5VN5VI4YezUlzLzx2PevcV6DLPxwdaS5V
D8qO3yDfYr7ajsIA7H1dsj6HJsz97WDQ9Ue6K9JJno0iuIdA2KwZoNzKCMXtHZmo
S8nupdBUZtjj+/q/GzkW+tHOvI255rCpLhG3C1qPdjO8bT3Y78SNVTl6te9yNXzB
Cx5oZuRj/w7CeS9MTyfOljUXcofxaTgnMevQOv9uthxxYjEoxw4bjVVOAEUKTarp
imfMxxxu9MZ/p64bleZ/1Ufh9V8iQBGTObQjdmrQ6VZf7xzG0j/dNo37bKWiIo08
1kwaiEBQjxBOQrP5Zt4lOXveBUDCTsicU+0p/TnFV40gd2ibPUKx8pcdVFKnGcj9
`protect END_PROTECTED
