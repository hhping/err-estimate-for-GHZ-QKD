`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BuRoFLIdUNVNTSuD0HIOpWrt5z8L/2hlDi12bicVTVbScEJApsi4yjLMNT0utiXE
bs6s/SSYBKt8s9h7VNqaoZz7s68jfCDb5D/cta5T6E82+TNvLjXUyn57H1g25DQ8
LBM3CpxyoA9ZwQazXeGgnqKNIeebFZb0FwLy0JhfAsYJA1lN/YGmNv5ojhB+wTTh
BkQ2wI+EZ5MbBBhsM9d+i6sIDvmR/UrIB/Ft1xSFrvxiuC60ujS+D05vuj9uqM/c
HENG4N0bN+awBdGaPNYGKLvClbkhk5DFEj25SaTja5FrzzK5L232KNz7qYKcmcB2
ajr7aQLcyq8N0THrYuR00o4BsgL6UgsI0k6ZGr+CEjxyvZdOin6+/7WlpbUzMEbg
g62E+rMbKq19IyAdijHSf8173x0SrQc3tO2Xxrl1uart4M4xT9G2/D8J0WIQDZoc
D559Wywo89E7qNCJ+RgHgvSJ6R6L3cfjIKpc8fyLNzsrZ3h/J2A17Lo8YixDCqsE
HzfdGJRDX4aeLDK/Br6Ky4spV/x7oEwvcykE5RLr45B2HfqmWFAWGjkqpEnVnn4R
QuTEbpovNxlBCaz/Kxi/7WVST3qdU4fG/O10UiR/fleCG9wgz1VXmEd1ojrBUCvc
BF4mKme/D1Dcjv9XOX7KNy2VDfuvnr4rZ6r3vJQNCeV8V85fZmF+5WtpsfaxGJpT
NHc2gMKHlYbTohWw4TotmKkJq3Cr90bnRbPfRi4HBrzN5u2EV863D0Srae3U6iFe
WzekHD0uKluSwg8vlBu/8YDhE1LMtidMjQVfTCpPDMWJKcrj05hgUB9CH3a9nOXu
YCw3nkW57+L6pV9MTggdG75R2zOsiIED5Xp3EzneExboArk4MIqm5cmgaKdkNfzm
iWHeiVpUnBvrzgRFlcspXGZGMeR8z+30aKEDOPadX6hoo94Rm88vdVXv4cdNyHU+
VIS1K0VkYsWjEhUGEQfRss69Jv09Z/PcRIgE9Bjtpiph0g5DJsdgirolS6E3B+df
4LZdKEQrxgk1M5CancYmJk7HXrY0fYNFlQqgYbTxzSBM1CVMfwL2vIWldZZPnTBu
yNYG3XGar3SYwCB1kIEhBCM5H+PgCzTSJgDbLG8DO4a2OiAjW5g+qdXh4mBLevSs
SwPCCvHXkcWmgMQ8NF024HazrWpKK6gU0+CVJFaM+OdBzkc74lh9Nkdcr4T87sLy
SxDDubM+ZJYGKKZoY8MJbjVNppw9QHPs7ouLGiATPHsdcUP3/9tkiSP8SH6ED59y
ZcZ4cVrIC5JaWaClwAzr3poYQ9xBVDaiWRcJ7cHxXQFWIz+7r5RhWS6APjCl7xTF
ZvyQf+rYkYwrc3ikHLrct41tJF/CEXDnZqVat8VLG4dphqaNywHD9couU2qTYtxd
ZijfVq008mOMkcqJSVlES0KFu+hGiIjxerC42Xaa5VNSd1NU1corbNGgdaCgeyoC
PbpUCw19iJ/DO0WOyhDAHfzWuwD3ChStkPxqERE7DFpotOjDPQnjw6ehevKB7JZi
xYiQObvgnQmcyGKMlToG2/YkU2xIR2nDvBg7fIqEel8qRcc6Hr84hUAs8Ybw79KB
/5FTKtPU4Sw4Gvhlz1zoP80Qj0zQhe35TQ5Ad+jtfQjToRiAbzhXkm8Ap9IhX0jg
GPp1hrmh8jYdKqVwi02eUBL7KlK+0e9sOsL8spd++z12BJci71eWZdjewhLdXI96
CkaPJevWAY+Y5bJGA3rB1L/83MOTh908aRCbj0t8S5El1pjCsOExUH5Elnp6zz44
nxRzahSuyy3ZFoyymek8cPzCPeP7+R4u6xUPj3TeG2puzfN3mI+I6+9JdEjJ5xlN
RQLM7v1cvz7oi6eG+n48BVA1anNwqPUtsaaMDFgAaY/UOhxjeZVFNd1crZE7WtM/
7+FYbVVQk7zSrmh8a4ErkTpDhL41/KQnSH6P753HuZNGcw5YhB8uVMDsduHwChbs
lwA5GGLVgPxZzeOQ2ivCz/D7YVMeUIFviSkR5fp2Fd64+ra4edvdQpPIXXkc0WFC
0XRHX+BlPsgqYMb5WrRux9Ybclt3uDDQPDGHbakrAorAYOjkGM3NMPHdAevE+DcY
URBRQjxOFpFR5UXXD8ArXxlee+w968qdqBdIEwCNGSlg8y75d3A7JjCHI6chfoTI
w53w/tLVHS44SPE5eDDjDFeRa2Jf5Z3wBsXSXBT8nfMLlDl+Zw7F/r44D22M2T2T
AZOVOy96wSAGa5gVmMNURKt3pwzqAPAG+xPvOxLsa074oAbr4sDmDNW4cNaKbisH
nGbVla2cdcX/JH92c8KGEY7bb2H7lteP5iujatLx4I6WPRsIdlY99fPx20c/8GZX
AgCRe7AnhLeI4aUviQ+gIP12WjHatT91Yf1w+e4I+w2A6mic5BoPt8naRqXUwhil
C8LrirCoNAHBBljF5XX+0phiz0cr+KrKjewsq01HvCSnsLq7DLxagXxrrzm1ve9h
HgugCNB63wI5xf5JXgF1ruuTKdF0ksPY0t1wBlJqbvs4a4cfebfHD77zNELWm9EP
TejCByv2c6A1Y1gclrdUGNuS1kI/ORsQEIyu1Wazp0TV0fzoONOVNN5t/7DKRZec
aDC11wxUsASMJ/ZbVV2Rc1yHCfzB3oSMQhWbo7gHDANs64/tPc3zn3nKOaJ8x/zQ
`protect END_PROTECTED
