`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hmsrBf0CdTH0MZa37yyx6uzmg3TK9ZY/ffdmRp4W+9MaqyXZLjQVNTvDxU4fhHIL
s0jOxx2nu9mybb3oB23gLYHmFeRz4nMKs6GSlH+QH7T8jLPdFZSIYb8RYXvWut7F
1FogjEa5t+Y0gyrIx638oRAgxUncOmDVBC4cC7OhRQrqWe/PCeth7qNBcaPsqzLS
3/TYG2a3PnbnrbW3zLqPNd68Fvkq43XeVM4bzhpfw0+gtxmZI+Zz6tBxJ30ofZst
2goWXzyQU0YHonWEsc78nG57V/U2VYuYJ/NA5QhLwW0bB8dgGvPTwL6Rl2ImDc/N
saQWcY/DTyvzs4TuwSDN0pT68vVJl/UbL1v0Eezh+Vzt8xERc+6ztVuhKcXhk4E9
t994Tkys5B+Ca0OqHhNjlkwvZ8qg8sSo4bkS1APNHrSvYAEvzlWk/7Ng2KhIFCXu
Bo4/5s87R/ozl6rlWjgO+g8ehhRIABwlQaHwgaFXHrFakkLiXbD8hEfJKPZEV7v/
OWLR10d3t0uY3bT+oNqFBi5pOyLv2VseTjq6oDG7ZPlD4UJAqKbNcrVZupP5nelO
4KVjZqdgAmpB5tBMn5uq8YLPmvisx12HQOR9cNmV9ZNEkHUZMWg/7yicJ56GVWR6
FdfwGVyMJ8V5EXkkj8UJWlO+0/FJaPw00oAT9YvvlZTHSRo0czqWhP7TMJNsKb6r
+F36vXztBIm1CfWc0jxvuy4BJRt0e8TiHzIiSBg5sy+qhXypkKK3gLe1wYg9EQ0a
8ibP/7oOugIid36msTORwT4lbOtxJ13pns4sGkny9JFaX0Gzzy+JPZ5y2eZKWF3L
p6DQTbN12bnyZQPFfRTsico9x0+d7EAL2FHHzdOqFNkYjmZb9jDiUZq0u5ew6QHL
d8rCdLkg2dNOFq/guPtFOIzWGCpSRdaVv0Gy9SOyKIr2JI6Uo1MjHcb69tNJDr0I
vZPgel91UYhasfq1vqaGPp0iSYK++P3mN4IhfblgvuSS1Syfu+jZ1V4/WoO0tlm7
7y+44LXFEdp6BWXTRDuLIx75lNoc+NAmpRfSXMBk9bv8YAbIUgWs5X97os+DsaWt
GJgR58/lk5laPgzTu7xBov/k7I3NV8dYGA9rFmDVutE2aqMvFmfBDHlC4cDXKcqv
TkccwIaO46E9Rr3QBNJtHNUEmsguZ7KqYqGwpqzAW0PWCJ51finD0YFpaYSQieIF
npVw3Xq60XNBkkml5j0cq530hmESMTI9OGPD79+grf45NNCRUWX4Mi7IJKncunBn
cvS4k3KAD/r+Br1vfosEPmX/Sg5kIPab6tNO0lZZHdDjY/kTXZf45P1nWyET5fI8
ATCQTYKiM7a4p00gUlUTV98WDFRhAhevP5kqB2uAujIpothSPiTObFOK0qVqMz/z
rYKNJGYpqP/z92+gBsBdK6mJRzqwjb1S7Xsis+YVeTIrA0D97qxmWxBGUWg0UexG
P8FlbQQ7lduV870qt0V6XCAibXwpR9rSDqsHCumleBGOZozyyJdu65Eha4avFkZi
WIAn8tyEDouZpzROysoYWmtom1+Zb4paUNf0FN9Dtaj9iCq2lgNXVWifNWx4rQ0u
xTQuu3D5q/Fvu9M5SdSY8F41TKoWMLnWXtKxytj/IxQv2zC9eCB8jKfiMMUuSeTH
ATPs9NCP80QbgjRzSpNm0Y+RbSvcz/cGdfQW9lSopqtroz0rA+syOHN0zv/d51g8
8VQLYC7C5iQfeUzwNSUHa5ouV9fOaxGsZf/n1FeId70DqFD/w7BkWMh3gE1kVUnY
wrvX6vW8KLG1WoA6aEVDL9BrqAZ+n75I7c0/HScsoD0ouo+jo0MZZh3H3DFHjGG5
IkFnK9wxIaVfzXnkacXJ4w2ZYtTWtY49WBLWy1JOcgTIdompk3d61vYaMJFftcRv
yKv5+qFpzNhenx3G9UNf80izmZPQMY4X4+e7rIn+4VLv0aNXoc7mj0TVE5fPjspx
CCYb0K/zG28NzKd1P3ZiqC7gCxE6AvgTB59Lzu/Y/FOBDsLOCr5h7z1InrptYQcy
BV5R3ReIsYaXhu5tyOreoBAqY9eL6mul90oGo4UDz9ojov0n34/+QycU9Api/cSF
52d9D/ix2Q1fmfh+AmucbAEm1tiCPTytzoX3xHxCj94UubKc9Wn0awU6T+WmBttO
2dLPqEqLfwrIWYqgxGGNkoXTsSMsFIIvfqlCN70jB962Mn4V8riRuS3NhEhdELnT
YIQAexMBaIZF/fdcGiCk1fZ/cZMc8H1SeWuuAA0ei9eCeCv4qTPfwfaxGfdwOIKw
QZQDM8k5NHrARZTFegEtuWn+O8XqtChBFn3OEGK6yoB2lJuR2KupT67sYrIVbWuk
ptohibwqsXfhQRR1P75pnp3hqC0TKwO9aofKkPYNiylSLaGfBT5DFLSFaWo81hx9
heD5nvaYCYY6zLlRc6UsyjnUa+1G1MCtjxKRC1J3KKqZjum8arFCIhSez5MM1L6Q
qLqEE7JV+0ieC4YtRF0BEkmyNuqiV2HU9wsWilq+gAw3yIbCxRQBEE4HG/LPC98a
LNRt1RACPlmhhHa0cpsKQXdMSnoaUdPHffQI61IDrYHZaPgqt90IlEKaup+rTcOC
6LilAWgdxh3KblqcnqFvvIdygEL7KvvOkfhTl8r7QXgV5trDyQ9afCb/YnvZq7am
P1jcb/kJL+0FTIEA8YAm/HqPo44I4ALf/Bg98M0q3/hU8TFGIQAY8MXkJIicP2UN
u3qV7uSHHGw9X8e73fxwDKMq7Iwoba/tsKojh44ANWRYfq2zxRHBJDAK1b5dGykS
h4/LvBMUGsV5R8kdvEQJ2hxI5RFxbPpzNeVRTwMVDBS9Ezza+AWtFOinzEiITlzi
xYB0cHgyWlLnsaFuzgSiTqTd59zYS/E/3rp7xx3XZVjiKny5/uAPduWqKY5043Um
N1l2P/y2bZD43QY1ftbkwKR9S9Z6owndE9K/NLVe0oFm9QMl+Alu/gL1o7wJPPNd
jkXNHTDbnT2TrSeSutZuitQrBHiOt8t6LVFUdhPTJED5B/TCCydY16JULbOHG9NN
zzPZ4T5QQDPbxjJ493BT/gQ638YU60JTbFc4/pIjUAAIPZddyR6pbb1kk/C0TEKP
kUUl93Pswof2wMTgp/iDLw==
`protect END_PROTECTED
