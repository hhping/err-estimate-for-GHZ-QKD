`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l4SA4KPbDtRz9DkF4KXAQy9vuG/pQ3YkbZsjDwyi/DSPGoSQyhYea6V3FW7y/hWY
zLtOkkH49O2bVp2YhTf2LKu6UhS/8HoeLUodkj5kRc1/9EOZ2edhmW7M15zLCmLj
vns/kdCnoHVFfKJwdmvfu7YTc2wS+gsk5kfjdhGe8nY=
`protect END_PROTECTED
