`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5uOxyOEJtyfAWYYNXsFfKkqXR87z7GgnA5TpuLepLteGREQ7jrEkJM1wmpqIQ++
p3kqtsbS1F75BBFPOC44vOJSpLR/Xr2nBRflwXdKznhmVQo33FrUsaRwzVMxPCw0
Mc5LcQVikLYT0fZM7xkfiwDcu9CTij4S2GkXaaRoawGZgY1xZ69aSC580rBOALCv
jkaXz0usIIEXyr03rRhoWjf/AbIOBZ1O1CSnsJrkFzstkNa5UBvWdiTV49eHxiA4
oHiCr038FDar5aWB7a6aGj/brmmOmPZuPUypVrTW0JZFH3oQxQHbJcB93NWFrh6f
aiNLwIhrfqf5vlVbUpHCDkCtfnBEau3RgrdJsLlDxnCV2PGkRBv3WxMkA0EQiIQ3
GnhGWtxsQDCLC1S/NCrmKq3dqf4xoNjjPpS/a+Psd2zJJ9y7wXSgz89pg/4DoRy1
UKglRl8fO4+RoGN/k46WFSu1ELZAHpEoBGwIP+7CRUopdsI+8CbW9bf+9bTsP6dq
pDy7CfnUrI258vCAPfDp2Lj9G3r9NH9Mnrd+yFU3gBwwG6UGU/uTiKbe2hRgYY5i
fG+lR0FN9uEW7bGJb88Q0qGsu3i0HXvhUthNBxB5HUpZAPMJoAY/lN6FzxcBzGoB
KO7SQFRUPRUjC1peoV1M++tGITFsZiQQb5kDGiphcBVJfgkz9i8CRi+mj1AryPIQ
pIjEaScbAtnfh3IAKOfskFglRTR8CR+nlyubhoBDpmjN265nnvRJW16CDJk0ByPp
N8Im/qCXWWayLp6Xqor5acMjQMIwh2lLCVVaqu0F5SSI0oIlozvaABUE90ziRKEc
rnF4G0bNGzTQtYIyN+F1DZKCFC462eUEevyhpSG0DYPjv9hFjcX3nBNil1xdWtKu
n74oJ9btSHL8NbeR3hb8/GTcvKJXYlVdN/K4xhw3LCru2aDpXxFWneKGzykPfKpt
6/C+9ORh6FrRbdexTZPVKPkH3jjwxQP4M3r2/Qg9/Z8xEKWY946cQUbWYfJU2P90
6nFKsoitF7sXb0zbcmq+eX7mGXdBC6B7L51FnPruve3M9vx+5r8cdWlJuHeZoyJO
qQb3aqEd8EVbKIIh9nADy2X3AVNh8VLBVleTSRb6gWpdOWnFwwJaK5qfYCAX2FNW
5YT9OYf/tzyKAP4onm+qNK0389l48ffTHCKuNguspeNx/6R5WLOCwGuc/D6W1ewA
xUhLOtAnU5YQfQezCVg+pjtZL7ugELj+JZpt/GUj3a2zziqsNDbh6r2lmWhek/NO
wCTteH+KZibF8cm5BaUraI8oWHLsBK42Me+mahdtQzx19do9ZKR7h+/idExBG7nR
vuUQR8NtTKOa6969JrWNYuVt2JaiNH6XYLwi5GK2Ai5wLk3FhPITHQ5oajWDF1xR
HSIcHyY/+5ivYtBH57U/xqsY7ArYwB4aozbMNOMWzoViqXOP5fbpWckgVUbfl0bi
ALls3rwy3V2qia3yVcitcAmcm2uiSsGYc44A+01e4O+21vgwYi4KE7NdMaA2U7kw
Li2GlRuS3m3KDQb1JK5sUn0qKPuW+Hroc2TvUPG+B2kNqkHk/KfuVVhln3gpyRbl
SV0sbBCJfZC1pVWh0/YAzg==
`protect END_PROTECTED
