`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmYdLYNyBDHtm8Pq5HLilVbtdDAgUzWXBSRbs+IP2Pf7TL7raI/BDsOz1s2aNnWK
TrUHbuecPK1WHsCDU8BaFepvJHbChCXZR4fOY/1xY70E3DHL0Vk+76xOWRaN7puA
+z/5wygkmmKDDrCmQyzbE09iNGq5xRk0fJzDl8xIcL229tLGftfNPx2HqMdItpQ8
K+/2l+vNPZGOXJoQlyfdiJsg6CLnRZdf4Z5ZD4/GBKTSjCI/zHUhJtad3yjhW+JP
TvpHW9awG2t1mhZH5wikcm8hx4yLw8vx5Z5KabXmAPH8sDBg1VfyUi+t/R6sDEXb
NWYqUYx3QIQw4zYSgvTU8ZDpImS4a7JLRFBO+2+ftPpR0z5N1j5uzNARNoH71UNn
ifz5HDurNI3m0YvdPUA7gcjATzmJaacW+T6On7ryGuejkxu3CdVqJ4WvA1C4QaV1
4k3P+HIOknFcf9nVGMHOmYzj22blzxBtBqSzFUP5Bdm7dBzprxShfG1Q7UdV8HWm
DRpTp3Dis1rUvisgNK/BpDjWxFaSo7aChs5f6gyZ9+CzYQe0qRCtB6q79s3RZLdn
HQGjQLr4YZ3kBgmDpuw72SWhkiPKEzJWyG9uM4eHosf8/EqfDDs2Z4R0vlsW/1gi
ahCp2tmgTsBTcAAgJQaHzSxSer742aOA83/gYGzInjBlHGJ96agl65fTg9dwEGu8
HsZ3BOWL4rycDMOny345muNBddNkR9+Er1gInetMqYZSv5RHDNPsSW16S3LEMfHx
ryWhT8Niid85FMkpueDEpaX3nvpddbkikeOxo2fxaIVihdeVA+L6LJo7f80bTYHa
C3n3X2ibITJk8UHK7wgoiKoddCB7yPGX2M6O4BsI1xDj5NwALXKAyCx8bpLAulWa
skIgDq8bW8vww4DqKjitaPwHxZEV+DveBl9+tmYgZO3CeExI3alqrBI7Bq/b9730
ELOIaIvUuVkOKl8p1bBZJqLi19vzG02UPIR/6q3bTUOTvsa2AvvaZd9om921fKd6
PWETwRbgd3iQ1WKnqIisR3fYoAm9Kqqxjmmw7zqBv746reTn4vi4j7ZDMyY0Uhrw
L/9GHcYKajdt9EbERVwmARYWYpqCi7rd0i/jireaQMGVxDvpq8u21QH/JRK8GpwG
U+QWeujzx6NisA7l0zQYCQE49/y5mnZ0XR4gFZijScbC5SJIONQrC7YU6/SSZRDK
PTR2O2mxwNyoetUmiDz2isVhNjuRK0rwenjDyGYlNJZcEjvdHLrYqV5U2J+dM0hz
OJmtP0tHLLpHs8cS5Wah1EFX2ONOH3mC2uBM73cCOq4vt05HupR7QkJY6RhHojj0
6TaJ49lDu6ret4G/yFgyF85Vibk0lWadFXyk62VxoAUMLQ5eHR/hlwj0E0R0cJFi
XxEuDN7azKMZ0zAurleIHNlxfm2tpSyUu0iTGyUMTxHqsTIfi21BkjQWqkBLwaVX
5fcACJ31iQ8NSzY2/rzE2laZcY7wt+bMLKcS8hIiPwkMgQpbNyFlTv/lCVa89YTP
iM64rEvuvck2bIkLM1pVVkLcEON6oQjNgU13M2oxtjT+Scfd+k0kuqb0USY7jkEo
ylVw0kYmJ/SiEuorMQAP/pIHPGGiul3Qh+o3qY4oQRlWdYsh7kJPFByIXBFqDhuc
MjZ8AZpvU4w8H+MztupYkKC4dot1aPdSKQJ1LEog9qTZrRW20Dlf8/q/8V5+oKHB
uZZEgBf7WGgBGEZ2eyxp+fIHijlU8DK72XL9Kd/4uFB/s3C5t4EHZKdNlG2Kg6JT
VTExBw+JX/8Fs4cBJkP8ychEUTVxfTzampwIEiN72eBZDk9B71loS7EjqYUpZPx9
KYdabBKUDvxQOVWsLLQzfKWkwLp8+FfAlm5cQf0ToVL+cgwt03yYo9GtBZIiwc2N
zFCpb9pgnGoRUf0cMyp75Z3BCi0bEUn5GazCQvVuiIONzvxFsxKxrpeKd7V/MmrR
FFGOgor11ubS2Q2X4FkU4WTUPpGM8gsgIcV25AOIIsEDuYvSnNC21n+Vd8586PvN
GUsxvwBrPP0+nW4gdFZQfIAlgKUkof4IN36Rjrkx+FV2dK3UIR0cESbeNyohtodH
KbQYb96nuggWMvn4gjk7D8GNUZr9R4L5Xc6PIqZNMNmU0L4usgjo7hshP+X2Jitp
kYAMn7+AL0EK++7z8q5hvabKOvFrkSt2ynMBR4/oaJ9o9DmjyQtcOT1AlScTd9wI
d6N4NaOQw4/xtBbzTGeTHkFj097h8eWjdPi4fItZxYsvCiJlcYuwmAYO+mmhoiR7
kjMKFGJDC5nTTUyodQzNk1Fu+YmUsTkg8psWFxmhkSBxOscvuifbf/zDlnp5hUtL
lkJVG8eh+UVIV3ltrTjIY+aSWQgVTSWIWMIXRhq3vXA4jBUQC9k35Koqo81CkZDa
UFSXHm28xPO5yBbuiV3KmR+Bzjybx6GdyBtkFmVIoTmnviJAWdez8XJKIVmJkL9c
SAMp3Os9Rwde9LhzqGJC71VwzJ3capEmi2dTkPZ3fvrc20znW8y71SFyuNAZP53z
eUdI5Cui7g4d8Fr/ozqFnyAhedGjQ9FU4ZyKrEZsjNOeoirkkjLjJxglxltUO/KD
5EQx+0J+hVC/akI0z4sgJciQ50cXAkIj3NkcEDXdZ3NUnR1Pb8c45kSRj/MkV9up
6WOZHC1cQl7klbBJ6c44c+soqJcybS9dzHnPkmaCY8o=
`protect END_PROTECTED
