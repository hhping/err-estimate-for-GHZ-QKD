`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J6k0RLr3AdGBomUTLpVapO2mNhxLLr/WANZj2SFz/zs1DysIC0v7Y3d4ygJDTVXr
V3hAHzmM3LVfa9VWqDarORse1d8W7XLPh3LCJwEr6ZqfcZu/++CL6CJ9P6lKHFHh
j6dapEY9aowBEcL/qV7tidpXyLzKv1ah3CVM2/O6VF3dupqGhYtxYLJ/wKmzk78I
Fp4P/CqWCA1Vwy5HLArfyRnLx7dFDn13Yvr4hHqfNJPzVR/deOwlPyg5z0eif3Yx
1NTlNhnoJe5Eihzt3PfrCCbufG2XPynE2dAPnKnXV1/7q68aq7kOe6jGFn1Saa8/
TThIqIjEwHKwZaH0qCiFvx7ilA+CHAlM1S5PyHc07/t3Lxv7eul26iZGfnx3A72v
xY5yiC9+YigEZUfPtIoRvoq46A8jJMju7gDDpc+7CZslBp+K0DKw3m8gIDIpwK3u
Pt8BzxpthqjfkVTeC8bxHvEsailPZSFp5AdpgPzgs+kIAx9IY/DS9Yikw382kadH
STVM0g9KCWxC0WSy2Q5Xdg==
`protect END_PROTECTED
