`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0e7JFx4w8oSPjF7xvFlOlli4zaGQtNuB3dUzgy755g3X/bw5vw2NA+0OxsBtsLF
G9GvB7kDG5OGSEAu4vrRhrOj3iOxoMB35RKb9GZorYe1NAwdg8nvJCFPAQKWvwu2
+Dm2wMowHEkapKltmeMkAL7wfxOEHzYfmriKgWqS3603iIIG0WuJN3BgH9OMxZIK
pmLSlcbygG6H5b86gO9UhBDd5mjURlWYnd57EyG00OpxgBSqLkgvUccTOMT2dDJg
ovykdAhb+HKmsoNTmYMkYqbsJccI9VW21A81YobUmQmDUJSnlgDeiKw2REIhgVRM
tPHwzAvgXu23QrqyXxAn6ZgiE49rIw66fkDyGAopWEZ3r4JOAr4zvJTb4goZLnGb
YR/qCOb7Dc/MAfXZKjJmrpZPm5Csb/i587lz7jX6dHvDgcg2DUVqQnR5BpOxytUo
xylNkbSOfKasn5L5Ct9NksqqG8m5qhMsvQ1CL13ybkV3ndPJqx3HQ+0UzDgSvYGL
EnKgqU9wgnJUbnvWRwpb+IXolfIOAd+KKygZ9/a/oTKHmeZ6mcwYGwzngJhOszPH
tN61OVCAocY8RRVKy7YKKaGRIX1Z0xkE5ZqolVJk/GdrVbBgoSQCON/mq/Ui3am5
r/9lX2S8fFByw5/cNquAPU+KspCkk/0ZcdG96qxga0gmH0L2I2uXygibhXZFzgwj
udYU4XVRFS9SWxNtGqeBFqSeFc1l0Oxp5rweLyACMAcGtds5LUe+DfTkrlomqY1i
yp+dko33IWHwtbnHPrAhPTCvpP9nTqZ28aTgFLIW9E4MExpeGnY+BVq8tFb9fB6r
0p9yt7d5luJphZiJsJWseT6zdtHF+pqy9wO9Za6+OyGqGFvFCmIryBEDGUmpN9k2
TaqDmTYnjzqhF8KPk9UzuD6KvLFySDTFZy19vRNOEhJU2YwApR7csWz7P1PCdAgz
evPgeOO/P0InzIPWiMRenEFGB1qimWyMkHyw9/0t0pg=
`protect END_PROTECTED
