`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNlzKSO4xeFktmEDqG/B/TugcAFliVhoq3Wq1XD6vxT6xKG/4QKxzEEkmZ8TvWLZ
Gtmq0lOdxcEg5c0CyT7vc3SNSzIvBZFeYowJwjNjcnjkgemJq9xNwSGQCownm97D
XJCfEbDVv5XkXV525tDJUAPBjMX40xDibRQLWVyd552l+m2cA35N93HpJZIedXpR
R54ib8xYf16aahO9d79/xX5Sa+SEvlISDVP0CalgNXKPA+EP8YSWUmDiCWywSwpf
c3nJQIcqqS+jzf0sm5f1wRMxwA+1diQtQv5ORLqB17WIBMvbR5R99DwKAv6cDjrR
pcWbMx3xg4vluAMvVUYCgKZbGOzdNd5KVTczOb/wOKHHw4IqwT1y5/3newXgpXIY
vJyQzIaGv7VQ7yXWIkFq/EMx3F0aZmO92plkUj0PIwFOLbVa6sBofgA26bVBkdrd
iGnl281yp4OlcZx4lw57wLlliA91Z4NHL4ukdbusxMAJ8JoUTPkGQkIxgjA+3hRA
poGlvpeFoZ5yyFCTCadk3zoBfNF6Lsg2Lo4QwGKDYRPv4HmKqKaxbi5YL92mx7+q
cBtttLt4XhUnK1cJdPYfYpCoH/vJHJjFbvlJKz8AwcqdA4LwJ+BwEZ/8qI5TMZei
dxvUegNjTRUEfi+80c9BryXjdwvYMHGWYTvFN5Y/s53FiWw1yaVMggf5SSQtR1LV
xjbuLYn/p0u76ZNSA1VQ+6909NAkpfwEnZme73zI5d1qxow6qvtGXom8K9TUEG/O
JBSc+lgcoX7DXXKZpX9EQMRq0Jg9kYnQvjT49HPGWmOZBuRD+LtkkgjCkdT4Rhth
WQzqcX/p8wUoNVgJbAU79nMsa+dOhmxdgafn2I0mzCZjG8OU4C7BLnIFpby9G9uy
tqiorNBo5jIbqcswmoVpdZgxAVt9LBOORToSIPnkAOPnQXlI8FxliSNprqikOR05
g4I0L2spNntk2uWF9nqb8Ry3CssXWqIxTQ5J2OMA4kdpMMsbfkG803PjzU32ONIY
tFUnxkRH/u+JPzA/ot98lGf8/n6uuxfbHOJV1weZ08g/NvClkDMRWizeKSK8i1yF
1yheVzCGQHu8lzxTun0zTGPiwET+2POICUNkwAjymZ+Xg7u2gFGFUHnWcIQllHNw
UePjLuV7SH7M1oJDkQgnQaE36C9I0xqeaMdrcKyXR7quWfXOfbIGC/xyQ7HE+37q
8YwK/fvKHqMftyu1c9Tztijpo7bw5b0kLOvJ9NWz8WM=
`protect END_PROTECTED
