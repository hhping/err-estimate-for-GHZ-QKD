`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1i9ppnnd9tOWF/3TIIWF/Zfmmj4xttkGJ+VgsWhB6f+64Q8zk41e0574n2Dwafu
RfVP+Aus2JsA06KqdH0OPLn5Ra9uHpoU2Zfaxs0P4TfQE3VmCPhlNGzSBvjTkmjT
q2yZApdXx4aNoG8C0014n8uX6/VlRqdI/xhePOjRnRi+jQl1yq69oIg0kNfpgPN+
Ob7DlXdPD3AKQ1St9tSmXyR289hAP9u82I8ID5cvXD8cXw3PqRfB08X2Y29YBUGf
ovOe7epDwfwjAfO2fqec92VPPkJ0U1YMqfHVg7Pfl7xsk0UqGISMry0FIkJk31bZ
PyvkLihySI6nuKOjNM8NZCyRfsDUY0oOsTiHgu7ibRXYh9wWwPuicnGWwRdhnpJK
C6qg+Zu/c2NFgQ+/pSV2ZBJsFcFLb4k/y9s9734LO2NL5eQt2bJhU42rns8D+ZQS
2uHjPCQLsrKwsIWizpoxEpiqJivApfeatHiRK33XnUA0TpFqM/Ms35yqTIJ/ORpj
/u9QX79YXA+im2bL+UCVlwBnAXQ3PeT4OOXTjIiF7ASWzgynIUfA1zCTCXuqtB84
sX73bCoITEKm1qh6t20wIQzMs5WHv5xhANlZjebxIjkrJjBsvxJY+9N4baRpeGQ9
GFHltSaFbRuu9shwBveUQRA8Cs5LcJ7jR2HHuL0vHCfTIWedzM2Q4ZB3Ms3nkZyq
cEk5nkY7LMu9cB98x7yH6uWGcn1DEerMAtwpgXTqHAzcYAsrJWxFcAe9nHX2XpeT
+PkJzsX9kaD/FE2ZdY0qfNL14+/awtoXo6vY7JsmZGNeUzl0dg45oyQBvuaA4nNa
NP7/8F6DEJkFJeOrqHjH6lgO3x8QPp4rM2nXp+7zTf7qCR+bnKw4mhCRsTx5QeiH
PxcVml2Nw8/BERa6qsEXuOxcvOx/AR77M+rlMkRb0dqIOCwf+Die7vJ1VA6ZmkGx
1PsT33UT+rcoC6JddiUD//swOqVD9zylBr73lA+8n6E7nHI0dV535O96Fz7jgFQt
4rVuxCCgdE6yyJpJMi/2sxe8/bwJl7Guj6wf77rDL2+uyPU54S5agCdkmujlMOzx
1rfDbI2LqaL1A5ZW7DX9JlAVloNRnKJfHhYiYdGo8DRzraJndvqMXehhSPDZnM30
Ekfke0HhUSh0MCQHIc3BMdUERchocxJ5FZ4usfFioQbawvUJM0OT2qDcCl52qPFX
uI2Xgj97s7eON3y+kJxnPlg8ddayRSlGpzpKYDYD16cOG0ctVheWpChBS/MpjdDA
oBBiuGSSBepBMoGol9sMIhs74YSSzLB0Z1UERXtItOj+N+3RCqicG+DFf3iqAAy8
fCgluzPLVatCt62cjz6ufatMWaPRSmjMAHtRWkPlF6Eqnzc0ZrC80MhhXnTcI2ru
ToBvQGcUJNotKcYshK9e7KeQcasRa+N2p/wWmwIC7KJrQrN+dF43T+tKflidc63j
2GQ4ld6If0KcQvPeammCecWthCXVVTBSwAi8THCEvO8Nsn7KOTMlJ3Rj2YnzSqdI
T4owJAummiw4Npf7Shzug+wxOGFpUjvWag5LhSSUq9HVpYmEpN6NuY9b1C0JP1N0
KWFDBGZ0Zp6iMEpbQgBBFkKMHpQWKrjs3RDKtGfkLpzn+7ijOgkRYRKdZccw+BRq
no4XRaGTyuak9UEfPkiRBj6rMSJBMqkpn5S4BBUJmWqf6RjlUTgjrOxycktbe7eC
9Sdwl09B253jfxJK+O0yA1h106ImnzlNmk4ECwvUz9nwYT6MOgqyxBsiULPOOW6s
Os4TGG2idUUL5omfHigKJ8ICH/JzKAKWfXnPewXvj8vMjQ66GBS/FSnbo7qCY3Mx
YRDiLJsdfu8L7GdBVPlfDowdW9V8fTb/2i/u2bvGA1IMHkqnLsfPsNVNTFN84tHI
F7hORgrZQOdfdCMUx+1sY6hdsEJjJkgE63937GHlmkPpDCtkJmbsQ7TaBD1v4qaC
2xgXlkrAPABWT8lIX/3sJFb3OmdxTxANmJKW7i2SRV/8+UkmydvTgu4OFjPmO8NJ
lMk07YVV5qXub+dnESaSnJYDOhIlvHKlOdcpLcrr/aOTVN6rpXTk0VW0mE0UufLB
A2lf+1p8sLFGLc/h4dgwHMsD0hR9KSuU0WPkztu+OnbJ4nuCXW32n1ec9MPMmjzH
QGf2Z+nueOzeNOM7ZANLva+yKz01QVP4iM2M7NAdk5Z+vNVxcpy058xdTy1ZnuzM
nJT1WjDGACUkcXSI/Ta3+g==
`protect END_PROTECTED
