`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O3BLaKhk/7WukmlV2JxBIUKnAWZ7urRmUkkdsqeIl9J08RPYe0yPrzCsE1GBNJXo
gWGuLYWSH+nQn5TJI0h3evi7Nd78vxUnZ5gJ1pu/2NiuIolY9JHbRB3Gpc1oCFoU
Kk3l3nos02N0SKr03VCMhgtniJ5dRt6fE5SS3qemXr11E4yt3F5Q5G18ppc5404y
a95UoYA37NCLKzsC3nyXYHH7hLHkyjOqAF9eObT8r0DB4eY9+yM+2axLAcVUlUmW
pCCxrl5TnJz5fsJb69WeC0xUvc5gePuFSt2/D4zQ8mSsASaiNuWdJKFqz+i6qCBr
eD4zVvW0dzCnf7QA/juplXjzkurRCDSWGRY+o3WAyKanVgk5xz8SdN9NqGbkX0/M
+HpoPz9lgqmANgIYEZ/oLpNnkMmk6JbYGIo9Mx2Z4hb8zdC1/D0pesyeEReUx6f+
Fqn3+uPcxMJBIcPta4QYmSjAsWTkdUqdoGhDHPSQL0TAFkWfupV+pJ019IIwNAqU
vqbtVFU/FJ1NPOk+7ACqiDP2MlMlOFJ7/JxScxxWvp6EMb5q7lkAjKRSt5TcLhrP
mO/zDGRPvI/jFQc9/B/AzA==
`protect END_PROTECTED
