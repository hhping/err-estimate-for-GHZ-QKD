`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LqyxU9RbSuoH0x5mtNskN7v9/+QOj6GLvkqXYV1UD5/Xj5mOZqYHGmE9RjsktzQ9
PfL432vFm2LNqt0zK//u2hIiQKJnCBjM2fhJMteVqXomPKBty4+2gznFrPF1ivLD
wR2DWXFf9JEPIFnxcexI8MWURCfMFo7CB6JW9oAMUQKdpOABXjJqLHKkwxCSDgJY
nkdNVjiXu5LaAMMpD68af2GpobKHGr77xjfzWl+R4B5KqHJB1WWVM2M+m+/rwPp6
0jjS++nlBiW4JjsOYXluZPwQB8i2AdhLDpD1YDruAPtmAaQK9ZnT/4mIjmbSdIYr
rwvR1DFT7RgASAYqxBoUVF4NcVTKjVkjQ1D9YPoOG9sOmRTnCU2fKRjz+IGq6tlK
nyJ6SqRGp4UYxpjaK1DU8ZVpLo6P9ZDHGeB+Po/pINczjELJ1MWFBcloG0TcLJBV
7oKbdVkRDgcyJwDom3fqazZazOHgG/yTv9EapVLowboHW1LTu++vcNl/CDna1k9h
IQhrlG3wR053j/ivgArcZOgV6oBLRchWoF7LI3UwOAyFFeuW8+3GR5QnYePzXmAd
JjW/FWjKzEIDtGZBnyLLXu7zKtrdh1TKoLYDgrKTqfw=
`protect END_PROTECTED
