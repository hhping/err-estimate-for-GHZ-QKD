`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7WzPMqSsI7pEUOMQHxKTja+djkoVAGjS3hcd2mi8m5SgrvyZdw/gX9fXEexWmWY
M4Ol1v2i+OhKqzoFpwfkj5o6zya/V1eDz83VSSUzIZ4mhAlIrVdlcWdpaac5TEJB
VX32xIzVI/PbcykpTRCQSqxLi922H1oQCDqhZbEhfu7CVMuUfLoqXNwDgVqiylHo
wDhtG3yMFZnVHZxraM4HQiQl/CdZWhHiyLDowW3bsizWiX0ALPLwvVp4awjLE6LV
tYyZu+kICQ+1cZWpVyGyugghiRzsNKPUUDch0CS4ZGYo7hmSlnKgMJPX/SYMurII
cXB9qOOCADsToqyEPlGDPVzhSrUdBr0/2QYyH0n/4T82xoCoICi0DlGa0AkNjVJD
2LAa239kNKAq6DNI7ME1fx3BlwsY4mGHjJgA8piukAyxj0KrGBih6rQwEYxr6iIr
9sDop18CDJfB0OxRBB7MP4O9YF4vHHaewHekloYH9MyBvg4RzzUvr/+syqwt3thg
vVQU167T4clZ6W/4anoewkto7o8P0K0BUPfB/NXKolfiw2x3YMnzoTQEjDyAWs2b
7vE13cDV+H6rInLeow6pi4afN0S1G8GoTrVe7GX7Ex0dI6QIhHsXsXIY3kkQWIvR
Slywld5FNamhNCoD8gERm/lvJ8VtjBSsqH6cqJannQU=
`protect END_PROTECTED
