`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tp9N//tk4S4C2hnmrLbuvnZnLMsOSjqkRoA/euhZvlrTfywK6NxxUgz3aKaIzq+z
EN+PXXMNTpHN1t4Mq4E6c8v+nVhUS4/624dgv63kyugo1bisUSh+Hxdxyb8yfPiJ
FXDq9my9E5g3nRmuW4TR/go8//T0mwPoOP9or+LL7N8pCxPvB/TA42yuAxFv/XnM
aKpa3K7eBCVdEIuw2bvLDeevOVcA8tQ0crq/nIuKwEy31/VCEe86txIdgdo3uL1L
Q8fUIXY05/YWfUa2gk3EQ2aWLZhkga2ZE9dl7Xb819HMySZ55VRsUPYSU5N9gdzb
NdPZtJueYvnzTknHeLkF445bZDBea/2yC5u9Jwx4dMiTxbW3svCxPQuhuqknsbph
uQiqGCMAzrMC3lJe0MAhjOSxxzyP1/HFQK5FOxxWYhDCca7xf5QtE7fWxEahuSw1
CkrRtwCHdztttxygv3ZUlMU/EJCMj2OV8N8qqpk4AsCYOZhqLZ7ZIStM4Cm1mTRX
5YGTt1kpbobY66fRAdSBNGGJqgFU9UVZ40aIEeyqVJmxkZAfJB+kCtItb/0UUZf9
CCY2zKfxKSMVQNGlGm9S1JvhXkj9mpfDkhAxaOTWUuyiF58zzesoD0XXwkiNBQoV
OUmOB3ZWKMOAIfLbe++C/xbudFHhT8kppt6k7kbrstc=
`protect END_PROTECTED
