`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0//fVCM1za6+Qvyb/KDXVLXfsSd2xz3FpYACB8Tb5OrWS5c05YScFb1f1c9mkI/L
rwT0aBgmUPdB95j3i0Onb+/jYgTnIj9/gyILHmwrTqiNtCMym9dG2EZuKmhhzfIs
WvN2IzcrrWf1Cu9nmFEJSP+uqs3r/XOFY/BdpeF8pwosgzFsO4djDtHyVRpEFEYj
vsKQCkacGaicY57wnrZJgA4txCFNo5N6r1iL/mpohyHE/p0S7zPLWCyG4s55EaT7
QIJVADj/p0SXuOnqKa9Ed6+hJO4g9bS1NepyZOcPvzzsZrnXo88MRZsd1ewSbjXF
XKsdqMFawWjigjnAFelv7bQTZ/wdrDwlInigXr6q7iYkvY99ijto9BILdh3jzIy7
8ShqnPC0PxIYC5a2GLDfr33P08kPmAqUyWRcSVVLyOeG5PwxWTQlUNixcWfLY3Vy
6ZI8lgkEwVnuAAgBXd0KP3KZYo0J0LeqO0LUfFocEf9wzHZzI32gbDg5QHWPW2TU
+DxoU9D2woLRVyb+d4gbx8SgeE/KWI2cYdaQQV9lDAe0uCAysAHaedPhLKJqeujm
IQ04Eb1x+YTHhghIb/sJywKoxpnplg0ZDRl/bINWrqeyA8JkbBjsiEp9E0sNWcRF
j4raGZeeLhPC4UdD6kQJXVaM+/QSRri3NYUDuV/o3LDMzKjAI4u4YJgROr9uzZyK
3VRsrSKug2rzmeVG61+nqiXvEOkqSv+aZSnBFo72JBEhBde5IalqSmgq4ndpUlgd
KPJ/iAV6w/6hHMJ6jain1APPjrddSuyLzwNHNL8DixNUNFEYbXX5+lFeqrtyuaUy
Ehe45CMEKjkEyCNDXi58tZqTNaKKcfoumaxMMz0tWmRiapDj/hHA6c/qTRgI78+P
O1XoDt205kyRlX8l7OtnNLE8CZoNJf68w7mhg/oYpqfC4j4L1DLjE0QcttP65jIZ
2pSzSdwMOK1QFtNvfK0sQQg9L3Y3GXbrUWAbljbvpCk9sKnUIZvFrERJQy+MihDG
Gu8CcR88drxrjJDsCDkD9Vqf+6wUljpvOY7WOc71sw9xXllc+1xlFYrF1qJw8Wtv
74Ik6XQ7laQgTPkWngzZOpvrBgyoeSc2kD8Wirwsc/D2fmQUM+Y00oOKuRbkEi/A
DCP6agHRNQz+RJNN1E38wqFk6jpAUFc96KUNC31GFkyroVc2gPIGZB9CMwzNol/I
VIPJbUZgacujKF5hMsCgw5tZIXOSUOBb39VfehRJH1ErBUxUGI9+Qe7/Rzamva4G
ny8Ec3ni0XRjbeTsInBdqb0ABaFbV07XWegdznYwBBxeIdC+LwFLvUM2VSBrU/tc
rx9P80xVj/jSOYPKjMOjzum7Hf5PFPvSnbJ+MZ3t17Z/hrwD2XwdiAfkk/bixqV3
aVne/VbOI0fqYgJd6HX/D+W8iK6L3JzXGfibytBr1kl4xI2ogD5JgVMYSI9mtYbv
Gk/hdR8D05fgqsER6iJHaHDIlQiHqxUkxbCTneJRKi6C71WveGVliEoFhWfxKdvp
RglDFZauM+gS/8JmF3AZgHEWZDJjcd79SpAMcTKqfS6MhI4aRaOmX1NIo5GDXmfo
iJSs+xTAFRPTNXA7NM4mndC/UljQA6IB1UlTM+dtrj2HtMb4uOILHhIwh6stx/eW
Y4k4wJMbcG/mTVBwrBciQKeIaMxKcjidnVifJwzwd/78UH+DTxaSd6F5iHs/Hx0I
mlGTk6sXiyqXh1mnKBfRfXD+SBe/AilFWMLJyiT6IHxPnv5Yc+oCIKmvlSu7jIyY
pd7+tqVJdhPl8NLlIMzaGc7JLUA+dm/WD4XjNylZmRR4jFMnWh4jpmyroiapjMZJ
spUfyf5CzlDf8ka0fp4XtFP9fFuvCjRtT2h1d+a8YMVUtq2sJ47eXu3GiheGzUZo
Ana6wybNWefbwfW0tQ4U5ImVJ3Y1myfQyzZtczyhyR0C1zbA2N8S4HwKjQkM1ZU7
iK1IeF0HQA17T+c9YGYFQEexZizfTCFSRtofj36cIoS51mMEcKOiNCw94F2DVuC1
fn8tY47K6AWRm81jdInNGLLfat7UUjjJ1sqplcRyUc9ibR9qhPVaNubYVbpOW/EX
GDbgaDLKqhvvLFdJUE11uohpKPtNf/SdWH8geZL5FUHA5DvsFOnvkGAY1MFybTk5
8+a68SHtX/mN/DrHl03xTcPOVCd5mChVddUklWvGtwrLxLN+ODWPISJzbY0sVY+f
S0j71rdDcFbfMtUGaSoM28O8wJnDu39t56gcYrxkIL/Jzq+fmmhOiGnDDxvKg5NM
Vyxl6Jvbu6NBcH/z9hs1Hv937UhqJS5bSbjeBOfiQXxsOP6u8/2LOIuT5qSowYOW
wigfQGX7ge7yLxttRXYs6RKqp3Cdo2e3NZOL1x/8PMwooZtAbBCOwJUy4qSwriK0
SjljaUw7N3FUXfSK+Q9Vh5LvR531kzzO5inp3/gBocOgfWz4yKZ8DhQO0rU1cSLm
omTHEFq5nV9/E6s8RJWI1akpmYGsYURHo07SqctZQOuYev1wZKZ0SAS9qnvVrD5g
YdOIKxW/bZYbxV/vOvR3A9Fl5Tr9Lo0s458sPSPw+KyCqf3yeLWFhrjVODvwjajc
aqcidwfJP09QfEG9UHvQmLkWM94Ieg0NSAJKSUeUqrLMvel28LS6R8IlDTkKu2rN
CAR53RrMmI0h5C5S3J5tTHpcOO3InKzxPyR6BOrhsvdtygEeW6QiUR115Knop7Uz
Fk+qTXDRoSCiOQM528YA8uxNIepFJuFq/n3NaydQWY0ocRdHbT2Yi8X54bHpmct3
9VvJWgI1xWbsyyVq2K+uazkohO2aEwXI8ngGlw/LWuJHhV7FGS7DVMtbgfiWw6kS
zVpdX+K73YZcZ/xFAyCQhWzAzddaqRg4/LgxTCkhRyfgObr5lonNpabenidx+apP
8GuFbP3ypdv8LiLXDe0OGS19DjcnOerK1l8AXqX/dRqsDzXzIAdluwQwj0zn6KMv
FdWlLsyMV3RhiC18u/ZuMIeAOfJ+KdflRBnSeIw6Woq/3cwo0BjDaCnozXxWh+yi
GhBeT6e7iVGFtEEXQlnATNT2itKqgc0LVEVkj5jAOsv2fiV3Fh6IdN7aNpSobA+v
wHCnPRr6QzdypYfyMt2lWpsdNgdu24airMVVQCxMAngWpTaSefv+VObmVeSJQHuz
MOEMBXyDQp06vY6S9MmYf+WxqjrTWBYqIQO3JJArSrxayS3eLsKyTl7t5NNcXvDC
EwV+9fuiXgA4ARvc0VMWcmZ2zG8Q5vnKZ43RqCYJnDrURrvniTJ+c4KmeXUFhnOa
nthM2bbVkOK0958kEV2PtF2Y6o97KvWFHatcrkHZqddptGlKrupl0M8hZb4SIhVE
2w0aRGaUfMUL/qf8P/LHvfawQAG+LWxtMP5ujQQioGKijU6gwiNal9tSz4QgBfj3
BjiYi53c/QxRAeqU1i4H3J+ioQNE/tMwNSppDzybz4XMgOo2I9bWZr2t7nHT6Vl/
ZAewrHhPaLBY0aynwW6OYpSQb3KqSWqTatCi+rGEANKnQzz3EFSTUhsQKBp2Roi4
RQxsWZ3Rr5XoAw56m07FHbyAuhwxY2ibxFzhi97ogKfYztvScl/DRwhywlnyLOqF
8acxH4jefbpROWptreTaltz/sspy5Xl/skhpKCYCEmU0Zbv4PHDY85SYqc8oc0z6
XQk2BuQ3yKx3Wv9YSZFu2XA6F4YmNWXQIZt/3pqb21a9yEIogUUIIJECu1avTkzW
FiDOiAAB2Y13sfl6N6s/j5RouVP+1dqFDT0bjutPejh/CZaDrQH5nkhN2bFs0ssW
lyd+d6AorDBDlIWqIXY3qUc5wo9ff+96Il5If/y7Ucn8p++mnjH8P4Q3f0YCYe2e
KFnmWaQUlClVlNt/45E0EZvn5Wtom11Ydt6vfpZ7FnL+pBxLQ2a+x+1pMiaMuBnd
ebMHJJwLPU0ElxGqoNOwdpXPe/84x7gGHaTFAP9b6JDaGwa4hxpcFI82dtIcD/yg
jdaPd3WurNtVLIwEp8hJEDI1goPB19sxvXULY8U3V4ML0XsOZwfxnZCV5M2c2bJX
nIhkp+4GgXR5T4X+sJBZD4c1//8BvtgXtY727GJAHNtz6Ceivvnj8ZwIpzHdO8Q/
H9K/xsqB5qI6MLTOCxtCcMxlcRYzLAuVqbolCFJY18+XO3p2JXLrMY3rl8HulktH
9RCuRVZdCDe/54tR4mAubaZYg9TxunJL0NS/VhfNjrIFSCPjMBYgCAH+whEM7g8a
oZGdlOQmRnnT/GrySk/Nmo+9LUH0J0PYWL1vklUKKdJPliKnnsh/rm1I4fvOZGyK
TcRL74WKEPiI/f3JT2k/LrsxLxde+sI4VKsrQvrczDei6a1sv6OyR5J9z7WYf6DI
CakJcUY3nZEpxf6k3hTS6QZo0AQ77lxnu+nfZjJrh3VQgyr8avCd2N9dpWpNml7x
M8eh+z+PIT0FBCzN5a1PCHu3cE23lu8NW4BzhbK4Y2kf1F6eGMlOh57f0uEO1bNu
nk8tuOiEwmrH9arxt0oCdMqOtG4BJztRPKtUfRTEUOU96i9Sj+Czp+EjGOcXyOhK
EhlaQjpFIGQJh8gcuaQKdilyt9CSHyluYpMMvHjk4jSOGPmd0btk78UWTdUXMEpo
rXiqNvRR53nUE3ahAnGIzRqXw9yq5qSKb0Bwkf90lG6CJ+w3HppfF0/7FWCVamU6
g6B5lNWee5euT4W3t34O+vg4//ZwbKY3oY/yueL61TzIl7GLSk/RPueGVVTIZgTo
rgelGV7sS5Iai2U+s245ht904hdmOTdOxGR29fmCmBGN67goCM/cpSQupU4LJkQH
cc2zhuXLz6DzAto54/jNN6bNdHjPFqM5y/xQ/Omk8PJ6yigatauUGTLlB54mIHtI
u3SHBI7FOtAQGD+EnBi6kpg1lZaJI4/qRq6Z/bYNO75rEYH85NsiAGmWQFH7JjMj
sucIJBSAOl3Im8C/k6lDngo+BV3JgXh3xhT6izC8xH5Oj7+G3Vp0VsKwjHsEoBMM
o3/gVdV+iO7xO3pYTaNpKoyc+KO4RDxoAbmbIlfppZrmm+Yy9rHF7/dkMZV27M4s
GCcTYQRHLzJev8o34GtVAg==
`protect END_PROTECTED
