`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0MRFbBAQuht6D1e+LUBDcsTJNvskGWjkRYUaqwpcE2GHfTy4TNSaDPvhsCNhPaXR
crqGhnf9scdgU5Td7kgWlB1mr7oay2+lB20QjHgIAtQuwWMGSp0MZichivzzNEA0
AAlg1Ilo2W8GcXaGeEeiB188HHk4hpjp1Xa9BFuk3x2c3ljiXf9pXv+M+gUmZXwD
nlADrrgCjBjLWUtqhSqbPIxwrR6pgTmMhncmo7iSKMj8RJdjdn738BSMbJhJ91Mr
AsPnr4/NpxyFI5rUnNL8kWqTiIpiFW+vmUS1Ahpqvz2wWkdwjsovgqlTMnSUATc3
CiS7xRKMMFbOL9kin5scmPKmOibdSJz8+lsqhLnsyCQEMsRFz+FJgrOHqvdBHC8t
Sl01EVL0RnIJD6AgPqDDyvn1RNZEmjDcuSNlKDStkm23oRE5ZiXnyRlp18d6S1zY
mZFjEO0anBgQXD8k073qpQSUSHB0gTLyePcA3FbeD2uz7JjgU8jYeBtIjax5hrlb
hAocGHdhWkgZ5stalJw4eO+wAzn09u9sA6TgUKf8yIy09aSrbGcuKwphlBZ3bxkw
ofrKEoUQeqCRnlOHCfIb/NmkzxSqhzfX2nP2OqBvrvoPk7phn3IfKuFLNpMN200F
KpAtJWW0J6X5BV6b6O8HjnSrv8CsSnI28BHuIyGLEWQ=
`protect END_PROTECTED
