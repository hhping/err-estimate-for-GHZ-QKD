`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oN/PZwIz3Oc+dLLVW09wmqYdS7YOANcCbf0GU9WNfZr7wuTI42bkJ9p3263U77RV
uBGT3TUkbG2obCHuzxRklUAcXM+VKLSdIgzXZ32zWXtWIxnv+IXGZLx7AqR0uZil
5AV4jmYSHG4v+NoI/4F+6xNyZbJ5bAMF6iQ9iTIJnw3o4kPmHAkU8kZKZ2oe7DYs
2tJhZ/xiLVCGcOpskDvqg//mCfC80G7cvOmCMl6r0YW9YPiZGF+dFVhwGn2ufQrK
TpH4UizHLN5x1P/FGfcod//p8ys/Yd/ARDAabnOhBBfsbK//tl3aocmXVDaED2nd
hTJvfpA29NgaE/wBxVzc+JaNr+gUY/Oz5Z4b7SDgAqaI5HHMp00f2R3VrlHOoMas
jxGDEUmhDghFX+jN5Jdhtqd2IOrHl38d0c7cHpWfwEpVprMnWuC9JBcb6aAzQzih
GZOfOHjxYnJNOIIwIeDHVDFFRLLowGSPRJAih2ajP7BgiMMTQ849aFO8swSFe43X
ahaRzgecH0jYVAFGmdWtO/psJT2ldIfy+hmwd+zeZDftEh+vAJb4VsWsFQtXValM
ZV1uVjmlbUcJmIv30O7Pyv/ryqf7oWCKvSHHndpdMciGqGiRWq45OgDSFJXbSABD
L9/2CeBSPElRtuTT7ZSXVoxeDUeawQjsns8dZHQ0DEIMJhyq+wClU3azyOulU/Zc
OB6j7yOds5dFJHi2Zt8HBurlRQlV5LY1mFWPBGEknkGO05sy/oFXNrt0u241fFbB
zwTioqHPTMIpDkt4YXLlIJT75TZ3g30f7HsgBAK78uuZk6EkE9q6E44xmFV6bYBo
s01hm+ccTBrbRRiG7S3JtQzP+pOY/c9yPIjY5HreaqT3qCcDoJmBcbCXpavIBhVU
XYBaImKSZd3+j7wGHA1kUFvv/UZQdKHDM97PpChdh2ORCDnVHvhfsxtxiIAnar3w
2jyhwGpeIEEjw/BAin+94l3sMi84iGyGwEG1fhK9wJIIaduSyGujP/NIXdVPJP8u
T/jpcl97T1/520bUOFIivfZgvfRBPc2KJRBTQdnsq7bs0AoPGc9Qk6WxpM56QvRJ
rwDerCOegMVCeG0Q3r3pSBu+V+iBDD3l+bBHKLsD/ww1t0xzskBWeU5zVqfxTzMZ
Va+GMPKNfPk5jomYDcCw1laWxV8LyTA0EnKAHGqjIKMHY1wOJnhWm+sl6o8anSAO
OOiMSa9G7eKbNLvWWi1rq8n0Q2+l8YhpiJamBEhRArABvBVTukQjpGk9W3KqJKsN
Xz8oJrqs3wzmSw5VIfXVrpDQJyUOHw6A/TyEpoJIwXGK0yzQmA+zXogWaai1NxrN
N2fj2ftB5v853DBXbg0BCoMW0nHE+y8WwSX8FhLr8H5DmOkmH1kg91j+JPV0f4wb
l+j+KANWuPF+/NBkcGBYQNecbjkeWDOSS48z/K/QO1c=
`protect END_PROTECTED
