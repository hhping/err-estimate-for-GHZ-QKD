`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTWTjcppXox3uR765h4dw8uCkQZ7Omh2vCyBhDYwbAwpeFxzPHY+Faj/+UfhB4nr
c8arPe+QbzW9DfjuLYP66P2bTathLfRVmVgXMSJIWvrt9Gcj9kYGOza9ByGAgADv
t65U2lcVu7Af2/ffIcoHoYwze2LeU494MmlqAiB9YnB75o4x7aiLHrQe/vzSLY2O
1f75D0MLFnqQ319FqaNV2pb7fWa4gOJkz0ExMazBss2U1nMIDU8UsBhtcg+dYnVu
hbj+trDo18aVFJPpmUPsyrwCe7bdXcxEnnTcug1J5LZdjCaMWrHJ8b1AuPhmJR4A
PfIM+99734ni38jmX8a7N5LUWlv/4KK+VRFTjDevKzrzIc//mck/CVdznq2lN2c/
ES9quIkoBxeCZ9gQmOFMJ21P1T1/cMNRsK/FQ/qWXk9jZrny02PgH1ySIsoS86vF
jVGfKS85rCMgNWSRpt3uPLaW1YOEdn3lghdMByLid+D1oDacCCQ1fWUHzYU791dS
TlGShivT33gxf/EtZziu77dZA87e2cHeEhKBr2eVZtb+W4LLYIzt2wQ2CTvx5b/6
rUCxrxwpMZI+VJgycUUgheO2cG1W5K+/nvRMm3s22aE9EUq9g4XrpM9WIWGyFQh7
TRrjUqF6cTkKeMYZgXv6oebKsFUV+cEk4MVkh7zgjKW77Cmc5rXqV9cSfBsBcSe4
FDrZFTpdG6RrAMQLD4k5RE3+wvEqhziFo0RrzLL7htbjkERnmnUhO0e4z1jnI37i
BlXgaHMUgVgBXbFstofycCtoi1lqcPjNpZSQx4Z/nCVICzPPf3RnNROqJVFCiBcN
`protect END_PROTECTED
