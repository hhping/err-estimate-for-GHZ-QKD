`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dxdj23THecGJJAmbK/QTfOkJraBdHH/HcM8MVcfabkKVq6LHEv4ekXgPyrZbU8kB
rHJdOH6nj1gdYtpPc+EYHOC9Acj58wL+1GbryaAAq8eIU17EtajDkachemWAGL3K
RhfSjTXNuXVrVPpHpHZObbIiIRj0mbFCoUVsw4ruWoFMfPc3uh/tcy9cjP44FAdD
QtfJVod8P5EjBz1Z8lLncy7LcOesFGZ86ztUKRLN4Zm+gKYOabCvDbYoMTVHBROz
ZqaQBP57tVonV5edZPImwVuSCNFsG7wq9LEi75wwsqsFJNh5Ppt/n/sJ4yTGZqA/
kDeYwTbooaofhv1b+4YCW4AHHEgbPqYcBfUiQD72P4VOFXAW9wVuF/3jrRv048Jp
azN3mBIblQw266yvszAeUJnzCULuhPIoZS8Ieq/dRui5Z4rw4/xA2imwA5q4s1Wu
OghfS+eI7tPO8WTpFQ90Fbxy5sJbX7sHHq3V/Nf/7U34aUYXjeqYZLgKwkSTHNXZ
epewJKLqAu5W3e62nIJ4B0StEUTpTpDWw5nEq50E1NdYUXd2hQzaLRcJ/tIRDA3X
b8M52jt6u7nfgt6J1zmJ58VctdqW4AZt5Affl5KW7Be6OU/6E6yapMzu6AI7GPaW
OwTW9xL3y2pNSpKHh0At0RKpLs4naxh6H4mbLhOdxva+CLBVxUSLVoIpNYuVcH/W
IA4OvSQctn3FREi0SzbyZRQGcL5Fy8UEu1O8gPjSHEO4W5GkTjCcnapvYztQV/fE
CBH+/TBw0C4kwev20X0fo9j6DR9A8Mfi9Ksr0yW2Uzb2ThyBW/EjRo6laqmo7ivD
vHcCxopSow7vh1GudE025lYGAIRs0lBwcMEXOOHxafawbHCAecuHL3dPDlvYylT+
TjrY4jkUvnG/LZPVU7tzM0cZ3PR2bvwBX1//Rmc7RHlwn0iDTl+/l3cDZ768Z8vh
c+UiNUmKTi2TK8poip1Jrs9jQtn76t0ntrMm9yL1OI9e7giw+xuWq952r6W/gsXF
BFc4mPO7P20XMiksK074Qg==
`protect END_PROTECTED
