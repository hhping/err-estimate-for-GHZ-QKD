`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TN0Y0dBuDIvhchp/ludUNcyqefSI7SG91e33x5LN50tFxspLV8GHHX22E4Q25nob
Xqa69c1dQmyCdO9/hf1f+MPOLMksp9h/tBYrU/FO5fCaTO+842IHz6KTkhR+qMxv
rOxy0sgu/pCEcu2SDTPNEm9oD8/YSkTxtbFwUa/K47cJ/XLKKDwelmd0Aket3dhb
gOUPnd3jfPsqqadk8kJVVWMBSEgxJ8ub12QubbKo7NQAy1ndCd9RY2vHwJpKJg8T
OKXGYdIkitHziKS4hCjZzOUbb5TwooDS9wT/hKQuCRWV3jdO1EQRLsqSDMC1X4Qp
0hFmbty7f4XoKw9q13T+m/NI83XglL2T5j35EOxAzck+zXDuerEy7dmWjTqsfMO3
J8jUdhOEE+OvW2bit6WTGuzvP5xCG55OKYVE4Xd22vifcdlRrMSyq1LyTDCKha8w
zbmysKj9DDxhctA0ac57r5VbsYNNlABfLw9pgPstWqR+3/erAChfxpcQMoH5Q4e6
yilvWcTtQwTuLqeYNfl3oIkWB5V++Uk9UfS4X/zgdoy9X4dP4crFmrgqF2Shenc3
vVO4LQT9DLh1Tl7dDo8WYQdRa2ERIWQVyk16nPt73/9VQf9F952tE0oSVnLw+z4U
Um6Fnbb6JTDrt3ynA/LV/kwi8bHFpV7Dx9cV0u1fTq+EqRifAc/M4WdH5nF17zs5
DVLxH6RsIoxCHKlAp59dKvCI9e4Hi/W+3V8h6Smn0qfpp/f8h5P6Jo0l/EeUjVu/
EJrjOyVrG7Nx7ATS+GkjMu0Q124F3w4mK+8zDSfmUeVuKq73B/jKKKwScQ/2u3Ye
I12ZzHNp1NkXhXT4u572A4V9L1hFlN1p3IoCSFqKWyqxwg3YELp7G2H2imneZDe0
4b1bpQNeqA3SgVLZCmwllkzIy0Jx+/tNViUvyhEzfs7XJCbWDBtBu/q0FwMooFFN
`protect END_PROTECTED
