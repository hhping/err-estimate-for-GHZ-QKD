`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
maN8yO3hqgOC00nkWWGViX5j9HzxHjnWaVx6fKYm1wvGnFuXl8KD8BLp0221Dq8Y
fcPlR+wTgo5KX4ePfvup5h9tkaIbY+XtcFSnnPnO5lsgPGH9anNN1qlreLRyd4jQ
gKWo+HjRlS/6ihA2IN3QxuDanX/31b48BG5HkXClulX933MffpKvR6EKEF0fW0s6
PmNL77Ss3zwfVc3x6aQCbdsdE6jfPz7OfPV0fn/WuMFi0+P99zgsX0xh5pY4sKui
x7ZYQKt1S4q8We6uu4X96GaJIQ6O1QZNfn5wUhcz5Y+LAJ6iqda8fKWAsR4JpT2X
k3xxYIDFO0/NaR6SrHtgsir1YrbGk0CpmZrdrrdOG5SNpblZjBCNhQIv2uwj4Cww
L5JuMcmRj7gTtPiNEH+WoZEJAFeUj5UcRuI61lHyuA0JB6wjXCD0JffIM2FdfqkB
1Uc9L6viRPZVaepsT97hqFmx6jwhpbsSVP/eYRhQlzOPl8k/UZUpQLdUaoJsmf/N
xRTWjfyU5C10GY7ooyhHpXfmVuGSSCF0K4MqH7aFhMVBdYPp1q6qC4khp4kCPDb/
hRWGVWr27JO6y66KseiE1UgEoKTWzeeyW6OoyvASVU99nm6YqweO6Wlkibz0ekft
5ren/8bYPDgrWLYV9xNPTbUJOWdkWLtOnLFBSofyhA0nLXaS1UvN+/1CKER6RlAr
uR6M8Gja5u3eyayHx8WuO6NPHC+UlLEnXqF++VoV1D2Mn5ldD8P9E6dWpT56Wh3w
uEdFbiF4+Y19lfD+Eh6yMfCEBsKNOpsPXUBTuQZurTfdWZHCpQwOJGhiqy4wuJOA
uXEzW6E/2M+gKxzpJq+poWtV/i8Qfi2d5e4FQlyibGNeO+7IM5/TZIDvqIwgN4nc
5FgL3VAywG8suqoQ6ZCvywnAfNt4xg8PrZ1IgD4fqQCPOq1CzdrjZvlRw9ZqzLT8
a0F0D6JNp3aVRxp59527p1jvPNvNtCOQQkaHCQAPHpEU6r6Ufkk/XbMpoNVm1yO+
HzcbgnqYvPMEyQry8gw0gG8inZWA1Gj3+U2junTwWvDCbmkO6CNJtg2dOhQcw20g
Rye5So3idz4zMSLWvbZX1c19GUTfgGejXpDT6QLMYlQMAm2xYM64THJV8jnsEY4g
dtUS6Qky+oVkjBu1E+4GwMttq5Wz5k7ejirsYBbNvforRD8FovKPIrTPCFgHrmSp
uNaTJigyfDEctLndIkqjwkby/eWmH60mx5ZCosHGM+zEseWTEVNR+jjvdqxQvga1
o/Z8a67cOLk1/fs1Qpv5td6pAmmXsPTBgQxRP1ZjtdXCpgbJNyWYwtoLHL+hSThk
q27EeD6mMphIeg0MjJ1fETLr/51U2wNjsaUQgrykx2V0j5DAf4TJ4/Z5h5xpWi8B
xaYurzdi/9CwSVC5B76YV3syYH9XfUMHyoUnt8W0yckzwXwRi4ZV47X4ia4DQvv3
tPlcU+yWTNQSLLLooO9Xbj4Wd9ad4K7poCbMuFqrHF0V2/ttKUrGyWJdkLFQx2Xt
edeRW2lyeha/vKiJCwVVkNgJrEjSj1JY4j7b4mX4Mk/5IUjFFKTqZyf7z7K6OezE
IyRuakHmjxfpVAibmJBlM0Z2BT6KUyly00OCkfssEDSJXvMJkece291ijCCBkY/f
PE6+6YDp2gU/TSzvMghGiHUq6kYoVU/ccM3+8+ncEFUYgeNDOV5QWEEl/W0V5uTm
/YmByLeIxlwkNANH3CfrOPhE40pxE9o6bQOgla5nl8/scMtSlXst0RtOWcyvuenk
P4J+ouseD4ndGjQvqP44evUj2O7NOX7Z41305+C6MKIZ473L181Tn/8gusEtEU4D
HlZhmef+OMBOtSN1W1T/sAIHHBzA/AbYqGd6AeN/skeJseY2Z8z750nrQT/fTabf
00FeeSBz87rceq05YfIbThSIsNFtupj5xgSt7xObZDsxqQk+2xQJ0W7SOl1hJruz
6+VPk/bq0wNbifBvsQDJXSB8PHxmQpuGI+t0/ac+Nppj0wEvsv+E4O4UF4FmWXtN
vfNeVReDGpsLx02A1IWCFWM3U9mUkUArHWZvVfFKoM6dDrShwNqDNiK70ib2iO9k
nDzBv+Jw65DVxGIKJkpC5QzTaNBrWBAdfpwnZS0nkaVn/jMMgcwjzdBnXS/6Ip90
Eh4wlc1yEXECcCMD+euK/1rYxusWQKpiRnL8rrJjnk3w/5ojX8RUpG4PvqHyYEe5
6sDl3it++PmdrKNVlk/JIO3ZNrzZ4LL4/T9+7f2zyXf+0IPqYliaMjF36Pits3a0
41TeXtuI6BIT72sM7hHabBWozTf01rBUi8xuTgWp3Cmszw23QxJoIpq+WHFQQjWR
aNRpmTcPeKyOjGuzciJr8q8/LTTy5wqX3GKtWx9qW6G5iPCpYpTcw3lizHFSDT2n
EjV5zMEQeb4sfEpamu6RYbbHJaCeCw+O+M+n6FSPNceR7K8YIe1Ibykcjy2VjkYz
6vlZO2bB0zWNgq2pAgWNJkNwDSlCaxefd6fhFYs/zQf3PLTtF5vjZkjuJW4UKPcn
rZtAxLpVPlsJELyQaVsUVMJc/OMf3YkKFOY9/Jb0rJs63e1Hv6U7tHFprj1XtFvW
UBW/VtM9RFv2xQustJeN+QZAtGXPwpvk1Lr6eRcqjyVn1fg2PtV9JhB6G+cqljxT
8sBMIlfqx/nIraFaXQJ69MVf2W+aGEWlw/HidgJ+aVifPW2NVL3Zs0Cnva4RS8gG
bIQGULbiBWNWhfatljAu+aanfJvs+2+/x6OoK3eVxuYcihyku1XnbxT9owE2lsi7
hSOXS8POHKfUMSc84+N/y3svdRnrgO22E/pQ2zNO/rYmiBFbdvT1Krk0wJMpM5mB
Xsr5r8X1gMWMLSVcqX4YaF6jOcZweG84+g2tCSog4ZGvVKievhjWjNOwgrUkSstV
M3I256x8mG8o4YVHie2u7IXQcp+wgsPwvFd/42xl/zFmEHj0Cke+o0Nvh6kfMukc
QCY9wfoYsNkbzX7G/d/NUxs993SPDJwAUX+lcq+sMxFegpnYHAiZRuTzOnmvdbrT
smhZm2NWTR/F9wCNgQY3XBz9K1Ye7QVE5l1ja9of5/1LCxeK9/Vmyvh4OwVePxWA
PDS+hL04rJt6/JxtmSeHBAN1COIZjEb4vYe+avIWDQRLqiHkigLTPVJeaEX8kqZt
/JkYsPGAYC8NZEkR44aAt2Icx9okLyXbUbMvLwxzMp2oWnN72pBUqyRKkqunCX34
0hfP8DAx4BjN9k12dZXTn8A7ekoVcqgZUD1rXsqLRZXeDNL/nug6kFk4oxqTOtP+
+uguapdETUUq1ahSBUFF2qjnrEuPnkZ3JUfQWEA2TQQ4Lt5Dl/ylzCcsjZx/ywc8
jY6guOA67MDWf5eEn6xzdWYInXROZAS122Yqr2ZqbkgJDUKh3+FN8/UThTFHab5n
wnYY1QnB2+GksJ/a8SZzcC3qInnW7/Jx2BBsGIlkkZgV4G/HNNrd18TNSnjNm79l
MvFaKqewPRx7QJSp5I8VDIOZh0/OesvgA70QCiRDQQp2+jSIq+pmGuA15ol6+Z40
Szvha5K7BQtVOFoTijJ3AkBUjzsZk3Eng4nW8jP8GNgLpaceueO6xGoJhBqXRU56
bouYG67ON2xXHZtosxIWckKCvlfynbvyn43qbNvz2G4pAosGx0F4BrzanyzgjRKE
ziZkqclOjeXMDBczSQNaN9KmA4V0R8ZgbK0ZphhMj6KBMdEtTJuy5vVxey1YYDs4
Sh77KYyELLHjrYNW7SGNu2DfKRNWx7LmCUSOooKEdtFjqujTW15etyJ85PGvGNuW
XmymWgnXH2kXzxEmCViPPwx54atQ8RgxzToNL9jptmd5uM0xKPHzNHAWaFjaOZco
W9U6/0ajT4I71RCgKRZgvnhkHYEwRVKs3HVOGLYuvUVAFsolFHWPMoSHlQ88l41A
Frg2x4OwKXJZ4W+Fjx83hVdO7kTIzdoD8Frxv1H3UUJ2vb3lLX5ukIecmH2i97zw
YdmBB6ZbG39gZSQT8Teaq3x69aeyL0F7QQF+rp6dEXpa+3EBiqUgscu2eqiQjDP6
fCu8DyszgrrJo1dWp89aXUag0ul3e0DPzY5cVesBKClClbrlrN40s+fgWvi0xHW7
v/sTEHvS5NHqFenukdNXpp2Wtg1guuaYAQmQrIEx3LreHalacDPzAelHTZvQXh4Q
KLpxsBFDVgcJ8iAhmWUHCxKqGdDwApzQ+O7NAbDXjwXnyv+whn6S7yUejcNvzePD
yD4RIXWnU7YOvXMOF8qxgGTTFEv1JM6W2I63ZsV4IWKghyKX3fHcteau+P+MZ8OB
Csl3a4TGuibIdlZKwGqKXqV74PoJ38w5JOBPeo0637Pxd8nwDIYWeI6iEDxDcFOp
TIM6/Zssd5/N1DQCY0nHxLmPoa3JEWGr0fZZNDuaCZBBsnY2em5vBetbgqFuH71w
Te3omD82TVoDMTyyESXTHudUybIeH6clL+af1SnOvXJ0uoQBqkwITFteLapxSvMv
HMxVGCq+2TbbR8JqA2k0LIElJKJYHDCe89jnBHvg6CERZHgZ8A4EIL8raTVswgnk
si72uWitDH/hdAFsVDaGPkdSIjCK/8jCddYT8tYUpguYOnkR6Tu3wn4+2fgkOaLb
drWnOlZeRoRSOdfe+TJ6AVPuR9AtBAWGHPxT4/T2lfckdwLCWKRLNcqEmyPxQMUO
IkCAF4B5fIcOt4X/QxpjvLIBh28D27ApPvenGviI1+ULGJmGaxAUdJK7BrpIS8Zt
RDxCpHx+3QyAscavfnz3Q0sLNzCjvjAS256X822aDABCnZ0aTOI3YsEeI2TQQgXt
UFbuaVMENqYkMmaZT4iUsEO73jX8qpqI+6pccExaOTw738c/2A1WejQd8CEsXStK
WYcudtLU1SydRUuTWX1uRDJoES4r2zJnojtS0WY+QbDOLr7alas6TnD7+WXjYgAf
ERHrBLQwskv4mPjHhmYd2f13OQT/CyznesZPNiuJD9RlnKuYZ9igRoCQrHIJ1L3d
stm2LvfuHEVUmi2uyrHkTfVBVv4GDB4P7apeUygB8wzLmVCv+WOKdOi/MvWDc52a
pDqyCqPJhoY7qDy2jlYVR4d+cIUJVy9LlwLHo6P7zUfdUBL2IyGPPxCIkewzhaJi
L2uTzS3Xu2pHUgX/M/qgTGDbGMCuezGSOU/itrDfxyI8dhTZw7hrX7jyCna6RjpU
q2htJg12Tykll2t0THzNBAzQ/dZ1VgK+j2KolIRrRHBZxA6gQU+RfB8u5saxlDXE
QKupTr0wUE7lOicNJLde5zShL2N11i/WOPqBuTXavZ6z70tozpnzAKqFZbmLNPWr
rSNHS0JD5YAtbivfRGSNqHjKnaf7j9Uhuv6re4RQOrrBUAyZnH3SV83HdXSYqnan
fhoWlxd+0NXIXSO9kdDpBzdxnxwpqwuTOykfdmFePIWredfibdAYnebP5L6YbUSG
WZoTl0TIARC73DK/ThL+KQUwxSQPmJba8WLeXaZCN422pyuO1NHmH1Rdq2O1iQYN
O64rvMtPe70medZ+Z069nVbAxbODbnqtuONsWSVMdvTTICwuKEY1fq5N0PfZU58w
SnZpMipaPCVftXsVq2wshRPMc8mahUoo+HVjLKsFj61MR1BKDB73Gg/70AP3Nv2n
vL9xwMXAU/KI45HvrERe2uu0hB6xvDijBhZhSxSddZuA2ZzzlhYn1fwYljwOTEZ7
BKuCRk5vaBuq4QcmBxooUHVDbQWdj3sAckHpY89u2D4EmCzFDFCwAV+wL1MuXNOY
KwQANz4up9dnSF5Gm6KLdXuJAM+k1pKBuKrDenlU4wbmGXKqxjxzPiucMPZlpWlR
QAQndSJdYIUBkLmyPnOhrGcJox7+05ZCSLc/V/7KUrntOIprzZGH3F1Eeh3XxDke
BKJ1gEvU/TvTINfMMawsthBCh9ZfecykFefAa9HlYjk9fRqTcIHi5j/1wrPyqS6i
XwV/+XTgb6Y0b4GmLWOMCNxcJ0JPZ8qeDM5wfGX9+Ubzd4AmHxvp73BgnlqwWZCC
FoXdIijLAoj2PQ7TkgkkeKt0X8Eut+1AI1O6Lvi2/N5jBVAIIF5WKOpf5zBsuVbF
zRmMi1OlZCLtqcZ7ls3K0XqbpCfROTtcEa6aKykkpXXIz8KHXSgw03Foy88QtNh8
vnZxWY21OyPmmU74WrioEd6Jo1Gh0lbZ7nz6UTDiyFWdLBSwBgAilE2A08rHtODl
qnUXrpITTcicCQ0tTJSEvkuc4aFLbYqmpKIT6QAD+kFpLQN8JGC6d3Ny3Qeyv5e+
QA9ScdlbmVTudI/a1lKneCQKZ+E/V7p6+daU1uyl/H6o/qJjiGA5FmS3DNZC+5eQ
jSdvkt04W8ycW/5KQCyi0biXQI2P/Enjsu3XJ/6rQyUWaCfROY/Z2dcFu4rT7LPD
Bpq6cHdZ+0OgIdUWtE1fjOZINSk+357N5hB7N+NSB52E5xukov9NJvjPxDVsIp8H
Xzpx8X2VGM5nh+dwxh9aEMH3ME+YkKZzll0ixUdfnMkLkD63XKLIQuHtkxmsDFAt
DZktGhJt/1wUWSryVi8AQbvzI7SuO3E2VrcZWznYp4bMafNsJnN6L4bMqWVIbPxD
UgDgI9sOPBsmFSnSH3ycE2wZtYBh+plX00k1gIYmn862fKUL7mlkwFjv5BKbnqtb
o21cq6EZUKSckyZeR5tjkAl3d4LBWnviB2kOyWLkxPmMwDM3sA5+vAu/qD4gwmjQ
x8kFZpg/JWP45odkIO8e1iSbrMInbm6M3xl8kJU2aatRe9nhZnA6JHF+NZBWQDFh
r29XnVXp5ORTjaj6iYSEfVRbaiEt5WtXR8VuJT4dPpmFvYDJniPMzW4YYQpeipLH
L+TejGeYZXhKwRmGWjRoggOi+Ws3MlK3cTCUaDelcFdBOnOOcrJ5DwGWxg9RczG0
rKx3R7uDIIQSEChrKWR4sqtCwWMRntuR6TQJyZatYWJsn1uOm6WuyNoQcN4be1G2
e9rOVmitvE27WWNi2vK7/Xn+F/XB7hX25DWvQ1hsvp1af4AM9afDj8R6MJs2eRM0
WTRy4yA7lX6+N8euWiG05J99WteK523pUVtbzd5eyym7NwRV7S8h5B+dORsGaG1k
Aq8RR+MUgbYvC9K7eTiVBG4/rYbv/glmMtHYF/K8HJYZwYExWM4DKfu1gso5fODB
EXkE1xwkdbIQyJQ4/eMsmX2/1bvWAd5ANynUUi+u0Sx5zm3jNUk4qTGCtjPyjebP
xIq1Rat/1y00/kcpE7nrRHbyJWhg2KUTNS5W/+9BOxidHqkNUGDH+CwC0tFVXtZq
mc5u2WJ4u0KHGCoJ1wSyGApG+AHnrMlxlBNgZ2pBDyUyji/DyP/rlwCj3sMYfcmN
n+l2AVB0Qux63DhL+d8QgFRU+E7EWG3VfrOcfxFpzQHIARuWuldhQTpDcnK8xOAL
9K7e91bWtR8zwdZbdllnkDxTIbEglQsl95AFZQxuttRT5PD627Am7Wz5iSg1mgQP
aM6Fy9Qz6WRz2jUHOVlTSE/9BfW4fDWkzkGSZ353LPM2URD+5VQpP3TVJerDEumt
uYAI48g07UUNCaBue65OS4E6FHB92miTRmlpZcwMc6JLNN0t1uB511os+c9doi25
BQKFEUh4pH7dmrSbNW1XKq3RIslb/DzoBulTd0Cmu2BDZv5TJxv+WMlxf/9iNkhS
aUDxkJjJbKReBZdhdXg0BhX56vjZNyWS4uSsD6N73j5or77hZbmKc+8jyxV2zSt9
KNF37dzViR5gxWg3uGGurjMHQ83qVF540uCKyOlRxMu9+mKaf7UCv4I2Zl6anOsp
HtIEACecWmmtjjNrgl5uuqEdA3M7509aaB0+krg6qzlXOVVB1PT/ZoamlAbTVoFE
PH7FDIPn+tp4CSBFpIGF+tpXZOy2WKmBnWShqm8iZloTxhZSH//6SVY3Eow1jAA3
HBXnRitzqScZr30orDbT0ffE0x+K8kz/nOjmXJd1fpPgTs+iI78dibRRsEDKRTPL
4yHBcg0CTcTTDfe/u18nk8iY5Ys2hU2g31RgFQ3E/4llrpPy6bMsriHjtcBWZDKB
9rpTeAgpLhV41XBSC8GLAp48nm5H3PRtI3YTgvqauC3uJDYypgwl3Ckya+UQINb0
TCJyukGhN4SKnFGZEzkXjAJuTtZteCYDRJ3ORURDasU38jk5DLOqi5jAK4AIHLfl
Nc0NmK4pHh14T47rWrr8zmzadVYhEZglcs4X1cq+duWd/XiXg6EbUJcazM7vWt9V
8cT+EXhrNJswXspqEN2BT/O1W36gctUnI9TPI2GlR9n0ewwqc+TLHvxIT7Tg0oF1
kFO+Z7ynql/9pxX2c0nYoA739CRQsylPBkz3cJ1jEDFRI8Bi4ZGwdZ57XGloZL2Z
gwl7+85BT99gODf14I2Ug+//cY8Qj8NMnKYMNesuyieJBVAqbJJPPWC1vyxg/UBr
GSh+iDsgvqc0ruFYze/atVjjqNgCpdO0HSlne9CwY46oM2VRP1uPWBafTTA5kIxW
ow4rjXger6/Yuvd5uoTviX4A0voMf8G6UdaXv1S3Y5rqTSdTZrPWgn8c2Hy1t+9Q
WzSm4x0JL48OeBSsI245elhNZbRUiHaV2ziydOgOs5KHK9bxUWRXwMNeUAfEd9XX
Wr1Tm+iM40w68lufCQziRzkZ0zXh1D0E0/lL7gFBAShhUjczSVAsHSsMunoUOhOY
Zv6umprUg2cbcUmeQGxVcRqvbj6T+hwsSElPq+vk7WBTKjXg8sxo5WmHZ3lBgpzG
CwjKugtTbTK4nxY80XP5NogRnYxBmK9FAeTf1Opwqjw51neYneAcbilkwT2aJB1Z
E96j044tXRPDgxBlTsRSeP4t1XBWjAkMNj244hv2hqaOlYmnfe42609yf34MLa48
Wz2svFl61+Ywx0616tOyKNYnO4Q2AlvMMuApj5R5mKZKcdHzKQa6EPAGPQ9Dhtfd
dHbnJzTogJaxJgylvbIMSJl+0cbH9TowigC1HBDRPVNoDPiteFykW9ODx8G1g+/+
liN6ZY+Krie+LTDdmALo1axHZYChnVFJ+wZN1swtYbZVNE8LS5JEZ4XNArz+WTCh
8vudrRnGRjaY3kPvrK5ARkLSp5aOymxvcMgYZRSQK0HJzRYmFGHNtcXV+2LLQtFD
`protect END_PROTECTED
