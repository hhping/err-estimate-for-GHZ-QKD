`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eIoisAkG7mFGXY27w4dJW0oMf2Hx3dPp2EXCivS2ZM4oWbyPVz9AwYLY0mX8HovI
m7fs86WIWueHSttT52uhezXdvTu7Q0MehE7yVsz+bXdOOLK/GBNLZWEgUkiGyhvH
4cqXIGlbPdKznObM1TRHCXRGdM2Ipatvttdr4JpZBo1q/6AuDG5Xd12/iUJOCDl/
uJSH7oKOwXdnpriDbAel5eEjp2NBDWFoh+6ieId2MqdhqqK6qLUbDo/RAqRh8Vl7
/JdTznkB9aByKudBROPozS6S0ZrBlma+21e8AFcTFcbGeOdE5HKRJzO4ScaBwMba
DHDPiPqufQ46LgBYzy2Tb6PClfBn/6HuiMBKygjhdC/iZ2r9iP8oqm+Z3r6dL/9s
0j/WLClpQQaD2nqEwC3dfUm3ETtKGkpsETiCpVSnfrmnC7/4B6gEEmQ70wlSNfVe
a8OkPpZEJDOe8fXWkAMshTWSU//KzFBPfSB3G52ykJ/RiPDkOERNFd8eHDqqmClf
c0eYyaGmgJkv6EWu1bzSApAABU0/4RFpmUEQyWIAAqIwn712F+XAxAyBVKnVJ+B5
IB8KclFhdfFeGE73Eg3wFYCWxy1u+nON9tCYql+S8GdFKSdX2C23KN8ypksgFS4/
Tdwnq6AkYlN75Nzlz63QQygWDalhBh0l76s0geQyBN5JorGsmXS/B/MhBU1DHSNo
`protect END_PROTECTED
