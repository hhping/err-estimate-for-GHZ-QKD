`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMvJRvc4ZDgTmRIX9sRejImvnxiGJpubQpwQoBRAyFv0JbyEywaOIWrDZ3WWHvAU
AlszW1Ofww64vwX423FSw/qyZdzvunlbWE+fjhjhEa0mE3fJ47phRaAyF2LJQtE7
gsS95DEA7uz9M/V74sDG1JJ6BYaRH+lbZk5TP76MHOIvIf89uj8P32GPf0GwURqo
XQWssHdKi0k33i7+BpCpGc3HHKg+NaNo1MPADQHv4iigD43aKyYJRZtevS/iwi9m
oNWiLBnhk0+Gr8o9oKddNeIAGAbCpRFY8bbqktwc+5l0rOfb8Dmc24qtF3FTMVj5
fMajOLvVYOn5zslygv8D4z4C0HjKqLCCNuO9rgqYRyGQgiyp2A42n8IJv5D+lj5+
TqGpki1xZR4nS6GffmhxN8I57jAAVOOuAw67+TaRjGTTtIJCgPQo4vl2r7uX62ay
q2FDDIMy4LfAXi6OoblgiiYHIZPPAOHvQLy9rFAOvkkMONuBblHBSz4FMtrVLxfE
21GyIuSHWZVlJQApOYatld+2qxr8zkWafDQDyYUB0vh5dHOehMa7afQREBx/A4he
jQtKNXdNwPvzwulvQ5b3NhhvCmFUox8/H0Cvl/OoeeUsIF2kL8Ytm6hOwKtvkIex
j0J7ZdiSiYNAfEG83fiWD4AoKcup2WQiJUP5HOt+khOpvLpGIrsgOX12mEJuNchm
tuUkliwEMX0imLiCSdoeKf9aYACRZ4lvOPf9Zjp1VfGzJlb8b/sP8o+bfDJ4Nt1h
egNEhlGTad7YZ5XMPAZ4PXfJOgzyeeuPuay+aaXRxc0wNqMnNiy2oBOG4Ddhi6Ng
K/ye8hUkvKQNDEsRRKcGuH0n5WyEejga3e/c+qmvWPYn0vd3B2cJOkpWFtdng4gZ
AiegXFJ5WqIAJXA2bzUAo3atyABlglPoBFO80K6FDOS1GiGPxKfqaIiKMj0DUsxD
ICz1MKZb8591IQce/gQFPLQQyf9NJDXoXBc1V7US17rWSre+djJAsyM3akXVK0iK
11N0e2lUweA0Scqs+EUl5DY4cfHWxulo0djZNnZ8hgN/wPKyIF/9Fmu3uhScJrGI
dyrmbJt1l7k39oZFMQpw5dwHSbcKxtesout9UpS5RqWoU1oJ3M9jhbl/jEaczWOH
AFaW0QBcwf9TINGKl0aUb/MFjzJZ/welqf2MaaZvDR7l2qI9oWPqL9iR/Ttv5lYZ
s2u4Fp4PlyIqN+FTeZgawka8uZ7qlNctChljw3q7KSRY4hlr1lrHCWMI1+tG9XYq
ZuWCouCidOH98xaEsFbcGAwOaHmplgiMSee8IANo8zNIpEpR5Dc8WFKdCNC0Sdt7
pMoUFnHUpTizcWGwyv77OKqDyk1Q1rBKeo0VRwXfhpuPiq/Fikost6jTnT1yOFAg
jWLghoVKB5gUQs3re0aA8DsLR5wYTE4QiY7CXmnEjteOsNMFfsaVr/zRDxSy0cih
CyAoZE6sF3i4BVzHgVHWStDPbPlKk/uEHWRPi8kqfiTZuWNnV2+Bxbs2DakH8T+O
IwclYYOQhNglVuGCoHIfIxxWLA0ayAQw2ECI3dJ5+rLxPdKJHuIKIvr22FBoNuba
c+uls+FocFRtq9A3W033weZNDkRZf8+pLqJ6Nzj+cVSFWOx1DCmEgK1MLkHb1h7M
4lb1rePbbfVDD4un+ZVJntRHxvFD3PiDaUz9PqN1uQIvyRz1h0J+vQyEUP+MlVWw
22qA5IVYkbxgnXuG1uBPGEqzZiIGDQv42xrIp9LuHcnzdZtjh7Uw8S/hWm/8JM2I
qcaH0iMYsm6L66Sry1XPxdf8Od3in6ohAGwYv8kXATDI+ptM6xLhCVouhiArlC9v
Y2EgJlKdRpEvJruWdV4gRlrdO6XTsx6d06BQPzxSUzh+dpmVtbTTT/QLfBYoi+QG
6eiKdkmtQmQ7SVib8CR6HvHlNZc1yIvSQF3WGWX/vLeqAygfAQU0iOrquOmybOhX
RX6VY4EMcdSL5qwqdHu0XHXQUYQa1gfkKmXeMz7rxZdunmqKgwJZpIKbd9eEcogI
GIoYDnSjilecR3iFSQMf5Atxt03b99UoTT1GU4Os8008QoJN1w5CLWmZ+KGZx9Xj
fQQ6F334VPlEhBtBbsytOFnrvmfbpmbfNQ6VuNwZs54E8N2BYxE7i7+3/iDYc7ZE
FkcbLvcsmC8Dmexz5N/E4WNmoB7+iUGaONyyNdQjLwWx2n/Yf9hJ7F9zuyTUxCDJ
E1cfBwsJHM1Q/vKaHtnf0j2on0Q+JNbh9y7yDET6XKBri4ysKpRjDaFwepsAo95w
ySJSnB2J5fhoFt/zeXu+1flpotoAJLZl9NKvon342nRrmIAa72TQ730bDjDPCdiq
9GVZ9BG5F9tMMvwy8jWX7MAkrn9YphYSxsVo5/IS2ETi+yPyP7WvJIGGgSSgYqxK
W9xfdJ+AoN36yLbVlpiF2tT0G1t7tXSxCNx7DQK53y7AXdRaYHhdeOGLYj/ZMwxr
15JgL6kcQCpS2JHX4hLPvAeMcig1fn+x+/09JK8RdYF5kPDZ1ihFD6jcFy/OyzyN
GLR0TTqfvRxBIDNnk0nBvxEwI0krrSZKCPudH6EGjk7DBfB9qoN65yKYpFHZf6gn
YOaom2uGOWwLH+w3+1Xciq6czJesHSeCezYsvp9iDCBS3CvVMd9+sL4+Rst/04mP
FTg6FJxSunld99In03vzJChKgEfBJ8FFgy15zaIzmWhxbo/pudYS/nz4kL4vKP8q
9xF6fWDe2p3kSK7MCrXymm7ePU6n+qMrS9fYcsV684wiwJsGBCYuVNEK0SMb+RAs
IVKrqnEEWD0/jBAU1RnnqF+1ncy1dJ6KL4UrHd4UyC++Lqug5DcL1mf+2YmlFBxP
Ouqi5rLl8lLi0wLrkfHmo0LUfSZIOdfuqRZDk/av7PwFFfG9wxwBtYKP7WSE67yJ
Rh4Jp2tAQgilZzriRYjBKI3hRBi4rKzDz1n7N2JlMloHd9wJHV+RHBd8d7L8mdnS
LsnECLyOBK+wjrI8Gc7jSYi9FUZNorVeCfJkP4Tkl+9MOh0fX2Nx5KcZBqUEnKKV
b2rD2ulRLQE81y7Jjoep/TEIfngttojGIHxbfcxIw1fVyNbOcLP7dI+RoipOLZo7
Dqy8ADmsCtRV/Y+eFJBDmQq+oYJ7JCgdaWqvL6TS/+8/0eEHzMTkQvEYhux2aJlV
QOa/74OCh2Ahjvh5KzXEC69WDAaGtg7FmZma7MIrJYOZrb00LrkGEeYQyBIlgSTd
56nxBbgUKBBVmdWI/nW3yMuA8wGF4AUzlHQbjUqi2hUw7oVJeBz58aUo0Rx8MpQT
E56ZGUIDCeR/PCTsNCkxgShh0hxezokPaol20r+Z/ahFiiGAtFZxfPpzanBV6SH2
TfMPswgPU1NhYmV+wlGhQUf/MdWXhproL6GN7VzZsxZzsxAqO5YF6sIUWcnCH8wR
fcue6puvL6avyirNIvxmV2YZ9qSa37F6osMBnfPDucofLwlH2gVnL0p32mwd+DaM
2mJLQiIcMBCfdhGCEQ4VF+scqoqXVfxvfdYpnhkZcLOU21ilAqQnNLmbQooxjXGK
9AWlDFoeuhjiDo+JrNYnbVVRa2xWHrQkcsKkRpM2PdNyxSxh6ptg46YypXIYkQwO
3VSjA9qFjFqyaT7hCWfnIrxeZ8x6ZUPwBXfquMq9Dq74ykNazmpdEueZwJDiW0bM
i3hizzrFkPsiZCbTkTZNH/SzhiuPBLnt1ySrYWA2BNgAisWomKNNVAMcJoOVAWte
+iVSI4fZpl2gJa0SMwhDSu/FtdvnJ0FK63MJY7B8u65ISc0Wz4zkJo+F1rURIp6z
DcJZJcbqcAXmYLxiNTLXrnuMLB0qiGSgHDT88g5/gZ7+7sFPY51Kpmwo7sLb5IuU
H+2WjYX17UBxRLXPc5ht4qSOr85SWMx7Iw14m0othK7UngmAaGgdx7jycbDZr4fg
BFfvB+iYinqJnDT7w5GJNtEpJekBRENTpUnbDb7c3h+I1/etD75h/xiM4R1JuCGk
1mGidiRbgVT+1VTkien2dzB7L+QkL5+uC87hNwW94aPreBqruZiV3ESJXveJMREQ
xszexDXDvc5Ja+QYHHUW+7FuPyd+ZHwcjOa9Y10DmtgGh2McOKnXvQp5wDPBKfnW
hxxn0lIMACb5u416boGdKhNcvjravzkVoD6gyd2KbiU0HHbuSEpc9ye3HTAdKiUw
dEfISiN0Jum0HjH1wHRFXxBpyOmIt1GOARXO5QtwJZG1cK7sVp98vYoS1mVyySrG
/Naom1yPyGuiFvK517WsvbXUs+ULoJO57rtTFpXE+W1n19DQVAC3j/dMLwN2LM8Y
PL9fZB2SbJWlUHhrKMQuJ4huOpPDwzNWqZwVFxrsEUOgunZDl9n3nK06G9hLJjFB
iROGEKvk8EpHg9K3FiGhoJXmcxF2EJXmc0l0Px27evfutxKBy/Pdvg8AavcF8yMJ
f+jU0AkkGbdLBp53MXfe7p9goQ/N8LQDQwz4ZCrDxUJ2J6y8ro/g/6yp3rIf5bg8
d6dtQhUGO3l/ynW7kub2Selje35xAPu7yEJaIR17AlvPvnRez1h5Et1xdVX2kcBU
KMWHK7KiAH8SoyGZXmUGJkACqgn8mWP68iP9dCh6TzYRQ2kVriijMN0Fp/WRvCdk
d/UIOj/zx3KXNxDx9vzz62zboMvlwzzopYlXMF4+EwFbpsIOBwIFHi9iH7R68Ezt
jKVJnkEpTtfzKYBHokoo1KWq6VseWTD9i+HjMckgm9TSrcis+Cbe0fh+ovPk4VEB
z7GgAGMg0biffxm+0SPMpjxWCnvNLfOPb510lIv+cvqkE+3ioJd8COQZpwcSY1KR
77n+X/AxbwO2PqYctDeMKuF9EkGgfb6cR+H7rvFHCFH4CdpGuReapF3XTBhkki1e
vuvGrswjkKmE3NogkclD59qPtxFTnBYOg94SX2/RL3vIMixsuG6cMmB9ypqbL9d4
lm8yaRiSNw4wF77LjrWwbqQWogITD1IUveiyVG4PMQ7akfPQBVsE8DpMraOP/0w1
Y8cK0M9+6ulWcR/Zl0jJUJxF9LD/ETvLcA8r93XznYZOESwdUmkRPL/d8Ar9r6A3
IvoHAvGmtVtTqi6YVENSc3W3P8Yi1PWHNKpvzIKRfANANLUicQXtDqDzB88kIShQ
rffpDfTpSAHIr8jLORreMw0GhXRYSV1uMZoJ010Nhe9xkbn+CeOEqN12I1YuZgma
YZW/FlQyMd11bufNr68wSmDobqfrK+i5yCTRZHI92wDxVdyHJVLuDxgUtYVanKN+
wUaL4tAESLFMDn3Qfe4D2OMMpC+taGfYc7I7JZ8TiUJWjbnYLRwhyMN5KrRB5ku6
dcQYpjI///YKrYlhOdrpTKsF1qceW4vM3yPNgxvziAzgaUYtUh0KI6iw48FsDQrO
kz7u64q7MHDwiE6bwzPcq4LelzGT8lN7DExcCLUinc4Hzxm1LyTl0ZlNioirGJKu
1HD5zx6g/cVYu0mETuIQmFGhqFbR4e4JgXPfuCKHhORUmGb/DDwC4yIcyH1fSmhl
ZS6EJrlZyUBHum23WKTscfnE/Mi/CHKQshrDuFjtrnFgloVGS1T+J5vMsJ/nQvL+
AXvFb+IYTqnx227U/j4DBysq2xYlOrqSCrI3pIf0v8j4Lkn9uwJr0lz89jU+AXsX
/UE4qHEBnSDRFNS4nMsdXOeAqp+hJ7RYJvMeG5j4MgN6EdMqxkMCB6Y4WEDzv1xy
xoD4e5MMyUuL/mthYgJMs4mUCLviK5eJk6BLoq2YnoRfyAMmlBHIYxGNu5Urt6GZ
OsvDFUdKYV42g4pcT75ybe45F3df40tAVPWI/n2pBeKwhjieVMv6+yG2lnKZwjXs
j7qqFAwO+CPoUCXd++AlrBtWnchbkZhePRVpjZSHjE3at86Nix7aHsoA42oWl21y
A6ZFR1uIIycScbQdpDqSUHJ+4vjKkpXNKEDju20U6zbsBnaz3uNRW9b0ELmtVytF
ZKIf2YDpLwmTjyTuY1xL1uiZUqVxYZO23fx4Gy5NvrA5WZ6AnkhvULeWd95qwVtH
Pr7gc1iuhiLYqQ4rUjmfrNw32zSneWAeYdMbFPucwyJmyefGTNfsh2VGHe2yMNXT
nccplyWnY9+Fp6so8Z375Ig+E9EQrY5sf00zmDV92p9M1bq78LIJbEsqg53dQg+/
nIIysicRZ9TDZV5hfXYGTD/r2P+ZLsrx7plt6afdlI2JQQwbYkyTDG0esNA1MAp5
DUqNGXokEWAboqNuYaPvFV3miMcgTjDtSK2lCFYo9Kjs4dNi92rZbEyQkxPv5MRl
JZOJnY+32WciwCl311HHkHKzwCqAeMM/PvOwxMce5kC6hu1T0HYSObLmYtHvDnPA
r2HPngpGdlCPPazratIIgqvaiyWOz6yTSwLMfC1sFTYdMVwH+GGqaKZKvCYD4RRG
hbWJt8t6uYdoSjI2B4S8V0LMAHpqk2tY4MOuLXwUg5vNM0jwKmtZNmbgrZEnpBIn
O+c6gJTbpJOE81UtDBXpW/1XUv4NoXjWwXs3ddiqa7pftpeTmmyQZCx6NEoYJGFR
4SeceEm179hc7Uw5WNmV/6b3bPDXajczz8QQZS6Jf3HyfHGqiKOzmxvWa/Oltwgx
Kl+x7Zyg2/0raHGibpz8OdZ0EnSARiPOvJPag2gVR0FwiQ0H6fOs3tlEEb3RYaoJ
rRKux5+4iLNBJI+/i+mOww==
`protect END_PROTECTED
