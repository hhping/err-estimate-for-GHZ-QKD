`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Tv5KR+5cUtBA7koaSCO7SL16O7ktl27BCcHn8gmPl5mMkZ/QZ5RaHbI3tfGUnuW
93+47bEB+ynh1zIg/UU+kAlmW8vEgxsyVKHyO0HNlNUA1LlYIAP21i48eSH/CtDl
+XcpWM11tbduZSAVMpMehIbnnLrE69q/yMtMqnICMmWaxKNPp7I9+AXqSuqtDIP1
SLYbCKslUMHoFlDIIJxwp56BsKbDkZAkShpTCJXTUUCV+xLZl9LOKuTQSffIUcdE
bbxSvCA7FL0d84cCcfmk6/udBDfaF7lmEbiMc2iZPlupJQR0deRwpblOWWUTIT0e
8dzM7TGmMF+okY8MfA0c6jwpO7kEMkRi5UvyWjm9UOykseAeyMWg7Vh36nWziN0x
/OL0WjvOiEujhMlJTj8wo8c+wpE0H3kqd5j1Nv10r4UdUqw9xW+c4XHd15d6MR1F
xbTw2NTewXzwwkSl10eSGSnFd/jCxkYW0s7cdpL503kclwWMXYI9LN3L3+7Nfjg3
sBohjPN4OSkMK2c+Bg3c3LdHPfmCSVqntD/TaLtqXDY6jmo2VsiDqTYjBBatEHzc
OE/9NRwRV+JuDXF4FVFapJCcLH//ODICaeyj/c6xJk1Ta5QH0VBLMedEcPwBWdBQ
Diqtgo4OlM7/DYdhPogH8wJt+g2U2ldZaYoP0ECl5NkVdav6KDLQQc8ayohl6Pmx
Z2YTK/B7pL8y0M0pDMegi7CqzSzn8vun3ys0iOX8oJ/eOc+3qQHJxKiZqCXeAVef
PmbSgNxpxOBBjH5T2YbY99Hr0oe2fD/gvaggrnqHqJ5QRLGGNTPD0L5ToQ+CVrdS
`protect END_PROTECTED
