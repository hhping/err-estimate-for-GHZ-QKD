`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c77mRyx86O3TOUCeqULS94jR1xqUk6HjdvZLhj7WOUqk2e0I+wxCMO5KZSMMEvp0
2avKfLxLNXlqjoce+b188FP4FL01wMdkc8ak8m2xzmOCm9pnLbtwlmrZKSjw9ovc
U67KeZj1VGAeKTMp0Miz9pfSDVUp55h9Fx2NrvMgnGpUBfyPSk6YKusl4heWFept
17IAq4bYSNnQtfvjSoz5K9An0KWJ1U8+tlRkQruCwf9kmiyDIPNNE3P2sr0WexFr
qRa4czLXCS2TZEVwrGZq8AruYp3ouR+dkB+zfbwJDuqoJHMD3m7zQ89soIThM5TJ
oQ3zKb9DDSxYPIEWJinctN608EMBcxR3KqzSmjtHZhuedAOHOwD9hecPyAZLpy0Q
+dtQOtslxbw8c3UQO3XuSwWy5rUZ/+rJBcxT7+1NR9BHJiRk3uV4g1XFnrpfJR6q
RHKwkDfqbh3nlu6SLCH2arXMwPw4Z6/ejYQ6vgDVgiFn/5CCjoUoBzniA6XE2TIw
LhZ49FnRK8KzJQUlsliI+V4WtTO1uM3Q9m+SYkzp6GWpXZANNvzqh2osDx+4huYX
S9qMlXmpWgA0+lojNhQ/wtNy2t3zoBX0Lce+WQaVAiTE1CnjWIEN24yr7Enbaygg
IFInqwjwLSP7+J0TZbBzpWyLNObWYmIw+ripDVC8SnZSa+puCRYB3BQyi2kgGS/V
YoWbxGTXbgKG3mdcRw8M0UTFG9xhsDxBb3byBJ9TBEjz7Sa+V4wfm2+zOeOjwqG/
UFfTAhlc4mEtk5Mzlem8eDOs81eypNQOxf0ezPZUDiAFddfFZMmuOhGy+LJnt4Je
AtZz3XRvWeZt9Mjh+wD59/BIlPFPnbtfq6BXUTOxTRO9uS1agbINpwR1iOcT7AmO
FMGoG8bCo3huAXyKxfj2DUTMQRImy6MiSonk3STMMc7o+/UnuQ0TzUER+MPx+LDn
Km1bCQpwDIGzblU9i8g/9/as8m3DTSr2AEeRjAQ0jowQvZ0bIR9NRONXtTIlNQhN
b+jMEvJS4wFSGJR9AgKIjK61Wqd9CNd18mysorRU7FnRc/70nG1rKciGNqgBjQWs
KF6BlKSgemS9RPS6+zx5D2vDL71+1/4DR2vFcxfXkpmNSjxDqplvVtuuN8eb1j7c
ZA4QoicbpsRqXsIbYHdLMGe+X966A1vmWUkFOT0hHiFFcCnM6HWxmsXGExR3aHIN
1PHP+zXNmzFburxVHQH6ypbjozDELFtAPJyfQISf8hwwX5+SW2MmUJ6IcUtTQ/gZ
Dm4PCWLQNXKokUydjh3+oKE4zPXE8c+UALaxuBy5wMSxm9TpouACjkW7mf4D4NZ6
HpteKm7L+XxcVpCVBeRopn6o+5rIxp+MyNenlZ5V3vKdo/Oo9fDNwget5zfQLGrl
+abqeaAEj1AyipdaQdRsMJFyp50HO7nCOBFAxt3vG3KgEzDMJYmUeCU3OFY9Lkvx
qklBtpGDDTDCPpaJd51P7A==
`protect END_PROTECTED
