`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiHwjMh2iJ2F2yiH/3HY2NEH8RmnoIzRpkdBm6E05MPwZ3skZIu9pmOg/JVH8Xl0
6ltMnPrFFGD0SrcwpW7oq1dKMgd5Kygkx303qUTbGd+aZEMv0VOOQARYsXNuF87I
Z/AfXH9wUDlE0M83vwB8odFkHmWbPdl7uh5OgOmoPKSX9E59tuV0UyN4peOXFXeW
BdYyrFLp6VwoRjWa3wKsDgHxe5UP1Mpj7N5oZiqmOw91Tv+NiWMMEIuURZtLkvMe
LISs0ZpsWXDiZPnZ4WKmy3KL1BhToqLQJKKv+DsDSYZej5o7AvbGRGoSssuS8+f+
IIQMx8k8ZrWOIb1CnMCPLYd6h0kT/BZPZAFkXPn7ltSNa2cma8d9zR6Xyv9l0Jfd
h00mZ9Q+UF4UFzMqXsP8YWel6L83K/b5Tw5LLCXMPde880oKTAQcxdIxnBE7eH2/
1emBYVzz7rZ6TiELgT1p+Mt4ao0ZYXUabwh8R6npgao7KRLCixjOkE6+IOu5LtG5
Q1iwL+6XFzpuJr2p0ZYCewXV21j1fC1MAsl9aonZw6IFOwZFoSqSjXpvLmmcDLc2
QLuaFPC3HkL4JhMIkCcOKa5UqNQw84WD77MIH3X5WZAgXRCGe3YsSscoYUOpsxaG
DMiVt8Xi0UlUsz07cZs+8g==
`protect END_PROTECTED
