`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5C01q589ho+gXGrQN99f4LqAs6LFq0zgp10+uxzVaFf88tQo9oe8FiiWYv2hoGS7
DRVfd534GzAQ7CZXghw+H88rOv335uWCM/8bMi6SjCS8BFWGb/cmm5UAuoLWndQh
8WtACzq5svM9W7i6Fnm9/cgyVmNeU0LaN2cc2xhMV6eRm9r7FzaMPDndXMTWXGDR
Pp0UtuzZu7jnDE9/vOPYXJXf01/jecgA3W25tuOlQb1FYjSm5hplhUGqw0zi61x8
53NbKSYWxh2krZbEO7bM5FTgD2fLikxvWM3RHGhp420czdOnsYPg3lochmWlGaDS
3e479Nkj9jqsL2KdDXjFNn7NlP1imV3dp2sU8QvF5mjd2dz3U0HYLY645rpC+YzV
h9q8fgE+EMEoKfSOli1jzVBlhjHzWWVCDQgyE3Ob8IHG12UMvSu3xgmWWLHKNmDU
QVViF2LBw0tQF1xRAhzoBUcXhMbYvRMW+5cjuTWaYlrbxsO0rzRS2YTpW3sk3T6N
KPsWgKLfa84Xf0XPeR7Cystuy7vchlZoLE6Egy0//LAYLWWWxYSwrYG6m+XI8Bs+
vF4zcz3jR9wfoPW21pAnKFpMTvxZ+wez99kPipqTMImSJeNL+9F1JfQwOhYR2eoB
yXuknOqJmTxeFln2pfySXbxremGt7Q09jmU0MTKjaXj3zAbdN+H7PitocHx2IBX9
jkQ0ZN9SQgT4hmnTT6YkfQ==
`protect END_PROTECTED
