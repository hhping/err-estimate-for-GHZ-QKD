`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpQKlm8JoadkQVJrkAG4Bezyx1xCGQLZnUKhMA4C4ppzKbT/umG38mBAZjEF0K8k
OXjDMLikLTWFUu/ZDghExc0qVkfms0FDpj6OYlofoByAB90W/sWDuFhl8OzTfMNa
Vn4pPJLdmqEfTkHhcMCWgOPsCPmO1GRCkpvzI9w9yiyle5j2KuOIj6bx9XJV6DKb
qxAIooYW1LKWz6kTGejDQbZQEbjKRxdU1Db+EK7Na3EOJTvi3ZGt/PjZw9+ob6M4
JriC6Paw5jdsLjXsvptnT4XDoJr2yL3MOB0mSKkQ02qkGZ5VRRBq28NuYw8i6M18
Y2qfExm3lpx3HE6+MVfcL2hTwAZNxnu3hW2ejl06l8gUaIlfwS84wqTpAydxSkdb
7PT81bvquvinund/6cX6lIc8ZOV4LVefISUjU+IO44qkZroAzd+RBEhfimL87jWE
DTvfuAbbclEUtRT2lQuFH/IvrrXGe5APm3E+9rmN9X2ucJLzROx59ZHrskMWegZz
Up6X4+vZon9qJ9hIRo6n37NG6LNdfhlyYQDyKl38m2h5lBhhVpOwnWmd0kAtbcbV
3yw87bgHP8R44fXanHtMybAL+aStmpYo6mY4dtfMrPreU0kghJMlURvvRr7w1cBx
1MZJCyWHdZNmSsHP1nJcaC2oVp6FmcoSL8oTwc4CBgvehrBGoJW9ZBtoeNvWawt2
hdD7EdzvI8TSaV4KPeoZKRkRm6ZxNkSi8ql3OiACqFVQHEEDBSFxH9LD80PeGR+W
t6ZpgDX89paNhX7BwOOp4krefqqvkyPlnVwzBCUltDaVyoMj8PySYfHg+Gr5Vn5F
kTogooIvH+570hDtHJk7cCDtTyivy2ODEcD7/WAIyoJ2GBt5aUMxQNRrfK/0EAA+
hYLoLTcmfqIDwtaaY243pj34gFVrgXyJoPNm/Jy5NU6W7VVFnu0s6qkW4t6Ql8CL
u/ln572K8jVa3++DE/R1SPuu2SSTOcKOKdGjPPPB8lXd43DHhHdsc+RDM23rnXy4
9orkuOhxOYd3vKBZn+/c418GgE4qROOAzKhS4Uaoe3lazVP+l165fUEcQBwhQo5F
WhT5K0WMaV9PJL07WVkog9olTdIG7Z1S7FLw+37QyiCnlIDZN1nCqIP8E/Zm4wcW
+OaQaict7xP+R6mWh8cQuSMbD9REwsabvxflb0bY+xWeMgqwlp6nW50GgW2ZKE8N
cgzuW4If37YJPXm5eVyL08+gA/Q2LznRxhbVNsb7/3K8dd8DpNjsVV3JsjzfkQ2I
I67N1v+6B6OdKzWbNFmX9k8Lsql92CKcyf7A1UGym475aKmrM1XXJ7hIC4nwPkHQ
ALluWgLRKeA5dX+MmZ9WCc9QEwvAuIud9P4+oT2tRL9KsAcp1E5AZhDUb/2Eadzt
rglQ4407ufHB+/3s+z6GhQDrSuyFapTQN2KqbyjXYJ93cEkr6yGaP2TUyYR4rqdv
FKZCNL8VIHGmNdxFaR/PfN/0QshGDn78y2rqrzSusaVzlzjmCxi1iLzKPIOmU1hp
kNNjBOo7S/jkh5zsB8cRPxr5icMvQoiCMJ9BVuytS0FPJ48u86SUc0wUJiGJet2Q
c5BI2vOl4y5bgd/fRqeRNKhu8vmyc/m7bfJo1ZD63GqcBYL4SPgficms7zFUi6h+
+iUXfqasJcjXr+w3FXxhGC3iIRW4ORXnHi+gdNLDrDMkec231wwrwymrUCyKf88u
JtKS54LUJ2tzRlo7v52Vsmt3Wa0YcCtwXHc6uqkn5BAobyIkoMkgWPFivLL6wYzS
ev97mbMlWUOKa+wmSULpONbkrHBWQVDPtCof8od6jVI7HkYcpkKNwCC3u19MrhAS
jQzTE6w2rmukJ3kcTJqqFkVsvBrWK5mpX9RGFMNgYSDdZ7bLNbe8xlxapMk/Wilq
Cxv1JgAbgYTeZdSVZCHmVFpWLCbxaysHw3dHC5QirZa+WvSQbmgFNz9jOYmSSgCx
AeYLZf9nEPaDQmppsnLASnO1t/5lDOzC2Y3+IAOMS2MKQPPwSpKETUgEfzuDOe+x
aSQCUWT8D+y6Sq3aDPVnHUefc5Wg2Tnzo0X+wcWNDzIuI0AdM8aNvbjjMJMS34+T
9N9Nv/V2vrrBcgBKJuvQCBlidO2rnnAtC5bpV5vhUZ0fN0t1JH9lsho8mDkp+l6J
g4hy/0eCyDM1KExDi47G1S4ACskEYbOurfwrS8S9g0rkEuAHZr42h2mNj1seCmI7
tfNolwcq9MOsx9qwP3x21G3lyujWzDbMK6BE46wjl0K6gXN4QItpF6F2ykLvRlPn
lhaC8ZRJpE79vcNj5HqRNAaCZ/5uL2SDRXRwciG4WO7NctDMNZzCQAvuMliqgjaW
w8mf6Rz9OWzwu8ky+xWz7RH5aZI7/Xu1hM2AOUL6RVpwe5mTYMwsrzt9xkL9QrM7
bprdlFxfv7i8c2hL8Af6mY7rlc5Vh5BgQSaGl+Vf6uZmqUTVmaTtrI61aaOt/Lho
N7gld7oEt30ufrDk9JeS6DZ34HhPS7YBIfwGMhlO8edJpWjbrGi0YsYAiVYYLUni
NQ6U9KsARC7oKxvutqOOPXNeiyDTPVu3btUg9FRf8ltavKtktcI93/ZkRCCRo25g
Di6jp7esD1CcTJndtrptsQztxgF/pbQSblPMgIjlFi5HGn/Bx+qS9xCSF+RPawUy
YECHHUjC7SehD8Aiyju9mtnmtWj2jbaB9S4Ve6r3AZN23LUauqIGBVDBKO3ILNDm
aZ11KFOnLFj1CkyCa8UkxLd3wnTPS5QY5/WsNIGg/QdkpHNEX9Z8esyxAnzI508i
v5ul4IoXaf5Q+ciiqS2FiU72o3Q1dxSQQw78wT1oVRrRL+8t9otQGuWW6F7fP7ar
Dh4UaPB0bzAahh2jNrf2j/BvwA+kJ/DQCVPkl+BZ0M0CFqFON0tTrB6Aqs77XTdV
gncp9dy8pMD8qk1XZBKT9poaVUG0K3mYBzaoKHGWDYiJ2nU6vbWQS+wy7Xr5/LAT
bRuRhY+xqCqQ3BxpiF7ObJA2621GQFawitGXdofJX/HbTDhzzn4xgIdW6poF7lP5
biyMmwEeXDPYSxvT1XNpAWNfDg6PbGFQRxTJ/1jG2k80mT2cYeVDi+PjshETjtyu
r3JVUxvlG4fivEAQ2EcsClIsympEPa8GfWzleeN+/09t4q2Uy7lrIlC2Pz9tMZBG
YOOLiH+KUK293PwTtPkZtbcOfZU4tpsPSRWHXGUCPhRCpFj3Utht62+siYUJl2Nk
I64oCwYlNysHyCm9LHQ66uHbIH1nLEDxuOi+nLdUUbKjsSCgJnYYagy2YciUlWUa
V4MtZY3aVGsiJgJgQ5WLhhpptwmSkocjOrWKgr6hc7EB1hshmjaNoktVjWpVZKp+
6C3Weh9L5xrHCtuAFEhoCmR076L3eNoy7eyyKs4WakWyzCkFfj7r10IxncWSzBAx
BWHtgzTsbdNgcr5d3EpT8XyPckMUN3bijRCW3Q2Tv76zFs59V7U3sIIHB/S3Bq5J
p48XE4orrUnObSUM2/RkK96bUrbOdgayxf1Gkdv8s5R9kRyY4m0iGzeWX83rsydC
OL7pybp6ziRWEBAQZxcwZkGF+RLYic9OwPVOH/MpGhpKmGmS8Cq3a6CIGlwycgG9
CI7WqgYXQIb69zjrWiW0dU8ymqlb0Wu2Bqh3RK8XPZS/2GlDLcL3Q4XBj2cYKCeA
EMGk6McXaUT9o3TEeXBLYC1Dg/PKwECADNKcwVv9c8KYEWltWBa8l1ypBjb5kEzB
16QjJZFhijaDdfTHfj8dv4YqqcHWvo2+u9gYjCbjTS0JvFQEu341FaGVqNeHcPkF
joKFLRxHRxKK5Why9yHneYODr3xjtUpMv8KKIkR3jERVROiVVm9ssYxnOfbHuKEN
NZAnDFrw3r56sv2YtSdvynHX0/mxptHq9bQeSj7US+iB/wQjotAKFdXuFYdNybgM
SJS/0BjWeYLJJviLZPv7nHHXw5Q+dEOzmv7KMYLDdEMVqVlX55E02badjyOS4+iX
eebN3AdU8yZ32RyTayBS+z+AUsqd5aUktyVq0UE4rs8LMEWSYY6JKuUmwETU9emf
0d6j/BmCk3lFo2tE6vHOstRs9/iqzxufRdjBWxbuAjgm6ucJbQ9sIb2sodW74DYe
mrSeLR8GJCKYrX1m9835hrycfqF9FnkyJtWy0FbH0XrWbLWmyypvnrYEv2B76x17
amZfhEu0l9mv0onbB0+r/L85Yk3hL7DicBrGg/dixSzDFMsKEagVB6pOdRT0DSq3
IIAaATgpX7PIIj/qSDWziBtOb+o0IwPFg8TtyKNPFRtbUwStffx4eOGWK4cluBKW
0Sd/IG6jjoLTL6o9xEEhh9KkS21rPVkEHqL0Uw4mksA1NneXXrDDrDH6RoBoe3AJ
rhPGS3WG8vdfT8EYpENqerFfnb3HRf5Nj4xEZo/JytOsJOa3XNCbvd3lwityvLEr
GgD6U8Blay4JumfJ1mpKcqN62ItGfrRvA8yvkgXM2HONgzpIIGX9r2jQJEGVvrla
ZilvJ/6ci2tgjqCsFg463wiHVqpadUjBhJlpPyFTGCUqGwCJnUzrYgGjqjx+D24X
8A/q+hy/EFM3IZJGg7CRogeNmXkoA/KVui00VJSTSnVv86vIlWJV+CZIGsa6ikZ9
F/IlGBfbSaYO52J+Kgfmk4CebrWBcfto7Pd/JiSn7B4EyJ2TMSxmN5f4Ecuy0qLk
HbtWxoJ5cK26mdPWY0d6yfX4h5osgvBnc6iJzVWYOzxnbQRbUk5VehPCmDZsbldl
YoFSmTxG6zhiH173O3IBaLFTNbP6rsdx04acv0YeGjL+PnswoUZRZW9duttIbETN
nGTi52BZ3kyJz3A/b4Y1KrZXNVoeJ4eQFJi5/Pg3oYjOGQI/79wcOjF7L09aH9gh
+llFSUUdXrOITdUDw4lZbQ==
`protect END_PROTECTED
