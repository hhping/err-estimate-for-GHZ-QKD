`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yWRLJ3Q6DRqlIJjghNZLc0NO3sQTDnxk9ueL2s08HW8X6B09+FiwYVK7R12ZiBT
dx65j4bQQzzaoHS98tC+NaRVfNExr3+YBVT4OCPSAc9T8+DFKfGTWlqxldM+8D+l
6ftCnrkdYKybBT/9jZloS8zpi6N1xjnk2Vwtxu+mV70vZujcsFkUDiu0pABoQDLx
bsaFN0BdV5xVWnKnM0nfFu2F/puqNkszSqWXnUwoUsKxLrH99uiusDJmilqUZld8
qyFKbWVsdA6EJGxxqvw0QHAWWx69bxOT+RveaxkRKymXA2smB/Q0SxTBJKIBYR4b
oFs12AwWIlxvucoNh8xXOi1j1makW+/8jQ6KWhuIubkZYReShEDkBmvqPXBzIpNl
A9/9KuNR2wo4Gauq/VDYFioi+x2luPhSpce6kidSECV7ctduv/Sz3dIZOwDTdnD6
eyNQTl+oX9IMY2X8dYiOtt78QPPgC7Elh7qiMqDTmvLur/Pu5Wps/8T+UR5yO0h0
`protect END_PROTECTED
