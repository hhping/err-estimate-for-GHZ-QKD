`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iM6bRDRNjBpakJF4UPI5eHiiBQWYufYsgO8tn3B4CE9uikAhZQxpv02824Kn4xEd
OHJQ9Lttbddt6zchCzbzF/pQfgBaVEOR/+TJZTvEtZlpLYGMcmegvZ3/aDGSgknO
iaNssbBjsboN9SMZ0Y6J3nBl8fqjNaVPUFMppFjhBncQAMwKpYKdVqor/I9/X/Dp
UFbjVaX6cBEDUHcAUgFrOfI7AYogRsjnTRBZb6gmJGa7TY9d8HO9knvR/u1rTF4f
5NNfMmAjRwAiypqOa8VtK1MdbTbGn7pvwmAt77BQiCYwVmitAtHX/YZ8Ltw3XAA3
JXIfdze9gd+WLfEXvyzrWWQIZvy/4N2gYJ26KYV+Yc+5aFjzuPpaNUcGN+cNfDky
YLpPnjMEu0My+s5oxYsyzPSxARvExOabR13eHqq0ttI=
`protect END_PROTECTED
