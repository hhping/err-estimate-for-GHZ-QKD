`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+JTfjC1bVL/OFQxHolsew0rV+68niEn1lK1z/2J8TV8ETCvCyUGAYVoVCVreCHjI
sOKiQhNC/yJlMUCpbk5zdf0u+NPSYzw3hz1SIKQfKr6pYFpKS303qBKtbKdrxzEZ
uYTKdC+7U9VMnzye945xPjsDQHW7t/aqb6l/pIjE2weHAE5tQZm2u3gemH1cUqE1
zi/q/B823ptfG2TnnPvj8tuuUahlym5c6Gkxmu7p4B1qQbZyU9bRpWLKbA8VSrcy
8KJC+n5O7Zq17SbjIHbXuk0Igjn9lHc45SJ5xku1LMm3tzA3Sryk1jdq0rqE+U7c
gjIjIcXTX+ZXQWQ7Z6zS0P349xb2gTVPT8RU4lW/ELfqMhf58UdUkA5q/2kZTeFE
AGMLvbAvUiTg2vajAiZ8zvjVO9PehG8qpKval7X4wZ1aucXD0sgA5FY91ul2E7Qn
SsOTK7XjqCVuz7LfZw1xz3b0pr4IlfY+WqTG71QzDC+EOVFv/lX2R7mltw8gxHy+
JO9znDipr/6uEhee109THud3RwPLdSVzaX/qi/GRpvbZ4m6i//9BeEmXMj0/vhyn
aV+JGZPWThO5Hmi5UZTc2BiQbuIuYfOIuB8FMF6QJ+I9IzwqIFnt4grdbL79DHLO
BEFE77hV0g+cGp1h10E8lS116/fRz34XKSzAZgfJ/Y+OqTvfYRNRusyuGjX62kKy
VG9O7gl6qQkf8478rbKRopHNzodKDUCXmOq13k9XBWcrVKlONZPAdNixJXe1L9PF
yaKEQfRY2rI94GMK1njpf6vaNx3SvfOYM/3/k5jnI/xfhCD9SNLSESXfBN3/r2mJ
9/u8au9cpPwKcTq4uN7ZuPlFhojYLyPPxWCq+hFZ+ldC/MEjAn9UdAEAgt9ZokiC
BINhqlHlSeuRopqxGpil6h3JNF1wIiRqG9fXzDA+aqtr72oyx+W2V5KYSkj2ndzm
iY/E2DKCOE/jjdhkz342NRlP690uKIq6yeenCySSDeT5EpsTklRem3+IyVVKwnfc
INd9cxiKU7Kii6fH5vX1XFb8J23r4RRxEXi2LGC/je+FJvgZZgx3Lwl+rkWDH/Md
RyoRRzxpT/AbcfmyzIkOOrCc6HogLaNs+3ce+123utabcH5EUupYzRH1OsBYkx7o
cGWzU52/7MTYmlM4kkEOhs7PgdsGSb5LI5UWluCtZgbhGKIA7+fAbcpnFIy6mUC9
IU2c6LJ4n9uurr2Zt852cV6smdYCmrq8Uch8vffkp+7L520l3MpaLJS2nAAZzDGF
J56HrYXGYyRvYb0XywCeWnZYUHT6w01ZYs7PnNMtkXAL20opRUV5lEUKEWP6/5Pi
`protect END_PROTECTED
