`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v/a4Bg0aAUpiEmkCPBZO+lPZ1ux5vicXYN9Hh37EBhdm77L67AXEE44OsQij00eZ
XzpvIj3gzWjBVqt3WSCunB4RuatUTn5U0alnkQHkhsk6dq8324nXihrG1jLY36Z6
uCrHMn28pMFppMI8za0oIVqlE1jyWuO1C3yB+Vh+jU7Kt/JdtwdEikSqxebZieiw
CG2CZfWAjwTbRUlTqzWhVYDF/+rR6crNkF6KogVPzIB1UDQP0LmL0eXMOGSe25YV
3Ql7DICVpI2tMhDVYvMcnX0NqO96mODdAoOn9xS/kKK11NOP3a2v+wf2uGPsgxZf
e76aMrJ4wb/ITGb8ACVTp7N9nhAjyfolySkRtIzJFdJbVcCLs4eSzWDP696DRH/H
KdfkQcKZgpr8oFE5GW1n/nsErixHnHFzbOSzmv6YbEWrXz4j+YRZfffVB1SlPj+j
OCgMFtFYyRihX2j39CT1LLUgu/K1uFowSK/m82d/qjrdHf83msHOM35cMXVviSE5
6s76wiCDNFQOaYVXvpGTfYpReHjLOw5cJZEYvXM7r7EDvuDemrF9jQ3JkdGFEW39
ckgNjYoL9GI9xPIC3MwZ8WRad39TLGk1DBjM8FdM1WOqQ3AnWWdJ4F3AQudk//RQ
G4ixDx1gOR42tyyv/io714s6GwF6Oeq23m1lr+nnfZoDl7JT5xMJHFclWGJDmrCi
Ge2fN6B2kxrTl+VPVx14GLTaGyEENGTUe24yMIch0km1oCmhcZvrLf5xlkdG9IbK
k1biZHy6FreaDG4RFcQy5+l9CWakFUjG18AyKd9K8eCwqLqT6NjBPGlNtN6YpiWF
qMKlUuc/0YSkR6hRMhqhUzjBPDL744QBQ1KG3kyIVSA+G7s7wJfEL7UjVwChPENA
9fqu1ODl+uZxvyTqWLcrym4EoLFQV9ruHMUv2S596AKEbZZzsQMK+DfbZJMxerQy
qvKq8qGk1VS6zNgQ0Y7NEiur0FfwSe6zQ2rUgR6l4JlRj9hog8NH1aj8nm/uMMD/
3oEvC6uuvccT2Ya7smB2FhYYRmrMHMKXps3hLBfnJh95tI4ajUg5Oc0iljXLVQm0
WJhBhyQBg+vfJQdBbnJe+X6DXcq+p6OZVS69HvVs2DFAP5RGWBTTlcbRvsA6IDIC
M+d8qkb9fWNME5Nf7xk4jPG+tmyXFngEiBHajQjZueg3PbnA8qt5aVfraU5D+h/e
bV7dlwwEyZqaKCesh5YWPA7fm4/q2XGEJ3zAvS4bbpZwZAkg7QtDOJ5yrUYIjvQf
gofriidh6i+6DYj29ps9pAwrM9gZf9dB1tAZHQjK5D7/v5LiFifOfHyRT17dXTvR
3ZCS216CQy18CKzMQaOWMSevQRkqZ6DZC1jceFd+H9fhzqdRair/h0C6Y3mYnz56
skRIV/DO7sEK8wmMJJ7rTqsLbUPnyowCt/t0eUBiFJFz9AtDXFlG+72imnZKbdZ3
4/T4ZfJxZ10FboLiJUNqmw==
`protect END_PROTECTED
