`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RiUpLQJfpjd6uDdPrL1q13kvhcOu28/U/RuXWYmzq9so1LhlxGgYCRDrqprirElp
ID/TbFxYTCM58kGw9o/NkYMQCNZ70ddxstmAsbl6hfUFlRX4tsSicFfNHWVD4xK6
TehZHNrILenCXL0vGtScmWUYsG3AEL/oeiNZwL/DeXdviett0ORhNa9ITDcuY/yh
CS71Aj2K3wY8DZiclMhL4akKcfMIO7Or/hZ1pFLv6seYUcGVkQxPyta9XQz1h656
9u+8caJ21Gvl8gc2EPnq507dzaGzDkKCJHYTw0Mf04gT9DHy4/xUu9ChLc0FNILn
+tZ8GfkElxIUEHIPk03SI29n2hobIzdkv2tyI8Krbf2niwvLNVFDGpFfF+cB3SSc
jWBttbvTyHRgYwRE0irsO3cBPp8cSmXL47EIdBiSXVgpbROr2fhHpYwFY20WcdD4
BbstXLgt/7yvJjv9SvyqVP1iij4OEhg7s9CU46Sc4xIvJBh4iH2cPeGZ6jEAaByU
vUWFMKuQ/8ICvInAnJwLkX3jIHse9hyv1Wddo/4lMnDWTnFhwsmtAllpk0KyVoFm
JpuSxQ9wv5FXaaaIk9POt/nCRdVQ5ITh/r+Ao6HGXipl1vukTPziQWeIKpyjIejH
LSGselSnREsFDO/d0uWTMr6XuSeWnt0oLXmVRH69GxY1yoPaCgG0LkUtnexyTshJ
xOW356ByLoKVflqxCmou+QfSoo3LJgqLwTxJaMaaoNPZkBDt0D8cZbbp8nCstZgy
hOaDaIzgPMCxOQndRdhDptswXQLEIKZOJhDYafYcXiTA5xnBfmOvVaikH6PjyQof
H43rx8bxLL5SHxfUh1jXeJN3ReXOaHEIJ3kbV4rfRcf7Myhuoju1Vwu0LLpDTM15
d/yFhK29eUzZMDkkBS6ni4Dkx9bFlVvbr+0T9DEaD6cXjiWrli7+DqN7lwCe2OAH
s/Y40smLP7RwNzERk2QIg0HvQEjjyiT99SqFrvcDwsKMSpHLb5Mo9sLUqp7Yv6nW
AT6hmlJl2MRxbNWgxy+JQs5x12PgQ1DsD0U9ic4Cb7KKHbFu4zZMooyI6tyazbOT
r8fIqTLRp2NDQNS18ByuHH/K3X2JDKVvKwqcDV44Z+T6gNeVF+CsSwix0K+WbtgP
4BICm/MO2i0wr5H9Itc7BPGWcu4fZcXP0fTsTJpFm12taZVcojHyoStxYi4kRx4j
jsuqDLtJtcizgo3shjepC9NFe6LjpuI7eTgsJ8U6TlDgfN+sr70gkqpE8VJmThYl
r5W0xBnlEqq3y2sRZYBKPtO8jvT7F/b84lMYbr75rILF6A/Kp++IJ+dYdNgQjWvB
d69YI5z3JEXaABexP1EEdXRvsd/9ycd2yyY+F7lQRqrphWqwV2A3RyuMXUAvMMkt
VTL+Hekr8rspC56oqTlrjDypQrNUYOr/OUzCZoYlqTCNq0en4AhRnCpAGNOaSIoZ
kW31RrtvVHoj5EhImfTfD+0KMjFcTH8el0fSzdYRL9qRdqrj0udv+sCjcbe4ZmjA
zykr/gw0FXQBLp7wI9kyCpKXtf5FF4D5VPJBeXBsbsjNtNiIk5549/HfZW5JZd2U
FUGK/TKiscY1X4a07VU5oW21J5hPByRKF+ozC5O+QXjSDaZEshgPka+Je+JGBWmC
b4oAXGGyuMim+Z1ecT8TglVKn0K5i05H25VEkKaAgmZcxJePuZ/E4TykZya99tvZ
Vhc0SCj2AkmmtCuYJYTf+VJYVPyaPqEgUKzNNu2AT8/QBEOtyuv3uy6V5aBw76RB
jpNZwqcJJAhwh4RVzl7w0OgrgEgfPdsz2u4BWDIIgA+NPG+cdos+wSIzKbi8BRbv
uB9+Ujy3iVtHeul5SWbIBcxjA+tuRVZVFi4v/AZRWD2vl6UMG7NMlPYHIWvmfzo7
SLmBMMbfZD3YCsy1qFffliu86PlfG92SV/CyZXKLExZby1zXMgpOG3Y3UXGM0lPM
5SN0ZNxq1B3SLk3/yEAV30v3LpPY5/mBvYi/cBIyQwSonjGnFMflZOWPk8/OtqqI
4IlbDsn/w1hWcvKXDBeBiPU9ro03WEwzBEnYL5MyEQHpQyeHe5UBaMztDz42s3WK
mIepsOv6l+YDWECPoqS19Q8AWoNZZIR1Eo5U2/jRIJ1EbaZUFzmkv1ZC8XSYgfy7
tUTVMNF4/WmnTnnxhUV7YXjIf3Z3i/MrxEU57I2Rg/uS0xjJd74/WpETnUtd0sbe
sALBliSpZN4bAwlBQmM8qGJIbQmgH4kOCBQqY/sFleh7jzPwDtHg9HRpc+9kjOB9
zoTYeuh0/mboQBXuTvsNd2Ebd03rNscbTRrV7HbM6oaJ6xunZzh0WDOp9yI7dTQV
RoeJHFFtiufiAyL2VT79jwij1JWODZVZVyUI0DJ2UyWxHjKm24fg1E2WeyLfdEPi
7MV8Tiy3tsbavV7SN0yNY0Zg+EiAPMgKley93x0hWCABs/os/gmnNqDGjI92P+vB
9OxIg89M09jAVrR53mNdVJhAZRLso8xoMICMBd2Qpnp2dSHxSVLuJ80ZYazBUsrS
NsKtsvayFddnuyOVBRPaORlH4McpIfc4TfCF5iQM42+k6qjwWG8U+5pla2DH1VNA
HBNN3SiR9JKbgWpdOE7a5dV/sjezO4hiNEGkHZey/vKVLuKXVJq9PXbUHy36b8Ct
0N8r3LgfeCgVEEgMNhUH3b8OjORLVUXSDdRjQiHHzzzGmdWTocFlJIrBFxYd6W63
iaYJbSUzS5rP9oufi4e707+Ncz2btn811IlCE0yQozLrY1i78+QMZr3ggjWFpidT
LxSlaprrsyHovN87UniMNVvZrzvv3exiynpRKnr0eRRS/AitkFW3LQCgzYesTv3m
fIg85gaiiOmU1L44foPKK/Tyg3WRV9webJInZqHSbRsx4l81J58jzaCNRwRO/jfT
YlFINUe8X4RSF+mvZJu2Z/ZBd0vg2kFFBzYoijI7ktkSVmooiyP+C5oVhQ1AAKt2
HJ7BIQqKlBrOgt4oGLNN25qOVe25uReVCsTc6sSRkVFKTKZ7hsTBxurzSsY/gFjz
3McZS91HdV4ZQwbUqSlgyhpWvaxm5Wb384uqv49TuU3aP+PaSOrcdxPecra+sBaV
+SPcv8alMLm9wfD8h8YKlaHZH7W8VXwMbKq0wOCsGyJR7C5sy5oJhZaHJA3laKse
dEy3Jj/QIzCvqLK9L6p9aLzdpJ6dgzJt+DxiviiLy24xDr/oB1iH+DqKJUKz/HLF
G4C7HfPN3K7eVJPPSlRC6FzOZMXEIXKVzFXJD+HmY9uPiQ4euly3Wc8dQoN/L3Uc
NhuXQedrFEvRp50Quv5h1RVaDodcmtVGiuEMvuzpZMkPf23Xvo/dl0isWUY1JrZ9
vv/SI2pf/J4YqTNp4/ze2NOhw7XRiaSwlsQciQ8jY2OFP2Y6wxbw0fAw4ic0bb67
XtVD1T+hoQ5penkb5IsccnaHKlpKonOLVqHXrCkKjJ5EkSlT+/wodD2+V8BosNw6
lwbYax9L6KQMgb7/+HSTotXnMdiWJZfv0+O7Ho1p/87oZhydT0BAuIDBgHK3CS/A
0uW13Q4hWippU7TkzLh/tQTq/+/wZ8fGB6ZvU1rToat9RBpWt+5+vYorYPqJgwNw
phaPLeFhl8GWiUq5ingAiTUNIldAi9XasmhavSrNmbxpx5T5AjYzYWuGwdZXxIEo
JLfzMZMGHLOQxG0k+4lwZrVOjIlDblFOULKrOs3o6iA59d5bCeWsGfEeAViTD3vv
eY7/2uBAn/M8+5QwNfqJ1Nidyw4A81is1SbFjdb6bu1WCSI9SCjmN47PZtSR6EGR
k/rPAIV7cl6n2RqH24TnCC/qYugWQshUGBaRokjcgevsu2zpijBZTa/kW1T2M7cU
j8G61UPnMX8tnXNQCw/toPkH4YYf3JvxMc7/nYswRGGGeLptW05FKbbfDiz3OjZI
lLgaji9owqQt7l7PDnYuqsvRpZszyStERMowMUC+Nzbk5qfyD94pKFscQEHUkpuD
5uT30tAF6lRYFyUS+IgSR1io4utBPx0upHUjL8Sq+jmAoiNZaf+au2VEO0R+V1uC
AWD7BtKwABEEmRiY9uxsrbCRPhtMxffcdRnPJHpeoUCPNr8sQ5xY43R25czLfrnj
bT2hluQHG4L+21KfUSMqe/sXwIxt08YsM9//ribl8fGUKqDH2Ycb93j9A6VcCZoA
7G3j2n361/MwOI5eEdbPK6TIwhx38v8F4HXrjnhg/838MlUKsFAXjUb3ZyUa3Cfv
O0lP/OjvavmmrIS4OGBOxU48cjghZ6k4mI7v0QkD42tck5B4MoNrksy07sbZKii7
AWfimE3Hvs9qTO6bW/75xaMF/VJpA7cbLphNFBuK1NIIKASKDK4bKQqXI+YETplC
N4lbavt7gywjG2QlXsW666V2XXMcpATXTs46Fn2Pfw+/TnnOZfbmlO/4URerTsBP
qYx8JiWhpr17iAAB6+WeJH5R70N0sfR0hChIp0m5zZpj7x3E4oMwsLvs5IbtN2JL
AB/bjKnyPP63aQeo48UPdjEmg8sMGYAuTC4vDQvmHpgptJHAJ1K6rUY66L/0TrrW
2s7VsGTswUtLGR5v92G75ZOKZDlVD/DK1vvNXcnB/IL4TyVG0hdww2gxSvWyYAzn
lTI2/gBeyAi+/zHONT30xA43GdKg+GP1z5arz3u7l4ZPyurpYDT2TY4QclMbmoNF
8tRMRB1YfcYT2r6D78XF8KZtOXlfxC4iVjtBky6qBjfhKn728+tMUwcXG4F94gKD
kSnOip2sPfNQUIR5W7TKDzukDwe06pOy7Eo+lHvbTwEb49n1PG/xI1TLv2bv3e0P
ZNqk4PTKherfWjVGLKb4ivMbAok99xBRewQYjAdvMkka8vuT4D6SAJchWcs5/M5j
ZriCbJm0BDJAyWfjLlqvnrqK3Aaobx5hN9mbF/UU1d/+fLRLmEPoL2Nf3VeVKAc6
k9Vmtcbso6B3lgguh0qHLCJXq512rMd5h352Qwwjw/a0ujek5EvNJ7am8epO3OT1
sMb/7/rQytAfC/GvGCyUB7ly2WGHAw5JLDkq3BOIkojio5TN0oRgjm6iep5XOyUG
losWjbvVQZnSOKWM85brArpRWz6Yn6Z4NI6WiI/O6S5pjbhKA4eI791g9z4F4tOM
wRgOBopDsKHfUK1CWG0SUSoy/Nfm3aciOFLUbalF6B1prA5iA3zr3vSUUsFwmFTB
UVW1FLP+vGQ8HohnNIp3pV5O943e01T30EBuPYhUBKtJwbvAQY8nm2P+LOmtL42w
1W6bwXg0BYkLBTcpeHf480f0z0jJP+dI1/jxSNDg53WfI3ZZKaehpK0zzo7+Y0I7
PvqCPt0NsDT8RdPhrmvWmaVRV7Dg8gSELQj3aAN56rjhOLY69pxpmo5t2yCey/u+
A1DZR7uONfSf4koTIOEczKbW7IHYwndmk0BHu3QYEQ1vwufWaGzpWX6s1+70T3pe
syjopgGBlsbS/TruIC8YQyyprC6R2vTLc43zhEt1fLeFB0iMoBAnMjxjsn0GrS1T
uktQqzqifTiuzc9PDgZRq3ymX4sltAdU+7Sjf/3ASjA/L55pEV2nNn8BAykYlAhO
xN0Ba5fhmPl7kLnmL4maXjECr0McQL3hkxYCGLzuUT39b0s2ADVaZcwZKCqNLnMK
2Wvne2TAlgK48cQ1yPM9i/bbst7hMqD6ihzmpEgtP0lM2AFmIJ5a1qjuNOx7gIpB
IOE0Tmu4p1NMKfwfC7rKUDhg3rlOWmvwkqN3g4CNsaQo+1czsHBusgqj+d81rXXL
Vfg0xMxp2yINxsaG0y6zLisEeqAztjT13VAQeQitcDkG8xveAh8fcsQdKNzgKpH2
qmbeNgS8xB2V3NHfp5lHPwR4WivJ9+NP2mIvzYdJibC5ggZgL8rJbfwTioBuGspK
t9ScdmFM6EfpE8dJRzZtpx6/Wpm6HJbgLk4Ze5De2wnTaMgJ5a4/z+dvuqrxnFpf
WGWx9Es4Y2WtL8TMXvGnMm4poZBM/UYehiTI360t04F8utZ/vF5e62nKYEKssbbp
9Ugjfh942fGIYmhZ8DQZUlJswbKKhe0Wfx+36oHn4Toc4TIT277lEwJXxLLQa4PJ
ZXxHg+OqmYk8lGEiQ+MYQ8+g53wFnFS9b0m/Ef9IQ2y8Bj/gMxy4ngeiTsY6plVK
nnq/dg9m0D4ay+EG01ZMFNfXBN4QCQi4+TJzy8FjJKxNpDpVw5bcw4+Vr+SnzubT
vZSpzPq7Ac4k/ZlW5LVyvIy/5GWpuZLxRkeYuhfkuUvLJUIeLwamntmR1RftnPuG
+EWqWpudf+CznENTKxlwbOsENHUi4ac4Y5sIHBQdoGGZhNOrzst0wEwSsDF5Fxif
LjRAmMbKvDEn2zCyJCOKsMu5w/fhYwe/KbE4WhbmTZDxeAAWL6k5tHziqlC2M3/m
rtzhqGSU7DmxNdr4AcDUv1M7tffvwUh7hFy2Oxfr5amdxCGRaUAjLcoVAPsRm07d
BauEE6YVGdKi3HL+jSWgGpd3dSH0M6kqQtZ2qASQ/DOvw6zAFxvn5XU4vnRcwg/b
hHIYHPs1Y2UF8cyeFKzo8eHMgibNgv0PHtqGNpSon/PQLrAvUkndW3D4CvWNPSpS
egzBapoalp9nLXDynd9xCKqHRxr7kHyW8WwvarFR6WXMH6GHkEDPUe9oaFaqb6ir
ZLPqH8nrOcEGZaoByXpLdAVUK0UgZoBogy40wuf/YWZm6UcgLzMJ1QLtYWCovfeS
5WOHBlZaZfoY7VSf3J4eVjwQM67xzpc2Q/2KFqaDlkPCUEVosxAQOQoovU0Kny2Y
RHlLUkKwNcm/4zCcI1EdXbe6WH1xQZhknF5PjnfPIfEminE7l9eHYzqGuub10cdz
352ahNHnxVTd8UZqiWkt5B1rYaXzG52UEIN0lhnuDW07fWpIkEoaNs+XHm0z0IPS
Dq4F3HYteJXV+Ix9kXEnCHlS7waa0T4Wo0N+zMhvgOrCuxa3iWnZLnHUk8rEi8sG
Gjjph8PCgEPXCJrXg4YFH7YDtR1BOQB/t2IMAH3LAO1azePkfEipYJsM4Ln0QC8C
9XnamcqTuG/XwSsy9jcY2imE1BIJxKUa6iqTL6Ed8XnqFauqSVvHcHY9UJixPNbz
MeJsalNsnMc0qORjl7d7NDmDhLRRYEV1TcF5AiKm/FzY248WuTEm4RlJfD+NOMAc
/2UY+vpseSyMnalMh/UwFAll3nHQzmGvA8nIP5DAVPCd1B2yrt0PsS9uDvCLprB+
wI1/mj5Q0G59WHD/GdsKreDKDT+wG0B75yKkgyYZD1POiLwXJ0hGEJus08xBQfi0
J4BVzw+X279/txUVpmfSYoykXmlZF09cNYS9Yy95ueUQIiwR6Yh4J9YgpSl/KWNM
9T0Wxu+8rrn0jJ5HVTuT7JB3Nc6BBI3ZZGNKQhmUYdtDI/AeUGFpwLwEbTwth921
KRpjdH0upsTiEAFjeOt4VLX/TwqpSu+fpb8m8JxEmeIL3FOvFbJyJ0wB6Cf0OAiy
wVk5O/7dOCPsgIAJx9u6nbLz2jIZx40p0gi2KRaKcbtVoP4MySsttc4pdlFHd4ze
4zxxzi2yxBAze6jWhGXKa055o/dj3eeJqytJXKxHfr8UzxpMpYYoEghPni4JBeNv
ADL43idZrJda8Af0wBHrBIb5v801t+8ZV2IHBkyZeb48P3jV3fhui3lE3aDTgclp
e0CKNMGmeNolcD8pr3fn+TlXuPnMzLOUU/bCfCeCMClodF/CzHaIuAm0BKh8ynXf
pKo3kstIQ9TvHcqfGPnrnWCxNrSZeLadynsM2Qy2IByiKVYKJvykUeOXwMo+bhn3
JO86zEM6X9HFHcganvUWKT7RB486xV/wgyDFWPPJ3ntfRphzttXDOYTwbLbjjGXp
sJupcYFsyYH+tEMPnUX7l/4w9TRk61Hn6P14+sI2+khF4PlRbP8lhNDolpZ1jBuJ
yZgdhZRt6t+Q+0nu38VSTtOANJ/0aGhFiipO01WWNXpZmmEDOjTONq3yEK7IqQCY
4RBDkbtHTgCyMuiRRDv4NI+sksl7/IfW5GBgqqga0K/1ehx8LgSgTNhSrafUSuIF
hxUii5uUYzBAeoeIXf+lcl4YLvSbr/lq9R9969uuEll+XVn07AGrlo8ooYbBQb9j
8DoC+/gxf8YC17ZGUJtcOmdhoCIJdzMnW3i+0GFEFDrFX4aMKzqsDHwmHN4ETM4Z
CkkN1ao2upSVbznslNsbP3dJYcMS0gLSC8eB9d+BODu96d3z24tyqS1jHRCy4OGw
/iucSSAERrHLOFQ76cYQSGDmMlsI/cx/wGHU4wUGbpIG2yio9LhlGzZZmDlA9ZZn
rNnjJUVEjdYmQffpHV6SN2Jq26AQ3D++lyG8f1wC/ErlVkuc9rQIZTe6LdWPchYx
566s/5rn0zQmOpjCxP4Vcfn+IIIS+1qAG0WdOdop8+Z4TEf1eTS5TfM782sm/9CV
iR+LNLnZg/JK0Hkzh3cXA+o88lPUYw/GviBM5fzxfLRB9WwKeGjyUkICg2A4JRL5
RJGQPzzgHzlHx6AsJTClX/aavriBEKRju/wvGPAOiwjeNE+eATDuyISyMGZi89rV
n24t2Z9bRi2eDzi3c4I5D4kEM5SUmPxiWtlmgU2xle1YwKLnr7ev3VJO6scgwWRt
aPZjdB/0OH50qSy5Si9tS+NyaemEilnuLczWOMhcO8+13Zp8zB0Ub0zG1UR0uaaA
7VFvR0lV/UaaENNr2JEulMuHVTeusEg/cVdRvz8L7lrE1c2viCIU7onwMibn930J
Vs9H2jJfhSL5SOnDT5JR2hHdirPOjSM3nV3aFRz7it073DxlY96wb7gR1OBIGqOa
RW39/l+8d0N6+9285mqPPGzFBCs9gZVxYzEqFZ46yYDx0UMgIq6Ul3+W5vfzTjU/
5YJJmnH2eCIpPcwTb3ySC2GJv4ZPKN6tAHVq/sqsWdtmgP/fvK6r1esUEusE1SQE
apB8K2PtFzPV5U5KzpzgDr/BZG1nQNTRBrSpLvqjvlNLzdi5CnPEKMQ/6SbGy1w9
XBFwGj8jBTRP6SPH6oKOMTqN/T3cqlHQovdsIjZ26XDlkKZND5JRoRJyyqb/Uwu2
QyAuLAKGP+O283AMSjgc5RdLPyZM0X2+lgg8E60B2CX1GdTp9R9OVoKeOeh94bc1
Ugh+Ou1eBgl5djyjWi42gJ6H+HCz8JMm9nP+c1pmQyFyI1JzF4/zQI/DT6srX+Sj
1WO5NcyDCB175PqiNitziP0i8O+KTwnsdgVlqgWAK2g7TlyxnExZTVWvie9vKwiT
47HZvuQw8ZVsipBL1w32mgTYFbmNrUXWDvKnn32iS+i/6s0vBDKvDi/vztZo17r6
E6q/7Hfi/dS626OBnWnlZ80eXiOH6ysmUjH1nUQLrdmHaMOtJiy/5+3h3v6nUz8m
vAq3iJXAn2faaC1u8UIcjVJYrIL4phuLVfTS9T+czuJXt4aWQ49EgVkt3/wJqop8
leCh1pjEUX80r9MfrfcL8DTUlZXB2iq8RDt4XawxHlzFxMn98yVX0HdXDHGEiofV
LGdu1Y0X6zTpTHYmP6J9UhBHvGKowP6HAwm2cN4z19ILKss24isDP8YeIoZQIcR1
Src9cZnJXKl+QMhFqx28KH4ud97GfnrxyzWip1tjZkZ7qdbIU7xchoBfFVdVHrW/
7sMl6Wk0z12wolzJyQN+VAb9ulPj73wGIcZS8JVD+whKbf8WVCR1+WcBo8aJfYWd
yPhzineiVy/UYtJE87jnT0N3iyabMKKSbqfJP+IilOznB81JjhOtltFaxr8j0wZp
CXq2upozMniJRjULyruANRSI9RgO27xMZT/yQGditng9xp/GsazJR/Plogk+eALu
bfxBoNUp2ZDtOkxUUsLVCElbEYSAUXYzEdz+R/gk6QSBWf8iLdrRaJ36YJLrNjAT
kIDS504i9nhExxULakGjBdip/KP5kUWI1BZ2AjR+nlyyBkqyhcq5PMV1bwZIw36r
uY2RrEg2d+ysh0YwqfIQoV4u+HtChHu8j0oKMCxGUoRBQBIEofBfozXzSHhstGLv
/7nsciy8hFvtSzcTeaZRnmRkQ3WfgflP6ePu9K1p5gsJECiSy4HOChKkRze4sVhh
5+PNvmA+1h2hZI81k+qISC8GVxUWZa7pQzRbmw/8A+rNNycf2YKrfBx5KU49eN7c
X3zUGjsOzxGyMSMERJ8PKKllnAL0MV+rbLluPW5vr3bzLx2j0HdFSevCzYydkRrj
GC1zVjHaRHweLNdaRRBE29S9xCOBqhZeP3IBuh/wKN/BFvAuOtW1KotM6R3x9C8h
8VDmfa8iCY/Vfo1+SAw0TzOcDBEcCNO9bwGDpHaESSu7bBw70nYY+th1g/79d0rq
rutos4EDGJaplpbM+P/p/VzSHZpiZooEj7LAQ3Ap7A7qXxflaDs8MMpxybQXk8vB
369nyY/PWb9RX7Uq+wtYDa1c9JYzWHPlU6EZkW7tddHg6bll3XEK9oJBj0MqRs9Y
ZhUsYLqQmwkbNnLGx9zfTSXl6STft5W1d/Ffqh6teLKtJeYsZGjpnNVN2MwNZKvt
DE1UTDCXDvv+LyCa8ym/Dzkxwn/uTkXlcMeetkHYioBFI0/+UYp2xIbeJKtRvZdP
MGaUDZ7Y45bzxFg9GcnQbL2jIJFzeTaWQtCCzjFoKm2rv5dZhBZbZzlrunrxTNi/
P5gpsgvP26aYgMpswCoSu3AHGtNr6FOs/OTgGwu+J1DwpH+pcT7+PFs/wQRLZEGL
auNgFVmc9dh1+v/PtGJepv+pRjE+UA97Td5apCwzUhHfdodctrxHdq/js6N7e1Fp
WywfeZ7STaOdjRxpGWGfvhEl3QtJklfp7vcRb9E28LWBYitkVkfEi9/wG1WuhZNQ
0Wj5rrvnfbW7GJwkben9Apa9J7//6Y8FEv80Bocwk8xMAm7OZqejmLI29Ad5z9ae
NCY7T4t1gif+EBX5Z3k7qkT8AvmpxNK4LHROVkJU7yo4BlIc5C0Ek4rIAEy+Hmcj
MzJJzErMA7FInK8UytLCPjOHsSW9S2T2mj4FWX7fYCAEqxHXpLET/wiC4696rzWf
APJtY+4j10omxfKGkZQtC7sDFmnISgYmhNgzKIUQM+W1OALn+10SkwLwrq8tOin0
L20quisSQtYZb6+J2BrTuADiijWxvxKg/+F9ipCibLcHjXI2wpCTbM1uyUVjTZq5
/MUz6TpV/cPKhngDXaXIdYa14Jk5XlAOIcU3cvH7Gg/OapipO9BXX//abc+xLOBZ
3Jt40YyyQEnqhbfkR9vYDKY4uoaNBOxHHXFdfeHmXiShhZmrcyh4bTR2uGZNMuwk
8EfKki5gvNcIWdryvjzhMapnMvTshd2FrrsO8VONSmnVoBOO+CdN9932XnyKfoKY
JYYQYCLm5oRu8liGIuBlr//ZPGx/5GsgqVzRitajUiTU5y1xUhSVfs+Bw4l2KyC8
2iWCiAA/yawbyijDfyNTP2D29k/kaB4MCmDmM2aTQyzXqT7Tsi4Wr3xBkPCAaZZ3
W73f6LVav/WMyijSZF5XEfaTosqgCqlcVPmriEAfmfaImpqPo6vVPl1QSZLYIXeA
o2Zp3te+Qr2GVIMqSIZdTXcyiKFjMkUv+uJ6voEL5kQmKLgMKbC8uxkupsDLZ7VF
3wmx1U7mRWXKeMeluzjv4aBPv1proULMB16mmhc6VKCEV0xvfOVYQeEL7t7SxYTp
nOePJLgDFokH/sZP9sSh9oAzYkvMJOpj9sClRT9l/riNiYbTfHB+MuawxS9BSDV6
2ID8m4yuMfKZW/pGN2ErgHaVrS/RxJyptUCEmpX6xjKv3NGAY/rZZ66Ee6HAllhd
g0lld/N/05Q/AYwlOEkau1HIFclEzaD1RAvOkEXh/iXCsdgMQXVDIOTpSkVq2Dgy
ph6JtZgX5YHNxUeDa342fCMpp9FwwNPz6I89HVtxfjAnljL4l5j7DT1cCOO1KSxL
eVKozXVL2LpCCUTyQ8KPaUDxO4lKjmYdeA5UEAyndGDr4jHibgfmc4vx39/z0Dg+
pE1sDlu+NlkyhtTTBOAryfIW1pUuE84jfzOXPwR7fRoZ1qOj7GyfeA74KdlFMLNn
C2TMlv4GykJWW0hPf39qzeIxb1Y92MkhIg3f6qgAZ4hLuoCxmpRs0QpsHBuEYbmt
c7pYHTr3yaoFTa3a7nRSmWLEpj/k/1VLfdDWS7rzoXYis2waEQo7RFJCrXQieRVE
E7OxsD5iPeXir8uMWuwrnniai9UJuScJevBCvwJ7SmswfXdrTcP7LhycKzlMvuCa
gYbIeHJQ6WZB4jpY1bEv4um/u3xY+zf05v3A1iRXvruYyifcHUOseWVLYFz0Ytl7
2eTWCq+Y0DgPU2qSep4HCOJAD6eF9F+Nb81RecTmeYt28SkcyEUtRUrNiNGixqBi
SykE/FLBpdU9kMUzB3aQgpv3lYRMcrXV87+nVkCvjhnpZAVA3TKtB7uOTkxK+YeB
gZoGF8cMfyZsvfo2q3MWJ+maACJyWmzdEAFe4Tv7JroMTkZ6L/HyAgHZ/Ic9UCJd
uhgYlDrzZL9V//IOQmNw4kXhr4Iy8mV4Zmvc0+4MRu1IBUwc3ntIwjl5mJ6CT76y
gySB8w1recEk0vMK+QthnxooRn3xiTHqG4JXz72j9S1QVKt6Mw9vlanwz7gNubtp
lOcnwqC29utTHYYpx0USrz4qXdw53HpkyaiVl8ijYyJyANbSFqc8jT16Atyzpvnv
sLm4W9aZhKKpZoDsAw5U7zOIz3ztFxF7rOm1eFcwT4C4aV4zDeGUANU2KHWx+1C/
bkWbftfZQDDwfMGGnE9ULtRyxiWSYf9y0fvNp2fEf92/im3R7VwmWQ2hHABaW5MQ
/V7HXMuuJPqgjeXIGNhBAYMB+zd2dt8Ubz972SuqmardVow9ocl9fx8qq+d+4QPU
CVdfRU8aIphfZXZzpKT1ZUelyqxIK6aJmIaNRSt3m6XOdg4/HMrVql2ANFknWPWy
dM/55Yy7FUy+ToRBU+mxKZwM2bB66SZFLIogy5b6onpOCUHHKiyuCXcF9Qas2QT1
NQlFC8Lqr77vA7HGHhAy0pl+7ByX5PK+ztZtEa4xiKBgtovNl2/R0vb4BWYiI8kk
HY1b5SX83Uge1lNghuWFs9l6NdJHKxr5zGFDYhXAKneQSt8n/a3Iz9jgSpE4X+I0
K9BLclZGzUGIiPwn79OpSAWYsIm9TE9iWNp8aUhfK0mqk2olWo7WUufd4Yb8GXZ+
4T45cG57sNPF4HOxjQ5Gknb5n1FXMvy4YLinRoDvLBhc1dXPDXYIl5AJ9avc0fXL
fXlMHT+F2UTThhAmgkLaq2z73Rd8HDwKbVXqWYaUKnGRa6aQOKXDFhH2s3cTq+8Y
azplgt1fdg+RTQLBNx5wR7v6pkvTW9YyqLNhgPwhLStMzSwXg5AgbIcEzE0HibqZ
Tzm/JXuNW6N58nb7gbRHkOJngLOtsz2tNisFWrT1+xQ7i1GhpVEZj0XbI35uXUbk
aH4dTTLcW4lDetyQgmGXshiqIovUBzs+9gC6rPEHCW2CfIzRCb2YZJQyKb4AM6lq
JAmgBDLOKqizeuFaQGSoTkJHfwh5Rk+QJ3i0KBeg1O3lZ9M9hy6ewsWjsnaQROAT
TFnmUwc92Dfyvk3AefXg/JiUz2I/mg/M7g64gGEdiApbboCARA1HOSMJlfhzMJC5
IguJuAPwyINg+C7Cb81rZbpfhW2rVncydRcMa5DW3sYKK/jJtRRLp/9dFRxCSxUr
+a3kcZJEvM8F4MFeNw+lSh9/BABrW20PsnxdIayVZGW+pIqGcKPo4tAZzd554CE4
7UkLgW9FtM1rXTuiFPua+hwwSVAyewRuivOMavIa9KRgHUrAmqMC3FcItne1rixD
CdDKh+1LHeY97N6Iv9h3LsARtAKNSguMJp6MphHi6z/mBy66w1QTAGusevDBLn3U
WPr1kNIkikyhMPN63Vv+n5/KRR9IFZZrkka12Mvi+mZBgcf4dYc54WE+lzB2mACC
mAqIcxICaoUriqSoB96wuJjcpekwsBJidZi77KMzDXxsNP7Gt8ZQJAiOInUhfwXZ
RjQJmE/6ZUllXKixCh99GhkBG6TRZGYyfFuK8XhPjNzmK4czL0doEQ35d9SCLXHK
oLIgtfIOLsu5DiId1VzjenT8KoPdlDWhNvde2vxptfZQ4N5eEdqH5Q5HKtX/zvbl
DLV5uZXBBklyovrE7/wfqGq0ohLQJ9kepMEY27DRwHAFuER1d1QaRm3sNKYBeJQe
NCnu+kRZ9pvRojfzbD3kiPZ+EZ7GOg8dgD6o4JOul/xHjjltXiPvZ3KACAHrSSui
nXUs0RlKvS+AC2PKU+Kn2eNJ8vcOQc3aIIpSgbtLYHXsolKguvoT7x6cWDLa9kn1
mxSgjtRoIXROOwp/JiO4avFCNig3HXeiIApk9ECI/jqt01ovrO9awNdhAz3S4KWv
EpjFhecZZPybGqgXw26yIpZHrIr3zqLNmCIOniy4msuaUXiPF0hlxZy8KhNwDMTm
2gomihhy9rCzO7b1f8WlcLapRLJDDt2GDuI6TaOdvwfU4DFHXPpSyudEt+aMybkJ
YcPs881PRQo688mOMI9lJscdG7t7z9uWrntrkpuDjO3yo7UYX+cBUaRTaPDSyAHk
unCalOGxe08wMyUHkQOb9NG5ktraXNpka+5vyh2ZObT6xsjnCt8pi4qiARQTFp1i
VWh+zm7IXXiUf8HvrAmVEdGL/aZFhoQh1rq0/acgetGELRP0qtz9JogviAdRY0X8
FPegub6yci4+2Q8SAFdVunhzvuSh+XGEt/Xc7EAb1+KJlVH1sOOLu37f8A7lnIND
3HX7BrIIFBVs9FvAyJI3rBb3AKrN1H+DWTwwFBIJllGJ8JnyHaJmITpfJ0LTEjdR
HW5eAkwbePJN3GBNH8LMauD5TGQPKXdNKNeHxBE9p5fd1syalt21UEiIDLjMvxFs
xL+WPKxRInFn7WfZ8bDPGM44RRdW34HBdopsX4P1MslL4JHtF21erDN06Jy7Boi7
2XRgEaS1Z4cWhaUfgm8yws6+Uy0+PlP+2mq4FnDGXhGI9/terSEr9pdO+swSNKyY
J9wZ5uol4jS5P7wx0vk5tCN19ArzK6RPIKF3jRCzC4QBDgKkXuGTUZ2kb4/+pxxj
yc5lJ5GoBNxDpLHnJeMAPMJJ4w7RRzD4i6K/gZhjKkBZr0CjQQMgVWIAc+9SL7s1
Z3ZB6WqkjDwuxyOmr7sjBQ208IzsI09joNiZr23aHD8/YexPD8inmr4JbcYADfZ0
KEmqJ+GxwJr/sWbRKkrghKUTcbxvaKK3jMOSC8wFCH7v9+/gKQ7yMMxMmQzNkBWI
Z9cCk2k8c39o/yoWgljk2lfbKbQQQTkvyy2TnwDXWqDd884p1tv/52HvRBxsX7JX
8GGnNquYA0oJMhgW4lC0uJNkOczq65ALN56lnZ2/dd8aZJxt9QBc2OqMIfptXJ4C
0dvRR3HwdV8l5gpgj2Uw68Qd8FtgWA8Bi8Yb26kSSG/B1vghVYxPScCq5BfZO3Ey
EzF1bb87s8hW8dRtzsxqXf0S1rxOm/V9qvbcxyediCw9oj2dsbEdyImWlOsoi+Kk
rzFiFb/HTwBfHzX7L93aX4/rORKHfSMuYkdAIS3m5RGDH/ostKY9zn7m2YySOKuA
1Pkt+1/qSDTceDB+BIOwv+tuQRbavIU9siurNI8IQueXLyKzY4I3rgnONNzkADfw
hNDwfNTsuT0bXNeaVZSFUeXHanDL1eB+8gNL3gIoeDqfvRzP9YIAEl9hjd5R7Y8i
VnmIqOhWZpMOHyFFV7UhkBPjU/qh/dcwcZZZuzHsUJlD70Vn+t3b3OpCQ2PC6yyg
nyVj9tHZL3glYq0wMQAnbH/0WeoBLr+dzTILhaWmAum67z/3ds1pHe331Gcr062u
teoChuzB+JceDpa2r8IuFA+BEqDUP4KW54v0ULckJe2wQN98Kl//jUPV+TR4jvEa
N6I9AQRwuarvLYtbtr/4zQzU+L/+D1Zp4LT7JJu++4VwAEpdhLC/yuU7Vvhxd3TG
GmTc/b8KZGV/9ZwlGM/5wO4iS587XT0YBZ8TVB8Y0Gsex6X1UjlpfP7oW47F9gNc
bcFOW6TckzCL3Tcq3/IT7nlNiPPNW5zxpDgZiMyqYEb+FKJPVlIw94NUjhYc3xX+
quPaSZdJksnMNVEsOAs+EobO506zAOfz4AjW4JTyqcDmiFIQg24EN7vr1Hg3Ko0J
P8+fJgu7tYILstXb3ta1PO5Kj3dJlljjUpqwkvg6vD0kiqjeJRU+h2dE/Cmq2nra
5qLuOHh7ISU6ItgBjzmTi0qx980mRydvSzHrgx7JnCFFf+jycQpY9TkFGqNySVLG
ubI7InrjRKGp4AmMkxkOQ2+qo3wIGuRhnn4CRy/gUNnnTlJ9jmr25jSiKGLf/bMX
DFiu93CoR5bVASNDJmy1ZQFgbI8/H6w22RjAg4OrQM6SNa4Do5SQa2/u19nEZuJz
XOpwW9STbQTjdnaJ6ucTg2b+d8jw3ymMng7Ql1CcDZ7VSHd9J63yuJNqkO0cJP2M
xeqhevjPJOyieZyY6OeVvrk9woiabdtMjQCF+rV3iYEZLuxRBDSUtpIN7Oqu+/QN
kg03UlfwO8zD16lyFw5gGXWYbtCOayqZ9CHZbrQbj6YXR5ixNBM7AGXrntAlYnC4
IpuWTxMMUmnNDfZEWpkq3wfzvj18I37bR0KocShZ8ar0oasmjqm0AHN4IQ6KDe/M
AeFmMIR1wx5QpuI9IG7q1pvxwjOy7AVQ0E02ptYOT4iIRxl8L9QssYBn6L32RCLl
435FWC3MvO87YtiWO8gFyP+9XBx7nG+VxMfpx4RGzAEr0vFB3BJnFEDftTxPs+iI
duXFz0MMLBkgaofF8jxwTlo1IYrqesuNZ7sm0XkFqrCdXN0MVZF6uvJue0BG2ZCs
x/39iOIdBnbqIQRCk6K1nr5yHzpX/C20GbyjuTOH8yLMYN/FKv9ajJ7RU8nyO7P/
6Vjqbt7fx12ltngH5sM+VoDLLUaX+Z/La9l/7vi2B7GQENWE1TA6iRkc8Qxwbu8o
zeaF/yFqdHdKDzWd4APLDNya04oZnh3qyXBUMVDHMRaup4f1Gm4AS76gE4q3KQXw
IOBGN/GGuNkFYA0jBmzqFgO5bC9T7mw+Y3WFAPunUhCKIScubRELz5sWrDP8XuYY
v/dD2tenNSREsOg1TYl5v1z07PvQAOOqduOQhP1SzYRKsVZtAFqHUVE/KjaDpMhj
HcFNhFllzCw8Qjsvptsx5ltu9qe3ZGcDUbEKNKF/LQH+Z2M7clTFox+7PM1lPJWu
J3Xy+ioR1uk/7ehAh6fmHlgThQvXVgN5htrKTLYT6HwB7df/nwPI+lo+ldoxOdNu
QyynkNaQddeTBy1pr3vm8kuI+SuUTXiGWmalfmkano9PfHQGFSAi4eLjfqS6g7Io
KTzqKTHL5TKcc5CU7JmADpsZlIPSFP3PymaircomnrV0OAd73r2YhxRWR/nV2nD4
kuInBv2tL+6tQPXJY0u/+z/esUzggXtovXZfaaRGJryMB6hfGPzwugpoOYvHcn/2
wiW07lMIwM5nj/sEharvbj9x4vT7AELD+BRjO4BwXTVS1ZmnGJvfTT05JfB/y18S
92Xz4qRs4vRKteMmhlOnVe1ujbkdsrdmZyqSGAfoTpkq7CwDPr4MH0HLgqCqzAiK
Il32AkfKQnfOCnrPrXx54PXz6V2MFr2qfzCHqm9EsfR1dO+S6H1ZvNvpAvCT8qcQ
8AoacV7dFCOFKpxemLvBu+K26bhGcP69bwQDauPOFGDygItG4mAzkVjG21j+0wzf
HK15I0hKg7W/aj2T6LXOmmxqX0zhXRS+XHoSeU3in0t9fqWEcKYczxUxCIdYwBhE
7N+Uj3I3yvZgHiSwxPRJnkbADK8h+/lPGj5iAZpnQqb+FkPNPbMD0hqjbD6ps1id
8wPWcpA/JWUOtuj1dfT8O/9zYJSnaajr5rcSfut1RibJx8a9wsMFCDJPq5u9f4du
8D1n+gSUHMgMUKE7dl5YBRkVkdU+0+KcvNAmR6+Ig0xK+7LoqF+oH/BCuMeXygqr
hTLyzQmxGxut4gH9wyAx1PzLEC+W8Yn7qL6uFj6VDgQmVf7wnx4Tf4sBoOUFTYSZ
cTnNZn1ISxzk2AbAIgd0EL8EFTqtC6LELVOOkuxa94/Y0yCofMI1XYJWG2k+seDh
nW7qdomGpxQat1eCpgvyiGcKoVGcUlQsjlc6mh+paNWWVmTKIPMpuePcwN5EVkKK
9AXdRAAOMCaYEbuv7OqXSJ49AgetLEMsv+c8FT7M7CmvoFqgMO9roQWnqIllyJOA
NuDq8U01Fhi2cKSHAgB/UqGhRq/jgNk42oAsNT36pH2eY3oLiPhv4fe7uwnktPvr
Fd61Y/DxbcO0nwIuBoJrApAklScao3LTdAhX+H23mShM80MeQZZtYs8tTM+fmoix
URk4kyXM5S4GLe/S7/TJ/BrJIIkQcTNukw3qt07md3QwToQnptWMeRyYH5JkvPJt
cR5WJrH2CrHUM61slF3h3NHjMj/QIoeRGhbBnEr3Jz0JnJ5v52NwlMBKSpz7zdF+
hwV53/79NxUn1YigVxJ27tAHhfbwFLs7FfwJqONLqJZRaHcD1BTHznjoeQvpJD0A
nqXAH/Ok/1po0uvJhUqkRGQpkhsr4K9phr6GUzVqzRQNqRvkEwI68q/797OrqKly
oIPeGpIFSmUOo2nSNOpYLHq5L1Ke2IbUkBUbzzgHVIINSRSNo1I7Bdg0KRnQjxaY
Vp9SrfyXA4m1xsOk7gfTnwdndVAL0atPtA23OsvaWpLwukKudGXC/wdZicvgfrQJ
6BrP8mmJNBypDyea9kmLN8sIO/zPJEP0RzVXwJRebJ1pwOoM89ARTV5ukjuhTKNx
6iO4n6vYxWcO6Yx+dhhODNfaPWoUmRftf2+e0sVOnt+/soCfDxHZYZ7lwcYDTfqp
Rr94rkNQocBKA6lLcSmvg3UQKfOQfZzysJOEDgvrri5ZSI6HNSFFP2NEX6gUgWkw
bejuOwuunZ5Av4Asr1aGc5qp8USH4q8GUrms3coVMBIDE9UXIyQou/ZybvqZ0f+E
zSvfg43Kosmerimu+K30ixNhPQqX6NcWEgZ7w/2A5sNGAT8gdv7ofW+eFfT3m9D9
B6uqpuKPGkKPkcXGhxRPh5+IgJv3dj9R7pzu2w/9FJM/1+Y8dEGbQojSEkY2PasE
keqryGXYAXUwbgmCKV29v/dv8QYCcc+BY87Xqs/PTSNtwibgrQQ4mupRoZ1KiQAT
7SrL9TuYJn95oqCg22QHmKJEoLudE4gJYVZWLknuJ8OqXbDDXfQHp7CzbRK9iVKL
DANzXdLm0vo/wE/czCfBfeIEQKjcdkrU0PSlVXVRblt6rP7G1kfm5VNGyRyA1/xp
WgKzmeTlokbn+CW0RWof+7NI4WSB7FFwvqtDPb1SPmPefd1B7FXZgONRK/k1fR5Q
7pvPTiHKP3cratl+ahLTjsNGgkbXLDauzUGTenYJcQ/dbagOtQ2k6NWUGBelT9+c
j0H/aMXHz5RXdDPkdcxDLTnXwpx6TmxKp+Zmq8O2V/CrlhXxEKzsO3I3O9J/qi7H
xiKT3ZYL2JDuHvKVIK63SqITc4hc1oaVyheUYn5fYI8k+xqimkGS0CZYTxxzjmpu
ARNCagNqvtSakUZv+j0Cd4CtzsKvFTBO5oDSaHqBz9b478R+ZK4BRPLAxUFTAb/M
yFrXc7ITf5W4ntbnMIrSH3CIlUAJbYpbIDgtfpiV3EuUGRTgwei+RMCfvad0os+R
8mwDkI8sdYXxYQs9tfTfOMfHH8egmmu1+PyGTV6i2EWict1wHCNrCucFVWDIan6/
chU8RtOGuzjw4vQJwqgDhUVWC9PtVlbHwW6Mb88BsuNqfdSOW3ly3/sJzZnBgT+L
9kXDJVXPBGOd3QH0mjF0afE9ZlfCwArCERWlO8vKfawZUrsbx5rLLHSZ9ctJ+pwo
aCDooo8gI+tiQVR+Ip3eUgKxtC5ZaBHa/ImaR3hbhrdeQM4uynegLJQewY1UzBOT
v6f62bKZS+xXYNIZ4BPR2cOf8KA8L8fnWeA6FnyNBbvG2gP5VDkHRcFq4broXJHS
s8xKWtUPF0qbPDrD/wtB9SmyhbbvPI13r3HlImA0UyIR0HUoKnDwOUPkgGeIkEFc
mt3JDx9fdVZXrfSX5wR4dINHvCPZgsEKlF7HuJH/hEbecbHecsWaoyGne1BiPQnM
/Q/fXGhy7L1az1kE3lpInft61IBSGEdws/OcUzSZtNNR14qwwlusSGqvdXwzJnS7
hGljQ+MT5f+mFQzqGf2VSFy4yhx5ZWGtbYfL5O5SgmFiQbTzLxr562+xUGTBoChd
qIAFOFxIXJjfLn64vdW8Jzfo1UqkdAqVmIL5I5dVRmYCtLHRTSrZmQD4mAjwgBOH
mcBzT8jrjx9QYijZrQh/Hu/zcsVt6eDdEsJsC9ws8olqfAyqTCXHPsTB/bjIKxoA
fHKDR1ji24RmjkAhzs/yKtmxyH8hxwtrRt3Yq8cZo0+SNSTIgv6hPqgvwmNBL6Ry
zmwKUf06zwnk2dE4VPFcCRohXAwV6+1QNkOsF/4NCJV+VP4wFVVl0M10r6oHxcZT
+k6B99dr2pwH+nYkjiO36xq57aBspyc2ggdEDAfna+h+9cxg7nO++A9U61rmiXHe
vvGqzqqXngCU1ycwFLDLnNqHb6HCWZg4Hm01VTEb5xiCcJp1mp2CxuE75TS3QSPQ
i26keGShZoGzZ2I2OO26Jv+S3sv4nlb+7deUrzkaYMYr+8bWYbxKYPHDaPNQkqbs
AtMmqLhzbMIrypn7TUY6CHg75PapUE2CjRo8l0CktJQRStp4C3X5HINc0u8NsgjX
S0LmUyriwp/Yr1EYJt1UlIdzo1umaokkUflRFa3VvBiHCvL8Be2Y/fmUcQR/26fo
NQr03kvkpmlPbTg1LvkpKmyZsBNns9hhOvvVveDazZSCRW7qrRBHH3I6+sKb5oab
CQtvvtvv7Cml8dIwALyomt0SGiEE76sHpWCSGVAy7CiUYs6lfpf2s/Z7wAW2eXjM
yjMv5cWk4zFnWs2FrV1CbSgPOaY9i1/zYbnC6uR2+HnaP+NDdK368pXf9yuOLMQ+
ujw97AP+tY2L1bxOTwLz92jBVnWueaqNHYAZvxfu/9ecTevVfjHiBusgCE68ej71
m1CQimYMuUBvFnRIzweRrn3JsHdc/V3T0wnXBgJ+q2FLo+tryltgYdvXxNNJsxse
f3NTrCwW1jKqBu51jSBhY1vuUiFFSVZpywB0HSJdSPDY0D7hpyD8uZOwLX7oepai
N+o2muytEe4UdR41Dio/vGB6Hz7KzfL5JGfGT4sndZRdsaKBXX3iFTCy664K1dQ4
ipAPzWYFhSUFsj7CDp8nJ2+QG5y6cm4HdKAOs6Feb8sde1ETw14VpcWtpg8tca7D
K2TBlDW4Ko4o3xXYoAKvAygCd63bxGmD8pNO7uZ/uqGlrukj6GrDHyMojY23MgdP
2/SKt3MuwimcTfxDd48u4sjddyQL8v38FW4+fh/FrIC8iKKxJm4ZHvgpRyfVzJyw
zyEs1HjmXeXvZTAKXAYIOa6rF9ODAuGR/vrZL8UD7rUm4E6sVlprHSw9v8O6YlWA
qynyI5UZJ35SVpDBtQlBwBRHL2bmRpbm4/0rGi45/vw4o8sDUV7H3T5bX1CpFdGX
p5X3Q1waNmUXBWCGe1mgAj+93Tsf0zf8yxs37wue4325MQ8i99Vv7k9F402lJVxG
sR0sYEgk56HFyDBw6JkU5uWyokR7JkUi4zuSclXPntf8F4pWm6skGsVYxQ3Ww9gT
IDfYEqzhaoKTODF3PpIrYbbyTg8aLW73LlTb2w9tKU/assnB4mTIvX3Jstx9stnw
QEYDrPsiIIhOMyQbGB0b0gxqrX36KqqFNsb8NuTiFsIb89hgjNqatkj5lW1K/TMh
B87jRRx9fHlz8/io/2e5TRj9wtI6OLkxQFA291xP/UJC+NX2U4MFpBs8if0w5n7t
YzEWYBlqpwVLmWGKOF7t2XlKkkUb3mk46kL4Jsj4ycImr1G80BrRQmEHid7GnRRZ
umPXe9B3NNQ3hOR3EZrTnAHsHOp9wQxLQHwO7LgIzmlwb9YFwyYWWPwj4myitBrQ
bP6BrRu0vtrlxu2nSJWFnVy9F3eetCbId2QSgsJ/PFWQ7bfWm0NJrlBaDl8U1gNN
ciIvMUb9uDpbZujGl0GZMU/wTKuN0DB/Vj7RiS2J18r8PA/2hT/gOEfnyI4PYOMI
tn9XX39voiIm1V57o3h3f3xrwj7mTe3pdxH5NyRh+5Hw3glOSDgroHwQRSwr4jF/
wFfHQ0DIS47Azp9DSU5Zw9xMvHnP8WpcnVJgThvoch/gCoQAkJT+pTK38eGU8Nrl
FHjJ0kcWgC7Pvagdkixmu8IW2uQs92+uRWA70V5D3hxlKYolgLvTYgBTtJAPCN82
Cl/TWBAcpMlBA6TacxO4tQL+lIc59dwuySwSrDl66XTN+0QorJ9D4yfhJt+2zsUl
hqGUzPn+Lt4N1BiIrVop0u9yCM9OfUNVVbYsa4fphTCUipnA/sFmt+0qaetZCaPD
yjxWf8WngGFwiIF7rmYysebC66qFBjxyAJ6MJyxSk+Z9UrxJhEYSZCpjYUf6HtYc
1n3UH24+AkqOxYVcm/mKfhzXZ8DKjViW/VToLlUcv01F0xDMGYXO9Ap8ta9rZwnC
55p9ShxKJ2HfZwWDSDQhAkRn1BNTDZr6v3rhw410tCEgnt/FmsAw3sHNvNv/3lgq
TG3KXw8EDFFKJx6F8/qWrm2cJzM3l/xEWlbVfmwD0YInTSIXSKQ8tF89karLPYcO
EiZ1GlMM974dSD0Hh04lbjktlh37AjseElkbSBqgruJLjWpleHr0rM2YZNV5GWO3
P0AyWYwAi/W+37BD1JI2ewZiHziZcuiflJnWD2zdZVWAmIn9iHq7BeCmi9OX4zhK
rARD2S5ENVw6oaOl4ZoYgU+D8lorsh5So2JXFLTJoAnsCWAinOO1aECzzP4bcZPM
VMgObE5wlgUvK9NRXhHeEHbcrSidQgzf5u9rJZjLc2c0xrZwhzQL5V/oFz7A59ZX
og3G1J0OQ/iZtij9eM7+XzSL/x5UrRLRj0AwUO/peMYNpeDTPWo/Rt8hE2MaoROO
uhlbQnan1WE5Y1yJRGfZye3++QxXSh5CelWKjkN3XGsfvYt5WVRGHEXOCTrl+Ypx
79/3suLMnWT00JdVPbOIFys1i3lNLxlHyWhK+OITO5dXmgXuhp/3P5Z5QatJNa4j
rXPP5K0+AIlDzYnvGn6fJK2NX4cUjRfIaAY7tmFgfkcEwdlmBbBmYb9myWJyOk9I
B2keJY8ecEodSBsF3IwxSPXRPvsfs50cfMH6i2d1EakPxw6U4kix4BDK7CODSqMV
Jtt34XqiJpTAkG9jT/zjI8KdmOV93i/kqbbDOZA4qBwuBCVWaPTnA5tmXj4GzqtB
dMryvYyfsY1RGuguAqGtkDtMWMA7Mf2DowiB3HDQ/19XuhbFtNMlTXOZ1ooH7gJX
qyv0EK7zCZ8UMOojviUaPDyaYrwwBm6c9eF8cRyH2XiC7+6I73VpLtWpbiazE1t2
Rw/Nzt7xzlblE2cytGmTLvoXIOP2gydoMRuwikqTRoCBA0rPDbSoitYBF1Ojgm6X
lNbjoCaDSHCi9PLNwaIwBT+CjbCMj05SS/1UA3H3yTown5nARGNm0uVGDgZJ6Dem
0xcppKG5jq6vqLSoSP2vEnklAYcN4BX+u4UHyTMRlYhi3p54X9hXbfMsYoK30eJf
YwJ9OtFQ/4MfEJLCj0Zo4XUCNh9OukPSBgOmCyJBX384gOqgG3rZfVuIfl9wZD8m
+R65Qc60LrQQH9bOWdqfzdtv0Yw905L8sso9KRtzUj33XHlAYzgwOD3iBRZPY4l2
kJA8XsyYzSzLQSe06CwS1Qkwiasa5QjZlQdu0/kb9RlSOa4g/0NfTkLhXVQcXoll
m9YCMCbtyGoeBI2PitdefLvDlo7qzzWkMX3VNf8eo9G9Voxw3u0ZDlg2HBjqUo/j
Nd83FWbX/hk3DjSeAekWj+490SsUV6eXpd9evF3h5WAwMw8M7u0LCO347MyemQ6x
yHOsqmq5mVMXCDio/LjYsVSnN2hexy3gBxSznCHPoYM1ckXmQ+9Xk1TL2UbSwUAP
2ggiZk5MJ3WV1703f233U5Luhjtz4+ZtioofkA/U2n7Nd+Ksq9R6YrDjX7vF/3MV
XkwhqJi2tEX50dhi4cajQY5exN++fpMCkwdi+M/TxN7iJGGhgGBk8zJFI6hTXHVo
37mHzAHZnaNcsb6HQpbn4qzB99hCXhPwT5hzPOvjZWevAstkymjeqPuS7eZqwzB1
X6tXiZ8qaYiD6Re+M+BoXXbQlyLlbav04f3pXU2ubIrv+2kzD6ebnAsDVr97mSwg
o3bM0Uk22i2FGkELuEfl4sYxaOIl6OSeyjpXurwQVGZ3zb1VZYoNa5HzQR5BtSoj
igC1tQ+M1Zu3RYeZQe+ezTw7MX52mt21OQTi/sKo7timjkHLHRrXGee0wN0b6y5A
t1U9Ym7qRQ1pU7bMCGuX+cNo5mo5feqW+epg6eq3ydZB2V6sb+zV/nspgtZSU9ro
n5SvYTo6a/4feFWEVafFEdvHWGoRXg6xgLyr/nPFtnqh7umg7iLdSyERgE4/YIcQ
vo6UdCZiKGrBCL5PyJQIevoDTJ4C32e2Kvbv1YdaGPq3eqs0zUMlJsyFp/Nz4zkl
G04ocCDkdUP3Red2GszwGPADF7lUAylFF0s7tS/uL5xnhRmnvEoecevAVdbYatdh
vU8V6kgFIZNspIzHA2ZLMqK0DY6OfwR06bk43zaSQcsO/+5h4622Vfhu7rg+SDRK
ingj8uFrtPLzp/Gamjn84edVdGHDzUjbXY4NEv30cE974C2siw9T73+bsekt3EQ6
bdOrwTDiC+NbrjIW6zLkrVPh41FomH9l56hbRICCtFUomo+Je/hR+S+ZBEOaD1th
GB7hZapOhiO7xhmoQGlpKrbQ2fxAo0hTfwvTwkVgyWq9dPxYBjAMn3LiwpUzVgJr
RyySqSoiQJygsgKyM9P09u69fMAz774hTJULBmwvi9WoOx07YjUSMn9z6jAev0up
0/ONBqBUTHiHacS8xouo4k5TwkmoDvMSyKHGx9BS2RG+j5otmTxY81k6METe3s8G
jih20Tv/OYyYUxB6Z8vMhDX94EiQ6XoPUIEDDBRp/37hJaaNURRzr/7fTPZwbyMa
hyg/rAWje0xxiT/HbREEVgepKQvYqA3ntsBxR2Q98RXA6WWtcW8kePZqDGJCTBbl
68vrVPCUF/8q+p/soI+Mt+nJ80MwoIdSkZhDCKpT4gflCgOe9ACOVRWloy6E8UmL
LhsbAoXAJxFnfa5+ujgwJo7/M0i8GTmHQX1oV+ij5CAqNdVSWq1Hjul3srBhi9iO
ytUYZdCR3gB8BxjvtWB2PQ5P4Bo3mibE9mQroF8xxBli5msbTHjKUIDtNN33gzL+
f7Ijwhh9Uxhx0mlvmy2Fo+yncQoKp3ZGJW+7hL6qAwIZBrRrejntpVf5Y6dhsSh1
oSaRQvJuSdJ1hYXuXIp2KSFjd1WpO8psXtTlaNbdLuZhOjqP5Eg6YeWbGZGtLjqR
8na4417Kmsc1CunwvjICna0q1MM819ndPtRbmXwc/ihmgw2h5ogqTvtvmG8ZkNvH
YcO5ponneBI1ItkiL4dp9X+y70F2OeHv1HXNj9QhOhoSpwzRo0Q0aXwjfTqfm8h3
k1CW6dfh85G6a7hX3L1ulytHIMaBNj9D9vPepLEP4KlUtIlzbUKzRaMMVrwh8tQO
n0FblyvxnnCCjoch80jBi1KsAnZnjcamgWpqQ/zXu7zyd9/fcGziO7xw8QPixKYe
fhCGYm4NksLYPpvE0/MOfevavjvVZpkqyLCU9e+eJ28L3jR0XEa/NXcCJtVItumV
hjq0P5lK/XPmM5UCrxoaZIvu3aeQ86efV6j9MM7xxNm5buM08HGL1C8lBh5ukCZv
xLGSq9YStXN3CRUm11DR6jQbCaDvkNFOD2DvplaMg7Tw9p1ZmAmbhX2LfMspWV2a
L0xOVc3F03x3l6sYrHSpHEvNyHKJbdnsZ3TQX//2RxPwXR0l7h+wJQX9ofM1kAVm
l9oU99ZL1Z84snHfpzJOEkw6QgjoXPV9R2DpMIWIDykxfrih0kXhXeaZ3CaMqGCk
1pxGa7myt/3pghAaaIvAV3dRtiAIs3WLzyKXezg2bKKvc1PISWIfLnFKy92PPh0L
mkkdqYdMFK5s2afXsCxUMbTUr5TGNfzMOHl3J4NuS0KMwEh5lRJapIrCU5H/akvB
xM4GbUNXpvMQyiIKB0VFZLaekZfsR5H+T7Zuyk6EvMIy2Sa50ux4GuDn0hTaCO+R
Ly29x8fBBMvlpFukYG9QeJPyJEvjVaPkoU2FvtYPSiCVs/ocNETf8afngh5bcwX0
ABPguCtLRynsoWbz5/XsVnZ6XZc7Y3/3wKYXhO5QA9QHT8POZQe+0LfCGuxaXuA/
HR2E0nSRw5SNZ0wLHyI0b8jNeo5X/qsXgJBHy598pQfRNoMtXx70yBpoM7Os0LYi
s86hTKiSuKFqStT47uy9Hu+41snqm07QCjQWfMn2um/xK+L2xBHKV7d3HS07I6vZ
E3DEdXakTWwgVmpjM8Iuvk3D6fjNcdPFvIjLcA+v4mxJiPDXwiDiGtDgr390cy9b
Nf8Sh1pRgEyO0X02eL23rO2UMBjOWgeJGjUbuxLyShIwEI+R22xrI335nuw029dP
x8UDVrt6e1MYXT8rXGfgBjuPQPYyWLYKT9FYMVXYMDAWVzj84aEf/CujlHOsZaaN
/Mt+tpzh0Aot+JcdO0Tqjh7r83ZIMLti3yvgCol0G4DPvwWF25jVomW50KmU3TWu
11umOTtnY8DlmsyYTgjzn/lhmeuht6n+L/P6pq5Qb5VywL1H1LmBQFYpqh6NztQC
HVXwcrErzI0yJMu5upbAl9HkF3riOq+CD+1d0VNMyOKXbzV9f/BdaX3vvV0cgDP8
q3JlWW/G77mk3GE5tNqS2CokWgvE7p74opAEDPHxoolAP1yGzCArNXTjsQyL0sXq
CXbM/pF/AjqJlDbk6s+ZQHHjk/4tg0/0aGp9APAI4ss60Wmstyz65PC1p4ZXzg6l
CmUuoQYWBlEcWi0qNM/IqN3KcYDJmVS0+L/T9gaD8OS4PifHWvkRsNH2gowjQubS
0LOiJf5zAffZYuC60q3kn2wwrkZJWGfjU8NJmnNzNKk3xyILsdRsNVrMdRRhfZ1R
xmlfAbVdgEsiI8fa8gZ8AJ8vL+lvUqvSkOAwog33bfL7ueuSOlcSh45GBRp7F9+7
gAI8MRzrnHTBVPcML7WDhr4sHfvmv75tb+ptHdKkDqpJw4bsXwdR8ivfaOQaFGIg
Ri5tSa/sfXygMmvhjVqwwJmctZrfjbHeFkgRz2HHSrdtncdO35MYF64eO2ZkhTYE
XeW0MvbPwCQxEr73NOrBnDy3iupErz4A9IkiKwMWOqc1vkXkxvqQ39UUvhEl3HHk
Lk1wAKeLP0Xq5aWc29QD+Pc3tzxAokdAJff0g8W8SkBHcGc6jrH5NIxWS+boK6sL
eFOkIyqVe3oOzrmw9OSCDLLQezLXMdSc7J6KO3twoPNgqOwh6Qyhq08Q5AiHrlI+
wvKs5AyuFMpGE2lUTnM4Lqok0ASTsxlLP0QWTusiuRT8qpj3STMlSiitFxAL+eVv
T3luezy6fv6vZwJ5zG+UA0eggvlvthcuRgZ8ZubCs6iZbUXgtKvQnoMYNNtsqciw
xhe5mGTElAt9Rm0ibhfsHknk6dfR4pFKmTBWxGnhTzblXqkO8S3wkE2ZO6Fx3xdq
+0P92hIAdag4rpyF5J4Lnfw5qi5RF7BsgM22bdL69tg0CtR1OSlY671loPRz8o/I
xYWaIkQ9Mt28CcuPLMO8+LwM4zQZZeWTCRxnDBKBzCleN+qcNIXIa8U2aStj4DYA
gvJM2Okb6JuRUlBnolK2z3BrO/5MX5tKKUdX1oqAxH/iq6nwB+Xal03y/GkaWmTL
0zLCpANqHGwjWwl0fb/TSmGMigLg8w7N852lLnln9XMg7WoZc8mtuIqdSA2MHRgc
11enhCaYJ/ujNHU+pyXSEZoHC+DJqnzuAw9e1Z8dQgcMNbv7qd8/fZ9AgIKYmkQV
YOI+PBSHqziPniA0CF2ta9MzARXlTDTVgfz7bltLzuGXkhM2EMdRd57D/+WRFdrW
JxQsFPNOkTXuO2vq6dmARjHbeSK3UcPZacbcO/JG53suElSkXzRzwXu1Fb42WD/Y
m01vdGJiRII4dHozc/hDa6HuMwO/gTWtaGN7fgq9OGKdRLIcceMEgLYD4KNQPqbd
02YsF7CZWdFGX9IoAw986X29l9bRACwFwEKqTNImir3PmUcTA12L54Qnk1a2drcu
/DK9MHxZ3qX/o3VJy8p9ikO39jdmlM5dqIL5o4ZQLwCmqY7OsoZmbOvlaImMxMcW
9NS0kiCQnhxdL1OVtzCLfpopoOTlMxQ6n6rF7BojnzhvAsEL5/UDOIZz9Milqe/B
joCJwF9Tf0pD5pLLQtUkHUh1Pd6GVOmE+9MWntsg88VqAN2wzcR56YnQ2KB+17EL
U87qgf19hj63B0TzGSOwyHM8j8yyvJRukTHZEYhlWDSROmMVpikaJ1BmFdV7t+WJ
59gMF9ad9oo5/4n0qZG7ZwaeNfk0y68iF8eTjy15KUtOsKaFg+/aqw3znSWGr4lp
zoO9NeW20BK1EVrzCnWaPfL7WIqIH0SdhRlHJfUE48mAyq1MFVyN+HjuUl5bS1Xo
C2ay78JVJFbpcAEKdlBiyvTTMgsrM3/XNpjH13bYY0BrCh4yrDCz7llPB1BW0xMf
CyXhmO6YNHIAQoOehF7+gLmeD4vp8So/guZi8Yw9ox35Qmw1Z0UAB7ur5L0xXffd
mjFi5Q85yxOE1GWVVSE1sa2en3FwWD/gKHuC98EcXnZo5VbtTuzJ6OpQmR0XdNQY
xvieqrPcut7dnX7zgxSEqZn/egfvoA2fZ0qsF6eevq2TdW3ZDZzjpYqVu2U++6rP
ZobslenHpEHeVW/eKRFk6Np8v/Muj9X8QjeWLOxAHTuhBeBTIrY71IiXoiCmImDc
luA+BjO9pkho5C1wM6PQQN2LcdtZaTt3xZZ3nBGpKI+xXcJ9KYonvAHyrrEN6D8/
Qn4ND64Wio/PusDdIUXyI6xpKhg7iGG5SCh4EcJfqlVqx4otte2GaRAihcckufXt
UrxQok1fEVIldoQc2zRDuv/1lJF/xTZxWZbMVr8a3dk35zuQ+BzSgGVC3cQVbU6P
hGHgDKz66CWbihDQt81FeHd2B3Pq4GWZPas4Kl96QdZg4Yqsij0fOig0a3kEERGW
tpIsNG3kdIBnwE80M2n0Qy1gBW3ef4mWZPdi2yDpZ53b++KN+pUiCoVOF+oPArQR
Xvo6WTH2TLmBPnx9b3rHeSTMavWbhM4aDM03uJrSg5fvb4lD2znOIBBHXVIVXMKB
hzj39P06+3PS8Cdpv/EIBv+LXX6ARlYAYcK1V3CkiOny2+6wduBVBkkY2XggfbD6
AkF1y05LczWYeHaGNtutDeURarUGTLq4I4PHNg5Qx7uFbfmbNPzqqWtHn1M6Lwos
DUeRfHPI9gCnJ6YrmS789A9hYGo2h/tKBfhzKTZxYoPcFC+DwoK/PHzG40fkYPEw
j4exYENAaeAkojayoY8dN65nQ0eaG2fmJhHxaoEL8Tq7+l1Zvhs3WMqmQ9KbTGUS
RuyquT/vw9AXQ+8wVHfyXe95tpBGKHRuv6pJ1/w06w5J7BVZhoRQ7phMOgXksp7v
4NEzLDWj/poa0hNRUeE1ONsxUcudRx8xyBGw7Gk65Cx5Th6qN4rPiQ2FZ4u5jgSr
lBprXpzsD5XWasUiVpAtRtk0rTC3q3o1OT+6m9uHwtAwlQGnulcu3mNqs/ZS6xJR
0KojiFFBvzu15mP0+qB4ZC6C1Wrc+x16ME/pHlk8xl0vN7Wj512lPkjX1EGRvP5H
KLqqrbEKtainhjxutqUyB7Buk52wwmTeSygogCN0xvBD6BVVCo+dde5hvpPVsgz7
M/yMR1i/zGzYh2dM460Y+gScI56pUgwxVZFrbFYicX7Wjs3et2t8ePocUyyVf3kL
o1LpER9eJKUz2lAxJU+DdhaKvn3a2NCtMKlbyASauFdxEWt3PeNqdxPQrjnv4JgF
giEGEbPh0HQz/iAsCidMF639fOQIaRF59gMq97ernCTtTmmV6e0t383cEUL5EGSg
PPFzxgQRJ2Qk0QL5AOTN42EiBroRMkw9ryKiSRMRrp5GliWU+65oSFaWobkPIcy+
u2uj0LN3TEXc1/3ECKAL8GUHovgDOTBdPushRwfnkbEtOCr+uhLQlW38zOfIC1Wi
My9xUv5gqdPPg+5iHXhKegVa3NAmhxzIv2FXD5eTRr4RdeWjO9onHuY+MElKn4S3
vCL2m6xU9BhkAijC3xH6NVoA5jVMdOEXgogxl1caUvssSAKPn0XUzBG+eYb0hPuj
ShYYwvuh4gpmOeqbKbpkvf16mRONxdhUONqm6xUk67qwYJ6ANS7zXaj1mSJ2pQxA
VGpeKJGrMXIHzns80hVH2CL3p4S0+4p+VjO63W73/MoaGxAqVn+SZJUerOAkYQh1
F1xvgQTvq4CGyLDNcXeVxVCGwhaEDSmaOWDGXlMjPCJZc0KvYg1qKOa+qeXZA58v
zvmkOiKeo6AKt2V8mEhk5lNhgzQAg+DsPHsAQAGlbw1BkkkA2nr22i5o8iDROT6u
YLx13pup55zNHUGvlwkrp2sikJB5BHGuPuqPRcp2IugP0ahPm9zkkzEcnKeqPgEy
IXZQOjahYBGoDKJA9TgoZyj8AMyOjgud8NKUAg/+6W50V3mQ8lmRcUqgC9vQBK62
9Q69PEarvvhSUf0TyWU8LgRu/Ih1TnFWtlc8kfifTa8522t2uKzikeWXlczaQrzH
94dECH3sN+6O0NKFaw1H6trDiFoI9j3tbFNxm/x9PLDoTWFPhyo+KtwCdTpj+Puq
wLeZET6oe3ATqm1HQzKZPvyhsCL3s8JQ+2Bej42WAmFg1riBDT92UzxZG7YPHJ4+
xQrrSu3n/JoTqaDX9kWpniJhcnOIOrs5xcGboFm5smDijrGyxzHcXzRwUzaXAFdf
H/Md0nm/pzy/W2SeyPcsziRqof+gNGa12/3pIZC+KUx1GDHNDgRQwPaokO28+5hq
vUXnMa6gzOe7qqa9jyEJh40ls9hK9Jfc+V5RukXZVN5LNwSFt0354jEZYgUmZZ1R
R6OGXo5SlrzXNLIttuW5uUvIomtjeLyscSXqlmoPb5d4nHDwTFJ1T78MevtqB2YL
2Jl/nQbHOmmuHFk8gcYxqYlx9a0O2nX0b79j2xI3aRjAMbtlz4RBWOor7YDv8APp
xZZGBCa+CcdqajrBU4zRPYSsK+xUshfkTcyaYv+aGmcKg31FSZaDIVg5UA3cyPrA
T1nny5bk11Lo5Vs59WXQmJ/OHtGktCGJbpfXHChf3wYXA1SzWmiio+T8mwZFhZMq
ExHAJRskuszjEfXCls1iv1xtLmEQy8qVSDVCtUwO3IosKzofqP++hoDpPfCTXn5b
ZxSBNuDDVgJnWkBRQxHAWM5ZUqs9B22HHVWbOviaU5v6LUxjtGPZeboL5YGDU51G
Fs5L88thz23FQX2tCn392EJnKZtmeJ60BENskkUkYemcA8Q7+3fcJG6SGuBd2pM3
MplQ2j6BgwDbwIh3bl4xTBeDUZ7mnszl/sMkQECbgKF32NROdur2lPSCbtz/mUnT
98/b5Efkkhsvrg36tev7vc7Ovv8CLz8Mu+sqD1rpZcr5G2dgXQJrct9rLh7OTTaK
flB7kV4mpbSZlADNLQ5/1qKeTkgPLbrzM3q4Nu21V92+NaeSICzBM8ccdAKso6Dj
BMT/lyDyCLP6BWA7T7WkaX9Pc0iwJCxd/gTf8v06TLbuHYFrMrLDfjo7BUbrz233
ApTjUcUS9l6Y+xeSXf09f3N/yJnZPtXOXv+kiEH3ETHyxxtP0tf1quTAZmWh8p2u
c6f2srRy/7qnzPBSiCnFM5gXlY1y5aUFTsTusf1cbuJChXOzjXgELl05Z7tS0rJU
Em3+V2XDJSgAx4nMRiswcWATzFSv2KJofrgWMbPufPxnW+mmNkrOau9SxnVFt1vF
lzR/5m3Nhq0PFIBFYPQ2VwGelWIJVgStysx/pRaLpHfZC+2hW+xevWQ7y9P7anSR
Bms4wWr8Wf5MveHa7D2FT0SDExXKN5b5sHSo1mIWrHTLs4tPWHvKQcOOfqyG1SGn
MiYDSMYZ0i3ZXmK6qb1km2O4maIJb/IY0tZuj/Hi8ApBIofFJRYQWZMjOyvfGzne
/QHHolTdNUqvFOGd3G2wTuZv1tztZAYlfGGU418Huttp64g+v7URdzgrIM4s9TwW
r5pzIctbWXCY1U4aJegkwZ6HOoCjDsc4Fry4VUQOHEwF2VSzZwjmQRLpue2NFDmY
Qc8RLsI34dag8WpQebk5xLr8EHTtP9l6doqbkWIl6fV5UaC913J9o5AJDEhH8lHe
u0EkbOTzUoWJdZrHt7R5/CcuE2ss/nMFdKpcuG3B9WRcpIk/1RENVHCcG6l6PejS
VwNxWO9rauXyQrTmqYNWnOInjhBwjI7KTSAcUy2wcQ6Gw7ZeT2Mn6Nj5T2TNhf4Y
8Wib8qo2fRCn+eIee6ZuA5xRMGmCPxx9si2O44i7OSAcxA4ksXlP9GyAud1qlksx
Opkovc1MjPGXDaoTHMXnBepRZU2dmlfrbt2GQ2yUOpGiSvVL5p4wqQlfqV3NAliS
ARlRMfjdRFDWqu1mDd/cm34K8uxBbVXY4Xo4YzPv/8l/kk672uAY+a8lARDqK/HF
1rDcRxVRd7R6CMzsRDh7GnpLShhRKChCYDrZM71bHWLNr5r/Cn4L4hsNSsjGQFpz
SqwMjQ+WncDd0mt+/PkGcm7MeSYTJDmAin8R9x2L4OUj1NCTYki1XM2YUt+7wdoL
WvyPq8/fw3AaREHJr/U5Mm7PfYflScQGlXhctq8hdQz+pZa2Etji8mMX861C9ElX
Tjk7kchMf59kaehSe0Ag8x+s3jqxHR5DAs7uN/hkGZGF3EOBrp3Nw5PL7YCGpbAo
zt9Pr9Gx+fgXQnZDb3px54EAM/327AUH0lj/ObHj3Jr3EjpJP2O1N+yo5U6MfE+i
dBVXYPOMva4qW+JP8i/sNGPdlCAIfOlNV97EAY4mk5Qpfl8zMrXTgJp9tONeDGlK
4uwXB6kzZBWPUmddwZuyYPW1a0pK7P1m8SttztSgN9amXFVFIlliBg+B8WzAr5Mv
B9DK1+mjm8z0H2Fk+VesE/7hBKjq9eEN8/NyLA6vjR3SM9YF6R93AYCRjqfx5HLJ
2BOYK+rClPU71F3Co6HLgQDyz9Hd6xxNn5Sc61+h4d1EhLl8UIUdmfswNW4/YkzZ
MJmkf5G7aXMPYEQGzRofVjyEmqKXyBHHAnRxPOYQUenRS83EGbpk8+gc7nuD7Bwi
lx2IqOjsnJyXGPwXYOl/duBXZpVlux8Dza0VO26t/X/LcAlBVOfG3Qfw79ThWUSz
Ea7ncmJUTdKEONUzRlwWHBgY7lXOx2BUyJazgHQbQn/8SUeQkpjhOBm2EBPHnXgP
vQuKp+6GuswM+UizFp/OIEE7hqsxVqVuhbIbhx8YxRSmNO7KMgNx50HU2SSg4iMs
0Df/asXoiFCb1wmrZxfZYqO1+tLChncbbCjDfU2/kBnwMhQ9Dd4a234AqX7Owto5
skgffCKqkoRCXDP6GQ4tPrM4eLP+n4F0kdsOCPMYQq82PSau+tQULSWBZjENRDV+
LKRuBLrZHTZeQbZb+H/Pl7nLrhTcestZ/vQNGoOtVMMKII4/YZIgus15aakMrh+i
fvyCcjLLzjMRiwPkeydG+TJq7lFe0+PT0xc3yFq8mSCMrzuUYPaXxuVtQiuPea5r
85kpsCfnwnZbT5wyjFxY/pwD5P0/JC4WrgVza0GMoTilKbnk8vBEOxIR+s8+/LqT
TG0kDM048Lqqju/jpLY7RWZqv0o14eoMr3cUjvcSOEskHspyNw2DzJvlyXuq3XGN
FYQnzGLDKO9Ys/F/58j8nI4gUJ1SCiSvFquDbw2UksKgwiV6v1WMO7VccHgwaoew
8XynkN0QRWo3tLlLoGynFHzsUy3bcp6cl+dCNsDrE4cAqk75liKQRVQhXb4FrtKs
tjllafkqd4sHh4UNuZV0AIovkulqeGWZ7s4RJPH93bjBhBlZzso/wvMOK0b5bGc5
oP1Xp3rVw7rODryPLRuBrFGeYK/194XYv5HGH00JCQJcroab7nEYonLmSdd5oezh
i3/Axzocw607TZ+yxof2w2wdiGodASWz4TBJOqKctNO+ZCFn2XmwUn0oZLe2s73B
+VtUffTdLunOYSiPM03GUip2TuJDxHj7vVY+Sxv0czsFeAbrDRsvGIbMAl2oLNDD
asI+LvHKhaDnEE60/oP+E0uzzDkOiBSo4tEOy7VWRSXmvUV+JdlQ5AZI+fPcFRe/
LFo8YWtGSXbm5V/jFaUs7rz3ZS/TKSt+torU+mhX0e9ZZK5vzd/ph8276KqfgbkH
DSGq4UiXu+7rQW+q2Qd+nCCfirA2BWQ+/qOZnOSwvP50EmWC8ezfFDiQ9I1u6wBM
95xFGSGC/pf+zAu0LY5A+jVhWyixfOugmrgNaGmM7L+MbdvaHQqlVyMWdbV1EyiD
A3Hqsary7AXPXxg23t7FgFtjZ2qr7eLcnraj9LkmNPBhcP6IVXrj6ESr/d1XspjV
bwlT8Ze5+ZAf7AdwVBqDS1HbP3o4TpfxPMP/5Li2qcG49uiqZUt5UIvXSVpt3Xai
BMx3E8fM9t7t/rKnpY1uvSJfF1tI9sX0kr2jgGc9hLwZpKmjqiAEjhhxR2vKVZ1j
9TmQ8L2QHzJaWnsqLdLrxgj6ceuZ3iGmo9gVf2SPiFms6Zl5kJmv9cRw5tRvwEeq
LEcuhJs2OdLTHW9YWf8TR37HDN1A/auQI5o+TtAH7OqUbiOLRdIhNJTUgX6sbsiH
bgcqh1H829NhoIO2MFl2N1MgcpA85SeZuv5BWfv9SAc/fOhmGzp7efRRnupEcTaX
KgeWhb63NAuEWbBght7wv9jQqKThIQiokT5ZrX/8+5cQds4bfJ11UttEBJoMK6e6
IccyCui9EMk7Ds9pHFS669Dgyu3bxPRAhAIqYn1N54vXKE+iBcMYpfYi6oxPIwBa
ESRnYce0EYW1aWPa/1ucfIAwCiaUwFigpeDXnEeTz4g0SvH5mwET6ITO9Kc9jpTH
53yfsMq6FOlST1Mh6CpwXQ==
`protect END_PROTECTED
