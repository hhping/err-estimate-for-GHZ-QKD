`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dT4sVJKs349hZ31fLIZzMAmr+5m9LUcIXbjWrFC7gbk00Yqfjr2scJyAK0tBNsyx
vlYUFfd6cmwcKUKodfFh78iPiyXkWUo0E1Z74OBEdCD83ub+XQguIPUTB38XHMP4
nmb5jFxCrQOSrnHPzk0+felN1VABqWgY2Z8RGjMuIATbcNs6ekWLYRecTh+IgeGQ
bjvnwDE/o89c5iwSmGVXJN8SnRJ1f6c9RRtYqyMWhkX0kpjd0zmLcgz4/+4biE+T
mmuvAjJjzDJOdKLdOSKLUIuSxU0mp1VC4JKk33EIBg+dymmH7i6obOSdHLbStL2t
TId9Vk1dL6h/znJwfl0JHav54Jt4Ziw3iX/0mXTt2vki47nTDs+/benDHt9HPBKb
jXKGzfQC/YKlhloLqFdmDE7HQLhRX7pwtyIwaLX6j9IDd1buWk4lCul+hYqMpF7M
cUFzaMQljh6cvWWrKVkatfSgyRfkmytbV5vqenuWRccCNCXcX26VYlkaolrofLJY
IcqWXX6hCfqpFs20SCidffE/F6lVjD0pUsk8SyT5xZrB7AxvT/lYNRq6dWMTPe5b
3OwABd8InK1i8ooJNHp3YkF5ypUN7UylieI4dx1PEWCRYvsDXB0GIUd1rHZfDjHz
u1gi3f4xxRkKuVtwTOByZIyF9EH+rCYAL0BaUJE3n5OR2fg/h+naSS6g0Pk/OsKF
GXmy0Q78qXj7zKuESQI1BjLYPDnhXMkDnmeZB7eWy2senWkG/WK8L9Wuazp/KpK/
rBPJnY9GReoqbmnsLedtIfOsXxfvUIA/qG7F1yd4W8I4sl7nMGi85NZHw3i8uuBC
vSHM/Znty9AmZAi1q8BUYwrS/MFWp41rgWAEKXYxtKgLvecgtn9KHA/7JwESc8/D
8iUMdpjDYXdyEjTgVmtCMRnGt4M2pRM7KrOaWDgwRHH9IAdTvGtLfe/48CUo1cPv
`protect END_PROTECTED
