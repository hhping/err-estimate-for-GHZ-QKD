`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJmhAS5rqYKwbLpgQ6zostfezaz+WpV51PZCnRsnX6SPZ+EQTcQysiFq6y2R5h2Y
J9nU5HvJsh3OLCoZC84J5t/mTXx7uZCCiSAI2wP2jpEqZCzF3yLfdCDhXL0rG5w6
t/A9WLG3z4DGYQPYDEYC4/v+lWCmUCSnVuhCS1i8DLTSsixU8AGRw1+yOskTtPkZ
SqkKSYD4iTmnHE/5OPWkGOcXBa6+vXjfH5u7qebFvUOHaZSR0jnkiASBKRU+4bmr
arLWgaxm+yN3D6q/J0+IVPuiysZSbahY2eHpbdsOfEMHjJkZLuJLH7eRLc6ewRPk
b5sZuge9Q4stH9Ho3pbER+6pdrh79iEOmbmM5+3rySuZkGCrn7mxASXeTtaXeqUw
tuXxcL+0NOxJtbgJrYccnRVazxU0zh0aqfixQ4MIGg2saPf/CUlqmQ2cx5Jlcw+X
H+KwWeX8O9PrYyx5fqGGoAjHvxPZQI8irdi/VTN06MkrdGAVTEBEP0GaMsLKg7Gq
tMp13XsrSg1/Bfz0DUrTARiLmXXAz1kPd6hJmnKeytcmM52yPo0rhJ4csaY1ceNy
uWBPk6FaWBQHp6OsBxs/PCQPgYasv4ootcPAG9j0W9av/O5easLyEYTU/ncjJ1gW
fXQYZ4/nhV9fQGfXBWyJEyO6TxYyfIbgGM14RvMKioHk6c9YeVZhNQQdhFPiiOp0
I+ky01pOmMJp//LWEud2HDUgpSgjl9V72nPttlngspsDkNp/u1Zmt2UqJTmc8O6e
41VojG/a1HPyBq3kX5uaGjPPu+subrp9B1VihNP7vgM2K28GvKPkQar0hdcHc+VW
B9fkc62GWEMLpCmBsMKltyVcL+HpzlQjQDdT6Onpxnoc3OHYDIoK+6eU3UND+Rlj
HmwX/bNukAiwdcIDfRPkbUmDIJym+Xoz3IDBIbqdD0bMB68XLU47uOHPE+iqntIu
yVAQQ7o5WElkpmbP67XXkB4VqBtWPT6gjaXJP67JLHaRWHKY8jMFy3+CgC9CJZTb
kSZcbuNhVIYReP1+rmqFMmWrgEJ5nWZcwemOWnhMb0fFbYUK161KKuYeSFFgEkqE
zxTY7Mu6dCuCdpLqkkz2/HV9jPG+WsvBTZ9UEkEw9vddbMOkCYuqSrVRLwHLqcBs
dchc+79lhPDBHLBF1RRwZTtWI5DzVhQdiQjmVf6YjDKxOtCIkojjUEQRTfokLrqL
z1mBBVVwrtvSA9rTNWjKHezuMd85xGrEqgs9ClaAFD10yKMNMDKVUI4C1wsyG+JK
k/kK+w0/L4uWf5UtRnLIH13NiyyMR4r9QuQqlOAbfjGcW5Q+5YmGkH8AOwyOrApa
BLJQrFY3+fELuFSjQODI6QpLGqrsgOq2BOwOO4UIrTc7BbpBBEXoPIiuzPpa/39t
u8zGgY2JPwcvUU7yTlVV9uMkTZ4oDd753tfKYIJAwFNwI6Oo40GeWgnGA9DC7eyb
aw8RjEjT4C+K/Vzj4a6mVYDdPNNj2vE0BpLePcBuIaeccVvCZTbRxH6jORRmSwe3
Ikomi4XmtMP/Dy7MmSzIzhP7WR6ZE/9zoXftWxp7NlbFcZa1qHrB+xjauS7BY/9S
dhcjCYqUy0klObjzcgxael8scSq67CrJA+AgxU417WOUE2O9gVZiSk/YqeqUXKeW
AQc6y0RCmXJcrg2hGZak0JbSU/mYDhRFBmHE+p+YNtbLMyAxPvEqNrf0CrEJKoFC
XP5AJT4WuuYVFdj6iuOQWH0gz50Hb34T7cHaVRWw4wASSgbMQiOF2jQETR/R2D6w
9LfJmJkbQn2FR8+V3dQdOcBzdOrbVKpU3PrLr+wKT/zR5wnByEUnM/zWcisEoKbQ
ZPlofqY1SUJt0zxsTPTHVtKRelwE8qw9polrrJIhdZU1CpN9Ntxi2D4wodQVQQ3H
OlqO4hFjObwOHQ5BaEbcTQ==
`protect END_PROTECTED
