`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPq0yGYV+9ooWL2MP+1WI0iQdjQ6lJwY9cGE5ceBACzQNvOCzheFThgqVQry4/V5
vn+vO9OzTvxy37gfEzhKSeyGruA5Rjasm19TnUMYslSrQnrV2BbmZojQrvY2xavu
wbQD8wneMnhIM0EpqRXAIXfJ+LjuUJSBJbvUSRs+JEsPmFjQYiK1jtUXJcXMpMHi
lHQvGy2Z1Y0Cq0TmJVpnh7pXE/QdWnTmxztKdWpyucsjRhX0rlIMuDirUNWYj6kG
STCxDIy91kbjp57TCbTx3bWYiIjBPFTVgdt7VRWbGBe4FN+g0MoJJaeqsbQvE96W
XQiTzS7R9AfxMlCaXtcAPQH04/Uja12W6eh6u4P4OCi03RwVgKlFxfnW7tYK+/P4
5Gnz0hkTm/ic+Xf6niA/u2bniNO+SXWAp1ONghewuEeXV/QKmiDUyuAfkxjvxnvV
H4GsHUQLfb0o+SedbVvN+hjoVNg+GeH0zFeoZfuBRuv8Trzmg4E95eJSJUv3NiML
flFKjhnRJOnYK+vEQQvxIJuRt/QGs5ZCa/3ZOrI4cBOVZ7AmfHuc1vLyQqxfX4lH
Fbdt1jDH8pCCbXwOufaMbXlNjeJoTr3fxLR45LJ6CWD35gPua34EpYxJ00H+Y7jp
E3FzCfN+i+NCcGbEkAZNSoX8ZfFX5C2Umiiz8C/pv/+ZBSfUEqH6EuoLhL/90sL4
z8dKaJpZrx9SiyyakLbNXkck/yqWmF5Bw3ulurMNEiQl4SP1PIgR93dlNKAI9QaY
`protect END_PROTECTED
