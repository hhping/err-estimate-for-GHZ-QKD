`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sF6W8WpexHjhypqksma54/H0KqMC9W5E50kE9inoFoOhUKa5QsFDbM8qwzgksf01
xF7jDi8IRPSHAkGib7xKjjeeZP7dEcAcDWPz1f/JE61LuNTH1j3lBNysRkokXOKA
pV9y+lpQM0sqlshhGcxrQoBNDRfWqIw3PPCSPH+S08YRCOeoUs39FlBewReanQaU
jm3Zs/7KJIndn2F8wwZG5a5u0X7kSW166fnxnIBHpOSZQW/IoRU9js9CHrFb+mqD
KrSMJL49QA1H1Sd4AAv05tZGzZ+MQTQ2AdXv0uQtS2UzVs6oPHsYYDXPq+NrbgqX
V0u+eTcMO9Zpz+ZrFifqROM4ezvNZuNCoJqP7Ak8srp/KTY+E2FJwsgWsQ1Ts3ux
oWWBZdI2n7k0NLVI5+4DKtlgfwVC6TgTMDaTovJYVjeO6HgjHseFAJY8rt0ENqQh
/WXC3ZiC5DdqC+0TSL/1wllaOCS3YCC/w+/PIKOYA+d9goI2DVPhlWllx7D2CdEh
+pstgYKXJ1Q0NN9S+L6oDVH/lO1HGG1aY0b4koJhF7i3GUCM0+ADCdcmRUTiKuF5
qh6kDvoWPf3DVnYdDHprVg==
`protect END_PROTECTED
