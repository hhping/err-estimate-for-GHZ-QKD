`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5Xllqn5O+mzUXjGaJfn0Bf9yoQczFPcYn/TdLvecJsFK8Zy9z7dBGQjfwbaJTVy
cah+zOjRixhVdz/pIjH9MXKVGj+6ReEl/RynTSRZRsQwT1gaq9HSLQiFGTeDr5uD
9Z6ZAadLuIDQiUwyNbZDut+4XGz7E/c+7cRU0MtRJe0YIG1cO3xNdhg0Es7Ry/Oz
JtCqAsCS0KObSIByPhAIYGWmyrOJxAQG/8mj3O7aCGrhJuYxN8XImG3BF+/WjgHb
op0JXWA7NVPFUqiJg2oGj0hUA3folR2aQ+7pIMr+/yIp+hQNrJweq6zZ2tAG8fzi
wlLPElle574MTzFy6MuDzBvl8UrUdgJ1edNE9m2XPnPBFjS5ljyfZ6Th85DqlEYm
h8NEoXIJp3dWQ0/inZGqdP1JSRXHDs/7V/8jYDTlK4PYqyR0++yGwVNl0w4pgs5R
tYE7i5BZhsW179CVRbeoMOB/vOUTCvS3x/+kBhvEGuKqoiWJeZAe3sTfoUEuMdBb
TTsAPWxX34MKdZC9uvdc9A3qrEVPxbWU8i4hS4BwEMTfkQ6a7gBbQt10O1XYc2P9
7xh5oufZVw7FZGhVQsHUwjS6mWwOkygEw9KHUROnFswdtpcyWvrPWbX4guxCb0fr
RwQACLh9p54obtV13RKHE3Gw/QOnDDq+KmVIgv9KCulVGbKuupHD34cAt/VTcU9k
2nRWgSjkBbVedEbKPCw1qgIIjGpj3YxrFXenPE1w+PWmcjXV9sxFRHdqKKge9B4Z
H63Ax5VVw9TrKiqbgAlR7FytjAMOC4LLgL4GbFgmXbFPWWlsC2NCowGOaBJKl7Y9
g1Glhufz1tgE0+X8KHoTP/MKeIN+D6DP3DEVx0jX8eZSm2p9vuO5+TBORqAFrUMj
gc4hzlh9jZaebTWd3kETNg==
`protect END_PROTECTED
