`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAuoXxiyo/Eb5xE8K5yssJZSIVaxZfrRG04V8SMjs3eT8twW1HHfIPfc3kcbp1nU
ffqtjQ7E9yuolII/9yQC1MOwm8yeKwNv3YszSeZpg8a3ikMPShqYx0jLXo/4tzJP
kdeW0gFpE/JjIneSLp+lB3BD+yXvYyrvMoIMMzPyS4YWcUtzdGbPNhLsM7cBHWYL
YrkPW7wN3qSD6gb67ZniHV9b84TD6zXqj4W5JdgrBaMssOD9sWGINOSrGADvm8RZ
SLEcRBD1UKy1Jym1bnd+vycBBapfq7uDwR3bHzQp7CB2l96Ejn8zrkIeWBcZJ501
QMQFSB5p/b2CO2XuFCNa8oEcxGOmqdSsWWfBslvpEf97Q8UxbhS21uu7kl8jAkXx
wIryUlv6ZAHd4wFwvRSh8mRKwgvltO9gUvsKrzGhUMYnWzQJIn7/uAo0u1KNmElN
5MPiLfnwySVcELY+6GqUt5Kx6oVmCJqRwUZlSQCQ1amF0M11REYLUdF2YJ9XKffu
`protect END_PROTECTED
