`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NssWUIuB2hKOnJ4O+CMAbVGprsflthNwz4puXnV7/s0SD7oGz4B54uuGBVf0jVW0
Urhgq4n8zSaO/pqTT5CBC/houtTT/zg16MFezX593d+nh8J1Gd9mIjrWhaIqZp/8
6YDRs9e5SyB7jM5RnplGSyJLqH/LK66uamIMMYqdfDnOgHH24O/jKN2G1o3SLyoX
r/s+5p3CY23P0GbY3X/ScakLAi8h8ekboTF8+T0XxtiuwnZMtkqJM4TtEfC/E17c
wElENs+qzXUTLU8tMXzCBSKsZqzNv/W4tmlOlAoXiHv2BsUFp2F8xETsNaXA2rz1
SACvK4dZuPPbsiGTHO8sCiVgetyN/Tq6waIfpPQtmZAkVviMd8XwoNWTEk/UHZ/N
jH7ylK38X96tdrdBxNn1gjAVp7kA4JeWAXRK0yr8acHv/50fhyhqrWOcCqjQRCCn
WGzytg5xehV79oz/v05hcWnJsBV8Nd1sHoQESazIIPkGnRnNAaDAZW8nt30nXL7w
w0GDZxsGXoDbGyVP8hJaAN0zqugxTEI5N73o8MjJcAkrR9dd9opZwUPbiaPznguU
Bbh+vn3plvHTZRVSBdVfj75yzdLd1M32zzYb3lSVJZE3eoijN6v3kDRi400z6U5e
6ZVt3jkwnvi/cgl1W0d3J//Y98xR9HfqhN4EOeN2vn9Llz9EKEZihKk9HX33QLSS
nhNE2nSr/bhkgDaR1umJryZfCTzhUA+q/lMdD7eoO+sxFi6KuTgl1ys7svjAqoMs
cA7Qgx1YogyOWRzQrnZ2ILx/ci+It+Sl4Gc+36qejes07YTZnGVuhwDBJP4PwVt0
w40/xHMbvwZvfNS4WGB+wiskAO3SbMyys+74Pux3nLHu7p3cmbybyYq4sft2vz9g
Fq59CIzTprMK6WJFSnrXsTubeRIa0ZcrgJSOmCYCom5irAVporE/AgsIWqujdP9E
Qn/K/RDgDl18mcbNioQB4Nv0cZicf7Gvx0S74i+liD8cWv+nmxByBDIsGMnC0dxX
5iU/GJyz6ZDxOIYlcsfLHwVY6AkFC5YnSlNmxp9xDhR+EamZsUJVrPjFUNUsHo2G
EwsPIfyoBKxrRyohtfcxycBuFo+lZjPuCpB+aqclDvHqcOX7dV6DBg98NjQuOxpe
W23goTVtX7ihJmSL6GbeEsPjQPfD3QYiXoW92qEpxil9rx/qQ7bn4+MLqLq5NS4P
mR2igjGKDPfHlYOmosAJXw==
`protect END_PROTECTED
