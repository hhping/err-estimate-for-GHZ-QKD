`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNpMAU7Yx0O5FlVP5UkL1mdwF0PmoG9IOR32l6WFjLniddaS1C4lBPvuxV74fMMI
d6yRbiy/0ZnxplWshSvAZmes0w9mZVYrS++a2tvrPI8pHvpRcir3+VmneA80aodW
nVfp5vrh6Eve9ay/EhqzvsS7gOidkI7+BhKvETND9sHGvYKh6hhzJ1j2KQbmP/vY
5283c7uQdgRhM8u+wsnRNAKbbF+cTNlid5lhiBzOcJBEUk/Zg0hPx1NzNxBpXM5S
VDypLq8jEm4drb2Yn9Z7Pg/i7Hk4EP74u7VQe/T1j6z5nfu0ck8GBAR4uM2xPzBz
3Zw4np+Hl+AuO8KrmbsIQgv7Xkp5/7/h5tFBuuX8r2xVqZ3cQMUr90q7ksn4e++e
KiMU5+z/U7B7eiI/XxFCLU5FnOeqWT9xuIK8jmKjuXYozIlqTnYDMXKyXE431jh6
y259dkr+bvLdCdGyhXZtJ1dVwlBdPxlKBtEWTnhol46IhdENWf7gZk405C0rUnRz
wK+869G1UgIqZ2Ck3nWWpDoz8EQpUDzzvEAgsFEHEuriL3QpmYZyX2c5Uu34+Y6B
MJ9+XeYG/LSlLcGwoYfR43DykOYKaZW84u70eksHJDk+2wf+xws+rBf46z+5keo4
1NL1WrtRuMSHRNlEIeBFQMORX1eeTh0h5lpb7QDdBkG/M8O/8drUWaOmE3A7BmBq
X3+eF8NknvcvpMXb9x1NMfMpyxH3j7ouc3A1wSV4PgRkJEYgDdmOBReLIewIZIKy
y9CXIkaSKHc7777DqK8OQfbvp69kUby6yKwbrPHEwdmJPk+F2hkzXjxXmsUQkm7N
9ZB6a0bmFixKfKhH79KUKv71r7Cu2gNiXIJGFc6ZXJb8gnX+QNn8v+cRnhy5upUh
GHOLSc8j2m6bJE9oLdEY7KNWuMkDcK2ulWTbwD98TzhUnVUDY5srPv4n+nIMbS78
6ZmqpbLSqSaVbW9am4/hpyg62smTPu3mWd1Q5dbIsvycrW8xZx3r3f0XKUe5iKtH
I/qOGusdX3lTPRrKLub9a7rZ4iptawi1aWz5T92nR06ik8uKV4CbDgCJEbp/pSZc
XV84UE7fgpJwRjaz3VA2VLS3lqN+sMpFWr1NsSz++TNXna9/3yTlHPhL9ftXPmG6
usVxoEzu72iijakifiArakmGR4sxgB1rrdiAnyIJUUHjCwUe2zGMautOlysezOVx
MX3y/bFRDS4kLa2UbNYtC+J+dtu1RB1S+ha35Q2i1L2MYWhMCgd+pwW4Ci8szCJ7
ByoSPmocZ1vLS1nGT8ycsqEAyLclRYQRYc3Q7P91qNe2mN63YfBkUNg/qbcOxemy
QKQSHqQD5nG7yMYDWXwl+7yb/bx2jZNm/F5tV0S9BD9LMy/J4EXy2ekqniBy0xzy
vKibPKz6FOUQgbfiZaBGv7NlMEttLxq79eBLikkGAi20ScitmDcuFJmzEPUVwRIW
aFIsApifv6oZxolqbNLLn6UhXXgQl49m629w+/Nx7a3hDysFabtzR8JpseJp825m
68D4j+jYzAInq0Qs2QVWdWbytyDUjD4lma4wc4mCWIqZmWGwnNEfEL/CseIJFwhl
FMIMMH28xxBXmWDjZKrH1JxPwBi3G+LtRQFGYO7mYACVRu2L/9y9O4bb0GhbeSu8
NF/FkSHyha268/3ZwgCBwcO2jWAQH+A5DxJe0REoYAQXDFEZ6A7E8/OfW+Bc5Fom
oHLhaHpykkHcsd4JoFPJJefsQju4Ls+bCEkgU6mtNNERafwBnt0QlerP4OaI21GG
1hDiLvBYUu/enDvLiLTr39gYGtEMNV909dn2kaQX95aW7TqLhLW/J0+zov9vcRcc
jY/ZjDWsDXcPhMRWsEGK8VC9r9UcDsfPKSbt8eDf8zw3oOc9hv9I+0HRdcGXkCfx
sNQLIJ4vRCw/1TaQYaibAKhhwoabx1C3bKCjrAlSTGe+Emxlntxn8NAySPY32KBW
Aq/AKHYvNoKnSUpBx14COkcM1wrpKXiL/3DU2akrRTc4TBpbaBaNYjpNVMlP3dfy
wns2y7fSNyEgtZcPfhRVb3c8EQGtUIw5+ES4y01NLJkjgh1SZaldmPhkyDa2czKj
2DCetQPr0ifKXksiVueyKQJmkjoU4Ci/4nFBdUYFwzKzkP04o4VZrHLyS7ODYzpH
5ii2qyYyXohGzWIPi6VObmtSiBAt+yWJhJhAYfLoN0XT752TtKD+597PVIYQhzmF
AEVU1nzMZlL610ijcdux8QYdtNCvHlnpo9GccqQPYpUBQWLAnDlru5rFomPIu/z4
HnhSo4YyXlVItphaWhyY6kgP2yzqBxokjjEc4smglrnwbW7PSRwj9/RTM8Nq8mQt
5jUDsQOKdAqomvp/9osRTKjOyD05cYd9sS5zlVgignCaaqYNEWvJOAdHylgtxpwL
mert9yQRnlCPmEAMnjmvjsE1Z8OfJi0i4TQNAD9a/CNUach3/xED38iTNW2U0SH5
SAllRI6GBXnxxALVg2FyxUIMVKY/lGk2kfUtqcNUfXSnzsZn+lFDQ8w7GarhpF2c
AFd2nbuwAjFF+G2CTqRcVj7PReX056ECJ+2Tr8lXIl9VrIG9hsxyqASBv1oYCVsH
djifb1YNOUMdt3Lvv+3IDdvpc9+Mf8ppNs4dBE0Y5n2LoptWa/sVgidpt/rGOPGH
Vqwz7AG3Sicm0LGpYuUY/HFipFJ5BT2tzZAWUIiTAxJGw82h2i5LXoVZWfFw6yE+
xRkBz7aEBj8Bza0Y1DZrtwGOzguKV00I3+mOkWj6qUhNxWainDeHNrfN4wszA67L
DNBiYqj63kEUkQkAWUvWDI5PbsCJ46j9sVjEH9R9pebgNJ+kRt+MHRV33OMUkHOb
vMaqaLFrsQv/bdSBTwttJm7qAV/JB9DwiOVRfpSJfDbwJrkWVhKVCtQVtax5I+yF
O+GbU2+m9X8q67izSZxSfRfaI/Pw0zk7/vuqcFU6U7eoPsFQ0q9sgq6Gv6ysF5R8
DRsSODFlKGXAYA6esr833qR53V4wPOIyZ26KlKs+d8c98UlbGfey36pUlYu9oR9Q
LkV+TnxHRFOSftZerHJmpoJDY5/1RQ8j7fkqMN450iGzHTdGPWoV5rRlC+z80Exv
SeYMj1r4UFChMtNgrJ5IuC9V5nOxlFHwg3MB8KC+vxeth5IXMUiWXz3jAj+lUCdT
SNxexFTShkQycCD/2DrGYL5y0ykmRFc9evskhu/oWuWY5yMUXQKZSD9vQvtLYc1M
G4lOikog/6uD8+Hjo1AJk9eN5SH8hYOOP9oCCrjeB3yPPrPBQFWa5EAyTMu/XkGM
/YmNe7jkh0NQ7sVIhT9D0DJ5nx0emaXsRK0lCWmz8lHAR0oRMS6NgbQ5vPdcDrgU
yZz9EeZvX1T817zu49AcVE/ayiLoAuZV7/+adZtaeln50WBsJyppCgwlllCVD5vp
p0QBHh/ws4M4DyKN29Ir05gLTCqWRlntOhuN4dM21+lP6uIpiJCWKzsnXtWTMz03
x5h1Wk88WdHv7knMmQHz9vVB0YxrOQ64gfEjcAeZxEw2v98YRp+0P/QVpMN4FARE
3eyiSVHsC0yKcN6pMoaMkgBZE0RcaKW4mwQBLnERDlxlR1TvvTJfOUT/yIqmy3h2
CLuixd5YXFrBxMDxLLiUGv1gkwcVVr7ZTUlwQIGulxBUZytPRn9lAKbrnSMRdE4w
+BR20DW9kg2Wo8SxuAlG6zXqf5RllRggKQ25x3VEIobOOGXeOOmaCSizQ1SZAW7h
Uw5mSvOpOWANsGDLELHWDSCHFlqgonPgM2Z/CKGdnwDjFKZah3npoNrSz1BTvyO7
BVn9m+UsaW+8MgJpyj7KjDyj3HZvXchFtKJIJ9cgQT0PXUYKzxuqw4eS+8mJlVyL
LHkVZqGrdw1CH8FcWAzSoToQ58HzICYnq8gMXvJBamiweyyAqRgl4vLI1MEqKlfs
f/OMBBDHs/q3lySLGl5dbiiVQ2fuQckiYZvkkniv9qFwekfqbeHnRaYsQRyHlMA3
mmTiVi8QUDF6CUGQ4pGX7dX+CIvDwcHu+NaqiFo/t5TUO0UDaswdHWa6EVWXHh6x
jffSKHbJb3xt/NDvZAjFDCQoceUOk5XX7SNCLhl4EG/mdCSZ482+cUyHR1eGv/wJ
ZzrcOR5uP7IjHE4SteL8coEmcoWI0vLMfTUaZBQn/oNh6zOcHwQElZ3HwU9D6z7H
PaZNJDjcbXSK52vHPNe+L/IJkO+ce+1K1UOjp1dsLoT+ihmBXRZ6eWSlUyr7HYKd
hRd3hWnpYe27wRupqpf+xpZxvGpFAxpf/TPB93Xxb2YTFwTiZmtjzIa2PyzK8ZvU
/buRMgPkwwsWGkBkoH3FKuvr5lGMMTvuZlBkncoBI1npTLxkUcc12GrfsGbVLTvf
58Ynpyd43cd2YsL6J+3NUZbn1XyrGq+/CgKK/hBtf45BQl/WHdFmENnUPaMjGb0+
HKkCkwOKV/uY1zThrwzplRRkuWXJWTEfIk7knBHRCra3GXjpj/b+YMT2tpB85EfO
+ryBHKXTu8RsRvnU/7PeFaJtsEVrUXWxQYhXuoLuj8vFW39asUNlL/VsOVWlYvMm
7ddS3S5O0hwA5RkGDuViyEjV3AgWGZnYiQ/FVRn00OdJjOwvUxTgOB+V9CYRcdYv
vROiHTRM7Zb8bReZjsikZq7yiejjSq2VXr0y2JFwOF2l0i/+UHrtxEkoLyhufJ6P
thKR9U/Agmy6sbZfrw+r7DwkkCyVKlNy0A9jvLYcHOAW/Kh3780h1nzs3Y9iUIC+
SzkGdGksA/b4/P9lj01MMNjkYluU6QlSqCk1VNwHTENLzG4zX7g7mz92D7M/pCAO
QLIzXrPG+eSl7+A7okGkSUWSs159cN9MxavM43STa3uMjSH0LEeRNuWg2sm6Mjhl
3ZRPhz6tv6UnMLHOrLUukmbiD05RxTvbSC51hASNScGmfsD15tKQPQULi7TTczYb
R9C3hVgRwXuwfkyuPHhSP65DffgTQ4hs+3Mz8rpd3lFuHjM8sPRfuSXeBUEipZKt
cBu3qcV9i7MsWy02pSaToQavB5ADoJLgiFtOp3o/tC4PE4qcIU02yHXqaGw9ILfM
ygfzZi9BztHBvMSZ2sFfQ6b1HvKeSacXWGS8JRtji4C7N++Qw9c/X+T+THzIaoGa
cACFzMQWAL2Kt6matnjyuJZqsANxK8Uv+tvMEQASozDJUv3MZ1nEAD90C1va0avK
4flDN0aNbqOZdQNfWLDHF1Un2VhJSwMbEXziSElNQIODaB/TVxfIEpWfMeNIoqBA
Rp3ZWp1jGFOeulZVgGDvrYv3RNA/8gjq6diwypuL2sGSiYr5FigZnqtHaLcEi4FT
hSZMvhR7nF5gN+0yxB1C5x763+0OAy4N+016KhiP1R0ARKU0EUSvDz9Zg0YCTyDz
N0zH6xYts8qH3KGr95AEZtOZkvizpCpuwUHtDtJT0ZCz+bJLo1gn3zdjWaxchCZF
I2oWfnfKbY/1MlqyUrbkg8vz0GgdyUludO/g1ezim2VmLsO9DIF/D2JHeWEYNrVU
xVJn8zdU8exBY2/64RwMvjtdla0mr6kv4W/0C3XmPMkzfIx/wqqt2j2wxiMns+eV
Jx8xKFO3kS0/loamFVH+t8ARTXCnqvwN2hwuk6M0B8yrNFpHzcHNPFo5d4LYhSh2
pmuaTM+PPN4xqYWrYt0uWXi2w7pIjUTrZwZOs+RV2CEoR/hW6CR+kke1Jg9lKnmw
LFDfoMICqrkfWhh60xdc25sVYTkwFCzkrQnmEVuwSa5CVpx4K4051DmWWB2+J69L
S94W8WDsZZGf8Ov7pVrCbZ2S+slXpNooQHMSgwMEbaHc+ddW1mug7F1uloYp+SEV
1RdqE3tdiNq5ZQONjJ8uVIgz6AgbsksUzCrZgmXmP0DiUxdndaDbbenHq9Wu+PMd
pBS1hKxzFyncojpr14JbMAlIIk1Zr49v/48c5g3EYn9Fi/MRlb+4+jgkDeJ2vUSu
F9Iipgzo8ynx65MVj1MuRoF2NC1wLcJdbumpFJ+p0VeJpLgOd+B9t3BOYwWVu14o
vmX3+8hIb4aYF4nSNwtCT7dVlcz6KVT1G5icDuGtGffN7y2MArwLHndfvkGE9ANb
rx/JxavK5SAuMN1OAL2VijBAbTlphD82O9UnMyO03/iQO6WVxZxKzOaoXr0MVf6q
W3BP6KjB5xxKpNhBZIVVJiYlXzdGSyP9nanrNxqW8XoeqQhMAzrp9mURJOAOCCks
CiZuhNxi7e3WemU8ZecCyjlQLQiPakzZG5jGqCWY6qYusV/BK0PmbAktv3AEtKBX
hYZGusAuMOa4MNShQ4nS9ra67hdWY8DbC9EYOv/RwdbkVMy9Nq32e/yaIn9Xi9GJ
D0xbbEFiWS3DpjyI6Y+oK8ZNPEIv1tfF9twEIa/bROEEY6JSAIR8TcKmR4wcuuhq
Oz3EFgDE49TwWsG7c/1BLfWq4ejsoUHUDnVxih4O0d1X+QiaeNTECsJzV795wga/
4lwooQY2AM02c06rFeFgLyX6LSqq29ue3fFZdo/9y4xzpfI8ZLxb3Tl7InB+FQBK
qMcROI0WnYDPff6Zlf28GbBOevPIgjIR25sijMaQBINO9E+VppDJP1XDe7eO/943
JTxl93wTeKXhc7ayxuBgUPLKCUl1u5ot+5JfBE/196bipw7zIBwhL465ZK0cBISy
jv0JAazWC/u0YZjDwhI0thhP/5m56Aqx27N08+FnI+XT8zpuqF81Dvd9+T4UrHMn
L8NjOD4RPnKvBelLO46IJqhIqhTcSOyxG0TFPdhHiMOVWT31uQYK45Y6//rYmwQS
B67R6vj9crQRcj2Mp2X3IVbi3Cz/zBRQSLamBanDn/bcoEcCRRm6bxxcoHS0Vx8k
c65kU9TqE5vLRB1A0JWTusrTaP/bcqVEHSGwXlSrrNVSun9YYNa6lNwWLL/vTGRD
PmjqVK+UNGmvrHOeWatXr6cbRc+FpZEGkmq2F2lRuMYYRR+BepGYtU68bkLMhAhG
G/uotAOO3F+O1VfxNPXf4G8GqADlOgpBQrPByntkDV9MV3EsdPUlqu/+OnB2KawR
yxY2mZoY5bgbh/Y5lBA0HRVivg7V4k1MsMs8umYxRVgm4uB15lsA4iW6IuEkeCMb
TZkpSatBDgIW9K6pS44fsN+fv/nr3LEhBSNnTUzJ0FWVSASuLwG4w5BMIPXqaXFW
cUosSbVKtdueOkdHVuUPi22qhT7+w3XJjUr+HDyKLCLE0dFarovTHgDrPEftp6VS
Q+O/gyDZxZt0NDyYvL1Y2Mjk250GgRgS3nKRpy60Fpx6XrnA1DHUYaJe9qXDxYA1
opF2X0EULH3KtNBHoJ2qzs5/UU8B1yXhRQx0L01KhlUX3CojZJzQ6+pumKm0EJbY
mSOU/NNUiM/jWOjajakZinPBrrosXMH4SkeCm7QJAlSpl9Tb3GuGhNjZfBS62o4R
8jXC2KONpTcdp0KJt47yvXS/+9UUAwxtqfCLaEl6mVLn3nP3nFC3Jzff7fxi5dWi
0o3io2S7SIqgzeX0YV/lsJvroPvY4I6GZiVzHINITTVXGFeTGXX5ogtiyqpZAy/v
esyJqDqaBO1ciovNRYERcYWhUjzehyKFKVDMqKcAnpV5u0cU1mtVXFl+Hdp9o1Ja
a1vIRncDxUYzTkoiLGSV3r0DJhrNa2gsV3g2VZON0d5cSpFq0UtM9jQJLknzBWzz
RAgEkNr7JzI6YOb9N3vOlkDD5MOqsdMbblvWvdDStva3fbNaQ6bKsDK3hu0eqmA3
9jMlsY2KcTCugcQ0fGf43DsAYSU2+Yi9AvVw+ktljTeVcg3qusYWlb99ktcyZ/e8
12aeGm21bj2ZBnKB6VVr4BARz77R3oCv2oJrOOGq9IBucrTxHSK3aP0QelliH0V8
V47CfozycMTD5SqXPWjFB1pWEsPm+G3RnzYZX7lcfrpRMPWASXzBY3WisolNuzAz
9C/h84hdR+OPh3vfP73DQuKZPyochBwOoUIWjK3r6lgkV59beJRKDuEQ1OQTGBbW
n9pWe+d8bV798Us16hweGDfA7ec78qvZXFVKHBIA8fdYRDcVgXbCzcvZIaeVEeX6
+c2+d6kI5Cnm+PyjlByGWGeyBzPM4D9/ZY3Ec8pla09ftNykxcoWll0poMQz3BNw
Ks83RBAZh5r1olgv9MDppUftxmDkIZ7Su2+g6aBu+95aYWC+g/p3M1ejRECui/0o
ubMeHeyrhi0uf07WLpb3AWnHT5gbhRl0HaSdTpci4qopFKyTQ7/LoLa68QC0pSTf
qt7iVc0aDAByqzHubHBxWoBf50O8kAgk7iEUvL6IAR9rDOzIDNDArCEjn3R1Tpoz
R9j+YJqgD3l45+9gDRi1FQ1ROaVQooauQiNOcif7WOzj9wbx4fMmnjhsLadbLZ1k
QxZ4FfOvwOQJnQqmMpwd1FPcUiZgiRdR2NFUjmPdPGh8F4J3MRQSvEcYNox5nqec
HBayCRwY9Kvyk+jpAsSqdJ2og8UsfLIrTMM9IcqWBupSGflRue3o1DVVDFXlPY6a
2XeyKvnbssdn+ww6b6vBHhJrc2wqGdL82mytb+2L4ap0v1qRtDIjyvSGuu6A9S5p
HAGY9PluW9Fgnq0KxnecStP1rMA0XGhoBdWi7ZGreL+2pd9cXuwRWXlwJOphxN4f
4W+1hyISM0DblfN7FMBuXdVA1AJSC8crdyJe/NUg/v0ro1SR4kFs0K9tyX/y9+oZ
8w2E4NCv2wn2aDzBrznMJwXoduiP6unpLhigS50o1Dyq0bh0hPjFqLdYhdJjOUuL
KTKjlMyL5cGiiVna7CX7bvU2UUQCxbRsw58k9peHoPIHZuveBYWbljzjefLL4kKk
KH9ZmxkdYADeMhUF47AxyGEUSUHb7yiGn8BoijyrS96WC4x1gQ4TaMeJgeVHCXin
PSj2fZjE0PvdTdv2Rwd62ETZtDi5QHbJpJ2tV0fwZVTs08itu6M3rvbQ5WsKTver
DL9DO0vr307IhzZ7MJui/spqVOq6KU1yomnfU8VFFiShMmXvL2KY9a0S3K0fXUmW
Sl3cC0MlEi7LFIJ+054jP7YofpHqdNX8jh7J1mRzeN8ZPdn5ALO7OaYe8OhYbolh
BMp5caWVxCn6MKnlAWdzAhasyXMvmy6MKmvRIAFtdGPTi2lmrt/sGoY5/GQn7XEp
Di1ON+C2ngYS/bF58ASBf0kRiRoOhoT3UY4ht2DS/aTP3D2qybi4qQ+1Cnc1fDGc
vY6Dzj2iEuQd/UdH3D4BrPZucsys8B4eirnClafb65R0ffa7WahwcURjzfCaFi8P
AZQ+s5eSIefOrBJsWSe9y8NMua7qFLu7e3vUmfRFH+grVT1ABVUYEexJtL3YDHu8
h5kDx1nD9rryZrEbqKkJ6vof59ihL5rOKKpTU6l9aHLjetYPIfelcsdvYxYdFBnW
wUjISG3B1nvBOQA9w9Xtit23MIjmWyXDaMiTccShfsaTi+XvYg9tj5k6qrw0pPsL
qaGLtANxuqTj0NSMeBkDpRrZtWCIlvzJuR4KDi0asTg/sF9i5OTnW8K73BISN3A8
4JlZj2AfQKIe+ErCP30iuC0R+/57K4uyZKLty/iXGnEhRXzW0DDMGOlZyGEYvPwN
t5cSEfJfMVvrTaGIy1emiL4i97k2ovlhisiovUbgX/l2xhMEpy6zLeLe1ce35pP5
PC1NPmyLNMjg7S32L37T5RsRu/RHvMTcA8rgvrA/LDuRWBpf6NEGzpVZahFJ9upB
qcZG1M7Hk9bR2OeRNF1mzaj8QeFmCXIsL7L1t/QmPwFY/l0NZ9jZ301cX0VrnFyx
6qXBrF3TuHemux7e9EvDp1EP/qI9IEagCq0hU0auNj4q2Qhzb+SR05LdNhx76aKb
rsJe48Juo/bNuJStZ/+EpQ5s7KjxG+s8Ljbvd2W3ULK23YGjrxWZZgXrRrWOuClW
ToKDEKvMzUTQ3gyCnZdJs/QjSGvO8EpmHGPDuDd26HJRZqGARKQkpDL35HyuKDFP
szD3LiEgPa9DlawTczZHNuXC5H1Kkpeu1QyGgKJ7h6hECarHCIWWdgfXA9X8Fah4
L/p/CsEBR4TmJ7qrH1yKV9410LPDHAHd0QjD9XEjhbJEGF/ipZvqFi2UW3C36LIn
HqXArbNFFGcpKoqrYspXrfv+qbSOrIUR1vAPXev2GGTo3K4rkER2lFS2pidVomXr
zs1Ph13Qvw0EVQsGaD8pMrwbCQ2rwDnivpVpPGz+sK6hE4H6VnZIg7gwVWpXc4rh
3YVuqoi2v06fAyburCZNu+ZG2axB73a+fhWWvJCbJ6BdhowDwGO2hVM+LouoEDyP
9xXfgtLcetmnkc7Ji8zxst4e0fzEgO0Pkl6plcfm9s8a//oMeW3v9zLmKdacy5dP
e6Jyf51Nu5gwvZd3VOZGywElpk+/fLxoSrIJmJ/qJ+Pkqp7nMdF5fW9b3c7qOTP8
t1cQhcEOs2EmmHTVgQKGUO6SMa1bIopvbOvXvlmnLTajIpXfNdiSpl9LtavlIp3+
35Xzj97rhhI/h3Huf8US+kYQaCwoRmg0UuUWGsvayi8MxKfLEpsUf7XxMV4TG3Ir
79KDWgkDpPl0Ds1z3Csj3M+OiFNRf4PpsSWhnW52zRDfZJz/ZgPdCbcf7bjO/u13
P0OzKcVcS2PLa6hi9kDQwMTscz5bQRryuLI278C0IOu3RERtscg6ZlqGcwZEomdG
7oGYpoHCOFbUQ7LcegS8mE6A1JOKucoSMcxkLFDLS1TR/nTHss7oDnvnBRxnLE+C
BbeAOt0+H/Y5qkAdNpeNnyC+0zmCgiNhfJbtXhajjNFiPvK/oQqINGNDXaQhpaTM
ri565OXL6vyE65xE4b9jecwGSqWuW1Cp2tkD7BQu3Qedh3+O7qtApIbEAlIMEbp0
xM4ThldFJsG6CC5oeLfcSv+rPWgr9b7HQPaGUPqTK06avXIFz+8pVj0slAWMTU3Q
IIhXnsPnFKRxU7bALcuR9LDZaW9o8UIibKHuDLoPiwPUSJ+VjZRWSHhm1abmvTpi
f5PKf/ADP9cOO17LC1SNsLuK7LJduOL2isAyDILVCIwfIIOwoKhQAGYRVgXczUX9
uckiaHjfMvQDle5otKtfIOU0EOtkVcHRACF6guu2/oARGI4QpK577/ML5qaU+WT5
bobp1K9xeaLEIjF4kXE6QmhO+U2il4AV85UYeFoo0q50ZHDzdvACpE0mdeTha5vU
sT6PRyh+H/NSbTP2wBk+qV3rtd8bwImU83RqCM4Ilzg3oUCZd5gbfhWKylTwJB70
mZ0AwWVa6bUxKdYME9q/lBmg4APQWZ2Z9tjCcu6fkEv/kLIeTrDrd7/2ZdFCp6gO
VOKxm9cwYyFygzWrLTVw2k5O5LFf4IW+5f4vNa2R2eH1uVaVTKqJQhgR0JWD/agj
p70pCcNNYH6t3h8eUae+Hjo/nuo4QQgpjEvMivAsG9z6wtURMByM+ELfGVmU1tQj
xJyEkxv2qD6SQ6pqlLhve/5lk5a4qnqVGnEcHOcBbqJLaDUhFcRzfDws8v4zajPO
8jw5ZoR9ZKwJJsGo1jfrBWkivaMnOn+kHQPyCO39sc29OoICjMFsSuOs8IGAmU4r
AwgaHLO+sdjXYTHKk5oyy7KSvwXWsFsVenzbp1TKY4xp6jdF10oIilbT6Z32wGX3
Mi5oglooYdYeQl6VyoowhMlUitTpcmqxKWRFie9tMStnRvaQE9RG+tdEnyRGs/Id
N7sYRwsHq73+WW/CtpR4yy/JJC4h6dDxaoeIMtqXb3Xvvdna3D4g4n4LBhRO+IN2
95e+gjdD30ZUmXrSqS36wylAVADwnUEwUjTSxpGqGH6zGD1o23iWlfg9sG4U8J1j
2tIBC0O6eStj3OD5sRP/SYJo0S2vr3kIvz4qgz1xlLmPGouOr9DruuP1ghnTYO9A
7pV5VbYr7kgyKFnK9tqp8peJ05zuClpv/CsazECoyq1e3Dz2TesfVbdMTmuMZBNu
gjBuYxpcsd3Xo4g40u9UWeA95xBPewWqsfE9Bw+bMV/BpLohpxX2/qu7ctF1QJBY
JaS9L/P0Y4VwauTg5K7cDN9nl5cvmVrO4cwL+ODqFP+4igb7HbuFBllI3bbs5lng
1cdTR0sM1QGmap0moetxrJ+jWZluSQKba04llPyRTSKOkU9WemnWyGXOSKCsSqpf
pOaUuhYaMyuK+FXMLlr4aaITIaIshbSICoQ1QQ6zaX01Rlv8If9A6twpugpjuS2a
gBkyQbD4ICcQMnzEFo282/J9t5NlCbA7jQSTThIwbz9azdgJwn6JG+/xTAhti3/o
mZZ9jBga9QrYf2BinqqDGHk98TP0Q5IqGon+M3QTyXP+HjIhGhZyH/d1pnv6q9Sr
4ylT1hK/VW6TGl5BdF4jYY5b+r7Uya8mo208vUK2u9TazsVU3X3Yb5arWy1FlMiq
6lwAltRSbIvxncYm5XxRgzyQ3tGQxPa6/khLh2CGzVbbnnGiF1+NTL/giqr6j1Cv
7Wsst0kQPdG6kJwReNFSbQ8HonVi1qDz5dvBiRsb+CEB/5KM7wFyOskMeBMrK05Z
PSoGo4Tano1KBpmnYfO8hwl/k+fFCQyt474MuSkqr4kZSRAj9OniYSkiyVzx8NpG
6OSsUG+zcWJrtQ4LrhN9TVhSzGcdwpw6qJjmZlo1Sc1baaZW5jQxoHv+GC3Zh9TZ
nqpReiqYdpgBHzOMnf/EwRicgUimNE1V0Mzqb/Kjal1JdrrrZNFZR+2f7zKo+nKp
6873YZpegdezGg5jg7AfWc4MFbhmSFlp8EunV8LncUZMT82bLwUXXGZ10JZvLWj0
mv09YO9dAuEMGxHneA1JeHt3qABZV2Mnp4zrwmQ7KS+0ad+lHzDFBEX5ASdd8MVu
NFO4F52hXWINNGq72pkmbolJm78ki2u1dFOvh/kNvJYoOw7plZiBR5HFqKtWeHMu
mCGg2ijCKArjvPFt5Bar+dpdYarZ/PcWb2D3bRljOU1EV+zS5n4atGOl0JDZmG34
5IVeNKK270V7phEcxUuchIgzk7RWIApy5gx4M4k/7S05BDwx60gC3ftl1kd632uS
Hazv8dPaTK+xLtZNilvpt+zLyZRRcKG3l/cN+5jeUCyLJodCZ+V/IpNERNdbAaT7
c3xuJ59g0PwlVFPqOdGKm5r3BqanrQGkn8yky/DmrFL1jKVQsW70dDynCsMUUqKt
l225No6gDS2UkoX+e0phUOY5hsN2PVWeEYmkW6E9z/8k/JH87YFnUVv9527OdaXL
T4YX0YSDE/JEOZykoaL/lQzDmGqYoIXDOY3O+sXJ+HAmCTHTTavA8xPtXWwcl2o1
nA8Ju2AgqvbHCVJKqHGjt2vadnxrw2CqWQma3l0XYTRsxx3SCBBvl4r/zUzpoegE
KTlng4H2RCQvNzAzzF7tW7j9/oode6RYb22DwQSHxhr+Y75uhCG7V/eADNCYBMqF
a3WuKOg7zi/398mMGMN8OHl0Uz8a5AIy+jbgRXeUU4hb0untHKbxuIdn/ilaf301
+5JCf8qeU22Puq/sOvho7TpqsExP4KMv6zDT5wJVQPHXgaEwhuxKoUjbfzcXLKC9
EZmHRQCIVuM/l/ckFS59PnF9urGjpuFMiH/h4bbyHjF/5nN7j62NTWSP5ra15hXz
fq6iOqS9t923IbtMgPsyBWD3NxLRWJk8A7oZr2r9Va8ydAk7zM1m4Z4wqiOOrzZf
v2Lkln+gQHHlB6fCXnGpmiQhqdXmHcXWhEOUK894UKJBLVDLcFIfgEyPybF0aXkE
DbMknZmX79/x1/CB7FOJ2GNoKzTd6iVah0+BhNO/qNu6BD1OvtG5W41RGZAlfSaT
5GiMDWiBG1oO4aON7E96HDmTms6P3P5mNJkcIfXNh2ODSIwcuhs8vIShlFDPrZAa
fyehPKSmrHTJ8FITnvhYBAx4msOc5jP0wL0fTJ0M1SygOTWQlXHKgraNM0eFpHcC
/dpY0J2NTP84+ufe7pVq2YbJkmGZUJubf3czc9V0PguvJ+ceLRA5bEjvBt+2dNlq
eTv+WJ/lEJrUQUddRaqu6VoHy47Y/cAP4t1f506dwrbpRMm3grPf2tYwMFTVVkJ6
Xl33BkVitNZlJbrgGozUS0ZqXr42YWrtjgNeDSQFpe5WsasKwuMAGgEvoSt108Tq
VTbAszZo2MiwaxdkmdbGcGW4z0oLnmPVhRlzWcR0knLJ2tNZxffdj1tLQMqygD5v
gKRPHyr/k6co/NTN4ZhUR9gfGZbC73xxAY5feb76qnISamiLoFRoooExJijWYWU9
tDpmFmfbnL1zd4Vi7CmtKKuGgDusskKkUbvH9uMXuP1gUT017jctgcsDuQl/iqmo
ZWROASvUY78PdGAbTPn0F0maMf7NSACQgqcV5aEohehqsXKbnJ3HJyePJ+6KEtqW
KSRALcGo3VDvub8e1DStIC4T9aqby/2tphX9JRlzSYt5C6SGAdED0t2FWSOY2kur
vU01AFcTJIU5pWMwngkHK8qvog1yvR+enwIAMNMTe4xiEOmXesutCm9SXjCODoCu
H3Ampjp5geOga/oB8Mu/KQ6Mndd0hl4DLVv+VHcMsUbJOoNlp91HRvD57L6CrzZD
BBPsXmCGfKDCjR7FDbbHggRxUV7u/yBu/KTeTJQ8e0KtCtS4JCOROntJn/p4/2jM
5adajNnP4Ry1owJCzPRz2WZ226Uy1s5B2wdFX+LOZrEPPqVLZngS6P6GtKW+Ui6N
SEHyR+TG378TVadOA/fIpjRgykAQFiw2MGb7SyBJaJQK/tu88lCHYn1yrLHzwlAj
CJ7FZGonuH2AuR2KRp5mmzqpd7X9qk2mjWLor7vU5QyX3QBkYom9Q0f7cUrexLGA
i4Yc4HKz9vDzeVS18D1EDHOmYjucMlgvuxblLgvKs42Qcu91JYRdUB/hLEDg410g
DDLbz1zrsLkJoe1v5Z8bl1GXNbq/M7Zo69QH4BbEwgwW1XhaOE0tWgRzQwR0oYz/
j60RpdDdVRsrnUnw5zCiPi5dQJF5Ii/Y/SIfNeikQi0G28gg4qEsw/HE6xLA7FWt
2FlOE5UkEe5hJL0x9pdUXXYC4WvB9xsQC5gYUS+K6xDkkfQJ+GoLW2P0AI/s8KNX
/zfBb4Gp7UXeEfJXLihN7gnlL4reg+xNFp4Y03VJqBJdqazBFetQHwFArdO3rm1/
PRtMv/nQ+oNmnHCAKiPXEcZe8IEdxqrs9AXDzVH+p8DeAxXCdtsgg36nHeFWr0wZ
sYSJEi0UV0pMYkEbUIZtsgUOpQoDV/tRC4L+NXTUivZGefLHJWdBgYoIJhwpJ70G
VzzWmMCr6yiFGv95EUCEl7nu4PWD2G/7HjkhlOkjWt7jd/rGXqx7QtC2Utnt3L/G
82CfzV7tVgveQO/lbURua4wAaAVC221UK9QsGinHwlA88aZORHGQCDjNJg/Ks9X1
yJ68SPGVpVf9GB5Dgt+YvwyJJCZ20lr9akmL4Xuknre4Oy/wUiha9XcticcC7mM+
mH3aBhPDf5q8xrPtPIajI6IGj8GF9Ec9sJzgJBdOGoqFFhiM03z6a8eJuq9nGXQV
4IZEK4K0EYeBdxl3QnyC/00/w9J+d/mMWJPjyDNTPaS3fr3WGRv3Eu6AkJJdS7gV
/i6rXtOiLylEMmBH/FgxwyWh1a8eATxi7oM1pg/03KRFoR2V2nSWskuncLuGy4gR
NDLFe+5wH4Q4lLEe4e2DucrfUahyjd2yOdCVboBZUijecxYtC2sgFmPcS/nPiOWG
GhTpoXFfNe3LQ7Lf015YbnKy94nl2Acedq5jS+WQXdblXpWePKCtFv62FP3RFk9P
7FugOTW0vbCpHhV1shngvcbDtYaSIxNjZ9Hhm07cX/KM2jvGYdMNinS7DhaP5l3N
WDLvfABgk9TVqsjpNNKP3PzlUjVSOOx0OHsp8pZDQ/yKE4izHDPtXiqnEefbTaJX
aeTTxPBuNcq7cstMh5P2o24gDdwJFG48Lc8lo8/sudnmIYSorMIVCSkQArRi+s3A
IyEaPtvQEYi4yC+aicKXgaYNkCyOgXRECWEvR/gZ4IgY1O3JljH69BwhX9Ytwp0m
QxMf+n4Fr9t1noZslEE0YvKhNM7QXsW1PFK/KEJBCh7FWFfczaxUErp15OEpFkaS
JJAd6M4jpX55z1mdWHnpSA+p5zkKuuB4qYUFDgJZPJHcqnEW31gLBOrenkXCZk4T
wFtiXOuxLGSzoiT9vBrLdNhRphnllYa6arLi7YYWrdinGt0DxA1SQvE0dFPW09G0
eTcJO0874Fech+kdQ0VYvB6I9EvZaOvcsKLW4n4OiRfNe653CHukdcSUy5Ij86oD
iLoLxXVrPPpPBuqqRmKYmHUerJBCn9Inom+CWGbTKUvFLtK0RKhJej+FMO0qxMUq
ltojNUtdKE7ToEVAzvzInxxuYeUTih6Zm77ydBjcqanDaxf+EVpKNbCUWC1Sr1ys
tTPM9q4ClgQd+9PvNyrWBzpIlkULBa/4Pcgc9YKTQdbDIDI6c67ZU+PrUeKw3eoP
9GtigIR9V6mTYXlcC2jdEJz9go5LaD3EqTvQuCnB5tM008xIj7uax9KsL05v69iq
VqWxXnS7F9bHkYpeAqDJUTQxDScVk5Q/qMJtJqFzFq9ElW67cFofCDc2dPb0FjN8
QOq4b/k1APHgfQIRhB1aa8bstiWp/+Tp3ta6DZ1VyvLJaXTnvWPXq7i2Vgcr9fQW
zTZIfl+qvL5U7aqBlI/kyFKU5NoO3qJT4Tsw1A1eulS5jfG0aJlQXEMnjUL7yML4
hNa3KT8i3xFSPQ44SSjiTNc5vtW004isC00ENFRy5EDlTrmzuqMOyhQVUT25INPl
S4YZBAZ23bR5lV/XdzvWhhHyqdwoKNMSAgz1m4YRYNbVc0HjSHgARXWuqojqxzDt
qmuDSBkFMA8kAi+kWJSWYSqMlX9XIcy0laNtCZx829Otb5oYk+7AFvo1Z2IIuztl
V2On7HOVnV/CagbCtojPdyy3fs45SgfLnNLd1NKkcTGEgCvJ/cdloSz4fr3b9dcd
RuUaTVP3bMcvbao7+DzbCe6ijc0mnMnOt3N9Oby28duL5VB1NEgXqVIpT8BYL/H3
DQzmSET6Vjfbo304N+WD7O4SUe+DTIzgIqGM+8BDOpr991ShUNitC4SOdw4U7F89
ugNdKcJ/iihKdgZ+HVHvksCMfvotfoAV7D+huG89BMJp+yVxlxN2KxEFyeYBHxHV
G9Eo40ZtIcVuKLz+n0OimL1Duv76uGqWjUz2IsoalzHYqr12HqvRFUGERT7avsoB
Bpvv3qM0VJRYRxf3YVBbv8jlyPvSzkH49mgTW9pBTMII05Subs2mTkVBUzAw0zGv
cUVFqK4qxGDkoG98fy10tWWRsPC/BEpdGi8gE/vJTcbXB7Md7+x6uzLOg6Vcxg/8
y9jGXvpA4QsXEnb3x/gD//e+29QQDM85Udqzjs2nNz5LVYlSEUKc+Fr/1CInZXqT
hSn9Io/RWYAgwrnRSdUYu6uimqSFURU71cbvuYb0y4/3jHMpEdYUA043fpTQ1Awc
+1zKD+m8QSbWgOgz1zZcOL3sCWfqKv2hiIRjqLTreyAWROjvKfY3HkOGvpS/cWvl
GLrj47nUQ8jJ053PASy9/9dM6yTUe8gNf9kM9uKihoJMWRvjAOumzlPRdK5xqplA
c0TEcbHkTa7eW0cbxvMWNRaaw9zZzmz9CJGqhH32gzjIufR8Xgd9qRF/xhzbKT2X
YX1AxF96nmuUcJMxomGVvLwzkI89HSbQR8fvMftq9E2wN+/thI3JnWDuvJ/y7PjD
UXP0FiZmCd0kv/f0bhxQDJSPze+OOSy9zLs/XYGWtms0ga4LthWn1Dw5rOMrwoY0
n0xhn7OPbQInVCB4x95sqS2+QqxYaGzocD2k6RIL5FmjrFvL9WaBJ+jeEtKUt8F3
G2F8Q4rET4vxXJlAuv2h59gbepJG+CM/vdQxbxxNPMwTse2VQrrfPNA/gZ5XK68r
u2XHmk4OhCAZ2t+hsxnh3ppt8zvn0OKmQhab9kojdZ+P+beNxptwGAc8iCVNfF+Q
Bj8LwjUM3ecIxjYG9xz+ZqH/VKDDay3Spsw/xu7DxyQJaNBXW4fn8YCToIhNnB5d
NAUOYKAEBYheGAJz4QAllbQyTyCMVn+HK90m4TK/2c4GCgwQNlKyfytMJlbpYr9X
nNEthUA/3i3tTIyJqdZrgoHjBCwR3Vlh9znPmREqMZPoKA2kdNOulPbCyyqziqwx
nRA8KQqA/Jf8ji6qry+dvRfVKYnOHGPjti1s46Hkc3sOJtXtC699NQ3JPu2xTqlE
tB/f9T/UOawIZGpKZWoADeFoRIjwrVCtbgw19mOU/JShtFRGPq8oYejwHHLlJexb
bhSUjvxEcg1R8LM8nP6S4xTWMsmN/+n9olNwEpzGFkOWQd3dTjxrqT/Zxhr0C5rd
mJKZhRpzY6BaDvbV9scIfr3wVLv+GSoJEeXVC/2/+By8rK5O9ga9Dhr5FkO7EJtw
pp9I5zh2GgzOeXQn30vZ2+/OV/zD9vJ7Kv8RvZY7yjjxUPJWck5fKscH0/+YJsSs
N9Nj5gH3l20Dp1CDZDyVZXXaLxyUFSY0AUH0X3V8UNSMPn/gRzCIR2zqlxEHfS0S
oewD9Ard2RoqA3a6sC7VqqaSLfsaXUSnaX5TpEqnFIR8Y1asvLpAplA96Z3KxBxx
Jq3B4JoL6iW2tve2wRAPZqSZ/gTMivHBPF/dnHQSMDDPTf+NzvZotaZ0I0ZVTr+g
dzNH0wLDqAGtZitCOQ9PrgiKwnbEdNp4Po4jYqEAuC8lhenRwACezFp87rIYtbFW
`protect END_PROTECTED
