`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Wipce6a7TSp+yKlXBU5Zb5gqzUOeoxvFN4nHlEV3z0SEqW/5f5DIKwZ23SNn/X+
00iFpTxBhvPh0TD7bpmB8EV54H89wAx5oauhbg9vRwVlW0wLmT9jGtLWzrhMKpd7
GEl3mSsA9LVpjW8K0OGSLoAKNgcuA+9GsN6CXyeOTXsrG2VGsr7DQr6DmuKLkX1A
dA7NQQcu+svs6ZZIveOueuTeQMlQiheOmRnTZIZjDAYLEFKNm2hLjhEdAtUJVKuv
DYQMQ9kS6t5ItDXnbNfVYXZIS63zr83lenK1U+Ho5yxbsW8asvpvCD6iQLo6VbCs
rpRZHmcnPvJ56obaSxCtFv1SKZE/I9PjAnWId3O04LxbrO3bnUgHEEDB4sorn1m4
WyEmMcdRsOpHjXrOlun7U1VlOQ1u/2H92BYoneBv5S09w8Jp0s88YdMSCQYZa+z3
rUOZF3ltmQI+0sphMtCWyBOen33hP2AN4gi/JxSI3skUdbYm0M410HVdQ6CvQoae
hrndmjsrHJU7HInHG5QbUMgmgoaGphXiACiLzw6C1WJ+VCntxgaKYpAlQdWpT5qO
S/4LULLSix5NxR1cL2DnYXSM7SQswenpGR2fZWQ4/3zPLGGOHkLlIwT90hygp8aI
ixL8HIJ9CfLmoH9NDdSGWgg2TNL2LNG84jH+3BqY8vOHRAS/lNrIrF7BSk7t/aJO
ipDDuXBaWtmS19bCopBY4D38POb6lAYV4I27ySALLpMKYAJtEQmTdbX0ibHwM3AX
6Bw8MgTkn42gP37kM7QHBpbx2O7nza0V9IDkEiRZc2RxGYsmPnC1+IIKWmx0JsHn
/OyIpbNB0++XgrQ6StNSbw==
`protect END_PROTECTED
