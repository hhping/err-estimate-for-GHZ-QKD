`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PWjHgA/fX6yAkwNOb4MTtYOTV38qywPDnIXijm0dNCO9IsMOsXH+cjc2nzfowtF1
i65S7uLH9dNszXduV9mvZWL2pdxZTyCzStiqrmm1DbX1W9X2t2gihMB2r1n5L6nP
8qfkusisk6rhjYCWlU1DHhxvBGmY3mUWLpMLrKnZm3aFuKc0jpT6e7Q6l6jLuqvX
8FTy35RMasMHDcI7KegOe3KSd5Fo4RoH1MYFKG40wc43wEpUs3qz5gzFOiWHHKX+
U7mv+3jz0in0DFO7EinCo6WDsoWAJQL1ZSLB+XsbbpNQUhfcCbJPwC8OW7szGniJ
x5b03PendY88eFE/qd+213P7/y8M8SC7mFylBZjpfs1BXwwOm6uI8OpzybBo3YUx
bExrna56GQF/VmYLUQn6bRm3zqweLej6sQM1R3u7DdU55RSW42KOg5pCN04pWCPw
e+R0pBhoxmZpA5j1b7tFmpAKoAM3dK56nYE7LrOnNB94oj6lqXauZhC8xEhoYn3l
hN5wPAKsnIoo9OW4uZrDlVi5mmyGR+5gqZ1MANQN1RYGZNv9BY08d49bgQKcp8kd
09WgvQAolxLV7dxMJz8sbaaUVWSnbNHANBNPJXP2lF0lwhXSx+CvEjYyFji77KPj
OpKDuAMB5kpE/MxOEfwZEHjfE+Zofr8iv2rSobaw4MhRdELbnX7Gd7cY7doEtWAF
shPqoEYXRzq2zw0DYekJ3e4dsbyHVBKRBUmCsz0JtmHiolBJZXeYWRaY81DbT4Qt
DsIbEMGKF6Ssm8WcFHSWtEOZOF1AS6DhZGECRYO5hKIlnznrLXBfuYPelOC98ELY
z+u36VeBkXQg5pxjkoSQdIsVafjEIRbxE8upwVIKwtbA8M1OxEt5GBO2LJ1Afn3X
5YZQfdgrImbUo49keV3N/hyO/yQp/MP1KYgP7BLkkEOQwFsDQ6oDx6thB5lr09v1
PA03s4T564tOyjpmLzArdYM8w9H+xa48smmpDCNPLB2VmEgYP7rgKLLgV+bQQv4x
RqGLnsjzAAmHFNpVM/w0ekR95/G118eDxrHkWei5xAVCtqc8Yc1H4Yk+qOfbn9mg
QEd+Ljw90tp597hAy5fea8vGPmGZgd9/nRKAFTEtlv0De8N2lbHQARHPTHphGSus
j7nxofAX/meZD9BjXSsQxsTkkH9zgD0OksyyWtbcg1L42ojEEJCMhMddSzC6lSfa
HV05PbObWNNMrCvycS0DIoyv9Js+ZzjCt2GPJg9Pl5r24HSZM2O4iC1BUPEi9/E+
FQ7DThYNzr/g2axq2Hz5NnF3sVmW2pd25Qs2Cxnz4PpXBHfK8QHquqOS/WV+Kkb1
VukeUVKVuf6EZxylQPe9HnIA//xiSvyzVdeM7XBE4i/L4gX5MhX+BF+jVhvFl8Jb
bssZjd6BBuaT/svgnIbkbn+4lDuX4zoMAliGDn5ztxQf4JbKykLA1CZUa4itkPhD
X0e7smwjR0fLt5BSLq5hncKlMCZ+r3F6hOZ+IBVIQ/+C17rNGQF+aGItNrB/EjbM
m5sK7TLBlnhtiDzMMbWfYTgyVACVcKqp7TNFUZOw/SBak/5kCmnQ6Mqs7TBggWy6
tG3R5OpVZs6zY0XhXGeKZmF1o/L1Wb/2Gm/bXrAYU9solzlZIjwtP0noN8FXIKw9
nWEUUIqMxmu1bNG2WyN3aeWwZc4Ptu9o821ZF5oZ9FNfa6g7BSkHR6KoXgqz4/FQ
yT72wZ0hZ13bJPygdZexS/T/E73TNuB3GMXSyqLhhEIbd16u6a1x5rzYeIx76ZA3
Bmyf6UB+k0BEYUsriLAUbpeWBtrGu4cl4jggjkMeVyx2dM7gr2/ysbk0EM1rdTN6
WjhTQKYJC7PUvNZqY+OoD4sI2yjhBEOYZNQqHTwADD/mGCK9x2Xhoq7PNG46j1L7
4cnoSxiIc08XRdgKNV5SLjYe0w59ekRVA47t0UX6LcrBN18aeZYWNHNu/vS22wwv
IDRCKt4XOwSse+ftEfATHDqmx5LI+Z/4wH1mTXZ9FGrei+iiYQ9v7k27Yymvxc39
HfQi/4KMGim3OoNYUKYOBxENy3EU6/bu2CK3mR7M4KSGf5VLGusTx9sQeRb0S6D6
J8Y+zHBBSUmAHLGzN5kVq0EpuJposmTSQFn7oZVvaMdO/rHWrERw8ubaFmDwp4+b
+oouM6SShSboOqM0LC/Zw4jChGC5H5ThFq1bWBt+fO1XTBAlS0DIGmjfsQ5KNk23
59tTSfmXkSQaePxpg6jPlnyYNx1KCf1dXObxCpwLZkb4MwUVQtFOf4PNzbSBWlx4
WfWK0p57i1B6lAqTjkA543blZvNMM+maADXoBJ4j8JLWqP/TQmxT1iXJr/8Ys7Ei
mplbEVdFNvrs9JtwMIpLe6GhFYPQNCAZJZ60syA3o3jld4+WKByfZWhggl2Gb2PN
fIX9RovYvPoLCj/tB1l5IduQD/jO6wD5FV9NOYxEmGVKKRGbV2oHw1xenzA7beax
lvjtQ5XOwXsUVieFdAS4QQFXJUDLa3Y3odvXfFnfXu50sfTlxHA5WdQJDfCxJh7R
Og4RAg2errj2lwhgeoNuUEmaCHqTVSlkSaPYa617ygPCmbOCTS9oUev1a0Y3qkhg
bpPl6ZswvYQH8cCZg2Hc9A9zuyRvHTtbsMHsXXn6ZA01TDQ2ChVo4dswdHLwj4Zd
QcJLCmAYTb+tCvFL1slLOK5DZQukSDPhhqe4RWxPa7K2hG16FuTxuTEbAWyFpCn6
BOcwPbj3mFp1GoNBXBrtcUmG9CY7HemhusoKHXh54SE5+7F6Xa7GynYvzommg051
1UPae5ahAAnxW4fxDBvic73no3tnSkOKdL3M2SMhqH+D9sYDTV/LK/2Asq/VM5j/
UeKj44gJbKkWSU/b+7kfJK5z54/RxSVkgZZWOi7GQqlDOOyJ06pkUHCGPtoLl7qc
eOCjPW2H7seliBYV5aP0zVfX/sATW6XLSftG/qW9+BHdlLeFhekvBn0KYgmggSuw
ejG9MHeVZhQ6fipxhjeyPjOQOBIwrAzG12im0K6YE1DNpj6fdNkudcoQdt2THCbH
67PdwD8b051jsa06XjZHFEUK4gPnWFc7Kik+XDnjmdrBf9eGFux6d246NXczyNHJ
d89EkTOpUO0YRMNn/yYyFNcMFnPLT8k94MY29ysGEOWbR7dsVGE1CjYAz136N4Vc
xX1+8eeEkIeGffj5pYdK1LgjvQH3Ew0I4SyJSu7U/ND8Rh0lj+R9em8VizU2AlTU
aFGFDBgfkHdO53koNgqpoS3bhiK2Dr5umBR4igcgrDgJ+6UWnq8uGlmI4aVPU7V8
hYU1HDRFIuOyr4uWHPKFzg11eWbIUcRdfwGAYlRJsu6GrW/u6BwBdoiWCU2KAnxL
lvdWy34Ypr9crPE53HwttAFCJ4ACw9mPYP3rVLHgom0jVqKyo0TkX0kvFy9iz22O
xoPvl37EZBaf8hKYaAgU+RlDYUx8nzw7ZphCKUGkCzSEON5/fRMQfFRFXYq9k/2M
Oiz5gfQFeFw0uQ5BXtKrYXlSb4MOtogp43u0/pMsJa991snTqsG+ybbDu2DSevyc
Rh+xxOSJw51Pqv9dcIum0JG61IawIKxjzpDMrpds4SVtSMLEMdsTQt45yM8/1xNT
QJlQY8weYLGVVODWINKWZ1aRiGPEZGXLxCdhiraL7Z086usnkhmfThvDo5k7xUdk
gad4/wcnpprpuOfOANsJAtJT4lBL9/T9k1IMu4A24jasEHIphdEI+aY86PBRXiqD
IbTeVs7+55g60j8CFHCNYY2vReZcpuZgh02UdKGgS928CLgCgUXo1IbyC6lvH94J
4GdiinGzqcjL/Sim73mbh1PwnWmarAhxjzgw1tXZaPrN86le51g+jowoJlNWiM46
KNh6KTpmUTQ7a/ZdhaFZwzvz/+KwY4BiTnxliRJHJF4mOwSG6sWT8gsdpMeLr4T7
ozUJKI2QQVyQHRr++hyEsq30/IwO7YcSZQ3seQmfjeikbHbV8TYs5fqViAsMaxd1
RjZifXRZAX++ML5lLaVDIQ72mEe8CL7Ej9163yWSmWmXVuQnMyttEma7M+k10Rgb
Zc4Dm7AiOhd5+MoDs5vov+PJH6iiSzM9+LCYJ8f8+Lu7/IMhCvA8DZt3uW7uiDQK
mM+9H3TUDZY6wssHni5KjZohFncetoKaowaXg21OTiwKbpBj5kZxvYUZfecdhEtU
RHVYtufi+d4h4wJL7/JcGNTs/VUV+S3fxVlEVR2hxi84/8iLUzlMzBLpI9u3viAh
tBEymS7QSAhXVxDiT4RBcZYYlvZTXHF+m3CIYcABqrGWWPDZyUM9Tbnv+P8vAlzK
bPAnp2BWvN6b+HTKY+HfO0OnKU+w1x3EW2hbDXj5jH/JCsuL0uAsav9GWS3G3yGl
t2+1ErpkQiRi7/M8oylFR8/8IIRedMDvR59t7+8OW6TNyMBiji5waFjBpwOSnDEV
mfG6zklOc883j77YnoINmiwhFqCX7/ZGSGe+uXVciPt659qNzRjSX7kG5JMzM8k7
jGaUEfA4AofVvSdZMSlL/m2IbCEmVWJWzS4VR11anv+ESYfLktvpoKkIxBFje9BO
5roRy+WQQhYr8HQHEWrILrn/ZXL8pY7Bx9IaNE4wGmrZTRCd1gow5BYWJb6sVBOz
ZwpJjTZWP9Qn9cFnApWRK8rEGsSp+n0f+aiz4HJe1U1C89VnsEO68gVejBew7jE3
ktJFS1EUI4bFWrBoQBW4zD4Oxp4cAt1D1jgKLa5/P0YP+MUUwBEBhReOj4jRzC2h
wIKU0st2A4L14GwH7Gn31/pf+0Vj6RQP0417m+jvucOIhkpf38qS7uSjMir0wlXC
H0q9GrXokHF0l3uFeO8XPy/wHuqY/+gpuBQK33M0307z7zgkAKXAVfxWhy57hVZ8
Dg1LgWBL8vRuf3t0anbf7mLJWx/blrSaQ5V2Sbr+K9qr6vOr0EC7MuOuB8MBpYM8
IN198MI5wyTwEYp11iNF9gBCOFvrwZtYFotvbd1OKwCqq5RuduR0/dYTyePv1lLI
yJrSMO+eSk9ziqJd0w6zgmhDQ/8hRtGCXB1dTQx3AJs25MUXWyvJ7YuDBnnsnoGf
qs9oxBwt5nL52KU1178jCn5zex5IvVZGAsKwcGa9iVcr6XelYbXPWN4LDciJpbUl
tcA+tOc0FI7u7CVJNWXz9fH9nUyoLFb+mgw6NXIR3TJ4Dm0vCjj0k7HxeDVa4xoC
Xmik5zdYtHdYz9Z4st4EbDPX0BYPe7zkyWK1U6Vbw5DYMSD8RUMYKwUL7vmnAFBy
h9hYedhCRSWmCNLI2mcNnWYsbStOeh30Z3cjjSTOGgjgNOUl6xmsBZRV6Ld0zHnb
us72eoXQ+eYAvchoM8Q49f0u8BzW9udeFrr2mfcv1Nl3G5gVD6Vpbwd9DjqxO2o/
9cL+Yk7t8PjgFjPsn/wdG2JjqYO7LIKEg0vCUYYyl7C3ng7fiuwbth1r5S/uUxrT
NMmokdTwienaxqBMI/yvtTnpbCMe/Gdbp++8F2M+ZJjWj3Ub4/rocyEyFKLV3oqZ
sT3MF0OnFOvCeny8kK2ysJi02MTBvM2Egb5IEPHNxXUI5hHdhqIaODUHw5+WdlBm
jcNFJOWZGLQvcCMYeddrucx44qBnaT3w3uJ5WVK0TSOvZQyoC1Eawpvsunk1Wa5X
ibCpZjecvXNz5ni8q5wKofGRMW/4Tr64E4MUWFC/X+JYO3sZZ5klBj4c5q2kdObT
P28mGn1mr2CHv0zqHFJm7Y+K4aK+cedm0YAQxSEt5I8nAFI3b5Zl2FoSUHSzTBXf
onCEUxkIlYE0b7Hm529CgCSq06YDe9Voavz5VSI8fd9jfp/a2g2LNUcURkvF8KLS
SQ9HuV8+jn983ET/ODUfzUYZlW7ydqatLVRZ4l3A8gbu3Qmd9yUiiviOBoExwNV1
Za+7SfMivGL69dqP4UTutSldu8OwHGWoTW924mz8zVq3UJKW0sRc5ElFAv3LH1lz
5UouMseISwkz0sqjSOnz/vUILinXA2SyulEMViwKsfURofC5ZWO/mnvZVHkjZtDh
jDe2utQmB9I3Sn59X66OtknVNqsmTHm/UTr1VfzQkkCm9/M7JHq0Nq6JAgaoPuks
zZY5PdE3u+8itafbBT/I5GRZZJt1TVR6HvJML1jTkRC0toWP2impA5/oBlSayePx
gSyuFAt8Jld2i3n2nIT2K7+1XJ+QLJ8OAEJ+Qm1MQwdAipzs/E7LGvONu01YJtxc
pBu2IltWft/+N1gnSeP0/W+deTXS29WooYvQ7IYqAImtpXXnyOS4++PMR5Xww3Xb
WR7A90ilC27/cl+munxJ5a2dcFTLriO4plUhhGfAMtAjxeejpCJTOwB2opPNLkfN
Lkp9FU1piK/cYEHmfO3j1+fHykAnq20s3E6AJsu78YIZhvZYcmR2CkAb0QFhrbYd
pGmT47nqs3Rn5YpqfAg/V5fPRdDd1l5lbhj3DXMqXrrYV4ZqIKduggPQ3K/O2WVc
sMdj65rlVcRiB5ZGuqiE9Iya3M8TfUAWHCcUbS+FBI5GzUyHlybiqk0pjLagtWvg
Z5VU1x5v2V5tEbC0kREaF+fZMjmcSdzlFm+P+GWuB7+gA/2QsqjKGUzpBehxlcA7
f+7lSzewwQ+rO1VVkOuw0Cg6o3CVXBY8r86jCzJHEL8DbWXXMuwbsUZLC9G7c8B/
SkCWEzlcd5ByGkwbyg1yrAJCDP9oPZQclZ8+dJSyzf5lAB31zI3KRNoZX2Fneymi
eJWSo0IKo+EpFCZPaFqL97dFb8gDylPfnH7oyu+ajjeARkOwox/SqRvTtUmKuMqA
CE7Kyu9BcJs1Y/gfnLnnBzgyWI/Tf87qE/sk2ml2qhlUIVCF9Keh0zI6+KjJkmUt
RIc/fnqMQj7/Rx/iYu9WbGDsrHv92i4GP6+0byPX2cbRUhbBX4XNX/1gzmRImvrN
THMetcBlzPZWVG5q2jZRZx8lI9JjaeYC5YK8dpfzkqhLQ7Pc202yzxXC3WWIGMcN
HZ0NOWCmE57WOsUgLviVUXK3+7LMr4+zNzZIXDHkE+wOats1T1V/SlopUrALhUfQ
fQGNU2D2f4r04DFAXDvLTZmeED57NqhRg6TTY8aBoB46ygI0S5s/PdDvDmS3Wxfz
3ZeWBB/r5a8Kqoak72SUD/zIKB8IFymwANEx0VmINcUP7ZAUbSEznswopJTl1b6C
S83EYAFHvE2EebwQCkqshmWttXfOALxkTLq84CLpA/4WmagoBS1Qx9DqmayK3Fy7
kxO8AGOoBYvDLHyiL52EKuLL+2NZcpn6Fzc6kWgLoHZUnbf0TFxqomfVDKBMjaK7
2imZFATPgPR2Jqwn9aBtd4yOmj/N7RNSVzaqR55n/mlWevbv/CRg4oLd9lV5g0Ld
QZLGynK5WvF6QY9oR9huGfCnoadVoQeMyk0+viMg2Mfr+t2li7mTv+X+qGhSSfBP
geB3H7d+1t6X4LiZ4ew4RgeUr8Yf/wQRrt4C9DOEgfpw3WcjK3efYl8qifnir+HZ
KRbqh4JV6VKBczvInkQmRDaDkIsRCAu7Fof0YRSeZB+2cKjDbfBrMkC/gxPBJ+Ve
JZlwDSggDt7ZIwaHd9kjXkpglPtHyVzRHYIZoMiAj22nhsDJ/wx2hlvjIz07RInA
rPjD4x/QNqSHYmyt9sFQHQmbxHiK9J4NtZ2DSfo8A5eJ1ZXVnSPbcmmyFM/6xnF8
878ItrUdCllF7kGnW82Ui16ljPwhSJZLy0VMFYzUkikRvZzWsbepip7bd6bc/mWi
KmRMBiyzKUaX6uhcc9QfK0Cuj7TYGdox5RE2QAmBBO1g9fDqyxXvM8uUPJ46YyMl
ZZBgpuBGkcrJ0dEL4IKoz616mdNMjFo9/M+evLzWj7BbgT7tc9mPMTcv+wYrZa5o
Vl2hELGI8lngdYsO/GIgrkZoaE/AOsyOUhZ7AcS2RLlodoFBFKWDDchBx4uSyaer
Bb+am0YnMpJ+NKFydeYeBYVPxazG1nSFEV9XgbitnOfjr8wj4ukokfzWtNxfAKyb
MCyof6fjdXJN61m+ZE7C/ReGlCXzXJPKCrlzwnxOV+u50Ra5UN0UJ9Nj9LjmlGE6
w1ZD41NBgMyLcAnDlTKJklUArv0oNqQMySee0rG6XeGV+Qgp/W0EVVxZIAH8WIdA
cY/cL7dWvMo+vyzEEesy7x17ScYzo8MQ6HAKGEhpc7sEIiiniTOcapG0ashNXQEs
XoHI9+SAtiO4eMy8s+LLPOI0om4TGwmzesa6E+oqLjbcWRpxc+3+poREcPtJkwd3
JAyUfRLZupxh6WgCzI+s2m/syWYENWDaQx2jBu02BepwZfI/aqVcjhlKaM4VCQrQ
WaPFR8vi8U/PJkGCFLxGKujKHUB53S7HUO6wKDyCpl1k29153Ssev4OxVS5zBXoc
KRSJOBmP0xTDjjquOqTX7EvO0ihQ0CH3XA0br5GoLdNyH3AB42c8tdnSQh+etMDh
QfZgekIaGZt7+w0BF+6JxARtz49TSHEJQ/kBE+tsTEsEx5Jg4jtLEKSs2hyXhBj7
qQD57VnsJi6TJ0od+C/pwMPHdC/eCC2Fdxgf4+tdy3CtAYr9JUHOIFzT5jlgP29f
pzsxFuzhh9SSzi/OAUyjSKV/qJnIQ6R7k3Z005Gus4Cs5zIizO1PnSUkh8wFu1vd
L4Je5c1YmXrSXRwYs8Ct0cA2/ZpZiKzVKSeZl6fk6xvoW4UcvTZ3DHqp3nYgTayA
CLkz8FcxMtHPLaT5d6LYMnX4wLPjbso9gB4TAc7WKEle0Kv4msGGf2Id211rH5+g
`protect END_PROTECTED
