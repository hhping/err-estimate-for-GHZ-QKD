`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MyIft30zABWKt4tV4sULHXUyKAITMn74mn0RZFOYHoj6N/c4FpcFduSrNwGzCne
vij5pQtdy7zC/4ZOO3u/nrPR1vHlwkAhUfUTTlnWo5xEd8GXIBUWIXC4qCghu96A
hFdWjngrZYS7FnOrK08JQuktpo4qKcM0uHpY3ychJLbAl+z12KWIrO0LwRHDSjvR
JRS2AZM+kGJrFxghH1lMpgcLJ0XNYEaD7uIdMOAW8CIWGutJTpO3ifNGorI7MyLR
voyqnycbVESiUCarOoxPBgjx5/8nJYZ1XhGBnyfJ1dtc8r5Zcu0myUHtoye80nqg
b5JGDADyoC47JnLFTy9jWNfdS8ftP9g0qkgCTXP1YwKOt97U3IPue/7/1Rer7FqY
bIcmHbP5pd0qo8i9v0/rdc3qX2XUJeyGy9KDzE0eXMbrGBOHKiH78e7FDBlNKL61
uH5ccpWVcTZbScyZkvmzjt77c16KYXKVy1huWOHUQZDYkI/4nexVFiW0wJnMuwRT
zRaero6eXbS+eR3rL/MFTB7/EMS/FxQdR02cGH2PLJ5dyIGxw3DDsfFVHfBl/tNi
QpddBEvb9+kvOcJC8yxJYaD8WuFVgXOWPuIPC8H+J02/fqTyKeI+Naz6DNrrWFp3
FMKpT6cqaXqZ9cuVXypqrpdI/ewzhLElhVm7btTbZkrAovDvCzabMVULLaeYPPFn
v+vASrjFKpNFTnbNMTwn+wZtfZ+kPZnANJmHvo0EJ+zN3xVXY5FajtXAy3/PjmuP
CdZJVkLmSefvBWQoaSDR8a27uchvNis2meDVv4ef4ypBxFPj2npuKzFv+8JmQtKU
lAC52txBclhP/yHGoN1dukWkr5yuaz5PBoG8QaXyaMUw2gp6SAWwWTvDyicXrKI2
5Nto6ERQj7lWtquPB2NnnKQQ/K74WUZlhQuEwOUvgfpueEnu2bcmqtHrAZepEtko
Md6HPFuS4Wx4ySYrVfEuyfzwDcFCDiV+vm4fe2aRAYuyhHrgYtMO0tIogKbetnUm
BSpxouPs4TGi2ftQM1AexodtX3y/5Yyvec7f+WKaioyw4mrY48Acd1aYO9DZYNUy
Pa++ZMn0l4EoF7v6DnsKL/FQ7s2ZIw0aoai9tQAOsPvlwxeWlNbKHQEHrJJ7DIHw
5/uOOLsoCBT4u+WQEcTZWAJdRHatRIISnCOUFydVPTUe3lu/4wwdmPn1i0t3lf3T
+VOvRqM9TkvrK95bzeN2Euo8b6qrGjTBB63RmNVvgdNO4I82MuJyd+ssjYR+HTT8
2QPJT48bgL8MjPlePBRet7AZ/f2u6KplizZ1lpNnW7g2O2gniU5wOo2iqD7pLLSY
WqGnntt1YkhvWbJZIDpHjnVh/QAMd3vtpbOejZTdXPEoozyNfUSXRnqANZBrX9sA
cK4+4NSvp+F2TSofUQGuXLybOKTR78Fggp1geio1mJtaDAwlSWMxswsBIa+wh5l3
ZSXaUGaH610hYCNWICuYJRp2DZ8kGlT1V//ROtLouau5q6+hY+qW/srownetQ50u
3pv1KE4LwscrcrzvKEpHqMkjVY461oYQ+QqYnmu7uAoBQBR7RGRYZYD4wkNJPpTi
nQFqMYlIYvPRTMXbwLGxsDJJeRamLdSqBEPs4v1Bjpa7yrzwuqsvfjxBgHu8pHb8
FV5F8PcGERkVENgjHexfgvVIMPIrZLnxqPZ8E28UDVOYAXdtSu3d25SacjzYtIbA
FnZQBo2Yzj1JBryYG1n4QA==
`protect END_PROTECTED
