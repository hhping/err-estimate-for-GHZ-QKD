`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJZkli8YX2WwZ6IEGNBOreOXqpngwx1uhw5oOfwlxlvgdSdunl4d0Kvkr/J0h4NH
T12eSs6XnbHN8c+Vbv+kZRIOE6V/cLlc/4rdfmAuKL3apEk3RCvqXhIAslKbskC4
Tv5EWjRzPTJXvvyYW+5Bv+UjnmwJcGM/X7B1heCgZ+rU68F0p4V3K9y9gSee8iVB
enLIA8gHZvMIk7nP0GxPzu88ZPdLh0ehYLT++JhQ2t128W4+z38SQc8YXSozZ0Nf
zOarOgdRGZyqqc7917zobYekuE+VujcSmArGe7/Bc7e1iAeheinLbqEBIPC7Xrhv
5KfeQO+ArI6K4Eu/HV0AyyFqOMxISFan9FPfB0WE0X+y0wgW/ybvl6bPLdqhMLhO
+7q3y3L1JRWGyD3gaiNywWYL8J9c1HQ4fu6a+MuKbL0kaF9jK36bSR03BCd2ypIX
t/yzJIrxvUEBHfWilVTNKSTMFAMwm9mdUtwv7MO3OsPuCJSaR7pGpGkWf26APioT
d4us8TbGfiFRdM1Z4grOFa5BJsEa5CIvwkd6cUsgkFHWE4YjpF+iBzZUnV14clwD
Sii9zF4AE+WiMuz6VoqzqKiK6o3Gaav3oq+4CG+DL8Edp1xLlAwCXqa4rJYEW7qY
teIS59gLHT9kTDlH0o85IuZagA0loA5Uwyp/uvro03Then54TmDEYMxgMPYrLOV4
JQeSBWuUsc5L3CdGwuycoZONTpiNPmTvmkwlm2EsnitYHG5CzHaJOT/FBNwqhaI9
qfhv26rGqoJd7B9I6jZYlSqbwQGHeQ+BS0SY9zoWIEKeaz85QjLg34Vl6d8diLVt
0psD8BKuCfpe+K9IEiy5GKZfQY5ApyjmhMmuQ4X9pHa8mYDWQRM0F6txXWUitiqr
ckwS3n/EMbcH+TomlE9Pz1HbegrfM5ZuEkYlFd0TsRJn3lqH6RDsFvVXDmtI/Wrq
6PVHjdjGedl+7aKMJhimZ419F+FrV2bQ9oHqmWJ4y1G1EIRNLIy3CcdRi7UYdxzU
al6eeHpW//eKH56nlcWDmZQQtGdzp6xjBCXA0HyNqQhUfTXHXHmJtQybtVtOPSKU
ckrvPqEaX0q49q5mILWcPxoCAqlnHt095Nl6u5sxEkSr5ZhvlS1rNRX6V3z587yb
AREi8p9Xn88HDxmY65+V38/yMLYxWAw11+zumhy5oD89/DjiVs63IkIcdM96nj7D
1dmHDVqsJEV2YNx26nSWfeF/5x+GVzJk4wksTasqVsbld9zzu9UOAqoJcI6NJgBN
U1JpTH5lIp0YR/kDzdUFc8N2n2FT7tFiNpWL78xYBreKSLKQGmSeRKNUv+b/0BOF
+8rejrQA6uxDXYbyiAt8KS9xcZP1B95LwC8yDKjLrpV78XROx3W/vju7BGLHpBXN
UmX2t50NCH0JGCt77d1ldP87F/lVHR4CkDTRj8BHVBJNwnyRdC3l28JFerhXvEZm
0XsW3OKiyGiHLNvBBj5/W2MuxmJe0KT00OHTk+aH9N4bYyw/jrEI3D1cH06bo0Zr
gnRj+y4fhCuku3nEcAPKgBlvAaU7W4Crhx7UbA1Q3eOK3nrtWjurSZYZeDb+qJXG
o1tWSDRW0PNWMPJADNquqsy+PmzJfI0QMJboUKhS4l7Ze0gBiScyJxbN3iz9M0r1
4R//YgivcRWJcJz/AzZcouiBF9hGgnYQL6yQ1t+/tKin+mIEtgvoM74mtcQaO5qR
sFQlOGONIpw3eu4WtxF8Q3Pm/QyCCHLWZSBkZxVBp1ea9fkoIlAe2DZSQZeKb5NL
0aBN4Y36Cx8tBXAvuhZ2eeGCAX8ujLgOFfDzWjZY2gSIU8xHru6NGxtNpLrspOUS
qTzr/EAqlfSbaG058BPi/3/9JNu+BnuJUBbOkNxK1Vfp1N6pnWPIvWWA22f8smtU
64FIrfce25ADFvAv0vPwekxf/HwqYa8YibXkgHf0o9c5n0DJQWvIL7GIokK8q5Jr
XRdL4nw9ohIX3+tKWEeK01QgiREcxiTi5UGKV8y8Aluv8zqS172eYQXxosYqkjzs
DAab7wCuN60cW4n7PA0gaLjZysuEXiAW9Nx9SLH/CYDpobbj0vee/90Dh7H60rFj
T/OVTQgy/YoCb4qPMO66JJwHodLjFOE1VUKFAhDE6hkUd7f9KDfW6m0JFw3BlYNL
yRiAX6v5zfg5I8NYo5e5pKUHum9Gkgi7Y/H4rhGZHwrMq2tlNxOdxnI2+ejmnjMq
HwCru+ZWQ6tpancgLIR3D5vW03/9vRJFn0I+J64dIcuL/tVLeq9ws6LOQ8UeQ5Ku
ZwNRfw7e9B8jDAxnQjf569qryqD6kCDAynQVgKMyU81dQETqUSt/4/7l7aQGFxTg
JczfgxO7jcvex8ybETiE/u+wy9zwmOef+Ji/GzUFxZJQ2IU09RiljvFeqb5CDXdI
ki45TwPstEzo5BwoBDJAZGFq2bUJKgf0ko2D5hZsbfKmP80QNZZscNZblb45Yp1l
iXdnIl46NsnrMcAl2L9IknpEXZThytZUNDj4lvwLRojXWtSxSj1oEpcXUBFPFa49
oPd3cGqvjRPou+PAZLzk2o0XLd713tT0HFO7ORA7JEz60+mtCnv8jyhLTwtATl5P
5KI5w84Qe19B6VhssxnkPUqT6lOG7ynCcSsLCUH0uc+gph4LHt6WVb0frfIUfx4P
zgVqUP0LWFDvgAT8gj+sQgCK2FpJeGy3yr3vos2fTiMnxvIdTVg2Vv1mipeoFoDQ
aj8OjlRePohwu1IFJQsbP0vM23G1Dh5VeEFPxReczR3Bx4Ry8nWckEq4i/jUdki+
q3LkaedE2Wr47u8Y2BBrYn5urlSoe8N38EdUIgkr25cOM+LKdS0tf3YTT9N1Q0Xa
75KPT2YjbPSeanHTrxQyPcujA0o6CdDW+3Jh1oYIlUyDpl6apGCsNbcmWew9LHjo
+SPVB0d5sRQ3h9hYAjWM/IWoV/di941296b3T8I3vLWZ3TC13HpcGJorNkpeRjrX
UJ/M9mq3eNikTKDjLF8pBJH8IUZ87Yk8BMPdXUsoi6F28E9cTG9aE6+yMGOETC2i
+B7xEWTLeQ1Sye4Zj9CRF45qFBF8vZMLXR5G21zZR908jPgJzRQO3fL62QHl24TN
SzOWDzhJBUja3kAb/tDX8HH42rdRznFY10CfWRpIYKysMr4J/19U+MljWinP+pUs
b2NVlIejNj3L17YUiHuFk3ZEJnTjILHUjtQmBXDijNBdE6kyzB8fOTtw5PlMmt25
mNK6qRBlwruwBP03ZBD4bPrwdFtWZIQlTLv4ZtCiGoVVjRl7FUD3QRzpvRC4ZR55
6E3YGxQbKoKiA3XsUWC7zcAbM6/6V2t4XNBqpbvp1z2IoxsOe8g0+pdCCrtsOn22
OLSNrSiuNs8kQTaqrg+hl0OFQdLf05jpWHwO9r+1oZYIRxwQmV0eZx3ltW2mkOMd
YV6fBX50fhGWkKUKg2ZuonDQYjSoqiAA+RSv2rlJN8/aSkQXGsWdjrKkxkFg1SB0
fXA3wrLlAS1fmfoyadg5jbJCyDw+Q7T6DfY2qkkSk9PGNQOMNX973BHe/8aulq+8
GeAHK0797HA016MK8KKCJJ7Up1zzWAZSQd9QhPE/1xuelyeCF+wCDYZzQPBjo2Mh
G6c1QPyPbIF+w8YLLADxQc5nAeDxYA55oXNQdXljX6UbnNwpHwrxY9mm2eQefjiS
gW5RC8Bae8/mjmt63e67lhBpVNyR+b4vDJIacDC0+Jbd8lG9FfjR6ibNMwB/rdxV
+ut7h6jq1J3RGyZgtQLArtpTAFn+BDoHnNSkiTGE+bkvnHlRh06u4V88X4l8kg0u
ArUofAx9rQZxMuD4NAjO867K4l3uphcBX7q8MC26HtL8e0An4rWG6YEzSVjT9xop
Zkt5RpzRhRJb3x/BPf3bQ/43JdY/VH6fpCiSIylM7bCdYVi0q1k9X2XHGj0ZRofI
0LlsycOj1HU5diG65pKqgs7tXS9pxpv0Hz5rwwciDZIFuDlBgfns/W9N2i2oPE0M
kcXClXz6cCEHRtGXu3+3STfKAiRWYoh1rF3hCCT/1mRIFvA0rhO7G/jrnMpkroBH
Mpo/zAR+bEVfdWVYux1fCi85KEIF6t4hQxFHpfNQRgnrR3PVJhqxaI742eZI4lKD
9pNCybGbf/OnEqdf/v9mTrlDfJr1KWu3zCMfhwktsG8Ep1BOK3BLZRBtg+Fel3vo
PvH2+EHv37anQPJIh4xkVm+9wPMZcXJKR8Ipu34VGWMVOTQfxSSqayma34Shq+kY
3LSzZWUt64e5HPb8tQ+k9+OtyxcPTTc3M0vXLiAmHL6JVqMdGLd+ORnEwLDxTSQA
lXDX4UrXCdRhhkCYQAMfGbiPJn5aMcCjc7hNEhGT0JeXOMVBTbiKDXjmWaumUbkQ
EkMaPgGR90Z/VxHNxkGWuJplHCOy/6dDNdnMtiWqfUPz/FH4Ft1heX1eQ5L9FOD2
V4toCNu1WiHu/FzVptM9TIfH9DhCkAG7ezHSNliq2dfjo3j4imcLqhqBGWWkxW70
ttk8+OrlCiGW44mzB2Ks9u0WlotY+O0W4byrsceDUhK1IyOdzRK283r0HZ4ak3M+
5k58OrP5Z1iQ5/ZOla98uEmhakKywvBGDxr1mDyKnoBHQKe7npDGzBaZtGxASkmT
8zdr/6GiA7uOZkbJR+bJ+lrhkvZKVvEA2YpC1WYfJcAPHrXpIQSDVo3nTlYR/Bpo
y14t1TT72I0N9Jq/Aio3hu+ylZBb/rwQPud2v/E/Hxr+JUIIEIovlbQFDBsQ9JZF
kYhoOtq0sDu5aybvfhBHRIkOBdb0d7GOboNhQTWkEWWBsDDF/jtqj5uBx+ONNF2K
y6yol1mhX0vRKcJb8OfrqUL75v2G6eV8RBkEhUUaxD7QscwlDhbTpcNiaQ9VQ6Qv
zdtNvIDzeeSQvGesEDQZV8SWe8nM6GJdtVK6iXJJnu9Tqd35EfR/cgFXRktu732w
j3mYoiHQoU6fof7SIIs7j9DBSV4qZyNgSQoaka9eLTBHV1M0GqqYI/iPyXNedbzM
0DS68wQqTRNClg0Ym5EurpY56a5RhU48LR52nSh8UMxvD2sEPmOgoAokK+BLnepp
6ohBWKBwFexag+k6fogD9vzDsq9qY1J1R1Vg5l5QEAM+yfuKoKpL7BZfYA2VaALq
h3Q9t8Bf43fXs7YFKOsCeGXnnJdvlQKSztNA3NtNW72OY963n6zQEwobqPPgfdeT
Bmv9l7toBVpEsoQbX80AF3/NBJCYDmceJ9FBcaM1mI4gXtJS//IgWdBsg7bMujjX
MztuqIjitrCs66oKhRnkIRCS5PbVSq3aqStcac8PJWRPsd/kOJj7MFAyimHYq5y6
gMGXHUbZOev41gXkHxOUsd1oj1HruY1skc/KiykO1eIz0p3kXmliOAYRx8urYi2f
PolZ2qxsZ2c34+mnlJx6Wx7ULlqGe/qN0yyu22VV3fsMvNYufi1xjdUYkQLsqMHp
L031tlp0V7AP8dVgeEK/flHolU6088NffKNXYx2BGQoeZ/7ipZ8/7+/SOxfA3YeW
pXtcjNHgVW/+033dJKfbqceycTpLQLMnTo47xlbNMs9I0qsmbwnfx3ZdIGs5w9OD
/UJFiQN32dEnRpDvgQMIhGNd8j2pu+yDzh5DsspalSreAXUrei+EvwCwPcjIAsff
easkSzcya4HDU9roGOw0TWQ/tdvsslRQh+j/sYefs86e69pVRQew0VUizwK1y8PY
DQzEQabtiI7uwi6PI5EvzWbyTRYjwcXxPF9imyrNufAph9RvNz5YL52HkuMIIaw0
6p+RBvmP7cDy5HYj6WZhCpTWeRxwcYccC5ILwj1X3Pr2FWWmjmUBjxugMAAo67XP
Qnoj0OcnBaFkBErqb2Y/PNQ5B+aroMUSJb8tTi2x9RlrnppvybBDuzbW6djrhXBH
vput7vdeXgOOA8+yLkUB4vYjcTidPDxvgVgXnN4hQo0v6QQdexMA2MLFI2kiW7vs
3RiLYxO0g8Q5Q3ZmP4z31MmBajotpsuvi90PXAU0eF174jaMmhlK7wl7vAV5A/8J
FJvU3XyWk1mIlTCuo824lgIwz9tATNRpZbYzhJ8wz9ms9Tg7AgYTN9A2CXpmi5XO
wdTgTezpJRZ8Xm5EFAoOp9KHMdLR4Qu+hL1fG7o0aoSUmet91xM2j/x8VvND9u+X
IXw6NZPkLnBLFnoghD9HtBmLQM6PQbdL7gczECoQkmDf0l4FYR+y4o38IwgkIufP
b0RRIlU49nvr8iW+qmGkk2eGtpfXbt0me1oEIj9PVDUMeGMVzAWMo29OFE9Q3gHG
4Vt2wPl55ZB+Vr/THlhYpXHrop9Sx3dB7KwZPmQ+84/msKSpznEsjrZgo42WqMJt
cgL84bDVQydvKquMwRuZTYGC53XA0hFOK4HlZWT91RDjyt2Fg78C1QyGX06WiyXM
N6l3Ee62qdJk+pkmBbEOTfcBSb02dD3SZP0EOe7I+G0hhexpzEOvb6Z1+it513rs
h8HQ2ifki0znAbHHOLghb4NL1PTiRYo/I5v3MyZ3FAnVIVtxo7K6bIq6Rz/rDegQ
43wXn+sz4XeNp4x6zmfYjZ0tTh1Af78MhIgzD4hMJ/1vQI0x6aTcZiaYFC1Ms5ic
8/v0ygFPh/pPFr12IdpgPiuFX6rSuxyY3uLvAI+hO3sp4Y8+wKIvrRPf4wkZSTOL
jLwCzIf3Ufe3ZBSBPhFNS/Gorp6rEHCGvb/gAdnjkKUOrA6+j9YCufWU/a5dZBoP
ohwfiA6w6kFz8s5wY14B9uZemj7/hqpbh1WWzKXn3/bYma0ORclF8qYVlsrbRbCV
yWQXe3gRimQQcjMdLjoOELxLaGy4Wx4M5rZ9wG7dvSsFfswvc+6D1vqe931csRZs
L6ApNh+4CvRlhsYLsEYnAOzxqrpWUFRIHpcZAVP0zEpjWCWMLsZqqQT7K5SFFFSZ
fSFYoc99wKc8ixrEbsFaYE8gDqOpBnwyyhfYCI8qOfu0QqY8cy8i8rX581D2c5Kg
TqFU7718heRto8DuvR0eOpN8bBxvj3ITM2lO/RLHijixAMx5eQzPCp/8t+Q+xE7n
Jvz/7DWBm30liwnSIlQ0kpzxu9WNJWsR9vZN/rSORmbkkxiN7gEOeT69WBat+swj
alYdrZpHy2mCg0Rf2G/q+TcQ/FLeXzZIIRVPKb/52JqRONfn6HTwHKN54jFh0pR/
XJOMixsTLGebNmC4A/UdKFtYU0QG9Zueh8pg5ns/WHQD8paTZ+TC5h6zjWdA3/qJ
oBGno4sEF4N/dAXr0xJZt+gvl4e2g0HW/YG2o8xwRaTVXwNgteRrnO8wq9wDcns1
EB5jq5Jtv+jAIpFkeSrpzYt02M9jx+nN0NBMnNzOGDfCx/IKF+N6eHS3dHcg0JUS
hVboX3cO0ZHvGyYI57avxNq2772ZQc165/ikJ5isPOvPQeNCWQl1B/4ap1VV9LIN
Sqi0eWsbZyeQF1ahPzXzBMr7s9R4MQxbalY7Z0GblJrT0vwU00/BUZaKj0Wcpu9t
7pGAe81asbKt6BHx5EektoRs3p1sYABGyyfH5zhUxzXvyefo/52Vb+dPsdnGmiXJ
NjD07yrze5mW3M1hYCub26GeMBM9XgKikkdsjnfxAQAZBfHQQ2iCxVo8qMCaxgW8
wLBDA/KT7oj8JgRCPwozOPfzE0P1ydf80cTneKe1u6NpKqi0uG8qFqwWa1ZErYeJ
Vqq2EViDQiorrQE83crIuqsoEv1rga+f8ZCJvQf2dsLRjE83uqG2076LtLcsF6jT
meVgSlyWRBAdjqEjYYqD9aVlNA8ipLJ1Bv4INb81zenvJlM9RzDWS3rFXi+UkE/7
VCzzD4ohS2q2ZFBJGFK5kEdSDIdbTAnUrBpoCxtpiQDBWAVYOj8Bt2wZNXyDZvY+
o9cSKIXu6LbFeoUWsQM6f79V+2A9+rq8TIPMVfSwPTc+9s1NsfChQwo6nrHnCji2
z64UrsV65GviLPt9oilrpBfqdECyNj9A9GJBesBmAjPrP+dF8wpAnbFcLkJmxUDi
GHW04G6BvZ6fv2IZFNrrg4Ma0AbUxwP76Xnkk44eAl0d7S4sjYTGn0obcmxWxQK9
jeP/IYkvyBnMGR6YM4oVlxPJXD4oyA560jcu7p9h1UXm2YF+GNk4utBd9wgMi48N
FV96/FMUZQVTNP0M4lwDWoELUMdDzR66zJY+es+Z783irWQixhgak1nN6SGnqulp
IT5KcTmSLlQTm5/dNW9n1XyIa7a79k2SQK246ylbrLnseeJ3SWh1Dg+lEvpDFq91
9ca3UDvFk6QzENO5SpFxv+IArMqTl0qHbw1N32P+cO8mV4/BQaEbydJ+TrAgZtRY
MeP0799dR00Bj3NYxovYfjl6FH8c2diw0gXcOQc7TRmreNp3Al/G9fBSbTwH8o+I
fH/yJQ17NNMgmbhwthdnG42RD4v+r0/BUV1CtsWi6jS23fM39p/wNeq/+cZfy6jP
lMH0WWoCQA2jlpXfg9oQtuouyRJGe5DLuE5mLXRqdzL7X/fmHMdJNiEevtxClOBU
Jj/bzUKRV9CvTR/CyhYN5b/+EAmoeAJpHBZDEpqmqw8ImjOw0Bo9FUe1YetdG3tH
dIvTWhv1sYjmbn40UPofpJboCNB7uoxGv+aT1xJlga7Q9Mmkzv8eJVfGY9QQaKtT
x3DxvHrpcspeieAkm65JMiuza65gfL0gRuGQ7FHF96TpXjroe63qQDZS163ZCsW1
cqrl+hf9evV7xRt6Bo+Jw8A57RF34jNS3S26Klk4cRIw1beCEL3n0VM41+6Rjy5t
ss8D7HhRWoKqHDQIaqCtnJhdSRstoT3dYyYAkuH8XfxkqGjNUK3YeucPr/2kEtQA
UjXj4VWIp4FFKNxkQJqLPqU6c2SwVWm0o7llXgFWtDwgD4m4QgpIQjTafD7Q7kjD
y7Yy1/tUNHxHPaWPgJYL+jA8QhUx7yrFSU/zWXOhIMXmeFHK+KZMsGoW8K3Nwc2P
aJXs26QyQ6K1leGqHsukf/hiAc6kHKMVC2l9xPcEyxzSUVNZMPJK+hOlVj2pZrPy
mNSCHFg6bGn+Inr8GbsKgGwX0g/v0dtIUJLT5huwd75OTUYA6o8sPuXbS/iNxuRG
gN1ybMaQSxVzLb6A+xSB6pPDD0k7xjTT0KNKR6yiCr3U/uqcdqLZSb9mnk8h9L25
ktbQdweig1l2uNINDwV315Sgh1ywBdyWsMBbEFX0RB8ZO1q2EyCuQeCmCUf14JUn
qY4B1pYyeyhIV0I5Cb8Hfgb8LCNeVH/y1x2dlY0t/yeZsDCX0Itwc+Rvs8gTOzGO
z/5dS4E8ncI771MXiu2NVzP6Pf2b5Zco3U4Q66IWpg926LnEnONRoyJbHX5kAAoJ
0c7VT0C6p9s55/fSbeMchh4/ufDKu9qK3KKQz+co2Y/wIw1vqcrDa/n1wuC6/GoL
dIeJakymOCAh3Us19ZytDusnlmrfIuEbQSnqsZfA0MXQ0ch7ZBSFKxRNxvMPsg2W
2PQGQGOBK2rBgBjdSrIRvXcBtsXsK70rZE16HxOshYxMV+PfmNUJqv/d4yYjRWZA
cgnJ/yz+4fXf73mwHbwUuNcRH4Tq1lzHQ39YXrNLAzMDjahqcK0bI+RIBECSwkOn
YHD33p5GJhXKZ4QfQhqerP/mGTLY/HYC8RoXBbcNQic2u6xh6aVefpItDRlFP7yL
dh4oN0dG0mJvyLO/YGpEQkwOXTutaWpfU54wCoUaPnxzVnk78qOFcFdQIzeTxh4F
8/FQIxCoQOnYPdsk+gO8XQl/CByCwPdIEWBg02qpN4zRRHwtxqcmLgTluxSSwhCv
sthGMZYhvey7JrrlP7SFGWKSJ07RI0X0RcKEW+nWIGzDH5okT9W1gfvYwoRzY9Va
yNvh9OLg7EPHF04HNxhI1AGKpBOuZ4/swqo3UjVGQF3rffKURgnGhYWsu9I/0ud4
5BTmYZ87oUdBdWYxyxWNhV291kimp4+vXbDN75OUzjJWMlRcYniBfkfLKm4Z0UhF
u+giKGrbSfjpNWkUNKFtdjy+JAMX9FVBkGti9p+weKhkG20PQPy3aPdrw29CVabU
RW40OXmh9qNfsJsSTKs6iFuT0L7NNMd8Fts09m366b5T/TGdS0agZInsQcvyUL4l
HEjyvbHlw/EdFGAxVFTL8tBsbkqI3CNVrWxKg2cUQ+GuNvUCaomSLxVxoVuRsTds
Tg38EIujLX6NtTuE4m5syge6/LDT7+1jx4eLpV2d2+fZfFcgkNFcO44GPGalumeT
aqvmXO/xrHA4S4jGlvkuNWyMgsAhpR5yWh/lGmklNQSNOtC5EWmhEWsfjUR2kov8
vP+EB6BDUCl/fmFGLTTiXT4WGNtKYL7sPYaSKcHAcw2yWgrDh4x/Ki9vU2weIupV
qu8H7oBW1Kt1fmma/blgyOy3uo3cFAjoZM4ejfsz2PDV5RuoTbFtfgenjvewxBjw
szO6AVMnSyj8dm2EQRutOvtbJBioUf/l/X5vsH+gsIlxkcpP4RZ/6wo3xBD3pbUC
3F+KbigARhI4BS6wZWyI5aH7XXYPD4CB3Y6VO+Nu/Pyv+j6twdBTGjdKAWV3h9Ka
aez0SBWm6/qzdG6GRLHzNBUr16pPTXiiik8uNPASdoUuzBbLKBG0j8RK4ddZhC9+
jfXrm1S/UHEhV+u+oHQavzfuZD7P0fTRV8Ky0yL2vmp/j7gCJlEdDxxIsxFxXKrO
A2er13u3cv2FFT0f+n5xQZz4wIIJ5jAGL7Edl0BRUZwRz/J9gv3GIkE70C+FG484
jpnluhcAMYru3g+CMSqcxqgLZvPbLAoVSHxj01ajg4qVKhA9KgktP4CyyLn4uUSv
sqf5yYF4rEEeo9vyJMf2KJNLdQxYLy+OTqfXNLIEY8qa7YRrPKCS3NRCUCXRySmj
PBxR/eDL+mhWR3bpctkFojNCKSoSrXswTzVumcQ+hA8ld0P0K2rlKGjYF+OUrcgp
6XIaILq0bIGH2M7wK7pUbHgx0kfhwoD/Kcp2PEB2aBmPgUbhQc5pfqbdAgWcyT6c
tCJbPo1PHBe0y/0BCYK5aHQTIJ5oI+vC/kPTYKcVS54/wwsxExHnuOawV/mrf/7G
ZinRIGUdcO5TC4Bmx93ETRjgIdGIrmstLW5C0damqYPVzx/p1EvtwUTKvD4KIyVL
7aT0U/W9711NGDhwIFBYH+8Dy4VJslYKAD5mhfguV8wT7BrJFvW9hzEF7aazkNW9
RPOAzo+wDHYAcsw3fJJHnmZCdhfyEVeGz/t65OnHPTJ/EBz+EK2RpZzF4WvppGht
hhve3nTtdjuWF+HsXPp8tct24WP5jrwhrkhvb42u/Kz59eJtlHy1IrWUSx10mhY+
S/c1TqVl6ebsrasWjzY9VhucHTHpMY6UypH5N3PIFg2pp7SyLiYFbWNKgWo+GASC
7alLAqLuJeZPFVyoRBnO+T+AsNjHGZ9Cbm+7XrAXEiNxq9m3CkzqKGJmI3j7JLvx
NR/IqhJRhQ1zi4hL/x9iCfgtVCDOwy4IJuIpwtYWuwbA5f12QhwYffk1vaZdqhBf
GEfbGmmd1nHBfUCwOjveaibzKruzTvY48xcD7HAJQphXVvzJpsv8uVeb3WogOLHG
ldwpiGOA0uXJiJTDlIxSLL23DF1WaG/US9qoA9NAVUf/gZT/5hzFF1efCjr4K2xT
5bjx1xP7uga4aiDG9glLnqTCjRU4kqaFfAxRFLnCXtcLLsEa0JJEGztwO21lWpUn
79css5gy7/OLSWs+s2ePBFiJrtFK0/orcZHvzj2BBFXNnrVPpm4RphQk+9x/W1/V
RNemz/eqp1Gm16K53NG56C53pzf1vDXgNwpDltJcFb9R0A8vz1qd3/MSLFcpO8Rx
sCWK9/UXJqdXu80sukZsi1JMiXDZUQkpIoyUcTWvMkGNRWu+AhgKbRigwc+BNonL
ueajVT/AjZNrXWc59/IU6V8N+uE6pQiKbobm+CfWwggwwHqZ23BulTI2CLNt6vVV
npiZc6hBi0i/i3Ze7U4tlsL4ODAiGSw1yUbz2Kkj7XRM106SMO/Kktb5Tfg9fdLI
0DkaDLbDsRdl8NH+9AbMCnC2MNzeX1zwQtyj6QEJ2TfJc0M25+SHRoprj7jqx52L
FhUeE95CrGHkJOrZF3yeFlmLD1f5qxwaAW8J6WLVUxw52OgsF4VixUDHn/VPlXba
04Gl3qj4yg+70YjwHxUc/SeZze0axpUgei5HGYD935hBpocGRpavBLhMm3nW6oYX
lFPRKCMzWxrUFAagkRLdCo0EoDwo88dhyeEqkZD7hTz7lHb3+uUSXmRj04RwNYo1
1fkeRtIPMAzJQhT4e/HhuWRD120JdLOu+cGaiTDfly5kBAAG7pd9tIFqp6TtB1xi
2QiIfI4UWgN+DQzK3n0110jtqgE5V2bXUOr3tPDQfp/2dUTOZ5Tpg62DxZQRmawV
h88fIUN0Qy1jx69FqXjpUvUk6fSEiymLcj535eVZbkP9zPhsHf/3tvCr6MmlUf7D
3SzV2VUXyYqGF/GwunEMorwo1U76YhkreccmchMmHjcZsrsTHoerQydDocgXJpDs
Mc6zqGXgMU1WD7o8X7qMOTkjfAL1utKkelohcxTbH+qY62kE8XWfLwNpIkC+6BRk
6JullKZ8rCRfYvaCi03ip3ivoU+nEf/0ZgPDN02NM3sBciE2ARhmgXHkrKJ8GJqV
eQVzUyaA4PSbwhKvRN5ekpxfb8Yk1GNPrtMrC+VdxdtFySLHhuFfFqkX9BH8+auu
zLQKYUJchEGlOlR2bu6UdR5D1UVyFpEJRCky+zVAoD9YGVEbLngN1lkAPj/ALmKg
ao0eeGoPxqF62htizJg0y50EgB0Ca4LG1JoY3TgiAzR6crVew3QhMiSZQPEvUoGv
JDlE2lcq3mj+k1kB+sQ+77SvWocWQq6Rc05+mvsscj5AaVgEAoh0M3Zo+74bBL6c
rVvQryAHdHii5JV7SiTEn1rHr88wTQVg9jtCOXDrEIxbe1qGV/Vjc4CtHFNVEivj
QboUh0ICEBdRYlV/hkyfVqcOJvLq7s5KIhoXobPiaqpqWPQQB+zRMU+cgqsj7ZBt
MgXRW6Xj37Hgy+NCVZF+MVs2BdXDEEwKy/vTD+kTklYMMFaQqiT4+kdIwNUFoUu6
ujeryFth24V2Q9g+LupVS/gyMVf7zwGnzksIetTOCwcJcu3HQXqSsHvv4WcderF1
EqPvt1M6WdyePGoMNpt70ojeGnYGQiREceRZ+acQrwMdRUjUm8//ieD+aPuF4nGJ
Jrf2Gr9+WseGJdwnn76NXFhyGbm9uf3FxvzEsDxei8FF8+vbcSQUgJRwSSrets4/
Q96CnKMObF0t9NHHtyIHOGeFcIvez3eGxiiAzdrlbuqvhsRlTZLw6AoHUzgW7wY3
Z+ypKXjdD5DuOlu7xZDWvophFdqD3ttZKIyH8QtVfcXTCltUt6LGmI1JclSLJqGI
Qe5b6bPK++qj/RGGmr22+x8X3tIlYK5dSoclUgbmCspS7Pd6m2ORbdwhm5MSzgLs
6V825+sNOWE7xyOMLhtjlwvrscUzR07HmBvhxd0XFe8Je6M2dtBhrwvNiah+YxEp
bKPqIv2Fo51Hul8RZFuirpTH15PudmcaveSriELN4+KClPYIv+wyBINbQ8PSngiv
jL38cEODWq3FQL6ypAlx8zXMJdab3AEkDmbUqgBH/jplJPE2yrBy/AkzAcJhKsrd
FgqB5kCinrtwF4sVUUFyFBqvTAM3iBBhDx7PQ6jAUkCovA9vhG+3EaRqvfO13NfO
wp2gzG6e/EfrhsBtLONGLxqhojUCi8WLPi/k371ePcn7Q7iS+jPv9AQt2BO5z4nL
XtlS3Ly9w8op+aLSOIFAnoffLauTsFyAHqnRD42shsp610vv1EZqRrY0c9dYtYq5
f8W+UTW1Os78qc4ANklO9fSlsxX7KZx1Y9a7vw9sg8HNDtm36QI1V+CAjrUFYFWf
rkOXivsxVfk7Lwslr2RYMrewBjcO3ZcMjPh/lQfiz0mGP4XgQh0gNvsymHk6KqvE
ZJDzYj32O1oBgcu3acHl+X7snbU5FJ25RqF7MtCAjEoGTCxI5W2Y6XcUbpvmMOZJ
9UXew29DNvIJO3pxsxDxO2+8Vd3Ji7yqYzwg7dmyKDtKQ4d6AWB3Z4HSrqD+XcHk
BHM03SFgAQpiJMSgmtU0p3yRdHqLsx+XDVu5UxugjwIIaZk8UuwsemT3G3qcnp4T
2no78SUYPoBGdg9oYaTIjAuQhBpAtSn3qi5OYWH0QzrvDZrAJeQzR8OdF1YUa1YB
He4KtnDUy18/viPV7XcaI3ATAgTCEAbLtkIQ4zJWArvAoumuhZ/4FOcWIgrDvgZd
7OrfNqSnjLVNlpp7kBMZ44rWHmQGpiNmTQvlEg3JhSLgWJ6+7Q6gaCga+5KlaHNF
GeJsKF34umFKtSXpT2NczN7VimADUFdq/pgSGZsSoYxqHLsO5WfDoOn+YbmvwM1V
nMsl4Pi7DPWLeGvaug42JSUjKH61HADO/t+VzI2daGHd1nH2JIOyWtz7gdd1XKCD
YSwTbi1NugCoRi+QitIJ9OWsILVMDDGJf55pKGhRttIFl+k2CRD9azLBTeoJW9TQ
4lhiPune5Cwru7cBkvJTQqF7xXHl4rLeLN2t19SVbc5zntYhryhVa8Cq7+uloFSP
GnbBH2tIul1le2DVx228D5LhzfRc/5RdY5qXMt1An1ikINRjI9buSJa6RFbCgmPC
mLq2+qEL2x+YZOIHyfwPg7tuF/KW2fnQ2P/qQwbKGRJsi8Dg6Aib2MkKvd4fXYzG
MU3BRG+Vrf/QxCH7q/Opw9QGbaWXWjD/Bc1amqcHAX+mgwnfRioQROC+c+X/qTq5
nQ1O/r1Kny6Ulq8X91GAjlIccmRn4NhgvLBfHFBO7c7vSepBnhRmFyMOcTRp+i8I
GdFKPfIoy8z1akhBmB7tasM7CZiRp+0gtRRxVmknFffOumpxPQ0nGydsyLT1g+Gl
R4rYQ7m9WXGaqbaTWPXzObGCWtB1SWSl/kuMEhhpFX/LO2zg84KxbLI99/e+Uqgx
AXeVeTd+Tyw5AwptLxNr06uKUAr5/UKgdk/g95YIr7OPvXnhoVy3/JVcmRzQpIQ4
qRjtkeTAGUC62ceWz8yJYfgB0jXXNV7l3uWdmEyj17t7dHus8A6xaw+/k9nHzhsH
6x088AYsmvBQaS0OyY4nGVx/pOI8TPOSMdObtf/QIUtDPFklXFSqX9nGw3VwRdfg
YxWqSRa1Iao6/QiQkvxqGdScGM3vjHvfeAnBfMbg2TO25XEVkDYz3KkTc5a8JDQ5
dfqQfepj2ra1LsI8XfXT1OmBDlCZAYKWge1SsafbZY8Nnv9aB+xjZGvcE+y2tglC
swykoqWsX81tA7drgaEr9jQ5m25Ja32VAcaVNBYgcWUywe5aKQLfnRLiStkmgTbu
G1DHqVVwYDPY/ei2f7xW3nl5VjMgwkWZLRXEk/1riboTOfvhIzBA+cW3ZRST2hQS
/3SI8EHb5pbKUsMHFH9fPzK4uquGQl7iHwKa5Y+3PyRsij+zILQwNG5MDSeGze3A
vufiSA03X9Mwe1yXsqJWoFmZDsjxT1MDl8AEISc2gXFoyYu4DDyaYMH6q1pfHvH2
TVpMa8zThAPG4PqFm4mAJSjnB3S5L0G3Ha5WTZhdCUodHmAPfl58wqmqBwq4QmPE
3yr31GbTBnvrP4ZvXUHXnqdo3U/sJ3qtm4Wn1deYpXBvsENdtUIME7Kd82URrtS9
owYutE4xlDnPzuHZZKdkLo0NoKx7eSyREvoAE2zzW2W5dJVgHBBOg7ZhJhuANph9
zqPwUcFzQ2i8Ed4NX3BJMVRv+p05V+0ISWqD42fNmDnOkIAoRX6/2Xj60c5GR+zF
Xx0ka7PWsGZRCqSNiwyi29U87giwYo69iW8+eZJUOXvJn+z5Pv2vdLIKub0P/HAq
mt5zcADm123mRk44p8RLdD1UQ9lCG5dn2Lt9VVsWGfLnLmM3o2ZGGVlcPAbl8YnM
Rf/Bjdu2CPw1eZ7DXnq2nBl3et/YHULI/RtpiFEws/mnGefkS6/ydpcMov5ltGXN
9WuBPxALfKJoTQzkji+h9zz0lSeFf6/L3VFPj++NBz/zexOZ+pkSC3EShaIoezvd
PI8YzfISa/U/+6xjpHhGT6rwpH9/NX9/+UrI+NH5Bd5HwJ6g5LyojLIn5DmD37LC
OVE0Vi4AArGXXLZG23QsPy6Hcnk/Zq4xMhZSAfGfWqmskezfbO88S5QV6Z1wvENk
WshcVTVh2ZONWnc/aYQDWaUq6t0Ajled38eR9PzitN/dlthJi7wveCFS+JB0sKCX
UgDa2sCKahCiceWGRIuUKNd5tf+Y5RMtfqNzdAQ9epeT4hrA0wKtcflh691G7tu/
Xgx8h0QWou+OyEWwrq70HGBq1mnRtpbDwWxeFJ5vnRyaTsKcRX69v/tv7LcznpmV
lgmwrC6rygA2X3YzMqZqssoQZMXu9i58JNyCA+uCfQgtPtGe3ouUgbVeeUGSjpPs
a35JyUKWjci3lsJUY9XCtEc/xjiZajYzde8mhmoWlCSemP1mEKVVdn8h1UY0FVci
WFRu1nnQddyXNHBRdYcK6rICk4x3QDf4EvOjxSkS/bKJNpiLgVQq+PGsx4mAnIBN
/AGoxlQ8I7eT+ekP7ZWhN7SyR9VbApOoJZg6kgohj5IZWZhHwkxgJhOpoDkHTzhJ
g1Ev5KruRcoZWppshm8Q1hhSHYW86+sqIsi1hqYdvTj0sii/PNGWKTncDWlIe6KX
P9+jjGezdr++GdLnqgpvRUbHGR6gEbkJvoiW1uW4O+X9FifYAx/7YusPcWMKj3hP
guvMwQvd+KWRc8lCP63ZPjJZpyOYPSE12wpg8QpZMCYlpdShJiMcHCZEszenjwCz
aC++AWVxW84bZW3k0se20ZslIu7y85OJ3jhNoRgTCoSDXNNaTeYJVQT4B1lqGxyS
lTuM75HTw2R7+QrD75RSGcFQfbMrRp8Ha4yReUU/HuA/8XWP7n93oMVSi5vxhRxv
lX6AMN7OkOLj9HC9Aftqb0hpCwT+ukFev+PMqmkxd2e8Iysai4zp3dHlXRbtPQDz
DfmrJqGIDhmZh+PPAf9u79qey/jtV29sueezFaZtWh3BMWfiBNbKc7evGdPE2zb2
eFJQOccSNoGc4rFnwtrOkdo324jl0mpyZFDsRciv+f6tmcZLHFyZ3mbxG8lWvyMI
ZKjjOpdYi2w1eY0e3azRgeujKwPKgQxZlJ0/GyjHtOlS6sjokDQww59OJ/PR0jqB
v0GU4JEybjbRzLjmSAN5/iXMfnmb8Rr4Kbm2658XQOLCbBix+JEipdtFQHzi/nkW
3fX4bW+dHwM19s9mbj4gM++GDanNolMreAnLOCfOp2tNo20NSYUncmxFztftsY1p
0HOZ39/ZtxaTy8l1OChwrW00FoI2re+iMc6o4STMKpHLJRVZ8SI+9HunAmpKLJZw
NFo87MB8gyhEsnWIDxVctTkAa1ky/3d6rKSZ6UhJypXI61wh9d4LIxb1H0hGCMHi
o0kAcStaOSJCtrVviprrj5NUvng/b7NSG1umcTL4m5KCxOY4k+kHaoT9YPuSxnfv
uwCtEwpJY5bq6K7f7joymNlJG4doyr9NnHdnlcSmjegJECnhlKNvtTxh+zCRal9/
TmGJQLaOMAvOOjfU7M34HxODmevAjwggl+irQxkSq3EFUWZ5whO7rDGENUpPbl1F
CeQq0Zq3siC+/PFnwRuPZ2CPC0U6kUoJWcrUwE5nivyF/2xYFvvzAdEEGCgoMgHj
oD7XgdOS44Qh2zRurIx75Z6Sl+/I6i/ZyAZtwYCzgGxBxi7geNakLne0RVmY196y
cKVH/M9OyR0K6RvV0O179mvFZ8yALVioUt5Yc6WTQVlRAsc88VsIPlHG95gJS6y9
N+GKTN1mW9m/hxxiffQioRg8W5nW+Tvq27h96MZFaT2QzhYUWuySbI/xZU7I8X/X
WMFEYASu/v9yghgPAks/OIVTo8JvWb1+YHkpkt6wQ9w0aa8e6nOfWf0tuNIrr4lo
k1g/ykNKA4IIpzlUrRM2sRz6Tj2zoHdtYnWFhoLCNG7d7102dZ3KsWj2q4rZswBQ
Evk5DWD7N0bA3AIZCYBwf2V7ekRTc7+af8UerJI6vz6dXDmTqLcrCrxtv3KASZoq
47gYTo+AdKv3igbjnmViOGO8DncOELqnhlb0k5kkJA2jswcziI/x+t4XC11KD/yj
BVr1S3BGdIzUOMt8f3ISznKX8lhR1EMShCF1+LTVWuyr3dzLCPS4jx+Kdlg18Hg2
OK6RIeKY/VrXosvYhVqOYuwJ6IAVzOBlDyjErnd/LLfO1pG81W8EVLJMrf5BOSHK
ME8RYJbVAyEwkEwH+TcivEu3tttreB0e70S6o8JHNc4ZGKjy2eOZ/mDRo+vuJPjN
fBn2mdEZmDGI/eZRQ2+qTtxEPRo0AjlbMmgvVnND/doOFvPTLUxgi08DpD2sT0+x
5mxekt5Lmz6HaJHt52Yftn/b7Ft7W91vlrsCMw2rNLMPT9vllNu4+4xsZWZI07lj
5MeMagdEwcpegRcTYIilL9kKNYg7IZP6JnRsltMgKfDDQYwt3+rTct5RyHGK2st9
dbuFxAbjUjSIOyZ6aVEzOg6EZslBfHxgx7HtkQKczoL1QjxY6/f+mxelC3EC9TZ9
HZCDOsYUxEapv4G2Tx/pvQ4V6KveBLlyOlewtiFNYljTgXwtHRab67qUdrST/WA1
Cxq5ico0tgWZmNdwKRFPb7wcqBFPG7ed1PA6yDuoS5JmIsd2C9bs09N91w1BLgkQ
c6wyDiIvs+RibWnr4iaDTZFtzQDtBEJwrRk0oRk05304B35mdhspJxkp4HgFzp+r
jKFLSh3xdfQbFCSXSVs1jdmCfO48c+HJmgjQviBMt890pPe7D2q54jCFOFsAjAGL
17ZYAywG/cvqE4MgKAq5LI5mcAGkef6C62XsmLYx9ubiYH1MO+hcgb6sbMebGJH4
VOY6FPot2FDEnfFBRr8HoGDpq7aaab8arBlGOkn5pp8DoyClQD47joqMNaEDFhLm
kqwtX2gZ7JCWnN0iptvDKRVr0eQMs4xQordV0rO25jc4xULhGB1zWYwtKuQsVYD3
IF69+YpKLMTHhyD6Zrjfcwt09QGcYllmFZmUqys6P2upZTgPZ+UXCy1TBNVJtRE1
Cwbu6gEnSMd7723A+UwRIgWkwkslfX2qD9TWm0tbsD+OtQtsfD1BeErPVrhrWOkq
MbGA0WVKHoyOVUGnI7IXQPnhrb+kWByppT8FenjkZ2L7cTHkokB21FTBwt05V8Cv
n9TXAfo4kVqnkaVgRklWjq+AaSaNJUP95N3K9rBA15HPHZLpgR6tJO1hR6bP+rr9
Ay77kF51kLtDl0nCbg5fHOoi3pIPgxB+V0Y0znzv6QGkFJIuGKOSJU8/niBUgxa8
n5fAo9zJ1VUBYjSwaFAngADhn6YICfGBXbItiX0lCrp83+2O1ymayernUeFOAkPk
/hejEjaYa/hyvKgIRuCXFCXIG/VjaCKLGHk8zLP3BoqXNdgDrIClR5bgx8dVEJIC
i1LzTB41xdpmK+9IgrJp5R86/IMutnTIVcCCq3/hjXx6VkqXGkOot45urniGACUU
tLTUch0T77wkAszqjjYfluH4dysvx8rOqfuJBg1ODfKPxmWh4zx3JjZe2gNOKtgP
+A02ZhauFHQ2u6excd4kgSm6G99WNA5vct7CrxmmXfGn2XkYB1acD6/deI2+FlHL
IZ7iHXhv20TD+IzBKk2mh7cy8s3BL16WKxAwg+NaVWwAHuTgoeHYuCWDfBcgV3sQ
My3O085nbLODvUehplil/t5GqbEDQEmKzahyOSMLSGk0A4SL0nlN99/erUa5Cq+s
U4dyEt2rO5QSFpiA/bez66R7/QecDYb9MiEuZobap87u2zTzw/CHsWGcaSi3BZov
uMKL0wpQEIXBQGSRWCR+EIbixi4nMlhOZva8tsbDAPXh/3DO8aIq1yiHH/DR49O9
Q88sgmK9fAfR0qE2ct/NfbbUJLiYrWzLDrlu4Jc4oC8Hw2eSQmIc+nQBEFStRKRW
8FR11eQ6rchCatLmM4q1cObg9wkGds7k/g0vXSNxNZiuzIMeC2YikP8TpHeMGMQt
2ns2qbTD84J4D2TUwpPc4ya1VpsJT/rcdh4NR/xo+S4kmWS0hmJTTv4u+eGzxEJ0
uTezuDpWZ7qzpKI3j6J5+RgE+3GaE00PYvYXA7zidHO+8wTnbnPuehUNbn9mcDCy
KK/fa00m9OpEB62q6klkj5Jic7Brk7emkfqSsJxh3/8ZtPOytfu2FvasXObAso+d
NVxi9zd7TWJd5Awe87hzg1AlnICc8RC66ibLfnq3XtYKBqaZ/aw0lVSGoN/VRSCZ
K8bya14PNTQnp/m4NLeAHNa+EyILCR1ab2lAKy0FX5WDomix20uanorwFWOK838V
+erQy6wnCvkBpOnWccI+0m5z4kOWtQ4stYuYM0Gu3tEDOQiluZ4M16zrZBBhEznh
999WIuiVIvvNXt2hGP6C0GRoKoGlsDZAdK2x305iB5An9W/PszryHeOSloAcldlz
1lJqEz/aG1EepNOPli4EoeZrNbzylM4dXZV0QrCGwd2zd282cJqqfp+F3wJyDQKF
hAkPCLYO/FzbEXi8r0S1cnSh1hnl5jZt99ctW9Mb68IplumjHjbRBhyZ0tSlK4Qd
Uitgr55++Wd0O+T68SYwfm/Www2i9ckAIcQnoRZ36Mq5DkPbPoO2Ic9ZrgHRQt8N
ewmvVgQD32kl27VmUVUJcAVLzcX47fJj6J+moWGfEHTFnZfgDHbJCLqDz5Z2p17G
gEk897VLj6ImlYNzcxkuqKqwROQ8Y7HhJo4wqr+542/0/SI2szSTEyUj3SF6N0Bs
53Cu04h1I8VRkVmcfgOM71xkk785Uoxks8S6IkaVM/tw34POouUzNEXtXVgqPdT0
hQlXoRx9I7s/+oqWymhojX2eXLLRz07rQGM9B7xwdueRFHenzNjmAKb5+OUa4VNW
vz0IjTgaomFNCbdg6Z5GUtDi1+HXTYM/EexT3XvmiKZMCAscm5C6wM1qfooPXZVE
qIAoattgHjLik2SVffG3Xk5J7egLvkJ63sevHy8p3uzuAPR1kPqPjv5/D6h+SMQP
0TDsfllokyIu0/URu7JqEUrzjQ53QBZ1at1Hy6wzj9A7kYpQ3GNospFeuzxRxOR9
4vzXfUM7HKfl7icKnCzYwgLa2rgE3jgciuYPvt9Y3C9y60AJ4ilwY8+NkmxgMQY7
V/zxBGuht3ugDbpN08Vnx8G6DHPHNKZfm/Bg1Cbv+Q/aZtBIIjIGxgZOItouc1ne
JGxv8u6KG7vxU2FHBt5sxLOm9s9D4/5L5fBTjSIch1qHqR4EzI/Cge5zpsENbOR3
pS783k+PdVcnb9mK7yIc+iaFxJtuTjd4T5MCIYrq7qZT4OoI3GEC6tFRFISiJz2W
zRA89//jUrsAWXz7zoYROEDIe+rijM70j6NLLmGLQnC51paKnXFcUinruvTo7nWO
7WLPZw1KoMcU4WRVa0JTGVaJDM5Alx/Ee9yOG6x00XkbRZHS7Wl0D8Tr9sRpA0gI
0GQUqyARmtd5LULPeHvSZpqkzRNYv5rtO8ylFFNq+zq2iFjU8e4aAI8UYZKvPREs
+GfMFahxZF6Och2iGQ5OEqNrKTCoWxxKqBGjqbtdTDSrfLNm2NXisXBAvRHer20O
3GDlfauC3fKqwPdfSWRlcBQAl4Rpxd70M7ak4cSozEUces1RCBEFvyBRT6GtRNHD
VUDDrztqscnrMAqM47wLSkfGyfXHuBfdKWm/dTD13/lgEUv95Ajl3BSXwch3A7HF
EIpcN4/u8G39nhYmBTYoAGcn8Z68PsWJ3+083CE0LpxHmON1lZk3dn6Vl8Y6yxCd
7UFLP2SDgL29Rkcud/WwS6brG0tu1AV0tHe8sFGiumpoSx5HsXBqBR6vrZWMKSVP
VU3AlDJiUeuK9AZ3qVzAYIWKiIoSuWZqCniN33Y7fbb1KrneCsIYgNUyS4IIAaPh
HViyABvu34VsYvMmwOAwcvLWc0qM6pQF3iT2JNLYdQBNspoxKBZMb15x9Evu0DVd
dVj25fNRAEa+bRgmvtgwcY/c3oXfHNcl9Yv0ept5HTtROKZklqtwCGV8dFzlD4sg
Cc626o1aWSSG0kRMIkRMQvfRCInFj1ibl/eL0vKoh9DJ7L7L93KOaBy4/spJvhZ1
o5FMB6WdyKcBIBzbZ+Fqj8ySU9dlm9ufoPCGgpeHaty7ZU5sUkR8OSsTNI0m+Mcz
2G3M+8tNssQ/s0vj7g/BmGe5uH5CIu0s2FHZbuuYY0XCqfTaMSJqwkhOy5gzJNoA
dhEzVzEQ0CdZy88zm9vbMJmByYk70g/maGT/1Rj+dhBQLnAi+thOacz1ngbLdwg3
O9Snt6s5AdoGO92N0SOpnc8TpNfhMkQfVNac4U4D+qxNkIOURf8U4jHlstxXCXVz
OSyFB129PjAAfuinv1Ao69RzQ6z/pvH2k9tjCC63RoIRkEmhuQq9nyuObVojHs4L
smSHZCIAjCknX8sgj8A4OSUFrcNXrqDlzEDhhPDRAf/nIq+j5BHHCUbv+ithLrsD
7XmhfCWa61AkD8a4z1VWG8mZR9Zj1Z/xkC8nuGbRTcopH/2DtK5aMiY67JiCUnYv
PDR54DfpOulGTqOQeD3l7krcni9xm1E5T/snhaO+zyzHKKxDrfGvzo0/q3xPWsxS
fvtd/qhjeL25cjqKg137g8K8R5LubqFQK2Kd0vvEKUoxK8nmSdT5CSuGb95cWdFx
zLfMjXnggGV9ls+5RZdD9BjEXr0hNqlojuKWssP5Wg7SEJok/SVweQtxFHNrVw3l
sUeiDhJPn8i1GEaT4TPmoAlPfA+SLpjAozklXsloRPlfo6HYdt+eErk1c+BPbJZ0
XpTGi3N11Fv3u7WEoz6Kt+EjFBnCfzcdTNFfnVf7YCICDrFDMeZzDn9tAuMODoJg
ZNUzBfS3zaCvq0d5hMgUpVMHB9T1+u/WTSvTzIMCH2MjxZtfPHUxRBt03xcx0SaN
pyFpcy0hdV3v330ZdAlc/M3p8xmrtb8S5P7QX0BJnLXYJkOTphgiwdnpKDqjEje/
bMdDpUY3o8ul0NcgUdd8e4sIGZ+CrBVl9Y9sVdj4ydJP+Xk4IUU0RN6oGadEA0zt
dmTlT0luG2M21q2Su/HQ5yB7e8ypa+a46ABRBGVvUoWFM9DUJoEgg5vPjh+XZerw
10BS1NblmV+m4QEDVHuVmI/BDhl2ih7uqieQZcmf2dgec51IQglvrdALZdgnaq5e
5hGKNo3ztKzpn2Athqlu3+VqFn1oUxtWQjqMURjgw3aSRmQ35DAKTGaVzbg3Di7w
Q2TO3gpWIStL9gmxYFSmYcOxtZodT45B1JKVq5qPdSfF7tglAmQyh8KkO9lQPWJg
35JY+UFmNF0gsDGncMahPlaYmUFq/a7FSyTOtco4udYTdp4MyC2cRnEGo/OkoaWu
H8du3FeBkoNV/TLxvG/Bmrk9C3cO4OlvflICuR0oWXixbYEdIKFAvZ9fv4DKkT0I
4l4U6GEYf9+OrCze5yjQddT5VdjL0mUK4KNJr5SVJjeKeu9DFJH4j3BPkz1tmL8f
bpQPZ285HdD9LsHX2ge9Mk8mjbqB9XKAXdW+VWonXJoWVWZkID61TV9tb7Jzzu2u
HkqIZwVoTOpUoKd0u62HsghFc/6FIx8N2gPuwDyEeLQYxRggRlbBmNj3LQ4AudiX
oI4owhzfKTyXpHJasOEB0aiWKNViSLaIxawOjniuuja66eQ0UblbySM5Jvad2Jjf
slcEFh8irjh8DJgHyM3XJ+fd0PXR+pJGNYERKFIcwz9Ir/jT6dYqSZjqbMqOIZb6
hzJSM97bsOtJH4kdHs3+lb5zmCRfDpIcmgc6YEiU9uLjMRe1eIv0cc+4baibSgGE
8LP0LpMoUD83ifgS76yYQzpgoRbR4yeT+BQXc39G4Zeyiq6rIDtvUxMTCEXCWE4x
WgYgfN/WND2xv7DzaPTkw6Oy4Iy1cWyAHtnq6ZRKBB5x6xRujY/sdQpyiSbUH7ZB
rIKapDKL1dexnfWkGW5zOrH18xwejmZ0uTZlj5f8dwwEUy9kEuSTMvMOJL9Pt0c5
OGdUEnV8V8MHKukUtA4Z/FoYJMZ+0NfFzwZbVzHHLQOSPlPnexqDGa+sx0kA7uiL
2HCJYoRzZe0JK7gIS7MHo+YFx29n2Zdvri7gJANLQMbMshsg8MT8tP4Nci4hbTUZ
U47eH3rC3+R0EU+WGBuASlUbptdNQr3d/ZWbWxf9EDfTgVV7j0yVlM3G5sbMpBvS
Us2/oncYXWkyl/sQPXzzgDqo3uAPMnux0T1oln0kQlZkyd+zzbtp90Z7y4u2Im9b
ETME1DelEfkXpE5M6ovAqq8q1mMLyQcWREYgqTzdElCE2Po/WBOObSkzXW+ZldEd
jgVjUG7WPYIi5Tc+njrSgA7JgiYNgAZ1MVsBX81i5K0vlekvozwfEJ///TzIpTaZ
P89yMf8RAujvZIiMe89ALsce1WNhWJ0XprMmaXPdIN/zl68DU0vi/CBdTBDFbRyj
AN35vi3mhOMJZKWZxmqlk0ozyp/rBS7/a1ufHeOAM8PJdgUhcP1frGriltzS4P+U
MxvldczwBEnPD1yQPLHYqqfxf97K5WiM3EwngQc6a0KRGOxAU2qVmuWPXNnOU4wu
7zxrb2Fl4XKrE+25RUImjyEHA9P55UEtJd6Al3W+5MzYmUCeYvR8raHrojYGIUhV
9cNgFd/IGn0Wvhmw+jYf3VHLiBezUGTIr4UmVZ+D57HluOIaSR3jcssqfqGylgAR
ebfDscPcgvPkE45Xmv/Jvp7bEa3onFRJvy8ZMsb5w1BZ/HdIiL7mwdZzZT+ziUpS
GyJvTx9DyiN6gYsLnd3y7x6LXliPV95ujH2RYDqwQmTZcDUO+Zd5uWfYgFgwAw5u
brAPNfkJJLZiLs2cR6cJsBEuHluro4/DxNS/4MnXmgg59pV0hTUw+B/hQh1608Vg
TXIZX5gChuXXZ8XAO4N2yJKJwbPlU8ldZOjYzh+2bKKNDJHaQdYvu9oxGzISate4
KfQgGfLA0C7ajIRzVCKcvvilaGhaHSMAmpDep//tQrUNBulW5yKqg+S8Jx2lbuB0
wOJxuxnWzJG+7tjUpYGOyagKPmJeGX5GWh1jMa5K0aXYgvuK9RzYjYkZUzYyDWgm
1MeId6xN8sSnf9DtmUPSbj2kU1RFJ2AMRazESVfMT28844jURoNVA0C5VG+4BxAm
YMO6VvzQGfGOw6eraqnThKl2de/platkJYEMMrFOxgKIjIrN6prbOiL8a4jpj2uL
2xvlcyv8/Yc5SUgsHpXk2YrdZXfkYFedwc2BvIF0kQdlOnxojrofc/pHL1TeGzsM
5hCMwH8el9ijzlY3uCEd4OiqsU9WSI9UQd6hkYjHEU6B5+gsZKTgMducaa5sEU5M
G8xYyJxQ9yoLzA3IBlZFywVpoPkAavEXpdGpvp5lBl0a82wNsUhIg8UuXzh01/U1
GZP2eeRdfwiSNV9VCIxNIHdKV8XVo3Rq7jyre8VDfNYrIKr2av2ZocdqLjL4YJDC
wlx4lUt0nHe7gKm9MNrU5ccia0i5WYvaZqYBKnpEMx1dOHufiIGO4ArDbne7TTYv
PP5Qu+wiU0UQWnOi0Yzxkm3O9pBbxspRvx2bOYYC58DP985Ms+TiSIER0ubGu0gr
yukxDnXXCwPRv74aEAwHTXuKvycbQqdOU7heFxQXlPyNggTrykzJCn2nzT3Br34C
M2rlCFRre3mNZ83aQruvH186vbyWCZWZjxTDbnSEa+u7Oh5NJl90CZDpxuOr9/7j
R/pNIDtHPU3sxbPm4H48r24hYaHBir1AZLS+oJM/9zy8SEdJlOzuK868uIihswdb
Jnb3cRp7E01wkDTdX5zdbTiHNBNARPyQb8neFUXDBsCfqHocv3gOKIAwWZ9GDqQd
ji/kRadkZxbEnVeTniC4Dale7UADOIdW1rdxw6rS9upnDV683G0CatlSXwbHz5ma
SrfOJEepujqeGCcJ/gRQjSYrlVGRDURRx3lvvCEDa/u/+WYJEJYoDTdjmUJomfSY
GODQOMqz9j9ne3IgVlzWCBFQVQ4qY3mhFknt/mPB0Slw+6I3V3dwXOnHc9om53Xr
sDG5tQrXXRUJlJiy48FdyGQXqH60yDVr1O32xQj3HvJCF66RwgNiS26hd0J5J/xI
ewrw7MZNBY+qbOjXKgrthGaTNCU9AELbV1Ef2619VI2w34pdGmEIicQOdS3DUVxs
UdkGkdyovuUvK0N35OgdygSIKOQlS6eXQT7KtA1T+sq2C5YtyEXDoq/DujcFAaxG
HBgsvxcfDUQaN4IQs+hWz/5kWtLVEg1vp1pL6lnEM43XK3fK+sVND4adAtJuv86d
PLhV3xvv9It08Y9bXZw+pypj3+DYn0E6Hv4kv3u03AEzlg/oH80vs8GtBsnwomhC
yKZ1YMuNbiaxQ0yFTsFksYJIOa7Sg2Uw2VWOsCImx7Nd/hKvt2etTfniL90U01+N
ID0Qvpv5dB45xXsZGS/0/G0Xiw/sJaVVAsCCXQ1VfoAp4Fgu3aCx+x8zcwf25WAG
CFNbX8yyY0Ej0G11AF2lDuMLR3dSJ0AgmncsgT2HocfsvqDp4xdfsf8dswNtG7zR
X1VC7krMAI+vNthsb9Kg1hCRCV07rPlX0hlsdWuo3kMmOUbfxgaiUaOWs0tLQNBy
DbDaokwjN4ewjQKWnjqn6vewMCjK3YS+AP6Itz1OW5uQ0eulHw/B4I0A8PptatnG
aPmlXoumFzYIs1N/4/6dMOfF6ewWUqLMwuG7yvgdNQa5wb7z1d5bZodRFhO+1GKm
nC+wgmjU+pGnR1hL/iQG26gOIgVMz6o41m2B8AMSnlOl9wpdPeD8SmRIhRxYg7k4
SaD4NXDbLpszsYvCKTY/zkKkAHcIs2RWJmI5TnaztWwuku/puOa2m0pLmQPPAFrw
eSin8MHrLK5OxNhuAuBhE+FbNw4/eMcZfjh3H9M0/fOVdXPKw+VsmxXEjVwrjwsw
Lj1XdT8H3CCVoIWPGufpbCt9medbWdmrxSbi7ApIzd7QLTikhXkwaFFNSj3YH7ij
K6i9IZgfXILnhDRKl3Co5C1s4Gi6Pcjj0rSXUcxoeu0D/mv3fbuioU7OmWUPC/cW
5pBvnC8E7Q8FPmHQ6//b2eOAd4KUY0klm+cU9aUM8HlDjDn41T6nmHPL1lfpCfPs
doohjq5MNKl47o6V6F8jT1juiBC/JeT4MxQvbnbBHpzMWELV0K9pkhUxHdaHhcAq
noJLS6LaQTNsiJj+0lcJ+wtLpJBFEsspwwHx5c2rlTbfuA3AWuVDjHtFtIIs4S5L
OGepvGi9n3rosrwbWw2YcO3E0/z8TjZT77owrcJ+FHZ5Zr3SIv1SPVjxogQEkEYU
jc6aPRIWyOGx32c/Q86AeB6Ygn6HIBhukMVL0eqg2gJ6s4MRgZSrq0nAgN57D9qR
7Ln+vaHS8k4Ki7/OaPGrnVnwa4TzBGeexP5YSGa8XO6veqC3G837AOWmBa8oP/w7
iXGa5oT8f9xFj5eTjdyF3TBeQuro3uTifiKO/0ihxKVkByDbV+/eZQHpPeBqAvrL
igIKwm8CnHtYJC5ofE67j8NyhWL/sIlGf870Hr1KU3629hU0Z8kcO6VG3NVJYsnD
mQly93PuzYPkiIDmrqd3SwTu1KSHf3IbrQlzxB6YUVGjQ6LuuEEyiaCXCDFnxG/E
IJ3YI4H/DEHNuRY9rMVowkDxbtPShHd538vxpXn9VtmRa+OuGnXpYVuVuu0OPRV8
TUsZNdMBiE/QfNKMqgQ3pZjw4lu+dgsWAicGKn5YY1zddEQKASD/wC/luy7vKlGh
FR8W1etOxLjDE1v42vwpfVSDsKq2Ba9ouTMLgBPfjLb70rTy4eP0/ts97QWORNXy
IGE9uE0zSmUszv8z6XCywWS9GN2MGoKOmc0McEFfUff/J3WIKNAAwYwx/d/hQAJI
t8DrwMMXsokfGkRaHI0qvTrvsUFoqBuICE8gafdG/KuPUTimg5J6SCYMtfE0dujT
rIzzPGWJx9z33KTNGUBR6bwku5og239vBHj/TIOXyI5vDrSMoYUSFDeFar6cC3bb
IiuScmEIBHLHNu/BtUHP7LWSv6aeN3gi31fkMMszPYx6GmfCFL+WjybS0vhE44I7
OuP8isT/vsqHOcn5XQSOcLIyp64y14nbMZLIQr+pqAswa6nWGLoz3L36pj7JVAwV
qtwrlUa5Ciswmyh5l0q6EkjWzwnT2XeTDNgcjKz2GMHR239uqpSSERu9c2eFskzC
1q1esyXB/jejFN386jgd1hYEVw22Puqvp4MS5O/lMIGTUZ2tMNF/KBmlWgBP3NcY
wKgdfNw49hon9PYkdpFGthaoEhKUMKt2/TNHpbvIpZodYCtyKd7czVPL2u/63QZF
nPJfPfel1SI2dppGJsdqwzV9khkaEonENJA1wbZKDiqhHzb5jnebKhXiRuYgmFWI
WEXnI0jQbPwUbLav8mVHDhh4S2zwsbdp5hdoRt1KSV4+v+W0fUDgo9XyGvzUljRc
0HMpx4/76BaQqybZ+Yw2MHRLzgrZPuSYEixsqkZIUQb1y4vyd+Ou6WX3gNx6+GLm
JGU2hobYpnqu3FCzZpjo7RQt/stusNs05Tk5u2MSj7OPcXEamxSlttbzoZqPkgZJ
2iXOwPLukqv7ixbbfZ7ulL1ATYdV914kfWgxoGKvrbBLE/OE0L83r48PRE3ZZpCC
qW+m8+8BwCUigsVlNL0a5xaxQg9umWCL9n6wwLEnM/dIj2p+DJDbxii0FDOeTXYG
De6OdNHLdDmj+4pTeeQ2c0U7dRl6eAje50HCJm/bIW0L8r6jV25cCVv5NbW7CAk7
P27K/OOcM2cG29QebxZQe3bqR6peT3KxoGyAGRtjlL6q4TeLwKTzuoE/kM/uVQe3
FQxzX0wuTzUvmUIwgo3RO+Xg989rQMqL3xUKEL1DPPImuoPMiu60nsoznF5Z6Fsy
CekY4vS4BUVfej+MEngb6LCoMPyTepiJhNWggEeij/Ih4PXII4VIyUH4CCu8B7Gb
vguF3M8myXr2jclmDjtL0gsRzmJfeaXlMWfoR//lFep1yNMRHfC9zpgkR3uoBHJn
vtLmofHVw/sYNaHPmp9lmgRciBQhn+/plbucv1Q3XxkRjFpWzrjDUx6G76MeX30c
+9fAHeDuQdbDjydeAVfB1ggyVQ/TrvltAbbEp3HYKxLRTLlwqzUtvRvGjYoaGE2c
cBmgEa1OFzx7jXtUMApQQt5Kk+R+L56aoVEisQqSK5A/WJm3rPhCRUCmMJDv/poy
M6WVXcY8VmtaljcxJi0my5RbwEgmQREjyY9XDlOTbMDviHy437IKQL0i750HspfM
Gxk2a23beODkT6AZdk7QiFqNjbNVT17/TyWOhfnjVQ7BlEgj0obne7Dry2uDmHBu
pGhYu0bpLQnm3pJZ9+NqWENtr5QqTHyHQcSBjWoMPby01/UN4Iii0VXKcYYa3Sdy
ZTwK+DnThSuz5PsC1C6JimJIxyMuDtsKObpOx91NP1UeFI0GhTyMz97hcvquetyw
0nH5DMwf20b3lSFqO3xS1JFN00VUoK8k5349gtgodd+TqZnZXaIkiWM0pCTOB3S2
RyIbW5/KrZ4VHiQc2D6UyZXw/zJ2OoR3yZuqNNyHdnjVamuL3Xym6dvBxti8/7Q+
y1Ae/IRYeDfY4Pzj/y0mBKFaxYyyrcQpTr5VXCQpgYuKK4FZGginvYeqBJXwoVah
gPn236icHDmIQRKWFgaTDppwdnWNe1IEaw7OxhWwbQt918+7tbpKpF1oJJ6oRms+
cNyHgsPTmPJgCwl6mjHZVg/cY2C8putWbTFGb5/A4HWJf4rvbk4pgem+00F2m9Q4
TxZdeE70oxXG5HsYY/+Lf07sZG6sI8rskV2t5z9l61H2q2LYsgDvVhmaqYngjtOg
1caNTQDYClU8n/DAnbgBbHYq3esmoVV5TrgVlVYky2hwaI22bz51/Ch8lHKwC9u7
sU9Jl73T1wK+lhgur1xXDtMHeu85xLcn/UTpuUuCTOgaMii4ZN3P2Rzq6Ybvd0lo
ndxgjh9+kGYVbgW1a8IeKD9GAfIgJ2LiWkXPrwD7p9VZszzJvNNRHdpqt0wXfwRd
cOZerUdcK05bfN/FyIBzeUctveU2LeLfzgrigKZRZVwVUadhnbas5wbHZR0e3Cw5
TUHmRDPrthNPGyDHgFZuYSh29Yth0ihwxbxaf7wbAeZ1IDCcu2T84uga6jKGKdlO
PUZj0vDxjVihaOWwQFzK6Z+bW9tg6ZDhNXlMQbea/vdabJEAJpsr0P0aD7UC3uk/
7Q1Tl4rbU9fyo4M1jP71INX4+2mx5sHxF4OdvN4XUMr8nsQdDQL6eANNVeIZycy7
+dh5BjhZPQJaS3lmvoMRrKr54pbFQcIXnKcWmOXIzJhA5otKmnBxJwuuPJlJ2H9h
Kk6Bgy6JGzO4ADFIFBYPSGHUpPZ0hAgKJ5P9iMIuKCWomoW5A6aFGRSIF/nCg5uZ
mgR3jWkJDi5iku4aI6wiPEjDOCiiIMjG3xqIG3+lYEFKRrxgMILrDkFssH0mw/kJ
5J1fkmGfIHyB6q5Thf65aHuY3VfsLDx4IsSfcJSJwC18iG5+Q1JW3nv0+CDXyJxX
t4vnCTyRSgnaDKco458c0QIadAQyLMFyNZvoM5Yh9l2McDaxTi+tDB0b8nevoqXy
zej3RJWE6DHQURtm0crF6ylACGNZIqShlv7CckvW7qKQMGod1EaknpCwjmp+fPNb
vvSjFHY88FgHaEHEZ0QU/0nAJjJoDLE27s7349jnxBWv5f7bqW7r83ba3xrws2tw
26H5aTkoQKpFx3gwtPVWvTS245XBXQrzo/cQGn8QBSpP6zl7BUEHP8pizb8DB2Yl
cq+YP3R+BenJGFnBNW6lgexhUYFJ/cPaz5au+NLac4jIKyndKNhVEZ0HSGNM5fzv
UpPZNwIZ6TZFwzpeQKNyWgc8YnJouN6C8zts4RlZF5cLWP2ZrP33YAim69X35gZL
ybNt/Iiyo5BbVNEMlZlpv+jHAcSFEHFZHaoBc8Jy/9XmFcZJ3ChOWwGtNN8asfYj
IVykIZsm+ROKx98M/aachgPr6LK4qOiGi5fA2c6Wzq5NEcwq8liMsn1lkjyOf6nP
xDebeMKLaCEeGt0CkEjkmHRq128V+iVeJCp7wObTZkJTGcnCyBAR6b2cHOeqVn67
x45sILPDo+MG7u8AE+Q7hhB4UfjDXPGuoveUK/cn/HVqHHAQv2V/BLVEWxUOJB7E
bTxgNcJXbVLuod/KwWP+UN5IE4mls7BIIiK6ezuwzIgNrQyBXN9hFOmv2D7Nfoiq
FaVimAL12rJpz/lb6FnkQ6E0bjIgR7/xRtqB3WnNE7GJDD8O0cg60IRSR8Hj5xA4
0NMXAK3Z2gXyNenGfjXzIgqvR1HBn/LsJC17Kx6H8LxuYry36N8A8AFI172xaaMS
A983IY7DPr/YrwHeAeQA/CMFdtqsLGVR02kdsdIJ7n6+TrdOuXb+jVlWRCoRV2/l
l3dF1fUyy2nfPm5Y1xC2g+I6cRa4eD7LxIZasDdiSxUTF8G/h1KlS1Q4gef8vmaz
EOfhynj18nmV06/619KcPaXJaVjKlNXrPx5QikDJUhudwpVAHYne8C3v85eKvYZM
i/2Pgk97e7DfWYUsQopiRN059IzHsNaUQcP5DJMP+JmRzt/jwRPRb+ULr017f9ny
U/b5cfnLwyiYbFZ8vWgpq4KwS/7/03E8q9aTocHy3M1PBnMaF8ytq8DS+t18sh/n
MQqkEpVHm7OL8D5o1NMUw0Q8bEr52vuCQbL7HyNcyIy3ZmC2K8DRbU+9TqJpuIW1
EAf8QsJfKyjobN9tOk/irW8ralmcgnoaDVfGz3SdOidpnXeoxoq8kWZQ5ynPUxY+
rDgG3Lk22zP+XC9gQMftlwfYM7CVxnFGSEn3WNrOHrdr2K+eJX/KQpAKmZC8uA85
P6yEUuvRuW/6yWzJ7ZMoJtIj+/+naL+1+Hcqm2rrony3B/uzmVBxytB0VRQl/qRM
IXVAOkMa5kKAH+k5SwB7Q4rqCV+MxE7EZZ695B3NhwUCShCsBaYBf+NCr5zfZV9O
35B49yqdZByYdDO/qQmh/vQpZs7ceaK53OvZjLzAY6OX+ztoSEj1D8JLtYB75kpZ
ggQFSPGNNQHH5Kta03vWNlmAEw1cTpg2YsBS4+G8tZXdoaFqeqgAADUrlSC3eRzQ
F0GB15m6EZtYKSsfvc8o5fe85vytTkRjgHghBkh0JVpYhM/x8+5sb/ZO4fiPiCLP
cNVj8+GcjOMulqAH/0wpqQ168vvXTCp8eOeJp9z50wqPvGLUpW4KhbddNaUdvpsB
18oo7CPXt+VYdqRaDqH3pjOOhEaMiXEYfhnaEeZya8mLws5XjI2HF/BBys55V5vd
HRLa+XmOmEuCeOdORht+NDIVg+FILDKjHLJckD26iFxN6KcanpN4hTY4V7xgx1WW
nqimUWP4DXQ3i4Crt8/XaW1/7y4+hjLYE2bnJhcAKmTcM5Q6A5QSXFplpX9sZ6Ip
dDyxuphqRVbg0Pr7G9Sp4CEMscXa0nu5ok6UPQ+oUUnj4kICd5rp0MqdcbE/XNOE
V9ehsnueKgCcu6GysVed70zhJtjcJ4KYi0eoU1PaLTITwGssEDE/xL5jwmmfZ1eP
GQEd1Vat6ckKcaBOrjOFpMLYpYNCgsY0KGFVa01vtd+pHImXQUYsJ4qtig5UG2r2
NQo+qAK8hXkkXnRgubLUTd/vdseMkVhq1+HHNYlBqDxV6wC/EoXZiep2dtgkXmS+
Xt0rQ6HKtP880Plco5RwDRxx1szHjc4AclggZFUa31tV1MstinPcaUHAbFJNhxsA
batiQMoe9fnRhgZMUaiYVM+IFcqjcSnY2Ufz7U1zRPdCcckG+f3oT1b5Qz21MCen
SPR8qDxUgV9wcvLLgnsiW3qzAIHdI0xQ2NDLApFzyheXRKQ/6yN6HqePFl3tJbZs
MIqFD5XaJXuFSrHSj6shoymMale7WsrUSgXXg6kB1wv5rz0qqmDGD0kbLnTY0o4/
YVWcuJ0uens4qg6pn++JRZcv3Cp9f3jctlI3GUAdL7JoiPYa9vdjEVdOpcBoSEGx
jTwtP84+RhSBG0SaJvyGAXP7Jz4SXrZzK3EmjWVTvw2EmedGYc9kJyBSF8LHxEr8
BIeKU67PnIgwJGwuaEpbHfzyePNWO87nJ1NY841ExCuYVKldp5nxUJQQPdTgzdR0
qWO1vydNQd9hnIcZKwpYh8leaMR6429Obc8cOqjqz0E7TG0/ZnDLrYDN1GYAjPHN
zuWPbVMtX0YJFqaHxq/DKUAy65VP2IJ5A+TDGiDdThNFsHufcrJ+9KNZJ0cgfol8
obDqequaA11BLhEmJWozvtef7BjX1LyRYl3mFMY34TWlCyyp8FEy1vCzECkwlFx4
OxjEvTMIn/0yJQiYODc5cC1j3bcK5I53NpOs60YRZ75Sy4AIliXFfChqNu39tTKV
b1k8hKgMWUhU+9wHnHxEwaJOT6CHzjjuU8W9vRla8sCpy4TequsmG/K3rxYLk1N3
zMrpjgfel6AZMmd2UC4FnVJi9I+0ocwICSNIwd/nAVPuJiU/MShgk6ANvhY4O1mB
/efaPZadTLe1BcvxwagpmHYhTmM/IL2BfSy7hrng9vzlCTwbC83kcTCOdEda3w3X
A/ctds+JHmn7KwTM7gy27u8gXmchhl46DPBoEUYfk+0BwqywcPNkyJJmzFzU1zlr
MGH1ExH7d3jlarmIXroRwclMHrcPkGWKo0ezcIJJLEk2K45i0tv6D9rgdfE5Aghy
35nqF43DaqI6qSLG7P7i2h0IVtITMh6bimc3fcxbk0c6ODu6Pnnebp5oppD/eEgf
r165mKWdFkCxdFeApev4sULN/raBFQ5JB3ZG6TYSLX3lGf3q98bHWruIth1Epc3Q
8dhG0BarXYpycTpWWmPy1Gh87C1tpmnU72rtC+dumIQvkfeLxEpsyEqfPFdRe3mf
cyti4AUIrAmLn0OIf8Yd29+bHdRDrkCpOlngeESY+Vffd6YDr4NI2hAzFcnMM2e6
yHXegBUzxRmYvkFv0MBjPbEOY7xkKwLyY9irmT+jLfzXxAHW8Y/BVy0hmamarE2Q
7gedcvNe1CjhJep0SfgqpdvFct2MeiAjBcuByxtqsQJDDbrNVRBowVBneVLZzX91
bPynNKdKJm5yyHnkaieourXeoiPPK6IfOWlL2aa5GJtf5FjVeF7h9y0wYXTZRApR
H8ZtuNwg1POom7Vmo+UYkSR/6/F41ono6k6aSolG8oAqe9sD8kIrVgfkZynCJs+R
PCFmgVAMpB6cfrZFuvP0cIHBBXvs/+FA9Rp4CozThEoWdOUGPdsMQec543jv+qD7
FTpKwSHABjvrbgKRx7ammQaTL03yJm9oS6zvk24gWCF8p4mMAnOfqDZmJnODqY2o
C/7sz2+YViFt8a9BsiqF7zqRY7EeDUIgDWccxA8d5SWXej8fw4PEvN/RgzNZDTKS
ETi5i7EHVyWekZuVzxH4Eaq7kdVSW3GFhb9peng7jcIsmibnZLazm9yGmrROFFRp
shxrPUzT9+HFuRFjO535G1hlbx0kivVjrO4IvufZBucWNNb755rZ1kQ6jS2z0yge
PPvaO47Wq1QjnQH0jet9ftfIH0adT9VugkYUjhLxNctp0J8mw1bgZy5nyIGz/q2t
z3MINJj/E65ipjyu8DOWis/5sSGK/x06MmKD1T9MPwsf3knsoNJSAcCqtzXNMfE9
BB2QHzkAdmA6fsnkFvbSMn72mjLkrjoN8qr4EeKnZVHHD6SH8nX7E/YEvNamEdoR
fD0vgfZutzxRWCSqCD/YutT2gN8CRq2CwZFBhjEOZUprPnKyoMvmJI/KfEe4MBZ0
N1loSJqp//OPhcG7sSSzZFtExXEz4dPqlOxxTCEcNZlgbr1XUGq4BA4wOWA9M7r4
ZC/SlKqB/0uUpRAw6p3rwVCQzBdjIn+fAgNoGKfokWmGLtH4L7J73rQ2/iEfTRLB
PSopqnWRlpQBcu4XQPfKYcN6TfhWJE2XDzMbL44X941Yz5vRqMOeVB4End4sNZrJ
tDrPXpUykmi0forI/yYB1n+lQ0s35H4V4gTBkGGejkDrmmkeiQn8ee5zCrCzbHS5
sJsYQfHluixIupB2jtqpMSiSvjqPjVt9OHy7DshLGx5rwveN+Xkdu4fnyitP7LdP
C329rSc23GGLL3qpYtuOunA3rd1EAU/5LnajHBAVIc8FGBMrIk0cKLLEbPaiffmy
u6JdKtqtq3NWMT3xVJIA6cdT50CS4Lu1mUUw+YgMn/DvR4qajNoVCbG30cliGZE6
0ouBryaTrz8/ORFolbf2boUIPMQCvfNp6bXECu/wMoEp0ygFBcMmjkXUSvbOmG7A
F/FTcZf9s61UV0Mo4AmGYLrv8Zb+MK/eBA+rEKDtcUhBYPq+hQXRsv569QonKIty
Dz2up+/JdXdzGBIwBZAY1Bcu8WPVspfRknaetG9TrabWlfWrdH6GovNABysVj/qQ
oSe/ViISus5W3LRBRZxjYC/aYST+n3lOpk2nDpwhPURHqRkdfu2ePlln29OtDd8E
+pzpJ4IfX7F2EkUBJDE5shqaGJf7g2XyV/MDFILBKm5ca/A1Fv6UVAucjYFmKKzx
ScW3eM5nJf5+Y4VOKnXa7IczCLefXISo4GrETvPunBEc0/08M+OXct/Qi3IKkvZU
THd13j4kJjWatLYEPmQ6c6f7Pb8kkJHnMlnqZWFnqAkmkmsfJokhcV5Y2na8IFEp
X94ImP/HniQFh+V+5g5ePSlkg5KKVvoC90zgKO54IB335gPjr5+/mfrGjYVnK+1t
XqD07oax/yelK2KaMuPHPvjbAJ2XxuidUEhVBa6c24IB0iZ/CC5X4op7TPD0X1Qu
SXKttNti+qShVbXH1hOpWCXjv8WgOZa8v6dFt9KrTOPAzV2Xh9Dgt8M9rtie7Xzu
Xj5+AQOv7/mzcvxy+cTP3fgREpN0J58gajTW9gjhMUmVWAjxYQY8rvOIa6zvjHkJ
cMYGxqofxKs640QrbM4nUkIlgpkZDqq/csjgLbrSXMkJOKxG1+Yo2HmATgVdqnbC
RGHexvvwIaS6fL9xAybTWOuwoeakzxcxC/mnCD7rL+jPi4Ud+bEwitWhMaln76k4
PQjKilRzWQf6rJ812zh76PuweRcvc7BNzsesRfLVPde6cZjEaiGVrCcYrb7Ovf2R
gPStbkWtGXHU0dF6A0afcpQI2dgD2FD1rAwvqrEbHTT6JvkkxKWovU1m1YHB9mHA
m80oXys69QsRm6cSL80a/ldWmm0pQb5xVxq/R9Dz8ZdtYhE7OsAeA6ajlaWQQ1Rb
wO8ZlWaUlEtpG6eXrZIPv6SaCCcRAx/HddP2spHYVs07zo9mKpWYjqCUV6sv0lQI
zu5iPyorEtTmyBKjMB/9jRzrJP5n6yKDPZsCCKi6ATf2kejW4IhGB8G9xiCZY0Fg
zurqT5lHu2jlExqjPFwzOOxOXuETLkxHXSsRHIP8hreZ6gm+a7PtBy7r8CNLl/NG
04kU9Fj5/Q0/oqyFlQG1Jtmh6d/unvpIL6k8OOSGLw8yIkeL4Dvuzd0ed6Ui2M4Z
+mAY/tkCKGEeWmBj3ybLCnwC6q1K/D1kb5xXIFDraMqrFheuQqcdAVj7qwWLQ+qr
fBQmkz6hU5WZOXP4El264nSHn4c4GRmhvmrRL/9Ih9BTkgJkM+QEsSBH6/CIB3mb
Xe+rOs87b5LmnkaiMce17oQ6jyxzG4orTVKH8A4eJBesAjfvr1osn+q19w6xPkQu
30YLDVHYMNssWMq3BPEqoaWy39N38yOkNcNd/k/DyUeA3WLW+5CtNlEbhhks1nJP
OAsASxwb1i4qQqbKV82rMRWn7io+y6WuOYcmO1XHY3JtqbCkjGJ/zb1l+1ey+6HJ
moL3xrBu0mTAP5YBWcGjAlI1cW4bu0tmDkKWj2ZvN88KVIiaApBb05o3ErL/cokw
zDooIaVs7wE8pjy2JvCpv34B4OzDW8Q696hFtbi7cf+X1+Zb4NFr/9EIKAsWuHpP
p78Yfe9kL1W4ysdcnGjL5HFXAqWfm4ZUhs/QJ6BfJ1UqnoXEsSaIq2pwYLaE9XOD
+hsbLz0XiIiZYpssV9rIX6Yn1FNY5us3pJZ+Dc/lKCOYGUThk9l/J2a7vD1PakhZ
2ZzbPYQv4SLXVJubiJnjpgnoA42avhJvQVvvdh/zYZOy+lSve+Usa9o4To3OULhb
h1NGW7JUf0OsU9svODekJ4ccYL0At6ZP8FM4QL/+DnVN62EVVkPQcUqfXg9nfV40
VP0g+Nf0TPaWeYTXTsgTaUHJlOMlyENtF+NFD4EmzYjSLQPy5HnctjG0tS0qI/oG
WRSWwGtGJ3Aas81096pcCJcBJXlUWUHdsHx+FQzg1wZSLBrCgZDw6gNpG+IQmEOw
UoNQllZLJ3yekiqdqMsTpuPREOU1NFh5x3CZ5q6UitgX02fulsZdhMgkxrr47ZIg
Go5TSPVJIARwqVRBJGziq3O6z5CGEnGgryxnXzovHibIPPVRR0ZbN3ck+GpNptqD
b0zl9PIMujzl/SxvB+UiPwRig/ESMS4J7WFMnHMqJkJXq8pVrbx6V/dzvTbWpzco
75Xf8yrE+zou1kgOfCCz26sWhUg9f7j1wjQgizUlGSmFpcjdrmiT1rVitkXgk77L
NSPGcfQlppsoF2qgt8hneDejbS7TcweNXkC93DsDEr8qGR9cVegazuzl1cpoWOky
MDTJCCL4K4J9BUbPlWTxsIJiOi55iYOYfLWRwBgKJ6DV1ptwXV0L8qdW531ANH6i
lE1iAFmSLyIcTO25CEozIu78cLdVXYuWUTJyuPPtNNwUugmwX5C55o1Odq+2K43E
CfwbSMRHemUJIrHHrOP8hxrTVfK/83wQmsF37AZIohpDWu/la0a4upSQi3SqPGWW
lecTeEEpK1+dqRbxRQNHIbzDG79HJLqmk6zqi6p16+U3RLS/kg1G+fe1XBuS5TxW
qi26Uk7NZsk0hP+0PMw/D2J1JxKS2N9SJBVcUKmEDzZVUi9RQb+FnBz77Ffbm0pY
VUdRtxJSyiFTaOmPMskqmBw8qMeP/lPM4ObMVzSIlm8XS/FzvHlWqznxCVb2J526
Q2hc+P04ehBDrtVRd2wAgmuEL3j9OYTOKQkVg8NuriFfSOdM850+OeH1Kkh7LcFn
WrZLvVxuuEMjt9PxxPfdhTwOcRpOTJnz8nRmEbLsD8ryGiq5xaJMk/pIakSIN6Vt
CtezBR/jHSEusM7uiF6Uh40GyhMp4POSakMfW39jTQjBvhcUrodToIHYjbDNKqp1
NMRKTsiykC40bu4tEWvs5DxmpEBLh9LA+AjrHqHaeSQ0N0JPOY9BYAfnL1gUXn0t
qHY1c1WDzVkf1y0pPU+N762pJJxlOQnMxi3LFfJvpcQq5ajKcWPTuMOO4aQb9fuX
KXivryGuiyaKA1CBvBeO+ncCD5wqrIIg6/vzzgHH5vKbjTizyX+pPpXUh7nyvU4r
qimDm09ucDeK0RqD7HcMRc7o8T0/Vnp7r6C9311lwLss1bkniWUbRlZvm5jGZmAv
aqAZgJLnE4BJvke1Qbzb5I5A8VI22CuWw2+POI3ESjaJXWp2TPOmUASaD/TRm40W
k7Wurb5XW0C0ucIrUzFIfaTHi4pH5BWoVzirJ76YstIk5tIBR/2nGzggRqcI+xHk
YemAMrCDiTVijF2YV1IHMiSTJ0X4ed6Ku6Zly4XgsvsyQgR05roHwAbJ/OMJ9YUO
ydt2KW4nxzRqz2WKAVbBy2mRUlH/Zyy2uMALJlLrH0tBT4cJYITPrDSAWIUOOhVx
GLNF3Pk/YnaXENnrn584q/aaXX+aRWHROpl4kvPDBis9smEdwb7tVx0yhjeM496o
Eg0CjEQrHGyxVhR7Wb+nbIMXya1wYaoHkM+0BlshPln3zdS5CQJl7QYTyDvEB1Z1
fHWt9cMV2Qpp5G67ulE2PcpBmKDyxL58C7KQ5O5XZBesVQipwwrKDglebB2r6a/V
PkrKv/rG7/vGEnOUuEMuF0nNR2nivHHzbKRDB/Fke6H8GQgrwPlUap9PsaSONUKh
LHezpwAQsLkdyK0As9Hs8JLa7VvZPv45io8zneuaZxah2JEq+qc5TL1Shgn+zCR1
uxStj59NOw2W38+Vw3LTTkDZ6kyzltKm+lFPQF5H59KVjROairseq42obJn4mYwz
2s9EW+9wNia6VBU+F3JhnCrVHSDhE+0u/zaYgIxduYud3I3C4F2cz4ywyzWDL/rj
CAeSWAMU6gA8S+PCI61OTWYzKwiHujJH+Neg1NiR3eQCZPlo8PTQsbnjOqzSdAUW
InhjZyrdJL5tV3DS1pq9NIqAz4muAiJZ7QdDIASDPd9u3jMvK0xxeDptaiYABTVE
QXTqf0SOScd+pf7XEzpn5NkRI4JTnxeugFofr617a4mN5123EIDFBu0ndRGn3fU1
gdvE1o98iqpj7pQptsmw9mv3HZE0YKZMF76wzbpXfORIg6BAN+iHs0r8IadVg30E
a4oHQovwquLismCAxh6WlVDdDea3yDZKuHEvIvXzdgyOk9HcqWzdY7CuGJLnqiU8
c2bKZ+ut0BXIpPfcF8/wVJG8/GiJpG7c6ZloHmrFE33m6+/EdEZx6mZ0zzMUxFkh
qhAen8ztQhK8S3o5Eurlp8ZroJ84SzTbfk59hoLcztJlObKR2X9m0/U4a49xKxpe
3+mzhJ+pHMitS2RybGolH0v3umjZXldXjePufCHkapPUsqE3sxiD6Os9WDMfVy5o
E0pjEUaVbNZf3KiwNjc7oI8c6GiKWS1oQDGbz6InBiJ5MNkou+3ttumI4KWwGtPr
R6r1CYEkBpGMrrJsZS14xbjkOs9B1u4sGM5x0eSPYmQIXEcHy0pjCE1DFR/RPTy2
Yi2/duWci9WZskHs2NI2doXA4GAUnjkLXHVKBsQABV8gpaXBGZkPWk8O7CoWl37w
mtFXaPQJG69dKgSHEAE9QQeenXwOusekn3QVCux5Vl5fOtHVlJVzVR9hgmh54RLN
OMeKn4PnJR480g8NSWUiniaezERoZDQ3sKd0i0n+7sZlo36cK0pqRNNhmbunkNH1
0EYnURQnKcM+tCN7lMzLq3+vLUvF5lktCvnFuXAaKkoyRU6sjML6bbtwaVbHpp1N
97Fj3GR6mFdWFlkNNfSydNbFWzOF9OtwQLRpcbGQwlFfK7DNZ06HA11QIJbF4zp+
KPgpP6zCqVL0RaMHaP3eqJpX2M9w77q5Q/KWlxgdm2Y3+EkPWMswHy11OmfAOl3a
2mwfiQx9X2uCHV51gVEdNnY6r5T+fRyYk1bHuyQus7Rf3KZl6+3TM8JEXokDRoQy
9+6p1FHFYjrqoz+ZNrCR8YZSvk0jYNmfuRPUURRW6haUTzXWKl397+gHW2lX/FzJ
cEwSnDsY31ZMf3MgdkvKn3Cj7L9XgIEZ5O7u6XKBq+3NvuAdZxH6CJxZrD1E9uIl
jPDBHYVhNX+w9oVkGtqOyKjYet+0+6tqyq6E+oODdsdmy0F5h+VxjbLctGUA650Y
fAQWWClQRV49cGhLqu+eGcr5JMlMgkR9s2bvekc+ISBXBF6ZPfs7rSx51eUjRUJa
C8fS6H7NMgwBmUC7SFC2/pDDXpDdsEocrilRILYQrcWIbid/mydDfyBiW61nTNyK
NR5rLc5gMrcTJjQH0vjLXS2mJiESUTweuQgfa06iJ3Hr1aoucJmSdQMKJ4LzB99M
HmfhKBPJJOVrIL34Qba0ThFcTTOuT1SacQ/f7ZpiEKrk9PR/eXswQ644BBimipOZ
KYZdimEKXqpWf1yorJSfC3NqalEp4nPJpdDIdYtyj3OL42vmUdybKbaEMBYclf2v
/OcE+VO0mMRJp2jSCmcsye84Cn8WcZGCfxVPbCvE94hMWqaVHpkRvhDe6Ngx042G
MAat4AozsnApsuleKkNXZkDyyNjMAAzQ7t6XlH7Z/b0XheB1v5ili0jFRpJ3tZx9
34qS1pZq+9VW0Q4eVdWAKRX3KPbm4d6vggrI+3xFD8a8nFomP8d6WEEA9sOFhm3v
XRWwiufFWP6+loXDP1Ld1DyjLosidrmEdbdWFAZf/aX0e1qgaCbcpirUmnNJV4oP
xLnNopyPC6qc335Qab8A8J/2GCCaztD1ZTas8cKVCx8n8vN0tzRwAjAbEj2euWWT
J0UK+IysymEfWLQGSqV8zkUUePKL3daI9ErIqJgtmL+1EbtmzymD1GTsU7jyKaAE
etiYtjLYkbb+pqm2gAsQ9wU8mt7eIhDPDegpVf5Eip7aEDhLHrMQTSOJ4KC4oPfo
6DJye7xEjCRtfisw67UKMt25PkG2waHzMsZ4dMLOF4PFEQDmh9pxyljfIFXtXPIp
0VLnXqrimKwMeY+VBka0KsbPfuadSFKXJILYZlUE6Rw1ETZ4vLlXB5YdjpfWlUP3
iks0xz3UFbnJxGXu9OsaCBZUcc54mP5rLUCFjPu0SCUruTWgXdS4yaLyASqV/PLZ
M2uKzr+j5IjVwO2OxI86E9XWOll43n5m+JLQa5u7EYdkqoBL7CYK592NgZb4K3Wt
j/8gIOJfYGpwrZON7VCd2WLX9gEfBSLqwGKt3EY+z+WjREQ9QOJWgb+xMSm81wWb
t/gncPmNlITDP9HvH+f/DKGI/iaJczZmRmAsSsRB4RvxLb3bBAdrlb0clHqXaO08
6I7Bu9a8fuEJ+EAMT/2Uf27FNsFu67orYffwKevvDes7oJ3QVYt9TBZiQYEiLRu5
emOpr6MSxZ2Upc716y8PA8R4OsIyvHUjwA8srcslT8nmT8FxnJP5ZQ8eLGsovcrc
rKK23pgGSXb5EfvVHN++OqmxTvISpN3SBKMuSNodmxsKcPZmN3pFs4pa8KTvJky1
dFaioQMWpWNp3gheG4RJ8p/tXPQINMOlAm1jzFJn5LsBkk80z6LXH0X4jwLqYq13
gDHMokoFdI9ZXQKiBxvILfBfZFXmCzDj0DGuGGX4hT+t69r3PEyUdLOe8lic6ooJ
DVJEF5DL+stZfpUzhnpnbDUBFydtrWvIL10p2dZQEw6UPVpYP1HOXSHq7ISIXQmW
rGFm/xFDgSUo0G2lRNL4KKy1VxV+FgadZdorMXmIcl2RJl/v2aPRaHFGXSj6hL0Z
KMRzNK2RbxU025KBUJ1rmaTYyZdiVPK47D9X3yCXJmz1ogKNnyQdKGq5Kry+BPk2
f5Sk2CUTKE2CfN8BnmD+U3XJwyiNUYDy1FWlqnRjLXuqux8i8kJgftwDbLH+iz76
7pBFZiPNo82KD2EbSs+LgD84txEpRQfbs3QwDDPdVxpCZOLIqgX8PfPbkNVKwEUs
l5MI1VjEFypozqKzxj7HSOs18C62O3mDKlzoswdJlz+L82mgyIE1o8sS4+r76syL
bNGmagXOdYDAB4WBiy4/6N3AO9GOA+St3I9oIHXyTKQcDwOZ3kRK9iSv+jae2Nhl
meqsiCyBVR8Qjc7IwUBtwns8CECvmIYqoGPnIPG51zCRHK5MwkotcuvLIdybyAPs
L5XYoWY98J5jyU9h8TlzqPgfhahm9GNf7yprQ4XA4zJkicSqCtJGGlYgqbnnv8hB
zdng/xUupLYw4xpRDC2xohYWkyeZrsMJTGQW4FNa+PdJyIlyJI3NmbAmTMR3Pq7e
bXG7YePVBvFDU/YFIkFSxNudMwuwN6Wdj/VTHG4KuInKes4fJiIA8Tlbjxc5WrsB
4yL+OPnrWBNuhT2fGb7eD313OKl0mqxHMHFI8qgYsl2GD6hPXp6ESfh5YZpUCYjX
AyyLKNzqi1RuEZkJ7bH5sDM1lzyXfSfMYWR3B10ezSLLTx4mdEuaMkDdrR+ieS1E
Tf994+5RO/Hxw0VsQzdOfYQcd8vkpLZCq3o0odx45ATk9ieRQcl+yT8MtBHrlaVT
RqRyoavRmreOcAkAhvRxT9M+wo7W9Hp0jFm8q/I4xU1nZwyU0yr+aD6l7BSfA8b6
D9ZfSbtLNZNRcUiaKz/1/YiuFsxgtgLwAGV8SMeJp450Z5cioDOhaomJ7CErXLOT
CkYLyumCh+mYkYveICLF+v0DSVpzx8Z73y6sz4Nb2S+0s47zTgrOpH5gDgTFTwI1
+PdXg2UGRPslvof0kuR/OUgt9UuUb+6Hp6nUgLf3RsBR41ElzBsxPhXeN97VYFov
LiWL/uvZqWXO1V1uc1JI8ODTPvZFDZ+xWd3BSdCU53YEj8UqA6DiyL0wO1U23L3V
mauVqt5ngbNVTiRGKflK6XqUXW3nl6ZUqHA5TPQHeZ+4xLr1Lv43mj0r+4yKB/XJ
qsGa8ZOC+Ul5EApn1arAkXNAqlHeuEfrsvQ2g2lGiAJUQu2XjrACqjAo2El9RKSv
E2BJ3uoehExbeCoCQ/WCae3GkwzvIRzQbOEgfAaMih/F9jFJBz87+GhgDMLfNHgX
HseExnUaUgPMmyypRe4sm1pgZATniCyZFt1nwxzL6vDyyNe8OTUV77/97jZWZDU0
gAxyQ77bXS9VrW+hSt/fGHnU2CIPI2SKzVAVgv3+9fPpjHUmrRsnV+v09tl030+f
EK9rpYQPfsS4Ye0xjdc/DIva2TMoUUa7oKN0Nz/EWWVp5j6Ei6n9DvLaeQiHL8qk
Vs036Dfzb0+BhSAIxYJAgTzk10dbj8TuXAG3dZQ50BCATv0rqTDJmyu07THQ1m9x
8dDIfPGVUo2xCJw4jV017RSBxTvzedG/oz813WNgwAPUxHyktg+eeESgOF+gAXvD
o91x7EMfkPEojAHPphllEDxAbO8gT/KOoIslSPjThRj1gsIYMeOgII9NsWlKJ1Gu
jQ7FXZf/4f3GNdMtq8BMOMYR6V/d+wFVVq1KqB2Msu07gUbJSd9nzkSsNv3s43DF
/xTEe1WnFtcG5DiVTvU2fGj3YSPkuh2oY1qbg7b/VohA+8oaFATHJdCryaFVS/qA
Oo/DHW4L0tjYHtu2at/bLWKz2sH6vx5TdEstiLBQiuJUKbS6iQ+FMknyVOdjrN8t
td4i7N4ggglo71UpsqhyYWh+G+SALhuIWo0MJIsw9olRpsS3No3QdtmIhgov7eeR
rP3HcbdT/NzhNKy2rxm135nMbMALH8wpk9XwzxrT8iMS9VJzBPQsFItazIjZ0hHi
6sYQcip4lbv7l60eh5bcklwyMegUrhIM7Ab4uhJ2H1DZHIyaLsAYMaH3mgLIueEg
sdRYkoXj0wFTNOKHz2+nKuTnsBhvbJQ2Ta05twEB/EpwdDgd+ayy0bmSLx+FMLDr
D9Xze4CuXr/6JxXu7KhRH+saJFpSqJLbypBxKkhx6+14iSyG1d2VFQhDdS+n1nqD
iPf5/cenAgtzWDBvF4n9LgA7MpgzPfSVKbstSpqNujhqjE6JHisqrdHde9+VVgRE
SSeAU9Ujr+XhW74Pc4jlsyZngHEsS50Y3+5OM2zB7QlBuY6dCJj9NVHU/W7CSzwh
jtSJ+U8pL7AiHMIiCuO+go/U55Dvo7noLq902UiioI4iPrZFkx7tLUjyodt/RGL2
AVRmiQMNO27i6KbyDfZpB7R6tWqpRHYcG5Z9M5rsLaqPp0mdkvtuTfBaS3N52L1O
XfTXOX2DueSKRQbPhXeA48/XjAh2zT+uEujWroMop6NGyP+5+4WgnS80dQ0o0ySa
+N2Qdk91sBk2cikOsU02CcAlr3P+Gc/EEFkRStagfYztA87Emb8sHK1LjQtgzJ4m
hRj2vAX92dQUyv9sMu14pqu9WklfRlC/CI/DADxrkW8ftVm9mjABeZ03srPvfF0Y
HUoqEStqWULbPlkBQuhrcIFygegSoC5H9kVqftJdxIQ4aTMXqIdoq0ghhE7Nn2Xk
vxe1OKepUYmj5QcmyxG+9r4Wct8Fsvwnyf6hXcRV1W7egiq1/Wa5ZYrj9am5SaDj
KQiD0q4lDpmyydINWq7ZRFBwwtT/RRiuEOZXlv2UdW1G5rz0xUDe9blzIzu4feBU
sgtivfa4bqjaXYHldPC+zF68LKlCE6mSpjhhgPoH3tEsZq+fnGGydlVz/gOebiNY
f2MQXVo20EMbmodb4wc9UsB9zvfcX9/PjKPMu57aid2IEAnut5yPKm4audlngy8A
TmGmy/uxWcSriWykjuI/c27WLYcVRDHvtxiqBx9ryVZMbLM6R2D3Udivd3ALRht2
oMFF0Qa7YsctCPll0boCZGFOEmdg8NYosL5938h4+2HO6RmFGrzDp9GdHc7PnfwF
7xIVGb2c97yVxB8kbXThj7d8BgOoaIU4MrJ4umE5AZFiL++5sB7sHcLbMZMOht0t
cBNroqDVZxIX0YfIcuvi9+See3s8vasRXIJar3aOSQNu7jiIFyB7H/piMxyEpjyk
IEzpdTyEyCaXPizGtJnFC0c1TuCy/KtBzUVLmL97sPPxFvWQYlTcY/BxQlAkrjAX
87qUUEdvdgzkmm3/NtpzlzFMNjpu3dWhhKjKTSkSS9nuQThfLPWRgp309SVHuJEw
+lM0EM/kVSpFYLr7mWBBOI+u7d2C/QLojlR+c4NBg4l5GpVD6LRewlLeGQ3CMddQ
Doycb5tlaCmbV470vNflVT/PJqGhUJuN77LaHAueQlDFvoeBQl7x16pGMc+P/M0l
2BwvQqrCYb7+LTmVxsyVvXK/XfHPDm2uccUj3BeSCAozZy4VOcgin+1CwhXKj8b1
hZwpzLhU2Aja/eJoU2SbNgRg5FiqUDImm6y7t9VeP7vfNPQoYpB2wr8oLMs90WgA
3kkbYI/TH0YEPuCS9/HQVXkWmHyo6lnArREsLRhL0+gJRbZ1bI+uqMG8VVyOmv6L
kVCiQSEZosSrsIDoDvZYFaCP+9IxqS/P/UlNYGbJ7ypD/ZNNoro+GsRlLbPFNtyO
D+I88guYLY74d90fjjMJxC0RCNSDMKHf6sBn/+TY65/B3+yrJX4ukTt8TEOrFvIN
aJ4E00UK6L9vZmIyKCrFtgI/TK+W/Pe1A6INWJTt9LtmZipzWGmsJHGc5H/p/Bzj
8lBxvXT2Y2ZSRTtrrhTP2QMdRU3zYAqmNJ3+MYdWEsJu7EZH8SwqCAhA3C3I2990
QWcNoiA1Y3wv2EvuaZsEuR6/E7wfuD+n60bpFhjBdQ4CSAbyuMcOtq2MVk0u+MU4
MxxsVH+NBYyTakjTAW5W/mxa2+wMIyha9v+NxEn6DtJRrXGldXrduAxwPXKnAa6C
VPBYWTPkpsd0m07/7YiAejImGjNIYZUmxNmoI2ESEAwWXIx6i4Z+wmfHkobUEYLT
XqyvujNCcuPiLiF41ROilDzcpNhuQ4VU8xIQumcVkGGtPzZeMMxGi12mmszuar04
eAp5UTlcYlPMFW6bFVuiaHJCJNcUDQFQ+gk6UScz/6aEwk5xj8x4g/VxpRao8vZQ
WnZoMlbfujmeQPxfqNLkPd+2CNZgmcICpbjxKfGDXzCkJEIJkcSRrRxHnZTiNtko
SeqSFe8BhSHWa0nEYiAvczf9rNGF7vTzyAe3qxMXjGWUp6YNQVRERB0m5yrtxT7H
UlpKhrT3wY71VsYI0wnfj5+5RQI0708D4X6UuqeulFD1mxn+lOvita+smhiRhuk5
XA806XYKIB4Ye6RRuTknvnyQUWg3nTW70iRtoOqwupwA+AYvQ8caivSR+JNQS/mL
WW6k1LcWs3lpzH7X9k0mwHx1HLTBBtXNWf0zPSoOo5HNSEYkNgPDYnoJPvZvqFQw
RDYcwQXDraLRohuZqheVN17lKjlxvgfR5POeQxn6BoN+KvhSqP8BiNNuVr9AquKO
+LAedEWX2Zd4/3hIastCuWItrO1ZpaMbiUH3oMaKMkUQzq4fNGwP+A1z9DUW87wX
2iGKIlHw2rXiBGE6d3GDjFD3DegE5VUI0SGfsKyz3fvLZfiIgQRl92XnIZ2h5ilA
/bUX/G8jZc+jJRujhTYcoZhxewZswNsdwbzyjR0P/vNKZXLTzLWmo3kry0t833c2
+X6IrTuPUj1qcHVudPW07tYHfrJtmhnMHipVUHTx4MLJXbTnsp3SMN7C/RrDmBLG
y2z6ogsia7PEt2N5O9Q++3YB2102IqcbtQuPp9L41EayNs6otz4MZVZs3xedu3V3
baxUDpzfQzo7+KKKoJs0WtYpABgqogXmQQ6LrNsrBvXqtFfov0jznNfl0whWxZvf
v8dShWybQdBRFn5fRB+E+BBDe5KXf7v60PHS/sCbgjmC6KdjtMUwHu/6tVIciLSQ
oXU6R4H02vjVdERVnF1U9FBdIQUPTALs0g0ter0SNfy5teNjg+AsnVBygu5Afjg+
kCln5u2M+jd+TgB65ZbIDqh7U1KT/Rj9htfPIa8eN+lptzN2wIJ2ebtZUCZfe4FR
eEj1EFlOJTh0iPrpR9eYrRgHkUDqaq26fc/zmHqITUAoQWlLWgQsM9r0Ry+kgCMG
mF4Fyw3aqr5MSSNTbreWj8XEZk8+zej442GpmhzBriexVAKNEEi6umPrk8VPRIEV
lkDScD1kbWhPcIfzIVIT0DKEx/cMQfW88uMTsFTIi4sSaOrBWv9hKkRtnw4lTQOI
z5jD7UD9HH2SsnQl3pSuhvaSkOc+x9qd+4cpFkyxKqQKIb4uEMIk3JFR+tOWQ3Xh
N16cEbqcFjBcAX8Zlg7XWmm0IkskCj2USARJDKYH48de2eKY2MbO/QADi7roYZaZ
Dt4t1qaYGg3eh3dAio9Xa9t7WRtTtrC7ylRXnsYG6aWnfFPrMP65bTFcpzt4TkKq
An0pYE+8niH/Bb5RTnadH2D8GSUKpPZN1IOLVUh80qXzLUPvLtDFYSCHaIv1Y2dU
psubcmZVS8BctsW7D5b09GstzZUGfsPejIvwqDX3HGnfTQxi8uo/fYaD3snVR8vH
zoD1n4oO3OvGgoB0PC7lebfj1awHf+qeHJ7p/n5b+dST1B4T2bTW86mySiy85gAK
0NBRhPqE4ugNf+kaWuhshaL6I3jKNJiq5mS2jap7Pp57NI4tcjyUZtWyVc5CgZoA
BfjNgNOA8GmV1pLyUPmwFlf5JlymRodCimtijYwNcnhlWThbcQi6LSaMAtvfeK+O
3v7UYeRSv+L6oVYl1tSqCaYMXtho/m3CvigBO0d4sA9cTKnfwNMjPOrBDn6qr2IV
P+9sb2xBFUtOD+qSRu3rQ6NWuBwFy0e3iTay1mBmtomECIjjTdfNFZVWXEBJYaJ0
CtcCaZDVdpvZL9hSAA+Zo9MjcVdgtL2FZKBosW1kcZDLckFYBOft2zKARwvpm8Ep
Zn6tGQxFX7Fr+Mar+3VEeQ0jjPE3EpWAlAKk7xrwXZLHuP6GKiBQhtdTG90zYwjZ
nJS9mmdEZCDw2eCIz5PYLshxOvj8SJZVV5R86p6robKOjcy6+lz91Wu41UWwweBF
nyOH42YmGeIYVd1MGSHr6NUwXiYgXsxmKfUvvjM92Xia+xXWMcHVIbOT0wzPLfK7
IJOUHjQem8xHjkGVmUsiHbq0kfZng+elHCGmEUeZyfWXPrdr+lrIjRS72eYY5Xjn
V25lqLeeyZVrz78KNEFpui9z6QzxwtNeeZ1cV48ZIHgbVz0W9Zi270e1iSiNqYNL
KJ7gPEZyMC8xueeDk5qhD+vPVjyyxmGEbHbF13P+VvJu6aJ4rPfmJuJxQDYutKV7
haA8rysA89tWyLde3+17/vY3vJCxpGpJxY9Q5YNidWDAT2nbW3jU1lLggMjM+bWV
7ryLANqHMU9hcioSlcFyI8jN5OBjr8jneStVQU+0xLerlI+Z1+5EPTwB3bFsqiEY
34PZmIsFfeda4rS6UelxBadYoUQF1Lt33gW0t4QcOdABbWg673ABfLiqQ8W5aYxX
6GkQjGvFAa8PZHNF9b1PGEhkHhU+INU+p1aq7xJZyYwGdpQtY4Hf2sOsHaLXK56v
Ss6Mgj8Beqi5sbvk8eUsa7PZeiwfPZrzxJ7+++fScUFsA+26FPqP3BE7BDEnwgam
uOvcQRhAC4Cqu8nxjaacxJq0jw3Y81aXivHMYRPOKQaGPoxnEuL7EnCouoMVZzGX
jXP6feLODl5pS41V3yMefYrwRd9GqynLw/t3KXdEeROQE/iOqNhatd2X2iG/Y9K2
ecxZBymnIex57KKplcJzZGc6bQAhUP5bPTTPkH8q17oZQjSdg7+eyQ1eh8Q8pSbU
X4ajb5ELtJtg1ViWq5SEbdTaaYnu84np+MqlMvoWVUe5BNpsareLn6DsXFrYOhDI
DnNnxbX8LKyZ8/z1LO83NerRBBJRcujJ50Qdsmhzc3i082Oyp8gEhhlY0RjZ3gDX
8p/Wh3W4u4tbU+eCp0ZYw+d+Pf/JEeCTdr8cIeoQapQpQhQR2KBf9CTv5Tm8kjEW
Qt8pMWwFrdZI9zO+cvry0HnYmbllzdbbznXqaTMTe/S2c3PoFpcIVm3kr0htm6hJ
yTquMtFubciyLN6FKo6EAb7ZhWN2ZAfKl3IJWKUjlsxRjcrdN/RIKIXlcjK0O1ij
heUPFb65d1myc8YNCY3TakY1CEc4xKoedxahKBa9JB1qYqJvlGKLpe1w5xH/B+qD
qN2GDiPICG8HDgH+VEnGvPZERFvyPGX61jXqNB7rhzkgi3sU07eKORXAHG49k3Kd
Hp6NJA5LLpiU5oNaauSNkCTheX2bzBJKHYtUS2CGsCrGwXUcySHcF3WVOhYM8OTx
aFPEKKh+Ho30XffZoLOtcoKLZV/G3Dsbtb8x1TT5TAxMuLqpOtYWvXqTOpguPK3b
dcSue/07OumRbS9Hg9TxDJ5J+ws1TtVB0MaqS3+jnzcrJfzWfwsjGXsMOQztv1d+
wS5ixg/2ca2mXDKzCXbxEpLmKGQm1bdBSXK431m+0OUWcaWdMQEszgCheMSdpi6s
1Gx6V/Eg58K69psHOs4kbbN+c7YhD1PIrI0o6b3q+oiXsCyw/fHH7s3RuYn0qrht
GopCYOPNa3KrCVdCPXjmj6zFiBVgSMlh4ZHMx1JziastJYqsgBzP41M6exRr35w4
B7Ze4HusnRX+e8fc5+yVORziBm0x+izU4ZaN+VFVFUlzEhw0VH9buZ9epuD4Pzca
37aScVXM1GNpFcrKR7Z9XPzOOlTHTGn2BMEx9hI3t6qyHJAxF0y7CBQ1a3Q7kg3P
Sarw3UOYKoIOxci+/yKdNdxXmXloHo9gTUHlipjFIs986A+9H5q748hxdW4h5RPW
HJ/06XeuhNudrdt4vESyTyaWgdj4QjnRgXPppZj6LF6C9RgB8FNNUDCMLFM3B9/5
EJ5BytxbYjA9HpMdUdQU2SaGKkRiLM8JxkLiznlYi4kb2OFF63O6bYB0eBbSluMe
XCoPjqpsD0LGELMS9GHgE4MqZTn64XTkY/FYrtfXT0hXqE0/TwZiENl6NPUIKG38
oYFWYZQy+iX0PjAAJpIbnSJ4fHuNZIoRU6VS/YUV0cYUx52DLifl1ymwFBUhkWCm
vAWRvaeVlBZF4Lb2DAmCYaLr694fJKwuH/BXrGwXG4h+BDURXApd6bpLvaTTBHqv
nbF4vChkcHpEdtpERQocku/wJxI53ZNsSr+O1EEfaQcs+btGuxGN8GQHEylmlIS9
VMnxjm0TzXg/XhQRfhruIXP1T8PqndUxcMJ4xYFPDpc6wT/MjkRbMk0c6iQInecN
tj0EqqzdvsqZJbzS9SeDVLIWe3dZtxbBXucIH9NuMixyx7zG4NvxvFAd8XwHgoC8
FdDXuq163AxXEacZQeGuU9ZuhMWGyoIJyYzWLATHWy55WW9dNUUlej4iVTxheEwU
7kBa4VkhDu5SMULA29nVzvkbuWMQjVIdRrB6DvxlFH1xXUc1aG5lQDrxoRtM91xt
u3HImtVYRjxj6HDUbQbSx2IlBkU1d5i2v5ybgHBDfXvpVAlWwYj2wlq1krRm1w6z
TpyM678Uuo4kMl9NgvjsS4BXR0AAdvaLwmNC6b/NFESVkJRgZ8VK7/R6cmg1GlJL
JCDLadYJu5Pss7NAp39o2MTzdrr51HraEa3kpuJI1fmAfBnNt/X0l4kWhEUhtyDp
i48W+6Hvt2AMPnuNv8dlOrG4rsYuYssq224rxDxVVHJ8bmmpic5yikyrFIsgzd6p
eWU/Hco/2rLqLpxzev2uAgo03hLoebSzlqZY5Ief2ZXDW8ZucRopK+nxvqOFnYRu
gMwJLyaf2nRbCYXf61Y0Su54e7tg68sNWclTaG71mN7wxJ91/OPikh/ooM7KdenF
Ue13JyXY3t6S2U4zp1ovn/qJ/HGB1FRyGvS2VY+hbxdl2Pw5FDnHJMnWYkYOD8i5
Jx0VbUnISwoNT9vgwkJbPlDbwObU2ezx7eqKh+azSwRGT0+KQt4pTvgSf00ejRv2
AkBgGwsFmAIi9kfeVyv2DwEJNHqACY/Uww/lKRS2kQ0+OME8Jrm6eCU0ERPBg86B
iCS/CcKiWZe7RTx0jtvCTiQjN9Gh0u9l/1Y+sTRICssiHwPBrAAXsgH0KYDVUm1J
GQI88gOFe2Nk3k5fSGWTDrKLeY7q60JugY0b8GyEgR7RIpudcpXQPnRArTM63fz8
WBJaYpsixxscb6GtMMZv+0UVTDxSHgdnVH54jc7VD7DgwrvmC/vFh6M7+4beUeJM
bk0YpOOLXju0fAytbnWtlwZ9JalyjcRSQ9zwfMesYy44WPNDcnCYsUkZgGTjd9OE
qaNtNY6oVxqywkLY3MxgFZymhJwwZgKo00lNRuHKxFdOUBxNdFEQeLPTNIFpwKLv
ayO5hLHHam7jMnv0/asTHsJ62KJWXP8XNhHQtBQqaelDLUNpEYhOetU06l1ZbieX
uy3y3RLcFY7KdcT1PQdF7Niqkz/3UxYbd4FT4Fj820QxFfEKjfqWvVYemZ7WbMe6
3NeSoy1L6STW7h3nTwLBroscJYIYufcNVJ6GihA5xMO4dbpXA0RgHZt0Pv5cJGkh
E2azuFVr4bK4bCDOqOuAPsnKvAlK+RfCg7hzF7x5bVMeUjoloc9bP1LYhxbjIURz
4/NkYRRbqUfzQr5q38OqHRrPlhXib76AunEpC5hAaRlyQV8YKJ7cauewUCaDAUJu
8pfzqVt+QkZJlk+rUDyXdJM73eFnQpl4CUrAtMiASohR6ym94NcF9GHmcxJMa9aN
qUGFp8dZYrX7RwG46KZmjue7gAaEekHx608Rpzu9G+9ri7UUnkOMnQH2q4CLFD3C
T+crI3HlZqy2YRRsnDc/JbzrAiywKWplyO8ZYuD6vmYeSz3bhaR1/5+SVfHvKXYn
NLNVi++kQYzV65+AjBTwY70+PW9adKjU7LTg3tdeCGnVIStrt2JqY088cdjK6g4A
ewx2TpwLIhJa1dBS2Hsba2yQjnzFx2bzDk+rhThr66BeBk2v1jdX9AyjEEWUchyB
cBSq/dYApidCNnMwKYlZ2tCz/Fo79WYl2rmwuLCKwnoqoiNZedpuCsSEYC5BlCCG
I30ufzkQe02373ye9JZhMPCt9jqlD4cTXEZ5vKW+7XhMP8TriQVsxJkZG78evvVa
nxkhEgw7u9JP+xKfBmaKWApoOhyzdhV7On1tNB0A1WAiHaC/HkccdLrZqCTTO2uI
tMrWW3DlRfLG1byKPSOkCscjWQLH6NVm8WpgfEx9uJqGGapejs9S2MiXnRwVmLtx
bryv3anMsX9HNzgpTzR8K5tC4s6Qaad4fL5hCjKj9kh3vDDRtZo1QhXMdQlqkeSb
G6ZxVLUb0mBfPyXZF8dNCJy9mr46PwcLd1L4mVKAMOypcwx2GD4S2prz0kFlD/18
J6xNFcUKpSrQOMRgDFUgUbJicio5IJsBTE8hgWvmpROl3PJrcKQ8NODr76Cs/NgV
Y30dA7+J15xZ0ODTVEMDZSg+0Wl9wTHzBB99h2eeIpMvwEbu19G2Apxm99/djyyA
UciLdtk4iEghzZyChzcrlIQSNWYgK1ljH8MAFiXRtPz527VvC16l6/VHvWih8WGr
xtJJ/mJkUZKbVd/vDzQ6hbRsDWduEDAxTUunKJTOEo5XEzovSFCNDJzKcEsqxjv5
d+yZCBavY00QqetLM6d1KLyxvMZ21Mq+iXyMSEQpKwcMkvo6yD5Gz3QTqs+YcqSH
iIhrrlOwkcF921yVFRUhAYPpG9+5wXgID6ZXbm3Kt0xGlij6AiDEyqCYFprDfg2N
N5uyQSVbf0bkZ4SFVxJ1BMbO69RPO72xx3M2Mv3OGGsSYScmADUSsX5YPbWWWgt7
X2gkMcVKFpx+CKHnparKtg7iGIT6YIVvUl8Zs4F9oGuCKjuk77r/OUyurhp6SnPW
Q6qUAOJlirao8Eu/nLkkr9nBsiw+ZcdLZdczOeY8o7xfEQLwoLfuP/gSLkIdvqyt
LSbM0ehcl1CwqNdlPkZ+GbUp+kUvptkqJjn+VZQJT1WFMyeSefuH/Dksca6FRDuL
pWUycc4q3I9tUKIJYIfbsJHL3j7Kqnaupbz2x4yqdFUDYlgUchIPv/QNRwMDTKe1
kRamTF9z+6ZSDp6U/tzvG8syuMsbSESEnP+Dz3T//b6711MCmon8B/02kxnbgdMa
fEuJw14dL+94M2aKcAI3rkGaDMYgIym3DPdI/hl3WAaxq/GZFTBchZzJOcWQK4bk
2428jyGYXmu5fq4FWlLFTBsAedISStHmkbKPmSd2kEq1FBA2Ru4FLaMxvsgR4w/a
grrvi7Z9uN427mWuxiyo5fGJJ7+8p61L5poNNJxwPo4KwTudbkYMx1BT5hypr94w
6pfDyNAVzK0rDwHAbbs6bOh7yLU3vH0bBUx35Fwc3htMoJYbbI/ng28EAJZGClM3
0GuY9fn1wEKARnpn/nkCsxFr+J+vVW8RJ53XCDdY2+5ZrxqHTQoF7oPVv81VJ0n7
2CNcrbxfUgJJanPN0As3NIRugi9tCUBHqcvk16c6TjBZn5UfDRbRN5+mb/UxZLUu
9wJYi2A4AXeUXobbRplTWzSZyCqlGcHaSEgVXFYAoOpqArNGcAVoJNkvwq4j8hiB
JS+p5nohEuSYnXskEilwYux5hkcJ6trqi9cc0QPv8ajl6CFmw0xmoKSOoxp3UZQX
r1IqMjstpXOZ6vyK0SuugeEv4GIDOBKH/TZVwCy9DMxmnR+u+m58JHEH64helcR9
gtxvy6Pj0msulOfqq4KmMihSERWuz0eYqA4wLYooPdAbW4NsGL+qYqfx1teUVjus
vHdcXRxNEmGgnJfncKJZihnBbrlMxNLTiajmwdKyXWpsoegzfh5SvgdVwaIlDfPQ
XXVF7AYQy20iL04tTKH8COPFH1/Z9ed06mb0ZGhKchJOoU2o1b0kJbzeVlCrVg6x
DrC5cSmxhhE4UL5X8yfhUWjnIZoivSCh5KhsRj8euCpYBBXIPJ+rUXhArgXBmm73
QzBV7QW6UvZt5QpK9/9hnxnQ+GQPj2wLVIwfTDvjebm4fhvxPfu07ts7B3YEEDNa
98vidU5gmyT4jvjKxuOGoGhF8mPym8OjhrGzcdve2y5Och0ajO+FwU9JCjaC2nEG
pEye8Kd8xN/+Y6KF9/n0wAWj9LFQvbnda//MvZCQbmjoovSWUSi/pFmQfQLs7NHT
hvaxDA8wSkYUBzz8ujkX5hGPTLFSPwrSmsfneB5HyoRYye64yhzFT5SsZoeJe3e6
raDlGK0otjSRlT8Fw6eSifeBznQEMS2jWtI2BmtgybxTn1ty81AyvhTYWmY4LiVr
YkuuiX+v10UkpI2pAAUwCl+EVX8h9R4nufVcwZSZkryrjtHhBqveCTFDdDxMAXjv
u9tqDy3IzvU6Yo1wJsTAn+t/eqfZ/Pxa4pZ3Fcm6P8myj1XODX04T/Ldi0Zz61cp
9eMDHTyg5wRmuDGJ9jGc/FQka50lpx68wUE5SPIZqp2AdNUyHEhbu0n+PdWXbm2s
1MajMRzVfhB/UWEqCL248Wv4s90Td9zffKbi/W1HiMltPrFScjX1mgHnZsZzIkqD
fv1wp2bnbX9RZ0CM5KM5NY8EeJREZwwT/tk9OQjv//U+rXMNlI7DBtD+CuUxUFj4
nL3wNTPiXfFQmxhQnDnE+kKnTMYM8H+SyViVAXSge8owvEAF8yvTFQ7Q4GCoyIl2
xqBOq5QPluI5Z6guc+a4oKRapAitV3QA2oZgQuWzcH0j+S3G303RfwtGrrADTKwa
zA2nUCrBTGzYwnxe4KK8KUnGGD2f4o/x2IEsn3WJwbWVxhEvnr4ORHjVJGK+Qxxb
zcReovhdtgPt0zrF+Klfpiu/tYV1lgvuOq1RGxeBxz4/xPDtaY0Su6QU95Tavs6G
CvSrnQt1zg8bxeRBElfj9Ec9jZFqwS6IE0xGzF/vsafARYXL0Cup3fmr8DvJRxr3
gYWWsWwcyAQq7YmEDSmQVZhV6CCB60mNq8kVLlaI/L+cOdsdCEd7YzTuPamXAoDb
6h4udxc5yZkDrQZYfs/nd6n+gLOAYIIH0AxH4CnsEPPnTL50ck9240Cyw5bcXgUh
VG/fzpOQbRlab+KKaCUZb4hJrtv8f6HAr/9k7bWBR7qJjPLjGL277B/zL6hzH+Yr
cU6G6IYP9eY+PjS9hQqmQcQTq524h/SKRqH6fGBsspMYcoIgCJg4WdhyUTP6Kw7W
/nXIQSPlMDm/Z5QbilaAI8KsVpwpcYQ9q9wtynVfaX7fk+2ZF6JgJ5Z7dSRllmbV
BmYZIt7DgCIulwGHH3hJF0UFFjL8LnyYREdirZnrv7TsQmAB/6itSytqOhgjLvms
eb6DqD7aEdASRZNEWCd+nhOUbFNpewwVRbwTligWQEBwOHaloXWyAYs8o2Vhi/tq
KrvvPJ0ygZc7wwFnNnwJRtHYqzeG8WODvYhSVr2xgLI6dbHsp/2zmablh4ljRKGy
+HiVGAqsYLYOeHb2VohC6bmLlxyXFPlz7rXcAogkTNpNoPkr9Sdl1HR50Y/vU6RL
g+ij+D8GEmz8CZdvtbzp8Iv3I9QFF7/umRZT6W46Tg2D7knB6BLF9zjzahLYsxLa
861C5BqLKvnZBWwf85VisQdgVp99FXXr4QHcPbVPHulwhqHcv2Yv82t5AtGHE7dV
I9Kg07lhJyvQTBi/pd/70VosJlm/Pl0WeHesTUN+E6Us/Zv6YBIAKRLGIuWwuNab
q9DNNAl8tD+QzobmKDcHYKeonqjWFEI6AM2prWz1MBe+ETAywrjxR7wUwuW0cHSP
YjhdgT84yDriV9n0nkkTCDwx+9ufU+yij74yOj984i9MOSKH9fvj9N7d9+e/+xdX
YP3aYu2kyeATB4Co5ib4tXXKCHEf2GajYFMJ5pRC70IjdmNhdS6eVPCNGiah5cFD
pVJlZHtXpRZD5gjIt3FxRP75QgFqOqKmfyhSkGUSkq5uhQPp3pW32y/ctEz0sF4H
3N1Oo9g66tYLqibCaoQVqrpl3si73tzAH5W6EANDGKcoijWhy6Cp/Rep7wy2FC8/
zlW3AVmw5GvUyeBFCupNPbO6jk0SDTDN7pJpnwqTfEVDbtV+niBNwutYcALgICwu
a6IGxgUkBDrFdxkYE3cuQet8FPHPQjhVLyhEl7UBIVfTZh7Y1CSZY9wmoeOS+aIc
j1AayJ06ohIPk+FdTuYdFNFm7wPwQmDuqjL5hoAJbSivzzdUl8CYdWk/fXdFPSAY
N0ERLBH7+P2RC/IASdit9OBvDzJtMSKNYmIaOAB2w6B6XMylfNJnrD51Dq6Zntq9
qAISpSY7eH/whancSJsZ6FO9a5seQHI2XyFS8mqI1tBU8D5iYFoI1aWJ1XJVp6Wb
C4HVLVUwZex/KD2CT1fVpjLGXKb3qWTr9mB72sRIEuQNV/PjkkRTvELc1KNF21V6
vWWUvWKcT5e208C6bf+kujArsdXgCtLeQ579gm4FBtcbBG5yIXVioCmLyqjpZgy+
DHr9YCxK0hGRIXmQ/gxSHGAzws4Rr/mO68FJuh72Y1g1sBOefPxGehxBbUBkvk5a
kB4MmCMNhRsC+Nk5JUXKDKFug6t6jo4JZHEOdRuGmo+X1Pcz475/OafPvS8N6DGD
/ZdXu/5hVdN0c9EjL4zsCuRsefnz+Rt9JmVNVkXI+4MEYU8cNHwsnXr7RXY9gOBE
TqF2CdYlbbq+FgTLYR5cD44WrcerBCe7HlGnEfCdU9QO8kdPPBOqHPI45UVNCtSv
VJ2d4+bG57SpVJDOrpq1uR6GsufZ9Z4eMAqbav/S1UKEjvUV0kyGsUp6+ArgaOru
vbWQqOVa426AJwSP6rFAtfXiXCtRqtuofJidmyLgKIc=
`protect END_PROTECTED
