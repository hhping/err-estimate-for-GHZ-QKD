`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v/SxY5rc6VWkgCkW3hnuLSAdlPbBAfU8fQL1MMcBPjP8Kp2oCvmkKglteCeg3k41
ObDNZsBPBq7Zq9YpLBPlHKVLL27HbahTfap8QTAm+IYaGBe/3YtbMNs8j9ZOr5Fj
Q5p12pIvwap+v1kietQQcvVU5QJy3XFqLFVT9SMfOXOa4YI2YXWjwfjKsehI/qKk
y2dHCla0IxxkwiFvSi9BI9ywMW4JY1CrdHsYyXu/hD3ENn7MWMm47vYMcNda49D6
vs/QNmcQw5PhPYH84F1NO3GlGfKxHhSQdmKYAhBWzZEjl0uBgnfk0rYpT2JSvVwK
UvwJKUGPNRu26kcVpUypbgg9okrRRkYGRUmLZWJg02TbUWuxMrTzitDc5jcifLMR
32pYyxWeUBRN5TkFomGVDkN1Uk/aUMlEvmRYi8bz1++JS5Ox5l6C1RdUXlTQIgLp
j1HJTULHXUQIDLmGsK6BkYQm1XYWbcKed6zs9rOBJj5Dsnh32ZvhaXC9GwHnJAHD
G6jd1qHQkjpC9aHd7rwffBK+7ZF9dGrQylQgRf9Tt9U1C1hGv4RNA4mKzD+CkuVN
WJu5/heKutCIEBsSUvyrOUdvfwbFuzpg551P7aePux2H05geOJAMGDTZcWmR9Gca
ypdCpuC8i9oolTz/03F2Kg==
`protect END_PROTECTED
