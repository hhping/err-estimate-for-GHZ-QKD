`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOb1L74IR2xQERInf3n4gj7S/M9c0ch8voCUWokdXqURsCbxskwQt5Hu1uHKYkVo
yGqy+AueVJ8Kol9qtOGAhLjnBZ39udXifV0lBP3rGi0M1hqO7CW4So45sOBSV5e1
ajscNACo27hN4F11nxkkG2U/1qo+y/DYldaPyBbe8yRen6Q1Y6YUxC7qvLwRGY4q
/F0s8tWfJJFmU1mEx8d6bOH89F8+gL4lnquoD11IReKDMcpjvcnXkKkJxbF09SSD
jxRMUf29ZKoDr4XEG6aocfKy+HnNV10IFP4PfrVMEdLNtc1ef9Yiz5+7oQt00Doy
KXass/3AcXozWETYLJ0xtYZfCy4jiykvlcCXcMHCuPsDq8YorB5y0DuzOq9F/tT0
kJ0Z6L2GIIKm8wNWnjVyIZHoZRqtHYFK5A2ixcefYQB0j2VHglwDTrU5s6ps5EfP
zDZM8AVBMM10h7kYBWa80COBdyufdriD06yYo3Zzs8w5hwn6KEQpKeIFq6pGJK54
lxDwRnDljC8RE1KdofS7EBrthfbInGqNY6o1BTe7p/th73dM8oKrX3jTKWZ7noIX
IhCK9mBYTRH5Vu55TLykUjKbpv9hyeH/v64hgI5TLKsE2uqkgV3tkeTBiKoBQnnO
uvYzIyVFIBg9qJakXEY3N9dh7A8UesYl5xV+Z/fx7JuBnHzS6QHyKojiBMGifky0
idC+vItX0K2Y1PUBb2wV28G0bR0wHJW3t1uB/tBxEzHvUXd32TcN8E2F8eKgfYES
iuRk6DrwCGsd4i66ytaNKrglMqrzV6HQvj18HKO5sb41upN51XmLMunlviZ6/mNf
tQOwDXLYikB0kAakpzNX7tQvfcYGO3Y4HLClxzW4UeCsWsBuU0OqJWnJbCffKoJN
FpaBjMMmJ2PFl+AHL5Ie1ccHmFK3F5t9EikNGIqlkhHRdHXqQr2Gj7irnR6qypQb
`protect END_PROTECTED
