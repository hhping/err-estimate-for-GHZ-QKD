`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iTNhlWxiAyZIJgmn2ajHnbTouIt+8X9ggroEnxs2KDN99XAyetNfJWXNULhobMD5
MC677iuHgfEJMqUpzk0e9dQcL14WO7PB93vAU5hoqxM3xJKcHrG+wUe62WJXtx7I
bihEjc5tWkahhWMlan8rBr/Aj6QE68UgpoHc41fds/eyhEw8uMxkqjCD/Z/vLnNA
Ik4EvpmI6QWkPIfoFLjiq+OhbUnRwcwDm07xb1CIb0Tojdk2CSjD/iuSMl+agw3B
WOdFBCJZURbGPwLQVKcJp5cRByf4oOzdw7rUiRywaGWRpMNsQvdLIfMgF1GJSoyW
05o0b/W94xisJ7/stXgWG7x2pLfs+rm0AVfk9NIrBPVGWxofqTs4yytCBH5xyctq
A0kyk65r72Po2T0vxJkOimLGOrM6XGvuynoE4DlVlsm/BPL95B+0sTTeGJ1tl8Dk
flrAhkGXdzb/pj3ubU0KGjDlfetGmqHkM9/Y/pIQWP14D9R5o5/o6XuIWZHuP+L5
rZB+ub9RoMhHjtdBt0TtsZUARmXfci+gMfxatLZNRg8WiR0wcG5G9YMMHeCVJat0
+nj9Ufp1Kxe8zfw9cVk70Ro3KYSpxGFN0nAM5j+vseXXzMfAH+Ig2QWUIGPdM9uT
hqaxPCpgOv2n2NffjvFtuI85Cl8mPxu1ADCVIAgb9NxTWSic1koYWx6M78pMSNQG
g+KYoSPXN1e9Mh2Hq5sFtE7RKCAGVAl1IlTx9l5zDw7ow2gRpXT1pmx0ZEhDr507
8K7EX4joyPHCdz3ylvaJyNA2aMaPWEoFN22rtLwfcEJ8mj8sof11MwQq/qC3hne6
bYb1v4YffjKl0BA8ZdWu0IH3lT/kfOk7i1clvWePhrpTFX4ozQAblpK80BgLQxqx
uVFfRMsfqhyKWNbOUkEoNXGRJQIP9aLOstz1D9hZLSOgSUOZBsiTh3fHSklyJq0W
uqoYpJRc6HiFKUY2IZhnKM+sEh6KLpNiR74XDLJ1U781cZODqHyIoWUQvBApFBtb
m+pOuTw9cFxzqR5t+qYux7Zstypf3XMgF9Wig/MsxSpvfHQk8Ez3KbZs6D8/q4io
BKy5nf02iTMdt6KARaM/6eX4mbagn9pQDKnboF/mx8+RomRkWtCoWwlZcvZ/Yj12
vhgWBTt0zUs+g4ork2ATImRRUSvniy8aPXOxI31NUZOzZkR8kPHQxQGMuwWICl0l
iiUIPt32iN8GmNDGMwwjnZ8E0L3qzCN6p3PIxsFIUReWrdLH4p3crE/W2cGN3Bp7
1XdnGjabxCPygHrBAPhxhDOfwm6n8XuCAwB3TbD6zhuGQ2bE0RrFpD4d73tHmtu1
VB3gDYFFQSfSBl8WD3KxF7tkd3fYrq7Jl0dDSxqtMLfH78wyx9dcO16wHtGos4BZ
7UjgnO2D0orUeaj7eJCVNCTDInZyZ8E9EK5R+gs+Qo6hO4QgeVtgw6gqXm7+YSew
nqqtMYFrmji2mgmir4d13Zn6+DT7Dot6Ir1Vmiyuh5ookS0Kv788WnzplyLYThRM
2Sln35hiAfDo7lAN9rRcHCIuITZZ5xsh8iMkBeV7W7GeNZLNYWxEnOvtJoG/Iedv
AxDQcLz6J7ckb7QKHXKhFr5XfK6gHH1QBUnK2SL0Yd1gVtY7rihRJCLA2Z6Rp4ou
BNixk8MFseXhLUgrfQRx0PaWuknYL0cNeFobsRnlZkjvs1pFC510SSeuVRpxnYEQ
Czx4zYa2YTdidtOfcAG+O5vfjKoGjn9FSCi8sesAt9U/nRnsAa4mgzTTVIVQEdJj
+IgnWJWWsEyDmdh3HqsEC3V9mCHO0d1rM2kVq8HvoBRxV1NNq4G/Uly/h+pkr4GP
BCOG+UibInNqk06ItJlOlX2wMS2kKmj0ZsAracqL4ZUZAofWtR47158C3SzgTw1N
0BslyaFVVxYvJzGK8D0+KLre1uBl9SrvrAuQFQY0XNum3t4pevsNJXgFgIJ1Xo0p
XLeSAwfHl5pBgPVN5EuqfIzZa1hJHXb0mDjBD2MjtG/XXNjbxgRPN6Fzakq/aciZ
Fp+Sdv7SfRErMfJWjZZ3RfDEzOMG3tSKgQnHYURijsD3BW98T4rWzeZ08icKv40D
o5mTkPeFsvlFH/iy5V4pgBhhyl0HGXknYRGJn8I+4kH78B1WhmdUw425T+kePoNW
ltWqnU3c1tn/2ghrnsYQOewlnULOBqBZkTmyT+N+hL66C5LpcvxRFOqr0fQwJJF2
0KZKoKO+ar7lCfnjPqII1j6yklGn5igUgt3SxfXIELw/zcH1joesgTAcnMXn/nPC
BJsSCbFldlxrsZxOGz+nXT1LQp4vhzkTgayWVxgC+FQDWDdveOywGEI1crO+8Zuo
JiIUJsbELmWYnsdnpj76VD8zowSNpwfOEPJ/dM4hcCHJaPHCu2dPawLwCG0/dQnB
NU0/1LZlCImjleVH5Z+25/li7CVjkwAVj+r+Cv/FrTwmoMiP3JCdhW0HpK+ou9fR
jE1gr1AMPeH66IO/lwFovRbQqxGSC246S9HlRVN4i2Bk+DRkoZds5EgO3rUEyqCy
eXtXGGCAtfFB0ATmLWs7+J+Zu6eW4DE5D1/LGYqKDO5tkCVRhSeD5xoowahzSA+h
crhA28oOxdn7MUrih6LvszkF9ja3C6OLxRkH2v2DY20+0wNheh7DgHiDDVSqbjnK
o6aA69dvMX1ctsPdmzlBtdjKrtmJ22aLUUQPLEXMEWNp3W8bsi5gR9NAXSozGXK8
xntCtl51QgV7uQsbFEv/9uC/I6w+sjvUio0Map6tVXyhHoaJaSbi90BsWpclSDZV
JcE+QASvkh7+SDxT39JX1BQUI7naLeliwTmau3MTihgADZTII0fjtT+cuuQXPs31
OUW/6BTOCy8CAw9PFWiUpEE3YziaNpN2joSbpcqcxZOJg69UiDwUqfgPO8aUnmMM
yjEnpiy8qPBKOB/PL3cGLN64ZqWtyokELpCHM35n1jSDAmkYIjWjpKGqs3iIeIIu
ZdkPMg3e9pIrMDSntcJT0Q+WsMfbKImvnxEi1uxOYTevNSbeLmfwDakHqg7zuraQ
QGX1GWMTr4cbjyaNlMqsaqEJc72+L3ppx0tYoSRi+60=
`protect END_PROTECTED
