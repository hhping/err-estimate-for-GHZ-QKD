`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ALYSZSW9gcKYHp/7ia0ZPFHottr4zygUMxOEW2hgtS68JhfH60pqAcdROxXcMD5Z
nOxXBFd1j1OwJsKyUyZE21oSKMpg3pa09x0NJJ17nUHgH/ealLyKi1Ur4rYWXLn4
5AJPcBDB2NdqVTgkyNXlkNz1+rpDuPrTtp9bEbJKizVsaJKp6HckBLBfvj4PwxyK
adI3jCSp6kBOnKSHoh9o9bOOZOGIhhU9ENkOYEqofrPDrmH9OmPtVa6JG4qog627
Z57rPvFpSvHSTqV/uJt9ydaeqZtniKt3Ekzph/X4q/Zim+2JF6+CO9FV98ayHNWq
dqRTo0k58k/T35/B1SjR3aBTVUSXuOBciWsRPlDCm2gVq8YxXvrALiCNlIFg01vd
+cTO7Xz4anBL/lQeBy/V2nEE84Nq/6rR3T5mbFqJZCUmWJRvL43sDHZC8PKvUBf2
X0om6+0jjdZacNguNkRMVCyXQRfUmyIYE6qhh8nNtGakrJuj/bIp2BGmawAtq9t6
KuEjKSFzISmVoWqXZLxHyXUcNyqRjqInRKBbQanNmGdRUcXX0oGmRApIpRGwXh4C
vxaRaCfOxViKHQg9ObKmlRQfBDHr3PsTG94WjlLleN9ZQMxvU27h5noOSC2oT0/W
uf9imGen5Y8f4hnwRZ4/Es9tmeM1W3OAMIJfF1D8QsE=
`protect END_PROTECTED
