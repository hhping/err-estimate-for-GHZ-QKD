`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IuWHpja97hbAMIsXcNqCqCGOmwltrX2QDike4JKOL9spTftdBIOKZIX0LTqlgUb5
9I9ftQQ35gL++UR8vc10Sepg6aHEJwdLRpVpniJFZToCqndOXPKZEYZnNy/dIEiR
0XDsmfe8OEs1ZTgDGDmS4KKp1j7wsV5PVdeKkUBAyoqI2K0kpLbOSKpF6on5ghMh
z30Y/XWsbypM3HNFm684l2ds8W8NllJOfCeY3+a+q9QLsDWEUorZJukLZOqUyu4o
S9O9BU8naibBsHJr0RjWNuyuaOQBpNMTTGVfiZEkbK5OJbccIfZXAq4hVZPGDYzj
Ftb6JQV8MOpRnb1AhaC11ndxbUNd8G3F7DzhP6A4mc7qXDHCvSUiNRBBaIcM0m4u
ssdvTJgaBIAdPDy7cuD5OriFT9g6TYMEtUsgL/097fbvvDIUtpcFpvmsRhXzkuCM
2DEI8RBDWmnuDXTpVGAyU5CIGfYVRlOSNWO1kWRLiZLd9q5OW+0dWP30drq3IW5e
1kNzSfDOpvOVXvmKESKeltf1h8O8t/N/DfBCsR6yYpBBHIKQ2sYSXMRCxuTz6Nmj
+nlt/zMwB3XhklykbMvCEUOSiEIfdn2orY3zdcIK3ul/nwrhAUqem59BZwqTVnwC
+jSJH7CU9Vs/svcv0KTSinj8vrngyVJfmDG+A0xg6gKDafWFAsOqH+5cmn5IsFfG
I5HTrO+yDek3ruKtMTIx2Z1FkZ+QEi5ww8tD05j+CPyarTH1X4630ftmQ+Nl8pVx
cmJr4zs1xcPl+asHvi+YPjIJ/IIGFE50f1O0bKcv9yVHVQ0u2lbdJX0I5Y8TMxev
s8YzEBr62Ot6yHWvPdMDzSYAB1W1zfzkYI+czjx6PgC9BlgoX1lVcUy2bsfHmbz4
HlEnxTHdrK0QA8ISXAHFphtDkQn3/eAwZWcbwAFk2tqL1vmPW8TeWQOj/k/Pv7Pw
Y8Quw717VUS2Jh2Py3o81XvXEI5zfod9RZKM9ymze0L4ev60SjHUfclbww/xMk3m
efEDScmVWuMnXzan6OsWo1fZjyo2n2KniIsOW+2IMU9Wz4vfxChUQ3g1YVPBIOlO
c9BsKZU4DdRAZdTwQlwmih2K1gL+K44jvp3wo1kHy+bhOgcJDl/p34YWvMc7VEZs
Z4KQLR/m3Z29gtnTM37sk/vpELfuatqU0G49K5P41vb0BuGwmuJ5tVlxlLuO84Rn
OiUaDvvvng2BqXsHxGJlmBX0GmZlld8JFOcqC2InznVI4Cr83Z/9VSpWOLHoLJRu
i8dgFLLSXC4JsraNaObkhVQRrsfwuDgNSGSpLfwq/k0EJlK4c+sNGErH+BYS4doc
b25P+BSHzFyeMsMOPZXBaFyqEBORXJHVFW+1lvnm5vME+HEoaY01aKdmL4WPr5dS
AOdVzAHuEtk/xlmuVIuU7kkldLjv5+s3EB+ZdYtnhXaXcKwZCn/G1wJXP7HoKJxi
5quMX+y1ntIq/FBPRuhW4ahajFmdBCD7AAIaJUc78sMnd4ji5W4AWMW/XquCKFqh
wHJyOgDJM3rX2XA3f3bUHIyL9VJcowP/CwbgqmxvQP+V2wcANPCiFJn5/Ssq+YuM
CYL5iHLu/4xdnoB+ypUvHNkEHYJHGVy2XwyoseH6F21feVr920PODKk0kQx905sJ
vE1+hGd35tf5pSiPTGEYn1QHR9t+YBOe/vB/AeMGbEUQnrWYQ04k/glG4SRInR4I
5yol4Qlb4FpfmdncjwWeO0MKxjp+/WMGAD1kuO1TcisjYtusa+3VoxjcIAVGHxn9
DfVIv/urpIApLwshFRFehA30y62esJzRxmYlXI18LRSAgQH6K37fzoXU68xFDJih
+QjxiXErmEg/z2g6BOFl3v8r16ai5xhP8wQF21kVAc25IKHGB3s5htl1EqQTY5Rb
q20wGEHG0olXI1PRE43OkD64bVlaRUIXgvdivPeT5Hl7AAib8c0SxSA9DTPu3B5D
VFSV8FJDzYPwmwG49e2T8D3QOW4Jp4YyDiqVwV9IiZrXw7VQQfao5gchw5IlYznL
Jv7QYYQOuPdsvq3JFbusuiAgKUQw4rmLdqnwv0uu1Cl/Ob+p8Pcu/U9IMofdCp2L
EyGVo6PyRlj1L0gxjK1vqtvQD7xpI5UeAKoUc1TTSxJi1sBpDOB5hw4imIxaxbr0
LNERKE6z9KeWAh9YZcKdgCYfINb62pQnFFOkWkLP9Bt8dvKWE6XzP9skuoiAgyGK
6SmdZQ8zsAJcZxUJGS2mGg4GT/KuA6JPXfD26ITJUdmCdvHuFerS7NL3VYAXsLXR
p6pBFwgemoEpSYn/HM/HX07LbK+poNB/ilwBeXTC2DE6B2JGzs+XEqumNE6FSHXH
+pK4Hio/9SyTHA9s7ClMwyoNDHcIkf2oFWw2mETt5ccS3GOWdOGqL/irb70bSIbs
j7Z0h4tND9Fu7oQgGADyMaJTn7ov+SoGzyTq87EYPAm2vljqivqppNyOA0S1svIz
yjoolzgVqoDobcuwu7I3pkcNgX/o+nj7E9EFdzIT/B72sGazJIeLsIAZ/aH2XLz5
pOocvxji0zR8/K6pYZ4cUM3AFl13syodFuQbP0AFi0d21dttKiaWpXfIZDG14QR3
w1VknvP7UQ2OfiZfjglN22Jua67QRJi1x6SIuqVyfFEA48r3JfOBWoGnIOujgBiu
iGbGCK93wHIa4OUP+BQ3IMOT9s0Wy4np2aHtrxWkdEhvtDX8iZHUQcLnbW4BOq/u
W0QS4B8xMjVHW0aHaSf4wjyFJWef2kRLFpraroFrUNJVuEYIpEXpfmbiymIBLb5g
htuUq1GsEhkeRpXOktDdVMXOCRC05BrMDCnR9PYMsLzy36nO2cz0GPsZd7f5OOSd
eMkBM471tiy3aRh5tz7/FTSuvGVjxy30RGgbUzjQopNlaoIP3HQHjmu3VPfHGu6E
C1C+gjHGHHTcEcJ5urEp0PmW4lCxIyxdt03YZAFkS1Sb4xP1U0gb+ObIkMQvz3it
EYEHL5njdwsWTXgNBXPM7T4WFB1Apuwzm5r16ZDvVOxZXRp7erFJyZ1Iiku/Avpx
ulKeKaEZZLsZS6PgQAQHY+KRVV2s6ngRtL0utWPtNoejsgIU5r8UZ3yMbskPjuTL
2E2XSSotq5WM3h3PvdYsulPrBquoYVHXwXaw7LAABymAYBU94XuXYEFONh/s5ZCy
pbYrLVFYOBLlRoLXc8sCEU3U8GWiB2lLMCMSShgMJzLOqmOF6CF+otEPUpvAhna3
JgoHKu2GLdOUFst0uV+yhH3QWhGJEJ82EJs9cgSliy9KAJLs/gQLYPJT44DiM/qx
zmVriWC1dqOnlO+2g2Kaezs223PvWw/67wN/SuzDsFYW0FK5bQp5s0IBV//xBzhE
3RURpZIzZYjTtnWel5gYW44IlWoPwSyHo7+8hqYghF7dMHb5qQjFST7bkNfStlJp
b8BFD4NdpVvykSQmHy4TSUBTsis/t3zqhgGsWVaeVB0hKSDA42av+vyqV2VrDUQ3
xxrgLoGYFxvPdygRFlfS/A+FYVa0noiNYkmVncD3U0KjeUdia4SqLePJ+HVfgoNa
PA3TYw4s2zQ/K+d9T6rPLweX/v30Pv3CkollO9i9LxlCktmc9ndp+cmFOiEn/c56
fSRSaexnLfhXxWGKnoSZlNJVHwjZT/V9s7i+SSnlVPsOfUIV07vNw1iuvsroQB7Y
V2JjXME/x50YD940tv0Kq/Y+/H8kaxNv/ac/pKlgmqsfjfQeM9XxIeKk0DNDJqgZ
OOJwBVPmf6Uc0ia583TjPNpKwVraZFKYfy2yGGkGyZHTiUEt5IEAzVQPxT2lner8
EUe3ZQFLfC/8jM5/02psJM1xonbItR9bilVZKLHb8RCAv2ABIebsE1p+LG+PwpoW
FWgok5kJ7+sURGM4GAw9SXQbe5UYIXciOpSoWhffnkDZfLfP1pDuQhsqH0TkcWQl
rolZxLLXRCriYtnX/kqinNSqonIgBGsdFPxq6T9DkaKPfpEmeMWS7How6nxFmk2F
Ks2roLRmlu70fCoYwvC8kkqa/Am7IE1coacKejelwXlMy8hB3rEAtxgdKsPyqMvT
3OefS5EDdGF6veh7RZsoI62efZWMX4nvL6hwaM2KVqV8EnvWgQ/wqrQ272Jsrmtb
P1+fUYYzwu5dBUOeetaCY9a5pM5aHyfJRMN1IUjg2QCPkLlnkkItz0e1nJb8sZLV
1wQAGDzz9U2kWGTZ/CzpNRYuj4HTY7mghHMXlqLUBa587iUFGfhDDPjZXxzLpVQm
ZByunmfi++EqUOXMfmzFhgYmQf6F1bqD4QzEIQ//peMgTKrm/cgAjpDDRzq438lh
SUDX9o4IsjwEJDKYI8U2hpJw1aEHA6Oa0Ds74BifsC0lGfYeHBkOdGw/RQPc1AIa
JPlgP1N+E02+3IqaPDl3Tw3O9gd3wZZ/7K4I8cfnq2rlvSPDFJLEXSRifdyii7Ki
sbCYF+yNoOLQj1OIBCBqw/F6g64hzL/EE34hKL1apmj+zxq6FkoDY74d1uyXrfP8
PLckUqNuskSh9h7etAfUtH3w00j08NbHuAnYjU38C5YuCqbqwNjRTA+M+6FUXXq/
FqLx+zwy2ijipxh7CFc7Yk2PIx1S0tBsYfA7AaJg4o5UeYviOldYtO9ijVOr8VzA
41yeLYjOY/RsmsdqGmihqCKXvLxHXiCbCkwWU9koaggDpjYbJJqLaMpmMasIHqOZ
+cYfNmT4YENMpqB8MGmZOj71XibM0Zwh8pOQt86cMf5agfFyup8VA+e25JzciKm0
MXAEE/6bdjMM8HgnURMrsq1AoJWzO1dOIEt8yx3rwisvPzrOVHPXaifEd/Lo3dzr
EvsB+2DaZsMRfRPGr+koi8wAzGA+vV8PIuHG6t5mjSZhqHEb50jf6m5LH+v52jAK
7t0OJ8BCiuIkHU9D4k4M94PpHqB2PInfWeJBdJcN+RV7Kk8JAFL14RUn1XWw0f7s
2wtWCZw9G4EpJ9/voUxKbZLhVYm4LIPvuI89gIhlxlJOb3klzHUlQjrHL12PdL7Q
RWcrUqzbcm9QHOOiSwTRYJ6y/O0krzAGROap0PUiu6OLblM3z3QdrUy2rSTXoP2U
q9xeLZmUmKR5bO/P/pBgL/TmCPmH5J4rUc3HWgy0dlF12ovSmh05fU2c0FEQ9x5N
9IN323orO0Tv3N7vrmUEbe7zCcLwm2pV+lkg0+qA1Zn2IQL9ztz7Rgeuo9IU+r/i
V5ZNHO4lpeEN75G4W9FrVdEScW/ghFd1kFcxn0iFScv5NfqEympwSQyRluE7wAa2
lhY2Z3a9i9L97OzKS+qky9hiHpfjRrCjGwb0U1iw1raZ+uPbrUzp4zJVc3h941tB
W0JfXNsAOAfiTknHN+iUmLRbPRp6CM4IBKhI0Z8oHyTfReOk6zUBpKYnVmMqpVzE
Z1o2bl8+cF9ja8GX3HY4NA4Cx/tu/V6MRej3GjWN4OBrle+NVQDMNkAfgLgrIE4Q
zMT1e/sx5yOjrJBIKuD+oWQYsQiy3VjaAM4R7YtKWnP1unDa6nX5yTbLnJrR5Dd6
JG0c1+mCtxbyIOAWy2b/4R+8xHZjFkuCgeGeqS30opE4dfaSCUwCzN4+7MvxNJ+/
iKiVGE3k3Tlhpmr7+hlzIhnAKYstLgFMGpM7xyKjvueovfeFePYvFvqMrBJ6OB9T
eVv0CftnWFzpy8JBNtQSlkiamGik/lguUAkvflo/kXQN///WsI0Fn8HCvGjA4UaV
Qj6dd30axeuKDrwSWVT1HuBK8MvGDIUWhkqcLRR0KMUnBqKzoWpnzfNCYp85GjEM
dh3k4VfJ1kLDK6wR2lPA6fzc89wAvOf3KcZtzSSvOEcc/5ld9UQneSJQ1Og9+/r1
sITOlKZOLX5e1lcWkTGyj/tEQaFLrNwX6HTSjIgNDooqpz3h5rQUzQQbo8642UEz
K5kSMW3Avj4DIx9Mov8er4SOoWEaZgFy37m5V+xoYBbKL0kQw1kKaaf1NH6rzwme
AJHGbKtET4RdFTQysA6EKqBq9rfPp8DK9Pe5nD25pZOLSW52sEOQY2wIITV2k3Lq
yQhNPquWjdKWYaTh4OILuOCjPtgC8m1Rby9xlzY+QsmShW+hGhs30zRh1y6+70lU
yYDdXI0j6D89C/3VQDzFpeX1F4y4abkqry/pKDvXNSB7FWS1mQ8W+7ju+0WicQl5
ndPdGVCiUDg/xMvzUsEGzbN8kMWbKK46CNMUOzQ71BurgxkXQwiOZfetrmyJqe0t
hGogrKrivYHz91La/lRyYPTLcJ45Cii4qPVtpbt2R0iKQxfs/QBj1s2SLYzAzEmY
0yIg2MfyHzvzIs2mOySzg1mBWd1uyHI0uCtkEMHwUKi5xvERx9cjXdpJPyYORxnb
3UezN08HBFMuLckKmRKBnJOtjIX+eWRtFw6TB9SfA/ojUgCBe2/FMUFJhhrDJChH
dSt071M57WOWw0TDqv6cutou6KRoaeYGS5rr00pQWDyhwSOmlaWvqGeTKny98yjj
rI5j3alwT946ILJGOx8SUooNa3yAi6WNH+QyuawAbZj/C49BdY4d81KwWt1yzqLy
bi4Ae12/LVfqKnKfJZVygiPit2dRqAmop5PdTANSFLKQOcrZDjGU8u9CXz4/GjwL
6mWzJmTnas9GmzWJgmSwpzH9IFooNpmtpgNS55AUpBNSmWYajHOR2/NxC781bV9t
vK+1zuOV5B0ipEadhvB+FMV60fysXw5D/TXSoaLoufujGpjUTDNxszRoQA2hN6Mt
pnRTjJitTxHY/pw507P3lrTwuYnfUAjNfsh1uwQ7xsVL3cmtkoxTfS5u3db/6VC/
y+o8n4mCQUmpzs72G/NUYtiSWJIhEZyLxbfuv7IivvjEpddJWh1pHdEm68YPWzcW
Sp+LsoYMF+EeClwThC+4QCrQtsaqSU+uRqcPZ7flhBoyroXAUCHmubjT1MzOqkUu
A9qyj0xYabZbeg8vGwoHTJyekDMQR1AuJZTe6/LJXz4KkXVsjUkXIF+m8bDxSx2P
Vh/R5OwoLklBc2+K8uZOlVBD+ctwrrOSg8KKkxikg1/BRoqtFBzeB5Z6dRFfiPo5
Ab2tdZ4d1aSEhVgzhZVs5YrzWLpbJLvijkgMK9fG8JWxBnWsCqRBpxKt7ypAgbaJ
Xw9SQKxD6EW6B3C5Y2iH2ZWlZt/kOfbqY6W8e393v1E09706Rs2+AU0IrNrdv7jL
zB8hp1MVaxA4+mx9aIQ1XLKNs+HKx10fSoR20o9UUWNEjek0fQBIJoKC6p68t55Y
viPHwBy56zEvTCoT9O5NcdQcMsVhwWlVmh9MBgiqYXINBzr+rTgzD7fR3lDwNj9r
672gPC5OqnBQH8dLkUZHZ/8oOAdTUs4s9hx5XsPRQvb+uzYdVxui3xrucxcuERHW
VndI6h8i8amj6wTGRfuISpYDYfrNbUCGl22J4121N9OjrOsJWiFPmDwUOSW9HS02
HbOyaTrXUjIJ9clBmd6HZDiiRgJqX0huvhYBiXrcjIZ4zhrdCpo60tpIUvgbjFvK
LERZIYwSgU4R+nkS1x/SjrSr2jd7psa2gpYc7TH6UbFbOkaSYk8MGa33BoeZuTXC
snyihvGFirfvUFNyG+ups0qKnPXZf55HUGO71AdP0+q5cRo/9Y2o0sBr6cnSGJ8Y
/ELuneMR4KygdYbPV01cKazpuieXoaHfBAKwc3KfBuOPtnvI0r/4JS2wlD8F2bwm
p3S2b0oUNTQbPl3+aFfJ+fA5RvNi3HhEMPIRyPqSQRSlhzlKy+4VvZvA++X6Icv6
tYqmvPBmcWLIlVLZveC0V4zMcmvghYMbVjGmHDVnKjhiPwwoTCURqjcfT5IK5yHr
bK557ovaJvcZOwrnRo9xpMsQXDklk+8bEdd0Uzuy7HAV3XoejZFezBVGbF1zzg3q
6jRdz3M8kgAdnqHbWwF7ZdC8GYyIUTbYxF64xy0dkaLSWJOacQqSQE7HoWpRQ0w1
p3sL9XA14ytFmyShlXBOgD8zrG+ZKrnVMQ2nmuC7uLzFCbV2DfER63qXRR7oWBPr
qdepz8RgxvBBCrkeW7AoVlDR6wVAIcAtdAMUYOlrNMdDTas9JS2vnVJPLLZQS2AE
2IRbFdmCehMypU71pZ0mzPDRB3EfAuFROYZWXYp+Rpkd3kSa5Vvx/nr1/P4L65qf
pzpILaWfXdJjt5a4LDK62FBxDbzqFFCjeZiQgAGLbyrCpYqL9qwFIGUzl6PSaA3T
eu/WnK0ZNqsTeoMtMWd5STVlWhCzjv2w/NBuDx9nJOLNpLK+wFFAnM5DvTFL5zyw
jhcJ4krLgEUrMDkS3k4h9IUfhgAihTYioGnn73AjuORojr+kZWenjpL/3NSGaDOL
+GpB5D5A5E/OuEYOVOPYLFVSemZsXlnQ4Za8YHFi7b/E1zpNpW8ihuMlXD3smLED
4CRyuJYorXi1gpT0yyCBv3KCpcCE1HgjmoRageTJMX+dgp4D+PZBf4hhXrdPoOkW
7sj1EGNnJv6rOiYHJcygDpc7Ej6/uUUDZi8NQO//MXKklV88buN25IBjacysvz/2
DgQeHhlFXsZSHaslmyuKXM6ihYB/r/me85Zols4iDTaVaTUJqXUITaHufPBSjGk+
IEGZd4DGgXTCzOiwqgVWy5XsTwFcmqX8NbC0Dgaumi08HSYH85hUNdbz/GN6viOO
Dl6072cwoR5zkUswzHkrl9gqLrgqmtnsvIPNtlNB4ao1pYKT7jw6x4dwR7ZLNErN
t5aknBZacDrI7+/8T1qYS5opPY1C46Y990ruW5j6p6Lj0GIMgJsvaeFgVVjKuBNh
h1cxhYFZTNmz0hAx/IevwSQIsbFg5AqQvsoT+ceQw8ZlmnPBCWik13El84Xnw86v
FYwmZoCo30R7DApK4p3IydxTv0ICuKJ69jof5mJeTolsFeRibPWl+rOs3jFoKIvO
oK2QQTf4wCMyNnr/vjYvKgMpHPfya9kjTDkjR2+arCVrSpu3c1trP7P3m/WMP281
L0xjtZEoMsVWFGcn5j1DM5zSyVba6gZOWAUaEDuJqgv5Xs19UQY+q7dJcYVQWYQU
HWhgqnxwkx/85INmX+/dTysH53e+zmy2ux7sPccNVVIhT9BQfLGKYfHiyJEHAxA3
qkO+U9ACaJ8kY7WuvAH5WMFtXVoEsl1BTQt2nNHpXMzmx/cpbluhNmH6KjNukKPC
yFAq0OSxbktZlfncWaekYfc3MXvTSPFPwixLhFTzt9QRz1S0wUKJ8cI0MrBAdQiu
09NqwwzPrxsyq/SeoLhE+/2r3ld6VShZf6ouSwhQ80QjkZXxzFQGBBGVyjF0b9ub
4SSdNSgkZ2K/s1kKQ0zMXcKdZ2Nc1OOw6GI6aC6NY4xrjOCIn9FEKv3W4lZ7bOPg
bfiBlBHyPmo6nfmLIZQbWIU7HuLruWpEzcrZcUufA9O+uSf0ZwnrTz4xT0SXG9eQ
zcRMpeT2fIwFKQO3nIZKKdhg8YU161C3247uOdMUhmPGTf8ljyuqLTupSHiSx9cT
2Zr1Vsa6VTv1wfNxlEyCk0L/2xlIZL4NU7hjCMQQdUmLRbEAeqp6AGShIRrjPF3/
F7fHGCT9arCuezQCmWXQG7mciy858Q3dPhpV6FmE1G5++obht4lnRXE7ebo0gbmG
okRUGTccSuKEsNhqDUh7YB9zezRfhynY47dJjVg+41E6N+tiabyZ7oZYVtKTssiJ
os4xBOrvB+0O16ljlBfgJW7pb8Bh7NjoLxKwXCBz6iSmCaB5miagd+1UoHJr74Wo
YEq1F065ftq6TK7FUt5AKqJtiGRXFIeBQrqK5O9jgOQMA7uSAVtuzUMmxvNYbX2h
X29nkTW7HVuLxziBPidtuPI23kn8c7uSjV6vveXMS+/XwqMeg3AZeoViagPrH0DO
1yH2ifSErwbirloW/w9pU2b9FYE0yqfAOML/hG/itWvq8ReMI5nRANwFBZMF7cDl
HN51hgyi+8d4F2sftynSPR7jXTr7Ic6geu1HwMEhdFI97jzTUFhExP22Sjmu1cvP
+NzJoooz8nXqWEbI5A23+Ma3ROmIMd1dtZAlF+uEmhsaWDsJhjc1bL3lP3QHIzZQ
mbBsGhcgKYOwzRiBW5RczFkq32EBAKngwuzCnnsGe9JClQY37OZPQEG02pUXdCra
/gnMlS72bShOcswRLDPSCbpSSwGNtyGnfJl6sAuCyMKz74hMy2hsFI6Z7G6rFX6Z
3dX8AjSCmkTuo8GIF4JSbRFdyt9+wlNmFCZ+pq+7wN+7+HFDonQ4ljn5Ra5OBajy
pNahxuvl9YxcDbqjOHc6pj+fmJvFmldPhEicFHhtgCS5RoQj4g5XDFJ21vFS302X
GxTYwFwN6HK7J5FQFg4h96jS6vQ7MgnkIjFQbY6Nu+KIxf11lQ3JHjSUaDPLDIk3
r5IR1cTqoHHEKpJ1iUboGi9u8KLhmK17b51ofMy82f5w1m4Smvw3cM7MUKObw1G1
wucTSQcBUXkS7gpTaRslQNKQwLJaZ6gg6UXNYVVh2kdqtucy7zIG+BBARft2c15b
XttMldr4B3Ku+RWQ11Wxn/Rt8flUQ0rQMBNsj8JUEvZkifXaPyFNqh0Got0MH4ds
Ir+zLqES3OmxSwF8Ke08Cybl/m/Sf7Puf02gXjCJ8iU7zpPl92yn+9qRs1qE5Mnw
zCDANS70iKnFI3zS5vJVRBxXcERcmGeTvHh+w089W+4wlft2uIO94gcTuKuzMUes
oAh99aDm16w55tVDj8Shn8zvM6lh2Kq8EI/ZCF01ewQ5QIStB2WzMKNkVOueLb86
7E1LYJ4/e7XXJtCoufBf6RVja3bk5s/rcQn98L65SwICY9trZNDX6WmyCZg0qnHI
AMOJY0EjzOKnStWVbGwJGrHBPWdBZlsUHmD/8zx/stQPTXzr/HrA/LU049yq1YMJ
Zy27N2s8242PMx6ZtEOjpKsSkl41XHE3o1bCuh5ctBOFVlgPTms7ralntPBjbHFw
7PMlJqfQRKOoXoFRPdtC4jyO0Epy6Qd1af6A06YlvU4WdQOlAVcEHWaUYX+gpE13
nlkHzWajjWcaID87uLNxS0KfBfZYNc67TMUdLu0mqFqdsCKdzosxwc8RbxuahWfV
dShi4WM0RL6Rqct727aA90uLI5OcY1eyJA2R2kA585F+axDSMMi9kJH3MwtukD4J
NSIZ3mhnAWMEmJ2JVc2R+ruPr0llh/lQhCNLFQGabrgvoV+ah7COClwKESlCgrRu
Ce0MiVSzWl1vbZCtz6yRK0Ke2B2DCBrc5URygy1Nf00hakt1tbP72M09ra/DXsE5
0ph7mMqwvCuJl915NuLghCHn+W0k3oNaYgooyKpq/L7pSpOoTDHGNfcnM0ZBRmr1
eq+LDOkJDrUauzcvUcCu6TP7nv4K939d/uFPTBu+a9oGqnU/XgWx4WvLyLCXiZtM
oRLZzuPgKnuiJajS3IVmXf/csG7AyuEZpwTdYTsK0s0B1A7WZzDeXSOcokHYhHr9
WtBvCChPjmd/V4VSeDgterI/Nqzkq+0Ciszf/ygUql1mcc+6ro6VmA87SwkHt+bB
hpKyZAbAg9ML18+kEUaKzX6u6GRnIAB35q5NPwqZzoK80MUg+eq7sl5YcdcMBYnr
ieBmnIT1kUXB23CJKlx+0lA9YcklU1JcX6jYEhQby8SEqq3oFMvmgexb5aNf9+q/
qmKpNUG0477ArW9AvcraKE3rkXZp2kl5lhcRJ2Elmv8=
`protect END_PROTECTED
