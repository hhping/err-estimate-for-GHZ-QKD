`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZoqT1//s2pKYdGwSTAzi7TMY6ynMh5bqz8QDk02P3criZ+dFZoXjQL2X5wHi9fo0
qPQ0dPUI++SWF8s5SMwtJ/fwVxyn1ZriuX4kxK6Pu6CMAZ3n/PZf2ibVMkiT0PEK
IPF0xCctYnTu517cDY2zeNGaGmDQ+doAGQk+uVQU5S6aT3qm9hxjXPKHXEyV7Wam
/mXZSQ64aHcSjrmmaItlngX8R5ig94zgyEatsgF8zCg+F26ty/5bySPSE0aiXUko
gdtRlzspM72GsehU/rKn7HJaSmjcQtmrEXgULxg75g8JczwhvZfo6mSSTmYGId/a
75l8HbDeXTt11hOZtYN/tx1q8v205Eg4mgtjD0AUxJOeKM2967C54/OcLL8OArlT
e6QlEotiKEUu9TlghBULwNqKLlpGiSy4h+7XV59+AKkVYTruwpALdnMRG2qX2eK1
1wGKQoxi3C1zXn5tyGMx+Xrx3CTAtzdlLJYiCFMV6aIiJzwaVwGaSR74v/KTDj1u
Xik2b1mMlNNE9iBwuJ/iKVqGL5g+oK/UA562+GnjnfR41UpRQy9gEe0HpGvPSBMy
kIsjin7CcEHZtR4QGNSj2F5PJIVINvY8CZ29qbrWjU7uy0gGHu1+y8K8Nn8tR6HB
Rj2cXbFiu0bCqNoXnjLg2NsQt/TkpxWTa2PB0GNDBUptf5fp6BhDzqBvM2SDhQnp
asVzJvaNvOGlvjQHN73ot52tZtru2lIpbuI/fk/ztETVd072EpOroy6OxlVn4mtu
HdGCqw3JT+J1ZJo4h+MFFMYmkPVmL+GnoR7x1SxkH0kLbrsgruqUFWrVaj5GXpNe
JSAy0sOoIvFl3HBdqKiBbs92QLVguWylPMDnjKFBEEkuuTp8NDdeD+fOrQJj2T2i
6D01C3FeL741zJ4sADmatgQBhwi1kCDU3zHKKsIcdAsRAste/4lV0SY60oj5UYCp
24SHAFVW9J5Ragoe/0hw/Q2jwi1yjMKthu6cuLRuyHSwWUFzNV5Wz4IAsvtKd4LV
ZbLECP8ZbD9g/9+FJf2PayHZR2tx6kFgPHOqhmciwpuNivl6t5T4hwoSHvJY/dlp
AGwhET8BUz/rZs+JYixPPRWNbjBWiy/Hz2ZeUBI2O0a4imkm0S6LZ+1miAb0nUl7
QB6UKlwiz27fHWwMO/9YQpsjo6VciHU+00Ke2hCIc5MNZkKJ6EyMpWoyPdbwfHRE
6qkOxUgMqz9ArS4xb/ZF4tZ2/4l7r/Z8Gp/3FqfVB65ABSGvueQypajdNrbzeyVv
foxusVOYVyLIgVmuHfNcCRYsiwfEm3rMxsH0ezMSCv4OGLPZu7b9Va7rQCcq1RmQ
Th0qtOMItT9751bxu6uXjgeRhTIT7r1O54jloDa3M6jAdu2++nwggA8xU0mAvqwA
sDHpEouDuFvfw0+bNE8FVdlUe3TKbXJIlzU0DJgquZ+KoIik5Dr6FDmK8KYz04mf
4w46r+4UPU/aOseuhk6bzAQkbIMV0juleaLqNuCawW+FoN8oTx9AJdKwEufgStLq
WuFub51SIHybEnnn5yeLLEj0NxGe/MnCCF/gV9VSTyx20xvJqob4Bo7DyNG8eP8G
4IV9EsgAxjBg24JMPDvCEdAeBKd0sbA4uz3uyVZVWGyciKJLybsKuKP2xf43iLQE
CB1yMDVT6F4EDoRi0sOyrJH/KE7fHi0PrBDvL0IAWErCqm6PKhi+64HhcvD+BI8q
fNydMYrpXEqHde4DUSRbR9wmULRi5qUoSRfPTTISLInzvo4R+ZN5hpxDSzd+L8/L
MhBXpu4Vkcya042bcYB9zWTPFODd/S4X50snA+1I2+DyXJ2kq5pWxLshzfoVBFpq
rEY3HAV0G21XVqOeH3hHoKyR5nhWtcWXp0RQ4ZlSznFuGlIYolOLYK1gVEo/IfDt
Re8rF+f9jb2DdgbeKLndwUVm16MwOrZASInbOdRWDDtAAFCEzMHr0uh6YNLVdKV1
DCI4WDm7tm05rBFpFyno5aEQRV/MjthNlBO4nBeMJ6xCvl8J7cCAzqaisvoh1+xc
vmDLYs82uM0CwIoTiRHZq2N6XHHAga6/xxNWdoIYeCGuM7CU3BjXX0Mp3bs7Y8PY
AlkVzRmGSdgQ2N5ae8vHYk/hPmwABZlWkOCVLtD4ePhUvx0Nd+LwF7vfnM27dkf2
uCZ+Tlau6B8LWgfC1nD6Pe0bxHNDXx341OFtyxc0th4lMQDCYNSTTogqyDpEpKjR
RHcsn0eQOe8UiD/gWZcx2lEpWSFNfDPjBFo1fI5cch+lXup9qf/3mhjZu99w6Kdn
xMxxaTnYutVv1Z3eGnuGwuI/cb2bcp1ZCtN3YhwzN0w3SI7rA3845UxIT06L8mXb
uXjM03+ihOlJ944TbqWGyl/QunbEEg7BN2AJviuwBXR3I4A6kjlwzrhN4Vw+876z
taOmvlhMwz65kJUIY4nUUtPIXa6cfwwc5kASSPc2BFbT8lfUbtgAhqOAzCVHXeAB
iwOLP5L/EpOrB2hEZdFMSVloKI9d/YmyqTfbOZux6Y5O5p0c/4YUm1eKsUJdoIGg
cyIwH7HhCzCTITQOjEDZ1lE4TeHByXmAMCjl8ffbKyRq0Kgk++W3xz6+Z0zxiguY
iGtOVbw/5aAWmN9b2aKOoRf29lWX7KMcMxmcmHHtOEMwzmYYqlbwed9ESAMkrb5a
M7inyuDaTI0xdCAvIOBvmPWBdiKkf0fcu4Pyi83oruWwBr1CRVPxN8yoO8QxscYG
sYiazmB130K6Jf7dsUqhKhfVY4t8MAK+53FbBsYmU3DPvSSS/rCoGslvm2vpjUHb
ztSsHKUwa40XaGlcRWLR6BHMFthlIeEvZ2zlWhRMrTqrO8V17aqU/lgOkPcVO8ce
8ASbYktmkHHYs0TEeRWRLngoV/rKoolk25iOnO/QOuIxqHQW/TBPOR76N60GyzNS
3CGBSAwLp+N2DSBdUR0LM/+H1EMaOYbSAAyYv0PBuSsIzsQeTBX9tEoI5+ra39tz
/aQZfyUIoe4gF+Mq8oFVUQ/kvKpjDHFOe9T4ATDWvwH7YeyH6cP75rw85J/I/c8B
fQQLMYnr8qSIhORLcME1BRcCi3XAHfzVCDtfeqpuxxOEjrgiWbMWiQZ9rrJ77KGT
iEWmYLy/aQZoCgP3aUhyVpcDA6hC/aCb4ESNc25a90s=
`protect END_PROTECTED
