`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wO4lgVgftB5+M07tbKMnQTfQK6FTVnztxIXMQOVxEd/L1lU+yozGvO/d/v0v8glX
jhfpbp3PjLLjWSPJ58ZEZsWQNwLqvR9aT9m3i6mU6sQ14Jj/GemPtAdPhoG9ID/H
wqRzMrhTojUBd9evHCHSdofqZzEHHuJmLlmJWBykeYV+XMvViqhYiQbrDD78Gbnx
bc3mkFBqCLf/K7vnpAimmNsD5eJK19UHlRgiEKTqL0Pg5J52eTM2O5DJGuDiQqr7
3z+NoXbuqYQU5FSTNr4SCD9VKYWpGSLHAxNnp8KOtjhn7ujg+3hU9oZkcVgsVUHE
57vYnKyKEoQUoFKNt4QDsWtLsPfa0Skiin24fIcyek7SJFj8sjID9ho2FBJX1Z23
n+IvtYccZDZmFzUy7RI/peaa/wRVuQukVS2UgmYjXedBaltUOQ1KycyOJP7XHRFY
zPrTnvacxNVe89D6UozUPTuI0dFcPQS0icOwDWi6ADRmtYJSUK6N89Juo7t66vsF
bfPQeJDR3OV1VVlgk3b4WbX/8S/4N/Cao1Gel3CvI+Z2E5D3jXKUT1sJQ1zmjZWN
Srq9nfFmxtPz2VinuZL9aCmApAcW4I9uIHogRaJn7LadU1DqDOrSIB65pZsuX1YU
UngwT2Tm7wd+xU2oivRF4j9EqSZWre262Q1Hbt6+iz7tQ9NjYRmiWzgp/93a7NzP
BeOhhVtjehnthrM1mBzf7vcmoS5bDet5z/Zhbw1Wr6ZoV9xEMqAbLWifxT/7KgDm
O0740+bd1iGIJZnJFsPE59dUkz5HNdTaZ81hWhzU/3shQvS0aicujSH5tqAZHmTC
gWmHypFewZTnwdB268g9lOBq7iqQ0VwJDmxnJpBLeZ/lJ5H6i7YqVKUpf9JL+5Ah
Q68QgB0KbKQfgS6JNIuLG9BHKcvTL1HQEJNnlFf/eq+4TfhXbis2k93NP0f61vin
zeBsz/6Tb4AQ9qOVidTH0+hnIqXXAJtjSltMhg6ikRxHD5bGXb7eNzcLDBbHchmM
0WUYoSBJovkhpqGdQX++oEllz2VDuAXJzbSpbHBNQEuAmWmiGmiBQW3tVx/ZQoGY
eFTftVNsmWjRZ+09zWDL0O6RkpBsZVZTxye3ZHTi3T9zcOBEeegzhjQrzY9IXqzS
v+i/uzEBYD3pQC95CnVA1oc8HwvuIqZk8pwLD/zP5llCJvC7g2eMMCaYftDOHRfi
YWBIXOVXkkOz7wglRuGwqRePC7WJm/Rn40ngGon5RiRFOxgw/nbiHeU+HH1xQaxX
VzMqkQ56wV/x6YrJ02HUUxcAm/Zwyxxy+Cl3VaDWkMFBgH5/XvNYl5f6VZJha44N
6riqU/XlVWtVEVSxKAF2Dga2SEpxXXvzncbdv28OtO2iHSLz8HqfkTHk0DCbHNjD
n9GYI0Z8ORtLyL3czc8J51f9b4HPSBSFeTax5e6b/68Y/2vVuXGOhMd/967bQoUs
rGC53Av5Ozpv1ekPInhzeQxRfg6wdl75KDavMxyVoa7H8ZvQy6yHIj8PgdAUdkNk
WMd5ylEPMYMu1yysHfPQ84qgj6fMDmDKP/m+xQA43j3Lxw/RMc7ykyiG7vk6NCoK
5HWPpb4cTi/HidpbBpUcncxbNF+WPFz7XmSyemIY8RnJ8gT5OmrHbwGAk5agXEcF
w9KdP14qlKk/EgEP4cqGY3iorV7DSju2z+PFBq3aWiPR5bBxf3lHG9+P+5QpqriK
JNyGJebSmU7ekFVEJVowfi5Pv+DB9XlnTf0w0wip5L53JrYZjfBvFBb90TvcqIJw
eg7XuTxa6swqIFD5StZmuW7S/tpAVVjinQXOZtq9HiXcdN5H2NEWHy2A21JRvnWa
VPRKpAAxX6tf0hSo/2VS/wGhqI1t9t4SdvqNQP51hlaiPjODtn5GQTE8DtzKb42Y
lRTB/Q5/jtxMHOnA8N6HrpMwddFjwT965RIDnIgV5AsAFWGBkMjR4MEhrRbcuCv5
cy13XywA30YiG86UxE5p0sWFqosxN0dNaX9FJ5qYBSYvldw+Ar0TGZtdHuOyJ6/O
S68RVssrWBBW7AS5EHNxOoU2Tt/CBEbAaUJL4V/ipVonoGQHMCKDtZ3Wy2G4Ifhw
kW+t6PKjFVx/G1Y4oWIi4cMdj54qBHH4YdJAwtBQXBPIwgIQyuPhVVYDL3WpA2YP
vNqCuOebjqRWqOpBGnMdLX1x3EV4f2o3/hMjZ47adEWVCSkvKUMjRtegHwLMSOws
4hbJNZTnKjDSwHLlB9U32sAvYS4MZ298ehylkQCCPcJbnddnCzewn/lIayik+70r
qvDNmTk/tP4txx1EpkJbS4Y3n73jQsMcbC6j08UkSAhg0fMtAu2k8mN7yXq/8PUi
J2o41FvPQsdMzq/JYtL4i+G1pfpIOpoQk23b5XDDYAgLEm2y7fRzUXeA//rZaytW
sV3TT/PI0FHFimJxy5F5lDBNQpdS1aFj4CzXBnwsWJziPsjgDYIG6NCUAIL55KhA
zeTZnvSzLDPplh5CvUbSpadCXHYF7paiZ4kxr8vmNiFYH53YsPj3Aadcx/b26skH
ZsdYyGg64pDbKtWWqxWms9SMYenEob1DYsttpABbcmL7aGrWHveU05oHH4Z042K2
kOHLm9cghO8ETB6Xe7BH4xrXiiaSkaohFU6bUMO0vn++P0cApujjo5X9/fuuIhpG
VPy2bTUcdmuyCki1l1gFhpT8YeW30KC9dEUf5mSFKjU/hT5U/jG1krVug8/lB5BR
lEre/lyonCrPLjoCulxHnPCtRFqaA+bSLi+xAMBphYQ1omTwU2knY7xRlk8VxB6N
pbUT1LXSYK5gRGQd6HgGY8ciRmeFIBIwV48pySRp4eyFBaQXcRviOAvBey3UBQ7H
oZAwfbwY2t6aLWr6H9MfYyLGR9SZsrJMPN8SiXEiaJu/KDbafjvcpG/FI9MXZwJ1
IP35DNPQrRlCm2zW3JsoZ0iVqEA5lC7FFQWz2SUhH99fXnG7aZf9AFxnyOnoTf7z
prNByMJg6EA5P+Ym0e8fDmZB+xTuM7e8wTPOTmA0x8NVar7Oel5PtHSBYP0D3Spq
Kv71q+N4LBMh5//Bqt2QNpjGdVpk6zodZ4IsFn0ZR3DPR2gg2MK2YCFUf+g1duG1
qxgHDIStEPXLD76vYnfBO/RBMMYZZsFgo2cvH3j3a+ZAVYkxsiskLSK14zqe5Jhu
7r98Y+1THadiCCFf0eC2/JojJt+Mmq5Nee7B4Hi2lyVqSlmBU43Vf8F60490mYax
6tU382MOLvENIxfSBGAjqF9eydc6ABJmi52OwLziUTN9uQKcrHYrUxZxyS/KaZGw
AWOLa9Rs5z21F5Ydb3pJ/1rHMlwnLit9R3lSz+4rqwbcB6Ie5QniACCLB2RRDiGo
fjiaHm6oDnMNA2izDaUV5vRo4NSdmebK6Im5Jv6ziGJxjJ+UXGhOlq5hyY4T3el/
JJnhjYYYIUTnJWYdagIMY/2G2iV3CVwkD320ltjq2VjKrDbVYxzJJrHW3wivocFG
QMXvODi5pnbrF/Erety+tegog/c1nv0uN3VQftLMoqdMOKYbxutPIEf021Tosuso
/WYvnB4Al1UWJDPI2o+TnVHiIf3hVrgXa3UMTszDfDeIN+Uj+VDmc+PoyTG02ilU
1Kj+fnMHZ+YmASM9FGBnBPoVqGYUtaremjXrgahnn/7BCHdq/ytLmLwwk4zK9vn4
Rj07YvAZwLsOQ6MXnpp5f17xT4VSWfZx6oFnfNV8k3u0hxunwY9CBVc8PW+dyNCJ
aXRzrOSy/+xnf5qyHEwYKFH+Raw6KEkPirk1eFiPnkyXdN5B3suJsFY/r+wycHNG
eeKBdNSUO9e16WSIIE8tcarXvITHCegPV9J3lZ0ZdNUREbizVVnvLRvL9oZw8YLA
hPL/Gvkbxy4o184svIz0S7MSNWStAVJ03ekC1JbZ2T3mZQxj+rkfT/gddOTamH1l
DTZftknaPMLwfzY9rTGeyiQ0M1p4cHFjuICmrlYNhnij8YFuniegdqPnrNaCE5LC
t7NhDxfB27ObgeudvuFWTZurbsdpuwAZ8AwTMZETHNgrH37e7M9H4dzdkov/1WD6
VrWSxfQ885pz8hh8ruHjp9uT1jv8ki+wCR9o0/60S5xGWwA+VyccP55FpL5W/TVT
v/aQMAc5ibnAnqjF6n2M8y0P54h3iIiy72/wxON7mEr1qGS+DDPFtc0j8x6ZJj36
SkgOuHLqFSp6SKcZJxXY7SuQpxfT8u6LRoeY3eV3Zm1mLlvZ8SF7nrMKAUKp+yW3
U2a9qDNL/4cWZX+yiF6jlaaLj+5yEvdkYyUgXOHXPjKi8TT+a1b6gZwAGafJ8sIZ
ebcL6OHAlH/5eaRF/Ela36FG1kPVBPMVIEm3S3X+0Vc/LiRxNErpB8GWyzlg8IBZ
+yfB7YrfSBNyRgGVgS3X4zEhrEoJqFyJqR3KhtEg9Jd9QmVTjwh5+jB7Uc69PBLf
nsr6JBJzgWTGGuKSPne28XwNof2NW08nluVIfYO0lUCDcT7ONP+7LS7nFlP35Ced
mUg2PRtf6jjkBs7oeKxvpipQ4vfDce3DC7ELRk+g9Fcy4ZfNp03cgMDvsYywsBbg
wOTCSWIJF8ExiDyZ43sf/4rF3K26bFjqUdmO92nLg5Qz14zCoDEIr2jCab/daSdh
wAzDdYN1x9mbrqN6dQq9dA==
`protect END_PROTECTED
