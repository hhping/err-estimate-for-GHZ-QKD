`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LJEtZFIMgQybH5ppn4b8bUr6zTaBjelZ9IiBIBGY3AmadO6G53oLnAqRr0CLXTHz
bTcL+yG+k3motDoerLYZtRL/iF4qKvJLEteSRDyb+IBman/hLIbdm2myWmzPoazO
iPUx0UszpjAZ9P7suRkFRSB3KLtzgfCe7eT2NcblfkZCb662LSE7vNYtCuJozOiB
z69Y9EI9NY/MdOIvpepVr77tplhP1xqbgIuEPtwDzYvNkOkzUu66S2ZhbWBS+BXS
F9hkBsSno/G7Z7HKIHfD1aKqS1qyuwxa61DLm/K5YXNZ+pnfRi1BQ/0qbMOX1UdJ
K+Wa//dJJNfCz5AH6XVeKpMJXaYk/lt6U/Bz0IyeiNEz11UBu1ZmEXG8BYF8gas4
za8Cej7u4ppM1HXIsY/BeyDR0x+ufVqVQKPnq19DmQr6ZYWpsA3vxEwpfZpOOm+2
g0y9cZLSSqmNJyM7DH/DxfmfwEbDRJpYfaR6lv/TO/IwqODX/80WSvcNcP5pVChS
HQ6VPbu5uuJONp7w2Twv9iWihVqvUGAG1/aXGwpJFhH92AfNFMJP1KaX83kRkENq
7wjhd70uZx3qZicdkV5E+vspQ6MGA9aut0Mw9gzPn37pTFDE7CHzVwYdIb+X6wXW
CxhCeLZ7CzAYTwyCxE/qnI3vCJW8rGe2SpeTyTvrLwiQ0+ZPPXQxqOoyitzYTCG2
vNIP4VegfQTHYk3If/ALBcAbXoFF3b+bnSe1/QKxBehR2F4jLd1ryWqb7vqacLZd
`protect END_PROTECTED
