`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1N4vjWxQ6ryxbWqG+7rR6C1GZ2vWtTa4vg/D5sFHiHI3WS6io3MUkcUxnfoFiSN
DxvtCPNAbT5j+JhzVKlfC8P/O3fvp9fPh6Eiyg1CFDQLAkV25LhNVHSTGQrjHqjj
FLjZioFALZk+UDu7oPCGsXRX7U90sA/CHCUCozBdihq2Is4mqe6DO+hSz51rbBC3
Wfl4ubOHhuj/m2KqcNolR+m8kfxVKCBknY6w1BWgIWweV5EkfAGiW87rnlGn9MIQ
btWd5+BB/U6iniCxHlec8JzJD/ZuhmqU3yfHug1wzMesxJ6S0ZpQ6Nt72oODJDbN
ypWT+Fh3YNR0+2e6vtwUd0V6pbUxoidFywKn9velX+njebH7HQYkSVZLlPs0i2S1
1oUgm4lfw9P+aHd/iXAK3A==
`protect END_PROTECTED
