library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_rx_pcs_pma_interface is
    generic(
        enable_debug_info: string  := "true";
        block_sel       : string  := "eight_g_pcs";
        channel_operation_mode: string  := "tx_rx_pair_enabled";
        clkslip_sel     : string  := "pld";
        lpbk_en         : string  := "disable";
        master_clk_sel  : string  := "master_rx_pma_clk";
        pldif_datawidth_mode: string  := "pldif_data_10bit";
        pma_dw_rx       : string  := "pma_8b_rx";
        pma_if_dft_en   : string  := "dft_dis";
        pma_if_dft_val  : string  := "dft_0";
        prbs9_dwidth    : string  := "prbs9_64b";
        prbs_clken      : string  := "prbs_clk_dis";
        prbs_ver        : string  := "prbs_off";
        prot_mode_rx    : string  := "disabled_prot_mode_rx";
        reconfig_settings: string  := "{}";
        rx_dyn_polarity_inversion: string  := "rx_dyn_polinv_dis";
        rx_lpbk_en      : string  := "lpbk_dis";
        rx_prbs_force_signal_ok: string  := "unforce_sig_ok";
        rx_prbs_mask    : string  := "prbsmask128";
        rx_prbs_mode    : string  := "teng_mode";
        rx_signalok_signaldet_sel: string  := "sel_sig_det";
        rx_static_polarity_inversion: string  := "rx_stat_polinv_dis";
        rx_uhsif_lpbk_en: string  := "uhsif_lpbk_dis";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        int_pmaif_10g_random_err: in     vl_logic;
        int_pmaif_8g_rx_clkslip: in     vl_logic;
        int_pmaif_pldif_eye_monitor: in     vl_logic_vector(5 downto 0);
        int_pmaif_pldif_pmaif_rx_pld_rst_n: in     vl_logic;
        int_pmaif_pldif_polinv_rx: in     vl_logic;
        int_pmaif_pldif_prbs_err_clr: in     vl_logic;
        int_pmaif_pldif_rx_clkslip: in     vl_logic;
        int_pmaif_pldif_rxpma_rstb: in     vl_logic;
        pma_rx_clkdiv_user: in     vl_logic;
        pma_rx_detect_valid: in     vl_logic;
        pma_rx_found    : in     vl_logic;
        pma_rx_pma_clk  : in     vl_logic;
        pma_rx_pma_data : in     vl_logic_vector(63 downto 0);
        pma_rx_signal_ok: in     vl_logic;
        pma_rxpll_lock  : in     vl_logic;
        pma_signal_det  : in     vl_logic;
        pma_tx_pma_clk  : in     vl_logic;
        refclk_dig      : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        tx_pma_data_loopback: in     vl_logic_vector(63 downto 0);
        tx_pma_uhsif_data_loopback: in     vl_logic_vector(63 downto 0);
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        int_pmaif_10g_rx_pma_clk: out    vl_logic;
        int_pmaif_10g_rx_pma_data: out    vl_logic_vector(63 downto 0);
        int_pmaif_10g_signal_ok: out    vl_logic;
        int_pmaif_8g_pudi: out    vl_logic_vector(19 downto 0);
        int_pmaif_8g_rcvd_clk_pma: out    vl_logic;
        int_pmaif_8g_rx_detect_valid: out    vl_logic;
        int_pmaif_8g_rx_found: out    vl_logic;
        int_pmaif_8g_sigdetni: out    vl_logic;
        int_pmaif_g3_pma_data_in: out    vl_logic_vector(31 downto 0);
        int_pmaif_g3_pma_rx_detect_valid: out    vl_logic;
        int_pmaif_g3_pma_rx_found: out    vl_logic;
        int_pmaif_g3_pma_signal_det: out    vl_logic;
        int_pmaif_g3_rcvd_clk: out    vl_logic;
        int_pmaif_krfec_rx_pma_data: out    vl_logic_vector(63 downto 0);
        int_pmaif_krfec_rx_signal_ok_in: out    vl_logic;
        int_pmaif_pldif_prbs_err: out    vl_logic;
        int_pmaif_pldif_prbs_err_done: out    vl_logic;
        int_pmaif_pldif_rx_clkdiv: out    vl_logic;
        int_pmaif_pldif_rx_clkdiv_user: out    vl_logic;
        int_pmaif_pldif_rx_data: out    vl_logic_vector(63 downto 0);
        int_pmaif_pldif_rx_detect_valid: out    vl_logic;
        int_pmaif_pldif_rx_found: out    vl_logic;
        int_pmaif_pldif_rxpll_lock: out    vl_logic;
        int_pmaif_pldif_signal_ok: out    vl_logic;
        int_rx_dft_obsrv_clk: out    vl_logic;
        pma_eye_monitor : out    vl_logic_vector(5 downto 0);
        pma_rx_clkslip  : out    vl_logic;
        pma_rxpma_rstb  : out    vl_logic;
        prbs_err_lt     : out    vl_logic;
        rx_pmaif_test_out: out    vl_logic_vector(19 downto 0);
        rx_prbs_ver_test: out    vl_logic_vector(19 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of block_sel : constant is 1;
    attribute mti_svvh_generic_type of channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of clkslip_sel : constant is 1;
    attribute mti_svvh_generic_type of lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of master_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pldif_datawidth_mode : constant is 1;
    attribute mti_svvh_generic_type of pma_dw_rx : constant is 1;
    attribute mti_svvh_generic_type of pma_if_dft_en : constant is 1;
    attribute mti_svvh_generic_type of pma_if_dft_val : constant is 1;
    attribute mti_svvh_generic_type of prbs9_dwidth : constant is 1;
    attribute mti_svvh_generic_type of prbs_clken : constant is 1;
    attribute mti_svvh_generic_type of prbs_ver : constant is 1;
    attribute mti_svvh_generic_type of prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of rx_dyn_polarity_inversion : constant is 1;
    attribute mti_svvh_generic_type of rx_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of rx_prbs_force_signal_ok : constant is 1;
    attribute mti_svvh_generic_type of rx_prbs_mask : constant is 1;
    attribute mti_svvh_generic_type of rx_prbs_mode : constant is 1;
    attribute mti_svvh_generic_type of rx_signalok_signaldet_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_static_polarity_inversion : constant is 1;
    attribute mti_svvh_generic_type of rx_uhsif_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
end twentynm_hssi_rx_pcs_pma_interface;
