`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNxrMxi4iuOsqMDtcOarUdWaSJcPITiXNEl92uPjyakvZrw8kAtoVmHxd+FmCzDr
3/4AP5shgEmCT76UMfnIOGDbwlZtu+GmaW3xzxd1w4ldd/q51eBtapk70cugU3ei
sroZCQAGvHpEPmU0zg2QKeQQGBmc0zGtctkmowvYoiBpFOxbmHiRvi8F550B6Se+
FKRnaJcMjVy98R1/H/1WcodG1zrdFhxLQkcw6Ex3LlLjXtmhJyEuXtlq0qAfFRWn
WiiQEmgnsNM8TF7OXyrFDz/eRpQCik3Dqbl6V9MWObfSXwtIbbOACjpncw1XS92Z
yrrm4sgsY4yStM0lZJEINRBZGHWiwnJW91WOlNKv2nGmTmdLmxuwaISGG57wmUgm
kCnS1KvqKOhC/LtrTyIi3NmWtHFI+ZJZR9oGUFL1Hj2e0+w1a+Q9zVun+urtAqys
nMMiVD9hYPRcBx/zxqD5lyrWOdmC+8HflXeRASj5vJlsd8wrl9oLue6iCGZT8f68
wtBaRjWpaUPDSE3dqdV1cvxWVMXBXFAxc+LcJLXAas8rgWxLP0MuD236HnK3diog
zdmQ7i6ydDk+Dj7u7nqteifU+UXaayjbOh3w7OC6JuCSD0xw+HJ5qMDiww3JN9gd
Cx5UzlXco39bgjD88GiDCbYtqHKJRhCDfovUcEkerZ9bJvyP6/vlMwG54tXD0DBF
hylj5RR7OUhEyX5UBeTmOmLR0C2IsdfwJwYsejPOFG3g6vIRjoca3oVkPaX/d2Nv
kC63B2Hw9g9RvkCF2RyNLcY8RH1KwdBjAjDph27Oi3CHljS/7xGZauCbn79ncss6
hB/nQ5/m4heGvaof5gnXmzIiXPgT4g/O0tD65ZaDfl04OKfb/WWI3nGpp2lFJSM3
1DtC9zB4c2LubdnDxQGzQSet0aMpHRL8tu1bLs3OEIT5hy8PKgvwsRj6Cd8RGdod
o2AQT+oc43v+l1jHyU9j6JeVDdEjaB4fFjRMqbXu7xcNzYimZLBq9of86cWqCey7
IwFCeAonMRvcvG+4DuM3sqMubs8JVUuKOT/8hodVN37UdIoq2kGVoKomp4sUOTRM
6hh74u21oHhf3BWXXZI8PeIXPzTaB9zjjeUigsRvEHvfVlacS2zpjsBnmohllkWP
veObiMO4l+LkBh8eD2R+7H6keCy1Gw617q7A9KvWzH1/Tn38VUmROxyd246Z4ATE
L36x5ql3e6s2hHdCccIONdStdBCU4J+afAv3qpwOKbKPvwqnp2RWp94mGqXTEz6o
nDvXkalqDD2BTSUfdDDZUGvYg36Y5PYQW1nNmB9EhCIV5mQ90uL5KaVdPgaJEn3Z
HPryBwCf94FG3Mm2O868X7yS5E7pf+wmasD9xXKdLinQ0l6+u14V+X98r0Q2f8ea
f3PSDYR9XwMEHOBZe+DXFbXu0/qOJ+iIBYPH7RKU4hZlcZnRydx1psz6t0KOSVQw
YDPtgfJ+IXDulW5QXWjDZGPHnRuwmmAFy70kbNJfEK6czfbWc+Go0tAHwn35m0fA
AA2nJ1jqUlgZ/8GpOPoYkWzNVca3H28xsDj83NQYt3YbYUHf1qg11AhckssA7MOB
2FDbC00noc82Ut+FlLTpRwgPgxKFrJIApsQMIwINk1Nzx7QhyXF/PaDY/kIQ7rbq
fpZdqyvcehylph53bmgsMbzL5Q2+BH7lzuJ1IRgkG8VwCyTTOI6IXCG6H7ikWwUa
vWkYllq1hLtByqDlcWFmceFvQnppXuWSBFTWgaRt9epchX4eDrVjgfwxZ0EB2IWt
shrFZhY4siP5wUO4G2mmSYE1bIRCPkEgHUzGMeaOnOEz8XBXs1UKsXutQnKO5cq/
q03XxJZKjaKFcgjgS9FFUaWXmHJCzQAHOC0HfZ6I/dyYupp4vJk6EcXAE5R0gaJd
pOAcuWN4fpZi0Pt/MDBC9pvwIiQLeGZK47akkgmJWvz96zqlPYmejXm/g9X0vr67
ubrpnsYfKI5caRQr/2brJcLhirrWqBlAXeQ4c37JwWhIan7qnc5Lc3Q1r2rBuzf1
Oj364dC+cJgZALw1BV/MJVPtvpW4mOOmLiFg7kjNaKCVcao2eKYenlo+Vem8HsC9
VxekrWxhcj+9GdkPIlviKe/h3Wq75O2CG1EOadYPRv9f41XZ+73buBmbVUG8gPX7
aPLrtHTGWEbNQgUxRYNPdiIyd+j8agBM5bcKoB2moINYj6/d0i3Gdvwo1Ik3XolD
xTNBwjXnx8UEEjTtSqYzzgtyqK6nVkPe0sp8OZSd67ASjTyarmN0afPgGCfQegSU
nzYYa8wnvGKesEYALRUIKN7rOZDPvwY8I1ejiB/1mFfPthg1trSztCULDp5Q2kKO
f7y4Be3jgAFqcw02bFxCljwOSXypokKLJDwgLEtlz1+Ve6UhHUxw8aN4VkJIfC9P
mM0XGYHVj70mMY4cKUamfbMe1LOU7jm5CsGk04YFQYep1lbMQL8G9/24tkMHgMgh
+gYAonGEuyd6QeGFyBw+h6gP7Vm/I1lxZM8KWP7xYn2t9WClv8ZKQb+VJFRCrItM
GSnHZszqVy5J3jFVZ2q0RiwmavQcJ4XSXYMbSKL+oTRGZU6I/B8Qut9X2Vp0rdYz
nGRvebOlksT5nwM34VumOO0yVVg6h5THTZgM9mEmdM7ARyLwqaNuHA6FOVKBETgb
C5fGo4QpPWKlr0+x/PULESY+sUBu2dIT6Oe5VYjCBT9BinPpon7SnvbqcalrZCQs
Mg8eCXTaB6Ut+SABT73pirHdUIneK1ER/Qtbit1Fi7nkcs8D+4WNzrJeIci0AsMI
Gqj3CaO2vOHfX7Hm14Qz/BfdDmYU9zbn4weOkxwVqdgLMwOukERwN6NWFTqUGc8U
ApNp1cCVt77zGiLn9jOMiN0cBZ672SX/f45FxO60I4gc/yswjhm6GtU1xGTsZPaG
cWIcD8SdE/J6+QeamxbYy1pLLwBsGgq3IjI0KdQGv3l6A2k2YOtGrDUTGh6t9s1v
XlG1aYyOLX4XZ/zGhKtfM1t2MJk6mEn6StR1nF0vLD/s1LrZLGiY6P3ZI0lLQT94
z5rseQmBNAX2r2ZEr7xidNZFFPn8KVQVJYqY0W2+ON4UBL57mPSVDGilxUnJ6WaP
bw1Fx3w3C3YGtgJ1fqSM5O5r+JHylF2by8+xuOt9ZUqL58+rVEPHz2iXolXa91Z+
/t3Z7be2CHyrpa3mztTl39yBhlbanoPPBx8ob+Y4HCCH3t3wInaOvLL3k6xJk8vH
OmuNY6zPb9fQSqumyCm9ixtKoc+27PRmVvZJOGW+tC9AA4CaJPLZjuqWkgv6jU/w
FqO0DDzuf2zxBn/mqm/50eX4vSjsNZ3tsqwyVfl2RzCWIzWC3UqVETL6PtOMjvNK
/HsaulQ+xG4uOxu8m88yI7fgf1dtnx8FblnH/V4rzmrDFbhtCxFl/pUEwhnwz90W
5P+LWgAd4d1pSqAAvheQMo76CbizcdevOjXmB4Ly53CPR0aFhgaq2oA9FLw72j11
Mpx6l2fqnNRAMciIFP67lVcKot9MI2bop/lSzazRFZ4nGKR5K4KV6nAjnvn0RRrk
F/b2SZMOj+SXt57eiRCbSxau1yu8a0DSyDXooAab2ppOB7oIMmIt5K0npqon7gnh
CCRpJPGN12TwIprOavSHHMZKToTu5MaZbucTlu+4ba2iNGMkOATpYByHHEdOXmlE
7+AUWH36NOGnNvUUyi2IuMlp3XDGojw3l/oACjuOQ7I7mAZiEFWKkG0SH047L5rV
XagERNklzg//HmS4QNItzH8UTAiWvRENTzkYgxzbQf8+rfJQab7xfNfqH0/iDz/7
2YI+S5hSyZrTiha7SH4LJUgB1i9+YjXYPKPdABcXHShZJK8aqMhw4aya/Y1pZ3h/
OEuHWDpAvcPah6D9jzXvxHRyYhZk5cEFE4EFClW6xNncqOlBC66y6hZ4stCeqk6H
mQJAPaMxMOCSlx8W+TGknqLzNrHcsv2c/DzcW4D3eYC2ecNOtBPNZGVx673y3z6s
Fr0tpoQCDRVv8i/dxaa9il3XD0Quj3BX7eP473kd1CiQs7WgTQBtkWgSLYcIOVTL
MmSPBHOTCKkbewqrr2VWPVwrxgm1+Xtrms4et0T1x3x9UWZo0VPr9sNYcKdBK/jn
T+EgHhllx6qVDZFHwSwVLDUD59lluQsmbEbjJkGkuGXKlO9owMcWo+W5HtqsUjbA
Z7Pii5iksecIThNwagUU4gE32GcQ5B+rpodncWAk4GZ48mPNSzzKqb+Fmis7oLbh
gtoRkrSvfQuekki0SB7+CqxmjRW9Ot0tdIGdSLXXCIkXVG25N7lJk5h0+Zg/P+fv
qQUJKkd+KQ5YxVeRR3MYuMiYLONbm+luvD/UIKZvf6lzAbZvBdbDe+8wT5bpCJYv
vGA+V6NignuM7nOHpefoyW8/ECPelKrbM9ucl8NU5vHAxV6cBpnxp9+dGeSzEAHu
+e2lavrSBJnHm0MAv4nC6gY1AaFBZmuSV2OwqeIODaHWlOLByi/CjDunpoU7GUBD
dDTL5oRT8fRThqamdZmXA4CkHLaV9YS/EewlBOKwc0UfhGjs12G0YYOBy8BshY9K
vmMdmon2wI+HOAn/5VoGj4jbFDyj2pryFWCPbhcza7jayEi3wjEEhVzY5VkZceht
APUp/AxExcA/zm75CA60HfCY0ZlE7a1GYg2ct/PRXoLK4myeFacKdXktBJAMhT40
tBNFKD3Rh0Zum3YGzw5HpHPgngVMARvFZJ78nspqT1yFDkGlLg6WYQ/NWrkpmT8+
VDPBFvp4Y/OOSXtlwv2ZOMsjSk26zVVe9L6o1Weickh8GTjHkDxk2U/FqtlzAB4e
c9MtW19SuHUDR1jvzE8hNrOEpRgcpo8LGbpSvUXj0+a4hd0QPWSU4ROxr6pagiF4
19rx5nKi4FWkXBx71E5hIJBsoRS/LrJkNZWfo8x5mX74ujk2loRWply2RqkB1RDS
duVUP3wFYDg9meakHxYwV2AipEvy8qZKWljd7yjENjf2yPUadi0a0GzeXvnx7nJ2
RlOCWYgIL321k2AVs7+cthA29M9D2mff0Eq/AZxegqBI6tz3JhXh/Z6jXFSR4fMu
ks4j65SVqIYmyAXjBR+xkCNqQK75/SHzC8Z9fp9PnbcQwCWygb5GYEcLPRR/X0ZL
qSdpUzD4YojKb54xh8aOSyuJryK51ehA0E+n/cYz+WATCc+PDyCpIA+F1eJjlMCY
+vTIUQmMTwrouzrYuULQuPDpBiomhTbP6QMdMgSewsxG+rMRMny27P3YGpHUrfvJ
ADoHIkYC2R+BumqvQxOcDJn7DcJlPcWs2J9b0rjOASY0pwlhF7VX8xMiS3CmfCsa
bGsF5rw82B+7tTgjf7oV8yq7tmii/dy+xdcYJ6pOtl1MzOppnQUSjiZcfzPyVgpn
RRGHljYGkT89SinRyjfv5JUClUJ5P/XGCTUtkqsAwhgXwfzcUkgGrtU1U642kS6w
5b2bRbEuYkkdqUbbvGf0NUoIFcfj9ayg3nQ/yBzp6lSc8P4+t4DmKxaGWfXNzYuc
iI/W4zxj1QK7rzklD2HVka2l8kBkWPB19CuS7eFLSfnY0gp1vAM6UoOZrKCBeaHS
VTdreE9VaE/X4dEw1x2iokLaprP06yPjC2sYaMRpgrUqe3H4SqSigzffJxGsE3kw
vLCdVi6i2ufNikhpHgxenxUKC8DiIiZCAmOu8rVDJ606NYqcURP2q5CWwa2A8KOz
zlvftrMq2/yLXIwJIsikWC+SoPSnMH9zyGMK+FB+bH2G4pRDaplVAJ7BYgnEXLj7
cM58yZ+uX7YjF4r0u4ezS4VpBXtzBDT4YpRfnUzTUMRD6myP61m02Yeq4gIeuGSZ
+jr2VWzTHKcIbzs+yeuYT+srpYjbfAhmODomBBlmeBzwoUFRn4BC72NM5mTOWI6v
znRnycQTUee423op5bX1XHzeUhJTzOZe8qW61PT43azQ+2uVk1YaZj+rH5vaMh56
6AKF7RAOebBvEYquil1KZvVful/kNcDWa0CMzkO9hbFrm5tkmP5xaL5cQYpK3g5k
3UHYpEXozfhS8cQKOkR95PyOjMQlMWiMHr/RsVWOKn+qcA33uhCZuDhXksRM+MAG
T8zwJWovi+wWQVgPQ+3trXHBSzx618goaa0IzB6DOYqS6VzaBgKFZZHx8d7eTBm5
7aldAbS4TTkVhWY1UIqDQyYt4o1kmKglar9aUPDmtT4LO4hD8w7qacbuGbSKTNgr
Wl2JGFrFmc7Cf9vpa2lzAJ9atPvaU3Y+j2ONQ9OVRgxRWhcMxKSEwlICFpR0XLtp
7iUTmQBLfdl+kVlhKW2x1hRem3MENpCxNFO+/TimxvFaKhrPCy5MPOyDS4gKv0wf
OR9eHzRgqWvpxCSzc+6XOxocFDwevj6EWAr+h9oGGtfku805EPezm21tOcYPqotQ
ks1NI2se4cJ1xUSTFsYJBihXyrMa4yN4kFe5QBuBxj7APbQIx/JTDzivkQn2R9FD
r2Rv44nJ2VhqQTTgDE1PBPzAVdvLGxA8uwfrWiryYOe/a/IODk2wuEMxdY6PG2d5
HO6be2kOoK4TQYlaijEOgxGv2gQ08ZGd9p91spfNruEgP8fDUCcKlSsMpzKQXDFy
FkBjb038I/uPhTSZ4O6KDcofMubUINADQueT3f2feol4O47eHSZtXmL6KzoKFcqu
9N1mLd2clcuf5oQvClQ1aRMg9qVnKYGzNa0IZ3RaEUnykkbYgpQpdR2QeJ65Usem
WI5ft4CNiKCSHCPLvxeD3zvhPSDADMQLlN8W32mBe86PzVOicgwY8aynE1tiVigE
TUiW9QkAc3Xy0Lo1iVNOef6OJ7W046eRmQCvogyGrefteffkeDACN0pAF6Qd1G1A
6myXPLqEO4mMfqix0CGzx9qzWIVoccpNfsPL0Qm7352B8pQ/5CbEo+H/0zNAjqPD
B55aumdbCXyJjWWl1mKoeK4Jk+vEAGQsX1nTxe6k59Eh7bbrddQ9KVo7euCpnyHG
me/EValoh1S55bah078XitQgU4LHAhxWN3H3p4Q3Tcu5hxuKrLTlABt6S5yN55wa
ByKCRXATHCEfRSliYYhzaQQWvRubl/UimWu7RLH1IcCoS/MVM72XxjV83qhjGats
ClfxycQJwhwvolbYucd2MOmql6Bpj3UxcE+2+7mxvo3sfY4REq67rJRnHwWdglfK
LHuvbKHxuWB0RLnUcStXltqChzVe+EgH8/q5CEWHtH5GqLXyCLIjyPKXxsfRAEOD
EGUDmiXsnpkNtEb1DnT9lTdGtvSNX9xYuJL5T8NA3Z65S2QlaLKaQQFTI7uQZ4Hy
WOw2oAwQZ0blJuDvl/22wz4rtqf741UzmsH5ZCOQU2BQUupIdNK5sYmWdr9JAoOH
qAHULGkop5JTglEBFwxz56ixp8+ljGqLKxLJgP4ZaP5KpB9KSoygcCbVsu3PqRF0
2H7jPvmPdjQie7EYmfSBFX9duCHUIylvCd+FMfrczp7GxAx+KoFGSIrdA1A4t7Fe
RTTwgxx2uN2v/dNjR9At7oGdxcVmidRJt77ozAkH01sXwDmf9OCGpGLkN9wThf60
USbMc3y9qU8nnYbXY0+8sKe90KTgGdvO+rye6NZtgOw0+Cu0GRtmuO/oPXTtAqWr
jQLaPV7I+h39GBiIaCSdRlFPH5LCCcJcqdIIDVkQfwZNlB6IyY0I6OcSUtK1mTUD
rz0Y4/VDjxJOUeRUa2lJKNlDMK9WR6FjG7ssulUwroqXc2D7Q/keaGHa5WDwx9Hc
WDE8DKrmUjHHQORUqNMuNsrlPm4D8pOysvTCdMj6wdO1GEcA1LEPJjDGlKYNpPNC
p+sb68hdQq0M/L5AAQW3WEWqBb9n43RlRVPJNyuA+Dew76e8TcBacfDlfneT8b+C
9bJdcvip0AqZf7N88iTyLgfQ0KcQg4kZKcVsYxb78eWTXYxl+snbC9EgMR2l0frH
Dc49yKsfhbQA9SnHQM9YmJNcX4fnVdzpMyyG41DrNFw1tludv5qoj3leZpm4tP8F
/UimR0JgMb/GesY8KIoWhOXmb4IeHqZZt88mSKIag3HseOWHG7STbmziazbFTM6o
zmGONbdXwh0SHMexIntoMAHOQXpiP6fePyLtrezSinkjMHt0lkBrKUNhvONjW1op
YP9iTp1CLNObH8z84gNNIrNf2FHsvAXOrTiBgneTmn1kB+00t/A7xBsoj9w4iry1
QVIsgw6w91jGaHD98A5EZJNrA3fNjZJYcqXHndme5BNYi73/3sHJmvhrMT8Ty1U1
iu9gZci8wk2Ct/EzfHJyVojbreL11Mae/y9Kh/TSB+1mAs3efVSjk6IwWPIJ8MYP
hP9wRNw1h8KOgG4JjPfnayr+TeJ+rDOLoIYcIBubGOfNWpXUG9aWxqFoq6OXxCL1
wWs5G5BquywZCgMYKvdxJ2gzA26AuaTrkQpWJcl4qTjFKLF8ip9a9OwGxMat416Q
a+BtmxbRyecUVR9DZx2/vkjlPRgXSytNUOoDgs30xGM7frlox3GUWVhGfLyiza01
aNKylWgHb60gUYvshmGqjijoxaqQpewZ/Gs/OWYptjZIktfS0Fw4RIL8Rik2ykwg
E4CigoSCQ/9GhWr0j/8utMTMkLa6vcBqjU9V0NtehePbrVTsN/F2kJELU4DJbDbn
qZggmqYv4t0u/q9LwY/gxbqKbygQfG4DL/FdaB9P05/U8H2qISCSBhte3pCIbXKz
Bnm6sgz1OGwxQtYuAaZUELZbQoYPW8Zr7Q1U+ZQNttNZ2DKanLAddYepiR4hKQfh
R+WGaJ88/a1DLEkHPrCF5fp2QItF3dgdT5jeyWkD/3VzZBeOOt3080N1weNUf5ge
YDvxPClVjxr06kksTd/EDIw9yywnG0WOmt2eL9pFSa4sWp4+5V+6WAo38Xs8qZta
tpA+9aBu8jpRicGmxShJXvUov15RJKdGPpozPZ7Vzdktub2MeInC5Ewqi/05onfj
SEJIRI0WwDX4TWfSxkyVfB68FpT5xyoKDqYQmCy19scAvu7cdHGbQjJ83+o+NNie
N6zYOvKawQflC5COCjbIpizbEEhlWOSdz+bPRtff8uOtCJpgDM30LtJDtt1zRi0p
HSSiyr/DmzXnKrU8IHfVrE9pw6niDaTqCSmJT9OApQ6Cx/ta7+btXTii+1W+0vVc
fdZetJxGXSQhqWnLTYmL4t0lzZtIBuyLwpb7e0jM8YnqqGk99QTPfli19DzOs/l7
oVmv3STmfszzM8TuXkN62398TK00hKRyLB3HMmOPymKEDD0CaXvr4QOjLLpHf/lo
8abNgXB+/N/yT73YM9vnkZ/xDgNiBTckjnno8VcF3jPwCVLB2/VUS8SRQfQaRKDG
84veQ97frjZBsK21zwo+D+TWlw7TW2U93tn4p+LDWEaas+E6s0dv53i4NO+90P+T
kq90vDsz/T4Qq4kTO74nZUOA6n/YdMAv++4xqynix/4ZzAouPEMfvgS4mg5Eblqv
Y6B0bWAcvqLQRF//N3WdxAvKBSOyEsKWVS65bT5HsMOkIQDc6IQ+OGAGU1KzV1Rd
daiG7FU96ShAmkb+1iPmSlx6DZV805kHwQg1RZt6soU0LRV9wWgoNnO8JSkgXYjB
BtW9XE+1VFLamqQNT3QrbA==
`protect END_PROTECTED
