`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B/aOn2/0L1Ezht0ciMdUF8/0e6Ax6t3xAblJjNl/VeXz+MevXlONEtzu/GFSfAGg
Jk0oHJJ98gcxbcTTax9r8UdHA6yQTG0vl2SDzbKO7kCMM6bQ8psd1kySZhqivcst
mcWyd0eZJ3uCgLzu44k82S7jAKZVoy5ew/5Yv3CDZI42rJhMOLUqAJd+O6EiO2mA
cx/XgancGQFYyP0hOeJhNpiIjLalo0PSkeEJQ22fuONvepkORnjq9M+rbO6WcHrL
CTB6pmIoHjZYqL4tZm3kXmfXcPowD+66K5o1bB95gKpKrKxdoSZZ5bBHUXXPOxDn
CwinPr8yny/T4xs9G5D25+RwB+kgwLTLltqSqRjfFCF34KSR5i89f36jRMsfQO8Q
XTWbMRFBhbEADfts8Yw2b/YdesPRsAtTARDHi3Ht0ViikxmUnqa/2xq4Y/d/5A1i
pE10A/mcYBkPAfrKsOegftQCF5+vYvJA96OvzN234MjguZg5yvl5Tt8djfMEpToX
MZlcOE/bMI2BMe0W59+J5MgUuDn8D4hRD77v2Y31twHELb++6+Jr/FFXblpM+hOG
8MBN0W/WdLfMCzRFmVzY4Cr6FWiJYqmcG3ohS724MBulBwk5zZLRwkMJF6ie6ClM
+hqgBx7/6Mdj6p+9KpyeOrPihA7rwFarPjtz7JMdhRCsaMtoxudmaCnVko8FzvcP
EjzRDIQOBuHeDYAU9ZX+vQvAIvOwUx/+ozY1DI4tx9cwx4NuEi0HH2O7BMFtZx+y
WqhIeDCMaT35LYgvA+OZ5UMcPq+WlXfp+6+RrRGrPpeLSmESqVuDGTkGlH/p284T
0C/LnMJ1V3Y2z6ZKAqtLPKxGnUZlyXneNvwmC9/lT7R8SygHRqNKqLALCBNHA+yo
Xk4fWu6idh/+HN743yVCWA==
`protect END_PROTECTED
