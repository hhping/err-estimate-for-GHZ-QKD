`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bP/ISNKQkRLD7R54CSPJSZ8aFNdgUQCPGIUOkRNER8ZRqXyfLGsmgn6YYn+XN+mo
wVGHrX8zM0HBaxotyPfS50TTGp1/9HmXX53Y2zO6iY4iTLnu3sUaP7lNfBVnFZ5s
BDvjmEwsTEzkN6CN3amKXRK+QvnQfDV6poreAzbQpCPMTb0y/Iyxe/FJcpyUzl1j
Z06jyrA+D+jzn8LGFW9Ci8BvaGWvJ/BN+/LoVrTl2M2GXqdrHkYpmJvahHW+GcB7
hJXpGXmMDOG4SwcanxsDJUnx3Vqk9xDACObQDurFGh3D2bVUC7hWo2dWAepaLvAj
atMylSQa7M2W5rNPixpBjOp2n+NcHjvC8gbUfvltSwK2UBRobxTxeylOY4GQvWne
lwEIyQvUH8Qvk596aM1p4HSx6m/wF/THLpjTLYjf714jUoBvn7NfgUf8ISWbq3uu
TGN1FszjUgg4DUfT9wPkfHCJrkagaXm3fiN7ezemJyZ0MWFtO0lA50N5eRcJ9jbo
oxiVezrZ2tvmMjTDZjEKCGyMRiACDyhdMte7FLUbjTQzmngomgCVvrciWojY65LY
d5D2thhcI5s1x1t5+2KELYpSLrIqXrXD7jfWSRnbKsFhOlRsBTpKOZXslMOmEncU
sFDQ50OAamrpokRhqlSq4OS+b3G625nhGZIw8U5rgCMKey2YH/Yv3lQFiRjnt51L
1aJMwItaqEfXxq1JKLBBUScYSdyR6qec3tNrqpiO6ihTvkI9jyBXq3XZFYmG2FlC
rGoQ8Le4ToIxy+H2jeUDaJB3VEYavpfia7wSbf5bwi6LzQBTIlkqHcLVL2qtofKb
+8/19E4QN+1BJ3mC+VIONneuVmB4hTosUL1ARPKCY9HST23QyrewDLAjNxskEMSJ
u6JfocequV7Yom7Y2XUMR1pSYGUAXGQ8Zd8cp4E3CU0brNNRBFYmyYRoBs5Q+tk4
mRx097xVtJ91TxnXkE6+kNBfvkgkc439nZ0MBEEgRoQj254t5kuYnJ8xu4xE2PK0
EX9nBKuiU0qtwJl3tdto6Q==
`protect END_PROTECTED
