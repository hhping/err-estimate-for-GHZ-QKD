`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QIwaxPwm4hm/Ax0YqwIPPwwnTULDfGv4kQ9S3ViG+cizPbaDA1FLRRVh2aKDgGNQ
rwWwpSE60BtG0GfRou3/lXPyA3Z0C7SqqRrJjjo2epjS+tw1EMgKC7574irVHA/g
cRKInlgksawbwm1HrD+dmt5CB0/B9aI/L98BHMslaH7aJNnolr5yAZHnHBbrEWFE
qfLxX5/Hk9b9vAuAY5jVv/lr6A0zwxWV3nesR1hjMS80lbBHabz8wbQIuZtAttn7
qFIK5CsPtoM7SFK2BCnhyIyD6/V3qncmfRDDPqqjlAy4ItPHJbbIAUooeoeIvL83
9rnjbXwNRMxW0R0LLOWidrVlp34p7U/HF6v9YDDXpyUnegK2+EY+KNxGGBbRJdhD
iVdQLMQJle6vP+3sOajtwOl00cUyEyNkgm2YU4Pn/No87mRO3b2vxWQaR5Mp6QLr
CDNNBNB+/oSUOBLBkPE3WOHg6btmRaKM++q0C/tlZcQTdSZrsQLvEQk5MK3b1h2D
l9VQSgCRi0R2mbbUjolPRngTHdZD+5L9guaygIQUj+vn5XX3d4+fXkoDRyv07hn/
17HLaJ2q8xB/UmlYjwJhmAxpdmpXeOmA/qwXzDxFlsqZSByjjZurXzmdcFN5+cjV
clp8VGdwHj2hy7QBtqLeM/30bplbatQKNykN3YDf1+1dbrWQro2DsXs9QqSjhSLy
SlUOwU3BlmDaHc6hxydprwpUzoNAAUmxYWXHVV/CxqgUbTbgRqAFHaA/IdmABO/9
Pu1QHZkz9KJgrfMaQkGtyts55YN9afB+fntenHRsUDyjQZbVaXpYAUNjHrdW7dIG
P+cG4W1KbEgfV5GjR7Tg9RqJBr1dGGGY4Bqg8/um+MmZM155/5gcAUuix5dsJ2fJ
WkZ2Vx75rJjkcd2nan7RkI6ZjaCljny0Cmlt/XBhhlcB8aOuEOHutnkmoNc2ScrX
YDVazQ70s/+zzGrVZIKGZyK9xzTusHKglOvpqwp6JBl1ZmyLCSWxuaqcltn7TT5+
ysbtQTySeCwiID75oX2FkPMD4v7YwWXB2fQazGi7ot38QUEK3BW//dsD4+yQ2sgn
DRsYRMMNlbFvnbKeo/oywmi6N7UfsFBwnbdnjG07i24hkvQoEXPbxZm5DhdXYCrS
qdETllYjCdJEhnhzIIGhiowkYG2utum8zQcN602nUTAO9dnbPIVJbKhJF1S1MZ37
WmnHyULGLfW51nsW6rxmc4KBAhiLxxYqvqk/SJ8mF3lY2ddoFQ5jGjSU2VSJZ3nj
nfvQcjAjrGfy0z1buu0AMwHBTjtApmeajHO1IFomfakyJz9me0movfzzer5hVOiT
12q2b3sTGj6t66ObivHm9ujPMRzEfktbEqUDYo/SETBAeirpWts0LE1yqiVEfV+e
kmjqfcovTi3BtOwL4MAs2ARbIa67bykXZ5vxE7gtUCtWaAKUtWjzrwF2ByTqHyBx
8ECXIjHOBp+TXJEsSM0ui1MUdQQlkScNZLpuuwTnw+dryBERJxUGBmvctnPRSCI4
rXP+XvW0q1jE8HgNUYA0gPn1cnf1MhHKG89ZlHEo4Cw5R1wKTmEg9a4/nRDluLl7
LgYC2BrsQLP64K1T2VsyDOkO+ETpcvgNOtRUaUJwfkrtuLWKi+8RAO1c4zdPn5o9
/X+ycx1dXqX84pxNmzfg6L5LAYm5VS+7cxM4UL4hCoI3QnPesQ4HitmPfFXITt5P
PlHjC+UQKVNojbDbN4y3cpM+kz3Qv3D/de0VBhX6PtVEcjdke7Nz5804TLh9xx06
qrlzNKm0ddTfBeOeZyc7jsXPPAltdjjEsYdvmDqsQMTaqnPzB0xDPEU/L7tzth5w
pv6MVoZkKbx9m9f825yaQGQSQUUGtdlRhx7NyaNpciKcggSifdqHBrehIu06sR5W
TB73GgARsV4v75Utax8iREIV3hZjdgdsjald/VTfNgTItVPtgMdeyMJBg5jSjJIL
zMxSoGTBXBWy8GtbePIlxBv6qQIoD0VU9Ui1OdhOl3T1sqHgAyAeYElIQWgn1CHp
ixVnQmTQjJGNnFd9cswJhiLRtOEuP+AZpfrKJuRmRLiIGdoQsigtzds9eiv54zk2
zmLqCRWik+ngr88lkTwe06XwNtW9XiUmBhyR2TmgLyj3a+q2J7gl8PfJ6q5jrIc1
MZ2SSDxP9pVCaC2ahVafWl/WkG0JFY1pB1pfPOLb3DnpBW9a7QEZxkU+oNKlsgzn
R+1EisqF/TRv+Xah6wz5ZbY5OJ+luCvolpimzPFd3SiHV5gqtPq1AJOoR6Wbefiq
wPy9TpKVVuSJhy7tfu6lqfyVtHioL/EIBN4UUVYY2a/3CJTtFkjDi/H1cZpLNlkV
BWAYWVCD0tS3XrFTdYEsgbDgA9k0q0N4yEkNzd8JqlgORmj3wdWMei2jbWZEuRLJ
SCZ4sggfc9t8RQJNRd4Xlu/ckrcVy1ckPUKiluG05wiOPCrFfQ0GX6mfR5YOKLKq
4eODu/9HCJdkZsckULS02qqiMs8E7wWdAA/N3pSB7Ed33FpgA8ApETO2dXjmfpOy
P5x/7Ywn3uxkT52/GRewkDCM7KTaZxS972NFvjgJzc24ubEBeJw7cbrEI5ZJxRas
B+rLGNuujvsxgahxyCU9WEuluzPwYlTVz45cr/Dbd6uD9acolapyMruyWaRHC7rn
naqpmzud6vSo9Qv7/VxNLhPHyD0YjRi2uiuCxxXYOWPtkJiEbXxdkN5PrU/6BL1s
o9Ve3bR0ce5jMg1e0+fLs5t0AdJqfr7bEIgTjJEFkddgYaBySI80lgyZCn0Jt+H9
WmjEcKnc8UcZd7GyIiDlgYkCHSNNXXDex8QnRJ91Krkl/hn06DYLnWx71j3yPiP3
I42z74n8y/76b+hHQhGlD2EJPleZlWlYJhUEz5e/qY90oxoXSfX8zHvZZI0LaAUx
V02JtT/pdnMrMkVcLHUAC+Bx2Q1s5IABwpyPxWs+PVRHEmZRTTQkSHjZH6LLnduc
Qi6SjldrhN/AK0hC+RbDiMqB1LdNv9r43gX1FisgX5Vy1V6vQ58sI7hU1tlH0hSK
21pbGL+CCZgPJr0m0FS7GcAoUGgK8aqSM6MeP9doUG8ghesVsFNeKm7dysoCiJw/
4mWfm9Qqfckyj+o+QvVvvaRkPLiYVPDblE784HOvCgdOqKfDAvo5nLyKauJzpXY3
6hCY4c4AUpyzPbxMGU+NoE0tibK+yc+o2oFNYs02QpbSt7wZwzPmZOrGTdEJu9gl
ajWgNZfC4KmAYICI18MGo083UI7YX/o5478HeCqOQfrBzIdnHTtkP9gc2UygXCy1
JDRKHWZGOJO6Nr/jOIGwSm3yt6c7XEkFsq6Iuq0LLXtfef/CUZxSluYaZZwPr5VD
xrjMVVtCcm6oaxhk3Tqa9/i1Oyr6ViP8tnvKwoPN7P/wS5+jvwjpP8ZCde4OaPPH
ONqF5DVOhKcJ+/l6SaQkYaNtHVRjKsZthxU3jOKF+9OuqItsUN02gD0UlTgQx6E/
ms6bUOgIhgg/aHphnHM/3key2zurjfMekvERDeTI/Z2bGLTCk/wyFfEHB3KiBgRn
p85kwSSjeptG2bkttz7Ow/ImbS95h6O/HtwmglfO45MIeE5iFrwMaHwWXi+yvidr
hd/ozDSSkKexty07ORmKwMsXoPdvYBPksQWQcGPqgsTnsNKjfQ/fClv1ZuyExFEF
LD4gvbGgVNtz3uwyUp9tjImkkQgnPMlZgE6a9ONwaXdfoTpLPMPxF/GDDrlDwP1B
uZBrWDicCSx3x0UtXMRI0uMk0sRg62SpplB1PgIRnD7xy3wsfhtk60Y7P3tS2t92
cbCBI2DndD27lp0/P8M0h2FsLUHTrKuvC/CuvWNURallVbI2ZEZCxFecBmrKFvDc
/+Vm18DvFFfboYldY66lvlPRkLDuOJEI9/MAfWHGg25fWnhgawI4sYem0ghRvRKd
IX2R45/Tx9lLtYoPng8lNsnTxsOsk/yO7/k6IaQsSn4PX/GkDZ9D+sbk/V678P81
PA8Ge7vqg4NY+jkLZ8oBJuYxu4yQvba5CihLN7p2gtJ6lxnoHlPd9j3fwIAYTwAA
N8Mt1a0Wh+XEQscbwgFNWKVO9h2FSEpCMZw1yvsSNT75LqyWhvSXkRiay6NTbnQ8
M95faVJ6tMF/So/RBauoiAvs3TYtZt++ETvcuxSBZsZI2WHSyKvuTZR68haZE59H
6Jc7kuLYDfytyZCIfg1hZKmOgKe8MuRwKBT3aTOfoKbxfEElN6qyX3lcW73vC0fk
NHxqMAgdXAiVuyChLNq0QTQRhitZ8dJB60PFwSwNn7WAJ6YIYHNAYn99wHUcpPdv
Q1R1rrj2pBOvoTFrZICt42v7gpE5BIMfcLAqg/oIfnc8LVSndnhF8FG8G6aTBvr7
S0ehQnfWniJIMQP9PRItS2ybPPuoCxZs6PEq7eqVoiIAd/kJQnkD82k+h4iXC5HV
2zW5pb395YgerDvNQT+itLy8DAONnZk7dlRdkBX7unwMlSS8hpAksFw+edA2qtx7
glq2//tIDjsBGFkTZjMvQ8FdbaQgkgwPuZvgH+KBiWna4VzACLZ9HLu+qts8R0fE
zBZTrEx07tMQxGTRhNylA/crfNOy8zvMY/JtliDC2q1BuvZpw6+vT/0IlyxCcz8d
1fe66L/F3r69mx5QxnhIWTfORutEClWv06a5/L+PMQcVCBGU5IpCIFZxnwcWAjnB
UOMHw/W41i9IrQnIODH7VxY9TIgD698IYvqzXEMnb1/J7lrx4UJLLXmYLHz3fplA
NLS5SWCT654fqLKxHL5bafLaQ/QIXtrsZNJBIuRyM+XUfnTSO0nuXyjIizNL+uSR
jgfzMPxwzwToy0xCfAMyPMns+cDOeRxzk3N9YtvChhhFZtuLzhAC1lywCKmGS3+T
ECP2hSzqcoqH6VrMcy728jkBtnsTUrkZXpEAf1cowAmvdDC1UWe18jSrl8ZQ7kgT
iynAO2GAJ7h2bbC/4tIDIDbwq1gR+F9eFgleeaBR2SgjHpZpB6vHehOi8ZS2VqW6
XlchFmDZTmtVzAUg33sALyK2qGG5Z3fLDMCLX9kbjGc1Iq8ImnCFBoDioJTrn9gF
HgKl1hJeZPt2eVWC2AbyTKEkbnW4TxgvbNnSJ3Fglis4aguGUPhoh77fD+Xx20WM
/1OvXIpiQ4epyB8RGOgf2wkbGtdK7Pc+MjTznEqcBuRylsdfqiH3LaBTQgKb+d3K
i6+H/FgvH+03XNcp4J4/5XC+FPtduCLDdgjdp87Q/GaZ2bNRo1y91SonMQ0F1p2u
Qxw2rP+dxOw85A+fyroQd8QuNulGIZNVO1yVoEAmkaccuXYLZk31OE3UuHy1KGLz
nIEX9ZSf96STCTH643rK+dmWAsdDQT0xzidugl1aZzDW/7dwf5KQPDlGX6AEwOtJ
S3z9VTlk1Dm10yKdn++HNuh8+3DYLbRJd0CO09xnY+mKJF51mOJw+LAqDEfoqZz/
DFrTbxxBu8S/FsmquhNfsCXFokVZ1mGbZfcBlgTGYfXCfjmu/gelBJfq36sGzNH1
u6kV9rcuHZnzPUFIWJvDXs+mWNFc8V77NcFzX9BlXTf1Gm3htsIKml0QPT0Lqumc
U3mj2D5neU/GyBVD8CHBeq8M/a/agj3kYHGMFDvS6sbvZsxCInLn2ozYFIynRIh3
suaJkorieZDpVXdcSxXitDm1HDPrLVSsNIkH/O4HIs8Kempz38bFXMuVoCfiO4x/
45mD1EWMqqA/S3DhZzwQTo3QaOIQBfyVyqDDqvu2a+R+uZesvqmNHmdofPvD2a5P
OxkBIEJFviC/RsbHZXivAJF3MmvbjvnRj1uV6fnqUKqCC/CSDo0K3Z5vfWj+WG7S
/txTZVyZ7cFTOBW9m2micmsWj6h5pBECWnA7/kGOOsEApzEGAVPzvK2BwdkokOf1
+t/tBn/i1Al+fcqAi5SaDuInxAJbaBpnGbfjolOkKxla2V2rK1CbeiwIxhwQwtTu
sQEJYGXmLnRVrPj/bgw02vVAvx1QCF40NMhyINgCmY9xhv0X5x+3JVJwnvaNmChT
6rmlEoE55F3toM5v72oUka9aWBH+VxhEh/s0lRtsxtd325ZGogJm2IMbsqnRv04S
dsJmUWl2pTGfYgeXd4XIYRvg3+X2ROD6RW3GeX+Jxo5QhkFApSHqT4nC8WLHwPAU
lIJhy5e8QJiskc3laDUpbrzgfTmUVy9spEAiJog3B2LmmdsHkowTP5K05O0NHiGb
wahjpSp8cpqlqLImNRc7GSfoiH6dcUEdL2DOoKtP9OrgOGtBAlKX4yv1HDCXnQFj
TeiSREFUuUVUrN1TYLRVN3Z1h5SE17DJ6ojgLIjNaDFE8GgOumpXFi2aflpcOaR1
8nzqDavbrtTIdtoZ78IlrrC4EhpCIrHt+Hv3wMUYHMuRQH29y00PZStkKONvT1Sy
HMvoxrslaKmIFrQjSZXCDAvhJvuqf4fDezkFSmhPt9xTV3qkDPAMZC3hKHYTbqi4
/gz3ay55c4LPc0L4N//7Ln+uEd3PTxdmgR81nTi4kN2sWYBK2O0lJmzwvp5bcGiA
o8XAn0zvugYm5qIGtAF8qwc3yvQJei9Q/P0z+BRs1MfjAzHhTMDLRZ6+jGbmK0tE
guTgdofvpi7uYf1Z9WpDyR94O3jgEFa4QyXg1zqU0w87XGRjgeOMKv0uqAWga8u2
bmMeFmhjVEcvdZASfadBrI3vHM1hB55JWXsTFfd1Sxc/3/Noax0DEySBbiY2Uaqo
xNVkQt0wnUk4m2uuKL2niij5r5b2ddOS2XG/JosAvsBWiAmeR/Xo/nYwPpOSuD22
DGaip5Sk5zeHkMfgwpRwe7O3INXsZREjtVNZ5InTXJiFxuaMxtJ6vNgpJzmDTnQP
PHfU27ZJ8nB86QXoGHxYPR/RsCqOr+iSwLcpYHVa4UbilggCuRPHWcOWYQ8kXI0x
YVc7nrco+dsf1dBl2gF6fWEOQJiy4QYd7JVVltQVFlWVtqwC5EWLnyICSC9ROe8d
AuoxnyIlWBx7y6iGjEXdpUruBcVY9HS2nkpBSWnu+8WV+rmhRlcyhziorpDtNMqN
RNRmRGqqBFGoeyvmUUfvdSHmxzqj6eMVZfZDdNjiPLp3Iwhw/GwHsGQRptI/8HES
3qLggI0DNlr8jAvAo5Zfl0ou1EFs80fy+j13EjGX5/Y2PdEyB41DLzkKL65a56OM
MP26adSOp0jNyks1b4VkT4ND9y7v6+hpjgPZaFDzBo/NNvAnlYPVF2AFtCjP8vwR
1a7/bxR4nFeaSd0eazD+e7Pel57QvQXMFaSZuJwPjrvmZ4WNMrnf66b1rYN7ngLt
2YgQZXKlgdhoDUOjN0ZhTlLn92JKT6+T93DMuLrEl4hMftTxDQTzmWGug4gView8
jJ7riujS4WHhCmNQlhVzSCY4f0kk8/8S5GABal/CNswTYapQEqNjSku1xADUkF0o
zzW6KLf8jFgEhVbaJIGMuA7tw3p/mrDMQHE49Kpifv2eHYCl1lvHCLHzL4nrq5dk
ZMJ6tfQOGtFtJxB/QrLa5XKGucjlUWNXKgRht3nr6RlOMaWVRGB2ar1W4A5AptyN
vGa6xRnsz43BXvQhOiIJ5oDMUwJZCy14MaKDr/oZ13o10M5COiAivR3GqAeMeyf7
/yoL5K0vNbBKhFAsJYsV81EDx7oWCFgVQH+HUqrJF1529CRU7K5j4hyz26dCspTd
sYOtfgvLVwe8pgIr92Pbfi0UiFzl2lOG0kQWCU1BTZMaOprKV/dWWDx6FVOGdJsg
9UDHeJWHhlnaXbUnVdGxLwjMyF2PAM5bD+sq6ZodypF4eDL0CHP+fzB8RnEjs/Ag
XbwVAAnZRikm0hYYo2BjiNVxD1Rveou+Kc1kFSdoaxyGfHRJX1snJgDBAXHQRlGm
GO2iUMXjV3Yr6lcdGXyGJD7AD8xoRUgHX51SPACe20fNI9l5ebKgnkMN9ca1WGed
+C9CQKEDDu+ImJ+IhPpsee1WnmkOpnCKMHNz31F80GCHPyLroiPWjVvPhSL3H38W
+07O5OdJOP1pgu4g2dAJie3V4BWX7sq1SwiRqLjDeL+8e5YZ8Mj+fJT6ysqyXewu
65VaZr2Qm3PAInRbRdGmrKUMu3U0X/cJlt7cLZoSLyBU2y0p2SlFwtF+s7XgOE3Q
o3uCHE/M8UwRXROhqpyg1wl21s9vM60E19p3SHw/f7dgOBHnV1Lebs558gVGYpss
5zfNMOcvsu7RoszuuJPB1RIc+WGK/YSfavqprtA9XMpN5aa+OVLMiU+92ltNwCds
Tulbrd5R8VxjsCTyFfG+KZh9dfdJ0fMV4CrX+VFEOCBGrhnpRFKzOlBHhvRw6bNq
cBMo34PS6nEMXHcdO5BjgQf8rdERHpQ8FZFGwllLBiPXZ9hXJwvA1TMcNGMJxjKm
U3Y5AQNuJKu4eKWFLNtSIzv2vXw5YgyhGZWV8yw20CVmPL1KxLwSz22SmIRtatJI
fp3cwvD8PFbRyvMMfAdFSdnOjmKjvFM9ZGp4IwGOFLLxQfqx9hoMnuShiA8IgIso
LIXvTzevkPcwCp1jKUF4QSaj1UqOv0tJ0DRy4mbA+gXOGzv2XBM367Q6CWOG3UfL
Fa/r5NFsYLEmlQn/m+hOcLiFx55eNNln7nT0SE45tPU+r7Nr+fBk8/yXXPmNnENG
P8hBwXBfSUmRGSYuEf+xQ8jq+SUu8mCTlc+GxD3Mr4h0UHTx0ZrP7gmXYwcKLaI3
Uh0hVOTJ/q4X7QwW8QJvFSoLg0mHkUorh4Urkze06iVURKocTTHcFplT9h6aJ6LD
AuvxnMd9cWoWUN02cGIS7NINtgllhHwNVXCrYw84xCE3gGBm9P/4bzC/2DFzj0p/
PWioNGGpjhvKxTEg2InmnQYASNLjEoOI9yytaH1nnjKSZEWzeaNr0v43KQks1B2l
ULJpAR/cWwXqD2S94Zzw9w7LsdFkmodDzJL2+0MbEg85xtmIvc7wjzO0WoJHjbyi
KDPC40lbIkM42+C2YYJBcyqRl0HU+8E2II+by92Z9+K1vdQM6yuhIef8FXUW6coH
WxbgZQ82L7oehu+tpiA2ctxy1gPvzwX8yidKngFavlQB+mC5lc1pPMGG36jVvwDZ
PbMpJgpfyk2+66b2xKT4/XaFmFDxQb6fcgPZ0QSKpkJ5DLDGABt1bLHGq5yBgboo
ejEHCwhEDVOmpv/+LCSdnV0dzUa8dU3VcfIRiJ6yp/ZLR5Ko0SeSt0mNU1g/P9zv
kweYaWZjWVVT/BjZfHXHdzpUQx4B6O5dMi+TqSkPXGlZnGE9XKDxRyPtoaGv7aKt
snW+08lTR0kDXbQNDGVFK3k4r/HLPZ366yPB+gVS4hpZVN78FSEcXc1Oj+RAzhnR
aEZtnLwmA72z+YUzNJXoU4Nop9oTc1vJB/C65zsaPii+iMFoEyAY8yi84e2dJMHE
lSbvwg/rn0/l9E109HMtv84gegzInxcUR76lrqkzZBOzP7s9S+XmRBNLN+RwBoFh
bV7JMQb/dGQYxWhaJabl2MfjURDA7u8RpJAxGWKK3y2i4Qt6qbL2wQv29zDZVmQG
8/qHrSGbpqynTEhty3244laSUC5lvF0VH9t1t/b5tnkI+5s4fEC0q0bpeOvBpZ63
bnskOCSR1FLRUh+E65jj1VHyGn5Osig81UghSO4Ul139L5zndbpFTKBw0LXbhP4g
q2FNyt6swxXyy0qOqWkultoVt0uUDQCKuY/7tK6MK2/baHmy2iq+vTv4fKbnoU74
jEJX6f5pH7K4KoAUEQDyi9G7s6/aSRz6RNwHX/M6G01ITZRKEwr+uzGs6vAEFUOz
0IttvcMMhSibdcIDmIHdXoPMsYTiENj6RDTDLtEGztxvY5OqNf5Uhio9oZEv0wTH
rh4+CI3Orf/kIeCykNiYxz+jDzjg16Iy+incxGC1tIuKogU8LisA/GtG7/KJG4Bg
r20kBqAtx94GCjc2BwbvG7w682xvGJ0XcUeIIFRA8etrorZTQASGUVfAIvrXyS0l
wHHTg4asFQ+lge9RYZrt8dLfp1TBTyt+B1iKAqSI9yJ0+FY17rzYOn208npZeTkV
eVT/A5wy6j+N/mkF99ZeQWLwqA/6BfSsHCHDfhIwMLjbZq1myz9aTdSCaq9bWngL
/4FWlCwbfWlvgE1/oxGkED7EMLNXeZgRoq8c9uQOxOYdUSqhuq2519vmv2uunwRX
H0jZWLty9XExNQD9+P8Z/UOec6Er/dgkWEsyjGLZIV70iwQ3kwDYe6OBsZgfYOAy
H5JtelDu0T4trBMcHXHtUpTFExbG3upp6xfxGvt2Z400Zg7jP4R6EEny4Ke/79YZ
hH9ePIXeuIdhweGvy6W2jTL/XDxuxHYXLiRkR8+LrUlGewHrpWnZ8ZEVG4L1Yewi
a5Zw75tbGNO2lsarAlzGko60hBOfDFVqaipJoivV1ts7jfNEMJ4H1jH8yW8lR+Oa
TBEmoFtHmylNQ1D3z5j+1PA+uaYb/OSUS+yNBGPSxKVfmZzB0p59Fzq8jP+d4xME
D9NHhh8MOFgjhP5EmIGQ2T8wRbAwWGXqsYVgovESMB03N5sSYP4wmpjUbgM0XC2o
AMw6FJ3WQtKpVL/x9Na1caVcHdsBxEbLh6BHg7urvIByk1SwCQNgYFSzRqufUoqj
6XrSH2hgztoMJU0q1PPqxs2a9iwFFLSrM1Jay1hkfKV6fAj4DCtd4P3ZLIDu19V5
ybP2EtrmpLTwyJI5LqNVGGXJAwQiAh+TrdxSK3jH0+5Rd2NkGrIycuznt/AuYNze
1aSucujrT9wY2y1cN/jJFy6N5DQXM3JLy5MXHqXWJHyiRTt2H89uRMyAh5Htu89w
M4zL+PoEMIPE9+MRoanFNp2V+jp3FcBDXRpOomiCx3tt/XalNonPkJVJFDsQZfYQ
xs7h57qjjhdpy6bIMzgBNHaTqBbnzwBAHXpA8olPf3FR/SEW8foSm7fj18qqkVya
n41Od/yDuRW0++2HWrGL/hd2fuUfda+ulRQ6ynlxAWEkVT0Ng3mb9efF5FDSphdJ
beqmTZTp4If3NVhKtm+r0MvVxb6LJmUDdSZQm5V/y1fO+Ah4/w4cONgUuRm6kzac
t8h4eg6JV7Zy1Rvp9vh6HrmiRThA3qcltCvy9GmwUJxaxpEdhKo/LpcHxsIM77pe
c9pY8nMXFWFgn3TZ0CVoOoFYNPpL1ke8T+KuJtiyR6x6GudfTbCswruXZKRi7IRH
3wJgaBZCIveV76Du5CmWQ8Vws6cnhLRQVHoaz1YlWjXNiPQtpwUtb4fLe161u1c0
yQmREap0OnNy6YNVxdv34g5Qzsthn3gBmqr/3KzQTUVqcX+dcXk66UfpAiJsn97m
dL6d7TcrDbPY10HwCPF5dNOwcpTyOGdSPyhdiDzQSfJPIHVVv/j6R/4VAp2l7TZI
57XRPbSkIqfRL7eV7CtO6Lrx/6Oj8iraalAjq21Igt+41ced/C2zIqnY2mkv1leF
3AA9KDNNilzjKiCJhiBfpoRw19fw/hWtweCbdkSaBpf98zrXuXHEc9PcEDf06kcS
i9BxFSW1LqC/UoylPJeQ6nHyCPqd10pDxCsg8QyfApXPzs4t9whMrlBFP2KdQHQl
Gz/JxJKvgNBjNsg+TcM4xaDDh83jYrQl6BJnxKqeDyFDjq7F+evXphWQ8x/lyMyD
1pTpkBelqnns/jJW2wu263rHfIc+MCIC+089VApiAmZ8zsBec797dDwul+rc7aFa
75rvd08yjT6omvDKWKhwKroeD+diQRejSMf+0SMn50xE2nS6NEBAl+WfoQwPcUc1
LBoakr8kksFjHfWsUEjG5q3ewlpSEU3qmLHMOmnsXUDtYv2uNoLipZ0kzd1m8dFR
ExMTovSqUAc01wQYqg+6xsfTM+W5S8ZlhWVzEVRmIB3mnjPo56tBfFKqwWDHmyP2
tn6fV7VyMoJv6LR22mLKtbYsgU4PXY+M5eUuJNvAY0fOgl/xH+eKgODlDzrS1kp7
wNrgSq/zj5CeQMwnVkfCIuR7uZTQTKv/Mhu06kjqMqd7ZEgbpoISIRtf5+sSOB5b
X30g8WIu+jCiZyAKBjipItg9nEI7ovnjYFHVo8gZT5ids9KWWqy/ii3gInhd+Myt
v1InTaubYdi5mrylQIwI5YE5qE8X9wPABA4BS3DRUttukppbyLVr5i5f/uySinoF
gbyrexdO0IUf/9z+tKTSm6m73G4Z1/r8hkNuLARZ83ixuS20B3LaefsjT0w0Mc86
drQkLQC9OZk5L1U3eIXGgrn60BhWKCfpd2CT9UoK5LE5bWlF3j5cIzauy6Cr2CvO
Bi4L+4fFqz1obRDF1b3Gx359xYuU2OShs5qI4Ty5ozWUN3i3oH13Gned0gGoy9Sv
FsmPVJIZVQIphXG3CCngDY8zre8QIPxq6/Y5r+ud+jQ/Wbai3O63xn++egOTKqcp
SxIZh7U4NmTtfT78k7ZggI++siQgakyeahk6f7EjLp0ZHhB9Geu4B6Eq+dR8rheO
VEhVlq6NR4M9huG5ex8MOHEtrUUj3y5XhvbRYVifnNT89q5dqs97Lq6pfINYsYHZ
IydjHvGNUHqTk8u6z0pbOmSUP754JMbvJ5iFvtbEHJTgyFYNKS7t00WkmymDp5aW
xnX4PyJtO5Dcuhlza/ApgyaWAXdCMJnTcjRTg+9qsUuBoiE9hTCdF0qkTCyMrAQE
4cuX8RMulZhFYK3J9hpUovwLvF66vXMYWLWKBNL1uzHDJf4vtVw/DR+mVZFu+Qqj
s78vdjwNVpoMLNNDuzgjjq10RW6IjeqENBzM8DUF7Jw6Cy6OAYZYdiZ2/3Cc/w1w
VrHrlxgPFcB3UYgrMwAcCswlMaDbceftxPd/zSEDtpt2D8n0+xHdiRUtM7/ZIGSE
+u3v2+v66HyS4p5L7vdG2AFj9P34C8yHRLdoD3GLY4Xf6Q95OGckVd7SCJkvOC9B
hRgHkY2L+qYkVM1CjJtDJszFZHVj9Iz8U92iF31QtHmihZUZe6QTMbe2dLlvidOD
gi6rdbVgJ/wLWdM7ySPn1qr+IkAqBn++dGpKu2vMf/h5p20N15XR1GJlqUHrmwwl
BiAAej4WahSdeM/Bx6loxyP6WLakmX3h3dU5cYhPvzLdOiBvPUd/QATAzI1Kkpot
xWbCmaKy5gQqqnmQQKfBsLQqQv5q9dII/h99ixXKhn9SKde1MOjyX/YBo8WKCmEQ
8Rpu8rPn2AwCDkVMOh/aZVgqVj+lHQmRvwhE2Uiyn3TVu/QOiMyR6tOJN2644fgv
ANmPlbpdjyb7XoaLTCPWvX1IiJgKfiTndZDSWMaLyrIPLzTQYa7Dv9iRcFQcuhvI
GaGDPR1+PyXTRW5mqxgPJuZAHocEQKx7ON2Gxsu/lmBNsrbQo7UnvhHUjmihlKuJ
9l3qrrBZJaGuqwT7ycZMLLbMtrfdO8gA3u768rq+4/jQvjhFAE4pmCXuUSczuC9J
Qr6BQT5wRsY7EVSx4Gw6543/bK3CJf1yO9okLBottniSxkPaQW712KH7yj9Nv9nw
GRDjDKqj932T/NOa6/axVAsoDKjFHzhf9S13u8DJ2WC9EeWic0s60pXJt8unJ5wQ
CZ8DXQ5XqkmedFThbOlKri7FGbXEmf2P8UqP8ucchqSC4Bjl1DbPkyynY9kbhPzL
zdpkDFwDBI8kyxQU4Dc6TdM6JJC2yQBjOFs/swgEAUvvt/cO81Rl6pBXqvCYLOke
90B9Vs4WQEdxLlaDv7ry1lFJ8+5ZA/AoRB2u+rKap2by2RpmeF/pTBT0fggfewhj
Xb4O3DhCekQ7oMAKSRDHf/nR5Fgm0P8UqG8OeBblBUNfCeJEqf9sh1xJkZBPWpkm
q5A1hJUIIpebI4XcxVKxZt5nQtDoAkXryCcd2+FCw168esPKsLEBRnT12XlL5SRs
fWxqN5ItPamlEDltY5IF2KusfDVpdGosdNMFbJYvDtXOEkMoncwZnhDCpeGeZFdr
VA5A2wSPdSIBJrGcmiY4J8FoHlBoB6LQ4DMOVrFVNsrTfwYuFBVaFcC7WOVCSWO7
KZ732a3w+NOY7eKB6Zkm6VUgTLnJklZxR+Kv53fbzqLRn19ZBiCYM/gU4Yc3Yk2m
YC7/wrPS8cfwgJbQoXe2Qcvb4XbGunDo8v5FszvphNg9BNmPdaIt5dhE29lo7mLA
/8+RWYIbmhUxl9yBgnS9ZxZSDsCfC9OiO6lSryt0tKgDAyXQAKugc4vXElW9Rc+B
hE7x7e/KKwQrzZoUXQzrRbcFq5rOT8gEAeXo2XJh7B+iBDMyJNFmkC8PaiUBLIix
oDSzcbnJs5onx2MZnuk6cgLU3cEsf7+mu3L2X15G2S1Ik3MWf1i0HOW1eqJzRLaH
L/o6gOA+xXhnkLGupyNH2Dl+CTsLd5fGolas/wPV+5whSH5UskTN9bjBNzOK+PXf
HmdOrN4qptgJyoucpIdmIG+a2lYlh3NviPYCnU0Fzv7tXznvH8fYwlwBoIDlP9oa
i0n0mRATkUrKMM11KHHRk1h458BIQr77Gy4RL5wbQAsusKbplE+MHl5+MxvSoMoL
fZbPR5N2h+fi+RVpu81MBpFJ/Iootee+n+lhqSrZXpAxlXp+gAUaE95TZgoVXNZh
LD/PC1XkF+5NjfAxM5VMigqeU4mKuIDgVsYtune48uLp4LbwwlfHfzfoE+xiqu0f
KVqyGaqEdF3ua4+oR4v84C6Gq6+LK6B3x13lm4NyqptqLV2yqWuY4I1i5chwycde
VKHSxyz8CO5wMTtgAC9O+WTPnL+vkfxxFMLkezxLUx2p3G5mXy8C4J3mkR8bWcm0
8ck9eGsWcFAcat+4VRjRzO705/LjHQ07Qf0J/qm0mIiWOZO0v8QfbNDMIb5X3TBg
i1pU69+QF5OYzp8fQ+4KeXWF4oJVfcKWSTLT6H49dLqkO5j36UmN5ce0PDyYyd6o
oS1VfbF21XtaWJigCfvTO2Mx5T/400b5aLafDGvdz2/IFHp6CklxuC4kslTRcK/X
e/lIDLVH8F7vryiF8bgViZv5v/dORfYZ0PBVIAtRDoPdvfcAbPj/PsuQLjLd7u+S
gdwq9+rA3R2kYB5ukfdnbcUw0o0Uar77zI/EZ60ssZu6Fnv+YEwvK65lgnxhEXL1
LMa3iHioqFmk3cNQ2PFH+W1C7HE3UkArjlWJMuaUIM2yFHaZ9rJUtc3vQ+tjumHd
6Yej2wQHP8+hldk9Qd0sthipX34I4iO3OK8gSqNlGDCYBhNPaycwm+hHX4YBuvMh
KicA5ohmZq8W9zn7iaOQV/0trG9/VssM+HhzfV4xsZ+xYwgp4MEgCrPJBp41a0KD
CKLyuRoj2p1ypT1M2aYGCvGscgXkmv4xN0qw7MBOFmT1Z7ApIJLEZUElDBzS5fv2
dfTvwPKqGXQJTOkPgHs3v7ArCPl4/znzYHL2W2Z020BKyOFHDSY4n6q4j9HwzC4P
cu/uDpgZvAVOo3YVNmKpG+pz8ge9j+4ci4A7ddig5iYLZ2f49FsjjTi7gUrlF6C2
OA1AHhIl6UTYWvxMmmuVSMDynYOBaDmqZIXYQkCBGXuH278UZ1xa13WWhJYonG2F
u8XZEvl6S++8IASkNl1LQsmU/qApvwui8hbswrDxNoOAn6QUAj7x+b+s5eyT6Zan
tEhcMcLWY1ADL2y6KeWZaesSr0c9KEkL5JC3c02PQYoVKHfvB4isuczq3YxXGriG
gzoN9zJIkIypkfSiZ/YM4YVseJOK6AJovQDzoPuk/TzJs5v/7KdfmEy5O0ByiaC8
lN8Y0ZDBPDH9uLTSPcXPXdbeqs0G7ceylO5FI16pE0jUl92dZOOim+24uRk3VBMB
bqHsB6hgKVPcOGOx7c9uQWL1DwVOBaNLt125hzUvZ0Nju7Uu+Sh/7dE6vJYaDXWB
nWnNfp3ZY5Z5ARrht61HgBv4lB9AOBlfprUcAvQh+0y4s72ZR1l6FkasXi+FXvDj
SqgDtUX/VdUIohopZRT5qgLYQQQTWfZ95pJn7EPuYeC0UjHYVOYS8qVyQBI6VfXb
OI5xp2I7/nIdUmY3fOW7KPgzqCQI2mMgEL93Na30YckeZ496l3lf9uVE1zJQNDQd
2lgcE+Bq+HWkqk6h2R8RYr6Rq8SBzTUtL2Jhhlaow0Kk/NAEiepQN0D0xw/GOD4u
BurVd0MemmGB3lO6kOslNJTzr8fYGNmiMKJyU0rtgx4KQ7aXApXLBEAuOLQmr1J9
bDnVDBxgipqsspT5XcYo2cehJtg4Stba+YQRWmmj2T26ZADTb6WF1Lz5Io/SFDQn
OReNJIA4fFVEccTQErPINbSDkH6rWD1sScL650/TRb+IWKqfaCvmspeL6UmT6y2R
MgOicoJuUTc0SDYNdeyllPyS9ZE1X6TpCMldz8ACzgqZeYYMEjgQkGgM1tLZwYnF
a6sbD+oP+YR8h9XEnhec2dtNe95/e9zEk11uLYvee/9XGZ7e8LihK2O+pG3/Qrei
mzQkFB4psRF4WEr/o8/HY5tYhOvNEYqtDIppM+24MaxW/te6pEXaq3/wOSHXEBzA
BL3wsVwvFdr3VU2870T0Olwo7EFX1wCaIQJv1vcqDziA5hapgZ6H6J1f+8phXltD
l8D2pL2CbhuXXheUbVZqQK1LJm/tfcNDz8QEpDVMF75Iy6fFgXFYr4y9NWCRowz/
zPeOCCkj5KWg31eQ4TGfRdjbe05JRVwWdrTXuS52tGFG43ABrfzl+CpNL1DcSPth
uI0rrm9A/6gJVG+pT+o4AWZCHAdumZGx/AHHO00weBlzPDpJN+IS3+xQHd4bphl0
p5FXA1cbmPwpeli/NnLIRlMzt/GKcJTMe5kAlj4SbJO7/rhqxIRM4NSE6e22o8Yw
4hpdDuDkBE9sqBhj76ZIANmIJ6/gtb+bfDNt0ZhKbugKXvWsyt7UgIimIUrgs32I
GCgHS1+kvf8eDF+4IwbFPif5oks0LkxXKT4gS6r8A9vLPRfWoidgWwd9AsOwSTfT
G4+N9JAX3SIL06Z9rPPXKKxuhsK1cXfS3YbH3MfRrzAXRKcTXVmGtbL/Vv7loQw/
GEiUqUMvsIROUwsPFgb3/QFwLSj0pf9Z/EjbawahUbLsHpVHEn7TiYt472wgGF9w
Ms32YJC/FNpYj7bPtFh4u1DW4WjP8f1BBMY3H+7N7g79aGcj9+UIa9WLLUvevU4S
lucnDzjcwP6EgJoPqXXrvmFrRNlFkLkIKKV62ixnjteFc6DNevbLZS2Fw3geR3Bt
CsRsaMlZiWC27OTdDz+ZzLbtQmr4bB8DrFcSZXHzBtaYNay8K7OUOoIObcMjQ4Rm
rTiuoC3G4lZqqS78bCixKdBpw59jJijJtjCZoZGNLSxTfEO8TMJZJJU5rJbCPZze
zIfSNqaiA+8S/q9/+42Nfivt4xNLqT1bTfdPUShyjm9BZbo3mNb6Dc77x8eWY9lq
EfnDdE6JD1fdiwE0ESLwCEAMZwGD/9uUw/OHve9MP0Pr5n4r2g1gWhIvRj8CFGhp
X/WYcucfBXGVmHhsQxJ4LrhLz/+DUT9KX2PWcDkOStcY3iHbSn3qC1z3CD5xMKyS
MN3ervtmJOl+II5aSrIupWQDj2MKuIc6QKcW8ZWqg57qbRH2vVROZfe5H3RK8eln
Zxhx21pn6kLhD74tNEy58jHAddelbu1+uTYvUBH5imNrQB8Mk8a1R/qUE9P9RR0B
/gX29FY55BANspzOSt/OBtQfOVNosmhbQy/taHFup+laVQJL7eDY4hTEnPl4cAnz
TS6nIvHPx6Tq9rTRXzhJPXNHWQCvJeJUPx5rrcWuM/09Jy43yNf43efFmtZPNQsP
1qVNt5sJ7lAvxVkFHveqSyKn3Ppt7i4lQ+5j2wJemAxDMxSBLsR4s1SbOVm9z1ko
dz2VeJqXAgXHTd1Hr92SkV511zM85z0PPm7LjzwfEnvGTinkpfZ532Xa5KiqLsNH
EXZbQLOtjwC//DwX4bVXNjhKtuUsWnpkmqO0L6u8o/pYTlfZOhFY/QZq1D0JToul
PWGqkGFldmGqqXzuwzkFidUKwHjA2ks3Lqzsf3lGd1jXxvf1ZfgdDXDYR353B4C0
LK72zAORJSctlQNRhmzEzEcfGUv/IrJDZnDJKHk5m26yxBoLgQpXp1dnoOPME0Tz
gUgk9GHAMxSK/q0QZm+cldHQILMYLuNl1m/hn6jby67TY7JX4D7w4qZDYNjiDadW
qipy/mCsiHJf2/ExDelby2jGTALkK7vE020ZVTf1h16cp2AnDqAk2yfNxggVPvDc
LbAEoNPNzcwcgIkHhcVwv4lUdsO1TgZ76szo0jluio7ZQUflOO/UhzdB1vAB9JBd
sgtIruOqWKqW+ndAaN6gYTDgNIY/4TdVuEFCVk5SbrccmVH4WIth7fbf1F2rBRub
3jJO06nMEJfiL92t3rbEfKNMuQA1ifuYHObgK0UUD9YvZFsehGvRZB2e8QbmfY1a
ZbGLLU51J1IChaRXGbD11v00+XCNwDOYj+7dAW4f2joOtYl1M7u8ES5+Gysr2H8w
eZhwbRpM6OkJeihH5mW9JhuhHUcofrNAnKZMzEvEG7rNP8i6f+ybZgOU9mw2oLIW
Wia/8U8DqjavLe32V7FLMbqEZEDmkwVFl8CXDlcRp2VKTAh9FDCw2GzdvihSAu/G
K4GTSS4Q0yUAJV3Zk0Wih33CPvX2MYwGv6zNzNVMxl9tVNQBY7RCUsTZOd1af7f4
8zYelHpH/fS/wDfbQDIjzwhreZU9YBB3XI29k3SEhIw21e99a8CEzjQsyR5qRg3b
3PS5LgaQmsMQPJeaPdMjzrsghBcoonkGLJT62xPhkQNJI6xUTWK30m0UxxswQnN1
Ei9M4iciksCOU6XptlZu5glWdnbdaZISr7EGcc+ahpqHQX0BwhIpVO7h+rwgZGsB
KYxbkh3yvyKMWaL/IL76FgcHjpphfyx6QbiZy816jBb3/xOPSPbHCycVgWHr3ng1
A51OFreWy0g6hTX9fVDbLBJtMwW5/hMot7ahjqvTQAWqy6hCGaVdMFnZSzwJjlqX
r52+q5c0l9wOr34s4V1g5gbLpzcYBmxG72gTP159mPYMp4/ldLU5CqvYYTfwF5XY
e7ct7osUY/h5EoO//m7Kehe7EnsB1KxdFN5noBWsXyyIuK3tdY6MDd4OGAHgrmve
zsirDsfZHy8npKrqnaYcPlUdi+o0u5XnKpOOyf7xoVQxp6nIUeWRzHsU/XJH+uF9
PmjMA+a/nZ7SX9QJDUXNCMS3ZmfBVZHxJQzwztFb+Q6MaOBSudumAeV+53b+VGrE
phcVfvq1ToFwi8zLvMVwyI5ZTxaoRQ417yZppSOsuTl/IJG5ACNWW3fBdzDbfn3l
PBRDrG/WJc6eaoE0IG8Q2ciEvPcy09bRaQQhXLirnIETCswKZAqa10lgb2ZsgkZo
1tyzADVXvu/ZzZGLhSrsY6+AKKilKyJ8SKNfhPcr5U4/tR40Nol0d/CMaSmgIsti
uHI0P2LwOCEjTmxaF+m8j5Jh+80UKjhwYG5zBkKpUNACnc6nEyh3LbmCrLKogwp/
J6GEj1HnrNrQUyTgMWXo5hI7uf+mun65howCKretQjcWlIA4A+biQKp8XWIRZ26t
V+HXuGUxXpe/fkTy73Ew40xRKghMOuH/Fy1Edtu346EVJFDlJ/Z89uM/F6lfvRQJ
7R2wdNK0FdsgzWkXa+XeHSkrNG0HqZf12ThIZ9DlUNGIqKzlWSzjMNtX8yI0E6Ig
ywXewUcf+TIOlh75V0gBINirbrc+WNljlb8eLPTGEJvULUGi2OTCtibpbrk6OUTB
RQ4kwafjScyOI7pbKIDZLrev4hA68pXN1m5NwkDVXHWtmObGMHdq9F+VfVx6M7yE
JONm4z2DQOTxU9Y1niWSBvJ36oXUXy4vrhSUQyXVbSFZWDopJc1cWPi5xBsDhvP9
9lm0R0g3H8xdUnEQyNB29cmfRN3nf9bbbUU84g25auWJ1f8lXrTtZ18ij9e2SzT1
ai1HyljMKklhHcLwysFxug0m2+UzktqZOzvk84mxP7zPC+xuNPnLc64vuHLA0vaL
D2+L9HiB6vTrNxA0lKAlRNLMzg45IXYz83KVebq5vORgN1fNuQ2g1B9yZl8WhAdh
GuUcajez5hL56gwSl6WpqOpYQKmnKB6Za/xcjyYU3cB2QB5/9LFvHi7pCoWtQnbr
zbBNYiEyJzTj5/zRnhlREjQhboO/zpelvQgYmmPfSILsgPiESxRyLkV6/EWm0/8d
KiansuTUYHmPvSjokT8RMZOrnYS+w72Xr6ZrgYQvLefcadl3XydvMvw/TMqIzPV0
S7OEBA5TAcTE4ar43O5n+prNdvpDDq8f737OLt3zLraa2E17jMmbP+dZTbsRSmgP
mXWmOUON4a0k4x12iMlZTyASAFSXE7C2i8UWFqlgOiD+xIEKWCTp4EzkIte3qYw5
NSRe6DX6AsSd8WiD9bP3JRsdRjpiSNy7tIy3XT9WOYqxxpvGxhKShLy8KTf6a07R
h8AaiTxK6aog9HpaF6cjf/SIA/RGnociOq6AaBMSnWItT6DBq8CQ07dS2VDHqRgy
zDwMrfd8l+trgLYlbvWEcFbzSkNRGwPgXx57qZZK1sxVOOJx4LTQ3vK/8U13Puzk
Zgm+PDUGft70ncMHkwDHDJd+XULmFUw6Ac/WUhp/HesmHI7aTEKZsPJkwLP/AwW9
skc1PpzM7OHFVXdmjezTHLw4iDtmLHQLlEEroOVszWA7s0wXitwzASKGQ10hS7Zc
DRm9l3pTsQ4uHCCcqnMJ4FQATE3Lzpge2wcwUV/jdg0wXxU5I16ZbqXw1tRuO4U0
St1ysN6VY183lRX+6aQ5DJH+hE7mXQXT9yBt8gqyDXjSN7Surwr7VtlP44G9rpuv
in8Bzu16FVARh+NyvWPqqnW3xNXXkGi/VE2jxd9LjuqaFpknPJtLREbS3TYHiqOU
mY2KhTsm6B/hhOVSMqKA4xK1PJ+DbqtnYtCu8XCzm/xGGxhV9aWYCWs6J/cDyq3T
qBFqDym8ylVD6gHL73nZywFANWhmXwA39a1ekNoAZ3LZmihcUawTV7TRORfOxNyH
8ZjMMyjBpvp4xpjHCiTaYtQcmEr59Ne/0H4t8e4kUidxpmlvATACDaYmiuNZZS4b
bsKxjUs18AO9JPpkMhLbO10NuCu2ujKnqyVhcEtfrTtTz9DzydPIeCIr5H3Ryn6N
4eDEZthLpAZ5UHoLZPB4u5GwaG/WRQZ+MdnJPhKOjXVyezrOqssK8ZVaOhl+ofr3
3MW2fstmTdkx6B1pYOL4Aiy311lR8hIViF7nA8y5wrXeb9FAxNVb6i9emOckaP0i
Ff2wY5r7qUo8bYHCZz0P+BH2k/DyKgU4aidE32CBmMLd8gasrLV6cwRR37RHrEMM
GA1G7lWnSkgomUanWrswJNwRwDTbMQCfcR3tpVMqqJmIqevQaP3spFfb785wTYdn
76tH1XA21yD84aA7F0sZD4aRloFW/RerycnxtcdYZmTsZ07x2k0AiFHL5VGLtzXA
o/zT/4+KDwk3oJPTdPuBJMHYHGRoQUmUyPMUgoFnFaDskJm2vcYMbWWXTPgbwhKz
CAFN2tPnr3+QrhMOKLsFQQDmq8b4drGEdMCbqarEmtXePoju/dz+vwWJgNYLAEzE
rbZnLVfAY1gEuAn5wxOygo7qOaAwmw9GBkqmWv7pnMrKGnFm75mW7LtXN7B/b5KI
S+sd0vm7To9f919dZJv8fD48r1uK7usDjXSSthbAr7Oy7/IBOXBVWrCdplLpEySL
U06N/hN/GWRhuK7/NNwr2WnvrttY3PoRN3Io3zHjg9kyhyv3n4GCrtgtCg1dXP/N
kaGrZ7+I/bcrUCWlZ39np5w4AJXIGpNC/BOyu5dpjAzmJJ1t/smifB40s7UM5T2c
dSBCDi/UBR16DlFEizU4mZmwr4PCFWkclPeXsq1yLBDgT3PLB/Y70JEyJcdtitr9
9PBHibtFwAYuPbUYQRqhTCjSMt/WPIWMq10sLER8BtBF0vUCHLd3vF5UvkPT+zu7
WuST2KMQpXHagwo05VtUUJGAejMQZzXB09rbwugJZD864Oi3K4FcVHEoJi0LGg2q
UlBjn6lCHLs1bK9q3DbogvcWfar0IXSZdyXbf2RI81z4rusxxrbTWztgoy6St+3c
r1N9uOB7dNvbwqQtZbjNOfKpliUdFcOBNa0sgF0vHmA9lC4dsiNxAq8NrcyqZHg4
Xm75QBsZerW+357hZX2bDGtDd1/wOpCiofWjGFMPoUkMICxsRTPWm/vifgB0B6eK
pCDt5y0n6t7HOzwDzyEeQvedW+SxApfWVQSd8hPuf4PMZXEb3KJqPE6fFoXRyojX
TgHoxCjiide4Nf+uKmp9fQGd8dbcDy1EL8ZiP/D0JUBuTXYhQOBj1DqOoU35oMoM
wYwwNpmwPkYYDGYpcDWuNrlr2VK2gViX5e+Jm35GD6Ack9/BhSmOvToVwmJ8k+n0
u0iulpZf29mSRc5UqPdABlYJ2hD2TPZFDhvM/LyvjjJ0vCR6C9gA1lyxxCaBW+2A
hhlweiaGW0WtDvTReQkr6w1m9157lMM6xULqAkegdFyD+oCWWCjj0VnS0koxRwZo
/l0A3rOkRMt/FvA3M8zZOt9880GhfV+QdZPt8RacrfGgFUt2IBCzUpt7pWqx5SI9
EFjddOhPRb1Qdnn2W5Og6iwoHxA6mCdLXey3ShOpcWwQyxuWJuz4WEAMGqr7mFkd
OVajBoNkxdM/yT0312LeBjOGGHpIH4ui+1TYrzklXhwXtSiCB3fpvI1OoLK/WPWS
af0ATIdBksrM7qu9Kajg/a0sSHnlZFXiZO/wE1TQueCzln2nUykC9RgPFuaIYAc9
9gBuEDQP55aCrbgTjynWZJx/t56GrIUuuXrFWj8LaxuRH/gUJ5di2jorGkixW0X9
uZfFTJkAN0DKRsj1nA3ZrMOxvEdIm+XDigZ6hO5vQk+uNlW4T6IfP+sxU9lSYlEo
nK138G/P8FG2abBUFCOCfh5+C/PbUAj2vVj1jzq4cgjhrbrjD1MQge+UGgHDbKXo
4Lbw0JkMkBVmaN/YpUETX9BXxVaGQnMOktb0PyCsHMOsHAUr43gOBht53LVQLwoQ
GY08PxVEMhfxWBuIyOFQUlzkLwKDwzaccNdZ3r2ZIpXCZtV5z4QaR06tZ1e/QAf9
VrSOoJAmHWUgCpmvz/NtAuTRn/RdbuMRZdMxRNCp1FSLKQpvo66RRSj1TlBsZGeN
iMj38RUip5cT1S6MsX8qQAkVoTPubeBne7tjMOp55MLtCDpwQkRZcIyu9CqPSHt3
X3VFCaIdUQoS4LPN38ZCnFFqC5ZbHAbSNOOCgKwlXRLevrC5v1lxrKi23Lc3BcEl
KRsPoOihfTzP+WaYaUtXkM8huigfyI/+CzyWQw6p/93oUBfBCBAhCJ8uNR+qJvYF
GFehWLsLzbiakyZT2IX15fgigeLxWGHFC1beb3wbp/9Tfx7+U8G9JA53QGx34JM/
HctNAIU1/fHCbIHinAjalc+7gxD4nShLSKj+E6fq4TDITXwMTDbfKbahEiefZJhP
iW+tW7zLBu026Cgt8rhlwKJxqi3kzrLWlsA9B/7RZjYWqe+FMuHSMJhOFov+EH0W
92BYdq5Si26dFewzS3oPxXZXWzN2g3LEuI+gK5g9VxtGSPkm5yqDp81ZXuw4eyvA
GG9i092WtTmwMAeRpslZo8tdDfHfEwCoU/2duFNAwJ2XwSfl/69wKJ6e2QA1E7ZJ
Dswl6+nK+gj9r8uDY30U8dFcOk6+EJpj1549Rk3aXgQR+b9ERxLhCt1Bvcqm/ZWQ
G8SLCZgo4GkM5CPjdnB9jGZ624yLv8AqSuuiK9oRTldChPXAdeKQhklgbfqfN4hy
tP4fYlm6s0j4MhKniey9olcp+kseU4b/3wTgQ4xYwZKmpuNzhW7xii0061WZigz8
SThCiL1re0cyEFX0c3VW4Xl+1ov1iR+untClG7oY7pHp4K27qmuxxrXyUHayVcES
Y9GR7lr7KGd8Jh4CsQ+rABmzY/Ej1mjNO9yoJqA2Zmpyx1PtVt82/JWtglsCwEfP
88GxENWXKUsppSKEZG5z4o9y6TmVmrz6jOKpz0vrDEMiVHqY3QZUnnWOpE/bTEJZ
5SCRQrsl4L0FeLQstIzYWTWTxnHmfIlASpyGU/ZTUkdE7CI4jH8DpPEszEo+IWwR
wnpNMYQzk8Pusaxth0FAGJBin9JsIzXFqZwoLmezoq5WzHkDxUHVOyUYOXWF5dmm
flA7wnKoOP1flNiOpxAb/wBczWdG5PdRcPhrXc1RR6J2z4MCKAnnqSvZFE9vck/h
/BkoGIUSaYPUSdVHJJcY2TXB592N+5MMS5B0SbVbnAZifIWifY/NmcaYJ0A9HqA7
Mg7LRao/smnt/gGc5tJgwcwR/Nnnp7tjQqZhB28Ewn4gyx1CV4qzPzu7XbwUJpBO
Q4MyLyI//x+5ftWIUSN1ZBuacvvQXHSL6NQtbNP6o0jHR79H1eUjMvFSpZYfTobh
q5e0LgyJa0gV5RnpsYZN82Y5ipxhlXLJnnv3Xq7EzSas/PeVIRV+xyf8YTlThqAC
6EREExRG4wdCNiRmXdlm3jHfvygci1NjTpc3SFgrbc4XOM6eT04WwkxazAFN5rBh
Xt7LlqLsvimkHBUvydefYLP14C+auOosgzzPz+H0Swk63FuLgt6L93pjNRkgSGfD
F27ZQRX0micfhiBteTWCVsyNkTApZcTbxIMgIRyoflq9LNaS7F13NKJLwA5YMYwC
e4oe49n/6Lf1NpGanZRsK+/LPZQ/L7OqjLj3TXyKrX7wZaCPayMbBEo4vx2gmowx
fHucvabYsDiuY4329FZqtCWaeAQtfcFllDaVLgceqPRwLBNDbbW+HwOvkuIvc3Oz
BrwrVoP6ln5gL57KYD3gLdS07SEEwZBHTO4RqIz4Wv87QGIaevQ8Tv5+GP4yX/9+
ro+qCuDaPUpdmnYn/xFW0c5WvfWtZwUh2ykeBy9HipuJvoGJrt3npCHPDtqw8rcx
Bcrxjlul5V4wiW58kwVkmv99lsio13mMzpk9HTjKTm7IUuH+27cq8fMj2oskmbeH
Z6v4AvirKePiVp7fOHfCNx/CE/K5rOrRygwFH+sgZTRc/vfZa2PC/IAHuUvHTtAO
6p6zfSKaKXjMN6eFS4hk7WzxvBLDAD99HTjAL6YGQ0vGtN0Qf61RVe1n4A3PPebH
HNSQwlHD5xpkho7qlQd9axJaWSSTOtO4iduzqthrOg6jz3dH1wXGJzF7FeQ9eoka
j3F5JFnF6aPiVxnXhxOoEqW949dni1ag4Rc5LbiyplaxS/vcDhXL8Llcx6dzGofT
httJgCgGvOraxd+da6j0s8Aj6Zt6L6pP/UQDr2cUPiyq7p/LVxMYXAbDznzThP4l
teS2+Fj8KVrqqtfUsD7xxrd5k9WpjlgqoJ4Snq9JjfoDHkdZVqn2Eh/HA29Wbak1
pixJ8vrphL8eKg9nmRxp5X6AzSc7ynUqITHiAsNzH+RgcFGkkZ2k2JZu3C9/ICyC
imWlPmUm+l8X6Gm7Jcp3JH1eh1zrsENyMcYAgb260ke9NsQlkK8vyOhlQnuUn3VT
bA/LKBrF6FnLm0Fs3YpLKBG91Wth+TrXxds5+pwwZ1HfeSBZHFVbmmFjJdXGmEgW
aOW22Wixl7HM7qhFnrTsz+rc8cyUr1NBqNKKh3VC2TkMJRh5o5+R+WkfDMEc6Jxc
ECe+cktS0aP3kRLGVFo5EEtFVuPjoDxSWcIcWC5WJO2cjBcGetfyyHs5ldUT7L6g
KVzkMB86GXymIIG1sREjxLEliQEN/FEYdqTdYiTWz1q6BqGilliGua+5ec9lN/9a
u6E02rnXTWdIAR+AWK8RscsWJb6O1ke+VrA+kB1aEz9uty64MAp7nU99nUXrzcrP
gjU1CMCWXB8pJ8rDAoeuOaIJTSm9L0QduByCoeCy1Bst1H1ReaDt0JKu+rRajkD3
zJXBqiwtYNw+4NbFJNVYfuYQKFqhPmkxQXJxbAFOSqdfO5j0fp8lNH/xVIN0k6VN
O8LdWd1AQfgANNnsCz0YL/pxuAZ+0LLDv+gkGkXGf2dmFfLZ8SpHLwaNV4J5d3q9
tKoCEQ/jIB3itjucfbTtkPz8hNkp7dER4o+eyWvWDHhO6FOa1b884ldMhwvgs6Pk
xBDion3mvrWLN5ysLuIQbwjgaBe1N4q5ZA5VqO9MfjAsjoo2IT2jmLOmOyT/46FQ
6xPZpJCzsUmg/+7rS1mN5hPx1/Q2TF+lSj9W1CKSI39MCIcM3m53oZQ8gUV0buEy
RAv6pTNYmn/Hvhncpsud5WJSiGYfzXkrAgbUC5J+F0kXJA7FdTQahCMDAXXxSiDm
Le516kijs8VEDNgE6jWzrE2spBkkjPllg+NfmPL0HJMPtNjM9tZW2FE2+L2gdPqt
n2FW7aNmVmPPbxj8xgPr1lsu2wZ1WB4hwSg0y0woM7ILd0E4HL5DnhyqmDvrxKB7
galUYEgI2r+CE/uydMSwdu2hfd3kV4XRKMm5tRY82C3zsVuUI5rLz8e+wnfKyJaw
JnV/gth0X1yPlNfL5mRYsNaNyk1mnhwlTxPriH8kXGTaIt2hXpKqIZ0/z3FwIQ80
FwelE8yfXSpn2zzcnCsN+ecxDXFIgc4aP/iF94AQesVzZp3iHtMQHdJs1uGXs9vY
kgvuxznw9zd8yTt2wBPavgBByyjOR28i7l6XtB1QW+BIq7k+SPlKXUs0qDr0UEjU
AtyyKt1GtGfcMejW7afsfF3KufV5mw0oGZPvyOwJdZDwtTPRu6GHz2TZ87TFVqPj
eN79AXL4Qq92emK3CEQdrpOPa8Uj8KGFhCOs7Z8DyMjOM4fJHU+o6yq5rOR5EgLQ
vy3auDbLIU1pcSpnJmoI1TeDmHPS/Dc+Ff1l8B+DhEjt34uBEeNehFjNTDtE5LQC
taT21f8kLLKhCB3Hb4K9umrVk2IxgiZGwWFIiU/zCSqfHQu/fwHTaMIAbiPMJm54
+kOx+nFVoXEy8+qwmk7MJCY/qqqzTZhQ+4Zuyvcm/8PTI7IjjDwjEpfj3b77a+h6
4p8QD8ZvvZz3EpbspbHWKatuuCY/U88WQzutJVfc8JzQL663W/Fzx1ady0vgPFxt
od5cz+OmqvWGvkNkcfJ4R15JDAA4uCxT21xqgQGmKKV+lMgApRADV/+igvGu5mwA
gkHxkvvl8GFT5R56RZcs+0O/m75woEZG3DCVGawWeRfbhdy+mX389Gx+SVA+NDtp
FQh6GAXLwm58qrXgm7Cgu/FLstI4spotLnKP65Vb6k9BapYEd7Q+WwxjkkvD2712
BMkwYHIjI3IibjN2lPIIm2k8bEnyz2UIhc0y2JmAK2YojNblBm6aq5E+O15GFD2v
FNHNyDwjFkq6LFh8y7F29kPYTc2PtAAmjfKwHOEtLLo5p8xSb0v+8bCjbosi12xI
uvx/DPEVeG/AeHRj62vwSLQ9LlK0Nx8pWBdbZ4wyDb4SpI/uKu2MM4xuIKnyqJ0v
rOBqmL7n7dWHMSMFYKtrPs82oZx2x3iG/LNPlnkMG8U5Jmu7vHp7gNWFVzBhqi5q
zL63iETMZ+4Lcq8FqqOKN+5kJWqHaAkcIq77hzxIgD5/tnevV5RwjaMK/x6RJiiB
ukEts/W7xHEkJFcakT76PMMcZDbRziBpsTOGgO4eKKWZHDXoa4EG9hKqignxoCXE
FQ2OnRArg7EXZuQ0Rj0ysCgPpqYytFSRF5c3AqU+YdLaj8cRfqv09cpw9Zt26aQb
UHTuS8Lz12GBr+cI5L+jAAKtux872aSTWfqJHZ68/TVeaLoHFVt00S9pY0u6Ps+a
o7z2FJ/j09emeRYQDXt7HTMoTsRZO3IPfpsm8pt9onln8cSDVSQ8q3aPF/nnWnon
rRl8MemjUYndw2a6IZHgvvWP8joozwH2r4SN1XsanvtyFX5KcZGvOXhiKfjPhgDs
ZjoOaLbAP1M6kfysNX4YQqfK/FZqIqT+cYc+p/qFsgqfIi3VfGKz97c0v/RHcB1p
MMhsIBZNIdqtsFttJ6twJlmHt9hDA8JKeP5Zit4u1KwT7bkScIi7OCeDFRip7Emj
kjjjgBmgqR0FnXtodZOEUpSJmKTLb8OgtLvBzTSQSmJ4Uz4AeKhOBDrcC/JoFvFX
7O5CHOdWAXv8QEZmmgP1C26EX5ofBtsk9BpBFt4Yu4dX5XhpaJSDay5gLTnoxcVz
pENHqkycemtdfpQRNCZ4KYtfKaopwiPbK3Odjep68bQ076Dw/5KIF5DkxxmT2+FA
K+SVFOdRYMNDbcOlsezOMrf4ZRIZtma/2B23Rs7xZIMdb5gv6OXewweolOZcDYLN
GgEWEvu2imVf35QEMM/AIyX6sc9WfNMgMwoQyjDGZBVvWsV17uwsLT/ocjOt1qK8
CQCczWLF2slZ8rjrxx4ZFIHz1NHczTwOyyhcPhguDxjhfwPCpDrTgplNYMenEcG2
vWNPnDz1nwPW1DdNK/PoQ3WUMHt8XFgpX9DybNEnys67v06PXiRVN68jzT5eoirJ
6iQuJ9vnFkcuw7vQAC3DSu9vfJDIW4sJZxfbvzJyMKVLxps1Vv9SPoOVZ4Se2UVZ
SljZV1VpKUSn1lbVdkqVd4Bq7GBTomQH+uhFOnWYQ6IM1zH75P3XR4Fo3Z5MyYdk
z+/UUkKZpG+lV77hCgqpTSYn2LloohP1NZ8qL0T+VzoNJm5ldE1Y4dcbH02tI1Dk
DXXCSfoPwPsMxPlkcgt1a6rgklwlmAGSTRIJd5YLMFB2mB66vIIl1LKffSlfbyOV
Msk8G+jq6qCRqNhkLJpW+lomOqCHWghFXtn/wb+7Rkfeq2SL2V7aRMrcCe9j2QBX
bwcbBPrjI5gXbzlsN5u4pkiKNkPlihE/HxkmEgEuo4e96itOp8BBAXn33Gu23l+e
AmoSy74CZj6VSF4GBhBkC730gTxdP5SaH1bTEmuNnaXgB+/RH7TisYKZvJDnvPMB
on8dZOsfNTF1/cXbf2VK8pHZSiLLNGt70Ld9KiKsd+Ip4Afotyk/aUPOrmpbQK5O
FTUG7G9Zv1M7bvhYs9DgxikXgEdeY7N0ma18RWatPzkMTBXx7hN4XQ0pvYePRGbh
0pWoOEJekL1uy+8Wk3DhDiyAY0Y629drQJNcKkjjNlf3ENDMUs7zGZdDxxmHfBJs
LhzM0v6bklncyIG9Gro8P7gRPT9kB/AAnyjC7+BNFQrVKhWojjdoZNg6i2kkBQI9
mv0M19SjhCAdlOVu2XCrCMbsMMQBUIh0+kgQldzjA3o15BECBjuD2mjoIA4lpFm6
RWdF53SKx3mFSMTmdc0we/my3AJfAsnneAyNPfA5JELtgUmNZ4vhiNYJCr7gvPKj
M/NcV+6R8PfMgdRiNlQpYpHl1pxjGLSo+FwiqapGp2qKaj2Ie5owIS934d83pwda
DufhCLfLZZaL4apv4iKiviEZP/aYKjHvA/N3JK+TK6Zm9qzNcILyCuumsk2Q7zf4
6/7PlorS/Lrrf7XceYHChCrLBIuqoQ90OtGDBzKEkMeIkgDq/kMezSHStqyXuF9Z
g0SUp7VGHHQnRmy6SVEf7+XxlYJTt+P0aOOIUNavQZFzawUFoVJc5JwBloGRVpnJ
mSOZ9hHRxJfo0b83utAPTo08hWMDq090oIGTYZ08JnzQHClUbKF0Dj9Iu560DgLY
SLIFyFHl57u2jBWwqz0ZXbQXzobEj3LqYerkY9258SPdjgMaD73J3OLnACM7DLR4
c7uxEhDGU0zAMLE2znRrd5bj3aiHNLQehGlCBRROybKUD/PS0AYvNbW/Ez53xBns
+7AtS+YWeToHjpp5kTaWnoLq8txLic15kr1qd1XcFF6Aemo+EVhsaVD7FN0Ps3Rx
Na6Vw9uJrKhPHicv9YYiqhbNG2X3OeflIWOqjFBYwmAxRjkXEazuHKKahCR65E2t
JyHBOW3PSTh1aeNtABldfukscoELX2KTdmqGdOxQBWCb82pQzu5KJLyvcEkSTwVi
plyNwvMQ3kKS8XnYDjRlGbofvcL5/zzo+4Pti/p0Zo+jeW5yCREQKOFsLSX9Xv5K
BSbg8MMuvWeHMWZPce1CscPuus1nhc7TtRIVJ2R2eMXdgAvtADsK3V9uPUmVQTun
cFQ4f+zATn8GCshInCJcAOvU0mP5XV3q80J6bedWBbVKS5VSXh6AJIxr+echMnGW
tWL5cgxhncAGugmvvMt54bJm8nrpcx+w1axOaXB+ZE5+w5rZ97s5SXc7GkZUv4Zd
HksHuUWLQCGFn0DTj7MhxKh4FcKc3BngkqdhRwyVtsJaA2ShL/pmG+iIR+8b6T2X
YT4qUT9eHQkcDeBlphgj8Jcww9ti/+sCFf0+36heJn3iYn+pxbuiKIb0goOhqeWN
7wBTIG/AMf1r4QEPu3Nma5jOP9RxVfZtqzXU+/fukc6IVESP43Qju6Ywp/gmRe0z
ZoFJJATi6glGmEXvK0a2NmfiWS/FeZWiUQ7tZ+gc7BjS3tzt2+MXGerQPjNUe0oT
F1U2DNrwCTt9AOYL6dK/9dL226VWBRhULECYydAxeBXc9bJpU+8u4iV21cbu4N7O
VBvj0S0Ax1/MDB3+3aS6Z2UBSrDrRmKD+fkNdPGNzmlfMI4lAU2Qcaw87zZSknIn
saZe/ik96D4XQcOuk7UfUkSIHohTOLiTlJ4kRzqNg0TE+XYsDiG/81rme2jxD4k3
b5J5SU4J7dWSregsneauW1AGS7QJ5ZSgl5uDm547FD4xILj2Fepjl1xTCyif/CnC
V4CJ1aQvUuH0lioqwL4bkx4Y/rr1xvE51t9/3xyqB2gyC/9sOKNaCD9dRKcL4q47
2/jCuzBayAXQuCMDO9AQkgeRdADCXp3ujbxEZvrVLYYrkE74PJ4w46Qy2fsi5rMh
3XhsSXAkvtDYQmsVxgTRFZB2m9MXLGmgf1naB+hoRwDewuF+uFeOFKo+aL9pjP5Y
Y6xF9QsraFWoSldOLtilG4RT8wxisULne+KRc5IJacgWJXDbQn4TY1bLhm1Qvk0y
5PDE/gOCN7/MR159/3Yw9cbWlZEVtKnqJ9MQF9UF0sDc5EE4KmEdKdhtHiWc5XXu
E21IXEpjaZZfHsbPjMET3dIMGZexzUIwTWvRt7QSic7J2zhm6F7/2mSkO3TinX/h
jQVEtyAfz0aFQeTB1aKOD9WS+eE4TkxUxtZZmtzn5KbQtyWlbOI2JmPmhPcA5+eL
Qx+iTFSpVyGjz1Zb6oMkxh87r7TL7XE1zgqLdaviDklQH2uZjtP3bMgF3nK9o87H
Q3kY28oDlpFLXcJ5UOpF1PSersX59T8gqF3jdXxzBtH7fFKbe+Ilu8zb2lxnsE8e
qmCamII7EUC/dkqiB0Hja7gOSWX+Ibl0b0SmzYK0PVs8LUthVlgqrxU9PhfoPGTH
7HzzMfmAKZBULeO6+mdEXIsS8e4xHEkHZvtxJHr6bge7dYj3hylHH08e44P9XQdX
hjffVo9zFcwZLTwQZDAAC1sfEl/EKJpXXwMnbfAT6pva/ZAuNHr8SqLm/MDqM4LC
HyHONrmvsfPXfU0q0Q28qteJlJVpIgFsuF0GP2CM2WX7icNi7UBMcbTAbnH9hHZ/
57kTx9WGYUXVw7mat9GQ23mIWl8IcpRKS1rL30ux2WKZ/9ZVDI1J0FQ/VrGpQV2B
fLleI0P4YCYuR3PYAxAnnuQab4+vYXaR0awvMwhJc/PSGVdJw52FcIgsE1QX+D/0
G64KV6WFxzSQUkL7vY3qULfnkJTTI3GhsanShff8i1DJ/E2UwX4a0VBLUtoDepLW
HNAIZ9QF4szGrDH1nhNkzaCXaC7uGapMeW0oee+KfrSBmuXfMzDkNSf99pCj+Gbh
J3PzMHxB92XIWMxN24zyind/TpWmgtztHmS5X4Kvr+uPhmGcF40jF/vVnWfVB1IM
hfcfD5hus/NEBGpBYzn4lB4t90Zd5zwf9MKljQx/eAcOHKImmPDlQ+Dk1xoOS1GA
jWwghdp76EbjZoDi3E4zKrHwjeOBgwazaTX9o+VLrCieXUHgKoYn0pGJ/jps74eT
1pK5dw3hfv04r0LRCMd2k0WNlGDOF4gTXm5XvjaDsbsrXwQ1y7SpF6BCmSVo7WrB
DPaiWGrhWWS1sCA3Gf+D6WNl4djHfEufjMNFna/y64/2StJTU/Jje6N4VvcOeTzO
lDgebCBFZrMlLE5O+turtgVfAWQv/ZU5B152Mfu6ywdTI+XkVXA8txuhEo7q39C2
NrGCBd6VZW54Iijxw0xT5NSba32McYMYzkLitW2GE5+unBepb4xGjaYURamgXkWo
UyQQtmk7gapmaGTLZOM8K1lPJy9ChbN1DMheQ+85qfAcJ0urBHCho0I1SVpwWQ7H
xw7JL33D+0DeBb9D1MT+3uI4eYoMNaupufWIgqVK+45A8sxYElbHCbalfzfPCLij
jmtneAonWEDpLt323dt7F9RkGebiQvDK+rompU9XwLsFNIQgrr1eO+G9EkBYgDNw
eVad/4XjMvZQMgb5mdCmbCYzpxmZSWgef9y+4xSxCzyBNDBMoAIBlOp8EKet+DMk
6QV0BhCPp1u1UxH6V87/pH4yFM9DecKrlbK3BvGMqWppSbDICoO+rl/5ux//cqd3
BB0kqqMuLKi2eCuLG8+uQ+9VnKSbwt+zchkEoaRrFW811umnUIhz5Q7jK/KyAhRC
v07n8se3byGIzVJ4uC8ZYvToNNisr0FTOrQ7Sk3sgITXC/7nmmCdxrjNd2X1Kpgb
al4E2w0VuYVFMTGz6pb32xRthsvHk6yE+wKb+5zh/NgZvvdwPm8qMXDmLOiC8ny4
IP5cEyxZxc7/h0s6mHy7g1PWkIEZ2qBErTGwHJ40P2ALRkR/7wNu57l/b47566Un
jSINvNPITJfdMfT8DX3TFhU7PjNoKtbssv+1yWNcR3itjHgDn3LEZ6l83jG3dR0I
ElZOFOOHxTOvGZrEdU3fnEGbAjZbyHuATrkqc8jkfsGGPxGNOODMvd9H/2abHI85
vpTkD0UyO2AYH+HFAmk650zWbz3YPS7t7ebbiEgVfknD3ZE9GCUC6ZaVIgHlAXku
Z5NBWajcJz28BqaiNhSPU6SgT2R9MJJ2Y4nwVi0gWgdTCwCEq//VaMGhowKRzeeX
2NjcjHttt0vpXytQnzt5IVy6Xzj2n7ET6tcBbmy7+AM/SMnIhcQWwh88L4i30wXG
W3izMhZfwy9rOz3cepIeXQ7ojtOxOez91Gk0vU8ElxDjAUiX7XGZJOKJFF+iMj0s
P5Uo32jfaGkKyCu4lP+GwxF34NRjX4FdyrKst2WlSLPIwB7ojChDKW9RHivr0BuB
kDAc4c514bbuXxf1O/U3wwYW1QvNfuP1tqQwGr59h/5r+snYWS+QPV0FEZiPgPvJ
2YSf0YflPADfHEPyhobSnh+dpHaGzQXMqRjWbahrhyHaWJfUHxGIseXfrzaiRsqW
un21WhPDopAiYbynAeTXAzQBlIgQW5UtJ/IBvw4WLnnR4ujNBHJKJ98dpuMsX6Rx
K+N3d2BXQQCG4vnWq9nVrMXjl/aF9+CmqMTJn6lc0XRIpQhst32pyTHKuZU0FjLe
m+iIL3NYmSr9JzWoqwIZgkSWfe9bnsTueFueyrDgfbxaSp1NJstlqkncr2vERBYY
F7Vo1jBZwz+0VujpdqZ0jlfNHFDKRWBY1Yi773QrDRGPaZFgteSQEk3a3uuE7tL2
LTxLgXTWtGdOGdwqYs4KG4v68AGUB1kFV2dD9+LwLuxTgVqpz+MNRm/Cw5YHuJXF
KrZhYllnNKDBk3QXu+wDLelfgyZ7svr71H/oGJ1d3Ye7kPuTv4cEpRXCI+4K8Ema
9ot+33BkpEgEkpqUiio07btNtHp33VNPmFbeRa1SQ5f89ep0Y7Hx1fBzRW66/Avo
/S+hJWkRKfVP76zNKc8gn+OD0rNK+b39muD3b581PdpG3DGLpZ0jSaDJ7zx1Mw0k
FOgngbGn7xyxtCo9m3zHGobLoYpM4dh3LMPygt8HkycELdqTVhRieWQ09fil9AeR
BUo5eJmZxHO5PEuaZrGbjKiI2X9hirXFwcb5qzsrbs5wdYTib2rvgvET9XxBSzEa
YtOsp2JJUzFBqzOdAZvJLKXXJtUdnYBa/ROpNxYPYYNsmNMXYJntWCC2lxm2CzhV
gtCj97PcMNxFan3Ff9ZqXbOYaNaWmtVgRmVrPk6yHsqHOrjxoSqEvbhO3QYPiJXH
kj770jisHg2kSWJSkDGYWzOrskAkm7q0B1sKk2YfJU1S7K+WgSZOjSUDeyZ2b+T1
MVyFw4GPHp2QvqVp8LG5EeaQ1ZdtfrsZLCsBWFlcXvSX6Jq2sgXchaj6GlUkwpDb
4ygiB1NGZ/nG+PjckqBv4/bQ9KksN8C4+5C8pUcsGZqme3MErDWNsadG4lNTUkcu
iDaeuJ572huLLiuB5hPkqkR5qtE//kQNUrK/1pIEf5UHKSoc7NGoky+XryFPHfAG
QDHKNV+bJCwJAJ+6b2wxafGQZ0DvSl8fVrk1LT9sRkpOEKLhC5oP/88IZWRTZN0q
5Rda8SplXQrFUzew0egpLEBbvKA/wYorwuDaePeiHzV0Hmd9BeCOkKWYmCOy6bM6
sWS7EHqTj5HmhYEaHgyDac5WQSsYiAZGOvJtJKUHStUNC4lfEHBmMPmPAwoh+pMO
uF5n8CcWMRMc/qJewh+uqVW1gOXHfwHuatVc/3phLDG2NtNNjmIp4AlS+KdWNYI0
4Qshs2cvGpO6q246mC/y2EF28spzuM1ud8jYdoGIufmPDIaJtpWOYwZMGsurT2Vu
BCphFinnx3WkbF14L3qe8T0auFskWZn3a9+Hj9rjZpoqR9F/muZXcYO1xIELAoYv
o1i7eaDlwAQuVzpiTt3fXM9Vv+1lecrOV/wxvS+WK1koEMLsjSvabhykfY2ntrvu
MCvGD/6rQFeKzMcB4Zp8AzhphDF8UtbxveAHfKUuDScJ9hISWh2cSclWRX8RxhFQ
EzWr20O/QZIyQozJbegrsY6rfORo5QOgDgLUUzjpGJLADfNhHIUPHFIExIndBvMm
RdopzHUZY1/1ucVZSmvhe6yHe5ScUNLs44apikpTDWyN20u+4xlmQBLlOKyOFo7y
o13+qnIh6axigRynkwqJAqV0dIlK0MRN/3sprMZ3NBTTAGI1yLgezdHRxyIOEQvp
jMrZ+cVPg98sfQDmZrYEi6zRbc3VCKNM6AUKgLqAjUSLlA03XzKPbG39F5ZE2hzr
ZZgKmkVousVgkBol0qVRkwBgxD32snRL1n+gyegMYPqM8/HhfbY48/CfIivVTiLy
r3knxQhok+GyqlZjouqgnu1Lt+4J/rEe++mRa8k2dq3CIq9kO8eoJWl+I4XY1IOP
t79TYefSx0UU/XfZapJyk0yxtlsGKG9NeCnKj3HWhym4toXh1lXPK5BSV/ISle64
r+HaDV13H3NmOHcBgLD08Rj2/cXdDSdjfNckmKiHe8nXQ3uCjFj6nQXQhaSwH9TW
MkXZSgr57T6AKrKao6K+gm84MNTSPpe48x+SmH80Zt5xiLlMEGbc81nohbP5TYK0
NUtZHiVv+ppkj+0qiWqvWVIe9Ukgs3v5ItUHfOF34z70/w0vd0WdBjdPsOhcfIKx
RGRy7RLtedTw2i/SqFSWsDEUmKzcul5bT33H5bcqAzrlqqm6ifhPnrAjepYX2fO/
n4r83fPYZ4ysxuNDf00cbv0OxmaWOM6TlH89OAJNQz9ivgqfuhRhdY4Q2TfBHMFj
7KnyA2ncRG2LWCwyJowF5KUJXDGnxH0O5Q5dT/LIH1Se6iaZRqvhauT1aD1RJf2g
tQK1FAbxjV7M3jAysyx967p9FWyy3Jw+I2eYtiZczR6TssXJjQut6W2u0ambeoVw
jjA6ilyj4kJ1JeWgvhO0bRvUFj6PJ+72o1PAXUTR6VSo3ehnlljQZXYNZPbY3N72
KpZPTFTLP6xQBorLeSgTSkTnqmTkI+gaWMD7QwiWKsIcqNnWExP2FuPHBHh/aoJs
P8yHSNhTgnkGs8uHYSMwvR/52CEthp0zy5ben5olX4nBRATmtNZWMVfF7UD5+Cjb
3wDYvHetAHOJYNw0ORbx0Mhi/ZHjdolNl7jwcIo9rRfT9scLDPB6ZFRUBVNlQK39
JMdHLk7JntC9O9+lL8UfP8KEanGtzMaMp2OcNvV/JnCYmRXXwF2+BAa7e2ntm6U7
VL7AexBjFE3l2z8vmvHrm53fEms11NpGkdbld743kbjEgX7xqaYotQ951BGz0MUI
jEY/i6Sz6hqSA2ZtD0pFMoENsF5pGO+te5jgdUcSO3Cg3YwpvZUYK3u7ZGnZSUqL
tE1fpq9UQfdwDFswifj/+SXyYSW8exBlCgmlxNw/U5p0A4ODV3LInoy66afV3ClG
G7v1oESDH55UmbNrxvAyytrd7OzWjnmWIdZYiHA/0BFZt/o9qB7kYPqywgx3EhV8
NJqTev6DrploRxyub403EVUhrIP++sHeC9qtEu1IhvovJ1pNXYK2PXl+7rqOQyBN
57AS8qTZHvZO6Ic1YCw1k4SFIXsszWVxWhE8R6rWKngHEtjJr4x7+T7BMVaqZGSe
HEkCPjnhPFUPmPalicakDD9PAqRahhgGFTLt2j37vA1TZEiqwK4E8l1C7QPNyWLC
RYZaVOgLwZ7d8QERTBubKdLFQcJU6yeEg95M88Ow5uQxnr5jlbS298xi568+OhQS
hnEllKbTehVYFZpbChXncAT73hgRCUz14nu4NC1F+wtuvmCO+IGErjrfk2vuiUsF
kFtJ7q5ZISunWi+dH2eQYg1RlsenOhT+hTdLeEO48hhwo4gfxEE9ulqV/VpaH+K9
iaoPenwcf9H+BzsgXglaFEDJtYS5mzwlE/OS4agqiU0WYVHqoJtx+Gojc8Oa10MD
4lqaxUBw8eVA3qLSM0W5E5wxmDNmGgfgYy0otHTj7916AeXNlar9XW/GbF5F924N
arA/eroWFZ2GBCwJDtHVlEiUnybnNWXoPugyQNGVYYxbPiG2Vx/fVx6LXyzXcrLK
ddPOAJxUaeXq8CXnzadmSIlPk7mpQO29q1Igvucy3XQG2iSyfjw42sD2EJvRlNrk
8Su57PoHdJWDzPlVEIBMBqLKomlR1imq8NxUONnTrUqa4CT+AQNC01i3VlmlPY9T
QdFtyZnuJb41tOXrTNQf57bOcuzX7DAEem8JVda0Ud33/91txRE9MxIF11jGZvCr
RPxjoa3VulbtXfigpj1Tr5qWQw0jcccZmd+SzPQFVKm3LSNbAlh+mvzRYb+3UUTp
ZH18QLKalUK5ukCEj43ktNI8PQfVtcWYLytSNyEy2oQUoA79fW1m9bsC+O8MwlxY
XmLwrHSYAMJBPyow0yHhOX211Y9KavXK1bNYg0ozHteX5vK/pA29q1EyJ8I9QK6Z
b8ofT4ZH7GX6AD+C7hgItC9isOW7L+498q7auPHvkTpuzc75LTd7X1xLoF/3yXEM
FT28Miq2O/DaMFIVHg0IYWYULoRaiBGkYqtpyiVOZraVoMXyAQS4n/5zhT0Hi0nZ
Ih6v0WhgafTS5p7ZFX0lMOcflYAXGBattRMXxWnMN7iKkXO+csKALP74nsu5RzUg
3DOEn3qH7mlQHW2dS7gBk1G0wxSet5wfDS8dvkEnwFF1WDf4+zI75B1bPXVv349A
+W8HFVZKzXXx+RaE/7wRFPYgKhA2yj+J+K+oPmgaIC/ueUxx9UdNLNE/sXOeDMny
X/0nycbwgFJLXLxK0kWyeZ+wdb0C5T6eY1wk4YvAK1sG61f17thIGXeBYuKDT5f9
/YiPOhILEcZNPOvppv8e3Jgke973CazzndnLie/21RKqkLKInFTpGMNedCoGmWMD
SLTZAma8PhtrUC03I75+9hptbUMTihZQUAnl5ga5arpGTS/kerN4VGZg3qiIhava
ZyeUeBgSlh9T5nHvl+Y6g4EE8nCZkBg3gwjNheSKEPECljo25SxXmuZ4Jw8+B4zl
jpvF6ZD5082R9deH3bGTnk7NkZkR4ORjJl365YsEDUv4L4JCsiX1WGQ95ig/mi3h
Ca1ZwT2X1H0PnHElroMQUbaAM2U7luBqDOfYAf9hCCmTLWG8rsopP1lRVrIFK69P
KZNBvvshbPiG3Q3Rn8xz5Sq+XuoKue8Mrg9XTxzo94XrWNUc7pykVYCYO/1uitvm
8eCu7lt2FTmhm7LTeU8YLIxiUw5rOo14mcsJ7ekeS+leq0NEZj+12N2mMt7ZghlX
k0wnPcByhkhP+X2/uR7La2YpbvIIyqyKxOQ7UxU+95WPlO5opD9OAvvjSHoERlDN
agqk+E3f1fvzzI+c9+r79iE4DOfEIETOKnG1bXenB3wknqyto2HTpbverkqpB2r+
4cwUYaUI7QGOpEfddNYq5Tx6WI0CQisA4Iufly7Vmo8n663RJjwsLfQtrXixP+Jo
KG7+aGli/XmOZVi5erLf6Dfj8ndwx67byulDOVCc08Vr3yNpX1QDpFP7petQOG92
H8sgU9ka0Dv7OEVpJiKLk83c+by28q0AL7rt7WNJSDg9hRll6cQVNccVxqzq4a0h
r2EzkNVKJB2wTGhw1cF+UIBokQl9RrpY9Wg8fVbxSrYhEktYWXGgbbUSJPMFfmUv
txRuX5mXvCM6RK7iDSjWGquZuqwBlBmH2DoPQCPkvaj8IurOmsLZYVNRsf+Dwb3Q
fKnhSVSYXdN3oNqDtz3LR8B8OU+Olc3D2HVzFP+68FSNrPq5AsqVL8dUbqoNJsMt
bfTy3VlGqItm0cQ7ypu6GAx6VMXtKyilBY1jj3972W6su45HQFKSYlcYQHuDUptg
4UbYA7lmB3FFnWUD3o/jGm1jtmvmlQBnNH8sKpA8AIj0L3jl93VOlKoT+BLJROZR
Oi7zIakapFqGxJgNMF/tq4bADGTyMT/sDMehJYDLMsIXHPM75I1/xOzEpOq/O9VB
Spcg+xq0ePsSLUmw8SN0S3lQxqj9V94y5nqOP25KS57voU24m5HHOc5PdlYyqpL5
7xC6bBOMR3VhglObKgIQ2+Gm6zsXahd+QPvvkkQ5dh+8WbQSdEUw71F5VOaoUYh+
dxr0b2r6nL0tcjfTHpWq4CMsa3PQbpqml/JEDP4TjbNEcgd82EY1hLf+ikl5XO3r
Mk5S5HlvxD5L0/UllmkdZrdYU9MAfKdCKrr/oarXNJdVSQGCd2zpI84/h5+P3HHX
7HEljQez3i5r8R5H6B4IvaUFZ6SxP9F1qhJhQb8iCd4Pl5jBf+0V9uMk3CvTDgHt
zrlE15/c0Hd5HxMTb/OKWSQM+UTyRbNDx/t9LklwHP7MtKVaILuSQPHKe8Z8kxWP
/eWrw1CuBBYOyQxY1QjaJ95tk83H4/0tTdsRX40yqFNGDHk0kM0aBqAGS16pNRFA
MxOITpJi1oHf+ab2SZg6lSv9wCEJUOs+zyOz8mE+OYa76ido+c93mQRXAnkGfj+Q
P5ClNB+p3TdIqrQbc2tsavnnRYur2T6VWDbf3V0p9HHFlM7THnpTEx/J+5X8+zL2
Kk3qI/77ZXmkKW33v+kDhcFfTmBbe6ZzSleHZ9ih9gS0s/2XJdQrkFFItiW9RTbE
XfhWvL/ZCsNSPvhZnV3PDUrKr2HzSzzbq6d4/vUG7IPEV9kW0ZkOHpVcTiPIz6Ee
xVwz9B/d2ZYsDsuii6JDjgLhu13nTFI5fz6iE4Pmey/kZ1qA+PxdcBBhjUs55XkQ
vCaFubpi+64GupOnxhxjRbGalbkPqggnKyynB9I6Su1e0y15yLm2yjjoYSoBXaPF
1iKlX8gg5XPpJoXg/py+L7vS2cngwOQbZ7rJTY/30FnuIOymg/rfd6fDw78Wuwfs
wSJN+5x3JGsQH7UGwfob2wRYmSyqI55OYYX4wJP1Mp5z4aMVWCesvuDUPcrinoAR
PTs1T4tVTBzYL2MeR0XPJzhcW4umQGM5fnSE9Kjkbe5bItszvnY4gRv1VoGtJWmz
v2ulR3cuJg5FqxY2z7/8w4bXMqDXi1Bhye5eDW8BcEcWonq9VXqgAk5/iQtiH3Iq
1G+UnGsWON1NSVT/JTQpc1sYoq+OHxEDOFtQeX3FL84kZMYLYiL2MqUjSY/d8crq
QvptqJrjktmPOYAN0/xUCGdzmekP9X8K/Bj05FCUvKytOSPGCSbheVKApKJ7RcO3
qVII6wQL5tFqeMB1hPDVaT7Y6nbltWap+39hvHks5VPR6YXqjQR31CXyb4gtwUgP
wAcSuMQ+3fE2aAuhcdhLn2FqjrTvtDUAwuTQV1dS4NRDlM2VK/A/s7mf1A5beBc4
ngdhqic4UlRwfK7Zawq/gnpTubFL9lmTjTUmbFnuqK+1ixAIrGIZvwClE/nMZzBH
HpIS67QmUpA3D5CZlrVbUB6LQgTdL7hS7D0z3zYAwvOteWfk1OU5kr3rj9FMG9L5
wNCl6Hg3eqL/Eeq59Lsy8RfU7sNdwu4N58BmHAZaC1ZYaZgBpsEolUHP3qZs6BGJ
5g0EV4Bzb3MTUFT41+47sabqTa5e9rTaV4QNYAIcEM/0yLbRYQAWFWuDy86O70mG
Or4M/YHjPOuaipyF3Wu3yCA1jeRxuXgh4vn9rWd9SnqCKWDiiNmED2BcVX5OhHQL
fZEthbRulp3e/dgWudcnc4A4zrXqQZUVzaTyEGbHIgb18LgITJIwR1xq+AG/rDx5
RS3v5rVjYNlSuQqIbvyUu6IS5oO1/V45b3PugU4CDRCuEox2OyL24OCpxNCR3f/7
wIBePzMaQC4BR5IGBVDpjoEYKMl27b+3F/kwf/02nmoc/xIxs9EpMp1joVD2vs5e
V7+du11uZS0CoCdZVxsA1NlNsLnPk5bMvMWEzXmZzU+jaVQhTijhejQUnp906rhg
yIUP7gRhc0xvQmQACun9U43VKOW2JBGAvvtXOtp2PVOlOpMDDf2KBQ981JfSAmn/
K4TbAikkjwu0GNqNLNaLmDOR9fe/mUGTF8Lk9eRDimImuOCOXSZjDWGYny4Pmj+n
Tkz3adPOVJgn5qoDRtqafmB8uh/kochkC9EE0To+5kgbBiBgdo7UESrJ4G3BnXAh
O4LzNSvmcHZEO0kZlSdUMdO4yJe+KwKFkdoreUnCsQTwuKqVkyw5JuUirgAn54i0
HKg//PSrGPMQsul1yiKlSt1gtS+BLGV0bxP6nEMm2Mr6k4RPXuaBkYLPh9lnPlid
2t9L0yQ/EHGlngj8wV78zlDsanmyWQQAm3t6mhMFvqQw9s+q49+GKUvTZNOD53n8
QxPgLpI8U+E7/+SYQHbAsq11aKEc23FWTyShBbacY4FXSxAqq8DRbkGHToykKYwi
wjtbHW+BLhxBBfDuyFnmjcImd+TZVDSxJCqBGwwTIlekEcTFBNhspYTxuRsK5bh1
L+Z7QpNamUMO5/h0xedObfrHsCNtcKtjGS0ksppsA/7Y80wRp1Ops3pHUVE6qQdS
mgOk1cpC//4Sw/dyvvofX9e/pgYqdb5he7SMRFpZzvbi0/wv9WhoBKHjnFIrUmfu
Ru5jYgxFoRodKfsiQEtCa9qNcF6j6vdvt4MimYbQdbVxQLzJWj2kDgMGvJO8zSFN
vpmRsYEWwYk00i3qqsMQtbXLRyAQUKS6PFVHSHG2Zr7ETjLlHN21IbKqSfgBkhqf
kZtbGHik4HivB99F59nUxhC2yHEIkeTklkIMuyZJU9dAilic3uQ+KMJn8/Qy1h28
yjdoi+Rx2ZaT/PQUWeswk/Fxtn+LTdjXqGBsNBptL3AdNxiS27S/X1qoUsuzNXkR
C+WyoMNCq1QUqX6Ai2RIAkfjtVxzFewp/j4LpqIIeMl7j8+o/YP/pAQK8jONJCRC
qelhnhumJtYqT36NKJWZtFjgz8GoR+xCIfWx8O5g9Cp2tcrRP/Ys7I0cY/aJuj1C
jSfwc8ZE+K1dySWWFw4DF3WkW9Hdi0ad4mkIgXk2/OqschpQL7NZZh69XX90HqAJ
ZkEtMrz3xj+knG8odllx+tZtFGb9dFag7iqkRNJOqdVEbtfOaI+84JZHzmvYt4ty
ICfbJZpXsfKIszwCUw5PLVClCybnA4Kk5OE9xRax3iA4inmQ4YJlMbTiK3KsJW50
iXACp33IA7qhWZwbmStRr/FzrehwftP5tTrUc3oCFmAB5MamjXhvg+bnB/LOlywe
YwqD4b5vCT6Pp9nimgwXsUz48shFpRnpJRe6Z1F/dwNngRW24CZIfLl6PWsVPAuR
RIVHOdoCqKJzwfacAnTXQ9JfD3PTp8XDPVFdT+DNPJ6Ld1AuPBt8V2QvUNLwGpU2
HxbFH+ik/PY7mMh8T5y597h152JMDm/IzW4dIZ4IQypp0b0m7SRgg+HNQXEvxk1U
PHWpFnh7pDG4g+8dskldqfxg/0wCEqt/1AnhWja7JvTlG8e22lV3kHvAJBDb/InN
rXau+Qayt7c1DmpdAdo3tMWji5+cyvf+ES/1YIY556xAkY/DhC0lUVrTxNHKlKNc
Vgnvj1+tfM/a9ifMo4D8LWYaOvSGyl0V9bompY3it5OwmFo6W/DE7wG0NGCjKbF4
dC88w1Hq+M8nud8VlDgz2dDNALGpDc3EvwFQawz832+piyKPZ+NPf0/XIj/ApLgR
BgvqtwywvwOuCHpiCegiwOM1T/SmvU8/TfHalonClwxTlxhq4Wo4AaiYedKv+Eox
bUKP3FawEc69exNw3PnuhOqo0tXEez6rR00nkjvHAq9YZNs2iKPvffORDUOkYXDS
3Kzt0jkPujd/6n0hvRET5rex+Iraz9782AUtfb5+btWDqLzJGzHPqwTR+BwzUEND
5Eg6u1PGeTIRcDmtVw9pM9j9M/zfFDPX+0YyQAzhXE2M4O2L1c34fO0axeBfXTAF
8y+zg7gISrlmEDKPpe1F9ZMsb+LQDsHIOsuQMfb8saulMU+bIS+8C4jOHQWSFVyx
hqFmCwDNiqndA2XSkIQDx9WYP1073USULTKynGZCvG4OZeEHxTHNSNUalNgI+vlb
mnDZ1XuV/LAupuBC52EC15ohvLysQcmuZu/xHiiMLk0EL6AdSXl9MxdP5epxCGR2
k2BaN/mtb68/ubk6FqoP/szipHM4J7l7VTNSBzDRlrGrJPfqg4AJmXq7gCYB8X/5
vU0LhcAWx2xGhBCGyYpZTEmgALgdzKfWDM4XI9QagIdmrZv9unw1y3LHucijVsI/
iDJbgCvsS8AX6rQAJZDdvjvng+cGHM2jmtiPId6wmyxtpnPSYTyRKzx1hi2oY6+O
fvN8CqczDl4Pj3bwqr+478xpsRtunSOtWecTpFIEvgQz3OLWCsUZxoQrNGnhTeun
vWoJg5ZhW4tj6kDB8KODGMMfulT31mU+LBVaWoZzuinc1YYcTOg4vYkseLdOjSqV
dWNZYX6Z/5lY2m0pZP9jRxN/wK9pCz8sW43HkJO9potZrxmhiBk1iOCTj35Fqw+V
lBzVGLFXt8rMZpSvh5YD1BUq2GgtGo81GvqUyZ/oEpaffvXLZ32Nlx3Otu6SWi9H
9fuiAu0TnqeuEA85fN2DGoasA5XJt2nnUJyt1bxk0Kd3hwxjF05Gs51wI0oZh7A4
B6LM2SxioYUzTGJBDjtWQW2so4QcKYXNZ6vTQIcuwFK8P3O/cN+3njR38hjeUGMg
+oJti19j34rvqn/tLYywyWfz0L8WmBEH0HJrkzJeGkXMjeS0+BPGaW6V+ntS0jMs
bu7GnnJs/KyUd0O2qA2UdceWBTc6tK1BKVXBOzmcsYM4aE9/JvDsFYim52mbblim
n4tm8FN0OogTjDRRTyzxr7HBE11OeSBwDV3WPfeQtzxCqB3Q59Jo/IsIfn4lRxbo
IAfqkrwgfNvF47/vu8IHVA/ALEv+NP/+6VTeEZVkN38ewG8zug9NTXEcWDJFKWsz
A5jCRFCs1lORGdUKpJ4opPEzZhN5eyGaQBfJGHWP8NbuSEQmWgfeTAqiXzkXAX9v
7T9bnR8/jgYntMcKzLYVBqlgxRJbc15fNfepwkBeKIV/vhBxcHBTDLVrqpIQkRbU
l9xdeDLW78xx60Y/BroekvLupbpReXOMU0jJMpM6nslvSbwAVruytqHPB5sdbmwo
ThFKwdIAUBVRU90yxgDXq4lFdSh19ZKbbfgXR+QvYAAhX16i+I5UVnwKLZFsrShq
ogaAM82Q+Piz5ImDguod8p6DatuGpFu/SVv7PCPuP3KwBeWk57SXFy+AiQEV7NhE
8foChPNc6GEblBu0Mw+os1BSQN+Lxr5ejZRHPQv7J/Kn3exMYJixPyTKM9bm9GhV
qx6tca5RSPg0Eq1hMMswNKPnvtaY1fM/1XmKllBSHVNa9TdCcKTrnzXtp/tMiobj
8kZtcxyg4zYzM8TOElD/z6oQBdc2GYugSisOonFIAsTfbQLjt8K1+vBso92bJqM6
70MLIh6gg5KJwcxrjb0TQDLOQvNjSEpuT5ZA2j2T89Yw/gKDLVlGALWi6bYH3mMp
JHysq1FmPz9Q/XfrmTB+UMlceX5GKtGfXlTwU+95EghswcGQyZZn4vetN2PoRn7o
6skUTh6ZtNqUv+ci+uuaoaXglgHe+XIlcm4YyiyHoGCuvPBwG8PBuECmScXIrcRR
GCyPAqk6X0YOCKSFbx3HmtRafgS4fovz+ra49dVldoo/oEMWwvYCJYwLZoH/tBbw
SPyupgtUQVAUzzxSgxHUtYb6HK1YcA1UnncHhFMusrkbwn2H53CDGUMKEToUsx/O
bOe+O0sZTXmpxEuB7yE7/vYvGLL7ZKVXPvaEGABjb+gkt/RCzOH16xS+WXC8VRga
Z49w6as4ARpEja0gyRBW0fXaQc5NuHtE4bu3X63tcZ2ZeiFer5uQfjgZaEQSsyHx
OnrLqSV6tKaZk4t3XoILXs6cZ63SNioA5/l86YTkoqCvqO+ilAAq7K6eaLYAdfpv
TLHcPDK7zrv+9YE1K+suX0wcZJdv31E1pxvZYmksE0/tZuFFixBozOkOn/OBODPR
O+A+fRSsqN9hXb29VBAos7IZ6U5JPSOog77i0JvsILjxMTP2OnAylYGjAnYVpSC3
tZPuf2wLAqV3A9ZvVppVrA4h7EqA/3EkOja/RT6W1Is/WfcLgkNnWmQfaLXBxdj0
soUOLY+CUOdOGyChUARzmp8X8vqPFUU9PXGsDIj001v8p54A/DldeUfzM6sT+OnB
doPy6xxlkwYMoq/Qv8D/hR/V8t1FStzTCHHLG+4bnDds0HMG9a1+cxxINnbWPhyG
2DBR83EBu64IahdCthZZkvm1FnJ0X4/BofEa7zShbJN1tcAc7OzvURh8erzLkaJ+
KLahxSfEM6N6FKtaNHXznbOZIQ4gkFdTTeWRy9168XM/xHCZDSzZzUNWGVTMF8Rx
SFt7d8eikscpJOBsqfYNQlpWeCKpMBRoNxu8PH/VU3WLFRUgb2dpSftOW4XKbT5P
Yok8X2pAuYDGE73p59HJGQThPK6GMUUTZeQWCDyltZchb4hPQiEM8XBPnynWQY+6
sYNjGHwtomhvIjjgQQGlC/fFdKvzOJ5jsBhy0z1Dtf7UwJv416xJFUV8GTMKbT3T
QfpfOA9Fm6uUtZXvklFCgeyHASGHYpYkWGFrMt7pfWaBlUQp5stkWkHRs218j/4z
s/MVHPlwYvqmR8AfowrHKRmTlvrFwZL6zXbOOHXJz3Suhy3cMPvntds0JpZdZ5Ym
iE90rtbDhq0HPOilZM6TA3Zk/dCAMLPtYveEQHiiAPlAUAZmkHlkwFYjSAvxv6BV
YABT2mYeKRAxjzKNjMl/E9cVU25mNGOdjpy5Df3wX19b4eqO6YLHdFRwB0Bf9q7g
DqUhWxm87C9Xf5U07vqL1LlZIKZWIkb9v5NsOmFUjvkhL/fD4Cj4DxOSIMKh/i5/
YolggPS6ZhZXMpRbTdZopmlZ0XCttoENN0eTbXIfwM/m9aiDiIsbiRiAzAJ0kvnk
qXeDZaAA3/mE7R8TVEc1c+4i3208H/xlwBa+le8LYLIQyP/32KJ+Iab6BOcK5v0a
FeQ9BeOvPqGTXagG8O+uKCJx504ryvKyt7dEZOdiypTnc3xb5/FVoLEglXoh1KEc
jPIeUkAIb369ffCP5ex2BByxFhB6FVlqRdTbwqLj/dhBJ6cFMbjqZuD2/A5X7s61
Nq+IvyR+kjsbNwZGSO/OAuvD0FStflycYLYXBqQcBP1FNnV2YnFJ09w61bYsiNz6
oooGnURXVy07+1CzfXO6x8725eP9gMhAYOk4ccEIyPVpgzEV54lfXyxC561YoOJD
6nlycyXNm526LnO6lpxnbsrOPo6HYI2yKxvk6CcxcUmMStfvYHR0tG6N918gsqS2
HAC7QFupwbAE3GlNtH8F2d2/UrC+KwvGzJL6hMNE6TY+vb1jQUwq4M53MGrmzERn
9aJ+CH86gHmUYLHzzANY1MHn13gKpi2LMPLdwgGyJdnsZSTi6DSIgDecKl0mYTO2
uPrxjT270Vg8FJlGikX4r3A8n64qBWLb/AGj2qfVUYPBhlAA+PmrUDHKOtPDUZ9U
UxAACLX7WTjFm4HNIqyPOpzCL7xNC4TO4o1vrlFcpHNcAkC1KkE124rQzycaCmBo
w7LEAhAI2EDiaotYqyJNvHxlL/YmTHEdPJq3ryt8pZLnsBlKFIRnYvRDE0tj32lT
Uifs83f+Ty1YYL5uw4sLrc1SRpPV3FvklVaBPNd4Mut4pCWvhhN6cCf1bRi1CuHN
QNwuN93lNCvOGrgHs+vnJc1D5Rr3ZUJd7b2C92qD1U01fcGR8bKbzCryLffFJgMm
JZm8obYWRWlF2mVYY+wOWyWdjYi+F9w3uFA9SeqLy4ihkonok0hZ36YIeHmlo+7d
p+CAS809QlElM590rvKiL1/PZXqWstw78hArY3J/ez4m6SmDdClP4imwNZcqpxO8
5BmhTOaE3vv40JaJrdodMPvvLEUIh5poYuTwX6fHBCxHeCmGRMZ1+Ld1k2VGohJr
S9eHKgABQOPrwtCxRPaJXXY9raEclbSyjvciJER2aEysOSZQV30gTVX6jEc9BZVx
QlCK+PPU4eu0Z846Gq8D/1hVGnLtiMTxe8/VpAb+dyf4sYJ47vMdlrk742Eybc7I
6rGzb+FFdHB1dwubjbezTtPJX5VUiaGYj0gKuRaA3y2J/50j+AhJ3nUp93ZQCgH2
bSb8zVz3SMFI8/evquSC7mh1xRhRIRmh05x6annvX3JDJ18TQYtzYVQwE2v7oX1L
uv6+KOZRWwq7arPm9NTlPE7D4BiDRSSg2ov+56K2DNdx/Z0HdcabcLLhgD7qvc7f
b2HtBc+eNvg+kXtk09OVHV400L3mKTvB/Ifz2xnmTjeQBTGlWSV+2KcEv1BG9HKz
G6dVhn7iLqi6HCYdquPVqVzAtmxA0O4n3nNwzBZfcyvT7a3VpQfz42kc9kWKiei8
2Gl+ZU92K3a7IiKA7q/AIOMFYz4RIOX5Cp0Pfo3tufcVP7a0nRjiKLzBUa7jRlSX
n2sTC2gU26wWAZcqnQDZ+26wzqxGgBdbf5EhwayPDpoQ3ttwReqNl/n3Vd5r8bm/
3Srs/hWH316QsrxKRXNq2W+sfzYdWkUR+XHuR3OdbOorQv0muaf2Ux5m74fjx4GP
010dvsELqlb54Ta4S7ZV9k4k1RBkJBCY5paeInVJFgTqtFUshmaY31MBOAHFP+p8
eT6Tr2P2rPCnm1S7qSy/iR9gjrbmClkHfYIMoKaCPbhDgpofvVou4OqVxGjiECW0
Zmic3wAAD18saRjDnL7idMVoJb5w+24AT32KEhX2gch8XsqaoMaEflkKwyw2zZKt
/cxc5Zi2Jjtfo4D5k7W7snAZ8Bw/cOsHHmvkPgQqvXhASMRvP63O97HmM7at49Yq
+TMCcrN6LlTdC+hi1PIwJfemlucS+U92T7tzBW6FbO0KBII2dGsHX+qgVFRoYpuJ
uQ6IRki4nAXyZN08jALUHZVUbI5AzuByqAEbiCSMAedR18VnbpTt88pr9Emupng7
ppNlSyM8IyUGCvjbX4QgFuzkbmFU6RkSGIDBeVWdaY5CmF3p7keqZCXdvaCFFYA9
fygK0gBx5XvsK+nTp+Ct+NTXomnTsdXSWNMslgPb8k7gaV4M1S1xrWjIxOoNZxMh
K56IMhPzL4f+oTqV1ulfuRpamVo/R+oUHF+IqVPCpyWFKyWxfeq3hNeX47FBdfi0
GW6OBBA/nOr0BWlIobl/y9iNksPaccQoWG/nF0GyNvWPEUagWuD6sh9LcWf72NB5
R+Ot5uQQGV/HxR8KL/iWsfJDlAn6Vyzt/Spx/FLANf11T8hz+geSZaIEa1QIUHXw
MUK2KxKLA6DuKVMuMgitZBHN+rp3C2RM3XIkOqNtvuYKeZvTCgvvOJjmkZ8Ns7sz
06KptxBuuh0ixlGFfocY8cs1l3MGsi5g/nhc2HxvAR3z/Jr67GWoXA/sekTtGq4q
tkpuXafUtLdcr+OaTLhf9CsuajzrGydedYOjIPCgCpH+rvv45eCx9RJoPv74WFEz
W70/9tYdUHVD+CnugtMOuY3nCjw5jGca4BTcRtir0f0I6yhUnGaeTCZW/hbQ0hHp
M1hLBhA+SbIBXid5E2PH3JyS1dNeZ3RNCCO8pwCVIaHFq7+v5/yp7EEAaD/DwOJQ
f/5VfI0YojN4mEN/OxQuwnmVQizMkLf/N4gywns3eGGomHPyZxTGILlh6L1/b1bS
nnz1C//WIXObVhc5wZi5o7qxE8KrKBUo3XC+m4N6xgqxoOHFVpfHRTR6I8SMNClj
Bq5ovos0hcX4vAA+nAxEr7E07euC7RFxOKxwza6LHxYvJmGot8UQM6YiZ5nUacCG
jLrkiPe1PV1oA83+/3VdUb/LoINGTd49qKJn1wfFoWDIXMU/NGkrVWOXkxZ8y5qL
BwJAJVVz2MLgUkuvnE6Pr7jzZ6k+jmwnVzLCyoWdr9OVv+GMlLBRD0s6oDE08rbM
Kgtd/4L1LBua9Ymf13BVTcVWjNRGkf+GEMRZWY+mFFJHiV/lvL4qmXsC9ExtNdNB
jJHmkj3POOwjmVC4gTaXX9P8JaKoIR+E9tJ/SOmqrxyfHBvQ6VAFm7pU67Il0c8Q
zmpLcQCNoYmGPvjYF1dnXsLP/fDs5MOEPHC2vIGOJXYsB6AgIqnD+NVVTAjfLtTZ
ev3wKt0jc5tkFAfLpePlivcSuCMUney4u/CsCtY6IyLoACEAGv/YSJdD7qJft9Ug
AoLC9sGWtY0hnvnRKtppUuoZpcUJzN69rsXHLRe3/yFOWP3qkJxMfPayMWZvOLcg
RR6CLI2FRDngJkcY9jtk3bLjvTRWJu5Ph1inS7x9+bGSJ5yElGKjWXTl2Nl4q01K
olRRW/obKX54Ffs2UYCvRxyfea72x5B+iulm6PlHje1qgT4acE+BpcSHodjXmW0i
PuAu8yiKuGvrvIc8YMMDSJWq2KiCqOys+qsDAU9AjCm1YqB01sF9kpItlFCuHgH8
vszn/DWJxg0cYZ2pLI45blDXJTMbva+/47Ycm0SE2BFYY+QV4sKCDB9qPxnCBA/W
EjTit+1AuwgkgK8tJEe0gAc1e1HBa17D0/QPGNqXroPdsctg3DCUV5XwuT/UJjDl
edIXc3NbCdtZe40VgunZo1/RTAxs4RNZHr9dkWFJ4xKe6rqdDpLI2nCfJDO30jN6
qW9yWUJdThH8dJAD5JA3exLB7q9wfOatuiVY8ltJ3KytHDl1Z1PLrwBYpeJ2238N
+MMSM+aEibjzDmlKYi3Ev6lNc1a7hafHxlgfVb5FSmQfYFsSYADKYBWc6t+/zSbE
j6um91bD4mAd5hsMKHaRIQjb2UIEbvYEe3lEBIr6E+UERWVRxLkxQzesE26/pj11
QYfKPhUBW3DDZ+YhmAlOqxAnF8BMBfR2ig3vkMHzNkvzGDcYOifG7oZkhDDXUzKg
VORPTcbPIlzSYbLNxCY/sWdoc0wlTVgK7JEww7nNF9C+/vaDhjFLSWbDKwbQK+pA
eFbxnLV6oH92mN4hijZvaQclrpG4pbv/OSsJ2S2NimT5G+lxEI3kr4AX/TdbjZGR
ynqa2mUKhYeKKUWr+T06QsjI5IgQ7aVzeCdepx5/0JiRG1CtU4XpqRb9R5EJSsoP
KlbUMEJvdE9QhXyecF59znCiBA8bX1neY+KyDjRNRzwAyKIvUUbDnQxaXYdjEDn+
IV23s2NDqIAtzpQaYiclQ6YtVf8FOYjp8/88/JYYJGZIgkyacbK58MPRVH+/9cFv
vhsDPlS/11OCmkQWaptbfOyxZrLn3sqtFOoT3zKXB1X4BVfzLh4MVa7rwjFUXNx1
QTXMCIMNkEs7+Qn1+Fvmbzr2uE037nTiQunnEE95BiCwYtEIYk4+zP5jl/Q9osW2
66vnr+yCF8/VuQEs17s++u4FpXm9eb4zGa8ai2IE+pL8xYuP0gsptijtev3DF7T8
T6wv4gktKQ2iAPhovz71g+RdlI2b2DKiZgGQYsMUHYYmmkxynBX728k+UghvOZ0N
Br+2hVxIzR4NcrHK3uG7PBIImWxINSwhkVh7mzxFvkoCfFgzDTtXWZneEg+PSyxi
/Ahhjt4SnfD/rkM1o3+G4Fi2pSxeV5v8tpjAEhQ99KciKqg19LgcsKFE1SbDRJsy
w9LF1Fmci2+c4IpRFgFTfisSJsrHpcvGFm1CxouvP0CRcd5DBqD/tclEHzo8uHHE
izot37ulMZPpnOOgAo0ZB7V6f9+RGCN8PeLoHuhJHHbqVaVd9dH64Zf8sSiZ1yyX
PkfeS7c4qiEpugRJLDSk+wSLCyOpXi6u/J3DeTT8YEYXjwCjr3iOU5HsPDikSr4p
NYa9f8FRpk1h8uzsnTYuFrEkndmiebxEtFJ0oSQpuM3UrSjcMdKAIsM08fyLOxeL
jJcEZ+30vTmhqaeiPIKoEonCYPUsF81h/lVaNvXfreYCmmeWB/pGxI0i5EoZ5gfj
x7usgBQta1wPDsX1+rOX/w/hktGRbuF9MMhpkzAwyc/0m+6WQ3WnJa++353M+I3u
SfFufdPjsGGDkQXns6ucg4tNCxrU7IpLLxzZhw9DOXSoi7X2MKs71MG/00djezDR
gcS7Y0tdfGuIOkIy83c/t8tlG5aUGx1QyzkS2wbgY4EBp9ruX2vkG+9kPul1qDev
SzF1mLon60cbn//ZXh6hoBS7Mea08WkZkFQTlM1Zs0TpLNE7tk2NCgdOVAny9DFm
po8OMaDxP4gixujQMKZRcwxRmU9AyWlHTkor/joJfDSnN08D5VnKcsPb5i2H4Pd5
/HFykSpJ4mbq1ghmU67Ua7PecrJoiOPtLBcDLuMUCeUFKuuUIISI9xpVKtyT2v77
xPjh64a+wumJeYpDv2UADw0MpOyjF0R5kC1WSXBc79ahtIB8T1ghHxE9UKe/6EDp
htT911AgyZR/bT5wMsR+1Bd3sbJJCvaWdPz9ftA8pQdqqA1/cDv+UTZLA4gBs7/9
XMxpY+zT7GMg8eU51rFlONm0PlyVIbLtdKAHLNJzuR1jUOEGw44/ehnRVenXVgFY
qegv/y+kiJqnjpvRHJBbQX0NF6S5lCI9AgecwlruT2as3d/fhtR5prPaHMPUWKCP
zWNAzJNO0e/T475AEDkU3W0aBMaGQNhveT+8JJKvsjhLyqW5kFU9XmpViv4KOC31
T3jHZLTOUxVHz3s2ComJJZ2YZSOF4PpY/bfVxftK17v9NhL7ov8d24oPWgHTgzYx
g4ooXvf/bcuatA+6JYbuLcKKiCdUE5GtObSiT+wAgruGVTxbPouagA3fagtsHzsg
YAmYdwnMr3bvlULTTnxZS0qVs+MIdkywsC/MdDtzi/xZV2Ekg+Od0QzYiDvyvBuZ
JQaAiKIaAjdMl/PBdP0QSngmn/3kk2EBmBpGWFLqIS0RGSrq5D+WkAJkfjeEJNKG
jwrgZWyS3lS0F15goIwz4daq44V+AeRsJfM6EZvTULyIOyF3WmyvJLQPwmmguFZ1
wjMbhxb+G//ITIcRhC7uwzjNPZQvq7ok1I/QzcR/Uovd0SF0bAcIRl3m6B5uG8Lk
4SS6XAjqMs8C8uDS1aYmWaAcynJ9sVYsDzvFTy7D43cO1IR4IwQmX/S2EZ+8rDvy
JjCXEHf653yxbdz19+bUbSuWhUIUgHNe6Thh1S6N41Lf23r0Xgb2ybAm39omPkab
pqpsSv3VE5DBFBumyvnoIgt+CLisAZT0YDyFAd3JazDiATfh5+k0HHTnDGQkoOsu
QmNySUTBXXEzmg+Y8MLbBE+q9xC+PGfIXzm3+Q7jMyw6zGFrTj4DkSWrXqResJAn
ad7Ms0df4kE7Q1r1MDJfk1vskogsAq4LG5djtTlO/cKIblVSRmtBcMPdnJxCJwDI
m3sdTSqdHupgCqvjWLvX9cQ3UHwMMuouw2zUIjljRNwOM0D/rtlBRZ1C5u65hJbN
tL9+1p06j0RdeJaCFJiXcWz6RS4zj+XKV2hKWhpqkTUUK0VJ7eZudrfQHiTya4J+
DssWTi1cMq2CSKRtIwZLbejAIFwHfxgd8w/bzFm3L9FdsFJ3cQBwaOwzgmiMZt9k
K+NYUWZ1NCkhw4Bk1zQsPcxzYeyB5TPelZOA1qXylWl1CdX+RJTjJV3Pg5wDyUcY
lDJ2fEKWVOe5SRPQjLkbwKK1kIpOLpPPuTQ3lbZSFvbKHd7+RFQVi7zKGWnwQUoZ
uCCpiKuRM5nus8rsQAUa3+gHot6qUOLP0U/v18fpti73vaqNb/AZWglMu0qkQQcv
T4mWsuZGfuKeyuTthKbrcD530pA+thQMap+OTquylQ5fYQVGGLqF2+q+5/sZoTy0
vAK8/YSRm3khYIdr7d/2H4fo8gXJHQ36uuwk5P8FnfvxSSmYh6u3Wb8u+VVx2nxH
bB30NNz+X9ZsL+D4f3Mc325+hpS7y7CkJOFcVYXzIKd46MO+lpDP7WCf4XRPM1Mw
utYiGsrERTyIol+ALaKyQwHCKvulTonlt1H4pWaZCYeDHsxHEqrbortoOY2sUIRk
4yUTlTPMCEYXqgw02fSbM7bZ67ScltlhAfKyi2BwlGKxgKvp1Ab/uQ1SP20AqJS7
xtYENyLVRm886CLD6he0LGYG/Zf0zk3BjURQ9QOSRaf4dNd0P961UgXN07o9lV0/
dg6UVPuPepCDcq5lcosPzs0eLz0X1ATB99Toe9H8TWGSX2nqcm9nDmSq/d6SNQKd
skAqnceuA6y+t+8v451kTJWjG8lF1eZBuddD1CInQTK7q2hqZ9jqgWHzV+85vkXz
Pjyrgfrd/C0GpI7i4FozKZ9qZiiwxECLHJ07qF9pfSmVU+64AQkDDgTCO0PsVXe0
sw+fwZdvOyJcSUiYDdXbVi9CMZYYPisQYb11hJzwhyfZmqVeCInpuPx9W7yD7Sjy
qBHVGv5G5rc20ZCtNVCAVykCYWfkIRGnKBCmMtcURpFwzshm4CCm8WtHednqiP+B
WTlz5MimnuVtSjUvh/hWOzIeQeQKLIWf0Y7lEzE7iaK6GldpJXeMJqYuUOjgkekF
muk4r4GDsqSwZVPDXMRML7JBFojK2obbVvxDgZ/3B1rY7psNFoB0milt/aJJUUFb
Ogqrp1u0232BRaDL6ZYF8HgCk1IOzO4+S4LU2pg9ES28T3lrkM9uNABp5YlQ99DS
XfdQ0p29htX8ATuAEg0AKPhTOtihb2UIZdsJPM73nlKVFg4DqUJSzn4fRZo5u1r5
D3NhrXShssyx0ocMShEQFDx2COZ72B+xPgApYaAHbF+iHpW48sa8hdvS7TMN/XD9
vbFL940/KDqBg9s/SDtqy/mNZjm5QBXGGXuuAk0i/0A3saxKiicsgTTmX6xjU3L1
F4EWMAXTBvHy0l0dMG2wbRs25rH7KEknO8zcKxE0dA5YJ/s/mFGADKUm8sjpbWzL
LsWyWVeo4LFgNcs5ci+wUS/bfpKv9bQmTVptQE2MGw/aTEEwM+IWdVcyOu71ZoHR
C8lk6wC+bMF36G9W06SlFfNIeIYsx/USssqi6AJwZCHup0A0L3eXsEo6Q6yP3m7U
h8hNdTzvNi9m8EBYNxnM/Zx7Fgos7WNCCN6KqwXXo0d5cD348RWnEZ4z6xBvLA7P
TCLPNEU+jRFTgZbMm9B6jAj/yLugOpefTzC77PYSfR0mR2AFciM4fyIUUTShlFNO
19q4LSH248lvPIJptxwjk0eIusvN0cYVS/jMxepEefENzF8wkQY580daaAJH5eRG
dfjBQCbW+b8gIwIDgvYE+Sc8RYYyrr80TW72QqryoU1z4mJIAMqiTRhF1GBKcGlB
qh4Wljivv+ifKl+I02vko+gLzQWFhIALEg6s0Q3Gs/YXVh/NwF8Ww2cJN1zqRAEP
Ksz40gjKs6fVVKX3vo5saXwsm1OdzMbxqKRfsh/i0xroQIeI5UpzwYU/3awiM9fJ
QQmwlSpeT/msGPniGVYfNYKGDqdpq9mHCe3fN5US9xctN9GxPrJellFiZjN/imZN
uLOFkhEnwey4NKbdneR85S4GvI1AvzevHS5S1j5lluQSPtj3+wZHylJV3Do8oGjP
Vh+x9RHcxutU8zaOSAVz+leUOrxDil5ZMvvOpzhBmKpCw/Z6+Yw6ovQDW/Vnh8WU
5+Fmu/2XSU7flirsFcCQ3LTb9XV5ur2JmnMM5ODwMAgOKwZh1Q2rqzcltg56Fgvj
Rkxi0Kta0S7tW/kytW98bUKR4kLRR6tT+jqrLgQ+pgz/zOFY+KlMSAQtjOqVUwJa
12+obAVoygqHoauhYx1/ClpPICCDpUsMgWn/R5GDsLgDahRisEf6T0sP3rdAuA4K
skLZ07V8ZIXc7S0j+k8zvs6zubAGLiCWEGIKf1jKJhiVS9gjqZNt4Zs8HrFUPQQl
eifGmj2jGkICeE5SKDfmjE02bdnkzjx6evhSy19gaOxZFtdkNHVLVlG8C2fFSz76
UgGbZ6mv/+ccFZDLR3WMfLP59QEA42Vb5xpEEfaJZfP7Pj1vdDHcJ+wkUlFphMJv
Q9BdQqdbGNt5I3CXfTVJaCVPAVJ2lpSTjr9RCu7NOz0rrl6Aj8jvOhxOKUqSbLrY
KIrxy4Qmuj0eLx3jgAuhhbKaK2TD0bpBGW8sv9lNAe/IacEFOIgBUJC1gP+Wkavk
VaJo6tUhtSJECYAlcY7uV9PYzFN/1suS5waPdXj7jg+jlKRC8f4kQjkXv5bRMe8z
Jhg2V3ovNWsrDfHzZZY6dF/HptwVnNluzQRR7cN1B+Mfa5K30Ki+aLgxN2Ark07Q
TbmEjt66zNJ8MweKZHOWA2uGbuMOJxskQ+/OPfmtpQN5agq+ojvoQY5lHDEygVlS
bnFgvH43ovnFfpNDOiCL+eWe3l0c9RZdjcK4qWNZ8HY3Y63Z4n7M2IgCZf+vMQPF
Mo07w+upMZDndK02Sr+/0bfk6j3UGqVWkfGs0y7iWN2Ans/xom/otOp1v/UBZDnZ
0uwLypK1UHYGXHrscQfZN45r206DWHHpbsvP9GTlBShri7VL6o0c7CRgWRKgi9cv
YRIll9dbIu+byNu1zOFBrFc3Jk771LUEkba7lkdYI2MYCSwpN70mL7ck2ROT7NRW
mWF92kAftHxormeQfTEuG6WUFYvG7tQ9p4xyHCdgY129bpyvUNuksi6gRozAIwD3
q1Fd4AKXZZJfxTgQguIbIOOLeGZtUTmZS8JRETo5Bk2oMxbEZJcg3zYHgI6P4huh
n3sBea5EofXIrboF+AElpD1tFyJ+sYRHm5NhPr8vWSlPSRoQmOv1iwz9Nlh8sJGL
Gt31/GCSFwL8CIRelfMC73Uwy7L8FUrwZFGtnqB+f/He9dB06YdEKmgJrDK/FTeS
2ZpyIub66V8eBKPRAQ+73jgAqI08n637l3eW+qk5W3OQ06HunhnuYqnS5TPaNiTG
x57KXx2UsTUZrTwF2pNWMnF8kfpYuy72qLEvjKTPXmlBfR8FBBtCPi2mkiqrup2s
WZ7C/O4INj2psP/7JeL+yol+MxM1ohmdsUp5tV3lfw4GhAjQkn/xkzfIJEOal0ue
OLiGobC+r5hpObK+1CaypCoKAT5FU2tzpwgmx9Wa4KhrvJWVh7dwL4o3zPMn7b/j
y7sjND3SuGmJpoRs4toczcIWRqiRSVQ0/1UKW57jDr06zvqK3uo6Bz0eelSga01L
bVRe2oObuqwz+tNsXSIH6Y//3rAVleiMopJnB9eWQWhAmpNEowaNxU58/M2mrMuW
mh/ZJ/0LP/xMGTs6NuTR9ehf61HDF9qojZqWIW0a+pKiWT7JtUGg6z+CFx4cc5zd
zw53H4WSFi7L2ITsO3IOzBz2Wil7D1j04vL+Mn5WieW5MiyFSM1MGpqenQJJncto
rgsp3O3UAEFsW7WOq7lhSRBA5yMF7Zha8FeijcRlex9tntF38pbtANJO5bMzdxbv
ZwzzSTFIFyaICTzbSyuuAeftmMTsx+R49hizULd0sJbAriDFjYmwFg4+ltjMkin2
LrTBODUdcyPO3qTrRp4DOJ5tOuHPr/vBB64AcQNMVkoVn6nkObVoDn5HGmwj7CQH
xLy8cbpjhYQLeUkAJdUHezLnPRV6POQ6+s5I6rDxdIg5AU9o1K1AkB8K1XeqqCFt
MTgFuBu2wnWtPKYsOn0FzeqpogE1XHjgTnifPY0fIkEpChB54m40gvn3wkDoMG/N
4oPAfpH73lZV/LZ3HCeJjvNtYLJlMk3dvLgHPyAWXWvUaZ55Syjb2Rf1u/2Hpgyz
emqn/3/gdiM/0DUQ6Cqh79zt19wg8E1aKiY2qTu3S1hBsCPEVKSDKjCxu7dInVoB
vVwrNKjXaXJTRKjx5qaELZ5r+BIvigTBrKAhopJOiaN7ZN9+dXSBkGSd5KCCk1n1
IhjvjeH6Pyc85vPNr6vFCNBkWjgWZ6RQ5Nwlb/gAmKW08T+6aBawvX5P/CTqZOof
v1f9rt7MGUbevAb4O6tjJBMHtOY6oan2I/hGPcNXcbNoJ7Yk2jQAHT5WlZGWdzO8
w2C1XSc29nY5BQJtmyGDuhHvb8eyHiRWgXoTyl1eyAxJ4xaN1ptzb10+TKd7UUsl
Qn1tKQ5LPta+8kzRANpKE+gq5v3Ljl48VL0EQauT5DAnjTGqdxrvrTgzoeEkJ2Fj
51ZvRs10WOP7YOnfd0fQD0cwyQ5m4Tmt5bUHeCqHGZv30EdlwsnmXCB5FmaPXidb
h9REfb2a47q4R2FW4N1GMVh0qCfPCos7wCMxPqF3xjAZjhe47jJB1uHDlBT0k5mS
Muim0KMm3qAeEiWApidF9HaojrXR/1n0uFPy+bZrJZLRGL/rKoItuQp9uzTJ7yUx
BycyBOMiJuMe/i0WuMvERdU10Ib4YxeQZ3hk39OvlKXUK0jBfK7foKBFk0eUpht/
gylAFekBQM4Hl1lPsw6AvlvQQXUSDidpUNwRdMX5lRtspa6Z9erVOCCSLlBB0q9b
ruJ+2t2qO2+P8uEz9TzuFOLMc1Vo7L/Bh+99hpLnNH3fLoYcEOIKmLf3mpwBAyLk
e1xFyBAzCdWmE+qqNAml1R+0apfnHp4A37m3oSZBPKPWy9Fob+AoY9yZOdEw3O2D
`protect END_PROTECTED
