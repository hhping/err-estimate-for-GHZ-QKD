`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uVQRpOxuZ5CX9JMHGiRKC6u79RlVzJHq5kBPce0WPvSiBfeN/zVtWJ/AEUrVnqE/
yijFjN/jMYj2e2i9Kz67+vREbbfUyvF80+B8Cc6Xq2Wpv6dEcDF/abnqWsNw/BO7
0Az5O+X5QtHAfOilrCZMUBNGGwojOtoHstfxEQT2gEOzaCYqf3sOfWAKusFKXQZ6
4/W4ABm8gk6Rli/7B03+oP4c/KONTcVFTEa82MzhEsjWqAp+YaQAVJPJ5P63HGq0
xyoNqZKYviFyORkNtLdOQ+QP8Qbr6CAyZNL9zTpFLIPvWz80XflL1ncTDWVxKI+O
0+gR4PF3bxkgzUxE93KIEzvcTcBK9+rI78VL3bFWMt90D6XP6/Rmhe0fnIGQ+giw
pIsyh/87UMISNezA8SeKJRVlUu+bo/wsLUZg+qHDBiDGWptqPtC/h1jZGpiaHR06
pBGIv0qUcW0XuLaWVpDZ1BJy2qQir2nzIMSCtpWwMWeqwxcwUtRltg8pR1/xhw/r
AyXJnnTsGYVUlswFHyfJK2uxNHw6CKA9g7DpyCeUMoMP60AonP19z6aeMOsNNFWp
PFyqBYhIZ92FjABuRZK5hDG/LG7hFycW8MAhSbjy0FQoi7AOR+qMsJ6ZxZ2JfYZ1
JrCMsqRuKeu7uk15ubjYY9VUg90YthWiVXX3k89t3Hi7q+9O5kwzwn3CtKZHFU9t
juCmlgGuWoZ+3TQCOQ/uIlivbEWcucIPOdDGCh/dsmkLYRdoBk6rwz4yrjTJ7kyD
AiJ4IjOX3m4LiAac+7FA9cRDzlltcIMiWSNLstFSBPjPXbwjYaT8JipZ1VolG7we
lwDjLLC2FzBTNKI0xzgdc8zoAkBMEUGE9t8GLLRQRIY7WHfO10TWpOgV/nI3zAgG
I4aVKbmYHZRM/juBlD/HPH08xdjHiYwyo40GuGSdrP95tGv8rwyIiM9x5PTIzY+4
y/t9/oBz9B8h+1SRwJyuNxcS++Q+ELr267UZ464pNuqFXVFhFRLbwQg14+Sqq1yn
hRM0THsu+7bjwi4Yh7T11iGKMno4Ecx9Cs9azLnrLIlCSwbM/G9qXPfmCYvFhK0F
KlWNhker9YBloedPC7ZylzLhqRm29tZkRocLxP9Lsvu3Mb9HoSH4iCe9dre70D0U
dgAI/Y/bV9l55hnOTiMgaqi+Pa3klEfQHZ5Fu7MRCHuSKlYie9FdgwDwG3h0UbUp
3P3u/SOFxAZw8qxDOKnsr/VLpEHtv4MfSL9IcHa3Uc3AzFIZBQMFj/z6oImMepHe
bUT+tdf7bwtwPp7XJ6BK4HdkwPZWVJyShB2eObyPh4rAu803nk8SBrIrvrQU0+U5
u4jN3b6hhGbIeTtdc7xpGIfUYssOdL/1mqP377IH8bAHB2gHfCVxp03Hg8W+ZgpG
6i78ny9wK8nB0wl3P+OivZ8zIEz8R+uIjgZGFrlkYM50EXAs675CJw3cH4ktnl4i
dyeFpwlTyEEmbAXBjBJC7WcymxKhvKHgpvHrITP8xH4lQJXJmLftAt//FS+BjsSb
WeyKn2tlMQigmf35+amPwbrqwMmFLlvs8RZQm8FpmtuYCZv3f7RJMk1a7AYFWiuD
XLlRP7xhrDNmrVu5WZMkNFlIetdXKMZZKrR75Qp4cg8WsiKuAc4+36mkCeOvJZy2
UDWEs7eZoAaYUD1vc5MqzZrt11Sm8U+MQEoCrZFBwelt0Gkgnfi6Kq9GbOeU8fAY
x8kCKcpq0QL+5wbFmezFSAJnWgYqzzN+cDOvtFYY2pBu2PEMdRY6tDjXjrIpt11x
IEVninzibAdbGr2H/Mb0udR3IUoP5cLudEhkMUbd78DDFJqWBajapyokQZNqHIGU
rgoxE73X2yjcvUhx4ytLJr2htNUCIiCjhAHXGLXDb0va6e0/EzbWkGDNPZo6ActF
cFQArDQa9SkjEp5CX7x/6O2xX28BYce3cRT9fGyQjDr7zqu4nkqOp5tEdnr6yqmK
/R8CKrE4b5Lf0jzETimNxDZWtCXkYejehaXicsrVQPJQ1WHHWyS0vvEs9zg/axMm
vhGMcouEc9banUxsCfptoYNCEAqNhfF5RqrPbNo85Y0RS5dejcZ6naV105/QCPB8
rxY/4rxas18Bd/S4Rf43vPc6HXorNOoWWp6RDXkqd/ALH2cWLv2VU7foIFlOdbGU
/MFbHqOSHfJEpgLueauZpGrFJAUDuA/Y3+SBEXoV1eY=
`protect END_PROTECTED
