`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nhsxZqy6UcDhbO0o6SkiGIJocg8z3vYK4rIlC6UPmvM1+prVF7EAlDQ9BtDEUr1N
N7toGVmdmGWsHySHIP/BDWfVsPHZz5eVZ6ZrgPWaEnoXaQsMwzSIGuJnekgR1/1g
s4fOvJMn6eN926Xm6LrWCUJbZmDC4Mw4g42PRUjh4bDJC0DVHitPyEjmkD/cd0S5
TItBj6ZwXc/y6Kl/aQ5UeNY1Y2l+t7LWk4WityW9wP3MyYrLKwjm3HQS3wDS9G7U
l/w//oTnufrC8kJCGs+EWA2hlQkioiDa1RaQ5aiuSi4A5VMHKXR/bEocj5ZVcxEE
BZJGBk5RygIJkyHfbvaziX5IbFvfRo2piNeo5FlePoWy1asOAtkGGJLcWHO/E++e
9cNZukOH9R6ViXiBFMYyQnvCKNHxiibqAnPQ2IYt3pn3UWhJ9jyqE1FfYh9UTKNQ
xzEoZDcewUaPCTXIoZ30BCZE/4aNLCbpIbO4Le3Bey2NnCyTYU9k6CP9zLab+JCp
wgrrTLBf1XKeVeUA/1ouYgo8/dnxwQZnNYTYpBwMd2HwrbdNDOEFZIo4KeY5gRYn
YdZzxoVOus16YH2LvQogaA6WgODNthEYBj0Nif8MyiF1i9CFdKZdk0IGBmBL2cvH
`protect END_PROTECTED
