`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkEtDauc7vkIJLYnznWAAF8QhHc2Wf6bvT8LswOpoNTVWhVDHwMkWwFdzwCtDPdB
ufL6g9bvXnaY3YUBnZvqvuIi+7XoHgV88U4ALDsSab5UFi4XodlzNwh47uu1QZf0
HDrGUoq44a95StvDne8ja4kaj4AEMsBp2f/bz62VXNejvBDBLG73BJkUsuXqZ/0Q
tnqsJPFg89QiLcC94ldlhL2HzoqdQ0fqMM7X9VjzwunK0Z6GOC/sP6euSkIfBqau
u8uvnW+n2Ctybwag9n3E0Dc6CyBTUU089KwEd836GcVgtS55r3DZl1KBj65NeIK8
EY9A9Jm9UoG4/4FYUTjmg1Cgxkh1ripfI0TXlZ0CmIQArQYOeAxOIjRo4bF3uCt/
bGo/cE506hI5Rq+rBNIGKknUuF6YVT4e0xQh/1PYAwQME6z1tV/8aSVX7y527Uen
6ftU5YBRbeXk93t0InnmYBcO8FF4/VUKPQ3jyxr5+LJm8zQnhdurM2CYrgXrygwj
GhQqTPPq3jZJjWT4Su6ECC/G7xop8awuR2ThlyJIi1eu+reNKcRLDO92+zn9Fbcw
GGLFKQg1kG+CSu2+8w1tP+hH6gAqp+xYIlr9mGuzo6q1XsKWLHqSUFmyTPiqmXag
7Low6oWHXGC8YqDRz0KQrTx9ANdJxR5vbqNNmYJ0BLTbc7Xu3SePeda77WanddZ+
3dCyCjlMQkvWkELfoFTctw==
`protect END_PROTECTED
