`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYN8vAbqgblAI/+3FaiQeJUSImvl4FuvQ5ipLWte6nxn7dG0hs4u1GFL2bIuwI4C
st3hgJV98gNujamaH0bu/OqMPg7RKq7028f6Olmw5f8UBhWxx/vbvGMXnecekRa9
EG+LnABh/z8uiI0Y4wEI7eu6/ymDNKkWmbBsMW3ymcaNwqL5PP+zRymzu4f3nySC
o9R9ZJY2t3N/H8F2pAoTMVbHyJp4suYUq17sdP01oJ3NMHPS8GvnrgQqYs6HtnZc
fO2oTKsWCr0aMc8EsmYXsDnuGL1jNjSfQHGwzHX9O9TEFGO1ii14NCqmS49+muI7
If708RM8bG3kZ6EosVc/9Q==
`protect END_PROTECTED
