`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHXSFTzyCmV21avRXC5AY+v+xWcvv0QxiTjk7jgOeME/iZhqSZRMPoYyUzgEue8I
YgmBetJ56GxaDo8x73yggxNFCkt5P145RKazVb2Vd0Nxap4VCPz7rd4JYr3di0Cy
lFXCPXsp9Ich4HpnZ7seaQg24Y0T4/LjvVN129LEstWMjpcjT0aCVg5kWV5Nin0l
c8EQn7+4qZv3TJMyuafRFPz9dpTRcIlv0mWSR7bz9i/KTy9xSZF5KbxH7YMzRidz
uqo809cXeK9fZOK+P54cUmy22RUQJLW/CnX15lPqlleMLVytlG3M5bqEeSU6Sbym
tCgI3eUlRAAt/rhrcWvde+zhmqg3idN4Nuzx4zGU4Cf/jfPuwo6KYPHrjj2lcWdl
92xGIrutGUd0L+KC4wIBYpFQW3hGdqEvJ5q3he9FjmgrCLtAcmHYroQQ+5636Pfq
KnmGRXFEWfSi+uusG65cWLKQJmkbDNMoz/OKEccYy87kocsI/8kEP+EjOJeVxiu5
TBiienG4kb/rKH2bIHtr3eAPqdeiutYhNi/riUtNUfgdu6yR9T6VUhottybvuBRI
2jUdvLjVOdEPwcIavORgu6SLdi7F9swTy7R+xu+3YzsmKCy+HSFGaDyYMZbml9fg
gHGCUvDx5kPeveG8laAmMlYivnIZh+sHj225gfPVbDE6d20NcXhjlV9hnP3U9Tww
3W5qE3Hh4Pnd19LS3eJRdNjILoKe01n+aD+UjLVGAEjGIf5fuvmp+OmH0NJO6nY6
4bSm440ekaD0iEyfTcT/+eC4XsbahujYgOBqX1YaXSbKKqYwDeK3woy2Ya8WJ+qa
YfpJ3waE/Vm2iuBD8qahWTrVTxfn2z1yCLhhmdefQ6sv+iOYbZnU9AVhttJv1Gf1
hcIje5pBFNHTczNnQEv93aL7oK+bsWiQWraImx98k63Oi1dSjYh+tsM4ANJsLwKy
aoFnTC+lsVJLjzd3Ul/CENaSqkf9jk2/3vlL4QAS94dQTQSWndM/96XnULfaepV3
/h6i5onTFCHBIUi55Q/wgv/w+29UG4k3rXp0VHjEbYvfujgkIpqzgQMmiatjBZmN
Mj1DZUqZEKNDtcpD5X0851LLAQzg7dV1PCn4JSVAWcR1FWosCkZM+yvz58TZg2f1
iWxNFuZ9RN7SBkQiIffBryik1gl59xNpq0JoSdd6vnhrAdaynqKztYMxSK++YenU
Myez5KaDARgg+wzTPW4vYGB6H93tCs08zeXf07whT7R+FwmiSHM4Ptup+jxjQlyG
KjF6ghCgj4OvEUylYIuktYU01+VPH/gBe0exw+xdmOJ6oQoTz4NkZWj94AEPLGDR
R98Rn+mtHqcNf1sCmJ88zX27AyUJQYbFtK9oQMlYcUFO74VgBZ1l6i5HjaTj4LhX
yBw0UdT42aAuf/oQQbisELNqR48ol5Lyu10Rc4fDN7ibCt1UwF9OvED5K+50rJ1v
TQrD6t9W9ISrBOM3NsQz1jXa+hmOEIF+IiE4foM/B/Kcnu13XScDgRXK12s77zj6
1Y0dM4QvILlM+qJMlx1QPZAbuibwfkeY0vZyq9tuf6/lqCQbnpipbd2XDaAyILtV
+lQLuKDMx4kSdBqEPPQrkLbL8Vy+FFOErKCpayScnP8X9UXqNJ6lst/51eQv2x7v
xrG4NZtxoFll8X/JtPNeAXS1Ld794vVBkcNITYEBmh9ska7HqkxbpL1OtpS/RyG3
HRJoHjXo2fw2sj2IOeWI9kjxxPG0mXe0UAayGzobRZ0i9OuOu+Ab8Wt4j/sXnpOx
bFyHxtqDgZn175IxbIfjumuyx8vInjk7pl9U23fVVnNcaag2793e3CRfVc+n1V/l
F0u2oPlWggVvwWg4nwbd90fQZ+chv3AEIjo3tr7Y1t7+kgoAoLwnuZ6Kwlgodr+B
lZIVcMF21bDktkmX70BiKtTZRHgK27VCVWHU0Y1R8IWXMhKaptPQ+DGlBr4gJsjV
pg52R5aguN6ibhfi1G1lLjO1m0A5/VdNH8hnhv0HlBO54MKFrce/15rDZ4gg+Jsk
18Rk0OUaF5XXYgTZqgktDv0dRELNcCdEQKFzwUTRy0FQti5BlAqZ9IvISnULJxRK
Kvs5sII9cw3MKFSH3PQn4oLiy6EV63L7CJj70mAxGEN5RwhjM/s25sEc05cJTP+t
FDPhh2eJLJUiRg9Ye2/fGV98+me1wYvw1JDcPbM2omHOejUGHuXaFTI9uoC1AJ4X
uO7Rv8Yy1yzgYvQELiNZNA0Z7NJCSIQmIrSzK7d7hNU=
`protect END_PROTECTED
