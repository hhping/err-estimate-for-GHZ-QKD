`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6MDTESiwo3oEMsk/2k6vn7u3NhJaaBTKVOECgy++nbpQNmnF9JvEyFSUJJe8d8G
DluW8HDbRnjB3UtAXwtmaSzVul3If1wK/oGkVG4ihRQJSHY/z4BwoEkmgeTp1PuC
kM4/kXhmWIqoSfJszjH35XpvBQ5gYkS6xv3RaKZ9nnA/RdEPymrMS/WRCRKXxGUe
fnEH942rSejo8tJBYG2QrTqKTSQWtxTdGGz7yJWFnJ9odhbGxVeEwj4vMpQcTle/
xP67glFtdAuRURklA2/6bN84ZitJTABcufLq9AJIkBzLnN5wtqSsm9ebz+k+RG62
UT/SI24ywJeI8TjKDCl0evDzHuZtdPuFuG1EhlopU5VlTwm2sH8ceQPEBv0RGUz4
xHh6PzqsFVdP0Mt/uY6sXljbBQbx+wM0uUtzuq16JgCSMurd0zAbV02pAHxDIj1d
THQY0jPS3gXVF/VaUkqFAnmrT8d9KaZYW/bLGbsldjpZh560jgaVquDhEDC7FhMo
Be3DSDBqHxDux3rGllclYe5KSkzMPwLAzbl5TIiweKBF7IBrJBDL75QFCwjtgO6q
D4U/X4ak1hfWwEuDW8rp+rlwIkVsfA8p8PalfQCYMXjPY7fG//HbFUtojMol57Y6
0a0e/SKK3VJ0OcwJNMwkJLKIiUB7LuhRhDBTE7aqWRh6n0RnW15AYrPQmaWx4ArW
QsoM4WPTyOhvDFj0F1sEz73j8HQENaOJAFWshz55GXJ8BatjKSuV/blWmwLN6VYQ
PLUiJsUe4J2NXEz2t5HBPGLXOFP4aWd+EOcJWCwWa0/KnB2m6xvGZTV8HFbwfCUW
vhCK2Xbig3esqLvy44OZfGmakHid1Ia4zKsSvPQJxe/cDxXkn5tdzD/eT54O9P0X
5x4mp7F100yqRt/8r/93bYtXcXYxQXPXlaNTYmFD9IZAW14BGKb1EDTbiMl+bb9G
7uv40wZIzjqHPS6ePne/YLW/jOWp7zM8GYfahkQc4tTsl+rOhPI6YDuVM+/ymHgJ
hmaF4xhUPiIjXbFGF49VBBV2uRWlAAz9QMnl/ldu+aqqQ69sTFKu2BeFbTJpibu8
EpAWIlTyeSuG64KSeQ9nIePcWAYBTv+HblSFsJ3yQ9wXrwYvTBR2+b1fOu4HrO92
Axs9vr+NCCnq7r1mzVqEon4gje4oTbJzurjZk2xHeeABuN6rRkgrhxe1SAzk/Q4o
UUUAd6GjTipDXRs3jcUxXIkW2glrTYJ9WGBuSZMMHDzTrK+o0M3u2EQ4CVqFlyrZ
smMH6FIjabj8DTTj+xBCTLvWjDwHHomfdQlFxaoU9bujGeBNYou7o6KzLBoNZPvW
MiODeA5zT1aD/yfgAHXsjftg/TXikEiSXZa0jVwmehEZISAkXwD4X8ra/M3C44Qh
GkIqxr1r4a5mJp0pJksIIu/glZS7ROxasHfk49+/ql8pR9PtEXqB+q32ZH3yu9O8
0VC7qdLWxxSaX5O9jI4JExy9kaW+9r/if/d+dAsvd4qehL0dfHBOlLZldwId6P1P
V58g+d5F2MezsXOgqSFfIZHPCfWMpM/Waj0HIJTVWZwdfBMrNHlPAALD7Wvz4egq
Dj4WUCf0EwcIr0F1QCkPHnCjdou5Ckwidyp7Ic7x/ju+/AW3Zq/V+CKCwwGYygXW
glKKrT9NzgBTmFK86mG+f66VKMSCyd+lX3YBZpF9NArmMvkIWyQGGGChY2u+pt5M
AU5OmS1osVRiPerX1Bv1J695Tjkrc9Fsm/5j7yzj3ddssSJ1FtixgZqcY/c3OuAh
s4nsqI43ahaVV2IDYpTFQ61eEgoXYRkbUev/sYC/s0ooTahD91RvK1F1Wsdhl73M
4Icg8EjKAg9Hef+aG9gOeAmyWQpjUvPFZ9D+v6VM+zt7Mgx8nWae0b8mBflrBMfE
WyCUH8M9ohGYzRcIrQdD5aHNouDQucfObk8Kre/6ilTIipjhTlR3XMOfCcDrgpG3
5x6B4M13IPaTqXRol5vw52ICF85zWS2LhOiYlIvT7I3rX2WCCi8GIiZDtkaafdYa
LYjxU70UZ0UVtikQzA0mjGUfEUm3NdtaA9GjJwFdfp5GPJRs1Yh0X+k9kejH6MOj
+xHc4N/vBo3XVeLr4KUhuAunqViSgSu6PtCl7FK96GdsUqZ2uO6AQsjPO/Q2Ym/t
g7sNZfuO46Bbv4ozy/S6FnOVhizC40uThgVj8QfUU06s39iibN+AEWemeHNK8phE
JZzWWrYjAK29EjVB4JJL/louj1DsnFEHyoRJ1MqdYN5ZanXCBo+b8t2R7dcO8hmi
qLBSA6JCWbjsEKcH0gecGHkwUsId0sZm0vErShyl7RgJ5ay62q+PWAtN89BDSTKY
ymlyQ9xuhuWD32s6dZOVUcW91EOONcrY2YsRlDDzZCoB/JLtfMUftvZrCEjbm7bv
ZUSFHMhtqQiCO007MN19wR1rriZ6GP4/EZ7Bmjk05GrXV2+XaicP+K1T3oluXsi3
1IQn7s8IalgsE6xRMJIgoK9dyf94HWZ3pDiGSbTK/vcDpV4mHFW1AjklTGrxReBT
UmV/WgxbOHhLhIGEBmEpKdLIsZJRi/377fGkl9XF/nYJ3jpXfSlNkWf2gzoBLsMp
F1jL/hpCoGy1WX9bhr+tPnjzB3xhTqjsii4ar/q0tcomsfFcNDnPt533yX7FNPMi
FMQEOaEqm02T6ep7V9DxWpQYdoBWodSRrttHl7yVP1jn9cYOBI4gl2pQfqpds0lm
DR5QAn//gRJ2JXFXmDgm9zK5dDSsWwnQ32HuHr+E0pU9hJvI4YQYuBdO7THHs0qs
fpibUo59MrVzvZTtZtyBehtmh1i9hNXg6vsd0XLMtjEg9rdfuAcrqQmBnm2o2TrB
G1oi1MAVtEkgOhEP91Xoskkbf1GmrrUg3D4u470ZeVx7RgSQLxrxLS9t/sJc3bos
gjSh+msoAun0F2sCvdQbIlvwmhxY1QmO+DxR9F6yCEmeUMARoVZbkaOlbE49KR4s
yOiGLOV9RYKIsxiVXq0b5+MA62wWmDBmjcBDgcPVjWV7zmIkVp7Yp/l07ON9kMKJ
+jxrmR5wj3NOBjHWp65lZ78O1XrrCQn5Uz7ixBEl2MKskKKdGOB3FFtWOFjGycCl
Lqasg+shAcwOpmRaWzNbWJ76JboBQmCuy6n0AWcdF4xlZv5foFMKyDJLljjU6wPB
RxT1z5xYxCKnwPZhTWJShzkAQXYB+0vC8maAzYo9N+xuQjtTZ6lONWX8ejXg78qR
K2sVummVXnVI9OZZMmLAFFKHvHE1JZAeeFFs99LWMWY/UKdTbqlMW0g+e2Yh5mIW
6hdlqsCtMTvgcyMaEjCshRce6QEyQzn7Ac3Xb+ZMhywdcoAqrUFZw3Y5TSIDeLGy
vkuZ856qb/5ZWYwqsJseY4fPmfEX7OsETUGL2st9Zp2tolYNbwj/FS9C1MpQC8Ek
lHsfQ6M1Q9Vxx2FAOD4sZ7LoniPIFxBy21MPhzvPxO4BHh/TIGFihj1Ssq7o1zL+
L153HJhf2GWh08k67XbWNwdCiFjtajkjGUflvdQrKOxj9YHsdCmptVi0MhHxEX+I
OADgQrATz/hQZAGiPR6ITHAxCcGbF/eEoVBw1VOWmDTwnD5nWIRuOq1MHhqGYk++
WSTCSgi+hjjmELVr16LDdd+DU/mj6c52q8YiO0NnHI3ZV4B1zfivV6ut4CbHu88l
pTzyGhI47Cz6KvJNnyC1ad6QkGPNmlKhBCU2ze7hfcvomVcz+2urWNHkNOxmdZB4
b+/KQrOdzWoAwdpWTeuU3RrVdLCxn8jAOOg+Cl2qg8PJTBp5JSAywNT3gm3iwOZT
yTItP3Ke3DYORtyGFkSTXOLjaNCzKuPu9lL8UGNslNG4N1QA5hfZqKHr4UVHG0gc
f1QVACuN5C9N7N8F2ZhlFpUttHPunEE8B8kqiE//HOOVskwZETPh/iG9nZydHJn+
6TpdeeADvuuiUfzBy0CmhzL18C2aiIRlVxP0gZ/KFJBqoq4G5H/r+v+oOfLo5N9e
9VE2diK8VfJYpujQv6u/5/YywJ/SGCMTtjvpiJ9UGFKAMtHeGoJ2I8Z31xyiaJgP
MPUUZ1n8nNaahtidK/m+SCpYNRYz558jNhGroRTIY7Vy6nJkqayODrAbCJ6LEFAM
YpmEZDrfUn8A3WGIsDzzxSnQ3MvGSXdniKtngacEhDEpiK8bqel21ynGPPkxmo8P
MlM7j7wjxuwCZWGDz8aIIKxGs9WG6jN8GsxbnFmUIDvQSPGPddUxEOfOckzm3igZ
q6Av4T1rx83RxcLUGe63wza04Lr6z8Rbr4gYGmqRoqNXxA1/6xfiCdJgn7Oj4FzV
mI/0GrzMwGDR9qnAq67YAK2sOF+mogLf/ttWwSAsBg4Fc9h5nAvQcpclm72tjfem
a5Whb4nNlkEiereaE8eXXfZTu8NCo7dZat37nZeHhuvRjy9ZhIrz2u1uC0GXCMvZ
YfsFlL3uTpLFuKBnIBTJ354A12wZiPvWsCLaEGDK7m9r3HuoJdjxG2I/PfYTVjF/
LL6NU2cGTZvaJGQ8HH1DUmGToe956pxByoLwl6g9wPyAek2DfLkGD+8pbYEu2LUK
bITqlrTw/8zJQScfyoV27qFSqVyzr4UlxFqvroxh8KDFkHJvnsnl1bSC2yRYe3KF
P2Hr0XuOc+/KuyzcbE7koOMhDgaXyrgX+Z6YzgVIoGuk6cy9zY2JMhg2vACMaeBs
TBuMZZXd1Q3kcQhKACpDqeluftuKG5IMynhk8VmN2rZHf0zXR6Z5r6mHaaB6qAH+
lnLvKK7N32PMDeUpHdolYaCJNQr9VhgkiW8xKqwttASIy9QU4Xi6yBjS9x0wVuS7
cbbY+RAdnehQMJjhu1VPKXYJHt/9Xnn5cqyyQwkSM6/i93VELuPFvZtpAg4oBOoW
k+NyzzAUF15bnNsN+8AOjyEFEtBfvARRwSyTM3VOpLCcfCFBMJ6EvcVqeNeFPTol
Jj+xOSAbaZhePOwnC7frD+6T0W5PLxMvKBI1nanlSLIB93GvCW34Ak5ovSKTttE0
zQnvff9M2qefrjgO/4dpuT/8fOT4FhjCjks10ktdCaFeeGI0nDlJ3b/uJtwWbNZ0
Fn4buNtbcu8faHYPZligap4P97HaKabOrD6zvw2Vr988r3Dg+M9PvMhL1AGAW3l1
JJw9Xypd94CnD5f9f5Fpc9Wl9h7bKR+GOqRWI6NgN7f79oGHYb7yrr3oSM4V1aSs
nDfnMfGWEkDAno+OLtEi7ZvPIDOqnsOS8y245g5XwOu4Ipej5QgL+mbaH397qmGC
MvU0/HuoS+odnmXhuTc431pfcesyfGoT2EhihTDzGHQWn9yCspAYPMkIwqmQLp/N
UYWNoGkyq7Yi6S4ACq3hQwE+P03Sm67eWOMPODjCLiK9B+jlwAB4XmM3YONeOSzB
r08NlILe9S7slwaBroyLHuydRkvI21DDCSuTRIDG5YKohozt0vzxWWahtoSTEVo6
Nf9Uwr4da4MRCKoOZDgocOKgmBCmEgVsIwGhtySfcv4JzmQ5nDwtTsdSVVokkbTd
cUtG/FSE+MoV9m/D9siO23ZnZalBukiX3Vz3L2BMJWZe1XLT84Rhfs+p5XKdaaz8
Huet0eui3Y8iehXahqwnGeg/IJb8XyE9PvcRcw23gnni4KZwPUwXUYgtobbyTgWf
Mn2fnrSMu3LSx7TOmv5Wl8q+lkMwOb1RP8ySEUDQdlc0OpAqtPACFqaIbziHFpfd
WiWagIPJqDZfp/kLme9Oa699vW272lSqW/6CFj3NSYFOOIhnfDxkF56KsmYSAqGq
ye4yQDI2pFfS/FsHHsjrjXPK0FN9StaGNaiqIPKUX1etsSQW4Fq0cYR26oYXtjvJ
W8lwyJXNVJgWAcQwSxAmk0CYjxwFRHYkW+LjtaJhzjQLjOElF5oyw7JvWsHWcTBh
Ak0MylPzS1pVg1yJsEXDAosP3EbcQ50jqNxshca/vFrLKdcosfZVrVXP8Xr1MaEv
yvpCQ3zgUIUY4+554kvLelDsJenVZzIKTSA2mryXhBBazHOm7S3jBW6a2BAFFtGN
wCf9yKYVBgQ+AtAd49MYg+jJ/VHpam6QehflDkZZHDuNLypwO3eEOj49nM1xcBNI
SuJUZfL/w23Vf2gWHRsehTU6qWCezX/X9wKgPN/trt4LmgePQL0cps5mKA0U+49G
kDpzBZfd/IYOF4pRWYk2lARb26ftmXVATDsHzMKy4zmpbmcwkJK9CDfRrSqktl36
PczrA3tBq69ywpGorbDBJBPKrhQkkcKPnq/2gZxmSPJNWhX62xk1Z8CS5G/KGNPz
oeJ+USU8GNUbwh3f0qONuj3T6oWnRrEs6AdUI+31gQHWjHf4un+4rgsMxnbaIplK
dyEfZA2voVaPgRimlFNQSDwkJ8ly1BoeRwWyPk+SMlTEptHEbH63JzGEO9Vc58KC
ZD3X4q41DkuHTFpYVXte9RkCJ6TX5xgec1cuRlhf1aeFH68A/HDCehVtfCzrzxD8
dnr+R+c7040dYXP9SzXAmZHs3RMaieVfX00hnvB/uUfGgqadcpQ9Vyj79yktH+ik
Cqe593OVZ+b1iApE6nkPn3GIbRdGWL3wnt4y5YP5cPMDUwijGCgH7Lrgb7fXlOg9
PtU4Awu36uKJpJWXPICx0Eu/x0H+YYuaBBweBxpmYOZBEs/ADfwxBhIEcBqAQXO6
MuPT1kU7bgN2vZ2QIKYJWMWQj9EzP2NVe6604gJKrTcxPQP1AnCYI/VBjR/BF67t
B1iSTgn91bEf0DY4yiCVEohyaOE1KmR9JeSJz7O0zr9s3iPRgwbVkhBkpY8uljX0
A+wMhbVkcK7xMp4ka/CRZvdtuoXpsUXskpQJ0hmDgvOQqc8JyeVzVzf+sVgDkbG9
N0Ah+r9jiZD5roqmhZdX28K3KkPU9uRhvQmaVQnBe1OmhGuByRyy35wRPTnQtYlz
rqQD+hg9BVKLCJRI/xEScobIMSm1tVnwrhxbwvNbLfxZUr3hSz431324tThRKHjd
vrXziQtmF/O/Rx5f5GINP3xOGU+U28b0aY95TXa4NbXVEr6u/1/glKhV1mfqrJzQ
vNeyYDB2SHPfNfd/pTLkLf6t2+ICcoHdvAlhETxpE7bmhI0EpD1mE0sH2yGtLgU5
Ibyj5qSFWtyUUm0dv94iHYGnxoWBbxJR1IAlNSL9lx6R0F0h2l75uJgT0c4fuNx2
CqJy/ufr333Wf7PFuX7dV7mObJZvloLqbvrDcNMaUso0FyabY3mui6dPnriaw/l9
P/90oilgCwaLHITfOv/+bin3e5Y/qfGxRRfPBkRCrxQ=
`protect END_PROTECTED
