`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiPK0dvzizz3Zcm9Mx3a1nvXH8fzeRkzjfh5tXqenWIPqMRdfrK1JpRCxgustZK6
x9PrOcrEOHmbdveGBGtdKDnXsujTbHGOC6kp/BAMY9OzJVCQG7V3niZK5Fw/bymB
qCtPtRfOH0oak91FzbXzMyNt66ReUMwTcEkx10qqzCP73ZiACmp95hIaoEbhCutu
2sEWdJGB73k3BWKgqyAt4ody8mG2J9Q4Kuk+7q/9kJkAI6LoLMT8biqm/bHJufVk
jOghHmd6hkNw2H9CjNw5hTKjUoNBhJBFMPAjUULdUyLkt8jCn2omSj+/TcOQv0Ay
BOELpA4Qy5hSlYMNznz+FSw95JT7KUcBiYCLdUQSa4g3lXFCcpQwM2ZQ8VdFzmJ9
/4FLHN2uP+/xAUUQmzkFbqfhzgEj6+gq4J2XZODgaCmOazuqn7URmy/5CpAa7bS0
usLiG49sS95CzU5RXYXmECKb1wJKvYYoVFF6r4n+aBX/nij9XOXLixdgKZtM1fHb
93ClEdhU66V5MpY32zfWpd8x6Or5Xe7pUqcmrmcd+q6zJDZmarL2iJYqlh1Wnrlx
C3mchkf4+OSfxBZn7/u/8v3HZjJtpSUM5mEVbu3Teu3lK0x2fJTPxcYDwoon+Fb1
lSMR3mcHsk+PKhADb5AsXPAFobaBuwhHVWzN6CGhVOwrpXpFhPwo+cBiHygdBMTm
vhoiSwtk3ItUX841WiahpVtYCLJ4rvyij4SkjV4uu7xz7v8ZxRFYvvH+H0h1+q50
ayOPJLIC9lr5SRVKHhRJX8THbkqHiYuJfVLI4sP6BTy0oj5nElKdGxG2sO7Q63PW
SOt60vRbpo20eY5HXMfBo1m82GAOT6/0fuMgO6BxdZnuz99JXv281+wgKrnmjQaT
C58UGyJQsKCaKj1vQv/j0VCsufYLJkTm4RfjTc8/Hm4TOzsnnGrwW/dRZKxPNPDj
wJMrYxCBkgZOpyCi4HzBnzrjk+bYpgrr3iicyIjRrSSRy0JdiVLDZGRkdpPfKt4m
I64Yllxoc9EwkYfwF6Tn6Pc/Zx2J9g5GcrCzt3OXGljJu9K6FGD7ISnPLWj3Z8hY
IJc9ii8Pvs+o2I0A50ZgTrC0Dwy1QsmqbOkfiEjNA2AdAZLE1GHDoKOo2fOknEUZ
hiNyOw6u/UHX7JVtp+xXs0f3qTnzq6r3KqAwwc99pach2fZQ2SN294XPsa087Xuf
m+Elkt1/AHouOAMeJQ93dAYMw7jBUv//9InE0E5o+a+sp3ffi2vanYJUHr7Hc6Gu
gbRtWhTte4xMo5lrCXtp60TmBvOBg74PEsLWPKHJbZw8qUMA76vG+8a92dsAdc5x
YcOKGl6sQzIxoIobBhdxL4SWtcYvWxHIfXpCFFrM/yPWTTy0ggF3eBR7wjd4f58Z
MXj0LWTt9h5Wi1hsfL2wZq3JvSPMOz/Dj5+hzRtW0ADrwpXDik1Q3ZBVJOIx3d/u
r/pghUzM+/9r7dqyCF0ktUcUhhLJZD7DdPbjlVIzna3kWEgpWs4xGaDuit05o7a1
o6lX9XgjziWT9pgqmh8/auhCpJ7O3NYyauXqnnlFm+5qayFASz8EgxNpXe/eWIsE
ogB/8D6jvxBj5AQubghtN9QVI6griU0SbWxGprlAbmZa4Oqp/dcveQ/+zQMaxYCd
LV4ndAgFerLohhlQdCM8SSFTty1G5LtVyg03pRlnEE3vF50cqx9//JJ0uHLfdZgT
A+nIhloe9fX+4NCkdPjPbT76ZL+UX4869SmRunC2YetXXcnFKyzcOzqlTWfmHznk
amp8Tlz3J6ewXy7E0D+3xj95lXuAvgdGGyZAmYq9DeDzQeHrm264xiA9XCOeCP/A
xEdWLQ0k6gRJwsvJ4RKc2z21hrun0nU8TTJQNCcvGepBccCfvrEvdsWko9JDwnPu
ffQzEW3LeSh0UmhmIPx8AXboEqz22ozQds7U+3FZjN4KEIOylk/Z+AmIA9b1ThRW
7Qp8SvvaCNSzMcZs67tnef32c9Z2F3m//USpsYbERD7IKi1rnoXnOXiKpqaIAQvl
9iTRtXL++Vkvd8js/Uf2H1kx27AA+5WVk8josbjE9UqNdgaFlvzR+lkePs6PcprE
er3NGjl1C/STPvIq6pAbDpyXZFgfwCydLKJ+WVjQ9EZCaBT97ov1kglp9XjT8uhQ
qKKOkqRkcOUjJR2mHhLJGGbpnjeGkpnm84u7Uhp+Ps9VW6PQ/x5hD6/EPpaIH1BL
u/LZHdWL+/0/BpGzg/Sefqg5LA6yQM+JD0oXPQhtsV6yd1J78U3FdDfenX5AEUxt
8uiYI0V+8nMpQoXX+CNKqfF/Mp+FF7fgvN6INaUMwmNGUBYk/SXCVgoHMXKXigHh
j33DFWupUna2cx30c+wy4aYrSWDQ4gAE1uP3op4Zycz68XNnaVxPg+Y3CUdo3Mnw
+38v+hPmwoWmoaWSXOKyLyPDekAmQ3pLjLTyxs30anc9kSLcgeDcIlB5PfdMFpvZ
Xn5vlBs8CctFG3cKjG5Qk2BeU/AmQMaHnnmrqkdjU0alLMaoI1dOcfe7tHESquEb
MQgLngKRg3CxQNq0pxCzcayNNRWVZ4AomIPlZ9LaxrCNqI8LiJs3zD1iMXjws0ey
8K6hziYg4VWltWpqoMDgLhkkW8+aDAdDWt+F8/qQwbbYV5vXFuMXQM3QqiQp7Cu0
dVeAz5y82AlMYlPTJ8/qtJGAq/Nx/TFkvRLAaImeS5Sls8mLMQv7AkuPtP5UwaIV
yunAjXdr/bTJWFg4daf3cIbJLKKNgsz2zL1X8uurGKhMbhLeC3kj2+W/MVIqLZb/
TTbRAgndn9jMX13959riODdmER0eIQMaxzZ4tjMyAbN6lDjSnZ3DMk5KzvfV86Gi
18YpvEVs9uzwUPkW5SofcYGcXwveu+wR6xq5OUJa3txQrkvlLWbioI8YfavQvTJR
Z2OZ9JrndUHFPJcoUZkD6+U8SaNk2cnT4foAcUnqP80PGuvOZhETX2xhivoG1SAP
q6GqNj6hKjtiktJ4SWDQ6ir3L3Klk44x5clhz4SXH18Gp57ggbXoSHUzUUQ1gn5y
M27MTJi41NKZWhK7Hsph4aS8aM7Q4OLtKWDlYOn2NXOjZoySlaFUFkTWiwkzV16U
muL2QVtQXnfQFTAa+xCLP9gPVyDnm+/QWmRDigUAgcTvyNnipLhjHa2kCIMApNNV
fNNY4sh28rYYXKyP+1nvhR0rFdTUbSA0vndBLKOXLbHXdlb8ywRXn17qP35xj9YE
4DTyFPxvwPbPdT4x9eVN4QX0hkXhmDnq9AzIQ982djz7VoDJIGKEIDSKpDvLPa21
IZNaIYVn3IGvrmD2hVDCAmYuyPA3A73mol1pJlWPvfQ0G4cR0khaIaDpdaHQI7iI
idyYbI/iRXavAuQbR0jDMHZHpAoljqXpftb13ruVXw6ubA/M2gx7ANOLaDrxylVl
weCdGX/yf9oeyA/d3Y0Y8XzLjTWxNt5fdkmBjlg84CWq1a6gB7JO5RQB0E1r9wJf
gWfvkHFQzRPUerafhUl34fRk2o3xFArd/lY6UfjRTyOR4sSSvCQ7prwWnkvhW/dX
dQhCQLz2j/2dEvWqWD+i7CViDABhBUHWaZQktXTXXStnmhc39lqurEKhG1NaoSbD
krRcZcF+qvjH0+/Q1JaBySgdgJzpbzpESyqOS4Ffyze9MPAL2P4tR91P4KQELhBG
/9NCEUpTau7KT19tMkAicFuqdgRkAq7OD8RtS2kUdl50r4zaM8XhTeIi4cA7Gwv5
aIewX43uxn3DXoTQJH2kOBcKonxvP8J15XPDrBoYXDGMy4oicYQ3w4YAxgKFiMzs
f3FZFeTNFSJdctJiSgKreVfUxFq4Oi6SkUkDyXTRraX1uKFz0IgiPcbxCqJiqY7v
n1lHcM7NfWR1SWAVpxPiNJzGByv/ps9yV4bEF2hDUziR8Is26p9oAXJSWn+BxkKN
hSOH8F6bx37Usumvr/jCPIACtJ8TfDWApTmF+dG63vw/ucLA06yW4E44UFcmRv1K
uYBSQ8grK/O3hvpGVBxCT45IDFHUlIaKQExmoMpRJ0xp38nS/RHTkHPdt8LeetV/
XX1h1vxoRrkExkRTaYP8xnq+Urcbu1ZizClqLGO9jeAzwvMjYZdguld6XzJBfgp4
Uk7BNW8jSr2Z8l4++a6n2STb0M3Xzgu0avQu5KgX2jRr86HauJyMetu2//SQCrd8
CP1AE7YOKY3aaEb5VKrhijnfsXYcMFOA2/G9MscBCKc/ghYCCOmUIm/Gu6qrV5J2
02Lw9BQsml2K/qGrNM11QVF3x4CjFvIF62r8lmnOmdIgC9uNi/GvGR8GZCqcuixj
+LPEWWL8Hgwh9aNJg/GQ1v4494hk7SRupy4DokZVhzAawMZcQFSObuwAoPJ4pGcZ
EGUYTZYGywC7JGizrjwrpZf24VwetxO6R+0MXGW1qMH3hgSwbx5DgvJOS79+uMFD
2j7D7Zr01n/A301DWbuhKqN5y9/8hR8HKYzxCKxidKt4u2TcSWeWx2PipGbKbX6s
cQFvROjBqHB/0k6ByUFSJ3q4Kp5qnF6AIDkKwQEXXlTCivoJlNpu4iD2biD9jkdC
l9wEIB6IuvI3+ODGY+u3Nhn/3wLBJW/uDoF8FebxymU1XMUAf8kOHxk/AjA/OhBY
z/n8tRA1KyUf2dcmS3oCQ+TkW3WTX3F6x6o2ltChMA9qO9L/jNvBhSjUqjOXaC92
I8qmvvQpEWYeRsjxZc5yLLL/13aVWm0O6V3/e2462nWK/GV6+qFC2EJkP6s1iP3x
1BwIVXUhJxx4xTejc0tBb7r+vAgNqVBmEHnULrPlyyR0MKi2O+A6c+i8YHbv1msF
vOPVsQvvZCgbTEKRbiSHEsAMeiXGTKbkbnlGpkO0vqswmJPaXFPgqRiuh6wuRuo1
K7op532I897sLZYPNzrEo3seeTxRIeQ5DhMhhXlcHssW61Fbx1+9gELHkZJ533uH
Re8B5rTtaps2krRrLdMDJ1KS7JRScgQ9ltCG5AxsevaQlUvmqiBCTKTp7r/4MvAP
EiDzS22Rvduu+TARNu1DiSQd+x0O9pzuFqNM2pGY6jlC1wdY/lbWdYoxNgTPaq/b
VZ1Yy40DW25v0rrii7z6CGc9Bc9PdgQrHGFwZV4CpFD43tv0P0xfYeyyTqegM9Si
IPLuXkVA59pX6lQTC9GXAMmy3DnRTXSD9BVq8WRs6AQZcfCtcsgKxOC+72OoxFtY
8TVw2JSd7BdudAz2Sz+Z70F1wSbDj4rhqZ+CLpDTtFuY0ms5yy3Qby3Wa88vSUif
yKJ57eMmAncOXCiq639TXgZ45d4+0mC/6VFWiMkd5WYSc4liAb3JKcTsNx4iVj9s
jvJUhObLFAUyU3u1JhHrsCd0lscumFGk98x7MsJ0clWdKNBbl7MHWmc0NYcpvaje
x8uWUiMazbPK2fctBibInE/mTANCM1Pmz2qN/J0BCtsBjJ8L++L+6pNaCyMGJ+M3
/n3oSa1lfTK628I+5ElOAWGQhVjBJcogzibPTYqDdy1/4tq2yxR9641pmBnOsOhD
5svTCK4/XRV/Vve+U3RQ0LY4RgYap7Il0/tXPgnpIsBJc34ZGzD9QZiy1Ipjn4u5
CiT40794yb8/LipZ5q4WgH69VXwmmUhpmdUe2YnsfoFR3R3ADwD9UCC2GS/GOb1h
BYMzhpr058DX1rNR/3MP3QJvpk6rIcgzSQ+uMLt/FuvF6zzlCqLrcIX8joma4lIx
C6Md9cT8EzxCmsmdEugzUCABHO93MaDk9JCc06FqnGs3V+7dXUBZ0UmH3+Cd24A7
+HW/XzTds19SMuUxVY8kSU3ADkR0W95XKQL9AoBzYol9wQLwnalMD+Zyc96MNOEy
9ImXAfehF7aTr/ZqVAax8v0PBti8/aOabDVw4GWhTlzxZvcSgDjMI0NkRZlUu2DP
V+YXiW1zqCwqPuE2SW3XuxAOxnM80mTYleOSBJ6B+U/cVMYETH+Fo673yFrATBGL
tulLlS8ysYLaqUY2KNYr7oboToJ3MbbQvJWXRCWTNMNbMkILWK6SaogcP1qnS6OY
R8cAx+Jt1+HqUDhJOm1TjEVSjYo6AbE9g51zERMRVLGpjyUn4kOmhRTtUVGXJ0Fn
6Zfksin6xNP6jmJ9J6MvaK6QGqlcELVBCwyeWwNZUNPezFRxQM/rssO+sET/YpAS
dCPe+RX+gUsA5Ul78KAHDNq8bpxMwaPfh8ogNIXExp5+gqjzyfMBs0VJlYN4yiJH
JSdkHqUbF/h2KstVPW/7XhoJaIF6ZVGAVRaOq9kNhm4VrCGpl7qi9MhKOA5XNshk
QkLyR/nN6CE2KWL6AOdDgbIxcYZ8axO12p2NU5snYFJFeHFFz0s7iZgaCLBzGeCy
bKCvF4X9HOJ/gcTLS+9sYjXFThKoBoIXCyPqxq9CjtS6D4PC+i5/d6ICtbNIn/ks
7rv/dSObhAMKguQMfsDV2zXNMFyplZFp6bLMeBZed6icdeseZTcrGlJ3sWjHOZqq
1grb1guWHoZjEw1myTeC8PYlZKZajKZ6py0Mo1W+qOTlw9PdsXwN4SjEJFJKBlM+
+XhxzzRO0ura9lPWFiPZb9GmfB/4VkrCTf4+zQavLOP0HLRRZjLwtzIPLu1EpHG1
QcW2C22RwBsSxLG/QQ4Ms+tdSRBWlrvr2JQM25/PbpQ9kYN0+PjQpLj8/ikaNqpE
A7qzZDkOuPB9a3urNkf5x8leB2MknkABFeKR0m8Bj4gKGNLeYjTaeTRzXIHQs07h
fMcIeDCF9NhsXOTcan9Qh8wzRg4GlY47HGXsnJ4lTBH0LXBuv/RM9p/3Du20EmzK
gaBWiKFprwNROYJIMwLIiuJPo8w+qmZdLDLuifHz5n9KYNoGGQFiYVEi64pM6lRS
4Ib0+rfLYJANDjb2GwPKtCgb4d7ZjYrCiqJrTK8fvUcRtttG1USHixN8iQoZw8Nh
1oWsK4nMavj8zu0BNPQ8LLF1gQ6SJ79ozRhnxo8JzcsViuaSisLz91V3GaUdvQQS
OR71zCWVRj/C2DlN58jM/lV2irs7EM2gWPdavo8apBCY3+PoMQd7EO5zpX8q+Vkv
/qrrusyPymH7Dq26XdpG0R276ykzVL1RzgNsB9n3ntt4XNjGG6icN6+CElm2Of74
WaNRVUxbzwpsUpkT5KXF823sVyPoyCfX0yBoY5jyygHgIDejdjAYKSh3lXl1Yq5I
qj9vXKQviPfhZLT8vRrLuWrxVyqJZn/2TKibPVByjcUbm09ziwamLhYN91S42GJi
u+nl67359Z1Ql6UOyolPLvMMIU5ElP1cMIA/SSwQNYHErYBTPq3XjMt8Q9g8yW+Y
puNAelJ1dp5nqhhBUk8SZMmgJMOz8uLIqu4bH6oZA/uCH/R5KqyL2abKNpdpIeE2
9w9uEIDP0wlAP7CezJ1ZDTeeaMjmEVJCj9U9vgS2tevt8J72l2V3fJ8Yp/EXz2UK
HrQadxzMSRdnP1+g+E+Rx6UH5YeV0bVn+fyZXg6q9T6gPRAREk9H77Z12xHvaiE2
qrWdyfqmilOYOWrOkjLwHa8g7GH46yEs+8lNksx6i/+r9bUiiWqHfYh8H6CAHllv
if95bBfFhsWfajHH5SGY4sUFyrOqTdj0ZQPIW/gD9dMuIVrKG0VLeszYsY0cxOKB
dm42AcNJ3mEZL3QhNE4xLuBkLEGpy/rxM/CAIfD00NfSA3CI95HN2LVYmCElHi3Q
CAGZyEUKYySEX/IaU9IH+6qnX+LZzxlz4WbaczLlSzZj4+wvdXIHt/oJx+yehqrM
/Bk+0f+dAQqhBWpZcUALQWxWB6DLxA4pUwA0ywIUi8mA2mZLaDtmwQQz3GngUKqi
ZnVBzpooPoEu9d1tNs901PckN84aeuBf84bMdoUzRSPLfl75mSSKgKv8ImMIjDJ0
6o7CLxp5x10oS0YAllH8gj6xLfo0pPg09h+TeoqjfeLw1I0F+Fj2IrFjOtxjyN/M
skPqsl2NQHEORHu5EnyGXyIbt8bQjsQRvxYNPp5e/vc0UEeVo5wQ9WTDQXNOl3kc
fDIZJ3/5tDq7up8Vbq7ekjsTPiSE1AyfCfKfvycY9iA9+UwhV5o6om9kzfj2tO8f
TWxnVXs7SFNN3SHyvr8M0zk7mxCxLli7ywUvjKSjUV0lyvy1sbTpl4zKEswk6zHp
/ff2IR/hz61811xz+4ymmslOpta4ovFrJtzYL1HqztsgH3kQ5bOpwhkcVbaD4zGn
nNsS3jMdOUrvwHFFP6XsbS9Wnex6apXxPVzvT2fMii3JLyVWWMfz/2Du0aShyF2P
LqaCY5jwTwI48V/+OD34O8Ni8p7FvSM+Tf6BR4QUPK0ge++IhGCnax6wTJNUissp
1CAHcACDMc3379rQ+h68Z3DQlOFAnFkU2AA4zw+X8rbdvqjogoePoGR6nZsN6Jka
wi3YUqoLuA3/j4zb1hucW9D80XMVIaooRNYJwkEZggvGZkzscBQ2+gPRfE1JuUhO
NXzou5jaPwgqtab4gxiSwbyDT+kOYze5bRyq+UFiVv4f4Ff4X1mRXs6EA3bg5qzB
2CAS/zWQmVHGWr4wJQBCShgIGyj0082d0xLtJNW2+KZ0Mpsr7kX7KTnDt0q2TU6u
TVHquGJshZxt0KknnB+N66/QV5fpTU4Vme7zGDIfMzx9ab80TXRfIyOzhLye+gOP
8Pn1/k6NUv2zAcTzjHtB0TsXGRuc1rXH2V/IAjCD7+p3r/DqotOU9TrMmu3RO8/U
dO+QBVY3dfqQkDlEx4F31ZXPlNt85xOE+eD89+wJgizDe85j+Vb2sIqLClujXtdH
xCeLYmaaa1NzX1qNa0JKGjWQfAQLdZLBsfkeDCvJUQ78kB8iwFgctPNLN/ASMkAw
xO5ryOFU7NxqJLCxPMH1MUPJ8jYIkvZNNArDrnesz0F6WMlQHLqQNUqk4of0k6Gu
wWS9XgnoBnAUnyuimEO65+c160wiG5Njc4xgz2hBSOBCMvCqF4IC3F1f9B/rE0ea
YzmRayZ4C4SSJeVwwR3NRKVuHr7BNWmuReF/nedRp4p11BhObZjpalm37ZoWO7/p
9Q6YwZfqsnDj8AdhCb+2BTR3ApxRQoOYsll13Vd3oiUOxarK6Ve/ilmv8DkviFxO
ahJ/IWSK1Bugx8pl6LiNMGglmH+/1pFXp8ZORNILmFkJWgoHlOY7Qnd/uf9se2/O
V7y8HiTBfH2xrPFBMmoQarhbNh9T432FDWFYepPN9Wxq1F3+Ay0WrKkCKSQZhyO8
NzxFhXXAbtO+PiD345w1nAekjomnKjEi4IGWtwv7lE1dYPx/8w25GFFaF2Z07aFu
izBipB0nY067ussOwsMsvh+1UjVST230Cf9llrsGMTx3sI0bLp5xL5NUqWh22RJc
dBsF9TzqCcvtvJTSMKd56FErUS1tHiubjeAuSiE36Kg1RK6Cvppw7RfHZJLHlbSh
n2lJfgyFH59elt9EtcNcNRm1IyhoAB2DizIrL0v8BmOzZlmU27FsbQJfQzHJDKgy
y3tRC4IlblqpnP2UFd/mjH4X4W1+5LsaGYqSwqdOpMdj7LufHu5ba04dC1PBTI3C
Hj0pp+JY5vZYGh18z2z9cWKxHD2wX791hcLZlnfCEYbuxzQUke+U4sQJps/XnSlW
ORmfr0npYp6Lwb6rbbOOHhB8YBNYPoK6A2oxh4zSqWOIa2forfnmZwaITL5obDNx
x4i6lTUoJGss6wHWNoSxaBgNZrmeZzOl13DGwbG7j4U8NHZf8rU63FUNCi5Tu3/C
kHRlQvU0+92aGoRiXmHa+ugAJy5KJjJAWKZsRCoEnHjoVyaeqahopaz10qLKjeXF
mNesRc0Ln5tFeI5v1NIrc3RizCKBkclPC0fNrlCFjluYRMwfKwmtkDBLkN9Vqxdh
ZX3/+EryC/kLBJBPTvErgjKBEeMYjh5DLuFISy+1DD2/lVEVOWKwedS0mQQ83ibM
ZySxFtxBLYeIaTSSddjGRCofmp+CUEic9eItercGcuRoGuY2lYBmHWj3oThrcNEN
1I0vTrvkimmlABMO7rjaXK6uoPk5w9BYRl2qA5jFil99Pc6PANEyC4UIYVTVVdDX
KELreSlAjq0AmBxU2aE/qQ8q/MihNjyRSTEtBthbIB2Dc7mn3XQzQEjUDgN/kU3H
2P3+PX6lf5a7oAUDJrKTuMm8ZFQNTGSU+EU7QWIL5pCjFXygUo+E0R8jVx9t/juQ
ytsz/2G4xg/8+mkXd/u6MHtYn3KAPjpHv33OzcwoMMUC4sp5llai/homxw/gK4Y5
pwwP0YAi5Mk3h4eOycESQko2LLHl8wuHxDRs7MLeJXEOtKcZsDw8fROygTOoGEyx
wNv5krtV6+jdS8se3jPmgfVwo0eMrPYdKqqeyFXU1Re3MX+DZiz/ieZZow8lSv+C
6uM8kuB+Cj/uYFq1FbqqeNqa6sSuPy08sWKnVbY6Nk72osAs0NcqwX8CoSvnlOUI
251uEFTRNRIwOoe0o3A5eAtViYRKBCkWbxxqPBS+xpvTBDdy4VJyScE2zpbOHoHh
2OKpzNDOHwnpGigdgU++SjXqUPN7+S5jerkFM0bXNAM/h0vrdNC7vqhDztYlVjyv
mouhzJFneHNn1XyJAxAlCUK/mz1mCqGupwvBv0Qs6buueu4jtRgHJMk8DxKsyNN4
YxNUdLavX1kK4V5JQC6rrJ5ULKWEMPO2PSQb1KfHH+jbMPANC7uIr4H/FGzqfHOB
3Li0f2Izm2jqxcaewfV8CofNX91srDwewimzLydTz7+HipveeR+sLePCNBDaMnRf
t1HPw4VBCLSec+cRK4hnRV9tDeZzAe5lq25bOvb144RWo+VNQ6xtHZcYZGXXB8nd
K2mVD4DC+EFHGx8p4At5gHsGgGf5DSULZYpUkAbdem3gEqnBMz611TrjtXGt9h0R
xy1gWJ2peWTFixJMPqpaU39ufOuRvt1lblIp1/p7n4k06aGaeq1NBXa0zwk8ceSZ
ph0+ABXRzPZcoKbJHX6CWAHsJ7eg+JyuvMWCeuqnE+CiQn6M3g0MjnCJ0G6eZM34
IlGjKYydYbyBGHpoFtKlSBv4TbIli8jLHohBitQQ45E/IeVZ2AJnMQUrqVkffpa2
dyvZIotWSd9BOZNpZIwRh1iu8RA4a0RVSonD8GgxTsegGEJratkB5W+Of7Op3w5h
zNFdH63qC5mUTVXjtlx9z6AgT7SF6EWZ8LDdExiocHOhRBcWPuZzqiMT9Syww79o
xqsIimrP9F3NUgLFzlX5pyjFL/a3HUl5VWLsd9KLstZvzIk3SyKlZOaESVCKx/Wq
MuN6e2uotOJQpOsA+RNqi3GbbxN0SWsXymq8HMyL6FzLGx7mLIy4QjHh5ZvU70bs
6evgdUi06FMKuVgTSb02AZKTzwQSzA0BdYNWq4ViEsTicVn/THTDLsJ8MLDdWuKe
fdV6q3MF8e3J+A5EqDevno7E7qrGmFMc5bjs84GuERFxoSv3aotiIjNj451sMzfS
T0cIpvdHxttTi6Hn/jwjq7PIMnqB9KFd0B2x1IR25RH6DIUGXp/xlNSnnlQRGC9v
AjNAaOYFPuSvi5wg+bmV4QJSEP9BHmdk8iaQMV2CPL8D1DPyhDngDpbHu7IPotD0
Y1kNEkyBLkm8ftRrwlWjCy68fRHC/qwlUNxD6AmFxs4ZSmuwjiyjtT7iyh62R/NW
Kn/jtbw6j6ZyknaCTyFqifPqcLshf4AOJtQLR7sc6+R/m7PEp9Lzra8Zuffd2lKB
JFWl7fqIkT2aQJIV8kFKj/FErT2Owj6hEAmzrYiCzajlWcwvnZR7tXRSi+xh69wU
jrjXCK5iHa16m0HuGfVJeK6CB0jd+uJssyL7lUxQlshqm86E4WnY2UFX3Tsi1csd
JkIgCic7CLLoNOpTQtwTO3dtow9K9eIZEW2fPjQyRNGR16DXvq9WCNbbMJdG11ja
MZAzZY7C9JRMTBJzjFUbOiP2zG3vy7vUFqm99Tq14AkmfWiK0DbA66853SK6QP/S
4BuEZH1Jv/e70zFTwM5fzBKOOjPXfkCXsHM4esuLdHRzqSVEgkUFI0V7mfHKwH2d
sbUAK46GzVnyc32HTGqEU/RiyU54E12+OUkD5SpYdf0wtHCX2XPjzQWKWRhBigYH
rzRRL/llNJp2bEM/2Hmxu8bjmDOUNBly4IJB+XrD1XTV4LRQGdwnYdTbL4ZTQYH1
ztJW3J+aZ0B+cyjrAVSDyzcprqovGhIKd+e+wYhLFpLUqwU2HCeWmHwtqCuTMKSx
Ro/vH66jHVQIoEN2Fqi/7hBwRg8GwRpDa3XSXJGmzIr4PyBiEVPO0zEtVBDaVqcF
lZL+irFASDVCOO25wEjEQNKladi7hOIBhzEGzaHRaxgau8BTLgvRyYz+HlPMv12s
0B7OMgLr/eCuiwW3BsjR/1Gl1NdupV7Ok5ZxoPlAfVSGnPpx3v4XnA7Gt/uXpZtH
EVOk+Z+ehpJljBM6jokSwhVQbZah2LeeDmin5TwkdDW4e/ERKLZEq+UkjgPWm+Cr
k7MtmXCEG+pWdZXG9r0LRE/YKRgAN85iNDzVL78a1lFGrMdWS/RNIhmy7DqFmhCi
Eu1rzVxoEpBUvsApanQO3YEmTP8zpM726CnpG2ewKcsJj/hQAhjNiDGvAMnDJFoQ
hhOEit3RyhAFGKJkDUy5Qs631xFtSJD/rvHoWtS7G6g1aDKY75BPjQioIoHPUyLD
qPAiZfr+3EjHqChbFjrI2vJLKuI2ci0YWvFaqoGYeOBTjM1ilcX0xQcQMx3AmAQx
5681/Fq9dZcz5Sclp1KeHoBeHtz/z6znFZ8SvDMNDfMJ1Z8WGnF92KjppLRsdXjw
p33BmBg4dhrlX8toMQxmAXFfbqP4WfsrQG+E43bGGZcOStoXMX2VOSXq3TQ/XL6L
Svhn4KnOKuMUI0et8//AXqyTHm0FOE/C1s+70VNamiS3vj5wEGmDHnqh3aiA66z4
pTjirDiSoE2bJxS3daGBaC8d42snTRcedeYi1e0nYjk9PDICPaUTJyDdY+peXXR8
ETN+pqvy3TwExu+upg/riqCWFdS6LeNZfnDA2Oo6BqVERJlFBbi4BRTKCosfbUy/
mY5IHpo6cG3nGusVzR8eZqbqHDULbvPKTWFOqr9D/oldh6ZLtu7ZPFBnBkg6QIkc
Pphjjlx7sZGhjLRW290OHdjbVOK25alupD7u9SlrHdl/ksYnoxYdTjXj3FltWnU1
XTrTtt3CI7Yjl3kSA+NGd12fV+mII+5NijtWcGilfUHyi8Go7WzTG+5/+/nsdOaf
6X5YOno6i7b4HKmwPCb0IZo8rvevW5AnCLayhbkkgMlIGfDZlFkibKLtxlhmK0fn
y/oCfRk9/h4PTJ+babhdkh6kZqDUb1n5bmuxWgB03Hbusl4HwNObuqEoNaKgWX4a
9zsX85vSFuZAU73NqoOzjOrJKZMpG5G4PuYDJTC1Ad+Zz4Jnshu91bdy+H1v0qA/
YbGGTjRzb+vpN0vxkoQW425eZTzqLQMQAZme5CqIAiOTk97/MOZGV55cVn2Mity4
V0ULoGevKUnkW/SworRQP2z/Zh/NmwHtRzfeDO1MzT4SFo1EmNfZh/2Ejz0zEAHu
06ACwI9LU1mRsqZwJ3PHtBzaN/kBs7sh6X0LQ9zm9pY4IodGzXeF/gbc3h24blM1
GUn+5//ENddIrdkpDtXlTdJGefX/qhWoooYV2Q75NOHK4O6gGwA5nkC9RsWyvRd/
B4GQuO7nzoynRrgz/UPdVa1JvJAeqZWJrr25MCpAJs80YQfZHILl8e84FECzT7F6
j+86gyRVz7noH1XvZg9TApzLeg28wZmYjh/leKS9Ps6krVXoNup+aHdg62H3/aG+
g6eqqJfl4FHh5LMm4YsfKQrj+Tm+h7KnOUlqkupaIbR9Bfc0oRTZs27aL7ISTIYC
rTJEN8nhes/X6bCF069d8RypJIrsweIQCowH/wCbtVKsxyPJl5EYXQX66ckUArW+
zxVjVIYDZgQvV4kfMK5/w6Tx6xgq/fGKXkdiDlVjHFopLLsS79ZdTTCxQNGzKSSC
ftTRHoismse5FOjWg9Sf/q1ga/fcmbBq5H3ICDM13+7kak4GYHDg+xmFDRdNHrYL
E2BmAPAZL6/M8Ct5djNCdcRo624CEbLCeM5RCBGf+8AjJ0uQYn3C4Z5IhRsQowEf
1vaFo1SnXL6vSaD6pEUJN40Ys9RjCP2CqvjrG8jOi9LmNJQBLJor0aO6Zb5T673z
PWCx6PVEWikbSc39Q+rtGEsGYGbjg2zc4T9N9I4ce8a2hFkxBncfsYXtHauN8nfS
6n0bVAmHKJmvM6IpvsEtbezzGDHNWH2ZqdBGTPFRpWT786qCZd9VesJlkErrrvEO
TZIgqykVTQfsaqUmY1djfO+rPCFY0/RyjQWXE/UkFYdtdT2GPcnePr/L5G8h22we
dXKaF2kIa2f/H80KzchqJkXbdTtw9LXqq1YTCTHHbPsxE8AX1CsWojRIKYO1kFU8
7ZCDpfh7JovATY+JrBXkYyb4eqA01/brBJwIKCdvEZDhx7Z9OMoCOqY+o0rhlyY1
rmvM7oYxY29yWUtcRUUyYizZjikFl1YthIjA3PS3VjEpd+ryy4wMOigpIdZ75ssZ
7IZ5RcJlQH3d5g142pXaSgYzjYxQubMN62luhScry21lNE+7oWXYz/rqf1I+Xmxz
+x4IqfTEXKnuto/XaqQoC2hB5SiRGpZLbU8KzfIEzk+JSwyuqjhroCm6DzNKXe7E
Nqf1IJC54Vxuk7m1oQYWJav13grfMMBUP57crUcEekbet7G48N6NDJuoyoJJq3VW
SE45lzTlEEZg4X8yaz3s5P2AHybJqLB7rydyIlornOcbHCsWXeYRCGJmQzLPJHrV
kAqGH9S12ylqLDCKQClxunGcoQzoH5VcU9Ems+0cTnkNkBwdp1FGVoUZnJS3i1aF
k8zy0YDqvWaj5eqy7O4xVlxg63Cv7amLtZMlC8RVYLr1GkhXJZ8Psh6qlRg/guv+
9emJluwVH2KOJDv44TCLxb3MIk1clawL9X3o7G85tml417+vKg+uZBaj0JwiqmQv
4MK7m92kporgRj1YpYdrCV5moaXrwTXvEiGNq0OSwQUyfVu1/gESnf/BkzyXNbcw
TGNqDBa+aGNFnvXUyOH52ayPrXzfJJJwlRnZDjXZaPEKCN6cMx+ik0q0bYafZ+l4
Tz/TPVn/9ryyI6c19jW07r9r7K0QN0zdcOi6Y0+dvfNyxYhKc45cDklNsm5htjF7
RZJmECZ5H/5qs5Y0qpQ3TFMZI4dS1QbbbO8MpYsO9YL/wDD0TTDlqZgC8s3kZyAl
CGNV2XLJtIidjuL4MPOUye9hvmyY3yu8wpYBSN7dROObn7Xs8Ir6DWC78Tb98JVL
VQ8MngvInZbVPqH5ntK5mlzxfQVyFWCcoVxlGiHP2WAvQXDbWJT0nSwLCPGDg6PX
2Bmmt3jvav9VBsbG2IPqXAZbd1F+Fg0c4A/TQkEulPXEJQBDqCS4tBqOt+X4o4Nd
9dG+t1VwlFzN9anOyFAfOe21TUsqo5MA2vCsAQ7QEdvtfqxQCZdSyOaBWWMtYNJ3
WeD+A2JbnTnmEncY5va8MOkatioWie4JoYI831IOoP8lNkmbW6Tn/mb1J9v2oly9
I9bR21iHi8cVTjMGAdi3BdEl+0xxWw29yXqRIOr3LIAXWrm5Yr6cQSWarf8tzYK+
1gHgv7oHhchkx6degVWGpT0szNGCu4H1jsixern2zlCfP1BzKvsGJbIqLT28RdyE
xjUJhpeoApFTWLOuOsCFRXmxq4OZ7MiufFtgHgG/KGrhdkl0J9YCM8q0t6tSEn2+
LwN6evmOdUSC4ZhFLRDT+qi7S+TnmaAnrKBZ48ihhl5vH5Mvo1OT5N85KiVv5XqH
mMVltSEmVdMAL6wd/snj2+uDwg+5tYg76hiK9vAhm+GjR6g2R4sQXvue0XhXpDa+
ILoUdbelUDWjsAcNyGtRl4lpTT7S2iAD5iHoRwmshl83nldv7Ke0Uktco1aKb6Et
FDYUHv0Odvacl9M2salBbNyAGQCVMsFv82PHPAZvqJwjzc9pIPLEzG3wDiMHmTPH
jIZCxy98V93ErLW8hIWkPsocwgSGfoeW7ZpoUhjiFrgZhQ556VvDHd6VdNh1NVyS
DUaKn54wH6PQUzP2zkW3q1G/pVnQcBmuZMOSGY1gIyU6VqktE9s63J0SRoDKQxqq
4ciZBwHIO39EkujiGogao6obMWKGu256PlM6xJP4owDXna4M4SkE9Py5QPHCYY4n
pUA/QmwufoFVWfh3bej079s2t0DrYzu3AktnraDwfuHdiHhuwAAcMBkJX65fq7Ux
eKRFLL0/YWtUxsMI2rRYdheOqDp+vUgnuV30+Ze0yMaNcmSDTac6gqJs0YdUwWht
N9Y31+0/3qNIu17W3MvJodQAwwWnqzcM0+s25jw6ZCgx8JWog7ltoNRcKUj8oCGp
DMwwxrWNUWuhX/hMhfD7sV2lEuV9cFRGZJ5WNzbnDyrd8MQjs3tYV4pkYTvXBrx9
8nMujbxgEgMYcx5G9mEv3gZcbCQrf70mwZV46L7RjBs6t19Veu6pl9mCCnc65bfj
iUWmCKlW3PcWZ7FO4PIwh+qpAbSY3al3s1BputazDDhwmUnk3sNrPik3ow4LxfsX
q3DItDQ9jGuXOqGRQSZyriWoI3dBJ0vEYaCFRaJlIWaLzKLqm5/3TVLGoEzOFEI7
kdCR7Fq2X2i2dPm0GthZwEpigFCZW0UWBqjv799JGORFNTFMjJFVehZ9sKHNbpZQ
51dmJUJQSdBWD3/Vu30unTx+IschfR+FCSxvxpEjuWLRt+OEdYaeV7PFrKRV2ptq
q1NKzRByY7CFmHi2lJGgEpncdzfUKtZH+JtunI0wqm4frKYwRsepML1vwQz+bfzp
Q88b/P0xnVIqTgpnrwfE/ztbquTdvEGRxmpmUhWk6ZU8aZiorJC/v8El+u7g5tIn
5FBV1R07Lw8yOacSuxN87gjw/3SBFhZ08Nw5+mJNN4e58Q1ojqkzzYrZwnPUdxu7
o99mjSBSlD9pD43fTxlbOitXkY1YTpffaUuv54b5tVVRyQwoPsmClnYEkKE9V662
cT5yAzQdzuFoCn1pm6Svmje0hRT30CJxXCH73Oj0QmAO7iB2s0EnNxJ5rmIWwLu+
NJKBIxM6rI33DFNrTDkdAyj3k/BsEQJ6D+LoF8AMHavyK62msBnjwnoj77LWDe/s
6JBhq5Y5XjdnpqE/rpNzJQIeSZGJK6JrRQABCVJuBLzAOToHzwZpat0zeYJ4TkKq
LldKZRNn6SW8HjgmA1O0qQwtXNY/AIjBE1m5sZtiMzkPs5rCPo2yn6HqFzynQ9gP
Ewrmr0LmVojjfNTIUuW8d2JvyOL8FHSU6cwCV1cnH/SGA2jS/QYUgUjL2hFnYB7P
y6IRbp9WuPMUUjoiihGjFEnpDBxf4XbTcSTqMlem6W71JhAaiGWnGMXTst8Iht97
t8cIytbfTmY3/+xehiSnz8uIoe0ia5O8jhtKY8E/5cimaxTw+i+MlNqtFvxmKnmT
sMzI2GuBF4jx85I3Dl/+4QzYdbbx/LJ3Ul6SRxJaZiINSakeHsAImwD0wR2A5LxN
o3xB/7elr6CuYdnfh+OSRiMU8EYsCa/YLrXLJ5eX6JgTLv2R12P+S5f6QJWfq41A
dMC4QxNK7p82E/ZOen1eiqvBUivpGhfPnpqpUU9/PnUago5HxpeUq5mMyQMiJQPN
GBytkuClG7u8eAIMsdVn1v07ex01ro3/a+ELTfZaqVK3JNgcGg9EWSYWFoUEji6X
/HUsdv9sBGXLQdSa4GBfuHlWuZQtvrhIcUZEez+3nW+S2qM8rRAVLg89zwy8GD5A
DX4GndNX0pDHVt+ngml5lzaNoa5b8YYyOm/3uzzOkM+ZI9NtMWGs7vnUWuFHrdzs
ocszmIwN6JE39ilcXvCPi9weidPX8Hu0zSD+qyh5VEfab3q1iwGpeTt2agpbZbV2
5vXWQVD99UleuQLlzSGSuZMswJr2Y1LomTEiIBo6wU9JMkmJTWXiv8GqrvDC/PP3
lEWJg+CXoc9Od7LAMNgAlPpN8jyMQUxAt/cts6p4nFsR15EaHEJzuMtwM5VDEiEX
johV6bCD6QgmbtjNtjnkSdsfLe//QbaQvNwz1ZXycPAzLrCStnBGk1ViCLeG/rQW
Xa6m4HfvwdBZxmHcOHA+tZ8Qgq4WGKSAyDjM4e6eOrSzxiAZIPuarw+CWKhZbNKn
szWiVut4ZmXp9O/Pt0hHGfcBNJJmQsWPyabEK0YP92LrZYZjaZ3zl7G40e/mYTAr
4teLpvGZ0qkOFBLx36oR8dlFraTdBGn0TlIkHp92e71k20nMHZhrlZwkdJOE0F4q
ntapLXW4OI0siBdirSyv0z7El2HqUyUwLPXZN4KsxpacWT0nxRvh3BlYi6/4LMRR
WNoQPG6pOZPZXzKP6EZscuCAZYtoP7AsY1iwqDqwQRgNg6KuL9ru4ujJKvnq/vVU
uhzUSMgmVzxTNkDCbfglUQewvLpfPeIYOif484gT546pEFiXqZzsy2R1dXRpRTjO
K0/P/N4OrCbThUSMnyUOH1X7nL0hWaw5eupuXDq3QQZneDWSz0Y16dAJ0t8jH6a3
9b5GH3KonrzqjYLIMsNpcd+t4E8Q8XjqTF8nQ6org1NaNNXrMQI4dLUi/CH8jAZ+
zrKfM3eVqgr6Set/w0ce+Hy/rNtvqEj90f539Vk/hQoFEHOVZD2caDnGfLMH7g2p
FnkQ2JITmEtJtMtVOIQ5LiMkv09XSmyp206T+qUrAoMSVlHm47OMdzlIqk29uGR/
u0Qxya+YWfMCprC3QSM3MgqQII456OjHDIZeTObblDUvwSZh3Q0kxvigBOcK16ql
EueaDHuFnt/Z5tsUUQlMSt9A80ALwggu5G0E4qJaIcK4wccnaVHSgGl+yn6jU1YZ
WpWh67cAgghMv6QeDKzDEppZ+Fgg+0bivpbJylEdDSbTel81QcCXcXHao1B6/lFM
rflIhsktxPktJ81R/x7d2xTI9vrC1/3vdia6eVFBtLUv7T+gdsA2ziJoLynHHRZe
+KTBJB6gTCvd1hrLROk2L5pSUq0C6jDoq96WpKfqd+ikVaJmMfpgupD+sMYmLMoQ
HMd9W9rE21qUKLTda0QxjW1r9+QAXMnoxBAPhfGQVjLR7GzwuUOmKE0vkja+vd7S
jTNyR13b/H1W3pEG/p+tEHFiUHbM9aK7VwlSX3giUVCr/mdIHZJmB009i9XiBKjW
+YJmBZquuxZ8Zw0ke18afum+dzfggW3GFDm2aNAFqK3EuiSN3VBNNDKKHvZXHkfi
8ciBtlSNz7LEdQh66HCFlD1vhEgwM1P37rJehFwVESnJQCK85H88O1zbqVM5Vjqx
l+DUEJ9RQJyaPeSNzlo1ILhEHBmLkXl+zwRxvBClN3ihO8nIn485k9Z91Edm3kxd
yotCiFMmtqbLMFA+O5XU01RwshwfdOnu4cLTURmbp7eEdYsNVR2rBWJSZoSmYgGu
Ep20v3S3/0G0P4NGCINAuJTRQT3sN6XMcrknG55p+vRkLEoiwNc01idCg2Nn0s+4
X0974nBgMISa/JH6Al7Q/gYb1VfRnvIUEsS38BAFuTopCBAlZPlMS/m7OWwbOZ4p
wF2M4pWGTRp6SsBNR0Sr3KUXncv4KaaA6u8CHEFaiT1d8+w4lSl8zj0o2cuD/bt7
uyU1UYmdi+xJ2/qHf6wjQrVvmR4WmmX1d37F1hHnFfEODvzWfNio8PO3ds3oYrak
NDth66REEdFGdBiFKecdatXWFhoWnL7/ZgL8CZNWS8lojjuEh+TT84I0f3riiE17
Z8MprNMRhL9aGs4Y4MxNUw7wuYZ1qcoOSMBLPUjlBQwJqoAbP49zVfVLDSPD6r/e
qsTknVMQEg6+V2Xc1L2W2lWAo4B/VrWiV0qHH4zFbqgo9IS5Ab0ctQTMVGAu9Rcd
cqD1lYyIn90yM3TUNy784hb6C40n9wqV5wO8mjdGb85mYqOqFE7D6PumI4ET3UrA
EdRVgpc3tBqxvjDWArFwbgB/KQ+sXlffdjBUFUfk20oZBXm66AmFYPe5sqRDR2a+
zUHTc7rMZQWXXQUhwCDBPRB0KWtuM2zhII6fb3E74iJ7ocXx3/37hBQiRGG9qPnC
EB4BQesy4KM7kZM4kA9bLhCxkQLSZqHcRXAMpsENerSIz+M4RvRUGp/Q17BBaIsx
Zkp8jdEpBsVpqyn0x1jF7iFDIVl7UBVSkybHa4Z71A/9Ms7MlHFIuhxjHZqEN+qw
P2irEp2x03XjXJazx0efT5w/tJfk2WFhj54RqoO8bqMhPE136qbGgwOIp8CjmKq0
NrnLs8+/xe/ve5AABsLClt9779dwaktNR2XgC6kVRprkZDudSSoMKfy0d686qUAB
GNm0zCbd4u0bp2Vs9KSgshZYE+QiaeUhtbA6ZECiQMJbJmW/HNRFR9GSI5N7hkjj
jFOGdndXRSE/ERxaeFKNN5Km48jQLyt/ylA5kxC8M3jk2gVjDSFr5SwpcjvgV37u
TO/cAFqmP81KRZ2OeUhzXSuKlODjRT7Ifb3C85oYy6JG8GNgzMSSfaqOcNJnTpyv
7BWAyeDjTpBLwEAEw5x+jmbr972evS00NusjGYn7JbUKDfhg05b8INcxgRGDfhXE
kHynpxRxuaYnAdKKq3OxjAiBkJtjuBff8jF2ryNQfwxKKaz84aoOsV2tXDOawCRP
Q6XKlKRrp9J6Yd/4dww7EsC3MKuHZxlLek7WV+2a75qtDqPQLaUH7sLl219lmmnP
zw7Zn2k+kpWsi++mrYFazp+vc5Qfr/m+wuyrFRAgALu48MFhqQSoY28sHMgyPhs+
nece8HG8g8h4b4GM9rjirF6o0xCXvV5m0z4jQH13VrKfj3x53rBCB7vVg2LAt2gv
p4Snt9L6bpSQ1AcgSW/jxSB1K4nVRc02DX3XybfHV44kvvWakIzb7DtmZ7iKwZiT
a+dmBJiDwbWl7JID8aKpYL6ApiS2MmGgG9k77kdkx3C/1qji9c994d68VuwB+yze
q1bqA7kjgNA3nxhqQzDayDzo+9JORWXR5qo0htwdo3mDvAUpwNPcRk5oVOxDKp8m
83R3KUxRvmA8Y91EfA/z0LhBIzUSgzjuyi4l9kVv2J6GpD84/HL3ZGzMlgKhomsG
eItzEjIPhX4ZJv0NiTjfkT+ueTMXZjTNiRDRPXMWJQ6HISss8RLjKRzW1I+sIeBn
W0q/kgKXHnMkeVMOqq2qLLlBUpa7guRromMGVcAX0nL9q60G1SuKVFs+REmiNxF1
hvAVwaITuVcpk1gXnMcvXCnevTLqwSMg5PQPXVyu2/jvg2t9ERRfn97nCVaTu2EC
v4CTit+b4XtWltdselckJGfjzByXUsdtxvi3NTXGy8yBXucuri80GetrfAU+7pAU
A1DL8bRAZl0aXpd2L3dBh6zTKHBUR97r4I+qUg0JbX55SVduPSVCXJfJCIA+oUIC
8WG1C0SjuZWGw0bF11xQVW5rlO+82J8n03nbg/0oW/d1jED7dlheZ/hAvU0sqDhZ
+se5B4JMzdvRG6CAlbQW57Rqbt6UNtMGJ9WRyr8N20SMx/MNo50E1aP+gTOL9f5u
79NiMtzQDueajscRR1VIeIJl3MBjCcDRe/JUuR7aQvewH6rugiHJ9z0RbiHcZLvE
YUNtQ8U0f9qZOxy5yZVS88YWueCmgCfsKh2vAwSeyN5oCxYuca63z+IgGlBQMhio
+/HBZa7UWNXoIHvILV9XIh9wYw2hvuIGmaFTTkOFEiV+0yl2S7jC887GPCHaRV3n
LOZASWoOf0kyvGGKnZ7sr1oAWMqWYK3QjoNgaMU/rLzuoUJAOH1ol+WHsOEK/fkt
adjZd/OLa5HglmPjKte3XvVkXbrXSTUQHgQviEHx+MzAm54E3q5Zp+rednVtqcCP
C/9tIr8gMom4fv2clCCra6JK0sclryq3htJS3FtFRnGGdW80GJi6rdzB0oKrAdyS
kz8DOTPZI4XPqRKV1Mc/L1jrk5V32De4/MqTdX8tawVwdmkLg5TIlrTCFdLuUXwS
YN7K0mYvhfoqKlal9oHwpvJsnj4rpwvp1upr3vPqmu+t5vmVMIjIxtH0RgPj6T8/
rPr1WZ7Tob/iJy15m540hh58uaXF7VJUf2bf/h7AkXYOZz1/ojJfLm9VkGHNg7ai
7HXcNuHa+u2Y18k1N3vpxL7UZH1pDnHC0ataGyy4KEdaEyZq79XDxu7psR2aa6nl
xI7IsAxsfji9GKQ/LiSJTnzhkj9WskygH5Jh1IQG982sJFWxnXxGNuj+n7cL0rnq
j70EV8uR4Lz7EH5OyvTkvYVKSLomki5+2GnXcjAdfTMl1krDulrzJgMaotbotEqB
z1hk+pk/Rj7RKI10o0sG08egOI3cp2PDrpZRq1wqrJ5EQjmgcjKzWfAUN2u1W2Xp
Hmrf5cHEDE+RA41O/ljqBV13zmI39LF5mkYN1veQr1HNc+/RqDj1EWbAbA40KEcm
e58tmr6E5FjLuFTlBZVkUkltgtWuOijoVNMajnpNCcWcdmJVUD2ab1H7KKKpX4Bl
T//1DF+INdJrSLFNMJfActRmtoS3N+vILGy6tIkiGfC6wjq6yG6Fo9HM1uGdgyE4
ORezbN3ZMwDilmIOHc7zwD/aKOhiSgXCCMizLJcEYMTElzXPcMnWZ21rdw1SYsDX
sRiwRjL+MWpmKdYY/6eak6os/8pBxO76C7fCTB00ccwrgNzzo8dB1aWIu6g5wIK0
WSVjzjPOh+ipKiy3qAvEEfZw1P280ciTUvix5eU6/OVbILtALa6NolyqSnVUIcO5
mg5TtlLGtU5WUDXtltIMX+69STwTDXlen9KVhawp9VpLyAO80I5CWMD/oPutgxBL
pw6nI/N/E4ugMGBO8RLwpBZYwBoHtyobN5HWjLlgdLZqCbQEpV3w1TUk99G5DOI/
Wydsuz/bXSKu4Oe4sFKn7qpMdXcr0Zgj/8FpXCgU9tpCywyy3iEVbLTGwQHDAF5g
k2gGVAcCRlaZpVwfjMDH2mZchiLKNvk+JzcUvvAMVc/HCNSY0OeTuMFb8pQGuy0s
dXRknkajFsATl/pEv+aEvisViCU8qMH8RiR1J/AMBVi0INcGYrt9repkFKHvVTgl
+NChW3CNQ+O3w/I+cv5smSMGV9MwXTiFSn1XgDkbKYlRL+2Hq8IkU+6BSLq3JBlD
ESBipx2eRx57upS7Nc8Y4f59/n4FLNeleRnyukOCtAqTNkehl3mel2wGkaDQKx1R
Cc+xLZdUfpJAi0vgZplRFqqX0GISZFr+cpVzKNk7QVj0oVBzzh4dOTt7YTP+fin/
aiyStLZY3KZ7VZVntL1THikSL3Jh+bNu2zGbFrbr9HMs5taxgbYdFi/EAwjtMuWh
BuDNVWDDly6r9EAutm49+VPZDZwJ/+myxkWsnVzKlaiF+WfOoENRNkwI63OVydjO
LCgTFWNVdJ4Y/T+JT/evMkWxe6joCvZsx6kSV/2UqYYHe+ORCh/4INVo4ZIwdrQd
m7ki9ERIgGWnFlXw2e/Xicn/AXCPdBZ5/kJSIEguOsMABHJWQfRiQuxwhs7ZDx2V
JHd3iH3ks3D44mmSIT8IFZRjYveGXzetYxkqtE7Q+pnfCeLLbt4e7T3qvedej6oY
PW4ppl6crWJkiQs/HChCvgPKMFDZG1P5EQyXQwLSzumVy6m8xi6w/04qlsQEAwxr
H2MjPCnIVB5SrV1ssXAXaV/rMNngKa2ZA1gkj2DTdsFrFBQqYxepf5mLjupjqSoM
Kvqkz3ls+QTuoE6ZJH2IMIxf9Qbygnv3D2Laf0SW+Cwtn9UQQPpNxYBUMph0bErL
9wH0jF1ZQKiQr8ahDN0kuA8odZqmRuQq0RrSmZlGbeHgSKRnzgG15QO8T3vlPqyI
oIPb5rpkID2nQG+INjWLdCK/ZiPX8OG0WUH7L6AJ+rEQAt0RWhrjxGxvsexMnh46
ClylenrfXhSJkWIrMVmEKcgX2yapceSHC0pr8Gg0ZHm0n5LZyJhBUKi8p7Boa6XB
Ywl6wNYy3wNLXUInXwBaVTxGLBHSN3EyKkLHm1hSezYsC9nmGqSbxjFdCdHIygrD
KYje1zY3fUZr9sj1LDnacLgvLzoCwUTjjVjV0bgDc+y0blb2DVjYT25h90bkcJqv
cpO8MDoFVpHuTDZH8emIz81kOAkvSBLjpqsdH6l+oOxYzLVvwu+KguwA4A+YAdY3
t0kH0leaQY6m9y7Gg+hLfO+KtRCgupIa8HZ72rrhK9BQAzoA1O211UO5Shv3Pzxu
NG8eqJ5XCEhcxWN7ueqG0LxQICT2YFDkhkHUgvMoWHWyTF1x7nYTXEcZkQ8IHrok
FFWsqstMDPDSQwka/5fJxTXTAv88mlkS4kZ1poTfCn0BMCUo/OXZe6IGNDlExfJH
yJx6Iy2Ype7eIP2znjiz3RPuBkKcekwHoWW+1dvzQ8VhQgjWMgeJNEKCtIartDZA
WeGeKYYFgqu5in5aZQe8DIVkBRHcdbxSMwT/bKYezyLttZEd/UQvKSl/iY4g7kJe
hFEOfQUXTs0/RA5/Y89fjmzB4K7gMEYyZ8FYO86sbQlM9lp7S/IPYuWWQPjH47+W
kS5UwcAya2t9ZSrla8F2KYjdGYvidBF6oMwT4Ubo46iGj062Z/L+YLgVbhy9wIN4
do0vVzqUjb3pB7zzGbhaBq/lOC6EgfeWOaRa8BEYKV0MjjhmJx+ma0EEVgTnA+4+
rbo+uC59ixYfe+gDVRF+vVVUzeYvvnM1Ufc4aI5PcHLNRu91PRbIzGS4JgDdcdsN
ib9XSIhMo9XD5T1/xWVFIbI4JFmH8LH3XZf05bCn4VTwOTZ7pJPVfLCz+5QjFz8B
Qwe9c8P1mttGzrH0+c+iP1Uq1KOWBNjPj75wR/xF+tUT4zZHWf4knjGACqFEOQTS
4QSzk4IJfhOKrArJ4xxB9J/C5x16iDRnwyjtHp13qGI4ypTFo0kfT2s2dF8TAdUQ
Fcurs7MdcG6ep0fieOD4mEIjEam9Q6+TnHYIfv4/P4rA2ulJ4dCFul5ayEBELwZq
puFfPIY+mCRT+DNX0NTj0s2bWArvi2E+uue17SgxvyMxu32zFsv4Sk2hdz3+aB0/
dUHmqElnTS3ImiwDi5oJTnx7kDynRtwlS7XkNkNHWJgJ6RoJjDZbG/o9aOYP6beu
Q7z9b8Ua4N8KSo68tUJMYmaPvwoIcpE57yqLuZW0M5+w3K9VgXU4iJkHOMvWCgO1
961kKRRw1q6r8vMcbZkBFss6s8g8Wm8zqDDjF4GjP87Q6nsOzfbt9Zf9HZ7+7ics
OgNf7mlxiAdvnTas9f6q+td178ePjJjMr7HQLleaF29j09Ow7qiF1OjqAPecnvOs
0fjs3/YyR2JrJ7aNnczTUAcjKhrTK4FCbQaQQSTEThjTOfRzOeFaWf/8CZc11xAH
z0aFmZlu7D2J/jFa48Fstm1dnRJtK/mBFcwfC1WqF+iztIOYArBVg0C4IgIKMjuJ
DprmjTDDbyXqXNQPljWiA8PtUO8Cwvj7Ery9iYpZQWFTJHCBfEYkLIvHyMG0U2Xb
zO/PJN6p0F1py6LHk1SEPr7hYFVExgCqx8BKJjYOQhAFoZ/nH/F/mZSLR9SihFg7
EFX3lwrUsWluCrMoqKKadKty7ehGsmT8Xr7h4hnIJu/NiZqth5pBRiKrtJEVk+eL
8peNRK+8m5htirC2aFdBJhkvFFWk3NyuYJn3XYAqZCuayKp30eC1YEJzf0UcLaZh
HKHt71bgYycXymCedBEX2rkbl9bH2jRw30rm/FHYMCyvBZD7qdht0s6VXIJ7oym3
30g2hsMUoes/N0knmE+1XQ/CxoWQAP5+f924aV9AiW3p+f0Q9bUFUOkYfjMtCU7r
tUUD24vO5rQIg8hC5Q6IfcxBxu3R0JEml4NW1IFfW4jFLsOKdrpyq16/VfX2dtET
d//jJ/KBEc++6Dv/v6ZUDC/M0Psw9MOm5qHbA6WkJpzc5NKv4a/jJKJSsn4Hs09s
eOzRAieRlFmsmW/LxJBg6vThqqLDgvFgPRkQEs2FilYF582DxsJ3zG/AB5TmktMu
/YyT/XzUdTZmC6vtNboqiCor1w7N6uc0O1sGZ6Rg6SdaBzy4IhxMnsUVCEh/UZJg
gTEdHIA6+ed10W34Pw1IRGS59MxKcq//6q28ltu4FlrnPul27lIMpMHtVcXVMZJu
LTz0S7ZKbUCiiHAo+ijRmz1i9onYTtY0HHisTpUZGFRAaoH5s89UXYIHZkjWIKL2
cWn3cbgxNLr32SBP/lC/HgfaL1FLD6eGHnGEOOFqK9CKU0ScjdcRr4aFyzGTkiy/
uw8Al0NWEyHa2X32i4oGOvr9WGc/eRKrqzJdMNi2/PM41lnn5jG8FA2J2ui4kk1W
DucuE42RlKeunP/OjoAKxQx/reYxn6X4NtIQz9mXi6ZjzVoUazqWLS3YVfH110U7
IoN/w0JzvZrLwoBnhYP0QJhNJcueVERp/5U5fM2TI0S9ZuiTL4RGWd4INqg55vSK
84ucSTSbBlpZbmieP2IAWZGvfjm8UxHZuEyKOuC0062lX4tgzqiJbdRu2A2MA4yX
W06jSdR4IkpGU2uaF1i5NV1tKKej3Fla5YRn0J/+omWfmNJl9WNyPHvwuybljwlj
+9gnbR1NkZyNVHulB5IWozmBQwn8qhoNZ7DtIUucOJerc/+9NtoZ0gspoWk9tA+o
gn/UDQCMbOpCRs4iM3wtBT+3knR+YV269/ybXchp5lQP7ne/clzOKd6rLnTABvvp
DWzeYacidFHYNqKFeUMX6njFyCZuYthCvgUf9oD98K5nNoBRwEFJ248z+luCFdOp
+auupE3bPXorh2iBU/KdY8DZXZ7HxzwLMLSzeaUkhg/DgG1EzzS7Kx40eM66fX5j
pXdgakLOqZ8565Vu8u6fcL2bV+P4pprtMFU9TTkvwODbPsSsmH+u+fOJ5z5gOxyu
w02I+npxngygpp8iSXFoZ00PDQDvCrJ/gcxItSjNNN6jvoQiVsQGIS15t3gvTf5A
hB1iNQzmjX/agiRQuNxq3/9+yAG/E6dW31Oh6pPp48u9VrJUaOzj97jk1ooHITpC
7fqdFduXEl5S26ZSaDV6P8BhztlBp6ZO/DYaKT48BvMRNb9wC7R/ac4pzb+x/x+j
rXs+9tiIz7dP7nDKGNgQCaAjp6En4ar3BvmnFUETD9CX1VvoLeQ7QISOiM+2y40f
1KNEt90Fyabp4VicXbSgmbxnCkkleqv81wuixwbSy120G+orWKzu8o1V+WXcZzSE
IUb5kABUWJCZ5oYpTEsaunBeh+F9fPj54Ag6cxLfaFRqwNc50L6hUJz+FjkwIbp9
AKgDB7XjdmbF+CaNgdHEHynYFsfVlfgOeP77UUN5ppxWxWmzmO7wvRGwGoVRdEkY
oDAglpgJotPzLCRNfYFkqFsyNJTvaV4P3TwCjLhJXQ0t58Ay+5p2maSumO6PGLPQ
PcCMcw6GKniJd/VXShPspeD+//ZtfhUzxq0Cu56lDCNqU+nIFNuEq9JejR1SnD0X
+yWJ9wWfgMDWKq0PklIuk2e164mmM6GiOdN5B5H40h7jphm79OfLeV1Dr1wqXMY/
Jqp8AE29UY/8kU9UnsPRweJpoSd1WOWlKLDnYkBno79IgiUgjza76Xs7O6EAaQAy
jOwYL4M3kbagSYG8sn9n5SEgMIXXG0LvD63C6x5+q7VLHZACIAEwTEXPVJr83CzK
TXQs55gCPo7k1kVEghSde0k8SVxQegJkszMBPjm8Dia593Ufxj1YwzZOCcSupK2n
YyRPg6yBCwOUxwlKdQ71EMyZN6yM6sRb3EZ6WmEH9gdRcMXb4yM6VgntdV9Eit4U
xVeodkMcY+Jx74ZjpHnwUR8HfVMAUJ7lx3RkpGL/UiM/Fyfey6OVadyXkTUppKsp
W6Qk+M/gkmBHaTggIlKbW8i7RaNEgl9wOi0TBvJi4Y/0PwVvkgZv5xpKdWWziW1p
Ayauri4N6I72jaSoPXVpkgSok3wkwe2NTNnVPpbJuj1kBxuVafaRkugL806x+2J3
ixHAHN4ZpCXzcUjcfwqeYm+VKltKYUG42+vbe0bI4lWkIdRIc7X1eM7HLFCNc3xG
brw5atAhNgAYczemPMGyK25FWIce4SJe9bHAIRlKCex2F6Yc9JYg2d+bRy063g5q
RF7eCN4ykePDVxNxlxdv1VefpO+XMtEQJmjlt+2/8B6GMzj+9900181BQa7G64nV
nwqZprVi2Q5emtMBHRKHARsO9zrAUCj26H14vRtJniSRBIfCpN6JSPSKm/UCzA5P
fOqMUs8IcQ/ype6VnOYN1qTAwqsr3nIpQzxOxMva9YNky+F4JGIpKz6Yc21kOU47
f/kKXqnQBQsi7AJ+DswkaJGEUF1eW3eZTXIiCooGtaEvw8qDRg7g5eA7ljD4jwmh
iTaq2Vv9Qj+NPFWzNad8fycWK2weTjrtuUNzeH01KV2mL5+5vOCAMtkIAcP1J8W7
t+5SAqbATxupuBUtaCgoXDvQvAylB/CjcLxPP4JDtwvw+n8pqJ8EAaj4LldKNXM6
Dy0K4J6yI0uxZT+uj7b5FZq1GlpHa7BZn5iooYIgnnXkxI03ro8KpSKnSia/PmaA
h09zL14zOX6BbFbXoYaDauXF21WWutEOxGxMAfaGQZgbvlQZ4UYOE4QOmbHH//mu
RhaBrPYWERRl12Sd5jviyo4bT8Zq0Ak0zDbrMApIfxHXVr7eavVb2VGMl/XTHtTc
QV0EbMYlrz/wL+U1X1EjzH74dl+ttPFVzASmWiH0aRzM9KytBr6ZCLoVOOF92mRU
5YDaigDPsYybf2ayJ5dsCDIoWCF4bYQqUB8IJeR/HdC05bJAaPnvEsEkYYqDpY6N
n5dk6zvscjBraqXe6Zg6l4ZzA5T/zPMZ4YZqKUH8VIl65/3r/+LYfX4PAaK97rNY
/r8K9wkQovC0asJEwe2AmGobBcmGWZItfDBiAy/KpdVETu6xotcfGYycPbyMrf5j
SDO8W6M5pFbbaAMt0wGVAlIlo7wUrILFVhir3N9EqOkUl/CkmxF4xDQlJeJs4A8X
fbVWIKa6/fUpzmWI6JLLy3kCIYvDaEj5Or0U1tmCA17rXLcvBpu3zbZN7Hl1Cl+I
seGAc07L7CD/yZt7xdfUUaR125wTqc40aZ4wbCfT1/E2L6JHH5/c4dvPqz5c3tcK
qJaguBpFYZPP+rcpdwHlz7kNPwg8EGYmdHAjYaegDHDnAlHYWHgPsjjYA2YYPc3N
+srs4ohn8+Y0ThhJbcJphxIp93isilMCC+4jbEA16SIWOWnZjZlUpevVpsuc/B8X
zsF589QCwAmLxx0uiHRCwvQ00LbGqDd45TJgcYo6bNHPNER+z4/cEnL/gKJ79S/Q
CK00HBlceweuwvVjhMf4KlK+2NoC8huEcGbDAiXduE91SkR2A34e0PR0Q7gKyIQT
X6iFD38NC0dqZ1vIhgfegZIypoOh4tL+JjsugiCYD7XzFfIBVLeqAjTrMa4/dLXU
F0VTr4EOwu40jYdAsTHAArWkIGaHbOg/l9XS39OMojgX1j9pcexjLvdkazwuI6Z+
apBYxtt7h7ABMzSnl9VSgePNEu92ZXE4saiEWP7IZ3Jq0lnQf1kB4LUyTxoK+B8L
5YKZTIQKgQJ/iNMUkmOmDywNxFcmueGwATQZFi+qF/WYtxd8h4p/stO905i4OE+V
lIUpMeYLnmmgrY0SJPKtWHR4qw/tc5lCfCwqHq09+6sY9067fHn5eDcqoNPovRjU
1mEHdwfgLj/ZuMiPj8sEB+YYakP3HX2eZ07BuMFsOW0Xyl9Hfgn5cfVu/6K2bcVZ
k52egxpYjT7HyAM9zXFsQ7hNAmlz4QRrthHGyVJ5/utEY3joar7bdtDzFe2xU6mN
BTl8L85lq4t5Y2W67qirytkH8hyoZ0lM4gCVbgbGySG8nJKRa4UlWsI1NgKUf4Am
hxQvi8XLWyMRkGyFQq8Tx4RAxXOi2HvxVtskChxdO9Qf6U2tqW+3aRmiV10OqrRY
Er6LwD5bGmn/YftEE3C3uKhSiBTfbUowRrFW8yrGry5W+ViR+h7fSogss93nyGkV
yZDNVe+Vj7asuBf5lzB8EJAWe/76wRRat+jPFLW7OagZKbyDyNhvCH3sq93i4EH8
mHOO11LYxGiCWliqohE3/K7hn73OJeLTlvjjInA0TZjz7oe8tQ6aN+f6xM2EDtQa
VJs28/RpQiQkQwnh96LfmOJc0D0wJvajg2Ykck8CX1cBXjUxtz+yQaqPiRHQYZci
8wJGfXYnVqbTTVUlJCSo+iBBfEhhnotGqhPoUkkMkD7awh/6+AKJjECv8S/FaZHW
Hx6jxjrsM6iEvjDDCaymnFpzY8FiMykLUTX3gBlkLdElTXpArvuRSFgVZvwSCoKP
93sFVjBrn3krtEzS0DL81BR//LKnzMp0kHKzWK4P+kj8WDSy1d49oDxRVPEZMBW9
GY3FtDzosygxj3dc9Ce5/kugiOo7WtjjmRGzaIDRr7N7+HNn3/VYpIMDdAwnG8/o
9KWUVNPanKYCJxGGasKMC7ElS3dnLJTmyMq5tfRgmjsomXrWhThIzwlWw4i6ciRk
0KlLorLmoUpcuZnkvFcR8TRqOLy7zyM51SckXcsTXPGolh5DWjQLEB4YrG0Wn/Mn
r3ZNez6u86cJgAwdtwMIzHUjk9uErPCHia9lkdGmfQZuQ+1/LMvUYCRZvPJlgvnZ
r9nZNYmJ5KrU5vWD6L+Yrg9sf+aAU9am5BXegzjQoKLMJwY1iNLJ+2ZDbsdSklHN
A9vhWzXNmLp7ffPtmHl30xDkGX9C+GMJpmbLb2vf/BvlPoJxEi/1SA2TGb8CPfG/
nJ4Sv782mXqXyyL7nQ13SPxR1PpKdcRyINnSxykgqbNZiN0mUIzYIcIPSTF8T+UL
dsbTrF7cmOZB6gcjuwslqP+ALAd2bUGJF7RhmWn2uo7nlZcF+GggZ/f5oBucpvMS
xKO8rqyEz7hMUSu2TWa2MmTYGJpaui9hHmuScLV651TK5VfKzqvMViPMq191OPW5
b9byqJLgVJNHuTwFeGtpIP/5hc0PpTQ2OeTeZx2tso0UMN1wUbwp4pFZV1S+UsvL
DNGHQtqjKZT2gbdhiZulGl665RcDpyLIn7IMuc23UeTEdkF9R5tXBMp+DkpMq90/
x6xx/N2qYfRVLjK8x3cX/mHGntPSqliaq8xqGHbkvtF85tXhso0+HT3am2Q8I/YC
1reRAjlycNL261Dq8+T3AGvglu5JDGZqHTGpkNm2INxMgWsMMvCsnfTAvIwFMd24
tnq1yrx9RPpcG8Y2B+Yu58tXcz4IoUg1gTkzfmGsPCdcDTj5mP+JNfek9oBhkyg3
ihm5IYLPtQLMn4xiBmwJsLbZ91HkJ0oM4crgLS7DHNWxXMo3B+mJgTmvTBomUPB2
M8nJeXdkbaA9/cEH620+wgqMXtqs7ZzKZS2J/9ee2N7T0G1d0wlb7DOgi2Bcc0aM
dqdwT0KLcQLmsrTVbQTHN/LSgNYVfsJ83Fhpw742GZF8X4aVPnT0W0dp8kV0PEuS
8Ns2eXqHReYpctWs/t/fjwVlliig9LEqilCykKKBVB8Qf4IOU7+nN7nMYWLNjh5d
/n+VsJyS/jjjpsYiCrfklNvSrqkCDu1nzNyRwIDycXFdPlmjEwQZcjuXsk+fHDKi
dTYF8d0DjWg1re9cvbg+czjYa6n6R32uiPn0xd7rkMbji34jo+jMWaMYF1FlHUQo
Ju2tNAuiyZ7PzRbsXeUaITyeYdvpCL9n8yfOIEXRMhhpDIfLkkyiXoWoCjobPtAa
bLDpHVqhgmhgWUM/pnTlwStnFqDqFLdoaSUF8P1iZIFBrK/xf2fBLjU6R6Pw1kcM
NKVrg/qP2eHlzIQy0mJlp7G7hkHJL26MvPBRizVMpBXQ4maypSN7DQRs4Bc/9RnB
RR69QMXXttOgTOCvmUNZx3cpvVmQGl/L773dQVMLq/VcnNmPDAFdxqp9CK5IbWah
pdMeW3RbJ2xgmcc+FufTJuY2h6jUDLLzUDN9JvD5VXryQtHM3b1N9p66v39K8juY
tl8OVQcnsLjwuUDFwOH7SEgLeREtFCEKVE0ms87fpAvB2RkpFialLkrd7dA2BLvq
IV94ZkXwM9XxQaCo3C2LS8YPR1oE09yIStjGfIUj4guzZCbL0UHudQpkgcO10I5y
sin7ikQKhkLT9sGoWBhc0LAtS+XL2iRAFY+s+P3UT2eV69h3fsIQZNvr/3b+TjfD
f1mUS2tJi21iYiKx8spV+O00cBehhegUl0YX2/QZW0tHZAsPoJi1I9GQb1pMJWzt
Eh0UYut48vxp5UyMZoqTWrGs9hpFnbyCc/hkxCUdMbcLsPNDktitv7t7u5k4TTOs
YRY2u0zNdxRZl2r59ONYpmxfC+8rURqnprg19kcGADAmdVf5RX7UUKBTNjXd1oeL
XrrjypycIdBjuldNpEp4b3ZTcupF26YuTGy0wkrpjdbLEtkUpK6plMVfXuoohuj9
4rZiPfzA8r9mjIcgJmB9w6sUSobD2j7ntGLZ0d9ZWelaypKwNZ3ht96g99zN/cyG
Iz5i9O4g/DmXx2M09jksxSiAyBFNcR6ShVg1nce8qnFFFZZbpDZMrV9JtJbv/HQr
J4/opAsg46rUbOFILBxvJBAwXdE0qv3IYf9/bZygaoZ1OHzo5yJTrsY2HOSOyS2m
hQ5xot0Z2ON5h7iwFPpbiMEUcF+dEIpp1y/iyv503oNykcA5WI1eMwJiygRkR6DO
Pphda3o44rws9gKpDzWORd+MGYsjfoROl5jnOYxy/17D1Mdl+gGCdtHD+EiPsi/B
3wntjU9/XaCydGMUmMBz092dDZYxkOa9KxyVfBmVNlweDEIaRrlTvW8tOE3X/DFZ
Z1tDNGTzDV0blleEQjBeu0L+qtDbGANJWPARt8lzpevik38oULv5rVxpqoaJF5D+
jcCguNcWCy0tlgxuLSm9bkfa4Jh7CeslnqGSS6CfxspmIwF+ZfrqQ7sz+Hc4cVHa
Wtt7jCDyGKJHW19E3+Ixn4IJ+usJjJVYoK9E6mwHWuvijGPy4R+5pUHQvr93iw/0
FPtqTMQ5WTxtWEokoUieigtl43t5D04sK/vDbTF2XC2Mgnm2RjDaH/FMsBfxAcST
R8R8T/E/p9I8uezYcGC1KR/44JC5/clZwWPs9NarVXeCAKcUvB7EJ4DKn/wU98qL
AVV3bodn6KRmyd1V+krRqB5wizJAB4CL9L+JY8OJe4S8/aZjpLCXrU393sKgasJC
nwZW9w0WnldTiX0N63HZN0O4AXH54ikEeNjpSsvbdO7hv/oPDNCZLBO006+uAPik
U8GhL2Tm3BeePhIc/QRhkZyC2vc63FZHVmZKAupm2eJ1cruE6tCV+8Ox5BL6I9DX
WXG8XJ6UQdP+ULPr+48cLgI009TBmOv27+lbZ6/4Xul4pyTuCSHhV3MrLjI3PajC
gGxxpypw+2Igb/2WG7K/IetV+/DdFcUs2gGJ1O42mMf4w0rlklKU7CcqA34sbMDa
p0HRsi8BhoRnByxYfpOw+i6LPHC/rxq5TPrgs4oG0zfDV7OeiWVL1KVmiEQZsl3G
nSKfjEYV/O4Zle37hu85qf1M4l/ca7g4tASiyYB34Yq/YZk/yQwCbSbvSoQdmBY1
Ej5/GIg6R3EBdl9AWjF7zm27bvbbyNvt3sHPSrlAtZyIfXFRm6YJiAcWXPE7tqd5
Jr8D/S5Oa5xfwuIllKkkIvKeKS7aC8kuXXb5QsLT+AD+cfWwN8VxW6D0A64KqSDi
0nKyPwtkJ/p/lQlW5sBicSRoXV2IiacZ8zJhDzOwofrFnCUYu3z2hdSNKOl09HEZ
u5DW/W4QlZ0uylR0cgthPYLqlPSb3LXowX9DaN4hFv/qPJWiGRBu5JXIGQRKm+HN
tpCjNIhQwTiwhdQTujjCNqJX55c4MVeph8wf+5MPqSeJUWjQQ99+81d4a+ths9tj
A6vCPL1IxAa4MVgYkP42ACreNxGReQ8h+JxU91QysId1gmF9LEEVhSwPDgDvlW7E
nBYuRulouZD0+kho6WFfoPWAGrjEQgUHHhdXWsA/4p3CfyqJ6ZZHN5eC1Ntn/RbH
QObxRPvhsj6y9XhwF0aeT5B222Vmqgv/+f8gad8s0Ql6/SHkyyPpkijX4fgsBkSQ
PUZnSDj029Hw7kuTvR9EYy3Y6iR1HtCYcX+q72lMDhLHUhhfTkYfe/is3f+gKtEX
YmtX9Ui4+sXAkHRXUIlGnTmFa9flK+i46HoVjXoK7leOPUJKwVpG94RBbZpTjG+F
mMf9ZJO7hZz0CX+BKMfmsLD1AnMQA1t0urCoKU/QSiQlMs9Ij/vyUE/ucwi2fTG1
ezSvvM0bjtnE6r9sT7Wjm7p7Sz/EdTqwbcEBopOlCNT2mhuK2hzzNEfY5T8Km9wr
mPwsnqu1F6kwhwH6OB5QrAZWyrA1XT0GglVa+nLIDsq0w3O0/fmp4tknp+H3Ne3s
leq9aXcSsHi+zVslpHoA4CKAC4dQi5Vx2XossoRrEpBrMbGoxa3aMvnBn+LEBHhS
KeEiMyTXcsGTmLbRdBi9PHYqK+cky5S/011mKsNcq2OBkvfw5eHJ0DUta8G4wiFv
AlDxl+a4psQvlxF2eJzgBvwC/y5+eRayJ90jdyb2VqLIP8JU19sovCXXRkRvT30f
8nPHoVGC1Hg4NfuNGEyoHS1HvBI+v4NCBIFiL8yqavxDqcTttoIOOvf34V95Qx9z
gpUSPug2S8wFN1SB1GLnfM6iCslBN9y0UZy+oARe9ul2XnIUqNlKJJAsAqXDsizC
uKNaAi14A2W2REtWYtGLi087BHDbjLsUnILF3dtDxvisXLkVgvRzmN8vOJPooRtZ
1FVmAikjtwNZlSMPr6K3yFo49MFt63mQEclKg6ublzgwydE8Dz3+Qo/px0rbidCD
BGwYbS97b3tztM/BDAc6r5ch0HCeMZ0WAQ/GyoI7LVVS7NeCjRb2BxWEiWr5vfy2
648uG6F56lpHFWp0xLJ97GNb0Fbf+8yzTy2zzZpdQNCFnvMsPOTacILNgxPEfs5J
DA61T+MHwUTayzC8g1R1Dbf/jQRZPvgp5SNLvonfC4un9QfPZxK5X32vdlOxhVJH
zZJQL378Sp3khuj0ddLOfITiniGvsf7RXUPuCMPsw2bNq2FVe4lQUNkZYQrmAqcu
JfGEJ4HexDHditIxUbO9d205xm9H+WtBP89gHd7E4H5K+9iQrdc/Krn703CFrj0r
EvMqv5V4NcskK2dgM5fSB2rcIYb56vFjRqIET9oxnuQra5S4mNfX/mdlaP12Yma0
ecknp4GdCQqL7ftQZYLLUia2SvqybQvx4JKETCwbR/20Sd0vkdFejYtGVfXEgTZP
sS23wAog96sKhDwoQ8JaqG6FdTD/++zVVy8vE/Tsc+aFjwZ7v9bP5U4RRLV2hIPR
PR5p/+4/lJ62nmGOqvCe8aKBiDo+KWjnW5mRZk/fwfbt8xqkgjteNOjOyDr1dqqi
fYKCrV5Nd2W6TK5hYGSqNoLL97ZTuafOyr6DAHg2qLaozmTw+gSizh9/MmiE0upw
jHCVl8By0SRTUXjcNvyIzXMzeMb5WpkzlQzYsYMHW8V7J1froVtgAvrKd1IKAi7X
mKJe3yLe6ycwqwd/Fjq7BzhpnUYZkbwYuVoAso0+BN/IGNBK4xZOscpspevXSp5R
QtwlqNuUsQLBaO6bcSQUTBFreKVCByaxS8Fcbd4zZ3lcb48ee1uwIIbhf5wm6JfA
P+KEYkYnOLKmHDXseyQXE+wfu7Xb1VmypVO+y796uxkH+cvHuTBLQEVIAX8c9PCq
bFF/NOcYj1DYBepn9NpYuWBs7XmxicvHpxGpGcVzuQR+5AENoPBnYENCOWzyC0dO
xOf+R3Y5CcTtE7nm6YpZ9FPTY64zvcuEab0Necff2vS3wKEPe/GzxQiSaMUbkxFe
/GoU5Ezxz0tZhwPnjin8CKO11yQXucF8qWQFsa7Bs5gEToM2I+xULS5ENCYRUf64
zZQb0I371FlatHAtxFdlN7J1AVwU1UyHKI4mfkhI5iG44iaeRAqCpWciCE1F2eCa
J3oEY6PQ6n+0Zcf383naDtigG2gxvBKIxaDHvHT5Yem+noEkNNncXuGKu2xyXgPV
afXsZheuc5O0ioVlu/Y5OJvDZ5+xlDPm5n98rOCKfySCPrfg8yq4lhtsZmctmgku
/EODMfRy4rfFJ26KjPCfVJoAiW3ycMV7jyexsP/+WTHaCRqZv3KQ6DT2GRec5eOL
NdNscqdqcFm6nt8P+y/uZaMc4zyBhZ8xcqzX5E2HvwWoeqvo5CMtDJHZcl+7bfVs
5ip72N66mcw/CaQ2xIKqw6+uCOQ9ZEfhSYEP/9jc26r/PDugTVQBZX4ZZ0ntgyZ9
FC135FIrLUM8AGc5CUVk7mLF4+2ZYgafyUCqgp+6cd+LqBtneg0Yo2zlanLeM71k
/69AZqEq9el7G4siFFIDS/jpaqAYYvxemLJChi5RVyntfrVzxAV7GDuy/RKL+U1R
tJfJL/jrVYfI0PIu6fTSFrzlN6fzc1hn1J+KcMvI+MsqtAz1ANxLTbYKHuzriUB+
EVwk+1z8sBbxccfbP6s36LHViHPYD1fq8NlwC/+I5mU8PuE6qtQOMeH/XyXXmbqi
s3ZPlQYOR8n7N6ePDNAtJTVdtnv7ZX02/4ySvceBO6ER6Nl7SpxfYhCzRORfcZec
HboOA0g41RhW6jQLlnLNLt/e5xuPzv1VXAYHi45lse2Jbon3OHgQnHdl1w0YIVii
ogKsm26s/BT883PyZCu+h+9AxK8OgG3GO5sG5IYH484zkASYfdGDP/+6f/+Lxpcy
vIrSevkRN0dLLtpcoM3eqiBj0X9OkbfB0i8ad6KI8A63Cr9eM1V2fs7B8IlwUIyT
R2APs0+mHDsHwsqBCjffH5rK0SUOq7iJoj/zcvYAXmrqpoTScqFmIZoEhSyumz5l
gxwWXEJYRKgrbDbOPExuHdSH4QpvEe3rMpUSwyuIoaE5pzmP+W9ivScrPXUY33e1
Sh4aofO4moafRH65iikLGdjRx6iwy3sPwd7A/XhH/twUyVs9lNxlDMPc4ijUFQMZ
UVw/Him08EXp9L3JAXHZBz1y0HazUS/UbC+I9T6xYbmjx4mDCpgtpOpWFhGFCkcN
q72vVP6j5hxlmhEE+bc/Znx1OeHqWhqfiDmjesc0NG10ebJ/FasqO58z/UlHFgDW
TFPx2Fek4Y0DLeNPwpYsEPKFD6V+8cqB8+eYFNV0+hnXmB8c43TKU/JN1TNpKQiA
lhalU92HXvFtsFqPyOj0TR3oMcU9QW6rfH6c4yGlzB/epR3XkEeJQeH5OueWZpm/
+zjhUNKSLrB7c4C2aIh+lB1OiloXexEFMCZFhD5KRsshNSOu87wGF3OJnluNnz5u
keSrBFhlFMODF2kF2vf6OJubqkCZoG9XW+tWHxBlfZOxjIjtVenDisyvwq9fysYF
v+tViUgIfG0jB5ghuIAxzM0OqRoldIXSdM4STFD5OwwssdsxeRlRgriqpCrfKRYX
KbKcr8BSFVV7p2QtkouP8I+CQ0qM27Gzuq0gGyPwbjSgm4sm6+yS9mx+YdywOuLb
2pLZJ9NRJ2wCfP7BOTdqw3WadjQ9Bqu+HNaKLvqdBa0ZK3i5hj9cXkEBGAQQdQ64
2ZuKLuSVzaDKkRdqfr9RKbMLSNAaW1RWFZ2qD0Nz9eBhF/Mh751YftI+QQgFDDRW
ZRXBuMgYkmCLB6FB8vva7GZyWgxNfZzoWzTK4aD3i2mXbN75GXHItG3XnGH0SsEy
+mxicQ0loP6fKxRXxHd961LVb+hKsqGztiVWh5vtw6FHC4upm5ccZ0YWTeqwWfTi
m5wK+zogG85Itf5w1uBcSsNBs223t8AGKhA8ENkWvj0PmyaePhGK+q2HPiUWgjZa
dv5DrUeTt47jpI2b+/zxmlnUyfuz5AufXPnSz3UlfZexz63YT2qqhoc/7r3PTIN2
gGSvMUJqiVNEeFBkbxJ5QlT81Ch/7ElN+2HxbUohFldGV+CUj2YU86BPzqZVlvvf
DiliGpFZbWjMgghcyvsmMWFPB0f2kZ1uo/7sjdSpHS/KO1FY246PeFbAbPAaY71o
xcDCio4rbXAitAFx4HGBeSFOqXuWSxyVlzTGhWn6uUB6JM5OP2p5KKhZBZ0K7XOL
2EBlYpQrwl/rY1zKXbV6b1Z0/rPuQF9NRtF1Nv1+FUCWlWH2arZ6JTw5D/iJvzld
C1oa3DC2cCRaGBABtUw5HhWhOf6gF2GuyFA5dcR81W15/DUwcQcq8R/tXtFWDCEL
1LWZtkrLnKelvL3mOdSVyKzJzBbYDPFWBsWGEgnVivlYoIBiHNQGl1BGRUywxD7T
uLVceXRVXTWkoN+QNVbCLXblAZcwZ3Ope2z/2a3/UdZl5Igg+lUz5rP4AC36CKMm
GAsdXHWmM2HhxkD9EFeZUPFPTKiG0Zufq4PCJMXHbhIpsYNnsXcEg3XBNKw0FKOT
xcEcKUD4zd6Mwza5j8xvRc+0mfOd9Ya2jvQ9MATxFg/wPHXuNuhEc74xpFwrJRkg
sYdZwwo9amC3gkURKpwLZPLMEsvNPNOm+/FkZXMGr3VOwPanDrzklqlhw5FUuDaR
McUHHAjyHFimflFd0u9zbF2oRCXqbLpaxE+ErVwqYuogPE85+fXKk1YzsnpiLrVO
Ddq44Xhq8kcRbytj1BELHI4KCwPhvzEX36YBM6Mt2KMEA98nH2rrgZs5eS8kFSii
DljcG5+DY2ZMevrQF1Fcy7soesONlLgtlw9DBhXSqSFLiQUz1D5W1RKv2EN9qqTR
qomLGwemeTm0sEGMNmTIFUZ8Cf50u775pOiGXnCAJqM1u9reR9txRP92oFhvMhD9
8y9bhveESalBKYayB8EoiF5Zlq/jC8ihggRbi6GNkg9h7dlo3GWnGfWz+23qgUKv
tSmlZXhTdPiMuDblq57o7F0Xvg4VC5n+5fKlmEdIl4X3IIH9n9PbEnDu0vSw1bJw
rnmfUznW5USK1TsnN2UsF5HOLfzHk8638eAUNT78j6UrMV5V6EHiXt2wmrYEicPd
UzayhNHFEaRXdrXuuATocACuptFjurrA6mEKiVN2X1In5AL08yjRHMvYlTvOuiQv
JuPY/lo1isU+pM+88xF2coYg6XeuftQgOMK1GNt9+c9Eh+Kaet8KnQmYRzqvmiJf
IH/2vyIIjVcyXO4qzOHOS+IxHs6CNP6C2DnFSPHntwoEJjeN++DMptaxF2HEFvY9
eMsuVbFeidiMOaW+w9Fgh454wjtdHjbx2Mp68RYsuhdNuNNRLj2GIbadiXwbM8nH
WkhEGnsfHVnjoGll3SciPKR3n8yaSEFZzh4b0xSOOks5HvbYFpjJFHxa4uN7QL7I
V926qK9/EoqoYsWtrFa91Uvq9eCAJ2DGWi++nJzVw8h7BiSBO6QXG2B4Xz/sOoYd
7BOUsFmLitN1BAXyIr5bevWsHgvi99mF403eFkhYDoMErDmWD/Z8fbV3JK5Q+eO5
eqwxUvRJSt2JXwn7RCk69+kH6VPlrdhnDJc+QYzAwIlhyW//yDQyH9psbJEJFB0v
3Oy7qZI5gpzXDU2RKLXzfqn5Tu9Ehj+6/n9Kl15/A4v7OM+gBYo72GYBg/rxVh9U
O3Q/8UosXLM+IxIeBsVXxM9fKwm+wlRRHALJ8L6r1n9vyWQ9WdD7BXeq0vaVIzUw
scUb4pV6KEHHC53d/ixAJikaKRuIeiIozcBnq/BMM8LuC9XRqRIUe70RlPemu7u3
xFA8rFejdPGHXO4xOE66tlUwGkRCMcnIlP8XROlePmYy2ihR0vL1rYmAh9SJJjd9
4bQJPWn8o0xe1s4b6CWO7Qr4l/563GrIqbq2AeEUcxircRed7qn1a4/06+TriKNz
FQAvF1C26fZupUWdMiff6TcRV3WygMf1nZTv6ji9scHZZ90zwvS7gHFE+zu2zYYh
/eLezdVCwJXpsDLg51qkXu9PIbqHq071qCH3YPjgYVm/zpG8saHvQYuIvyL9Euhw
wfBtPNw9VOXg8xjRTxJntnpv9e++lQFll/EXUsb+Ch/SP0Mq1FnuJ3QhoUjA+Nxn
BEoCxTxEBgIObLG6hssx4gumrqJQKVI920sIEbIrD5K5I4tbTGa/GY8oSxjfKV7Y
LyDlJ+Ir1jcoNe2MQUZVLAxGD7L/uGAodRJCpEScqzH5WYnxgnrSONbsAqtNYtAn
qItVn262xsEBU5OUhfr0vZljKKwRRhpwSb1ghbPBNowAad4ht+R+AfDWMnhJeaU7
srE7Yc2kF1nbfjNV/v2GpUvZhTrppHjMGHS8w7S5q46z/p/x6+pD8DXcYQlzwwkh
ixPJDyzto5lxGVZS4QlDJiPN2Xo+7IIt+odlcUpPT9Sefh29D614+1YFPtF8CXMv
CtGG9fmAqmlscyzsMOuAOYWKFYug9VGqZ1e+jRhuHGe0gNXhggRovRXcbWrBEUxx
2MnkEcGfhOcI+hwbzS1ezn3onUFmLqq8ZP62LAu7CZa3Mrz3zD/fBC4DffIUziDI
nqcL9jqC+UE7/HsrCH61Cp5+si8OWvQ/EM/AkNzFaV9f3XnOjh2qBLp4AeEkzhQj
rbV9XVHygg7s/npkKqlBsfGbKWoYiBSVVC2wSRh0OhneGEIaAdIRnBqB3Gr+XGCK
H7dnlOQdWiz49yytU7L00wUqg3Xfgavz5o/sajB8t1MpF/Ov/lfbhSv5LR90Cj39
M7ej3nesqifshlLlHjL4wYoQG7w1Re2aSS48vavzMjhg2GyREEdpz30BWlA0rZhi
mxjkm3cjmqTZVmtFoVBZAKYohdIMiPuBJwEcZPFCVBUM+Tb7q+YE/Xgh00cs3xMl
DaqgabkEZvGhoMsUoU6KprJZMzcwgrkdbuIka1ioEm4pphvk7m5Br6UD9ktp+lOb
3YF8CMyn4+ltCo6/1S+lE3MPIt7XZE9YqlSeIr8UF7oobFtNV99DsEuQBsTigQFw
JIS67kZIUgdR/Utj6JMSxv1P3mya7Ie0iLbBvITUWgM2hBT+rhx+Y6oOjpcB3vCX
SnGmxWiJee8SKnmy6BQmwbmoYuiGXiOv8QyfKy3pfGMtTVp9s/4hcsFfJA8LnUfi
RueXTv7Qz/+n1TMomUptjug2WJBP1d/FXx22Z5Ai/cZZnbOaMif+hnsqiZpUXHCZ
0bUJ+uicCZMC+jRh/91huhwLZhNqLDI5Sss0NXOg2B1cAk+nEpYDG4IakxE5QRnE
Lq8IQqCSQmctf4RiHB+87mKw2kDgWLtRHjA9fRlUYwdBQOg9c5H3RUekSCTAaUPD
C2kpMnEkDzeNwdr6ijkaBMDXzgOXqQOsZ8vAwSIrk3MDiOp56fv4xkmd4ctiEoMQ
nzGADfvgSxXdi6vSYCAZcQ8I77a50tO+Jixdxag5DqxNe/oQ+g9XAzEJzo1JDYIa
R5J/w6OS57gRGyW0T18+Jm5aSH551vH1C+EbWETgJ9UZ931DVrP/FbP+ai37zcM2
8lxQMD6OK2v+HzmrBGCxL9IVyse4bPn8yhgRlfSH/CAcWspqlxj58OQvCqHMBXwR
fUylrX8XNpZ7r771G4YZMmUHde4XCF7WoHGONBi11Xbk9Yo6LkyJY2om5YztBF04
EAybei6xn8Xv8I+dWi3eSGYFyw4SwciuA+EvNLcljfRufaWI1yMVrn7fIpQBcmmI
lt/XedJDD21XeJeb2831iU9kr+FxMUE2UwaSxqStghAH9BXtugzRJHaLxm+/Lcii
RqUqdvkpuGygDU9fGIhGXNf9dZlPC38nvuuIgaWQ+c5E4cXYQE8MOAcMfpIuoSw8
rBh8QTKPrN6LG+XtVawnkYPqvN7Q+YwqJX5HYMBXGrtdKeCMPFSVWws/U/rvV4/k
iDSn/J4ljdgviYlJRvLgAWw3GZCB+VWzv8WndDiXi5kWcezwYEiW7seB45T0WS8+
VFxeidjMpDKG3aCZfO3FXj5g0uf9Q/CUkvWn4rQUaStU05ZL1Wx66Ie/Te149gzu
BIq55WVXzsEOCzK9mDW8e1Rrm0Xgz7IM/vpu8YLkh9fL82RLziO++82dEyweILUO
KEmVGA97sGMlxipQTltPr9qrx72tMBogexat8z0hZFZ6+HmAVTwNzVlGNqMwX7Nn
WDsPen//0JB6t/VZhMaEPEYePZyVaUMr98aCBC3hxg6TMTHeu46OHx+FswbxMF38
XmZfuv508r48koCtt1taxsKkh4ugAAq9E+B0RYLzyyk+wODMoyC7U2jg1jQ5drjG
93G+E16MD6I/PtW1KBCb45P7btDaYQpLvj6Y2s/DRi0MzYRogcxmGWd5fhKeGTSg
NdRlbcGH3trj1m/GdEcb4g/ZDuVMoPCvHz22QpDCZfACuq5M9wD+0kG/cDYrSvjg
yayRdU/g5PJrgYkhnIDVpGoS/j+cUJunSJOVuO4m5vnMqqoSdZz0cltNAtn1zSsk
s4JDEus4nqXBF1CxUkLnfMsL/79sOSprHFKRZ1jsnDkumYudexOwadzXru8sAbqH
N64u4nR4bP9czIIEWAWDac487vD1I21dc4ixHEOXxyaEx3OVWEWrVVVhYiMg3QdS
OnJLO7mapt2cNapNnLUlRUcE4fBZjtTfLN0AolXdicY4uFVRortqyCFcA9eHXDMs
hwhh+FNqTtC7z1NzOZy6TrODDAcotEq+l+LgAJlvKyCu3S94htwrx6oggJ8z77tu
9ziOt812KeKr04p3GXpU/WO22+qz5C/mKqgE9qFDWFl7RbjHvgWdeYwhKa8RBoIn
m+in1NWDCUbES7ZOZVAwQvNw3OUZ7CpXPKGP/uRzjhQ/HA4D9rUrzu1ZrgQ09q+K
DyZPpbh6fycL7cc5V6Q4Kiys065Hkp2RlKcYuRQQtvnJnYwhX0yYx7vwRRvHV5aQ
hP2uZcxfiCCTegcJeJ96ThDoQdY9IXrnsWzFN5SnxfcftpdOoLCbe2WZS5UvtJDL
aB2JrKlCrYk7ZbCwYxHGhoCFtJUmGecJzPSE51cLzg/2bIFpRUGrL6+3u5/P3yD6
svkfd2oqyIxxP7ipHqnXq5Hmq39IF30d9msRSDI8RCzrJ/5BdQgOh+ZDD6bYOnU1
4K90cagKU4n2aE0ssNIzFAnVC1w5QsEXCGOEKCJ7wYbYzz5T50voCTbJE6n1IKIm
y7KXprYr/jShvraNnLZzFpE6RR1yR3tpEAN2QJs1TaeMGzsHQYgmyPER4FhfqNRg
Kdrn54U1H2rQvJVBQkYiyoTFdXCjsaF7iKrWZusYXfOTTLRFMFZ1qRvt858eWRPC
D5thJd2QXpObItZG0x59SVnAOQ+UdzPbFbLaevA96sx1OKOChjTbvwJbZNdwOBob
QgU8+tcDprARuMjAWhfQnubqYCTvUtP5WNyZw4yuQm0za5g6eIMQl2awxaUuK4Lc
4EFFo/1qlGsoqcBIEDN+r1hRPzWKgzIqv7yuBZOUO1ZA3EjkxhXtLk+vaAiPFA3N
bKyN5KfP5SCRuRRiS+MzAjsR8OZnJ/n1VX/+6s8Je218ZdL2wAwfD1Ah66VH4chZ
NefKQLRoZXmR/Fz1PjJX979kSTAGyO2Sy/QEMiufGIWD5rM01VRp9/ZJBW1rbPIU
i0TThsAwi23Uo3gedVPeHulrUUmMnn3osCbHc7txlFMzCqd5NVFjhW3WC+Ed0Jc7
CdNNXwBJDxH5if8yyz923RMOPWYtwmUVJzAiRS6+oEi+k7t5KN4fb35DtFuAZRTv
+EUQ4/9KF68G/Gen6derBD4bcWSqqohRFG8reZyAM+p+p4pfszz9HME2DqeLVUlQ
zeSLTxX4beKVxEGf3w4e4rfV1pj4iAXGSoMjMcpw8xLhU8mPbAfWgyGr8sCBNKtu
pOs0CRD7GCO4xF5DdiXMTCmPkmz8QBCDlGMd3x4iM457QD9asWXpfuxH7C2ZyApe
W0oxiD4MJkMqAD+12PI6ROtg/tryeh9hyajPghZc7XBuK/Z6Hh7JlkmqDBtycdLU
CuC8n111FS1C/k5WS+2ZAWb5DpreTWBwKNecdPZfaz+JtJwh8CTibwOdZKK3fMvQ
qiDK/yaZ2XBYV7S51oXGdx8+E7F4cWqeW8aWjHMtzfop+Ej6+S9M1JX60Aw2Bm86
vB+mG3HEneC1qDjnKpc6QhAOhTbGr9N+P5XnFFzLqSt40gCXHk41qaD3G6tvF47A
qLU6OZzPBvA7EzfvOSzm/gI/ncpcy6zjAohI7cj/JnMR9IvOX8QTbUoaZo4Ol+4I
FwK/eRpxo6k1okb/xppuRGTftEF077eHa9na3h14SE5jvEx8JxKcUTTc1oQ9oZkZ
2eoSc6n7+AgtcARJyXwvC3p5VJKnrJVWCQwHuUdUiaLXQK4SbtFeqwUUe0tC+W89
3yU0q0iLZxzIaQ1fi/UcFxqX3fEkz8FqSbAqIifzAOGwGwUjqKL9lzS5OQ5LmBGO
5OpkgCVsECqMu0X76GbLi57b+4S8+lTZqEwp0TMqqdckvqzCpkHl6p/Nd1pcJ2cS
G8EXGnHYmo4ugcoC9t7vctcsKBx3gCMh0sGCk0jF5ED95rIPi2iRihO4mkHGNY4E
9WLegv/h16isQMoUYJ2E1vutK3lbfgDxuSzZI9YYY3ole+SNH3Jwj+9bhzFdqafQ
gxvLNWgZLkq9LEj6wCX57Bho5hDYSVgm8bx7pAoiV7AMShVI8qEaViQMggMn4/Wi
yHk9vlrEZjg+ycm1PsiY9BLDp7M1s1Eyz6AV80LPGgWjJkEgmPkFaW2C0yRGMv7X
xWyk5z6OoG8QNNsTcz4GyGvnBpo4IknqDaSXoFe4ZGQEZy6FmqSAAyc+/b4c4uo9
p11/9ZPdUlLzKFuIHtfvhG2OB9Km28TmTZeRfk/oER5sRoEY8qUmmVQPpLpcUeK1
nPS9HICiZmkf22t4rn52f+JK6nNgLFVqeQEM3GNztmbju1xgWmgh15X6MTbyUOqG
NpxP0P0+EDA0V8XwK9o34YlC2+dWDbz7VYeTAK6HNavhz+uzCBC5fxbH0DMEEb8z
yNlhQgRbsAdkJBlkXr/ED5VVsLCnL91VC4Lp+J9JqH9x+Sv9GcArVSHKNq8LBVRC
JQ0ToauWkeJVWl1Ps3eqEVkrKLsWXCRyVLqEt9keu3Q/ZZK5q4/Uc/O+JgCdJyt/
4PFGpfuVFMxbxtLreRPioM0bp20Nos4zRfmW2gH3DzoyTJJBag4L0pAIqJD5QIOX
89UINm3oJ5KmIJgvvqP5hUymVZyUxF7azpf33IebW401nUzgaadaAB7+ju97uU3v
lus0EkRfhC5zXXOzsFkHGUa5XQOW9JVebbkyaktOY63vuFpGHb5MbncvpEtKWTp2
GIgHgaE2kguPjIkg7rortn06g4wNf1A7dTuR7k5bmQgIEy5gvikW7h9WJH/2J7cl
FZh2xS/925Iw4OEA9tI/XXwhJGqaxr+OZegcJ8WN8I6LHbUnTuKZ0yhyKSPM1Xug
Mp3tNsNp/mHYpSkJ5eB93bIn8w9D1aPAl17g4Zz8Ub93yASEIpA7wV8d3Cx684Kg
uDI/ayAVCBOB609avHvNjoKIc937N0GnOLg19n+UcwydVmA80CxDfSsFQ3rPLyCb
slP1nBo3ir5vmKQJgCLvv2Wscu3m6llci0kmWokoqmQgPpqnV7qbz0hALWiSNYWo
hiRB8iuFFkfm+sF/vDFqmZefdEufDuk98QBM6yRkSJaWdbKdI9tA62TcuX3piir3
bJQpyUy2/K27B4tTOr2pjr/W4GJhH9VSO3NGeV+W+xQqNcAbuG3lfDjpM9HTjdqr
wMg7hj6+8g2x30lseRG4hnGG2mPUb415LYCfAVZBUGDXLlXBNFRsaz9EJMFR1sOL
TZjE+qObFXm3F75UjFiMGZjmI54kSuIh7SN/ZNAhJfc0sN6dgjTU/kU7Ng0o9Gcy
TJquvJGLqtexyWQiJP7GcYKJx96j3Ffhisi1wCXJuFZ3VHS98Y9qlEyvnHWJJsox
yYkMkkyfq1WBQhSlylelJXNrpJX5cIm7hGV/v8u/O3IxQlDTPbhEVfZRm14uzs6U
dEKrxVhQJ478AGjpgDdnstLaEldf3qkfcGCs3/jaw7xrndtT8TtCPgK+GIwYUj/w
hgo7v2mTfgeT0j9gj2SLn3afYPNzgPnzmi/UseopKibAL6rscyHBKbQVfVoItXvw
NKaA80c1PED/0VTn8t1VlrMEfjsvepQcw2m7u2jqkg1uznmG1ghrWNYY5HqpAmDq
rzQAZXwJJwWLjldxyAEoQQ/rN5KAF8vankRSOewBfHUEwCgilnmrKf80peanYI8P
KqAq9+4xqVZGr3mORQ3sdjZ4D5gdaZxsqk46Cc4w7SfQPDsAcOUZHQE+RuVGe9vB
Lts9/uO6Nnh4iSMnxOr+0x3yocwwF3OfpY3PZsAIgymeY3GA+/TORZ7mDq1rNxDy
432pkaMoWDl0naD4NtVwSQtMrRiFbCB6XX2bBWJyHvlssHNpSjctRbRGFKb69Zxg
m5FZdwMjVp3w4aDrhlroniqwlv4BQI7znmg3ljfmGoM3GnP6RgoESlmSkHk4S06H
yyaPFvFHtv6dwxLWfgTPKq6pSKqdXfKk+DnCiXgdNTlECMgdpLUiTXp284+qGSYO
c/Teqx8ufEg6OsiNr7q8QwTUHO+eT755nfEc5ebT/lRAfat5wm79M68YrvjrE9CX
v1xopmNxDiw+ux84upj7sNqe/V0O5bpKxEgkv5Wk6srk/pEMn+sP4FHthIla0+mI
Wbv2Xl79JgkIDvRM00HYaY/K8GKNkXBFL4cyMdCyqJ6j2fHgb54btxXC5PG14kF2
jiOmN8NmM+PiRTrlJRUfKFvY49Wdr1h+FUghAeEpJ0BNhLWProatW9vW1P222y55
+7iH2ZU5MwNKFaguidF2k5j9bF0sqpPEMi6nS9g1LepZMLDqcUPoWtMJSFgfbS/L
2bfZ0YLz8t545P1W6+VheLBeKeZ0Rx7ikptYOv8ceS9Nh8AhoB6AoRDSgrYm8pNz
1UJbzGD+/rZgdoDqVK/7hdVU+t0WB/EJ1EmOjZHvzAo4waZhdG5Q+oiC/yvCXwze
VxnvDRUeSQAs0oQbqbscshlxHhqklX9XshCkqnhmAb+mBBBczIKB1S53npCoKDt0
55WjLodzxRHzP6ganL6D66Tr98MgzVZ7tbEeePh8A6ZOmIF95Ki6ybVHohV2MC70
7xmpXfC/t17ehaelxiHDvrrBbEEolRFdbeuYOP7a4iolmC4b7/aA0DzbbAXY/Ps7
HUBpiq18raHkh+99jeldVwvmjLRxHvlBDbeneyQH5ahEDvKNLvZdnfhHIdFTVV4E
yRgCMslRJiywY7QsNN65chbvozfpN9vSDgLdjs1GpExML1w8n95256y6+NaCb7Rz
ik6LQ9pJATXcqZLuY3bGhwtBdZeiMlhMC6icd1E7jJlYKf4jeRmjqzgDx8Ia6mKf
8MhcDRpq2T3DFapwr0Y/H18z0xW6ocLerkJMHu6rkzsT9SM3R10EU+Ea6lbH3K4/
kvILJ8BwwS5D2aVjwLAMk8yfiIiT0Zz3drcbbpbSzQspFPCNfhHIOs6HeBuIdV76
o3NAKWDwMy5oewBCCFVf/fqAPzvB6NZOeTTd5C3YBkbJtT92nj5gZmXZ1rZQMa4R
i2N8w/LeC+HmREZDkjibFu5CcGLQ0MFaLZgQA2LBHUrFkBE5MnUn5G6qijkxhVxM
fLGnF/VuVe4TGBmZQWa7mtcqO9+LLhUp/W+v8b96Mb5o2+ACqa/Ayh66ftXt0qjP
HbPXI7/ImhlxAKQ90DApBbK83xqoQcjHZ4RrSPYftSM3sxaxvUgCcGfByVEK4eEU
RKJIdE38XjW21PWpbfMXDbmS0B6f18FzjI+6nBJ5pMG3TYrFBMVKB4+gbAQI0BVu
tIQptMNjWBfXG2NrKv93dbE+0My5msrZlq8sWNF5q2JYWwetgHOM3iADebOCzkwj
VLZS9n+FtZ5k+qhL331E4q51G7TkzyHRO8BzHYSBjKDu3D3mk75nLL94zSGiEFPV
XmjE5WF8kAUTVRs3R4pLs7L8nKEy8nAXdpKd/PrVHLA0R0HDvJ2rRjIBZtbl6tiw
D7f/dTuXJK2w7DhvHmv3tXb6W1JcFGEFWvFKx3lqh7EyF2cx2euIvkdsI8nzNyjl
F6dCYeS0QW3xgme0Mdzjk79iIVb5Vej9UKTfd0A02RCalfOVqPR3DsWol1VSCaYR
lvNaGHbi5KcUNLm70gzad32wER44McLTsppaMnSlJa4kU2PJUwmxF8owFYJhm1rP
MLJc8gsxALQ3GoaiFau+ANVuq20C5vgz2TtLuECW7QUdZ+n/2GZwdvmxQg9pPrQx
zg0wdM9Gs9Ctm9fKuXDoGxTRz8V6KAP2KT7iqjoMkZ+i5YZgcPvPmIA6CludFVEE
Q0OLIcv+vXDdqcOVjmjCVtK5lWlMlolIx380F18FQJRdIdkyaxZE2ceiRWtRHP1Q
V/kAZJ7xR3rdhJs3oBEEMqPfKm2As4ATPoHqlD4UFdcDP0qsKze+hxzbsvfK94Tl
AddEgzJS5VRhWkYG7S48+tT7gPKR4Ymb92VP8P/fZeqbVVonyMbQfOzP9H84o61k
StQoxP8afT3ESrZBHZtt6WsByDCokq1LJu0Q8GIu/JZujpibMJ8Vl90SiaigLDhK
e0s3EBckrCk8K/znPAf2BhXX5pCMkaGLfh2YMOr+FbMzV3C3jeil6l5vL/pRKz0o
pSu1HyAWCor2dRjVkU194IP2mbUSZu3DgUdz/j99l5S2koHVdrYlnKCbhsoLXsH2
Q1uR7GmitiWwfenWj4yfemTvxMGZu8e6N25nmbuXfgu3hDtUOSPSSBgsKPAaLSb4
nUeXTV5kxupfY4x35K/fgGJ15ZS7/yMEYF+lhmEC6Gk2BhYv5edgU0COL6YucfOy
qKjXKQif4FF5eoHG74hwlvdbVt1uvTLsSTc61Md4Y4ki10KppXR51PnF3Ov/yWOH
luYyduwVI/MnaEQF2HKDyC53BoRJTqsXJMQyF38d+EedCjjcESrxPQvy4tQLW/ep
WTQX0TNhhmYreCiq+tH3D+U1Gmc+M0p7bqd05kekdADfy+qpjnLXaqse5/0O+GjO
vzgDIHhPSvQuV5uTlV8WpWY/rlUi9VW3b68Ilg+6SD7DteEXstSUhNk3I1lGQI0L
jx+PevL98vI1r99SDp6Orkdaas9oU/YbbW70uAfdq9YRH5b5vlwUthWhx3Vh0vjm
OFnTVoczlr1tyBMLLf971TAIWykX2/rfNMYl6WI2FOnstEeVeoCA42LERj0SijHO
78o/1rq5qibYV284UK2Q6DXz8FpnhHaDoUasehyiLIKw5RaW0z4+lNahlbccGcae
imvLIk0bLhgEDBnXG5IQGiXI+sEQz1Tijoser/hMyOY5/7xyttSwNPbQ2exO4hTd
CJBCimwA6eYfeXIlI0TGvRcNz7hwJroSAjTa1Pz7p5DJWizVVSfr9fZ8ltA5pME/
ykeB0mvRtPA9oCnGufttxGImYPjHPGwmc5+A7LLK3cOAYAO2YnZHvDmkyaBuSO8q
jJkoZEv4omT1mUplZ8LRXjyZNrRuoEeWmnU3Y6xzbqAGBUYT8Q5Ccm3SsLX71zZw
mfG0PFdL3Q5DdJfIGpgasw7VWj5hmafTAvlnX2CHIwf2DoZEIzNonqNLKIXJrt1+
DLiwS8nStTANipL/PNQ5ihh4gUG06KgL+X7xaES5rh6FouQ5BdBWmGWdMBsrDpaL
a/3uHwRW0+sGsyUyE/PwOsI8fkZecOeI5RsT3XEd9UBnURGZO0gqbh3ZnsoZ5wU+
dIOvMrkw7nxfd1RUfNLsJHXe0RyvWKMVYV5zgvWclRZb6/2L/7zERIIn7s14I622
FTQcmIwvaJgLQoU4kSfd2iTrWGmEo3ePsT8+dOH16uNLBGA3YU4Rzq10hMAdAHus
Q8uE53ONUkuA2NHEb9+JAoxepNCMSA14xZCgGXLKdoTRvtG36kTcMNZOLhyRXBrW
kKDlHMFXN8XeMK0hqR33LsFkygaBJ9rfuWRhAZ1Sb/AI7mgRi2SJJhKBT4aNAnzf
tXyfGQGMB75R6X7/0HStgtdHQlpGWkaeS+El0wSjeEGZnFT50EQ1LvGBL1pmtiJR
S3961GqziVQ8hWEqQ1habwjH+VUd0O3Obe3dXVZziwoUi6oKpNH0EuSRDbX9AzzM
jbIBFqNkIVl6ffV1p8irj40n1+Deu+V1S+pTF6n6vk5m8kjJ32X0V02MG/g9vSgp
nj+2X+EyoJnVaQd/U5XsyhvCX+QVWrQ0UWKTmQtyEmZt/XwSVb4brLk6j5IvblYe
Qa1EYTcwIdAMwn8u4pTLhxLHK3fyctELYcKisErdRTGltZIFN81n9wzcVvYDqFBH
5ZEZH76Ye/Pofqtb6580VsaQFUJtNadYQ8A/tWZG07ee8tKWgcMHlnr7lPyHJzb4
phIpOhhGcyXTm6Yke+1501QqQyIcd4AdYIzg93CKMyus0atZN72n+Qjakd4m84DZ
KYoYeTBnLVEeywH7t54GCwb5DXzz6A+bXDHywc1NezrN+r9322mX93gawU9utxqM
t/BQr7nkNSQ/Ipqf3I433bAbOAj2vvoq2F7IgOBhLykogZ1X9/UZT79GCexV7FW7
7DRzzD4G8mdT6YjCxINehpBHoZ2T7Zy4nMewv9GfcBoXu6gC0hCm+8bWlK+57uiJ
yDyjZRfTnMK/kjFrfbMlJ+je0JCK84lYCwPmPVu2WRZmzOs1lOzXhI47k/koxvVu
hgtTKVLSHruJcS1EQ5BIAuziEyCNMS9B0Hsf0KY8KGyityNBJoEgJhYBPQxhLu4c
JH2g89IwW5UXe6ivqz1dR6/Oovunlz615Fl7rMH39nm1j0HmO0QyoVgOMMSnBLtD
8s5kDiVnUBTwFB4PzwfGXGA2/jM0YrBhu4ZkX195NDl2JabEwuednH2Mzs7GreIa
JEC/Cw/FTpO8dMbY1gC4Xv6zs/2ayhM492QuOYs5/sYn2LdTXMPYQx++afDjJ/U2
uexTGrrQiH5ZMcGPskj+hFy3BzC9Kp28Kv7Y4eUSfGZknm4N9gfUKaMRfsQ5YCWp
GkYQezA8FY1UzdWQYAyZHfmaBk4IqXib/sITYQEjFa2dCS9+hLN1VuS8UErjjWR8
wA6l1RL3n2urPplFPf95f8eBJQvJP2n0BT4rZH3WsNmOJbfvM5cP135i25GsKmdN
z42XivJmF8mmKdVPKFUDoY9xOmfwEIovVZriFBmTIMqTiXcOlheUli+G13munIpx
j4GAF5JbaeqcBaguhvlQhnr/Lo9DQuHcfs/uKjzeOs1F747K1WTvW7ZlNm7FYFKx
Kh6rtOISYBhhcDCavYqVkuUI2G3WNwsDtIppD7pSqY/H/R3arXGhR1tvCqdWtuGh
0ExVSH6/TaMV9V3sjyf6Meg7Vhr0BaBcgF24gE9dwcZQFSXlGYj8rZP/EKi8eYaq
AeizUf3sxWEz3r08BEqVfu32af4Cqx4Pz4WqHCzoO7RIqsCuKUnyNPqFS5X2eDIX
RAmW6OQZPpv5h9LIEFs5uZS1xM8zAciUHIvaETxpbVMvhp8qefsd1M3MRYsOZfkk
p3179WYNKQ1rs1GeHM+usLxCODeuWNNdaa6S70PI5VliPjW3MgVALQ9qEwgSR0kJ
CuXnLeTv88FqwxtELxnIh1xx5euxtU5CB94Zk4NYYWW6yoOMgFZLWfY7kaFs5aSL
I2N2d/hgh41afUoCgIiL5sj3SRuhUvRvjzeeVqGJpvKc1BjfYGqGXtDIU2dIQ249
qZT4D2SgI/73YgNZ95zbfHRpP58FoCzuDDrbUIICYcgw5O+U9fay+pyIcWwWdPxV
rUgNuNPkUr5CO0TEbcj2NfSCHFAaCyX1pdYETqueZxiurr0fjibrPE6XMnzUeWfC
w2fZBXHGDbFyY/v8C/9j38whApmDz79QiQIqmplMbB7hdTQxULLo4BEa5nep2aPx
MU9OiCIGgiDe0RKLlcRdaH/Vb5yIHCH5lEKnB6zeiTeKMNAFBzcP73xtfTM6nwl0
cokr2rsukJ4AQY+o3TmwRcne194WSsPle6nXtfqHd2e1SCpaoLclGvxlwXCBqWM6
5L+oLbguUbGJQcUEjI8Q3qgSBQM44ne0h+ghDzpcB29h37wkX1nkT5mLnp3ZhMbA
swQY1M5a+mBX2IIwaenEzUls08HK6U7zBFRTbm6bfnV6oC0MOi3SwiHHX3BgjZAw
1+lasBz3ypif9t/51m7hDBj0GoYP2ldUhIm9rctpkxFBj8+E0DD+sRuSFtAyTMvS
1A3FZXIGMBc5kwwGwU9o2+xxATz49S/M5t2OM3vkIB4E6WbFmM/fITk2qTVpUy9N
1CvmkU08w0sbLCX1fZ7wWWaQFneaSKycjNm3WqZstPbNxbPKXmYw0No9C2dmWTV6
zs1Mh8H474cKUJ2jbO7naAFLrFdpSxk/hQTj3GPC2vYX5YzHNYbvR/6FjGHzXLn4
cjnUl2PPQMaRkwvBATJsJADoCu7C0SkqjdsPz9ubZXkuGVLiuubSNBjLvi45KzyT
YkWDCNnQzo3uzaS/YgvD6hm3EJILAm5F0BgKCkO9P+VUzOeO6M4pVwJplCl/V+nY
RObcqrYFLGcwdFn7PRj4OQS++3XQoNE86XUhSfhaEZar9Ru7mqM/fFS1YvAXlNPN
9cXvMv8RCWin1aBw76OxpVFqd6HD75j+d639tUEU908efMWA9txnhOd9js5+oyx2
3gjy+dLoSVC8w4yTWy2gSDUNTwocN5I3MDt6V2Qgd7Jdwi8NdhcD236SwYVTHUv9
wfGkmOI5G93VeD2dprJfsbiHghm/ZczYuoEbsF6uJAlw3t8aWBiCAqVDfDXQ9U3P
cd0iHgXEJxoWFywLRBFDumLGPWEvi7+ErC2d55/x15zVXKnLA9r5Nr0WCNElMb9H
DSFfQ+3a4w1KG/FR8dqTjksrYnlfZmnoSu7TPjyqOIbKa6E886x1/vFiod0cV3Rw
Jey77aXYSeiMsaqtQVjQ9pnvZQ3xq2oHAzt4zRUtPI2W3wuf4sqwlEMWknZmWFFf
s8ZmW3/Rv9JZ+DBWoo7DhCUsqHVt95QJmH3GTk726dZDjADpQf8IUUvwoQQCq4WQ
X3dSBp3slVy3hLC7bdEWECed/fYVWakyxJDTrX1e7jLvhjFdBpFpcH7aaJDj+8Rf
o5/dJ6c9YO1G37vjiIgX3ES7MqT1to1oC0rRldemeMzt83pubmwf/BosyYyCxTr9
Zr2tj7HS22/SiMhDLYk33VxA3MbcRbWDuuNpuNNLmT0CQv0JaQhiyVCnwsJe2OfD
i1xh2SmpCFHEQh0h/mqvuBmxWK1p3ecY6soq6gXqDuGOl5STgahwF+d0Z5e9WiQA
unhc1/l+Vcci+64YYGuI9L6pf1fs00vKEopiTqyjEpjot2Ox2x1ALD9aIcdOyxtR
CvAafFCJM0jmFCm5FNt9kkXU1G1UEhVMPFyZzu6mQ1v7WS9hlFq7hhhA5+ctoJ/8
oKSgKf0XoKgjXwv+p8zwfWXm7VO1+IagcLXIJ4LnvNSR9n4p378tHctuwj3HDa01
JVme2lm7LD+EetN5IGBKmnHIbN2U8txlEyA8YLN1qU2hrDeLzb2Y5Jg1NZxBtBTf
I6xPiNYCSFoEa65QNeL1iaoMdwQvzGh6h+O816j5qDxFVqhL6jgJoFO1pMmHwgC9
vckQ1a9tzytAa62Jw8xhFn+TnhT5MkWWLPMwBeaRuTzgy5demtsOnw3VcgPrObu7
O4UrQyQ3is7eZXVstTeSiyyf3urQ0OpFWqL/75mzi+9AtjlFnh5BQC46+pxPlaW1
hKIGKRBnFFOXshDsVM030G4eKLOFYeR4lXa+dXU26MqhH1L/i0BirPKqdnNHZVgV
Iesj4jSgHcVZ1Ws+9G7ARbUCCCSAt4c5baT/SqgaiFRqzqyucO7W3t3u0+sTtXeJ
oxduBtBMJB3QCetv5Q31RMwmdQC60gs+iUdALsL6uTT/+F+Idqg6BQ4E6WWQ7KgQ
YLfh95wi1wg0oL+GIyTVGhL1aFMNeM+bo1nWXlti+2hhjWDY2mx4x5prg2ez7WIc
5LPguy1biGrW29T9Vo25dvJSRCE2ATcD+uXq4h/SKdSSbaHjUywDa6S/W86T5oGo
LjpakDFlEHmh36bZ0AMU0l57kHziRfUFfSH3Tn5rYAA2lfki3ZaCQs1qAtHN9KbQ
2V1Crb79h+dnX4v9++F1edNIwpCKRHMIKJctul94k9so5qIoCujvAPaNtUmGSaWr
rkhq5A9P19HYxeXXdpl+O1T6fjwLTb4jN+Uv5ekfUwihnx6pZ+wcpehHLwChOyMj
zqlQawQxOz8y4GSCw7hO97U/N9IxHHTdJeoEvGpqO9qX/w4bgsDI+NW3//xksbDA
JYYd4wpzXQ+SvT+U6zTvYgVG4qrwAwcl8xht2jXNoobZOMr+5TBOWmctfKpl4/Rh
CuRQUUKMBFQy1bipn9Ipyoh8y63mUiqng44CMTBh0DwrqkS8raCF+z2XNI5mNB58
IeAj3OCmZi1q05GcgEApqxK2CCKqZz05VrukuJ/hY7r0F/eGYi+sSaCBr9qJfFGe
2+Hlc/B3/CtgENiMPXM4OxtP+2w21edeJiE2NhZblwQEGEJI+M7hmRucRKV65KKW
0+Sn5iNg+Vww3TmorL3GyV7RtJOWV6xHdiU8vQ4CEKgJfq38dF2qA5qgF+uqIBRU
c5xBjwr9N4ZJP3ult657FlL+MpCCICgEhS+txUGFOmTMDKPowyNZ7nyJB8f6Dvum
p65goAZJEvsp5w3DrmybZGgKtVh8ajjj33nSNkzhArzTY3LkFOZ+elZX3LlhkauF
mrEz6K7j5qihvBc2Tv0JD9P7cVZ+gpspUbeiz/1g0A3JwjIX/KW3CBqGXz7EO8KF
I2sH7p3SBGeztPWvnD2XzCkv0IVzTpFGG6B+iDWfHiT3zEblFd9+XN40ga0HEcE7
aNoA5M3eSAz3sNa2FtSk3EyYNQstQUOTx+TKM7CQC95Goie13W/Kvwonagv47FHb
rKLS9/W1PAzuih8pj4f5hMWqQDhE5OEUfjQVsM5nj7c1EW3rFTBBtT2xHk626XzT
lAvT4E+QAkX2Uum6oNxtMP3GDmmj0YdvsK8NNk0gaBHIvLp/xDecjW12+nVe4jj6
ANlExlRqrIS51dD8mB6Jh4SzO6aZ0nqRDnnKzHII29nu0fAkPvONxwID45eJlWhQ
KR1NVbMLPXmQS1DuUYJ4YGORB+bHvkrI1PHVPNLU/NOC2+qkI8sn8HBFGxMLhTRf
dbNhkhujBFqWZY4R5qG3eOMe13+Zub+3lygAtzlscwoNhO+UFuLDHIyswz0G4Uyr
qyV4/4FtsFsFaiDZbUh2FXrJHXUZfTRccJQChqEkRp9MgRB031dcfVJUU466xc3C
2ZrsHtgYb9beKMVKdiFr1x0GY1AavuvLTVwK7860Sd1CFbjhn6yxpuFWI48mRFjU
bmiaae25KTILi+7H8XwhbXT3wXMN5SHL46b/fr3lWw/ukFEqcW8M1qD+WEFmvz8K
1heTytx0XgD491V8XPhyFqoztzqKAzSO+v8ND/OSUR+U4ErlOm+XRUt3YnFd2T7X
0l+3o4d9HP7BrNOMGpoH4jPLugIlgHL7XasWM6nPMDayARr5X82r7Rub5PqrNtmP
9L5EcY8JRu4bPPY+H067bLVOq1kwyFsgqxA78GWuqqMIbgEwtzfGJAjy0qaWxAvV
R2Ae0n6GmZohUdMStxRmxOalg7BaMAIy+b9B8R2y9/nA2zq/L1rHlmC0VfH5K72U
huoZ9fpF09gN6wb/HazLdTs5jUAulOa5bsXjNa8TqD7fA0uhqCkVZzzW7SKHBjM3
/x5PYyV7d0Z/Wr0kkZ9biGa499hKyM+rJZ1XCMoSq6Cvtz1QBXrln/KTx1l67ZFx
VIHe0j7DPGixFZ9E07Naxp5LycNn13kbERpndzVg5hzYDuAHaHZz7ITQhLI/ob/Z
EZTmWI5+eEqDRU30he+L1ZhewktqNc2r3er7eGacHNR0cMs5QHUeMPuW+zWcgQBa
CMyCw2kYQ5GLD3j49FOEjEhAFyA+yesJ5G5omleVNG72FPDWvTL/sZRq+RdToSNg
7xzktH2vx3sD5IE6VAts03zWMAXZieq5/TiFMVgazeG27Z6m9HSjFWILdE33bx1u
4zbrjCub/vC28i9Voc8Ckj/oTiDLv6K00djZvFGkkMfOVryKF3qATsKGogzeH78H
ETH229lcdRWIXEMreblDNPmowoaHAos+SBwbV/uw18PK5WjM0yyElShNkll0Mhs5
fjvykyaCO8v4Dl6eDw+uPPcnw6PtvR70d6srqEI4+P+VyY5dQ5RK94ukPbCSl60G
3E5Fc5CmWTZxpC76+/DH6my1Yn6nxKNOu/wfw/OMvofv9D53wbXCrixsnROjJuyy
JqaB0jW6m+cZ7ctMqy773ZFYRPskmNpjJz7nTrCEe9KeBUfv2sRGlVJ2+Xp3S9+o
LYD/vaWDQRz39dsvBXaOX8txfyWtknNcui4GXSKYXquFpYt/Fd0q+kV/is/4jIKl
uFTyWGIsq3XKF8JWkP6HYnXpHrU9kPVWviH/chJiKKoc4QAWAiL4fwgGmKCnH2mM
GMaDDfCqPU/+rH3KH1iHevfxbU+IIHnNLJhQjMayCr2oUCn2pVCevDjK2P7PHQJd
nxYxW4wRKsz+s14DQgc6GXPKm2KUDJx5XvVD5/M4SllzTWoyBdyM/G0HLP+4sukX
JT4jwu1HSFxytV9+RhQXSRQ3r2JG+bjEW2zUJRhFz81yc8PVz6ARaXQAx4PIbJX3
MaN/Bdq2K0Ea3ucSCuK9HMSMswSvV54h1HXL4L0FDOSs/kByrN6kFDkRTMtRDJ5x
O1KzwPI9eKmN4f950lkGbbM+jh6q9JKMWM2ZpfeUayLKbRa8q0jqcELqI5AIGkzX
/yHkqSflibdBZTupD//GLcg2bSyFHUwrQs5aakpuvq41cQog6ZZ03aIq7tdG8rVC
q1M5TMy2Evi5+578S61R7E4aAPA+D1+5PMfa3Wg4YbC5fD3yqfaSz6wWWOmjIz8J
jK2p5xtoBAStanuCS1U4UDS3j2iz6K83Awef1Vwhxf7dVjDmVU2H+5dRcwQuX0vd
KX20KsCt9jQcf3XNy4d3ATvUYqmlkSCkKunP6Zvh3K6db+CU8VYly1U8mhtBRRMY
JQYbgEO5mCjncnz5sCL8YBIG/n5pCcqe9u9mwuMVZ5eLfknQjBjYtveiCehXROiT
2HZnVzXvIR7hgD5HsHdj9QSLa++nobW3Zj4sCQwYtQG5QIjPf2hR0GkXLPqAR/xW
Q1aFJgbqZJwvjRIvWFsMaeHKlQXze/1yyN4wFsgb2H2unvtjb2w89y62bITSDtpn
h6e1XTErk4ZyN5vaqxbgmh0M3PneOozR4KAIsVDBEfqepPbh29V3L2/ymx+Kgb//
Zyp+80rEbtO2dQ+ByzDdd1/smFRRMYbRtEm9qz73DvK+BtYRI3eVjgacyoeDhc8N
nHb2HOSKGbITsWonIJGo8v7OMRTEazRinohvzlbjTNhwYmIVQ/jYgk6Oe2RI9yp1
WHwEGcM0OpKNh5UpxmzE92bVG9PvhMIQdNW11fSRnKqyhQcX2c6SSnIW6cac/7gr
IOfBrMDYhD3QYS1aq32ARofH0a//+FsjVCtMUSkKcp2vO2WMXL0R9GsEsELw7t9v
puE0TNzzKTbv/6bjTy3hk4eCAm14DG3bsXlyGIA5mBTzWDh1JAsdJYyu2NeadXF/
/AxvqiWXEAItWT/CJGwzfH//bgXute3swV7Vxb+V155s4/eepbfMdap7g0oZMqDN
wbQMhFtL6x9HaQ6DJy8ss/YICWgFgZskRx1qpkOdVYbE+dDLT+i3M9XhSh8B9M6c
S3nSPasybmZbrfVlzY3FTMxRsb2YVD83bcP5ff5LNzi1gJHThyDfTaewrV7hFKyj
snUxamDcYXv/qFjtvzMzHSCQLZHxGzN7xwstwaprzGDlZGUZMh/CDBKpDLq95C1e
/dSjE5yZ1bLl/NJ3UHKlqHfqr2kz0htQAkEvJ7VxZQe/Yf3cZQ3rhGVAvdWx9GS8
/eNKGu6LP2JrB1TuoC0C5s3KaCm7GI/jg9xHf0KdQD/7SsWEV6/zw65fmquDna7i
5b+uRUG3nbFhdTmQ11bYgVswiGUJMCF/dXpyuksbx+YAueNl0kFe0Ka8qzIUV7PP
1MEKNV5G6X0yjRgfDYi5d0ncPfLRUf6MwAGIJ/vFDozA59fxuqL4+t9M7vtfu3lJ
lnG3kyeEXb0AjqkN5crx0hZBlMt8tHGORmP1ciO0XzOQrrQnJu/jW6Hklbzr7wAg
c3rSy840eAg5OE80fJvF1MdDEQw7Oh8HMgYw3DFhzHAPt1oMaIqdLjQZdyA1L2An
+v0IVobgByN5usMkiauVXYYP1y3LgpB/9PFluBG+5XdnuWFr6iWg/6p4Ie6CSrX0
codxBZuaB1vNcdKSwyreSv6cIbzCitWi//YpK0xjZOY+GW/djxJcYgurFYMjNyJS
Cl0JP4qSuA+wFksWRFWnm4RxWHIG99KZVyzJs/Dp/lZQ9sB4x9wGPl4qWGj9JfeZ
aJ1NV5QjgZzXAGkoEjjs471/hIeZwRCLdeEF5pmNqJGEfwi5a2PUkHjB42UPFlOp
GQrZstUVS+c4drzHGcrHcx966XIIyO7Ct9qBrbjcTx7alSYCz7/CsOB+c9aRTHPc
l41FJ3j9XMBc2UNK8I+35b41347I92+GH5/07YEmeHH2tNmUvqmoMqGmpLU1WvTV
rwwFiKrCh8cz18ZRqGMrzIAElCAbaygK6BNOLTNJ0z7sOCfpDDN7y87hpTKk/YSH
1oGHR2zei8CbPXGnu2H4D8S5va6SMZhe1Dla+8grr2JZG6c9tvjEFAw418yI6f8y
uTpEkcUFY45YDboyYCHn7f+ZlplYsvaIZJABt6weDlIHrvqdJruPx87ihhkOEkfg
ROp9Rv1ZwDr5sqDxST5pUkCd3qA1mVjwtx0c3N9Q5vZo2STnBNYfCT2DHSf0Hcw5
DmrPUWcA181up7o7drx/ZfcKxt4ucOXHvYX28nRykdX+jBaJKdXFQZxw6GpKQWDP
DCSh+fOYpd/LgPdQKQhbkt7TCxV37RpuI6YK++99FmqpsBdcxRCqscU7+Xf5Iyr1
LRC83mDkjs9+pav/RStXsJy7FTasnu2YoVatjxEpL6XT5aETYCUFQCGvDmj6MOgv
SP2JHWsjf7rpYfZcl8FGDzf5yDrqcUYjOA1MwtRt1GJIOLw07Q5HxF6jSj27H5sZ
w7v7dJuAPQ91oL7IxtDX6tOL4ScmbddMz6uoxpuPo34YjNBjMRuUEGYXVonphxxa
6U6Q3hXEWlAfAMYDZuttmV+OdPi+jBm+8cFfuC7gUbfDO+RFv32NsQAFgVTxUw2n
cPCLWzUn1LOjx5ioLAvLqGcY8+lVA9TaR7OLBinmap8mqVj0rZaTgJQ2RdwM3Nal
cGeNnKUGz/xrNYaxCUAns7gjE2bE8EG7vEkR4w2DPVbqrkNIn+PW+IxzZo0xzdkp
NEzZ84WsuTHbi9Z0B3m85C2DUz+FRvwu2z+lwFLAG0zn8R3nsHsCRdGFIQ61JehZ
D9Jpq8TewTU9e7I6l5Q017tkRkplJss57JU1t3aw0mLPxHnQhL8Kt2xxhtjZKAeC
wp6tqbiKvwZswAtTG4cKSyuho5+5j+ffq+gyyzgxk6fHT/Yk0rJ/kTuj4xOdB/zY
QYQi6dV4OEoFwEl+CtL3zRIFLYDwW0J+dWH6yvzh1OXoIyJtManXZgrWlvmcpSS/
ELA62aK0sRT6GWbJL2wD3rwM8d/6uN3X8cOWSwApb8BkSoJcJ9Rdz785O//VyjRA
RhOoGyO/YoJo5POXI9OFW0E/ZIGQ50OBvNbMGFn99lJMlqAJBEeTdzQeuNgyrAyL
3hq+hmpJBPEnYTZ259i1GqwFT9qwbM+6SESNSkCIW37qwb7sA5fTGh5wryFkyKbi
9SCRr2nuuqk7/1eMNHDYOYYXbjEhsS28rxs3TMwVk3Yn5eY64r3uI+F0uRDQ6baf
rR5nNzrBH/Gk3EK9NSZWgzEKzn02giUeCvNKttLcIMd7NCRdM3/QW1DvZbLtnUgx
zevr9OV71oZpQgNZoASRQ5l6nDOweO98QwA1tQCgLVHVU61MTbmUShqRZ2BtIwPN
yJPtt/8Ce872FJdVlK0UQNPDAgfRKKR7J2NGKVU66e/3x4drPZSUp1LK2+SspwEP
mXn3QWmn/b4ozcCnGC4VztIFlwRF0jVJrdShwThiZ99fMcA8wfBb6ZGmps82s0yQ
44JisUKNZgtyGa/jhg9QTDUP9y8RZpipp9WEaAzQd3+oB6DL9vb7/4syJVUY29ui
7yU58ZWy9X1jMpnLOsD+qbY5R8ojGNL75zQVmzPIUx7x46W3touwMytwqb679xD0
VUrm1XEEOwDXudvKCD+IVa2t/k6jUawJ6dvOsS6sJQID8QCtjh5pCuRbu3iPE6Oi
sy9d0sR6YJlpP2FS7WHpgVZEO6M9yezfH8nn0HFj3vH/N6wwjA1T5d4mDSZKh4qG
ELJgKQcIbTon357F0eitQaejRzmNwsFrYARGD+ObtbNYheTEcsMI+33t1yHL7lLw
/LV4vFhPKxWZPnsxxbRShP7+rZIFoHfGzi9RewIuLc9i4rN4nhUk25BZavqJLkZx
ipRW/yaCc1husRI2jgC4/Cu67P/B85ygRMTV72nkSVFDVpVT/FlRA9jleBa5H+fg
3CXqHO8J+kd03/9Uvvb7NZoETi3eeaHLLH89vpMJQT+A6HZSrvBsASujKY2EFHIm
pgacDG64Fo3Ad9Mnxs+HgrrYnyf9IoHHTQTGvEw/oTXuQJKrTjnZD4izO5ZpF3QE
yQrCRcP2IUSHuP6oaUpnnAKXmpHsQddORd7cVjv2izZwjkzEwMcQnTdOipR9rinL
SQ5WVLsXrX5qDrDtVWViq+FPjlo9co5fAKScXixoUKbmCN1VXM88Qj0tNS3LAYcG
7WWe5k0Yni+siDCtZ05RdAuL0ApXVWm407U8qhJqlNCIxdOn93YCKFWqbZav7Ciq
plJTERVvwMAYlnHc2VUjGPkfWx+T02aEvkmq5eczlc0VGHv1bMhDkS0LvbLIyQn1
+6K6jL8Niw5H4l/yCSmXMs6ujagyFs/I9iBEYT1QH4p/v98kd90YSxEWjRUr8sSV
Lnm1xSg46mZM7/7JSLUoH+hNjbMhcn9vk8i33s44PRBnFxBoy+JmJy5ov87XNWid
glcgWeBJQwXFDRHco/tfCn8Cy6VYRRBNZ2vKMQ0yXrCJ9lWfeBs5buEtUt1XywJ6
ycX1b9R951KQbaB4zgBHKH6k0ZE2KtjPvwnI40usz434U0D0vKDehKL27ZDvBKRx
OfRWWw6J3ZGzeCLYa1mGkUikVQZ8kb89V7bqRUTT/8031hOKT50l1vCAMep6RJJe
ocb46byuHnkPxNAHnamHJM7/Fh21pCn2Ar4Sf3FxCVEuV7yVSrvP1g2FAqbeX15t
jJIsOQyT1SrXvCt5NfEsQjTU2EPcfnEQqHXOdT6s1kEmveZrD7Mj30nnWQsIteOd
JpAyKCp2rePLHEQce17N50I9Do5CgdG27U/v0SFYaupPTetqZb2GuzEx/O5UPG0Z
m1LJRi9ItfzY5SwJfR5SMa1zvR72zjygDja1MuPFn1+yrqs8KeUWO0gKo4maFpOd
AOBr3iGKdo32gMV1wTQMvyA9BOFPVElLm626yWmfi0iAoTMGkWyTlGrgj8m9uKgQ
/AFF6tNSzmdShybUnG9MQV7emV/KmlFOXt9lEMGNlx8f79A91jHzPUamLcQrAapG
hr+uQ/K0PSrnfVrFVqgsk9Q6hA79tZpDy7wrandwbSpqXil1ESsAOc732HO43imp
+s5FImjGNLWR1xQCeZptar9QuC1uF5OQjVjUF4ZL5D2chR+C+E7DzdxcYkUowZjI
Z+VEBgK5GDVkOPpVNKvd4jgGSF7AIz1iIERVW9/R2wEghdFW08jKaDiVfItRMz+L
0zRvmRDNsxw7ZDwgwC/hethQSovCUzly+0UG41iy1/lHz26Z/S2ZvEU1ZFAo5ybX
OvyrfE9WYbrPm7iRGWpNb7g+ISz2BDlVSo0VNyFh+1P3mAoHTs9v9cMYFDM7EEQC
kr+swFhW+nHzGgLtLECbbAK4Sp1V1ncP/B+CabSMalDkHTm+5ZAa+Vpf2vZvsZ25
cu8UkKX129zrxSN0Gh0Ym0tNE62qBThbcMAZitv9DfQNnUwTQlX4YfXz7dag74Tw
ppsstj6ARgghhVmQEIWnM303AcbLMva+cN2HFXWATMFKgfpH/lC3kBleiTMqLkRv
oPM2wUq1bEO87bUmnl2QP6oVfagCkg4A0F11Rf40aMEtyoyfBM70U6fMgYZkBNJw
4Il/Yn/7myzMRBFedQa1F0IYsq2xfdvTeu336qnAArvzcpdVIQC8kvSQo1aKeDdY
josOZX6Pj4/ej4VqeNqCZvvg1h2qJ62Sy2niiHVM2OeNH7o7DhbB3OPquSoIXFvi
ApLT4amQd0GkWdf3FUNRNbwrui3SR5QSE1IEql7YfCB5dk1HLen90Y0yccyonpqO
g0wS1P/bFsNdg6KzpAkUL7Z6oYWe1YQ9tbNHw6Q2hwAqQZ9ihA56FtHazbMNLNLU
92vOCIIT0VDmMbWMlNzKJfjBwwappF0zMVSFkdx6fn6W/8an+bnhwnY4OVvUFQ0k
/infXvFU+J2S7Vdxjm/O/yqpc6xuIJl7STwGkm2Kr9hC8FCtQAM2SIlHPVUuxOVH
kcCfXlya46O6ZeLJXpb4NfukCinp3ae13enSKZxneoyf9meewn9PmM8teeDqorE0
kRBRBvFa+0F1KgcExm9kLCw4X5LKqpEp/NawP4vBQDvLcg0smV2A1+QZUny/QK+s
f6LCtqUdlBu4T/egcpHf2zmRpH+wbuJEbV4+B77rF0t/7tZaltogztxIE1nFsbzz
ScCQri5/VRaam76jAbJAYcVP0qosMv5aXtVSVcYTNuHVW/XgYS6Au3n6eD2pqW+S
Lu/vncSisXHA9HnKSe4ZYYKp9cHZzw99yLIkXGZdPWQSh4oT21mLgDFhH2/q85bf
HPT5y8Tj3S+E2RoavsOO/HgFMHgsbN/KSMQg62HMLjp345A0Nmmmnd6BtT9AwPhu
igdZfKxUi5WGtF2jGVxtmla4d6srqy5Hdw38DOHJkg9+IQB7v6Xw8ugtHJ7Pu4PD
C6zgiKeQ+YnleXbkobKLEnl2UV98fZueUCEhGDvOw6JVAyrRN5DRuUkPsLbsKm+U
y1/Z7SY6FotleK1jRCjpQWEZ3Q4eHBqsz9OMpnoaWDPYvNasaJSTMNonUrLp618g
821yJSzba3lzNpE+a8qXHF5ygIiwqoC+biP6D79maF+F9XsMQgRUt2M9KTTDCtcy
nZFsMrYF2PyCmAdCV62VBWb2K7z4do1nJPqAdHCacFe6NLonaeF6jKFgWrGjOlou
jgE/jXzkMk86jWoihiH44orHN1Qin40K+Cu6a+rAkNjzeKADPymuJJ4zqywZjAKh
lxJxwCy6UaRJwSEQy/JtQGoOtcHM6EDLgGyzFgVJN7f4kpIH5WQnjaBs6mp0lu+L
U4xKq+I0+KXtwa3+1pnAf3uqk9bCrnsQmYl2fk47tTMnu5E+6ugBBol+KHrFM2av
GMiadhkwO4bi077kM5kuIdXO32aPiKUUFDVuQvLAZowkxENfTK2EsNJOluvU5T2Z
/Sc+7GCjoLxLZWShUmXKi9HOfEjQ7GP9u21gEsWZnribdBep+23egWrUQMO2D4D7
xymnh3DoODYFSTjXp/MypzHKl4hueCxkuUefIDfFCJiYgAfjjutS0MNkL62KcpYa
bVnm8dy4Y+YFUA8K0SOu4cGqC5pHfuZjjYv9J9HLQjrARnJQJ/yxoHZu8DWOgkIk
pAPe0GuPsZnE8HTl3EFBiZTSe/0Dmd/PVUzRVy1/M7zKgrNdfH0toY/KTRJLB9wG
ncjHVKmoEH/Rh1ewTUa+gycqavyXnoFL/UmYvsRQUd6uLHlb2GYyIsuCNABoJC/u
y12PjLggre0mrWvUGXFK5Vph4mXytJJG44ESRRkq+QyW153IMbf37SEFf0TLiZag
22MU8J2NV9k6OqK6F1gcK1LZnwMWYcpYSCs3ZzoeHi2QoxPt8idgAPv8NsxIc49L
KP2gnni3RRFmJVWdVMKwEt7S9ivNYEFrrvk8835fv6saflENzqixEgNKbw/xcCmF
LrPVWdG7k/faeDLe4CkgSw==
`protect END_PROTECTED
