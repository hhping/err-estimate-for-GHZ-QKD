`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NB4sLHILi6EvQr8xZyoTHWz8FdMrpYFdrlecJdQ/2TELVAUf/WmeZ/Uh/gS0ZuxT
TEUQ1EOiOH/cwYrhmRRcHOlL49W8F6jX02BHUJzmhtoL5GvB30Bc3vBndUz8nbQx
IAGQtSn14VzeWjvhAnDQcO5dad5WDTrZDvo3axv/smlGKOH19NzhS1JxtZkH+nBS
`protect END_PROTECTED
