`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L40VLLEzr+s/2yQCSZn/1JdZPKgGufJ5WbSzMFGn2UMO0lsOx6JRvhAHTEPwMjqH
porxgH8rWklh84KtgqM8JOukjGX/E7wfl46gu7zZaS6VPHmyUwey9MF/+ygO7Z68
3ZDGDFYkmfmwSN4lC1UA+RvNnXel7vNU+g0AEgzzgncZ0nIaWgCD/mweAxy9irZw
iszJ4K39cmsyQJh74v2b+oHLIoZL1gm2JS3pG9cISletqEn88w2owaqtInTAzmVx
mO0Q2Lsq0qOlJr4izmau2VhhDZ1umbCeuQfp/eI4Zu/Z2Qp6NTl5X+mOBq9hiaJ1
/WTRO5IvJSActnxf4f2suJCfoP0BLWq4/8JRYqTog4xPDuwZfvd1Zt/sTTndydde
oVBTYAkrYUHgawPr6YUFB35R2+k7EVtycfVF0l8mf41AnVapNQ+cNa/OrRghG4q9
2wzXJ+QX1r+lGPp/KYvoYw5Bt7Y0yI2pYWk2B5bLqrRt75O0NO2UrOs42UK9Z4kG
qQWi1nA5jZPW1oDII8sct81BxbitxWzNZM1iCEkbXm5NR4cOG7cbESI4hBpklHzY
`protect END_PROTECTED
