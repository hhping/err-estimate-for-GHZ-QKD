`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGtIEF2bp5DtMI9j6xhDQMWtTCCCek7SN5UqhctXxEZlhMgSvHK4iWBYbvjqbaHt
JWAigjv+TxZ6p39bYFMS5ExG38TnVoSUM/qLsnlmDfex+MHQzlLeMv99wQvPGj+t
QhJcWx8x5qg8tp1mVXcjSCInA7paksFhgfLw05JFlzNT4UjKiVF3msWNCxpXRgDZ
dbM9NPToxzohZ0+hghJ5UqwEt6zk/Ka4/qz5lT/gYiR4ovcjyCezyfZlQg36nJV5
H3ZUdlpVqXkX4Gn0pBQiwR4Y5uFTBkJQdVPtK/FkEVsKFh7hYL+zPTOEM+awtdj2
A/dhn0U4oX52prF4N+S+XB2qIK3IJiWBJz9zdhEsedvGsmLefKw+7H+s+EKmntOZ
/pY4Ufy2rGDVq6kbExL2eri/jflbBp1ls8DHeAStYa5uYiOjfLcQdD5CSw7NxDJL
9LsQoab/jlKuecsH8mSp4yCceCVPlkNLZ1HXhoP9DlV6VCW7TMkixMClEGFSbRNZ
CLFou7pngpL5KT09mmTw40Evb81ZCu5pC5lpbMG+gCCCLWvzFZwqpSs3OWojQJtu
mjIz6LjX/zD+22eteXJm8PN/mn7ozemS+/M0ZLIWQb+X5PgWLrn5tffq1KBB0yir
apr8CB6if/3Rj7Wequx4rgBC6TqzK/OvIt4KOMBTFAH7Z4HUf2NaI+ZanZ8j7djb
BWQCt0PcMAX9KCeHe4UeH01kFIh4bDjZ11364PBfo2O+U7kT9W4PELVRnTWeQlk2
T3tOSgfg1k249gjOjAVrUtPfrRJoOeJ7wB1E0SRzW7k9ZqywbRmA6ieGfG1j/Q/h
y9ULQWAge3JSgVr5fEEl1gCvS6MATM2bQ7Ie5r+BCf+mOtC5aoP1lGLSJPDVaYsu
mtR310JTQObXnziwUEcVoL95OcTt+jobr4HuP8bQsJ2MDamm4M9wiRKSrjqBopc8
zfGVpFBsDaWPr+QDE3gP4ts4hlhWxxcW7NcaUR8+H4MpC2U+7euJh8Iy8/UuQlKU
zddUlKOQ/7031hdPywJB2jY39VcRSaaw3ep84uhslMDeXRWqOFl5dTa73zXzDEMj
LGYOlZnSs35vRBUmr/oS/wpuMY8Ubrb/m9gsLQUbvk7bMVU7j9yfOkGbNHttC+wd
OSqeWK1ujClw2dDJzFh48D9jrim637FE6yCZ7cn3m8pp8J5x8Vgp2XouAXF2nqlf
VFlxENwKovXHVS5kcRZstW/O0QzUU7ZLVe0BH9fc1+db5/HWk40WiVTFLTdeDekr
mmPxVz5OcdnS6kXw1NTi02HDV72i6eWpFgvU7J3jnoMov0NEMnDJDWjt4Sfzzwc/
QcTnLVfKtjwfeantmBEr/zg/tvPTBfbKL/1tIT+ggYnNvd+7yzkw3dT0YWWb1reH
/VWKW6tJdVJHoLx3SWsHdzsf9+bprJSMOHgy6U8pjiWNSweXv/CCErwynxqny4as
`protect END_PROTECTED
