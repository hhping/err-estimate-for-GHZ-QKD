`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JcXnOtBkXjmKgoLj8uTQHgmVHiPH/42usXJU+ZxRZ4Nmc9HeVP173E1vDXQlHcmK
HS8AYA4dcFvA5W6rbSywY/UdrX+EaxGH91bGxtMiWF/tsPbzDyAaIHO1nFw0htaR
hMjG2rt0Qh/B9FF5adofYFTFZiSmCKiEsFQ7u9s5dUt9fnaXos9c5UpywgZlbS9t
O73nQvYzUMNJOpZ5Kh/2RL4IZC1vlmMV1EO2JscDwcAiNOVLsIuxhdjkOcyvYnh8
zaju8L47bDmK+t6Nffu67WNVtXxQq7+fGpdSGKlH/rrH/8ZpRa/eX9uJkLUuiSVT
TBThm/ULKDowZBpEUU4u0Em/0GWFx5vSIHFWkZNCLQJAPVp9mqQXmg/AB7XzT2bS
8dSPQypdBfE0SjMPh7zzWlyULTQI1+Ag5A+mZmlCk7sl2vYZ9gTILtSzvQIqTx2y
C8yMeqgoBEgqHUwHlD2rr70LLwb8V1iqFgt3MTIQFci/hiY4Gu70jRUVxIapdy0w
ARKdU4toKLH+MmV6zAhstbmSZQnvG/8vFHGrLbxnw3fzUaJCcuwJXX0hYJb1KXx1
XltgeNaDmF9i/8/Me3gAfRziwge2p1QLux7SfsNDn7UDNsIeJzmWhXYjD8ZR4UCM
ieVYJIqwOwQWAgOeYyM2Jk3y+uFBjiVUb3xkVjeqMamG89yO8V7Salfv0iZzzyvY
LDZvLvrnkqmkCSiNHB2N5JknKHQgt3hspI+DHBA0oCD+3BbyTFkHeoEqnXdHrolO
`protect END_PROTECTED
