`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5TmfVCdyNMl0rTnowAaw1XDW+qHpEpypLoZDAyhzTtrAFqun20IcRHrQAYFNu9GA
KhYUlbdY+P6+IDAy7CTMT3ITCmi4Xe2mms1JAfS0mNx7pLeffXBH4VlDaj1tyCsg
cltI+K1+iIlV1OmXPs/F4sWpxov1a9v7ei6AgvKTIznUYNNn9mdQtoTH2+s9tRjn
qLToeUcMgiYTn0wI6QQNeYFrfXHfXu/lxEwwdQ4bg9QDZuizD3neM06K4vUHweN8
FWrKyeZACDskebtAbA+1DbYby5TsHlR6r3WX9RV24PWsCnN41YgXrRYc4nVYcPF8
GDTK3uyPhIJ7yik37mLRcvxF+BlEDXVbRdruRdx4m1P6WX/3Ry6Qos304UxNGo45
EhH8MSg8oryvgEa6p0bfN9Fu8xFWO2SNQTLM0mrknvH/3ZmAFpVvShWWiaYaad9/
9NIO5vEPiqeY4TRPkxj6DdMX2boXLkeDsN8QfgHXnongl06h55HiU6OXUX0f4It8
9zlF2+mTr+0pPxqGKJDfpnn85UeyNmRBXEoy7Dhr4SzICtJcT0MY4htysnCTy24n
bBhGvxdDqcC4fAD9H0g3Rxs5f8kH3S08SN0RSDzuvO4jJQkmdXtKGAE57Icp5rK5
lMazjr1abvbgC+nDiSX5uEz3dTOC5SBgJgXkNIQhUQx0wZAPV7h/fRXyz7p8o/G6
/SvRTgQ4z9TKMexOnDLUv2wRNFri+tGuhJaPqEbJcEHMOGIJCS/Gk2DiJNs+muyc
osxPeiQQsK/vcmkd8t+if1oAdbS5euceK94ZtUigwprmp5w27UmqTt4B5oP9nSEm
wOPDXBABnjC/+1958fJ6SRULIdB5VRfraUnAIl5azQl02DVTqucAt4d9LhOotJ3Q
Rbf1JS8a9u2iIuRYnbd1LrKTtUlA16TJXdpiM5h7dTaa1QpTeSSq7UKpjixql7gP
28QdO5VcEyxkkussV9CSdjwAx/L63MeNskukiIlwCWGyjy6nBVsVwJE7LD8uTN9d
8SmIoqmTLWYWu7LOoedaFq7upaEo3HuSmgBbUgfS0B4L8UFkh8g0oXEISwBmsJ9U
yQ61QL3TNjMPZqAP/9KOhDR2A2+Af3I0BZIwGAaBISFEF+o1PlhKSlNNEONvHeE1
MmIE/dUmIieTlCtQWrYgIqb80L7QV1UWc7qwN8ThjR2GmoDEbAHkrzo9gpdNn+rZ
shmtfqSETxSU+2Ejra8RH6axWUexH3aFkGHaiGoAR1GGikttZoS0b6fF4QQwtnf5
gpx6TWYI+J+c7wSSTAr9nAHJTkAT3qjOCBvSync/by7w/QwRZzBaGAG5Ja4Gf7U8
XNCtZNM0ZqoeFOVEOs5nvw==
`protect END_PROTECTED
