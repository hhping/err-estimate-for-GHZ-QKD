`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7kmjGhOQqBnNCUd+5jWzihkIWqPfDHfzriFn4jhgyahz4eGQ03wl7C2qBl/qxoPq
l7RkSr+8uMICf3bd0YqB2O6hw9EKwNIVCkIVGgRpuNY0zMcWV9JIx9hUniNSKHOk
woPqYaomklPm4Rcc3NOPmdirixKenVXEIo2ioJED2+/ehS/n+nm6/cspPQ6N7zce
YpkwdmxXuBwMf5e3siQV2BCYZUIdYVd1iab5LKdzgbTDsU6NazFpbPgiyqQO6mwU
9YR9zoS2uVx9SzoEWMfwI5vtN9KFcB6y9rFj5FickyAc2NvlBQeAb+P9isr3GB1t
geCNQqN9Pv8ryEh/DtSX+9Q1Si4t4QZOKd6T/+Ig+GNUwCoXfC0NC4OYrVcVuPQQ
JiyTbygnihvWXxCm6Lw5Ie0W6Zc6qjkuN/r05gYKGdoDE6Ku3KH+4EHsAG2fkH8M
CKCFf20fxeV0DiKT00Akbe1BhZdmSzJoIxuvUKxqvIyYnYPiWLktgpVo2pIiIKdi
SfcUAvzQikavBy7NbMfIvIREsbmXdbzvvNiZSW321PzKozq6hMS/bWvpv9EcL0it
cu/uTggn2VAJH2EKpQWGaGhr+ZkWpeWYxYWrIDbVwr/HDsBIAW/ZZgygws8+WBEp
Wq9awVplE2iHJEdFr2ugBJNUvkRR6ONIi6fybmL9j/8Qmx99XX+q9zqX0Z1RGgdp
j2h6Wdvy/phK7tA7AXgkP3m9aiswkUxqOwHOPVaOseLFplTbyaWI7Yzd6Kgqh0aH
tpIUz9xKxflkJWfj86jUYl+h4CbC7GDvSs1u2XtPrl/YySSnrAe3Rs7PP12P1sHS
uJq/owIXawkpceco6qR9llVYcYebm7YMK9+8buyrewP61rNTml8B7gFgKCTF+h3Z
BQnTSwWXvTDG8njjb7uXfYywdJnK3/6zvLYUFb/VmciTtyQXT4BaXFWZ+vBF2Njc
MgYx5lAlf5bxj+zSKZQhdLhs4QQDOOWjxjBhSCXPZFDMv8/2HhGWpZ6qbItZQz++
glXDLcWWeIDV8Bmi31jd3w08K30miM3svr+1/lN0+gT/CgwD0LM0yj+hGYfVnJwN
hJ8UKofCXnr7Wgcr2OIgD7m7Zueh2UGqAYqi+MR8uP5DHZ6IaDPtUzBq+fyodDnT
u/UOzgCVTKESTevQORHQtr3P6cFH3Yms6vKkbOrNNIJZrQD5NvM+NiMVQRoV4FNO
L67pU7muPnqDJnOiNJiQWgeZ3ezVCUVptk5hmeytmeMQy6q+1Tk992Ub5dXFEZFB
BvHFNdMZBy2vOJ2wW7XiE+XfOWUF9l/3w2nO/N5pZyM5ESVTiuX6FygUkNyn5Azc
1pDYiuXDVq/QEkiwxbfAOkyAHO00r30nsDUOCWaVbq9HtNKPYqDUFmULt3hitLH/
PLrcQqQjL2YZxxh/Y3Z4mKvrVRvq6GpOAMbe6em+1pavlPZq+nOihuLhlQcuxnhl
9xrcOLB8osFuMQDur/ixLRhKUe6kT5+OiLgL8aMAWgSV1gW3JULPos6q039SZ8R/
dJuxz7RQxgKfII8ukxfYbFVHwerVTtzAyfrlceKJjcq1DNu+y/wYRm9woUGWpvrQ
hRt3Z5FGocYYhTt6ByscC8YaCbG0EGg/DrlaDc5BjhI8VX7L8mxZGfeG9fuv1AKn
s1u4SKbbFMvVglXSxvhcPuWrMfc+YocmNEJsFfBBZNMGBDHNs0EDDCkesSytmW2k
KF8cwQ9GLXuTvI5S+jqifKl2UiBS4CwQ0WUINcCXo4OEK+QlninTL6wbi4RIXIwG
cI2AsWlN3+vpCuY5VTqK3aM3mz5F/jeeJTwQxBPR+Oy2og7aBJkXiQxlf+XpCSv3
6elxqDO4ZHk5EmYbvWUzBUc6LGwkw9b1kc/v5N0Cp/KznlIIn6Ym1reOWJeJANzt
wk+YgNd9q/LqDu/IVoTA5owLiIZHptuXcWwpl8/0YMohbrX7Gv6oXzEje4/dmjdZ
Vi5Ya48TH2uagBBM7lCu/sH66PyNZxX+UluwAhaYbpQQjQIDdnjmW8iFNHoDxGHZ
DaBqYrFGyWSYXGr+majp9C5qDj5p3OWI2eSo7NU7mD+T50odS+baz6bHl8GKqjUg
Vq+IThEP48l55ibg6zbnNbcd0RROxOb6AcDT0R/r6RZq/tfrwimmdHQuFoubmYxI
hPEhVmK2R2TAOiwEAF/fF/bB+Nz0pW8MAwXK7rSLdX7o8n3EQHW682bxDE8U4F0I
V7cg0Hym+oUHokWqjA8mURlcOrqGMQBNCUMsg11ItmqzuKEShBUVjx4UrpD/xEOp
+woXQSsomG3liW255eb5+QUsN8rJXj6QH1qcl0lJ2GeYyWHEz0MftATI30u7WA4h
/3E8EF4sC5e+w9KDKmXTWHKIbh3442FmIbaiBxiVXrh9ERTFweTqakyAShUPgLHA
hiD3rnndKp7ofyAwCCv+vz513y7N6ct0Pjr7ahOKGdL3fyuPck1ZOdFL3q0dKa5C
s+ITsx9TF5E7fnkwl5Lg6uRvWyZc5J9V8kK4Xe16wROBT+l3O2P7Nu1JKfTNExoQ
x/6l3sXitMfgCCKvAYzO8ZmcA/Ew35s+iBKnavyDqb1EgPhxjZB6ZVfvcXTE1nCP
Dm8j8HOKi/VfN49jkbsxH2eU6hjQdZxVdQNH2hmjIo5hM1ODUgvv/ak0ED617Dcj
o3pwqzPYkWiRzKtIgCx/28UZzJ5quJn+hf9l3AfUtPHSzF8d0tXWAdDGsIBXyFN5
qUWB6U1vSh6X2jrNmNFm2mJJY4Gggz76F9v46aWFeR+LDZsPHZXhgVX8u16Mp2tm
KxmGsp5YB3W4gaIf16pFSDP0u28PHx9IQeSbR8e5ks7dwPWxb9rBFej2fy+/UzXB
oA3RuUIrg99VW1ZPKk78a8BXcZMYkxpt5hCw4tltjT1aYtGup/r2sPeqHnSYxami
qPsDho6EEgwR+nHV3veGlSrQVYlUJwXhatdH2pBlyWsSbRGOnOqW7KTSM/8wf/Sn
2TL8xXuhpN4uV5GUvf+4mgoxqZqL36MRDcNfJta/5G1IFL33NyuzpCSkLlYZkMmU
gJHcNQnt11DLh5VMRUvxFZ38v2oWde5/ey+aXw6ZTzLBivrLnLDxgwJyT5pU21kh
djD689fdjeiEa+2JfPrgU+uL/ZcOfZmC6hkfX0Au4wTJJgjaxxsoQMgRmKKFBl/1
9Tc0hSvqcX4Ord/IW1t1GyU76wsJXp59WXGbl1Zrf17A9ow1DQOynXBVygfkARun
YYqKW7ABACaqG8xpsBKSce9JisZh8nicBR8vRjTMiGjoHYTgp3Y2urVLJggDCGnq
GvIyVjT/gTuLzruyPqYsZCzuFwYMa8R5sU4Ou53J+z9MiaxOUDrHI+A2wbGhGE82
ijgR7clYN7onOdD4UvJEP/zA/bVyMNXVXx3OrDNl5qkNlJhICRJqRTQpUjTLj09u
7T9CTH+AbcziNJwbL/+i2RoMULDvG79K/lB8KEHtpJnZ1UpETxenkpQG+FQREysm
8SnHOk063gXd22je+Qfck39QRPv/xdtRUo9oEiq9GDbFZ20itaVI0X2p4Fxn4Ckn
JNg5Ddtw6aZQdMNG4I+O9lc1t54bwrWPXs5K0wJhS01LzY+H1HSsb7IrtNdt9skQ
QH4LVjCXZSnh2bLG2ANvAG+ZE/tcRvWWWWAKIvQJA4qPtwtv/8UEGpYQk+WVXcHw
cGbFdL+oi/V62UhbDE08CBdaER6hqmIKlj0SDBb6+Mq9SQqITHL5aZpGQQbjRWhl
vhoxQAHt9aksuBtTIu80BTgKnolN9e/Rh6W2OgynbdPWxkWv9SqrwQtzqoG/tFEh
R/5zqwcl89GqFdrY4+a9iimbzO29DDy0k8+1lXnMUAriTPeVz1E4gZJLv7rKrrVa
9Cuee9XpbNWqln6NtiV37kqPcec+gAshsIVsyrR2CAKeiQvVt5bZvrtMsRDi2J7y
nsjv7NoshYs0VUWdGyGDNucx1Sq3yz0CsSoFVhhdDICJL+y9+oeHOHWluEDeKFeX
qcwK8MmmCjY1iiaJwbQUkHhWpaQU7Yj14YIfPBNdj9udQfw5e+UTAmP6RmreDIvM
I+xD/Z8KifWwtmdyUk+w0WQJ2xTFaJ1HffQAvZqtdyQL3UUbSqRuU10obwuFDxAm
HinErbomxoJ60GDLv4Edz+uXY0yeUxIXE5/zntey9mFLDCESawOEUwky5Rge9L/K
vLY9rtMKj4hVMJv6o5QbMKAulJqB57QSZNsGUbZQeH1fmtiTRbVsHs6R08QMFeiM
tBUfyKBowvLMWfaKNQeNny7dZi9NahE8W7U5vuDpjS1WMElRAHFI0MlaKKPbYrsP
j7RluON9nVzRyV8hS3oJFZib8S0RAmEzfIJ08UhTXJj/gWQulWVUeaVnTWfr9tp2
CeEt6oNrvsUYC4ZTEE9+KcXXwL6a34VKSgF9wxh6YVnQcNSGZ7QGF6SZGyzKJA0O
xR7aJHxHKlVoBzqgmsLweoRI5CUTHniGGKb1O4s8LfXS8rKgMG7C5JGepGCI6Au5
p6l7w/OL2dYvzo4DUB5vr5YhiisG30KkMWktDdyxRZpwiJWNVjsmjhuQKlPQLGod
SavMhWdcgol1qnoq0kgW9HqMT8cuHiczUBmpa5+NR66gIdCdOMdsWi2h5z5DDT8w
+JI991vYLaRZZnUwITqIkPyKFrE3HbhghxH/rRKbePIt/AelApP/AHjyn2K8eMWX
hnRuEh9zNsJsoGgZIFP3tRbIslkvxOgpkPhZA8+p+Uilzd+XNyayIiSElY3PPAsf
FkP1sLQ78qmGxbXvsKNwrX/9RdE1qpbGd1j9d7wI4/93Eo50EmaXUpArI8Pj5YZK
NMK21EDvE1Jv95gZNaqgi5e/qB1nlsijBRCswZgmLv7teFYDWsoiMZxH2jwUXLhS
mpc/4d6LmSHLRylv/YLSWC3otE4yNX+SZoU0uc/XcKxFupAEXLebsreS4MO4uLM1
9bA7suq7zGbjc3jzVHuP0q4JfZl16QpQiSuo13dzMoc97TGSA6iPEL/nUGh47Mum
MfKoo8LpOIAGEcRvi6pjDOt7BHcsbCzQ0gGK2fZyrEUEhuHjFg8Tt8R7IpvUI1lu
su/Pz8Ho3RSRHV8ovWiYzi1P4Emu11xgxIXvgJ9rRJ+hXvbhv1QJnUcaJz++JAep
VUXmpAgq0ZZmGhxw5wHxynkOaTvSw+t/AowknHeyrMj5f6snIVPCIc+AUX3/z5xx
x0SHUe1dSrjZupSnf4Bx4hX2TuI1cC8BlSY9fpUW8Ecn0sOwz/uTrrRHqC3tmatV
e8aTQIk5yI6rcpJWhJ9EKeNTc3CD6h1wT54w8i3zyf9NIex54XFfwGp7DX2A6w6a
YR4ILi9HXgD0s8v0gYpH+sMUrPDzjCDlv+SIh0YD+YI8eaQ3fEP1z/2kQx5AAIUM
qwkBjXz1Lcfg2Y/CU3+JHme9x8bas6BO1aqwvzhg93fii7uDi4G3+WvSsIzQ6K61
UkUBCI8zNkfLQHXk1l4RMSk50YEEtXcJNAHD+OZGIP6D0CtY1YJQSwmk5WqQDjh8
xY1AwUR0SZe/aNPXA6wpmlXDNZUxti5Y1UP/hH1mPI8WzdJujiW8qwm+mFwy/rVu
OAJte/i76WYh3Z/O47CkeAgk5AVLeV/IQ+G+lBQIycsGQD3FlZoPbTY73XSvtxue
KcafwbrqVw5Sbjd43CEdDHnKCDKEmBVyVCFBVxJ15DLRedu2b/9Mw2m2g3SMzHEB
xCsSfRLI75y9lj88Z8jkeqWNbEMTF7vCMwKCiGEW2FfJ0IEg0XYRh6DacJx4pm9/
3ndSLmN9wPKmR8woc4IoPgBMJCJqZ+ego/AJFol+Osb417mW1OwMB2sX2kWKMbAi
vxH/jyAqvEb3nwPtgZggi7fU2hVrIefF20qtmfXm3COSXsP19lx1OiDBv5w039Us
c0O1ksQFcg6pLcF46fZU44BDZkIAi1RfWngzd6PRTGhkS9UoM/WoYh+3+ZZ4RkIb
GLMHNfO22NlYVuXg/AGRZwljCO74LhfH8gADBM3xC0ITKXlVQ96XLuAcriLCRhI9
okoMa6PPJfZU3aeM/rj9cm864XxSbJJJvo5eXN6/Zz0NKnjXoIRPL8jTg41gce1V
EkD4jmsMWPCKvBRwJjanbAOktnnQB+nX0r4j6RrNpLR/HYXsG3xgggsTTLxEzChN
Ijd7hMEHiOiAIrc6x6RqTmHUjTQiABkSVQsWk7ttZRLhR6d47rg6IC468/rO0SlH
kbhKfr1+I0Fc3a28wDQmqUHSrNEVghqH8CQm/bd0HQItwC7fFWNOSBhoiuhnLFNO
ENkeOuFxm0hxyDZUqoH+cYumZ/jn8wU4q/6SJX2DZiiPYccCG3ns/H7TWHQLlc1s
J1iZqxV5KSvpGGVUJLr7IO0fgySZ6rESAhM+bFfVv8QQUDtS0YWHpeCIOQOfPEiY
4bZXuFrT96kB9OiunSzhPkMVZa7qRHf6Ga6kIHP7oNzWApfx1YOJlTgDXfwcIfpL
uAsBnbGZyZFjq9wnT6JOliZ5SrzDhQCQWkKesc/Jg2gZczcip8xejgD3bn2qCXTo
rsyG4QnDb+H5HWCoULAbG5cWxdMRTlj3z/N5v/ZLuWoIeeDFmNvcMbH3VcJtICPH
JDKopipF3dnrx5L/OmzpXrqeFno8A8e7rpz3qL/ZQnDL068mdAoSRT9UWouGB/je
teyk/cRjdPOih7HlU3cMNuEbSixYyXrLz8um3qf6IxSX9zQ1y1y24/PbeioPupKP
oICOC+snqdXqpa/SD+l5clHUL9YyjKa/J+hiDKbNk6v+OKF6+PzihrrdGCWKroEp
iZ2i77hhIl5ucISm2OE7AStLmHB4Yf2ZyWR29pB3xtiATAqTX/A/MTcIx8skJEFP
OoefDt+omkvP9LVc4pINkR6h7i7SSS8Gt1zHP6kHU25fKJpJ/aA0/R0GouhcYdc+
dPf8F5eH2wmYqMLF/jMeP54TttIMr8EYoPyLpwwhdnDVSsGtnp6G1PLGzDmByDR2
gt+zAU4K6+3KdjSC/1oLd/oMhbIBC1mLiFxAnljcAa6cYFbXpEE4ecGA2HWxzl7s
ftcNEpD39KMSL+qykHbgGuTxP9hpk8YZNZ+C9hfW7LE+VZrxkcvZGoHsSw4KDQwx
vmfn87EBKPxGxJDXVEdt3+EEANLZiQetoenU69AZuNE3IY5VGQzBAvYIyzWzLOsA
H62TJYLE2kdnh0YQfy2pxHBcYXJNGlui46K2QuEYl8ezKku1x4oziIu2aCHK5MO8
hfMuGR6YpkDQJNNPvUe+Qqzobj+fBKLyiH7jVS3v3VcbiJPAGm5hWQRbaGiq6qmp
cwa6Ef+tREyLK1jkn+Zz3CqPkzjdbHCnTiaq4j6GcLLeU3RYCiZrEr1K1jYbT5Hw
M06eDQLSlwd2el8uI7vIhcazJmU21U3ddnCGesITwV9nItMHlsCN7g90QISTgrnM
7eD9hYvmRS85QEDTDK5h2z+w3YQCvKw4WnQPrdXhRJw+gHNbUIDgnr06KXxLTZRV
mu+mcZdZOqdfx9juqhikWtgaqaxUVuzecKosgP7THQHASHXYZw27HdHjghlS4ZE9
nY2YY0PNAm8skX4uDmbp6wIfyZL/IGmsYh/vHU/mn3Z2aNj/NeV3rXhH7oYdh7Ma
FG8FVUsrLm8wbcgcPVC0dS6d0UCSmEvN8aEfPlJV/8BNpA4NZd3fBcO+uFVbu70d
XC6E0xZrJhCJhPYgoj+NSUnq00T74dV1NFOireWnt04MMf4olQNIpenl+enMwI3D
iXkiJIALW6SBi/16E14BvuzqbEmWlBHWVdHFIeSevH0kS42eowzQJej8BMarLYOT
Fsi5sLhZ1fme9MPRu8CH20rLz63LWLU6WrOBBMlTHthKq+JVXRIMffwPRT79hDFM
pZ5BoRUBPU5ZaPt3bFy6kLxydZjiZuU04EkOPfNdNlAyVRzZZyAnNTLDQFXkozRL
QUIS6stlaAbHJtNIoth8xDzc/gy4ypLk2SdCimAStJLTxGNCRTtdglHjBj8+89Kj
uxI/OIcRk0iH2yxFc3P8blouJRFIUmp4DFeaRn968ReIYjlb83IjnrDD6pupeKK1
t4DHR3L3jd5/7aRMphBweEkN1dMDhpmjKVN+1ckZSzOPVxXklIdzils24C7Ucm4N
ufDgd+dq1HiatMz5QlDZbsneaQLwrBny/6H41l62R3t5NL/+g+ms15noHXPjNq2X
gBeGja1ZPj6pTt9p9THNLKUjs11G6T8lfOSPOvnFQxt4aaYyVECyXXQZxttNhU9/
kjE8l24l+Uv6ACSPSYLMsYH0fXPIc8gtCy/m2h80gUXYAujhhzaJhh9G+Yotk/BC
29fTUSc85PgzHdUc4ox0BobrGyiYDzR1sqh9M/b5flvUNQZCv5b4kCdqk2Suzyc8
TD/PXnIGHYZCrdTDmlVABIGLy7drseSpIxDDOYudrlfQOUDUgfkJatIfzrK5O7mZ
udlWWe6aq9xko0wT3TP78fruI0ZDe7w4rpIWto0E9hTytjHXu16k1N6BjNgzwD6n
Fa1TH30wwAJAscSZzw9pkq/hstGJYvCxQtThqXt/yWWE5UHpzM5BvtKRP11zqE2o
5+PHSeCzxjF6zC0qZokCKRCOsWyaH28RUucpZ5WGZrnc7pRYLaPx5R48OZnhvdTP
zRLRjs8RZV5K+YbpVayji7omlKejZ0rzX0O3lrp8rDG0kJwzUX0KNrZsjUBIJg+2
jrPeh3DcPHI5aet5rx2P1tr3isqiEmUFrASWXXBLyGsVapg6k4Rn8F4BD7XZjWut
eOry4Vk17X8rHvrYFcCbRL20faDzQ+WUE53MoqIUFXHZ2DNHb+Ezw/l64OQuj229
Rz9OyrUTnvs8gP5OWDHwUaDQPvgeq4t/BZ6V6OZel1GVroQmsnbMEuIDwzUV1679
xmgTg/6d8eHz160XnptP8UxsG8qAgQiQtoPed5zHhibDjX6MnfppeK8qyDsIYrmz
E0trud7HMhIWGdqAdzrRajAygfb215r3mkNXqoNfkvpB3ryKsFvH9nf1qzhzFUIm
2qRZk6pHs1CrJKxrJQ9D9x8efY9RLj8awlpDtqNQ6Phj1W8HTLw93+2bdQm+jpFJ
P2mnTGxqsSB8Bq87wfvjpVeTj2yFY20Zi2Xah3u6cwNOwVKf/hASuzrTmM9zc396
NnpxmB/gUEy2/+VXQbeKWWjvfYkp7Ne4ugnd9jgqar4otDdOBIlWP/jJOxwtYwPK
0phmNtF0xN4HljoIGMV36r5fue6gtyoqawB+xQtyP17H+ryUpFB9zirz8Cbx7a6b
jWx16y4w9QsHU3leiJ91nzjf+ceAfMwaFA26LhrsPWDpiJJXmGWpMboJSinkGtPT
lVw6Ps+Lru/kH5kS4OYoQ41KpkihNxa6H7rh0tnXebeEqTQ7sBYSmOSurQ+3uHMY
FalPQtfvZlW6pVC+jzPM9a8pTqQRMgt15DrbJn2rEEmOjsvwbMGPrB1fRqLsHXiR
rXNBF8zvPM/hZL/NtaAZmd3GQCrSI++qAYIay1ajveR1m5T7FS0H3FaexLwhStE2
fXjqX1/hOhB5ql34kXCBz4zpPKhLN+YtH9Wa7iFNt3/I342E1mZKACVSRkAdYO1R
X/xj2Ap/vShQheZryV7zGyXmgoqeGM9aWpvZ20W4BAsUdsAG5T7U7tmdrZw+wpH5
SghctA9RHPmFMeD8YvUgAubJAL/ieYMcUckQ3q3OJSWxg5Nxv7XjA2mFiYZDLJCw
WX03hV6qdFQ57LxTwTUaL+mQWpxhubAWqfbE/ZB44ltWaCmlSBJPKMRto+qNyfW7
l4zRndnUAVcznPD3PJJ8hCt7P1nfqu/to/2SDblyHOU9XNV7yZ8q0LUE9hzMKc9L
7LzbUgrsYLQD8cwbbGLorGI/Yhg2Q/j9NLrs92+ZyNE9+EuN0lNZs9IFwLUUlvLe
UueZs/zmEZnyn5dau93xxR1PceBSR99YB5RmwJuMalWtVhlrV48VpT+xYQFpuWmr
lXWxnFebxNYf8oeGnxwfoFiXwdFqtyr/HImPd4NAMTqQ/O9EMkGHVT0v4zSBopB4
lE80TgI2IXlS/eIenhTj15Nb/BSskgoLcI5jyav3WwpB1DeHo8vBDEFcoT7HHw9b
hg4e2AwkzQ1Foc98Lp1U7fEJy3qH3/N09uoTdJj5SrRLyNn+3oy7OuPHdT90AcvY
6niBAr8iahypnEkMn6KAEv9WO183haDoT/vlqZ2qKTz7amhmDa70y9i1cc7RhDnK
G1+oQcW+fA6fD4Yfsc/LFPBDKP1H17w3mWdH/U75BieTTkakeVdeX7WwQMjrISsV
6ZXhS7JFyl+dVPQI4K4gm9KC4ttey2Hn+5pF/zQnDWfLS0IYFJOsABl/nAtgs7Ys
uCO4rqyX2DJ7qH0OsZ0hdpWe/Tp2hC73LBeKhTkqsOg10L9gG5B4PJsZ9refh+Iu
Sos+sX90BHYax/f4x7Qw8Zt7zGVGLcvrmUlL/WBF5hqyHfmnP8nhB0+N5yYgJbvs
1S11ZXYfCy062UGUSCcu5/ytCF0pjy8Pqvu571sffSjZmG6kB3Yu9/ujxahHoKdI
emRo0mKjisdcoejN+sJtnB87l5n1Po0CPQInSCEgsi3iBKba6sPcLUmWXNlUMvSg
lnO7Yg88sE7RBi/3eB0wQZT5HS9I55EhGoOKV0qYx9zcY+oP53QHw1nVFy1NL/iI
mtbaYwxpIaK4B9joB7i26Wo9rZ3JE4L7dciKhUWaO27Syr4pY/8JP1Tt04h+ggIX
cHSLizliXGnRXC/xOHHvrnc9VE8zJayxDCGqEa65/LqTRTQuW2f/L/xCFuSKB3xt
X6lQUcR8rEP+6+0VP688ANY+1PKNLimyg+YQp1OY7gbtLLWST3pNvNKnzKT6rB6j
hGg2iSPzr1UKDSdymgqT47F/qCrDMtp9aMH/bSGIS0FwlwmUc7wLbENv1GuptB1U
7Ky6bFY9ZUqRaIcZSJ+TSxE4g+h5S91fk8EyAC6e1cN6zdjgEkOgFFOuLxlbYYSQ
jMZzNrTwuQP89zxGGJYUDSO+5AuARD+7JywvuUMnUPcXjjARMPYrk1N/HhbhSwbi
0N7xMFArKUVzTgik+Slg1lcxWY6UB8OMzWiaXg1YRQR53XfNF+UzrbyTgU0+Pf/1
IK5Yh7NegapN/RzDL+jHzEXN2b2Ksa6kOCP4B6yieGAucszbGqRqzd9vjpIsqMX9
ux/kwWvxv6e00/0C67RUAGDd8B7ZJsHziTOlRYZBn/4i3/WGNP/mfjPOOIONYkYd
48aqMoLR/2b8AK2hOYnRMDDXKozuTNVLOPgSPjzYWbSsyBgdC+oRVst7Vn6VRgoQ
qVQL2LJlO/to2v0f0v452+2wxtwEosU/v6mJSlwJsv/vsOGBxLV4MjajnngIhs/4
iynUQ0/NeuZxUnnqN+DQOZt3QRniRSjvXqdjTX4g/ghnBrt9zhAylDWUsafG72/i
broZEdPQL0m7lBTS1AWrLKQxXGH6mn0FYtUG7PUGOninOzUVOfGdBZhUFC7/a6Q0
nAYP6oMNY+eRE/ON3JHD/0eJ5gH1wuFOMcJf3C5QKyMbOIqU6m345BFkkMGwlqzM
d8F4YNSmO19y4kwxbPuB6CYDweQSSCc9EvrgfMDuAooTQShO3P0gK8s1MSebkxdT
8LzikcNmZcIGU9qyuoIDGs9cdwr2a29tj6xswXRcKA1/Qj69uPk8iFOzvYwjcd+B
6T29u3mKYZI8i8iTwMXHtDKWXcnzxF9sIbAA0w7nCyQIPIzW2iPnfv/EcnSD+zyV
go8jm385v3PIKG7mlfPN1AcMQMT6U9Vgj/KtUWrVqz91EnH8CO0fZcHtaZWrc9To
n1SfoHEpJ2pifhW0UUzf/iSnh2LdeqcdSm3l7KYFiKzyMEBjyUMT0cxSMPu46N9Y
l1k/Zz63ek2+0ESTrc5wFRWAy8SSnNfJQmaSLWtVUsQ/DxA8cXb0zQ44s0o+iNjA
7KYBfAxNbVDFF2TG8qZAqZs12lexpc9xAfWEiaBmGmT+cFzHJtGu4E3QqhjZeP3b
ROXGG57mNh/b+CqKvAvulLOC92n5d1mdWiiWAfGXaQmXPRNz8GcXX6Bct39ZEmbp
stB+pH05AdmLPsdyWUnLo0mrlh5FFuExPJALEoZu86O7QkT70yjdYxTdOGJWLLJ/
3hdj/9Y0r0IQEF1Wifz3P7jxFHDzIKnxP7S/LgfPaFKYXHYzRZelDUoJyMuwnP85
jhbxAMUlxnjG181Wph89HrgOUl+YM6mDzo/8+y7P10yIP2ORmuoJe7M39m8XWDqa
Y3keF5Rx3nO/lQ+qDqics2aqmfEN1xJHrUdHmRPJUCus+0P+ROaTI63/lT9H9WlT
aqIFy1ZgG+Lc55/WSkCbxz9sF+1ZQ2mqeFcsn3EYiQzn4T8qOBXDY10REys5mi0l
EY4tVWPOlu5cDF18oBwNmHJEKD1/qFbmK1fkw/fkH3GO1JkkT4F72RgW3Lpja29Z
Cq/iCabyDJwrVeO9OAfbBYNlxVMyjDaQCBKF7O5IFZia9TFlu33kXcH3r06mLbfE
OQNQl7Zicrs5rQmCDKJN/VuNQ499I8RaRjLR+FaUnTGqCbCLK4Op8tmjswHLt3ph
s17F1XrwiZgvEbe97WEKGf+tao4L6fpuFxLf7IVprs8KKt4ddlpYFhYyCsoCoGUn
BcMDJSxyMupvJk/cIu0JwN+kYI42V/l2q0tV7WQlLojzrbIuk3BHBL80zWuTSV4u
l/tAZ1Ioew8OGBX9htH3Md+Gx1BLBXoN4rODzfAnEb45izAfujIkYg+gpayTi0P3
/kcrQ43XFyB2f5Z22Ri2ArMzDrPTVIfinJsbrOCJ1opecJyoviDpwZTqyJ4r9jlY
rgxzRAQceo2m6EN6rof+bM9tsTZxPnaHi4PRv/4Qf+vd92pECrSPvMCVZBH6EaDX
bM4Kn0XBGrk0j/MIdHD4hBAALGoSyigI1B/LuBx/lxeKWkwS4MnkDHklfHQgH15M
Ea67m1qehKNuqpg/ms9Q/XSts2PB4uh410z2ssWwtQ8nq5Jz0XNuuLKT/s+d+Fgi
7Q5WlKwB1QStDNk9a7GHncXQdQbrGAwE85gDaQM89bTFmsVlXGJOsKCn0374sJxc
ts5HG1gCDUPB5Ai1FlJE0rHwV8l3/PHRxWFm2VoYbLXSDlvZNN3ixaT6VdphbbZY
e5EJ7Vg1UwivmBrJFRCEuviEtUyoxu3r9TQUg3/NvaEHd1UopOfDAcj7wjI7P7xN
rklrikogq6TbYE6urcqcZAZb1TxaS2iBfTGAauDqfv5R7bnv4WMhmbmO2px2lFoM
EGJeLTL/0CDGU+QDlxXh8UdKKqZ9PlAMmYd8g3xEtS/8HsW3uIaMRgJLjNtAIbZH
4bunNt5/PDGFo+QWR7sspdqeJuSvyH4VniWlyU7PKtx97twjNe9UP7GdhLC96WOI
bngHaeZ7UVP64yvfRICHYO/WbQNNqoBHA1qqOXhB5Dvf54cDsg2Awh77Se9oc3v4
QJU0WerG1KcFXhOW1+kXxmV5d8VbiCqzSH0IBSu0XOqNgR8J+Y/IxXMVRB7H22u/
FsedWDk+lQM9zMkknzH6IUsVcAcVx+TsQH+21OzY4BBXawsLqrXsJyCGFnxZYASb
CV57zqY76JDs0e6B7KiPnC9C7P3j9xh/EQIXKB3LB7oq4IowIsSlbQPX3aHVVPJo
WtzEk4iByNZVAH7mWTjNOZv3sBimYj/T0grG3lFmmHcugXGVtrt4H41E36l0v/Py
FIZLidQ+JkzGEShygoIktgpecf64bAaIwQTQX6SlHHwsotzVdctflt1LFSebYdtn
BIYxqMZQAuSb6USBJZpYKNNy2ryuxG3+um1E94HtiD70iXpoIjRHuxbftgqqc6a6
S1wquBzUHeekbv1YDY26JM024A8T1CwUqR6a5qrGMJzWq8l/JFAWAYpx642hZo/Z
ucHYdFjI/Y1FI86kT94/3fJy3NmFW0Vqd8Ni1mmlplJj9x3kkz+rZTcXjA4UVqJV
pl4paKX7ViVaDMUuxTtrhPyWfMLvZCwKnThwyk5LzgXkLqnbwkZgTkUyFMa4fSeV
t+MKnBm4uLOqHuo7omON42ITbEa28iQ88X2GCEdNJesjL4vc54TgCLBXW4GC9LOI
59ZsGNwk1Uk6jAQ83hjZvkC97+8DBqy66GwI8eAkNaB5DYAkXZ1LuNZqEdjgY3Hf
YIuPcXqN75HqQQWUQhZ4mKEdS9UViEt6FfqbmuFCpCOaULrqmZDFAYnMifW1JsZC
aiVVADdv3XzjJ3rGS0ceHw8+5XL/HFUDWA+GuCw6bOka+4vX4CT4OirYqek1sl18
qDpRI4Z+T67kbMvgR3hdDSTTWdIk+QhCkEYaG/w4qUSRSyNkKQhkl1225Z7PQik+
3HlYJLA7nj2SfLoQzOLfx1FVixipk5JWuzci7Db9mmE4krfIqjKsaYvC+4DOo01O
yAdWrGLK0Dmm3Blg+GTgeYYI/bX0Qqj3+PMynb1ihxGQCANCf27+nErXuDSLzQXR
wDR8x8lXgudh934iZ5SVhX1gd1iH6c/cG1oQvmjQpsoa7PO1TkRDJgMzyg3sl9gj
EQXzLBemY6dsylZ0F4vWKwVGX4v65pcUlzaID0H76Eg4GKRtd635kvwxJoaT3BAP
TYtY+KIPWeqxt4CnjpTQH8b/ndaGOubtF77wohnXVosDVvPOmAN4kBpyBqy3Eofe
CC5EVrtM/0y3ayFIoSk8IdcHZlEOkG8oLtSNG6NAckXBRHubJySOS0en22nJILbW
GzGCi37SaAxZi5CDphtcb+3GO4l1iZUnX+gbaCSpSsuQtN7ZoB+2CkWB0TfvMIA6
rjaKS3/8FAGDFbd3T7+m+P1CfBo4LCy6ytA+f1waZo33Kd8YBVYXjT0s+1Svgs0L
AvFqpFokEi5IVuWQB5K5qSjCiTjmKjeh1FnBvER5K22vGeB+mJ/Ye7GXeoXtBpfS
FO+5yK7uKtsvPCj6rycniNineGUXzo61ff+IjmEA6jydyq711QF5AIwU8NGlTw2/
Ulm+6m3I13r7aqpep+zsQidAzLu93eT7wlaBPipK5W5VL3jOlpyXCSG10DZRqCcH
CMwQqdsuDoSY95zLsYPUu79m3rAdC9ix7pyFHEsXcBPXib7ZjJ1JOsC56lDD53R/
zftYLFAfMX1pRFo0zVjUi2RB3eRdpUdkvir1DgYZlYn64fJbTwvt8HByeCwvOuPY
dyZDhMa3XghoRLPh51ahUcIs/bpq0Slt0m1cqtTB32FAXRlh3p5IzsbifWwW2c6l
7a0T1ziWGYfLtGgI/zbAkWYw9+EfbeLSACUHHJvWp6FjFIb/TX5ghRh3mEztxuAI
00p4snT65yhotQyh+OS0PDHmWXrLZy6hXB28iBnVcFgmGPXXzMUdsu3gPdj4KG5t
hZHjyFnGi2A6qqSOYNaFh4TpcExMfRtp7gEx4BEZQB5H0rCjzMmCFibI+8XA2nNt
9iffW7mmduStSS9wZ9DV6yUGiCgqD7cb1M+GKW+PePmx22N1s5PtHGbTm0+oZ7Nt
CYbzloeVEArqsMb3rVbAHCdjhIjk1K6tAA7BoM1CJ8pojGTal64cm34LrYl+YiOe
vvAyZwPi4YU74Sz8qD+r85IskEU06O2wx+Wy5pVZwizsnsupGFIyE1ZzArTUj5pw
rowIF03+IcU5U5zJuOu5stFvTfn5H1fUC0LMBmcjRavKmj32+RKKm9FjBhE5JgqK
0p4jIlyaEaj/HIg3wl6Gtg6GfO8mTkJ5Lcy4SHbU4FGNGjyXM6EWZAjxq/aZ0tzV
heqxX+OL3WJWhLuKSdolctoXdb7SKuvK6F3krgQFKLqUiT5iu1MnR9P5NIjmGEhV
dXsECOgIanI31m470T7MdCz0WyS4WsL4pvvf/9+s0gafB/JVM80DhFo286rYCqft
wwCuPfE8v2bHFcieltPtmvH+Yyxa4IsYK1alLsml+I3GR7ORHINTFQu1oRORczNv
VlPaSuN/MULZlFZbX87UJnWFEyUiI27GcmlwaJwFVwU6DhXwQm1OSlGjIMUWIujE
FZNDb6h0xXx11xI5Q1RacixPFD9qi+qI+h4HLWLN0nHe1VFVr54sMkUss0t5dzdE
uVaREW2dGK0CdCGp68k6oqLkDg7900PYYUGhGnrtU41GZ7Qgjx8ShnwcUdLIsMq2
6pfvUVAnrpBeD4JMQnJwGQCCSDS7QLU1yj33dD3w6Thslrfq+iUdJlStknKe2A8F
tqK3+CDrT/pFqrK7IlwB03i2DobJhmpoM9B+EuDhX585OrSBvXS1FEZ88q4DXXV6
HNhELybD5dkFmlPtRzu8KcPCMgwTJ8419KSARBYzJUZqUa9+kJcoZYDTESV0UDbH
iiikKpYoebDJ4UM0Krk76KybMWaikITx09h+Z+z6y3lzTXaoouGDQAfhtNTo2Mnh
R6X+asDw0vHY8tlt1oB6u+GT4Sp//hQXGUAf7Cqq51nrgptLOoge0CJDHuRUeohy
upv+fcrL6GtuQo2mTqIcbcrTyKo7VAir+JLiO/p+mSAipe6p3IZPXoo+plk1IPdI
0jGLGCKWNVeQ0AvMrnNc7JqKNmW+Znp56dZE9YiJ2I7hn+5S8wi8wpXa8TXGd9BA
zstqgbAX3Ac9gkU1FVABpxvALKQLcMuHqlX6ULBdqnvl+27wXrkStxVs/T1zmhEJ
cXo2yW390iNbGE/mKOtIOx2qwUQnFytYnmZgQY8X4m8hjv8scHDSkOckXG7siXNt
+0fOC5WyXBN/z6rQqdhP0HOL66r7Eppl9VH+XZ7L57m367pUVuxPAxelKyndy/71
OrwPbPfNm+RnNFEuw/eT17lGnEfdS8G+102jZ5Zr7pnYhZKkAx/dpFKPOFV5fR5E
bbgzupb+S048uLuEvlDCBI7BuyNZONK3KPRnj6jJif40ISgPExagxeeEkoC4JOFv
wATGeEGC1TyUFo2Xt6P7phxA3zrwINuPOwAW7rMLrXjHJ2kZcdEX6CtMnVpFc+3m
fZu4jAsl8hPWEsCu9rhuO7+pQMZLTHWpJgpfwNPFYpjrUsfVNFfx/H5pEBnZUod+
4Fq8HhKykGTEQqxW1UQJ1b9nqF6HFSgUT3pJsZ1GJ6yooL5HLD7jwnPlnmMfDTzp
NEZF2xolr0TdsMUJvalUQFHrBAGA5698yZ23rkhcxOynDGYSR1WXxzB9H8Cjgp8t
RPvf1KwysSuSY3dL0N0ycs77lyy1fPuUANpeFYUAsiSr5e1WxAZPsv3F2cGERNVa
yJJhCbFNJ2yvyp488yuuMxc2oK1hdRD4BC8LtedsIFW25ayhrIga/YISyjoKjOa+
rj4ZBplNvVhzLkZOa9gzSlBxJQgD0LE01sGRNOJC8IYkA7/8kCOz+fV3RJbYSZvC
Kvi1CVFd3h/3ybwqJb8ZLLi1A5mEFTsHHGmjbqJsc7W1XxGz3yHV3+KDhqOgD68t
wfR9SOw9NuHzAHFaMlv47qgX+aywHoFQWhyf4TfPWDOTen7I17saB8Rgp3pIyLdD
xgg3xuO+jyfNLJtn+saa0AL+5lGs4UeZmK2tr01ASFTSYnBYja3RWVmNSlV4s4oK
tOxOe741/npW6JdUc+vFvAOHlsRJpRvtcgEx++wXfdHqQanQYD+YGoX8yD/jJl39
YZRp7azqg6D/hOOLk/S1ZCJ4mRRM5Wd7gsNNfQLZj/Y812yzF4n0lZ/FPrBC6Uhj
zjy0fcsS8n8XfJaDkN9ghEbVAmnbAgVUubCnD7EluOjvATj7mLOkb9JTq17a7dum
dbjpFVSlqXjUT8yGF3ODUjW0lVdFABD6lG6tYuQm9NbcFNjaLaUaCrfQ+eApEcHO
ehGuuHA+Ihl74dhqvZrH1p1tmqCpBMxv0MavE/qTe5r8idrN9i0f0v98rU1jvJEg
/1GQywxtDPiKQwSb3gPThY5YL4M+4FdPA9ct22cBcS4SS2VSgRnJPVyKMCL5jaPI
zZ2sT0OAZWRrIU3eCor5KxAh5xpSAaaz//i/s/ZSeg/OalOnEEbOyVQ6ugOa6IPf
J7rG7IjVT3iEt8rWfYBT5kQYTBxmiZ2PR8zNRe5gwWjoGtory+nDdBbsuVZsIPfR
p8GfIBZkHv/jdsfdUj+9/bCdN9o7i87fz7x2sqxufFp3+bS2wa23f0DcEGRMH7aS
eYHKTCaw5Fu6eCV4N5UIN/FGNoooxisQZm3F+O5jq2PT5+eYIrJ5fq3/lWT+UDiR
3IqFt4UUyYExmMEjsKPlhKa8mPrU4Wq3tDYHN7ReGSH5AcJ0pcCfakubEiLJeGqR
40i8n1elEq2PgIskkdH+1OuiQ+o/MBYoLvRQs1I64D4yvhrljOJDdBkmGCsaIb9Y
nsPMSukJMXyoge9OONJA+vQ6YP8STwvWngG+TKuFEDrwvvJxAo4vx52ZhOi5gPca
dJQiNGr7XuWTnBVL6p8rJk0JXrJ8m8ReJBwESCk+pVQZgk5rCkx/WTeS2Z5Xbfv/
VlikwBCA0+Jy4C0qb50OuqdTiw3DOz5Osf9kDTzI6VplwyNQAtibdipNGjrfaxZF
fHwOtgZU7unTab9R6ToGTZvfn9qdGvvjHAechg7CMtcYqxM1Q89dF4U4y0goBJxS
jUGvHMyTqhyIn95UIOhTR7yXIwaTNAqE0WBOUp7jkesT5qzA9R+abFzlMI6cNuPW
BZNBIvM85TJCN0pwkHLug/MG8GK0Zln5p4xHnDf0Mw22qf5D4Za+lsXUOvKzlIrA
xD25zj9RVDpNKhz6yFyPYUlYVLdnP1ZNG4xk+HKVY6WBOFFks899UCbTvCJ/XxhI
jHap0MWjTIpp3KMrsZPTgiTE8hW6epniAhsd3K/LIHW5ZBoJS74jbDwlX/moY147
g6l1WTNNcofZ7m4NWHbSA9rcA/wJUDvWw/iwoNgL1VAgEfrTjq+o5ZNqnTGkGrgf
FISvLZzlWrNomlCCKQhSBbja3HqHLmqM/fesbkoH7MWY7/dgACVd7HFQOCj3dB6K
uVIds2/IGsFQV8IGMILMO6B48mDUzPyAp2EXTyD2a1GVAghomiffot/9sOKipTl1
7N9KBLywuD30F5iUSRc3AUNv39xt6Mi0d7cHa8RIwEbWAQEpv8nxEdwCj/6zXfEV
JZ8+5Uf7GHPfW2n1sqE0hlwn+NcJGn56Wg1v6XVS8Gx4bMmTBzT5/YeJmgCO0daM
uxvceaAuCFenNf4btw/7YncE7XTYHCKjH4gHVHhdNWbGNqJDEloDu5N3J1sYyCRV
dKVcL5NQsGSopZRCyBMcU906U5AL8dhJy2lbvBnyX7tRffCBdrvANCtjwaBNUMs6
l+r2h9ed+ocPlyPjhcdAx0ca/yB9yhKIxY+jZFkPEPytNeCm7/OoqU1J3nevelm/
Nn8UlZGhjBOAlg5cX77YExsXCOAUzO3PT6R/t1ihx/FH2O53/dUUTM2GnCKfD8iV
W5/VOWgAaPU9Xz9LP8Ce7eeng8162shNlDqM+iYJ0T9TZ7pX4zCg3ywv9Zg+pb1F
x/wxHcGMHPSdux1Fh7du/5jmCNctZDed5Zws26un6dFHXLBLk0RhFJWZKQTiv/ug
8zXbEsEgvZ+9mf0gFjtkoUY/RCck1fhN80v3AboicqHtbmeFo40YwjLO+dkB+KJ9
pIV5ontDOxustxMryzMgHRWagkDqYeOlTlTqvxEZibnADHiHCmqt2hFbykfDb/Aw
1In4p7Domj7Yt8QmLvLjFA91nvPKTXemywahuJb0WvI+fc6hF2cheMSe5bB4VPE7
l+rREhhoi2PFhmUeGmY2iybXUEvozjfZtEc0wGZbpbBArtDU+qtfZebpx/7Ms46E
GO64Wc12QGkSy0j25JjYaQgM85CbUlR61f4u7n2zowHmKuE+uzAb8HrJ8+U0GmAu
ieQDReqMk+jzVsNAo0FzW3gNUi61XGFOPeM9YNL1OX9Se8MCzrdHRjtHHYa5ZZ/4
IR7yFjJ/Xe8cukUv+Y91uhk58qXCRoi2a/X77R+13CpFWscaMPQLku9nZQDnfGNo
VV4ugZYAUG/vEcA6ZjcBhOzXD28oiRCn6E0dN+6Z8E8X+BAWt9C/qKl7RZMSY5zk
XUeF1auwS2FnIUDjGi2sg6elShJZou/rAIt5SVU8RLp60fkvEdQ2HaNJ4zz1oXml
/BP2rq+O/hKK08dR3yMerHCxElAwLgGf5+XhPdCCQ+REu7HwD/c3jEyn1xZukF3/
YK4R+G/HlAfZ2oJo+D3GryaZyVAhJOne9pIUcqW8t0/h+ksK61U0yi5iBQagUoeu
kogzOtkz0P6mjwIy3egL1WOqDLSlBd4Wsj7B8EN+//A6xaECdXpWmxl8tVzJ5ROb
ca4ZdGZfbAUQiqUtkH1HwOOYQDml2+0RnHCTBoMRMPczOLXH5lNUHdrAyYETJoXS
mrcVcF959wiNm00Yz6IktMyQUzJC7QtLe/7HHfS5RASDMUrqF5/vg7YGI3TDCATB
BRKWUsnIPTJV8xqIegvHB48YnY9MT8wFJk/PerfdcZ8rKIni9qu1AFXFx7x+oU5s
jNFqld8DgT2eYe0ZC0gvAkEUEDk59paeveXGwrc774ZGfAspxGn/aD0PUzi23LU3
TiYHJEserJpYDjPn5NOqS/x/g/fSnIaLQ2hDndRBt18+uEqT47k2x29jgRo03tZ3
PSeI01/MHmLCABR+DfpuFdT8ogXkTD2pDwGu3UY67UTohbwYP5SRQwVbv4ioEOlq
zFWWh8PNs8OEZgcNZsOWnNrzFRMUD6t6Nw1g4q9H+TE+sQ8jdX05+siC3+Ea7BWb
nEVykq9r5WyJ7vv1tuhNR3AZzo9wZRDLZUUV06ByCsF+XKT8ulf8IxT3/Y565Lx+
4LBXW6/u5olOqrHQ/8p29ODBVUmccDrFi+/vlGufzGNtyKi4xH5JNWT7NiecshfR
IRI3zeBJ1Gw56ordRQSGpLF5BYD3E/piHaTDT3UJQmwOE9wtn25iXHQHOqTI+ZIY
ASuHkawCJ056Ncv4rOmG5VQl4Qu5+W6MXDSrnVnjW9u4ttix57V/bLNGB9i/Xrfq
ax9QIWDfKNzyvxMCrsOT/ERhNSxYoN2a5AFwjMDHZcO87IJ72bZpu+PcUolpykSZ
cqMbYhWGhtkOyqDCBh8HDMeGMIugP9q6Me3N79dbBg2mHv1Nkmgn4wVUkVVO/g0E
wjLhGd0D4c6jaxtyZ2ceJmsBoWMEyOE2Y4Ox0XKmoBf3ZkBsZEKM2ltEHSkxt6ps
+tBPNb3VPB2Fz22CPPN+k4seG/Gg8Z8MWzIkSCxg1m/I3ezx5md4u3rR4CPXiXmz
hscaDu/w6im1oftvUwUxQXEfe1rzFMV66eG00cSAcZk7PZyuOW/CSYHhTWgS13ZM
FDaOz3Hdq1R6JkWE47+lsWmQrxkX76+iP5pSDsWSOG2QeHYaEMe3FuhvEHF4PvwL
PEaMmEBuIg2RsC9yf52d+bSbdnYvmfmk+bNaKxtQpVEYnT5OAlZnO7U00B/cRLs7
Gn1W23Dzvbh0B8s14sgrzvDBTtYj5XosceViiVPSVtz72Mn3kaN74mwdkI68KwWv
R2FFbBmA69F8c35rFcdXfCaGlMXpQZ8hWrcTmi0QUoeJwXzBwaHqO7GvIZUhIYwO
ErFi3G0p5f3xUglYdSFApIjWscY/TOILO5llCJjad/uarJR2lK4dU//XGTitPSQf
R/l0gAkYtTf/2ybKtLMrkWAMvnV9Cm9Q4BgEjtI4ScPWNitPWHeBA4amQbaplq3f
j3xkjHU/6N/+YWHaU4Gz0vfolMAKrRJ6t5FCKn/W+NX+sWMcit015AK3angrVOai
JnpUIJIKVW7XSr6n/JlTmc+C7XQ+1B4d6H7FoCBpCB2Yf7yg/BmFTmRxaGwjjKRT
jYGrIxfsv4ZuiXwEJNEAfyrm6L3LTupzDm2PC2cCrxHdNIfOsZkjTVPejZlIQzrQ
gh/lavRwFz1qCIfsUh6ltUNLJhkoxUMZt09rYWIMLMLGG4ITp1QogPw9OBN6ak56
XK78G9VuwmisEVbQNORDV45SA7VZnrXWoHM8lXQKKqpfpnyYHocxBVCUk6Qemjru
I9zn4Z3Lnsls8j1yIV3+EYCE1fE/WIJqtMUX9qsld5Bu/R0oq9ooPf4V8dKkUwja
3RLlbgXrVqrvOBU0b99wZGN+q8spz+W5XDjqD0rvcg3D33yloFpEj6grv5YqeQcF
BKQ80ML8g5WPO6TLYRrJkLKsGAfnbgLuwOM4sGSCjljvgV1RMuefGBxLcwily1eU
1rv8ZtifVmzejuq6bZcMGlZJJl4tmZT+ujxSxWHg8o1JFCS59TdUsm8+qBo6kgMG
nsrgBQKqRis3DU0ywOu79CfBt1ZWi5zx+aBZmVUA98ufGXQlftBRo+DZdqDUhl1k
umC1r0cjdvaN9v525pdmDNjHpaOqC8KZun0OHdYYKEoa2kYhYQAotW+LAjZtxNXu
ucthXsLLyInr/bXcohKNkMBH4cFXwB3VliljkPXxtedQBwj+LJd9uW5xkmfYmhvN
iEVcj61b04yjHZYFz6Kb+CfpKoxQX5FAyr44unHNjXeoOAjMSCcCsxSHGSNePCY0
rFljsOk6da/TNOaBMLJeOnx6VXBtird91ZPJD02Cn1B7EuEyl/Rq8HVGR9m6S4Qb
nfnT4lEDx+QNegluP/OR80kyLNhUEgLw8Rifgug9y16NEOmUE31Id/FxwmarxLKl
2a5gzafzTK8J2/hG9yLg2klgK5nTWCQYV+QBVec0bDZmhyCHg2D0V8XjVT8rJaV6
NayaDxX61Usko4m8FPt84fy47r0FVe7RoTJjGLNMITWoJGUtXgcpIGA7824oJVuL
WlskGZZD2zF9Q7FMo3r35EmeRD6o2FMVa/Pi/bDM+2/QegHBwDPHWDFZunzKi+WZ
4jt+hnk+v+APntGubKpRZvOamVCDTmCFOwHfl3ylpEb4ZCwVoE88BDERcKoEMazO
UEG7wbaBr88twXLMAWxAgdvZLevepL8fE/tZRcBDIOsP5Ir+O590vC+8QpKgZXtV
pnsmomqjkWSGewETdYOQtjWAHmnNZKHoW0KGTcPPJgc5o3/Uw9Lw+U1+tZLsRy+m
JIhESBtVuqUM6+Lkas7OXLJWOqoReNOiA3u1tVC06mOeN45WVO/qA3Um98aQ594I
uyyLyQ1kfZE/Nswfwdp943CQhKaPXuSa4kmGp2Ui1R1u6FvcDAMe/G0+USAYO8wE
lJtE9wqiinRTUQLRUiA337DKuMZFm4Zpx+bSnFaudOg0mU8xRtNuJvNjiX1psKx1
RYkaaIOOf6GUAsI6DP4h1TEoqg6MZaAwbNtCROEtw2DQXUDk9x19vO8iAvpeshAl
DuSYqMFOmbLWCI+AFvlxksvHKWw18xMg79Oyv3sNjkwJX24UldiP0bn7Bdm+EU+9
uothr2ooscfIDQQWv20crUmqz1iFYQyY1bSLSfCGG8HElCA8GgP+UnxxHpQ1CIMP
IA0Cq0muPDGmFI1ItEXezbLuA46G61J2Jao/2zH02S6RLP/xExePGTM7b4RwTcUG
o+eHBSnD1BORH+S91N2DUQiMPcd6tLLnglkZ+P59SSsMD+ZV4MpcNojvg4hTvDTD
CgUHAdzNCRso4/YlRKV0xPD9O5uFCtETdJf2AydswQGbU5JuPC85AH9H7TBqAqO/
sW2BUXb5+17zToNq/nWU+P/ffic7snJMPsk2nGZfyGNRPBSkGdCbzza9oDG9w/J2
nTGOj8ezL4eD9Z84rjv71djJxG7PCRJFn9x7kYd4B3Fjh7OjGgtvr+p5DZr1EI66
OQx6/aA1kAFwmr0BaQGlWYZJU+4ghLTedxfLqDgCHn3eC6tpCRjfDuxWwEyxFhjX
mMzBCmCsHbiT/2hR2/CO+aEkkNSXozgLtF4nkm4reDCbsx85MByBElv0P3aMm6Fj
KQ26rA+SIIxDzNZidEUCK6QvcmosG84NT1FMB3CQgRkHdpKY9ztHrH6VPeL7BTu6
+MMMmMTtzRtx5vqLvkEz0UVVv0KLyeth2ggFrDFxDjCVAHedo/x/uNIVcVmsPu2N
2FqXBheXl8V0EeQv7UTk+CgHRdaciAHf2gEx19q9nZo4EU22pSeQAgU0OS1vynXv
KrEQpY11HYUBjiKR60GRt2MI0BCN+f+GQj9tulz6TPtBDuVL7+b+dbtsaPGQudqa
U8JhUvH6+bJJfN2o0+whMhY0ZsR9CpSwxXmnj128dw/AjC3XDnw/MQGQOWpp8dTz
FaJ3x8oWacs/2++IH0cuNyxYIAgMSmlWnHbLvaJ4h3/k3rkl50wJklnE82l6MpzI
MN+oHq3+841FIpVj6XTk5nC7RTBK5VGB42AoM4LXkNfP3aH9uN6p4oZ5G/iLnmW9
iqTGqGzyWpVkxrpwyehpbhO2eqf5QTLxhM8sx/YEBW8RiU+sak8mvLgKb2+Qf2Lj
Tuuu+FgS+QgtEWvWBg2rmKTTPQPxXLX/US9PDtHxhbOk0+57bGsiA9U0PWHNlAoT
30OdB3Kqaos/VCvK5YuJg6pKgu0s4cvew1rkwXH8hXXKSVVV6kAn6CFzAE6nC4yH
t1PfX8J8Adu398R+pPN++795Ef5yq6LthPbFzrEdBZ9puyYDomr5c0Z+gTnzQ/8k
FFnvYD/hdLdTHxoQ9g5XYfEGqYW59qHWMWFj1WMlossYwyn8peps6xKvj/am55b8
HTqupSZFyaKRlI6VYInYB2wg/hnORHyIQ98hnf8Xh7jjITpPAoLTeQMaZx99CSrK
cM4Bi47ryaRXXWI26wmRGaOYFDwedDLO1yU4cJY3mIaHJsiqRT4xUTLVVndepqIS
qhQZjloNznHW0ILoQcS9D4GIgHMeE3rYcRFhrKtOvNBLBZsvh0D7qzfk8YTygvc0
nET2Geomh/jp2IgqE67KSsdr1+5su5uewRxlroj7damdxlr3WR4b0S6haEMv/waB
uMmY9OgyyNJLLh7CSy4i5cRZrzLuJyniuffCsbHQRMhsx3jvJtuY3/VSgvr5veUO
Ed+uxlfgeKwFb1qZjh8rcVnES+p/13u4nhKm9NdmleF171jzrDMaalVOrTXTrEXh
02dXLex9p3d/HHPOuU10pG/E/ayvSwGgkCTx5Bq0yBDE6P1P39Nm7f1QBR8Xzbd4
3TKUsrLtRoFctBFNCUSQr7sc8+LA6hXd3CTXnE5uiXs4y9f04wV/YzMJaiyNQvxK
InjwnYnr+bXKmgCaTcnxh2RRzzcmBG92CgVlrWifQ+qlC+Dy2iLxOzk/KrHo9R5j
ID8bWU5EDahdzkHzwM4SO0u7D6vwEunbK10PEQvgWAjLx5PiRnK0sAYrTIMS466j
MCLL1R+DiIS5k98y1DXiv3b+h4SdE55wGPtRe2S3Gh1dU2LX9V0oFOGT+nfiI84L
t+8B/aNejw2MrgjlqINzpJNH/HcrpO7VQfHIGWAgh8gFtqAnM4PeBFquFeDPt+6m
kuBuRPhW9+Wt1qEpiH0yuq32HfFHk+91whkMjevtl7gC0BgDGWJsR9+SDzyWF3EE
yEx9u5F2ZYEkLXQg00fhJWwabdP7hpeI/WYMbnw+/Au4P53SL2nWS+LJWmIjML2I
m7F2rpN4K0KYdXFjPdaAkwIl1OBFl80p6BC1yyT4TWKFavgF3/8x3u66UVSwE+Yk
L8vhL4D5Pf5i8PhL6t8NIn/oi9NqlKJ/V7CtIeqPzxszKWCD98i1FEB8pnWK3luv
5YEyQ9II3EfyJW7abFfSdeZXZwJ9Lya1R5vEO9NxW5Teypc35nCuyhOrny5LkVUW
x4+QZzNV5j81SyoKxWeCqYHIjD8pgKT02S/+Ti3jlb85Tbbt80D7jAK2mwcQRPo3
FCoS6f5XqwEFcuTpj+Sii55N9u4Zm0r8TOIVDaNJfxFd9aOu7Xvo3x/mRrkctR9F
GkT52q7ufsFsFxuUWO5iW6kY3WC04RqiZXOoF/i6buBXsJeEncl+H8Zmh796FoZK
U404IUSYcji0yHo4BIQ+dgr33efAixMflbLlYbfYYrwXa8fcIKxZrN5ZIXNdTjXa
0O9+AwgNY5mNwF0b1sQlxY61qd3LeGTUbktc03q08qs2chR20CNldwV0OeMcw4Or
8cZuyHTfV+Xnq18qhlcSwI98Yc2RTWjp7/1HWHvrD5Q1khKStB0sOHHpXo72cMP6
xxcEj72PDKf8jFyVZjENktXpk0q/sZyVYsZ02y6VyNwlHwTDuCNmsmuAvb5yW3Zg
MvGjFZkw4tP2z95W5jQAJeECXxXzoPWxVrZb1psjMAM=
`protect END_PROTECTED
