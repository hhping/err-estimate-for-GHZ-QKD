`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1eofFE0/YzlRHaWGjlIvtpLI7ZJjRTOLeKfs3ciPKShBV7TY0k1vz1LPiP6aaYOq
9IuW5O6JZ+QUAo05Hxou7nFH6/NF79bHOsQ3wcLfITw/KxhEx4NHvOaEEWPZHtUG
RePI0KLGsXwuCjo8x4w3SM0aZYaSspozXEyH93FmXkSUa9QMF3OQRtofVZ9fFxAf
jWDJa69NjmFMhzaMKn0PVf/wvZNhbkleCoNAfkrwNf3ZUP6rl7n1OemOdR9pe5FL
FX45au7jEr1HvzdDqL6ZZaI535QG7/PrJZI7UHinVPG4SlGgvg6PQypiZ258ikEZ
cH/hkIqgiA4GbYNG5sekc9Ixs0mX6MT7SdOeEwjEQLJSlS1Nz/Gts7vKU5VbWpRm
7FPfet6SGcIpfj+ap2osYw9zUdOfQu/CkMXVxK5wqcyz+mzE+jYqJesolLEh1+5Z
IYkp5bS7z5pxn6hFOXKfRU1sidAZFRQAgUY2ieL28yDSPAOXELz1/pj2SIlHI9G4
6iWx/Mm1tRYm/EP8Tn2KVmIeLidecsvuZku5yMobwajzxgzY4OXomcNot1+bwH5s
QOBXWTIwyNGypkNlno+xdis3pQlYUplg+Lpy42Kopm7UbYhVmDFjkpxe9GCxI9t7
rIjaJ6L4rLBIImp+pc/twD21NmktQ1qW8vHTTDmON+9qMACNvUSX/Sw1F5Wh0Hlz
fIAb4Xf0KQYeDaXmjoSLfIK0O9D4RT5HwAJ6KlsKX6/T0z/jRY+BqmpJ8XRkPDhx
UeQtczsTgU9KOxOb64Jy2LDlJexNxbzc4FD9JoY6J3LoOY9Q6qu80xNCk1r8Dc+f
L6bXUxrvkc8BtKMRkT1kffqjizm2SsOloYnsBL794MY+QXlTozo+49fu4cQdMnrC
BmtqCj/1yqrR5Dj6tl6rYW6xXsSS06K3HC0aVTkO/QXUQmEJ6Lyf1lx8al0E5UF/
nMV6LfI51hj5uRyA4yq9wVezJoX0eVjnHp4ue//BeWXLOVihzxf7xWiNJzoIOJk1
6KC7SZKes9XKJkZEx81UNQHLMdi8fAMTB0dzDEskriXtUusTPI6YW+gEY5gzZMer
nm1Yp30usdPYEYhHLuIs0e11dD/xQpbTB17ca5apOiXd/3vKURXskt5IfhZgbWXN
WMqkBlLT1jVt2dgq9e4wsRMUF/XmTj6tJ8bj9uDgLOE7N7zYbucci+C6zwVa/4jx
+d95boViNo2telVzlhYvJy4JHDVZzoXAmTfnSlsEUW2p2oq2x3eHgzMYFR+IK9z2
AbhtyaZ6fIiP72mQFQHx83vkPOsn8pa5KfQhLGoxllpO61mG3yI4l4TH4G9oCihB
uDs+wALBXnzs+AxQk0rfSyD8Fv3LjK1ZTRSA6kB3xav8xnvTaH3yqcl/gZmDxc2G
yZBlD2pW/ngd+KRnRs5Bl8Rt2DB/wvRdsZ8Z590NYvLFZ5UMg2AAWvoUZ/Cu1FcI
gYB902B7ZIyaZvdzaeAjmEupz+D3i0RgOsZ6WflDXfKrjy8fterSOQ/rmPdfzzsS
HLYTRaH/olC9Uz4iMvdRB1uTcoN4XPaZECyt/O3lVO0D8N0EqD+/EEo7kUKYxHi5
UpT8Rh9mXkdjRWFAZx1XnnR1gXapsjkke4Wq/iIfkOH2SwWazDRC9vXDlg2JTfCp
lab34IkU1vpbGsnVbO410ciz7jOa3C4hEjwGbin1IIAum/eQ0lnsQcvnyksgDqUA
sbyrdmOKF6PJyDyWktg2+slz9tYoaAQVwgdXP/2Oclu3p9XbbVQ0rr5UoSQXSP2X
q0tNhVFjAcUdVaY8O5kRTGf43h9i7uyzQJuCTfw3Sszlw6q6qkAdM5f8ISiR+Q/Q
uuKqrtSlcu1dIcGZoxGR2eiH5+81lY+0riWPevplmxHHjlA/m0eysaO2+AIIfXTp
CKCzkt35vG8ydkE8SjBz903GQRX/6VS2GEF/2ypixMq+jbY/tFgz9SYlcms7J90z
w+AhNikMQDGj2nvbxzUrcvce/juMyP5Kqro67v2Qr0vYw52PzImAiCdBdi9OIRTd
wlskd8eCBhoVqH/7i2cWtdbZ1DDCsSS+wvJngaTZUDw0raplAXW+iUCsxIiU4sL2
`protect END_PROTECTED
