`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjhWAT9i9WlnsLlUbQuonz7SbgUUSn1ljXfwJkTYB3S4F5h7vJCgZPzlkRBS/G+I
Gx4x1PV1mG8OAPrHnwiBSfRcr1Cd9JQSXOZMvMr+rJx2/cPhDR0K2cq6W3uazJYa
YnBiMqwevc4CrsWVf36V11esFQmL0/S01Aff5vxhnI7/kqawPj0C5dOEHPXCunD0
cPNSfkH1XPIUNx3FZKYsnKOhRn80wYfG4BqQL1cwZTLLoAOyk3ZE+YbRp1c/i8ma
HEuwPmFisLAZJ+J5PNS38wsQ4Z00/iMn05J2MABA+QQlhe01gLTEV+ryNlFxixud
q6IikI/10kKq9U0d9f9OHUZpJunAW/4fLc0+Qhn41YteYUvREquspC9niNY9cSrn
RSREeY3DZprIWq9Y5eMNET6GoGiBdiT8IN7pAyaPtXn9gRRggtejWtnwE7RXE1qF
92Rbw4FMp27Qdi/G6BH1/Td+cwlZ3ZTQaz7nUzFV7jVYTmo3G6B6ijYak4sj8y5W
0WM/jyJ6XyQCyDGhkvocZzbg0TqfAXLPyZLgxeVhra80F/4sLDsLQHJ3Y7TWASCk
tSvS59K9jWpBzKW7A+mpEA==
`protect END_PROTECTED
