`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ly+gNZcSNr1QvVJFdPPs8M0DwWlmBB84FMf2y2kL/OzmeK1lFo1Xtc1tCJIM1RC
mtEvvjjjT68Wfd3rnfb+fSsxeklWxMjZytzeGLJw2Seh+ZL4Rhc81htpeZi5ClyY
4vUEYHJC6prKOG8iQ2dCODbxYj937upzSyhcQgKDfyA8JUh9etWqS1rpfVy9ozGA
px6JZDN0lxrhXqEvyrCNIP9zHkzMHT4HsoZzYTBB3gXmwi/5Bht9NXz88b8wof7t
RqVCG5a8TmyR9Tdqve7A+fLCU51htHeNg+w/1qCD43wYNw/L7/8CFI0+kgRS7ToN
m4POaRPuDlzCVUf0rNAZ+HwfLiv7qT2gBjbrWzWldRatDGu8QUdr0KDfA5m/GUau
YNU0Z8wdohoRXnKE4fGVY2ehFYD10kz+6eECUbeu6jW7nPQZUuh6iiPhyj51+FgQ
HJbKyxD+xGyRyI7iPE0BonYaduQA2gguIQ8WpNjEUHIWzX8yd2Af4BuIVaqpegKd
sCvYjotvJ47v6EyM4ox0WREPP2A/3X4Dpnn/giXz9qHNsMq8an5FuPyPPx3prVHj
jlhHtUKdBjaRZ3URAo5Zi3e4HZuJHTfvQn+SKlu+2tL+mh/UXkXW7ZIkX8VbR5EX
aYsl3X7sZN7vMYTT3OnYGsmLGmXqz7n5nSDPd7oCcWMkUF3ZY2HZnFo5YCpngygV
eDTYwR3VsEo4U8I6Hbrac0wFVdjJD6lTcabc+IwtGsSSSEUC52bpFvO7HXmCGen9
o33LG8TCEthdi51TzFtef2RWUwMl8e57+6W3VuO7foWlv1YhV0HvfS08QV45Oo6f
/iV/GcG1Dq81/aXrlV22SXjr+9T9zoE7/MLTD8lGCAS/WWT5qzp9KhPFM/EL9YQm
MFGKWbuupoUqG72NKR2tU1MJUH+bNNFAMoZBtwotytIl0mEQlLI9j6aaA7O3ibZd
d6jcYLbZ2Kc0cMGaPGbu1UAbtoc3QJocZdXwk+7H6fUHZgVOpnnNcsfUflIyPRcl
zE2+bRsyaB2Beso5MaHJlUu92Laiu4bC8JYQPrmt5iPvLw7fB3YxzqQkXkJ5na3d
Y7P5PdXz6xz2ldZ9Srb+hJEX/9YARkaI89o1h6lKyTgCXjfBbSET1GG12f5jpTvw
8gw09nswkmHvasflKUe2l/NwEk34vxT+5Ri9v4MRgCdG9ibji4KpVv1ev9rZTBqx
G/OvLFXw1iJAftDF7fU8e5YbW3tx1lfiXq2Q8NtWE87uaas1p1Va7Y+V9qLL5RV7
9wicvEQu8tlqBV6HC+TsEHhFGMT0WjCjbU4v5yF+19jwuXDPpz2v5DSidZuDMMsS
Y0yRjb+05moD5VB0+XhCvNxWMIEbeORbuWrRIGJJv+NTP3PDyWAjLVp7wMkL+GLQ
mtCFfgU79J/eRD7BeS9Au+eDghDprYeOhflHNF+2zRmw31AJ5GL6bU0EvEHV9wsF
MrkisKk+yRAmZ7AFUQYVej+3GQcbjsMFlU2uOy4HPM5h3OGdw7CWghK1A+a1JYId
0hM4whTChgRh35VU8qQnlCbqferJjzHT46NucSHNslrY231w6/FVfUXoGP4SZDKv
9eJfMESHwzsVXuWuJuqyROKKqEWqZ4Q03P+/x2/JwGHfxJ0szdspkZ/00ixBUYHD
HG46iYBwlBk8Dw5V2YkKvCAB7NuuEpH7P7H9dL4+B46u6FYGuZu8bx2sfWWF5Grn
vr/NQ3A77tw/BkH22zz9FIop9jPaKDI9yuNeoTBayQeSahnZPOCK77X/Lo01N/lD
7mkI2RRaNytFfriwQtTRqOBEqpOt8TcSPA/O1jXaddzovRblu6XnO+MQzRjTb9tL
VIhqAk6URyYARwkFKogzBqFJHoo0SSD0GPwlY2s+fuuwkkI+IaWx7RQJIahDcidh
j7kh4b29E1qRgpE5aPNPIJSJsxqRdI/Va/o5Y92FEBQQa12aePux3Q9Dd5AyFPxI
3yP8Qbs4STzAEp91/arXgdn0/fHJG8KHm/jwPDjmjSCLlLJsDA6uesVifrKZpiJL
Mo+PEzsGM0ZVuj9+r8t3zbjBJY86J7SoBcdr3c+doZK1HUAZxw+7+aORILftAJmF
pwffikUZhRbA+tp7KEhfpuFNkQYhP32CutzBFkXBfx2qiUQII5uIm5i4m47mKXTC
dcnLWd47dgLMVYkkcw1npC7Wck7nuNglYnXun36WYlvUCYXNYWBlVZt2Y62ZiBfg
JUX+A2E3CDRjZ/eId2kef0gmcpBQGHtwOK+t4hJg+u2oQBPlvW5I6J8I8kyKQKAq
8pHNTId8EAlCnu8bSC+1bAnbFLpiZlPIzoe/A5vVrkPmd/Xf7gFll1VRQDMFMDXe
ka76K0vu8iJ7VCHMGO6ko4hIz9sgSjQRijqq7Gn71al5P+A7scJlfKmkROje7cfR
GKazskQYRnmFj3INPBBk+DJY0XfTeY0wbCYwtQQkcFJ7qj865WlAMw/hlp/uIEii
m3QqBd9MRiFV4xMFy6zJaeBLT201U/VwWZKSUxZctB65S1PEwrXgEZgRzSxng9Pf
dgM0oQvhkq0ugoKg7VmxJOLfyoNnFT9hPSGaKd9d0F3odYMn6qrLR69VIz/qvd4N
RQDZlnRjJRNrDuimhUktWue8MgY5zW/3fG/+IJQwbAY6aD8oM4YE+oFlzgMlDt99
SG9jOr2s/yyYSb2IsX+TG9BpdlANtT/bwnid2BKP2r7v62AGexDXa0glyNb5FCHj
lA3fAVgZCfY8LJtwX1yHy7rpPUjMQxavan7MPwdRrOZaEEQjyNXbnspdzcpQhxIL
McgSRj7S+XQFDFDLdD/TxGmbUm9xSOq/U3zeH2ewBOkIEjF4cd3o7He9puhvnCMP
W2hC8otYGB/uprUzmlySW8o38CStHvA8MVB8mPBrnnXMSb+wvc8k3sq/R2P0goo7
Ld6iAJCxY0ATlWPYjEUXl0vjaBH36nc4qpp0qotaBkV4QwCHCL+a9a5K9+tEaIPh
3iKS0nS/Ffd5L6AcQqYYuGVHbAXEvMVQ1j562yLW2ehVsJhEJL+r++Z48Qvq8GR3
iXn6URqCbw2ZXb/fELo+myJWbWbUiHN3mtVv3k2c2zKdCyVSGdr5MIy1uoathk9Y
R9sn6A7nVjubSW293zxhHMdpv7Qt+I64xW5JS3lCP5qN2FEdJUDMv7ivPWxCcGIP
fSrjWQX+sLE1W0IIiJs6VQ==
`protect END_PROTECTED
