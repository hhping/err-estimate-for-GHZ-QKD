`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CPSbUMcnW8RwVXmXFZzrPjlj4QNCUMr4/HonofstJbG6qD1xxYgkoMCZCMNaGKZs
va7ms9ugK+7qbIVcXuc/OxXUvU89rsQAHrEiPeF6aMDbQ/4pRnhe3hoC30/4spgq
BJRcXsYWbocFascXv4NnOKDeRZ91GEP0f2r4Jb4r+3PoL5BUOAXGV06XavdMrkTz
Ovy7ES0OIQnsxx4ZXcgYER7LFchVlQUgJi86U7ZcJUrV9Y51ck9ne/+CIJtn+VAi
kysvjbPrQHlQtnpbiqjWrQf5etOLpfxNKP3D9haZJvHxL0h5mYFi2ustMHaPh31+
wPzmb1Ymbed8ZaJ3hJum2beqZukN7UcBxoP4+IxC5OYHNgAL/dqH9aPjWCaKbvLC
eF1hEOjzo5DxTD6XElRmkstK/JjoDX14V5jx0RSHIMwe3QsldBR/SZ+sApudaIYp
kdwZGgB3e/2/CTLNrmMuh4ulV3IQrjaiHWRM/O4QXCpUfQ8sIEQxjlsrPLDkO7s6
TkYTRNSu1PbOdhWKJszH2s8EOIhETnSAd2xklw6nHz+w52pB5R6h1qGU2UOM6E8m
LNooXpjRl6pYie9RDxik4ksOIMARbMtToCR9PBCCIYc0MVjlGUcJwANBkyP9Lq2B
p6dO8ccuBnaBftqLsBeOyqjwATIYA8rwHc5RPUbP5cZceIyzonbouvm3yUP/p89S
LDQEWcHiDw7dzO2Yqp84cC6qvYTuDH4zke9w6exT+huPjtBv3Wwg9gIJvphmaTpe
Be1Zq5jZkO2GVsTJ5rpumiD//IqWFxO8Go0YwVkAQyj3kFNRpH2oQ4p40plEETt5
ter+QGvRR8hyEZ2ClOwn01B89udhJSqBN318HnLQDs6l7djrqfq/MUjzA9dN7DXc
JO83W31rvu0TaH3W5BTJIb4QjtJZpjYP27lWbnIz/KAWKhZnkX4D+j1ERYpd1ZdI
IKf7NQ4LRZBW62e6YiULsVlUpOPP8WUZmD0zsdKmhVHN/3edOfzHQZaFxm0y/Gkg
fM/W28OibeMFlxuub2J6S6YhtU2ZKADuSGMGg/+lL958/wWHDVwBWKBplgODZ4/i
acymjR8E7+bCk7jU867a8mEyAPxCuTVjcqjppZjFZFPQO8Sb7z+cFh/nDgYJFyIs
vIKPKO/Z0Kgt0Ee1pLLihYp/fVyvk3ptbJpPe6lh0oJGbdcG9719bTtNH1+jZztA
edOm3gT55e9M8lrXFLm4nG3BzDuzbvYaGwfcWzL9DcdXhCLVDNWLg1VasHQL/XyW
QyAmnFsQV/55XLLRCOn93MqTa4N29Sm7XWaUwufjzABKvh21p+wZH/r+lficBitU
qQRORn0f4BfRva1qn6TmMfQ3yFaM1n21MY9rE/oekdZkUeREZLFfaxpRYGQPs/Ii
7Llhvs4Q3EZBY11E6MvHR5L8yFUDu5fvJVmFFFKeMqMwP1Oygv7OpeE77oYivE4h
XEJOmHiiEIQHA1zEQ0Id6AYBML7Z2cc85RLXzXHAbzSg0B+LnJBAxnhV2yY3FwMG
Gh0WwfTbiO8yqIHBHC6TsvzN6mc5VYxJVkXNj786nPusIMFWy5/poqULq9HN6Bq0
KYaY0Uq8VnVZ9i3oO8ODi4VX7px8CHWhYG2nV0Uq5ypvapOyuOJzZMC8Qn1XO4rO
e7nIsl2QJisTecbANx4TQWoBDFWTOdea0mJ/PZOc3h1AiA/QspCgVhR9NLihLLJX
+NRX/g3YukFXpj7a5oW3HytFQR3rJQGh7g297htsXXPTuV7m2pNCWI7YeJo3ws/F
uGIFI8k4SBYbzXbP+rYuPjOPeJxl2EJvzp2QwXfrklAnlCg58NaWYZMxM9wNPzr7
iN+6s2k4RjXI7/GGra4XkpOiG8KmNcyWEHulAvaeNzpZTcRFvEjR5NtAirGo9zOq
+OkHVYZlXkMPViT7rSepZPg7q6+VotXReJrfrVwbZ2MGYs/XJ5MZpUvFhEnWfKdB
QKaN0gb8jqqmbUc4fRtbFqTn6olZFNky1ckm9jY7AfcIRP5BMHUH5rZvDTHyvgGT
/NqIdM66WaC4F2yqzNzdpK5+tWvWQsklES+hnVqhTNAKpmkueKR7eOx9qi51GFgG
cSqjdqB76ODH86k8GbfT6HR/CThAuoC68u6b7vRmC72mR1YLLKyupQytLnIa5N9O
x7/ZftkY3b989L27NPu5cXbaVH2QmT0Rb0ZQuVlqX1RWE5UKjnCF38z7G0NjNzBT
CQtukB22UrMiaok5JA/Y4lhwTw1cg1Qm7gDKWQdYfqXa5mUFyb9QLq49xYt5ici2
80OE9FNCxlC4z/SgwYYQZuMuqdXBivdKuM1heLsmL+Jl2Ya+t2yKDT4iON10tKBY
eB2bhMZaUQM1w/8FvuEHh2gY8zMeo4LPeuBmK8JhPKd+ycTVce5XhIqNVq4K8fM+
hZuLzv8fu5wEsT2yitjwSLiDMXEY1g3sUmiuVX7WC+oSNGOT6MEAjOUgi6Za1kgx
TiiIkshrAk5Zxf7pqGS78rZXDO0irZH9QbWd8pkAjRIe2HsrokVBKfE1CVFI0TWD
aVEPEyxtiefZ0GVjmSsNBKbxd05m/GqT18EgVzAacttv3JRkWLt81KI6IA1MyPrz
u11CLr9x4wI9GjMzJUINegARtjXjmJQOw4oNx2WGlqu1fakeYlD9xlrewuEAe3m5
G6MYybxDtJ3XiBg4gmDlZIKXN2DPRWpg8/ag7ab2H6HLUzdbRk7+NAHqVOv2+Fi/
UG4pKVQs1GlJnmvShedyrEAr6w8x9q+s4vKWavY/bb4knUx/PAwaB8L987KkIb1z
dj5u8lgT+PEt/dxTpf63Awu2gCx6eO/ef0kosHA5xrKGjY0h4ptaJos91veQN41x
8BwBnamxgmEG85EkbV1xziwuGFaU6+UuFvi7XtetyibPj04CHbJ4ckf73TYJ+cXo
f++wVSJbXOnTYfRH9WcCAeL3MnSNkvbYTg7wbnczjSEvIJhoW3BWZr72+ITOi811
oq3ZHxgjb3jCFf/l1fHdmPkGYBaTEV2rxa/Iq70BwwzDFJyaBgtt0ClSkP18pBMn
/8MOGY2NWHHT6Q7rn20b+1zsgvcPHz3h4XahTnMyTctYNF02nxA2nCBOo75G+gn0
VTliTlDuORI/ZxbPu8vGXWlaOl3F1SjG2XYUU1oYEwN1kI/2VjkHCdZAKK7VdrWT
fNc3VKhh4zIh0h7w2Yun8h/w/D4aeyp5bURZX99v41pcZEWqwUd/KO9ZcxOnZ3vn
O4tdO6BvmeG11zLaSj3SvA8SDjTRiq+vXihLtUTJqrUTlJn104uhTJtET1ymkP+W
XMrJM1e1E26FGwPpSpHasqf3oxyR5EWKaYCNY3aNBANOJAul4zLeEaLpJl+GSeLu
4vQxhi0M2csN6IUDD5P/bxsjcZMS2WgHAFIW2wDTwGsgg2njhkEGzr67Li4AHCOj
a/0VEVB4ntK3gaj0D/w/FXmmRtHDND9SC6TzWDfo1S9O8LFeaA7/A/raX6ayIke/
R5UEXc/k/GezOvzgfJQCjyFu6wjwNcQOZa+NjjNH53AYEIOOoeNRspWquwkC20oX
RQq+kk1FhmWbs6Fx/v0kGvxgElKtgXFH31AEyUgK/Cpjc9pd1p85lD+RiT2wKIx1
6wzfqkTJ4EREzUpAOryI/66G2b7yyP8KZUAcIjw+tIJk6OEX/C7cDN8SrQ52QfgX
53cNgdF4LRKIqOKCxZ3T4ZEyEDXEHGsCEaRsUM08EeDn3GBMZYlLPRJ+0aSemCdm
dsIHoEVtszmWUbOvX62hA2qYaOyijoT1x7U9NWF+wifynqpcHOIk/Wpc1by7dSkQ
yaNLXq1Y29ZgLQNt6eymACK9II8CGEmkG5D0gDnkrn4yqb8qZztjtYuFCbxtuMb/
udkuNnwhsqkuk7dstjM/QT/5YttslFzABKO4LR9Y6/Q0QBD2HXFcTPIBP2LpYPVg
nDP4Yi+AWqhu1kqSU7FV0TYrhNa8ZgTjpR1eDyQJ8SpwEOAwKgdVh+HUMrTruKkj
nWf69ZVZ9uFwCLRs4WQlLf5UjY8j7lQyO646OjepP2531vyoUDsMPViMXNrLTfM9
ZRyfQQxFdYykex7MoEnxZdimqvU/HVuO164WLMpJ5Y7kAOijRJ+30O5+aueZq2uZ
He9xq+946tSDeHknQk4RgbEBeQVAZntewKfaGgIbmdKLuF7lYyzGlgYc/z3lHNDd
yTKrJEOxFjr+rmaM4l8hYmirn/CLPu5LoTW/0Dmj8UabxoFCF4NOVepxm8Hi5Ohz
a+BQjk90zDmNkwPIGYvyx6TXv87gJpMx6ceIs4/SxnXmjzOPR9rNKJKzfgcJla0S
oF8EPXQlfX2RBbpt938mG1QVw/U6TQUPZ4XZiNxFjiv5nGcc2YofKapr8HK0bLi1
bahYBlX13HLZmz4ANft5Av0H7UEhAQeJpeC27YADE8CJIIh8bboJeUttdHJ7WrD6
dEICYGvpu5nCoFUVJWk5HGhesK8sUotjXMnHk1rg9FyLJ5bo0+kGjIpg4LYkEYKX
xt3eHgorv49KQnXNIsfZ9GAouqX5OvUBwWE+5JO97+kIUsE0v3c6UVbEdUns+K1H
US7oHmw2FK8v1D3MkXWKN4tiA4JOrAyzeQ6aKtvljOTi6enTnzOrXXsfDdLFIfd0
fO741zdRFU9xQypKHKoa23fy1XuAPFaf6OLezs7VJ3ZYBr9TxHGOATiionyrQxTT
D/8A1/iLCMi7JAgYPgGUoIbsvBSfRyi6d4MzJXLsAiRa5/TAfVSsm0guRXBNJJ/N
wZWvkcsV11PB/RK53jNDav0z++smLr3NykAge+EafaTRRXoyXxqlaH4xzp/marmQ
YBwMEwedimRA50RlK8D1edKkKSmvnXpYs5KOuaDKAWFfy1WscxPo83KaP7Gv7+XR
bRlVjXctPwF8n/mQ8ZdAAxM6djKbTdOegHTl4aY6WRddzIyJi5E/SP7t1QfJtuZk
bYJuQm6N4yhYW2XVDSpj0pRjdhwqhKbuBtK0CBG/5/RpXnP6bBTKR9VU99Cndeu6
YZHEs2OF5Bv8LrFrnZV/p1+yz8U2jXxLUzikYX4L4DDttOX8Eymv/jP+SOAfI7VL
TDeE1uUGj5kvZ9NU4Qe0FKU0k7hIftBdzuGg8BezwVWeE8WBZ6ZEAcERKvJBjD5j
rxdFmJIUvPwsWgbeRF8W/fkgAtkfO8f9YdIr0t12rsqz1aHFaD2dEsg6cpynjNH3
dZ3lZ1f9+isZD8orPe41prguFA5Nc89KvizM8pBgVGGHVrWjVZkmwnUfOQh3Ddlf
tAWSkwgtheqCUri2WfBk6ftrOSy2FTiY+Ch7Z0Vs+OMzxKV6XMgkW2l/1ppDHPen
o1JPhXnQR6P9MqeoRlLZQPyb9r5fkaYg6b4ZP2p8rdg0E4tp/CD0VPFAT0LZYRaG
w8Fc1dx0cRi4qP9bgo8ACPxmQk2AHBENWVZvQUI/vWdeBj1OuD3ku7uRltMkqQGl
1uBhICZMvuQK50czUKAUXYyFciM2R2sbuzJ8G6cWa8KpQ7gT48NmXlJlhajhmODW
q9oXRLur6en+R/IQAY/N0EKxFv0tRv7vWSeofUONDwvOxmGnntg0169eld9X1/2i
joI2Q4ZRhnOY+ZNlYYbqZSnWn93zJnIWHUWDBSoEed/ysb7Q1RwvVRLFvY7+4/Ew
lstGB09EIWzONih2QTmWgn4H8IxO2jAlu1ljyticteM73AyJY+trFtNNP33HluFe
aHn5n/2JKe8ISRMFFQkSirAFuxGyiKqNRgHuhyGImZkEHim+gGjxbUTlwmG1OgRk
08NJiRocyvY+ha7iLMe8iJRPDyplhHeRowSPTd1NDHD8j/IH4OhAQahOUkumL7PV
/YPR4G9scl2QRM4JgW0Nr4nOGeP9XCoe3IRf4HdGNswUsmNg3WUgZ+7hXNdb7CkP
wNr2EVf7Pl4mfGDPrqWQw1oUlBIBAdS2++JtAkzuJqvnzEHP1fveVVn1HRE87FkG
TmNDvIbVRH/HO4KRYV+C1m8nzWH/NcsgiZXRpSrDSkyfzKsoru/JYl0gfkptY/rM
k/d9yyEathi8v4oWJxP4QXcNBLgqLUEoeqIqBs9xgJhkDjowHwnI+/N6tInFT28G
265s7kt2WCtSH1rQASfyiiuW3s8T0VS9lPD/ea+fgrqpcR9lG58HbE9Cycj9WZ3q
elVduOalePIlich6OoCZeAK7Y4P/jaWq6BH3zgU4BZQWSCxneOVoFjct7ds81Boe
/Ykr5aUKGAVvJcL8OXII/zKyxDpnyTZtUhRCQHUHqyxyam6/CezbUfBODPhaT4lK
So6/klv8RfQPIcTDVrbgX7366PbB7txmxykH4Ubww4zXnEgfLC/hmBm+fh9zrHzf
mUh5Z2un6Aj62yQcG2mRlrh+2H8VgbiJL2qXjoe9VOlgxSeJ8b+5bwA28zRe2FD+
T8ohSHsYrd/zgVi0hSK4pHcn8mt8uAm0esNZ8z6QO/TzV83R5nKEb0xHT4yQdMpk
5NAsUx67/U8kIO3gDDzwsf8Fo4B7KMK9ReId4/v9sk8k3jdNml2q5Fz4CkpbpE+T
6hKDWPZUUpHBJdlI0sFhj5Jx68norSlPSZYMWWXtsgzSxmh12AmSuG4r2kA9naFG
+UQWSVaJtWvUC+7XUbjFramebcxrV1oIhixkwzSuAu4ILVvmi6axrn2fjnZ8xiS4
REJr6JAtRn+of3qumebPM6QT9ahHVmXCvorNJXun8kKtEmK5Yaa/LqVzqbUPsKwX
S1jOv5s9m0dRxoybUd+9Shn+vI0X4BRJidFPo96r/7dSqKIsHD3iHVpIEk91zg02
LsFRPwxfnUNz1WLyEP9Z5ql0LArmnQFjK88nqPoz497hXg+bklBUCGtTYPMC6lnx
YFfEzJOTLLmHBx7ckifr6Nc4lBUbW7FrXm0SJmOAYr9mBbcuwau12lRa8JhkIfwV
n/oVnEBJVF+rbnn4tlh9QCqveG7IGrrqzTDIOBQf/uEm1yuEnfTej3tYnDxYcef1
c96p92hE2MDvTh0wGIRlPd9nZ74jDQZKqssfAdoYdfaCFjzxDe/bT+6FrhUvUQ4n
pBzwqa06cWI0TIvi8ZXAsgcCZd+sgYwIsnwaHWCDpwfmhRhionQ6smcbxz/WTrJb
FJFx4fmGBg2wHWl6it6K60Sk3JXuUXKUfWYH1zPlYKeG6J8NbHnlTzv4pmd24rv1
BYkg4SxZR4rMJhhP7+1QWwe0d9y8Lxtu/Yxjvuml7LrYkzeTZonxpOUczXNfW35i
+szwgnLtXvLl243aH7d/MjMpqNB5kYlLmD/0QycHCU8h6Jo9PDNSvYt/8wZxFs79
FfYiMqFIIL1aGzRTJXQOosTT4nYQubvv/ium9qW3ciytlIAXaaBhsAXIEdVKDLXO
OuvaEx9Nu3qNw3EGnNIIbuvYPzj3flEtxiprr83lysXOmdfz6d1I5s65eo1LdShJ
jEZVU8uDi3d929QyKAl4WMWKSLUpOfxN9yV/HnizuQrbuh5wpHiuULorrH4tOBzB
PILWmebm3WkIi7/NsByjzmEZFhjwIt+Mc4Ix3QSZiOv6LPZHhGPCZSu2SVXeb+mX
yvvFdciLUWk/pS1fRSu5yWwjL/bAte2pVz40r404DelMajfpCkVM4aAv1HBWCEPs
mjsquFnOLr/ftB+cTYG9hsgcD28cR5OFNK2lby8oLOdhu0zsL86o8+sA8knFPQD9
7MkqzgWrTlozWyA9eufhzd3ZTuvAK8XTpNy0zCuuKqHqc6GwYZVkrPbm8dKKQL/C
ZmUPiGIb9vQRpVCCOFZO9COUIDe2kGwzbYSaBqsA6VtZlu8n7Akqp6XcfliocIdh
EKiXswi7qyPw9U1mftryhxkr5mZdYo5zUjo/bX5Mh3m9HdLkvFXq826OI48AoGJF
wuF3gvYeyrewnGHLKQxA9c4Ey6VP5mV49dZc0ylS6Wf6M5HjzcrESJuT7NLCh8Uy
yMKqeyMtSFhuV1wdjT86m07HiEVFCJ/ZalqlVqxHPmOmUVP0a4ddtKhYIkFKU8y1
Wsmd7LV35F2GBncgPxxClZ4JWjITOrK4V3OEuL3H5f21SvHxLjHRq7tx1nYnW4qj
cacxBB2LcFo2tzmi51/YjWrP1xcy3pUPjIWMZFWGk03vD+f3e1BUI81g85q3Ah3V
RZH2QZXMQHArK3vHG6KagZfLGGb+XoL0P0kI1/81GFrbcoq0uO2y4eGKsOtpHiK7
dm4d0Pd5MGJvAOe5jdb+pK3vd/rgC1YH0TQcKP/tVbV/hOsPcCoKpcIRrc0S1b07
DYPUCTKDlvGnQhdxYWkbqnmQ+fwT2wzvv64WXGQ3ymS/tRWGGXIp2ExLaO33EUcT
EV+gwqkbQhhHuOisoC4oa/wfPRCmY/ZvJEWo/Us2Ia9nooMOUt5GWZ/Q1hMGGKSi
VKCMLZHiY+d26+GqM+TxnoPwKx/u0MpewK0kRy2mNtiYS+9lTcekWpc1Ew1rjkhi
8fV47Q6evXm8moOrOuBS1YHyTuG27Fpt5wUH9N4R6Coz2Giud3UqH1Rmq7n1McfK
10EeXMUjgFoqJ4c2cQBgCnXrj/khhvIYxBBgFDSs8IiSS5CfK1oZPqlfCd/FVT+l
qi90nFaZczUfAeo5zyOdtTvzTCT/j1tQcTqcyH44l+F1bYXsJLNuybSWVZUivpy8
4onr6KboMwV1b3P33lBTc0SuYPd117EL1D32gAzHp9qKXLYFGji1UfB+14TWs1vm
r3lxBjReBolVTSdZxk6Xs2ZudTu017JqanZT+dnIONQOkUlkYrhcqelX5gGQowas
JBR/9fY6Z2yh5KiYZDpxDn0+EEVFkTqr219RYAXw0Q4to8TLTLI70U2wwIJ08MaP
Ev86wfSj5VP7XkhDUNoluv3enn3zl0HYT6qra0LQyMrc+VJmT4HKJsjkOFhWKGtE
6hOAneXbqIVeY9HGxyBdfCv5FFlBX5cTG6+5LhnFCMxaj3ObhWOLhGzKOBILA7UK
54Zt5d9A/08zhXBOas8a4ppzWSehPivup/Q5670qrtLvRgovyAIzePdAtyCrpj+4
eq1L9Nm5lKsYB7ScQQ64Ej8kGt1T8HXvX3tVYmgPvAdVHFWN87Vi1aHt7TppV2Tu
IQ0AlpPc99YNqb4335YlMlduyxhif4iYl+87qsKqnNhX/U6LFdyTVCTDwVZI+dVs
oweLWgvAMdrnU7cIh8zkLt2z94Je2NsM6VTds3eqEaPW1q+Ck8I3oHiSbB7ehzWB
U/MAHd3TydKTk/Nj0JgUokZqXlPr7XX8znYn/GQQojHVDAZzBJLQUYwKI9ZdKcHf
9k2KpYL4CsYvJWO9hkkxvzV1IYdLn3w7FyB+A5APgObPkagThTucVkync7D9m2HK
HRowg/RkyyoV+PBJ/0aB+xOl6hgDd7ctkt07G/k4PGKlxr41KN/GMsrHwRCmiFJA
Pc5A7fwHjekZzKPnvdygHo2PbyJgeuAFxzf9faAd98vrI/Ca+JmQ+8UcGxjvytdc
JLM/ya+98Pi8nNN/eoEhS6XHq5pT/1rIQaU2906zhTuj8Ix0t4OtTe0Ovgl02+s8
u1eJjY9kPifaqF8iV9C9KB194RQjPNAJ9URlg81AZfDDX5I5G4cusXYazTuFM1B1
36WkFwwMWQ00OyhVbswpL2oCZAafa3pjPvO8NzUre/Fnqtzq0DoPXLcdNiAKRpJm
m5hsvULTkLlpBe8AzOQx4Q+bhV4TdBkmC1IBStOcMneIRk5c2lffwFoK+IHocrOl
d2q/s1bM4P1zrU5fTPWqxt8tSaPSk7hKXdDFuc02uToXfpkMNuAs1Ud+OJv3rSCK
IhhoFp1EceI/bPvsD93rUZnz2d14ifuhVRF/ctK6tqOE9rDqQbcPQtWl7v6Gmkt0
Pv2Y6mQTkLGNKxRap/AD5JswxyWk0Ow3OkTo7w1vCFS2BA7fFrEAN4IyvA6/hsJ0
S6icGIWzPEN5tCcftP/IDpaztrR/DiuMYYjJVR36+iDmlvq/204cWcVV9pnsNwfN
l7Jr7ldeNgj9UiFyDjAgAbDAkeqOS2RL5eb0AhoWs6Kqia7flxRp4lX0riDM731r
InFW8K+FOydcbvRglRAwm+ObtrocrxAo8j1SZ/1U5z/TUnKzRPI6J/ldW5qEA5VM
OvK+1/nsrm5Aih6aqWV81Ms14etNnImm1vUdRzOFvGz0VOtkhzPywWCZRsrpX0ek
B432L8+UHhfiQX9fKFYdzNJTCNkhBvSbQOI4lWa7m+t6QW3NWGLpxnePAoXPXasT
sBQITHM/T5zmN6iNTyUDQfonrt36U7XyWA8nKx4bRb7WIaWe71tRhZB0GUcRIpMT
RjyaIdqmxuMj6KeR4NZG3QyE1jEjlukz2qSgf6pw9NOyour6JLsKLAvPcmdTwiXt
hPpClvFyhaKcun+K7RbmFnOVCVitllOq2VdKGEFIvDvFVaDKIj2p57DaOPZEujK9
LBBtLTi+/E1+FcyfWKavtKucAuVp4YctkOwBR6zifxVDfwBg8QoeqFp31dZaikQm
zXkS1qX1lIILaz03pFcZxtsW+s9ExE4YbzP+k0WzmW0507ir/Ufk+JLxJhkV/dB4
Hcl9HRAiNwZp3I/q3sNnROUKXlk8IWmXpPT/bi610mX8PK4eTosvYoxRXoUrRTFW
L8AkOsCetnQTj5pFC6aYzfUPQoaOcKc9m9VnNgph1ajj9rSdcvFFBfmEVZBhiUaT
nXwHaMDVgkZY2+9qGWOFOwz3wW6UiJYuSQkdK/o2Ya4tEcfAYc7pmEe9d8fMICKN
BdY1n0FgMazkRqH+ipZoKYO9LZCEfbsN/KZ3wL7oOP0nNWzxY94kJP3xcFbScmjP
S2ie251XYm4w2rNVBuDU/qIYu86vBe5xMLUeRyOwBTbXhaZHAH2cPa1cEGwKZbRS
AsmzwJ9Mu1sHtu6LAelHOaFTDaIO1DpfPunTKXH8wlFOg6HJTfcA2LLLFYua0qhu
LPSqQJ9DdcwlNq3JPK8oeNtKqZ5GoDv/P5zvSNyN7vot8LlH7twpwwMp4WmkiWu1
JgccgOuVbKkY3Q7VHiz26w9JxUs8B2tZjGArbLWh/nTm463Eh+BI+qvHGXrX1SNX
gIClKgFGeudUsdlykrNNIbmkVkVxFt4m859g1gR6CFSf+V+KPznyltIv5/wKcJH4
gs24ZTL+s3byk2ga3A7camLqyruchCf0Icx86aF5P+SJBQbV3/XGCCYpUZPLMUlx
t9b0q1yhTCHGWR8lFaZjwGPKx/0E0VR6kF8SEE5nqzUgjRbTwJs+Cu3VN4kcG8mc
CDNt90tJ5fRrwPsKZb/l7jXna3//JSFAot1ETWfPck3typrKkqd0Jm9QGxysVzen
9t7Ay4WfYtM4pSOF5N3VYAO/89u4HteJHuuo42uzY0610oT+aw7TrPZ85pwwWjmQ
wD4sw4VoaaqjuG0J2GMnb9Bg4VIE1XU7W96gvY0fw1tnFvGthyB9nj5LZ6ZefkC/
RlbrKJIc/oOpL5p01pEzBTXCX3l6/2aGZihdVOFdSeSYsXydE25L24bs6Oqy04u5
KqTqzyw8zp8XNrc7MYwcPtAklsUVhpzvKdi9L3OX22gwahNNjA1TI60DBiDvEys5
+cC/aK9+oFfpg3FX1hahibq/FSirPZ2b4ixs9qy5rBCauyi7/sxVC5HzFe8JDrij
vx1vfB8qTcO4p03gecidvJ/uE10Q5TBqlt1g7p2swryc1aUhaEGcZQ/Iby2K4TeB
XUb7xTdWL+EAyy1l9F09B4GwxBOoh5xzThgZ4wELKQYdrImFKRT7155z1ApUZTsu
QwIfiurPkZqL33LA3SRgFlX9c653mRYttEN41gGmmkBpt5Ctb3Epvf11S7Op6fwn
RKrx7E/3Uycsa5R56PrvPSnhWRU8HRkgWAtaaxQV/fb+8AdVANI6IBOvGh0fwRbC
C/f97B0sQFB/xOwe1Ap9iyx+VQbQzK+LjiR4SOb4oGVgcd+f1IYkbKTfvEgWDjw2
N1Nt30kYlIc7R9ts5Y/+mJJl8CD1b/F64TrHQLc1pE0BDTpAuJ2z1c7F8Hh7UHGd
EOW448sndCHjoqpUVAKV1rBTdhhyoP9Du+WBMrfg475TqnFaH9mJSmaTWqBH2XAl
Q4QiaNGsjjbC9iSWAoiz7MSluKINbbQ6lhDbo9s4ueW1dkgbObiiUCU4A8WMXgv7
zffOz3pXkgDxFlq7l2LhxcHD9c8viSNC60DZc8p69w0+DsaiGylM0XwF4Y0UhUVD
xQKaZ3qVrPlJC8VJw8+zFyRPM1cD4NrZ8wADySn6VGkSgCF4iCdua/wzQT4zUHGU
EYEdd/QNAu5w6PNqFJjjZnVcm+twGiA3FsgeZtFiflJdWH5JDJbXpBQ6WR5p/yaw
R0RM3Uyw+0bTABPNAvhZVMhEVUL5wG4eZp5n7LiQTXXvG/5BYqL2COoecGyX7oNN
yP6NPTCScOUB4f9DmReMqQeHFleIsWushQddLHt+rweB8ae+HC9xVWMQMOwJcvHb
L3gYqMpL2qt2pp47G2kOMLDxmOHZEyWDeKmqgI42tweetziqVbatpBykTnlsaMqJ
ddNZgSa46C4KTYKLI5k6pX2tpCPs3aYG7/0QvWWDMpewXh6FKCZyZyt8UGz67Uy7
w1yijBiKtgMOP660kGoPKWmvnTj5jmkPmix8nDVG8pCDLQtaHaQuVDpvL5Gelhb2
2eU3yuDU3rpGG+umK3k98dIXv/DRJtk5Lx3wivO8dVY8Qy/eb2WBK5hivg8P0fUq
yeDeHtuDwu5pRWpuXpfO3ZnRFGa1aNIpsll7YY6uMIFhkyVReuUEgZsQV9+ppuH7
+konDlj1Xmbg064DUMKQJZf+fjy5IMLtsAys4hH+8/oHpopyoH8TnHRMQOQRRbqn
BxtLABN1JGzoACabzljCQtSvdnPeLQQYsWzGe/cBJC1xmWZOdg1fWwrpI2kMcPRZ
2EPhA+evlf2znAtSipbg/iKC1dcL83eDoM4L0o0vLhIbrBI97j7vmtAIx4FJCfdG
Xd7mHxAMT/koMdcgdpVyRgrkFBzlQuZ1K7xkvoJhyvFQyfD4lXPNkQubNgGnQ4Jr
525eAUMTLDaESVaMlBdfGoCDL8vHLjldd69SNv4JOZeoa4eXxI1VAPEDjCq28HEy
eBqUDbX+3l7dG4jlpnB+joYYoP9Kbqx3xBQKjPUOKuMyks1GtKrT+AyOM9/3g0gS
8vmP/iReZ0hbKAbsVxUxMH1P0EfoOrHMdM9Toq1lF8wxU65vfdUyJKcRcxrFQkfK
ZNxOvl5H4rVtAvfv/hwQw4dUoaQzfovXs+wAliYrv/4+EfG6nho3vf+b7axHCpFS
u3oewzRxrYtJ+NxRSBo0SC4lS0EpOCkgXo999y4F5Nn0cSmk57BT72gmZ7y2CYtZ
9HhHS16JkMdhkKenOYz0ZCgkDpl6NHwbz2gyPXpQGpnlgc/npaVR0pkd59B9q/9n
oDDzbrFDWKciu0RUVBI4KURBfmaZc7TaG+uqnAZZQsnmlAAf+Il01h5E11gaVkzW
CkIpYH+qA9v1+/c0KS4J+CD3B4eESFmQxjldmwryWzG8wlFETlb8F14jvvwT8biP
b6/zqovti85ZJ/g0QmWiZ/b+u71/AFxCerNAl2T31tFJGTa9xUOf7Fnw7IFg4JFA
`protect END_PROTECTED
