`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4vILhJeo1nhEMq4o7JxxKSoEhFf3fb77r9tKKkf7q/9bfE4Oe1JspTsR8/0H6AYL
Ea1optSYhOcwHalE+tdTsGNRD6JdclERSbojxXB1JxGpBeLBv+ix3n+T5ltOT/ga
J4+uvXDMAsWSo8qTFi2YREmft1UThvC/BPJMItlAdw7nuQGzq3J3iBbcaTIZTF/i
Gc4QMu+L2DBjvaKBF1tJaCYQOcC9BIXAx7Fht0gYMRBt6VTMuY6rpL6ThwlCS5y0
Mw+TzAG8dRP/7TGDF6srlQUS1qugRMkR5u2+4ZO/ZT+t8w2PFGzWzMp6W/I6M6or
z8M9pnR6xs+rgVy9aToTkZKCRJl2Oty4BsbyvjjlreyCHzIIaPIk+Nd95uxt/iN+
SEhW2QzoTF5l4CC/cZG/hLYPpIEzbkMqjpoKh0E4k9mxUJvJd+rND7MrjzysqqXH
RiM2lQKwiQ0thvccegn5GrikPEzk/5eDFm9jKliz2Q8ARpUM+v7jVvlqUuoLWQw5
AJILfxYCGLccKWWWswpGaeRHIqJqV8a5n/YpUgTlMiESrBYISHtaZxYjesrtPIL4
A9FxoJ67Y+bXQd+xWcAMSIsjNlrjIVbCQcBSh4kBU11Vihdpx7r/KXuqocupJZhH
kAvKVJJylroz8zkIugR0p5FIWkzSUYR1nm1eKD7wZYSDrHF2z/sgNTy44wnyLLCH
7mqSbPNMVA+jp0CukklszoR1BSrvvS9Z2w4lcQrfRnKvmwTYtzW13PuUEy15bauy
soJI/NuCYg2Gwnr2MSSAE4LpJrnL3h+ifnkChOjBb6DxZ9+lt+gB21hltblcRDG7
2zwnblW1412IrHiy1UwnsSkpxbnzSRLBR86+LeeEyxRwvjnf/mhO5bKwPJ80xwJH
vTQi6FaVA3YGYv6G/Q9wJhIQI7z17MEl3bAGY7RXdFZncyFH0e9DgxXv6rd35rb+
dbvzVDqnQGtCFjc89N4BwEySpsZ3FDQirSwP4nnm2yGf4Tx4vpzUWDDhhdKiZvYg
tbThRmR6sEaI6RmvGkt0Zb9/8DknhzMCQF14xYI/3wor26wlh3Sq49wqFjJUt2qg
55l8XU+T2ut8nPp7NuTAE4GspIM6wY5AyMcQq0aMisqZN45zxoyZgjWjP1KSJ/YJ
962aDWdsZQGjK21NabK6ETbizwSNKRq66Oaj4/t5/09sjZS+DjdrZ0hZ5GYHDkBR
v8l7FDBehUkgtxoiHOLnPX6khY54YC8NkdczvXo1uFSp2RboXrvq4Byz2KXYMdYV
oJ5WmnlwXvub/vA9v293gEPXOzFUYRvHeZ8jleLssd07MmwP6+ZDCOH6hBkK9Z/J
Ap6E3yeIK2orm7veyQIIOK+faLutun+xzA6e3887F/UrZNuz3o54p/uiG6pVjla/
TSY6F4e9pXHQF/Ce0ZjbfjSnwHEBmFLhzILfW5o3ki0HJ5P/tLyaRFDYm35fIDKW
E0xIceyOCcQpPaMD/NlCd9wvkDuMsyEF3+7fiwGLfm8DKbdipPwc+tsk/b6L+w+k
2+wEDjl6kS1SRKXjtIByLlCTuLvkVswguSSV0ytGXdMBaBqp3w53PHthDc6djuR7
nvT/3mT2+guJFTkZLIJBUOW4D0K12fcRbtvTMvfqraDwtuxWytdQWe+MPBEGIMnR
rZ2n2d7DdTHYRSNFFU84gsYjS96YWN8nwZdDywGccD9ZQa84rp8ieN9hGyePMIua
idqsZRKkl6GV0Bc/c4STpb6b7vE6ACZm9/1swsNyxf1tr7WaRw5OlH+qaewmJnJO
Mi7Rp9OGdR1nS0emjFZkcraoO5+OhIGG2yYqx6BpFRDkHnt1La6A6CXseNeqCBCy
z1ZXerfBg3YNoPkFBCBAmrkWT3YWuxSVlDmv9TL2aeJP391sH186gvpNllcqrW+E
g0IH7pqsHPNc40pGPa/Xq5ofO/Mj8+HKSTHn7SID8Jm1Mx6kMiZsAvRbpZPjKX/j
Cyt/NepGBCvEU8PWJoh7/ExxUgR9Q4crorbJfD5865IFuYGP3ku9ENOgvTH1mk1D
UADmmmyrhN8ss9Se+ECVXb4leBwaiVuUUllpYVgpt0wgN7xlKfTGseRRJAw0MtY8
OD+hy8nixgMTD3MNm3zLenzsWIzr9lEyMJ+3kl+Z9W9DVYyEt/qXc8IRDyhBuDzS
s5cKfq9JwTEAAAu4vDheHeLXNylNs2e668dsPGspnnQh03RfIiKoJ9Q0BL5l0gxe
rpAllT38wLXnS5GhYEKNH4rKCpzha6UGmRkZqLYAnHgbFXha0dcWLfeJTgNICF3Q
maEWxVhkg6HHI1rLBvxwc5UIAzgGeUaHhCWgxCc5foh3HStNvUxt96T2TwlZrZt+
0X51UPIAVZXRlOf6j5SoTvxVv2+WWwv/PXXf3nN6kBUA+fCM8nAcFKnDRrQFavH6
PpWTVL/S4jgN9TIHzhZt3xCudxSq4O4sf476i39emjxpabfuG+tdHCnnU7AxEmX4
4ja/s3ePXBgLdkgj38ywb6xkZdv/Iazym1M7n7w7paNrz3ptVUpJweAW6jwZpVNW
oVkD/uy88jSKeJPLfIAzQCMZ+bZ+W50fOWOczR3xHUBbyJi/YH5d4AigRfyCcDYE
2PpemQChVSiI01G9lPqsrFgVRj6rHG32Yg0hID+L33bl5QI0hnHlHQRMJSO7KnUa
uKV9EbYdc7TtFdhPBjvmPNI3EbAowDyuxEaoRoSneWX1kozWfByGIbWiNl5B/pZy
6oTI1oHgqKZIZ3IbJ1WgxQMIKgoAyQCRo5tPvxvi7nEeMHTm87K2F9AvBfYkJYwu
8cgSgCxim5pBRHOOTf1VvWXBd38naOc7W7a2C09cU4jwjmgwyd/pfi8PwnmjVYHg
Um20zUwrgtJhbJmLswcoapscOM73yGJBUjbQl8px4oOAN4HN5L/jNsFgE9rGkTu/
H4bAboVb/q/gIX8seWXkUPHAjff0I/ad3MWIN1Gs5Hck3RWFad0Ft9Nuee+c6oNf
D6hs+nL1KP5WJMmvgM5NNgqXnUb1ihHiAewBLyK0E5UgaSbUB0C5iLn6uIkISBBS
mLXfY9Ua5Mg3d0oEM/Oq0VikeQRlojMdMZkD7GPFmQtvlcm+Qa1OJQ7/PMnfnEJy
MEsJITMm660shIqFUDD7QLODG31NhgIgvJOrCRbDzDaH+treOr/TrswnsNmjOXjJ
DlLRUY83y9ycKpwW/NxvdLrXX+N7NgpNwvHUfBMonROTlP1kh7ceG/EWiOQuHjfe
54QeLlTzXbHhjo9vFCirF1iHGvTdKtjQ7Jqo/3DQsZLpRuJiMyqLU3nMXGyAJlUk
3oEACVE0qa+HdOzu6AkVahrBsAbr3CQU7m6MmwsT7yKYkrP+YztUCukQ3lSeYj2v
webmhRNWtJvQoXH89ceYsUUnq8WaPBvdf5AYijkq4vcMLzaPcC1JU+qYrOBT1+s7
3/wPDR1ekEreaael0rkWx0LXrsPP5yyW+WWHYdCN7eIymy8w6x5w5dC1NiZjjLQz
QIzFqdNGUooON+CLSFNJ3ONApgtDsvJmNSBrbP8EphChZ5md/1+jFwQ+lgTvcwHE
ZQjZ0ApAPJFVhYJRHk6hjIdlnPsQv2lz+zIZtXnu1ofYw8rOltZ4QQLeTlbzcA3t
ndPNJDfa5LOeSsD1cVK8BNWwD81r3CeBR0GqF6xZAdY712z1F4mLce0+pGYVms4c
nDK0NbbwIvedZ6rFXjK86MXsRmvqxqCnuWSXNNvrilMvUQkvGnB5DRMGyRHNQ2gt
8tlBuWcu111ygskHYtranJLBkz5GWn+Rk6Xkic2UdRhg1X2q9N1JGuK4xgTdmTUB
FBR9bZySEJ2Zj2FfwqhIvE+/a2U3BXVFLbPPsi7GeaCBKS7775tCfm53LZQdRQJN
l+8axuggRW1udcZIrAa3bkjskhPDpKlInEbYv3PRFYornbbxmh9XLlq5yImHy1TQ
UJfxVw94kkfHvRnC7qAU60pTC8CEV3da8fwZrqzTcWJYAe0aDR9Yxw/uYy5t0zd8
r55Fv81O1jDAwB3/gemLvyDALMDnyZ/02Q+R8iL7+1VaM71+WLFLpoM2SkUjMnYE
qsDsXSqhkvJts5rNgYo7j2y+FPPFck0j6O5rHQ08O+P0CDlQAZ6RRFPMGdst7yei
ZQNZ4uc/ferGHYWoHz42Hbcrz6JHzZXJKj3wsIw3bL57hbeWqNOG5X470nDzQR7z
pSNj5mWPVg8zqhf2P8yNWjneEAg6FxisvTOQbds/X1q6hwjMZXv/ZdjMxLNz17q1
3NDdv0lmedl2fX0/T4UnyDPW8LjPnialv6LSOQI40Ag7puM+dWX16U/b/Q6ASi/3
l6fHuxr4xyl+c8PNyPJvUy8iuGfVYGiwbJwyq4nfEBEj6PgkevGIomAneMBbtTJF
jZGNHQ+zSgfDHk8SWgqermDErDYjTN0cny86///juMAr0chrFSLoehrdHPODCN/7
QDOs6vvpXovBQ6xJRrtNoSoZAomR26v0jQ5HFC04OBQkTp4oUBzm63JXies6qzR7
seyk/GwDmLdZYVOw5PH15cpbMHN3RTXcA1IGiWhfSeippLpwahxDwxyqBFWuV3Xl
jdrQ3ZKKdBQhTfookvMVOrj4+Xr4zoDfmmQm0joT9FkVVL5r8d9uVTVZWL96NBaR
J8xL6Pn4+9enIfRJZE2KJ+Flra9gh8vZNOPs/Dg1sBDsO7Vz1KQn77o4n1PtLIER
Ka707ZxXq4ZpLoT4sWU4G2HUXh7OXQi+MX2jANBFMKtLKCAJ+H7u86UAbL5BS65Z
pbDMDHCoxWl1ptUDdWaaE8VI/UQ6t7ssguNO+m7BZY8sCjdnugbkSYfDsUk7ESQ7
t1H1p3DEUT904neMTxDCa2pdbTBg/LRrclxJqVAwG8PoQRCIjZJxVGipJXZU8iTV
qCGpb6v3UwEiNg1Zq2pUzABEKV9yksiKO2DKRtGFuEMbtphINipdncyfmh+3JzLU
z6Sh/izaxYRD8pXmYkfcOpskilQ6HImh1f3+8ZmcvWLRb1Vw+v3J6HI8X1wo3Wq/
P06HC4V6O3WFme0dHAZ/tzJPPGLf7i9sqkps+b6Ze99u5NZa2312GuyYfApcGTYe
QmGDIqbA1apOE44zFt99xA+jGjHfyVXRBj6DRlPNGouG/LLFiB+g4NAYYZD0F+NQ
fjIpIMPR9AE55ZWqEvce8wtZNoWnKkBTX2wjsr5kSu6y21tspBcldHuFPH+SPAf9
z/FMOIc/nCz1cE4aejiM8HMlNfQCwbmCBJYcYFSI27hHx8WA4wAYq7mhB3wS5tnM
oOzYQ+WY9leKGkIYuFmuG9hjs46wDlcNpoSdnvuh4gZqeTQNADFltmR4edTnwhh7
kxzisJnp8sFIWpQY0D9LAu682+gHvnA8UWQL7L3ohnSbw5HylpczExcFJh2gUQ/2
2z4AuWpoZXQ0VhmSe27Gzifta7oOORbvCLWXxDKrqzrrMvXQRadqD2CO7mKDUXg+
VH9PLnow0AJKE639fDptRov2qyCEH+ztrZp5mkTNIQ7ntNymSRPCnJLY0A1D+60y
nEj+el5uQFFvsVE08vdZ14znZzd9kuCugh3w5us4b6BgpRGJcOB7dSASCccYfh2W
LJVtKhBosEVrd9oQuo4gAIPwX6yC6PNgVxZeT4VdUWWtqlt26Ibq8SObScSmqabe
jD+eK+GbmTvjVplIZDMWpVDD7IgTGnke7jacvmIy86ci7pOiQ9eLTwvFC6thQAxw
bXBGNyu5JLdkAtE8gqNRwP96LfMbJL5IEgxUBelJ1D6xUoJVHUyHk9VXojqJZaS1
76kDlKoDboSYPN1Ljbu8Qal9+2lJ/wtlIYE1VbOGCWrS6+DhBpJaRmO3x7sLSos4
SlxbboENHuDnBoDluNox6OqDttjvyU51QPM9TRNXp2++MneMHLu+OQVONDA1bcDJ
OM7kgTdgTB8XId3OSAbnrTr6TKv8kyAyydOFeEDXqV+ggfDbKb/hjrSaHyS/3FDW
GvMyOORBwSR9rTAqye37NYfl59D8/1hwKxMM5ZayTD8inxrYbu/Fmj722h0mbaiR
0iCiHF2B8/Cl5pTzRNwfWMoYqjA8monvP0PBqhz6o9UBQ1lqp7MTigEbDi0z3UWn
ZQCbT3tKI7vRn0uNMPLgs4ppuKwuzT5Q5iYJGkDLpopJdukYLOADGbJo2IM5T4Ir
bLHSvs9jP7a6pKbS5k5Hz25mTD0vgVLiuvnOYOeT66PR8Tu4X9T+DQlnkaY3OJuE
R03AlCcblATE1geDbYwgmAAQ7JV6BkaQfW9UFRQt7hn2iDanS8+ti+sKldYnOo2S
qMePjeeT/G2U4j/PVgWryqJfPVUEWuTohK2eyQC4cQwXC159utDFgd+H5JHzHTo5
dsJYwZMeKe2FHJlF4Ov7fEgonkwPN2GtX2RrVBLJRTRI4NN60k5AX7fGg8Mzv7VM
bv2KX79vdZfMVhyrflYLio1f8O8GmVPIMVO4hTbGpZJ6JUGOqRdN5lUURzbGQwx1
M83gRX7qjL5DmH+4bj1ztlBKXQwgkrh2yYfXTi84j6xhLufLpgNPFrQ7V4zMCswe
H8AoCC8gV8PpzIKbPlRnKXsKYYbw8JDTJ/dz82eTuI76c4YSF2o2d5nQn3K4aZ71
rbx2OTUYE0vTEwvR6nhxihcznM4kio/EgAhUi+cG6kjvGf8P5Q29CXptfFkJuDLB
bM57hJJXYoeUqISabFw8Ivt/nFeGH8wfklAyYdbPwADkduM9t3mbz2ihhNsD8lr3
tXpHXThnnAJODRBl45SrWIEc9XF1jwOFHuUdd0gwtko=
`protect END_PROTECTED
