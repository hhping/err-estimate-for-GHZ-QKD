`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MVQzheR5zcvWZFq6fsoSNk/ezauYPDPP7DoStMX6SWkv9d5xqiKwercvw7QhBd3G
m7cdLat19gjIfITpjrT9ebR2rBFGWmZaviy+TrJowJblEcUVcmHdOAuTtYeHdEze
W2xqQzHlcz0ZYvKEedLIAKIfcmP+PyF3bGwMTQ9ZJcKrCcMVWml570/kKBCXNbJ6
jr5jj2T0XoT3yk0y/oS5P9X8+FzTz0n7k4SGbmak/j/nRHALR0La4pSW3yU16mR4
KqqbjwOl/2GUEkTSOdjqYeIIAE1sh2DSIfV9sU6sgPsoVRB5vxRSIrvfT7RwSfh5
+uWXk4n4AbY1tyU7ZFXTtaTv7z4GjXUnVCnm4s41Os6XpSZiv4D/6BO7Zy22dAGU
gxT/jF31QHoeAG0tdexj9d2oR9/V80UQkrWVTLT7vhErjlr1Trd7xJ8tK64SBMr6
sPsim4gR/P+YM+L1MpG4GTW0gDdReXNOAkTQlCpYPugKIZdNqvXdBsA23S53Y/g0
f2MheKcqVlA/h/dCtLAV0p9+ix0PacSxKbg3aofEQCqTOp0uFNKhanJ/n7uKAFrx
dZYSiehOl44xmEO+8S24ToHVGnHPZXofeHAZWZ7l/qZLp9UbNLWvzYyAhPFu3WrF
PP+hiZmxF0GvIbvnb+y7hcnKBBjB94EdzICE9I9tL2gUqJCwSiqvyIeeLYFI1cIf
zUw2vExWPrTJwBgdMGRZN2jCpuqr4fgbGIuI+oI56KrkxiCXQjSLZ5ohaZhNtONS
l+3oJ2DRWs7xscZxBMKdkBuZ8iXy3GxcrbFgqP8NK7r4nvJKzqtSSY98sAYFmqZr
BJuUTZEA0+H/OXhkB4nOE3msg7tdukO8QK9FRJNzdBNc+b1k0KouMfWdRQgg0+Ld
4FpEJhdRQ6cNn1GsBP5aDBh+uFixzhCrh2xhPd3mxBo=
`protect END_PROTECTED
