`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84QOg8e0Wv3ukcRX4djvIoDkbBHigMJi9YN/0zp8wWIFKcoAuQJgU2PyAjoWWGOk
F18TtzeIEzOMrTreslFj+XMGPh6rmqV2ih0Pl03XQ0JwEKwmRRulRTj07PaoxnVn
xyx8IbWfQ9T+AvS8Mv3+lqk+9Q7G/blNhZG476Rl8wNT+GZd3aS78OKvNCpJ33wl
oKK++NI9yrzHCcw9K6+yP9Cixk9eDA0/7RsvUtOWUVvb78U9maCqFSSO9YtSvqxU
aGf1wHpMrs5WIIHKWmqtDOz+Mth5DoOVVJyoEJIOfGmY0eNWgUoXTGg8lY1WqPr+
tk7x7KMBPXLftT3OOuVbwvccUz11CwZQNQECFYlnzn0hclN12OShyzeflO50ehl8
3ZZuDRByBJFyeLxbXfChcTZ/crtAM507M5CEyFe/zbS96QDc6dg5mljmFa629mU8
FcJ1G2IZlAYbI2Fz7YXmZ3QCV0aU91WeKaLwgT9m2rjT6jn47zCLp+qlthAZ6ITa
meG9n1/yJSP4Uqwq4eZ3+MnWnq2mS7tVU1l827qM296RGGsVwLlIO/Xh2OK4zYzN
aRKUd+5eOdLf9xF71/+5pDaWYT5y1nMaBOJ4rJPR9VYLm8Mtv0sepDFgwkxz9+Sy
J8UR/c14ylgfiqjyUkrovA==
`protect END_PROTECTED
