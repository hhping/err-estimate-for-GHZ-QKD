`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkLu7vMlAme/G2WyinwGdvdTrRfYp0SPMlCrGBx2sShmPsuvhSrrgyEG48W5YWYK
tx73lRLx/fdC0bbmNhI/K8iCVAmaCeqA+R2Ob6NbbMkIo7Gac316FlDqz3gxLqfm
dtTOZqchZKfCa4M6nzXuf6r5yYn/Fz3vFe8CFvk3Pa2/nizumsys3/hJqh+UH9EH
VlAjGisqhVu50Vc619fV1x9W/29kMRIVNhfwPWvvnwjOsxztbstTp+VIoxWLRpQe
1UKgWMnnT4w0JJwQOzGhQ7ki4JKxrbUhFirKHzHgB+1K4p+Psrj8aM9H0tF3Jk3h
Uvkr4HQpAtBngnJ9uxvmkvfyCRgdNhIQEctst87ZB4e/CYSbuQYqrvK0mXG5Vpy7
G5f/4l9o+JyfzaCV35ArBJFgUArwdqeDjC1sfMj7uMgjcCcAihglV0/ML70VUkFM
g7ASXXe17GD8gRllyQg7emiY0ZowB4sfQEaJUvpHSfBLI9FNQBtlB+htnS53Yk9N
WkYHGRtLz0Q2Lpz18fvO6shT3urqhcVaqotJfAVxKcEUTaQGB+UvJOgNeWNY1CQU
Qg6KTQctsNqZrafx6R+TtDWLddSLQxSEAQSxIGfs0lxTUBvJfYq7dA5Xh8sUWQQI
6ZpnNyPmjFplRfFJQ4wSfkoWu9TMNEfVlH45t/hTA3iTt2tSQkI6kQu4N/BmoQGH
W5YuyOYJIh6/8aX4uNw7fWo0XH8lDQVmBVOykq/jC8KznoQbrEMUtqxsJtB73Kns
SgrT8IQJ9OokLG84NMPzKAxrBxDux/8c3d3sHmz0faAbDTgZaO7+YjBWdkdE3iaq
ro7gVUe9h/AO27P4pDl6fFN3/h0F6Xn+0Wntx8V0mMXCBOD++dAn9goXXMTlR15F
8IoZK2wjRt9DnJFqQT0U5X2mk9LX7eITmHRM5U9mE/Rj1e3zAvuc9g9hPn0ZlaJ6
iss7eBIOLW9QjcCK/Hf+GRc6F0IBPH06IFeoJ3OJLMVta6fD78NxlMAtByAGNr/+
Zq6uh5dUCil95naXSQF5UdVodzR7iUJ3Ukj+SDd8aJxo/xApHYB1qJ0XuBzuUkGW
ZK0wHixT5YqUoO9ZhSfBSVwuREoZzwrU4CST68gTmomZB8H8+ZUOevNImvQLWflT
xyRXYbNNVLdexKXhB3WLykfekERvd0WLtg4Ur40e+s5pNQ/Obe7t3F9T5M7V7+UW
T/U6UhdDM0z3kdZYFZnYVlhKWV2uXRhoTSz+i368u1TO6rmMkP7Nqi1O50pJgf4X
FaGeASAnHgTeCP1QOXy2ctzfuyykQryV679OVpsweI8uIeWMwBHb7iZ4igI/hRmz
cgdQmeD8liPudHH5LM/3jxmAXt3CVHUxaY+Qxwb/20la8mCrjPpv93azfyeB10Wb
IGgbuBUz3JSjyp/xVEYhvXYoHYfwFoC55KN8aGfMgq7K5mA7OrQcRiKkmxKemE1T
m7UVVINHdYiO/pJLH9Cy05PKB1+vvEYshSvI6tfWxNLlZTE4oGhFu3S43gEVejit
vlx8FtK3zusU1jP+OhjbX/uPOD7dv7KTNdZCJMPr2OfA6oNm/jRd4m7wsaoRcSsg
lj3hzXwaa6nJ776ZdEVNB61h+0fKBfUlrST9Oxs+UKq8tIQdJ3DhxQJ4e8BoOuGu
ZiiEI6XOJRjgJgW2mHpYvobHOyDxdvNouDC3mLYNLenGc4x5bc70rpdnRG0Zb6n/
fwPxN7GyalTJa9DRs6x6KnazTlC6EEIwTZ/kk/N3olRLlZL/Loy0SdsOVgLCxtNX
g6SdeiPakm8hGh7KUReaz+FyQNL6+R8Ud4aIX/pJdTRgBTLRE8fGu0IsQJFXA/tL
nzYogC1vY/v97tc2hHPlsjPT7hXA+QSHZyuOB+bXmVMx6AGrbCLF5s2ME0I2XlU3
dhpTAVFAjZ74slUz1J0lKjkQOP92JF9F3u9YkUGSfbwtkKXf2+mq0ThoKaKVa1h4
k0jB9amWQJ4NJUglM86mK//t5+BxX2el9BSm/xEyKWmCdNgyXtvCElSGRNV8v1o1
NOoqxdDhDT/cnH4201b9kNEFUGUYjEO8lG9Zx6zVtzxnhTH0E3j/BevRuecxrHZo
YeQaVzhizoUKAFaHZ1AGluLp6K2ZvCjRGE5wCQ1x90Imen3Fxt2F4PTvGUlO3OxH
L2A+ZXEGO1g2qsDKE7Gycno1jNuxH4lx/TBReWoWp2zdCCRyuiH3Qps+7Sfl/4xM
eH0gBOI68pna/yd4Lqq5pK4F9FhsIUdFlueBQwzgiibfMYIXG1VhH14rh6hdX2yF
DJwE8hai8WhGX4GJtuu5xtd5ZWJ0h0CQk20mCwo+eWGgDxBDzFbXcyAEqbzOoAlR
dcjn4hgMuwL66LW0Oq7S4+bjA0aEsCsxssO3IMDqDYyFFqFfTEYU1rrRqWhYVaSw
XokZy9Rdf+krmVzf4N24qfbxrLXWZZjPUFwbBn0q3NEv80VND3SFqjpTnjwZHdtw
fGM/fW5JAAEwZyC+OeEI8txjkREcZ48FGbFGeYNEJAWouK5YT/fL8LCRDqnrx7Nt
/j2aue5Xpkdm2TC+WTwe0EbWaecuMNNyZdz4E5TYYWvL4Ykv/rDkIt00+zAoRH6I
TianriMMG3GdU0EYz216zfuL3d+1YygCp01tOhE4dkR/dt6h3Cqo7DzJWeJEYBQT
9UlYkV/ohsNquDsRmP+qF4PK3/vhcurP2tquTwqRVUmqIDerOyXySC3rAXocHXff
C4JM5B0bH8ZFoLsC7FHFcG21igczK9kFgXe2YIxZwIuLapTdvVniSxngzShcYiEc
LKO4hhLWT3Zbe21vba02tI9OGiusEU40UY484XUt+sIJ4GCgL8wPZGm8zoywPBlF
4mC0Vh/E/i/4y3MkbBlDEUeoPtRoPkdvVSvX721+I2gtG6jaf3SWXP3aPe+8sHQF
UUHE0wVbhhUYMsmM1s+S3CjRXl6j0oNuT3pPP0dcek9gaiy0r0bKg4NwGWqD6Qit
JagGMjU06hE3yVCtAYNbO/OAk2crpKziEXcOQJMkaXtUv/nokBvcE7ovMVPS0esw
SjdsECe2nwoWj5mgb1LiGBwQ+gSKH/JSoXzWEwN678f6l+XbG4ITP5vpU2DeFaWv
XtvJxRs+xBNCjBcYdl1hzjusXX8GQrSm5ZYRZG1C1SqsteB1U7EtEJ0vSOUazhzY
W0l2/AYHcPrXx0wGQeNOBiyomFC2N8W5ecge6eXw8r8iyYbw8OsMDK8uu4TEmgXH
mniGbNbeE0K9RB37AotJ/s5Tvvo/r9J95kbSsTgguYXT6bOSvAoskEgZKA00qev9
EAggjNa+0EFRCbPFOXgVKlBRAq+Eq8dmwrxV7JHbCRwU1tcMLxI1G16fAxLowsxN
nm1bei1TnpPrgDtTNwGFKGkPFSz2UoidWFf3J5azCo0WSgLR6CcQIbCVL+uZI9d/
G8Eel8wg7JTzGCSyeVuC0hRNQm2PwFDjecxp3RluV7UilTa54+QZpZcYExw8R7+0
zIRncodHNod3QDUxHYbEkXwt7u5M/imnEzRaYpSZL380tQ09D6jf7nGB68KKavau
bQCJ2FVBky7PJVe5sWGxf4T7+MVk0zBsfrYnCN9FdCeQHZs/yW4Q1ZvP7cIhvyef
ZAT9s/cnqHEZfFM+S8HZcX/W9jkgC18mQITm3nA9kaCaRuoC6jsOYekoI8NTeDEQ
kYzeVvFo9Z9bssR9FP1XaWkkNaYv5oky9vFfkZKlsltdoWwNBkUyEoG2b+JrxGgR
Meg5JV69XzcP1cLX1G/zwE6LNZnbE2f10Daj0mR6Xx/zMk33Oeoqu1DEX7+zHzXg
0xB78h12DT5ULDS5E9QLloAFcfnLus4CFw9dbJhJ+AubzFWO12oldPHYB8nW4FJp
lznN9tYGGl0ZxeHF7L0UzIBZKWwD4a+oD49SmvmIja3pHNhy8AhKnjDr0yRATbc7
sPYQj5Lj+GP0LTm80umci/8d0fvRJBGGN8CAACLdfMyae8U/xioH5b9jk0vjgrUk
H3LOzkDhUamHqFNbrj/Xjwnh2nNFP594eEzP8Z6vRbyG34iiLo06lWbBRWO1Wtfz
Grd9QrS07S01IAj9C5kkrppHc3AEmLEAwDYF1vQ+hso/qNNCTyDC11nNZlnvKGie
L93PY2eP/D5DXVuA+/KmwFwi24Q7ByrxGbXCwMBmtGgykfQ1tawTroFY1DAXostF
B4tXFCrp5mACISTjTuW+8LXmwnX4VP6LIYeprkvp1aGtsuZIHg3RZjeuJEyDLrfN
g9yUYYLWotKWW9OlS+VLU8NU3dXCVmIpatg+DoFMLDOzql4sEbsAxaBmhQ7RptHj
fIppud52utfFG6DpJsXikfr/xN8ANt6PRd+pOkDWRitF4akTTdeblHW5MmxgVTC1
74Kplrj7OaptL/uTYEzQvLc/Bth+0LEWZoNUa880Xmu3TaClaUMs18lo1FjWEESf
eafkCWELwdtZTrlcq9aHguMKHqiZtrn5x9H/r1rK5xE2h8noOC/qW7MR3+UIr3fM
qWCywcKkBg2PAE6kN7IBUK9gRzvWk+/IU6zjfizCx3F4q79qxNCQcSDJJhVxDGnn
TagS94t/mIXSPUSbSUAd4aRAAW2cvxsCmGaIwAJgcSK0cvNY6Tbf9wqyIormN/9a
tupJ2mUpzm3tv8Lll4v8KMXivayGUWH1DWwdAFnRoCxECVkE/Rt6oqEJxcMtnW9X
64SuXkcv4KGQxq1rSGpCoSO5DEKO0ZcIaOWnuZyj7n1Hkm1GHp1KIdWIX/2iR2LV
4gfQELhd54zIAkqTB61nMWI+f42rgj3Ya87qApsfSqrIZ66V0NOOjmeJtEVPx4oh
GOlr1qQV69oXo0wn984q/jgt3rUXJLsBzQNLUDSaJFR7KL647zRXMj+/q7ewGWkx
0SjshWL25cfK9u+4o6THoVG5OeYp60JJp6xCNbskcT/OhAjpT/uoRV4PBA42YG+x
1+SKYc37JVz8tBMKvS2VJYKgkDqHdC3U6CUF7s5rS/saZOjvtBe8nOvhTP/aA/F6
ix8Y7gtv4d10VsB/HmyjOjDXptVav2W5PkjjUbi1oGKR8Umf5pL2NbsHA26hSlwl
loiicd9HU3xPxVoiMDL+Jff/8zq076UFvzw7+b4/eDGRpCK9B9MjAjBqNb6HuMj1
1bGQqSdNrlerHTBuM69oYhuvsKMFApFQKrGyiBXP0fW+XRSXOwSxBLJxgH5oTVOK
CKZBWrsGZjkQ1Kx8e9OIl1x9h9mC2RvdO2cTNWIbiAl5FumZ0ObT4IQi6ztynC1v
jHF2/cL32+gltjHNh+QuXOQfTkItA875xjfX0Hu7bkPU0gXhG6F6PQRYox53FEtK
caSWmZy+tVjN9ee3tn20Sifvh1Dzuav8uRUJEhRlFlUnxsYVIOt7UWgUJhx86zpi
29lN3X3SNAb/wFSdl9QWxlB04AKfEOpxpQc+6ACxkQnDJUOOEJD5lwy14WfZNkZ5
sNwz0+TsgGOPp1suzWyGlzCJFbmzhl3u+xLfOwuSWz7C2wtfv978Iy6uIGj9tmNM
z38Jak9sKKPgFDY2zDyhVQs6FEmLz1ovtwLFGPrrfeWLPCVoDBNcw5lJSw+buTFn
rcUw6fsWyQ/IeeD1nAkY4s9xI9KDZX79P6jH1KbqMUgeyEUVXRJpd9lP6hENJwRq
itY6oWpFUH9DR7dW+c7yEtVQnlsXT4YRTX7T6ehc95PLrPTjH8hx+Vw+uRcwTKwE
LkvmmuIXUugLGIlk4SxrGjjm1BLE/wbktpnbuv/mmrsPn9n1eTtUTPm3ftiS/W8P
F8vmtWQChT0VWAsuUbkfTk4IYnABMyPzHCgDAqSIzh5kdJPgdVFumnul2Dtxyn2r
HJfjCd90yxlpQS9BdNPR2hXx7/AYYoqWAlc+4Pz9gS4E0W1r29Iy1re3dpKzdoJK
VxP5HZBfOYNzY6IoPP+jDsF+df7DtK8aKLw3wQnn7mxOrdxAl0Jm4dQUNg5kKRVv
rT+mGy4cPElDoLVPkpXHjaaRo+ZP1z0JUhULfS4Gzh1XArzme/DIHq+gAbArGS9f
CLsQSwrUb1rFxDb476n9QqobiPg/P/2KmOuX06PffPATMKEJOQHNJaae/VQCQ9ds
kv1YnhxI3fdHJzX1aJP6/haZjMU4Ax3V9Q9csX3xEYFM2TcGg7hbQwVbw1Iivt0Y
Xf/zytYYbcWckLZBAC2ehG1ld2/x416E3l2NYSiWNs10xbV4cn1En6LtwzT/Ffk1
2Bii9XsG8Ea0FuJgI7XyavXEcdg2fO7CLMpWXSVq4ZE6BLTc4eIch0s+y6AeVVLe
uKQMKgb+NEBjyUj3O/o4q/8BojZKpnMBvq6ON/9oxW2D5a7DYHzAcTpQrARJqHUc
Npru7Qmkcm8VnzVRyrFiAjf9Eg48Czp4vqiMwB+kWtb2HHgMjT0wA1jPLsb11kVd
wFGjy7Qo/VcH5aD+KcVocyZYkoPD85ivSfebNmzsHmkX8AThwraoA3pxSfswZznm
FOmHi8drdzdTx8E43jpNBNAIVtoZ+KWWg5NKXvwtxt0BSXbV0SODg8DEY40fi8SB
4SZv1vxrJxTMlqP6MHLnC/sSEPtLY5wNEBCk98MJzCTZF7QNkdhxOKBd8mHQMLV8
QXXSX0fjcz6xSc/owTvfFS/79fiwQ6Da7cZn/twP0z11cqnw+cncRD27rqrE172a
7qWL4giSYay1/ernEiUQcWItFptDwQp5ID5K2265Mgi+ZzgxfeBldOVoQ+mvOIUG
/ETizDb1T9dIPej56Mp42onWG3Q9wtqHD920G/NFXklUpIjTceCpidvEVNzihAMi
vPRUnbiUalh0E2T8ndUGBL/5Uu9bGlxScfg5QpJutVdRnnAVx3PXeqGC0NmjHuC1
CQxvVV7jjdCqbVPkYGhNUJf5iUVenWLoVxhzYo4Jp10ymJ2uP7+6whiIAe5OtFVY
G7lUrtu8ukEuECe222RUwy3O03//hS9I5Acw+cgfy0BR3rMwnXu48yldTUztLQB4
xWsoYSuzvGSOjeeQIByUnGzKoN+gJdaJUO0nz9fQuQCcyzpaNA9mu6GeRYxIk6UB
TR54QPfa2O9CT0vxoltrry56UvgxpV4tnGOzrND9dtaWkOv6iYf6M3M66lkl1R9h
us+LiUARW2561wPl99rIZRbmNvS/M1g/vSOo7GfdHtUJ3XaoXipmWxpudbA7vBX0
zwBnwWbuk/QWwz1ViguCd5MFX8V/jHN4Ey98W5q9lQ+i/jjdTweMUlXtTKIvUG3s
QpJ6Jwm74VgERHTYOVHrukYdpxvE3TnU+MRBoySU3cXP+1AVFijA7VoVBBkeWHue
oovIsg2eepduS5vEXS66NbU4UUcYY8urH0BeeRLGYSPETyLsPms/dp0yBzpRF+ew
JPHuKetkW3OsiZnums91ec6BdkAs+tS5sY1hJUQCcZzrlcdVu7JThuAKayYvTb8Y
rHF1Y8Xzq1xiyvIy2lotek5w11A5mPLY57PHVBiet4ephkQW0LrHXjBlW6ZQeVD3
Om7eVSzMHCy3mCL0MGfrtHPGIMn4E0l/ARcM4zeVwyfojwwROr2FcymCcuKepQbz
VpHltVYtvA8C2Z9QmM56R6eRu8/pslCK8T6CSM4y/xJ5EihpFbum8IQydarTyRNi
wF92KRJXhG9nbFnOLMO1b70rVkNqtRwlZFx6FyVloZvu+plA25y4QwprnV7bGlJt
Y60oyQ4yThJKF0rYiWtQ+b7Svod8eD3QGmgNq4smHq+bFjBZL+eRXNvMRpJr0IoB
N2C+qaBWhsblkOPZlFACcFTrXzASv3iPllGOe7HBDHye6lSaA6nbFvG4LAndMZAR
Q/lbzaTH9TULGqN14u8Wlm8ev4F8JUAzEvhWGXtvQapEALyuXeTIj1TeoeK/TsNz
GRpU6npf9q81/Gz0ZfovR+w7gWEdtKIp5m5UsuiyBPqgsBm4lXqp+YTfHM0ud1sX
dxQeWSixJgEYTjsyiLjrqmn57Y0KUV+IgPKYypxTDMIKH0b9tZg+pEStpT+8E2GC
PnUSoEa8zR2DjwFAyyMlQHJcfMusOpiLHZdGU7EQGuvXWR/WLryHQP8WVfAOKWfr
nmRGdu5ahv4SflFN32zM8NB7EuLn3/bbpEaekOIdnnJmsRN3OeNZhv7qzVnYbeXs
fK4BJvEwLwTzHDG+r+F6PvFsrOuWlNwMRSdDRufGm4HPklC61ZlzLLbqnEtM9+Ih
wu4eAKLt09xK2OWlkw1r1RoOuGDPBYGSe/5HGTMDD2MKw6jeDzA40Tqev2XtoSCa
4GYwk/jWB3jC1TIrqhCfv2qMRbcJAGQ/qBMFO35xqp7vVtIBZP1Q+qwqhfxiXl8j
N+2LqmuDTc+1MSjaOxwzJ1aQj77D+S6cLtT6F5GXuNXksEqQmrnCI5bcTvxbGN7J
VWu+RPZsYszWGNoQHXT7lEi60zVvHy9IOHzMzMIL7dGBp78Qgs86g7mJR2ME8Iva
asFgASjWXZ9zbDCpkyDs+L0GCx/CdgKRE7PUz4cVOmLunr35uaA8/rW4ebl6j3sf
0w5RRqLy6MUJp9qBTkc8+oMcA8QeYlZ8cCAInT2PWnGuSOu2W1js3dBfmwYX6taZ
3KtHhFSLiiRYwaPePY2+y12Pj8FA7Kpzu6ZecIQf2bZQlUGIQNVn+Klx3tbK4nYP
IDi9gg/rsydjB0HzTNEMDksxHHoict3xy34AlSOmujgFg70Og2bR5LLsYh+6B58D
55/mBhy7A762uf860rVn85TWH3u97j9J+LdgaRLXLCAbn1EqkUq+7uebsA7c5TTp
P36ZsFztzE0ypUCD/zcGHwilLMdPjqEvySMqzHUEJzALVWrUjardakJ129v0sKaU
jfRwfDnSFdn+wOSqj3p+hDkQ+1MuqZMmVteYGglkcZTWQ4PWLObDjkC85yNV3pkN
PSlWXrnMa6FUEPzng0DpQ4v7fsArlw8E2LmwgzBIyLhseItaQlQVKvPdkGf/PtPU
7lbKAMZnXsmFeVcWkXIFABDj6dfM1faOa6l7Hpdit3xdQ0oZnPfthqXpXPavfvjJ
Nts7jn1F3mRMKWZ35+QdoxLes04LMUrMNEQY1AOeBlwpy//udv6ylan6JdYBuPLv
PJfmNK1AF9nP9n8t+r3F5Dtbj6xq9PpDb4QN0HBFDaxQQoKpEoC9uZeopcRKkpu0
hIv+/SZoec3I7juEwQIMIGC0KSFx5Ei5W3DUoBM11n0CvTOKIkxET5+t1RdBHaKl
FdA+p4nk6Gi5aDkKlReD+BlK1Nuj/GVEnzOUQk2b5MVnyxpChbZW+TPF1+w+2QrJ
Dy9rR9NrXRdyBOLYAUbBirIRYcPkTEN2Iwk08Efhldazyo1fhviK8ZVi5idf8+FQ
LrL28LjaRcwUs+FIWdvcLtPqzHRglN7u5fAtpHdyMk/2TGMtkxfqtmwjK2UGfQwo
5Ouc+PJEnrtBmNEGqtx++uduFj5CQ3GNOdXkEIaOTwVhiWn6wMULL9f+Sdyez9XZ
VSOMR3xgU2FZjrfjojkMT9fxc4aZLs5RVTUjQw0qGGDyDHN6+8LO5AjLYNtwM085
G6BD4oDRnoXds20lhh/4cOhBPGvTWwurZqGGlIictZR40UZFHrG7YDXjRDGrrEhE
Y77s8GnSDXawmdXjY6SxpgQftbqkAFW7fDbRMAoUDWj6VBGanKy+LqAw5bvhC5+I
KFIAZR5D1E0uyt5AqB4Achh/ThNOjFVrVIjDjQWNu6o2ioifU64cQb8hezuSAJRu
O3lxnAL1pimz+veHssfRoaBbesdXR6qDxD60+sZB2DTQsfXCFZJdXN5OXiyOcn4r
+r4ZqjeFSeNTBmhazmlxMBCRP6OMM3kNT2RFEgKWgvZpHvYjASOc9eYjbD4oR0XP
NVhPyiUhhi70grSmTf4c+qYWdTr5CeDTMoINuzQCfZAaj7NzgSEL9jBcy/JkedMi
7xPxDjtvn/nLRaLJxK5r/aj0R1uLiohxnpYpSxzmYzF6Cd9G8eJN7PpsepINiUMk
lel+kw4FW8LsPDaTfGuEJr3TDDdvMNhsxexNR5HahGrGO+aMUN776b2CGxYi65Mo
HHYubeadPVrE9vwD/z0IykL5ELDylGw6THVJ5Y97SFf8AC5bjMPef0tEo652MrtB
i+4oueE+uFnKr3F16cg4G4mbs2FW06DCINF3LKuIYiGOcSpN4d2NN5+7Fi3ILhiM
J3GOCAU/QZEb/RcKFk7tCQkXf4nK6VXe8sTz8OP7gqeuhCRQjpxJq9y3rPOFIKqu
uu2TCJACCs2ZCEMJJzag/KqcwILBPxdmQZOYspa13hn18XjGp/M6Os5RO0uq2GkM
qHNN91iYSD5l7HkVGdL0+9E7G78aGf+7JM2eQdKGPEBhscPedw1dzzLQlDL9n4U8
KQdEhx1ezbBtggTG76XghEyQgLTv4ehpI6DGdiIX6PasQUp2kGyqg+ln3l173TXd
ufL0teFBQKcPs4IDaB84NKkwKu2zo1YTLb3FV4zRNPiJoMoIyQ2zr+E87uEutmzX
BtQKJ5ElI8PRBm2Jh7CWFaVpwnyFolcCg+EE2Sfj3GXlOcADBV7ybb2ZBoLLJqan
Tn7vzQOD0y21xfTwgZzPXEsQWTAxTgB2EGHs8pcXG/HtPqH6/r8bw1HMdZusI3JD
FAa3qzedrh5vqQ7SoMtpOteh2BqmThhYbJLxUcy2CZgVlIR6YAiHBzWDMpfl4GNe
ZIbQk25VVDaBW8oxA3eXvm0tjM/VXxxVcwb+UPloiaX3GnW7zE99kK7eKjy/MFpN
+qrlQRvKrmPXVOtKUba0Om/9XL6t1Q0Ai0N4BoDbqiLE7edD9dtkq/dzJ4toDEoy
7Qnp958e5jYz1Ixb6KlSIstm+PwfmbOpB3/JS6iS769jP8nV7JnTokkgZOqLFJqa
BR97/tg0NGzmGrwJLG24h/pJwVPsdVJ7L4nTa+ew1KSotY0MgHav5Q+NrCozNsWN
M3ZOeARwFGzm9Cs16ngy9mBk/5tqapMNC9SsNkeoJI6naqEbmJ99y2cPIUxMTZ9b
lKEc1S3qDzS3r7NbPiDOYlNlX1WTafDl6Ri5QTd5jvzdszSBMIw5J5mdp9rAOSOM
gjeRVOo50syknkIxGDZ+3+8L2a/MFmLxHDlgpc0w1+PI/xy3jJ1VTx9eu57gd32N
+JLswf+cZPR/fDfLS86/R0Gh6fTgYHVyiq7IWVv7SgS2q843uI+0o02+FCrZJJXo
tNJRXeiHiTAbSmhKIEOop7odk78t4zFTFEPWpKYYbzbrrn7prVCoy33mof0WGVCp
XO81f8VwB3DRcUg7hF+10VrD20Eflex4GYWbt5z9hpCg+2ZXHQbHJGhWWkoM1q1C
mpOsOI0MdftpCQlR4Pq16A20Ci1m4c/z2AGiP9BuToSZI6lkRWJ66pn350o3X4d/
FFfYCdOpz5yE005LDr+c0Be7HCwgiPcsARlxOXQXK8P22ytmYrHhNYOq89HhI7+c
nI+seqpqIow1arIKkjBEHTQS1SntzC0hGXnbK5SWZvauqGObSxRV2uRFEKgt5uKu
DtgQdQyME8x/tsLiOknVGJZJij5mCCeabpYS1+rxv6lKt8yz6rdNyrJ4+Qp4YnmM
Yu9BDByxXL2mDP5i7qceFS+BrnaNIMMqIr9fUPRm9VQYQIYRkb1uLu+j4MEdVPBE
9SSWn44C2Kdk7weaz8zKzfHJhDMXycVWqYR8k8v32MiFh3dRziUW1LzjhNTmPmdZ
gpge0antvQuwgIxsdgcKvCPvCJKBoi0Xt/IEW/4XFEvQQV6AFi5T6mkoP6APjpIR
6TKiGINZQXqYA/sB3jJt49K0p6l5p2syX/bDaHJjnEX7IJjvaA+YqOmhq4rZ4q9N
C7UH5XNzbmMOLJhfvH97G0gNz/L6qbmGl41mdEgUghX129hixjpcQyoVuC9ADas3
bAetChmrlwdNqU+OqU2iA0HujA/gtJOrx+VWIstr7kQ/E5B9R5/AUiGW1OSpek7t
tZix5D4D+c7+QFbX+A1iwx2GTVN8Av5t1ZRtomO7u4qiRn9D3ShGCKftiePJgPOo
ZYwTbqOc6Os1ffRQsLGuixHhlVddmJUCJdrBwkeS2l99sS8qYM+lA2iuugiDtwhL
0GrIdR5Cy1WjzQeWSEAJSfjimEIwRRVhSFs6Vz/lUgyhNqFQ0jcI//SpEsIEsumy
wStfd1bpJ/UJsKWhN39oAwyngABgICUPf084aoa7wWwqVW18o4UBeOsWHaCBYa/i
/5hcwP7NX1xYhVy7fzc5Jg++41alAPCag4WEnbWqXv4egNq5LjQUeq4LqCc/TlO/
gdFFofnTAgzEidsY+bc0n4F5pYghGG+kp8yfXj3CSeMhmKj70HBinanK+nm1xkh4
LnvXjy/bIvELbhtnnZXqE2gBSR4QgBEBAy4p8X0ZB/U6MtY2MSlO7OtkoBaZ3FUE
lkhAU54azGySTinv4xuAcH1DP7C9ZCg3gzOQsTgRAZ4V66Y0Njp/3pl6mweASRVy
vGH3g+T7LOWBKIWAaaV7tsKt9uJP4zCom6gpjM54Q3dLlPo5BV5ZX1bWtIh7K546
xLbLWqpMSYt5eBxGq+Od4sN85MFrdgr5TcDRJH5C9iehfogoSEmt9Ae+XkPoKYUa
AeaaBLxOVnvbT7Tvv7DyM/V3sldaHrU3+PNleeJfBuLRUleNcwaWBzDiWd5X6a1J
RrraQXTQ8dIZZXmZLtyfcuxYCyBlD1b+ZZwdgvXGUSB6Wdt1zoBKv6eb/84lQL+Y
YdJRvJKbQL0+JMi47bTC7HVapy3pVy0tVP627m52/cEFPdjZrZdIvjZhJXK6iD+c
cLQfB5oLKPj2nf0Ui05Gh01WTU2WNwa0cp43wYhti6IGAO1D7vbR2/wV4C92glXB
4plUe9uyoFpkcE1g5Qch/wfxmJJmNvZ2ZTDgT9GvaDoV0eI52cItc3yPU6CBK8HS
4fsanin5DrOhhJvuAKB/tLPwxw3DrSKMwU1tM2XK1KXyBGxRBn49hXFMYjQLRDNp
AJjRN62NynU8KduyKIembtZld8wZjgXOMaxDf+mWLHGxPdWQuqRh7ehNLq0CXaAI
3tUW38zZw7OoSMZtPJ6wLresSVewZ3mM4pIgEk0fPYzuonaF7S8jHFA9z+aq6Fnb
NIJMyjZZ4jKrvZvqn8+YP2HYfEi9U0vVYaggxgb9xMc5W8I66t74DZrb5Hfzf3es
ljeeh4HWpBpZYNU2Yl2LgyA0akfLDQKM0qG5gDsYCV3VXElFsBRtx96oK3OXmiGY
9Ctk7zPkf9dPv+jk8vUWQkXageBROYYo90YlwZMJ1Go5ON04+t87XPSARyC2r/dS
HTiLGxKIhv5y1qUz/fG8y64NAEaSS0fbS3tlvik7H2XLpyH9gdwY0ehANz1V9bxA
o4CFGR1gVKgfsiaQ1Wa/MDNoEn/J/EpQ6HJhsAJ2z3TFsGnjSTtex3gcm73ISv5H
aT60G4Cz0/ibwM50ZlLVoreEbmBPiT1rKbJLrhL2PKOulM6nFDt3H/ttoaoiRbTD
bRnsJyx6KEz4Z67cGtAs1JJNM+ybDz2SouklF1MF6Vjriij4uPHbZD5RQZMDS+14
iZsYu4Wl29swvphYPYzozWsbpCZT0Zd++sAoYM8KKUk2y78eOA+Dt1wRiCniu4QE
OCwsgerC7+p8IzPtwY3Q8G6+NrVLJsqg8shg9Nf/nC49TlZHUlER9Z9lZsvfYpgC
lfMdlU4coAlwefxSMqN5+FlgYbWOI+QED8TA7USJ4gmSJRRnkuy1RnMjJRKQ3df2
mJyu7WkirF6Yrt1WyCVKSf7cnV4Lvoko+MZ3HkiVYOlv71iSXsOw0inejW8AOf26
F+WDopnQuImAwxZrsh5zdu9xR/yyS9Bg7nu4yCjmm08FnbYksJ/sVDZdG+buKqcm
5ZMamUtb/KCiT6QS6ehcLzyXRCUYnlIIf++8PTHG+ElgMLqDrQZVYpus2A2hJgyr
OYEMSwaYWjVvI4lITrgASlnEOFiLQdgbERDZkVqpeZS1iC/5ukN2uI/xC4iTXKtb
6OHcrR7sO/0wntWB1PCwDqkR51hHIJmy9A477XNdX7NMHgU4BY+I1T3X0BQfJXwd
/vYfnUNtcVAqfF7DUPAB9D0Z19IPOv/ejpMuBO4JwCgbJDY3w041wpwPodeymKul
0ISctd30eWbcDvPZ1ikv/Af6xi1QczC5gMabf3806pOfo2cF7tSdmuZHFCnk7uoK
Qs3Hqe+w2CpTzlUf+9XXQik5El38hQk0RNy98FWQwGy8YHEN6WT9C1p3QYYvV6lP
Adnf+uGjptPhm3dYPA5yOsYHbo+rNYdM/E54AdQItY32yWulFLqUezjlqsTghAjl
RRrBgjdJxSk7aH50bJVy4sbnyi/2LH1YYwPwo0aUUvagL0nN3B0LvUw8biA/yN34
8RkQvONYtJl72SSsd+45R7FeemLoHGS675vRhNZUBf+Rguv1aBPRtqntlgJGTjNb
5mkVAXyVNitZretTVc746SOagzjxaVdyBqM4HVcuWydjYc5jssq8kefs2kjHsAyr
SbIJfQBTrpBnJEiBWJU2MwoYwKglCIVucF0aXAmkni/OaaHlAVuxXbSMU31y7QTo
MZTTgFs6yfSm6vZIqDkddlv98xutsXNzvsuiLI7W3NaGRjYkZWPYhPSq9SJsYL36
sttmLk2gc3m/juol0UxjLf40ns8srLQ7P7YyCVGNt6QcEhpPYpSxOEPWj8NtPfTe
Jlqp5NhPvNPqmYqbC86GhQ==
`protect END_PROTECTED
