`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TF0qh+UW5QkTjkBDsI7+V6l/bcs/tJ9cQfTP+oxD9pVkH+shI3hPDUPvA7x+5nKw
7qaCa6uje+oTVayfBktWnaLMrLtesyC8FBekjBHHDp6ahe88/kFGPVlMWaanJ2IW
DIT9J+IOFbY1Mx91vTPgKzYJckCInVLDgexZQbPzvnkFzL2oV4ZJyqUEMn4FDvkq
CFBAGHvR8+MTv83klB7z7ZoewcgLvePvgtN3/1k+fHCp5BgikiUYPoFqHJJpRcAW
CE8GfHKvY8qskfbw9gc0k1AGogiarl2ExbgxfQvMROfFvvUAQY9ZmMfw+tAqT5bY
GVN3vpol38sdSbE3RG/rW44buVa99BsImVYY8xQX3j0rz4dZpbRMElVCw3KI0EbG
vRIIgNR3YbskHvvXHWwyvWaqPU8k+rR23VO/1gwOC0U8aztI9N421n/Jut6sS+8n
mnV8ozOPqJeK63hhReN/QdhcK0tMpm2+luv9IpQtHV3/d8yBGUQiQbz4NOsB1waR
EY4rPyxLbzuxx3CBZN7k6LQoqh35JZKzXzxJYlr2x2KFS1iDucxbg8TmS1ryYdHk
4tAA+S8qSCYU4UAZX+5GfG7C376BDMh965Q059iQFQRF/tYBFI1cSdlmZMUQtj32
vQX/b+QHArkU85HgSzOkJlONCU3BaaGJNMnP8mbcCQdgnoPOvo8n1Gfze4XmKqij
Mv/5vjAc8Yy0+Mc3XonAA9CGKhyC/8L9K/cIGVmvyfR8CHBg/gaQjYzCKPLE7J7S
7kFc327UkIECxiWzI+0ukvD2565j82ahpIflUDtnIDEOB6k1AzlJcCSt9FzfsK1f
H1ARkrntRqj8iugb6YBp5KRK16+Pm+74wD/vDOxOAf5eSCXqhPAy+VJxshH7Tjw/
kuO8yxmsv3qY9Pt+Dos8GKiBMC3/XkJTkJuD7sGVBY4l8sbx2XQFtqt6TtwtksEz
cqYrm5UxM9anVOrerEnIWREtxBOS4uh0VmSwP9dgN7t+c8sMc2BRb+dOmi8qdPZu
I15cV5MEngDFyhnt5E0yLXrHHnJEB/qL4jAE8EljawY+r20uZoI5XMnzOSmcZDIm
`protect END_PROTECTED
