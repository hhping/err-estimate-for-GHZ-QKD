`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WuzonqTgAaL19CYvUSZU0NJp1yveXjzStRUUWkcuBSKnbejvhgyka6+1OLytT0vR
0Jix2DXXVxQDZu9ZOhfCtN8kAaza16Ss7b0PQZXSkbt2/yVJ+wHVlLMhf/GQKMT+
lHd9EVSNC4kdo6xsr0vB+IbVI4SAlIzwKa7pbOMurkx7T1AgaKwW8ZgD8EF+UGzW
wiaNR+zpJE10kSiIN6a2j/6IDcvAUXy8Hm1GpsIxkhV2fQyshj9sEyPUxQAd+T6O
QFxb2BLZEpRxNAWfcuLqzOwKRW8+lKR88eyivKZ0gAws2DHR0QEdugT0WqF5ubVZ
jTxUJVwtNn4BOJ1+DDufFbiWAMqrHWUegH3fAZVoQ/4jrcyioZ++b4iXtU5aL+zh
+9dJZISsBu6NXZ3RVqkC1Q/a0Y6MvSGTDSTplGdnHhYKQgTVeYeAPlLNt8y4pHXv
nnFAzeANL4kstMQqaccfb+7d9HsopE4mti3IplDKNVLDuJIVMF6TYnKHWd0ipXXY
0FQJXeuQAvnHM5ZGxlTjPlOE1CYjQB7iYjz3Xbz3PTFjJgUs5F7pItVt8sfLHHSp
fjWaV84uR0dQty9s397yxQlLgntruJFtLpXRpEtxqTYPQPkgwjbdZy+Mlbtdit8g
DQ9Lgwzj5klGgr9axVcKXGYK8/dZpoY19UE6v/rn0SI1wd9oKOMx8V3JOtOAjGpg
sbril2oOsI0lUVsNPRYK0tr/KKJ6ExpAFVMZ0eKoVXxYN8AsSqfTWH9BbRgbfH7u
k9vvfTWDfyLuTDpZwgdlDMYghfQMk89E5z3e85AWNSz6KN3MExptOAQm9KdiI0Wm
GDtYH6SWac5VzgWp8W2QHX4uR3DNG9UTjMvTREaNrT5YvT8HIy+aaIHUQ6Z+Up7t
vtBsFXrFNUOcwuwI/kvOyLke4DMgloZtCzP29Z1q5leTbRq0GmXlcbNbZZM8hNnj
`protect END_PROTECTED
