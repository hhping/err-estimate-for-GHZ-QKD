`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nn3/7uvOsQsWpvPtNZ/bz95pUxYfikpQluRoHuRHf4OdFW9SOJVkScoZIi9DdYQX
gxLwgnroZkqoYr9ViKJx5GFURx1vc6vnLme8uJKcc5X9g8vk9hoE+Z2P3EEhuiux
ciEd7M10lGnjv7ZTOxcA/wcP3jfHnmmB8zO9LZTFOwGA2MdlmzPQwCAkf+SUTOHP
gu0PIR2xTJxWYlF4+vAfzFH8IIhC72W+qXzE27L/AWndclILoR3z66xI/IbHfKPR
H0kbXc8KclpHYlOt4ZBtuUq5xCwPVYVhVrBaKisZoFEbdnQXu8Rz9iL1DZ8o6JkB
klvN1+xHpqM5P99fHNGD+UKyzdZDWTp7PMJVtK+4TBHkMBSAjw6ER9ThDx1O+z2W
aTu0a6XG8hXyrAmJ7jokjwTZS2foBazAw40aPwO3YToj21mPYyHjhJWgKx00AlN7
1OaClwvehCM245XaDkZbc5cw+4FcQBX4de9u3QbIclobSb6kZmOrmoqHFrsSBx2R
qCb38jVQVmtpxsFW7j6LyAWA+0hKB/HqH2vE2FqcqRZ0NGohI3nuzdMJALxJzF5j
yNEhhWQmVw1xqDPgMRyw8w==
`protect END_PROTECTED
