`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wT4Vll5A3vUBlcy5o+WQBYuaeeMScJAjr9F08VT83Tb7c0XyGfiagI6zFacRKxY+
14+y0mhsKmfI3yzX/lGusc9JFcpoXNXqyJl0ZQZw1oH7pQfoLc9cdCKPdlr7Mj0h
9QQhcGO21Kzh09Ef2LxRgeuMvC9Qwn40mEBQSr93U4Pd9XtJ+u4Jkw9ZfMEX2U2g
bPSmO8Fqecr++YsmWKc8kpTiB/TaMF07y9sQAR6D+gMzRMaWG/2OEpCv2Qr76Vmq
zshpIHhTBRZWKR8IlKkgYq2ERbS34NswVdgeyUYe2YkZKCwmKvUsryQxzyqzm2Zg
R8R4vjEubBwH8wiBOhyoSbjK2IJTkmdHf3i8ybADsDBNoD9amPIRV8wp6zekuexy
P/0HB7igQ/g4guaaCYoNepBhZwcX2eTpNPlZSEvGFjuGu8mDoh4ldRyYtxQW7C+w
KDn+KRI0Nm8apJFH5ucsczjYn7PIlqaIzzmLugO+JwH1xXVo3XnbZDhiocA7ckd6
sRtmBtRo4n08C+3qK92ao4ZU4vQ6NiMjtNw38tR780wyM0HHrCU/tMqt7HBJBlK4
CzCAAlu5Ug/wYqwt+xJR+tR14nPAA9Gz6oS4eEhsS+QHFf0g/+x6XjsRihdCOUYF
y09oXoGHMRqrhyt5mfEkcaJkCv59SBCaiWXIH1wLYcNRYk7Cd1NHcsKQT7w91k0P
BZnIk22Y1PimJWb1yES8syLWxxBVc9SCSaXmYZu2kINP1IMSZuJalECSifKEIXrX
RzQ7mD2y9H9B5o/Q5vmFRMOuwPPEq45tNWU1uyFNI4X29s5CCFxcmv0RlwldNr6d
HUed6MFNUILLWnkt1ZTI8cazB1mS51OENm6ADf5946BSiVeJvFKyaR1TaTz2ejhE
TnKF6vWlyUkdEsjimNLQNteVzCHSnk/Z+PmPYj193tvZ7aE2s0BU96U7lBElZ0Y3
kIOoRqE5MpgtKpjILQ33ABNE8JnwceEnyUHoiTz+HKtyelN8fWSuKU9Vb2Gi+KPF
LHC67C2wWV1D7DLMxvry1XNKL3jByNH3le7w/7Jrbp8=
`protect END_PROTECTED
