`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6xGUbjTBn0v30mp2XJQk3Ut81h2hLFKDGGNoNAi7MdVOUsEbcFsusK0sWXUjbu+c
ieazFLX4NNaPnblZaA8sI8L6JzxAumRrXx2ATPY00QA4pNtzoI6aVejhNP2x3v/z
Kvj+7sbSvxQ5SX2QwVFMgj7uSgwIAciHwBKoNtvEZgwg3TBoyqCQg6M+Ls8scyW5
qZtcywE4Bb+NTxbJF2G5acWRhRM+OP9y7U15qFtE6GsMVcvumEzGaB6p4VWB0+o0
UuAxwJXQKpXaWdHhq+RutpOaRVKGE/q9VIYdSLhq0w6WPgoQcvV2NdM5d59q7F2e
RwxU+3qoYcw33ANZmI8EzbzAxjAGmxBVw34eKMctjtwHVhX/du1XEkVGLPA4MaJX
2cOj6IyDfjfBb3FH/StgIwxw+QJXdLcL2COk44F6ERs3dM0kfAaSWOx2cz+5ZGVq
dzNDfWneQrK5gNpt2EJGMUiWDVwADlTysAa4FV1JGJdz62UAA/zuFm60bWFC+xs8
ujO+GIDXtj1OSKtmklLHxRdYl8XMW6o1ywmkXmGQfPmoZfpEyqEDRmmMM3e8oMBU
M3+J7a/XMQZQ2K+eMZgHiXEL/JuB44XpQHTNQ9awwXv8Iwb6srDnEk24y3M5+5At
jyVfPCyee/pgb5lbKF71otLTIWX6uXZjT89WD5MtESLczBlW9+ZPquYTg8IGJQtx
69jfRJ+QE8Gqm9g/K5rIscKM3rWxBdFDpkvgcDXEmxn6UMCiQ7CoRD2C9nhpP6Uj
YQ0liQo6b7rN8HeQHWUPj+zt69ugCkL5peh9U/VjAaJNAZcuhNNg/53i21zGPUmb
ynoN9ZcUwUuWl7CH+v4puriUNhb3lFOw/mGoREY7uplPD6YCCPAgB55HGp07n0x1
CjdKHMFUC2tnD8a/XlFEP1P9kXdofjIbu7pcu8iZL+7JtAIc3CPDsRikg3qJr4rw
Dm54IVgkLP3CxWzPQ/k3EHHikpEJygYBRm3FnCTtZpMGvLyX3rZePC+q13FnWMyw
UFh0bGMJE6Suv0H8GBEy8vfNg6befGRDxnZbJHQVdOICwz4KOCPy7ZOJfdgqf3AU
Jw3Nan3tKjFMvAs9pkX8H8x/GnH0wWz+PHoTF/2Te1NA5fX9GIPzm6Oq0xIRZWx8
Xxf++9ew/YrbD5tU5rNvNl4Pq0ycFGQYXwBxv7OdJCXLXWomMN2kp8jpLdtVnBae
GC7z1hQMi+SPMjR33qS0vkFMoL1R7sMo8o+PCe+dli4+HiLKye6CL+uTA2cZUFVJ
10XOK6yiz8VC4QG/u0ZXYvKkAPI1Tdf4oZXDQyQfLM7vgebxQQi9BFBeQwoWrYC2
SkkoJyLo8fYmYIwVq6lTt3wy1XXJk7decQr7vly0GZxA05mWIY+a6Q4okBSDuptO
u+H8wnHLVF1MOhV6J8nZW59fesXDLDrfODpbtRVG+I1nKiZb9f9EQfbQgLmnN4xs
fwDKWIk5PukjDhMz1Qg+tAZhoeRYzZiJPDai2mMiFP92aweuZ5zn5XtIc2F99AUb
NadtpgTuSs7c9QnaDXMinbo0aE6eRvbNy3OSWmES6hBicYnU+pdzCXYl0wfhfz8L
wm/T9kNb3nu9N0dIVUklfht5rtUqfVw0uQX33RGi47VZbzVOhy2mSeZXmREKc1Av
d48XxfzQlsxVTRYVaow14x9r/TP6MfsLdgHMk/YvLP20nikwIG6HGOWK4no656Y0
7OVj0mfZYZPjVYYd29G+wDsLDmT5vxYDVqQ/+uzRchOUVxMQS5xe1+mby2kNw/gM
4j37wld5pcYdowHCTJVLwF2/dFasEEpP8tyt2GqcHbJ93NzH1SmhpzqDJcahI2ml
mGEdTOfii9/OJcVjfZFWmtemf0Aha26B6dd2XSzxH3fyMNDhk/VuMkf1gTYDaKaR
QJDMjyPxNIHB5EBFXf5gpruAhNJY2OGNDxO9BpQRCpCuxigAwFz+/SOaZvLa/ElL
2tv4J3apSc0Fur4DWeIPoyZC2JHVIoQ6S6SbSymk9UjtupwLjnFKn2Zw5JlI/SR3
DDSVhylordrxtgConl0p8So3inwF8qaAFWneSr2tnqn2c1fTaTf2yoT9lHPp00Bb
BGZUShOsT+TfEh/khPPefn1Wa9kjDwCjOEF/tixPRhfBnd6yqIHZy0AFA1WZiFBR
ouD/H5M1WdVpOO4FjySYQN3p2J28AYgONfZe6nAlpyB1+5BEeafltraT5sCTNY7S
3IPwNbWpe6MdtBmZ/w332Dd3+/B+PYTsI7wLmHha0pBZEJ0XeF1r2I04IyWHobHg
5+IbvUJmk7DC7sBwwuOHs6xaLxRjJe4GEr3XwnxaiU4hCkBCjemY0a0I8oOh6xwY
+uOtx+UTedSBmmGj3LtEfdjIrS6SfAPNm1nbZRPLKoxIwNrls58Ln1viVYXU2E5+
T2RFr8ogHGdaXHZCzxTAZzoPQaava+LsBRfDUGpQhTuZ7P8p06vBwsriRCpCPvm0
Do6yNpV7v7IfjllN6PjG7fFNAQl6QoSk2D61GcaJxbVu4J6qS8uoif6VuMhBwtTc
LZNL1QjnItOBsMbqz6xpivglhuitD5P+UJtfqE2k36g+BP2ElV1Eg6AQfTdxAr2f
VxFeYKX5wEvvKir2UdXjCJzHyn1EvkFFzF+//dpn0UzW727234DPAJJ1KwjnDo2x
VXAX2dDMKvUwiVmvEpdZP4oH203DqTKHZgWeVeaVnYrKgikiesz1b7+EIEm28hx+
yRQzCnsjx9EwhPLvhsixrFY6AJwmWfxdZI4SysHBuK2IeGz/7o/Eerz5MLtk9umR
6/psenvZo8QVvHJo2sxC7RMUh+sHAvF5TXgmnJc+Ma9QSPHn/GUE0e2KLRqYeprH
l3XJO6XORmpGzX4XElN+2apT4xg0DwKOIbSdP9KqPnTRbjcv9Km5GbldPosyRjcP
UYINcd4XBRSRtu42MzBNx+izEapA9kCT7tP/Sk5BN8IG11Mc06y9g3Lzs4ABvoUJ
eGf8+BRkz3EIZp4R/lenXU/RoT58Y049dcRrv1Lk/7aOMWEcjc3qesUzeHD9tPrl
4My71o9IgIAcHfLHLi9CMH7mNkwRkk7h46iZoqKiRDOQs/YMYGYKLN1xtK2/58x0
nWtyuTYMVmhS+LCgpgzfVluExMzuoJ9IRH9GaO4vrx6l71A+Onl4SVMjKauwqIyj
DAvjgR+JXm/teVWbaGFc73U2ZRzD3/Q5nvMgL2pIujMgy2lJTYIiySkYudBO3/ss
nka8FwgeudO7boLERiEKIuxzrCrA0UIiAslryAfIs3G/2PnKsNzZouBTVf/YrVgR
Qtrb69KnEq7Ewp48pBBpV4Vk9vF8hx2QZzGeiwI18e6pBH2tvD7eU5sKlyOY8ZL/
1dZwmL9bzz+pIR5lBShRstDeJ1SfIFEQSpK4zDzX01Ba95lmrLKKlVKD9XanwAmh
ROgvj2p025lgraCEheEXx4hq5gO+ahTk+8+9d8kx/0BhkRNnqib8gJ85igB3dk/v
GzxKXXf0L/kXCJwY2/EOt0deySSkDKq5bIpShkdrj6wjPQjsPXQYMGRwpnirChTH
5sJZsGNEqCpg5r7RVmCEFYvyVBUEDOKBNbU+V5ibnh5oCpDU9V4+18+kJCPushON
8MtcMhKXkDx180BrYBbKvvurLPbHdAcpHZZ+goT/dddXWhbEp/B/uE2TU0UI9DyF
G1qdF9HTBsybvvMyGnwq24dkIf2nPN6Sb8oc6lvM/36oziBldldIg46UEc2wiehW
MpmFiW+zcMccFNfnTIEcW3sbq13K6JRJTMjwKq85WLJV/HBx+bne7XVGBD+lXF5T
iLyGkQG4X8zOM0TtwCfVYrIb2WZQ4dwX/6Bg3FpuQ62eZ3EsXSMfiDT04YFrizho
DmScGIdWFf90dkr03xoi3psZJ4HfZn8RFhulGdlzNv70UioiwuHpq2aBgTG+0niD
pZgAzBnPNDaXf5XGQWjjocEHnKINz01aLoGVpaC0fDakQ7iJlz+2/4MXvyZ3g0Hx
EAKMYeTpVWH+bAunP6QzRAKcN4yukUSnLaty1gaTZ7r+b9gXK3iEQn99dZ1ENrWN
60f9SjVXVar6xOS64XYuZGVI8v+2zvGzLVYYWAD0Hgb/8Qwz2BQaJtMIQpfRc33A
ahG3PlcWC5/EM9fqUgp/ci/1bvqWVZFgi9g9xXxPOaQW1G8uEcRhnnDL4TFyB4jQ
6Tz3twjM1zbMRjwM0tQTQ80SzEEVgAS8K0WUxVXMQT84ZhbsK3EOXSI8Ii8SIsOw
7rB0nsOOwvNZd4wEmmumFdueiMEBWLjraumBfXeYX8X0lbFNoe723bXoBgLMVjgk
mJdfLw43cJPZ24dwFDRlGnW6cp2V1C2suIM9n85e4qqxJZaWvIQ5KhlPSxu4mH6Y
j+pyRTwxqZKkEk0m0kzDVx1CVtBbKUbBn8hVX7ib+utZtrTbHKaH0ODcmpupJR8O
qibpwbWfq1Hzyjtq2fVDL1XSXk1Ij0hP0JOGGmnjU+NrTdl7Ck4EDs8PvkAsw9vp
9AvkRahTa5TdEQaG0hEz1RfX/RK/eQVr/3We3SN1mmez5Gj7XZNonEYs3SC2BtBW
8TK9sQx3EOrokA/wfBozun9fabJe1b5bfx194zCY3fL9kTde2xBB+2vbbJPdngK1
TNviQ+a8V2/X0wr+oFOUn16KwnnMCAKc1Ro4TelFuWuD3RWrWPe/TtHgYFhZqgiC
J9AZwr8R9SPweZ23wLUxf+3miSnOCbKadmi90SrWVtPAXwCc3TWsBM/RBPOYZGNw
UAoUGxON7RszKyPdDlkAE1VoeBzvlYwEi38qkMpZgWx2BwISZOMw4zZKHUh6j5NA
zyTNZlfCk1pjOSSsSOeFFxT/3kji0gdo/mhSybT/8YAbtejGzKnYX3kcgxbFW/MP
aGgKISChV7Hp/nAppNwkt9lT76KvbIZchpVwg0IfoE3t27bKa4inO1cDxtRh4XaB
OZXAJLgm6Qn4Fw+xy9QQtKaATN1qYl2P63cK22u8mmrgLKis2o2cd1xf+xpdSt+Q
I3oaEmVZQdqkwmZt/WFuTJjegfiThRfmt7z22FIGHB4qGiNIcDhDsadR9BYD82vs
SiQduE/POJ/DepMnMZzXml6ug1e3r3rLqtV1BizNOU6K5cjfz7hXIwTqVnx57loY
kFzZAwJYRdUbAOqii+AQifl0YGEoFA5+FXTZE7UUNS4UC7UtNOAE9v9GhApxjnB0
zmLYgyOrLLlYLMD2yxgWQrKe3j2Rcq9lBIh3uRBa1PpTt5lQ5hJd2UEX+cqE7M9b
YuXtuowltluV7iN6LD+ZcHvhMHbzBFMLWC4eD+lw4NR2ngFTt2xYN0ms9Fk8+t5u
fH+9089QvtmdPkyNnvj88m/9xjxZriQSTR/N/C0iDpjqi8uhCsKDGhPT2LcfwLhE
QwnJ03MWQRvGThSz2IkhKTf/nxHKfZHbXjf5KF6k7DqGCnApYU/Y7UskOs9lyghz
K4j/mMwvUbq+D4kAfAziaKnnUavlbxItbhrJoPsyflOWbAVZBUjqnud+gBvxSBni
8sEtZuhvUYDXDVd83b/oFnwKNeFXX/qZawsd9lDa6Pwq7F6hIFyhW4rdr62WB7LL
hyp6uWzMzbd58vVzygpJdDIL7dVRh8ynrsVRUfcgIV+BPcejgSepyruh7s+0kJgu
252tqNwbBktrKejDALnVMyDzrZBigc0G3bTAL+Sf2wV2Mbr/cIgNRpA4Mg+/Ccqi
n51cfWjo2KEL4K9f58yeFw43LoRc4hIEf2n8e4V+LMVMSNGpoY4RKsZdtvowoBHL
wjGjP77iaozj1IR4cCJeIjlhJ/8JT5UsAUWwENTUm3Dr3741egiUK6NeiXAsuhpo
65kh+UTxI6Fb9/SCGGxHcmVtvLBLEmcw4wwt4vp6gn+OqCZRNnqQssR4zoDQt2NO
PmfYe7mJAqjajp4ZJ1a5jIzneGu76B9ctdWEXVT2QOlT6BZAc8E7RgWmmazdwqAJ
TDeiQCaEPPBtf9uaTPEzgWHQowJe7kbXmMY5+VTTr5/Hrq4ZWr6Ym82JwXbYCqYA
9a1Z8efhm+026QjuJPy0XXSxd7cw3De4YIRWDUAK/LcPJG38YDTaVfnG7Vp81NNa
Oq+y1Un3DSFQzUZZ1SpwXp2kvHMNH65rSZTg5LM6Z9z7MnroCQhX6dNE+UzqSNAE
X0XnOwCaQU7hHdd4Vy0Zo+kOCkxvVyCrS9zsonGkYcTV/hDJWxPnERdMpD09UGUy
OIocTsP3DbL8uxxJgjSM3AlPDHlsQKfYY8rQKcXQt8d1ZtkEk3UlUQ6axtaA1aGJ
SkhGo7XNUKO0cyqxxDd5955TJUQuV5AOr+XRaIVhvqOIhm+PvwKhETZOxTTXvxz4
IZwR4tgcN5bBPSYpWcHt8nndVayJ3rZOtXG/WFPsiQd/vjFSQD4BcwZXKU1ouaaD
loM6I4VQFkvPPMFeRFbbOtFolKg5+M27+mSkkU/+knqQ6ym6yIAM/+tr4FIzvJga
mo6RTYlNFAuzivbkO6XW1mepB02Rynl0g620M6Y7nQFmKyd3uLi7AMYvUVtus3YE
PTIXa5UNazClPzVgFAio3wBszsr6QjsDe4XBL/t5quQU6l8GZSB+SQ8o11JeCIEa
/hxbtJt/hi4bxK2kcv+sgbDzvBNA+1xaya0Nof9sHF+FJvRV13gVM6XQ9s9fA1CE
elk+XVtmJGzwjJWwR15JXiYp4F2Ypww1AcGKZDHFkkJ7Byu772ZmpLQRTll/OhS/
vN4oUU6udMpZZsb07UR5MIUdLbFN0mDtxcjLMU7dqsVBJzvv753Xv3EynCl3H1M+
WqnA0T9PD6G89RAJugogpl+ztlwikTmb/gC1r0iQaTw3Q3GBnfXPOtyucJdxOxTJ
GC5bBJyNqg91YvjXWY4MlGvMWv1bv+7zeJ85TB6udfsRdeYIuRDxpyp36WEEnW58
rQ6qQ+kUiI3jH8cJGMnBTQV+YLhQVQAMqyu8IE6aXQk4qC0bgkbK3PxMAiq2l2PV
SyGnnJ6tT/KKtsL46oRbUv4MvnPMDuIGu3VNxWCI64QclAVNkj2mrrCJnmnFa5sw
GiKl4jk+jEM6c9+6HYCa6T55fv4xQ7jb3bct8lJdtX4TsYjglWUuuvmyOHeuMn9V
458GIDn8dmZWCetwQ+0NdDauRKCOJYb0tjB2QKRYW3eD/mQcODq2jU3QiAPXTSgG
0oIMGSwbS8c0uOfZJcOc9Cbaknc9OcyvdF8Wym1jPoTr75SsdpFEPycm+14LwjaT
56J8qAAplrt8XHdXyO0uxemt2qGuqGQSny1azcmU6Ur80gRjHq6LwzzkEqQA2MHu
RyYRTeDtwCBC/dcqTDK+qVt0n1AIGH15kwpM5yFThU8m39RZqSsM878N42HrwNsC
NZR93zQGAU6E0A33RBdVFUywdNZoyRH39K3wMNSLV8njr/bsqeoX8YO2WlaUeSTH
sCf29MJ7g4fL3Tqq4BEpuit2ijcU6zgoJpQnBw6Ra67CdrDkJB0S18EN/yQIjKsu
nrlJkXHdBh+i6g52jC4/OBNJde3d3ZCcrJF+6K9o6TsIs3ONooqw71HQxoeuMnWd
HOpVdoFvNRWketqaAWi11rmrnJ6ZAM8vwhN4y5ic9XI08ZwUxDctSyy26JuDr+eE
D0/yeXI83AxXdkAO8Xk0Rbb3uObejnPyJBEPJbDFbMqrujuInQMfuxsG15kYUAgx
Cfix1GUQFdwnScqSofI0U4gy6cUpOcUtEREV2OzWuAq8nNCn3hsunDW4Z1qdDgYl
QPeBKlqlnsijppMQLqXDWEjovIz38OQ7+3nuCSJF/ecrHhoYGCcvQVzAG6LqNlBO
kUyYxX3KF/2eeB3uESSxzoxloafFczUh9fj1vAegyYKRN8Q7RSsQrDIrth2FKXBH
ZtVBpJCoAqUXZhjsSy7As+PRqN6tHljXtpSd7qfXpo512iPkScvi02VexgHcwO9p
Hu8oXKCPLgwpkzt0KFJfsXFyUWtxQ4H1FT6wNzcjb6E9ou3Hl+KpMaC/CRiiVEtp
M9rf/zDyOjQX1CqrhOJBBrE3NVApwFh+lEfE3GyncoL1kcFDnY412RtRYNKWF63I
OiyhqXN2OCPKtYVaERx3bD7Sgkhl/DvXAJ3fMHoL/ktXk2lzSfgH3JAPllyH0MdU
JVpUTbEeGKQHUE1xHUE6mKNPqzIXeTqEk7eeewxChkOrSjeGpwLQS8LXIdoHneN+
b7qVyzDT8FHM4lgG3fuGQ9nGZ+WFuK9zlUQ83h//PaPOWY5fZCdWVU8xzvam2kyE
xLDgX7RhIdp5dACVufLlFAFUo9LKiv46VpyjXn8uOjvt/w7Fd38CydPFByiR+/XL
+FE8ASGl6P9PqGhSNT8PT+Hbn8MK9TJdp5xQfkg0XD/o+n1yO9cVsgqV6v2LydcR
n1Dkk4tahXEw6Mz8E/zoYISw1u6yAVrOSXV8ko/obvjzl2GgeeaFe0lACS3MUmSL
KGX/L8EVyQSMIJrkbFJMQGP8qZCABqoJo9NoasfggqO1A1+xctpSGsIgAx3fX1Kt
NjFsf2ymBw8Abczyy0b6oS0E23uRAw+shjTEmsq7inwpoP9ikYfuIPLyQZGBjO3G
ZXIEjlqMM8rgc4atkqBZV+jAIdI+q+0pRdZOknooRR4CLPNZP5FxgKPsBeaKSPG/
SPhyPIwxeJajIq7KIbeiy1KaYYBox52GCuP9ErTALLV7Q/s+lMM5YaYSH1DE+gQX
fhBI8ogbXfQmLTn1RqmxoOyM0vKz84HxNj1UEZbimvy88ELTEHPkGzNwjwGQEGsY
BuUDqhkLqL/Tn5qC86NFmNA0U06rK2OV26+qg2x44VfWlU5aQU0UX6KtCAULEMIs
bLF+97W1UuJb8gA6AmXh2LoTeAAPk9YLnwseGMUCPWEOnWBAkdixgTLzA+Xerms7
zbiRv/nb2bV3AJQ2h1/Hjwrwy1oS4cCSynR+BiwXVGbLSyfMFYuHQz4ZwRmK+1KW
VcS920P+bpS2F2qr9RjUZziD0t5o1GYK49nB7/LlsaSpuhDYfrgb7LZ3c0hqRMnb
C3oLSluhs6yxUo/rJzGr+KfvST6AumzqcK2rRDAa/kBRs+TBIQlTW6ZlBTTVajdS
bEaFsZz1xzOBISUYKl4rfQ/th6oCZ1L/X4KKou13dhaU4+6xyrvMH99riGyv1xvt
AG30MDJZune0kNBaFfaHzP756TNVs7ylrhbmINIE3RJw4uY+mqpKh19xQjhbDQJb
CU3P+xdDymnaw8KZ5u6idL4fk6seT+nZn94d0Iekvp7BIBPTiqA1JUBzEcoYYDZn
fOA/sT7EXul1JsyusJ3gaJ7KBCOCsrZdo+i/1No78YGjx0UngRoQZ+SHdPnIkX2N
TdDahPCuVFfjPe+cpjZJydZmtfgLZxVReWXOEFb7bKgN7moBCbszOKyrj0av45oo
PR6okpohhPMHGt9y3DeGb/1Ck/V3dAz3f2XpWDiPVxMlm71cYXhnqk0Q9Lw2W9R7
K2KRPJhUIWDHN6eHFG+fwQc4FJ6rpBfCZaf6A4kcFgbd0optTTy71N14oy25qEMM
lrJa2WVE3e0/UooKVes+/E0k4UM3LBI9hnWKeIQYEzRJCmWnotDl0bR8mJHwDVeZ
VTbSFddSgfLH2/hkNHJIlEqTsz5fCXtbil1vHxR32MUIIMM1dUf+fAlHDlGxxYvF
kE1K435tlh4tW2zshp4UZK+QXJ0g+d6hhyIxw3nE3Sk7opCi7YAdAY5KwwFswWV9
a4DAfDgzfAcqLJW3M2D/7vzpsXtKMQDNwsTEYlVpkBRoAiko0CDmgxOxMu09XWl8
tkDQJ8S6zJR3owqE3sV/5XFUqfEt2OMtIO6cVTnOyFW9whXaF3Fn+uPpnPl1iYHZ
fgVMSuM3NVZXk8qM73cyLj/2bQnaGaYz9GdN7hZZqgr20fY5tbVxAvo+J3xqR6n5
3v1aoVT0g3g6vYQeKkDuRNShd0QQp+Q8PkuXyI4/z9Xkr8858QHBpR57UPKfSqyF
2yy+fRjuYKtEbY5NABnLjDkMf2smyP3QLTvW6sqq6bqUEKTdpMxqHlieceofMN6L
IBcVP4aQDNH7Xhq1uhw+MT6Cnuza8LBsdB1Ysw6k60Xt7FZ6PajAJ4e1NxUsEg7a
6y9Vbgtj7OwcPuHuaoxE4Jqpjz4Q/lLMFM2+7b3shpWaa7mDv9C7iVlO8ZtuOGsp
rPaasVWBNE+KzgL6mzwFEQ/ZPMQxjcnyX4ST9cHPxY6Dd6/f3pLhWMLbUhy/A+z6
pL+1KH5oGxbp/qw9y+JaVvArwIU6mLgWtXRoaT/v1KrkUTyUlxnY65JLXKST1VbL
oZo2JiaKx2bK2mao8u7l7+zBH6BJUmkk1jHzLtWP9jaUibUZ0ETkn+/Isf0EuB9E
cFCcIOi247PkSlw1OrO6SS0yZye8NIDnmajU3WdwxbS1yg1e6OE+MBp39TF9lwN/
PybjJ8GveMarUUTqPRMJbmBTEGvH07NdySJChpIRqCw483hZGG//94TigXpiooM1
77SxSxXglmlJ4Zbh6WVRezS2G30c5ca+7ZQDUEjIZ4QYKX75qlDwd5fjj1ITsBez
Sz4Oxjyn0eraHUyq7KN6rzs13hKkPdVt8Rrg48Jr0OJNlWos8cVifdlj/IiLcQ0d
GXgGxJVY5pNKWa15DjneDckKT0A94w9znw/eZgn3MBWAhxx8XkpBpSNjx4J19dH0
rcRsywMYWK8clOng2/zLtl8GKOArbhX6Na7SbVWlcnUXrMzanOQ9DDoZo2jD/OFU
U+uO7K0z2pAsHt7AuRcj/rUzbBccdHA8X5QdMpjswEViRhMWXJ/2l49eYGwN9Hqv
uKaFifZk8mX/wbz2bCPzsYOAo6sISW7GTgFTQFPL7h0C98vZGClOkLhPHZxi5Gj7
NepmhRbNjWMJn1O2mQYH3MvB8WyuFXISwXHbyh3AD72hSmP8mtV6YvZbOCPywTpw
eio3XDLRWfwKqwpsuLU9GrEcY4IRsqEUTqcIJa4j/hcCI2U98QFz+LJiDGxAWRvO
mZHlt79c+sMPANQDr1UaD4Kt+LI1IDIq4GJpWirYTuGv3HEntco0/IfGy2JC4NKA
GnNThkfVs/zz/oKAKUzcs33D4SIGu3ZFaGs/F9zDyzeoMHbAU3Qaz0clPiXfZK5h
5I6HhZFAEmabc1IZ/DW0pHaST7KPrRysZQOoNqxG6vPo+aiMS/cLmMOqr2ISrE6l
ostAH/ynlZjq6wWgGyLYC1xKXsrQOQb3JJk8XhVagE4gNdEam5zOpnF6slzciN3h
6TYF25lt/FWoG6CZ4a5Kx/YxkL+/xa0MjtO/3ZbwoDEeXeD+JOVzM3nl8LVSUX0h
U+eIC1XFhkmRN2QtJt7kiSk83Vwmd1CmMIcUIjLBqkDNcy/JoWQaX6sRXHsdxNI1
D/LcElu821z/HpQyOuO/BvJSB/Tl9y1+gz6hAppSK/k5V7jDfYuPw7C9BD0z+HjS
ysaA+KHlbX2hYiEbbVd7b86UD+VvWu0186Z0DJ+GNW6DcYyYO1ga00yvKKxCCq4T
kwDXDSHMJw3LDy+QZDi3GGtbBZWUAYWM/LqELL5Nmtopv8bQZtxj3m+7ZguSZmDs
ieqIuHDKGm9lKJ/NWffeA9M8av1ptNBqacg4GZimFJndgkpDZoKHngg9NqEsvvEt
3qGOYImdgRgAJvalKTyv6rqUrxChoAJAhrvO8PIm7JgZkgmpWMHfyJrNbWLNNSFa
EyRJWwueFz3MKtz8tGKL3KHfHCOOmAzr9Oh2yeDLHlb6vJVTCU4//sb/ARFpSj0T
du+2X7KOgv0AM7S+Qpm/vo4PgH0X9kis3GMjRx18+wcBsODLAKu5bJ4pTFnmmYMs
qrD+l51Wnmc5N/2vRUpOof3pK1NXEoflvxyA+MxzOPuq88mwVxXGGFgWLtKQMBj9
6pI5/TDJBNqbgNT886uH1VTJy6yDUO+Bz5Rx/6V29XayJXlCLWOjTHBt0KhbF6UQ
tjrtRPIQ3s/MKf1YP9FNN1U18ksfImzbjq8s20UtdIpEj2J0UkrQuDdX/4SchIxq
EDzgA5nt0i2vjs1ONZhdkErsyB9mTVdGOa5nc2MOY/Cq2C95eBMT8893+SauRa8D
8mnr5BOSqCy/LLo2zOgNbuy/+O9RW2vaaCNZ7YdGlvLqtHu0C7jpFCiULLyXJxyt
lDfN1sMB84yaxP9miG1S7tGVEgcWAORjXrMJ+BPdSzwuqCpx1StoudhuK5LSESuL
Afoyu10lnUlcBt3qBpj6DofL3epQdQwieHMsL8dDpVnRw1caeHxWV/HO8NqLDs+z
un/cgCO/FgUslWF6x+BGQptHLvtW9tXM8uRL5cEoakrsbwvH3Pk9wNHL6vp8jV7y
5i4XVqoUeHlJiO3FX1pcG4263xbMNnxIt6XVYlvA2NSK/TYf4PoH3t8RN7YdyEQh
T6UlK3oVviUgIdow682ksPapqeki1kotUkKxIqHRhrLgKpe+i4pIfZKLMD7t/JZl
kc0zoSgiSBABPGYV814bd0i6mqob8cDH8ba7c7x/m3qM+W68gzFFcoZKnKk+gfNL
Rq3YXm3kXXM21ZGS3GZYDRcQrFRWtuJFZjwwwyno+6OCqoHbEbkAgQWteP5rt3+2
nkO0tzAObYTVYYAdG/Mk5VsEgGR5mgoJigJHn4Qavm6/0CyYiwAb+q+P18swpHW/
CfK80aoJi9TIOaNbcAhTmDGH32jhSrrvTH0waReNhpeH7F4uf0NlnT8XLNuRIk5e
ZBNvDb7JomDUIJu2wQSkecd7R/tvduGWwol9pDPRAOdAArkDLDRyzDaPUZpzahHK
wH15s9Z/tMRw9zvCAWJWKk1rlZ/bf8uE4LvpHcAOJ1WVwrI87uHUciKE0GJbufle
px/o6TdvfqI/NEeFsoUOnfUIBIYEbDEL9kwXsSaPPnRr080989O8E5q3FEW45DBy
a8agnslVfqWEbhFAXH+/X6Ej80SzT6EpDOXLSyBSUbxXRidqGTka5Ap8QHdwRI1h
+3N9vflsrBvS777s0Jgog4oktYgfNNltV/cwHCfjklDhNJRJyfSC1t7xID0ek7Jw
dOI9twroEO76izTYUTbwcDYSpHuaE3SDa0v/WuX+LBlANEr0aJxGUyeMkvHMsxHR
suwNmXBpWFkHrMIfwWClXSaqKMH+4EdKAC3fFquW0DTYeIHqRnZYkFe/jIGbPJzC
f21Rl6r4vVBRXhOzfuKkpFDhj+pPPqJV7Yse172cQ48IviYcPXBT8epD9hsQ402m
yphHzHY/w/2G7BbDd+WN5HqSnoLbviTQKd0vaN+Ei9SqKVIizVlmuQj2nIu9yNzB
I5D8BMfeIGYjt/YChWwTEvNPKSzeSHQ7jgQ/daAcoAxs388gg8y0LssfzrgYNt25
eEGLBgJPfZ7G8cpD2t8SV66JMqpZJ5UPDOVe3H7zzvcckjS+JLwN/zpi7hutYRjz
a1l6+LFQeYxXnj8YQ9C1Rnxe9hi3XlaSDPaesd0LBT88D8VUth+tpotkFsIVT8OT
7oTiDAa0xAy/4uP2lPFbQhWnmraHc7ZTrPU1R96HrDjp0UdxAujfdRialEBXkT4Q
gx2JmEeOYZ9yh3OfufvDKF0X+I1pteB02hyy/wpQAWilAxEuMNcYDWNUE81aMNEs
mzlBgfSc+M9cojeGAeV/o5Vsct5Ew9LKkNeworKFgubFvTKfcIlebDHhOtsIdwsN
cl/b+h67uKUxjcIFQYfKLkqfbdqcrhqF62TDfJep3ZwrHajrWNJsKSD2A2QoZW8B
Z8mKV87Na1jWaoHZeTXenOPO9hGZcIlPe9PdXcf29PpjBz6ig06i2GsFZunrS2zl
n7yN153sNd03ks3IGiuuMabJueciEvoqQ/ERQ2F/kdaewCxrU89FXVYwUtltmWvl
l4eEeVOziZVvSS0T7GGQoQuHDw9+JjWj+9K8wHXEOVv0XDULzej7MX4qb9yaBzd2
tTDYoFOYhG2YfkyRIC5MSfDR6sHp+GlmAjqLDADkUbsPizqjTO/MUFSFeVHunnUe
R2sBz+WfBgKcp/Lwj4nAZIyln04QJiouxdttKG4NTIQ+trZRcF5xRsEDfUnLYEft
uiK8H5EFwWIqPe0BG3Yn7FVhruHAqgy1hOejqsN5WvK70GB1e9b2XzwDWoYJe0JG
pPBGN8fh2vBM1Pydj9grsSS8Fh7SlicHl3c2Q2/+0exNOVLRhNzAidwciiXyFIXP
zRlicyp2Q7DgxeXat7QAUsmGxHl2CIb2cc5AKZl9jZZq0ikJa1Bq2pBaan3AkLZ9
apX+QcSus2ONwRET8hu+qUg3bvZH31AvCTvX8Qjxf6st7bVE6HgoU94hDfCF/SF7
iQHM7UruGG3du3TIYdKiT6GOiyUuvgleCRXL1ELE8D2xZTH55MxkO87O7CumP5CN
2+VVVOfI7Q1Co4LZxCgIWxllEwJ/sSa7Q7Q8UCPVTuOcz87KjkgHNDcSgMBWjgrA
VHLI1HNQJceWoAr/uAW/s3U4VxcONc8iXdGkjljBnTGZrI6m+GLSeo2RnFuu6Kjs
NpMrF/cxQzmMvriFZt+TpjiXaFs7uBZqbMuXFbZWJ6k+JDnRiovUWqaC171RXVTq
LSeEXt4mQf8S1DmjjkCMI0PxKpzXNuBUQpXdqNX3jLWz0IUI5LydgcR8W+vbthd+
FQMbNensaygRT7VpW42LeBAOC4JKCZZkeJoU7a+yw4Aj7uqnV5suzVwS72GdEg1Y
VE3yFCKYI/VKwOazT+7LTbv5MaXDxWPS/SYb/8wsM1ruw/hVThsMGvjBZLX7lRgd
1bf9v/VBux2Ur7mtLCRWV4GoZ/GwBVJtOayvT7ZNUugYsFjEM/w2ihMepc8EjW7A
YGGZhFgtbOUGfu2Roo/cqu4O0pI0ZxInFpVbQr9KMa0N8LLaz8Tif00mG90Pb9yV
dTNR0OBOK+xFISFM47PrB7g7pMJHABkVztLL8Cw8rKX8A7N+kvZl2y1Z1R84itMt
P0fYxwHYZkkthDWUJ5rKD43rqSYo2p74KRUgwFJxAppfvCIgaoOGFViZnV2yye/X
e7cDk6e1/3ZQaEyooKBcWX3plnexEoZ2ZsU4qMm5UVgMJk4xB7JFxUU4KG+olOAq
tIuk8bZjNpxuGjdzL0QYk3HwlGfZXnkXsJ1vQ5A2q7eHknHxpz6E37o8fOh/e2pd
DabCUXf1G0jiwp0VV/XCT390aQDF6IO//3Oaq4IhAAwh2wtEcvRtkXE+NanMnWB7
olzLN4RkO6jRr5yETtgGqbXjpdTVYdDY2+Zos2uq4gLXvcQauP4gUjLm9Hpj44uu
nsetOP21dae5CLE7R1OFh8Q3FN6ZYmQs0Ou2BzU4bPSZ4oKtuOTmb434+cGrkFUm
suFzW3IM75bVuNz2h61ksOZQ+stWd1ufIKTg9UhnHIR47GDfIgem71rFq4ofXwn7
t3Ndv3e0pYVamq5AwyBYaQnduDy2Y+VCrjtHO5F7mXe0AtkxI9rlxacfAmytTGG6
cMa51OzHfO9C7V81jK7RmSXtCGPg2SVHAW2tyWxLsmUszv9YiSbTObi/VSZH7ehC
6MkwuHXGL4lD70S6G/3giRc0ts2YloNz4IS7JylSMm7OI9apD+w0+VQy+op/QHxM
82aE8fO4S9L52L56p4ZGN+UpHz9HWHIRgpbLCM3cxR/U2OIT4dFcnfAkmro+HrTe
HLCKabN3cm6tfCeY/+8268jRmewIwOiniktLhuFYoyHNtmSTDOu0Z7a3j0FFZt5L
RVeV61kH2PCzxuFzBIucOs3/KFgQEpnPLNcd+uCeO1aEBHfZrovgDny9hUI5pHOB
xhYH0b5/i12k40W6G/9x/uH8pTr4ThhdAKEGBn4E0DxPH9RpXHe17HZkof8HIWFy
DQkwPO6pMKXVF9JdEKBGsWDVcUw/EDFlcO6FV5y64/P9tLNv/tzAohuQ7GaS5nLd
uSgaekdppK2mx1PR6d61N+UDwRseZp4JBxGOs/K+ONm06lgMf0nPgvGjNKjc/CMU
tmQSOVezUvmgWV2xkpa4c094AiKsYvgx9j/+8A4FJhv5DYRPzkL5YlRJ7OiVrax4
fVE1cZcWp2NvhCgUiyeU/lmjtuupqIEa10fYTZ1FDK0FKUoCBgKLoN649/Efz7xf
QbKtBP3SQ/6mRHOjYJ9VBuNYFe07r53U6FRXnXKta/Kmm4KBXooM591NNpa6r7j3
FVqKFf1sXjzKb/MbfWMYc/iTAbZt0JNCvai1CatiAl9UJZJ0e8Hgy5YB4xBYkM0R
WbKhqLP/vio311qhj+F44kMsjWG9ps+wQjzHyVSVl0ZbBHl2NZ2aVPsGIoCgMV/5
wS1y8Ibibw40ZpvXsRJxw00/jpdJ6gmXdXMLXuTxejIhrqjyD4WnVHOWcneRUmt1
mfvgPxtWgrc9TbVDI6KgWe5cly+v00RaW6kV29OUjQQb7qiYwj/YiJKfqGhZxKFJ
6vlVmLywxM5HwehFRbKzu4ZJpZ/XVVuRw1KuH+ZdctA6QuSW7MF/K6vAoQfrZvmz
3J//q1GLR1LVAG1i+5/emegFbS77DiKWGENtgTVn8dIorIn79wNGXnAKotLSgdVY
XWObQggt9f2ity2AoeEluvYsBih63COcY7Lnglazjw4RLJWabZIhqbKejeFaT0Ju
uxSA2OP8C+XtUqtOHaCqSuCm7AmbmBrHUgF5RHGqquuMq6EOA2ZAsZwAAP127RPl
thPQubBo0DwdmvlsDhkmJRyMJayskDSlQEogv/V6mMs1wR61i7behE9HmOgl2kuM
kvMlNSeilFAZX6Ahf4iBhLmlVLP1zbUj8GtMYCqyMATFMRmLoIGv8IZ6sn0Izq/0
0sYEeVGdwe6MQNrYuUrhi1ztb8bbnOrPnh0S3LDxPcOI6Znt6sNutUbgj0Mv8bl2
8Mp5vnEGg/2ZNBVvdZMV5voLpLesOSHJ5eGsudgMLcjMlXRgS/+Rwj3oBIkFnzIW
VCQi+3MbgR4gKEjZ+FUEXCgmccaJpYLsimJdJK1z+XdltV7vkJl525hKiTTisJwL
yuM7rMrk2SdTwPRRXMjAxZGtgMgRFZY2a8IPHDl4UW1R1wzwDZ9DMVw25e3mH5dG
/O6iXX2wznwnjuZ/zkzXw93mMNKETldpQpKQEGFSLv8jh8tgOq+/xKQOpzOh+7k8
YNsjGyRbFkS9YvwN31V75VIdy/IfMkQVtGD8be9Z+zQ7pO4xkTDVMp8FKMRxFToC
oWXEm8HTrK5+yp3cwcr6+aOO9t+xJ1cf3kGXiy5EkSpsAr89UcaUGgnEV8+DRkoZ
TacO9VTL4Pqj4ey3wKYa1l/rD8w5o9Z3u+XERf7kpwkEPb1QgCXXlygzsEqsCiUl
ufzfKRPyqgWTHa21/g2k9/IftO7GWmjgGiLjWW48bPFICWnKj+igwotMfhwuqT/p
e31Ym/llKwBah1zUuB33xMW5Zy6ULEH5Bif9LyhPj+uScVxO179eXGjF50ARZA/B
JIsdxgwgBzKsDx8MMylMlhJk6uXlR9hfHO5AZP272wLjSMKkImVfMt93YvbuXLZJ
3mMiLX7sLIQBE38uooiQ4SeRjoWnt9p2VX1rmWRU6ifyCXP+/KBinAcA8sKGY+k0
qGS56ADtPjka9u9KoeYxDL2vEfu0owJCaZG0OfIV/GtYDWZqU2SIiOR61As8/GKu
CuKF5INMxG+CPzRhKOJP3IKwuHw+oqefmZjywS2DXbiPMaCDemgNr8vV8R3W3pz6
kWQFqmgkdniDPZElpBMLNKc9Q5rlzLRWHyqtvCQuZxEeuGGzHA0yF0yHGOI7Nz3n
lYtlCUveZA/vk8ju/sYL6rp3J13m47XR8Juk5+bfwAF9xTSFtuj07g9G7pCB4P5L
bbwub+nhs7HbykTfZR1kLI9sdQM8vgDwk2jnd7Cc0aion7G/yQiZ0eeSUelEjGmY
c7e+ulv/hKZLoa33B3KQMOFoglOuaS1So0e8iqw+v1Fy9AOnwJOWgdY3YTWO79EI
EK+5PlXnOXok2SnITs0zSW0HhukEHTeL7KRfixKfGnvVee4XOtVfh+ncFWP2DFiE
4iX79275tF9vDe2wMUtsMmY3YM++YfcafWziIgZGB8Dl6La4ue/eWdyrnreOeKbZ
kpCTqJIFK8V1di1anKEau18Hv438eM72SacDqsjNZUpkCA9NtjpHkNf0sezuKAuX
I6MeDldOJA2z/gC7zVbBfDpFb7YTot3tczJWNjD7Eku9pwPwJmLypDZb9SxsbDi5
yYPhm4mHWsWgbFOSuE6aP54Nd4h7q9704wZfjlTqzNih2OF7Kv6AHnY94uQ35HB3
JjFXzUOJPQY8pbNUMypsZpY/WtfwvU428kKh6FIIJVnRt09zeEUii/oFurzzRlQx
Pw/942865tqqFnP+qpeVyJFA+YDQiZuPEsKL4dCrj/hbZCepinIJo/xq0nbg0pq1
Dc2nXKkECgufk2//qhrSYeokjNrrckTUKhcBJkMlwlb5sMGYJ1GZtXmhdK5UD0zb
nbzB9QbsjyEIYJRrK09PekWkPCkH4AlcJ5Hd2Ev2jq0MC9jlZ0kkUWtsHIy+VWvy
Hbta8E0dp4shMIYv71ZGDuUktxRKR5hedMzsgFyBYdL1w7bQk/04p5AzFbWIHETr
QcRaIYefOfz6XdzOVRAy+NsvHDFynaTfBJLbq/cD7uaW5/+nS58a53aMOr71ZatK
HiwWhfDOi9RCOUp7+Z+We+SgRXvirwsGb3k0OWDPXvcMeKuFOSk0DxEn1JmA9zQI
QGWytEFTs9qjseSDrNQNnEn+2GXatLWLgcABiiiBblmSEaIuDgJgCpWpwvbSlf9e
y/pe4jkGJUAJQOwPrmb6zKR+Td232wu2b6V1gjMobiGSiKmrCUdXYJlyKh6jUYk6
g108vbK8YilbAVn3cqPNOTecVUJ8UW14hblxy40PdpU/IKioISwYqMyAA4OWM2Ft
/TsDIiSpL4oWBruXy6VmjJPtsg1pdH44LXLswDeIQ8vpAEcOKJRA1IHTW15bsiSX
epDWv6ClmpOc0zfWY64cNoccNwsiXx3MspWpXfSxXdnPeVR0fa5jwsCeLb4K2b/C
N9zVRi6oor4I+pN4eLzOYS1DDgbo2CO4h2LKGCfTQZpI/D0SqSdn+8vwinLbpEem
4ADPLFNv2K7UEMmmVTrCazlUTgbayUYeXayO+BaGu89fzlCN2CS4nKyMLHx2rY0X
u+pe9I8R6kmEoN7ay4nZmb+0uao+dObzMoPLe3w/e/Ny+Ykv/FPub0mE2FKKPghw
ZZZNuPkGPoEEa40Qb3r9nLA0lN/v6MH2FlpvQRKWooYTDPnCv2gkOPl/oYQVvTUm
InAHaMvUx17UZoAHF/LvEWxG8pp+tqsSWxPuaAxgs9q17XsRiLBnCJWsz8oUijfN
UKc3Q4chUZWniTvPQem6WsRB+xf+PzRs1BJSQueIPvHBL0yU9Rde3x3r5QSwpgPz
Ftq/uV3Fuc3fuVZRs2rgsaJnxgpNrGh96Gko529nDuA5rt5QlFXUmUXPVa9n7heO
bkONsdg7vCHQi2fozXmYx69Jk5ekceYUTSR9jbml9Dj+jQ87rXChXJCFTCBxJXsd
gRGrVuZL08tmc1+kxkkmzATuJK5EusgzDEQc7gi8J5OVh0X6XRDp/zL0w4ribL9r
y5fti3ySTwHLX3VirtecwJjiGHcNsERQWZMsnZTW15siz1kzsxdN5iXwzZM4N4UY
rH2La6KpefBjL+AYJpwLrtlbGfFvxe6qy5tCcUU7q+6kxWdw+sgWEqIZQ/nTWvUL
XpO19Y3PTgRhqbpWxkWiGPG7AFnvgBrAj0kcgUTJQ2zn6IUtpdAgYBbr1n5RFQ6I
Cx47v8NWea5dZBth6QU7CmXFOnvAU1AnKdOh48RGtDuy0rwAItxZH33uTf+D9jon
0Pv/x1mbB+TTA+gec945oZB8HXDbj9uckkF2V619Eqp8QRFREJ2JY2YkdXhlDf69
/jNl3akLV+mVt14VFNtxez5tVG8Rq9ZQ3bNnG2/jqGFUS46c3OZ3FiC2PE3pqhJj
86uc5vPCZSoZD0vOY7+zFXqhr3V6h/pGKYtNthtZz+Z/OQEQJ6vJnNKr/OeZFmVJ
+g/d+7ndxjiFZ/mLAiIMB6KSjieUr+ARfbLQCFZ76cEVz/E2I8khQjqrkOQfqp1V
5N8w7DQ8/5EIyacrTbDjhZ0Q/NOxD8FBdNgVfKK7T94Wrla31J89wA0dyDlG/H2o
92O26hsXDwWDAp8yEZy/toEmTvxjafc5pai3n+vwy1X0NkgFJQrSQM0tA7kt3jVb
zq69U9/kpLOEnCLFefI/QNwGjsPuhZ5dCdUlGMA0X6B/uDJEy+IcQs5V4QkyjKqK
0kIminOkZoYGHHM4hOKMRhYO+zv3g5z5Vuhqe9CWgDOPiFrAU2MePm0d+ddhOULz
kwcRVzag9v3pXXEayCen5eHAPi92Hqvxm2EDSirDgRi9a79xU9KXmQ0PMVeHH0g1
WljRZK1ZhdPoTu6Qr8PLapfTDrYJJpdKM3N9ZJueR7My0USQoURJZ9C3uhUktspi
NmJoq9JRaWMkEYlhzraOgfWy9Yf8ko+14mOc+JygjCU+7bDgCpKfWQJ1Kg8qaIF5
Raxwnzu+OAMqPfn9zPeAkO3QdPboXnOMEzROGSciZUW8lTLDw2bGFG+dg3j2CfId
a1LKD7V0iQkYNxi0xKOIPoigg+rzYRa9zS/Q0cuZ41PVODdOfwNSAfHAnuFM9YFZ
m01rRbsR1eWps9Jy7n6fy0ac+kR2ZOA8ziGIJDoqGj92VuXfm3Jv/pPxr3C4pGru
KuzJ+X8T924qZnS5gWkQzDzz5SIsNm+aJSCPYWZLu0CE6TwjdS+3thjL8ydcXSof
wBA0mqQOWwESr4RALz6+X+hE8rykV1oTbp8dmZIGdBq+k1yBJsV7nFQOH1Yh6e3f
135GkBo1Xx1RtGynGmVGA5+ZJjIIEG+VuFyOWTM/yd+cbOZbbpmkL+0ydhVR+oeH
KnVKgPc1icYFzfKAJlCqZCJ8t/KGVc1WciM8G6JE9b2jfkvY1C+iNwV3ZeeGKHwP
rSu4oIG4lOklkKk0k84Dsf5vHr4cssiwEHqpq3RtS9siQEcykTIYKGn0txYKYSYH
PiNydg5bpv9KRO5orHlLCTxqZ8bU6bOpZOfm0BEHff+uF1ut9rnfPfaCcdWu8DlC
Fgs2OATyogN59ycW+3OUCzC0i+gqoxspJneGGy8KLm8C8VokleC2r/akJFMfRzs8
mRtcifayHUtoqGESIIWLkvMrBxzVlPcmWbc169qvktfwKya6gNPXzWJoI+Z2XX6F
4bIYTYwd++GirIS644fcjnbtEsEOa/5AwBQr6tBfif6y0aM5jk4ephbebzpDMeeJ
yRQj3n5FjT0yYi2vBMF/J7fZ/BhoNIexqtM+nyhU0KpphEmpO3ub2G8He06n2FX2
K+pHb1wp7X3LK1PzVcuEkBkvkFqBJy/1igFcUs9AHAC+1cV2e7AAkv090P11qH6V
a3MIXaSgUVOTcLqRFTs0ZB+uq6Or8fbtI5S9p9zng2LN6wr3WBE0MuAxcBchOqZX
HOgzhFaIu8nH34IUw7ZF326rbifoMuFWulAXO/JkzTkXJ8M+64Bn4y4RVJ/xhLmO
BWtUJLWmWSnUmbgAX9/uu5qHuwktIx4zJkYVtZAhS5Fa8TpE5bgaSUswvbKLV76t
8+o0VpcCUPGui7iCsT96krnDV7aB4k/489iVL5K6SDVPSHhjSfAwyUt+Qu2ddvQU
DdyqiSCjsHZGQHfUU37CzeJOqIXWy+IH3SLxldIhduuOf+Do5JMIYsUAmtzxGZAP
ELyDWA6atBkfCyp4kpJsHZG0AhPlH4Qk98iBeaaTvw0YZEZPYA2igVvoq0Fa2re2
rACQEXTWfSPrEVj1lkvJNEp4GHB2IWCbNsjfKMXZYnAn0RLkzS+Zscy210aq+D5m
u1ro2ci93ToX5J4RYYRt96zkWiqeVECcm3M/yXdbRwSnpN8AMSH0nNPuKkXAL/uj
0F9ikn/gIhVQaKOQUggcG9+OP7F5IJsDQD6getnhbe6ZXp5RSJkAD1EYPu3aVLKZ
vfvwoZ+X1G+dkPTAmYOE7/U8admO82ftyl/IHKktlLOUcmbu1/vs94zb89q13s/2
1WCQokpSqbUBR00yNkjSE2Sms7uQaI0tHOJraswnGm+WSC9Bdg+GnGNortXkWuFc
zGlMWGo6ECyxcL/jNxjc9HfDFQTD+Wjbaets9aFTPUXg1EsB65Erhy/w7chn8vQV
iHqJLA6qTpKI/ZrHRcZwLfW0ydTznHBHskNG1Gu0ykwuCtw9bD96+jc7inVqG467
IKdiCFBd8MmE+GLyaQAnD6guugwSQM4zvjwx/JnFY79iMxpxXPjM0ehD2wVQgrQI
i7Fs6Ygs3oeR9j9qmrpmCcUBiQT0Hq2BqBiD0nCRXvJpjEtj72INUnL++pTQCmrY
LYGRklja+73M4vv/v9mYQNG556RO/wQ7O7ZFr1HXCg2F7EtpQlHu5VdeEsrBFv80
uptzIIGG2LoOw30nfLdJOaGAYYnvZfY4Xqf1V5+W8zQygRE4oCGt+snkxLsKMJ2q
ZbzV6J6ZVZ5zneMeYQmZ5FvE8/ZLwsB1isgsuUWNOlK2iPmAhZVDY7KZRUsC0FCb
BpI7jDjX3XGfsyR+cP8iCN8djbOP92cviGzpV5Zh63qezr3v4bElK432iFA9GS/B
Ah+3onMkPHUBlcAYurke/WcAbpP5CQrVHSjOUif38Xt64XaldmF4xdN0GztCcdob
/VfP/eT/UbLYo4eU0HVE9YQP2IMWPqEQPoiUa35SRFNed4zZ39f0fKmfKNhVRpsE
IFPw6E4PysaJFMMob0jWUpw9tObDiBjiuqO26jFtwnqnZiZTD3r6ZUr4dZFDif4H
jpf7wWB9zpmwz7e/0SqyA46J9yiK5cE/38dloERxYjvHwB4Wff2K23m2aV7yQfCi
D/CR3Oe6+4uPw9uyHKo7+wNHmBWieE82CQx9OBJRlD6E7zIF7iVD56qt3y0YSVSh
ghkYdzccpMWH/DHD3QdqGjjwb6eueBXH7ds0dontyhLqiy1eVUH8RRFD6mIDiLKF
zfqxysoGITRcM0TG46Sl6axR8whEmqejMjfkUvPLHrw9t/P11vgUvVBQ9pjaeoa+
UgBeCQG+rvPSg2gaLGA2O5Jw2xiByhKwi2nJuG+kMGfT0+i5kFJAtNX2Tx3cvGM5
3U805o0U0IiY3J1KVBjWa+IPgbPC+Zu42UczzpNIHtSGMD2AWJR5P42FLN54sq8H
8CLeHbo9xTUmTsY8K9ttyTRJ6G99ejc1PX6Ds/lH1GjnN3y+XM/OScY7derqlZWV
pj0oHjzBGKfrXobf2KwNhDOJ+6p3bcsq7y6LiDzeHPoVrFScO61JjTutjN9U8v2O
y6EMU1yjIkoRSQ2cqWq+vnJEbQYRvgO91a9DnxeNL3F6QYZDieFmLaS/EoVEcfX1
XfPBqXOzHkEFPnaax3RbzNQEvyjLGz2Sh/gPb+c2D5NPwH5rL5+w2BJkmN0/s8xj
q4TAsf+jaN3R5aGQQ+j45zlzdyttkWcvGCP0TAMHPEGqelHUktDVwQgefDJMT0Hu
F1tAENyzUDm8D4gh30qb+Dz2UpdbkxqkJe2GvSOcZu82j7FXVGGYFa2qfJtLRhfi
KIlbqz8RTg08qTabvKAyqazbVyNcAN14F6O5ayadU7wcAnbMt2/L5zGfLP2DEsL2
D276lT1vdymIy1TvqhGHPXf1OI1mkOTEs23FPIaE/sIm0BARCQLEWT7Hzs+dgr7W
ibLS2fUFDuzDMytt4iD5EE8ysyO7jVKSEL00RsUJGyiobHm15jaWgktKs8lWcllc
s7HjBaKAEIghKg/d8CL24fd876G8k/8Ve80Mj3VXoEB9Rly/TAnJWnNsaJRMSdAt
mbAFjDlyCzHR+IMHQlFx4Zb4cr/8jjMkt+6Io9fZxN+M2vP1pBIZcchN0aY8d+PE
WjdJOx+v1sEZVHoLjsAgaQiYHfHuFffyrtZ829GWodAFdqHJG9vED5choznEfl1Z
12Gts4mycvd20p2gJBK7d0hUfVkXCAAc1Z0PuyT1F82eupMd3jTrGlFVFfPBrhIA
tXQFTv3r7tgTd4ns90d/2Hveu7UGnYOtvKvaMZ7+/tFeN6zBCnK1gTAFRR0QvbCm
MzcvJIFq9ZT4ArAM+tO3OiIe5CGsUV0gh4zUpRq17KUgDDo7pBaCcsymDkH9+RRu
Q4Tc0NbX4nQR5na+++U8XJHiZyUZZo5y7CJcARrL7p4fKwtsxfMEWYOQ6SAarylO
/8MtS8oj7vNSNM0+kdhfwErs8P3yRqfRuQzfdo79RodRpPhhFh3EKOqGOba4Euck
oWKqtISzdndvr1WDYn/tszDY20q1C2Ea0DgKbKQ8f7x9dFIKH1UOFWV24Pg8zyhY
6O97HI8ipbo4czr5afitZj4LhhAb9GI7AtjqNvskUd4M9dCpLh4dlnySkh8I06db
0W+nKyFQ1qME/TsY0JM13Vzm6ICnMHvG7J00tXa0atWL7Q5ZfIDeksgb0K2pt2XN
/45oj/SfZWDFQLn6LtJ2jHdsRzmetfcmKLxEqKoq51LQ3Gx+g2QkAWUS3BUI/e14
0zarIpsw4Z6AulkkCi48tF2rxucN/tcF4rgYUOr4rYxc74oFIyHtxFz09+ko6pbh
BZswRVR8A2rSmBk8h8xdTdDCSKt7MFNNzfkIObj842m9TP9HIpQ0E+/d4UHPLpWe
Nzx/d0jr89y7+A8MskfWpWlHhnqe8EzPrEqaYZEslVzaB/kvgNSm0Vuq5ZslRGGf
7e05av4l1Doo4Q8585UPSjR+jXBJbdW5VkANvufZfKa+R3uJINzsUh2B566fVB1z
wxK4wumKNZhtoIrnMyKPQxesDt41d12beJf4DeyZornQ8qlpsGPopLRzM2PA+If3
kaSnaq+sUD39upm+2Sy5xeM0c80Rc+hnYOBz8vtCrbWXFb7YsQ7eUE4CR0Tm3fEA
OqxpOHwI1O9FMwj/vQ7ZOY98bKn5tnIx37ZX2/0lWBT5jzItRaR7bzXok3076Zm7
rhLo73Enbs56E4wCPzh4YzLUtOtAB0eyjXr6fO59wB4e2TnArPS/LJOf0dvOU7UM
pX40LT2J+g2HO2ojYK+cMV3A30f8zm81HbcfAol6K/gzWWUVLWB1U3B0PpLMT/Cx
seXRuCfrznqbiE8N7o7Zy5JBVbsVkUvlnaPOnzUqHsQjbZUu77ycquDqDO2183YW
Ytus8Uywekho4FnKhhj4bFfHVhFJRwlEslxM5J8n2pqhMfMtVtjI0cU0Zx4uFPH4
QQh9KDvei0idDMdKmnPV4bvZpClEdw79gwNRyN/oEno/iJwCTAG+OTnrSwwKHQCf
tB/KfYceV4isvLgp6w/RqQEfaAAfA41cEpNqDoglN7tFPNu4a3nWbEMAJr/YVMne
BSxzbmLMgxDJUpTrZ4vYodDuKZyuT1vp7ABEM+n3sSE+q1UVbp109EfkrSh6MWoH
anhN9ClrFwiOKLQKRlrHLqdgRCtJTgioaDJ5QSIzCpckRZtusxV19H8wi3yX3xHY
P2njyLNFMCnaTgcy+5TBBn4dE2gPBL/dkwg+cTm0SExL3d3S0KzPHQ5a1/gpk8q/
axRPjH5+IrUcPMhi0G9RbVXasvsml9sevtpEs5cefWhuaKy8MnHesquIoaKDlNwA
Ty61AhFsD1UY14v15aWnDI0W8eQMk3qE1X2CayfzgAjJ6LloFBvx/5zMr2E61e/d
L8meQD4/5xXb6KvJgFJ36yKx6mLPtgC2lqSSP4E8vScyG4++KY8dxHW7wWYCFzAE
0dAsUm+u139Y4FQuaM5Ez5HtA2jU3NXWSH/oAae/0K5aqE6z9dXZdzpOdNreH08T
TJ4MX0hpjAuHq1hIZHrFMqfS3gznC0kXOqLmopYjJlPmwHkNjPtrnZzeZdWaVsX8
nxGqxrFvXyvTfUrkLmlhXjhUiSFQQTE1Qr5VjW9gIgDJgJYwddosRf3xolhcjEaG
+ILtVeuu3u1fGTVxOT1plq7dxncHkBk1AgzRR6Jcxqt3mf2gGCDTwa/BIX3P5MiR
otSvluOSakifk2NAcQULRGRUe4AXsWwakEMz9mDS1cXlhkrb4km0eIABnlwiFYNQ
e88S5zWuobsetUznEMUNfYUb6B9yu+m1KfWMQQUSxaHd0eQMx8mDPIXh+fxPTqX7
CYtqDp83mD2nGSOzUAKcSWVJ1sunJ4snpmd+BS2qsBevwfTw3JfyNpAUVl6niGVb
dTf2YWfx0nyU5khI8FU0/y6lOpvxaGg6Gx4NYN+tjpGnk0e7OXL0bnRpSCc8V6dO
5n2pq3oPbW7tj9/not21VTrqLt3PRrsY1jZ9zUkMUZhvLzajoWLudMVcabx5eEBz
sxC59Llzy+IieRqtQjMs/gCssXapQ4GMtNaTLkyknRNG9HQTq+aO5fi/wnuC7xaH
ixVmQW+AQfFD/Vv05Ug1UHGkrjS5QfZXcEzKMxgub8Q07svjo8ILeBBuyb5qJdxQ
YK62AaflmJlZPkocV8Xj6APOf/32zvsbU/6kQj0rM9Jho80ADjZ11ZLgzDBBG/kk
ws0sVxtYzs4OmIoI0Saf7rCDiy0lSzJPqzFEl4z1a9jeLbnsQGrr79MHxB9guZwv
EEnWVFPGgzv9NipJRRnD0no3+Mer/4JFl8Xea+RGnWAjHR84e+PKUHt7nC/8Q0po
raonoXol/M6YTmSzRD/lRr1U7ZpGapu9wkJrMb6xXNMdYQM0OZBjSjBViXhfD2JD
J35lE8UAB1CtBpURTZMkZ+nFC+4z0SaLlpZ5HS6lQJnV7p6brKQsMMinGC9SFT9X
9RikXcfxNyQoc7+QSGVOR2jPC5sMfqn2hs6C44cjhAeQigQJHHI9YiXf6Xa3VN/T
Ri6jp3qeBteV6gXxmiZmk4QsPFtEGqu7RB7IGOTnCIeSPvaE8jte3b7BslXZdJP6
Jc64EMTWcudjD9qKDECBw7SaMQP+2usHsEgu2rJJ1vYY5GTFVXZ2syNGux6acv1l
MV0CLVutk/SH7QfjoRQUT82ZRTyUoBY4icIR40vO56ZMaE5VZkPVSdmsZAuEJofE
g67D5arwooJtcnqHyiskv8P5mCR4a7CBgkTXo4rTgsz7rpiLXmRVtT3DyCsL3/iG
GQWAj6oeX3g8mELheCu+ApMZaEfbz3dM2pnpmw4udFr82Xu08mguM+W75k6fErIA
VFflEp3uta18JWgpEVbkArNeAB0yzu/sjLJTRtT5Ilo7Vw8oJRvelALs9HAcGmvC
Dnv1ThoMS5w8hy2VEyWh7X5tfza9cqSkzqJSwN368G316V8apEQ64xtXUY4V/RDn
EnenyB63cPp+fyP/f6gxL1txt0q2VOFkjY7+Lg1VjOdzubKty8MpELr2Bu+9YlFZ
kKNRQSyfy61V8UHfXB7KQOhQ42M/dsqaSR8wWZ3d/3xlK1Ppg/TD/UxxIsHcU9yC
Gaa0UrxBmGQwZZwUELG4gbID2u+Wn2Ha7te8t66lkjQ7wIro7NRebbNEMoOX91JW
VeWoI2KRq+pso6idyIUc9fp3hJBFrDB5kQiNlfnenlr3KaKdQLAUi8nNVdaMPjvU
TNVyRFxAa6NSQVmICNVzfDrYHI7AHCoRG06ODyLlY82bEjrK0KXNf03uabgC9Nuz
njrCAT1d5g/Jptj6ok8IW6mNUk5OUoqMKtDdtqTgQW+OC5JheILf1gjBQ58S2u1j
IKzclZ/whnyAdnOPqrR8AAF1yNh3FxHGM7+hgfdx9sMv7mC6hbA9iihBonGO+chu
aWFKpiGvl2I0Oq1L/gC6tyHqnMlyRlErAUL/+0K+u+Nw8mwdfSUehhAbftmp4gKH
WHc7/6IVJQngXWV0V7cgIV5q8ebdl9EVIe9wKh7Bvg/8fQ8aVhXcdmj1rP/mItyh
5JCbXzhofhawgCVFOVuu+NuV9SOnbzKlxkPGTjq1T0OlweM8NQTHujO2hR4tIQ/t
Sy8tXeEwO8Vc/zdlsYiU3szfbORbkwPDRtqdxAxwTIoQAZLvwiIpnq1tt3zqUKDL
leWIH3A8K1T1NIqaKO3iqmVArswR9ts+gUOqcPShA/bEKwbX5n8g7/XC3a9nWH6K
dhpF6PBN87W4Bn3xmNrDNOfIoAh/rL5DccbyiqewrMRYz3ccCGZizvlc6UTRYkOX
HaRG9wkZTGNb1GHfSlxq9JdbfSuP43EOoFCdjLij5uiS58ANBKBh5PNZi+Cn9AEk
75LnfkNl3LeIOOX253cIVfuC76fXEIiW1Wn3xHYfBEtDpdWOohnsJ0Pb5A+s7Sbn
5GKaR+9JvbPsjCdvdYZxmvzFHG7vtuy7PYt6B9Dl+vu53F7JUDQVnyGnPjTvycUo
sDgOgjeWrOGMbsr8vzGztCEmwQG8I1Gt5zdPF0OwxY4QACz4oY0Ep4e1H0t4lp/0
K7RY1Z1SsrnLdzfc4GhydvtiVANkfm5SMwPzHyCEDyhwqSDrRKkGdaYSTTbFC7pl
QT8tC91MMFWW1j42cwCxi2yUijdTHGa1aPKxLtGiBZ8jOcwbCWINNkebeeuyOrgi
Su0PgGSPo2BDVqcvyL3+1pZyxFrXupFMNimscDwcaMhMVT0RNex7AiYkMM0vrQse
hx1p0kxh1EP9iFEUqK6gaUwfZaL6dwkEXyIbtHtbqx6sfl4mD8E4gS1C71SqEXbp
jsfIwYauWLgmTYWZ8UHvtOU4KybZ4MnHzn9CJOIvWogpN+Bcs1YHuKNjjmpNu+Ko
d/w1qxO0CURR8lQvnD9fypGeAlGFqtgkmpyqc9jeRpc+cl/YqHK163MikjPyHZ3O
QZowSOLR5kNtvdz+l7Z/Rn0vs68sx6s4L0tjvvO81BQY79uOR1Rw+vQ/n3ShBK/b
0ByLf/N712eok2epKWZyhrD+xJh3qeUasWqf2r1i5wieoYBbOXgwWVF8q3Z6SxeF
C4oRqeX7JnANd0wNsM98EqOStr0x84UY4meXjTWjJbZ6zDZzWT5IiLeGPh9h0EoZ
/1CnvMpND6ATNhDR7NIcFXBLODyWJmKSK/QdhM5XnuKys+I4I4gE/JwCBcp8jjAs
fVkLBmLKU7JeMgNLhhUOE1Ac/we8a/wdD+daTlOUW2vEgDy0EVyDSQaQrL11fAec
/QXfWNZlFHdUPsEVaB1JXlCVCh5ufViwDtQZXBGgcvJzUEDK2ol32Ln/Ed2j6oYp
4NFkKwpWMtmwBj5E2+6LdkZY5TGVoDNsGlbeRIFpP5W28nsEhfp+gng5OznigjyY
Sx1s5/yhwbSjmfsgIKJShZ6YEHigCxzMjYIVwwZSfaJ/XCMuG2rM5ALZkh1w1vLA
DGBhvYC9Dq88DTNsa0MRdEc1HMrgijhAiHdYLhuNIbM1kw9/s69finUMCvCXMdCf
0YFBEuvuRW6JkgsJjRyHyowzWnzFsDoqohiMkpSs5LtaNj1yniumJpbRO/1KW96p
aa9OZSvax2W5D/8pSLDCswYp229x0BlL10L1uAqPDLXZ5mw6oMT1YLlnjWO96sbo
0CWCsNcH+cdkj9ChvGkj9fFM+sqfDJXCgrmiXo9ya4MsRI9DOCgkvWpt2KkBE2lh
ZPmnUqrMt+N3OjShMB5ZE8Osbld8rmuHbdfSET7GGA9TZIsfGc/Wwqgo/ui/J39n
V+YZKMXEnxB+1Ybl3l9F+q1qDLit3swiVRUi9NIfj4rkcUBDyhbjtGUJnTVzkNng
TfK+b7Y1elXnaXIPz6KwduCn9mru2eDiL+FbY9DbhOy5eBuDqDn4ic9fDv/nj7XL
gUvDUBR0X2WrSWRvZ7eXJ86ZqBJMKxi33L8fmSa5VntFgyaBoYyz53eoAD5KRjOE
ydeO7DVagCDsmB9ahqriKB2HCnSWd7RK/B/Ym60WtrCFh/6m0DufKR1GysflIC/c
KnzQhCnkDLf1jImgeYw57VfGA5mHorX6ykIGZYXJPlpGNFIz8cmSrTTj5P1mm+53
4wHFkpHd6XVMUs7R8WPk4BWetutHcjF5xG2keu8pkOl7WHXp+DovY5tuldKLSWPO
4+OLafEzKXZppvGQUyOk6d6j1QSEHML6aWi1CIVtde5RwIv30aNsZRU6oFwFBj1T
SdvuvtZEPbJiIimqs85MaoMaOckXzlTl568/eFGL61a+nntQ+MzQYKTxv/aAo7YV
j/hTquPZmngd+bIflaXDGIiwp4KlbuCgH1OhIeX6T4xS/lFJ0PoSfzIzr4Cm64dV
RugBCVDqfTQz7yLhWDwCRDQs2cC3NzJppo21RE618AlvNWQhf29sf36o2FfSbZ9T
9kUlS0wFztMkOqZ7r1Em6DdyhpHXT0tqA5ZJ5IFp8pzcrGZ0yJDsEVlyz+1lAsd/
O2i1NjzYDoEuPn0ckRfVScrvmKY4tzYMowYQGdgIAw+6AI/qPe2oS6fL0UbXMvkp
nlcrlqzlRNqSvjsz5DzWhWHR4pMfvrCi8TTcYoLSOyJUzyUDP4mtUtyYPpkvG/gV
ZsRFzjCAZ+sstZXuQxaUMPR9QKtIZ2PmYwtd6rr6Q5xbG1MMnPKsdARKQd+WIwAx
GMjtOp5Mw1nfTaAn396m5idzfYm20sER8V2EbS1GVoPF1lluG/Y4DZ3swjgLyACm
NP3PF34r36ijy5Hpuc6xjc8ZdwRNxYWQgW4w9VZJovgXppkdDHD5v2XC/+TrmBdd
AiR/r+leKQXs1by+w99PBGlttR4LHLmN7WcUIuttbl80oaZ87ciEZtAyIS7Pf2RK
V+cxN49wn4OkTczAWFnRXxUKAxxfVnWpa+stOcxqY+D1yHGuzMTfKmh9ACO5OUx9
FoyOdQmekTJnc0Z96odOsdNsVqlWclAsDlW5WoM2M9l1uL0m41DoMx2wa1GV3gLw
OWHNOGbqEOiUIYMmKQCdU18Gjqy1ulDXNL11mjONjnpLvpIBQMMjeL+IX+snCH7n
sMUDcRzZ8e8KXzS2QmrqfCWEiEBG+RpFdHv8DliADoqSy4srja1eh2AG8p6NZLg0
Wf6RVdanG2cVzoUj7XTH4IOY/Xv2MNw4BG6Gg3cJlwkNeFHDUeUOSNv9o3Pn1V3W
nBIgg125wZMWVySMmbJBF6lUUeRzkebj0ofKnajj2q0JD2AgpgC/+igJQHvOhfv2
BdA/bHYcvcm4eyIwjXB5B1CEMqWeU7/2R7NmrwIVMzs4ul55fbMagmfugr3fAji4
sSglnTkKpoXtSb3sR2KbjtXDTDdrrQU2opjX4pCnOdU4NMOPZ96rRMxGxN0SYJYS
kX7NbnQtnMHgpRjIaomiUdFtujY19oG30I8vVBAWMDgaNe9YT2giuVG4GbQTYmAP
33KKmhg5r76pR9Ooi6gGOK4TQ2xQBbAsL8KyXR1G08czVfphE6xXJIqiZiA8GLd5
+Ssqdk/okHx3l53j+0OQnucqU2jhj1lcCFPGGWQouDayhfi7gDkgTuxlJU6TIK4A
GVC8bj6BXFr0UWYmf0iPtwQ4ihFUj1j8mQ93OTfeK5Hz2opG5JnCAfK87CL5g6Ta
99cThH40XUW1p1J9xe9yNQ4uP4XpkkgMnHhHQOvryxWr+XNw6eKzISwBeSw07Sko
TWDZ5GIjREzBQ2XuDzm4gP0TkGEWQONHuPhDIditjfZSBL17aDP/ewLxOTcjiNBk
uxiLXY9V3IOOgoTBhnZ92PIeW6OPNNjS2DdFN6v51WDH2mkaPjvE8PwocoBg3/U1
V5yVHLOuyASidywIFdYo0uHpkg9knI+leJwrIREzXJKr15MNmPbKh82aDUykhmyE
WsUftxSlUy/TMpLfSaw2lmfWq4H7e2WTX6nqkPVpjSB090zl+4j6UmMdJXAmUtyU
9EiG2TOgoCj9yVyBMzrtuoj8W1EnUUZtoO41r5YWTI8fyVeCDPb+wCmt176UUyG+
Dk8srxIzt86UsU9GzT2PNFuDPd6hRbU0INhTHUeoZYoZQOsl45JwEuMITe9dENHe
tkokhsk+MNzU/F+aoUKG7UC8n9y7KSsRYqDYupg1eB1WAUM7DKkVc8kLJnGaLDBq
24p2hxjyzjUvBSBjSxZWZEWDJHjMRONAFvOQUxuhSv0Dw7y0VzJDoL6EYp0QlTxP
+mUrdfE2WHVs/C4klMm1slmeLy8cJW+Sy7t3qypMsCrR3uLg4uiKDJ1haoty/WCp
C04NVwie3s504Dl1DDtWIz+817Xpv9HsYhG/Oe7etCNYfiCBrvKQrVD47G0Nq417
IHIzhoR4hvzpPFcSDGiI9Q6BEcDVl91BqfSGmuPNoWgf5vcuAHXeMHbuj5Jgq+yg
aUEKaS2JmTND8BuXNgYuwPwpWlOoPvODo+/WaONwvuymVcVU2iIIRGvjxV/DRr7E
jH1Hnqjuzpq5nFnWpOPIPvMoSAR+yrBZo8zAd/qG9x83VKxCwayiNxjaSx7VzJH6
K1SOrCZ/KlYybd4F3XjVgJOrE3Fa/r+ojSqa7Dch+bvU975qXHmWxtgBKz6CziQm
nhXvB8tIVidVpYUe4somPJHFqQDc6mdP9xo8jEIbq/cnvSsjrr552FSfX6xiaCIj
QyL+Y+Xg2xLnm0PGjDLXL4cbm8OgTl6Yv8HstplyiIJZNwUyvA5wO3xhWyVfyHzT
Ns7Ut72tgUkG0j6DDZ8PipQyIcajdpMQR/PYOqnV9YdUGYiA3g03YHjC9F97HFMX
FcO5sG0NQbQ2JzvxC3U0bYHShbUEupXdrhSEoqqLOPFN4Mip5WMc3EYMlQFs3ljv
R2d502S8fG5aRgTMDHSqM27YQXrxcoSoPKcjfNvF2g6MMtJYZbRMF5JEZnbDiDE9
L77PM1D5RU7GlxX3+Oq+k7HmyV49gRpKBNs8za+PbZXFnk4SCyQm3vv7qbKRKC7L
LvtOzJYOuZksk/enw3soYQbkO8OxuF874ifN59Lj+17nHXlIF/XtcX6j/xg6PazX
MTfuQ4bk5NNF1h7uoCEiLs/5+zfAugGekgudyXBLMTfMyYL+iUo+ulBJeZJt+b9j
Edhx4mNcVYkgmgAXbRK17uU4FLjSWPb130JqN3xWmOouWD8uToUHssZgSoMuBvSd
ZiG8q41f2mZGe4tLVQ52HExCNQh70kFJYTFVrr+XgB26XCXJZxpVHrDjEfsO/flO
Bp9nlR/dyi0Y7dV26fKUsvi0fVAdU50zajImvDi1uHMlHoz1Inhdbuqo34s+X6y6
FuL/lVo+VAf2f8ANupVqMrFrgRzbmoa2LAS5Fz0dsYw+gCVH2XNZMmfVZ44+oA1B
qDXOcO9j1diE2Sg8yswnuhO6cyRSJRL+roGF5sEzqjr51DhEbOx26mgJeqvW1lgz
tdeUz5UR7sq12LvOKOx2AxV2RtXC/llUmKnFPDx5pSo55HnbTt6kjRtBBtFJO0rf
U2zfBhrgMTBNtDqIFik5h4j60vOqXSfV2oVColHD3VwXLEEicfqozNVf3IqrdWTN
KSKpo/qqk7V98bifnVnaJT/7M9DKnXPq5RwkTcBOebPs+/0ON7vqOBJhhuquXlDM
cKsoaOJWFg07W88xNpXtINHQPCHw0JxrhI6BECJejvmNn6muPbW99vgX2OHZHhFo
30gICatZ6yBqPN9XdLkFJZ2RTDchfTCzvN1tgyq+0GjzHI0RspUpToU385G5B2Fk
LzoOjKwvKWgiQEyn/fUkoPGGtND+ONkYPOu7KVAy2KzxQalCTfW3WBjH0N1pf1cs
kzfsq+jUEC20YCya8ZnIYPwrZ/z8w1uA0qvNgfK6A9KdfCAip0mGOFN/W3/yQ+Fq
FNsOCy0mIgLtE+S2GOeZTEhi48bInbyfhQA4u2CD8KcqTiXy94V0gck0t+opUioT
ft3PoCz1vw38KPAGO+vQTT2fV9v8P7SbsfH26ljjOFjGFTNwh8hcelNnaWoYhSzx
GJGbcGsAxSuRZdBoipMXLH29qrnOWqRefuHTAq6kuOB4EfsLhxMplcH2lnI/Nzg9
Ds/xi1o/5r/yxZaTJ9sKv8malJSt2MjZDc49tVEooP2kzu/+WsBkqQ9bR9bnYuJu
qTjladeA+c3eou5jmnyF9oNAKfwlOhlKViBX2LRY6CmkQshRDNmfvPfaZReHa93d
gLyP52VYTlIq3kf7mZYtYWIYiV5lc9xH98X4CpoUXDK21JP8QBs4F1NKV1I7QF8h
ilZxTmQHQjT5g9J1daSXsBHM+XNOeqZrYsmBUcHrSJY52dwg5vW02ODeu0Vbz4+D
yyelAXTZKvrdPcwIk2zx4tCqlruzx/fwcA5aUFumWNT9Gbsawh5HZCB2QH8cLc+N
4DL4FdSDvL2JVFhMAPprFbaNBEk//efhR76uN1r2mHojZmvndrDoJVJ9oXH+RO8W
yNgKGeOrEoqbbl05UQl23RVDIwlEjwnIIjg+LYiuF/7izlGOPy3oUPtI/Z+Q8pmg
GvrlYMaki7rGnYipgfxl5vS2KfFI0yA/M+zQdxjALuT5Bs3TQZvp1cwHX++YhvwY
dQ/3SQTxN4qZz1d5VSnIlghKDTIWn+fobKMKk51eLW1ZMZ9cF5hARu1dLooaVmoP
NB/1HME2MjcG7Xq93VjkKuzRwhtpJaQtvHl4KR4CvedoiVbjuyVWSX5AQP0TifEi
LqI72tAVOm0/uotuWgMEvbQ0JIojTTMjfYEbfuHG8TAYY7F/9Re77l1D8qy1u3TL
zc4XSM6ac3hVUEDkGlz89wT6W9+FIUGGz3pvWPs4/WuVUsPXIQrzhbAsYkJYRRUU
Wc/D/cMgyAmcys8tdD8t6D+0mzdHX9EjdggBv9fZth5SIe68ttdrJ8DV6aDUGkEo
pa3t3QN1z5zEq0s4vWbDXeFT1g49vu1ttM+9D1LPPjpjJ+kHkwVD1Mh8lFUCHIKV
66z2lIIeiv0rgVSErNNtUFeXkqRZ4hDkbVaXxN/aUiC83fwMqTbAD8gzRdpYcqIa
1axmcrc8h8RzMUgena15HKr/CfYbEbzmSRagtDJoeRaGpTegk+DCbIPxxCZhO9y6
N81NOmGHXJTAGf+9eLEK0HiSqqbCFSEbslYqElZrd1pvVDr99pgv2MJa3fXPT1Bz
H3OnrEf7ba2KAtE133pywlH4lTDha45z8XIVPUzA5AFtP4nBqlLywdB5mH1tJB4N
Fu/SwXM6BWlVa9QPzzwyoSFC3mRHmN9WRNR2Q06JjFdztIRN4mrwyu6bP8bWIuzr
3OoApEiWfOIV3SfXJMHwGDM0eERtuvv+2W8pKDnujMYy0mlBaeOtpoMHPLHtf1HV
cAEfP/BeQnOgso3lzYgnSPxKagzQXSiuHUoHg8I8lCe0JxHwInYPWPYDh2N9rxP7
5C9ShVitg1mQ8Xk9ye2YrlyRlFsIfYqwzXxqiKvGwc8oMeiBdGoym7EqjRuRQvk6
0OFnvZUj7i+HBhhPDAtzLXgcQEPUyEn2vyScckGQM+uPxGyd5ldN3P+o+8NDkB7L
c+5qF81i6f5MQ8lhOHnOtccazplgIBtt4ZXKbyxljBc6Vd+jFuKr76ILaVMMAiBC
Z4r26e80U22gxbTRej6DBKXccnCFrEG7B9gGZ7WEeK3oBHUqQTpHVK9noR223Ntu
4e4hUCh1pcbKS49R6vS+AxNmJoRamqb/lpRFar4ya/cCqqYKY1g0cjVlfMmOyaq7
iZ0Th+R28zZ3oXK/3gBwtnWI98ElG1a7g9Bo0EJmMSq30FaCo4At01lDQl5YooNn
JQu9Y0kNwawxxkSo3yi7aL4/7wAvgqvPZRHIrAXKaaaCfKWW2T/TwSywrtHpVqjs
hJ/oItX/qF3wVqyiaKpiPLPv903aFwijhcJxu/Yfvdw1/YOIwfieKUiOwgx54dB/
zLuCl3DLWsZwUWizxm6PdsY88QUwX1E9r5SZ0CMPkYtwpk0HnxnWln0hsNqpP2an
S0A5DNYDtWu6q8ux4s0dGbiFFxThf7N2gfDS0cUYFhiB/aHps+oL2LvGN5NIz0nK
9Vw2TEM6oUbfk9D3AlSduXv0fRid+r++92/T+v0akribvIVl58PACO4Zx1eGfnto
72ZMXUwISxZM+t8+923MiuBZ3zixMIysun93bIpqxGktlcgMB4jDhOEACxecMpnl
kecjp7A9TrKNR8SCQXXYZ6nqO3m8NSQ5zWcGl+j+KHy6siUyXTv6GaIwHnUQcreo
4x70xLRel3gGvCbwN1DsG1j1byVonPkzgvXUtTcMeT6mY3biTf38wuBjsDkwFObj
NPxdKuFpag2hRYpcsebozRVnyp2vpWX1X/qRyhh5q3FpYOYORWc5BjSHzp2Ncf9E
fG2T9AsCz7wOHJgPCkZupN61tJPIXoVRDF2gnz2AvuKx2TYDlkjIsgOJuE5ItIUk
5t8ZKUg7FKShqmdfMGS6d6Ih1EK0AF1YotsrjOMalqCB5yfwkTpX2galTS/2Rvjx
i3OZGfHlu0JDmslpbqbRfPvvwLB3FNsX5p9cggNUTSWIVxvuy9lx6FzNxzqx4eXC
FUXcsV7Zuc0ENh4g5rrZ2IEcui6v+hm6vNbg9XwUhnlYDyM/1G2RofrOkgdkj8M5
wsjrwTR9CF4pjU8BVGD+g2J518rP0otDwb3NoQghS/XB4T80VfpUypiSnFLhUn2J
//kJTmO1lCet21jykeCHxXFAAXxcWeSrjoXwiOfDT2a2xL9HG0zkAn4cnoT6WWdx
pCVS4h1iCbFm/5Qu0dQzZZlnrNE7jDFgoetswPeCfLXP3Nx542yfYP/3NjaVsi0f
7Xg86Rab9eaE9LmxF0Nn6cLzh3Lqd1sbpyusj87uejY/3ogI06UOMzwT+osSp7qs
jitKWlqnem5qaUXVmB1i5u7hV7yJJCXBRQ6RatOy3sMhJJ9w+xfBe7CcugStyWlN
lRRnH+VSnJe9OMOv/ommZQdDyh11N1cLK9kx4Q5iWx8ykYh51+IO9CZcULEzKQft
ngoakhxyJLcTNc41FuPVs0uek7i3ZC0xVp0K0Jhaqj/j5OwSiD3L6r4EMGqEb4Zv
4YyoYt1HmyHZlyS5xvul4C3ZwucJrUHgISPWjjk2b4DL9FYpp0i+j+VueZl4ph1U
6d1JUa9WOhmRcteLCghU9cPVDoIgA48JqrWCfkboo5lzrSh7LoEPc5z8QU+HcanC
V4MXdChSudNWrq/6ijJrppmuQZm5Bzmy8oXwqdh4Z8i3zWSQqxX2lXgz+wiKdwBq
fAzLMIWhKdSO1LrhYmFWf5djmjELzo3tGJt0E2Uoy+EYecm9a3upOE+RlNLbkBU9
GrfJ4Qo1iZVs0x4Kyd1OmrZvqet0+2soGZhfhxEGnCKgJLJ5zG1vvzQcxlj4MdfV
cMqD+dIWKVh2z3Ammi7x/KJczMhrZCbMwMm0GpOghmMilkq1b1sbJG+Y4TUP+GXb
PbF0XokIAj4kL35zoKGy5g3w/FuuPTmivNuCeGamNyG+isSrR6A1VdM/cwWADx8z
oZrUYKdq/e/5iwFQwIsapj/o7nYPCIMEAH6IxcCtXPZnY4ffJ9rJ7m9FyKL0wprb
EnaMQdafQNoEwBnoA9NCyakQ4wAIjMiAs/q/1aVpKaQwj7FKnDGYWKoiiX9unJFo
AQPZ9/8IpsxIC80R8KrKb9wRdQGeLNLwoc3Zfmqt4/Egrpm0LmdsOizq1p7h9EPg
ny2pztqBM30n59uKHvN0H8Kq+MK37OKbONZK73fCUmmvGtSV+ksltV9oToEbQBjq
dgmVCLpfRgfKUbx2cSKgsVsQ7+4Gvm+Zz9NWGCg9QoBDduDq2jxjWJSyWQiHtFuD
u4iByfbzkyhmWKdtLC0L5Uj++3VUvg0HDDuO2FxTCE+YWlShv2m6EDm0ORgEG8dI
/7zF3th/sUIDDH1mtAreQeqamPQJWwTay1EhAwtZDdkivrNOnhgFyb9lMquqVO9k
68tDel/8X3IYTtPgV0538nWvKzDAN6/PJuDrn3PUpb3EP9v9bmk29WyCQusRrUdF
AOKuicTVfvneLOun6p6ySFnoJZFo5AX+Vd01JU3oh5ucoZ971SWz+HGl4je41cuB
KXe6jzexzJBupzsp/Hw5OTa/PwxASJwvjBlUDteHFvT+cJgqEkg+nj7vfDY/SmfX
7Gn/RuIeka7tjyjWAeuXpAeVDQrXKizkvfWBDptLA5y8K7FhciBuUTK6HYTIqf/R
eMXhNK7Wk7vhmbNprL6NdxFvXyJKSnHDQO1jKokO4uOIJtIUPRIS517ntwYlGnRq
LLRQX4kWh2dqXv/vklrXTWGmfYwWdY86QDNkH5IXZyG2WIynY4rwOguUeRWiqqA1
8q/1haNo/jDavUuo+sQcgf/kXgcTfgmyFHHuY6wuRco7t8t/GaCtVm11uAb5R27a
KTjoYNHeOcytlm4zwD3kBc0MMRJl2D+sEYKUyKBeUFTT/h0KnILHhkgnWcmqz45q
CL0ChSxqbFtyyU5p6GMREItzEYlZ5+AhS7kIa6YTXwrlnvFErm1GlTa/BsU3Bs77
y+jOL37Xfst8oDQoyEyZWmRFMQ1eiaMycBOda/FP6X4ZVlDoTOnYK+u94yBmRTTj
yRTcmG4LYIl1AT+SJ0XMwc6gPcjYHayfCr/IYm1KcYAq5p5Ryte0+ZDSgTVKGiLb
OsnQQCN48tPGeZhWT+g7yz62YR8dntX05ZBu7YUroCYjA472YB2UH78ojAtccYnu
Lc4An8X03czcsYGhMttnRtCSTEJ9ijVHiQGn3QKJCH9yqn1OyYERnkyWjTmX7mhG
8X+1Iv4KCqPh0NNazuJHSBdNOy17r4qpS1Kfyyd4KJVy/yLEevO6f41g/sfX81k6
5VZtj7i3toI43yKAsdQzdNf9Ge2ZsNJLoG1+Lbxyd24ZlAp8hNE8o8DfmD1bmvDC
P5QKtoNC+6YY6hMdDfE5oi536sfPuYNuqxRq1lv4nwHuVlxKwvLu1RTKK05Bjnmg
GywMJ7OauXWwXx+7POAaUaee66sGPzFsiTgpA7CKN74ShiJjSWV+aHMcXOnWs0Hz
buk8RROl4uF8r4wXNlkGWM6OC+axmEmHFdKfZdDOPLDkgdhSxlJjA2JoCG0BKjqT
Qm6PLwR1i9WipXpvLrDdTxpY0zEodFQrOR1ynBh5Az/PlMnk7r41RJLnv1iiuQXC
MW9RV0DlW0vqXEnYpGZNY2Oplwa9Co3Mk9gLjN5ZXtiEMrzqNIJclgCV3OKEyowg
BM73D/0EuL26D294x/CtdfMK/Wo4Jx+180BUrECyDx5+LTWwBny9DQ1m4uxrjvaD
EAFZ4qyCLyCa37i6v92tBFT8sEHcXwuf9H97LalLgvQ9yHXGeXnRzrrr2BgYUh8e
QQJtcOTWOzGF6aOWGDMjFV6qRiJ5pqM8jsj4fauPOp00ppvzYSPBb0m4cMUgf78X
Khc9w9QkOc9tfII9UlANO7EMHNrefS6ELc6lrfXxJR88lS7h4p7GIfeBV+HP9OP9
MZxtVu4Dh1V2OGS204ZZniCZOuaXQP9fv60Bo/JGVae4Qe0CSCgZaVCDdy0iNFi6
2YSjVZMCEDDG5dvKSpxEcTqcWXOso/CQ8Qcs27iMU8P/1pHz05HW3GGGtxjB1Oq9
w9ngWoQwymtjJDh1Tf5O7b7Wl4NEvFVDFnBVsHxulEMoy5e53jeGkRBaaKC9XmUf
P5V5zmmBFhaWtfSLM0SiKLlxmyMSynT0x/mKvRuGsLAExOTdAAhpEcQkDMdEfuTH
njxDoFQ7qloetrgsvmgjX9lSDNHIEt6S7676ox9aqXPWBAmDZZzlndGIvNJ3owMF
QMlM/l9CZqmlqKjTJKhedlBHd/J+SkDFIyXYE6/U0gbjto2eNmGJlXhH++4e6vXE
gAf+bTqKZx1wd4N7z1qAyiuXEPYKgA9riKfQbB5B4VQJQDqOYNP8yk7pseMinRkN
Hw1MDsDjHMa9U+kL+3G8Y72hgJfVJmovNktmaDNuKaeiUXeT+ry2YeDplkz+w0nN
IReRcWfxaZqDeDMARUTss1VLfgrR7AnZDmy8FOng6ruzZlxhBFAwsLU73G5K89oQ
WRHiSUie/TXa4SaU2VH3R5zdXT4qa/HulfNdIpob2katIoVK4vCv+AqCwB82c47X
uP2K83L6hZcjpuBLnQtfmZpcEMBuUXJ5NB78rSNhyYNFR/wa9lkyysY3Jp6RLIE8
4ERH288nptde0SQCqFck5eOETN65gxRYhZ1PHGWUIZS5hcFoIijQad6ou312wt3w
CHvf8m9LfKQzyg8A+3XTb//LKDy98lg3Yngod7m5/Ez5QAC6YpShGCyOdaPeKGfX
QoosguLW51ftT8DFN7KfVoBxo0RdQna2oR2HAfjASAIF8QJNfdJNRZTJVNQOrrt1
6Tk0C601liKp0Q4kjCp1jbEuqpa05nhMxRKFermB0HkNE2iIWjqaUJyxPFU6MzH4
I/sIkVOHaos6QSc1SarjFCZsDzRJYBy3of29mBZr5FHN0+1/awD5PNLLO5suxSn6
1zQSV7DefvePAv5P3g+tF5yvQkzoZWlirvQ+kGllwsjSbL6xJLGWRdSJHPnzfnu6
6OKrUcIbzRzq2+hibq4thQojiMAlgikLmVwK8fbhsMA4AJJPuNfmg6bM79qBjCdL
vQCyntf/U2uWakUplwTKfnPKosbqC2AEUTt7x7/qXvTpQPHPbuNjfxi7uJEjdikT
PvakK1r60YsKPAviZE0wedl0dHT4rJqmr4LsGHG4RbU2i5+ozkfv4vPJtc9tpg/f
q5q387FfCefgiDwy8iPVoXl9dahV0usm1VDZDHf7+GwexVnWoFBdXK5SBP142sFm
Qw5lt3Is8FHzDdZN9rXcQK1n3in9EAAbuWTtUGdwOHu9lnU4BOb1v8vqF77eR2mB
O5ekrf1vFVaeH4KTP/HgxhGRmrxbFcTmwOX3voSgV/WO3TmbuMyrfsU9eMt7u0kQ
uCgjzw/KvhskehhHSS5FG5eRGRc/UubbGy/SXconcy+EqvRBsTFN3gPDz/i9c0p4
bSejz/gFW32bLtf5MogroI3lwHLgUBCrQnu2mMB33tfFAphef/NWX8yNLiGwqQ1l
SD3Mc2dYOR9q9LvCJXdUJyTDQRYNNbsZOG8XPjAIC4ox/Vcjfgw0QzQDvTkNv1SQ
rva666yfSCsukQbMtDyafoGXyQGcRBW14fdrK4Q93b2pjYmuaCwGPAMH0eT82jT5
kPZIbhxvGCKH2OUtZgY3ue21tWomzkIQwMO4HPLy1YcZ2My61UC4uU1gE7VDJyPq
YypxQgLr7an9RJNbibzd/sNB/nnKDPuO5LRyd2mGyjdZJX+WO66KHjGMKU/fBPCu
02o6UQlWXQha7mBwRJKgWGYuwZyyDWW58hQ+RPRV9s47d6TPhHciY3u8tWKeI3oB
SVJaB8zY8+Js+UsHSmGlxeexbyCtnaYEKEKlGzNW1rr98XEVie/vTGGnoKv0oOzx
u8RaLgV+ftaX49J3uT9OxNwIh2ESbEiWCwWWc1Neu9wZfetk51U/TpTSK07pLkCs
NpTRo4DtDqspGIghy8F/Bxlej07PNFSM0GQ7y8gbLWoHFLdddeluJTlChhoB3c6K
dsKAJJeTPUgyC0PszOYsemoXVmg9ubP/DlHQF/2132+GtrQWaMDcG5aXIzvo5Rz0
udTxXlpvaHEryswlUaeopROw3+Dua+3uuoD7s2evIYsXKaRhL0kDKILZZNmyNC35
jnkcUXzNtTxsQqp0yX2zHGx4Z8Xln+A2uuehIwIp58dyLE9NxUUiMQ5Mw3JUY8bT
w2DekuhN5wDWG/C1k8kAusWspTB5i4zYbJxaZ+8L8aMaYj3HB5ldI1jWrMKtmMFe
U3FzDW9jRmfb617mqxupx8NloprQ211x39QS5xjL5HEMc9HpPsjEEaaBmKsIsQmG
Oph4s+OKGNEAPNUe0+DrQfSbcJJf6dmUsrLysEc39kIKycnaIL4BetB48x53GuIk
eJCYWXJDbxljkXt0uVZVvVTIyzCr3Xk05KxbTE01tv7VsWUgYwlaUEN8HHdKHUgv
fiWfYTuaHHFbv/O3lU3JIqMAGMj9rAMUT13D6KbnLQuHZqtjJBmRhVMl+px4QpV3
2FFMJ8HuwaAl32luf8LN9D8zZNvt4jwyE2Iz1jK4WU/JzYdoq9M7ljqShAyFeCbz
FMeGjOlB6YQaTEV3pRxSC4D48TBqa+x7jn70VfpHdtpqlGPW+SV9JWgUO4UUg5KI
iTacc/eaK5y0Pw0jRykUm8cv8F5uhjGHhf+5ZaXSEsW+pa5uOOnS1KfunM0rMTHC
fHUhBEjR2UoNcDRYjkJA1YY6otFxyJMQpcFIEBILqEy7uY/UliuCJCKTHso5Clns
2IsE1Ho/kBsZ62X/W5Tmu28TyAEuqbJsvHrCqrvGHhu+0Cj2pic+AjmyLVQVSuux
WaHGsOoQeVbPrrhqdWThQF78RGtVnMe092or7eUm57kx7l/om+5vu5JVFzGeT1qL
6tPHk4eMUZlLChRFDbWaJdarvGCplw+wZ9VovjG4j0HadB1mAxEEwoneNSJQrAkR
y7f/kbNdTUmhZUVZkjpZqgvsQ8UJHwpHw3oQnagJ4wpshsDdqT+nNheUlKuRaEy0
BXJ4tOWdQ+cJyVXJpWoL1bt7fQ8ZJ4ebcub1tS/HzdvZuJareL1UEzDG7Py6dZtL
/AOOlFRW6YZWAzmpuU/qaJeNiO/zI7AJRiakcu0hYX30AUXO/gqX1wReETDzYg87
Z/Sb/5xg9u6YASibPPOce2lpeNQ9oHcFnJF4PsA3PNfgeXeUVkD8/saTPa7pWuAW
FfpXrXdZzKqXO4Nh9JtxdsbPoOgzBq9RLi6y3VG1DMLbBPvIVo5U1FEdtwpH7wUC
4NovkT1OmmiIu+ZEkDZ9qUsw4mHk4a0WKwwyJ9aZKH1sau6xpgbCs70DKwAplwRQ
X8YI7b8FTlIDyLud1WG14iRBhuiLjs8r/kpmFy4gJQEvxK/MINEyJVo4uejsJgQU
2K2JcQ0gMcE5BJ5DPKQuXzeF1C4eQLtq1gwhX3YjcGQDjVAaF1AlMpjwncUo4odT
p6Pg7OCowLOVFcywRdca+xXxVFWtPj+reOSHx6zUGljlRkRWGXiPJByUpwOIJJWM
1Te55bD1nexKOrr2D6mV5d1fFJJYdZkQmYYH2iQ3Cd+FUQVy8a36/HA5Eka47MG+
ptrWYoI0pEYoXlGEgkRIfd71v8siKxcErdbZzkiN22wmi68AeuMij6cn9N7LWTiu
CeSW7LuM48Tdek5+VpvXlKeEVPnW8PGbON4Ff6zsk4JdzwQ/5plGQiK/UhYhEuKR
oq97EQrdvbtN3J0fPT1VCaePQdR4pZq8kp3A2PALNvwPkNcz5cbEpPNKp4KoNU+R
Xfu16A2mloxwr8HDDy0HxarbOeD4OR8wzcagLMGSbs9/+wKRSYPaVPxvLeg0PdjD
akiA6+2thHBbMW8dkSsCiTvvX4ELpD/atvYDtFyhp7pCtrEk4MPrCJdl3M1WR/fg
fIM02UTqAmDwIsJrSYaqm6OX7ThaK5Qna5Sz+HzqHSEn0cSEgVjLO1c04F4mWW9u
HXsZevqlxRCwfnmOztwBa44qJrHo0R+gfR75gv4+YRdI7o8o5jNMpxs9VrojB2u3
B2cKW6AFAhGgx234wJ2jopde5OWhPjR8Fozm+8WbOLeJ6ezzKUP9fAsoMlL7apZ8
m0Bt9gfm10uQBpHR7CFJb+QMM+LXzxwMJnZK6pEgjtt96ipLhAoEUY661e8ipp2Y
ZxNHH3qLpk9v0UDohfFO3ueBfxfAfLGR1SRG0DlvEJ0GQ1BcCryA8WfaFp/X+zxG
Hp8ZxLJLqcr8jX3lLUHld9Yaka8gsAZDBDT34R2+yGTeKChSp9MJns4iK2pIAqdR
CBVTc0hL5s+dzQrDlATjz8Y5/YDenber+FcJCMKIyP/nLfWAxmRYZ3yy5f4dGvQ8
JhQdn58HVcDUwhlDAxHfYHyN3hRalBIVAZ4itqaguAyIpYZomhoqSLs1ASo4xvRd
N9qJ+HfLw1mTUdkPDw950oLdHfCfd/lQM74rBn1Z/Kgv7zSa2VRezNql5YnKvBwU
3FddjCuCInWST3MkhNgNTXY/9ViokFI8fiGUHb0ijEqXmJMJlvZrztvnAKd+ZDkm
dn0qdp9oD7NgYu+UXtM8Y9nkKMUtrb8z5W4I+1BfNrGwyyHyz8z2N081Pryz930w
sFeh6HjkuLt+XmfN6o8Dcx7OcCiE0I1bMyNX/vcNPjz/4/EgCLJ3jEYMLCgXTXlK
/zv7H8TpYzQC5IPS8eL9XFeFlfnCxUPPrssO0pP9051xNLZDBYbvTDjy+7d/1JyS
3puffteqKYCX+BVV+6U/3IsjxiBIhJOMnxUG/Ly9Uv2y+oUwpx/rHCJHsc/jpMtx
VMImb9o6l5Fr1eQgZpj3M6g35aoZVKgP0BNplRXk8lXWwQJuWfT1Z2gS6O59hLuD
O3gLGTm4MwMr4M2ddXhO0PkOQ7EkDC4hapXbDYf40X/wThRXexUNqkBhJpvlXFgu
+HF5X46H8poY/6jOKsm5vQs0i1EgXzm3SIxG9JyRz2F4L+rbdjbunyVor67tihov
97AqB+RwjPyz3opvzy4lbsTZP+Goc2DuDdoaOBa8y+bVG4NrDV310Q3CKBphIj39
obV6pVdywWf/5nGXKTTNsHHHi3Wv4xFSMTQEhYQBY6bimQEXfBOSE7QnzGyMpELA
rTh62nhgyl7PDqNzC8TEQQC0vcxyecdFUdtryAe6GYKJIeRFnVJF0a5ym7C3UCao
rVNLGeWctQXthnLgOXlHgvJR3bgnkaiYJ/Oz6ngO0oyksjLNAs3BzcD/kVfp9gl1
irIlZvR98Xa3GLYJYWDwBUVUGpQSKb4KlgBB8t0i0LLZVb3VJ0116bhXcffklQPJ
6xphH0+O6y4WH4wIU5qLTOwYG8S9YP//RK+IQKcN3glkGZGB4JSOcgmGc1vioptt
IuUBQlkaLlZ0Aj2kgySph17S+m1EBXqNxKSmrjFErzeGmbdjHEug2TisXLJ1N/QE
GsbAm5mrfXh3XXFjafSpqOs9JMVU0NV+NzmuU7NL5bn1q9qSrwTnUUwv/RiJ+gEM
cOrzABr3kjYgSFDl1lmo7wN9nF/L/s5WnmWGGJUjYRnlMJhPEf/2+FSC3st/K7Q2
/y1K7O1UI1KQTI0Tymvf14zjlWPilH9ToogI8q97WpgDR3Pt8BCSzXMhKERd2GLa
6eV6Iawvd/kr0WVD3/fa8g/ropBGbWXxfFt0C19O+XFB1LU1ImxiRSFJ9ec5T5OG
BvY8CJOXVgQhATFVX4wIOFxX/sOuBCEB1vCQaSy4MwtLnSxVzZnIuDKzfquc2pQa
MZNlVFe2BWR9Jbq7m59VSQcH2gePzJ9P/7MgMYFc4thRCN7mKXN0FbfbU4RV9fPR
ZpxxdJfyYUJudibN3SY8Jljp+PPpeTXsXyO2bxoJxXVcc6IJWF+c/0e4gFol7884
9MVsIuDJcU/S0BZfzv8gCD8cWjuI4TKSYYeYR3XabYYZlFaBvATB2bgz7DKFDjo9
Q2mLdkA35AjJaEZY6x4jEb/GVxqFrHrA6a+Oa6xZKRrQgSIUQezDfIDqFa1TFKM3
xSAG8pGPDzxU2gqTUpX9WkylgxKm+HpsLSOaoIeHMCCF26dywcOv0vQNWCZBNKyK
+h1Wym8X2CSecD8omT/ffbkv0aeRtc1JyRnuZpAR71j7ZXcBzEz1FIfWCco3FxXU
mKKStGzybPbkWnTAkFAdZdu0yIEu48bZh/LR+mq8BaTe/qK0WQAmJYW1luVmpzoW
2v8sB9R0CiICiQ9brZBpTiTE75I/rLdN2bQGsaa55u2eMcFSXYuCuTmCl7f1KBOX
GrcvodsR9WE2cdG8CrHyYTw4wQN236pSHeLokvZqRAcT3b5QuXJPQtH8gJXeGFKt
4qm4YqeN/fHChWPDi4PXop5ya2v0rvlZwLywEy097n9iWl81AK0Wd07py4CVtkJY
jS6NWHzuoduOJmlb3QLRd+xw3vUjikSN7ovVnlonWIqNKrbPVBz3SMtk5lcEp671
S+mb/LeYlqfWLhd2n9g7Sh5FCveYCJlMi6bBGbYFUsWvfo2uIPFVxmm8+rnoPlj3
nlabn9yBtjj8LMQVxmWz4+sgLntcFPzhOsDk9/dosZd3nW1C/xAN3dCSV91bt8OG
STDGO7MRcIbBYS1Wxfz2+sPKTgKaYpjJM0i3Qdjht3nDJff6O3HtiPq52WJ3JE5f
m8vRhV4JZgz7f9wuqpZuknwWSplp8a2QN3ebqzMz1s6bk2I908fLXTap1FmduWhV
K7nMUecgCLtxtIVaA71OnpIzOob9uG+NkM/y42+JtiDpH6t1YyzWDcUg8A2Kia+8
J/QY7qCvUHuRVuBLN0FPVJUQmfGD33NzVunZsC2Todrxe6NQaU6mhu+jGOau5fbG
k2n8Fxp9h3mSv/+19T4Yqg8OO4Uqn5mzSA9pFYWv6RuSXLHbxyrMy1yiUPV9R1WT
dQMgCxNgH4Eg2acWQdkSch+7b+Fp3ZpZhrEEcXbUAbUl60h4/zbVcv4Yd0BQxBUy
x0Y45xlxnDl/AFQ5UsKunY/4dvdJorSeKN+02p9SEtMY66G3lBGfTPjsgvXLk2mR
hQTnWskqJVbfvPk6dj0psELlb+joRlPtAGpWg9Q54UvedE2qIWZo+aNziOtVtr9x
BVoBLETGJZHNXmLvgqj/ssujiqGGE3NHTrDkfb8lsvQ/umndqLdH9dsjBwwjHl9t
D28mGPHS+vThHy2kDGqlilWKwG2smKyWxr2zJuzxKl3whD9mkmP40RDeLZlw3CN6
HplnQb0uSVCkbw00Q4KH5cwmoxL9ZHfn9H02sURVL/uSkwlpVUKVCu516GRpt/dK
WWXcHS82728zXJeUfCSR6L+YlkFdXM7sbr2i22UDBlOmYp92XyaP72HD9XJOEYDo
cL5IrRj0N8sfixRhFrGmORCsgf7hVDPf4eJSdia49B2uv2yaKJr3NzEkDKIoxw14
s6ESebtj8BfUphzQjwkLNj+Sya22AFfQcoUPegqTsxbLWm5yFNp/J/kgBUw49f5u
+XZO+fQ+M2x4STso+LJqVRACxreWy2dd8xILj6xbiqfib5hr7oEcC063ksYehQIC
j+x/ilZRy5JfuLiKw05o8l8S1vL/VYoeDX70NQaSXnlFt/57Th6oL5zDkO6Wvu5y
12sFAuMNHS2W95QqGPOR8hetfxple3T24BBHKaEO20rhds/qxk+aNLkJfcc6rIo5
SW3ifE1lR70JdoUtLdKdDDasGM0r7YZwMDqmd5aQu1FR7V1onaAXLnEl1wKptuJZ
/CsxxaPizmtCbugEhGG/bEA9iyCkTDS6YPjqTo1hntrszZl4/Ece2Z646ZudzgqG
iEwg1jkvQPmJXCeDDsvjad+Xi8Hpb1d6Pcc5sC8Ft0UcTSvx8/ymcM4BNuxu3wg5
Aj5xYR6i1B+1ZfLs+8YXEA+10q+Q8Kz1uvFV/aSoEwjmT0UJU0OhonDYo9F6AXjH
dvjZnSRaeJqxt/Ta6tevtWfa8aeb+76DZTq5fTmtxMAUdv/YsBjtWzuWF7yXJAqb
NhL5Kf1++8a0BO99axOYHV+/rD8T1bmJpJq5mCe8g9c/XqAdh5ZFMs2d2WwMK2uN
t7QFyU6MCyj7s6WMz0ni/LwuG3uW1VxISTYPBZOBwKmrzR0I5FqyqJISBG5N+WIX
PWvHhnLQyJimpzeZivWuZroe7cYN6h7IXa1eD3x3eVf2YqZnBNzl0E4mOzJr+zau
ZM8hk7DdCMttvNn0CelvTvb7CmRko7la1ph0DBgx2Qrqzq6j+fKOvxUhCqvuy5TW
xIs44DBnkUou4fZsx0RzZEXt5k5G/TnyVUxVKTzW0JUV6NbzA1Qt+HhmyXQQwKjJ
VZ4Sb0D8tBosUySEGltpnQbcKqfFdN163dW21YQH6PcaLcbeVBrlBMX2PVojYckC
+JMbQVfi+B2WkKG+cfTSUw2wJ2nfQeLGeVNOm/p46BIIXcCYQUBXnfdGxXzPMa1N
rEnFLJNLGqzPe1i0t7EvqRlddGfdoynOkYVqS3ph2EOZDiLZebFgjIfNClx2yhoH
UGmIY0Xutyn1w8IS1k3Xm1meOH8exvV+7L2YexKIvtr29wnBS7n3lrAuoIJQyGro
58fojEPVZy47RSCiM8rGRch+m3VgnGv3cci+gM7IOty/ORNqoyleaUhO3A6GRxfk
jNK2qTWngvAKEfDpBK8Z4LrhXfbTUOC8ZeCIJNt1MUDyH8vNeDMVyT4y3cWmN67d
RaqA4yCXk13X2TbR7EmG7+leQvVBd65XUcd6hb0U96bKPIadNUqeGQDWL6PE0Ber
+23rqZr2YH3Mdn94ZnaGU3MGXPzG0HnH/TFLpImruyWrR25vn75j+6I9z4aQGiAz
+yAY8HrdDn+JV1YOqrYfvOaG1KNRLwzGnP9HjjX6sRfTlb+fgq3tmCP9733KjqpT
5Uu4IClHL3x+/6E9htYRxYIJAkiGWTgwJVuKcMtMG7kLG4EApBujxcdSSVcWM4yl
Da0/a+sdTjF3LRkqvgxhCmoeVzttEjns7DGCYbZLvlkRsShEOemytx7kV5Ji0cK5
yzjKhp5r66LISTwt6shA8fwbJip4r7AtG6Ow9rD0EPGtrQzBPZUHBjRiBYmub3eU
/9Xq8mDdT0mBW6v6W9gWccBf9PELVZUd/pFsPzu6IpZeDL4s0+5DUNrO4woE+17f
iOK1tSfKgB/jTEn/Qj9tAMWTDoWEWjzBtApk4UVahqfRijrzeq8Jdyl7sr1gehqu
w1hIc8DWJG7dkejIzHkgUdHZVHGybQGBz4XJnjHDUoX/4IvOsdVKhZF0oUJ2KlBw
wxwQSBlqVO/ZyYkT3wXFba2UgRs7iRs7nMJSSmKfnc4Msh/2ThWqBWCalPMgeHNW
DfVQnl/uTYoXlE5w158qjDr30R4J1ubPoS+piqJmQgzgoPyC6RwLVj9ePjdQ4Fvs
1VVhJsKii9Uuw2xNIuFk2Hdxm3ku7mqC+i/6pPXj8XEMvoQn13mlJePA8uJ3D4hY
urB1ja/Uaio+065jXbfHz/bAzPoZHUPpSnDCS/n279HZaf8zERYW67gsHiSP/WoL
RUdH/UInD9xJeevsLuVS5oo8lU+z5KPWyGhhIX/FEAm44r1y6A7KSyVRdN/WrP+0
ay7dVztX8Qt8ncU9/n2vx0LzEIrg1Kd2VJBKt6RhhjasYEu7SWERcXNrpIZbU8Ck
Cb7x7F7jFMf8OEL980DXGVUVAg7sN6CVfYnIpopk/LA3FQQYMFN4Xbk8CMjZZuzH
GfqUaydK13CPD9espDVf9TGjzrjZFhZOeOyTAflJWZgsd1YYtdK56BF6i7TY7G70
q5+SMd9LiQY1Bfid700Svldly2mJHfD2Flix5Ba99mggEo+cCJYXLtskFmPvMpxo
4vLwtOKv8ZbT42HGu5R/XHD0yEI+rjnxE0sS4KgC3rozVZy+q0qEPUaTHjw6BL1E
LtPb3o/0N/5lAbF8NV25mzIf2Tf7rM2R8AGQ/Mx6aSTm/cNgEII2STQEvLrVfcRh
vAoP9khBW0O2c5jLPNZsR70Wsy+SFoZ8xTunBxNYyP2FBEOcp0jLo4Jw4mE2pp4q
vsLe9oNEZ2hKu2pmUca/6KROnOWuXlBicUj/gE+CXLpXY37++aN9gpKT7kWnMy6d
si3H+HMgj6s8ujOSIzA4xz+3o+gXctTxNvwDOErcxfrWGX/8Q7kXyL8CYR02w5EK
cxIPIMFKh/iIH442go8CMbPaBop+iBQwppOZY+YUkgu51P3jYvp+o/YiwMGtWXXz
e+74ooxguHuD7Sd2Rb9ZrvpWcbFNOlGWvNg3XUwLBzEUut/+79u0GMLc+iUinshP
pyGKv3aQhvgAcrTETG+txkOMeRzbGcfNCTZaxE/5br9rXDeVw5RhUe1cAK5ZzwLh
cnagUKtxR4qxnIWdWq+5niI5S3sy/4gf84RRVWFbYOkiX0IfLmkabuGJt0jZvWPI
BIS/RJ3qr/oYwE7v4wPavHDwI2rgtxWORuj5iE7VP2rUUBIuKz6TopL+U8qcSUCi
zPfdvGMLNDAaRV01ms6uTlWWkAsrP8lE0GL0LKKwjnnb3IicbXyJRN4hVeGissh7
Rwi9qXl/QmtMLzbNGtjfxo5JVSgXSngiut2WMPaYIS8+UCLHhyJA3rG71p157plx
pecLeyLlgxJ+hqcUrtn5HXQ5JDFtBwgEvBvUODbJoaK7To9AZ0gQi8xAhK0ONKtO
pqV4R7bL/MffXNyMTJBUsXA1qChsaF9pJ5+zpc+CJOtVMwIrnpDSyTGMExbe1zB1
51cyg/Haoe0cmqSKhlopVHNO3bKjDGVTDr2aHfDWQrKcQ6jnZCQegAMTafmPW+Zw
p3RSvzcG7mCRjxc6msEyH4hqdEvhP8MqDkOaPRinX5hET2GAli/VmxXAZh4hI2rl
qIt/Z+96qqaHMwM/IFIxI3ofDwYNoKzJ2uSrYVXWJYawJBjWJKRSNkMF/piAUpaL
Dlfqn51PVUK2IHY13rMV8oIqBF49DwUQugPwDgUCOKrwxZJhZvhxibjE21K3rAQQ
ZCjFqZqWMOfiAOz0g1apQnOXq792/fzAh++G3i24Rf7EIJ58V227h8D+A77mvNtS
hmqrXCP1+xrOAb9K8jApmyqTcfEuv39GMtGYqkjs20MWrqJeVq+TuV/iBSvwq3Di
EVfOdJXAASn6WxKjD18H85KRPXoKqGDjLVaAMuLDGzykdy3S6qTDJZ8wjbEFnrSH
4lLz30k9Lv1TMvBY7+c+HsH86LYy5+ULjENXNhZ4x7BkORnM/ebaOJ/vD5//tY9p
PytM6LfIxgq8L1A2r0wyaXAeezwVBhu2ny4wCXcyvvnEvqRBxLUENBCtnVUrdyYf
6fFvwwMlGJpDC1clKDxKchH5S7xWytlSwB4emFeyYxxgO0FM5UQSgtHdgBvIGG2R
zNMlyS1dRjeV0zrDN5vuINAawaXi0lhHhdBNwcJL/d9Kw9dNO5elvYoa6y6mtIg9
/VAzCOEhyl3UDbQhsmu681jM8knJpgoVx92ayC/gCXmCA5VMszx6B0hVQVQjc+G/
ACb3e5k8bE757I8IMA8FRHC+aKm25up76bZfLxbEvb4yAXgwWUHLPvIxoSdhDKam
qd0uJU316mZBq8HKCUucf29wXxccIimdofc2KblfjmykyV7l0JuRZGnnXOUdrocu
QemW8yeYtrRczCRX8ATmFnwrP1Ik5dPfJ9hCGpP6TFMzY7tvEUxpF03nu4dVS5Ps
GKACJZpxAHjBzPdwg2FrebcHqqkys6nTESGCg5fq3VQC40+RQNDqz2MG/sm0jtVT
bNyZjosDnYEEfOJhnoUp5Qp/SdBocYXirVqtALroP6ntnczsgeBcOzA35qBcNrS8
qMl9MkFbZmzPNM85+seyNM5S/CL9FZScaJhg8EL/B4pv7GK/mPKvZOAqzF2xrvYM
31bmIOAefzPLVpDbjQm9hgiBDXpC76NLkj0yTHowNM8WBKemdHNvD3AYNpSsewoP
ovMYcBm2IEA/80x72EAnPyGGtmy3IzLjwaW9AVsSPkWC3V5TTgwASXwQedl5ANhE
pEHERzz1cVjkSTw/3WcWqMRf8AleR+he/4oZz2jxiecFEUTjrAxWShH3B/+lRGNW
YfOPkP7CoML5Ec+NIoGRE7FZkAZcudFcovAoy/lFbG1m+LSRxCYMiOmMH7UNfnuM
iTbKQhWuLs0gyHq1VBVfZuzlfqhAcLjRfWtfaPebmORnsF4Pw6/smB06QBFogVgG
v5S96i8V7KX1JrK2gnuZVLrqC1KgukOLNuK1DZou0nOPY4bnNqEew2FGDfjAmbnX
jlgrehUDwNjvgE/843OUJuogW4Yoc0KYQszN94O6Js7o1Gim59kH50HOpTblyWGi
Pr7RyPgAJReOCQQnWxtodnFZHy1LVGaMF7/qcI4+n6t0yE1AwnGFFyzJ1Z/9szv/
yDZLWTvw5MOCEIatlWwN82yPXEUikYVH9KBpZpAZHHUSoFYBEiFXqHGroib/RWdP
zHD3gJNM8R2VRcPn2POqlkaCfOGf+Y8L40U2dq2jo+OUcalvMC2WUnxhkXad3suR
VC3azH/PGnmCI2LLvdNEPo0tJLkqJhr0PTTw47LPvAX470Ad+kpI0KKhvZIFovjY
aZ6J8ioRe776LUI5KjFdSIYKCISUMBldZx6a1h7agW0wLCqwT614vPdV0tj3pqzs
RWuqZkSd9zGGno0RVPMYtRYKaH2qGI0BFL+lsCSNrCFBh/lWNH3nlPLZCaR16O8L
bf8QcSGCkgknpLzkfu7W21ozI87rm//RyoUU8uBfS3b+6Mr+akUj2ybWnI3BoweI
R+EYYCO8vyTBvlUHOt8dpebj+6PSXmgQIsgpwIleNPY2hMfKMY9wp9ZMKTu/TJRt
2UZz+Xs09NdlHzwKRstL04gF//6+sR3P3HQ2kgjcgSw530Ey1gs+YJfKENuNa8pQ
fOvIy+ajFNucc0KYDfDKvSFEHd+LExtLancyXdf4AAcePWBrpKPXQXXs16kqHXRu
0zaAfE9H48WzkswPAVQ50VxB3Kevcpa3ms3xQIFo0MU9+FAxABMYbzg8+4L7bxgi
sXTDUDhLks2fmh3NGJVtgdwjnueYDOsw1yaRf9LIdXr8iRQQKEfbVm+NCbwT4IOB
xHc9WbVoMefDUj4vtOxHJ9uLKxsOxzigXUDJpXbhAYnlBgSf9MaPyUoV5QuggcEQ
7zwUJ4aN0/l6a0ofTfDsgxv4M4VNrx2h+2YiibN7Z4RSw+7w30JjynvFh0WNuRg2
xws6orMYE24D/OPR0ShZXyOUptHOeQJ1C52/QT65UCLhTkLoGFKwzPxS6D9vfOHK
aENSeLw/4RTINSoQQwJUuyJIjjDLXk1gGjV+i5jnF5mDlGGmtYgQsGCQr2FCxd9Q
iLd6MTc9+QN/Mhl1f3OmxFNazaIAN/3lIS50DnxciMpmHZ0RMCsfqL+ILQCpSni6
SIxMlbGuW3Iidt0j14jZhFZ8fhsh6oDGHb/jNw4NR4yf2vVW2BNqDMP5fbwpPa8A
xrbcddSWAgFBP8u48io/YhHZfkv761fvkR2Y6Bcm6wSaf7SgOLylhwSx5rFPEj0X
E94prOjagEPraVNrUQU4HJCmz9Ca8ZBzvBojsuQd4EvJUn7L934SEss+T5aiji3m
rwr08heXeCRY3uvLMV3N0jZQFiN0/EH9A9PrzyEAXXe0rdZ9jDy+vIK/d/zUmuB7
cRXh69qzUh66cR8qAHko4I3R6XMY9QtTf3kXJYlwq1hWiPWYPaFbhaqxBNr8ISOc
d9qR8dAKOZqOJuwvMQ2zReXrK2Yl1icysJXndmCkBhmgljJG4RTNynQFHPmiZ+Qt
lvOOwWN9S+ysKrikgXO4wMbmpLBC/G6Dq9irU9+/zwb8mmhhCqEjBE3E2rud+U1U
UGEx3hSJpWCm+OSXhMREEnJ7MTY+2YwO5xwqnMmUnv24Yu7EvBmJuLv+cEUd4FrB
/6AaIuxi7Pk5zOV8eGU37MTGmaJRRMp9G7a/HhdKtoTvY/ru5t3hiyVRghO3e8Hn
s2JtH3n5gyfs83ki8XBV3dkwzlPlsFqcdImUeony8iJXs1HnYlTkKuwPjEh/Hh0U
pDwM0SFnaZGOGcP56fk9V+8iVzhNpIWQUb9uOL6JVaQyta77zZMfVjp22gEbxnBn
Y1ZoAHtdJOSzu1514i49dls0Ty+OfFvf/v4ht1vq1aR46GsHsdGZXWTUqAt43zp+
j60ss0ag4U1eqEYblsMK9AvIxD0HJJJ3MO9gca7NDiDAa5FczVV1dYL0NRIcqu2v
eLtr5NP54F3nUHed8adhqyXuNAX3566rNpw7fb0L3R8mRZ4zGDVXrWgKTR8LgudV
VGZVxVt2v14hqtJ6m/HCfpwMEdbFn2J83rJqxvVElPT8xwmnLMkvBTSlZ4XbY2JJ
iuyg6z2jHj9RBLuuwUKLF7UrI0OlCADVoOPZilzEQJK5zlrvuq828iViVq1TLwFj
WEXpwQQ39ecAcyFkUQvY9y30+P0+vk7TnI3okCZgzfoFfdbnaTDME2yj/kHz9Gsl
j6yLXCpd9YfAC/Fe2w2W2xuJvhAOdRA3FIU4W2/xsnbcYsla1o1Jo7ACJdJKf25I
dcgO3fKemGtNxYFbCF6dJK5KB/Mqc7ok6lTYou4I6AWEfEnCXfPBB0rXbwoxNNB1
dfViDhWnk70XjbDmPD1Q5ULad65HHBr2pw4uIL2EeZ/jR/oMGLIJL9VfifLFWb9F
8wm0xvjzVUnSM28sarD+TZlK0JA9naLKXbYNMYD9Xi/1moKLALM7nQGHBKIuECpZ
0Uypw4TEmErpYW8GlW2wD/3/bAlaJzUGOCuS1JhubKAyi43sQN80SpfyQ0bOuPHx
/ClCDxRC8FQybM6eX+UhOUo7b9mVsg+0sQVwdZd+mYacRVOOE5g46oZqKfJWNeq4
Bm/DkoKgUWMX5udURQg1wTTzdEH5jx0N8xWOBv+ZlG5JpkgqQ8H3AdEwdK/c6K/I
67gw5qaH4234X5k+HN38JbMwDGMoTKVomad6IyB7lljV92+Cv2xtjCMgTM1pOA9s
AK4B/RKxZ1SdftvpQ5wTsldOnIQhNbbp9H1ZHkdtns+cuZPcjKurXbWbxNnLdlWe
X+MQk1f9AO6IlikhGUohuAcx+nQxvIbpgZYBa7QaeyMsLIpOaoEysRjG8wdisVFn
xknD5WClndyEEJEJhv1xcpVH+JzSr7+IcylS5/BOHVS2YSy5OtgYp4AsFryTGdP2
yswEXRERWDu9hq4lE4mrXdfoMPJAmga+mi/zZcdJ8Cvynqy5fXcdhec9D2AHCNqr
09txgscpPqQsc+Vx4vRRp9DYIKkaqQ8/pnrarjYiJWdTHSv2ZgM2QOq2DSGSfUC+
qMIM7JpDQGNtxjZ76YMefIgc724NW+ol4OsnVYBSzgY1yg7/zWhSq5rcBDecYQVE
tfRmX6hQOi2bFnK3PechITro6v4OVhLilIeMZMM6NocK5cNtsK+kzxY5gi5Fas9M
sF4rjDlcJfxQ2c9frwN50qjiOJevudQ/4dFlFtk1lWA8qh6sFTSKzIzPadyLp9pC
4O3YDoFg5P61Zc/WVyeK5LMeDPyuBH78PJWd89LqFdw2bhM52ygJwbGeLqyBkM76
rngADJa01zbIU8nYtnVHA5XpjlqYLGx4eqCI5NLEj0pe00MXWsaEQ0S9G3V7yJXS
8VhSx00D9dtbyKw8pWCeflhIQibj0CjKC1POJevhq/YCP1pQYNqaR/Lvd/gojL+3
PhXe+Fy2lP+r3SOMtfuDwtVKTF2oFeZR5aYx2VtccgcdLD6oxRsErxHE3hCzm/8R
xnUBZYLmfZE7Igt3YpswTmdapq/uexQ1lQxUq8CwrIAlzK4vghIYDUs9L6wiXtUJ
WOlfY/epKYyNgh9MvPvuTB1ePTCsnW4gere+16E7fgEMsT4Ahxg3ydlt5Buyiw52
5Bnpe3L7ZijAfut0HjSkUCh203uxzpHMhhyFTECsNk6JArA6Olsx0Hb7Giljzx0t
n3JPhuNTOIg1RJkTzFYfnyi7xF/gviMWdZy9Uo39a4VPCqZdo7w0v4kp0/fnTDMx
AxPE7ffjqtpbEDHK7Wk7HMD0d3T+A6iF/6H+N20jNAsZYFrtK6gPvFoSfoxzRxXm
zEOG6G3wXfNtz6bdBuBrZXbFkXE4kYHf92c/ZqBMjluvTMT4xiT5iCc//w3UKzHp
OkY6CvOf0JQkv6bbkMJ4yJ7/uZJz9s0KsMtkDujrn/PWpYOYG4yije5eQMKtIg+Y
QeSPvMDHbRcC/n58b7NJhuLowJngbPA/h+8GwETGlTFPCZ298FO9NyfWxM2p8BOg
f37u9wvIqWzOPnzXvJzo3V4AKDEWkeG1Eq7YHQ6JavDQaxOCHW1Zp3oaP+6HgRE1
6dSD1ko1jUDV2CmX2apOBePRodwwiRczGyMXNInB6PtANvZg4UtrEZOJRm3+3gpK
M22ebjqZedH8yP4c7OTVLQt/qzl/yhzIuKxnpLhQFXHO0FudbgShxvsSEN6f1oob
ON6qJb+GuEkuM7W/utJCenQnHNtm1m7Vj1hZNoaHK88g8sqmGld8TcWKh0uk9n4j
Su/SAESGVbKGvODF8JA8b9tilL5xECYayyVx11l3ak1yQr9/v3Y9WV5cxOPR2T54
Ptw9irJpj2mOYIOIyXG5T7m8cNpLjXG/iVXRXLWvJrZshq1OvzZ0Mx7lCty607hU
o7pMIMbRJ1FK7uUJkhorH79plCYLJcPgl6b4iugPhBcBg8zdctPUZlQcL6DQPxKF
cfvSzUFAIvEwfd08rgplSI6D/6JWZzSBNr3nRJlz+0vZi6cwFncspznqn3TT1RCz
bbheWm4MhpiFZ8CRyn5aBx7sQRKfG+lm9HQPSdEvaKcCIXsuCWnHpYIqbD/VHakQ
ZKEfTTTbfSeE0R3VQl4nBTAKxqmlp2IY1rZbRXNvmD9ovFNuYiroARguBXlDuv2G
xu82sUEQkD7unDi0FYuFqJuT0KIssrVJDa80AsqlUeW1/5yHWcZgHnjwvTPrCw1G
pt4/cPY3/Jp8bga/PGEyNV2qIQ61IwxjhCTklwHrQmRJMtf1QJyqFnTCNax6tUqQ
2WwxoprjYEobOXvb1eO7QI/OLoHElY4A1O/CnU7CiBuJtqzearepCojxnwGD6wC3
06wZSUDsjpD/JKxFh4qO1OZ0V8VzgOy/a/uBcVEKbd6Z2xkduG9badTlZo44z9EN
P2fF9fnFqIFaefyqaHcTsLAZ1xpfGqXFh7BKP6mUD6LmJrfcaJ0o/YvFCZ6y7AMh
OJ4DJclbt/HHBcle1xiZ/sKC+U2o1ane7alOFL+8PLRQrsqiuacIh8TDFFkZVbK3
zzWOnpC2cRX4bQUnkUSoh2PtDX7QIVuMP5KBPBLO6ZZldOSoSsjGWjxifhMy1sJe
jcX8XXPthWMWD2b+CEcuvooSa+kRD/WM7MeLCN5X6IH4TjSvQZNlcJK2L1FlklvS
kxSYAfRbNvYEpWrOyGUBq2i/hif27XmtIWRrf4hYMS/NtixMFWTLBZMHaXwvJjEA
ln8khLbZihMGpnObRNx3gZ/gDPIyCYNmd278FypGcjXKFR4tQxOGHykMYo0cMyKK
g9pAYb+pwxzysytDdIPNkKvctcR7UizpRZy3U4fGEKNR8DpjdEA2rQwwEGlMeYVQ
XuoRvFccf4hcQ/8J7oQ+hteyNVU2WhJHHMH80RLUp3MuirgwCTql8NE7IDjyq576
YLv2ZqAVGdJjMiwXB7Wn8wDrSDC3/fXp4IvURH5PjRYj0smPUQ+DekraALVgHx3v
nuDgT9wyspj57ZS3YFmbqDflYfmiLyVqXK5QBxMZhT0fLXgc+o2yffzF+9ZHrbMs
LTbdZkNeX8Bfb/T4lGb336QGpEI/pCKYnd4UidnBx0a03xJhyZYYeObi8fxIB6bn
J/HgyHvbmaHTFZROmnodwuFUnAS5rrvwCeSUhSlRdX5HB9RZ95L66JvxCSX9ORCb
jTjnVwGLQ0+kLt+v6RAveWwYDrgmBtHrG7ZK059Vd+qGm/vF0/jnuoDbAvZuK1F6
oEemuW28A/JnWROmYCdwaylENPw8povQcxy2ujSV7XRoSqUG8dFfk1be6+8tV5ms
nCIyUEgO7qcOjhsoMljcUIKv7frt4mJO1uL6CF9ZmaaIrWXtclyynTBPtPBGX5WD
SXv+OeLd1QnrXHBJUzUTCREg12Od5AS5NE9GDY5uwFDaLc/4cDjXTzFLQn6jSydM
BEFWZFfWEcqjaKePPiOI6dsK/Zu7dwXxkr4QSy+0aObzI/bLrUj53NH9yN3P6cYF
T6uTxupEvYABPWlHuRzhgzeDSDr3544v5ouOu979ObsTPixzAVfkhBIdYrt92KPt
3KH09BLKsHZ0C31XMFvIPDpX4XOfomlzJnT4fdNXo8+HE3jkAvkfubz/mCmd1CMA
wmO3kG3ruSOBJFd6iByR/AdtQx+XxCG52tidhkyBdjk7f1VlIufST95d3Sm5Eq3B
aqoKBclZYnasVap20cKRf3mN99ukflPWXdUKjuNI85ClAwg56RBQB4b498TotGOz
neFQLjCXqyGiAQ36opzWBvXqBD4pxrzkMk6U/asAG+RJ/2309MUEBArVUuCVmpD0
syCFx7797ZUDWWmmvykO7/I4ptWEsNZ6TGjq+wQRCFgW7xe7P4NcM5+vsPsyVlUR
hZNcXNYLvkNxs+1UetikY4+ep7R2pSEG97M9u6vbDKoGWGcmRNCV0xv18PXNik9p
hkqegVwO1iz+YDimkv8MlA==
`protect END_PROTECTED
