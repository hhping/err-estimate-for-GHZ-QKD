`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10LHvWUdXA+7ZshyfnU3W3G9xYoSY2LQWTuO1nnzCtz/S2XuFZ2JB/tVTGfBlnGf
lFTbLd0NnF6YviOfKgYt6J6m8fRsov+Ml8fjQCmbUNpdxc8lXfuSACxy2IOe27+c
ibWkJWyRR6NdDIimsc+4HEJzVlz0GVA22WK6YBhoDqkcBoNEBygThFJBkYsM0dS7
auGJ0dDsCCJE5UpWvhiVaYtZKJ9vgJME60r1/iecKKtnZla3oDYTzfd2q5jNzd0J
V8uiyLnfXbzReifFwUvdZh7cy9NPBVYexCy+tFqQ+r9W+GKdREt6JfCmqXT1XISX
E7k6G1YY5O8nnU+CMgbdf6Jik9vBGzw56u2DQdtzR/c61YU+nhuFEeWo+hZQCOnr
PX1TwzoCVt1VEo1gvKhVaHOxMDfWSfLmveYvJH42lTbwHb1iAm/2ITB9hZ2klq45
1E8aeNx3DsUlLlt6IhKTopxwcTMZ8Y/j+LYwbAhLqlc5cvNSlitX8nkbU4J/eonC
TnedV9Ld9grW84gWBnf9yB5HCiFL+uh38P8lTTP1E5CFRl+OiN9Vx+hj0GW+RGAz
rUQ9MfFJmqQ/hS1ru0UcWaLqrgI1DV4ZrnxDawbcmZQ9ZxCSR4ZSjy7kyed/G/YG
6vEkE5q0i1SE6E7eA3u2DL0dXVmVp7T7Fzh5yFhlzgAzShZqlgliqtvlRkGE2lBc
gdLhrvogUlPn282wjE9nX/ycoYatyQbPmHUuJcoUizMdbQ9mngdc0qNw3+7RP6+V
OJYekYIMy92GeTIX89pnkAn92c175GluYZlTBiORVTSAMRXAUw6/q2MSvAjWDlLI
sn6XX45SKmyDGoUIPXFOXWYLq3c7v5Jh0k+6HCge9WbIxZGB/8cJMRZrssF9KAEF
RPBX7Eu7h3ExVtniNmvbqpFtD1Y9WPCXAN/gWjv392I7FKJCDF/oYEpWpG3CaUX1
hzhAAqWZK/WbqSovheDKxWjY13KJOezO47MK1V/0EH/nkCM0Mz0FX2iB4lOCDuUP
5QL7soq59GrhcrVpo+PEL9png7kpbi/1gM6bWg34jtMd0azGRLMgHnrPaV+0ltJI
6f5NW0bkCHlZqNBFhZGstjsF7MrXnGYDjR4GCzNnh5+VIi7Ypcdj8oY7JcFMahwG
LgEGDst8cZDc6+wSzhVgmGLVLynC+sc6BYJTMJENgYKX79t1TdHyTbv4YhMOsotK
aQA1qRBewESVSrcV0ukKpfMbr5VW8yw9XUO0udsTABP6N/JsSJyTVlKKqvNuIWjd
4IzUGThfgoGAPDHZYA5xhxDez1X8RDXUzlaYO9opd5EISb/rVQG7Mv+HsbJXpnGA
/o+eONgGa157YGtaYcJh4sBrHWA94xKDJeTEXNECb+Mhm/tZqufAsviyTC8we9us
NcFg6+O5kyFZbBbTRXu10UsOKAcirTuVZkZz2TYPRjfN9ia7QE2Oh6tsCy6cusCv
T2QYBOeh2H57N2XyK1S/jXntrYYkc4nzASgB62cHFfILxFFOjN0ih8yaS1Fex7Cl
Vjk34ng+PK+7ZuAmI69SvgwPtcW7TgZ689dmdLHqECawA6Jg8eamiEErcQ02dzUy
XtyiKwZRAPpSZrv9n7w2TpezJdcmMCJcEn0B18sw3MUhUWJLt1FbMiSa4u0ZSpll
wt6oyUtG7R2SA9JEE8ORwzWn3O9I73MXwtHl3CtjUT8/Wu+azuir84bfZ4o0S5BZ
AcFIhOGKikoJzw+COG1V9JlAmtjllWgfu02kqSlpV3LRxbmssqvs+FSDUn+83row
vilu85a4OjOxMN60yhKk1TbTMQsxshMugTdUpjNSs9ptB8kgOeB3H1lkDuYEhqjB
ptBlFTj1br4vpEM+QnIjuVRHUnTRRspF/SaSdXAXFPrgsXNT/fbMe7HFk04QBhlx
2h6L8b2ZnyM5cjelsZ5bXdHvl0iIGLpV0yfwilK8YWtWTnV4N1txFEUkPypaJE24
NchggN54XKGMY+UslCooBGXa5k7S5OcwAQ6QRMurS8rei1N0wS8uXReRJReSNAMc
9u1ddOxRVXXL91nsteKkOTZVbwvwgMyIp0CsqmuhYQ9iqXyhzcRbl7Ko5ML4X+sG
+BMmvUgG0AcGhpYcB9PtoiiNrM+zSAOfPmAaGkc8AFwmybQeXJ/cBb1YbNV3gXup
hKgW03O8ZS84t2E7Qx+onlMlBGvDrQV8W9Fos/Ww3VJxU509LGsqQFC3gmpwjgCI
67L4AWw6qZuXMYx/x+otRoiyLf/RnL+0DKxJwJcb4bdyNg+3QdqDvm45VsE6F6Ur
THimLHUSEdwuglwTxQyZtEAszeLT3kL8CF6bpWdTIMFF6BdpOdtbsY0hULXB7exX
7NVi2x/zbnLKw0W/6g2YDeeo8ctvqq4SfIsdFEGPGGX0WUkCAnKBEmoE2WNpeTQI
rA/sogxl+RsYYRa0SYMtqVxiQNxY950vSxCMAzghtBiTUHZqdFEkawY/tvTDGLmu
STM4BO2qkBkuHSxrKA3Fh0C3iPZVn4UbfM1M8ADDMS+BuX5XFWcCz6aD5XS4nhEB
Urz5nPWXfc9RngtSaqoEIQqdsH7j8junCO7DxEbna3RgIIawso2wpdOjRPYo3aUz
Yt51ts9yAL8BxXMx/RCrgqAz80KdjRpBLqPRlE2/D5oJJYKSXWYxdDbb4mgk13g6
Bv3s4jiKo0GaaMQ8QC2XiutTFPuApkiMXcM5hfPLMs/pW9O7sIu8v806CpSB9lI/
I80tIA1Gk3O5EDIewhPz2GEK3NKqJnj4uwYwztM6sbksBKPPO0jEb4jvW7P9P9vX
yJGIHDfhr1V/99EZDL93pz0/b1qzysMLxP/JvZGiyN/wDGwZOo5Rp6bvdkkifigI
Bb0EjTkIcK8cV71MsSx6Edz43bG7V/jcg028pJ3yc4zaR+f89yDzucugU1FMd/VP
meRI++jMACGg+dlR6DvK2FjrGkBv85OXRCCmnMaa+gy+/ZBebupXBYrbIDNESFmU
hEogie9v5p/Hs8/Op6PJouMafjYR42pa8Z5o0BhmbK51w9u5jpqOYoahVp2yFKa7
c962u6S7s6hc1oZ22iglYXLSNJl4pdYLLNu3uShTJQzEillPQOM9CLvQ+mhHfVHQ
PtpbyKY2qniM76gI8rmkMoXSrUKeTOXhJCMNBTIsHykT8iZSv1fpARZ+cCsINeOJ
1g15nMo7a/2YmsSuoTdSlHH0N8D2zGtPprNcv4Mns45wVSGUuu2Hesw/kggERBJy
mNQKz1rCngiHvaLfYFw5zdWxn89fwNlKT+WvBaL5EtiC854c0xHKyBbnmg+GcqJn
r1Ob/Zk7wcMLxTUxO4yBF3bCGwU8lRIW/vZD76HxkZsWzz3IKrZLPLEwDBv5zD0v
Y/pXpSNqX2D36kYOYLZrdHqoaX7RY9KotftbHEZGWKVJaLbNhkIavxcal3K0q5l0
UHZYCUFdUOFCm5DAsnzYRcxg3TyTQPtm/eGEenG8v4ekNZn3Q+GNa/6AjHrfvUTh
zsQwP0ALBHWSmy1ZclvwNrBCHJxdBKKD4AgfnZ3PphlLE4MZJvvScTy3oEockJrI
HLhTF3M3xiK/fvNS7tDDhcLcXE/4xl6QZh8b2pqcc97Sd1QeMYLhfsxdX49sLIj/
5/x0n/pTojypLTttJBykPd4CDP+4W4PwENiKsiuOcENppUyUTCC/P3ijX8bchXu2
8pb6QTi0iws0jzoxL/AMwN2VGzeRBEiFt6lozxi9eY5nKuOGDpypEJuenrP6RorU
sTKPJ++QoCx0w6opMh5Lk2e75Vhh03owkpW6M0TMPgDWH1TsBhW8ziaXSbCntGw2
B7wyjPrE30YojwAlTxSJ39KHV11ijMe0x2E8f9vkC18vdfszWyYIPY/hvqO6oRm8
rjAhKrkuuvmIvGHVcN3tMwLIciSz+a5HEE/HP3plNR5yoe2WqNn7Lx3m9JrLOiAt
RFGsBFPfGNdSPBZfR0X8CMasO0ibm6N8PN1iIedrrXZUQwY72oCWi+yCU+SqRZs+
dvNDT1vEW2yIL/BPYtea0Aqkh5J6AuWIkqJZIkRKYaRviN/RuV+8dwiGVnFTWyk5
LctRymdBUCJ80ykzxHtKO1sM2S9U+y7EWh+7OqyY/gppsrfAMG50GcM73TTpxRBW
`protect END_PROTECTED
