`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+knmnSA88ed3rSPVAhUZ7L6hXhKLqRoYrjmNn9763eg/3SwD+y8Rzv4d6caAP2l
SnqmxjuyksUHsjIYqXGzeKVnMiMYB6MaNQE0+uHGQOi7fNdhH492VCBrnY3mhbF4
kY70P2rrMptnz16KTw/OEMdFWhXotEGXbdNmWQ4rsPDgk+cW6h/GVP3mokNEa8Ks
n8ZccKOQAHV8y4prgSSQPuMF0v/fS8YJymUN3bq6HSsMlL72i2rcLUoem7QAksUH
UFJfiig9v3v6MgJy17kU8+l3YwI/y+O/UXqr6hbPIxtkokR2AsRY/yUn2HJUe6um
CRWEhrrdA0pdWi9+HI9yAK2S4ovmwpn0MGhreyzgaBQtDeUQRIFJzK+pF2MAkp4T
WUkKXayVhaBYfISYKZltehux69UYvS2tWXojxZsSsShI0Yfapc1UqUGKA1gAuOXT
anAKwl9SWbXX/JCgsLWc8w==
`protect END_PROTECTED
