`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZilj0crJmwDoJaIPUYQYQLe0mf1FciXcnHRtVq8gus0gYFwrnsATr7WdKAr6jQ7
KUJ4Q6x5qOpE00NxTQrRp9DRWBr3hOFMR3ll80CiZAhOVymPfbk4mAWb0K1A5+Fk
ENsJ5HC3IJfq9RqTegizDuhhmuh+QjYpIcOYh+nTOUFr1Iy+nHPLlfDBTVGzeakG
1RrazshjeWjSE+xLFQ8ozpHvB5kTEGGSw0ya0cDuigmB9bpAy2L/HDJl7tDNAbW1
G1AF1sOzIn5aiotK3yhrMkGnoF+J7pyP1N7CpjJHNH4Qu5Ff0wj6SAJRamyoLjUp
NX2bEbvbmMTzUUZdB1XdGQZkcCDmZanrp13xiCWENQF1bMYel4nfliPBIoKEWL7l
SUPog50ojGUKlwR6LnEqOGKYBgFwFXvoh39tsJxxvxa1ZvrsLWztEvPJl7D78zbB
GAMeza75VAuFt7lAB23boEPVWTYn42JXbsTlUnFcwcBg/9vLIZ5vl8EjDxKoUQvV
GlhW3RWGvhcwBNCH6NYGY+Cish6kHuCH0GxRBaAZT9mHvqbqGF8/foDzeNzTspMC
lL0vDzW3ixBU4HDQJD4X6zaEGENinpGuhTx7uqi47qJy3ln0jCMnYA4fg1MmxQHc
UXXnPrnCNkNlskCJfMuk7Z4UsDdUjZoDJRSJKiYkMXs5uomEpgYuc3nq4ENq2pGY
35kEMBkkr1SZjuA2j+E7ix7XYgXA5MF13QDSBqa1l2JJHdORAezu5AQG4ZpKCcXj
dsQ6AHTCeyVF2Cck7GYqsQGpHqtz+fOJtIUc73fu6yHb5sIpi0Ryif/JVDuxfoJw
9BkjgWsUeCw2gzywZhcgxVhgTcg5tBaI+evP3ZMTUpAixZeRrJvl4SmPPTEesddd
QWv+t8ttIoK6AHpA1424kHMn7SrtxiAkvxTMgnQW8MG93XLyMoiR07oMc+DtOMz1
v+BA7uTeoORIIgsNond7z0LleGBmQ+bSLtJX84pgeMv3kDCN1hBvQkpgEdNjwo9u
MdUg0+yhpcWX7aLavfBoT8u3b71lRPkay1rPg5HtZD6p11V9zf90JkQG++TCmr8M
K6xnHVEoOhVc+zhiejXO5S7yssYNSBSeU5iXtq4pLp2XaARHUJ1Srl50eleoAb/Q
DfuVj0zWxy6pec+cMCoTYEo3ugGvsLDP6G8QmiM2LhD1ndnaoGhIZbPsvxPWIQdn
fx6d7bUJb2rth2srrgogIb0U9bTZ2p47dBAP3TE0Jk1fnKYOJk9TPYMPsrFRY3MJ
HNy73YdqHa3oRf035incDhpdQbdVoheIJwiwyAgzNtTM5PTIySlgEdNbGMB7kmNR
76ik44diMP6mapCpXtDh3wnnn25r/MVrFysxMHGdZy9lPtcF7FSUmWKKhwpp9BTf
EGW7XBmjfAXCevdYL/n81t6553xpVGkd9tOBEwbV8FQB0Et9GbgWPF2E3OR6ZbLE
Gd0XlrPTU7PtDS11eS+gy7hjKx/aiGO00VBGl7xlNvaui6CRXnMVK4r4JUUhNSz7
lrhsgMDaHjwZ1vg73R/1R9XC0ZDmihOvNTnWyJrVSRPNeVDZLfggU3nu38h0ic+T
r262Tkuoe9jp+pLHPtO2wOie6hLx011AQQf24c5Euory1qjob7wt01+uJnVHyMN1
WPEMW/C3QRocPUhlq5xyETmrqD93VQJrUC2RerrqzQI1c6CXcx+50GGxH1aBt8Mf
FbGQsLtJ8GvJqYFHL3Or0n/lb9vLP7MJ+jVIUWw24WoCFPdo6411z3aslni8YAdT
3Qm+DbrcAH4beMWFLGGWg7uAjEvd62vYOUW7lTt32Tg2cTbQBdCZRgwKRYUUSJhm
+WtrmvhffBDm/XigrU/7tchvYyeYcBtB+7i0rrfajcBy4WGsxsHLC3Ucpsa4y8jB
3zM/TYGqIf78JgDNdydKgWOYwK8HY5JfIVGQzjx/xxzFOF7heMhP9Yp06dJct8xl
gvGQv4yb69wS3emN4s2OwYb7bCOp6XGjK0KMZH3XjpmwcRWqgpA5UXNdcYUTdGeT
O0i3htw+jzgtqCNAi9OVRz7geCKvnl/LGhRDwuvwTUS9KnUEQCDCWmlLhhkQpYYv
ueeyPl1jHGPenNVgSeZZX7PxX6/LzRQKiXJig8OJJaCKoADuVL7nTclXEvStCQh1
urjMhKujcH9zezntF2LdomzNn0BC3qSiUhDteotgUM5vsW2uZ0fiyaFnw+nG5eLP
D7qblZ0/btRB+3YCwfPngpYp6UIDg3WX71JySYf44mrfO7xXx/S1hZOrCj8g1rG6
33RFHd1+K2lP7qZnFVkRs3wH31dQMo0NIDgA4NaamU8taCsdSjxiBE7Kzzg43qAa
tWjS6jx6bXZinZWqFhrSd5/hSeEoK+OGazyMxHX4O4QKnpXf8dchAAgzx0C/AvPs
Btbh8OJxINI4Vemht5IXzJdquZlaPS0Fzu1jtVNpFzBONKBCir3exyuhV0LztBc+
YMpS+UT15et4wEaUDZBlEM68FNzFgWo0Wgx+Oofv5bZ/T9o55AURA6C8zembKGHA
kfkoKFSxtheENbJ0hxyqN04zo6EJ8BI7DWRnQOgE/88KuXfS+snC0f6n9V1Ybuxl
n2CW9PdkMNkSEoLNZyqksPf09TvRvNwueBT+3tWugLuqHpXVtgO7ix4e/qt49lzQ
KaqkSmz9mKe+2RCnwKYg0bvTV47Q0STbkbGXBcRTgf9EXhpvIYR6tKmKwLmD/+WS
b2AwIoe7ls4zcZdWXCMVT3ST242SpZiYjJ2DPYaD5MsTLuC0BmjgsmgEAiilBq47
vKflTB+LaEHwKCBSMrDKlKVag40KkArowm/W2Ccvm8x8ThyugKKiTTn+cJ3Zi06i
OOI9iMWud9sdp7fUn3T0B0fNwXw3X6WFwMeU/j/nW8ica/u7Xxn0nISwKhVCjU4W
P6Ma571GATxBMqLNJOZIZtbXJ8MIhiI5Bu5E+jS3kVv+fU4aylUxFzoqv2pQ+3fU
bynTRCASlyCs2dy+o9tCQRdiraadgCrjgGKHKafR593gpwz/IQ6nDtbnQgarzwK/
OXFsXTQ6OyuSGYEvvxtnSh+XClWqNM5wUfneiww5DStHKEwdYmz5ASkd6d+Ds2So
wUnLTNmb8DLEMLiawlCOF+RaZTJt9AkA2/a3Vwboc+Zxsb4qS9pkYYWzaCP8lp3W
sXyAnhMCWrLIliz+6GA+Zy/0HOy+EYSXd1vmgy3fmGWYKfntVXIz9gyWUGVDUJ2+
yYrLA/EScz9erafNcySrOTar244tRWX1lDNaK5i1nG9ckMzRUH2lgm3P2J3nwVXB
zcnG8jKUOzfAKPtFIyjIqr70lCFGx2Ggl/obJKMwD4k4zC6DmGfBM7tnTUX0y2kG
T8A2m+1BxVJUoK753hApYzl/k3pshzX54+WnULZORYd3nIwHnuOZQqPBXi0UIUUQ
AjwVrwg1dTt9r0PNJucGVd6ci0Y67bDZq6SGq9rPFFRaz3Qylsp52ywH4JtzZ94t
pGizBIyUU6SWsVAF+ET7toKQ8UkN3tEq9WPVUTTmnv4IAtb3fSX8Qs0UfJzQS2sc
I0pQji2CIo6RfJvHXx+Uv9322Ccwad2DcY963U6zoycYHnTL1uulmMdtGOWuROyB
s6g/vmF5AnXTiTzmcKRnBmGynHAU0QbGDffn6HBw/3zYw3yTdVhtj19P6c67vrB8
B+6HGNYeAokTQqbxH339BjpHBFzTn54Msde2OF9Sqe/c5nX456FFRQQp3OxajLdO
MM7pDOF8PEdc8MoL6rvTc3/NMDK5/vI/EsWwjtV3wu17TszqecyiAybCzAAs2N5k
jNSsQM7+5ibSfUbE8D3JJjlavJOJhRS7LUflQu8U/l5wCToUNlOJgILw5HIrSBme
jjBfQMfn0WuVH0/ytwvst1sOk18Q0pOEZl4gfg1Ux/g1uGO3olxl6QNzcSfprKP9
Rk/coHrEYfLQ/eiNsmLiuBfUG7+zxW5tWJ6BGi1Z2xUVmO3TXe1DSTsYbWBZR22G
VqWH1Zpm+XjTarDq9JyLpx1CgtUYX04pz89aRdH+ZMxCx3OSPaNhrYhpKIGS6W0S
yWFxr7JTZvpSrwBV5c+5BtQkami2Lptq8waJauAWtEEmKGPXMChJDPgWh1UGb5Sb
mx5Ledj2SCSywrJIzDPNAGdIujJVxDQSqk4lx82e2iX5Fe7Y6d4JsqvE1KrTiSBH
7CKhq3VtYEVZbtxemKpuvWjeeI4GUdYgK0Dds8mVIUywzu/vSTvM30uIA5fN7aeZ
rjuPPCWDb+IAYtX+iik2Z/LUSzbfApxeegqAmTC8R5EiNrKCEpar0QcZOCX/XL76
eM3XnKUdEUD6hppjTCIW/GaYIjr1PekJtusKIz/7I/vr+1c/rJCnz8xFfNmHFBBO
chl+T96cTEcSYLKFpp+Q8tuW4EYlWrUHCwRqSCvd+FQKEFZFaqVG50qIMjXIXv5p
b8596Xo+d77h5gAI3ch1fD+fp/N083uh4eaH5SdDkc2uP/wJKXyW7X2UXZw410HY
d/it96i0UzoOoPzJ1e4i0wpwj1zA/xxnzuLfyxBroiqM/U+h2P1fXTJq8tuxfiAY
cqyV7Zwm84QKDQzGvLvkEKtgIY1fopJIfJ3Cm12/kmkGZolSCzjlVHb5hNE7mYLg
EFGCMG5GPxP272SBBB1XAj2Gnb0K9ruJGZpPANUIfmy3WQgIX5rcwCJQUXjGyot5
ibaeQ73TSwJSB66dGUYTj7Z/qjy0IYzfZMzb+kZQFYnowpFn4zFbAVDqy7YroDrG
4wFDd17vaU2XS6FuV80kgxCNiHzDYjQCN5VUIxZ3+CuQ054dC3MHxiHLLsXfER22
BqGIGdMvj7K/4yuwEyvOsHR8hOtOwYapP7iiYA6Zw2A3ewEveQQmG6IvuzApFNOP
9cQJm3iz9l5lzsAfYEf8YbFtciU83pWe5e77OKdZeii0iSYv5GiDRGVJ+gAOrbn3
nGVSEozEZ03r/zG3GVEp1kDYLFlAXPUwhPxCS0ne2H8Y3QJxUlMW/NSZB69NyaJc
+4KAwYS16e+ZO83z7vdP0Xyj0YSoTepqXgmmFfve0uwVIZb/vwvGEUMIuGdrK1y8
ol6N1MnMxyAacdO6oLUaIaXkoWOI4yOs+urBzwvcfDHIVuzELVPl244s0wBrzRau
r0jCXUPtJ7994fCrO2M11fm3yuaHbgYz3LknvBGJV0ZQUc79X4QTQIxE5sRwIUzt
YFybtfYgEeUo9/LYiY+qkHaESIH29wLEjTxNor9/XRKmLmScw6JlE54+avQrY3Zu
W3qJz4+LMQL6pybQcpTnN2R1mym3QM7FH0LcIYVSaElXoMG4uZV6FPEnqGy6BrgZ
aP+qEZ9SZpTELIA3OvYiOqarhWLywHc66U3h2f21wp4AQDcpo1AJx84JN3t77/Aj
A2I8UQL/4pwiy30YIvwCTUzgd+78vAU56ybu0S9zTEpYK7TpqPeVOvmI4K4yQ/SF
wDI8HZTm9WL97POUqc8TUPRG4h4kt6558bamqUzkekef3IZP6NtOLnw96+jHMXh/
DW4OGZXOjV7KaN9R1nhcqkNm1bH7xG8N0CZjf7um8A8ku4MsgEr9NHf2NnAEeSdx
LRTdE+HYBuM5UcPI/xS7ZHP+4X3CfB8vMlCaNOSr6SBkne4jUinPHtdtu2yeTfPk
pBjL46la+Kw1vhKpMV1vAgNIphG1aZNQIx/T8o8pho3I7wnpF3H+Zvi/IgQiNRa7
`protect END_PROTECTED
