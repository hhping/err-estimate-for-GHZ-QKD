`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zefjlhRVmYj41N75fSlRzGzHEZZu69ggr9Jp+9b/fw1XBDq8uT9MHtCtb5544xg5
TeLQVthWleD0gewFzWqJ3VIXBBAOL3zOOmSmaQdKAWpTsvCWPea+jF8XVVLveKMu
PDvKqmpt7JwowiAFmHWU+0ldhPBtfxSDi6yrgzfk3xhsXU6cIqqIila58uYustRA
saANdvojXwgR3eh+79N5Th4TuiiN0pU4sz+5tnS8RZnaVoNr6AtpLy4KQlo2r6W1
HZcDWVAIZsz3JwedQbpsPmVnQMr3iKwil6Gii4yCQWvh3sU+NsQUWm9zljH4Xs2w
yX97dmG8rqDTCqFNFbBsG6HGxdAqeVDgvjkjptxOHe3SehWupb7sp/2Up1d6GtoU
uADz1WXPMkYwK+hyjc+dcIoUs0J7wjZ/BnWddgEysCT/oF1eb09BcL1gaPXNMZiS
+LgxGct63L/7s6u+ubiN4Mee6nGjjClBrb0g7hAwvsEUt4X/l/JgyCCE2yzsZy+E
TN4XsfZfRky6qOSigD1+hcDcVLJ1kyanhn1VeCbp0KoqaRPGguQPITJQDWjKs+Lr
+lMstQcHNT7jDNmRFuI5EP39MnqM3kEYiiAxQRoTsuQXJ5wa3AlG0HBq4sDr7PTm
hxvoAAhTdw1xFcN2T3yBR5xeDodFXWbMGJko+s9AmaJp3LwZFxxG7fHX4ODP/NI+
qCQebKTXzRm6QzX1+XYVl2TLVsJgqD3iPPMjhDLk5WLV3rrdFUxsDMuaPS8cPEsA
8opBggK2Fg/W9c/u3QTMbE711c9yn1JhMozgK2vgE0seBFPVBKcy8lmNBzkuMQI8
BbffuQKnOv3QCBqRbz7rj4rmjzPWfan7mEj/03NdhYYSDH4AsKbjz/VD0IEQyaQx
g2AmCLYZuOnt+yCXGkiXs1k9Rw0++fli4dhwFhj2QDlP/2gJyA0RkpjnqQ/YS/8G
msv7Qr+9M2JjBNz2m8thSDNHrk9jNLdXZk/PS7YXa09DgCT6OyX9lndiONwwrqdB
8f8R/7f+ppGdyTiy2K2Np1bWkByNj6KImOj9bZJXTbj0+wXjVTiv3vFG1wnMFLOj
ykNj2ahpWTOn9PU2u6R9Oy6nWHHVVc90+QTHATMPe7PlYsj5Q4CZi412pAhy8LFy
wj/y83Ky9veqni9mME0ZmNulNWKPVmJIY8k2x0GPKmdZUkM1HZL5kW003nBOd9mV
pRmL/uZlZgmaKEqgVfVyoyhpbkuYpFrHIqYzMqipnCjBiuWqv7OjrCGcAZpRL9s/
YTCY4uJJENrT+h5lQGheTck4YQ/UfvFQjCHA16YGk9Pwu19Oy0Xvfcn8Zb3AhSxc
efQ+BQ2fQK4DxFCoymIQL1nl9Pv+jWObnkLf+Xsj7621CK+mdMB07fcxGPBDbRjP
UklmHRNUIexfabn2VT6/s2usCjZIEAgh/M3K0POC/0D1nq+nNsuGu8OYmN/g+H77
ovR1WRg/gxKpUCtH7q4F1vXmRy0kRKHUoAhpl4pD4m/P4ExThHP38oDOVPzBovAu
LKPOfS+JrSEHCTAt++HtEtwtn0QEuLUfmW3tK59jMNhEbFGL71aq/h7tqaAi+vTK
DLehPDqrbsxV5ztxvdQ9IiUC/pwv6BUBDosgXeel4Pu8e9GVDKxRhbdLRTPp3M8+
SWumptShPUnYCSFwp0d2MgS/stYvTPssRkLsKLzvlV4XhNPWkh/OxzM3fguTpF5z
/M6Sn6yWZRv+6q+JR2uZoMFdnPMZtJDLx2C/0ZeSJOzqznniG/bQCHjOxHwI6rlA
NdhVqGSFfZXkaoZshC4kM83qUs1dQ2NpRNRGR8XhMqyovA9WK2RpYGCAC+gmuuG1
i86SiAjDjpn+tv+vUmtHR5tyTwP5WPyw7Mji9xEgv7/hvIDklRSNUrdVGRL6w1WD
peP8R2X8fcU4hxEU28Wz59tpQzF56Xr0++Wgj8wSJMBJ/6fBFQZoogrs1yekO6pJ
MJrGZJqb2sAeejxRBal+2nrNIdM7BI90PjH+GqdmCn0DT1g7xMZtVZZlqStL+JqV
k8lJLESnm5gS9SCPRbPJvFda+pexlhov3lpK0We3s9SsngQaZNl5nqfickngf6HB
ienw5PeKV2yif8nwxGoKz5QUuqPOoVbg+MP1OUw4FpYAzJvO8NMFcYwGJ0evp85R
`protect END_PROTECTED
