`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mR+1Gc+KOHS2ehQ89HSti+YuvWZw/LN10M/MlgpG7SY9DVOjfeihMnyQ/A+0EPks
oPjtTUhNhF5wDZM0f1bOROf8U2htaG3svLNOEmDEtfro1aF4SqAiDOYQKk8fuAjd
JovgVZlExOGBBMemlDScRUPVWth7Y5ohfFXgdvJXugj2jq++SSElZuetS75em6c+
3unnXf2sY6hZhqHJpH8NzjkIb+UM2kj/LtBzBNPy2WLDwz81QhlKRbZih7zfy+07
cCkUDFxVt7xSzUM62pRdULCcCXHbHlaElsU6iGUHaV3/HdpkC/emGm0+kNmzJ/to
bi2+ItJe9X0uRMZpYVqOMDZlJpV87N3Igah34EijLDPx0gMla/bb9t4UNokMOn6J
xx3unIFKxVro693ZDbXW9Cn7xAdT5ndAjsfxLPCal2/YOVc2I2qp3OdTahd8x+uA
HQ33PHGtmNwp7ZENHYT/CghTseoWDa6+FwB8IoF4VNtbrNzYajEcUf7EolcgkjYd
gOjNAfJ3BC+d+c4/IVtke0oKQVaOSLe1dD86ncW+0lh5KOcpQcrst4S6QcD5Ir1U
7nHNtUzwY49uI/yJN7l+TI1MfRyzsR6IKkNVnWl2WiZtGPNuewFTlwdGyVGuFhru
de9sqviIgkXCUpLEJCLvvqnJMtXkMPn2Rp0bjxVBofwLHrsK8vcu1IQRNAf0rMGk
9GR3mFYlCwTsOeJAITvss6kxMiP8C88JXaVHKeTtte/tbsukTGZmAz9uZWRlgoCU
DXs3EhgyBDWTiv8KakZxQpeVJxprMaviFXbWPRgUhLg6L7R0oS57s6wZWaWqCICi
G06NiqkPZTK+sj4BFVs90WQpKTy1EXBBhRwpkHjtn0YH7+1JJ0ErPTzPX2wN/za4
j7pa/NuL06R6IkjEx8YrKumiSHXSLFOeyn4JsgAMLNRm1uBt9ux9vGwgonstAVdx
v3Cudb9b7hl+bPZULGprgEUB32BQ6BkU4lYQLn6PLUdkSgcbwuUyIPEm9dC8YRI2
hp9zhZcQ4MRw/4Fx6guH+ukUDkKNBiGHk/++MvvzqqEXWhYaSOJ24qtWmNQvZBYr
pRVQGpeVJH1LrNlr0Dvs78N9vQpXx1ky1RaRDRmriez8W4lfoYiVzznXrdwvNSTe
IDZnV+Ad6YaHJ1aTryGCRpggvPG9aXbZ/2K2lQSBGM4=
`protect END_PROTECTED
