`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/CjlfUiOwGEJnZz0Hvx0LQNRdC/PjU14zY/akanpbibQ5Tds0hw9Rz2U0C9JnR+X
UJ/dUX/kPNe9OZ8ByvoWIa7+Wq4RbI54WoOl+7gt7S56GgoQKb2OT3cIqF52S5iL
gPCFt2vecEn5rPFIJoUfb/JtJQ87hGDDfTxUi7jx9Eepa9/R8hYh6Yr+P9XAoH5G
K2MSW7Yx+tW4ViB8zMuIjQ3o7+w7wV4AgrED3/+VQzJUVJGw1+C9bzizPXrS3HfN
YSvtl0rZdvuObdtcPxfL/kXE2+YtqrZ9PlpAaMfIxeMIIcZbMi4i9aBVHjhKgzcn
xwxKnYHZCY21MUWuAk8k04PAV7ZPRHuh/HQF71KNYLjM/dpZ3IpRM4XvVOieW5jJ
2fKumJ/WB5iGI9Agyc29oz+CXXJEaN96crmuIo2puQh2F1qeR9ieVqTvtJQToZPx
xWh/Mg4RNlv7W23UYYRJU3G5H13qA+6W6CocvFRRouGs50JiYlMfNSud1DQZuerN
d7AHhwZucOtigd14PyQ20sPW4tuYdQTtljO43HIp9xnZirHPSvxhVG6Q+aW0pK21
3PopDt3AKzV3lC4aFKbj0NZ6UPUEjbvEkfgrMzSfL88eepNLhbBXNNiSmqEzSzhQ
pvnu8rP2JSrGuuE5qGC2+9GnRyyn3wTj3zBpOK86OWi9vEKSUTGvQd923BTHt4KO
YHr85S/eDajFkB2B5PISXAnb+AV4OlCeA5SBPddV4X7DBPFsCj85cYQ4A18Vn9nT
jPt23bI6LlyGUETxmMzrVjHva7//jndgo+f1RHZshOgld45otl6aYoQByjPoRAq5
D/XJtuZ69hKGqkpX3yG7jKIY2Rs4BXm7ruG1W0WQq1RE2qFarCU7PpnOAixLExJX
YE7GAwY73CgmPvuUgDQPAiBAaKYwrCCrH13S7NlSrsNUbk25qiOeT4DrmRkBYdFk
6DtOJNvvkAU8HEnaX5Y0eI9qrC7xrPBU8W0PGjHiEflsXmADa4ZVC3GZJpneGtay
LO/O+zi7LiRD7PbH43jazhyFHm5KxOC9OFmH8xzfyyCtv36aWDkaJjbmzDOWFS9J
KCb42wHUbT2AdlmVS5B8PoxWHZyeiQAgxBSgxBWsQFJUjggW99KfnqghdJ6k8UzV
lMPnAyDdZ5bMh5pAx6M6aWwsMuejfQ4dL54S+we8x/EpNFXiWj5kVll0e9dhb/+N
OTORhHdNmi42tN55yrdiebxeC99HPV3K+6a+lL83VzgSL8JZhe7LM0+zUBYo4G9x
/mcZ7vmY068RBOs45w4tMGFvd3ha85bxCo3ZxhIqT8PKCLV/Bf+fbUfF1wvU13eO
pOfHANQf1HUbndELUAFM/SR3B5Mvm1/T8BSqy0+kBUAWglEESUb1Rt3kf3e71u69
rmKUgBkv4BUMaCbXhvY8Ef4FvmHwTMfGNH61R2WZw3wQdI8UWNH76ys5aeZaRtSc
6sMfQL+UAdINMAsKNEG4BvnnVj5dlg2r/BnYdiq17sb7R8mUE+BMFbjL04u5bbqQ
//xmeKXMqEt2tNMQNTbYWxfja1BPnkhfCBF063AVpzfxg6rRy7J89wvQLrPzkaUv
xutljbKrowLqF1/dCXftNNBqGtw5YPf9h036K9jf0PQ4NOzWGn1qxugt1DrWdTSx
VAFTIYt/GZp6+7OKB9IGxywOZc4XSyE9EP5Q2tfQgGWqygkbDwMBYWVlF5hwL12m
iFAEwmLOz4USNZZ+7r7chqLxo2UiIUGKWfEDrSYPnfBWi0/cxkRQHnppoR2Sm78m
+bxI5AjADxM/OzF3SHjqU/MbcBwOEou5OZaOvkIrdIv5m4DFs1GyYXdoLonhT/0e
LTQ3Z2yoztVfdZH6woiaayunWPy6VeJ+/l5CINScspPdKTxIGx0qeAyHWY+rqjum
X2yhDvwSdQyXy4VNcZY2s+d/wTdbrG6mHdPaHd2Nhb3baPtPWSm9z92eEmZhcw5c
HFnD1V1O5JLn0P4UH9qMRhoXstJ+p4lE8uTFr5NLyMGbf7YULqA8Q+gIE2u3g5Sj
F6CgVyq5u8KQhOXLmp3Ye2JOobqXDsImZuFRvA5ZL8ngJfdPdHGmNzEJa+hvGIEs
KqtO3XOL2U4fIvMQkVNTtZD1le6I3mjfWkvMkHFJUld6giDl3pJ3SkUmXv2DwIXF
d87tPso+o6XDVbk83wK+3bss513jg+9DY+Pg8RFnUBPLZjVo3wHYv7Co0gDMI+XW
LNWhLE2jEJqSBonqhGBJb7Wtcz6JLXaRU9UDgorxBDXukdvTHQYivFLZuPVUNn14
9OYuIwhQEPssa2oEFN6V2ikzrue55PFTkAQptFCvilCM6xN82q0ixaGAidN4pLt+
/VpYYGFgECAdtQL0HJagTQ+9WllgFDhGeXW8fSb6XrOuwkLWyQSwElJOm1DOfJbl
wxTgRnZgVeJ6brg7yaFWPc1CH0EGWv8kUlFq29bfEQ8SGol+nbrSIprvmlni51cd
Ld7/Bpo7ZzAbb7xMSnVQOEt89g+D1uUQylauaJOGuPJ1wYrwdUmYem83uTv+eJ0C
odF7xeXl4AIcIU8SIAjDeQoJbBkgd3gp3wilmOjtorVtrq0oZLWWhO1W7B3aZA+s
mGPskc7qNLJEtjR0rdKHTb0s+RHBDQq+kz4VhbvgJgiFnSlh9OzxTk0RG7ZCBfBb
/L7bZDS688UeAPBb+fDT6tNutSP1nt+AIH20CTPNT6utAnAoEWAHIq8ZQVi3c5Nj
durJW+4JoXxSrDJo9kvL2tyUTBye5/LDrA1SE/JCoCLtvCzUyeE6uqPXp1okI84t
o8tUDJ4l0nj2jto8DckhY1OE45wbxO++HAJP/PfoXmNk42v4WT5CrIQtSMABnSPA
KxY1hanI9K3gzRCTqHn3fTyBfPj9ExJcqx178XgkOdIAJx9LZoIwWJ/dGe2OgAGV
FJte1ZdY9HZWtUzmsx+SD5/BzLGE4KfVWBNS1+Uu6tbVkRIsCgGKaxGu82wmEhrU
HL8AgGd5gXEWuoZD37iPG9NHLuFR4O9GcN5/Cii+exDkUXFFuYNd6FoXDqCGLmyY
jkDjsXOrzi1b+m6XrUxdzg==
`protect END_PROTECTED
