`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BrV5UHC/woFWwf9f3qpSHfb0oxKU7pTcXk0xDoDDAJ4ngozpFAJvM6S5F5erfQnf
kWJsHdeZUmSO1J0cjKm1GvzBN9krcj6G1BDe2P0AdDXr5CMOkweVx6YMsDQONErU
2Y1OsL21r75TzYsnZPczhRVNRQqDX904FmrKGaykwBjteUqLCRJBywTZlmqGZaFN
cqoKBY8ag2ObTQSWATj8Ol5fm2i1GW3rijMdy1wAjVO/3VJOJr+ffPWy452IZ1nY
F+2vxX6YEf09XzYzYovyCvGHWFzSqipyY39HYh6ViKQgTPbO6jhqqFMujxDO6L5X
XwL7gisxJj1/dcrzs69u+Nnfqk+5m5ooQ2hCTQBIJJfBTPZ9YJ3Ck3+i27dyPxzn
TN78AtVhoFvX4jwZQKlB6ppy+42PBYFu6OcwWRWwS2aFnNAvV4vcG7t3wqBvttzr
POLeS9vYKvKiFocMJ7zs3D1mr8KzjLSWs6fYUwtAtfhgP6HlYBBzaOc3MKo+/nAd
CIy6SnPJCvBBHSupPlY31GTwOQ/USgW9n6VlXh2+KCzJsL7nEni+lCrFVQL8lOoz
MBdZxA82L4l+o3yVxcuSsgWzTnXpAv1Sh7D7ow5O6cNj9IG5NlHnlYE6rKWxi/aB
+91ihCRUL1aJhrWLpEe/EuG9uwP1ZyozAxJdqFSFnZYsx/ERxnXjcIQtoW//RwLK
TZnnKx7d+VyTMJR3rxxNMulhmPXfrZLJifKIAhjcQHI2iPeBDLUIeUdTSohZklZu
NnUHWd/k1oYGD0TA8RMcywT1qXpZlhfmMlNKD8iBufUFQmj1gnX65OfGaomuxmQF
bjn2jMO3vypoB1qVnwKoRhW3r9xZ7lyWqg48Sriaw6Otc0q83tGq3vGLpWTiY+1e
`protect END_PROTECTED
