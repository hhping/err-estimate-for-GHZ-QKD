`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNkWuXNauIQbiwkuJHcdTjFb7jd0AiNPyXJ9+Z6iifC8BusWVbvog2Q4SHz8LBD1
eqizqjNV+NkSz05uPknELCgis7/ma9MTOXP4qNzTB01gb/wMpvt2kSkhoMLI6LqI
2NivtRd0WMXYoCKgb5bk4hlfPcW/r87l7ikdPEYFh68c2zkiD5Fu50jdJFIB1Qge
zjf07F70s4CnDLf78A4hlKjDM47WGYacdn5D93nfvo5XFmvyz0ZwU6sRB9c5hRF2
am4B6uXbWhA8a6WPTpx9UL3k0EBpOjQZfBLPxw+xLIMuHO0C9OwMWbv+d6n2GAYA
VSqZitg4vGz501AxkJsholqMW0wqGWAftnBl6Q8Q8HTzcj1Kd/tqv8T7ed6ljcW0
oljM9ylHBnmZFGN3y9/uJ/9Y/Y5zoLo8mkvuVOUbgd5kyMGOokdEj+1nH3BPDC/6
raA8AdNd5kADLYBe+bO3oUbsqvQ19AciQKNZ3jVQTmY4F3inTv5htmhZKqzrHZ4F
psLpIAEYTCIH2MErkw+utAGMLx29PzIU2O7SO3JFwZOBH6fyJ1FJbXiFP83YR1Ji
mEaaIXjriBQBzsjr5cky9dp3PxelFyWuay2ydO7OpfSzFgW9XEahAE92LBfLNQov
4v0PxG1KMqNDbzTrlqHMukxgHY/Wd37IBq918wPZ53yJmvDE+V8XgIST7xV5LWAj
5ZU5qVZvb+VRJiqxNuS+rEGYZsR6iLzo4Qp27TUd26AbunG51MpGPcRMG64Q3t/H
0wgvyGBYsZ5PB4EpJaIiCObmf4lpzMhddqaR3l1PYD5CJ6Yb/fSt/K14qS9kreAK
tV2oGzjlSk9PlifWVlQZStm/QgJY6JUi0LRPwXt4qzwBvYHy2WNF5Da6jSdEpGdl
eROi2oYmIceLq4D6Rc6bea3X6tfTNFuSSSox91+3XAsqccqBaG/GKHeBcei5y5JZ
bIOmMSS7SBNJzoe3hYGKM7lcgeu39VHt+jBNTIxRgsBOMWMHw4Zo3CJS/jEZUhCm
Y+KaY/5xVPKLHtWG0MzNzva/YfbHMBPsWzLNaKHwHMe3HlLJEPxcmVj2ZjLKXiaa
UGi3VnGAj9KKMJCSXBXEMB0NryrcALOfLC3D84KAYc/3mSVSN259QynqaVZxXZaY
zU7aAGeM8jaAYdTtQ6ZENUWb8PzU9hXur5PinDYzmdYVRwj/EDuTRA7Z/fvVVVqp
Qd3dgt7aFhM+qjcpp7hV2L9XVOKmm99VYegXt2XvMzLh309dr96Xv0dPxCAMy/Fa
aS7m2gXMYPDa6aQ1EPPtJ9Ke30PrznqxRF6aALVXahq8pt9nOKxuPLPzQ34K41dF
k5eKVdNb5Ovw4wd4f+AvEA==
`protect END_PROTECTED
