`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bjM+wIjJWqb7vZWosC5LPOIh2UcMuvxTpaFSwbw0obQAEr+zJK/TiNbzv7Hc8vXp
Ydh7HLSFhRiNy+XYcYfOW2YuEBGIWfmqKPWvK3WMjGTh/WtSYX8SIJ7Wa4tF9454
LIfbK9fBMbuy3cOgXYtZ/60xfX+hG3WZMpqB+G6yCj0jtuRLd47rzT3QV50lkJvi
xGQbWcmQCB4YIAIfqlIGZFtGj1POw09jQG2RqdM8DgunMCWG/CtIs6LiRjJGIWaI
H1aq0RAZi+QxGyZ8I7yZiz95UURYRCjgOSiDl8ljHfGCNyx6Vzz4AW8g5Kkubgh4
KrDpfym42aY5h+6mfPueXi9SHHW+ykdcg4bFaIzFIcnL58v+xJLNSgt9FMaUXWT8
Aov9k4bLEYaS76F54wDo5kHA3tseYzQgxBe12X47TmbW5OElELAiIiInCzMBkh1e
nrZVfLYcjycdT/7w7EQCwcnMq7yuRK8x9mDOQ9ELLuD6owTC0nsHN7RiAjjo3nn5
uPCQKJLNIpY3iouwxdNSAVQ3JWv+iOLx97SYAKwVwqziCAr63Ojwaf7uE5unVGtI
vOnZrlriYn9IilS/IhMmTIlAYTv1fRNpTGQG99Uu80VX1BO6LK/IE9QxUgIcEnjh
vdqC6Km2fiQnxkUoQ6YMlrtuk/vnzUyjLh7g2D92ZxzXctuv9C5cHc3Nx2/8PgnB
hRbsfninPffy0c2cKX6jOYIbU5DH9ZPvn+isOcwx0nlCnFhplD0/CgNS65tSr2Zb
3EsykOGekZ0m8PWcbtMCBvaLVOW9/dR3dATo+zQ3Wm5WkeolHY7oBi1y+pvqbD3z
hGmPgJQkP32RTAWlyz69yWcWN7PP4zsVd1xCeohbuKVgb1hqv9ed/Kfb14OjLXSV
NCqD/PcUJSqXfxIHG4pCRFaLpcVpJl/htqTTcVxqB2eNARZq7g5rPd5Czhzaa4gC
cFFe/W6TF36wRFEpVQztRT17lmPMduCNRSUh52zm+e/TbBA8HLuKPe79+eSlhA9c
fkYBaaLFsIYL3LSRTHZNNhS+Ad3mlapWODFuOsr2I20WlfeySUNsH8ylHks6SP1I
BZ4TSP+CG6l9yyBMsDOlj45jxumJIdxzhbLSJxZh67CQnEIurkDnN7fUYGQWWNLk
e8rwptZOu/6Uos5vjbvDpPT6I8DSqkNcKvgaESyxFvHI5r3pgcTfiEh0l89ACdxy
l9m+cfOfDg3uunBgcmvCJe3JZWvieMbzAnIGrTG40M8=
`protect END_PROTECTED
