`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qglL4k39zwBUKPYXska+Dfge7Iz4o/VLdSXXfHs5KnHnV4yUppdqBO+k5qnzhM48
53BHalBumIiSzvvHq9o3hKra8A4JgoZt3f0OZPID+/Qk7Q89TVskuVZqTZxNgOh9
8Cer0lcbdqu8+qZQt5KZrjCECPxAtCtf4TgAzdtXrnvaoeiXZLqFhavF51IZUqZd
9ghw0Ax2+yA/Zaq3RlTxPoZYdxsviFgLJfeLhWXpq9t8tMsHIJ0UZKle+Ve+8VuJ
hyrszVWgqWibda9dico4BFO3N94UjOADQAA8m+r/HpCbCHy9RRtUo6/M6bDV+d8+
RICAqakjyDKq1MH6wqwvn1+F7jQ8ipyr32/qHMxZCQJ9ji7ECJCbfvBcNLwch4i+
UdB3/3MgEyG5SI8BWsd9aqpXe4KA0KwjCINoghrNW69qOnXLaJ06jmZ45tgNSg0J
7ni57spVEFmXo8YVV1J/tCrYEf+8G+IuwctWXdOpxBvOkusbjCWkEdn8B2c3JaFc
FmafM596MlhUFvpXszB5/Q6BLFwWYNqT6/SsQQUi8LjeCsjIvzw4FOnm4HSD2EzE
rf2LTdJA05fDiBg4DVuMrPNyxfNcCI8LM64SNIJNWrctS/pzUGStcSt3baJXQPVO
V4XqUOhrNNL3MFf60+sNAuM0kEpHPHeJAzgRWJqMgR4l+zdZ+QKUqygGOutrsIKx
wMJ9BILT7kG/OvsuMfzwE26LtkDXJCHJuV+9ywFofJtjej/lP6eCyVubYZCyBKO7
ubAFw4gnrwl67uD6WCeoB0o/4JVMvXmDg6RAvHnHQmDvVTKrbb9UWEni1qodZ2ko
0RMvyzODzHot47+TxllXuCVvMMZGDwb0kkQKwRQyh8WjnnVPQGVUZUYRu9dZWVjN
y94lvaw093wTfH4NTJP91U8S2u6zDOaJBcR0h0k6vt7NdaBTa9advE51QqAT8htW
P88ZZ0fU6Zaj02S8tY2Go05Shv3vay0sFNfuzPupBhVzT3yx4Rfy5uwIApzllfFm
BQsdEUzcWTDglg4UZqZSarPigIXP5ppJ7GoPxZutdzVYBtaHb7vz9BXSkS7A44Bo
ayc2OQ+toDsylRsAoU0a1Hueq3LB7L2G6QjGX545aBAN6g6pX66h6xrdANnMxr64
+eYFILXc1AHfSG3kCMFUCsYeJmXLbfe6JuOdpyPvM+TtcrI7+cKnL6bffoPLHGwi
68UveTYHu5kdTw5QixXOOkRreqhr6RwXAumC43AzcJZ9O19mRjEp7BaUeJYzNIIA
jOZjTR8SsaZwfYCRsDmaoj0IBdGeEkFE8h8FpPqDtQI=
`protect END_PROTECTED
