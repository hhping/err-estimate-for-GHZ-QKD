`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WW7lwElLD6CRY6a6NIC0PWPRrsLc7K3QwDOgOv9YXSaA9H+YIhUgYOfnWJ2SyDaa
uZWNuzLp9P9+GS0C6efz1ExWMO0WDuASHhCWSPiQQacfDb7F0xVaQA1JKzrHtLow
Xz2CFrmcRmPVmk1WMAPo8wX55OzdmDjFWy+PoKHjiJXDxD/+1f5Q1hPP+uOjZ3Ov
sLKGQbvuEnrOFpk7UzbcYaE0iErkCNEJDLM1Bt2gTh2XRmebbDcqJhlgQ3FIwHJr
1TLbyHAZlHptgTQJ2TUzEcSlp+u4SC2QWjZqCKTmWVElrhyuofXINuc/jkDGXiht
8MoPhaNRVGnl50M+bd02CbyLzVwgU4bGg+tMdwikdxlFV1kGo+g6Rj13CfxKQCZd
f9eS9eAbdZ34CANjKujWvOjzkJr8fGfuUAcigXqVP03YjUe+IUnGxF6NqJsiKgkF
zHdr5Ef2w+Z8iwxU3DAvfElncgQuHs8FPEfQ0N13hOAe4o4C1uBxnzVQSLcbM/8Z
fdtEEPrp99pFD9CPIEdn7aKaWoQL2o+S9xxDz/sIQDHxIPhDU9SXvRLCBcsVeEn8
rSIGff1HTcRd3F73+gAViqAxXPwN6nt700xD/rVWsP7+ncFDPWCNi6RFmIa5PctY
ArRp8Zn/TyABGtAgGPKTeGzdCuxr88ZPnzoMlxuD9aNGDK9KNhqFXOCUSdIbmDIu
hAHDjDE2IL9PbUcsIaHiAmU881fPsQSrJjLn3VLFriepPylQXL5S4qmyPhCK+8A4
X3brEhf92XhVz+dWYcRDtX4ee3rUYhFL47C7FDpwD2Si16/1sNTtOOUdgCPpumFL
3rCtdsG6//7RDqGVsws+MY5KiMh1UBJCy0hSpvOQ+/PaW7ueMBT2BMUl6Grx2AIe
Xz0hdk3OCGW7eKY+zqAkOlQDK/JvDEiQzb97HYBW/wqrxojt9SBdJxK1ku2ZttR6
+PTsr7GElft3TepjMlw8eGUcU4UuyNmUk9ZAkQtUzcFeH8Lp1hy/K1reiMI/f4+U
dWyw/FyZIW6zR0EtvOfd+Mqcj9zBGTydvcHrA7pPl6nDy9NxayIwsRmzGxDD8ZAe
CWdqLrZQqW82xAdZz8PujVivU9L0LjvXl0c0e55x/dVqM7yF2g5EKmuHMnQ0/bB2
BqgbAi62VUP5BVYklfLubtoz6BlDpD3KqoLPtkEGOLQe7ASIXWo2nn4UjGMWb5ms
y/1oTr2SC3h8/sw6szYF9psutcIO3w+PP/Yy8Besk+XiJD/Ko9tce9ebccbyMm5N
cLWQs9n+kksh4gK/4pAodzA0CsabafzBRfXYn47Pgz3Kt7LIprJqopn+LXdIS3nR
YDUVK3KXqoLSZEbeKnKwp1BzydP/UyiJCl1mR5pJYNsOx221Oo9ZRotBBeQ2TADj
BItbMePolokPJWqnkUn95b705k7HPw3OrPEn8Mg854gqnD4piI+2atJhtE/i2Oht
glkrWpd2oqjyB7Od0quaaa127Md2Kma1j+L3jMkZ2RH9sO1WPmDuuaJQnj8UYVvn
U+EnRwLRioNk/FZmG+GowY23qM0y1YDAn9XGF6OwGzPUngYY532Yuuc1al1aF5DE
ATFbCnXk+Pt1KsJ7qGwcyzzfjmhIyLYQ1Ujo0ZrYeL/dstB8KViSXArKPhifgpDx
ZJjImpMqA5AHygWQg3ckNNd2phaMFPxs5OxVpauWEcvgjTQC+exwDFA2j55ETxOZ
8l5T5uc/x2ODx2IX7DxOjmbHfaEYk6GdbvYZiMfJX+/EdyXcuTrBwnIKww7uoRrQ
kTtWsXMFOugc+7wmr130SNdlqZrZq4kImcXrOiVpT2ja51b2ANd75bFhByyX83Mq
7tdIUIaBXzzN/M0zoK1s9zntMstwkSa4aJ+40/THlF0IvoZaYW2D/IWxIReSlqR7
N7RGrGaYYx1g2ph9kGH5FwDFHNco0SiUW1uJYpWUIWrLpwCJUtXvSAQ7dcT0UfYl
jNKk5VYoVhNMdXpRiNJ2g6yMkzHacj7NDixgpKugHu91P/8zoH52LGj8fy9X+fvp
/6WONMc95qh4O9GBoMPyYbJ1ePsEiBTxmoMpCjc2/IVvqXyeHN+VS39hoXCLEuRm
T2E92J8nWkJcR9Og2bFZAFWbU/oTPvWEI97VCqO6S60iT/vApfD0CXHmcC2fChr7
51ThzSz6J0H3l4sxPpHRyq9VqKiUxViyd9YArTwz9l27CE8uj0D8KTGJ5aAdg2Dh
JyuI0BjSqlm5edAb3AkxiCTTeENs2kFoE1Y/ZsSXqfEjstMU2Q8M4TvP7NuUTtqX
li20cD/RRBW00oV+QETvAf6wiurMbGKOFrun34fT39sxmJrnbocw05EkBaIkcy2r
JmPVHc8iFTGhAdLOJpLYOFMLhOHboDn6bqwHRBz8nb5/32tzZnsIV7EyrG7WYJ7e
107MpmKL4ANmPmMNkxPfR3Dv2UfbuA2ZXlxdGBOLho1WQJA9zlnH1WGQd4vaKvpB
dwAIqeoMHBIa6zVU2YVSM2cTN0PZIfkKPIM4v5YbrcbIF01vAoLa0TLnQJTRGeZ9
fApArsgePyMpIEPmvAcxcSzhJg/ICPa8n7qUoC4tCqSmN+LykNhrkXzZZhI5KWiI
hym5ycxZhiUHeuobiD+aFTsFQhZI5YUy53Q/QX5QcPkvnOUmKPZ7H9mP/xYEJS9P
TsfD8ve2jXoDZD6QzoLz/Fu3HR40dT0GyShDdJ2U6CaPD8gKEhl4N1o5m+ayP2lo
5dlhCyog3Ouj9/rQQ0Oi09V/6KlzCd8Q+YDH3ez2WNhlLRUYbI1uXhedGBs6XZR6
9+xeYmyQ1feYJkVWe6YbLWw+CS8MNfzWR6PZgS60uDMsPOqINOteaK4vKhLFIf56
QdxzGn0aTHN1Hg4oPqhYMawbcsjMSL7HigAS6pPO0IJLA5Srty6Aw5DtdT6dw2aX
X/1rxP0EKB+UmTObX7OIvwuHtltnQQMI4UmuxKtfoUhOIq25NqDTy7PaaIBabR4I
Arg/V9jDqyR70sw/XKJ4wICHiUCtBM1wBMYuowOfZNjHMX6Gr1ShBZGBtron81SL
bP3X+GhKToY5Xx0Ptmp1T9gC+/0ZYwmOZyzu+Dj3alx9MWjY8ovC38WyHDEHLPvc
lUwEb6cShGVZY3jr0aOlNlOu+//XogprqlXNyWOYWXQZFs34yfCQidKPryZ1COp3
0PvBDLo4VxqKsUPLA7dCyDZkUOBH6VnwF2KLOL9lxpSNB8NTHDwjV+NUiYTo0BbO
W7Uza0ugXHb6sXSFj0i1OHu/l8FJ/Zb75Gfk4OLXM8o72MJXQNIjWQnmbWX4Fv51
zoJDGBy62vEgc7ZrIjyLIH1xizKD9ymuKLQY1cJCujx4moJaDjYcHe6IEgP6vRCT
SFMCCTwuGg9rZD7lzIZYe7FR0a+WoJOE+X1DqCyxkta9DUjucq8nrVHpGYuhMEtn
RFgsyABOK1QORYaoOiPeFMC08XL8bnvUAVevQjtqItQY1Ietn3yzMmJMXkcRYgfD
23OtSX/iFqgCVSv4y99NjY8qDp/E7ZS0uNCtg7wwuwqFww6LRf7Xetyj6ZN9PPuw
oBr2JfOA933Qg/vY94npZxRmvmgHWehIbDIhXpgRztViR9xNfmGXsdPfmI46EHY/
21TByrgNzwCMwg1Ovv6GFUNv2zOQFD7qvuPAN4Ay6P75QnyoaCo3jFOmN3TnnwpJ
yCqwuCnwyxAqC6PxqINsNOihvSmhj2GuYV99SDMLNZ04fFdzCgYSJs94e4l3Q+9O
Gh1CcBk+wavkpIrshaxKTlF+26V+omyMlAcrhVAv/IJriEsOUtEjfuSstnpNMThA
2spcgmhA4JeiXTWeyXlQmV8kWcDv1T+82XzBHEWn2dBlpY1CBfbUVnOm6j9KfkBw
OOxXWr99+jwg+BxJIy7lwJ6rKhkPzz6Ywk3jfhTghmvMBFZx5sHz7PBAD2arbdqZ
iryyrnQ6eoGgqKX8TFHLxJWBTnCTXQgbOwHz1fWmiL+5GE8WX/9xz7Y8yi290ClH
15xGevvdw5YUFJ1gDRlKhWOEAkcXNkRYISnlKpl+Ug6cbHpwFroV1DP920BNFExD
Gmvk4y4GKrnc5BpQkYRn/KX4jPM6fhaBQUCf4VWklTJBuc4P6XDob9vcqa000FZm
p51pwU58BIQMdYB9hQYpgntAPfeznuuRGU5j4fOut5t6Da+UTIU8XoqeHc7viRVw
fxjKdiMvu2ZbGURf+6I1KiD9Uj4BfTZyDjaQvu7ePaE8+oyK1XVDUi+r7MAlCEV7
Qic/qoLudJ9uj+vlOwn5bNT2xLJ/QZI1utJpHI5sjaT4k02lF8b4fTKydRX0zuWS
WAi39PJLy6HXm9H0gGgHkqsBjBe4TFyfiCqtdaKsbor4kjkfJD3ahIFx11JbMGkf
AONVJIEjHvmHDBZy5R39ARUqYKkplLPpudOsURZOpu83hlcXgAvy5smylG/kbCZb
kx1jdZaRRCFkNgcDCs+LZ9TX3TjGxEk0Qaq276p3kRRUBhavD5aCd0H+w+dtSjGt
V8vrZli8kGjifoy4a8oRGkn23+MeS1XRcS/g4INSVG+IQnHAR0AGw7k1P1aqUnV7
h0IYK+OTljH6hkCO9UWN0cTHx37MnwbSnyWRGr1PJ8+rliv5sFfJzivYLizbCOp/
T+VRHe8r/LJoJWYY5a/tChMjRtBlNk6GRi+NO+nNdm1Rg/RonVeXXPvZy8BwG1v1
WDJInzAj4gx9yjV1gxNfBGlnV92ePMCG0EpUDHkL0PNDYR4SPcTihwzuW4/sAIIT
1uwDORvI7AfNySpHQlIJNL6G8m8j2mwd/6B2rJXSbjm1lNVoBYqU0/LNjZVRFM+i
/JT1SlZ1Hw6AFfEJ/Z0KrfDghlEIOmMGM4qe2aqkxoxAPkILuJ/pqwaMhg5Jc6a1
ud2CiBLUHxA3rZNT1bAqzEB23Se5l9eQ/slGhJIn+TjHERm9IzJcTAY8WoIHCC/d
6jg4TAr+4vr6WJsxxJUd3GhdG6B2TfSZ21i+ZpFRwQ9/tTb8d+1Yvr6aVEwYmlbb
91OcccYfqdhOiDnxhldn6FJ+6GGNvijhFHTB+5TOTwVm+guBtjiv6xOAgs4qaUWO
xhRDr528/yoe/11HnVHKCIZ7fqGS3/YZmCkdlYTZrfRAoR1zKOskxPV3h+v3+IWq
xrQNmue86HdtvEj8/0IwY03d1mrdoACppsRoTuOG2YkzDjlK0tTswRdgEHfziLaa
y/bY9KqQ5JP/n5Ykkr0ipeZVhZu7Hx18ocMwrCJ7PORcijzdOipdVep8zu0v4QfX
icawW7wl5Y684tJH8uwrgZvt4A1CEVqwKQ6Q6z80tuW85K1INxojQvi5b7Y4s2i/
7FSFXVPpiOVxhxjdALe2lzEbiniyknkdBYUs69XD0kstJaoseMRE9XrbAb0nz2tq
STVphm7cj3a5YWBNTdmrlAanvjkKPpZHxioRzP4JYuhrcAwLCCZ6+gr4AwRW4AMO
VxwDL9kWybDfYQRawAnkutAkxf1kd6MzahAjMRrQsmK3osZdUzO6f2Di1VqV81+U
OVyebdZi1/wEQ7+4pL/qoFQTWGLValjtpnM/sVfBTW3PHOghFfnMa9g1zcvkhdpT
q+WDlwG2UHBsL+OE7vFXGzuPkoTJbPKlJKGBBglCN70opAXn/yz95MF5dBBNNbHm
4q8yCEInsyrlumuztICBlCGV5stwOzbJOCUU58s9InGZ+bvKopYWJAATfW8SCZJy
A+IEfw0shGra1+ZPyItz4amcPWeI8FtDPlmRKe3yb2PHaQYNO8QSESRbe26ylmYJ
IGwIuPacgKOBRd8j33qBLMNE0pV8vcBUUxCI6cF/NJyaq3H+U3DK9QP49Jvvg1kw
tKx7KbGLbWbf+ndTLC1MEhT6jpaBHdtXIvFycctaKJwe660gj12Y/ABwIYw1KZw8
5m+5ED80LorPULK/NMncePXBBs4cwD/bkAeI6plysFlDkntl/efTsZNChnmHmH70
9iJ0P+bK5fjO0i0uLbYnbWxvy1CkWhJI+eD3x3E/hlII3MN8cDWgXkVktT4GsBFR
xXFFI2SdmtT2drHxv8oedFbRFvA5qo9AbSJvq2Xvssqbi3OwWiGTOSBCz1U5/ddz
0oZjuGPUelmapWs7qU3xCTXD1kAuAwww+8s/lACPdaeMquiApHjlA//A9AmXZsPg
QgN+NEC4hJzqqEjmDs/9PjUN7yhjh/v/JUNYA/2LSIhhs/lyMqoORFNfk8+c4DoW
oDrX5G09EIGPYNWF52p9aF5r0IqROSF1+hKH4/khLfIhfLthzCeyK0L/XKE2rrrd
t6tXEMd2UISjmV2BXfJF8yxf/PuseXgHNn8Z9D6Ag1HxSaHWt8CK8eY/UplUp8cZ
Ulncu0s7tZ+B9PWu8TOdvWhneRGuccc0hUiuGdxLH/255OzJ+GZ+T4kjLotn+DNZ
13yBiKX7j/AhGWUq03PldDKUxwAZBl2bAsmq6TvuCIHkb+TPAxcZ09vtndfMbHrS
1BUiT4KLlf8X6rsuUZdnup8rODuemGSfd+YEAEvr49ZiqPEY2IfQfjQgbJSz4i5C
NDzO02jjwm1hiSy4pig1zFGRSoJiC1eM3pd7bl8ilY+YocAplWwVoFGmd4wfI3en
c3zQWgUqT+Nq5d8ruqgRQ32QOFZQKC+vgHz01+mMVEX1Bl8MCJo+tFl1ZumHjtEG
NfTMQOiQkYYVjTdpH1qvPFTjs4qH/Pahpdf8yl3Dpad96Kn4tr5olmpBGxr438ja
xU+NbBvNqj3tIa7cqi1d8SGXwooREPMlQy1iVDPdpz7/NuKpkH7/Sk+n9k5ipOFL
Zh8t7k7Uc0Mxlv29X6tGiP+181p4ryHyXd71Whlj+RvhhVd62xVp/JBYHgoqfNJl
4VuioZ6asqDr/JYGqtwOxenwMm9qNStDfgH7owD10lBraPkLzze/Nxx5ZvuG1nc5
xxvEORcOROrbp4tk9LtxIozAxRB3lE2yfYggv61OKekyQ04PVPalNTkRj6GB/4zC
QoJI+O85aQXwUvgScnGyWSQiHaT1mXQLxz4+9pIRuFhFQqPr/iniufr1drTfUrGx
e/5a+VZiSTHWebNvRCit76fYHX6kdKPKy/ncjNmUbhslwA33tMe44jhR937nfe8v
eoNsSxgJkUMghzahkSCerrVEyGHeqy10Uqb/LH1itzgnu5ZnN9ketUKJ9tNz4Wts
qkGnVf4vypWY41vnsq/1f3XqFOvx5Ua2PWGB7hteCpbfQXtUw2PCDT+kH1RuxC5f
HvSWzaNtfeTkhqOuS0LwlwoZu7ssAjuEac6bbTKp9EwMQCsSUYpFeGuEOo5cBMHg
dV1wAcSMVJU2OiOMNgxxLxrSeM1LL9NVcVLvhoWr/QA0ixPeehb813Qh8T4xBv2X
0k/E4nWxZSzENr+7RRZEktdhmOQ6iPgDfPEwQuPHbC2pOyz3Qd8Nc+ppaHX+/maN
UdZXwn7nypWuqIdr37nzub1y01FKJ4GwG7nUG31O8ManEmWWom3Kv5FqgbygyJT0
qLW8gdrMIQ/xH0/YhjTaB6eiJrF2P9gkh5pRUCHU30EGUC5wGet3h3zevdvgJvIn
C5CpsD6qiT/PJpmRZoTKVUmS2+D/ROuCbCFPofE3BjkYLlXPGYDm/6/9c+1nUkb4
rseZzx3Glv4v8PrciLaOYtKpCpyVY8YNw0lPC1F1AXDTwVd1K9mHdEbWoX5hHxAu
eqxnH3cWIvsucMqDI6Lxx5M/BIiZChPqkcZhZlQL2MO8nP5mf5kXLF/DcyNrzovO
KFLMMNZaz+mjwEdID0ZTOqLKLPpIUF5Pshyqz7aLXE+XgHlj4zoGU4gt3f01Kj7Y
Ae30B2XthS0I67q00UQM8pN5mjduYw3bx8N583L3MxC79DSEcla760buLQo8gevC
Hav/Bc7XDgeBrNyVtoXGsygSwy6xcOSyGxBp8uuY0CMT2rqXzLxBCJr0hvw4s1WM
LG9/sdTR6zM3bMcC4Q00CLi0b9RTNIM0xeGfOWxi2oQNmr8hFlCFxrhJjW7JI3KZ
BKVd6nqrs873Gc8BNPEq1Ak43fdai1R6X2dFyd++u6oYDyCJstUrnLX6SkhUHtau
Rphoc3Fom+/w8Nuc6nb413gDWEpUmEEEvH+n2wCP+Yj/GNkneZ91Urwp/8FYol90
J+w99nGJDY9IOtc/mbKcjknICJ1zR9QILkGI3hBZUJBLFlmC9ZRHOBcONNsAU4xp
8e/3LKNu40utPal8kM2IRMPyPdV1v1DT1Xi5BZ5UfrxGPKZyCCxPUzMNKuMRc0cU
TDXm8cbxmQS357TK4ePApxSVbpBzsoTGxxyj3YHj3CObvcmOEN9lgHKYs8JXfs8/
IrAFN3+hk8K0nUB8zQKFx5iEpnqpKU0KBZJcL6P9Qvk=
`protect END_PROTECTED
