`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNlGVxaOExg5b+JHe/bZS5WDJoFbKdcdHJnO8ZW8koICH93mRXOSkOSFuvZwat84
j2/JHc2L5qmXjmD4sNHZXbuSdTjMg10RZdKpyqxfyKhBsKeMMjD9eWH1ZS+SkhLu
XHFpuK8IQ2cb08xl5rYswgH6ZsHwldIHxjmGhdAZVlVV1OdHRZuKzKb/PDH7czzD
EEbMHV3uWyEjtT7eHo+7LM7HT+zvYrCa2pBNxn2SSFcu/E1NG8IwxGcHj5tAiE/6
qvOm9xEckaUdNcweJ4fU/pb41nJQ/GjKGCLiC+4w3uLEOH56jtip6wycNQu9Ckw/
n+tepTvE86obqXI6ET+fDhToECBlCCaj5jF7hxMc71ChwRXGxxOjwSGaLZ8i3bzY
BEuyRhkNn1G/tabxEe4vylG4fn7BWrFBUJEjELjDT7e38wQuIYOsq54r4sVu95nk
zcUi2LxPQgAccL6iqZtBfoRNP2VJ/FvL9a+U1yaoHlA/vygSdx2BWgtzUoMpTy7W
nU/iReq3qpgIecMZ2eKUEPDLtPxDoYHrkBCZHBkQ1pclQRCDbcqf8v8mbtiXCKsj
ipPQddZ4TIgkGF82NYRftbTCOMjBLSYIeC09LSuu2uwVEREtSFiii9FF6D5IxbDP
wfWGVI/3xMySJdROFL4bOqenHGD903E8J1iofLbA5ZbgSmbssN/JRoX+ffq2G7mQ
0WzX1nczLzFCnCe0prtWh7IthHWpwuayXLYNp0hQl1/aSJSl9q23p2dofzUUYAbg
KxDjjxnYD/VMFO3RjScpPQKqkBpJC91VAEJZ+WD5fwxiU/8uRBNJcfDcXRueHK7s
H9dQ81G0a/zzyFoj63muTQ/fw1QUv47YDkrEksWmvaUgEhWuhmpLvOxDg0oFTvyQ
K23kUIxwnqrgRg7uvvGnT9eiaydhauigncAZoRZsTNadKYZhMRib9Uq7aYZA8nr3
GZDnZvmG5ZknFgBbxl+5ww==
`protect END_PROTECTED
