`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFOu9joU4Y+mmKrtybvfWba8KKRHVdJrjtmB/F1kGvWUJ4FA+1RBEo0UqVtRinsg
qXQBw7SRKB2rVyZThgR2kTfCe/e02Wsf85QTv1TxsCfuoAazMeQ6L56HWKYaiHOS
26Vw5Y6syehvjKJEXSCxbOCv8UQB4231WNcQyzIIkx6fmJGnc8gQmylXVX3Klxqv
L1YysH7dDbnE4w38y2T2SXWB29q34DgePOXREEn/HtfeZObfXY7umDlyMsDn1svr
ai/2kKLM/ARGb26jAFaPyb8RI1YyO9JRku+FYpYwjYbqg1f2oitZab7od3V7Lrq+
sN6iewxFi3ECXU2ojYRMqUW3x8CkY333MjUMU9ZLfxPXp1IC8KSyYOCWNTQ/9l2N
D/omgTORL//jAvD2QZYl5Ah19pYH4lZJgZFJg6TX/ACo+8/rZcZvIFf+U7mtEFcf
KVBfbEb4aB1FhXzQyoCq7orRz5JSCPyiKhB55aKZzuksVyMZ6JlnYeX7mr849PLR
ZOjj7LwqBQCWgRN4fJlp/+7Okv9nDipSGaSqOoQqwsJkC8XVMneImsaErcsr+QRj
GmXRz9Gmqms/MHygNA+XFygAzWZauzL6lCyIZXLFVLl5SE1ub5bz4SFpAHnQzxJC
Dz77uRLTDZpxK7l3CmRXEabiO+3xEXdKAreO3PbpBBE=
`protect END_PROTECTED
