`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FOMtO5S+bck2mQS0RZfG8GsSpLyIjutKqB8KRszt0mgpRxnuU9d4WEf7Cf2Sz01
GrVfLnUp5OwSLfH7usz5C+sDKeof7jp1jUjZupK6frjny+F0HnbqdSYMvJCPwsRe
rYOYzF5C77ojFiw4TCIgFj8nD4zIrW2cwt/Fao7uaD5e9BLWPhRWAtKZbxiAzKNl
aA/Roj0LarphDeOLVMhg+DKnW0odxwqPS47QJtQkCBrv8puITEEnDpkKqIv/LknF
oeVYmraH6VYma63V7VzCqzwyTxQvxNImmNx8L00n3Z0dNlKjJTxHAlbNohaY+xwU
Nq/2qIJneRyEtowWCuVtZuT0AzZGAmlTk5yJ1uSRs2KY4kmo5Of9jJ1iH2eCoU3L
MX0wXTuAticb+tfcBeto1waxE/vEUcsDyoJG/nf7h4WU8rKFACHCXLFGpv43XnS9
FxwhI9CBbko+xrCBNhQgdw+NBCKivT1tQbuqsYTID+JI7aff/iAozR307/PWn+Kx
j9j/uAcWMFHrzN0kO9yhoV0M91JdLTUtM0Gz+AvE1GUOxOE7027w8PNpD0OA5aaF
PH1EIUA5nMSwH6tLTSq88IDCx5hXut69Bn3WKFJ5bdYeXeqVVO+6iapxIOlPiJRV
DbrE8LPTKD+beZTZPUbiiTVNCzY5aDgwMGk3r7hHWuQlCGFGFJw68+tCImhK/nfy
i16uzQrLWo6D7DkRSA/eKHB7KMIx8qeNk1+wegAWq79mQWM1BLYNTs0voidd2lq1
VOc2YOAit+NvPcMca049pCRZJioHpTiyFl85zqeaRacsz5O14gSDDnYvZhoZnoId
0ocmOPKtP/fw3ig2OC8+eo/D0K2VV0LNHELmgh5572PyrSKKhCX8OYDlpmBOf1u8
SAU3kz4aTwUKA3e5+ZikLpo1jBRU6bHQoYG6h4XK4uutAutOB30Ymm2UIhUH/klQ
LaPSbtXYMRlhMIkj+NbqgU3wwKOtYt4ruJtsUHgHWuQACcPfa2q297lczuooK85G
KZP1bQuxVs+0w/euWwLK1OSXJwxv2PhJNbsog7Be+e4pUCu4n3TMrujyjkEzdLfu
ILKYd0dSG7HfeMxR5sax2hzIQsQ4tdD4B8v/68xpe4Soo27VHFyDBvzC/oeMW/wP
bXrfRb7JlQbE0RvQ2og2SKLdHiE3vcDpbVPsMWdgfX/8av3f3wlxRCajZ1Wj0twD
sjqdwcrb6TlKe3Uk9XDk1EgVUl7BJQUBI/uC22WfMFTP6MjU421T/FajJl8kwlQ3
e4NTasbxeWxPRevdQgbR6fJgN0Xt4y67+3fHaIet08Kt445jLPVnlvFueEWYmAWg
ItDkKYHzCIk4rli6AWJDvlpxVI4DIQUrr8ipg5gy+L0/jB6zqj9MZKgqGX/6zWPH
GRVIKyhP+w7/HVfWk1pkMrt0APnBfpGKSLRkHXYTC+5gGGBgL7IKTY7UAMpOdTxr
feF7/Y2qngXZbryf91wmRt3axZBVs5atV0m+W4af7pKIRDOKvqzJfthYaOCdTeQ5
lm5LBymxNjG3DZgac7+la86c6J/qNfE3398axuqzB6xloO/YsOu1Krszz/bLqMPp
hvbZZMKcy7udEvQU4V/VRmtAHcfEh2TlqvCnXkg1Go8SRp3QIkDhP1JB1YfrxZxe
wSoIg2mIi6553C3xtmyH6J6RkrDXCB7dL9K4/wKwstvcpB5EA4DNnpXi+rHBvTCz
wvWUreCW5v/6+AUHfsvuL/kXnVF09yn+Fx1wpWuLZPL6mlL0LSh0bBl0wytunK6w
TOm3ko7CTK80eB/iT5PpnEwE7JNusgHoN6etyKB+66OwXXzQxDIojnAFz/mRzysS
Po2R5BGgQjwSmlGixytNfMAUPjL101HS8bmcGaeAElWD5QYG9MJG1DSXW4i3Gjzy
nuNYlo72/j795y75ToBzm7Vg6Kze7oEmBrGSvYd9g81CtdOPkx4Z5wULOq1sb9ns
EsidkbRCq+pBRc7IE3gJSWrTIFoE9cFp4as87O3NOgFMH4K3h/IGY7zUi+OfFqEy
x07ldB/9i+RMmhUCqbgB8qJVSguz9fKrrnKBMsLwB8bUFe1LGTflpEAfPwzDeLiR
qxEYgrKcDGwOjLFeSCvy0Nfqjd0qPqlKZcqugEUJZqc8FxydnCb7GAMGmqH+vlgh
T2emBfyiM0tuMQ2wmvcD4/dPP7hj27t1pTAk9hg26TWFQuIYX22PomoR4DX4CAvj
ZZjlqqxBQ3Dvqpv6mWFYzdnyn5c+2LLR6gOCWfqVI5zJlYJNp8vb1GWfDhcRvhhq
MDqGIMH2I/CQv8jermBx1mKkOkjerDWmZ0tsP2FT3/njgAahWrBGgXFYEvjl6Q0z
uTekBpQlwOSi62yg1VseQcABgkCMHGaa7B1QUKXuNUABLjkKDUj8xkpFepBlH9fT
/HiOM8Z5XQ3ltKZc1mf2vOFKK5BUoo+AtUDJRGDHhoPD1DkztBKrxEhmzwILo6gz
WkgMuPhyKmVslwQazFMhQbaiH2htHE7tzkXj66D7SWJm+cAAzmYwtiJCg4NyQ67u
qVfkwsMJWZg8SVpCFmaaslEYm2weaLRnM6+KtjOt5Rt0WoENNSecNk2VU131Ojgo
64h2i7jZ1VgHEryqHLzDSkswY+dyKQhQHczQwb1nMGjC+rhcV9nGaE7/r31EVxcr
7AGLJBbBEXxAdtk1RtFIX0pa/AggGDNDrFJhUs4EfBxeT+kmqIEVsNVMbR//6Skj
UoQJMCiGx8gmZsuADkd+r49rOvY4Ujzi6iQvyyP2+g447ENUlXRVhXuFKVsrOWd4
eICiBiFMI4v6UhoP1uyh6w/YZDAaaW7yOPijC6A5Z3LnmZV+Ww0VgCMe8wENbJwa
drykEhHWAkCrW5UxH+O76X9hAZmgY0K3pv0mGOMo4PAaJIIdYQm5zAghg5edgetU
kz/U6vhzWatZC2m6KrWqSENVPAbbLWlYU1AOnLN/vH66BaYBNOV7SrVatF5b5EAU
tKDHol98HI+cBkXt/jEoVTwQQn4BZyqLwp0b94xFBLJDw8h+8Faod1onQeGkMD88
cj2eEZLWDqhWVOTvv+e4673bZmFu9TgH2NJOuh6zTiS2Ou7fezb6NHSe1bmuFZs/
koJFyFa99gKbdePCUOVPvoNexVewUaGTMtfJo695t/TmOvyQ5v+dcMKuAzm9ADOD
2AouHSk55oC/cjkMqVmGLqIsGwIqHtmjjLc/Y3A+LF+ZAmWNe6saArVpzIu2bRwX
H+tbtdN3euu4rlJYzixIo5W4tGvflsXhY6D4DE4HO7n6nyXo9v0KV1AkdFnTpE57
pPHnz1jtHupQcTA2bcIpf4DLveayamhb0diG4LXwIGYtI7emhW0E6eCzsrkvED+i
rXbM8j+ySM3J/qomYvRGh61axgOdASjx5pZ43IY0LDBl6o/5eR7mKFu/tzVk0npz
LDfG4KelJPFDJo3cNRUINH8ie35qxa0DqZrrRB0tj7pKZhrK6abI7S4uyRqS2A4J
ggJ2Mn19MhXQQBa8RW73o86CULsAGytDOuW8kNBiMoIv19Oz1y+8EV1kxFvn4kvn
LK0uOz7kmC33ChZXT3NhmOHPcjZFpx8ydbMzHb+Uh96VNmMjZaG5TCg7PUj58ABx
gG+hRevZ/kfx9bDiE6t7M97jAX74/2OKTWfDhGk1UtKeAKPzEvf2yBN2oimkI8He
vYIej2r3xtEX/ymdFK0+km8rYETjAEAGs5ne2EIu0xZTqKq3lDoJHZUiq9lQ/coy
fpGgOhHrXnc+CAjww6dxPTuqff65BQ3UsRZrNa3mIkwX4gsRqSDjbUb1IAPOMuPL
2wS3P461Hs+8BjDEkyLWLLWW+6Irz+VgcS940QBdScz4/PIWV7KOt5cmpn+QCIbd
YSweNRBbMsgXWhm/PbWqEMaU0zseqeAJXhruh6AJs7KnVvxTqO5TWySC38X2Vwqx
8YEeddhyCIVb4cmMG6tZWJOiZoAK7nga3iLZTUjf/LAdaOplY58Ey7BXkO3BjdvG
XyHdiiBxEUM8lkCuuP9e0NOY70kOweERoms6xnegu4BaD7yajUFqZ6vYxFeyKJxO
NXObDC8kpqZHlf9Zm2nynwb6nYkUTg/9jgiyP0TmeRlvYMl84o6v/lA0OMyxT+c5
KStUJIJv1FK46OUDGxj1aGxCZmzWdyuJnp5uwAww8YP/eCVQb3a1fxq8ml2VBi96
DWtXNXVDe2BktmTnb56yA1dI3RSqzBiE6Zk6s/4Z6Y6WPVu4WuNihitM1argWQyc
NQP8Oli88D/YX+QUif+rJh1tbvlxPPwSPa6cJdGxw2i7ks0gYRNlTr5E5m8B/lrg
4JwZt57rqfJglOfcFOuK/g+zmIn9xy2ZYMvv/WwFmyEG7tHOXMHBnSTSEnJaPvro
HEvYnG8nSum3Ond9Fty1E7M9bAXU0RGleKI7T6dgnQ5XyqNmoAsWecGUab9NYZr1
`protect END_PROTECTED
