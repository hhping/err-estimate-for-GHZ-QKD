`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXrE8qJMpzsC6JHHxAGdyQWwzwAvm2NopTtedk8paxQt9k6KT0ycFICCrPYjIOpb
RXcZZmLielA7PNXkj1cXHPTU6AE360GBkizeNP/6U/u4+x3EyxwNuDxuZ/D9aM5W
UR2Nd7HXwUn5kM/XkmqariL0jc8A9kRJJABFWQweGGOo55LbyNcJ0LLadN54ZRqI
qjQumPAZab8TNTmDQDSTRGq2+UySGA6s8HzR85iWOoHVtB/ZrekhsWklzNGYYgd5
xpCPyI8LgDLaPn6yJRWPFcWKdoWcgVvfx5vid0ifYleqfAnkEP7/01zuEin+NA3m
EMckc/SQa1J5fTwY0aaYXa9hBjHBfKfi9uUZNMz3RDXUWH9kn09mSThsjUQg04hI
0+sEJFtDBJ8uXjlvVkCSno3yO3Pwu2Ljzktt1XnYLPMgnDaqKQ6kmHDgWx5aDx92
GDo4dPJ2EQvnOsdUze6ZRQJLyZP/ood+MxrFghgeQNv0zwwL65gthTjGyOaJi+Ze
/gJIJPYhBr8GcEtUMxDV5lpdW5i8OSF2rmlO0gr35wXAAr1gk0Y2mvz2DnlNkyCr
+LfVTwwfmrYVdpRs0Ym5Omx8pW3brlP7nOr4hG1XHRv0Xwvs3rEl2bHNCcX2bavO
dlccEwpnSDijc5VRy552YC7fpSEmobSMSRZ9XybmFmdaJqNiKB2Bi9vV12pSeKDw
5gNsRnR0Tu0yKkFw6Wh2DxPSKJ+7Gg0+hJgXzTBiPxjc8vgyNfYexko4Run7sHif
`protect END_PROTECTED
