`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7U8uGqjMde8M00RBt11Fsm4BItdrB9YglQzoVztYe5acbsntLEMw4l5KjUTD4ZPx
8+hFM7mVCLuk3zy/hrqyyPelkrD99AXh4/CWRLwinpKczzFrI3YHpygw51cPdg1y
k0vSS73/euB9qEdxmf4gD5n+kIrgfO5SXKccQTPY2fHwg2651KjJuD1p4augU4A8
extLdSDN7HxH5+qeuz3deVdarHf8xgQZLlC4y4M82x8aeMhwrHcwe5DV9WfhG6vQ
Uz3O557M31b/khVSTjJFoaEWRWboitwkEVXfCN5XYjkoNpYHnvXMRYH6BXJhVWwb
6jLlUb2AymQe/Gm1r3/x7lmVp7INYKU6WXDv6SX1rguj+HMpa53pN68gcoymdUae
y1x/fzZ4qOnr+EqpzHLpu/HAA/pcTAnkL9abBbTu9PCElv5eVioxFSpomAM08P8N
jjyEFQcZAO7SoUVe/dyzYcH9PWFmSOty081lSDzcZcp0LhLmm2zOmT1CA0te4pfx
Pv3Uo3Vwy6ywY1ci7LnNB4lv+bevT/CDlEAccgwTfXH/R4OLSxclfV/U8Z1tNgGT
Hp40N9F/EYM5ylr06xTUvyaVgFdQlC2byEA0bY9SSfaFkd+surmOo7ofUca0X/7/
yK74LY4qxtqWs7FkFjhRDfCI/NQ7Nbn7K/4lBW5Ug5VbTOAD5YV7YgdJCyPe2a/C
QfoisTmc6FTk2HEbew5zakXkK72Nuy/voxc/lQfivqOg1d3cIo2WuqkAJRKLQyky
ItU1vkXoowE5yV9P6rFMT1Rc6vuIYns/PJ4V7RdITwBJHQPrdbXzSlEkaGgoh1h1
QGk3V90S9ReaEozOMRp8V2Cwwvcq2jwtWlkntRyL3U7fmgv76FR7p7sLBrSHSfGE
yCfrOG+qIpNvMjfuAtbjlLvjdotwwSlnoe8IZS+v86PK3EDfmR5OeOa/2WSiUg0G
FDw6pS/ATXn1kjr9m4BiDncM5KNWv9yijAIOPDbOaCRzFyepkWhdyv9uUjZlDEFI
VHUvfZIZeee7Oa6soQksZlxX5CeZpi/p8yFOC9POsFjEu7M9p5DfS2imzILrpAR5
ZSvZ9yC3mPYrSUkM8pYvO2mWkOwyGHUtrkuYUKu4JlWvq9XQlUny7l2gpFeOLey5
qRipkH0tPlLaHt62eg/i1PLNicVqdplThVUXADqz1ZDmWWlPYS2q4xmtokihFAYw
lwD14n5arptbcoODse3VhOIUDR16ZeZdBgYIupUaFTdLfj4xekS1sz10FW2qixY8
iiCYNVLAMSLe9Nks9ricn455Zg7JErr+kDkijkcsnoTyYrwtV9itZ8h1tZcO5qxN
1GKup5M7OA+qIVdLEuxG6oTyCQO7bx8JIDcdzLHCFePIWXtBLeSljfgw78Hx1yau
PbuBmxutlp7zsy3WCmJAHw==
`protect END_PROTECTED
