`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UV18s9p2rUaTcNBa4G823FKa8ywVkVSZD+KspDoem0TOpEeXfoNGIjsTric45OJ2
pbSfq8q4FihNb9ZwKO2SfLG74l6c7NG/M4VycV0FiLourbkAgq8Buli73fupvKL4
5TovaeZtfCqZ3jAA8tSnx5fkH0UTSS3M+P3YDocI3nai2YVDzDuT9qytTLKN6myl
NPyvvKsF8dRcLanzjX7VqlGQF3Dm7wrMtDtgUDoiZghVmyZSk9PjEzg8deuCbgot
qHGNbk4H2snSUBIH7bpmHTPZX7nCL4JnqHLLjf/8KS/i0PFgSyo8+CjrPJ9of78s
IH2ZCIpa/jxG/EAgdKhv+T8RYpVZf9upftxg039PILXcYjX5FDw6wKUsS6xoFNC8
Oh3pdZxPeEaJFS5rDC1C6JBLFvJwFmcw9pOiFQL0wnTobD7Y6Nu+4ZpiDSlnMKC/
0Yoff12TBeGrKWQjAWV/86t0b96vTUKI/sMek9e+/zpusV6NN8HgyTw/qU9S8ypZ
dMQlzTZ0T3XHoCOSoUzH+jy73bt1JvTEhlSrWkD90vkrqUYqwEesMX1GSKkhLOZS
UOji7z7hMkQD6oGdBkLyCSsCCe5JwSbPzIRNXV3g+0z3y5lq9hY9fObO9FOtktYM
q2sxUp5ujNgtzibnekifU/If8y3NsJnyUI0AF1+8TBuSJOB29qG5+er5AEF4XQNP
/YxJUCp+d0ELLrVeAQV7bSqy1laXu5pXRONO8nEbs2I=
`protect END_PROTECTED
