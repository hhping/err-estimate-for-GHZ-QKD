`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWWZyUTj+u0j26aF2l/UDdRG0xlr967/lMcwcr7mx/+MPathP/jhqG2x9pzapY0g
+nZjbNROyJrMEydaB9CmdQ8q/TzwrtJRb4xfOQFUpYue4TzPylXcSDuMYFJ31pk+
jFMYLrGc+XN/M89xWcpa6b5WTedcZY3DLv26eRtLGAA4Tl0YsVOMnl6tes9tCyWF
uvn4vb+mB3B5xR1ix3LrHweREC61G2wZ6Y2Gl6mNmHT1l3WWG5yeRYU++fe5U4om
CPZ8UBqrCZ4TLJ3qtTBvQn3Z0MytcztQeFIj08Vk0PWvp/7kxg9awmUy8bY1cs8u
6Psn3RjS3QtKn9fxxNmgeK8ofgq+IM6pcEtTw2geoP35ONP9Kt3T8hjkUQmfLkEo
nA9PjSNLYxa0JL69dCAIGlaka7PBOrF1OeFRJPnOQzkzJhAs9y6jt04HLg10C4aF
A5IHvxyf85inYA02BpbyXvUemDflS3+n6zMSpKgNQJoUQcfwna1dNyEosPrEeJTx
dCkfTFiv0qjuF8XFbX/gkU/bift2G36EsjEnADobvknoVu6TG4SOTr3qjNwElNeq
lgvB+1sVjZ+9GRAKYRmJXo0RYDJS+w2jhoYaWdIzZAnscS84shGg/H84/h2bn9Wu
fYiNXcaMeg1N4AACTIo/zYhr3M3HrdHLLYN0wLUR8ciUr+RdImcL63qzD7/100ge
UiOzzh/9TOmLkLa4ejxBhbdwlRXYkmAFQdIAFD86Uvsz9aClp81pxqEJ/2TTUvrw
3rhz8s7iMVtqgRUJLK2Rlg6pgLAC96yAipQaHGQVLfKE3CzLbN50MkwnLWg4Wd3B
LTWU8DQ3pB1ifjp/0EDWvXJSneLkQuvUU/XJ/WjWurbCdOxHu8uNaZaSH5ZPmCVr
WhwVndd6pojY26Z9orm1FcAj9evUSj+KwM50JLa4msnFN0de+HBb2G7atAgzWO+1
ZgqvbpKS6zaU5UySa0fPWrw/rZcHfn7OC4MvJEJuQ0Wst8lRmNIzlX1ru2cmd8aH
tK6SdryHlqjm70dZb+N7nECWO3Qm7APfo53cxxCdtqiwi3+SzeuuNrPpnftJKaqk
NlUySSwdkCl0N5PMCBzaQ5BLnt0oHDsThOQlP57n6RdWjkC2Jf9u/Cw9mC24Sxb/
E5N/jMpfNflmAKniNYleKV06RjGkWZx372NHyU7gBW4g5pxKMpHIhK/A7dPydh1x
OJVZ2oiCymhwxgm9+Pwr/znI5L6IAuVzAo4HrL/eWmqpd03JAvl+Wr4qBe1Rhlcw
zWJ3YM2zdSAvKxDWMmxKCdb5DDC3mxjvrqfi7JMeWVqANKotxjIsbe0RXrsqiE7w
ASWVdb8jIsBvViTo3dYjglneT8lGfbxWiojoHnKy6wm4Tp73KeXRkCZoUnQlUExQ
1iEHxc4bU1/GfpQiCu4Vda1aF5S62K/ad4p1Ci3ceMfrlcHozlxDb0KakcSgy1d+
Mt85vBhOsmP0awVVJnp1jQ00EZGlarEO2bNcabAmUEsjIxmOwlkEY6WQrtrvuTla
xs+sbpp9bp8HcTCSznw1F97AoiMkMvejV1+7EebC4/7f9szJ7aArx9xPx0T3yMgO
jYw61gdSEwGQNbijVqA+gjU7tF0G3oIDKekbqQo8Q8SDCiMwlAYTR7dGiMv8I2pn
RWZJ+oeMA2YY9S0bocyv6WJrSJ1XTq3pzi15QF5EBbgyCGVRIDFliWC7avO+AKX7
pz2NX8XnOZ/aoCCCWNrN/mxSVfyR9MEy5AxMpF7Eb9Z0NW2fmdrgLDnP0ikg9b4g
7EDUS/neaYOQ002+Vwzq8T40NuWcAwxXvPhpSKgJChEK2EevGbkEOQ+n0Om/KW/A
D2a6j8cQtjKsjfu4vY/kWzWjuRou4uAPBl8Di5QlyGEzmbmEiYw+0II3XcCxMavc
auSioJLnpcgKGHPZA8erJoIc3BdEJi2Y3S1TCUTrTOO5+/I4K2Ar/Idu03aXoF/r
AUtkKfgwnZz0r3JBwfuBaC+8uL9K/TRSIrkYvAroOnGYXu3tROrKuN/D4GCcU3/I
C1uYARh6AR7hzcLGOLeldEhVIB4eXgPo6Jt92H3jr5LiMIRaxi9wMVXCWQEkrMn1
8cCq3fdkoEAAk6aj38S9nI6JG5brA8bQnmZziFM47MwPcKQ9yVYHHJ/UKq+6ZtOh
wzDm81r5iNnrYhxXT9LoNBQhGyY9Axx8N+fsQTZ9nUHDy+PddwX+m/a3RiOn5f/V
zds/WF0t+gyCFG1OfEkaOBDZeE4NUq6rsqhCBSj+jDFmC+W5OA4CTHVs6FObocKo
pW0DVKUoyqqezvQR1gUdVjtIVnGj0DVZMR/2BbH0caKLpHbbLxF8Ga6HB2D1JsBi
iz5UlPz9Av0Yl5mDax7rME70zqnPhqMTXKZLq+LmQLPngTw8y3sEpuirRM4EoEq2
5vQJvWijJfg9EyLQGM+d7c9bIF3bmhFvHHfJOC1TK59JL1QwRCA3FxPtej8n8sHC
bhGTrA6OBvipPqFQM7ry7nJOoZxX1cX8I2OIm/0aIqH7aQRjpZA5ScsrsGF5e8Vd
kFRpWw0qwh/v0G9jKdVYWuz9D9SNr3TVm1ZLlnO28MULauH/XIO1/qr4UnJP/rVZ
2dxs85hQwnREB9QaV8Ko0YEC1siSdw6nuE2anVA0g37l73jH6zdNQNByyR2ZdaZL
5Vd3y83t3eXRzRdWTkKnChz9EPAFlDyP9qZ0H/+jjK4P+iHQdnUYH/4KshY6Bj2u
5U6AU8dvKYcDKrGIZADdlM0BYEu90/TeiP5hnjawyz7C4rM4MbLjVV5H+puBM8ko
TMQHV+fm92GbEVY5PhZUp5VkR/NfYYKGWWC2BPCIPAyvtd+5e8NrZqPY7lfSPTFS
BonC+ZHluEPe2dKWnwwlNpqqM49WAUy7TFnTlMC/mF6fuINnUqgmGWl1Sh64jwFL
cAeGPqpfXJ/H/fu256PFM5M6vVwYhX62989gvPQm/2SJIyCqTfQZn0s1Nm3mtPeY
gE99hLTTy6zcx3sLQmQ0DeEVTn0tRsHoFMKAGqOTZIoIugd3Qb0gwXZcVTiB4rTB
Fby4NmEnaPdrfKDpgegwiHCMSrZepmgNuwPK/dT+/4M+jjxBUdyJuaaCeTs66LFV
ViKRpGemyOma+6R1lNbKhcX7J6U6/qKCk2am0kpO80qa0Gqk1/OhFsKhRDFe8oJt
XA/erlCiuX3jKsKuMtL4lKtQoQSzsxo9XxSgnnIyq7UQZRml11r6F7ts+b4i0uSc
K/SbYLXPNsO/umtlZ78uBF70DXL2M+XGk7IIkbjU5mEAYy0z0roNsQWueQjl8MZv
zpmk08npObujkF/KbbyJiyqIlEjHH6MAQH0Bt+zfRrIJvPf2/DlI1d19gOVplzHl
HW9cZXQ9kCq5waDssqUvxcCWUpCgncwi8H2py4+VtVBui2mqo67iEOghSsTa86QN
4ZTbV8C+WlnzSTFIiNx69iXYYzwRpGJ9k/rtyr4ndhSHjvlOI+CSJ8E84pQTMyFU
zsBIaW9Kr8RJLOXnjffOPmo1X0a9ElWahsHw+m2h+67eE1/ffolQJKJ8eP/SQuFn
dSWGLKG2vP3yLvn9QdYV7PY/LXH5ppu5SAgGsTXII3ms1pJV8C1u3u6lRvVf1TxW
wYOjCFr9cJOwo/vQljk7VHfi+XjeyCJT3vUogEIlND0jb+/iwvBrrCTCRHii/pOT
LGYpafxv0kgtHPH7D6z24EiL/j9CZ+mcw/W4NYmngiN6JKKVsnYNBv0t2B/HPa12
iTYU5lVsQ6OiSCNIak42/+ZNAybT93L9g4GnzNaLopcAw/deQgfkcrQyIskTP8Uf
nDdq6hVS6hm2NON8VpSn/h7+AUcnQJEjy5KnF7Ci7jVf+KVIkU+vr2pCDnXYfN5C
E0RsLrLTZIcJiwhpv3FuZ9tkN+nU5B8mmG+ffw/NKjScwDx0326/VtEB4DpRrPwZ
eMq/ksBgOeMrYwmPI33+AjVvuBBkXPEtOR3mRjIV5YKxd/Haw7KPrJiHzCT6j9ft
glr+Qjn74PPNPVwzSwAdXn8AI0lJwU/vD24osyqs9aio5XR1N0o88KrPf/VDuHXb
osvWxRRe6nAX8WPbPpmBMPUEws+46FFUQ0zOCyYxucGv7Q3GuVVCi8kQrseN3N1g
3LQSeiLA7BM2h5isfRIfmzNF8KBtLLM7BpNpSG5pULv8sktXiLG899MWCKxDTDkG
2Gr8ZP1LVsaCbMyqaTrbEJ+Pqwcd1X/iKjCv5cuBqlHEG5REGzujlj6dUcfdNvfv
qV89p91BeQFkO/UgUFbD7ZbQQ8E2sQBMGIxJVmzkxW/fQ9DxhJYSICkERkgB/psg
JlmgevSZrH3SzwBYD+hiYm0KBO61xxMJSVVD8dnvYYm/FZlV0bGGzP+vJWB1LFYu
KQ8m/KQpBGsmNWbCIE33B21UEzQzSMIr5o9kqF9NQcsT0YAtn50B8/b06cs9wK1N
9VlVgRmqvrYbWO99ZoFNLz6Wdg7FevoeOxxRKZCfNEXEbmkieTOcGadjHfmjI4wI
jlt9S/SeI/qkzOTC1NHqE80XG8keDeQAjAh80dCaIbtReTEobS/FBVKE9wiUuLbH
QSF+WyRvwpO17bSRgoIZbx3vhpx4uLzmoIf9ru0/by+0dXqnavJpMLtJApkQM5hc
BETQDZDpXpQMqc7rmjRlyLHIUMEbBHMvOYfljrnexg4dPThEd03VETyXXeA3fngi
YX8GQoLGC7yaf97KuXrVYEvCZCxHC6AiUAl1sEDqBFa52g/UFXxsK2of3n4Qr20x
mYYSrB8Z1aaOyBxob2yWxULpE4p5AFkTGwcKAeg/BKTPb17Ls8ei3GAH1j9HhE/f
q+aTc9ANtMU9NQJH4mAEuEGMzWI3E88F/1MdhlE1cRJ+nDGJoZ0scWeEA1OAm6UU
JU9m+mwVAu//F+kqYTrxPUmPGtsm65vzRgJJSjZ0IKahF4uWtpEfd6pgY9N5VMgJ
JIO0e7wQYRBz1+J5jp7LpqbbRy8rDma/fQWxpTCx983q5QRQRBke+Ws3P1JGbKN/
w2VxMKWeZalv/c+LoUf3qVqtzLix6zbWBU87Xt6j5dsGE/wW3kZ07duMIqyxojtW
yWbynOCHG6V6MYe5AFmnql74caED4j7QEsqBeihibDX1ToAZ2XTWcnAV0bLnORMJ
nde6ale3enNvtjvTbn7M9uMNL2eazjs6rkzOUMp204cTK3IbloK/H5HQ6oZtwL2N
mQX6hLrqwq1A2Tf8Q/H9/uWBkLWwh/BCBIzrBdNgzZbrjOa9AAb/lHwFk5nF2G8d
5OIa7kwLGr7YnKOrqSSMIxWRGnesp+lDuIYB1HEJwKFlt/ReldK5gEgWamfwHsmS
KeoOyIJzNKpvHlSzA9C3qzo60eUEumvYs9LUbrdpBtqSe8SklCNIeWVR5dE/jUlG
6NLVYjC3BLwaJdGjVEHVL41X3tJu74eYGZLUIrC4Fb48wjDb9B/TQ85zZfe87OCg
ILsPF0Vq3NmhmSdA1YUMlpL+LjyAKiM1izicyVg3CaUV5ftC0aIRdsKe35wUfi7O
KSk87WJnWfUgapW5beYlFvMI6AeVhzJND+OvFykE4IBYTzLT/R9z/jskHrys7VtA
811koPMCFOGd7WmhZTlMLowUERumPfc79y5jPHL6MLOqew7guFZKR+KaBT/mPIXn
RYy/JKcxYVKhSdzaM/zGA5wxfhpUP5zdE0Phzq3ReQCkyHYL5FlapJ8Sg3stopxi
92bwAc0Utq60OEboyUXd7uCetdGNr+vukdBayOK5FN+qVhyvg4JnfRMMAEHXCJ0I
76rfZV/QNqP71HQu08XxrNTSNrt6dlCah4fwlbE4xurGgyWxl7IROBMogbncYRkX
YW3F5uLUr5SMUusEvCQxB5LY2DBsGXPyRzv2hs/gpcZ0xgsuHWjnWRJOA+bavszB
/NMywU1wFsP041QffSsA4JKh5jk9kpNjRE1C9l0UMzsI7WzzpFgbqBeRfpZDQcmb
mJ3JBWcdRtrVXyytX77TjSLvD6BP2F2aWJlF+pphC0qPTqWWt+aZnnZqaPTnPQ22
OV8CMrPAYjzxokwphCWFyC0JkEQiRWpYKh8253WizwXjlUwaV8H2ucKi9VIJNghg
a5sStP8cj+3JPn55qY7HK9Wg7RoQzVpWto056oDNu3TN8V4kYs/tRWbZgFqrUqjW
PDxLQiYvCJyuGo4Xs75DG1nbl9YpYz42cqLRKispFcOFlEOdcSlSHSJa+hKdinZi
E23tsMmNcWHFj0sealtjTDtAMUPJRYF8TaIQOwkORcIDlPEyyrO9H2FjprsQxZrV
VvBPipcLO7w1ulAtOizB+vY5bdenliERslMDNJJXiZ/zyXYGwdK+JqCYkHBwklBE
lcTrvZ6LFkWDcabrZSOtI7t+xVYlb71iPMu60F08XosQIHjIRN6at3PSFIssOKsw
PStjr96wJxlhTg+JMTa5/oOcwYwiDlYdV1GXyQS/8Xvrx4lyvMx+kq7HLQpB9r7Z
780oLr4cRg+DFTESPsKoqawDM1fI22hCyLnvUYzpZWozKVwfe5XKANYOOvbJG+Bs
f0ykyRvBTPyxIIYeKIFLrPeM4ICorvAHdImXsl8lRvtcfmW4QTRemexmq+LGGLh1
2jADeGVZn25Csl15AqF8B2q3kbf6RFZuhrlwDnYh1nO7ggWjwJXkZwsmMUCCajXy
RxWLIhtjgWcXlutJhyB90H4QN9IJuWGKJUY0ktkx2taBfliK0e3PD3wMvl2/Kosw
5T+KybAr+TPOzm01xP+hg+8qrVCFNlez2NDEIOBUQOlfpB9h+tzf6EsuBpbc2j0K
35+WPqyzVMtVnkVipfBnPW7Bdahru47jVl2lHTxGKjUj91vo8VoL1uGH9iT9Jo3a
nYD/mszb0BZkz9+X83SdmVta8fZft6UCxxv4/PWpxV9KzLQEApQ+ZhBhAUoHpF+t
uPRdctJv7I+KZGHqTLo+l6QiyBpiwRxOK3g+Rw49IU7kSM5umsPO5Hs1iptyTBvZ
e4BLroew64v9Ya1dJULTYGJLu8sFMg/yj67XOpCvwkZSCxv9FXlR7O68eo53vHWs
srrMbzw7s9SlxTdsFgeTuyjAgsmTccWTb4Pbr5LWKcDm9PnrlvbZkez2bXRmUiw0
asObdaB5VJhTIuKchgtIOgJjT+8uW1GaUFoWIX0qvDDwDCwha/Cuc945Di2VBm0j
wZtluzNFhYW77OKtZtMAj/63bEkKABpxQf7cZMSQwjAH5m/N76R6yS8to7mNPSpZ
hzwnR0qOHizzIoPg2FlNNkQ/7gIwGvXDV4gCrxL5mMVPXs4PNab6FmUBRbZouhUG
eXwe1ppwR3NRSXaBKvNV6VPZTrpTNgiV7pB1baBq30iSW7Pk7BAqwrF+Oz2Qajsd
k42s3mrR/a2HXMvkEurfHh+Jz8QL7ybV3QiR1onNDrwzhNExjYlgOMPH9nIS5twO
d5OdMyJHm/hZYhoqC3lm7LHBpvjzyOK8ccOv4TndTFq86Wsrqjj/K4SZWM6LK2MK
OIdf2scsKRWi/IQcz0gcyvtGZWItdS8kTe9sJ78YaZGLGAV/NRb3xfQ2mK6LWM2O
Lj9iI146dzmdq21A9r8xXgBxRRGa6ACWHmpL+e+6asNtfhfUt0399tku/6Bh2vwn
HaCBgOQ1w21bW6ocEFG8gJYGIVxB0aXAcyBgbxRF5gjxKvLHROuqPmUCuRLB5bcn
hYLiTWDqMDpK1/YBEXpx3y3FMG63sBPFggRB3bNyhaUwrU3mzsD0iVESPkHS9Xoa
QLa9F0YtfRCJdg03NhFq3YkcJ5IgXPj2LYendNib0zd0oO7OI0R+qdX9Cifc+dwl
xlda+1lopPFqz/VhrEq6xnXqSlXvHBv9tA/ir6v6mA2v/k00PLOAb2GjC0CU6yb4
H64F3zzvlocd9Lj6wtZMnBBpLAtWV0j0s6WuVf/+zieVmvanQ3O0uy/ZvHzR4zrF
8OGqM6/piYFt+kjsu93D7khrZVQn/wVP9VJ5ycQ/ppul4g2F7wIGjYbzIhHMmrO1
tVJA6QMhPu+VrjlKMmJFfXf2ufarQ3xiRTiWVHLj+MU/6NmpYph93aeL4rE4Vjy/
Z7wPXfSgx0wAMKmp736x+2GLXjRPZkXst5faaBwud4hHXXTF7C+G03yER1eqf0As
0+ekCXCHgQ/uZiajK7ZJ7WZ+xICN+eFLiVndvXxhtnyVB/Ktb2p+54OZ9PZTY7AA
Dggy8vmsR05O4WnQ3Ycb+0MdW9jp0WA6UIBcmFsuY89UvL6PGwnipEZljHknexgB
NO37oU67IlmRdEAIG7tFxzuDx6aO7xrbwgYg58Oja3aw2QYKnrL6T6ypyJLB8xNz
aNLY+IXxF+jrxtB6gGoVJSFwTCkLPr42IwA7XhCPL+qgbcEYApcxXM4sAX4PGBli
w604pajYT+/ipZ4/lWJtTbSDoZJ1P6n+ykA8r2r5FHuWxoDtHlgTBgNtooabvdyV
Qa3hA2vCog+ciqMnIYUDZ4nlp4x6jmTlaE8c99wtl6teoQ5TOyCr6KhPboQsr0Xz
D0yCTAE/ck0GK09v2wUAVikYvCMsQuD5UXZlF1tQSDTXW/48bN7AhJtsI6q7UKOb
DTx8gVKMhLbR/sRkUwlAaFWNbwZkOFWG9gzxB000q27ikwqmNJDo14q3nxTdnaqx
fPx+YJbCwpM6mnzUcQpD9kXfNZdL5Bqj7MhyEwEBBPNIrpH+i++xkMavctU1FSCy
ZBfCBfaCQGQ6lKb2WKNcBXsJNyBp0FfAcqYwleRs/ptPhOQlBjsSdQXZVuco01IN
cV0agPFjG7zHh1GRIQD4nwfwOA9WnFkTOuqWFbJ622PIExsOtR6wdKIOmoX5JsYS
BOBSXkYjEFVK5BbPiIwGxG2lNIwClSDLrmZj1qjEJxx65m6hdb3trbK9vXQtprc0
8TYp9S2C8zccn19JEPj562ShhIVBvzQOSwQwMRDVOWdONKBu2KTj+01rH+0sxTVy
C7WbqTmWYCTc97TlQfbt/z4YM3ztBJg2WYj4S7d8l6zLqMlxkN7yN/S3zaeetlj8
LSR1jaz2OGrU83rXjtBvdv2xmzlcxGSYcueMuizclWrevqU3V2B28Dl1/8tDu4GV
nrWOxBuJ8TRYoIH8bcsNAxCl94jFgzpz0Dy268xMv/Jnw15o7VDQS2sd1Zt5LH5t
fGwplhGVra7ezHBnWScYg4pwLGQpGfjgdA2tQItXfB1w/yrm5a35r3R8Fk3z1DLP
V2kDYad2jRAh1W5YFhIh+lCiSo462SLrDsBOpgGOH1rHBOKvrznzeHWmIyAMqhyg
qhll0TSMnUkKZqXMphfSw/nmQAPFHRB8kX3VUFwSYneHQfq2Hrfl45dyRUKJsTkD
PdqjCI/yyEHENg1rjnfVlSZkuftpsW1IrgD9W41e8aE631+Sv3cMcHZtiMfgrv6u
OFrFjqMyX3t53s6F+0ITNoCEU5F/UY+hcSUI/748O0U49aVvGcklGmZBbT7b9HKe
pJTpNimqgAsSNUj8yuaiWAdQrP5ei8aeIhBkLzSXfhFbGq26uU7xLloeyYRFIpct
ydANq8o62ewbRhJ2ilM6m5neIPxQheOSbJ+5R3/31TDSahSs2MFk06q6jvZdxsIf
RIlIjoH2WwwML+jD6MGCJNKYNKCkHYpGoJPGqcTtO0box/N4MzteV8VUilO+TjkB
iuMVFgRy9maz8mEEdP/yO69Sma63/veRK3E5d4vrMLQiguwY5yhSaKOiW3DH/zx9
mZwJquvHNu3Vk8TnKeE+Z9omQJeQmaIQujbUDJXTyJAwoTINIk9Dm4iUCikWD29I
vn8meqXVKUK4LaMaUU0yfpogZST10eF0f0/6kcI4kSHN43pJJrphTMyBQkRGRlyB
M5p7ExDtEHcDsjlmaRiuHIB4Zaaux4fGi2IfbKtXLySsiD0yxaTzqKHhWOjJtUFo
6ekoCU2EC/WqeNNiYzXeA/V2FEHSP9vX9vT63PG2wlEVg9G9ferMQP8DG6cn+N4f
0JBWF5NyF/KifrdWRhAYThrpkjLpixJVOP0AZVIpHm1xEj8q/oeQlUOl8iP3i3gJ
a/7nCSRsYgRDOIKwFsdn78GgMRxyCBc0vxdg+OVq3nX09ftGlwWmxxYG25nLZK7m
uK6ijwQmCfDiJFrAD+pOEsWIT/HXFL6dcyNdOxSo1rEU3rJAdHl1zXY6LFVK+iou
0skMoF+PXNKMPKaqIesW8P02P1zczbPK9h/ysULVmE0y4R5gGUs8FAWJBai3JKtN
9c60TyyNNoWDcogps11Z8gwcbjwTgAcZdLuuCreXi2I9sQwakaqAuzJXYSIabAy0
e2atT+auDkpp4ougtaREf9GjJmRbTGo5g4yQyei06FNKaezVeEvBW7AqsuStmFc/
UFZn4RmSHG/donbAbo+DLCpMBZZvd2mUM4VcJEhBaRmeIQXj9t/1zhzU0H+Nn31w
p8h3VCpyz//sNTAdaggiWjiKVcH3b0RuJZ0eVp+ZR6H/clLTN/8Ivv0xX3Ezz0fG
82agVAXBPbn64WwTbQKqqnI6OLPU3ummLII7TTwdsVbGt0D+CkdyOEtA54zCWB5/
4wqRM0Y/1UrhQ/8OvTPjfafJO2tonmkQC+YVNwzkMyWRV/lMki1WE5DNy57NRynJ
2x8gYgTgeToJ5cR05cpdHyqpzNTNrh1zBL1XnxROrcFZWZsNSssm95KAWCskq9bi
XdWXabR/dcF7Gk1/oDxrdWdKPk863fiW/2ObUpNsqAD0Rsq9vsCRDH36Lx3Uj/N9
li+xUXxw9SJ0CrDr2RmwTYV/bJmDM6vujX2/33N3zDKhMILXUvgpzWSPtZMA33Sd
UFFVdU9amN4LXuyHSH7ywiKU29M6gNET/Y5+f6Eu6f2PSIyEff1c/TWNVBn6tJ9I
oitgwsTA0nek4GDLh0+h0dRUQH6E386VoqIwY4M59Al0CvR3EW/7DQwsNUeKMnyr
YPJimu6KigU33FJgaHWcMwWWn0ZCuEVNC6kcx95AwSnhUm/P+YkRDC3qbpCBYCWs
woXPWwymTGSfXdfRA5vZ2T3fXRZXfCF7JY2WqNp7Y1k9FAggRjWp2H5s03l6W+cT
e0vB8x8HRmhYN7XPmsybe9Eb4EgJQDJVMpObxFXOC6b+dhyR0835uDnjMXRYQWs0
Pc+T6Ux6jRNG0cmioiei7Y/utKI7tgCRfG5aMGTjzLieitBZXtbVqUaUtH+xhKqw
ibK7m/Maijl37aHUDaN2JpBPZWA2HjsKwN6cixyMuHLRvyT4THCM/x9pCC2CKMB2
S0/0auMe/F2h6ilusy+RiLfybgJZGM7b//l39UaurLmV/EzIGPoYzoaX0VV+OY90
S0+Bzly+jf/BQa4TrZpp1NywzATWi+FGhlWcKq6xHZQKqH8xSCKo9m7hJPsIeyU/
aQFaDqTx2mMTKM25XvHJYH/OlZzN9Xkhz4KCPfjp3hCujzfNVCMJqr9KbmdC0bNF
3pe1G4kN+sSpfvYzsCgaBwL3QbFWAu3oC2Ea77aElP+eUo+gkVhmbMToCPvrJbY+
50IbQEXO28Qy8yJkGosXO5ZnMBjbTOq6K0nfQJDUsEsRVndvG0o0OwgLE0jaQ39k
qxUc7DIESWO43lZxALqmW3N6O0YkO8n7v5SKLU0oaO5Z+3txld+M+m78YkEh8hZC
LG4p21G8zHHKPpChjNXfnvlPFFKuuGO2t344CydowmPdxr0WO68PCT4mEXB0E4k+
VhBc1SHGS1d1dKk6VVQ3w1xVBNfDioQo5U6mtAtvu1klqm8E3BC1boGd8AGPL9q7
iTjRinEfcALxKy2Bl4T2hOsoOdnMUj61i95dtZ6b18wFmwn/N7unljT1Yjrd/qG6
aeI18HSgosN786Zt8y960mAaSaNOgqBQnt4QPoWdBafyXIbS1bXZ6CSgIH+lkOQX
iijR8ApUIV1r4FG5wBE6upTBs0wrSLwD36DbRYsE6yclnQTMSKaYJ+qe/03+ULnq
NkvkRazjDm3WkY8N1YrmRU/Wzat2pyybs7/ywvhga9RI8lu8Pew5tvPLsksNkrEC
TmgXK5c8UXsr64kYiIyvVxoogChJDrv/KERFeNrplhwPwHwHKF9l1nWnljlpwfer
ifOOYt+w12NOSRNOHskWxuxTpJBzBUYOSRZDXrSssd2OBSfGCoULUAAzhhm5I+Gl
RHSbePqkAy5UvrxA/BjlzBWPOpnsaxdwKl+hFLnlIrrIpZrgQ2RJKC4y+3VVlSCy
Y7T50jvjUq3DeyDb16uUEgCBMCKU0pbE8p0I0V/u3HpS856i9MaONKwtAp8J7e7K
ZUEAaOWpBJ4wRASJjf9sw3JSbCc4wSkfOnfPppof57tdqc5dP2GntQbbyJ/XWbFZ
/yId/rx1ggqtccqhaQJel9KtKiIUIlBGuIKIv70zmJUnmhGpkh/PweOqLn+1lGxD
4NAJxYXQCZw/6QkGLR29ZFBL5uL/61i4NJHej5Dur0Ag9acVFI8zKxGkgKZJ4C3U
O13eiAVzn28eOeoYuFe4tZpR1euDEvpaXliSZwaxhVzEoleBNa0tsVo2gVGbepII
ZyPyGqBuznR913krsC0tDcb3ox7xuMYJzfvEyJBxp7nN+oqwIwidlnPPG6KrHxcj
M+ENeCj50J/Vix7QvhElzq5TTRoni5vAWJZOxztwmDOCeFipYEmGwEsvoWwwBDiR
My5tBOpfoA7H/d11zGUTDUs/he/BFd11JD8l5mDAL/1YbF8tBFo51ghqSb0bLbH4
brHXhb6ak/VEEtphJENc5a0BEpbZjx+Rj+pbxbUdSmLna9xLBa0dh4pbFMIgqNRK
RQcPQt5J4AtlAmp9D4SnFHiQsCOUX69xgD7jNNSOqjLD4QeQPm3AkpGDJbRuW1Xs
9byPWSa/SYJtm0lJ5jR30pfHGS0tJdyQu+osNeJ6OjFObrUtqX01RXX/HYDkWxsx
X9vV48BpHYD5aR3HXal8It8FV1RdhD5MmseuUFsWEDOwK88L4Br7Nv1J9VY2Byfv
gEgfUG+X+Q3DVLRAjtqFr23pTzvtnHy4C47KIoueU7zTSSufGbFs5jBlhsDJltV2
E32oXVzcswgK55HqnCA9NAw7ibIs1WCU2zD8zNB0P0RV3KBDZ2yn6DpH/Edrcv+Z
X2GOinEjg/hjYkdeRMvV1nHWKQWaAmHIL4PB/HkCTOOztX6Q3Y+cTH3XSQnuan6f
EBSdOlZDQal9HxHIEn7mMdlijtViKoIbZDTXe/pqSJML2WBnRFUovHsu5HOmNrHT
JzApE39kK3xKl4wtdKPCxxVR70Q6sW+BCBt1hnMRu5Lwlv/8l+4ggN7pROLEjF41
er9NPOlAnN69VUYvhNEiEUCXAtqR8jldMEmalIHhcz2A48EzyJjBa9zJ+OS5hpj5
VmDd8XrNpwM9g4mbs+3Ko3mMnHwbi/6tskt+/ohy0vhtJeNXNokkgLm1IySmyyUW
HVw9pzmeD7CyApiuC9Wicg/dgLQC57qdOiODoabnfvHc5OVzHpL5fWMxxqDM3zfP
ZcG5/xQBMc2X5emVVTvBCe7aui4AsA6xLLp+5N7eNT8qCARnbLtS+COHL5vYGWVs
RD567sCbvUdXdyEC4m1G9plpAX3hhw1KUHxauyAZAnBpRkdItmGYW59WZGe8C+j8
VjuAeM5CqUZGgQ94rsPrdtBhN6Wn95ilbskKe7KNJkHpbwjGUTwaCYLKOufy60JG
ZjWOZ3Zt+XVeOy59azY4WXAAD4E1t0/q8p+6qQC8ZPgQtI9V/fl2nT4/f5ZX/ggR
xnakkpvio9Qj2TfZE58RXaOxiDcoSZGuIUcF7XkVMzAe2SLR1ZU5NrX3OSUbp42p
o2kDfWkgMGSruepF47MTlQF4KBtnPzwltbMLk3ljQHVk4AcgK3o3PFF4RmUN09rJ
PHy8uKhEFn1WdGqJtiQ2A/fFvU2QXNTtOinh6ZxMZ+yzwJ87l8rjypEiVtAWT5sW
Mnq7ngkal+/9sk+yeOj/ythp8QFSXZrjTFVDsFHnVH9ni8mTIFl6KpLrlEbZBtSy
scvJTJARUUcLRFwlh7FHDjzhxiWssVIueNRtSomg0xuWTfh45gALPnLbvTSZ4Lu5
YXvd/xm3D3qH6Rv9EK4MRt46idAr59cgWImSb3+PC0HzAXTeUSKUW8q63jaxFovk
zLXSnc9NgGxwJ9c6gjJQiSF83PQlURx01sT7fdta5l7V9AXW7sg032a9vAmGQU0x
KfxWVaEnCDHIGaNS1AdlG08HOtTYB7dHIZF9FUa3SDT3WOOfTsD3MBkBHNTsfcXS
drJfylW96zDmTulz3dBhN41FzGiAlz8QQsB8P7HHFEFcktt7MgIpUESh/ujJR6ZH
ocduS2liwYVB02+AjqZjUp5TFDzuUdZhmnyAnuNbluBIZza5V23VFISzunIrqRWT
83v2bwdm8/V+XnMUSjKNeQXr7KkxHXE2qiJ7UBFfUc3c/EQhxpRGm5p5Xybt7Gzi
THm2eWFcX9nOk5Nda7N54Cx8yFGjnhiyBmc8iQnWQFboO8Luc2G62WhS2DrVk1CS
KjoWCp+5VgqDIOE8/8xNwM2xGC0Bjg8cSH9L1dZJnLyd5oFYbvqXr1PVVDckdy3V
5PR/Urxj53FNJE8Fs3mcsP64nmqw5i/X6XNLoVohSUG68TA6FOxc/qeT/BBEkHus
XuzZuX9tJE64V9XRoDPjQnYYZgWe7OSB3aj9G+o/lkYZu8/T83kmWU8ThyRUH8ci
z0Dkt8PpQHybDtYdY5e9M2CH1Alf9KJ1rrt5dIHBUgXLt8VZh9LNY3Ir2Z1RCb2I
IqGFxt16+0AcjWqWIpVMjyrmRgCE/qMmkkSQCGAI1uaRtwtUJ3PSwvNxHXRF+MyK
g6u5khKhNPO4MkF7EO/IVYT8h4dvrkroQ5HMAfk7AQa2XUxueK8VHiyBwAXLmg0k
qz2u01jmggjhBTVK2Qscv95StuDBXfsVIonQN9k/d+waSps27vgIPpK89A2nNc2K
RmfxBVJ+P8Kz0xYQUfnZQ5c/kqZQxiDvnp2Sn89PS5JKV9bKnVxgQHO7RqQAJjf0
3HtPVdZs96zhQrA0/clU/z/7D1AUiU5NeEdFu561NqTPHtFOeLOH8fpbZ2/vKUV8
XZQmFR4l96aZP9eWCYXczP9Jl3q9n1sIAS9lpm/fqkjQxB+224kV9V5VB2cs62PK
LYuBZyMoWQ7CxGb1ZHsZdFfmcgzBFKSIyI8HS2zMf1PO39+RPJEh3AVtfMzXWbDG
pVZMDyVMmztotrYDQrndJ37T1csfYxURpkUDkY4aY4N2Lb7oNAAT4JCjXgVagjLU
Atnrz6zkaaL4tV/qopPudrWLBtpUPSIGq8zJrI3p3u8c5RhNtbjOX/u1yn+Duy1U
V+vY3Pth689jSZgk+yuLgd63E+ajBPLGu8YzvSZ9X5M4rtlKUhgvngt15q+qSRNp
DG1sKVznsAuDX2hkYyQarFg0KJ021HZMUTdMzazPzSBAq9VolHX3/kKOX8WRhr71
23NEXHMDSfac791L42tts5MpJbm2u+ib+1cNPtXfhvsihwCnHYxqecBvqdL1YvPI
swlDiPa4vLSo3d5gVjbHRE9WgJqpa9OosTD/k03S5NyLxcIU8hOQaIXoaJixQMj4
+cGKYrM6WbIpGuEO/LVgWx695nzwQohI9hTqNOHUHjamPU9YTuBulv/73YzYgNHB
vik4vHuPIHUKaPIUtkHKQ46Jec5qJCDGrcZ6ADXI29q53uVxREJPBvO47I5RVQfh
LgOgaLr0nZYFvW4rPJrcw+aYIP77ycikgoBf36W9hVAz76StttcCxC94Gqa4fNi8
Ld8DzfMXEfdEC3URAZOXleNwfm0kOPwXhJlep0q8tiBXN+JksDZgt37n1+haEsx5
szu0/n5laUuWq8kSxW7+sQZLS+UezH7uusqGU5yN3k/pEe9ZrtRN3kwrnMIJIz5U
0rj+DoxM7Mv+OAX3OjzruDBiPqQmPJIXKRZJi9ZCS9B+BwNdAfQs/pNJj3UF2/oY
ai5xwzzkDOfryaUfmvDHTNy8xxa58Aoqsxk5LXALb6RZP5CNxWvhePIyjMLK5/Dw
0iwvgsmEM7SDnxNIL9B1T/iXy6MmJ+O+6ZUHoG9KZGGvBXuGcgmaP3/khfrQ+U6h
E3DJ7u3HUd7vNVzf0yW1Pxp9zabFuxMDM01LI8AxbK6jO99fjkK6MNsNfAKcIFoK
zVn51cBbv9gjbyxVq7vTqSnn3wWctufLqiFA4VwUozovqz1hBDX+L1/NNcXy+OLZ
pAtDn2p2ccBwQohVNEIs+bcIULkj9bTfEdUHLuidLM8NPSa1vABmxulGnqAtda/h
wPvPhT/atHnEGqdlddAMKViR1/8LJDiOyTuT/MWAbhr6MsBJpKMIoKAOtPX2LyyU
ZdHML4yrzYwstz8yqG/D3oUY/r+l5s/Krd3YAdyxfMjE5OSbY5KU55pPR2byLBPv
lzZN3XQIFcIQcNom58WzmXbTTguFt/6FGOcmB2MGARUqyxS5qmVvLiJ3ZlRohl9w
iWGphU8d/o8nskJnL/sCycxnyjz1bq0xZo19aTSlJgS4GRmt1EfpfaFQW9vBLHWM
lc5CutN9YfkCAjg1XeRN+QSJtJXRJb7PLfdwudmn2ez1ZrzLphaw9UuylJmaz6o8
bM/6KBkpBK/Ehxyg31h/auWBR/L6PDau90F0g4lAC7U+Jij+QxzQBrSZjkkrUcJs
4gNL+Mlt5pk9D5eks3bamu4pRYNjDIWhyeWgb6qV2Qt9wWXYGJawcpIocEBqeEQP
cOig4fzYFB6Fw9YsooInXoRPSmCRUWb2H/NQlzK/rVrSSTfDMG1d6CL+kj/mD8J9
B6+U2s/mx/bsXei1ZZk5wrAE2If77QzQ8zGeW9CnH3/CmUnqNbXB2XnmMd+vPOUd
Td7xprHCNG2rO7vrF8uSXoadpHxHkrgPJDaxeakY2kGafuYO4lwggzfu3JR++4H3
yF935o9HLj1Ri3NUqT1Rgp1fP8gptEcya7mID3y/2spDaaMd6h2dG3DkHyWO2pht
xpUG7p0QsjJR1nRxJLxTWF1ocSwn8iotzW9tHv//7pO9xcKsCrGu7DCyzellGHSV
AIiRaTtJ9ObN53au1ULEgzhFdyoJG6Q6qT+1/WbFpkemQUZLEU+B2v6H+atShz8E
ejBeu+QMzR62OeNbG6Y8SJLtxVPEegz6H1gcYcula7Ni3iFzD/RlzVspe4pbZQ9J
JYly2urtcDSGtrpthI8fchXV9xMvzyDIG0AQOtkQrbwWfApKBS2BPaoFj8Rt9xps
4CyKG3mtV0qY7bqGW2H5UOSL+XJdUNWVK0S/AAjOBMbeLsjbS30WIh70ZytshHBf
pxrM6DduhhGyB7syE8jHJfZ6/MfoZAJJV4mbG5g2MlQjmGzOTD+EOcf0jed1zHhq
JUKMgpX7xRyE68OMkPRi51sdxUo1BRDCkJJEgp835E15RPANFhxhodTMy5zf2jSB
UgYI2f+dlg0904pRmcu/szZLjSSrN0lHhA5x3+5MmGAshsDO/RBBK/JZbjVH2kqn
iPqxLCBfeMT5tFmPsYu8e8mK8PRtZj2KQiDmDiqnxfbPvTZa8A6M6kI/f/BqpPSi
2CQIa2Gei3XHZLyHnn/g29vjn5OflDxWmLa1O+07u4px0wXAHYcJA4PYinBbhSJH
5UohoIZAAV5Yv1WHbuUSpaG4dbHgeQvdn7p0+7pIUWnwUQLS5jSlzkNsbKATFg/W
MFFyowHXcqpmjEXTpaDiZs2ih9WzwngfyP+1Bq39q1PVsBwXgIfiue+5btueitls
eooLxzONJ0CyPeKO7s/DjVebdFO8zJMi1dcLuaL6JmgZ5hhq8FC2PCE9lqXActy4
yiTcBoI/squpWH0kV7MjSReUSyDWHVZcM+CaA0UM907X7OX6ihUqNxwaOivFMnxB
U2mGJA2UihScyWUsjFCybMPBgefEemaY993ZUgMHKrQTR6rEa5MnoFQIavheo69y
P+kl3cuBf2UTzyxzt3fUvwBWBy8n8iWtOk3OVEGO4N9+/k57wC4uplcY+ILBlh0I
7c8YWG4gTHiukUt+h2OM2UmhisJrxZN8ov2bXCW5ynAOW4TjlEmTSNo6EWLf3jmZ
8sEC14LEFVHx/iUPOoTqDlvhqS8fqzlALh42+Epld5FkHTaV+n3mzfFakso1UTXI
yqnu4W+rOheMQrEYLcP/8myFE5PjwGCMrkqG6SLxgr8wWzY5aopmOIC/qJLJX45C
K1Lh9aLqIUeHZpRy9Cl21e1cav/KR/E+xoQEWm4LubxaU3ZF7KkFa1nJdNcjUMzu
OrmPrBHijuHYP05IugdSNko7Z0X9dBIw4nJSg8YuUR2vQvI3F9M64i6n4kYuKpu8
kQzRNaqnTc/q6qcSyo65TmLfELwHv9hr+Sx0t3brsW5E628hIkFKwshic5DO0Otj
g9LascqXkyqozJk/ScxXj58cxAJk8XRrakUGKNId/JQYUuMuysB1/m7+icKDPmui
/FeEVqaCaCCj04AKdHv4qc+NgByASYyoOcCJaJKEgJj21sJP8g2CAOPIjfWiwgHR
8V7Oq/yg7eJ6q0d/inqV13EWaE/259U1fsnS/8v9eHBiUMP0xkjDmtt3ChHeESik
LmhQMGubqDTBuhhDNNHqG5WqRuIFSv04/p9Dny9BAnCies7dhOfYAX28/Ahm5A5d
M+UdboDXXUGPOKtQUkjbQL+j27TAjrQP+MbSFxiDL3dhnadxVXby31wrvomMstB/
Hxu5ol8DAR1TiDnQFQgQv7oPQCuzC1+F1I53YXejTimriSTUOyvSpvCafKOsHCzb
aE6N1gZc96NElbUWM2pRS0Vr2q/os686UNaLxzdnrT0OtuvB0xEc/7jwiQpJw3LC
U1EmZsFbZj8Tczp5uk6MOdMsCfF25GbdITgtQGCG4ABHqRlSKMerwhaam1mj20gm
PDgo9/cviJJTNcYCHjsHGU5ani4QKgxqQS5ZqutpoH3/st/HanSrMpLMVyNXS+Fx
AC+cgMCHVtc8bmtoK5ej9gCODy2p+l8sOaIqB8s5FjowHQHluLQ5D6xVPEAe918k
5unHsJQdpyzNPbjUPzoLqfJsHIgGg3sXeLj7qrSUC04FxsPPyn2vyD70HcQ+AayB
wYlqRg1EzQDShboA9FLFhtl0X8DyDAi8NTIXvVh/v6NKf1uOwfeKWOR45UBy/ZEt
fKTrHZHCB8dwRKNm40dXnEHRgSKoZcsB6ozN/zLWomeJ6aPwf73mZ0SqdldC0GEF
804coyuMDYTyArMWRjggU4MuhHKKNXc9idpb6t7K3hzyfdkZbYZvTp9907KukLN9
wCLKWVObyyUTL+Jxthw8HJQYI/reIE12RIuZMce4rWEZSpKir/0MmZhcjOGZQGte
lyIi7SwoZCB+HubBoGd+nF85hy32LE3eW92wGC8bWS3VZ7wOGjN0DW5yxNavHmc3
oRynQkCsyf69ydMkVzbbok73DCiMlI9a4rLTolo4ePL8m+Hqgce1DiwgykE91AYC
Ts1oHp9RpfkRt8j3oqnIwRL4TLme5yKQbQvAKEq916mXR+ASiffCxp986n76H061
VZ3A+NNXNtAGH3tycI2ySMVKFAB8uYOorLjQU4QZVTMoCN4k9/xI0kRNk5d++6og
q2BNzoO1AZuaFl7MI42kQR3eyXPGcsRXNTdMUdFZLsRrfJJT314JuJIQ9YkMf6BH
A8Ek53zbJbU/BcWQkqr36IvzvHTWDDMiaoIBbTz6FX8AXhfI2YztqhlW4xt9IQic
kK4ruAOUcbdcH1T6p3h2sI3TptDnvKbZs31ZqeRM90juGUf0iC5ruTJI79nA8ljK
txRD7ImZ7mr357n786sAV7sglCluHnvGXdzisM5ztflMaY3j/GnxkteqnG9qGvwd
UZ/aWkjzPxpi1mYAPNk5rJkHUsT5qxrA6njKn2NBXxly0QQV8pKz7yITKE3viR4l
lO27Oh0A/KCiwNdfNw4Z6e9FSWds7NDVQUYbgXBgfLOLvNwZPKlC7JE6abq09H14
pkzsnkI2YI/k18V8HVPDwydT1pAbAf6GfwAOcR8wpIAVixkFY+bYakZQXpJrnaAN
jIPJd0FVTPUpnQom4pLGXNZPS6zmMJtAOIFz70P8AXKA81uQuthgJ+ZaeRRrYthr
9+9HL2iqXVOh4PzXZMFOAs/gdGtLEj5wnggkW9dbfxJ7udY0kZacJvnGQviHxtXt
OqU0/9adOYIjlP3Sae9vJIrGbd7mn8Zbg6oM2kbVf5w6ww3mG6EV2vcOQjoCLfkq
0BJTNaa9J76imlBPDc1iFR1oV3HvJ8QCKwBeKJOeLEO1S2B3xveyZL0cUQvaIDY0
9C5pdXZWlZyPo2n+fuNKRuu7pgKOA1Rm0qivk9vKgcuQRH15XyLyErwJZ1avVQ7C
L5SE9jWxw/U4hbyYsxdIslbXWB8Qh912yS54HMZtq3StJ/xxzc2oV4oQ/1ywALcB
1fpiH09rOzpfBuF08tu3WxapOgKVfxV++jXV471C2V3nygCFaX+bYQR544gmbxM4
2l+cXrigvH5Z92d6wGgjbWxpnQzn0hpvyLQ0CEXjPTAM8uToFY9ugEIM8GiRFrxz
DQ8p9sCfNQm9Raqfo0Og7vtoESELGkNYgDpMRWOzXIf+cov8XNaWjSpKT5XRxqTZ
5UtDPePudGRFPYUF3nXOr8zdQVtsYA8Nc2LRe20seYpCEVjzUX5Eghb185dox06i
cYy/BVJm2xeZNTguzr5DgtfKbjpk57+XQlwlt4c4derSJyLVhv2LfJaNGrlYZwzu
08DaNkuXs4yFAYaLIsi55Ges4BKzhluxdk7mN9AcuyEDkKt2BN2BowzjatO5zdMh
4tadu73TaD3E+YzG0Wtj5b+nQ+W6a4ohK8Y4kC6EcBy8AGas/YbXOdut+aLL4xve
SaoovkbffaoprwW1VJQbzesKoHZHtGNiggEEMRd0WX9iogMJsCOSfYKR32ISjg6r
qZm3aIAy3mf4LSGBxfJ3vGuo+1vu2fQxqwVW9i93LLHz/cXPjbNXbUTpA1T2vjuJ
B+ULIxgwMcww2yX1MW2aouyBiVQxepCFq8LOF6X80m2UB3cxJkGduvPe7riJVacg
6hCR5vuXvXbFDQ0PrxcpZhWRHuQfzU8znrxuuBaCPu8G2TDekKeOd1GXov0EPDi4
mM7jyDsd9RLEim+JeK1w8Uwy0JAfaNeAGkNBT/6A8+DT92LgPaNNZ0TUEVS78A1f
JQILpytSvceFkT2oC2FH3PipoV8tw9d0s5SbmNYBA7L+hw+bqcC3Eb+nEtbSiI2Q
5SPItsjMwHaAjT3fv3fCDt+TbCoSDLGge19TXVktl2lkixEWvWY2Jqf77CtbA34o
Q+h+/WOk50ZLh+KnrNj/q25LR6Uflw5MjNKjcU1m23/GAMStkKyuHeFCitPCFfoY
E28zWGhLZlw41QbEZLfhacks3xI229bZocN/pN+vKr38hqgNZ8Mp+HTGCj0kqOXo
7DDQSJEC4iZCiK0O9WycBGpk0Ichk5NuQ/YSLeHf90cig53CERiwJNlDAit+ilZn
Tu4YQvP8ZCdBxjUPelJLeyaa61OMEFc2NUtrP7/9TA/DHSWrfzYuCpkUql3Dmg1+
tPZd9DjbB1Z2Ga3aaRXq7C6X9/nOyCnea0VOntE0ko2OlJycTF9BklMK4M428H54
o4BBU0U4j/ZsdqCVOM01loF8P6vPEP71QW5RVte7SyuPtAMNxix72v1a8mqRLDS5
3hxripmvXroG8Vw/8fSAzA3HQlkj5JHXl3T9QRvFh8GApUakOlnZT4TWlb2XsIq0
SnVyJNRkvhFnHDDThI/5V5cdCjJrRossmTQn254+WlIndkNLAMagFDqBLmnHXPeb
2wcY+SHGObaopxZo1SYFMnnZBhbxnKWGlLStPu/SuJYQfeq5/TDbGpw1Kp7FM2tF
2QHka92iFYDLo/j4O3wVli8yeQJricOeXckFjwoAT/YUx6CwDx3gMm+fyXHKh8Xj
gi0CY/wp7F6EB625erMXpHKKjhLbbQ8V2HRx5stP6IT93n/FPEJeg510Gtx4wePo
PH0friwmEGIbNkKhSMBsrKRMy/zJGD/AU5P3/qrg8Nb15uUPIKmA6c0vZGA1tIgA
bvxe0DqHSLKEAfxRv/Sl+voCrdJ9AXATrMxY+opPM3JyYZwztvZk2DoEiB1Q0fXV
yR/K7cp4/GQUBcNRunfwXLXwMB9EozDGK4bjDKkueNC2j5aes5vUwxgyuQ7RIYH1
r7Rc/0dpEP7U4Qlb319889JNEZMfCV7da3fu/7ObUKFF5nBsrEUwZbWqt2HdStTO
Py/8Z1DYKB8XcDdHvH8iJcEJJM4U0hZOx4l4cMwFRv6d6ey8AhIqp5T68s83MJ0P
c0kyWxCXsrbyl5TxeDXkGyOi7GXFVkNnqjGLgom2HRmDDb555jPxpVJtWL2BFQY3
3s2+Qs5ElfOyStOHT7KhiuNYwa0E59EBayCsBDgq+/PGDTe5O56doiKaYd2T+FMG
n9KYXo31jbs2lmHc+hdoisHtmT2MkIgNn1G96Ej1lsp2bwnoaix9dn0w32slPRCl
przbJA75y+cocgs6MyLIf87t/NotstK+sIQDqcqO37VdKp6QAM454ls2Cc1IiP4Q
t3+I36qdtIg8lVxe/uNcjy0aReQXsWQ7oXpZk+2A/ExlawuFumnyDTOhbSztBdQb
GklLcbBHig/mBZeGji/Wvgx1BAZFzRhu/PD+4MyozMMSU2MDgJmzOdTl5xQP0PFN
2WT9aLf8mNFhrvGj/Kq3PH3gJ02+H5wf7hJF2FrVYukcK7mSTvFd/aB/Cw6NsCUx
gBWadJiySdGzc1pjChPjiJzRQw/d3kp7NsiNvlV66gQM7cha3XtehAgPaXnzmipo
bw7mtx5C43wfEvgufqyh5LmpX+D5DE4ta+VlgVctwmiwTuS3Q/mYSJIr3UfzslmA
ZT3wtETxxfFm1N8cR4TWOi6gi2l5FeypQWmi2y/pqLgPIsqNqaNobt+qWWEn6RHr
+iB3vOuqdBGTFdJUmv5e+jlWz8S7nv8Ghl4LKzMeHERBXgG46wQ9I506eVAg4MKK
e8k8xMdVhA7SbJsWV9Gc2F704P9Eqn58LVS1hAWbrXylG1f+JzWyjsZlRQNhO7GY
hHi6tHGYDvgW8n+1VejPvm9Fj54h4phucQMdhADG0j40o2A4YPpf+bdx+UunOBxn
aVjW+gEJ9RZ1KyCy0aqSs5xq5nkuDF5o93RAI2JPgJhD50hmEr0WhZyNm3zkWOLo
rn3iqpPUZcBL9NtLqK65jHlNu0TBaP0DtAjhXcr9fsk75AHIPkKRJRF9zhzRdYDw
iV1iavVeH/vSy/DNJoUlJmK0+vu/tyun5KI+Q+TV+LduFN+oNAVElO77t9hmqRSo
3X2qxVXVsw2k8syg4BTZ3BRH9yKmQj4hCsBqLR0rwUMa+CqZm9Gv5ANsC2dnPhhe
7fHXFf6C2jjR+vc9psh0wi+rHHeEZZzz2bi9ba4G+tVFueWdUMZeyqBs1CxfmRUR
eqhr6U0G6FFZLmtUop2IfDEEqXnCqrIU2j/n3YmjyIv9lhfEUAT5gZXSoVbqb/Se
lcxxHpQyjC+fr0QRGG2wcrpNBmTivjPanCy2w6oYO7PVsq+wOtvar6UdaWx5JjRV
i/D8gp6cQpFSl0vgqH6BySGLujoLigniXxKxzflf4llGz2QPZn0i4Lh50XiltNpK
BwJSq1VoAM9Olm0zBPnHq/62T+NQFnmXr2D4zt+9ZLgLZtyI0l+rQZ44EjcOXSDs
xnN8llL4SZ77qYOyvWtPFRnZJHitNMvetJzXDZdOQiGsIbm/uq0l5jujQYdr+tA3
crj0gXZczpgrdPSLMgmC6NkdpqzVb9UfEtcC+Erd1auzsuGR4Wr1JBNnCyMpyXoH
NtcTjak9MtcoPM3CxmCFWkZ5XI2E12Z+TnIwJ2xcP5k8R2JHN2wvZPgsjCf0SuQ/
64mJ8km2JNZpEawrUljDXd+Lj/vQqCG4DBJPwaLxrClCskYX+Jz0E3+a1E9hDIGw
4pPgrzoy7O/Tn5xhjVxZMMmtXtHbAvDwsMX5TkVw7O1J+gXRnUlVhBB7+Cr/ArF1
HA6vmwbM3eIMWDjv/bUgLRbXumTyIt9JPtFGg26KP7b4/dAoKvLUt0GekV5dlKvo
I7rqiWSpB1m8A5Xz9bGdc4Z2CXCOSjOLrBxK45rNbu0cyhfn39v+Eyrf4mGzMeRo
wghyDzyKOMyukrUZ1GbkVoCvJf4LrKUE8bNqUyYmeUOHcQmTGEv4POfX0Lc7DSLT
1pfEq8NZJGdlPeTTNLYytwPoJQEeDzFOfhRaP5fphfr501DUjrkzPAjSvCdmOUbb
sDrBgQ+I++oHv3488su3znOhsHuof6KtqdCocHbJ9qlzKjGNKSLrUYxwan/lLNa/
Q4GZD9HX+9zOFWnyF8lKu2+OsJTe35boLgnaDzMHNi+3aIUeDHcycAAxUH/J/irP
WyS/b9d852a6SG4Q0Fdc3k65xDGuIBFTY1Ns7JoZjAxiT0aoRSeZPUs2n80ev8uJ
WhDx/kIfbZs4wG818x4qxrBhuniyXEcinqEO0uo6YvAFpW/o4KfD3YVcbbzK11MS
d7LbiH/LQ1NL8boESZeHAZLlrSDCf7ojeqIptajTKojEf6gDTNrCafr/Oxai9rJZ
MY4UO8ZfACBXtwCq47tqp8iiI/hWORoIg3i3nWBYszQggpkcmvGDbcZU94vPhs2T
nyHysPOLApuP481Q5t3HU1+uxbPUTYW4lGNbMY9Pl4ZJXd3o0mfuHfP7CePndwHL
wMbsqBVgQgEN2aNzAQ0y6jeoJSFVlNirwlJ7vFE65VJlD8+AYgY8fNRzGjFmusSZ
lmrzr4AaIl63DkQUdAAq5kzGBdpfWuKiMaTScw1tUZC0Ebstn7XuOE78v1Xf1zcA
XS76S3NwPiYpHUkOMYzRCiwwe4vaNVLRKH3IESKWqVGcZen9XgJOr2y1JN8SCu3V
7mHBqWf64vLrE6GgJ9VmmWz23RmJ6MoEuNGkT1GtqSi6oa/h5I+iWpA7iVr/lUgJ
2eI/n80XAdEWOgN33C4XS1QNQ9KNTFeDdoEuM0jzZsMUgrxJNDVQe9MjMQ84uiGf
OeSkYoKbVKwHyV5v778hwxRF7tu3d/JfQro1HyO38jeHa0yu0DrpbxB8ASHx2W90
TbrVuHtnbnlKj5bZfgWoxEVHinsFdzxbr+dL1Cqu9Govb6w57r/4f3GObQfgBnA7
+nF0CVETlqh1wwWkTJ/St3SftITmfitAD4tZx6/IWAw4U5qbk07o7b3hvwIxDqCM
fB4vDn8S6C98cisIP2ozSSYhTsLj0GPKA+2vhXYYbSKN6cAPrAVgeuT23Mu+tqdL
kFsDvgVDga3klKY7ddTbmAE3rtNIZlQcdRqmV0BJYYqoKeMHfig4qjbPbL6xApKJ
zvD11FS5/08bua78nQu2nx9stKnF+Pd//GF2GgD5tHxzqgkzP6zUw+gl/k9HecwG
WN7eigVAdWUu2rTao4xGBeU4BDpe0U/MBXyq6yQ6oNPAN52KIpmgHurLlHLA+5aJ
n71011t2887bbK403Fs1xxGpIScxRMUlqfAoj+9ucPCbZL9JASFMaULCSwNlXvr5
wBDiPDlT7XkrOGk9kkxHq6h+zlCiR0YOsL5aNZpvsT1dBSgatmPILVV0rQPH53xE
/JVPRVX0wMvEInvfxIG7O1+gR0scgJGT6netHrXC33jTlUH2tJCQbrYa+2n07woH
2A+GN85Ia80gPI0HpciTl9aqTKGnrWEgmCmj/uoHx3+RwIn5fLYpAfI/kxZfuJRp
XK/MZfIq7bv/EHmb5TBhVwBx2gKLM2RaotIAx630jHs5cdCRN2b9xumzXcLFVggp
gBSReaElxdTrZwgMrjjBUqfBuBQFhXRHwCVDOYzKvsJpvuqo/R58vNgdkZm93CxE
bOIsWXLdcr+TfkwiaJfR8DXCCkrY3SL0irSYKGo+ZvnGtwG5b5RsfbQCXRcQcI5b
dmQTcytfWPcGt+RgNAQ7QQW0miVaUt3vhe6YrK/e10yNtP6JxeU7Y7SmQeQDNLfZ
Hq573Wkpw5xVs2fK8FMHwWeudbTofaHg7VPPHpiD4II6IAuOEsx3SqKscC7Pr24M
OnMPwDFBwjPQvnNPta+M2k3wILcVBea884mmmx/pd1kYO2TBzHAppKqAb1lDy88n
g5F5EuRexlsDDao2U5o7Ff56CstOE9RO34sly3ToiHiiCAc4vsMUMEkpVWKwvyBH
jDIvxZPjBH1+bzbDHQwVRzkJs+DTwdJIeqMYKg6jDZnYA1CcPFGvku/zVuWTKHcu
+8XK1Rv6Ko+G9adHEG2N3ziHzXNPaqe33zj+I4pp4/Jw4DHn85pQAZZPpWxr0Ljp
wP+yFUKUz65Cm0PIEp6wh9yKbrcoK6jHMjP3MywvZ1DJ1tT/UjzYs6UE39hzrUyX
BGHDeANoLXnzMDwRsBaTeRwMfsZ9D5RlPGahGl6biqsnpLWbPUlE/8kqdHd4CrIw
KymQm7j3LkX7Qg8ZtAuNgpSa/IRqLq43r7Gi15psc10AIA6HtAokTc0e5oW4Xm4d
/RHVbA0cL4X26yBMQ6N4WFFUfgk0lan84nTepmEdmifSLmdilyyS02W/bhYh+/uQ
56IIsUr4bn0lmxqpir7DP/QAd/Eu5DAGgdZtpM6uFQS7wvCCg+QM030dbollqfIq
te/BAYb0mvsKBkZPlb4ppld7j+wMw6JyZmDJqndE0G8JAlQp/BLOegs/C1ocXEJE
jJndmvjy5KCQUInaf7ZWWie7riTju6h1uRsA7ZAdEZ9dFmROgBE0UDVfnyQ0Ppgt
OdFQ0gy2D4fIO8U7dKcoyJ9j1nA1B6YVHw6WpBZjTu4o+tWZ2r+QEqWOOTPr7D6U
TRtqquza8taycq9eEdRqm26QbKTuvfYS47sTx61ag1aaC2j2UQx2lzpjAL3eU++L
xJPs1iLfVGQIfYvYPbVCfffdKulZftKwJZ6fjtbPIWnurVWK8iYygPHFh613xv8Z
XynrEiCGPT62SOVIu+GW0YuPP08F4riw0MbFzDjbIsNe+R5CfCv4e17Ejb6DtWPr
tf835jiwPH6Qc6muIwbUY5jy4FRB/leRzKgbYpz9EW+B4sQ4KwrxwX+frcnYo1b1
4gCcquTW+UgGwco5enO1dRIT+8ZoWkLlC+fGfxn4RxC74sdzaPEB0mGiBj+UWFSZ
IHT8rJfU2CSyr7Yi/waqol5OffflmKjCbSCwjbwH6VtMAia0snYpsDh1TeFiDOMH
V97mWllrRb8GDHgAATCkiLZRaRZJIDEeuLWMVLFyXov6Ikso8SuPGpEQP3xtBAXw
hqwkmQN6S+Nqh/nWSBmwwVXcF+EmJEd8EAhacAPAV2H6ZdxfXxLewVgyiSKydC88
hbifmHtMZCoOl18EQpC4Njyt6g+U6UGZk95/QTjtQ4iWBzoewEcM6GgHqa5yFlo1
pMpzstxmsIrokJUVPXJGyIT7F50JXbUmycXt78IFbD8KrjPJLGMF9Yvq12QcunHj
UUnLDbV7+xlto3DtAmQLubrALrA7vUWrvxL3WRNmLUFirK9pvQ6N8oe88MEX2CbW
tvMQeo4FOpxecH71vBu2yc1KlokCLsZ8lLSxdnsd2sTdlIlvwopWzXMtivFyZ1r9
4OngD2AdD/6NBHmvF+klsFT/rSDqn5N7Mna4M9OEqPldxAodK6W1BIq2xqa1lyw0
iv2qLDw7JJn1QDf6ktSiiwwLUa+Ll1CqSmU5kkzqEauZgfdSn01AuGOX/hLUyMaA
ZRRIUVcPTN9/+GnVKmJQXTwcfN07mhi4flrSyZ7+uy4WwS071/oWkel2y6b0XRzy
vuK5ZFBzy/i2kgW79jVfvAeOWz3fvghpt9TnfkWQYwDQdaIf+zkAvE2S9ehGbs4y
l90S7F0+HE/nJD5mfGJf61XtneLXTYgL2pzDtFRjQMiLXL+JI7TkUjH5I1fVgpgT
SvJNBg9Qj9CWsOdpaDQt6iPqUhFENF1ttInsevZqHjDlrbjoes+GtTnkidOoiDMS
3h52px64o0j0r+2Zxp7+V9Vbjq+YDhnsbvvzQ6ZO1mgjmhWAQJDeT995KbrOgHZn
BKVPyX19N/+Rc1rGBJ/XLFjjbWsFLOyBINyHVlzJu/118u+Xl9WEjwD7AB2Sk5Ge
ECGklSzD+eSocdETMluIqHLA/xpUf4i8X64PpBPtP2cV5J8UGJjFoAsCZ/d/JHFS
Ojnv7Nk/7CvhkMjuVKma9m8d+WuCI5cVcrJL/YEpfZtsH0IoM5ZASmO6cY3O3ph5
5RYRRDenfk+NutkXDNBJUy5UGwoPxGQTroIBxRvWBVWJBFVzNzrQn/CJUcVHUBJ+
8svIPffoYeE+Z6LlFa8XKm57kq/FxKSZWmtmpJuO3mp0x3trTwwa6awg/kBsU7Eb
/i3VjY290E7oC1bfT4aqS/JyqIx31OHOpNUFV+5KLEeKiSFhAtV1Uv6lvyrUwZaU
lpWdTPTOSTYed8CLaRvUdu8NMFu6Ks0DiTMvppN5S9AkkWVpGArXIb3yOAoNE0ov
jSSaF+/ScBZC/88F62HRu4pdhql6cusZKLXS4HmRtEKamuKx0urfzqwNJzQ0RAoJ
2HXVmirlSsyKOuEl9UC+LLQ2ZDB3qAFF5DuviguNJRBmWY9H4YQ6KOyF0toKI6wF
p8ZG8+zjE/0riwY9ubMJrOJp7NBUM/dsMXhs2XgdCgeMfe6xeeaNRwC1bu9+85gJ
0Gy51N3vuSFeKIKX+IpwKXz7MnBNPTNaslGsqD8OslR6aW3yBa+uA5UqKkZwkfjo
1swIii9fiPzWxkSsGmSwbdas34BU3w59HGjeco5+0zDR35aDLQCCcT4ZxH/zLSGa
USug8Hi/LWfyCHDwBAcx6z9YKWrCkFox8rc5WVP6jygTnuUsS7fsgS7Ij1xQFjWH
zOCsNIcbKWbV7YKZpmD7FY2FOQLdpZwB4k97CBzU4zrGdYXclwFR1RP1F8PmEsQL
2nXp1XFk7WM7SCaWm4iCxrFKR4CVdxUQtOfe1zP4JEvNr4W87e7fDV2Zo4sdWuAt
tlGl8xnbCgm8n2xmHs6+a6XbWz3rtL3EM1zPLj5f0uwjU+ub/gK/i8aOI8v3X6EM
1ZRwV9yiV/hasrWhW+drNaB1E+UZCxJpy1lJ4KdmyKdS8oGfJvXXzEDTSPKj1k58
tp0DWvbaZXlCRl4USTaexnkaioLbRaA77mrfxb6GgTlqgEG6DHe84zVgd0rRHFJ7
LMyJjGSVLociflriAP3BFU2J7SHl7SvR1rrtZp7uOHiy22HwJ95HGfyygD/Cgv+h
1NLw9SIGdQA+bCEcHzxaJthzDreg+E0ejWIR2tSTt/yY0rg50C4Hpzm7bXMtdw92
Fnthh+ITpL3/QYtPf6pyyQYB5sHgilz+vBZu2uMXnTXRQAk54i7S+MPKN9buqDab
nyCbkjVOKtW7ZHOb2ylPweC0DyHfAK6/QqsIDYzdAtv/7VR265kzDSmzMwWQDzsO
Dwa8U/6NDqNRlGzQyrcmjesVWswzxflh/3TNo8XbApvoJNASdJdVkytVUaSErNJD
XK2PnT9QTo9FYU7wy39htQQpXOvGX5JGIRuiB2SmgGDDquTxBDDENqASg+WDu8OF
UuMC7eKrelUhyOSpG2PJusPTkmhe2Dpznv3hE/HNmrAijHgm0dT65UIUp6t/ec3Y
t81OYeJk/wc1NGIKlK8vPU2+DWmin39IZTtYFGflo48qOg7EL+K4+u9xImBk4UAJ
oJE04k/33MZh1Htvut/YTGBF5M58m9qpxeMq2sS7ZqtcgSlc9dt9u+3l+CYqQNXR
xu4bpPu1MS/yL6Dae+ES9JOp0MA3HP9KaSamuzmPr+0RQptgrj/Pt4bDy1t0PUy5
vaZcMfB67W398c77SUsUwoHXnofNEsi0wMca6DZux/pZh4JLtW4KOI0xqROTsnee
LpQb2SH6gDGfL2E3vwPnSIGERcp7wM+ysCyZqzaOT9+9lEqw19O8SHkcb19enB5A
e8HXKn7dC1sVNcGH/fdBocwILoEFYq0xUEx0JUJM7I4p8FcQb9vIZxLEl8RIEXKr
BV/t/N+fREy87OOo44u3snqs7tQ4qv+7ouHAfBRjEUCsIonVigu4JlUl+BbD/OvX
lpwqKRNU6yuomm8anRfCJY+p1Vf90sTaDOcS/MTffiZqWLiU+wBEgAcOqt9B7ty/
bfAARexs5oqXw0IlqySX1Fa4zOT28bLQTpN9nkJ5IVUgnIBVK5hILKGHYUrBnrWG
z3IkZsGCZDo8BIJ9x6b41j8/uhHgQTJkKc2YZBPV0NfdfkTCiqfiMZCg1mr4Piac
ca3zLzrt2cFnqPc7XKWyns46ZqCn09RNhJDtjUYaM+gjqOKGR+PjqhQ23Y6tGXK9
ZozzhDPWEd8tdpwP2bioLeKqRkZLBPCfGBAsg2yv2+pVqvHKQNHQoZhKLkt7uOw1
p/+1MKFrwwYkNanoSbfX0h1RKMgDaItYunQEEaX6kGNj6UbNngm0naF+4YAF2Uwm
rJrAGBmNgs3AiOj00rBqY0V5Wy0Z8QyxMjm8aqDoip+jvVNHFC32YjTh76q8RLFU
IV1WMbaX2hosXPM/FN291U8ZpL9AsEioX1dEDGBK81UBUNyHJtIB+VfIGfDTlfO8
coN+y6CPkoTW1NLTjA6bDxyeQ1kWLiyd+LeMhYSLZ+cjb4Bp8ufWlS5MhHRMZnhq
LLLbXztZX/3GpFrkgv/dL6NRz0pPFxnUYKL/lzbNF9hSCzkYkZ9V8R+tjJojKzhq
Th8tjIisSTY1aasgaSqg3edPJVX9b9FHRctwHXa0oov48eXxk8tCDC7IcGo3XhP/
qrDCQ6LDYolrE8et8BWgMmjUuZEga+3g8ImEwj4cFBVyjPnLPDp3sE9EukYa6Bhm
7o4T4IBoxtpiK4Uoa7wcH/KXjC92EkpTmdeUWiWhDRlFVG5waYHg29viuPrASN/m
MgC4i68qtemDTcoBWJFqBD5jNj667ncp0JBaiwiqSHuApn5NWDGJ4W/glvNxTK4r
qy6sBOFxzyV7e/252xDLLrKtC5ttpDu5ots6N0bRcsrwdY/A+YqBLbYNxnV8Reza
I7PzKtnZ54Xo+kDCUb3Opbzj3w8m3i+mcyUuV8OYDwSVImtvMA+hbki1ftU7JV+T
9WF66fxDtHRpSP4PrTepqVrvP9Nm40xQrXA4dH2/rmf/u6oMgoKyA75FkpAosyPL
bYiQLXsn4i/GH+Yv4MCSc3G4yntGmnYBj5oss79MInF9FXw/3BtslXjHFtFpRUaC
EOm9+4nFpIuxgoDBiE9uxaETmlnzwd5+suoC9twRSNxQEs4h0bmCQYbV8oR6keOo
/Fv13NzUCBafnjFBJxUjOMsru3f+ibQ+FlgUJ8xMFNNf8hMoq7N6lJWVAxC7HvFX
1LS9h9HFOi9fpeBQYaFNihb6JPuWpL75f9ZHc4IYY5qzQ7MAy0pfEn0C4eIgH0Wa
23zHQ2vx6f/61muf5yOI/SE82+4TrBusgRu4hk430Bdj87Fzu/7XEKRlqWM10TqV
s6pbUiNlpAIVh6d5Hqdl7V2Noim51/t+0nSykBB7g4M/+QJ2Kdd4zWOz4Cf2Dw29
PapQjAdgAP/bFcroXhB8MHuAmt8IOTYyraGlnWx1nW3kpYqYZZJqhnv8lpbteeaC
L4DWm01vmgmZ4xCS5WD+ySsbrTdN4VPCn77p4XdsoKGPTKHgtDx7cMaGd9572J4f
YUeIN13ickuPWOI/r2Wf1n/QlUj1ko9OG4YWM4bTJARphSqkR0m7qiAT2OZRnLan
q1YsyJ180TcxFqJZ/eIbXA0LKGrpIB+mSXI+5BLCwwT/vp87Mpu9Np8IYvQhhwHQ
LkF/Bi3dc6twDQf1EiuibDRK1/rG0BJkCS6H4FgigFpjN3elQHMXzdjzDiaG+zY6
jAH9Ce7BJ9Rv2P4YTs0LZIekeK32SzmFaMDLV8QKOwUAFYjZgG0+cCo/5BZTKEVh
LB1U8fFDCeZ3u4gim1V4fG3T1GdpBF4BqvP2yTfJ08zAk5PRRgcvU3OIYmxF/VLs
tzRCpuMmz4UTEtym8HS4bER2Qn/sc8WJHKsyagDsQMM+piBimqdiAAgCkcMWnC2N
w0ozarWezdbb5SXadpG4Ep3N2IGRx9Tcph62ln8wC9tICt55p7ZsSmJ2lvI470j9
E6AuQK2N69RmBrs2uTCpTgdoZpP2Ut5owDgyQRKllx+btptExXlA1ASA2l4w965x
IASO4VLTf6Wb7gwyuW1jTc6I1dP+C3jaPlQISypEyQkb+BmstrR01p4X222gRn5W
FFM3UuNhmP7OJvpcsjs+o90ItOLeLjpIqh6SV6IDp6BAjQ0t26DjTr7M/5AtkPK4
SZn9ZGn1OBR2LwPZ4U9nfmAARZE/Rh6XuppUN9PVa9R8jJb+urCOXcoLgxnEakuP
sisnZxaF1FleHYCh8UGWxaMexwEalPZuG7/BYpBuMy1gysRCa93/sKwFQ7jA5l+w
k0ifZfx6hRHcsG1yFPhd25SJ9KhaSCIaGvYtq0RYzl9yAwIKijX5RXJEN3SyeGIM
rjW/vNATFcsAO+ZAe1igHWz+FzPwfzkdoyERqudb9xSOsQdYjCmMJZzdvvk+a2sI
h+u1Y7e2wBN+RhlhhEEOZu4+NZSkBOiSzrvyPR/pgmJ/grjs0f6M3X8R4HgKGT+C
9qYt/6S9DBuz+tHbwXJrNdWeNJ9/oRf2GiGNH6kEJ4DbRQuuU+2KhAQVkZL6LYGi
oHsTab+wKVeMSRu5yrUBh3jNqCbCFWaGfSFhweO6PFlebKfaHkbvY9SI1RygOe2Y
NGjUnSPAG6z/kZEUOKc/9VdRVpWSBCWbO0v7sIR3dEfFDte4OXIJLj4eaoxIw+QH
kPYwt9vj0GH0NSV6wRP3rmO+IPty8yesIL6Oz2+TBylt4fHV/jV87qk8O5xFq3P/
HL1riM2BnxH1Daf/YvFRtm+5SWnh6FAjWSVwU868yLRatyCjuiwYQACraQATYGEB
KU2+axHFo0dgaRvq7qyp4r6kBWsp1EwdZX7WgXIjKzq/RdPz8vAwT6MTeaH3rIaE
B2ByrfZ9zsuno4cDmz2FyolNgwRLQKY5Hm36CBeDdQ0nJIvz76hSqo6QFVYoHuEU
Qb540sUu2yZzkdO/XXwXTI0NPDE8BBOSlPL7QsH+kKWaLn10ZJY9m5wYScA+gSnB
yHpvLJVlGEPZM2jGkTHipvLvaZiw7FWRqYivFuoqZw5Pu6HB2CAvpBt8N8i8eXV2
6r1LNs+LwkKra3oR7fPTUjbu9zwy7bFLRDPPBgKwMo2FLdzH4CBOfKbp2Jxm/YqM
kI/XgOm18f6YNJMGBTaby82IlvUm0OH8DC8EmepePnoSa03mjCo79LiS0JMwJ8oc
+IIaGk0UHxlf5idBHW33KqPDW4O+bH8LZ9hRu6oxwu91+/tOKoZWmiyHMbmvgPMm
N93aJK8FAp1PttOQAYEAByUnK6vwhtM/gB4Px2bIkbsNmGcIgjXNjPWT6BOgiCdO
tCHL03sQnnWABFGstH4XrHUi/UbfupMaHkYKRRdodqu9URmik62wfQN/3Urs05JI
Xu+mz7SBTQRpp8N2JFMsaI5Z7ioYnsTJp8qOw6Z+QVQ8jIvmY/SNOKAwuqPK5GE0
UMd0ouvVKj4OPrr9XwaA0Jk2Fb5xqLImwzt+X2SSsdbntvboMRqjKgEtAnBjV/mF
+qE+zmJiRLeJZxJahYjGleCACZo1Njt7anP27OpFnGEzmBi90U8dkbsgFB0J2Taz
2qC2uS/Cfh2woDjVrHW192Yv7TtpiqFxflPBGGUFYUxCLxxrk9EbWCACTi65QzBv
hcsHwU92E31FybCBtQFOUc/du8cNVtDmOk7H/t+A+p0WGsw7C8G+Fs01+2lDz2UE
v0cwnrvFo+hn3jyDB1tUhNf/4hW6x4o7nQdbPOf9aeUikCnpEp7t66sxp3XCGIeU
2M5dzaIBOJWi/BlSF5lX0UHWMPIWY59PHSey2JMkHG+iHu2OPF9q8cRb1ViY03NY
OCzjt6MxQ0QHgEeOTauAmawMLtzDNDgYUfY+yCAsCXtUcCHlLx57pJ/kdZmKRzVh
KWm7F9MVSa7OPl6+K292zDQNfIjuK5+4vmrdn+kLIwca9F4vb5KdSBQmwtdAdSIx
Lc8fNkoMawCpNe+Ip46LxMggV9fr4K9RO+aZ5k6QNRS2RQW8MwsJg7UuCFs+csMA
05e4GD9byFjv5NNx3/MP/yE9sPIAq5+7G2HcSjYuNUvYw1CmXzAEhV3hP0BtCYgr
ajslcQS4gLTMGi/AGXd9wnCsXwz257OuaTry2QcK+MEwDsITk9xg71bLng5qaKJS
9dBLShBkTsnP3GN99NMvKZ/6L7E/vY19z5f1kd0VLaKtxzZ2QeKCospTCnY+UctU
atEqigwuBnGIpitCXJSbIrMifkmSFhHSEaAubSizYeb4qH2JDoIvtqIODLioTKqw
KLZmhoI++ue0re+liTA9/L2xOcS235otkV0041dueUMhXoe5Pscz5OlVR6PglQUZ
86CUvNOG3Aw+gWaor9BDYeC0AbkjyHdIR4fb9cv/UpRQEFI5h6SWbXrbqXN/nGdh
fzgMYCSBGsEDraDtMlXpZfAdbea7aDfCEfzWTAyYqBxS/CLRAnbdzhNkgfgkf8Jp
X9hDnu+NM9oZ1sPZF1GuZIRd2OyvBfTzdqLSld8IfHSRTaqIv2+Gr6hrcmKTIUjX
BOlSJ4vK8P2EkL1Ot9r4BNh/13N1/9kzIb5agdOrH6BzEYLnRHE6rdSUuySoHY5Z
AjU5E3fhukgOBiTG5UG+wVFbob3tSzhWGh6Vm2zchjp7P01RqSc4aTJVwBwVnckR
YEujCiJFMw4HJ8D7GbGHOHNhuyPKyMC7wemz3l2M+q7v/r2xVXDkALhjxHV/JV1Y
d7JMMj58d+vckHA7MvGSt9ia3SZnXhYM8/clQBuNjvoMwNK8I4PVVQjypFcwtsl3
sxcTji+31GGZtVKDT9TmjKkFJ6re+OVLVqb49O0+UXknCbvDr9CEZQASkwklshCW
mldCjXdzjwXJsd9IlmpbhysDiD2SP+R6wVq7tHDWdzdui2MHXXvtQe+yNuHCg9vI
b7kkRHSVDUDh+Z80wpBjvBDqY7kVCHtJmMV1OVCweAmlllvt8mP1e0UROuAJQC93
UOSSegqG3nxYjoBjxFYVw3v6dOBg8WkgVsSU2qNXQBOthQOyoksWN+xlIsFHMFQK
8QssN7AuRnKMV41WZZLILfEhFmzcpzyzggtBCKg9uokwmOsuS1H4VyfYR6Jc7xt6
USftysqCGrG1bxnATeDfHgdm5dA+y+k9UD15k5qE9oL0Y77ZrZcAZMRTAj0PAiUJ
Rkc1u9qpfBTaJYkoHgJCFb9kdqYFE0ae5hPNZvZSuu9LqOddlM1XXBRps2p17tLi
Kvnz8NHwKt6wtAW5KhSgCblk6nkQWO+Eyisj1xPcL1Cad9paRp8WGFZ/jmhfTFKK
Yh9OsMLUGFkO1cLW+8vXxhvxMtGTwHC9Evzow4nun4FdMGidCny1GbSjk7IaE+OO
03BA7pekUsWix34ZJlYHVEHmceOWYwTHSZzQb2SPUPtWcXJegtyuVOFx99TkbPiA
/eu6oipNQ+cv5ZKa9f3DboZaQ766C6KT+WK10ppSXmWKdADeosouboj18cmZAE3D
ZGLlZiwXjKT3mJknMqpbA/84TRLoPlIneohXuonuFfniofb7C9y5npBnVn0chlrD
2gIIV54vDKCgrBs9q35k31K1ajtb4wnVBFzCxeBlpKkehhr8K/Z4fGnFWBtpDUQv
KMrszQ07ovkBNhoOXwK18mw2d3vHq3hVEpQB9yowKMQ74Z6THc6TIDCSGueKj9UP
+cnqsxuYyQXiBW0nYYhvjyDfb4ZE4VL3E/LYjnpFGmP/frbNx2d0/GllskJtw1s2
g3ko+lcLCTKC/JBGH2dN+/Mq+4AVqUK304LznOxsBWUwDJ6K89gTKHOEzjMvoNQo
huwPfGUHwif/ouyHs5KHc092ZLvwZvpCE+EtppfWMXu5S7AEVq7vNWlb2Nbywdg6
qie/Dh/oPSWMIXQUsxHwskC9zmdzwLNwzA8yAXbj6P2je1Xp6fvyksEKumki2eoo
BjYraFKXfi8zy3coYSJC39vDT8+Y5428CbFO5kKzU9R2l69M1liR7avvqBBYewlZ
41J/sXWqitcqK/9m4CCecT+2X6HO045HPx3LQ55h9zfG7dbytIlSKWxqGgp0B1o5
/rO6u1uxmiyiO3pJskZY+mKOmbsZ2TQZC7fnCXtSDgby0gSSZSz950U+SoTqCldY
dWD0N+kNqMuyDaDjNJyOGcdC8jniAeM/5jzNTGbcA1mIj4+0X3e8JLKzY0k26GAD
In3AxvmQztrCyAl5lePe7gBwG5mGPtM5htbI806US9pNGvvzMBeTEIkp3Yzc6xbV
HpakkjFXl3W/hpGOaqASYk8QuzYTtdMwy6YIvBCVDorM5E+B3P+Lt57v9VX0Vpmf
CcnSZkt/92khTVeQMQHB8EOFHBB0ZWmmUDiVdrHg7bhvmAQwYDjypTJklokYmedg
clKh4Jqp7fkIXFVFd9CLXdQXhN/AX8LzN0BWsbz9OSN4OgNf8sQcRmr4SBOGUZOw
ecsPxY1B+BgiCD935tvipcI/RPkAicv2/n5mI4n2cqkkLNmmxup+oeHujuj81X6P
NiT73ZN3Hyj9Q/mPj+DLAVwfpVW1Jsl6BVasTr+6d0UTIpLfhue6Jl2jWdZq1W2y
SAHFrecdoJCzJfsf7tTwkGYseUOh59hiYlh8CsuJMYBo+0/L5swtBdWaQPfBWCzp
SCdk5bmVE87HhfF1YREZew80HZ5C24p1p2xbB1wU2/b2bhRFIZhhg0cUUOgcebmw
aCKi/EMtqxos23d0+i1EAf3gMUJrYQ0oVBTFC+hiQxyqbJnalBsPfP6fvXm5RSk+
l3FPNP16Q5CHwjLvFnKLhz/K6x9LVRURzrDQarN0dHjCXWK14hMUD5JKWPw2KPe5
zB/GwluMwXY7lOKuK4aDl31t23I+7c6Ou61IXNQpbn1oHEsbAEyqMFNo3kk9nBnh
2soEUtesjQgSG7njiMUzwnIYdDAzvbuJjmIAM/5/iX2Kptn7sFal9Wev3QLfVvYu
H05FkoDEXBsKpjTKhEhNNMy3RnvySLAd/Hnl3VH5qxToGKoTf2eXBNRAMVy5U6Xz
aUVLZvdEzjr5OTMa/3jrtxZ/VPvoUGL/Av0eQOcBwMMruDRotSSJ7vpyI0sl1Aqh
q8MW15VS/c9Rp+xPsaYBQubF5X+zal+AidrJ2Yir1GnTD1qCYy5VubSJ/EjjRkjt
JTNHhegbwG/sf3xERskUg5bZobksUx1op9o9T4i9Y3i582BUv/4/DlQDHWiDfOUV
G4NHEPXKNtxEAzgHOG+M1dzDP7211B8j0JDqB/GMkzsFAuAREW9EQltKqjDDtRFR
ljNFx+FrfmAliz3/NXzPNiWPfNhP+78R4VJJ0NYH8RJJ9qXmlJUOSKkJafQ+uHpd
G1+I+Yn3t661mlCreNAh403ME51NNeilH5zryJY6H7XzeiwlxSRtmD40wKe6VuR0
91LJROb7TpuwjprWJHM60p6nGYTTxK126SHseQd/Zunxb2w7p4q85i1z2q5rO+uQ
3pemmPUJVJ6/In0y+BqVSwmoGrl+OsKIh3JIAxDkXWB3QKdIT2XZChLqs9rRdZaf
O3784k5mapl0BHLcCtk3pNliJI4+dEJw7rmfJGoUcbbrcPRT+zRnkUdHqRC2JNAp
VJxxoiGm360Iy+jTa258NZSbAe2iS34v6PQ15L8A3rZgyTo49U7YKHBhNKGoDJsV
rQlokinGt4NtCh0ceCrJXTScr0V7NG5q61jPq3+RZbY9MgVu67edlGX75M42WAul
uda7wda2Rdwf6Y+hqpjDvZvDFtFUFSpl3nw1ZiB8S7MeD/IJYhBxjbtx23gcrlmv
L0oom9UL+uvjpKS31tampoP9Bq8/uASY5WGaYg0kLFJoaPT+VPVXNzecJ7kBQfNl
ngfbBNmoX1n5rSevd637AbTacOmjmnM87tCQg2H7682RiiPaCrn03PqWAJiCg7Xi
jvQDi6Zs0bwGHGB3dmxvP8PJzBb+V235aIqcQafg4qyQg3yQ9xzNg+tI+KT+9HA0
rNjzDEN1JSfAWdoEUydHe1BtkS5Bff4b6SN6/uw5M6mgqbYW2dUpudzu8Mu80X94
9HYYmADY8uStBxgq39U1xw+nmNjCEcg+4AYxctRBFRff/OaHRaLkhh95v0zUgR9s
COcMJwEY7SqV+SGQnqaQ3FNjT37Q+Tgfr/kF1l2ZsGFRs+i3KYik5fIi4zHuuKgK
8eMqyOwitlXYb8bjRGR2FF09pb0uS7kA8PaVPCggqz56knwk3OADGLXZhBDw/d4H
e/mIjfevt8jNq8MF/z2jA0ACvR1/wKvFL2+2BY0E0BeDg62AncXEa0voBSyGNq3k
rD9FX2il6Osd6+mLKQTrLIqvoPRkVbAtj2uY/vNlUanb3JFS3S0+oGgKzmhmMxqZ
njQR5/sSRYh9h9IobMVEX8O0p+S4HW40+nRONRT83VBwjy2osg9mkpGZkTDj5Xaw
n0CDhTwYeL07x/CCVpcLadZYgYq0O1Oh+n4LhLOBAfibc4cMyXK0HhpYSYKsAAQM
f82Xuoc5/qqLYHg5ZCxKxTitydiWX4fmy2zRr8YDI4af6cA3JLt7yvUduDKDtG+F
4/ZIpRcN4Muhj/Ad566U1/Kli95TR9DGE2xCjvQuFrN1Spcu6rJeweA+lD8cPX1R
5XxjOtJUHlCmCEGMLZaH8/OrGWh0B2n6XwopcSLN1yNSkkYJH6HOu3d1RWvrimU7
WMh2/RdxupB5OkSPmTlkdz8DgzvSx7i1i/PJ92fWNAiEp+mJSkD2b7M0ZtQTrJdl
t4mz/995a6H94S69KzxYosgs181ESP2KDNZ8A6po999xxFlWpDOvG1ry4FABP5WF
I3BWLWO8caXjsDXXKWLeIgjQ6eUMVJ5ljEqXgk3LlJWjsVXulLKRJkLYca7CUA7z
Jkms9cABl4gfhPuhk8MncTyCETFLiqjRhkWNVt+0Negp4nEOzLQSpK+W0eS3rQiG
4PDNt4mOHHUHH7fWcAPchKdxwb3E3KK2mQr5RPcXGQ3sXLKw/iuLik3zBpQfuHjv
jmraoC7146jWP2U24j0pUk4v3t+r0kNX9YzrbyW/R1bqoqtoGTyr6/ZJN/fpdxs1
c4bLkkK+FaV1YMN0a7cgaLAaF0mQVPZ5/Qc/V402igEM+5hBg5QZNmt8qt6TEylq
pYBFQKbQCv4wp/VvyYwfVynY8lpArlwpvQgN0SJ9kmJUkS80V0ojMf77W8oLXo5p
enY2bBFT8YvJ0WiWsYJQGOiB8AOwjagUdKv7PEnY2GvHA2bnJkkHSy7MuTdXQJhQ
lhlg1lhQnmQIGraJqr3j3sFvVGlVtXzWK0Zeu6XYRNJmGi+AsLme50IuTuFh77E2
0Xe6OSsXeLTKqQqWcQwBISPEjwe8NcmvhgUOpYi+NDgxUaeGbj8ofGl32u8z5DsP
xweN+N9sE1xNNjDt24HkRLuH2SVCy4CjfV5jwP/MbOG/5JXdElfR9t1tPF1WRsgO
NIMcDuo8BqQpltSJ3FkCtjZq8q5pLADDHnvgv0AmE/IzVPKr9EhKCi90NHu+18kO
0gqa2lcp+Kx13lD8WUEfDKS7DwLyImMWEbCTvojlIvBSCu2I3wdmgT9Na4o6Yjq0
I48CDFM5Eia54Zx86IFGIktG4FaHhiB7pwGJv3YbVLVidMTboGjo3IsCcqFCKnNs
JUH9kYRzNiAK0Zg0IibSXBp/5JJp1VkojnSjfWbv+L0g0q+hnhP0nBR3puj9Drha
fDu/oMHEAJ/JstHKmVPO73c1wL8dq8ZN13yJHjAVoKtcKhTmVTnEYbugKsT9bbdv
UTnhro01ohcBh0LQHHc5yDLksSecHi6xizKg6XWzn6WT7/JHg2vEjPz6PKYpRzV/
JeX29UWCrTrnvJ8ZUXzJ97ri6MAiNNkI2lhY6M8AqT3WP5kW5msJ+YXJ8t5k7tx+
m4tHuF3NkttZKXRxVEg6UBEbNeAJsl8HuhdmLI3WGojbPapcSYLLRiSbha7AtUnV
6amxwwy6hifn4sf30wfyUjZNMQqYBF8vRgLq2CBED4hLdwL9dC4z3WRwO4qTnYDj
t2B6POy3iGRKYRsHFjS9xVPIrf1NyC3hIvhxD+GQWRzN93AtTMp/dCQ5TYA4KTKl
4APpphWrMRRkyKnbIo0ORDyUrpuA81x1RspV+qwE83YBC62sy/aLBLydxtm4cx1B
b8yhl1qgn1BZm7hgK61bvmaaRMEB38IJZCgWRHipjfFnliBzrQYX/ZgOdYYO0pDE
BAnenoqLoW3QQztSlAQMzpTYLNRncP93rRiIf986R4wke1EqGZtLtUxdeXrrkGvT
V/CboH0y1Kj1/q1PVCMsra214jN5DSWM6gJ9jTej0S6FaZstrIJ3POyMEUtP0rwj
bt9zti4+WOhTlw2h7SF8HOuABApurDZwWviR+cGTw3RURyIUWqTMTNEVOUqH2zkk
1wd5PHGk9CqyPV5A8qyjn+KuJmsGRFDekOKXq/YURamCLRnRp/mjtkeZV0PnFM9o
hTd18SS1V4DnDYJ5LaMrf1j5907aAY+jTs7FsDLEwjo1f/UOteGyS7/tTYnzYOUe
7aDZlitWsGLZyu7DR/So2ckr+PxWt1DAD4QbjfKAgLJypqAxZjQh6rAlLScUMZPE
YaU3jJ2WW+1j6q+E9v7SQ5vef5NIvseCJZEs/zNX9M5DDzaXe8nm+IxnwK2IWgIy
mSz8/FmnEnWd7JzfUEscB149AD98YMvSxfltFwku/lLLd3wqKx5Y6UXrwLEgwBgu
BISrenLeMQ7f7iOy718/lFsl4bOKPhQfV8ETGAntOAufqcLS3mtUV3L9V+QXyHsn
ih9dlzAMNguwApyNCBxJGnz/Vk8skGHciwnBtGuZezsDLOVc9jDnrHagJd9mwUl+
uvTo/FyUTghX8GpKC57A+tsqwyD+fQVQtmaxKvjIQTwyflk7B1jNG40z05NX2ASK
6neDFOCUVbg8ZAVccIQle2eXee3nDYyfUzr1KnUSFSO2xCdyzDBK5BSjtckuQ53w
RZHcdNU1IA741sP7Qn5jBAjPn8wGjQCW2I1SPqA4M1mOe0vmwP4j2gCxRNzgjM2G
C+x558Cr2TBsNTcRMBUtcWnJ3cXADLtBPHvVN4XRZul9Tg7aH6LOXuPO2exTWS4i
ksCNOp//HLq7FFEB8LMYd1D1t1awGwvi3T89AdKA4DMmsr1KNlOE4AwGDhnXUEr9
uft7E40FNKVRkGeAwXic8tIwxXtMKJaz48BZauJFvUC1cieoqPyRYxePGPypT3s0
2qrrEb2B9FPLzvBCUZ1/UfqP0T0/N2JTc6cJaS5HO8hzlS+FuDhauqVPUn43WuSM
IpyVefCdlBm4UV6A9AH94B0jqg0GYut64hW/g3ARQ6G3tDuTDgPkw6BJwFBtS5F+
upGymsL5sRQrjK00EyfrCwrPhHvb5goYoAe5ezN/obNGUW/LEmu468/Lkmk0MNSc
pDw/3leLe375NNc6foz0AxmcRgbLaQiW9aCX9pBGExdfckEfew41MDRz7xYYEEUK
Jxukod6SCUSfX4usnAVFphHmDrw3MyvD3DoRICEcZPf6vV5H4wVyclcDcNI+cohk
EQr0EJPVYptZDrPRpU0x5TFu0v59LF2dQpjL5QbfTQ40Fyb2T7FrBv5M0K4XUpwU
c1vJUNgRheUQYEq+VZ7mGAGt7TEzeoevBsQuG4NBtpPEplgNpbd/+9d6GHtvDGx0
CnUSWZ7geDTsXWpnx2gcJPNDse4Bf6qcIINStp1FS8cAuqiXidCuwiXM6FrsD/wQ
h+zb3KGYdT+KCN8XPEiQe+BwneqyzQH+oJg9sY9T3uIW8Jq4wuR42W5Ah2AeKL04
gB9jPLZRX7gHukj18V/li2t0qkcB7KLiAgBf77jkRAaZXilvjwC0EgNEaq6xkE7o
6VurC1SsZEeJNgNUWCcj1JAd9odntKiz6167cRlxf3V+Sd8ADjXnej+HQ5c6PlZQ
UQcURTUTLVpF/2sDOAaAOVX5jXHU6BQIG66SxvOYMJfzNT04ZDPPfNJT1GgyLRtd
uC9N2+cl9xjb1kAUMSKy8VlosrB3xYnVKEUxTPXlwr4+IdeF1nCTlUVYLh+zzezC
Yq5YUiUtVbyfQm+KUSUYIqUA+VZrcMcRyWuUGtl3ggKFxtbacfQOjcuBoJ8Vkhs0
tyPvlA1v8QrqsFr6xfCKS79EHY2gufR3j8W4ZRdEfddMBqcZQ29uAhtIjRIlKgwm
HH4K8TuOyfKppE0uo9/7+jIzBz1tFt1Sn5BtpaXCs5O2Sbk0U6mf7b67bdTpoQX7
zMhtPK5KiPKWOn+cSq9S+BiUA8h1dFy2B/Da44FTRXAtogDpIxeyti2DievUWJ0x
UxLe1o/BshYlA+gkelY9XLijcCzchVkr/UhSsel19dA6V/+a2Nyefb61OPI/VmBn
MvBJrP7NSThxBiVgs3+Ertjtw4nQ87rL8s0O4+eGnswOSqclSdoh0iiGrCFVccKd
5AVoWfQLUmlY8yrQcOESQYAMSutCOHFKQpJ5LIRpPOjzu11KiucO8EX2BPS9EGP/
hnNfbnbDG9CeoOnAD2lyczI1MYXGSTx3aRTCM/dR75DNRlhbnqpolkKGVgyZp8cc
evCtXH+89PY46Q4Mpb6+woPO6QREoaSqA4pRXtjkH+2/M6CaTvnrva8fxS+hOdJy
fy0btMHf2sniBMODZMBNczu2HfOFWL+uEN5S995uK2SHzdGp7YgjC6+V+UidxYwT
3aOZ/z5uizI4n6qLrsubBJgN/O2jAF9bjcyIz3xXUAXavGy2kpPBGuMUQbTS8z9R
LabO7MGUMhkGEKM1uXvzpWXOQ4t2v75kDxeQBLjsN2E+z/bu8ip7OAl3VOtD3QBS
SNBOG8md378ed+yey2jeI6ZvMEcBbjtbhBjnRoId0XNUeHoBl2gseKXHwNuWFaxm
682+B4TKHHyxioNzQToLBJ24bXe4IQDox2d+ddvOTO+PTJu6scAPqEZyufCr+7Ml
gzrgsmBmI4OXydICXT/OKHDU3BwhqvsE8pieps0jCyDD7QkdqOdKP9bDna0FyDrw
kRrgHdGK9Eyq5W4ZWKUGBi/mFxfwINXo/d6GmQ10Rt9TFResK95CoBmkeQNZhqwc
SxtJZoPdggL10PrTq4Q4H59Oq7BtbusbhKPH6iV/tzE9dXC+f/9DJkqRyGF8uolF
nOTFW+ZrIgSw1atndzpH7MLUAK2OGbUPXRoetxcyujFgwgT2q8bRZgnZgOX5LsC6
X8l2QrEjIq6r9U4qFWFKDzTjollWg5wFik5qCo4xXY6GnNUtrabjRoN+JGvlEq5y
W0gnbkjTBK4fV5TtvbbQ1rSo+u3DrxVfbwc13hS+KYvvFCAAn59ODKm0n9gms2DN
us9nBkrBArEs1X5I5Luvj0MTHN3kRhZvBHsDXhjjTCi6gySaXrp0p1iGpulQmdZz
GuriZcZHDddEEyUW/TpShb9DlcP01ZKJ7WUogsQlPFT91mQbV1Hjbw7YMUI7g4WY
DgjJx8kCP35d7I+vg+Emsn/ZYjv7HTl8ZSRaBUrdM8DiL1EfR3jjvTXOlFmxCHwP
QSuRDs/GdBoAvEFm1MKV9hu9uTReOqhb+E69etnfhJYHOcl6WNwur9EJxuc9/MxB
it72IxBfDRIcpY8ZDR0l+CwRzgSlvB3yV0S3JHoHcOAY1ObR1A77EeRtxjbb4MS2
msBm/hI0jTkBl/tOcC7VY2tdzYWjhoc9CwY9s2LunsRZHpXZgIpraO8uDV0GevT8
XBEl4RE/vVR1VZIhopidjJvHfhQg+jxGeKUbZLrsQdIEKg/zfJu9ZhaG/3XIZmN7
SxoXeiM2NqrQ0w4tkAxcI6fA3oJcDMTv0EtEKoQErDJbS9K5Tf0pVWZRfE9DxUqu
RQHmhsTngjE9Kx/ehGkYn3yfnTfAc1RQr5Dyz79GRX6sX2N8DrQQyc39QqaS7Gyr
Y5gKSUtjk414kgwvNTsAf/PGBDe5r6HF6JSOEV5GhZuqV5Y1oJwMORQi5nhvz4kj
Czi1+lr2hL4GNDmtZDziWJ4JJr371JOz7uA1ArA8Yhrl/Q1iclXuI4ukVmfYpJ6Z
Mw6BCBKg/py63V6SVzIx3Hf96VSUp14lndUjQhz310ENtiPPhsik+bF/uNxWi+oh
i0fRp/sI89H2Prgni8cJChovH+LiBw2mxxgG1iUlBRCc9zfUULxKT9GGtFXO17wg
BUsHgVVRwapeM7yC6JlCoy48iJlx1PQho+h5RBn5dgOErbVOG2I5k2+C6e3ASDys
EHQSAEAi6RabadV7sMS1sZBIwrn9nt8kBtKFu0CYnHYtJAWHcNuwT71U8nzH7Op5
A11QtH2PblcuVszxnxQEHA==
`protect END_PROTECTED
