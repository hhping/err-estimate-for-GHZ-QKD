`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiVWzFHMfYASiMy//MoZS0zO1xGDxK8BXSOCl7MIJZAd9oTevQbrku1Fi5UsREFX
/fuj6+yjqNNT+0PX/tmwchruosS7hEaRCWnAediM/dvb3TIxOuLz3PQl897WV6Fz
Ju2kAk0URixjIRoMlNTwygvpIcoYa6Ip7dxoyvoYUG/QPK9W7xtTDBaNdl+uhP4w
C2oGneVgg1GzFZGesyUh2MGS0dUS+o9jD27A8KsRdaZuPbAekC9fMpddeb0E/iVq
Ia7gPcfgJMOhh/jGWB2/QZwPQroYsqktsOO4UK+WCzXCNvy+G1MRp5UKxbfpbInG
cD39quVqK5MMJ1HIsMp3apvnqXKZCpfxmK03PCz9K5tSg3+2L88ylswPukBqMN21
bUQdMhD2jLP1DEXKldSoGg==
`protect END_PROTECTED
