`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
45TU7azk0mKm6ZOVjU5YgiI8vCtox2uahiw2ivV/Coal7m0ta5HJ5gaMPnNhnyxA
MP8S4suymdXt9Q4rUd7isDPuIUywkVWtZiJ9zv5xY8uO0j959WyIuW8VNapKlyXm
tljmITt0aInOTlOm5/Y1q0oegoEsueXIz/jD1TEsfykkyfSUztAcOKZNQaDT5X9+
myCuVjWFVcXFfK6av+7dMKdvy/e6mOF09lWaxL0bsYtZHiu8bIImSjDGw/8QFLjh
GgAgJkqRJN37wuPvhDK7G/PSphHo14x+GZaS+x/IpYHCfno4egcadk7f9etZ/ypS
zMYy85QTU+dV3ZIxUwdStbt7NIQkn5NEWUtjISLkf8TafD5lppf/TbQl8DzkBcb+
dH2uV69DNBhOtPpegfPWPJrd2QY8SqoilwGl609iyeG7lLMQym5O/Gg5hy5u0OyL
4hy7M4aSPoaSanGIQbSXW2bHGoNxDT2hRYdMYzqUMc0ziz96wkoFhXVEyY2ZJ5qi
NnXQJ0z9Rf0yg4XWxMIpHQXFNV1AbGmoqe3wuZ3WOSHIVbGYlP7dWSAVKN2P3NHs
XJR5YDmrFd/RmbgE1HmyEK2kXN2g3nJWX1Bpkn6zT+OvA0CUZx20VMj14TkIbJbD
WKtfxJoyBcO2g3pdjN8As5Kdcy1iTzy5iElAhSZQB7JA32DDXTkv0TAeKCLu9yx5
gp8lZNqmZXc0dufhxaydDpYb6fVYjIgznkP06+xSkwjGfEDpZQ8cYnbilWYEKC1V
MCFCH93fFPcJZxJ/dIo8zCUCly1gzaU+Jko5E+/ZJ6MVTc6yAWMnl3mC1u3WfwgJ
Vx4noyDReYKIvKize9o/KjoAn22GRua132IhfpJ6UccM2ojmUp/Cusce+HX2mhH1
4tfffRIIzOEPtJuONQKDecdAUqZmhu68e2sPlBfKHx9QAtRJLHX+aYvJpsl4iQAY
g4dnA1DOD4E7jjUCbbLI6myLlKzJDvp25nFgXjtQwB7CgTuQz+LOtE5qNKaCDLOn
lWE2rh1BlWkTDcuwt4U+n2AU0hbS5fu+ccALU3J3cn9b2UCKcIzmB4dwRC44nxCY
Uadagjph4GAOJPsb3giLpKm92f2OMKjHmv7x3IOUhJxCA9UWzjlTnRsqQc3Vh5Q2
vH+4QsCz8R+vL9Ig1P6X4tbpjpyxnxvUpEQlVaiTE83oqpHmIoROldJnJq2fdvmw
R23WIixD+wvtWSBOydveFfpBDv5njyqsy8XpN4auVxD0gT5XfuehNgo7/7DcIsqO
Mb+IUpY5r4kgHWpYe0YYniCJflgp6MFzGmK5jPfaMRgyVv6MXJfiHum8P5llQo+8
QeaRX6ttLUPJBxe8UKfirvb8w3ZLP/ba/g9Tdu2jKA5rlGdrzzS1NIi0XippTuqg
6tJZsijeivdB2ncY0gAlv08frmg4YpPpBEpd+pWWclwWtASZzc5uBAOclw5xi2Bi
MSX3lQFU6OgjdMfSyBOjADqnfDaSVEIIpERC9QzgERooZaPqOaZ6nxgpet9LoM7f
5NxLoM0j3B7Yhr8BbdKB+KvqPvKSDAN1yBj5pLWtHyI1M6R90jnzfTTS6UVy+eWu
C6a1dwWqFW3pyffifdJ1i7Iv2sjMTgNTweo5+7iUlyf6MT3f8dQDRXakoHUJll41
7gmXIjG6IhBVFfUcFvIU+kZK5XWtvMSs42MhJnPSDhaeivIL6CsxP70zNCCmAcB0
2tj5fu6oy8K56eWQjDrCNfcGgT2F2qJ4usIIMQhwC4W1ygMbzOdiJgcgz2wCTv/X
zfLvzFePo/CkyYIsbApr+7F7tOub+Cs3XC3LafEkn06AI2klru3DaFCIM5PZQTF3
DJxkVE6rSu2aGxrreXPwhTP3H8lWBWgR2L+CmHfMGCeEZhUoBxbFCJbbPlV2Wc9i
op9c7q0nHxg5/nSqrQMoubNSOlYwWuUDFHJ3WjTVD48532b6ADnTAejRp743xybI
LadL9/ISybdG1RTnTFbI97gc7VfrcNoPmOr/8UgVYdHXSbUPS5ghAJqcnc5xJlmu
XkVNkwonHAAGeLVyBTfPhuuuNjSMZB5Bhm+FCB/UHHu/pF18e1DXP5lsLrbBwsXm
1Tai9G/x2yz6oLhzBNyGZP1abVs1MmNSjf4GJWZD+mxZb+lyhjLEPM8VZC1SDZog
1RJqCkSNdbhzL0CoDl4IOE0eJ9WFozcyqSIjH2ZoOpJVMnAes2ZMrIVd2uOtm3v3
ENlwOmAo1w5jbMt4WDNVt7z+Uo5jQq+Lla8n11CR55cET8sHxOm1MJ/gO0MYn0GJ
Kje8/C5OLLjFUlyHCw1ZeQ==
`protect END_PROTECTED
