`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ouB3yGwIB8WeNINkdVn4WUiUKzRNB5L1DVSpbmWecoPU7kk4xAT7mfWmCit90z21
lZwirHDOAdKzy2ViaH2rDzmPYlPEHFSRP8NWPZeIZzrmjgjtM6wLN2Zck0G4/ALj
d2KgWba01lsq01vt0oW4zYM15RrpF4ivVwi0auabvGaagUcBP9RV2usaeK2Xcj9x
FjfC3r2Seesb4TCaFgiNK5ofqEs2nx5eYw50POYNHCboHAZ6OQap5HnC+TVbn1EJ
eGnlkWr4TiWjz+7kLiZ00QWiSV+PhyaPyS2/aOfogIHiNfEny3k5JpCVrEkY/g13
vb4k5cT1CiQofnPZsnghlzlJhd8knbvuCxbZn4rnEDC+N7GdtpM2D6GkD9VRiEnl
WGT7cGhMukgwXb7aNlWefFMSuV9gmSnW1dULcKIlWxmXoBlzTGhxJgPyHQmZwWVc
kaTerlSHn6Qj42xUtTnQrHQPMxveffKXYqPRWDJ8tFL4g/dKYXwP2koRcaTrzr86
`protect END_PROTECTED
