`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dK3R0o0/hCcRAn3FplJN920jXs64xqI1Iwjvq7FbPEwL2lmKb3N7+fi3j4xw1PnD
QfROeqskJnuLmSlAdmMGbAAY+qpC1p5bdrLA3EvQF5Tuvirp7QvMIR5eiktdPcXr
MdFcOeUWa4hRCx9mDpDCdFchVuk/hrpHT0To3GvqVdR11Zo6NAOYE+LzWHYT144E
5Mqwnx5DjYEEs5Hn7dV1vAW+Xxo3Wn7GkrM2gqYGpk2s/EGUF+lwch0zrMeEBc6x
wuz3he9IR4o4pAcapk8dBV17r8nsYN1TlW1ouNIFagJqscx9vHzmVc+7IyBJUxYO
AcyiSAIUGZ8eb4VU+BGhOLKM8X5YttOGqxQbcxhD/B7gnXkG9ZMYQRsWrGhU3D80
omcf5k/7IMh21TZZr29sOVcr8eV33WyqXOSXyrWlWqOfRVaCWtXFvlyQp5UlRKw9
WrsSCL/vpGuO+r+gOJMcmEGY193rMJuCXveyJ85AAMyFiSEls91h19r9tMhSmNpy
6o118lxfQJYg2OWf+psabXrbITXdWikCloLf4HQBcg9F7z089iqVI9wZPqQj8X1e
4GzXBIOp/WGEoYOiCKU1M7sNOGU31nDAXcpM/fwEPd8uLDK52ORhujDPCF8SS5bL
a+qQtc6wg1UCdr2/LN1nLiLkYbdd2jrX7YNhHERdNYenuhsWhhAkQ1g7Y1zenQva
GxMvyg6S3nDTNJz0Y6S8R9MuGPA7lTsHTVqD/N4fjRkANXjsu01Y9gC9LrUe0plW
a5HSOqZwkl547jKj+72NsG4Q+OTe6ffIKVdsM0YFbajk07/ctCDxG+BWQNMEUd/Z
D3b2RZQypyQ1kn1YQXxqlAvtDrWMqgIR0wP0ahfaCKY4u3qPBOgV+KL2ez2XM3Q/
OB6EhAlLzQUlJUJpg964lSjX52A30PXgRm+GR2NSukF4MPdGS603lrZ4qo0hX/ge
J+azUhCCtpmNBUjYZ2qUM1kbsMzA7L6aNXJrAxA0XgMA42iMJ8JtTY3dgmT+DbOJ
engs6BW/83EMo/Z/c2UWPvvJKO9qz8JAnxve+/2Yui/xv+taFeAAFRS0rCafrR8U
vnlgtO3GTDoo2cbF8rhFpYqWxcCCt7yFhnA4mFlaKc+MEsxHx3ElbFjFubGHrtL9
I2DXjsRg8//m4RWUVWTRCmFrCTkdEW7k79a66/egXd3fnf88uefAopmZ+nhfGeeu
sArvUJWYxOqpHMBXBzwD+mWhiY9heb9xFgmAY9sHD3P+0cOe8URT9Wq1UeX+TF7V
y/zPKEff3gMET9EIvNkKOJUeR/4hD1DeB3Y/H7lxLmVIROW34d1FINYRzJ4rjZIJ
NZNwuW11khyBepoDPhaHK8uGAGfBnmSA8x2jJ1r+1KwIndbzFaQQ8SI9Pxm5hVDh
9QBUEolBlO/ZIQPi5/eGY04xUWVX9bZcexxAV9bHngpzbbiHY9ETW4jiGslfSpAa
s+iOk3HzOxnm34PYsWoJDRWRSFKtVdPcyMcCKIjmoc3ILqq9urD6pLvrtNdBmMTb
deOOXGRgAZTtAi3suwFS3MZaw/U28E/AfEaVOT/cwCQgWONeTvtdyPapTs1efy9H
K6VnNxHCDob+tkQGbq7Vn0wIcRyEy2Y7C995hAeiVVqidF/tD8W5qNtUOsuScQlv
5kmqdvCaUk+PPpij6NEd6tNPOexcRA3EljN2MhgJORqEt4sL61eEITg7Px3rHoLo
dpw//JF9s88Q7s2vkhVwmRtdaOiqeJbJI0IF1bgfMGcVZp5RarNWqCsdi42NcJdn
+gx7yGta9BI6i/7BVw0GK2/U5rjzaQlJ90EGqKN/hROg0tQ0l86WE1l0OGAd2nX2
rP0568YVXjouNtHGzFo1UxudcWmpSawu9XaFKPbJrlBU+2L88NOg7G9vQHhRzbom
cxRk0wk4uGnMY9LxIZ1zgpS6ErLlnfk8Id+WVCIOi3XwmvkM8lGG1+/VYWolbU6V
jP2GETRPyYVrjdlcu9W5VmzQ2ZkjrBMWKqxWFclogPGaJumrNVxiHIHBtsnnI7ni
j2+Iw4wT7VEn+ly9OJXorTaCpZy8lNEbJJ46tFEnpSojwsdcUp3sn4N5YIB6f+jC
Oi4gmdCWY1lyCTXsbd2w9szt2VUdEn9L7nRe2+sy5hQW+AP+rybCn/Ua4roeu4CQ
eTUKNAYQCbYxswrUK/L6PpLIgYDVZo8yaNBpefB5sm/TjtU5IV+9nn0R68dyiDBe
GBM1KTUNWJr7SJMs9gpb9R1M4Ag9qwfi+5tEvOUXMuBxGy08idtKdRQsLi3OMnHG
A92ZmOkwv95B2Do1exc9qdZLzz+L5+VIQIrFAou1tkKOpXdFHN5gd/AGsY6+c52k
tfYUb4liTMcnyOOUNzMQF9OgcmCMAHYcurfrCRM544LzjSKyCtyEzfx/lq66iqh4
e0Wpm1KanuWLm5UgdQqUu5XD91ATlflUpzq6+oY4Hn+M413QxHtbXcKhIzChL3Ah
YvouIwtT+L6/zVMi/F6z52o3LHkgc2EBTZsnfjTu1VE4XgIALRk7A5ogdgjBmu6S
obres5F/5e7UhqDvgHe1rA2lVu2ndzNV1Hl9mYWb3okecs2zDZN3MD+Ge6ALWi+e
0P+Rkw26xQHb8Qj+QvoLMr3Zqf0iPbDv96tv7CPRQh76q8XjDLxmsjWhUopsYjGo
3PxnQsNmQlph/nJ52gLyVsNGZkjny2pnVwo16l4WTp+jvfPSHE5OkY+7+eJP5m9/
59UqBAOpFBZAerH4uiQ0T1z2SG7ZWpymIiVV1Fx43J/r4XEcF0JYFG84K6GVUC7J
VbJTO7KdF8+9uY6+DtvlsRQOLCwjdnVnW0+7eLF+8DPEhnkzNID2VH12kFE6ghHH
VZCPqZUYlsMrHYk32wPkdwsVP97OuaHh7OgvIKAJDKFO/GFsr8JiXH9y6wuhhiJP
2Uef7XD3vnnqMY71rE2JKysABnwOfrrV9naP5qaG8UyTRlYg30wNxn8CL7h/U2O8
K0xXoXibesRZxepYsMyby+zD9+PolZVqS+EDIBPwPtsJVVdrcvUl8kwcTZHRYKTp
xkFRbrklkOr5ELQgeKG45AyRhVKEB9EDX2rX5ZJE0fJ1R+svL3Qz4MRSoOe0vHSl
absbaXzqvwxCqRXHj/53XXvcuj9oyLzusshl3EI4wi3qMqD7PWK8viEiYwhLVqhq
AtfD6efNKRprfareH15+jTVWdP65O23hMd7sVhTp6TQFQuMKpReCus2wst41Dwv0
UPuFJMfup6llar02JHJPJBXFoTKuOmVSkJBcj0f1Ok/UVTdhwbpTF/3pcjndKt/Q
nm9K8Nd5+bx5QrFXBmyog/Ybm68ZaC7iQ3r/R/OCM0hk6aFKkt/OAzZFhqEJ9muN
KcUuQqy84lUdKVcfyr800s9RNafID3nr8NI3jb54/Pl2sMLex6oWKOGxN5ivyzap
WVe9IZbrDcAG1DqWCujGGP4IEaZo0sAskrGozWgqwbuUt9dndBGjbudZMQbwI+EL
PSQQE6DLjhQnHkD9FnEJsJLrUyukLxQmcWT4sJAY+FjogFJ7n8L8IiQj/T7gTmFe
UrUTg1MhM9GAx7zbwIfHk2LnGy3QtdCREKGGfHm81U4VdcnnEcXGFeQSrttrk8Q/
+TM37I3DHerJtsCgYy1hj7AoJhaNoKw91m+oY3fm0lw8uRe1qSSXn7FR4q/TFTQM
7ssY2b99Rqv+jn/R1ZpRlEQ05PfcV8ubwK7qiikjOGVz68mlvrOaXp0NeHqquk8i
inCa+FQsSr6hEhxeBDcK/s4SqqsUOuiNiM7kpFQoAcLdYHAIDJ9Je9K9NolaiPEM
4rOv5ji6EObf2qAl9PPeMpq3OROPMGAG4zfFbZlfyH/nSB7fbMjQuqGG0fYSPGMm
Y+Hsn4UMEQTxjIPFBgh7876557AsqT8tVRV0CxvIWBbaFEdRNlK6AXyifDMEKCIA
GdOZwZunYqLmASHhOLJEnfpf9IQp/vuyFv6/HAQynvKY2yqvRKBLU8FUySWP2K5o
TEIh+EF+D55dcYDK6aiZ3mLa6U2y4AxAY5MbFtA6bKRKd5tqTU2KaYZUP+vH6043
oEuUsCXkxaRV0mYeeqmxLvHkz7oNF+8ywUjAWnXbSZPASiwCVnhameg3BHNVWCbm
8bZs9fylS2kegdLI2JokMLBwDADSOv4C/zbt9NS6ioWoa15Uw5UHC+4MHRvZ8bvm
JAXPAtws2nNMU5U75sdVL0ZhY8Qftxqc4yXxXQFJdUKcf6R9SA2wBhVZkVFcS+DR
ovpHyHp36tVC0HaRs6qx0YXi/U5gHMbqjDaor2+x3Mrw8GRfXYYgHm/6J6T/8vO1
+CzUbFnGFCzqiI53G6MdWlRvuWiBNtkv62BHgKZctIqBT9M19/qJEmhcrmdnn0Yp
VyENGfPbVY6G7YcljVIorYZyfhMD/hTQzN/fz/zOuT5NCbI3yodNfVFaHOrhLdO2
toBqN8a9f3aiYalQaIZ7M0z1QfTQpPwQ/jmIizaXj9cqgatwndVTJD0jF9rnUIxB
QFaAp8itd4o+zpei0P55gDr6dTY1W0AAxxw2VW2zZJPRxd/ta8FAFJOEnpuAx5So
R25H9sPPf26gDkoa2dCCCdSyElLFcm1o8Frtf0MuHQs8UJjRHCWMjbcvdhWeUqnn
RprZg2uWEaPUr1yx2u7mxfH2Dq3B3jaxM93RviOZ9+vZ3sj0w57bqr8InaR9G8N6
C0aThiD9J+A9IRi/xEjrjDNAkfBUJJR+z6IrYxBm91oEnwrZ9hMzK7JSHgfyK0jd
LGuBt520NI8adlIsKsoh1WOsierV7ogkUaQuCkOrYfu8iLdW+7Y23cVKr3RsBQLs
uRLAFThvHu9ipXhSne+aMTt3LbYmxmg3Z9Dq8vLsT64QpyasfIcd0GIt+ZoYYttJ
3JnTg5WmTw5qW+MKG7zpUCCUlObtf5usOHpp5AlslbO6ITtD2FGlriK9uUErbG7P
iCty7RMakVQrpR/UBYxR8NHYbpdhDJpw+fO/PrKLTwZBCfui3qBhehq3u57LtWYu
4X43OkFCZb7ha6pAF/g8oqwEnWpfK2DJTkADM4f7GAv8ygcwmef+PmUcrSUp5OnK
z+Skzr4rmcklyTJsPv2DBFLD7jDnNM4tdtrHgzm9EEXfBnuTRscsloxg+N9zW4o7
oeO96pYsfjXFQ154Atw4mtk4wRXzSGHgOGYP3RUoUd9BAs3ZDEtiUwaZu8crD2mu
YKrMwa9ZVa3B1u3MpYIifNHPm1BZMl1XMu+U9QrnBLTOXnnqHvEvMq1nP7Eb3h9H
+6qPSTrvGCeQlhPNoDFbF1i38gy5vDCSQV8A1fhXdskSgUirxzAsol6M7vxXx3xV
uiEJANL0hZfVwwG7nB1vsNudNPm1bm7Z1kWVADG3fmyy4Ek5RxNBETodNSTWVXv2
OO4ohC5turgf81jwpeKwQspmkh9pcK3ycPCB4nr8jNpmVFNqLuhwyQjBlmz/SMaY
DfWs2m8jvvEpfV4f5C2Oh0pqTAxkZPpKlE39S4BuLClUPdXQfJHCrBA8bqLX1WKm
x+TRnw44/girtLdkttEAxAcS1+Vy0HAHNP5PnhDKcqeIGHyTNjBFozNROxlnOHta
Su8xif5orFpnhZ2ynPeQRBKl6VIow66ZhZTkUr7muid8EjdBnQsTKCVIwOSnIe79
Y5DMgwap9VYTL7pCbIquYsB2+6vxIYtAgl5MfrF4Bu/0dhyaocVSNsxiK0dpZoVs
WC9peear/ciKSdn1HFRau3KlNOlBfU3PhdfBhVJoRzdus/9Wk7tN3nem54nkl40Q
1YjjSTjCaYaATuV7h2GkI5C4rp5YRS9bQtIP8sxjVSlvAziIJ83K+k6Zt/8slsyl
yMMlzLMe3gnHlkgkBXdK9B9bnxfkiQ4891miObMtgF7v9c69jxnmX29jaTxVS1eX
z66KSgXaGsvQZIlOaOjg7iqpxrYkLfbhjQiPOiM94gTXiTL+mBWHpELyKrm5pzjq
spct8qIm3Q2BWc37NYOiL6T9E5tIwh/MuAlDYjh725RFL9ZKKQpbQX8M9zitUa9y
1K2C1HOIj5yxozxS8OGZQueFDP6Zn69y03mENX+f2ry3WbYqAD0V/1LDglMS8Cxk
80GphuYbrd6V2pGiLGsABJewAog8hG2qi/no6EeksPw2tksUQgutbD/JcO9UoX3z
2EJdsxgqx4WzKcRD/g+3TpSQtwntXNmluP3X/RvD8pWCpPqTbQmt4aKmGqIw6N7x
DlZG/xa5eS2zP4ha//DL5BXyzCwBNuIwPgXs0Uz9/korYSz8RaiiwPvQI+UAM3L9
RnGslfhS1p29SurYF0HpKelO6Xbx0oerO6gQMChy4lN3gb0IseO8dmln3FLWu9n5
Fw0dOx33hLRy33MGdBfOuL2qubeG1IfL2g8jED4OM0BlmODL1xmkaLmIOS2MhR3Q
YHmJwuQJ3AoU3PMzh48d2tQxnQjcPogsf7vUEceIqc6YMXcESO8D/YfRSqYpCnWG
MA10rC3HrfEEHJBxYboVbl/MBw4XSZhoDEjFfAtmsO7rlPfveEFazuWw1THsBWYd
NdlarmuBXqvQ62w2w0nFhh2ENpTk9mekDfXKwKwa011kaxm7KCuYBRFE+ShK2KS9
B7DJSJzKcEydVhKfD8ksLgrYcN1errjOpO/8opPlmVJ/9ic5KXRorVRzkaGEo/Hv
j5zzYqgz5dnrlJndPKUKNA3638DS2z0MWCHiCK/C7LwQPuuXrmsXhhiY3WxMSB49
X7JzVxgTtKZ/3wLFQUD7I2Q8G6rkmsrZiFmezKSiptlMbj7K7BkHw23mhlhnryys
yveVXHFIAXYE8UI/spYvHx8OGnefzzDYS+vuxAZzhj2LAoj1vZlbmOB1IWgfAIyC
/2O3IbJfUEwTNAp85ZFkpM9PawZRDn4glCrIfPP3ZwOgM6zOkGG1S+hRaqQgbIl/
PU/Sy6wPfuwjebJ/KZtHbq19IDQclZdCBm/k2cU0LkADZXj7nXewT2jw/BVpunFO
rPthrLVCc2MZM7G4ahfiiKgFpLK1/AZzwpS9P33Hv9hwXkw8PkLeZpCapFh7Q4qJ
ETGUWOQYCRRiAYC0U1scx9lQ+KbGAo5RdGDzAViTGMreJ3aRCqT8lGH42U8V6HZv
8nDQ1vCbTZbYWynPnKiTdpMacJc+IGVBI5PE0me7lNsXYAODuKbsfnT1j4MXIHGR
OAIipg1LG3422TuLX4hHbmvroMTDaTud370dVyB9dH2oSL/Z1GJnUymDBuraHQ2t
4FUrnXSrfG5limAXjOPJlThQDd7YGbJdYZ0hwrVtN44IxKXO/EqL3/p34wAODN2i
9WinlONZ+mEbNhpdXg+ByFgrG+dJQSvayMv38qRYdn3W0Zc2lS0eM+App0y2NXAB
zHUNI05jAfOtXBpCrbm+E71WaZ5DJ4VBgCgjkOKHren/OOEhNFYvOeOk2qLTQlgE
UOZzSwwDCrkIB4KTVR5scc8U8RGeJTHehinYyTiy5KY012FjOZ7P8NJwUIgRirxP
H3P5WGqwXHRMcEU7EkehFjB7xOafnCLy2Do1uK+KzHN4iM+BRrph+actKO1x9xB2
t7MD4hIOlVlUpcJknQ1oowtckpqDyB9D2MNa1Ig18GZAyBiT+ifWZfOZBRZgdz1d
XAW/bzADgywj1PM92VIcsH6fUcJa2J9KxBEmMhrlzgv04mW3QbIAU2bbn8V8qvRM
2PQUu/o1r6untU8sIcP/8k4zcZ0769okIHV53xVvCHvRdZkiQJ0ALZ5dXlGecuME
9EZj9Dy9/C/DjE9LUqyCjNCj6TilQ2R6R/bmrL1HV47UaR3udopUa8CggxQkLToy
zpymzi0keuTeqiRWRvQk2lLQXYN5z1gT4nXocurkTtCxFXomlW2mRmhW7WSbjHH7
lsc8Fxu8gbRepiF99Jju8Hf3/HAcLtJtt2JlGc6FFh1KHCb9ORaYi5uxWD5zW9Rh
M0ha7VLocemV8iYoqUuWQD7prOah6U7iRIhSavuh5J/KhsNwvOe7ehLPpBSwgITe
rsP4Iejkkif/LjrlaQCwICO3nPizonbKVJYc/L5VZtQ038md8gBas5pmi5dEWGJQ
sPPIBkqT7ZEfqT2PKh4PxfNll0clYDtyufKGpD4T11fwxwzL4PRVZXi2VjYNASt9
68qH8grS0Cexpe/rd9zro4bPXxqkvkFha255FToMIZcaZdjl42ERe7oHk9N8zdE9
7Gqz5FxlIFIARs7K0v46WMTbbAWBT9yVtcWvQbRtJP0iyn/6znppCWuXTLN4IS4V
YQHKW3IeuaJ0XEPt/jNiJluW1PdENCeY2QSYj73jvGuTxHmF8J/AP2RmbL4TT1Pw
Oh/ntOVpaGo+TY//1nvmahZKNwyeQB8OCVPbUOtmPke3YTMn3yc71y+/eCYQHpr1
zrB3210JcIVi4If/m9TBJTxdaCNmfx5/88lBSnEDHiXhsDB1Z9/8fwPcteSZW5aD
TW1FWrEiwy9AjF/qghp7Lpr8+5K0jhfwevTNcPSA096a3YTRtI5/aTNieIL+1ouj
HDkZusAW6Jm1fI90I9pzaHN3otrawlkGo1AU3T211iaWX5SIExQgNkuvaiUlYZAL
DH4/fEhwjmpcLomvbgbQDdXNmvJvtE9Hvu3E3BwEymhjpvrn7FoRx/QLmn5G1ho5
+wkbP0XC9AWPkBy7ayV9Ss/PSH+sU6OTdIMcydXHQAv33J8c3CroJ07DXOf6z4We
dmwXtgThUSMwiq6BRZyFjxEObx2O/daoNidJDyrV5b0mA3DYEkndHhQ275+65cyv
/mFJr31RFRFiw3Al0DwiP/xyIn119w2BTc03YyYklEqCGMhlI3nG1Ya6CRneFGFq
kCo4gVWgUe3e+HR0c0eCfHgw6+468jSt4jKrcOmtwULM84I/L0Q5/EU6p7p/1Gu2
kkIZiWZWYQng4ahnNech31haPDyW0EIlO4MT6JQpdHbNwfpiwFOidf8ixv6dNk+7
xsbLhwAFiqarulbQO+gkPV6Q3PJGOxhdGIS15Ym+6QrI02dwC2E2QtRsRtq9eCB+
b5RuFGGwbR2BXvJ5D4H7LBLyADCIm87vNkm8PjDqvkw+vQfHzU8AykdQnHOf+8Sq
SE3OufVFQn2sn3FGDCYMNUcw8ASxjRMtY22MLneI1Rwc57uxb76RUXy+ikWZ1KvQ
vXYQOtOGwakGL9SrzLCaawQksBRtmcB1yhewZjn2F0yzi2qFjGC1k6lXhlVAZ8kG
PctxgNf/xIgg5fmNuiFbdjLEwlMH4z3Dm1ntAxjA1d8/A1AWRd5dOuaudciNCYIt
/OBClwIo703VH1VjKiw0B1/tsS8BWbUhAUAC/3FxKYwcyGUl7/vELGefvAaZvm+n
MWCrro/1zbKFbfctV8nhiuq14O5tq3KkQtt7vGvCQA4nc69GhS0k9hlq0c7yzGs3
aYiOYd23+a5ohZb3S75/4e/oCALZlqhNTKsgzZzEeFMgw2Qd4iWAscrCXy6ugDPs
PzGS0iGZAVLn5yjd12L3yp0333DV8t2w/X/gfN+0p49LYIThzHzQJHMcl3pcWPGW
XBZgmPad+rCQoGQVsp0nc7uJGak5FENi/W9smYWFUdMfg3NoJ3wYxpBTWUfAfuro
Abwo6N8py/XDL2yNBJff6XDUYeHr8QzdE0IncJ1X+p082SRkTEScbumYbp8EyQQS
s4PJM5kxbjz9ZxYbH/ak52QdAoWpXUVYLjuzC5dpweXEHrpGUu1f6zd+e/kdGOEV
W21mRLu1+mFigfzsEbdM53UbnzE+69M6aLDrQxu2j/6fAvWfxytFKt9ww84P0HMJ
x4nvGsIWMyJynP9Qrb3aSymgLONfJlyUEWLiRefiCYiKoeiKN3dbjbXDzBG7Yd/1
2vXwNVziPM2pw3RqNgEGbzTyfygHqpwd9H4Ece35igC9xMLYtX2V/GrdkcTk5ZDE
3DLg90NcSBz23iz1E2+2TD78jRKzD3NfKGxER/vVe6OVUner/kNmjl5nDfw2MScL
tP5Jfqqp0IQZbtBJ4nuZFFQtG2wIl5nFdlTHVxO1CCIstujYdTLzbFwuoBeujIhk
t+mtTCdNMV7M3brKQv596O4Xvp6zFh1n1NlyLrB86UZPD7sen/8N8ts3sj6NZR4w
f8H0emuGQePn0nZzL2jsZwsbvVZi2BTBCBJYyVQQul3RuZF7DZFEvr2eRRHtmmri
np+RmgedNNjT797glpS5+4NOz6F8/fpaX6UK+XEIw00MOkflCpBbWf1oUBDN9KFp
ICuTK5zrbIAHwxsAJYr8viKAI81BhOJrOHLz9FNpvTfebTwM/DXoLNI053thTK5l
yh5LvrLpgPuQMv3niASlKibKjrZXW2lVepi+tzgLHSuohVAWPC1UOB59nz/slqpc
S/2deiLO01uo0VcBG5+D+b0WPmQQQl3UB/QlqfF0jwAMuSExKdado/mo2yCMEfxJ
7P822Auc7pl43hB9tN97FcGk/UzCcG0BzJ2Yuptr+MhIw9QbYrMpDtXht9fvUAU4
O5ReZxS6734uBSnCHilFq6BCgMJcYWvA9fMDtK5uSjrEPub1fJ8L/D/lQgEeeMIj
lSe7HGcyQsTwdkLbrvAU8sADohCWyvlP305ocKoZZBFM9CRB75Nr5tRHRKUKCM0s
T09rpKZnpbHS84immOiWjHhaPqUNkYHUMkBnxED8MhmzWQah6A2u4X+yc17zfBqd
UehabtoHMbx8xzILabA4RsOlBjXKAW9xIDXj9oEBK60XTEa31azEA453m5daaBK3
idiAM5DFN50uHMtTqkOEQ7MS1ZJgsZ27bhcbVYdPKnln0zT1sM1l8l3gbCGibovr
byCPfmiY2phB+WYZ+ZoqaartExDa7VLguCuQQc7i3WHgC4SZ7mfR4BWApr37sjvr
mG3e0+K9i5B7brsdT4QVEd0DHvIlINDwNL/YDmkjnA7efK2VQNYrUmzul3zdfp0i
W/iDsaq/hwfINSr6mAKUygLZr23yMiyKQQHTHkaNkSoRTzuC80gtoV6Zt7hDHE7m
FipXLGQcSMvFqIL6WwNmm9afJRiidx5wCvlPagukKlgLQzWlAhPhWtBeqUPEpQUL
R/fZ4Ur7SGlXN79lCatBWNc0Mhvm/6jtSVsSTJ5aEj7Kf9EWeJx2cAu7WBQxjPMz
U2O/KYTPUs6ECX1ChadSlfGNOe20CClQeSm7Y+sPlg+MAtuQYoo9ivCQ06NiSCuT
39KC+tH6nUYus2sPGyVFfPYfENQaeafo5BO0MGinkcaZvI7+0OcV4sXHL73IMqQW
wyBjL6tCO2qysbDVZS0EPAhNSytczXekp6XZmCFEo5thFQJEpeHt6N2/73E6Auer
mb6q/sE+rONsbQHGkgwYJotyxgZpfztt6cF4Bu6428XN52JgH7JYXsZf3yus/xk1
T63CEOewsXNgMOEbJv5Fdr2Rxld+ZU3pD1Fnz/NEFYog1YBPZPGwxUGJPlhDF1a1
qFrpJT75nVFW9NFsJOg0hG3BPh/UWK0mqNKfpXjE2PJYbMo1IeH4y7986YHC4Z8q
nDJxUrYBk0buQCPzv52m0sdKz7/2n44KsFr3ZvCFzsUb7oZ9m16mbNklP/u2JwSk
tXeW480tYWXc1OcmwWxJkToTMOS1FmfJ2K07Ru5CTUPVj5FQ187R46z4Q2fzaI8D
oxwiyatHVRE2yOlLg4Q8TQ3HI6HNvIJI8u20CIDcgH/s2WoP3WLtyRpxrBIMam5H
itS6W42uMJNyvGTnTB6YGz4AMcsotCu0mZswbaP9DgGetcGNqDmHyCgfCCaOMq/j
ChUdNaOZvfT8TgmlWg32tGlXqn+9o6LiqFOTY1Ecf/Dm9zWWUJFwb3XKk6spEN0c
kCXqAvKm08a+U0m1cUGPHXnFbeuIEu8JtzL9VbXlx3ZM54jomYAwrXCVQ1cyUeim
Kbtq8Kns2Vm+li8EIM2XmLrw04sreuAfAeCdCpNaBtXq2BfOQTojUyLNgGHy97e/
msvyhLCICnj9YrkU7lJc9MfQn3xwAyOX2YoRMTbXpyO6x2BFuUr021Q8MhcQK8TD
RdESZjmuhhuOup7kMZgXaeXGnaz1HrObbueerK5BSJn/9irW6z+7g4n+CW2rlMni
6rQKL/Dcc0C5vQ0V+J96XY8b5l5DuFLwcdBomu2KScs8DlTs+lwLE25lWDBhfuu4
ngYGQz1U7RaMWzqqhzdAg5d0qVnmtBAXizlc9sY6E4Nm+H7J/gCsLGrY7n3dOb/Q
WzDlB2eSyhqdpWCky+VakrXq7p7kVEid2WD/YseE6KEnkb8Hqe5Ln8UQipySV4XG
GePAlG1UkuPs43z1MevnH5U/4GGi4Y80JLxAWisqIWgZiDe+wkhrUbXvtSvxiWWv
aIbKTkQ4MDOdLnZxF/I3Iyds9/IPV8Jf2E2T955ZbPMAaEUdUKZEmx53gl5+KAQH
Q9zvTrMqU9IlaOlFc1slN5Ic8T5XjRSqAnGAxlOzI9Xye3npJU02f4iTyvhhXa3Z
yBMUOU9tjPEIiMPYkVTcn/ForeFajp3LNaxjruK7O2li7VSG+9mgc2WIlUTj77y6
+GmYmk1MCOdnbCpaMFPdxe9eNqewrUCzvUvJQWYKfDtpHg/zfpcsJDTMbuXNbb8r
SP2OncTiYjWuVDK9594mESsP4j1Ag+MZSqsipp9cww3w4tjQWekO6b/GgirK7BOa
h43107QKqklrdSk+7LYPy/8fg3o8V28OFo0nAPUJTt7cB0+bGGUVXjqBVpzS+dzQ
0dc3o0vtLgZs+uyYbcDshS6w8ZTZqC++nuzp/gRtZyjZI1U/lZO5HSOMuu0M7rsM
ZIP+Z024dNMKvQyLtomCxjB0dQaxcbUUI2Aef+IE6LG8E3Upq0ClOMgeHQbYPILv
i/Gbs5myAkvzbg3prkpMlozrIGDdfETJkAUvdERT66hIRbULxSGZfrnSCWagiMo3
5/87FADTNqFmK6ncToiwgx7bp8jFBBcbQYVyeRY1IQNOa3fMmwa6lSZA1BU5knr+
nP7Nb3srCdUQcFY2ygIxLwGkqbEvRO2s2Jiflq76jqqNSiGokuKC7iMRup36bmzp
hSeSMNz3+gOAB82yXnzDGWklukrK0fApQToZGnz37D6JXbm4ggoIHoWhDcywdu0J
K34oMLy0bTUQmTmqXuLtjhiHw19m+mUUJc4UHeE44VVOCFAyu9Pw5040bEolp8ia
0p3I6oleu/xchsncPtuWOAcXIxVEVjntR4jiEul3N/qj7aK5YC37Fi+g3okIVV5D
q6D5d/5gwpAOtLwydol5ufC1XpUbKBiFw+lQaeOKCnf+N2B5t29+v91WrOulxJ8O
ZsjLB63jqfBJaFGunymRkBNQcE+g0zv7DilblB+h7P7hTBcHtdNbtF3xMHqege+h
SKPqfnQVf5kL7eZY12ePt3hI4m7bpIt+My1vP6kCH9iygM1yzIvPlNHEtUozFNGP
nxQeFIFY6KOp6CLfxr3iNlLhEaphbV0lKZy/sGXQ+C6uJpZYqUeZDROjXQMuudn3
O4WIp8QQUaY2TDFcKsGRQk0sxkbn5azrgk8ZR5dmDXUEG5BRcalEhmhIiyPTzLZZ
JHzsqypWldEOWzOIoL6GQUYkraJVqjG7QABdrmdK4gmkV7mWtfOsIaX8uuGqun+M
LwASsBl3ZwJh9O1idpIDCcVALsiP7PoDRlYD3f1xHNtgQjbK/z+7DRLspCHd8E1h
V+EZsSXV6cxWaullLr0UB6E7REI6+TqhTYghMgnEK2hJRbp1ITjyTeLAtvL0u0el
fG6n3rlGZ2KLxrtHjQn2hx3p6fh3dy5l4yNrjzIbfzB3r3O0H0WeJ2j7lxO6uAa7
v870DgTDnX4SXYYGvO/0PvcCXD5ote/YmPcSzwZB4h28sGQaz99hPPGBw22Zql3p
5uB7R/caErZjLHubIYlvIyhF3yBqSoWH96nF4Ur84Oezimj1zgVoDPS1do0/MkcN
/pOSWAghUBZZwSgaPUkmHB5f54N3yTDfQ0r3ihRUhkOwLsf37+AAi6JzazHbgQef
7abWlX8EYv/wumy75sLkWewlHJTP7SeEbbyK/XN5sC1sCt2ChX+C0tXo5U0Dn+Qg
NdIrtv3iDZlewOCzoH6tAM4APzugcVzMOGDA9BtE+3PqGuOWVnSLK5ObMtqBxfh2
CC34F5PnEnx2UGB8u/iMS492nuIsSpNBrAFb3xojjDNpb7ayop4FxAw8gKNWQzSb
JMXw7xXQXI1n/9ah+VU4I23GqfcQxjTCqPVJt2l0FgwgkXYJTXEba1ppoElV9kTH
HuuOC68r4qU8mYgejhpOg6IHoX3iTZM472QgVGuCSXlloQUb3V7cBVQGRrJ1fR1a
/KFKaQb8A7clxatKDiH8zjiFUG5uM46HOIjtHkHcS16BSg6gYKKuVNuClUVOXdZg
PZu5tFmJe6Io7XsQtm2y/VUoZMN5OxARqwauUuetqFnOauCL0+m2i5cSv8W6KtCX
kkOQO1SXETjTKXzGRWt8Dmh5SZVq+SAJ4IlURUhqemBFp6KwkhgW/yFD7o1vJ+Y7
Ez6UVJrlmKDb6nQK563HSmQWeIXz6KtcNrudDHFsrttt3/PlBCcGZ8fWv68WOIQw
9xUkApK5selkcErNowEeN+jHORIwqXapj4+02XrAXuThdh7UlJGJwxlqdlw2apWI
xlTDdCnPWjmT5O75tDr234OjpWwzK8FhsMciKQyI4TiZYFbD9VE/bGq2k3UxgvKw
wnhA7AeDxQsjuK7FTCHfUBJ7MSmQawgZBh+kvm6loKcdYtTg7Ig2cJSvgz4hh5kS
UQzDR6uMH7OLzHjBwOXjQ/fkUyVeWeHPvbHVdbw9Irmms2XTMCgVdPYBiypy8PZn
PE8e3qIiOLh7ALqfnRqIKyQkCJRrEG/FdxqaEBty1KW/JwbUaC6UWJWcwb8HbKx3
mhsT5wF9tc2WhzDsHqvBcS9CPCy6Hx6DXYCqFHqlltMYrYvn2DxlQgPMhdTn+Io5
rU+aeZxEHIXIORoic7TWET8oag77IJLoBu9hgPRSEVinx7Kv8UmUBBjOJfABYObT
MTCjruDkHjNpH1yDGPkWk0ODDVhmrfkLntCucvGHudmwF9bYSaJfud90JJg13+nM
Hla1z+rzhz7uxySSyVcVcvsV6PtBw0njU0T5uaaDAApMikuTFFUWCiHSf2ey/qwA
YGwUkR9S6kH7jGJr2OOo+kBGT2zS59vR/Xz0AxTlsrklLWVcRiCHwW7zDygrLcVO
bQACVXMHLVZ+g8ldueF42VRqqEtsYZm08qu+UeHQaAUwiOBTGU5JuwlWt288l3jW
oC/Su/rtQaC1GQorAjwF9iljFPfL+VaB9THumXyBiwftswxXvnRo9Tuur8+AxCUt
g69lqtrZ+BhZ7GhMprO5m3ED6hFvgePWnNxjTApEwwWd78Rs1tBnRYv9ur8kkYJk
THhGmqw2iz5itJ6kpLkBpEuzDGIy55mbM3dUS2T1vurwpbaHI/RHB1w4Qg5+YONZ
EcwfjKaqkNWLRaIkovlNnCWrLjXpyq3h18QYcIkBTzx3q/u/lkxWAa2V2GtTWoXf
IuKn64OkXDrgLzQ6CIoC3u+DSavBykeaJKCFzWm8qhZOFc7ReEcQDbHFPrHtoGHY
mMHMLj1S3dc4SFpHZPdTuNC58Qe7kG60vU7ygqKU4ggnQt9dtTOPIsawGSmCNMba
1hxS0UpRJLEqc+MwcdAPLJ+ztTighI6E8amBW+IeZGtZqbe0PpVwvi53u2nUHLWg
tU+LLMr0LnR4b6wpjsoahM6PdCkTC2LdhxmrV4hk746npMMEJGwPBCMiGfDQsPHf
xUUx3WkAedIs1NjFBsWdlCmPPafwX4rW2yUmdiguBREZMzybBsrf03BzZaV3MXI+
B/Q389Sm/LoDRjoshRI8FA8NkPjh9A1tu054BOtiWXiiDrZXQ+MDZQmZzprS8ykM
c9UsPN5H/K+87jKXritgjMhBD/qYq6PIPNTIu8OIX1IEXGw4U/pzcAYYrOQyogGK
f2ceiRB6dL7JtTNXVBaG+TytxBH3ijie1GOSWCGeObcVev5szISa3pjLRkZUwwwg
vrW5KLunCw5J9fHNRWOknyZthEBEu6GlEArS6frWO3iwwxZP7gNTby2MSq6GTlNa
XP2ByQhVKVu0UUn50N54C5FTsNgUs6IgmvMytKkLuOPXYFEams/rY2Wi/17H9xZb
xaH5WxVcxz9WMoRww3rEGY69Of7cicE7Ue+S62Duwn7yGNEV3L/6Dqr23btW0t+O
9twi1PKZ1LaWBN2MrCWyv9TbhOIQ1nCbqfqh9+f8+6VNC5LJvihSCwVABkP36QvL
lhMOmF7X04thwCIPabNn+4hx293GYgMNYVdPb2fe/ZVr3xYixwYmri8t2rY3CBWH
vdh8NLJuQMSryx+Tel4MRSy4wrMDW38uhdQH8KrjA+cnI+IMvZSGUUcy2zN6pu1J
S2Sihy6k0J97BOYU5PqXlqF/4+zjzZNM0Z5r3V1f8TozE6/58Pugg1SB/zI+8yru
t7Dy6TiNTIMvuk/5WVZzuAgyXtRY5fXQSN3drIz3/3i8cjaweZBNkcpJ3xIIcBGr
sH7vAV8x54XWqsVrzeXL61qFtSgJYIWFEi+sRpRdcotYJjRVmzVZafX1tks+ALtU
IoCkK+hHRBH1l0sQdRu5pdWYynf+fb5pm4T21TDyaPRpCk7KKxKR0ynFbNU0KMuq
SK6h7LLusZ9qozf/z6Vw3OFyKlsJPV7HoZH2KjFH5xIyZbPbWb4PX5AO3GwkKwae
Tnd5E4LaaNJh0gsuoz4hKewA2MOrHwSQAKZDXs9KpIgaFFcDX1DzTGjYvFDoNgm5
LgXwx2KNr9sB1iX9JCybFTT76EFcwhu2AwVe76a1UZ4hhn6gzFAEGv9GLuCLxemj
cUKCcAwlKoqbNpfroGL4hqNBBH9YwTo8f9ytAtOqjfmsbNfl7c02Kh3W5NTLADFa
8Ow9/zVLiwnvFET9Lfqe2mnj8gnWfC2QspDPD/8MIyhMzqcOE/SHY96WNDHC/zNk
AVrDZ24vpUQGHTkfYIoG3VRBQYvlPotOu1oyJjRbv5BhnpK11aIC2FsR3R6TrhXz
guIRoTx922fFioQs6+6Z8jrFmbFrO8Z7kxEsD7+1I/huiULY6lyDBfbO9eBYc50D
5VFS7O4A8Ih8h3o7LsFMcKIBT1hCoFdls+SLKP+sBe6sqdYbnEmHMoZHPVzdXfUK
zaxnRT7ikCWaa8u6mDOW9AhtxJQzuV/7ZHLwctV1wQtqgTpZ9hxdUfc6ZieHdvPd
aRgZEv1s9hRHre30g5eLM5nBach5tkVyadD3LfOybWPohekmhxYTpX0p2FobJCe8
FqIL3nuY3cJuSnjAyQhPZgMFCv4YGeDkv/KPT0H/Z2isMWIVjzYla0ehEBIk6B/l
Cd+Ltl2WUe5UUkG/sJqD8UhRdFdMybMDNgePjF0vhXzaTu2YWnYcIFIdqG3uYjHO
hi+8GekxX40689mgNrKtBzd3WqjxZjbzriEthNQ07DLD6uZM59waAYWtOxlu/X4g
vfqNh9ia/2e5afSLO9G+sLe2Cvau7GSoxtZBnsAELi1+PG0PJNEp2t2uDwuHCaEd
vX8N1NyGluMfwqrM2NV5c+Um4N4EqkdCpJ9wMT5aaV8vVb0iTqQgrc05fb2ritQ7
CKBgW0zu6dqbicpeXnHWw23JN6aaIjSwWufjbHK9Rr4InTa1XitirHnpdr9u7AcN
RShabgG4CL6cTdHao1hckqVd/PK6AWtNXtb90K/lxubH35jAHwhBucD4Vx2NT93q
svMUDviqJY9P4H5FZggUA3mmc9dwLbwOZHSfu7HqhETlqfLrpaUy9W2fHVoBcTsW
zlhqrHl1ggokU4H4xwKVxel5+7avlGwe2aR1J1MJEhYjbyz3VJECt+SbWDs2vP3X
kiUc0oMxoyXffCegDV5Ti0Urfo0HYRoKlcjuxTODfj2nwo8yozqDj3W5boDNRUkh
qiJHMru/ATqrQrltrFj9sRpg1n0RqYBPvY0kKyRSaWMLEJl29D+0Iji5a9jxOMTf
PiR3/BUEfgTd0NmoHZ6oQ133AOVlHQAERefJsCcTCPCQge/WuR6bsm8PiV1mttIV
acMF5bcacEPXJZ/2y4b1tIqYfLDmM+IGKZ8ks326mjznPuPJY5DxH4/6T+omhOmx
8Zt0xqZgMqAiL7zqDzt7rd5ooLyv2sCtNNnm49ieVf62J0LIHph9BEzcKr+2LUhR
mEpSpg3Z+ECxvmuukToj8sn3rfS3lFsRzlvRqueFRT5d5hTy3jlVQAJpYecyFGLB
3icUKd8GpTvAegZPOYsLQO6ic5b7Qu2LCLSV7jIwsefA887KTDmkGC8kUAxA+GDj
k0wa7noNjlCTz7IH+Xl8NOM+umWSycYNzU5LOnzpa88X6P1SUDIKqw8h3zmvrEov
cg9DqpvFt1s0gM0YAMdcgPSaSToLKPckKJYrS/eWdNakjGoltRpPLZsrD02OG8ba
b2b0bbSPawNR81gu02igdb+QDARz1E4Bd85FzMaeK1PCEO1NJkIYgQx7Mo+jpRX6
37qEDQsV5diatkXBFl6pOPBUIFsmOPJC7Z59bwk6q9ydbrxgYN2ahRBwyC16N2ML
htD+3qrxZaHUwdR9Jk9v97T6h+rtBw8DlnZtxbZibhWGlle/AandxMtf5xH3OcKQ
RQGSk6+wC/FgiVu8gvcNMu95qw9tfjet6s7jAxC3mw5C38ucCBfjBblZB3ongFMl
Oh/jGrYhM2DBjwEcYq9DDU29V+zh6gfUemCX+yXvP3K5g6FLu7gBvIxVMM5PlkUW
cu2WVByEIK81pkdQr6LLDbe8lw1tEoxayrqMeyQWQW5+0oCXEbnQTliSkyObfc2t
Nn+C9lXns1LImwgstbuPgdpVbg6WeB50+k/QPIk+Wkw8AiARY4XvSZOIgJ+4kHXZ
2fjnPuchzCtzdTlnBLoJaZ68pAeAEr8v/ZfcHcSgto8ZU4Q6ElDkclI3wGdzgeAa
QV/vx0RQxYRj9dimW6hhGmaJ2jljqUl/I2sva6d1noOcJQ1NiSglc11CWkglU+Lu
X8eVDFH1sjfYyfUWq6eikBleehq1Qe0bC2bXnBJrlqmRorHxxDtuHqDlL2AA/BdP
POC2GCTaxpX3OnDsf7PaRqcCkbCY3j1tUaJWsjdS/NlgkoNkFW3k7i272FgMo2YX
U+MzkZGOTIc+kar3Dqq8PVZedow2wzzKK4FeJjw/jGLiLThHCe2mLsxLHT6n7bO3
BmiEkreuZiHZsZuPx8Iz1lru5E2F8Hg9piOZRVB21ITRLBiGv3kGuKHkLElYiz4A
9OGA3ZcyKV5oHLuy4Al5LP9UTs0+p2RIU2xBQ+imAtEXpwF5lYJjsZVnC52pkU9g
11FoDV+NsXfwNAQKwJSDLe+2nW6onYm7M31BGd9sx09kSg4y/qaZSjotXAkAYNpx
nZcNQbd1IlVWYCMZ0z0M/NV36c3+IYzgCx+7jkfQTepPfM7R1Kc+oWXrIy/KmfAB
75hZ4yDo1AdCMqxyVXN9NiVLSl1hBC6goacZb00UV4F9fKsnKqY8AjybS5IrePJX
CepYtWIUXHaxX3Qo69VeE2e/59YLF3Kdar18zkRFHLvZ0GGGtiXugzlEqVf9USHv
trRxZK7G865FZ6xDYX2KD7kS0YLLvgbctueUT79fH0a58ZUcWDK8wcrRpMU37V5H
/ZzwbIaUfDMUgdkifa8M2KteHjudZkG5O59B3Cjebo8w8BC1RtiNIw5V9SohMTu5
jDeUWLws0iSNuU0oVBOv8lBXGpXby3PxbvYPFvyoaDekv0bdXfNyK/5sd02zWeFx
xeQ+iLHfJ79cxarrkOHbiy5DluDrhJOqmrnl72IsXcZfvcJhC7VBetNyFRA6IHlY
t3dXNfHwUsNdsfFFQF/kpaLwgsrQh8CPGBO5wqGbkihI1jLyjXq0FHu1JsLMCon9
QgiLzXy5zIUHlXi3IPyXpYwoXYTcF4dLDOdRGmfKYIoPBSAlpDH9ovb8cukd5ohg
dHnsdUWqr0v0lsCEcMn85wWG1j015I86GJh5viLSAzCNmQBP6WkXUxt8f9GUYNBF
OxTV0Bd09pH0v96sk4WOM1eCa24k8OhbNRmryNsM1t1/rQoYVPXJ0acqd8VwBPuL
wHb8v8T/rnH6GAWe/8c5iAi3+iBik0nnjRgPpS1iwAr2KzUWCRnl4svaU6GzweiG
DG35O/ZU5nmG/FXZyM8cggMvb7okLUDr7CtcY9nt/ibBA5SMooTN1K6k0ymj5eNm
5iOjjlrxi80/I+MDwqm9XTTI3JLCfZBLX7XmKb54Wr+YILOn7Q64m+RlFCEJl/Nf
RsuGiSIuKQVlG1CAgEc8Fj67pP0nHn1UKszgI9uhHCtTL2HGZIO3wv7mcT0X5Iom
EfK0VR8MWStYhj0rsX1QshWwqpk5R9Jy69o1pvjtSuxsGFZb/RJ7TWgb0RaA/BjO
194OEyBdK2EdlgVuvmB3aYdEGF2MGd29FSn4192aYrDi0lj4haSr/pUN5tj4XTJ2
T966ucigJLGEDVK7v78ZdN8BjgfMciQNRYZHZXWvtFV6xKXVBU7EooEGu/00gvQT
sY1n9YDhRiMnckj/ka5Uo974niYvL97XLxmp27Cb1Dhloh+if5TNTcOVzZPl8o5Y
bmVXUkNaiq9kMNzW33bHNikbhl4PUs3jn+1efINHV9pytnaoJ14DrS7BnHbOfPnI
5+1CPCSVOn5Z6igthfX1fPRMLLGz83mVOqYk2rINAgmJhBBGhYXW1xZuzZniefzp
vwjv9i8uKQ+ufY+f+0Lx5TMbqbBfE/gyMBYRRjcZfWPnFdJbxnIZIk98fSi5g7Qs
4bHX4mwVABjlZpNvij6K6b+gk/8UG9tiSoTSD7ldnauol+9IwLmrFAuYf+6urYyf
DfqDV6dMQPGZuVvVr/r2YFr5Ekz0fw9gGQk9z7QFJ50snaJdsin6VnMSpSdKG92B
cfc9UDs4AiaugOsGXLjldj4sVhD9MQu4FVsf1djfOoBPOLHJwsPIGWKaZsQ3Zg/3
UzgLtKlWqx8LJTuL+mtaTeDs0k3WH/gm4jMUoa1fL2KT0DDQgU1A6efSeqaHwFkr
tgyro9VcAqJ/erpSJWzJVQCiZHWUrxXy4iptB/db/66WYNDNRWdnP1rrbDb+LSij
gjP/sfs3FvDrzYVmtRvvadVkJ26cfnq6Vx3L4gCt+AavR45tI1vhKkV/mYT77vyy
1tviWKMPG4LYmk8OplqEJJ/ZH6d5BnlAPPccEtl/ZlJWUwtU4NGAz3205OzOViJs
/YiCVbdx17VA0p2O2qaiCPRfXSuiheh3ZE8z3T8YpnHRvIKG4G7in/rxeORf09cd
ydspj51UqLGp+P751YUJtoiJ+LYwVsN9hVdJ0lHH+nG4dHFi96S8ly4s6QnXis5T
atK8xmCfrXZQKs4kw2CtG83KPOfjHzqOtwVoh/ZjAbCNYtb3xRK7HGnPi+ykmyiD
uYZbIYOYhFAPrGLPgyTSZT/CuJ9nmX7DjjAEagS0g/mY/rIRjs9jCI7T0kMNsoxy
kb1+mxTXgypejzCNom3LnOumDphbdsgFAkWu8NLm3BbKXMHZ+Yh2QMc+xXN629OA
OMX0aIvnrXKU5e4urFizQC3d4I1HbXg7oU2fU0aI45OZTL9CGi4Injt9sXtjQyqw
i2JahZshdnvRrGTal9CYBlbeTcyM1e/pTQOHAv+0LhYp2E+dsD9P7lyAheoTNMbW
QWsSbo7Vk0jhXg54S+sfUbLAmSuCbSaM+ZYN6aieIlWaEBcfP5HdiRNTehm51vNa
XWB2CZzVDBV5HB0mjnfCVYN52Oy3d9gV8Fd57cPmiWbeZeLKnFD3IelVFste3iBz
N6iwFOZBZu8snCKw/ires8vetWhzSd6ZxvAlmnoa9XvlwGLhNTpAU5uvIOOApwbo
TsYnkQJTJNKuiw2bngVx3wZVIby8sbnsLGOceAPCJdxbWDR9SLYBUqVvOmtYqp72
hc+5S2hTn63BtFsAZvwU53rH2BElfZRHU1Sh3PjEfH46v82r/gyOYCSdjvzGol77
C+EORtb+JrhgfywvveG8mh6gj14SxNyBwLfcrSrko2bPTY7cRbcDCzWBG8Hcnf/J
dsL8FVIoDoX9+DTHBRxkyNG36afey4g3a33AhIfyD8+wHZqIEvSD5YKkWhjvZgRI
SwUfSWN5C5kusTRPqskMsVTDP3RyJBq5xwpSXj7MIw8Yq+NYL+AAOxeocQUtvd3N
7NDPXZ6MUf/TEIqhubbCLPXkcnxT0ylcnZFDAp0BAwpBLdhnKQ+jeuANWsJQCGR+
Bd/+U9kO+vhe0k7HuvhRiv6os2CwkKhtKLKfySYA8Z3rVvzCPm9L3MBa4/Ur8wie
6d/QUQDIhyPdg1Gfr1G2Mly8mBYOggUyXct33HrrLrmmMUA5ajdauQF+EL1f9cW4
H2pnPxOEew70bKFm4wCTb2NBZHk9XK/mdiyGqRuBqHc48q6skFaUEtRE1bFyTwot
8ZlDR/FeFpnBApzAcLfq8R1nDgf0sf5oYIG/4cM3Gq3+hwuXTMfvzJNWCykGArRI
R9VTfWtvEswZr/gPonMWzx0JxbYD0r51Lc62t6qtQDXPKupi2qGSsZVOQ7B0D8Xi
0nKVsnVJPoYuTcpBgNTcysCUSXl4YhKuFRzoGtYrcuqYIDI/pEcejBsv6YOziIOq
LrKbHMhfSm36aXnVjt4K34dffLcoJaneoCTzCD788YXAVltNR60Ssedka7WIehmM
OWYNcGdaR3Sgz0Dkw73yUPhXuPX3A+pcVeRtp+CmkbwcmQN1D4je9eaTFnI6nyUG
mpTlFReOAVcqmp2emUZ6DT0TFeiiRtsiG6UwrUxt2eeu2gZ+VObNPd2RXsbcV/ZU
FVKqIFVc3nifJJBnhUJgCPFHD26WT7SBW8+G/ywTYzPQlqzmMempXRWRrWv8hcig
atdGDmlcpTbn4eDQkTYHaImjhWz/wrymHRCMft1dJNogZsa9FiEldcU1yCfJzLEU
debWRx2XibaotIJBfPgHSI6Z69K+u2tc1Nw7viabTDJp5tTbZYKcHMhbjFyxSRy8
qd46/wJOTBdJpwE7cKjKVi0M15dsdQO/VQ2r4hRTYqU3SNkleJaQ+rflwXVtdGcQ
BZpA0FJR1dUZ2/FKd+59jsYSTeUMODLEU3F3gTZK4jgtm4pMge0egPk5lCeWpyOF
jbdIHHE9+8UAneUk9d93vwjeWjK1V1XSJz9lwc+eDs9R9IDcS4Rnr02eKckXHGWU
ph5lEqh0MslxwnrKPRQIhdDw62Cmq5tPdcfgqU+fbj5mpPMy1IXMchsykv2wHvDx
8Cc4vEWMf3Jx2KKdPTe25+l5ZxbkXcskuRe1FTbFsVWGqbvhMTMs6QSM5Ibh2stN
Ri1yj9AzPE0r5nJ5F0737Cmua60F5wx1GO1u5e8I0MSyvJXfI1LNCXDmaSBWJAAg
8ntWHr1oNCin1oeVjfQ0ucXuZ9IW64JnuaS8SMVMiSxjLE3YMGPV8WCx3w9gwiKR
Mihw6tIGruHYAAIb3YBsYKMQXJ/aV9eSyc3kU8X3AQBCXLLG210LdzN+pptYqXes
y9bO4J1zBCzVkgei6q25Dk0lFxeM9jQHZAlZhv5JFA4zWkC9OrhdRKvlrshVowKl
5+3mIuE/qSzTOR/Z61etZlTAId0mqk02w9Nzk78qN8qu0Cy3VAsaghIyW1zLJOuw
P6GsnRDHo4pVoEzaApjh8N4UAxCcDy8+HuNpQtrq3Z/Z7B4WKonxmiND4c51bUTC
jgpj5h8Rzcr6aiwZSxCZLYRH9LT+/8rp1B6nVUF5ch+o84FDf6czPmymCyAIvPPV
r2CiTthFZok2HfK/I0+rXIEbiMTDtqO3Pyq4Er9cAZWT8yAXdc3BiytCwZWq1wtp
U51rHb3WyZjwpnfJ9bVLllgv5oXrKARhRrtMRM0y03KrO57ayUfNnlwL8kX/XCAT
LfLrZUDiw5N0Q2jtpzHH2MA0aCYM9Cvr7+yqxcORyqXLU+5LmYYZcxxJTt67umTB
Oms8wT2KrxZFumzLhTMnnUpoEQT779eBrgK2yodJRDulyB1YX8dZ29tLmA7At3b+
BoaiLyPEDtkckjZYsz6RjhLkdC/OG3a4WuO2kXCdKmJubEkw8WhMuXH92FPra7ci
VEvHqGAFQWuK3kxBFcCSzznOrnCkP2UJMI/90ZXXnBJ26A+pdf/aNk59Pl6In8zI
1oh1+XSGSHEDiu7Hi1EBi0yjBe6hIjyTOWsEOrPpIzv9SM8ufGpKN0KpiXauMrIR
rKwZzi6vN9QuJy8Q3JgrDe+04/+ncb0oXe/AQboyaL97f60ZK0DlL4MQdDuqBbyY
2T5/itJq/49QrhslLjObeKlgdwM9J35F7lWGx769usxoy8glfUgMKZzMC/ErlObb
n9txTKhFG6AC02hnp7Pp2exoRaf1h5/nV0Ye0UYF2CMiIZcuJd6+ulAKIDSb/0Xq
xF8LkFA5h18BZuAyqSzKQEXDDESkLaNHBzL7jAaiPn97N0YRYjk5Gpa3/BVmLTYK
2ESJcI/LoFXvQhdOnvpN53w+U0qrv9WSS8uzZs0UUjhERLdlVfCuR93Lox9ibnMD
5ft13tP3kMie+/ZqxGUF7j/s8iud4G9De4Im2IGJioxgbWqRx0EoCVK9k6/3+UYb
kFJv8gQnaLzV2H2xxNSWGxAFREFqHoRlDGkIbDaoFVWOZTmVj5BQLVEWmvLC2Fm6
aJdimn7AxBkI4A2Bo5Ge3pn2MH4Ix6dpo25A4MQZwP3mMUgBZh5Cysltet+CHEgt
hthAvCwq65v7fL4Z6itOjAdUkY77gNHyVb4wyfil5vamLzW/6SsL01vOPt0e/pqp
3+seW2XylPFYcc61Blh7cYz7oGcql6ArMJX0l7ogQ5DdG7iC0MorzaR7wj1iqr1/
pcKDP536krDDtbmbcCm/kb1+e2KgB/wiVJdmp2JgizJHpjGQ8eDYe7yqZhKFnRox
YcvV5NFAYpGwUWw3Q9Gw+gDyyjUYUJLyIYgcNxtyQyNAvG9RhnRhk7/1Y2FgNsMA
KY3qYvUcLg3Slm0/NZezX63oDBS3E0HWfXRL0dBb44IdUD1eKH1sQjSACaQgWXJ/
DfeGDpmaPgBBh5KYs8zq2GzGrAywTVnrTCQTcrY4feA6g65U3D0WYzOM4dqTkhjR
+Ps7QpM0w/UAvetBbcDWTTJJcO99ZGqcAO/8FODNb0LEAEpDQDRb80DoyLVblBFy
lOJg5wNgfmul88ltqwDixtat+emAYe1XQ1isD7MwT/uONwykfduVe0+3qYgV3UYB
WeM3rYf2z2JSlRbpIfixvUz4Vz57nZLeBhfBhC6mhly626QUCeK9Y4aksTtdxKz+
rF8OcrFsRCgLx6RFSssuBKUgkywBbCIQ7XPMZ/sJ3r5YtzSKuFXr7tmiM3TbyKbC
STS53XjUMh9GNmyEqsB8YBGFR+DNWnnrdIKnOKWA0EH6R2GEfPV7uWWzEKAYM/Tn
0lB5dTHrRq3Q7tfM01nAQcSXvwGd9jNUUEABn4G8TbVeaW1rxG9tcQd6Q5RPTZkb
x6dkX1VYZ/mHNSnKK2bAisypfzfIOvXbwJZezCFIZFzMQGPnWhQvJmk78VP1bIl4
kniGC7RqM+QaFp9WmeGPbFazil5wig8R/FK0S1BuirvpmdUbPErXp2EQyE0ipm7I
8e6QSko1RSAasb24KhzdKiDHTLhkmO5ITROe/kRaZ61GyMXfa5yhJgaU5FftYOZW
dAtn+nx2bBX0PIK61rx5eEisUinWS1B8MC1u6nQvYMyu8J6VEC3FT/O86ROkIj7u
ohTRSEz7ddtNkhlDqtlxt5d6QFSRZLJjjjvxiaUlWCLpbqYLxAFmmTh3iveF+4Zl
pQie9jneb0hL3EE/o2WPivLLgJNueukTQu0X9Rdow3m21CBDZQ+QRzLSFAaR1G6R
9lWOmiV8YeCMZWHZZwY30OWTKNDiq9LRFX/JZ8YWOz4dFhuSKrWHkVty7iPZipb+
Fa3BNP1H0Af8z/jy9WrKYP0MO4GIIxd9hwOjHDIhec9sRC7Q/D+E7/XMLRurZhN+
wSYpd4+jlpujDEnV7urejq9tkJVhl8J7cW0+mEcbu6+7HV7bK1TNDELzDm9QTSfS
fp3v20Y4/hTlvPuTNUSFewllHCbc5zW2rjSSiCGVXzLRrlTPYLiqpJm5CZOX4cO3
eS0dgqrtGtfDpj+gDwIQO0vc73tLlYacar8Qv4VmcUwcVK1t4AXkmMWS5QM8DEDC
hrgKGItz+rPt3xWs9hPCXAHFa+TBpouZZ1tJyZn47iNZCA7BIHZ0X5bs4x6l/IwC
e9gF1hKKr3HMPtfsUdh/Zcpa/ieG2cwwO09nnN8kKNo5NVNn0fau3CUGDgQIJgBI
M0ATsgZbBwFMximbYOgs4fuRQ0in1J2B5Uf3KwnAJ9svy3jHKERrjS/csCphah4o
G7UCmL1do05cekfycEwB8Ya5giqOPFP4Fl6vTn0lL6Zta6jEjqHuTw4yoz9ko8Lw
PM1NmFy3tjtUO5J6m2kYbYtTENZ19fTaZz5AIrszSgvZD/wT5iHz9CKcEyME8X6P
BvizmPIxbmzgOpdGYrLvMn2yziM8NLdczbvwPPGOYzypUqB4U1RnEXNTHOZAQNKu
dcPTzpaY17TE0uPDrj+xVGhyXk/7RnWhaAlRGjfQ7yEX19ZaNr+baiXEebevgIeG
JAXTP6mpIYzzw5rm6lcmwzljOQEyQamtQMvmeLXfjwSI/LX+K73VmQp4EgSF+cKB
RAEMuPwW2BsuHScOyJKRHCIQxd4A7DbIRTKruob4AXTTTSVlrtuK3lWVd3LgeZDI
OVExC2giFI+Pdo/Jc6Cg/CwEjjBFC0tOFxDZrAvAKVlU1nWgfG0YG5wsFYR1HuBk
IDyN6xiC4CpL92zGCPb/fnTUaoDgQE84+L9Ki+atXZxgKToMkRY75m6BxYM9yzKS
6+HWnBcVMYmcbhKhFr76btl7pGOPQXAtR0/piFkcrjM74xLuiRdCmjCmiqO/cYCw
QkdPkHZKF4DFkcmnDi7Xv0SmTyHDRIdTwPE3oVK7pPXNYdEMitsAfxx5S4MD6QOv
3727JxbM7nd2YCOCk3M4wJKZwbjpdCJ4fdivOzEptGdeDnxCGnJ7CRdPQ6fopkiS
QrY5aRle/xEMBD9OGAG/C9F20kVUbZf4uS1QuHNy07jASwMtjwYis2JmUJ40kGrg
1gGUzx7L5lvI2znhRKIv8aTBzPzDvNUF3mjzQU+dPdE1oZxUtlUNJhBNL685xMAj
WmqZWcMwyytoN+X2He9bjxVumQGDkqA+PilzJ7L0IDFiDXreWnn9yZYZ2TDp/TeS
z2eDGqhnfrphz+XFnySbdRNirr7syva+d8JaBv2I+eVbiZhw80RMch20bRsHkc6c
OUpuJ77pYNHyO8AqN2ajC+YGWnhZMmoYVNwN8uGfF/afFvYr9Fh9Y4+rExqpSAo1
1VRl19evVuQitkNCQ0yLkWnaw1fzoYeRZDBD0F90G5s9+lBjUtA2OTF2fSEqQh/y
ZcJBcOUFJVjsEO7cwq8Irh/k/ZHXXDoybPG/CNjF43fwR96372X73PVdLL0EYyQR
F7Q7bNeWpDdzjIyKbAH1Snkh/j0k9j2Jgepr9BsYH00l5OhkizHd5QdPpTimcN+p
AOv7V31BhcdUmH5EPPwFjaN2AVc22YO5MpnR4C00lAQUQTu8wTrsjSIEPbfStYmi
jBozbQvnkVW3FHTMa047O1CQDGkf7B2vAdezwRCQNuJmL82LuzTAVYHiUq5we2xL
oBGkmxRtBQx9Ay8CTYxLOkJQtI999ZR/O58v5O7fUrzQaEEXQePgsRKbWw2qfJQq
s19gqgQZgg8iNKcLRHV+bun6dBAwSkliUOmFzAWVZcmwh8Nhow4GLTEhHuHtEdUf
69cGMlbhv6ECMk52pQc/Gf06AGkyFxTwA34qDjyNxN/4QUxfERzHzd8FKwgI0Y5S
j/goI1ruutM6Jb/YqjXrVKIbQaZBDrQ4YNgWa3YXEG32WRL6x1MNo21yaeicL2tr
TnZsRl4yhfQS2ndLhuI5T6/FrwGPQhNmKcBpCnQOnpqSR6ss93y219V7/1bjEmmi
Ef7MFfLpVsVb3B6vVf57PzPiwcNq7j3ud1T6APUax9dPk2qqeVUNghcCgvZC4qeF
D6Qz83Jq8X5GIiXYxAtDIaluIqobAD+eVbqCvYiHD3JYXadhMDiPKPoGfHrZzENZ
p3YJs8i8fes5//6v+4/4Gl2Ksqu5k5igwTJT4yza3GeACKT/jA/dscOVxGFQbnpj
x0pCfmXmga8vWCN9rJsdl6V8HwfpG2PFrsuJrir8CKBvgOwu5olXDIjMg9XphsZ2
74G2ESq2stCSDr+j2TpylqiyXYQxBz6dOzD3jiqQTVdkIwsHG36qbUHIhoGGQUTH
ddR1Zzjj0sQJLAq49uReWzcQr4m77YdRVuSBlQxAu5Wpfrepwsk0CSOvmaM/IBfF
8l12vt5DAIo8L5dL8+6GkmEYAQRjm5vpK8XAP8oNCowciz0v3dqcOnqmrQgdBevL
af9PpnqXfZ64B9Arg6zZcajTSjzA4znfoUu3foqGxc5WL0P8yfA5ZWJjGU7+5bbC
UV46E/x8vzNKN2G2RU8S5RFzIQ88CPje/yLUFsMnWoHgTSf6Tdp8LtrRhKYnD2gr
3HvrTteDb9tV50tZGiJWt6QuADsuZQBLFjJ87CutjCTu564vbWvucVDtW6zkdPZ+
bjbasxGi2BYq8d05rTSS3bheH5M1YvMT4EFDzgN8uQfWbSzYHG0xmQ25GkAuLFXD
ukNaexhaHI8G+MAYvCuYM9Fqhk4/GnBTsGSlU3/CP7T7VNSA/UtzDmWbKWnV4wD3
3MQ0WVbuCNU8wzrqdDKQRm594B/c0UbdYtTU7i8htEhbGYTUUTUaD00oWRNIhWwY
D3tCzzv4/AlVqbxo6/ZVUyfTBui4JAxZmrYwiEoPz6Vwet9fS+dhHqC/ZOKMEtfK
TgyUxEGQ5sCaQOiSggEKiQoGlyJrM1SkcIdMiwzxLivVBGaCyXUZpVLVhuE0TuCF
3L9avDqlNQbzTSLQALRXYjMvAsLUKV529Wz3Ln8rhZ8SuRKk+QJ4imGILUZlbyUM
GYUQHgu2o67emCRRhyW4F9hUkp11nzb6h/QkU82UUQ2ejOG6o8abCekDwMD3PynT
DmiKHdH9Yl4EeovliiYDlpp6fnOqoPzYj3ECkwmlEp3HG+ZRSbNU+AQzyIiUumaU
6Dc87T+Tul48yiD1z7X8M8FdKA2nzqRLCTxRyp4pb4F8xrRxOhogG5l9p6u7/g4d
UFllnYHafDlmEKGRM9lZQiY9A9DeTmuNgFQvwQtsgz0Vwev+K0hnHjHsK/SM2sIr
IaKX8OehI5takpSSw1VqOozogTYnRkg4fvsJ33OAH5VHSh8tWe/X7ozpEihgtVte
DZvvYuRc5OozR/VbUnmfGCYJcjVHJJ7ux/xjtgMFq4GhVRQIY03F3Qt4XofN3yEd
jbYql4saRDBh7HSKcO2BNYpn4v3r76NMKNwjgEOxtGTDgsj+VbEYg0xbS2Q9yQ38
DrQwI5+xZGUzM4GfOkxvFwE2KS5XlockTjh0oXCp3vgpwSge9spNbD/VO+utylif
ZsUlsYzCT7+/Nu0ZReH0+gDmnuNJlIL0iLAs4b5yL9x8jipGQkAK5uAmsGZ5P0bf
Wq449r1iR+udmUOlnzc2ky1OGjwgKw/yIR/kkpWpG9Pan1XshTD9f0Wph7/xUdC+
xFESWrog0qQ3tNmmChmExEP9dBSVWpYOj4d5vvj4EHeEOV8Xj7Oemq39hJSD7K6M
MQcSdrQeNrVuyZWJudtW9NQmVL5CO6f7MolD2kSKHdM+iBgjLnfSJwjdzpbNX8bV
uoT7j8XfVDcjeIHCD/k0NlO7DziQ6b0YsthNNi5LVxmpotCDHZGns4NPjhUm/wQu
MtPJ1IqsjCvSnoSuH7z6HH/l2w2PoKN32D8ogS+MDadOy6sy0z61PxeWGTYT4eGL
b7CEM+QE1eg7h6K5GhffIAALYKOTsfZynR7wURajxIsolAoWzyrIRP2+b7mXERE/
xHP8COPvUO73c0rnQ54+fOEmiggNTg4+1fHzvC0e3X0wpDpb1udr2KjeNMHTBZSV
YZU8B5K1SC0bV41zK240v3oDzxBnYjrdT4P/Gr7ytBDsog3BFQ6P7VNdxrbfYqfS
9I5/r0SyVBD1HVDc8trN6GOBelk9o47gpXL3DkUA/CJM5caUkr9Q+GrrBbhrGahN
t+VMIu58ZIJaHMUoq6Mnf0R1AWtaWkpgB8KeHY+7IY9QMmO+SyTQ6wB+kLHMpqn9
wwkajsjrzuiVTpdAVRoyagLu1XpKcxzdjems9n5NzkGXQfM2X/aFEQhMzNjLdok1
exQs4Z4voKefU6oeJjt67FWND57x2PVcNTbgUG2a4bKd5zS1h8wd7Tn+7Jhqch9p
ljVSnCSR2gdPrDzBjk2xrQpk1s+EVami8/qAlvvosJxazMRvceSIQOc6umtINOR1
S89qMV2xJAcHlj1VmJ3P8JmCvIZgiWoxnZhGZs0nWf2Z97NFuUy7Hlt/d5YmLPVL
WNa3NNRvQ9GQIo5rcSb4Nf5j2Ur3eEPofLTDOpWcqH6ca5X1i6WsEr9ke7wyYOsc
h5idABeTwjfEosrnxed32x8YWxSupw3yJkJnKxqckrvDJQWZIm//U5keLFk3Zd/5
URtYZTehwFMsXrqz+Mi4W60NEyZv+JFPZJlo+EMLe3wiZd/qah3hw8EU9skBymHD
sM67tQ2a8D0sINAiNv0YU59QDVh9bzqTtUZ+5re7Rl30lFjBl9+IlAL91i9/ly/I
UcViDgqtm1rele45gPsa1H+wTscK+nxJgnQZzsRm8TmYIncSpoQdiBI2LwUVokyg
aHE+9SvOKBqonE5wFABvobMzf9VsSWcl7NOFVsAb3KBmBEHLLuOpm2rCRF/IzMnO
I+NbONHnXi2Eclx181hLOa/Y54Vc5FDVsSD4OuA20nGsC828bHwmnDzhkH4PVX+8
PCaYHNmrHZqvFbhDf9BKksjZj3bzn/ZYmTRBmXBIs4UI9xRBV/UEIgdP6ngY+O93
vevIdzSm0eJRwxLxboO5Cdts29px5VZSins4VIJGmEaDPaqypefixA94c8uQY8Ky
zzPLv+Jel8yWTFktkrSnoasYR+9o0HUGkBMPKz1E0YVdlWw3QxcSnzPUnQc3jC2p
02d8E4Zl88slBKGt16yYTPNHCHXkH5XIn98XB9mf7os4R2hNSBP6y6oFDl7XQbMf
I9zPHVfa0hmuF2doxP8eOe075zY5TwoUNS2t+j6OcvLv6HqEmHrLnE+Lw8dTap6Q
BFo9nU5D4XIlhHlXEfZWJlrtA4+PjbTtC8/dSShKPESj5acZHG+Eh+VxQl00DixT
FCLXLlhGlvJgeJsIC65J12/ZRygnO06v6kPNA25V1X/kMaVCGk3gsKP+8ffMtQEi
JErhABPsnRHKf43+mBxwBdNHwqZgnggMArD1F1vzAUfDGn4+/8K0twmXFqsjpWPq
C1z+jVaJWtYviuhbsYkeWBlz1zqYbod7vxmMpazTGQ9ersx4xSQf5xaVhpGRH26c
t9+L0GpLrTgZDB39XW6AdUTDA283tAMf/j1EsbxiLRtwDtCotiYrw8ARJrW+7RKo
/7t9DP92pjJi2Cq0nJSX5DLHOTg30qthbEz9+71uHd2PkfysdSimMUfgouo+6muw
MH2oyr0vlkqceXOVIFAI03xdk2VFWhkdgXxCSGOJKSqvwZ1BJf6pnQ4XScJBGsB+
/bJxxoS3T0/ZtLnuiB+E2OE3XgAJXNTns4z5i+zLM115FkOpiwsa4sh4Hp5iV4cJ
0pXBk82Tkon0mXptHSDihe+IKG44cy9GohEx397uxS3PaIS6pioUINRH6yK7oxnL
O7NJyshlQAyvKnlNhW73rejF++bIV37JYGSBcsZl1LlQLnxiDaJzjDKMagry/EUp
Wc32s98+dodXH5DDfSa1JvUX0UUf8B//J4aqSk6yuBC5Nu3ofBzpnEqlNPYPz+is
FBf21ErWA+xKgnkFMv9ztzdo5ody1ts18xGxmNWl6zlbqwTuv7CqFE5zPkV+jaEq
ZdGIqS5SyJ2bAqU/fq0lPGjKRPt+S4oiPP7SeG5otPtfzGKpV5537iV4/y8Y70vj
K8rMMxLWocGgz67TeY9H+6DBGILPExqzN24YfiX4xd6gQqh43gUbSHcA/ywvzMPk
WI+IUtZY911u1oM9aO8dmc7YlAWaLDWpQWEM5ae9CuZKDfHlw11Mxq8hA/Cdo9t4
gn53HBbDcu2VSM8jpC0dPrd3OurUjJK6N4CR9Lr0hmvwNddL2qpn/1pHDAjKMtNH
40TmWJQLk++JVNVL2JHRHMuvTlc6ugziRGOUnLnHdjp9h9SuDd4RkP7ojw6cSGF+
pESFennv56gCXzTtK1i4xGASe9aRmWApTrXxUlShR/9rP1NNMTxN28e+L5bV5CNt
h4cHcVWz3CGRPi02AFCRQni7Hp6pABYxgp5l27HkPP0/fEmJmttxv5Kql0yMo5q4
odovgJcfnTVXBc43hI6eKjI8XBDldNlnn3mPnBPWhXKZgYM6M4fAYI4KNfYtAgqK
FshEq/0Tyu1cJdKBSa5YZdb9zwAfoPrY13AJJ8NRnoS/RsrCuLK72AMQ+GJmwx5d
F0chjl/ssaf9pWoWvuCWzaxfmyAUIXlxBUa3JXpGbyID6p+7IcjW3HDxp1EdrOuj
HrD7+2fhObIYfQA181mTTSBRoV/+VCXSWPy/kW82/OpHl8ElC2M+xs4qu6Jj1rhz
smUI49lRyKyR+cbfoiZqch46UyJliZ+/S0QmVOI2rKMeNr7PlWpD8qC6nf7XVGV+
CHca9TOkhzvRegC5DFgHOgqEJklRHJUsi0iPn6PG+RsI19f92YflR5Sru0tWMqiB
VpSToPo0iPKUtsm0c+VNWDwsSikFLjFSiMXYQDZuhZsIeozUt7aIzxg6P+GTFGME
x5dDe6jVEAEaszEnL8pvVA4f2Tt/lEU4iwlVGcTpkrYDAteaGGiSzeEeTU8FxLo7
74ojKBYn/bfVw+hPwkVy21t58LtQcv1LUbxIuo+BAeZ5XFBIQ21vSRmrSxFGsbO6
69yLSU3u8b0tVSyhw5usNTr865MarCD2DsMGsOaLNTCGdrY8Nbc0deG2E36riwql
Lz/dhd4vHc/QlmgDBWTeN+F3iMquhv1YXEz4D6SDkurxwlPCeZ0Sq1jUdKj8ShtW
ePjssOzNfIhc2A+PiDjU5oP/PYSgXVxXXfR8qp1jFBcx6wsm0qVuwcUocn63ndfJ
uBSbC41weSAKRUdHT8dxQ9YH9Ul5sV5CLl0SsjcR5ieBOhHhFKm2u2F23deDfVBs
jwd31o0K0HucPq9vlfhraJdR01dF5nKymE4eGy694yFSq9iXB/8XzssewKlXnK/t
rZyKLdUbGKk3cHuinjXZH6TTz3PzouuDqIiTgWwc+xq1CktFsvsZRgxaQuIhbM31
4i+5XxePMMmwbNoeTpGP6lz8AaDC/fcVeRmdh1GqD58nh1PfM/nsy05QEeHLLlpI
voBIHLew7E5xIZGrsmmWPmDIyIayMsDEi5mFjnHpsOjEPV9nG3cljeaxikIYWJME
dnFkmrKjmFTNR90RGDkPxIlfUUUpFrLKU3h1lgmDwqWc+8xcgRUXpr8nm5O+TjpA
hiJNGdy+vzjS9wD7ez+IRjXQA4XuNg8T80ZD/Tz64R7qq5QdeyYT6Ps21BYx/sRi
9UlY2nr0Gwh+0KEt0cSfAC9peBMkTIL0iiwo81hfs0Yu0FeIqkw/0uHv5z0gxPo6
YRw/K+clK/Geo/E10ITD8V8id6DassHUNh6rJNuP4AbZ3FCqL6zSXqu6ARVb/Unz
c9+PCt9uhbGn24PDS1jPJksyM4JBmXhyUBgnz8nEqLtENktDXKRFko/9VlLYITTg
Z/XYzMlm/7mezyveY9E3Qc4cdHhCUCp2hTw2K57XgfRNu2LJluKY3Qa7gJhcOkow
buzYJKi4lOs/YaDGZpU6O4HMZtCZZRa7NOXZZSNhUb2ObV89EhuQ1DJBlDusUH2l
jEwcjzm7xFwwNB8GKVccduu1Oj42X9hEqPK8AaqWOo0Dfnkg4pVax0BiabuMoVCO
YEoJNpyS4SZBS+qhIaySdB8wJfeGJ1jYxEbOe4f0CGcdOfLsHDmiOpa9A2nLxRWR
CViEvls/tw7bQGsI73IW3GVFJrFmY+g3XEWtAW8xL7aDz2lNz5T56c3QAc5Y96fy
nLVL3zwjb2yyvehMesVS+nHQeZEAUlpLDcTHZIwxkGC7rJ/Va66DaoiiHl9uwb6g
YAcmJ8KDYnvOKZS5vhWWSmCiuaNh1gMtxuudzCQrcrOXxgwQpNS4NygDHlaXKmlZ
Agzkg4e6AsgmmKzv+VCwEYpnQlBz9cZjQ33SMh8QT5ED7b7lQnopr4LNep1APipU
gkkXNEMmkQmKS14pQp6qmGt/+KmyhwB6pWosPxx85mO9KEK0sqZymfuxoGmAU26s
NxB1NiZOGSwt5UN0+zl6hqqSnA7bDvQ+yhcUhXS/F8Ly1J6IdYSRfRlmKvftKOxE
4TwDFA3CYYSx55LkcJ9VbGRnBBzQPN/pQOc/wARzfHdA5EAzz+OjPhm7fd4tdZXt
vz7dduuGJVfCQNIff70+y+r4W2BGE2rKOOhagUQTotS757s9BsRxTixCm/Feygfa
mL899QibTBG6ILrkzLABAe5NiJtkrfl4GGjTCGsTpjFPLS55eEBk18JSDtyTl0F/
F+i4+Jw40hZHj2xjnp1XBadWQop+DV6hlCVEY7K+fdN4Y8IV1ihN3UDrvO+YZbSJ
zBjoexPhIFEMxsaEwvDKbrkeOwrdXVqUBWQgilpMLnTQJZLYxqWCuXxBMafAAwGB
UuFumXVqr6jqOmcXCVZ/ydyjJihpd0Aw8ngCtLViQz4So+LZEMl956mfWsl8cvhP
z7aeLDOSwVRbVykpMKxTFJPiPZDKZr4euQ/PWpWQbjkSjHzZ3wjXw29Kdj42K6lb
hnD+1gx/ER9iq75YqBjCQE+n0894M2TVBpoHTWngOrTwGL/FTziBXh6slwjeClwd
F8WLxBoQhJix7Qr+SSLYj3AeltZyhDUtut5JansH3Pd1APmLYnG2Q709+CeBLRam
ZeeItXWBle4ASdg/zH5nxtxd9YTk4sBP3nA6dB4cRcQeRDGE+7SD844vUyxmQUwC
ovabR4OjWUmYncU2JTqzHSrHN7XW0e/eIiL834VCY1EYvIIx0GVIoNp1EPB5r8nR
JV30fS6tfmjBQKjuvbv3GRcOQ4r4MWU0TOIqAwmSdm9bHRj7cpRWRYtWV4KnohBA
dZ8ZPB1BXqSh1i1XS+anwOVsHOokU/ytmhC4ZwY6EvKtTM6j1Wmok6D5HAdgFJIR
fBbfhP3UDcS6oJjhlr2g8ENyUlpYxvwTATGl3Zh7FLp4OUebbilZ1PGBPiG8yYR7
JuzAMmEGpyCSCBgk3Yu7RP7+BIoHbMKIF718JsUeKDsBHXpE5xGTb7C7LXdPaSif
aTAlCbGohU3S5QCN8CSOC8rjVSbOEki1j0+AagLGeuETcg29yEx5YNIv3yv+z4TZ
5EqTSD1w/C8d0eSjOZMZHppxo4cMXmO84GqwVFu2xPVDjU5jn+biA7Kp5JWYmZBj
JS2inws0cxoAd0uinX05UfY1xJDQ4dbpHgOJVJ5lWha1iuRzqrvGjrLtvSwtblON
vt8/3pEut6OzUU4CHf5fdOlbqnK2o6GgqslZwEm5PvrZ7709VO3btg/VYAsPHTNy
62yJ4elXH8dIhIBHmm6kmUl0L/mobbFrkP/728orAlzlpd82G7ndT6c2OH4HDGZW
7k2S1Ar843zlLlJwg4LAn3FWivMv+2wwSyXMVKwJvgwb6IxFtw17nf7/1NI9wTgM
WzDxa6AD+y851/dMT5hEhsMmrtmPaSyyT1vqp32eIYJsSTra9hcYfav3Oh5T0BSV
XS95ibtpgLIUPpAhHYqPPDqsZsNOT/4BdU+sZ8ZxbPKaDcZ1BBOHpSqLU9w9RDaF
qmpK8Y6x3pCYJWsvcWVCQUG9t4elTk2agb5sCDWBw6piXQBMd5b8p+z98fEjwd7D
TW5j0SlH3mrvkLujLCNnbn65JQkBHBEKs64SEnFIQLYPrvdY5zCzffQqJnwCPVJO
2RcB5DuZFROIC40iWHlSbrEHJswya+WBBjxMUIsHVPdvHvjc6oUtDUWHnTLr16m/
z0FxGSsKHWjDuQe+A4XXXaNpkc7EJ5vUkO6hzKsU9jRXHhYgCtFnwAeRXcXtkLd/
C2diQDnODO0ffrXypw5liLdJh0No0aBFy8gMNkLEZPIKAUlo9Soxt3X6tWnwPLD2
/Xj0JL3V2zY8FdecE2J4yGvKDyt2MDkfxxW+oei4F3JuTrMmvCjN7VIQwiZ2TU0G
pKj9MIndUiuRMOwWIDK/BTvWFWsRsBfpg5fZjI0fTI07iBuTE4KF/Wu4vQGA7bLA
u1t4dgQJ5PkMbHYlW43XGaR0Y1l0UoLHSxiIfUzEVxBn6m9zhOBz3WFEFyeyr066
iaK9B3qfPEJ74xll2dgyqaAVg+Gv+pZnY9VlcyGxUu2vltdgBovXA1WYRJBI/UHn
Hy+g0D+H8MOjw9DmN7x3Y6Ee8nfZ4iRZ0IoqNL6ssC0ZilIV3PlVw2niaYqYxL+2
SGWLfSDiKw4sLFX0EddpROsqGmbFXCAVi+pp8+l+vY1OQNZfrPgMuTpvP4TnuC7/
3iKyuEdMW4pv/c6NbJQ7vV0lY1pXMHbwn+9jBT3FdAWR5vLDaxUvjMs3yDyfyAGK
qm8G770ev6YivMjZ6HQHcUp6eaz1zzDuSdxMxxWCumc3d/3hraGmwHwWNF7YbpbB
sTKI8EdSu/X+Viq8g68uyOvNGIgbGrtceCFrTO+lciHgQuaXicsCn2mGSs+F6pDN
7OpysAWwrr8J/bq5R9vPtTyU5VtUpgzJhrGpISZbTxLOxQwkSUv7R7TQss0QkutZ
TT1BL2F5acaA2Eu1Rx1MtG3Q7xUOrlaMD8Fwf9LspgbJR0qSbtJCUBQJ6EPfryv2
juMQ/Z8fvUw7kJCkSrya9ObOrhEinp5jncxV4aAVArlbadTU2Yno6WzIYcO8dN0y
xF0UDywrGU7EZ3mndP5SuKeJ82+SN5n2KsIx1/95Fqg/pmK3yAr8CLg6NrdGA00i
tG7/Dpd1h8nlunB4ASkoOGTB645sCWEsWj5VWBNvsiUqdmf/oYBznhaj4vOXr75u
kylZPnmhXbEDQbaNE8WoHSsq03f3edhgmMjn2zoJCG99R6XZCyU89e2Q3JH+QOu3
9TkVgFn2M4Fgd8Y4opCCY9WlsfV3MayxxiEXrJzDbg52Vzyb9ScY7RLJt2WHyGW7
/2pBwAdPf23MoWW3GLZ0JbfOD7qCaPeUV2TFRcYaFBk15i07ks/RnsHWTbyrPHiQ
QcF6P8j2PtAlXO4TQKp8PPQwR0Xofu6xGsMTSinl+swD0UFG0ZAPQ2wHpH8Q8wC9
33ClvUIhTsm7fqsas5DKn40C+EGCv1EIOQcC6eYYrchsUk6Pzmh5Tg4/rR7aJU3y
Vkxm3Djke1SQpq5N4ATFi98fDUicQLoq7ipbAtRk8QXAXeby/0wAzhEuU4eXn/wX
J8+wg2NBV8HKpjoFP6KqZMTVSEp/gdvUSOIuSIuwVNn2Hkki38WGkCSOK/OiZ7t/
qucJrSpHqEUp6xgplcZPXxztQZ4GW3AowjIurEbLcQ70wUvjdEtWEpbI6sBLzNZF
qaVjMJqhp3+hcKr0jLveogfVyQVlkLWizChhJB5Z1iglpTR6fbY/4cpxGXYym8Aa
JUTIzCS7wnDd3gnY+aVqO1mPBGRZDZbnpt/Jk1CsJRbLg+qXCz2lC54oLGmBHX1G
Uvtw6V/77I6BmoM3zzXxJVtvbmJFYfruBryjUjhmM4W9n7EpIQCUDfdBQZDo918t
vF8KUdJ8wOMIIUNsdx49oqa9EaglU75LebL71KEpHzhMK3BPqnt70g4WUW2HFyGl
xTS8B6MMa7TuOU3To2VMjFbBx6nO7oiT8JIdMpKk+9PGn+T6HFqNataHOWkqBxWa
A3PTTypT3m9e261bKkw08mps43lsuuFdcQvo19fhL0l/lgA0VHruqTgZrn1dw4k+
pfCETGdEi2PZg6gqOEt5G4TV0egh55a+bBhlMoiIM3GRV+ymdZKYqUx58A3uOloc
6VQmD52xdM7Q+Ah+XwJCV64G5L/RgWsvrJNyv49iFgLySv2OG/RqAmo4eoDOS5BW
T/sUby+cSBA6xPIzTUev3UTujl1b1Saix4wmoBBCxgchtalSCQQ35I0V7E9A9oD5
LJ6PEnqzgZmafX3g5jz+nsWcnPxdP5uS66lIbcc66j+taMotmQKxibtIlyP9oUMz
EHCVGph9IjDVOjMeR6WIqDO0xBbodelxs8ZnGfJbe0zvtmqXnmwVn54VKMdefZiH
yfQWReXlkXY2QtwrHVC5LerXxGIz7/PCLVq6Jv11NRWrf76SRoN50WrTDo59kHHM
Nx1KOPZih7grxlebZv0lCofaZv4aYqJc7iclGtivRt1URfKFUefnERXIIHw8Y6BQ
DJyQWnpTdvvdymLPLJyCgtJfPsf7WC9vHzjfdqDQHcrGnN2VTmnTIZWcXnk1PVGK
1yDjABQQ3aRhETZQQ2QpuwDpoBQrYjEQ+ZV7j/hieTeZ2+eo9UZcDQxVuCDefYu3
if2zRUt85Bzc9IVEzHREKV4XPvtCilise/MA6k7rAlqBgpRsWcS3NfEgjDQDd6Ia
rm46J8E9QDGgIC8nvAU9+S/JibJ+6iID/dss83Hzi9YlCF+eV97PkNfpykoXuO8c
AIfsUBmO0Ijptrv8JPy2BfE6uuHnVSz1DXU4zAx1pYNw/LtbJ6ioQZ7J7mY4ms5y
f0AjxIqu8CdNcbiLdGyZw71GSvYPxcEBc+lTydMWmDmLLzs5Xd5zSxXlEX/+uAyD
F02CwTbGF6Ff62Ff0NFYV6zqs96nYNPEPPBrmxT60h5/oYLXa4FJ3jpz+h2PPrFX
BhkbbGudI4bURl53OsHmzDwSE5pw2ijEkGPIXSTT60wFubdi0odhMk8DevNFzVRR
h/WlSWr+6W5VC8VdTDubORS7IXM9FdEvL7NYWmkC1zeuEsFg6/Bx5YBz6xOteYP7
WAAjknZIH+XYmVmbc7TwVRmV8BYmC/927JyFFn/e4AFI3uEvidX/M7otcsJsM9Ix
yV0xhrhM2LQ7tEtEVAW3LfItFUS2Z7Nir1G/x8x5sy7VhtgTztRh1HgttIYdQEgH
9T01QBZ1Zl1oUcRjuT9iW6SzS6x4xaUsjeIZCCqGKwNKGdiSIOO681ELl1fAxpSh
wfyX1PVMW0y4HPXNR25xZme69q8YQDxxCMQgPlaSB8cCLR7FwBLK7wAZOmzFacLp
D274uCmnH5PdnjtpCa31/ZXXOpSIpC4y/cx7s8gBBBVBJk7t++qno7ALErD3Bh+9
/OmbFEPTpjLZ31eLgfSTIzr6DSgjM0PMpvZnZrpuar4z06HNr6LCZyzVMw6fVRyy
jBItnJoC861vN6Uv8to7MwOI663ijK8DuHYsKYPzw1r22Up0tlHpFL3SBbHrioei
5lIdf1y4fshvrqUqwxIrYVILmTxLDpq8VfdL1UlV7YILZbJiVtTrWnIpiR3nPW+2
tjLVukK1tS+HoILtBjnkhT3cE432V/n8JJnJjR3+nOEELdRrv/NBPWRTFLC8pxu0
QkE+cjTEZfIJAdpQd7KPcmXvCcfEGnSizg1y+7UWfieyRQZWeWCyizPJTz1G6qH4
EhNIZ9m35lm/GaliSfzfKbRDSh32sQMekb+rf2umV0dy0sngv4Ea4S+h5cN0pEUe
COZOKzfc5qVcoPJJn5XN4YLL958CYMtFOtCSDFVm4TC9LDvZsZJGZdK7Kufn+1D9
wBmmbpGuN/NEbFvFktcWD6CpcgVFxonhyp+1Xr8bqjGyAbFGVjvc367CPKRzWEu0
00IC8teHShDBQSISCVF+lOS9Xk2ouf0j970okue/64huHV7u+wpmF/XGJ1H9ZJOB
KLgagr5QK6Y2jAtUf/lTRQY0uNS+8vyPF1ozaff2lIU8Suq+PC+6055d45E8xF/N
q+ZXzYXwX0ZzZvKlMoKtwmDAwnzSF/jASyLb4UlidjK8ZFINlDXPOCnDjm8yHoK2
vbW2ijLdqTnq8fQ0tNyYm9iH182AIkJtO1DmjWvIKS7bl5bQ9lw2ALAurMDh/2ff
o3MeNst/YBez1JJN18W+/tRmN1g/doDVt0ib9bU1wOQBSP7cvl5pX6ZpI4Giwk8j
uT5uRcmgZ+/jL5ZIS8TndTS0Se2zSs1olbtbHhBp8iJOBzXPMPHRK1oiG39YaAj0
XzgN88To+UMCB023JaSzbqu6ZyVFLUSo/duEQx3QwqCANjM/l9SVjkMWEngRBKD3
uSJuIiKQH0H0Krq4VmtTxOLCR8L04Zc86M3wNElvUCW0dq2iK8Y/ZjtCeTICthUz
3RojZGgu4T3/HUpFdHKq6TsUuMDH0TV3a+49bEg0ZStBLSQzGnsxdxG5lwHneRMC
3xB79Bs4UO6k0YqJia2bmtMEQPb3SjMehPWUL8Wn3u0phsxTjqabWPWVm+g9VDuV
NyyZviJVuuF7ux2MXJj39XV9eFnKiTu621BTvLerNtvm2yXmh7pwzC3DrM/s2nNF
5yTMQwpb8M+ISDAhB9JDFsQ9tQMpJWpK/LXpGe8f3lem8vNh8o5W2soCZz7J0kv3
2gyvSfxclongEdaYFs08VZanuDLCalWiyf/DKjRjhu4sM8UcWRZL+KBx2LmJqXqC
PTV+tqn6J0Uc4x6N8Gv++TN+xm8+OfjVamedSoet+5cmfWMYJp8vUB+HMImYxiPN
YFRcNO3L6xifo02y4KmbwdwBQTPdEqhTaVIzNxvV4rI0exiLwIr1gwip3J5geL5t
IovMJxutoRUCAODuciGb0lqzbWa3bpl5RvJc/ZWZKq5zx2TlyR4YoruWyRpwG1Rp
INdAiBlnt52hhaYlUM1uVPlTMJMq1+15aQaB1IGhgcWBM2mFVBGL0x2w3kNK3nxu
3/zJ4/MOejtayUK7c8rZRySd/ULmUeQ3CElFjFlDy9MbZDDtwkAGKnVUlJSigJHk
SwoX6u6FooQqwozSjkJAwjqZamedsrbaCuyPt9mAUCajHKzQHK3msti4PGkJ16Rz
uTD7iGT8BcgbU3OoeoOc1L0a3SyJvxnrDwUciKcR5t9bTPIAS+481qMhi7JSaT72
rN3DSeMjkc6lZbbKg4RuC5LCTSZjM8bO+BBi10MDfD3vWaq2haWW/Vicy54rGjYI
bG1XhvtFOwK7FM0U7C5Ki+ap4JUr/GgkL3dNaD10n1Qd6dW/oP7ggd63CM4eGlvh
N43+cH1YL60K/EfWtJfXMwK3SN9D1o6txenSyZVWyUC1zp6n2CRbQa7IZWfno7th
r4N70OUXDfp6ZExgnyTQ/Kn18HKCPRT0tR+ZqA3jHw1y9R8OUuLCcRVWZvZkWczW
z2noFgSppTrZfqt94y1t9ZKPWgbvka2XD3gLV0wog5tKt1pJ0xaotfpn+rGgGI/y
1ug3Ri6OEK31Sotbs4B7fveX7D2ICfF6BKT719/zOUnwnBaT7Q6wiQWOWkeRMZjY
AD4qNsmMaBulgJm3mZ0NGrkxQS2V6kYD941nGySqj1rJyiDxMip3j1MDgUB/oAcn
NnqkZufifi6n7arRTJBxMcpHZHIf12Br9rZM+LZ8j8R6pMf4T7QC4+iRE/035pkw
TY45GPe34VUmhmxZNWSXbql6Yv7n3YBbTslsgMmqz2rWvj27hOE272DlkQhADnIJ
TVeaRZkWtaHODD+v5TcAp2rNGD3VUcA57XJZ+3c+0pz7bsuH8+uzrUChVhxF3Y9Q
pH+Ct2ZeRh0Dv8pY/KkbCmNRfRyrmpK3da/V0t8c+EoFiiLd48WFjmTlxenMrkGW
kB/uTkHMwHdvbN0rJDdLF1vctLtBNjHjRLKLEgcJgIesa9CbbtcjrUVW86Bo1Kq+
A6/cNK48bu53BXvwPfX1c6l7Jr9xx3aKAgV3ad91uln1+u35jQgnm7BgDhyCXWGn
/mO8nbHlCgVRVmbjbvq99yprub6TQZDmJF7tSO/zAFhY5iCscTaOyAE9i/jKhM3I
29T/ri2aRI5NzOso08HqzU2nvtqPY/bg7Fg3dG9DlFFcON++uJaxAnajXgHR96LX
WEOEEZ2CVr7JY48sCinT5vXs4iIyMLuoz+3z/j+91137mqccI47UtidGL/Oe6gqZ
eP7Q1XYadrA4o6xc1m64VzW64pLgWzKIv0t/yyu9Nt9sj+BCfHuHkGxjdPoP+TsP
ceWkUV5IeXfUJYDSjYgWMBtWT3YWl4+gqWc6taaUcHfnzfttxmyW4+SsEyOV2sTy
pE3UBorF+2yNRubftxSRBS+aQs7PnhrxJvB1Z/rqSpXHxrokzkVCrVe+LY3Kz0aJ
ynyOCQa2cxPxWNvFH/lWPFOeTBIfWPv9ODLvPxw+Zo4zDI76VoEuyPc0I6GqDJJU
FBcSsDZ2VuLY/+tuLgjmenw1VBTjTaI4XWnZMi5ZAcNa/JDTRPaaKIzlnVrvme6i
c5bmBnNYqDb3kJfkR7XQEMXu2HlOsXFnEgfwZ52cBkB0xDbsRmonC1Cp59L01C69
hwgSL/vLEN+XuV/54XQioUdWNtrjRDNh+mo3uwBGEUvxoNXqJIZr+rz2/YXSDcqm
cTG4FFLjgcCWM5G8cN1le+nIxztoMw0NoDR+OJgjH68lzQupIi5Flb3WdUSW69O7
xi9PlM6VeuY/lzNdzAaJW95Lnt7FmRVZRRdzeyGO1VW2xEwZZmdfRfwq2p6GeRmF
nfE296ean4P6Urp1ux/g0WcWmuraZObtHpd90yiD5nuXfj/I8n6FUwzlnEXnKjmt
O5dDzIxeIPw1V5ZnsYdDnYYGemoWQZEDVGtAauPteFaIPue//IntxhVbMVKuLZ7u
2/4PKADPjtN4xobDuDudg08W0PbmXpjJ9fWlZ9qHZQ6yLeWeEBlz+E9zJyJuNxhb
0cjXOdSOfXSkVcq1ZVwK5/Id1GKcJz438llDzOKNGuX8kJfZEg1YqL28x1jblRP3
djgVCTj6UVW6jE5CbZMlqKKacQs/7y5r2V12hUzM/ggLOX70XBHw5CLZnskys/tV
bhVEeBBK6HEJgtIii1iDMjmx3l1Y7nGEb2rf7f6jbPgpWN05393kIDagRcEiSWO6
8yJEG9teQVUoPSknvw+QIc7/8aLfgr5mNIREIagFbvJZe/kaVhivFcAM2A32wEe3
GyBDpLiq2ZZXMyrAr89d97+7BJdWALBUFoZkGWeZfoeNGtrtLm70GYYVXpE6kqnp
hBtTLQCQqJlMu1c11pnlbqOhF31Jt0PvchAw4Q/Lf6L/gh9czRzRFDPUiqS1kawA
oR7RQF9MPvWIe4gltL30w0iCxf8ieiMjVW/42uhwXJlO4uO4c/RVXOgYUgQ/OI+A
NRNSqBNf4kYMOryjxzFZl5+EFhT7RL1hbgNThtnq9z9FaocCcUq4WOsaYt8MsDwH
6ncM/fdUyiDYAlFs9PWr2+yn3su31PndUapWQhcskVGCYy4vp5+37VXs3A7yMMMg
LqPA0T+GAwaKBxcvVt+9ae/AKTxh/NaaEyPbi6GVIj+Vt4eU9OqvGEBoSsRaVLMN
rd4/DCE0LgbWmLCjiruvmcQTvLg5N5AVTa3ZXNMUcCyq8T+H+nExJ1f/HZEXfONb
k/jtqVTIcZHatDS8BwSu8NtneWovcBLiNFxVyMLgt9V+C/dLLI/ORw0tBR85ca9W
zA5Mzt788eYphHBgLxdL3MEZsgGZz4PJ/YWON7JW8T7NU+k63VK0J0GBaR9hJy38
bZuRKV7/WM3dClC9fT05CFlEuoiDBXOL/UOUxlSAqBNxEC5wcRn9yVs5OCL9MVoW
MFU/GQ+qFAD63s7ssbc3OhIdCjjIQtaq7XUUCFYJhA5RwqeIZr0O73tkuwAA+hVO
4OkrKhxL1vo8vUV/4Hx5GV5/1CH0DVVliwpQXCFz0A1ItNqqaV701jqDYCJcVmOo
TOk9+45htBvZ+0QjZyu6TxozWktGRIQJyZrjkDDgRbgw0ZPlU9h5Wa3q+e23cgvi
U4G+/JyOxx6BkXKjgSory55BVc2ssAIWtFpFh6+FH/B6FFVe36yIzf6E3ARUZyAh
3ho/DnJx4Z6v77mWYgpxQERZ00PQPzVSfPQW3P2M4OG8new8s6Hj+HpmUJ57axTC
21rRTLk85Wv6TJG+/kGu0fr6OoulkUX9pPa1cwvBl16uZOaUDeo2erNLTSnpCUxJ
OxWGudna3szVZF9bAwA8P0ogmozrQrm68TDNeB9A7k6cu6meRiHloLLQvclchZTn
yaMIw6weq0oZ+pdL5yKt9G11Z1sl798Vk/Yam/AOfYnC/C/z7umlioEU6tRPQO4A
Ff4PbjDu08irslDHJPbAmELwByVYvDZ/mdgplNVfXFiSj4F+SHkfQeUAqd+beBOs
LpQM/s2VG6xKCHDwNtmLqgFz42lv+c+pK0KfQZNcr6MoX23mBNGyca6QvbCC0pGd
0L/4BtJrkrXek4yowTL9VBB/URwh/6ggKsxK3zNVtofHcYZSdSoFsqnW04+VW7+J
+xAcZh5HfdPJtGBKXyhQJNuV2XC/uQprv8TpdYULSRAPyP4gDIiCUEQz/XgEbBpl
PXzFo9DPW7kmJQgNjoYET8GPdAsoNLC5xxTQazthPvy60rjPonw7CH5i3039BlEN
vcKX/mSgOjw8VT5tuWM+LRqI7svDL+f7889KiyTgIlnPwaSEtl8juvmhds+slIy9
FRRw0V2xeSozOnIUPMablKkqagDYw3fAbmM9GmlSYoF5wB+tXbESfxVNgrhFDFEF
/Ea1cAzueRNM8y9SUgDQwjkspXmV252sMpn/Buxn4wXnbQxAyQkkqjOvQwJ43cEH
Z5igVefzr7z9Qd7ElwD7sBU9O+DcNiOMHZx4icVeACSNqOE9xkwJgrMeGTNa75Yt
vHPMQS8nnt6Y/35QyX60GQf1yXNWNEmlu6yuqhFVUQUouHYYni8YqSsUC9FlgvCy
CQKVzNEqcf98wKhI8rL4EYTvfvQfV+ynWm9yqJybeBV+aRMhoVXIotX/aK4Hsi0x
HcnN03STa0e6QTOz7DutZZ8s3bhicUq5OkgmQ/FQ2+mYFvKXe7PRuelAmbxnvyvy
BGB0wBRsjP/3P7Zg5S+ikYumTlnJKa2lGLtce0/kaJwm69nEoY29sjN2jsyKNVIb
iAfS/PLHw616LiaQG47BtDk2kaXHqHxBonP9VO9621mPtyClb0SEZKBPBzVC4jNI
of2Ip3Dn0LVGwlwFmN/B/NTv7PeknU4HkhdEgW7GBeoWjKQBF0pitsfFZqPtY5Kn
kpHwqxz/tfEusXgOIvFnDXMbWyH4ZN1ZdmMsdNBSrwXIhHLrH1r7h8tX4R9NYoVm
1YrKAezRVoLbW/iI8MOVUfDJdD2nudNITRzK4tSeSf6plJd5oWjhgNrhz9uGYk+C
dUj9EWyb3oYa+s72k5MtQtwlsRv43jCnJ31JRkWbZsI7wn95oASJPbnava4D3mF7
dHHSg/FdAWjjP3f4TrryT1DzHtZPrEywRWgGGCoGk1poZyn9zjvOhr5Kqjh2kY7V
MkMiN6kpHQrzuUeTICM8W83gTrzX3tNa3DfpJABVHHYaGcOy4zopAnYXInVkmQKd
JF0wThvKJ2hwfNM8J3ewDDFJD8Njhm56nCXx77M2ncsbH5LYCy2WXE32mY8g+MPO
q6QOlBeENcJr/Vd1Vc7OrBwmHABVUyDdgZ1F/wad4krVXrPtkIfZM5IJpIqxt2Wr
WzfD8aJUsUpekvx3w1TCMBGxOiCaFifmrfOkGHrV2AeVdl0pAGf1RBU4rorg5aUn
kh5LJ3ABCoDKenWEg6g5u0+sqQ+XnKpb3A7/volX6JlzGZV77S1XvBS9ct6MENLV
OhSZ2n9L4eh7sVSEFRy7pY9JReK0d55q56ezsCazBzdQvxJ82Ccc93GNxyQ4oceQ
cGmpn8fSwnk9VVGyqUGcScZs/Zr5Vvs9kHuNpwq1r78vQjOMzdpALm1miJjsJLwp
qcA5Vwez746KyqCP94t8CQgpsWaDD1iSPKbPfZzSqS7IdSj+mMCLJrY7IjeLD42L
k7XXK3JKlYLJxf47SGYEDn3grEmIVek+4Ii0QIO51AvTude7HYUADaB/CkamrNFb
3yHHV9avnj7Cat3ywpcrEQNm5qFIawQ1ywjFTqhVicQ4wbcT9WG5xT1giA8hI8UJ
4NiFclFyZA2LXUFGfRunJzQciyq1Q+43SLTWY5RZPJw7Ag8U54gChWndGGHFPZeU
dBEu7hw9PH/ipqr7MdpSNDqy7bWVpGWBhFWh9Bfgb6m39zwmRdfdgUqv8PZIB5nV
o2dGf8pLNP4NyKIO9iCs28YvApgkiJWP0e+w/PnBvs4fj7YdiwTSDt21zxQOT0Ox
n0Z9mZ6TM1qlTlkyJc0sM0+U6j8gVU0NGNZGfWlqZaRLNVQ4AU6a8XhPnsuPrG4f
E79hOTaoWYdqD6dh7d0lBfd41zcg7NO7oJeDLBtfhS3NPdk2GJwHgZeNwlCLY4ho
Z+nogj0wkQ73ojXcnd0HnPnY0i0VK+iwY1Lta2R9d+xZZAj+8XFfsqlxweO8wUnu
n4HgMr6aGew9mzyQ9f6I3paHxlrZmVGW4m/aWySPi9m/JIKQfuYzCMYebBpQ/3Iy
DtbP3NTiKSwlw1KAfnS9ZsfX8/U8IMQniw1NysI3uy0DAF9/XoKEoUgE6b4CbJvO
iuQ5SMkS0JqF+vOtyGwno2A/sr7B4GD4yfM0A0HaOqliVD/gTlrEQRFnBv9baUaS
xVfjqwEJM5wcVQLg45IMZ4fEKXH1cTKF5xS6PRRbEPIeJKfUPriujzXnSlFt06uC
wDZPc+yn7IG6+ltYNwB+3MOFOg2t1KKjAwFwlFT14oc3PlF+CdOABpAhhvJEgI0+
CtMXcm+y9bKHrNlYwncL9QV6oTAPlbz9t0oAK75fyM0iEEqQDGU7rRQIfJk6RcHg
s1BVwUBcfqFyRWOSg16wQZ6TSXTWW6crDUXozOfyjbhjSnK1U/t9AGglgl1hpvEd
cLAu2IZhzC3cIJrDookSBbqNv9WnYe3dnqbGiGFwMF/mdm/10buE7c+VuWU9HLAN
zqEvcMBuzoD5nraC0lUVjCq8U5DX5ByRk9uVN17iQT72LgIBQpJw0NGa8okefRhX
+6crGfgwW2HuIpbX+5WJj15sWlWmKw7t8SkWRdmv+m+F8Rgj2TgMFfY5GO6a90Ao
Om2tQF94BB84CQ83MrqYDH2461oYt3HbnhAjX12fVkCvU+TmYMJpM+3LCE4WsLUL
VRclIkUNFyU7PoRJouGUfisC1wv0+g4xpzS6Gzwy48aLnBMEU3XAW/+NAO5MmbIx
8MlA7u6rfRv2WeRo/5GfkClvpnpCWZ+zlCSGej6gDe2XlguTJIO1JdjqL5yGtQPR
GNUX2WEBJdPSp/UrtY80DpmqpXBt4kq4MrRS5rkNaFgVRWqLs7zoDfueBHCGFzyz
iS92xIhIusjICme2j557Fsybhu6H/U0Cgv9Bn1h+5xgG+1EjQ1QNILN/8xctZZou
9PD49cxgD35DuTiGKjFwn3+CybC4JR4hf4eul2nIWNIyVDyEMCyLfAoxp8B25AW/
UbuIGDSwltMOp/89D/pguZ3DTBECnewg0C70dqLY5q5wgSokYuUdiQy75WmFIDu0
89q9KYAgoP5RS2r7uUpo2iuaF3hjc7vHTfWPOACMMD+OGbapYuBEnQRHN3M6xFLo
KUonkOYGGYaefCnI2urMWiL4BvemnxpczqmcQCtaXpX4stJs5BKTOdy6oZ/G6YPO
gtLkpDg07M0EvMoooaLD3/jap4ESwl0nYDCZuzxowlMW21aWH0JHWgMMASDVLxYu
EOQ2Q+gmz7B0171M6/yEPKWgJLp3+qSyzr5cTWsBPoNVEnbOEzShJeKrIUoKfS84
0YZiP1sa+PJAyrvcTdapbJLRfyKNY42nGlMHtEkS+m06TcjizAS6bDd6F7wJj+s3
4FMoEyr2of6uYI7x2t9nwmd/anex6BU/siLTJDD2zKhW9TCJfhSl2wsixPpXOJOe
HVVyju+cC6bPKdtDWKM/Wi1EAaPopIc0axnTsz5wFlKmnChhXAcr6eHbvdo5/WSI
QXP30PKk54LcZdEwyP+ZbR+Jg3gZpsylxfOHUsLLKvF2hvWooLQ/EL3/FCSo19Cm
Mce47ukaGk+h6wHER3WPj51CNTEd7rxr/5lnFrnUC2/KGclsrSncUf1jgITVcRqt
j7cZRqHrAlx5pfrB2eyKsqeLvI6aFgG89jYy1FNiYn8kVfwdfwZseqFE3wqIwTwr
qlj7J/l46cmnxeJhMW7KqhifYi6+lTZbgbrbY2xibuAz/NcqFCMXVAU4nG6kZsE4
n70iFjofuz6NH6SbezJE0jkFNkPTpCMOXmWsoD1G+t4rpKJZxzfqbr02IqpO6H/K
XzfGTRoyOoMvYU5x8vdRiKjNnHHguB09x7Ic8rMwcfIyoCw6/JJAlWOVrRW/ycVB
cK9SjsYnZtj7jq6BCklJpFvsyLNjB5Eneinl6lh5YD1XIeqcmOCLbVWq2r4mFama
PAL0lwlFxW29AhUPvv+EzQSqcaGPfDeM1/HIxKRbvDXLV6J7yV+55FfsFkADMygJ
a3cNJT4OfFnzv7tKUVmo0F+DL6aEUTvaqHuhFHyoDar37IJLK6GcWIWDuSiasGYP
6G+iToElTwQUWZUSdHpyyFGh45zxbOWylV7ovqa8C3gTfG0UX6Ns4OsMCfo3hv6Q
/S9zICt330WrtN8/YhMpV9ZUBCxvA+pJtssJNxP6oWCHalsLmB2deejGoex7WCma
WQQxbnpR84/k/kTWt16EL3icqWDCiTPLgjAK5NYgcESaAmlaA2IOhyoB2+C+jEEd
GOgKdXFtAnTzAnAFftmO5kNwlS7D1M606M7KOjeNc5xDV8JClWSW1XOXY/biUrkb
uYepIufKgDwoq6KZWsyanm3fpZ3c9mbMDKclTQtCnvYCfXFlxWqUipmSyaNGDtWs
yhpyEaC253zUjcwBMbC2EeiL+AlJ1gspXU5NLwEXmyh/dbZu8WzzObTQ6iTt6rky
LaCFcMhFg4BOyhG4eA5G1XryUi8UFVxrsFCR8Cd+QD4qdP9Jp1Ltnxz3Z/ZqAxj5
29eEEAZvLnJ+XutqAbvkwSj+2iZihTY07hdwiWwG6AX4TJxeJ3UDUThNKQq3lB8A
D5O8vL1TIZaYXCRPGe29hmM2ivyEBaRLy/BFUsiKsSFbzZVK1Ek4mxLOvdMNw06u
pT1iwKHf/lMl/TxmMyhztrE1zQUsIgrSTFFnFtajyWBakIEjB2oC84KMJee5niTf
1nrv2pe2D86sTDjge0peDagqYazWLUUy1T8jKdEje3r5cHfaoqfEGiLkmZHt9AZi
9n/Bs9UX8AtWQ/eCWbqieFW2yQwaR+jjFmqxPcLhKDEB4HtjhqfVfR1Yl4JQ0A/m
8WK1q4bJdCRNT57c7XpD1PHdIPjm6dqr/9UpSdQd67iOn/shBMBsdsz7y7/X19wT
AP5NSGgWS3297cMp2pOtfqij4suKj7k403eWv99WiGfw+GQBj0XxUxibgKJ8j56y
Q2L1R9wvyqCzHolDppuIS+wJ/vsoSRe6WC6VMwj3d+hMSkQmasu5vd+wy3H3jdKb
mNoMD/uAFH2Nm///bwJ78rYya2KFQ/fsfjHbLCIiGz7LoGtbOer3xac2X+iM8gaI
oQHYhtZxksOYgoWn1E/2Yxl0qXIFQdOknmlHruqvQIBgF74RrGyAWEqV/eqsxeUt
CkVdrOmI4f5JQv1MbhUqXrsKqFqM7k3omtwGjWs73/WD2JAp9FxNm5ZbVfkaMOKN
q0C0Jw9vWwyoLQBUIZfPljOsiEhll/8E/HrqoSsIDlF3ildrSu2aAynLuVayoBw2
RxBNWeJnp9NRowx7dPXvsdXcj8fbD0m4Ce5qnc7FmmPsBy67nahdqg2OvtTvlLS0
jFkNSObdGDokm584mWfT0YQzW7SJ5Kn+HJ9uLNKxfcT9o0rc778iyGmnc8wmVbVn
3YxVJXTtcaLshMnxx10HkH0qB0OPNWU9chTVgeD2WOzd7y6aGr0lkHV5IWxZAk4u
tgEk/rdB/Fm8XzCWc+hGDAqdSNpaNhgsuzl0EQIAy0TGyxBeL3roCyLukLadLJmw
nWtimScHT+0CZGqUZ/yH1w/Txi0DIEFyV+Y/4vBTyjjqG4n/NW2ZC8eKPiLCUcEo
mlCg3kGJ91dUO8Ldjy4dXwlP/w/JOhVhGR0MiJXN3oIn9ij/p5Y4pMWeIfh1gK6N
7d2SfHjmgRBLdyH2croPe8+alzut1TJJ1S13bebZi/qWTwI/f9+6evIU+5uMp7jO
aTe8r5xbpNG+YGePTrZdm2s2UTlI482+6lSNyNo3lqjTShgCWhWeRdqQRBxiEnIB
322GlNZSE/3lgXCB25cGqM/1N3DSpcbOBb1COoTG41YFlQzFKnvXhUW0YfFwJO16
/EBww/HwgBbC0CalcA4KqVlDSblfaD3dcajSMqtvqb0Gmm28hdjhzgGfLQ45sNrP
uGeWcrvjJCospYCAwCiR/rs4v5PgRSL2z1AEV5tJ+3O5r0+dkpDaJDPtJfTAvPjH
TxMDrPkiIpf9o+MT4twR6s0aySepjXXj2TpRWTptsPPMSSOPRedohZQWn/ghNt3I
0gfJMXbXAvyfKLq6spwYihB+zHjYpnsh3YcISz4Vv+noee1sxPjoD/L0F+7hs0Lr
EfK813+LaDuNJpGY7tFfLO0uYvK+t901svyt/aHlOcEcwF8iizchKEAmp/9PEZ8K
nPsNfyYuEWyT/odFzSo9uk4e7pkTLUuP7/jX/pRgVw/G2NXi7phfizEEvVsDG4Ta
SvoEcnhGySWC37mIwfbuRabB11II6drqsdbhrGekXw8V+pE3W0MEGpD422a3meRu
QuIHLm1C+SgJxcRruNPSiBcplJo01+9Oa5K8RP6HvNx6rwhi/3rVdaiXcRryoHQ9
q2+JU12K4ATutVqskdhJs8hitG4s969uWl+MjZiDOuStiDzLqKjfxR86XzZJ8Scc
vzC0SrH9bnS1rLViRFa/jDCaUAokwOcjditbOGrGVrt/qZczy05PBEnwWep37GN2
GH28GoagB6TIjKolWza4HbYFrlM0xzKP7I0/qssSkVXpA/zBFlZV3qdGAZjFbShQ
qQO4nHEFO/eHO7uppSCiiN7/xDiKNMoPYzjtAMqrAA9K7vV8ODp0nZPVhGgm55ck
in4NOl/9oocWmJ0jkz+Eg2eQGQfU//fJ5zX3unaRCStw6zFiPxUimTXFBVJP0ghc
KypfwKo/8lTi9ySVKEURJebeE7nssRgxRZqy10M3y3CrU2Kuj6I+ERB9qJbM11pw
bGxh45cksh9Z/SzojZu5ZW8RpZKC+Pi9oIV/74ZYMUOomgo97iy5Q5858eFFFmYm
ksrPsW5hC1RCMlYhmO88VwLgqfCFsWgI8uL175hTZASXZvoOAecKVEz7CUy+0v0I
s2YdRUhnx5h2dPzSKI1neTZpmokQ0cTiK1FeXCs3aPw97HB2tN3OLemIK+VffNUF
mbSeFOUVqZLQp9BKmkN3AOp7/WsD9kiUsFeltlMDn2gi6mCsel4XkRbi7kSXvnY1
jBTKKqTPUwrrfmiIqfCabjTYiAt4+ndV46TgRZv/NaBIRb8Z7kjJpfVh0/Z1sbfh
Eo4v2ZKoPQhABcx7EnZqh0Kp1u8bxa+45dcffEvrESwSeLhk8G4B2YzqtFS13Cl/
LIVW44F/0sQjdRpL2wXGW/dPhLAszKFhBIqcFOABf9FxboURFqAYSmWnooaD66M3
+7AD924zp1b6zZU6Do0LZxAdDIvSXakKSlbOSpwxAeFFldcvC4if9J5qZIhlONEl
P1IggxZp858Y0TR2OHAgUmNrazsbDtBnhkcNrTGBpWHrEQA2PmUrRgEjEEYxcksq
x11yyAVxpy7rxKkHDenYI3GheKeGoWQH7NpeK7hCUG4zyO0ZTh5tZZmCB0Q+4f6i
YMrIAXUiDGp1svchsGcuJeFcu3BFc61bfvWcAgUMbrXrzKbmimiePMBeATvoY0DK
5+vIazPiHdXCOewRCFRXkcy2lb8Jezc8XDgARU/YV+eenRwUN2FuN+XTtV5wl9pn
ad651JeMrC+8s0WjgWBjGi4phl7SdBllZjyWT7flc2jQ6CxI5cHDo5f+jJO1jBuP
Kpd96voMDscQ7ut3zIz4TRuItKHa/AAVlaS80reDwD2nkl+2VIrq2r6xVGH/IVin
K/R3pwpSKtpfxJIPm8TKk6wqGrl8zBakJ+k/CdKd0ZZkEfUm7DTRRLehL5ViZ4n7
FPtbTNFRVnI7E352ogHaPgJ9g/o67DSUeM3P6jZ5hPUo8Zl9rKzqz5f1XLmE6uJT
DwHB+4DN+Zajng6D0X7pV6W/LgsmXD+IcRmE8TOp214InWdugAMYRaEkbEoendcn
rLrbBmy+R8X6PWB1kDti8YTRr1Nh1bLF7dGOrYdle9HjP6LlB7ed38qSOpijYKVK
B4LwTkaSPehUFJ/21Jsh7n/1bZcaRavBr0EpRxpDTAcpjIsDZ1WMYi2xtgHbelEV
UsdIoNwhJUYcLP7nYf0pXZRncOKuUOFpyn9+nlCNDz+gQSQx2qx/EhJFfcLR6un7
IuTrNbtzqICh7EsI69iphE70JTRj83GfE0xoC4EqPmvpnwWrdErR1enDL5gqAmN1
zkg8RXoWeWvnherOooX4O6rtOs0hae9rgqZPL+LKHVQf+HhYpO6wad/GDanW7ecD
qviJ5cVv/vUUx8dOtP3JtvJxKzueb5D99xjimjVjaTqZfXa//J8Euw7V/eGOWN92
Ryrz3XMdHsvIUOG09qxYMZxavq56r9hein8QIO24ru9NSh30WkNF2sWQhTn+st21
dc+OqqN39UtypVVZql8KFv+mruOpqT9IVsDUV7MhnNiUowgsvjmmpia5IdsOQDol
hWVyszWvkgYHjSpdUbK7g/o9X4rzba4Qy1Ku4CxdH33/RRI0tfzkRJxTeceHXnjg
CF4k41Q7pLreQkRv9sV8PO8S9aIFbpUKDExElLuW9IuEXjeDTvY995CTXkwUiz4t
+Wig1ki9nxUMUSD6EupdU/bnJBX34zW7PPIBwNevxvAzURJrlDs7tNhZJJJwEidR
EfBSpvj2E5i5lKSG0EJPHTYb/2nMBWdSIMrYEdqAJv3ZkbSx1Swnu7RBsTMWX6DQ
h/LWddc5lK5ED2T30dV0xUIWHq0vP3cYf1gFBYbSjL4/fwr1oWL4S9P4H5NPl82G
Ec/IHdE3dT1JNWo8RvhaatZU2h7/4aJMc/27ERw0FfPFEX1sRah/USCqB5Q83o2P
3q56xB48E1lmpA2xFAjkpUCldcLq+RYM0XAX3JXGSfcd41Yr0E7cicIjXX45yyNi
PMwiDdwKn6t9SJ+tEIwF+NpwGm9ERuP+HiFal+moZbnlsAJ4lc4mU7w3k/+z4Mma
gjjbwoZd0peHWH8zIhTxDG3HEeXGT1vAIIrL0nnJc5kU0bR7LMuK8Di6LW7CbMVR
SmtOsPf6SK6pzUME73UayWUpyjNRT6Jp1973+6I3EPY39IEkSXSdO2oALq6BZoqx
kMPU1SUY5hNfWzIo3sj9P75Go/peB92nK9dr5KN1QuHWXTDajf7JNBHUb9RgPZK8
fmbuKWoxJ3zSVxeONeDcBCrekn1WEq174f/6MveM7d4TahxZ3NFctw0+/fIfhth+
9VlhFPk0kh7S2VPyV3Q0Y6AoR7oVx4mpER8/0EPBKir73nf2HhJF08iSChGHsLqt
Whz/ypdwjPTIpSm2kLbThttSF2W5ubKJ0EwDvJddVgKC7SWuZq4lYDONtS8nS9b/
+Zma2BI6Z3TpTzGDx911cFXZ0eXs9AZPJDnZgMaPV2eykDHYSy9Yz1kM4r0Yb0cK
XWYcoujo0DhadLNM7wcFJjp1yyLwh9EJaFzbbsQi9ufAKYT940Uy3NVVCz8CEbkX
a3jUC0xXzR9vc1dJ7Yup6/4H6ofvkbyT1ouAJnmpSK9fGnrnB5KopZaLaYDTSpce
iBrzy22dd0jNu+YNZPN0cbY+GmSEvbkmzqVM+s3CLA/rZvYCISBM1twu7wdDZYso
Cp6UBUAfZhYJIY+ruqXIEPLhvDmfi8FtVTBsA2g/zp1316euDCNV/WQwkkQex5es
IIwfrVWEK2I4a9PPMO1lZ/UlZ9hn7k8HuLGqEDDBm10GCNXK3+JOJK8ZGIYYsBBm
nDarVkkj0TmHJFwwKqpKS5J3WcQCL5kvLAXDotG4DwBkp1c2pM9CIVLuqVPjADvd
zKADIsP6i2ZFUMgxpxVr9A/oeGd980lbZaeHwf9JDIzpz1ubIlKiY5zF1EzJpVo/
fmdWunOWGI95Sj7kiXwvWcINI1fo3PzwiM8CgQWrCkuyoj30ZoQXsQB5jCoqTeiB
paAykhL8fayTDZFrt+VowckWC2t5RML+MrE7GJ+QfvY+c/qJbj+xIyggxY2RJeYI
KFyvNIlLC1gR1gonyrbz0wz1RjSh0FiT+9aaPqTsPtmO/Yg1TwDhUHR5/ffSSB5P
hOzWOXywPNwEovCirO1urSAoyGksBrLJJSZ8LyN8P+pkHXO+X5rx+JXOhhYIMC76
tqPg9msw25XgECxYDxnDgHuWrj664oIfiVQXrr8xq6p0VRVkRAapXsX23BmlrxIP
gkUtkHW3sjExtp+tEFYngSu9KvN485uXrNEwsqFsm3mIWJZZW4A+x1esNQclji8C
38iJyJvmt+oEtoTsLIXM0RViXJTWqDHNc5SamqRtRtriymNSXSZCoyRzNIo6lkFY
AXADxeJ0eFn0Vzoa3LN65jZbOIoX6oyQ+a8hjlc03rv8+sl90KvceC38/0eYnHiK
xMmP6Uz2I04jmUUJEZEnFqtbgkRmHM4wpO1uxbbIWaFSM//zysNMF1hjYvaV5zpB
Ew4G4FKzhfnbaIcKQejxnnPQQKRKylJWM9Yv1+ZEuqydbg5yaOr2nMn5AkufbWsH
UNDLcqhstrEpCoEd2QOvqZQyE8MHk3qD4M31j5Ms9CiWIs4UnMrRxrTRM3TWGLZE
N07+1PTVcFBldGCEQ60qN8OlPXNXKvXSSxaomnpM7/L48dfQEbjPp+82o0iZKmpm
QySUuemGrMBrNZcalCH59D5ZruNVE84Q2vfvvPgrRFNqvDbBausbPc0nbQTESjSJ
DpthG1oNeZkqO+b/7DVbCraHr6nvHA5kJ0fpwBpX4U+aNdLRSc83d/E3WIEucbPb
qJCOpXrrQSozSSk0nngHjdPrD3VBAW0ekyo/SEPcO/NgXSAknoIR9UtMkTA/BAyZ
gspiRpP5FIQgGMNbgPr071jdKlg1jsseVbg94IGH0gnMCvmK+dm3XQrllBJGvBr/
rtdbY92ZhLi7zfW2XzW7wgoJ9J9/2gDsrQAhVzJ3BovrPME5aWHj5NRlt2OJF+dZ
lrCItzs7ATvu0IOfVbR0e3IlH1F4CSU50sW5ipthGJ1F6ZQWMx+CHxyYjUPoltUX
6Evh63u8dhgMlZnMlvrjOrR/YYVmREzpCO6rfv5uhpZU6dPakxSNuERFlV7WN0kV
ioyipJTw8Oqyvm7pfC3aKmzlbhrMsgy1OHdjpddy1nQ16j50RgdqN8xq29AsaotU
5wnK6UDXp1ChvTy29VxtGyfxLqA5WKvqOMBNSMK0aXC9Y3l7h5jueTrFWm7l09Y9
scF6V9N3XI5h2oSzsMHd1oiBP8fzf82up+b2WeqbDfxW54lmDI7nSmrB/dZ0A8jO
Z5qDOFVHa7SIsDabVjJZawIeIEHgoVu1xhp+Fia86mjCxObtWU/il61bA/WRWMAK
sEdCj4nDDS6y33SYF/G5I7MBLc0hW+O6udz48JctBOA97sL9g5O06PQa3HpP7Meq
BSxhsuJbLu5KyuPJMO7f+cCb5atdQeGvQGTMY4EFyZMVW//ch56VBfyRpcORoL7G
`protect END_PROTECTED
