`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGK41H1p9dzUTrZJqvpX9h0ultHcmjgDXEmdbIR7n+gOZ9vLqJVMICTDZB3xllg3
9yEKTWOZs1LdlutTvNtWXZ5tciXFPYfyTiVeSkWKC8CVqXuQlbaxLFWouKlvBf0R
8yc9OlJBmL5uQZ5lQRWb1ImNfun8MydXXrVB6Bi/hmfwsMbYhP4MdCbr7IYgpiNC
TQIi2QTWsyWu04zchzNI0+0fqcYRmPFo1vPFsonZAId2DcucrQWiui0yVCD2/J94
UJw25Qsdpi4vSqe6iXyZUdYjPHkaguGD4mNMp6Pd7eE+pkSA17VqRnCBnRegzJmF
31Woue1GSZoz9KaRGduDcE1WHaQ3qO8OZ+ZY+I6n9WxZBKDxumvScfsTpuge7x46
JQrigQ0ojHEwJw4B9za2OHWk0Xgp5ch2vLvReSBivBWmtcU6rwKIyMFbbB/ok+oX
f1Ca/bOTyq2EMeXoir4zkZAFgdNB6ATivSw2kwNwDJUV486XQWpHUIvpbA2WhwRe
HrHb3/redi0+ZDEClX98DNlN0Qq+Bi4bvU8w+hhdurpbbI87wuBXakFEht7WsgFL
kitGSCHK60FiY4HUBTY39aWt/LvU0cn6R5QhaFDH8iQa8yChq8jh65IHqCYShFO4
zVy6UFJwNgLD9I8Ct4WEWuefcRs6fZkVZWKqeDp8F+I0/2fPaLdKmJIW+zvcyR77
KCvtj3iHI85hT2h/qUSHqiJWBhG1jTcW0GWWJorWM8K1CG44PG3zjk0NrqKlW8UT
IhTOHY7Ogpe5wqjTt61+yOspFe82MHlTmlLVwmE+vMy/w/XBa2yjzIG/DU8f8OwV
/XVXCaM/seJfukzvY48gffUZ+e/RmPWokBDTf23JdZQkP/PTDhyXCtZwCTa5B+NB
n2JvzFdm49GPN3QCadD+OTndXkkY3XHpNMw4M3B2j2SUTEiJisArukr2o+jemRqy
u2Nd+hO9dTAlCQyUttgJ2lLgw/BzcJ+7St4a+loI0Vi1OFG3xriuQtlwUg6d5633
d3sGuW/IMbOTDLbWImjnDjsOkSQan6gaF+4SXdeI/KXxsGtn7LvIiYqcFanFRfUt
n3oFrxcQo8oElrxijB0hQFpxlsrvjX2bEL74nLhGZQizw8W+Zwqb6ymHMSnZSjB7
gmCnAuwQqTQcvmg7c789C7DuTk4jgmkJrAKARtjk2zPiEy7GG5ysa66KrLhACpIA
2VjYB1x38COxSs+MLlw4bzkckyYZF1eXaHsnQw4ZKzVInm3NryGHsPPP4GmUHmkA
qWcc6qFpOpcbaEfAz/ruWxWEMWFY8kx7S2BwMcCapyJK5LnB+Kr/59Gu01Oaj4uE
34X1EOGPuvmiYLuUfjYA4ZFMw1FLxJE6KSR3Fi1NQFUXw2YGESseaQG8EBnbAD59
phqa9v2EI0U7Ko/6FLkNXdE9avLW895Kvk5X9a3fq6thfYDa2BByr4w/W2oET6cH
ri/8usMqC25IPSSN+e/C3KCbzd5VZpuWDNxTZekntpP4j0gtg69JnPcabUchlKGm
BHoewot3cVRuj0xD21dCqPEdcS0bJANRxCV8ksBsE2a0rSR3BRMkkMigMtgl3CU4
VEoV7xtpePeySmvadg30hDqt8QLUm1G7Wc7axMZ2jNDgvxFs/oICzPob2PFDp+oA
+EwKFlTiQy4XntjilU1jh9tgpXoU2BhZCZkdJjVQ/iTEx/4hbfeP6DhH5lDLv77u
SiGi8SUiCEsxK0LiqjFSydERIifRiSS+VNTHU29AzmeRgDyTuPoVEzudEJYMZbp6
zAnMFLqTHXmCOlF9xnqGadMrIMeVaOZvTrYH2Qy2h2b+OZWPIKrNh6VcdkLF8MG5
vf/DmLi83JuPcwuK/nTX/HObywVGv+PcgKDwsS7P0MASvPXwVx1uak+HUMx6JLnk
BOhILE4B7Bu9gU9SWtdKs3+ivyXJk8Mdioxl/qkLrdP098ukiMZs4ZkjCHj4GKxg
6ThdlyUXvMWRDLJr8y7mcQTSIWliZNZNfp/i2fM7WhYy+5/LEH+P+H/MUU9s7rU9
z6UfzuVWfb5pmfJ8plEMF8GRs0ISS2yCQJBOOplYqZCztbYLY+Vt0D3RfWIGUZms
HgHhAf+fjl/aqugchj/5TO0LTOWsEtB5YI70RLb6G+fO4JAGEDOaq1tlRdH5cltr
jL/g2Trb49Dq4aaIX0I3XmQgmNXyUBh0Jf3RssqFsDnz/yiVL4npkFw0SdmTB9hn
kalbL6dtZETgBSkrfTIwRkv/uPrZU/yXmaapUP6CpqgB4ia/9vIudFgXsRT+o2Jr
4By5YL3XMl0Hc7FQPOrGlUJ3j2YYwlVHuYjuRfqCLdP99zttZ/BZ8VTLJPFsSFUg
glQHxCeGWL7JyUKoKHv+S3OMUbVgXkMtGSbEOhwbO+hB7h9D9oOwyK7XGrhrcknb
xRmVh6mNShNQ4yx+zVp+8cFnPOUoiqqdzQ1dDq7xpS0Uk1b7wU2Ft3zNzNtEL6pq
ijxuAA0z/t95MjXsjD+FMO4gx5KsCVlYdqB7Vgh5wISWiVAb30Vjqiobq49/SvAz
0ECpbBs/jzULD4oJBIlH+/BLqhcI+3jD4DsRpFoYkIeVbISxH24w5NG5Py6D5TkH
NEPJxea4QhNNVMH4F7YNRPzmBJDHZjZYMvrHQpu0D7YfCt0rRIE1nJ/CfJXbGm39
nSEvRRl75eO3vtTLQatpfKuVEjvV5botXz7STa7tJV7xJPS8fxlT0ir8Vu4GSTSy
j5UtZYdyPvVPD06wD/JCMK0baeB0vzWfVBNU61X++P967A3vREQ/NCYlvPBfAglN
NmvCPuT6ojV+bLy3ZhfMmAzGkgUdoxE7MT/JJRl9oDVfe0OKEbA9j1BGZZT3a1nI
Yyjf1IjKA/CD2R/ut7Qd6v/rtGTKKE7kC1efVFCE7RfSz8iDAhhPikEK4XTClJXO
qOppsFBas/8JfaWd5FbOw4fJdlWAt0HPmHp/oMcDkR9alqUCoM7qXjzSUvBQf9bm
Hd0yzEQq04jki/NQYOkBwi+NjOB7UPeQcGNU0nsh5W84ztJZMtoSVa/P1AEtuWRV
m9A1LVCWxjleSi4GoX/q5DlAel5LIQ4me6ZKeo7ZcogWto0vtUhHgBoeLzre9iLx
n45EUDwN1WgrWT4f/rlZTbM8h6O5lDTVn7gsY7/+bRWOCb8nnRbWBj5cZOCvazAt
b2l4GvMbaEZKZ9vgV0niXCuqeLn5/3sacMEaRQLIxyv8QbjSvoIN+VoR7/B7oPNg
VrilPTJVa0LgESlBakseFASkcD2Q7JraU8nlyjNLfY4KtwSulr2isxlDf1mo9L7g
5ZvLUjg0khliv3c0clWfL/GL18FszETCPtrrR7CocaBZS2zamHmd8Gv3x5YufehV
EbXjszH7G3T/YLLtxv4fQxI5jsG2LQG8NvzRFa9xAueOP4HGWGlJe50xAzIj/Jp3
+tzeNlIVZ5BriH4qyxtfu7FoHToKmq8e4kpUFn6RzbL8/UNEYQYRrsOtTP3GmWtE
jxqd6ccwNMMFRbdDZvxuyYcPxT1KUc2jksfZI+OLKROhrC2f8IYL+4myJCsD4yxl
7bPleCTQmX1yd7ut7Rn7xApWHt9fx3DBlJlONpaWpDOCCEdOOqFisku62J+WATij
1geOAb9rn2U6qpGUH/17JTz3rYflH3kfYsO8T+Km3YRX0NyzwJ3W5tru2Yip90aj
ZFn2YRMWBSiL5GgrxBMPnmRDWFEdjnQYw/CxS+CFdCGQLTz5YRzWWAg6q600Dfen
G+PBQti64XqN9u+pAe1DpF1jb6aqS6v9r5X/E1CBGg848NOHmjBEH2q78UpE3/Hq
PDAZuSe9rMb6L4pgcoP30Jft0jOi/lAOAv4vkS26RBVsT3E9tZc4fJFFmdRoRUGA
bSECcW6hsgW3Eplcj2au0AS54lhI+caQi/FdYrK3g5916zgGNUnbWTaQVeWzCmpc
IunR1xM42gQgkucfGdCDW7iBwOLyipsBg7zEbGpidtOnXG4XeKmW55wA2PmhAIpZ
zMe8Be5JkhjVnanOZ87zNH+b86ENR1fWxy4t67Q4Jvp33huXW2x5rXQ2V9kCLT9X
MeqePLn+/IMMHRYKgQQCSOb+ymENpM90f5fslwhukGWqOdPkbFdt/74LzhnKoM/E
dpkqubqjdAkMX6jtv4p7wXqZWEifdXDd/GHH4quUDjUSedOWZw6skC/Hj/fJ6Y06
P87Vy+xeCtCVd0TjeRxNDqqlq1lxvW4qaDJXxSxn/NR5qpqc/Ai8j0UuKtOE1hv2
/tR/zIgo5PruUpIK5sYflJjuvlLb4n0hugicWkyqQiqFcB1Rudoacb0iuUE7CM94
PtffygMs7g0TTDXRuyv9BnDXr/5B4A/2c10oHCyOhUEqhgzLvpk5oXFDufE3974b
gEK8qkzSRlTUVPsEX7F5KVNi3NniagDqamLLIuJ43eajvoHLqYCzf/j89U9IQQ9z
zb/HDM3lIRmgNmo4zx4kU+bsjXQ1HG/AmuN2/NgScZT7OU2gPZz5zzU8jvscm/8e
6OsA54bzqfQ4060xONMNjUXAQuoZqWk0eY54OzIjWvfmjnUGn3TOX+9DJseTMtqM
FmuApXkFXAZ0fra9i+MTNw0Mh0iXLZpDsrTEUmlL5Bz31BYbMOnrl4QKsUYJSNHk
xNrUHJYObFyKO1yiiq56gE3nQFrdCvPgp94eN58flNpACBnAvxag7bMEmBh5ey1E
KAl4qCZWyF8gHXsCrxJdu1qZmm9SKiF3LRPxA9R3jARl/i77DaLNk4G0xRrdDIsM
xx3RBwC6Vo3pirH8M8tM/4WsmyJcgiJr4lMdWWsN24rZEm25CJ55jG8TCc2+r/+4
tLrX0Fn7FKR8G4osF7GQB4pmr1BFK4N3cqcwUyhN1g8+b4iRZtZOtUYcYJ3jIvZY
SpGVCNsu+3mgmdRNK+aG6D39iww5OCWGw6Hw02HLpD8e5e2Ak+SBMNVa+WzKE44v
VfnQ5kzh/h14i2jqkXiX3IQxHZZs7L7kYRvn/bzPKEqtGxEUpnrm4Jd+2wk78gPI
CywbCv3ax/0VK6s1aRgwprumMdjwAaBewvF7k662Bk6euzUWh+uBfkLHSh3rfHgC
abQ9es6KhV6bB5iNcC8If2t7USLOKRvcrN4xq+C83InvvajC8fvdP+HArc/bA6tf
UvuT1RRKgaMYeLncma2Xd+yvAgduWH/s/1JSLTRLdVT0QE+Jfiw2VS2jqTm73t14
3Qq1cJyrI7EmK/CjnsLg0ewp7guLA5LApxi0bYiAKZBh8QIDwVJnf6i0HEzmqly5
o/YyaDi7sDaJerhThxf/PHxzqclGz+QVJpYoGCkuUjod7xDfPK+4Pl21W8YVmuZv
0d5DBK3bjl/jUbh9Sb8HTjLuHrQpudj4ihuEWeqNqwZjytQDk3XdE/nJTQCF/tMN
kpAGiJRal8opvoLYI+hfmBhOQ7zCcLiliR35aMe1lAZ/Qw+VlTgiVCn7GuCuDstp
lPsE7RUEC9LRsqNtxphpFJiK/pTgTRbUSy5hrTXnMIydhlTpUqTS1JL3XZpYBnA2
E1AmAzpUcJlp1SRIZsvbOzA4FCChQZgPbIf4cT6NnZvCNKMvj+arTnKHY0yoPSJ+
dt7Fry5zHiCrR345ptKkvJbgbOnIVPcOIQu6f/GVBeAnOE+yo8DIVJiScqrFHjQh
A2+jBB8bS30f+r1Km7qJ5rJlZ7z8vjfLUlLAnYKu0Rfe8YcMeRFCnAtknccLkHG/
KK4nWde+843Ss0FJ/l+Z/+KtvszccDSu5SUeUNSPHVtHweg/ISrKykahH3k/VN9a
4MJzebNFmji7ejdUmprfmjrp+R69hkg05qEWRSqLgoBwCLNYkEn5Pn4LZCt22o+P
ouAZlRc4VXc4bm3OO2U3CxUMCCRgX6+d5Oe8sqguCUDwcNd91stgKqhYIuUrei9W
AvImUdYaurNuUJBEipXufuQNZs39D+utsh2QdvrDARwQIt5FiidVvFNlWA1s8pEz
j3pKak2OzMvnczFUBg4dFCXvZ2L6ZSQYiG8sxBbLVBuhxXNIWf//RoAtaqhk7YLF
BnX2bKCLMbFBG1dH1rI7aQ0HfB7R9DmueRr/STOSxK304zzide7lyDSK+xBC02d3
aTPhJhCf6QFzXVWvsiCVgJBdM5w2q3zGpUl8Rvd5bmbTuWHAkhpX2ZjCd7O9kuCa
aEq86uWGj00MlKPYX1HqVLe/7z9GwKJENxce9gKALLYoVjT2OU7UZ8cYm45T6gze
2a6QVuXdpr7sLJhxuKA5tftADKXgp14gC8NJXn+cRvElHd6y6E0+oEODXxIRxdJX
7kic/R8w83UVNXlMqdvq+treO8MOgWSlvxOGm2eGd0P9gMFcjBcm9h3+j9qX6fpd
wpSbr4p7WuZn1UKB/VSOSP8wbvL4Bx9HWIzFL1GJ0bWLraiF+ZZG6PXMTwvb9Vut
HCvWmz+QyOMtICRC6rbFy+uuE7QcyKKo9eobZh1/QRy1ubPE+OBSRbpnENaXlkUi
Istfj8p4c4mWByifBuQn/xF0ICi4FtD0HZCwD+ySpvfb48EotnhVqSdcBymG+vxt
4nesBA00s44WJsl+5Fy9tRTIgrVqcoo91YFI0Bbmy3MHtZy/1PmmByaP7Wi/iXF6
1iG97Cp/RsG5MUuouLJdBHgPuqS3JO1tDXsPlLSotOl/2y+MCY1ochMmiQNGtYeN
WGq17mGil3pBGHvdGt8xmwxPcWlBK17TFHrfO1Lv03wQt1rP2KnohsNhiAU3lRbD
8ocK7RaGXIm0Bhh6HPNeCPKfj22F5OkTDD7rQX9IPRvzYenwApmrGeh921sTV5ZI
YxlbI/7xcHxaC6nZaqtC+MYV+gHVJBAU04sZTfocQ8SmFLNRV/2ImzkahmjLVCdw
FPQZg6qgPir+CK/EyeN7b0Cj8DR6o/CMc01nMs3yvtC00ZN2h9234iZYuc48DUDW
M1UeoSFNxxCoWtGJvsGAynT64RF7g7vQNH5RYvydvLOTs3Dplj+ee/QMiOG7FT6L
EPox747x+JvIf71gM8EW7EdLeNBNAi9R7YRgv8TeetO+wggFasdfoMPGMMo8NgPl
FhJOfLLIG7WvJ+u1cBlPWd9vXtYglbzSZz5zI7Dnq08VTutmcPrh66ub3SMVLTad
YGxQN9Hh5BRyw+M4HDPdwg9000gguNV+OyWsLrSug4Ds2wMjWIUanmiuVx3GfiEB
/jP/G814Dk8awbHtPS5yt/Jccbk/Sal/5jcjJ4Vu7w0=
`protect END_PROTECTED
