`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6W2WV8fWdq9mZFxskvOf80cm1f4X+YzQM/I5mj05AFSVKH0E/2aC9TOyCDs/GvuZ
OhjBWGO5Yb85nshR/Zo/EWyqaPn5/ix26In1fhKanYrR1AR6rUKNN4xiYbAuR1Wk
MDPbzbTuZAe1w8T56ob2KJDaue7FLdO/Yj1XIWqkO8wfNzniMS/G1DE9a0en7M9D
SIW9SaRhe1w//EUnAwPClrViRdBzP6Gs4Fl1yWU5njcI5bffKJIV8kspUxLgltVi
DtwBTWWfGPcldDvze6a58o+jcuW1NWz763+rgdS+7xMBbx/ujq2My+8dy3M7LLRx
7kqp1/Ar7pl9SiHORvzL6dt4FBpuKz3bkqDaYfb3yHqDxFBdU+shD2lXcrAKSjCA
2QFJXA35LytHQSRhPCsueg==
`protect END_PROTECTED
