`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a68tie4aEbyfSZ+Nu6SwyV7lR66+8eOQCUqoR5KBzJON7GG9JWya+Q74/SuYNx+N
ln6EjvdVUjwlLKMsZIT0uxdte2gyG1+sSVcqHgK0jlfA/ezel9wFbidWq3tj18l2
KZ7q0TTg7pG2rUvNAstTxODszm9OoOzZanD+caRVw+a9PcUWyI0o6s3zI4kLpn0/
iP3IaXkqU2mlB2WDuqIBhuypBrTxeicy49k7qEdT2O60idimORC7gemr1wYMzkRw
9tENgI0tiMxmbXsxexQ0vAMAXBwPoT7wCT7V/lFrYWah7WbuqSPX0ngLe/O6sEaW
Ud6KW2vsRmnlWSRdHSGaUUSMDK0TpuivREZUNpC/u+HXqMlvWGm1wjaS2v6QLsZU
7/joAlhBBHrFtikdV8xLKcRNl6z74tApfzmhM2GXcWH3IxsBftgp8igI8afycn1q
RzzdfKiMTt+KP5Ljy7nMF1L92KlFJR2MzO4TQ+m5fEzIS4UDIJ0l2QjRNZkJWF36
1WdkZ0+LynfV1X+OVY8mGEB4Tij0kcMv7phPXOc/b4Ciu7891B82ZGzH3QkZg6VQ
WlG5LyaBWGRlPOaGxOCUUGiA0AQkn37fvlfRXEZsPe7Bz+wG2pGB24qL8XZrt4qn
Jzxyj1yx2FzYFyAU3XWuTyDHDHbDFxWxcY16PM8ta4s/EkigJcbxD2KVFTjsESDL
ImXt0ZmhUET+cmekWSWaCZTddPEG09Zfaoa6C8qtTUk5kq3PR6V+fhz1pN5JkVBV
8Ke2KOQ4FIYw1kkQwSI/4OHS/PiipubAzCx0E8NwonnYGUYlXV46yGAceJbcSLfp
6RY0gC3GyFsgnnkMl7yqOdgSPb38ybKEjK8tV4MiWa2HmAHr8kB/MzfVknNnVNaN
JRGm6e7A80KHcuEYVZcT7rLrUHBLsFiFx699fu65btRo0SvWK/+/Yyxdl7qEHSUG
33qh44LZ8Bg1Ku/g/a5rYwPJCvtOziLtM4rRf+KGWnf+lSpPSfjV0uaOq1jcq2ut
bRfPaOD5Uvk44obGteLNP+lfTnRN/TByeaPrpwI0UW/fcZO8jX8FDQJbbSbz85Yd
gRpM3ejqLIiUEsDHjj5ZO996iPSW7rujGdYLnVcj1UBaWVXevMTPJTNB6ERcfXpE
4hs/CVqGZMYMcWudgbUVLyf074Mluwy7gCDdgKvq2DIOqr6JAJ+VRUs5PCBmcpMb
umfHnJMhbjTia0EeYDRUIKpVCSID0Dp907UIrzqOzuxm+HVYpLc0K4Y3juNkWBGQ
SXMQ6aAUTsPwVzHa+F6xurDUzws338pg4SmAxm0LpDgXH/QR9khc2fVuyXnsR21G
gTQOCMu3Z0xLxIfApvvq6YTs1rtnaaZd3XK/Ijp43QNthfinm4CoeWfnqsdQ/eEg
cj+l3Qt1IIzpfkUs8ynQZ4KUN8IdQO3ok1wMrwMwSWtKNRulIkZ5pPK8a63cfu+o
Z1k9J8/eYX7ZIgIne+tVmT1Ri548fvtOmASGnCv7aKkWp2gj6T/WVzn8GVRyiBim
NkFNNPwF17ofbBhzTFdW06RVMSPwVjjSJM+aU8q8oUZu7g7fZY3NbsBZhrXsPK/6
1qZtQOveyobu1EPi8+ezk11IPpap3rEn46r1qkbYf7CaL+9/5yO/7pKQZtsK0VrW
fL0CW8i9iAcxbu6TprKWLKGVqHaGtBCX/wZu7IUZY/y/rrm5/hGCvC4HY2EUH3Xf
5e0mvdOdivMmGPVBUst9K/1GK5N71gCrLqFITY/dl2f1Ty+l/q/DRQ18gonSLMu8
YYRsfLuc6rVPANzYzOcQzDZJUdzOlrwzaSO5B+cmzMYVDgnckAS3Kamy1z1Fdrol
klA3YDedZEDnw+xXDG+eu2BmgmZ0+Hkrqf3BCgTChWpkNFnUebKejgzmtV/d3voc
CrgzMIeTxPtXBoGcg9ctRot42M9icV642wEEPe0MqUIi8fawsf1jkAUgoG6MZi58
/DouDHAWMvzmClT7yrSxOGkBkuql5svNxO/0LZUP5/k61sp4eLdjupoTF/lWd36A
Gvk+x4BJ9NkNrZVlDr5VZAWbSzunzSzXnfyQdf7An0G9TaIMSXnsW5bvAZbjJihu
ww9N6qA51dl0nJ+Dho6bhkGrrelDphJ8BuUyxCJs4bxM5ci0pPStswsj/tw+bJol
JL2U2OArpUECmnbl4xTxLF28hiIk4j29z+Bp5C9PHA8NTPV6CwlglKfo68Gf/RDl
xIny15ZYLNDlAsdlGEkzxi8glatmGyt60IIJT/iNGO5OxWyrlfioaAaJgAiDGXYT
apwxxdjdLXEndk0+XhHbHyCsiFUDmcFK5yyMZPYddkdLq5BqYEO1bjX/eNKoXcjM
fw7N0efjOFF1523ovCLfc4mOWUw5+FILWLPKruAisg/UXC+3OzQN/z/AZDVe5rZ9
eSxeg4OIYRfFHegXwEG4sl+L53fEB6poqarAA2TQvqL1tZwy+l86HLXNjTUdxi6G
H2wEG7MMZ93xLaSwPgErlFdAj478q13+aj6UfY7VEdqY91bq0mOxcLx5TDMohUU4
HNRzy0pvs+9TZRSZgJp89MC31u0JZMijQoT/+esFOFXhLcUuGKSaLhRkEneCNDxc
3So6s7fssoiiF3t+smeOLW6w7q3JGHLWGL6vxzvRgSyX0uD1/nUDg8gioMZ39dvW
WaXzyVahg9JgT6oXdhTzidCIKulG+u+KMcbvvC8Lo7agOk2FldPeYVEadJ/ykMD9
4gOJ6VxjM1HZUx2StVUXeP39HIM+9Sh+KRvjUJqSOaMwAg9x8iybykzaJpeyMx1K
4MSbhLHcD0ssSzqHvH4f5+lxzz9ApjZHBMsS1Z55tcqDn+Q3l+N1qTEPd+XFKMIP
24nc3NEOmWTctkQNXuYYw206PbH9V8KbXiM5jkv9IzNRTN9dwSaAFkvtj2iLmikO
Y9uGlMMevajNKace4aVPiZOoG9w+hus0CRzN5zQ4f7KQl626kxxvccTuiuSWs47D
0SwQGwvLHbOM5TSuwosaNCZHW/n/kXigcIinnZgXxPwzyQgiwcWIYnJOJeB1ipyy
JD8rzQaFz2wNmUJGcr31urslJFZt4ENYgccnoVMgc55TKm3AHUwaDKf/dstPLjn2
XtArxCPpelz4McrfX6uZDhYTUgncVHQkPKvCv+neICgHtttvwxWBpdYFfkDPIeey
z+b4autWUEA9f+oA+U7fU1CLAPufO5XMnUZ+pfoeQvrQLw6hdJMvU1hmabu8wRjh
sJUHhSLUwyUZ3UthiHzKjivTpyynJOr6OzaRYhX/1qySkdCp1/90Cq3jfYrfPZc7
wNVqmAsgJFf+pGMcJM9Hrn/NUELhzCKr0dtDKnnwj4SMpBQFGSTuCglZX/s00QXP
20ABXI5WNPIVqn0ft2T64HpHbe+5hyt9LoPHs4rnzpgaqkNBTAhlY3m9S2XcVQqN
eg8ibKdCk4XrOa8D0P9thiNuabBDYOpFiQF990LOpSPQx91ch4eRyFrO+dq5UlLn
lIoVJYv0je1Mm+t9NrGivtUtfLJZp6msg8oK5Y0CJIAQsUjkQGos33GLkFryilv5
sv0MfRI87/mV53nsJpRgspVza1ACxxWqNwPlHMXFZpM/zM53Kqk5oG4hRYSR3rst
0ac4tmhWNNt+tTKXq/YfLXU8QjZyl2fZ8LqfX86PybexnCNW+KrEn4fyl7++emLv
3+n1qDmQhQzz+HCYN0ZLTfOod4aKe/y7/EB2HzgyFK7vWJ4HbCOgl2X6+YB/qWmN
qtUEsM9qFSt5e9sBzvP1Ef2sePbirmpXpxmr2dQeRRcNHB2JWLPK8TIHPtNeTIqT
IptsR7T58G8iRfANtalNCkYbg8IA50P9XtWUrw6Mv+tpeolQPII26flwodgZl/OB
CD85jwBRaR8ohC7NBbA5kGsfadlWN3phuu8J2STF1t5c82yUJTxBQKdy7hXaPfeq
Ar1IVG5Z3WQDidV2bMFzvucOPHu7m268cN7h8FNNTiBzzA1Tvao+fNTVtuqmR36i
boaJPIK82G/0WJGWj7NbrRAS+Y5B9lsWNVlK5TvzkZpnxO7KJlq7hl4zmXEVZYwu
8KaSb49xR8i4BoEFI2QNwLFjXhFvz+DZkcb41WgGLLT0qduL70d4docmNY+dxhmP
ES6KNrno2ROIbkk91t+GbUn69lBs1lbMj3tdEhREssTB0/7tAy+6o2SCKQZEmwOP
+anc1kA5w0HS4WKjMk9yv2VRF/rzbZyzv1697zib/6Rx5fJm0zoZtY+E9NZ9VhgP
xAWvfEKfUcCXqHR7Def/8F/SUdxwKd8Sj7lBMLIUEFetCzxhQVHaHzpAj3iY7uO7
e9oIN4ceOaAososVTXplH5NtHmtHx3AMRem9H7VDXNxwVC8KQhG/ME5dA4aF+wSa
70G0n2bkw7/9WLtLsQZ7zvvLh38NGCvO2Uag1dM6oXd3lQrZQ7/7GC/QR+ME19P8
Q9NzeKJf5Vo1KVd+OoNrivNFRJcb+hSfwTrKLTiJjlGEWwsbKsYT/H+xiR2tZSBu
wjMlbTzjj/3J45eaeoShFkHAxnmYhmU51HEGClcwwDCR1v17X9Rnt+jYN7L2Eueq
8ieOXhG9E7swuCfOTcz3gjnEcUkN9K8mo0WhsrftK+Tb8yjdXHPBBLZaxALqrjf2
nfMTtpVryU5FOLRFwM5rcGjb9mcqeXQl44FXG/gO6XKJ01J2cK8oMmW1aSr9cbmb
gU5F1i3SoTNQiRbXNFqMjG/BXABB4tjLnvvZfl6s/E+OIW8oc4MP/Dz2m6CpZrZA
MMOwhUnutV9G2x4lRfHABpz9pFh2sH6j6SIyjfnLdoARa8/CU5DMflhD1dMSCXa+
yfviB1jpKq2+hwtIWny2vW/w5R6/hARonss1GJ0X/o/ybcNMNv9PBuhZg+Y7PcbN
3LSBl2scxMCf0lY4cvYNQPqI3fnFaF9kCmTbRv7+xo1JVpII3tn1/UQqRoBJkCus
9Ej/QO7G7xZCqR3xo4wg8Ct211hWqkuCluF0gA0rrbde4h3E0NcZgE14bIjRtUTH
gd92EbZyYfKzQyrAFA5i4/7yIzWRQAAFauEpJscF8Ce2rQPWVr6KEd+Y9tdiiCxj
EWJXaiHrcQKZvCJiJseXya9hpmgzH9/AmV96hLvYV+y3Ah7/6Z9SGj5e9kzG13Rx
frjChnjwepEmSfomDG9nKuPec353RjWnS2P1ew2HWbaOrgvYnlvwBvq5L5KL7xDa
k/WOjveHn3QZT2MHySWC/bYKEQE0O/ohaml1lNZVnDpUXl+8VrGBNVTL1HtP3PXn
9cULeQ7gqkIy2oDL+JkrEA==
`protect END_PROTECTED
