`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhBefONFh7rI9YuYdmOj647UiR1PvLvnjS2k1CgY1EqtKh90SkeaskTTEcqlOJAG
b0H0v1vgLcNTB9x0YQexvYX0VlG5QesxyUqpMdmf8xYxT71CICe3SPXDW9m3xip6
xiKePXy6RMuF3G/0LrkO+oBPCcJnIoXIFLcAp0IWHqyU3/1fGK/ZWryPiVPpKO36
9DCrKfKvBThV6Rl23OUmzQNuRZe5kvq2EBbkBXmplDHBbNbk+E0pmEEAHPUZQtXH
z83qvE62RJQ5cNpE133LWZcqjBeDiRZxtZKdRYfWct1RA46ifM6LaDdwdzFzbzgb
tC6qypUfxdkGDQtlJvY30H45cqMgVB8okWgUCIdc2KIjjC47KOQpp9gIoT1P86Eu
pBEjuH4lAxdjexzc4ouBmLiik2RkgdK5rIMFnmn+6iwtrmebXFQ7vvQ9zWKsFkhA
4t7cCwgOLfxXZLnpxwzuK1mstZZDt5TVIwlaxznpHMf0PGpG8HZ+I4jZVOlLueh9
MrJ+qdaLuETXqWuBUnlQ53euQm2v4DkT35+fxj9Gxchk1RfArnr4ugDuXEpPwpQg
2DgXjifEl/9ovqe0+NX3bntgO64ppha2jTytwD8Mvpq3bfglgNTyRp8qxXZAtRHT
qeW9za9l0DMeIHDNpGydx7hxIMqhRbV4DhLzNjFfRS0CSlEiKmzt7M/GLHCHw6J3
vl3w/4ynfncELGkgrLXh7GjY+DWy/i1Aj+TLMcecJBk+Og91znvBuxsV8ISc1NKE
AorhlbvXoiDbHWbDTEFKmas+oZbPpqbLG7ldLOX2OOEuIRN+F9ow70qCzanmhYPD
LjbrOihAq+Uw1COVd72o+hNYMYtHDwf8xNzNCVZxHmny5of4Mhm1+SopQwJdV6kl
EqgWmZwfstfoKm/dfIaRXsoOipnxjUYluXXjg2KCH7jMgUd3LFyG/0lsM2sZzycB
gwtMSS1752yOnGUVgt4AV6d27eOvBnJfMvHWR7r7nG9DoMe0r523/7AgShS1gd6d
uxbbOjGHXPBsdz7Dt3CgN8kvFmlEmVMynBRNs2PiSuG0rj8cVBVntYnbprnwAs+8
DlB6sIG7eoFAKYN8sgQQU7+xwk35yuWtSInzgnRsupiK5f+sTKozlvLFozGbmVqo
mhX4/HEJoZ6o5NmxWOCSDXc22VhUB81LbtoLnkTb198lWz++4wGAf/7E3J6K+zn0
inkbB0ATdRn/mqjAZ+MXeH+ZOtixyq40zlYtiqRi+yE58lPkajePxydipjTdTkQR
mDCFR8I3jquTLzfRmKA4BNZVTvjO/WzVGf4Nz/yVVMQYB7C6UPHhhNPqZBsCqQTx
2O2qtQl36kzUktsseHOgW+oBLsTZV0D3zf7TpvlqG+TALZpAz14aPLVeOAlc4kZf
QhoMwp6NWuZjBm5pmiBEQ7FtN6aPktE9+ipa7Dq9A4xnJpw3kwRWQy11TLnty6Ca
3cHm22KJVH7qEWP208Ysa8fRr+EOAJgPFko+uD3R8yaXa3ejNvwy9lBBtuIL65UG
pHab1zJW5w/45sVSimVqtykTV/ucfUHxy7uYmR5soHeaeh6s0C9Pt4sedUd60FYo
aZu+tLT6KAHdXIw0nzzFaNYUh1PyDGs5PC1Hs2n5jIsaP5uLVxmxEPKAgjm9F97M
Xhc0Smmuh+7evfprEmo/sUSYP6k5JLbWjh5z1kMQNyOgnPuCLSr45rWtyyRO65qX
aSuWZSi537iNjQEIcpMRvgLOHXMzapBwvADAIiaSPW8wwQwhdArUHBoe/L8rud0E
F1zqV9qrIk38G4ZSzl3CLB7qfELX7nSkdE070YMcsmCL7f/ZTVL5XJCp3JXxaE+z
CMlUbf+MQVrZGTwK+RfDGbH3kxIOBwnxLUAyn1h90vmUw+1lAwS09ekdG+/+yWNm
CXLkZmmV4RdK+/J3O/mdY8doE/pRdBScqQUR76PIYQQKGwrGfJLA30J7Lc5c/TfG
mfMAAQ3fJBRbwG6UET40Uv8E/hmEU2BE8vzzoAUyJGhdHhc07LVpzNHT7Zx6eb9e
atdHDNT06i4kiSNh64rqu/wO3eUYvhdCrOyvgbTVzczL2xs2xCgiuxEPtjAQKFal
3vxq9exAIZ6qNk3PdN6xbQDkhFLQCq2z+t/nJLVS3Qs407icq8iZ6Z+qVgbtSSqU
6V9fj7+UdR9aSG2ev32uG7LgUBB+b9fIJpWR/bxTEiNNseUvQoTERRrM1O8DeLdq
SmjgUduiL0tVmUuotQ5umZH1C8LuUpCh9En8h7dVmnALzdUHdg4GgDgAoBdkSN1T
Vt4parj+qcoIt+SbAkOe0NPXF5m/BQmCn6Q1q36lJqt7hsnk7t1SN9cHCvpXBSWP
XB3NQzLE++UhC/PlLFzPCXIYb5tBHC7bntBaOVbzWhLdLd+vavSMAi5rmJGmoq6x
v+XpEL6KGMmfyMNA8kKQWnOu8mltljll2awuuZMDpD9hWwgFdDQEb1D+Sp7BTUaE
q1YxNXk2bGSgWPFM5OqmOYw095VdayCAZp218HC3xoMmlJOMk575Fbb878R57sFY
GfBNjQ3P5GvX0ZLuNenpBOf/mEymxnShIU5v3szcpF6dM1tg4sS04sxySdwpdfam
OPr9VZWJMHk/V93OfvNI9OFiMFiTST8loqdOdrh0O3SuJIdnyHNXzO8f/NRGwhFg
kr0aAnPMlgFTzid8mxxItQok4LMjcdglnx6CSe5DqSsuEZQSjI8J6LEWDrXB5uGy
x67rG1w3P0PyLB73SR9YhuLFk76nW7vesbNyY1X1OOZcKg6ZzGq22nMrQWTfEjFw
VByVXXPM6VrOfbAHnghV5AXIP/5Xh7vNl3e000CmLgJqga2nJ+IUdxK6/1BU4kNy
KULR8ul2mm2TFdYkkN9fMh0n6d87h/OedgQEFbJX8QddlNlJkLd7h47NEqIZ2aHs
pxPkXW+BAI8/PMFXLG+XMwdrYv7opIqCoLRHr5KS6n2k39QvjoarX2oZYfbV9SMt
NCKY0Mvr/Ri9kTQ/eZ88VmkTg+8mtwGlG3GyrNnYjdAH0w5WlqtxkmZM8EDWpxV8
JRXAg3o2uiokpwvlSWvbXYP95kYOobZdLDUDZGvBRkbD4QD1agwJhrkL+7lN9OfO
ahtcEU6DMEXYsiqCPqH655RRZXjZIxv1xxhemj7P/F3z7vPI8C6ji7oyZOqNhd6E
`protect END_PROTECTED
