`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PRg3Nmm6ZHjZOttvSySkkl7JYFtTivRr9alAs+FM7JdRnHdWvS+lG/xblnm0VNkp
JnpSzYcyZjyVHe9pLyr3vI0Jty6NZEBtgnPVc7Oj6DERdZwEJK2NBagmfkJqoFlz
vPMLTmJRx/BiOSYIEyuwWF9elsXdVPpOo6tM0HkvqDyUtX2gScp+O/m+dM/UuIJl
FzUD4+B1VL+U40b1f5E2YQxQcD6K22tHQ3LOMe51BbFkInxXwbP81dz9zelenQZS
7O8KF1dlvSXsJSamhRPm5z85khdU/kx7jsr7vUjKiPYfoVzxbtAgrlSJwa2pm6tN
FBCCOJOZWvXJTKUQH7Uow4LgpfNzA4wESAismN+OhtFXZcGTrZOvZ8LazyoXboc+
imt+Jdlbetymx3rpC4j8594cEx/kiA3gQtBhsITjdX9Lq8BHS1HoSCfAnbJA31Cp
P4AsUB0WakwQ5TXK2ER7ji5Cu/aG+hxgXrKJvZN3VqpQeai7DXWedc8ESCboF8eQ
/A8Kqvxh64wykzh4vdYyn6kXNoZ+pZNbjMR+fX2bY89x5F+/JIyfIA6IBKhEVrrO
`protect END_PROTECTED
