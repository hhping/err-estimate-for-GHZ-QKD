`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KW6U/mtIT3f6CbwqIX7Q1YY1ds8DGSkEI5UA6e5TP9RaCreMVx90rzxoe90fvmZA
rN3x63CElxeRpyWzcY67pwEQ+KokK881f0S2YAmxk5+i7lXpNOu1UjphGO32eWZE
+VAInDPEqKgAZIZTD8AcFSPE+hKC+jWgoffjfep6enc/WL2ngBUZ5BU9P29BQYZY
nr9bs3iee+mwUlc22rZ/4b45paO5fBUtMgsGHaG8NKcbZHdlM1b4T6Imc1E++15W
yMA462Rl8z/9DCS27H6ZSrUbLzoGU8ChwzBODF7jQcaVC6xV/F7QTrMCNOyEWVvX
V8x/VVTanhzjAfqTo//KaNT0rmjYsQ3AP2e6Fu1WFoUbDQ7tRBRVrp9CAk2s4yYz
6FtI6JmEerXZmGF23STEU7YMSy9EXu4vzmji8cfj5G/QdNYy7z7OwGa5ZsBsN0CZ
AmngQ5Gl9JJByycpQqWrEZKf6LG/zhySoLIEmI+JogGSVVsn8LG7d51YgjXcnUYn
/H6LyG/2HZzudef2mHLORh7FLYqoOVO+cXaBDumr+33O/63Il0PSAHoJs/VEc/9X
AudOKFJRY0xfEdMtZVPGo2DH1dPaKBZ4nZAjIsFAlebt1gZhBpl81ewnfnBBj6Co
RAIsMzQsgNN/HN1GI1tdhRYEv9DbU/filhAy9NK0d2U5qcW8YcFe4GSuPiQw/jzu
uHBj7vIK4ioWQrKL6/THEsF9kwdweQ0ugVsbMFuoICXKnD8MvYdJ6wO5WjKoxycH
x5mXm3X0dgViapLut5uOmIr1xGqB6DGEeId0q2n2SZLp5c9XUWCtRN+K77A9X0MA
aDkCAOJcoSvplKjfnT5ueUoNUMe9m9oQMyiIStrpkhLus+3OJGgNLOrZX/TZTlF+
o1rTFKZjU1ZL3xFyoDtzBrlLOoRZN8T2A5BD9fGtWJymZBiq2s36HkwkfOLn3tFv
b6MKlbx3hj703FyFALf0nvQyfOFvL3gUwuAdJS25gMEhQ0pxqVmtXeZ1AuXE2cbs
6ZyuzWzLJ/b2LncabfOZkfHBfdxnEs6h48xzNg3sXxXWoU9Q/Elw6eCiRo2G8AGp
nvnX6euYUX4Zfhbdje7FjHa+VGxUFuojNemdkuYuI6Mm2lUE0SJTFDsZPLfvvrBl
CMuH1ktne9pEM4bgAeOgEBzEZQ4RIbaLfdPBvG8t15hQXdCs6GsTIcJkZI1nxz7Q
vKPJnUHQGH/Gx/ZylxduFqIaApFRvkwmPSi1aHerxvJzwwtrju4xzRLeaMCUeLXc
z+U0ohQa5env/5i85/CaebAXJCLvCtYGy2fdAGq/GzMLumGE2cNtawPsds+EhoZO
6zXXVYDkfUBbNI1+nBv5PaYmxhXvDG+eozNWTqrCBegheikVSkXsyN13B7Zp85Sn
FWtzvx3X1t54uz9GNf9CxaZ8pgAf7IPOidACjuDQS5u0w33wt6a3sUW9J6t+KKMZ
QGl788fZF45WbOG3OOSzPS5gygErfu9XKzh5Ayb6z/Y8dlvKHM3QUhpy3/sAvFWx
GWpQQb8nITFzX/EfO8X2RYVAjNEHpncuaAfxwVYEasDGVgaJdxxwsdXSMkHGSGW9
zaOYfLx27QFDIsgJAn/Gjy9yvJVHtfxJMzJm2gcd3hzUj+Orzg40+l3NdWOo0P7Z
PFNgMgP03oJ6U8q6WjWuK/oIqrehvLAexEWoCn4oskT/xjPQ8P0Z4Lt4T5yNZ7xC
9hZu+MMebpf/tAfsd0ET2wb0SFVErNq199Ky4eft+CwGvoYW2ZlD9EXBAoy0VEiv
DN8AGp5yhYpTEPIO+bkPwTQpPUKl3dXx3UXlVQwtghNnlzX+H8XDlqg05WrRCmVs
tNFCLi02q/0YyQsGkP0f4ndNl02hcPd/+ZvWvvGjfZHQm3i8IprnSMoB3bF8PoPY
zfM7PhWkP1wd3WK9dV5CbnkN/Mw8zsaGE+r0lUR+0YRiuIiqTxTTVwWZiBMPeQS6
QFzHGwmC0D1OiMuwAlxAE0x+OdAaa2qeZTLuPtIhpkrxAlSJ1ghr3ifm1Aos8NbB
5TLPv0g/emohj3QNr3/Io14eCcw8RYVtrQ1/f/Yg2iHaCRJVTuc0XPZM3ia/VCzf
g97hFFQpSILQIlwkqxmYzzqok9QBjkCkEvh/kI2Vd/bbYzzAwjJMIwWP0tf2AOSN
BnqSycutnkHXdQtpAk8QcQ9sKyTaPEW3hf2w0Dd+Er/x6urEidhkGhfpR3jBDnyP
tfPGSynARhb5R89RlV5aHyIxqhraMH9FFWgJDL/3rJsa+c6XtCHteS7MN80bXfZM
td76xWCISCPWUJmw4EZe2NzX2r6vLu6GflexDbu6s8VQPeCOI8rbTRgIvSHwhphI
YTeTUWH5u5yC+zoPG5/8ftLCmqXxi0aG5cuTbnaXnLS95/cMqfH1lVIPhlmLSLOs
aZQUGctCOO9usOjnt5rF7wPfSzY7sdFrg0y8LjBgYQ5PXQs/ixFv3cfiMwcKukQN
UZc9ZdStgyP9KFllJhhDZpbjKTAiHUUzcrndledOqX7GHvE4/Fvr6xIz1xQ1clwW
xq+qDCofAdtwemCdd1jRoxSGr6BIbPG2tAa/E9fSS8upTK6qiXIBr+4a635fqeJG
0xvESqTYIJwocE7DwCCuNyyyskqaKePd1Le8ccuewE1XP770IjOWXl6VvqaADQ2b
23bguKyadAMf1GjNzOfuf+q/r1hkexWIj+qk4dU1N66CorbdQK9VF5Yab5hHV2Xb
RkfQqgRXW/t72t/pEVXDMIMfdHOf5p4EOIal387pW6DPkK1YE7vjwstPCQ1B4Hjk
kzLW5InVCq15Fktvw+O2lAHihul4Bed62m1QAyRiFGBUKapuTD2H+WebQjHp13NW
2QtO7dJmU5F7IGcHXHDdO+f76VczVSOxjgcJPYiD30Tez4lDoL1fNni0Ohe77SvA
RiDiJj/81b+E3lC8V9Ni7a4bgUYoGGPhehCzl/HgpP3DEIAK4HgnIHnkdtcrREd5
wpgn66H9z0ituH5K07G5OIp2mKkhD6wyrJZj+77VsYn/Nh4iyRhxFUfl4p4dNfWG
uqbXV2Mt1C5pnVF9U2pm0hzh/C5FASiumXNMrlhDb5brZCGMV0XMdvqHaa7xk/8c
CGp6Bi/Q1bvX98HQUhRcj5gPNGc3bx3ZlmVB0E3FeuTABX49Dw1xiOVubethaaDY
EziyHRXqRcjXvF1EHm196Mg/TPueGWftmGGe/KNkVafVzQ1G3c95YnFNK8Kc6CJN
SuMs7oXvinS6CX73ApUVa1JoPmeTImoJ5rcbnWrIA/lEC4ExIOnkwIZjNOSP7MAz
3vaaN7I0KLGatdIrLCTGb9OVHeiAo4DWAI+tdnjZrcuEJzmkR3PhjMxpEsmnLv34
J+iFdSozYs9vUVT5sn/bRyD8Y9R+7HMqnirtvXGOT8xokijzKAZP4hDYz07DFJGY
B6GiAcgoXAFoUuRpcK7mIK5U8KXL72oKfFP8MD+ieRYPE1d6r3V1dKHrd0X6zbD/
ekmYzZnoHLjVmkLaEyIfEvKN66SgwIeB5qBbeU+05qZgXDOjx9te76EPP3Oj7Yvv
PbrbrLcKRnVcBdGBz9XIXOkDRwcUAoT3gpOhLFbvMk7OA1SpfgE4qQa1I0jer7Xa
r7xb1ySbyV3bg6ooiyhV2pl1Z/AJY5wVTh6xUHdv82d85o+UJ5HhmjxPsoKJVqAe
pFnnPEIOR6jMSD/HaxxFi5JXUxEsATbho4LkW7wt0zSH0poZz8HedgVHTts6nX3j
apmtg+Go5vklqWLlwn3o56VoH23mEDAehQtx00vdnM4zVNHcH0deaJu+Z+TQCanq
uHvVQCNOuMH29meXLPskns+sYTzjj0CGalm8rn4vKZkoPZ3RZcWpjhdSK4/nGG7x
gY66NiBIjkDOMjNsluCTI2xz5fUdLY2w3GJqGpnFK4JxkBA2yoa5Szm0QU4ogRUz
rMMJ8Em1A9sqXas6Rg5qRSE9AKCbQ7gN9SYyaIG8BtjOkXNqopDpUHjIiQAvJyWW
NFlA1n+OU9mJUY2TXMCBoNXK7zNfbmvige17aQF1N5H5w2u4rRsKTDTVXzDEbof0
ICEJ0fZ3UAE365oD+1qGj8E9LyU1bkCyv5v9/vpe6r9nMuFjgNpT81Gu6E4Jfuo8
fJBQGGvnCg3nnBW90j44RTQDDqggXcQTmwJRKptchMP/vqEbSIig6vnxp23odEDb
Cr3GYhYVs8v4IGviVEgmPxjaX/+Z55jGvMAY8DrOEvpNJZ9N1Y7fChWXGzPLmsu0
TUMj/8Cv2vM18G5cHgNWWXxkLT++y9IRgTNmiXAPIe0zDvZRMX/OBAU0m1GycTeP
prATZcMAq2wgz+grm3PadVrrmioypDRfVewFp29L/IBQ/dxcpiJueZ6MtANQ0NMe
IoUcKGdGHhvc0Hy+6SXZIuZtl0+iqnhOYjrtQnrIS3sq7b7GubOzswjIKSen1ftN
IBV7ctFu+eXIyTGyxI/NWqLpgeFwUi68u9duuB7O2L17xEFoHqXnSYVPrhfinNCR
MwsYUjWrivV8iRHP/YC1MtTVnTABCA5FFAL+p/KoPg9U071Aef2T93aaxIfqWtCE
xXpWG/Iz7V1eT3obzcMWoKJMp7VIVgse9w0mJPnRsI3CA6MGPChotkwCU9ex9Uks
54uKLMxLwmiHOCIxw5Of+dmP00Egcyzu8gteZr30XrsSTbrItzNxXATUwRZKB6hZ
7/FhsOIrTnZp2mb8pgAapzPj7q9YglHi64bTKtAGijBOivVbLDClN3f4trzVR9LU
JUVqFmPoSFOMr8b6OqsJtsVShZh5H5c9BMEUogi/CbF6/t1YS9CI6xeQqs9j4FKa
49Nl+1aTv1xyvC3pcsLPxVl/ZFdQ71D73D5zcZy6OBWLQu3Z8V4Y9ZbhKZuClmJr
vPzTaPqEVJWuQtN2XNDCX1TYsUBZLOXL1x7+taHGcIWI/rcEhArOmPSUhF6yjQWo
yPcyH3St5/SYAYYoNF11c/MEHC9bu1ooO0XWaZ9Wn98rL4elC/JcpfaJwk535/sG
iS4B+yi0lJ2HcdmgCvXUlYnA/splDto7Rj+buX0AXY68lGlx7gLGne4bhfGTFdaG
em0BDqQfaUwzWkulvWerOSnAS1izn05G5VEbY8xkQF8U26UlnveMGjlTd8uq6Nar
H+lnayzgXSgSEJRxX6Bp1u84m8C3xeYTgybABZhvWCT0DAUfn+63T9+LHuoi79gP
zKmjdTCbKqQGmFtkaJeaUaEOhXMQVD/Fbrs3ZwWwqpOEnXQ+1aqUyJ5epvXOdkvF
3qF/w3If6+auuHbAXuUJI34MuT31B1O+B8cDEbXFPlgmXI0kOB7prRt4MiWbqENQ
uDTNnjR3TmHg1HiR/jUStxkT7iSjMc+sLT1gqkupHQJZG/q0c3Bn7102Efmmgbxe
WeqfXZGCrQcU7dqxyWxvrX9FBHoGzYl1OVfSeCNMkLs/m7TQCzWjxDrEAeZO1xCn
F7i92elud/bHVGSwh0bcpAgkJOJeKZfIIHAhP1uHJ7vgZoNwAwyzRgtoMhtBrY1X
JrXhPX5DXitB2C5CyR5HmqmUbyzU/pyi/xZoveRkIiq2Aa+jR5L8EJQ0xPkvX+pR
g/x6tm1gnIcdQ/Bf3t+3ne4qZZcUctRQO8BbGVDqHezq8eEVjS1UfmLN3svrYVxW
3JYTgLxnLAYHj7bWwP6P5xZyklLbC/vTOyJhjS2Tn7s1hlE83yaTn9GeA+kKpgys
06vW1j/VzMUheQbT6vZVYwapBZJJF8UroCkWuXeKvaNxBbSPh14k7cVoxUoehiCE
xWl3yb2vJgdq4VqwoKQZ4CFZulAlLNUuJyjvUr69V1+YULQVvQSJcxm9l9TIh2+b
h+iRr9rLvYILiqKYIr4+tuO+aDegOpOstgRe+vaG/EKR8dBeIC5+A2EV9o9gBsfa
yIJpVkb9NsTIt3HY/4p5wwCFsu3TmDTpsu5zZzGxHBXuSG6hMjcYGQz9zWi0yAdh
nL2Ko8h0aXiMhc3TidQ6I2hWb11AOI8SSeH8n4//+V+Uect1U4cLn0SPMCY3dD3t
GC+mTakfAFoEK4hSU7Ef4Gjj1Yxq9nN82KJI90xAZj/nWCJp+iJsmsiXYLe3qcAU
Gvi5P1HZ0rpKbYe6S+ULh/F13KiS3g8YL9sdouLdTaFgqnfoY5BBcrl/MNNyLgYZ
NXh4R4hge9Ysrow4crgYnmp/uT9SBxDlO5w3kBcLNbhwYVmWzcBjn26oLXCJSI6g
1fLuddpc1KTYi5Jq7s8U/q3O/yNBiSl2eEPybXapsqanewkZBQE/xssr+IO52v8R
bqF7vSvHoywilAP4Nsa031uYO83p8BcBt31mU8emg0tUy5rjeN1D0m4FAKzhQQHJ
AXE3ETZgcHRNSzGqUUVKx8I5NdrHjRPLZrRwzGOdpObvd3wzZBLOoaT/Wfp2xGNr
O2xF/VyWY1h5BVIZCN3qfgwD/DGJ62zD81ZbHhas5hiTZiEtJs55nqE3TYRTXbfb
o6HeR/as5ou4wlOQ9/zBwA7zStNOmsJtCDJtNymMeZjNPRVJzvb7SCE9XaYBy7+F
nyTE+aC10Ny1lh8JO2xhQaNZJEJ4ct6Dma8LBnao9Mt4u8LeRfeUb7wpQUGO7ieT
Q1mV5DejNgSeuADrSMOekSA25PPHt70elwQYN4B4b0YbjAMe8cSSDFCsh+upTVUL
eLz9gJFf93aGsHB2Wy4jqwHn82uLjr9o1Z30k0QXYjP+JHJtEhHzuMA59XBQ7WVI
OPmaFMNMP38tbXXEjSfsE1tmJMDJPYCud2yTu3NKuKWCmASUxG9zpvQzoEljntt5
N5gM+tJvVq8Z0IUrj6Ra82MjPD4B7N8T9WOeld99EWUsl+mwluUkhCcUZYDtG+F1
akJGx+2x1gRHfZ7hZixWe5qtBmTi0BTy4Te3AunYUV+SgjbXRqg+v98ZkgoLYKwK
8bvv5PqeecsOIh/1Z05WSOiIrNBH1av5SSO5F5EVrtYZhzdb0N3S7KCNy6N0V9E+
3xnd/Sr0bB1XsJ2JzO43tI5GKTe7ATkIHf/NcIhCaszG+lcKDgFOkO8fWISW/TdW
I6jVkW55113Mo5yyM9azD1bW+YWNMQgjwAsYyl+1QhbzdHCPywl144sEFow+3teR
dG8bbeYyqylKx/A6ucq5HKx6I+6on55prQ/WTbRaWeiJSpQTuvueHF3RP0XJZ0no
DpqDdTfTvv26NDZZRsHzpiCIcov58TXfU/i4IrVhAla/B5uY5zlolciS2yxFojo1
GzEeXXWuyMrYjULTO2Bpfi6iAgmwS2UvrrZjVoR+lj1KVElvYuPXeRZkypWLLej2
sxVWTMnhEqFnFuTn6gBNUnAeRDh7RAx6iA2zmYF2m3OcmPVjUqDit0uV3lfL4zr4
vzeCWI52hqt+wkZHOSDN+b3WxSxRnNKoTJbfPf75Dzd1duvPIrsIqwzIH6CHNOfd
01tr1W88ZFIzu4O2VvNMWTlhSOokckdtCsID5uS7RKtiBgdwncRoauHUzUvBGUzJ
wZEMs93OOqyQXnQZRUU6LC/4cO49zHOPrR6Cq6KjpzqsmEomLUIalftb7+89FttJ
muSwAyrikVxSyHoJGIJajspot4FjSdqy3Iejf57p+Lz3ip79DeSFkp1w4FVdoKmd
h+QctGBAy8nikzgDlfK7qw7iYfbO7RGtm4zifaMb9qoYD5mfnfjv2Z+iwTonfe5l
HxhNoiGNf/QOm+wkli2K440/n5awae1EyQwtjHJhBtnnkOnFBXJ+JBU72KSMb4uv
OUU2btvQZxQ5cEfw/jw1DUkIfKWSj4BbmxNgA2y/r/wSpdSC1DG9eI4msReLNvkZ
yFGRA6EsP9bYGczZ7NS1tnuaxeEGRH0QjSjNmAhF9xWDP4a7hBIZ8ZKMbv22DbdD
++O2g2Tr8lagASHktV9BC2PXVHyUXk8CWHxWTvM//LMrHdmDiUCo32SxvDTBbxqa
cNKGVam5zExgIhA+HBPO0E25Le1qw3oamJ028l6rzutXaTc1MwUtaaj2KhqLpgtD
kFfRhNCctF4QILPDcQhTauRcWMxz7WUyGbORFvM+5UrkBWG1zvuvvHjMWlGRR7Nn
rchqdTI5cIk6qWcWDMrQt+B5+zmlT/l4o/dLeLv30Svb8ihhh3Yh9ExqAjztcFaJ
T3yxt1FuwJqFFXD8EgWPWleFsnI0FDuKNdYrcYGhrABx6hY+cCiaqAQx6gvAbjKR
fCR6inqbh9yPXNOFchL+wALTf1IO16nweRschyqGnwG1aVdxBuavJue1ejVjET0P
42QRYuLvQkw6XXL6xDJl7dKQCacaYO1fsa7iTYRYsv730434unHIsM3zGtH5xGPr
j36YKe10LYNA7k6dGDqUJ6SdXse+B2rwiG0i6/qat7Ix3pAe+SxmXUnVgVVeZU8m
OxeoKi6agAz3BioUi1jKmFvLskGZ68ZSuNGrv8bkYsbeoQFVl8Z3DoASM4Ia+0YO
33s2DJB7GGPhQQG/kdsbmSwbuqdpS8KJFtRcpilGFRBLCjrptZqqXq0ZzL79//E/
46CjEdBLRhG8PH5IBBnD8DFJhcuLLLfQ4xtBCbPvp0cZB7GZQsY/i5MXmFOGVEzj
1U6xbHdRcQ50LiiXv/eB02hKS9kfFmdntn0Awm/f2L3+xldB7vk9yLqJ3OcLSlBs
Oq7fySHQTBfQ40c5cLzplA8NyJsFygYtxpTdJ5+NiKKQU2/XaAjbCXNoev5SV2FE
H1mATrn4hKuoj3RGEFilW3JnnaRPcWoY7K8J6lwdJnIu9HlLv/7HJ8rjYj0JiYpJ
Wh3MIiDUC94tKjVMIiwxf3rys7gqpxTaSNUqPcyGIEKznegPiTtndVWyPLPY//UY
rp1Zb+jALXq9YwCKeZGyJHRSNiqNrU4Ma3VYS0ZvNyoOtQhONI89AwUyXWirdokN
ELQy3D47Z2zcsig1mKa4SZZ6pgRKIi7bQDcc3C85APA0hFY5pwmOPl8wIuKhZOE/
DlFZMYesUeleYdq48fc25SQppB+iOcPeFro/2q9f/Jiz34Jhix+cyyWWbm1rUN1B
v2Rh3+2hwT3z57kpamzgjkNWByPPQCTIYmGR3kujvRbayjiocJkmAkVtvFq52xcB
B2/d2wS7WRbiHy9DxsbJOAv847kieJZH0b101H79OkkSIAYNu3UWHyHV851qG8pP
6fhgbeakz2vhkjUyDvv5UxoR2xSxHOPbEp7Baec41h3n9CRhGv8YaYPJC/6JLVRd
hBJtebmdzl5m4qvffJy8e5KDkWGVIgOz4cv27cnblW9kGwMdWCF+8jh7IdU81u+i
wD+rVvguT/iIo+Wsc52cWQMnE/ljbjuMD5JRxjMCTx5+GoamXTk3DGI9mB1y7ciP
tJTxKkaIOw0VpXI3STdpLOejqI76mtwR7+s2kgP3mF0aEPo8XMazxiv4sKSMS/3y
ibINQR4rNcjEcSUhCUTOH0VpMSs7h4bRsFuN6QRm6BcSWSstpQkDYENWT9EJQIYZ
QIK+nqEbiI/CeJ7Qkh8I+z5yxB/c9ZQpFFLZDbwSqIED82bATRB+MJy5fQUzwIW6
fBmolF9CDwGaS53GbF6keC5gm5l6FIbU6Oy2wK1TuZGJDBaTdy5EIeK28cq4mm+O
TNBJeXwK9qQX27MjFWospJgZFTj92G0EJD69CXIP13cyOEhRbwpLBSylfjn8ee1k
agzsjSJ7bOSdER6KXmrwD6/asIkWqQEyb/bf/j84QeHtl0e2QM6QJ8CgyvAIcUfc
lOW+zcKE8C8cSWldHKMARbaeL3S8Vvva8wZvBhhRYSHc7oGi/vV3+dU1UkgRcoyT
n1/ASpGQBrWVhzDIqRl6XYxpmatM7FRdis/dMjYAqSLa+9+AhFfHtd4D24hhETlC
t37usPTiFP0xRKxpaoTapq8eeGM8a9HUbU8eKG1T7SzPXeMDUJsZf0v3bKvslqzy
c8RGYoWR+2yV66uJoGUjXNjYirpR9JRlI+zCzdaFYkE8ew0oCr3yI3dDro2Hpmif
VNNpkCrWA7jf8kXlT1YMvS4oAYTQjy3D7XrESwhxsAtmjfhAhuoBysDL8fLbOe3o
hcHpRCzDCc2G6l0shEMO30vJYiiNyDiEvlx2lXkIVfjTe6J33fKyd/+97PHilw5S
NbNH5r13e4nximhADhYcvdjOcwvbHTas5hu4mhshI6RESO9QbQPXLaxdlBo/Z4wT
nonmqeXx92HrLK1XP0j8aoMWDLw2AkuN0D50L7ReswxWFWBCcpQrbw9F5TMhSMWm
QQLYgx+Z340qnJTOTH1zcPeZ9QW8HCPaCvgSdREvQZbJNDFNXwxF/dRV0gnP4DqC
b8sIjMmp4E0U7/9yhdvo2dgEusczd2vG+PzbT9mEadbmWo+MZjFhhDPvRYjbCl+m
WrMQrnQJiZcN2xYuDMDtNtPtM4cd1rOtc3AyGuIELlT8okBlNixQCbmi+k04INfb
2nvF9G0JHHp47ALtXRt9KZnmU9qA1BWsZ520e1UlOf+6RINhRGOeaPSEylM7E+J1
fJwtVTZeIxOHdco9O3lyyaLbU3KMAYGNinGt+7iyXSt9FjR7H8qMXiTpjju7TLGc
kE3EE2rrLCYLQJhl1W+7BYbshmQaKKf9h+vQmHfJLLwq0JwbIXe8l1zaIYNuqUWW
EVsEMP2M01sokl6xEI36cEvgVcwVaJev9rC+cN2oRsr9z8l9nhIyZT/PAw7f4U0T
3PovDZL6wUyfePLAl3GrgnYyUlDXNdymWJez4CIcJmbJg/Z2PVcpEjnJglpDhqxw
Dtko9qfRPNAfWjLoPsSYZO4RPb1OqzYUIM2zcpB6ZBibg+WXDADd26vzA1sH5iT6
0YJtvJTIiRHXVv/IU/G+wCjAqOomQB/vxooiPoVp+qcOzRaZDLPHVlI/pFcNnGIC
5X5PImCPOWcPgtvBA0Gay4QLXTGebKL24nfMhmxVopWxdvVih1TBk3X8D4ZrLiOJ
Mp0VSJ7nOk8XrXyyPyGT5pATyZBgMKI9UXehDaH36A6yp9eSnjd9i/B2Zy9x7Ejp
ibNwUgtbRMAuDrxZ1gHUb+UUaLxb8hyc6jg0DZ1QUEqbYrkVxCdvpZ8gFWDwAin/
zB4WothaSlm0I/5ytnuZhBF+g4lZsFIy4JHizENR6QoT6LhfNdNHrwbJgkmD4Suy
r4rxKNMTYqDUOZIAr8Z7GHI0Y183dsrYHw1Tbhh1RLEvvuOD57AdooVfUDZVDZwr
1Nm2exaX0AhkP0JOHsEMaMpgvkFkuL5RzKVAtXiI/kjqXgEjTn+lIcYkzwhvD+tl
1AJ3E0TKVDOdDXK0YiSM5JsoElDD3vZavWhno31NHXC7COTWPrmhfEMXa7ZJMiXP
XhN0mzOIu8alo6MRSJjcKgWlEsSErxNfVAwxplgPthcazM+eqqcjkJIbk8swPx6z
FOG3F9f+mXcb0rhsQxrPEN0m7c4LW7K8xAprggqJnmRBHsS0ZKFA2SGK/6e5aaDt
K5MTFDjApB3H1kEQkalk2lmXb0SLbpCPhBVI5ReuaSOE8C5/Um0WsvpaBs6XwjBE
xq7ekTPoAmKPwiE76ST/0gkTTxyC8cwZkKqJKuCm+U70R6NRNLadFskE2trVuKxV
BRt1nRM0XQ8n4/B8dZSfJ592Q3hrYEb1heNQ6wX7ARrufl0+90HefGaZYULxrBw2
Ik3ghjZHLtAznkxXtWxKfIjUJGZ974r6oxcCqgv52BEtoMLnq9g5tOIrXh3Ojvp8
HMoWUZCrBua/1xKhjjip8ONH14iHu8XfTpjy4bH3OpoD+L7+sb2p3Nz9FJ4thA/C
XgRK8in2vBBQ+/v7swhuOt5ht3SIL2HEJzp6J069V+zaOD8135PB4HOivhYuoJG5
HEzS6TF94dPfhAyccibO6LueF4+CsduOrePhb8ZCkt6nqmXVqaqxQuCuNZlj/2dr
ZAl851vW0AIotgtUeukEIY/mxvF59K53rAobD3AEdF1KwQ6zzjFgF/+oeW1w1sSh
/P/Wq4dWTXg3kicAsB49Ug4yEu9KvjTppuqLMiEwM6Bm2bgpEBW9Oz9I2mwVl2bu
iuhc+d4+8WSINo022R8FisyEGKRLO/e/6aAIYKWcKu0FRARZPHrVOdAA1o+3KjQO
SdQvOcAdjPNW/0Lbqw1OkaIZFVnBDIeH2RtxbTF05rRL9SeBhIrKp1jplamxrhQz
pYbWsf8/NnSCEfTRsuKzsoUTqS7kSX6P4xxdYRi2J2mjiWUCXqKBbynPWK6mWg92
xiRGJhce9ztQENCJiQa9p0dx8CxvP5guIQO2+Uh0brNpBasr6qlKTZtTc4WKJxif
BLlhECHc40xww3zJ54JwjRX6GsTR2XdC+oZyJeJ/EVfX17JnuWeF5s3LfoMzdmss
gLFqGaWOODPqUsScrNoJggoFjFpMV96d6fbb/Aw216JmFByFRnqtEX1iOKGGz2Tv
F+34TOupxfg2PJlnV3c4DRHKoxpOiQGWCc3N2cCyeFWkmOIlEGGCr0s3n0OXxqV2
NJzuVzNU9kXcujqQdNRrzSKtLiv6/YR8sidMsI8ROdSaOBqvdb5wWNRtnX+jBLcg
HqQT97DRRrL7kgQUkbrMQt3B6oBvinBT/7cwqFnjM2jTvTcW9+0KuhXFqV93fT6N
IUmCUmBvr75jVCbVVR60yRdoF7du9GYt1TG91qVZCBqqLAHc74jB9p8XvQm8d0kx
iSNE+wK0JCntFuXXlHk2rSb9jWcLro0nu7NVGhe/hGUl08rQw8qkPqoOwzyA3Tu0
KrVHrdeSuYvg14u8I2QNKX/u297cR8MtbUis8cVzq05nMrqVi5gD6NQDt5+5JHNv
4LL8AhOG7vdHyBOPBGKUNAk0tc1Cukd/znIMoeD1Mi0tIKlhk1+GDo7/bUCMlYH2
6e9LV6IzUV6777j7giCUGf1x/S29touXBgr4geU2W69STa6TP+S0RUbioo0vvUu2
dLd+gEXz4uydypG8qETTGNCmgH3EUQg5MQwP9n2O/ZXBTpjT3dPwpkEHOUkqn+Br
qGGJxb4WTfjW+hcAxc26v3591MCNP14R0Tkz/TSt+C3ECvok4Fc+Y5FH37A10XaS
vz7x3WXkYF9YVK7rQr/Pm99xkVrHgppbnL7zI1u1QxSdQWuGm+oxIYsxr/2NfkIQ
vpE4Q97ZAVXLJgbN8+3/NkUsd/E9R+lvmTwEsmMNhCGZPh7aSC6JYAKymOwBZuOo
H1oqKrDuof7VH19asZnsuAU1yX7W6Ka0wD5UZzqB6RHI2UdpyQ3KMtlk7IkeDaFA
OBDEGEEZ7MdkbzWNrLG/p+yTEfaRVqX2D29cZ5c0sSpHK9xhGwucKnnPlt31sgCK
ouulRUeAyPaHNRtlcDEoqtyYGqEj8lAoqdj68+nc6wx5NQ+VjbrxtdLOzT4hqpWM
2fR1lXIsuaBEQv7/xHa0TV1ik6SJuXfKVRlYU3vUjXnd/8A67uPF9avhOeefq4ir
VDgW8cWs9/he4ml+RjNOzpJK2eAex+xkzX3l3LFtAqnSgVfNKF90kDIJxdfnSxov
f85xR6RH9naZfE+3h7Jjb2bmVuoJ5NwVweBq2gikCavCT8QSNcYt0tJU9DmlNmy/
V67bR1t0TpRYj/2JHKl+WZxc4VAtYzeoAa/KLM8CuUmLKMIzY6wBC+8TeDB5rVQK
hfJSdSE4TjTg656z9Zn4/+Rqg6dj3E+ygHyumvVarzqO9OVYy6KQ4mLA95RzSABZ
/vWf/iwStucic0vjNy1HyMIKnSgHWmedb6BAr7Zw4cCeNmvc67dFVY0JXX+Wqj+x
miceEqbJz5kPbeOCXgzs+XI2HVrSHTcm9P+7X7xLqRgtBXKUIPkFxJ8slkZuLPV1
jmJ2gE7q5N+ZznG78tQXQ0k5qRXpO7a24L+7v7T/WtHFLhP4AhZW+g/71V691LIz
DLIaR8G8/fBXmej1EgcUPD+PIcrXSDGMzh86tWBeQclyXoTFCz20eUSKV6raACtK
hRibAKzJSKKjOIS9Pc53Rx5rMCoVN5KljFst5WSFS6fhJ95d4gFOi2i7+PLL9cTI
8t09TUzeiqyOH0OtPUA2G6gN2CmrRf5s8/X0iGg0wJI524VmYGo2EXO1lBzDwKLU
7qeOVpDAA69gMjnz0TldW5nhXUhWOB8I5K4uBH7fyn32fn5x78Ey4X/JssPM2w8z
ABNdSV4TOAximNLxXWf6hEp9Pi3oBIAH0bD94amNobAh47HL0eOuMOVAaL/DChuW
ulUGEtTtx74GRCwfuKs1vBrccHi4511rW/0sgGLDws0gTBlzMIqp6RrV++0elfRf
SLla+P+7E7p1BY+LNkqeOh6e0IhefW5v5/W/QIrzNAi+ekXvXdUookhW08exIvqL
Y5bi9awLDrxSdYB+CpkX8nsBydZQjmt/FEwqLpAVMYuTOEsq1Nf3uiN4S8lLdlyr
E8v8iz67JT3Gp1GJxMfYYBhI3Ht20Go1p/kA1XU/eim4cLvU9SRaN4qSEwReOB2A
lpdFm1Izs15BXuUVO042mLsNyujpe7LjJHcJMoXfA1ye2jxi1J5TljmOk94s57AL
relE/yLN3kM3LNvGW70LwzrQ1UFVRYgpHi2CeROHjq9vOjgZQDv6Ej3zaOB6hHSk
fzEUaNUqlOmMZMSFHUeK3o4ryxcV8ZIilefOWwgN+OhFz+EiIGlEFs6XwYj8vTAE
6bjnXfYE3o5iEFWNYdc5Eytn9YGoXKMg9UC56qP1BpLIRFiKgA2IRaCp/CB6Fdt9
C4usz1MkMW42EO/IsksrZGN+Gm01eWWxL9kxayy23dqUfE3CZMJqOHl6QjT6MldW
utayxV2GFaRNFc25S0qYII7G/OZcNrP10MwyFYEvD3hSXabGpMR+I2EdmAKZGGik
RS8NpHgvfinVvYGq8aAzqfOERuZsVhyt1lZNSw4rSLN2p1U+wRk8Id4fwktEAP+e
Dt/LHNKQt08PH9MkYFpTt+GZvgurUbLmxsk7LV3X4GdDWZw34BoRR5uJR1l75coa
QEWdrr4U3izMdBckJmdl7oBBAokZSiLLzVNLH2GSL89tAIJn+Prg5hHv3T4FBWl6
uJ4gxUKCPYw/vEtKQdTCeNWUOC612R88AZagbHwl/nXhekJnWbJy3brH2F8YcjDT
0+yvmCeuuuUlSpH1GFzTQEGxfRoKvsHqG4oAHJaYEKM1cFr5vbpfk1X3CBwrIkk0
DAdze+WyCsPdtII9yyHo2ahVvX2e22W2LXzTdM6aq2HdchJM19KEo2MCz/SW/BZw
MK4dXDGjsj9Qlo92Rt24sRPstZ4VAQ4pfp1KP7tGPqouOKIo9S0g7xql5nHuGvd2
6HgDSlvJla50gRXwuVIL6NCgezntBhkJ9VHfVbNIGFicv3cqnqFdAOWkpMzRuQ4K
R2NOj4coyk1aL1qsbSy7dCZrci3Gtu/osAYlDqtl9AZ5zf10PvGuo59KWHasP5FE
OHzLrUyQmDbH1FmFYsOflrNu7TG87y2W/84ydqw9MiPAPEnEvWrpdD6A6tQ0sWNH
cbl5R1Y8OKUFRj7KaIc/x9sMVwPRIII9HJisctZZ3HLeBXuWAI9N//JyHwD0lq9T
USSbkzs++xg94c33Qo3JVjMOvrCBvqlJ3TXx9Lze4pUJcvwhxykfUbUDW9KA2C46
og6z1bj4VD/xwDpac3e+riijjOGuIWC2jitncrKxSTjX8fX6P0pc/rXj79xsD5PJ
GqtThFk1y/o8KUcbfb02IjdnX8B/JEuR3RmKgPbIFwxMZkN/OIWXgSI1VixMPe0p
DRzwmUNbcY0WTDiJjdCXW6u0JeQnCaeVokWPZYSreR8d8ZKmD1EK3bP3tmdvEosY
VXyNtSaKnfg/w/QB0pSqn2We7H0BLeH2n0NxpJkMRhedTGaYIoIToTcQo5bQSAzn
7YulRlnuwz3Qnp2uUGEtv2OYRx5UHWJwTiqf2sfQVmt2wLf1PcMypjUT3sNVmTXy
KJAAGeS8KEctCHhYUqYK0Y/eN+RxjRaWHOnnVzY/11JSPHs2uhRR/CLHyoc+IiOs
vfLtd+ffXr7ODqEl4m2VTGIMA9XUSSkfQztOLEwtOXcpWvMrhUunMM6aoArDwbyF
TNxppQWNPMcgXB4BaY5XqISoYQEUf6eRsj4aBCmBSepKkUN4juEbU2IzpE7CsvUV
xKhyOfUL6OHJBycj8qiPQ7wglfCFf4DWIlwcqd+N3evV0TGt7CFLzQ4fzyBS8Nt5
dFKt+kyyiZnaRLkSyeOwGQQ//G50xhp4+7CuxYOxzNf1dxN3a9tSpmml/BiH11ga
M6OQ8Oq+oREyR0OY8NNm95nrMYbVlerzrXIAP2ADLRnNVKY7bRLxb5TLmzuXC8H0
ElGCECpJK6AmAD1nctlqwmR/NZk9jt+D6Z8qsdXrf3UoZWANwMwcL+DOHuMFWnbg
RHAP1TNbAqDcR8Otlxqq55esVPzINy+8wklah6Q5/YwMRtiDgh2TeDT/evIE3hEa
rf8a9Jjyr0jYRWSN0pyuqkCcCB8Fgu9ApPAvfYJWXfrd0x+rd4cBiakvh7nevAln
eqDpouBrm9LB04eqdqfpRNMQaLdoP5hCjNPf6aXiEs6lBkl05AQY955ctjJH9HNV
LSPwlk31YMgZOuTObp03yGWnA9Ep3nJsslePsPQxNp4Bs6c7l+yapQsmuNK4dBnP
ieaCI+P3CD+a9E6Afd4FkOx//WJFgLWQwp7ezOvfeJQnaekevmW2kKNyKDe3rMP1
pBn9tzCz9vgkmB7DaA46FGyAG/h8ayzAO+K/fvvCYlIAIsdiVhVrTrE3XMWvg4uB
jpac5AZTVpkrV5sR5MC+s7Hbtu1F+i58pxtw77aNlxNVnmduXx2E6Qc+kjrMGtvC
nL5cWcawGLnJLiizpXF8f7+NXZYOowJpBg2clwHH8jVHe2CzG6Fs+3Zh2dKP+b42
NVdiogYf33NUtw1IT4L54EZV6K8VF10xlPVPc59zfxgeYkf17dq9+DESUGFwL7Jz
C7aUaxI2lunUVoIsRKmOU5b+Mkc0kKrsBM7FXbQaqLHSVLe+FHTMwPJE1JbUDAf1
9Pjl65lr9WSjIzWDltWtrf2Q60ig2QUPUmpEeWTE/gK06pD1wic1fPpqwTlMWdrF
+APlo52o6svbyXRH8p+h5X51GfF8jcwZ0M5CeDKgstgQHiV1vV65GQ1zzD7Lzcks
A1E+YsUVC/5qdFBL1H/ON45r4sBWFaKYlUy81/dPnSBhftNUDaYptNOZRgBdD6FT
pjQiG+/OmZor9ZF/TFUSUM+Ldo1vaxvLUIA7A5HfWbrTd9m2SKygEYAs7wbQaYDp
iqrkrE1Rllut3rHOt0U6y3KSHqjb6ZLQk0bJRjiPE8GgdUtFzSsrrAyYKFugsH3k
RAHu+LLeKvn/Fg6P90joC6uY0J6BIG+6jO3XA4sbKHcaf6Bg2Uxkh5Vgaij3/i4h
LKM8JEl8vNQnulnoYKjK78XQHz8KBrhzdy+7AF24Em7j3R4yedWyrkjHeBJABVjq
kfoK8uP0Wf+sVDUnjp8cvEeHuTY6SRTvUMMbYL120SSCOblmzir0FAcOyy1Gbj3N
4sScDTXVdtFcA0QXyJtbplspYEEqEozsSGVNEkZ9vE4L3WB3Is9gdk9xEXdBE0S0
8+RKYqvPp4Z+RMnjsxfEUISv9wtdDmm9rIuUARuBIPLBEaW1DgEVaNsVgPVta5lW
enBroSra2N2rjRL18ArC/+xCzRRmq2UP7QAXWOR3JuEc4cpeeDW/w6XXw2oQImrQ
ZadHzhojJslLmIDzFKatyXUoDmE9BtfYLUnsNWJZ7vRWWhV3WK3RaynOBgjM5hfA
qDKGbbW0GLY/JjeSe4pVNWcYz0LqxXzL8WxeuRyRdWD6/mLHdU3QcwG3bMyz2LSk
CXJBoxk+wdKm7qgXyeXqGXG3RyrJFBMI45eTtL7yev1WTKMQgAmr/EDtIvibaw4t
JGARTTYxu9NMoRc6FQxGXb0Mo01XYYYL2JydpQBRy1cosfn55XbPicgKI57uBi9g
yqhnbRvQk4BK8lUlFZJCRXK5GCg7UVize1wWUtrRxFVJry+82MQ5hnkcwfNykEFi
c+3B4xnn15ED8V3WlM9eLm1JNk1ElYtH5J77fXtVXkReI/OJ6grNJ/GwYkkzHElz
Nxk4zilkBggRdMLHEDK29O9TDq992k/W1X8ww8MnBg8O6CNAZVXxNqzkZjX5ZPw2
8FmmQeJGmj91WuOez6Kc9v5S8RqLNX2NJk7ma6gUy6HeCV0ZVE+XpnQl2Pn7aGt+
cLDy2X86Qvzr+0gTzUsHHxpLiwfZ2VOFswYo0f5SuLPA6rEUrKSnnH219ck7SqYE
UMVGxG5d0H/Zt7d3404kY18Y0rL1Yfw8ABx310JajSeHE/gU2k8LXjPhitfVvzRA
PsLlYBr4gqD/xLQZ3yLWFXVTtDx1wm+/d1xnL8IN7viGDpeQ2noDULJ2hpUV79H9
aIRQ0T8iLFw74zsPtTbNLbS8SMnUEf5/igmXDdDVrJihnMbddGSn8pT/R9nufbIL
jo0PqsHDGCAchvkQW+H5BDKW5YM7oikHbJWIO4yVMtOCg1HpGMcMs1ad5ekihGTd
dyRTJDawZGccxSCC8XcenT6LbAVM4kuHupR9S2raCnxNxVA0i/TDAJee1KI8FebV
BW6kXTrHswt6cc09kcHjuIc7nDgekYdeHQvP6foqSFQG6B78WCQPAUipXWXHP0J1
pzVICyViJ31tMvEhw5RuxccSayntEpnIOAXiAMod0hhKJhVm3hISCQPes0rsNT1z
1fkwEkVOi29XamOwDktgROKDpUJ1wHWcqcSHULTSvRR+nd8LR+xpsVKavhjEXb/K
AQpoELpQ7lA4UmOboRSMhHhalRitXC9nC12YifLsCL4ukZidHBmoRddXbR6JNiDc
58VI4UIRbmX+eDJewU6vFKW2t/SanecPjAEczm1yzhGXv+9a9b5IRqlHDTsNVlIn
xo+irpSR7UPvj3/rTwxOtIiYAzHiKzh/86BJAdyQGp2IH+lgZfDQ452hPNUt78Gj
dJuVc3P60tFTBPTucsEPazYJMHBRfolL36+NoDirWHxMQth1wDhtBPkGJ8y8Z8Dd
JAJ1B9oYh0Sg95j9P5sClOAVEsXx7jatyGTDL8mzFqa098IHz4AN7gliC5PW2HP1
DxtE8j2QKop0wgjv1VamTCajtqwFvYUOUDeSFBw5ovLwxdudBPJuAsvOuwWpd9+H
T9V779N7HAvNwb66yIQldNtjqvMNHqSjog2RKPEuX1VeJfikfIRTka/tDIYITrC0
eNCuq5Rf6vsCHamrWWzvxLqDE0PST33oVCnnqWsYo3ytrNVDD6rzUdMwBm9yub6p
IbE+wSBg6tgVcYq3VPshfZ9jzBWOMoqlKf3AEBf3KD+G0QPWxqQ2Gkg4IGKtFFl+
/FMb60FXSZjc5iuqsK0sFybbi1sPBVoZNqlvZPt8kSUO7MfvP5BpNIRDhPfhkRB9
uO5B2eAX0xL+m5kKBZy3Bh/WtSpDns4j1ByDewc5HX+rQ9Dyu/4AK5zrxIerc2al
hZDNo+z4yz6r2JQwfnSvy81K7OlAC7sLBJsnjOHCtn7Li72GGkuT3C/2T7T67Z6d
J/wIRiw3Jql3M+KvHnbdV/HeKroHax6v8Y8x41C6xgFUlF7ZOOwlHtS5PvCKrIeo
fFyHPfW0GrQ0lANJ9jZ3TgOtlBFnITpnt5nvip0Wv5As3dn67BntRs9vRNlFX2ds
Mx4jGx2ggdDMaimlTOB0Fn4WSA0cnW+oWPKjekCexMi5yajxoZGEqnGZVxBH7jvY
imKi9E8muK98k8QJ0OWxc51LxLBoACW2N+Dj4wnAZOp4aeRTK8lH+GA2XxZVm0Ka
2+1sVFsLdnwAnQ3pLnb0xrlG2pDGOlA0EY/CqoRNU+dz/Lvya1u9RXmJ4hUbsb8H
5b3rx4p4OesFjeYIEVxTlZVZ+w6v4fvXMAJlKOcd1BZqnjeA4wE0Y8i7ScK83Fmf
5cFNhpREy7g1ZVctX6jRWSWfA5hPjn08TPXrjFt8RvQo3Vqwb9EW4IaA/NaX7Yaj
g7Rl/OHaVp9Ru8F3NnS/6Fh4v0HNLG7jDN870c+PDuF+v89c5SLcgaVFNVgVw+lU
hLGU2L+REKqqlgWKntUQYO4dWPE1TnNb+U2T9t1agyhhKUkn/urAUHbAtgMGXRR9
bq28TPOMfrWFgzrYVE972zBbv01ZzIJq/lqOU6vgZbc8by+WdtodqXXQvM0lV6G3
4kB5GupojIvKhe4MNFsiNpqvPG/UHR4gL9ek6Y99ireBUO59a1ISjoBLoEY+fjVg
jJh11v9qYPYoWB/1rDLNxw4XrOpVsHBBMHyz80jORO55rXPaKj9fh7VKttRtT7KS
+UqvZ6e5vA3fllWE321sk5bqgvLrVdGhbWDhyO3O8OfhBqXCWFf4+xJuFdxeuCUq
DKOWBTcJTdNkK+YAwU/FxM21tg/BzAhItEnx0EojbPdDBMo/06B8JkPzQaDp5Ayw
nJGAiyZt3/bS2ohqMQq2FrEqGQ/P+ROXE8O7Sm37iseR3r2VDEuy8nvypOUogiWd
ri+oY0YFau486jtSfSNc6uAxICKY4HTRjUf8ltAUA5SAYk2eYWBEe62cW1R5Ekmq
/EMBKp6xF1pzixJ/Sw9rhsurlfMNqtxPtF/CvxBUfH+rgrnWWrY/mA0IIqfJKErn
PGbAl7wBNCDUZhVDlqwE6w5fCHP0oepIE9KYheowduyRrW5NpsgHd3SLfOhBzVs3
r/lKtiSzvwUrEM76fr8J4ZSTVFf+t2ZrAHYyWx81EdVLKgnuUI6BLH7OKvOFagnG
Eq8VdWXUWBBfM5yx7zRB8L6w2BFuiUr0LTtAPj2EQ4A7g020Xwdhe/ZeworM3Do/
C6bcyNM4RcFTK1PhiYMi0G0on6WCoT40/nQLetRM2gAeiApJe8aXu0ubo9m96Lqa
kQq0U+NieR1u+1+HcRcU5XzKquuqZZVtUnw4yPMgleLqIv11c4/OjMsyVmxaTpS+
8sMT0zXM+Km9/F9t8FgKnRBsVLauTzBeSBdVwpmqNRKdot+7K0zk96cVbrl75rkb
xIqUbqimM5ihRGLT48MTBroviKijjBAzkMlEP9H/2FQxjf8XbSOB01XI/LWowwdc
W/MIKTf+ZLqjLJVVaxM+n4rlLXqq2yZzOfGbPBHqAQHfUUjrgASw2Ut88e61S5wp
10f0QY+AAQl6x2zd/w1qgELS2DBNDmfPIQWp6gNQOWM22qKVeIbeepiVGTOykfrc
OnFE4UA3x+VqvIPaESkX1AutydutdLcPFZHwldC9yFCcbCH8iC1a6NTs32xFqvxh
5uWK2fUB5hsEeB1I4Naecuf/otFu/vaiRt/Q3DL3gPM9UqWFjPfPQQ19itzSRKag
2ScOQomSUrfNpZTd7RhphNL+Vc0ep9tG3zTaHj6wfZA1uEq4QJKV8LjSpqL5KdDH
Bz58LjFPd/yydvB/U8bypuVZ4Qmt+6iPPlWtZxW6x0na02M3j59C21nOmoqMfc7W
VuJ61Lj93y64qdJ9J8gOl1bIZqHZFrhN99Xx5vNDFt/bP0dixp/JYjyad6Pi1qW7
2HBeXGGHHwHyVfGXnJPihTyN+8F6F2sXWWOYYv1kPlI8nV84VJ9/ANimnwnT8ICf
IMXoENUE/Z4UyKMs96W3KBwWeqcyPupf+gCd0gG9Op2E+QZI8dO6PBv7wy4V81cx
aUtCrmswAPyC+JV0bDveVekKnPgGWYWDWZywxkrnpemH9vz4eCQD2P5pWd9kP/Ho
Kf4/7qNgkgikaOzesm+GbMUjwy7jSCl8jbNVijUNwE6XrXc0OIffIGDJO5ern+nk
nclogzWZV/G0gvxe4j6D2WTIXIEw0drRwW0f5+MfML9QtKMpnRTVbHx88B27+MRI
o5cHTbKjqA1XM23BoLinTEs9XjJbpEELwYz2Hi8txNdDzK0FgsG7xJSNVA+SxgGF
nEdqcvuFWYfp1WcKmwzB8/1Iir1KAsCBiSe/CalsCIUKIXmp8f21OYlscQ0fIvcW
dbw/UvgSahJ5iVcjneqcXb+mR7vc2q7S2qEUrnBgtP725Fz22wmQBoQSVRrVdPLq
8GRaWkhntEfze2PTgQJU0HaK9V34wNdfO/hmOswgeLuyvIy7QSzQxfW4vNHIn8zV
iVtzquEiwrNgYS8Q3aLgcxUjGbkQw6Q5L6U7EgTFo7Vz87GUIqgjc8vd61UtbBKz
KeDLk5S9bWz3rPW5T5+fPsWWk3GnZlna18pNOouiPShg8lzT2p9smdYMLNk5jOyM
12bCcTY50pL00wcdb3ul8sU0SKnOw+etEH2gX/R976FFD5TbpLNbY8OuBEtrO+yW
5fT6bBuk4Te5h+L780h7qTSqIeWk/iukYf1tkS/PGUMgN5j/fAF1Iv+ijWZkl3Zz
DPdFxrcIoNxlihe8/tr+eIPA/Y/XmWlpoI6ddbK7KX2bjaBMMFrHt80sKITh0R9L
pG9PuU1YDl8gQcR3ZLn/kDDTtvNz9CTgQMJDb1MetUM6d6RkscWUc8W0/CuKcuHp
qciUD41ehBDO34oD1TOMApuNSM2/ubwmR1tBrCZg8PNOI9znP351kqP4Mrjjzwld
2dPd9w/CejlZXDLGUp1Y4yKlTa+D+uvDHldRQ3/EUyHf0Awy3oJ0nbpTaNRHCROo
wPJuIsaP/f+XRR1wQD9ResFpPfcnXrMaUxuMn09bj4l3BGOwFJGiNvawVTCDI7xo
78tD8zIpECnlP5JuVWs5NW71JtmvrvYjMde11DW0Mtv3SteayelsPXpRMNACmeLY
WBk0CFXvPPfdjGaIykOKr5PcaITNcLtkQsO9GdOFw5hUX663LdvH2EuLcdO6HPs3
ZEo4I+UqIEsiXAtgs6ftaP35Pka7LtcvV4H9Q/YeVzTgZaYTB+IRpbcYZ6AmFFh/
gqdLzsWKk3xl8NiISUA3EXatJP0HR4653uFatmBXGNvlm3+4qpy69gih8nvtjhd3
CNzZjPtOqmAYhFhM6x0qhAXHqfWL427qBt5G/K/3aU7Z0P2WrMhdH216PBalcLdj
1NKdBwb1APS+DMFYxFTioy59F7OM6T7AWbgm/Kzc6RejgVFklKqxnK0Hq9I5qtPt
ypJ6SY5p5qXrxQScYwfaPoQv+KCkp2o1IrO7Xun9rvfXkJcZeUKPcPksT1P0+T2N
o/cy5tzhGyxA0OgF4AYc0lliIzuzXsoqg5vD3xAZBvLhx0zlbt3eW4kKApX8i8ST
rnMjPtCG6lINlyGYVKnyHEEFR3DMhnthIqppkGkXTj0RrGpBzGBbWmxbWqqHFaYV
giLm3zA38OS8mWwOstGkyYHn3GIB9mjZgjHecV1mWxsAsAADjn6bfNj7pk3Vuthz
NFlF85r0adnhHgUw0H3r0QPR1tMO0iYL+jFC/9peK2qupORLdsA22Z2EDxpGA2ah
SIT9sjyScoznsTrnEuxAAleI8tCMWBuL9Kyy4t29E40HoRbN1Doh6lEOgnHV0Wa/
kJhzrmsP7W8Vbd+uwAXg8PYYQuAt1SjYgFWOMqtDLPtFSOSIMCo74dE6AZgQeiy/
OGkEymeo7AAjBj/tkP8rpRx4Ucg+EocX2k441N1biYaIiROsxlv6ba3Zk8bf5H8u
1a+DTEYbL/cE0OA/1NAJN1bJK35J/2HciJQcpZiMLd9Sz9lLuekH//sxUW3qAWB1
feHlGdTtEgaB2BYrDy88ER3a5liaK7Ky4qItlZmpz65vLwFed1vcYRpeU5NndKJj
ND9pzQKCQe+60ADUyDdWTIL4n2B3H0uWiCqcUlL1wqz9DGrv0i0jwhcV+eS7Mhmq
57ol6uGylTAPvtFP+N0J5MDA7rzpbBpPQAjM3PyQ8xLjb/Zpq/MaYVE1boGmBNDO
VIrafAeOWnCl7+6fcUCHI7ysXXPdfyUfLkrYrioHgb01hFDIRSuL5KiA6I8XUEq/
i25tu1Uxr2DOpCzAHmyX1QbnsEcjZevOSuzz5Rxy3F7vSHYz/nGvLdqEYps0WujX
q/P9qRmxPNIIpAEtB9+Ipz/e9oLLXZMehLUxvk/txykc1ruhK1N+BTyolKeJxY4J
IjY1KtuBpBONPFZxEO6bRhJUtI6r5Ii3cqDH6eh49R6TAP3ikGYHfBGbGDqUT3hU
6yM5yi8PDvFQ/OsKyvgolwd8rqP8hTQwdtJAFLOHTGWAAHsGaMBmn/om1B6G9FMc
+3rCEGBzrdxZ0hMREx0VeRHDSxRHI0ANvnLvQqLJ8AICgpOcXmvoUDYhMvG0ugf6
op6skf3SBmYnutoS6Wgb238OcLXScwNh9iaElQUDg6iiPxFXsBSCEG3p66xheKCd
tS0l3gByp7NOR+BxCa0lXF2I1kXXOoaxpkEqO7bqzPni3A1YDrk2AIN//iqu5HjF
SSEODUiZmc7qgjH70GrilV3Pp8vOMEyEra/XkljZMMDoheq7VQG02b2nJnN0yhD3
1Q8vxMWbgz8y4yZPBpEOVHovfQ/QuJ9Mp1anKRAmUij1KC+NroJKUgJlhysomXRQ
ewxIoQIp5hO0hr9dul2d0i45t2k1iY/50m0HRmrZngxf93RV9Nr6nUwKjoYTo0Lf
3tx+eLMjgJ3hz6Q6ZqrkR6F4znOEPU7VOeU+0/Z3iG4DnwCza9DP9WFyTn6zTNuH
5HKK38VUVf+HdB/glgZMksePMgrittUdfRV6m4vzwv7V5XabGVdgV79BIRrGZWGq
wsEo6qBW0L5zPmJeMu4NuPwCpzmgryJGGZdJILG8S1BC9xmqIHoACDHUZ45d+FCR
ofCVADmZlxVMtEcz/en8rknjog2HX016aufjxvnp4u/TaE1Pw+I++SryQD15v9cY
xMFS4ZNz3GuIVj+Nr/nL6g6tUKF3l47zdG4etpeGxbHmdTII02uDkjtr9wY+7JEN
67QE4ZcLzUjh2Jtym4ztbHKQkdoSbFhrQ5oeLZc1EIWjhX+Oza8yFhMi9K91+hTP
BWLkRgV3+t8dbX3YOeyISR1IIBobKvZxZWsF/0XDJKijuqlqjkoBztl9D4zhJUIB
L1QU0RfLsMHl5cK5RSLv7qjOassPLbTLGiMHAF/1Z4a4JgKl0JLYONMTIdv9qUfe
ihfsWqKUIHEWAYgqk/vHcJRgQeXw/9DbyIgIMvkMxCvrdJkuHhPdFSfciplvaybz
67NIAHQaLUews88/iYkSTFcayAZcKL7zgORNbdR22G+njz/7E/w4eWQkX0sxytJ4
3CPgfgicFfVVPaoj6aH/4Ayt3LDLZBi9+BUzaPjvjYK+nzJWE+4hgi3jiuEEwmQ/
Z5b0wB8InysCGiP0nSqt40JFNnIzbvmsoWkQUJpayzez02mf0xnAe+m0WCqN3sAT
dvDG5TrYl7P/t3ug4LZiBwdF2pxfgWwWox+VcKiqIUy1lHi7GrYUZCGPxvnB300C
DJxCxgcXCaniYCx32OTEBoupyaizVSe0Ac89an2xMcPi2pfoqEPFLT7ohv42JF5K
JeAoobXY/g1CeeuYWq2/uj8/1IS6drRAVfEK3D0Bkadm9T00fjIqtbMo49XRFyVc
UKWA7x6fDIWDkBddwIx8aWQ8dPh5qa4PnS8iT5jdDceR9aJ+PwUIGc2q7WSy2mO2
MWdwPnUHFdknb/4QovWeHWt/LuUGEuk0zjQ0bYUoJEvcP2g3sFDiIf5Y0sVPJsog
PzXiyj2K1UohNoUAxKWz7id2nN6UWVQ2QjL4tzUk74GMhHVJDq/L0EuVDtmmSB9k
lfaoWxvA6sDplK4DMRQVMtoY4I08KgTKhAg6LUm6EiOoA/i0oZFf+UfRZ+DlRahW
t5Vr5EdtRqH6AzDN1tnqmjRVrjNdggs9mxw1t3GjynyNmqqc68x2dIbDC0suZSKU
/4NvsCF7paA3PWInvgzjI+Sed1dW1iU9F29w7D+3IKfAgTYBANJ9gWbci7yD5EaW
F6GA75Rqf9POTSNbR1MiHJ5T+VrxE90y1H1hoZQgdQjgZpi6mLQzAoy99J8KfPXy
46uBedW2+28GKCX+TvdL+yL3blRYd9xQCe7yjTFhb+qTGBM+2hH8XuBzDtIgw+wD
R1pn5nWBzxj1RQG2qd6qfJJDy4qGMshiyy+aKslGosV+TN69/km0Zm0I0qaD/pEV
4ZYz3M6rDllUtUyjnVQk1XyeRp/H4vKkKRjV+Xat1rvTzE8FVxre/jTe3YJsJwmx
ZD2nNKmq5UXci1Tk8/AiDdQb/CvMjYD7BksFzAtlOGZqY7b7M5LyzTvwYSA3niSr
TlIc4+80b1dALnXsnEUiWKLOQtWNnefDojlexsFrAwhlGvRbj97PtbEMq9MuZT9b
nBGf89Fq2ej/JQrEg72SX/UfeQv/JOzl4duCnPGhtrjQXsiqsEEVRbyoEGqUrAbK
v0ggS7VklhXh3HvFO/NZjihcYG4OYkzNI/G9kJiWVSgYMpqYAE8jT46VPrxCwDzE
FdBuoc3Us0sxODt1itEMdFzqq5z64VgJ0eNF4mIwf4Ekgq51uZPvzXqXwHbdBHzx
bsYHv9m/Sk5quurlMQLmU8IML5amloPMybWwvorRt9EgbBJ1lxTYSbnFcJPAufBN
is9GyYOsJFdZxU3i4OuUw2nolLB9fdF6Alx+jMoxguKuI5so/pJEZCJBzRlN4tcz
ubVQ7zYvQwRLIZmrN9e1Jao4je5zFGd0LPDn2umEuoBAHJijWGMCXteyZgsLx/AO
mmZ8cXUS61d0cIlA4I61lV+Ba7CxQxqabzcQtKuZCwm3h/omoLpE1IqHxjjGcE2K
EgpWXg2YVflUM/y9IrlhTUz5F8abkDcZqKM0bgm1AyK7pfrq4CiIKL5CBh0wbfML
49CdzVCkHjDSPHNqwdYAsjYBSlahTNpseaFLq4oW01N8cvmkPBnShXYijUaSaQoM
2z/sXFN66K7fzhCTcUA7wu7NlHzoSvn+4my1nvQoopZzisk0FLq47BpkujZsR5ig
28w1LFmdbpcFzX0i9t9wqiaBBEg52Ri0fFhbe/lpi7xqAHZuZAIIfqfX/5+wVT5b
VG12Hl0r5GpHnCP7vwebXXDHLf73Q52BwOMSOH9DppuQ3CNgm+ROQld0R8ngGEMQ
gEPkHClqo6BoWRf4N6wMKRZUFxeqkedZ6GSAMScieVFB71GQspaoki8IVfJ4k8RL
ReWIejzvNkauMGts3NeR2h0EKNhYxhQWtftm8OmqrJOvW6QeImeM0Uutd5RWSzs6
aH+ARIW6bjU3qCIT7N/6i7wuGwe2cmDUvxkx+rCxUZp8R2U4kS2vYahsDAragWh9
nisqpBwYabPxH0ShIG0P5WDgFL01SPiBeEpKb8I50bk+iF9dtoWtkGiU2qbgbhW4
H5zkDuwzhSe9fdrqXPGnPn5urVV3fFgTeWazThwX9t8ww5nn53/hpeJV6nLjGIaK
9+CWZWG+97FEh6Z2vfw3KmMIDE6qDz5WqzYY8VNWCiZdSG7MMgKaVIAtjIfgwZQc
nlE18lvXxakHLgdFU243Zh9GKNdA7rSd0HN87hRaU6SJ7yAZAez5sazqhcSvDYf0
mgHUqeepDEW4pExMtnRivTbXZSTgLA0E68ZFf85LyR1qnS79EbysfFh6dDP4R8Tt
qA8ebfxEgKKP5jk/+dxZThn1y8x/XgnZcxWB99vdyeENj4x47R13eXt11uRteBnR
+VI0V+YxQEkgx9eks68ATgLhiW9nrF/jaGx3pUrX1FPndy6x9OIrP+TYs32y4r9f
FsSOLQv6IanPmBEkBhu2IifLIBgm031BQf9bYbS5JVT1910y9Y7UNNdYM+NygBTO
CBgjlYR1b/nGAMvjLk9G16JAIF8rmt6JQEZBSmq3L6feqIkaDdTPid1U88vOFr8v
Uxe1bUgWtmtTLdK+gDEqPZx8x/Sd4Y48pG9YpGsqauc3SinBH5zmqv3ku1Q7vTrE
AClowlHNq3uP2owtdy1ZBSGofPkAPM4fpWU5AcZQxGnDTN8VzHjtEmlOy773I9Qc
iAuqURewsOxz1DZyHdZ9rwtP6TZHO7YjdCHs+7rl35/rFE5CZRNAri7/LHMtrepx
5KgwPeVqArBZ1wlVvdYMJeaJ3YfroLQ2kAGiGa1O6Jxzd1J/7vymqu/ZyV6Rxw0+
6mKT5UEk1zbZiCaAi04KnEFu0U3ScV1qZ+qjbwgq9FVdepGeG5J0cZ6G0aABrNPS
x6cBz44/EMBKTNn07FxoUrZhzs57/x5cfpwrlXpU4B6lbCQmmG60oAh1AopNZzvb
cQG/6gISSAePBegXIxGgK7MfXSn2wCHHGfOJzYVghau55pzhUshgzi80vu0fy2K8
94rhAJTKMSPgjrhDhJhY6GmY4LfOujkN6y7yYgRJUrXbWMr9VzjAVnPdx4hbI3Vj
F6aqR5vDBQjf9npWA2YNa3eiskcA9wiY4aKGucnPzxbbkPv1daSVIzpSALQYfwkj
IRLuAIo3IoX8rKIUubwfp6+pR+5cl8z56tISYf6i7LLCM5MxjlzHmXQZ5UvZ49D7
FVcqacktO8fuDr8ufYDbDxsn7FV/N8AliMO9neIwszDGMtIqlrYeSFkJt1t4nZNx
leYghphXQ8F+VCZm2zD3jFqseRCvNOZRJBp4aKXk9x9HqAWZxL/7wBpfM0/mu0yT
PgVBRAZaOJBuk1iD5Q/YslndVvVcoitgxZzvdC8UOeo5+fZHZMrz3d9K74blO9Lg
bAYawjnKcOog/SLiqkQRAgTqccpFmu1DAqMhSImbcJAgJbGe/AIrtRPZ+XJaDNW+
n2S2sWfxLlsTYB9VXBJyC+BZuE3ACUHP+x7d9Yiwf3kBOBIf+srJ18ChnP0JaT2q
9VCXm82D6g+hgSbPSdJcPuHYF0N8KU3GN5H3Mdb2Q7U9iVFQ3aRcrps5czVLpii0
zKXaQung7/1z/iZT8E3y/LPvGdi0jTkwDWQ+uxc/UJfAgCrkDUZkY0IQ/if5vkwc
2YLSiqGk8zhULrn9MknYd79KcJyHibFf8FZQNCRl/YxsimP8dq5gro0V1Sj27FHn
NFcaWmFh/Rvws7lVnA4q9EXQ6+Q02OVJysaUSi2xcSrW9rHQWbqsh7hVr5QZ5HsI
nUCTR9wVyV+QrHyUBQId5tBLNX5k31mQdSrEvRG8DS8BC0OXIk1i1cclBIhRkPYo
Y616QQGXIgRSmgFTJNZsmkDK2sZhKpJLUcqaxi/nWhrpP/e4IKM3pL0+tIVpY5wA
+kPf/pzpryBBs9DWi10BIfDvwTITql5ClWooRth+sdSCQcjRp8wd/45zJggfkuae
4QJRwNq6eV9e7e4q8tg9LUKzBr/DQkI6t+5dS3S+46YLeoxADhJNmS92p+9DKTeQ
y+xZKtZJs4uEC4cB3xggvmSGgRrw08tf762prDa4h9KQ+ZEp1NcyVLvpKo0bNzVY
20uLHdc5LsVmg/R56wnWftvVw/N2DTOd9PwvJSUH4nhvO6gkVIeONTJGfhmFqPcM
BAtNCYJXHpEvYf4gtyHxE2pIxm53p0HC+T46russgHaZ0IRGV2GzIqJ/37Va+iro
MsIqVXHbipbJ4zp1+I+R+P0/WjXs90dM3CdZ6+BUwNsH2FCdtMVUssXibEA440Wf
FIxLzqSeWrZYK03Pj7qvAYdQQG6BzX/3m223ppfAT8ChDHFXJFtdfleKw4sBc5YD
35nZm+L+IX903jmhMZY9Ab5N4m4G3v2rOgTFI782FMdDoSN2jpR53imaK0guKBvD
rRzWsDi+q1CbA47G9P0IFueFzxuOih+J35CyOHa+LGwTFIcwvY8LZAsaj5WM9NN9
6GX9NRXlG8rzX3LMwVJRRvXtOz65mzetYUhGhYRkYxwZWs9kYqW/Ez1JWi2SHbEe
+5pWQvH19TUxjJTVF5Am85VDJeqd7wPyTyq+LDGWGCZ82NDiEh4VibYqbkqVz5LO
D5AJNGdV3ivjsGPwXKeNSYSQRzkw/mpS+YYX66afCrqZkZSMXXop8t8nCppMAuqk
IKPeIUY0NzaaJKxB1mSY9z/hcLe3cpNXsISAKPBOW2kvU7hs+m2jv8KdSBuj2bmo
oZRUM/2Pwl6r8fNU3i7284XDj5L3uFrOUN90Vo3Esr4EY4Q7kMUefY+Gx2NC8g5G
lNU3SCIpJ3DcmbJU6uOD3AtM5F1MigpElomyOhgHCes30zEowId12FNs5BTgo7Z4
hDyBFooHhxaRX08UBOXuYck62Bfx6dq5XU71qFet5mQb84aAckfgLz+N69TGNcym
vSkXp8u6o/vI0eo+jvcxOcozCGvdWlf4uXMNdyHkaZhwQ4m4h6iujmlIrhOt4+kX
1S63qzCw/cMaMNTdhkH3oJUcQKHBEu1QpkjACmJKA2e10pIJQVaQ0fnt+W5sI0IV
nmO75w+KX1em3BkRizsBFCeWakskJ7EBnsfe8Km4SO18X1/3W/UoUoEThJFd2MzT
lHyd438jq5LehQAkA2L1xg+ZHB2nRe+MkQFHwFtwVoZlmh2VTl7asdejFWVsU6ZG
uCjLD9jKj3jmB04rfLMqjntMSgMv3dLTEcB2n8qqzEWVEp8TCzSZ9FEFVjvVl0Lh
9QAcaZ0uzCBFL25dpa7ipfqWoCWRU78iw++52Cug1L1wq5oG5y+mvZJVwUnzr/ya
9NRV9ZE1odc8IvwFDnjoGANfdQkE7pVVvcWKCwyBMu/56PhCiO1/U+XYRoegBU2x
waeLMzuHPbinpiNWnuCgqb8G7T7VNFbsT5dsqCoUFdpwyX0E7528SZsLHJNxcVxc
Qbs3r0a47P1PF4u2XV9U0l2g73fpSAk3++6zhuLpkPetsGD8RKbWkIXxQ3r2Abqw
LqvUEj5Nrf45zAMyiEeApCcxhBrtR2JQ0KvoaRKAJj2KoJvAV8Z3UQUW8avvC9+I
X2vxxPRSSLgkj+6iSzioCeXIZAaGfm5KUi8pLkbywy7PXQKdYVtXh54GEsT36itj
WKIk6wxqI7DLFrf+ks4oSb6Dq6q0aRZuzZZR6fLtWKIfMM6EP+3BQ1JReNMl1Brw
Yd/Vrhc3HyPVR526KyMc/Z3YOtHKtlDqA0Ru4yCCEAmR71ofwGCnwHp4N0vVb1hT
x87XvfeA4HPY7Dv6z8XWy9Fdx4C8iFEbuPnYPeXPj4YWcEDPob3RASNRMg2JlzJL
04+FsznEE4Jt8ewcGM4b73MkTew0GGzvqp7zKhkBc4PDUPdQS64BWS6sJEx6CGmA
VRyC+8eTEdj4yFsPAHFgBAyCmiX7QS+hTkNPlRV78JGsKy1v3ZNFFiHeDmXB2b/n
fxs5b0yqxl5wFh3gigeMOLsip8s9qQkxmG8jXfTbCqKJcqifmpJfmrJk3wm2re67
Uidf34qn9cM3OmNbebQBbrUMxVGo9WkIoy4VMJFt5YByN6karRzoX0kWZHNoN/4U
KjogzVtvYoDrEM3HR+IQVYo8gNIigBH7ZksiF+VdPnm53OSTOcRQBOaGtAVUA2os
Xbc0+vRP+Zn8y7M8L/FXYvW1bfuBXVvM7Kp9QMA0I7pEXyTh08VyEhQOnBWyFkSl
fmImYDTF9ppiDpQ7o3loU0DGNc6TYjyOphGetaOrACyDI2PfNAHjKLNiIYdpbFcU
VNIi0eN5LA1nU7Vu7GOmv95vudD4VQ6Tu93LESpSJwZ8FhLYo9VR120sa7kDMOF5
yfyXDBZmUYCrMnqG8rtwgJ2orF1RKQLGO94toDpvEMGOHjoLJtBLgflMEuwtmL3k
OFEiW/74aZGvHGvMnK6cf4CHxP0BKyKA8q9tRlPXzHjZhq/TvKlU5ke1V+BTATra
GItwpLJQknmkiagR04kJj/uloEJ6vq6AzSfDFX6QRB3U1YGbr2HqsjWH1V4rGt1M
eCqZcXLrD6xrd6OiH4veGSkFkSCa4ZeIH9AzIKWCWPAizaOSHUC7RV/arNmKHiDz
eB9axA9rGN1X8OIY3YaJfp1mTTO17yyb03WNa1Xoz0JG30chbG0QmlZ7xxJYR0Np
/4BPuYLzmqWETLT/jTvRB96bHLzyQBMpE0cmbR2BRYLSDQb5gFuIIvO8DZliiYEr
hwEFqDrAtQN/OFRHgTJ2ltUIFdgUSLiLG742DopTWmRU+5GpPrYd52xl8F6zou/y
rwLn51La3lPNshMAvbbshiQuVcXS3GSycbblHFR0KPgtmM9ue47h+FgAWXoOGg9A
GT3W2Kvw2+f5vBEAFIqPulEolYjbH1XpBtwblYmpaFHE/iFKjsaKNwbZPfsqTLb9
OwJwUnpyX3jqewpiImWoZKjaCRp4KaAbV2kV3EkovkdTXQhUSsMqxJGl/AyOQ8LE
3ITicQbr24wIbRFcF1/39XnMkaoj3hG7RCv1byQtglqrs7TSI3NboO85S8O0aF4o
OGnk7Hr56Q1l1OwK1UTXLzUSyVjtfTspFeCUpbU0vQV3ZkiA49ZW/DITig+QN8og
/jWHfNRUK9TOz+GGHBonyRM4TClDh2ZLW56VqFEZ2QWTBWMTyJeatX15qHMhBDnb
l3/YyiuhW8uAy5CXIESeKr81X5bGCGTOBo8gi80YmyBl3z/3dMB1jbZwYH+HCqyL
/F08J/Y4VEczJcM5m1dbY0ZUVBJTDFbyVMjJsbE6Wj7Oz7WA7/P8421gkPcm8RTf
5SCUCScc2xITkUGVrzTQWT+WVyls7FQNMIAQc7tcmyDKJM09GNGykys1qN654B5q
cLlKQyeetpeixqaHy9WkP0gUjSN0phoZMvxHNdEJ5tAi7VdaSiUsoWYFbPyj+/H0
L54+ROA0Pq2woZCcxL3RWs0g7OC7zhulZj1RdOue24nAj4uFaK4D9rJbX0TdqLh+
LB7h9iPgztK6At/LZ+yLmU7ZETb1Bt0whIRXGVHbRMSVcqXEoyEif9kH6hLugHTT
CfGgu03YImylFiD4hXbikxKfwtMRsfO3lMFaOWMYVqgRP5jpz+Uz3YIZj+Wm7Wb8
HKfKn6wgy4u7JBbyRTnTeBiyP9+an5HxtQTQ0lLY4gfWhiXzqyHClbPwfYFz6rMU
6z62sz12bc+GCSv5tHeS3RHLhBT/LoVFOGANPLjKFOV8iJ9RoUilxbx3HdQAQtiM
Kr3fhQcO0/t02YxiRdMcJ0pSJb/57F90wxxRbpJb+ujqR4ZrjwH0eMVwdgfMZ29C
XiwbFt3wq4pCT5BKM1aAzo6I6z3nzpvhHWJ/4Cr/P70YsWsSDUVCkGT+FUHjHUtB
x6eYWK+e8W9X1PSMNatZulLBCnRkiYQDHs9RnvZQBPCR5q637mCAhY7SkEGHXVi8
LOB+EB48JzBNsjq8SzGrS43y9R0jnyooo/qyOSGDPqLqtsJUkCKEskyZk7rbGu98
t4VbcS50Uyuk+BrmnO3uW8bJAq97E5KPz7eUDFc/0eRj1GSDHVS1JW8aKcP6IIdy
M+6c9x8cMJnsr3gxKWs9jXPGVyT+sNhVEDDQlkVORUEEXYLzzXcZKViOLqXZzkxg
cnNaPROPIxpnmzpwHE2Z1H1D6mbsaANiBd6hZtIT/6DFFs4KYdhjC7thlshCNAeM
0N83MaekbW5wOdcV8NQVmSNOIdK/DSir6w95n9TfgWJm05rCin+LR8WGuyeDqiLp
EViIkNETHTp/Yo0Fn7rhdouY8fMMN1wXpb0yh8226z2jKz/CRIWQudrUI/9Y9JzY
nqkePFqeM0Z5cdlA8OJxgkWmMi0PZvr2rTsvhp0vXyASNJLM4tanhrwptc3K+2r7
sy0RqdOVE22hWaTvFj8QKCMaI+3h0eZZ4c/LXWmVLCXGsWAC4Ht6J1A8JGkhVK9M
yhvXgvvlA+3XNsUnljlzYCRVYOepxfXdJjUqDpIN3ITivmk7PyY5jqHbYFrjgicg
Hp2fOWFV1oTdPgZP+kxBCklnI2amIK0Cz1YnWmjJ0guDl2AM7rbwRYuziwKcMEQu
D5IExronuJ05uIlXm2sFfXTQnxCdAqgSsrKUYCrEvM3W8AdltL5aTIx5XT9L3CFV
mBwaF3tApHp/MnQAs8Hku3q57LJBjzozFyw6avA59MnNWrYySgDPR75yrcohZd3B
luHSEBVmqK4k5HdLiMQBppvpTRKcjXuWKenimWKwJ6leDCVB4TAuTuruDXiobr54
m5N6gtCDpw9iJu6SG4Arig+7ksDWEwksMgaYF/0M5+C5WlmU5ld3G2IANFT0pnQO
m5y+mw3WCBRow60VIuuFhzYQc8AoCqrUj9Sh3XzrfnnRRpLFRsWYTDNK0qQVfe2M
WsQe9PN0We0Ti3ueoeCkhw8ZmXBmbuDrkWWpCda+zDJzzSBbHyAR08N4i0CJL/df
Ku1SRIVIxa8b08LczDNgNImiQ1EG24grUnoazq6uvx4UlLYhqpU/MqQMcVGlwobN
sSY4LUQiEwPDmxiLBADsH37RSqLZBwsjbRmXDYlaP/AQkTKaSXIDH0fA6bDT7aWY
6vwmoEVBx00bjBrW6TweoZHbkiN45YizCKVNhIuxOPNK0HRxabM+lmanU0ZfiXB8
44hVNITqGaICJuylZJY6BBT+uAf92ITeeJo7YeRNQNtG+KMBCQ/4pVtsKVjxjr10
40tA7fJj6sQsQ4btPPGROP296+Rdp4n+Nend0v2iQ+PGmURy//TnDwx2ibnHjQ+I
fxcoQHBfW6i/OEFDDXNIYW9ahhnviRTA5t/+zMWkJXUoC1MML/NsOywzdHmQ5EMG
JQQH5GIE0b0vkzLQ8XZXQcOvgcf9atPFGABNgDExyeA4CuioYFCBvE5nH6Lx84O+
+FqhY7Y7VRy5cfqC5LWCreZ9JxQ+J449F5SnzEM5DK3XQLBdrFZfeZNkvP0octq6
T3MWzQL3z2oQK2YxUu82sunHUMT8KBIywqhNDMpc9+r9tPbU/adMjf7V/iZU8Hmc
/RNx1m/H+nG/c3i2TyYapd1T8w9yDNnTy4wgWuflVh1mBDOR715Yg2QLuRRSHhsd
zpj2pf6x5jhGJGOFwqBbHtyWF3rEkBRwc8n9IBMOgUCdLCpkXX+BEQHLogR4V/jM
jX5FgXufleUPOZKLiTyXVrCL9DViFGXM+07Ay6J2/qR+uf+FwmnZCOiajeWPwPTa
ineRL/lUemr2sJayOnZ4i00CLdGKid7mFLQad+im7709gY1juByIrnPCF8TJIf5k
1zDV6a0gM1ce4Or9MxFVX9cuowmqwEZG/go06YnbrIwREy8Y8Z0RC9OuQei+fNb+
Oz+oexP6p7GONVa8zwHgltT1pdDC2AVx2+k41YH+N3S4TaekR7jWZG4lBlihP5J1
cc8BniJePMy/qeqKDRaemFC3EYFjXNxg68e06Q9UQCZP5AI5BeCCBTfGiLz+1YxR
v+dNpWL+pFOH8QKQkGsBJjM35op2025GZ49986tsEjBB2OI5TC8S1nGFVDQRzdZ+
DJ3uDluLU3Eq4neSsqKUIfjwsRfmaIlxs06Yz+2AF5QSACqy6ZnUkcO1ORi4fHTv
o5OvcXNbKDtw2zvkvX2AdTU+EvZYJ0oh8mrKJXx+OBE/dDdrhafre6UjKAg/eexO
xsQxTy06ycSFqNPNv2/djB6pXexFVuejgRTWkW8G9twurvay7uPUmuqMMnyOQRtS
cDIreLq+cgbYMujrE5HL5e0NoBQoJVlauX+9h33DrJTt60bsSIYSRaDBH6gngTvh
1WCVomyJV3YB6iUaXYZod6QNs0JvmGcJdNdBmwFsIAGcLtLR/XKk04sYOEdqdKbR
Fv7Na/4uRODaUlb4zRU2MUBRCWQc35IlhjNMCjZxCCtDDkCqF1akvrcmzgjG0zSx
TLPvgPVtO/AZ6C1sk1qD3AQqUkpShoXD2dOAFfe8xeIHR1vOezMMKpUj++1upEa3
qfmFTfimHcqtQDqXNnbwhYGEWh/XqjAJMx3aM7wpwDhYVnGgAZiTOWZdtSntT6Tf
nvsVzGDvhL6ablfVqZJ3AF2XIgTArmT1XAhYdAtw4NMrH9Mi0fmZxKAd8R35V6dN
Z+QXhcrRvny6iOqMsthxrzL4XcyAj60mhxR4fuHHLLPO3k0ggE5QmETeoFb+pEMn
p7HBMDL14fbVvDWtp9w2x7CfINjHOfPiBSvnkwabLM/pxWJE4uGS0uJnbeeyvOZz
XAVJza6PukRL6nhBeZ8K/TqNWkTIEemgoLNsIG9IUdLc9W6dvmJ0UDOSHQNkn4pv
PdNFWS4qGscA7n0ihrg2zTGaTSHMZLwuruTODSSuu4WccPQQ2FjFu+8zUBMf7+FS
+LEjAlIyH+dTPpvp3+Ojj1GnEi3ATS+UEX5q5qw/3z99Ee6Ae9FnQPl/fb5tU2D/
mvYl6DBaMJZ2Bh8JTB6T6s4LzfgAxbvK1z/PtbOVkmJEXpijw3+pM3QBKBMUz/xO
ccjW+Ln710jMbAchYWYvZhGx3FR8ci0Ul9J0jxrEC9iJKL+5OKDIcCc+g+VtB4II
7EPWXpPbiCg2GPGLkX4M6VLqsgOwikLVJ6wOQ0s0RtLwy+tzPLL2wQk4jexBc67J
gWdsZ3Eu53y18NJW4qbqun8WFpFxg0saKmDNwUaOdytDBFp/pueZcu3V3Do/xZLX
tZvkzuEFlrlYhcU2TJPszFbm36NLRKpWZ+NFrN1cSKdm5Ti7rCoLLt7OuboeA/TM
I9/3PLPzB9O3I+rtRCQlMCHJKC2lLtJFbZJLrtim6+A42vip0Oku9PoOniwd/Vf3
UN0FLC5TEmXPKnP5d/q8esb7nlkG48z70rTAbdIT+H8e3DdqDjh7G0zcypKYrn9A
uebDANMUFWqlfBtCJ2AngfkMNcRTpy9ziuBKb85pWwBLNa1IfFuhlMBgh/urcCFg
Y7gmqD0Gj/Mv9Fb27r1vI8C69IdCflGuETVTU/9x2Alnqdl41NFcC01CUkLyeRHC
bndBrAv16xD5mKtm9Bapvnxs3+yw3PSjUWS89mhNYZfNT/siLvGAFYJYBl+EYsuT
idBb8PvHuRJ6ZdP1rf1FFOVDlfW/DVOtqSH+Xrw+jyIvUTPuQQFNQbxVjjSg2VRB
bJ31JuPI/qlm5RvyDTfIHrXvxn4tVdBynH8Co7uLRkn6XOSGyYG0MLSb4LhylwCt
83fGN6DMn42eyrzuRL4Jr189ORrFgiecXTwHfe8+Djfa8jIiBHJJ3lvNGwq/3/e3
baeCHqX/Qqy17byyvd+veQIdYm+FNzNcZL9wDEvQZjRethOT/MNngqPPEtjG17+P
t8aqt5cYxh0UYgVX06FGsgOM4NURvQcKU5xS+kolSAcLtFwfU1B8GeYz2+5rPY2Y
AkzN2yM4CKF0S07G3o3DWKVRTLz5tPYC5+FHFX4IydlQ0d/6KYcqYt/7gvmaZcHB
rvPg6DHwB4gbNnEV+2YlHhm8ovMv1lmvlf/fs0gbIoWH1yOwoZy91Ib76G/Lu9A+
cNLcL7S/oDOl/HfsonGbyWDEe20H29LQsG7qij1w4IphkBWxtiu2v4h/v8j/GtE2
RxKE8JN5h6HXVx8TX3/g0fhs/JbpCybXKB9P16D842CUO+GCUfa/bo69ResmtPET
7SIZfHJZhdkYx5E/r6EhbdPwKthljNTeMmK64S37+Y+s3e8pKEp9nCLLDcC6v8Vb
Cog1vysABcgTJBOv3vpp6aN3f4swj8CDVC4d8ZPyRm3NI7nZ920dgVPvAymOdS8M
EyQ9aRjniA0SepXUlsk/HwQghwubK8ExmWSxUe0IN031ty62IDYYje368zZbjWOi
IPjCOvpMaXssDtcXM/T9ZOjhfaxRWZjQa0eakJfilZRT15rBtkznMg+JUYrAyBR/
Wf/e5lEwFef//tylFRnK4P9sty+vq82Xp7AKSsKvHg3Q9mCDUkWrBcApMb7vNUr/
H/5wzkp3eb5pCIOyqXVQattH5Xx1oXB2hjGNGUyRRlt0XFL2GBO+yMKCGFJvcKxv
ATgfY3rtTdogjqeag9tLXV/9vEPvwqv/CAx+z9+fz8b6Tgf7LUT1jWf1HFEM4sxr
RqVgqXHBT3HEEVWdUWMM154EFqJuExhrAGGbxMo6AwF51nWou95LNOx+atz0yVpW
xYIuevojmFttLy7S2hDjXNFlPHJ6hGKDU+hD9DSxD4Gi0JWLYHRRK7W+EE8TT+nk
uphvc5jC9lCWRHj7EHQI3cCLHFEmjs1IR6IAa+pGjYSTGhvMzT5Ii7AQX9cBosuN
oMjLaPE7Kzeoj/ewyEIYd+VRToszpdXZMKci73GgyfMBHPz/qgxl3XJoRBy94TgN
pyseAU4KULQRqrNmjicinuE2uQAaEWnYdj16yvmy6K8/FC+c1biS0zxnnb5Z3G5U
voNOoV0cmYSsFLB35ddttNOrwW/6Iu/7Cj/r1g1UcY7Gky2Uw4ZqANd9QhkTQK8s
8FHGG/ceoWXXIEzPyTm0QY/TysmICs+F+/SzDR37aKCKlAkRAphGpL79kd22wB5u
3gzsc37iHAAyVCQMYKCR4EAP99lZridYgJ6YtKpmFPeMV2X65ZSTndA0ZjRVP8h9
3wnBf/qIPKmrtsiU7wDqz9spAfKE0fk6du1vW5c91DFkzPym9Lz1t+KT6SoNWxjP
gZZaZx6EL+XY2IrFCrG7S7QKy9eWe1YuS4OUUACdef0pmYJnVjgMsQMkOD5ICsyH
d1tmmC3/fNFZdVQukA+HnVm/V2SpLdvvyGxEx3aF9mOxmC7DbYxR/wha133OOdhk
+Z/fIKdP5H4rvQHbq4U6rsJpYwT5VQjw2W7uZsTpPOvoWOR/FAJmnNiItKvLWn9n
9cQDPj/Yzs3Sn4ys1jmEprd7ulkBTDNcd4KouT6d3CYMDkjSXz7NcIhHOkWKEmAs
LAamRsO5vVXKz0eQXKgwLAmPId906grr0RqBlT1SgcLalY/U0LcLslZl/jSb4ARr
aPJPxyYyq4FyEyd9KUVwzzMO9lkE+Y4KUwzj5O1DlTJ3PrdqFe8yp77pZcFW9sei
JNpag+DQFfPU3MmqqYfegSVGkTK1q3LJH/JgERmukrQmOlxq5fziAgKzlYxig3/L
fwmj94BO8Q9gnUIKxKGB49RCtXQ2Tf70mpRKe20At8Wzq2qCtzK9wLfQgNFXlTpn
wufVz3ofx/XpMuW86v1omUngwSjOS9/w3sicdygHvc0jg1WT8VnxPC7Mvh8MfRw5
5tVoEFLOfgMNntHLMmWwSCps3hztaWcDeawqAxCh/jqIekhdKV3I9vs2GPzKFapg
/EH57EI3J2cInBps/kXnTO+u/Z5CRmss9MSdRcm+5LXKlpr9pHiy/J+512/MFAqT
jY1BIs2BoAcPVim3o0K6GawJRR7Wnq/ruYn3vL2B6EYs6whN/4mlSkJ1VRQmwQsa
4XxNiamUGPQfuhHuSfp/XQHlJVT/x4/EaLJtoR8tMiPTKiJ2s8LbIRGJS93cCJfa
K11g1QEadQyd3JS75iIyG7H2FzwEA6MaFEDOtwJz6F8tNv9HG6cMJUwTZxp+eS43
D+oa5sLolixcBy2tm4k4Jt4gYqmHK0o9kJgKviTncT0nQLcIKifs3a/nKKWNB/pE
ev1WBMcqPPG4dClUSZre/ASVLsgukkQk41QQI9oKVGtXrfp5qXfdKPI55f/Ph/3u
4BvHxdZD7DGHCHzXVECt4PSn+quoNVXPOztVj9bbCs2FOZjF9bRRz8GsCD0lduDc
jImdC/2HpeS0SdPkGLf5LK3jLVDnGpoqklsLTjXrU8aBqPJcFHXHl0BW+chyq7++
mJ7/f90iiKZrCFmpU7/+wyo57vvBEpGKiuzi7qdGRIkRxdWsUYzBqqF0esYrFq9X
DMtFJmN2XH/ZBF/Vm9DWf2igIkPqPIrKv3v/wN+l/z9aq+tOKmIhwgTBnWnxku1e
FAWzuV1JLpwJ54se0a6KbSRNN4SWiHwqtYKWn0X5SYIwmVN3O9kQWByrW7zgkArD
5SMeq3EWVhl0stO/JketZz/dJ+Q5HyzX+wr0D1jGQc0qBEB9/U35lIpTcK0OIb5e
+pA/UxklrQa6aPLlzH7uVozvC1/ybBgLZoQQVRL6Y7UKWxBTpLXrUi/EsEouwvVq
peXuLVUoYn9DDqM1mzjqg6aspb5g14MNCGTdee7EBL9y4p7Ygh16rDwJYIJatvE3
L4LskxXNqsT7VYJRj+SK55FZawqr902Bv1QJsGN7SvL+oGbzP2ipUfFUesYFvaQ6
80SxiDsqJvBmWs2S4RRod0WzdXmG7KFIEtkv7la4cqY2bb/GXAIVWMl1kq1U1hhU
wyPfRaH+YAe+OJgs3/sL3CuawvtgZp03M2o7fvkRYpqLF5U95wu1YSHM0FQVKtxr
JtWm2070IoRwqsZ3DyQrTZEGFb5PDF5FxSOF07Lyz20M7cnOycAIguakuFNSHh8q
2A8Vpd1YpROWQff0UQr+SPyz3lzsUvz50tcA2F317My5rb2PnJOWH/Ff2XgfXOH/
vubjrGL/swQn0dfhVS/nflSQjgJ1rDP78P2IHFkEK3ZfXtfRB79XmMTtkbhqLXCg
bdlIKS5gdHYf3X2y7nXBjxCAUd7xSQh+lnAyIyC6Wvl4QcmExALWwbz8jarR4/Nk
8JF10rC+eLWbRtFyFq2aB1nVEM7KqQQgni40T5+HyscZqGKzteZBU5U0Lz+KXMvr
s+NeTRIJgB8BGkYSMe0qZQxLPQ5omMkvxj3YWeiMsrX0f4BHT+9l57xlsUSPoN0d
GnXUa6Pv859E0bec0PUu4dNTekaGyuPg7AjDpnXYMdvHTvZrk/FK4YQzYCdpX8Im
18mFB/nfSjWixzKyxXr7c1B84VXK99fmvIZYo86rq/IoRjs3RGrUlFmu6WYofdaP
p1Puy1ka6GQi0YQ3WzWu0vQRt4qv+4UARynSCJHCQt7NLRrkEmkrbhJKZ1+WhOeV
c77VQlEfL85boK3W4AaxDzjETp/Y46UxMxK5OWqZqz+b2hmI3I4RFcVHlxWBBVEu
0yITLnznr3c67AppGu98ecKFm2OF8/7Qsbf/+0GzG9CrKHrxm9DYf0Yyxe+lC4li
fqPS+3JK/mI7deRI7SSJYzEIvhc/mEtmPJW1y4E0iQPSYTDos0tLVan8+ikDx1i6
sG0X1Y9QC69q15X4jf1dLhMoq9sYQQ2gIQI73pXgkz40Ys0ciu5Nt0ZY4niq5itG
r6O+OR4kPliJCjTL9jJ7XPBCJMe1ED37NqJA4PbRcBhlaH3k2OJqf87rxnKEQLSX
e13b5w7bm/pscuqmWgCUhAr25UkcUiFRdUTNgaRbZ5rtrBXtqME1rBQECHyOacnu
c+WgCS/C6iTsODTei3f3WeO5/CoGVXq0u51Kgfz1v3aX7toCmjhs0okwXkfFHiVq
q3V97YsZwLjfd97d5fkc9c3hGYgA5uiNEYgbY5Q0GovFOjxHEtOkELCbmu7+JKMN
mEqaFMBS88ub2R6JaZ6ARUoIqGgZtsslyzzw27Xzv5VWPTtMpIgRtCzC/fdOwGJT
ErKrFHzBrgwIOX8CcpMn9fMqFt0p+cEogK2DTk6K2PvzvYUyE3IL+ZV+DjEqzmqO
hmQ+gyAAXFmnWOB/NrnOyZxTX+6FlBOUNIAWAL8vO2/VOp/wNwOnzkG6qRquVMIG
9QPsWh80zzjiKdnAvM5OwgZuhT3XgNv7xLtUKEGCCwcIBXVCtK5SNnW7VjssdCnp
nNCVHaBXOFzWf58KP0YfANm3vpZYZf0KQ5iDgMtmBHRgYxkd+6ZWdUK6fIneWRnd
HnG9YSyq+hr6h3XgRdfnbYwpHxNkCoBEm2zcbnySRv7ibJZSOLV9PZVAznq648+P
S7lW+ZlqOKYqTiTpTnx5nio3ggjI2TENLDDANNlFLFQzrtuF1HVdT8vkyTImuqm0
fE5dAjpkaXJ3p4f5C0uW/BZl/+zsdGDw8I6BDYi6/vuVRtjI9kZxj4Vz/haOVvjO
hO+PZJ6X5HL493Au6rusjc+mPuhWOglHQu9VO7g/ZWOwZ0/++U6RNr0YAlmQ1urW
nKbvOhKf46eRHGxopBBZdg/wvGIUQXQ4wg2Kt5DF4CRAkfwHsDofPpINsADVNJCz
n+mspeiHyieNS0FYYTY3oOBl5HoFOJabT24nKS+5QPJDvlFx/O+6sISXqGvvhOzw
85p44QA7AdkzIR6RdwLaHwmAFOzsNssofGOUeZifbvFVlW6A/Axs9MXudIP65XIc
RVdkJgPHL/nw1Y3DZi2egSki7bWUX7Re+Mq5KkWP7DKntSoF6zAwIidBNVfo9ERs
7gcdG02ickxqwZszNq1R93HnYiyTHA66OUffTN7EegLiAVIV7bWPTYZpdvQHsnsW
IO0i87psem3sUtki5i6AqC6v3YlC6cKXYolyUNdyV6FTBJ3Gcmzg5R0Lds1xvfBo
f433lLQojAl8kkCpvtJyfS11VwtarElMfjBx+7oLRCNYKtx/+m57SmSy+uZgDKnR
f4NmCJg4LNP38Svm9mdbF6iO8q03bMWtVz+Tvkt3WbyqJzCDlpuyp5tGtmKk2vS2
8JGZp0OaueO/q/MmXyX1/hDPG0ucZokyMQRpn4Tbipzo5QyUompOLH5On6s+6NKo
nHK4/AM2g1SxPA7i5dqGVOF6/yN2Na4kpqsxKu+CnEXjSu5+ilZ61PdZvLWMFMp/
WuYk2dLO8cqSBnX4Spx3nwCuDjsbBzFflEpw3icl60bG1Qlytf2wVMaWoFmI342q
ypvarviDCdGpWZHuN1xTKQ8ZVQ6KaiLbTpLoT6aX+M5BRAPC3sOG0GlZEKRBTKKK
nWA7UuYG958Si09PniXoh1JqZEVO5ONOye6GAmB4ZumAUXBVWK9xM7bGDwfeY15Z
Ta49TMIS8Dm0aEU6/4t3/eub1jycasKCCQX2vyHfKjoN4hZac/aOhal8kT/XFE1F
cnn0hNe7DFIXskURtZXtN1ceHA+rkSLfkJBVwAQ+Holj9zM6c9RlWobX6+/TacoI
aWt191fCSmX8z9F9Kp6MsnPMsHaIoIGqBE24k3WQUAfFw98O691H3bCr4i/kRF3s
24niyQmOhhB6NyOo5CguvFIfTeTVYsoN9qfGQ7mO+KGWnwWFegxw6VMOHJzOFcy6
IpsDulVmNEZTuDg8RpZzQst78p+I4Sr6cUqN0U+X1WdDTuq/gOxbn6bwFu6p2paZ
QxN6gQyfGc5fplg1RTcOIINaGjMTQcGGLagBaZbsvgYT31jgKHRHBnzIIs+j2qSl
X5njByGSKU8/TEkALI3T8Qnuf+N00nSs86JUi2D0qwykuahNflj+ZcxlN60Uh9PH
uyDlKxN6sks7i0kp6TDliy4GUMm/m4cxb/MamX00zC8Ci7k31Qs28qNw/YgxK6hF
ROJ/VGWfto8DH/WdeA9Enin/PwAh7XjwQfHFgbk1xyObalurfVYn6n3+1CZ9E/XE
qn2X89naXnWODl+d2BI7C0ejp/tPbL2T3hkA8npKXRpg8zVHXk1mphurzDF+pMJ/
vXuanlHH1ta0GepMLjzBjcYN1bVhF3utjlIgqbDx44eNFRuv9HTu7KJpKGcReC11
1lzuRVZ8QcsQUAiqxWGg3SrO6Wf3f6/pwRUQ5gg6OytlWfjbeGH2cJ/Hf5N+MCAQ
gMM43A6ui8SR28CXMudhoEEVK45n7MvkDICd7TyrKb1G/u7rKbTUmJYjUU7LbQmN
7n8mrwbsvTM+cf+EDyikxfvhTdStvauKjU3lT2XJfNvghFmMOVXyOuRkvPNWyVEK
m9xcYDPkNeVqalEqSDsVpH155AE0+Kddmd2/gGjZSc81gDzT7HqTY7DAVhZN+oTv
emoWHzH3q0sEg5hmjQ4Z4OHoV/HHgwzLprKM1oMujG52Pr2d3aAVGyxZL+kZF6ri
YbWTWWK9b2sZ4tGGhur4cuhHYhrBoEhfESgigGJJXktcDMr2HBN6ymNkcntTnCJb
b/w3AqRVYMUwT4dQyA9NuFlMltcFvLwrk2l27bPovh3Jjte683gJCtAeEy207aR9
I0V4Kyzgv3WYi/yFA8jNYLENDH5ShPE/6SwkkJjHar6uZUhIMTNyMEhdmV64IKcG
qD0Xl2MDjVG6zrigETxyUMuLSpY2VmtZaZeuWNUdwJAReraalKVgrdp4g848q1Dl
4yvInyo817TCWLLNsRcT6hb9VLRA2gnfaxVu7wYgzkKb28h2+3LMTpatkQ9MM+9s
cllckkEidh3t3nxydye/QM5+lH/B61WveuA+Wn5CINdMH1jKSKWjX25rsH2jYODk
rCnIf0grPvEGFRUa0m+rklQehr1/ffpL/fIO7cTCoXWn4wBnrrG8VlPRj46JjFjt
95UULFgJrWJN3/WjlxzD/28pAmhHc4lGtxIAvVXSL+SteO+jZP9ih05bgPRXmiCJ
dBfEi2g3pFiYoP/HfVTwjPSWjZKF3ch6P+0ldNNyVhGBvsQ6xm4k2Kb2pGoxjV/P
3z1vkTa6DoeDKyGuG9uQtWdKwSmsIO+wt1/HYDcdxMYxq2PB5gIU4V8wb8Alm4ex
7guU0VBMs6KXaUhi060FCcMXqJKAUUJpgAcqAz3uoRzt1pANy0anQS300ARc9DOP
y1hOOjuXtCRSRzrJ7f8n3UFCCOwWp+F6uw7I646TARI7x63gyOwP/I2g+S87GhZb
JvVNcIQH4ddsBuJTpPpqrojday09vk22n64sUgpEeSzb/3By6YX10+N5aWtI+4+1
l3MfiArY2wkhg2FcvrJDulz9nh5/wipgVhII72xBEayofYb8wC3j9hjJvNIWN739
J+R4rsw2KLwVw/J7AvM35hpNcvAVCR8s34CKxqVZaOoOVZAO6t9pFMvhvMZrRdUl
K+/iAyXABUJrFTHBoaYHMV9PlKilSd3VoyBTUHTN2Zyi9cd2v5jvpqY4RGE/cFy7
fLN8kIc8aGMO/Fca8YuZV6vGoh2FXXsT+WH2Yr+J/KmDw35ACFrDbWa3jyTczj9q
4NopBE50nOD3Ff0KF2TXTeiY50hlPbswpREatI714iELu0wwABMmuEwg+hpxjcwp
6p8CpQ1XPpVP5qEsbC6pzkhAbo86dKRpD7dh9kdgSGL1mO4NfQh+hh19G4e13AAD
OK5rYywno+kPyfDNIVwmdOF44IvCM94Fi1aOFq/LUXCW2Fdq5Wc9uivNCVQOkCOF
JMcMzQDQieBcw1wLi281pHpvXLbfB6PZfkeNIO0DXu1oZc54GZzXDJuzKTEfVBmj
wLKT37NJgT5tNMO09urk9qpJJG18/cIS9h8U/Oh0b59Pks4VMTXS0yFqphrOoFtp
tA0wv9yhU6ammLwgmN+2dTKObrnOEMh7NK+RjnND4FcjJxLj15s4Xmd7e/W8VPnm
ogWRkTJJ5wVdHLQW8rGLCrgXgkOmu0ByeKUYey2hxJguOvy1odH+etrwqRX1Mx97
eECH7zWMjtUR9klL5viEJl/N6ittZzXl7vMUEbNns+mMLdg7/EhjaBs9bOcQG0VK
rpLvFpE9f/ooVBeAkPH7l6zAGE5vs4WfDf7uSWgVCeDe9xO+hHk/pS63zaXPWjL6
VslrPSQmD7xUx+/XvO+YJpqSnAZX9kSUAC1xfs6W7ygFMS09L5+xQ7f+iT6e28RH
u4iYcXB44NtEF05Oz3q+6o/ocoyRd9jZZHNEdR3xlzo1+15uDsbiVDotUMZpRjx5
Z5GkU4Z5AsntF14ljzPFpNPlnu7tLUzrFmtYenMENIp2wk/iNyDfG3pw0sDi8gXA
v5mrNEz9brDZOuitTfZhXstiagghNRK3BDg+iWF+rFWDgfWQ68cEWbLvwRzaew+4
5zhXUjV7znIs+XnS46y+oiCGRWRr9LthRP/G8Fm+jTgHreUWXBMECXsnrgN8lP/U
2dlFH4BJGouFSoifbYbTJDa9ma15rImpRDtkltCho421H9b6v4gOmeto3l9PHwd0
GlUoUfkUkaiL1mLjZYIXMbq8EIVL1ijOXiTHSCcSP8KxZ3ERzR2Gc3CZUxzBfRlE
sWwhSFOHMvKrtGzTLo+fcajc6wEV28k0kBA1MKa79HVjD+/JTLSSpf/wGnPWRdK1
6uQhBXzDkGx84w2A5rk4EiaiI7jbvt66ApRXkW1zThRzxe1onyySIRFTaGamYgYL
T7w8FjuGf9RGjTL0KWrObipWf+mHrYgTRvKDsUdzgj1DvSHfl1sdSJEmP6NMmMEl
V//9AnhhSdoQPZsXnvZlfVFFg0MqZC2DCo+agnPW907zqrp54gXulSXjtLXEQJ/j
uicgD0A98hh5htv+03dvide3ZOQ/mFRuQg6SF/ts9Vf+MmOi8sZ7+rwky3YXEl86
/DoH2/jtsy/wbiiPtV+RAkaADk2PHBqWHRJwD4Rmfy8UbEu5kqOQWfwORh5Opup+
BeLGZ0MWOQ+zwZtWpZGi4ivDgPBw5VyOqChWTeNnGguqFFwtWCQyE3B56rzwGXy2
rRKBqOQmb06Yp5QoJ7QH0bNxG1lgLQFaIA84Ao1UXiu984BNJfpuZgP/QwBxf8m9
GivrR+X1OL5tFHqfWSyv/H+/jfrVlZX+Xp9knEku+1N5A8RwHMLDpBtP9JYT98Eu
jIiVj0IW/jcLOF1IXWdAXXK6jE8y3EKF3ndFNSe9DlOeyLeUREzLsYrmDMGqF7bF
A7NTs7V7y9pr14M4u89weaak5LqvFeCInZItvCQdVFjUg2xq14T8vfvLzrhJWGdo
RPjMbOeobC1aQPJMTiyGByxANFL8vGfbstdKN25uieo1hDZYAOetfp6ZI2a0Angj
JPwIb8lVm5lyHixIjKdyZJ1z0P7d7YWQxmljNyE79n22Zv4+792ke3+EpuFzjuOK
TrZsSV5BJegbC98banmTqCvdqqj+D4deMV/hjVn6fpTqwNp8+ZZqGuzSEzJjyb14
KI9FONgaThBdBE9kq0Uc7Qj5SRgI1jlqHBOT47kLfFrQkt4V/rLvTmJ5p6r4PjMl
G4ZIDeDoGsmgFj5sNHtjvWCL3LmGY1PVT8A2Q25gY4bzO6VP6loGPH/7RllqZ1Gk
+NHniEJpPkx26qLDBU2vv54vnmOShQOj3KOQVMlygySMcKRKWLSvsOdK86arV+w/
+P4gNcqSdTnB/gAprdp2pQoJL0Sl4LEdCTGyX8wpo2p9CN1ENmbmrE4wDIYYSJtD
Dvlt/MKypL7sYfbU1suakURY7hBoYjQIiDkMViXU5mOUtxPDbSG9X9lUabWyQ/Wd
F3V0T1WTfAa561H34jm4sLhomS1O+erRSFjSdUJd6vht9Zac+1gqzbbhYgP5ZwCY
AuAWdnYSaKdXJNPTBYhbQDtYh9sTQTnW0DvEL+9+zI6Lpr1ALCwFaIEnLXGcQGtV
CXgG7HDKZhwnMae2TWHCRqw79uEEDTLqXiYNDgD8QQnGnzl/wo/7VWAJLy2q089q
Det/xrEjKcpemeKQoDUQoILvyKXXK1wPqM97kYjCgDsBPDR52VLlQuLr55quOAOM
i1sdorFcwukNRrv9vMQT4qHb+s5NWlIcWXhi3pyAfVqMpqEbD0Mxs0E8JbxVnVlb
zPLiql57ralz7tmr1RH/oiq1WdWjbDDijYC/e9HLx86yLPRN7swnCVFF+asuWPSz
nMRc7LrtbwTMylPDErdUxtkR3OEQvKC70sMCh5ca6eMwwSUeZwsveUbuXah2Ci6i
bKEP83v/UCRiNvrsX2JMUhS4f+zSTyQNrwJxH6CWf+ds5y1HRs0UiVty0J4i5eb0
IrijH2TwIcSz/CLsm0xX5+IGMkFsPp3sQv4tXw2VzraeRA3fCQXvllZ6Et2j11ba
E02bOMiB4rNLA01nyuCay4La5w35/JKIBXmbHQgtAxpoiryijWamX48PlgU0eKGi
UK9WJoIiWirhsGFHuua4kVSAMv1kn3JlnS5SY3Q6VCefVtJo67/VUjW3L3OCuOoF
BM8L8u+J4gmIIUJerIcLYsBNr/GMro54DrqlwuuHx8dKt+tJT07C1TA1wRBBXu67
5/XbXIJIikW5dDo6juiDUSHLeSynaqNiFbPV5Yf44XUF+nwT5F9iqQkit1H6AYjs
4cljw6s01xd4/dBtgNFk1OLuZCATHHpG7phU0ZyZJHWyvhnPEebuSJg86CsYN4cj
9VkY2ZJz1keQ7+nAxpKNfUJpz9WLtf1GLiaqIeYOYoifPByadC/X6uDjlJlF0Xtr
fsJUZVkk/VQQ81KPgXiUdq01DOJx8Ji1T89BH0p4ZRcx0AMFI6WVwvRIsW3sLfpo
UPcsa0S+8cggWfsbbzWFvUGWNFHCbVU3BWZYBrSwmMtz8lJ9QZOogrJSJKe0CEGt
9VgzsKkF6sNj33tGBDGxY+vG9BsbaDKeca1363w5MZQKZBSuR8F0XTLP5aQu3Wno
DBZZpNGUwPCtyIpvTzEoTJ2i2IoFA72ZSOUl9wd4fc9P57667Nm9jPIJ2b+1lfkY
HiJFMa6tgXPYDiqneOYTH+8LhnwifdmIOu02pUzvBeJIPETPFDGYRaAVfSi4Slrc
HddIQqRSShNcIMabTHc6vseiXR+1mnUnoSaOfu7DxmaSvR49VfaIm3aYcdZnWk6f
Uvebh0cOld0koUWcind9ArsloRj+Cl3DWtYXy+zig6J71qUFXK+BWchFnalaZkqp
s4ADaMTNoPUVfjeEH2XyiK6x8ElvHtwrff2uqpf2ArZe7bZuZz1MGFNVMb4Zh+yv
pg+6K2nb8/6+gFYy8DFF/J5tz2rA72avbF8ax5RZg6lIDKu2i/gQV762YX9y8DGB
W4gI0WBp8FPGVSnWpcVUhfOFfWIenN7qZub4hksMs5aOwIMOIEumSaEDDefm5upI
MmWcN8VctCfa1G3+2na31JH7yJ9v9rFL55vKdGohLHqY9tesn22Q9QRxqFk5fPwU
XN55b+iePLhpg40YxCN3leVyNNCH4qlvHHZJScOX7iLPwCQSbRWvy4tmlb5jBp8C
ABzSU+N8Qc8FU4yzfuy+9okFpnpW3ztF4t26TLjoCsLlKehiiNb1Cj6MZ2euqbuY
No23xFAjEaHwLui+DAK+fz7LPLZcoIRttafVFNRNG+cl+PSAm6xwSmu8UvJpdjg0
uSfsK55yThdbx5phDxKqw2bEEyItyWhcyMz14mRCNDbUQQGjCvk9Cv8aznrBMRl5
FfJIFE2Oi4GbwnGW51F9AoSQ65J1VIm0BJjeRsTZc2lJ06a3KOQnLQz8peMNK+zy
09yN3RueMeOpRej8SYN4pf4blEpIeAKtsi9VIfFV8hPfVrMzZqabX8JnWzOqld4W
QU4pSJEywxU1GrWIQ0SkhDKUasZtkzKl+wEOYYHLuzGHb0NhK9xx1+lgOMkpM78Y
JUEHclUmSEAIYfopf8AtciRV7dkWrgaN0kE4KzN07V/w5yuOwFebOnRqfLb1cOQi
BuaJznvTYU21moTn5K24N4x3271qsUc56eHTqeJsIKZIEvYHeS8tSNN2wl1WO5Mk
KiVsWMlNtetnvfZHapE0NYHqy5nLMzQAj49PWNe7fro/k4w0VC5JOGQeFO5gJTYP
CcwL5W6VC7MWtT2M9Vjje1M/hFHll5azj0m5wQIhnB0XXkhhx+wAkoNwrf3myxS0
l9kenfUya325OY9DvRmZjEIgDZxzuGyheagtCNN67DBqljv/xmZDex2LrTWk09vy
AoEABDklxA20dssQGX/M1Mn3ms5o8h4nNLMCqAvGBgJ+pmdtaXrHPOGTuwyDNjVW
exgwnAYZKBtRU1k5A2n3BjP3SwALBKbNf04IIJ89n9bAKSzvI4KPqU2ZGqurc4me
yI1I+LuSgraIZ7DRexBgQJs3qQb8M0zGboY0003Xiz9dSXzAgrQJJzxIONLZL9pR
6Ya3+Jly3bSF4DlHCIY8UtsACrwOjlThGZcj6/aRBH+30CD5I1ihPs83YBgKn0Rq
ECHTdoZEzErfkjwWfNFqPxW6aifZG2ghhl1DHzBpbV0T5vrQG86CQwW4QixyWSUN
8jhvH9voZBjywx7Sj9qK5pusn8XSHIcHvhasetgXdGwdd7nC+ZBcy0FvT8LUC4k4
U//ITMwxG3FMU1wLE3eXH0sbOyHiklWdKJ1/KZy+aBPpwjEUbSUU4Dz/+F9Rd0OD
fNBDBCw+cPo2Ist6PdPQ3//E1y3TzZUT3M6WaI/t0GQAXbOgJ8aKOlNmCQSrY6hd
bBs/aPTRTLk6OqDsGOVTc/7eFNa9DnbfnuYHVfjjNipe9jAvxaeuuxziA8QFk1XH
p2JcseZ+krqmr9eqGY9/HSWjx73Qaaz2fyszLaEWHDj4P3/SKUAyhBRtMevgzoq5
SqBLw7janGD65ZK1H0D8C0vxlQh1rXddfYtn+2p24gLJu0gxWr4cvzleoLHDoIqZ
Yy5FYcHqzixfTGIizTwcxmC3jlecLuqYrvrSVGzuUiF57QcI6V8hT4FU2Ta3ZwF7
WQgDX6gSqQDx8FYFT3HxObx835j1eV8VmhCt1lEqroHZndbosMrxuDywD0N/TyzG
Ea4zpTB2+OiyzYDHrmoLhZSKKGpEBIwZq02yiu2J9gKbx3G9gGN06WPK6Y5JiPZm
MIE3sf2Twfa2PbNOGQy/7StpxB7HKfXE6Bsr0R9FRoagg89YTMxJDTb7uZKRs0+M
AcwUHBsbyrfSU68dF8NbGG4FcABTikL1rj9O4zNTj9SPq+vaICGR9eqOKaj33SWy
43znRYhymnErIvAcT1oAYxrs3qe98xEf9+euRERWWnRY/6dvTdlTRuhtbUcpyQd6
iHRsk7l7Fq3pfQzZi2JJObrool1DigUTZKxWre6zYInanCfShm9VQrrN9vVe3a/T
QknPF3VU5LYX8d4Mop0H03LMYwsi4ysqXRhe7KpjaxIydKHPGmGzjnE07Tk4WfsX
3XFJCW6eQJXjSzD0oOLX/x4P40MXZPakA3HUXH4XSi4zCFvEPVRHIJT0f40bTaB9
GEY43fAmUuwklKJ7ToN76E7yKFEbU4JOFZs00g+53514izef2/L+o6+Q4poqHsz3
wbQTE/8BQdav2v7aRE/ykoDYVSzDoZ85wWE4f2KF5aNK4eCl21hFCvUjDPt/QhoL
Pyy4e7gZW+eSbZSbVXQ2DWq4VcFxgpSg1cRqSxHsibOaj3ULmED0dlJ5ulQK4GUC
IV7lKX3dXbQ83wzzwg2FgWBPQQhXJqje5L6q3YypyIcLQ3aef9Xm04yc3CKWJR5X
nbmXex5E50jEgUJTtS+9zuTPcmkzXUr1O3QLi+DhdYwVmGOOb3Z+duspGZRkLiop
bJlV8cdh/1XhwJg6BTZM8DNE0fg5yhD372yy0FQkO2dBCqKzIuqvw83LfpaiZQr1
y2g60uwdk8lPTEsJ3mZWCdyE2UqboeUzG207J7/O40hOByKowCgPWXpJqa3MEE5d
WC98RRU0fSfk9OLlwMF1tTqrjp6LZXVCt4UpWvyTHd02IVdSOAYrIlt8ZuPxj6BW
v+zH19Ae58L/7kIa3LisJMoSDXnbzByMX1ThQHkuEtgQOkkj5ji0Attgd/YSTIxs
z1KXf9GbUbgbky2Juv3talgzoM6tUZU5TOQmYkka2XIgj35U4WWzcVV/xztBvdyr
KDuhLLg7QJ83u5D7ryZj0DypGf2OFm8x/7gtA/NHcVxny4Xg9UJH97iTdAa6MKCw
HnCFo20P8rvZb1KNUd+EAQoqK3xdFaUpMEzc8EK5U40AJqJ150HRQNWZIT3tW0fg
ovCYmY3fiLVuaCi/Xwniyly7XRjGqB4j0tvLGucOeQv0z1jVeOczrf43ogqWHnE4
0Saazs5BHy93CFLvJpQ3mr2xhRB98OVYx+7Vcn8MLqqCvTazsS+YbUG2o/Lh6MFo
u97ber3FpXmMrJIEYPd+sZb8YoHvr9cUPqklBtF2jpFJtbrnAJz8GkUfotjxkLdE
gocnDlOt0F0EoRL7F7Sx9vX+3ll+AlvfnTch8P1GS8ZSNXTu5iscXBxgZVZ/fjcH
fj392HVj7NJFFMbz99zXlTDHjNF9Z22cK3vTQM1NsY7zNI7WNT1nyvts3mi3gJ56
f1wcArFiNzHPGIFQho0WgYrnafvp+q257iT7iz7SMugDqxpwSeELi+nnfNX6UUqZ
i6YBptWHvwGEEJxX1w8p9I9kb73cXMiSB1uKxBlfEtcRtd0QBsCc1qR5+oGLWf/u
J1XLz/i4A8I02q403arNnSt23HeEKoPO+y0leePE6Wo7ngJTB+PSoOBB3vxojHUH
vVf4LqIvq6pmIkX5uUbtX8X1ZMA+l+MMKJDKfXVwL0VCUnSGLDrMa1csb7q21WSV
uWUYZIhxp0ssxin7m/xHNG11qQjM68SvzhahS3p0yqt+P8sSGwzlTIpERJ6MFVho
IdJwLIloizOH1aL8eflNbkt2ikZ8szsAVHBiDG7zuzNtJOaO4JF5c1TCB5baBwfu
KFQGAyN+6CIdkWLy8gS+7pescEEZULI2hBph/bRr9p7LBP7ed3BjtUuElAz0UkTf
xr73UuywyPgAqfdeijWkiXRcltfeRBQXt6AtMNjMgkkBQUeVPcviaNlbuU5FNyWY
pcafuXeBU9u2Rxw2TL/FN4smm/pcXYRungLDiVvWmvwHuLtbaockhgbLi8akQaUT
APbfCoXDKxRx2oNaDhAfzfFfI9S8fNCr/eqvyZ1b6I1qj8rsYZVTR11u2NX/D878
DOw03TSVzMsaBYpOo+uc//zZ3U7DCCfbK3PJ+I0f74TNc3Y8zqeOEf4KnNmw8rxl
2H+fEUOP85wECt46BZZRwSK6jZKtJTqIZoeGv0dPpnTTI8Sd6Z18st7iQ8U+HMoc
E8BrYFXPbe1AuvrLG/fFbaTlge00bfIVvwG/VzC6RekwMSui4miWXfHZV6JdZEX6
vEGOKztU0FsITbZOrnOmsHnCsI7pm+q0Q729/PiCCEYdA/F1TPtv8tBwpFhJwGh0
TfNk0ZvCGOEajVwG715sMuNrzx53oDuhoRRI6pzSG+koo0aYkgYHqNFWylIVqQ/F
RFh+oj78r8KZsliPip77/dp9sHF9Lo0Waz5yf6jveTU1po8JIkvRZBrIv79uUAs2
dUNethu8wq8+WHDKbuHxZQcPmMsVmONnITR5QMdc2OqWO2xLyw2vv+P/EZvH6P+v
TSfmTQLZYaDRalMDZAFhcBnxvGYlREqG33e7mZzZpjU49GZakKlbEEOj10BmLjJ5
gWDvBMHnHPeH+RYcmx5cpINyeHnWzmQqxMs1urOnJ5F1Y6zfyg0qs5kzrnOLQh1k
WkdIcbep+xYZ3qGf3oLuSNyDDJeIFl9hTXn/jjDPnaDm1cAw5HCLySNU1I37EjJ0
Cv3h+manctmQwaQE1Pmhq33+gBEo5i7mRvDCU8TTAZM/PyMoaKB9Wz75m6issgo2
787ez47I63QtAX4Z5X24318ZySQ+/z904RkaL/tmOazEL02N+I68tazbxIYiHDaD
MJrEpD5SNgjl9fAV/ScLgzTK7IP71mGxK/A7ty7UkEiSLtf4Hij8FpEReGIX4FmP
6o+iIvnPNQXW45qnSjkeB5WETe7YHK7abU3AjC7Gk0zgjA8C9o/q+k2SgkEXc0fC
8Vs0Nglaw3t6WoD/elFnyWfDpMgRGtqXlCWlUqugbFnSDW8Qyv/ETEWPPpJ1ddie
4Qu/8tD1py9KGJ/nMo8+WYaYoR++vfCLElFvxi7wy0tMfv/UbwsKDVPN9K+pL4Jc
e9dnFCCL7gK5bS6lTVkkcYkY2/QLxp+tM/mmxHVj5W1+dKiG4EIOMDMJQEmhxlU1
qMKM6WmeYvcXIOZBglWPVu3J5QLPTTN5mbN8p4XvUGxw+Xhy9mWoN2eW9glLHTQk
aP6UOkDRG32Qk5SNN7yciTObMX1yioibGb5Pd5G1CAzZtITVy+AnosmFhGqgZl+e
mT1UjrLnpdZ3WXq1RPCOtOhtrvZnl8zemsh/l2tAXNW5oQc0b6mc2mU+O9U321Im
5FlGPBeK4EiJpl0dm3NUVk4QGUVJ75bPHqRpOhK5o25zY/2iqO5rjuxd+CbN1978
PzHhyDHI929W0sX9xqZ5ecAKK4j2NMXs7cVbhgYX+6Pf4r1qpNcwQDQmGrku5utS
IUf/E5uYyPTh1fE+bO2dV3U7FUOx7L51J4221FaDjjM4+F/R6n3dSLDXZ8uN0Ds2
s7n4ZRMMRspffHQowuXKEjKR/Ato5lOyyGFRShurQF9b561xZniL0B4VgTLlPGjc
ik1N4ELfOt35qNA40DSBeKrltgy9y7inPcQifNDvWRSG8zH+czDfPNy4Tye+ClVR
Wk3HmSCvprQ5ASrdTVALqQDlS6Q3eJ36vZDNk4uSVs6SC0ZrikNlzasduzRJX524
tqOSfLewdp7Lg9Jhk0TI7PT65ZAeZ7sNQ0FFZhajK4bRpc7WjE6FfypWLIeZ+aIf
MJgJNE/q/CL7TzejBMhMlIgdVkj5EdEyiBXnAoc8q3YLikxEKAoa01O63ZWa1q7t
tfzk1+S7BIoROle3lRXxfmq48UaM82m4pdPSL3/TcT2IDXdiZVEFp1UgkCsaRroZ
5FoHkkf+SdJVDTdgezjMt0k9FENEx6XWVnKravkKchnynDFp+YWkaS4UJgXnktCW
QUgnPuT15+qP/gZUrL8hBhUzT+xHYU8Zko2KzAyryZalCskqtiCSHGP1e1GJ6HYL
DLMcVnPqptCGC7H2uXwgxhoIVboHonBbo4vfyTSd/8Eoth6cG9VCwwIC6kCYFnF/
HTT76qvDzIaI+YFAhjC3AStwDPivgtjbIw8l/WJ02eKLZx3CXuIBDxIfpVPn71s0
bo8YOa4JCX88eRnnswPbXKrBKcxa75coR+DWXt79HUuHpAw+WvupNJj3AvctmI2O
Jxte3ziyhPPCW3tjULXhB/IJ+bQfsczB7zMsZqWC1nXD3h0MGViTm3+4/SN4pgBi
r3gNcwWg8UFRbjgybnFgQ4knajfPMHbpaJu4kE6kMffvPjAwiotvOgpgDcmpmBsq
gextIaPhBZjy2/kn6wSUN4JDkrULoj/bYHN32meNGE6Cms4OHcgRhWT3ad/L4NKw
14trNB4mHip4zYCP4P5PItQb39nvBVYMBrg5jyXx9FuyuRPMahHpTecYdpqZAheZ
5lBt4UvuRLS87xmzMOc49VvOhKoUbdOiR476aj5tG8Z1Jb/p8yJ3x5pODl1W7waM
swnY9DH3l7RsIcFC3aImqH9gDpUfEXFM7JwtzWYjF+zBwBF1T9Xkjtst54/77zhx
vh9527Udqi8ydaqgQe5AJ1oOnMMRWCWK+G/ospbrlIq0EYigF/KJchL037i0fRGI
Wp6AmOz3AN85DVlL30Kj4j7IDzLvC1q8nPd2hE8Tpk2v3apvZ0a33mzUAFzPrSy5
kJ/Tcj8fD+xDHBJV+73cU33hsxfVqY/d//R3khbvh3fT5RXWLzvFQT9IFDSZeMuM
HnbBOLUormp548iAX1XIeNiqaFIhcccAeiF7p6Phhyyce3G3NZ8SQE5Wq0Bx+k3o
Hko4mWsbnhpGAellcERuMNRZsoY5V1utBo3myAc8+6fWIM/eg5GauoRW/kGRT3gT
Js8zwgk2sqdBNB8mBJhjbHKfeokJH7c5VAFzPsZv5flujan4t/GcPO6p2pDyNzYb
CXNpQNsyCK6RvxXhbGi7IB+VVoIkh7e1D+pSG4as4l9qEYMSzZKho3OJW4JNf2R7
oYlf9skCkRVQojbQYLc9PXgly2oSYBIb2ewgYlbSuGr+48oNMpRmyKshZR2VY4CT
poj6fcEFTIGYZc7DM5EsLoGvOS4Y6l6lAiT/ObX2cr0oGJ/VN5fW6+44+IsR+cEM
GEI4u76DlNOrmoHXHKvK6hFDCKcmJOKzkoCK8wpKpHdN8HxdH0Aze9O6wGwvoMIm
ux8EBNSl/PYMNaiSRp0zI5/I25dqXf4iKT9afKfDxhBSL+mtTafppdX3ZZK0gdRM
9y8taC+TaFeryoC7uJTtRJoO+U6TXXQuAMDbHtZ6LdTqZTlFAkL4/d/kWw1dSTRI
17rKUlDEb7hH8cWMlpDi/cnyjRekLvME/CFfVFJhUOTybb5YBPMh5WzuoRoliiGq
KGCgrE3++ud3xi4PaCiBZD5UNdKpImgtqLhL7Pj8gEBh7Hx/zzpulx3+uQZZSkhH
cqe0Tmk+viUCLT+hbWbucaHy3qGT6dCY9r9L2O95r8mueqyRl+i2usI8LSK8+oSx
Jbg5EtgWLi4hDL0Zqk7m0we8Ctth4EBaCNFSlIInPmc/LkfKl9SdGf6wAvit3jVQ
fczalGky3hcsBAPQOVLUSST71vT6s9BHF/Pbb9yYTYgUppoiDhNyg5YqXpS25Im0
t3U+if6kc+M7ItHyW8OJ8+D7vgpkqTWQSS8pFYC32YdYKuWzqcG+Wyax63/lGfTM
r+u3OTWrhmrLTol4OXz6WQ+1Lf4UT/68ok0+4OJAmvOUZUbg/XhVnQvJIYzp686J
R8xJ1U06sTSuBqXPzxEpvW/jNJoGBNJ9cmeGVA3sjxwrI/tqbD1u4/9OESDY4YkW
1T54UQ8BuLImwfD8TDg28yrQ33u0s9MWUTq5ekKq+bUL6Tw7+IZL1RT7MSLNBAGZ
CnmeZMGAKylOzXOi0W5jdK5HMz+q+XwvjYu4JXpNyHGWptyd277d3Xbc9LGNzy78
VpgvxFJ7VtP3gT9rCAGoiWzt7vNTiAge31n0X0yPEaMKnyPmhOo/Fb/20q0V2CHd
whmEiSdq28UbPi7ajqG5d5CO0ivS8fQAVP8ZPdq8bZNZ0pBqw+9gOdi0XpxiVknU
BXWItWhoIw4tqaSiDcU2PmfqXOGPVNl79ZMfGlTgMs7lvMRKTz7d/XsPQ/Rmg3qE
noqyGEcNSNYbXh3kI1VJosLpjOlIr1bIUInnLGxWyp9dvyXqEDIAEOC7H2Y2IcDM
jZP86BzOl+bNHWCeWtH61vdZUWWPNhe5PIsTyR1AWls/m67Rynjau8wLC+gRZms5
pwOlhYXKGgJ3W5yCswpeIoB5bITWoC4og1Q8pHifKjENspt/eW10Z7/7q7K8fyTk
nxR/xpOt1hWDmQDolz89dbNc+qZvYmsKLOmN5hKIaAZ36mXYE/IcFkqEKz3R86+0
u9rrPPm1NMy6LaghdKdpjNQxrT6QKIlU7AO5ypHZtrmZDrvjnEtU1BxRSpD2JtIN
ZAIZ+GZlL5HKj2WUKDEaK8HhjXvF1n7+I6Gg0Y2Ti0Q/A8s96McZj3pnecVlvmZX
FiG5jGCRX4hM6ZpN6jrN4jyoi6tp5pEtVxuifcRyVMuRgylxqTbx16Jz5x3Ex2Lq
yb0qXpdZMN/DUXF77FmMeCjwNUjKHvWrZLpqiwKO9dSNuC2aXwVibef9DUQFBWaT
ilB0F8NpPzEGZJW6jRTHzw9oJQnbYP+1Z/pg2BoAlWv4LXzDo4eWyhvMHA0LE6tQ
4Olc3jWsDVNm9BF+F6r7ze7oFeTy3kUY8NI1HFbJeAm4W9meUL7AkZejx+Tg2iXl
dHVRJz4YJ7rI5LttVMDNPESTHWt03c6A3RjZaWD/JvGYQZPg4PqkdrYARepVUnvR
1hO3eMzgAeQvOcn2eKKqQoZMGiYC3YsLFI0+3gspeXwaXwAxOuVigEBlhpACEegb
o0m6vfEy1XwQYEk+wtJ6NrT6+NsVEoSCilEtf4pSe7Y1CUPcRvNVp61l6QYtUuiX
mrGQ1eWYnL9jBHwjGst6GChjDVexXsDJyTpfIQiigYz9/TU4XbSxw3tj6/q4QnWf
7E1u7R33qrOdWteaHEXST6NT3IK2dUknykWzyPCzV4KHoO9dh2BpIwEZysGkhXi4
aLUhCnM/86VzF15x/vpF8g2qKX2XTVwI7DjoYfkbzrtfVbuykE1WGhmKZvVfuvfl
w2hG14kuJXul73E+IJpAViXWJJDs7sMNoD+fzNdZ+0hVjSO7kqAZChFHtylLkXRc
LuopJcIt4MWBHvmDPVGAwnyAllufmguOeCGPklPTYqkCw92eXZMZkwTIkwJaf/YD
rz1c2Jjvozp8eqlsIWDc3AWkPjFhTZFx9Mmizu4CNvwBakz07KoSJcoFq6fe1Xdr
cNchixWUTMCpuKQZH6qOfAqnNHhZq+CIMwX4kuPikprBuBBMKPFzzGnYmyhyXId/
SIY52U0UX3/XFz3icT1utprR1hPKy6M2K3jyjibFolgFVzKpeLfPJp1XvUMJZjIw
nNRm8O5fRbvjyI87KhUKeAXoDXzSt0lrkRbojbFnGVrO7zPVEPBp1/4qCLkgUHc9
wlAMgezIT7GTt/KW4rTvhN6CsXy9E+ERfPtc2jy2krSTI8PzTKxasOrh7O0wBMqi
EF3e9TNS12QpJb1JdVHnVUT57Ma7JSeiVN1iyS3aJV6ly91S6yKjydI1eefKgh95
zWqvELGfZuLTYHihosX7CUbCKVanplevXJ63HMszzI9cXcVWHOsdDLI2ulUFfyzV
Vp0basZ00TKBmbpM/RRpeDGYgompqXmMyMQUHtFPRBq/wquIC1JxIuFRJfLg0sYN
NqUI5j+hypn1nd8FwLn2Hivo18nY9lwf0AablWVCri0fFgIS4vwXjVOVT8wtj0ND
mc28AEIkzDS2HxrV3DfRqyeI2Y4o44ZQNABq7/S2Sqj8EvMgvO6meGZQrls9fsJx
Mi3J4CMaCxXom8jnmBAV6Q==
`protect END_PROTECTED
