`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ITOPBtTyrijKk7p7f0GRbOSoupRik62I7EWIOMH0PRVsNFzRNnCLLMZqlfHpXn89
sgaJ//xvJMAy75Qru9NdmDB7w1v0PkZ7rbNB1Mjuh1VP0NM9oo1N32zYdnZEi519
1lCkMF1xLV1fMLSBbFmMY5aS021AwT6MsKn/OKMys24LBjyBohcap4kElrcTTdlV
s6XWIqX3nA0u8czGZU0XIt5XEoSRQ/ceynonIEn27TkrxbpCutxxg7WxHLVf242C
9qGnKBQ5wh3dF4e04zDN5SOYEI13FZOnO57lyJmkb/JeuGsI9ffrj01v+jzZHMzm
4IGCWkfUbDAa+i194w3N8xPvkxSBdda6D44JJ/fRgCjnXrnj2kG4QHCv7H/q/1t/
UBjedR8wFMpk0mVz/r9uBoFwOJbA0RQSAkPRpnOdYzU+VsMi7a3uqkORsxtU/CEb
4pfhTyhKGjq/KC4OEqvLT4g9H5wlDLtzcyASq5cAm769U5EseH1xEOJBwLVvB0H0
gwO/LBvJ/Q2FCixB+ZcT9+aDrLA4Pbt7zu/y0fHipMgvCdLcn2RHyPuqHvCrfM2d
zJEe4JYx1sHFby0f+4JYxWoOsF4SYJmkC90H4Y8TOEJX9Q0yQl8FwvM2cMaRfsk2
wKVWrOM9xrDlnjxmF+0GRn/hxZqBL5xOWFXZ9jnNWEyGxxLFF2GBw9Yk83eGJBmj
`protect END_PROTECTED
