`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iXUfQFvuvxXQLAYh8DLsG0QIax9ux7bYSzl7s4xjX1iQYsZW63iI7PFaQ07aR9ib
mCXCEovDu/drGnkE4XIkAZQnm9jI1iWT8s1Hp/AgaSD4iZBPfOLFDChsh5CZnISH
VrZGyr3maURTy1jm6SUdZzW1regY0Vu0SpIjDiKWTKHA1Qc9+sFM5H90LaxqbmRF
n1/QrHVG3kqFD58NjORupgyOJ6Y8A9br+ZF8DSxdmwXLqgYbvyGVnys6S2NFKHoK
oJwxPGQ3tVZ/G+cYfq5fPgrd7qIFWvSqd8rMeZtfVrE8HDbWmxSvpmo+nPxaw5qZ
ncr4XipLil2EUIHkhabk+OJMem8pzrl/6zkJyA3cUqk6xbLhg19bdw7jPGrXIa0W
3nQfU8FE29kZ+YUssFYyzFdH9LeF8Wk/eudNlfdbtqQHbOb0UyJHzwB0aR9j6slD
e1Yd/wUN6WUVKZfXsERXtrEMhxIcW9hpaMWLybr5RlzMKWwvYRsEs36gLq/ZWdN+
xMKkDICNzHZ5Tn6tjwkfL9RzzQB7O7TFVrcQ3pglhBDgy0/Ze7H9smGlhzJYv14s
A3OtmofgyTaRu6YiChIPJUWcJCiBPKm+46DwXJ0+1Ui67mWx19OnOHrNB+ztb8bM
WDwBqKEIMQz3RKxHsAsJlVkOQhIUZuSc4xtLvRX986t7UAyd+TdneQmX49xQtmSY
+IVS8rsrRkTy6VhncZEz3SMRaMrYZT7UpkOJ3vWzPnzmH7guLqp9MNJL8SP5ZGxE
l/N60AxQaNtzhTur+VoMBZ+1M9nsauALqEVdB1wZGlXRkT9X090GTVcCkuYkttkp
2fd/qTiGFGynLPvEv1IdVD2NhysAcZmVdqUe2+wNl2SD0/TKtWgFWTZmo4vP8nat
MvmL/q7negpVdd7LbD+f39NNWAH4hL4Uucrl92nliKxqkE1LBR3qWX3xLpdMZWJo
DgSUo92nnu/WWtmXHx8FV/ggmOsqKto7rPcYF2V514+eCyMi1AOyubV40aEx7nkb
TrTfT5ji/f1J9JEB1NToHLLiVHbCvfBISZNi9nq5TAijLT6Pk4uwg8JbKrLjHIJa
`protect END_PROTECTED
