`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKLv+PyGZ//tnmRf46xp9uO9iFY0AaDDy5oox/yv+0lXXZ7/PSpTjKCACHyq0yj9
MCKbjs0Vn7M1n044Htffa8QbWghMoQ+pzveFHQ65YEMkbl/+qJrkjoeEtG0piy73
1pjJr9ryPNkVld9FpQmYp61RdIDkMvPwfjZd3ZtFth5l4+tk8TKbjEbqe+RI8Lc0
1S4JQeA8HZ8UBVcJT4wc7c6yxkL87S6FIf5qPkmP3JbdHBT4VVbZIDzWb9lOh3ix
jpmjZpx/GI9VvpCZfypeA9gc978YHhjbeJ0YYgmMhkWg+9sR8HHcptxULc7xiygN
NHiYDtPw0JV+n46Q/IAUWozfxKHk0D7H1H9roI8WL8Nv7UyBPuDZm/wqAzxtXASx
x4Q8W6cm/awShElQuQJZM7dr9JhvJMGb9Qod65wn08olA+XQ73keUEWZKx60cmRg
FyrVy3wjvM2Wep78qFn7xd0iRkywX1X/IJ8ESafeNYGDoxA5VAzdUvNciOP11TyV
pWrSCa1v/JvHxxxu6sJttSfVXsqbaAn5ozf413T+WyUcWSTpW2qeIC5iw+5mIMAh
PlZ9pg3xa9JQN/b9fepkpk/RCvp3S9+6YXabd5SKEgja0gSYPD3oEqvX+AvXG4dE
UsaW6LpX3up51JXzm/YEtCLF8aPqj5iHgr3jygyFOthYB7T10AJlWCjuB5aRF2Ei
ER+suxALMjoXs1IkJhM+Vpdl3fMIG9x7WgUghrZVlGQIm8hQJyvx3Y2bBC914PnE
xsNH7as8N9vrxmFgeDoLDk0dNmn4R+0TbF47BByGs1YoYmrwl9nqHGZ6woqh7mEZ
/BpCAykFU0uV4V779r1jF8YAca2CHf4GSS67aww7dDOTs1MLoNOIOJP0sUMr7S56
sJCLxR4IjPug1scTT0RSsafLBvgXi1GW/Nbp41M3Y+ENmsqLqpHM3AKc8qFy7QKO
L1EW2RNY++TIWHJdnrnMcv92u1qi7Z/hEFSrVjWpP7Rt7KmgtSnXmDphv7A1FCM7
dLppFQfRImLP8Zl1kT1pdVF0N1Ob03bNxy8EKs8NQLiPFXrB3v57kmE69HDEaaUZ
GqU7P39OfS8bEpYOrkuPOwBamlZbY6V0+sYtRHIcRr66LPUIXmWLu4UYDVFgFJ9x
6qEMc11lT+zLGZ67XLOfsiL6/lam/eONGs5TVa3VcM8LxrUB0gcKmbFQ70Okgx8T
BKgHwcr8fMKc50x+C5cIvVJsKQhiXNwwEEwrKtoGHtfBmGk/2KagVily0ozYkc9i
gncBaY5K0SnFa+kPdYDOEYmSU3k3ngPCteD6MFHWzqZAmmlMaU5U+BGhDfIyl+40
Xb0VUm31UCJk9A0Gy98aD86LTxeNU5I7kYU1UWlQ6mkaSa5ZbN/Hc5zpA3U5FPPW
F/8bZU7sHbNV2zHAw31ICLJo04iUu50VR+SQB0PZ69oFgGqj7K83MmOFUhXtpbCd
AHrt0BpLzY1LVeR0Ue4wfU0uPqTHs8SqUdtNiOacm25aKQ1MlwxSJC+V8kiafs6A
h/jNlrfhfxumdRcg20bdJ8IrmqEIf//oVyMymTwd1vTFU7cfL59Ygfj700H+WbQL
7iAyB6U19xH9N0Gh8P4BUKwe8LlN/bwvYcNk/OZUDBJpZMCjru5vDg6TH1IqR7qM
YP8AM6i0EBF1cxt0MB51M82qRRK8jeD/O4yWA3Y2x1JfX9xB2qDP42rILTisPfEJ
+R249jcF3qIQU+sGf3lL5RJV/gsyXL4TgJ4lLqVk1rcaISJuyTBjeox7U0WrmO/J
RTCk+RtmGnbFBg5GIE3BJkpzrpyLmLe1QqAYJBUWfcL6BdqwxUz8F2K+nmEFV57+
pv/Ul7POyNSNmSPkq982PT2d5hCb9NCCjtDRcmqX6hIs18L8Ko5lmivUClo4SYai
pPYGvIZWiqtKTZG0GzKZ6uYICG9I1L6cFUQD3jc3kQXxopzYbY4Iwy18HS3O90JR
pdj4MiGO9FzkQrO6wH8EBkp95oPqPmRMWQGvrImrTi27oluxV32dqjtegp/wpowT
XDUVwOoX+4o/HaunSjFxq7zmU4BdDmmN8Uwpe+g1dtXXGRUMxnNYLZuxMhi8cAKy
I2QOeE2T2SG0SuBc9k3g9QmPtfOBUI48wodWi5/y7vwDOj7xSo5ePn5zB7jaD0+y
yi+OAXpqxgg6pSSXWg/RIx/NxE/wTGO42Px66pxhTtMkob+u6N/z7E9FnSORRnDG
HVpfH7B+LmXLlnquE+4GT8zGPnrPyxeXOBCCx/MkW/NDDp7l/5Q6N3Lo1zxzV9NP
v1OejVk3hjLjyWXGX/d4Gd4vaGOb3sj2ZbYVvOR0HPESw+zbXAndLV4P58/qfckY
/hbuRmdXDUlx9vNpxCN3raBU3ue1ip4XpEXjRwmO1u1o0T2lANzNog7akZoldyJr
yIcFaYFGEeVbOTNKVdXP5t4BGtQqyEfGs5tTBdU6BfwZbZOz/n2rvHN6em1Gt/yM
FUVVBeWEjv36J3lnNGCh2Rp9LMBDb8aBgzxm8aY68ES7zb8gZ05fBepXVWIMsrA6
juZDbU1m0zPoO/lP+ynldwNwvTVoFC727d3aZjt6vltGwoag3sGdSVuN+6gX0teb
YaVOBYXrzC/EClc06VlTTdTsm9l7ccg2X5d3U/BxK1cazxBKhUsIx9cD83BkZI7G
1SG2lbrkn6exjhXFlbU96AwDervoNxmNPJC+WiAlGkVhZBO0wFWk9A3VJ7Vwo4/a
hygpQHmH6gl6rdSfHdlq4HSa4BUgsE7jrLC+0CE4WfheYeBd4ht1S8FF/wbcCiP0
ogN7Qe4kYb2TL6PbQB2YIBhr6EwiORVffsRNJPmxeDPu0vZlahiHdN4Bn8hFiRFT
29Rjd7sSTHIzgf9sTo+hODSiaXkq3kChrP01Z4RmxUsYqMVXkVLoYVRTION8iOrH
oDbruS78XKa8upry6L9VcsoOrrVrTasGFx+9/zVs7HZwkjpu+4fz2w1V1PSCFipY
A+59upDlDgnzxvleZTxaikCWo4C6yR75/uweiIxAq2ysVM26WZmmcAbw9xZsy1S+
rWt6f9Pr4V0G9HjSZtPQBsmh99weQr1y05qE+5vgHbwx8dF0H4ltCqc1Oy4wDsAi
ZeXPMziKwf4PH69cHnBYaj+IPPNCghdqyycfQajGSl8fYFuHY3u1FjAK4Kkk7p53
Ksixb4/cnHeOq9TIJbH3/0BFWtknIqgDat7+uTnTzGs=
`protect END_PROTECTED
