`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78yuZiRlmxE0RY+u6gsaYjbvxyxvLMT2Js+ju6ti+innb2SyDkpHvgqIeHmf4y5f
7CU8jFSN2K2lTXI0us19LjiZS7WUKdMd/3IeagcDAX5K0gATroVtfeD+yhz9O/oB
pLsP0vve3Y9//TOTKWeCQH7HGxb0WCvJ53k2VxIxdexR9eccUk0SzKeymOKw7GIN
qncdum2oKV0Nay3liadXopB+As5MHpOUO4He6dLIzcp7n99pHOoGwAINyDNqV+jM
7e8m2O7aVeZeb1mjxW7qGKc1BnansCNCf1Kc93r9qWB4R7R/UggKoZkTR4vVRFSb
Gfv1MFwAl90rHlIpTZSa266wp9yXKPp/cAk+rtDu9Kf8cHdI9NXsqqhOau3x0xy8
F2/ZwU+OwLgSVQiQvli7g6KGJ7ilJJzIVEF7/Q8pcZ4hg7Lqw2cEut6m++TFOWDI
m4GQa3wQeabiGajiKNZppL8Xuym2T98HQ86HRe0uDbXm6ACI7PZnWUCjms+aZO+0
LCgVCqjFWsp1EvheKmNWFYpmRN4BKfHz12r9mJNmTGmoeRaSbHm/D8AfotO+BptS
uE6hb+VbCRwJg/yYTVwJ/Wf0MfR17Cq05D72I/n75/NnkrrisaxaCtuMqiBe9eYR
Ee/8UxAYDNOjY1Hr86Q4Bi7m+kKxgFXD2xuJttt+UWNz2H541L5dmaMYZ/oA3tAi
HuiXq7tRruqpDSX5+7lYIt6cUzFK5mlYRRcCORwaX0DWHzcUM94VaI28IFr5VYpX
n5ws37CZMkSMZ/6CiVArHbmKFHunYj92g6NDhBfSxu91+4o5f9G69SPq6kHq+zOZ
wCLwTJaEuYOJDccY1cD2f8eRWfEy+sctxvOuglUW55vqTXIP8zJTRodAD6sXAX6x
NcrwI2jHyvjoZfHysRLqKHA9jRY72GdmSX1ybfUhssjUWTlmvkMzPiI2MpVY8u3R
eKEXJXZVAsjSFTKZ+ZSUrvnm8Yk4+DCtNuojv+dtUnTeNAQv6UIiE6Qne3mahql4
Rh3ccIgT56mxkVo52C2mjecEzu9JnP4eyhCpeTqFG7YdBjAD4nMCy7Xkii3V1Vi5
PXaPSPlJRu06yr5EhqL21233MyKCtYXg932PNght/3xm5PajnhJqK2xb6b3UNGGB
NeAcRyRfh0FrPBaEzDdiY8sT0hr18ue459SrWbyx1U1IShpDzl9eJ7QTCSibEqDN
EjD/dmXO5gD+yKV5fjar4iuIYAuHf7HBJu2tgwuanpxPZpU90vn+0DTtb2PcfSAd
WzFMjxmwUfj0CEpXCTzFVqWrjxc2PIhhvfBcHGzSMPXyhteDvR+jJ79lEmEfrXHB
`protect END_PROTECTED
