`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mtmYjF1+IB8rFX46yd/ed9TlsQ5w88hAj8pzlbvFjTWWHr/kozIHdK9HbiG2uWGx
Q6CU8p4Xdohk1apJFKiQ1JXLWw8eGOTv4mlfEGOxpPnoKEQqsUdYjWcvT2Xv653k
Ki3B8QYQhh9rUbtKdsU8/d6pSn1cY6mDPpb1iVZeF0dGgf5SJcw/dp477IPb9zY3
BwbM5UGvbyKF1SnvcaXnTlf7iGrKCG3AxaHRx84SWZy4RYLwc4y9bx0Gi0fOHF9y
hiTPifdq0cKZYopMR3pYyLIXaNe/sTW4h4FEZuCfecLc3kvXM8tUH3BcfJ/b7h2u
6YhSGmW00lYsrzlY//kE3V+C1DURzxjQLq3CWeDnZMAWgQyVz3aD949KMztOIM0e
y7rq7z7sx+5aClq+ekfTMqBrU0x74UjsimVXQn24cu20qHDgwVesrtcCaIajwDLD
a98Lol27p1kA8pTTy1TW+l+5lwsKMWwrCxWfkKq7nrsohiESDv9S3Pqa6/aF/g4Y
N7kKiKcQ1dxotqgx14AJf301nYLi+wjcqX7y9aEVLtO9bjwwA177luBVzt5anDYs
/AXmjj+Tmn9xHLI1bVLTJObYqg1KyiHMA7oEj/UmKi/qvDVp0HIH54LTu4C7Hx23
RsVZLhgZ3MAnlltB/2ycMhfYEUg38croeoCdHtjhuJCaAENadZMRgJj+IBLIJuzQ
QL56hK2N5aDHacPAaOu7lZYTh8+eefOCKtAHea+e57uu7e7YRPDUSd7VTwAKeZYV
EsZYFP+BHy3VYd2WHRgiO1Oi3Xu2em0W6upL45tiToX/UeUYm+jUsxSut0H7HQI2
7YShxf86cBr6YVaW6kZZWSoTPTGvnlizN/8T2Gu6XXIyxJRnH/wxlmZjXMyNnMks
fm9/ptWunz/MOt3d0X2mW5i4k5WXs9nssaTIdclCU9fml9GAxFEPPo2T8Q7XySqN
zSEy+vSM9rBGF9lxDPrbqRHJ46kahmx+10gGuWgtIOYlusv+1OP+KwgEhKwa/PDO
LUT7eDTHLR5xFdARsB9fApirx5CDcAtkwvg/jUfAlZjsckCiVUBPhTpXqykJPY+Y
ee4q8K/pEmijDxS4SWaQraCkOHXkCtQ3wrgKH17HMVpGd7OVU8HdumCp+7PEbRLP
SOrqy/1xzzfWwGWOl3NGmAzLvAPs3RA+kv5ygp+oZ7v+87dHdikS5pIxWxCwu+L8
/ZPYnEjlW9KeOrADwoY97KVkkqyIS2lGu8x13Wp8xu3sIDqvjKNl/Dtyf3Yzx7h/
yyV7KC938MhCJBVd+QyYKYjb8HJUAJ1ChqWwZ8jf3QCwoYHCwIUJoSMfJR16E0Ca
r7P5jxud2TRN9F3Xj11QhfqW6ofknzS90AnIxnnc3vvuJRUI49RmlSEHPuPNOSwU
tztm8Q/Dzl4K1gIl08C1hja0hLte00aEWye6sKg7T2/pbN0M8UA9T2roU4tezaNk
cmxuXUV1GFBBhDI3W49tGq3RLW6mOiRr5hDLitMd4hHjBko8dLKqKEc5atrhaGcr
0CASuw1kGhYCjhzd7VhPTCLFgleoS4L7lXmHYwIHvcBppsM8jkjC2Y5f32kMK0HE
LpSS3DD5F+1b0Ly0XMJi0U946a8dl4aj9JA6j4l0It/n6dQBsp5ny/PlPVmvOmnw
aoL5BG7JhQaWMcX5dKcmlMB8ZbmM3bSaXs6DA2IsmQB8dO09rzyMXmBlE9H8kX5T
pwxxszfEFUb+KnUIOL0OKikf4DhQGOlbMTCZFSYn7v8IA679wQUOU5IKCWylCB2w
8Gb9s5/+prq4PSvmZO8+gPNquedwbCix38DCeuGkgp2q+eihJSRo06hqgR91Nl7t
7BaWtbDcfhahMmloQ+8EPyE6VRNnCnSGLkm/4WhExEqwJ+NnSjsbJtEEhhRxaQS/
zLaoXPtafv3uC5y4xZuSMfBV6PmeTWNir/ZZVAcNcoA2In90cS3rfvlYFD4trj+9
028jeGTVMywK+eWHfibfVj5BHEmN9ewJH0wrp8sgPXTrG+qAqrJQgW+a8Sk6KR4V
xD2IcY994C4eA7v0+tSHedBxpJT4//FlL2KM+KcFoDpCp3jrpcaQQzr5p5T2hEBI
OfeGlkV7ZlsisFypimYNqZdmtU9POI35dDXGmUy9EvNnz/ZNQp8u2f8mFFBwxBIv
tXDUIGz6fGNr0S8eYji3+ODPG3U+U+/W++W4qgL8i9ANTK4uSwX3dGCa8FsUtPaB
hnZO7tx4X0kbBhdUYPc4mxd9Sjrx3nlxm6fYOXfU8oxpymKFBlEXNHAEluu6x85U
e1hz4pHRPF6AOPzBniPr0ohs5aB8vtlEnDF5tpURbnpzFVXQW1/Y5c/SAqUK4tP3
4DkJXE04qBfIfWj9xmTtUQsiFPP4cUI1/90jV6QFKZUGXHXAZdPVdLi/J+LPjKjI
FdtwJcp0KuI/mwWb4CNhN0Tz4KmyrkkKBG6yEPKbXZAqBTwfdLHQl1zh4V1nMAjG
Yzh1YaxAOC06nb78K8OhqAAzTp1Hrpqa5dU6ifFQoxp1ejG86dhfgut2gDxw6TS+
Wk6S4VS0rIp5XA/1gFO3uwbBmdiKXcMRnphP2wDq1AzQkxP5PWve8sFREaTzTNPf
fGfd/vZMoG8j8atst3H8ewA2mI/V+Uh2ovxoLZgVR4HpdIO61mZJHHse1j1KZ0zV
Ok3m7uv4xCMYwoCAEB1Z81ovMj3XR1Esr/Cb2Om79BOZ4iRdQCGmomklmttaYl6R
xyGsBo7aryoFbXgVDSzwKzihx2p9tPCEJXqz1RKYFQxvSMOnqmWVFlXcWeejgnPd
iH95JyUKDmmYTfr0hZuIPj1kS0sX0HTyoITObJcZJ3PRNdp3s5PR/R/LKddbRGhJ
Rq3FBK0OVP9JDfK2oiNii9zXM69zHl+DWLjNFS4waYe9uK63kkPrFISxYMVCEzYh
D0jxORKrEvZTSfT6fKTYbmoGW6YS0lZ919RzLJzhPFupeqITENYS0+Ute3C1MkLR
vnKYDUcTuyP0c2tW5dl+i78rYHkt/xxNZjBtGj8bDKfPze5x8BZROie8mkZzk+Ze
DwnZh7TQwCnuCDZgfoaiqqSLrElMsDAT2dI8cruBy10CHOqaNvgsPJKa9U0bPBnk
Q1nIwYphyYPcnY6eu7MWv6X4YpsCX3Avno770cmLiZrsHodDGZWr9Xr3bmQYAd+x
NuFBk9TfH+9S5ohd35gxzjgJseExoTDTawXzp4fg5wmx8ie+ur6bpMwK2ZN8Q+wc
Ry5df5+oevOALsYFGCdkQ0xmAc28Feqnk8YuYV9+9kFzurkoSITEa8dbj9uhCaQl
h8yy9N4ws1uqu3OmKLYWSr/OdSaRcsedI8LQ8lImFQemIEOPbtAaF3bNQ4ZUF0GH
n8/Cr8tCiY82+hyPiKklsXUieq6OWX/RpYNJHNfZCmSfR2N9PiE4gaJ2iTJi3YH8
ByPs/3UnqrqDvqDruLUnxhpaAIAUsw9+7sodVAEWESZIC7R2w37o349afzRAW22v
j+u2oaOtWKPL1IgFYds9J0JO9zrZbiYie1mFVdqRwY7CbSdOSHHTFqVZHnTVvDGc
Y4/QO0e+vYDlLNEsW49WnzO74RO+NjUQRJMjCb+yrU66EODmxXRkZe0dFrllSYGE
At5pIVZ42Nw8nvHUMR8lDTaw6JHIqMrWiw3WMWk3E0Ytxt356Y9ODKjdnMHsTaNm
OOpBvy1IUb/SEu3KlQ4xb2lnWWrYYW2DEQFKyAvBUV2wbnKuHIt8dopxN3qfM6Td
v65LxG1+X8XCFAaaw5Fa/x+a+VpBtgja219p94qRVVz/UUxwnBE5Gj7fjktpvNM+
ocLxWC2avTxu/ylLTV62K/wDvMKUU4VIB8CuBeZPF17zElG08UzMOpf94TwkJWT1
aN+f2oiuUNrSbVGc/9JS1IFUgffFODhVqv5hZw+8pz7pT6WwFled0EfHk4LdVStp
ICep1bbVr9nWS52aLXyAkECyR3Oa0P+fNj6AjN407d/t9CC7B9abx4tFWwJvIEEi
iF6DMeyJIfaOnDYjrlePodC1UjIr5GqukeWJzXvAxaFokYUxAqAG5hz2bxwxEK3c
L4yJusy4x0nKsELIP6No3xIFkTuesuYstOJcfiOpm70iOjUn52yOlPeFvtCsGGBV
A+VQ3eM/ENrcc/zynfMibofzVO3VIe38j8ICm83miHswMyFUhN8Il27xcKGR3w2Z
Gg3la+43EH9b8FV2X8gq69r3dEKiasSmEjiuheQY9HXM+hEFbYIRWJyX8eKbpZcP
+pLR8QQJYwDMrZwWVPHUKz9EAsIfuX6KPuZmK2Gua2j6fcbu/JjvCvrHJ0/UL3Ft
7b6gZYVkFi7lR0e2HVCRbZUYgm62fOK4R3W3Eg211+MHvseS/SuwoKQghcP9TAFt
Y/26P76RISQ23/e3AqAgvZAwmNloIkjK1adSUxinRDIHAzo7ZCacwJQ1UARCRJbq
8Na8K+nhCgOwKdFsyqoYGeth0ZRmp0F5Xgm+Jy76l1StDdVxaJYr3dtYQxDvzHyI
E5rF7bA0v8d0FeJLZttUf+RGRNaGiCi/3a7Ll55BS9/7Ks3Y/fAqMGaNLkbT03zI
eWK68bHgUhxjuevz1TM+jcwTwFnItIvtToysAvxY0MIDMhcmQUQ3I7zMw7Ouauq4
k9B5MgYGWmi2IOTM8UX+66sJb+/2l37uF0AnwYN53YbferxoRf2BgdFhd2H2LUoD
i5w+UahSEYINJXm17ZIrDd0yHfaLdviu+EFqUdXk22va+n1iaCeDmvSCtCTi6Xqb
5eRfASb6vpK8Ekfdvpd6Bw8WIobGvVbPxQCusQ64riKJ9KMgsiJ1NlwterEzRmNF
Saxh9OKpedNrHvVKSJuio+nzpNwL2HQRSbD6iVwQzwjcQxyO9lUBd4iRvchR9VbL
PYkSaNZs70ikvtYrB4jVnZ7XQMw2CTSuqaPxt+8ouZHT1XwrEPESjXxtRTvD+Lro
2bqgGMd4fMSchXDi2TUkfdZpRwAe3PoshLWSg9h/ODA7fp7JwHMyVIvQ9xkSn4aI
il1TVYrbnNtbe/IKgLrsFQh/0tiSFfsZ2F+4VwTvuCErUopljJ9tXewv41ohXhWf
4aP0I2FLHSsfQ9CEw4NLEJSs6kPeSmRfEKcx4oEHTP3L65xSYFzPvXOZY2TlgSLh
OpkneZrZvkUDOESBYrYKagRsr5YO4DEXvObZA4DXFUjsiumGecET5VFmnWKfDVrZ
ywJsMHKUH23F0HrxflZG5ZnFYgqzaRhSqTAK3uYFGXNr8NqAz2yP+3DDDbX0EWdg
MTGFE5XE8w5IDTh4athbUabfqhq5VSYdzO3IkgFCBZJPejP7Te1W7ZFpynUTiA4S
Z7p7uHORnAuGDEYAw2Xbkog9sHjKPHSKviWLkLs54EnB0YK3Zgzaadz+ATEFrsmK
A3hasDITAndtKvh+0GqwenxsIQO8h3WXBrvpo3sZyuAaKKUlOucv93naKInPpdKe
Hks6Q8opRwLXN5n5oINPAh6szmrX8hpND1aMLCvUOMiXXGbT2MHmFh3j2qculVNK
n4a4BnczWgpeHt6YK3oeCIVy2lmqBs97IH9cT5KSe6K1HD3UK9gyfpYQmwAreorh
vi2vphhyaq+T+To9IUK4KoXj7EsfNLXL9iEhiMslPudwf7Lcgl/TbDxj98sJel2l
+x4SiAvUO1ENYK7AyE5dVaNAdsTO6f/sa+AdlzAV2VidW5h3vJU3Y5Mmne86z/zM
yjjm9OWigijrDDbxnsSVtYcVtrFmLGXjR1rsqSyVNO87laRW0FYQt3BQfCQaVCG1
Ce/+HMnkOMId+Lyre4S5hWGnpVrfJU17jJIKp+1J2T5JzYWzVxtS0K+XqUzCufsk
Wywx/TFxm/vIccBSqCbjCpbEFZ0AiXXXzp9O97SnWlUPJPzE7LEQcxUC9aazng1z
ACMatWr4JrAa6A/HRLldBWJCYQfOoH2vU4Krw/gg0s+deHkrrwHQWJLRcyI7ofBf
hF+AOykfKwjTprWBN/ox97npVriwJjOh3MStx32AB5DeEEBRMgj4DdjdS1RKzUJm
BafHJ9c5y9/HdSH/kBaoMLwts9+7iPxTrjn5kvYAzhCZQIGv5/G6V2Z3fyL/56DN
rahBKNMUNHVMj6gIi6GkqwJ66a6yaLdovSN0Wc21iVi+bGGC2WTl5WggxArugmWb
L3SOYBO1b0NDxlSqEC+pjN3FAD4nUGdDvyp43wCg+WH5ugS3Rfq0CgAQv/iw8gq8
9CP1BxXzmLW9aSNUxnNFlrLhHJDTI9Y1TtWwwux5f1MVE4o/yq/vd+OSCsPChuR9
6P2w54RJd7lN7JutJMUuRG6KvuztxyIPkUhv5sV9G8jr7FxrlCZWCvCrBb60FEWz
9hwCoBCaz3bwHEf+JO/e2gWl5mmbJwIbbrY8CCjSTnH2tqGIPapvA/S28hXWk0fq
lCWiMSQ9O9lZZPEqXz/Ua5hE/9zsdjPYfyfFdEcCbOJgHG0nbXE+4W2NVMm/hifm
0RWSGfD7+jSHcon8OXrPlx7xri/dV6UkbCSPeulsKfLeJvsHF/9p1Q4A5+TxK1L6
YpFGpa8yZVSxqeLWlaS/JAct5U9xB8Et1RGDPc5EX7mNMV/RUrPEvsGfuVc9YW2W
OXOQ/ig3yfXAcpA+KDyOmG/yIjYLX6NbJ0/gjAairR7GKnAPXZbGWJO8X7BG6Fw+
EmF+/0h6PfuuUW6D/nO51uutqx0dU3lsUDtgHQLX1qkNsjXx1LSoAipDEp8iBiFD
smb4N0hvvWnmMLZWKZDPJg1C9rE6qYiWcUTJFFYtU8A+lI8Pl2WMO7UVWMsccuQ0
HLRnar9cSviiGZkfJzNHwTJIoZIZiAFVLLbU443oLq6VFJE2HZUHZSCRxrFEy+CL
wrom82WniRGFOWkPLWSFtpYOS1rU/nNiNhxOreqpoXZLjTjhVKOv/biU2jNADIrC
QkyT1Q8/O471q45sng3FdVCEzUtXYA0SEjX0ZQgPHA6v7IROUFuVp6qRwbqmhkHI
uJjLmtSfSKLGX3FFhdUOxPR21JWiC7wmQ4Fa/uZxjaioCLqZHG2U/uR98iFgWSO8
JIS7eTvnMs/chercRYDTjInOjwGIKIp8CLkqoD0SCjowOc5bXAi4kc48Vs1wEGzp
6t8ZQgBk5KMMuD+pfG6arX96Tt915b7dPuBJ3pBJsWbwBJNkmIP4o1gj3qxVbTJy
Hs4sZ+o/I49NIKZkKRxG4SkNJn/sKqr87ZbAIjfLyFkQRmUtElkuIBuK5mcTBrth
RMt16GuYlDUgBVuUJpERY+LCzcaTF5byRNpZmezQCy4SCjNj3Nxu4oNWhPzbnIOv
r6iSNplc+jTifGHRyuQ4fJThYD2wSRmbYpf28rqbD7OIcIeIAOjVhwb6fthwE4Su
e4S8dQtod8OzVCcNxsrPEQyQMioYimy5iGl8NvURZTC0mOHmRLQqGeE/YTXsEZDW
EzimsZUGsLAPSWye9dBbub+bR0yXQ/+CNssHfKwKG62QtkZnr7jZhSDgo+wre3Zp
zsbEC1+FauAdXibuJA1TYBjXtREtymViBro+0UGYDVhiuysEFxJlfjMq9lNBiEzd
ycx6dSSdMGC+zdzxe0tuGNx6AMp0LCxQfqhH/zYLqTz5wFaThBVvth9h6Go/20OD
PgCYFgpJ3dRF8tUCtbjo3VWz7PMwiFvLjWsALqu5A2eZR2sJbRe0MIDyf3d5v077
xghVTRVL4SAzPpoYeiNZPayPoyQG7kfVzENcd4bN1KV2d3yAsO/0yhG2GcwfSHxF
BPToYUKjC5o/Z/9A0EPkM1t0jBHHH+JyDUp0x9uRTERr11HkqoTpq+d/Ye72xV+7
XOYIa9GqYRnNYh4Fr+uT4T8iNYg0EmXpSH85PvOC3zci4Mm2Joew+qAEoKZpD+Nc
QimebNAc6L597DRxuZcmEyx5kZpdDGSJGjcGxlTcFIxg793+8iRuRlkldgkFqano
IAJxw4/HJgRxWanKyQRCvaGIrjIdpCm4sSc2dmu+VsEUEXBzA2Zmc+P61exmajTO
LVrfHRLS2g7FewsJvqjyELpakxk3a92HT9uMnFvo/Gec8X0MZ2mMkzV9qBtZsx2m
9w5pshKFc1R4u9Fafls5caraVSxe7RKoEwJJahQj1vWJZ38Y5T7bS01LZgG+56Eu
UNhGlBly8vkOOk/Jyeys9DNaDOfPBtYE6+QzxtCE83k3sWHagQol9/3kshchdr3f
33yJyd3BkgOO0pcduqgxWkRn6W8gbAZC0pFwROWJ9rnhqNxlV5R4XOCD2hIYrKxO
tnQMQeCnQJt0ncyml0ihshi4/tbRDRdEvq1ZMIrsM2H09nsrkT9G/HnPavMz6LOs
waSJznx0pqAKrf0SUemXkBi5jGyLDkrvmam/2ZwNbenASl5BF6C5JlC8ZV1PGAvo
ZumvFOqw/E8DqXfqOO6oeyhReVBuGvot5uGeuYsUW1D1AGUw2TgsqrBKRKH65Z/8
lJsuYuxMvHvn1XC9rgrii0sPjwpXVZ2DgdX07t2pWpubaFA5Tocx3urELTUZX8gV
JvI7Ly/0K0MtPxLAE90JUrluUiiDDAoLkXOfg+0ntgjfAuQRudpkFhq/LdqV2F95
IrFzsh97+lRs63qhcOSRxZrH0Od4htTBRzI0d2Mf0rORCFLRdsUHN9MtIZJ7Pm1I
h2HcMxmIuxEYtMa0e2oUFOHIbqfC6WEnnBny8Xo7cm1VtpXKbEdZfH5RUfvJA4YI
dvujS8o7sWLP2DISCxGRXJRV5G9a+YSjk/DTOKlofLCtrhDqx7aBbacknGso/bMb
8EiflEfUPh0ma6emadVfJcyEccK19JeFAvHJSZb/Hnh5CNPdSdDJJ/l1U/AYsqIw
K+VadbpVJW36rBbmBSVXpQZjzQz+U783f/H/2tqffBRho0+Ww1hcBuUzo3K6FYIZ
nsOQW9VfXIZ/AJ4NK32hQY++MXWwuW1y9YUVQ0Czx/lD1SoGsAIVZA+mw57wl1Hp
j2z0FyIlKIOsGrTCnLv896U1hCb67ySBBXI7+UgeDT9IOqZYcr+OE3BmIORqF1P4
Swtdutv4Mjy30vSaT2HAILqn9HA9ttdowm/XDQ3miNtpuTdYnYm7oWI+sNcbRFyt
+PVcBpexnmm5FAHDKoaeshuo9YsEmUxudQjgrUulO4f692YF2yYdlZUQErkeKVk8
lR6no+UO6ewW79hphepvvkIgHnZ/UNs5U7cWrmlUX8TTIW1Ps2yTNLzFYgkVW6h3
Jiaxo0FdUnYjISsOKZXPUzCO1R4AdVN+e7m9ox/HgFeuNHtu9OsQj8+nlNrOTkaf
923f3nd7WFMvZpjqCG13wqQX+YlQ6JNc3sb6+Xv/xmc+SAutIcjhPG0jD/uc3gnQ
nM2pBqus0danGzvO7Ftay5Usq69k68bSc2MpNgfOkkt5Bx1gYW3F/VH/zz55uFZ7
jb9ieRn5nvzpiWSzs6WCnX0Jp88mkhLbsn3lSdwYNLiYA4FQn7+IzImj7aRAdCIQ
3b08kZqdCb2D6lvtyrISRpplfJuYnytqTyCql5CA0QUKpDHq/X2FtlN7yjuamNVC
kTf0rvjPoEhGSAZg08gz8PlmhHKVK1v8o1RJZwn9MW9jCSzyb/lN0L+AC5Wm9QPi
TR2sD/dq5yVf7Tr3980bzHxfW37g7UdPKl0Oqtb9saee/DHkkJb0sNHezry2O4He
OXJONx0s+NpiGyjcZDF/WfGgC2KbdILiWaTVQz9G3MQfhQMXxsiXbywZvaucDH79
jugSM+e7uT2TVk/OiRuyaqiT9lsbM+3mq5JoAooL7PgQWLY0P4JBgZUmM2kIGlXU
6j+9icRJvM8AvLaQwyE5kI9itn0Kaz2rbS4BzRghFtNYaPAm/PQAhlfqh49gUzTP
rkZh7NFE90ney6RrBUwFcDE9QOS7NxQtBuD5VkNBZHaqc8cuKNk8O+h1PO4LgSCw
bcljahKfl/zGP8xSKoXm/PHyQdLO4nhdFdBgWwtoC5GuJDlsp3D7pqPMkVHWLoZf
ItP3Gigw+8G/WustjsWdUK63sxdazjcIUwt1UrvR3X+eRaDI7z1Bx8GK8AUSs8ci
U+2Eqm7gzZ9B9Fu6Kw0TAdMgCXSItntfBFVk4Q+habhoiTR0Xs+h/hB6ZU4LO9e3
MVM/8ltvvOhf9+pqxQveeN+dovjnNKivKlcMZqHzZ7p85aECJt6XlsFqz/vPznyg
TX6jlKkqISL+RoLY9JY9+UwDimwp4r955Cq98gGnAYKAYPL5KPpNuMshEwRZCub/
HRNF9Pt0QvLmcRJZNzqXQxrY8VFIoJwyYcfTV8U70xGIjjgx/uofFnFaqeQS/LEQ
XpZkDSVJTGMEgfTYvTql2g8lgNbvXggw8hF3VVD1IrBIA0gWuxUw63xgR0Hvgh/r
jCr/XatNjB2R/I1WppkiE/Rc4gk+5OoYt36zreiNwi7mY1cEfPsqrmg5F+qVg5AE
/jxttGnpz5+o40qFZLuXmCdQmRZiodByL/0WPgdVXub982zpwFPsK1tRequ57ZLa
XaO0+gQSiM+MyrRAVe/rnS4DyyUsbUTQWRpWUA3/xNfZdhTIagLRqm1QiQvfBJ0J
QqTB1LeRfwh0v0U8NaxHsvqBTeBbVaCcvMKE2Bbj3L54mvKKf2t+W/6k1rnPRHau
pxnNQlgdR8GngcyJHbRz/78mFgUh7nSwe1tFzbLlBfGZ50bgOIBtYG2c7vvbFHIm
SN1zRp8NWwZljzlyXxWMvnMH/y7y9USX8Kyj8vxdYs2c5zuiiVbH+ut6H8Gc4Njv
kF2+pnsB9PuTEpmRuE2v4D3gbjSZvN0+sD1HKNeEUktmvr1gPzsV8uArNiIniF1H
2qeLd+pHzb+c8LvfcIlLq4kmyNlYrOtQvoplzCepVVdm5HPuHwSS4sK52ObdQEv/
qkJCow+iYjCZcZaojhPhsxLm7fYiivhrVrt23gYTTUo/bX3OhYD5K/x80LQtl8gZ
CINJw7DLuWySkKIQPbwwPEji+oqcXY1FNWtjF8Su3HZ5yqtLTDAgAfvd8JHhcfId
VohIyYjhPwXEMfStFCwLSEHBHau+b0BxxA4Cj+KowXO0CxTdY+cktxthXt184CYf
PilbFuMdOWsB0vqwt6/aYZu3PBxQNG0/rMIJtlsAp5f8E1Dzx+HSKu5vqqaChcVq
axag8ibowQdIMr0ojRws/di23COt6tLwqDOFv3cc8BhgU76qB9FJj5L+fSNy89lO
Jtul8q98mdmLVFZQ68Jvvjl2BK2B9FXalvypn9ntmuFak0tq5ioGGKxC86J0GQBS
0pcODiy1/adXk6WxSS86HfXPmQ/HhE0HOM5kLs2zMzvW3/Kq2BHCjNVjlhOT2ZV4
iiNLO14Tuph4wD6XEtn2/49E9uBVolbxUocTIX4Gr9cE1ws7q6ic7XMFYgyMvEED
CHk05thgLW1nOIfqx+be7fFfbncddHe4A14wIq4zUSUEFV0Bpg1V0bCYVtZhenZS
osXKUjyZFwXWDzLkxK2IU+nGh4RuKGByP785+eiNWdsz7TYXyiwJww/dAR74LifA
uCFXBB2wCP4eJaw+ZcnulYD5mxMHCikpYTV1Rj5bulfC9PvuOGwEPt2JHNiwDMBg
QYXFb8TY7Tddm6MVZ1rm/Ao0T3d1yyAdWaVVBmGWJCqBPgTRMC326UwXRxkukIHt
hC0rbXrFBXEhPipXO7FDz/x+wR/NgQfXyi8gtxClWsyJUGweb1NiaKc8dW4nvdfN
1rnUAa/zqR3Vdl45eVA69ABVhAakOT9vVFi1a5cRnKtDxxybhYZU+VBy0sXwjUD3
l9bJM1XRBoQ5PkX6T+HJnL+9a//5vKYT0bT0dK8tZFTrKCnpaJSJ9ybIBkLtvrW+
UwKYNPgRGHqZqqXEibd7sAF+wp14Sor7djXhLVFHI0CTJz0cXK/Bl5y5nym0cpAF
MBOiBoU/eWXbW6Bi7pXS/0D5QWhcG5uiD7nzV15spS2V6guf2FIYjLIBq3tN/e3j
RGdODfnjKjHoX4EltzIGaGrMfILvDhir678/0glbV6n0RIkhUDcF1clIMfAX/+JN
OmnyzvSbyKVfXh3TmsAX9nCNOCyCYCxuswY7zrCRdvMSQSvXuxFKrjKINIM0YepU
EGAIDl6PHy2tdWbcrgkMiJPknhDVjuo/kpM5NCInCWIyHpIAXLtbSob4+ZMvQJZU
dTX0J4FFjHFCS6S/1oSA9nhJyjf9l9xLQeGZksJLE5U5cdN6rpgT865Okey4Z1jx
R2RDsrmoWEurfCYL0dBPf+58YPJVIzfgu/UO2aJzM3c900udVzzBvFxTaBAT4fN6
9RvWhAAp4Ig/TNJtE8MwkEIOUyXpLghfoGPn7pEoK40sMOyuB3MdRui4FWKdUXC2
ByMAAiKE7r1mYvxD3uUOMKX1/quosNQ1vUUIm9vIETCyvtiBEeXVkCVdJjWTB2LS
kSJpvb/g0471YZDAn2qsznSkpff1p0ELkJhoipPx/l/++Jb9UgScQm770/LT9EWY
4RNVuVi8FUmpT+rdz89a1MAz6pWGbu/dc/5Ua3KM1WwJ5XQ3xUttBsJTMvX71bIw
OMC8yyOBZyBwTvTLK0lvl9airGOsXDYYdbo8lJHmBfFAOwZ4KcuT/hAP00r2O6zH
iOHFQSQDBA3GJePjw4h+gvaIvUvCGjb6KYMMg0h4IvEdWSCVUtri/dxvv2GrJwWp
ZRbTyZv6aMDRvjdxJKdTgmPNMwbVyOGkGGm8IdQafnw9bnSKIDeU0QLhvpZriJcr
vyI52s33xpWl/LLdPCmlqKPU0WPMBe6U/BAQBAGxHxnFx5R0Na0u40y9Gq3MWX8m
sBIYbdbmwxGTLRYmY8KLVTqBqwsPkPhjeihb9fOvGn0ybsgY+daVcGwMsi4hQNa8
WtvN4BM0pHHNLCeIn0uHHe7RXvkAvTBcr/y1hJ/5WM9JB8JnUeijvZdImf2u/qFr
A/ma91K334cSQx/GcoPKpBqFuuIKALnmauOfEbt1eR3d/xx/VgZ9hViw3o+tLSzA
z9cLR2sVB3CMaHVRp080klZ1IGnKirEbh+JYmE//kw75dMrFtg7B/BL5I8G89DVr
lBv7i2XNYTLGrmtQb+1qc/ef7TvTdlLAQFfzAEt0ySemC7y292FusGGyWD52voEs
kCt8EH16NCls3o/HSvNTTIBdJfFrDVPr7dqxRNcyq3aGNeexNn3q+ZbbusHtBeQB
JJU+Mu0ig/gDUxPFKi/O4EcThEc1d7fGNgMCVQM+kSMyLf60jscuDUTzFVJ/kklU
TWrIaUzZVriJvVOA+D3A8leGPMyTai8YfGxDX2qQD0E8p3L5O0haqkqPvbnIgqA3
m9UPggVailFehLIXU0RVIF5ffTcmKqjDc6KtWrjMflsZdb+4KjU+XS7cphy5iO5+
q2EZIZQaP4rn669hRxmUgoLChOtzJMUBnRUX2Gt29DBlv7UjoU7iKoATCzLfgcrL
KEXCKvTDbjlBtgPJPKbu6VjxIt8N3pMKkkm7c23aAmKwAvlRWgS94nYJeki4mdGL
biCSt4AAYx6bqYzXsRSO2cpIlpxUjvUwzStFkeADOmp2qBntVxLLW7kuaUAOeXwb
ek6MBrAwXPdnkL0BihgMhDTsMECMA/O3K8pN+HOawlC6+tTU1fodcBPSv1aHRE8Y
seyrAUOJqkIxGdnodSNOaFLvwOSjBYWxfUUOQgcMbLIXmemaog+ZyE5eu63TA3Jn
Hd8u3QkR52B25yRw0L9j0nSEHZoIYLm/JYGdG4qeDCy/siIo+I5k1U5SG1X6LtaM
IGCJ2+rLBFJlMKZgg0/Rwwcj2jFV0Xne2a3rFjcgBntlhpcvqiljdY295ilSoyBd
rNa7DOOcvooMtwgKspym/txfLN9VBWjzi/SwQCy7tCQNvb1ryV8fUd3BbuP2E7wv
mSmGq+DI6GAr+HoEvk9H6LVrzLQaPOMV2ek+IROCjTBCctPa57W/YJNOYX9Afiku
/3GcfzdDL6t8rRy2puEjFiPauIZ2zQgHVhytzYEtTMjtw2TMVhzWVAh23Z6z+BHH
9AjQWL6m4qOBW9QQr0Lx0wwZnhXJV15Zw7Jgj3eunyPNQcDnZ1rv6tEq9QG1T+Dt
EI1hs3uRlrK5Pf+nW/3BbFqOdML8NwN6UL5991fjR7x7zXJxpOrhjT0526YyIOMH
d+vJVaxwQLLomZer6FqHymnHZZhrcH3j9QgbCeZPhLLqJAc5kXaQYmI5iggBAJbK
FGxbs1rdm34LH8KG+GKvnt2o2AmlrwVHqSV01awxf/WSFSjpbXVqrt9v/04GWmd4
aYVGTs+s0/3ffMMUnHxjO6EoBpHywcmChbeviioz2Wnquut8TK7yeD7SZDOiUFnt
ntM3YFJoSEbw5B7e98fbe/4oc3QNOfNlGpaN29dlgdVaEPBbfzbe8b2/PAauceYi
8ORAp3Bdj45Wvsul7SnYBB4+5rz8qy7Cl8ljrFFsL9YvkwTzShvFVt1Kc5fMb6M8
ADjJaOGRrqrZ5FdhLD+JRNCxgwJ8Xa5yEdg5m2SYaA8OWPNf1VcCFUib/NLx9zWa
GSKyoxGzjTgL50jMdNDLS5AKGqKG5SXshUGocnTyFtpR3MndVK8l/Ypwu5/Ed8I9
lrySdMKuYVdx6tRCcBunz0jtWZQQGrK/+dFR33PZJnopZxrUYcujz4keB+Ba9cKj
D8BbzV3+jSmoAE9VSFEkOzCP81BfK8T3gu/+QvINjCHWm+AD/h617H5/1Kc9oohE
vmRNTEYfPmmwibFBwuEz/0bkp2BpC6uA47DVBBN87n3LvtuA2/fAc2EQ5ZM7USOC
yxTa/56Zqpm7FU7seDDM5wD7w2if4RaA6Lfh+H/oZptPYxP0X3k6X7819NWz4Mbo
K5DI8CdTRETDmojM0yt7m70jV55yjPlTUWKPGpMV1UKuV6ClTl3ObrxahOjeikee
aJRM0ihDXeWKK5OmNs/lDu10K1wK/AhIS85faBDxlzLhHDUxPbJyd4hz8FbTvLTw
hz/IFC7+CdOC+fK0ZP+WDA25jE009jf3DcMYnrIqm6VikE3jXybiBbT0vFGVn9AW
u/AwqcE/49w1Z9h11pKiCSW0EhclRTl0th3WKjlM81Wk8q+zfXmwG4KYYVopttYC
bOx92yHaO6HKkwm9jsQ3dt76r2mt2Zqj15F8IQfrtqt1wFzhcTu/FC4zXDVdA5Kt
E9vo/vlRjEGCRLqjM+mZmQkbf1xr5ajMXJoTauOr+nO8cHoE0OJMYDWdrFBBHZTN
eM4CnHS68NXHX9M+iTQGDdGCzJ/uIHgJgrW/DRsepVLYfB4wDMMrmshFzRpAwPfT
ddpRWbIu6PPeucO1UCJbsRp38jpdd33PQU7BEQnJueGvr4U8cAM6pIvxJexlZYx0
YaWT14mf0E/XAgSvAGccre6Wn68k6h8El/PIk26qSKaXGuQLQh619HEGXy3WIURp
vQsXVnDU7ehgwC/GzyDZdBzmL5gddopS9+JUY6duE1iYU5/Syt4cwsAD3XDg4RqK
zvUDZ8P3nLoQ1sHl99ojZg==
`protect END_PROTECTED
