`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pKJuqQy8H1wdIFAw5U9StvLfhf3eBxeOAqbnbmCLirQN4UZuHcM+RpqWtMsdNNfa
LX23E/5SYcRKeApo4maICE+Af5agRixEJlANSn7cWXVeeCBwBczi5SbcC0FUjYvl
0VXPGOEgIFQ5/hG5xvVMb9c+2m+pgWV2BTDT5sIzzZ/2vz0jPg9mSEQf/+uil/qO
8pjJOnx2g4NlRVZrhQQQnaeHI1dVy3ghR8KQQemDYJle5ldGQmnjNkWecaQcrTdE
FxHumWjGPwx6V/5xkcZ81r7gde6zTyCh/+C3H2DuLbrx7KiuxY1wjeciiUfJLSCF
7waHpdPuCOWdyFk6ja91gYY1lmuJdLuYHpfRqGINv/EoAR9viIgtim/Dscm9NOAP
S8psll96Nb4CS1xte/ZDVnl6sKS9JDMMBh9kK+vSyxGMwSHWEKNr9rOb0TVYD/Iq
jluwlUFqHcaZKDVy3cyEOPhv+GViUiJWjDHRKH7Dk5DXBsXnbe7SLE6LwmTuch7o
GHm049BoUQVuH/h1tmk7zFYiNljwPOwOOuqbzcd9PeYhieKPEWkd2g8FvXTjV+mf
UmzkBcPVx/TP23xtjGFXe33/kivRSVKiE/mp07+nso3qPI5qwuI6Qty8wosDj/QV
3qFFWIGXhGk1veLI+nzOtBoDngXANt1BchgqPyJyFHWlKOLg+p7P2NEtaQqgORgr
rWWGsrKAWhODwIhRwri1Rz8hWRwnO8EddKrQdvQztT7umZAPa0cu2S+oXp72xTkd
Q0Bjj3Nj57FlcJga4IajX6/DhI824kJtAshxREUkUHeE1st1wdS/7CNc0wg2S2oo
T/pgSaNV1B3eNkar6LXeEbnn14nh0qEV4EYwgfBMWDLDEq0XnSZIroWBsELEo/vR
0DLGXDAuXLql8BoTHSquDzkgRLCpB+f5PUQQwHwsFdnN+tm4c+cAMop6W1JZTfEM
l7lTHaLNKBpx1bC7Bk6/X6V31HHBHXVVGCaO9sb8z1y/MhWN9ekW1KeMN3DhXiUu
`protect END_PROTECTED
