`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oIOiccho/2eYTjEUUuB4l9f/ukPi3QV8ySHfNIR/B7qxM3GkA6yDZkp5XelGniF0
EYaoR0al9SXNHQv9pI9sLU0Su/1mZHv8S8QHaTh0zumWInK6ier2ZmsPhiuWF3Eb
dXABydMZZhGhS6e3COmpuw2bNNnP1qEn5kpKhXHQDXbH5lAi14y2LuqJ6a+PpwRw
FXsnEl63XZB9sSfmD2HFR37iZ9/wkgNpXnDRtGmYi6rRvqbNZ0bt0F+YL8UEtnux
HDIxbxN7X3MkYpIxAqKCVTqRaoyEV/eCFCqh7CpaUIloljQzu/Y2LKS5GLHBuev2
3G6bTm01Tn/JL/AKNFLoknspXRx0hATduqyWVIVORlUJgm4QkmjhcU4gDRY3P5g4
y9Vw2HquOPJAbT+k2X36+18KLheV2uc4o3pSoTjZo+DzRjXi+CYnyy8tmKiWzirA
D0/C9fFMEHy48AdyDbcMC7+MKOB2L6DYGpVMD/VPF4kiN98TvNphO/SViWIUa85S
sDwjEvDkdsiCDCslPfmEJrJQiSEYLGp4gChfm68f0qK/z4oAOjOgoJkQY43UlLKd
OLB9lCpVC9IpVDITtnu00t8SdcHOFxmCf8ddVBGEsQ3GcHqWJSYOtOR2mRv6ggtO
Bvz6Ox2HisfXWiixpXdRHSVli7v/PW0h+OYI8m77dxR2YY2Vi3UdfTyPzugaxjpx
FHLv7WjBMOYw098D2Sbt3+uKZy/kKFcnYIwsgzryf0hhE6sHh4M9EfLIlv1sQqXj
EJfQepHy1hkaZSLHJoVswcPGdo+N7hz7QO9Lkz6qmDDtWeXDMivSq+033ACeiMHa
a5xzsNmMPhjETe/9llWf8Exf0Kl3MjpAd566uHWylAPRXHxUEQh3IJUe4Y9HF5qj
zs+lxdoA0ydRzormz7BhlbT3HlYNSQFtupyxzJHT1c2KPXy5CnCHTL+m60cOkfGA
CXGZGS8C037lg328opMKK85Qf2p1ZPhW7HuJvIjFePX8AQsCKBtLd2Vf8USZyDWR
sVfNBqcBpT5i4hoUhts9gknPmMX5pPEBHGiV/z8oCmeL9rZX9PpE1IeA8oh0e0Cl
uMUxxKAHfU0gjl2+fJuJ5UO9yHVYdBBkAqWqUjDV3Q7ZyTRq+iKIav7BSYcOOEZq
cVVfeuVtRTrSbqYpRsrdkCREsC32b6sjzXRGW6GACYs9khUvkYR4g+yWKsZiUwu2
oqcTGY5sEzU+thidE+/KsyMyVabgoyNp1Vi8fT58VSo0Rj/92iiqxiswX2f/W6rr
yoCek/z4jVjPXjqar/jAGu/Uz/XP/6dkFcFr1faYNPI36u22H9OrYJNTJWpaAiaB
yEnNpJdrTT1fuHqQnq65cQ==
`protect END_PROTECTED
