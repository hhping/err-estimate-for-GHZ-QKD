`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D8GFqRfs5ujs56HXXyUad8gvUN6X4qtryENq67c9blP0fQlVP7rk8mNXo6i2mfGi
/phWzhxScIpLuGJ6ypdyhuqj0FWXfVmf8jY/QlUUgEno8YsPdH3tYpLCUiqQi7Vn
ZkVUMC2WpdfVbG+kHmZ/q6+7Daq/MKz4imfoXYpbYu54C3vvy30F9VjkwTl5QAaG
XIYQ0UQQkllGse3TqAMHizx8wHopRROJgp25mLgO7RpbhRWhVaOQZ0bheP0yLcil
1kZpatJ51OBDhczvKhI2OK7l5V0JG69GpXaZhKgn1iySz0EOzP4ELPQyCOvTdcU6
UWooK2vb6QWGXEPURX20jlFEGhhDxHJUD7idtrJ8KJV68vb//JJ8AJ547pko1oAk
zvJOSzqh3xQRz/k2n37A0HCVZu3B+B8E35tZ4kEBpYHXuaYnJ8BICaR19uWyzcQr
CE+J7d8eySolPF7gS8rHqw==
`protect END_PROTECTED
