`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0R9aRdC7PRM/vqZj+91dTt7Zdjpgmaf18xPBeu33ydLSJKnft9xlagE3q8HrmN1s
AOnXZ5Lm+kU/aiSRD2pg4DAqKmhusOVfTKRn4W/Po2IadfsIg6G5HpNxTq6NsG/P
VgUJDlZ2wCm+eTl89Qknt6UtDFu2iTyRFr8CuhLtMXlb3nYDqZ2ux7/MhCz64LoB
QzF2z09VQAw5tiyoId2Yrra8yD7O9HD0I5oTwOiaf/kg2CMydjZjd+7uDdW78gSu
72sFsfTokKrLEaHpO73XIRwLAtHDbO9cM44EF926NFsFhF8c1jSZEsRwaH5QDVZo
pViQVJ/miDHssabXsCOfWg+qte4weegXJxFWWeg2A0+Vvpm07X6GxxegvIvlHUl/
/Wia4voBdUeqnJJj2jRw2JPfwKWyDLNOXYA2LqYrf53BLTUxWjzjMWXmTnK9L+Iz
W6huZiLGxVjeyCOaZZt+lDU7qaKNw8+CFZQ+gkeTi2+TSqk4Fx+oBT9IXHu+ifuc
vsP1E2lARYuUqDXyWXYZlqcuu5uAz5wSUITUINCIUr7+sL+OUgRp8OSHJYKCKPLJ
DpgzvkuaCypzjpcDERwmdpwxKy/16D6d/hzgucWfcDO434IOoZlOP8wNqmN0ybM7
znAhfGvUkOL2u0GfVcpRBMHFnxejKvd2T2L837Eqy+Su+eowY6M+3ZjJxcFK6SX3
xYhvFy462ziNlYkJwTp2HOdQyTD0iL4sm/1WlAUeJwzmt8xEJ5wvT7SvAVhchqL3
vwe8b6dif8HIdX9g718HC9N86i++L2sfMkHoIzk/bDD43HXhhH+N0S7PMMnpLao5
PUYUUbhNQfhTTHjHVph9A+Gmr1aUac12yhHvVZKpaByChlu3sVzQcSQGEjsADjBy
Td3QaYS/IkI4i+037T3l44eTDHu+fhzu3p6omSTlbR7iIKFE8vzatenXOByLlMTb
InZMA44D2jTFeg/iWr2/6owZ+8wK7DLNWcoDXSa0LXON3kNPT4mRomQn2gceezPU
VRl/lYIT+y5zKB66bDVr7OQU1EKIuznADQoo/n/WLZzlbIXY6kVGc1oYFQ1Cxsww
pRAqbunYzb9pbQk2iV8TconQPiNJuP8YrbpqolIFwq/oKfu7IwejBP7wzmclfM/f
Bq3f8DY5CH5DG2xRfmR+CGbNv4YQ5lwHi5s+YZsiIlioMg8i02210ZUYlKx8a83O
WKg896gxYXGzSkNdP5rph2WwiCK3x6FCH3EmkbHJTEDojzYhzwsKz7BNftnpC6cT
TNW6i7DUDRgJKBuXdftC60FVTQYRhbQAg6WAeLuFd/nZarTnrwVQRWEGmWCGUG8G
BpDJhimbQUAat/uVShE92O/2sYnKBFAg7yl8eoSJiGnTxqmTkcUNbM4c2bdLyodB
/gaxXGndZm5IjEXdWzw8LGIABIu72SaCVBl8ozAMwWe3CJaCTfzqAnAjri2Ab6ug
lvZOIrv4j+FZBRX0wqyXEydChj5fpNYfpWkey1eChCZjv+7xKLeEUYZ5MtQeNPGm
q54hMxmM3rZs4mFVB3HX7ZQwtoZCThGWf4FoNRkKa5FeNehQ2Bq6bJvvrrbzT1Py
FQkbKloZB9X4ox3+/67phNEKiHwkNOhXNRGWnJiO1+PF5wskgTcb7VtARyiymHPH
SC8l+kfwe6zMqBTwRdg1xVZNKrXuUTwHpXUOkILzY90=
`protect END_PROTECTED
