`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJWpPzDobAYCey4y3w7hVLhY2ts0O1f4zlIbeMEbM/fiVTuCFoWNtKWnB7RfyRi4
mkNO5IvulvmGbkshW+ek6g1s7I6I3EmiDJBS/VhpLGrqUyYJoTtL8VcgMfBvT4rr
7oG+lHwbNIlmnxnjmxFcw4KvrM6rTBBCFYJweh3WP2yQFXDmQOrZxuRRQ9Ctowp5
ETDkuqZ2eGZQSgtSo73zGVK6E73uHB/2YkOKJfgIahFKbK3SDKePRj+c7i+MhBEu
94CjmAMaVIFMf/ynYFAlSauO/hsUWtvcvSXmtyUmyFiqj93ulH7VTm8tnEWazcJD
9uJxTLOmLSv6DUU5hh4LpE0qia5NyNUjvAMVYsmrL3Lk/gICSPY9WxByTpIf4TDo
5fsS9HShMP/5pBsdffmJumQL9AZfEcNehflXe1JDNrrP317t8oTGNIaBWJiAvUfM
TT5qQbCfoyTYKU2LZWy4nhMNHqcp85NruHho5M4nPhalhd/kFZHUgK3eASMe2FX0
v9RTiym6gxF9K+zjctnUZphiPAkZNsmbn/ygxg4v1hIFH9dBZU3MhwrZz19bBPe0
/cLJMZqNZ0JD2S5v/mSpWlSoE9NSoeZYJLSTfwv/kPh7PxYvftqOLvGRJ/HxHCxk
AmD/8dBNXrSgK6jjOPHTr4q8ZUZ0lOSp9+bbM5ub4yZHVdf9zJB6KZfg48Pe/Eck
qYOmKPduZWo0raSlScjHPS+HsdCbZ3jGR3bByljB2xUywMkAvsDNS3L6JUgxdcvT
PGV+gt0P8IGKN4A1gzeeljoMCqXnX7q3wvqU1vnA5cb6hQu9QTegN25eQol4ipmn
TGv7MW0ug/dL8Q3Rl9odpyT6Un3FLuzmcyFwnDXi7SpT01AvFQPl12cJNY6iXlFV
0xe+1kuP1IbcgZVeVhK6sIwoPeeF43+652wPF/qHVZSKFv7dT5ta1vP0Hajj/0EZ
SyLslFZT3RQJ+vtjh04NpKBdlNrEi4kC9WIw2aK5v0eezCcXUDvDGru3Pg1h5yzQ
3gVewE4gweOFkyjmY8g1OTN+GjxX3h+P8YykPD4zMZonQ550aL9odVW0WyArP7LD
fLRWnvecPLNSdIKTRRKCMUzNKYDgGznmmqxhqXEObPUbajYRK8NI7dmqxf4lNtN/
LJnM+ZdxtkgQ/rmDAvWQOqCL9eQr2Q5TVxiibaNU3ighGeUBehvy9GmFtxn/P++6
9Nb3/uEEe1G+JN+oKcfETj6RgoDvX26Zs75Tp1wOy6UVlf92OWo87b0IVy8f20u/
JycZULBYnTmtyFw3XdHT0PIlHlOPqy/usg0myiw/SPKz/oumBb5r7qnGA/LmcoNJ
DvbTLa7Z4nvCnG3dzvj/ipgSrzWVCPe97NLgd/9oI9qy+8oLujBJUWvSqiprIQAP
o6PXzop8Hk5Z8qbKsW2qdQtEYAfEzsZVAqD+dfKOHI6gSiSQqZnLUXbve6prEqla
KSz8v/RLz2pnAW5AHHVhGcW2gjn69wJoNaw2xX1cleBbmFMc15OA4smhzfYVAI5o
rOUGHqlXkDuEZlXSF8IK1lBEwEx6BIH4+z1xDxv5i1qKvpuzCHB4rPnTCzYh6nE8
3V7OnGTSqdD1cqi+9xT4Qd/4AAvg1rUyV8gD4/ONhcso2yrFAUfKvN9nkVozU6et
4R8nNX9UJdYYmbhDP0w/WlpV3IsrRmqv/tsbb7dhSIoGS50/tz++nv3aGA5MulIh
l+cJOAdbyrXPyCV1aVvh72bSXVLySVtAmoxTt4Cb+1PrGFLvWg+iVABCNMYywKVX
0do4LIjk7i7GK/rM0prHu9dW92esg51/ZVU8TxbVvtqbOkYygO+sdWWJiRlXyQL3
QTYpCkSdKmfkzBXr1EASGwbhwSIVETTrNUH+HnpPDg7aXy0G9b2IItsZdKIoS+rP
e6P64X1dzkriHYPGc5nlPnvl8KTleG08/YafVAB+9jhZuwtyb85ajqPEugNtxeGV
OQEoaMwi8F0cUPcTBXKSrKnjINcbcvrTiek+75l7UT/PggAz2hsV1n6BQZOmhlOE
FaAn7lPVRGf1YwZZjgad4FfdcFaF3E8lmjyc0emyLNXWvy41SaCaPSd8wIkcSrNP
8mtrLxNscb5nbAb5FQGYJ+2w/sDPtHSldZ8Dk/9UKv9Um+5IZTtGeLnq4+fiBvOf
XrDMqSe1v8gAV4Dg7Mkgg7Oh0och1YTSuJOHdW8jV2ymoDc7C6JhZsE6u3nGOABd
hlDDRcadfFO8Daomcew8y5AQ57O/Axmn5J6r91nGy+TOQgSVb1XNDKvkOxie0PmS
2ugO2JT7MvEMrwtOJ4i/qCWgqr3gNtSiHRXIyBgPkQ8TDDGxWrYoNP652+t2b5Zi
HNiYIUhFiltN6GRsZzufO1lLqyqyyuSxi5jeZhD7/3ZVlvzrGRQYcCs0yOdLQbjs
vU+GU7VSvG847rfbRkRXf+FkKwfLLhrLA3fDeMChSqcFSbv7KAhJPpDlb6ujbn+2
SN2B96X0Mmp7NzBvLxwVUAXY6ixy23Yeadnh4qI+oOtCzNeMZOTFcfacXnxJ2psN
4Sd50okrd2udluM5EhLml/n8toOFBwpI60b42ix5ewboexiN5BTVskh6WfkKGcru
OvZWQiNEHOMeKxc1YjhAlXaPPz0gh3l5tnf9GlRJvua+mwnoSNkRCI8YVu+UwPFJ
kPwmcBmZFhR3znVAf5sN9PRBJlGq7z8TldbUp/mlm4+raG6WjRxSadzq2GsK62/S
zGI4pTkmAguJW+1f/Aho4PGCbpZ4JinFUWb5XlNJsGsFiYaMy7GKf4SiosDVf1Zd
8LqnuDHstLLq4jqAppvuUda8tGkMgIiad4XPpCPxW5/4UAJ88o7GDqD+w2B1qCWr
/NPLwbeOXhZDecXKoBi/vLZndWIA19gTBeUW8RJGy3fjG+Ey0xJrUnqaC9mpp+s0
2tOkF8/ViHmRNzOM7FMK8WaXy6Gqsxp0JHLsg1jpGOphgmTHdrC/+2M/tbQx22iL
1uQUw4IXvfFuWcJ7c3q8tGAK2khY5xYE1g/C9tOfH46YeQuKN6MRDOcVnTlPdZCD
hQ+X4z0C+BWYr5UIxme95QDeZ60TOsWt6cPY0Se2IqFltZllf+LhjxR2pv2VF2WV
5SYxNVNoCrCDmUepawRV+lrQP1+wJDRtybWuA6J6VE8sQLxworrFuFo+9tY6QtRE
o/0AygtICZ33GpSD1e28VjBy0DkOftwLw/UKn541LGrynT+zfPQK2Ry3XmFKDEfy
a0xyjzaDniLwF1sjnhdwWnqBfF1HFA0VIj80adPv5WHUjSFzwIaZCoH+yJVz7pxu
9iZPmMgBWtZKoOBSQJoEg7h9YzxsjJOvuGB5OY5v8L9R/nQ9/RAoQCaUKp8kJgwe
MQPHZ7h5gDBHVbJXGA72KXFlbZBIX9FsK023eMbd33mry96lLuH9ct5CgCow73iK
yFUdwM25Jo+UhakhN6hQmVR+0u99GaF1Ka2jfWxOAft3FbUf4HbA4A0Wl5SjkcKQ
cydaB9tzxuj/g84+tsk/MeCKGiEb7oLzHJ/WGRlyEkjvq8+dpTyIcLY4E5pnW+2+
PHiVdYoa7UXCzSDcfLxoXeyaQ0TgRGdZkJfvd6ZPpVSoYeQ5T9zIlnFyaNfrXasu
D4j1kXU1nWK70+oCymrjUd5edga+DYOxW8reN65vckuLklcKkKU1kOOBh1YmxLKr
dZVohPvNMiuxDop6+kxFFYtKTQ7qGjhJYFeZeggfYAQiNxHJRd9CcLY45bZn+AI8
cSGXM4XFKasdlvEHB9yqTKpooTMyVV+fwR6Qex51Yu2LtPYASfb7+WgZllMCjZDX
QK/SkP34Ny0XZgzERcMOc03bzzHzXzDNHh8vvz0Kh974M1wwm+Ztj5sI4rJN8bVO
sI0wTg3FU+CKjBsFV1RNqf+vRBDYj/nnZGfh9sc/DOc22BYjZv4NXJie9J8omlt2
G96I/+37awsdqIBwtbV93YpYNCw+KD9DkfwEXDxAtsxjq/x+RW5aMMq64gCYv1i3
3AaqL37Uuv5YJTSo51LieRbShbEn3qqQQ2AaQt/YhlJBH5kmXS8GBfjhn07zXWWz
3z5cM3dam4fNuJqwRR9Q2GFk4E/f7PWrLsH9Wt3Y67gRQKT3D1KJ0TazhY1hOWeX
TBB9BN0zEni6x6wAISnbOtBVa6ZiVj+ueO/SKsdIuvfo7/ARnWaJdvDElsRDukKI
bVyIPX4ubOiicvDt5FLm70HbnSI3Ehf3PQigpMzz3p03+eCRq0yHKaS3IMJnLqVj
Z0C8bnRupZV5+vFGh80PxmjNGQWwSvrl056GQr1Z/3Djr6hjbXRmXj1BYZFGDaUG
8qef0ZzKP0Kb+LIBEhfvqxJbSVjBOtWcTZbkq15Y0mk1791+9+S8ludyVU5z7ywv
0v5k3BzDgvVUYiCeRiLNioXE6JmWzejBR3nH4V0Bm5rCSpGmphCXUvRB/Vj97NXO
g/lYKJpOTkiN7m/n0su7gZ+Blb3NFVEfp1lLynldwycnjOE3I8XRFXhKLk5lnxJG
1LngD/gF+kfRydyAR9Hi90c+HSm471fjyYtFJIw7s51nrD9F7NxbmR9WqKJB3BXb
jOM1RJQiZOQlwB+26tu+cmEIIBMfHv/ZE8NqrwP3pPJrKgDgXuNqcoZPVujvSVxw
KjdnAQBeO9OxOYizB84qrtnqI+FDzhJfRETbRL1JhRJJV3aRjHRinjvqi8n7rT+u
w8R3b/RJUTvV2r9SYmIG6vpkBqB0NO0f6CqqBcFPhXfmJ11UuWVbor+w91Ku6oVm
3A/rTm8VvRm+RBXv9Ec+pVYjKga4Xjr1UMAkmI/Kt0Uow0ttul9Wqb4L45ymRgz3
4QWoXWm1iHHg3o451PHqybv4M489JpRF8mUlmoXSKkOnFy+E7fzjkyZYyqEE9Yzz
2lTejSnVJuvUezZrrENbD1NPDXl6P5pXwZ14t1rg1JNw916rAw9AI4GgygssbZXj
jLATTv9D1kJ67E2R0sTZA7ZJINpo3S8GtgjwbYr/TR/EpCOlFPgbh+Ba9Y0CYjCt
xAcO2u4dciTcXGBPDkYSrXkDhPjXqBWy4wAYP9w5KqonMMc6vn8EJThqWEvh1oxF
yiltDsC7gdiMM4jVWwtCwvXsKezPR0qKgfexJxRM+E7fDQxCcXERNQaUPq1N5OZN
HzveVbocwvP6o2h3WeVD2mu4VB0Esyq7OTf+Y+JX7uNbqFxiZFkLjNRT2Dfvkklk
bU6TaSJCT6N6ytR7SUJA3CD5RgnR8FaMpuSrxrlDb+/6DQR6l7k8qZsGk5PNLhp7
C1U6cf/Oza0XMKvHmqkAx+i4WZ5FfmidcrRrgA05R5IeK2xLvfDzFTN43klyXC41
UF8Z0YqVJMrmxP2RRvrOv/aqwo6Jlew26lrXINnJjIIqdIUB0Trs5/W/ggdhSlFe
BVyv/alATKjO6W1UALnC3M2y5EejL3Z8hMudlUoHFDgRaePue28AfpE+IFAvygCJ
CP4RT4DkC8zLXWydwxmT5dVInlp4afN75IjWLT3sOiK1RjId7qoG2C7zOeoS/cQI
WN2zheBHtoShyQf60W+w9KHO9hnc02UYqdb4YyZJkmRxL9LWvIxIJJdk/qLiF1Py
DQUmGIkn6CtZe/boKQmGWP4aHxSdYxfTz4F0dVr2XUN/rvHFydjfU8/pnbZj+is+
a7z29vcwtAG8Z1CRDvEphEWjeL8joc51+rrH1ox2qp1VAjjJFc6V/WyUhbtmIUiw
YuR9YWbPv6Hzui+XR6DCypP8gIUUdO7OMY05JN+adFp+a470DecA77hCyTPNpzY6
+xfqVm3ejyn7bK5/vCD+wcZ9nmN8Izqo+LjJyxKzF1H85Vvnhz7nzUDRFupXnJuZ
P9u/1DPEpj3G7vpxZkzaWJw48Dmna2OHHrcF/POeu2NZD2ZZLf/B7yHIVg7PMIJ9
UubYusgNmJWYHmO+67otngQa5VC8WrVj48s7FOY2VeAgmKbwXuopo9YChInO1j9F
F4FjhXevMsOMESXo9a8A7ajIzKBnyxJEvPfmD0hBk2s6yf1/QAkSkiE+549RFbuz
opgbGNobD4SZHtXLpDTZb80FhZxUSu4SlA/RZmkvJWdpfg8aVzJubIDfQ+9yKbDN
zsg+BQlg9G/cQOIA1VUSy1ULaNqPK9dWew+XA5QhMrtNlsV3TPf/Rz5g4hGuHWXa
lvgVGVP2OUOdRM+DrZJFj9hKTx8LsTQl7RvjtgqUlSvGk4z8jHNzw0JB2j4t9ymJ
xN90C80SXjouIRoNvQUXngKu5/JognKSmYBML6gkp695tyw/+o0fbEQa39/Invlv
cyurrbQ7hRkfZzbGXFL/Tl8C8utKUttNe4MAV/CZEhAQxQCVkotYaGjqxkPeAXPe
8jfeXK7IjogYNu9sRzvvWxKnWy1BZyVdrIZuSpAWY8PkMdzMXlF7aIO0yV4rhzZ/
O9vDMRu2rrIZ98jonLPxb0lVbPguQPKMWZxVzeFeyD/8XW9nyybplv0IyzQk37PN
8zPnP1S+Qcx2dv1Ph7bbf6FfL6+VNnF4sgcr7ZGL2QTZuxK+sPbgB7wdWnfAkCJ+
YfgXuUK9QvyKH8lEr4RM9E37YPh3Z6brOK4FefJki4z+bd7e7gOn43VHPpEKEzIh
gwzwaZlDvrlvVYnwmTmDF9WjVHcn5RECXQ2yo3Cpa9oNzF3Eo9E7wNIPb02Njzgz
zHZdpq0hPpx7mklCmdt8MXOQjA6Zcg57rJ3pof4RU/9jMeJGsrdeGX7WW48GITOP
nx8OLB0ASJRD+grLm/A19mPBYMdkJat9AQsHg6/mnHvfEJHBn1ExXrUoR066on+p
82uGoTIXboRuPx1ezX5DXQHA2OYK1mH9cWJ47f0UsatJs3B9naB7Rz+hgXuOQjgq
0ubYgof9Rssv8CmB82xnb4oEi4PK75ttVjhUd+Nc/PBA79i5qNK2abbOh4kicyJ0
+8o6Ps6mfKtT5BZMqQzHddzeVuUpZx5HEiWiCgFuS30ENOavexBUvnBcz9fDP0lE
NsHVM3f3H2Qek940o5M5mHChK+ac3WpRJbRTbJt5SFVfdk/esNxJWupcFupdZF4X
868TsNtHbGRHw0iex2qbaLBnvJcApYn3MrVsnUrR48kb15DMuDjjJWKti38UTRUc
W0I6r1/5O2NdiW06MwW7dJHFuru7DJOD9nzhf1XXeKfZ27o6XP/fIpZLRAnN+pXn
LMw3FyOcrJBuxyAfYIoEHli9sFdsvUrM91s6UeDSUJvOrfogce1vg3OCjGTrW1h4
4kg5/N8WTnLFEs7l6yHSywrfjYp04kqhQeJ5kx2m+SKOEkk0ldo2e2PDqplLTxMx
kyFOwgzBRWJn0SqHveyhaYYjOEdT13GGfKL1p6ecK1vAyG5+Zap89LbGkhV/3gyM
HNlU05upaXpIns4RuncY7wcp6cIFqVpNZiMmqiRr3x5VYUinrY1STDmspGBszA2h
NiA9k7Mwbl9MhrTWHxIybl4kZarMDl+GAC1S7//InKPnM1SSUgdAY3JD9mVBH42D
90YQiV01sr2nqWuvjUwFwZan00cXbnl/J94P57XPMwMG4XuBIDufsMPvuJpfIh47
ghlXExdd6iHUdvbJdQcx6Y/6TT6+LI7wlkMaMp80CLyMhMGiYVovsbhwn54CIGHi
E269S/T/XRAs8ODHNRBYSiuyI+WL2DWn9bEz6DeTBgJt26Jx1WcsuLEyKUCFiwaV
KSg9w1d7V0qLg9Ft4ZRHUpJYjgimdGkDDGHdWv/bWaFQcHUrj9ZErINzZ/mp1pn/
dYoU1O6kZ0cex88YTTlBfH2TZojDaOozikFVJnGOXz2LHAtOlMvWMtpqA67tAp2C
PNhx5Rh5LdlzQvOKGY4HQ6Gp7U2/KvBGkSoxhh9oDbuIQSQ5VfPg1C4Lqo2LDy34
vcdijKdI1nhlFRiWagmBYWbkxlS9JCclHftL1n0FSy9ZDyMmUsrMS+DJvW0yR7EP
lNghc8gflwANu3Mx2kaLJM45BmOyYNg/IluNWHCusYQoUHs8FS2NrKgavgsAMnhK
p8eTENiIRAJHiO9rcvXS+rcTMhYqIap4Yg0pOr03EUzSXtIeAUvlwoDZAXyvOo2F
t2wqjtN8j6kcvQ+i9kRyVleNHS6N2TdxqYfD7Xks8A55G8LJK1+COgxnAhpByBRb
V0XYPyQh2f7T42CXAgbHKCAQCKCcwlDNnct8hiRWvEJ5BioIkFO5ZDYc75AtjO+G
wZ4SEDDI71KT5PQiBQf4pvotN9xFUJ/ZQk6i5aDVW0ea8jzGCXG4Y3B37Zjn4NdP
WxDJ41sl9fY+wpdBp705sMwon8iiBGXS6Sx2GuytVZ4xI51ywUFfXaixRbjq+F0H
wE4RHmuOAi9s8JAXf1651he+cyy+nRekbQmPRa3hiCCBl3WYLSE1MNjzpuAnsCYT
ftVFeu/V5h/r8wEOd88fbfuiHAegUJSqYenfVN58mPRC71ogunbFSe6phDZzRZE3
2WARtNa3AG/6GzB8VIb7C6mvW39ld4OQ02FZzJHgN73c3QCJwPRXIXAHxkx/tzeO
p39ofqn188YIFRaN9qzlrgtBcBRvSnHkLC17HFQB043GRJ8IpoAWASXLwP6eB8Ir
1uBRYMfbNNE2F25cd3eT7bMS85OgMCf/w8fVu4FcGtM8tc7/n+M7U6waWiBu2G3R
146+24Wl5rPXcVAO/+SOWb34LwKtL1UN3Uy7j+XC/EcD0bGtfkGT3m2VDAp16jpm
JExuKGgUOg7fvQsM+tgccnZ/XlxqNIDjo7T1b/V9+tdeW5+7VvpYZz5hjqWdIrjQ
lAIHyCiCEi8ogW0XLlznixiMqFHdez4bt2Cq/lGExCTVBMm0sxG8XTiRh20X19EO
NrPDEtKo5JuTj5W1/deBXFTcF3kj2cjWeA6X6lj5qbuJvfKPscBmq0uATkJxgy/3
cCvN6+jWQtEPkLvXKZKwFyx0Wazr29Pwpycb5r/YvQ889EOT7OCUxig7LBYph9jO
rOIg5d7CsZO/xHigf5hHDU5QQbrv1o4YL9+LS8v+DPewdM+fVNDweC4PZAuKHYfc
9hSeAyLTA4UsvCmfjv0wwooElG6+IO3CROGc5mv0cHfRE/UKBHH+DS8bxqgg3PLl
WMGrYTWQoBLTLm73Ys6KA748VfM2sFlJUL/HMtOmJx4W1dCMFeYMyD5X0DJsE3HJ
d0r+9z3pj2/RhlypRwrjfcYVR5EsNq+QY+Vr/0lT7CRL5N1KVMtjapdkTJTC1x8R
aYk/5KIhx7r1Fuc2vGSsKdEFq1xR2o6WMQkk/ZLzNK+LhiDOS6E2W+SVtd6hBz/X
vy7HMJta5ZJw2v7vN9XKeG846FPPjMLnSpk5Yj8uGufJL+2N/ESwEeSuyT8HYe4K
Ga0wf7cQNXBULWBazM5YBQWAeltvB4p53TGK1a/Hdh1L3ebLOebHBnDP4P1SLvEd
CR2wp85AsfnuCwtrPIpglDJw2eNGqkGa85Xuea9piu53zigSg8y3+ZBX6sR604aE
v7ajC8SgwKLuErzboFz4T7a5ZWyijOSOgtZXDWy/NV6SdumblfP7T2zAXlwRGi3P
M/SG/LWv2mchT8RCjkSjJGhEcQ9l5oAr+wfMmEKnr4SaZ6P2g9RllnCz3IUr75F5
TaxjBlCwbKzsT8ay8moFk9vCfDtJPzySu/YaXOgsN1pLQ2lLSIMDOoL89nBde1jV
eSTwgKpzNjp8T4pce9JFG4rCcLfZJPt9WSWu2bz9VI7LJe7mFGI+GqWPZkQcf54d
AR2fNuy4WECbmfHv+JXgWoUSVjsdzW3Z8NHeSzAj+IWwwrceJtdWg4nYlLYVMCQo
bG7mB5GfE39wpLySIh2ZZbdstSsbK0cqHcKSv5QA39AYlK4s2DYOoCKuCbL3w5VN
MEpYZxePyjpWAjIN1mcxPWjyqqcJQBVHBlggjzLI0mypb6CnoLYbKo7XxKK0XIcv
SpmNUpkgOuo7bBv61/burBkdM/FcWYHU8abYhVUxvCpmTbW4WK/ZSUX0rJYvreeT
uI/pR3vj2nIjMjnTTAYWm2q0OxcIm97f/2CIHFxneG8lMlZQMpF1cdvG2a7DLneH
bprSsKFH1iVFOLK2YlFtS1Jn7+C4FfS3aelWT0KKNxAtiG92npBvfx8P5DoSvScu
nWL35XLckHZzmXF+sTAq5SmdzAYp5Yq6EEhJISTFtFwE6V/iG5SSwRrjMsf7oxhE
g8ZfUWTEoKOM0KgZzsLzqylNygmtd4rvyArn0x8yUe40SjmUe5b7v8sG9PlQyv9X
hnrtzR/ZXQS+9znSYGTaRrMjdNQ4owmaWUtMWR5Jkz8zHsrQVzUeSmE4fiiA0OAj
Rvo7x0xBJ2/xgGdejke2benYEC9zhGixIJNhHLRYuUZQ9e2NZja6PCDf0WnRyUOh
FkSO8id+LvtVvMzo5MGjZB25NsREO3X5gtKhFVK2xgXpPkwhFdaFrvKUDDfN2nSq
fP98ubOP1HlHGK4fgf7VQEXa8cdWpuksZKh3FyMT/jQ6ma37HoLh2jgiL809nPZB
ggm9z/GHwLdv0UicPKlMf9rX0TPZmaJaYABLZ64zEHBfIbf+wp68ddBE6Lc7nXE2
Fetd12OTi/TL5/IMiwLNyKa8L3RNboGgbkSuOqc+/6BwMD0S4Gvn09LoAyO2p929
2pI57mX7RyblYlDEzciBhSb6bWo+PWYl/RSsgjXKsBm5mdXrrjRhsbo5NcmCmVnY
UfZvSIy8NFHK8OtGq9Sv6WClU43ilgRezndX1Gi4369An7+Q5F5apMB7en0J9IBw
ym46gJNpGv3PMSdnJ3i+OpHaHlRUQYVnGdIZLCoy/Tp87glkCP0slGzDg//Puodg
jCKT2raroh6NZixtjDi36qDzFSuJIk6Eg+P1PUYHfwQ0649yKYNpZoRutauB4t5u
uREtH7v8HvCzr1UF/ph2ZoLMjxVuiqlEXLSZ5Za3JD1+JlZr0C0DZcep/Edi/w5E
aqCSi38UqhMjLFvvUjwjQCs5YOJLZ0194aNAsH3tDVAoEpAPGauN+CpVOw3SHzlq
6ljVe06UbUFpaS2OwuBCuZX/Qez5G5dpxyGbS0sxMeHt30ew4QQX9MufXxIr81/5
bijj0Etz6Ml+/O5OJYGGuavQY68PeGjAhWbkUsFLpmWKmW+DXs+qgMguXkR8cN5/
Q/HdpjlXeCIb2Le+GdncyN7R83MuqB/x3MkZcQ7hy0zs57A3w2TrGX9YAHAQo1yf
64ieNGngpmCIm6JfLfmy1pu55r2FPGyACU9TzaLX9itzx40feEUsSBCdwUvjTZgM
DWSl4ZAhRx6dVwqwe05NEb/i5tgHfZRhfU/n9OWPx9I0jCy6l1RpHLjpfThUNgPE
Av/1S1Baj1rBaeevl44l7vDOiZi+Ym6k4C71vUKDPQQs4fvdsEQ+H8tIEZvNVEih
Ev2mC78QbG1g3EYQo0iEG8Fxp79NEK1GF7kQJ4KdP1auXQuwD9i1fpuFPxtbND4f
j9/cfrw4bNQPNiF/47+YZJL3WsRxCfBVovc8diAlnMYbxFH/R0+mr5R+QDnvAQ7b
OczBf19x+BCMEqOoKvnzKiYIVFFYKDEjeQ+pXAucXXUI95hQpDdysJ3YJE9jfq1H
XWT8fNFVZOtE/Cb/Dfedk1PGPUA7u71RTOQ/+0psAD/7pAfJkuqAUeNn0POQN6nR
iNeokC0It9KkqPlFuCO2oV6QgH+RrPRg0BuiXvPN3W2VTj7ERUctt9+T6pIkcv6A
dJhSNbYHilnGoYOdoK2ZSpqImDZSxpD8aLCcBVXk6Sj1ihAywtQcKm5s8dGEiI3a
wV5USRSIgn6HDbu52/aoeevVYiars/aXrbxd9Y/AQamzDgiY1PGYesNSK1zlgeWL
6IAd6pRsw/1ll+CilWrkyC4eEhbMY6FLbgG7Ehj9ush7A3hl6qRpP3z74lcPtTD5
vDCMeKKV6o5nY6hz5FTNWshVOV5X7PRwte2MrUz9o9zhO8rX85ms7eT1mooawKbG
Jrq6Wt/n0CKlP+ovmJb00NlrIDHUTh5sayVuYf4HC7Y++l+7FZi6Air5b+Aedrpj
rGuzO00t1qHhjV76nmjtO4fJ/pt6VJvuNA8Q10ZLIAOSToSqVlw5MKVMD4ShHoVA
eGZESl48fDjrilcWaJaCSROvlQffxhCVuXeHCFljr0w8kQXtnrUgJF5g9G2eYH/N
YCttsnnykEY/P7c/yOFvglvqcJTZRiJscQncYSQmYekX7jR9Hmi+A98hbhD9SF7Q
9yhiq3SpeU9OPUb8JPAmm9zjoMM7gpCERzFEoearpKtAeZPTbvyU/YpiRP50ahv0
LbbWsTQaP4bOGne+D7dxxaCTwHgqnh9GOf0VaKfNunbKIxBJNASMkQKiSvibgNsm
dBt2kXXH5nAKgIxR4FGIhoESndwku3rI8DhyZvIa90g8L9VZKpq8Idd/E5MBUdTl
WwO6m9/9/71qG2l7RDFzw5zThi1nTT0TqcB4BSV0blZ6XDa6GqiVF3rocpbnyMzR
UMSoKrgxlMaHyjfkGRgD8wxNxwFc4Fb6iPObGdid6nMe8fexquF+s30latLzcat9
7wOHvTCQZnrs3I1UgX61F7xpzRsvUHoHX1//uN6ZKUnyLj3ATIGZzSIJjPfYpWvR
4eGSuEsrUj8eH3wk2EOOZWSKL40gTaktER/QfkO91vGQGzhhuJ5wVmRn1D/s0X65
/atroR8UBRf7zkaUKaqV7gmyKWfJA6h71BbvaZCeVWX0iUbnJf9PuAtmdaCSJlIo
fy5xSpTwXTaFKz/zJrsmOKwqcNF7uY12J8JANlizuKzZ68vURRUSGlGYf6szbdv1
y/CS2c5Wf0Kl3nROYK9CQGqPZ4Sj5Q7kse5CZTNcAYu7yZRqJJW8Eb+cqUpmnxuy
KYQY8SmIJ2mAEDoZ8TXC3daK4TIpz3GD+OFCpkcNA7khqqLa8VUeI0iF9x3esWAC
nPKh2J54Z55J6Jlr0kr6JQ3oP7cbeineZLbdcEmnbl2nMGAGDCpjAatS632ohYK3
uX0gEr/OQpnZ29W0kFvvCdS3xU68bSI9L0ht4PvQEc+Uh++dunjzXzDz2RjEw7mh
v9WiL00YX7pXxkk/1AlVZqjZzpQ8yYBsSYUD8MkS039h03PIBoUT/iuL4ejryps0
/PZTAd3nEqJ4e92lQVOMu9I4E2JGxu8oza20nEi0/9Y4iXEg6LHlrR8pn75t2NeQ
y7VtOeeN+bF9JJIU/nHtojZoi1kOK/DsokZ19zWVwguiasqIX+bqY3Y9BYPKh1A3
/GzbFW+XX0QVuQVxwBoIGVainCqWbgVhevzM67oQAODYveQr+W8Pyh2uXPkf8w+I
GC+ciEOtdue+eR3m0jIy6agw7oDYrrdQFxdIDD2Uu9Gkkpdjncj6Hu8wUO2dbStQ
NPtFrzJOeG7oni6+AzVFULbGXiG4mGmQK2VgNReZsEi9HBGvCIBKLb0M7pkTP/x6
/gWonJByAsmbVIDwymR7+Ll1dV70r60WoJ8IM7G3UYNLBWHKqW2UVtZ4FVm4GO2u
Gmxtjy52gTN8snnGybFEhCaAC8/PtjsZi5+Uk/9GnuzluRCTZJJH+4E6l8BlGBc8
KuiFaaToxRxKeL/o6cR7EeU8OGzHewEKry6XSqlA4HvByrR7/VnqZqHYrSzIDBnX
cIMy7YzPuqKBG77xshlZg2nT6N+MNq3y6oDlK8dU592LU59mXM+JwC0PRW1tvWJR
EuIMacc/hUpEOv67G+GhQr07/as3nLyudeKaRu1903RqMRgtNQuA9S0FPkyeU6rd
JCoFa/xMwN/4BH+6zYgksop5j9LYfVjhrKoK95tOSAw4N74jTGjiYQ/EsaLv0WXg
cCaRbsgzgasiRo1uuuh8DHSpI3NLf1aK6yJDInRENAAI8QmGzwmVS6bqv6QrdRrC
kbSGHMYPMuqjp0bSRHVmWZztQ2h+DzPQR47Au0fGDD+m50NJo2qIfsm4NJc6I2oh
w6uK8k4ol88h5hH9GQ4TtZ3VNKkewd7H5qByyd+GRoR2B3wqSLwGn0FcfyO1pw7l
g3Nx+uQF9qtl494CQazDEAeN7cAer4DrgmT/pN4ylSG81QREu7RVy5CyssxiZnTv
eJ+ogsqt9c8ypREyOGSOTuQnh2bVciygrIhIZW/MkGSspg7I+umfikBIDqU1SZpA
5OMngz3Ax+AlcCNhPjdDMeYZkEJxXPn7V5CFFWUZCkmiD6v/1sCZ9RXKtsL/LVzG
XkwqcsAyaKcMFCIHyota2Krr1fiNc9fhCztpDBFR9hW7E24kQm6S57APurEMYpg2
4N6EqW0i7xsV/FUnShKh0AdYlYBzrnK2LmTEt9ZHK+ik7aqvg9UJM/L7P6X1NLZB
vGkJY/2Gm5ZI7730k953aPI4H2eZSQwQJVSsXoL+lA19WictIfcmsL5WQqsxWq/F
5U/qBCppoe5s/d7TOrDnC89eChppUZt7o2Ugc6cMojVVt/QdCBXnzJrks60c+ndF
+4VDCZiu3/vqrAv9B0jxX4N1SzAR25E5mHZ9mQaXmCHSIN+sf6RMrCnzQvSvn+0m
ffMs8rnsaR5V8Crftz7dXQxXN6L6IRqb9UxPAVpk9KvFHhJTqU5N1kDgCkgTMvlt
yMw/dvfv8Ow+k+539v5wB6eLCtbB4mZEo/IHH3coyTMrnp+2iGyBkNiuKqXx8hJj
jlKSbIjWU2GXU0qRVSVGFO/VWRYHRRpecEF8rIjxRWqlGDsR+sd61sZukd1Z9FNT
T8yx7i4N+rd4jYD2/MrEkdK1Ua+7aPP/q8twRdoNiGuv92Tu+XyZQahl6xFWT5IO
UXLi11vtLBFoFWB64/BJ3YGT05Tvj4+s6ZzaeZk84vOdyKGlnFuDzJ01l9oI8TPt
QOqLtA0rVVmL2nZFFQRp/e4UTeLDLLoqFYrJwltauNL3OeEzLPpXXFMGyMk1991R
fHoQXCVKaXBKR1PT/SKnnzgOQfb/6m3OI+GAvuKxvXLwc6uxUW5yrastSv5hqyB2
1BV1M2mqN5OFhn9lQQ9+AIrgRAEccbCbhyuPL7gkCLOunJJH6sjgJ7FNvFENKYNC
U/9Uh50MtZ3LxzZXLNzoHsE3CfcL5Qm9o+ZaeS4lhRqCWRSWlnq0uqsxk2dcMXU0
X9IW09Uup1vO+moJF9Rz0KoFtHoEsPakE1P0bQnk4HbnKSLXj6TylCUaeAsNBFk8
gQ5bwFFSjXR1kynw7tVkQ9Sh/YxTd+jI6BTSWhKqukRcGPvQD/HmpTh7K7NMH2I0
6hqE8BfBYxFWx6osMpYWU7QGPnYoJzPskeFH+CSOudV6N45BbJ+gc5FOzWEqpKDd
WWMswAPQe1fXijQHc5j6cndeXoIi9NbmznbmkIC1gZMLfqNcgQAHFgnsY3VpbDUl
AftbxM8jlF3bUnJONE4k/FFk3QF+7wxE55WdpiVMz4pP+Dt09DclZCaJVDIABxgv
uuYtSgu44C5M8mlt7rGHhjNfn85yZfw24wMEEDuOcZHp/sOVotpZsIqGS5ZGpFc2
8BUHVcfZl/sBL1WdxXkcpENBmpQxCSPH2rLWZNnUXrjMUP2WXWnR5YLiwzSW/jpz
folU40PzQF6GYS9NGuIKNTapArfgs3ojfyXtRXbfGSky6qBKjmX+HaIH4F6k6TQk
SzGSp47Lgolnl25dW74qrKTaBzmoYrFdnL39MS7DmAMoSG2DAVYLjkvMKt/vewE9
77TGCryesxu6JmzRYNNUanE7jgB21zKyDyh//Z5DVAwSEe4ODKYwubS5+t9dSErW
WG30d7FQo4wwJbfLI/L3l5LuOClMaHf1CtzfsAr7/tjqvdRtdKrk//VTqZAbnh0u
BN8DoHo21f/QyfMusdve8iX5gQBiK7OPlhfjTFVE3I5Qnt/sNNQoXJGrEsiTFfMW
LS35HmvMTeX1aS2IxqX0onlTHQpEFiG9ZwQyG9BaViGnx6OUhw2b4MiBFMewS9e1
8E3MCYVo78SqDTkhY7PNeW9sEqH/coA+WcIk/gBcUpbznmhcOuyNNkws4+JxXiHC
dM/ieHTuHCZP209tYpsXFKJ5+OxS8cjLB0uV2lGav3nV7jziQJVfetEuGWyOktBR
l/XkA2voIwx+/mvm3/yAEqPbMxLoTwdZXuoJJV1i7nRKDsFJcrYLBEg/QuEN2NNA
uy/fzqvK4pePU97uPP3aDDL7cdlhJo5hHdlIxsjXeAV2ICZJPUSCiuaY4HQ3Eztu
v9DwJkXKWN+LPNhRuW8zMCygfCZ3GOcn612dHdtRbglhsiLp3JTZAkPiBbwqr28x
yE4+GxwFhpC93khJWrEfDME55KS8YZ9o2Tu6l1/cnmiWo7WMX/JU2q2bI5cYJJEA
GCdouRrMukco2TG94daW+2OVMYw5f0SpmYjpSnM3oJiu0jIImdb1QPOqVrFBq1qN
M+talJw81Y4EK97mimxrDTGMKDuyEGF2Y+HtwV7xcySO8XFL7rx9sVqlYwUZGRR5
FoOvo3+ZzVLO3gA+G8fjjLpxnrSyKDLHmcpmd6TwdCpXhZXkbOr6gP0CCOWHodD8
NAarqiBFSmLBq0g2KYuG1HxjAmv48VL4EK4y2kaMmcTShM/RBNFdyDmwbHmnaPGX
sYhmblKMMfuLyIvGrniLzFvoFskUE/Ypvaq/FCgux9gCOMib4Xriv3JjvvTgGLMZ
J8bn24fBvRPe6jYpwn8sregV85Cbaa9AMg0XM1lTL2Ur9PO2IIU1IBdznogn2kix
9140R1ZxaV23HytfHEqYnZ4/eEFBdqI035lMoRDzmaCg8ryLaJg7v/YIrTBWDAim
HldErFpLGBrvc12fwL5hJkqTGHhBBDUMUzODa+p25/d5S1MUiNfFh06sGEoiaFdL
Ey1TgF0j26+XO9LJzDu6MS4TkPy0Cm8noLOW3Xc/FeBbwtQZA5TM3SqLxpUMTF8L
MGYnKpMTlFvvezcPEyNY5XkdAKuGGE7am18aULrwbKlx3PSoP5BSCsDYD+9oKL8n
f89nbP/e/vWdPp3QdZFrOqIaojWMNCQ5Co7nDKPxKgzs2TCabjex1mHCFLbSgEmC
DKLwWgtunLxSm4qO9HcQw4k+3abj+5nK90s+v0ZpS7qdGoq/mK1JbOOn2of//VIu
5WakDsxRi3zHKNEZHwZ3CpaNhAkNqAcP3f10EEZQUi08WYN4hXBXj0JafTApyAje
APBzzoODiuh0GjMRvTRQfR4sIH7nrGQt0Y+sadywtHGCGzrhf+JJs3kr5ukEtZv1
LcSJC416Wy1sj8pPWWo3JkqLmy+qXx1aQdBGnGrQDjCJ8Zc3MBIU8QxM5w2xDbc8
/RN92Q6sQdp2/Yq1Twp7ZqMvmOhz2pP7eOOmlKRBqISyOADF39CQiiAPWGGRopir
p4OVcTN5zq6fXRzNNUvKjGAcHO7PB11WFd801T3jsORG1FM1m1bZrx89IjNRUKsL
oarHtoViHToDALt7ijCZKqPFJcCYWVb49JOpczqGTrhUKAAj6/n3AwHPhUpTbB/N
bSqt/yuT05uQRY8WAkHlXWF+0cZbS70cR8pv/NZu1g49vrGlBfT+9oaOT90GdT1v
dd4U4xOb22tPt9GXoBpBI1Z5kNUUAeoAjPS4s24qgaz20DrDtiNwnor1yFaJ/W2Z
pJvPI7tA6zP4CSE2rTVxSLr8pI7IaThJRtY2nCKqq4SLSOLyO4xcFsUcd8/wLBq4
rUnnR3TvN1PefGTprDEn8SNsOoEubD+E+90AwKZRxrWX11ZWea0SsYx6yFvPUXNt
zjUHH3XuTcF4QHZKZHSSeD35dbiKBuuR/brC0HbVau/yEtUPwibcLYOg6aoG3KT8
5yqn2z7MtawdMbraPd8L3We+UHXMVrzrlQDSmKMYeuWEC/qek6SiDRTlUc2flLdR
yPcgcR1RQZGv1apqsVdkmY4Kle5M+AqrXqWSR9JKWnsGRtEV0YPk1rITDl4RwL4e
XXOau3YLRITk6KzneRbB8vJB4p6dXlGiR6R7/524S+re4hdhVAz1CMcDR+MVrsP2
wtEs6BYX1R4AJ88394YoFmSAPs4XIR1xHoCLVm2K/4J8TT8/8rbROP76zbp4UsBx
eyfzx05M4XrSpr7dLJA1prlNFC2Z/JjmWDy/bUTzJWgI7pCylv/w7W2Fs8/dMfvH
91b9kfZVWTQbx31FBJWpxkH9P/SQpqlAkQdgy7xObEoQm5QOaKXQLH+u3zA0YXmf
h5NtJN9IF4SBt2DSFVji1tbMYvpz7Ph0bqqu1lLvG/XOLDH87rC0Sch7zgpi19fl
+et0cjWe6UQ/tJt/rlzpan7KUB4kF6PjMWS4qvwEq2M8qKJ6lpFvl3sF7TEw6kPP
oPEHVay6s3/9adksOR/HP8roNmq6aLStpYjcLnyBICSZ5nqtrChuDuiIQaMoA1yt
C/h5WW97MkJksSMfv9qu7gP5vFTaYTsZ+56WliZd3ZsQsVOi/TPucM3WIs30WH8C
X1M9EeKQJ0ZmoNlD6slFbAmerjzdNSh+41feF9FKtSL8GmluQzZGIEVvydlfflek
4/OZMVutDWYVEwAt/1GuLBiaRtOEMDj0wpkcgT9rd9I1Xz7XNqdTZTi3lMeOOmYc
cbQv9gw1RwtR8qJ7JXxSFGBkMVBxoIcOJYk0fqTVJ90VsoBA4ndSHhZobdQLe8oY
LKAwMeNk4wEfUu6on2S50IWz5egsthdVM++fDeL6Zm/GZg9XBQTn48X03sRrvRYa
cWnOdcuJRWOSkitWujzUXj0mRqbm1GaOmMQMz1i9QmXu1scrxzIBV3rykBAq7gjb
Tp8cHXFId08fb8STZWIRVOOgocGNKhhBHZTodmzvKh0vC1FZl/Ua8c96mgDmWTZL
nvz7Bo73MXRR21CwWTIg5n6eDVN6Ai6BbeMuq9Cycojs2rgIUJHRWztSI97LEHHE
Wn6FAh1TZxbluhGQV6vigc1oIUZQOXNY7w+6YrZmF0G6LZI76xpDGCjIRqQB1NAS
cyol6xJv+cVfs5t88NBlDPCXa+ooGPnLUcnF2p0rGNpm4O5DulO9JYvGzuXoDtBH
X+vIdOTG6OqkR23zPj3MvJ65RAKiMarDZCn5dIWA/2HW2cffYEjr+mdeKsaUnu88
Y9wrfQIIAV9qw9QcMF8wS/BQJ2QwPk44m/UAvooJ8D4KuuWEAOLipChzV+H2/gYe
HRSzFwHvJ1xiAEHHe09Hj883XFgLNWM3/OPqc6BI2C3vH8Pogz2LjrNapeTjfqRB
vvCfZJejcCnLYgBaYnzkIjmFcuwAsN7ZthGhUDZNK/a7w+YSXTPvee9im/LqcvoQ
+bbpniVA41X6FbxDWU7WCPF8bziAsllPQtxIsIvfFTuD3di2o0fethXtCtIDg5zV
KezQAox04hG45zLBuHHL+vwZ2WVCCHxqBiQh7YOsS8GvtoNvTD1sOk3LHNsVmuKh
XF/78AWruGxW8+BLj3R09A4gqP49Z0UqDXdMOqMDbXIYeXu6N2EBFV1qMBm/ley2
aLgun/+FmgxxVypvNqyCbsINu0ZV1iMufG446QHoti57DlKqoyyHat3kEXT1FHXJ
mZ0IAsVg0C/vHt50CZnRIbmEaFZWKTZX+umbA/SI4aQYWIeFQT2pkYKF6xh+4Vlt
OmNEmqT7ZrCYUhZArDeMXIFDpUMBTjmlmRsp0W1nL6uY4odzcg/70kbClrwJaeDE
deFBz39g8ENKAi3LUvSF+pi9uNftWcjgIus6eeIAdmv8QcfEFYjWTcZkj8gVfIiY
jin7eZRWyEBhUDx4L1I1RP83IPHmiAMBzAaec6VSAWwlVp8EAM5ygbXsFeTtgI0S
BohJyVrX3Mm+mdRAp2kDrszeo6glWKX8a+qp1QMgn84Xnz5JZh+rkJaz8xgpW/iZ
9A0UErxucxN5g1nIRtGhqX7dtic8wMaeW1wM0IFv8/50KBneR+x9FTw7LKISx+DR
ZqhGtFvSIRN/Ep8Tg5t49Db9gINY9puV8GT/wcFBaeC+Iw2dg124HeaiFGzT5axC
p6FTSW9laGfUTyIDIDn8K73xm3VNUZrSUXyxeeHo4xtqn2q2ZqT45Vi6hUBTD3OI
YsXky0Weqzb1j17Y8oa0QgK5AKS+g7YUx0kMu+YdYGPWnSODt6M6SGhaFgVOHNAq
k/mUlQRBZwYsxcWs3yBRXvkesj+3I7+qgj+atXU+luwOcBzsli1O0ZfVYG2LilTR
rQMrVvQVy9uwlgvcuC0d98xNfjBd+mke9fzfbDfKohKY5Qs4PdIFZsjUBe30p4PE
9lRSxZP/arnqhauVtH44WlZMF08BHzXzTKKLtU8c1hhRF7cwp+Z2Oa26nuZ8YUp5
Qh3mph3tdHCtX7kxjS65UL0MXQRGUhbBPuSjsT2lKb5M8K7sa+Qe+eA5CSJjuhct
/X06a+pviangJV6Xohri5zNiw36tpMYg5Jph0LPNxaCDmmPal6vg3+vP42oqN6x/
GTAE4gXfdijAjTvQKIgbVWRlgmzim0dD9MajZ6xmGrm9bHUHzhZqGpka9ikQRSOe
q37oryu5i3mbG8AoXijHsBhdyt3Mkcru5uzk6hIXwC8Zyy3l8bnolsKWmw5bi+2m
pvBkLzPTN+tYnO0meA8pC4aLnxDjGyBwM3hL8m5wE+J5+B3zkLTNHTptM3T7JRGO
bCOMSXrCPFYnM62DpJAWKKhmql4H4wtaVBZ/6l4B9N/ZgELSJXoHkweuSAsMOfb0
EksUaP0+TmVe3z+ICLuE9iSDAmniRPzWuM4Hpj2Tjl2fJ5DwpI9o6O0yWKJyx8d7
iPnwGKNUN2mSxsowWxleliA4Hqqsn0CkeUVcZOiLv6EJr7rWWQvd8GlfcCz3Tt2a
/e0LUsfC8e2JGQWEiMrJtVxftA5dpUVVzudvPFYKuR2XxDDt2xg/X6hHivITG4Ne
4APgTkcWzxkdMyRwkMj4NMYLGfk6lpWWzHm/WddEzDZwruifQQWm5oWFaKubyE2i
dAIbI/1QT2o+8a1McuTvdQJG1Hcvzt6VbVtryIhpl/WbWOndPZJ6S33tenebY/XE
6/lzFM0ieSOmDXO3f4ziGWjFNuijqPf6RJ5U9sL1UcHZgHs8NTYAYC709kTj8h0Q
3uW8R0bZ6Ra5PRmjI2P10UMwvX0Ro2lTsOJZGj3vzJ6k7o6MW8mhDp7tpcjJpLou
Np7JKPppve+9ZLTIJCe5fjztSYzP/wnv+ugCiIUAP49c5AT76vUlRK64YmH7HQdK
N+WXf3WIZDGLtwzfgGEzk7/mx4yBLx2yMjd3Z7d8GGXyd8uJpuioSnAIUJzrlVna
To/O02WrrN+sMxUN7wn4b3Lci3eeZ9YX22zAU6t5a+SadT55eZr/9s3acsmzjm6C
WnVvqvAwkI2jkTUXFvR6DR/+9gHxnRNZBVfbP7sCcKm3thjZ6NENm27rPwtSQK42
f0nA6bjlxgE3Yl1gloCUJdfzKOb1CrBJxGmaMxw5wEhl3pzh1euXZn4s2xSClKDm
3vwk94h4dQtOVcyk6QdZ0jYWLVU5MzyiuUU7kzNuTrM1bgiNxBlUkblySP3SCFbw
7eWevuh8XmzPamQQS0ZT06KNmAqcI0gVyxuCJ/Odzzgat1IlpzKLroXr0TO5bCpR
LswDp6JcT0o2bWw8/mdATC9iTykEM8YmNbpqqkyoBOJjsiBrXJgijAGvM5CDANth
Mk+qjh7aWMKOrI6aTRcfoiF6MFDnFxBd8+6znG5EhFn2klgcmK6O19WNb/5qzOhX
RChkCv+LakIAuONANGjVMtQbsU9IqypAFGfAJuYRwHLVgyHnQ81gAVlbyCrDcGWr
HaUFjc8hmF1UXeLVd3OWrt/5ZP00Nt0bpSt0Xud4RtAMvHd/sKBDKQoE71mvtUwi
1BNmu1TpUiMLtqK6hPcr/DQBfxOYPvkkeaDOLuByufxQIhmldCvN4CZLpkkZz8gc
zLLwd3qdGZjdOOcK2pNlXPs3seKAnapTIcGkiIDNp5++v5/JQ/RmB15o/YopjHbj
FvLPweIyvBVG1PYIdJg0KDUuOjps7BZCuWS37G9y0KFn6n5jRNWp9Hp3IEATyqRj
bbVVeVFaTCCat5HZO28kBWQHhSVaQ8OHTzvjZ0zWi2EHNngJMkOFWRXLPDbR+nae
ukvlWLxWTLMxR7fR1s2cNVE1gncLfqwWqBN6xyKxvYeLrGVTQUsVwk2SBj2mJ5Np
8a9N7uVktdUXuzluMQU4DkpwAdPbE90aRJvbaAzxoywQCq6SVECl7YN/qyhy0UUp
7I1i2geXtYs50Nz/gYq+JA07a/kznUGOspfFww1zRWrUAyyYLy+XZxhaWBCHLF8J
lFAwfxfOE/+/cQsS3vFy1yfQ12u0ksgDw50KPsEbr5sQScEidEnVVtR0UD8X4xH+
PgqjnLCwxwbR3JVbXfLftDyN16qe943d2wcyOhYm0DXlgDyAHBsbXbLiEmsYQKkv
hzT4pzyMl/0BTh5dN7RZ+p8Pse/FVTddG/jbU10jOtWpCXEa2BcVyAdzlzUgPpx2
Sga/RCXf2QCoeuSZtPy1OoSmAofAP2yoALXKYFFA4cWmavoYgDpgwASBPz+K2MHu
YCD1vDORSL8KAFOYQKMZoRM6vnxIRn47rWY37oMYMwpK/beEnzAHm1UxUAeJ5Dpc
hD1NCsxQH6f3itd5w0jhQvHN6OsP45juqThj4oJ33jaTRzBu/yLgEGBzrj/0xXjT
XbALUb0dfQvs5VVEivwxmfR0IYGOJs6k2MPt5lx3bAJIj1rue4cZlXFaHTBeBppu
z8I+k0MEPrxCnoX8kKvJyUyHPNwKK+8GE+vRilP86kjT4Qh4Rixu/taEk5qi0jBz
hUzKzA64dnNtNC/QJ6hF1A2kFE3klqli6U1Wsv3lBi4NP8Q5TgegKWEnG+oxn9/Q
XNDo1AMZK3TsMZ3P4/3as24oy4e9dTMG+iZDsdVOEpXhG+SfInpyfjG47djHX5en
EsDbeDH2xVaITiYfFuCxZnoF4jRVkOITnqQUDUj2WKwvBXgkara2FDfnyl/pSMCC
wK4cTUQDqFsWQP9v8d6VD6G0i0rp1iQIy666kc8PRmMsZe13/xnBPi7wPKuI68QB
4aUGY/zWSFFVz8kSujPQnyieBijM1UIx5k1SjnJbOY2EznoJqsnfsDgHE5tlFTC6
gXBy1hSHa1weqwHDAa9kkdwxN6GeyTIdhbNavYXkOeH5lVRnky/4QQ9fGM7kgLdF
/BWBoIx9pO7lJQ+CxtYk2iAd7n+jmD+6gCyvXEiM+ceJx18o81ncJrKw4kWnhKbr
92k/64w4hz8ManPVCvblozWRjn6+yxUhnAMJfKzBNeo1S5KXRTnfQaY0JarewryM
tglilpb3vfc77GR6G1zhPLYCT734FODMaNfnSKg/Y3fycPiSq/gVv1dnDqF5mIvu
TZMELId40iuidPUP5sDWPHJZmVEG0IWj8NlzyNe/lEHwxpv91C7JNpHbN2SNcC6B
X4mhR+7NWEwWOFAO3i6VPabaWtuQOyAZYUzuih/DhziiXueqoth2AEdrgxTIz1fN
EgfWuG/Ggk5HbS9NxS/DMQ8DO8Juivspj9VwNidvtXlvtweo9tjo8OVynqE7zJhg
IGTfz3EBvyXjCcQGCNX17xIDUuP/o3nlYla++xD16ANPvxq43tsptZUC8JOhAamY
GXyuPyr2MJHoKQb2mrwlVTsAr2+gAkLuroQ4ann/84+1VDUxC/nwe9gVTImsyesN
4F86og04//fI1XBJNl8wGurVhoi6RYHJ+veFtz+XL11SlWDP1iz7gUzHb+j0YJ8N
DbIhhrZHsew4Q2VQdATOaFU71Ykn6MMjU5UMSiJJKEcTIAr+5YYeTF7z4saqTZOZ
gK39GZEvq7Y4/wDyRMNeBswCboRBD9MKgrBJ1Bwcy8BCCjvImxAZ22iQnjskqpVE
AtSHzz8HCrnGfUw5r9e7eUwIfLjb5bzscq2TS7ghnDJrvD8K4nBc+WT/ZN/u9JYu
SnBezJ47D6WHHXR9ZnS1/GV6KhJKowylY4k7JQbkXutE7R6whTxzISM6xMlwZI50
0iIRq3V8r22dusKDspp3yH+LBDUSTTsqKlN8vcpCLswQoozze60hkBLhNg3AdsK3
1jRGsGh/A2F/3zYZuII+QYS9vXgkd9yLWoSAVMtQevTPoccom7VGf2JNbgvx2ywv
b34dTEaMjS5wwNTAzMuFrdkRGOpHT63va0LK58J/pq905kthM/UxTJ0GHa9AlwcJ
qrOCNJNmWDzrcTdgHMflUPDSOIySSCIc6J9wDGsraMUeHWrpkLAwQRgiMg9jhySF
oMfqc/DjugjI4jDvsfFLw489b3q9TBLaSL2hSb6NWRP+wbpMiiBrfqIGu563YD2m
/pIPwn7ooRUj8AuT8g/d1q9M43dThinfxuNwkcSwRh/z0qjKXRvjO35H0NHCtYz2
ENxBgooBdkwa18MzJeUWnQVzxh1gedIjUco7iaQeopqDNYUN5HjzXRoU5mMc48jw
fb8V0ZEtenVdzA9HH3CTEdyFUqw1aFM8wITXF32YWQL7Ckk3UMw60cE33vrbfx5Z
thGnYuZQ9GBG/ST0m/Hp72krq4+S0LA9v/P7QLy5JZkOXCxdmXz/Mjy8DTHU5uBZ
MTN0oSZNRXsWnC8tyXEfG2YB4eNoMEQ+ZyhACl6bSMFai9mKRbv85UqiiCDX7ZEW
zM0QihokXCTF65bVei/XF+yG0Pkm30h+FGw2XoqBuLk/0Du6yeFW4w/pnlHc7gC3
IPQ1BKzWIP1ZZLr8a+t/cA47uotjiwP58lTvsfO45DG4DbN1Ru6vya9WQlvFzP8t
P8UgcwvDMBL+R+od4V0l5CmJkZaerr4HByr0XEQ76alggRmptlIqQ8cqjhKGpcrH
N6v1USZQOPvf951alzWQ8Ka3Gsu5DK4DFMSLjB9L7ySUL0SpcYijWpqlQoVs4KL1
md4EMxo97MaECOLfAELrSEwV/LyxhNxGA8I0EMAvncPenIMAHxfDG4C7peil3f5P
vrICkGEmaJo3oxKMvEc61JzTzgz6/qwtA3/OL3Q8kNFdpzADh/eeGdA/7g3Cj2LC
fGmHyYShwthK4fhQYB/w3VE5+G+fNA0b9Vx3C5r/Z4Lx09ifOF1S0+/glsEkv2N2
SzjE1AMQ0gNLTxAaEPnd+9qOoJ9U6XjRfAVP3aMoS0G+fAKypV+9traHZzb35T4Q
uJKzXa1OhHwnSCEj6AkP+VefohljR1qLMfO+6S45SHGHWZhq3IGSaWtrLD7iGuPw
xKIwg8r6pNuZYgqbVPhVcrtZKJ0ot4rNXbPUnjUfR9ZWOFBbC9ZLgZM7745yd5d8
LKA6r6o6yQi9X3joPSQOisFDhk3jqiM8GQdweE5rp5tVGwRbNBdK4PwlBaHrBdKq
bgBJ0pJNePObpg7zzdP8q7f6qwuhS1JTXhK5zhhLhGMURXL3xx+KfybpC8zwo2qA
xAB5E3zcUvznRxWetjfRs3EUXuAIBKsAIizgXWm20DyJOe3//1jcI7rm4lHEr0fw
fnMB9oY6gVSsAYdDz+MZXPFRAdEkBJxPwbPxqsxLzoIxYayfOT6yaKKSMUega+N9
V1wk2vc3RLatcHCmBZufdZJOM9cbTjR6EemuUwZRypW5LiCIyYL3GRpzs8vXDLpU
7XAl1EQFUXI/6EGFpM2MNiFsBQOz+R7h1XN5WZgEQoPdtAiR7wW33V0DFVc+ap9u
3oh3EL7jAFFanwT748mMoFzvejXW0l0IIVAkuON0nvQ9QYc2tryK0kZXlMpyAVgk
gtUikNA7ruz/DVpdhshKwDjYcUvn6QkQzhk03RknW15BbidegzYxcYFTo9x+8VRa
72uaYxVIHwOWn2hI3s9qxy5kjscaJQSFTaDhuTE5cIOjGn50rvXujIcy3AkzGWlh
xzJtqqrfMadlHOmOYmmFX8bHbqKBV/+y/+msGfFdwNglvX+DWeQXT1zR3xYTx8Or
0gXAfH6OZI6W6j6mUs86JngAFjOybrM2xLVfTqiE833iZNVVAgqCIbaIXRVA7SaT
tkOpbMUUEpxmfJ32uONCg2RXn1TnePG6CoTRs3/0m1unU1begQIWhCQBZDk5cCw6
pmLRg77xB4ku1hGPMRFNzvGSnnNaIGERJrrA1hMLeCaszKEfm5fILN7ATmT9D1a/
OlkbAPFqpblWKrMgTu7wAkGZETM2hNo7XR8MmSyBXZa0YSUSpPvqJE5pIWxfXREq
JvDdgssKog2CCyVDESSgbV3YzEZtzUYhMPZxrsDiu752IyC3Bug1bJ6I8oMhBHpW
tJI/+KfuquYD8lL/2SAhPTUaaMo9Bvzw1VxWMh7GgvQBFrW+HcbIlkREvH5eZ5E0
lrivJn9DVxmYqkZGfaVjILTv/F9qx8GroEua+DSxx8r998yIz9jvvLNYZIDbXI8h
NhhSrpF6ekNSLQNrgO/zBC0Sw80MEB6f3P0C3cSwqHu0wug6Jil6xsh0KWxBKST4
oSBbtDn2A3pfloMRaLmrunIvaE6bFvIzIdqHfwp/vXBhuwirfOBDhcAwaZy7Jq8h
4wBy134V3d4YmkC+JLUdJrcquWM8SB8TFkxTeLgytvZt1UM74Isi3gXOF+zV0oJZ
X8z2YjldLK3TwmqO1SyQa0YXbYEFoludXh1HJ7R+2rGY/dt8Wpf4S85SEHN3UUGB
ZeZGByA2QvkCfdXYe4dfeSTF9FwBnXK9ygqCf5OIMmNsyP46RbxBdEZsa3NB0ss9
gkKlmi4kOZQ0kXW5pD0d5JD85ZlLkOAPF8WrEemx55doZk9P0LqdXHrgbtAnaIpV
tV7xftx843gQ5mCEo54U9tfKIxSk/QONEFDMRbtjjTslIP8eXpHk7N7KCXuEOdux
rIeYjMdkyWF88AfjEMVPRsmW6k60uZFXjX4okVpNUdDsVxLcOGtJ7O5d7yh/Jy2C
lH1AruXT9fQQtz0HwbLIUpOhrx/cUdeLenRlQwsu77gCSRHNjaUEVaNNmg/4Pj3a
QnXBtVD+lrHyp1hEBLeS6pWNDRGFwSWQjRS+csltgkcC40YVDaqZ17lb3oT8gZpK
jEBfRdRT1XJlaoA8KLmmjVdP1lYujAYtll/BxpLxFnAc7ES0asDhGw+njZJfVhAK
nmW9st6Aw21a34vPfDlqtZDW8DDqtFKvf+pZyJYQj0wk6ZU5xk1gDghjhcFngiG9
hBA9D2eCyQAJ0rOqTlzGL55z9nRYpWZHZYic++Or41v5nUiThCU5uV4gUfAYZ3R6
v7UHJBjkbaS3PVXTvYyqlHcVsudpYMKYC55W7W4bMX+zOjQgB0TyhsPtC3rHttfX
dgZz1Ycm/lcUrsloFeUWeSnU9gxQjxi7k3eMTPCwt7GBGyNIiCJ3RTjVi6fgb8e+
AyxVlQS9R+of5rM4XcnuBQ782foZYEutMAlW1wIBmXZEUrCEZq2kmubCG4jUNp6s
nGDVSqz6R2cCAzqW2kMhHXVN+X64JNFSBXPNRnwym1RLaxjH0R/ygpYMfw2XgYTB
Xk7hK1PcZeQzjpXg4VLyp4NKDlixeBapgspdF9Dnk2I5ssr+X0kL/7zBjx/GBaC8
x/1wHpOX8tTtVmlvL5gqGRP63u//gKyDpPVqU1+/unKwwDMPtHRF8r3Y6dcpLMxB
LAFzB6hs9ZZ4D5tp8Nab22Y+5w9++ENCh9wPXN8xlsRmKGiP0wOzxEFRnuRrQu2D
X8bvPHh0dt9x/geXbVeCoWpsBmAKhD41Kd0gIYCX3k5AhfQusIlOk/lzIRtjiBhC
kquja5Df+jCMg8FAM9V+Jy7QBI9neZ9jxpCZcHrnZbseX6Lk0F7h4h41SrnqlbpM
6OFWyvKEiIfKBmXfCzzl1lYvIsbuyliYTi7nti1+TTkNzRWuKkoquyUEed2LvSLr
H/IWTOYr20DIoc41Q6jTpfodj0jzyjqCcsJnP/jC9ZeNUWB7UjYMw/UisSJ9BL0i
4XUGkvj7+Go//3Kw6lNxzqL1FWmtOuwZcYhEEPxLHPa+pkurEP8JzMljVKz7TL+6
+bn7EqSq0F9FXAmgtPGkKlWeaxhtLQN5CAhS3b+M1+cGkEta78pVR3S+eWTJnzk5
Y9ebneBW3tZEH82MbRKVsPZPjmST1yabjP296KnGjKdtCkk5sYNWttsXOpepe6MI
CnpJAG8D6Zg8c8iiGJFoGUiDPWWILYpxwc9ZdcN7Nzvx2wCekmVQXWRhw3rBw/mk
vNCiDiH82N4dZOhg++2sMiW6SSDdbDpKuPe5gb56atMdKmD9PGdlzohmyO33pvpk
Z39kZ2N1Z76YwsqBkCzRyxXwsdPSfSi0ay8p3B7fRGrxcy3Cf+nulK7EvAc10A85
4bdh4NF1+RuuuypVZdFfZ8i3hOBHRaGyHRsfG0QKUdzYIcf6hbqnNXm9KBeC3Mhy
Y6jJsBmpPd73FP6ftoaF+XOWNDUYqudSLEi7+TzEsY3yafrBoE56bKWOTf6xbgRa
YrTWphWx6F1MdrmyVOxPPaP7lJCzznJQzV32VxYlxg+ZdaZMgFh8pSZtwJwVz0Nm
YVy/acxNHOGvmTA7fA34c5yqW8s5RlcHRvBK+APtSr7EQCLiCst7xPpBfPAxOJm6
KexDtKR9X5KgvrL+AN56unxNx51PrcDpHQVfoVuxzOjPnVws6vQKVsBWpdM3knYz
ZpjUPfJR3v9zNycgP2hOH3PYJZ0U4iGvM1ebIVE0n4okX7aHNkp9BdNey2Stsyak
qX+gvHvpoCNSJWLaVBNJr1t5VSyif3mpqJsqkeS8ZGsYlIHpQ5cm3QJQt0QZ8QIZ
fbfpJbnZ13fP/UcPaLkx3WqGQiEQMxGhDkGt/tpE71HnY6v8R7apF9dC8XKqmlH9
jOdd0Xzax5bzd0ww26kTfGcv3G590StWS18wdsMKfKYCbG5AkTx00Yi/y337lyMB
Q/+4ZORlUglRVHocH/GUw2B3+La51SC4kR1+FrrBd7dX59MrIvrid66tJjT2NUog
nfYR1zN6tG+AfPzGKdgOq8cglYB24RDU6kOq1BUrkLho/wHagX7okLDETLoUP5v9
oK6cNKm5sGXRNKWKhNLicHDIjyVTo2vFkLUV1fT0CiZKJhEE+mVO/EB0Tzjq7v37
ObCOYUebIMPzvTxI5FGjo5RHJChmaT0vZ7Ft5mI+uvpbhZKAOdekk1bzbUeRgRLp
ALB7q/55OlcGzXmu336g0QvfVIJbFRohWnmJP1KHzWCb28wMDzBScJW7P8lq4LYo
dzYQcLd9IXpxIxZeSWw3uUzVg9CLleWivZ9UddjSjhgVGkTM7ymw4u+n71tX7w3Q
TahCokP3zbudBWeoUVr8zffvuxygemhYkRjbPLxQ5IUIDNIUxuHrk16n2nkCSYfh
Ai738MDd0Ul6+EfW3HsE2JPW7Z9oohPkzvfrJJXf4ISf10ts5KSyCDZrwQXLYJkU
rjak2IGaoYx88mme7Vljl23DekuEl1/IV8bGhT6zhYittfQx+XGynguW3WfYtQFk
rrMZYVpiSHIjmBdN0MTQK7rVwtNHMNkGnmO0sB3S3XNOHhlZKajqh2onEqJQjSQ4
5GXhK+ifx+lZAV5JkIcfV0nEl6c+aEc8uAAtmCNxpge6EEsAJxQk5PdrgVs+VozK
klAoqN0Rvr7XxbEp+xk1nsY720v6VmwpCmfkdbeZksD5n3QUZECmaMIVeK8pUt/C
YOJ8r4A1p9a4VV6m3K3jerM8JA1fEAL3QZbT+k+IbuzvZIK78UziGok2q6ca3MZ7
Zs3/QZLcZAAB/0UQwjwQQDhLCmFMXUMC5jTeMFvpSN0IwsdARZD8AzLfXolw3Fhw
WxG80qWXj4gS7KYYccw9y7XrpH7GWQACt8916vi2B6QrRXpULjxv0+Za2fD9A5yX
25jMj0O3htBYK01VP/zL6Z/d10zMtz1gsTtImSmdsi3TL63BAwgjLGWNh+qxmK35
BHcVHEJdsiqMGgUiZOSp1Ojltb8wG3Gz1o2VqvI6t0F6AYaJj/qldVEWD8rJZtTp
fHgzTChrNhiaKrVtvWNnkOHuH3O6L1lgrk8vPJua6MLF7DoXYWUZM5oES3+DQmdn
mPyCMMdG+cWtSQwaukIFB5xCb69z1ZxlXMQ3HCTqcMa83fHQhq3JbcMFBr8VSDcB
TDbqP73xkuLaddRSFuP46oj6xS9bo9y812gYfq/GdMNL25EoC2Q2OcSwTrud3Cmy
u8Q8u2gjv+w/hDJbRdvcXO1hGspI+WZ4fDNMMVvCRMdLKfIWnxSKconTgABb6Sha
pXcc5tvxhsRIK4PQ/3pRfyzT9XqOY1qjCMKh2CHzAZB3SHnU/Ptv1c2nked+zyoE
+TGar0IQtEW5TeGRosGC7yxjEUVP70i+w3AfNPJzrF9tEsiN9jO0JwMkHQOgg44l
dn5g+QAgSI/YJQHut5qng80vEdHtwWRG6MhJPfDfMtKqrttPfGeIjHzCA/mVa83v
P2UXec/VwT3y7MIJjf29fVtYYgs/MStmfsvR9jEIjX7vM9LbjzTkNOdo0+9pjKGT
Y3T6gQk6EvEUizwzSqlTsZP4R5gBIYoVG74F7SM+RBP481SOnyVHHWtcPpvhSXiS
8QfEHrTVNv0K4cS9bnk6GPNXywo1iWFWXIGgAps81s2NimzPxpkinsErQ+UR37Fn
rtPKCNqYfN2kYLU9ATbmFAKvapWcliYaRR+ZjEtDIuP82n855iyShylWOEB9viM/
IZ2nD0MsHwF4WGTRKpSChBKwYxEA1EqOFvup2BISWtE43X8579cMVO3TXq0aYOAX
FLxkURrX8C3QPMWZ3JKBoGKmF6UhTmOMUD+j4eSJDf++turyrz8VXWVlme5s0xJt
On3XKm044xvC9uG7eSIVH+QLuJYr4FOnEI9rPbkOHi4qrGauPGa/ZFUVIy5xxxQU
LObiA/iDeWPmVvf8YIDVWtBqo1j+EieuupIL5CoAgwAnx4bMvMrws9pyty9CT2S2
PXW0QnIajXeLPyKnbkaozLqUBFXzNnv4nTxKawdfQqLxu36i/Q2Go1pj/IEU3wWl
D9G4R027UMAzm0+igcmdYv/9UNYjwWeeSNZP3S2pcXKlEbMyaOy53xp5wZC/Ooqr
1IVkSLdlnjurhuzSE9q4aXoUCqPaeRXxzD4oO1eisF2YeIrGhB/syH/4tDsVm4XZ
L5mhfrRotm06AMAoKycTIiVKq4H2nyAU7Jk8xXOlaE7nYkUoUVLRqrkyyEUnSVam
X/NcZ+ODBlhtDum4xtIhJ5ZePaPiNn27MYnodU0v/7UASbB1dJCb3806QgCGRMno
G1NRjY06dKZkTGRJjqDpEH3hvlqJ5Nzp0cEcb5u5jXq8fZDYlL6MRFZ6idK3KRdx
+mRLuZs9tsZmUJH565VK+mbZ6BraP8+wBgkisCkaDJbypwGyUyE7A41kJKFww8Hi
nNy7ETSGp2lLlMbMY+ZH8p13hDnHA6NtdX25fNBW6wfSpEzXQx9IUXQyaFYNxGuu
V5ZRao/B8QJKZqEHzS6uYxBs5NKCC7Jc8R2lyzGqO3Kv6rJoGgs10ffKqmHBRErt
AZbgkBx5tsqyjHM3ZrxWXxUHchqYD4sG4mrbq1Jt5NhihVBUy3HuCegEjsr5V8Mm
I3Z88RxNV9Jz5WSPkLHXd+6k/0oYu76h00fNtBDqtpP0cQMprYrIYj58vhCgjQOW
QCk9bMEJ54dsGBh0evEH5Pw8V1yLNDYv8L6OzLe7ZUMlE4gBrqXoWSqxXU1gh+hJ
yESdyq/hO28K3sUFRan4BkxWVgR8jWAU6Mwd3KXX5BFukDpamkmnJmFMfiPLnacb
3BDC56Jk+dVO7UYQDfiEwNeWC8moiDkYYGMhhT8WyYLHGX11Nv7f7GyPz+2p4Hta
4H4uOzqZNcAZ/SdAml4REQIgIrwwYfGS4FUa/NEEHfYrOTcOVAJx/VDBxGLvdHkJ
LFCTOs91/t3GlGgl2ZwNfeaW9JoU/UC3Gcrcna54/00oBV+6aOULkUkg9FKviuAh
Gt9/eiqCAq3PJqHcNKU9H5pJMBWdXp0vKXVOQiNA2K2DbRclqXHiTPrneCzYpXJf
XSm5Yyq3CfMXGJmNIj3Mrc/OSYhv4GqZ7yuPMlNE2GretPCjtl0Zv1BICVXXsDUT
w68NUqNvj58iVW/3kBH3d8MnvW1eiUsnOPxamrbUDBu82VYDTU29C00iL/vITKxa
Vxtb79/uHSzg5X7rfmiga1x9n9SmeGq0C/Jv0fvpt5eBjpZ3gKBNyXbjVL3+OsUL
+g95l/QjQPXqNVeuUIJcf/C/tQf1XJLq9oUPS2yXho7CaxjcGKNg0yXQKGYkw9xA
J+OOm6J7jA7BWZyF8JbTDJ1lrnTOs1O1x3ygphJNUGEAvkjIk11WblRMvJxfLX23
WSlvlymkzqtLKm4KhI53O4K5i3GBDOP6JX0JkVGw7V8EOxeQKcunDAaWg3J29+rt
GJAuTymAeI/oDW2VRU7qKNNKbdP702ctYSlWOBhd7eRz+9yu2rS41s5kA0lAtSp/
IZIq/D5CbsxUVueN2k/ahAtRxpMc+rPl+0gauzD56n1cyNsyIEbcUxFEte/n2XJ/
bDS9hZ3Q/8boD7g8MTbhImYzOpAAhKRy1OjRibdiJUx16gIkCHqU1dOZF/m5GJfn
DBhd+Xw+2HhLJER2sgbLlVod3cDIeeaaXuEhmZiTg7nSmx5mf7UetpVsPcQuTieX
Va78n/RsYy9Ldp/rxasrFh8y24z+sSVH4fSc6v3v3rCcCrii6UAVThPlBMUCiN1u
dtSNYlsMU93Ut1ref71otEFIlvv1IKq1E22TQ2x39HEvAYGYb5Q5SbiB6LitvyLf
we1Ix1G5A4qCGbEGaJ+6lkWyiN/nJRMaPVCzXUvN/GjsHOt5Cli99Hra1qmYTHcC
hnwwn+ebVg/NBsGRN25vus2h0lparG8t2bLm0ddOeBET3s2hwV0B+R+z3HH8te2k
9TO2yro6bvDvfF3cIkLV4cgFYqNgiSBFr3DebuzRxwI/FyvvJk4okF3gb5rp0ulX
/eNI686blGwIknZG51q1KpVxVVnE4ZsdYUmXc2L3z21m6LSdPNdaOTwkF3Zq1KJC
EzxZaMUjR5R8NOO0WJ1OJYOTD707gw1j75WWgocX75dyNAooaoLZzhhIpKxaZv91
ionRzHTK+MPEZrsb01/Wxx7ncOufxlmFOoYyEuwQeSwKBOHYvCfw2bJ+xLwt6TWQ
I/Lah/KNNa4ADbCwuZ9s9rGWUiN5uUYtWom36ovptFf2egfPUeIMBdnV4zfzjnlb
3K9Jkl6BimINzOJiOyFo14Ij98V4nCyLKjXjWl2zmw5bJuh2CCJgT1tuItjvzsOG
tIX17b5lYMFqOyw5zLJZvTd2Iu9LvzlzZ26kE1U/zVrd5BunHkr7nn5Y9QzjSLLK
5F7y5o3xzHyOOIo/YIVAU6+ZChIaFlpTK4z9OkhJlFxDx2toDAQy67YYOHCiwX/m
VF3CSJlnT7t2iYDZ2+h2IF8Oz0iN/hJVfiOTl/wTRRoA8EdU6oTfm0yGB/6Gnk2Q
OPqMIbe0WeiotnygRsJU5IgIQmlWQPc303wmAQ830LIJc4vawDEjKkytT9SM4MNT
As4rhztvKFC5rz2CAtKAT94UBbEs4fjp5ezUZBKUdUIkIgMBp3gzj9/lM4YGmvT8
Hu9uC19HEEeSxI5uvlQEhSR45wyXyc+EDwNZPK/MXHU8Kvek+zIOUhNwKrE+jsnh
xu0TvihxWa6NFyafSdPR/A0bzgb4rdr1+fE0ZBWCiOOvsY2fbd1DjVGsrvolWp/g
7IMAF7QFb8qPf0IgdvDSH4n0iTesChXDd2VzofkGsLJm2Gp7MQGGJsNbK4BXBxDA
8Xl2MXvWxTEjwCErEun2QwJUv8uIrQ5edKBMTl5x+wxOJh8gaKEEeyCBp/ScI5m+
lYRee8fA0QzkSWtD2MwqtjOT47vDpL6PjhG8z8V83t4UZOoo+WK19qIhg4PNA0Lv
G303cjTcSl1nMplqmpfLHyjh2mAfJBDXMcUpRpSTs2Fnu1TaJu071fjqERopD8pG
uJm+VIhMKEl+ZKjFeqMzAmnorvx+9qzi8vdY8az4hs9G45WhKMug39rCzZ8xjScT
GuFfRNGuuBqrvIEnffMRYUt7xqLaPoDS3U9/lvLkI9CIqGH5azJRpj0bMR2PTAsJ
3BVA22L8bTwqyVfIFMDqACm4bxDDHPAF6EorBaz3o4+UB7cqv0QauXLGvUsrLKfA
VbaKR554qRxTqMtxP54993To6T7V3NTpjV/xW1UsRxGskaKFdquM2zQARimwW9YQ
vxAgef62R4cvI+PQQ4ZeXFTzwyMQm1KysUWlQuxyCI48WMcYPqnpmFkOorJcFhMl
NAm3SpHF3Fk4l7Jwv1Koho9WW+uXvYlWdes0vvbTs+B2k1H94b3nLGyGczXH970U
wDTchBqXadVXz0VhvgtMdRjmZ/RKEpS9OqpYSTuPPlD6DTsT4fmmW/tkb9tc2Yr2
Xn+mrU0uj9rULkhgjDkcc05R28yb2BYTcLjB2EfsqRtjAa2ELkpMkZWsPn7F+BhG
7auVvwm3Q4amB51O6wfuhPi80sX9AK31bIN166SgzlVsGFtKtG1nu4aHfUeyTk/Y
MBnSyUd97/TaJ6Q78ptd33Qv1TOMKuJMqzpQz3K5P7PUAXCzWhgIPH7e9gkG7vBr
rxmKzgWdRbP5+IaizCZtvBrSPn7lEmYfGjJjgRRCsTxgFv3yYiI+MIqY7YLR1ooK
uQ/s7BXTeXbgE03NyX55zsIGFS9mASK4HX7Lkxunc7i83BUhYUKQWQmy27QLYkGM
sK+LHIN1jJQ5NchHzzDRnI9dYPSkxP3VEYQT9fdmTT/FMB4qom+97EIDFkb/NWB8
S9XwsbzFKVffncfy03l7kMtU3T7Ddn44WAib7aVA+62T6eVSXsKaf2dyuln1tGI7
E40/f6EJe/X4Tzkl3QpLEiGVukViOZskScIKgkcysxZ3yP07U7MaZwrWUDWc12UA
CIiCCe3rEizD0dxEXy6FfGuLqnrAGaH5WqOIxutbYOu16c3KE72q9RNUrYNbY+Lv
xcbW6xrbR/H6wsK5at7tXXiVAW6YQRClFmepXtP2FHceIH4UROFp3GKeWvhwY7m4
UTZ8h7eCTxQYeDh6d0pUS+LFjcPNKXbhjJPu1woif495WErCQca55agVrEPTe+6H
piuLVVVlhOtjdICqX0RoFnq6PBDLiVHZjnJI8ST1KRvQvop17SWLsrf6TMxmBw00
pXq291zMpoUAwVUPPoFYRAttgsGufybuDrSbZGyToQ+2H+QtJY1CXjbvmVfMCDAy
pPvoiLXiIE3wkG0zSNfW1Aw7spbDR2a1NXuGD5te5tLrXu5TfZrOHsn+TmIvPXX7
LbssKoh25Yy9/D89NLN4W21j0wCevhY5H+k402ZmHwWuwB//PCnpwMdpm3fX0Z7o
So4KB+3hpL0ZfS5dzw+tG7oH26C1z8buwK+15Q1CdyRGRetBDf3+qlVt3XaBsJcz
6/hBTKDZYGeysfE/wONVIddg6q9ooHzkqPtvl5UeroeMAlMog3CdbhdUq8GxLfPv
lKzFMZkL1YTjNa4qGJ41efaNzIMUXS8O0b4odYVydxFMkhbefff30wpSaplcGhRO
B5zb8fyMblUL4IPnpleiuSTESNEBHvWdVlLggsLowiXZIFMMaqZi4rNiMPe2niFB
PiMOQyeUiMal/652OhCMyiJX2BtWfw25ZR0i2fp+aZ33lGhR+WbBy8oa6MQjGWwF
T42Li3BMZCjsRP6inIXNeK4UAi8kKeQBkHN4dNy6Nn4ngznPa/n+Qa7asDFjBk5O
zpBnUZg2DbuGMdzjdEWwBPOLkTVLnEVsXTowkM0C9jVF94nshNdUhB0aoOL7Auhw
JDd89MY6laFtdQUme3pi7nKQc9AJJenUQxwIzkvOgZpr2pLyBA3/LB2mygkPNUQR
G891QfK9IgbHWbdZyn37lLyFR1H1F0Gga9V8CLW8IhE3y2WT+MYQWyBUZ8ADhRGK
NNkJ7cP8MwlY/9qGJ6cDydf/kvp5TabgmQIF+1fnwEhFJRZMB0qil4V6wiXnD0NN
9Lhqu7SnOCwuuqyo8sAmXsFDaIwoTihaeK27lQV384jNez30JicLC9ZHouVTpHrH
sBeJZdhFYN9Db9WBDx0bWLkBCABz/xIvxoaCdjxRp9fa/bKo251pkucUC4EZoMmt
/Ywk2rBniBFZLUuWhpWcat+pp0lWOqZf3cLrP224Q/PHqblGgJYNAcdR0XWDTCGh
uk5Rf/FONu2+GEPLkP4UfPFOLId1N/wAnWwXg9ax+sK3L57c/p09FbsKS82ldic1
YaLs72w/Pnz1m7NU+RLahUTZpcJVV4/ItNRCp7hliJOj3s8qINMXEh02GmGE9ktT
2NUVzzvzsDM7MxmU5Kt0hcc7NhnqVt3KLd5mQcKXhdw6MIMwbRaUuma98gFkQNBI
4S6RKzAKWpJF27LH+g0w8SLVCexT6Sqi45ngvynlSbIQlPUmRSlk6z/1M2nFMt2w
3uUdNMqkI04vILPDE+GyBm4QYs8GaHOONCA4eboLB/qd+boSMmNQe1lgEZjrzk+B
buj2NJlUOTcLOw0696MMNLbvLJozTXGa3uLHABzAmRERJDjEzCu49uJ7JWI3VAHG
GR8ddozC/rnJP0SgaqMZ6PCXyE3qYEjrpYf7D6LaPKybIsPgdQAEaPx5qqTkgz6d
b4MYQSynJvOrbsalzV0e3XkvS31jGixLWbtRSRH5PccFYQPsXP/4PWnmDXVoZbm1
A9W4nB56Ai1cmrQIYLHyon39u3SZeLUxxM8hokgWKwtG9QUTb/MjXvHqYcbyuwKw
76i9g4Z2WGHM+vJY7EeN7Hu7NeiJHdEMfGPPySRiiQmrOa9zg4H2m/aCsAtxcMkt
Lm4XxEjyT8QeCTBq+gYgmXGi3TwpLYi5s3D0eqwAb6aeYOHi5AY3BW5mxCUwVSYP
J152SQ6d5UYYZcIf6wb7Wkah+ZoLA8wzzwCSQaYvB+wZGJmdrnDZtPdeQyZ4DdqN
0xBLmcZw0hYSOOWu9yu2rD09X0elw3MNhDzUHFzNjl7Uar4Du6QIV+7aLJcgkurQ
O4QZfV7n9XZaaVe92haZantZJMG/gCwv6FBIKevH0rILkkP2scnr0vXFznEvTdjq
oFasdAj7cuiuTwsiRoaaLzR+zn1GFG+OzGx+29bAFDGHm7YUsi9fWEm94Fj+LozR
jPEpNTE2UrWWX9H0ZBU9kgEtmWzgKvDPRd9+jUE9T9e29YOD+Ux9yMKqOZdm18mN
+S0DIs3BbLl85Ug7QIgrI/OtsaVF5cIhwXFzTZA2qMTn0EGiOwlIi2ILrzMlkrcL
LGG8ydmIyeDNxcWWCGYQxAnnVkbsYwFJGQ6NsbirzNp+cT6nbfY2qp+SVnD7vSSD
2n69/6rjQ/6s3Ph9Zlf29VQ2chgJXgmMIhALiM0Iln00C6VlE7v8qEURGBY7VzuH
78RIRReTw+AuphPmiKSj4DEy8GnA8MZbLnW6k5nj9pvLKkkspKsLz6D5D5rMtXLt
H/7WZ9ibK5zIpMT0lINkJlLkrlAMTqqI++NVJrzGE/N9oQAtC6MmcT8qvJQkbNkX
1PXkDHJ29Zl7JnN8ubtPMrR9FJdAe6GL12C4qcpsB4AUB3PXVEKKltVYQAhjDCCH
M01DRKO86KWU4nWn2slEcR3THR0usm/zohw2klv6m61ZQBWjkxF2hpNP3WfqDrv7
NlQtulgHYRL3+bm4D5ZvQ9EjttaSmL51lCYcsQH7F9+QC1vtnxorln6Za/I5YYzP
gNTPTK/UQGQF566rQtrpcqyh1q6hM2ZTZZ2Wk1RKKDkrOibmLnaSWdmGjJkwOQfz
4qpWl7MW+Ra2fTKrNHJn5Bcs+h5FtNo77ckVUKVA6rkfurU3Va/OABO7j2dLER4f
qRjdUzPnFHxLVzHtKbm55+O5p0pvR3Uv4qwG3iA7BsSMQds5bBIoRkfkSkWRPL2Q
YUU5G+8W9p27JlRdIrs2W13xcULxiX66YNYSsndH+mKuId3khyAlfWz4NxNSty7P
36aFl8drJ0iOmlD23mSVBxK/vcv0KB4Iw3KdcbZ9CU94lopvxQ5FGNfrI0rzPPhE
ITkpowggb9DkJ87X+ikMO/oWK7yTvnIiX12geAG0/VaMZzeC5j2a7fjfK1ibu1+W
ZyzwlUHNWKxHAW+Sk17IhE9fsKwwRmJUfLUDtHuOlCe1TPDjyZy19xYNc5DJdkgD
ETxn9V+9CYuc31ob19XDo8fGNqHCA/SxPglAqnBJ/KxCVV4o7ySbW9l1cgCpGXrx
3tmOfQ8tRnCOcJXYviqpnIW2PhRkZGSoYmzqDCrd9pWFImOMyNQ1NHN6bOGPNiFQ
KBnMcLDThELWrzXOpa5wbDJzMgWaVIokcqopjXlUPOoP2mpK75M7cYKNS3uJADfB
5xVUzSUhtp00ymG1klk2rx6xaU9rY5siNMxm2VmO3ayxMS+WkkRyxtuhofkamkcN
GzcbQb/6zMyBJRvszsCQseG2trtJhXcazD+TaGjrw/tBGlT9yDEos+8QGhkTTa5u
Vn9eD6GZ8QAsqGNk4Ao60rONRDkst2Bl4VjzJ8FOdx8a/5K0QPQxj/WrlaPO70bn
81QgW8uj2k0KQEqEhiVWkgN8y/sE2V2MoYgqw6+jIxx9EAVL0jHbWQZRVzXzUogj
pCBcXQZJ/8eVlDxu4Ag1X5MbwscFAHTS2Ac1wRAEe1On9FkNq6EKQ24Yfy65hG8L
JiWdwH26CfoWNMAQ9qaGT74ArnyNGSWZsnmgYH9qengvTT35vOJ17/4sUffHGPQs
4XtIhOzOqmk+LiQEhTyqh6Cq5wiPpZa78JV2Q0jJrhUIfy7C84xF3vVd/c1nbvnX
tU/z3NrEx8fxsaYpc2YUTSWfgQ8EIdYTS4Kr8sC2TAFYcBCw8opsfnLDnF5sxKB9
owiVf2csvIR1m5t4qNsNhCJywPCF90GB4St8B1NpIxMhc9QUVPsi+CHasLqFIiep
Z/SNgk7PIledStNvtrB+80Ve0zaf7ZDg/iQqThJWjqjUwkH7+m8pGkBFxy2eea9V
iXDmo4P3cbdGAtVgL251VIwJhcAGlvKpOjE+/jjT2qCqNEJ1C+KpbIOEXefJEWwm
zPpgNmhr4xSL1AoyjLinrYdn4iPCiOWzORUplBLQpUJqb4GwMLQRz783kPl9L62g
yyiXcj4wkIJOLYzN6OwjkopsDOVWb9W4iMX7K5PhKORH4/FeIPwR9iQlufCOjZ2W
uhPl0un8t7uPo9L/AT7gJa7ha7j3tUDCXci5/gJcer1fwl0ZfPBVm2E1co5uRJ3q
cRkqQjbdT+DYbcKMMwRSrG/INX4NMc5mYo8GKdhVo9Qqjq+RHwq+kPbz7H6k4uU7
tYAMppCST1C5DfSlMlHBENE0sI1ksykkj2rR2ReJwjX8ssg60IHLbsM4rUT4ytQl
27Pr2vbOo28sE1BY6nQUjBghV/+2zRurKsSqVu6ulhYU8FHqss3AwVHJkHiweYWK
0IAv5SocRip6w18cPyeSCHq3CVFD+1ZEKD7s5GewTXNxWVJARJ8YjglWlgg170QI
lG+VIazgS9vlt4Q2LLXpG+pWCYO+zzTv28AlFpSRDjYbQ4pD6hSoyE/v1GHT9gZu
Qj/hqN80r7eeH6CYeKZ/nVf9x73cV2RsOaZsRmDlJWN+2Ap4ixpOdxoyLfRLHJ6d
m2ceERgH9n7pFE6Jb7/3zQF/4O5llcHDVJ1d3yg8kkrgVf0tJfo9GG0dWfCGNq5g
b/H5j0NBxCJs9OnsALbmHSyvN+xQkbB245SZRnCXMzRz04BnCKx1pH0QO7DhR1Xe
4LVC79iWL7aD9QO6jlwpPzAKrpNYIIvl0QGKbvJuPXSv1FDc1G413iJcYaMKxb39
60uP+srgk7qNqpIe4G/6ak7g6qH/theMdI1euVeACNsRtmv5gS2YE6aqBCXYoJXw
1bjERJ/G426BiweTwGoroWLl2qfLGnNwoDkfel3hqZrAY5c4ikAnMOf0ABixBR7/
PuSekdPZhn/bAy+TvntgDZdWpiVn+K8N/sqOS6qtZLE6evZlIsnXezv5ioD0aQ/o
8D9g+QaJE3rkLsn0lSZtYfDKGD2eG4v6vL4MPv+vBhaJLROwXzokBX55BUdc+Db/
CYPq/wtEfzzlTz7G/Gewehb+bQUpeRC9adrd9Qv359X8MHROnHfRyUpvdVtjnPDn
O/bWoinSIChg8pG9qUCXky6hEdQhkZcG7pizcXDzsFRJEfZwwJlrYa8NJq38h23G
XAifO7f6YXnmqylJfVJ+WTzoH0n0m0YKqxyXvd33V2H19cBQHhaaJTco2Qqnry/2
v2CTNWBaUJe5Dhg2ksPw4Cb7bUUnt7GY8yotcb2+CpckImVq/okvMlz2yF1uGaxa
cXZJkjmzbnK4kulEsjrjyYWzmIPxsD8Lvd3wHEmrKfM16F+JmMB13SvKQvN3eZ7r
s0KW1uPGyEo09zHyd9H1DJoFDNU8kL5UvyDS7bDFt94Vl6X6UFpBp3mp2JduxHa1
VoBGODWccDEHJEkTbUJYkm5BhQxF1UNp/K78WukYOadpye3ihrGSlFzHIo7XcLnL
Mw7esQ0bpJ3NXDQZ/QdDtgUg6P2N9obuZya0HdlcVMagzjW1NZk+9E0+10ifIQ8m
TgFRwq/vQgwKFmyOtdYk4QQDBMIAjlHsgqkt42cV5atHm8Gv9nGeD6e0CN+6Bekv
FSkJQkSETd1k9GZ8Cq8uFr10v7RtbJe655fiLlrbz9EPL1he3AeEjRIHViWHnjwq
PRiYf+M8BiLtatArQMrG0bJll+gR2swg+0xhPzYYN0ffhh2203/h7q4X3bS5tmbp
N2qZgd2adzQRXTslirKehvNdwv4kGRTR1WxSEqgYGVJ8o7+DFPIwPFi2ZL6V+ApJ
mj5/AHcBvO1D6trNvYZbnGlSkJUJ5EHlwc7g0y3klLIVuvDzp2el9Udqf0OD4Qnq
TAU/5lDGISZByEY35Iekft3fsy7GxAX7ulw2Xy3w3UU6XxBvWg1lOPgICCyJyZpc
7Ho2K1Z5ZawGTW5W7yfMnZFuUmlmbJbiF5UMwbzhfQOYH1z9xQphhgAzO3mtbcig
xitXBugufy47UNxDwfUskEqH8akhlvvYjdi3LFgOqhYO3HKxwTxvooKzH0YwL4LP
Q/MCo3laVrTJGwiETpssgKcHKCgBzrgdTd845955uaA6u9jBPUrmDRqqp/SAy6IV
56PnXRe5gsqp+9p6RYWmfqn/LhdUqdXsC4SqtyjnaWJ2atL4821z8YC9jDZJ8JOE
7nOqz5TA91Zq1pon5tpn1RJA/3DcDZ18uR5Q/zwhOIhqVnhOqoIbV41HHg7eS43Z
n+Zdw4A54+gM3LptZ12WZ5N10J5S5m6aEIUV1NOkQZVNP1zknqXFsf/+P+sOi6Rp
N7gKkcNhPnG+uv/WedYyTJzqHM9GJyjFdj+T5QvjoariDkUqNpmenGNN/qCx+3Ge
P6Hbu7Mz8NElGs7JLeqX/fnTE0INS9sBY249euQxnMT7ikjZW6xUtMDKluSaWJek
rskR2h4McgLIS8CHOS3iHebr7FbpOVwVWlF2bR3gWAiHFc8QGPxiSeLRoo0PfElt
J2bwVK5flfctcnquHrEV0QoZazOFh0PtwVQhLvXE6YxUrtOpv5GZKXkCDlcJPs8K
Sd28d0SLkLYytyxVf1zNvaiXRrFrkKCJ6OKbQoLsw63FCQ/6YparkkG+GbFhCqAa
mNjigpgXl8hq9WCo85MziakU0fa8BAvVemYBFYNwrf5/WF1ruiRsJVYBSz6ZVQp7
3rIwlM8kyYBgMSggJyfGJJioY1spEpo6zOt2vXtRjApQs1BwG5ISuZ4qh8F6VQ7t
tUB0qDwVp9QKUn6L/YPtBrgtscrZ5IeTrQT0XxnmuvJQTnpiEERyspGlDxZhwVdV
4bd3T0x/Qd3TCXSp5BCeCqbCCDpJNIlhZD5aZ1APfNUepIRT3APe0c0sxNZQ897A
dwFG4gNb321jgh5u+u5CphlEeQjwz7GFfGDRxPOiKUVudqaQ+YK2rIqHEDCkJTcM
CbTr48iITr0cLI/DVg5Au2gsy0iA/I4lASoTnUTF0odD8aTWQu6cvn4OtG9dxyGv
KYJm9Jb1HadVtqWVXBhagDzkS0vstQeYEcdjNLVX/X4cVQtN2t/RQLIc4tI+85If
u9Re4r6rjCWEdIB0qg4V0BMJjKb65I+ZGSV40xXl+6Qyb6bB4Qd1t/CSEhWVjkOD
ypqLS+OO8PbWLmC9v/UmoQpwIVDlaEp4EngrYPYgbT9Nzvao0yaCjhESgNLsyX02
Ye1O5PTOxqZHOYBU7UEYTRBDdvbYxH5EnzeFt2FOQTHqWVXq3pAiuMS+ZBQFcobg
O1t4hf2ev/GgPAnooFNJD0EvV6D93mbX8P3GjbPD4sGGjxpPhm6nqAQ7X53Sbf2L
A4J+vFc9kUyzdBX9ttk6n594WBpVMuK2ysTqGrtOJ5aDfeLPsV4J56sMysKBh4Tv
RY+1mx5V05QEdUGe7b1D0bDHGPM6YwsWdHi/ttaub8GLALPTLMEZJ/pXNWw6vy7L
MY8TUZfBQwQ6F67swcFA8vb+TwNzs2FTOFv50stggjXEyfS9Qg0NaJTxbEKuSOsS
WO7Tw+NDTdjJ2klYIi8ukLCK6WsjmjU5PaaZhEPkNBLDaLKjzI3z2kciuCs66Yq7
p7NAc9I7CV6vINMUI52E+/IbM2N3y59yP+/nr2XqgKyhdlMWxWdaB1ykU6FUXCzh
mYd/bNaZJQkSEB/f+ov6rohqQZch052Fo66vr+FKIoJxpBuWPz2TitxGYkc4UVYl
WwqQZELCxT5OjQupSRNRmxXb8HkRQqsaYyhXydZcz7q6a1WT7nVqPz9Z3N9XfJKH
WJeGTtQn2PCSCEH2OgX0ZUegpHXevF5dyQommmrrzrwsoiS0vYyq2YLpsi7x/WWD
VT3aTdieJDh2F/Kyr1uOb1jQ0EEJjKhkLmymr4GtXrZGrALxO1K5Q1xa+epRm0Qf
L23jqxzJFzfHtzfegaB6ZMtKVlhODhjzkNsCSgH9O/WuyOFpApweJetAHrR5vkTR
4+R5Yf0EMP8XHML645/Xb1j1K2kjOMjjwon4a1np6owahhPWHW6mtw6VrLF66z/A
Vej38+f5K2J7sWyhbEdOULBsqdJklxQMz889scAUx8DjFlpVTr80LoH7APBfRYCA
fvo6r3W04LKxx6uLgj473WiSsgxSEXt04eY8DpFrIGHUbMVeC4l89ammF773PKzk
MkLipI92M1Fc+MIIGLV3tk1q/Jt1yHgKE3T1AEH08aphg0wYZaMz2oArE27r7zza
tzjZ9MRMQ++W6C4SttmoXPhafKUd0V/Oxas/cWDql50gcFSRH3fRsLYJPRw6y/rx
NhAcNF1iOMtalOFlqMVzMbMnZaBjMk1ERuRIaVvoGBmja477yOB+jMnwSHF+bGiK
ZNU/epuhkbg55NdTulpyu9ZGMx+dui6LWGZpFPnnaPJ/vovxyGxDn9JiLz7l24aO
ZLTz5BddAmRi77IiT9Txt7CPOl53ujh+XFtC6ZM697q0oaYO5OtJrq5jdfEyoswJ
8lfZptmGe8gvrlIYWS12FvbT2kcv3k9cwUKgKcVtBGSMVvI//Z842n1w+ZJNqHWF
I8btBXjVI+uUVlfZ9OuHU4gmcV9+HyG74vhx2gCG+0LxE/P5cykle/I3ZdAas3t2
0ub1nFyxMMhwLF10NL7LJsC4eVNpgPHNa6cTjdjaNZ8pC/MgCrSzZIuNgCJ6no+T
UPhfHN31O12AVo5DxZb3ropHDGwued1LxRQFcQLcqMROmX/g5bOI3BRXUue+cVQL
j4nwwPdckz/NvSEbDwPJNgt1yyNKjm+U2/7IOo8PNP7rVRIwjyflyRYEwl+w5Tmp
IDrEM5M3uJi5sGmV32MLwz57zs7Q2cg2luBSsQz3O8jf5UVIxqzVClW10d2/1Cw8
WbrUUzzDiny3aLvT8QdFwRBQ0ysXJ72snIK8SNxGoLkrsRIMeWrciOFFUwVfAtB5
wg8pXotmT0Gnbekki7eMqQ==
`protect END_PROTECTED
