`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OzgCjjxKk9IAQEzl7ER8CJpG2keSz+ayOFdZFUEATnFYevuhYqwdagi2skrh4snY
nPEd+joMut9zBM8cUs7T8MZazgzQcBt+yB5qgSUTgpR8cVUQ11iKQVpVtmE31MAk
eAGttRBOAfRjInY4ZnP/oim2k4P+b4UD3dVX+xX3eYc22Pz7trOb59tt2GA4K5oI
S7GQmbBFoGtU3sjcgMnjnaH6Ei9LJNJZ3qjDZlMt0XrfP2L6m2YSYKyceUL7NE+6
Pvo4d8+JD38nmGVMTLVDwDQmuiHzaCWZ7F0E+z/Ec4z9OOery6jmgTfTqCt/y0it
tF6UQ0rKOQKZGVvzYFZ0XxSb5lDuIxpipIA983byehnnDqeAt03q7d7ffAyoqwE4
MC9wStyhHvsyz5dhySnJMSVt9hpV3lNkp6FmwK1yi6VcLDTeCYCWAmIKouzBho6O
EZnkL7Kyjq95tXRfqEDUkWaRYHGOESxatuQhZJCMUSBU7CqVCvCSHma9+RZ/l3gD
y4hhh55y0M2cjINr+UsySbmHQcPQvXxoEqc7l1FOqBFT+ZSPQSw8TTxPd5Cv/zDo
QuEKm4X/Us+J7EeepB6W2Q==
`protect END_PROTECTED
