`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZPVfKH7WIezRtxadAc+LNROB0w1Sl2rcSdOpbtOSHOUxDTNsR6IFJMwG3CwqjEC
JIHrwLHphGnMxoGpBNPZ790yvY27ebSv//bnNaUxFXasaBy/c5wkAvvpYPj8Fm3t
HOMmr9j8V9cW3ZUjlrnwVpyCSKDotDqRIJVO2EWeZHyTrwlSNYFEoY9vQks1akJj
XCfA+AAGi25S1yhmiTQKdHGiqfu26SLLInUu5Fy0L350Q1fvbfpN8217DbEfcJR5
Odg3fYYQuFesoXB63lR23AKRZfTsnS8mycWc/MFqsM5+bKRmEwpQ+P3B1dguYjqm
PA0GibFemJQanY5WDOnruv2ypWgqMVmmwTQpklxWpS12qipexKaULF+IV5sJ33FA
sopquAKtAb3QrFjCSlFYfMbp6CoEZv2WmNsaobEn3GXD17GpKKIMudQlm5ZpUPtC
n84qiRbMbmxcGetiL8gZe0h1YbxHlk5rRr9kem3aq4lI4ob1YlijfF49jkIhVRoW
2UaVpG/UUVBpt/8EjfFbWwd16mi8OGjRq/fQUhrxfu4vT/6PnLxubsA+PvCdpsfj
RSV3r1yLKuvVcx5ZbqhCxqzu0xVieSaNGEH8UgT5pcvaLRSFDGCNiXKyte/udcE2
zxVIFA93gZcFE1h/fLeeqG+48qlm3gFndJDbLnrpGFX1OXjq8BrrzvTX0aYWp5Oa
jFXn50CrFySO+XmDQMkylvJ9nnxdt8ACgGhrPkTjjFIUO7G3F30pLjdyzbG5Pazj
KZYMi1fkEk1gYORIlGGUV1UCwqVPBFBA8bAGz9BdEGmud+Sn8tGYqO/IbXui4+ky
+8PWG1L/5ReVfTQc+dcOG/5uzhlI9lqqnqgGUsCv5zioXMYLtK5D1eHPbbDFhv97
bSNjVtDxjiy5oY6afLZrWUGFr2AKoxL3REEN49esQFbKZVHKqrwcfXtba9r0c3OC
xMz6IWOFHe4MxR0XkP0wDsMPogfnqbAvAcFED5jG4TF8yDh9+iNJT00yu4AnqOum
V4M4NuTIsKy73yyTg5hAbODzQjqVDpr2NYWcuAgbykA=
`protect END_PROTECTED
