`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0q17b29BRy52fJ7UR6p6NzgxW46AMXOhfSkQSlxgrBbs6ojcUU3lY2XAatdFxs+
bXBuryu4M/Sy0YNYNGzZk0DL1uV7OA8Zvx75tb/UN7nFt+ZP/Jt1+CHOb3gylFmg
1snqs+/pzxxV0a4Cvtyf+ZfMFlxCMx6R+A5bp9LnzqoOq/OyX5wN7e27iXrni9mp
3hDeRuWoSTa9HUyChVuHe3tSQmPThJ9jVHjmCf1T+JJrtsM//TS1ayTleNN+Iqpw
T38wQiK+7N2wOOc0K4z2G0n6mFPwb8DKdbxyc8fCRV5E5qwIClHv80+c3hvIlTuP
q8i/YFfpVZ2raixTcMgnidVYJ63Om5iO4UFsFKa4Y25oBt95dqW9t5zhYpcbmFis
Qwn0G5yW7X0hm3Mp2fxLSzkBnmkOdRkfld5iONMgBR14Wtovw+x7LzJbA/m/aEcA
1tOJiBdTDoibC0i199X3HD3amElwnbQbMGpokE0exBDtCndXpJxGS7Ge9iPxO6rl
7HCatkhDVX5yhfA1EopfBlqFeL+UTH4aH89hscTUJTnCaXemONMk5fvuBUAWRSIZ
tG3aLMaehrAyTsVOCbb6A+vqW6BfRiJOWRUQSCyri5k=
`protect END_PROTECTED
