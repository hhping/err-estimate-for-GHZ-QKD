`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYLk7YIztpI8+zrjd2LEMp08pMfuYVH9KZzWeVZCTwebxcLgc0oOWqmBTB+qNNLe
yNSvG7NJHWsRpNHytxSSUyRyR2rqPlNgTjAOn3fmHN/AoAJG7Qb3rePKBA/dpWRl
QXtWxBYASkh5/Z0zBpirtJww5Lm1wqXshuAI10/0b3d0wkxJgBRlFQRrqDtoFCF1
VTFMDeHKem4AfwDjZhfRH/yaWRTcTlSJkVq+SGII8OJYp/If0sijtLEtZCmwxDGb
rGrGYkJUO8zkbelrJjbQBY4XvvBfylmTACxjMWHbwcKe22QVpjL68FBeSsGzyLaO
VMgrd9kb7gIT3+qlPwfnvR2Qdz2WdaVyxLNK8IS0ox4GcelNErdgcnybk1msAX1E
k+PJmsgFZ5XkmoGlj/NrL7DF+xAr8CH4HIOIrq95h3H1kFcsLQa850JSlFzJ2Ept
8t/KY5Uci6xgWC6v8sLuVip028SA4Lz8Yuz5LGN56fo/DZI5vbylYNenvS7bl6qJ
Nd/+JuTS7wglFtwBO1uWjs/MIVTmn69iZu7T5JeK6gm2cy8QfDZI5JmHHq8DctM9
AJyYSMNfZ6hJcq+bXd5/R6/5wpthdBw+4HR8m6F64u3XXrqiqCnD7h6zvIZwjbf/
VKeILwJ9ZTO99fvk/cMqdg==
`protect END_PROTECTED
