`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnhXnVdtpo9YDfPA7zXcPEoHpZjnHaoAIlOYiIjnhI+BttwZoz4ysMg/DbZYVsex
tpJqUQME5G2NqIoN7YjmAjbQ3wnkHsd4XVv3xjxcpaKuimGTe2I1t9l/XigwZe8J
ucBCoEc2qjD9hYsR5b4j2vOzQD9f42oea0CDRFge238EhAyxocrBuSi0Gq2lUncH
kRoAk9eAbZAKMjxP/Y5/IB6pYqYLMeZkDQEqcCSMxRRPWBLCyAF7XAshthclkKyg
ERaE5TXWU4IlL2KusboBdwpDnKHpswtoIxUEzlj4OAwVDRidB9AOOzvQC9MfthYX
BFhdmGBrS+SDk+JtRkQ4aqLJWCSFSSfHgw8W90UUAS5c5Sx+arBPBNNDpdlaBTp6
AdUM+BbA+IHbP4l+GU8o9rETkMuLSnLBfP5mumSTG3rJu6FXS30FDgtmDBk6SHGP
oLAIb/fkX99izq+CRknjUn65spjhOSkurHrnpTOC+7UD2joLg59l+5Hd58Syr0/Z
tJJjc6n8wOQJlb11oCVV8JPuZL8KkoYsfqmN8wu7A7QS9eyfyJJKTTcotsL0Vw/Y
i+gvbYYXaE8dnYvYm8BeuEbZ97Na02nPIWNyccMMIYZm6CbITNpaEGwMqk3NvsSI
+pXX6itRJiInMO2Z8QGbab0z6h4VDbVzyQSkogynVFF1Y4PU8M2GZ6fHWovyWiXG
0YHyDrl2Ot9DwpaefMi+1s7jJMgrpzF/IfzbrhvMqvjIzTGbtEaHnG/ApLa6if7Q
f5g415nRU2+2oDMlKXjMzd2n60OsX880T86wKaUU/RFXc9pnGbJ/O8UPryRudqq1
O9PELOq0svecpNiG9wEfq7lQZISmbno/zLj4c62i1AKxV4W7VLvsuI6OTeQvkTD0
BJIUdi6mxECrADiaX6GnxD5BylcjGUTXWzi6zlJSB+6Nt+I1dMv49EtMt4EXiPZr
8IVVekMopPPUwfFPBpbVhO1umBpFt4vF/emKtElLqGOOg3SK0+m5/ad0XcgEIbHd
ooxHzrSHzheq3SxxyQO3kYCGezzZ6THeT4ediwUGtwuCZJ+XS1xv49Otub1zvAIx
7p99KovRuTzNdBx/pbCZCucSYoXT+v9svL+EP+OCLyxyIsjN1xJqPmMSxh6u4ACp
w8usjnGJP4+ekNPXi1dtb76ZvNwY9gM+RfDcLBc5Myi+DjXvtibZKQF2muljwX4s
4Z6meqTV20S12x5UFXJtGH5Az8d9saaRfv+tW7wi3Fed8VesCAs1OasDfo69sLt8
KoAwfaZnAeHLXFf1KC5cJeLI7BI1FyreQqvv5QHDlUNCVfZBCktO4krBZ6zguRxt
mFVWBhibh/fZcmH8v1xuB/tiw3lJoPf4GlAVsx7LkMQW5EgLgFogXNS7RmMFY5c4
7bLoEsambL7h5RPPLG0grmrZ6mn4mj/7UsHzpIz+4eayZ0VnTzJ739OSy5VPHxKV
wUdufdK62fwdA9Zbhn76iM7cW0q/3CA4YdrtWd4IcaYFQPm/14I+i+JA0jEwV8By
b4gwVfFa1/AJjVlRYmRNFtEvejHsrjrJB0ka84BmZFAYKKpE3XUqNsHbZaoH7dz5
OidD1UWDn+7ZK40MgGKMp1I4irDDncKXZymHKkVhtj1Gvfm7rhIK7mPwrjIdWXp3
SYjg19nnyjfDlRzwZWdHt0/UzlhzAdrRouj1Cp9VyKSKR3HsjPbRjwlWBsEOcswJ
s4MYXvSeG4qwS54s3vqY7uqasDKb2gMCQRSOEx2/M62va/i5ZizKzX9Pmdu+OE9N
NlVcbTMf2zPdKDbDkfvRLOEssg5b2cPPY18XcdaofN9eoGWTdDqdspsYDFjVySWg
eZ71Y0M12h96rOhX0lTyF/0JOhdDt8z0cjTvVTMSoVaBVlWxskmnY24SYDVlxS8q
pcqhig5O3jTACCzVXL+xNce8fOOyLJ/+des2YhOTWaK7LD4PfQobcZxLnbMdPKDk
hvTmRLnFRIOz8Srt+bQPX3hRF02evINvsDJK57wmvdzDjSUwT4Tx9aOZf456wSBg
nNUQbQBeXcLU54YFwa4RpG5W5B5nWCeLnscJW/OZ5SFCpAleIKHMYQfWNQrQhfTG
+Z1l6RuZGRMdPWKQie9yrZpd37NRvP8K/Sy1u9zBuIHVPYgIPhuraBP6An0bcIf0
bwi7+YnOQq3tOYMzJ1tWttb4aEPKuYjJbJn/Chzdzqv6YCVZtMy9Rwi2AzYTkxw3
eWxeI9bp3hudtvGkY0fyeLFzRbbDCu12cHd1tF1oV+0thniIYsuoSDimk7xrTDrY
db8zh1FoZSxu1zVzTZs7/rpGyfPL1YUeEfr3RumasT5HCMQvnjgH0mNkvBEysuqE
nrXTdjPkJw6GFf3xSbh6o9iSOacyS6f4amCZsiPXu/ItGyGy/5UOkTkTsJ1GWLWa
9/6YddxNBx5h+QIj2bG2ek/lfLfBWQJ5zqcSPsJahxLlyKTaOEBRIJinJaBntlKw
JDGRZgmPmeg2EtGpLRTbaqnLpp3kCAQ2eSKNdaDR8RHGtMcSluIjsNwkTA3fu9n8
m4mKToMtnzADM3P5LfR3qqv0DKDIf/8ZPYpjkpTOzLtM6ockH8DLJJE/9ds1t73P
Rl+iDVSND01bCGeFNCMVSXPpdHlxYcKvGSfuFs8vocbvNyDvh7oOYBLvgVDoMeR9
aeTi2jUWNfvsyJ+rjFtod9uzf7qVxHiUeIrLtHiTjqvQtjfz2nLDOo3bunbgx8Xr
qPanbjPtNEMoPs4gKDT2AKmt58r9R0YsVFvyPcSJADCNjGIh/4cGfEzflMeQwJmz
a4OAeTL3IwBjzzQA8eN8vn3psQ3UhEJl7Xv1NLDRd2M7erfAjIEsG42YxKMG2yoR
z3TYkhaGo5H5pK3eZ8daGWY/xknmvHwls0spmY1dkSSQiG7WeWGRWCDWyqHzduYV
54f5KT9F0LifdAbUi4j4d7v9kQtOv9yZtRn8iWQyJdf6BVBilwCTn7Hv40B+jPof
z+wSyjGqogFu8wb2HexZltmisptLGn4q2vDCgO/pw2GxIEiK6kBx+CrWnLkQMhJA
Wl55BsmaLdOtznqN3FDQgQ67TF8+M7Xf1jSgcRBsNxlBaqFw30a8p5bvXZr3FxQw
CwpqJCOYttcF3evGl/ncxLtoWeZ468Q+bBboClOV1VqXgRdTZgTjl8ttA6pl39Su
SGmyeGqlo764azlKomLq/sebta6XTuJDjIOX07gLaylEbhAbqLPMMQ16zRk6xhba
QPRvd4wFwzjj2ElJQnzYsogOoLSVhKYgmI7a627+nOvpJwmvnCYVoOqqVUuw/2s3
E4Q3jX10ZyYNhYW4SnnIFUjd1knWK1cwfCQToAD8kHvfMQIDePYde99Tqu2+30VY
OHkjMboaKhdOOpafZwDvs9Ym5ylGDQzYiY31r1VAq/7Gxu9oAC+RiLfnyRXbVWJq
+Ghz8qI2Pcq/+KcGLrjDwUE7r03sZJHgvOAagkcKgDifoq7dHC3S3OIXKvup30wW
nSTyWwf1tddyqb5/nw28MR7/1zSNhawn7L45J84ZzAX7Sgcy/5EiazIyG8+kT0C+
9z1mD/ozzveUFv1tHPHwnafyh41WDeDoJyA0j8K8Whl4a17HHrID0iEKuQkLC51T
IYzIzPQ2XReR11/K8gbnyeXH3iCTatOMBQTflNzKpA6q0WDOM0/R7MYPvk0KpLrY
dlS+CmdJRjtrUn1gJLaHcUMC5TgKPiMvMXykabCVdL3ksTXrIjMLvDEKEf5mqNGI
Dpi9rtlIppGy5jZ2T7gAlA2hOd0CrUB9Z22bXKeVxSrwzjPoNV3VLkp2NRlbRD4H
xjx700rVeueda23qeLnKnBxCi+PfwUqZmulPLdakWDe3Us285O+w9wXv+WRXrYvQ
G7o73Y3/jFI4f4ZsCs+p1mzTW248ngAALaLQOI3lmpkta8j7yFE2Q7eVowrfh86y
jewgXxXzfB/eO+bHStQLHCv6NVrNzE0HRRawnVTSZbDk7vPbQYVvpVvye62BXXVp
UQCsw9evf3x3DvOD4FGaz4agpueH4UqxgaWFIgHGwPQuol2hWzlgROwiz2NeHx51
sXTGKvA2P0KhvoCRiTtoQlCiZFSnghjCqkOXptKdE3zqp6EU0qHaEQBsESWDCYuY
pPpG9NoqHYLvuMe9aubZwfvRlRwEHg5RWcIRQV8qsvDFhQ9RVT6RZ0hycJmtKpT3
x+RM1bWPB/VS/WUqkftZBebeCrRy72iNGQrxmM2+UCwqTEzecfKc45sbmcv0z/3R
QOb6NJ7Pi6Q6+mciRJqDnJscOuu8+/k1tiyKEvhrx+1hud83N75lims8+JUDL5Yf
vt3ZZRK6UO6LSer76+14BBtFQz+rIvYHZtzzH7ja3CmWYjbQSamWxus70ARB0rWP
B1BDDXPNZKxnzlN8AjxoXKwu0jOwLEYrXWT63mR5kL8fvCMKtkoGuj1EFR8OQgKB
Ng6jlgb9YoNlfHk1ac/hoi7MTt2FKz15HnssMSI6yj7tTJ5RKw5bY3+FR2cAsY+M
fPPEdHXDqa2lGyAP9m5f+Ml0AXT8nssIYrAkW2ji064SZXQHwJsYBJJuhO+PT4WG
jXvCY8YtKKDEGDdS62RE2i1CO1pNdgtRJRVCeHd0Z3Jz3us9MLKaI38YZm2AMXm0
rhXoXvtvacM6dZzgIfxBwqTCSEJbU3y5X35ZwUlR80ELGEwjUrmDQYM4pS7o0ymc
S4hhk/ajApWjbPjx2XcKTgPTNZBXam836t7JYd23w6vk8KIB9AuvFrMQeC20a6+E
cWtUxoho3rvk8018Li4UhraWxqarfCKziG0R6uPrVf07LDoPPRppEzjI1Qr9hXnU
iG+zKvXjfLip3CVErjDzoHGLcJWXmFPM8MbX0yi8Wx65bIXEJjTrBDnlm858l+Kv
JDA7HkK2hkmHb/Ja2E2FiEnYgbyzibG4jEeOeo1u4XCWS64ptR/CbFjbp4wQuIEo
QtoGfc8gshrR9PsZzDw3Px9VG2IGsNvl0a2/A1um6gls7KxcdGGc4J0pKRwkpaGU
4ZzdHXXDXAugG3h2jqBl3CQHzag7+ujMSRJ4dZs702yY8YKE6xhKclVUWPBI6LPc
HNy35+66oE+PN/RTxhGwFp1JRwRulVcnMFDexXyZYUO4w3bDS6NWsf+mxhua2R4C
DkNGwpSpv1l2BjE8EnZu+pUtvCo71tfRKTPSjsejYj60WVvs3Sjy0C8ikZvrg0S7
6tAAEbY0qAWWcQ5BRBC+dlD9i/DJa+DBF4Kd1t8uVGVFQwUM50scygWfCzF6Eh1J
Xo7CnamTzJdnpNVCXJsn/vUBNR6FACVi7iQLidk5F+0hDuODvMQWIQul/SUAbY8N
I6bte7XgKU7M9kejsHoYdQstxY1wi8duXQY3qfAKer9QDmB0jG0cDbtjgJWV3Bn3
XsLzbT6FpOTwQxyJOlL1e9YPdA4X6lw2K38ZJLFNLuB2SyWdjHx8XhXHpItuUz2Y
HT9xj1rDKTWhFzkAdeXYpBufbfCo2F5hDQC9t2kISvY=
`protect END_PROTECTED
