`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+YnIpBuomigPRIugRgXyiJgIj5EIWkp3EL3vfv5uz/VP/GsWPCti/ui3avbF30D
5XeaohswFjZeV6owy8mMaJCpMc0kuKarJbT30NIuWs38/BQBGcxSDAPnpFzhA7Gc
YxnVPftQCrM5U3/znK3t7ttqY0NOMoPfHAx7+qEFuST1GnVSkdJ/Elvr5RZsEPKw
DZW1OfJXaG2GBTLU5h3iODGk2ZIGh53x8SOPLlwnXuPeO8+A1hZOJmqKgNRfRwGo
p7fgHAi8pkG4kpAyx/+tXkdiqlQDacXOPzexJkeNhQ+QOqEieKFkwx+CwtVoJis1
VF5wKaVeQCLLsddScP3W8dnSGG3zFaayVZnpjKZKu4bCPw2DSfWMD3OhjFABbl5H
Pi72nV92ATvBuokMRHSX4gFVbu/L+And8Qn2OTbLpnzlPtstc/h0xdbAyzYC6C74
/wTrOZ9Eppx7eh7tQcS6WKBsfygKHOuq/rp1ztQwH1iROIyD3HSw6OqxAjg5EuUB
gPn/nVx1LIadBF/eUqfenm8HM6T7+3Yie4P7urDzwUcxEjWhOfEzsqemOi5Er/gD
sbN7XLDaF9ighFuZSeWG5Gdyismsn12PymaRRa4w/R2klFYYf3AHXks02Htyp0aQ
fOamJa5in1twwP3coVFYWPBbdW/tyhwvVDyC6XoDcWPFj2Akcq426QyosXk2oe7n
2i98lP58hX/s9uhRGpFhnvMmMURh1j8/ptWSz/NYJKQztlkon+k6Viphzkmkd61S
lJdYluqqtA5voRa4HTy4yfJSIcQo14fDb3n2khttYQNRUtCh8mtffZsY0fkoR2Bl
rveM4VXcnb5uUkqjkCBcNHSYl4yX6tq8F9EtX5COyAz3bCCv+cR+7pIOS51QWbOU
3FhCjKy6V7y1vG7DmK5pONeT0cVa+PeBaCFbf0ozrhe8YaNIqDA36HWIWhem3Tlu
5fS1A784Xp6Ap00C4+mLfEw7vI1OkZE2wzs9PW19fqSuiSmwgdz3jQ81RtXHlCjz
VUPBJ6BP26sWKyzCTG9DBBkn0Z4QwuGx7kbOTjLLdl+H0ugr1yDVELehexviTSA/
`protect END_PROTECTED
