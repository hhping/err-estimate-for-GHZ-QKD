`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWB4EIAMnBaig8VCGv0ezWQkE8KmLwyN5En18syAxShX7cb63i17/7Xl+uGCkmco
yXfCKC4UIEtf7EOxLEaerjS/40vtwCF4BwPbG/dufygi4sAst7w2fr9Rri9mfJaW
+wrvVAPW9jauOJQtFPb6d4nZib81hWWWtigJ9L9VoGYkyXJ5wVJY7tXtv5IfVjcB
FbN6df7/avLQPXnmvKVwtjlqcOo8sJdbkpDM8lNCnQdk3gpQL4/p4fVo1NlDLK8r
npPbCh+Qw7eZAqfSKIIVJCt+zMd/jn/t1XritO4Fftuoc6G6XS6ANbpflfZbBwdb
9YP4JztWL9AALiRiy6EPNrMsimc60+TBmdxEAet09aHN/6A3/5PiVUPkyyYgMPbV
nBkQ7oK5ZNTo9UdNIar5fvyaaFpo4VGJfORF1Wz1Pzg8TwY1nfXntWYn1r6lb3qZ
mjOuaC4pyu9JwPgHpdSLFMBJNvjfOMeLs1831E7vxmH9UtUophg/TiSNMdLTWjpW
6BqO6L4pKpPK7gn5nYGXIkb+z66mAHIZqNUMN6Wk8sZk7f+1jrsQG5XrMQM0yxnN
CZwRFM227UmRILUeMFDBD2ule2/PNd6gLC6qFHe0WKcfZ6lGhmsuO9/M6zlXafMV
CeiMMfChzVuSrmRhubFT0VZ6u6sKIehEdFxeOw1Eom6GrEK0tQ8/rb9tkaq8MKg8
oKEMmqpbRmzBBSLSqM0TLfefB5L89T8GNrieYqHIiz3cQpLUb8syGboEsPOhOpmZ
MoqGUJHd4UTjC/+XgtSxKdFE9rcubelQO7RjfEha+PcNScZ/r/D9jkjYD87UvnLO
fWVlmeFJlvytDFGQS+Lg2xiRLZsaNs3ymPYRkV8H0+qOQ9FZ4eG8vG0aRVS+Yamc
fqw3VxQ6kda8Y63TAXTRS6pZj6flshlTdJ+w4ztERYO6oHF1+txZ0OalsTXN72aL
7gKzyd6iPws6mVS3tZ2DnCvcSqBMFOHQunRNgCTZuyEdQUTJJmqewRo/dEIdOdvP
35BrvHxysXP87cTnXzqmoX7n6kIMiiMbsR6H0cwI1zasoAfma+b51MBv97VEB3vC
gmwstfT/rCylvaprNhTD9Smzmai3RpMVDlmwUNnCSH3b27gN9ncaeJiL72C+2hmG
5b7YuUQwfHnt1HJ0F8/D4ERgJhXs2U9ovdWCeAMTjT8C30TxhXD+D6qPSas2NJie
TFxteEYDdzKSlrQT2ezQhinXe8eJMUG/PZYfv7lkv/Volh1hq0SmgYmpjxgsbxWp
2LOYJwL/CNjXblarLGBAdkdozBaN+TKTloHLVIxx45jsweF3FTX54w81mpVszv/f
UnOECxiic4zXv3fiqFwF+aT/mdh8iSzPJS3iXvHIZs4qy1kwuHeVXTWlfIBkbEdm
A1ui/BUZxncpol+mBtf9cL84YPnSudhX0r7vAX3apo5oG/ysr53kSs3XVJ5MoZrB
iiDg4sMPp6CpZJb3IzTJ7xW0xU5YNalh/ZBKdp7ELEXd7Cz+H2ugbCpMwnllCXBn
aZ9d9scylpu6OI8C2CDF35Yr+QZE6vCoFZTdSaBP15k2jNbYgb01FXdtCVHfzDeK
kTz6KqLrqlvIcxRokvL803wuxq7uvBWfblhNyJczaX0kNu05qgwm3ZGVmgHq5/wW
GeHT//JD/8kXL47JRpqbaPPk5mpnLzTg8rhOraV+1bth5CI939O0fkyeru9t4uKc
b8wdhRMzSBneaip+6J4yRzNJE6XBojx5b5iSC6AFnJRtrxw1yDzToEaV9bsOXY/l
a38W7lZJs0bLDXz76m9t6iGSiCndtM7WYM1vDMy+1mlzLKQGGUdIeE9CbfTe+QuO
V6DUa4mavge18GZKXdB0HURRf9G57iiAPuhaop5JmvN081eh5C4Gbygl0tgTf9LX
/wjyLiyAeDoJt3CWuvgAs0QpjoSTN9zeDkE6H1i4taTXqnGbKLKR3qZ/NkxLecGT
MkbLuTXAjbhgbsrvGKW3XlV154Op0zupBG5iD9fWJQN9Wl67KWRJHAYgIrVkh5Nk
3HGPxHfAYDGW8HaViHEaYnKk3GUKxYYfcoNcKCO4kcDkBqlW4XlPNnwjKm43v8WH
PvOjp0A2LOHKwy1Z9KbCDOPfEYCxBPCpDkuBzLaUJTMrRQ0HAPWr/6FLS3XUK06Z
fpbdEswCkFImNsVaYmJ01mIlmn74iPh9MJxZac/NCqMK1cGXjdc71jxFQPZ/oRsm
VC/+lpE462qTtYfRaoPxRX+i7QqN82aCoNG6o+14yJTDrsMYN5cVJp6vCOI3WV8l
NfUHpqAiYyuaRKBrHUxqXb5YSY7KvwESq2SegMKM7Um5hY2224+S3UCT5CvdgMoH
yKuZGoZjdjMycZEU/DRPYlaGcRC7325Rcmo19h1gU7/46XG9w0M8ZSejZfLvszgb
enyQxfKBAeDSvmlvC9LlYQdkee2gqqtERUhJVQFg6tDkjOhNllGSw0xD8iw9iv5m
M4Ad5I/PGmp3ka8PV7F45fEG5bSPaFLGvmWvxcoLQ4+PVjbg2g9Rl426iiDrvuQX
3hcnYfgs3lcpqYo7jELVwQ9j/EPVJf69P3CC39Honf19o0+NRYHPw0p7RrFAKTlN
T2XL62U9NRfJWYnmhEQsHc/nppLIQBga/lQK+HSI3RW/d9+8KnAhX6IoEqq1e2Te
ikkjuS0YN/6z6bimksKFwsoS/f3MbkYVVvSj8ow6EfYh3JRvkGauHJ97xoThKQHF
kKhV9LScjDslR1NoDQUx2UeaXXYxZmTeHMHViR3MSxLcMWEAnYUWQXia5CG2sfL5
e90e9esy877Aeb00yY7OzJBiRivph7t9/ojipW0u9gm3Q4gHOn6A+MUjgx7edaxT
SSlLquXdaN4xlFNWqhh9DwmnRXOrFloGQ27pUUGcRGP8VGkncMfo0N9IZGDwwGM1
PWwRHoHI6Nf4f/II3gcHqw==
`protect END_PROTECTED
