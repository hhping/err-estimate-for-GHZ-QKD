`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5VLq9hPgkbBwD/rKkPRO5gOCG0sooZTt3gXZZps7mKfC59kRDu+zDBDJg3/baM2
ThzAeAPCKFU1fNcYsNkmsI6SsxTmxOlKEFRVeUSARXf6hUIT4HjX+8s92u72zliq
/iKl27wJDiRrft3EcBu6GDQfmQSrwM75/HCOVODBr9CF9IXD8knEWn3Dfdhxqpbn
OaFjV4lz/DQg0m6DE0mAqJIy8torEgZy37JDDeg0fr2M1g6v6PJKKOehITZHH2hO
mzPufr86VU21/ebgl9980nxV0iigNK1ziWkxZY2LjFBmnhVuXayd9BT18gcQ5Qnu
OtNkG1JFqX2gYquxlCN1T94aQbtLfj1CImKQimjsC+AGd/FM8Kq9DqNYvWsqQM3q
u/5wDy3ugjUdAqD/7OS3Z9Vv/1RkaXHWWJ7xHJIZYgEQtekjFBAlUOM7ZXHFAQH4
59oFwjJaj9DXEhZ3ciA+K6X4/BgId+WnMO3GBtORLPvMeprmFryoHY1/KlUSLQfE
zqjoEIbQwqKd749N8VcOzLua/+6w/xPYPr0UpBIdNt5xle7RfQjCf6EuUHpTuDIR
7zx19Qep8We0VOwiMeMCeFZNT2rUiO5brIbWxsW3ZDHNef8tajEGB3CDb/oOzW/f
wpn3UzJPsEM75UpT92m/897oPfQHQnmAMmpDKf6HveQzin4NGnXH9DcoU+z5xNSv
WDwjPMoRuk1bcxr+CxWsvhH3GRiIF8Zhq7SD/8A23A9xnrOhF6vGQEBBquJ9WjW+
dk9JmROizCROtLzU7RivrTPzzqSLBlLgcDVlneldHRa/nT9wOxoWrB6CYpWtPYVV
Tl+LKHv5R0wiY+QiESOY/dCJ4I7h3A++mJhWdN5yrKPW4wZOKAfWD/k3zOfd4rDL
+AinNuLOhZTrWB3Rxu9IaPrWuIHd6Ygc1cXLL23P7J7+RXlXaSpxz5aAUK5/lg1b
xyRGpLec2G1EIXrBJCjn697wvzwAni9W58scRGHL4EAdAQWzvZnHtcstb6rL0oFp
9vRfEeYBuQKbF3N+wylAHBE7ufEDvotj1Enqiq8/SCWATx+yKqonmn8/5M9GALRU
Yb9ceIo7eGVebrKLkLBYa2OhDlqvRijNnSUyeO4vkn3zc6IK+BuyKjxFfwntcMrY
nvoVMe7QkV1R0Hh0W1cXfx47GcHLQcYNw2zPBY+q5HD5m5wGg6KiyKf+U19SGfBH
OLPphtJUM2CEIpWnKBRUC4cKOFSalu0U8H8PyYLs8hdSW0+mwC4Z6Xxg3C2UtWMk
j7oRxHgX4OsELIIkzH7pF/t1loe3sR6h0y9kS89auSbI1rjT1KByCGfR/Gm0o1I1
bbUMfK8x7M5YYAXe0JuTfxsn8XAlwU8f71eRazyMUrZFgEiUDQYkK3YCFoO34uPN
7jr+TT6a4sCjrTPr1s1ycQccizBxYKkAuBT6xIvp0KEincmmdB8wWY36eHh3ssPH
hhgRxJwCa3E6wyTN+bn9P0csB3wD1elbzRHu+dMO3mPwBD6Ky22/DUBk3VTpDFlG
oiSzJz0oGkYukclKFofSF4uEYQGOxq8+bMbvn+9k2wHlOIkQfIV6Hf2lfTKHmWoy
d1YdNoLBaf9SyLDqvybGrP6vG7moUsVzkkXVtI2a6jBm82GlRWzsOUC4dGgjHL/8
N1pvweNqF42alDZurh5yp9D3+uGRFZ6D/w+oWMIfMK9cNTbrn5C+8Tu33BgmvlJ/
VcmSFhJvtioeY2bUr0dAeS6q3CK7deCaFk4Pe6nnLUU1RGQciGwtiDRtdaZP09Wn
Hf+3TFHKT57q985enzSawZ4iVT7gABluEGxLoS845NnT47qXidEtnvBKlyePkyb/
LzC0Zm2Oq1BllGKGj1ZgvAR442oCS0jfgtTJz7REa62tJvkPSjM1csEi5m5AR4q7
xuBf3rTH+KRwqhE2mFCX+XM4cosZSAB+ENtM/odtqyWjuGfr2fenHr0pdfnuU/fO
qkRKeoosEzcKwwShit7Keqxz/J7KQ28LkCHInxN1c+eZFYUJUj3bjbkf8UbT17c/
ispOW9rej3KQnKqkf0fj29pY5Vu5AWByPTcxV9FmrXWe6NAV2GEJycadl2x5rQqj
5L9krWJ3E3t4v0O4ORZwXmMEjNtGu424n+voR3q/nvGB4IxC0tPauXcfV2ges6ar
0YyjCdASwg9vOxHTzE1hEUwHMIue7k2zHQgYHjuR8FzUhCKnWeLxeQ3DVSsitc9p
8JCAQp76o94MYlOV4BqAj7ivUPt5mtIGhItC4n6T2t5k/J+WuL+WTmjvctIbNuGj
/eGwNUps0fQk1hFUfi4lqFFqek1iXV9Q/tbuR8BOraQkGQt5FM+K/0aXsIyHNi2p
5MeBQeuH436lvqYNSlQWjef+wNuLEENRKRiajx5K4KD1Y8qRcVnKs68tdsNYpVX/
7FjQv42kACEmX7RkIbyZQMWRKBXzv8mvOsggxA6+KloDQ6ATxe8XKZsOPDsEuzcO
6lNNixCoYOAj4VkENMcZ4A==
`protect END_PROTECTED
