`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l4x10jJKzhYQFSBpOAMzU+0Pr4uwBvKiVebTQh1+BQ/WeRuJb5pppiBgNc9SB3Pj
cY6GpK4yx9wJ4v4JjNDdECz4fIdMPpkUhl10dU1sLIk6QuRcFP48DpgwlcEDxu60
Zdz4eycL/mb64p2DfVO0w8t3m2WGzTSYRPXQlhW21ovvyDUwJXu9Of/XrICHRR3N
9+YOPkwFvRrCA4m/sx6FdSSy4LEMR0HTsNZv4IgymvFoTsE4PcbGOwoTFFo/Wsji
Q1cP0hk+3twnOYmm7lBWqEkW+RUrc3OJTM+uH/GnvL987OBGbx310Y++itUIBD/9
8phwWaDr24HXQVY4ICaybFXKBgmRoQj0uHpzkm/IOmjV9OqvNO7bA15Q+W69pfAs
FRGNDllT8USM1FxwtOa3aSQ7EdXPrq4iARVbtX2HIhTRewI47DVCshbp5O7N8JlX
Ji8rkIxXjFwa0wd1iV8KaybWraq5YZSGMkvrzAvLpfy48l0VNdBmhV0qsICZeoqU
lihcjcuuF4e35D1MEXO0Y6zcPbQBhPXxf1nw3BzfP1crJ1s1eOgqUQMTYfPqPeY7
emC3YqhaI58JbtyLqCKUm15FRfVGjI1xZj/IuGrtyGc=
`protect END_PROTECTED
