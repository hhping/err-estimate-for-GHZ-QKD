`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEQ+i8fINpmqSLPzhGz0myrKToNW3SbR+2mwedh1N/B8GBigZz5QS3tMmjVrSNNg
mkXYZNekQp3sOBxsnPMoT+OtqCxLPvrrVqIq45os0PGAHGINUDi5fBiWlRyzjUua
G3snLvyKIZdE1dg4HVRHlxk1WdY34YSS8FBXeHUuMxAzpvgPHv5VEhmajX5mXjby
iJd8naAxMYXsKZSWYar9Lkfn+qRrzaNP9Dg54KxufWRVWTEc6+/VbrD+bTPYY9bI
evZ39xjZz7l2GHHyMDpvtKk8ebsrOcZ8w17/z+UyUqeqJNqNDpAwmrMtW1R1lIMh
74ZRg8/MBrsFaW0CF1E7IM+ZZyt3vfXrOQbnXEV3c+DJtR9EsglhslMhRqm8Usab
AeakIeAeG2ogQKGcWL0QUjt8inWP80BUwljbr1ROHAsMMy33Jyz4nulLJRdm/w/J
jG1v+MeOO0dsQeIXMIP6+F/qByN126+ZJFUBnKR9cnPGYLfMTX2uRmu+CfdQqnmh
KgdvMyM+JYHEGDWKgh7xGIvbD4aPfETYiTbxbI0xmnWNEt7p0k5HYYTeLAROj/Cg
Thkdjsx2+yXL481TYKwuF+06tS3zq6+FFUZxnSCHWEDy6BkO+Ji7AvzJONIjep4k
VgQiLSZsN6KxTVgir2aPy317pBiKuOkMUPy4o7w6wRLpRQrxWIGM1P+Nm9rmPvfh
DP1NCPH9NOeSNk7dkFLz1eSEMWEVUlmmmZZmH9g33n8TPlfi0rMyDWWXiWz1wazp
Bb2MPCjP5NNXgE0J6Nu91u/ihXhaIk4nSbapqI/1tr/ZBRVFJhx6MA1Tg6MbIWGm
GZXjI6BhTV0qLqBDonJuUTTP/gBBxFulZVceLUWxnflx1uDiY49E3DOSj6I4KV2/
0OmvvxbPK4l586vFFLtpVTtsVZD8Z/NjKqi/P63ytFKXC5g4C9giqQKcHwIp3fHX
ViGDjuJKck3w7+XJkU9xiVKfoTvsz1pWzXyI3i4ysfEyRRk/t05u5tJdOQucxGIn
O/NDYrZwQxnsfW8sTRQo4pd4I+/dBGUHIOxV3VSwiZJJaRrjR7XgHd0FFHXu4I1G
sALUvz923oNKUMGzc1pX/w1/ZRZp48AgDOQciTfGHWioxU/9SYV/hD4OY//Wzr0r
yZGiY7jHXkhp/bgn+MwNcw7xDxFA3EwBc5KEIrRnLBY86hlMsSPyt9DlDzWVYVwp
MEqmzOxRr/Xadv23lGgMJqE1uwdUI9dBCkF2g4np4xrvjT6vCSjGpLdywlc6ZSbe
9Kn0zSUwUqQDCtcO07Ek780dVxa1DwJtS6VGUkUqKTaM5Vr/a/JzN27pg+MvV4SV
BRTEaXsLzNLcLxrP6kSKAc5y5DgnCVfH9PmU3sYSN/zSpISRQE+555hFSilplEDO
yrbwgtxeaZJh9Hi+nP2fprcXs/LGAkc8hQ1oOGnOwJa5yYRnUkNBMPd55XSPGLDz
MNh5LTrpKINRzIAdhdXeLDWik8Lr0nNcxIkaKQNXx4okdL2TNqT2QCHCvBr8J548
hZORATRK02/C/Ulo/MyyGDC+E4X4xJW8T235fMAVEsoXBCpuQaphl6yBzbobRF6s
4+LXcd1V7BYVi4Xde0hIWzlHUaOEA5bqTIaOgnMlZlvStykXoIsCm5MrxtB02SYK
4PyMtBPUC3cSwYOCMj7vBsk/qxAvRXsMwG+PLE/LBpLpZO24XNcLqQb3Y8vQdZfs
V5nqCiKbWBr0kwODthwfb19/J8Y5+NUdjVzvV4ncbA1daGJLxguOjQqUbjjRQqVe
KokIEsF4pqQCZcmYk4cfSKylKWaHgS5lpXTaxqykE7U/jOo5LzrPo9xUFzV3sJyq
AsalXksOhzKOJB491/qK/dFfCx6R5/K6EixvuVyV9JrKYHNrRK8DK5dIjr2b0dLz
HWtGtb8LwBubKPGIO5hCmv6qQQzDS4na50/Y/xyMyg2P3AmPjDiZjpTcgjAsXiEP
TiU9RZM/sabC+ofScWEb9VfxDr5shzO2tJEBi4K5HuRuy/UIY6Ciyzv8sUdwH1bK
DHEI2uxVbSEId9FSxiIdewqYbR26MEZhjQzFsq6H9IERU1uVOOUFRG41+xun/8VY
zfhFLTdx2azu5gsmif/00DjrmaPMyikLNSkhkv34QnpyhTfGCZbBblIP6ZBt6SnJ
3wh1ACAjUHHdd+M4+M6cYR7N8qZ/i4yVlZD+daMDPpp7CPlHVPwvTMALCBu/KxbH
lcqMVFhbYLm0KMSEAXon15W/Semhz0Vu8D1in6HF/9PDWixeR/G1G+ukuVunbySq
`protect END_PROTECTED
