`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpRQ7dYw9xtbVXAUb+1r0u+Iudhs7xKvI/JeoAxVf2OC6X/4eEb0T78XF9BbY26o
8e6oE2EFiw/lsLt0lLvF6FKRhJxT/oUOxXkBCILne164Ek82v4HN6aiGveilMU81
AnyVejUOtyLSMdXP3OS4hKBOMQQ95+p2YWa8BQd2/32K531sGWXYU1yRXfNfFjmg
Az38ycQryfgcOP1+y+A632NbHx0T/tzXVwODhitrVr56NU5G6eYEXasrSO3o7jJ6
7nN6OQPVkDxTW3B4BXePOvM6ZNRp6cnX8we7YyGebFgl3Wsm4jz+WgUjR/W9bd04
YydKrULPhUFRbabkXImbL6qgoy4jtDr7f9GQlelbcUrR1zNCWoABUrA8Gmj6TZvh
+TRFsnw4avJyIKk98fgpHl57ZawO4VlIPmaIcRC0TApvNhPKJXspjnqM5im1mPpL
L5RKYRuCEP6XthSTSyZgf5Ydq+OuZVrqY2ay5GjuE7ICMFnBCIekZfz3P1pmomIL
yc+swx5JMnlJJuoYjK6sCc1ObT3UxjF+zkFjK5rmsURpX1Eyr8iBODwVSlmuuX4G
k7OovS0gykxNXX5wQUQkht/a8qJk0EKmNK3zKYs9ik18z9IOvH4stxRj38Ui0vYp
TxosxECuANqx4nORmWWUxndl813XtuoKbln39VBlrgeoLXLLDirOc3Cj/1sVaCyy
aFDij/TzA1Ni91QUmFQBC/eyp98eiW3/8GTtWVM8uhc=
`protect END_PROTECTED
