`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vXXmgKvGSNaCMO0u/cwKBVHtIiYXVmthmV97n3tNkoUwtszaxDEOttnqgYCpFyG
GFrDT0cjl6Ulwl4B48nSruvuMvhbKLn546yOF9XyP/ZGiVgwcud/LSJUgVwIqiEz
KRc+X/beANK7cBLkQFMpdQuAhJNIMzg3f1nZlhSADxuipIYUr56i8OkR+C8kylGX
Ty+3lKhDZwowhbGuK/rmiTk2OucZw19t9/MXSvkRCWYvAzgeKsJ4Ca/GLZ6Xl7JG
Umc70IYLoH1tRwfWEj29l0eF6UPIipFvs/TKfhWwDtZoZ/IbtWZ/33xPNwIu5JUw
B31+TVuxvtI/5nPQWNwTrm4+LgC/x1xw/ARWqCtW1bsKIT28QrJUxABlTwPuuYqR
XhHGvd+iWoK0O//F4HaGId83brWpss/Q8ep55JAPMvraSEjU1o5mqCPxNNuBQjfz
7grjjQWnljWQH7nb3Dm8ragxONgbpKgLrrwT/WPj2R4cYU/XpjYmmPmk4jDD83ex
R7Ap1tKws7VHDXHoctD8wauPaG7/EabVaMiafFN9jrgwqH/PZp15APeI7GN7t+BA
gakwivMgAkzkTJY3lw3yk5AWGOwKxlcZzt581ksr84Ko7fmHk4pDNwsApmqH/1Fj
Yoe0ocqLOE4la2Sbx1H7dyiFNXM+nwUJ5PtZRpwtBzim91WHnr035okd7zcziUsL
cArY17Kbty+2oPEQwQwtC1a/YDbpe6qOc9NhEDt5+pJ2XIhcRRZb/H9b35SbEgMm
D5zZMK1dZBU6NnPYAtl4TJ3EV+seUblTouXpdnOfNfHF+ngY1g/TDkrMX6JyuFOr
alo/I0GhKKK79BDVMowhAjSANPsDPUhDBg9UD6OdH6Dao2a/zksoEsXXxg3conbq
Rtj2RunZXJdjeVFQ9JemJjrzIWSjlNnQ0SOI2fAYP6aIf7wSRC2IjKIYXkEIA3X8
1T2Mp4xwEMYw0/ek8IztR155rRl/B6EgNkkpmqSe9Mr52M/qcu6pEi30tFI4qu+K
pL+zgCjQAo4t8w2zAZk6jE34ZY/o/1Xp9lLyqD38ouSanjXlzCzj0AxbwkNtfOXo
YcqGeaKCQ1kmk0mRS1dbd3bWrYgabPB+xByPX8yBiSob50YXgqOhw0JsnQhTTU/e
ifa7mYaSSbfr7ueuY0e7bHo9LeTVeBAm34p3vUIMtRsssoHLakhjdsxhSD75NhKR
EazybMj8wX0Z3oq1jlF/DH6te5Y0BLkNt++12bAHMyeMQS0WMCERCxbwAyIV9N2y
3KVrpe81wlSdOxTgUSea9vVeoKgC7fYQxOz4mA2grUAzfgvU8EM5buYtS9C44/xe
XkeF8g4H1njjBPb/uqUxF+AhNC+XWKWmXUbk184MvANV3EE+BBU1LrHcAuEpufYf
9b0mYd7GtxsVSfd19cyWDhzcFR8htOFmlE6bBXOotHHUMWyvWHG+o7BsQKMwoQKC
NNpmMzWy0CisRLGBsQOBd4pdsPCAViNW1WayUPNwT2NWkEJ6yzYUJNZGy8oRRJrM
/2n8w7NgKoB23haJy6xvCY94AyLQa2f6HYbDLPDLcMOxBqPLul39ibPl8vO2LlvE
6ZuQgXuZu/P1sa/qDNBZxPd22AWLD4jEa9D+6BiRoFeD0sx1VwEpZxB4uaqAokrO
LgaM8ZhNaNxLXwPJFEMMdMZdVXVGvbdarKwfPuDPdiP3wHOF0wLsPjBmPXQlwHVS
CrhGp1ZVTTrSdMrHQnWSLmtc3QMFkY2s/rnM8p+quSgx1s+HCNF27yU/thpxkeMh
kXOnxFo2zikOCMM+TUNJiKXYIgfZTaTjFVMc587bd76XRB9jcEGK/dPa8U9tAFpE
Hi2ENA70mHwVZFwomjWCzL3461SCVLrTXQayT111G+khmy7bTQNiAE3TyglWo03Y
FdeCaLTzTyVvirVcgIR3rVZ0cQTJc/+vN3aPqMLdQGvBmubehs4r8O3OxTLrvcvg
BGp3vonyLjPNs0Jgk3pwDBOSe4JS+8IHyi/FPRb3vpSujXaGfVD7qf8KRJGSk/TG
uRRCi2dQGJTh6Vh5gT4WS0m2xCI2OQ7nbfPfGXhmXshX/3yP2Vw23C3c9E1AUF7g
LGE0dmBgOm6tLrZSGAyqd8ajkrPjMOnIQjRb0tarfGXPnHL25cvS3RzlsCqQLiEl
GavYQaoRoZ1zMOQ4U07n+WuiJjUSrSEAuU3TRiruUxuBpyAOgTOxf6mQyusgEPtw
65Ajl9U7lSbdIFRDc5kXJe41CKhSjRRHS3g3XuGaDbf1e50KcNtJYVYyQ6Hzv5B9
7MXMXKi11HqbrH05S2msnPe+pSrBXkQYMzWbZnXW5VGC2K0gIwgO42TpUHFTILfB
T/ZHuGNUiyQqon+IVt8Vz/TWQPsXOOqk9TV9daZQHo6IfJqzNkCQrGmNo6XjnHsx
vzEmcnpklz+b8Q9WzEWtJv69iNSOWQ5yiz4CLVupgEod3cLQgQtEC0NJzGL38J0B
qRxTNq2lJ0MsGPOBMH7QsUJT22vV4oucfE6iVPTlKC6S99PhEBvZ5t1PHbS/gDCK
9peS5Y17s402pA8jhWQPA0X//9Df0JhQmkx2zn6pxOSolCh4I0Lg+NUKRHkalX6g
hpEJCfrfPJs409uF+zEcszXJEq59UfXCrYwfwHl2N7CV4pdni+Kch2zmVIS0j3nR
yckZUJp92IVD3hRSdu/Us+zYqphEWsqtYnPVOvvHllkzB6etBH2FM1TIV6vez3tK
OLBOBNh+hEzkGh/yjo1/ynxxU+TX76Jpafg4DRzK+TThu3bWZ4YBPxcIvxK+mD4n
tRwmxDiDY8WfWWf+H+a/oNJniIlJC5zHJgiaK/udcKHtSxkk1m8UOLcj4iRDRoHe
U7UUGoY+gnjIupgTb2y9vlUzUkCb54FZRQEAGGbrZ9RyrNwkgLqK1fWfVDV5zRa0
h8NHw6od4CnE3D7vjcQEQIvuF1zsWJ6DFTSSfzM/6j2jW69djlbOQ4FHgOaDR2P6
yMe2oC2j2I6JHRl9fG+zEMw3yYpsvUnq4VKWqcVUXJYV37C56soPniL4Lz3NzLHZ
QwAUonO79GnO/WlEI7gQycnjJ3DnD6NbR/CRtyvAg11Kizw8RAlyzf4v+Gp7++pc
TuNbDcMEbckvmmoHGYg/fT+f0jymlBIrcvO2nAU/DujDSckZlGjdQ2tIertxXiwT
yxz0AGgMLaBGb3a7cgh83mdbROJD/qDwfxitQdWpSgTsSZodVz5A4FuOV2iwkZjc
Yy44pE3qk9+ymsCq+c2EX+Qzfmu4tP5pbyNs1w6eyReNm/mm4QooukwAw2KO9dz+
icDzpugq3QUjqso9sm8utK++8WjQrWT3zrU/trngz/1DpeupIpp9/XJx1PDxneki
oAb4vpvP3loPGzTLNMKYAsTmohGSfdMTCjv+XRHXY/k7zlPBhF+nFgGJEriBF21g
eqSJmnf0yB4fhX9S+qSJTPEex8R2+0GmWZM2oakyitiCZgsbpHpUPXIrKLhLWFuh
cAU2Y2BAa6ypuNjm7qoPmv+ZzX8oxCXkINSv/KqOVss51c4yjKss1oTEg8VbmTxR
+yboQmnpfCS7LCB/1XBFOW47pAK4Ys7QY0NT/MDwb8jCNdZClUMrdQjp0pNrIZXT
cMpBZXyMb5YbhwPPhWF+wybsPJwsGDkEonMuBK9nrjgYRcN3zPXIxK95Pdfob44L
h+b1GGYWOOQFUB1PwQHQbX1yUPH7Epdb0qXJCsfexR5CUqLtGSwsMftxqwYN2GJZ
zhVVwvIwPsuUsjopbg8+BxorAyRfdzDTB6U6JHUoRLPKqGQigZ8cHzQj3wvE5tTw
vWWhUFt9Ab6QPvbMRIHhyg==
`protect END_PROTECTED
