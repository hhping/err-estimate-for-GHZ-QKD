`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+v8smByho160iLbBEGHlVpdHvZG/kIjhjbNavSm7g4sEjH3e8yTXNcsY5AfgqD4l
103PvjzHllYdkL1lqE4077VEgoKYOHzyxny7n6BWUl9arE7M73HYQoyhEdkOe2SJ
iY38QkuL510S2D+jU3MR97Whkw4nqm5XGzB8zktI9zcH8GQyfIpiyrjOljI6bsx0
YDUmTgOkOCO0HP+BoH/dPCUDQzEmsSVi/LjEFPMEKus7i80OMp06o1sHLVjRa0Ct
fanpgFLBvmWBjFLtL1+okKnNROquC5FGtty/Fpurg/hCj8c1S3epgXfoOtSUOL8n
GKi2LeBdUrbofhDAVJ7PfvPArc32o+uGaFZNhn2sLeKUdL/V0mGn36Y3UvVBn7ob
kh9dz1g6hcCJsAQxYp38aIUMEFgb6guoV+NHiSKEFRJyWM/THZKxeCcIcYUf65tn
ZMhxfTxuyk4YDmd6GpUjXTZjzzqZv8eng7iybX+tF0BaE4KqdyyHVfaS9hnMGL7T
BaPZ52dHodhrMluQoDGppjum/sqZmfYUO/2mzhixjFa9rLG4zvu1ZXecNUtVeT3R
lRZBLWgSInGloUGbv3A6qoNa/4F5oVCNT73wFXlO7tb7vO7pCun+qKpo8ANLbfW+
gbVzCGHOkZgnyOnJcSvMnj0yWl7PfDjKXh1bG4BjO+DbTtO5rV5lMGhzFD20+xdf
goVJndsauEWIrJS3zhvsa+xDRcMzOMcELzAbIknaLerg1e3z+nkgqVdZ5pngjODz
toSbQR+cKo8iis5yEcE4QKl5dPc6x6gm6I9KUj5loHUzdkVPj/NCoUuwikiUSM2q
5F5eH9AfgQRcIIZBtPRL0bhJDXpJNAW5aEu2qHfx+Uwe5cIKgScfpqG+WEhRqbhr
cucWu7trPfDrwmZaJWmqowhHXnEjl2EXPYmILZRECzORrWzYOv4X4MSHSNmXr/+9
05PyLoMW4b17AM9RJgU1l3XzaFtJYG+rv//hCyl2amc=
`protect END_PROTECTED
