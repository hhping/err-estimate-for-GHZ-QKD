`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9E0xSyl8QYZJymXWfv64lZhwZzblBSXi07GUymPwYNf8FwvIBBe3qA8RdR+4KgAP
ghc4aNSFSjxeVJdkxerWo0yWBBeXdSD0YsauRXPdqlHhx89/kz3kxnsCYx+HhfC0
p6fNBpabzU+MxM+NRWuUYGwxAs5aF9EQ60q2F1ZqX4qC0Wf/7Z8nPl+TBgyQ7OHi
BHHT/h403rIM0gc1vyVDbFydu5s8ikwQBMkz+YyTmSMoVUpoCnJBMGLhV1restYI
77x88GkBtVB7nqgjlRT7FCeQCPfobRWryYsw7ekQRjJ9Whjjp2GCbPejhbpUAaVD
Vern+L11m/wf9u5vNP1znpLzK9NGUKnGfv7hBeqrhWauvxsIM8TOHbgeoIMgFVg9
M8hsRDRclOa4KsHaA4LR28T6WLyYxO1TewmwTzaAjJW5e+xgN0aF75Vd3tWSb/Ll
Q2gREVFTH3OZqWiy5HoakPZmvGT96RRIce7ACsFhmb6yhZq1154mCU7ivTuKKS9u
RIx5CxJYioER7HU0aUvutJs5n7qbGLaNAe+1VnetWcFzMMNLs9Y/cPk68v5EVhFV
nPSyhr5SBCEnEj4CkAZh8neThEdcygXFztS0fKw7qJ4QgEEMYSTlqeFmcbsmOI2p
71NXgNVjsX7/9d7zKZkUYjgIKnHbe6azC7U04XGgqA/TxV26hxyz6aCNE+G3QC3F
8o1Rz6IkhMU+mA7rl7EyWoDOgkCBO5g1Y1X3So327fE/YoUTo0HNZwm/RvIxkgd8
Uj7//V4sY4y99CPHYQ8+5AfICXC92YAdPejNgudNOCrCugYWZ/m8JONJ5yWIbHW6
DnSNS6EQCr390JhfFEpKQ2pLM/XDYuxk9okBBmAU7OCwUQcwMNVM9VOXDI/BsxL2
`protect END_PROTECTED
