`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Rb98y1TighsjP4GufyMhG18plEcoGVjADkwg8xS0SsiCFX1+HK88qqNaUG8Xiw7
heI0zkJHw7ONpovGeeKHqFY91YFtOIhOlPc0ktwoblEfpmPfURpsNOQk7ijG3kEU
MwcnhCnSiw4n+sWE936wxs9/CUXtB487QAzC/cxTvj4Mw3JhHb9Y6BGPmyGi8Xhy
PrDPz079I+LwaqbtkUGGbDpsVEY+lD93jqkvY2JVcB/Ol9vwm3WYH6h8hcoobiqt
cE3HdQf4/1EASAGhXK1beP8jRw/FNz31MIqDT+3p71uYUe9bMTRHHiTCPHepQJWB
S7/dnqrvi19E2pXHCrPrxc7h4lb7wVdOXabZ0uRvvrcIBPVWLyugxnPNqTMYkDuy
1GMDQjUCQR/MhCIHIGRkzUlz9uxwx2HE7EZKi/4c8U75aUew8ja/hou7iiSLeo42
5A86wZib6Lek7JD9KnB3eRagF1z+dtTkAf0tb8ssN38OcovqcolTiROmK7cUQALj
B+zNPGCan8Jynqoi/GNNHeTEOylKMiwpfHzjqwIipqWDOJkCsWB0fMXJ8wlwlWNG
GtsFBB7kS3VGcutbFcgN3NCi2GbvnDW+1Sxxjf0hAYM4emrYRtKdU7MaGFRWQt9+
kaxAhXbiGH8OF685wwyK8UJt535ma93mXTwFzH8tLfdYeA/h0mkV+kvsESxhTWWj
7Xy4dwbIr6YqCx+VIKPEBMIXZiwia39FkzDfjmnhAoaRTTtsXVmTK43OmZpAv+IR
64UTi43dYKkNAVGPHip/JhC6N+3cZKR65hXmxq6nd9ZhxHlpf8RASwcMXhAbd+iF
OwC8onaHqM7wvtWe90HKNziYLC6RmyMIAE41eN/gPbFxHOfCHaJN7Ln6aCRoAkO8
mC1Vayn4MRvt2bKq1BjuTUCBXMCq9vkxwIE00Qhv+xL2JJKxPAPKay0grOgTAb05
vEM1e3Kt7U4Zz9dQTDJRmUW259avIPBEZZ6ouwYdf+Uy6/o7bTlMLj9AWnX4Bwaq
k5B8hLE92b4FMlfOCkBXG/QulPArY9bqgeZf2JbasW2MoCO+hg6KY32XrF7KfS9f
kVt6dcigjikpjnpX+J52gjzlDIQjTMnNkTDkAUEYJWbnY3bmBAzioumnFzGfdlW7
kK6TUW2arEeexn+3bpyF4v2WLNzc6p8PGMJ7N7iCLmsLMmGsKmu+t5x2K7IK2xiV
4leTN31tAeZ7XhZdLD3Z7GtzTJFg/lF4XDvFUuRgkECRBW5ir7KBYN0Ybs/FJgvO
7TY/MJ1VaGNMP3nCCXEL8Jq4yFgyulsLlZUfDlxHnx0HG5r45oSrq1dxDZ4IyD7c
8ZRgvO3taxdG1DEaq7np4JPayKT9hdXnBYQu8tE5z4CPqGEcYyWhvyNR8QJnvORr
D1KHFts3WOQtJ5FNyvscV0TcJYRNyGIjYilVw5EJWa9sr2patrzy+h3zyDdiXB0k
sMxZOaHP0cHH6986Ej4MViZPYRFhjGzvBDzDBw8mk3Ee+6LuBf9Eb3sDEfTpTDA3
DyO4N9iqK4a85sA1e+EJ1R9KyZIIaLWm0gXMGYqz6xZs3C93Cn1tq3bFaeQvzTYR
NztU7DR0HCPiQehsc8ki/eErldFG0T2qOnj5bOveDZRJtZi2v27WI4vDIC2XcZ7d
p9VR+fnfr1SpdSH/z7CBfFlmvKe1zkZYRaPXAKNxjmnLl1fjXcLMs7JapJi9u4BT
xLxnzHexYubvCbYV4q1MEY11Xscz1igXLG+4PtNPYGj+rtXY8J5uiwqmthl69e+7
s5KTqkAbteEBPmFomPnIcwLsCfzr3/Zwhf8m26nlteY35FmhMFibRbH9a+1JIdA5
CI1iN1GvRc5ML48gvnOxWVVrguhhYYG+vBfhY5UFghL9qYCB/P2rGiV4CNMZ0r3u
2fAbwO+2UOcghd8jeGxwKdIU0IMKWv1ZZJitA7/FXabcFgDRO3GI6csedBwBZ58F
lbqwOrWXZrsnsPUYTlszBViwOK5WtX74BjO4QxMvZ15mo5oNjig1VKJpcAK1YxnA
0mR2xUOic07BdBsEUrTbt/Jx5tuz9tTFRXk25WeC2WU0Jef6LUN5w2KAUw+AJgbD
ovT1XCrR5kX9gxQO3QT8un1M+MsVa7oGvsr4Av0qHew=
`protect END_PROTECTED
