`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ox4hmzxjOweY4nuPXacvIo5g4XcJXYuJFkKvKHR+abJ4WHF74mJgeofyIsGc3rIe
l35p5+E3n9sOCkd4b5ekFxo4Sfu9SBcaE9LCNQdJiaMGjjmb2ZZKIrf65uOdLzID
tXfls1c6yb9H8lAiuP6ouAc/arzUFyB21La3k+aRA3pEAZBF/nLXqTmMMdVYPs25
qke6B9IjC3WIid79X89C53GyUobN0i3NjWAbxkp9qCISU33JjIz3yeemmh2tMysC
WdCoTFp4bp0wcZyjkMTN0n+rseHt0+29TTS0FUa7jOEwNGwOCPkyz+DUkbcTr6Jy
6NEiOkjzKr0hSPxKb19DqUsAmdYVRH2wac25tSplYzYvQkonH7cwrhXp7JsTc2B2
yki5BgRaENV4rBYc0jW7WnYmNlgUaBIF7zFoEy6+3ZUT+9+o/Mcjn6EW6J0d7ZDY
Q8FNgyec2d/lkJpPzeftnjpMpLPFu0Xr6qrmcDV5GNVIyg+ji/1gEjK67MkOsZih
mElyWD6vUll3ZylI0cR3qgl9zpzjTYslX54Mpa8dfhHPqQv7SmI61ZoSXdn0DgMr
5xkylKYgSsjwX8oQReuTf9fX+svUgpcj2LN048ItV/73zHRQPM6wjmejwvJYTOyA
zarL9t7ZJjSvm4rU+pJFQF0OQSgvv3HF9r/13Il66/Ozd1hOnxuekvKfxRPpmGhK
k8OUfuW8bOSpzSTjdTsXC/h6FcG1zanMAYWE3PzkwDBMaUMiBYa45oM3Y8722bCv
CvqdhtNeMTOhFh72r7LK9M+9IWdU+XVznmW3Nd6tMX/qjWe4/rCgXpqVVNGGHF7A
iZNcghQzG5iPPCJsmXYHVfVDPnNzb2IM4DnJU+thcwo+UQMvArArLGzkw3kwKaQA
lkucqtEOdmf/v3U9wHNbC163ZUXCvlws6qoNbEftymyg9Z3+AxGx3LzWIRa7u0Xm
Ygqg+fg8dIt8joP086oCKZhsqLssc1Q9O22AwjMtp8Bc+EOd23adkPcAYQvMHgfy
UCXYWq/EHJwfNkHxkQx4sUoPzasmrSxXXCVtvj3WnSwFcGfuaFPuoZek+kItXq+e
iDjvL+PEqFYhraKJomgHKrTG2XpIvo5Hgu1vUZ9EYTQ8CP/+nPKXYhC4Hfn0c1sc
d3+5u6xRbOhLrxg8hFQIhdJejXQ/xOhZnc4qCu0orz5xTey1pu4Csf6cTtKdd4al
Cwc9+EKxi2o3MAavYwaTuYW0RaK7tnVaFzYuEC2m6+lo5H7GJSIi6SO8F0MGFt2b
g0aMQ6xfPxic7eHWN8okFZkWs3gU0HzjcQJUZ/F+NKhx9K9ANTN/Z5jcROdXnNsk
d5o/qZ4v3vONg2voh96+UBhFYSaXgA5FUD+xkaf3CCfuBeQUdr24nkMok0tP+Nhb
0vrOp3IsYfe/g7IyHbyzy5WeXc6z2Uq9KLLHw515mLRGvqDeEaGIAzBhrkD735Ea
aRxtbrzliV+hSGHx4vgUpO8MSXAP5DkCM1quVH5/yrxqJJC4jWe+QkYN8ohJwfJn
1b261KjMK2c8dBVfRW51kToS0XeZvCjI2X/7+YWkK3975m1cpYEpwpF8rcMkz/X4
9rwdvlY3t/f2TYthb9Fq9+s1QyQk3adfXIO9b9EzWIYqIOvdV9IVLYtCSekRR4wE
VlKF2xczBIuVIHOdXXu3smvjsSrb16PvEI5S6x8G0G6FGTPHuSPScG2W0zQPSVfr
OrKPAF4GWWbN4Vl9Jn0cn760vAFWkF7BWRyLzPeNibP92ULjTKg535EHv6ySDHTU
5qNa1S0eoYPwPho3Nu3Hc2+hhsfewgZadJ0yKL1uleNO6IRWfCM71UqYZC3/XKSM
TuLH9g1Cmb27DUn3GpHxjyDPxPo+9JPwjz93bRBDYEk9yj/N/espnMQ81sx5a2vX
zsY3jb2f2qrbHn+ggjxDgaVitI1ePNV113aErXUQWU8xXyiXf9/pDDbpcBbyGaIO
mbF9dcIkVn0W1l+qMvoSy+2o191+wD7dlt/witiQP7wkFPXqN4QS/fgLqWpXaMe3
0fkfQsBaYOLrTMTITIhzZST9ocOCN2NzO16R0fKT/5bBMBqFaai9gIJuJn2G/6I+
QdfBt0vMi/LcIjFPbAQsJb1SAKWOZS9VCe4QO1rBDiz1pMu5N33JGgYDIG0YNTkx
4QoR3rM/XcWZl9U5QuhUAxRdhDfCPJh9xVwZFnDQZPI2yGDATessTMLfIMMUF58s
XeNxA5m8ayyYAKBYrIhOcs3bkeUxM94HuzVZpsPDuJPIh4x1tdk71Sbm5qliExF8
6vPzU2W2kH3w5lpZGhT+VTtD0xCmNDwap2SU2pHuCpmiM+AcnQUtUflLp1ODN4rs
E6X0hepB13w8f2/MM8pkdCe44TBhSJY4wie2bdYzJ5RBVVonObvYy4z10EDQ2U28
lPOoG6nFgtewit1b0S6i+M15B+sfPtjmgT55Rq6Yyc0FX0atRtMmBkzFtg020SKF
6MXipo0R7vA60S87eY+Dg+nkgIzo04tY6s5gCTZOiYDssf75pnJIwr5EzFkbR4Ij
GcZP9i5W16jM0qqv6WqnVe/QGjr/hrh6MiD99ZAJlm1PwYIvzjeWWDy30xmXsUCv
1vHSpyGrXny+GxBkbjvEn4iotGXW6cAWIqW8x3R0KcT3IyzjfmxaGIjMxvVwyr8z
PjYTwxEEUGXLqiO0U3Jh9qkUUzwHCo59USUY8WI6hhPTzX5QePxdi+x5CfUAtCJx
EcBd2soP5CVKEQM/r4G3a7z0MgLV2FVgvb7IuqQrL0PgcRngdx8T4P2sJ88C1lIU
DVMJRvGb0QQShAReq+EY6SVINhPH3kCA0WfkY6n6q9iMQ5ISynWLpfvn89INByky
HFcc4+JJZzvxnJPxaGWW9/2yYF33zCLQZIPJmWrWLwA9cvXcK6ZI0KszoWw+gf9X
ncpOhX3QC9YQN8SGYoDtEMwaQ6bKnz4DxyBvIdlTjCijZBnXAME0uUMBSDBepTFS
elkUSHwPO241hjO/M0DMOltYlzsZYc8xACqpWEyNTVBMdEKG2PLtYMXbdNLOzSe1
AmxHD7dQ1UQXJ1HDqKfgYFZHuz851nMGCV1ZYRK5bcLA4BnvFrycBEAIFon/3OxF
jdPheUc13nKWBABAsNkmM8f1bcdTYpX+pmJ8YoWZ4tUyAUc1PLbwwG1n5i8Tg3a2
11t163z6GKLJzE18uaZpvHV4PzVG+zmtJCIG1OQHhdiLXJx1aZgdLYvGZD5Q20sp
z1NfNAtyirtqynYsLsFdFLqb9FF0/ibKhJBVFApI98jKjHGpBLSxH4Vtu1t3anFf
QIOLfrRdTnvT2LqI9bi2W0bpTyBYVC10A6kauQYfxDgMLFfiu3v4Mow+6mbQia8u
R4V1MlOtaqYN+Att4iGQyUnhSjATrOFF/OtjMaPFdZ6CZASI+kHCjJmN0C4DnHpT
43VB9D8Thsn3hucT9/P6fy26qhL1Tag8tsWzwGkPb51DWZ3VBuaufg9t4g5uCwS4
RgS2emVvv7y1oMHppjrksZ3t51W/XGVL9Txfoy6fTgG/4szkLsgnyemY2dw80lS4
6YdOGHSCtSGQOPUxQT3e2tU1wtTasv1H+X1SxNyw+ewkprvK5KbyO27qZbr4+Zth
8NU6v9D4VklZ6d2LhOXUFo2Z+FWe1MykFxkcQoCCXImtoa0xIi5rNHGBa2eJhrFl
Vvn6gbYka/2poFW+vJRl+2ZmyDrOpbBZ6RGQ9LTSVPnPywALYMc2ah+Q2Vym+xc9
cvPaB7PEesQezHo845BuRijHZ6ID6smx8SDY5np6/f4rVHnIFQnIZNnjSsWAIC6G
F6UUaIZWGK7i9I14a8OIHkIQsUt7kIeJGaUwxXL7/Pq9B4UCaH9+I9/bGQiMyiJX
3baeRImWR6quWLDwnY2dylF3hsODH76Y2xvfa4BkmY74sM5wiNQ5BXc8im46UHFC
jgXzBgI19Dj/zqkZl62pGClfOmgGt7OX0S4hisimzZDcuQ4a1krBC4bBx3IEFUfQ
pYCpebpbiYwlkpVJjUL8Yjyd9JtUYcZHX9cs7X0H/IJ4N2RSU/2++B16QYgRa3xm
9q4emZlb5gM2XWQzzkyLbxwRh81tl5MgLp8aLSnzR2zqyU+QRURsvLs/rweja8KA
OA1fRUEHwtpUhUfr+/RG/wvdEp/DE4azBHFpX8iC4QY1Ixd1uoPcMwTkZrMJQvJe
qyIWiklibHCb8wNlUC4R7ZwzGdls45b5BQZJtyAjAQmKQ+Snh2PEMpYi65uOT6Wp
ciq9o1TTRYe79NOUVNMzdpVQQMw877GXpMInKsvATgc8ah/i+030qkm/hYZNPpY8
ymofhXW88mooy7x2o4L+dTt7jKtJLAu42QGhTAsMz7cEobqVZqC60oexgOUcxsoC
gngjXniBzuiNBHZ97RXp7tLOmcEa/L5q+CgEbGBTlcovHo1VK37FXhi2VD8jIeCU
BHMESpFmlkGzVnW8oR/DbxquudHvDl+qIFDCBlsoSFtbneOGk8lpSiJPbGrJVTh+
Qt1PtfUYIy9zxeXH7np2ilNQoMHn+qUWOd3DAuP7+7Ze1d5CemRMVplUYYhsU6Ja
mXU9yij2tJAQT+l7kJUcqJd7W6qa1umbAiTMXNKofesBDR7rIBimr8Jxk1agHwLV
/BVxv4LpUVobpKm9M8oVUdPJ30u0l3jVl6ghHcyBln3So9xZ9mfWCh4Rp3+nKx8e
CjuO55j6BVRYK8ZeUcSRdyYYp9/vDtQhNvRYk/4ibpU5QJVV7hX5RoiSkQxvKOH4
DGODWbaztOu4Tk3rRsOUei1/w0bgOZ5lZfRYUxW4a29zMTaqqSgBd6gIxrau1rHx
yCmnwSMgHPj8rCiJBCq89nRwTaTLfISb3dksys2EU0S8nc6dEzN4LjKrmJVLty4K
zL72nBXjDba9ywunBJTL39nlDrEMPR9SL4IaqnYtu1YGaK1VNg+38fmwKD6g3yGu
EKBRIksMWZkYbkmR9eigNNnoybMnSVxPKTNky2ZRypxKBkA8uycrQuTlZAjaMZXz
VmBtcoaKO3+xAJ8t1kjgAg7GoEPq1C7Ixrx0bkrCeg5cwrAeJLg5va4ve1Dfehyu
mIB8W0kj/GEiitDGehnIbYFclmwyOrppYw5Cn7qStztDNSfPwD2cIL2pvq/RO4+x
UKwtYMArBTXgE7IOFp8aru7zXGFD8lpW0O72R5zUpJG20hsPyiqN5zOZy1DU3jo8
j8kNM4Yeyin8vtUNquCRrvXpcRQzDXIOSmw5ox5Y4g2PHPLPEYyXhB/lZZt9US4U
QlYj7JVkVK0fzgPmzewRUAy/ihr9Rk+UoVtsT0E9GYfxYTkxPRmMLaox3M7ytq/5
B0vUPnwPs5iugvQm/sx9t72Ix/fbSG9moaKWX+P5jafB3a612ALtvHvrYti91rDj
rmJMsQ6dTZN/WrEnA31Iff9KcwN7nAvBwqmM8TNzPQ59ev+m5M++FQAtTBYvLiRS
ESDUAYzUMDNXkBmfpkEYmHWDQ0ufRXoWgOxNaDT3ls4ibW4HaTcMEoUpY/qXww9z
kNKPFQJvwYANAQLect4C2V8d+RO0biO1pWOa8eKcc6gRuc7YmxDO79irH6U8yGmG
B+qnoDuQIFtwc8T5z6e54Q==
`protect END_PROTECTED
