`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Da6x5vzpBOXgjcV1caGBm/93SQShBL358NohAzmgR8Vki80Aw4y2qvegF1qyiEXN
R1yLi04D1zjhs3yqNiI/NbamRAZEwu8kzDXSu4WVXt14tmY20f04LBhIOmpSiWvk
eV0uAORQExeXcDwkNN3ZdRxALEEkUMbK7sxA/xzO/G1emYrMqQhrWYbDEndBBeqh
QZiolVup5KDoKDWHacW/eW7/ZTov+JUg2e1AWectwILHdH427eaX2ReJhMu4J4Qz
P1ujWNMOy+0bryPwYxTpaQ+PdoYzAAmcXGnESb7nyygxfDLLHbBl3Krl93PrMaZ2
C0Tu1AI6XZBesY98LPzJT5a19AZYTmczZGiY5MCgRnQ5Qt6LGf8uX63Q08GRzxKf
gvZ2KVI9YFJziSzjaUlzgo5+cy0o0mymqCsxuzgqxtm9SGuTUAAvhvxswvi1+1Nh
Ap6Uicf2CTe3m9aN3GJxvZRqIKCGTrP0Me+G5uDCMhm+UiANnMIGPu2clNV4jI+W
5IIxT4O6IuF0RU5RqNhORlVl+grKXW9fJB4M7LSh0FpFLqaFnv6fDm+Yn/D3g0Lh
mYMq2njSqdRZiUqaBVzLG5I2cqJ+pNdDmmHI+zn1jYImUKwhNzXts4WqM0v6wUUX
f2a+gWP4ndKC8dMCmRlCLwbXmhsBAr6l64wiLHrnBJV7bxve61Zem41JxBteuAgn
fX6/aFH1WnEpqkNsIrS/ac52uX/CFIfEgslpztrJWODMeX3VIUixfjoicMLe+eZx
i5dfY+MdWES6jBqlq1VSR1TQVuNFoGiwpc2kxYJKTdKF8eASjXZPTbh3lb4m5XO4
D1y9zM4vskf8RlKM70I9rmXL/4MKQr9EPAsPJFa5gn2RFWKvO9Acl4AHVEt+gO4V
sPYuCfaeFdS6WMQYax/JJaXWlQuJ1GZAK+liK9pAOo9eHKhxJqEkSEpJoDSBw8iK
kwl/imnoHUgLMgtEK0Vp7JIYMtS5JLng41SkrwOvEivfIzHIHpORuNZSWqDAW5gA
CnPPF04atttCmKeb1n5IDqZxOC9zmowvi4bjvWI7k5m1QNsx7cJNpbLlbQJtMhVZ
kxODO9lB6wgoV/Iswpl3f89BRBXLvzb0RXt+XWj7Kb2KolDvDVqnGXH8A4hrcLCP
feVZy8q8d17yL/HSzXC+hiFRtBSKbGjX4CyKcbT/bUtd4FA2fHq/+MRfDbRLYNxn
YqnMHiuIYY9h+yRLonjo5TA8MH8zX/WDnMEEK7wpbPQwtlJvPlQfBUKB0BSkcNKb
0QiNVhGcPevndVpf7qCeJUzkGh0VScUqMZM+st7gEtHOkMfUKBv79ye5pObvDWd2
qJIdOwB0GdyEE5Pqf60cWhDVfrXIxyX+T9zLk7SofOe/+cKPwXfEXShF55KrFPu8
zZG60BEwditobkQrd+aStt/NavwfnDwcABhP0DYoOUGL4Ls/IV22sO/uMEBZE/TA
t3RsbKuM0w8mvl7TYdH+fwOS8TYVjiLDTvwqRiJoTVFQxQYSSgP374LygQia9FkO
ph61IVvQV871lXCwLBiWeYY27jMMZ3Wwp1lWKCooHsc/3WOmPnN150PBHQQFaYSf
urQdsXyGw21Fhj7JHnNTIc/w/DhTIQEt7Y8CtJkiffXTJhn46+kjhXa5ZXzfmOxK
1PzQQFr4bdgt98Y+nbv/Q90j6pxnJrCdaBEsjz5Y5Vk5nL8Rvkeb3uwxcEy1qQmd
tJ2V+3FgbO2HiH1wPqWzvGDPJEnFmdm0H0pjC8TBz0BVl0CYf3r+r8W4MjwWZH4G
agmMHGMMrg9O7d+yXIzuRyZN7FVP8RkR96S7NG1KqK4s5ooMCXyHuf4xBs4Ysigi
9ZiQdrgq95uu+9D3EgEjv8TsdG15qGxASiEXWfgnFxIQd/2zQ4actnxxJZypvCyq
YW6nYOcrMN6sASAC5gkybqeGLHCPMeojQfoi4sumHWtGQBTTZcqwn0mRnLeNaL51
0ehhli269thp1DXtZkp2gV76otTyKdugM5vKUTwQiXlX0jV2UZL7MB/sH8xaYJh9
XGZogkbyaPhn0nqPnPmxwgWzYEFdjIJM2Pm4qAjBMCxHXZ73Ey2Edd3iESiqSVtF
0Qm810xg1e8odGCDkO5o1IE/sYtpjeJ1wpFArBBShfzP2q3Jpt8bn3BwMNJ6mZm/
1Qk1KKUglhm1X912KUm1jZJAYUWZIH7Io5prBu1wDjyDUGBLl0uMtmFIzgqHmWRy
KkMTiEZxGNYLqP0e6f7olTtlPdDjq2W/d/IVdbEeFjf3mRKxnk+kwwq1z/j5X1PW
MCbenW1Cj8fkKBjDEbVcEntpjhkd6ctO0X4wtJb3vDhNu9YRNG4nOO4jT6BP3ZRQ
xZXjGiRw9wp8HCL7Vdj6SQqM6YEAg/PhSOrsQ4lC4LYQZGNsKJlNk/CRHPjWf9Vq
tHR1CVZVX9hCkEWaM3hED+UlfzfZq+WyVJTvRuPUccQi4MY928eYaccu51ePjACD
oem6uYOVSKI4MVvRyaywaYnrNbCSwfVQTFl6bmajyxjypLvA6FnLcTQhdzHB7OdW
dQD83CsR97kOwKlFDw2OfPazH2X2LwqjKB8lTzBIiOblx/N9ZTeuYDBFlRfYg2tE
wj1i/uAKLe5BqNHJvaYaM+U3T0O3ACztuOYo5QomTsu58caaCT/k5o8WG381SbDC
sb+KSSHOdhHyvTNk0lX5QeIFhWjzK1ISnVahAaW7JRdGQ1/aOTox6zCOq1Nz07+w
bPmucRN6bLUEIwWxLk+K76q4r/KdRvyMfx7SBBOFPlJjxFkGu1X4FNmQsXHcPKLl
i28vPJ6231kwOFUEu9V+5dl6R1KeWSN7odYC7EXewjZW6REZ6j1NgGEDdh9UN0vY
Mb95mXUT1ENDuZBoDYbqcT4BM7ga1B+IDbceMltWDXnFK6N9FtCZCXr0lT32PVG/
cr6/MuH0ffOUg7TNaKyVD0wyDAa1BaqUC4kVSutlAaV5kv9q/R2e8IHjU4JPmzGY
ZH2VgzDDpZGdt0gD5o35TioY8lTUB50C4JaW6S5cczhanVkxfxdNS5BFlv0GOZv1
fS7SUT9f9/DETOn4pIZxik/gZcJLysEkC9KEtV8M3oxSte01+tATPpTO8U9gSmcL
lZiOD/l4xAKl9+mDqCL5BIXkFDJfvHXN0UY5X9A0J8z5xLqz2Jx35Gp8/MGWvLCN
+dt/z7Dy2blwGdcnh8te+W80+1xZVeP0NRYD/iJdcf9glckpJ8X87rdjPOYDUzUo
D1IuT9aFYU3kngwMTwls+tJpDC9AyBaCiIlNJIVGuNKLwRyJcyveUk8FYuppsDKa
rESMHqDps3hzsvJ1tdu9pVLzyNuU92PN8+pEOPmN0is112hhV6VpoklOjtjoFHFI
dG9Mrmf64nPvLCE4BT9szByOGAPd2r17iAG+xod1KHiZJla9qpCHxq54aGFIlz1/
Vj94rIzj62U4RuOJJk03sQdHOdiPXv3AepsOQTTpWhAfp/ZOFXpBqvHQqZp1cSzG
2O07nVTyA+dkTMnWYcOAyCxGBRLqrDI5JbgqCqYlQ+AsXu85v2X2SxPH4fKHVroE
4UETscL+FpTJnNjiTq0/LFJyDMHqTZtL+rEe2PvcoRbc7b9YiELl4jH7hCPlmfaa
gidit0Zxe80odkiukN7zbdmEtiT/O9jb6IMu/Lfzwl5IcTr4Dr0mwuzzkZFDF7O5
ijevHh1Y8NYalURGIIgBkh3oEMsR2vlOP7Hw9GILCoCaVgsLlX6GIpL5xCtlgn6F
5YMd30IArfoK0+EDLu/rDiphOPRJ0qeZxwS8D4uH6i8tmGlafOORrI1+trMk1VEJ
FaQ4cBGiZAcI8JKc4vjGxboowehVUrIe8PIw0x7skhtzc1popmJn8qqIldNHfOO0
9UTX3/KW3XZHRZYPRJ9QCi0VPzEcJP9Yf0lDx3TiJwCITUHOKaCb8vYizxyoun5C
UU6V8PDpTjy0zqz4TOn4H3Osqgwt3H7rJ8+dbBIKYl5pGaaxQ8TdJgTa62vqS8TY
pO8hMRGzCDwxcBoa9hrLk8bk5Pz1xcIE4cHgmC5/AduHND7tHFP9V8g7M4kvPOgc
qXhdmbtMv8+cgDOp6MqTf8PsUn4YXQM9GzVhVFHa+zt4uH8iFjuGfmHVMrTxy2eu
wMbO+L6XlA5qfgJYsNjc+Qx39k50Njwh5PXurl75tqdHWYZ08hRzcMTop8NYY9DL
SFo2ZyMBZLQuEadD+Y80COlL6Yyzc72J2CI0eE4NTWJWsF9BKicGP4WxPh2vGsgb
hGU+XKf6OgIEn7/yLe+7DnIpiZW/qN441LZ5wLt8cUDeu09BLFJ852W+Nj5HgftA
kgMMDoimazY2IksxAPATw0jnAB7tqOBjU1CHOtyutZVn42scZcfZ9QvVzyLsToS8
VDSn3tV4IDTYwdXcWpzFbNwRxgGWUOegPbl9n+9x3GgpZzJZyP3uZQz76wFMRo9p
LsVKicrocMENucjn7JgZ3zmVn/wlR4OktQawwhC8mXO0AbvsgzUrFlcHrYn/mIuS
fi2Ja4TrCZvy+Df8zmMjC0cBIEb4rwIav1d2K13FIXIp54ErpMCcx7FzUb2//Bdw
RZZ9Re1RqL5d0k+AP+lI8oCtMRC0zM9V7LOWJzSRxuIflqEutoXgTC5LiYlyseeO
mCrshaBpeV9cEp3A3xxeDJRlwvezWd/vRSRqIfU8cGFf3lu2kZhFvlIChXiPDSY6
x/HliXXoXE6FUAvGiXDalUKu3lUH/LIp28V8TKHSPQb84KPSIneASwXHaOKZtasq
4iKYknwjLMTJpHXOsB5iMdKCZWQyd1JCYAzjQ0XQwcFY0K74H4ae96KmP6waMJOy
Jr3KKST65/YCzh+vhwnDwVfcdVpppF4ibGzPCPXcCn56fvtDKtUrK56NaGI0zbBg
5e6/12OrOAxUAYFDcgMOKiMjFN6ECO0sLwr+EFaGxhOk5wApK/3w6dyzBZULt6Ca
QGy8HqeIfq91WZL8sfvizXjmxh8qtCtaUHA/CMx2hx7Lvp1rmx6iAjcGBN3rVUnl
dX10x9tEnmb993Yx8hikuiCNUBgoiKTlGnWPHfxWfnPKh37Yb3J5JO0OMzbUkDBz
AsOGPvWlLC8yJkW82TTZClnJbRpDDKNTXs20N06UQWXY6+1Uc1Eg/0dIy1L8XaWj
TYxd9/LFe2Lx5dhy0+yrhkWRyjBtPujcGUUnXMtEMBrhU9TzQmk/uQ1luKNVNoCg
qB1SO4ZlpG2HMyPLdtxDrIXucPSKrEyU77csm6kll4ljHZ76vu7dR/HrTXtmFTf/
cy6O63cxZf7RktLJ3r0DJptIMwCH3DQ5SWP0kGiwGhNc/7ZAlFBNWpE4VP4Ueqt0
0TvFSaUm1o5xaSpFSR48c8g97H7V2WvFlAScCla4DotZEtk8HSBnDZdx5D2qyZSX
CWtxpqswtOvUODgIj9aWYR3yL+YErPkKSq5Q00Dd5yeFReIsuLXIsKJsTpUpXVQg
CzxvbT2QSCNrwOHahDqSIBCYBqlBH3IPJ6HlctwGo8CDJcMWxGMknDZQxw0SAJcl
0epGZRDZZCtWyABJC4etSvtFLOS10yJdDvqsc6gisH0fW9DgxmGNBdL9GpoG1uF/
O6I3LA8VLIN6fbg7GU/Dm5cERZy3MSSBr9h4vUZKG1T38beS8Tk4CsRCC8bJ8DEd
FKjJECrw5Q1FKEreQcbu3lA+llqgtbP8Z+9wfqn4DEe11w/c1bDF3qcPxnI6JaW2
hcFBa17Oqhq5m9fJzvZiKjOz78yEnKhdB2caOmUbvFjtVWHlD81o1jzI8iSV4LNR
rTsz283v5qJfCmoNnFjFpt63dZnu4TLEmhsqFW7RkrvToK1ZNKrhNmpas3oW7M42
4avAhbHdXW3E8XGYPIZpaxSP2qZXXTxJcZ//g+5ToYKm1m5yz5NOke3K03uOZJ5M
mj9p1Xat1VXtG7M4ZRQEu+ppXIKepKHpmp0zG1XAmlKxU1TcJ8NMbPnxdd7Ygp4T
9B3TosQDW7PW6E7m/6sAQwY3ODQM+SwrAMmsLx/fMn9UR49H8iHn5zJ4g7c3zqTK
+aJEUJ83DP9PsgJwJw6pSrTR0Yr5IQyc2vpY7E4OJpxNmFE9tRkigRGKcaRTuN3Y
nQP6Vj2Becx2GheUzj90T4vjKpl8CV4sR+0wA/e7uhS3h40USpggxnXh5ryJAeZc
C3Utlef/W8E4GZjCkFWAPDxeymalrYHIb7pDcFVVffe/uo/0/8xyRNpl4c2NX+pT
roD9C9px6mXYoPS0XX80Y0AB+19ZbuaBlie1xk4HJXEWN+uaEFppqRnhzDFPv7PI
S4sx6ApnXXdgsB9qMyD1tTcWdFpSutV7grzELmEoRrOOozvLBARsGChC2ZAaHXPW
VVag4sKyRiu6u9VdOvHhMtFA+spk9ERnxKQKAbCDdL/D+DDlSdfKalurZkqECCcX
2QKCYGIThkvNy2c2wGro3iLHzDUmleRt37gDm6BMtrYaZffv4k5llDtES2XBAaxm
rIJIgZ+2wInpVrs1x0pGvsrCHRuLEDhT6QvEOA4eWfNW0VZgAXV6mNtttyYnZGqY
VcIr5Bo2gphil/C1bs+UtEpSVwqppTWnvrzIUm77R754MEEs8NU6YMyHRq8vCtCw
WsLEET3FOfGkyj9/xbdqivH3HJXmc+CrUwj5OQoXYLWohZPxD7Ss9UVT1ZZDVTTa
v2oRMuAgjDA5/dTGuFtUniv7SEOzJTd96X0X45kz6XuJGUAWMVUL2MWf/O5AEre1
zAA4lrJ6MLzxJ2e8kR7CWFEXWOlCraF5qIZ93lWswIyIb4WmiFpIV0sY3liHkj3k
jqBXmv96MZ0mujJCedwHQtOn4giN1CXs/VWCsPb7ylqe+pLocUfVl1rP51CmKeIF
VcIc1dXPnR7TSxq35IRtvy+coeynacGLOzgVT+TE51JHJsf2RvIEAaBPwkNSlgIZ
Cz8CYwUKFl97rMIhdkhK+ulTsuOZTG7+o1ZU+pHPQI7DhhcfOAcQ3R+o0rjvolau
viSIsCx0e4ktN0rZfZb1DcpGH3r58sW/2tihjG3xU5hq1ZYE3xHiMmdKlFX0eyGP
bB/qIjc4uGKmclz2/Pjz0as4/dYa8pA+3x2mUyIUJ2ulA+aI2QxxwSDW1IgTrSwf
DFOudk9xsBdNP3tfBcW1xFRqhPd2NGaBRHpHADgZvYpfIsYLEGUp4GLpcytsZ1TH
C0pATnCsajU1+XdXKJWVbpO0/rMI9cpFCF6DCgjjObRVKWZOIHBI83VwBlYeuPD2
IkvCNZl4LFciVB60O8logFJVqOWCch7xhf611zXerkfAA5p8qbpESvnLZikg7atk
/5DBHTY2Gs9EW9c4O2j0fRuQMl+Qk0SAM6eMpKXaARqEQJip8pP9gdKFs6gK0p1X
yxsydFk1U7gSOOchYevdg/1VVF3YT+8SuxZQ0/jGdoQ0Tzol5+ucH+1BTvqmpGOb
zaIaT8LRlEW6e8wuB/JDLVKaMg3+dZQrC4bSC7LiI1JM+3Sxj0o0Q7I7T4zUdzM/
NkkpojcwlWEvcR6uGhoaFRwP4j8u4cOmhlhKSw4FiaxxzlO1SlXXdVA0+BptBvf0
PIIDobld8Y9b2Xi/NSf/U0V2YQxXcKAeraqCDvmhbvf+yh9Ja42qfxsnxlamwI4d
+gbiPKYoZ9faUy22/gV11FvzX8vEOD4XcwkTdzmZHXUUxzq7Qdg+xyhqRU8Cz0aL
xn6JfheAzDE5kT0AzvEwwfAXbKXH3pV9UpFDH942+EA9MHNK8gtt7oZHrt+X4xV8
7OevMdZz9+NXVKlKn3OR7HNoXBx9Ud10BOsk4jADH5viWvtU/nuTd34fOkD9m1Xc
zCZcuaLH5VQFPwJT44ADJhmihelvWRDEiJ28lMtOmoK8Nk+i2TSuZynwW/jZJP3a
LaCUJj6DWkXfAFYqZ65UwnkSVAvrPyZfvZDYJJZ0wCLfNaRcafN122uf9eGrphSe
MM0DgTyT3pvv+ncqLm4ldxoyDhyXz2Bbq1TwJByv6k/dl0iRZrwProuTn8CqCOED
SopMCkG2vcUC8YvoVBc8eBGeHK/hlvC7fg//gQtQ1aSMnXGFb5Kord6s9AHqK9eV
7cjV65JPg/SpvTYCLKIHMhPc1U6ui12nyq+EsnIpl3U/H7zRb3ku8LI0zc4W8KOz
DrdEd54o8+hFYxOVVO1J5gs8rVqLxQACfdcGprjll7sEyEmdNZqKz5tMLIhCodJI
3AZ6H7hS0bMJbzE5UJ1WjOb2DYCr+LkVsH2aDEMjfbCzEuZ438xldejbOkjT+/AZ
TteGYZiGbQuJsrY0IAubZc32FPR+buCffN+U0GfVi4/DuSnpfds9/y/8KNRlkjHn
GcmSlXi0TGvadtmP/mx01zvmM4Oe+w3TOia5Ka0vMVn9tpl5wFg0qyAg1ZuuUG/l
tiVi1zK/a7J44bbRdGqPzH3QRK2NoscwLEo+wEIAzokX0Dlk0Q9/IFhvyNr8sKpb
ATKpmHNE3XIGhweBeY2yMXAJ/o0q56NgoOLnz3Q51dnOvFA/kzBysqaWM1i7v6Pi
PQcHLPzvjR7zcMQuVv3Y5AC9N0szBmi7pYHtIAHtfMuH6O5DyyJB2Kep66OSSxum
JeaTeyl7bZabTkwprdeWkilik72HN6Fk3kKUMRJXUhiCPk4F542DI8n04XbPe0WG
dO6+iaG9LvfWcXvUtMSQMmu/fmJWkEMOVhutQ37I4pfG6nEDQMtZWzMPQwk7tPAp
KCIbCBQP973LvK2RnBp7P9okM5d1L+u4HJ+BeF4Yuv9RWJGWSqTukCD4CWJfNBLS
LF/lBxmpYKG3Fh8puAJooxCBfSUxBR20ktTPd2g5k69ODIt2goKFgbSRpC2XHAQ3
VUbmgrPME8yxLocgvRz1K+a5C9zeIEsiqtAOyniKl8EeIH2GjprekcGtXh6trQHD
JiWwmdpa/DjjKorCI/JtP0Bbcx8m3Jx7lJnTXsvJIyUasVrOW4F1iA5TTTrx5sVe
sbRZ2vPPJ+NiSLJTBcsI9UkwSS/lXkLVLYsk6b9U0RN+mHPAKINZLG/dPEDbVA04
RQ1WmwVURTT0b1Nb1SV3fbksyk5AhK6sOroEkH2SqJQlvbQtgnpf5c6wiaOSu563
BHNtLsKChJRglJJZKdNG564Alc/3uLz6lstxeB/mpvU6bJTU5I/FXPf3qvpKKrYk
5eH8YZbXxHtPY4t9UBMi67tOc/dqGKD1vWOXpFeJklkyEg3bS3VdgoKohFLI8491
MR9/7jk9LPmhz3V3Zpfx9o1LXP1DUQMBS4RHPlIL9dBYsxJl6nuS+HuUxjQTfcMc
1TFwUBT5O72x2dwByAB7YB5bu4Zxezoqd9JUOcVQ3sP5NZcSnzXgSXjf6DYnCVN+
zXNln1UiVBfwgGb68OuIz6tEfBw9Zcph72BctXIGQqmh7UNTxNtPD3Uo+7n7G3e6
MvQ+z/WyBerTP39iSQpMougrBcJcF1IQvVMYDQtX4YmMtKzJ+27WolXghkBbHALM
fjuq5HPq0jdGaUER+PIqM3k55VtBVh9Z52fxyVlUxfnQhaba7PoNPbPCJ5ltolPE
cHpVGEtpYzoPgchV3wkBVO346oA3aPu6EUJOaswcHs2h5UExSIZ8VQvMeJrXUsnH
zQ3eSRG9Teoc/MtOduz9K8/3d4lo4ZtbRk+vFSG+J5IEHSz3s+WBIUC19gM4zEMP
vcH3Zq/98byJdJy/zHEL3J7yVafoEK5r9b7cn1V5b5aAvLZ3Y0QSVvtt/uaTszWe
QYsuXfkWW45zk7o83l1WZff3FNOtoc9XmwIrSc5OAZ4X9NdmTAeBNRMNayCQhy1d
NiIXwD1wVQFH0mMgOlxVzXQZiXQ3DUVaUpo1NVYYvNJDEmAFOYJ6OPW6v0SHumoY
c8MyjAYPT1OvSALN4WcKw8N0VnL3JavMaMIxXEGcfhaeEGl3JAGl5TV5SMXokhLe
U1yVSRduamaqv/z/G1xJ9OeuStD1jpo0/M4tv6ipNthu09HSDqSDSJvUuy8TBxHS
h3O/QMsbLxzqi1HYMmupk+OltRRB6X4GbIznBxSBI3YdlAr0Y4gcLPjEePKI1Iyt
TvfrU1ik5dazU9KbseFODnHfQhRqvQ93NB6Xmc2+nWJSosxMjd9NNsjyL689i15K
ad5ecRaugaSEHCFsbNc59Sg+gS1z9xxATRItzSwu5qICBFF2jIyVK6TahTm+mK4E
Avwyr3wGnoMFJGyYjbl3dzqNZ4AAWy2iYnTrGG2VzYE8YwQ/YKyrI7i/XxumLDrA
u6+yHIzdbEOUcex+kWpw5FCHA7coNmGnr35vqEvvq0XOfWTxRVUYKcSnSA3g2vgl
KITkeq9DHPvaZTwNlUzu8cSC0B1jBy/rLtKNPurqwB66gK99skv6Aw7yIdILpBUp
sn59PzozDw8XUyNXIVtzK1pWYrCVI0kYxZkTOyiX8em36KO+wuenSb/MvH6xXXf2
NgWM7m57QLgekPYgm1eOFrqvVMRlJThQsmc5goUsGbdS+nfI6BM3D/mS0c8K7uff
tW0pZ66WVcLj7oOS/w8LAntJuR7WWhYAoI2LhuOa8rNEJqxn4hgKC/q3SNGDRely
lWqq7a8TldKNhMCSeB9sJP+qqPZquzW9y2v/aRho2QIeIdJPO3m/HNh5h43T2/cn
h7jarMGb8K+F1dtvIUKeMPd/IXBoogXbDIp5I9VUDAYtR4ttPOJQDG7f+GyR2D14
FFSBAQQRG3BogdxNjuwaM7gDWOfqZRyWnhd7MOaBMG0sT+h1b5moHBlo7ycQvg++
/PqVGbImd/cJM6UAJsGNdAgoCpmuPgymh9gnj0ZGXpgLKnNEOofzPiC1sKqK415L
mxdDpGGcJY5V+mMQvuxWmfGnQiuNV5rGQ6jQqLc8AW8j7+pWM+BGQmGzWXinU4pi
5+kMYHD0KTQQ53aMrtm3FiPxg6Dd1bR/X/3NIH1NcxjCv7pSG/PLzjEHenV5Zwju
R0IhI4Ek0RGjd+QK/a8NykMrsSIYM3NgaflaY1CPIDLeu0ziVI2q558D1TBjwGLd
oi+esA8TJ5FKnoag+b7U3MVeXAjn22QN/7SRAiGL9y/3/0WFgetpd88/R+vX2FiC
LTRCgNl0ExwWElIAlvNnJHdVqPlh/RDlATKc+f8yQhqfR8b2lEwTHTJbVsCkOoC9
ma5D1NUb5tealJMjIpJNuislb6CIeJhfkP4eMtK7ng+MNN1v5LAnLhXZttgysKG8
1vOCEdO4KfMcSiHNt+qH9km0mzwV07/2ICD0ToLcyEYAugRtVnNWf7IR7XeEu20S
+UXyhiKmWR67WV/M7sgu/tk4BQYq+0PVmNS3a80HDNqN7DWwO84HROP1S7mzv5xj
Sfe7mB3R0tjn2+Bt2GHCel4csd4ObgNhvCFZnM2UmfJUhCOd8twGgivSclhK6gYE
nJNUGB7084bYK3wVhsTxrLez29rh++a8suoQmXghfguAe20cSBMNdAbZvWBJ2Zoc
xGlG0gxu+5r/82zFY7okxA67+qM5Bjc0SbVLVafPuXYNMhW/L+pMNXh0+dL+5Hm/
gzBhE2YA/K26CZlaSkr83zpA1dzPFHLrc+Bw9fHP6YMQCfurjIOuojl96SFoNLNK
SbBM/zhFBNmV1pxn4riZJR/Ghiy/Lvfq3OLppBDD3sVQdk+mM2QqCZbnoHllvVlg
q6JynTa6ZgwgF0reSWvYzPOMpd1pptESgzoRB1gHWCYVspd2j+wZbzAjz1Y4WuRq
i4COcPgtV16UuesoeYdMuY4Nrg7rx5ODZrH4ivN35C/+qn+4dsM14y6aQkIGIAS0
TXrTYWCwQtclvTpSQoG07k1+9P99IlTQYlrxSnehFCHx/493wAaHyXuNfDK+uml/
ddbH/vtXutC9iCW72S792r/lQS0R4x4ThZ4acYbQCvaUN2wCmVdcMNIDXlb1idz0
eKiXfEhAYbGElpNV/zOGVNKFhZ923Pa5Tbv4D9S1ubAu3Tl6ooPqAWCJgYifg+/v
z5LZ2gkBqMVm8hWsOXV3EFP373aWtIrFmuZQdk5Oz4kVyJzTMDSXH9n1z22MZ2ml
lOLqiKbN16ZtVJ3tPaVF+jVC/45ZZNZ1+4w//lOzLzpp/KO+auVrJFk8wkMt74AV
3O99FcrzE5RI848Oy2bmQgnQavw2yNMj1y96ftMvvu4bxOfZbHYw3T7yuQvgpi8k
Zh8RRWXbqVVecGFRh38XVLs13r9iggR5N8fNr8t4vfV6ZhYbrnc2tRYlnjuGvafE
nweXScZcXMotmz4iJkSSOZhb/05JXQry3Gzg8FVUWuwnR8rRaOeOEa9xBNwWGgN6
nqNzrNtJD98oqtMPCFq0Mnd/eJo8OR8Z0Hy2kJG4Uv7/zwTN+ZUVkMiSmx7c38rn
26eV7hD13Zv73WKj5zinGIDTdAqmnWqunIOvKUDaqE55CA9jyyKdJWaBkRacOzGv
VUEldMSLSg1p5JAo+JcCeXsVSVIXaqc7M5FRcopnsQQWCklrTCrZ7LMbmvfmA7y7
Uzfm4ahN9+E2BmqCdKLP0dgzCSj2RPS2qE1NEYVuTiLlJ0MZPwczpl9hqkgupjqc
ndcree1/EbRE8Ex8ES41775di22YihBCPMICxR/zkP2oADN3oNpEGgfT5WTvL++h
ZZEjbE7qiWhOEmLZKfc5nb3jHSa9ayL+cCTa82vgNTopQJ25bX5dn+NgYqeAe+EV
eppcl1zKxWfaImeNgpV46pXKKABN9nrY1gnMkXCgSadiWtceHeVngLbgvze/DUYv
eYevaw6tNWPiiHHlMmlCPuM0xp4Rr6ZgAZGRRPkM0pKWKIuNx1VMLQBq/XBcA9Sk
MGb6lIFAS7z4HEk9CwMDLqZbwMWQpOxhuB/Kv2U/6FqN36m1kQXlZdzkSH9IRn1d
xkmRMAof9B3GwO+25d5AVzqNEk5WzsizUXXRgDrhjhH1b+deKq/bapn2Rf+G1TyE
bvGsN485mKinH/rS0cjiv5UXuC4P9DIb/AxOUHxvixQwxRsrELHrHs7YvYgS2vfb
xkZCqdVfQnGRA8akFlg1UdtTNCVUxXn0rpp253wZrsDpVOVvZU6fM4vNKp0elHOn
W/2GEv8FKEwSziavo71NItGxiccUT/Oz9bmkukLsMJ/tOE8KXXmhKZ8ISBhFSROV
wNM4u1KEzSYcY3ARhI1iwULxq76hSzCwo5zt9L85sc8TJhUj9reHfH9J+6AM33OF
irb0yCkneXXYxOyQbJg+YaACt7I1p4bqwqEypUQ9E+uLa3JbgVRWBmT4YGMGcF3F
5Z9gll8vP6uC6jrWn6u60niRJLPd4k/xKMUafvhyZ5a85oa1FhPWlMsPfBevYnZo
WL9zpZgVr0N2becx26QjMGJ4vowsge8kVuV6M1CmRi2seuNiS8oE5VSCnMYE6OON
S0RuyZ0xfgd1/Wtdj1effUD2OLW9JKwzSOExYFJaG8biE78tYPkIIyiYO5e05Iob
ADvepOGREcKnhwUY2zGp2u9qAT7SJOq4ONlKVH0/IPryjVLtasPIUuRBAUw0y9tv
7FJjdcVljzMWzgIglLbRByN/g0+cbPsbI/JQjP8vZXsN011AbMd/7UZy2vO4hHRu
drokDwiedF+Ah70T7+KeN3dx9MlWZ4RYRQZHQuIjt0zC9Lxm43So/AiT0/NVzLex
IQR6lIlabyFqqsj2/qbORpA/j5HBVWdfe1kHyMOWdoQ0npKMBm4A4AI+V2z1ImaZ
r0uE7r7j6vtX0G7bXkXO6prnWpCUp9EhymGavNYAnn48WJnA3XP8FTpKkaehp6Oy
TBksiM7a2SmpTedEKdWJ7D9PhFhZNBz8XkRosjVnFJgpd4beZRxcNZII1B4qQcB0
bqeXp/SMc9k/nYzL6/+fM+8HxMrg2k8lY6+uMrn8RCNXIMT9ISsnbVl6l+50RneF
WncRwzgtIo0svqfBMQhY195fydYxMgQxYLG709JDPqYpt+rWnLBQ0lgiT1bLX43W
z1dUyOhyYeAWGwGm9GwdfD//lAMEw/IYN/7TqD8Ype/CuR5zbT50xjtkXCsd/PeL
BzbnTOK/UOcTk9horUsE2e44uv/lccfvlpO6YgdOzf/rIVfBFXtKm3Bb94aS5Ijh
VwQYCtQxo3vAfXd4rTg1eM484V4fiCx0bp5IvbqErpibnnclz9BIS+C42zhjE5gB
Od4rsN8laC+SG7NXdNii5mX4XjpOfh12Rp7JAyBvJ5/318bmY166AzLmu2sdEN7A
bol71YiDf707/4dcE7QeaTV95yOtIrfzBKfxeG/qE5kPEs3M8RoX04ZnCzENEsFV
0gBH6hc6Lrkbyn9kht/IbTBSKOBadNwluvrUEFa8fK/IBvzYKGH5rAvhN0O7G2Da
hp+fsJNPn7XpCF/oXok7+Fknm4EOOFnozhd4W0GfreMN5CXrWKiglth4fA4ptFu7
OBoT1dR20k9XnnxOYjXxXHUca6xwP6KghpoSupGfiOVD5kfhUMUUxArgk1VW2vQj
UR+5AuB6grkoPwOqsYmFa/v2VUikteJdtYkrJel2SIIHB8nDUNJXMBUAR6kDuU0H
f8ZQQQ8gri6+f9Ym/7QC/FjHu0S5h4gICsfqb9cHYuNAIQqstsFW0j5dJQcQsU8E
XPfOMcVNKREVTjgx80+e5ajqUVbt70HDnbwbVLXRN+0+8Y2laKdgMb5CXE3gtCKz
/ZX/ufbAI+tsZWvNV3IBhH646hvxA0t0aUgZBeWN2QKxVhGb+cQSJs7ZL60VYuur
hbh45WPjROR8DxablL8QtKvtTkHBHNUZj5mYMOznn36K2j2gsZ7iua0/i2vNnixa
9WI0UHwX5dpDrdB4hb1M/Ulfl9JKKAA30eVpqbOM7cm7XlcuGctQ+Aq+hHI96HRk
NqL9297oeHqk4WZtmI+iheLeVS7ZXfew2glXGEYyq83TxkoxkSMYIluZDyaoTnV3
AhV3nYKAeOJTkZ9aelHhhiLevmEDXrrsvD2jQVuLsmkbuQJF8RzXzyOCCVMHRhuw
bAiIHeoq3YbYJ0Trd8wuzkB+1y14LZgZH0Rr43eXrYJtKf6XBS2H5wAwAKOPYVvt
hN76HWDiIpwe+5PrhDUiOWL3TGJbpVc9g63UKTCofGbTomu6rMzVAxb379La57RR
WqC6WkP2knzgtXVumrOy2Qb4XNiNYdu91iATcZMxYpS7IIk+S/uaQ0GUOZTRzlKK
y4wAeRxI0Tif9lv5nJx99fWGmrsJqCiwiqBiYYoXcpNn7Q18tD0wx60Zj0RYxLWU
lkzCiv+jy4vgWDBTgwlTaFNn8y6ORlb8KWlvu8sEBsJsPJLlMUHvMl9BQfyFPMEo
hAimoT8vhu0PFe8+Qzvr+8BZ5msVzeVEd69Rn7OrVIzpuZU3/CciV0hZjz8JQt6F
ogB2qjTRvxpj3Ila7AlLl/Kma5Kv4MDPpVq58zuOkT0A8c0/MJ661BqjAeWgRfEY
akL4YAwm9mQtcpLwVVCvevGUJXaOqFiRW5u0AaPSGe78RV0JZ+BGFed2DR84tvai
ZxUgxknmdvJZWUpMyH5g4827PrEtCWy3usf2eySimAQv/Lxnj7AohG/sEwebtIks
jYB7crPWARURE3Z9BKZd169rTauqDxnZG6EYABFXqEuwgsH/lUi+nyY2vEGwxenX
qLrrsgCtlwR/rAq+j3dvdZDy5tUVlBstho4fRdAlaGfsqA781sczT3ut2Rh9Gpun
XVPRD5v+TrthT9apm71b0lPa2MJZTKqzZXeWalMODboYuCitG4pTfSScQG7cMUW4
JQPsWPmXPfLth445z3Hmm5tzpVh6vwQWenAxkgKXPpyC2QY4c+bEiZ8oxS6ib6Ws
/KxJbRGG6YQO9KnaHkE52frpr1hp1D1kD6VSfDfEpzAnxtuL6KbwfO/tN4ipFOCW
05zWAB3hrWUkeneyJisrX93zQoDhEAYR69wxB15L+Rc4jd+QS5CLqoPeWqTAgtcv
Mo6rhMgcPQfSdWeRqXaxW95dZYcxJFaNJm3YAYdiZId381p/TSBz15eEsMjV0IKT
Bq3MGffatvsQFosQovxg8rOkYZqDJ/sj8PsX/ei4dJKG+xxHhKW5kqyDYFuCuaTK
WSaHkzsstUBqrqpVkeFoO341+U27wvhTlKDQUbu2IZs/LbRgWjhN9DGghnwY9Oyf
thB7x+zP0q7uJftDO2xeZtxl3Iz/UaQVd9WV9sEhtF9PPwUFvYDARZtqxiu1Q17R
jHYmonX4smNZlK37itVEaYJPREVmb/0sMjWC+By+9jkcm1KsHWWvK66dbO3ka+Y9
JgIN6n3J7O8o8ED6Tjw51rbW1Vde+lc4jw28RmQnFazb99VQD1xUuuqYNJXq/I8p
MoRIIe8OtHlmyA2VszWUh/o/SXmLmVP1W0tQTg4ddG2OSEbIvLowXuNDiT2wu9YB
t4geRkKS1Liz+cE0XhFOsq3BX+OUJExknHsXd5a03XSNkxw6Ohnw38/+U7s4QYud
Z3t6meNUG+rnXaGd/FGQ8pjjtZjuViAk5Fh+zUPw4VYfqDe4KyHPykMphXK8fPIm
fLl5mZQZZOVsVUtQiCg5v+d/t9AgnOCeum3iNF/SeSgSW5fi+R0oDHT9da+LlTVD
yv5oe8eyaZEx8oxfYOVvI3J7RC8UOb8rnqwWfEpwSWImZarZr3LfqSaYbDHz9Yyh
LV0Qyfiz5WQy9M5v19BxPjsG1wJkYFWzc+sKDooVcNW2GUGIQ1htq3Kz4pqiS+9M
Ydo9YgdDn4EYga+ITWZBVHQq4ZnjLvPDDMjolSBYB6uvkdf92813ubT5Ouw/9t44
gLiWPKzONu7UsvfwSWV5DDhYfHxF6gC9e2m0eYka4LOp3J5y2VWu14qrTFvX/zWR
Wjo+ZUO1K5FngyPC2QtQvcSasSbIpWjqtZ5fyGxNS98GrSF67NkRfYIhYZdUbQs5
xsl2lx++KQPg4Q0s27fSGz6KFg9KuTJkF0nxywbzAZsdghpVPa6RJz0D/8GKxRcj
EeJDIWgs374qmwbVfUTtkxIdw4BEHD3QbS5fEzMw0Jpx/8pv45XVaZ0ixTLvxGiO
KGKEQSqCbGf49itJB+7swLJMkgoHBro1ePjZT6UsywpU/pXkwC6GE/txrKPFdkMR
+rH87uX3EvBl6qn8QSusm5x2MzOUCif31WG5pUEs0FfHP9cxmQp1zkMv4RRABCp2
7rxmIlcrLjov/DwWODUhYMayYIovTc7fYL9vERSDlaSzELurjh1MuOSqLyxzHUx+
UhDNtO0gsetBzjQNrouoxesB9qVVwLb3TsEmXR/SO1pOSmOBrlMEvp7MsqvP4y7R
fYevx0G/wf2Jb40uzh9ZsofpaWTblH/iZGFcw8QizrNj9w8BCCHMUrnxL6yu983T
lIALM8RwPdr0UlOHgLNsgpr2Jeg3U5p0l4y2LOX7TdXGjuE+9eWrPsV/cggmCCEI
hBZmMdp+qI6SlamdeY8lL1O5FDLFtxHxV1MhMtHUMb7Spda2SVbmJAKZrNAIVg1R
SJpQTBDsam3Ir42mbPu9t3KTeyYTvmRUqK+1GshWqtQ1/G2ukcUSCYxWxxzf0y4O
fqkRmuDx5hSleb10Dqm3Zithfoh2Ikb9EAGUOthScPn6/BEqlzxCeFVcS8EsAR2n
Hd3uWc9um/EJYYa8EsFaXeBHmmX7zDWdC4iln3XVyV8GDmILAwPQy1qEy/9WlNLB
JNFASgC6HWMetmOT5fRgI0qRFI3cdv+kXGbYwDNcauCm5rkLd45imKA9nTtGXpxm
EG73gA9CI0EJn41Dqq8le3k5zjxUOdd/Z88VDnGz/xNDOcFB4mUo1vzbbRZz5t49
nVhyicxaVHBafg9uO7QjS6JkNh8J3QMPHY5K8cqZIX/3QGo9tmXCaMNj5NkwkTWd
tUIvFEGqwCuKRZMz9WWEhZLZ74oUxLR4aeE74bsmpwZecWTpaoOHJQv4hBwnQITw
mvRt2XtRzwaUP66OtNcrVy3DBiI6FOVHckyQ2p7SC5dqWbPvtTygx/CUwrkCeCbs
9sOp4cqinI16Tso3vvh5DK/JfoqTDOIvw6OjcuEkZQBh9WeAS4hzU/Z8twRrzQnB
9aEgKfJN0eFEIauI9shYQmvGUXxF43lkajLeNBXwY65lHGuFNKfBP/jYVpPTK1mf
Y4Dsk+VAMOiO+xXy8nPgU0he/IDjI5NhOgF1fE7zfgSqKHRll9Mtj9I7RBy4uUar
TVrDyC42z1Flt4ep3M/nrJrNl1Kun49NltcR3Smtsy1IlCFV7PR0j/1LcoLn6xdC
L6jJMw95Vbclfa4UWLf+Bs7Im+DBxM8NHNxozteiXYPVI1AtM+9cLOR3bBmgkIhV
cYsq20OBJ94BLP/Fhg7Y64J6vQBSkjDOqJoscC1waQ87kf7yBrnrk1NQOPTnLNA4
/RfV24wqhpXe3ZHbziuwJud2KZ9pBKf3yDZ11SvPCIAxCnCOP7wEkFkKasSzur3P
rYwUjp0D3BIQL0Zv8ZM4EZU2w/RgEMy3ev5E6GesXBcB1sa2e7xdU1ES4uzEE+zY
j3fKAbI5yp9PVfEaEnArWqeVaOmRBabjcLUQJZs1MxQAqarsiKmpm8GAEyyZoo4P
YGmeyOfCI1XtXOGJurkkk0fgLSfKUm/Xrod5wXLreI1cV/RJ9GWxSvfi7CeVO7eB
E0xzXurpnjstrp28CH9GOcXqBxh6SeEjDShVffgmnmvvw2uA0sgzCbSw9oVZmlQg
d2FxS97QkyCoqaJnt87N+4PQifa+8fr6ELUQn8mpGNbrzobUOhEDy2C5HqxDJ1+r
V97Ai+ue4w8FBZYI2mk73KMxPhyGEOKPehvn2TEf7zE4g6flO+nN3IKzsDx5RbY4
+sTBcs5HBAwBnx3YzPAiGNoUQnccUkXRGgXcNlejEWi1SvLd+hFGKiyClWJH8nLx
nnKRaYhLN+MlVoFSTw3iW0Y1neRCSU6slzTDIdf9wc0/08D4ryme5W6zq9I5wGhs
rarOqEkrxakdmXjCWsfbDXXI8um9ymBDJzYsenBi7qLN6An8+1Lf8KlFzFB8QqEg
nOussgGQLyNRuBYo/H+SQYP3gcX1rwZU6ka3U/tBiQLEX2gZPAgBtuodhSM5Cndd
7VST6WY+BNRiqGCNmsD6yJwZbF8lmylOSa76qe7KHW1MBYTRHsP6TJuC0QA+BRb2
m9b3xaLgI2OSX8ElKG7mrQrXp2HwWP78BAH0H1MrgNM0r2Hm5bPneejtJuy9hK6L
oFKv7dUSoAvop+h1Cz4j0fcCXk63KrbqqogwTLG8W2eSzy+g4N0mL2aRSKYCxUHp
SNh7Bw7Idfofp6RtUPwjqjik8/Kzg5p89uz7WnS+6ik4GoTL+lLRUAtP4/c2N7cf
fPBcnI+PIUsLs+KaQkaPKrFhMBbk2mLSdAHtUddyzhlsODtFO7axZjFSgtxDBHvy
lpXkwMbWKPyMbP7Z2Cf/4C0uL9YX3fVjpHuCN1wKe9kgyzQGQ04DL0MiajWcLkKo
w7ZPTcA46V7hYXK5axUiC5951OGLvrRlPSyWGw0hszEhZmS+QULlGxB3PJsicnoP
Y0rH0ilRocY1uBIkUegK2w8nIxOSZv5+ynZ6uVhRMaH7L+pPqGMyw5TSFTMDiTM6
Tucg276ACD+pM8MlHOGfMItm9h5aSZURAXtKsXyzcB37AcGDbNJGR6b0Fki6WRgf
S7tgL/rFkmm6Pw85Sa8QBk9AuHxDxhqil9pFr3ainpVQaMcYDSujJLIV57d7NlmO
eicvBtMsqcrxpv3JONWudNJof5OQJXSQJ80tQEadrfxPugEudtzKdhfuYlL8B6k5
GoY6Zt+UjmHRTDKU3XHBS94x+0yEuwgiNhS4I9q8tco=
`protect END_PROTECTED
