`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J4/xulHomqr67N9+gaR3sRQerP2dzRgIAUrs2kXITat9bIlXVEmbo3XLiM+AFQV5
S+8T5C6qZrHqztwjre8ikG1qvYAqC/mx9VqoCkSb7BYBNwPzkSfuAjY7AHs12pSz
uUVsZibTh8km1g6EJGxmqF2zosdhNc9uUXJNY9hPuDX2jtbUuCOK1OCKWs3xv4P2
JmoKfmuDvA+fK+JBnHp/rc+zZ49Yuc2FtkHaRLAZZm4b3y/oaVKnHSxWJgznCaN3
7EzHk8MrQwawqraCO9ylDN/L1sI/IuS543CmIpEU1PKtvrZ8xS8LH579ERY6Xq2c
bzNJ5JK8JWBNnw38qfX9d5kZy6NLnvIjzKooSygRCpxpWFhAsvKf6L24rBaXBDvn
nAysgEactpKAcIubBnZ4tfpVk2dH2OZXGEiZin5Yo83d3sAHlmDPtcF8VPqCd8vW
81qakq/qPqbzNgIQhlpILbNfYrwG4r8FaCjeXxnpDcVyZ8zS4R9J5BfROnVOG1UV
N7r2IMQ7nMrnzjcjo2zxBtwmKq+vEyL0jf6P4F77eapqNxjR9GbLja4+XaHlFdgg
NrvjswS3jNmQZbJgf5gJwE1FSxKGCsMcS0IYfZw4u6OjjjHtZcjurhsbFI9Qse7B
OVRMw0Gfc5DcGdRGU7BHSvxBaRBq7fh3JC9KmaLv6qC7YO3W66DhGz1A9Icpcbbd
MhcwdSkA97Ppa0HcxhnrHA==
`protect END_PROTECTED
