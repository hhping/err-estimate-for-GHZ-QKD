`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4vMcf4ZX3X5MzEcUn4tnFsUW1bYB3tiFDWX/WU44x9orja4QVNyGbp3qbTLzuRMI
17aKtyu1VaqSRnkW4C0qwm/5w34+O2kRF1WkfQWQkt3fxVP0gIiQ19ImWyNT/+N4
Wi95ZeZfgKO3T8B8Aw/pse/w5WA0yrOmtitKjoJ5AuitVhWQbb8Hkfc8YSE4Nx81
a5QH1Dr3qIxiuPJUETAaQVDIASIaUKLqiEu0IwXfOJWrYcK85musozoEluvpD5MD
eMiFgAY36s3Qe9u6Lli8Nqx7VJ0Glf7wsKGB0ApGqfA9qMcvDbD8wKnKWIHv0t4F
KUWFpI9iupepgIsN0fdLX/8oWdWa2Q+7DFk5N8HFBMT/Jjc4KgCIWsixZo7XJu4E
Z2aYtzS/RcQbOMsuXd9WrIR47LcAUh2gkY/e74gkgyYzm4tofXAiI6ZX5GHtd1pX
bj0/9/rO/Ts8LqFS4zZu3wBTleWLtykFJgJZ8s/HbiThASmiKnaWvzgJJtPDj0uj
XEQbI+gf0FvQYU8lMB7EWcSnU0VwdeV2dYVMyObKXdTvtUqMTo18BiCLNgNFw7Sn
lve1c0AN8wUzYDQfiF5N29U8V7bFUr3jUkoW7QmQjAeA5PFdapZlIcBjUizcIeK6
7WMUCyFm1COcbINCxpvSKaeiqDYFwQyQ5987OaMBWAidV/ZO6KKAEOLvb7mzMcYX
+SBwvszmTJVA7tbpGE1FHdvr45O457Njgys3z/p7mrHOSpHTadi2Z2iGURsseI0X
is6DrzrU5xMG+yhz5lXAATCGSS8G3oMagtzHzEThIDB8p58DuLmQBEDqntQ8nvFO
B/JhDmObGPpcf+I3xD97mgSyXbPvHXWWot/nC6FogDFI5ZIjcPD/N5M/duAXtSon
dKkwXieiuTcQUTnKv1kQoNhq2FBiqW/+c2LFXTglSIbqOPFpkpj9wVnrx/J0gDEI
elWZk6U+qzchCLxa/01zgQ==
`protect END_PROTECTED
