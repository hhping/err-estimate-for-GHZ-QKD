`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzAyW5Gy6xHOAUzo3Ks+9uQ4baIb8yzpt/m/4zCBlcqhOWeuyIIU1z397E+P+SzX
onysHSE1SmprITosdK+PTB09bdTqR/jf5yQZdjSa3gc3E3hpXxc3gZM3sdh5TKsg
UPFLG0DiX/MoIJGXD3OkZofjOq8d7xlI9SlpOyFpBO9Z1VP4u52GkiHm72IwnRKi
C+XMTgtOkKJD4+iwkTpw0HyEPMbdIlSUhCEjcfkLv3r6UV1zznaAHMSv3t57NcmC
bQINmyxnzrGN7V/G7rvJ14qdSMPrGkyz9S8eTlvXe9j8M2y4J82SbfKxtsT+Sn2R
qo9yWjvn2PVJGDWkORwv3Wc8pwTBnZ0MpihUh57Fze146lYnsITXo80CARSg6er0
VN+2LNMjm/CGP4bDNSLrK8ocoTgGmqng6MvO84i1eft4NkLIYQOcPn2a18Rqn/Q4
Bnacs9kmZxWFXwUMHBsVjoWgmpLtaZl7HBwgYplmSKFKcD/dPptghLxNICpcf+d6
ISL+3+DA4eI+k3A2ed03zJPqnWDMac2NLaXoeLOUqVRWTzhOgxOVD6+DSTtqHaBT
uHjD6ELSbnhTYNotT6hzjqATes7G9eWvzu0ytKbtRxP3JpYWPPbBCISJ9vZ/4JRp
MLIh9JMIbiYHFxje3oP5CxN1K7zdiXomSZT0TbLSkcF/NMiQHTBHCsgiOo19ohQj
pxBVCfS6aLq1N75OedyoMTTdrtJ+GzZQWyCChR2aOBzgtFAHow4G9iIJbilNDgTR
bl9p70fZbNn+p79Z/W0S0zJfO92u0ccVdcN/MtWuhzfrV6fRDLxi4sE6vMudsYOs
795WAnK3aQE8va8lLVMkaQ19xAvk39/OAQ6eZEmhB8r0kyn2tUSpQ/ZGBwmV4d2N
sZjyF4aWiCAEqQ4NXMqV+7n1dZaB0EpY8TL3vsSa4ChA+pLRgZeXqmfoV2s1zUat
n+rH6TrCasbmeAWEKrzXan6jY9IRat90YQ2dJNQyWUf7fmQIxz6DziNZjuZIMmb6
onp4XO2GMTsgBaJ0hhxCqNsp4/exYBDs25U0zFVT6JskjSloBY63mcW7OUblciwf
LOKutOMWmUGwd0lqTHhkiu4n7CgNfWCvVIyB6uvw1owuVHHrnZIox8XZe6dCM8VN
ZK2dzCBmxvzhNVF2z0pH0s38Rheu/CeyDbzquhLq/syRhG+7YIhltU/hZsZpcWk6
QbKFY8ja05yIdHDAbnYvv4OO2AUm+POtTb4MZ9wCry79+6j3ZRdwIg7ta34E/jsS
6rMxQSrezmmIiaD+begJNd/ggYWQdt7MLDftgqJaY0+pZohtTKPRZ4yyATAS21yn
sKu4DErjM3KJTAKp4DUG9+Ajgf1O/SOh4z0TusWIA1VPslkyaMmwLMYvKFMIffr1
XjuM/r7X8fHq98m7C7qqXQhODRMNrhWa/cE1TxRa/PvqtQj+POZu81mEuAf3G6Uf
so00Z0oHUorhcmoOcikvg9uj1ZUDd2YhNepEI5/x8HvOjcCUXhXd1oBrg01dZtQ5
KkrRpfRJCOh9ayege2RWxq/KiVL5miu2jq1uTMQ0mKZNhNDZf3BqYgi9T028EReW
TwP2n6zwZff2PEec2DezrFONi8l/9ZMgSf7zRxj8PDZeX7mvyLxJdbGmAWG/9o89
r1u8EJGUleWOCUKfyg4IvDkfeuO++b/kFN70wRhDrmyDqDaFWlfhywfOBgWWDOY6
ky0kUYZc48g0nr9QBq2Yztig/n4KbOxhxeFhuIqGCqm5ksx3QXGOy+2fZx7jcoLH
28z/Y8pMqbBUck4EifECl0eNzFrMw5YJppkf5tf3A/UJQ7gJoVEKyTw1BmlBlSj8
4tKtue5zJ14RdplLATeRwyOdGEgT3WcP/qE6aAEOpzbxWRcJyLi8p/sijDh3pqTI
EjZggkKAh5xxXd1GhGDOtyRxp06nIT2SoyqjJgl1CoMdtqEpj6QzR5KgKKMlUBG3
XJqhdNNTQ6VmlUbMSxNUHFapPQeu3jyTXrxUd1JWY3Onfb+WI3iILwuKuZ3x5Poo
a6x2W8SU0RxMid8wkC2xZ/+xSlCMc2C1dm5wn//y4GYJYvDV35Ijrfp2fpe6H4a0
GXFf5O8NQZRFKYVqO3B1sqhE7Kb1MzWFYrsYcXGL/PGw+HtbpXsGHiJlKf5ggM4G
`protect END_PROTECTED
