`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CjBqr7NJbw3o42sSv67lI2NR1s4yfRFor+5YoqsShshul681N9/MM3ZthUprLQu
Btz0pm9R6Sy5KuypDKK/3oPQqxs59RPmITGaBlZHXYpjf7fZQXKFSWkTB8ZekY5S
babc/bLIx/71VtOpV+/bi1xsRXJAHDCUwC16UF6Og+EEzdA3PYcOr6t3km2M7TEK
+r525GM90nkzWak0jYCn68V4h9MzcitXpCZZ2+UYZuT3yLvpbjqt9Prt8t8N92nS
3E4LhOIQk3FuzjU1vHHQrvzfK5H3Owvy2gpmIL7JaAyPkPtZ1Qqr6elruCu6pgrK
3ZYPHMHfg+A093vVDEY5crku/t6ZEQSaOyzB6yiC1NfdNxEzZvB+WfMWGnpraCvX
ijfSMKdiGHg8x2TwWumzvBvH0DqlCkkPsAcArDg31Ah1HNmqO4kS4VAAKrwDBE1l
HyGOcKqQzjpcVkug9dx6aTdjS8hueJTvC6QptTXbnzMR9IiE+F0EcTs+e84xIeBU
TRxxsvo8eUJRXD5ABo9+acU6aQjyt9WTvEpnHW3A43vRabpbJQPAmMBV+Z0ypub6
rN2maJ1ZifOQyYX9gzmdz3yOsR/E6ayWOeu5Ofk4MKR4lNHj8r4VrJFpav6QSJpz
Z1RHK2E9fJggcUrxUO/7n+QJgWX6eFpJDCYhkJUw/Jz4QfqWyPOYouZbtS/pewNs
eOZK3nmie3U29In1gG6F2sv+B0iRANqub9sCA0qlgqQQvm3IT7uqy7Q1ivqDmq8y
1bHUFnvG7G0s8uxCThRYPtf1h7E0Dsnk4xx47VZEapM6O/+wm0Ux9cj5C2ysOPxK
/5iZojM4Gy9qcrhYTy+pgYH6Lr4h7lpsIXVf/DGyC+5pbpbXNh3zkwD/UWUjJXgT
hl7iHjGJU7EClfDlNLT7HD1TxoZok/D+H0RRHnVHN3QN3ig7Mcj/J4dN1MREEpsv
aaduM4SL+52ePv4oYQY5nGNsT8C9XV7JlfkHtP+Yg7Ntwpniybyh+O4P4jz3WJwO
P66+LgmmQJe9h6wK7VxGF3bZsHSX2Xp0h78G0iLCsFuQOYTps9OyMsOla1ZQHMsb
5W5tY7HpV/lnUjB5airdRKuz8ti4/90ZU9ayqylVnjIznQ+M8hWbW2oyAuf3P9nf
7ZE9Shg/lXqx7o6TqLR6XghSjM8ANhNuypu58Bj0Ls4vdE8d1AA5iVPk2hFkt7Tr
vpDiJWEiKkxZCWUmI/CkIKPTVaf8FkLjSS5UIHtqY3MLGFxJD97fa3w9CSIEmhPc
ydoeZTdwXU4kycq5BIBoEhsCnIMUEml/Gy7+1SLv7IbJ0K4YwhvN9ixHctiBys38
Qyn7e1CDNc5IvVA/2fB0NGkVU8fJpFcFsJliwViPc97q1P3JL3CKAQqmmyL7q8vl
xPv7gScUgTZ488hcBW4KMdPrExfvaB+ec5cDtE/iRs8RkB7XYcm8ZEIPV/xVngPL
Gc4v/Fv5r60Mt+S5frgF+MH0uxof9j2KMsKL4mQiTbQj2qTd7RsG+sMFIoKz+T8W
IHWkPGOmXcnxHGhOmK/Rj/qgwD3cFDcKsTvdx0W5OGno1HPYff2UD1zxROU8ZA9B
NqKzbgO/v01EZfz7H7VfMdQQlAeFULeBQF4kSmsuE0ygB5OI1IjCKtvkOnWFL5LW
UQLMETJ7ovslCb25fOfO68MpdhNiDMdp5kWXoTK4DGeOs69q4Q/hf+GJ8wACjytm
wwTBRRQUqyHTnbXEEwFApQTcb2V4DrUsSNBQ5ZRxk5/k2FBzaccjev0Pmz9UO5C2
EqaBYPU9s1oCyM+rBoR0HlrbG2rzzmRveoYl0XwqLe8eXYK0nKxNhf9tB8fahu7A
LhAP689sfFUIn3gyyD4qJAV5VHOpO07Gp1xlNq9js2OzUUO9Ezmj3mU8+AQBCSsJ
wdHItFvWppkklbJcI5fEPaXUAIxmolfNiAU3oLkBNJl7hdT8Zh5KSXdPqoj0V10Y
Sgy+3YlzoyQcTAtmI3f3CFO72f910VC9DaN5FGIIW/iWNzQ47MyBRzrmGfkIaaZp
W56VGyA3PTJMqHM7fZ1aO2u9aysVkOsWzs6VNQlLWuGcFMkz7HBCVNx0Ym7iG3m9
e+eR8lG5P23p4i6/Hx0J8yOWM9n/w9W36x5JKztMckI5XzotKf5D/MfSh1bBPCJq
rBbgcNmH3hHABhyl7vhrGyOFkri43NvojKsC5G+VIXYyFsuIsycpBupxQ/F0bV9g
rbKdT09XHh1/zM7hQjlD4eKT+5XuON9dKtU83dAK4La9+yoCB9vsgDFI5vGvTTTv
UBRAc1gXmN3Ra+UuqKtn4kFYDCTGhBiK8aH+nCG4p8FwquqjnH7hFYYRn87fEkLX
g6k/ghPwDqbVfQe9zBttO/Jd42BdjIu4caisUMrVHT8zAL/p9+YhDLeIq86gXUaT
w0/3fpFGqP/2ZocFaeVxcSzIREN3uf3JVNNGsVaHzgCLF9YsAc+4SvfcV8g4nis5
9wbvm5Ota9mTvI6EwrgN8Sngibd+eqWzolOcKjswqoW4asrr/W0FntrT0fpd9QJe
GoigOdd6FoUjkNFLNTivR172Tv2sVQn5RcNeHJy4y2n4HnpDExu6aeynjOuF48gE
rf+41jJojkisPfZREiM8EF6Z5cGo2vZ4meAG/vzMmd3hO6+eqrcM/ASjKlwqc3Wh
rmHHOn0oD+lO5gkL2s/jhOzpv/L16eczDCZND43qPac=
`protect END_PROTECTED
