`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JN+ffwCbteGefnQS3NCOeVPwtxcUFsRsVVLylIYYKkl1SSD14sJpiZLhKYpfNEZt
cS2A48mBw9hrHKJlcrlPBCxFLTx3xBOblSkiRD623qi3zI+rIYPROFa4x59B1gHe
fdWxz8dO59EMcQko3w6/Hxy8pBL3rxBVwgorG8uE/GEkt6RM8q4rZeKdJYIBTAc7
jc6xMOEtxktMno12kiMVYzVkSk1yUwKOdxvtC6oIQvKEiUBsGNO1zlKkjkpPQcHg
Z0Zypp+g2mHugW+s5res5ldUNRz75XBiz+6UWIeujPnbl22OfeDmTU18rLjSff+k
PyjFSr1wcFZuftD+iOya7PvpaZ7Bzu25N5xFFrrt+OGI90Wjl3YBDe7v0A4CeOid
jpmHrhvv+jK1DV/y30TEpJWdU2XjCCe1+w06f/e8ZxRhKGjxHlSrcQ9thK97d82r
HATJFJCv+0gIOFnb8FtvOEAMjpKm5Yf13KSr7WLGQoXYtWT+jitZml3jYn0iJU2d
f3B8VAXy3s7FuNlZHZMn8QGRorXvwFUhOUO3yS7+Y7CBhIC9Yk7UqCBGWv25Qjmy
+PclpX4wnZQgBvjyRo1geMkcmKm0RtHb0V2AF19BJ+9KdyH4u6JCp+RxievHXhtV
YwivQoRjVL3NstGdYueoC6XD/LZUtgnx+iJOWw0mgSm66V5zCpnIC//fU70bC14a
YXUk8XLN2NRhE0iMT5iF9vhZdDMMwrJb6PUQ1Zy37Ru1qYk/L8KR89r5EOQeni7y
Ozg/UxYYSWUK8/HFRyK+oAZrAWxuOt8PbxwWHTt7ltTrombGW3v1/SnyVy2XKx1O
`protect END_PROTECTED
