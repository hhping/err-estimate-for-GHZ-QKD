`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjCFWucRZ+0iOSGVI5dgGaLqXUV4CRt52YqFx0sGANaSpulH0ggPtavRyqAdNI+9
CIPJTxGqIJ2vgM+ZyrqOGwIIeB44pZIib091HcK8WvKcVsUSU4QF8H5TN9RfMDWC
EO+9xOxM9JX48IkcRsYUS4Me/VIwaOKO+LbKtYJrsDxPNibzRTwCJo/LHih9BaKV
geu6MV5NsGKNIvXZbdS+r72mr+J1RH96dSn82WsGaS2q3m/dwq/4jX9kwWjM0M+W
p1i12XnVIO3pF3NCk/2XU0QmR/hYWeDpRy1fuZGCWmpPZEELsF0/x43u2MR8nl6+
pmj4AUfkrt4dAoczcSy+VBPkphMWNZdv9l0DPCtAxv9S+ClAJpmWt1NfwuoJCiH0
HUNaGhynFNlrujyraEt9A8vVUV/oyu+u8e93ZCGzbMaVw3EjB3a0qsI3O2eThbEd
pJSSExoDXt8hHshplPXboPozc8v3bmnuev6g5DMQCLEhMs1RuARTtoLHPVmVjmlj
rqnkyjhmQUZPJ1QQtUKoW1fJjTqcMqDq+GY+j0/DZyfZne4f/PwFFjDL3pWukmGR
+IKsSWaoCwNwFo7c+VyfLDj/3+MfK5IBMw1gqu8FF/IQF6J/58dHE6puZvlfIvm+
gx+qYwp6RmLtLcCFt5kdel3LAaEZDFCFtTZ811T1hRYUYgT0wBSi84dml4+gUv3C
yiH2rLgjsQKgCVImFfYOepTQBGP2fdWFmDmupTOG7+On53FbMJiFZwhQ44p2MIT3
/t1o6po/0sKNKXd8JXCNgUUWYRp+2p6MgIMX/+OBwhhBX5mL4VAYu76L3VtrGVbu
GQ/kNzfJSIRzC+rB30QcKRGltnyhm17EUqI+uKJ4jEdikIDSc4DiiFrjLzvIVA0P
CM0NzXx+HwrTJWDceV/ound0zlYFI4rU/UEUJ9D4SC8QFC3aiXl+eqvVikXeDhpM
q/xFyqAdu9fumLcWRn4euAIs0SNK0qUyYS/CGqFH0JCzprb8QZYqQ06zwQLg0hsQ
D0enAwrZ41e0CWFszrlsezhgvOoZ/6mtvvFshZLjgJJUwDulsfiQIl6nzKlMA0CK
hWf892SM4No0WbIMvXuOg+6b/HtSNs+GnwHcr2jNOQC9jKwwElfijTP3Prb4zIdV
ap4tTkRnG87wczItyL3sJzpEyXX3xgMgZ0Am1eNz5c3i+fb2LVmSSYnQMmcBXyrx
WAHD4p1+tOPE6ZT7KO188/pCChadZloBMXhvqkLlt66ZXrVvniU+4o1wBQT6Gbqf
aX91nfUwx6PNS1LyOS6wX/gSUhH2jsxTTmrcPJyIlL/0hkJcNVr+Fd7rg44WlzEz
+vv6kJL5mlCcRKed8gXDkt/iW0Q/Oz5ONo0LBPRJMkFq+Uf7v/rf/iNCxVzJs+EC
5czpC0kMFlb/fnyb2HbwN4Ry/1fZtXwrY6i6FVMltNNxCGakr1wdpSQZPoymCGYS
VR3bwIanTIYZPSkL5JgJnd+Xwd12KxdHFQtiN8/czwqwxfAoHFPXjwXW7/mkz5yJ
yLH/wEwkXsJLQS6jmhiUcePZ7d8tq/Y1B6mcTpZIIokrzzQ0q9oVAlTvb7KVv+/3
E9A0a/SuMWcaxOVaDNkoQmqMjPqdAeB3PDXcfZowCgzQWV3nrO1jWpuUZh2AkGik
fUQhO1OsMEiJoVgD0oFGbYRPFJQyGTNaJSBeifK3bCOjOI0470GXC7ApE7n+P99M
5ug5/zToG4/g6Yu9FO5rrUwEanwMdqZEeGLdACLz0+Jp+AyBOpapVLnjdzLdH+br
+/uxnURQMM1tO1skSihXQzqfkGr+7ReZ7+ShCfCpi6Xrc17QFb6E+UqYH3KgVP8T
YHfpw1jg7We8bM3SP3geIQbqMZ5VpRR80112XAvIySLqT7AlwtVJQNtdmTBy9fPj
lUplBDfRozWFcFu6+/VnXZgSDAa8h7o3Ydzbazm1Kuln1nqu61eH6E5wE9lHBMEL
YuiSNl8oRoQfA6vSIRVEKFmqRnJCyWaCbFT344KqtrielXNhGQtd4R/Q+63Xi3PI
Ip1SEiY5V9joVUQawHphv/DGt1ZJYcV9jjbrqXbu2VfjqjGRuxEl3PQiqf0MH8Ma
lgQQLlduLXTWQjjAnDNwnyQxonxQbFnl93ZrR5s/a/A0VyRt2Bux6KWorlAzo/Fz
MLsWn0yWcFIKV8ezoM4r1GRMs2n18LTfDeGXG6BPf/AWZU/dYdJ4p2ZZyXLEQNu5
s6TFMrypnkLNwunle0LzZ+UX0rxw264O0B7q4V0YZt2G52lXF9ibV5bPI5hr+cbA
AK4HDwnvYsgQvBpwOCzfclHt/HI9RLvox2Nf4BPntisBcS3jdJ1M6t3xDJa3E/kY
gTyd07JFXRnspSLZufsAKJ4YlECiISnOCfArIKf7hN8dURSjpTQ0ejG/lrE6H8xk
kxxYrljaMnav3fz5HbFPL746WOnyxWk0JvjKIBGC9NH48ZVkaOS47VkRnwv20EIT
8+jGCYa0UbqGOxVHiYxv6SzgI4KAi/JHmpAm7lUfDYH6HUFDqTkiI0iQ479bGEKU
ygj/zOC2ywwe+AWcpU7X3R2AcyuJRJr2Hg18cXBJpdGn0TvOtJ6amrMb8ioghxjd
BMHQYUQE7UtnEht/aEcytpnoDVBYP9KCcnQn5THKnpkL74N0rwpGJl9jRDgaTITO
3+xy8Q9UdnHMlxFDUi7jHCYT5d7w8yKxUe4JtPG5azJB0gENO+8+xcNbl4tRilLC
Fak9heXf65a5lxz+0aBIVc2OST0yPNH9UhikzdWyL/pRRBipBiImqDkW7RSfW3/s
qPaiDie9zE1kzbuqv13yAZlZ8wmc34zYVVoqQxCIGoaiZVo9sjy2yNxAm6tvgcjh
qlGZlLaYPTekAQOJ9Jjpgpz43yClVTxxEEnVxgYoXyduNXp5ZedbyBXms/ZSHr27
9IOF5u48N1jQ6ZnPiUQLWaAlaMpujqC5LKLJwoFuwVkItmw5mI8uPjSJPyCSnpYX
rsvwFi5rCYTg2LtuQF2g3aX247A4mKigwFdY1bjOHuIRb/GbpiDeHFUJSMwf+czb
CruTM2pu5kAEAS5Ng1aTqoBotpTskKhcjIkU428QQBUzNChnK9F3O6ennyFJInNM
mspKT47wcPI6Cl1aeThQSx+2cfC/fMlZ9fzBXu92Oo61uOvIVZkFtUsqimrdFH7K
aNYgei4Cn+SqUgmtULHol+9Mcql5gR4MAfySlqAAwijJGvMWsjwDfvT7FLtgHOMj
uhIoQU9Ofy76X9QFz9XjCbQ3idozbxWv+0n8qL0PHDLirKjb57mOxhEO8j+HwENg
HTPoq/j+GExFi5Lmtg4lvNd5pQUPebJ9uL02983o6L2Nc3HMXFdpmoaQQHAJroTU
VCJFw9vlVU1wiBf2b1d0var7Pl+jWlzYI2yhsDHO/OGXnSqZHQLfenXctW1Ke7Qa
2dcG/04fvtp1K+NmXQPJOp3RCZq2FvyL6GUfhoFgw3A4F/st1H+ZWf13thuYbpPu
oE8zDRTsl3agmx7yFrufPw7GTPsvxaAwcM2YGA9V7lnztObewLmogZA6sP/PonPV
+2e15wVXD1y/5MZvPg9Hn85M46Rshmw3f9ir+TMyVLwrGiq5VUXNAKNmx+GpVkzs
y3fhagzohknqOT5mAZGWSeiDTQmwf/Mu57b2cfb0HsT/n6DV5ut/Iq5lQq37svtL
i82p8N2f823BGhp3WJUrI9Ink7hwtTZpxpY3cKjQZSMauM4c2EWOv9NkF392ISDL
V4CbYHYE3CjWEI/JKc2f9S5SH3z6FjUXkny3zqqARSKw9zqBdNnTi3bqyQ++hDj9
26Ct7w8OTvBX6/mkIMBcm+u7cjNsnOMWDvj9XRRxsL//aHkebR4CbvPHcVJxmrQj
8o1J3dI1p7PgTpQN8H+OOkHeVIvm2ZC4xbOqtzt8EKOYMmvEUM3cgNuou4nB4yr2
n04rukCvysyOXaLoFC/rBTfE6gqVCjpmo4wp7jJc5iZCHbN74e3oyxD3pi0vXab7
WVcs4T278U53IseFboM9LTNa3FSmlIjjO0Mz3FLUMXQZAgo5m5XqgENGqv7laqLD
1dxxd0+dHcrVoGCwPOZsNOL3GuaRPAnS5ybkBNQn0B82/wDZDYSEyDDjreH8/vjj
XL3RAqq4ZB5smhrysQK3up87gHo/J8bEnS3X5MOtmU4iWrn4Lia87fE/E1LYN1am
eesmzLTh442JYMCZLMo4yq1/zjwY7QFwLCG6ALwqeVQRPeOQhPHxeQQ9X59wkTrd
Nb0IQoNO7yFiV1VAmX3VWov4IF/qHW8g/npJX6INbrwYa4WxBEZ0uUqqb7EzoQdT
nHjdXFoayt9wuIGtyP5wtOYo8dRw62MRc8Rv0WLhrJosEfraxaPX8v3EtYlRpU7g
doAK2Gvaw/nXtCiduUN1T+Sji+1910IiblWb4PX/5taKmusNJlmepz+W4FGqOw8a
GH5fjQaWv6H7qOJiukmK+9luXqp0ZSG80QwEHwyXid0b4Ca+QKjDlUM8ZtmYGKNQ
U1oUbE3wvT4xjeTT5V9qF32GzF0OyUByXUxee5ekjYs57q5ll8dkqRifN6B/WMGh
++fNcA0Lm6eaBjOfCkhwvVJlZmWvAwMvRIOV8cGN0bMoLtDnLhR/0WJVDS1UbdXR
A6lHexj5I/JmHTslJwv5y1RSo+cl1HGsAcC0+i9BZMFtR90Kd7PYTWc1YDWLguB+
DKTinmX9j28xcxtMHnjUHcud4IDMPMY7j+fzsrwS1J/h3VP+sw5ucBsc3lZ0/y+m
0pZkbXNs+jHoOJiNrO1C0WuiS81/Llj39zEUpJIkiCieAwGx0lzbGNFFk7RSCCGM
VMccPxfBv8nXoBYyvEu6pLxkqNxdUDiwQYikFcXskBKMtrWDrDDlGhcixvVZH1gu
YjOO2vk5QzTHeSU9MsqjeE85oBnwp1j8pbgYHzC/5tmZCjOL3anOq1a1wLslCKLj
3JQxhj3hHxnO2SvcoDsBHCKMiPgDE7SV6LRpv3yiKj1xE1C1KHs24/gW0mKDEzGO
m3xyX/mZa91rD/U0fkVQYg48QH9o4ipLxi0G7H9ig54XPYYRK32AHiwAwIklHs4c
ciUYYcqG5YVaN39+wLA70Y61hDAHhmR9jdA42MdVO5F2xxjO79sJf2TIQxv10vq1
LJznePoDnfOd1lLIiZ+Ms09Vr0UlzewUnEImVY/6CdK6312A0NTuvsfY/1+UZL1H
S8MYVAOt9uM6HG87/hi3t0Qoq2jjJI07dm7NfCZS/A2zdYX24Q990UoQ8DMaLEM/
bTrDlmD0zUvFWJYK88uqfK2D9zWBc1BpeaT4VVro77iH+sbmu3A7S5Xbw0t4RcV2
PjcauG31Re6C2uWyDWs6R0H0G7avklwsYDic9SXgkzJzP4iBoSAnnzZXvYQXYosc
A4C9KazD/kc3C/gkAfmarmgak9rdagdKVEBn3HrZCMVsac8yUUL7EKIYLL9a4DEt
tChO1iBV+/xDNVdCmyCZeVH2XLbDC7esFj1GAWpRMJ03GOr74bIOYuFJ8AjtfHbs
HtAlow/aV0QXovEWt45MrQhbfRjM3PC2ynUKMzXmYplaKHC6RgPotFbdE2IQRvF3
ZT8g1WpHuG4tClyB0odcSHqENxrjkLPhKuiPBkBMcK+0tZ2OL0UNFtS+3TiriXr7
W0QggrNXQ0RyF140O8ksGSvn2WdRehQzppglABcsSAy+wtBqiIOq/IWvjiofgcu+
9eOy3ypZwnVyReRk3wEwCkzBfPkdHUki3Snt65sLJe1S4eNVpuTA/Oup8F0Qk2k8
4truixMxa7d/OvF10YyXNKtSbywsT3OxdfCxjD/HKuOmXexa5TFBCa9yvXhkwYrD
mDO3xlcX7gQkl+6DfdjjsBhr8WXFcHLehQW6mGCxnVH3zrkHV0Pw3u9B1Q6m04Om
NJcgzlLzYC+h3fOVDNZY01XSgkWPmgvivn4xhcyKo/TnT2Slk+wKkMLzCebFfjk0
qmPM/uIu02IgmIAsmvMS9O4d3jN/aarQOjZ9o5MzcMo7WRMc/F/w6vcbCCjMn68D
2DnwDcDw/GUW8MoDEET6ZzxkDS6OMZkbIpx/dTtKLx0GuEspgi7uT+DkHKsmapNr
6AAESa99dnMMZFWMsdV1d8XbtikV5RaQplhWANUYbKzcM8jNu+p/VP7OFl1YAAK5
fQl11FGFWlq/KklGcRXvwUAyozrwfRlZza98Vi4V9Lz6RKjY10GhuryBTg82ivVn
vqNmcgEHWV4EO6b7Wlv/TMIc+IQQIFwoN4UjBrnEsqToZDkcN9LVdn1HHG3CqyKA
zgoec4TGAWntX2RDjTvtADn0oktIMt5VC52qa0UZsPuGhnDQGhdREZKOZjKh/xZ1
Q3TfsRO+jlP/ijAAuUey3RQoSkcDm+mbhRFoBdlVv9x8DwGi4zjl2UGOgH3Bd0vn
etpNGm9UPtMpvRpNdEB8HBBaYCMAziJCrimsw7ORvgRO/HC4R8O6fwzRlUjYvW1E
/pU8bBTpG8x+Q/lNIARLQVv737Tl1VM5wyfo5ENPMydoi4LXeMxVgyTfxVj5dduJ
5CbtPC0rTo0hmUqMbtUVLGhB7QhndfKbAp1vU6soq1ch3n6/Krr0BJcY4mDfwjKR
DvVbTEp9E1Z/kB0aR8DonzUMs1Ldrn5A7oNVTqLAlqTWn+R2H1uSTPJ3u3qpkehe
ZyD9bbzwUREw/BwGHBLZrLY06y8NUpxhJGEeGACksEmCUBZssxMIfKKH3HnUTejs
YXvMyOB0Qxi80PZ1he6zUVu+8p2pFKjpK3eBjLtPR49WJHypUY7/xTqL5aaxL0o4
gSMvVineF8UvqZb0/41FiRhv+3N9PaVstAlH3GB92VjQoO3XCR0BjlwHTqufhhF2
1KMV7Qifpf0OBCoQ5+e8mYgHc3HQ2/vceVTv98v2uf6/vMYGI0HzIqEERJ9v0FhP
VU6I3GSnNXBTfGfdmHe1mK/Ex9XliGhR49NlsjF/hrbxdU7oxcHQeEujITt7V1hT
hmvnhKA5XhJ9x5HXyA2xmWEbiWuQnb1NleXgmaDwQHyOYHsMYWZw/09qDkw6s4TK
KpMyDG20pcJX902vSAkXefVt+Y27k6tffpElxWVuKyHS+02v0csGSUoNOZyZnYpR
2svcOrkVM2ItRe5Y64iB3nUVCZmAPGCY+DSXrzC6k5OJ61rIt15/YlfLW8XDi8JI
c9zMvimwn0fg7RV7fZzk8QkWuHQSbxwYiD3Y8OKArAY7/IUEWw+fzUcSGKhOr+Ws
tcmPVZ3MPDy0NFv3t3Jq6p7oqVMv215Fwv0Kl1yyHQOASvVe3xyJipBR9yekKMde
gyRTL1tuRY9g3wy7KrJaiiaKkYFFn3qW9a4SRpd3hzGV22MyheidnWRWsUOq85Sg
uvsFZWhNYQZ7J71WUeDBnpj3/W0QWrfi7WkWvu7vYGzGVkdSlcp/e65x90UhsKbK
c9ykajPygNhjnSFxC4OdJsvviYkUkxR9nAVJZgnYVV8qWbSwHP9Dm+31jGPVAxDn
QCM2dPL/m1k4CJ0RD8w3AGxkQWXXb7xpr2Vw6pjJmwPd7QMtm0irjuH/kP4nnWMV
CxhUcjXo4Q7txPmt59QUPA==
`protect END_PROTECTED
