`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggBp6aBvcLJsoRcnhD/9FVmN/23a0vJOrbE987Iy2rt9xVZow42/A5l6qH5xvGqI
dognIxnugaWYyr6k/CH8cBs3Bkn0UsNl7ljZj/xwtraMB0WX2gSJVTkedMI9LZXL
7H3Mui0q2XxV5lH6s3hfHbcLnGf9TKKW/2BV8UOcIvIJ5gC4YXoDkSu9Ocjp1iOE
zXQewf0TU16b8Ph29N+PWpYucmFIwlvLmtBAI1bcyk9uLg0RLAcY3I2DL7xbZPWz
NPSiDlXVenKJMWb3alTUbpHbP3qpogo/xPiRlNmbbA3ZnDckLliQPKxgUc2HXkqK
ZadAqFaX2FDhJ/TLP+If/YcQ4IIB56NRivRau0pu3V1A+JdK8wMpmY+6qusQdvh0
z5u2ZgQW641SkQG8ZX6WVaDF4ZYb9sxbCrSu2uZmn+gLrG7F1Fp4Oa70f7QxGrlg
2x80dm/3mzaHpZE7QIgKBqu+HQOsk5Z+5syXzhgAMzNunojlUZE/rtmBDjKfhnOZ
OiCv57powrxMo3fY0ni/i5dIldNJ3eNi7VsLJc4Zw+5DmkOv5Zph70z67p56xAvz
OEchnE7fsz6CZYUM3jybbpWrXdAzdJyDWhAuS3xyatpaXxg/Kv7D2qhzzE+BBkCC
CMTjb38Lt+IKYYCoKtkivJZaZPLlpTQTVnOxgLtlsR6KqW35r8h7ZymdcBvKfRPf
/qaW9arnwAOQoaygKzV7WyP4G0u24UmGZjqcGTPizUtRgkOOLDGqqG629LxWAx+D
KjRcXy0YYUHG2/3CNw9lOBj5pRN29I7y6QkpDLwN7Fn3/lDyvz0mWTIR8jHuFiFv
g2kzQYHPi6a5ZeINLyHD6lzWAh+fpeSAXPe/tTilAZrNPZOjbWnSZh0byf3qaU5C
f2er/wt8a2IxQ1K3cUrJLApKpg4hoiAj05Iux4Y7Oxgona4C8OdlupxI1LwcYBHa
ODL28jer2SJj0Rd5OPF4y/5LlTPpKT6+azrWGvxJJkr5qOqafA4b+FSVsxoNlA8Z
pu3SyInw7CmGOCE656ytyrewfWv4MhsjvobgTCQ6qh2SKlVdTI2+mvQxGXrO24yN
ut9uvQYptFJslPAiJdV6msHUjnCh+CAC0iRxHJ/MQDxUiATNUWgSWwCbyWjZJFVm
dNEMLb98UZeO0Y/JLEM0gL6/XialmB3I+ZO2iBSz60iusgRXV+RiWwO9ORV6bvep
EAD46yeyUaxt14vxk39QBiXUWWMakDJvBltLawGdrj5ZAYvqAjJQuPWWpkgqTQTW
RjMshLAnThZcFfqfPe/nG28LYp3b23CMn+I/AlZLJd1wpAxbOIci6go2WVNUj4jX
jwmTL7+Anwuhswu3amTy4NrRRbmSZ9niZ449LKzeWYilf0gZR7bMVEBbUnThpzI/
PizwUemyJQBwvrZUAEFhCJP3EJd7D0mpi2txoSok+82mY6bNGsuxyJDWG/03JkaE
sArhxrLJ+fU6l1oYAeds7HkmfRwuXLKQwVWiJFQGARPDl3WNxYbK4lj0aswOglQ1
5dWj4qTduckrZC9DezgZyjqFIIlRbdjKd1FB1iMtssQaSX0xvDMVog/InfFBpiiz
ilkc2l5OqEmHuhSgPDbZnDBRp2aQcpKMRJ73PfZQWqdB+9/mRWVDT5tdqDqGktwZ
m4QJHoE948OLOsPHCDCgH33m+k/J3BCDTYN7UVnLqHKGmB1kojc8lXTRqhtrhbq/
O+uoHZzRGKLv5BnPXICqk0KWovtt1pozmma9xs2GibtkwdwkhkjmJ9cgf/1dVCDj
De2ULJZQV0zTLVxX25/B9ZL6n1PKCQT7Ii8GGCdwlXi+erctuhyYKxJ57hlNeZFA
FMEBfpiEGxRzM/HhtHzBqxC007QYKEE6NmhExz5qPhT+JlleEFzhz7SOlgFO2ZFU
k29gx0xK3RiN09/B5Ae4Jd/AyTwV6FtnLbR+PgUmnXf1KgrZdtNOzOZxFbD0uVnI
YecjNVIdUPVBqjI3BB1F68q3NAZc69mGMqZslCywlu0to1qgNO43Q11hfPoogci7
v/x6OEOT1SgG3wwxp3NoTFZ05Vg1JSEqSVfCSSZKPnLlGPeSPHN71ssmTt1Jx08V
75JKEXWaOmqluZqjIPtjJqCnWgAtkqbdbNETHWhQ1IVKUz10Cd9Ar5gHs5Zw5lLD
oOevY5pfknHIpIzRu31g5A==
`protect END_PROTECTED
