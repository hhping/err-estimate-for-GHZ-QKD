`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWl0u+x0JaR9KrP314fz51gVDl0pyl0NN0ZBRkVHLxoj0xEX8XqTManDzv4MSCQe
hp2YPHfALt8KN1ntr1dkOpJ0SudPDWtuBgFKJ/6JC6QFk1Ppc6Gy2OESyAcYykjy
E8T6mAwegHKnmPaXYAY03urS/yKH1ba1m15Hli6Nx9OIPcPYukavyni0AcicIeAA
9sjZOms32LlgFyduubyjwb87xtSVa95FpKAS4tGnJDbRoJCvbk7E6T1hyklhYvz8
w1co4b4w9/6y5/x6IKf3sHwhrkvjhq491abJYHR+I51kele4YCe8Xgu0BFRjbDD9
V+ZHMTXDiLn9qNq8oJ5aJyIikveakqSe7N9sqfmy1tMGosbm8i61WsDGnIQvr71W
qTc7um8YXyu8JZS95VEXTzpaFA3jsRE1Sq6bgWwYfwXLpuhBFhyS1IuIWZEiyroi
OdRU31VF8nqOOr6dyLbOyi9nX5EJ0g+5qwxaAaOFBkmyW2ZDU1PVb7eCung7Ku1D
g5YHKqMtsyZ7kP/wNK3SKkjmpP77m6vMUYEwm6s4UUntYuw/mL6+N5kUsdcC7vh4
nrSJGPpRBWlgcacGx4mlnyyiR6VSl7O6uz0wPH/K3CYZ2rZWekAH4MQH4dxFYGnD
eBCBp9GulF5lbBzP5K1aGMFor/Iq7gXEOBrpzDltTMY6dgiTeMVE3MjBxK3m4Xu1
Ain1PsID/SzY5CP4DCEvzuGh+Dsgg3mDAlR1e7dkXIOHNQcwGO3fqmLPoOALCXrS
np+QXr5j872L8nuMZsY5sG3/02lnAB5oiIlRkjnHLeWpA3b84OdFFB9J8gj6+qwr
ASrLtYTwrrOtukGwcGCTMXD+kCZlNwsCJkhjRDlzUYguONHo5QJDX8hZcQERgsPJ
KU6vipyUeoSJyjYYvXpg9m5Qj1F3O485yiGy39BGYGPF99IJlu6rpOjhcjdDKehc
kZUmtMER81fUTMKP3lH0jlBt3dsAEfYpwJoRwNqKXPSNOAAPHfS88J5l4kuqd4sK
CXIyeiocKDY39hG6myceZhPPt9FtBid8q/M4WhcqQGWsupHWCNO6bh07ixloBE7M
EK5wIqwdXpLOZvsFxJKMwwz29rdYIuQfvFPhZV/AxgONG59CoDWd9HNzZ0NF5yah
LBIfjwax5MYAadqHnywEFevu3a2RQ2DUNBefQxHzQ+SatqdDzrLWWUwFY+o8y2sq
fapDuVmBvDDsSIYVgOe3qO19OP2bd7FDWj6xVvdEA2ir+36jLH/XpLJeH7WmM7oY
Osjrg1rpp3TD8nMCIqdeOvmUP53BKWiEpNhNNtcy2Rx7u8M3gDPq+HgLT6T+SWKC
caaRTh2rp2t6CG8CY3KQZpZK/c7NcSosttGQmXGuSYxEeUOkJ0zu8KzBEhfeXmhY
t/CVxNJxVJXreApaWh4RWhyErhZ1BamEaUJyvfyGIoICbBcyQzXlrwFLknDluYk9
DlOCPAhKgMD/Itd4J7Rj1hOkU+DAU0+f2uU5eFtvejpT31stBQ1UGXoCfFAid5ab
T/K47Kki1x/j0qwx51XcW9rkxfD6ctS1rX75nAma3VraVymx7Ps/Jkg0bZs1mwtX
hw++ZLjcs77zQKhLjWFkYt8eCKay9SXAUz9LHTtDrJ+twyTugF44X+X04uiP800i
OgZT5LnXjLOgxv4+xnCU7UNjgu5XvdElR6/5cOKXNCkpAaKRe9pnjrTBkZXFq6+N
SFmbmAxkNdCyeqHUTQ964T8eQJXxEUvXpCViHcrFrquWsUi4KKajwsf9d8DPR8dn
pxF7iKN0QRmqOLG2SgoAtmqOcwvW0F8xsVIcHQOQjzOxbgrWIt7H7cfZ9POBM1MX
p9K6r+nX5TrKsEoG+n5GeM8xP/lO0vfCl+N2gxJtD/bsztUk5K1XaXrDKY1XGSgW
7FE2hK4cFU2m7CKmNQr55A5c8Ht0JlHwPqY+8G1hJvrogHNvMvUgg2nVExGPZx0g
wiAHt9YAMmESw6E5NJgkWpsAVwFiRs9FbzIwuPBuezTasB4q+VeC5VkpclSqG9GL
sqil7MZK1FcTF9cMxbPzMsfskYz0HZb0RPmQCYa+tUbM1qPP2GWFxS0YdyUp8QQR
P8ihHdRJymr+ZwST3NABQL47AAOR35O9ESQ1JzBk2r1PVem07ePkuduqpsmIqrbn
ZW74Rpaq7wnPULWblTjpweqheLiqmP6d7NEC9I/VIdQKKn8jHthcIMiupyuJ9+Ah
JWVOtmYl3NK4kywaQLThJo3wgj2UFGW9SrSLDzoJL8HBqPRYTLVujukuK5Mp7ahh
Pxd9O4pmUEzr+04GijnDqgR/ZWJsuF7vXJFTxgPqJIkzAmbk3exkpiIJvcgs72Ln
2EfxTeUqnurmH759dzadLbgvMM9UKp446+wOFAiYxUhg4fhm2ovvV87UfrAF1vri
fMyBgpT7U/OMsK01kVMgUbdYxCgi4yFf6XAVg786sZYwtvVv9evog6/V5fO9k9ZQ
N0gILjRf38Yeg0dK+i55oZNYMyaHBPTgW4cP0fVcmFEo7YDmpQv/gtpQe0l75GmX
Y6m1d6JfFz4YmcLEec3cOPFTWrK3wu1d9npPCC5Mfv/kFXb0yqxgC+QJPaQw2wQx
/9ckRro5JXZdLydXtB8g8VAmxHa8vfoioeob3KEN/qQsFxWIO9MJr8f6AH4ZSKP/
/wzRIm7OQcfly81tqXtVH42gLTJ4PVLlyc5V5LR/J0RjIrwnVBEggiMSDke7Q0Or
/Mz/AmPBMeyl0bbuEtH7XruIqO9LZHcPV3PI/9qYmFXzc3ZdqAQ+zNOpXfyAqy10
s8+yijZFj0Kf2ZKjfo3z8BeblwL4it8rIYe+ekbkP+9a82W8uhLXvy5VK0GZVmCh
s9082PT+G5FyiSAJ8h1tTQwAqqrkj5YS4qC4HMzms6LE+eZj5ZKTea5txz8gnM7W
oie+nqrVyu7uE5QJ7N/SxQc8o2hEZaifa5Qjap2WP/PLxVXMju8IAAYdh/r5s+gs
iKekq9Yfe+N41hZXCfnCcr7I37DyADGwc2oZJK4TIpAfTjIKci2rlPFeTl9tB+DZ
ILSLrEe0dgQg+WYqT2BSCl9/fzy8ddwcVf/RxKasghz+yNttnimtKkdzpAADv5ZC
JcrFpIm7gpm8U49gN4We0R5f8ZRkp+c87uztw3uKtYfXji79l52cufE3vB724FWH
gVvS0LlKq9Ymh6rg2cFjUdodKke/U5Vpo4Tn68+0IlFkdiSsxnx1/jFTKvIpioPA
cLSxfU6/DiCTiLPNN4pNirklc9K9UHxNzQE1rDmBUNh/lV2A5nTzxVp1dn2zU3N9
szsaM9EtvQ0q203J17NPNdizCTEjpw7r2XwWXNktSoAV1vD5d4ghYQMBOk1OX9Ky
aZF8dPkHU4vCk0X0BRELjxmlwU+a38AITcsflcBpA8pFv+L6pT9WdOzeCNvI495R
8FOiwOn0rg5Ef87s4/k462GZs+NbVCU/aL2rg53eNks4I4/2F6YTXzJ2VCCcuu8t
PyZPTqZRXq9VeUt+Pj3ClcTDOAVonERegZX+hxa5UZDDi2iwn8RaqGmVKaiS59tU
xKEvBRenVApSXXv3slgd0puIA1dCLju2IxUPsUx4RTzNxDjVlHxTDqgP6qXQrss1
hFN2ar6eXLBpl2SBqAh1FvY3goWGo7xCWW5F5Qs8A92dHHTc03g3jbpNiEIF+CNh
h7xKS3Q+xZeyI6RiOvy3HR+3YH1+hzrvl6g65JY8FiU6bYKs72CrOE00mvXCsfrB
xgu6tPDIf32cjJ3Y4w7F0Gtafgbzr9mOXOd6U6Z9FXffrCG+cZZ6OOAOKrxf2VKY
Rd8x/VpDCdMxD3euyNJeM7yiPgWouIggt+/LBiinsIrwLm8E+ZEWQ9SklgI441gQ
GTp8gSjVovkzd912Y7Op8GpZW0iQnPSiA6C+wLic5x1D/Un6SaTI3MVDeyd4ma5p
YUCVs4I1HtF9SeVDKdfAUbh3ZCF7rrEEod5PPznYz/S2cA6uTnKnXbJUdjPwNWtt
nssqKqkyEl7Njt5P2N4Ov4mCCGZHy865O/3QLKZj07M9MuPGb9VbUgaMMIPHe90X
vvwqRUvyD2exJ7yRccMZtImh66rJgJl2t5x32nVDT30HV2FdORwJ1z2kifcrOCFD
PJaXtWSAbuOJFJt2Z0dMlN7xWUHokvHkIOPA4+3+oFbBtI78NIOc1AtkWBEyeQpV
V5OrsN0T/ATqWz6h9oFtmuWj+JHagpXAqPaCPmnidMuC31c6D9jruZIE2+O7THI4
NgTHtRNVx459yyHINpsdQnamC0v9lWmN1BFADfpmr9QbEuPa0Y3Y69tf9z206skr
f49EsqLfbhL0P9H2Rbw8a7GzdQ2LWDMMKzP9GYVBoUT09D/p2d6sNO4xKob3FvzT
ptI3+rMS0YZ9ye4PE3liHxdXnuLjtG6V0Eg+gBvdMONf4DyUrA/vyS5r+57skhxg
7TvIbYsCw3lURrflc+wPIjXC+pDpD2KcqJKSbJFlaQ2RXHIOju7U6oIIqLmQvkIO
QtVe4s++Y3U+wU5jJtx3wIFmU7Q34MIHekfSohdf3u3KZL97I10YNOlyt/4ZjqsT
Lht2HMLI+c/dcjtROo7u/FM8Qfv2hbZGPZKtxWGKXR8m6MJRd8mzpaW80qWgYGIw
vWIYlCYZ2/7lU74svZn11YJ4DIJqA/AFsvXjyTpsn/U6tDBj5riB/nkLFMfbVfr8
jQFYfNtdGoGALHTEmPaRrZ+NuMlSBskq4n0XDNREW3uFH6KTn/reCYBcyrqJpnrn
0xkefQOYVD5ZQ7qyKb0h3vBrsnImYPPwMXUvGTl69IQI4qqkV2itHeez0DjGnJvw
SOq3dCPGXcz37hkz+A9bdPu3zEXqgE64jjiCgxk01g0xellTP8vl+WRvcqm7EytO
wzVdCXWPOwI17+7rymOZbh88rTXDP2XVBVVhgpKOoM9EyFMbn4d9J9wNP7qrH2gI
0uU7ylFPv5rkynkn4pGqWbwKuTWGLHCL5hFosx1cicQJEXw11ZUZu+6qwkP6lwnV
6idy6hxmk2vtEzAwGTv9B74VZsP8QFMEsaTwfb8AffN00jP1Z9uUmfrF3f32JATT
4xxjxkaIVi/t6QMPouyBwaq7tao2ChUV3IIdorQzyCaN8m7DsMdXC+QSZq0hMlVo
EXvaolUadhbmmEuGfLlJU230bW51aMZ0ahl10HxRSIJd28xTyeenSt8XziqSbll2
Zbyw1VncGHzs5VqmwwElNK/Msq5Yf8A8utVFpVBPnPPkc1QkYKji3Fi0SE9rECom
ahQhdfDrGUIGrzydAQ4I6nhiIfVGRt6Fbnsp5b6DE1tcVnp+LUN8QRZwMkLTejm6
KTqJTdyzRyi5P+35WuZG0XqvcxD+fKhKv0Wgp6K2TwStZj+Zk6VtY4lax8Mh5FGO
MZCVHRTtBDYrqnrHRfKJb0iVA6c0pdF89I9YH/U0AMnln6U6YJpnBWIgDnCqNRHk
uKkoJrMUbTjXFCwZGsxx7bQERTIsqCKy/2MVLtXBKLfX040vfzL1hdnQD7ndkTen
FHMjRx6D4zy3NpZIIozS+Op65ivOJIAnxhbWDCQLRwqIzmEtkUq+hMibyNlA8dW9
qkBUpBl6t7gsZi1fTMhGcahtAXbXZEP9/ifXmKmvWbL8s4dOaQNyDds914uXd5q8
uDw+mM+0xDm4MBB0FFeoiBfAEpCcVH2CtE9bP145GKnuLvJ8Bd7oPkt7IHRFirC1
2WVC7G7vIq0jU3arD3qiJVL7b9NWSHYEE18A7rzabwKrw+1CUh6hq68E8nD310Yg
cq4zmV90a/6mfbyL7fyNe42al0qaTamVVewvsFWALX6o8Ws45eETEvoubKXCzeq2
rEuZmx74MrToTAumEbgPOKR4BieUELAJh7ikp8UwAxKEjo4XvA70lz/3BlE0H0jP
i/XxY4a3QD3waXQIpaJP4Ad/SzZ5WDBhu4YwWlJOlrpUfL7XsXvadbp0TZ1bpRVe
QroSCBnnYMnx5SlL/iM283Ttv8Ic2OQHw9/TNGE7Jp8uHT8Xyj8bbFbJRhvaNtjZ
/HlA+OLR93OoO3ZicpFMeRux4X1OEAgC33r5HKTFH/5eW2d8rpie2UMOlhdbeYaS
yV4gmS/IFWwryMPns8W8QIwq/jyPDOwg8FVweaIfJxHQkXIw+79ac0pG9k8K3o5l
vbVDH2YT6Kqk8FztREMdaDXDnxKsV5JUqNtxPsVHU6UZwIQlEeWaTQ/bGsucA8t2
G/3PEkiwawxTEh2PJFdij134ebp5Q3LaY8enKPzYkoGCZSWQtLBdu7ND7Da1xnKs
Z3Ecm2PapPKTd1sGP1L04raTC1hWJvTpEQUMVNgjeTlInXUEyG5VeMdGdO9uKgTl
5Io6ToAsvby9ALCK/AO0J7rKBVjWL48/Kx18TBFdREx/xSD40wLKenuU8rpK82kD
qLrb3/Gw/H9UfVbPEF9MeWPutPv/L561kGOdtEVPipUq6Qoiv0xtX71DRquIAYHx
lC0RSbodJ+FufVZolCG0yOf7Xqvfqx2j7prySptByT0cztE+MDcgTxkqJkSWvPzj
UOy5hIcBzohUfXq6U6S90P6/Qqi+No9MQWis9NADevrhzYrLz2aBySNnDc1GlRLO
5phAU8ZGhffft7yckj01m/S4QRI608kc9T6wC6HJkZV8qKCKyXrefI/F8XZpw3z8
2EZWWnbj4apCen92gDor+btfjmlRQi8JdDvc0YsdiUWhk/SEQ2QEETBP6eUQUPB4
Y2HgJX+YqcNACld3A7itaXQ5fFoFFcU+Z/C860hEtslwE5bTYMb0ekhzdJTEIgKK
e/jo+OK4332hS5W4c80d5UlICBk6cJuooQG9q3bicsBwehNBFMzERANqcLSSTOYq
7uJVhj5R3FZ1bRqRcFqX0yJECpc3R2jxm74kKy1O19qRpPKkGLH7tSIfzlZSR3Yi
4YpmiJWfGtO0kafOgNl9e+gga7FyKP0w2xBDFXrkV3NI++CMq77GctkjpH/C+xp6
Y0phjFfz2MXT+BreY/vNkyRZZoYapBSHh5TkyaXTeLxyASYIyFJeXjUnTu+8lbvy
44pa0GfyJrWJgv0JCUXqcGuY8EO/nkUEFHDzzHSTwhbaRjzvwX+8kSlDioZdmRPB
ryMdAN1CJZbQwLQ9WSjOun0SyKxMR7I8DR2MUVBMQ9/3OLCnRvDz25gfnprQq9kO
rgQVFocRM61+e8229kjuJIqaeINO15kVnYk7n7lW3vPjxrSCyv8+1nM8DeRdVF9p
P7Z/hjd+NbKg3oDdblkoUjMfE84fXLsGgiBm4bSWeSHbE2S4jeyBtuiLzjq8BQoc
SJkfR363kUyT77w012fRzJ5U0UpyxE4ABqDIy3xPFQ43SZiZkcHB4pYhDPH7wLxT
aHznSxEXWO4/A9JzH0TrwIDQ1qFhPJpuKYMAnKuPpDLPCZqIaYiVAyMvxsZ1EoUf
aUh1YtxjXQVwAOmlK7t3+gXqZfljrTrV7r3S8XgInisL/EpdqX9JrfG0eJ6rtf/s
FQhzDSSo3o/hwxx9cueu04YPLvs6GFGHm/xEbaAyRcGtWV4yZ812fzArwAnQxQp0
QGiWUo6U/cZ49mXf01SLiI+Kjpuqh80mLn3pQbIM7CufyJG2pUMm+EE+dmVccaXN
Y3jb9xlTAQRFLuM5jS9KB15UNT0adA8VggmXqU/BjzcjuPYUWwIGb/bjGcl6Ljdi
GsZRkdJrwcKKGY0p429HsOqzun8lh2ULMzq+rlNZKe4BlsIbz87++GwCOAsWNeKm
IrhqsFwgL2czo+qYeUtYWziPtfAqh/gKk7/SWkSHe5LVD/wo0R180V3SF4jW9V0y
fVfwOPqckKV0baL6EPds+cVhvYQUqV/09KD91Usz/ycdILPpX813NLd1MTJCGdos
BBM+jMBoZsfUImtLu2GAQ86rFNv4hTky9GVbO+T1RzawcYp39ffzHXH3BBQ7hwkO
E6KEf0Rl9hwQdoEmxvh1oYrnakEiY+9xIsG8FJaFKm28GA7lpRn/N+NLed+mIoX6
KfBH+wh53XVCu+o5WbMWuP9mdufocvWU9rAE920UnzpsnieLiZ7WLdvFk7n4T2CD
B0WdUMiLpqEjnpYL9vgbM5+A5fJ9a1tdA2ZdHmRV2S53jFsgGxYnvpHR7FdTh5I3
VwlHhp26ASyLoP/E89ipjlwFhEeHgPQVr/VMNhz8ot6u5108dI6mjQ1nQNc3rSja
oJjH7oDnMeMs0gdWQnioPH1dpI08aNdAqwcTPJ33DJZDOspyPQCEIBLH+IhfwRQw
E1Q3/gn5HGKsCua8veEwjq19u5T57bpkolwm/hkUTv4G3QX+lQy3kBnFX4sKd9OX
qh1+zKDXfIdZ1hFHa1uzgnrrawTDI0eJ/bNoLjfbzqTkVWXdsqvFWRm3V/TkLs+W
MH3AkipZbG+ukZbQlqLTsBqxakgvCmLzyv2CH62FDxiE8Lw2nQdIQuuWhNZ1a72u
5Ob5dBtmdg1OsPknNxa/16gOp+iBZAJ8z9BcOjaixEGJD2NYPMcyCvnDYgmE2P5O
ml+ZJfHt60dtbSX0NN4rzobDcUPqTNEBp9M1WXa8aVJ3pneDScMPsXCQ8hqYd120
VO5dKdPtL1EAV/OBfDRkXLxZCDpLVRzjO1yXcq0smNp8tKmFraZrSl8Kqe157TH/
xQUI3RYM+TS5IJLdY79RhwuLGhbVXOxhEkA+iq1EPrUDqhMy8+lVfygd4kxBSXY5
pZ/AZ0fQMrmiCvpY1RuggIB8uDy63ym6N67KtK0rvqzp6GRIO65cpNdfLytfXjlA
aaqxwLzrnlgZfUHphgx8fvS9x/NbSynDXKbs6Mfo5gp28/FthWKjl7TEsi9q8/zn
cw3tqDS1hUtI1gwyTenM0NM6fKlKsW9IS/EBG/tUubTuUoEojhNQG2o+YJSY8h4O
gNTP7SN16kzbI2iypW70HU4mAfdhgmiRX+q/FLZRbJ+HCJmQrDsSfEVPrWBkkEyN
BUQYVKcn0xQYZBMyNbr0Lgkc98ZseBD7W4vNWcpCCDZBBP+7MC1PcNyIaloPqC18
mrlofH3LR6PIfjqBf98PS9KiLSmt7Yt8/aD4B7OPsQd2SsZ63lp+WEc2lr2KkqxU
GnK8fzmnXJ+2HBZPOCJlQ9GyabeaQLpwcGJ4E6EOK8IWAbnc3CuF3LCxA7CYTbj+
Y7jfK/IRDzgE608T4wPwTf6LCtHBxC7eC05cM+R6Mj59Z8eizU4Tx2J+kLCo8RJ0
l0RJhh0hsyWp6yrJg73RDQuevjqVFoA6C81Yzd7mdezW9Ue6/DrJVaOe3Iebus2k
GyYYldCvShHasE41LJtD6aPssBoKTmdcTGB09o4ZhXIC7Yv38Z3xvviObrkZcbV6
Hae//oitmwKi4DAs8xwyjawG9slRAg3/xZQoQ/IQF4rMv9FdPqu/ZSD/Jvf2S++x
AuT6glLQdmaF13MTV46zowbRGbydZfo+IWOAvqOXOOS+CJ9wiSglkVa5u0AVly/0
yMHlm/NwDsqSUDuR5T840GhnOfHyKC9xvp7r01+5KkAeP+ggLttDGE1jvnXEUDUy
VCaRaSx/ty/A+MewKGsuMWiecU0WB9hkcGPcmlf9bNlko6hpXzBANaV29bZz8qeq
SCA2unipXE8PDe2L/nmIv2efttonVuVvjEHt0GAxH3z76bxoNO/AIAbJT8Wz/TJw
r3sjsdxD5J1C8MEZiGNrTefg5hfYwX3zyoVxEHnCXGSrWUIzAWp7lnqdj4Y/i522
sxKb6Qktcg7wYbtLxsfdQmS2wi/KEKAyFXZkY3b3N2ernwlLYn1WXUFAIgeLb8R7
1+06X8Q9PAcMn4u7wIBuaU4ZLzXkCE7vOCzoCyceiHLTMKgq7NCueXnqZrB3WT4V
y01aGYQNWbVauylvJi10LM2Yp9YKeKnD2wQ4BE6O99d4F7r1UhZSLi4akneOMENP
ejKFl9KNLtFO2z7i7nYDjW3o4eE5pkAfqPns8KseyZSeJMhY62nvsFQBMzAWQyOT
MWZI2J4+kmyaTUi5Gwh+reMUgPdCSqDglT8buDsq/OqsHSk4dmnJnAdFtJtDUW1t
GP5884bUke1+WHEkNNcjTGw3f5ypgb7BNU2byGkNufflHh2lDmRV/9E7uuO6DBKq
rlLavTt6b0TStuCUeXf6hqY9trAXQkhhKdBuofPqHCkk0bOxSaVdzfek6VJmMT5U
yOu7RHogopPrt/ygYjq9Pt6ECTyUzfkwDOaDdgttHjY0Z5Xy3QdO9Y+FPLl+4Rpb
jz695kZOoKoN3+Abi8L7bi7jK/uN73aMtvxHkdcx9Vj8x8c8eilaN2m3Fca+nhrF
lXlcw9h9gqH1Ce7prHe3rfoxJk2R5uo8imP2XIRB2vnvxSFdqw2p5/w1A3eZpqdn
U2n66ztg3wcR1Eu+HwCh5t32SN/Di+j7iOywHVQy2lj9r6eSbY6CFzKl/KyhqshW
dIsOZ9g4l2VuErRFYNyhoC9cHOw5GIMaX4oivXcjwV2wGA/3BtTZ2dYFpmQkMzu5
t5OPw09qR/Bo7jNu2HvsS6I/PHw4AR2GSe6fqefqZju996VHCBjqV8azJupd4nDF
PD52cNzs5oK+oyY33isPOYISGlJAzzIfBQqITGrPe4Nif1TqJldUAhT+5Wf4KO25
SzCh6cYY/sCNF9aa+7bqYxBBdGjfmJIawYr9icoQZ5O6w7e3jaw3QO26DOIBJKlZ
pLYr06buwaniAFt/ST7QewxKa8mzdMjXl8GfgtsgOSwJHaPNox+pl8J/aK/T+lK/
YV8Bbcu807aW/yrDP7mhrmnSAiB4lySe4TvgOflHYEhrOfUnhw1G1hXTk2+1phe0
5USjeecMx1I/7iwzs40y+0zgZXP3QuzhBkx8Qf1JN2TmVb4vmv1qLjOdK0hHJTZ8
LrH/YHhp4iaBxwC0dcKwBg88aVMUlJNELWEYIvXK0hc4BjiYVZB+AfYi8hIHBA9U
NwAfThMJ+KV3xx8pVUTkP9gF2LEKa24aqQKy4XtCGOX3Vr+JVRhaK3lEqXD0t5+8
wuSYIrNe9qavyXLSILFjDFlqK0g6VRv4hHzReU+xhfd+A1aMB/oGuUQGlaqNwlVK
pgEI38Rq4fXyssaoHv0vHooAaIC6NTKblHGHRWQWFSTqHf3rpRujzXTJmA8/ZoZO
nrQJzCCGHyp2zN/H1cBU4NIdjR6K4rRAHjIPZ03tErTiUC7tIx8nYwpPTF0ANODU
unGdRGUj5YwosxE0g/Wt9n4LBNK0g7mKg6NyGWh6fv35nfB3BeHFetZ+LAqGhmfv
HkNuBeq4VjHP89kb9IGbeoqKMP0wMk6RgOlBh+xl6/PkGaATEBKZNu2lEkDE3QGI
ud5eksb3H2hXrl60aNgyCZDo45cxwhHqEsjbLOIYmNGCL2yktXflLbX3DkvoJWFw
PC0NcuA2c+5LB4MUk3ShvkWgmxvi6uGbATIK8dgN67Q7iiBi9t00CrLzJvHv16Ek
aiMNm75XrPFlW6FEVCvQqf425A8T3gznAdTj8sBjRxrWks7zw/zmxqvEVYrGpLHf
JEGHSpXCTfOS9WMmIXL636Fg5/PxzV78QGAwHe7ZtublO9Bun5bGIzGMSWwacO6o
muWnz+Ny3edTzg5f7ylRfxo4M8bw5RA3yC9h1GQW56h4tO7IUmIIyNnA6RtQcvDZ
n1ulz6kUMyGbV67mreZuMaUobtITTZnhcZVflAGf06CfLmmywxDWbQSlOWk61Vp1
ilG48RDRb96RxKexexi+Q1u63OPNnOXsULIXVqynUhfxKdgMIOZUrYg+TbC+Iwnz
fPjtlfHN/m4cw0c0bbRJfU+YZD1qxaJ9uqAm4iGOcsi0Yh0gCafSPhCyPCf9ECw0
mFiU9BcTnSl3mIUvwegqCeCuF1XWiUzheOY/x1NB2cqGvGkS+2V6fGUgFDvAcv5K
l8NEhUnNIY2IhIWU0EOysiPfdTHh5P9SA1r2JFN9xPHFgSeIKba3h7bXgdth00ux
2V+TL5BAldEg2AtacBS1mV/uqLEvRDfiyJslJ4U5s9CZB4opvWdawDrABTh3pptf
BuaaVUbDXXMepU9n7KshWUG9IRdaKY24OMU1k91Xo0QcrfQ3533ixmmEuDQtvBJJ
djhM8ga7FqikuuG5M8Jq8NxFd77Cpts/dEgDMlIpFwF8x5LEtbUQHsvWModnVzBC
fh6oo1n1ztW/boceg9MEM5OKPuswEKtD28yrDH0Hf9BNrd739RZVQzB2lmT6H+J4
q5bkVe21oKNBT9MHsae4TGc7pKIpqgNiql5lon8ZDJId//Qsxpc6uSK3/SMLLXKC
V7OshgzY/jyiSpKYDDABn4gqWe9USimV6/zbYBZbRGbu/4erYZO4t3p/TKIcC4Qp
7Tos1qK6iWqTYXc3ip/jNugVB2MyM3j2pYwA4DoK6/IKKMF6QWJdSKoNedch3FJh
BZNUcYmkGj8/R6Nt/Dfy+Cf3QSXtpX/eAK8x/hTTUFv/8PXvthcoGZnqfIEYySso
xAaYEvILX0TbM9iJCnGjQVcGKUgI2zyCFtAOc/KR2Z37g1yxCkAW9wItMjI0P6yv
fkmx+VS67UtmuP53bznqzXIadDoX2wDyi778MO1iz9+ig5+SfBAm7ux2s2lB1Sm4
1e3iw6wrs+BWHNsjCUyOr+DE0nfoJBrrLhTKYeYRuQaSGeEbjIeYfNkbT+qKmUCf
e1THaQeGnRih1KKZD0RFyqun/LndiG2556A+4PbWmV4cMzc1zcRgrBkBC7wPW9Vj
qB28bC6zQJCmfFjgeOQuDb9otvKf5qkcXxonelf32T2/nNBKPHja3rlnUU/eIUZ9
/bsRYKF5sOwA7ljwV/VnVDGJtTrZjieUglq72o80lfdxWC5lDlttF4/zbiOcbDZ4
Eryn/bBKvXtQFr5vBPPLar6hkL/Tw9r5VFgma5KLdBrPxgtDexYTOQPgqqQ8RjMY
cwdtiRhErxfScx2hAmAV6nWXow8UsX3eJK144tb8ZxwjoJ3alLxgh1rUHkQtcoeq
Ogsok4WBLTl0wGdxQawRXc4tjmRs9/vFz6dBJpBFoLDiVgLCB/r2gr7CW/nB3144
eWF4v+dSqEkGca+aNPMXb56a3ZLH6EwJZv8rC9b38tsfFV1PShxKHvVwDxK2HVlJ
lvFZx4xvTNfpqq2QVVJCF754IbovkcUOTRESR3jntYvG3JTIDZY9HUAACWZRUgZi
FYsgAMLWEFt5+kt/kyw45hWA/eYLNKaEdu7ACAG3VMTZ020FJbDkGBLn/WQ4zHZ9
yfN/L2msxdTZcUqtSbXx/Y19JFLG64bWaGQYD9TU1aR++/iUVl6NYnXFk0wt+Hr5
JW6I4XNkYRks4i5/EbcS4TfEKrDn+8QXAyyFU2TzlO+CyXyreWp+biXDssJGwHP6
WyXAJT+L91ZCFshV+iqcqtINqH98DcPOU+qN2AF9WVT+ug7wPqP7v+FZR83KK0xV
Yru3QsdAmm0WnUuxHkRz3R4Fopiyae8KTUiMaU/0A1LOPutMjIK+zwvO40hdhdvC
SaMxDjRmSuwM9TsxIsyls3Bqy1S7P5SDRLnU6d86faRQwGBt5hwXZDyfXVrK3QyM
xxF/yJBDozv5Jzq3QaMT6VjYFoRWjyWs+T6zgsXeXYyJv3YUmu87nOBWmHTw+YQZ
q/LnLvOVS5Xwj7fIQg53jmVFLK4AwTSrQh6L3UfIA0At8q5pe7HkWKEstSLFfUZT
gIVxjvu16xz3fHi2m+EBJ/69NHDS4ZfDCqVfzNbHFxFdnJ0WMUA/KEh9O1K84qRN
kSB9pMzPF0+vT0lNDI8WREdFf3utd6sf6rfSiNF5inbsDcsYqNL0iJQbIbalHlT2
xe9vQ8Cna1jlQ5bWXRTdsVP8mZ+yZ72FJl+95vqKR3q8TIrNLDWPVGjAo7asRJGw
gAsyANJK7+uItMcmu2BnKB+5dMKAgUM54FQGM8wsSIrPKzcM8ySzR1/0LPA/dlC/
Dzlefx+y6Z3SQQb628A6sih0iMrCC5jhqy+B8BlEts+G5xC5t3toNsJQ+XimraBL
kCviXKnGGoLLzx3joqitRj5/jLGW/5FsW7GgR09ryQ9q5RQm3OfP29ScNoOA5jYu
sfz3L9DZ8zg7UmUoSQgULAmP+Sy+nYpjPNC8pSg1E6ZfIlKolJS76wGCAYm1pcMH
ibkZ6HEPpJuYL3j8MEw4plDxRiwU8IYcszIVyLIME1WblHQPUDNTfTJRrStJHF+G
eo5bD07KivGrR7EX/r4q/cl5FSxgMzgFah287skgQS7VabwcuOfKT0DiE2LDnAnR
wHWgizK0Pe01k1zsEFtQ8aLRFrmx7Bt7mHBLJDsyV52yk+FYj5ZOkeOIFcN0MrgJ
Ve+uuvpWWuHrIjjVKnzVVfq9odkdoCFQ5b+XsEucnhWIR9aRGnnfPgMZ83OsQ5b/
U3UACABbXUWpBYpW9pRNaBXM4AvVkbnRTPIjTc0i9avReVOJ48dlptLMb3M9ll3N
lm3n4pZ9Ilsj/8lJw4+6gSrMvW3i/FN/IvFRQCaZMF7GKJ3G8qPD4QRh1Rfc00SF
Hv8ieygrIO5qYcK8esMC70DmyJD9YHdCB9E5kZEdSmJmlACymdq1QKmaWXZmiBqy
W5az4D8cR9v94efwkwg/Z56EYEYfWrcz0AT4zIALkGUuqKEfgoXGqamRy+DXW1BF
Z7GSMOlDS7Lke2qzYGH5oE95oSzf9xcM6qfzsGhlZaMwXZA0+dEdLr5apE4+ZbUK
fihx4W5pBhnjOADR9LdJRDjCnv4RBeU5O+uPGLkakumyjx2fYg4XmM+nkxoTQ7wQ
StFYetyosoWRBnF4TL7Eh21lsqQpfisc9cUveUzj0wK2isAzyr3tw40r5z9HwMH7
zJPqTyNVNci050P+kypGNPD6GMlCc0ktFPzxMbCsBuMYvb4Tv7XAI96Bu5N6THzM
iMoXukrQE9Zr9B9nzN7dmo08U3kLfL999xETqV/sI21+4rlT0tpH6Chvz0TJ03eU
h4u7myonikdDXjLeSWOmu0Z5COOH4Zsc5xtdfPYVPxg5hFh1xA3nfak3CVHK87Zb
64Xt9ciMS08ePoyU6BL6ISdwS2DuVTYIbwvAR4dHrpPRKig0CdbLInd+ashVCGwI
wQHNiZu2gq+f9lq+bwusoT9/cOSYrXxpFBB0U77pSnZQ14qrqYR012DOmUl6iP+/
ZXKhRuqEZeWW+NrgakQYIunCLgIxd8f7Qd6dSCW/CojNky4HSM4C1bWY57xuP0ET
UMTQ/A09CsLXE4XlKpxaUhGkWrpWcmQb8lxgDdOrsCLsm24uXr/QACdmErPrz1nK
q/w4ul3IS1BLx4mcJf10wZPVSY7huWiaEzsdPuAtyPaxCiIqHw4fV5SejvQaaPgz
Vh+1lge2eIBf8HM42GvgqcwCR6cZfQ+xWt77lIvYQUHPFZ97cZbdnnn2eHIIBcko
NKQbVnrtRhTqSRK+y3L54JAx73dog1hdLlH+pzYQi1KD6i517OL2l0TFTsXjrjQp
3B7jH8KKm7W+VNSlexN/BiJDTreoMLtjh+h81i8wPcVl9GKm2/m2gHMNf4Bieq2U
kfTzwqsin+jqMi15x9KT0fhHRjOOWP6yvt603M3psu9HZdq0WGGz9LtCGMDxbEYW
zaNquwdO++2pFWCRvcuVXzB+7/mzKZwxmuh1F5lFuuaN4pYg+9JDcfphIhX2c5MI
sqEG1TNIY9dJUmm0YO+Kkpog5BpSFck7cufIWmOg50Bnr7QRKi7FpAnWiPdOe0d+
SPVBg3zy0rGlBHZ6N8rt9683QhM0OMOwDzYXwGTS4ftPqbSjYZDBu+9ss5pUOODR
g3r/bkFdZTDB3lIybRgDoE+qVROjKRT+zM04RJfaXrPFQ+vTwsny5KB1W4UBgW8M
CfV4J/++QhXuS3TkwfvQSEA1k49M44H4n5srFruUqa/OBQMjti4h0+d0vyVjBhm0
SO1BNdKdA5p1FsYDXjPJK69XGh60iEsc70qs9J+CSMMl71JNspIR6TPfK28AGpPo
aV2uSbAUYWYGFQcXGbFYHJfoO/3qIpVOguXrq1BN+Z6DZ8QJRW5anJ4osCKXfSza
PdWVa6XRmvXJlHUycWil03JuEO2DOp+zqZGpzbZz3LQPU6ZlzulknOH0sSJPSIEZ
h+lgrGz6XgJNFp4y8BUoFFUL8sF+F8ZNiAs4Stg+TFymKxEBpfs7CSx0lXY4hsFJ
okcGKrccG9JqL8L6NprQ71pEb0Qltg7vZF9z8U6LnyGGPVo12VlMEreEf4iSHfev
KRrx58EM9tAGwQBUbBHoqV14uC7OF5AIN0bUDx53L9i/6S5ndvmLeXlhEDGA1mYN
/eVpZvD1sG087Io6yFzfulNzkpg7JUKEfn1u52g2IYGWEmN16PpE02uDTOxGMIY/
KFB1jb5zwQXBDQBjmAeyLrgAJh7U5wF+LSIhydFrS8FbbrfeMJyhN36reUuvKvZG
prrEm82x6SIAPWkUf+fZTmIMvHXt8hs0JJ4EI5Ad9qE9DR5LXHIK4GYBQh/3kDud
omO4fEW2/bdr0aPttRbfU7hdZ/xhJzCXjSU81SGrBiDFgyRM+gdjx3rUaYPlKbYz
YBT6podlt2b0/2/5dM0RzmWtNGvC4/pPRMiEduePw7ivhAiKZw2d35oraWtIzNxw
7Vl0g2pF5CCwIcf4XFl7fCANGtEt3gSJ2U6v4OG7oaj7AW+S61a7aFIz3fTvJ5Ho
TQfE7MgE/UdyxdmLxLTc+mo545Bds4MSb32b19kMitjq71mzbiD2r2/gO68Awk2V
VkNJ0WagdR0qXO4oNQTJeUD/zBVBODl6s8/9SY3RL6T6vmGcB0yFto2rFYAYIcl+
FwgVK12/deBzH63yAcJP7rNhTFxI/vhUAQZDh/99AKTV6uVpU1VWy/ZTjUcsD+Ek
ZYTgFQdmOW5IyC0YW1g/33RpfTnzlpqwU2P6Tk25mATzdql+5i/QVWxtYc3uxzd1
ITO15BpGOB/HvZAA8FpxmGd/Tjk/Zo6JMcfVESQZ9tNhZCbQaprM6jgBr98NBNgm
FV/PhBQbmtaTUrVjBNSuXyRsavHth9uPXso4LHcNMKf9JUA5Sxnn8+bxO1Oz2YjB
i/1QW5xya/ONLmWWHxdT9mnZVloTuMzwdBY2ZzBGivgvD805guqw5XDyBUa/unqz
nT2G9IbcZktHrfkbY+VDbZkUmFEe+cvlsXPhrk5cgBi9P7cs9RV7SaWXoJe0rgRT
sLUlkp38DOotomD11FZd/mdgM7DusH/68iQexKqlQ0jHKP7x51kJzLUXMTgUyw0s
RDMQkruxXfVbL47TK1tr5xdR5RoFAdMOljAliiCR6JZ5e5rGjcXDjOpnCPFS0+mN
zewZF/uwwVKrzySDfyGCgdFPYEcKm9Fc4cRJs/NuKQPLrXsOPmSWajKNOSL7bCFf
gRVqmOzfxAl+/ormyC4iYi8BdaHCnyI8OOAm5aASnPIKgQyVFhn70+inXAYcTyrn
sJCHUeiNawzrf8Drj4IzvgHEanlHE2HSm66fbrRnKFoXHDl/RfzxdOdVi8Dskma4
stM55tb2rxbvXrN8tewkwYKNHGi7nVh6NGfRfHHJ7XBfLC+GcizUs4Q3npQ09sa0
+nT88OcFehpNqQZjNAfmqIGOgO5LR1j+ebaW/FnFfe9TO7Ujf4b2EVerg2HMFyC1
nQYWYwBOCE7F2eRmxLxe1h7DH07iM04pPWfWZFUKnLh4JicLoOGR3rs/QnjT2EJv
DJ09xrwxpYjv1lLnlsX1/EU2pLYIFDo4WE/oKDZUaQ+usRrGWVOquwpcwroJkD+Z
a+Z/gIzFpJJ95dua3CupqWCKMIoPLL6YYEIobYoGICOA50zuO7dF07piF7+tukRr
3VaoVsMm4C1RXPHhGCkYBYyn4UNGK6DxnyuYsxc/TJ1m3h21eWNdhugkazaqD/T3
pXhTtfiJ2+gU++eeQyTrujh0ekkt6B3v2JiEJCLpUHZSrutMtm3tEhjdQ0OmSQeb
PiCaiQApyHkoBBWeiTfqhyhcxmrcDU6yGcONZGQAei4pS5B1f0ptz/Jb0bdzZZQm
sD825aSQnmQ2EtTj9dW01lGsOllXhCf9DXMZHUbKzbyENg6KXuYVppsp8dg8EbyX
OrB9OXiokTe5F71bS/mDuEkCwFevWhO438ZK50fSaPIOpmwTq5WevT32xe9lqc3c
AbllM5xXsvwGR4WBHZfEacTS621roGy4MvlT/7QklcNB5yyJSlMfasCkMfcJr7Ub
pbq8PSQjyzePQGICJIwn05xKq3LFsNgnpAS4OZGEXL5dKj+HtFApEIEGWAqPIcvg
jza6yy+hBQ6AdoNG1Ogkw9k0dW1uSHZSGJdW0RAN5wwvlTr/2waZlAj2HAvQveKf
uzLnJqlkESomxQz0UFp+cl2dgaZfG0GMgGhvDj2b4hPIDm8giuHKvUWQfSRQ7peV
bMarP/Ikj1VthDgNOkXIlhjrTrlLVJx+2lcf1F1MZEX/5fKxeoSRA670iJtKd/iw
DDYX3OfVzyY+4/+5US/cj8RWkDDcfxa/HrqsjeX3LlhR5aCDG9n3aYDwR/HU8mtU
WhwbeJj+wX6qenv44IGb6O5219OZqUHuiPMQ9aXm/cbzIdd2Snzea3zuEk8G/7KB
oEVrWbG3jyxMhpxUvuk1P6xECoYwuX3+Wu/eGJLXxyHUjxqCHC7rhh+ACfcUmidM
kPww9+KKL5Ua6bVr87pE6YNTbY3YCtxlTcTCrI+6qw5zV0WTvsQPRiZyMeHA6W1q
XzmuZiYtk/suEOB0ZnQPeoGCHGVUUmN2A50ujcKvJ007G7hc8eA9xwGKiu+IzjuT
EQbZxnY0ulTm1qB18nCaMKeetpFJLVcqA1pAC093RUBab1dhAu6e4Rztt71//m3g
4VOXiAGH3fqCMhQ7Et/KUnXx7MJkC2xoN69SVfSF7uw1oIOLdqruC81UJaKnx++M
izsLWU53ILIfPY79LSy4ufr8EirxfOH/iTfsvrSVmWX8eXbVf0S+NrT6yiA7NHj9
jNj1eCS+efCbwQDB4Sk5RcgFY0zMkQjsyYJrdVpCt59Xz7OCn7xT2u2rpG8ZxGUv
VlrSiB92mYr+D6AQzU//3rqTTSD6a0ACJZAxc+nsLfUqw63la3/re0w4KvJs8kZg
qcCR3o2OvzFf3Qi4crBf/3qdAeV1RcsKkASLtZ9qjXYs7XVTr39ewW/ebcK0yy1l
Rf49tvahXhq2iCgGk6v5v1vedSN8kgRU8UOwcVc1L9CvKg5c4Y/b58hl6X93/JKE
Q4Mo/hYRfB5ljprj1sWoQTMaNjriniaszajddi4NETlPdFe16Qj1ju0frZm06+l3
sA6uFsnJ+e80LLW1M+qCt3DI4DgiYjPjgtbVpeR3EoAK4uiVzrEXJDlhLTkSGV5M
G/MwLJzLZ9h6cQMrIpe/qVuIY0C26WfAzZH9lmEyelsD308BM4E7pakoMPdSkF+W
CCuMLQTdqLT58kPilzjbtoxtvAUUH2OcmnuYhNURh375iZDbVMXDbVOJmMneIyZf
CwoTFC+8F2MuglaRha/twG7X5PUxtVLHV33CYhVsIP8e8JzOHlHIwxo4UQXbfnAT
pEyAQJmvYE52D6S7x+v07+XGTjrbY6IeAqefXt5FknJFREjYniskNkF5qeboDSOZ
jCE6Q/rVQPjzi+LjKQUDHpWZ+pqUTZeG/+MAYdTV56QgYAJvEU+3yjEARia65ESZ
gY9rq/no5yUubTPhFc4f/CW9x/y8CPs5e3SAj9EEyNDMcz7MGftpmRlzHVSk4D3v
iDW2Tnhl5ADt/x0DUBB54WicEkT1BeHIRyI6golyI3dTqBF+ujekagYPrB9RrwzY
+R9/ss0Fs8ItG+APPW1JLJis9Q82fuFFB6JqZZG/1iiWBgb5Ss7c/Vcddbfaadp1
t8YpdfBPqly9blQc1Qolcn6BxQElG/HZQbqHxlx4O6d8JABszbgz7q77GSbsMKGU
TGDM1PTjQ5aaR4Osi5rGOHITxi9T+aXe736DauI8e4v3paCZ0SPgnFn4NQt4sWog
XCqfNMXvzTFAcso1BpkdxqeUjQIem/FSZeIiFMEGP4AlRMi3crJaIMJXoN4ugjEc
wODtssZP4qKtfPept9E1XC3tz+nt8Bxk75KtYmS5ZQCP0yusNwN6DWuvfAoLnqgZ
Ia7fPOLB7aCfx04WaPE/948yT5QNY1PYpxCJ0yrA8TWfys9JaOBImsxqCqytz6iY
L6c8GY2JlT+geFBOUdwABTfok0Pt+Rl2RqUj3FkuH8wgyibNkb7G1A6m+nmITUU+
KPJDOEQeUKSKR0Onz0o0XMwMWLJcHpSG3m6fF73K26okRFSgWWfXXlh3BzLQZmps
5jTYfyNWJ5QpyHqfhTe9LVNg3W80swzuXYGmBvN7T8wLu0dXmBRI/joTk5xshu8/
BqLgC9hA73zHZ8dRRpHhvPI/xiAVQTlKyNmQHJCLKOHvDLmVdFGcHHIlw0lYfTgj
2+aCd4IFmmlkTvKVAa7f2MCqUfXtK6mznMKqdqATMG+mgZc2RsiZAQHG64gz5urD
urG5hETwFi/kQyLrG9O80zBbeDbfp7QhB/s+mKIpwnWkaMsjAfoJZgTTVG0sBtBB
4sE/sIhOuVBp0i8W33xuIrYfOa18teEMsDrhBvZHO6139OYz7y/xi0i5waOFxj1G
GNUqqgzm4uvRqQTRHRWb++cfGlSWciCys2JVlrSg1JXmDkFOCDc8ftMI9yyv9jys
DJhlM5kZiebpLI5vwuJubOfU3VjTge67cB1taWDYJGlbMyV+PIZTuMsEe0+v5Ht+
DDdfueMX7VbYikeeuik8GaNBGuGe1Swlxp7ADAzikVN7aIlV27IVHlqqwZ+bXXmA
hxNF8qR0zeI3ddz9dm1eeOgCOWcY/uKh4E5rCG27K07ot0VrClT0ud44O+E36HrE
BkOZVTL1SscjtQGp9xo0Aqua2Al8SEpF2EyvxQ0uxNXoz7ywyN4v5cDYqzTa6P+7
J/xWFxwFUBBYt4k25MHoJ+p8lDD63+6ohPUu3LeIKjUFaBw86fd1tyYL/Osdxvn0
54Mb+8lMjgRuNtgdvzezALSNrhHuhmpuP/hSfiTvJav6KLIURHWJ+IK5pivcYkYK
/aRw0kmIdz1t8EuQoDCQPVn12Ryn+8vgpnX84m1ME1KtRUPs1Nm44TbGEoGpO7b4
f9FM2JmDQZaHRXUPOuRpcHjulwwEqsi3IM/p9EQnkQWzCsqiThkEOOI/Ae++Npvx
CEjvA7ufpQuKIn3+zjXnmTE+FMpnEib+GxQI4KynXobEf9tE6DhGzRBVTKxENqat
GwJuzilyKjzd3GsQ3gVFvhm95OrdjYCrLqB6CEvvvIxDLN48tM6H1i0+Of+GFHfH
jogPOvPJ2TvCpnObePYwik9eHNGwpbGvZBK8nlxRYsgys7Pt2k9kZx2wdoD3R9gx
NuAnucN3ahhnpm8NjsSjiGRUPKUIoUGa4aqsofxew3UkMLSCeaBBnOkqSSbOkeCd
HhexaFbX+3bXTIjvUKQnDMrCA18yhDOUx/KY3kHTV2lPfOxM0X/5WHdUHXhXs1Uj
x+DhyDq4Y85CR92zTVMa5EEevDB56bHm392Ij9w9cH+btsouYEIeAfMYT4AHYip/
1FV7RLP8/vtCBrPOvuwACgzg839cA39sgcZL3BEiux84Awca/wSalVP/EcQcRyk/
rd8gmHumQ30Dt+vqu8BWIEvrthBIRPPzx8y4/+eog+AmzY4d+xygDWMPb8HZdw0N
h+82cKpli24MKt/xEj7A6u8U7HeBbVPYWJlSh+U6OCuaLZgNXF9t/AG6JzkDli6T
NQymrzyUcKIYZBsuJLE1FR+qUWS8G/dIpi7YrKSvBfGOOghW7BRelKHLlcTCTHaf
XjueeU/DiHl3JlZBoDjPJhZlXf6jR27+qjqVu4rSBYP+tdDcbV6crboNL4XJlS4q
qTJ+S/9CJQYSv8hWckF8ETpR9whGYxvnaV/jcDHZHFkkCrTB1U+Sd3C4+SUXFQ9a
lW4ijedi2zdcEtiv3Ti/jAtxKtPDzn8rCmDvUYJBDX2nk7l2fban6Z4CZHf6RnC+
fhFATWfWjrXM0Iv6v4xIxhN+1MMdcrOB3YeiKGMseYqBmRp4Zv5hbbgM65fHBE3b
wQxiJS3llU6RWvh6GIfK/CrBSlEpkBJ1zpJApPyFKeHAVDdj2UCRG7bklhyBPgeF
Rm7kVtJyTzDW2cSU/LiY437D3m8XbfOkyrGQ2hJBh1OOjbFqs/bGHGAztqAVh6tY
TcsJRmo6XGdSP6OKYcdTBkVdp7Tqul0pU7wdcITfGGyukp+YOmH123eMFZBnXXtX
UMIvnzhw5jLUcN96Y6two/SQss0QoPOv6IN9mPLWMtYsLV+WEaHIgmYU1nLPMAkE
OXnR1TEDb96y123BY2hGDGbzGAR5dc8rZnLHUyyxZKoy31zMOlKRZpobjhPJIXMF
AQ2JekLqPRFQFwP6RCmSUxcm5nLjiNDZdbZCcCgrBjcHbC+K55YLxD/EsTQjEdRW
KigQwpcGhgLPY2fH9lJmPnYayQBbdoqMuWRQe6MzFoZYokIAlneOxuGU7E39TpKj
o6q//6kzijND06OD6g6ZIzOtVQWrj1mhXCX05pZFcX2rm3XZLd//BOmmDSn4syea
yaHY2QOKyhG+YbNZdUrqJexT5WH9wHvVQVIM8PNb3srgk84vqkiuO6WBLuXUtKnS
Vpl/dlrx2YeX3ddboGUqydiyrkyhlmgxf3qO7vIHxgTA5ilmmDfzAS6d8jrzecr6
iUpI0RkjuyIyxBx04kAo/HP4ehPB7RZDsua4dAeVGhoshmtQ8B+W9RHIU3pxueKw
J7LnmwHH2gEKlzCW9OyLbXJcez3hxLoKAFvcS7iUq9iwIrMkCHNnE/kHjUyB0qdR
MBs2l3wOg+K/xUWmkUclmQ6HFY+9ZMClILIjVaCiXYxSukUNNiOmlK/K2aPnM+hu
Wm6Z9vcdsWpFp09JHXa4gBTQLduFytY+Fezh/tmfGRVsaYxwZgSoJS4+y8BNb2Yt
CRPszG5TWItiWIgnS9Ior9isIXzqkVP09YiTIyj1sIYkSR1UtcrbTeZ9OnHotu+A
tpez5iUAVAJDLX90zi+/cICYJnqtWI8eIUUpZlFH9xpzf4a7X//k+tp1SQDoXVLU
Xc1ddM80ZYDYID5moMNnqCM9tx+xoQXdp+1ahDQ7NsUxn7UNQpnEQOzo6hU/oRD/
84IftSRc6dlnhv9jwbQc4xgvL1RPAr/3wGJyJ4APvnhbMCHpIQwZz428hGCjFruR
sFvRnefZjXwIrfI0umwZ4oLlj0OEnlSP4qFlYB7wcoqc6w84FHly1Yc10mFuZqi+
oYgN4qx39klnZArzADYXctQe9GBrX46zcxz1v16w/U7nGHMBg1ucCT893lBcG/S9
fweFldLtQH1v2Kd6X4iaHyRg66MCgp3A2Wb9aspSQv/3GzY1Kuun0d5rFHeJdoCr
IGdaRwX23wmOj5A/9DI0b1FjiUOyyXpr9GxoDmDhsbk8J/U+3gEbfen7jq5nBBjt
CzK2nwzwnBKQEg2eqXlJ1ucVlNLpiPvF2yKuslenEJybkxoqL+ZrSiIN4STLt5qF
kxO62K9KkBvI+ZzwH2jlrnFcdYOh8iaRVzDQSAdSissL9CJz6KKGecVZfYvo9qN3
fjgeyjqtGUv/qiZPsNCVtep7k+89/7YVN5RuzubVY96OXnbDGWvP4WXQUpTtRXDZ
6qWECDAeMvIyPre/4Q8EZYQV2IrxFT0fwSOIc62YFpqpaP0IdPBX68X+kFNuLBfA
1c3EuNllJvh4UUaQ3IVy9B/pNJuWl747D+XZd0gD5Srexpmo2OrzYfYmc1H1P1s3
NZh0ceL9Peo1OyNhfsjQ/0/VMCepKghLbDuvxIkuI0fpl6GssvX3HCXbu93zFkef
pHvfCpS36UaWP3dPjNVVaOwi/uIalasWJOut0Eunyme4ZGzp4ywIYEGvmMI4nEIJ
z45t1m+PWotX0KqIaMYrHvVmII0wOarC+u+eHKhJW3tzUVad2c63HaOJ8fnXGCiz
JENUsK3KuzvinH4Hq+h0CBlsqyvQUhHLc51q6qzDAWZ1OipotLY/wQuIuTWhMfTq
K/lVzgW2IuLpQQ56Hes35n2R/z+vQ18fCgEVanTrktty8X1T10ENii53syFkb01H
LsYA0l1TxccpISseMsxYJY25KYuE9nZoWFE5pu3aPH0LJVrNAzsYxcOnv97cgt06
/D3xt4t/ZZ9+ywu9CiKFO7p621MTrLWE/PgAGSMIJ+x0cDwwZhYjC/R0R9oJp5Vc
/fQbdv14AtRJ9j6E1kNqKLzINpZa5/SuzYB9kWErFJC7O3rOYZI9k4/SIjYPBrHg
gM5xhCDDIuwc6MkbsC/BpQCWLt2xz+8OuFrQrt1HcU7j734m0Nn1mCrESRrI1/Uv
1LDKL03N23uPyBFUFtEbHodeXTi6b7BWQA+e3NDkCxbkRVQJTH2zrMKV70zA9EKU
ju1oMtwdHy24PARWGip04WIbwEQi/I4URDP2QmT9yhBJFCynvoIf5oqLSYIHqe02
pxNkIsmYgDDmK7CdUXVxE/1mc+h0lYP1FOn1fEHijZejvuDXsoz1GMS9cgnAxnpx
AeL3lbIIyqktvZ/yJdq3NJh8bMhnkibYUHRdfHT2lCuogf0q9f4b4aWouXARWw4u
7hD4TTgXwgb9OEPchmoytDPdbwSOzbEW9W9F8HRkpPs+7jIYuLeYpmViEAXe2Jdt
Uhiptkb4hAO3W61zHUOftF0uBNwVHbfzARhzdLQx+t9VeM7kN78MAZeBW+8wNUaS
ajMkIuZZaRdESysIDRJwi3oOaPn6h2DoAEzEfDzbZSGXwZdIfBFgI+giyQFgY1Rf
0rPv7+ppVll1J9CUf2mCLEEKaBJcig7MecYMIQKtGhCj0dRTjFYgRrieU9/6DwAS
HU1Q89KYo0qfT+8nXg3reN5yCjv1zmJghMtgBh13zzbndpXUbhSaJ0sl+tppWGjP
TFHuIfAFK/KkrM4d5GBsgp+L6yyU7v0HnHaUWyJjN1339Uo7rXM6MLrxE4H1Q30p
5e1f+bMBEsV/JzZQSZ0xT1c9tNyyj/81aiRLL7BncyjG6OXRKdop4LgOMvwSdNwZ
TfmJ3JQ3FT9vuwQGI7gwUD0dwb+5sfBZrv0WT5IPH4n1UUkVepfgzJLRQriO0d+9
2bsgb7crCTk2mOtBJTk+jGFVRhWmIFeQc5wzhYvMKetBOglqGH+rtcv6QujAP/ys
2m27q1CfAEwOCm4Mol+AHNhtZnOmImMk000X00zNojf0TndVZG4ogdHhXCP7k/HV
MlABfXEcbZYZCnNNFTMEYieWsu2Gu5GzOCKHxf2GjHMUnWdCgWrcifsbvSvcGl1L
mK7jsqcwd6n1v7/X6OEYJtBFT93tRiVtnDJ1c+SwXGnfeZGEyPoc7ITAT3NkAqWC
ZFZzqzovo41BIY1Tk9FezqBcHnxeamDFeP5SuwajR6ESylXGi1fOcMeRrA1BzAag
LCVLKZs7W8tbMPtTNPSL+CP6VE8njTMx4z7TPGAzXsG4Wi/JsuMaaUkWwhJNnjE2
m+TSCIBsgfjy3qytg8x/k3woGK9SZK4np+snAtYJCcy2d4uR6Hl1uFndWduzC5Jk
33V2svL06bj5mLwwTbFdlKRRZflD+9Bqq++oN3JhvaNzQ1HRqlZ8SI1BBH9aBEVc
g/8XWjVSDgQuPiq4Z/lyjjQSohdyJQPFdO/ZBF2iI2cd0Cr/TyCcl9MHs4wkEMb1
C+tovB8E7+23UNMMLkUh0EORuHsdfoQJK2baGjBxD8aE7Lls3weilSz1850SIjKo
mcgBS9YFMceHn78CR0khjQKrsk8QREuOlTcL4bz5vGLXDmIZV3VJplBRJ00kryPi
hY/M36Fth8C3ZKzpfBn0ZluZG51tpdsCnhZQ+x2DxHdVvsddJ0lKNzVoBgc7LuP3
utg08hQLMlwtkmZArxEHWWk3HEyr7/m2U+KVyoUOCxoNpyn6RbB+N/R2YibgNEhP
M4zqTOBBob/XlGSy4OUz+Y5ZmlRpmYLnR3oX6+4Gf0rMvneP9sI+R+TbIfKH+BsD
By9e5F6E80LrmQEN/0pVK27i8kN5wL+/y1Xkp3TwImbd3GRI9ZE0FxnGr8FPlr31
i89wkKjYxQY2tOkbE7FoDtv8YP1bP+AoZyP7av1B3XD2Q2xqtfvbi0U0dKUy3ye/
3Y999rGo7o8qijiJMNjMHMGaaoT0YN+GxFvlvuZii5dmwQ3nn3YLSZXVsqpeoX9n
aFg2QDrVUJlDIvdvbNY+6LXIEzTVBtQjWW72dmj7RVIvUnv4qL+A/+YYJtP1R/Dt
tQWqZFgwP9AiXjq73T9n7F+eU15PCzhPARWqd4Reg3+DDmyrWNBboT/qpZvuS+u7
4Ocvr27yUEwp8XFlEqJnjJAx0d/Ipkn55dg+oV7FIsXslmoGvMTB034UpG1N56Jm
PyffcYUeUrxV3Z65ZwUh3j0k6C0QozBZHmis2hVvUbCf1SxIYoIZ+MLHCoRolc+s
Kowkz4+dzwkCAGDVid+uOV2IuO699+IyA0aqE7xIAuoAFXrRO7et44ANsavxDm/u
UOVhT18375lDd6RE7bPDp0zOqgDkK5+u2TRBsFdX0cfwH2XHA2zbIJalZu613x0k
73ezwyaw9m/D12O2n4vHR2OyxXp7VQELCkU71i6RFGimaHua7vhqpN441ECgbmJz
PWtDhNJVp0B64x42b5RA3vg9jtJUROZq0JnrdJZF4zNi4CzpjNEInGqTmZpBjbTD
6OCPNK2u4rzuNmKkofHZmaHIDBrVZmdoLgrOanoaV+TuZ2lYgrP/xzdOFDkE5OT7
G1DkBoI51ZE47qqupH2pYFQ1dhfzV3q4b8+X542NzyPeKrnpJQ9YiEKvXjt7kA8v
cEIzKldHO/yoDrfwak9A2JrWVLMER151/8e0+HKYzjg2EYmUk9BHv0/rIFniuwVD
QpTVq+Q73hhLYS69UN+dQV7w7faZWk/8ydq2mQ2/JZ1Bhnicv07FG5ijXaRK2qOe
dtyD0lx/1jmcUEBTYRGOPq5VV9DCS0Aco7yO3RuFgK1cl1uF0eKf4N9bLuPXom8W
uuPL54TvhOTYLHpV3LbDgtOHEt4Aq785TJumzsVMm6wS1KqayCTaJgB5mnTFAqTj
m5RcgVxgaF7b+UYfTWgi33hGZ5387cRWN/V85hCZB9nDKXHMFyGijX728S57cADw
cTWCdw0ZyubsUROxVYHI0mMatTI1A8+pvWriaLM1d9sUcs/ylp5sTPHosOZknbPT
x7skTF+CnUqJnEhLbYI3Bxy0WfeSRHEBWwtyxTCtNUsPSKq08H1z+7sWneX4iU/J
GFPEVPF+qaMwEAorvZzNW7pZ285XQK3tjKFN8H9zicqmSwYMoQ/AHcBje3Brs8qu
Zd3tdSYS9wYdUUAR/FQaq5/ORZJ/+eDSLcGTsgIijvzPpH4nOGIXNNE4ErxfmzBN
zNZQfzY5pu51N8oeXINNQ47WP4aPDdrms5RglubeFA7z9g1l9Ab3ytz4aBjhnXDk
MQBPpMUhrsyK4IFPyU7ZdF6hBi0/6XeZwbs5daq/lCZPLdwL7V+jjw/uF1AwM2Eh
+Dw7JnzjHK2NaTeoid+mzR+4H+Uo/eJvR9K1iO+Dnr4JRldv3BDmADHkrUJHXDMq
HX/aLakrNHSsJpdZ9vKPVGfWFoMZRD/l4PVG+sr5KfdvxM0iavLXFiSw+2ID3PTL
iUM0uqfFZgW7zScE147sEiuHjicVOPf5vakGBayepJZGy4yqMSn+DKyN9lXVyEWT
fzszsRnh+r+8z0I+OtcqorkfQsISFk0l22rxtTzsUh7uFp6t8OHwlPW1hpdeCUdk
F73TEOgcI/qsM+j6xTVW1ka0JR7/WfIqNx4hKPt4OWEIk8r3l5xgZsOwuRnR1Nw8
v/6nZN3fPhK2tBYh9GDDUU3RwvS5Nk3UhIChp2njLrO7ZHRd4gP8Qc71yKG5oysk
t69aS61tI/5jEFYAqUGu4L/MIHewGtrdCRqaSvR5pyj5XrXVXKrDItrA36LpCY60
emQ8TkF1ofKMrDVTOxl4c1MmwQTbxNFleSKSAVZyM1Kz04Nx/btZ59LZ+/y79GiH
M/gPeanmqHmFsRXQkZuUsh9RKJRneCWei7JdvGs3ZRgEpi9rXaHQsSw3oEqpz4PK
OVorGmpPA/ZcN+qfn3FKuDkJHVHEIgXTVWiH+5E3cNgO4tJ3kqDQjDEiHYuGv6p6
WIXz6X5xN76v5BtDLNC9IQFQCVBHVX0kOTdExwzJa/NIyAeTpQWpXRr+6GDA9qn9
i5YtWYEF6B/OsT1v6jEELxHbsWTtsPk1ZBcvKhxJKN6ZjPj3JJZ+qXC9rYZfJAly
iTGHrsUSDagAYYxto2p4kWXlIRbelAwwaF6mZ0lMq/R471w+EMSful2Iv7+pd21e
AzF9btjOrwoNCZkykfIcksAWtnczr0cSQG1aJmhmIhWsMSAKmAzrRooxpzaSbPrt
6zCXva0gZPbomadUJpGqlyFLQOKExUbAVAhjRisp3ZYxzfkTEGeZNXeTDpm1yAG3
ShyEygVq+oC0uZzr0XvCoZnpqnu0rhXot5G4Rm8lEkxSuPa5/G41hWbjtSnP1pB3
9a1NTFM5cvofIh0pr6KMAsn9s70/WU+J8I8gLS9S8UqQv4cXpbDn88Ebev2R6FpO
o9xRqMCUsNnUYBd8JLKC2WKZOE+7wZ/5ppmEfPR5BKfot0wDOF+j3aD7Vh3OnH/7
r1X7oSDeUbDNGJN9eEs9x9zzJXyH1w2o+HlYXx/E+PAQ5Lm5qIozpeLEcWYJHAAD
Lf+70JfUjgtm+lpQo4+z7cwSdFdefv1rSG1/Mv4MOlbfan/eXWJBj6jM4FoTVEsH
EgoN6WJ4RslqaD2fJ59+ikhNAhqgnZwkCeRXntSrlWIdFDiMHyI/e7SRy9V+U263
s/FBk2m2LP2NkTm5NzOA0i3hSnDHPthFt0d/1r6W0+LQ8laQD04E3amRgRvIkJ/e
WfCcps5zxOgCRUJ3poZAi7VL21b7NnhQaYXIr29+PK1cBOltohtd1lvSHW2hcSlX
q5h65vrq3CNtAlyAC5JJuLPbIoJZnXqSDwE+67xd5ZrzLBhOlfatW7F7JRGbETFt
HIEwiEzvtkc/BKfvYIj9wPITkfuz1HpC/nLuWbYkdmLSKgn1AhZi2vTInBj9sbbn
bLqroYL13QhYwBGLTYsY6s7UCHvduOlPyfBSC4FWbl9m2n7s2TzMsF6N23L6zuES
1lEOP+ZTXeGHyQhXd6T0rVtl5l8ubcYcklPey1qTIlMykzexMnwuEQn+Emeovc31
KAD5nWc0v/MyiMsni3vLMfgr9HUNLDH6Ymyk9V4tPZIlsB/IZg7lSGXVHvadAG+H
RjjzGHznOEfj/WUMO5m5MlgX32cTHs4AdCCQxFYl3F32jO8J4Mnwc3LRP2O2LgE0
k75tOAbXG9Lh2QKvCp5KLtnoCSi/ijePt6yA1pTERzxbyZZd0T61pk9qgNRtCK0s
I9RusOGmKvE+4Ko3jaAc/KWQ2ED/+njf6aILtsboLMWAJr1wEQ1kXQVnJIO7qJqh
g3mF6wsLZudUABavEfPrwcFcbBAicDEACS4bKSWzprC2WCQlNazytb2bWOfPsZFX
95BJWp029fW3dPFXTK3W45KrBCg/rx6Veer/qWhzXmUDGL9oZuMFqjenI3W7S5na
5DxZKM4EXnWl9OIJrGl4joIBWD2TfgOFNdYEb2k9jzyeoMJtN6WQNanVpw7L4M7L
9PmXZkDbnC7pza9dg2bm2r8sg3eixjghJ75kR81b2IPugHqgh0J/EPbhO78soyhp
eaIbapCYZPXVppAiRYeXQGlwqoruK/de1PcBr8ZW87X7aNMsgn+iiW3QKo+P6BZx
c7o7LPQX0XIpEi5vrUW5Jy4ZWazRB1Gfgp2wvdaylKagduitiUYXplIWVqYYCV4s
sn7PMdx8kriubE0zwD70BG/EkYZDW7wx6Enu6PsGuP9QZYiixZWQuhe5CoMSPzQy
/nt6iiWo5Fz/bdWn0pc3N9YcPbvL8rx6Huz+2q/AWmexHBvcmvrVdqSNB2BEb+rG
SEDbf3PH2IAYVZHFma/EO62mm2QNVySJzM+pwH5Sc2R8rOHBPeJoSJ+EeuppyVxu
nEpJldMENNTTjV7XC/LKGp0BQowTRgb29da4/nnLnsHfI85ij6eDAABWADzPKD3g
17+KoIYkwyuj3T2ELKrx8NaXtCuXFMPifFZ/byuNB9SLGio2WN4rtNsbr3JR8V+K
PyNM8Y1/L1MGM6HvQNrnqiezl7wUoj57bb+nIIwr/9QxMSBMKbA6H9MVeRwhKfZJ
OnqoFbqv+1+3zFk33ZGw6pLgyO2MPhg3V8Y/zC2FEZW4bxp43glNU2q7Z24Epir6
pciKboVmTGx05fAyR8C7E2XuNzNnZT99rzC4WHy+eHBJf4yOpQ4zhuB4LSF3EX4R
YXzPlaVwxrXO1tu5VMHjMPPCkSsZSol6Dgs+TNOV0zhUQgFmq4e5iuGWpjcLOyOY
N9gRM0FH2eQu4d0fiKYSjHDUTYyUlW39dWE+MJu/iixOYkrriATqv/c7KbXIrwJH
tL5bebRT8Uwfty6dzQdJZTEzOrLSqzDq1O7/i0wAbHUlI09zGpBJxbf7I4AjexTa
z1XVV/GpnE9VrCtZUsPOEWqw3h2yjaVI4/bRBrm8PcdkaqkZldbdBn5G6O/IyiGi
9aO808ZbPtHUYkXiaPJZoLoRQJQBYmmoCJZsphlOhbBwCYzx/XTXFZdAf5Ro08lp
zJPyHTSibc6c6DHpmsM3tVwjQIoehmcryy7UkIwzoffSKm54blMd9/d2P4F4qdUj
DvnjUVazzvEUKiajnTvpHMHDQ17eJ1cJoueqWqQWGls6+fIbYHgZxcSddyJDFOeS
dQiMB1QNAWjRwhJhF6p+5VD3Y83+5DEFtUYEHHBvZOTNaVxTSBTJX+Sab8J+CeJi
QMwSzlg4R1KLJwVfWHbgecxqthpym6/omlTLRgln1nu18UsUsf1CyfHbZo1Eo7P6
9HsfdrNvX05FOdMPwf7gcsbSzAUYgEIx6TuXflhddNlIqP0fnQIDqc5U76wk5Rx5
jbSgMg+aEFWxxrLGvWdFJb7uIAnTYXHZ4dRgp3cUYk2mUR9mgxPNGHNdqyzuUlUb
45MwcCyYwQ7mPfTUjmfdBLgN7GUFL0m1/S80sEPFHqnOHjrb3f8fA5eI//3BYIMg
n8wi7DGcuQNljOYIlqKpIVwKUK8UDYQuV7oQK6wNREINg4NP1/F6fv12YUJ/6hX1
qf/ii+ODGefTa8kjS5IxsjLiRKMbGB1d+UJYiWjhjRWvViRoFLG4oYtmVJ4sc1t1
kF+oFW9W3gppw73zK0uYTmsEAL8Amy4ipOsP7lUrlZrwutEHV9aEnnN2uXkgxOLH
TZtaVacjZdiHnDUN5EUtW1MJJUiTwgksMWsoLq93cr4toQ7p1li5d5ULA2a7+Zef
rGs42V6Cch2ka+LBl7BEhn0HEUyirRSduWE0J944IICJAUjW7FgqRAyOfIWIreEj
IWe8gtH0U2SqlQB1p7YJlHUPc1+/D12J7yb5szJ5Q+YkVtEihR+Zd9p3b61YQ0bx
lmUXqsjJk2m7ILNrp/HahtT2qPDrBD+jGCLRf/mg3lW93DA72RFzEmtxhsEMh0Dd
jVSWx0eeh/l7oGhDf9+3XkXSioUL3QE6+9IK6FQc67OpZhNaS/cGOzmNu6yC/ldN
JYz5VxV+euyGbwH0BYndHWJbjlHx0J+b3P2AXf1rOhh/PUINxZTommTr2n9paBFH
G5kf6/JftX/+lTIotjL2XTSOYHi6WB7RWzCpSDm3kENnHJaIpEB02731Hk1vdVdD
zGKq9RfLvt8PRaDyaoNZ8dLqasTlbUXY2fI2F/GTj0t0yLvDHNdM9uOiBjH1h69z
2EiDmuaSnGihN/C+aUvmyHH4+4CAIdde40w/rfhmZd1I7drD3D/1KUVNy/bIgBpJ
fty5eGcb1geS+DP+7pBKxFRDesUJegyodZs3j/xQjnsNC3OJ0qRFveqffLmF0My9
kPdeBLHL+gmNHIkddRRXw8bsDq4KgxCD5fbSgGMe+pFAz9zNgBVGWLbVXxHSGKeP
BZenb75g5+V00JO0ZIBXedVIRgVRH/3CR7rhfCeEbKZd7tGAmGWVRyWY6RK01qs9
Iuq84sDufHVIKwgH4/ru1ucVVMf97l3wSMs3IWNRMcM/Qxs+gPy5uC53LUl2s6rl
VGijAyCwM/wozkvOoJbJolue68TlELaHKU8cS/4+a2rEfspRbHbj437Jo9cuaNvR
7g6qrBzZX/XTR1hv0ayPfflItQYH5NSlFkdYW6ypSHaPFfpLcHDWBgYgTjRa/b13
0LipbZS/X26gf0rJml4rlkj7FX7PFGsDr3bBoLV5s6/RH8Eyz91+M2sa82viFp7k
RWesC7nk8NOYLLTDs6Z2/XXHicpk/kcbw7uAO8ITRL+UEbIhGk24wWxK22fJawM5
Ih29OIdXMA25IlcOdFFP393Kb9C1BsNUmMfPXoPEsUk5SICqwMkdlaJ+usaZ2zL+
C6dmd81ZEUrOsMUZhFVs/DQYdRlA6frLKGzjMlvzfaFuIH69KPuEYdmtd3oNAQ4n
P8pJRVT9qRDN5gcGuQc8ZAZtfa917f/0P88AszUmStgE7edUZm901Z+RnIIMqARb
N7jFJmmyjxQ96glXOAG323WKUQFeROo1rhS5Jvg8zDOEEFp0MIDQ8BuHfM0qC+zo
estle71E0HxaZb53gsjTRAYJaAnH8z2x0c7Oy5mzhMWINE3NUHsd/eT1zjL3eAiw
326z9wUtY1Pz+jrdCbrs3RKIej0Mm6oQkD70/xiO20XKnQVmGhrlDguPVgUO3YdX
2RWGoSP+zrMXhDrl5uXKJGktz6X+kwyOVCX1rtY9zlT13Al0vF/X/c12G1doRQcB
DfzXunXxAjBC/hv5OUobXRnEd8hcUbacYyqzdO82mQYdesCEbtwpwgzUAjXzXId3
/fGo4v/06DLj5QLttYLQ1qCGDHTa3PwhZGGjBKZ7n1FC1yrdp9a2jw9bf/zpBw0D
YnNekuPfE3i5OF1tYuWtrNHM09zCeKT6qVWWaah6YWRxMrsgSS4I2UkaBe1T4Vj8
gz964/AFJFlYZpCNiaEebrfRqIq4SmEx0oxLRO7YiHjeTk4flU14Jac8EeXFXlag
QiEu76SuiIFyMrGOdNVKPnQc97T8ljM/hEH8hicRnmnP7Ue8tyZAVQzJIOryQqlS
wf218RcnirFGcYzrNNEr7i/POrILTgr5KGqQ3IwwLLgGNl5u8BpvnaEUb4Ef7X7j
NQmxhknj/DAKKjY1fznE1R1rvC+LF0qRcgDUKCtraxnRltuD81Vvwrn9NqX5YCk6
fcNeIHQXs2SywD9BLoRucywCfn4+NgYk+JWFiKkEd16h3I4itMFZ/xw1JzkJXail
66LV2IKgD348H1WPiTBnuRsR6+wBEjfyndK5KoMHJH+kJyNyc+wTUIDuYhXCXaEs
yD4Hb35kpTN9uL/vrlpPKlfBbEGBy34rU7m1opmGVU+/PEKb6oz/D50W8yIHuGpa
DKvK9IqGyxV8bUx5PfCmry241VbE0aYov9kcOV2RvbZTjlGEJLIpHDf7GIYUHVKu
TbFb/3e1ZIlLBpqpmPGTY/VNiz7MmrM6bHcKnjHl3KtrsTsBnKVrDrrby8DtGrxB
9WcFddjQlUHmSTvW5hlnRLySXvnuWT1utiA0xQ9ojjM4gxyWUCV7odOyqUEQWbTi
eTSpI1jwt18rMcyhAvnfaQvPcY8FH0KX+eLm46rUtad38QbyqTAarblfc8XxjA/l
OGDY18fmPy4VjLmG7DQDb8bwQxU7fig9SRXFYSshMe0w5rvoI15s8FcAvkA7NKXC
Ax96ebBC06gZ9uf3i6sOWVSPLyQiEuzMi/mzB41fnk9fYOnM6Q3AfhFY+ztIPLkT
nKuqCUDpeFW11CkuJHxGyInkvlSoHbrQc5MqJ2OMy5NT6Yg3KWd2EjvyYtOUjRaQ
xL1aQnhJEgBsQoMefJwLIcYqU7Urc6AzpTldpfgxpYhGPLntkH0uib4AiHxYsWNk
gj9efCD96HkaZzxG4/4jJanl+TgAePMiWB89M83DOtOPvYvqZ6dd5FWbkYUasq9O
PZ6E9y0t7NXuC3DeCkxF3iicxqwmohVsIuRaAvxr9SyO8UeeNMbIKyPfzFS/v5TN
7xWgdBlXAPT/bns5lMaLAloJeH05fKJsDvy0ulMIsahmmg8LfOTMj/KHj2hjSBBP
T0k9oDqkMjVlWxkBl8A6OJpQVIz1EyQBN3pB/9YurUM3Cbc0lqjySfTkpPeKVD6+
ydoh3EYFkpVAfkIfC4CxD4h5Lu/zSdYs6pCLeghJNhI/GEOdt5FcnmRPhx2PoYA6
mxYhjdcLQPtM/vepcCBkbWo3OFRvLfiUtKzCF3DU+c5lBk11QZ+A1VJexwP4yudC
6JPaUlgsxw8ZZgfv9NufY3u0PbaPTAN/BPIQTWdf9mMCORZUwoiIPg35Pqa5AzQ4
ZZkaOp3rC37DDG6zQukRMNXyu2Et/r75m0hOQufOmufnv31IKyr6HgUi+7fKWozj
Ldlkjj7ksGv/1kEwGQOrgoA1AT04v7s2X01uVOnRvrI+ezKu2wEE54arEAcyqTKr
lFA6cozUfa3bWcjweT3jvJkhjF87DFA1ELm990lp38tMesTlJBJnoEv5BcERgVCv
dn5ZvINTy3k2OfNin/Z6LfVvnhxATFuoJaXQ7eVNel4OoB5tiuXUSR0xsIVNIjpk
ugw5FIuARPj20s2CrPLnBxgP6OdhCg/Bmz2Ne93jqcgNwN9IgZsYyjrmDtjD9dci
I0MKz101P6jP0dOviVW1hb42/AIeT//qqTaN5Rb+BQNyUYdfS4mfpt3aT0ZWCQOL
d/SpS9gKIyxh35tQpC4chH2fw76plXQABzl/9/bP9Rg26mtbRV7WyfIgnkFJYUFI
ZDcLunYhUkHXQ0jjHy/Te3klOp4cU9XQvVFeYkAbcelqDUdSxUTWyTvaR67Ud8q8
4nvJ+2+kHWew1UZNrdUboDpx5TUFwI+lx/2sxdak8T4AYJ6OPiPcRFG5XgYuLvaC
Q4zGxA49bC4b94FPioQu6VVobizxUOKTeDoE66qCGzLxDj0a5oR83Gj+Uz+FL8Nc
9ZzyJ1OKqRe0nNonFUKNB1nFOYKNnxSzKYpBO6cQUQrACKhAV02PoUK0YhQSd+Gx
Mpk779zm3iA8obwryyjnz/klMzdbS4VPWs1HHcvEa1HTdhhMbuMrpvaD3eljIByo
Mt96rS5ivU0lm0GIR5pX3SzZoaPHsqS9Bk9LZcQn/DeBO7T/qZTokbD3IlUklMCg
fO3Fu/vx5TtI2C9X+juV5k2sMPFmy5HhUMcONfjyhc/tJPgglG+GdoIUhZYwrLpo
zvyhNI0Rfm4AGWjzDTvANdebGJ23zjj1EWK3/G10OA/2SZVrrNMwCPQc6RXvW4t2
cVc9AQ7NsPMyGDDaXMXKu+F1Y8bWVrWG+jTEeHpDzpz9rq3N4SSoO8ekWMEVWj/z
aDemClYo1EAaHLF2h1sI/uIXr27GM/JmENeVLcLxZ2nSKADUWhxgNeMk7Ldhu+P1
COvjOsd3AdkkFAU0rj9hwpbx7hI6h6KY+q7c1pgwcjkYhREdA0o9VgfZuiWRJ3LT
CmLy/iejJUen2vVG6ALubZy/ktPXbiRn5rlCzm1EuTRyc3p1Af2KiJ2iq+vZjvJE
tBiNs5hq92lBFgPv8eQa9zcUwD89RMCVHQ12zPofiDgo8wbXL8DZfZCmyReJAiEj
5hzPepZeuLHIdYTrbzETa2Q/HjiplYD1m+hoKUA2b9+zgsl5/lEPv3JefGva7Wyf
aPHexje77Ge1RZUZ4CdajuXkDS+GXqO/J+Am2xdZ0A26npLnW7IDI0TqqEUJoat6
P9ERgpl61YUrE9n80Y+luMk4it6bcFCwWqLT5xRQs9zIk9/FcKB3ybn7jEZTbBW9
WqLgY5IgJqCkCVNdx1ZfSQZeF/vKekPyjciwQI39oTl/mTX+HWljYpLl8NasAAeE
6O1PkRT4U86ueXhgQuQ5jDRIYm6SYlfVQUAPCdfkT4sIfUikNm/RpGUcpGr/tsc3
SdnMhOhxc8IrfqujVb89onyO0fnK6uxB6VPuqw7gSyrIELJdA3bW5uSgqjFZW2dc
BSAnXGl6bI6hFMxstw2g3vSRNCM8myxU5rUiv57ga+qAzappcP6JC4kwp6T15VaM
zG3PaEfTY0ckRgqkq44SZF8zSOxwy7Y8Z45zo4NHbcfOiyzFvBM4kwNZw5axO7kP
epXqUmlLgXd4+tbxwi0bnSyiXwKvcYxly5Uuqz2OL1OGcPLyL89vH8ce6UcdFnqT
6obAwuwM5yJ8UHJiYH63VJ+yK/eKY7QAWOrFym3dSZ3NgY0WIAm+ygtwuBMZFNYD
uAOPQ5f5k1McKSde+4chpgv/+UdCznFotKATN70xnTYlHAOy19z33UdydgPFOg1m
YI0X7m76vfH7CBv9TGynmaR5yQ8PZZcCRB9uhhtZDpkEmvBGYBGKv73jp9kIB8NX
J1MamxOQ84ERktWWsX0zxsdsu7F8L2t+GPx3kiOubwy0KKzmxSTmIaDK5BWznizJ
ZhfoWgxwCNJhwbD3+YRZ+KwsL7TC356faZvqnhxAPd2u4iF8rO4CkzBSVeREyGdg
fS9ldG5q1/YSb31AqE4QjBK8FeoITSRj4bViCbWSc5Vj1oLZzu7OtX8IuV13hj8+
XaMlUgD8LtAI931jkdm5yzsDnLq+y2Lu/HGBoER0fZ0LGVClvmRaAGmDZAdItIBw
ZNSLk6Hhv+l0yR/fP0qaHu/6iJFPpnF50ilp6iPgFT8wHtMiaIi0EvrjShd0xxJB
+7KVOf202N4nVNTQAL8pflk41dL//CgEfiWSZaXEucRy1YNCKwpvFtG1U23HOQfc
0Aszr1uarOKf4VfX/LBmAiOUR7p/pH02Un3dpBr6idGKuaIq9y8e2lc3lPtW70WY
n208AhpJO+IpI9Q0EQA5zggs4IK5CI0v/f5CaZ1Cv18m3uEE60AZ+AtWMVqAcmeL
TwGBRzZs17ZnQHUZLQPMkDq8qoQ+m7u3iPYD2zUweppkhygE9MQxlZPg/NPFtY/3
BIPhuiXBhtzlDcgwl5kfvN17ZR/HrpBYnaOir90GD728BPg5fkCfJieYModtU+Dv
xHZadCUAoyyHzYG3rX5CatOB76l3IQ08skSIfTWCvaQ+F6HhmfEsFQmHvbG7TBGF
dwsObWawuf2fZ1ktML0dwzlHIsbL6zRSsnG3ztJEQYMTAKblt4Z6BoAbRgTZnWgj
/sQ9peFny0eBxtKO4dNMmlMrYuAYcy1VT98GlpxXh6lBlVMInezwQRP25+vY3pvx
Mn5YZTXJGU5/IsufxBIDtT7PpFdReMu6+8cYj9GF3pPxj6PV19DPSR7LZWSsL8o3
ktMGZbNnjDVRm4PKKmTsB7AT5SU/+J1UfgRvlObyMQgjc6B8daLGz/ZqEz1dU3I1
UOj/cwyU7G/IvSg0CVfXwASMmzwIL1pLiNWvgx1e7k2KMwrAMotMKKpjLeDINrvN
sVskAV4UyUXvwzn+RmDM+3AuxsIHrrmJEbkJJdFtXbV4UCihbYSO0gl7McD67E/x
H+F72hd8Dd8VuUqCQGbiIrwd1oPKVj39USpQ+UwhbX4MfTkTcaHjqhEbYrOs/Dl9
igIpxQgBh529Skd4vUxlKyKTRQ5LWcvr9Io/qisehCcUMfIb4KgAoiZLw7z/QnR8
Gb4oYDDRlK3jgks/xohaZSfAe/FLn3LopAlmrcxhPHCW2bH14zyDjEkBhDh7RYkJ
2dQ9SoybLaPewt+oeRIsKIoZFkZEXENFy8fQ7o7ud9e69WyHUz7nm2e09KeipBL9
0ou2QW1eT3/p9uGND9C6w8F4tJyZDsL0DzAmgMfP4qfsHvlcWI5p1Z8fHAJiFlwI
qg2Ndg0K6z2HMM8PB15PEHBCX2Bqn1ngy+zml5GezK8Y3VP/IuKtgG3849w1da+K
+rq9sXnXd4LmCMvtr0IxgdhziMUZjkk1qqEzrisV3guTfsH2SBoyGmAUiHa5fLuB
tnnXhnhtURCTGPa6VX0AEEXcrDUlEdrcxoEQ+dl2ztoHxzrUi+1H73EVYhltgboR
BJ8tbwe0PIieIGl+D+RHUCZsA/i2Tbf8RzMIUR2tycbGrFyJTau/IavcmaCaYhaj
EoEqvafXyOJnTZH0EbKjieizdApeGzOpOCnfTLsmtQelKG4YgjQ+JW4uiBAXcmxH
bstEQOU1GbLEwKZnQeF/tvDv2PbeMUKEJ0C8rBs0ZcEarpNA+853ZEJQHQib4Xdd
6YIJvI40cAoGJeGrLvDOFskXkG24sxjDRtA7e+qfBHDUn55VSwfOFYr1MQRvht8O
hCX/5zHFdmbCQ7OG8qNCo0rxrnz7JUgxrjovUgRF5v78qsPN8OX6Jy9FvQxaCKgR
YWG0swXYzs25O8hPwoTZTlihItQ263DnK56oKGMGZ3O++56lhMaDeE1u4PUFuBTq
hu21/R0J+LF+3ZOsreGEi2mha0n1EUHH2tCjvZkBR/+YgubsUrp+ww7s+r9KjOS1
AB3+aXR0wzbvJvg9XomdgXNEio9E86Ori+kQNMcyZXgt58gw7W4p8qouqXUoyQ+Y
DJ0YPonHCg7+XbO126UqEUIf6w9DWeAWRagQk0+eT7MDveazjkSEOYQl9ClCVyo3
IuWh6RkbfX9OxILcC7rYsk3oMJetj39YTY6DQrS5xUtWqj1dFSZ9QU9VchoZoLT1
aWvf6P30fk6m+oLqQwk1uetoJeuDXxQqvx8hcfdeifxULD/epWzx8Z6+k4yOGyhE
ZiFRG38SnlaRLx4EfXTvfrV5b++5hSEFa20C5avlwSRV2sTdCAEjasY3fmEvqW/P
xYqCUscFMBxnrEQRVlNWvm6o4MjqF/bwKYOcDBvw/MOsKpws/PhLH/UA89eVO8lv
b1DdjbAVzmf9fxTetO+EF7o6I6ayq1D642TAUUHQLQCW+MX76LcV+KfkMqb02Gdc
w4M0c8g474IQDfzxDBmowyPfkJF3WHQBtBf2ybXpF1uX4cbtnDjBm1RyumNLAX+Q
CATHWS8A2tCOOzk5MgwtsD8/k+g3/s4Z/G/kwWn9uipjpWM3Vlg+SMuCpMUIwiUn
wThpQFJnCC40W5gGm53rVfQKmkXXNKGvKhwwOCWe0TWhmEtgdsoeHL/5WnUtu+P3
JVCAranGALRy8jLlS6t3P426cuL2Lme+e5fZj7OKj2oPOWc95vzWWlS6Q1/Nl4Kr
sdsN91t/+9OYBKSq8I7/1AZbvsqOCYaLpmT5MvbFZm+fcKkL4DbSO5esxb1slukn
gbJFqIwhNOGPUwG6c609X6B1hE67oKim7pU+ZBKVy+WGtk1XpjS1UqUC2dUcsbsG
3CKayZAZyub8f5jLzOLNJrplCYJu0npg3m8uyWeiW0MS4MuLoEKZprbzc6lx6IgC
fDa1w6qko1+LINn1Taf6O6YnOEnKMdoEh7u0EZ7MCu9HwDDNCBpP3nkQeU08cJNJ
yhEIp6UxYaN5BDPE2MG7XB/YyqQLg18kfiWbA1A/zwsKYC1O3WOn0avlpHH7YAn5
oqBpATtNDsbNf1dfDs1JjWrDkWaQ58XvDCNPp8t/Goof+JAe7zIL0dlBFTjn2dlk
k3UfsYcp5VeYfm+lSrTst+i0f1iuz7T7p5bQ8s9a8JcQZ0/5SDVzzXo0WVKxKmLJ
sOrxPp06Yzl5LLtHDvSsWIADyMQWnnW4bRsfFf5+u5lUNH7NgCC3tt1g0tvFR8WP
vMxDONQfEUuxC3zsZ7P6LXPxv3vpU94jVWeHaPJ8+Ht7gGcVWsozPyNqcobvq4ia
X6WD60G9qI7L1T/rRWkqvfnfdi3ZW3Jk3zDhkwSNEC3177PL+9yqayg673RAATW5
e8FF6efm3nkKNZLCNY9p43VB98QTTzql18fhBPKeApCAW+/dAfpOYRixLNF3fWvU
foTV1QuRIFK3OsM4OfKZc5wGLY3fldhbMsSwSpP36kxNdHP3q+/hbfpIHMiZKVth
WySzfMfbr+2+gwgaUWoi87UR9MNuGNa6W3vRWMUvDqTcV0mqlmQQUsWZYUBa1KF1
TsLxirpCdyXsghZbdVf7dQLAcKyQjEHAjfGp0qw5scjIngciVo2assoppe8dQk/r
iAzwcu29EZdxARI36mNyot0YtEbQ5ykI4Y7TS2u7vGEJLczWAntNCdotgqY7DWTu
aTbvscr1qWCjk7HtzahXHO5s4XrWK7RjLmnOG44AUriHEXbXYwE+98070iI3ZGIg
1jHfmmc/thU0wXUskUFUGfl8xqK0JNPVmOVq+qRULwkjM/OfIIk2jAGLwFpb8kqm
DhJ3pG0Sp/iyKUcCpJl6n3WYOw+41+w5YFUER4lE7vDHfxDBS13cyYJKHTwi1nHB
bss7fPl70Q63DksTezLuDxkdZPmzwBq1OIdi3Z96yUNmh0SBi5kDF+YyvmfIslvQ
Dr3SXGFLXCvwwdUfIPXGhOcY1SaezT/eChI69JnpirWKKDGLk+MSpPQLavoUxb4s
FhxIMg5o0AxTDkR1GAbBl6W2+1JgE1wzj7vZVcCvYp3MPzibXIhz/KjoZEVyzq1R
QCqcBKgr5TGel8t64cvzptsLo1zJhAHhOMiZfGbC+tXW49jelc0Qad5Y1q7tNB+V
HULehDwB/Bl1BwGEIiB7Jvhav9LrDqtdhb2w1FApABEEqswWvQ+C0Eixf0lgwx6z
NTSpdbUzAnFtnrSybVA29TwahB91Vj9DOdnVPzuKJaxjUInU6khyEoI1QDx3HJRV
0MMI9oSteO6/Lw9ih3OBswvwgk8p+Dx18sJgubH4uchqxTbz5ppzlV8Y0tAS0J4S
qpLFLVAqtkcUeFX/9nNLJarsdGse+3naIWitQ4rLrdqrErMXlVvtOi8WQaH9vcCT
RkkAshzdoMJOos5zI8Im5MTbruMGTAZ8OeRwy2Zobly4HUFswG03YXjfWnue+mli
zCwL0W937RnqDPNcTrlwHqdfndoLn2SsW8+ugCzEDamSjZSGffClku/JKgwss4Fa
75hl3BpVWZua13l8sGeNubz/y5QgbBjVqj5zqsPHQInu0uhg68RARRXAEyTTbfkD
h6Xj9KI1Qn9V/0nIEATJ0Y2+nU8a+mMELEXIl2wXeqzH0ypYZZgl1qZn+E+/xgI4
dNI8gFpSaxm6znTFScnShkETjec2BFhLoamzqsHPaXY95XDWuPHgerDioGwl1BOv
gp/5NHCy+1HZ10luQBqcMRUjSjGtngTjjAy3m8xHl0D0d0ZmtSWjN8Jftr11kuXX
CsHfpBgsDaYXwXw7Zij1jEmw3JPY9WRodgc6CBhY+J0oKf8Ifi3iWff3BZDAM79m
cr1KN4zWbyxrAWY9LSnRkfk/HMy1IC/9oCgmKOEBGgEX9lQTQGE07oHGm1lHWRA9
foHuBccCUTYoTTsM/6jvanSeHuWBnni23tTWVwWPZ6xLrFPeXbUu2lhUZgIvvVRL
o9XZkSEd0reS82ova9BWB9E6411JUVp3KCNhJdozJGHhwzR8HSx1Lnmd4HULoFaQ
4/hSdWjVyScFUpdr2XF/jnp8HSVVncvjjExcLZSsOAAyCq5Yi0dS2pEdV/v3R3a/
v25HhHSaZMH2uhYAjWvbGgV6sjS/BOC1Z0XeMQwTljF3u6NcCHSa66oPfu4J+6Ki
qcrb0G74VAdToCR4eqqyIOZWDhi5M83F9+OQrl31jt9Zlb8P1Wt4O2AcJ7Sc+eOo
YxEn/UGd501EH3U5u+4Z6Q2jKSAKvO5O6vXnsy+Fct5MJDsZYpZR4KkgVQPlDVqE
bY85xrhz8rnTPI8gR5EEXyLvDN/u2ieJZU6l714IBoj7fGiQfwCHhZWmzM7/MGyz
8ybNSRrp2rkIrhYepybpcvyvFoAqlTDF7JK/t8NjYBAK3/OaphTzdw5BGacjWlTH
gz6wKhQjDHk+m2aUKsXmDa1rLqgdbHiG4mVuRXYVl2Hbad8SDXflHRIJJ4EpcdWp
dOVxthwcjgEf/+8Eh/euE+9bbkTqL2dnNrEkZ2C8HkMiESmpvZ3I6uaEkzI3Eg8Z
3UTiJe3CyqYvLRyC5YQa0eYXJZm50lUQYvrBsUzJxf/a71yd9pu6CQrl016kkkBo
IGl6uhN2czmxBhumF6QDUXIHQ3JAOIR0FkApSaq9NNwveCnV9cuqMEHJaNR4eBhb
uFJksVsVb60avqQX3biYn9FX7uFrmDzVIbRJg96jR4hBGJy9WUq0+mmJhLmlgfOX
q4mug3uwWOysIzG808SPDIzWCV8bVDm/C7DB461i6RWqsnrcd9BzeF/GRRnPgEf7
bRHF1a6q+6AWjUdOBZOb8aSwHSxsL91mDaD9cJGXcfvR39D8e5XudwDMiaX+LiwN
wio01zOJwi6s50lZL1JWmO1KCQw5Auza3eYwzpJK5ExgqKrMKe7R+pxout5pC31X
BKVdM7GKYQAkwUrGfMgq0i0pi3pESvyDqfPKXwrwtmk1GBEhCeUXWT9adCYs7RcA
sLhxtJoy37SeJwXl027OdfTCjlM6+DxoFuNPbP2qpmMUro9HScrhU9inqVSuRbs9
4eCEM97J9PZFJHlceCruAJepT0F30Wy4G1BKMZGcXf8orYLQ+YYACxEcxd8W1pFX
f46VoAtGZCrmoLgJRtPjcbBo55pJTpoR3MoA7J8Cf1PAFcsSrpRLEEZQNtL2C/ug
Q2mXRY56SKJPq310WdzCtwfYnxYhNAf4yIpVBzIqZpL3fPp16SHKWkoHJC9Rxuro
/g62k6OtXVC0wbhTT1d58KCuGeik9PUHGPt1VPFx0jsNHe+2BncAIBKjtHcqx/8A
RuOvXlcPLLqX/XaHRikD/8hLELs3TMQDUbc6qaJTFgV0PKh+ylbXv8SGFTlU6pnV
mbfR1xYncdEev8GUIcGYWa1CDhEjDUKfbpPt95eRS4czoqwfc5cdoCBr3rkYdP0m
dBEOGqCkHzeI1OZq7nKZbruGPfZfCp/kj4lI6e/nQma2Xkb2hChfvwU2PfLv/chl
22NOZ3iMHY0jS5odRNeFEtjD6P/L70gOPXRnnXDoQ29SrYV8bf6qUX0241J/Sw9x
qAOWYnPF6hHxi6Lfo2avgREu09DB0/hKHoH5rSnoRwyO3B4UfnFqv34DQl3aqRwJ
pPuNj6vioYhHsWUBF+L1glTi/7/ABHM1BCKA1vUHjxbko6UgRPOXq8ziOe4Jh7dU
x3+h1mdMsBGqf+sTa9KCHkyvMwS3SJY2SU+B1ekhlZ21/FOJQsrIHo9vudLvxCqJ
Nz3Ohra+RrNRQ0wH1+b4Rm0gj2tngm+FcIxEGKbhTeECBd2LmYMF+kQxzCokmqXc
NW7C/wUmJHSs0m67nZ36L8zRI9fQUoq7DDmpAS2GHXXLs6VdiW7oKXQFnmAYHtM8
o5aUKSt5ZoTgJUw64cD/zPmUzgsvgmjlldnVO8uQukKdOoKw0cGOIFWVxV5Mrh6P
IbaWhmcpsro5GIw1/TRkikgpw/8trgjO9ZlXKI7/pCul66ROKDq+AC+d5WAWOjdy
kztAyYTy6GBGTE0IheE1CM3tZfbs+PCix3hHeo2mmvVuAGsV3qLhKlWHic6VckmA
aATMQnQHwMwYThMHXqNaRXPrIRs7QNFBNkG1vzNfCvfzTEXwAlQVCQSNeSg6k6zO
OGZKJPXx7bVvAIZS13eMDc7RAj8wvchOS/JGMRtFt6fob67Em/eahmQ4igD8w7j+
1tY0RCJN1tjIGmBP5k9gG0ioIhaTbn3wgklLshxqRzPltPR8Yggn2NDD0SR1wmB2
XanFMxGbgckil+f7KlqW0lo3ziX5h+ViAd2P+P5bXVC5G/gFBb6nP5cQEtl67N+2
7sDIW1cdMFjn1fNT4ZGn2V/7izuYg/8L3FXkhnGDQHXM0eF0V1IfqHu/jS93Ffk0
j1bY/RCv3S2JOZbtACsGMDIX0ZJIH6fRefbTjoFmL0OtHVyIckuICTzt2rpxazX7
4FIlHu+YGeWbUQecJK6+vTNDydDbxghNPrQLBwdsVYmbWmpJJDeYsKsWxkKNKx66
ULhPmImdDTj+64iFKGk2jjr+ZFzG5j1h55x0bA0qVD+X4ewnjlBbJFlHFfERa6CE
3kKu4/Vd+DCL0i5KiO01gx97Kv2mphU2kl1vd2AatpFuQZ24ztG7i/cue4o+kTGv
tUOqhE+OdAZbIXxUnKTjiLI6ZLzxRjxQhKsGhkVyo1fq35fL1hKK8VS39zZDp0md
g18ikIrw4cMyQO0qGgjOapfcBqp8yvwr072IJzSZwGih/b8HXEeVR4mptFNC9pNt
rhAMOxfXBbXqrXmvWUCWCSoVo5SORF+kKtva54tBSjmzEW4pi9ylsGCSVQSKWrnw
gV/gOmiFq0JCAEzl1AT0R6U3ELa2bnEJB18VOmqhHerRxdFlyG2SJ6ubCqN86bKy
EVdnYDqMccFzSfGkW87q+gDxF9VsCbBuSz9squTedS5FnKa7GfDY6doI99ZVupJM
uzqbxqfgSJY3jKzsDsAq+AQP5rAU40r6kA9MwQ7gxEiICXZIpRJl+v+jldkzsHHQ
fk0YXanJgdYZW7WkRL/WpmqvFoscefk/YaS8xYDJiE0ahM0pJaulzJmJWR6NpBn+
FhGPt1TmExn+J5RtQOy2BEVlc2D+UKQFuCKjuymQTI4Cgrb0bVwPDIvQqNarOmKq
ok8dUIT4SBOeytI+9XKEUQ2wiDoVgnOLWZ6DwKOnLBFJnJmSGJIcKHqZALPddbmz
yjDm714UtGLPC2yP7gR83psCiwnpV4L/gwE0pn+d29wKwNEqkBleKLyEp5Uxc/Qh
Bw8xDQre44LjjL2a7fFoYrqTuxcqYPu0ymEbK8Ve82b7HumUA0ha8xiF90Q9cHbh
I7l7xtIPCzxVjOBt6L8fV0enolNv537v3Ea0xpN3a2At1qAqI68eCCIgBpto9rdM
GkuMk8kHX4zE4raiz994VI67NrJo9eBVLvW/unoUurbKDMhuPeF2ZKGfzTBAw67k
vt+SnmIBq77S3D+m09NdYPfxtHAJyny4oCvH2NWHdi6JD5ITKRmFfgDpytuv2ZpA
BAyn5PPnmIq2QBmTPd4BVx4YEnZMGTOu91k5mHkTuQv36Ej0lPi6kzIhjAWxx2h8
DEq6KT+u8BDyIrfTynU9U95859qS5f36Bx6O0iQfLl2sOWlSf8a5qlAS091hKHU2
flanigRbWq/boRTqm3wUrv0y+/y6uYNpKnY98d8g7RVpW5Ca3Ec+g8Z0gWAQPbFm
kTul/Kwb4eNJrohHIUGCdFIF44tUBMoFUKDj9XG+Wi3UjwNDkdw16uQYbFZE/fm7
ZbTzL5/yrX/0RO2SFtMDgE6CLy0R+n/+Bu0wCW5KftXVEzs3YyD/Wgck6TTRNDFq
0LRXmDIziq92XNuR99Z4n8Myu3DVZ8Q4IEiZuUGktqKYpKeevQvDQinCzHnPCKbp
NVIji7/V1Q940mz9iSeu5WQIVOxN9nDcR/MXUs3YYfYiQaCLyYZd1xjsfYJfHnO/
/M9h/1vYyRx2XV2yMQmYxLsU2hXOZIrncB+zU4YKTdQqkk7wqNB+2Ew7OiHDrBzs
vWjBagZ6YK12u5GFcP1YjRoDD0AUe89jvw+YDebKVvRzFZJFzMue5RlzpkYVBcbz
+G4NS/Gs1K9btGHvmaO25s5ed7PdQf4Xipa0iYT+fKy3lUyRMJskWMW0N0/Bv1Pc
RUs7NnDiDLui7YqnvMc8XnnjO5buMhDcdisMIj5CF61DPNEE/Bc5LpoEkwoIkNDi
y8WhzcpTIUEG/2UjT6PsMMzV0941zogp5LgpjrBbFKLUkRvyw8Fu+l4YGKe5Qxwv
AkZh+r7LrLGlWHCy09mw8mHFXPAK6qEosLcYYBp4ivHqFpvQ7x+bHZqu/rYjoza7
Z2zmsrfoEape8+zc4+PrqLmJL+T1F/UOcA77yw2gQ+Y7ITgyEBpDO7R6/jhDlYOu
8kskWxXU68AuzHX4RroQQ32ZodpLuN2zx6ckMLdHFSqy20nMZuKGfPDz6HJCcaIz
MYNM7YWT0FBSrf/iue6IkUeC08fIeZkfXlhyYT2JxmaJ2WBGo1BXyr4nlbwJFsD1
tI6sr/9JUEeaDWV/KkKcFtZLgrdZ5i7uLm59+2qGkwE/ei22LKqVDuA2gCEtY7Xh
fQ7uCeRp/ls+sSvHqtLlJcw9xo2i0N5wR0oTZjb7PaLyIJQVpGe9HirJIp9r41Mn
eIgGME4l6OU0yK6tx33Bm02scZc2u1yL7UvZ4vGxS9xJL5lI+xZc+gfdp9kc7wiA
IOlSQZwL39VnxOSHOl/SWVz8FtB8loxKTLaEtRuu5MFTzmwhcMXzy2ARrKebaYrH
UPRFc8T22yYIYF6SkfJWXTaEraLEtj3DqIEyXgHz7Rr8EOQn/6fjtRs0UEbLLaoD
WUmc1gAI7GQ3ck8y6Ws1bz68zzBMINYn4TkJg6hrtAgLuLukLJD+p8n6GIeoPNwW
itQmFLBEu39bsk2HLR8ZTCiVw6baC9c8F0jsGsaE4ieilGdeEiizm57vjmY7Swow
WCWXsQnNf9Oiv27X6Cy4co0N5dus2otb/uWXQryzihIbj/iS6b7vqlx7jTlIoKji
OGUsCB3PEeuMcFvyC39TlRmedIhd/Dg7nQks1bo1fSVPn7rO20njP8HUuFRAjT1+
YotXxUJuT0XW1WQ3LKlcd01RRA3L9Cc1Ko2sw3qn13sUofGtilf8ixuxdOirrXEC
N+x1N0XXU4ej6xynyEyt/4AwRoxmzAm2VJgWD9OiOvBwHgRBEEqdS7RA1W3/XMe0
Uy1FbPdoxH4+At8O8XW0MfdwS0flL8WVY+7WSTvQrRnKtbrJ0M3w8dmb0wNA2oSb
WSD/WML9h3vtJ1fGTWZS2iFlu2MTwNiz1a4skUXZzf3cr53KT/aNt5ClN3ethC0E
6uIIWGGC6MSrkwktaMf9OjLVRtfKJuONDgT1KU11yXu8jWcmgwZ1Pcya7yugMQE9
UkTKJ+/pam3eV6VAF9MnanJeUJ57sKy5AjHVzSisvq1SZhvHJ8qfXQPiqrx5i7ps
cPX3NkILQLAMt+YyY9Yh4qcHu5caHXmuJ8zOoQNKULndWXyrWzG0X553WTPeHAM8
0z8qcTtkxmt7ii8xa2PFF/7p5clfhvfQbl1JdvLsWXS8U6lSw+4vghKqEhW3weAE
VZYRCgiDJFf7zcyKwUiqVQUnNJtMm488270I2oJ3x6u0lIng/glLiGWSugPpT7LJ
/CNZBQvujHAv7omt5biHSMoE4jC3ynefLlYYsghc4U8/nCKa+I9a3itXX5i/UdLs
DiB7aRb1DtBYKG14SB4O8OpxQIQgVVpUrvc+flqw1YuK7yeKc/z6X6z4NvnMNcN2
o2VdG4oHUwRTEJWoH9WcnWB/1IFx3g26Y3DWDfVVfaRgHfy3LC2v/8xgpcOxCJn5
QJyWvcZR433oI/Lwzw2LZSRl6rq4Qk2a8gafGUASAkOgsFaTsQulKjuIPmYnyIBd
rXXwMRcBopxOeF2pGQQxIn1HgWGijifSsATJtWUEsbI+D0RgQNIJTqbnrYdwHZMj
PHspBj1FRo00KFGnuxlLmKkr9bIJubE3BF3SM+qhgk/h3qRiIeyDSXDx/fRDewMx
2FpKPkUMrqg8q5Tz4rehFV65lRqaAwmilfzeilKQh1pMxiQdEr0R63Fp8TNqeSo9
YeaUIMOpwsIID7u9LTH8Vp7ME7At/QC6iVsJVnbDtBPqzUmBVcsB52aAXxy0zGWb
z0rgnSomsZymHS//n4/Eo5dC1hSZjjPt1v9rIVezp0+MK+0ASi0bEIw6nqDhcrzW
//FgF38dO+5TmIOz84aGbT/9s/hnAeV8YDhkNf6I4kxkYCrzq2ojVFRRBVR4EG9h
Ur8SFEhRWsjsY3YCZLFbULiqkvWWibBpVQjNSKnu1RZX0+I8bipiSMfSrgc+jIh6
ZxEsqYzQQqRQUvBIJynSDhVQsHe5LPWAIxJdhhL+aYo5Rv9TZEoNSzmFUP00m1tK
2xJTuNyL3wMWWjhH4mhe08fofbJUCrYftwRCcHyhtJ+2t97aSp2mcDLsvnAQW4kY
lVosH2qt8uhDw32z4cT855JAuVuwURwAMtMxxOwsmsiceGFs6EQx4FfcVIxvtpSQ
ickmtXsA7MUFDxcUobgSAPD/mDOfCXMjPZ9edRhM7HBxXXWFkmvs6ORMEjubSYwe
GshS7HDT62LFGjTup52IRib9cFh/2hNQWJShzB8DxI/ovdFUhI7ev2rc2TQiizmr
E0R5Y8ufM6sJjwOSb+xKFvbRPABXL/E1HowP1pchR+VeyxG6YnzYRR/2eqgeP8wY
vdYRDDL4TTlzdoAiTF9Dtem1PvVE6HtYQJ/vYFwUWRHRB/z0Vrb5uVeU3eq7tPOl
IrpF6R/BUCqav8u2YoKE1tbinltTMEvmbxfmmop+PbrQi/AetNvzIBW8K1FSAvVg
pgp9bSm3sHq/bBXQRGNcAgPFiNcN/riPPGSz6TJxdxjm01hd0ry2JWdSzmVlJ05O
k3ukdtePgqk48cuy+/rORxRVtunNz9qkzjgJRGReLXujEJV2N/P+B8G90vmsqDIf
J/VjItjgZMwBhaRaihuVSUDzPH/TjUdouVWGYAbEUQ6C6zGGnk9JI68OHKMSDmnB
cIJffX/XwV04qC9lE2KU069BDgY2wtFOp/t7uYvHsd7A6VnqSEarQgRmyJBzdWia
muhX+UgsT/6bmtWM7rb4OKp5bJAQg5c712wAyZERvVUc7DxSEcbt4Pvx+2WyvuLA
+v+zbBgcUapxheVyuf8BbxSXadvruMVe/rJnJY5qc8a0qUN1CN2/m+CdCvikoNTC
EwN/tyqrfFkqwFnFEuca2KdxtT3yTvlTDkLBPtSGZdTZP83QQy1tIV2KOdyw3DI+
ue1t5JEIem++tia5Qur3v45sUO6wDvOCmTUsiekC/ngMFlt+hYqS4SL+jhQdjHQO
oOq9u2ruG8j5A4b3OksTRPwg+Ml82pZZb4JIRoFVVdq+Oz3hyVHOye2vRN8S5AcI
nzC3RMReD85ZAN65A5niTxpW7+dxwNjVX5cg1b0BpZDM/deO5yeKxeDhVkd1eBho
ZsEleUMZsnTEuKFkMPy/sk5vQ6TCSYgqkwXxxcUMrhS5aEGU3S2uSEsdBDDs486h
NvNTYswCSJLwZePcBEoifQbZh6730kYlJT0VaI2aWPhdHTjLJPKptDvUXecI7uv5
z54LdAzEESO+ygNqzwatVZdbNO7PVZz/ZyPbLaur+Nmf0m8mSUYsOCSn2mguZaaT
vifjssyEjptlVhFYNAMHWG5MU4XbuJcogNj0k5KLSamj76lwdqBZ2gcshqE5lduJ
j/QR+/NzGZdR+nzTQe40yvZR5aUSr88QHwWLCafcr7E/+IdzLkcu8iZxEE3KgRY7
qPfq6kKSTa6MxJFII/JQ2XADaMUmicPjyzDC1cbzeD3DnNODUXnsLM/POtVzk5q3
1zDRQ3Ugh9bw86bfpLQ751vA2P1/DaeECkNcvT+LfrWknJp7zOMNUcZFxf9qYb1Q
m8DGMLrqLMfssdKydhfRVZZIJdqgug8V497lQDgm0Xs+3Wxh7id4f4f4Lpm3pXgF
mPBis0waHkehLrkt2OwoHioAXwdGcBrBHFCtoObaixk7iUyi8aPYRGoPa6KYv4PN
n+A2dk3S5VYw8y+0+eQyw91P80myeuKj66dQ4BSXQ3/7ZmmVrcY6UmfSx2cCJ33G
Ux+wh+XQB1KT3uKqg+31uIR8XOYIBbXwpXDT8hZITetwKZ8TYlhKeBhUaMgZ5TAr
Q+TElk5fU2nMZY48z+p4o9oUo3E3AIGQFy/AZny7BuA/DFJpmAUZm16/CAPWfi+8
LiDLCCWyD2OyiVpskbWxhFEgNt+U+lv0ni6w9jPyucI2JVpYrTN7P9S+BP9rutbo
oSAm5zPdccQ0Y1qRHttslTWjupK/rGNj93kuI9aJ6ovYGYt/uFTQdCugdYbXXN0J
OVzpeA0RErIvqQCZBT1gb3hYM4QYOlTMq1WaKp2dxbQV8YXEfY8nf9AesPn6c4LE
K3MbhGc6SnYciUIckGX4CCpVhXsIkTRsIvyD0xBswfQC6kdUAW55zQym4wg2076X
VhcR9A9mzmRXMpcBIzBOhph82WL1PgHYYtq4Ts01AqLx5dN8guxA5tM+09/R6nuX
pXdoNPLz2DoTLS3DPNXL1Zr5aCRCnrOaHIy3b+afp/Qu3nXxwIO0HOyURt4CeA77
psSf8fjWWqf+AAMiq9vahxVolgzqHspTzxB/+Ft8r92fwfjESkM8Qp287Hiz4BFS
goMi9o0mwFfjbfp3iEtzmq1qF9+mnt2bkJOOnGxsTevsvqWdK3As/quT3Z/pA/fz
BkT4DBPDmm1+T3RpvUn6XasXlZl9wW5pvPaOCp0DdZeS86pp5BsBPOQY2oYB0Cz1
YsC/o0wPj5n4aaWfvGqG4bCgDSbe0KqVlLYtge7A0jkDdjfYK83h9ab+E9IBBFWX
PkQ3myTo5XQUOO9GhnAS+NNO1YMvWTINgABoaEaxHao+lobzryhL844DyhqoGWhk
srQN5Bc6MZLC8RhVm0ggqhPWDIVkwe9b/TMSTyc7iKHS1iEnftsiJI0p66/zD5H5
P2P4Sz2brwledLPEZ9MrHlFnajZeiwCU/ifJMLApW2l8UBM5mowuntzWNMGfMCgP
LoPyaRfSmwmwvQdRZRTsYQrgVfs7scww4Inj8bzTataMRJEBSzc+hP31KEL7s2LQ
hrn+kCyVSDMRYdQwCdebOGAfhxC775JK5Qoir3w/YEx+zM9vfzXk+82ZJZM/Ou7X
5ar08wCdGFMOnVvpgCZzsA05dBEW/LgBHOpTA7J0LerDeEzzk7KzLSFR0REwkG5n
SvWu1p41UubVQpuWtO+NMIbmRWory2eFnF2TqqTyrqbBfjeiBN639nT62ey97r18
XzvKWYMQGncn2K3QYEdcuMqmAV9FtIo9JbfMsBnMhlAq4FfGZOTdJuByjqB2cL1j
xiWvmD86HiuCYqmdYe/wqGDSLwJ+0K6RPR78YCM97uL9tTUE3Tc2olluZhiB6mGF
aZ/lLGarKJ7HCfA6YYmnFhhYEprro6RlNVkqNGa2JSyX5NmBuU5l0IG+xI56fMNv
F1N4vEtzYRxcfTMziRc6WbUFfGS4sogiO4vRDd/Vn6wpUKkWxtQMUD8joXS8sC0e
L2WKuXDhoU2a9b4wZQl2F8V1ifFWPeoaU9tSAQ4utlIMESrd0RKbeRPzLgsaDbx+
MC6bERM0kIgGx5Cjv+VKgmEQNx7bGMPMH24nhnlm5+pkL4D6quQKVEKsRhK2Vx19
usk5kxFikVFZaoWJ+LvzolP3Yvqi63vnLct7NetXLs2E/mbiPDUKmW7G9YmsvZZr
aOA7SNt2tE6Gsz0byNNlQ7ahCiOZ2iMZL65YjrNRWTRyjqrhZTEnVQ5Z6XYPZ1Fn
wyvYfaZcQ4vkFWa/DmE7p8X0OiUpN5dQ3c1AdvXaqs7BkfGoTw5weiP6/H0jwrz+
3JPDlDjA73WENSBZKHJNY0mvRAUSmdkcDiv0VNRGjLe1BAlFSoBkPAtc+PmdVesz
QC5GFIelYLTPn06dc5kC7t26GTJRkFE92M8Ick941eZfEE/Gd0PRfvobTWSij4oh
wo25TLoU4IN4Zg92KUjFN5bxcx1hAjjmngqpL36q9NsCclxFiCmYz7BGgpsAqxNQ
9rphF2Atnop4T6oQI3MKnI7JyERgqH124bUM1VUf8byWMr9E2EDYF/74Bk//BOYM
oFoOI6TPVVRwNmfuVYS2TOTmD9y3P575F+A/WKNDxS4eSSmsJ2Ep2SPm3csyWdDc
jxmpOvEZ91palcX5pgnrkvG+EF2Ri0Gio0klPKyz5ucppKMoAluaE16Zp8wPxqsS
jGBcfGYHqP0GIhhxondksLxFDCvfGDLYlb9ZkQGHAm+oahUypfDkGAkTVgIYguos
lC84aIQzmPBlmTP1UE1adO2lbE2Nfti5z1jU8VfA3RGt2xYCMQaq3sRn9JFn6oNJ
UJOymxKGByuLx+OmrJ0Dv0BdZwZuS6E07F6QFEQr6BsotG3JuJU/Vf5BtaWKP0Rh
lBU8t2nNTgnPXHVgdLTEsp7AZFL9P057zCOfmn66EFjOGLW10slZDQdqUskpL1zy
DQ+pJHKo5iusAc/AhD3pW/TAM/vz7HlRIMjSiMUHrlFP3sJPGRmdGRf63hgnn7Nm
ieFbN94PLp2sxWkj0v1R82TO1BnpwYd3EC0VBxoL6Rfbo3F/Hw3LmUmbWKFrUrzk
HHX8l9vRBsm8+CHKCsf7QGb0+pv1u3FSWWPwqJ4339ldcIECyhXEujrhkJGOLB+i
LYqz4ZgUjEbAQ1uMRkUUTRGvk434eg1TJzfx5aeUl/PpOb75Cb5SodI22FGPbCvu
81Ju+5/AJoSk8it7SZgesnLNJM8Y7+7doiBvmCmTT0CJS6Vc6TqmuYLY6yyox04t
iK/IUYuCpVhNwkhvn4HOvny1OhVRTya88/FeANmqcvDDeJi62IXd1dGMMF+Ycvt4
DphKZaU+PFDWTGos6o1kF1ZnZPSUfSo+CWRCBhIZhj5tu4v2jnHfRzoK5vS3gEzw
6TebhR1J2gOqLdopOkplzZA8B+tr/Y5fcxV7KARHFwn+CwkT55tL8ComIZrrSqa7
ZQrpV1otk1rLh+cEtp5D9IhkToyjJgvXje4aBi8YvMvM16hJb3JHyuw1kG3M9MpA
5+iPVwFpYYaZ0Ec1tlJEPOeY+nZ13iSMbu7Rsi1O4ZEJJd+teQr3F35cAeyqM6TB
DHHfPh295uhwnBQR30kBukdXfeoZkBONG3CwRuWU6Kes7S+W3i/4w8e+gLlUYAaZ
gfSD9qmlHPxRWZ04oGh3E8SQldEEeUQkXh9esOaMuCG2ubYlPT/y3JRGW7P4ImD+
OiZLG9SZ1Ebs59fUky2HonzqIYsUQFI1YJ8zVhtpwu7LWjIH+BIAqa6Ik1Mqg5wK
fg3appjAzFY/Tc1qhYQKd6kgj2YEI/ZzI8L8NswyE+YtY78sRHQrnCrCsDL+Lyt+
trgVu/vrvciyaoJk39rpsQZfJr5HrNSIIambYV7EPei6BKnT3ACdEAEbuYHVMfzS
znTyaVzwR70ge3OzTzJ6bwa7Q3LzXqN4/wZ6So9pPJq82OFeDrjOLOdXIcK+HYSu
9JbEMKXT5ZF2+lv9BF3Mbe80Ugb3JxxOj0WCs3h9jGxq4gtTFnH5JgNU9F7l8rEK
L8BUrCI3Ox2DHx8l4waHjdCfmNbKoug0wLU1Vnj//S64hWUdzsrhPT02Br3hlhmr
kw6iATq8YJFmMQzlw8In1q+Rp+PhF/T8nnjM16jgjQWeDxE/3dy5+ahG7uKB/7Mv
fZpTqsYfq7ty84hUhhpedbwRectLvuYYxGA1cQU3dGqX2f8zyrZZvbYDHO/yNmB0
BkzefaG3WBu6BoSaE/MjFYvapEoFavvxTIwASvrf+jetplwYzoCojXIu6mMPaa0j
/DkJCNRDuiPT9ccZ5bFY2s7Dqv1vzR6CiPsjFJWhEJn3jsYNiVGnbRuZXSAGtN46
oXo9uAc/9FXxpOZib5flpjLHqr6Pk4/Hrh+Mzs+LdeKVTRpT1Js+n0mLC/XqjY7D
q6knDKDlUEIoW+no0iA+QkW+pvrkSJpCTl6VUYmpGYIW8b2VTR1lpHMY4gfWkQ2q
F4buuxkKaqxZx5+GkHLolr/lNbPD44eXVOwz8qitDF/IJkA6yu0UixIc74kbxXKw
AVtxK83jWlqZrBPolKiHkAnMNyhe7ZvFub16jarxHMn7xzPiggbs1x2hewdNzjhC
O9SmIqsLJWZTor3amWLJDVIDHCb/WirlFx+73PBMyek0X3ubiGog+OdTZwDSVus8
Xt/UHvkVlmeRTvLEOOytY6THYlRYFFyUTmxedkIfl3c7Xwie6OMmT6MkktJfnoKe
nqEustEsdcSuKsgrOvUloBRCkf2SV96Zphb6HpwBnfOCrpkhuEVLM6RCHgm4j6ol
OHdYFd8+FJ4yFL7wyXEh0IfJcFiPjyuhBt55Cf2iITgH21Tk1E6qsjvMsiCQzy01
tpFD9IDWXtpWl+JZ3vGH0XyoFX933qvLldl3Ux4uBtbrDXFCtEQnuVahl7Mkbn9g
GU70mPCZpIeO2f72g2mu5EQxZM1OrvHvjjKwABhHzHZ0dMTtBfioEM7qfdbcruNX
Jt5Qp2rgZGWoqFFizh1l9mbTd9SanMCU3tn49eHRWEdp2dTdYWEJSPK9UA/ohLHs
fH69dZKUTW89ys4u3qJBh6XhkC2O49Sp3bA0P6KiXTlUJqEKbdDkF8T/xoNFJXaE
MyN1b2/lWTCsrAXtom3PabRPHhKaRYbpiqu7PiEmM6n3f+YGBLDWOEVkWM5tzvMj
34bt6zUOmmPJyOjAPacmtCQgo914pyeXcNUZ7XaoGZQrJAnUfrCGF/KddlqqzrTr
LA3QnGhndlyvgxgI8aau9Xjy2FnItFX3Btqu7ks0/j0C7VNADf5eB8Mx5qZy6dcX
DfhyrfMkAwHx6ysUH8iCN56+Vcl3RwgLa3lZVHC7GBerMoM8j6jjBcWTmj5i09h7
ELA0kaMP3ZeqDF87F4HMPcbPZUeo2nE/r1+9tYOQ+7xyc1Ycv0aGoYBQ652HC0g2
CQoY/WXg2NBfn8zIEbC4wYMegUgSxg4refUsDRzcgNAtf1wevz++0ARwD7hh2urh
wGQKULkGFcCRsE036HsLAvByATpPwW+pNuojWadI/LdokCnvcNsK2dyTuC8NdDWu
Dkov1mLTYwpyFRcwGff6uLPh6eHuUFxeHToe01TUeFhmPRl2figmOhcvLYRbiWSt
zwzVwbYJRHoT5bse2cZLXho3GRx4ceJmDDbeMMHopNKmBYJvL0/jmuBfzhLK+NrB
WQvmJKwKSppxyE1TwXW7JJ1mlay5AENBUpjym4OuYlVD5H4n3v+yXOD7AL3525rz
i0KGV4BpIrdO+c3qJCeISUmO6Juj4nCyBPQRasggAyRudsbbtKScsoWiA9qaPtir
Vd222LaUvuE2LgscOFc2AO+OytQ1F1TlBSlD18hfQikAsfkA5w5ds5dI+Lp+0Xhk
EfDC+xPtY5yjgj6WvSuN0VKOHcTu5stsnwsPS7ippTFxlmOVibigpbevdxeQQ1lU
2fx2I2FIoKc0O8MSpV7NhsW8Is3VTmLuu6PQNzX6d1WcTE86ujiVaGG8sS4yXCf2
I0cty6XPfT8xEWDgRVhSwkqJdA4GC7rfCssuZiRnLg/ne3bNRkDArsJ5h2jpIWJZ
F4/ERoaRFcA4y7mBikerV862SI2PtdvKFBSLAk7vyByycH4Lp8O2YNyKNgdAtvyF
4k/3f2xH5VoH+S3SXpf+RbrgMR4FHLIUpzhmHjnXemGKnc0T4NQGb0lwWME+4RsV
3+yfB4eIQaOm+CpMgE7+4GB8XAfAPbC4mZVooZllx4wcvK9iOKa/p9OCsszxaPck
TOLx5VwZ9WRd0jdCMabmXjXtlm1Yon+e7UrIy0/tvitsFiWSv800vs5j9fRXdugZ
eqct6LV0o0aZ+zn1/Ov3aB3ww9Jghh+tRG/41z0Uynv+O5FPRfnmRQZlqMjmXwIm
kn8zPKOUASkUzKDhaLw0CGiYtyLBZA8Nrh7L8YZze17vS/jUfxUmNTQKXRoQbdhY
MIQh7A8MKypFL0nV01HoCCfWHgDT+0wO+uDffGOhfTELpOpkmVTa1ivh6aY0xN35
O00AyCAkPiUKNFiLu8u739dv7pXV5ROd4+fyn4wb6YzjcjFzQxkpZgZ4JhDSEktm
nk1r8aGdP+0cbxjYG8xFuTuwkzsuB9cCggjpGrEmQLFK8CUGVuyefKvyHnAcdJEy
jlwq4iCaXNs/JPrKVW4uDBI2SnsJZHDHANJvB3ghrIxO9YkyAdhN7d9JrRSwDLw8
6D7AJMOrljwMYYxL2NjIdnEW0P2SoYasN+dy4vBFMWGv/jySj/cmOpuE4s8zMO6L
3MylbDNAB/qcRFc4wIb/n0qTxs2TRfQNWSFqITgk7lGlhg5dhsvYKBTxNQ6JkA4A
xqx4sltE3+Y+gH24sx+wNXvnFraGeQ4rPn2y4Cy+WffFTNyZO0dTecl4Ij5qL4nQ
MlEqokyGu+ajSETrUMghq2Mmz5OlxcOY9R7AjFsX1i7KdCTfCmRisrvzaaboEe5y
RVyQaSgKkLmvrpPvjFQ21MVF5f7yt7v1hv6Fy+ppWSPP2Ry/kVqA1bJaoLKraR1q
7uMk1E1op0CYOLmAoQUkO+V4f0/iZrA15sTi/DBbKOCCBLUgYKO8G/Ilgf1O70vo
P1d9HAIxmJELgl/3KCNaxFAiZjxrNbpW30Q0KKVwFSMUbYj1VRJgIQDliuDU8OD+
sq13UjObgLxAqAslWpevfxsOZVgkwZFBibWE6DlyxqxkDTn8vyuExyrIK1vx4L30
PM3sKxvL5zgd09iiR9DvZVCSj07j9n0Qb4okkEHcUhR5aCnGwv1CVsEy0rHyCAhD
4O4EM/McaGSe9z6wzvupayKWyIMCWkExzxFD7EDGhpw/gMNaplOo+6ybga9LAw2I
CmCrI5ebqq1DpzM2h1qu2QrQdSqtzaqL98aKf66o+urB+Z9lbbYsF5S6S01ohwVV
zSd4ji/V/rw7oNydRgw8kXlWPT0VNPx7vOuzGk0D2rHx6xSAfD3ob4hDhIr1UkJm
VSGVgdPgBNWgC+NupsZHslzrTiPMwaipJaiJ3e3wNvB5N+RdKFogKXfeUQsc1yNH
25KoZkff1wGCXt93ALAp47vjlZC3FWpo2KnRVhBkxhYwU64JnuDEOw3D3RGT9dlZ
bJ/fYDL/6LQgcU/mFZS2Qg5zEZvW9DRiZ0e+Jfy1nPjzcT3MTfyu7PZi/JVUoZ9z
jp5bO9wUENxV/PbimKpcZZXYtIZL5qcLkVXohHuQqOokrcv1g3n7UZ4twCEyd1tf
LbAW3VogzsXz5jInUta0C8EACVivq3AjJS/4rFVPTiJwVyk5G4S9ztVG60LOyYqx
YBe7SxdCDif4j6c70LWt18tLbLV2mTs0yPF20UScJINkbbtPKirlVPnQAv8ycfeL
ORsK/3rXWq5F8z8lL5fnecWyy+Bt1ObKiX9JtFrahr++n9rJ+VWVaPYsK7MAlgwI
Ieyd/rAF7BmKh9PHHEOyry/vMCQhpUJjZPA97hYg/aD5+HsZAhEVFVXw6G6JzcVj
HjG2PnbMQN3K+ijK7sZdwsBR7jQmwM0wXGwaHVDFtC2JNq421fO55PuEb2vo7F8j
waFblxkp8A+sVDkRbP8sJQgzH1CQcrRs7VMjeC4p6mSd00vwWwxGzaLi7TM5pot/
pnox1TxT351CemF6zyVqpvvvi/wDDjPer+xwsTI3KRbCAuRu/eQyYunPqEpCJxse
MZJT2t1St8N2m/sSFhUQn0jmonPTyoR/JzkYuIzn1J6hDb2vxjNIlFBWkZ7Y3mgj
Uk7vmfTR/LTbwecFsXmUatHitl8lj1LVdDMvVS5Fsf5W6krnHEPl9/gMRlPJkW8u
rjsaW/UTGWU77UFXB65w3geVLhEqFjpcSFfcArLMLTbvhCrkokMa92ScQy4hPAMW
DrYLdzkmq3xejZPw6NzcfhdMEzu6NxGusOziMf79UWoDJkoLo7zQmmwM6yPBoj3y
LX8uCRtYhFqQqKbzlmBJj4/NSxdczfqjo+atq/KOuXBOslwB8tahg6Faa16Dfg2X
gYRB2D8W5ILCJgFqUPHW8brvH30QRLkI4H09IfGbjE2DCg3+AuENDEOoX0uXiHkz
NtWkJJW2xaXQL+B7R4diKm5bsOBrlMdye4jZ57VemyjUeH+Hz+htqn6J2B3p7K4s
yr9JiG4sGNYEKnRa/nsNS2SlRsBrMjFpFSn3cI7WMof0YVFQYugcTJeBGntGQ8a/
y7ih5Wfsxt29d2mHcAYBrArF3Ymd4+F7f+/0kuU3S/y0PaILCUMzIHVasSzZuf7L
9+mlC5qW22BxstLxM3eIXR5b8bCinanXItPE55Mel5U6XUp8vcKbXFG4pq5VOk6B
cb+ZwVnVsK2/D9nBsJ4Jley/Xr4MiwVRhR/bdzccOHyWlBaFXUNR4ohJPJxKvgi+
wDxAAK2jUYRsEWbCpPTggVAh+HWmcEcg/U0LH8WBak1rpfL76wF+WxUnh70cRMoP
MAH5/nZCvQEfaTCYquvCESOUJ8+g7VvNN6p2oNoU980=
`protect END_PROTECTED
