`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7i+0uglnswEEglnIiRwmEZS5tZ8bPaGi7uC1eyCGKZ/Zg6+qtMQSK8n//w6yVhg
TvFZ9HnQcvorEaawiWMa2x12t+qnJPccc4sJJcoUuZWXmyG1uT4FkoezDYuD/rt4
0HgLdEnd9bf+SCAC0RDM+2gXVr9wWu0zy48dMruJUiaU0WEdcMRd0LinRsUxMxWY
W/6YkVuFjXsi9Dw7dQNsZGrrwZiCyD2r+lpSf4F0KVMeDk3fe0zAgs7kLVaq2Ieb
Dx1q6EHS+KOJc0a9+UiO9UtZbJ42Rv1j7BdkqsDTcTaXyFrHWZFEVqBLdLXe08UM
c2FCNOIBtY8Gxn5JMAGI7WJmXJZcsZsgu72/DtlJs4ZfHTXrCiDkzn4XHnQn+zCR
OMNKvkPdeTDyqZX5+0YzcHSAUw5DGVXyKGy8EvqyxJ/cPJ3/wwkOJkHR1YkMalbY
RAShwkRWo3/VtDM6CtjMQwuEXJpYw/EdKzGrARNPznXnSO2oyENI7bCjljmexq0b
7OZuf8e3zWb4Nw+0Elyg56OKWASe9D2zQMxkKb5DipR5X16AOFIuaRHSRAWDZaeV
+AdZJv+Jeqq7PItp6h+ffufciRkmiF6QuzzNst8hpWHz+1zklfU7PJzVn+99F4xo
XRSKi1t3mJ5gythe7tneqQ1dLLoqVDjZTc7S1xcR4qmP37IHAE4NdE8b2laPgbC6
NL3pIGozG6dR6I1x5RZAcMh1/aYbjbOTBJNV1j9RLYX9T7GT21Cz2Mz3lOrgLZvk
cANMSgamkKmjYMVhAauSRVdGyDXvBns3yMm39QvzMz4Zz+LEl+y9DmYspPSinaUD
cPMC/EC26FVNN+dKApMs4dyd+p4ibJEFixy9m1LPtCF2hhU5cvSbDZJSQS5/fXzw
wEHF+EFqbBLLZVxH/KyNw4TMsBW9t1m/QjXNLDBeSBQuRfT4u/QQczISbZ4NvGE1
edQf8/bgI6LbuHMJXBu0tEK3CaszzaWcfXtGMIvaiQ+mdz3OF2zQ5E1QhRKA3Ehm
/rgcY9diDtaLh+ugrmMSO+l0dirMQiJ0SN2q4BCcf0gH3awQiZHSxGTxrtshyA6U
4ypkEWmseFT/wIWywwbICLvKKWFwA4S2u44HLfs9qfdlmZ/S1cjvNk4TgBR8D+eB
kKlRvZyjL/UEhqJuTL11HZCzswkJ9Hm6Aw9nXz5J1jzXtIVVsm+lBFXk1tHEIKpY
xsuBKn0qXYq5lWC/8Gl0QQwRrhwkEefrAave5MQcGGIL5vKZdTv7FCNeaNVF8S/v
8fl0SuyovFSu3idxFdt2guAMWV1uj9umt/R2UUd7EiKY2SJtqlUcxl6lMaPCfZzv
01mmcewRl95tB0/ihhAxAqfd2qnKPi2qHF8Ux0aXYBl2gERPT9q+41IE3xHQla8n
etn4jnr1L/H7MArKJAGrNp/IbpSpFxmO6lUt/9KUs2U=
`protect END_PROTECTED
