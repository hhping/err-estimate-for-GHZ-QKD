`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JasjVAPuvmaP/3hWu71aL3UOei1gratSzXjhdJPusNZn70gmpzDHZUYlbewonAd/
nWBPVnuEmLwFVDrIT1OoxSweLWyOXxt7EhkSzeBOUu6ErtkZv175sj2FZDd+aqlS
+Yao+Ch20NxoGHj9BxpBi0QRFCvXuxt+1LsKSCOvTVBH2zpK92wW4QM4W+WxvzN6
fQyBIvNg4rnYFaAUbtq+7VZRwzOwomfGvd5Vd6cbbL2i6dXb4j+WVZBkfEzL4K7g
1nbxPzxgqLnHf+2EiOLl5J1z/fib9i+dUz91mEnXiNr1fLspOJwZZiBuCUpATXbm
oZfEMKzIigAL60DbNWawwfBzDvDRWKj4ORHJbAysVUjwOnep24anNoWwMHmcWa3h
8E3h+zgfEDyDaGUQP0vC6S/+TiBC7yfeCX+xl3B4Cs9caO7emAfXWTblKJl3uvfW
rtTlPWzlWqAiR5ebTlucYj36j+LcCTxy3pIhonZ3IQg9JjqP/8cABLfet3yladYV
at8wiUonB4D0PVTk6D2s7JUpsbLP3FL+eYwX6tcEqA3uFsYDdCOP1sHhPWXQI9U/
7PtT8ws6Z5/iK1Ctb0rv0MooZNxFqV/LwrwDlkqSYtQyJWpanS9GNqo6OkhD6+sd
JK+ugFvAgOLpYDuaePX47Onseq+iYk/kQdeIaSBVfhQdnmqAngTQtoUFIOvt3i7s
mSqFT/uS4Jeh5SaR/Q2Lg3PDVvDF1FlrfttQyVpkqYehPew5A5MB3FrR2J1moYuL
P7dR6lJLR03KK0fV0sCq8RDSJghyhX1gTYjumT8B8Wl2x333YjHxjSpn1H1YsbSO
NlQuUo4I61C78ss1kpr0qU7B4coMFEcMo7bGrkkUgjz4lXBaU2yie3ceT5722JOu
eCXJH/SBS+vut1nijlYBdM+vus1Zu0rjHTAMTALmhJ9pZP1uWB+mSU7wIVokJeq6
eyF3nDNq8hp8dFCIM/6DDDfHHCfCnAfrlbD/2MlhJuY1q/i4KuTAmjEjg+OVv/Ev
ooGUTA+Pjkx2tApF2ksK5hbVSm4HYDf990cpG1U7+3w8BMU9LhB9K0SYUxvF+Sp3
bMyXRm+ssB0qh7bQiyYlcgxtXNybw4d1qiJkWox4pKF5xmXG9se89gd56BpXCz9l
YfsB1onwtW6O8Ru2I+hQ3ISlP8OL0bQYqssJVyt/KPnKsw0twFR9tqAOW7ba66BE
ZaLVDAxWhyijsLRLT/JG3aW/ruN2NC2sFFIZVFnl+Y3VI87m/nRJPagbvOpUQkkT
`protect END_PROTECTED
