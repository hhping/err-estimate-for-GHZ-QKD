`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fK4qw0YGAzqWo3EyZRMPslzOKGiw7D0OjXLjmBAvTtwhqPYNSGMXY/bwc2g9WUTI
1FhE4cC0BaW/yghwJKMSDVsCaLKxq7pt3U7dxBPk+0PC7HOK8PJShPTyDUVVA87r
11Oz3LMA0vqigr1515BHVr7M6PlfyfHQ/aSk0eufpTAkb+oC8uE0shKBoPTbBDri
IPkIxjNOLCV0yfVjoVmZgTrACyK2NhoO4SQvOpcaQiuKVtisrVdWIZkaya6Re7kZ
cHG6X4yk2TvKkqec9u6tHPK8bNnSPUjq6r91606R4ZsJ4bvPqFPeSBSEGZYSIFtr
XzDz+ZceyK7Lkygm5OoU+RK9hYmDvVfHeOdOy+M0tyT9qq6O1tkOHKfPV2Wfjg+u
7+UGMY7gwCCMoUljnuDI3UPWrpAETgwxwyycBgDnXYlCwdJ9WU9tjEOYEn1gKBJG
GWBL5tOTjU31s5wd3wAtB5Tasm+Q+beDUxMzoVVUFn2q4WgeR7aOYtkSdOtZHgYP
JcGe2vem+HbVZxk6b9MRVLzJpcuY5mRrdy2S31NCItLbpTpBSVD3vGeWGLLG1Lon
uCzvMaSYO5vUaDGhSZfAFlRVVC8VWjdGwiHtUsazi3hlGyh/Vf8nXxkLTrSlB12y
i6H0L0sET/0Q1uByf092LtE9VZhG8E1GFcneI9S7HG7ysqaIIcn1xyy38ifI5Ldj
u7w3S2c9R3ZgK4ZnGIlNINlSk6wR238EtirUT0RZZmetzVdcAD1sHcAV3xUHMNDg
Z8hebVynAI3WX5u0RfH+bw==
`protect END_PROTECTED
