`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NAKBFghgs98Vj0bplH7gUltKZs9C3AzOy0Xm9hyPDjmxioZwBkTrEDfxwEfabgbu
87uv/1FAoFf7PBTd5NZmbRTpnZCNrQWMQb+dJm4uV5bT38CkiOejm+w0LbZFPLLp
svW/pqpkZdhxcKs3Fn4YiuNy0gV+mLefxZp1PdD8WJRQrHMZl6XBRHQtTbuwHd9f
CT4henwBQfxolf3hw4OCxhoWqjIe3CTkB0cf4EpA+H7VxFi9joLa9CBO5CrWo3BI
VwyMJoYervQUPCt6xb249NmL3ZGEmq9pUSgOTjD4XboLD8C8sXKxgRHuwp32SMwr
/1Eu6AEngWUNXGQNRzSxuRmLQt1ID+9HjETQxzmn6trj6HATfs7dObTZCkOc7F+d
GQbCl400YbFFUddalHyIBHWT4ZBZfEH9FSBVQALGgLaYz0JLXK6QCZoWaLlixMAb
YJ7Yba7iIIE6NuChy17qaLdA/mIkU7hkbI0T0Jr7bryobzYqx489L1ukcLathmiJ
LLZJx8+qCw3CT3X4o11vEzhiLCJv1PdhaspQidYym98tnB55X0BGaRyG5adcPU1N
fYZCqntD64LQ3VKflspRqnC9Fjm0/MTqU2eFScz0RYcV0TIWD82sJ5s7UqivV/XG
Enio7fufqgcH0A0sZu8ZeU5I87450yfxmlK6BadorX0q7rzrcVqOhrszIw4XjN6h
ogfFp003EWY8Lk4U8+JtbDHdPl97HrKAnjaSp4FwptavapgR6krdpRo7fcvBQC75
afv1guY7tWNMlutDal7JmgFWfyl2nc153LzjimJM7uxOvtap1tenJYiTGllMrbMh
o6Xio6x6AhFqejP1xt1+7eboWXMXQ+4lzMA5WyZ2TkTKudbc/e7i1/CRfAgjClOV
V2dhrcXnxTfSyD6abiCUtvJPLA3WwEMQi72hd0IN4CJlFyOlAKCxI5xGlml7NFAR
K9FudPXasecQX+WkilRcPtmXXuKgZHRQetXKqQmx/lzjhjgQUe6nrbyJ5Zw2C1v/
Kch7CZdJmHypGr7m+krrhM6hu3cN/ylj2e3N1tgiOKlWzYejUo9SEPuoD4PoSgy5
FFId421zR+64SiiccZ+xn8l7sUI1PG7HUzZDqmYLbMpreTMnKBQgmlkoVHUjBiPB
rinSaAUWY6jQ9BTEyzjs8aPgP6m5X5POF5RJu6xoo0nbYvkNfMzamIqWyTVJ/wlU
doLi4Q06E/b1xdyUSsMkBriFqdSdsxT7/aR5Gzlwv1Rq7fJzZMBp5yZXrmUUm3Or
HenRxaqOkNmCfqZddoF36bs5WnxH5Ky6UeSa+H/0CFiAo94+LbhTDrmWe9XLw5s5
gRODJs+qT9dlFLqG3t3aHM2A9paunsXEwcTyePjKXrTaVj+G+MUBpg282sYpfZoJ
R8A+uyDFbXfhWtjSBKO5K3J4u5X1VGQk8xdPohAz/0IJt2JCz8mR8cvGmTb+JgtU
GokX91LnM1usqJ+qiLtU57ugwT/GnPUNYHV9qRdJIRkyrtz6ZXxWSwpPYGJeyb97
sJbW5fg5y6zsqGYx3Gmr3vkuzR84nKcZBCs2uJSRy+VLl1/tjjbQ38AxZJeQbCg2
gDNzHEBl/oopgXJKDwoR1h/mYYtXonCftVy/f+4YEsE0tvOYk2YblcY1Kg0uuWTC
GVBH/0a63u+zjxmvrmuBJLLTkcV030MY9omh4GP6wraSe+VGoFsvH1Wy7pdYH3Jt
rF+hPmAOU1ODOpLsxZd517XUD0aCFXmBqYfv42QiXAswo1RaDpgmjSdjej/ZM68Q
+3wUKugag4HgBo5kaGviGElZBqBEAzQ0Nn4hCXBdc3JEQlR2AFGY8Q1VSrwY/78N
k4M/owsHyru6ZH25lrzDmmgxC3veJmdP9I7KGu11d0iLxg1nER/DT8fCDLLNViA6
qpQjZ0LClLTJiCvSMBLhb1cYnNzBN9U+5S07uOxvRl3eCZ5Gel+3GPY9+sbU/DR1
gFSPjE6RT0nOs+tt7VzgkrrB+n0TABYbQxIBCH+tb22ajJrELDJQDHh7iDTXcrqR
Hf0wVNtD9wmpj+dH+CSXVc1JTfoLcosldLf1T/JQVUWewdAUihCPvTDdE/LdzhxA
rrJhfXXaoZCvZDWlrS+bH/Rm6uUkyRDX2KiEFuVFaIt53fDyKz0sLb95mpZmeuf0
s0/BDiqgJhTxcQY2m9JxslXV0QJoeM+pH+1hlg9ZQ+snwSgA+OOnzszHsMDJ1XVQ
huthoeIGfwyyAUSP3ZOcMHRmlsYexdORJ3uaGu6FoGAD+hKJyTqAlxigeuI9aH8C
4j1fovrPXwvo1WQldjBsJYxXO2xNpCu8REJZt5CX67NZGgrJdzhjkzhz2t2rv7do
2It2z+3LStZP6VRxAgmbWixgMpafNFQnMT5v8MxOGeK3p2NpIDnArap30CN2Cpxc
rOZkV9etrVZRb0eXIKcUpicG/2rJaZRkTavYMF3SB7fUfNnx4qZPnfVu+nhup0Yk
Xue9u6XaP2LEERzMPCkn2Q==
`protect END_PROTECTED
