`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yz8qYbLnIRLH4UPNadV069UZPvDM7P1918Z+cBKAZjqndzo7GWjumR+FWFWAZ4Nx
vXZmd2j/o5fVF077um7suJ1p5kQbI5ciXTUcwP5ovJ+dmS9Nto0e5GHbDSzuMin6
AZikbbMv3DzSk79vt3IyfxX3RST6MqNl71U52xjemv9ndNlYIIL0h86W59d0YDBs
Vqm2ywoM1u2kAD6NaD8QjqRTRcsfjvhvH14MsLtHt+zGpNr2aRawZttIKW9golWR
CKjHWwRnCEhc9oUvftP5azA/8xDAeSE7RUwHam5rO1k2jsFFoS+9mqZ9K+nLa+QK
zNCaMTVb6WPuInMGjh6bZZsb/RpiItB+42CXSd+4g+9vJ+qqA2bcyM6+4umuJSS8
vO+CWhlmdjbQvIE3qUqcDkfbZJdzD+5lMrMfJ1PCWd54pSJ7mEFLh8pns9cFbQgS
yzIUxc/MyLVZ/oEfsWD9Rg5KIOp4hATsscNoGqYZ1uzJhuSvttLa3Fpg9baWStPV
ljK1kaWkkGwH0ZGYRpQ2HjwaqOD0SyyVbRwd7WCJo/F+J5kCgrADuQ3u32hw7tVv
76S6+FKR3wHmfru3Tvc2aFYGc6GWxiTOw1O0bqS3HmZJaePmK5O9DHXCpurAkc4U
JTCK/2kl0vOIBcPP/KiWmnL00Mm+tPru1YMfCt2RHYNcKPQKif/8cc9HAvzWUCSD
6F6hZoHjlYIygZ8yn28uar/Fs9PPWWPKrvnt4lHI3yz5y4m7sEDPHouvmJC+P7kt
4Ea2mLZNGWXGMrvE0q5A3GX9VSECx8Us/xoHTpB40EQ=
`protect END_PROTECTED
