`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HfYgiQl6ytMf8vBDJDgiRmw6pctHhIiTrLVuTV1v996Rc6f76ZEr4E8Ilt6Q9pVd
fQxWiG5Peaj4lBJ0q1N7MhqsNV7jKvMJUMNkv1HBUtC1fWyD3/J72LaOX5rxJw12
PVH5yxwnzm4ab247vA5OSfFN1AyXNDD2kxG3SzcarJ0RrxsOKEYuer0nmvD4q7JB
HnN4FYabudCnM5iy1C2WPjsIKotUQM+6S0Lt7VzkLYu8h0OhSfpJglPo2/PP1H/S
SviA/mb9krtvWXGudkBJCHxhKXQCKg9gN4gH/21rJdWE1z8jpZp7Sx1rCAS5D3UT
QvjRZx09nd/+Ezy4zLipPeW1tU8gBVuMa9+uqL0p5/x8fy+YVnOMDJ2uV25dDqxi
1DgZb7P2o/6aav6srpKLLRoIZNjwOAm8m56Jow1BovkRs9B0WVjlHQGMHMHy3IIw
rAKjTl/xCCIvkwJVb5mIxRE7qU1nvAbLnh3kmYYUrfkYGR2LlunxO99W5K29c11G
Kjzm6cSnP64oPZnn5kMG+NxQppTUT1NbM9tDe+9QzrMBzQHOaGPJ0lxmUr4bi+Bm
6n97z8MM7btLbypnvOwpv6z6ns45hPW7HcX+oVl1FDbDyD0U0lzqpvTXJDCG+Mn2
CS3jK16DfV8hE8Cl8eah6TV5/DweDGAR5uzMFvyz2Kecg44NMCpNK/xvM63i/Yn5
DZ4ENfyFEi+JfVZCN4Bz0vOJWZ/VNO+GHvJnK1zR08Cpt3rDMh3kRxpREfKk3wmH
MpW/uxAFQsHG7xL0E+taK4/JSL2E8ymfwkEGQXl8FlZuX1ZyiuyVZusx2KkQtLF6
TRGCUZwuv0xbMJ/2OikluDck+E8JnLIizHRrOPhINzITU0lrDBv5IVNixK4a9CVU
S2gzKx/p5z2OOWHwmQ3NmCJ4CmSNxCI9DITTuOU9Fm0PyjEYqfSezYAATFRpchSM
B+GBH2Hnz1qivV80Uv4YD92G4dr0clnf3E4fbuz61dEIYgyLsfqznGqprM80q7Ng
JBCXsHnW88RkkN8E3jeFnskOPe4W4+s4e566a8wF+NXaSajW3Pnc2C7XBt/qFB2U
OyrC8wBia2V6brduR+algCjzsXDCyKNRUcifcc4MZfozTs8m0ebqEJzj4t/K4LtZ
KcoxoPjtvLzKYBDspAbJCZ14NBQW+z7q12QSW+15vqzdq0jDVM8tgVyVn7+icXsf
kSOm6bBwGO70knNQTO6GKmr975GSPgPIQBusZbAuZOpDl1UBX9XNHt3cLnAxTEpF
ITp0eJ4Q7F8iyglvIdAlxXJuQsBufR0T5qI6f9Q5i7hHCKBoSm1SToOYOMHP3f8x
bVr3kuidmh14ANEmSoMdzvDxLy0rGLXKuwBEHi05ANW295rD/dChZsYkEYvEifUw
6niedUnFW5yBdDb+lTwoRoPdg+ZKYbPsSkUZKGS9q0w=
`protect END_PROTECTED
