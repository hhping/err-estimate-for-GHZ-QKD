`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hai7UERGWOwnkEqbquWGERfSIucp1XTwoLpAygD2y+v41b0jMnp08uO5ICaIK9ka
xbWLW1aNjPrQt0L00abEP7UG3rPvB6MByH8+XMmWi25hhs/utZYdJo/c0fftiKlb
1vU3vtKfCGnzqKVCZP+MyhbtxOiMR1bbLNaurt9I+AfNsMTd57W4YQkHyS7ntDGm
TjkPaCisaPOJuk165cChrtzf40z21b1mV8BPHixtFGyyHXIOckO129/pzqGu0n84
P0oywd37KGjh34n/sWXDxuAl/f9UTm2GKvgl0nD+qM5sdquLjBPyI4n/jipeemZp
BfnILQiAM5mYKT6QbFni568J+GbLK2fGzFpnmITPSF+s2O5XjAWDTOmNvKcY11MR
ZT0+xCuq6X/KYc55Azd5Iy70F0w7VPr5g5cKAjOQ8TA43sybYXvlk7COf3l+v3rr
ONJF/4sQlzHSHurlsZheZ2GPaJu6F508Xe4k9ICkD/hJbwmXMjm6qGeqbl5VEWX/
Lss4215g2OVhpku8PD6dGHktlygo+RD+lerS2fTOj4PIl1V3Vs74hUJy9BkVjFqe
CfnPeC22QSInMlujnRPhAbk67UIJIy0Ca9CO4ALitNyNqJYK5uBLCDyNiICsGcpE
C120wt0hMckHfYfOQxpoGZBM+b+yvxR2tpN7Zj8STRl66fl74/ioFzJ/iQ485rha
FsaYIZ0cpcJ+ITdqza3JFJtYiyZOeoGMGdWHjj56MXRDisQFIBsg/k+ljv0op2VU
ZVRqDQatx+AQFQ84akich+m3I7buYsoQ2t8tkAOanJMyhWJHtXfq+v0TR72g1rBX
HQWXcoVkrEkt1zm3iodCTrHkJ5Sp0g+XA+cknKRgUz4oYqpdf/T/F4N/muwi3juH
oweMn73NToYoMCOnw+xdfi9/fwMX+9WL7neMA2sqFcxoW1wvoHbkOuQqOVdEVuHp
h2xHuSrS/e5HCrGx/31zdckC+IQqazG5JcfbJxBToEKa7AOQ09zNzaV3di8XGd90
oOOUPwvrXhOyn1H72D+n8vk8RXcF1HBX/pnn0QEtdrs6C5TWZc+xSrbIPT6uuxFV
kpRU1I7Gwtfzl+SmiNgITUAST0aqfDHAOfzK697NTIUXDZ6mkEFW/0OAwXXO7FEQ
cl5KGHKgUo85I3llxbL4Ybmcuem/zj3ywpdGB8NRZvM9IexVvYF/LmGxYMJ4K8YX
asSnxfa0qKXo5/KxU992BfROmwjEdCjy1Pafs3iUqNOTwLJY/jaHXQY12j0ob1B2
Jnm/z4khhYigI5izQN3M2uUzzeYmOQyArWlkyRIeaMNSazhClNGIJzLxV68ch8TN
PDIaGKiGTbCYopBleskr2bebQlCf98tWPR94OOv3FtrQK+1LnoUnjcKbMIc1sp/P
L7+cX/GZotU/4vez/Y7CpvNUYQQPuNC9FKqgQj+rdz2eKUMGfi048y3lx3AzC60X
QK1ZV4+xhw2gCBpS580w5ovjC6Ej1OMajLFZdD2eYMyFPnrfeEaw+wO0AyTYK/DL
uiSMhIh3UKzEkfZP/YlUWKz0YMF4uBd/P6nTNF6BW6SVLBqGE09d7wOf43SFU648
1uCulvXbw8n+WATnWkaMRhksRFN22Dx8IepUFyZ54itnhr7JM/e+uY2VEpScF7JN
NhA6CZroLZ1ORhvP9MGezEnL7UAJG0ayzPTWO2Jn7ewq4kTlu/p1UwuduRYIjwfX
YvZWxRxN6ijz1do+6qz3cuT9+y6bJTNsdy89/B7Xv0pb3950BT7HImKMvWimgPwE
zZ9RXdN+l8hq00i1zBCgjfxS2ST1voaebhX8M0Ao+ggcwzy4DHLTPb5bjo2rBP+B
2acj3TVPV+lSf4Oj5OvziX0/uDfY2G1pOBpI7Foq9r4jWKsTPFiAAs6KN9ShjHkQ
JuciNZyaBEShhgILwJZ1fnjIMkTKTr8mGfpS2SgbCJ5pXWao/4lNJYX5IAqTboJN
mquB6FXs4x9c/IDx//9cic7EVPNv1M4MyoE4ksSB+h9HJubjrXv3IcUhkvWxrHWD
DMroxCqfo5v/MK/roff5SgwFSyAVI66z8EhqSEJaNbs0quR2hVVxvyQY53szetqs
PJN1XQS3MX7XzQCVEJEK1Sui8xdM39ag79xIvmGhJ7E=
`protect END_PROTECTED
