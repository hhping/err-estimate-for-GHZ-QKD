`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39NGAsAIpo2HdU5xbbwV2Hasl97wSplKc1dN5Ujw5/NWND9K5W2/SkbmFDZfEdLm
LyAfyMRAlP6SRuRCFH+kI2VTpy1YV1xd3mv+sZ+8onWSzUEZUWPSdWYu3w3fSI7l
G0mq4gtlwMnR6tlbelXDcTVG1cAROpWs23RPWq55wYB2LMLjp43ZqBlHGtXbJa9t
DkfKQzDqC8fqtNecITPq9TD3uB2ICossqLBK8GK+rsJZObKap36KrWmDso9zKYil
pzElh9VlWsti8YlbgZf/Og+0LlRPbtKeCfhweeFl4airoCTIAkG7Zlk5RwhR02tK
zqS245+2rD/uIgRiPHhSLuIxkEF9e3hA9l4xg9ZUPK+C9BfoLnDlGaigZTeOf0iy
M74gKMXTV47Ua5eTVZkWeRrk2XZK0knyh21lP35RAmgBKP664vidxMp/h0U7Kl+a
u5oVikTYu0MRFlP95qokeQLsF9cwy6ifsXatFs+e8wZ9PKR7yZtIk8CTkW+b9yI0
VA49PwVkDM0cDKaXZ1zdaiTv61WTmtJATFG5zBtG7Gg=
`protect END_PROTECTED
