`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncXwjiQmSli3eJLPXtAUpp+QJZCyW/pLdAftjkAaMBrH/nUg2k8B6viO9fYfdd0h
1kQDRo6J13woShhE8bwuXX4vxBibHR2Gz5tVQUeF51B63+0jwoqx/ReLXv4bXo+a
5X1ZtAMmh6o4hHIw5fncegXbyS9dQuXtwDR4+0mwnk+MOvvdSe7Ay6leISXrAriI
kWuv8mSyuEM43Tr5hmFcTJvJVamSrdbh81FG/DOf5BmS9m4fLItrMbI5KH7iaO8g
MTLEgJA/Q0a/wbJpBBCRoEsxuDwpGURDV9vyw3+vAYoihbXqX045/uPCC6t9UgWO
qvBd96L06uHjvOnuGAe6zgjF9Zc7/cCw2wNntZObX8yKEiyodQCJaYlb6WxC0sHa
Uhu34TT/+BmH616+TVtbO/xz63wgml2VLLsCu52697Skr5udPq5cu1w91xjgWIyp
2nguoENHRmX5dWp1MXbzk3kvlnODJXGFe1tl326hPjKIVVzTq1LSrmyWEYgkxn44
bhQksGXdrKZ+UkPGDg8pTLUrOIwBj7vZUrPQYfw8IYbn6LFaMgVY+lovsSH1/1WG
BW0WoFjOl5Qtcid+bYqQKtzJp/gjL5sisFO/HW++DkSM6i10qSsltPtn/AKxdgCw
Izt2YgfmChUquh8JLcb9rjiXGLMKe3L34rJ3kFsXBq2RI5ZKjxW524uYuamBIq0m
D/9xD+QSZaJnC/tcgK2OzStXE2aqBKdNIImKb+oi0kRUUq/lRvKo8JJxdRxT5YVA
UsTDNXfj7swmOHEmjv/uTPMwq8VQSHYboILzLtRUQzATP+OCyzyNpWySRvrSOMSC
z/zGA7ODNJpQ0lAkERM3wr9MajPCyf6uCc+LFbUV10DQ/5woZBObJHnNyD1XiUfY
0rKev/2yOgrlvyhnRWOQtXOLiz/PxbACI7dSNx2P15e0d4ef8D+uvTK9w2W9Hbam
LQpYFNQbuE+gPVqduGQZGnocDOYnsYwlo0V0p26drAeJh10nGYxwhARZ8qjjVnkE
BiL5DD4JuBh5sLbX83UlIXNw6PedhrFcfXtima2JZnDSb8IcuGPnr4P9zJtUWb0w
VJn01P0aOq1LQMIo+KU4D2zKpxqqzF1qLvj/amSJPurE2uXHJK7zwV8FHlbdO8AV
fVJeJ2HGG4Jy1KvE9fyLHIiDb6yVMI4AjPxGA+xbgcj+D9Bmam0yU+MqXoG03BfZ
ZW2SycYkBF5FsT+Wbi1b22y/nbT42edccDDq2Vzd2dl56eQoKXUl+h1IhzthM18U
Kha0stUxPPEJ7NoCmFvyhyYFBX8bR0Lggp2dlZzHVgthRL3Y1nduT122hEkODobP
xXoMzpbF/zrcnlF4uXDf/ENwzc5nhUm2h/u93kXxETjz6a969HeGxtQ1DkzVLIaV
PNdEK4Av54VzP7QIBeT0euRrjMg+I4gSp2Ppi5CFMaP6jzZ77J+nQgpknHwz3uGS
nh15o96ft2sk2wz1leRPNnpljk/7SDHcUxDjzLGbGs8s9a/ZGN3+1mgSzrnvbSWh
vo/r/IgYHmS495GG6o2hYUxHLFWWD+umfYYta1rpHsndSR4Q9b96sm5+s/ae8nte
6dmXLkNG9og0ptiEFWP4Lnrr5UuL4TO3fEigcM4jDAP54nCZLdAl7AyGQBB5NaJ9
DIT4jfpBeQZPRduwtvrMomO83RA+Gs0a0yUrg7o+G+IJxAJ9AcwiUyBFwROINAb0
rwv0WxVmCkIocs5zO0W1bfjjmkklIA8tX0vqyEDNdoN4/XwzOTzBHuC6dEjL/u5L
bkrRw5UJDSFHUgSFSh+/cHlGCH9plVazEx2JSziGefGHUeJoffHOyYNAybsrpmGy
1Enp4m7pT1cqqpj7/Mgz4VKvXuLVEF1UaknrdyMfF7bzZfIvLgq0yxgK3P3Bg+Zd
XYKV70plHisQ4ONou7WtQ+ezFnOFyRA13DAjeKQyZs758vPFpObcdLRKjaerBtAi
ce1+JZAvwhrRCjhf6WDh7zdIlfpdNbj9AHJRkx25DL7J+ySuwB8kbbAxWjCREKHX
zxOgWUQpcZZ+1f7v+TB8CrPcdddbBr/FRWP33blVh9qsQ8y3Hl0AwI1u9VaOqzvE
mN/FSY6D8o6BHCrlqOex7w7Cy6w0Gbp5toYPhKQDvgPVXnqg3btY36zGfTyAy4ge
68JoEhDb6DcY13bcOw4wrjRs9XYE42NJlL6I/V16J1evKUgAj3mf5ruaou/yv6bH
ADqCWU7dy1sndQmJFDoYWtiB4+WYk3w5WV9AJ0BTISHetPhOsKOtidKidKdq6hd9
mNWo8WxDU6zcAw3DRHAW0gLsDDSjk/OgvOE4isxUmbcZpspG405dYH3PmO85hHFJ
OQp/A9kapm5zQHvwlpQyshKsfSaiZ/UX4xdEkjOpQWvjW3+z3YRIwswynL0KsVDp
fbGThgsxGh/7tcBnnFHrWrRMroY3Y/FkBi3QVsJZDM/yGaqL8mpx2pWhyGTjUtz/
PmTA2p93WoJBmjukhhNmyNYw8CmGxI08BjuQ9znQaUXRnd1QIkThL7S/Rjl0vn9+
W7bRIJzRkdJUYf6llsoymZ2c8zcWm3qqXbaVwknz3Xffs9Qm8AVM7wa656byeJFo
3+Tph4PHsbNhz7QJmfqFnOU3J8HPG4+A6LZMAhXpKOJzLDj972i7QNPmoIAemm9q
9gfgFOEHPZxmm59yft1AyomU3colCSiAnmEHZ0ZiZ0DQtnqI7oYjWJIGOksegC8g
yNowvkG8pSG5Nor5RO9D+4QMshezIqVYpRCD9ncYFEPC3zzFzQrU6kDiGatHmyNS
EaPuJnL5IDfPwdgppJt/0jSHJel17hcehzIXoR16Tr2keoAxyDJKoAjTsICqSMHH
+cgkSulMLkOT9Oj05PUOYivIPTs5C7zNEPz7yacZBTfXW/uHXJNucaSU/RUsOzuu
`protect END_PROTECTED
