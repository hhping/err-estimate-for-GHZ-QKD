`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KG8VDkg3TLjV52YYaPvuD4/xMfWoTkIVhgCqrcCzcFkFFNHqzP0xxgBrm34gAmS/
fkBwEP1mi/7bsosm1hV01oVifGde70LRWe52pEJWM53l7fVLWCR10piplfc8Zizc
wXwY2otwmjOSkls0CKOWbSSG9cRuZn334TsrrHDPpr50kkSqiHXu9grPsW9tZmHg
EIfAYQwjrM1UqVgLQV+SiZYh0NfEm5VNqNf1o/lIwPuCaiR6LQpLpgkoSnFIMjhu
5prDzt0abUKtvLBThNusxx/47p5kx2w8L+GTzruE1hKLW4ydiQAuRprFs726vaxX
ZBdlKEcg2LTJI8VpB48EgDU2XviQ2Knvaj2z6s+P6MEihOz/ig3WrG29r0zY2ABh
YHP6q2nOXX2n/D8r0fCdjT44Tqik7CuuYNn5HpQI8QusX+lAmOSC7RCSB/e8yPxs
lwwz/atPyLMOkfyB4Lzogu85ayIWeE2kjcmdXkbkXJXRhaOrlDy5dm/Js3ongrq3
PgvYGNu98fOKyR5Hcy2oTLJocXIMxM2jMRSnQC2L4EOneTSjeFp7JF5pfWV4sGqY
rsuMFLIoPmWxYQRHeh18fjwZCtmFWK86/0p3JkbeSdgyEi2eJXlSTLo/K21lNrPs
cYJeCJ3PRXyz3aUcRnBG1JtdOor9FPs8Dx66RHApU3Oqm/F4BPNjWcCW5EMyuqgi
4bT3iWTfQnSd2V9y1G9jdAYLCCN+wnceUP9Kj1ZiVgmxeIt/5s6d1/JGwK+vOphc
B6jqaqNbfGg74vh8DWWMgHXBB6SfEQBaq83k8wdVFPg=
`protect END_PROTECTED
