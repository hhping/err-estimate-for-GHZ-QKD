`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XmhfdJRFea1rqdsnCZOGJYlU3M3ShK0DwGnUTA1WFTTncZEzPCOiHaXN8/qaNNJM
Vsg6q3UM7d8gUZuD1ar/ldU54sxKp3Ln+PbYLymwNX2uFkIleZiBsliUgD8nJnW8
rXhf+SWTS1fmxCNSHvEFzHeNHH1VB4J2KVCqZi6I94ddA4B12+6ad061/rrumN2I
GeIyum9m+pvuHx5P7y/Qv7wPNNDnRFqzq6XFjM6RXLuGdaD3o3u3ZhhR3/MSYw9J
zTtId06wivwHArTkA8mQhzLU/clSV8RFt/3fNo5CtYnC0Zdg4vaZIg2LQZFE5KUL
5e0YN4XJWuSvk+7MC+tH+ttwu3svij8bz0GzDVBp/44WDuUqoIcrxABGGDG8BjH7
gcDo50/OJt+f1Z6C+LYc8uLHLzTlzKajZICYAFJ1/0RZot/AbLT+YP1RgZ68u5I6
2VN/Qa4dJNhsWBDtKHWgUrWIjUNplYrsLn645M9Z2+kec1hexN/VD45rxtElrHRM
hxgbWaqOkXKWJqnsBQmFSMZliszEd78wfYO+7z2rYqvG8ZNw6GS6QxXfFF2x1Q0y
elHQtklEN59se/Qz+EFfEEjFuVU0c7V5Ovk7X8f9B9e/5P1GLx+tYBqCDOC1AxgB
5kPoeIcBWnjZZTCPfEHAay/TJzLfnbF39tBtRto2Qx3SkNRdrpgQXx84o0Fd+ihO
uo9zS4XgnQrE0qNR/rQIf6QzbSBe7e/fVHpNtX8BwpUPHVAdKGRHEXKHfrdiYrdE
UULBc+9LcGnpNYW5oQZDUDNcwZo5VrUkG8N8J79a72y3vsro9IZ935690AU7y8VO
PYzFlJ9Q0KVQbG4+eOa7oRfDfx9GweC/NfMBW7gpe24cnWb1+rlqkTRYWsjkA9gI
2xyJjyUYotg4yYB0MWqpzg10Ypq+t8oZ9WB8EhYnahbYxmrpCCoxSIS99BftsEPO
XvmdigW5OxsjRu+ifgcuUxI5uYrYPex1Z964lMa+JBU+iSL9d17gtd/oryj/x+yr
kA9r/vozfxAJ/1anvMnIc86jkt3Ca3l4XHT4HGA/evpdIwbTgHt5v7YDAFd/cas9
ShuaRPZXkfKv+mjpcZskoYI+6cAocCFIrKVMi4+Vej5FRMxXYzqCOUgveADouTeW
F810VnsXLc6ZLfTdUeJ5RAFz2J00MuQCLl6DthIKgQYRbWmzUubKomjx3mp5z0GI
yq0IhPuPE9xnvIQ2az6oHrZP9hmDOSJr4UFiZSltCT6Cz6/O2rpJ7YLiaRPiJ7z2
cSnEsKA2u7PvybmHkOWbDY53ka5LD+pKiDZ/OfDWv/N0EqAuwnfE3g6/q8FcU5nn
Qi3AKvgAhqszRoU+CkwW7gZX2mIPL0Ho+XE2XH4a1f8HM4CDoSX2YZI/olvsevcT
2/QKTRO2hdttd8sB67YlahC1SFDxj1tewRAsREk2C8NZcN3eJ6rttsfyh0i6qEZl
O33PiRPsoPjvnYuzW1RSeBQyhh8rD3jgqup7HbQ3/RKyJMO1NO/cOQlHOmPouIf8
t5bsusFGAMjtD9MEnAAFoMLWF+OIDX9CivYEKhwWbU04dNpXj5EopdjJyO48caRZ
MTuXDud03IZqFC2Fm31eSxQQzI5WOUgt/7RYQwJgloqbK9fqZy7j2m3K19gZR2ur
dumGqAieoFUI8TxKU9A8OCr9VjpU4rfnmjyPxyWcxPxpC7p7IPDVQAl/dJkQJP0V
RgWXsVqun8H/+6r6v3J/QbyfSjKIkpP/+ZIiaEnbnwwZvy1iF01AQ6zNCFLof93G
yEWuMeXZCGmkrZkNOtMTYhVkmR75PzzAYbPj0j1xnHGjwCNcBrxe9IZWAhDbTKYN
xNyFT3WhPZwkTYq/Uf0XMIxmWpMdAnKqF6MrC2Y5NdGD/SrHSki1KIaTdR94XsLB
gk9UEpAKq3newee+AiD6TdsLLAh+FCHCkE4L8rbjG8Oqs+957+Bn2PmAvmgYU19L
iL53QdMsB3P5g4eM/FwjfC7245OHbYOzWV6fWffKq55WLEGvxLzA5Qd/1Sk7RgtQ
jah4HeomZPJFUV5oKX1njaKv8RyESBn4vXtTFzUkyZOfqw1PSYTnfBrsOc0Nc9au
7I6sytjlGOPxKgDhgHjL9+yuWdRXGi5wvMLWFHvdaRaYAdFxUHwMykSXzo39cPGG
Zvp10LMd1ZW6SPyJW36cYpqim6SoNF4X8RX1NBt/sahE6dxfM6XrtWjYfjViPoz/
mPIURVvo0gjL1NS3PlnjnBfReL8IIf+Vs5tdz4nuKl/Qv7SlCwIqzv82Y27mqvzJ
qkVqiuPEA6DXyF76hqOD5mrkBJA/UMcrlb0MGZptmShHe/RLgRbATAAdJy81fUVy
DXBOM5I28FNX/D1r024jlHC5d2cUCJIMukvs2s5Xd4yXmbpRN3HwD9JR7Tfraz/y
MM3J2n+lLV1LF2wFimxMMbA3foCiydUosZv8OeHUFvtRAWtgeF1p+U1MGNd6hMN3
L6iWmismhsbdlvxvR49EMlZA0xDJax+s9pb1Ke+2iHVIVAxAQnLp9Pp1+2xCzw1j
dlfmhCVNlwBMS+jvz+YeCXA0ToP1oQTwMqr/ePPKWpriWYcIga+RRO8JMRst3oIv
xFggslZlS7ltUsgIg8rZfcvZodrKKO5SO8eRUHAZA2v9kGAqhuAQrX9i0HGG1dEx
hQejQIylOjI1VjbWwYhMJrfQvXwRLa2DUjKXxaoQWQs3Iq/UgXF2fgp58K5hD5ou
ECJMR8zk0ruIDI+nG13m5RcbnAadZYy3aazZrRY1iy74Nyex1+ieRIuQs7wpukzq
y9D1GdmmGxwePfsnQMDQo9yjfUcUz0P1OWZrPDtJrXXo6uVd2UFGvbv5TGRUvVC8
sml2ciAsutX9TFw+/y5H3/dClsVadfl1nMRsjwXHXygpkiXisKY7TBXgtow0nYof
/T36g2IMmlBcbG7gO1eLd/q+7f0pn/g6G+4JqaXrwbfyFN5w4LR/pNBTrGYD+KAU
n+XyDMDMfRvVLcpPPiPEp9c4rm1jCqVXs4EB+IrgyrRxU6BYbzNhY05DtmNNShAE
wDsBl2Qq1Cc+2eW4huk4FkFu+dhb1bpUKPHN2tbApih3HKh1+dm1hNTJOtD9E1wm
22xpReiS6G7RhFJwNeyzOkOtA8D/odfpGsKi73P5vOIT6y/XVO1ko+NpXXCxCe57
h4SG7riUA6MHQNzhYbODutVuXnAyk4hiD34ez/T1N9AyMebybPmvyANFiejZQVby
uHC1VA2gg3atc5pnmGHJBbjanrtxzvwnFes+rVwwqUCKWEv/ng5QlN0R5JA426mZ
HIiI3IolecPvZ3xJw9yVpSKiuH5C30LX54QKG/li69U2CQB/z7WG96BLlYRh/THj
M3yQac/unxfm/fx+92izUV+lKzDUxLigH9jNF/5zrIpnMYDfsT2lddmG2PW5OzIP
Cd8B5PaihIm/w9AnNeTxLRVg6PnF2NJDDEu/YcZ/i6pkmGcpzrHlPskmtIlyfbqC
6nSSwWdSaZeAFsRBVyA4hpcbKTDxdytTNscBOFI8WPBm0sAzPhifwrSqIz/q6fvZ
NymKa2PZFipjGQrq9MKbyyYOePMhbGRo4+bAzP55sb8EXLKlYr/qATTv8pW0m6AT
nkfpU0++h/npUyaKpweUkXSXoi+9V0hE7DteRUhh7EDOLpMKwBYhG6gFKAGa1XgI
0XxzWpkxgEa6u2C9aKu4SoZAZaIWk75XpbFTjFWvlll2r/rxN1zYt1QGHwZ/+yGA
sYn8V4PXlR7RQZRaHDI/sBoaeAJW4bUTiUBKcARpkZTTKKh24j2J5dk5HGckubTE
g2/JUwDylvTahFGMeVB792iH9KrC4HBBUeIy8MEniQalBMqPl+IjoZj82R4+IuY1
jDem/K/AY8EAed5UZF29n8jbMzn0Omx5x24zfK2moy0D/L8rb9eLfXSvR3W/j+o2
RKSsOGxPTD+yltNEfih1Pr0Mzh+TO8Aej4HWAqPv791S1jmnc28PpVc7OO1Ul4UP
RaAlFzefDYL6RMTjIdWTLAlbzHQ4mC3lBpn0imVA71H60QO0HLcmUSQwT2m07XDW
wmtCKEear3wbg5wqY3FusmGXYZxjJXMMl8yRZlPuT3UcPw10BfYeMyAsSvqP7GAU
5k9Hz4hTgHc8eO9vs/k9SJwGESvaCsi4bE9XhxncLCV9IqSbVVDPDg0795UQsOxg
zsXoFMhtK7529SKb6io6WOoEUe4TT3NIcf4CJQByzw9HW+t1ZVTyarADmLThqRRJ
LrXaRlW3FnlbLdqwaaFnnlgNl+1h/x+SwtaqJYvvyatp4gW5UkgbC4ffw2ue6l62
Amj5FQxdsXMJ8c9TVp1yykdxv1UluE9y/UCUJX6o2OHmzu+vltPj7mM65MDPvgSb
JkqO1PFQPXp0P8X08VjI8gfTM2RpJg417gx/DAYM/bAMpE3YOJhNEB2xrSoG+9Rk
BnE17BxqKoYTq1OtHDfepH5U4Br5rmAfCri7OZqYneEL5aVQhwGugQNvhsvO9ok/
c5/E/R5baghU6tjkgkXLJroywEozFiCpXiJVxh9/PQ446AAEQxwJv4XbvJ8hw/Qi
ex6enlD48MPqDlIK7diVUHsd9VEnOwbMLtsPDJ8w5XEAmYyOfGXHZmUu04DRTlze
Yw0Zo/gsoEjVXlN/sSEov0L6u275q09VHhfTlXe8E62uZwSLpwl5a8M+nh38RYHj
BNl/L2cdN5j6y9sFDe3bQk7Raw40maliwxgeF1RdifjdCElUDRxmnR+iH8JgUzz1
DRWeAiCR6V7Ey5rvwpxlGAdEyS8TyHgPH6i/QjPP7rMT8IULbxa/vdgtxCL9teJB
EaZm86c07XtNo1j6Bc7NLSG1YruQUlRb7mqrTSkrjC4CePf9azEeCn1w+VKV01Y7
6eeT8M7cqPiDbwy2Upe2zEg8pR7go6ijJ9qFFZMMEC4lb8GcKb4zdKzZJDM3h1A7
N+hYAbrhKRHP/sarqqvyG6sC4It8LBwGGTZr9CP6u5jQQJWQitfoBy7oRubIIePo
dCPo5PVK4gmjowTkHZlNSsq6nhZFk88U0baH4+cPWb5tI+BA8xmf8S1p4L2vPt49
FGRUYfJxNpD9wWBas0RzQU3p09wLmNxun/Ub8elVL3oObq6q7ohv2XTqHKuJPwPO
J3eV1AAjoMIayoO2IOIyqLej7TJfTOWing7b8UkMLoREKcQb/WJmUToeTl3s/PSb
1KkQSCOuzVbPg6znqxyFTQQvacjbwxxVVIw2M/SvBwoGKjJM6772wHxFYSWGjQRy
A8TsMFxjHxLaCNiMSvKCy6XVFJiGQXShay3U+5JusOShM0KrzNkKBUa2EGbEU+iP
Vv34EORX73efD+fN3eJ7f9lUFXDUW2oKhvejgHXWairoduqlZIoG/mK2vo78DMKI
1Sv4Og8To+K1PnbrjUThNMm2DG8FJ4/fqeJKEnKrE5vxEKZElKr7V33UqIWb89uj
WzYau0A57NGgNsxEu25rmvRjKf/Ib2baW9FrqzHKY8sAMaVcCBTy26OgA/aYPDft
v3NuNmPA8rp4UBvyKBEFUEmo7SbqPx/N/elW7MeAC5Bn+lLDmikDj5rJRHo3QdTS
y991YKVntIox3eKI7EG9awoxG8jNHyPpRGDu/c87zGysUHPBM3JzTPSbx6AEHJj0
aeW9m1ThT5+OQW/uUABWXwJ8tOzNMPeWzjn5N/pbFWqGAK9EIhztwVw3DuoF/iBy
HxweZ+PuQ8LCjoF0htmMK+dkfuao14aGRvBvit8MZuQ9iPg20Ifs3Mp90QjWsNHw
I0t/fiB7eMWMRG5K8y2XYgFxov8FB2WtXDErZksAqP4HEZTyl/AlFVKj79M0dzbq
Kds0DVhoy//RSTB+uBm3GE7gp3ckR0zIT+fKXTjM4vnM8AaWa11tb6P0PujykZom
OIrgkqhVcIWMjLFHOfjMlRlDvADBFTjtpLJQHzxQm5YGZ+LYjKcZd7M4KR54hsaI
lM2AJnZ0navKPSpMOUKdkY8v3n2//q3fJbA6gYF8llCLMwDebB/y91ieYEAynszC
vBOx2N7YNV5neO+5l3BEQsMyESMvZRs3DIcgKFpu2T3JVYagClGbORHvN1/glxgb
PCTZR2a0FbmmAGnOz1PlbD4geqzAHU3i0TCtVYiQJyirlmXAW/3/Cq8+62dIguZ+
ic5DM4XdX7ReWn+Smh8BtTuVm4wb1zaKrsOsiIB1KNZ2KxtrGrVB/YlGNlTDW+En
4qn37BuRjQiBZiNSaTG2SxzWR8CgCXsfkSeHdqB/1nIsxHaM+sw5I7VGqU9su+cf
FFlBnjKxHlGuPs/TDEWd/qevGJHRU+ysrUbcuQF0CMP2rvuAnNDWWpthDr7pLX5N
4nhVSJWdDhFR+Q2qaJQBUvmopVYaTVVt4Vpvs0aQI73JEYnzsHhRSBkxIh+QsLmH
iWBlGOhUAKM/Dix8UcgmnEHXgaVNuPybR+mxkOyWY2/ZYDXJ0z4qx11chfBSnfFA
/tqnOFXnr6azed3/bLMVarChPg/tu8Tyx5k+ba+MNXYHM9BzBgAcLllhWXmSPEPU
/sXi3hjrUkIDpl2eZSYZSifsM9ov1Oz5Qi82cS02TrE0BD5AFm9KMWceRaO9zbp9
jw9qgZXMd4laRDhTMWDkMvcFfzfV1B71vEXeWTt0p9PpOoUZVGXuAiO0CHESjbL4
WOU3DjlqIbhufbB1Hq3srV4/LdlgmyVd2a4JMVwVZLwUa5M2eh2KEPB8MdSk43kB
yWpy9IuvROYB0UwNScDMQFDe51/WPIxy1XS9gbLaXezHrf95JB8Uo7qTTl2HgEz9
q2Zmhx6XeNYCnkKi4NjD3hdIFcR5CdwpcvR1cYfleqOeYjE5IAuWA2qpnQgcHyaU
nDDQQSOHmi0c0qEjXJGHembMVVm7oNHNEXVOh6rlPdARaK1D0NibKVIohfPTvtUm
f7FTeJHFn7o9BB9PMj9iaG4P0CGrqDu62KzET0R6mNGW0JOJGejDoGRB7yPmiZBz
WElQiDgJC48GBX5rTK//4zwA2GdlPJ881NsUyhIle8V9XXGP4Tl3zsIA720INwj5
9gUDN5X/nBcU4nGfZlNlQwO3CsihZkMeipPx1rcJ/3D3U4CLzUBw4DERt2zLI5jb
cMfWjks0CZCtWHMUr026f3AsK0Wgais6QscY+n9+ZU+/W/QpFqEAWX3YDwSPigW+
Ja+AcHWlRtdK+hgOMaHgvoDFVOA5QJsZKyuMgLHPfPoJpURxz23IAnWssdnWhdN0
V8TO43hJksNuYrXJCKEGpuoW56DDMcsCKhxzIS2zlCasGqxPDe7T0OwD4VGd1iBK
zC2CPIlcQ+7r0qUQ6l8piO7MtcUgE3pr3agta6hGdEc9Ya9oYdYaQHmRgwyz3Vd3
Hum+cEI+0Bqh789C5dapRlrt8fMQr21SgPJySx4IkNEZzCURL1wYjFfvtv4nBsdi
PXsnD7Usegl6VzqNCU2G90SPA9yOKw6U+cflJpmx4gDgdLu9xrHkkOmDWf7gTw0x
CeeNhS77wFZm/vs1BNQC8cqBE1MwireX+A80CLw381eBRrh/qpnMPjV933hg68CC
070X43m+m8JXHjA9aZkkE5iC8EDbjV24iopnMNNGYw200jP3MheuuRDcMgzIDWe5
g11FhiYbOmHVo9qQREqE1TPc7NKA3aoc07e0TbtVx1ly8KLjSOyjCQOcZjGaKUaw
O+Nlc+5Vjd2wwB058H5B3AwarqVbfxvyUEGjpNw9lpkmEqm7W8dJ5edwYY6+hP1h
j8k44LhaLzDQw2APYmxyzSTuyvDZznRrLJmerCzR2K38D1OjUVBm/NHZz9uXryqT
GWo83cuTEO9PPsBhQx+3hulWE01BUI7FjtZaMLzqeVNcsZJvlXRUVyqya6pRHsKi
WEoU3D3BHMXiWZXNQ+rs2tJHsjDADoWhoWaOZzsdJQDN14UGhMJe4nTW18jCHkIk
mc1g96fTEj8HKGdsCnCQ2Tqq7OlK+zzUtcPV0U4nvUp1mljlTwP22DskkyIHtY+f
CpLGF0X4sJOUi0tIUto7r0VVmAwDBXbIDTjyGvA/sMpRz1KvcFXW44/6NatY+94p
qqYhbJb3CDEGmWVMNcbZcNSOE5bw4MAypMLN0QdU6pkjhEgo6LybWNhqngQCucXz
X8erX0MAE7bg4oVyq55qIfT+9FiU8ek+1j7g6ka+NtbzOIrUNgKf8IYAcd+IL6DR
tvFzpNQuVkE2VVw5kkQVI/p5w5N2B8QsqH8sWxsRniIB1X7mrjgBwzepxX0Kwc++
ROnpNcCMip+PvXT8kC/tP0Enpk7pxXg4pxvcVl1A69emKzcnS4GRZhnbK92yLtPM
OQf2RVDJFMrhoiAfnZQoozpkz1w37XuMMTYDOE4sIS/TLX4h+DAORc3XPHKV/gJQ
9FEU2VjvUDhq9LFfEhhIwnmFY7SIayKflBiPW23ZZ+EIz6In+5PfHe+zRORyKcJY
IE4aEfUTiAOObXLtTYuQbj5fu9S6m/2+kKglkbweyDBZgCYYpmdvb7Pi+WCIIkAe
rbWyczxHwJIFKFWO+mube3/5fKmR4zQ3Wwx8UxqRitYeoI/4xOOnUHT5GrvGGFgC
lARqRPIV9nwsX4IbylLIqeQ5itxrfyTgPLNGHJ5wQ5IUs+lUbBE4lSNCtoMjLlp+
8Q4ldVf5APmm03I9O7r18qELjOMbz0YFgdSfX558THhwZpQ8mk8ZVE0JYyTfi1qg
2IwxoIhzznjmAakb8jlW6FBnBcQkkYokXrYzXQuv6rNtPAM9yQMBKXo8O7/77bdE
DXG3Xg4bzMak6aWdt9wvwSO5pmrsUSBs1nbfT2by1KApytNHwAlRKvx/CTE1qQPC
rYlhuB/Zm8Ue1SRSIQFpMX3TM6E2x0mp7ISe86NcwA9xjPxiZynDC9Zg5AegNHQi
HD4XxfitnOFzHSok6umALN9FxpLckuOeswWOy2H8mTAKhNis3eZLeQRP6pww80B+
5mEXHux5zlHWpRbGaXDu/JU5qqlKzF25uiDRmSjwZObU2BC3IO8t7NerkDyFWquh
7tzhaCziJUJpq297ZXiRH8khdFA176bIPB5OD8WakayyFlcrGmwGS0G9j86q1d/R
FJRfxknp0ObwwwLJ0WMgm1Ojq6TcGp+SESPgA+LcSS9Vuk3MoTRuK/LyvgOeF1lH
p8u/4mRmCMgnPex+Ja259hkHtvDxh56Ak27Y4/XWK/x77iDxaqIx0M3DY7N4xgj4
B7bzt2GaENuUfeVns/BKSxSttltPpQixw5mKatVfmSz3V4UyLDME9d4xMfwhWo7I
3B5ukJ6qdbG/vHZQ2ttbxxX3PMqddJFS73/jpQ+/bLf7zFC2Kds3dp08B13unJH9
Tu9YwyWBUQiCRKu/9E7zo+vPLy1sutVVJ123nFWDOpHJeCkuK0SRBIvrq3wDraQB
9LLy0WqHfbzt7ssJS/n3zOsyLt5TpqEf2aKQqkT2WinvFGEFjUiSK4cg1wD+Ev5F
buOcpCVy0asjlc4MuiQ3rtseyE6JhGuoQYhD6WJiTkvdzfAR9wK9K7QsHayhy888
yaUh60SLejXY123JLpr+Ztx61zrDLnTFpLB1NcEUJ/C5NqEMhu6NJPdvLpqCh/+R
qX8oqZEM1cNAOtLZuC9XXsgy7XfxbGou1pSqp5xfia2HwWVGPMNe43w/kIlg533D
5by5OOwbH5WupraoR84zgBY+nswLi7q6herToilPKE5sSo8h9zbx5X3FoumQXM5i
pa6KXdPGkG6je+cFjYg064r5LCTROK9LaBZ9dMoyyTD9HxQ+nBYAjqG70IutuvhP
qwJtZHNjsQQ1Du+1mT3YTt+qNL0CxQFA6Wb9TllGm2R2NXmtCNxeZtzcFXnymto6
GztfTNA+oz934+Sxl7ryyeLh3NtQX67PTlLOILeqz9o2xcuTT8Mh585G2ITOKsfz
oGAqlqSabppVx/IkwAXYHFk2yVvvqw3nqxtZXh5eVaew8WxsE9fX0EoCKhO/x0vH
9UhMdFKPfR3sMNLJ+0YY6XSXEcdKVOLNwlSuGwsV8HwwHxwM9vRizOlcpWpw3T5v
ya78VRkNZbyVOBFD/JabnPeX47hIdIMs1Xbvu7ng1Q0LmWUjz1PTHB+SUEsHZJoO
eLkpjcF4v8ovFTL6i2sZITbJGxaxj1PbUheSMqMOFRtsEy0QLwBwwOo4rClxoGSo
hysRaMGCmc43onxhUVJR6aLoQ/ZL9GIyzs3v1+uqlMIWxPNbAgPK8SljA+roWwTc
F+3Zfq89IKN2SAE8x2PYJHQFVOsV8YddgJFeUQeciYYrrJ30ExzPt5f8DSj/CmP+
vARzgFIbAyZL9eP398EZa8yvuNhTF4mBQFKQIDSQXdo8zcjVpoJrH+/hZIQN3q5N
P+g6p8CPkk+GLdSyzfDvfEZt9E3n+CILqIcB+sjmV70iZYOmrsdi1ZkPVghRggcD
XqU+YX5qNYtiF5+w2qA7XcDZPaTWJ+eXb6jpEDCsOam88N3i24bng0HdL4NNSxU6
GyxG5QoVyCNxQ8JEM7iWWD/l2zcRaYOUiQGOUl2x5sXm+ShhN44UJYt54qidRdcU
ihwuur7vEtqpKnxMl2RGdzEx6IiNWREd64gGmBwejzeNHuesDXnL1E5x+H6wXz51
CG4CdiQmjaqpQ058veEoaG3u3mz7PkD09IfoelJh6QPCKZS9ziWPM1vK6ZwR3y3I
OZ2VFqRZkFo2+8WNCRMtYJp+jU0zL2SnaAR1xAWmaXCC1bAKEyPc5xOOicZ4FxOw
r0570Y7mi+MFiMQJdpQSQVWdp7sbW4EkkIb80eyjYtfOUtGtb3t2YbgCidxZ7NPj
Fwffq6mKPi3Ftb2DEvnrB4NAJzyNMVhktqMOEy1uMpWAkjUDIU5ILihThL7g0FMo
3FddHyvlAvBcFl0K0jo4N7xofyxVPJe5PmVBw/icuqfTnGZmbvWrFC6pSLF1Xgmz
FAkqPzzDnHGBkFaFUgZPhiRKxM7ccfik9TCmczPjgBO9HIzqSXXvKwdyLMnZLfIU
nviI04kPlWfmdt8V8Obg7hoZK9sZLI7Pd7+6HVDHq/VPoCLnh13fVPlDI1oe12Mz
OWTm58jKdSMSveDj9hMKAdL63tf/HU849gFBlOWQG0SBps/hXOj9inQET8JRhXbm
zB1kWOCAun4gMXDXWQbWEU/arVk5oDsclE6rmea6bL2hKlZLISxCmE9x82fJWDT8
9o54dWdKQUgkcfBwl699UXdq9a9MlBI610ULT3yYVJTJDdoGAeYRmdSGT5nXtfWo
gdGheRxGFeWRVd56hnmk0PKca9Er0WXVlYLklXMvLDEGaLEhe/RThksZKir4pkAs
j7yjjkWzLo7dxXcJ165Zui4VavqcUjXb/EOOUqea/W7MmFsoYv1YT3HBsNoLZjzT
LQX8kVNy7l/+k6khW8thZmDDEwfCUQgrgOsN2AOz16QkQQW4m5MTsCN1wp5tlZGe
VujBLd/MBQdn0iBpQbpSASdwfTU0H6MAzuNO6QEgfQFxDhe0y+SmzfWWaFKorHju
OPp7glomhpKc5T2VyypEZeFxwYPbRa1V5G6vKTfmEevH7m3Eemx1r/WS4eYJ03YF
Z7/bAmhkzlW8o/EhRoTJs450P7gXuJs8OymXI0GqTKGlniDNxtJPws+e9InCNJP+
IDuKyU3kCN2eYNUdXtxH/8kTdE4Mpz4NgsAq9pNK7MCGcjeS4BNgJg9619V1mFpZ
Winl6PjuSmBip3TTyyeQAVxC9SGo5z2P7tEfNeXRQE5RoXXJPnWe0rdFQ021C1oE
xsoRbbEG69Mp3Tb+5AD+Hi1C1+gJAaIPlID3XsigDc6/TVIkxBXW8CKcIDcJfol7
OHcciPNFqAaYJ5PNWAxU5UT/3/hB4ZzQmOYRj2FZlFgFH9BOK6PDz15ENl76CUnx
OVYwrQlIunu0hhm06JYimNcG+O/AYHOkSn+etizt5mHOR73+BcHRKfKLCyP2zcLv
K0yQuLyBjHMVqNUC+PHhDp+5I3322euWGsvZEyy8EKMX/TmItkwGZ7D8AmgGZYPK
rn0fbC/PU+FP8RLpb3d448xZSQfBjOLhiHbvU22jFWj+RdkkflpJ/CU+d2Sw6t9a
RxRuba+eKqAtRi78fQ3sGiYWUnuDvgjBevtwdcc36AyNTJ9fxTK6cN87YL1oD7Y+
MVnc1WLuapy3Uv1M805i/4lZED1NLtCJZDPiXmUWwVJMQbqTIAd852ueENw24/Ma
UjQSMk43IVdBEGe6Qry6DYxaTrHcjTWyIMJJAcyn0g6SM3196Hyizml9TARzfAIt
vC+BTHePxdrJm7n0LPGVhT8yDbA0Q1k//TW/mFNGpLG3GszLAUaJrJ0hXR4xE/u3
u3/gTO4SXgavGA+qCR/CEKzifdSSr7HdeZk9q1aBhG8kSbR/bXy5CjDS3jFPHWco
LX1elbIp1JcXCJlAEPxsxwTOMOo9sEkq5xXyI3jGVAfJrZFhbiC/T3QKHfQhs6+X
EJzxRhyiKOK88QwFAbcvdXaOkUCqiepFxFvXrR2G5zVJlo1ghZmqgM871j1TIUHk
MjkgrIWLHqv4iO2ye/8cDl9QgaNcX0PNELT2XKJlCrtEqBvxhLdR44T4+k9cm3o7
hXi8J4cNh4RSzsWMpyGE5/hWL/isM+PXFN38CbRnBJws4F+5jtlcKvCBW+YIRWfB
xOppxeRAgLOuzrkH7Lw3HkkQlb5BEJBtGlffHmIr/9KYUkwIZsRsJPg7TwzRSMBb
OVvBz9Cl9IV86GwnmreveDCtDyHn59mLxQGw0xsTNcuZzRXdRiNXu/yR4lDf3ir+
fIpXDHozN4pn/tujs3PGdY2m5LR1r6XvWNaASruqu+5EM2fCKJyOLbIiPQw5WUqD
9Sn4WlCLkRD84SerJBV+aYmbKxpDPT7dTC2puNRnr99RTavyZknrkxRMVGxgNVgk
otyaPpjztBUfjFOoO1GCp7Z9kgXQssnFX1xe2JIHAW1/NqnQ0zVCpW7sSb5Ywlu9
fSS+2ucds5IfjGdoCVOprUqoFQZAflby4rTM5x8BjIlFR8Yr/ygJXZWh4Sqbsyzn
GAhxkbIaPsL/8sKHbOOtJye8+BWE5Yk5veu8OcaS/XABmC26FO+wSYhBayvI4kXi
cyPIKVZWnTSIOikqJIz8yAx5XGee3M+WRRTGjaNSnEFpzelfUkPdrbW8jark0PQq
1n3LrjNKusL8vMhI+ItgQLavk3wXMn2eERmsUEEtDFK5yf3ieMiKcqTDJvpDoR26
D15iKTaflIPiL2Aij9taWafjdrjM+RTKsNbTpBESDQAWGot1XkR1hs2DtGz4DGCp
LHEP8AkDzrln+zqxFOh3VxCMvRbYVtrWQyWkAKKWQIseuUXv/PsDHTVsvwoXwciQ
UAWa13bh9SRiRT8+8WZgrSkD/Dcli3e7exUbUOYyZhBSdYSRtepEWTsKawGyISmQ
KxwuIMFPt79b6Q2TaApPuGlsLcjzsxVEGpP9Lfy9S+RHybh7QZOWP03axHVthM1D
tvx5mB7asYSv2UworqP1JO+NHqYjO6BGosS6MDtLmovHux+C4FigkulL8uJAgiLt
i7/8VssgWz0GoEAtMf48UkMEhQPxP7426PGs1SLbyjw0yTNUZVS/h2YJQyLDmh/v
+6J908NvFwtqV7vJZIIl0njJPIqqMkGBhJjVGElqZTCnZsdl9BXkacLvTs+8aM6B
NX20fvKVZUat/cDYvb3m/+4oMmyAx9Of841Gxnmv9buS6KjRyW84A/1TH8cSutXG
o2KJBfjVjC6OALF9/VRnAv2braNiH+HfKL32K/R7kdxYnJy1LQMwTMjSmi58C+eX
EMNP312SXFEO4JR99kwXF2hy1S59ZpCaKs8Jk+TlVo0tvIneYLrpUaGrR0MuPKwR
XDA1DFg16O0Chsrp2p5at2gFZvc+XN8iIRbzUdQVZxQxQqtWPSMoE/dPawFgreDz
atrKi3CFuvt5qHjUmLJvXswQmN2Hg6YDkUbej29ta4jhyiTjrL3wGPpuX3iDLSSC
7ipn+Sh1sRLTPkTY0BUQ7Gfu9ANIwE1lTsBwe6mOcFK6SnlTrqKDyy2oJfpp2Z3v
9guRV/d7dYd74GIrhBT6t4WF+dkg8B32McRo4GgvRn5JJS3EmI3djIXeFGWaln3X
hBEWq6q0QvmOGlsC//U8dBJApreUITv9rjozYa+pG4A3X0yuTm6PeARg/93oCgiD
+orNB+c+pJm7KoReV3wubxEC9wiL3BWnsvkUc7HHtrrBU68jl+Rw9sSygp5tAzTD
KGMmmUH0Lv8BAke2elGaEMZRogdyTzE/3xjdzrdTxuJq6926RnshYsES26FSjV31
x0vLPsDgEcNjo8/WeJIb+cVAzB0Et+GhLZR9iqLRZUbUeN2+NJnvNl6T9a0vEYqJ
R+093Afo9HHmu3Ybh6m51SoYHAsQUneT1l/5YEZh04vvU9XA1SLfrAELrdDaFx3q
ByCKr7Et6PJc3IPjSQfyUpVRWR2bO63blwip71JWwJtl2LflCml0j0VC5Bqnu4r8
6GCIZZWRjzmQ0j1RgRF6G9b3IpNmIuiOUk4OX08ND0mVQ9pXcxN2Sb2tjuIAuTxH
Cie5XnV91weXzJCIdJrHoeKo26xtJeSBX5axe0E7R5com/fHS5zmosTyOTvycmMy
2jp/1PAaNs1Cd5Ui7IzXo8wmWGqsfMazGSF9Xu9arY2rxPp1NdSONsYwuUeSjS9j
GG/LL+MWnpmJMDEJmIYHC9mFJdiYto1PLHUwWbfTFt+trFglj8FMiC4nPx1vEL8n
s5ZYS89onq6kKdxbhoahD0fQ6dwmd+rW14y8SyHosMIoEWEcFpdudR6j6puN+Gqv
PL69f5DRCmMJS9uNswz32/g+qRnwj/j0kVlpOJ5tNNkMDaKRakjN4go4W6P7HEk0
YPsgygyH8bUADkAbt61QIpa2gKwU09oCzSmELMaEwiskcSHiOhOm1qMp+D6IJheD
XsCqzvGGDllqjZ0djl/bErW4BmRgwYajEgfmkW9iLXRLbuT3RRHxkLVUr/XNzBNI
BB9DEqh8OXAFNiKM77w157c1VEGl6JJU52GqTgO7dPwT2fztiSQPaLwEhRb0hFqR
b02A5xOhjDCDQkO/efonOOxXYtakvrPRAS9w7oo9sxWGuQQDGfC8Yc4EXqyDYOl0
orvHxcAM7mq0wX/cN93bpEn7hRV7uJoY9QzhcYcoLl9qhGRHbOEu6LvOhuIEPKYW
5Oz5gYS2PuUIWkZZ6Geqpmzd5SMqlWqp7txH6WYunkdrIGtK8xzfD/A7SMwg2ITG
ujqNKrWN/SqkFYU9a7RB9t14EQ7rlCWeco3FDTKBJZVXfoIffDHPxUBZvbJ0uOS6
Ti0Xo1Zw+awCLPtG4Ll+hPU/9f1WjU2K5pjD2nBlwZ1tprZ88xJ9gWyZuFkz9Vzi
uU+YS67HMdIGw1VQ//+SVpwiA1e/qNZYadzhXTv5QG56aGGf3nJk5kAF9jFffx8A
ejRSSN62xO2zYU/OOKp4XTJTYrNaDNEjEQbo7zts6l+kFS0xKFx0jMbGa/D+H/PU
oz+q1yWie+AtEekl58IeTpCsmHNVvd1GJM1QcbFfC7KuKOCdnpC9xHQuGxVEWH+u
JWngCk15ui4TmmcMSPbmt4d975Y1OWfr9niM+MtSsipFsoZKK2R1c388lPE27Yz0
Hl42FCUAmJUN1fziYp8gimMA/eNb+R35S0vEfhPbIjUu9rrJO+j/mjFVQdJ7Q8I+
6eCtYYVRT6e4uI4wrbNLFzWNKYftDgEKfJMi+9sflvpDYlz6saNOzoTxn1xeKE+v
bLYnTI9gn3TKlENNzspjXlvfRZLyv8xCECeRBIlqyDUMQBsz7Q6lERxc0ot5YZrX
kVtqN6ftjT7kt1O+70yCbOmlwKanKFi4MutjJGZYPjJPvCnwH2pfDSrmPU5dVaJz
1FYa/txpNbagIXNmFCnBm2W6J76Tchl1x57qKj+Qv2QgbyfSTToxXZrw5GTVeUOl
dQBnmpaOAyMEGOJ2swQHHCQgAOr86U+x9eNjQASY4pnnjui58VpblTqkIteEdqb0
snR9shKjepEtnlsAKKFuswa72W5i6jfb1YJ3seTE41RNNU8vlPezI5Qe3r9PcGT3
tMCVGcJhtz910yAg2H1P3OGP/5U19Yq4WI79sUdOeL9rwe3Bk3JcEj6azfBTfrws
ksbabBS5+iKfA116yp/xPYNSENrbeut9gR81hvxA+ybid6Sc6ZJtRASZpq0Bxy2A
T910hBQAPfcNwPka68PwriCoqygETRGQbkfcPEJwJD+GP/msjBHaVgQmzNLHocbG
BsPO9i8KU7jatNFB1jjtZJpuNUHrXGjWTuAwAQntfjP2AJrzUdm2UFZ2GwSeKTB5
lvytp48tQa0dFmur8oPvbu4zG7lFiGk+GQMRVP4aCgd57Xjm1o/E0uCMVG12Z+Xa
hLNluV4H1UbxZLJxNeHLtsueyK/oOSzB1lUXJo7vjoMnJrmEACVvIjZjD0lGL66X
n0VeMYZ6jbict1hubz21ZctuH1QtkpbPhC2veFa8bjQBunFk2QNPgjH0vJD04eMt
1CviCmrG4vSSVlMVPIhEcOcM1IW8tw9gJtpd5RSmih2ANgf9aybx7wUvyaY0LOku
ZL/Go/RHc5US4TqnkweqGOJjChzoA9wfyKtjh2QFeOu655xLQTjKkDQI2egYdyZR
ggPVRQ9dfZoC8Hw5B42paPzjWfkGCIakUM7ad8Djw9lK5BjvNoGKOrypF/sTAeqv
PbZruCrezoaZ31Oa+Gv1+S6JSnrq+GDD1gFVJD+LBf9bVhhyW0PlgeHHzoGKQU8C
CS5jsFMr+cvlRtpsLklaF5g2XVlHCfOnWDIgg6CzHBwNU0If4BRansNM0XbRpRor
mGOYIbY+Hmas8+/PXaGu2r1AYv7K2E0umru+e5lngaA/dswnho6p85u06atECsQb
A5RMmQNH3ZlESNIuitZe6uB1UaBaB2FJzv221ro5fvl1jyrtRiOM9QTlyl/DB+0L
OIBdFGmDUBrYkefzVEDs2dvUym3pAoq0IzZo2+ZTJ0zKQtiC3yX3i8Rs3NxJTH/O
t5oTUTcJmI7qIh7Lz3zM82vHQKnDLiYoip00Bn6y2ILh3WOQ3Luw0yLTL1OkNB2i
ONldU1ZPsSrIQ/8ag0QTew==
`protect END_PROTECTED
