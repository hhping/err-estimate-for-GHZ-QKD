`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQgLeGi+v4DLNyDy+/xCi5HJAt7x0dFx/4Aouscmk9V7ZX1jR7/L9XHXx/k9IHwR
zrq5YA7hsTmbRrhfCgDOQrxmzs0hCX+XhvtEtKisFGYg5S6dLRryMpDOV7WGiEPa
54NqdPTUIFvjRA5QOG1j76InjOMzzpfgmdMJf74pa5ZBuQDl47n3ZIhz8kfnPbN+
/q2nNYopZpCYYEFl10c93bOGh1nFgyuc0l7oKcBOdMKFfd/GqMB+KXlxzBJ+RXrV
v1oEOfsHQyOXsrhzTUaUp4OltVZtlKrnhnpBW4b8pHpvqt2aiK3hQnavY/CAStt8
COKsqzPzt2qSey7IV0vYlPDki5J8TIdcCOOYdyR27UWlxkTU1Uqk8rjxDCVMXq8Z
K12zp6SDGR3jWaNumhoSFArffOjb+pfXzkRLda/2iytactRXNvisQcwUqIl7P/9A
BRvXxgbX1lsbdDyVzb665ES8bO+1cZIcUgtTsnzTwaz1+aDPl9kTKX/h/4LgYH16
uV5W6njTVZalboz1+9uBpKI65re1wKn5OGUush58YyDDej0rm6tBzx+RMYXccq0U
7ARQvgglyC0+A1I4tlYISM5fUPySS6tJvhknZ+SVsYVOYvgYq7JVz3frrFBf+erl
4eFVqpmu1u7bU87IiWdmVKZAMFilboY7wF+Ql06RG3/cKpn44KR29edWokfetCrH
iNQ94uXxcSmtXQWr2YiXDKqLTDF+uxl35JY7lXMrU1cMlpTt1XgdaseuPYAMlGwa
IJTQsv1vLbj/2DmAvgRKJFOCuN3gHykeeBW1noTHhu8K4RLvMA1iMimF+eLlMabe
31Wkl5XEOGp3IVBHMoLM4qFy933rY94hYqK9OEZFo3oWz+c1beMn4G23NnsG6Oep
i+FisFUh9HaRBRKrfPOxwaSE6SNdkms3odP/rsPAaIdT7K80yM0hvdGNL8IFz9lm
RNZZNG3/XQmbcfGSe9nzMyfJOUiMRUv/qg05JbPbXm2epqMAGBZ31oLZq/flzlVT
7HQ7bsTeyiadjQRujZN4sB0JZSVtk8L6oQv37d2Vh/TibXYBnc8m7Oxrj7tEV7sp
21TQCZgLKQUzkNXvErDhXjwjEDfaSI/RzBY7M7FERJNza4XItKcGR8XGRsaqF12v
JP1qy86Vfva1cbFyh9Nck3RykwQvow2gCzXa8WpjEYS8hzxHlqEyYB+DCeD/B8AO
VniyUZ/AK9NFyXCQt0P0/xixQIW8deFNZlmgooMmB1V5mDZwLML/dfjdEsOGxxhM
7cJSPoyNiiBR+IOjHg/oErlckgaSqB3LILhWUWKK/Z0wSI0EaPc7uKzreQzP3hVk
tYYmAW667/hCLAKpcXisxuB+FwPWdhOLPTfMRh1oMRZATyVpl6PojRuJtpX3ixe6
v4kOkrJCKXXRCaWSJz+LV8LjT+3rU9i23UeeodorbVnvqwKvNGn5+dblLrCXQgvp
m4oDKKSyNk6zBuwXQ80ELajgeUzdyV4FcO/XQdCaW1qq3lCJ26RlRLmMxmMFk7rM
Ux1zaLut+hq/rLZ7iAhN0ZLLvhDgZkCKyLTxyDCueXQN/IDPKkAusZBwX8DNqfWR
6GvNL2b2qO7p5KBWGXneMbHm3Ue4MmPZcSIcGKC07vsKJenmtyTgi2BRD14dXDxC
FCa0DQXig4MqE7l9OCslDIA1WNIlKrcdYzFBENV28xzurNa438BhQB8Y74Rdbisv
IES3njRBEtiv/QO5BuiJPPH0+P7Vdw4KwCztZbXTNSm0+0B72Ohnv7f4x2vb+kSa
mahBSwEQvwdSGPwXCTRCGvjtQATuV6+hL1gu7s0NG8QShFhv2mIasxNj8Oae5MMO
2vx60MUnL0TnqIJjCQb8HQhHfo+buaAFe0EUuNyXkjElr5YgxfdwWnWDLrnj7RvL
8qElKjPgUNcJxPKhh5xsJUx6DVySK0TfWoIlwqstrBGyt/I6RyfxPpjTYK5mU0MT
I5YanFFHo4XgdvGiY15w5ClIqAEcQJw7khf56BbfbnTzehLiu/onoHTXOFTgW+mw
l+QAK0CkQzWei1tGn9OKy7hlPvET3AFAbXTp3lI2TdOwC+j6uTLnvXasAWNAMRQF
e9X2YzXCowMBFJZdZ04BG+inv1h/SUgqtFSxGegCRrgcgE5dfF+FUUYBV+oBOrgt
yM0B+Mj/slWOI+Vzxt5N61IOB4l68HKSv7Lj8L9SNwhkwt4QCliPWeZnFfYycbRD
tHA6iU7SRpZu0a4ti8WZeJChwmfXRVRAPg26Uslh0oqMQl/piWvOErayqxdojjUU
jEStiHJFXa04b+P5HVE8X29Qn2rMZCB7wWiWX+djzQQzPea0B+Mgl+LQGI1S5sMo
n8kmGB1BxqYWAWnmxlCvbzxJuj9fw2ylEK1eIAaz+sa+qVFlGxZcSPVsb8w9QRIq
evFj1zDJ5gZhvkZZ+7fAVeU7FHX6R3ZZRXrbXXHrECbSJSen94jVZjET4kb9OdT3
q4hYBQHcncUEil9Io0Lf/qVcc4VakryS5XlwDpitxf7wRpMBeli22nbZ2ImILfJn
eaNTWreoaTf3LtPZbLpv4X6d2oK+/MO4y8fcCHyA/JFtg664TdeEYuyCS/xTG0Vs
1RcB1cE6Jl7RA92+Ejc7tFoXSFJCwJxACLWreseOYuflmJ6ILrVZXsYO5VMG0tCn
Axr3ID3cZgoO/AuhADsDiWZeCrwjIzn0wDsaJKSoPa7iQngKTrN8DNKnEit4ZDUA
NtcOEIspt/TZ/g1bKAirx123zXzHQCOyjPUXTOJ7+WeCquKKhlfa7yrcNaszd9QH
ZbtSGBLJe7jrWYeKOXTiwdXsJdMpoUM72qd8BdYlSO/hJAv3iP8YFAZOoHPDfaE0
olfy4meC1GosQPvDbnzF6TFLLxxKSct1f2ygeB7xYkZXRGLreKvJRfs+pP8FqGjx
BwfPXW/STZOwUAfb6on42T4QplrSXDq/N1r2JZE/v+5wGCCTUn5G8ZdFxMxiHkXS
RdJd6dT3A9+QRsAIB+NevvqNhxbXHcU+xSifBXOsz2fgPhqZZAVuAK75rB9FgMnf
iuq9TtR4qXVrqeL2o20+QjxF2z2m9yWrtD+XVqsE3azsQgjj8cMOFtEO7qB8ztzW
krfOOLHPqDTmfEesRIJXWG0IqVe2TcuOyGROIjKpY/VqvqQ5KyjxB0tXPwAD1ZL/
53J5pAi0ZTSaZDgiStqU9tNAgPgBJw4QDeVV+ePETgSy/dGvJ0kaOWJb8RGum/YI
BeyQB/dtPbbhEl5LR3MrscFYHOmH3V2M1jTS0mUAGH+nHl4cJ1Vnl4VuoFi0++za
Yq9EWPfHcYo/OCRKTMBX0DSsYAGfjXj9BQx+wxSEIlnzaxI2dQNsdaEJxJUwbaoz
uA+ccdXyeAX38QBxj/U+T0VALO0uGW+anE6vkr94j8niQpcAIForvekyK0E/viW3
Q50m8ESKYV77KqeIlvqK4EKoQ8fup46dbx2mhqIptQCXZrtUk81nZw6s94DAKBy0
dtzoScWWEkPFGvVfUW4br2yxZWzku89fEpxobVj/R2KJqn+ORUUzO6QZBu1W5En+
Kmny3CPlB8EuMMsgihZZ8HW52oR4XBkEcucmtmxBZvm63TseZZzhbuLNGydYr3FR
dT1hm67OqNCfsNMTBBUqOq1xvHEk+ZsknJdgzwIu/OJ7T4FC8Wy05KogaUXYn/eG
ATneFdKggwtNgtBmTtv7DIptwTaum2Q7+8aIynlRcbvHHHlcJP3Dg4DWx244PMZc
Ia0wSDBS94bO1vK8P/Ypzmx6FRQFaXzWqFmopjG1RVi4g79VtK0rjjWqGv0Jc+D6
7C4O7R6U4I8hvp0oaN0ccGf19NTvTKbXMHQg1NfIr61tv4znSoEx5iOPjx5O0ghR
wtpwhOT4ngBkjjSzCorSXR6XQdqqXxNkvPlzn6WppEEfcPUVCuDuJ1wgf7h7MdiB
RY40Ziqp4WaZKr9cRjosKfleMZduwR/C5uzNOGf1ggFMk1TGg0nqg0dGIhsA4Pla
D5J2LCMcbRHqdP8JcFEAogHUwiyGZdeogbx8MySlW0hFTjtAUgC4QXwojYnSWf1i
brwMUok7iz3LKJMDFF17aMU8lxVmjdq3gqioiLenGI3EJQeOZpgQuYd0h0r1AlEw
gKLuKlD3IppR+0PmxMjHYlNHv5gja+q5QmIYvQeNhqNnoNn6E1H8Qd7nanFuJfLS
vnP/NT/6GewFdVx2696Gr/8b/sWdNUpHazHdH0nnwNk1YWCIe3MvX+aljQkbzN+a
UKNUXqd1rPy7qV3qJJBR28ayFYezA0sXO8wGDpqOwDIJQfiIlBACn26+dLryaN+8
/2pp2yghRG4ZyW4MsKFKzw38WFUpzfEns4S9KZ3lTCkvGhL/5WShm5MtSERhH61s
+yWsBZEUB7nqGCzjpn3Jg1Nx4AH2zVUKObAp7B/olrPgBKdaNk8V3bKiGjgA5EwS
Wi2jWaIswLzKvbXCoCdudBzfUZBBQbZIxk0rhwNxfsL6c0e/24xiLwmNrsNfK/S+
U657s6wflyxyQ2E9oxAk1IC7wFLpUl16NdgOOZTsnXlDg4sok6EPzU651WDtuyK1
YLe67DHwhCJmrFNkJ6tqQd/A12zAJu3slLjQrsjJS3AMW8NOdkD1rKe9PSlcMVio
5ET9h1RbEH82TGTaagxaptY2B1FarwcEvX0HhaNAb4oHAtMfscDOQwTHK9yw5QHp
CzsOoS4eNxC5/MIsicP6KlgCE6ThJ6lxkmBS4DYa1e2BhUR4/WtbKN78H544uMsA
v8hkkRKcRRpLwokgc6iaUzG2Xv0w8IZNJ/aYJ11QmjwMfpIKCt3A4QJVQftSaAcF
hIhG+bFjQPQIdpveKX0cPhq4gjLZnEg24I1AG8TZK5xeSu42ZXXfHfB+Pu11GBLf
hQdGv0fallvQ8iaGnlrshEM41+ynI0tu+PD9Wxkyk9CtIav79L/46Zpn7rv5f4m9
WzYWYHefQaGj5u4oGzQ9Ghc9Cu4GATIiW72AGZbXpQl9TuEecyaghjBeJWpupJsW
d+utRg8ALddtx9cXNz7yYkFy2zZqj6pWKYNZfPNtenNCL9igyfmAOzxc1X6jBjdt
QmXHTM+TYHJPOzaJKKU9OdmbOivJbXC5XPMFq/V5yldBxFsNJ43+ulV4F0V3YxtU
NHkkbwTBxY1sYlIEWjVmoKb+VochW9NZNBr4R+zMPB9ThalS8cQr8VIWcpQNumdc
MB2sKo/7Ak4GLpVy7KcgAvNB5jzbhWRYbDcNOfQY5pYqEB4PkArzRu1PzKRc3+p3
zuad8jmoGQnizZt1Yskf1zE28XfOgS+M0pFF8TJGCt+EFgN1LfRV7HQuyd08Pd95
hgsKzGLAyGeT6fKLH+jTC+9PqrcpzQROJtE39xWApbXQ46yirAZqq/b/Cy7PvcXz
w+A/lmmdpYDf1Uwg8ak2oZrkwXy7d2cdhEetCDfoSIXbAks4LtuCiX4Jkp1qQpI/
c011x4ZZbR24p3PHL3fYDGI3cVg5Hhm5TJ/2ipHEX7jTOsQXNCuMNsqr4u5aMFFu
qvHE/VTClqesqDgW2SjjPTci7HjbaMTRERaK5RXnaukzXAdPSBbuUNc2Xwl2qKLR
I7kFvO8zsQgN+qjnqtlGt+YTPNkETEBe4I5+r/6ffAkIr0XE+Vh0JkhmVm5p5HbH
rpTU0sJNl81ypBGSfF5JQW3kKTt6rPsYS/gjOjdYlWEsISeuedQA3LXlFNJM/4Aa
gwvUtLPUEjguDb9FoajUqyC0kxL82zO+b2uvVzIuEmr2q8rYaiJRJWubHq1MdMeq
iR0z05bDt41oU/v8iDb9Gg==
`protect END_PROTECTED
