`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDAv6/pg8eNbUcQcDn7j7EZG/QKGHyFWN2L+OH59rGqsVSQg0L9rHoC2sXIxMvfN
tyWOJfs93aLkl4WCdpd3sBQKXHs2GTafnWhNuhvsKWV6JgYV72tNMLjZhjpJcFbs
Q4I1K0NAxdqdtsdr6WSbA08vNb+jwHzZ9tludWI3Xkl/RhVVcjOpzSOi9C91G7GC
ckosjc1jBncvUn3q6sGa8aqzgGVNv5ePwPLXIq9uzZSkFKhwM32q1xd4mAvpc66+
FYSzItTjAZ02Ny4IQYbW6ELny22eanfudCpakA/WQQjybJeyMRYIMx0a1WA/5tqC
OLbfeFycScr2zy9MncR0OdK15ocbeqv/dUEMIGDFtICg3eEbl85dTedOsBsAsib2
ptYDivgJ9Qxdmqv8egzKZHvZZO7Cu/rttIYtDGPk3o+/FSrWMmwJoOuNr1eumiR+
TtjxcthHccoOAw6mshTpUmW3wlxaMS8bYBSTRx9Awu7Gkne9a/4LAFDCfdZmOma5
MBlY7Xj4Mf5qkxUFQELwOsIDM4NK37Htp9/V6rYfpXa2ERrfBTPvmgrn0ULu3G0M
1utbFNxw7ZOi1PwNf24YzjPcviKXZwYRTrA/k+xjaVWowGNYoJkKOLfKXpRkVXE5
x/urEZgGCEk5XY3g8ya7I2WAdzk4WstUBkQsBcU0wsk2Gfhxl2Z1uFbThRKBiY3k
6V2pXOhCjBXCoBch9KKxsaZ7ZPRecj7Fi2pkx5MdQNY=
`protect END_PROTECTED
