`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFGqwe0IET0ol4f/jYI5rIp5o+6AM8EQPfYMPATgIBarQLjiKG/rEottBpSS74V/
K9089+j1oQCtME3PNRWX6DErvQZPMOT1X7DrprXOlRwGpBNEGIKsWJLExbvt4uV0
dLgeSH+Ek88Vf10s2bfR4KHPgZJS+h6gF2SdRAnPeOttG3OVppENe4ucbqeRH9jl
INIhM2jKTyFcKAdEq3CVCrYTn3YsAmRlWSv0FsG6pW/x4+sEMBQ2X9kVmfJbuiIo
SwihLCTkrdMAjtLkgk9+PEXl1Z2NuMoBUX61OAIzFBzvyZh5ZwRbDLDoc6TmTc39
dCn0qZU+lembBkywXcPc1JFzz8KfBq8GZCxPcFitb3TWJ3PKZ+uNhcLU5swqe6Pl
klSsgrjlmafd1X+iY7c8gzu+ngXlMUJguoBudnxpJf7/cpRD7k/EuepYX8xbehlN
km0NTGhAAGfBv6XJDjHEwvzPh2HTWt3v5qr6sxJhrQ0/AZgPKaHdbr0NDsakotf5
`protect END_PROTECTED
