`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yoaJR19ppdMn+sY9D8n6sTQWt+DKPyVlJhSOT3Vz98ftRaHIzh6X+4u1HXgDSWqe
T6bnDnQQZADYmLHgBFZBhqHqxnQ9QtwxrqUNEAFBmnCRA0MJovzA2HBvomfzo/a+
lHvdZqQNE/PIRWC7K0rvdu7bvbXBmGJJxe91eSFZivdMElPA1EpAfGfrXv/k/Kvo
ikSs4qsiuqL6dZjrZGYiAvMQQipEy4Xq4SSc7sjPfs0J23cIpAr/yM9YiD+SRu/l
U+zfYFYgnHrAvI0EqiX0zoA8If2VwXtIDeCzYfz64aA4u2/9to7M8V3sQxFIiqOT
yz+CJB5PtEz2eoQPuhiYseK5MoZni4ontuZ2VoCfEzrI7nspsSnCYduhqf3kiZPu
8rcguCRbQ+XYhvxZPlTHGOqc/dilysEcNiA1asVEXmGpfLytR4mVWiWAJ5HlBdXL
MXiNTLmC1OE77Hreu19iliek1fGG1EbGbJafjF3UBdZ/MyeGa17AfeynW2FtGHne
gkSEZjS98ThyWGUebS0v9eaMS75NOHdZ1/tZEU0BvIdW/LLyE2dk4wLSw180QOiD
B3m/nrkzcjQ37b5SP4tg2ALBX3sxeow9Csc5I3xg/yb/OwS1CMfSCrGdnbcTOqPF
mIimETm4cqLOhbOEChhU6k1X+YPoxO+6zSGueBT4TePKKQN4S/l+Z1CnTRcKD5ID
ATnEVSJl3Xyx5/tS6dbWJpgM6EOlfiBKDQ2RGyYwh5Y++46J8y0VJ2RrQ0u1iX+d
64ADyIY+vRnJ/sW8wiaZD64LPKDZLQEinPnZkWjRmg+7epEdNexUtZ1t+yZncn8i
0wEE5BxRWwTn6k0XPONg0AKnvH/KCPRMDv+v+/46329ktae5Hn2CbKBi6fFZdIx0
4OAavHgAfPMT7lvG3ptdX8QIM5MGWVYgm6I5cvbnWkbj9jhF3IxVxY49q37HDCo3
mwO56cqSsCDS9l8K3ycSnxW8Fw4ajrxcprEUFmYd0xmMv7xGesj2JkWNwl9iGuk3
gFDeWSRK49e8El2AHwNBbWMPqafIP4glFMHGbCU49eRiCCTSW+hDs9vtTh1IlAH+
wXc4pYssQX7d7AmmVe9MSicuaN9nDVtjAXIoiMjTqFS7ATOGZOZBRFidxvp/7/DU
lZdfrwiRJfVcfSdkly9lKHZ8+QyKQKD4BxfCt9imi8jCI5wSzQskcm6xGD28JZlb
hIYXGoSKVhm1OfnOhnB2bhMCugpjD2u8SNv3xSv1KEdGBp/G9E25LqBY81oezoMB
V3eywUtvCRvLMtXoAsKmFmK//455lJKTZ/58jl+2GBc/oHRyFlsqlv5pTcb8A2Y+
`protect END_PROTECTED
