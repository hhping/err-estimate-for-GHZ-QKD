`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdMhA5bXPBEnhq204BYTk9OEdakelwXiq+8CirkG8HJOGC12/nlgQfC+pYFotlRA
qIBJOJ4HUdHY59AT3jgPCyeo8ZxeBbkGS6tA3JZFksmfa+hIyus7PDEXVTX+4cBN
oR7uIPdwwre9khx+uf2uq+eaWgL6S03vXVvxVR1L0nHsipXYB4Q6y+TEQOlLCwOP
04f/J1S76VnJIk6Iedqeb9G7TGXJase2l0jByzP/1lsYhtjPQq12sA2WPfM9U4OQ
1psHuBPmQegNh+eRWrhmCnL80iP5lxBSCjcTUhWfYt+OuAckhWIRmBMpjFIzADfP
byFxufTkasFpUkeL1oTBjw3ZwvdXHLRua3EJNCE5FR/VZK9YHo7Ljy2zGqdyHta2
asEPIlOw1GJYjQ6yZtSJigrQzxEePONRA6evO/WSMbi2g2X8671ZM2en3DtcJAjO
netCSsJvazo3OpdcPASGsY/AlyK6WFScIXNrJw9BJKK4WD/TQBNQq/TvQLL1vrPe
uXF2iDxDHkZtJqqJw056Sc6CXlFKqBGMa3Hf90j5pb+8sOTcws83md9nLi2T5DlT
SPTzi2p5+lbZ7usifDzfYd37Xh0fswey+A3AaQlkNDobZIdgReEV3Pxh31s0J2oo
fd31QKBJAJYvNjuwek1HQgbsmwHn5bngctS03RWH6qjQq7HiBQwWehXz+38XODZo
7lnPmlYHr3ArHYDvtt/OKgBCKxbBG1Cx4j+g+JWDO5kuzcqZJXy87K1YElG37c28
gX7jJP4MpaurjMwgW4gfcwtf2oj1klx4PxUW53PPDC6GSYsZuv9xlfq1Eu4faAK/
2bBUYtpJ6pU8WDrX/BgvQPwbCcVHtRBVNWkyZX9OOUrJZ6zY8l5dpmPvmXSMODuw
Uyv4crsZTOrJ4kPB/hxvfWU+WX7B93ZZkp29GnINQjVKRZnSgPMIFhdN3ZvqxSs1
xz+34ciANQdZqzIvKmsgqmp2XS1okbUGKLiI87hkKfHtEkimJAFj9ZCFjOfu3UYO
WCf/+v+PR3hcBfpmKwTpQ5V/9XfDm9s36O83HwXJPxxbLRaYQrcaBHAub+5if4uQ
UdOiIfYeQrHYFEF6uVPrkf7tI70zsHZ4UbHmTvKb38Jhsi+gGZp8F51qHh4MK2F9
Ksu/f4Sb7cYPysCmbh8QKJCi95d3t0TZNYXr8IPgUWX8XmB7TtSiLcnXTtAPfTqx
5JdAxtFc82wvDmWJoW6jMR865+X6F1bGW6I+TQgCmb7gTgF7x8jx0M9q0czlOy9H
7vHTSS/81mlkZZZMgyzHTBwmBBntGeMAGpaGKkMuT/WtwWB0afiM4tCpGlIgjU2h
43xXM3LaX4Iv2i2+LFbgSEjSSvpbQrHNKn8oCyLVOYF6o9BoROdulJzfVOVDbtdh
PXfp/U07n3Ii3SYxtlaPn+MHHKiWeu6bQaNE7OFX9EjiDtItMseL+LfXS8ed3NBy
ufR9qlpPtxw1CdRWGx/mXg+sggPWG74te1mtJ0NpGkJJ+zyuW+JiGOTmAXMbLCUC
yu1UyNPlMzeTP7i/wQr7PB6dIi91wCD4PNUbdi/VvqJ/BPaT6QsxKYOnItXraz57
UG3o/6pnnfTzfENlSKtxEKe/sGQru3ZZBzpnUkEPph989uBhEKqKBiNWVdPo49XT
cd79JZJduYf6xS4LxMoruB//rxvGjw09zvW78jQniALzOc+WCuUE9//Wdywm95Ot
v7d95G70/gzpj6Ymt4/kmMU2nIh3V1ySWpj9wVF99yvy2Aq0jYpOIwiCcnCJ0CnE
/MNeIdwF5Q0eobEQo9uN8lyI2RVWrITl7Fv+r6WNmyHLG6g8zj9tAsDnx8vSaXEb
wB2rx0UdSqwMQVtVKxw94JC0GZDmmdNpiNeVHHOn88IoJD+ulq9Lc+j1Pp2i8G2A
fGRcsiztz1UU0g8NZNvMRKv9tyWcCyHWVq8sb1jLrOECNEFt6xrmDT6DOpOjkmIc
HReXzX9GxkYxDWBAZkwBEbDGrbMVfErGHRACuz30g4jhDYWTdTyNwGEsyHnWetE1
FTTsI/eclj3sAbwGl7WsZAZe2bHZm54ZNGWNMhRqTxvFK05gwoDvkrizml9RMebd
xsQMpifyC0UR8ohAfuuT8jS21HXfr+MZm5VEf0Xy1RSzwslTqO6u5yvgZt5/vZLt
1+ncKFHgZsEjMme6z8tD13yZsvc8BFukKvI3AK/H3RqQ8j+XExeOw4yYwBTry0sa
G7PjuI9FoqijjEDxDl6kQmDv7oyBK12OUCkpQh23PbeHEr8VXLje67dU0YSirRFn
KRXq8AT+SwKz0JWRIVTInGvajzqFCdfEXnQ30RDDBs+DQW67FGuQepnkIUErLbIE
14RQ5CaaELflQykYLIhNsO+1VgzmscUiRqgdKpjsmPCwRsXmm8k7yehk/WoUm5Gq
QGO1rTquLmaUL2PSCxnGD/AWhsg0v7szhWpvch8Ufj+2WrNqAXwGE2oUdpomPWMM
LNEL/u2uhOy0SAVvexJReJMXTjAp4pAsgf1hhtaLwO3LAHxRYNWCtsCiPYnm7f7H
`protect END_PROTECTED
