`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIbYi16ZPZi43NGDNCxs0NDSSGh5ef++3pvxen8BVn/j/p8HSqko/Qn3I7B2T7IP
Dthy4lPtA2xz4xjshPyV1JmZ9DZ85oYX7JBYWCF2tCQvgjTfsX9oiHgfAzNblNmO
YMoOD4sedGF60UA9160Pn3dAI4lZXNf3yO3U+XGnN9CGzqZ7blSdgYpBJy3tFKAv
qfo/KyT0OJC5YyLHNkaDYUC+RwROE5L+paWwvjzJnNJxWwmaeKygcEFpYv/OMrkx
iBLO+0v4+GwdBj366nfhcihA07flslTLIVzm8lYShLsA1re2FdS/UrC0d/KHtciI
wLOMgnOcsMOZ5kLarN6EzgtMpnzEOKlAVXMIYMFaqZFDheEvHKAEsduyYX4kOLQs
hdQvYep9yPSVCc4T/Y9mfeb0H96LRRRH1YYsqP3c2PawRCJG0AD+bD59Tnn096zj
G9R9xLhaNir/BzbbcCXkejFKeHXT/chk6I4kEWawmYY+c3N2Bkn09gGZVvaQN6Oh
tVsqXfKXX24SxJylRAeHR8vXsHMhpV+vFVHyYCwQ78X98d97mx8DoDor2UyF15RV
RhUz5HbqJdBHsArHwIjb+qsmtTL/C4Q/8CAAEurQeIRG46e/yv9QrF9egXLZBZRh
nX+OaaDgYJUKZ2PCeqTYkpR8i7A0lFWU8LEr4PrX1I+nsI20akMQLu6T7dQS7qiE
57CVsV0axrJKU19tdDgsWNDYmVl1aTqPC5TKug+QrgzkWUFKsrUYR+DnMSDrCpxH
qKDA1TGahBel8hykCpaxBtDNaSfMB6gvaC1XdxGVXro1ql2Of5mrDtBjPQ9DfF+F
QDO0JFuGZEpWoADMgZlubLcS02sJtrJ5B0JERxN8bqNCvniI9E+JsPutAdK73fGD
k1lqnQZpCErzRLJsxZekQPG8kiyi8An0QnTAZ8M8HnLYDpGhKC8zyqH7Fpr7ohbm
FxrIf9hSYqLmpSvr5v9jChvED9fORcl3ao77+2o7Yv5+YRrvZtFmJxBGb1l4BP+/
PA5AxoyBqzuSM/l5c6krExlNJuXZudsFqPTFmekvTIJJbCDm2ofpvSNnbcZ6FkZ2
mk/K7R/F2semokhZ6mEB9Dt3AcKOXgCKtcENhp8ibNRL7LeIXIPYvbX+5Cg/hE2u
N8J/eqbfIFd+NVit8YASmEVi1nblsgpF/BKlLCMFiLM1cdvheFqUaQn5R8Eg5/CX
+MkFFk5+rABK5yN4UVWDvZC4D0rCBlET0FVV8V836O8apiACMdu2EkrNeFcBCOrG
5XEnKezDVGbdrfAzmYymic+WPd7U71/RCZjem3jwwTFlz40fdBSUFJtWPSPSNEIR
ddp1eQ0WFmODK/Xw6MOLhS8yzjhu5G2HTSGs8HjQWL/YXql3bOTxh5yk0mKwN9/r
q15Z/FHFyR8S+fiPQaZNzmV73W4jrsPWKqh5aJ60qPbpNkeoQjRFn4wKnMFde8u9
LqMFGApgYtxaifpAPcq5NRoFKSXA72dqlW9/fIHoG8lD6/COqMycMkDC8CNQA6GQ
yuM033a9TCGT+hK+4Gt6d2qV10W15aIvskedQW21kpbMaes6O21jchuoR5u/sHwj
dKwsPm3/dd8GlN41PAzPsYOuIibZ/XYZPEAXrdZSJTGJP2tGd7IqBEFVkDcaqjoF
PMrACD3hS89KX8hrjrFr/ZNzsq2rSj8asB/Dois99QAsweCRgvZG+3bLhLLdK2Jv
/DYh419htENDH2clWZwvZbAvzaa54VzojG0J4DGwEEApSPij157prV4b3aNX3BI5
3D2ygAUj6fnLHyJ0SrSBU32W4zSzcVVluK3AHxai0uUJXfGNNXkw+U7fwECqldrZ
NZbzRIJgDTUa3ixWMprS3bSzdThAhPOA5wlk4fKpXxxEhx0XMmqCuzgowGVP0XAK
tUAw7JQJ7YuEbZ/gIF9UAOMVEt85zKKR9Q18bzkb+2xYbPEjFiEBkSt2EemDu7vw
e/PNBlkkB947dfgezj8Rnkui+9BZoakfL6SKY0vONfBiMGV61gAO5hZ/PbkM2WRb
nCIC47ytK55vySCthDirkzrF5Nf2GcsVbtSPjtndVpgbqK4o08dDH+Y116lN+om1
hIUQAG39M74P75ezIfBbcFSkD/D4D3ypHFw6QOjBQkeZ8XorWpficI02aLicO3dN
Te/W/RVoCAcc/b641r93KXHMYhPIBLKIhpetQGDntsbIExX1An1CtHWsH+tqj8Z0
kmjpPk/l0YXkF43iwZeUIPXkxxvwJjY2Omx08g4JPgMXt7kekS+TpjFd+DmSLqn1
QDxJpNJxlgC4Ba51exP01JRO93OndRgARAhrc9fkVAaIzkKbLTzBuKvFaqus644c
uUhEwgoX9wV1+YRZT5ivU1EIzcXylzPEiGSUV+BhT05Kpb6IsMVv/qRTQ5HeNU/A
Ug0GdfojCfPp7q4IQ6FMdJ53sS8uzkK2iRf1jsQcqhSi4gbtJXIgTjFNCYg3HfE7
sEkuPm9c3qpg8eyylbHWpWJA99CKNaBQQNJSDu2EPoIuw5YxxdCfRRclVzIKYezk
Y9DGZ3HJCgW1oQCvYIdaYg==
`protect END_PROTECTED
