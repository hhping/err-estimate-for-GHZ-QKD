`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j4YnJBujd1QRCDZ54Es4c9JLQGRUlF/CK1vxvvQvjeeESveH6baYXvw7Owm4JHY0
xRVV+jU7SfLEMUMq9B90j3Z/osrM+TWW07WizrxWKxHaYeHCc5B16AYxilA95/Oh
kzH7WE2g63wXDKO7unAPov0j2YqGWGW8bOXgL/riW+2oG7+ECsQT77YagZSwrj1S
SinDZGBlNo1nOX/+yLlq0tORw152EtqbhGWzWk1a8gPUDv84h0Y2ZAELsZQktkLd
cMniurGCqUoYAQ3zIKMRRtxOaC3EpuAJWbmHvrideZLBB8G7IJTtal0e1BTlLu/K
9njYlsw2ac4oPK+ytkpZrjGokhtT3MMoOfCuLalTmO27qPxhLKN/An/8dfKPwj7e
7BigzBiO1IJVvNZOKSRDfbc+mH8qEjXuFlxAMmp36WHTUVKUdIFrKVnYhvcz076Z
bAJEzDgY+awCakWWVwoFx4n2hmXNkYjvri0BEzuIi5+f4hDmHiiuDW43RsOt17DX
TUheHeCO0rbGJJQhxIpz7eXN34jnyri/SA83IU38r2eYeUO94YDeEC/XcqSK2dPQ
HfKXcwOPLjr3Tbxxg5YeMbC7oCsbBEO7uZKUU3NDgixb9BdK2ASqoZhZbH11+XLF
PrjcrTtUlsdDlJvtUU9lbYpUfDnyruMQc2XiPyDbwaktI6kEgJhpjEls+ABeXaHi
ysUB9NrWyhqfJn3Z5ZXQiZd9XVXKTEKyF5l+1tvpBOfw2zDSXAAeFiR4dmKlysrI
JOL9O40DgXRug7ynZoBI86uwtL0GNBb1FgX+RrsPDf4nBfELbUcHkCJWxpgxAvYj
ynlS7CEV4O8c3ginTjhOqZi7IGhixGgTZfChkvmr7fBumQYA0Iu1lfCGImGki8El
ruxw55PWivFkdbl2iddDT8S0Ej3UW/NqpqjVjobD8BSS652GTHM67lyVTclhM9ek
s68/fQt7lGBvv2QDxMQKi+8CsGIF2n/phFj2/tdokERhpGMs04pUv3VA97TQU7V6
vDWBc/U18EzpNBGLXf8rwo58tQtMEb9rDmbDBOTxLg42kvyYcCko1mx6HTRpYpcQ
3b0st4d6nwH0EEq6CsZEkFnDyGTL8tWxFEC1gGijVo7JVW/4pMhSnTkepCzBB601
VO5sw4/lDsDTdGMakd1tHce08AtzgWTpu68tv3uZZI+GxU3dmkbwVuebyRHLcXYB
90kZCZU8bQPG+8+kmV4Sfli1sNS/HPIIkYNzJxrbmJx1LT5E83tWY+VeSZTpBu/L
RxpA62K+XuIFYqI51p1ueEygDVJJ2zBkgsw6fFj4OoSgNwCGzwa3/WNCXXyPEbeX
IfMRLABQbT7ZrNMCTC/ql/up5KCFxWtYhh6uzD0nej7mf2wZ9uAZsmYtwuxkz/YV
WIt1oI4ZL4xpeFW8qUxXL2Qnv/BnFmGFIYwJqq9IZm21+KjzumiGak2F+uV9fLSY
m4DLc1OqTvvGWAoxc+CzPNEu9G/v0ytp7f18ySU2fbAjwGib9H87rauOp9UFwy2G
ShI6XQ/A8NrCouLqt+U466en/qk6lx1iVOeq1HT95yHRWx0mWc5g3UEQkMZKpaYL
ZS3wCMhaTYrruoQ9fI1NGALKbOJ9FRa2P+ZDa7fFrMtDrGtavJg60yExL+/6TBtE
pzdZ/XeAuqYULdDKLYYCp4UX8OVy8y1CKUIRupQrU2pAueuRKqNyzEVln/Unao25
DXo8c85Vk5apurBLXXsgmGPWtR+gTmQnMWAu+IBhyfIGU/zScIAFHrt3eq6MKDRE
XXyjtSLiGQCJ5LQuW2TY2P9XkArk/vuQKsxBkD597K46Id4P0Vv6MMCjsPD06iEW
QxWgkdOw4z6C2ApKvHirN+DSRhmWkJ7An/NVyBc+87XMVbf/quzgZVWt1nYd7IhO
UQuxCWdd0pxLHwRgWFcvXuAJdto5fvDLJYoef79dL+Mv97W5I/NQKwQyuXGiomLe
6jFdDRURQij+C8mr6HMf33yqqpOcoBUjE0HPXnpYxioth4T6NJsCi6tbdfDKbQ8f
YyHA8PCK2QOFDuSaUGTeGpoRe2SvGIgmGKjeedikinCAeSYyi2ObZ8vtRr0RL6ii
03mHUuODPohV4rEI+U3or9VZr3Z1lnpdZsfx5DsE1qro6vAEQySdYzs3ksd8gyy3
cLDQXMHDpEhHkW4gFJE3DBSQJhLjbMd5pPxCu69TaXqyRIWo/3R9dCvglszPkVBZ
5OtohRQbfyixn/mfP2e8emuy+56aPqB6aZYYksHWb1GhO3jPmoj11nvBZhJJfLql
AkvGoaa/Sz/MJUkTie2B2vdig+pZt2pNUkAet7w+dczN26tgfz0uZU3flmwx4X+Z
oIHfKKahHfKHg494dUnXknEJ9L1GHq90+U/2dj7aQk/lW1BUz0VON0IXOGN95Yyf
RXa4COL/XYkEr8542wjAWqjteAi9bfGhFcJV5MC5Dgt5KcKk96UCbcONmy8qaSc0
VTZG8UNJ64oXZ3lkgrdUjCdmyZNuMj2LPLOVKW1EPREJzXqvhxYnHSM+BpFyKyy/
ycp6PTGbX8EvO37dTRG9i0SUg/CIAdBU4Mn9bkFaV+9H/tw1VOCcwy4CVD2VbzgE
t31kBKGkT762Ex1UEMJ8UfEp+vqkelum1b+PUmvwitIOjk5luq4OCdTUvwFwAH6t
VRgvseoLBj4lcyexVR15TRyX+7fp93FylYGDpFEPZvvVRix0C4ysNy0f+R+plzJT
jDA5eGW9gWl67keivtQHtQYQjsgg8HlcysFLqwdUgKTnpr0Odkz/txCcfFaPJg/V
ukjeqmI8tnh3U8NjqtFntQbwTh2OZqnmz+8i8uRY3bVPJkotiwpA450dnhZThjgJ
vlJg9Tf/r7bj+MqxL0Rbk9LqzU6H/CVXyTrvEMN24nk+cGGn8ZwjWqMobOLDtaMf
LFq5vh6Ott1TstREUb69eF5R/Prl7nzFgNf7jPh/tBX+yq0JkuLEb2a8NPzF9z7l
hsss8u9c/G14G+Bdvqs07D7FfZ+URh/qN7rGEJ3UEQoIN2kPIxY8/gAKPnZmluvK
P7OAeCzX3m2B8g6jIEB5NgttkUK1d3yFTxNNTqQoEACyYxsxMPrtPPePTeT1vFlL
`protect END_PROTECTED
