`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qr+7i6cmvqri7Z2GQACTAe2K9jgSIUpN2Cy0BwKiyjXjgFADl2Ew6wg1HkiMwBag
VFY3rvEZYWF7AhEvs3L7uFHl3eqJDEectJL584JQSVUvXFKeaEvJ8B0Aqb6bZcfW
n2Qa7Tiz59eCkQzdqVRwnLcaSKqbikQIhz3Mw7n5CN/Bvw+2HSZNJD04ngZWQ9Hn
VVb1rQbAYwCtQzOpyXfWrvUt3jklhpiWQe60M31nezqbye7LUK+zlk6g/I9kJlHv
c6wsfN68+srZyX0XigjUs6uap/t9XPjw2j1fQatfSA8DLZtbj0lpmedgqV7xn7G5
ZNodfrx/LXiSdm+MJFlZ6hRPX+ey7GtvvXhgXxNRXZ9qOWgLRE0P1Amg9aSzK6w9
G/4KclCbjE2bW4aFE1OV0gtbnAp6nqqn8z9owSqiv/UlhUtEtnXnD8IoneEnQqMa
dMpk0tfw6y8p1wWcaPCIDQrHSfzchsJ5BA5ScMfxYGIoIavdCpgzLHNfsT+E2Qzk
n6erxRGhsJx8PnyhmuoEeaE5+tFii7vHRNt6ZccoySqkMMhkCYx5SN1W3k8spnx7
c9KsRHPiOv7NZ+ag0hH6ABeh1B9eJwzYWU4RLsnQwCM0WHXXPl+Rh+PVD3TzYYfU
3qupBfGtrncyYZTfl4hnTS4isPrf2YKxHOQHTmwmv8z4kd7sSXPbQlITHZ0OcpiK
Ynp9HJzIE1xpoTNAcG72KRUmhbO7FVGu6JRnQfjZ1dpWEjAoOHDPS9MlIvHPIG7u
jhh9dnPR2n6snuFV+PtZGw+n4RblxNY8tBaPIEnJeNC1F7bQ7L7IG3KCStMvOamu
83RyOmjIvzcmxgdQb3WRpVylPxOKATsubeJyKz6GU8cBcFi83aszeCKi/nvvn4wg
aan1ym0oUnKkvsoCKajoKgJ3PAT0n1Kv/VCR+6wpCUrf4Odx5HQkPB5iHn2OjmET
7sVGqwWMdLn50L6i7KRfwGUgr5vI9pGMJeci9QDFnLLYrU1wGIJI08Gh5bUtYgdy
MFxshHF1EwsEEaFlpjaKp3A9sHaWKgWMYSmk8CiQc0gfG11o6d2OXIc6kV2dN1xU
Zw0OlkqzkqIJSxhsHSm+/iELBo1AxxbsmSbZA8AEsvDaUv/NgP8bEuIoPjQJ9kX2
08d3VcXst/xnZFkSWJcs+ATlsAD207rAdjRWo9HOb6CHurXlz29QNOwFUsv98u5O
Laa9I93rIPXdQse9FeDc7uuxUjeRhMAqJVmZYbTaSRhZ2fQAdXYyz8BkyYXd2NQK
Pcq31tZ/y1pd9PhaYFFGfm+zyIIrDfiUq25pvjrJqhlc3jXSG70bGsVIoZBsgjlq
EEJw/DYl+6tv9ECyE/x6d+wgZDEk8DaUdrrqn7hmlnnLy2mI7UlIJgUaW6X6J+cB
eftV46Hi3LfX9S+XLvzo82j4YzeNCNmfGETxQgjvw3hEOrohz9GB7ZvnKOAg7IQU
iSm9nYNWzemZpIlVCsqpdxQrpmUDo530tmY/LwO2f4RNWvT+7KVp0M3J9P4g+ZN8
fUIRrD7GUV3N0EQgn/bdAAYPVXZxHjo3zpYqQB9XOYoRs4W212a91VUX9CXZTqNL
bfD/cxNbKsyEsVHMOnhRpg+EGI83gYtsdMCBvBNQH+R01qOOZUQt9Zv416RuZF2I
x/0ieL36tCRhpoAyh0qkXQMFLnighMtkQQDTWLAQcUHj2LGBITZMrN1eXgHyIRt7
kv1uE+43iSD2YKhZJ3kXjGWdzU998uUFKuYm8v0RuPjlhDPNxO9nMGTNBXSGYHoP
eyL2t82NCQFSrEHq5fMgqICsiPEtzQkC34y/8WI/E+HKG4mutzDIxs4AiJLDgna8
2xrJH4MLAOXkFOZpHa+o7NeVXq3ymHF0xChS0NV22XUUB533IeKUQlEk2cruyEJe
hmeMhIr3BH7349CGmDjHkflaYuYPgf8qNTwaI+enEpyaQZSQs8Zh+PeQ57Yc3n3M
ooYrg98wtpJUNX2kdmSNevZTzCDXMew/XH4UA2rJU+Tl81eHS9ftXrwkN6hNQyIj
C2L8Hb5475cXD/2R4s0pYHu7V0+Nu5zZ7SLkxb/bg34A8QdCq1k4w+aT6mfC+M1j
n07yjrgWJYT1jmrlokF88dtDHiFc45Rf0wuTB4agwEMV31ulZ7SQoVJc9g01OKIe
b4oJHQNAsvpYLnS3uZVing==
`protect END_PROTECTED
