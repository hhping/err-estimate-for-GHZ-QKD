`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7qYfDXcnGfLEbhVQhYpbnQTnrqSmhcfFn6va6NWcadl5yQ0TvfaP3PlgqlzIpZq
gc6D8fsAUxxDvP+Z1eh8YwzT+g2/sC8u03Xt7bgDtquYlK6ItyU8QwJr1GWXIKPT
nuBlc+xhvIoYulD/qwr1avamOxKSMFGzn72K+qPEaq7lXO8L1Y4ubLN1LRm2ew21
4vQXBRZ0McUX1m3IhGRpAW4WxszAGSLE8w/7tVBFcDlUksHWbzElzeQjjssKJqdx
3ENiXvYvGp2FpKv99aDH0EjtU4fg0niAcjBTRQ2RhYAyOXiVY9I0YobqHl0HbIHo
9CAcdaiZ+pEJ1Q4iE60l+BSKn/yRZZ2S3UyXz2ILUz7Zro9P2CUDJlRO/5uBQXkx
5MCjmOJr412dA4cczyX97CpR96PMj8FQ5+eXMmIwwULaVjG+xDOw4UQbL9HHNFSa
oOKPkcp+LouI4nq0G82H13mlAubTMJxa2WyKjvfBnWAApb5ltJnkBSy9MTsRAsbT
XdqP80Hle2VowHm+KutyqmPeXX1Nbk7Q7rdwB3buoEvo5xFjBXEAXSgLvhOq3qdu
yOvbXgDu1/fQPr7ihLctOtYXVUDLF1X8VVpVSfwlsy4DZWNNBfNFjOrc6wx1q281
2zZaKITiADpJna9q5ybskW8hHQYd80RhG4rb8lFEA/u/rFrxPKhx4RD/Pju+QgaA
LiDuN5BGmKRsAfIT2pXX9NQjm3GInKQMJsPwqkZliW0FK8zFVaY8xaKmPtjwqeDI
35P+tWHIHrMpYXp1l3/smbvR5fXiQKGZjX5hi25deuMZCzCQnCjTLGxBZ+7U1FYe
NCN1Wmeg6KRzRkk5ag+9p5Vl0+Y/wU4+7gafiVVXK8bAQaSumDV3KiChTYL7k1Yc
GrkW3nJASXMRkLHsRulXAgR3ldTBq3VPi0U2YDg2vb/bg8RMxnp2o1ltmHP1pIGw
/W06DLxqIKgbd6EsOCdEUcTItTbbuxnwo5W7vlXY3giNHPQsM+nW4yQZtGI6Xqxj
lStXn+AeE9WbyP9V3M66xrZHtvzPAEG3Id20sccbI2oY1bzdnCvM0AfkQ/FmRbnG
4euj2ABxGRK1jVsI9gf4LfF5B2uJP+93ubxuR6Xe9FIGs+mV+dWnQym1CSQ1x9rr
`protect END_PROTECTED
