`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7LszpfW/vPgTbq3cq/qr+VRBXTYP5HKaPArx8WIq3KAtwZjPW0lpAjzy2qF1HJx/
9ORrGYpAcCZK4dUh1UYwZQsW+Idhx/hlYPqLjjePnk3ZislBpg5Z7zFKPstMTmxf
A0qeODA1m2KEY1b9qNVYKJS0XDsJlhuFPTFXkW3N8Aos+GSdhVafhzz53kWFspPX
nWhcMMgO30+LW2R45c0Rj2a6TCbJnblkVeScyJ/PBD/ipMgdVpGRtau3+Ck+/vbr
kLyB9qtzxLtTHY9QtjdLAOJuWpkXlRzmwpzB7SxN+qBzLVxk5VMVSPCIGW663leZ
/iWYLQdOhdKf4NQytaFmEn4tl0V4K7NgyPsO6EfZB1NfZSzfVZxtv17IxN6UyFei
g13Y6pHUkLfE2SY1D6XFlRfPrpt/2T8ZTuZqibIJCeahP5j58PpdTuDJt350mFOI
5AVm9SK6oB+jKtcsB5iVh9FBEftPYhgqrgHI8lFq5kl+00oatWOdl/lc59qFlae+
w+btmzDOE1fcG+iTFtQYt0/60aQpLXhkpv/thlYC8+MxUnoD0PibmSfWzrcSat89
OmoIFmIb33b6U7j2fMEe85rZ7sPzH6WBTTiOafA0UWY=
`protect END_PROTECTED
