`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoWs+BVrSZYIPKBLbAWWB16kD5Xkoi4ecmtQN3mtMCq9nZv18YePdhaNVAO6eHx7
GRNlX1y8GMHWBQikIbm9p2DpAyS0WqJv7/J3Z156+rxj1txY7v80I/LoDY3Rj+sX
qsNVJ1OLToHzpx4q06yxQauKL0vkKPg3P9et4PeV0kF0bLrFiqEo6VDFIgYyFbaX
e+iIYD2TdIBfx+h1lCUr+LeOduHlAs2KcublK0XoIpxw4LlChCcnLh/A8tt8A8Oi
o6p9/hrHN9mk7nYpWIa646Y6E6eScB48FbdRIBxoSal+bQd1SGxMXcFIgxFTn0HY
SLJtxg3+AYmNF0JGCeOvzk53zl9yvTKTO7963X3CdMFRWhP7TxamEEAOGDO9EgB0
SEFRIiNCVsNnbsD9Yei8UG6bbXH6IWrT0dtJLuMvKCC+l22ll09tUKZD5Cp9/Iml
LcpRrgZMAvxvCXU1ONIsUVjB0Q/jiL7GlC8uOmOG+9+H3bRl/02EDb8ze7CytIlF
2R8h3HMiQtkEqrOmB7htdT1OHU+ULs/fJSqYaggW9tt0DmutihpyNeJEkN2a0/u4
et0mY5Ar7iwGKhPgMs6k159FQzzZfbZwiGBzrtuqHYyRm3gg+62GeyRjVLIEy9sC
Hg/8hUqlm36ICfMnqZtcMDwece43fJuNAVc+uTnvzGtc02mKuFb1IdaXqXLXDV2T
Q3R4CmaeljE08D8M6eevy/FmMex6oj+PUcferUETz3TuAmqeasWleFkReXv18ZaB
VWaiDb+ckhndcBiA1433ujxscDn98qpavV1iJkcUkV4df77JvUv+49bURQmLO74E
4FkUyDMgX9fqJ2aOGY3tf3Qd39e0/L8smh3nfAxz1kGaVgJ7Ef3Mic+zix4st1Eb
SdsKag6jd+1Q3jZQKlJS356qy+5dNGYXXtTkhN1x1+6GX6ZcFOk3YYjAE5MEfZBa
nHRtN61CX0CSoUNWDCCsdPB7OCc+5EZby/YQcg8htIU=
`protect END_PROTECTED
