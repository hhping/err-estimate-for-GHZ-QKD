`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2vh2pSMBrbvpIioTbM3PE89F4w/M7xjxKG099Prv4t774+aFJ4igcMiIIUD4sS5
XZXC9Ml2WH0VPLH0dap5ZBj5kRhbLKNlz/MXnoYr4Ai38YuChIXw4O+UVbYrNgqL
b6kxDlRgldCzeZ9d8PKl/XMOSnGWFKJCvp2/qz1MeqD9+YCXmS55dzbIVVJNM3Wf
13Q+40/io9pN4t/NbCNp5ytjfj0dA3MfDEGHiJSxvJdqE+/FhNoD9/fMhVXURge4
PPwk0gVyk0jMRK6elY3jmcqy9PKrsKABUS7ViqjDHzInR4UV/qYJODGPsCD+a4Bk
LEMnRPCYK5SsqR1JMzmWfHHW0T7WuMe2MdYH9FEYpLLeT/N9Z4PcWdvwCe17XE42
DNdx2IyYHF1V9R6OeDb+BXYHN1siBZ7ZB31qYmiHNSILgFmUG5VeEuElUrG/6B4v
kcdmJHw4QfmDBH321mgZaKp2t3vR+wl85SnJVqijskfsCjdvwrPOYUE5gbsRec16
ThofdHNBOFBnuov/7Du654HgPKfZoyKeoTy/nZpWUGyPD23LVoIJjF0MthrJAgWB
KZOwBGW/yHFOgv9+6ZXGywOjmOh2/ThJbaW5Z+I2QdtakM/W3AxJukmzfgJfSp2i
sy/VeQ+HZU7ACzm414ExNeDsUMF8bbhfNBFuAbSEkdLGZr1TxFRUYPx6a3g3DfW9
ORhaK3B9rjZdXz1GcbaEpQ==
`protect END_PROTECTED
