`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kQekLFbHJdxcBc0cvlWAyf2N5Rg313nEwTzPSKT3lRGevLq3bl7/SpOMrhoSr1bG
j7xwjr5KxrqPNjBPPdkcJg5hEnNABPzGM32ltRARfUFlWZ6NuByI2cCZnvLGQm4a
xQqqqw8ZI3hq7o5BW2c5tNQxxW55qJcgAdXvsJzADXqy6VewclCAOaw4is9xWGpV
IJHmVEh2bue1Mlqkjgxg/mFeYJKduQGQva1+Q49zbcn3DDkqPvGAWJxA6Dn30+7R
kDy0kaB1rET+w+a93G0BzZm6D6TaDbqutd6uXV0cTzoYOrmBBhx6241OHNKHdGio
3peF2nBuxvYxEJj01IdIX005SlYbstUQT0R8oozf4dc1pNDvNHyFg6CVkDPxjPl1
xiC/QXucwgaHjWcHqBYmoZPosswJj2osmbfMjW1TpsqmRGmZyy74Tmi8Yqm1WKGg
vCsbYmtT9oP8C6ry7KgqINs9jZrKcQEBd6Fwx5pvLWXG4kec7ES+ZVgJhRM+KvoP
`protect END_PROTECTED
