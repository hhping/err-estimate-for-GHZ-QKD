`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kosLGrXgU4S/jLHgi1tbR5LuluKz9ZKvTYExbF4vDM4GGkO5hHgoqqbcLsq8NYbA
bGcyKD53ELFsFK7REC0N9j/sdB+IIvAf1HGATiIEf1H6ZWawJbf3xtKsaCb6WcHg
feuPmQWkjyj5HiZcCQ1Y0oR7oIIv+jtVPnwiCATeAp3VqIAHeySX2rqMouB0WgJe
8GGJqmnScHT6697qh8zJxpNRtKdxDnvRN5CtSNab35TDetcRzb55A6prVNrzkhAU
8J2dMtLqJN5U2O6IKP8wT0XkmtxGKUrkAvmqhLPJ10C+kBTkO4vFPfmrXM5jAl6e
2qxJRDt8eHQ99cvy/TdcGHewvpcMTskFxJxaZTEHD7myT6vnam3tD/b4WQbjqwgJ
SoV/BLGFXAX89tW8NFlvWkJNFtZET9RKygFhByD2gotgvd5iva43njJ0e73UciD6
J9AyPgneTl2lpwAzf+FNNQ==
`protect END_PROTECTED
