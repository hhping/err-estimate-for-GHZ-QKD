`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DcLie5c93cJ6yvUAR4dDBPjNzJsZvM/e69/1hZ3zshzxx9XvlvMHHxoWftJ/4zx/
c53fw4yb7/4DDRVQLV8UbNLElGvUknIlcNtkgve16de5LgkzriMOyCYp2AGVtVEH
NMwshNFqFBEaPwMRbD/f1z6syrw9bsAu44KGt0iXhOOw3soqeS+uLdp/97sSFNk0
YqOTsq1aRHZNAF9iBOlj0IC453b/zvlSquRfYPHWzXxMkc75WhaRuhrSWBlkjLQc
io/Rv8w3z++bpUd5OsUMjgE7oEQyELJ6168IUIbNmQVdO3uOC1joCSCA0YdVao+V
4aDjrPmEZjMdRs3qPXMi2aYaIb+MIYHLooWPKzF3qWSr0kXUXSzDqT5m3yHDsjq1
dLUc+wZXdLXEZ1rXPd+B8Moe25UNH6+hsPeDwRqGnlCK5v53M6CtfEimEr2iPJO5
rYmDMsL+9/hLPq9fs64qXedkwIJQU86To8QmeiVehFemAzBx9inK2SZg+loKLkkI
NzMxep7DHAAH1GGBxxc83dg07VZmtV5Jq1bWUyzVXBDfTE7gf4XOS2b38FS2ssHN
WKPgordr1fyQ9WpVd0gbmGoVN817RVy5vJjQZsAElA8Gi0YFzri5Lz4dGE6e+qWQ
`protect END_PROTECTED
