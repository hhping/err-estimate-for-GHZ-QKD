`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNRnq50nz7+qoNJ6Yc9dyHWZzrrY/X+UU+QaTWB8U0NPZZjFZOrk9hDshaxaSwzA
EQHqe+lw2oYDM+hFH2++J6uxD2UCUqFIOnK6JLK3/RMoJHTg6HWVE+Kpazq7ZI/I
iFTP4eDp0bHe9GPid/ViZiFKXuykx0R7Jw25dLA8wlk8b1ISB/ojk6vjUF7Mvudd
+WuK8KWrbdXwEHK7nh3weRNheS+sLhgsz52LJnJBQqHHfMCSYzyRYK4Xej4vn8t7
0s+eNtki6TPanxOY9tFtNlhBYBr+bj5k3Ooag9I+/dPjAm8jlhO6kiWyTZwfdid0
ABAKilFw3G6wOuPs5G2pdJeEw/SvZvSDvdgYOA0Z7V3Zut04WYi0plTsVaM28Jq7
2e8uWOxz+/40cwl7AhvLAkjhjCXXHuz9Ah/kduI4geA4rNtkdRgbMfvNsTWPKvA5
VezxnKQ6B6YFoN27vtBYM32FOCgttSXovuc4gPJvcuacNOwAPXFDzLyxYi85ygYN
A3+t9IIEBx20JrVLTX83iUb8Jb6J62eiu/Q9SBAtu/WQ41201bPsP2TEeiyDezD7
8AXFBuSqgvb0cHhB+pcKPokAzF2CLJZ8fl0Rce1Mp1tXeC/v/sCH4OipldZVUlJv
ILGy+YK7ry1/ZnwUPWN9HQHkaQT4uCB2Ah13TFse3Ai0HW0I8nJdzzfUyNKOG+gj
ujfc0A1zaOE2pJJmpF23OcH5/T58kkBMDepE4Fy/hdo=
`protect END_PROTECTED
