`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
emMYddatatQU0jox5IVbxDEMZyLb/qJWogMPAynW9okP1l2eSAAAk7F592L0Zz8K
/IB1r9FclgCSGx092cHnMa7R+k4wKzJD67n6Gd8he0rRxaYk7nQtGjy9uotJ/mgR
kCU4TWEf7cIM9QxTy7aY9UDZKMa7LrfaGiJ4gIivLEKy+wcBaPQc9HGQMHVh3tEN
D4vmqQjCd2o2l3/jFrCHL5blCMFbKd6QTetmQhRgZ1ZGevTHWeam6RRKW2Vz+ETh
h7zBzkAIyN2HEhBsKa01kJHSo8fAorJEIq8SMNl/MvaIeI2TtoH+k90NCS3cxZw+
9VbO7bY6HrMjUu7ankq1yreBZPhn48Qme9J4pJBHpxFlUo3uQCXVG/ydJ96nAnZ5
i8ksEGRETu0WPyA3e4hYX09POaYr/DoavJr2HeMDFLTyEAG8HFtdJJdC8aMz004L
M/Bd2Gvpkjs8BrfK3i97DyfzkoK98/W6Gd/Qo62FxCnxm0n7bB6cF2WoXASAxGiw
OzEuem3thwxbVVTTbf7kFFnk2qEolVIZzlKrYmEkiHk+r8BpzGBiWjYLdKEUtLqE
HjHtdNc4yMeJkZa9nm0AWTWXQiXw2xrqJmLAukX6x4PIx6cttMSKqIk2JWKjK5/v
kM6Lp7TItwAC6cxsnoFP0qTtDN1YYNuV1D4ubCspdFz4I/9cUSa9K1xsp48T5eu4
wjQv+T6VYg3tNawuHCU5b2QhdAo4hNzf3Md2XY+mrIoI635OcDLFUQ8OeaeGKHKx
XS51rF9CGqfY2EP8eFybvA/cfEgAvCb5Lb5PpBs639CcJRNgtZaB44LfLOZdQ+ju
KZbYzS61TyJ0QkM3LMVWsgGBL1pauc5OhWoLEiLhz2dFI4/qs2ORATsnO16YowpD
8bzr2HSdwpdXINX0+Z75BwT3ZzUKwUgNENsksQ41hIOqAXlVsYJu3nUIwchyB0Dx
IrHJoJ/bgP0I6u3jYTM3wEWZ+qDFoiOAU/WptELW2EEDxdly5Z3pKVTtnUmJR9xd
jhWo6WMAo9yUbhmZfuX6faan+WnDmkCiwKwotzO7+TXD2p4p4uVVIlzF9rcb2i/X
rhzZWrEu6zVDoPwR0BtdHgVRqf9Oa7+ig6mSVLS9RT+kDB5jiVGHwrQ1mwi4u6gW
MgyKuEGCe+9xARR60e96oMF+h10BKDm5CYF/s0H5xQ7eFKy/cHOjgPmY7EDH/5Th
VwcrLLUcegkc4khbFrcyFZg52hDSiSv4eu64NwuWYRK8+lSlcNH7pkHilEmo67b/
Y0zkdF3RyqFQ2clDtCW0iNteNqb0Cxn5SD7o0tmqa2COH431ZGeB6gkVkAlj6Sz0
pMJbBDTV74Y/euDrXoxsK+eEDfIDTHG3x6gwvFqa8OQNCsdSc26XgYXE4XCZegGg
jjjOL9mjqk9xT8Sx5S5nt6oN42t4CpQowoH06W/jcbAXLXKixaM34GyKrpQg/mU6
mCR2JgQvRjwg8X1z2UGT+E9A9mMFRKg2dMw/GqaDXf9wUq11H0hGpUVuMFGJUXV0
Wrh4BXWn3JTO3agGeED+jXQHTl0RgUgSUq0RnUAmTQ2wXMlhI0F0NRmlIoeZN48Q
Lue8I+5+cW7sWZ0MGosD27aBhti+UmfaBOsSpdMNlO9fME0IJ7eJL+9LDI7ExvfU
qTpfQbkJbJ6h2LUw7PkTHqGiH37/rjilNOyDyom7xwhU4SYPLVIKrqB+pD3yAE/k
QT9hI/UeCIt2jmod7g8Af9C6tCe0FRUWwDpRdpNhjThkN8Kln6+bowECy8AUe2Im
ECM4i0EJNJG7lm0fxI6Mj3N34X0i7aob7PLQ4Ybg9+H0v2ZE48VCJN/qrfQclip7
+Mpdq4lZAnDarXECO5Kzi+TmvKBNNjIZeCULuerAaVk2HeHfmHOxMwbG3IaICMG7
Ea0Ds/t4D0OMLqd+zQjZERHT380rbmL2weNGQiLoh2ClNbSNjVpnU3E5dfN92cU+
zii7GPXiYgUgrvmxSKj0WeS1ZfsjbJqww0D1BhWRkMJub3LvFzFh2V6fJBUpju6J
s3K/SvSj1o1LOypwIgmKQUEJXuDgaqgdETs70ycuk62xJspliLxVRP8YuJ37UvYC
8BsKXxPulKeCyZNXN2ThnSo5Ig1kF5uvDU/A3ScrlH1mcyki+ZRow8ml/XIDDXi+
lLPV/fT0hTDhJo1QdwzgcKRuNGDRLf6wT+ghJAqcf2rg+PDPpkRDBR+ejsrD1vVe
LPHd9ojzJ/teZ6WtELHxDVrz45PAeEw3JP4iFdn6v0wzPP4F2p1GoYwaUpYJ5Zgg
9GEOhIzLhHEY2Q/ykAii98Y3aHIGjlglBrbQqMCxYiXNFH2DtGKXpI9YPS3fykSq
TSmVIzULpJ7cTtXTkVo97L7wp7Y3MVwp8Tv/gogHzSW7zCpi1IZlE5WsP36E9Um5
gerP7Xh15808FKYjWWJrSB9tp8qodQ58jzDX6d5HwFpxYSCqU6buntEgjxQik1By
ZBdrFZVZGw4vPTO64QJwbhxm8Kc/rWz7eNkqCg7NcF8YODGAhMc6rMRTmzeU8osz
7RaZ6K1MU4AFNosTQ+ib9KCRUES1lb0QoUNK+9jL6smHlf2XZOP85rAQ/HYBA0ju
ZwfcQFTuqCfwvRgbSxLjiWCABhie7WK+MVHANLAVjFbWJkV1UjcNqAgpO2yeJFfE
eoK0PbYwnGxB75Lc6pUtsH+t8XFNvuFApX5Y8GK6g4oPBm83fM/iVQvL+Hcr6SFI
2LdQaLBwB0gr3id8Kxth1ynBDk8qaDJXIBSq/2oyVo4eAVStdGw/QjBs4Y5bGpAf
CHFEPIzCuhsIFuInKpV/AERIRn5MDWKTIqTUmW7vxZT/KU+hK/fJKAnwxf3CJ1Hd
hbLOWHclKITcwjx6gUn05jZA1Hpdm/RwyBwpy8hzfvcTbuTcbVCybW++hFQjLw2D
Gzgz8WYvKoXZZsPghOfk3MwyyDuw6DMJe8Uonc2qOd7sDBpZEyJqYd0YyJ8BellF
XwegpGabD6DmYMZ9Kcpjp87ZgB3a4uMtpNo23Ir7V4aLWBMOYcI+BRuTL80coyFZ
EszvwT42o8M771iDGUnSE5Ty/cHIu0Jgn9BviKJgbILEgfKlmw9AGePZ4ysgGINR
HLUvjpTlmSdCEQBk3G0sbU+sdYyc+e6J/9QVZd50aJBK3xP7r6VZ8dG9zSfyjTdU
WD/6moaI3zMrW8Wj65naPwK4hy+5owGrLphXpdlRXUYJj2dDJBCN8/hTv84fNB8f
Z+mr7eLpfmSHVQq6erU9w7vzmq5oxb5xtzL8gkQQcnlK9SI3XyUPj9GUamo63vSX
hcHPEzXbT+xS7n8/LHUo7eqGyt3/5qHPNQIreYPbJJJFoW51sTzwSAm80PaIGrU+
fG26PXElmQQ6EsSfjCqqfbBuOWKh6z6bEVOdSaVxRjebCKNp5+FdXI8j5m8+mNzh
qWxO+Qn3IwDDSs7C8rUIwdIVn95ShBAcVZlSgey385fheVUPLo6agNBj34CfM442
fMpy3Kn5qMvC188TVUJcr+3itT7K7FZTs81TYIYBP6gfino5WdNBnKDGqYKiKyOz
v4uhxb4dhC1GdjyZXJ9v4FU8io3lXsUBiSQNqijvMfMVhZg7dmPm3MQogYDoqGkx
6h1+gJEmpct1r4fknbrwnoSA9v1ywCcHpCpCR4QEsR3pB7iHBPCXRZh7M0ew0b7i
xC3n/QLWTd1D8+y+SMQJqPdpHZYmyhyZN8gSHWIPGjsR0trYb33SWkqzv/Kb+ma6
5E6gGwT5HycypFtQGrCjiYR/oH/egAUWPM4K/NDkauonB7OiN+tlwYXZPbj+ninD
+1g0/TvpCCEaObjDjlDhghrsJWQWHYDG6lKeyHF1T660hivhJoXvyKeMq2fzhw/t
ZvCvK5om3yTbjJ01o4M4/3JaR6OnMJ/Bsuh4mgnM2huT4qX2gYSohP3o8eqp9ijd
OsSbtfs7bXnbgOGKnf33j4s9ZH+2EPrbhy5OpdWfbX/cjIlqQ7KfPa8iY93Em/Nu
qL16zG6HIZi2YucNnl+WPp9vE5fsf6TilTAyvVcottkEMTJRb6MTpqwVFB9VzTJX
RkGNbvxP4h93x1FbvHcTvhle9bSUYgGMMx79OuvA4oo1H6dQbkSWuo56djCR0hMJ
Ypqy2c6jhYtFcSo7HRvAIjX6CXKoV0gSMXyP5CzuDaZN/qq+YJOj1+vNqrwmIPIt
q+9zNot6Y9R16Oiw16cuhutmAqNn+VEAjhK6a+OEzLx6aBmY+gEC4AYuoqYLC6vI
Do/Vpu+b5b1Gdi1fw9pGH+Kf5AJQb8V3TLC2g2Qu8unqRVoMyTOslMgYG8Lo1s+V
Ce+CEJuwNaoKQfXVdIQH5/JpYa/gl0lvqQUntjPZxYq8N2H8VDo+NbPMjExbBPH9
ROxHEAHFV9CBNUU9K0oneks74yG+tOHKhowT+JPWqtp81HoARN67B4Z6fnFqfX5e
VUBbFB4TsElbpYkglnKVUw/7I/N+JBZbiq3jV4roJUExmQp0ZrsvARIqXAiqArOe
9WDAEDS5U9cOZ03JQmU7Y9uN1MMqd6lYrShaiSewHK9ZYFNahlRi7PPkSWhN7EKr
EpI/N0DkqAJGGehHwgnH3gfqA+HdqyEOyQc1JgMjP81t8NGmto+2NHnCKc9eD0ZL
JC8dzpj1I2B2hshMlTaDhhlIITgsy/m66RNA0VwYDX822iVtQAoOWMAB9hff+n1E
7znxpm1V3BKmkO0/K7NhrOuqi5zeAwEF7iCK6w3l7IExbeECTyVgaaBTae6awaYC
FzPEUGBjwjxw7n4sPGb+AIcFqhsBwGmuKddjyf9+fnCakmpa78Xc5IvaiPLBQ4gG
ua3a/bW6k6HQMmk9isM0rPfK8/vzmv8vrKkMiavx5dwh77xSyjGj1ukYJPeiltPH
viIo3oB+fm1+mS8D25S6uKjAp5+quQpgQ+5352cMEC0XfWVWUBrchga/71Sw0qgF
1uSEfaypJCcuKEkGAcdYQDFVUT6M80lLSyzdVTV/wtSHm9WxwEZ2W0enPidIM5GZ
7JOXQOt3en2g4MRDZMqdKlzyHIKpVPp5YWmjCfqCmibI9JGY/OojdCiE0QT2XThz
mZztWEnBZyzJgfct7PnfydAQdUeozKDwbaWHTfTDXK6PYjP/i51CmFMKQn274QTg
UfOR6AqZI/pPWuN/JwIYq8vB5g9USDNxbV4Oe1uWKe7R+ydl69f/D0XuYIUU4F6z
4YpDzXS4ejNOSo7qF0xKOG7mpl6pqPuWndeiDo8YqJNcbZe0sR6gqiRnSLgu6NY/
2lT7TnYlMuHHrdx5WJIoRla5XAOVQaLvNhfk+MBqJ1NjsSkyW8oH7uoGEgDxMBv9
Edvf0Se4aBBTTO0qLjIfNnhBHAQqUTTvio4Eo5XDcFjEJAIlXkaHXjwrS3xh44j3
gNFsBiQ5XsJ0yrVNEf4aG//37qBOIcjSy6o9HpCdCcxQOr0I7ulD56xFG6HuvErE
Ds6zxcCuuGmiap3RtyxCnIJMwSwz9KBBr6JlOPfN0Kd+wv/uafJqdUYh7g6K2x5Q
ozGJAayk/r+Nqh/99EeJPAaHKULQJtuKqmnhRT10/tx08dxvKj7hXutktQuv4vbf
8Ub3Yt+o1zJDN+/2xXOFlwYbNymcLznek+XA9QMK+Iq4ONJP5wFOQpG2hTo4lXaO
k8tFiKnton9SnNdZj9y8mzh/jij5sLsH4NhM7yG7DOJ20cnOXfeGI8IXIjIIhaom
mbV5vlCtblnuEwefUhBniYS9DroFL+BF7yiG/HYBTyRHTOcVknvRuf9BoaCYhg7N
9U8Q+qgX8ZcpyhUjb8sgMFax9u8tBAL0I+sOt9Rd7ooqreQ/RC+O2NfFhOH3qiwb
ws5GlnzF7MUiZK1Rosky+GxOWPcJFeVNVEoCPxKzw4Knlqwck2/Q5+V9AXKopTu5
fDzxBi68YwnFBqIqxx7OWrNgbKLU4UxDECGXpzAqzKq7I/jlrVeghA9mPnHExjdg
D8afEALVGTmnT7OsbuqmZUUgUJ93ColQ2T/x+Ggoiv7AmVxKoFlo5V60Z9XOKirX
DpJ1yYnyynZmvgK8HFIikjE5MrQR9v6b+wcpewWy5rHai796lhurarNPtZv4bFUI
Ebo1Iq85mjD+4nojM+ut7naX41rFz2TTEJwoLc6kr4uvUSQLmMVIOrHQgmheBK1M
wo29b4MBq9NgV7ldYFel9OrK8+mod7OocojAi2uiurxvthXKL0tqzqzPhrz86bFo
V5cg4YJB6y28q8XRz9QQ8DJnm84sgZgCGnHldt/SfuCyYkmI78bXtLHOo8Mvm7M/
7jz+8onovu0OTWV4Xu4cadDLT3JXo6pEsO58Di6by+CXChRI8lGSkYkI0t87tq4d
Mv3LLCypqIFC5ZVYidNqq3Y+iyXTzsMZgWCY4Tn6F8jo+yR6Nv0A4Ht8rjrVvIR6
ORuyrJk0sJPFDmDECq0LBYMlrT3wNN9zdTOeClr4Zfg1JJRJL9waUEcRF2HZQNxh
nAi2jC86FOkXzuMTR6L6+zjCbHWuFW+nmSWRjEr/OLPL1h9+qt7mFe6pkQInpq/n
miikkqrEOSKhSmRGBk3mud82CoqOUdBgQBAJ77pyQ8RWRA3fRDLiMuxnNCG8tilP
eOuRow4ujOdgMxaaCI/JFXDKb5uKzGFtwY3uHVc0bW0apnFNUmSRi5z/1XH4vV1S
bjiABcSTZDtn1pApPfN5041b5wGkvhIWePqTeUBIb8kKLoWUfHHYQLLsQI7xnA8m
t8T3cysGr3FHsBEjVPdlpXdXxPu+Zgfz6y3eG9nkFaXpCTAFZGI++G8VPHvPlMSO
Xe+0r7DOTiQlOvqQGBtGs8rTrQq/Z2R0BMb9oQZlUXOMezFA6tlmqt0S+S6ucGru
OIh2XhxbuNaax5pHo424vX2UtpAgDi8R31MBgGQlC5idhVgIhad+F4SXsb0rFbYG
o1KJyPaRhU25ItVAQq3LOdM4jRUB6HzEFoWnSaFP2a7yFmSUZSrh7r2rwUonbbBy
7H05P4BgzVwu6s7Nkkn4ZG2nfat58vxSI7bWjegfIQJtQJqVO46+uCKuE8FiUMw4
Dmjt8WmndS3XiCsXNtn4QOJCb90Tv9r0zCMbwQ3O2BsNYhC1acwuclZRklujzWC0
5ff/+CnfJulV2TodYlzmA4mAevXeC1WGrOA1rUO37zpAo2LUVP8boPjkouQ1+Pzm
0EwdsCPQWYBXAAuPMZkOCE/cVJ4Jf0cLbObpzHOwko87jCK6BbhYHC+4mfw2EBXT
cH7MV+motJEjNqm1W+ghiMGhP58dSCX3Ek9PRbyKXLh8XHqfN0oHdC8NpBckE4HR
IyvkL8ZuPJxF7R8k2jUEMB8dPDsmg0suJKpJIcVWQ+0Y1bR90k0fbR6e0o2UumLc
rIOjkF+zFJO4hy2wE+Djkefr1p4VKaaWAOXx2ifL7UD39+f+z9gsj8J7znd3UZbq
Qwi9rQwsStJQK0iqTR9JY5Y2mk0bKfHc0nJADQyiPDPELILrmrbxo3SMyIaV9+hE
pibwpJJFarLGRjfkzMzO3kaqjuO4a2GXkfPcOmttP2Vat6EgoLXWoCZDPKyIUd0n
qhPkc4a623GI6znuAFag5KBgU0JpKHIUogYuqU8rhWBwB+kt06tWIsp7wzkmdzQG
XuxsKPbE8lrPGwemtFxFafGX6wiVKogp8LGxkN052Qrv2ZfCpBAWNc4qUxboLViz
xRkQ4UWMeFdli10Cq4GvRJPPCWjpLpsivZz64vq9UF0n7cx6liG//YQtSqy6LNrQ
lnZHBW5M/ePvzXq02d/ol8Zo0W9nS/WRnzCQlX4l7d7s6Cs02lZ2o/gTmxF9Qjfp
48vU+qqAR8kffWmwwpUzcDfTiwA/tWT0Uv3K1fkbo2pkFrJrgdMjhawZWDDnm/d4
jr2xkawq07XwG2SHPgEXzhLvt+VxyMMoXspiyz7Yn3WtGt1+7vojZHmAWc3wjpay
gQxDZbYP7bMChHZj/VGIsF8YR/iWJ4wkj1c+/iPxM5fLVGuBYDBa0qB/tMAAoVzk
9BapVvy4009Ls+UMzgLwR4gWMJ4wWkhc8fh0wpSDnu+PAQmpOP1mSkP7Z9bYd1NC
9OwB+o3Y8QP1ogV9ZLzS5yJ7SbiTA/dIzb+nxqPlNVV5maO8/a53JHoXXAHIVhWj
+Ac6H05pw3ZppMzJ8lQxxpxD+vQqmI3Py1WGTHsHuJ+LEvnukMFhd0+1pLjpb5+Q
ZN3NOop3Q1mREUdVeyu1uQMZM/IgDRyUyzpWoDmc9btNx8mDOZkavhR2x0G8yoIq
KC25CbQpAo7L6o1wOyoAUFEpVHXO4a0xzg7/9+wB6ZgpZnU/r0gsYo6mshrAdzot
GXi+hER3krbsDK8A9u8Ndqj3CViImhJOkODO9S86bsXHedtGZjETJB8ok+/zm1Ge
ljQFXs2WpHyNe5Zmxb+ajAoUIF6RhEBI3YLv7GuMMIFOyP8G6TXIO7KUeopyCsN5
ki/A0Gx1kF0LjRC6mteT1wszRxDCEVtAtPuBJhv5JD5l6cpkem4w+lPNsH9ayGOJ
PjysF8We6L+kg8WftIIGqmSVjuLuRk6DEkmmME5WrKr82MX8kjR8JEsYfYyaZjYb
Vr9xP5NLKPcoPYsgDmMjFkUO95dpX8/fbffsmSMYKpQ0wXUcHLXVQ3LRhOhC13+w
EkQ+Q2z9yNJRMV7hJagEDDgJHkSDEJ645rXebxh8MdsBH2JawvoQTLkt9c4AUUWN
2BSqWPLOgkpQonjgOx6GDrkdOn+t97Ewmk0fIYtmHpWjQeX5IfcxLb7gBVr6I65c
bl7q+GGNjvrg+U/OQ/NEr+jRE8updLU/s6yXabU+rCYf73pUcxGshiUaenM/B1Rq
VWL+yp7h1pOB0KxqVZSSRXM4ZBk2ggzgZNgfwaZMnpzCbjeqaKFrl3iojJZLvtRE
EjFPdIVjB28kbpB9ArG0fAiRf/+u1zP2QHQgZh1IDofXt/wsdOFlFkLZqbInHk29
dNAkSk0JasqSzlpGXosbIoI9b8GdVPMHB7nwPgyH448ZR66bLF0YdvOC16LCs44N
xHkolXSXtNEhrvg2XhB3dVewapC2Ht0K5VDYLvrCXvS+n/ij9ILU+x1q/8upw8xX
oQSRs+EF5sJy5D8bhnUkY8wFDbBhB3+WZqolOf1oxO7MVjmC6FjChibF3zlaoYTZ
eh/jnLKWNosv4iB0/7VsjQiVdDwAAYpPuydSoQbiSdD2ToBm1hk0R8eTYvmgs8bl
+VMSWxYZYLjiyIFNVIVVWFDiyhkuMA06ylaGqlEMiZsUMob1hOQG/GKdHU0h18vd
AHr2F1T0CBPyWBegG9tNB5PcIIs7SMKzmFRKW7EZOdzTdyanNFdMfGdioATTsK76
byJdWfWD+mB3ii8RK3KB9rL0CruYXvGzfFs8T6372QZKruwWpVuyB28/j/jv8tjk
hj17KXZu/evf8dQwVKM7i52ZQQUw1atz8Iw8AKAcvvWXO2qZiqAft5dWHBIG+U+p
P6YGQkS2aVF5wkJ636oGvOASjlpQlcZNAtn1hRZOMNKHg5RIF1PkojlQVHfDnEcI
kpBN5PCq9WdRU8fUw/wDpXR61oJIXZpiU+R8oRheEPh64MPCQYen9dRRz/+QXBTV
hIz+JcD5mTExqeKcgOvvQTO7uu5VnyrJ4XZ/dfyva4XlfDhgY8xJ7Qn+6d/FAfcz
YxE3T+wB3aiG6HwnKqElHT3b5+HORhE7tVbolz9d0YlCYxhjpJbsBKBQjcgTmDJ3
E+Ph40L4Til8pPlwckSXXqgcDqd888fDqLpRVJwkMyT9tPSp5B0XOXP02YfbH04g
SyexjqLS9MFw6WXyNs1IC7xvdCs5xYD+btPTfNxWUWBp2Hj8mMp3tqZJiYnL5Rag
7ENZBR0HPkOVWiR0f8leXa6JmCW3zMSRdYt/OY3a05RYM4+SoB3JAqLTxUPin5FA
F1+MEKPGs5IprR8bl/ALRKZsTmP4HIU8qsnZGalBGM8P303XRyFaTWx5HoyukKaL
b6pllYydKv7SYohu12bUUsw1UDhz/lY8WH9ifl53oJ7Ys3ce6xkYRIZ0U5fcq32v
ceCP+7pXJpUvUnlI6t/kpurYLZ9zMwkMFADPnDYnzxy53Vo+0oklNwJfRh9b+qkD
6casZFYEj8l83rBPkRd1slPGFXbHqF/3+ERvbtBW1q6gh5RvO764Pcv7kvE6qMx5
aDjPa7DwJGIOVP/+YvWaKj1mTIjkvquOVBYG0o4qy8Dxv6+iPnTGEIvzFItZQS1b
/8gBK4hnDT/tWNSybOhJvGQyJaUoYXuE2mu0MxRVeF5SQ/VBk6Uyw7rDsB5fcN8x
0FmxlVuXxwOG7O7XLAar9Aneg+Y4ZbKOeP2zc6O6D3hU63WTAMrVYs7Zt6E3dhmu
Eu35ybq0f83dmtko37LShegK9RycWENkeL+CGGnRJchGOeDLvOh7BIMOzxyBML+Y
kOp+IbRMYhdl4d8J50qdKOnnnkiL+Jw/i0kbi8vVuCNzBiXXZNAZRLdUbkDHudgG
OUzfKC3yYLEsByUYyCsd+mWY2YL7fyDDs49sS1L/4SMgbT3PrUJJn2qQ0Ieqdn42
RXKvVBWzK/7tt5x7sOOExUgRC6tSXCLv52R3riputAkWoGNpyIaTJeeTFGHn4HLU
9MiQg89KWUODi6lve5ugiBKJQ/t0I+OeSug9P7hD6pCO+7LkbKk/a14Hay/ST1JX
l9QpkmtGg3POKctC3Rl2MmFagmdnYupvAhNw6/E8nIeBfYKTAuVp2M3i5XhxZUIj
W1JU3h8SgBFhOs9Jn/gzDY5AsJCaeDljKpucuMkK7UA443YWlZuDAPb99FRBdn1Y
pauSWjIW506kPBFYahAhZQliLLlbCJ0iGLR7nQhud4Lc5vavB3UaRLcIO8TDh1as
0YrDdYdrlCTqgXdixNczJ9udyoSczgEX5sJCAZ+hvDjqxzzwuDwfXpUCy7wELQ7+
Pul+gJRclyMnrkcsEWKkIMDYMIMUULXJYqtoxLU4yTrAqT2VEc+rktzciNBbdBKr
3cVBC1wdpNaFmZnMPbq8MFSjReDHb2nFETBkEuPKnB8loRiFYbZE63CU70gVwaYv
xgxfVxBy1x0ACn0hQfzyAnLg13Qp38mHHRwfmV7qtlDW5mgG9PZ3Zc2qttb41yP/
IoIl1bXReUGp0X1VPrzxv0uXIXVgrkWZ1WtbXYRJSY3bD1O/kfdygskjxqD9w3w1
JddxjIL6ziujT6bQNoRZKO/yxQuxt5+F4Kb/S13UbCgnRq5/7qJVFSGPrv89Al8c
c3P+DhgPsU6xxV5optJpo/tDpCLQzvF1yl0qNGOom8BdJDB1q2o2XyII3X6BpgoR
k5TB1fN2R38/Fx09OYqCS6YtdYulOFOJCiELAph5L3xTwJzVemu/1LHACZ5Fl+O0
0K6QR+EbLlt3XbsM8u7awjUxJU4pv5fYZZqRMl+XgpRvblnK0onBzdgMMWZuzSg3
OvO2syR4PK9q29rnk7wcEWvxM4CK+edh48zWpFKuTZE/pRabJw9RuaIpa3xeJZZK
6Pn3N95PZ/Gbo972/9IqmCgBL/OKElwEUCluhbdm+MGxL2sifqg2/SU2xfGnzmoz
rXwJanEddVjBXaA6jHCFXF2gD8h7uQAtVFYLiluAeG0RSjKSopWX6GygF/1wQgfs
gOpW6UH7u7XzuhXE2Vako2b8ZoyVak0JExYiovnWKA/PoGejYoPQR9wzliT2oEI6
DwM5PUjgWHafuvXoUjYDk1Wt5QhmKuwBGQNeq0PNtROmYHjRG5WbduynxmjBY6F1
xjlKya8xU1RW/knJFQWLiJ7lZHEfinbgBycFoqZWmH1E27w8c1ToCWRMqfkuRJcH
U8HDnhyU9L74pc307fwuWDU5hCvp2HmTtWY8nKZrmmV8X8caSyNYwqZp7DN96baH
IQIAtFZKFs2Z0lj6vpwjmqTPXMiUqCT52Dpk/AgqXLGwjRPq7A20jhxAn5ytHcyN
MLJ6PfR00iunseEkI7dXvyLakgXbqrOlzIX0jD58ZAyksZeLzcmlme4PjvViBv4x
FT97p9kP6dpM8PpqebSpkk90gqyiPr+4lHp+1Pmdw3yvSqplUI0Xkrm4qEHj2kZU
0xJo358dQo14UNvKqiWnxWuKYk1JFtU0uXW9NqvCzqmZI+I+qb2eVY3vp0m/4Ciw
uFVOtC8uBekrspcmCG/0cspZkFLE02hlkIaJ9H859FjUvh46AMVq8BwP/+Km3H7L
OeGE2K2PqGJz3O4px8XhaiVfsmZND+pDuWIDcitrFNCnLygUzEgaXYsJHDJecEF8
MJkysSLKWd3s+wRxHIla5e/1kqo1/uP/DWh4RUQxRdQCbHHFF7nXCQBjzghuxRPD
K3m2KvivLx/fOl4CY8gHxkJnxPnXUpx4sFJ4sCkZYj6qIlw2+d19V9MT1aovQdVk
0yqnQzLHMDiTHFffNHApSE4zhoJnD4KbCCDtAFEf6ecEByaB8rm47H0nghxiKV/b
mhhoiRTj9LdwCG/W3BZaj/wVVBZThT3Y/IAy+2feNn72fQifXAs4ClRmbSg4/+8E
UdYJ7MLxiwA5bCXE98TlDxiqBaIX+bPXk0ItcWeuRLykZsq/iPx4Wy/2GDjMoXN0
sri5nTKb5upq/SMb7VvkyHQOCKRFCZRK+gOdc6md42+fFwcVh+No5KMj4Q6odExT
KV5ca3Xhb9nkyfFHktGIHAhLpX+reJK2oNpA/+d81Nvy0Ub6h0K/CIiYPigQTP2J
PYGgFOBfaai2a20QmF8VlkNH7i3o2c83gJaAdBDMTjxTeTgUcZ4BVPqAY5nIhIu3
QGkZJVDU/hKvBTM5dZZLAWNb2Vq/73WGG2VE2lv3tf1MIkRKazBCAMLodppVFenW
yMEI2AIYec7qPu4KT6JvV5AjTv4+4nSx9z+csnfT0Upx5kJjPZ6Ss9840lh6eVEi
9Pwh0BzPzlSBDv/kHL4HxVm7/XDbcA4/hcV6WI7gfty0GI7BWMdhUZkRPMRouHaY
Lm4MHJ5203tAtaOTGY0sppYSw5e5qGBF9rxLY9j2GitAHmzJdFZJ6lpulSMI7taq
iyIE6tVtSJnJveuz3NGhmhlekMBZUnfGeSxV+ameRp1if0W1DHU+ULS03EvxS9KW
Kend/7tkhbQoS+VlnPEETUnIaFN0ja6hJmd4PAHA+12rLy5ZLlq+lXj85gTKMJY8
jW6sYQmJrzcInnaaynuZ/78X7snV8B5uo/umxRLY+lTVCKEK+qrirM22op/bOVhO
M133pT2siyp/C8f31lmyStwtcml9nH+VKAxzOISs8kKGEQGW7GTsBcINFczs5HZu
pkzueeHxsOfD6r3rC4d61kfBWTHIg8ulzVrBxRuhHPVKCT48LRyhaLsFjiYLpvIp
aADzS//lAgIpSdBqjub9nXox0ddHhkIyL7odbUaaJgrmGVtMqgjvq6oz06IWyS3X
JjC63+DL6u9z7/LUgyeqkorxAKA7oIrJ0msrgfTeS+0mHULDI9jzZyM7TuY26fXE
tSTvcfzfQI3JPp1ga8xEyKgBjOnTZXtWtMDdESb15xSwMyKqwXeb5Y+o3bLGwSRv
lUvKcXv2WBTeYaq7X/anJMfPQn87j++/NoKkasILeto+D8gvneXrihZeBDJ32P3w
rjNLHEd6vF6Gv4ElgJ7LPx7ichD7p+PQwmlAj33pNTLZIgziTfrE+0/EQga6EUBH
z9WTvMM7cbUFYihwHcDrXLyasdI9c2nMYzMVg9+NZhMBc6SjH4njOgYdfd/NYTnq
JntiFf5C4ozZUBB9763r/5vgi8eGPwmZ0d7p4dhXGL9Mq3hvv9qsOiTuVXJGcG5v
WPOwRegzfWrcocLVaLE9uSoYlq5AqXUZJQL2Mdb9CuAU0j6K6Pn+CDXxZEYrynex
p3KkScPYp+u9C+Ren9AV76tRz3EqGBJ6Ttpt6uPEuZ/vxxOwjTIWt7jPtJxRQzoQ
7+9ajYN0AEMy2Ht7uVkNi6t07Rv0cj3J+oxf3Vw97lohNQsFr0PV1pRKD3Y6EYZG
kGVBIVtMYxjqGAMTRG0t9yDkPSLnnuG5t584IcmfjwBDsZy8XItaRce2gl8JBH7t
6Xr7EnKrCTPPHhSyUGz3KyUCaLFV7uObs41jFHaR79DHls/henog597vIxK1FAlx
1iEWs4668qBKpB6OvMkCWCEqbj6y0VcH8T7TSG2yqmslsJeebPbcLD6aRnVgZSRC
2QRyLt3FDBWhKGe2++bEj3kqKtYKQcrBgPtgiSGF24E54XhcKhoDFuiKi2bKZPNE
+LAKzWMwouCTtnNJjDECvVKsBl6kJq4hU1390IoGNAH+jAmbyEFnWr8xkXoDgfSH
HpC1GYChZIiE3Us+23JIik3IxmXQwesFOhjVGmjLitlrfGl19A/0Z7qr9lTDFYJP
LYAzyUUAsGTMIPJlwWR3PBdqr4m1uaTKLEl0EGVFOHTl41D+TBDI0kstmRP8Eaot
IXGSj/AO6mrSM0M+0+e3pxoyRD4PfKqlN/8NTdmAMavkrc05sPFOEjJ5FXRDYR39
pWl/nwGkwKlMEsE31RakMyu2kVfFOAM2kvtu3gf+RqVyLhzh8D6bMjkIjt6nC+Xb
kYjxlgFlOI5U1IjnaZ/DnnhgcdOb9q15EYWj1GKyBNuFGYwyJse79zrurDDbCb2D
8oglPQWPwszrRZGE3ZP2OtHAv67Ke2BxFo0NlFtrhNYlrADV0bz6qIQfkGwweUKx
3TLysouSLI1h5n3INPMILh5QUSugB/ixhzxONQWJrvnuQE68JVLY1g+cjaHitIUo
jIJSIkofMlFNQ3bB0IeEafTrqpOz/WoXBqn2q1sVaJGPF3mwYZcUodELu8SmZ9tp
DDUV2B2vQAcTAT5EYfBrJ3QIa6ypkbouguM5vi895kMdUIZo8EWlISEy0KMKM6W1
OK/XWUD1vrkt5yQUuS3Ws6eqck+mpsedfUf7ALxb/jVD29eyJKkKsAoLO2/nJ0hp
sHwG6i0Y7WUFW03bVk6BwuOVr1dDu2c9PJkzBn2gRdSzdZYnjI7V8J9zRNbsF78t
0ZkHTggvZgqyZGVsR6r4dv1bjzBppiOGbUfiYW0rbz9OX6+IKy1RTdcf0lFh0t5S
22MPELo5C3+ZFQ6J0kl61AVeIAewee+2izfVwkOnEYuDc9h8SpdItkuBkx8XNSf6
Q2cLiHPqggRjArHjvBrmCtyd4CIf0/yCYu7TQLuddRuuY3UrB0n/1NSKw3cPx4XY
lzZyjlJyPidB+8+f0U4zIMOLxU3PZUP259+RP3xavkOc+BUH2EAiX2BQ5tf0SHAx
Z3Yvi9O+es+7MhnSa3FClgYsWE5G4UmO8549wbf60wX/EvwC3zK2LIgIbBzFTwCt
skumOoQX6i95V4tBcVWetXleaWFTtY0B6ClYEVWDHoNmX767XLO/mXhRqSP3UALW
hyCimPd/XddK27zmJZQRZrVWusFHxiffy2iwgDTpjoin2a5k4YLvnWCzu6hTydks
MTuj/6pMYSDU9ytPvIFzb+ttDnF6gGmu0tJdaPKZ5nhAp8iiw/UFB+hq+bL+sCeE
AQF6r5zqdvuhytZOr0co2c1IdZiWOUGid5I8UCCoR6jnCh+hbu8HBkw1Ly/7oI/2
AZoYa14EO+8ZblXXGbQyrbqPM/Wkg6hw3netA9wzNarlm+WRytjpqyM9Iy8ghVxw
hjkwAizyCe7vBfKoysBJeVwbyXvwDXF1W1yUTGAP2KwfOKP+Q2lDm4/e+34UmFSO
cbz2NYLreWske4Fl+nSf+lme/pc1xVn0wGDtB2G8MJvk3AR6Mmv5FRZkxh6e/pmq
UZZ5LIL/2E2G0ZhNxhC121JG/OFWb6Un4xtIRkB/O+sRcYnfdXjeUgWc1S6KPyvO
CI81pdHOrornazIOKBFUY7AMu1t+Dr3ODLWqP7CrXg5OZOy8Bo96FAJUri+IjIbZ
QoSy0PPxPIsAdi6k7tdHbMHyWqDscpiMlDsIE3gn6VqsetrvU/QCY3/guYLNPAJ0
/MIfTp9Yjzh2NhurAYzk4zgDQ7efmUMe9wEfLRULNFcJxpo9Tg1YLLJF7jupDLwP
IT8DEdAfoLtEE3QVb/i72fKw9HQS5nbiy7b02dYWzUuXxTUULzaPmqYxTnvsxKnt
/OnAOb6jnkE6ACCXN6wvxhwhgQ0OmWn8aIGcS83L3ZOmWoA95umCbqmMfOvydDfz
FQ7xMJ5/FzRSsuDx9zrEuqwClg+Ow/mqHOHaWZ9JvzSq+V6D0KkhKA5B01jg3ccM
cM/N76361oyZRNCImkm0rHfoYb6jKM7UkglUbZoS4zNGr1eO431o8uEc0dd6KIO5
gB5HjmvIoYK3w2n+fpwBz2PSXKemJEDc31A2XrhaN6WN1CYvRXeGsOTlFqM12Qm+
5zrHA0njjyoUG3V0DI9bKj5BdA3gFBPX7OMC7+ta3F74As8m5xd5w+SYJQyWRFiX
PGJAhM2AbmmCQjewf6cGH0Wux5BFOCyZwue/iAgvSTT+GkZoZZT0x+wVWA3ghrJA
NLBNhGKKQnmaDbERCrgMIEdlyL+JnkA80Np18C2ygfx4AedvaK+EuHZuJP3GINkz
8qoV8LJuG1HQCsjQv4d7LA/5lTPoOu4qe00g6VdPU9efzyWQEiNsCSjYDgKoaxlD
t07z3bnncfPq6IRfchXM081sYtuTTcyyqE/ksgMJNmxUpGpWNilgkmTWBJ6khIoL
6d3eKlfkhrS0eT4XCj2uckhVsLrtvFb+8NP+XrHshXa8zIWE/dQ16GmlzNH+GjVi
A3WTliS597+jXza5pky2hkyyOyiWiaoeUi9bjJByJX2Mu6zKn0E2e+a1sZU6k0V/
WBBUyMIMHb+ps0PElJ4A491foZF1rf5dVud37dtZ497/G+XcoRfw6EaBD8n2dde5
2D3UvOYONFvI6znSfBYHZdTYGGBFKFS5hENNOVsr3dhWnAY00Vsqu5SbXwrxi4Py
vzjlUJKF1VozFHTwQGL2haYLX0jkKniN31HalY/xMnrbQxVbxnkmA98XckQjt6Bj
lAJsv5RZ1DtzDDUmPFoYAuDDPtQwpOk9LdwIJ+lhZWTWDmoUVHhPj5ibsGVH4F4y
nTWsrhewUR1EnLiipb2oNhHjd+7k4kxSoMKkegzc51yPfbxwT4Di3/M2iGdB6O2w
fkMEQeSjZoQaS2uYTM3sXfbTIa63hvxq8jPa9neQLozPFx4BWUEC7X7kSeMrcMVb
WykrohfeY2g1KpxeAPp/XmwgDY0aPJuBI4vBwQUZQp9Vpiy6e+dxmcKBsid/HjKP
L9/Fxlohmd4R1ulfTXPGNI8cq3UxeefL+elXPeHDaNyMVsJBA9T3WJU22frTQgJX
a/00qDy+6/rO1jphVU5/alszPvrs3810eiWNZlXgTpYvhx0NUkZAj8hXqQu78hun
WhPj0+g0HHMhKE8wGUAiHwmeoKuVDXRhHYU0nvfkxRmd7Iewk9HO73RgkrsHdhcs
dMMqDLEBX5eY15zAsoZTUkU4LC118/E6YuE1SnZf2xemDT9eMPe1em9WhTLJ5Wg1
v3hzMgwRsA89VecnVRk2AxrVliSsiGcwCvIcDvnTlxzdaxiCs4KMj3HddQ3+6owC
LPtK0N9NCFCtalUauX+MvlKwFONYiWqteScNnAfrNisMCt6OtDWNMhGLGEZJWCud
WKniVwJ4sUk3mrrdIHqyLNZZRIDp+raB3iQo1CB2tJHsMhHzFcikP7Q733qplvtF
yzNXPT+RCjjjXAjl8GHem6jS0P7JPZ0xfM0+U7yZ1AEjsdJZgMAtJNu5zoCYub3H
E6J8ouixjkobwAwpE4Jnks1GrRxfWuBGwXb9sd3WO9tnMyJwMRh4z3XHJSFofFSQ
L8jKxkrBanZrwsxOuPnP9UohL1ETpTCZUtGGXlb4jkcTBuJ3/JZQk0ExXi4gCW/n
/wbJ56o8GrOTo/U0x45SqjuBetJogrfH8WbRwpTgJIxs0D6DOJLABIjkssE8RSFW
FdiO0VxSezeeQcLDSo7eJXVVgUvTq18jFAHadCiqqq8anOzCe0g6FGzcoSrvACSf
ZBo9TXLSe4O+whFHr/Rx1Q67rPdjJ13nntWxzt9/fypaNf973yihmjKL3EM5hPVN
P9wTw42f+i2c4a5TtJMdib5THIuOMP0PCXMnr/ifBdOBAM7bqyP1yK0aFez/54hF
jafTHkblczSoHXDJrhHcRbdDWAGOoDP4HaIDyB3krwj5lDlMO3u8e1k0nLveLpKh
2jBG4GMK0mk0jsdnSVaZhYYNPjOfWW4P/4ftx7YewjMIsKo2MFVjXjA6mkN/4JJD
Tt19ZOJkAooSPXDxLWQVRIFBPksQ5CgNXRgKyGdoGNd6bZsPHo02KC1eRKE2RPpK
J698Hdmyw1CzPq92oTQveCtH11wvNAE3wZ/WmR6q8fB0yXhyJPFkIEN2cdYG966u
1pnVJws4EdAqQTot9InG681vAVgv4hhLUAc0qv3t+AnpUBF5v0yOF6lnhpA2FVvz
cfx2k4YmHE4EZoEnG2Y6f/sxNQwonHWFa6EmKQ4srbwdO9UtSDiFgsXW5IKwbIUq
qV0y3gQ5YPyoZm+16GO/NLqW6ZKewiy2QTNtTU5EWdR8YAy59HrwiEkfBM4Csdog
sCs2sFFijpNTfETFKlkEZVA2lQ1QQ6VK/Z9ISsxJx44hOjAbTkNDWBhB8DdTyB+h
RI8jipsUNpCbzjY/lKyqlkfqxzYv8PYxUd8XDB8nEH6V/1ySt9IBODol+EiEDD9X
zqoXMgvle0ayEKNuQ93eVDHcC9OVQob+HGQe7kVqFYhbXDm0kxlsDHiva8vyra8R
1zS6kdssP07ef0fGy7AYGcCKMouGA036uQnmooikuxvh22cX21vhnFqvTlGpT965
TznumwpRzJ+mJFf5NP7lZqxaXBd5XMlUKyj9MmNV5/XrI9oPToWVpvgC3o8yfy4M
l56TNOFkAdpwiRM7aJrtUZwXx2MVA748oMaRL8573IihJZSL1zMcd/feMtzlS9OM
k0V10vZYXGqjthJ5lL7B1lgpxJaT3BMjcxqZs+mG2k58z3zMJHVIfyem8mh0rhPa
2upVK6bNleHKCrC2AAnGC1MozIpnE5vjNHLHz7noZ6atWP5KhngyiByDU4UCHz2h
G5JldFotSOF3ohg0CynL6ufkJHELNeK8ZDlHfykEzYIQjJf+fW+7TwXXNzW5jWIa
LDKj2faCJnY3SfsZKv+YfZLQ6NNWZz8iaf3dARjKlbaqa1LmKjPoA4M/gv+iGjtv
z0K4/JjydyIplR4Jz1UoxzLWQMFs4kZIK+H8gutq46Bbt63M82E3iNjedpZj1TMn
mSt7pZAT00XVx7h4TvGJl4YNKF8rcC0JLJ4pPubno6z3zFMCf+bRWKZ3PpFuPPj3
AVX2kVo5bDZgPT8lkbw6cWOjmCAl7iMq2kehAhx1NU+HsfvsTjmfYwyQp1uLH1as
AqXmRmhyIpqn1CIH/VU+Kaa4+BccAiv9G8X6z/QE2tOxvLGiaN3E1IMttVvxKVup
PHYfARwRUOew2ceDfR0/UnYAonoXfvQXQsBL4lia2rPLbnUgylUx2Ax7ZD8E6HxQ
ED7pD3DgJFTlu1L39nHCBQJp0EQtKCg7ngFGqn0Q9PRR9cb+q0tUAdZhC+LwsUHw
d5/wq5Feq1SByG31ji5GqD8ZT3+ij1M1QiSs/1MrbL3YJNLsm/T2YtMFOygaThU4
fY90+QcTvVIw6PlUaPkOYrB9QIQWLr8QexJzAMzQZNkezNBMxI8Jh2yBa8lU6Ezn
9xuTroiOCB3XA7KzZQKkWS2csQx4EETG/ozm0stKzhm63kngi+tL9F/Wo+Ehtix8
vTi7yk0TcfV6iTL93Hh31d4eViUURIRjXTClZqx7xOaK57o/OBGoSB6c7WUqHWp/
1IMYJrRV7dWBqy7fcfWbkjr+ordaEdZFn8MXR2t+AJd9qQiDrm8uT2uqh4J85fBc
AQGxhgRur/7kpFZPLTr2SPnxrJmcO7pewJ310DTBGq2oK6xmn84G2lTY6cONLLLe
zWszbbnrh0hF4RKHJskmfzBmRxGVGsBWRwSNMpY5Gp4OxzB1yF3LfOiXdel56jcB
Awj31HghKuJS9z4pob0R8IA+C6BTk0Kt/4EFPxPP3J9B1qSa/gkzqVe3guPXAlwh
hFJWBYGZpDFDVNprylZ/m1XApBm34+rLBfw72b8Br35/E/R8/SJSdFw8vkmHUwVJ
bRxzfIkKNc5IlJT5GekNoq8Y1/mdnN7IjWKTjZqYJS2Hy8MbBd5ldeAi8gZO0s8f
/Pg+R9ap0uHT5eyO1ugU7kebUMnJqVRq8cEwnGrXJHB7XgiThFYZrdXfP8wogZxy
tkZJIERxM4QKaQbiZ5+LS0xm+pwZlZpt+OJt7nMAu8v5rdFc1pVBcBjrWaYWbBQD
0qbpvnKbyQKwxQ6iNab0dK34Jh2j5kP3nGFDSZQ7hLZrIHEi5SpRqtUFD8zrVW/q
NuzCTNGo5ZJxmbpJ4U+sZyIEQSTQi1pKjJAB1LYAEG5PJV4SY59BZsPYIVjXCcxV
O6+z7FI8goiAJDBlionrN4n7FbPKv7AxsORrOlrbORrvykxsbSMIglF7vrKw/5Vf
xGa61kouEC8exiS0gsgC/ZwvxWkTVarLkd389iWRY2MGJfZ1oLKRGThjg7+bfdav
84paQyEdiXr8UUUzuSNtAaCu/XWuQnyhLALR2stZCcXUI3fXDoTr9yffQG1zC2uK
13V3OU771HpTxPrtR7S9hrwmwggr6N7p6SDG+Z29rJYYpiAPFisHjCKGl1hWPVIo
ekNvZc+EIu28BwTDcwjVdVGjtshYHiuyRwJY38yUmZUQgxs1WV0YR/79pdFicb49
NrGYPg1JYqR2RkPZHLZE7EUBKqINwq0XO1KUsAoIEnhXCLvwuM6b5d2//FhQSKU3
2CwW7aKDgFURAZlnyywGo3qCUybCKbaFOWaoRN4UQKlJDDknA0NbRT11goUjV5Td
joMEMFYEX1np+3Nyknv9ulEmhaA/JKlVhpEfavNZPhxNucuO1pupnIgt0fWfY2NV
gsx87/eglIZjbp4MSKc883jMXdrmJMBC3uY5blxuQAcITK5a/ydwtd3kOeMe51EW
QivSE/lCdO7o8eQ3pHNjW7nRKBkgCgwu0tf6CYVTpr6FR/WIykxM7BaLJ7fCMizF
z52RDem3gPjmYrIfJps/99rgS9mu472KTu04Ks6BhoMIHGmQ3HiTY6gXwqrtBc+g
pBMg4lVf+Y6+1R8lOJASjU0hT/+LvcIMiofjrGgFD6/B5wmU+pdxSS7wqnQbVXd0
zbbGR4pcn+rz/ZBL6VuhS7yu2NG0TucxuBCzQ6mQOYbV7bO68VJprqDZQkhbha99
qM6HLQ8esepPyEy2bhvwQcUlnU2+woE6HYW89QaChhQYJY+67767JYHQpfXbJckU
Jk1WYZxUBDA41UIh4tQ5F13GmyuspsQazJ+56xsWXsgZamoz4uH9uMi+yIgCW/qi
rJF/HnRNEWsUJb/0Zw1fxVSwtQ5miceu2fMIjBmutVFZbgTEGbuxebW+81TlabMB
CftH+JVEkKGBAmv7PSKrqNaCY2bwlg51FFjs2ygVnPvDQAW6/BMCSxVf4Wn1DmBy
cuhy6QbtgXpAxIilfftG7SFIHn0koOsGo61PIL6CRPZpi9iY4dfobJ6V7W5pNaRH
K/7nDAyrhjl+B4vgMaKorsqfp09jqOJ/kSuvhIH00D7JZM8GURW9lYFyKkFyBvNp
sG/qPtb0hmDGm+v5iZEFgjQEK4m6RmRna+EqXeWpMjeLic2nUH/T9deSW+pvx2KK
a5hA8gsSNmKT+6nuLnBSFmpih30aqaaaUFhdqRfORAeS43W0AuCXk4/0Ip5KLXS+
apV7JnY8hEbpU0xtqeRKLWQdllzfG1MDYvnDJpqX7+t3/CBPbpmA4z9pFan/yHG6
Sx6HD0PzKg/bKn/upDk7vD5o4om/GvlJP7Dz4d4Ty2Nhwovg9Oinrtq8OQy3H3Nr
mooYMObCcAioqxP+zUgqSqLYqDjbM1km/4oFoBK7faaxMuGq6RZP8R0+mnM9ITxQ
ysfegh2yKB+jHjXt1jo3WGijriF6mpfdJKnE9xw+xp2Iqwx4hIe4hne3PAW8OjOE
ns9ElliITowh9GnaiSYqB42lD54+PyfUOu1XoJ163CIoofS0skz4OPJtgTHhUFgD
cKNL5ffLbKoBaRP5CHrsbG9dqwOxfhE8KEWeXTQTGCAD39g941/7npw8HJwcoXN0
Wd7Epmn2QG0/IxDwYfJwwd+5B45SFrHg9TSDnCDC3Xdvs4QPGygKa4KqDmZEhqWS
M4NjrWOmnP+krNyLyN8FgGKv5Xj66O1+/rBOk5YUq3IMXu1yLbcPQ8r6aKG9oKoy
lfeamNU6AEj0Byqyxz6SsHBXQf6+DG3N2Z1UrLm8cuKabkDOrJnTWtOBEXmpzK1l
HRm/FkobEsvdncs1Aqup9pSFi5cjgB1dBD02K/uf1JvJ5Lk+7dcWOYimSz8Q0YLL
rcpIt6+aVpdvfxdP/CDeHZXBlbCHjl31c8ZFPaqk68OdnxYFsuyZcTQYDffDWfQ0
zGRmLUkjWToC8ts4wgrLHckzWXAS8cLcpZcxVEasNxGQdBjzrdMjKG65l/KonCWm
+nPs/WWYclTlHa3BL9J9JNe3ezbuOTdvWQTuDQ9wbHQvWp5CAWREuUONyFuHfbbY
+oM3+4hQp1zRfy8lPF0+UynLAYf/vS52I7nTWR6a0uqTuLx3qXQ7jZ9FR0r67Fpj
lbTEPb7rvT4ll90CT4l6fPf0WB6xeRUxGBI69stsqwWLiRYcxAw2IqBoPSEU+2y1
zlemCjY7KjnrW1MyKZ7hKdCgHl02SLYF7bAy/FhI4O80Xp4beT02/WZ+uyyOqNBb
QhqDVk2ViDE8sZg4zUAB6Gqsq9JzixFK1ThpE3jcaXQx7i3113hFiw5cbe9/V3tn
77pIkqxUPQu45t9vGJ+QMlV2mxz6t10cnrHvas/foFyUJhZAvB/YFujBAyamWA53
tV7dMtx6/mWLS7hMC+MohZeRXoRjHs9L4TxPfyjq7+ZT5bF0nD3JeGWtds0sSup1
m8LN58cty4MUg8PbFDNbR3Q4e/egmBeJJH67NBQqgdHdbSvGXWcSmjOwr8vRWbWE
77xuOb9TcpBU9M48ldDBDHzOKCYziVXzbN5M0zW4IM+gdiUmRs3FQfYjQvK3rhpP
tXrZb0F2KofpNr7lGVjU8zp6C3cgN4kG9fHvpfO/hRsB88kzhaXMBiqKCjlw6R5Y
Wpk6KIPI2jKkmPptmQH2fw8kbG3xPGJFqi/hGeuBduPxP5GXJcR7cG3yuUfQPLr6
7ZubwC7NtUUGCLpIIQcz9DdNQC+PxhZ5+ENZJ/+OVWsf6UPmlfOlFqFlxbtTRgf+
Q9MKE5O3q6q+DlNcnO/0ZUXhfLu3GjOJOWvzAfkfIz2Z6YZvRW7Ba0ACISPEFbL4
h8yEB2EK0G1x5lo/PQblBjm5BhRCgVmzEZypANYCtWjlMh+kyoymqEd149VVkCiq
gL4w+MdxNCMPK6yopZP4+x+KdedAK4QyGOH6AF5JaehI3ow3SyBOt4raKb8dA4oz
9Bg46xsw2zOBx4DuTcjrEM0BSvm4Cv8xJO9gKDetYDGTTO1qmiCFLTC8CjJsvHb+
4Z5l1hqjZbtvpMpRRrc4dZ82G7Pn4BdbfGk0T8JY54NBFVweibTQMSxtAn6QzoJD
HLP/JdiSaMALOfBcFRZTuYP1VZ9VbBk5Zi+uBT3hBtBhuQjW8zsPOaIPJmT5DBES
5s50nnryb2y1IMxzy+8/9EN0FweI9lMeDYQdmhoaCdRzjvopM8alqlS/Z0QdyUTI
nsIOJn6oDqdcPmQosGOHRjdjD5fLjpwzM9sfjl3rFI56X1ytesMjpcy4TJAM+fCd
bCsYBYhBy65V7zU0h+HuPldm3RGY/KrojDJ4E0pqm0LQRXd+F8F82B//k1EyCLTR
7FwbvBKPDAbuSlByuoQZoOm6IW3FO1YlhlwqCvTvXq3SsrSmt+Go5KnP/WpVyq9D
ZdyBlpdy3I6cn3Lwv48a0/REE201BkLk0kelYFN+Kvsx/IxywpFoBPnmHzoOfPIz
Eom/m5bSEUnxT2Mss/LWW3CVMZ9jGEeSubfGX4jwFfrZxEAhHMojySYXT+5gFGPE
CKVKFC/XhMcucoCEidwLGAtMbadMwCiXvFrjdh45wHQDSixEhhYxjqqy6jQYg02H
FVbix3noly3I5eR0AyXcM+7KDvQbeYVnd9N9Murbyvq3tYrZ4WWnlEtwEmQRjsb4
6FQjhxq0xOE4lcsOmxNyOVgvGsxVD/Ea4cd5Rb/nzrVJPYRLZQRcrDrPZ1L1kJFu
VUaauoWwvzLQVJjyTBXR4olfdHwXsK7O8fR2wtvnWKKG7FjnkmtYQikfweuqpKgH
78ScjSq4hiFU0KZw589ChC9VwnDnJ+Gg/I8ehNpk/LY5whTyShA5y1DSj6JGxL2R
zELZS8LvB+J+TaTvqmDmndzRmMpAfBH9YrGSAH0LFSkMXoDaTnOFhJHmY2tHw6h1
RALhOBDQFe6WFnAGOSkzktqy5ud4CX/p+Yl77oJjwi9zKb/gt5COkKE2E7eUIMMX
+0srUmoKm2wszdSRCEP9Xu8EtPpNO3ghz4b2iAAx6hNHbzZ2s3KYsReKANWA+f2z
YS+nu/jlfSlzTIkN1n5r5/S6QJ8XJxiVN5GKOpBoLSl/VrFYlYOoTaINffBENq39
5qR36JwK+XUdsoudGT+8xniZDqy3y3uo+exhNZ5XVagPRH+zxPN2No2vkZkQGXld
6d/7aAJrRakPPEvPehXGJENfnx4wci8AsdxoIaYW5nBENRHci8X49yVsZ1O/ddNk
rX7pw+nUGK2K7iOuB6JKq1HsWhdOQBTyHP+jRQOkwD0tBeFxC/1Gj+cfAdCHd7GZ
mDWG6LQC7IDl+1LTdmR5oeFD5qzAB7eQEkPZSAKyfIX/k4/zBm5Ks4uda9eAdqDX
ionaiodLj/rGYg5EkihC3y1ImmSgUYxZXCg+PhzmIE/cdJX+T4buKsQaWhgb8s4v
um13T/5EXqS9h2XyXNbEa8PIUCwSXSdqdJ44ALay1FMkq5o3n6VxqsG/MlzWKC9o
unrYgqflagcjv1zgC2tBZ2z6GMATPty6spHXh5KmUjRhv76kz+HRjIPd4cA9UHlM
+XEjiqCOeeUR4BScAlMxpc53TV47mMtCsVzvp8+uWnXedn/C9qe/77zKbCOT1FBz
kwRnysn9aM/HO/K0AjrLFtCVUyeBu2N5ALhbDhgj5D1ehott7qMVaWsRT+4RuYZj
69mrLDaQMGUnTakaKDIxLwZD9jfzuAxeG0CusT+ZurfeCEW0wRVJp9GX9NbUKUyO
2pjRn2WwocjaF51CyubnMqNcQVR+UUGKH8jLBc6a5vY1QAUdGyGi0AJoOWGRCFXg
wWpA9DAxRHmF4TGmMsRBMwsLKXzXADCB1sarN7I9z9b/+ARMNulJtb4z324QnXaN
5DhmLr1ak9PB3rbVEgz8yibSdIUEgOsVwMvYHsBVvyVAxoWz6avS7eZISVw9gaAp
9M3Rgx24t/XaqazO/uti2tCfHPP70on72MrCXNRQnTgoTAYHomQD4DMKCrLagCDX
ox3o/NXzSqHgXZBHO/F6ywz3VmRBA1vi80VvGKLAoWkw0QmHyMOdB0wWWlUxB6Ye
Qm/JSP2xv4WPnvJ3TpbN66AKk3tYwm0pXR1wPB0YTC7e2gGxjMT9ijo63DDp4FaK
zDs6ZLl4MqE5M1F+GhaDhczEVO0oeKxh1kv83J34q9VDswINSAxyDUijQ/pu2ylc
MrrZVUcAiNBufpdfEb+u5pgxbU76gjpIcV9vo4coIydx3u9RP1EHTPTXVc5w7TbI
pRKhMOud3s4/yNPY852JExXgHRZaCx9acUJDLXrBwfNPVhF2WO1aaZKnxY2+WMVr
quT5X0j4eRa40EEsP0H3LGhWnG+QREyva97X69qDwDUXbKq9sm2jpSzQQoKsgEgm
fRtMbe5L9BUOGTUxZ697VygN2tlqG5UvJ39YiQYE+lF/Id0t/RewbhuxdS8iCTSU
ilb4sb6WAk7BbWoBHKVCeDKsMEzzCqMmEhmnLgf4SyhLo+tyW0QZhh/e52+oS23d
55dNu/AXe6I9VNG4AzFTS1WSjAdIv4X9jeJUIKNmRD7l1pRHFHHnAGM4oeEWIIOy
kB1ArXwi2bVtrjSMSH/lEaQP4E+22tIUQdlnPoWHRn7P0s2UdlHm/qCL3e5b+opr
ynZmPq7hI4XnokNOOvAWZzj13Qk388X3dz4ZsJfrGdTxK6Bm+oiw4dMTXORBoChu
+pPsFINwYWWxfGS4mDpHoEuGNhPi1tyysVkwXkmmB3zQGNgn0+SqiSw6eXQeiZqI
O+W5gbZ7+S2PsLQnth3XtpymN27x2pKhSiryjbMhsGXUaHMwaWiiXrmQhVLqRgpD
5KnMMNYK6KofswMGbNmSM463lTKNM1pFccsYhc6HwhPA5ET99lG8cc5lKcRvTOEl
ovQAt4uFQhKDPgR8Mv5skgOx1cBFw1vQj55CU7TpO1FLXdGu0dxszpASRKAENUCQ
dGvnoN2cbZAFvFiQ31TYMwYa4U9X/oRvFi0U8RsZgfPGq+SSjapRzbcvAs/KmQNY
NkDTpVmJQjO7pXRf5lHidWpbiepoRBpz4kwb54hODlmLmAmghODDMS7pjFPrpDaA
pAIqqwR+dZkSXdAcin84mu2OYphyyinCa/2mSEa4o7JoE+RZQYXZEo6lDkoC6vL6
48OP/qpwI8zpX3fjCd7NMAYbPA1qDauDrqCp4APs6fRIgeV01VDOCPK58zFa5nDC
m3ukL4iMu3JxU6j5gN4BNlXX3+YofmPbnx1wIK1RBT7XWu2WZAwsg72Zyk+rF8LX
q7mP/lmYaqjfDEffVTTRtC/VTQx3c/NTwRbl3HiqOIfTC7us5Y/vjdemFHP+wC0d
bICMIuKgc/jwAkiV6TMZ1vKGgMgnyZfA8gW2rOf4WW50gLqUJeWZ6HzSE2e8aLzU
lgTG57M2hicbv/X5TlNylijXtIfR4RNeYl55FsxwMkd+ZYNdu3dyhIkAVDZehrIz
xcqZcAr1zElzDX+kvoSUkeEB5DlthGgJLo+dwHwVrZXeaJy31nfDhBWoGWsfB6D6
ja4LjFxg3Cdi05qu1teuh2+3/D8A2Miy3RKgG8L8qCVWTX0MqDTJVnGJ/DZoiExV
8/1mduQ07JX5ZyrOUpvAfjZUSMnn3q+316Y2HQi9XmL0Dy374RbjZqYIKyGLDAQz
47MSnZhZJsOd895J1Bv6fn0st0h4U6jX18QvOrG7xcq1r3GG/xpuokceej8ZUEL7
uHf+GZ0kD+Gv6SnbRqiFC9/MbK25H9oH304YXOuH8YMygyvfPM/I/CqoRjg5jSp3
snK5ip3mCTv29duRsmskOzQoqxai2r5D8Zdh5fhWmw/9+TrcPZt9wmMZ1Xo5dqY2
3+/ovVggIGbiuh0HeeGa27+cZKUyppEDgkTngx8cFCTsBREK2ykSk28FmeH6JqS8
XD4TjaKOjY7bkup6LfIoK3HphuH7V+p3JuTTHaTGIaLJ3YYeQfWg7GeR64IORKG0
ePaxEh1RGDy+lDyr9qIgc6CpbeLFN+cIO55j+C3owXspWWxTsjcyyz29z+lcQhpI
3umYdMEDg9l/9s2OkE/KKsNYGOXvPD62qMJ63B+eS+DOwwf/Q3RsU5JeSHcFuqCZ
XQBqdmOeb+o/D+H4rce7Bf4XWTojbsYyfxV0HJrIuxpehh35LCqjlUlm31hXz9SZ
0q4oWAikcQXSRm3ktatn9rHDOCg5EpIt+LuGuzMXkNnmp3XkTgLLNU5bg2gwnV2/
Dkj2Drc+Om6b2TqQ07fYhkemAOFzC1Zep2iL7Rsrn24/emH6xZi/GFjMK78IA55S
4FhDYQqjtaPX3Iy+0a4tmlauLUYI6sCgeV6HcARQ/+edhGmIB9HHsLsc37FM11lI
iuzdmwjwQV5VronKMw55musDwbaQpfRNdKCjawlnRLJB5esYi+AYnoBpm9EZGwYN
l5RI5uwTagwcVkv8tzJGJVUNSlEckkj40uPiFTjqiouZ0/SO+HA9VgA4QWpGj8HO
6MRQ/Q0r+BKwQH8FYOrtqNLBINt4YwVTb+/BvFIoP2gL0C4nbAyZHkW1a4C+SBuQ
wI9ejq8VQUnqQ9XVuickH7xt2A3l9ez8QXkP626+3B48KVbsVBljM8qfJtAPLIKn
4Mc2FIMD4kFQrxFUAo0+EcLGV/MXxDW4Fe0Gaoav47GNINd/PFA09jUm9plNGGf0
AWY+AulF7T/aKkfLGyk1qy9X3UUzJ0rgquJkZ029vcmm+X8SY2R1RbBsYjxwIodS
Zc4YpXZaCrRG+F9cJ7IrAFzwReSeqJ4kv2dZNPGJOzifL/K3paL+rccB75JYJY1N
eowcov8w8rThCbi2HOaUjsWk4Iz/Jijf6Fm7DaoUMddAXzq7v1/oCrTrLrf15CYX
euZlILAVPiRnVXKWkRoK50U/CgZqU5GrkuckwcHxLbVhiyhkqwChZSCbk16S1De1
YlDuvWUGMI28pxVpPMopzXHWTIQoyMERFj1bYhWFuCxb+YwDBMlFYaQpv9ovrEjB
JwuaRNOEc3+UCCClZqZVRKzZ7NHSPR/9VAwIsjmnEQZ1mSu+5UPHdGkbbcHlg/gJ
Teay9kBD7BKUPOnAtUtdhqvbJlCJapBvboLHcFRWPN65OIiUV6w1wXlzfu4IwYBi
uKTU5ANuOFI+VZ/P4g7apJdhN+f42/sBQK2B3z1C/V5vfRu2tFygReS6CSVwXXHs
qXqCsmhmA4Ij94DovZeOeKxF0CqHOhrWS7cf3fHdkjSpjatubMHMqt4bA/fOinGf
Pc774jZ8y3Te5FyntYZ2LZddddR66gpbp4qqUBQym1MRqRa5HfEGeUPIf1ARRFDn
tkf7Hi00461IGAoeqQDObdwZGhk4IJLNdIsmkGpF8QkzS0eqxey4qcUp/H9Mvar4
vXb6R4z4VAvUVIdUhEsaxzP0Xvi70w9b1wD36Y6UG7hMjJvusbEoyi3D6Tl9ctsR
3FpcYJhvW4EDyxmQaITixkJMRCRXfgSKb66V8ZWgWemeYPCiPub9Gu88/WXvcrfy
93xlu7EoneSQZSJ9mQbuXG5qj1Yav0ymQ1tgDn7DnG/Vi+yLB1Gx/SjktPOMcfLM
SkWGQXv9ox1J8DjqI/J7v84gjRntxAGBN5tLoWEYwFFmhCVovHUQTFH17vea8q+7
8oFKG7uwA3p9n3JgrxT4DzKx5VSl4QUCEo9i8+RJ7C2apDsFpQzWz0TvUUlGDZyo
08hlE+VCGEC/PqjPP5qkM6u2PGtVrM+Q3BGc+JU7LsJH65vV/Wu5JHuKVOjew+3V
xs3bzsppBG3WWrdknwO8PWVdu3gAWfWcW982OCKUqcKpupOExpj2kp4BVv5ZSYbc
Atthr2PHYpY2pztCHdxtnlZpRITeWjJ/pGKUTr/+4j3uDo1/+68E2chWOmdIm5zP
WAf4O2CdYEyYqXUmUj9HgAWU3/99niqsoQHsZ6EjfUh3nvvoxXNNd+7S26KubYiV
IPE66KUMLk5SWjasddvh5nPkH0RAbFBon6qBD2NbmRq424RpN44DRo34JNFfGxfZ
9HMQsE0CFsWr78U6t3hoge2SIDP4nPkuHIOx/slC7V2zCSeD9qvVLVssXuv+JIr4
PTF57jHV4QhlUz+GhpM+mGrtSnD149NDQE+1aK32B2t2i2xcOuzQygtXJCGVhgyZ
FtnfxbZHouZNefdHnRl1dWysQ8jELiQrl9VIC/+THoGPqEHHG1I2hB6rhSTYyuqm
hS8Twa5t+asVFqWcYyxR9GyWBN56Sn2wAhi8+1/YIWIaFfegdp+myOlN8W+ctqTC
IaVDBYjVsBvne88kDN0tFyhtMI1hQLngeOTQ+otPB3hvpYJfIWK54JxoOzwB/bhp
SFpLN1125VgTayINMhM+b8bP0lQjdm0iD40zN3Nt43oPeXlXuVHbOi2blAhsexBR
58xVgm8QQVW+cUgA0oHKhedpmp7WTdeLvFwlb+xpnHu8RergsgMOsZymMMp7WRiR
5kwwAVBEVcqJKZLdAFQ1GdKDPQfU40PzrkYBDVitDnM+BxhiMiebv3M40zSVxi7f
vqJPI15F+9mGy8gCiyAwDvpcvxP51IF4k+EOGn5E0sQFK4hpC+x8Wfssx6vfe4KE
8sg0WL4VdXPVu9vwiKtyfgoAMWgQF5DouaqYyiJMWlqqgIIaBEQgQ+lzBNbfD6rY
rZtTEhUQyNCImd1Zf1Viph5FtHV1wts/mJkbD0+fXXvrB6VW3Z1URkvVNNRqqswP
zsvjmTOR5i6ml2riIbpHjXFsGIGECiUxbN7lsZ+of4d3FXrm5T+/5cqL4ZQlzXBF
PKBIIjbljQ6IScjFZIItboLYuM8s+83xn3vfmbDzjAg0bmxIwPVgC0VVqhf7eZ7x
3NxoSu5wgOFHAKgbmQspuKy+K29U3PZd5F3T4nCkFOMmspekY2RFRIZPiQjhfHLI
DlAdZ1klIt2D1Iz73mUqYL0SIFzFVGhNVZ/1DhWkHFYCEbY5SjIeZ0clQxxhITTe
UGX92FmqExr2GqOrQ4PZ6S6Yagi5/rh5Z8uvDfe9y+QkTGZSqK0QG5ZrNeo8j3ao
CqosYA4LG0CKoFJIbbsjZs2cxyK5ayjPPJMy9/v655MU04Ch2tCv3+xby3UHOXu6
xsqxEZROk46L8V8XZh9hmP3RMETCtOK9D0FnkOBOEvOIaO6WilToYsyIgoassiAx
uEnzz5P3K1T2GEPUX63wsJeAxoMiFcxuereSty1ey+5en/Cq1Tzc6411OJYx8B7R
6sOKCOZWA4i6ykLfURFI3auAsq6cQ1DSTw5K0jmbPSR78Cr55hw99omRccy73DLp
zjbc8mxQ0XLOD/O2XpgqKbJnuna4xRxVEqSfEdmn64xDrjU/ge4wutiskFHawUyl
k8n8h9CxkFaCO9y6kMoqgB4UkUiIEOBqRg9IYPkfsup8VOElZRglOy1qG7eSFwfb
ktS9IfuSoKu4OjTueQYVR4KrejdkrlpjXzTFGZA8aWVAcG+dYS7mlo3TQdCMHWrK
3QbtXoyvbuaaEpSXbhtK9wyE/Uip0jOSR9zF+VuwPBMtEnu2jqDHAnqXhkhM7rGJ
xdd3HrPluJcl1D38ojOxGFH18mEa6aEB3f32ceAoXfU+blimjBRwjJTKLa4LrQpF
NvnXxZYYZWCCetiG2gDsZ7VqEO2IvYF9fbQAnEZA8Rg/garuHEyUXizCumPFuPXD
EXtRkmsqrK2AL8LIR0K8MNB1iaCR/2TekxCEGoCYaYHcR2Zz4pmyTf1qMg+z5JgH
rz9Cy8WRO4+8/1iYxjGE5+t53pCDOfaSZuXr7+E6p5t6tP5KavlD4woObQOuto02
xJeGd0hKThclJ18h95isFvchuPWcMzi6xCGnLwZ8UINIoZ2cntyIxB6MLpmSk0tw
Akf34tzCE+kDGpmbtHkuO9DbQSspathVXKMz/P5XmMpEmxdfXTkgTjkS9b7aJ0i9
4R/P9/P875i24DxwUDvgg3vAQnqc2mdM1bpnBmtnoHjTgzzSH8XgMLzUlPS9Fh/C
uMtFYscxd+Gv0+4xtdNXKbnSGr6fnRQfXDxbw/CB7rrvpkerWNa2Dp5kaswZKxfS
477Ay++zfipfc7CGGvu7dewXNMXrQTVknrGq6scCVxQlqk3prCzjI3dvv7tsG0jY
iSKk7S084DhsGBTIVhWNrUXB3A3Mh5JtDXv+1/iRnd/1nzWwvHY+Qwy2h9Jd17qy
DiKzurZjQ0j26y/UquxgNBnqW0p/2NWSrVNsw5LNxaOCRyc1s9bVXdfY1etDrLBn
cZlLIq1LSlIt7IO2Ns7LzFlfzcOynYhWggE9mrh8MWxKb3K32oZPneAfKuGx0ZHT
1baI+QGvWqixNO/iQ2LSekWQaCuqMzstLVOppKkdGzAo0oD75mrL+T32uusiiKDE
/Odd74aXspA1MrbCGAdDiyTHbc9MlUCqjt+9gh/GowJgR8N4W1Uvc9H/nEqErrim
5e8I7pPYZYeignRHpcKT0zQ3WYQvTbN5yiUUY/krHACEWtxuU9j5dB656I/JaZa+
fGfgs4E8cwNVxiL07o7UfkrN2OH/pkev94/PbMjyTRmXf1YXyWHUZQwMbOl09R2q
ueXDsnSUMYJnF5O7XdAQBG1s6Z2Gtek5tlC5H9XFIxoGgR9EYdH1NjI8hxUZUykJ
ganih3I/h8wTEiBNfM7lixfy9Uepf4LGvcgA+LkIuFmHMw23xfbvpiLQkWvX5Dir
KcG3AhV2KOBCBVn2IVPUAdLdc8NK6+q3YkVvgn3fgn5a3go+aGmyuQUW6oEwNqd8
3HXlWrcgcS3ISho5NvcGEy1ZMkoven59QhFtK8KwlfTe6UZZnmHdgDTzmpBbJskJ
NKcYI5mEwYw3lWvXCZLsk+yZaexbPL/vYJeGNr8WSA0MCqyGi1tukipYg9PZmLJ5
6ezj6upjWgL6m2qhefrnW4lJJUgp6sBAmpgme0wv3wga3TCQi5D2vVT+nryaTjxu
qjk7lr+I4rag4gNyGBTKYZ0G/9HTr2IyU8+u4ReHRxONpTAtmOBmYFOkw996SQkN
dv3sEGN/fHkW1mye1LtKMT1xrCX/exqEgRWagB0wH+kvzybSDl+60dptlcL0TI7i
krwbXkjjhnvMPTL6/Kg+HzYXfYNX6XVHffog3rV45M9U3Og2av0zVPEq6dLz4qY6
dm34MMJO24edXjyFIWjyyzU3WGH/toNsRguiSR6Tbf5i5wrE74SkDaEFMW8r84If
1i3u3fobbc+e74dGCiBcaGabi6CHyEwhm0UZ7FPU6ZgvQ1pZDWp2HKbz9mZcCBNT
YOWNbI8DYVTVZQ26mKgA1hFuEVZKuic6JKgWwADz3ZZ+BWSgR3pyN58slfEtQ1QW
p0fCASoTE/aBro8Lq2x0rLdn2Ch1CapXhiZPCKK4j6GLDvBJzNuIteL0MltmzD1v
AW0yvAUiA5hFF70BN/ilttUM2xqv+mR82A4ErjdZaahDFcnu0wyCLMekTi5va6BI
VOXO4UWpWH7LBFaPq2yfEPwY/oO2jvdxmtyzaXcY96aqmGv6wP0/+QRiQnIUlhwK
XPEbDphwOZ64gF9vOvxx4IK9wrC1LoU2riVO31mDF+C8WxDjTS9EpqWrHjEb7nRO
BFrNsDgBeY29/KT9UFGiBC/3g55NuzZjQnE7F8Sz00pcLOLv+YWFllrK+0pcJpY6
9exvciwCyS1/LdJVVkxVyr8qCnnn8VgSzZsxFN+ki9rwHKibgKnWyEFE8nyJ9+bH
+8sqycvVdGYZa6ZiER2p+wFLsnD0JEKYPIGCLRt90nhiW0mB0qPctSiKudvjPCRj
XViswa6nRPHG5S6heQj6ggsAjf3ylgVZoyJvqUMAC1tpV/ZcervU3xQl7WoNemBJ
7tlcp0lXecG8UCFEjql1In5XiF7xaIa2OXrlfZWRyMXP9F5yh8yqUf+K3QcSWqHl
RIjyUFO7YrVpAEqG/moMacTUSq81M5PqxAxe12g6H89OzXyX2EYGOsR0IwtsbfAY
fJ8TiqbXgZXbsgs9UMY0go8WTPEAzoNG2P4LpYioYarLcydzZeNozab5c/SQroQj
71HNawYRKLHp8o65V8+wTxK6gKOnM4paSOio5jzjdBwaNV62YEnZXj6RyndjLJV8
5hJRzDF+3GPtes49yB7dwz8xzKkR5SCOkMn3qhUFeRDYIpn0d6ZL+4WH7IReOWrN
jnObiFditdKtUXcfv+MyB2HwkmCixHoU6zXN7HwlN1ORFu3voWu2fqyn8XKMPZtP
kG8t4k7Cy+Hp+15g317Dmqx17OPONnRF5mZYkBRX6n2P61n1Gj+n1+J4pxR7wo9L
gTrSvgR3GK6zy4SysqKG+OtNBkp0TwlOsuaOHbv6H5epfqabtvD3VJe98+uR728X
4M0GFmNdEagjhJSMwn8J9EweDwAqvJCiwLizEF354btBE9AB+uTJ6a1u/g5l1vGw
jvEfl2Q/EPZbUr4AL9MdmnMkUK/lq7W78DREd+IIZFFwMr5rj3dPwEO6v/ahqOon
c7HVzLNc7yUCTMYrjxaOlriM5/fK403j5RsM2EFk0WOl9Tig3+bAFReGMVfPQrLg
iaQQswj5+RY3jkhRkUNrXWMiTG72XtsMF8gooTDz/Ja/F6DYCzkPgX1FzIfG7cEE
KS/9HjiZto0tAXHhRy1A+L+/gKr/E2WU/3OmbNJEflToheAn7Qsdw0wqxKCveZQ7
ychs6DZdfV0cjkB9wVguW7qQCRCyHYCtWzkz4em0C7Rb6RFVSveRKVusgwQ4JL+0
/48+Kt/nQuIIt5yjYLH71IdmmZr7sMHs9zgb0i16cdc5iYwiKiMI+7xx1QE8hGXR
PlFdNBFl+OCECfrwsdHfXD0ZuteYldhRyvxxd8kK3EaPSHYRKr78DRqLY5ifTAJF
SCnW6LFhHle2SOl59Qm6G2eRGhfHj0OEf67HjMyrlzePBG8wuQO4eFtjqew+cVTy
Hyv4io20fZLtenO9tNv0ugC9oRmxz4XbELJmZlp0a/nun4oVPJxu8T/PQdb2lBeO
k8+XPynDiKHW2zyfEa5vSeWHzd7+PdZU+iYhBcnCmH/AZ2oXhTSNnqBWKDpKlhoQ
0cV45877VcJoAfMFQRxNy3wI0rwCIs0BvSL/KbL/f8Pg/RhSLHoYNTECkHZMkev7
4erIdu0E8638YNMrUPMfnifuPP0xl4LoCNgRhRA5cPaJyo9f5+9LMiB/g10C/UWI
KL60xP/NmugPzgzUGofwrvHZJewMPiH1tkb5eemvDbqBdq63tJ53kaK1z+YKpNwQ
snAj+s888lpZbcqcxcqBXdGTF76SMr1ouohBDGNEyYeuFhMa+qReh2AuwVbj9iLs
QhwoQQ0Dd5zdDADfPfxC1icCuNhA9VSs0z6OZQzgBnRvP7T/NZEunZhwxXRCvXQg
dxAibms9Q4sq2f2/X7iq2/Y7gz/iwpKnAI7+ocr68zOhZg5i3JmHp4bHWYAUlS2+
AJAl9TI8dCEdNNdN4QCCX7Dqg+VSTSYoAklEr7dQ2w/jo21rFqUF4WJ0SJZbnbtT
YBkRiLcxZnZu83k0JAS8p+1TGvotWdXWVB63lPH9e8tbSYgG0QsCCPlrZwd41xHf
jUrHX2DY9PLFo4uG4FsFzNOA95JDGkeEfQ4FJFl6uAlORRA2zYSl2vurpFnH6deJ
WysUwkSY6JnLo5Vda2EoZ6A33+WOJMy9KsDl/gAnZ+AKVjGA8L16y1TR7CUNx4TA
r1fxwO8Z0NVXwWsS1JcezOgvy2YqwpjohpjbymixDOHLGz9krNSCkHChjiw6XxcH
sbaTkROk2rZhC8ynSECCR73FG05xdQc2+ksPU2nBYzi7WoA6CyEn7I/rMgip7lvG
94vDicTF0eEmTxB3HD7b3gcopR+UWsWKoVly+EzPczvECdrCoQBJW4cVq1fk8BIR
g1mLFHBHWSSdadEbIGvSaZ/r4LKtqg0Ill9zGpucOpe9la+5O0rfsXsjR0uX1sAj
1xMMEadV5IRNdl9pgLwzsK8sGmrTfAeawUNTRN6XXdGPaPJVAax/H6RA4miASHS7
hFdQVdZAwdUMyQcnlaA76gJWx2YV7ya/dOFRlBSQdFpZ5awP1Ui2ZU+10UWNwggt
UZ3+JCL7P9unM7m3f27NqpRgatIKOX+NPwZs8sdzFpNgsnsSYLJKHhAfc2wMLMCP
Tuqe0J67SknubiQhZCGKC/cocVbnrXQij3Y2XBayLiJbJCGnCBkVaZDAbqBiO+oy
TjxiNlDPzvdbYfF03FYXNa50uEupyAsXkSlaOjj+nl21OuXYLAzAf3oTzJG+O/0S
OE+DSi3F9WnmVPMT0LZZ4QcZam2G++eXdJ38bdqr24JAVM93pkBg9e1KUlX2rdGg
AlzGUM+6MtwXVaE+gYutmH+sjUnP/gT8/KC9Jldbr9YMrfFMikRn+2NyVPUmxNW3
KQMeg9zS0T1gh+qDdEURuOqaGUXSF4phwJsKZjt5O4sEtVd5Y9znhmf2dOZdnyiz
hyvNZtxLdMfA6WGJOUiNdWKcrHIkoudPhfJqy+nH/dd6JqVMpKo2NX4Ln49AQcmN
oHuR1tdigT03OMuZqNSLWfaHqesZv/8GjBtDpLCiiqXzVkioeOHux5jrtUPq2lfe
iIg/QWrLLdxNIMJ2ddvTRZAx4ZYO4K//9ojeA4wVVlz8nFE2hHr7TtWLeEbeVVXJ
CffU2d1AlYGKXGqy3NPzb9zsUTVANyI26p0aDsm6FfTC0M7KcRwVD1dWBaE3Ghhe
2zsP5FD0JxyOjlBmWcOY6+YeM2pktwsriHxQNE9hVAuoIM2ovJijDtUGpNMXtjuV
degOtQY9BQY4Jz/+RFF/l2zghxlq3S0cTljWlieT8+3FzciZLX1SXHGI1lrMCN5O
FFqgrpW597g8GoiSbirBbPuuIUXPBVDAgt5Qe/6Dn592zZMTeoX4pUmr5fsIPcRM
qmb1eoap0i+9y1g19jHWdxC59VGmiTLSZfLoPp819zDMS27gxwsY8g+WzhVT1c2J
iSLsSKuxgmMlgs4eoBrqXaqtq5k5CyYBacYB09oGL2PYzGHhxzR2rTcURB4eXPZu
fOjH71PfXjsaAGeWdDwgllMcvMyn8xA+wbaAhmEVsvu7YHUtDApkSX7k5yRZ1Yid
UOOxJGyyLkpsdLjvR+lqYO+gD0tmssObRZyprpbhBBXeJXrS9/K6WVxBcOl2FjLy
bcEgZD2B0vA+HOE30ZEAqGhFP15k6muk3VOD/KWJPyVi34axN7QuH8AKCR4fJmcG
oWdKUpRbeedxhpL+VJfGbUuNYhta3FTh4HU9ZAYDVwSTbbYiaHLYlZx8xC4md1SE
9N8rck+KhNCXaa7a8G47oXp4l1HVZR3e/YkWF/OL5i1Jy9TY+drx946OvkhUYB4Q
BLSPfkrSyzAt6plFkC5FmeCo00Bu7yuqNGGhRyGQpgfDNKddRZMt5h6Q8HeYlWWA
nVPXb6u2wHARbMKIPo3Vzbk0ZZ9PYkO+RjjRhfFl0nBnw3vKqAlrPclGduQ7eLDN
rpMyv+ujxu1StjAaCAOzzRGeA5jOfNL+yEtVLOiJKPiKU93/r7cYWq5k83hzxTHF
S6stOIQfE+a1r6Me48tjfdQZp+vs0M0bFcdbtFs3Q5zOZ56JR99m9M3q6+oRgM+7
eWVr9tXjrxoS3i+5Hcle3sz/gMKIw7KAmJF6/dmLmcQSI8wxI12tBNxlrps+fJ64
vfuZqEgeBJX0KApPFwSW+woCNoTgGdeqIfhnwNQOpKOMkpdcyE98PTRzmqZmEnD1
DbFx5lX8aAGr/hS3Nm2MPdsF3xCGOVMPtho7+MF7qUMcjRtA2cOqt4y7xE6PWQ54
eaR5pXCyYBUqBso8mxemSyqawgV8t6CobAzqP+Xs3buG86PgklKjHL+ZWjRA2BPK
JfreSHjDSXNT1kVvNgFGRrE519GMgN2aKE6f4k5DQVjWVGI8DrAVfRM+zoPS0Tsh
PO4hjfmuFq5T3kW5QRemI6Z2jn/u/gxnks+od3zXDBh1Hwt+DgmSlkGVGGW9SnUC
OD0sY5XuEV3poyMQj/POb4SikRKIU24Eb6BTsqonupmh/rKCKzEaLsgnap5CZIZf
BgZKu7xucA3BQT5Kg8N3+CZg/AvkHAD3ViSva1KpzUGH5mIlN0SfeRy6HuifzROy
Xy5KsVUpLkhQFrj9pHMiFr7u/ESU41ydisAhv07LCShfZaGzmn5W+KJNadcKUK1a
+K+vAZSh2rnEBNOwMC++JKUNDwg+quPWECnY/89sZQcHTgLYNu8l/yruqS6thniF
xoAMoAjqVWZDXUbnv6ijC2P2OMliadfkS9II/ckfiRvXz/4ToX3zcq8deLd0MeaR
xzc1+mn4MtS7/ePzfsCINzjRyE4iKz7C+MSjKaqd5MfNZTe0NHFM6hNisNtBsxzV
Oz69sJyw+9YrvEMMbjer4iEQi4ReiaJ9lla08jyBa1PUkD6nomoAK/GE473DNSbq
vBtUiH5APaeFUTQWsCnS+I0KLZoqpG79FIfaeCVWtDYr8og6k8z6n/P3VDIcpY+d
ThR+JF25cXmjG1I0pZ6FAiytHrnovMjPIJWadSlrcm9hQ7ouLpY8YlZ9VFqhXRNX
FcbLdHdoo9LK+/MQ3iyXDt25VSv8DReLi1d8uBwkkPmgegWKUg87AI0P09EXrk8f
tgHA1rUxPCPIAeVAFDPZv2pRFsZkB4Q9TI6THLWEA2bsiFUvtAdPncuCD8VLVy+B
c44d6XEsNcBk/AALjM62YxoPWoeuJhH5nelZna9CoX6+ak4qWeC3LpFtg5XtK1vl
tOnagRzzT1ra9dGg3CKn1+/11iNN6R9W9TZyjyOBST+2eG2GhLzj8BaoT0T4h3EO
dGJMqzC8CxGiuUvSf7Erd26qSPQx6coCBlq09YfdB47QMY806rzBBzAtu/50fyT+
pJopQvPKtjF+tIjo1F7L+UXjstLsL/1pjY7YECP2W4vDuhY8Ecl+y5fskZiYrhAT
jY8GyWnObatLceCRD6aFeDqOYTnOjjkhdWO6kO1TMJ9BscGeQcNDB7St/5Ab1DUV
xYv5CQ/b4HSULRdymMpwG9PuN0ukaUvHuYrYpyueXH97aSG//8siE+IJ/wp/3T/L
mBJRPWr+UMXI62DNwIsPJJEgnDPs4dA8sfVTXE1zu8WPg7Pzqc9diU0GPImYpf+p
67NZ4wd5zlBiBSAKTjqwqfld18a3hG2hmit1m9OeRgbJ9/HZZDMWQ8AcSddQCDA0
jOzn2W9l4i2c7ZBo3YYK/m5CR86+IACwgdYuv8/BJyuLuCe3akslJzNd5CS5k3hr
kgAnBtkRTBM7hLdNRXAbJl7vaARkIy8WmKff2d6S3HU9YkdQe/vPwVPlPRj2RfNo
DuVHhLgPvG7MVXgezEZMUGvQwH2vMq8FATiw/Et1yYUicFISk4/uCXdIl6lwlzRu
JbdJsUGVbYDoevHNlux2XCpw5YKh+0QMUtSxxLkYdG034xO01T3dAvmR3uQYsSfs
RkdxwPDhPG9Npoby9ws2lCpGJFHstVHXRVkOz0FdP6IzlSN5lB1XDQihnOnGElUm
OqebHsk+M3iDE8xfcp9dv0tRv1romx0tcMhOaem7PpKX7LIxGPQt3LSaiQww1Xs7
dju1sNEkNUWm/H/nsvLFTcA4WILtU18cecVVu04DpsO46/jFZNn4pquHZb6wIXOZ
1Ic3Gj7R54Og0b3GnbUhoQrKCkQFL2vuGzFFDCdWS3AXw4R/moWumuteJozarx3E
1+C98YWuZ9NCcSokTEf03CPx6+W6aDoNz4XxLn6InvsKyggbSl4Xk1JjsbbOUUMR
edZQZdqXQwZq2U11WPog07aUkyBgVoidpSR+0VOl/Wxj0xj4chPFxxPduyThUwsH
wdbwU12rWY/QTr8iti0FR2hBifnpOmadHDz8tNxAQEc+r2rRqE7Zqw7YXZGTBvDI
P9FLsy6dNP59nMTTFMlGn93beTS4qDr0oCUTNoA5v/I5YJo3/gK9uTKJbVN+uRY/
imJKy4FiFVNojI8rGKH1QavD8O36Tt0ZGiwTN3fJu4ERBdyWILgiECSfKVVIZNk2
DGrIlxzydU112YV2hqwVYVgXEGASmlxB+NZWavzXLBzA1YbQkfw5p1eN7jUAufak
JMPqediluNG6ZaXh3u9JbDVwrVHTBKfvH6313YF4pqPTkdtTNUaPARfRTlThkxiL
Bvc8RQOd4KzWBjr8ssHJNVe6E0U6qe0kDMKRtCgcJCzJpYgfZunw7NgRKXleI/yq
uZlBqS0OdO++7HyFuphtuG4fAZj2E/Y5iIMaxcrE6TDGB+FtU8Ot66mh2PLKDPgE
8/D/NXTN3N/4x7STMMiQXbYUm8mRd5lVXh6+IA1HyblRGQfpwQwjWa73QB2p0uEM
cHRnevpY/5ybjaN2jhlNDLeQFzXGeSIWEeXD5RqwvxbwIicCCBpu1qcCMQYBESXB
awXxiBTj8foJcNmmszdu9oPUs4A4unR2O5+u+Ys4JSVAW9cx4jfR1aUxvbDhYNqc
q1CaZ6ina/TH7kKiBLhTvdcUFeW5p9q28TcbE0xHN62xiEG8FnYd4l7qRiTq4h7i
tj4Ra1Bxw7c+hCHvmpa8UWiiBGbM/FQlg2UeKQq03cTDbi/cJMaARlvsU6RUWRPW
M+yMRHuz1prhQ5PPvIBYWnV2ItS4c1BXnDZyJC55WmvMQYvWgyoHDqF/1P2uU/wU
KhoLwX/L4aExrAKpgEhI+jzI8z6Jgc75A4YQKWaJ4mq+W1QReIV1ae4LYsNQmr/J
XQjnyYjHm6CNE8lfNrxvIdBs6irljjW6Sb4+P9m9F7kVxK2WsSshqDydW2Vasehz
FjyE+cw55+aOLFrHYkMpdHsz2Im3KYeHa3UFG+kPmByHru8s9/j8ZFsTFdj6iOWI
EVSS3//Gm8KkozkCRrw5+mrEfok5Kpj4Kyy+XgGpc0OzQ7lmlGsslGyNLX1pevwo
qm7ulS0pXc7EiU0P4lD/J92NyvV+pOItp+HxSAfgev6BVsyYDFEukvrETjW4ywcK
v7nJfwnADaXsOS7Lq0L3H0FlSezEAR1Sriw/3hJeoDbdDuU18IkV7Ezvw7BRYZl7
B/bGiYeD2YXzJSdJrLiwn3I4VgUNB1X19dSo455qCCGh+NTSlaJ7vVloTPJgBDnC
g+sHFtyWSYIYwku4CkW20CCreYlKS4SZi4xpngZe5q7GPehaduviL1C1ddoqz3LO
Bl50MifQH6SVGud22DqW3zZp2JiZUHU0oa0ZkIATGE87qUSTMd8e1RlJPJj5kTIt
1KBHEs3wQ+VdBAXK7aNyep6mwTZebERdvzVjQS/E0wCsxUFxFhMK7DtQlN88wIrU
WrdfvIop3Vv3SOwU1nhcO85dL4YEYKmpVdwzANI2uFRDkSKNr5UTpXS9BCV5gAui
T+0N/S82T0x280c1shXpOC3m55yj+VDbnLXGEhiHwy1n8+b/tVcSON5JaNar+P03
lW3jkTJiBvp2RGhSeBkI7LBGUrgHljGrJqaMz7JZwOssoGvr9ULoQGrxeuwoOYzG
nrtVW39f6iLEoPTBB0oGgsjXlZf/ugihAqtn1DyaVU+oNghr83vHzUCeh51p40OH
h9g2LLGQlB7Bk5Jm6Gdivigi0JPnLUY7Q27Ozb+4ELTN+H2G1BtBtsyI5EJyxi/K
j67RSwJ/4Fwxv1dVoeLgvcx/LxnFprIyc/jNHM0QCepoc4fuCgarIeIPmyRSq56E
h5SFSvX39ZQ8nM2lffLIYlkpehX/td7KeL/bHRHQEQP5FU3W3ZFmBAGYcxf/6URS
cyInqsO4i2PjWtjtdspGz53TyCH9DoOe2pvP1xbA+ZjHWxc1YcIt9luObBoqFRx6
5+iRRDvA1o90poy8pZvD49UmSwDm1YMbEL/0u0Uibs6vyKUlMHfUKmRoNDMVj2Qu
6qmCEYL5d9aYVkFSl7WxerHQFLKeIsebvjIZZQFWIDd5OlmOUJw0g/0kIytOIfvJ
fF2+3Ajb/5yfIuAwjd/Y0PQ0c4gtaStsb5qaaK4KkuPiOn+X6kE+nzCyfWMOCs/+
W9ZQCaSME+NcryAdAeI1nVNkBVVJm9v019u1hclf6UFmmtktVgfAF8zcyXZ97n7i
t9haEXI3ltoLq+G/5TbavcWa60ec1850M4R+J49lReG6kO8keoZa+js4cRx2pCoc
8IIfLbTyZ85aB1jNm5e3aKMDNRKD0xBzYzKhxWZgtPCPhNCiN4XVz5mSWXeaU8qi
69EOTqtkcFsZm1uJp1XQQ7wWs0skeOCIOi75krqHXu3f9X6cIiqAsqcgIOS1ClLE
hoLfGv1l+TI4U6/R6Kl814EU5jS2Xk4NRMYw78/vLBIqT3adrVaaH/bxUb0Ul8qa
Xibdzb9x03gFhko6QJYoBzcNgnlVXdDqyd7nNRYgWxgTirb2USsjLshV104c9kKZ
9MTlFkdnDz98dhwMldie2xTAwtJl4qCA6se6CFt36L5w1fL3LW9oFyK+mEqdVQwJ
lwoM85segm5RVfdXoFBiPI679FD03gejUrcAaWBd8A1algJl1eusneSZwPDQvd5t
LVwtJhwAtbeRMROpi4ivi6pBAcICv74ZVsKH0s2IT6TdjhH5Cs4nhivzC8CuMhXr
equCPh1hAnT/yiltwz0fTlyCphDZv2ssa1Xb2nywf7MgTzDEJUiajrPOfN0BOfvv
WlOw8VVWSWjiDggm8ZM2iP61a2S+W9b8gbt3pL2i6A6KHC5I+WaRK3dHEAsM7Rqe
SiF7a/M0LfjqEtZsZVKjYBNDryl+/uP0pvM4Xxd/5vK6ZC8qEscitoNgsmOmu/ng
USnZoxHO0gg8Rda7s83egxjG2nkrywCWpbZyY94exy2RuUgstCc+k0bjmcRYt8/M
lAMdfQjJQQcwzyRaekcnLDTNU7FBFkJjkAHAjWS+NqMaVaMQVqzOQPkATDdfe7EI
Ar3BvFY8FM3eSfjGmrRu25nIfWsvCux/ovhfjdequjJBJW2BFqIlIlQIMuIgI2lz
VPu0WSQnZD3TDRdP3iggxY25kmvRlHZy/3e+zgcmqxrQreXVwACRbwqI7Ih7ZMnI
14fNRkzzYKBQanqAu//E3Sjez14DEXTbVAllgAjfykG6K6zWEXfoDk7mlQAXPzPR
vyO+LkMdo5IPAIR6Xs38wx1I425q/xFGpMzah3JZ2l3BnKgzzznM7jDAI20q+VU3
nUGwqvc1H4MpD7F5i95rcfLACJMjQp4hOJtjWP2xdAzVsLB5TsrIDE0weGiKR3QQ
nGUPlK6nfe13MBU42G6S9xwBxGBKZCQrmOFIviqufBOXJ/kZ2FCjww7b47O2x2x3
KlO/r0y4c105Bg7uwNSr2oFvRBmejj422Wu5do63F9LqnDSx47VkSjcVEdJC3uJh
2A74WsCTKruosNFzUwlT1Y9GcB97v98MbtLhbwSMjm7QE9PrsWmHWGMp3JpVcJ19
2IgAwIsVNw9IzVahQJ4KwzXj5YCokTNAVRYtWRl20h4ZMmiuDr381MtbyX8+3Mu+
BBVQZfk/gWyXT96Q7Evl4p/Xl+t/eRCq11/2y9NXOwswJh5Nk5jj9PSE8GCHaFqI
6Zef01S+1c+yX8hhUd+lU2at4j+KvqXVfgK3BUjmHjcMSX30fQcpL+7Ps6+JTY4z
SJcw868nWR8DEw0c/AyTDUj2yHyVJ9/LpsBX/ktRVyiEiuigtxsbPG4OOV9LV1jn
z2cPB+QAvzN2XHxL/Fvq5nm7RXYC5nQHkbMDXkUkPnMjZlzesLPZKDKC3ZJ5cQty
6bEsNHOuAfnIXzcOSO5DF7RRqGpwysHKvsYZ2ySB4xFC0PhCGZ+T8+Ql8NtUu7Hk
3iQSpg2WmH1hw3gPyee1BIQrwXlxfN3G3hx2qfXS1Ch7hG6m1hkmLx3Ws4C2DSy5
iWI7WTOw4BgcascenedZfXw7dGSQlQF7CtPfxLJAVdYbUMfS5A24AKpTzbQUJv0U
1QDsKc0wV5qqToCgYD9rAS4UMk9ECV4pDv6K0Acr4x+UH7PtMuQNip/H6mNRPZVE
2KtNJX1MSW6QTG+ULVXLZ6xwYG9svwqYKsR6//te5rAAdI4BOTi3IJXhotXRwzT0
P7nYadvnqNi+zAgU5xUtXXpxMmFcr2/NqCR5oKdKf9windAjh3a+gP+7JO64Er0P
wspSpEewDPUwmefGAQWIT3s46uR+IxUZQ6Ec36rRtECnXI6l5CcHrdA1HpOaLnE8
kBky+R25NgmemVZhVsI6bs0qz0x4OsOKZKWFirLQxfWdt9G24TdEAw1NVde1UgFI
uPZ8eKgAFlLsfgGUXKBLfGStdiFWUUwuLzh4DOMM4KIMT4Sp7iDD/1pxoM/btaOd
5nm03SR4J5i5JBGcC6tkd4rIV3bQND42vWtP/dFUDQlqsjK7uNH6ga0Rwm2YLhWj
+BaHWKJVbz6GueNOucxrUYRCbQsyuKR1VHbhwEOL0J3y0JGaRczm8YP7aD8GQCCx
2B0BSz/IM1EalvmOGhunrpGRd09NLPh42hKzBwS7BoXH7tPFxS5fIkz6g6SZ0Yog
kNtLMmuZVtNq6maER1Vruopvu7c4y+gd/MT5GgNoj00i5v6IDs7101I13FSdhezj
W5yt+qEflp+yp8WWlYf3R/lfe2WSkkY+g/lCA9wMsNus8lMrU6ZLYkh2jpd/VIN8
O8qTv+cMBD68iALa1Lj634wF6aYaCwyGJiOUsiFRMZt4oUcsWWEmJwJ7Cx+2HouV
LxsLXzXvNJNNhEexd7fsr3vSsMub0SQ0QwxgGIF4ym1P1dJ3O3Auqwl9AtZ7bZoK
p+WhOJ1Co4BgLiT5KRSlHt1PxVZJ//5PiphkQ3ERO3vE1DoWhjKMFRkqArXx4c0P
2XSwcG8n3eoQNqlIWzHThCXR3Z2sWnmvTMu3nVTnLFHpaK6kBrZzuUT/Ce85uprO
0A8+F/izCHRDKR/pcd2jKzkcUkaXBcfHasnluuz/N+0=
`protect END_PROTECTED
