`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6cxoeg1+GCUgDVCSWXdW235JHE8X1TxAdkLffweQe9k6UHP5WT99tPLLIsm+6mK
UTDclfqNxfMPhJvCPODgqRh06SzKq/xyC3brJcYPc5wFm1T0xEIKS1Go3Ha1MhCo
I9OgtoeY6iQGmArEjC+7IprTqC03kUGUC34WplP4eHLbCjPgxoEGjE2GxKHJHEd8
NSBFhAgeYuW9AojKqkVRcSvbIBIv6g5eTDCUh4YcXPvNP7sHk6cvValWN9G2IwRt
10Km0DIKGgaVaTywRzP7i0X1Qa4mjNk0QHZEZaZKSeooWAHnu/CYT0u+wsqtlM3F
aCxC/wRDtmAxQSxZBR1BpndskzD9tg7tcao6yqqQBlLRLy/c4g7cozsSbZZmQ8QC
10VGZMp6ER+nUgoq1exBS0l7ULue0I7WoX331hQAg8u17C8rVj3sR8TRl+uqL4j1
ADSXT6h8GYpsiKrXnhA6x2vzxmCcwra4ZNPy1Mr/TGTpvjl42d3wHKjF4ahPf01L
`protect END_PROTECTED
