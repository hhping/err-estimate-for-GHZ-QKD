`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iPPho5zluiMaKKerys+TPR9njjnveGt4FH1SFqpwTMx4yFVGVEPlKpLSB9jG8lgM
EDqu4X9plNkv6jH43hxh72dn0x20nnY6/mlAwz8D/6j1gWVUVHZiy5QfpueumI6T
IPm0PBOui2TRub7NwjmMyb6U8N3qTDAUAqRSiqW7KJdHueENcwg6X/y6O+sMAAwp
OUNTYcLMZ2UcdbcbY2aO6iFF2CX92qn3Zeo/nA8FXHlCxzIN83E4ALeY/yOHPaPn
Flurg0hJ9q1eCkqjyVjfXlYGK386OAzI28cnfv+NNUbB92ynnzfH8mwXPw9hRwKu
bqA5w58ycecyJQGzab/mvI3ENhbz4daq3XWPGvMV9N0pbfP9O0HbNlt4t02EPSh2
hK9nKEDrXpQwBKtyhDeYZW1RHUVTmxBSeILVE+CJZxfgLKcNcalAjDyeeob9HLf3
YW3rtlitoR6HasuIbmjmE8Ze5SW+8ruT+6gWQcKS4xnvKwl8AS9zcQNDzWx4sJGk
SqPNne9c4wxdIxLgg9kUlTbFzwjiakDGfPvBNiHezzfFf5bsFKlMfYSIpTxoXiG9
jpL752jUbJxtWlqNb3fXeeg/oQfYC7h81MB5zjhyhapv+crcMPZPgmSd46PzPPlg
GifDxR+lFXMCU01c8CqBlA==
`protect END_PROTECTED
