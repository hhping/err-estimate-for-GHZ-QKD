`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jpVlklLh3Q5lxniqtFkyF6GY/XKcpywDAFZRnKIRz2ZXaOH29Kh7VGxnTA7Ikxb7
tImIG84Yo2qmDYDDF4x4AGUMmue7rmDZ507dzTliIh1sSd7PARUqEocDk2LSzeID
tuz+yv/1oNU4edJxSGkHbRr70MZUpKY5ZGQtZlI+SSfJL4P6HMbgzJceDedsj3s2
2Yr7aw2FhSngtaiXsc/SWJ2UMRsAGCxOMESuSOEq46ltHIxGZNWBO5GNVm0hw+Rv
v5T017vGymVLmyBcQqGrMOA3nQQlL8/WzEgan2B23wkk/F8xRgoJYeG56YZeF0Mi
RpZEnVAq9pfjhOZzgkZUNnqSqHBBfWSFfLUpVVP7UTMgX8dgP1AJyiB93ardyli7
hu21wp1c6T71tTjB93tFxfr5WIpujuPjKckcFoLB0l9X8jROp+J2BDfGymiaQz6u
Bfle+kswqRIJ+TzN42xA/lOvUNFS/lkHs1EUlaX5pNS63jBoH+EXeyp0vmnatgTB
HURm4g43ZFX5EXW+T6vA8/TZBLso/YSV9mszfaxMS50/BmkxkiY+wykddlZfALWG
VYP2hTPBS7LrrHfhitHnxwTb4vAA2tSSUnGBMm1e8avbqO1TNZufX8UOuJfhso9q
1Tqw0GN14Ip/5AjMQldYbYKZwHlVV3YB98wkxhsKDA9YDm/DUctEeKjoTJLq4IN4
oUGnF9pzmxeL/J1O2zz5hX8uawKr5qViw1d+hVou0ShGgs59pF9erRTclBozusUl
0e9So/dRo+ZHbOvLuRNdOfY5hN8ZJomdBrkFJLjKiJ1kdCgKZ628nOMsn45vPU1G
jHmgNyXciwCZvNg1o7gptvaQIrTO4WaNoj/Wz8Ygsc2HCtGxg6yM4NNAq8wQ7Tnc
KuoKD4a5ggNIY6QtyBawJ4eoR0s0qElztembWJwoKqU2ZbkylnIKXceFiCGGwjLQ
vnMXrSYuN7QTcvUjFKzfdmw/Y06diFBJWRRm5sb+H9Ik6lm3QUY/f+u13/JzbsT0
kDJTihHYrY3VqLzHwRftJZGjdm5vJYJGBHk6xMciIQab2ARK0VmCccRME914V+sR
G2JGFM8oy9eXTvQTov1DpLlXy3HaM8Fh8RRsTMKNrqMxiTt/AU7iBopuUWsBC1a6
8aMUcDS8iOlQuZjFA62YhG/qiiHBc3I7YUhtBSEMXYxNx1MOgskQTGRJCj9a372A
HvWRXJ9sTS7uV8JEMZC8U+uiwnkaF1hrKZodb1vnPzQxQpVt/2z31ARErf81rBd5
1GVil+HrVxd5+31ZN/h5DuldKWSG3R3vORoC15K0zieiPQxjEAEN2XRdWSC6QfNf
HGHxwHoZFgryvNc98KuwbaSr5/gORGnl2ax8VOKAaigpYT7HsseZA1PWhsRPLUK0
QYGVzYxKMyDf1o9m+uaQKUhyJq0s1x2brjgtfF/7nIxAiBwt8M1agEYBB1fd4q5h
plrRSGEWS0DwqLZHdf6ovfSJKpBd/rfq28OeM/TvK48rN5WDFChK9yVaQAPVBHci
pE7vrY+Bfqh9qWAoLPCeMio3LTLXe9ooCplXXWi+DcAGWUvRY0rIP3EYKriPf1vM
v6hpYmnDvXg5pOgbx/Y6ZRC0aj2uTQFwmRVj/SQyfZcfX+7fIabf6GAhMyqs/fFh
ljbn6GMeo4z45Ywla+H/MshmftFUBW0FHLSMpxJ1ERI/DvbUT/IEMcVh0QqyciTr
WCChn8GWEBDB9CT+qLbvjcuWyT8lQ8pC88A2MDV5WKkkWNRizB9IEPX1gd93r5fh
GYGaaY+E8Y5k6gXlgu1ufgTBJdi3FtoysCWp+VobaDp1JnvWFi0wQTYKHdtZUEEo
Lzi363vDG/PzyZfhH+ygzkSmV0kYVSODjYP5OtxflJelk5LlHEkJXKPfsRmC0QpD
A/9+RBYpuJ4hfrD3l+nfgOkLwR2FQMuehohl/d9mVLM=
`protect END_PROTECTED
