`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xg5QO4GqndOAsjLOkS2zr7GehQPbsffb01f4obtfRukpn3GGWuWEEAHQyulM2EPV
YOdLtU3wWOr9xTrkPbP6/N1OQMCwQ1IyrtBgKiZytK5l2UtiVx9cBeL2JFTzZS6t
dc88c6o2ow0AFzYdM67SoJj5qYbPAFLcPbqfBYg0Hb4soqdHAvHUwK/CTiKJ3qOd
/TVlLLK1mBDhYwjYNXYGzfFcp1vo4sfmjvYYJWg1RyE087EbrmxIBDzdo6fIMeOk
+JFYgOJ0QhBjnYsTcIFzeLweom2+Ln94xvVXYJlbrFDdNAldCGjpfIrcYrQ8dNLu
+/qu6hy1ZLANaskvwX3H7g65BTY+q+lGwk8pmOcqFuzfQupu5VIWMg2qhA+K448w
`protect END_PROTECTED
