`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9BUml65WnIc/o34dmBMfAeQlBgepXZ/OITbZ3Rr/MyeTFG87bEDkZlsocmZmTXYx
Yfew6ekJ05dvya0StPRz2ShVbViMvO4V4NcSDw8jUYI8t0TLXDYmRfn7vv+2KGdE
uOGawLyRaWw/TAVSJ2DWEsmSBjF9HjUnjG1R+KEkRG6AVw+1stnl4NY/W/KrRepA
LimXgPsGVwX2ADIULL9jlDFHjZSkbwEP4QhYyzAGi2EGD+aaOXe6F1+t7E93BIBf
XU5ISKrPV1qOzLvwUwsO42Js5dU0WFARJsJQXh+EPwKjxhLAzIODefTJXYYmhUzj
v5j4FPPKtTDANEqPTkeUyisoZq7rsV/LsDiLR//LE//HrfM3X0ArSJ9yitU/1711
0DH7p+IR/i4dBbURn/43u/s8roHyy51JQq1qU3B4hIYlULkCRAbsPhq2pqR+AO31
K8/KtRWHBVOasbNo5Ls1CWiIY9zyex2zgEX4K1oszjReAHW6oP+suyFwdprglcFy
z2zFpSnIVUY5t5TowoNQlSA7GQXftIs2KbRo73dYsDk=
`protect END_PROTECTED
