`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QFlf+eEwnR8+0/90r5aNycImZnNI2PEcQHPZSxHUe8BZF0N75WjHbyNQAUAFgt7H
HQSEWWSy5u9n2HPOsAchJnGaBrSutSdiM+CjGxeVvxRtTqPMW8eBScNVce3MSj4A
r5UhtNdRxItDiDaNeZg9LPEEI+ix69rkRADnxgwsfgWXgieWVkOeIkby++e/lscp
1YmsPYN5yLO+bNvhuKK1UlpKpHGpLGKZTXz1AYqlniKAGhZTWaMzlqAOc/e5KRD3
Bs5ZO2ejMkeMso28Pno6UZyyfU7KAoLRnyz3hah/3MzfFrzbEWVJ+w9WXO4RQWhu
OD3UK8vWc++wdfcYc0jJfxdj0QG5JE0VUTIGoBy224s1hgLNCGj2fyZBIVojhnXx
/kmD5PbRT87++g+xTqrMnKU84wqUTM0q9LXivhMOC05yH0kX/4QkTdIGtwYlEGBk
EIom5Yv8b0dUa2Zw2qPe6J8oAiFqPUu+prII7/S0PQfnoKFbyFcsQIFGb8N/Q5zK
r7ysmQhgAkr2sj3GaQOjZHl0H6XzP3P5hTfC/A8HTK4nJoJTeGkAuUcWA3s+dlgS
I8MYdslTzMPppIoOFPbe97nyNu4sl7mp/qsLXvZeeviYhgOoEPxdjPBndqmx6NoL
OlQLETVQwlezOw6VdSKH115tiPa0Pyk+vvTkME27bwduDotjrBdWgawnt5at9a5a
N271+teLt87CzR0lM/kiAs0ZhDy3h9nRbNQ0L/xOmT/TRmY9q8RRCDTIALcHPeoC
QKQXhYH3vqlTG/kzX+WVyS/dz1c6EWEeejl7N0kCxbGwlLpk0Hzbiueq6Y08VgYQ
x8JA0n9tC7fjiHLVeA6sbS6h58Y9xFvbFYeybVNbjZbEOAa3IilKbxSSSt+UIb08
nMyzHkwvBrHKqkS/Gc0VevsEdcP+daPB4zljN0sIbqh4e9hGc+8AJvOjyntlFhGX
`protect END_PROTECTED
