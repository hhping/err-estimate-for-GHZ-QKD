`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOXq1uExYkMszzjwvyKB3GnNK9Nl4durezMGhvIsbAcX4iGgdZZLklCnml9X+2Ow
DhQwAuTbzNsCQp16aJxL+xIbl6KZCqH97nu4e0kGqKe1yw+Mqmu6tpdrEjEZfrZr
Rr64p/YLcteG8Ae1EJmFg0fflPHBHqGrwgsKxAN7jdVRlL6mVjrF5yZYUmbVw/T7
1lbtlJ8KsFXmmApNwFrslKp5chD3S5VkH004R8Gy4FJY36Fl0Ysn5Ds+s7e2WnkJ
8rpWK7wO/tGprnLs37MmTwqKyO/Y1xdUuwmJ52RApaogIeLNRkQXyG6qUqZKBUcr
u1aB4sFcG1burhq2qxdB1rMrvvVWbylrrpzvCalgssag2N/fYPpTMnFZw/pMdORf
hXZDt8YGPmnZryZ+eXQZ5lAcB0NEgfBdSzP00Fxur5TbjCWSboT2C/Pu1pDQYbJz
sOy5eaaNvImx+H4gP+GLJLC5T2URdKjw1CC7o6RNZGT/BxIXnIAjjSAwWHyyjNYL
WjcDMne6MBJgrSmKkm/OufF1q4LzMa3UistSPHYnf8i3ly2+Td0eEJ0Fzyfwr0fN
oG4cs07GkGIPR6VhJ5wcKJFpcfy2jUE6KBixQHn1okEjuTabuVfktGXiC8Xb4SS/
Q91PuzI9SB761KUfmWrvERT5S/VvpoclBvn8IrGLESiNQMsai0T2OL6wbfblgzNZ
yKt9Zyi/3j1C4yuBDuOg73Mseaxgqc8tzZUh5GsFQn2IGFHWr8S3pXXJqMlc6mg/
/2tLccHaBYeg2JFVs/zMJVASNhsVYZ/lYLKSp8jdc+ilDYHOdhIRUHOUl4s48i+y
bSTz9RJ34ylnEwKsbbHP05jEqSZ5zBhrLy40v0d7bXhOgeBGmcGs1IRlQgxI4rLV
REF4iKzg7cNQBqf7P8FnknYaWY7mgiOLiQhxW7rdGPc5zTBOCjsP5kcbiA5McKDE
mwMliTB+NXOHxPPte/2PkohH8YCKe83SWtiW8+F0z+kIfEX9Wmee3eBnxyLEenRZ
/fdAzEw2ltR7VNk9Z981iERB9qQHbq/jJcqbGNg/bC8=
`protect END_PROTECTED
