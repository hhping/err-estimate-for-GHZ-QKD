`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P8cU+rB7vlmGdYfqs/elLMqH4c1surqmZWjav1a8fOlxfScepIUeggjrTX9hFt+2
lA04IpDAh4tKBUNhI6VBJipor7cl8JUZ7bQKiXuh9hqcpXadLH0UZVevbG1ebX+j
1LdRgakPdczp5smYH/qF9uGLNbZKAvhk+1u8uU6JoVvMNAO0J9o9YQt5r7G3+ywO
HoG0fGbURE3+A/cBk8GBqTvr3/jc8pENrI/1ZNuckbFfr2bqoqihjeU7b+rqTf/L
EgFK/b7S/IkAQwgLAFlmy1tFMCgRux0JGZQ2Cx2nGwjIgocnf2to2j2P+H/kmLaW
McTPWaCj2Pa3c47FuBLm6MEB5zsM7rpjI0im0eNErXBgjkC5qCxkRWaptTbOVh2B
matGKdqIW/3EDIoh+rpuF4/hSmFValsHVdApwRobTpQlMKDVPNMUjSLMfWF4Tq6s
VL4bQ3BoCvHo/4HFLUs+hd6U//fxNmKcPtNniacxSPlJq4E7jHUJOwkNW9bbOhxc
OvMckxF7aWy/SpsnCp1ku7iN9i4ICEn8AeXSge2+iRxUJuKFraTe0KMqzQGEZrDE
ptamzVT132X7gGzH2LhVwbBR4SV0FkWzwB36+4wzeCq8Nk2pEw90ZKeaWvrTavUZ
fuXCqsxQK8FEtq7M2B8Kgg==
`protect END_PROTECTED
