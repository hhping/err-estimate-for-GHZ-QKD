`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZmSyA5G53iubQWJdylwPER7FI/a/r1uhuftrUFhFwvu0XUHbxQf5LyHb7aVncsY
+9vU6GcE4o7wfZN/AcwjyBTaE4v1Zpgx/+Y+lgSUT96UzvSPBywlTnR5t0ltqKdH
ggZpw1dxeCUCbRN+9L26DIuvZ128512FeNI2qyX0r/zABtysegesu0tFXTft1hLo
N1oEkiC+8mbsiWlIkqxpbMHvaaZTdrbdJ/FxaaUm8YpB7aah66P5orkElLI1GRRS
aDcC9wr475agnYv6w6vaShZ+TlDAjvd/2e4NVQdYo8jg+1zFwsYrrWfRBLrkKxSi
eZvgDEAYn6FuL1fJvcVX7L7swc2Atw8GQ4Wl2TMwi6BOp0fPS9cXj6YH/gTeySR7
`protect END_PROTECTED
