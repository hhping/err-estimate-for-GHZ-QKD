`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dAC9MfKccZl2ZbPYI89q8dccYLGHq6KmzCin1hHnBvg/F6BIdMQ+D8LzKFYYohAG
J0bpigTwnF6KWKqGcvYuJ9fV+E4S0lJ9g+ElnKTpgvclSAugrgfQMI/zSnqbHq66
nrV6Kqa9KE7iFdoyr/+SJkRUJAmO8iShnBYrqz3xBrZfZg1neGd6bT8465PzRrRb
fPChphCKrdSWYAvn6ZYAsSuK+Glu1AS2AVLeH115oJmTCddXl79JnlK/vdnTEJnO
5RPa344ulVQE/UXkZV+EHbV1KiQdBKvfxHkXFfuyCq6LG4RTt4ZvQ6sZKGAIsJHh
EtSeqZHEUE4r23RtJ+NQgPF3gG+BlJY4co8exhcpftcqHlmNVoIENw9pgzPxm9j8
CVpxrDjjmY9lA5ABScd6mbDYt84mgwJagMSmbwwk9fduRmbz0d0H9eugqox+Ih8B
D2CNYtSVqmalxkkTgaQlgcgsIvTsBUMK0zfzGBItMfwU2Uq4q3ph1Hi5HR2wJcrR
fb8/aPszqPHKJrTIdnwJKVO2A3RkrMXrLTel6ntiV3CvM4We/U9CAAp8xB7j50ln
e3V1GhDucZK7vMdpmjI5Q1ceu6Uxxd4Y5YXub18eQpVScqq0bDDqnUMFTihPoWND
AkhjueBNgg60TpFoGjmhn1lgg2WEOUo2WEIZJNyJ+/c=
`protect END_PROTECTED
