`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3yh5TrmEcoY6I58ft6S6zb6qyLHMw3d/AnZ7hyX5W6G9qumpp5R1Lajzy9vUIDT6
gbGZxqAbx2Z+hhANQPSLJY49aGZP6HunxLSV2EB6E/oMLPDUhbHm+iH6Bsz9gOfQ
wirn1PQt/Rrt9Fey71976n83XM+g9yoDDU91vtie4xCTP1Ii5QUlrxAYF1HWW1fH
oovmqVB38cTY/MOu/1C46DdMzrshc8PmCaZP1HiGCWiocEPQewgwUOXBuqcTY5/t
dGselsYYPz5oZtf/OZo7uksHDKOqnhUHAiilJGciyJgY0ZxT4fk3J07+IkEf9NFw
XBWA9+k+vX44PAisApuPN/LUBwyYG1ej8867OkfhmIuY+yVR7ffKcau5T9ehOXDo
mmA4AIhTaIR8JdeRdbj7bSiOWYVlQ9oqduGpY6bOEY9+Bdpu3GqpvMOoWyiCoFGf
74IIvU4G1Nh2HD1B04v/CkusMv3Wlgp5Sz/iDcRzUVy7F5q2WD6Ml3snssY1MnZE
mi7/kIlXmabUsjuIH8w5rLaVq0GYlYVYzSCQ5895Ttg0oeBg7yKMwlXMAxjvaq5K
kvoxtXDwagt1EyGcMFyFJ7p04B7GfGo9yyp7L8D2ELNUthrDoJRfMyFNHY4tx3g+
5egfnKa+5fNw1kzmdBGOM92mgRe+3zcpRvBYfOFYX+Zz3bgP6PeTtgpYo5CQKNhW
41pNdAv2hq0fbiNcbUYgd1U8RKcbIIkWOHAvA6zrkg79KidPS5rHKABi+YdpEqMW
qsLLzqFUhWXbzgXgBqpgIX+7xvMWJk4rVYgpMQrpumcUtoWkQxVR8NbP7O1KvXhQ
1LzaXkshWO4JXaA8dRZaijd75xqgTSlKGGV3hSf1N7zP0XejfBzYV35Vs5dRQH/6
SMSvqm5eUhiTbelrb8JCz0PRpw7tkfPFVzLSH1MoZMplGJCF4AzOBPNUxKRbYW0p
KlM6OPyeKb/I0gbPG1wuWA1Hq1SZX993Pt5cOwGsa8aZ2eOgB+uKy/rYNK53gcPh
+NqqSZ696XG7MdwT+3Wql/IVUhiTv2wZFLRhLytt0lbdWYsUjl+LNISnMHed0TsR
yH90TVSrgq/ZQOKB3yoY4LlfvxjHLKI2U6ma567ZmNXPWAnW7kV9kG9Jj87HT9kl
HO+t8Iou6Y5j5TBxHmClEKhsKPl8xeymUmMKmiQIKB1b5GRjzBCDMqBQP3iAr3k1
aJrTiDb9OE6tSTGHPmBF5DUdjmXyXNKLhcv6bLnvnSVsK2Wsp683Ii1guJFcF4H3
RNMvMUU85HA0631H3gebD798HiVz+PBtnVFuoMr9o7Iiluv6nILxXQeKtSOvhBpR
paN1NySYgAoPf3gvy59FIRvqdca+9v6CzqEFzRebaeQAW/g7BrF+bqRiTweIiIvW
u4pK865nK/V3pey1BSWAcsCym0VLm/5adXchcXXog1zCwD6p8sYvNLmoZliN6IPX
deUImq5S8HROs5HBARszN+sNvmoThb1cDcHNsokVFdjfC3n4Rz365wa5tu7BD8Xf
c9t+BR6K2tGVL4TmXgA7gJyUB9Nadp8QNsdwxSJDbC9IwbFfvoppCgd0v9teXq/g
TPBcdD2ph7yQDdLV+loGombjqLitMZOsE55aXEGZ7ihFdjtnAYPb1nNU0nFxEsKW
kV1GwvhKQP7YcAKW4nHGccJiduikwbBC9mRzjiuKSfXsUqf/Ml/hfDbfZmkoUM4n
DCpOA/WacHkkH+GvdrOmNiVdz1eMRpPMld+UxpIHkx8m0dSWjTkYAXY/DAL2EPEe
xXvvd3xhXXH/vXL4WAp7Rxz4GgOiDqP61bcqSSgz8yeP+QzI/nCJ/a4L1rhm0+oX
kLlxrLub5yvhAJ5kQiHbC45lhv6GbtCnHer8qKRr0Ksz/CfLlzig1x54UvNsJklL
G0GlYuqgjvpeDmDdSaM0iYOyWMRWraKmFBsIm2x9ihCt2ngYwpgZDEjl8LbrrhFd
3TOQ9GVyPozn+Mf6P8oAVn7TY2V+y3MHSDhoEW4BQpujyMCUkLb9SYm163KwGkOD
KWoSN6HEtVybCv4wqMpPLdYSq3Nyya8r+kURsw/oMFuREBNF955BqoiVB/9BH0Bz
MHOzObVw7FddEYSLKiZnEoXnOZmDV8+tPKuzUyTl0plTsGDwGebcMTFBqe0xVKCx
dqNvGNIP5IFnvifz1C+nNZVRiKfbZZpeduiQZbKDrAiTTeGt4lPfpfHSteORX4vb
HKMokkRrVS/oJTQIOTRlya2ZXQWiSW5Qz6TmiMGmUynUsEQYzMXEeS+7nPEsXgIW
mnu+4XFGoHu2WEOvvqKaM+q4H/sqTUnQAMQ9UB4odz5gf0fk6Q76cARwrvaU99yE
gfg4qS6EBpADgygVw35N6t7B8uOF9ELAD5aIdfx5Q0EQ3fN7hL8ZzZybZ/kF988K
9oXejrNR/g5Vmd/bfmmydjTBVEuI3cl7JKNU43SdHOCblUJ/UL1+9X35xxO/sWmw
3P+ams2g/ezQiFPT7H6Igti6IhrM9B5WOCEZQxpSVlNyPHjrc0YTaNrRlyM9LxcD
yUYEUiqztWo7AgtKZpDQxQkbqdXaRyxh40uowBVV5xgqrxhYXpNw49xkg8jQ0WiG
KkXJ8uDr0Us4vA7f//RQeUDw2kmYgev8MAyW4i6pFiWXjLUtMbljsChS80W72Tsk
P0l7Evd09Rqro+ZxmV84C4qmEsKbq+TL8HC2ekemhcPGO3e6ebfJvLgN60i97ns0
X0HtqcxGiO6URafMmErWuQQoHPywoxagMCdzZ1AqqbeB3wbS/+DjgZmhbqnK/GC5
eSCIZfRKISGW7IHyF8hVv+HAakE99VkC3owQSvHrTlcCSVpfgv0/S6Sr2w4wNzvj
/h2gymvXJMfS93vg3566iIz3RJ5izsKmrr4QrZPH+KlsAV/kiWSqGr5vx4cTbqvB
PI05HOaaclLAyj0VxpZ+PGbtHYH/iSq113q2wkF3LWjpGxzG+e0glrAIPVtgon2b
iTxGPEheDUH/+ex5GCZhfjbTdKGCP1uqmyGqLg+OfsjPw1KzrJNa0Uhg/a+G+uQc
3cCNjKifR9PIrBrBCS19zNXGh0elOXUZeoMn0HWlZToqlasWPeW8gilLw301y1Uo
/urJZwdNucObxotmOZB0pTU4N5igwXm5IDo7oLpHK/KjXRtujxaFh2KgptvDhJ5z
LAnFYdva0HrRLd/ogUR7N/Chd8t3ukXJDuHhlviEhT+c3Y9tYHFc5Zl6avgTDYOq
Y50Zpy4OQ0JmIRO7jF+7uLeNAZzjKzOc3/k8vLuoubAu5VfQf3j7TDqHcXAYHAaf
Evvwnu4o641PALdz7PkXDaxuElknnoD1KvkUsEyoTd9YYb7VrsJMQJXX3LXoaA6o
Mspw1P6QT8cV0OvseBYgJskFj6T/elL8BgAuQr++0decRzNRicCWz8flIGKyu9TG
90W7zqK1kCsMbCEVHyCDzI5H0JuH1aSCP+yQ1QmMfgnGeFnU7OiT3+rJI992QrtK
QXvoAwwrTkUVZaFvrZNLDl+hzkAJmWQ1BLJbSjAdQiQOl2HnuuEce1jLk8nm2EV2
Wj0tUlHhnE9ENtBRKeSMV9/sHBoxhn2qGaQicnlftJao7YhUBTZ7l8QczI3wfFop
bIFc2ZVmda45g/65Wb1Vnw5D5nRo4Z6YDoCq8+ZtCGK6InwWTerBmD7vn6SZ6lqp
7Gg7qHovUhyOJrp0N/9nfjC5+O7tMUJ548btwq9TaOLPe3l5uSV97FWsRP/WGu73
yButs343q+SKp6/sgCsOw4YftozFXXdRfRHE/sPuNvK8/ie1e7TSwlNonPZZvsWr
Kb3L7g7Z28mwL8GXJBGdw+wRZiMmOkPZY0CAAbk1A17VwxzATLwtrtuv+A0g09Xv
3SoSfwqrtV4j+UuXuz51matbDmUFK3005vJ4dywTzC0spvHe/4wAI7zTQGQnUYlB
t9bID3A06uza8f3VUfHqFX3r+vgWXb7KXV4cUiy6VZuNW15sJhJMXYNIf3tgcrQk
SwU/qovUjmQlIsHlE6RTCVdiiuUMAD6kMNqJ3zKSUl3jmTUYmmzgU0jzTNrVl/X+
y+jPP/z3vCAIzwrGD4J61WyWYytS5L7yWY9rRyVqoM2HmsfL2e+tQjshSHctU90h
H0TgKeFU1AGiKD0ubYzDLgVc3fdMqDbHmdBiiMGtuqU538Tp/T8jDZS0iNuqq70s
xqzIdm+qzy31bvtcy5fI3hbZboIUyq0t7s2QG84XlM1FUQSb5Zex3lWoKdQAPCeQ
gXpYdAhnZO5fEzcLDu0TOsg+sf/cTBW/ZfFBAcCJRjyznxc+UtJLZVqErsIXnv8l
lILAGLy2rqvqkH5euI7JVI/ChJS2qrYB/Ep4FY5UPtP2Zc2xI+zunZL72V8apG5B
5s7NiOswDcJwXwlw1Km6rx4tNzrVgI9tn6MC9LRf5OjUGn988ed8RPyTgFBJdsT/
t/zd8hRtIRUyV2IXgQM/0tF/x96aIdIyMmVbiYwJLqAJzX70dAKek8kbVpe+I7A/
2qG3GRgqbLae8Y3Rn7BZpvX+ol2usaPxorpPF6FYyaxkdOyi/iM198jtpTmEls9n
vlOw+zH8VPmoXolTrlecrs1muTeQ6XsFRU3nV0ZQZoeEl3T23gdriq4dTmHuLU24
EtzDsU4D719JVBdaVlKNwPgR0R0vhu6iU3Asr7GwHu0pBGodcWhLqiZbRXsLWJKo
N/Ionc8XLPgv4eYNk4JMzvBN5ZPF2wmL0IIzIAIk+vD5dCo5uV73FdXGBFtcDSc7
qU0RBYGYDO8eI63g64ASnQrbjrxoy3vutmVWBUZGqpjVJJSaRw31vLAreS02rpNU
gja2Qxj3Es/kbSUnYA9NDwxfGGVxowRiEkIcxHHjVW1anfC4rU4V5GyxF+hBB9Gj
8JcV0mXr9lDrwjGdPa14SI/sCALTsTNPnlzcmcujaLwUu6Z3wEDuc40IBIpzpXjm
JgEGYSbCF0VIFwG4Lc8teRfH/gjh9BSAdvqArbSffU7lE/LO7EWi6z0tjsrEl1th
hoEhMsRzb8lSCizQoievxbxxUIB9EIF24TH7IcYP5Mw32mbRJz/x/KI9GHOASVWO
+BfuwH06H4uK5C8N6/OxP6DDqazdrqtJQMzQK9NQTGyEzlomACT43hodeILwlCEC
27BAozCPw2I5CGWUKFU460JT4YnojP7Eew41+SGF4M0wzyhdgdVK0If1ACmWYGhz
yNLtc4Kr9OFQK0XouANqZ73rLJJzIetWccsroQ/Gm/MC0yp97O+ksqH2ChW1zNJ4
Wsbmbja7SwXW9rhdmUxlYrtj42BWvaI6l9v1VDSTnIrhBXpkYwlw4gm4uNRZGHYX
6qGP3dtqb/yrt91+SztIRg+lSd4Sb7+r/0WDwpiuIwM3wEhOsiLLGX/78mIMZntS
+tBUmmEEi5brQr8TITF5gmPaTtnIq2dW27itQ2kTrtDPhShZYnW1pH0cuxwlhA0C
HBfsxaDFpuJUvx28L7cZfsx9DnC8hwAB5DIuklAjCl6O8r4ER0yPc/kY4LOcU/n2
BKgl95aDGqXQPLjdx3LYeKsf0wfNg+mKRS/v0Q0U+gOvd3CZOJzC2NjjaU+IFEHY
MzKvLmkCw4A9KCV5Bjh9H0zPhSDtSUd06pabGrKwzZbV6gw1791BRggN7gfVIWIV
I6MwCdfaiZ0nzeBaigGLSbISvx+bt7G9BGlEwlfadb7BIdlKre7mRCiACdWlbtiL
rQxHjOw9ix6aYezGwCKbvn/b2UbcmUjUUfowpzNgAoClHtviCta5Wf6W2fGVophU
CDgmV+IpjwtLt66vGKWr6xCH6q6g5Xkwm4ldBFbAS9e3U5DTLFo8N7pM0XdcvAI3
B/u24UprQP42aUE0e4hUeqXbNb41Hk6qTXd3Z6RIUTN20dPTf0ZnpmOItqH3/8j8
+f/0kLFEFNSebLgHiDAwfrzE4gctSluK+EKdENjE6TDBuVZ1xXN9amKjT7UYFShj
Hgu0G0hXqTSh/Bl45A+keSlQevE+kcXeSPboHqIqQOmfT0FwAr5UQTlcma20anS2
OgL0Ny0pF0wMrd3QxaQDwcCkkKPFOznmldcs+TZzM5ULgjTwr/PNAE3ei0X4t+/2
hkfVCA9wCWLOGegiiWGhBEcooYok9rNE1FVC4IaNzZjOTqv3U3yc6lg/y2J07B5h
wqBQBzM/KrTebSmbSutp4fv/IrTbSARVy+CUoT3fRWWChTD0X1YsaifiTiazFvx0
KfeZNootfVosPoFwSlc8xyLmmJmqn2d/RukTuvh+VoAfSBqbBiCFPysmwqCVwG/a
utL+Y08BWvpRI32tshCJQs7ZqgszKW9DKJBsgIIG5d64LLPCQfS/F9OpuEwx2BcW
EGerr39UvnG+KbFqJiUIXR8aqK3xVjveGpdmCMWKbmIXZNmsZnNFzGO8A1jMLAPv
PHGlmIbtzk6p5xYTVhnl37Ey+5CCveG781oOcKyHfAxjikdlG4jR+2KHAQwyxcez
j41hsIhjBWpLdCxSEbrGSNLP/qeKTyPqKTM8ZYMC7hcqRSrZGL4sHinvR2HHyjCs
rlmtCcQXLqBmx04OemR8gcHEwNEVNDbnLKrsy0Z9ffIgphOCLAFkCfAZcnYu0+S3
zigh5AEB0Qoy+nIqMUOldcDpp15kp4y7dd+O8vw9OjdBco9hIsfAoAiKH2gmJcoT
WZbMqH4RmgBmXrW81EUX6rALt44a0rOGxzj7szQ+v8WAG4d98AjpyU/mjw7LH9JD
F0i0qXtoxeEGzsfG73JCYBiz+HxGMJH5ZiXywsb9/S9HO6eo1dvRJ3r+ybZxMxiW
aTJlk0E7u1w2K619pq54RugIvm913F5ZtgbsmRYU/LYNuyYdd0PV+iC9zMmSPny8
Z1vpN4IJU/XlwzHun33M6QQ5tuM7xdSTBKc4diwU4MVIlvdBUsEr1paBGwcUJidt
j7Q492Mcav/he88yC0rxDdqhVvEeRhb58qhhAdd/yu160M+xc9VHdLmu7YCBT1jJ
xLlgw9tTk9FNJei1Cy1Fmi+I+qrD/9OEqcFZPRWGF3NflgIxGSqq3NYr3M6RXmYw
wI0hx9gajomrboBFAapSL6U2leJNgjx7wrPCjHedy9svmF5GrTg0V63h+gHJjO5F
S6wDr3wsh6I4U4Lt4iM0NbIhv12BUsv8S10ckrv7ZoI7jAAv3YXkvkjiDMgFfA8n
XupH1NSnNEvHTLvFvpsDZnEEaVisNr0w6yi9dQjQnC0+7NUavZH9pn29oSDdFe0A
LUv6/q/kM25cI5EHPQBDYv1kCPrVl1s2A2QANmOY0Vv2GKoXDNhYpiwUEMyOr9Fd
lAVNx3K13R4S3t+eD9LDDcyyiACl+TyTURSOefQP+vgKN2UfQmN1fqGOSreIPd+M
H5UF1LgmubiZYIbRda2K9Ap5KrUUbj9h3P9JSmducZjlHT9NW+5CnSdFBRbFKbUw
aziFAl9kD8efDdcUq9YfZlHjWOevJZ6JGdbi5FvdYQHm/WGDbyj8kpl2B4S19I79
Q3lIke1KyJUH8vUDtZU6n96Ur6Jo6pDXRcnmdEvhokUx3Vsv4cso37ozuhFD0eT6
gG9obugs42FcHV+USNDxxtKSYHoGb7Xe5I9MFURY1wTD7D/PWYUHkDDaBaC/TDiM
KHKUVOfeKuhXDAR7B47nwgGXcXst59+cTl/oNXtRvXjB+O5xx0tR6ScqY3hxDDZn
BB2fqjlPHGJIPfqqA/rL4RBORAolQaZC4QyNaqYJ42WK2CeVeTVakGo/aH8r3Oj+
sQ2Z84/bRHX3rugEUY09Uga6uCUZnjFWqV13zviHOOMT8LldXgjK7QHapJoTAYfx
lIcSIPvrwGgKsomfTFyRjSxDpS6qHus5B+6Lu5b5ICf5Rh9yaZImzGgvJNkedw13
PZ905bCFHr5CWwHDNLq1JyifqJ3eKR7tCDYy4XCcBeVUkMyzKqdq8Xgs/Iv+o1Rx
TNbHcFEGhx97BMCg+xkYngsImDe1uO3UXutqf7zhGaIe0FNaYEmehXCY8A0HuQzh
qJKSuGC59TDTv4TuqrI9sUN/tooRKOM/VAEaihaG5nbLziIZIVYCVIxxsk0hooTb
/BaqK1kXPdmft9VxbTFjdDE1CvvGuWVpj0MU7UEGPIG9hPDWOn48+NjQGCgW2ncF
CK+VAtQLN1WX5frR4SccNnEaA0L6tZGAdZRdAtXAnOs9KyUO3H9RRzqqy4AJmKO1
Q9ABbuxonqAqUGBpe0bIDM5u7hoCiKxpWiG6wlQ9vbEDUHR0kyNtFyoKs9woauqa
NYhVDCOuWP9zYn3wp6B9nfP/o/6n6gwYWxaXriVxsIpCKQHeV2NAtuayPV9PxeZH
amtwMqor6VhYT06CyG/V+GnfoWOO1ZYCrXQG+q1Xhjl8ik3SrcFx6oM2xWirzENL
WMZNHyI+7yI5y54rpMvGtSL5256SPXRZHgj339hjLKMRls+ONj/fc6W28moTTh+h
rB9dHxwaJawaQ21yTPP8PMxZJp3jLm4BEE/0+rK0uQMse0MslVgNCadAeL0M+rBU
4nxcsYpjQ8/sHLEiCGBsW7E+ihSF/0/sbPwbCg0iwnlmn93XApii6hT4kfNMPKb/
qZyOggR4/2mitKcYUz9zVsf2jsmVrWVj5QF5414gGbx3QpWpejEdJxoM69/JqmUO
SN+W7GMT4HKlPI6YQooM9180mU2PcD6LFnrR3qa81MVNUmjpuU21t2tI3mP8zK1M
zfNr8EEFQYfXV8ODGy5088kaz4/xuM/trTb42PU/qK9Kkupd/gOBeSZWiGhebsyt
sdp/mYtEyvBt4jdvYnFgaK/r6/E3BhaEF7t2nAMUAeWpV5WHiUkTaE6fyhPok3zc
cPB/9/jJGWcB3LLL8ft1sSVyJfm5GeHPdelHKqUK+/pForsHUpTO4XlB4xGzPuAZ
y0aiZ4OEXkPU7OPzC0SuiGuhcECZtnTl/5rAs4IB5OnFdkOelKuyLaMxnWzStuOU
lhdFUE9IHr39wdOCxz4k+wEHLvD30QK7tEPeEJd3kL4SNK12iOKl19QRxwNVXawb
dXFC/NVrrLP22j/nwpJtAcOXTNQOQcj6qK3CvLI00WJTJOh43EsgRjB35+zZAkIm
EwtKW30KtFicLvEqrcbAWikBZ2Lxsv++dRS1WYpX0WJOgAPTk7x/T7534qYn3ruz
bIg9+kOCHm685yAOQxkQOssq7LIvlzE+izDvlZRfBQp/wwo+U4FZoPPAci+CH93s
xanMzz0l8bBkL4UXSIn5RGKW7Pzt5knUjKGe88HNHqR9it/CP8d1u5hjCdwZ9Omi
NuQ1JqKuUntcex9b+HjmM0a3yLMepAPiOjAEemk/gLWVBmIB2oXepVkQBTuKQR4G
WJUk9p30csSmzuiLASCdLkjQz0TSmU9YO7RRsfnDm/nJ0QZH1XSvUSCF92EA79sN
avqo50nBqm2YQZO57wYfI7eaJ5zrO4VJqV45lWaBoY3eTe1NmBhTa+hHNdttd67P
T9xsvFTF3wD8RJ4jRfVisqVOXei06rRe1c0n7UYr0eVJBnUS7Yhs9LBlrN/pdCiq
em67xpV5kTU8VUcH4Wk7mpEXusHxv5u1L1M2Zfx5F1KbEdH+dFD3XTd2R4BdfW2+
TGAd5Z/Cu/r4AO6Kw4qaG6evsc/LkDP/IDTwcBKHsHPnYVJd0SwOqApF0OPYdxOc
7WwJLh+vtQ3s4lAy/p0Mw8kMvhHeRSbHTIJENEP+wvF5gWaqKl7TZ6HD9/NU6xKF
l+DcUVjF3Z/Xht/yw2yTpR0dFVTvL1jtwwVXe9ILQ8Qjabcakj94h3p5YkfKoaBV
OMOnJcAlTF+udu1vcF/LKlUonDkcJOAq0F6YPdOIS+9r+PalGICUfWX7svxc53TI
FE3HQTO9ZOiR8PsKho3by23oo4BP+9XESlnlWNmBegfkLY9o1HZ9xBvAn+dGpY13
fXDanlYahgse7kaMjq7AfAHVLurcaNyhmLv1G9f/Cj4uHVJ3sjLzKm0JFL8RoW9b
Jnhc5nWGkfHI3vv26F3E3kcaD2xfGjFPotlb+zQSaHlK6I5x7e+OYtftwQJ5U47g
tjQgU9yS+fr9uCOIgJcFlivCAzMfUXRAfSYyuzxnLE/ffBYyOTEmZFmUjKnCuXIN
Q+c4TlonmQ3w/JmnwIJ5MDnG5dzL1C63p4+AsdFjq5im9i3KTolGe61fwzX7BoSZ
sj66BDE3Abgp2evKG0vY/Bxw0A2zmF3nQCuidEYIQz6VoK4+W6PGmdig1T1s9B53
FKl3R70a2CA8oBBOdLQZPgZj0aMyJFxFz2o+EPgVWbeu3QbI2zO7bowNrtIZFFFX
RsAvbMzVl4iwu6PafSg7daNvaF+ImlvmI0QHdregmVq9hSvVomaz0IPi/IQufyMk
d9hC+1nEPmDbfRBh5NuIn7z5CDW6y/bvv4Tgg+MiMmd6z1WXkCYBSgBUu8Mvyz2w
EZHrnFUjgTtU9kxysjYmk5gzwnSospfGaeQE91EUggiyp3QJK6WCDeojX4ads+tB
ON7BjCvt3ivc3YxyzjlOew==
`protect END_PROTECTED
