`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zpcznaKhy25BW4Fhh8MLvts2013lNEBaCPtb4QEAqM44lUo7IQj2T993kAhb8Hv0
/Ll0z3OWDsdCgPiAevxNzOFWf4aKJk/Bd9G1GwaaHrmKY+fUrjIVTHN1PLSJVXd1
8XThnGmB+oxLPXBvmlHJopRtolhyJXo4BQaJurIRld52iyfWlXBG8Hzc0Q7PjKsH
I/XsXo+Zn1YdBc8r8ZKdm7S/7TEVXAtC8XKqUlbSFkDvPefnvubdtVxpvx0RvsJN
wulXjktAWFZRywped585YMgKYbNMvpp1dZmntUxj16LFQ3+7vqRpV3ewnKvucq+j
MRDLng7IP/b+e54dL1RwZwXEJXvci1ggSG/UCRalI6gP6E78pkJ8qHbFzuufDBVJ
9NeyjKcmya6wnG1d8RLHLV0jQVM0RQGXUXzBixqf53pJuLIu+0xgmPUldDYEXoqj
Vd3MkvsxfDjAK+v02o0YQxY04e35FlVaZcIJpyBj4LXT9gVYrwOsFwspFkqT60O+
eeadz0CNvkMc7uQHbBop1XMzviyYQHjWHkbKY0bYrt5+HHKqVX0TsE1HDq8RejKZ
FN5e31jqErBiRwjDknkdikXT987lFKlUkwbXr/JXHs/sX+zNV8g+gcZo4wVVIo8C
aEUl/5yupgb0+IOm7ypmDatxINdQk4nVY5990WDCIOCXMpNuaELEwWBiGGHqLDpI
xZtVvF2/1qw5XXjFnurY0GwAB/WTZWCT/0GQTBGQ/vMUHlxYSYVjlJt8NVGPsZAA
PBAN6ZkbowjmnxhjGFENjyiFZj6oNHd7IR0RIGWl3t7ZI3GFvVpVzeDfwfy/qk9w
hkYNqc9ot+llNSv4PXtxGr4iiKiHjrO9+GZRXoRCslh2RqSHwZkin9Lhf3NC8rlz
zcGbXsKLWaNKpKlJjIYCpDEuTpUxpRbNqA4tpfqQw3nYs0ks9Y6mwRkbSKDVyjkI
o59twO/ug76aVNrhLoXWxBDFt6HjA8XSGVzsCYRU+rWf/kgRYCafuZqHKtWfsani
vz4fzkpz7IE74afEWbZ5pGOJFUEw0PA3zIARCbmhgHMHT0Uq2iwGjPX74mbPtWBx
c2Au3IZ4gURE9mW9crcEnPrsPfLR9yZr6K/XLqCjRcZbSlUKO2JqtbpwVzpcEiLm
f5sh1QyZv/rZOgyvrro9lzZzfZh0DBH4lB8UXZ26bQRiS1bI9jga0s/vx3uyAQaE
BdZ7y07wK09r0tzVFwK6qfCvflcdrSRW7NS9S+FCMVFRoqaJtKx8DvnmTqfutHQN
tV7z/HPyGMvl8ttjrfOfr5ITwxUcieeYPYxeJHTToOBgZGQDOWvGzyryir7t8Pv+
vroMuyIRDcDEsd4ADR0bwzE/tCwpCJQmEfWEbUVCgdtFAS2uO/mDuT94acyg8q8O
Y3ok3h5TTONdxtohaWDENgiWPeoqcNZQbPDCWJPoisIlLYjBpASGwb23nj4MhUet
wBT/KEHU9Vrg5yhj05YFFkVH5LnZiNvkRKsM/5oUL/GeHQ0dAeIArX4MlbN2Onr+
Wf929Uj5j7tUtQcCXEG4t6+BurVJyrIZku6ZuBLUsKaveGCmqY24onMUGSYbhICY
p3Io63GMTzG4podZDligYXg1NAIgYl67qUL2+XtoP/ulwAm+nU5+svpFOGctJhRB
16QQsHmXvTKE01yoab1clMexuvtztS6eoqKgzZ/bTX8kKKifNh3vHMDhX2idQHZn
+z2lVsizIMADZBpLaC6KhSx0LyPK9wPrAh6QwmvxoCiq4tDZ4GeLItcyPJNPk056
+CKnynf2bM0WsmCT8JUflwoK0XVN1B3viA2/YlajAPNYzusBQjquovrhQOOfO0PF
vWW/F6/GBM/845cF/k23HSHFIL2V1sSAYKqH9oMMJcDrnRLQGQ0rx9zTup1Bc6FX
x4GBEOShTo0L3rhNKXoIQFQKq01WhzaoCL1QvDku0LwufMl+YxrqFl3194AxD/Jo
7WZZYMIEs/pt/rxJ3HtD7jFw+sr3ZOxZYoTShph6AY5XiefUTeiB3qGGWRSlFluT
KTzj97yHiyldlKvR6rc1hsqZF1Y+o5tQR3Hx/IYYPodf4sB7J/6+qW5Tn2NKrmqx
xCF+6qGq9x4fDPflpUu4otukbbrZNhm6MQfQhEo+c8M0MWzzTXOl4/h4X3YbUPRK
+0i6TIA1Zy4fspmUEQIvnNkyhfpr3KjF7LAbsOmGtOsledd7B4Gsg6pIkRVO5RPW
YjoUhMHBlvc3xFCTrYvWOa4lIGDUGM2pwOC594zjnQHjAWKaAvM1WRB/Go8PXESv
KOg10cUo0imRyjkABQn/JYA9PYfY0oiMhL4wXeshraRNcWJ3XSJBVbk4MDGU4OE3
AE1TKsGsEEJ9JeaVeNQDNk3tptTWSTOeT02QvRkqAwdDPNcXtz/Gf5X+moz3hV+x
4PjNDKZ3OpBnhFr9x5N9PyNF7qRK9hxdzKnfftUloFHaH2HETMRJ9P4BaYfpZgAD
/OB3uMMmbT+tWF7uksyAGji4Kgr5iqdO6olinmmaNnZxnBg9IB+nSp4nv3gw08+Z
znLQU2mO5Qic0Oegy0ChPwFWtnQJkHVYY3DgmspQ+/v0j24WHQTu8c4N9VRX5ihk
a2fAxgP3798rgyEo6/e/K4SYUI6m1jIckloTmX5S/oRosauflk6pRbI5dauvktjL
1OP5hhX0UjiUGDwrr7CjOaKOBnpx9228Pptcv0bAZWQ01gZAxXKJIehJpzRBxhyW
F09hNFL6h6WuQCmZi6KskgrGX8CIOxiCuK88sMx4mAAY3ykeFElXBZGpUqc9RU8j
D9B9yAKahPF+21B21o01M9OrHTf5YEsccGQEUs/WGHnLFDqQLXjcEPPCDFIJXHiJ
rMYag5g0JCYzN8I2qsA4u19uW16Vm1YHNJy7BnHH6qzxFQTxXNM6P3lk3nhfFAfE
Ddr9fqYO6jKNXpT7PY2sPeSfzwRhtpq/BZO4yHrMuquBpypmq+0/1HO19KmS1fuB
l+a5TEyuJFFJqKUwS/xtWG4cew3fZCv/SFYTSGcO8qnB6pESq1/Bf0wxxwM11Q93
LrhGU5+c1EJJvZYQuaap+EBluWsKMDyhWLCimOgBLlORfx7xifqhei89mkkWP1u+
yBuVUBBCa+xAd1U8dkPD32xCgL27/vFypvYv1yJGtcGrIJsHzc6LqQ4WErY61pGC
khR6qEUM9iE33KLLeIWz0iDVbPiBsdktw1xKGL4LUe2pr6x4b7Qz/zS5F/+xo4xs
sWk3me120V8+S2VoGs67Q35dn9rj2XojlsOo9hF/suKPI2Yk1jcbpbwd1DuDF+vX
c8yB1Dbv2eFDsTvj3s+tIGEfjl3692l+5RVqFkFY8Y7Ea12bbhsGFAcA5Xl7TM+c
DCLWaCo3wrSHNoNIgIIyq9dHU1dmxuv6q6eIdzkgpdnmSv0tD1Md8xiMnJbHViPH
ZGvyZQh4Y1vdHx+eCl7w1ppMYr/Gghypo1qrV0o3txhJoTxnGQnUQWEF3cTzlkBR
BxIQDEJbFbI3hl3ph5d/LBrJmO64JTxYWLUUQpA8z53tjxOPD0nbHBCmJYI84c06
rMnueN6iZpHpAlBsTkk+OIFKP4ylXfjoS+l5eQQk25iysE62bH0BByw9K9SE5lsB
Uuc/E21IHam4OZ3nWonH9HplmUt+v1uds85AymZmD0Jk1oKnOvj5mEkDougAVMYR
NrdHSwb82B6wi+g9lydSMTuz54HX2MNO1toPTZ4Eu/6a6mQ8Jc5TimmqTnt33EZX
savdfF8dXG77e7C5tHL/48gnzJuLWrXcSMgZd0JC4GQ7Ydom3l3VXnjheRyJqvCT
RiZ90seq28wqdbWdLT6nLRb/4TGSNV0ku2YwruvI0DWn6SJRAzS5vJCoONEtUPuP
xmtLPjZwCQotu+pMUhK7Ded3BRwunztQf2rohIRaTsnz53mQ6fSqfPS1VphdJbJd
7gAzpwKILYcRzf6wuC4meCAIqZeg8jCGkn74LYoHauaSFSAnovzoOhRmHNa1lqJQ
NKG5YSmxF/cgQptu1tSTXFgNPHNYQPwb3qPauhSOp4LMByJGAQLqbpF++qevakG8
O5jnxuXKA4O5iyYwKEoxI8I3RC8kBZl29km7lwzjyn/ELd9WXExhi8NhivyMyExn
NIWTAiJ0ZeXIxZKoPXhTQoU2tu0+fkqSzu82jdZGO8BLv0w4XH1lgISsmM8IhTba
6DfW0H1bGTZ+MfaAdtg7tgEmhLArtvaYIncLBWqRMKw2ya8f9cIGhyr8eH72829K
Cq7JUgl2pt8YLopVoHm11+a0q6Kvo/7Vw+zeowGSQEbIusfK1x531JfD6wcF/3kM
L0HrvZn540puMzG87PAvmwIAf5N7E+DCLhqxgn96duZNqdggdmebXZyA8m+g8Z3b
JgtITy7NSJip+KOazGwIhbYDzuCqWeCBc87gNBogsxSbOhmdOr8S16XPyYmS/zOV
udWYTtbAonXc7Tms6abTVWM5ikyz3CA5pFj46qU/s6MOjSTgwc0MoCfvB+yTWsvn
1jl8gBbNdbh5G+fwj3OYDmhCkrhu8qHmdc/9sJahB+hSlB3zha/ttwOnAVpSnkLd
Kxtr/81t9cUfrNvpFozx57ei6+yMFXAKfHUj334mUeJX2zPsC+MtxhASyj+dIegg
MLfsxBnchOrXEVRqHTgDgOvU304q7Ff8tWiPMDVUc9m+Ncnbw7U9mTC9Ov0aEtHW
T+t03bhdemzwnxz+WNgPGstEcFv6BoZRgxkE3Dj7yhq/SSiIm+Eykxs/XGajr0o7
v3pgxUb4ssXs2/GgKvyxKE4sDzEpgBcHeWu26TLEZO8feiXQ6z+I3rD/bRShf4qj
snORzVIO8cgIlhrCJUs7Ni/ys3XjxIgLcRKz0nGiYbQZ32xVFCnw/Og0A6Czum7J
4lveNukRqggnjMdTewahOzez2h14AS6x+aVyBmIyinyVK8s4/ZpH4vZsjOk0CCu6
/0yj+TyoB5TG9Bu7AXtN82Mz/kL2BCOVFN+M6mZin5UF9XisRX0tUrWy8Jvk7g5O
4dZQd+j+Ej+1CbWy8+fXfw3il6lrv5Kq3+6qOU+PcVYrvTA4DS/jKBphXdcHh6f8
flnSmNiUBVL6FIGHIAkrVNnbeaWIZ26jw4GLqDYWN0MtPtyzVq8dUlN33kHzP+Ak
NsBJj49m4t67bVrFw3Cl+KaYLMabPud0a70sYNVNmLQ2FMT6vi9ItLJCtwW7x8R8
pVtLGTpbzGbZojm5KX9+08jS636kVPOIFkhnVfRmdOyTO7B3YaCrl5wohGpQuRtq
SAzUayJlZ4dWddoPhM3uyrSRoSTBE/9yeg19Wz7wka/JVXCVooM1ALRMv9f8EiRC
V18slInP9tSBOaQpRrIYmBLZE0WkeztOBtPQJcbmxCm68X8CBks3ZwsjyCVRXIek
9m5HVa1ubtFoADy7A3+IEwiXdK6Mx13vTtmIOhbjZeOG/vBSIJFqKMLyBnwEBBwn
atDcKF+5kFyI8fRcijsx8/vFxbUN4JTkOLcCJ4lFmMCeSFgr3vEfGgI8SOv4eheT
uNJoQDm25iG7gPyJhXDpFxp5YIiSZ1iJ+4fKhFRvfIyVjiF3nfHQfJyzWfV7UKtS
D3EDlHatdWI1RC/eAa/C7NuF4uZ/gfpS4pvM4y5kMshvm1GehSQ5l7fII21wM2JZ
C208LhmwGS3sMAt6pADOvk3dxo+w6XXA76s+I7V0WxNoMGx3Fl4n66D0U1ctV8aI
RxDc0hNCV0zQBSBwi4No5tfaj0JNvdWQGft+TI/Ckk1Y+zPr4VCrXb4Ndh8rQ6X2
MtmzRbpvtZMEFVW0XUTYpdPh9dtQbvNJYCkHxGHAazVbmunSSBlVh7bSWhPOaN3K
5XawhKaE6sS5MKLDhzknYqQiGy6EpratC5KywVk4kbdAuf2PHcvCB27xolA37LaQ
X2pwUKk8kw32+/dIWfjasoIMVIbIqWgq/zll7zr81BFwkvSyVtoxeZnlkL38AYJP
Y4l3eqhdJR3UkkXiTd9ZT5bXZIsUpWgqXG7du6xCqfnSxtjENM/uYCbIPNJOdwjn
05kHSBKHHEKGL+COKCqkwA6iv8aE8H8kwH23Hwemn8GkIWUnlup+GqFBeTOiPbPt
XNW5ty5L3c5gylYG+8Ee+k9fteXz7F68pDWMAVhY8hrmJquPU7HeEb5GMQoLg3tW
qFYaV4U7ingbGTSK7hKJYs0OdVPy3f70hi3nW4rkwgKhXwrdgfkXQlqtcUQGJiAh
6srqGX2VDOb6E+kLw7JhGUMSsLtBVgDPijDOn6y5wXllSWa9sSzy2zBDB4P3XDrr
Lk8oACaPvZoEz0YfS6Us8DzNmNHlK3xsUFMd6h/RinKPsF0obw6t8WxYqmAj7Sym
MbbVqdD7iYaw9iq+f8tDCTmQ900BuBwYRwPUG1VGhIKPFF0df59qWpeRP1wd/Id2
mDBT7DI4jmD9cMz2OT8IwjspDRl4BkwECdrgsFMzWvOUaTAoTw8BmfNt4txafNuH
n7zKn3iKqkKc9OwZKxF9R7sWqrt6+R0ZnGM8xFkZ7sEsAnH4GcCxWFAqGkpcUmjW
dDLRf9ku7P2L5GD9NrwCyKz7ihCHy9SvKIUHc/5oQqkiA3pysRPrLqwShBOtzGL9
mur8vpuCAseRUJsqJJvdELhfcoJ7JmXyGOlHOwAfXs4E+07kuL+JfXSvb3cCTF9W
9E5bsx6hhKaRXJdW6CL+fcF6xBhgb46GPpYzEu7gRymhEb9/ll74ZP2fXInPQ7cl
okNwb8R1uxbPcq4avtItzz/MwLdwVQf5M+2krfyH60FaUEIr3DNRMa2xDVFpvkDa
XguNmHzeT74L22J4pVRf/wDTudQFCpK7DE/0Z4aMMMB82AwIh11TJrsTUOLnpBYs
xbw1ex8LBeFlXSJNT8iaF6JqxVSFPdKVepCqJ8I70TcVl5DGFmDE+5CmqaRbkfGk
7+VNUQG6RbwtjHjE0PlplMs+rWuMKpIqbbc6Oi/fbMoUti0Rn9UYyGouYUcEasRm
D2ZdMDS4Lr9sQhRSsjuroEbMz4kNU0SUq3JLlFOkUDcPB0UgUKmomBxSB6beWfX5
LSHOoerG72elXTJpKI5xfTxdhRJUWJUWoJdmcTOg9fGSvLrDIOFls/IfiJMZFgNB
M/DyWCTDkBDa+wIh5OhHrnmqkr4vPwKjafL6tjh/IEiD7cBqMcrlN/JdZy5D1k2h
jM6s3G4BAc4sjv5LwAv0RUe1trowUtbYbdS8uSjdloyXb6CRA0unkIgRfsjpL+4V
v1pqoS54jE8/hCqLXsEuawtDjM8Q8Rio+y+sLHllq+9pko2j4LPGNCSXCA1vX/y4
NtLZs5PML0UoyWFlEMo3qeaHIIIo6MBQtPDGJ9NoDXUW0VCJ2qqAYUGTuIKM1YWH
nZH4mvtZDSSOajZ1++Qjaw0EVwLUfJW7mkeaXo0y2zAjg4To3h5ubY0C/yFhPVxq
6MuITlqYvgg6oUIwezcYPt2ktcheWqSDvJB0pftOrefpKddmqh7J5QCRcAH0yRh6
f2MddrlTlQWR4TqnVbJp2WSDL82JsKrEePE1bH+xmdEOGJ9jSd9/WwdhWkjqm/hc
ggpd5YSjNkA6EtgZ24LKNwnv1QdE+u34mVtoxl5ze8MHnEiKiDb15AEak6xYjhHm
3EGQDU1wmYhldRCNyqx+3mqb5Rml8lFqvDb7I1nk6EFaOB4qyDF1BKx4MUYcKqJt
4SnbTVaSAgAPLQb1JY9j8R02QP458Cs7qKUtBlVcfQlflA5Tssq+M0mooR7WzYkF
a9OmLMkMUvb2uB+Rz5ytn9+HxS/U/P7ulhaQ71RHsqBB6jv2uEDBrA9Zbjtc/0ls
wxmsqFJXPoLzbR2gDwRlx7HjwPXvHuFhPnbFdmB7zHB2OAbrAKbE3b/dHJ0/HHzn
H8Qmnd237NQ+70KnQHaQfz9LetK2SK7dnSgx5Bd5B13fIks7HEkGgHepHIzsfyy+
deg/R8BUEAJNCsD8117OQUxKsN1RFJZj5ZILh7ZvJ0RtdB9lGIJWB6VVaDFjkNb3
Yr4CW0P6j8CMK1MR5pYPWJcjw9EynGV9l/7KtNWe4BIsR+e2dm7vuH6KBZZPedVi
w/Xcgy0jEx+rZPU6DE4/PHP10ggk81hR2rVNyeoDg9PUDzFXT53g/qHHV5d/dw9v
+a4FhDeHRMKSNZTCQNrSGKaBD+yWfvSxcqSdxS8JN4CV6eH5pXa+3W4xj5qHEBEx
H892rXgOiOv3Jx54JibdLfNIedDCv/vR3iPccn33EipWy2qK1ZYIUlpVpdMBK32F
Gz+yukA9vrGqjH9wgdrMSj36K8oNeL2OrHywp4ZEDRRWFioT71qGCyTb6q+2HjEn
6Ran1sbHua+ADaJu+vr4n05ySbqT7uiFkkL38EqU0/78cZ7O/TC3Ij0/UO+CM89R
UZUrIH9PY7bY5bMoC3PCHB9g3/G1dwR6RMRwkGWvfRss2K71a44NUWWrIwYMUESx
04tRDYgIdVs3PUG0GPrLEbN/zaynGz0iy7bGhWvhs/aENFNtwSDD8YhqSiX6opiy
e5lYx2Kbzb0tKLddbpGgp6NXcqaiBt548KSakTH+i5u43mhKLjYmK6/z6F3mSUIS
FaRlKjKxsHS2+TPH4DUzca2Dp/TujdRHs1fILGcZJY8ax8UTL3fwwLB9te0Rdu4C
gmgjYKO+mST1G4WfsNYLGHVQk2bZSxPG3u66UMcoV6sZNyNPrYudjrDbNPd/zZoP
gduaewJKe+1hp20DVIDj7zmnomZjVBndoJMXdiCb/OwCNeducJ6p0mhsZj4COBT4
FGsh62gUZnrqcwyxhgyClJhh/Bw+no77Of1POu5tbunmEwHztJqJkqO66o7wjXM6
wkg4Z9LzVySV9IDSnW6OZ+HYf5GEqa8bYRgQIierFWcN7MFrwD6lGHLlpuOmNZvM
Vve1+k6AfZ6DYCVD+OgSkkmONc/5obnZyFEdWZmTkH6tiTWUw3vW2lp4MqmhJWBS
xZV/szs51jwjyI37N/Al3boYz1vJHNWCZ4yFB0NTqufjtAsDrNIhQz2NGlInF6oO
40Yhs3mSrGsv2JJc7rq9fMz245t9gN5PRRgGJ/dFG7l+5WKvC5wP3JklnMQ53fUJ
vK5O5LkRob4OA6KZ0yxTLqKgcK4aFIyhMlN6fWVpIlxLYqBAMNLXPlAXjAYcRYrk
CpBcq5tWtCWk/QHD84mQbpGiJO09SUUxUgk2OQ24SKGBb3xLowIalbwtJq8hEv8Z
I81eY3XNevyMjH2sYvj1ttO0sL4XX4TwiKH87K2qUj3peUSaxwWVpyzoptXZPDrH
vmxW+wdaclHKlNK8o/G2zKrnNS6H/oJtIiddq0MdEsILT0Y6DCvFNeP8zT1B+TQO
fPeHPqDHQolW/Js/bOS2d86TTZeJiOpuRMOVFoMxmx17m8C1UGA/OS7NHlho0uQ+
QxRg1ciFtftJGxQTKo8sHTXTlZiMikmIkDc4bk1ap1nbiyOaJhl7xmKrqKeRA19i
4zdiHmxEwsQpFDVjKAd4MkhFZIr4keylkeGwS7JKhUyfYwv/4iXykCa3btHFiB9f
DEXUROCJEl1MI/53zmfIcBA/qxxInzkCcpGC3vd6tYNEiftB6oVwUhFC5YPDLdKo
0JzhjsjnuoIHeYO1eqRV0He6tX0bhZilUBWGY3V2CcADX1wDNZUXwD0+wym4ZvfX
9HFYB9YFFqy9BRWAWhKwZL0MoSHBknCMv/nFwFZu86M/sqsfIWgvRKVUd4w77Zvn
7pPT9wnHFUw5mO6aV5o8G4d7CuBBnSe5RoO3viy+O5/LAhCkW97IRpgdJjgj4YCt
rz5ejrWSysN3IPhWJRqZq/f9eJngyiYzwvoFSYGcBe5lQ0SNDNA6qQ3RJAjGFK2S
HKOlyaF2eALFtd5d8t10cbMFHZlsQeN+855Ij0cJbggnrpLe4GcBWQQUymc9eyG8
0pOfbKfr96Z+geoqcjmmtb230182DppHVXg+KL+g2P0j4x9V3mC8rpADaTqCyl5f
tj+DEFgbFEmu8Ad2ZkIRw7QU11jnHORtMoBOG1Cf3x3bS1lHx+LTBXVIFCvYeZ6V
jIRadiEbYOpdS0StskCW8tTUzk9PKdrZl6Wwsw0bPlhJse+UA2whaN2eEDWedQZN
8SYL7Ro6ODoHRBOa7gjqhfg+SpWx9UI67mE3yISI42sajFKP0PMFM+5dgaGu0kNY
hR+4dCr7oEw809OL1Us6fyqwUL6domPcAqye7ErKimJ0xBcHpzikbEJKiMtndQz/
lNTb0lP/iPZxzPJ1YUk7QGvzhKXDs/tc1jakwn8jjkB557Pib7RjsqSQtGF7dXed
refcMFpq5rOW/uCmVKykTkKX9aHu4sN+9tr2owYZs24zI3FElmQUJ4DCYfOQHnHe
NPcsf1jxIv5QF+F8grpct5JR0/V+XJYfiVklR4ljbtNlSXQJwqmxF3QBIJH5jM3S
W8IQsUDHe5WiEfeLyEQjyyjv4ymm9OuYTcpaUbbaCrAcZ6fj7EixnVj/zZhS6wfj
bqxNeiU7AuzjJnYVFxfaEJFbW86rad2GnrCTeEiy5JM/r1vLgpV09mJy48rIJNYI
kH/9T43qBHRDZ9fuRzHusP69pu9tob57UiLzbDkUnVYnnQDyYpWrWY4FIDy52tO8
YsOzfEp3pjl/R6S7XwRfuUZ90uhBJPC+/rZt47MX+EgJC/l418RTenc1Z1xapguo
3kqiZsZJiqsktmNOk2WpUGt2srFPrH/zbMupDPDg9c8ds5JvV13Sqeso8Vff1PVf
cBK33eu3DgzpH+xbG7t1umh7JSQUrHjNDazP8WIpqbfVr1CSaI1PNFDLT8Xu5Vuj
ul3381QVonpW2AjSdzhJIrRRGnlIcXNYvy3/rECDNf/XVS6Qr0maAxL/cTPqLeUs
pz4AKjqjcFAnEWCQ/6NKMT070ZnEj69N8M26NvezON3Z4bpwSU5Deig805U2ayY+
WXl7ClHGUs5lGezB29ipwoA5BHojUQTsdr3M8suonsenGfugaBsQPxBtJi2uDKct
+8IXrbZigEV1ObPXHYm7Mlm31WHtT1XO9LYJTI0ifFzEfoDqAZ41yNddMiPnb1fe
jnJrAn+4PbkMEzQlvKsjB3x4i/C3eO0urMqSo7PDBsLciKYPfLfhc3hgR8dcTb+f
L2WHoUVUJuDqVJlX7kz2Y280I88FUOM/97QQ9aRiAbZsOVokHX24/t3EH/ijxUQt
V9LjXQ9ngWFUV35H4iQ4CQTd4TASMNMxV5wMJe6STTOI0nszNsV4hwysPadNY4pD
ZoCYl3tA8n5nuYWdqrlZFsCP8u+4svttAj342bp4WfZ+PUd870HPPJsB78C5bHmH
WazquRFQbME8QWo3YeT74q+wVzJ79Qn/ZVAvNAnN7QGW0Tk4Onysupy2mZVrVipO
09+Yu6u6PFO8ePrZkqVVvLbanU716VW2Bk3CA14WUhlAXkMT7CXuMl0JkBbUjnAx
PQnjhQNYV5fSzyu6iqNr8iIdSHx5TOa9jk3dC2WXlBNdopmkWIVdEunZ5vaQkCkG
zpjaTb08il9uXvShZ9IcpqDRXmYJLjB/cSbOMIY+sTacJNxwEc2wEWji0Lujuj58
D7ELkXawGx2GY42SOCD39SgxuJceU1acxX0haPjzCWMwVPpU6wSpVBPeky+f0dJz
Ky/Xfv4YJ5iGs6xSQa8c5khxnweAXYjKse3WeiiR4v4U9whyVVYob7uPN/Sf5yMe
B+J0Uli450fhgzhYtkPL2HVjDHN5kvXiTC7dIwwLrDC4Xr0VoFcRP7FCOpXcvVpi
SZ3l+FYej8ODMvoVHLyHH9MsqeKPKssH+tW2KMzYVqmoWLBkQTSXq0ErLL06wtM3
4u++GLwu/sOYV0CjX/Psscdgp+SfsP7K1+sFX4RTBQQA/mseMUm7m4UxdYTcC4io
6khw7fOROtjju0n7tuF/IhffQR5rkqQdm3kwHYsVDjEAe5o8Ocn1J+QH2tO/vIRS
cNVMHWlICiRYilEM7MIM/2ndvo+/hSKLO6XWEr54sfYY/mNAiBhp7Naf4yauzVRq
2ia94/QfQVh+8S7ZrIlTggxXso77287DLdO/WDqvv4ZFfvOV9FRX3t/V5GTcPKAX
PlHBd7i5jVNAsGYZ9ra/TAyiP0ofBdQpOX91d18Q0tGAmxECzxdPe65c+9MK1t6F
t+pIeigVDYZ2SBe2+baajsrsMpabMi5hcT2Qg+ixN2oPeNpf155Blh67XC3dgMvC
kc3Rf8p2L2nkfHFq110kBxqvEIUv84zInICE+Q0nu1mr/vK5GI/Gxyj1ckKaWV65
j9viXTw1Sep/+GUFqqV7LMLTnjfTwrH42QPg8iiCyyL2D542ke9M9Ckuqq2AAadi
t1CS3Sj8mAnQgdVQ1/nbOOqk2l0OyRrBEFyRuC+TAc9eKqmgqyGNdevii9G/GMX6
IjnASpAyNDyuyyFRgQYnX5Y/ssrhCz9Vo8eka74QkBanUb5n73+9J2SfJEgbG+2t
JrZ9TcJVTZbEj8T9dkK5EFQsMNYBGeobhUj6ZYWcAjXRkG6u0LgrzlmqUOiOzPFb
8mijquEMaZBHu+iRllz4gRNlNO13QAPCTlUZ4jIXSavrJ0C1xYArQQJjWY9Wn+jC
rlGdwHwux0PacPXD9DnA8T9STZVL5BRmGnXiplz/jY1Bw4iLTLgqRepWIZjiljNS
VHsOJcaHZZhrpQBo9+3Q2JeRE+aq8wt/zHYlB3+tP1P3k8cBJ8WF9b3FL3LIUnmF
bdWaKVvvRtC6R6koXcdfwlsldmS7vIHoYcda4Lc6qEi+JZKTSgaOEYdzGC3l2AtV
+2brdgh2pMxVth4FW+LA/mEmtfBv8VCB7gIJTpKbwxmzWflVI85RerDx94Vdn4cq
qx+/LsX4iXqO1JPHbjtNBYcZhmvbOrZX9hG0Ki4zJX98feNBUrr4jXDshqS0ywxL
7dkqMO+fY4kb0E4fRKL382TL6yPKTzRxsy/zzUEFqHPQcfY/wfFIKJ9GznHLGITC
SSeqzcnJdOPlWtSGBkNj3ugn3wY5jJ1mh0fuZYeyBklgz6ibcEPy8BuwWXKpV0pp
FqF9lBGobFRu6I0RmH+Wqc4f8qAIPCGP2M2z1rtm/H7yR+6/CFO9CBTa0qu2p+1P
SPnB7jswRkcERwGVc+XP776NuyXnqvRv/gy9VPQz7CfALHqhiBX8tAiC55qWQ3+k
fzKXNXodUMHA1XkXsIY6JcZjIHvnpx9JF+B4MGhjMcwi67ni+l/NW1Ue/+4ToEx0
cSXs0P6/n73FT4DHpKW81c+b8BYY0U81TLoHZTGEpu5froXaCC60KJl4hCQPZqre
VfehXCurCw69Qb4HzI+w24t8Cn9W93FPUqIm6MJGYDhlGOrbo7Fe+mBfoJdnnLdu
wYYguib1z4xD1xKd2DrKSAmcV4mlEbW1A/35LGs2nv/MWCGrdOP5olkaKA+YItDI
dRpIQfdRSTdxmL/xakHWJ+PYM2wLL396mHHHteAeFg05liB2/jtbGXYbbuFVlcjY
mXf/nfkzQXGqttdE3b+6DUNlvE1Ry55atac/qT9PkiHiyeRKze2Qa7NBhHT3P7p4
jd0SENEkLOLbG8TPzanB2g7DkRVZ69IpuBr0uf0YuaZjLNEpyCNIhMeY0QLLdkVP
96ofNDS+lc49bKjqP6K9zBWmUuhfkfEsmfS/E4bV21c3y+894wg6+IbfLrFHNxLQ
TB+SYjYVOQxNH3L7SXyuRLtHWWQSyDMoQ6uUrc/pN7mWCLjQFfoP0p1s6JvEk06/
CEYfpi6b8MBB4hwYoL6WSqEAZjM0DKr63TywqX+xoR8qJYP03VOG1nIXZddb5wdd
GKYF2MIW0H4PLfYQyoM5s3OYJmHroesJFwC21YODEncCrJbBrQcaK7tcSSsjn8Iw
TvQjEBmtnL6M/EhdLO7nbtf75ak6YRltwOqrn8Da25UqJQUh0+Npu8wFwDlVvvaJ
iPIiMQPuaa2WoACN4WM5C6zrlLgnl478xMQBlGi3PtszspgqyxC+m/A033lM4sVr
/mRw9MxHqmPYNx5LAkbv8a9tPJbbwVB2RWLnmSXrHDWVfqdpJV6EEZKobV8IcNJs
aOuHn5ordoJBCzr9J5m1FyNPbNvNGDpQj3n3OeU7pMwSiAXfj8g1d7qviXiMR5KG
mr3C7P2Kw2ffgyaLy7NUuo/KhKLcajojnNNz3BeyzY3gc1uRiDnjGQ8iKAZD/83h
mMuOwpc7SEZjaBZI4hoYZq3k3LVLFjM5Wppn9O5a9bYj3U6jIKjcTc9vU7vf+5mW
cOqKMC2CdQCFU1cl1vJqLOdinJLuTeeqN2jd1P/zlaIRk5yIHxLeeGPM/uCnVpaB
1o4AeYvJOT1vm7bE7tZAHnxHff1WVwVajMMk99ypyD0HtoFX8mz3wOXAyZ2jN5Wr
lk3f+EaHbIICUyZOQkr0JdnUUqaY0nybXw92iuIEMfCoS+dstcEEVMscHpDY55/e
NqPOsaRmD4XNH4NEsVarHP1tfkGZp+0ggp3K1vZSaJHipV03tXvP7Gw2r+S6TE7D
w8I6OCyGUrAheri5XPPf2du3js4Dk2KAyqpifZpJNBYUTrz0ig2BQtqh5PU5qcoT
jJ1Y4cc/Duy9UZOS0nQ4+WwcOogl28ZQXIPepx+cx17icWx1pk9O0wxT0cEq4epY
NMHjBOhfY/MMdNm49cTPH3BKC+ZGseY/W1mm/jb3IVbWqXFE1NyB64yA9kOJDzYL
Wal3kXTZ4ZX0284zlfQJnp/hTjxtz2/ZsHXgalbm9vmZ/FC6o4gP+nXP+yJEtCCX
uBqQIjC6qW9iv4NbnFIBOS/Vj5Gaiw5nlnQDpNrdJXXCGn1gvg/Iy2cXB/XpKKBp
zPxtAjU07SEhTPsXRi0niOaY48V/uO7NFOB2SuI06wSy++ysc+vNNPSaThtlo4v8
J8MAFwzLZhrM95Fe/MhUWwe5VScJuKKIYfSKlS36qXNvlDJEU2ydTeDdL+zhfxNE
zqvyNf1vVPlcmziqAyAys0C0kYVUURlPZ7xGa5ykjPsMxDal3kfCNYZxo2TYpvPh
oueBmVm1RvWq3YAaPsfOsA3iLifyI/ALDczPwkX3HCTMa8ThDP3/kP8FpZA51WCx
7ZjRxW2GuSML5rf+OtyfxVBPjQg1dGnGp4pY1PcWRInNSdYlmMRXC0rUElbuwsFY
Nk0a71HgGgiUkqsBIjJhjKbK5qtsmeatgwgaKhtJAYS8/YlX+0BscUrufyADcucK
Ku7OHpR9ou8NOiUY+iCmJ1CLNuCJEvFgD09mTBCyFOcqTL9CW+WunnEYQneRCPYs
vk3ZEAJr/uy2WNBDOAojcf/HhQXnF8Pnr6HZvEAy8I+t4iB7m9F8xhs1ZmmdALKl
n/INCK9a6j/OU2gqVr7ngbgjt2Bp7ZUVnrMWXUBxfT7kyuEuSTuJDVX0DTg14pE2
bGlo6oXXoJELiiSykmrPxgPVLSBYLg5kLyFejBop3QreCQZaRb+DAn88ku7Mxp+s
Sih4u5N269JkP/fUlTbaAkroVpoYHy5zHLbXcpH8XqWaYqJxotJ3agrtX1z3ZexI
zKmUxtFMhtTAoXUuCSdYvCilW2l2Mtf37PK6vPjAktOYhd4SJ3F0xk9VZ2q90Yhx
cf8+N228+Ug2qVovoFwBj0UL7ENUe5KORewOrmzEfWZRyPd0RCIX4gjhwN302fPT
iRFeGJc653IwYYB3BoqrhniyMkU0doF28JLSUJqDM76OjqPEz8WvYHpjXQTN4iCt
62tI1ZHEj0Odsq0pEejGpsNL3IPRR4rduQczaZQco6B+Dnljncpo21IOSS2N1R3N
unbtpAX6ojWmaDaRdSeoDSMUvLwyqUPiVNJwxFeH+JvMITZo5hyrBUqXiinVezFM
0rD+5Gx7ZX3950av7CjtYMpG/tpwDMpb74bGwXn1ZPrHJ/QJdNO8MV8bJGRWL8+Z
S9t3b8+tTC1VG/CCTRqqNdN/veY/NKLttEEdaGsFGVCWp/9mn0A+bVBEDFugXO+N
1XLLH9sU60/DHIicwf3tNY3T/YVMmTPf4xS+Vuz8cWdsE+FzrQ7dG6ysJ9xfBZrY
v1zBBY5hlBhvXTZZfCFRuTf6byY0pr9Vp0GdonPqQEE7OEnV7YGrC05Ue/KzKs1P
+NYd4N5h5V+G3IY5CV0bIqgqfER4fUs2jGgkGwpI0F/2K1uSPlj/023Ixo6kjerN
n/kybsr7xwusZd1G/8gQfigyJ/n2Uu4K3u4OSJaBl7IKAQovca2cJEU1RidexXRi
6Yc+vYff45gsNkKnDSArkgXYIcLdpuy9zbpGUGQQ3itqrziOM8QUXv7cyWp8WfEF
j+wS59Boae9vEHA/XYp8BEh/YKWH7YG2VabjL6TJxZZjhISTHWq0QwVzgiaJvLj4
wn4A0cP/+8EVNDXsb4x0t80/viHOkilIqIJXG0Yk7YEfZei+4ugTyz9UONPlJAXX
uwmHFXduhWgM+Se/3mVKGIceqnplbf3XMDBkgzI0VuKdEhBZG/qul8SD4ZBTOUL+
CHxgeW4bMkCzmRO37RS1gdNjq01JwRoicrVu2pFOPDHQbZyBhrRQWIMUKe2618et
+O1GWPBjqtnVbh/ru7o6GfQjIbRAUdJR0gYEdw26BKV6YuTDEOccxfHTJVKz7l1x
C+DiHt9bydUifLI/BgBUhjXGjYMCKUufeWgijGQ2j/WD/s0bVFqh3st6q7XhJxAV
HEweWLwmm/1lJwGCGwvnDURE0xypLcE6uKsNLlur2OeomT9aDjseVEFbV185MEvg
DiukDdUlZNQwkXWgJlL/vAHE7eJNfhLBpW9H/oVxyVXjbuM1alKHsJDYWVHKfK1Q
lozl9SZRJ18TruA7jdF4BJkWekQ3xKZ3Ez9sfXEcM/8HBJvWM4dDKfsQBv65pm4M
mmaxbQza5KhVe6LbVFZ6vXUAIEWJEEm/JOVivzD14RQjE0wSBqj+qaEfuNetnMy1
UTCicgCQ3tmi8WC2CfZNxGOiI4r1h17XfQhtU/QeZ8cVyNYxH/VllrEyqQQAinBS
xjeG0U+JnbHdWsOCpId2H4RbydCgtuivsRPdDVRIgU0gwquwgsIHeIvaNS8e/sSI
HnoAP9swQsjT9BpQsMa/IjJW9Hiq+K7np13NN7bzgjP/zidmxCBWhXRbcJ/ssgQE
MsWcFcVzWe8+F/ASaTP+ObWgDlgC7szJgj91QQKmoEtYTjjQ2HnRU+uw+tidE3Or
hBSqEfhWAYP19uFvYhWoyH861BOCyH6MIZTEgAnw3tRow2vwlxDv9T7fTEUd0SeK
Mfmy4joKsnUNnyeAMNd1lTpUjrYIUxL1KzIo7eHos+MaOQJc/ZXyu7/2ybU3ZmGd
d1s7hrh1NrUwMoPUDAUAkUTQwa/ICTszNI9fApQNcxeJkYVIwJ17eXBNPzGzd6ZB
FeHWNalQxPUdOVkiaHmf+3VGqrIG8hDJ+tZlZX13aJgk7wxjpvVcWfGkIdj7L4iJ
Gcvuka4pOx50ZexPNlk4ABmjCIEBP49vtA/8vdWBVlYG5R6aQ7IfBnkF+8x8i6us
AX5gIRkW6mtLpwc34z9CMNZDF1uKQpWCQa8KqCvJhsta7ZENA75x++4TbnrCwFEn
kkwnlAZPm3F/XQMALlUDbiaRkFnccEXhZT6TPJ26L/Nr6/rg6z+3OMsQtcn3RJkZ
CAzGBgABOO98epzqZ37s3GhDomLsVgLcW3LFpcLvVFtSgh2mS6E85quW7aO6f4H2
QlfwMzbtTq9AozF2Ew3uaZyhzD1WkmDavMahirWpfpt+Z3FLhJpZX/cQfTQhhkqg
GVx0GxAmGNzUYFtW3uDoWGN8IUyQaBfWtUQ0VEM/JcLlwW2mk4tOK+ql7+2pGF9+
EcDN3m4QGaJJ/7fCCj6efJ2ePhUcoYu7nzTC8qZ2sSTkOBcRSmG1XmGCT3VNCxVu
9gyaVxJ+It8URgzFq4M3pYdR+m3dbfIpdiaGUUxAd9CoeeNLFeXAkKdZwKpt4HAz
R6Ma0F//zxYuVdLD9XKCP/QhFdCzlhonZJY9LsR1ZPNFcLkQwlby3rEE7AaMEz8W
NHPVRwOe6uu5ev+uLz/4KmzSBCZoa3PlWCgY6ivRv+LmPX/gGCouEqqjqLjUtHd9
r41SuOHQt8y1Mh7sohKRBnYSL7SgkVBVRX/cHgBfbseqXicQ9pO9glxMSBv3lCLh
cIc3lwPRkwWzgpQBaiBCAql+bIpm9P2w97ta2y5P15WiqtreMWQuVcECyFilQrXM
iPXXAJy7f6OGTlu2+z5KyubU8AFONQ9GLdhDCH7yjDdk0Mp5FOQv4XOTJhRIdBeV
znGx9g8OBx3TqH7E6LWn/b0RIX0b0EWYHQykItodIN92ZiZtZp/QWhoz5sXBGHYQ
g4R5Orb465U+fin7dP737YDWCJpKlfZKkFeRXI+EPoeSMQvgugkSTvq+2Z5WPyre
MS94KxDcMnDmN690kmVyHlsqDUXjDpYR/5SJb7QsEauIY8ORPauJkC9pClPDLKm0
CvlgnJWEyB5Aw5Ewmcs/rdEtx5d7jDpsTQ+v7JvIFQx5xy58FQDeg0Ko3Q0FNHxA
ZQW3LxNZ4V00lLZ/F54lBGwdcfNvu5pIo8aczUkiz6YpEUg+GddRfQN+soYD6I+M
l8ZzxJdpR6ZLknPMiWrSdWFVpY3d+aFce7IQaVrTqM/a4CdmjEcitHvAa2n33BZK
lfoXg9AtL2FrMzHHkdmcecP9/KZit8cfhHad9lZjn2pRbqvmkwZ3AxOWLfUi/yBg
+39VJ5rnEdX/kT85XyqHUSr3giTUJz5HOHiISe3bfJdrFineqoafqhMKBR+VIvGt
XfLfqoM0dusWOoIAMDeKxjdrMFCzO+of+xolqJhvLe2roW/KciBY1UfwMzi+xFrD
Sfg/a8BNBP4RrF0H2Nb0XHUHwS1hXIKUT+rT6UEyOleaMwDw+1yZ8AC8avScc9s1
GYCwEwq0p6Ee98CpKIk5iw8+TXrS6XbTt8tPipIDpbNRqJVKZRlDfPavMiRnQYjk
hV4UMf/CfriuIuPBSoafM9WwXYzg5ZQKAVRunOroDdwUMGccDSv9zT0eehAlWeIj
nU5wdLEnxnALr0STCvc722+IsStZdlkHMPi6Vkd++ajBhap8g6E7WPn3CFsOqIXX
BHwPiGQ1euQOhpNwIKqrL+KJwFp+PJjR6LDi7qr1L9DQboLGkXxPMoi7X2UF57fW
tzgLPG9KvM6iiGFGJKc0YhsPRLqAxEpoVHrSaMoNTTxa4vw1eyJOxJFzTf9pwXpb
hDoqRjCOamxJ0G5WwXseMAC3qdc9BWHF2WznsDa7Y4eFJ9/yHcWpiQNyZttCEQuk
hi4vDGDyqrKfuLzH6NP3RqUiVZ8M7mmUP9IIPjRHMMKJFk1s+kF0z0AoLlKiaclx
fLLQ3YyJlnBKEbo7aFul9ctfd+DkvpCFEb5wZv+U45GPw1LRGsV7P5EVhGLfte/t
MjbsdKQ8aMvYSVtsaD9VHJXe8yyRYBILjiEQT2LNH3xmbXR1pEp1w9ko0KgFg0Iw
fP/tdPSJZEG7qtgO806Qcd1rz9Yo6bRkbGAAB+KPCzl2mWa2p/6KCjjeQskhGC8Q
07PQddFVTCkVQ+iy42T8c0rPATgCdCWAGK4STav1soYQ4yxwzs+uLQDHF9FOUlPZ
Ntrfop0ckq3a/Xc7z9cH1VtpMSTPpdKBCL91p/E+mRBI0VRZef7WfBv3tw3nrk1j
4v4kuWM5JYjUAJ3+gs7ZGJggJFcs4RhlyYlDUmXIo2d3aYtCKC9ojVKgAU2VKi0T
UedeyFTAnkNaY+TfaSoaoFAIK1Fk1ApTYM6Y/xsAl8e3svjWF2gGdj/N1ed1+yd4
+8cM+Z4/RtNdOXRW0g0dBLO2gAUU4/ln/I0BfITTQiUbQeW7dWXBYxNkFxf1aopG
/BNn7pf9LNZxtWLH0pUGkZxYjQlYsHJfe1FRoyTWOf5cerjriRZcKKnLmjemtc6L
q97Ea6C03dXhFBtcnffOnNy26Lp1U49TyKfkL1ioqm3IQ1pTFP+eJPDIws+bSwKb
c/MQgPWqz/PmQ2zU35+sgWQkVXbBQlcbM4kS6dtH4H8QH/qk+DQFg+bK/TxUU8wV
7U8v8CdclOeyc5dYzFEtt+DCesCyIzTgnbMD4CnIuOjoEUWtvK5t6KVGq03uxlKa
JYm/vP1OMi6lLBleZyspg2CjA+eshG96W4/ulgv9MnyFKTmYhqSHfUMjjThvsV8c
WNKMXmJfs0k9ObkKcYZe9zLKeBruI0TfYCGOPrs026KxBPjxyB7igXuNDLn20Kt6
q1/j/136HjcJf5dRQGL+fMpndV/OQN1h0e4Ek0qysYM6QDG7Zdpim7vcanVoKeJz
teeB5Dr4nrDK95Vli4F7fb9ukedK+yo0gUJLVjjlW8dr/yEyH2a44XKYisTghP8x
cY9vWHOYNCcz/GHHVPG/yR44aPDwd0YXhPGX67WktdkJFxHbRVKolnLoHBUfjjyv
tLK+rzfXc5syepvHDJxIwXpxQ6FF86aUXpMnEWG7MtALmy3aVXHcD3pDGxyyeOnq
FVpAkuUdIUl8UNFd7vo6i24cLF122IUCkaMAgAIMe2Jt6h2HpoFVOXq8pv8y64d1
4t8ii7WFMNlER7Bs58Hj1hE+2mztSaA20Vqhmi/Rk1yHr5v8qVXPNMv1pseV4v1t
lDaTWaRhSLCtS2ueBvAn3CVEuarfHafqYAGHIt2adkier+7TrEctm/+2wupGdG36
ZmqWeMvoMTviq0Kxy3N4Kekk/nvlXsqHnFcsKZhHVjAe0K+x/ZFET2qdF+EiaNFt
fE0Q0WsGCTAUIOqiIJJruXAQDVM9UxjlXLzjG3DLHoE5IZn8Zv4nurHdJg6LL0FU
2yvzXQ2kEGg18Lh35HLAgWuJJ4qQhe8m52jlOSlnqqCcsLXdH/su+4MpZCti9rXo
2k1MhZnAsTbjjWhlttb26sI8lvU9NIGBZSbHZYczhoEo3l0Y6GddJTXjAU05vmrx
Jm1Z0tssVEJ0JjPFbNBJKjLHDI9FwGO153tXmdGWlw/CLUTv7fdM0I2tIHq+jqN0
K6omrcxclgRVnpSVYnss9az+PdXP7phsEyko8fgLbl3PlWWCtYcxTvKcMmfLMMGT
3ddiFD6hBy44+c4oW1EKe/h3ie7llguVAAbQErJ58Zvf3Z8IycFyx8V0ZI/fpErJ
UpSsemF0dSGyTpt9gnyaxP0tMNtD651WXCocApLzB6UPXbtVudHVXVlQ6aFxXU7V
vzdO7mtqLCRSU3YchqxIpgNvX+8n5PFgUk/Zak1txGMYYV65som+IUPwN52xVdwj
w32lhBaTH+WWKT4L+o8wIVnA8mEIleXxOV9wHmnuJYXvDbsaKoM/OiWYVFyPyFhc
dwDCUlK2bo2Ow9LQz/46Pmx3UD+2lSm6ZF7Kn6YviIyw/iI1/ZjqNic5xOhHl2xW
DND42X1Rvcmo/zyYrfE0CmPanyp3o3yJFXEDQnHK9Dr+ZcR/l+N6ov3C0KHxOBFh
rfoLG4iDG2mSlYMXn50u9+SfiMYzgyDhqEnG/i8qpaNPcuz0Ah4JLAZVwv4eKIgs
7nFktcP369D6tyotwncSHr50HjhpCEkcwaAsGEKU539gXogBhXbu/8t7rtlTSlD4
LODHNWWyEQUZLXFTQ/Esz5EwcypAPTOOjFl/V3K+r8O8BgPWW39UKDSbfmufWJZn
hh+leGCsGFA2cIar+u59YMLNQzuEPrrZ2AbDnzCb0N03pbRQ7Z0CSUIUOjiqKLU6
LbXW2quT0t7xwRrXAjxYStAO9jMVsguogPA7YPkD0tydwbzeINjkYlodfOuDA/v8
Bq9XW6jtpWiVFxIVnytF5dZWdpSab0y2rJFNObp3/Y/EwSfWIqEdPOJwbwhN0cz3
7+ibDGi+jfrZ3Mh6yx+pMdVyrEaBD7ZpyOgb7R6PUyaxN8Uufci7KIcfjiFnORoS
+w5Xgxtlf19rBijWNieDDQAEXQ2qOhv9zcM9cZFXKRgUqLx3kKlgZHeR10RcPhv2
9z8N26kQy3s94ZubzxjZsX9MpajleP3HbD03PmIEUipPcMr0Vk79zJ4k5DzeIDoH
iFtBNhYmtd2mE1vrkHJKTewmp6zPW0JYWzpzYm8iL1qzkbRWoNxI/wRhrdOt0mTV
fPBfzfqNVqN8XIu7TJXXBqKIFPup/MG3Bp6sVq01uEtlRs47PyQX4lDWXdcPGle4
3wHOnFSWn6nIvLAF7LJjHW2N6G/fUiCJEyjBwoQGzFx9E4YLf5Raj2NMZAamxMk2
AIvcpEc8HIzdf2v6PvokgJWT1u/nSfyFg90TlVEQWh+QR+qjYXhk1vd2tvs65mye
a1ZvYh3KHlq6rYsxGUi9Q0JePy1jZM2k81XBFguA7bb7dDwRZPbZgSaZeaNBRkk7
yckGquZqe4UGfk5rWpPU26Mv19sz7UI3Ynf+mKSqHekKkPx9MW9xNIEE0eBJTWqu
RJPvgQilHQB6f8u16JpTIaQLaxh3dZA36GCSh2vOKMQwA2JavIv0RpUpKJr5Ka49
WtLUiMXMwCMXKfOZlMYvHgeCKIeW2hAqK1kVVm7ijia0jjIQ+fp887D8Q5NGGT0h
JnDPYZC5ZiGFCw42tiBZkkGKuYCr+o16lotBqXX9UREbhzeiAThntD7bES1778qc
I7bv+Vu6Bv30jLYLLW/uHYMjW7txkHG51KDh/Auw0nxBzITa9Fe6ntmWpiBOWYT0
p+hb0rgwIT6a3hQShcW5FE41dQkZF559SdjKWmS2X+9clTzmdfH51MIlyS2j6LjR
hUppJH5wUahaAULEmYF1q1k/5W6r9IHjtJsAd9nxM0XDRQZL85ivJFJkY80pe9Qd
eBiztj87LrSmQ80zqegtJxoiUauw09ZxG/SY69DXuLOxZY0Sk6m0S3dgSNMV4/AR
zu57Ltc9TW554mE/58pVtcmWSPCTXckJe7JFmYY4FXRmdIsDkAWR9hrNGFJnFV29
GdYUH4ifNM1VXj+xXgVDoAoei4mClO+I0gmqOr2KLwi9oa++b/ujwkw8LtzfjXmv
Cns1r6/7ds8A51jHAS8TxqB7NRTMMEdUtxcwmYAHR/bUWkyDyISTSv4uqTjmK/pm
qMRliLNJYwFGsWSaDCw0Dt+wpI/AjIIvGq4uTU+ZDcaQbtQ6jl2uuTagT2iRktmg
L7l6iLZBmlBo2BKIDJ90kuXaTLgOcEfvGRNJ0SC/ysc2uLI+TvlDDBeKRk1jeJWO
2ZgdXnt0ziVA8acbZOLJAl/mW/mewzOyDctEgKV2JUEG/LQ6LhIFtZsBLahxRzOT
9yn7zMUyDNSWsnSOVzlrd9BNBZXaJ3pEnp2CxmPOPZ63AD6OUqZTFwW11uf3oTPN
vgsnWwvx7/P3gRZvGpFFz+9JQPk1jhBNuMA/7pvptifVi8REkYMKHFFBHPfI9D+y
gar5HHl4IHgMw7AKG8q4mXLr06VCn1lqIeI7pwTG9RoFpbJk22taRKLtzxAoGoQ9
hdAaN+h0BL4Lg8xuHdhDF09c5oW/iMxLE6LqulNML0lYjYp6JuowJgEJx5X2Ayzc
o9VCHCObLuknQCskv4bUW+hLLUKH19NL4TqrvQkNBbzFCjwKLpeSVWRa9fL1qw+X
nYe9rR548AW4Z8IqljgCUSIsKfCbZP0RfN/X0F6Oo4WdOhrW3VUK/aAXaLDNyNc6
Rxuh3KoJ07D84dswid4YJFm66kTzY41Qf7+JAmWm84yo3qWNnf5e7i3G6HxxR6RC
k/gSOuNbM121M9dTq5Ga+Yj8uAsc3QgrAsnS/WYU9zYsviN11WQNwDzU9Fe/IiqU
mAxYZF/eFVixOo0vm37k65cB9gTRdv8hjRo8v9lhjmweu+ICPk8F1SkJ7DvYMiyP
InHpkSgGPrG3LUokjEIM3o7a1CNfhuO2ee0srFKrCUVdoz5dtkQX2a2T6FsDHF7V
NHxjzVtehwLXWtgny0btZBgYHI1zS4M/K0Z1mtcZ8/fM/lWZBcbikYKNpKGj+cTp
KRFx/pxs80HuH+Yy17WcC3qO0weu3BKtloTDJD2dyPSpOsKLE023N9wu9j9jXGXQ
oIQ2QUXuTYrEB3hONWtesb5q1oMqPgPJDehf0p1HO/0guexZ7ZukRbtlxWc5wT4R
slEmiUbvME25thvF9Pyy93BcmcGGvVhdTu5YcZTX3xEa6USntDgBZEPuzy9LZahF
1rYqGpwvAHMndSASSHB7JUSxTo6rHCws0RspufGpTtY+sbtA+67LcwKOlxBUbmQO
oJ2UzC8aSPpzIoS+JKyA2MfGGyGzgQhL0u0CKDJys7Vr5TmTJt6o/rqOpH/YZUVB
rw1LCB1hwNNhxRtr+AmC5tYQSfHd/HetFXUcLaZarStpwAzk/TBxST5Rtb27l0Mu
m7OpK4RqXwVAfsv9n7lJLC4OLJRhUCCQwJGt0bjuhgLfsKQi8j+Y8TaY/KU0xaa7
OHal178hMwvDdgSe76yrqPBRUIYFta7CRP5cv0mnKfLIoMdJ+jZzhg+oGkD8PV/f
yb5ZUpwbQbooHgFmNVTNkkGAKN81gqOVoMQU9qFY9oH+7I3TYX+Lwv8d2L2t1on8
zPcofubdSa1aMeUBYR6ORUTe8g7ZZTxbO2wxOZLCAAac+p5H4FUcHBEJbVy9cSih
n4i85qYQ0BJXHlupUsDx+6p0aj5R2Kt+ORY7UBE/CLrOE5sfA+xrRnjY6qdmhAJq
CiGu4N+bl6Ima4iJXlfX8gI16it9tgNMOe9w/hrDxOOgiq8aVtOuzN4dUfkiMc3I
lBeTE3hVfHYmB4FK5ZDxJKsrdCfM84AIfqzthIUe5lsrEMXSgKFVbxTTJbGKgBZh
SFROGeydrvDg+4Na8Z6LyEU6+94lyQgI7xrsvyngC38ZR4TYblc1dKZAHBFPl/D4
YyJ+lTZH+1i2Dmv0wM8W39aO6jnQ17eDZifCRRyhtR9gBA3UgyIkTNldF//5vy1j
B7yoE6e+TnfC2z+VoYhsq6w/gu0oPlcAkVedTPDRFYt/qaqS5rDnFHUqOwn7DMCP
nsO44RsACqF6mwaxrU5NNBY3HT86rt+8tsDw3R+yFQWsRZfWxm+AkI0V1NFdGCqx
J5SYMJ1ypEXEz8k6mv4tVPnSpZKzL6OE7/hBlgW9h/SkdAvZ89OOQkl1Ek55tcNW
ZMwABvjx1Kiug2f5yo5B3gLVf3oklVlP6wxWAXW2m77DlxTy3GT+r08H6igsxKY2
DKT0d4E4cOVfPItJt0dUVXwDCTIrdkuliBfY169KcW3qFSQ3yhtsu30B7vyw8+f/
3fFEnHKA8mXAZxYvLT+CQFrM6mu2q+pdU4d12wGUGPhKpE2YHd74xrvNv8TAAMxU
BLnu/HZ/ErIGXMtblm9m6DoGQYj43LyIzvdM+c0moPGzyQxFBWE40TkVKorAW5yl
FPc/WEPg5aZ9BpU3k1riKK3Kjoe6Qdk168WkmbfKThgvGbB9czWoBQ8Ds9mMusOj
czgD6+CxeEYCbhVE86cPyJrRlrjiWBshJaGMWb8mKU2foJqj+fkiUSb90DvI7wwU
8RaNOwnFHAAmZqAua+kl7DFX0DqZTFGUaJUv9jEzKu7sb5s+8j6kR7o1GGkAsRIJ
wvpZ0UYlFyAe4qiYUyuo36Eib64OvSBKUmkDlLuJT8lFwppROj/yO9PWWI3V5y9N
P+Ba07B2SS2x1LM0H8qlz7Tzmk4SNqU38gk7xe6efIZ5vmWVY/p/TnNGU1kCn8V2
DbHLI9OekvfuYIRSolfWAyCNSwa3wWpwrQjNaaOyLewlEMBYD4dGS0lYXdTSpn1z
AyGkgNB5KKrE6WC2dV9M0HvrBL5yEMAiZudM5eXlbAMvpSyGHpw7TXAM58TPFj/M
TytpL7gOVh1RMNPtdDXQO39Phec4SJm5R5DRzH2EXDF/MzFEqprFm0oGS1Xb8B4o
OwruQI0n0bS6xElfMgEcVTI3MKXlXh1Lj5+asKK4HwAv1q2z6gA3VeAPl+3AvoqT
mK4ijD/CymuxbjINjHZQNIHrk3rznQDZydDH4H1PYtZstAff+HeDjFrFJuXTppgR
7Vjnn6XK/oxJkCtk80dgDSzSyQrCyT2pnH5SIDZhqZ4vG9f9/lI1ROxDsmVgh6Pd
q1Wq0ZRaUhJFeM2hOOXAoCYJsI46PwwJsG/0P82bgbuEPh96+jsM2bjQLMplI17j
Y4H726PPm00UYJOLEw/aENqONX/SGQCwVXZaYL5zftPBiZ3H6j6TJDsrD112CxRi
0cVzCr1Tli4TRGdon7guehYxktYgQoFZFbCrCgKpWh+T+3UCP597RX7Z2v5MD+l2
cP3/RKinwaiscJBOtLM+IXgF8Q6+iwwMczR1/5vBIsi/ZzQ6+0+l0uu2/tyDBUQj
hAaR+5HwhSeZOeAB/HHQndMsSSHheEsAi6ununTg0Tg3sOWu0bhGYU59MZBfp5/z
5ICI2Xodx5vuASXUnAQ7VJdwPtLqCN5FSLWATn0n1ldlDASeYToHiDuujKBFu/Qq
A5ZqAMvz33Yf2y8swLEqBVBhJyPZL6SVolsobp+IRGqVy6qyvtrkrVQGRLZX3isr
nSdUbvtr9g/I5S1GbuGAZ4xqW8uM0LgDyq+XfPTJRrH/PgW+/vpHZZtE5RBA5Sa/
qngFzmBHvFFsATiLUvIlHNdgWjJWznazrnEKyYD1iCDPsTtZu3ER7ITpdKtigkYm
h9n6h41VNot6dAIr9lWlTfJZn9sL4nwfL8KvSFvKPigHL4GMWx2QiMRk6YsURw1r
DLdpbmoRNUO3czNoFKuEvdjzMV9B6K4r7VTXiBvdIRwCxat05ruW/DEMhRUmZ2WE
F1BvJjxN/Bli95wPXiBWJ6LTLefUZ4SAWPurMBA/dav9aP2bz5FgsMFQVUfk1LmW
G6FWKYNU6fm4qXT0NsxcNONRXkzdK3dOJYOYIeBvNqzrk8WDfEOwwmNZo05aQfk+
T6lvQ/1fIeyDoXqYs+fazD+fM7oiJPWzUr557DyASGO8Dqia3uHgIggvDlTjB0YR
/QtAV/a3iuB3ROS0xWHoQ4SKwP297kNqcnOqssROj/KXQGQ6EhyCcns0WfRHEl04
77fCpFwm0mKqy3KZVzb4dsvGK/cWB0A779vk04p36OWJtVmKQY+4pHKS4CvloUuQ
MPt66TAB0XhEG7VVBrjxTpGmQOg8npg/9rJodn/UH4LXvGubUazzzduCdi8FlT09
DW0lVTP8TUZBPNL2mZ8dPRMD+sUPjA+jl1wGU3R/gCZJ8l3eQ6gOBpqak/1di5Co
uehkSlXOa43tw1sI4UBDv3Y2leftgIF92g9wMRq57DdyNDbuZ3PF9dOYRjaPu6pG
+M6v7pxaFk+3vVPRLNGrvlct0+PaZ2n2F1hjjKXvgd631NOuI2cDIPwVRUN9Aydk
LqthjPoEr+O/n+k6MyZ7WQh+tJFrtjeQdsuqo+bU+SoeX5IAMmzFN50eGiKjM6Ny
AVHacS/uvxB0ynmgvKgu+63z8x2yEcqEfljy6YDCU5Ebt9wnrxKbrGikKVLFpsp/
GO7HR4v3qfhqtgZ9ciDjbwQMM3CkgGZ2SbSJLaeeUg1u6O10FFoXkjoBRuZBxT1K
UFfh6+1ebN6rrqIlsI6U+2qWxcu3KkztEEfLFELTr8FpNQveXL0ab7qS7ydKLpVF
NxNW9FDHMDZEoqpGscAPvlXC2qIO6TfmIYjvHDQ1VfRx7B1NBVP/T5OsnhxPz1Vs
OaI3dqyS4V/tI5vsyabfW6/+05suVGWECtS/HpNcCbuMbcU4YSoLMsiux3HC9HDX
xAwEw4d0uI+hq9A69WNOusDeMMwIHM6LA9qJ0HY/dbQDaPViL9mxWka6rX4zP8iZ
oHKfkmvwdpd2CZxucqBZiATT6Ge6Veh0WQ5Rl3kMvZil8qEj7/YyA1JCHIjQz7ry
/lRIM2+H/h+tAwaCW+jai7caOwy7hzmzj4RFV1gZsdaq0TfHeimnLdiLKTWwHjtw
EdI1/rdWQyNt7rWsT9eC4orjKjpMJzYK/+v2cojTMinFxUK6B0R4dYP13e3/6fcy
SzfpXNgWG4WzOTELc9ZN0fJD3NUPImSH0npNz6ZplgSxwzv6DMO/hsGKRnbxzyvx
/nChO534MxRj4jTb14V40jfhr6ptR2i0BNjCduXb4C6YeYMmkTj1KepjyP4+IdDq
fvEZUZVi0m3F/1L+0Z35rtT8wVpCeRuBPotlMHUXNUzod2gyR1Hf9TFoq7GMui1x
cRifFktEfRB/AaNVpfQg4pwL4PRIzU/UPZXK/2nGvtTv6svf1t+yM2T3bQj3zrkz
usmKynnAa2X1yihSFh4HzZJTdUROF4BnqwOC8Cs0icrksDGIKR+9QvwDlv/mXq4m
UShvDt2T4c+H9amPQIVLgWQHLQKh0VKp6vz5OJh6O6i5pqFiV/ZdtTXnxfpJWco2
50fteZ2q3qQwAuxh2rFZNNmUEzJeNg4DJ74ugEG/2pcULLJg/M8gtkQIBFGEhTsi
LxHj4LoNxX9+Mkb2r8tpwRuWOzT/J6IWmqEKHBkYs1ozAV/ctdC80v15x1ELxZk2
eCVQ9FSgHJWQ1QguHP6/wtz1DS52jAKkWPcD55Vs2x2kOmOgCAROtrnFX8Ljyibc
c8a0zqdpNvaD5I1DbLa4+AtVUxYJrer91XTP9dKWu+FjixBstZpW6ug1nkYtYDmM
ND0rUjnIArFqZvIp3vQ6XtIK8hr0ZC440qntTWjPWBRKMG9BhOpk199zh+n8kP7x
theqOLfd9LPtRZedd4KDgNrZFkO9MC1I4l3iNfHgfFj723mG3R31jtujC05juLLi
RrTJep629uO6xELuvkyZRA99JqG/EcRz3zc3sjmwSf63YiqEM+4SyqhZat0NGIPI
PqgxUIcjjlc93+wgWdtfeFSMC9pXSxaqvQ6ZBpZkhrhr8wPXS4QyDMkgfOQ4AbzP
dY+dA+cPcItAhLTCBEwu29I23+xUlOvhjN5jMzIUWaFYkgH3sWI9MMi1KR8hbNbj
hSQJfoW3lZqZlCOSRln09CqK8D3eNguC1bALvNk3Iw9f8bpRmMNBPxXQwfe4Zuqk
Ju3yANcX/xQyJceKGCm9JAztrhSTPPuKPdvzWS3bnwCI7BcZX24ObU4ewhLchnhM
r9KYpgemgz24a/RSm04GZSRmT51y5v0SsrvurYIJJ94fpCOd352MiqXg45tJ/8jm
jFvX4NcMm5UjXMt6bUqnXqv6wINV55NuBiF692/jp38rfKbraCsxaxYsK7fgJxrJ
mx03C/o01slKQ2tiLoGRmFVaq9k1pnEiY+1FYQ/BxvtSHGJvnb53N+WJQqFSx2VV
E8ZvPwWzd7G34LF8p32nrfUMcoXvl4pqu5ruH6Su0eNrPUzafKHn7vqBYxn3GTFf
RtFACfmweJJC6z+r1TG6Bxv2FjG9uYWVDKtexp9vaLC+8ljVEIk5Nl6UexgcwSeD
dmHlLkTGADvTmPywFOw9bVc2nfZEAiX9w474yB19BW9NLtN4dz26XGPYaiwAZ9iS
7GRGYd0LHumko96fBh/jvy2Y070TZU4ReOjEcl3G6yvfEsjicrmZ/Gi9Wn1LAPDC
Ki5Kz4fNNoSDHRf3S+ABO3miU32oX15dKJYuroCSd7twthK4/ywYTJ7axFcn2OqB
J9ZRXH9EV2IOTrt7t2EvvE7STLY3pEuDC0PhR2BSA9eo7orVhZ6NjuNa8Kytrj1C
96xAzJq7bIsN2tBhV/0qTHHhS8RQO67oxyeyoOdvYoPK7DtUCi7maQb+nYqK7mfs
qIjRkWv+pf1EAqebUCodcEakmhhNdcLy3QcSbbnF/29PZpBe09+4SxbOI16pH18E
0Fn2EFNL+G6R59C8xUd93xCE9TBI5kUVec11KV3dmjZhmVbzv6u53f2Ia87TEBUS
eKZUWuBGb+/YIhFYg3lyYKlV189kjkBZv2/yatygT7yQC4UtPlW/H1cr9zlxwC11
TQ3jl4QzoClj7GFF8a86gFCNdfvapm1uBxjseY4on+vguVLIE5GC7s+2gA8Xiwt5
3+XuZVwHWtFB/enqH2He7wt3Pl4zA+5IL6CaSUhu8gsB/7Eg+nCWVTo+QI6BfSa2
lusVMjnuAp4NCKvi/Pc0LbrCUqJBku2dvH7JPa1YuJWZET7uxek/DPjDZA2JV8zz
IcBI+xSPWOtzaG8p/jeIij4YgKK7li1mGPsistF2qUBvj9ji/bXNUxoJrerOnwWA
0GDP1abTYGQkvcvyq8vtMLzp5OPCwneSpy7nDL0ECM37Rezu6v+StIbwlVy1/PDe
i0Nt+KljNmXJoPAg79a81PjUiPrUYWoCMpSeWu/5Lb27CC2Lq7C+nQFWazdTx0g/
Cv/zLTCbp8cVlsKOh4fY9U/UbXCxahVdEM2KRgxT+Qbp8Us/AswF6ebZvuhYUJ0X
T0hkY23MRlnegwD+jQDS2TJxIQbUsfHKJMW3vdbE8jbmx+1SeOlHq1jv8fIucOus
ghPxIF/lPqLevPUb5jyFFD7vQyZw0MwJmXLi/pBX3aiNw9jOHyuM8nd/w9cBKHMS
q3fqNOJ9O4CbZlFRjOZ9Z+lIceFlw54Cg0quuPPVJOpEAG1l+ojn579azeHwsdwb
O5X/xG8biY1hYQhd1TOPQ8u6TfMv/HwWLXC8/9qP7aONBCpi5nBYMwrhfGT3AlOp
Th1cFdC0HP0VtdeYtydraPqXzF9DwathTmfeu4Awf2PjAL+rDWH31qY1SCVHibr0
Z9jDrPGi5J36c7DZ0kiLrPp7/OG513S7aQBm1n8+ulvxSIYzq3XKhowuPc9/oPhx
4Dexyck46k8orvi3Ay+kdSU+5kIwtiOSe2PbPT3xO3tIvGnrGthSvDJ3SgM9hBtP
2x2Z/hvX/DieNWYtUIocvy2IIhxcEWHRp8elw7VsTKW8uXK2znaICiEiYcJsuKp9
Wfkmm4KTKwwtuXaZpM0SDc73q2Jw6OIn78SdHQ0WNUr2XX3gMJehb9w5AJFQ8Wmg
xXQz2XXWSW2B3niqi0aXDJssAG4NGvBqGx2Hb+jMUvr6AWUJ3dcEwaYQf7Yec682
HYWZwr/Zp5wvCnrjGOqb7AxPfYBREonGkN0d44F/hI5frHIpA772xT+hGVY1SeNn
N/xGY6e4sQ97LrrOBeLJx0hUfxLLAf2525Rh7d79rOzUzPw6QqNfhf+SR8GHgOfu
PdLrYjR1eqr+aEP3HiYKHSUs09YSSCHFH9m2NZC1nRBvZhp1ccAWcxwLG+4Ol3qD
qhgCBtaRWVyfnokUuYwYdCrAdqy8hRGPBVCieqo5F4Io0wgaN9y3p98+QPzIv3PR
ryIFw8o5aJLV1k2NLljFXr2rrLqLYw8zHJTexc2vo1rkpJ0p9UP/Car6w/uc3K9I
cB55pWNb3uvXAedPhFWdykm5IB7ceD0JOX5dnJ/aUUmeF9c/OCs3wku7EfDDKYI0
Z7SPpcsMCQBJZ2BlN/W19IUx0MUmtK/80R7PuYjS1HJ38b+Dk6n+sNBveED5hQ8e
jrWYBKUZ4DuaCW0g8tnytg21fypRh9oJDbRUdZjvz/ZCXHM4o5pmCCsKVy/zxKXK
+JIeGOYQm9wI7kySLO7rL3E7MMXDUsgkKcQlzVOEQ7fulF3cLPnPXSfzoYVyQ+X5
96yGe3bd+t4UNOWkpIwOFq0JAyOEyDiRZCDovv+ZSymcCBdx5eqqcMTMTnYUChQO
BTvigR8AezmJzQz6pYVp5xWLV0cJYINt5Hf/gWh3Aar/DO9EkkKsf0ylcXks8+5f
CO2Jtw6i9CvlS5d38NLs0ZfqF1ZzAuzvaV8aRWAgcgBTbVoE/ztOiH+v/ncEHMB+
BitwGD5e2xLa6FyGU3mwppYMncNnoUSuoIcGA+Bw/xx1Vp78Mp7OrCPNjZ0IF7RY
XiLFR+q6kmSyD60krZpiO+/AiiSyz+GcuC8BBvm0e8kiX41JtcJ84UKz7agWg2Oa
pqdlnH0xGW+pKMBRBkoMOfj3D32Q3kJgN776hGS7nGm/dPC9GJ26KXE1LzzWkEoU
28B32BzN+aExGpaXzbvCaAMrWpCRV8Sw8QZvlHQAYCRnDGy5KxSACFHACje5P3wx
HGoafq1NdnD7lHTY802eWRV2yh7Kcku3ZK+JdW5CnPf3tWJVgDmHWzvlLvsYYBVY
7Xj8ZdK376qaFkQqGjNsmNogK18qIoQFXxorA9Xp5njW3QYFmoTHqL2EJI7PgQiP
j5L8jQTHFJLnDbO6saXuDNOU2HdB1Esq5orSqrmIPfiXoIdvOUFMRVAoEi+w0K6u
u+aH8hEUr/pfg/oyfkClxNgVFOIFhJ8Py/1oJqCV68UdudMS3s1o/P7AL1+Kr0mq
zXhpKKhzqiJAARQVK6FdkITcAp6v1x5vw8wg0hLuOS9RyJJ83axX227S6LQeyzK7
KQ1cXmGl0U3dHpXwKNUTj15JlG96/UJrSW+jWF6TN0xaQrpW1hdK8bFAJicA+/Ck
NNug99UlyGfSBfs/CdIFV0wE9o8ILkHLaI13ddRmlLW88/bDU6HuVePtwXultFSL
7SE1KRX5rh+e6uX0Mctwwfutel1PItLbZeXlEetThjFnQqdL7pToDt3fvtqq168i
5vCqYSUTLAY2YiZC9T3UxYqjMeS1YlIV6cM6lwnGrghrhVNpnqee5UWq3cVMvZT7
aGmrFkVgQE9iVCOpDl9P/2qIXbNxCUlyg4/fdVjJRJ7YaNYBejHjCZPAdV6eSd1a
77UCDidGXokGC5orZdVc7LDOnY03NJNRpkNPorkkdrmDK6kSooiEbRkIMXokJNq4
9uWahPijxLERqSnW8VO45i9p/5rLl037CllkA8yRhd/fzS8w+B8Mksj++EV1Yp3P
gIMbTtjmp0FNKivBvAvRqfXtPxtGRTpDaijVSZIFqpuW+Ib2DE+OEOfs0XvZ8gjt
FCUXnElm5I3MsPzdX4p5CndsgqgEgWk0eAs5FCPEdBD8HHDZU86qGOxLQj84HA2O
yJFCWZB40wt0i9MmmRHK0AuzsElUoH4yYzd3SWqh1l8UfnX8YXp25vBhX52Y+9yk
ZCi12Wme3SgKiWr3zw60qW6vu+tW+24DMbtY33oSmxpR9711fCVkJ6hTYeDdM2fD
9cevVr56BBGaUA9GTU12ir5OO3HMWcAU5cs/BA2df0/J9Erh2x4/lbItxKw9WhP8
+TVdgdug2zrbnpzj6VvlYlwdMvx5RLP3E0cT7GpR2m0yZ2frEgxgfIgLea483fSY
8hreWed7R2FM8APHVnK+hazvee3/9OAw0IYI26ZiVR7fQkH1UWhjLBAleqNG99+A
79FI3jfBc9jkJtO7z6mrlSRnhZHkn/sDER/HQcTw5E1fGJm/84K38NDc+Rm9bgqq
bwFMy1FtggwEuhTF5snp5dN/lXDqcC+CCwpFRqPuiMeRx5w+KqYIO9F+bGiJnz6U
usLg8Gc+PsInHN/nbbejog3NDsWRw0k5wOW/vzFbaLdWxCG9QAP7wyb+cUkoDBAl
W9TTUaBLwLaRkr0KwdJKTLaMiTjgoN6s/KHLMK4kCUsKYEBllJU/SMCOSKd4B5Kp
7Un5O2r7r+PiecOzUO/UMg5uNNQZmWDR2FfV4c6WyyKtHFWgrUO42cvoHVdhcNjY
sjbs0+T3NJHFNJvJo86474voUymPDTPQsIYCXKFMhEIQOsw52Oknxf8KioBsQXfc
6ks2ooROFVKHHV6rfohU+i6LA7zSXNMC34J5C+b42lvfHoKU/brGEqzCx3oDGLeV
cwEEmsg/0svS6COL4iP12VxH/3tohqgx/Xirin80i+O6vBawT6YYOr3f5J+2QVxn
axvKPHYtn8SnmsZ+E96MJLUvtZpq2YbhAAfOivfewJ3iD/8CQAxzzngmGJLhRAKU
x1F4VVdBf5LKMusGaVkUysFBUuGTTuZA3bdU9TfiQgm/rtFaMuAAbd9vvG8FyeP1
Ch05kfqVWMYVjB2G4wTDg94mDLQ5MaeAEtSoSmPxj2YLlc8s66XUanUL2151zJ4e
5474ED3iH2psUME/2zFamO+0Obq+7/ahTsrNtulPQkIlrGOEnDDdTzibJ3jZ5bRN
wh3Jk6gKo+625NoqlvMSEDH1Hg2fUBTnwCQN6P68WrgtfLg5qoSe3mrBgzfSa1qk
SQh1EUE3bLP8yC/3Xiru1e0kiRKOHWtNHoOL+NflZCHczam5N53QHzOLSy6j1woL
p1JkUrZ8rIoFi/KSYm9H9RLVKFqRKrQN17ae9ktWXWgaRwjEpoKR6IqCeepuIo2y
o0wrb6ucxtHFhnKwSc479RWEKWGvtERuelf/djbvAf2nZ+2+U9ob8JNISN1cXheV
BVE1ENtJ6FCIxXA3SxVpweIR50cNOvzc+hHopNdPhgTiqvV9HhoqlmaAdmU5/0MM
6Pu+sjnmsYSHCd+Qa8wwZ2ElXrAx1JSr4PE/BJMEXPUTwzMJ6ptbVLqATlRckKHj
66X39mr+a0GiLHUYMFNKqQlLhPMTl0QOXI/IOrSiltMlm0XBMpbZGc54Hl9WKcCm
YgWv4p0WQ0ZNTRlcPsiU0vQWu3uJsVcaQuYPcIV5V0o5Z2fHhsrmYZ3LiNjv2rSi
HVmUu+5dP3EOmSANlC7H5N7ARJ+yP9HaMsS4V+Xblvr6CKxPV5KQyAvU0M9V/4DQ
k5gDp8obXYK1Jr68sLZPJu8BTAAfEvCsAIXO1qK+Zh/QRx/FMWIwxUHoQRv4epKh
Yn4F2SqTN1dgh8+/0bAv7WDK18U18O2tjgxHKfCJRQd2R4nUaTxLRvJokmLAnu5b
LJ7a3QVd9WRwixVNX0q7HKAME4Uq0Bq8xTRiht2uaAETwTxJUQpmQQM0Y+9qAkLm
Z+5mekT+12zEEYi5KJppCHNNI3Im5i8shOBsB8Ew+VKEUuzllYaFx+CL/yf7G62m
FzaGNUfvG9490GeALO5XUUfXr/4bza0mJs/K/YlwFpegwoaOncPz0zUIJJFvcnFN
SmjIia/YJLemeccZthLnWfZWohdLGbO8Aw20Ps5DltNUJntoVw4zqDE+YpQJ48vT
avtfJF6Hz0q2Xd/H0gtmahpImXRor1Hfv6aUQMAaO6riDlbOt+ozt0znmoc6gv95
5tarFuDdhJ5KI+4aEJkeSxFcoBkDTCVWjfYTPrXobJkTe8+fHJcEzu6riXm2cRbq
A+Jm9p2K5iSklump6xFh1m6L12M21SV77S9qVnV8n76OlH/mKL9cPfnGDtcAF5ZV
TWDmlZZtYJAdRDFihTiZc3Z/+vUsapV1FWPam4XdQL9/4Sw/fXo1lvh5mI8g0436
2iy05r6w+LRoOugIUzwzEJlfDpIx0zvCyFW88xYSgNbSPkdbp9LEMNPuBikYoJ7j
LuhUxHIiXUZar5UJMizjpUEj8MXR8wg3bcw6Tytb7anyBS8yMdVEuDTXwEccsk7a
yh/giS/+bN2sVxGfMh3x1h3SOTei1NZcAI4bZs/2OfBe0EjeVEGBDN+l7k38VSya
DXzTXszE+Tt4wVvTssz5z21PVi0e2LDx5erx43q9AJ1Hsz+dFnVHtyRjuQCCyRc5
O1rEjSXKPccEmrVrFfD9CtaXoPA4VUl9+ls08SML5nBGyulCm+onAcCGFEto82Yb
1uN1+gcE7uSxu1ZX8yfMicwwMqqMdFbh3c+CIcIXc7wZL8WUuHu6M/XoqYU8NM85
DjGMg8fKqjiyQEwd3qqmsB45j+YBot8sDur0lZPMUeCHF0tkf6DDzpOjbeaCj2LA
d/58aykll4z0A3pH4wRuCSrAV4dZutOBpCD+MTi3fM1Ylb5jQ+uEx/oSon1K8P4G
hwJ4eGVoFw/IgAv+tluG3gdwNF3BOhRX7cBBsxTwpDXlB9hlm/sDMHM66esAO5RS
Mve02GAaiml0v7xggh3X2FNJA1r1bzPOkEjQxoPUWY0o9QWG9f0jwZ2tBGsp3duU
RhJ6I800uHBH7AR6D2goTRnp6vukUEiBRLXpYRpFr0cC/s2h7dMaEkCqKZUA3NHQ
ur7S9N4ke+d6Ght321W7uRhhpuvQ+Ff5+0QSHV/hg7cKMeIR+gnPWWXV2EEnCzsz
aH1SAk1hhA9p6Nn/yVjF5VH6pFnR3ZH6Xu80wiumN24IWd0vh7i6L7DmIvdFbVqN
sCypaVvNDo9mVT2EhPeAVnM99zRiBx+faylCk7ko1iTjH8jqXfnYaRfsRxwVIc8b
uxXnGadRH9GkCN40N4omTZU+k/CwQ5s9b8naeRTtICchqr0+lUVcYeO/IxwEpFdh
F7DIeu28ogmg1VR2bjgfkOB450YbMua4tK+qbkPs69WeBj1CxrLHerXza+vYsID5
GcTeFbsPsNBBIm7OYtY2r13pYgKtHUTRJdHfPdGUVPU4fHOSxa31l0qAP2LZcAcy
NuN6o05nSmUMXke5IQizvjW7l5GPz7dSJA/Q1eLF8x+vSoRe/thcHcwh9319iJSl
MASm65kP5G9aTCeNfHbfr0t7s2cK+MPtwQvymYTZcEzbk7hns579ojs7Qob1a86z
FZXJVMGySR5bwR6YJ5YUcVn/MMHQ3NVnm9BKanfAcrJ1CdyZkCyJBSazRV1ze521
wskZBUqRl26uQ60/hOQGXZe5NSuQdc9tfn4BJuOzatc6gEwPLWD58wz/8ttfclUI
YU8TUV1/4LwGXxIwqd3G3zOKrFZrjwv+zFrHsNNBMAqhqKvSyKSZoMTCRzob20xp
thso7fklVLhaSfvxWZ6iQbvrXq2ZKFAIaqjUuizSeG/SnyRHTx7NQzFEWyGOsFfx
l/QxRabgRaG0yrdZf1XYLsCVwVL8YN9YThCbzFYtIDZTnYYwHTM5JTLq2R4NLiwe
uQEukAimbGKPlz2edP3FMozEgmeeUT5XqV865ivPwNi9QsP1bHGmwm7B7MOHcw4R
fNK4p1xtkpTz0KV/HiB4MKUgVsuj/WQHtoElagWsLk3MzqHLL3IvL8xY5+LG5I63
pinu9eb9pcp5SpzvnRIADtovBDXxLuuHpQhI0W7R46fJsXOl7L0Up3gXUgUU4T26
X2rPFpHYQHbnjAVpWI+exQHZBNhHfKKZ3MM8gfWTm0Pgrg0oS/VQUCL0hVI8x8AM
MRV6rbrY5HlkKz82zym0QIzWRfmdYXbxnnyVVDKK+ZDxh3MeH1mwdn9tvbmq3Cb4
lYGcuUFhOeSeh+dBOI+9+ZWXcUqEOmC9r8tu9bQbQJ4Rt2LveYSfM0jFkA3+3W4I
j+CQ0RtnRGiZNKJHFBDXpSgEWvN5BSPRRPnmKGpkK2IAuwFwSCLmgyqtUdh7n9Ou
Glqt3FrFO84p7Bmwxx1Ra3sXEh/skCViNjQ7ZqONILJlmbtY06SjKzDb1yZRntF1
Mt8YxEGGRHb3R35gLTi3c4jE8Az111nIHHjokoNS9+YJG5YBbjo4/I/hTs9Ew43W
y/FGvgEGZ3kqbgfenIHhA/I7q/B1VS6Ij+JzwcDuGyMeRgITHTySggZVaxFzpW2G
qI8iLAflqd+vR8mwSKMfSLShs9hnDYK0D8Ickg/3OUVerQpo9O0NTbWebv4ut/gV
u+0d5LUDTdcKMHth5eaUWaMG4/8tLf6kzInqQJ8XJh4+vXMnHO/qrKtqMqjhDgmP
nL/qMwKFhxPJHdb6qHz2kNOOc7P5iTGOyg5euwJmgS/udAcMAYP3uvSptztCvIYq
KrwmvwewkndxSW6Zs0M2o1fmTvEWYkUhWSyGSPh/MNhbH0nq/zad4TKEKoeroBjL
LBzOrrktAwvB4kWV/96Osm210f+ks+OXrcefa5SwXzumV4feXoVqEhNRi5XwfiHu
fl6zO3G/Gh37yrEOLKbDBMEuA8xTTBZxh0t8w/2A6+Gtl58sGWQr2bUHTUlND3Yk
eiH2CfzzPe5qRaP7q34a9SEjvciMCg+iOwUK8cTdWYPmcq8HUoGaVflsPphuGU6o
EGnILPhuPZIcj9rkNn8U4oP5p4HiHgUI0VP4m1xPCXnmn6uGejJJyINtx5yjZ+HD
KswLYuyqrCV2FHIdGyMn1KhUdiQmzG7nKopWZQjnYyLKTOr+h88AABOREoMSMcig
RXkew8jX7Hz8WFf2eUQ3Yb2N9ygB7JsBqWXVGXEFMXsvRNzBGpeazvR5iRzYq0gU
AG01l40FKQiSwC0EOp1jMwIWg7A/WQF0g/dv+Tw30xxTjwISHpc7tARxjar+u2Az
U/ViVgqN7sObqG5glnzJt9Iy+9vpBoRIUt1qi+e9HpJtRetNnv+FwGGoeKrhJTgN
P52lEBHagXkNtNAlL/ijmeMtGQb0skLCE3GIIiV8PpfEQHGO3xwKAo3cvbTzwKBV
icjhHyr1p3pFAH5e0fKfAzLp3WepfYJwlpvIhOUVsKPh87FvrE1SAZ7K7ILEshpu
efRAbniF5Crny4sWU69OUcvZInR8Ciy9EEADwuCNGoRNO3TVUrP9730DdR1SiJeo
nEG67h0acg34VnM8fbXLKSyFhpa2gss+SPY7LvxSHEqJvSK3rAj4Ib/FDh1YxRD1
YAlIsk6LpG6vXlLZBpOfS1TXKDNGuWz9J7HtbiyTkQhCGKv6zE63IOjJltM1FZbA
xlpX9mcGGgmM8tvTC4KOf85GmIszQVv1pAyGnR2NSkBXZSPnPc3bBVBzqnX66U+G
hFl2WKMWsGLUm1T3XWt4NagLifs1JX4rT8QVZ8xNH4FYVWkgbsW2UYZ/K1x7rz74
7SlWXBC8Y3RAR0/kdSsCaTwgC/vanNq0d7M7N3uo6J4GSNTMhSnTnNEldmqDw5AW
q24ifhFE9ABUEAM586LALmTrIB+ULLps4HuykLPcwTl0NuNyZlaRszpiSWalCG68
07F0RxHFtbJvk/QhxT6ukoyacbBSFQSC5NYTZ0JFDL/JmO3Kxn+F8OrjIFK+SUsM
+3UKEQdXA2+G2oh0H2MmJ/FjUx5Yw0lgSOL4fwHPowMQnioJclCEXW8bxmaCV3xv
MRH9pZ485jbb/CjMsk74vXVRuiXfblRydyR1CNaaLpTfI2xoClnzDq8OZI8n6VHl
JhPbdH5C1zurDFBcLIWx+AUMzcgrpCQCTrBQ0nf+kfwDX4tmV4euC1Jx3UWS3dro
3spWMLMNK2Hoj5YY2d7U9BnC3mdc1LLAGwJlHqcH04unFkZ0sbpB7sdkMs6xdoH1
LNxNV8Pf/3TYvG7yH5y/8546Hz+b242xukuwfOzM5X0Xk7nkgGCqxmyeR84z7oB5
dr2zcc0++xvpts2wYKjiJRRVHHLslQ/XhAHqj45cTvs0kt3jpgWimhGkQPfHvTu+
jBsEdbHro/x3IpMYCPKZhmrIPzgac29xDnd0CM+YIZz9e+Il9uSCA8jrmcCt2+UY
q5f9Q6pZ2ld96N9GgSZLqeFlDIIHKuRSjSEP4jr+vilFWc/XmAA/KvuLXVVXzEjg
gKMfIet89TD+f7wmCK+n3dNYjZce2S8aDknUxcAwr8k7QSXtGA9W7T/aQvVMA7Qc
0bGDHiwUfFlB2vvJF2PwBFwnCcy/2pqnACbAVxVYJ6QFG1FXtO1gltVEMPdpn0RO
CoAJtyldRZY+H4XHOiOnUQ1GFZitvJibIx0wJ2Pb6f7pJ1JXrs7nRqKcHHuko+SE
yvDAvLUH4HtGKJDTsMbUp6Lv3MkoId+NlIy8m749fLKTAcf/R5IUH4CYPspVHJ4N
kTVSlP1uaxhO1zKi03UBOrDX8PsTplzLtVq11bzQ2WcsiHeNZXlJ2AP++P8TcGKh
N7vsbkMo8bZN4mgaXDcf+vVt4pfmc0YFfatvG4kqESzUnfPQJe/s+33HjamSe5Oy
t7HueLtI3HJYsLRNy+lDgKBzs1tloRl/cp+Dff7Oa0eTRxwWtn1pMNJfq2LwpYph
s2CcLDOzSsH4GAf6Xtp9r1eNjqnQ23WUnaXfF1GS02pJUgoxVP9eytJ/6j/V1txA
xRDgjFifMt0qyZGKqviQW6/i/DXINGORaOb5GTqyEs5OMFf9n1UH4BqMrw4Opxk3
MtUm0YDYuEfItP35C0ou028qnOBqaZpT9Mll6xBH8assWuTbdBD333UKmQsAOkVr
HJ6i8Qnj9g8Amuf6Lmc0Y90QxEaUsSEyBYtx80izWUnNiXENRbmSpWLmeS9R6ZcP
TO8FXsGwFfey2wDMxgHrppYZS6xMFYLAMZUczulknTprr6FLs+c7ZaZ7kqce6rLD
3GJXlDLlL36GV73UucNFLoqtxa/kRm05upt0U/bev4OKDW2jLBgSOqNwekoymoDN
ezaYJqjlnfVIXUh846suGK0kFfEo4/20ZBwh0FHhTFWxWiwpx/cQYGkW2hMWCyGq
9cSMspKc2u3OdX2GixilkFhuKvkfw78SBNawimq6dERqdqde885JcTjM6bXKhsLf
KD7G/wMagMEzupYxwg/sPmRZPn8xodJew8uBCCbYBjJtZfpp/uVUoNBr0pGbdfip
K9EE4vjGPMMzh1/CNv02BavUNzBXmZQQJ9MTwXAPrcZPoHByI2xCR4cxA4X+0Gfn
1Y4QN+d4afiM8bplU9F9N2+akk6E6tsLJtDliDLArXt1qgLIfUE87PRg5s0tn2rA
FA6WutL3+5cFKRms1hE/PNs+twbDa/zjlsxg3lLvJx/YnFyjo7poUu/9rbMyEk/s
rNCAn4hRA03asSYN//S+X0KTVIDaASLJ8/eXJrNpgTl3BCihu9ggpJDaO+fjmaRp
GmjftExGpVvdfehdkT08nS4PYCctklcyOQR8/digkrx8aRsVLKADwXU59MkFjTpd
wlH6EIoNUX8TPswSbcQR0Lj+LUG6lplVhfmpcbxTzRe3yyCpes4k/a+qMH9Ubq5f
e/PkY3DBJd8aCopBl2Z6c/Zw4tMl5IdkpdMXlqEzeplRXcVUaDWkfHQ0w3xDo95h
3qM/ej5xmGawUee+UxtqGvmCMUzYtNynyaD5f7L+MC/Cbqd5+qeVEGk4k54wG/QN
Wo2E16qIgsJN+xiI5r5T60yqeyuqqvrXpeMTr8D2n9rmeV/xP1cioJuFUQZOpwOl
9ykWnriH7wLT5eZ26ZzrfE5asCVtzzWjFu+Cx2tcZAje3Tz8fB8dmWrXZgjlHlfN
ayCQZhH7jtRRW9EzHZyxV+mNEum9uFncG7ZkF36fcntGetwjt9+sguFVUJsU8dxi
VW1lxdXd1O7og4ooqhJO84etjNOi8+bd/0WYwmOurjfTLjQ9HLwISJIcbFb7m6gv
5DIEhR+//D0mFF6Y4cy2nOvnPpe0e7MEGD/KaU5q9mMzsF2Ly2styZWz1JWXX0fz
hUgwSxRQUdMGnDqUpAzQCyLEYkgQhPy8h/goITGJ3O5lTtmxa3mlifyfBN0iXg9w
kYMaC+LYTwjlPYs68r2dhJmkNefmaIuUYr/SQaq3ZKZW2wY7r5rZ6Dki0EQOir/x
ZpvtNF9cxXNqgLu/Itez0PVf91jlKBy8VA6F27lMode64i8bRzMOvA+A3ldLoofR
0bjF61PnfbhIUXY6wt5N5mw6EANlN3iDqquyHFfVPPl7JeRqkXQZgSdX6ALfLHUp
2lOxRlwgApao3PxhAroVVEnVBJuUr+WaVbOy2qMaW2FQQItPWBLEmDnHcblBiN1v
QReucsnHCpKC9HuEGHLGsKkBBblqB2M3D2Jd9d3VdjWpPgi7Cz4K1mw55D5z1Laa
lxGJCmnGWpAv02nkz+vpxBLPqCInyQvmKWZciatQW4qbu0OzU13/aNSM/eo7cb+C
3pQBPpA5kIgtI8mPgql0cs8h3eSjXKSnUiRw0xVbTtdDzQjgfjXjwU7DLbAYfawH
/MwpGMgSkceKYEso57Z+hVr8wZQGc8XoUN2gti9mq3Kwwm0HH+/hNMMCUzJfU5n3
ozqeStsIQvvOEVqKbIP0Q3OdanTqE/++lDqjsnY21C09jTZaUUT8HjZf74rvsvji
yHYuzfEmPfh6SSFfZ3SjLPVUtEpRJKrXeoBVSAHqc+gVRons2EJChoIWMOP0Firh
nYTJ1/QJdUK+NG8j3ZQX3hN9mgasxJLT4fUK8t7ZyTJUk4efktDsUzSt4Ztafs96
o86Zuw4GtwW31sCSvmDN1lfOoq+3IPhxrdGLKOPYNj48slsKVK9uiw3zE0M3fyVW
4wHkrKdMVMzHVboqUSvFedEPJ42LlBc1P/nTpx7lDySGdh42AGgoOhJ+5eIpgBHJ
gAcBkq53XfuHixuAu30hhoBvovYX7bvAIF/pLuxCVcrGY/OLEqws2uOgpudhboD7
X2INT30EF6QLdyXLAoBs9lsK4id9dXN9c0u/49um1zktpoRjyBhHC7+WINcWoWuC
m0D2G1B20d51zzTMB18MBjzYcAidp4fVkvHfQsCK2GFpLrISpmpSwFjOuWp1Ev3r
spkPFLuBeZh2/kKfHmKKqyvK5fkkbUHcvusR6Nv3kPQNC2FdjNIknWCUs6o0lnsn
FJAWkr/YzjBBADLxrtLIdh5pbn+sr5BV6oXACJ3De7nvEVx7X1nSMyz5QPFf+IXs
ZE4fLcanoGvJa+7zCF8IPg/YMEnRU1PS7kVqizmBCJqMWsvLo1V/akCcODDVh9UP
leI2xX7G51XlUtky3u2P9vHM7zIFsWsZAM8NCwKzoaLTrV1nNRotU/aW7LBIpO5u
wqZzuqoHZeliE3jxCrhyWUJP+RMD7K8xH/ykC2MAbMRxM7Oiv5XCN0Fs+lLHvW+G
Z5IbC3qY00np45WBx5Mi6lSGEXhBs25Qck9oM6ARs3nG3t2jI1YP5w67auupum73
BkvPQed95mWOA8WFBsl+xFScucC0Ca7VTBssbA31Pow2AgwvoWAFqn2IoQLXkLxJ
O9qNajra1MhLlBVci1hznhVv/mSsFggTNP36e68CWVGBDoT9zf0gRShzmDDS0ugE
qjbwXGyYzj9yC1DxPDB4aX5bkvWX1kW852vbTy/vgbsyverKZ6HuhfFKbG6QnzMJ
xB3fnYrIzv1cfLkyc85fuy5Xu4ShSyQIc6XcUbn7AHUSjw63Lr5SpnQm45k9Q/CF
MwN7G7BfdqbfpJCtZtlvFbJW7viTPgafp1jcEkg+6rpE0Fn4cQgaB7sfb8oN0/DO
IWEagDqEFwicJqO9XnTsdCSmOkm07QSnduRPlKr8O/X4pgqJu4z21H6pCxOvRhcc
Ab3dsvxqW7MxI+2+58/D8IbmsJVJM5vQ71gP+iv2ANG2hl3kdL9UAn/3wcOGyZCr
AgxqH2uBP4n09eBCGrb9fCY4hg4tzPxCZcxMImW+9XxMrhBrLqxydFtem9DAUxcY
XPRPkLm+NnVQqf799jKoypvH3aJk4Nd+x0cY8aG5W/vtCrGLq7950DTKqeXIsVZQ
G1z/heNKNykA3FTdmXMkB+ncsJYfSZcMVQu8GQ6hXhpoUlvrce1c3FAUBq34wEz2
9hwDzAXvXAtr1BTnXPcw6Oj1EvF3gwx2Sw5bEMh3TXGasFZMzEVpJM/fmoGOzqcJ
GJNEB02WLJmOXKBrCRQXkA+IKbp9YxYlindDhyoRzLMoYDIbNj8/FQjqsZ/MSxEn
U5pa/O/Hc2d+yqc8kpSOAOc0R0bxyUgxwPXccNoiUtGyexcVbgVVOrbobTHSOH3E
n/RaNrskIDC5YvyNjpQWJumhZsJKENnwjVgkHndm4PpB6emxmoA2eVMQ5HLOAI78
J9W++5aOs6tinY1J5oVRNcgAXkegCzsf4KVf4tDymcUC8o3Q7oYePKgvezOK+og1
IUsDO3Z4WNbA11PvS+uSMoCA/rihhe6OL12q4kJapMxpJ61Nh8neXdncfsn2n/r8
sPnQ57VvgyYamjb7zXUJMZm0oVBYLgpG382eVLd07Us2v+ZtpJznakI2OQbNLp/Y
xQfYTVzSj4L5tw3oWEaHl8IWaCxEt2QtWwH6yGRoN2nqmV6D8NmV2RzPEFGN829r
o6M5Ic0kSqkHbJdd9yn2EcEDwKtlCo/FDk+GeHxM33Mbr0ldyEGG0JKs57ILmATn
NOHBIp2xNqRmliKyi8DuonYb+h+qG3Iw43Yfg5IXHGirpYP9oR21d3q2BjN0/W84
SnrNikOlEQgKpyANB2Y7ZH7H3c9+SBrvc8nuxgmrFCiGL+2sdpj8GKDtdGCa2Zn9
JEBBNHrxEGuhebwDHnxiw5/Rl39G7bRIKIZmNMlcZBCJ6NgH9W/VmveIAJzaEOwC
DAFGSjzD+yMDLRIeAETDkDxDmRjzX+YzhHzD6X7gikOoQWXL/VAK1hePI/2rt+ut
ZPe8JM8A6kJRT812rTPpICWC767RPp5DBgqCYmzNTSDhcNoh+iaGGixmNomplLr0
sPY+up1gtTHok70lxDYlAphyDhcW+W7YISbwN8eJ3K363tOLPEEuttCW04V8vJFG
I0dQhOztBZEDa6ORUbndH9Kxn85G5j9S01m+iwzoaFHPo1bJ/JTH/gvzIZuAvJrZ
nwUhk/9mIG0SNrdAzMBTMfdCzoTO/xmG0fnuCqMBVmcjU1K8jNqgp2uEfAkQS297
VzOrUKP4E+nWOo2iHTqAtTNSaxy8/Kwmm/tVbQ7ZGetYvUHBx4EXFvFGiXpYrSnl
n4UzG50BsSubCGnfmhffz5AKOFL0FVFRp8Tqm+AfwE7kIMstVj5Q0cDCOdDHJr5R
thsc/CtYkgTtntdTQgL6X8oXaB6rsZVhnkrhcmsR+Q2dfhot1+r1l+cE8wIXnKn6
xCnz2bHhQC5sTqtGjJEa7vHVpjfPwDZd6MOSGloxnKD469eUyEofSwywRMei4Fy7
WYj81NzOD1axGF6sMKpliAfqv0jVJWV/YJiTeyJY6HtZd5zyhbat1BQJDuoRbB21
AAzQzaghEicffl433BkkwTzzZGY/iz0rWzoq/Hsa8RXXo3WxX3zJoNSKLYV1ZhoL
VHlj6rb6zkDzUiRkMjAcvktGArOJWSsUbqtigHWf4V5+0QJNOQIMDaGDMoph1VQg
og7p09OLUAjKSn6vL5YSSktWTFnrDgOuoNkh62IyQNNtZw02FqPqTWcEqoXeYzF4
FV8A7NOQZ94rixTKY2HwvdgQHe1vt+COVU971dCCvtUjQCGmVNAmqpXi8oCd+bWZ
hYNzZaCGPHkjpv9LQ2l4AO5anQ8550yYgsRukiIenM01ko0T5lNd50cLzsIeDSLN
jjACP6OmF9gBFa8nYy0/UuIUMxmVV1uX4gZVLxxZMivSSu3E7w9nuL3uHaoYCLkO
j2l+Y7EGeZqUTBcedaEMnwjBrwpo5rXmy3t5iUxdxMrbPrfSMZ5ric8vjGk+qsjj
VqdywI5ms8IrcOS/JJnWNu02fkP3MoBl3gwoMivfzNt2Ruvkd7nA4ry++eNYApcP
EIT60W8tZivjElPcgglIIB0QWWamDkenVALh9hWwBAWvlfTK02+q60hMTuIMQ0Yb
BUxA1VYaNjPa+ZE6U/OwOdDUxLLjhIWF8uyPy+7NVuwLKkf+vTa/8kLar5/FnYjo
emTROaIsIZKWbo1LrxXrQ37FYKxGCmxLIzV3R3BpObMuWiSeZ2JqtL4JD6kdA/Up
L8ugh3Y/TSlTimDWjtQmq6pC/LrdFdpamHcshvCH6WrdqPLBR7rJ0PHct4pyBMXT
UYorj0MuhhGzXAm2D1Us7/9s7iC2Mbg9lPEO23wwt5rGmjsSbmhOisr/duYJe7Lb
PXKsj8ZB+NnIMy1ogYmCKbmJY27LZuMPtj2WU7WCiGbtpdf8tAR38d6PvjRrV5qX
A5/oyTtbufJ4YkfYThOPelJr5UZijki5cc2yaGaQ2ca1Wk+a6uRHC3THgeSRA5hs
aUSrHh+U0gehXH/GAOHSI+YKlBrfXLXlJSEvlexC8cq2TvP3f7hA7iB6MKMi/6ur
7hW4MNeCj0k4YPNT4EdO1yHiXsAVMV08fCYGkyZnenewhTOn2UjmnbrFCK8ZEZ2L
Xr/qoXPINagTThgve1zi+KrIY/qnpdcR4LRvTLQPGeOzto3UVuIEPO+I0o2y+ozV
swmzymGDs13PUPvBPi7B4PfMB1Jkj7aNck3zA7gJBRDftJwYoPPmfOtCwcmnOeQn
euvjZXl0RE3isOf1jlfLD9vu2qnFKgSCMWjOTzPEsSyGSfKw5DdWn3omVJcFnjJM
NQw+8JQajr/QKDL9/7CNoJ3gBBIvauJQcPFITY8qbLIEiIY1t7wx3r5gpv3m40fw
jMwPa0s3YWAUnhWhsxepNtEWWiBLWcjqw1KJSXss5Le3B35XLGG1r6R+Wkc5hD3y
zqKl55EAiHDI9Tv5mh/k/59uwOKMGGUZjEYidN/257jh5TRfTIkqzYjjLmwsNACV
83f46qo5H+LbmqjEz05GUF/k1PEUqsRHigA1Rv9Lt+CYWHvIt5rdLFheG/OFJYzW
rCcu9qLdZmU6CU/JbQDz5sPCeaIXIWCqfyeCF8tk8LEvP0ARANsb16BP2Fr2bAjU
XT9+UmVC++uz7ACvohcAs6xaVCxQrHDFNyYeNhEUHGTqO2KDfE+tbPH8riTv+ZK8
Upfl8wvMXnRczfaU+CBI4jy/5TJlnOZFfq1JmvkTSYI4ADg6MXMQjKFOpsywnyRu
3dZIRVsKTaVaKic3Zt72IVVHSHgnhl/eVPqTVoABlEYQNIo+s5ehNHEsAXF0NB3q
MCnLBjXUoDVzzgWeRJwbav3gudAD6YRD1NuImEViOHBk6bUKKF4IIQJuAmxJUNBX
I5UCw4fJwkx53YAcEU8hmSANCaV5ylBuAnmjdXaUbJBTLcqcMTBLargdY9OjGycT
xqcVWbWQcni7ILGel1JBbQLBuoYtnTmQUJ8B2Pq6iH/A5dZcAdFONUlXKA1+FTRy
d5avekcNaKX3PLkTFg1AO1e7iKOZLscQpz2sLuuaSEdj3rM7Y0CYe58v9f5VC+Dz
ky9C4j33yIH/6HkJ7caGX/aX5oiLenqDkX6b8lhLo288Wg6OZSZusV1oiOWPqb3v
OEQb1tGHn80nkXsgysEJYw2VoWb9sn+0warhD3wIdZMvU2s7/l4QMimj51eKScQ2
cIqaiB7Ixw+QRCEsiWXNHnH2IzkWTriBV8wa6aiQe3sQ1rJgTJBJH1kkTxchwezf
0zOcbVx+9Oqah3fpLIowtoamD2hGVe2JyBsi0lCqxV4uaHRZP3NGlShwOnT6DZeq
9xRmzPnGzcYgOsCFdZqHrmm6YkMqLm46oQ3njvQDbaTuSkLlOfTQt/5eLRu1scQ9
LokIyzt9vxef3TfvPsFnSuQlHU8jwdYcTH/Q1BEjxDJ76zimm/B0vOoRfWNnr/DG
QMLssRWjozKyvQ1NeihhT5WD1lyNyhQ17/skL9D3c9gdysDO2uEEE49p7TMz0SSw
wUW1XLGF7FlbzcLDzfzRbXj1wxMmM1PmxZEwpT27FWoitpvpVy0Ca3DWXTyV6Sih
DoQC8oTjoOlzM3ll0Gac8emvt3LXiEuP5lK4wWH8XEZMN1JJr6l2borsbpDJgErZ
Y1JNeZUluACrBDMRmuGEdHNeG5d+qbrDdMZZsxbjo8+ixf3rgYSr8jdZzC2Xcq3T
F/hx8+t8pjVYhPTiKLBLpeAFsroulR4GF3odNyQBgjuUtHa2SP4nCtf0/qFLgnQK
vHtVhUCmlMk+VSvNqq6JQbHhY+LIdXy19R8X0qZIy0jj3ib48ClQL6nqhnCscc3T
UJvpcW3nGxdP5/99ifdpn3TT8CsDSjgI1SFCKiYhSim6M5VPo77/2VsIWE8X055/
QOS1AmP+NMv8/9EbOtDWwFat5yNn5Rlic3OiN9qtTAEihEBOroHSipl6ajRLSl2Z
sbplvi5eKh3iStnOUwrFsvKItNf59H7AUxzwswEmwYk/FckDErO3DIIpQe110KGd
7bC7ClhKejxmEduxytxLgOpLYjcN7gsBREKSxB+YtlTOHhRJlaNpCONerZYx1l9g
To0pK7yn9YVlYueLUk6xI4ochy+wKLeO7Y5/LJYzuPvTLvt2lF5EXmYiHYHcOUEv
OYS0NGhO0G7t0bW2fNpYImVr2QPr4bgrnyWbyqzPJGSFW5rtFLWbeLJYWctOd8/2
uwqdA5ry1cvhWksFqmXgoPhXrWrax6Db/Vw/YM8scjjEVLTyTc8tYW3ujmGsj+fi
VITDFFPwbJB7HB6FPL1ZSZMoP1TUAol6S+QzJTlKY1EYqBDTt9yViIiSU5TyT18I
IpcdiQY3VTjhAAjJ0m2q1prnQ1uXLgLnb2f7VulUNvXpn1902ErOIcLXZATCopyW
U5rvSrZTUjz8OkUyCYi2gPrG088sKAJ6JiguhX4LG0HSDM3ne6UXxabDG0P403YR
s6o5+1tesbgp0McwR4M7/wZv7CVy+hBE46ziDnH4wEwojin/8Y4I+vaA1rd4OHrJ
HR3bHU5XS70z0WAspSqR9CwOVdptSe8QXi2dqdGXYQTEEA3cjlXCruwvc6TuC1Bf
1OkCA/MBJAz3i8OAyMfSXRqvpwmlSb6CNmFsraw5wBLDkCvk9d6RHz89z6fGO1QU
N0HwOxY/6uASZCvZ6YabRo2otwheUt+2oZ6UwgxhVXK1Nsktnje3mQOOOLUBcjXs
+k2qxrnACgNd3RX9OumnVuDKPwWzpAOxzMKtw8Uzfq2hfNCUV5d0T4F1io8xcCSB
s/57Q+f/1/af5S8WaLsl07qa6Yg0Z8wfe8YOTAaxqJVClOLv1eIjYBaaAO+qpdjb
peA0VYr4i+/RkDKTPGL8uNeHyVC4eMx0WC2ydtYslXqOTrJekex9421Mjxd4kO6A
3ZOVZo0h4tJU62qgHt3YmtY4iPSFoA9kshA09eN9imQyZREKq9jTLV8TI73Ah/3u
1hRr8KwtrExgzwBXoYRkDJ1/qjFpXbLs1NZPGwc/7suEfkiMoXbzPwST2p/LSlBz
aoQyyltvn2HVP1+Krr7AMjZxGPI//n2/khq92amzr3MLH0OzEnHBtayovoma/zNI
bAs1tL1uPZHFuvegR8FeAOwgIvOetbnxDbgH4xXT8Cc9nlLBxmC9Io4N+vozzGQg
iHuRRLPTCIBh241L2+TisILrneTMTG5w+tuuB87aaZMw10sSk/iKxobWPF3zbfVR
xik/IN2leSpCnmAUpbjlnU25NBVGJbfNH19rHMIZ3FkNdWD/NuWXFX6lzgsIkQ+U
tzoHJjX574aCGKBWUIGdVMgmYc0UF7Z5tKdX/z8rHplONV22JBtGNv7s8Izzl43k
Mj244m2ggY/zRvCVs1CAK9hq19MCMrQ93KWKNgS5m+HOPDiKQrZZLEiBkZDzYybN
fVukA7P8vBY7MSoYSzkH1BsxGVOkaL7HFPLgfy2rEJGRrL2rI8dznryV/0V2nr4J
Th9GKxiW9itK/B+weQN6vU70VVWpUjd05UEeuRca/22v1ih73ILkBU1O33aQ16/T
G8zXh6G24wJLq5H5iDCslZLEb9NloN6+P5sBPyOFV9ePPg/q9pA2jvL6uGowGj/r
XZVXjffCdO4Zb1ETz1ErNypoxK/IzHxvs7cl+Si9iN6Ft8F8MtNPGbGCalObTtQa
xvXdU0KwJ8kI6NzLNedZfbOBIpIe7zEGSXETnqM3trQCB/9Eim3rp1VCjp9ffbYh
QME6//iXNz6Ww9ne/8r4vGlO3fK5GasYFsAT7Joc4q0lonN24ywEHHtrwydQ/ZCq
fL7usmjANFl6rSNRQPsfFLUKddwVcsCvZ51twwCvqwwhCvD1QtHvXXHzVFk6Ulq5
CFCAaXrMNGhITFy8cmvOsVlFTAgNeFLF8VEh2+Eig2VCI2Vlcg/wiR3Idc2WJW6y
xfdjwXN9nHEa6XrEgM7tBtSj2RdFdpVK8TngVGGfuY/F+UzV/ZTm7HW8Q/5jEIf3
D7LFyEe/dU6Q5kH0dOrcr2HI0RRy+Rd2fOY35orMoMqVK8YIEefO+msSErYdR0oO
Kjed9XJz674O6UYykuPw3FlBqZUkjSXGhm/uJBDMkEgmf1z+njgpMH1cq7mUOe1m
pUBlmPxGOBzhGOd9Ej/WsTYMegYtXfxMyjZ3VJk4/gssXN9/i6ZSakOZYF8z2wEO
rN9uWKCMNyaFQpSRd93A91GGmCuKp9vTH44rd+6FHR43sUIpSt1gC15bIKRHZJ3e
AkxH/wmELwW8LtT9Pe/gJV5bWcpPG4Cn4167NM2ASzIk/xmaWGt959yIzyX+A//g
wxRWCmxR+iSxiNDVePvAgS1femZdiuGLbZ2JkAsyjuw2NG1T4Z6on45lxTWzEYIQ
7lEYrEtuLtLYYQC5A+MUAy9PlRR1/cyfw2OKdrlmpiUf3xrQd+gsWiFxcnPZzGRQ
o1tRRHkm2KY2gXdCIV5RmSSk3UKcmKj7gmmIDxYMv8RYVlGqakqoPNTWbiYKMU9/
96/fAQwoYxAzfwFxJnb2AUFc1FGf3AMSOhLx8wWFsJ73MKA5sY6Y2/y9KdpLliYx
W1BkFTKyxgwkMhvebB2V0YMyS4mC4HncyFMz5N0KPk0/jvN8uoUOligGTXrvg7En
wFDhVSs9vgL/ur9rG3ri32o8t5SCPMpb6htrC9KepOptleobYE7V8xuahfEn/qoE
H7wPv+vYvWVMl9/cijEGBTk2YlzAoNHejn/jh4NN5xvQger8e0IaibDJaNKHT8nG
mqo6x8cmsL1TIDCClZxnZ6rkPL/3UunncbxDEwky7jFMg1+EQm/7XaopbE55MSlg
vI+BWWOKrJ5VPpzg0OwdM64TuTWfPRO3zUSLIkIo8Ok1x4FTcATIjPNzvj6ObuDw
wKEVC/wV7dpQTQFXpW2EyfddjRrV7Bfp+mw6jHZI5T1S8jIdIAsjh0erbM0g2X7N
s3KJTiuM+iHKTScHxLKx5KnIwRVjS1zk5hCnHiyFbX/EMTerbzhW8JURyngDvrGk
lq3xxmoFwq4fvmc2NuJknWu75hrTQeAxTjyEG7jJQjlvdq6phkbp+q3QrshG3IVf
ULdFPbhkYzADwitheuptm5xyHa12cPvazU66nfExvaRy4oKW451e4ilKYAYctwj1
/E7b5yJDr1Rw+KxxMtHg490eWDCLRIKLzTeONIdxaWzZ2cDiK4ziJCMvN5gdmGx9
neIrl1PaC8WkjMAKzJEzBPBgJAI6rubEpHfR+yKbZ8PSDWXTvLiknCmphVs4kKkB
ekpLIFpUcjgy9120oQQxgdd74mJ6lEla2UZHmZnYobcn0avyUIYnRKCd25NRQSos
wUKh4KzRr9DViSgL8A+SdXMo53V/x8JhJtkhtYRwQzp8kRglFikCdN97NGRRvPH1
T51UXRhqwhDaxw3IJIHah5eRhahDzSDLd++Y/qAnUZ2dO/QyLhhLyQxR0b67qTsv
Wo3A/Xr4VYTUQv0wDp5sPdWqKePgwpzfesmi5j80ni2EEPCC1GBM6LfXIz8Owpw3
R9i0zg/QBcAIMKPXr2O+IGxL8trYbhrXWpaNSxpaszqAcgJoZm5KhzQhZqf7grJf
XfZ7S43tSTehYYzJtnmMLGLg4Cf3MaEGXcJlLIXQXwlJOFPF6gVybgXN1WgE6hsm
tNWoO5QnVrVlscKH9YPILViNSJUfozFcBv17JqYBZ5oUUo9stoh2CUSNXzvV6Xtn
oYsyq2hMKHu3iucnWzR5QFNJ9xBw2SZvuzqmC4GQklN1UTudW5yzhlJMZZijKF9V
vgQqVvC20x+X0JgzV6/BODRy2uKGqQ1FGULi++FXT6ocAZ81BOWUBgGG9y5EiG+O
nHU/6uNTrnj/gJiWNQDhHVBf58ZGfZqt+U0/b/YNTwqffeDaeWI2gpkcVjiLOCXz
gCJBUSevC3vuSaxtRZqQGHuHXc5C7FnkuBr6zCOrVhqFs6Kd014zxhV09DKrNxV4
8iaGyM7KoGoLLhmV6/sWidGwup9lYQ0Joe0vKB2gn9JTh2Yp5Cm48OzWzN4dBVOX
v/ba8OORkr+aY+vzTuTna40jSdGVXvqT23aR0WQOiz7YS2B6d2NOw0wl8qSe4TDd
Gar9rjg9naiE+SdRZ3MpBapu81rzyfLOGtNeCmJGY1IM2oZ4mkr9CKruK/51Y7R0
5BYTJg8NMPj5/UVPH7aHy49jY6f2NSTV+wsQQrU8cXUSaoYFe5rx+rmPfIHJXNjj
6fARhxjJJX/6CPPcAQer2cKWH/XZ9PoYI5hBYDuD8LWfr6CXNOqBZZqHhGKw/Hv1
HXx1u0kYCUrtgranfACeKk2GvG7/rV+TOJnsRN+nIztl2uz7dtzhL1ykVyYfgMgM
C+b9zzeRUZ+q3PcTmZt60Z2HiV2EZzlI/sIKK+SV5Ce9rhBhko5G+Qcki2hzNlj+
rXruESAB6Zw9OaY6tBRVAKDfTtAJJcHjUdKrizxce4fl7YGpBpMdy/KhzQvTU56h
1ERgEu9S8Yx+S9rrx2P5L49Jz5uYmK0fIknOvV9L9IyaR6GwKIqEEVztKgRhy36W
bYp7zy34Z3GzRtSCioCr1fYyBMfdjADRlEndTkmsTtwNJrLqDJwiVQLxoXi1IWkS
sY/+piF2jPVPZqmqZHDKHqHKXDp9fYIasP0TohtHyMG/w36FI7LvQG7WFJqDGkfi
0tx/3jEJ4RosmV8MTSkjuo3DPmLND27wJoWXStQRotso+me54F1Erj9xd6VIzfCt
3eQ/v5q2DThQJorO3eIFcr0VojFlsXHlgt6lXZCL7waCOntSSS1kPVBmAJXSQ/L+
cfqc9LT5sOxiHmU0YBHUM+MKC0sXaEXzNyX4nLWuTPDQBZt02gJyvAwPfoTIGegR
5ytkKSviWlAj6hlpf/PJzBqAODbHPnviLdQQOfTjt8+hC1BN5e0ZcqQe8H0NwkCx
Ro0oZ6rmB1D0Z5ofBYIlxMERmjxIhC9juusQ3vZX4+0XcP7ZIYIOsorXmxvZgXy5
x2NsKaTFgs07R6X1MlwREvIRE4zUMettE7CEZ0E8FqozzYxQfWSAoAVJ4GfxLaEH
P0E0uwFm1XziYq727osRzLq4Br5OKEmSHKJp3N3fSMBzq6U3md9YF1JERo1w1wk7
Vk6huYIf02PUaXGxRpFUeH/pFU8ySsRnTL7aniGK3L7osankJBDBtxXASFdDR3g1
jHCtUbCaVG3ieVOwVfcY/qh3sw939B/zIw0MXGxaBVel0zdwpNbKpzYGQf38ShNL
i5IHYffQm6QuI4BAw/cFaWiQlCdJ3vXEiC/afDRO86tFOXzSHidbuzIdZ7D1ziLr
fx+nN/z3Hn5+FpQOTKQqUa8JBGNp+Mixzrquyc1UTFrEoORdkOA02CCbe5WBruF0
ULgu2wblzY1Jeqpe7Xzp0kbRQBh76qmvcxUTgA9Sj7TJELGdYSMO+8s8rC4NEYE4
NX00YrZkgnw5s2lmrDCbkTSKFKyL8qWO/CCYeWPOw4wDVMz+YiRoXUESsTse25Xs
CxXttLrQS8/++hEfzSuRITMPej0e4ET+DA6oNOeZ2eo7TAjnPCCUQSBUo5V1oSKD
HKkihGPjr0wTlH4Oc1N48YDSCkNdIyn9LL/5m8JZgT9hmemxHOVGb6MuxR7/ehnq
4WNcnzPYm+6AnSWk0tTiu5mkj4kKl4d1Xbz5zQs8y81tOLseOBrcv2FyBagcEkkD
jttLq3f52lLYDTMjnwl35gTdJAIeL1YdItHRXrM3O8SIQtOw6rrZBKRZ9lFIs74F
Fvs0TkA2N3wBG1MCE98UtBBjeeYHR7Jr7cnnTp1vdBDvum/ilkBPPRTYtmpXFNhM
+j/RzZmZ8DQjMvrmX8Okh++8hA7eesK6tLuXmV/78+f5IOgbJ6FtfJD7ErWxU2Y+
LEMJCVeHNmSSNTNvol19diB+YRTQW1eziNcaCZ15hzrx6fcpbWavqE/+foDCL6iV
tssz8tR0JjuwtUjrTDw2DgYrMiUUCSOJPbWXLKNU3CT385rujLsmLbxDBEY8qX6l
vDZQ10Mk7uYFu9hMEyxKAMXKuo/EGcMF2xMq/EK9D/TPFeNaf5GJWY3rEf+1mxBY
+LXFvum3qYQtRF14cwh+TAGKUMQHDeXuSSchOQb9rxYtLSL9ixNrlxt6mC1318Tw
idf4yZM4niriNPNUJToVWiKlmESRcAOrRPhCAeoNBxrZaA04Mqv5e/3xFqB/LjlH
0a3eaQAS+rSt6PtyigM/Zpffmm0kPJ/d9ACOGjP3V2YAl+qITS253TzBbbDQRJlE
6ZwO/LRmHKQNopFM39wBUKUuyyJifj1ME5TghN35tiJdp4DoqLnydHsXCzz/R7qx
NCq+mCkKX7yCUjeaowLk74iUONXKYq65nq3EQdiUaQ7KKNLnTjhTHyHYpJtjICH+
eeSIhqMcNCbJwQIY1QBUsX/6fbYITZtvCzavKy1Afs0Fw1Fkh01+Ja87aTNqTZb3
QhEJZd9UKODjlJYgiUuCPMQaYRX5sAa6o8P2z5pcCw0SAArN0v1HqBbwmSbUGpc6
X8ap2T3WUvCxOySard6DJK3JVR3eiCM/0jJMaKpCMEtUaSF2y5X0ifRjXIDK/FlW
KcaHMrX5X5UvZfXzXy2WeX1MlBBCSFSf5eRiUhZsY0ZXje8xVybFOFKMrVA4a01b
WLECvVAchYbugkZ3pDkoU9RA2PL/+A24/v7MBCAd4Oh+HzC2GV6+8W7ug/prYXpt
moMXtsTWxzq6cWENbi8zMKLNDX0nlfQPufcFb8KGs2jkmcDbxF5C3YmTV+v5Tif7
VMy6D+8LDSh1CA0ACoGkvYJQHxgUrzLO8BHAsZCXwDnbGoDtCfy+auOpl5jeRSJt
pwRkzWbVKgPZoADxSAV4l/zYdPBdXAb77Fx0aIlGMW/OV+7iwCThPNN9yMIgq1JC
PrtaKIiZLUimFZjGN/FWaKvNpSUiLqRg8u9CZpBF6EdhM8LYhaCyv4v8LRDN9DJu
eM+6vKrBe2epHWAxSiVcLY+8WvK1Ql0xbQcJ1kgAoaZDrDl/4geesS/+ArKeuuGo
/XmCrORnOV4WvNdI9wtV3aE2Uh10i9kbnSFqYbi8M2KFgyzY1fg435NGnH6ZnPr8
Z7NGsdtfqDNhEPiM1Ifyf13HG9uMovoOyOd1YNMP4QYn1FvWFSI4ObmaFBCgCbHu
QnZz0sczpzxpfzp/W2eQdaxkQutSV/wIZgN/GHuycFhuDryFzry68sXLsksNicQ4
FWa0qgOcKe4sOqHfHvArCRYq4ZOnCanHwiFlW4jMSezBMa7uN+O+HSxw0JDrma+8
rxOhu5uI69BsGVxQThylPJnwh6mS4w3HERRzZjze7rqQUGc5mDqRHGVZdIGEQRdm
yOjROW7K22ecReOH3gYO4igbdRNGL8yVZyJPX0REpNTW19WcFf0nuwYeABG6eWk2
xmplbkz49IfJcy4/i44cpALN1KvAlfkd1wthg4E+U12J/B8DkZkS6JKAB4Nbkacu
dod50hhycTOHIpi7N4hliubzOnnMcfyYTn/RU1iQWFrNwN2yeG2y7qIKkriDBFGt
8SiaCJBzcpsTDzCosCrqmSb/s0RtwD6eSiB/RWZXMSzH+nMbXdGLUZ6GRGagtzda
SW2aqA+Sb+tr9prH5KbLUvRHjirTDE1EEKlABXTOal4LC3USByMBc0W0/7p5DCS3
kETFn6kr+xn5AzOmRUl4vmp1EXQJKbbEYmO+/QGuO6ZlhEeWnybkQd/X2xYBV5oL
wzzCNwULHBDD6OlYVIZKHooEOxSqAcPTUzxQGVwNeWv+ZuJ/ZMQfmlk2Ljh0PtPQ
Zi5B/o/CwxtNdaYKAfzF13uHZIhW7rPnb9lYqDalm9cmBRwXAJXqJYQgybpLqiZX
Vmp4Z+fCB7RH3/V77qZ+o72TROBQxcE1FGBoK/JuV0hwhJGeuSvVWWaHJHTQOX/M
JdCuBEgG7hGin+iyWU2qpEso57EtxCaIDeBDEy0C+LloTK0MZs9Egninj5gC77Vo
DKb+Xvfy9LvjIG4wU2cNCmxp+OoLeADG2ZhEq61sS6luDPPZf7FmJmY2GI/Fasf3
XKYWnpXVrNhDbu76sU9HiPWFNCRzjwXx2eC3/V5pquIMA7qAQgMMWqXATKECZkgJ
7WABbDnsH8lUWQ6Gga94PkJB+uz3wKpMVVbK/NBhJDG/z+y1Bk7wWhxTwCqDOtv6
ULRcuMkXwx1Vwly92hTAZQdOEqo3/7vlDzF/tfPQ4al7kLBlJxct3YfBYcO+Afv6
7p7Rz/copTNvGf7bGGDGVuR8/XOlD/OH6VYWr98lmRukqBQ5wuUPJYjoSgPiHzFM
2u29atvT4XbFyHOdfIuI1NLfSqvopzlYEe+KDBe6kOWC91Y6PGnX4XCoMIDB2Ubh
xC0EwfQJKbLYNqMHtFB4O+sT/1i3Hwvofmib34CSe8t14Cjw0vnjT4bjAG2SpgUJ
WcoCVFlYS+NxY02V2mQ6vtSjQHPhaHrcnmsEJCLF7WVTc/E4APpZ4fP1soxK4vCY
Tx6deHrNmu/8rMxvMkS0tIH/D9eA787SQu0sg1ydu6G/YQ01hLVXeMEbUgkyM7u9
HKiw0KRRFMXTiTA+HRMgLNo3gU1edXLIgtINtglTYuLgGKy1ELfeyFd5fgdhAc1U
TvucaB+NQqxXMUs67KbiP0E/I8zA2m0t9RDfY7NHEfyhgUCBacF4Tt01RRQsMOje
OyFTJWZS2qIIV7HEDYutOhH+SIGY7tu1R2UkcbaPdLmIdefXiCXMPrIwfsDnI3Ur
HhvDtV6DD01OabF+uy7BldnrwqrKP57zsQGg+Gajh6S8os9NJ02rxQFg5AysKgZe
wMevDQpqZGV2zKqDQVRLdQp5LIzbzhvsJaqxNc9H+ob8KOw8yjWb3l7E0vlcCOrY
K9PizH4NTCSe/+hv5R8b6suf2OaYLbU50rIRkeCRcbrBkmSDTTmj0LWhfmmZsZYF
k2fi6IASuhrkWkeNkQOrCeH1EDAF5H1X/RnfMS4bdo4aMNxkakruWW8b7eeSmj4D
BDyngDN2dtiqMx9FgvEEKZd2S/2gdiRAKrFLMl5dSl/Ci341J9XVU3U4DMMdGEMy
Bg2UdrN1yYAvdNHmQDGhDo8YSZmmT42/Uyj1zyAbeMiEqYYz4Ryw9emSUdL74ScU
xzdNyBUhHYsgjcewwmYrHxyj/QVvIQTBjBXEX9injwxFSKR9BBLhEr4QcQtH7InZ
kAh8DDFvXh19HZyWjPSXqrXJxl/F9uue5aTRWJ+yFEpAiZtiM3EAZgaCcgOAwke9
U+k2ljBTTXJvR+gtXFuT1fUhGXAlT+38ZNXXVRSQmKQNUX7oNl0MnqUEpN+piOEE
vlcftseWKMK4VRZAparqL/BmtbTonYBh0tNHVXr8A6o6jldQg9eONtRMbyBdxjhP
z5aYxrnFUgMuCMw2Vk2FdMRs1+8LPHN8g/ANrBsiVi4xpQ+JkvSrX9JHlNB4p3I+
bprf+SEcBGYAk70u/+z1+nOBgGQB0xZvETZSB4hTuCye3n1Yxpe30OQ8HPpB8z6/
GPdEy9OHB8KEWOHPbGA93B2STllF87Hy1RAyaePSfyPbvWrgDK3rNbtyGSlPFKtI
pshnkFimEm5sFo4aShHT5NLJKCAy4JuYtPSCCBULvXICRKgTNkrOOZz7HIovPB7p
KgE1xpfE27p/y9WulpebMTdlAUwrQo6H3rMRJkY3hQifZXxDdLyK6SnttCPwPEYV
/pRZnKpaZLZqIsA9NV6pkuJRiUBDyXYFf9e6ovgcFNuOPrTn+YVHv/Y3+KySHOEW
jTVMScStjBQbLGbwwi/raAbY0H1fMmaxdO2Gi9xRo//uAlSdqfnmU5KEKBiUj+KK
bxU22DDfGeBroAYhJKrERxuo6WYNaO1AuvuFlHXraEqczsNaRJNHu+GmMSU27Mkv
aGmuBGW57MeZTFiz70IlGe2rEMAEU/DFf1FjfbHOi/n66trjjhU4AA5fbqP6f9JQ
Eph0KtU69AvGmPs9p4/jXpO1IpWZqh1We5vUzdBbQkxED3BANokuHZ4a+gFOJtvV
5tBcqjPvNKiPcvIkHqZXvOSZS4PQ2OuhXKtsyBAcNxzT3LVsnrQo/oA/UoyjvFOB
LE8o1UJ5WwiwnNmh+/40TFb6lcFOTuevdmMZQ+ASNQnrrLcqk88uF54sf8h1c8TV
hikiq3d+sbHCCUDaYBeqipfwxPoyhmUUh29ahOJFqBPRcK8rZIqEAe8LoVjHIY7n
/Fw0C4TVm3a0Nc9yhItlZWOiIo5BRCCEQs/jL7Ds0zY4y3a8VXHgdWOY3uh57pJ+
1LYpQjLPgJupYas9H3/OtkGCfJ4q2eXVZQzk0GbK25vfy4ul4VhW2oW2coFcdjkz
0Pb9Vww3BEVQ7NZE7zqYNvGMZmkAohkOmNRJ40e+kNwKrd8yuAHgK2R4gYEnX3Be
zDQMhaz7rkOzWj8UuWZBB/lNbe1grnzRbgB/901TMPmfhsuPeP3G6141aoNYmcm3
wdeBoCgj1Gwbqkx8UPJwBqei2QkMTyFS6WmKX2Np7EpN3HzTmzbcRS7H6hCHR/OT
Rm5n4cHt49pV7Fjiaxa5qoJrWvhp5QxkyrTu8icrm9B++xkrjHmSGJfpRPAStPO1
FU6NbuKMMuO/C2naNJ5C7PiVKkv2EMncXPaIkx++9seYYzTMcxdyyUApoHaru1/U
rHqiBR1mdOVnID45H9/PpppXGsZ+r5+s8BRmj8MnORojkiw+Ic71GBkK7EZVf2KZ
gAHsvC9nysVNgAApq90hIjNYQHonDfmH04palDjcG2QrsQarNBo8q9DplD0w4sGh
Sds6VmUNOVkIpa6jBW2CzoUIAxRhytxKd3Nk9RyraOIZTD60q228k3kuYKYe1lex
qkTMjvBtIAEVZreLJMqCyEMezuztPVGm7Zp0SgRykE1gqLBk/mGyrtMyH33RlW6y
cb08LKAB8VKoRjkxlV5Uw3J/HQhB1x425depaqvuNw6eWcQFZfMWf/7Wa2pAVicp
6DuSyNgxI5bo5ObKKqXvJOsURUpjxECFaY7S8eYeT0kOEWfouRj/9ycpAVYIpH/z
Jlxp0ZP0bYyY3rNzt7Cnbx4vRBHMVYAeVuJGU6BwadGNAPMYwJZiC7Geg6DKW63q
FQzhchzqYo4NUPf3MPUHdynyEzazfTr3KGGKyyx2qG8R1joIyACvMFQtKZnAXgOe
sJy2phdSNsGNVwTuwff+4wqrG9w6X6y7q0IZnFXGR9XnBQ6zxcPdDJThf7Gn+wVH
bw3g3kvaEBEBQEoRokPaX48nYzJjrDjVoAd1oSWMYu5kAO6o+Yes6l1ba1V54t3p
ArBGBuskbaIPdcVIsTGIWPXqtN977IHe6I6XvIGlxYgPjDYfsJmgx1Ji+eYgHqZt
Eki2majMYCdjsjPc1fTya2HWzhTJ8OU3s+O/gdNEf+bVSx7NHiwkwca0Mrnlp39J
CoPUB+vEfItbifitodt3LNcdl+gVgw9JJALG9TIAOtsPmKz/yyLxDMkxaWBC5w7i
QgU4p/8HK2gd9oOfGxT8dXGIG/DZJUnIdil+rff75TVTzrRvnp6kgMiru2aomBLJ
bNI2hrUCze028oWEG0+bvobdr8glRC16YKBudpIlcmiTw6Z4wsLHeTo7EjeGw3gC
QarRoWYtxvTYi+PchYlNI/YYMb62dkTX6f28OtV5m1pHedPItt1fxLwow97JI0r6
jjHEUjXwOi4/ZZoP16Nlz2ccLj43ZsiQ870xyNe3G04A8KWPezBU3nZuqh4ngHZh
U+BY1zwH9r649yTSP2Q6oesXLPus25AP8GsijTBRPZugo2Czg0/k9ZU39J+FdrQ7
s9rYyTGiP6g1yKg/Ud+vMBfZY/Vt9oRQIp9A30S+8AgQNEqaf5L2J6gDLwVjEMUK
JmPkvWkw89E2DskGNMcDgRAqt5BS0vycmzT2WoN4CCcfPgihDh1JmXDd0zspkkSY
dTWzzQerHR0zJGqBvH8+72P0kZDAqtnPq0R/ZXbyesOdBICpLwty6OgG9B85X2oA
QlRqr3fOOY0zB04h+PjCz8s8FOe4UvSN3HbS/UlhXFGV+aW4KvdVwUXwNB7qer+c
ZOjLh1Drz5nn+soBeZdd3D/VMH0BA4J8wHwNWAj4pGfU4inHEBNlvBKZ/pjq4cwT
rvCF+VtnxkMYzoGfubRVMgNURwNeuQ+2GwqZE3rnWp7w+1mmFzLOkQT+thMsLXzW
HSPDbhJ1rF+92VmcU97mXKM8Rq1ST8ToXG715Dr/YpWzmH+buXCexJNa77HxsTRj
BhYZ3lKy8IVjFbFZFYV0PTHqfh1I0Jqw83ryOnlwYFOAfJtGGCQt+nr7hdahQrV4
sMG8TPe/Z/eVRiY4E82+y03hplIHgiD0EetnHpiemRaUebxVfZ8NrHOKL5elW468
a7LuBRx9dIz8tjlnGUzL+6MB/bhhvD91bW8h97AYOHFPO3yCHzrZGfdF4U1Pqr21
qKWVeVnQnbyBNXfFjOlbCYaoghoclr/MN8cQUY3Ei7PPbdexVKyVmOqAuEN2AUM0
2UVcwebT1jtuyRpkXG5OZBAqV836b5fkbiVwjsbBq1kL+XoTgWEQGqOwWU1Leb+h
PPoIgmt/Q+UHAjPrIJT6CjTDA3hd8M6prcecNAd4+E4QwZmqNaYvznBfL/EQTPuS
UcHtnjPkEGiB1c7dxz7FzSyOfMZTK9+vevNXiXsO7s5kgbGwquBr4eaUT7cQ4CW6
QVxxdA6S7IC27Qokbed8rmbyqRhIuaQgH6YZVVEa4EyVE9sF0Ws/fmb/mr1JX5yC
OAOGH6K/ZOZUY2iX3DhslZujTZp4VUQZz2/WRkIHo0qO8WSqFXGbiht4X+5O9Qu1
eut4d+LdRP5UFmXrc5jFe35oE6cwwD1d4RLY3E5Ko6OoEcp6tDJeaPtpeYb/RuZ9
i61xw9ndDVwWRvSWUb2Ja2xZWQhXy18fTOaLbaG/dqUb/bvqbztnAFer2NxLs/Vs
s0a8KQsNWg53h6AbMTU5KBk7XvrlnJcwmYvWEaNJiY88hBylNy/jsSDGzkhgcYHR
SdwkeORbHnQe2S53bBD7GQf58j6hp+Z5iGaJw69WlQrwX8NF39xmxLrT/7WKMGiw
Wb58phgS0IhCp23ais+So3lTljdvYMI+vrVifqjB4nYFfnB1M6mICaX5cXtfrJ45
VoYTsX4UAHHgP3m95T4NE+hRtteJByBrDxojqu7xV2fumEYz6dmOvEK94oAmrZw/
cq6PG1NqVDl0+0ZXaSDzpdxaYdoYxR01DfkYE03WlHzEohFOSlRztgTMKnGW0Ly2
wLnr2stFUvDuqJCFMA6AmQ==
`protect END_PROTECTED
