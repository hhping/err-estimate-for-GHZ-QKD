`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sen/GVdAfLbd4ZOGCRzgPn2DG4f/vCZSao8vh0aoKgc66ub8LS3/XQF5pvQNe8/r
Jnb94FMDw8eiO7Ad8hodWzXTNh6dKoOADkJA0eit6gQZQ5ROgYrnx/xLunMk58y+
W78kYB4zAEkpFGJuwaOV2JyyhEwgi43xzvWV+eQ4RIRHb5RwpXPLXhmXy1Y8c2B5
7b7DoO34S+re7gchsXCZ1aCngLJmLooRHAq4XdDwMSu/JUSgrOK8d7IJlNBKFibP
KYyFb9wJzBQPZV8NBAWcOWsDrReiffoZmQP9LbMzsc1w6Dcv0IYneVs8rRL9S/Mi
Qfp71kFJ5wt0/BdqbQlwi0JqOIUXyEi0SfLe0ungdmDdeXxQV/hpoRrLZ3oAMe6+
5MTJaLlsTl0CuAZBlovKe2kQp6WiQUIpkS0NvxMAHg8CellfOQQFQdtZGZeRmQlQ
dfgwq+Ml27Ag7v5em+G3zoiyuuxLzNiCCGHmsNKD4UBeyHTSKkIM7NwWpuzVFiZw
oDWjKG+bgmXHF5BjGQvUR3xoBNtpnZYAirwFzUZbmHSxkmBzdQP3JOTz1vfwGEwX
UTCAR+6Jv5GqD81y5Qx6mwujps/OnWO0GSogi/nyEXBfih9PCGukWvOWiqsjYzzW
R/CRcBp77szB7FbDbo3drng1RxopdRue8hEQnuGaGUE=
`protect END_PROTECTED
