`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukopUcynbB/6sxfVUkdxuC8ZKKh2fNvHicSMjgY0GgS/tPogYV4PS/gsevVL+LWS
u9MbTm2IKE9rlVglVDOAKZfAowujmlcca55qOP0YSpOVt6UVVgHDuYGPgp0SuyaY
azuzdumJcuzG0uwjJrcLNMPMRB+iN0E1e9H7ux7o5+FgkL2gAchhZld+Jmm3L2fg
dD23OJFhB3hqTsFeGps4NUfl9EJK6Q80sk6f2Ju73X5P16wtnvtT4PC8YEr+CocV
skq+TFueSbsJE5H81jxoQ0RlNXCFliIRk0vo3c+XRFnu4dWD21NElDjsZewMq6oj
8YCKJ/BrSxc/GO22L0M5/vq86f49tvgMaa5+ACbMLu6tPfJNa9FzK0Cuvwhprwi3
ZI3bqti+aJbxe6A4RHEs3iJaOhCoHEdocQvP9vY35MqPZ8tg8jdlRup9Hdh8NTqg
GZ0XnmAg4J2XXzrfPjqvI7Agobw9Ar8wpGuv6zPVrW2Yr+qq8Gy7E1cEgwTa8shk
g+EmuHZ5jY2QwYaIcDnYsXiYDT4EhtMbpqH67J17KhBiOTogKe8QtaZSgpm0MBGi
cD8KQVd5FIB8DGTQU+4wphimwiouFuAPpAjyV2C3W/5vAKcN1X4qw3MsSyn8jB8x
Lk0DRVaBEtEqfFFiJFbcSvx+RrVKYPjGYXXJ8RSlPadBHGUghke1eQ3KMtsU6/9g
4XsB8ais+mDfzuoKNZUBj6wrdXVkX4fqGfww1LJE9QLgPZB1xSDeliPSPRfgj5Vb
`protect END_PROTECTED
