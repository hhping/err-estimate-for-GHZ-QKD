`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L9HuJYW/86oHcjHTKXuGvg9ZC8SGk0VVLow9uDCHIYllo1AFwHNGTGrEykdiXfR6
+oMbNqVrk7bfpydonxDiJmbu7F0FqMu3VwqC073+iAxex6IjcrgOgUIQF2Y0EbTk
OKRKFkyE7hFsOvSpTZX/bGRnUi4uainOOwM54xPV/ULlRcQIr7oIotZp3ja7EOPC
Y1Wh49LpkW+bQ1GF9YR0KtDgPLWaEGLBpkW3DeYvxEHpI+xl94JXo1/wRnAnNVqV
3N0NfEUW814kV3zwzduHMq79PW5RNiT5RRL9YRNSgkEeRpMRgN+jI1z6kVoZ/seE
sfRhrgzwbH/thCMVu/6rkxvzUHIUA0Poe/F+x2wvvy8At0k4hKRtflgydCvl0coZ
Mhdi0RInqVk2aYK2W5myIkvIzVjg198o2olj9h3g8bsqdwJoZLBzb3iH00Qxl43L
yk5l0rYKH6mAlN8C+U8Z2RNrs3s426IqNbDt/vOBBzRGwzlaRzFwb+mh0BflTuMD
r3mn46HjP1+sEa2q819kSS6WgtEH3qYyS1QaNEv+PsSLKs5NdeqIJy9s/hPgFSh7
ibh/NbkqC8+0q2GhJyM4RjESQQmzcYY4GSBtO4KWwTKENc4QhkjxzVgHBKlX7oSV
wU7vc4R/i96zqiMNnW6CJ0bbvEivkIwq2/px425kxrIdZj5i+7sIXyq9NvSGapmX
cN95sO46/GWBmCoJ50dqiwwMorOjcvkUUri0rJ8HpZryBHypK28U4zNCv32kSWyz
mMokflpc+vTgXtc/W2smqbnMBD51DofjzX0+cQYz0VDcLD+EOC88KlzRBD10TS4Z
O2a2zx4n07yBw/BFVhZ86M2kXW64lJ4j//cwUY1nilTJbJJLyK3EdRS/xvDRQ+Hy
D5NacEyPUh797mcW9rNHWrds4WxfCvknF2pwBSuM4a0ZywEOfwYg/wsvUmey0fZA
QQL0x9C1R3tD2GoqERrnEfg6sd38eHN+KgiDrWRHqQ1NirrurH3eVYHf4fhfdHE5
ztkF9D9glPbj/tuCOXHBWomRbbzmdkt3I2/02RdkXJkDB9LovZHOmzfxqrP70ddD
Uuyj58qOiZjvDDX1Ax6SKCmPZ4ApdMewbmsUyjqjXf+C7jx7z2X9RRD25oWyO2G+
gEdVrtd2Vc3c7PrHrE+m/BSHm25U/W/Pb4Z3EinkkcsInRMUGV8HKlucx4nqpCXZ
gggjmyOKqQgmLO5hGY6L0j3sKueS351nHQycW9bmaAoGOAtQgBSQLFNNPLuXTF1D
0r/tPIiW0Cur+3q0NkBk90sjZspAZnC6zHOk8DxRCW908WEKJn4/rLnxjcZJph40
drczZXMTINQcs1lH8H61cJOHr2Eavy1WLUZGM+Sf3LWJ9MdkiKdl/kHNl1SYStZg
BTOl+97GOp5R2lGcwVxnEjXU/aiDJJdMssdGXKr1c8C/mEj/oLL6JSbBBFYmyIdA
uADIGXB75gAcZH0mkUMogPWmYPFeHfQqtZmCa7spOHshoZ7v5pnjVludlJFTb3qc
Lko9HYtJCSt56i63vEvx+tZw1Vz6WXUW3rmuG0hEkoLfzLJlq5NHJ5y56Egpd2Oh
j2zHc3et92WPmwbVPchx3eCTdGq9MKdlJN0hgdqH310XPppE1bRFEoplcJ1Wz3zV
fN9mroqukeWV7qRWIsK/4/R5J4SRVLa3kzHW/DxROYone51RP0Y4GEAGMS+MU7kT
E3cSKg6mJDJV9EPxNOY3Dynp1wX0l092fMptA+ICLbzu2UBuMxTGEc8yaeg5NRxs
hCNLZttu0bHUBc+6aTrIvsY+ci2RJ3Dr5dI4I3MhZhPFrPkgf7s/0/X73k/W6Vst
+XGfkFIN3KMu1L459Z8yVVVIaHbBbkxUpYexQHsKaxyPwibAji3MFfOo/nDNKzdw
VL8jDzNhbyM7vaHu2dNADCQ9UGw3LSEbRQcALk7PVU5ykmLH64r0+NR2JjLHeLe9
mttERWke0Hq6HAGahN8wY5y67t78YOaWnkm3cIS3vmgJa9qHBZ9SyzgHNTcIDvvw
HEA71Vq9cUK0EalogIBNconROIZrqL2Hf8D2xEGgSuKyOCTIrtFzuHSzOHWqWpUN
WuWFPCPCC0vBElHQf3duNK87ZTfa1qMbrXeYzTiUxZhyCQtZxMZdpzFjL1CPhY45
Bi97ukJPJ2ZFVngx5ilgHFZUwWi15oj1c28htf6oRtpF0qNo/+LRz2G/8+nWuXRJ
BCl+Frh1nZdVXKSj9qfKOZBxuhMPS9uvPmei6hHtufV2x/3yawDIDl86vI7Q9BZb
faz7A0d40J1jJGxwx7e4JRNrgkMDDilFVa+lBjep4TCKNXysNu9Ig+meUFbQVskN
l5M26QPQudAeSWxpjFAio3r5deZNuvoDqP8PurkT+ZtQjvwbH0GwUBc2ayvAOLLA
ebq4zQUU+EkwdPaF08ba+K/tLH4TE/Qra1kok/QswMWbh+SogkmHbiSdENQrfNFv
n4CF/if/dOHjDc1LMtmY7abLo7n7MsqhWkZYXwcrJNhfPh2kAFPpegJ8RbtMCXhj
MIlSxw9L8adiXo7tpsr+sA7KeSTRlGOsqiSb+qo+TrB2iv75LerCIoF1/k6YhMRK
48LMPdFgkP44zt1FqfZwGYqeFJmSTvbdv8ZkxgtfJK6qdrao56EDQoxxQHHd4bzt
2MqEj/8FBTxFqgCZQRsbZJTu14CEsnyrzMvFBd+u6xjP4sQZTbwAYRMbEUyUOOrK
1lDTBXJ8LzOOZHHajB/oaGOFbfiYr45qwWo+9raxTu83Br7VZcjMK2FSKOENi9WQ
RPUHZlEfOD/m36+ybfvnGxZfoe+flsngt78yE6jZd4n3hI/100iZ6eu5A4mPdmSS
oPC15Yv86vMSZZhNsDFFX4ucAvcDNlLd7EkeDhQc/4HITvKjblJWAgEzViEMD0ir
0V2zi7I6i/nlNMeBdblsSRy1kJsEoL/m9IHjZLMYnPRVHrUj2H/+xkZ3rq0WlFOz
xBnYE+pJg/OPvAp2Gzzl+W9qNwb8utBehwU2Jt/OQUFXbZeO7Jgn9qUSNwUDhFCL
KYcX4PAOE+RMSsR8dQ5COiCQhU377C52de60DJtSBGBm3N7rjjUBKrNxUDfSAC9R
KoldePHx9z95SEJVxNJ8HjqlXJGTpiQbysjQk8PiYI513hntcw19+UeLUPppMNRc
TkdPhOIpLRMKBNBZR0yfD9vRO7S3UdVvdlvuPWFMxDcmTyx7LpcTmfo2skFisKQT
RDZtLBlAi4lPCBWRDweyKEJNjPrl62ySau6GNgchIpBOFfGwgN1WnAphcceH+7DR
1gaoraUDK6gJt5LVS1R2iLYOzNxFlDUBrq1JSO0tcxCMOfi1KtQ7uyRdeJn0Yt1o
5oE5oSh6VB2SWjloyHMacC5eakzN6OVdSc+X6yJ1oEdx+2FPHLj9DDZ6xxeGsNeO
S0iBJg3L/o9X+mBikg9lmwqkM8Aqu0YGCbfFVKA/t7KtldPfIbKYKkUI0rKwJb0Q
lDH74cvnWpwzN5sEew4KDpfGTHev4JLmHGJYQGol5ofNbHXssnE4P/V5jnwO/emF
ust2wgaoDPpw+F1hKxOPJZ68yVdOZKSJTHuorEUulsJoLW+P2Z0x8JTtxkPPGXyr
gsY6kbfdN+2dcAvS9c/7QaTxyjX4EjSOl1gHtf4CA5/7KpjIdjCjqJpZMkxN+ZVJ
ElvQOheZnq6Wu/43XcxoOsBcDoDcGgMSOpi1e9HyVKxEYqYKRzX6HosLrAhx9nrK
PIcEkz8/xa2hYTzLOoCdKYQZ93f1IuT/fAVFGiChh6kklAk/mE38G3n91aasmO7I
sUEYY1dr9u3PT4UKMTP3owJtMCapQAiDkO/L2ZwX5oxBF51r23POgzzpbBEUSuJY
4G66cgEEQ6Dde4s9/dYgGLAH4y0b22ii7vl1VzLnv1oZt+5n3RNaAQEupvVD3H0R
/CPE1SBuE9sWfaobQ+MmaR37aKrN6bC2Hw4K+R1PuX0R2fzrzuOUHFK9KVdI9nN+
PRdA9Q5ZGlHHP7SQm2gTgPm3eXVsrij6m/qQ75Is4f0zXt/Smxknh3SP8JtV792a
8EGlDxu+UELEPhFWfrnTcC8rsVN5P09nBzfsrEiBlTA91fHMm4BhxuIH95WdpYSE
uUY34XDEGE2UOvpIucXKD41i7XyOK32jSFf9tD+h94uajGNsGM83R7AhRiCbzaBi
WsvPIEnUvQRACTHBlv0IDSG9hdpc3JyOHx+D/rgl0FinQlWtABan4NmizgEIEpQ9
ggTCrWuq8CaFWLvLxVQZxQFAMiKMVTa6fgYsBbKePuhis/mI6OySQcNowjXVCZ8y
xzvsF1U91I6Dqa0lW4iUkLI64PuwHgbzHOaefVqp0DC3qIbxbuwFoaGYctMpEls1
zFaAbGmFaSAhtcOAy1YdMXlmKwD7qcql73fAQJbezyTsZ8OBpz4KKQF55Iakx+WW
FhA2ombMrRCJOfFtmd7vFgiODr4nTuTbFxQHjxalvSjMoj7AIAmdzeHTZEXGg1Tb
FC6y+Mz+DTWuJ1LvaARIPah6/6GMGllbvJpLKWqOyLxYkeFnokQl/4cXscc/dYZt
a0IDwWzKYxuU5Ma5Uc+7uE2AhgsQOYBSHQmBgv/F0rhWz8XbvpyoFO6fZialgC6/
R+OntFDp1yPndC+RhlE3842+kdKBBf8Z6c+AMnbhoyvWK1tQn/5Nx5HHvPyCKTnc
h+g6kpiFhjGTmAQvOCnOrfFtPTUmto1j4PcFlaWk0xgjIMvLcBKpOxr3045Bn1uB
qMBOd2Ct9waEy7e1Bi2Zr9JK9/kkFHyvIMSztc5w5Go2Nk7MX6VGSRUbXPJkipvG
55CIFG0Cyrfz4+BuhT+Z70ah8PHw9cdu+0Ga77pzrTeMjahPCzwnQnFH7hobRZ54
n8hB6irNBa6CT+mYcDs3YB7Z8oEdWTUby4Hfh2kaHYx9BH2mfk4tVyvRYzMKuTLY
HKbuWpIq4ndx1mz9jc7MInnORwy7E5Mk+a38x1B7hKLVsbDA75zQUFQRRJnXLpGM
KFtArdGNVE6k/DOVFadq3I4yBeTdKWmLnyZBsKCJ95cDh+d5lg6S85svVNtEqoj7
YeshGTiFZMH7M7LwpnJJgcmu9wE1sjMpqiyQnIkosp6PIVQG+IjPB8yOMD5/S79v
sOp/RdkxfPCqBnB/YNM2N58ycdOxGzES5SqjPbvyWd4iOc6sJp58H2QEA9jUiyNt
znqtVYQQ+khON2/MvaRIRMuj/wRaAuFcXbhXjKgN0D3vR8TjpZS8Xohc2Mqe2tct
tdyi1sBq5FbGA+lhSlGp4gGqchdWpYfldq4XWOaVT51QgyjbBD08ZP/WxOxMmFjp
RyeVL7hrRYFsewsyr5RWIze7GwSwQ+qT36AtZxHkZ8TvJm4ee+rcYnNWfmfIkolF
L93SIDyATwEDiPYJpSlvCzJhquh7j7Hqp6KFDXtId2JsfKWkyoxxnAUGU4Yv9Hfc
VqlPpOh5KTEW0zWpDGqMGWz3wvzjsFY9BPV+I6s33cw6RKn5cyj8WAz6xfDNKf4N
Q9uGkgAvGHZ5GbXsrtzcSscc7DctWrnqJOloh6SB9mTGCAOlNTc9WdZmLv6eYa+d
8uTIhTSSLHGsEKj9cmQFBdfvXV9kldsoyhT+TTcqXEnARkcj8QSM6ffAstTjfosQ
7q1+dU6P2X81aNJvjmJU0iRJt/L1KuxIQpIF2yNtQqEM4VloDYiOLlbxFyS06edN
rW1BKEN8YDt1lsEWoApgdEhZGmIvOVD+fy2NWVadL3GPxobgEOAww4ikZriXuyA8
GONZ8P8E8P4QbqcXBcDLziizs3SWrCeDSeV2PFkxTlPj7MVERM6+cajYsoETH+lr
Wk6VnDMt5JouRhNkAZs/uWoJuMs0/gQa23GBDCPnXkVp1T6fJwp//3pDAptJuj5c
vJ2LvvNAiQqoSOlhRTm+d/hjaKFLlBLGep3jFXnHQRBsIp9YAA6tGMGbW00ty5Im
lGeg5va7UUjG+XQ2kiYfiVExbawh9oh5kIy5gcd8AsPS5uCAaQFJdP7oXLPyeBhB
zbbbDCxS3sAXREuaxalMnea2cNBzRvU/Qi5MgybYIZuZidGzDXgtr6lSLmScz7/O
SiCsmHw+yI1gl+kNCxih4O1/kdUBeO9H0MGtLMFhcaWQJeVLtWtDLVQoTF82JS6y
17JpWGnJvA/lME4FsVVEx+AV6dpXzqMLLJlQGYRIimFMGSBTK6XVtZfH960EkZf6
4tn9mMwIWLYgqRoCUkvBB2go6LAv1y4G1sD484WX3G599GrtkZTh2tdyP6SzB4HT
AGihhJmWDpvFDwC0RpRdiIHEJ8AcfErvt9NM8jYpHhM2DPxLTY2iMnz5YDyDV7kq
/0Nj6P1ndQ1gaV2aeLxceBqAnHKshCagzb6mUqk4BVAzV0TnCO2sNOsjlAoVUgb6
OPsD9lfeVLPSbHBqgED5AhKwHLwvfpzxJ2C04kTEG4EYsOgIqjM7HCCREx38xZRc
AHb3KsBTcSqFPz1U08D40Sc1xeNUltdPKF8A8zPn4j+Lu/oCHPMyclwdNXvsJPzy
b1BCIFt1HdUtP7w60Zpe32ALTBIw8u99RzO6Fm1kWqPoVqd5vf6oZS9boU936TEA
Ac3rnTskgXumxIMRAEFhS0zH0K2sEvuWlCQZGRtzUIuuLLFhbyo7wMLvCexiwwUt
JcBprs8DrHHYajAQy4KyPUtshMKc861NWDr78/QfqqHNLIamwrdZPnMJgMFpyW5c
YmuPSAgniZCHZjASRjid4NBdNuyls7CYanSOpzRma89kP74wba1ahkEjWd04htzq
clMs5feeWfJBgb4R8PKpMI3AJGraTpTC95U2Cb7NsrlFCYK5Hcw8Q6Tsh8TZZKGd
JaJdXqZ/6VidODRtzNWqueZHkNUki2rCjOaeLUnMwtBpYh4K8tg9yagsnH6G8fhY
KQslNVBsRR6wIntBAaaL6hpRNXDZ9avTTDzgC/HgtURxe/KWe6z91dNlMdPXToLU
+UYwzP6lwBS7Ilxp8O10eRIWYTMy9N2nyp/rW7dl5w0wei9eyWvI6lnJo+qIOf+J
PqfAiVvrLNkMGcThDcJ4M6FtLqph4p/LfDKF9/p7suCwla1vCeROHo2FO8J2QMn0
hskjOV5qVB9cbvUYjJah0SFxTUJKO6uKIThnuor6lrxKvRMelI1BamJ2Mc59bfAU
yMG4r4GjInQbg40KpxkC7DZgKaSqrv11NSjiNCfOsYk21kzI0qp6x26j1XUrolY/
sX0jsi5s9FT5aOagimRr2e/b15x/3W/Z+8/DcbuGcmSIJCpeGjpFPOJkzZBHl5mO
1g6hi2jUhwaT32lMq+D/dlTDDZ15mVfTiJr/Z1sLxLuMIP4ZaV4ylRmlKghni0Y2
tXTXJvFGdP+NT60ZP1yudjQX51KY4mZ8hdWahGJt2XTD3rHkz+BhZloTCK4m5Uih
5obmzvVtEPWc8ALITTmUtlXD0kDhVCIKvwnpAm8yCMB/xDaPDBeWYpjrUh0vVSlL
ATVehvVpT/vOXuKBXCDCXIjpo0hZj1ypbcvONL6ChNit3AeFgFoF/cj5PAmxG/hL
LoeUoiZS1iaGxq/fG3GmhPQPK7uNgZRo9dMmYsjCaKQGyuOlNOgS7csbnxB8W1ST
B56VU32UcIgu2y9iKtEvdV2uyYmYPhWfbmk7pRmNFq/I0wvo0yhxDNulK1HTNFpD
idshVnn9aqRPPNAgZMGJ1oulB+Jjd2hd+10XgEsDjskeg7UHwKT7k/c/Msi7HQt6
ggtZXf3/j6vnMeZ65HVeEYUmKOWRChdRFQQWFb1ga8Ay6Pc1ccoNVf+q6+CABDY0
iAxCRxZ4CR8dw4qtAuc1EBaeN7e2MKc/5IIo7JWV1HHr1ivUqcgD+jtP26MNuzjR
JWIluvIUGx5uGBOpnBtjRLRPhbUbQ9vv4n/PlkG0cZnsRiDiHFXk6PfkfXt0110V
SqMCiFyVOYeBIQh8znUGXmSzLkOLX327J8xNRUOuumUY74f7hn6Jeerz0cms2FJI
uNDrcdCXFsGg7orup+tT5oKtrrwdfFZnAE8abTryEEryVGBiBTmtXN2nvyRAMvWe
Q9R5RhjA29WFFeeT6JA6B2LW/qY8aEQk0L0w8O0HeJZVnPeQuDtkIXwhO/aOtgvD
flAnqeqhk3Vv0y4lhhnUMOsJHx+6qivuZZ3wegYKxAm5nVxbjdChVpbgtEZtxHc1
syDzCifuyFMQKuKpayBZ630xRueDDrD/6w9X9UhyFObeRicbU0k5P5XExZI5wdNZ
X/ijp6mTXW6yEUqzUYwQmTZBubvCFHhoxuw69Y5vD7S2jUoyKFlw3P4f59x6A5MG
gV3g3HWK27M8uwp4SUMm/oXjmqafXbQJIBA/ykI1gH7n4/tV8N5bBqXyPRQMgXcl
Hqbq6dtbO6LZN1BJXS3U8FS9QB2XbKwakICg0j13M/fRuX4gZFdZrITZVTdqnUT4
PZ7VGHdcNV4TadQUj8X9RFn6gYrKSC4u8j8OlstA3mtsn3uQ5qyGXtjrrGOjhRsx
1jIcrB6JoaalESDRPaB6sghEiHkvu9aIWcAVaHUnh2fYoEImBsnMEyoB6J9t04Zu
t//jEjk2wIfn9nFvwocg2obaVG1L/S1YbOWS+UI3Aqbae1we6zAUK9WbjdbFA5mB
7L+jC5X51uEE2yNObLgSYrzrb9Tt9S4Ult59jb11Wj68cvPRpPYwDhN5LTYB9LZt
oevDVUaXadqKTgM01/PButAIDSOi8X0F59dLQvPo6sORWiPwY54qDctYlgZwQiBl
neO7NsPPNCsxqfq3/F4stUjZmVO56uvL6+haprc2S3WmtQLi06eu7ncW8jO+Hroe
PkLSuvg9hBQ3kAq9eSZGJKzMt23XvD6PiBh+8QbazF2PtSOzUkt9Tom3+yf8N0i6
EPXwJTuD4YE+B2cNKoZyRkXDBZAKGr8yoWPmCykbcIak5e6/zbTW0KM1w2VoyDuf
GOInZBjInB1Z9BB8PQHW+626jHCMxh9ygnY9e+ZLhOFaZJJ5jqOXVhpfDbWOZ80u
69iOPlf5G7U2YZkpNrhqFJL9w0Pt9EXFCgd3SQOlg/kWcRrUwa5AKbkznSCBygG3
D2OEBAJqMDcikKjhRYDgZ5B0VwIh84qtydOCl8v2KgExLY/NDVgLVo/RFtIXq3DM
dVBjIDUjqqBlcl3LIltdalIaDc31Yrfi2Re5oSJ8VljQfGe5fS/FiQSiXGxzegVJ
M70khr5D/Y5uP0Xe/C1RrVSXHIBhfxwMjng3ZKwvw7CNtXqQyL4JUyG5Mpls8RG0
GwForjGvuAGnt9I5+iCSYxzCiZDBs5j49z0yr1qj51/ZnwfNaAFfCI+bAKUw7ltK
deyTBZZxIKMv4/CTQ9JNW30dB/1MihNEqEDb+AUXDv5XxAVRbOMEqN5PiF7RREZy
6oPy0eYO+SfDpo/5OKO7m7Hrsw6kwe3/ThXlQ6TWYeGdayb1gWBd+SbvBM0hMx6F
V4Up9nZO059tgfkycyfQ6E31/h9YLxF+Fn6uRrdMU2/o3zaJHHdSc1kXPq/mIBwy
YH0pgn7ZFwTVSF/AxdZAiwHe/wXULZReIL/OF8S1Qht5e+zwGitK43bRV5ickFrv
YLehok0Ie1CKaQTFt8+Crc6FJGQK2C0hSyD8fKwC0XNsJiYSBrPjCj7g76XIuf7p
SpLDtFm9GOkCpbk4cUYbLO+iu4SvNTPk5B0u1WV8F6RalJvvaKtatIxNy6OX1k8+
EYV+IPRhfWLKMDO8IktcFCldSgbmKhwUM0xhzJNndc7Aj6oP3ndpMKu1WCJMAqys
vhTSxOwzbtIeEAi01sFXTrtrvRn5/EJKPm3QHOKQXCtcKcCi4H7mTJ7NyslX2+un
3pwDehE+R4SmytESKbDJKlhfyYjgqWp+fDhMsMWf8E/iX1xdEftr1HcjgxaqFUUp
pWNwsx0lPA+/ckGSXv0Ups5Jo2Y6ukhmFab4gz5uuWMG1dAJum78URgn5RaOuK3p
VxdzAFCoxlHErTBZcmygnd1+ExIo5239DTG+gI/XjPfXkdQ05g+oViXq4SAuL3gd
BGWlTRCLhfDOwOdGnVkEEAeUWV9eWZD/NXtXhg2+yNMfw1dLi/yjMDCVzBe7KWpS
ZIgEaSY4VEZiHKp5zo4qh3xTfIQEVzwiPhPluX48W7Qy/kopnhsSnCwoe29wyeUR
KTv/by3C2C075OhxWrl+bowiJcQEk2EN+LanGfz8iLHCWpvdN9WhRc2hZZjNsjp8
Ru7rdpsDoAFW7s2Vd10CpR1g1ATje10y2f7UJGZRAiwpkhMMT+SE4LQng0uOV/Sa
adKd8+mPXYqWkmxpXL67TfZpFgHUn/DHv+CvTVFbDB9gWs5dU2oTU6dht3I28qnk
bKIVIuGHJ3tLSL0MfonixA51bLgu5Q9wbdVz0zSGIoSsEUDt9EolLH36W8i0IMPu
JgkUZ+W4AowNZge/gSqvJB7QGetE320RrDk6b4iVGilIWu7MEOja9mt9ChwriSRp
xM4u0zMNCaTEGgvMfbjRJ96Cplmrv2gM+2I/H0rHjZxvktFPnoNjFlRa0OqJpwqq
GNw9sRQB+H4GWa307Qyhzoci/Bz3AQj5NE/JBl/kEg0SykbCPfJUHHhQz/Y1w1f1
EGh5Ko3KvGMEKSlRuqQLIxbTxcivGOsRpA8ZPj2WlEqflddoiBGHCqd2MM1OghSt
VxHwEXAkz65FHnePyoJFGictc7SarovAZ2D72YeAXE0GWhgMHID5OhBGEVNzfTmw
LXXs5hewnH+ySU2Oxge+we1wA8n0KPEAPK3DncygzZeXXmRiGvI6eMZ+hV2X598y
pqNhELd/3aNNV/50+KAHmpUT/S1mE8ViOhnthjCbLsM8dlA45HiBNVcSVJX2LZUy
r7j5T94MzioLYNF91q08bHGSPpLg9Jauq63vvdIOxT7EEY1WELablPwDEhuLurmt
mRssEs0d+k+nXPd+TtxyD/BoVkzCfgTZsshFrWFL7/MzIqvISg6MM5zQbXX6sJNA
wnvjU0/g9c4HkjxXub3Is6z0mG+PsHzhxzqblNxeKra9sYvU/L2YqsJ5ZeydUD4q
O8bA6xOgG+91f2CYKvL/tni9gHZ0lh19l+EszDnyFe11DBwh6vz0Ul38ETstQuzH
8MkTIfTHo/uFFlaEpCIxpeiHrXRd/1MFgFQkmXjo3ZnStgfmnvxIjDL8/22lSUQY
NR3t0ei+3aCTlRUQN4ldObKmpJpHh/akjIVCqiPouNCU6/nZQmRPcu7AuSe+M3zv
ih+vhsn8GXhHsXLuq9AVVkNQt1iJuCmTnEUP9XrNrLvKj+1/LaZ4nmFF1VWxEq71
Wwzwtxf+N188lTSvbjFjoqEZX7CQ1Omzf6aJuZpWiWQ9EH0jXPpwH5Op0KME3xwC
vHIn4H+LYAttuh2Cc79bDiLNERXGOXFbFe2B5JkfFJNBJ8W6rzKoz9SHTkrdnjnR
j+HIrHm/SUUgtvkGB6ylo0C9/L20ZbQkN7SCxh8dWLE4NRs1I183A3sVSzbgmsM5
LCVlwI236MPX/Fp1RBhGNaR/nThhDv6395C5lcnLT4Iiuz9Nz8FYxgMKMij2CizP
rboiVJwzVpvwXzfCh+b0FiIRL+AReD5uCO2ropmJj4Izbdey6icdz+LVG9YgW6Bl
5ses0chMCmfA9rXrvxuRjjP6pUl79Q1MnFnkmw73dOwhAgPMHeQ+VZnPNeA4uZSD
RhNOlnoZp4jA70K3DhoSSR2RcMV38O2g065DWZvYhvpphPkpVaE01+YZOU8vRy/7
KoOoyvddhYtkuf6f5z43q7b/PxpQrgVhaGa/4OHnEPernY67KLZrZDyhu7/Jq+JE
v+yNzhPCZfeNrz0fFHKxQHbPOLXLWSbz+RiiJJfH1W9iaRPMD+ZsR6q08qGdjOER
fXvnfuNhaNkTMHqlwPknSq8isjhHDvhbXXHcMpEQRpRBPFJ2oK9eKjn2tur/OBwP
Y3fG2f0yJyQrqHygxMmyGbPzMku+r6f6h2vDY+I1HXdK6Xlsfs/yncY8W77lDBJV
zbMdl0z5QCSFSS2qD6tmxpVbCfmsrUUDsASyX7aszBBUnam9IDVC9qW1q6dfusZs
jcI+wqnwi28oCzlr0QtmaiKjCeykYXxiHvDZh4Gfb85GNtxTc6IemOxsLMu628Oc
Bwu6rCqEf3YkJt7bPA5NQBtwVqqlpfAO6cOco0rh6sdP5FOakdnRZk5Sd4hTs5+n
vHhhMigVa/sydL5X/QyomCIcsnb8y06/GDkT3JRUm6h9hny1UrgbwgQRzoyvMRYW
Wpw+NM9lNRfXNsEAG/NOEj6LyBJExjDZXfL+kuKIy+vuQQN4HL3cXF9bfXVqcMeD
na8IOxvzsF4GLeYyADWH+VXE8Qjb8JzgTJwkDYn7LrBilK6Yp7KvXAQEzXSrvuSg
Si69q8l6mzM2PPtePgNa3xw7Jq1Fd3rI8uwACAXin1tVPgmiybJpYrpoIxurxQVo
2/zAiAEYnVngDqJDhRZW7LVr6lNihCPeZ/HjzF5CybYfr37kj3Y+09IrzRdc7/sw
f3uucKrH+IX2lrEycl1IPfO7xqIxXbuAOVW+PyvcDkTqXalGPbx+KSkqcBBlG9Q5
rMreTzRFS4+MR4rm1m6gm6xBfxqrJ/MQnqMyTq83cFYAoLRUGEe+LJOehd75kNIG
ME73YyXyeI1bGsIXqBXMWci2y4KWCsED5tmR4PSdtw9xBhwwbEOdmZI6FvHXwqHj
bLAHsqtxHbQn1Ea4XUMF621W8f5+HHdn1WRbv+Qpmfq5LLZuMnr8P8NTTBb23/N+
VfiOYZUzxtfUdB6J7uaX7grQ49K/Dc7wU58kdhNCPxiQoK2+3LnKr40sZ5Ww4XLf
7ABAQ+hhljvfuiWEeHb/UXVPe0Pgb9630/EgHM0XS3YNZbcEZuX7CjnLu8v14GSr
CUJ1EPg8wsNChzj3IQW2rLBjlMPh4pC23ea58CCjgtkTWf3EzCBCsX+KB+AjZrCt
RI/Lgth1oG6z+oGpJ0Dqs513c93fCMytCsFLptg9yKk9ltXsymhjeeePdDxfPa/b
Q1GvAXj6RHqkB1idD5rDudEXaaPZ0V+bUpex6MiK7eXtzdUq1NXnsBARZLvNwAa8
9GCoNKs2bOQ90okU7TJdXzfzae5Y/u07nGpH8K8Epfr3sXAIIKuOJgjnJNn7ESoO
TFfnAdTDOW7LajjstAwEwfrNebbcBHfqOR5yuD/h0D0sLFRWwIjjw+Ux9EUPsMFZ
yfjrXeHRObFucSnL+CdHWhYi85S6VCPPqt6eM0bjQ0xPKB05yOt/M59VnXVxJL7e
dZpN+SDnrIEPEiatKGiREALXGxEP7OrHUSPBINopYuWDt0fzAg4O6b0bs0dtwEGQ
ML1rH+9wH2roafjkPjz66pnsYly9MZ2RLpx7NiNtNGs70u7ea9Mn4stx6LvjoroT
65U6Ekz/NKquf0bIaQFZsxbO/4hpZDyPeQZSC60NHRpEaetyJCWz8J2JLU4kBmlQ
i6bGdNIejTdv9TwTPY6bCWFHh1T1PSXfIChLsQLwK2swGXHKIcREh4UKsDPoPhzh
R6y+NVqSVdVvzKkl5QhSksIKNctZE84YF2+sFSP0Rw/tryHmlomzOjqXaDft9Cs/
bi9Qsg1a6peTjI6NqjNT4475G8sR9dep31qz8QNi1FHh+VuRtU3AtoIYxtN/3+Ne
P3YJ6cxk+VfwMdaRPAl5mw1Lo4yseSKKJVsaa+ACM+3Xv78GwIk4e0TaDHehqNKE
Mfddyr5IAmP5wDjL/9jgqqxiudhhLA1J5wJUX4B07gSh27DBnAqt8Pzbz41Zr3ut
FQ9c4ke50g4bcT6D9wnSPbY4CofsYlVipfpp5u6Md8cYlULmLdPbqY4W9DLzuTa3
sIEZCbdEcJnbgFxs+n07jt17Xw9WfZfb+CY0cHmW/N9pkvpFG7Ah6SDY88pV/3PW
FmuRh4a+gZQtzkk6FRV1y7urj9OswDY5qa+d94QLsYgeTNAstlf62FiHE5DbJsvn
VMLwZEOnQ/vKXGwhnl6d4I6kSsgiJ4yGgG4xyPFUU27WJrLo+inodIkOJUCd9c4i
Qy7xbSr7qlY0EtfnAlCOFx69vbAroH8jDji40G7IGn7+vwLxEYmACF9CWWC+T3m/
Nts3w9zmqn/rHKCOvlb7x9b8luEo/YY8Rc8VFQ/lfI7wCPD8PlReJY5bwD26Vmr7
wN0EIUCFAC+Qc0U4zW9u5thhgUwNjYyQELVDpuNyd9OYZ2fSn8QlY1rDhrGhlNI7
NSABk2Hhh4xokHzaPv3jsvZqU4JmeBSfVHOgTZynK25uDIxWBldrnEQlmKyzIN+i
N12nZJjKrNU/MrbA8cvxhN8Te13UAYL4M4cddk85AILv1zfavr6x05HbXOhgdgpp
t3oXBLYXfwcqquOaABbIvfxG4fGRlZWEqORET8xc3VPwgSyQncT+k+h785DNZsX6
MEbhVLxrxQ+RGeK71wRwNMc9QADTgmY0mG8bVQG+WMRFoUrWkE7IcXWXVxdX6WdY
PUbnunGhU9UKUTZSNTpWc2aONWZptIinjkA40Enlu5FubQN6Y4sCCGVyTodmzByj
2N/wNxL4pejj1OHwrmJ9htEqr2gqO0siV0UTxPfgqUo6Bmysm0JsMkRe6kH1OIFV
7LmjkDTQADxrZO1FWD2FyMs+Pz2Hr58L7TbfbWij2bDCkYLdT7UbHQmn6Dg+fZgx
Pjh1mEb5NhdRoacN2HaWbk5HZULnexDp9+kQelkFj7/rpq5qqGcFgl5Hddf3cgz3
h1HGrK+xEEDyS3nOYs+aOgYpSKmFqVKo9NaUpJJKIh36vk+y+cz93zTg5aUJOnin
iq1riCGPSVANCH7XpaG69qu1VZaFDnKfv6AW2cof5sl9n598N9vSeakWhTTeej5g
2VCZeECBRrcEel7Ihoe9qd7XMBK+iox18P4kmwRZi+XAUVI3iQU/YbtMUYLmD3si
VbOyFzxN9Bg/X3w3Bq8FkzokmQMK+l5pzodfuBk/UwJEuYgzMNUIjAPsoja4GFE0
jLjr+99Av0/kGGzXuLkU9P6hTnHlebu4A9a/9TAsUz43iVuLPpxDBcgZMxIX7wre
zI+vMbu2SXO7jup8r235tXmJvSGz7ujpz7yndAwuwDcrAOur+K+R+PZpXLAVrHJN
lUBcUAdIDUbulRD0luWAQCJw0mczO7nOChbKCsCwQsSpRf5EXjroEMdOgSZLWaO6
o0JA+40numBqUV8+PbetA9GV7wdkMgesGI/iq9NyqJXeSbTpbjSlpoqBdIUENfyT
zFoXGB8/jtL2HuE9BGvHXPL6JQ7pFZbOkPGSTn66narGUxPaXZH28PVCGoaOC67t
o6G7A/yeW6Fb14g/DWErGU1CbaaJKw5yUHTI6nziOH+Fb42W5qxmtIz0dmDaqqkc
DMC8+zc3NMtyYQ98xaL9kJxGxazTDxUjQItzOd5AsvazPvsh0XDDuZsoi65P/l11
YnumYObmaAZPcZe0t22ZU7G/3gEWL9cqNiKfZdhhOJrmL8lPKSHVr9yG2RDjqlug
l1/FP5Zoi+aVrxdUhBPqC7CzLdxK9gVxAPwQAEc7ZgNQILuP2Hf/wojZRWwkH/nf
QXqx/PynwNoYvyiRk/zXeVVTngXHcNYJ8btJAf1W6GYi6ClC+lZzjJTN8LfHHjMQ
FlpDmBETs70k2yVgJ37ctj3PI4cPJ5gpvh8mQepWDJATwMZaBGpRzHGZKJALsW5q
iHcIRKkA0laJXVvVaOiCxIASE0QKJJSPl0CWYLnxoHdNJ8jgb9nHId/TYtJjsPXP
JQ80kJUKTFjs+AM/vUpW4JGHul8p9EFPVqIutzT5qViIyzHCMwnZ+egiefSlLkm0
eEGdU/EmXhs1L0//DHwKZvBtYum38unHmAv0o77X2nHlxJvTWyqOrJEAORqoRWLn
K+0h1pTv0OrRwuqaPiCKYg==
`protect END_PROTECTED
