`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bu1+ydBUYirf/NMAGc2UbfQZH25Qe3sNlkpq1pRhOTOgB76pCzZzos/ZOKpP3eC3
Dzl6tBlTk6q3iU2GOu1uxIslFtTUPSbbzN2owoYiSafowz82ZJ0dORHO5PujdbSb
F2TLE3fR211K6ITY7WQFOp7t+SZCo95CAj75U5/ANOtHF2BRZs5/0Kl7d0xVMYMU
mXJYbuhwQSav2eVdEPEeuZaPiz5pml/Df/W+8qPOQS+F0oVn6yMM63iiuAwWiJ0n
WF37UlchB2tzrJvBZo15l6d1Yb13iucWvbzl6TZgUzoqJvpDD7vYkKAvCEVJamsk
PNt1xeQmobdCgQZ/LehZdyCUxrGKdDemHLp7KZ4klT2Q0SdA1yuZKTzpT7C7+sfi
cYith76Ege0MgLRgsgV/Q9S56jVYD1D8P3E0QoG2Qe4zNkTIXh/3OP0k0veLmnFH
lewRq8+39xNaD765r59HPLtfe33PGfE8UJ0ct/aaf7AXGZGpO0171ST+rwTyztjV
DL6QVv4CxPa6oX+FjdYdeiLS005yarAnHFvhoMZ3KRQQwRBH+dy/a6UuXDHnlP/i
P+2I6tQoTIYHh506uZ8v11sfnqt/clY24gEm1+sHN4VsraZwt1M5UfILAED66UKy
bs9qRUNgGxQfmPEhvelT/05fDbzq1S1xltcL2C7HPvBJSP3IiLMsJ9JH1YcRPno2
nfg7CAb9XGtJOF0VvdR1NWu6YNhl2hpX0vma+cLYDZw3SrhrVgFckKuc5foqHiON
xn/sWylPvl6/c9JUgaYCI3QYLNR0nKKfJPyDSRch6Sm0T5wOxL2KqjfuL8Sx6i63
ybcP4g7JbY3zYmr54jktKqEbot9ZZ6UvFvnPdyTd6VBHhgk7XDemsL48TxLJ//EE
gZIS9/bRlNrGGyd61NFhG/WEQehNdNnNUuYQ/lsX09uBGcYw+pn8NbIaGLLkPZa7
dDi74Q77H/2EeSi37sllwGboN1Bqx1oDDncZyPNWUzY=
`protect END_PROTECTED
