`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7B8PyiagYk9ywBgNFAja5soiYDsCn98+zeEF+T+9K4jUlvZ9bRZhyx9kA5d4MbaE
qj8TX7M5WElkMb+mRytYTkpByVES1fsnotcIjr9UreZBbbvEH6ikkpIQW5cTOflx
tco4f20kGHMHahY3pqzqDo9aLo3AI9WVty47eMm+Nhj8g4R2r+GfA59qA0q6ZIwh
OQb4hePilxdH0tPkIevmDNPnAUttgKvB/gchVUwWZJZXEBTYZCd3pTtbCx7JwIIH
wyOhwV286cgNCw/rI+9Kc78wXyukWqQ4YFHGruf8KF8BXCl22n4P94QpCVEGQ9Qz
tVsqXKVOSQjFlsWmKK7IUCi0CRSfD4x3xkAk/94slQEL09Jy1RHyTzJh7o4n7yfZ
vIZdk7EpbWgPezLgo67bkIUS0LwSIEejr6WqCIjP7KQ45vhM30ZCd7aRZCRophNp
iqJkAK2C8j011YW0OTNsL/HR3Q0qIDwJmVM+M11HVp7nGWPDLEuCtqH+lFKCq29G
8ATmh3XwsExMsHh2rwFTPrlxLfkL/Ann6LS76NkTtaE+pCn35/8gIYsMZmZf7bs4
Z8+RmsHm9PHZZvGXI0EG+WO6Mvx00CD3RXrTz6EopjImxKyyQFkCtPKU8SojQIPG
4aJxsMnrPM5rlu2LZWd3z2VqyK2hSdW81FmAwTdHagXZwtOS9P0+ffNL7nmkDVhS
DmsrrHYD3AnJ5IXVbcKeI8A83J2CSMk4U8lnXWLDOcJ72pzgVNRrEnxNp1oxgegM
yrUMvh3QeaNiGsWn0aVtgovdDjkEhA3MAfL8MROI4+GFB0wJguV+t44Vwjfpkz6j
yYXXvHH10QSxqs0o1n5CH85d9CYMOxK1RuBNkEtVu3xyVie70Ww/gzuZN8CegJmo
kEzM+AxBfe+qCPOOkbmIWribX3dRXe8Gp1VslV+/SIanKdYL+rB9xd0xEOKJzhpN
ASMjU3ko6wsPTsXdYMeeZAyKQygUZfz/fVzY4DV2ulUxutrUjPfqUBXEds8VCdsp
jb5efFUL41XJM0aEF/GxnGAT4tGgDlIhIZaxVEx7IqF6hxJXIh0aKL/QciAl0Cc2
BtEuHlWdO3Mk52KJ8NvPciWLW1FS8b95mHqjhFqiIqRf5yKppmMwd7CiE4XIN4Q7
3QJWyDbYpTjgva6lF0fEwmmuT6egy349Xdn5oMV2jqS1+pGeZSwnAcxKSbX5GmbJ
/m0bZ2sxNBjNrU3Gl3wBI3tbEbvV+2YvNpE6IDDL8Qk=
`protect END_PROTECTED
