`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiFqqNHdQzU/JPaT9C/kyagYeF2kHGT3+iRTnYkbehHPxCFoJmW41B7Gc1RiIzcp
1HDFVepZX1yBwN4KbKhNX2tHzEXpC2kgaQx+66IseNskzNGVbpb8B/hf90KwRiTu
2AKYx3tVVhWhJarBraawq8t27hsaRpp7FOcEvLsgOzrhyfSpDmWpYln4aIYmEeDT
4wiImJsePgtnIGI7hd8q7IfcnV/q4n33okffHnLTsj/dqvy2kOLrAWBK4+XSz9Dy
LWfHWyLt6anF7kCoxjXlIxKorG6ptx7mkuZsu+NyRdBWMeEqJfJW85QJXPHFeFn/
KRT6dWKefP45BVRev8Q4opamFLCP2J2p8iKnnKuA37ukvYsQSRnYnianU2LtLGmL
Lv4wPfIfKwgHYbI9ps4K3mgYSnQfnOQqaJa7CVUEpMjI69OFF2xPgciywByoEIkO
7o8GacOI3U86xmBwPJtDsVQWZ8DbMIjeMmbAt1YOfvsjwdsV6rv5hZd+VdV6NDCk
ah9LTcD3YALdAWFoaeqs4uPhjOagweNvxRFY4WxT9B0J1vBYvgjqLZIPHdnpyss3
JIFRxtzjf8s9/0ldGEgphqfvPmVeDup6ShoM1YGQJPwc4TxAOnv3fo6lI+5x0G9A
Y7S80hjd6/przUUPbXFbv3cJpSr3tRl5iaFDJqpVT2aDlHl7sylMJDSOTA1ed27h
849hCm072IlQ1NIgKp4LYauA4Vv8ZRRRycgiZ+6tPaf/bqueLsHKDno17gE7y8yp
0YzvyhUpzJrIkijyMQTCaAvi25JMvVTD2mNOG6hKwbmdbBeHGEh4oJBnLopQIBIp
Ba6GNrhpaYNBEORB/NMY4gZFRgCRRAkVfSgw90IAPF3MQ1sUvEivY2qwvfLQfDhE
4oxuSZzDnAfFrpSc/YbaYs7PbuHXsNd5fNsZ4r2QMR12/AQvQIF0KQLES5Cw+jpk
/U6bz6fBdgTBtL/ZxN7VJRYjggh6c1m2D7jmsjvPNg3ZrN8rZJILWGe4i895cE4N
U0JaOH46EqwqirZMtw7X+iRYuMR823dXpL0I2u1epju/ZvRqBzYTH9ijY5TbRQOw
ApZRk1KdP2fTllWJ8rUOJNAqdV0+un72pvWflhriW+w0O1TbiGuLV0Y/J3+AGbTP
ViIxsD0GOdL3yX6dGWwH61QTlqTK2XBQ1ecNvt5E83AFr8ZeCNou6J730Jfx+q4C
1CwED2kJpl3qbz4NWT+9KKQ+W8VEomcPGRKQTXX+fLgu8Y5OdfDPfJlbVkXSJLT1
dkAJRrxklehAdb8Vq3oSukSVHZhoUZTKSfayLEoDk2363LTAmAn8rhIgRR9y7VzF
yenJmkMK788jfKFJah7Nd8MsmlRO8X65j/S96+CALOOhuttoBGePjXEICATLQgAZ
8F/SUY3tDZgxsGM6sdPJS2SvW70LqNpsJj2Ov5p302JqAzrkfuphkZwmUppxAdLB
Iqzs+F+xsZnUUc6DCORl34oNuAawqRFs+iqzYYo33XHL5aZZiR7qUrCmvd+wJIcF
1JAFX0N/pHL1btmwWtsPPn7zXIrXMpaAvofpg+T5MnRFNhkc4fSqGgp7zOGJCt10
cIRcA/8FbApDnr35WgLB3aIThhhnzRewY4m5p09c0e7Lp06/v6G6T33XFjNaTQIT
rEhStsjTKPbKmPGXj76lOuoovjzAzs6d6VpnQnRKJXqVSY/DKYq3t8HQtJA7GvP4
PqByC1aCEMQcBT7zO7zlEq+ccuDQgVEcJWetW4TEiZa7ZS4g21Jxb+xCSStc9Bxw
SsH/1KuC5Q0QxbwILf+aymKcwY8GEItCxQPDhIO0xDY87swokR8DPoXvxoiaAdH7
8mtZWN7ZNaUAOeRBGEk/rARqgUgU9BRO0ww1miSdKSl4FYQ9vMf8B/8k3iSv0guB
W5cpyLx4GPi/UofF5v6Q/qgkMn0he0TrAhimGXeOO6t/uqW0KQGrnkaicsHKY++k
ItNimLhzfKaNQ9UUpIsO2Z1JmcqCaiSm6H8DlHTKn9B1oRis9zL6emYuSyrjDNpQ
IrglXRNS/Dd8yA2k3taAnIleADi+FxxWJBuA8Q4OdSrh2sDnooA7EtBDBAnG04+l
ZT02+xZfsqEM25GunNliMz6HFF0vqZmYrw8STxHftBFlVpHXhBLfmm0+Djv+OzBb
Gn2blAHFz3D7VZ9r6W4nNbSV44s6YY1VfNcuH87q09TvEEsndBB1h0KdB2iw2L4b
en3H91TONyJKPcgcuBR5k+oQt4YhaKckPTalWYd30Ena3lBZvqELB+gkhPirKzff
WbQYHEJ5yiOH9s50UNc1i2p0dNpY0vqFD/J+AqB98BbrAeX29wVmPQR5uA6wOMiu
NlkQPs4c1UQyoITx5eITLollJQPsFCscwZLm8LcxKWSp/Du4uiwo7kaL8NiakCKX
8lztiByLcsrDKBF2uo2uVDYUHzuSn1umOd5FIiUV3ena4qizo4cJzXqqIip3jDXp
0rKp6lbOWA+SCh9Zi+n8IiTV0GM3tXG+w9itgu9pW6msGn5t2ujslUFK0bXfOiq9
/r7MX1t/Np2UnOVbL10KTGYvzHBaWKbUN7bAAMdMtDPiGOQ/EJEt7bt2Z1joyH/Q
Ha0ltTYNnzHX19UoYI/gV2fR0UyweVl7DgI3e1fdHcNkuCSfNYwOq96MRJFhsVOR
nZbwec2mFjZX4nZM4tylA/KUMjXjYk9Z6N5f4OQzPE0hxVmxdqpV123HYSpaQaPK
ny2n86awaGXPsPY3KfVddw9BOXVkeTcux5oV7g1teFqkEYg3R40fCMdeTJsrB43p
/yzbvxLp/HUGDnj3JWK5Jhu84fKtBMvBSu0KIXUJRKeIbYv9kjKtFKBkaTqg14Ao
EDt6b979AhHAErd3I4jfJYxTT782CsKPmsPgrpf73UJHz0dE+5JpaOBwH0Kk2YyV
K193Na2WYNQfo7fkN+L50ndFcz0SB4nI3xbCuQ9wqR91DqVCIA9E9u6gauIEg7I3
S6FYM/yXhSqdqfC5Bk1BF0AbKOuTXsX2TE8gZy45gBnYlPkUOChJYOglcvFeO44w
8mrMPwvFaacRjUJqxWXhpYZtjX3ZlCL9Hf2Hx7rtws5z9t1YTspu8T/lqdkyJIph
8H6iInJTk40zfyDLDZ6mVapylnRuohQHL5VX1XrIkaXzkNMFSZiERnFshOaGTjCk
GMsnD4AQ4DasUe/z9zLeksTLAcv7yCbCYTEPTLU/SevjReceGRODQRxB7YcMdKFg
kAfOTITjAB5NIcZYWgY+DVCnZiSoUrflJjWxGiwwKz1twuKze+/L7hdT6YA/4vPt
bQy9+i9gN/zlYvnahmFOO+UscJGk6m6xDvERJC3BNdVOQSF/RPHvlcCrfGA4SAC6
4mxkZV52+jDXBJiDbx1cwdwuZsMPdrbgwOpPk8jthxwWn/onsC1Wsf9dRB1VcMgK
EVDIniRpLp9ypna2rA/48j6TaSjcgqcSLV/91BoUfD3UoOZIRYfTvDcASgb7cQfO
Yiqy4krom4yYa63xf8dcKA5FXCqGRGL7YYDgECYWqcI55O/CupgN3IbgWu6ffAuR
Zzk1e7ZtGeGkCA4cjSmeXAdQ5Y14nLfnBohq97EN3Zp3ulpkj8PEqlvfj3HlHFBC
DYG81413qzeAuvcMHuT0Vbp9D/Qz0TuFEXyCrs4gQkP7d2Xj/vP8wX9yIcovIRJt
dTwiba83rP5r60PBe8CA91YmrhuP/2tSLZqaf9IVD6sqC/zd/smk5qpSUiPV9HWY
K+dZbOpVEWjuKxTbqFZkqh4cN0cE4Mab5yqNzAs52/WjAKG8xD6YadXi5gUlCxGt
C1VvM+uSVkwvv+OneIvwbV+suYaB2jqfu8HxRYS9XOtfeq7Zq5pdM+iwFVocrPcs
L2vq6Gs0rqBhikew/C5CFhMLHjmF+ot5SsmZxD6N8Sb5Vs60oc8+XU9yxTixL3TB
C2MJZ+s5gh2noIw1G6XJcXzZjmBLrX6NIX35Xt5orbumDhRqI0hKOGI/nA1UtbrL
l+4AeP8BZ43OlY4qn7Zz1TB31voSCQoa6Vb9ZOPD9fAKbPqZzgvtgbEy/3oieCYU
ksbjSLYUr/DFqSQMc9Hq2f7ZbxipVKuIMGcRGWUM1w7hQ+BwxysrYgb7Y7bEPf/a
7oCj3GRjrNXdFomXMue/SYV0h9jqqY8LRazVaK4qomVtC0Kr0vhk24MmDtuVLCNU
26Cccfm7ThkuYBHzsEI81lbaiw5BQhJCqc742yoNlcgc5RogSjVcZu7iubUedtqE
601p8iD7Ph7C/Xtl9kVA+NOrNk8y0g9F57B3chlmQEkEf4LPonvQBLXL16N2xKM4
3Bd05KL44PEcZmC+a+zcewC7F8QX3WVtzdjcnpBSW5njRHcQCxfzr5H/SyiBxq28
3xxYglkdJmu00VClfkc19KdhwlkuCRHUDVsH3erTgCycRdRcMFahvykLd9RVV+sF
0yhkKxX42g+BphGBpoqykRO+sB68YVNpxZz5ymfn4SpHndCeSu8g3VX2cZj86Fa8
FoY03fXKtZVfQvc2mcRn3myHAPo/ZxhskRQTndE73moSbD2vyJUDwBKtSp3rhIZr
8SC/Nz48U4ABXpaitQbbMO8t6AHmplABRF1PeBPcW0rbNXPodVGCZgaRGn4JsWm0
y8y9yVh9LxMJfsESbt6QI+sQwerwcGb7ToLBW9ebRQJAUXEWTUcwE2mS1tyNfRH1
0N7/1O0jip5V3Y+M8t/ilivylpnopprflvJc8+ZcniX44zp8Kwps5z0YLHKX04L+
ATTMXoA9Th3qkzORPK47dv/dliuqo09AjVwxuIqPwxvh46v5THHTGqLsqZMJN8Bs
cmg0vktQE4vpECJ4gMFlvHBFXN1Cc2pzIpV6Bs7MblEK05z9hM5j17OAtY4kODre
9V+BScY2SQv3qlAkB+t4nqaUXEJBXx1ynrZvekQ7AQLWdQqL/WFhlQBtobpAprKM
eTfVaiwrFvhKqENcOCFFSezWpqIB3PGS70vtAqMj1BYJvW67vDJuPg4K45uLhE+W
wiNWA0cReKLkB47XEHJMdtkdQiHAmUu2rTa0RoTm5gx5D7yh5yOR5xaEDtfMG6zW
EPuU6YKv7ySRCHKWAs/D1CQJhBFpfyUobZOuOTv3SeUpmXOd5OkDRw1+2180Ad8D
CLN8oFcUwy8+Seh0VLUziFLAh7zU8hz1g33bhNVjg1I1P8pmTSTQDCoVnsqnKZoU
YW8bBIJCSjO5DWCcMq9dAS6cbfmMdlSSkXtDxCe1dYlxS1f2Y9AItpJC3zDVDcO8
Gk5QDrEet5Zk4Dhdsr46uougXmQKToCoCh/UNLU9c5KEjz5P2Q6H+C8mefzkLjMt
60JWgvImKdxDaddBQCkhHsNQOR8PgxxOUOT4nWUyWFVrSlYwGD7siQlEGiu6whHk
evkLkAmNMD27y8+ZoAzholP3NJfN3AvUP+zv6bQD1lDVJeRsRPqdQhXwZbHVFhHa
rWaYJkSmV4ldc95U+Pu5PawmYrLHfqSwKArUkqH/3GFAeZj/PjBB4aLSn3swz+66
lmvO8tNvlUwyc9j5YA/lC4wpNvXRyQ1WTSbuxYJ9YBGo/KybJ3b7TvZ07hQTql59
+7qx1+/LsQpSKZPAQCdeSCwc1VKnUKjgDAVgJLhTuMxH4dEoXb57pcuidUDhZJPu
smTs8Co4nuoKCBHcVbKTU9dxjU72AJ8bfY/CZb7HTZLntQEIEKrIHDiiJlAPWswj
x3Iw6AMx7IzZJ0u/okvOju4LdMJRPnlU/0vdOqvF0hs7PyTIOGYfjsfUrTdmdUuy
FX10k3VSI0otdmYNggEspWRGBpw3zbuhS5KgbtpwZXlHx1gwKPnYkshU6AqdHSRM
KB5Irl2w0qoEsiSpdqRdpEW1dgkBD6ullUUwEN6RwlPtL4Z0Iug06GPkZpQkMfyU
pvqYJ9AtwokQQgrnjjXqkCQPTpLxoETwN3+/XTshwuRt95I8EAs7B1ccav9ViAH8
lBrbs3F9hKbIfhpMIpLbLtG/UJFa4fHYdGQm581ElVBBQWnbngw21j413jtREeG5
3XUdeRt3oBDUK/nqQp4elwMQZI3RBjyP4AphDnAYrOF0AgfUjusPocu4VqmfV6Sv
dSHwAAYMJxJZNpXYxcbAVxlB3iU9hfjSjdm11SX/alPcadm78xi0ACA9X2MzpoSK
B9ck6YLd5qJ9Lvh6gfXDXcW/pAgDTtWDAwzoH61FLkWe3x3w/ct0/ozDl8YX8pIM
nxhiM05Tl7jq/FWaOxtiilSMmrkeBZ2K8KKgakSo8tclAtt+kVUsV9H+s7ilXvi2
K2clBF5oimqEmkNuzuuj/Qr7x/Gf5jpft9l7Fkf07o7li0UauFdup/IxVG1EOWfI
AS1xecLVLb3iABM1ZMBC9mloeJmu0n7Td8BPATfJQacyLV9vaDVgVOkyf0107J+X
UJYmOyQT74aZpHN56sSW4tMof06CD6d6z6SBEF+e3e1oce4nBLNy0bjabF9WrMrh
oW0gS23pffCPie0r6JLuGV7gZLJ6bVE0szpj840OHtS8GGW0RxJaqPWODuFDLgQX
kRg4lehfnCG3Q5Z09jYnKiAPnIeu4Gpx0ERNd2igE5RBWBVUO4b4cfl6QUiPO/tF
/vnoWr2mfKsB+Xq67yHVZ+DzdD9dWSshZF9EAgiFMkNLxiP/7HRUFX5+JJqop8ql
yG5wYrRA1Ps26Z5w8OX6vIZbht9AnnYkKBdMn9VWOWAgJ/2OfMAj5MWkJOSvitmx
Jd5/d+wGn+rsACfreeRuXLaeZgKxkGqIQMOl70xgL9E1FvBr8xmUuJ4juuNCLJHA
nJGt3Nm91jZUsQazRzot3fxgwNyK6tlTtsq4xSYKm/kKh2qSUI+QdfXXVp8Fxq3k
ct/SRqLpF04fRQjbrXqy5MJNhrRV8Jk0Mrubkx4QEd83Zh0vY28KMl3qreEufOek
+iHzwbMxj8ktYy3Ec02hYShNECmLNSqyeGAIujb7+O5Uw7m2ATnrts5VR/y6gNvg
01ljtBWIfJNBnyQ19Q+71qDw8Hwwam2wnQbh6B8lFvrFaaUoccKWBxbFYt2xjQcz
MFs8M/hJ7PSqUyfGaasX5xDc3zzDWHIny0EeceVN8HVL5LBgSVideV37wQ6c53IH
sVjo8kHcu9gaUTLPyagah3uHf0zAyNJOfHspVmDYwiyd10rl8Bim0MBdjE6KNONJ
Rjy3rgLYaHv2KLN8Lm6gOqBa3PWUYoBPHSrPVCPscVXFuOyA7H6sduZN7T3Efnwu
uh9BTun7tNdpJbuD/H4DcH27ETxqfY6/ZIeJWeA+5NIEZ17m+ddGMLdbke18I1fd
TR/xZIFpS4v/AEUcT+YO1cxRzuEv5aAX1GXVpIPeq9wrA7sYfpXRTyjfCX+3GC6n
1+fJU/y+mfEbhtzrqZhQkxSq7GcZy4AL62m27A6HwFaDhFyGWK5k+/u6QpjDrJpf
dsqPXL/wG0fw4l20LGp6LF0VzZCjI7gNctmYYBuOz4zQ+Z7Lf6yWa0oytK5vZ/k1
Ogxxy+BZvMk5YjuRpf5fbtDg0T+/SeRTiTmY0OVzghlSTN0IwYzoMzSwUeQg/iJf
kZljyYGGY2XewajTV+1BCnxxg/SenZGEy2Qj+Xre8PVimHSeWa1W49XpA1ipmT/F
Ta7uvnL5MW7gikR9Ozn2JqP34j0P3cEd7ZoUCWKdThoTJHm4mxUPw91d00BbIe4m
1DtF+YrtR0nBptw1j0oBxkuopLznZulNTdwnRbVNKJwHppu5tlUwa1ym0bBFlsAn
tWRv06diw68IjQ+rzugf4YHxLKbRkUEuozuexiOkdrwpRDkEmYpSzAW0RFkW9hnZ
GSmlI6xlia1wK+AzQgW4JZLkQKn31nzcII9pxZf/vLNJvBmgbHgVlPIxyBsKkjDE
/R2pQ/E56wiQAkTXz3DYsjqcMmEmJvjs3Jft1LtfBnYOpGJZaFG10/GQPHw+NNEe
le5i4tv+6D+Ym15iMy6PTyjYFgqxdkCwnu4Mr27dxn8Y6+qwXN8Z0sSRol13zApx
KhDhOEji84Y572gF1odn5uRFNYvX1xLquDU0049CttQ=
`protect END_PROTECTED
