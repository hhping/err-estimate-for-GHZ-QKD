`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TgozqE4XeC8Td49LknVkXHnnXMMjUI5sy3O7oVMh81bLejfBoX7zrac6xaqPuThB
aOLGCFDz0e/bttsm2hnIq+iKh2QOJ1GLEzWlICmuRvmdxYflPLaaIK8aDdIDG70o
9jKnsMM+PNkeSVDHdS5PXpm9N1UXZBRR6qtNidih2K2mzlJTxDkOYCyBXaaSxYw2
F4s0chVF5P+dSCaDXikffC9Ot4f9B1/NtcwZGkPuuoGw2BWWWhjjXNo/Tzgkgt2s
9vejyjFfbndfpJRaxmeesEv7SHo18uRUKPbN0q8SuW6eqMzOj3eXbdnBAeiOf4rP
ldL5neLMeVR1Gr7kQWfbexaSBvw33WS2CkANyK6cymbCvjd9+tCK3J4J4SiQ0q0o
XXHQFwGkg1602cK9ZPIgVrYCk9yA8GqdDvDoolYWZ4rq6TgKgnMY0xF2JBYn1Dwn
5CKTfRUDvot5ofDq2Gw5T7S1o3cwj99oo1EvO2eNTwBLV5MlPxlTk5W7aSg6NhkX
`protect END_PROTECTED
