`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/1LzyhLBfy2uN5Yt2pZ9lMrt0guuV60ErrKyiqBfz3fHL66jzpibVz3phrn0SCeo
yGf6GBQjr44T6MWWkG7Us9Zm3sBQMYRENxmkW8ZSbpEw42fCk0/MgtQVu8B2YNaa
X6f9F4o+pWV0fexEQ9TGmgwSCwjPZWEhbAVv4cYi/bgYg00Y20oCSAOepFDI+GEQ
27tq33lpwB270l3503+mniHlbZJEYNYFQhbBq40lPqBVfitQRuTomAIC2+hXM94u
jxVsSSRmj0oDbF+0gPkr5y+AujF0LxAEvVhdjRA73t80jUSDCW2Qi0PbCEfdOKRk
whkkd2uFQQEPMhHfmSf4v7UXwkhP0m2Q2Ft2unvXSviLmgNn/YpDQm65s4oQvE6Q
G5aBourRtCHVh9H534Ok3cT6LGVfn2TK25bOrW0WYJ3PWDVL7sNMJWKK1eqeMcNl
sVTX78ysbzyOB+cXy+azdq3na1i3/Ap3qmv0XUZqnh1Ikx9XngVbPZ4YOTRO53RK
wa7KGz9YFLqyLcWg3xvcUNMBcOj2F9YrwgV+HsbzD0FLKW6Np+/ziH1wJjNjf+y4
DZVskDw9ybH+6brvakpyPVfuJTToEnqQJb0qCLVT4wScZC938VLNz5jU9qO9g20w
X3mFePG4M2Y4qO6Tj+fskVDNnWAcIbFCFJD13Kc4NS9MKTxOnddeDNwDbZEAQsq0
fWDDvAeUPUF3ehxLFuVY4JvlX0U1/7rlMgG9qth2tsSy0De6DL45hbL3d9hkn6ib
`protect END_PROTECTED
