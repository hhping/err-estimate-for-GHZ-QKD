`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/s2oTENMmHdmWGRBxHa59444F6s52pN4zoM/bnIBEcIRT4X7qcp9NQq7ptX7zaKv
oahy94OCZieE54rLborX+iVefjEQ32juEPDdD4nofvwpjQOah8ovwgDMvI8DOAzF
zPJqW8ptasJlqFarRxUKW0HmPzxWftDAbInJLalfyTTWgdgq9YcMpL9SN+jGH6TZ
6ulaWm9b0JFzNQCxWElTEAo2md0Bqw8R/FN3G7oHKzPvSLNeJG3R2TOrqNcgaxS7
xsfiSFGRLwCRxBK+o3NyR9US1IM2uPE1qr6+Nfakd/sScrDkFBQjtHmZjj4S2qTR
jGhwNT2cDVuw0xfgjElYURkeqCsfSWdpbqxAj4zQ0yjEOXFmtI4hHDS3fgEN8jGn
dOwOZPkvyVqWVUNy6uQsjwyJCteRmp37Oy3kMzNHHDropaDwb4f8oZrnxCkpF3um
d80xgXT+LVLuBhLr9JDTOi+pfnR0xdSmxTfzsiArHGBAzALgv8JRRozg59nq5JqE
qpeeBo+/El+E1RHsWBfDhHoBX/DTELRQNcAL/HbmsWSZJRWeITDbeaGPxcDxEeXz
hzvhWrsjyvadz0vwpbujb60DByqHXPHBKr7qFVC3li8BnNMY4+czldQ39yhekG2p
0n7jlV2/cMhHqgdKuYtPRMwlTW7dQ/Sk8OcZU7pMofSgmUfg3dPUYq5zkydXmYDE
OML20IY6aaBfJX4oWjdcZwPG8ovZDRddtgvQVpcOqzt2w/Go+fM58lyZMHw3z88C
drSgddEZwigQlQxxQwaK9w==
`protect END_PROTECTED
