`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ib1ysvi9y6X06WdvgSEezPaFJI9BY5n0xRujGQL0rpEvWFD1sQkuLq+QvVwR9MAj
w3/8mGKRRXMSPmv08gHSRNoZM9GVnzigArYPWjzPEvMsV87oEJfnNUFcF/Ccu3W6
CKPejJGKfcS8rmM0yi3t4XaLPIEu73j0gmAwWBhIoMBkORDLbxpTsbiUz+/kmgKf
HEPqFgxJjM2E6VzDC/qHLCbcSshS9KgLfmgZ1T1hGtMq6+DiDwKfHAiWzXh7f49i
3bzLsIxJNQKHPnRXj61ygmDJohYGq8BZSf9YEJa5Z4DS0RxZgLT2N5dHgw8Oi+tV
s4IPfQ8cklDm4P/5EM8tXnL/nxL+U2v0bfExfMBk8XpYn7m+Y5ahcnAtuvf7aw0t
VcU42KQqWGJ0pn2fS7vOr8od4Pyls8Ys4NrNczfBycRUyMil9NDD4m+00SePdAtQ
FC0fFDJyfd5e8lwdyvT60TBJW8wFw8wvmY2D99YNS+42dXtDDDKomXhSHcbSHjF9
5eCqA4zJcXMIBqQbnPMumw7RhPTwK4VkRaIN+WGtXUzCOi+G4gUqCJlAADH04xCf
b8rjY0tk4hbq3xE+skjchUuk7WcIRfT2m8FZCnRCm8hwNfOdOd76C/4q61ZAy8hO
MNwl7B9gl3iAcsxo0cq1iMlMa5EXipYnoLZDtdAkwSNfpIotiz0/ccBC3j495FR7
5k9nrKZ9dE3/Mh/HqW4Q8hy22jnn3nKq5zuVXL4IFXJdtKI+hNk05GRnmuGlkqs9
WUzhHZQbdrbkVVX2Ay19nIhO4P6CHFmfAAIq/BcITHqolTmyIA3RNuSSNGERQ9+8
Q5cX3+owiPp9c/wuDVVYG01DskcUal6fy3pv6n6EOeqlIQsE3lKLTyPc3O7dsgcv
aXJy1AqqBKOvJafiok1eK3/+WnPXx52mMSH0ONkk1RWrsmni/yProI7OIIdHImpN
wzHwBkMNX/VSNV/dTh8bwiPttu1x22VMZmHQJKFZKokSBo+swCNgx8aZ5yQkBlNg
j/3hJdqPco6IkUXD/zHBEZFn8mzMOEQgIeil3eeNF0Wo5YAZN0K3XKrSa4r3oGhL
9J8HNmPy2W7VIUba+erxLGpvz3wajYALoN8R43BrXFXNgPtnb/QFHcqYYRYw2pYw
q6hGfonPGznlgO9O2aLJmaH9T/rJJgFewj/3RptaSYMHuKzRHrq8tFJpal5hFTfy
uWUSYRoklz+klkk60MC+X33ZBPvAasAzGHL134URr5x+ofzszB9bvdY3sF9CQcIN
9QGrfStufQGmBJmVwbXTm33nkSXJFd4fIlNVJY2OeE4PBgBfKgjsk2WbPnGvgrnE
c9omvQrVaBwX18YbFSQJP1+P2xmbppiRsskt3uvQRI7f9LBuPhG2vJHP3GBlizOo
5GCqa8AWoWAL2/cmXKfDNe9QvBM+VOGGhgdsyj/oJKDk2VZICLvXI0WDx2U2c+hq
g4hnjUInKoKqtep6C0zhUtwuRjEPUo/TFTzdgjMySqraZfclpAMcZeu8NYiUruWC
dO000PIQUiLm3CLP/cjCru6vGgom6ly9fKyB4venH+iC9F6IuL9i7ea06CTWJhdR
ZE3Y3bqnmxzdr6HjBZYpy67S9YkriMe8xriBPOqdTNLhLdAvDo7frv1XWWu1Wdo6
TUOxbmrnRdP44L3cup4/wX+kp7PnjRaNNT+CkTY+Of9rfVXdcBB9/zftxXJ5isY2
8cuDyYbAIlg86eDF9rofjaHtTSqXN2XdeWZ0576aQZCPNpta5HthO6tReoRghcNb
n0UD5lAe0rI9MLu1mA3mfUeu8avIv4r4zwz19XQWQqDwB0DFrwIIrQdP7E7Lb9VZ
cOpoOThSZ3tMhscMamEC9xdpbFl+wHmPI/qVfPgaxG1I7p5u/C6TgZoeQGc8Blvi
zG1nVcLQFyUzp7rKbBny/RCbqbi6YGXFybHhB3LlaXI1pLbtaYIJL20yoGnZ18pp
EUZrJmWNjildJvRbAIUC/7Ietq3q4goY3jn5lv2C73I+tfB6JLkGr69y+Bts0tXL
Yw+hQ1TumwbBrKf+0XeobLvRAlkt4CAxzkyaaWiponiwwR+Zyw7R94Y7krzMI6PO
gC4anoLeSzSCZsju1eR+ao7S8loJYq8eUC9M6MGXxQFuTpzvSxHDFDIxPh8NqDgX
KIAnFFZzY5e7hg9LLcrbVPQwm6gy/7NQfMg7XDQDV4bOtQiRe6/eIx1cP4kdr31P
LhGBWc+0CtFuo0DklK50fWl0qb13KrkNoNEJNPtVZSNuDZqqZ31MHxtT7lJGG6ro
rx8iBrpsTCtcFAxRc2xHzAIHT9Oou+d60Q28Z6tRLGUwfa1ubvdBKK8jV6hFkxhx
ZkX6QQ6K0byDle9zY92kjuSmajPTnJwA6kCbbZeCr5r1Vv/6RL8K72Yzxxj6WpQv
G3iVqEEVPtyVGR+Yp7DVgg==
`protect END_PROTECTED
