`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQngKxVwXZbA/U3gIowtrFSoTimpQ1l8vDADfM8z3yAGXrq8bP2du9FsKFEhyL2v
bYJUZW1GcR0AJJOmemBsJ9fZyvIJVpLodchSKsvi/WRhQGFZjO5dpsq3zbgq0LbK
6ALo0ohJWB+qP9ZhoGqzOKkLLsoq7Uohh9Tj68kqM7dIZ8zYFk8DTqzpOdSOicuR
6iGdFSLu3nP0MGb8gjrBwwG81hOXfuEe6t/Z+a6IgS4NI5JbFEIdWE3GfgHNUAx8
8W6vTaTdRlPAdxj2QGt0AF7PE1qNmpg8K6sNrRoNdIny9KkFuRk8V3j30o9nyRky
CG1jG8xr3qS1OAAdPeesHmL/QjVZ3xtvel3UPsIV4TOSpbzFGexsCpa9mBedR/pM
gXsMaVvZPbd8cGeymiXYaGUoco8Cpy9HYNVMneg3gh6Q2v1PlXXMPwXc+8/XsGze
KiozFUDym6sVxvC9d8GIed1ugKLgjxQDJHWWZCIUN5wSTLZYXz7/+W6wlAjH2ICj
6Acr13d5iHXVrGBGwoYy76TuCoKu5VFDP/SANkpWD9fMCWLgNIo3CPph+8FnWfLV
QkuGu2W9kdarKMn2qGegPzzHKbliVqUDNKxbt/EZofP/fETA0WvCkDnhFdLqWBVq
QzNkxW2yXXB80epiv7HazBtt/EviIwVF5/dN9Lt0kk679Qd5Ir+vK97B3PEZF6dX
TQm2TEbCnibHG+Z/anmhmIQzfeU/QI+xPxBSh7j/wZPRLvjsiXAchU8SjMGDLlFo
5UFkZ+0JmSE2LjWyO6eG8ni6vgRqU/bNOyBsVB6RDDJn4CKEE0OjKvWsKXB7/du8
Jk3HPlbPu9DERSwlVFDT7PaQrB2B7y0pIeAL+wVjPfIqTJ0aUjXtYbSeddUmkTOc
LBwFmRcDcsXP6FKJiaRYhrTZNH1G3f4FCjnMgdeGHoR4PnnbHCFxDBJQgpwChvtL
HpUYITbhRnrhD2pjwMoDAPZal0DODkZ6PeP9rUyl4qszOrLqFy4s6/IOQOqFLRxE
Acq7fxtXq00+FTFHIvl/cFNh9tMI3mU+m+3ZZJWkx1couA5qhAf4P2QL3TYt1mIj
hlXYCYbR00t3qkmWGfNuICrKPjCIjN7JtrFdK8hLGSc4dELjgZbm2SLv/WF0r0uj
6FgqWy4kRdRy99E5nl2gFZl7cysMvGR7mUMi+pRrAcE=
`protect END_PROTECTED
