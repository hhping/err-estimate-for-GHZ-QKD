`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21uEl5Edngit6xqwklh++uLZ/5jR9Z39RE5+ttZM0Ej/fkzPyTURpPzRx72VRisH
KSHGXFRx272eFnw3kfabFzDZn5B6MOC4Bpvu93eru7mJ2g0K/UJpyRHFmIR9Q/yC
g+l+AbyVVVBkq0yzVT05/LOBxR7MnUcACMPOYvAjUz4qw4eiZxmccENv820x/VFE
941SjSzID+uwnaV86QAZu4niVcKZz3WcHAIe78ie2Mk4n/NX4pZTK5aN47O5VUsD
SZH75GJIbgzZFOu2r3Wvj6sDYQU54hq9BRwAcvpwAdVze3/RGvm4TvzMMS46/x9f
TpnW3ArW1GY4BmKuLaqrrNTOqB3zncqowY5/Od3c0utsbK0qsLTfMz4ajDDKvoOu
WtRRUEofPZHIiW/vnIFj/I0VDBCNw1LElwboSWL7JEXpbWu1YOPy97dE4HQP53ZN
xv7wrHRZhcGJe59kUBq+dhSVpWm8NDlcAgGdbDoLNSZbYk0dkqnIZva3Vx2jSefX
kMrOxnOePYp0xKkkZY2qPYzbMMoVFiaI/0lDiXGVHhAyZ9XjmBBGJo3fwg6hwrd3
QnjyQnz5iZXO+bS9JQrg1jCv1SD1l9aijRwMudvpL0Wn1L8+nqcowcK5I/Lbxicr
6ppSjdfpp8uZtabM2NAhwPHco8JdrTNrTM7P7L90Nd4mt7yBYwlVlZ2EJKhziPVC
ELFTLu+1T8KCgIdxHK545jJTrjAZNMK6DQnML9pcPvsgFf9n3U1ErqSJ2dnYxcqc
CPM0dEV8NBSSQ/BM7RMO+QSBsBRY6Pye25kpxmQYiHxFClEec8N/4aeU8P8Px7rc
I3BftSZfyeL/4skIEzE52zPUWSFc5mabSzPuTD/HRhHJIJsshIuHhL18aYje2X5y
MPt5ecE0QhKnyomlDEPF9W/ZKvVX+xIZbfvnEFlexexyz/zVtUMDIHMvzqPI2pQy
1PBjyuSRMjB3/A2cwMBNAmbjcmcvghkQj9tnxbiBzzSc3Cz9SVvbosKKF120/+vu
etiKxDb2dFmYI/OLeVpKfG6GMiSxo8E4B7XYX2DVUdRj4ejSohW66LPjTkklvGBS
Qyh0wjBz+yi9IUP2tEzWVQpoYkPVQLNOZ1S9TX6Pj9hQcavztvM86bH2cJL0xw+S
G+xl2eh5t11Mlfg22LeqUnsRVzcl831dpXdupP5Hp0euu75xHT1dJ6YlGlz3ggOT
wphjfKGIv9QSFg3yCCeqBr0jUHEm+otJv0Mx150eW2TlehzAZWr0g6VDYnfXwd3F
gqJJxDUQbADoCIecAx48IIxZ/8IMzlGcFyFDLiOA5rG8Ah8rWK0rdKT+fkEO6z9i
Zs14IHlfywVn4wIWcGAbZgk4ULc0Qrav59rr82z/WVdhc0hGlF+lJh6qRvCnqZ8Y
kSInF3I5f3Z2+IYeZKTJraXyl5fNISUpvk2BrixqX10oDKFfHpwRjM9/+ezLjJ1u
xTqmhonTz06zb/QqB8AnnB0KAgSXlovHR1A9SBzfuCr2z0GVOxW0OFkHAoLS4Gkr
zN0IYj/5aaQ0j69qhCADSfEiX63ikq9JsUchHoA5CFFlHsaoJSVuNvBb0u/zglMQ
mA5cTu87KGnD4hsV1KOFmcxd5krl76n7k0tqRwRCt8m3VTVuFy5/bcReqtT0MaSn
8f0rZVQxejmNKkC9Y8SV6js5ngZQwC89L4AhZL6o0d8=
`protect END_PROTECTED
