`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmiDOMh9FpAJ2DQeC8KwVUEudgXux11zTRz82EgR3Kb2W9YIUtyB72vQJ14BH4aI
oay/s9aE6Grb8qXCrOP5aJp+2eXTmJvDV1DAHAlCFVRVwf5gL+qtN+S1B1MUGCo0
A2+k46SOhABDOowdo2bXcky4+88TJaoQCtuEhnpzNTNkPJbsTBPSOaQTcKNKpzwj
ZHZsjU8v642GafTGSAjYdrqdWSAK3B2b49NR6ZCVTaPja+CfqIy+ntqnORi7F6GD
U0DeaZ38EnIqsZLGRT+T5IiE6fyB2GdvIekq8Ry/DT+PQxpyu7a2Zhs9uNyN9l24
+CkaW3T1gPlz4AGtXeITzDfStjAUzhtvzV6Ieq2S4JwwCl/W7Fx3wbN9GhGpS1ql
06hYgdxgOMvqe2ISa5Dfuu18uPYwvZrFdUz72aZpK9FAxH7UdL55xP60z1xS6wuK
A2XMCilRzGrBVu5bvdLafvHk2YAqDpUKbEvY+Peihmc7rszdFUBYa8Kk/kvs+vAI
j3YdPZ3elYv34EhdVxk+gKPXkwER3ez1JAEOCNSIjFPbTQfbNxqMEgS/1dImJQO4
XoDColq+wKCojBz5Wz9qKjvOQ7PCKVRYSHOAylXBwcpy8U91jK7I6BAmYKiUux37
`protect END_PROTECTED
