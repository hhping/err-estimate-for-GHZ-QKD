`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5OnBJOgPB1bqfdqe/cUFkaZ02M2qaObyWnhen8wvxDia0njR2JKO48X/A2OP0Zz0
5Cywk7KoUvniTdhunAo6uDTpSf/zAnDQMFCGxyIsVNGQjjehaHxmwj83lEB9TRWA
SNa80LejwcmIwqJqBNVb9wRjNpKyehzfMSxkgb8pNsGO1TibI/l6HBw7WXoczVfy
hcaIoMZUL6eRO2BvOE6/eLl3K4kzMs8a5xlLlxGVwrS0SBqd6/3E44Wgr1AJ2Ynz
CioQlSj5GJVpot3cLR/yGLcfgqqLAVOXEqBnaLkvWO7sS8fbJ69iaksorNpEkWQm
iOBn+PG/I+GAWN15tlSVW/SXrktVcfMHttn/dgvudUvbOiAzbr/1Ib+V7ZiEbjjs
0ZFapGpkHWuLKhKc2rKHLWHEnH03UhYl4Qtb91bOFauIbrDjiAKVJPDAIjlxXSjh
vR8L1VJmBTvt/zyPqXFcrYTNnV9w5ItwRyRbRJhUywjrY5+U+5LhELlcDLOd/JW2
H6pBAeRajiQPKNTMIxayiLEI/BzgtcSzbZylWBO+Wg0CVLeAPcQYX1FXp96yn/bC
q1a3aiGqd79BPMUVDIQXBgY4/A7BzebqJ0ZB9U6V6r1Z1mFu2K9ENGD8tdd5IzX4
mNppjmPaC6bUnYeiK87CJFlnXbVPCI0Ibn7y0j+I9eUYFSAiIQ7B9YznmW7bjkWX
X9ZlmzNKSJQwlao9WbLHovJzbg4NVajlfXAj6x9SDGKgxvxXPb8MxSspPFYEGmOZ
my/0+cHjQC+k18jijQIs8OXHNm4SrfzPaPFT5f9yafEg+jigTXL2F8PLeGvabykv
A0jkkiDI9BU16phD5bahiyJLCc1eeiI7klq60uRvqfyE9hL2502kgSTCiWkAOJdp
kTq7pdyaKmPbv2djkOlPrngxcIXpGNJOg8IHif4TvJZkvAuGKJaXDMRVuxm6a0Aw
zrzYSKLUWokafEhKJUdJalzcZVciffri3ItUQAHAj72KqNMLrfx65bKtSVmQPTqY
40VrNOMxpe6R9yZFWXtubVAsr99ilrQXXYeWawSMxd4PA2RarCeJrBij0QTf49pg
kS6LcOmaG2DFPWjvbu0g+qKtAOYJn3T2Z9h+vweAC1vM3CmUkwkcmY0CsQG1mrBj
Ka4dv+e235bwNMq/7HwLgH1ZoHSTOiQ31BEy1NVAKcqt8HKphkPF66WNLMRY00D9
0nQ2OwQOmBpTxuIW33DVT2cslZ91LugMuvIpPBxbSxeFJ+AJXvHjK7LXzj64tjMY
H4nvq0XJxzER9MmJoCWvYfJYRF0aR9iNmTYVqsQJHMQ=
`protect END_PROTECTED
