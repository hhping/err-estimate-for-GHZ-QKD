`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fHMae33T6edxXX3AqsgrmynQG7H03GAPD+LClG91ImioygMBRO++xmbbZXVhi76J
9JsvNQuQlGLi1aKS3Yl4yrtip/+1AaYvmnDEi1c5Lac5cAO6QINSyR9pyMwFcAM8
abt42Ca5Ohh0IH3blIRvzD9e8VUl/k95hnZjnkb2J70ERT1WfIRDYQlCwGMUBDmE
mS3OaATqxakVvjYeK6Ch7Zcvz0nn9r0yaB05FM/hSIUFadic+mODA3SWtBGQFYqQ
OyMQyVhfVASO/2+WIr9mrKucvzYH+IEPZGUskkITESWb5en0QsOvVDapc388IOZ4
Kkd1rt0UerZJ6t4KkB/KEi4CaFK4S063HFyntg2v37nZQCVLroSufweMiabg2TXl
XlIrmZI+Vy93PgsasVEwqZupebAktbmRyln3eeJIGyGwH//UTcdE1I7qh67FYnmV
8C6M5gmzTFCDtZxqjAonQX6M3FcDOr1Cl91qKOBtEVfq5l9g0dc6x1sgIbMTHO5F
vi9aENW6lSbwvM31yq2XNfhVs7afX94NOWqA0AIP9ugMhu4M8k5DmCJzE8HhvYl3
yVjuD+YtB4dxikB2Iow9DdS3sg+gTYL+5AU95x2oAJs90pwbcSpfWrkP53LY5tTt
9sGSkUaXGUV8VknUWU9z7XN5316G8YPMZrstkyWEUxKSLUbrUP+5uFOFsu7l/Ffg
9NeClSLVB4Y8Gmck2EXHby81VINaHGVU0MCdzd0fMoafSAhntCvpZMj+bIqWjgGD
Msw/4Xcd8dN9u0/CSq4sU5C+V84otJUB2B3p5e/qZTq4d4iNYFDW8Q02NFXcaORD
skyJA4RrbEt8Fs3d3Ii5PscpHs3lFDIRGcIabjRBtwZFAqHiYcmgA15s+WoyOiyI
fL5j1yQrLl08J5ePB9e06R9/1bkQr7pPPCWbPNBMH0qINmB8bjlZqu+iDsnOU5de
vIHSbp2xEmoWDOXPPn49auMlaBkotYBMCB1yase9Mu7rk+N8BULXfQdjcxZRI97T
`protect END_PROTECTED
