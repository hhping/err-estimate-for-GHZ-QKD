`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8Vsa9Kpg6Knne4aboKnn1AQYG+okp41QCnxovgeZde/JiSrXOB7wDrBpjIRmLma
38tqIwGInwGklrNztiB1+eqWxiaGWfp4q85540M/W6FyAHunRukhjcdnIP+v8Xbr
JWeftfsjvJG5Hmw8jJn2F45NWz8GtYiLgUjcssIuv4UQA07k4I44EznBxuYXip5c
lHj266RIjQJiscohxaWd829caKb1xQ2G6KtTwx1/P7yE0mmY22u3eUz1Ri2MewmE
pBQ3Z32/aYuwBegri7Yb3DQSiJSt5inX5M3XBjnx0Z/GCtv6GUWJjKLqCWZcoojQ
3mLwKaidkdPY+qzO2py/wyh4LlHnWu1lGnEof7qwzc7SncAeid/EGkhUK3JDKUgY
GaBaxhFAACZu+svGKQ2xu5lJonVjvZvUgywjTgH7D4aiMUD6AsS9x4K2FwzyMVqK
7jfAQH4hQpITigGgjX9H7Ukwur3Mt3vEyFYdS1zb5/nZUK7hf8+FqCI8f0RoO9MG
8UojJ2ttXb2JlWfpcAq7h5iWacNsYVHZK/0nOA0P9uEbaRe12sFvjqk12GkA4cBc
dhpxq8nNn2AUScQKO8yB/YQWXSHpTIBbGqCBYwnQj0ALXAE1Ec5Yhsab326GGN8p
NW6qIE+dJiTr1q0pqpfpzQ==
`protect END_PROTECTED
