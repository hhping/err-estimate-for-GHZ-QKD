`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdYTe8UEJhQOWm17POrnav382uyjQLDcaL7j+NjmVHmXde9qis1GFEqRVdLOdr6N
1bA9TRJvNbXQ14qp+jWZxdWMX+TqldSFN3W7AlLFDk7vEwTw+TvRUPbGFGuo8b0n
n53zrh9kuIwdGv75gTcf577RLLHYRnyvfNOv1mRHF2QHXS5yo2WQxxuIySX0meYQ
C4ZNrFZddfb1f0JyvACKKy+Ed9WY7loYfDbJ7j+yZc1NWrkJF5NlW7XQd3t0Ymp2
1Y0WQbCKE5Mi5jSyPFVU4AGVk/NsXjmC9JxFfqIIHG3ZjGoK0qvvgNiLKLMkAXCC
idMk1n/Cy5UsgYE8aU1LUEa3bn9LviZJBHeJadRF96q/QILqtii3ytMZcrgmx3Hf
9YfVUmD00Nc8YQdTtedcpvy2u7MoG/u08ONCiRQZUxnUHQmd3LEnUB5+eOv1BYzw
6wgkPCxiKhYjBPERYgXGF+xqI88HlcCdZpYWPMV8+lZcamAPlhck1LvWaJzRwAPa
KqHVYuAUb7tX0bjR2yutLQwzSX+WRUe8OEIcN2wAcsXi5XsQgi1irZuhfJsHXYW9
5NkL98h8WMs9X3d8VoTRLT9eAoFJnnRmMOjJV52jwF3Rhliokz9/aCBoVJSs4X6m
bCwkD1L8f3tDKFYZCyKgp+6m7r63cpMcYB799IlAQLHooZ+W0IwfJOCBzaJFHHxd
40Owe5gDo93EVcFcShtI96dX8EWnRK3L+n2AgBMSxwmyIvBGiYgMKvP7oryBgaUT
HJxj4JlI5s50ekQslvrEd9rlIJi06DRhAR9YL+xK1KD4qKhy5+9S9BCfPyCIJq0Y
X97MWQ3n+2ltQXvlIDB2IfFelG4OxDF2XPl+fTkVsCTDgKeOwWyiVZtHQK5iWObM
Cbz7ooTsheY9OiPoo6sXJ9tXSYx2KBUNAcoC3lTARG9WUTVKcUveNXyQCIQi8r3v
U7uQxmKLCJbmrti4TqzhfqCnK4sSQdbj+Nxl6mg8ROvUIFARH//5NtqT+pkvFoMK
xoP4q+1n4oshHQVYeS57IOdcL8YV02Lmn6MAMmbSPyMi8SSRniqY7/lrhG5nEJBE
tryb9xlfQ4gAWDsi6JvUP+32wrlmQ1vRsAmgdRSgea6ZyIOo2Gw+fl7KzWMhDENj
xfUwwzz9zxPp+3fLSvwGFdy+90BYJNsn8W7KztBoI3oHqK+Nt9w7KDg44+XFkuOG
2JVVqvUj9hh3GDFUJGJhpp2xW+kcPzyNY3LSrKaP4SAa8F+6Az58sRttcAX9xNWd
ANkFzhkCxdtwhQ46hZNNWLam4u4AEV5K53/05aj4yaK+QUuu6eUDLZdsIPEKC6E8
`protect END_PROTECTED
