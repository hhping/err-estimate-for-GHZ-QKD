`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAoEZBpQCR4deNuamIOYHXVjOLvtb9dCeJ/UUiB98fWvwK0Fmkd0wFarZaTC09eW
VHGpL39A+1HbEM7NXdqzpD/Alu4OpYXGvRfOt8MtlUranASehORimHjEATYfwofU
a9Xp5epCGBEbeXljDz+p25U0jjVwIv9nA+vd4F9hYc1wcnfyXdpSnPkTKWe5qcKi
yIoDfsPh1qbs0uJAvmKj4C/NC8lt4oyBDAWNbISufQ5OBDumaeniu0jlr944bSqe
hrRXBSVld2t7xoypFcxCdncCjpt9aH1WriTgusaiV+5yX8jSBtRf8LmsQ7tVbwCs
ZjCItul2hgXPglOuRuh0rnZFf4pD1fULVF/yqeZGMae3atseZJaTxXWSpGxhIZJY
uQwqpFI+09uaqyWKij3LHC0OXXbi8mpDLCQ/Jaww5Y6FEYxZpu/my68ch49305pC
rlyHTFLJ/mEJC/5ui6YIB2rJL26iHZQBSEcgtNOUpKSR/fddT1RIgt/3D1cs7BK9
e3l1faw5INTV070Agp9zNuAslEsHePi1gwLp0gCQdUxNNeNRxmZ2ZgJP6QUgauXC
l/eJsFFmrE9Nd8++ULhopIxGcWAYHm+H28NKbWo3FV24B4P153kQK5ievl4Hv7xx
OZUruG/ESnkRKj0V4OSjIAxmCALwFnK7R4kWAIdeg/4=
`protect END_PROTECTED
