`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTVyM9ymdBK6xNKitlVbcxIs0+EzPTqrtDlcgZDZWagslKGs6p/y4jecFcAIwsa8
zheyVtoTWD4hz12mjEOgv4VmjY2d8mMiFeFKwAxahcKIECFBnfeWqejqdAKdqIQ/
ZzT0gBamIWc8aCd1wBcRQ9QvKy2g8107DuuUBMEOBHelEF2nkuEUTIPS7KFLjsBd
hKG1ytMTw9OlYj2jmvnynQvAwVSl3SdzX39b6keoJn8s4LXRbpm4XCkcgy8as+PW
ELs/ikPgmx2lnlZ9aFPSk9Hrfv3OGS+7BegtMggmFErE/aBcDUJ1jDlp6DnOJSlX
c8C6/VD5BQtCgGeTd/UE1OxujO1avseZVs/AruhtqRg6lPIGi5Og6dNrCsnjmKSR
fELd+0bOE49SxRW8dF135CwRX9y7n2o1XRJpLvkX/HVQN/mv69s5dP4BdHCvdJ2H
/Uu9N7BJOOvvmck+l84CMtQ4eA+bs3v8+RYB41FJlGbpjVEL2z75zTDljEE/0/0l
HNNIRF2K7r6EDZ8R+TJhRSdDEOGC+InBcLcLP6xlNBR/uafk0IlFS1qgAgEguuuH
KFJOKz37nCkuSWvQvhK/oZCet6Yj+TXG0lXVYgxLVioyT8r6KFukLT/Tubqb2QIZ
Nix6ISZzV+PNLaxWiRUnaVH5Ec8r9WFeynijQt89qci3kFZZAuQ9TMLrPoljQBtH
Gzfgn5DNO7USr6WU57qaqYr0fFPmt+L6X20wuJ3+GmVXUyZj0bvqUjudyd6mCv/q
InLP64YAaw6A6QnxOe/BXvxOA5OwOhku3t8Z2XkRv9g/u2P7leCdL0jg6/WWdYPF
nzVQj/54jnb+9bkfuIbFhloxABGzj25Y6ii9B1hx9MoSGVd92jCB/Wzjpa2pJJXw
dX8UhdkSrrVXJaXghiYUKHyCQ5Zntxdva6QA3TJPO983biG/uReO4gS8IK5fodM/
KGx3plGufFX0tWmPRNfHIwOyjMqqZMcHfa/6Q8AHI6E=
`protect END_PROTECTED
