`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74/G8r5RFR8o0BEVmOyuNWlf/J6Kgpq6o/uQ3jfxfSrz63rcsgyoZoZ3WJbdomjP
gYeyrnHNjz7f5eAyzQNarslSoPUsSvY3p1diDVrOIBBCsZ/gOf1J6ibJi+aBmYBv
xP5mzP/Vl6vH+tlQHXLKzDa1Us+8C+0GZPpShtBfi7/5ArBfYe6Zbi7YRc0I3CyK
afEkU1JX7Xo6dR0G5VWn/gnxk4zk5lWX2kjXEX4oQIr6bw7kz/mJuz1YZoeij6L2
AveCvFJ7yHliq/xOeH7gXFX4hcgo2KEST6DGK/ceG2MeWJ/3glJ3W8Ih9/Bklj0n
D3T6nCeuJkYMLJ1JsachyCXJaGWSpWQETeIb1XyN7t/rZpSkbx/x0DApogMVpHM0
lt8OuT+NvG4HwuskMwIuqZYhgCJMD57X9lhCZb+5vwwimbMFelmlwL2OYd5EdxUO
5PYBNjCwTt7sNoLiYlLgw/nRsM46cm8OVpyA4JN8WelC/no0Oow0xgZu+q6yCSUm
rodFbpbj+100LbdDyxDqIAhoCHcUKXBoaikyqun6uw9EDt4TI1ICATL7LtqELJMn
q4zt+t7ku9GZGkN1lV86aXrXGYmZUlBiDecg6jwL9dUNRyE60Ha46Bw4QqyjinqW
FDrhv0fcDIhglxK1zI80pgE0A2iut8llLS/loySzukgCKW1JdOQGqtvmHkAiuq5X
uVK92xkAi8pvgda+ax0nk43E7lM4HB2P8HzDDOgK9YW+fOhLRWXyiRlJWxowGaMf
wlJUEuiCgbxbCLLyT/n2wJ27aWww6CYcFat1DvCnPaEr5SAdj5T4yZBXSsPkWZfR
TKmPE0TPhlfCk6HtwI92EYgH82lUEvDP3ovcOkYsPEzDvQE//ZwQW2LKJsalpT/2
0r8mZN6vLOMAhk2GVYr4jtwYrLvDgY9OyWkzyPqtRkZJfLGZNKEP1MBvm9Fb3WGY
l0UdhKxa6RpageP8BrG2H+F8ONT4wNWdb5osaqzfVPBsYr/D59Ma18haMelorXao
vnTnbCAMUTgp0nMPhHQz1Zy/HffvEAUTMIbyuiFzRO3lJ86VocH39R8quiZd/teO
9/PhGnsy6wxZnMOgqnLmKtXkJ4V0Nm8aqzVUq37uxtHhLjLlsQx2dn1hUqt2n+eP
PWGAxbQhoKuYz2TfoRQXwkuWuZxGdPaiQEt99JZUghXHHaRbymXgbKgVBKoctZTm
jq9EJ8my8v37A/0Ht3dB1QwA0AWF1HU0V6GjECI7fCw8aqP26DkO1lx3ax4+2j/w
M0UKtF8EFithX+upP6g+TApHWWn4kxLdBZ2LMVas/85lyUr1PuA75bfiNJFZz3mf
KZ00cmaQtONivj46rnDt/fiW36Qh48ohC2LlyfhXMpU0Ah0+AOR3RMxFOyGQidCv
fFUKhdqx6wPw0DGEvXjsnA==
`protect END_PROTECTED
