`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QIe3lzDwk4Z1WyMy5FwXQ22oVBJ6QGm/2LntIbuJzp2UxflOtibaLuhuj9LfsutO
jqkPWS5f7p2OmTAHQcJZu/62C2q2dkQJtiKXVQ4dLhJ3buK5AlP8PdN6ijwlchGE
C/qmF51x0RzJwcLYWfqDuTyvx2u3q7LkLdjFxW0Fw+UyJPVq+dZU+jipByyDjvoZ
CL7lG5I5XvJ1Pv1/VgueqSCD2TDI5k48fiHNv6OhoHI6+fvqvT6N8rVsX0zCJoxZ
zqZJWmrf7No6Uu0Bu0Bz4OseKS+zp5C4GTovKPMtn/jbfayNkvVPrmOfyarkTnXw
vZXJvOHAKBsj1rqH7Po1xW2RJTFiVUaXjBKgQAgKy4wF5JV4WAtE94SlTcU+4M9W
gLA7zY2Zb5FiyBj96jMDi5GAYKS8L3dvKzg15if5uLfZBT7sR8+q/AbC2OWBNoOK
Cs496MZzikHHaYQ9Yz7RTFNk86Inj+d5BfkfkxzsJY/Gm0SISryHGS7EueikEMCW
eCxgY0b+F7OYMFZ5clo2Ag==
`protect END_PROTECTED
