`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FfB2qPy3PoRHFE4Jl26I+ksLnqpP1bVgIYcd4k571lYykNlOvC8U5UVZ/+UO/UB
c+Sa4j4hb9hETvEefk3VFFV3wJQZv2numqQ8QiST0klbs+jOUBu6cdF3QOJ9x1vI
NxPj4aAzklj4Xar2KzA3xWqUPB+HbPWgy7WrXx1eIpsN5DLf0NINaH3m0yoODT+W
LpVJFlWkzzCg3Z2/dZZTn/9vy0z/fcJlJKvo6me6Qv/RLjC4/vi8o+ew6vLXBwxy
tNgb9qM+KLhBGAL0CVWeO3GsEtTPfKWdcHoZzI8DmczGrLjhfHCG2318O+MldSIt
nEY2VpzKtKlBMwOibBMIQfz0whFHxxzJjW/sAvJLuCU0NVbxYnxbJ2hXyRMKuMF+
/UstYiA58CSY7KJKkL7Tk+kaeST4pHfUTVT6VZ/cqlVLDz+aTFu96AUCJttU+ahX
35xVGN5WZrbeiIRR1mwtLedBXN/Fg9gnnV+dZcK+CvRmsYQhiVoIx0TsNrXh/UYv
Bb4vTy0R7dkut6ibgkp1E6VBAWhqYAwV2X3Hfdqv0ADm7mJyNXwq4jM662tWLD/O
wQcTar0uzmWK1OnJTLXQTKAuOU+VNolAecBj0ot4X3UldeYfMZYvLzHGNIZ3GNOG
gBYK/ZuIF2Bs4t3wE24/3z1DursqE3HcdhNEZJtm5WJPGpj2L+PK29ROSkgwFAa2
yT1bKguAvSjdaqaeVj0VdaHf6muLJ80Xpo9c42ZloIjOftELYCOK/YW9nxSyg0Wb
yHEAzbpOP1skH7i2XU5NGX2mtCSgEpulDpTYtEIeKBM8LMxgaukfaWWWpArs0Yov
UrueDjURXAoyqCZcUVqQ2e2qJtl8OBiTNMHKm4b/lUmKXPxxOuh7ATgDABUotETN
C0HnTXaPPrV0ZTKJ0ojzioFblvbKBsv22AQcMQ11iU4HnyudDIZhfuXePcUm2kFU
nplB9Mfy1D1bSKawOFIQiRRqPM174C9RgHwfXjGgqePhPN/x5e0MgKIKX/76Ck78
rPdRTcLrIT+LNeUVsWg+fWSrxAfomjpG+Gn13n3HqZXWH0vFPFxhFOPOmSCSNFL3
5hUgWHdzyxiWYQU9DGiTcm9T/DsKuEsT8v5fdeehxXc9noppu9idsxvqeGDCcG6F
FrhbOUCAiggT0KJboYSbH8/COA3rGK5SYmBM7bQ9AbqqFNIUxkoR4uFGN0NSm2bU
0nPDmBaH6t+vvpSxR9UDLSc0RHvTxIIF7dCBnneakvGY682WiDcP9Jru7h7wHRah
A54FAu+niD+lE+UWaKlmLLH19hCtaiNY/m9FgaArSGcMRGWgqUsJUeNzUUebUXTE
133C5tI5l1xBqRav5Sjv6GJvPzSAqG1Z+n/yqBqx5xbk8LOU1rplVV2VL0LDIg+f
vYAfEYAYKQmlPJwWnzxRIKF1Necboiopf8fIXz257/aTHrvJJnUv7JgMshbAI9Xa
lcqei3GXz5+t6OW9y0gj2yaY2Yv5RXmBagTCNBBKkqjFbeL+CkM/F2zJ4cZ6BVkL
N9yyTH8erCxhKr4aSc4FkxMU67eBWKDWsps37hGWmAl93c+/Bb7nWnHnESpOEBQo
ZQlLpWhp3oPDxMpD4C1e8MjUu7TmvJ7xePjlcTWXm0gvyZUr/vxOlHbv292izByG
`protect END_PROTECTED
