`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VysjzT4K0FxkgAvWOoLBikZYK4gQByQ97TrGqONEqY23hNrtyY1oCNL5jrdem3ge
xCQP+T7rWfk3RwQpGfEsmt9mWah9/OkeiQk3pKqVW3sBbKVlKCqsSz9WdeNNJtkI
kJYj05ZOhy3e3tdTW/j3JKPh8rh2I2ib2DmuDeZxo+hst12tW5JgUdU2jazlT/kt
OE7MXkEAGRI1RqOQRxdd+Anwab1eq4eF4GL2QZyMhEF1ViCUscVyLGUXCYaePg/u
9oAYVvs0mVt56euGT4HA2cvJGcRGsm9KZJwLQycgWJdOaT5qEr4MvsMlj6zKOurH
kuN24qziq1CTnkB6mksV5AVQp6nmbMRre18urB3MjpcwlnzPMyKWJxVkAEuMgo4t
OcY9LphjMt9VC2bdzL4dU9Ol/0QA7iJjy7GajVY0MX6wXQytiVH0E0GSKoXEQSO3
x4P65TAhhevsl/m/+EoSYlCWDWgZo5ppvlwgaLEAuAhcDf9SRnFpcYWQSkTg+dGP
iyV7ZcIh0PEzq77FEQBXUev6rnOK62Myuwwc/Wg4hmZmBna31PcemZF9ov3BjY+S
xpJdfS2TY2oDSTJouLKdmP68e9Xaq7qOhf4OlgkbTE2plk7z9ztIapva4uvSqJB1
xixIuUtkvs0i6pBDU+cmuSjUVRYTtanz9NK6Ix8rzCD+2JEjnmO1K1gEXHX5fgx6
i1pL+lXddzKhTjthoHmxHg2gbRn6CTn1jTNz9h3lH9YdwUrAWz7Vw2VEGuFj1ldp
o0hcDJIXDF5QZ8sCUPjLav9/Xi8SharOk7mIjvl6+E/u7KSs3XL/CKY0vpXamKeZ
/xmQdzDY9/hjd8twfcfOvC+bXkr6gvx6yRgrbvUNRN/VrldYOFOZpsGgHA/HjkiI
PH16c9+KuHyRn1DGfL4zATU+zNWBsXDSJtfStNtZ+GeeuOiY3JpAQJXHHxcf23No
NJdaWgxFhvCdHJjyP6gVTt3W9TVmnI3Q/S1w5mxEOmjshyJkjK7bdqIocW/YZXpF
R5KCxTlF5yhwjkSjyMobBV7aXwC3aE0kgqQdpwzVp+T2iM7IPekpr4LdbFdsPH8I
F0YXCpGJwkLBlWt/lzxeMsjFpc5KBiruynrRnQ/5klX9NvL7JB7DAWO1sAP+D9KI
OZWMmHHRlbxrQKd2/G+/jTEaK0PxOo6apCX0HLiv2IPjAgTUOh/zZ6Y2I8YbHL51
QY2B5+2cqk5W+amrbf+cGdlM//c9xlhJGxbrRN39xaUScy9+Vb/HsKksen9JzwDC
Porl9dkPLQhCXRINkuXkE4Viv9RLjiHxxao3mysGfAibRiXs20c3eWAPaxOOe/Ef
D9XGM5whDtvoZWhoFo8wDudI9jsTfhYgkGZjFlchxnRdg3sl4tx0JpZfFhX6HvlO
0HIEN/zIH4oHn9SoSFVxtA6RY2kXioFiku03t7T8pcM6PaBSxecUYcJgd3E5C1Ea
bSBX5QandXsnKWiL7RuIic5HVgf5YKtKAL29+8fSQR2f4NznRGscXlr9sWaMFdYB
0iBQWs1oGopAUHSxP0iMCW98xIKSiQACrYE6Of31NY3gGBNrwFiSE1mCIsD1KZyE
IGS42+tL7zGQSs3e+FoL1J0jl6yrAiQ76Y17N9qh1mhS0XBt+6j2wT/nPrqbV9w8
iTTng1B3EfvroRCGX6QpWqYxa8yKAkx+4DCmSldEb7LUptfX1TuscomAVvrIzcbZ
hXDVToTeiPq8BET/JsbBY6MA14piHcbENUajGyDzxM/t3RR7DUI29PV3dS+P/u4v
jrV5Mx+nQLd7vfeuzxjzo4sicVhcIOnAvDaQ0ZOfh2wFaSksuN0upWhQyk7/6OJZ
R7mY7WLCxngkKEEwICLU525bGfDxTtr5uQ/5tVhmyEv58QxKyvXECNhlurljNa/S
2/UHy4LzeTQmqLmqYdeXGjL3Ux59X0ewM1krhEuFoen39SApFdRGwsBEhdiAWhAR
54yqmIqLz/lEFwnoqpUoBF6G3QXDNxxZNQpnR4srUBrfo4oR6jlzBNUL++QVvVb9
nB4jEJDTK9UdhvDV+OWGzK+j0PCD2rrrIER32LhL3Mr0U/YHVIkCIy4OpeWIsHvI
ff/qJhcl1wNxA2CwWldRsHEOKwNDyG7sEDhnu07hVFeJgZsS77hl4qicizYQ+O7y
y5azd/zWxe2Fv9f/Vn8/XkljBXCugmDdpYkzQdW3wMcqumnvA0mS9lIKS8Xo6P7g
XOPHvepkmRe0jP+mcQw67/QfRi7Zs9+WxA3p3DcTP9RVLxzsAvqfXN6TqQZPqAm/
nOH7HtrCV6l+ZXYIBPbz5gFjHf6/LcemEXA0iBJFQwaMTzxjgjmaW9swzjSivpuL
fl4N6kGVYR+IyTb5cWMIvyIkWB9ig2j5fARuTEEHXvXO0fGdbMzzjmm85OJJhVYu
mLHOG6Kv8MMGdLI17wsD9DSgMdXjr5FXtmRHRpSrfPGE4eIW6olz5Pw3WY1PwFOm
dzvhecDEI1hrjPEkmzY6B38ym7MQqvlLhE7BcA2fPaFc+cMhfGbX+Iqr7g4kNmaV
W6T7gTaS1QVIe5alEZzVX2u2/ucjwhhp8+iKeVqeeTZKm++3PQzQ1gCgXj7Ajjjo
nFWXVigTMpd00Jcbtp2yEAhtD86864NMIkJJmQltJivffE6iS17cn5LtumYK5dxb
YXtT1YtIbQMPcuXLw+ADIbUymqosgDVYAOwZUEPfrEeivTd/76g+FxrULs4bVhvF
gFrv8XUKbOsXaIglD6Bt9iGWi5ekpYnZKgD0U7ksI2a9pQS6IE0IjbhLmQjATPfh
UwgxqcGRdNosZ6V0GmR0D79nrb1xJJGXR4TTkmpkhkqZRaQC9jyThRRG2j88B6qS
S2clKE9lbL+ASi0jx8ab4n2wCFUGM9KOa7sbWZgYKfkA2yFSzVepCKDU5O+J+Nec
2/4j9SeiFgSJgl4OYI1ON7ydlFXDnVk6SJE1B8+1SWCerJT2sG1d5+oKWNUH4pWT
QTO0jK1U0OAioG8KAZB0BXR/m3j/wMI9FnOtei90vMZY4daS3PyXs+MZbphAdHpA
DbqVR9Fy6gQmzQkQLd1NvnLatle4qltUciIfsBIudyxmMRhp2vEp0hbV0OOV1PFx
w3EPR56zgsq3TD+mgjPr79qMwot5u5kJGEyc06RO6nRafTH3b0b0RNBY/XQkda7o
WCSHIxrX3FDXaoejK4Tc+wrdD1P2mQIiLI0iSp1nInZv42FNk1TnpCChdUh7xSWt
3xqjx3QT+QKDjt1vx/HxHz7lR8lpLfgzi/peW/aZTZRYL+tPaQbCIQcH4vOp+Z6m
zJVlR/Ie1xsVEd7GH90MuLP9m27k03CicEUmh/px4jpGE8kcFZ5rVIrYyZcqFuOC
pFIaXXZ+eSsvfRpJXHDYealVmB1svDjtWyXtXzw4zzzTm20CPwp0O7pqkg8y8v2w
5LMbySV1Cv5AsXqGejyr8rBzdeoFHQynbhaxft8UNGE7idb0fwaLfvKoe/UpFunp
Nqif8mNu9uR1gydOVq7n2aKy0rNkcGrMNwVT5IiNGciPav4TAJdNWa1s8243jWgd
2Vqw34GJqXMKY/561tXcXUq1GV+YwCcMEMHCUmH/Oc7Eu0685dN7kHBZvaqFicY7
e9DtINReLry6qmZHAyGWOWfrJ+HlaeQV8Yux8Om5zh+AurMGTAkUd2gAUvT/BNUO
s0a1PYigeRmAvefzoo/HnkXy5SxZYbd7zPXJwj3NohpQssNbtGUVQtANrzit7v4V
mFJ7IZ2873PeaxIyaVh9Xx/XdzUw4aWokpF7Eev20lO3u7AdyYMhG3MrhscSYIv3
661h+BTflU9M3Fsfag8pcUwJx1XfncFnYMrYhFcDhq1O144LpbmBHAhTJ7Qx+9pf
iz4jn3PP0lR6zDOFiP/WoTleNcBOxKCe20GG/hzwltfSMftYfBGEn7+och4SpYq0
23ZW5U62mzTc+nCsMJLAahGfgZ2q5jdiILM3264Z0hPb5DaL/sTbSxkxbo2kpbp5
0+w5yIaugHKoCAlgdiwNnmBohsv8sjEkUuJMXWPsWmQ0UEctWPJ8w4B/kQvAnnad
eoydqC68JhMsFBohH2IQz8dXCjMBTeHOLYZGvXT1VEc=
`protect END_PROTECTED
