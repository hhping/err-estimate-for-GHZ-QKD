`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mh7Qk5kbBP3CYlSLvNyFWgK0KOvr5Gds8U4CcSrexIR/cjDxySWtFO3Jr1lS2RJh
ZcvkR2FQSlkWIAhdFTDYWKpgtTWumHBHQEGexyjRjB7b+qpvWwdz+6OhP6jxtDoC
ACMBzakMr8qr4EVrZ6ffIm+8EcJdwcpXVFY4OvsIW+9o6nx2ScAw0AwSkE7JNsef
CX69V8HPglZv2DmRNm850FkK/MTHfn4PSypVPG/Cb3V+c9rdeJBVX05Zb/JHEFOg
vnhfM3bSA3M2/q2P1Y6D0emQEaSNOlEXu5JMnt9dutBCIlURMhvWMCpcnfCLMIun
ZfLSw4+nZtPaI3AXJfZVnwiE7lp+nEVOm8zqypaoFs66RvqFOway0XiE1pM7pTn6
t/nP7G+rGB8Ni0HQThAwpJgRaNqtjsziWwx3T3aOrvUPGbBDfo+aftABT7bxLTs0
TBXuw3YApFwu94wc5ztRV+bqy0u/s0KLoFf/W9Z79De+7qIRn7SsJKXlFNGL5vy7
4TQa1A02R8QERw7ppZURWwUoetOX4ISh+pL13GlaaT17DG/+FxKIj+5VnTSy+mN7
zhA4zklgVCmhA1mvIYSaFYxwnBFR8IFkVmyATDB/ppiHKAiDbCemY9giHHM84a5+
yKIkM2RMDICqv4XbELdrX7zeX+sZlgQpfjRHCgTRsYkKcT1jQkQHLPQ3zTTbztpe
cfETdofi87hSh95a/Nug2gtAJNG/flsw8FCekz7Ocn5MsTxmj85NOKBiHRi3AYvM
1YNKtot/kKzloQhkDCG1pZ+UDCRqTr/mwTccnVNmdSkBfmI6hL5URSrMJmUTaQkY
/ixqbn1BscYe9HWjXZFr992jrNw2OJh0YyC4Rq+FL9JLqmbvTj8YFoVNhf8vnLCR
oYspfnu8dyHXGXbFK/qNg+BqCZ7M0774c8SbOcqbFc7KZd18OHx9jKUEAz5F5Ddm
jXJZe/fJobEGhCVGx3TOyED7kER6Vtd5Js/RWpfG5FXDX10A5v7jGNiorvpSBRzA
`protect END_PROTECTED
