`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JbFZglnxgq+LfhQ8h/4+A4wx1wnsXDgbeXmi9SeGo+63wTYhqlVDFKRdbn7r97y
vP8UgqKDSj2kA3vPL00tJAiVgNW+TGnruliPy9MNMT/jDTUF8WaMZ+C23toMVIi9
QnjQoe4qbJJ+TQrdfEvU+zI8NwysAbx3qUOVVaI3aGLV78Vw7AJVcbBOpJz9IYRL
Ngft6LAQTn9KRRMOhl0ZDxOUokO0xlYYWgr4JeB860h/YHXqA6Tgrj2htMEkwmFu
CGtWcbXhipTDVfc6ZRrQdLXetqCm86nxfmuWDGze344gJlGJ0NwU/7l/qqPdbkPJ
8L8+aNPqco0Kq/3L0hyYMoZJ3sY6wkOsbcVPkB/PLNcneAPRGe0xcjaUiM96GKHR
ggiDLKadS1vlPJQFqHLrVeaereGjCRKAcY7V4z4a6cvR9vepzpQUU+MRjo0GBf78
+0dvauEJXWZkjC8xYoUuM4dXsFhNL6i8kFeIgdM0qIwD0RrhGmWTWGOIIt3hvSbk
F7fZRj+PUu5kTRM8/uDsasZkPL10tyQpgkgzcKWigNDkwzJ5f5HRtPfkIrRJh4sP
z8giBHCWVtbUNiM4jk/Zt5TfzLdN9P+SX/gVoktEFLAJhSgXZtui44Jfi4a3QYCP
TWco+LpVkIsGbdkcQyl9qVxXIf60Bfe5xIVdtkJNZA0dcmyCXPespjoblZCKLz23
InMEsYGdqQNat1WWHfef4oary4lMwaqxSSG0jGV/MZU1wq4knehyUABlLciSXNya
TIZVayRA+Ck4m0xZT99VSHNnz4Lvko2jTy8duHc5UtKBeAFvwHpJfSIE6Sk0hqY9
vqTALyZ8RP0w4V+S/5EOHU/8xrDmEoU7V16+SSiBt8XuVPSrFK+nEJ3hKt+THEe1
MyvOXzcGw9GsxluLw1ph/g==
`protect END_PROTECTED
