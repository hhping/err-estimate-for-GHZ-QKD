`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jW3inPsnc42gYH91Dm11NHndIqVKNjXL/e+Gw+nU0qwrkwyrM5Xy5Gqy//2CDbn
4CpCjM6J3SlsReMnWHylbCF3koYr+ekt6RKxjF1FyA2V7z/pTqtNG+4y0mCPUVnp
NcgJ6cySy8ZtqdDsaZfPPyy5pvORKFhrKHZHg27pDEx0ErRbeFubF3h/kgY97SI2
mGs2mAKySPYWM+r7015Y/+EocUQOSMqNbUoEMEg++spWlwwRCinL6LCLfLbx6YQJ
AxpEvLa5dIMSfs/XR5yVkyJTBofVa38rTFHv5iUvf0JH4inedOzQq2+cpOopNd9Y
kMbchrlnPwhC/olxtfufWRVvtfEzb49/0u0PT3FU2sKHoUQxAgbrtxxGd8WE+ZVY
NVoGRC38VfvJcjOJyFtPzPmI7/QKnxT0UR8z7/HQs5vWfNwh5Ihxo03yweOQIUh2
RGx53jG1F2BlP7oEJ96hdpAAB6Y1bEQFWMwV5Aawy9uY6Uj6RWaQZpZoSO/q5Ck9
9jzaAY2Jow+RKahITmk6O6gki6JAsI6pd5YIxzHK1eSvxC7t80b1HU+v/SSYUSIz
862XT730JR7YTCROrLijpuUld4t3x6XQziXkMYglI/Nxvg0G7svS1y9ivYfUPzgM
lv+22bwKsmJIpvbOaFhpYFPyH2G7fdELtHziX1svXUIsTlUPRoiO62+LogyrpngD
8o287NXFpRY8fokggh9jX8rTVCjyyDAmp+bKQV3Bg4dmmBFkDXRZ+O+zgov5k6rF
E7EZcUEuha9mYSQeM8dVImW8+PcmonOkhcMjRyxSjVLa39hT6qhVkZ4MDwzZ78u8
ZurH7BZOwVBluzphjX6BEdvzaVPlsd1NmuVsfvo1hdyiWn4AhITYqpOjWndZ41Vc
FMltm7eadxBT4VAKLEFjA/pK07Fj8n1YtCejFwjlNtByJTrFUHyGK1pwhbBqzjY7
k3S8gwSQFgnI7qvPiR1bMBZpuyy4K5C/2yVfUO6EyeEG90bYWw94fHW06wO7N2jp
O7ahx2Dk1X7vtqLznwh6deWtnuvXdoiZqwRqK4ZI36o8tKZVG65tcPRcoQUisQsA
Qk/ex1MJfwPzNErphBPKkb7t/uYVKdbMesxxEyWYLDWXblovy8reAq/W50vsmh1r
yThjNI34ei4kmwvtmYhICxQ0kDIW15c/LO40w6SqaNY2YDQhs/HeS5qAZQTW71iU
LM3Vgfq4WC7U6xnfb0TDmWu27IUnXx8fQ/swm+U7Tzpa9MioZmH/ZTJK6Hdu2/Fz
86p3VCJBud6HNaE2blHHc1iK5YWBiP+EWgtDeofyAeg=
`protect END_PROTECTED
