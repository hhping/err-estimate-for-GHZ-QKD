`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OR5qvHV5cTNzhPDwGv0Addlo1bLdfshNO0odRlSjyv8ujdH2of26rXUwzrnrjvPW
fJGfYtbyhoWD46bNsR0Az0z5+dNF6uLTU9w0FzMM69dSK6m/HhfJKv8pSiZwI3Uo
UDmsSwSwipDU7iBqrxZUKMu6DkSNDiKlDijP0Dd1MyNNaWoLOtSlaz1SzyIMggOz
LW6OqY93AKiJCLiCBaMMyc7JcJu1ITmcCsTgdz/L7CnGefoPepRvZTrL/SMxwUe2
L8XHEGNxVE2aE0s3Sdh+u+F/rhwnU9Ix6+WuXb0a0fe/WqVKXa/Mry7KQSsnT208
WC7A4HN/lrjrcK3Qg8cvTBBhGYVDhAMjkF0S8mQ0akukf0VYiL/H1axEW3kzAHBX
COGm4fGUboj9dIIhN5mrA7s4Qxz3MD53nHjJYnD85LQyeW6zFz0tzejiEZ05gcV4
YnBbo3uYA3xFjYoo4tSZZP9TsycTsef807vuW4n91kOWOZp+dYNVaVe5oufzexqZ
rZfRpg0xeJNTglfJhqK0p2Debjx37CCIZ2EVlEg1RZx3ef7U4+BqwxcTH+KV3/tp
+w2HYV/c7bT0m+QJtibPTuZRVA/KpsgAAHrcj1FT5Q10kbyw1bf63fb6djayp1Av
aQ2VEiRZ8xca4dq9aNcFmRM58PoVNBKq13qk+4wr6XpbV6kvSo8xJuq2dWaCS8Ck
qhJc6DCu6XW1giPD1j5GCsWbXEXjrwZMfyfWIzRoE7/r5Og5asmP41MZR9fbWucB
69kwz2HhPx02pebr28speLnvbol/H272+0zplOE2dvIiSk7x27KS3JFerKaJPwEH
cGbpaON42cz4kmvWdsi+0a+bgcGRA7IL2n5YsWsSYmQoyx1LHoGZC0QvdhhbTFXO
xpBUO/N0RlGEnzN2tzFYD3IGJ2dySGkL/qg1eGuk4jBpbLSBPwCXxjdsBTswalDV
VWuXWStdEkpLYH1sljY1w8sHNsPxILNk3kb2Rs+QRXhfL3Hc3tID+UIzAT8NlqKX
MdG/JifpusNHeuQ1vnY8fMX91fGw4A72M2qFN1qCNgeJ41Px6LkBy37cuM8L6PGO
3MDr31DccffeqjkTBwkwjRDvWJq7HsjIRgSpHVUXrhhiuIKONdyu3IjBbsAMJUyh
Bpev4KkA6c6W++Mef2os4cGm+ZpWcI5sE/gbJJ4KsJt3KfRiFKSJDTBm03KXnwrg
l3ATkXFU15XaGz+rhcBRJR8DD6lhZEXaDkD+kaLxLy5pHT89ieQbuphxI/BWLBv7
MJvuw5hkCbBx+tyFnDdRrBnjVtNc4XV9Yr1w7ii0cbehufD2RuzwaIu1iEheXIJO
SyfT8/dUrjFx1UmA0y8XPwjZBiXWfMTPfvSa/7pbi3OcJnRxxT2y5vKtvHJVc9d0
f0FzjIGZNhbRdBr1mH49j21WtcmjjnXlOmJWY70u4FUx9x6DkNYOqJwXqPL7WIOv
NMax3DklVXo5ldORXcwnaNMgJ3cCaQeYjyAGufMv0fLmr7WXD/64aU2wzt6iy2uO
pQrHtM4lO+n5GhupF4C+vCOfzLhDbYhoSy7V8gE1nUjQ/rqjDqfnLEzjPmyGTZjy
wwT2Ru7D2dqi45aW1f4RFeKbEz2glIQ4bK/MKZ8eEP5mUBovJASTEn/zdFsmAh5M
DHYgh3recPg+UWLw3F0HI3BFclaiqssuiMlweWy5FQirhxGj2DhC6+h0/DRYGNVh
Eq9q+wdxxabagr+sgbWGSRY0+DRb98uyMjJmRhQZg5sn08QmBW/i5eGbpyiyLYZZ
i45+Mltl5mD4C8mGziOQ3aOz80uAUh8gXbMaFegOKDQJE0KnfnZNjR6t1BMN4JBL
/No6AfTpvyXmBT4ceyxwme6PbtaCoC+D4GjQouIYTEVRc3Z2OE5CZ0V46Txtmmep
`protect END_PROTECTED
