`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XGZXzFjmY7RvjYHDAViwyryD8KEg4M7vZMMtjL9x5tiwMsMeKKczJYQ0GsW+Ulf
XL6XH9ruhMTM45jMZiq64lc9er2+NyCSPATdHezNvHB/YNVIbEhVt3Fu7SL7ZeMb
I8HrYTEJelQoJarj2ETI9LDNU4OiPdOY/kqbWRPfdKRRFI4oP6N/PwnI50T7nX5J
QIALtROU6JcUG7Ue0zGuK8KmEYZA7PI4DiDd+E0GxxMcXCuYNukooxmhnqKWYxLU
TWfv4inxBrE5b5XVI3/zbWPO3eB3Q848QnSCiOHW0Yd0nFSAoVWs8M3hsR82EVjv
3VLsSMfLjLlgN10W09zySSU6g3gPyIUn36czdBJNGcuA0I87t6fq2U7Lcnqb7jSr
c7Coghso0oJ/N7OUrLPfJAnATzzSHanUOZ3mMRTsN6myNAl2Ndx0yxc3Risgy7fP
bqlirB8fLBHSqAuOBLZvvGO/0CWqqrfkJMXG0WAxIZRtwO+C4B/cXJgiJ8fs0G1N
GbFG7NdS9sW+x/2MmAsuSwi25LyK+TmfBtokDl3Hq2rYCi1snVJpOa1ggeHxl7i+
hCfLWsSMJ6g6yVmNmE5wcKfzg1OA/sFayzDCq/BaJz8sX0SmaYOXlihHnkgsUuVb
rq8Hp1uUP8m5c/tMKpKQALHtbKeSeKaAvVNBSeV9gcHbDco2kYoLnS5/ksOxmU5G
SsgvrF9x2+cmM8R4iqCHOqUgh9mLA7BxYAn5s1elkksLpAZMkTj8Iva/6E/VuLfl
kYOpY59nJInGFSVd/OGNF7tc5CzTDkvY8r08vslx6IJuSN8LPYFxdYDB4GZMgTko
BQ9gpk+cqY83Yu01DS0UqRBLG3tE01vKOyo+ntvadCYIwz4cHUkF7My5kXEX7adU
dQSzqtYgpN0xGjyHBqJcC2gN+yA6KgKyGMA84P/Wa7fMa88LNQeK8obIpjFiLgR+
B3rVcQeyAnPPqOqaSlddKR79aNurjUYi3aajY+/QtLsgsPjhv1oM4Boq/subckFW
NPc2JvhMiA3hNpnG1pkcXr2bOywyPDjhspk0XFUB2YJFXdUC6PtuC3DoKuvW1ZHY
qEUKycmwkscnMcuWQ/NftkBPwxrQ+xK0OGBQpXppVA810GSPj2atFwXN+XMKtrdY
AH4qJXNrjh/gtGE5jGos0BdlqeOnHmkf2jrR6zPlosP0vOR3Dadb8VtKC8AaeyS+
hTML61CfqSqIncOL0f6YGCTPlsKObq5mMqxgVNZuxfCy0BtYKiqiXaeuMNzq9iXD
FTyUzR32mF+OgNgw5hsxMAqv4NWmkf/q9OnBY5236NMIKAKAGU+ER4o0M8LxT9NV
g5FqsitzMc1210lXeGUssAkIGTLtK1K8G4IGVlsQjM4aTKFCmDWuV06TD/dYYf9n
vF4S27GT4TIok+5vDgo/sW7Et7w0Uk9QWQnE64UB862EJ/cflV7o+/pqUH5ofPto
vdeE3WyLsJpmrRnfj/7CeIHuXNx1/MqfADchEySWwUz/eluNZcXaJwXckj2z3300
OiOgzd5soqt3+ozxys5E5xAzmdToi/p1xSIDMYdzIIBNvd2Q2DNvaqtuMOdlHMoM
DguIYfa/7i+K3mBLQhWbGhq3kbMSNUJkFl2Zn5tTpuPfq2qhIZgWVuU9zGLV8r5X
MoT9NhUQDM3A9Ikb8a9Ss/M7ItRdtJNud/LNQ5Ayjvdp2AhpK6EF4OUH8vJOl/4R
MGKUoNxG1/PUSCiVN5XFj3FpvIYZ0atkW3eZEcffPtUaHOKhGxxX2G0u4oxp90m0
eDuR+p2+E4viK1d4cy1qyh5BWeWV2blfFQFd0Ri+rjwH+3P5QcxyPcNgIwnyNWm7
Y7bDQKqMCnU4N6v+En18K0ntKcLIABZCxRkeN4mFe0aqGoKTUXyG0FMcpbJ/mDwp
I4wEO0acBFm57TOZqiHvl4lIAJjlHpU2jx2mtynsiyK/JEzJRUeNvKFujaqoWc+M
gx3X46kCUvT4TrV8yzELddEKZ78b46eBrE1a207NvwVZQHVdJCD6r5Fb8lQ5DWLi
iKGxDwVYbZqSSE4KDFQqwA==
`protect END_PROTECTED
