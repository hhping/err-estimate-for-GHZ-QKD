`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bdT4A1tqCHyMNzpuxP/aMJOgLnJP/KBy61J8TtWXlTP66Gcr3jWFi22rC1I+yEU7
iB3Jxs2HNLNyKh38RDd36VVAiXLNxNVg8FRhkUs6GWhWTMmeSOh794LHfYqFK9+R
1mrjE+MBEQglXtKtlNQxCRoeZMRMl1n94r1+sOe9poCkf9zkDH+JAR5yxy3NbfqS
9/HKKRVjNJU2WdA+hPjZ7u0jW6qggN79H9jxQY02BNIc8cL67DiaAu3xiUTbyCQF
6dD0Z+q0ldpUo0VeiSf2aeSVB81lqFYc3iRKSS2YE667NfB8q+GVaxUju4T9qzjT
j60+KLKwhRz+jzTHQ0U+z8xPIVzZiRKPH8/3TM9KNei3muLS48noOmBt5loyrZZt
B18waj4XPTK3sEVaMdeKqJpGrSPoCTf/QpDQV+ctE+dVyrIR2jXvbfkYk8Vsvc3y
ErTSJDKQNvDc0kfgipWMizDIe9b6aEi6QiINLML/cInjBMFyyG9km/CV4wu64RdV
1jEYQOzvLUWzZYPRjjMfda5pMMx/k25AKFqo+gfoUoEXLRt81D3WX5qlPwRH66nz
PHUFRw3N2Bhp12+bWRGl8BbnbX8z0tuPKPx3sW/5PE33c/YdNia3ESp6Nm1QoZMu
nwFGWht43GtKK/CPgnefYTv9iz12IUNycP/Y6JU+kzeGCkJfRxo4gJ0Cs2rEMQk9
Pp0HpO2d4XfZ5Xx4PSiRcN9iRByABj4ln+A1WK48sJW1BJckmwsSxgWN1NRVNtx6
PPb5KS6DOP/RJs1k1ZcOrCenIhLIm873FZGaGzwazEEINnMWV3lK2D2mcK4B1A3I
MN65zuJp7AwT8246PNuMKYC352DSv/fIDqCriaWhDdP+A4janYwzkCVV13h3VhqO
ximkvOshZpPPbO3B1agyndjAF33g/PtnAAB+0RQmZBq9Vijt9KG20zMXXbCFoTsf
tDUvW6SDxQXEgpOOc/uuCK5TuIR74V0l+8R6TmtvIC2Nj56KewaFZbb2hFeDGald
OwcmeyvqMN7XtUVBGLHJgOewl+8NcPdL+q2B22wmaiLg3bZB20cIIcuuNiE4u0I4
Q9hdXqu0c0S7y+NbvQ4jk3Rd1CoSuF5SbiSgKScV183s8iYyGqB7Gn1sjYxmr3l9
spdK1EkLzTOlTdY56+TNJS3wX8SXPRDVVVQzrJsg6V7cl9ZqowiOEXcJ0ARl/buB
SPrnM+6xwY2wZIZr9sySdVQE7UOyK4dCu4aJ9Ed9PGo2KkUQ0zUTaR/bIhTrgiKv
gDN/airdKOdTDWsxxAmHM0uo1UadhH6wJ971eRikUG/UbHl91xqkTxBJ1RxkQFvf
GDZ8VLk7lmAdyZptSLyQU/hA0zjdvlonkXOjAegH0FB/UXWp026bKEEYrC1nzDhd
8lFcsjtxHbwlcmKQxbPjFoAUGEQA8YACRVVBgj9yQPMv1dulvHggIGipCkgcXRtO
9Ze3EPrYukjbMWuVDkfWUxtLOwv1EAJwdwetakI7utoV2MuMjjcv4zOQr+lJCLyC
fz4sAktENl/s1J739bVgGNcNhKJz7AUIQC59080jDKykXgO7Y2oxqv5QJBkf3ZDl
zu+HlOpAtpgbA1gVCxJnXSG7EFHMJe3GzMENVV5E3KBF6VOsPE9x3jANu48E2F64
Q/k7VGv4N4mlI6tRcIEmdTtLykpAzRKscRhTYEJZBJkfqqoNwQulVNJnyNQFWGow
/5Sw1FslsZsviV7MWfxxN97MZSP2WxggmDTNvVPTYTbLksH7WweA+ETS4Q2ADmjG
FzQ0x2nlOUnCnC9zDkvbXrY2BYm2tfDOoJLdY810mWYRLMuRCwTb6DAZPYTDiT3F
+16kcVzh5RO64sBbF0h4gVEDgvOZ10dnQFQIoZdtegDf5IObalERQeoABG8ocp/t
sBOvVC6BHE8QOZ50gYtgwGtSDweupfTVv3chjMQAK9knyzQGktGPoHuPCMH+R+hH
1P3BQUun8VWBXuSJZKhPLScn2/WijucncuZBJatRWuqA58t9ek33ZeR8b3hB4WhA
NeyiQKW589FGoaNcoVyDHEval9zVmPPYbWdO1PbFI5VwNjI/H3w5Wom80l9ToJqx
GnyghJ9R1IDeDxO6oP8h2tDbG5YoWLaa077XiVHwsLHpUP7YtcMitoez6hEVipmj
0o1gkvJzz4dWsQfLqWrOLEeoNeEkgsh+KaTKIKu1ShOddaOcucZHcQ+7YXi/ekHT
2A0/jfDT0d5xjUcHf97kyT4+itOVYBkRlHukIS4SLT9J66O2dGi9JWOptArN46f7
gHgoE/BG4N8I42lmxQFsb80JNI4fTWW3uCRXQuUqhfpKAn0ErRdiPGxfvjXQP17O
1RqA+M8qW1SY2tXcMSUO184/KkoqGKxeJkvuwwAVGzTkW8vmRSMJQgnz/veGOx3U
Ppqx8/DGGe+tsm6+BGNNtyqUb0oRZIeiCmOYzDZBRP1vCRfuiaAgCU46y8zq99jJ
8UUKmVANKG/EXQlSZKu3BCW00V5tGQEol9d9U4GHoHIkYQ50aOj9qp0CfrbsMGKs
+gY8YHJTNUJeduwoup29tKI7dN0kjEQa4p+4Qyr+6yZoTvVKf50oi77D3CO2BDJl
piwQiXk9cEg6NVmYV3An3HLnQk2DBd1iISIEuCiXmkIWgqcOrFBi7LIGwqxtZC+3
UXQxbsJ1vJdWFk8GcM6jIvZjeQ9qEbVUKOv30pNfCgmAcpTdsYHlz6w06+yROZSj
5jWexHi+Yi96UGkCQkWA4u1EaxDIgYmuN0eCnCi6hegIxqsmo2hC4BkYaFJFGkPE
HuOGOX8cWVONEqUAhJahYQ2AdspMmtQDQlE2t9W6xTULqs428gLZDQcSb/l6CLdg
VR3gN3A2MnJON0lsALZL0wFeHSAJGa3tp7esgbbpWL2ATlnDmEzTMkKLSSIJsRao
cODrPx8pAB5NIzEXbIq8FTLHZ5AdqDbI0FMntQPen6KKBnPclKSxQoe9WWjrCG0F
3Rnn1TtYQm4ULF4orIAVSEf6ECbu9ur+64nrL6b3kXbTzRapBlLLPrD8wbi9hOhp
+ffIdFEyQalVLj/ZZeJCq1y2Cc4zscJwuD53USdoiEVoeLxFGN1X/OF06QzzjWF6
UQQpjC1AZJprZn1esMlQDRPIn8OrY1QmFCt/hJf/fQrKd0hO+pUTa8oZeJAZbeH4
M69fChxXZQIMetLNfVvrZr6bXpvwKSo0Vg5scMkyGhBICowQU0WlDyx2jTB2gH6f
RiDOUh8zzEnnRvnvlUpSBHaf0lJ2ud7f9htsq7uChIGRgI2+unhZ4Ph/CWNwjh10
aKL1gsRXgjmUn0kt8tTugB2fFV7txlO/nP0UkIVqz3bJayuT6OxWVz+P7jDBwgXb
16upqDkeahovydJEgs8M03h8qrNtmh8IsFF3Y3pIhkYPoO/XlXsdxwcltfr3liXw
7e/M4LkFs7mt9eLxBDPkVEj3dDTw2b/h4FHkUTeX0dJcMdWJsyT7mQoE2uZk9hup
W/oyuPFa+kPU4rCaWsRXS/GxgXM/klfjDp5u1vvX4KglQMLjffxmndm+I2+o8RWj
MX3T/t7jS4By4QPMjNkuC9cHaOB9U88RzvyEdwE1tC3yAm2pbtQyjTMmr/sEQwex
lSl7b10OAolDRPD86lVHuaeiRwX3NJ7db2L5Hx4iOIGJEjtIPXRIuhCnLbw03PAk
sQS+g1S3dqvA0YTHSUYkb8kRqVxJRADyuP65Nrv0veh/d1lBZFUrWZnW2/dtV4NI
YQz19bDQGLwSClL5IovyXQJ7mxg6945iN483IqA0XkLyZYDUKh1r4U/W9SZp6A8Q
9nmCRfoPNdRHYA8l/XFWfO77yKQusWkmDnpbSu1LZrqnIUJGEhbuGjuAdUQ8lBxH
swpEMI4VzX59Eqk5v/+GE+Y+ffHSvXvYhZG7zgWYfr6D3wxj8BPKVR0bi4rhDBk9
CLfiyUhnAGmldFMfwDrluDJiIf2jpey7SNHiL61i6ee7vYBRhEfOdD4AkmpUiMOO
n2yurct2X0Q4E7+wiQd6lhyo0KTdJ2tkj7k10zc8+XcZaf3Gc6/NyzaAtbtCY0BB
8DHnK0tMuhr5+OwJyS7Mkab488U+6jeuFCSiVFmGIVa50k9yACwcWhOjPjsm7BZk
BiuOLWzdotLrt5zxIx2xuM3PV1THSqO+po2pTm/ohsilwKNFlLCS7nSEVQkpzbt/
dH6MPpTkhrVMJdBKJH8n+jkXq+vevLcZUmlFNoYrU75riDrL+jTa4WLRlqp6ctYZ
prrq0meY8Y754zSHjayiBeMVmRxzmsA5mj86bUFccy6kf/uPmCu3AykGzW7KpnTg
YU4TI6xcB/F1clnYQHUr+VH3FlQ/kxoc8GrrcxcTi5CBWU6jExSDz+N7gwgnYNkm
Ek3zVk+3FA64K/7y0ATuQwo2cDqtNoPmvVt4+WkvGdPwx3eAvlJhDXOpBjAf7nhB
XdFSR27+/+2TngoNNdvktH6Gs6j7YviBX3ddrHUeKy3QA8liOIxD6kpxnZblczJF
hS/wXrKgqn3Zy9Co5rzQaEfO7glh/RrtHEzHZI9A8oSvrAa906yJWFc6tFl/4TDk
8zLgIOdc1DTm6jygmKDvbz7qPkGAJpYV/ggIPeOIsLrwe/H/JnH2y1rPinC4vD/X
oc/olBkEsII91UAH4hymdwv03a/vlx0NUnHzxytANAhmiQCQu5ovgonqC5Hbc2ye
kaCqlETKuZKDrUIJxJNvnCbtBS6qBgn+THTJTsAm27pp0mg7Rc6+JnZsvSAFshgG
hZYDFJxUM+tcVQNx4sI2N1vNbTBRbY+Y64pD/0AifFJJU58gL9mE9sEEGM9S2C2n
goxHBH1B6c/lYZG1HtHw1oyApDkWf/xwAAT57R8tPnB/UumAV6FjZ+jDf5N/gmZa
w4leIRvAL7+3xabw+qd96UiLCLZ+V8uelRQ5qBZhGayzVmaDbWuJHJp/gsc0sxm9
m9ocHivzkBuy+y0udPV/no/FQoCAoGksdHvY/ykwSZ/SoYDwdJtuhRj85tv9kuks
YdaTeaTYzeEyzEb+VjzNAeK92Lm5W4pfiM+m4hsUgpRL6YOdHdFrccc0V53KwBN3
gwC33B1YFigoZqyYd+a+zvBAC50Pj2VApWcf7OGDAK3uEeczsBhzvvWST0WvBpln
nHDAlDbSZ2Ct2/4qM7TM7t3Au6ef5D8XkK9mWhRCfh67Bj6ZoEixIJg+pDj8BFbm
DUjo0r51/AoFN5A6ZT498GDuTTwpaIv3W+N6TfrjOENzeRslNxfkt1B13+qb1U3z
a15j6+6nB1/1br3LAeKRexMKD9qJ9Nc/vKwb158mo6QpIi/TRgHr8Gak7I6hFRmR
yalQz2V3BPkDFJU836DDV6cgELx+XKNge1uFgDxFo9mbmpHBYAlLiSa2HneQ3w1V
U+30OXRCexFk0HkvAGLDWI0afZmnJC2UVw/CcO71+GaEPte44/6NUp40B6rrrQpg
KP1JZyya63mdT0LgRwFEVvJDCMpN1Pklm9EIbybuANRmSADhfXo/Oxd2W9+aodbo
11DCfqgL4CWVtMeQQLhHwdxTGOBgYqwLLdlyH7+qMcA5LURv+m/XXQG/l52zuFp9
P/znE4Phrqwr7DgBUOtC23G8cMcNOQlHaFQsf1SEBp54BZaSo1JczN0GNyl5d0xC
5+KXNn0lrQEvozbQ3M0Mwz2UiFf7e0vS6oj3aNodC2K1/rWy4xcqjfQx7RUxRU2A
mwpdSBopcjFRggA2lDwGXHiKgDzY+yAeWYdtS1fdv5ad1X4CCOmrk8r4iETkW8nH
wN+SIrKQBRIcQNLn7EgfraLqRs2bne9vh0DcLxW3FbQQpyI9DjQFiLM78VWtXn2r
cZ9iLbBHt9K1/Rodau4QDTQs3PqWLg4FYuEt3H0cEiO/FSFoli6okrQyJ6ql+Llm
RBBBI+MEOTEjpAiE7EPyb8Ktc1GrtYHUJvTGK/Vdf1CneyxjkU08jtrmcnyDxgyu
xtoy2/f7eVH9We61vIsuxfujButNfSl4IQrtyvQHbbcJZgVY+hCH1v0+s3/3T0pz
2LLtdYEwVW4990Rf7/vBfrQMSgoaSKee37Pv3a05NhpFbRZzaGWJIjovpbqQ0vTu
DyGji2vkG4XqkbV43kFykMzzOWSYU66B3T4aSdDJm1HGDyPyN8iPENDET6LD77FK
eVyeb21ZliiEQNWEXkYfdFesddhZxawb/0Q1YX0zoesv/UJGkkheA7FuFZh1n2C1
O0kancTg8kOMrW+CdcvGY2HfxPESHWsSyb9R4eTMYBmeklL8pdmChK/tYX18OtnQ
L10H02C9V2J210TcKCPpT3m/nGwCyOgcYg5DFxF4BEPRhBL7QnNPgLL/hBDZiJ56
RX0IAlal/nUPf8AacLOGDhQPopfjxAGlxBg+THZFSs77w8KuDbPtidmSSnjOe8+m
kg8a2Qqlw9O49ZtKi7jR1+7jqnbS2mrjCjo+stwUQuQcAhthNB4BtlFo9hJ3YdDX
b+iaonbqStWO77DjM/yNOpuRd+2/txkd6tpFiV4NFqPjfGoyTtPg9yi0+V9mcatF
Lpzl3J/QoJ9/0JtBiH+hhLWOE/E0DQVdKdYNXFKPUZfi2IU8yV+zfRrMDaSCk2WR
b+KUgEpWQQyTZzbt/YR7/x6ND6Z+xAWNVnirxNnFuhkk3022KZ/IEApJEipZiwMN
QNqvTOtpt9F8o5mcdq18qXm9q7KMbbxd71wULkZlJxXQDLjVBIIffG6lYwAadLZz
1M/CV+FSFYHdpwzxvsK7J3nZtvAwiKnqkBSNsgPahfaHpCeujlPFYHb8LyuprpT/
Abx+Z59if/ih7iPjYcmRmaQIjo3nXNimAtm/eDy/BAB5xDtId3eKoKWq7oY+2Pff
xecIE/SOA8c2t5Hk1H9rTcTtRq2HCf2guWfVO3MWyiY1qGExH8y+WShXxMWcS1zN
2krBovcjy0Hd6Ri6NwN+FaCPlTjR3uXr2rohWS3h1KcAilBJMcmuGuaANukdCaEp
HNnZnw1V4J6mCNTtGvySu5cT6KxYzt7v6AFSJujBexy1c7ZVJy0ietcEIkuXAY3W
SWUibeC0r7tA4gnOF9zzMHirKGxEHZ613eSs6CflrZhjV4LXL9jOXoilbUO0NZR9
tNdrdVZ+7VYJUTEMj1NKN10FjNybiMeLsJUut/O4hDfdcD+4xeMt140EEGijpkHP
/XS99kmmC0zrW4hr4EW5oh7Cg1Exlb39ayNl2g/uBW0PDWVCkpOUnzuNfa/sfmHF
9miUVRg9IioVXKp1kcUcYvhXc+9To/zqYbRTVVO0znzpF1hUbPMZtdzbs1nhz4u5
XAFSI7eYtlW6UGygfCryBXUxNsaQMFNXFfeL/LumWJNKsAL5E7ob7DqNElND/ktH
JUGJOs12k79VuY4qPCFK6rwV+p3dmU58yjO9/2vRI7XXcumMnGknH/8NKZ80ikpr
fMPGzfyTe4hO7P31YoMiJb/zfa6AFgqRlBc3l96NNDrNC9Dq6t8LE5vVehmBjDl6
XmZhW55K6lBjUxerPqYWoFz+1SheekaJQkzYuHw+QIF/IFyfNS962ETuj9bWCsPu
No++rD5Isj6i8xkORC8UxccG+u5nvmTiNjKukdONzes3ak0HhO0RqlsiSqxTZ0Wy
BobqmjOptu91kjWAUSlPJWdKXSm2OHKgfdQyJPgOyDdzVdxGDTIM1RKoN+MEuRwj
3YFxJ4AuLa3FOPJhbQVOju3c6U7uUsWAroREq7e5+9qjvigPsJQ04B+o4vAODNBS
+iQulART6wjRkhbg1y2y029Ca9PnH8ukhR+lz2V4dq3bn1HxKGsQrsT66vR4vn+j
DNDZXhRb7vsQlGzKvXc+/UhMeLcm7MqrXnz283SCliQOCgmQ/dQvya97gOuZDAf9
7BHD8CDR0XwMb3D/Plj722xEH1lI4Pd2IPvK4wPk8SLfOBUuIu9vGoHO7IP5YHiU
y5WoxdlUfhEzIVTcAjz+fbxGNSq9XTOo6WAmWrkKJ2iLpv0mRusps7G7BzPHRdW7
3WBaOLjtrepOLqVjRMho/8gzoGbuxRvRGwn06WvwPPot5Ryx5pznmjB6ujh05QAv
eEnh/fqE+qe/gAWdAC0s7WeWWLyjg148psXPE6qE12GKZlBwZ56RE8rgs4hmXfqj
4EDnOl0xqaUQ1xBkB5m+7kTmdoH+2WQTEXy6Bqnev3EIhFFNcuShJUeXeFC8oR2/
3gpH5gCn8oXc04EztPtXXQK2EdWanOykTvBueCs9dvr+z/y/WxK4xt9Cs0GwwnbY
YxBEVe+ID3q6bc5BEk8yS+plZdrL2ZxXWe9le9+X7yhbNaoAByMKc5GmXWN4U70f
FkixI79K7UoHzS/E8TjHFKGd4QSj5YWAZuRcY40l8KfKHFnY9bkWB2GqCBSPKUGH
CmEwoGhb00JByLx8vX3Q2rj8FDUUlUrEaQWwL96bXxddAXZMadNCgtdnUak0xYmt
OVL8ltGw9gyVo20+BhCiQ4NFLWAgaGLRojX2fSNITk063Xhg+G+8LnzaaF8GLOe8
Hz1IaoJcAt1Lhanm1ob6eoxXzGdyTYzTAAb/UZDbFhJFzXu9Q+pXIK4aVwG7Yvrr
AIJfRsorRap2sFhdLX+a6K2Dd3UKMW2qNfjnEWz+zSsvFbIwzXMRPCNJdJwjK6ci
e8bFCV+fcHEakEsYDMA5cZLnkMvRaDnyULEXt1uwNUrl5D1/CP6rC2wylwK8r3qh
rdSznguVgSx+AvQCs4sLS9TTgNh8mhVFL7ylcobhqygXaRWu7K+WBIz87Afv/pu6
ZQz0UiJAyLjHuzHG9jbI/Z+3q0BR/F+scwrJRTPeD1ExE32EbqkY+lls8RCkU1cq
MV6dTHpqqDTxNj4rnU1xcJP4FVF9ZmZHI9hH/zzfQhqLta6aQj/U8bxZ1YtT6dgC
yac6ZShfqemghJbUtWhsjaiStF9X1LlEUAV8NwBQMZ5t8rOeJBwFDu9nKcpHL1X8
EgTHuVuM8FqWUSM3cOpDduaSJyuD04PnTArabWiroclQ99VHuK2s5ckgZFtKGd5v
08iJ5NmZ2EsO4Wpu3QDItSsUjlIwjU/YTdEzYAfagGWMEFeQikq+gW69kKUcwMMs
UFbvdIj7e0lmKgNv96ByxYWYe900evagZ++foOqzynz6a3d8kEe30yVDN076gqoj
Cg+yMkc/+4oyrLpUSRHA5jkw2v0HQi5ykXg/LMK3NTkA1xyqG6J20jAN/VaHI7Vn
ObajeQwZ4zXddDoIe+psKljr71glo1LPFAfHKgFr6qrrezl1TPAt6S7skRDO/0/H
WatqTPzowaKiGC356gltBKEETJNcMYpqgGsqwzVn9Ax0cFpm2KP7ac6wc1sI6IP5
LFZLbD/531lu4FsVekzsfMRXvgm6hAVnoQEP8xrwx2tJmsp/1E1Dl/y/mEisUOXB
Z4+vHyj3wnQpMfmxOpkxbpuTg3PJGrsNLQpj8V5Wya1gQk+iDJ34Ets5bPZqqACW
hlaCZ8IDcL+Gjj1yc/xHqVcsJw1yXtrqDP5QkWZCsIHL8FQTH5M5/cBoZNhDCDSI
E0k7L0WkxvAypUuhjY0x6iGwj3HpWwzeMRJCoxydz08IIErlYVKwpNbqyZYD/sdf
rRflXPKoZYaE56ykcPrq/ghg3HBlRaO6DI1IHMVT6S3RK0ueeF5k1MQyJ8oi4E0Z
/vtcSpfkzYbkuNm+36glDftwxVaPHs1ysDpTb7pIFy6HywcV/XwYokcjZoBBgmsW
SwV2sRAUzEJnuW7OqveZM2ioF9JbSKTmTAzBJtAi3Ax3BgMZ15xUvqM0zLI44n+G
sS7hc6nxQ1bTYxsMegBXctWNEiUo+Kf+Y9hkTyKJuG4ahiiFN7WOXPi84Yahs2NM
Uyhsr0bM3+Y5sPMTZdWAYGTVbHYcbxCEBlih6q6tBKPvnfNxeZPYsemKSjmujDsx
yrGVO/6buXXjoz9/JSsDgxMDaa5j7dG13z/i+/0tRy0EdzuvbsA7YKO45LTSTAPD
sVuvEeNDJOvAhi3Hfkviw/FH9IJZYxhPex9Z+k8kk6cux7dJnFM+SzeTCMtdBIPP
IDl1+dk0eMsbhPRvWPFfA04+jUPzsL8OubXn8vM47idH8GZyBxSwFLnEh6CDW1gm
iGdrTkZD2GT5MzdlUMmK4OC9o3jgn0XtUZeIzG8MefE3gTnfQXcbSt1H+3rF4UfR
5/MLls3U3oDXjlorBAhg7qtydntjo3UFdd86L6IjFtq1yVTpfetBxwIhgDtMrSpl
O9VICpx7y/sAXDmjKyUHQf0cRpuTO12fix7amJmHkoGRAoIUH2oyq1QTH0Lu0s1V
UqHUyGAVWAfbglXGav18hWlLBpSJQvJWSofed3n/R50WzlHAhalLAvfNXW5RYGft
0JX5IwBrNlPIFT6UFc7YAODR3tsmpoUkSZvS26qDmRmGuYwpQr4aRnu6YxX/1nhd
iPKVORSoERBBEb3N6o0BzTCjIRwijYMC6q1Nrh9qEZRINLWCpJzYf0v9hGV3zwC8
9t5VjSRiePzkbOYBw/IbmgckzyI5Gv0D37T+ioDCB7CwQ2q9TmU6cMYJt3rwhBQe
KyAkja9ECSy2wYO5iiun15/jbh88L9a8b1Yhd/d3Jf+BXOD7AlOWLNEIQnrM4N8L
2dUDseZBUq2bRW8hBG+Ng7FrrFDCqnmicIb9K5nn2Rkg4SUL6910QgVaRDUtELfk
rmhAUTbk5z3yoroFISuy8Ek6sK6+Z3MU7zw3zmk7Nzbv8Yo6wze2OTAH84F40anp
qsWZsao2hctj9Tlg5zUF3ETml0bRjSzPboOqQotC/elDkyj/Pewhoq10FZbbwBZ8
IrTpSpNBnQ3yQs6SR8dKLcj9Kc+FMKZrctQJjQ9B+kEw8897ovmifrF/zqkfecyt
g9Ds/tzdAH0TVve/zYhMVt0Ns8TEIOytHJyXacsu6oFbjLLrZGnsZl8DQsAwCxpo
bu3o13DcNY2MAtbGCTXjHE0eCzNSBVT6GfVswu/i1tTOpuMrUSCF2nexc+f2Zv7I
OiCzL+utxKDslvNgInSX6giVifSiR1cU8ixVHk2FltaMYxyJbLzLU/oXWoZW9RKm
LPNKkiahwjJoCLGZkseUvLM8T6t37Cqe/VSJEiD1D6srww7LhiRsfWJ1jc8l8SxB
jFLLdXBk+1nCH+eGnp+HkHGPM+PO9a0AMP2lxB0hOgAKiogscsOqxMLKVLBgPRRk
mZrUWmpid3czQhYOwGgMn7/QCjPnHuRq72uEDHjDbuW+wklLa9tQxNuyXUMip5nT
ccCVf7aJ2rRhMd0FHB+An2xZpwj1y7TvCA9hLX9go+Wp91CkZoI6TS3fl2UlVuT4
txshYurPmUEasI3QQ1z4p8KU5C/Npq5lXIZxQIh2vXVXH3jDLUXNMkTMEzF6Xc7Y
selOq1rXujsecSL35uK89B9lZnjDoE+crG3ut41YYvmTfW/x32S1jbmR9dgYuOyO
JFt3VYIKA87wmry+9Hv2EWpx8saPcOJ/jciXaHZs/LOWsgdo8eNg/VdS5YKjafTm
qquhZ5mr/wuq/VjQzq9xcl3KRqzbSKUIzZK1fRz5ubKoS6B5CAwQOe6g1/xuw+GP
ayECqz6S2IVnEFmCLL/ehJRRBvp0p464XqJ115DcSet103ADxCi9OiqaUP70xWV0
eCCC/B3lWXU0OGbZ6vMg1z+maasu2rk1/nYtr6gF7t+/cG4Hs7cfsfgiXB+Jnwg8
X1iXCfusYWSHPVDE8JiZmurO4BXAphfuEv9571wSyx+TMWiD4fbWtuCHRgGpFNRa
qm0zpJuXUiUBXKhQDtXYYHFM1tRzSolUBYFsIK2gnWGG0TP4h6K9YOOb5rNR0Rbw
6z9lMIjFyXc62QhrPqFECsCzazuKCH0ncvL1UWyNiRI2Y2lhACC2ReQ40vVpk1xH
alkujZQ460KIaq8oNPJ2VxGKpTe/ceT04uAZ730ABOlRCDr/ZpHU7WjTo2ooADst
ZhSrAXoz/tXMJOeeOgkmXiAuuXZyYIpk5Wh9Bd8KHsm/uu0KChvMSousQVeYhXaW
YzAd3cLH4YVz/pS+hjaBAJBrGAcbUVA9yUOjGFVgOp1k3EFuTgAhplYTUdmrwdft
i+N9k1Ynx2J+dn76v6cwa8Xcq/xZUI2+WWxVJxSWkiivr+q8SWU2VoKzb/XNk5uE
kkjfILGcznGiSKM6yZo7IYO5ZFIr0LgCTNlBA93k9tLG/Gj0mB6nlptD3pnXqyj9
KP88f9GYEvN+zKTXz62djQooUv3qMIkRNV/utBy6g8y4EM75pOcLq4RnzBaYZoZ2
lm/VDzJUrR73EptX/D4QEQtDpmCDrdGQ0OzSflwo/DNZIicArmjagpgD23yZVwrK
eKpAuny6XNnidQ4NTSkYHgeZRwvRVELcbM8TJUlrW3zhqsoql0MvOtb1bJsOevxU
mMCkx/5KbmXDR0CJe6LduajNFGH0WmB14w93XRzsHOF6BotfsGVk8ZON6MjwtoyU
r60+yW2zUq/d+QctiXEHwJDXwHn1HoN1unQC8U/+cPgTiz0lHdDbqSyijnP4QueR
8bDv7JKyUWVtGaQscMUtAkn/bzS5id/8s91Ngwdcz/FlGnmbfUwID2/AGKtdcRLW
fIuppqsrtftGYqgzbBm3Z9S7obXttgU74VY5mMxKsoVAF/UhJTo72QjL+IV7dc2P
OCc/YQ1VwSb6KfUwqA0xW36p40oGaaSV8KfsTBpJc0EwPfx/ZoexOwdBQNmBP/Df
zTLHIXUxNcfNqa1f0/+2VQbKsY9sxs02dBg6dnqvb58mjlvFBTx8LKLRrMioNZRY
9Uc4ed6tqQP4gGaf406c8kNeHTeFXEYlNAwabFEz6z6F3WXPovI9+h4k0ym/mhle
5N+YsheFsTXv1noBmYX4qTU5ceKjXmQVcb6RgmxNc3+VarsPXKy16pMdnSWfwRqK
9S46oq97sCguvxj6skOWJoo+CgeFm2wVGpiAVK367ddx011q5g5UwTY8QP2oAatl
WbIGdfl64hZymWlW+KRqgfJ4vczjmUZBnGtyWbvXSBYJJZS7lTvMRc3LhDpr+EJ+
AgooRqCwcuvq5NBCKVuKSnxdbwFArnXVoy97U+q3zHnLrG/bYBRo3eaTi9F7xcV/
ku8OpUXvo9rG5aQAvaDn1EqHV6838axeX4xNUe8ZLTKHijNEqOBL/duSnM1t/mGA
zHSNd13Ywcg8FMsflHAbD5YE369ycNPFZL2whdNBwqHC1A/NWwxAlb8XmMdf1KX4
PN4JuLsbzhhwzRKnr/RRDiWxQddoHAc8MckXGZlUGwTQJBn1YOh/pIOP7NZk7QfA
RLh32ChdOfCnJcPT75el0hW8BXZZe2/RgKoG/CP8nVixVqypjE258kkYAVw6nduS
T/UerZfTaJDg1TbTt/PIMcPWSX2iO8O9JRHMlTfpTqg3n4++lolHx0TtjoD8FfoW
BQ59/GijEFS7CfwnlcmvJvXct/CnGrvcrKJeNoYhFLIFXT2lJ+RugaJuNYd65SZt
qlreQKVh0lr4OKKZpoy0PoZWHqjk4mUEBqc0C+EdJa40SBoKX+z/MMp8gQJwsxzT
GI25pPsOFbNDP1+DdR7pQnq6Ab/0sCx6d5vv+RPU/1hoEInpZJ0qf5djSDMI7r+V
LZ19LME+QHQdCKdgtzbr3ncBonpy8916ceyQVj+IkNsy0CEOWb2wxb96tqUYBO/b
J/b1OX8iBcx+9GOqR79Fe1td3H8Ly4ORDVi3lZrU75fyGWLy54jct0hcHt2yZmpo
iYxeidr1bEEG2np64pprNybgcp60KPix9eo+f1AzEvd1aYessu3ZwNnEErdn4reI
nqqz0R8KHKIMhP/qNRuiopiIi9Tzq0RWfg9YbNCtqE7edQ7Xp0z3OwwUg5hu0bcg
niOkCMoi9RCL/xpuXHN7CjQi2oHw7KP10TIMD4Z2k4rKNs89ztIVrVxxvE1QqJw/
e6ianBSspitNtwKTc6+dwq7q8ZVdrzxxca6UlzSqkbM=
`protect END_PROTECTED
