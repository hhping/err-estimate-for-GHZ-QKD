`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7y5FKrHz6PNRf3LrKE2X3YLH54e2uxlmcogdaMOTkBIF1yMA5Oqk/KpcOSowfRFJ
Sqr2gisOTGqnC4+iGZZOo/SMWSLsOYLOYA0YaKl4rUYjfSl8X6YAjanYemhD2syX
xamuPB9f4SSPqrcpUIAV9g8I5aP/PM9oHDTCcHv+gj0KSG0L0DRdsZ1Pam3wJm7h
5uLqQXG+bhtouXSzuj9NJmH2RKjtEJlgXIWA2gf4Z8U5wElEHbH8ptVRiPLSoiQy
TG3mOadr1nTf8KiyLsNbXgmEtO28J/akthxrZlVRcBD3alcfB88+pV082GhWN0ua
43ms7G1JW5RmpoL6MhaaZeqeiwmCCfv0/UO+lwC/g+ISKvgZ9Imhi0gTgWVy5czj
wYAozlGFkYY9mBrAL70RWxau2HoXDgbhPVCbErGjQRfjgpynaLam8C1pqrJfg/TD
oXMOT7FOQOM3pXkFtGfM31d5WqPYXa3BYmmbclMcr1hkSgyYp5Y9NnMvz5RzFN8C
ex8B07Xz9hOeQk3Cwr0CLG5R2fE+nI5OUrW9j1AVJXGAC6Uh1EgDuG/EwA4lILx+
bP1+5tSMfaDf1JOvtCG27KtXNiTbDXCD+WfcZsAoVeC3iRMHTvQ7jDIfbpYyp71R
l6vQGJrFMjGnNcK5oB2mSQlpzWuP99WGDG5JLJpqp00GrMk8oq/jIjZ9R34nS/gH
nXdCkhjeeuWhDWS3cScjFkhAsF6CmxAh8Af2eQwVKbD3GaLt1MwENJ1i0jiHt+FU
zRQehU3fxoFXfLROq4diibBXJY9jXU7amNaHMwfC4UAMBSiE3qyR8RUmWeHBxbvq
uQv5oLJsBvteoMRW5pYennVdnwlNTHcNkp7axjaQz8YhHuv5cLIUFb+b/8uwcoz4
msNwaXMohxYB74C1adM2rY9Rrw6ngnkfa4lQSU9hPAWRreK6JIx105V4kqqcqpcx
CUzqXeCq5ZTESYXScLQbEGYaUZjPmBORpN+amN05C0vxV9rgyaqyQM00nr/wBRcp
zdEZjVvDzgtNCDX6I7OhEtmL/Xo4QhjX+YzqD+I7Cx+lpw+nRV4PyQd6hUYrBYrd
bVpki/AlhCCC6r5+yzlWwNI8OK6gF0xq6C6qwBoyQPvr5FFwTI1H5prDEXCT6cal
RIn7NL9qD7cciVrlPo23Ih0Krrs0xse0OkQXhd4R4qh4x79UJse0tayMwlKrGAYu
hYfQIzk5WUx0DahOyY1DEklYdt1XItgpXkdYiR8r59sbFpZ2BGOc75E/4hB/+PEI
wrYC6mJpLDXaSBJZSdSBwq6/vCrpJxkVa91qNKXNmMaYSkadz0NBsVOL1kREMmFS
2D6xELanxlLoOvNyTpWehpUV1s3rd/JCp4JaP3GYcW1L3jTI/YDvzhuvSUIY1Hfe
yOsIPMB/X8Fqnlg8MRNqO8l7hUdO0/5JqTH97yTm1uJdd4ri/eN3YxX2K4u7aXTm
D+C6ByrnTPi0xfoQP+rdZ1ImxzEwlWzv0Uoy7r0KsjqfeUhMgulbu+igxEcgtMrl
BBMpQ0xZBLFQUZLOED2qSB9OTuiJTkdhnnuAkGYecYUk2VbVOL91iXNTZmsJdlh3
/Kb2raCTwd7t7DIaykSQoBh5oQm8zwiN0T/Ccz5mqpVAPLcAp8W+C1D1BMe8TzOF
lER6L/Cun5ELti2xMlnZIWk4r8xR+gycf0nzCU6WshLw4m8hTJ0EmnyoGeFVnzAm
l/bJ+NJXVDwsBPgT1eR/ungVz28TSHg7LcIIZbDeWxbgdHfshWX5y06KjZ9/xGPA
gFZXhbdkDm6KSG+zufOy+LPiEMBsHhI+VNxKLAvdM+5DnaKOZ33g/ko1rOT8V8uC
0u0Xdaws7J8Tyl4huelQuHhmZFbmOne6w7THBgaRCQhXmNNK/llBjhjkyqQqTaJI
UAvZ2ftTv1dnJq1rYVDVWgba8IeoX3ef+lGaYCugNyWKqFWpG3joZ2En6yPFBPlR
+xuj4HZtPut3BdYP3qBdO0axa7iW+AyjLVdpZUlIwy9jPXUSoKHoCWbCW1od8Ket
liakZ7zy7Ktp/VU5L1EGDGPVEZ5V+cDUon+Nv06NcWpZ7AA/uBajkZWoDCZ0uuiP
Xz4sG4cXSfuWH1mZC3YSuv02fgaz8NJCJRfxuctpKUsx1mp1mqHmJy3u/yR+7to/
cLKfeMXVAejT+TxgOBN4NVD5w28eZ6/SVwOCtErWwB8VkClLdRWst3B/Bdx/Ll7u
W6aGcTz7OI8iczGs2p+3bN5VKgAt4CHaHE+aGOoM659+FvDK9NQR8UllkPWWVscM
Q1l7DkA7YyvfOPvuPl6u19xkXR6WmRsUFtaNCwvqjAgQFTAx3y/PohpgeLr66A5q
a1UF1UO74ZLPOGZVdAjj7evIeM91eq0QmXdpeIiC0DbwB4OyW99vAzaBsatl88eX
avCBoAoK4ueGfNwNzcuA1nWo1WrwFMhVDngo8F3MmPiLvwXGIgRT0yLv2btYQdG7
`protect END_PROTECTED
