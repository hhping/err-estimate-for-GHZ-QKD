`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bF2dHLKZ37FYXjG+H0wzzCOJtv6VK/RDO4T3UiOnM3cLZfFdS6wOyPRBK7Fg8kSW
FddbkWXSdXK3qtIQi0vSKGJbt/Y01rth42ojckyAmr/hdhM9VvhjvxJ99+USy2NV
Kj8BE/emC3aRIK+K5ZAVeeB83YiFIdKhj64woYu8C+MNKCy5zbODvmVjpacS05ug
6mPjCg+gPi+qFn9+0UWa2TycTyn4wgSa4jmgUN7uoYJvxuey8zMDZwVFEtseuT7P
mnZnsf2hKJ84IZg/zy/8yB9XOw43p8fYO9kqNpOzoFtbDOKYhmwhi+oCvlTgb0ad
ScxI8EUglX+m7pJUzeCbUiXu6TsrACD8mh9VvnSgjizHmIHNHnUEmuIFFDRrNPjd
NvsalHa3bZi6zzuNPCWommnT4Uc0TI5NSlrtaOZfP4TC2ZPqFfMLsBOUyJ5VqXZL
qovEh6rBPNVmaXPNdk6bwPg9Ic1fQOpKjHo9J+2CFwt2PExsyFxtPPM1ZIJyjSSu
PvS9pVGZhfT1S2LckyF7V1ECzTVKnvxy+6lC0moy0tPnAzGYbsJOJVl3fJ956jka
ovY8wWbuBLMlyyTTYfxWGizPGI9mWVHHdmrLn99qP2dzTvT0rjf+T0rVILzJq8dE
8Ndi2XjfNQXnjxD9EbQWadBVjtaXqCVB4hybcSwUpatXHzit93Netm97uxxpg5dV
TiAqhd94lFXPZnOjgR8h5R/VJuLMScnsN0j1iF2fpBZcWajYIqoLbmfqUMRyKiUJ
17nRwtlqHGE+3ZIl8fxYptWoUOB6rI0aaRr9+NT7VDV8oOdqq/LsPj22xRI6hXRU
`protect END_PROTECTED
