`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
si37NC8y6Y0tFIbgync7EmmI7ZIMr+UmM5iLq2//3JwiY4QlHu31NBwOekTjOX2J
fY+ukrnja+rEfJqfmut9hW4sSu/i90G/OpJG6PIz914jG118vMP+NSxq6Quc7Dj1
tjhELSHrYyfRL76BKyHJIQphZ/CU3D+uJzXSIV4zal1N9YEYkTu3t+5oo3ADnmeX
Z3AQFknBdmS21Q1gJToNk2kxWWPSz4SURAoMehHWno8kmoyf2ScweksFV/Z9N6+C
hK+RH89xXE99TD73G+GcwqMWqqzfKfwmKNji0UDXM69I7kdeu7hWWqUdggKPICw6
oNI22h1NlzLx6OXkdNVd+S6DeJkS8Ki9i0hJPy5DMLQGPUbAUCIodrvxkYDSd6eG
6cJQ6efLsazzgYz92MmSGGGzNPq9ADX1O6I63ggp82MWTgnXQsp+K81XtwP6zwoK
v5eHPKbDSWCSsiZEagj9dAlIWUyurevCFWUqVnX0icq1eecsGsg2pdkyQVcpzdcJ
SCz6jVV0wsiUnn7RM5yDFBlFNtJmIHT4uSLbeWsOO5QRPb4MFRd5bO4sUhBNh0AE
ZLU4L6Yl1KLISxLAb0XnsfpUuXakCoAUX9dFeSatDkzziRkNv+tdbE7bkAzEJG38
2oBa25jRqfL9OlTftYc9GIE8vCga21GhmG0HXi0Qj1sf9WsJe5E1e47l5zpOT+4w
SVQ2HYr6vMg/AKe05D9Mh+UAuIvfcJpu7PCXZ1O8OVPcX1zYT3jpb3scNz2CPaNO
loAq/XCHnrbsCqBPMS/KsNGFgIajKL9cCXblsxmkWdDHA6nP+p3DA/Vn31D6p+Bd
eMX9wu9GlL+k0kpKEtk6HdJKMOcI8HMtbgStDCluZZJ5wjeoL775WRetzQo4DoOu
kOoEVOYnPiv1uTVrq5hY0Q4lyBugsiGwAHqMJ4lJapycr2mMll0SeUe4yk1t1/qs
Oj7AT8IGFoZvT9p0IPSzMy08ub7uZcC/h95ay3+BGIJCVRoeWfdeEiQCrMJM4NpM
IgiAtDUWKTTvKA4BF+VBipgkkpCgMUgPhNEkAynZ9+GVRrwolK59xd6J6x0IvMAl
8qVrBjKGtPE/peK5yw4j1Zj3vf3DShrUXgZ36HuaYE0k7iwjqKT4Q5duh63FkzKQ
zoPEPJTJOoJ7RD8zrMwdikU8H+OfuzcBdFFQUwdXTno1c7TWlxzf6EdhOb/a6IcT
kfxKC9Ll7Q3UNQ1XBqBtTeizA9ujzn2/I+B5EbagSLKgA3ExgmmhcUalrqHfDWj7
lXgsBX5D4WnNCBl0xNYqkJuruSAkiC4ZRJm1wjw1zDyW5blFymquEdGqaRyfpC9/
5KUxHieAAV4ENcOa9Y2R2aPhbqe5cscRKEcXXw8T+qjud5c2Z9Ni+iGnXxmnbon6
BV5LbBg6vYQHTA3T4wD4RkXNNJKc3hCnIXCTboyarDIEb3TalOikBWi7F/vvx8gY
S4LqpeDo8UZUq0yCMIJs1Q==
`protect END_PROTECTED
