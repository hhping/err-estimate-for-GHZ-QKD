`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rd9nPNgXc/qc4gIrk84AQOjHMdgqYwJV1TZDNpusKDpDXdr53UbAimMUrqg/5ni
eT4jbt0qyAKvSIn+g/HKgTT80G+g0KOuzJfYg+SDOXyN+JUQ8fKt3FRiBJMHMkeK
asxSjXUeWmglQWOBPPSVW7gM6wRpZ4/or6LUnjZcNPDPMAGI02ZKWdlOrlE/GsfD
2nyIuC3FYJIdXdNVBtlTQ9xThfMDvi1foUKU7AR2GmIlcdivGYvU4Tg2BHrOK+am
XCduwohXAm+Kp07RNGWi7JJ9QP0jkIPzBS9n5X1RpP5LVeaf7yZ3L2IIG7lPUNPb
uYc0N2mgEDMt4e3gBATVZzQ8OMLMqFmQg2ZFQ+qmIs/0GNPYL0nYf2BLDoRzTYqe
6PwdkYIiwfOao0q5RkvdMYxjVlSjM/VLPNzG3h7heLxYKG8pPO1WqriEJDIA5C2F
hp/p5LUbdRdYP9JnJIQX28AGRSVCdBE+f44zSNuRnrGBMwQkzCsp+9iXM02VXfki
z8PO6yMLQZmQ36zJj5BANKeD0HDxI0N4BBAQMd9zJB0zcc2/yU3l7kiwZLE5c6NT
XMkq2JcHRZuMXZRqQv3Y2wocQy2+Leg6lnuThjNNROvoGE2vkIsQkOlgK+UtoqXB
`protect END_PROTECTED
