`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IBnkW92Rs4cZAo4az6R8EE6lFB9B9usszDpqwCiPbsmegaVJlfCa5ae7401iDrO
2pJdCn5soKedSXQvTq4YljoXV/z3Tbxv4+TUzKpjT8MfwOvaQepbQ6ZzrLOuy+LW
zkV4V75q+9Ee3viV/PV5Btu/0iykWqzuOCRppw9I2uEi5M7L5VtRBdCC0/nVp91P
h5qIz1FqEMGF5UfsHckHhU/tyfiRcdXxFroTzicMcrTNIhzmdtbrzpW2UtQKUfCl
G9mWozBX3y0B1EpHEKuBtUzTj1HjpAXLyvdzBDTQMIXWbIEhCnSyiUzDlO/CW5Rp
ajcHGl3l5GW2Y5cUr4kGMtKVhZUi9+2wHQKvy844WZkSoE7yJWj1fWkZc66KFaSU
hmoeRANsOtgyNpBcVdfSug==
`protect END_PROTECTED
