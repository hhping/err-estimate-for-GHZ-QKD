`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qx6qpEa7V383lZTIv6e/QWb5nnz3EjDvJMPTNTn0kwdPYhAx9kTmeTXoZpsn8iV/
yZnrNtbc5Z190PVyxapwcmdxVz+GMm49zp+c+/hXjzcgDHWZmE0qlucc5Pcd5Hku
2MQf1bZBj3pIRsQVlSh6TX2aL4Xr19nN9knccWIhRwcDStSRitERyIJRKSQadcj3
f61wb6KdSl9b/t7UkuY1hiOZ8nPoIC7Rw2CAB/rRRXFOlNmNYrrQGjBl45+bC/kx
DRrAXqkglvten4K+iUgAcrp2K+CTgqYspNRJJSpRZ+FP861cCpzh59KD21vIWKa1
5+LKlY+Ek95251PdNZggc/iP2yHZVKpO6DYOOXD8+oFy879QSzF4AEDvNHm8msOS
/79yw/Cl5PfaAfZZ9Q8Afa+JbG0p7o/80soeIcyoet8EizgbkKfdFCqsDf7iCws8
61ys8KUcuxA7/LTg3Xje+9JZQcYqPB7AqQtpkleYOd03odt8YncQGHIXTNXpXVvy
hk4dfcEYNilLwQMD1dHvitQ7W6Utb2SamadTGWhoWDZCLhMOZP7mgYFJ2WyZ3VYj
LL2TCOicOtOdZeu//vtCSKkdTr43+ZaBK5XrlPf6hq44Lg6sAbbNgDzxWS5kA7T3
CoApsHfAg7zyTzr6sRURzsva4Z+tbaOLSYNf25BynQp/aRkNyVe2DVXV2jGVU16V
+w4QZPqIZwTJf/L9stny8ssGtPUAx5Z5ysKxYyErF+/N2I8rDLmeb6w7ZQ84Liu6
76H9cyvXjykD/xy0YnmJGBR3QJqtFbB7W+8XaA6G2REWOGtBmtiMgns3vRHFH8ML
nOpF3RraNxUF0xAoeyTmw1LoKggm8ZGU+0K+Xn77njzZbo+6MnHq2o7gCHpw1pA/
jhMZwR8Tx7KqeXsEBzCGZ8wbxHSGaL9tRdlG4WpI1a8rNYOCkrR07cxHO/6iXLpv
NkoY4fXSSp/FhlBo/T9PZQXyo8GdFKUgnAl/7gbgxhiQzBoFXi7X1jk8K7WrhK1l
p52PFTbhAcImwDAQL8IVbOkQqAm+VgnjpqGFkUU7eF1VX+uuGRDuk1e2RkSrTq/g
1bbq0j6x8urjVrCmRpT+XE1GBqGhT9Dadju2VyOVF0KocZ6eg+YN3+DqiynMRjDz
jOjFB/WuctTtCqFvZJxnTCqb4FDHpqdEHUWlXuU4TkHffATapJGmiUZX/k3v3wqT
+6BfhDySytMJenmSH+Gd5/lDKOtfjoZyQZq8y/ikLz/iVq2C8anC2RzM1+xVaSTr
P5lFQcNV48q3xWn8+Eig7gNXNIKLO6otC92g3GtewiPKiObTz3aKDcZUhgh0g21P
6EG9nXf4QFzPjiPGkHaaodR7ciRp0nyQdZ1WvrV8AWBQGdg18sGsSVwppBMgcb37
3Dn02GXy3FLglbIuh9LK3WkgOdmXXtz2bSSnh8RDNhYtq/8sDrv53AhX5ZAgc0ux
wtum0fE3TzEQkGeeU8DdWweKNKPWnfCVmBNR91Grsg3hVs3fsQAgWCM8KZdw8YRA
m0i3Xwjr9lKPFnJDKPA5Oh2GFCPGzV2CTcx2O5G495UheumpqAopHb1tulief5Km
hJKcYmAmHabaVCoejIzEeeiCofyIbxRKfD+UY+KcWFkHYpujfZnfHVNyY08unruX
z9sJThUuCpE1WPu8yRrqvPzBwO4ZkFI/P2F1XdJf9ZwQW7N+pSmiN/waBglqxnzh
aiYYZu7EYOVbOF5IloJ3mSklC6+0rBGNDmVagMTWTWbhqAlLqp6JUnzPGg6uGnzd
rtv/PTAsnAt/PlOSLyv0ROirT38aPRu4QpQy7mTZ5BzuxevcUceXxRuH+3vYI4EQ
+3LQ3CtpsoEFpbBB72/ndcobfi3lELxKVvPEgOhSfnqK30Q0JwJ5EAH7EyuUDMGQ
uF5FqXnpqNcrC0P7Tu/RYQSy9mpzE6zWyRqc/iujBQczGQdnXgU1b+DcPw4n3NAx
gNXAWUE5/UQ3Z6wYXTYBekzwD++vZBViB8slIhGu9f2Fv3G3lbjFpQ01S3qd9ndE
r2fZY07xb6RKZ/n9TbvJA2rz6l5LyKRGVMnX4jAhhD84LEb8wKdgkyZhIHumiX1u
Qf3Wz3vbn2xYxU58PpwbXSsx7+2bWZNTKewdIOcbI8ePxNPz1PLSs79lyPYp15MZ
kiZGGAX0X81+tGqtgMwb3kxzLSNaJE1/oGKo+0jbM9J7HMGFq5ga4p9MUt9awg1+
6MPbMA8fSw+83yCbESHOlerhSumeqFF6ByyCtUh2ugRz6wXguv9H/0reBQ5IKotp
xd6jgwkmbwvJbGMuiLgaF0ITHKs2MFKynHX1FH94+0G+c85YfR0viTx2ohdUGROD
29wavprYghUu3w520mozDeYfGwZMH4VbizXPC5zGrf7iwtJ6Ece5IDLXtRhIrX+u
zg9IZeL52DvtshFwacicDflrxA4dXDVkuk5npPsi4zogSS03oLwuTC78gPhQeTDR
lYbMfK53Uw8gnu0oiX9flXbXHIlj+evdRzpBsquOFbFzTxqPRcRRk/Viv7BpYPG0
H26EC2z3l5A3f84u1WQoGC8Ds4FAouErW/u/qIpyaTKqbPuMny0MXgKPy+ce+QgI
fAGCGtdNpnck56CDIEhITQ3BmAXMzS0as7H1rr1Z6z5vSEc95szqd5J0gGeEgIWD
NNe4CR5LT3r+QReRxmz7JIHtfNZHI8m8Y+fY6gSGj8BWgyDmoD4PrmQy1oFS4htL
/jiGNKSdf7otoj6wfXf8O+0ck3TVvcR5XAIdc5xQcq2n3R8gQ90/qIXTmprv7yvO
73RY7oGS3aAEA6p2EdnXj+Bns0fPFNxUFMOns3pBpmHGyjHSdmS2DzsHdxuowSOm
buO5TqazmH7ptuGugfNdokqS1n2eWjsPi45kEn6h8wjZqqxDWiUdJ7B6LDWcbBfA
4wjKjSPhpKdjcRsQDbyYI08MefXmVwiNjf7MAmZ6G+cWOXb+2PhEDGTC+2P7aTum
fQ5fZ+3sXkh97vH7ma9BJSFNeO0G778Tu6faCMTDatj1v5ffXfhNwvMx2+4J+MLO
mnys1pOthR4oL9LKWlLTNtThuOEm8HnDrZ2Ws4vclydeA/DKa19soi6YdtbVoDmv
CiTXPFnXUSleWEo/2xKKiBgXTphokMhiA6GqPCfHBaxEMEuQ8I0suh2Py37gpaKR
gc/0O60BTpGjSCxbPEO4Pt7nMjGFtuLdzJYZooqZj9YtFwvoMETvg4v9wpb2EAtl
fJ9zNbCZuZbFmoCbtkDjkIPschRn8PwBl8WE6IAJtr2E55MoAQ0wqIAOzJfbKxZz
NbSLm0jHGEQdPeiL12YUq4SpOeFef3JcWufGT5vnz1CP36eNOZoIq2cuP8BbVv+T
1EFGjceURW8f2QcnYSQGCi/+cOo7z8/d7ftsdrt/bckDxTbYylGcrI0U5gCXJh+C
JMcbYSgIs5duBW+WQeDJkDuZMgwr2EFZQRhG0+peh/Gqll2Gwof4970Y0aeDHLMC
Pv9jepqwu3BQ5AJQhOZUa9AjQByd7/KaFdkrY5UdhNNSRD+/PF56JQrYTiuOl9g+
wLF7YKanK1PEjFAMmCD9lXkDqfcQFzz7Di9qhDQFD3bg+4KwDoTDM6N+5zKvWdU3
L5UCQqI8zIPU/ZjWFoIHNQsi2Zqko2lWDT0366Z13PlwoepELqGn868FEOHutguE
PdyfTIOucIE1KwAua24n8Pzq8CjGXVOijw1m7MmgOX1gB+x9io5pLZTQKGnNIXqV
RTbN/mtnyPKwJPdwlEuD14z7eI+Rzn5leOwosGj6ZKuKQv5BQxAZbN6ixX9pHbky
8t5rhyxRuB3ZTjmRd0EmB0hvAYhDBwfll4+62KeIT7k4DrM4DvSWCe978Si6EmM/
G2ppNnt394Wb4IpRDXNBXYEQaEO8OLMVSmAKZ6EWN8fJoMilge24BavT2N4LSdql
gyCfDONP6mt+8VAjKEwbGO2glAN229FlBRRXzzguSVU6FQrGSlGjDcbRyFjoiSsJ
xZvdjfJz3pWQeiHvs8YYO0HIRyFDBB1HTpS0DvA2HSesO9rrUEShbCZv+bZfmFAr
IswE0Z/XrB2ntYtMSCNZtRj0NmC9xcLmRqqKEgSjiP4mcUD36wc2JUotLt196Xgi
QZ/w4GPPG9E8tCXey6a4YA+JNK1JjW8TDEMlpUE+1voZQmtfU5E/6w2EgicVQMAg
Gdn/yO6VhIGwzyWpbxa0TG4NRGuLMD2Qg1wEXl78kL2XpJG74UNbjF2ifUlRbYeu
egSEGlr0P4wwBNikJBMXikZpf2ws6EQo8X3IBA/1QHDLqdenYsNy9JuaZadY4gXI
Gg7RRp13J20JVyQwxkxR2+EJLVsLT2668D6jlRmqYlpShC9FHbED38V0bGV/+9uo
e3aoSZs/IvD0e6zJN7TkrBomgNtlP+t5/oBFwml206gnfjuKbW37Fhk30bj0JPDV
A+iOu0Nre6GCwk5Xvlc/ThhfdLhXnJDSYVYXegwgqN6H4BNBp97dRXbUWBUkPzYi
xy9RAl/8RY6ao8k2VOmWSrSeOlvogV9j/kxbwbmIiRihtnYcgkEYqHrcieGPpzS7
GhXWj8XWK6RA3jiPh9IWB85Yc449j2et6gsaFIVz8eghMrTa3VFZJENsH2jLp+BR
lYi1/zfKKkT74oQ/YQPGHLCaVNDGz84LV85tn72vQWZwCkWIlSvrs9iaXW1IlVoZ
+7IiW5bbToP0tf0/PyE6Wf8wYBfYvpTKfREXpQZqE6Ms+iEJZCrRS+230utRpkH3
avGnI4RSRLS1yjwEOdXYBIbPyKofxOt625xydfW5IqNWITUT8tNVp0xjxOX6hdG/
MTbOEZfEI5uj8xAWaCmIE/wEoxqaoeOV+AwjQgZh1L00fbA1Pwdhifz4Rnf6KiFm
dXT62kCPZ7A802NNQ6DnMM3d+T9aETBpHOl/XMd517V20czdGgyxCCwLNnxJ5qtD
JjqWTvb4cJ75933/8e4xZn82bNoto8SA4iMQh4isO3eXbGszgck4POhlCOa5lp1i
GGU+C+5VBYS6DiauoHUWZaLh/2u+qu/O9ywYP68/mxglVShTNe4XufpJwhubQ+HS
eYgD6pQOWCyeKO08Np2So0QvLFaGLS2CUhAJGAgMO8D1BaJBWNU8GekSwHAJZdrH
IpHs1wGVPnuPsDJg/uehG51dlz25jpiymyCtFcV2C52ZQuTFhcF7M2iNRki8qxOQ
rXVqlNPUVFxxoMCynpPJOuIMk6llOiYHQn4SWfsUfmeBA8ecfCKxhwAAnjaU37r+
S9gBHdpDns9nrX/XzOqR6nZWlHtE0+wggaSHSO1adwR9LK9gt/t8ki0LdD8PpWiO
eA4obnMFeflMSDA3dvSjyaQxpo8SJ53/og84WgGbDzC/yklDPWeVeN5C04O6f3IN
AkiGw6jLD1I6/xHcIqUvdnPIrnnNJWbAEDasEHLbycF300Gh1K1zliPUAgK9J61/
qr4OCecrKx1CaZ4eqHLCO4u1uHCLNGj7dJCGnKXGgKBfjUAerL17HJ80PyqNWRpY
upRXyHWenJrm305uKEiGzxolVtvfbqmG822BpFOEw8n5cBEVJj0EZaJO3qzpMAPI
SPW6cxD2w579ExTRxaTzI/4E8xPK7r9Vx6wiZYvzcsenH/gAw2Ws8IC7WkTqNf1w
Y2sqKLKZsewxlNh2/YBLngNaUuPzqXI3POc5yL173jhH7i+MwsoRU0qI81lPRj7g
tnHNML8TfHemzsh2ZWYvbcB4H+lM4p+iSQ4zr03C1m7TWLD2wCa57zKEPW4HsBsd
wlwG7k8cHh7Ey4Hxx3EAZZhdkF55dnEZGWbU3uLbR+j3+LJFMM8cTropXp2tIzni
UDtgp45UKmsAmhsof8e4KH1qI8XZOmcIw1DNFmgT1YTY7bJcVLPWl+J1eXn4J6mo
rBINwrRcyrecLbiotoWlwz76tDmCcFbbvQqCGPwv2PYZLRFplQKgXYERLhmlJ+I3
gZ22h3+2LPy0JZNU3lLxAlKm1QBRV8Iw7/BQMOb6WCts9mvBX5Aku8qINVazZmq0
mAzru7uQoWpII7zrcwrH9w2eUjWtDhRxJUHvZE8VwZ4rldDNKWfazRHiiSMfDg1k
pVxwsg8XeHkw+Q8Z+5JfkeOfIll/wT7JbCnHXPB5iyUAkLeSj3hjkoWfQ1zmi7/A
tzu4Tqkdbz0A6ikbbZYq+L/okoR0JMz3LOI7Ot4ewP3PilPAuupxblYIvi4WDJM6
ifzQqcMRCpbHyZdOVyzUWHVlJmPN3KMhZf+XA9buJ8axmMv8e5IrxOQGGp2Z0+fZ
fVsl5WkbTTgL17JuO2aDCFvLa6wRaw+jmyiGQfDsl3Y9bsVPPxNW/pums2C8Px2R
2djQ2O9vPixYQZVJi25UYdzT7bG+Hfqe9l5YmCqR8hDMKZU0ZAGcjMdxKsF7eeeU
6JWmFT1acrl7rToS6kCxR7ANy41AVdoEwrOUOZfuSo8GgaZyQQazgoZ8NWFevZI/
mNN2boKKSsL7xx6Z2FWTAL/xLs+jAv1uxOnMkHU4fhlnPjoqvdEWb2WN6WmZY3cr
pe07Rsae59MRafe39LfvMYIXaZ7JKmSnC6fFTqP0d3TRZW8E2HB9KUoYOvzeWZ0E
cr+bTmPPQdtSq4KisdAKM8J2VHE/IAql3axNWr7BCujHJgybEp/MkdGgTJMEQZL+
YcR+eXyufUALReqVcPWpfTkVr7NwFrZDKzCFOcxhurUZ2trP2MTORgls1aviZSYj
p80+WSRxWBN+wWb5BjmAExwVWqgGyBj8IsDEcVKeOQB9DeM5ckLFIxegK96YH2y9
b7OoWr3uNOvbF9/5UTWYfL7z8aRTeviAEiH5LeCHPwoCM/IUvJmbTYVqCbEmQ+Tp
DZRiBvakPUMVisp8LF/gNKZMPMZ5WKoAaNevhHs2Dkj0DM0HhmY08vCNTMGw02d7
zTxAoKctVFIlwcVH35LEWQHXGGkhNYg87Tn8iBtcs5WRJprUpYzCW3hLXlkWmk4/
bt6/z2ER+57PmZLvHUVm2tvLRze/7y45XG6HtNT4JE8z4M+KEMuz5VhmgxmcL+xF
KvU0yYEJR3EUFJCp60UJQ223W3Z/NKp6wTmTvXVu8Rk0bPEXpA+Rf+mget1Raf1G
+siPCBMpl0PgkHAgjJmiMhMdqOCVl/6PmOsCfWeGnzzjrw+p74q0Bexjg+bORMfN
lBdbBWghIF6k1iwOJg0Zo/h0lKgDSOWrivj/rdmzHBNHnsUN7b4IVWI018jt0qtk
D4WKs4ythkTc7QKy/+8OKb35jT5ZiQBR7Ejn48/jR11S8bHe07Znv/hRWgyBTrlu
/uBYd/5kmtnYGAg/RJdWAdTQJwRBgn4+xlYiqG2cz/Q731AxnX5IMECpioUJtS3d
6iw7Uq+4uvvHow0eUl6+ZNBOItsaEY15/z/s8jiDyXxbeZZnmGToKcIegforNd51
e3D+Xx+g/XP1pvW3Y3YGIYIBrhqjSc5UHcL8wOoqfq2J8OV9+D6v0GKWFw23MQng
2MPsPy5v9LhvGVQCx1YE93RaadMuWALO5PcjOZbAP9HtUOeW2onVZ11G2W+nz5vA
Mebdt5f969d2DI0lrExjjK5HzGU+LBR8sf2IJUuggvzNfFH3IUs3ciGHfwA2KjOe
ZTGqXFQ0MkVuc37h7uzyM9hdQWdNG+scU/0hkV0FvW8A06ch+GBYWzvVflQQ9q90
CusC63ZzptpLgFNrc2QB1JRqF4OqargoGYhbiUGo2p6KWshgU+JJXe6PGGlX3pp0
e9tW6G35paLYXUeNK1qwOb4pEYaUHOBAuko81W43qUeZOIn60Z1lkuEkNl5nNiSd
uhxInRnAX2G4Y++8qip+4AnIEjN4+3lGiHz1IluTaYsC03jGS/SZzOiElIVdusev
1+OW+AdYrOzt0dUrHLoJ6tHN2J6cgboMT4X0IA2XgkMfYyY7Ah6jfyq/+NVZlRLp
zhkw5kAkDzZYb3bCcNjVDrKwm8NHW6gQ1YfTxLEZn4uLyJ3BAq/CMQMtSXDo5JNL
Fo3sDhMPsi/OLUH1WEoTaOS4+RA0qsigJy9j6reZDf26bqSHhIaLNEvx6UpvQ1kr
vjUgWo2P6Dn8wiCK48RhnuGZe6ad4/xb8NLDcyrrp/8Y0OHGs2/kpoHYFXS4mPPG
Sx51C+G5R89hLu70UPnWVLYrz8Hew9PtGHh+WzaEARtKF3ZprEgR+0PW+zjrmuxH
8lo6uzsWKdPkP8iIVjD0WZPi1Lb6pDc/BBrAFMJG43p+O/38i22rgkM9D90fNlUo
o/GVjVctZhhjq+ZlNLV3/Od3PNNzWThCWJuXSDnJ6vVw4phkocxDj9+KtsnHrXTs
V6UZwLC3Lgf0m/VWo8Z5wPxeNBelsvJkpEloxMPpFvW1p40YXq94Bu5E6kG9+OTu
55CrZ2zOgEvqPL8Vc8KI23h4adeA0eBQYOutRSF2H/RRIBPUK/eHJ/JiNf0vrq6Z
GvGeb0iAmgDupb2k6SZ82eoOHEJZoLo8N+bNl0EHo8AZaE/aPkC0USW1WvP9JTEK
0gi4UV8BTCgCnUPrCHPhmIud1+DpGBoAKVrnvxnlK/VmO90V+OxLL4M7ajN2l+vV
WglndNSV+5mxMT5cPNK+qXLw19DTpIWnKgnWSUqeqB+o/q9wys9SaH7FliuXa4IR
lq2oi82WKD2HRtTaLH0TIc+X65Jjk78OG5Ujxwo8A5KilwdUjHIXU8Q1mo4izhwN
IFBGh54HdRd6ufuIJv3SUGH2eXWDc0X4CNtp9akT03ymTWpAjsva4QhxCRWecKn0
Yf+SJSmWrXr7Mw2vjp1qhB/WCO/cxJO278IIQjNJK8esaTvbLV1uuC2tooNxwW02
5hPEXLQVompowJ5r4p6smjx/jCnopj0a9YJXJplNRjBuPp5ZM55x+8sUrt8gcSux
cy3DEl8BiSIxECLgAPRw2l9IWxqmexnAQldPHC9ZV3i2osAqqfFKSHAQmUPp29Ip
GvzwHpEL593HsGrdJvUB/VsMu7IVWWZIM8WrPD7YCUbgnBlaBzhfNQ8A1D1tItEJ
PpFbd1rgb+kbY0bS/Ich2DkIxYnnzP/moIIEebFe2cUnpVG4c0LgS2cb0dKt6oIF
dbfyCm5+A1Dn73/89wJYb9hMGjABN4srXN81sDQRKL+SnD6QkzPlDFJdqSZjAMKR
EDM9zieTuVTmrtonFSxzZB9mQOWCFWv+i6V18Ei+CYXIYX1eFHZ1UnvGVlnLU4WD
PW4fZxQt6ezGWyyEtG6zP6Yrn3rLxpVeOUkHz8McoEk7oU2FLWbcpnv/RkcFCUBf
xBUH2KUZQ1Tx+ljna9kCyGqUxd2i7n7kkmTHwatU1Ja0HY9T21ujWrPR2L4cgR6k
WC9F3zE6u3qmJ9B8YMhdWKAI+I1ebFPGdXIdJl1QO7O+sh4GCXIG2KY4MTvxp2Wc
oC9Ye+QylmgGASjowbrygai0pEHaVMdPBTDZvpebwAABD7ORb3SJKuInaW1GlAUB
Kocx4BhrhSamzhMX1n3z/1HJ30+fPvQ9GwiXiZXRSm8OQ984bPV98qDkD7rXFMKx
ZStb4vdydD+mKdPCIwMB0m27+RQVQZOoY3I3yvPyGWFa4vcyfv0bDyxDR5MuFZDn
eHEDBJd5eQfXLTCNupxqSYQQT5RHd8Y4bNPv8gS5syY2DuuuVp+FUO7VMDI9/YVr
pwS2y++6cj4o2JNunEZ4lII455fNDRv91mx+b/boSz63vVIdDqumM4aIkvDwRO2W
u6xqiqN1n/UzTIqS0PTOPAXjdc6SrD7PXFJFbDs8zJr+VnndiB9r+3Dy7gM1wFBF
fApnzTzwwChY5yUWvPtjQ57bx4RjNgwvnKedb2lLRog8Vm1/VQNZ+ilCW2Dpz0SI
pxMN70J4UPqTwHni49SsL3v09h5AVVu6dN1UelpGkkP1W9HkCNSzRQA/uSH+rhYu
pvW6/O67nleHOVF52skZu4O/fA3bF7BFLbz1clDEnpta6Om9vgk3M1UkLLQQOfcK
dQQIywj9YJykXcgnaqMU/O9F7TQ9M14HgORQnd1dUBRIuBbob9m9ZLEi+LF2w1cF
UzfV20o8IOdzz1KCa68Mfv19gjdtb1v2NJPBSKyxJm/aHzgMDnDJWI+RZWxV+xK/
snOKycl/Zoh0MftLNQ2LER5iYMSQBQ7amkq9pY2NZgUueh4jpLE78wX1vgtnqrHI
Y25Fwvw2VJf8ny8mnk7rRz4D2JRtCCQw9j7GnKE6IdDySt/lG54QRgnnEWmeMZOn
sLovqOBvDLzwFi5NZn+DDlo8Ar3BCFa0Mebjoo6kwh1kS1ZFEPoMoq5k+Kk/K0vz
bXG7WGXNbpU3ZeXIo5vvQkA1Iw+7ZOXe50WEp4pOnM0xSG8Um2aHrAck0A5AQHXo
vbz4HpKWTdWlNv9fnvQj/CVF+Hep5dBjMTX1W+0ugquBFZEP9a2jvLftb44+b3S4
fOGBkpDtP20Qjk2igRGhKdlq40SiCUsHdOziixonan3Qp9PMGQyjVKa/UF5LUuM4
TuTBqZ5tbJkNlFzwsqQbunhmxMTfDQapHc+XNVFRvSPUmO7rvjC/fm8+v2KiOHen
2HOksCj7tu1jlw7hyW/8Kk+kma+8eNxEICiVzPXBmbDFLfnQyuWJyyKbqfBtK5G4
L808RImoDvjJGu34AIH5e6OwqZBi2nSUkzWWLtRR7c5oBx0KzBmO41Op99O0uT2b
lRTZ/ExmBoRFA9JtB+BpiIBfdZvRVH2q/cyky0v7TK+fiV1L645U5L3+L4MrJU5w
qWLkxvCibN8G93p4+VXVphq9KpRuiswn/ZO7j8cBVPc7T9zXsUHZ+pXA80x4/PLn
wmYd4kji0Vr9ZOrJfEr8C//83JXwI/DChvXUaNJkQsFGfuIYtw/NDgU2h74FnXzW
h1aI6p0QlxSebEuTdB6gpa6vJ4ewlf9OEB7frAAIp6RPGoOCm1dRS/FamdrdnwQd
XTJ6UgP8sNlXwsCDY26Ij1sua2GNy/Y+pTPFw2v2Vm0PqBvf84X11mw52YS11px8
JJI/+sTo78uPJlr9O4S2EQzlGoRMDFQAL4tHeLzzMNMbpVmTzvM/JxZJ2yLEKKal
FVeypGVFpfd2qvHzNiZidWowhTRWVNRPDMPmeKjS7ouoLVZ/Mov+ylTlUy2NA/r/
7YfNItsFlSgnRthDeNcSjwY5U+gyCoafRNwzPyi5zn+BcuPGM4IYbiAjAcKAgZCj
1OqcSwUeIhONOVbI7NvUDJOTY8Fe2Su3frCIPm+NF7HQUqsVfO/KComhwCKq8ai4
U7ACqNrn/8gmYgH4HZudTPL+eyDDcMS/hi4rOy/fJM5HGArvhAiWUz5WT1PL+BV9
LkSU6HNStZx8NbZiA1SCsAisGPbdkmcXkuWrfOowXpat9fJkHJAUuiyTeq3Mh3Wi
C8UglYjh9fWKIH00pqW9s00k3QqoR7JwG8BmLmMmOhlytZBF/gjo6qkqvJFy+E1E
uvFYQYz1hx8OVr6uIc7pyq7yUmsGUAJc35istao0uSjMj8gsL661ar6QrI2zs54M
s1s/o8iUFd/obX2Zp1zya5pcb4kFPnUOEnNaDK55ka8hNytIvXbvYmnGs9k1hJ1b
jV8cZB85dSNiCJyoNxiIDRbbRcOcTKQoVD1lAIPSCeg4X4K7Xv6hth4v8hIuOg9s
GSlqTHsNJMmBWwdrMiyqkRtX9tQE18pVEEsfIkFSnuj4NZ049EoCrF2GRizOXu12
A7E6OWDH7wYxF/FnWx/SX49PnbZgSO7VS3klYXWm8tAuElnayN+yY55aaYmZprY/
zIXOGJ06lx/i5vQrrh4wHPR0h6vP00TU7pP657c/gmfSTqiM+Hgsj4y9MEN9syjh
/Pnflz95ve17czQgknhWoRQFeEOsW3CIQUg3UZxkOUBX8ELFPzeGZkr/wjRbPT46
3mAy7cCTCfU+kYFAYla64TgvCPYpixf55Hnjf8MfW+BFCJbmtpDWgGKt5WR3LzAR
pFMm35sfpazCRcRv62r7/ypWsgG/Nvfkv8uIxHhk9dcKG9rSlvHy1VJnmx9hnO8B
bZDxkXQgHeQ3qXY2eW6xtfqu2fsjL9JS1DJJZRhlHoqq5t+PIAVweWowPhruRZ6Y
61anNryaLBrlz31bNcu4kPem4yOvuGTPC/bPYhPmJDkv4Mth3dRgW8J4ZqBFs7Bp
1MYljkBu2ekr0qEZeaXq7OvwD2P6X7Y792fIZUsl0JLG0ViyaBqdaDQivKnd1uNh
BfMpllKMQcD5g1KkSVfLxW6aU9yyUTNTG+a0LZ2gaVFz7NQzQ7iWQMnZ+n4qmjfn
f9KBtf4N4HwO4CYrqCxkBj12FDWq/Sc8jZuKqwg0cv6n1x89TaeKQfVlxSVrtjVk
OpZRj31UgJh8HnNL2jPDoBDVbLClwLhtszYNb5oE9b+aFZ4gVDzvNVqm6ad0Efl0
lWjePgY15rFJ+QhQ8OHi7gRfMb+gDQV2nyDgcJi8FcN7esaSR2j6oxFo1BQaJTdL
nOLIK9/TkQEq+wxkdotGl5xuhhkpbAnwY9u34c1zqv5vVRzLnuM0NbL1+Q7rsMI+
WJYdiaC5xVvHZhuA5wpHYyms51/WyN5IYr3hk/fLc68+A6DX+HvGqbBXJzDiTWL9
FM9qAeq6nzdOLKdtNMeA1N4rCzwtewFmRAFZ9XRMeWW16VZAr0iIO6PjmeNzuPuR
jS8VVINMB4eRva+mszPBYiPGBX8ns/fHA1LAvO4mEIE42uMVfssL8MNuI8J+GbMk
/ZLfTVgkgwGb70YhWOejGGsUHVvt1KBMmpNO80OdMAhYJwbjHMPIcM+FpCn8vRCk
Yi2DYM19CdWbJq4rAZrbCEeecfsrK92A0+PcWoYI3SsBi5sR0yDoc8GrFRrvuXcz
obRjhHVIDGtkG0JPu9gGABjG7L1tvr6SecuSTa/8zToLCfWeEVIO+QO8gAtbGSiW
vYAdCCEGV/0mJsz7ltwYbuQuT/vLuSHFWL3LyStUS0dCclKQHcBeJulYrxOZSJTt
1DtQ1TSvDee7TD6c1mVyu8mkPKv4LNPPsaPi9L//IRU5/5/hKJ/18AN1np/Pjo8N
m7Yku84mSFZ+MrTddc/GAJuSy2hC6mIXwBxn/YsX1wzjnTWYZZzmyM2Czp7lY936
9HmumIkhYxnap7HbQp/cmYWVHLiv7MGa+oxuXtzcLqsLZISrIJzwQHs/QnvfnbvE
PkMpvqS/TiPl9EVzhdeNsiD69CUczHmfopFBmvItGLi/1joB8y2cSxmGxlJygMaX
PgIIDw6RQRvc6z7Be7d0kqVjUjN6zYGCaUIvTRphfv0UYzj3VQbsB5ZXGB99etJl
wxDa/Z2drNike4N+zhDdxQGkheP7q6/uj55zTrKKINGYIWeua+nqT4zapRkzUIem
qK5Ozj/Zj1wz1AnmYcgC0Sv9FKAmBfKKyCZqTerRv9RE0OVr+TnNSneCv7kqMGpD
gxsl5lwZI0B9lfoQPESJl6xZyMCRpzq2O+dWGuAuRda3PL6vFLfOrCbpVLktSuC7
6nT56LWH+ax7UowHCBz7JbTO4UW2J7pt47vxMew1C4wK9ycie8PMe8bSyeAylMa+
sD1TLoGCbtFUGjraYo/Rbprwnzj5rvBgCumuD/5Pg6St0DsT1oRjRJTOaN14BHJO
KXFgpAhF2/Wyg8m3Y/7NGXQmjXjh0ydF4M9GUPInbgD2xaDIbuh4LypVjRTbebJp
qsoY7OaidUMYCtctu5uNMgdlqhJruRx7NBxiob9Dfm6LGxhhQT+qOCI3FtjgKvVd
/iR17O9qFrtUmVK1w6NO1c/GtsdaXDbV9opvFpeWjDII2E61F0me+5bQz70cvMQf
aeRSRjD/Umbf75BckmbQa419nngUerK8XtRO4zGM9ydR/phBemFNo8Be29CIao8M
bxVIRNp0BgCCNQ9J/kDmjrTcbSDjbQuXYl1RbFotnnvjoUb2+PK/2ilm/9O1ofKL
IBQTqmLS4JhnnssnfaFijJq7Rrm1pj+SVTKe8Uf8VoP1+IvBHVxjEzCnDa+u1clP
Os0hWeMNjavIgy2xZaJX5/eJGvkH4VgsFmdR5IvbMMd7G1Ew/GNzvpa5O3bvgigv
DxPmwgjdYAwE0KEsofmoO3t7NoFA+b5fqEhsr8vHQk+zcVISAJF/zJFP0nxfDeO+
tu7dNL9dxWTp5kBN126180mWkxZgxnb+3A2uuFvtxq2wfvyvLat4GPcbyVo/gF97
xzLB/EpZv1Az6hJ2BCbEkREhJWn6VL7bOa5gSSuAUbQsQE4le+VelMuEZ3s4Dc1O
ILACea7ZqL2VLlEGFgs1SavOUHcX2D2M1PAoQMGq4JrqjaWVQccJA8eJ6wWwZWwF
E0mRyyeDR6Xq/hGIIsPYLmDAbalWX6Tx+8Tv0Uj8Ykk6Cih/nkZoOV/2xZ0B8Aw2
fyd1YDDZ1qEQ8lVg2ihz3rdc0Rep3RazZORnz8eofaRQItGUK512tW6J996yGmCi
26QL7d/c0hKoxVoAmmrTkBpxe5G3GaBjVAM7voqguD7eelmkws8FntgNYs4RbvXU
f9jFcJRCiisrRxPhgn/hd9XeililPFTXq5oLP7sbl4354hNFdc/gPEs7xJafSmkG
Jue7tUwTYaCyxK+pnSIRZMOc26ZZ1vTBdafQDjOHz2p/QWav9EOMBFPDgGP1UsLL
fFsMVkgJLSCWMB+x02ytULIcvHh01kH3Sn4YARoiK0bCN++1BjSLpMPqQmfW+CUx
bNeJDIEUNoDaD/eXLT991hX/7ecgvXWGgDbby2aJL5JsdiIFjZxbBwX2e2GnmoAf
BZtyz0z7xuz0L1S1yi9sNd3hFqH86G6yQPM2J8ymUuauMFfR6bGS5JLRUzZMW73J
mwWqfD+BOz2BIWenXvr0bmtCUn5EtiJvglqRzNAif0H0EtK05MDo/Ev4PqWJDmi6
wpbixgL17O+DnWusgaZCH20/B0LlQFWFyZJo4XYlvhLWupesFkpulma9S3NrVIAF
iusump6lVW1dSbHiH7upEMu70h5J7UJHJ7XCKFb+TWTRbWCzAHCjW3FIz94W40bV
UBIMlSdtblhnOUF36jOKkBXLND4skx1MVqG7B8e8Oo9TgmvC0G4Ijc3zzOHPIDOX
FSG9JBYUbsC+yJfUIzwRRTJ7yH4gjzFxlZ3sNuZ2EveGE59Nw0e1wB50qdLp6R3b
/KF8zzqOmJ0qQkfHHymo6b81MJHIAdIZPlsw/PcbGSztAkmzeE/G1DpqLPx/6/Rx
ATO4mWqtis6W0nvU5tyf9O0m5J8sAqeHD703ChoqLj9r24vGvxcgjNNtp5ZqzBOO
vsQwvlzrBbJfULQDTlLNDrjf+0MumVTuyg/I15ArdJ31G9vSRg+9CMgj1Pquo5dS
Ox2FYvm32lXGldyjkyuqasjaeG7fRPihP3QuZ6e3JBL9qmHFtGaOLZwclELpHAFN
5HWA4ZG+LWap2kruuiXzOUg5pjHy5sPdQ0iP6A5BtV0pn9tubX/0e5q7R2gIKE2x
mhIXZsJMX5bsEVuUHCUYQEsFpXpRDZPxyQ4M1nHZR5SrlPlfeV1lixg1bwsP+JTa
duBvez2m+4eDyC9VUbvrQteUvJQYk8D+oMmeVoFflTs+mdpCnNVnOi6X27cOF+zK
vPmyyVlsvfVUE7ZZlR4/0ECbmFEYGWyM2xPruERA3GAKWERzHGuP/e3XNwe0EI6b
YYEgwO+v8yBptGms/b797TPqGlcM0kpGzC1Qd9fNCP8gxbnztHck9Hunzm80s7As
/cVLn3lffMcxShV+r76x9ibAbKEETY0SMTIind36TAm9ReLmcxjk03qJrdxGAMst
8aR/terlG1Rxe5vHR2KuHRtgHa5SdQrm7Zlk++SyPCmBvhdJZ5eNWVpVViVW1qOc
iCBqP5ry09fkA1aXB/Kq0tC78H+QDiEPanBo4krrYQaQcTKe7i3QfRRe208glhMY
Ksq0tDKsxYkwOnLHefDzlOKiTv85PtTjM7sUanHtULlUoEyNM0ICn5Zqyfd9wJO5
wOk4/pUps1dgU+CZB8r8Z312Gx1ZYcMvQoS6zr6OkMIPm3Fq8PiS/KbrFBr0HokC
nfuWhxHGUJs00xG6oVtgD/7ph46Hz6mxxzdPiH5l00LrvrmlNzLwPwc5IG9Zy9mY
rrKBRSGgIyShKqinMQx7UT77yF3Q1mCd6Jting995Ak+ALTN+q8WqdWTp32h+C42
BVCTgsPI1vQ8JHeWU0194ZdsZWMLA0cXYetHfCCOQgdBXz3Xk1cjv0BgyGQ1PlOO
1mBK2grOQHjKs5BedowGyModbUocD2jL8DdgOfPHQlMpJeWwAEM8Tj4QeaxtxIMX
5ee2E/Eu8SP3UqOnIDeYAUGS38TNvKBnYBZFjkZSwFUy5tSKdQbsACg/fhQgj2qN
9Ww4Rts/KTT6nupYNXEU0WKBJwSGVxp1OPGl5aHZAIal5w+s1KFZLI4Ct3+rHErV
wtueWfLCit/MQMjJIDePYrJCG1jCzLOKrP40aSqW+0WswbtAL7d/+8FB64fdGOlQ
cOkr//JliSCxVDbkM3nPiMbwLeFJr2Ik+e+VkxsIUZU7qxB1tieRDpOscmYLBbA2
+G3qZ0a8o++eEpbHSwKWQmI2YtqPQa3FtE5nbYU/7mq1VMtspjwL+28Xk66nInAC
VpK+CbwPFRFiFlKJBvyYTU+7uKcrIfu40GX5qNFTWGbgHByBfq7DPLG5UGDV88LS
H6o1sFIY7w5IdANEmaMq7nfHlIPUVIDmo8kn8c2XRUNXSrgifq9eEOv19oDOtBCD
+eP+3TyzepsnZPL+jk3fOfXFZ1dQUI9lIduwGNMji+ySps5+jqx0lDzux6VcWTPl
5PzGLMf0UN2CM1RZNYlQY65y0oECOWycscMbsbSXAJYWutP/Qbaa7V5n0cPDYSka
ub8puAYGCscTSiJtykt2az/dP9g7I4iN1FwdKj6/ayBA7rbOw8CuzbkUHYpVuxMR
LFn9QSJieyLnWafZ89byqgV36/Eu6wihdqceXNYTAYy1c8+03pi2mfIH+aBMGq5I
7EB0WUS2couPTl8ZBHHiHRtkXkTb5gwwWJenCJrM+ca/Dd8uyVMsnx7iAH4X1Ph/
Cg8uYI/YV27Qdd6l8vc4J4r1OvmEbLEzhlkP9c+vPnTncWXwdu312lXhfaf/GRhY
aU2iBIEYzR6u4SQ3EJQRR68f9JNncyEiL3TXLaw4AUp3XP/bqtc2GvKjZVQFaQLo
MloTwOhn/A45VSKpfW19mgax+zxblqx0APD+iTP6xhndUA9DkFe/OQ/qGFouZvUl
Xmc2Oosy1PpE/mgentos2YeYI/Bvna4kstdxPnGfZe/mWVAm62k6DKzbRak/nZPc
S/ssPJsPtVt0F5BNDTTm7FWGkKmoo+EljYWq6OuSGRPgZPi1dVuy9XOgXt5iVmvn
4AOuWzIYuHB/Q9E4irDL1w2B7aZWVKnC0udEEGR5mofY6AXCKhdIysAA4huAm2UE
onpgQAZSDmRRWs00w+rJwc8s/NoNyqOlHWd8M9A+wjuNnQO9THVN7YMjuHMqJLOM
qQD58tseCGCwz3npzd/eSn6Key/OEwlkCW8GxIoMgXmPGOu3XYMhCcg0ydD21I9n
hRv6RoVaTcZ1iH6a4UbTM/17CHMdQoDNZexnsQ4sqKcGGgcWA/1s7uq029mCs4QU
X+PyXVnog/47GsYAgVyq6zhwhQ/5rno8LMkhBrcT64nUR6L9oCpqtdmABQv1CUHp
yR0JPDwQKFvi3IcCpaj0QHqbzebbGXI0qDVeEt9oITYzc1vbWZIy4oYn2JaquyAe
XBPH+rAX1BubduVanjjtyX+Bz4kkYdA5mijG7bT4zU95WzlnFazg5LtK6e/4i/E3
cggoUvRQObJJea320jaZYFXyeyV0qPyB7pIRO16GiI6DFAoM4eRlVBB63AbainPA
8Ou1pAXzGIVM2k5B5i+D20fY5ZErPueBps582Ual6PXNtPpDn7ihyI7QXFSXqW9A
u7RyLObVajV2Oy4NH7T1dyJuK5pmlbVKOX67E/OOWrCu4IFoYrc/JPySNrBiY0pQ
CtMcO91imG9ba5FneVvBC5avBhEpgeaeztwvHNaqFFdBk5N0gC6tJa06cfu5Ifdc
4Qqsq3RmwesxrGxD+ZR/tSHfph39nEzLDy0eyzem5g4DQZ2Ux7cwVAFXsBcYf2yP
D4lWmwxfTnOckWG/UzbayGGWkmNl6zvC2nwoCIJVn/bSuognDL0ebuj5M8Xtld51
7vFGGEpFtjjL4k/6DNfPIwsH5thV1BZviW7lgmBZ/YKSxIJ149+SeMOOJE/GaM7k
LvQLWdhJAn/GuwkHJgM/kFAgUtnrPOS0dJMPsrTd+RclNAdYNxSYWgxiMDL5L1f3
HE0fJwCgx7t2BdyzPWq1qBvcw3FbzKB2kkRpy/Mmkw3x3RYuq9SWfDH23Aqdu5wf
wMLlo+6/8RkKB+NSzib+5bPD7aDVWKqNMbEF+Z9R6RQkC21O3h5EV63E7aeU3V0O
flI/PA0tQAtr9vUyw29K1mRv4pGCcvbKtj20/hBUfCqdiNWPHHFGQ3qcI+9T5Swx
G42nMtoukG4PqRcPy0ottU3DKb9eX8J8pSN87MM63Blz34I45qCVVYS6UB6EpytL
1Ql96ZTek2nftgVA9RoDNLtffe7mi9M9v8XP+m6iwIqwoatB2AmJ+ceEiTvqoe5S
pHXixx1mIHDhExo39l5mbmJRK/jP/tPzKV6o+3+xMHeTHc+58ON0OHNPD6881Zlo
3hebQQdYddxA9guOFkmdA5u3ORz/wMTdUvldmgJ65gSzoWTpDHFR8YmHWFxHXkU4
iRh2hpEG0c89e3GkpLo+3ZSiI7f6rEdzMziZg+ZtSwtZIB3UvCxwl7wyGytIiR4Q
dtIfz7TF2OyQdFsSy6721W23XcA8FIaYpiSzHXOiIlngpBOzw6DURRzIdfBUOSgO
1lNHX67lvGqEpT+9UIJ9cKLpNyvhbj8V3NR/FGI+bRX0ar+FmpCCsWysMxBbzMRK
gsDMOcuiRAaQwo0C+L4d+pGIihT0fAnE3iyT0JPH3LiC9kmMHjg8RxfwHwFXaKrl
0a4BNR+SYUoEpZzTdcQj5gMDAFRn7SUF0qcM7ULUcVtDYpdeDmLfZL0C+87RVTXe
iFeVpF3ufLImNIE18g+i+I0D5qcAaWZ62wwr9CoIuSmZsdu/mlB5qINu/t7j0pDA
T7WXe2nBQaFb9aZ7aOue95rz+OCN8TKbIQPsIeLr1JM+LmzrnvHxhhoeQvEtLvzN
iy6D5tiUcGA+v0+vjmiPeeENpKhmpFgBPavdcrffKujRg/BQNCpIEorfjNXTetVv
I9V0NdGB2KTENywwmppAD/3PJbP7qC8omHvXYDkaGnFGwiVclxd2YMAEt/V9hjNl
+AWUGTey0bE+A7bAyLIKKU9mxc4dIvAnQK6eXTNn7nLbh8bUJOahEDPGfk544D73
RhLFoMb1OlJBmxrXzP0hRivBdWdvetJfI7F2FgEDWKgJ5vivBT5Kth4ahtPUXpby
iN9RRLfOCtzMWO8IKjQVqsbkX9mlEhvOuh1BaWTAJDFaZ9d7UBM+mrdlARujdfni
StiFvi3Xdj/+4vZgBAha9bra9OzVg3JERNcozKkVo7XWi7Q4ylbOqpAeG7pzoDv3
kWO3AWqt5DM1MX9tS9dOHiJ7nphXoqxpW2ieuM85DGFmtt/5QqyUadkx2er9B1ZF
Kk2msFbCC6e9dNGCVE5yInLHVS5mgAmMJuM0qboz4QDelaWPeshNy/fqIwjULhle
By5uFvDIoEL9JLSf2vX+oRcWKyoi7pz5jRrGSeMT0Go+tECjbdUKAsod9KYLc+RQ
MecgLx1XKJqi6cVU45v3YJv5A4Flhr98PMRkfdV8HoRrckhNcl3p9u5Hr50gnw3R
nirMi39VEU/N1/byMFQT3shQLE9IkK6sKPD2E51PmSlnMPV2CFx513rwT+Ijk381
XZQ/NAxsm59wI4HH0ac7eknEPBgiAEgd+mKoEgLC2AYE6oJuFhpv8ECvhNKTYOx5
GmCHCxvz6u41q32D/WUxssd6UinFeL098NTj9tGSPA3BwNK7EcpwsoC83Eo/ssE/
A58K5HC3yZbUoKq45KmffxGzhA/3XFQbLpj2JOOy0jVqpO7Km9iBlv5YfIE/gPPO
v5k9fiaeASb2JwxQNB/vkPVaZYKo4v4JlQZUxU12AIlngnLYScho+NGN1H1pyaeB
uWKcQyld9DfMZrynHm9RoQKcupHrBWa+BQKfxI7tqYht2mH8i922sSCMl3qv8CE0
QX6DRVuOMDsREf5ttig3uR7lho8/u89JVoqOQ68BnFCAVUQGExA5y7rgPxEJ64xe
HHGbjX57ryLq6Yy8eeVM08H+LOmGroz/f4YQ1BGMlQTL6jGNaSYq6EChTe9TBZLs
h7tiB3S7e3vt0UlEeSyWS4FAu4VTasyFM2fTUCCHw532QCfsMbFhu5nhts1GC9uk
X8a5ZksYXIM3Mk9nNrqCp3nFNcjlxjuv53RzW+7yia5mP/xBcwoE1ac9ivS1nmue
6xQeFCFrxAs7/gTpH7L8UONhWKoa1Pik2hSL2eBKR/GTB8BxfPjq4avaKbx/xMEt
BSaP/XQjMwLfCduWnH4O7uHofJKFZjvEZb/4vf9oSggik0NQXd45ijXPSRXmQXYw
MYpTw2BE2p7auen0cQW+0bQVWjuFfaMVW8VZe4nLRONKGsdgwX9ZFhaXJt/41T4h
LUPDxsQP9VZJpzpRoXkZX7KOEcabBzLIYvnwEu/fElweBQR2UbOctkvT0hJ2VFuP
LLDf7OB+0e2GDYLIYgoz2jQXxOmaWm9pWpl4EcbANIMfmliYlRvtFzE4qwVCpqBT
dBPNeIYrokWTIGe28y3d6inLJq9VQG48PZQsEU7OGKrW5+NMK+6HhAT8xd4b48j+
KG7E20C29K9MH3oUhvoH2UHKEVdWAFeg516reU4rNL7etTEe2539sx6bvCO7RVNN
mJHjD/cvN8irO9qLsXR9aBYO7NcmqUKBIPbGCv1zH2J6uXGqk70n1SDKx1ETEbhq
d2CmrxB917LRjFMxd0BcpP9iK0sRXl+lhXC1Be8CWcXzTQjZ3nZ3oAj8xiA5jXBX
jVUL+60T9ZkLNQj8QAFHXIuEekvW372EPC3JS5anYKjDjtVGdosTx7vilFZVucTh
E7Zhd7u49hrVf8QdPM22c+ZMvgqJI+DI1Iu5N8GEiU5nCNeiBuxB6YcPpzyFJ/lQ
peFuhru+vsZTD+2XuOP2eNf+MhY5S394tGlFB6yHFaaNKguSadM+yvPYeJwt2YZM
Ou0XuCTkRQ8xqfeSUUWb5/oNwixFtok0U3ge1kAf8iZ/XRio4BMbWPE7m8AAPOoB
CuV/4qqohVy6rdc0tIiVycDxXR4UAJG+Pw+ykyu6eGvQrVR5otX3moSMOf8C7M7h
UrrTmm86SALpYL2vNG0KP/y6xmGo60pVqgJK8yP+Dkd1gzD9IqXngpwAsyqxege1
jATSqcln4Y6KRHKsLLGjL5wrfTpwEUbwyXpF5amFLz6W1CzXx38HNGqwCgE8AObY
Bbx0Mz/xLTR4xsGXNZECCDYMH0a9mwG/oB5up2Rd1r5DvnYrVvjJ77VfNexuJUfY
eId6YCJ/PODxmQJPnEsC2ZT38FNgXlOLKaK0+B3XG+SXUgiC9qmZ3GLKLCh3Db0X
qmOmTi27H7dVqEpNUaJin8ekNVZRIIlkTRh3ED4wpM6qSD4xJE+ZGki1jxIxy4UO
BMtAUCC+7HaX6d/DqeEafWwzj+7qeOVvUF34N/aqi6d05K/ST77DhMdDbJWNuq1Q
gV4gkgQZA4uFCCFSmHLNjmi70Kp+kd/m1WZuGACYOhgjw7YbNTZIAGk0XV4onrWt
jGmy2Viqe0WHFBmNTD9A19T37yb25MFiOdAqG4b3TUuyQfgQ6wYXHLeWKOFTfCSQ
SMivoVfulsH6xLu9wysPfNj5IZIlrfeyJFcoyJnA2qya5KIHO8OAoKxvNSG0zWqM
3BxrLO3H96BpTEhyGeW0RU0HvBzn5CdGlmQmVZ6o4Ge4v+71WalF47mnkcswDWkb
NUn3XaLAdXfNt110SibLbWEoqln19h6Eeuj4F+GlXHwXDRN/81LQyqFZaYMJoRS4
yBn2HeDYFl+xWxbEFpOLcLYGa1aeZi61pr9RhVK+1Q6luLaDXJ7w9gwoPy3bvOdx
LPrMQvIp9yAdJCgfBVHXowiALRs9ZlxChNnc+UrzWU/uhqa2T6IoQ7YOwLTAf851
83FfaizIfVe6xZJ/4DSrwaL2xwvAeF9ADGINBBjEYYI6T18TURqrtZphKE840NZF
XuNQp7NlDFGSZacakE/1jnVJ/1GSKw+PtwWBktEwvIgrLEMy3Y6te7cWs4T5yett
GHCdeH7jWcX050mh66CBGhIbC486ixh3jq4E/f4vooeAmlxoGnrMCVtj3Dhv/DE2
WJ4/4Urp+As1vWQIJX17933iWLGytupsPwtBNg7+MNRMoVc28AscfLrt41fqgVgu
B0CBLUBkmpPZRTG6kw0/A/aJhqfAmhR2IAWAN8r1nMzzTXa39n3WuXoa0oPZOY5a
7tdXwSbTswmYSM+U2J057xs9iVbmDtRRc3PsGUxCjfrPvsmgT2IRfXvttduYOjAD
Y6QoHcntY7RlKjqzZDSiD+zW9PG9zvDepEH2LA0vAdtqTPgoUgnhAEPqSrYOXIfr
TftAAAi7FiBB/OzkCLT/8lyBDI/O1I+1sn1inWaGuaEQsEjz6qnnrcIyMeqNvpiQ
UfzEJkg9dt3az/pt30/s8ANkKX/aiibnaPDSCQVxa80RD2yuf+/Q6etQLJLqEqIf
XntkBPliqrwUrouUYut1thVMU/UObh5tOlU7ivooNNQVLiVdQr1rGJOqGID5WzTI
4rOMNZ+bDypgNoyFPPQrDdiQbm3PGW3x8ToHBry6Pn0bA60K5y340acWdHxzoz6u
m5y5ByIOkoapki0iuEj8DRzWS7yxTreghP61bdaU+5DVN4TONkBJcvWEsUNIuJxR
sTIhEtFlF7iVKY71NC8VrSkEqAkw8P5kKzvX2ngkzmi1jOY/zw+PibMAQE4dgZWN
6zEA8OF35wKJMJ4njBfCjlz3pjmAVNZ1JFMRf9+lbL1ZCVWRYnGWGuvHj3/9xiZV
x7IA4i3iPe1x4rWtl1eDkSC7wTb2ZNXqjy43uSSTt5m8udjXcqxHVRLDZ81EKDaO
u5CW5UuSXUB3EFfioUNV26B/GdqCGmTthMRzpgHe1z686O8c0wn+5HggxdXaVj1p
6+4EpMwpN6Dcv3n8EUiTYZ3DnrNiVLI8zAyh+ierrqfymGoPOINXEPWpKRIJFv8T
Bc3+uEh451WIMkWQ/zaGYrFWMfzty7ZG8RlExtS9QD62YyYhTtJwxo3CpgleaUzU
yNgjtqkjSDNFb8N1FJBaURr/y/5w6RY/1FZo/dr9fjx229LUn8OamdDxnifhVOdG
MBKzEc3QY+HDjh9L8prbVjfzISufVBMkZLoSkxs7hQkOGM4Mzy9stbXVbcHoCoc2
P+7SoeLYW/cZ7mjdUTlXYkqFFOXVHXl/LTkixlmKlPaRjs6Eb1NKZ3wqAhwYTrr7
mXIaMBpHZzIHbIwjtheuDpgNdgrxAzbCvMrwQOAV5atv1EgPvDGuvMStZXKsKsda
Kt2jLHoM932CGzmnzZLioyCUyl8xkPMpNIJHNrAxlP9nGbFlrf5V4ShJcW7Yi1DN
TsnTvFEw0O/yF59wUobMLFF0dpxP1PCUwr4FrOfhME4UFB10cpmwfI4lFwoYxpT+
gpr+JuYZ9/oLvpXiXnCxoForhgKCVui9AqDce52zBOjpWBJ5HV2nKvhHrxwgh8tL
4cTAjvV0gx53EjGhd/zeLvYG/Bh9m7b7fY4mOPA0/rM/hVYw/cgWdKO4F3g9mroT
FT+3OCJ8aa467gQ0qZqNAVFjC8HL/V8Ne9BIohkEkSAXWlHsJNKYBZAQEVe2xJX5
ZIXwsT82occwMw5+U5NF8tblPD+NtFVExh7U9hMZG385+lCKmNBzMeH28yeQCgOI
vNHewSD0+tFSFX1+jyRunz8c2Nj238RKjFR+MCu1e/nZfCM1pXTJmrgWtlzkMLk9
JZL4QtlErD2jfGbKpRg7819qREU6Z/Sm/mZ07xskh0t4kYL5j2ZEm9k339teCOic
esXuQKOeFdzuvNTnrdqi5jqp8Rxef2QVDsN+Cw0t4c2gTcyd/U/t/5fq/7nkNiS1
Y76GUNRsmm/Kzsveyk0HD7QE3lIBoZfNI25arKi6SydUfF1bM3udqmrKehyRxz41
B722j4MVXJaVptkWAbW8Xcl+gxU8sGWBOOquyQUehRVS1hEu3QXQEmhVqr78bkWd
OAecd24KSf9SCd/vZ6u4HH1v3MvjW8urizHVEhVrxaK/bhsZTtLcqSxofDD/d0Vy
KUZToAymmkriwvCXhoQufll6C0BC9+LIA1WAA50fpzUpFjqKWqSj9yOwC3rJw0Gb
WoA7elp6c4wHT5HADKyiPIfw4URyRLkZd8nR+R2Ml33jndMYwK4cFt1xh4uc4jle
TipZVy82oPBWKp5XBNUszrIB6pplwayNgiXXmFtMxUDhfMP8BZT96jf08waj5mUd
MJ8RbvKOspk7CmuNtCfie3+w2x9h8ePcaShdTnpZto+do1OxUvBjyrudNbM6asZb
FUcYjsypX0cd9GN6yXbuZXQ2qHCTZc20wASmXhk9aK0LkCm4EQJ3qrixnsJgB1Rk
6dUaHlx2WoHWNcfjQG4wIInEPPXu/dDWrvgEuJ5mBSVCO4CTy0/l08pWirBKbbNi
/Zy148V5mfjGCzaRVTqb6GgXpQdV6Pnl8bQU/I5aX03nTawWJtrraDI2xduxK7e3
KUr9mcyyzBVJYmi9kk4U33M6Vz/6YciRoTPTiLW8kqw7D1FdoCP4JWBGDMEyltvy
j3vOjnaj9NGAF1+R5cwmiiqpfHcBFV8IsPGPoOm51vITvjxMMDU7guMal2wzZ/zy
+rZdBG2jfOQK9Bdoroj9D8INghsQLDJlUTulY5l208pdA4n2Wgt63K4Bc1KF3r4L
jDjbe4cUvd6Rk3LI6zpHzCc1El0e8ZnaFfHpMyASx2AigmPB8e5kGUEgp4JpNyEb
FStU36zxnoVtyzh0NagZvRWYakGzwPY7yj6FCamMWyPxYkXKCCFV56CemYqEDDfe
kFLtGR/84mIdRV4ShAYgGSTkzAud/qqDK4bDro85BeCYHerrASB6xpvqwfK8znqr
QMibK8HLlWG1KbsNIDEexB9Pc9FwjolpQfnI1I2IQ3ahhXSC1PhPsXFctr9gbiTt
ji/goRyAwQgHApqFzcVUV59qi0MaQ6TXugJ5QyMa0AF0Ho3+xmiDokhRarfdqSd0
d0OkwbPiYeyvpJp8GFjF2rdKyNGvuzkdNuCl4KFYPkSeaCLaEFKWZkQEVdW62s0U
2r5ugWFAkYnV3xgAllyXvWvNnKdnSvPDtWvlyC+Wd51aOw8AdQcoKyRR9PUoi6ok
iyLd2ItD+8QNPz+epm6X+Vcjz0aHjgd9Aqs5BJGzdC5cLjZJsMPCRiRkbKCMAlUo
xFJNKH4dqm29uJ+jkTtVIaCkfsMcjLUukQMWc5+EFSJBdxWHLzwUOi/C3nlLAqJ1
aeYQ/ZtjMVoKVn3qaTDAfAyBLCQUDywTOPCyA+rdASQ+bZPBHJNHCFg5QvIviJcb
a3DLo4flwoZDoPOT71IJtX4vB1OGTImulE+jri+huib5l4O8z1nPpqTfW6Szfza/
YLYZuOHCj9Y3zKU67coOov5AOuTsDtk087+c6xYnhf9L9jOK+ssZ3Pm2Sy8hfygP
p86N7O23Gh767atDNH6hpzvtXaBINvEmC2q5U3BZvt1FUGrSD0zOTXMISbUnMFqL
civ+zlzxmwLr26kAuhcWFkLt4m/LlaHNqVEyBWeh9Sqqe7Yzox+5/MDNRSRtIEjC
uhl/KAJmcV6ldNC3Wjv+5tKsDYikxcxoG/u7/tfcczHKWB1FB5TWze/cWyGeMrct
bhWTqPkLrl7vz8sB08RK7M8CODL+hPAYN/CY2/OVvCz/UXYqScGRqxYilxTg8U8B
ofTCN3spPKzA1TR+4DzHRMoD7RCIOAhB1wYehqBE80JSo3sukSF4zR5Yus5vmUUs
Wh/yJoDKE4G4LlOb3jHffaCQmBfK6+M11NcR/brLtSeJMv7Txm20qeOWwCfuN8jR
hF6bOCnWPTRlAMODV1OTpkNBbphFz0oIYJmQ1uKrFoyTU9xBmbgIlO0oTo2ZPDA6
hwZpMC1HMFeS6rG/I99G02z5YgRcfvtwZsFGHPrFzY78Yb7EaMDzez6mD57QJXbY
8qi+Rp16mfJc+xS2EhhJtg2GZDOoZU07dNznYbS1Kv2iy52T57koh3qHfNXmBfWy
3O8SOnKp+lLI1OdTveIF3TTSe2O9rqtPiAz5dbk5kJ4DA0+4YtJzUP9UUgy+9OTp
oooL7u90helh2UIjhW4WXMiDlSHq7Snlw9o6mLRBI7O98u4Fyflec3Py9onwaB/1
oNIeEp5vOuZ4P8ZcT1gvI1l17nq9vpVxCX1ZbZ9pE4Mq9rl3oIAVBzewp2lUQCd3
YkaJJLcg+eUkXSnSPqLv15/BriHvP41RmtI5GvoppQFSYwN+kYc9x+CB6n6vBJoo
IB7FiWLbtECQWMn5CBs7K6ukO+GYYC0KERFtNQJpSehCShVv3sw/I7T1VWkr70f9
4w5ArWmexsr9NwMnmyIL83KRToCgKOog5w76LycbNnqxXaN16fyzC9q8xOT21ijO
ie2W0vyf9rtkjKr/T6b+C6XGXMqBZI4Ew6honEHZkP12fOKIa2frMJoyvPpMQ3Cu
UyI7MlKDaPK4RxY5e35Lzzkyf3jzriiirsNPpsTB7nfRirAgtjfNyUYXNc+Al/Rb
qjkfjzE/0Y2TuFAm7Z0zvd1l0sEzHap35SqqJf57g2pF7BoNlMlWJsF1yAJav64B
iy+IQy5xoRlo92EhgjavXdryF1th4ZFv0sScDVRMZdFoBAdOdOMuHAjPLtNIugKZ
bVEnHV/NDKNcQwwtuQZZRlDmY7dH2NvwEdkpduZ8QFb3dswGQzpnkGmDVlZPPYAd
LeFxosnROg4K3WfJL6cRUcAJhuMz0pdldrc1cKRZxQeVnmTTp5e96kDOODSyV+/i
vx3pf48/6tAmxOttMGtxMp3UuYN9Tjn3FQmOnGv+Mm+ZS61z5Y+29SlzPay433C6
eWFgDuQcNpbUiUqHsqS/wtHQkfXcVBXirwJymdxXrhO+gwBTB16+2hdHr03gfCMU
7l3oZfoE/flf7OC4jfFY4yX4S7iu/6yVPMYvqkCLx/Ygf550Z+97M16g876C4xCn
E+2TuP+42hhKIJm3v8QSm3O4hBaF3wQxvtNdIvmLzSjqVh8EsdVmCj8UfEhUq+bP
xZYb8/S0Gn8qYhalGOSHKgskK9WfqWd/vIglOAL8LKpX9l77WT19FnxlEW6AWv6T
tzpisZSPet+7JQ8HK8HNknZuU8RKG7CptCMmMVY+xv345ME4uKBMVVl6RpNdUW22
AL4/DPT2vk9z5dxrqBrXgqiizPYycxY7iE8SRMdI8UYYSRpz+rkuIw2udLLW3lGA
64+IpYz+3tfLKPFrcRCO0yW1jLnNcy4BRpCYKr8g2MK5VtYoWRtw4vFGNlApWWS4
FHr0HiLOV5qK/S9n6fFQUMX+xphuH+z3S9D66H60RlbzMdQYHLkETrJSazExwZ5m
M864Jq8adJsLNr46Gno2LeCOoVCaVcdwZyAZJbY4eLH1zzs8mwJ8XE4zKhtr5WQH
R6yGYXVnZs5UUfOhAnm1OdVy5HauXTtg+Cq7Ba3uajQUs1+Khc7XD/RmMPdzvekQ
4UqIs0iknA3gZfpjiRWsq9BLDotpfdL+CyiYTUfAlM+1Jhpu98c73WFStieRy5WG
/ABYz8DoGwSPvrn67yFln08XGQj/Oetu6KnQV3fvQlkoJbq7059L9L7XBYj9Gkts
oYPLd8RIhuV/4WEASVLquJm/rh12be3s3Mz4H9vsgxPr1jloQ+1B11JMDTrrGcV7
6nhgfL9vGSaJdZ3pZ53Dp1YUBHrwUyAssZS4gRgdYQCjFT4pFncDI+Fnprq4S5p+
xVVbxZTz+vmirAbfdad06eYgOABrLiVm07VCBj6ier8OMT5ZmFerLLUDiyNKpsHJ
Li/PyeNFkdAAkOrT1BJmOlVJmr6sGr8d2uvoj5F/+lZiiMKJOW0ye6NkPNj4xguH
IoHUAF5ENcJnvMIv9huAQjzPk8HHR6g7iQxZEPaCz2hxBZgkCSbzecISEz4hNctx
rAT2rsYQ4YZ9WTGcNKcKEvcAQzvnK7StUSiRzMOlaKOY8x3BZdbo9V1Mo/tgk+cH
O8i89U7ksSXaX/EXMSKGjYN+wyGJjvBFOoBz8ielCP3PXY48Pa3mDuAGP3KW+eLK
b/ZKKPFH9AhGEQme/6boOhDXa+PLBUVYhhpXoMDPFHg5YU2qSW58SSv2/3VnrzSu
wAXTj87IvroKtlmjuexh6AjKSbxWb9+0s62aViHWQPeXNz8imvzqkPezfSiPPejp
BZ1G+oT/PjH/D2HnghJd9JGa1eOxq898ZgzMhbbVIvQLiGdYOVYF1qsoQYlmQAJS
jkNHxz44zB5NsrXwCzo5KylfMK1eQmjfkL3MaySsBmV8gw2ZUURJzIBAv2sZYG8H
lD5Uc4+mXWoFKCaC/8ie27l/FQVzDDxKQRQtQqEkNdFFlJ/GHfmrtaxySUWI/HjO
0CpM2INUy2HuWdKyVc1yLgfQTycZ5sBQnbryRZKB+sDuy2vYSzyHplrNCXrDlqo9
CFSceZJpdx0CrAyx+ul/BbcQvQXo9FZfz/D/lszg1xUQ1p9N2V9JqTNLU/Gnowak
mXBqBBISsfRb8WIxmhWPEBMFSO6x5BdCUkOuKeG2fE6jFtNKyynn/HfYB5cUjrlh
kETWwz2QSUmLUR0MaUTMAMG5S98cqc/AVGMo5heIMADs1fpB7Hj3IrjY/fYtJozQ
TCZT03QPReHq5AkJN7NLv1zkYk8rmv3lB4uAPdSALT7vLlJ5YiG+4R/wHohCc7gO
Yx9iLjhQVEjG+FS3a8bVW6rM/72uwLf7kfIWAebqf74+RmS2Yp3g15A/6lxAx5LJ
qTNe37a3VwVBV4tom5/ekjrVOdK3F66i04UulPG1dz3r8swaQVQrkywCOJ5bUiVk
aJ9B+vjw3NrStygAJJt8PPsPgx/4Hqx79iXxkvz+WeMbw3Y/MAc9RikviVT/LMBp
QhskxX/CWu1XORzvyusHEUaJiqsyQlZwR0Ker/x5JFGcvzzYxHdhlB70hMl2bTH0
ami42fl8WUp3v2ZP8swCC73f3NWbftxUWi8/YK/tCPRxBTrNjejufWLff7pENATF
8wkc/98sXHhsSAZ7ptfWyJknhKpkRg4oV8KoobRKDFeULA8OLcOWuRXm7+scRqSs
HdRZBuGsus+kj2elqYzAFp4uii8V8KgV3cZUEhNXCmb9JoU+jutx5zmYovWJxL79
m98ZKgejrqDxxdAXzz7zyp01aQC/XQvpVXL4LmguaNbA3p4ZoZ5hyVzhzxzj6ND2
asPRT0cDOuMPiAhIAH6307PA0O28e43JZd3jZ5euPciLAIEOIbLjugMiLy9c42y7
Xuwhko42HRTEQ9pQyEfeTfS96w2s3w+VDyS+d/WOtG2eF7OfAA7hfoolISj5XtTt
ujefd8iChixLgHm0b9ElPLuaH62BlmRmuzN2smve8GvkdhXFu/Sul8Zf1LGTbKgl
0LhDtkzEFc9hB5TU/M2svPh658Ti8HowAGoIYNSW3Y9X2CvpExxuliH1Ef6iY/Qd
+V34UXEs6VwnHTFCb5142/SyXhclnolUmsXmFW/QY9WWA5o0uJG0mPDQlBR2YXGr
tzFPPQFkLCmr/h0/W3EVVufe0JU70BirJr/UJ4NasMLmN1+vb73oDzFAoFjEzE05
wmnEeFv3v45sTzmErmYmmvMxwA/wjdFSNK3W62AEOhgX370wBXQ2vFtGq6vHimOi
7NAuihfmdl67J46hoEPbyj8e3ZMfbPTCyFRwgfDU8IxhdEBIeA0E0X7Q7iCgfV6w
cQmJUvG0grDDYHRQZOHM1XYSK6FNEMftR1ip2N8CkScUr68Qk48uuoANRJjQHTO+
fWKO3GWFx7V1lHmupI56Pud8F8cy4DtWLt/HeahjrX6ZdwMXC33+odWA9wH7K2wh
iwHTnKiXMOqZW1lO7Pk/9GL6JvDNnCZ4fcVmcQnjYP+dfx6whfDdyR35tZUt+ptU
JwrmBg89sMhO1/hNyXJ6P7fmz6RYDXhYMzlF0QlAda484KWZWYOau+uq1PRfEu4d
ATWJGidzT6c9l1E0OvRr+BN5vrfhUliH8jw28Nvv/Hngfy+aSFCqwAkugngRQlMj
SoCftHrNkFqyrtafAUgoHws6kNCIErLTYIc/dEIHLdFITA9BDFfJNvZ1hw/9Dqvj
UG+OuEmNTq4CNuR6OJPxWItVFy1KiGfaELRzu/ic891yZSGxX2kacEsyINrmmuDS
CXh+kS78hAJEDKdHCnA96t/sykL7y9nWT+kGo5Rz03VVmUUlCBXCNZsRzSWy1XB0
3BWokokRR9u7zquXuTEM9w1MaZSS8LewyCJOkAQ+aZL+YqlkYVWkRtAFRsE0+vvN
wggpnLHXmlE/wXJ6uqAQ19ogHxNHpQplY7C+WfqsufhYcQYc5MkAxBzXc3KrLqwM
DitBG97ZWlIySmoSzgCXe1oc8Jn1o4gDNpqqAAU2Znz6bpBmJR8jBi6kxKoDoMKB
nbGLSV+L2Jy0SvXgf0y55unoLJyeQZkGf9VsgxnzeA4rCDwDR0UNDE7/BmLCsUDL
kmKyYEOgBg+Zyuwx9vfy8SrVKOrZRuvRrDqkm6BLR0ynp4ZHgCMVVZC4G60ruSRz
cxekWJyzKk+ggjpKnp5hL3G1b+GHxW/igqqdPcxzjhdF3rzShQwrPzFlT1MYA4LK
nfcFHFsDm1Wd5c6Jw1GLviSFlxYRLbAmSqJqYZ1o8SquS/1KthKhTi9OKiQn+Nu2
LuooICAfVqRNULnRAPrr/lPqQYJ7IGeWQPPLuOajAm76dIDV6LgupgKcrgm4zxDl
m1fg4JSRTnhtHzpHYzzvnJSEr8//w7dUqshnfdApqylJsHrknt0ICTFbn+jc3g9T
nj4eWFTeBL+8eBARmJZ2P1ATz+nN8U4esNmbaHri8fBWSTYFvPqChdYB5ho8/yHx
kw2ABYB9cdzAU4ht5B5I4FhKopX6PQhbrWfZGzngnMTgpTygIWcdxlc2t2qAvwKF
L2u25F4JlRpTJwwNn9AFsxhmII0ylifWBjGQ+jYIBo5Tx4PcQ8WImoc4xSaNRF2j
q1uiImL8fNrQOhNDW/A0pjlTtP6oV3fOqR6N936EuoSDa6ercMBNefblviEfANoy
9TPtsuvydoz536YpdweDzcGBxn4KbyzR8VlIdAcLn53C/pV6LIcD4k72KfcS3yjs
zJVYvHapTMMw0VRDQgeEeGYWk/ITVeQVesEspCUNEygofJp15diZwApSlBOvRmNB
zKpMhdtveJ2HA9Fiz6GMmYSYN6bxzvtAnXkWhDSa15nfOS/MeBa+ddN2/O+tBgRk
KHLH7atRAN2nris4WBz3/Swfuoei1uChLWR9TGLqpKZE4T4qrnzk+vMsYKlZKWF3
LWQBPBxR3nQKGYanXspaLdpp6LMIklbKGWoJyCMGsH5a0m9u4e74bB+trVrg6sSm
csXR/3IGb8Da7IG0E02QFVONj91BU6V5P66b9vq6TYW/xhjouqUvt9F3BPi4vWLg
ncQrKK+oLuh1riR8ecEzqGdCYYkTE7HGCHD1PO/FvJuSKIv8+SwtI0CjfTpwBgGb
CwJf8xLXuPdSb6Xx7kbEBmlfCWwagrLbM3zQWlOfL2Vi0W4Ils7Lzi6Y2+eFgphf
gbDscgGar0WLifPMfzkd0nx5YCAQN2cNgJkHdCTX+ifZ/DSsd74zu2cwvXsQCZos
+nahylqDNiIbf5FYTkuLLuokeYuLe9LgnWPtuUVOy/jVPfe0HHbvskI/PJ4ia9/n
BnbLTncOvyRD3ZU9Aqhzz/4vgih9A6zQb6NqKIdJHrsfkzedCruSaVjxAu9qBlfx
BrIaJt5xo51a9XmE2/TJn5NOc1c22HViCFYe9ovlYaxcaHEIw4xknJMb/f+1vdCP
h4daxSvAWtkclrD+ACWhHfnRfC9lvNvdOIF+EZmW3dW+WHtfhCd8Jig0UMh6BFs2
AxIL7y9SLW2EiMD6UWRNj5FTzk+Tp8tU+UOfuF6C4v1A7Ai3vg62RHY3oVzpHJlM
fTWnJoE+QKBso6CO0wEoo6bR0OlLmRANvgiKfmNee4guNrzEAadl/KDBj8DW5jEg
Lg3C/WRU9xCkKAUBB3JGj1ZJEgkRgoPvxmt3bSR+VVH/zE0ndOxyF9xfwwuYMn9N
k+6JpwBSVF4nnR6NHfuPZ2lNGa5Yhk1jcGUDwpQI4jQU0rAPEx9exIKIO8p2gn0c
f1rSamVoNQRhJqA1sLVjVXQ4JAnsaetfDUspNrIgi2ezECJf9kLqPslI+A7eXZOS
pDsIQeGv8nsyRAmZ06cGsv0qS1FcH5UE1Key8FmL+XX9JQL1uocvBE61fpYyJ0+V
apspnU0RuNYT+pjX9LriussVhOUGY2QtIAUdA436UXDWG5974mUHg04QrYibzMyG
7lQxtP15/kOOZ25YQGa58P11hkFu17eKij5Jo7xE3OhSp4KcTX+zVUq5+GoMddyn
CBLyQ/GwfxWsgGWHORfg0miOJa1jMu+KVi15DIYUbji+EcrmsxYWoXN/F3l7jXVR
AMI+ex4/KuIxy5B34ZJXoVYY5aT/jt29CMX06UZdNo/UEYiot7it/6snMu4hAgxp
ffDT6DcUL44jvOIiCSZahjSauEg4nNCHSneqovG+ALro91dYNXfPOAlFtD8A4HBK
0GLoN46PEX2tbGfIkeQDQ7JL+dM7Lx6NaZPp/zjr/mXhP8rml3I7CuQvkh2zC4Hi
BbkHRXuVhzjHUg/qj9TncYb8v57xIjlvxhMdjrfRQXYnj7rfumgr16QCnq2nQBXz
4RcrW9WV98lxg6HtThF8BpkNhx5YzS5ZIkbeRviJ+spdzdUdBgsIzM69t2CXgUJS
LId/ANuap0dOKhO/jW5d2goTzQE5c1ETWPkOHk0/Fdm/mizvpKhnIIGKLVa8hTzK
dY8HS527qTI1v2nMOLQoLyRDv/joKNrNz0xJvun/5Q8HtFNIStGW8JmNzTbHRZ9I
ag+y6M3awy/jzKNn9E+TqU0I9mjjc/LHfD15GfFTzZybvhpz0T55xwoYu1eOsFuv
qhTFrdPIaOZDXI0H8SvgjgpotvMpwJXz86sF/aGd+DKLQimJC8+IxKXjTaI1O8LC
g9bcX9vFCZrzqSo4rXwHJuQZmTGi7G+RUi2OrZU3mMiWO++IBH+ehSlEw+7+XR2d
gsfQRDqK9STQiNmV8M0bXJQCzn67xilx4spVQ8E8G9F2E76e0nDH4FJ5J+iMRrxG
WEMtSsrq8L2ZYExiEc6b5JiAkktoA1QHPhjMNlKMPmq+vTcOd/X77Ch/35KHF5bd
cFEsEw3JWaWxIJSUVYlUKAhsQPUh/CMhdMwrNCvxGDFnuOGj5U9n1gnsobtUv0KC
SxXfkpX5Pab7grCNFD4BsQM0BjsWwgyoa8tuOhzMy2roXU4MkatsLK24SohauQk1
ah+jOR27yn3fTHaAaSddH4If7n1zsDXYZJz0EXOYHbpCTR0ZqZHuXnUlhbhtZhXQ
qODcOye1+PS9u24wx5Y3tSkZdVP9s+yUoOFOYrq6YDlNlubeVLjASq1vOCF/D3mw
XGweyBI6rHf87yhX0eBLkeHcJ8Ib4KQ04NtZw7Zm8DPgxKjEQWV64PidaBIZtDWT
ywcamda5oL01bMa6c47nE8Eu8p+ykVXFh0y7/ee8/+elxOSQr5LMOuVtVMzkbFlJ
aZ5tvxptCCIL4abQqtdiYWSj79PSysHHcehMoMWY5lV5h9Ow2OR8kQwBSbNngSMq
bchjiOG8+tX2R/VKWl9gWGv0fxsdbpMddSF8ImparssksIWLMKBc0Yd3N3EBGfAT
25IFbcHJxtsVJP4YZ6uqhBJmSuXJK00Tq3xKIn+XsHkrSKW3V7TeeNFGSH9KxoVz
m9vYtXRpNgPCKHRJbiWpU+y20JUU9Qf9wkhExmRHIcDz7mzMFw41hj97xNb7R6iV
VYf3gshlVmabGCUZ6mIW4HrSoYHvS8b79sawc/fGTbhK1zarB5qkKGOLcdsYpFkF
PEw0rfdmQ0EHMihcibaToJaIcxnOmw2nx8l1HnPShfLYimd57a/WVoM62MnA3bT4
Nl+uVqWacG+QQGPVdEhbKuu1viPmqxySUgdeozr3Jwid0BLjpL/jGU4x8qqgfRDJ
cHY8uCKcCdMvsNX/iQ28yKipv4BHJTZQLJdg+GGExzJe63m+8mg6OwD3JLIfdhQi
eiyKOxcufDfpQuNnw4p2N85IKLW4PuJUE9/oVulPR3rS04a5H87q5L/a5LmVV4Xn
ZfiHvumT1Y81WyY/moR97fiKlV9U45TRSaOGzU6XpC0aHar22vw3GNrYtrMxfWVk
zrGfAsD0Ke+cOXemIYfGj4yyzUalDcKisYL7em1NIAW5jW/OllkRjF7cSERh/M2t
3dWgqcbhNpWegAdihbV9WEv7dGFi2XSzCIfxmrCAOo0Q3QlJszEa+u7XQC/uOjDv
bMU8fiO2VIff+X1bc15Glc+JRX6tRQpKN4M17YcaLYUEB8F85jxPA8KRf4xgV8be
JRQ0x95Ed3ERevfAQADVMxz06jrkan0mdkoPEliuDGTUC6A0J3DZtZRbrlf9k1Ut
yisB2a/2DEOqzTYSsa11BxnOkWlC+ZvYbXnxvF3hgdMLJM8JusJCxie6gRQ4YWjL
QUNbBihLCo9+10GQR01QAuc9hxLlJXajs3jvv/+gsuKzKuoAzEcifqpRXF6b/ex2
9yGhEQd/se8OKWiwxnvndZ2dNQCOXXl/0Rv54dZzYdUbdPDpWOVuTVXertCIXlI8
1M7/vCDjUz9aBawE5lgtFxZUjOHDKnottaIx2rPi/EIUcEUAH0GDZIz7daVfJHq7
DXjKYAOuWP7Ce2JTeeZIL92ItnpRD/63u/9bOdgR/oDcJgDMBPa3u/wZW87nmieq
`protect END_PROTECTED
