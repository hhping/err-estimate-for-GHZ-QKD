`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T1DwkKqJQBa1nCsrVRi1sTzW9J/LnKXkDb2Ct/+SuBELZevRCyoA72qmSFPHmUz2
xN/hM73cabrM1cEPzPcncJxS0mL4Rs69mxQ1lUHqXtd0hVPD7srL92RCEAveIWHI
4IoZDz/uxiwT+YF7FFy6DeRlmlnTmeNBKQ7gpJVDp3Dvt+T1geFPGzGku+6e4zn7
gWIIv2StstnFIa2RybMCyeR1Natr2RXDwyn8+w1LVGqKIGtrmFtqOFryAv6eJMdB
6L506itN9ebyelGHpvVoeTPucvUkqzz/FrnWX8VfEANCCUSxxmBldYpAJjCjjRC2
x4As0nIqRRfayMWDViqlP8nVhT7Bkh41k8/RsZAGn03DTsseOsqr4HQFYyDD3GqW
4EIDtdZAySEBltfCbAdhWGpIFOKJi6uGhsYxXJzX3YSXzg39djiblH6FPiCKDnAg
NhlTeJNnnaYzqUTado9yEPWZ5uum2zVMHWjTnTlxCKELrYB/rM3qQzmJLNyCJ4Q6
lwK5Mgn3Oe7cU8t9RQq6D+Mo8qM1ZO2ZO4rA36xdttJK4qyhHhluqIv220pXmGBO
WghQxebJiEkWVXPPtSqyB16tAZlQ6/4mRPeweGrjBMY=
`protect END_PROTECTED
