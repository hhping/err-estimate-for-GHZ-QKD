`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m4a5se9lQsS7x9PDIVYVhfXt3FSUnDt8dlwBXgz/tQSegiYD6wH4+LTHm8ADjJ1h
VqWAKkuvxSdSswxefGPYeEsFsiD6/d2e/yJKZZc/SUK4/Lo+tD+TWCRuCtq/59Xe
wyNeSAh3qf5U+AH4sS69R2v2ePKn2SsK6HN3r7ClVfYhr65w5eUyywR6dhM7iGCJ
MA6p3wkB0ZY3V5qaepAY5dqJfyzBtZdbzY61Z3lxMBqWLEzhWQv9RxQ9k/4O8Ygm
t7C77nbOuR/ZlJJfUq/YPnmavINr7JPtb1L+ya9ATaXnpKUR0w5TJBPH7H3HZz2T
HgaBICcQNXKsey1dV7Hr1yb06S6Mt2fCzaDo3oc585NX4W+AAvgrShL7hzHSGotv
ZMpz3Iy6grcUqVzjyx+UhRQSpdXW0SgZPmeRSgQYVI8PNGzMh2w4GlCFsdOmr6bg
jc9r/6hYMku0CBBCH4MsOfU0dBEA2H0OPxZf/0hPD+KYCozAnW7Futrlqg7ipfYJ
pCjwxXRWphBhRe22pPSH9ibHEPv9meUl9H9qyrev8qw=
`protect END_PROTECTED
