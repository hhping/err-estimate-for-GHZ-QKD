`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5BuVx15E/QjMN6yJJhPSsZyPQLGG0O0M/zQP3+J/GGq1hjTNFxjqfBPFjQGbC/AF
mxjhmYi1MRylICrRA2E/ulSd5CtTtLGWFm8hs4uUqyHL321qW40YelevsvX2ed6y
kvsGiT55OLtlzTkT0RmqYC9uL29ZJ4j3c/1Sd2Y5dxTFHR6ce02ZoDM7aCCS1TMa
ft75zjbzMM30RFkGDyPKPYLIorG8p0ElAh4hsnFSWO6FsiYn0zo27ite2TBwV/4O
3voLCJpIuJGT1vXhhLtgc5faSlNjocW8psBInIF+khVCDqFDVmqSzsRk3Y5oc/NQ
Sg20sLVoQJKmVinba+C/KEWZHfh/YxG4/5ni+re8gDcdVvT5Qo+mitu8sk/VpBrq
CGBmbfZXO337ikXpyj5oyJga1k/vkjUtxQduXbpG4Nmkza5IvQ3SuStNHQCYmokY
B9ccUcnRBIsvAmKrLKp5SQ==
`protect END_PROTECTED
