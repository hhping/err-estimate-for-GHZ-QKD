`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hetcBP7sOhhDZ1EzYvgN5qPyFG4yXWtIvvphApPL1k03PghuYLo/U05C00xQXBoj
p5voANYLxBzOZ1ab9L1fwATPwxEzzA4OyOi4gr/YS90MEnRrKSHWauLsDqy4s5iT
+Y4ExNVzAk8hzo4eFw9ZXtZN4FX9DtZsVJGTz9A966VYygQcqE72BciiPOLqk2SY
w464tqE/XcbvIsuHxjG6iWC/zYu6Ei+thqcHfmoLzwH7eDEzj21zDltZpKNbqsSE
dMNNnwEldFOuh6qkJ1hCu+QsNducLzgybHpGd9A2ityRdeuIURz51jxna2FvLx9t
qovveyl6jFQ9Zr9XsDP3IaUOjRJC2NqgPreWTSOZ3HjjVPGbPemSVR9XgG53z523
K+N4/76G38h9Uc5taWzYtl6pHMGrh7Rkb0gQXzR9yltRhDgvUcZ4HoXk8KLpY8rX
cTjnNDRuHRowvidteie4Zz95I3W8HUjt6NbE6AY3mL0veA7rIgI+atr8yyyGPs0l
oU8zSX6dNFGpvI9euVDE4fqizbrblgAClXrw4Lc3Dx6ZsNi4EmmN+BcZxnOCty7Y
/7c+88Qwv3x4vmlzBdWoQPwaj7U9PzkQxYZJ2oEJqj+BrwJwpKx2v+bJoUm70qz6
FRLYGMgX+T5LJjJzJd5xlWtXkfGgSqSl0362rkH37xldCU6HIM8oZNbnxd4yvNb9
JbmIDDJaeUDGRx62E7pKqkhmM1qmpZfYBQIe6XZdEPq7wMtSc3xzDFH5D+4wnzKc
kXxDFQYV2UjoM9JPopOvDYBjlWwMnKE8Njk2uTS3Z0IuyWayyWtwID3RgosrXUdV
1rYyHRcv6ng+gMsosFPsm/ksqgX6vi7fyWjmNaCMTrTJ41k4OTz9ddQ5UsElZywb
tJSSxTygreDkRNNMIb/ayv3ez8RAmQZP1q5eDNPR2XUylcYUuhQUiUZyKirxVOS9
3Hi/x8GYSHFXG/g5LHa7lSNrWhhxCdInS6u9P1c8YNA=
`protect END_PROTECTED
