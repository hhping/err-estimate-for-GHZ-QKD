`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xfzfuOfoaRD0XAfBMZnNCBJJNQypu6rJ1Cexq4Zh+cgo/baiB89+Xat26e4csgkW
CuzkEnEflgrFn82AwsNL1RhqOn1lh5D+K+PpSkuOOEyKYIqJPae/XnUdVTdub2iB
95z5tDG+jQsy47uEfXZXyKEa75wZXPgRI+PCynY47NoZ3ppKbe7FRrY8xP2zL6DF
avWkbVUADP5Mwa2wek3TV4dHCiQUhTsznHwaRdx7HkhiocS67+CgFlEVofrJWFxq
p8zCh7sJpUk3sjJ3eAffAyTUU/ow0p8zJrnDn0pxKjmXnOvtT35Ndghl/Jgb1iNf
azZSFnT2ibP1uvgQ2WP9j9xf83fdEooeHliWC+dQh8TNkI0/BVlWDX1LjK17Iq3h
qfeD7PtqqU5BP4GW3buIwaY08lwfxdt0fEj2dEJyM52xGdU9hN3UrCGcjBA9sU3O
TJd+FrX8sraFYgp32Wdt+Aov2IG7yRwyc0Lw0d7xGoMYAL+3ENPhH6Mm9iKQ+eNZ
UlCb0cq65Rl/cXIw+oHxPHOC477egqH2egzGg9zvqKHnKR/dY7Y+yMigsTNOt5T5
/bBPDj9KX97rk9KUWEwaCLitb+20PNqKzUWeOr7NmHN0mF0eM8mhrC5HQLwnyLN5
m28oAtwdwlwluS+oRm3cjVZJ734WNaqR9PHmqNrFAHKsVs7ql4DcYSyj8UhyAsrq
reLeqhF4ibPj2ktRFymF53V/EuyQ4am9nS7hJpWx8nn6EPSgMNnXEX1b2lavhFbn
`protect END_PROTECTED
