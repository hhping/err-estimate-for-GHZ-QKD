`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
coG3QBPZmHPciARK1u9DyexK+48mmXc5Kb2lvnlf+O5ZMkjK0S8Gh6wJ4CtZ9jHI
Q1hTKmEUoA2dBT94Vdg7j3BkhCxPigcsEjzzYDA1/tuvUG3y0Ok1E0vwAfa98SO/
Exs+4B4On7irVJ8RKL4MGzaKelsYWML9junExsSE9QYIDpXaIs0xtxgBB5CBHWVG
C+ovJqR+IL6n21BjCU4EAcqWIz6HjePe9wKrFiV/Ky4NMqeQFPn+jbgck8HRFF3n
fQr3ZQ3sz83T1wMjV2pjvDXH3rBZMNrX/KOyAK521XTIg+P/X4eeYmjTPkmCllf3
AoQfD6eU2oLPkkDADclJyRHbfuZYm5QtLp0/Q7/Mie/Z8djszShgsGDOIw//GJG7
pBQfpDI43JbzMWZCYOk3CFKGcnuYdeqHhhoLE2uAX+K0qS5ul0cP55xTDS+YaQJb
ubVUM3iHXmnTM6DDduuMsSROYFWVQW3ez4m94p/a4+GvqyZ0bi7wXKhAijX8Kl7S
CAKxq4KRATIKjW69Xufci3K5+y1V9Vh6CxnTEWMTnZNne/mXnvYTN8wGTpuuKL8D
iVCubzK3U3v2SUtyIDV0/N7Pk1J/HqEUAO9yP+U4D56AZwZh+EX2hCuph2k9KLHK
PrwlwCUYrj7cJ4/DOgkMBAbnABZEuOlahSg1F5BpYrsr7B0ceGvlwligFXrC+asX
AZL5qefghA754snrICKdg9mmEbD7JJzCUySebE9y6ZM=
`protect END_PROTECTED
