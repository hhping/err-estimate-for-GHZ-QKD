`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POkujH6sUVFfqJQu1PRhBkC6zfRg5OpTraWzB41kMvkF+WIjnP7sxHZ8RO6ub2vg
G6+Wt2sh114TFzvjdvg1ZTp8MprpbUrdB6HzCvjwSZMOPyR/BeGlYJhYUo9A69IL
fXitOvoxOP9OklMx1qEFO5knF6fs/OpD49MAucl6GDrcNgXoYuSsaidrizFrB4Hy
Sk53Lgvwz16bdBK0zPQbBt21QEASC2BCbkj8PEj3CMTqVUrVtBUFmSvHUMfiao9q
2RTIyhHDxb7Y7E/h9a0y6nK3Ky6SJCpyMPYdDKinNUFZEAHxTjNDYyRQkrba95l6
Fo2NFE+A4RzEY9RyAF2zBVlXPOyuZdA1qapTlYDY7ZBmSvloD9APbIWasJawGKnj
TUFnAxJg3dYcNKyqFksb9DS0gFzn8rxyfV8SJ2hjAzE6jcrXyceXJsIyf1i4tlDH
3yEgx5hydmpdAlVkpkNO+RIO5nV1IxHBhe3z96sO5OAQ9UUkqufJ8ApJbSJZEn6U
38kzlPLKprrreNZ/goqMQhLOZ5VnK+SvHEkUXRaFUJGEjQdb3PE1ExMQw8I8XZgR
3tyDM/ir0I24bSTsoj4ZGyFOIjm0s3PHDVDZgm1WIJOuCxct++ZlNLSapZOIIxLH
cNROcckt8bRAQKbrWjSasMu7kf+/V23kCQMo8Mf8giD4evhXFLxVEmJODLMRusrb
uco6WBGnyhj2rTcW/+WxgnLPiVikZpsyufWybb4YVummf9zIVuQ7XSUp4Hicgrvo
IUgWBNsrTZqvcO4IaYLNm1mzYyUtM1/gNY4DBmP7BM6goG6q9lt+SlFe6YlEcf+W
jbAlaC2EXBaUVzpI4rHPdp+PS295v8V1mdiyo2qvICi2IbQBs6BEZW+idbmVIfIR
7kMWanFN/8ml5WdeF0C2k+8zG+JN4Rohf8LPsWKZ3jEunsiAr6UpRZRDo0C21b6e
5WGapR6XAMxMIschOq4t2+wBNutsIcABwwgdkddBuuMgdrtLIVOEcHHzG/+M1/gR
M74z/0+TqZUSSMK6COeX82JlQ4eu7DBvPHEW+dRn4dXUBV3YMIU6b10c0Ppogd8e
CCBWrIaGhkehljQcWdZhqDBfFRicdaeRypWlsoDkqiDIWFaKDKHwnk6C5sM0Pq1Z
pCOqAF2CSZNvV+hK1FnOODV78juqAFGLIJuAVvFbUIVIqsG9ag5a66emOOYEJxGc
gs14BukcA5ZgimVIlw7XU/GUAqbhDpkwLpwz4YBITaeq44UoSEVZqxnSq1R0UAAQ
By1g4aKAkupzqjZcab89r3I0mQqD+38qvi1dJ/884lDd/WrrF7AczfcmPLwwa+2o
KbH1WNfQ3jBpD8SZbh2tx9o/0kpefS3IPmSAAlXt4PoBCb7lMMJLXBLDlzV8+Ivw
TnWU0miDaNAi9gdmDzS35waJeuw2rFIVAXw+hbl33r4RA9BrswZN4321/2CpF0Ty
I/EFeXvR3FeBHUbm4KV57g8fLH5q9fxn+kwyeY97H4tW9ry91kMtpBgKS3E2ktlV
EQmkYYzhzm6imvBMAyLeyJJWYPFX2BbdnIKptiDdKrCLZi+JqQviaxA0FPOGVPjb
iWsMCIIqB8bd7iVYIMmNx51huwnZf3DX5EQeq9c+W/wNtBRzEI4XBa0HPDNmA8i6
00AAlnG26sUjnPcOxBsRAKELFhonKGhZz+gHXioRLb16JiMbmGBKusS7rZf0pPga
gM0hopR+nZJ3k0bcXfd60WqxbHhZEppXzHSJnp07UXgPz8BWvO/dqCFsLIGOT8at
amoVv3h7zESHw5BUnX3A3l7qLjTfawk9q62KQnG53KSlwnPxSt4ZFnIlO5hq0W9j
oK3OwoY7nYOnHLGbfCSGBJbyXkxDq6HKlXTHxuuev4DmRU6C2Ck9xuwH0Jbfk8bW
ZcRiIuuh8uEpYa63aTU8yFAiWXp4UfB7dJXLIlb5kvT8dipbroaNM4r74Fs6Pgl1
lj0gDlA08Q3bAVg0oqgpxA==
`protect END_PROTECTED
