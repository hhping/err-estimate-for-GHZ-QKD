`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63ignNsXtWTGnKr4cUnIcGHV4enHFYxY3fNiN49ByXBqqJxlkIF9o1+7buOwIGce
u3VgAmiI8hsxBiTTtV+BBUF5da/OfJTlOTXWrhvrUtQHnEpxuSQvnjlCMgm2vKq0
M/+Pnczwh018Wc0p85RY2D5pJFfYDxYozcM23llrpRzk642tIJqy22VM+/HD6IPz
uHsvTp6I4sUfEGEaEa4sv4JY6aa+/X8wc9mrONVc8P/TRRTPovXJV6IQBJZpn7Uk
Rjl6ZkQYEw8PSZSKl4RYfJ8HQmqoxPJvLz/055c5P6qLihgs2Of8DZwkS9q5aQhC
nlvnE4CZw3T80qrufAbr7Cr1tFOZjzDqbH/kEypg2p2tAMe6AK2INEzMEXLJNWUX
W/PECOLZwWcY7dnRVsrn1dj6JZWY5u2E2vUoLXhSlr/R8rALK5mms60A7NDu7sJ7
+W81IhAWjg95h2u4yRof4QhRjvEJxqgn1Ic/+pEPDblIoBg/5byZJDLxweoh9lui
vd4agRlEjW9FCkZfsxmvf6YC4EIDwXILvuEmXYBEEVb6/k3wfgTJHbNqPVxI2+DJ
Yhogjwcq709wbSvBH9/U0+TzVwm9n23RU/OZJjEIETBB0gFZrHi/3AC7LHkljbdY
aPk0XY8XQKSfNYWBLS2avd4YROVPXsxzmhRuaRwmWxE0oW9ud4gta4PfEdrJ1usJ
MsVU0QQdcEsuxztrUXEMeLT3e32cveXR5yzx/WhW0AQ6/rq+rVkHwBAcALh9vbQ2
H2HhW0CeAvNMzVj/AY6k3QvfV8blo9t1+Gx3BFy7hHxnBj4Ob04strAKhMDTdl+G
8bIhOPQg891KZomy2va8oTbXlOl4AHJMOUv7trTBhqWyJLBE9BxHnvs/0cYQCHh+
EYgx8SfV1d1LOIIu22Gl2wv51iCNDf1SXTPU/KIwaeI21gI4++vgJqiTLiwPnXqW
LGJnNSiPyiafhhO8ZlbHnCRz592kC1j+3DrylBd9K0Ba/FHT46OC2XtvwjMJQKI7
3l5+02BNIzKW+654cu94CDmwv9lR47Am1Fm9/diXgtDibqUn+n1jtWBZe0vhj8s3
RhB2bFmyoo8jtRurgani6NB6pAER9xehFOpKs7+IIip3n1kY0fOuy3arg9ovVIfn
1OYYuQGazgaNN5kziVZyYVSFG47ZlJeoOQScpgt16QvI3JLYzYTIOvbIpK9YYAts
lEjBrkGdQsdF4QslcRje5a+7Ev41aIs4wiqz7qjkrlDXgxD3R7WmoDnEATAF/UMI
lYiGrC+haAUXi7zywNgFGf9BmZ4m80DwPcGpCxhgHE0ksdHp5FqzkRhxALZDgNjq
DXYqNoIGkTYs0BIWTydDUgAlyddINwWJzwR+Ty5S348DFvJRrkf0KS2FyLDmGxAP
r31UY3zVh+bPaxhnU7yuyrp/0dw7fIvfDcz5PebaoRmttTcY8a5GIxUAl9OjISgO
2fqtomU5VWnyVBaBSwp8OFvgx1/HML+G0MA4VMETxlfrYEbdK6KpkmhrOiDE+mSh
Q+RL6l+dwALtuRvufekF9zyFhfZvsyUJj0DLdIK+gJN5vGs3qdQyfUFNhNSaeY5l
Ve/uPaOjjJLKWbGAbHRQsz9ieTm4se5tOErjrvK93o9xGdSMLPB/gqMNYHc67uJm
LfKJ3asl6uV4NA+kYb6Gdub4qhOkgaPHr39KqObiJcn0aF0vhG+tD2On2/3hZkWc
07tRspLQpxJcFsYX5TwF4mPUwqhHvTCN8wCshNd/DCv8d3fx8oEiDsCzoUvghvlQ
fWgP5MPId4b/TmISNDNTWhDGW4Z79etLNg6m513H9Dwisw7qE6acRVcfSh3Og3NX
+lS8JoLcm1HWtT5YFmm1lZK6E0MJ4mwG7nhVyKoBGXXfCLbSj2K0HKfX45sHyNRS
xNWONBHjmSjiw/DRpt/o84/9dpz4jKUJILo7xEjv+9U8NGiyzsaDDYnkFHa8KM4V
FbXWjIz50J/w0+fNL8ZqOwfBTyQdSSe67M6yZxaofrhK6Y2daFKB6rivVuwjQ29b
7pTsBkRy50GYVq1BEeK/uYkS+2EuO326gXopc8RFI9s+HJrfRM2HRn5VVLeROZ6o
iUhzHy4I74JxNsy7Hjb7BwCku520r2xJNIuBcgsWQMzsCpUeFk5Xw3Y2cOUcOddb
dqeExECSzedpPMqXFE651Zol5B614vCnSXxF+iXTvYS1nyrA459EslBLUskprLto
92QWV+f/KQwxBBOHd7IQC+m/rV+PPSLLlCSVz3gWoIaVvG65o5o+oxT3/VzZRLFX
ew8UUr3qFawoVSXQXtiMkbNKzFW98DyoEAfkwVBgCg5aB9aHTPDKgFHI4olY+3YQ
o8pfOmexNDMP9iKv6wEdQLHocMH14G3F5sDPnpiOHh4AZ7ID2jBvSWHWmhuTRzhH
c8c9Lxwy0uf9RtpFDGb9CkjZwmDq0k73L8lWYjQr4LO6QnXoNjiffhKMgQFDnIFc
2k8UUODegZr/BhxIKkj3ae4hlEU9TDg0i0kQf+iCzDPwUroATMdvizyi49LFk7gu
2PBWl3In+0pqB2V1RARgXoqrsZrJzxuXmYqRhMOllORFr8yZZmWHymlZ4V3dKdn6
75xnst7rHEQZnw72/hpqMzUl4sWlhzal6F+7Jcl9zt6+4jxjpF0Ec7gWTZAvhnrg
z0W+ReMMnzmKe5pOiEEnu3Ck64+3/e3YlIFfX8mocSlISiYfdo8bUUuHLAWBDzmo
uXwz8r/TFJQ4qKvAvCjpEwbbhihKCFwvj3Akanq5nV7eX+a+Fz2OUTe0BHo4qoXk
VM+vSJC6WIHU1r3L3ZAlPocZQtj87dvBwfwnhU12odF0IpdPON5LzFdVd+54Y6t6
2YGdufCBveFVKyQNZO6YxCc+KqTveb99y0cXsHTebMAlSjAoIUWrZ4mD4pzhbAM1
OUYQb9+rLzVbWRGkYg9XJ7y+30ntgh38OCnHZ0OrMKv2YZplFouQZ7m6QZfoqKuT
otiSoZidJSM6V55EJuFl+Q02wY/FYWrlpjAToMMjDbQW4oiMww64RrEBcslJcJVx
TBHjf8ysfvzgEY1upenuDUSG82gxwq2oYpLs1YU5TEfADW1wxNgqyc332Tdxa8la
Ysq/kS1hOHAXFcFsINNdTiHIHLyQ3ZmsVP4au2FovSw8l9P0uVgfxBZz+bfc8443
e/pmGND7IidGjmV+PVibl+Xw0Kxqgbyy2nY3Foces0If9pGpyyZfuuBABYFwaJe9
H2pL4fdg3YxzMw1dyUGqM4MLrtwV8WhQUG5SI8uqy9k4p112QCsH/pefrWy4yggy
QUVTDsdJpUYTCnesoSAiaRWAXMUWjKaXVKjc1JMx33lvuc6orPhi9Dp7kWTKoIbA
1R8ef+6riYMN6nBHOSmkc7flSIXlgpq+XvogTP/kD5TiW7MRfyzL5r9F4lktRlQK
CDTUyE8m206ARSim5Zs6DGSejtRBKnkdjdQw3UOVHoeG33O1L1Zx4fWEJto5lpq5
ekCoarBPJNAgxXrfRzJQeGpyQb+zqyrD+arabT3/s+oG3Nj/wsQReOmhJdCzA4F5
HROs7Z3uVG/796UVtgISjsM5HHoH21ikJfpY6ncFvvqqSFDalcqkEs/JNeNbOJZ2
cb+Ax3dIxeY4lmb8xebI3fG6IjJRWhb4N+1SB42+z3D1y5fBSS5VwwdfB9ADyavO
XSMrRTDhLU4M//mYD8SooGEVmn0gA6eHYE3ncbLXuiN+uhcxQbV3kz6bWqTlq61p
WQg20uiYbuzbSycou6jh6djrP+FSYErVEYJbZufZosuaIC3qJcABK0oXgQyx0UxH
q1fu3mhpFYQ/nv5qL4/MbW2g6a7E4ZRH86nn+nDMx+vRNUpIuZe3No/f1glI3Sfr
Ib9yGcn9CsAVHWe0VrtJwmTF50C7lL5H1tVA+ekcsSS4gnbRT/wtEP4ecJlBSkWa
l9RF7+IM1RLFDGD8dbrmZX9eimWEBT2LP5K/WBYhUJvLr7moetnK+biRSNHJy0ps
s8yYoY77YAlSL5Ya8X47NyuJDEnQgDHouOdoxYmDifvwlw+xaBTddJ4+/BBHeE/b
OyQEEgrU3RoK9UmtHrOjoekiuhj1xK395sDPpMczDwj+K6YWlCKjPmS1L1Y/QGvi
b9fgIfnLntyCLlDY8UxWqRD47IakJ5zkuh26JCvajoK2D4JShG3KYunr17ixmHuQ
KJrt0WOaIYZt1VslVcoyZD+UBZjjCk2pdZWNNDMYUk4slzJ3JP19ftASsfPmovth
SnK7UenW8HSmQLeF+5DsVEHXzIwBzaKHMPrZDCAi5+njmIOoECjXjJiSe45KTdUa
6Y5ytUvfQtZUOr/5XIRLojCCkiKpsZvqCYBWfxWs/npSodivT2zfasYy6ZHPyENu
8E9nvNIiHXDkNNx8BFLeoOHqWjUqttBylHidrchi495O2Z7iV3WEKW2V+IfxdamM
u3RLIZSMv7dGh6tB6aZGSJrOKw67MJTDI+lenpBSUXwzLKt0f/TpiBRX9DyQvzcc
+X4UWhzW/HSZl/liM2ruahMQ0DrZ4fPMSakTBcTAQtlUo6Kw8MVwbN9JOs2y7zRF
yD+FkxLccBfaKhrBs023ahBg/HOlyWEaJVgj8LV5NL2c34m+4/gRSNGtWIwImD6o
kpPhz0KFs9WN0R723pOorqnkKqoCCQ03sR2THkGZv5suPquYIYxhrlJs02RjvgLX
2Q03j7U9qO+uTFrgFc6LTD9RI22dXfkcvVzKHbiylOg1yxqlNLfcNUwqwWZvUEBZ
qTAbjihUTpnM0IIj53T5Ww8BjU0H4ygsI/DK5Jk3PgFgLBd9ZfJWYHGwlRIsPoz9
LxlNfJc/ksVYKk208XREhB8vH7y6N/EvRGff2i/D2ZqChISrYiI8mN6ygX5L4zST
ft4OsGGPw+mffyyA7nFtx2hQCCfjoIcnmyQSxKlkGJveayqHntK3fgk7RqtE4wR4
3OVlcgZxtgdJh8VFAAP5iYcVsH3Iq8upIffRCaw3Vt2Kn1NjgNKZvMkCoYOPPyjL
OERIhjUTc2L5T/Zt0GW4XUYvxBRmTmlgd0prre88L+A1XAvd4SuGmLXM+VvzwOOc
8ReLZH76O9LXxvXZ17CX1463s8ecnT2BumGhCD/gFwKfcGg5dEFSiOGnLh09q8MK
Yhps0u3C5sOV1sg5e9VPtU4oSUGUy/mIF1a868eGqFK6yoGS/d5V9rxBcIQG325D
+rfSO2jQOrKd6Mbmkd6tea6zn8krJF9/R+Z0pre/1c+B9vkAreRXCNBIYQRQ7w3h
iSD/zSKA4A5h2kYgtF6c+Tx71zxA38WfqhYcKMk8IseOgjb5YN+0Efeaj8ntU6TK
jxqgSOHT0Jjc5rjbQIBd6nvkWCdqC0pol7iOnfwmm4tznf/o2jUyOkbdRanBC5/v
e6XDlipRagqXdelZfeGottqnMNkVetvpHwEavf/bfIEbIIutUQB0GWGUj/Q/Z9ON
DzPcwpHDZzoNSbkYsG1Czy6j/XxbnIEQlD+1CHH0IRCASAzjSEQBZF8TCw1XwHBf
cplAsJP6YuXeIuXxA1NIdwGb14HCDzn0n/AjtvlVs80ZUg2Z+wX0u+xXDnv4mUZr
3m3RC9uu3VZ8WSuzkTcpI9zVV+H8CwGxShdfHGPAO4PqUjrNn2qxL5Yu+kYJfmrb
QUdv7GMsfnV35udNjgJrsV/ubKJHz5lTpnuMwboKfz0YnC00eyUDdN9qtT96t5kW
7GauHJ+EGXz+vsCI3Al2tYqa7q0UnpFHHsm3+eAUez+4DxIE72BJEu7RuB1OFViB
1xBtCKPmmCzaqEcuZZ8ztgkGcbqXkcT2oYLj6N65SQNr6PuIOepToOl19gAfsnYy
0FA7kzuGbPWG24xJYvYZA9YUg9/+jisJtn3dUH3Rrdb3qaL/gh1VNntfsnBn2VxH
6JpO9dGai+UZBQOZ3+byhi/k9o7fzpmEpMfCdLhKvotox6/t54vnOpjd0nV/Satq
rtS1MSlD6B5XpTLytUvWB4dAS2Kk2pbLFL7qEHXwRAFgM2LBO5FUI0fQpOrKuN2R
cbGhFxXxkTTyOo312PZtCsRIbIdmYOGkvdIELbbWAhwb2vMIqPWOnDA7T3M4cBxx
pcGMIOdPlE9lhMt7IiJdELsQ05i3FNERUmDmjeO0QqVpqAXh2YMMoR3GvDNAKHR6
QfnYbXvC8qZw7mmUC7WS8Xwf0TBBdB2Eh7Lfi5dKS2Ghay4xiix8DP0E9j+F+UAP
3e1OV+J2flIdFd+Qyjvr4RivrP/S9MIVjd17LA3Z/AgktrVIE51s1KD4v+RxFHHb
AaFPvbrgdXRdu5Kr8K7TElzk27wVgqTDTzjLMkcZT0A5OUuVkrYFgl29vRFRUcjo
50fn6LivimRgv5pOdOFsMcMcntCTMn8CnH2G+kKZu9ybPPyJnmUM+topqRqA48qs
d9HvxiRbyL2OA8rSB8tvzvuBiqZwnAIr2kOTHWIyMV9HSasaaE54R4rnc1h1/Xl5
KLecbBCHs2GJ/5mSqGcSijokgrChyZn9fZA10Qj6eUqqAQjXdo8Bvoh9Im7rC/xK
V5RG/pH1xR47sl8PTrLXlK00i+b4Ds+bGK9JNN1BrLVoJuso3G8eolJ1Ex6heN+q
DzZRIlI3ZnRpxjp8079ErwdIKWGuE/+7g1aJSPOj9DZRf/ltFKuPbpkCTfeH6jLD
g5pO33zwnXCgQFSiiFQXTjjSMKH9DPRdUsNRfWn5sRn1aj5EjYaCosCFaixJDhED
Dpm9nRjjdKYRNHAprs5Aumb4eAG552KoXZlknNnfyL96yh8g5eGJDIWkvnYq+R5v
w76dHUZDdOyonns0K/zT4ERu7hIIR44g0pB8d151WxQha4NI++HnlDEHRAVTTkk8
7kp8yTVH3NAcUAOUZ7bCMp8dwT4WZduKQ2M4Car1r9J1ETE+32nB0DOo+rbldNYc
ojueK9/If+xORhvSv1MyymM2vQZJjRRVcLAIFghboFOEbY3pq68QunmT6ZAS/RTV
MAQI9F5Bk9gj9UB4bPqyoZ5sXAIOxleIieP8oNWijSGPwTDBHTAMOgl7LZ4izyC1
YdIa5kSTo+STSBNnt83fQ0+D7BowMXrN/Y75vTQXwreEvNfheIHMUwsdo1l7Zith
TqKPPyoUW9lSM9rza2yQ5Rw1z8dm2I3qnsvWzMLqgdVb4jc9vkut4jY7aT4H6hcm
YqViIqUUfNzuModrLpMeZSwnNTanyuhQA7phi8ZyfWzD1YGHgyI04abmfr8Q6OOd
l8o8e7BsRPhYP+X9nH4nH+xH4J8QVFmhVjU2gULWkMoLbkKNjqnt+o8y1o+0PdJy
iR+yansNcyYpsJA6jkKNBnLMYbeLaK8K9kEOBAmhKlj/A9jAIALf2ZzNzd5I7Tk5
JyP9S+b25BDd1jrkjoElOIp8r3W2tCyXcx9Yc7PreY9Q0KftQ5P70T0sk0o7clvs
jUnstmwrPNd7HLATpuHRL98dA9Yc3getBBxbPY22XKlpLubBSLSVTKkYNMUsuo1g
C/LoQaHJShpYvu/tecGZPB3Jotj8EQhv4R6PTDIKNaMJS1aQa2/gE2YtIblFFi+u
/ED4PiVDiAaIZzpiNrZw6vOsui5gDAbBl5+s79pyXADotZgAX1ODw/2rtbAvUE2F
aL7lLLHgpSOWoQWf0FsEj45OPZ48bXnqfENpf0RpsSao8qW0ce1vwzIluSaBMi/S
JgCMftUI/5M8FW5MSnlCt2A1u5elbgYjplXXqcZJEDt8FCQS4lVh9Qgn0IFA6ODu
BaU+MBnd7iltEyq7bdJn2imWiiMhVMTz+By+vxvvDFC5wBsz6yftKAVRqq8SnnVb
W7NbW3WmddMxCq8+0nbUXO5yc5j/1DZ2fBo+mIalRKxcjqLOXfo+RWiJqeYYGpKk
4SY7UY+CwdE4sMLjvdTUIo6R8urV0X4pJq/Oo3G1r7QI6v0mZ4cQel5j8XbH7eWO
MegIuCOpBI8LuplT5ylPpWjAdqMRmQ1dIMtKweWc/BCnPea7Ub++I4+ufltesaK9
NUYrqgcoNAhfY0CKGxmT3zGH1BgJ9VLwYpwSd4ig1S1jfdbMUrbI/V5CwhvN6aF5
oG1CpGjvv6VpYERxg3buwONb9kMxxrIi7JU/FHsV/nGF2y2BxEcq9pFbhp1FHFVk
0tNWrMtSO5wEiapVXt1GxsXYZJqayZoG1LDTLNo9UE+8JA6rFHXbz6XYYWGjLe4c
rB0PW3ZAYSG1jpTx8a1YhFicwkpw6+h23X2GlNgNzyDtszTwMpRS6w/sVhwsoVa8
Bd34fNfHkuiJKf15TrnW+mjPNb9Ubz5CH+2AQ0Ryr7FGhag1J4xwwRJp2trwx9Rl
GeqfMW3khIiSDTz1sSItFGwrDfJTa/0Vc/2RFHht3Lu5nGZ9TixaTTwCuL72HC+H
8B4P1JRMbJqJYiAVfczlt+Bdxrych9yMewIPqvCKWPmNkDZ1SpeTAkIzleADa2tM
VRzg4WfCXJhyPMWYjxg+1RKz2ib+LRFysVZYT/QY+aIRvIQD0OWWT2b4U3Bo0r1S
EWULlECAc15eOcDm/RIOjlfl7xruigss8VY03Sp4Q/39t8krryEEQeXzWpN1tHL5
+whtdwHsiYMM4+qav+KH5Sup1vl7JejFmdOngm2n9jnNBqrz7iJSDhDE4asUG7j8
26kZU/SsaZTGCVUXAzeBJkVdGxdlNl1qs/b7fIg87FSIhFzRD7CWldHLBixnIxLP
kwFgWqcxBllHiv1k6e9EvneG3MSWkWhGF5DaDEQ63eQ2cWhdltcTGEehKXt1S0NG
uJMJvX/jLMy2Y6GjnCJ3uwsEddEhcItYbQyCHf6zL5kdIUH4SUWny3teY+0/Weyq
jybMPFhEO6ihXW4JKu3/yxytuXa2itq0dphVdniT/XG3/HRzx2IDfByZslrbzclU
C+ke+8+KgegNWkr9wkquRiFkCTQHvRQeLvUArCMuNwMkELyluNMNohiz3/1oym9C
1c5lxuJQFTRRIfRU7+jPjTkIVHMOPlHze2+Dsd+5WtCnMsWEdcGfS1d8td6mPuW2
B6O8EXCLQJnlejI/ycjXu3DvVudGdGpVzAn7l9GYCbd7anwj/9HdjdUtBRGP06QX
4XBThxTIX+lr0yVIOmTPE2qDkyck9/6KwmWTnlo3TTSySkhQo1pcscZ90PEWZyVc
6vIXxwvqv7JVRr3VPpFhTzqXz/gZPIzsYKIATBn3Eu5k/4E1A3avutJaUEQLRtU3
/nBz9k42NP1QEjIHQc0teihltmN/p2E1txdX3JfyqtJwssWwa+E9PuPby5k0DBxw
YC2tWJkItaYakL7Gl9C0LgGRr27YkXMkSl3cjeCLx8vBfUL/6JGlGPBVETwcezvE
RABOq6VR4YMQhrhMkItFZFVY3EUjvx3rJ1Xro+EThERufTowzwb3CtkwOvXKY6MR
CjeF/SX4UV2BKwqZVeNBGrwF/lLNYMgZyDz1XSTk8uLRFECJaQ2xHiIOsxC6S/Yz
aI5wrKEG61c3BTt4hlFobwNKoXD2YnzfaD+iXdMW1pmr9pQHqNXPZXfGiXnROOfc
Oevts3t55jJHlYRVLmJqCoLGwsaofqbfWn4pALcPbMIWrF9NuGtL88mXHXmrbzqn
gcYK/vdozh9EV7/JDEgjazMVv4Oz8aqvlt+22wZgM3nZrYle3TpYfFrNgx8aYAp2
/0WGCV/KXBojSgFfLqWxfy4Wcn0FEi5SNEMzANckzlcJEc2PbJck/buf40OdMOGL
wBNyGeq9h0zjT3IA5aidJTA2KAyQmgOrtRJHHA1Bs9cOGtxqRfuiiUji+1t4a7x8
z54hHcLyeDpH4RMcBFnsE3m7AX5FKroOW4umOwkINJsNdiPFKgG9MhOceETAQJAJ
0X+RoLDm6WwGF/cDUOaPU7Tn5m/yEfPb2CbWDeSMnrXpUsJYMZ0d3R1cRXhuHwWJ
uSsKKGliMxtQbhI8TRhg/sRW6qIYWaEESXSeBs5lcyx2pc1M4TmQDgEBZLRTNYJn
wI240tLacoaDWf/LMpzFQmdFLlZ1ROMlKkMajr9cYXDryePS2AmbeuMcb6hsr6Cy
pB4/m0FVFWK8gxzOQ7mgUOJ56M4P5fXDuC7pU4cTtf2AmzHioYVGLGteICN9tHOB
I7cb9TQF75kkVCDdFzsn+wIi4z3gkZiaHhY9jmNsb3JiBwHchMOjG9Tirh+I+K4e
s9k9OPvoEDvJE9NEheTbqK+lekPrZ0DyOqWGl2rpOg5iUgQtztk1GMO+JB41A8DB
6orYs2owqSwGjC+Z7oe2SXYzOC97D3dtTqJYJIu5YLOs3Pgd8kF9ENKOIwbuXba3
ga952yireHtS/LbaRv7M5QtOedbrIY6JN3nQ9ki2rxWQXVPy48t6YzIq/F3cBUul
PRCtPEWRvpuN7u7B0tYtRb5QTgQ53aGfhNWS5PKYA7rSxw0AeG7iGoMx1e/T/zqC
96PsnyeHzJdYSO0K1G4RMAqONy0YgNShyso+szLwg0gh+1GwS4TmjXKz+6+r2YId
3E692oJcy5zRpNJmQtZpj+UNg8wvEHoTQuFgQPugadAiu+XH9dd+veOu8l0U+IkG
/NJ0wEgDede4u7HjuLLddPSghN3EZb+UzhFuuHwe4LMKj1dGkSFJBG0rMY8SEDET
aTlwIL2ksbO8Y3dC/EvhZYnYPvLE8IVwwWtqJwfmsneKdNPdLhoeBdIDfdtsk0pt
v1xpQcAVrbPiU2VO9U3d2an62WCqs6rsrfjPw7ysfuj0xWKd7nL7JZg3EUtESzIv
GFGECXVZtmzjOyn1w82V36xwPlndfLyJC/kGKtR+GfI1z/H9jn+vt7YDX9o7g0Ya
yEBDEx7byZyHfObQaEUlKGdSXyold52T4lHB/BUqEVQWnPeEAgJb5Uqbar+zbMNf
NHyTu8Nax4/f7ZjEl+sA29nbM/xZl6GYlzKnQSJGRY4HwhsYX7/bm7elIP7Ya6R+
OkVFgGihjERMuSYvKYRdiakq9UO9qwcqL+cfxvpazA4w1HF+zhPbkQGyQpaoCVfz
jxVO4i1ST7RUSmKVaQ2qcd6EqY2lVNj9lKSPIOaKqDa9wrGMPrJQs1QpAD8W6Djy
rjpThtI9dHN/LPPGaLgK/nCr+GPTEW2khnKIyiuES4uyDojn8zpD0/eAg0hLcxJv
SQz2HOT10w2uM4hOUMr/XcrKNq8atyf0lFTlEk5eG9MeV3bg0kHgt97xB2YAcGX+
O/8chbqsdbCrp1epZMQ+Dwg6jP28AY31zIVtFU0sxInug7mUXktLTb/1FqMjhy86
E0upsCPhQn3CM9TWRjOby8+gsqW3vdxIUr80yERoC++p7qrthP+6qG1tgvkK04nN
DqTekhveK6hdTEGrT8LiCwAZLq2+srkO86CbQiTaH2WuA3IOFC9VxH+Y5O3pPM0U
Y0fQTWAiFiwZ8A6R/+9r5+gyUTbB+dOLK+Rb3i7ZdL7UsZcfmL3c4nfua6E79rlr
DxZ8BoS48io2ohZFNELU4KyiJnIuhuuGW3MV3NV3Typy+oexjCBNdnXt0s2Royk3
oDNuPSTZj38FgmkAiCYAqsNVGdPiBdl0HP31NszlpfHoFJQKcUmHaN4cIU2gPpUJ
zpawTRB1lSdlciKdRYoEE5FynNhZgfID2XNT02aUpLJHgrA0ZPuKRVXm+dQc5pOU
oL0IRsnBVweN31PBLbgHXzIuN8r4KU5+uIaTMpbWMVRunsrHIoR+SU5VVKS+7glz
kI8wIqEX92AhKF9AgYvtvx7/y6Onr9CBA1noOfS8do4hCz0hfDgauqOjiFjI1GUE
/63for/Bz5irSEvTqbXQqJMuHTlWhxFzLkdha7j/T/Vok8pnNw1fq9ty/DliHLhB
0hz2SHrtW+CAemK3EJLOObUR9DiyCfiIwAxLze9F1Y219B1rSfRkEuNKDa2qcrTZ
x8Wop3bobRIDNj/z4ht5zd9g1n/miFmdJdv4oEOyGlSpncglS2GDLih6ClyMFwEX
74PkkikOTb7lS+hJnXGlMhhpvB+IsrYaUh+dPo4A97G2lzMeEKl0p/ETW3Jb2K3H
PrGmyPZkgbgx2INPMxGn4mO2dyYT8+G9NnPCUS5jGUB92ChwDbUN4puYIUOY31v/
ucimlrvxOPHc3xxo3vX/uRxrCG7Hq7OFDhEeEMqG9i/uzRoXdTOnsaD3I2I8ybyT
Bg0XD+2qkaIWFhntB6ulzRNjcF6nRneBF6PS0bkh+5hxKpptZ4A4fdoxsLAVSUDw
rElhBOFpB9qlGQVXIAnVm9kwD3jwR6llpMzxdfRbSmVgMTSnztyNPG8RjIMVIIoQ
czNXxB+gg/dL/h65dFbpZdFOkj7+sVNjGYkZr/SXXBtHhInIsdxueyH7sEqgYx+7
e6cBkk53G7ZZddkhHOFu1q+5tPBpTaRI5XL7nTdF6+dXC8Q+uK3rCnwoxiPOe3kX
3FA8omWryNpAE7gVFSN5EPUbD4PhPoykJKP0idVw3XAm7Au/gEeMSAtuPacrrVFG
RXZSoZvkSb8PJWQOJtdjM7Z3JloPVqIQK0zojtbCV7y6/V2+M2JtDbZyTh6zyMnn
JVOQv03u64wrhOn/oLfgrKforYs91p3gvBBxRI7mg1rdj0W+yKSmdxPzb3GGMq7G
8tx4oTAZQsiWezkTTNNqS7kt1zX8U7gvQG0H0nA1/Mx/RBKMOiZUSyGDnSpFc6HV
WaTgGpSs0lIF8oUjPF6gUZ30ybDSppeLKp9+kZ6jxEcIG2JM1ejJLGp0kaPn2+WF
2a9QmdB567p3KrK1tjaz2Sx/DEyMgfn8PyEQdK1xHGQXuVshx8gGgRWJJ8vtawWe
LoP1gyTkzoyfqgZr881JsYyNfADF3rqHqd2Qf9n49jmncXbIemCw1i1r+9JuT2/G
d1IlViDOAJoODboP3dKuNEaz0a7PuKjPyn8q6eaJ9r10FwVWjVtQ1fHP0oDnZqMk
od5VPLb3NNmafFj/WgtZvCuGYNf47GjviC7oEZH9z4VEf2jqjTBRwmP6nHpWW9kD
eYwygu13dPYs2DfK0M3/pt3IRfZLteEMmyOkN5FqkHJfJT5GHl8gg3bfsP7PxWAa
rlCgqazxkF6qBBYkKrb3bRPfP+c2ThzOjQIZKJdbsSlUW120y/LKvf/Qw+VEzAC8
3is1BOvC+N822Kz1BszYhvnv07PQ2pco+EWhLoV6dCMUYMhpWJwwl10n6s2unmo6
pHX3P1wy/obzFdbEQ6CKdZX1jCPoI77Z0rgnB9tJHJ8nedfmEae7HD2AcgoEXoqf
Yib/yDWu5sOUuWhIik0Ul3l0AuYMwmsZNpW63uJR17PxuCd6Yparx6Nz8utCHs8i
/EZMa9NWkArI3ywTHrRBHWl/epIpqaMR5zFJE2yR0gB5N6qm/4quzBOR0tYvQA29
fQ7x3DmWTbRfmTWRmPGBLpkD/ccs83sKcnTkWdYd7cmw78s4vOYRrpottnQ4m601
lUZTlNxS3bNFFjwuyMI2GsYd305jVQWG6s4I/DAc4x0pefvp3wpZbzIVj5+b09Aq
NvLyF/aPl4O3hnIkWVgtnTKHW2qU97rugqST9hpGRWjeeXOfk5+TmbPDNcRSbjrt
JJngJ1GjbxZaTbUWOidGjRHChXQUzwIqwSzfnQi7heUre2W0pdKVi4W98wMvX4bP
YRoduEuChMoXO+LwvgYTCJDNSOQXzmVAgD0xNvRQPUKqd4fHtYiMIf8JyxSni4XH
eblOblUS48PK9eryDApyL2ZGMFrM7wKbnc9UcxJ1FSQ3mJjuCFJUBWGx95bTvcvP
8hbWMxkJIP3PGANf6l3ArDksp7NprTYTwZYRlD9Voryc4HwdEQaS4rQ0qh7rY4MG
eeMeaBqtR6EpIK/mjNQFaMIzGwLMB55oaLvLdt0j5rMnYmIAt+KfYVZe83CnLZOk
RIVUwAa5CPzXnzBXHekKOD8vwH+QWgeNc3bs7ek7DWAjM51aelk314oFwvcRDX1A
KUzFauGToIMjB9/pQL1FaAXyHPfOqouVR1IKtuFxcyQqpyC37zIwNMxIaNaJU6er
/emAfYywXrxUddlTrddo4PJfwhIPlWirjPW0nJb3dcDIvR7wjoucpqPrPw9hqEG5
Zf0fGQWePWYzdbfZWpWpq/HApmE6VPBUmXochCa+nDlh3U6HOPSx0EUTQ/MoSaYq
BH9gv8XG6uNy2otDztxd0StYhmaxNeDIzFw1mtctkCBuZP6oftoUO4V+S89lZPo4
wu9r6PHr/FOuDuRU0KgObma6ujyfWhoSoVWeNXnzFMhsI8mK8Z9K+MM3UfViyZCr
asGs42Riea/L0ng5qSJ8jf0mnezuirelBvoMVK4bMIdB+19oKO6IrL47HLQf+Taz
5KUNRN0A7ReR1wvUMQujj8/G0bfizFvArRMckzO//qcNHBlAIyc6j/HmBRbEjCPP
GpJIyRmIVJktLAfzU4JTgcTJZ7fUONwMmEjl5ygM6N0jWZILAl1DJ0bALFiENWlw
TxnhXZrGs52986lAPZKvivJ5C8gJZU4KBkD1OQKXBMj2Onhzyl3DQbIpShvn+0XM
90wI58Z0YOnXtlqzn0OXZwm0HtmMo9t9mk6jjyaHk4vYTL3tKDMXiHURg7+6xN+y
XUEpH+xFJrty2EwJBs1SOuKMcL1Sn40ETCvD9JpCVw6C4tb7HkMesii5v6OeLHp5
icPP0t5l+nFrS8ZXefkOfqaQxx7zVIAmztq0T2za9PQ4xPaHCJtvcgVpwHTviB76
1FbCXD7g/7smfBx3VUP35u+csjsCo3tUDUJ2XZGrivN0IOZVBYVn5EAqvwyH3Dl+
WAukntMnzU1YvuHll8radIMg1BOyCbI+MtF086x/HdYhoL2UX30z7MF1f0MGcJfs
logGA5hFrfwEpNcHYkYYhRjdeVf0GVhWL9EuhhH/QA6XmcJxEma1dky1QNQk2LFZ
nGrVCCGIUdsmrI/AWai2vb87Npb060nf0qsWbYhDEDx3g1pWQZCgpqkEvpMLi6vL
lrfvBqfjZIsqb/OXM8hmza0ZBGwR0EdnLs44gndBUqmP65cmcqrmBUyfFJ2QNvgF
11qsgbzAuqcYV6GB7MHT5G5ABam2znzAkDMY1snr+jeq/SdJ2sLGaexA0W4U+L7f
SfvabCZxcZJa/stRDlF7hjEG2omJDTdA4lISPKKUUn8R+I4qCgr3MONeP81cKjgs
U6ujpvVweZl0rW9chnjJ4FLw8gQXLAfh6aimH4KpkRJnlIutXoxb9NetfnBjodYz
QXsQ/SZPksMvzCrVXV5uEYgHu9zVBTpo6sPz2bs9IPdqhxAoJHDZ6ZzgmihR2gxc
nK/rucnpouh2WVIIhg/FXHl1cFAQ9DX+uMbcaXYfb9Ab+hCHhOuBzdIHbSu7SqCx
iUrYvMA4ne+vufcxaVnUX6Hcdl7AQUa0M6Ut7LumCLLPle0bwBT8KhJ7BSJ83Owq
SzcbtlZW9HswdTPkOITrM3xV45WRXq9NCqGOTUX2jwixrrj0UNkcBNChvBCMy/wh
1mm6xGJq+UEofDA4oP87kxvZjUw7Jd+83PtfjyRleTW9IVwEga4y4C+ih9y/RBMC
quNhj6XqDebm3CAllxjzB6YkY1k7yUG3XvaxB3u1ZJDlfbkVBnJHp6h62Ckuiq03
4BLyk73on7TSab0ngpQweI2y7eOkH2xZ1wRYmYHHVHt11sgMGEWgFpGCaneecSQm
7UzYBzsswNE8fJtmsQ67WzKx3uSQ9mo6zsFfVwWnw1Sx/I2lJKY1C/encNVlAqUt
OO370XstzWIloWU27MWlgvryDuqlhl+W6FCyfMCfk06fkLKZ3yYQ/4xKkGT+ZF73
QhoLHlDdHUWMYZghW8zPfhAKaM0Ocu2MbOiXl/i3uBg/4NLk4zFz8yU9Cb1Zyq69
KG6Cy++b3Dszj1o1hnXkuoKDyQvrsA5DEeXtdml/TZef47bLJ+33aurrtiwsq5+/
HlDrczawvv8ldtWPI4ABzKyJewWeWqUXS7GkYBvF1O3WJ6YPTdk3h95yVtcG0o8p
UF0vHK5fDLZnwP5KVLpPCvzXoG8VGEZFgCs8/Dy8t2d2QStxGHpWLcDrc5ICB2Ri
glt0Q2Da1WK2hdycAJtGaxfj2K15AvQ8B/sOz7KWrDJfne+hgWmgbgstEwDqGFkm
v/qfqijQS/1g4AdcIugO0N3ROSIIrZbR9hEagHz3oAFE10EbFqlRmRr26BpkrYsm
pr7hy2ZbiU236L9/CctRDkYC7oI56cS4qzkYqCGfVKwLa6X0wGaWVSw0RU7oNBCk
JzR8BdrX9IWQQpfs618JQYSBbB3f0AIoHxdzuG2DxBqGzLoNsBrWH6+xfh581dZD
e+Y6XI6+VtmUem8lSCXxD87i6WtyL/SNErrz/4vqvdqrWwvuMV31cwVMRzSkixR9
Wo63s0EAZVjJJ0LxzJL3ev8CNLzUeH3G8dXJBXP5B1pSpR3c7vFWPyGooQAvDXrW
wG1VRp1WBODAPuZ6MKSTG6iGunsBkecUHMjM/XDLTbbYbdGo4/zyLKgaGmgSSyho
4W6WTiz+spruYezF7JPRDRYGQ2q3iLK9a6/umctKfHtrd1EVbTPHShRUSQ+5+Vb6
ZTtRbzOtJ7UsznVA+5WKty0Qbq/tNnUuJhwIBrHXG4BYViiAURgC0MpkCIEgX/LI
uaMcPxvKvYh/ZEo6CZNHbQoLUqW48ThtF/xt+I+D5/mNE1L1uyL8t4nA6h6pndV6
4LfbiKS6ryzT7GtUjtes052MSqrhZcMazfF8xDo6btERZwKnollF1Q1v8rAdjP0s
CjB5ki/fsyDrgu7yef1kQtYYHjNhRSUQExW66N/0oJ3EOH/rAox5uPsX3mR45VR0
FVJjiMcdrGnTtCSr9GuX/a5TpGL5U9jYqa5RpjmjatKNZtbrwLQuy6bAnoae7ucg
3C/bruwI7Bpv4MvZgN1HOQAhFEni7ut4+88UuLt8mtcie0+pc0f+OV/tQwzwqL4o
YiKt1n3UEtzZvvpYmwlASWj/R0QokR+bu2xYeG65hrCjldP4WJZ9mgS1c9CUCtar
ez37o/6RCczQG4zsB5JJ3wcflazBIb7qbRYX/ofgZ9lii/dSqAQHow7ncvtwkGix
oGmD+BTXnUeoIYAAHvxS5akX6JI/ixsI0Osn/xzljG9kv1rMnAJmbtqC68+j6zvi
RlKaKYlG09lY/xMqc43PW6hf5h8eqmbZKKjp2txXCqIm/Lujyf2017g7Bm2ak/Xk
jTytXfSZ0tW7+g22QdGX55PUxZfevBWszI/uNgzNhhC9a/M3+oDRwtYx6Pam8GMT
PIOT0dQECo+uWZ0Nw41+RltDKNL/tl91EGD4QgY7QVEa58VIhtpFft7IFCXaMJP+
eN+OjFRAVvUJtAFYWKaz/s+plVrXXKSpJogqYBTxnF/iK474kW5TlmpWeiHjzi5R
yYwtbqZh18c4dBt6CHWyqfU09nUAe4Of/CscqPgKceBpbGhPFZJGRa1pRCWoODXN
djxlyRI7F3ih80/3OyvbAz3sb78wFJkxb+B8tlWf/OtgSfqBB6DDKU5lmreGqtSF
iCKLVsWP/yqXqMudh428eObTyuHj/9EEVljAsH94k89XgqMOmV4tZrPRRd8q+VZM
H5ZSI+WrBxsWypK2NUDOo80HFdJRWzV2rNr/KdotNLt+FPZVtOWnbJQcmm0cGKXg
b4E9kC0BCTtud4s00whZlMRCWuK7EoYpBI/K7IEzYvjHnVr0LugbxHEud+fZSQxK
ywKXW4hDtBO8lUR/wIatphgGDN1n/SiFhDSqMb1FMcuZaIaKg2MzLO0xrm9PBIJi
aVMvPcO093V9afp9WOfW0+Qwxdo94aq3mxnwSXl9YfeujZq5MeuX/1CD2gP2cevl
qy3d8005XZiL0rqR6bhS3k9+Ez70yLRnCIjZXNQg8JN1uCqTpGZSzdnGnUm+1aQT
uHRgquh3TB+q+I0ehXopVUGIFBKImYLN39qgGtqIUsmi6Zuz9nREgJwSbLExzMN2
U8y4mIx+6zynmtkj1wpfJRLBcrv8LAcH3wRE/YbpT2M4wzqSBKl2mm8fyEbIA0cL
DB3YtxdsyKFDBDeQPEqgcVPZnWAG361cGvLdjxWkTxgCBlKPkCpcUvQsjUtJFGTB
1AY8/4pCrogD7LjO5gd/FXL+WVN+FwrP48Z8qRuaqng8Lsc0vLF1E2nFGpc5IfHe
4ejEmCjzlQQATWQwOcVZEU2gs5hy0CK8PXjt8rhap8EJtQh0TNIpIMpxX65wi33R
wd51ABTK+dbVFnvJok7fEvCwNx9hcdu7XfRdmm4DVdXXSDKh8C0y3rrckpwEA8Il
82vbsIqzv6rqEqgZQfC+13WkyQAISlesE4+jLmqrpAZ9f2nhZOvopj86FcOYIkGZ
jHGYbQjPqSa7qlVCjhwzsFENnv5urtZmFK1IPuRDRqn3PKT4YwIH0i8bb+20HiYF
CLnG3Gel/eGice5uR9qkptofeGlpQaspU4QK7ODt1hDd7N6eV/WCxLtyaxcyy9Nn
/BAxMg9o+tFOOvTtxvThD5nhaxIuE87DqcDTTiKw6RA/4if8kh1ewJpLcpuxPWxp
1KVXJOf4PIcyMQ7/5+t9ekCoYjt0QNcfnhtfWYFIAcnEZE9v1jDYC4zB0rbyTYWQ
yNCvdwYkeAScPXxKla7MejA5jHjikkQTzpxjZa61d+7qnPuZ0LyjWf0CDlWu37IN
W+t8kPeQQnUoyp4x9uUlRirQ3ZGqF30Mb5PjzO7ASLJ1W3TEAaCGe/mUAkXLP3dN
d3y4X0gbcfAn5vAoJl6qLWkiM6k28FqErilX+EXhrO3mSdeX94RE5qGgvdpspLdo
bkjD/zDOabECVAo6Fb5M6sljGNDfnumMhmwn8j+kdl2RCbWyEQNAusYXFpn9Rp1p
b7yJCVo+jRbN7WXZyhRaAHSt3EKzR/eki0uZ/G7Ab3E2HtsvaXGX6MBbBhFYVwTv
NOaSYjFWzHLDHzGEOiloPvJoMa+KhLtszxQG/1j58Qt0h8n7ZCOkP3PZRcfkes3U
+1Q0D1T/iLtPuFVo3MmxPO5cu9sXbweXqj4rAbvi7QeAHRnENDSEmmebye5XjMGG
9tIp1qt8dR0yNmmQCsznbFeAIzTASQgxh9rV7KRUpHZbMTbYRdN9A7MFiMOSBPvr
FeHOxa07CTeABt+VLJLWMLZJomZLj4H+uEvPnnDe8lqBE+m6QUZddagoef3+2z/F
aeO9IRcvghDaiikETDblNaUlprUJQISTYu7GcvLNBoHx+ESmOwLzEfJ6q0wK1ELX
URcM18gviGV6aWODJphwlLdTHg5lnt33v0dseqSSdgzIeOvHD63s+PQAw7TPnmaL
AI4R5YT7QIsxuuAwD6Y1FedY6cmKefY0nqXbNRCGZjM6Val+gNrvDjnt7UokQX5w
lvNPXI2jIhOKwhDfEE6Gq5SqoUjVfugrBZO8BdMwEAya1KjZPIRLX9L/pKF5BX4r
y9vftAQObKiAUOe6dNS4aPW5Yoo5IKEBDgygkVakstJ1EYuaQV21Y1ZRQ8RaJ2cN
7JkXTq9FBW8V0c7bsVr8y2+nGtYJdZyI6DMLCmtIltrT4mLvA9E9ZXOIDwGAdWVV
0vw2syVR1nv+MB00Zuplz9fiQT/bKMZwnxZXaZgDjltKE6pQW9Eu0buWTzvya/Oh
kABFD+8ibciPkujQkECut/1J0u4t31cWpcb5sTRc0oYZTLKxmj83IYjoL+eQmFtq
wzZ3FJCkagwSTZvpTQ3fIxcudWoKnENcrRbLN7iQZZIlYTb+T34GqE7kq4vzaqVi
7y8kaZ8MSo91Qqbi3ikTr8MXqkV1X+97GT6x4LS7gmdaVt0kFFu1fN4lpc2+xHy0
C5jGs8GNe51tEMZqpD5Q6NAvdCpujb79lGWwbt4NaEDifVH7P3BHYzVX7mhvqrSe
0MAPOZqIfCxflAgeVrPigTlOUolEANcgcLudM6RPowOTx70/2ufUunEZVDliD+T8
Pk3FxyDwEz32PBAiQ3ko5/LRmNWxSJYwl0nkZHffcmWEiEvTCwSByPopXf+3FWRC
AvcgEbuwotEdqBwzfXgfSOJa4yh/72MffYM3DG07WhYvyJlRiPQ7bKSS7VBJayk2
mcPP8oarcUvYstpUrEhG/vF860/7dafilMt+EDSqCLVYp9BA/NWVkn/qdbkL4VZk
hpje54f/HZCIJfU4jE9EvTp0Mi16kcv5kXIQsYy2CYQVOGerEAnygH9vQDy6uP4s
V0U7jqMBRnHayYdckOTZcG+H+wMGnd3+UzPhtAacJ/vcgOqopvoRq7OQjFN1Di56
EdWgQdQLKBEABksq4T/jI42Q1oegBcZj7lZzzGpxuc0noTqskwf+Ju+4VMCaj9Ya
DSeMk4eXOD59aDgoe4qpK2n2dX85j//c+0mmTbVQkt1DoOggK1mD20FWksNrKTgF
ouoK4Wy8wEnNEK1cvy/KhKJA6/EG3xdGmUE/N9GEKbN+yZzWlCbzWheR+7eJziSP
TMSyg6XFWVjmStPRuLGFLDMT4NvT5F30JbZw9v5L2ucIKWMB1tB0I6y9+K1qQTJ8
hp/ApwBvcT3Aakdkovm4c8IkRwO3PUoqE7e4nQpdXJVWN9W81Z6I0sR+udghaCMG
b1Pl3taTPRbZdjL78T4dKUBM0BX/6u3WF1wsGu7W1goSn4Dl5h6FaGZgCYS1NgNk
reMcYIgisicHgAVOzBH06F4gsJvDHxD8x4Y2jQMovG234On402J2wazpWQS1c5hR
j//8ajq7cJq28YykiahFiLu+f47hVhZC+ARH3R9sLBxJqF+bD91y21E/FJXQILxk
8omwdfX/pIqX8dnbQKaQMpMA80OxbMqHneG5z5e8vZ5n+222hk7G8xXp69Vhv5OJ
MvsYSSWiZh4fnnO7Rj6F3ap1CWA8B180Dsr9Nvxhx6qv2vyL1A4KjI247+CzieKw
RogWOaamyZZmUtVrAhlrUqDf/ePRYgsfC4/sIcbT0iUjir60hMhypfMQ2H7YZh4o
MbcYsVR9DDVCCBc4oyTZ8XyeUQiIWjWG11UPp4ufFAjfzNEuTw5I25OGm/uoQboX
Tr0UbzzIi5NCzS1603vFHg2jic1m/c8/7PtH6FXRKHBReCv1U1COxSNspX0GYF56
ZvwT/pfrmAnXd4gDcHXRsUQe5o9ofY9uheurf0ZPBcSNvyHbvflcngfPPOlBwAFQ
BFgTEiJTFM9hqnkkfcNt6fQ+RJ4aPHhpUdlWsS0LM3P5IfA3udENBifsa//W4fEy
YkTAcCJDl29spWbIMOWGNnBhtS0sOtabTV0chzW3uesrSHNme3IuRXQHifryGODJ
gtLBQHo93/V95B8Z+BI6mp7qSyecpEV8XoMM1Ee9eveLnM16DFl4O9fHfFf/zc2Z
T0J3bTsoxR+s6UeeKc4k/H/z550sTyhk+AYApViZvNzkC0kRsinPkpJMpwQldskf
l0MuC1cUUV91pNqW3Y1FY8PZwmTStF+AqrQR1dC/9Jar24+/4V9+DoOj04+LRv5u
NVXKcyODoBTQUd8syEl0dr/ToOU9aD+CZVbMZIYZA5nPX2NULuwI6iMycPQFAEFV
6ake72YHXvNeGkDm7zpM/2ltY88x+uQYuDviaWXkyQajAzWnTKPy2xdNys8f1rqS
pS8cuRxBNN95Ky9hUHfSbx6PWAw5CyrHpz8x0ElUAfneENS7ae54S22Co9AE3n7A
WS81Vc5YDTCCe6QTUizNxsJg165otBYh8sZpR1Sq7ZYUD1m7mciGYC5X8+Kc8BFx
p9woj/d0q14+3f1xmoLQtBExiDSrtl+0GTBRljRatk+c3MwDp7P6K7oMRcgEHduv
bGcELEzSWsNsvfRCerMJ+GxPbw+8z7lxTbL3PhcxT41AhIbI2jTrgtTWrTkgSwEh
is0Cwp5QhUpZgiwpnggqyffVibozCN2kYmkRGlm4ZDSqifwSjXjubJBoxrWLzCGb
ZtfqUUoEETKpowGK4K70/M7KNFpHWJ1EN8UNgoFQKNS0l+uXKmnD/fGiC+ql3OYL
5TYA5ZeMc9MQdyJtvaNabcBBTr4WXAOwLhCoP+GgTiRuubvEdIytNqruPBhwv8hd
wR6X92jad0MAz5m7a6JRhyQ9nwkbWD7myfEjgYddMYrf5I/GUcZCUxypnvaXBhFz
up/TzIzj45Z7aoa3mSn+9FpRO6x9h3CEtuR/YnP1e4dKzIF5dWIgig2zFABD9pRi
FKk/GiHUC0hy6Sdwg1KP0RHz+hIRZuE8tF5pSByeKlF/grootcrPYT5pGzimIzDD
HTfQ0TTrZA9me5PpA5jDVZ5PSEh8EoF8z9wUMBhuvirLcSaKffxJsirHuYR8CIrl
afecT4RobHRRKb4cGWBcBZf9PGa453icg2o+zCscJRM4BjgsZG2WWtwzXVSCWU3E
/p9S6Th4wVikVOEgYaYKST/XUaQ01EsqzKm4A+DNjtkQz4mRLouyEvhxhH3cXVit
MaYkXjC+kqs/0aijfArgRF99lj4g9mkAv/cIIAr5gSMU7mOq7xBx4XRn7zCynvAR
0Y9Fz2JbFb26/dMK4h0RZ8zjsdoDBlIVg1U0VNehc5aTXFke0SMIza+jUVIqL4FK
g9pzQQLllsXlW6wYoCZXUH6XZtOrErwa4ymlpdhylkgYimCANGm/fnveYquo443G
FXTZOKBYsQx26+W+vA8jQ3hsf+A9s1e8L8Lchu+I09m2fG59ghyLPguElGEafPdy
Q4tlAXpDucrJ6jB8tHp9CORjUTQ+DEgruqO9d74uJ+pS+jIHGWWmMJxQ4UgTb4Fk
d3TH6r4AHI4DLg2ehIpuPgr4p6QxnHrWyd6MWN3wSrxbaSbefcKggR/sBNQXeLC1
zoz6GTxyhJqYeQT1EJKtdQq8wk64u+n3bl0TN14Fal1JMfGGGOvJskvJnQ+WR2A6
0XwL4ZHGiK7T0Gy8pJk1B3WqeJOWaDA4iSh21oRw/ug7J9xHXTXwgJQYQ+FrbVH9
qq2Ehm9+NzQAUZO3NTMJ8DWeokJhiUgTWOLocqFvZOr9RE5IIYMjaUX9Z63b6Hxn
QFJJWzOL3CGNWjAWV67O9VJxvm32CIN/JNwhjKcSuKGPOS2C/2B7ZQTeLnq+Wxd6
P+Ajtd8ogA/q0qlC7MV3XqKiKC+R7pxBOJzEYWtlKUCNt4XoYWU6IZuI7oVh4HK6
UffsOjQ0h9qBAvNN5+wdqOt/Zz5yMvSxw7BxMQxxDURxnPo0YnqrWfANLWrjvYGL
vIIJoqeoBkheCbzcWS2W6AL3iRmZa+YvHhdQHL/Iu56Hi3KyHapFbhwpLArfIAe3
Xla9uYCUhbozn3o5kARBpbw1My+3e7iHLbrgEOmKHeTyJFBJHrYImt/0CkfqudLh
jNWpL0MEBKtXx3O4XlbjR7Nk7RQPUB6YLZbWIstwqxOFNKdGjr6ziblFf7ooYMED
KnGMhCtUhuqGK3uxlzJRofegL2jT2cn7i9TpcyCdWQr7pSKiBniS87CLJcjj28W+
N/dN9jgCat8+VCDIl6hXeTSSVn21sExy7+3+mtHS/I+l4gCGA4SYEi4WJSWZp+Wc
i5CPTHfWhwE2TZI68TP1JD9NGIZd6G97L189nkU2JTfTlK3h2B1iLoR6fUpb/Rb0
sg1hisEmb81QkkEQhHxHtAAeNNbF3BJATjivOzyn5kDRh5UrarFz8p3od/QJYy75
Zg21m59R55XoK6B2YC3JlCRWm4IMWsbFpn9kGpfFKRsPkjwCvmzWJM6nU+fFi+Cr
APAaMIvRVc1qJalJNhgcc8MWvCd6CLV5cQiEi1AitvI9QTad4Dj9+YfMav1Gf8Ty
BChO1OFmcGJ12UqBJtoNM23RFqH1a4CbdQnf2A6F452eGgSNzrwpun5oV8EbNBM+
Yhv8BDK8bhvv2RejSK2aY5qLTxRIeaCufJ6AE3yV6FWM85DVj0YOWpkFYQT1um81
7GbkESgNV18cSEhRjbSdbtFPPkwZ3Tz1CoujBvkad6ONu0XWAJn8TzDtzwDz8J+R
lcPZ1AJaP1KBXigjBmgLu2Pem0IygCnu6hQ+g+tYM3uEGjZfqZgHg6PcXkUuH7/S
/UZPjzqUP+cBi5GyfvdjCv+qP2/UVwl7VyOAXKi9EFSWpMc5fvEVP3T9ji5Utbuk
qTyviDzcxn7k/W8xW3DA+1h/3nFCwR3FNUrw1KMusBHe052EjwquvYixYPOr6tga
ENxBz9Tn5gWZGLYALJGP1RyRLSbMkXpECVOhcVts03t3Ty4D55kLjS6dM6Zhxb9Z
ppbUP8+GWcr3s5EhsqPNzzR8Ic2oA7N9wVjKEymt1bI8VSNBgZzA9Y0LRNWZL5by
S2rwHf2vLNJObgq4Tu/zcCwbwE3Q3VvCdZTrL5vWnWljkr9Tanu04tSXemIG2Wf9
prbWOXj5+KowGTTorHaigMLAUcY3kBx+PXmSISg+uV0ZItOCGHknYT/uCcDdzBsE
Ja1Z6T17n2MHwpABKaVJJKlq3mXHnyCwJIPBngIYnsy69oLoVu7kKeMHOCB3L9nN
W9wGmuC0kqb2+kllN7jCSQvaEHkHSLYv0RuGTO4zkowejg6S21Poj9hjOcAcWGlw
5vJF1f4ur5pYlF41oAC0QT+zFzmB4gV3/vWtb0eWj7F/6bQ4mxN+7+Jm6egZRCx0
xLX3uf4AObbzq72guyQ0k4EfRypA8KyiL0DGfZpclfwqz3UHm2n0Q3Q6Rnk1Qzf9
P7qTSxn84j7UGs4INMTHSMtqZyQrB8dVmQJIP/fQQ8uaRBHR7tbWqwCqw3xsvmxC
YKaJstRtsNfqKg4Lglui1FuZiAdV2TjIJy/BNF0cZJDobyrL6U+eq2RZURhxiNQ/
VJ2VgvSikHFt0rtKX+DOdNIuDRaASRFJhxa9WV7KGTZXki3a88rkcmpv7zeAyMQx
4WTyy+lSZApHrogSnePP0bF4SqAcHVJ51S/dYZqPHx1etPoWZxE5d1nQANjjSa44
vZlEeC6qjCPgvg41jqHS+H/566kqoigkS4S3ZujzSNdY0Jc6aZ+JPtqIq5IEkP+v
9k/yf14KCwNgkYZP2Zw4ae/k10aQSVxkjkh5/zYxB1WIUNa9E7Bsbjsj9kp+9gu8
4onskA3R5jXbOvd1c3Kwdp3TkzXZ9Q8jVWKl2+BeoSF4gCA7OLJ0HMC7OQek3Lkv
NcCQ92wfn1FwZZE+z3FQ5AQApynxuhGAFyVldRvrRsg/GHxHbW40GNR46V6ze9Gl
hrsfvUY80aj65cz0u3kcJEe52h7LTuec+R/Q7HH1+ppH2xmidhBjgDvPyayLeJ3f
LL/3s/8lHndvXnyui9kcEJr9fxQA25nT1O1g47leza5OAt60OD9NCHSeAnGm39NO
E5Q8iQrv9of/Geor0NxQ0lGSN7iGIgwCR4wH5+tCR5EXQ94G3rxboyomz9EJjTw0
WlPtIZjhvwqH6py2tBq9UtrOXuvH5Ig/bZIt8ICJgUbS+dUVJnEY28V494aKAXup
poV+fNTE8mlHNivNCALyMsP5vzyq4kRNKr9GBhmoBIkVw6pYCenLXfTQJ4DVMVGS
iNb/OvdXaGSK4HdiPcoN0HtOjwScWWE4PcaJTm7vc97kb3B33qJP8P8RfgmUBExv
S1F6D7o3oafg6Lb3cVGBFgyCQ+tCL28bqRbWV6kmVixofRJ+OQ9cAygegMX2GdTQ
gjqwcVI+45Sw/euxMirqVmyf4ZBtK090Ng1PvHBDfzsqbWIkjrCwRDUPhwpP6wDv
TlLzeVAG60+tU6tqmMDXVM+dbqYfsIpHaSzE0/WADDynhNocSibzRCb/0CTRNr5X
vPPQ4wbou9We/84M045UjYk6VDBEBRkcunKweSQSYdkpli73hhc0HJFniPUkxDGg
rXzmMtle8R+TXKh2JCg05vw3hbFfRlhtTREaO2Mhf2+9Vt/hFDRcVJZjldtJ53Yo
jkNk1TCc7ajO7TrM6oSs/HF2OzUwwqk5fcCywZDAum21DucXysIxyzzEK9GhWPmi
n5FHlS86c5dNvvWH3t6Z8qcB2m6GVuO5KO77dCBMU35qwrVlN+tSYUZUZ+0T0tHS
godnGXXMv7kBt84z90GkANZZ8CrAgrkvneLzl/0SsgWdOXeNEMXuRpKP7R2rLvo+
yQmQrU+1F40QZMZEIQ9XLo+aYrFr5ZUF+kZcYhAV4y7/wtnzk8ZyImnkUgvIehqC
6dk10s5jwUZ59oO2Ew0Z/2MRSipjNn3367ZHxbnB/C+5wiAgUaQZfQbGBXYMCD0o
9x0XPzr7sbZgkQ1LNvjBYJIm+wPF2Mh4F23Zthj/0WcFSeLKOXvPvh0+WR2YZCn6
RRy0wyW/C/onJj/u+NvNcw5PUUGmMWUmsYDVgqvXMP5tEoC1ilN6fxbeYL5B9qw+
FD85qVIKHmjmWPW7pG2Wka2ou8Oqqx7Y5UrdEP8t+ifET/5CzXNep6/gZ0AEckuv
GGeEqWBYzSHxLlGetT1Viu2FIFnERpyTF0wWAg90kcznt4afDhvJxoOE6cQknf7Y
qXi688ZmMo0/T+UA/i/1/2JBvAFmIci9Gfv13kwbfg3gXUEtygPqJL1HerdvpvGc
+N4Tt8uNzdAQt9EdnrpfA6eLkVFf0Puku9sH14fCUgmn9iwQW7eON9Z3WyVj8/yP
PsdjmYYkxDFxl6DnVyBcJAg9uQs2FWIxHjxZm+SNARygw/QQ82lnjNYvSvt04Znd
tSJc4Y8CWA8ilMA8YILRMyNaQ+4qBPTQcDPSvWR9NfHIigeF3V4jQAxSQiiVarfa
McWSCG3padX5DNl9xUMbE9/O8IqbvSYZwvX63KmUpRLeDGXxIaPwKGOT5F7lHDMr
pjUoSTIC5pONJPCySmb6sUVbBw4Z/TD0ovDVtcnVHtFIekp4Ec0PLyDixgInGqg1
/B4X/zh+Zk1WQf8AYbCpb0pDfpduZW2rNrniZJlDaV0b2g7njOdDEdJIRYkKrAoL
iwoN0XVaaExZz+rzLq2qWXWLrIDuIWwvvr1yHFGKLsr9uEw6tAPLKnobjsClx9wS
2idQD+z86WmEhy6qK/g79pjir4UVXldelg/MQldsQ8glEEHPLAItItWskqSJexUj
Ohqt1goPosRSV7ZdlwpsrEGOFyNUleDsKBMOWvztSmVapOh9W9L+E1A6TpzpTuYC
HQ1XMLsyldThhaZ3YvwcyXv32DdQPgwYLv1yltOmfGNT6Drp6OdEPZXLI6iLtTjv
N8GzrGCwivJPF/mbsNc8j6Ym6N8w16ZjAVrzjQi7lKiTgqtTfztF7zTaMj3QuLTy
gBrjDnd4q5sXyPKeXonlhyhDQy2R7CTbz0CWJ3jHM0TXd8cKfLn1pJGFIuAOnCG2
A9MJsPhA1mMfmcTWODA4MYU1gzdCNgMGtCDoC0Zkm0GEaVC4lEtgc5nKB+D402aC
Po4pLsxosTz6LZ+iavhGpMA3ptmV4fV/MNsxBxo2neD+UPy8azRcZFSRe6smezyV
UQAbAoZq4UXqYMqbzNfxHX8oh8XxDltxPCt4RZ/5pZcrUOc8Cyue8h56/6JzMO8A
5q9tcYBQwYtX65jGO1mHhaNa6BV0nRABqbVo2aqcfRmlJ0C6yFxq/GTc97GgMa0Q
0YRb78SSfK4ZJ2G3PUMWgmMBlFO4Dhu5LWQV5uPRBszKQS8QHmDavgdd1aaVtwEr
rksz9jQfuZtiVrw2k7/xavv9ZDueDrbY+/msckdy9KAGfprkB8FUKgJJArYA5nkg
KtQ3UTuk/DixIoWA5L7o8e1BAi2Q2OlEAFVR3OafHPMyBSbk3tNRVRMTOO8EEbtF
oG+u5KXqfMasEq5/qcYN5zk41iuHbUh17XIlQhU+XfDtCUQj5L3oMK35marmz7qu
Ow4lGNxdsgdy6nITUMWkJr1sJ8iQeJWJzFhXCrq+78DcEtmNAnB7OOxJNRutjQ9T
BPx/+vAWxdBrXtHKFskXfOEml5TTcJLicYKK2e9im8I37K/jIHGPEMjuvn6XZD4F
yT0pjjXo1/2Dt6AD7DjkymfJp/Hb4ZpsG019lQJfkg03m/yfLn3spYwm88+AZop4
SEL00zloHnCPx14/nHiTDDNQEv54uu9sJOA/YGGNjfN0ivRIZ+PHzROpsYnUGLUo
w8VuExxZBtjTXC2rnDRAoNfj1YnEZKvTnKe03Pw2T0P6f7Uk8b8Z34dQZjvVJ2LV
VdTLESakiuQpLsK6OWc1kM+BKg5PFcbXIIsAW8UL7i/gdXokKVWgtpgucsypsXaS
BajFkaXZ1Is/V1mGFDa+ixe/XnH7QEsi+Cxr8dybSVNJdcMIrRKd5/OJ3xLhIl31
EuhqwYLMqpKlbCbe8vHvgDZzZ7KuZf7aacP7AnfLpKpvj4Q8n2Gj2Y2CpyDo5e0Y
4eYvH6ozZonz/aM2QM9wZq2Boci47S1h4RC+1kZr6FQ0SO4wyIFYW1qJ1s7GCpBG
RlaykTYx4307mw5VcguTub9bcRE4Zy03VWSqRc3fB07QyUqDxMTc0FJXPAwm2Ibc
8LY0iIFEo0Nl9TSQ4Y6Vhag18pzT+Vje77SFpP37rIL5sQE9bBSBEDBenjwSHkJ/
L02sT2WaGKq4NT4aWD43pf4/K8gIXDsNvOt0pCm50WaHWJW0TxTu9IKKOGXWmqEz
V0OAuPuv+S+Vv0PuzIwzt58U0ygLbkhN6eH2YvrS38bYQyimhmD6zyQRwQ/aH9My
B8cXuKe16LAoS8ygoki/Xyev3M9B52Ww0eSO6RSBeYWd+1og9fqnr6SbHBNbaIcW
EH755BMGBicsvMcZH8CpkOVlTfnTwpfcgGvkWkkr+NEK9CFIiCwOruqfa7w/8L5M
+scASMivJpKvrIAmdldnvFteVQmMHkiMynNJP3iW+SUGAepgUMayHsc/KH6hTJJR
IdW5+iSdPLolegnZ9JJm/7yPdIgnCPmHQAKwtjZWiit1xS26R30to0GABKjvJcBH
Ey/1WF4D6kFtzNlQ6oDOeXGFVTiRkgxucRgWBD+Bp1PO2AOdUxPykNwNTYEvbhAa
jErj2jVReBxTfNRcQ7wWvm2hSCirxhGaGWgFKCmnuMsw90kUboZvsTgav6LnVam2
cU+BSBy2IhYPGyWeitVAUScjbAvktVgiN8kyG/7uYlVw+LyX/zSTipgwU8h9Jib0
CsixNf3ZvKuXJ/0RYi0uE0anqzXvna9BO6IVeR3EvHX947e86m0hl/DsvsZTWuKe
W+rbU+/A4tQmOvs+yu0EyMorhPFk5i+d0+eiLZdiBrFK+4Xoq0VOlw4K4H5X/va2
wROttoXbsoZSayGqEqvcAealNyesr3RdziGuSZkIJZFEi/GnmjOs1RlqGKm2P5LP
R43LKjWfn04c9D4btkQUcwWve+7T1Vk9iZH+KnlRNttUWHnOGjAuxMdrAQxVQn/d
Lw0X2SShH3RP/tOwB8//TdqVlqxqNDS2pwqYAZDDhh9WdQwDRjPzJHd9mB9EzSJ9
BAx0b1CvAGE8UGMOxkJqY15xmKyR+H6i1Y9Iiy63z5Q+kA9MaqsBE4S8NG3HKuqi
Y7Zt1zPedvN1+BTAMhmivmYk5ogCfQdxz1CSkh0anetcg6S0c7Ph55wiMa0kPYwm
9ywWKtEp2bBI2p1kbwl6SmxHklSQJOOb8Mz8mQAHIyyLYNpFgAbC1ICv/GE18Flb
/8Y+qPvpyAVtQSWYMcISkwnU2NMJEH9QAJwSLF8J4bBI7WUvZifBAvRuZnrZIYfh
PQpbe/kPCtwsZyWwlGri72qs5tu8Q40diLtB/1H/TQWSPVDlY5id6eP8SPvVa5Gh
HPpKoHIZS2OkFNoU3UuWw/4K/99hoW4VrvcfzSoxFLCeayx39Z+GGqQoAGlFFoZJ
2AXqmh0Rk8VPpUvhe0GR6it7yQLYFFHtyrQrvbwEjY0mHdFaQ46Ce+5/3JCIMHam
fe0HM/nGlrSDj+e7XxcmXsqlDMpP49xsKb2H+eeRJtMFEaL+FCWDokTbjOLZXkW6
fZWTBRyFrDN7GZMJ1shiKWFozNE9FTRUJFVFgwK+z+MXXWDvmIXsuP+Xsr8P16aV
Re/mvh7sPwYkWs1IhixYVHfe6cSqo78Gr0RM1sqZbA69M+EblDax3qxmm129Cx7s
QJcq47EWkclsJB6sW1OOPbY+I8LIu6uvFdgWxVWz1xpDjUm8EBxnWzaCd1hXehyh
X7pEFcJF62GxgfLlPm3k7zAUm4okvGKGLE4CU/D04Jac3IZKvZZzUIdI9xj2k9Pq
ShPGIU7w854Q/Erp7NmAkdQZvC9Dq9j2k1LrbBnJjOKlYkz7Hc3vWPQpB0sCp0TA
uD2zsm2QaY5YFK299WQhjdO7bpCFh/NEA3HHLOqbkCOdD+rDx1Uy8w6fVhwDUVyB
eDGpUFx6+BetoJyvHHs3GUq3OhaDvoPyshnlJae2f0vh8YWDfKa8wSRhyyOhdE/B
703TSDUmIFMaUGihyVnIqCHJRhlvKRGUyX96jqIXm5DP7ucO+rZPt7IWBQy1iRp8
7Gwqpw3n8ZYKO22lGupswm2Nhg3O7eRbUBVrdIVAqbUXylRfwqYoQxYHTXI17fjZ
92A2Fl1ckSQ7/os1x8mpTyMiWrAxB9rCSlMOMam2Te+/ao5VBO7OX+mwF3PPeVwI
V3h365Zl8nk8Q+U6IzwW/5W/ECT7a8mK00NMh5Pcr0eKmoz7yf3CXtWGgqlsYyGV
9FpC1IUpJ0yNO26fd9luvDk0ynfJgk8W9CI1XuKWvtLIl0Y7IgpTTt9+H4nMXMoV
Ul0SBIbMGoArdP2ZU1Iebg9XqjCjd0LRQq7Z7AGW3mab8azyEkEiGz8CEae5tlSG
u6etq6rP7LaxHRqLw/MUPxp8hmrMfMYstkJ2INN5hoEPKZHJHhT3gMVEBRBjRlqx
bIeLtbn0WfC4tVclKScDHLZ/VFS09eaPG6khHGKmbfwx3i0Txw3A6EUws+4hPepV
rAskb7UljVeaulOATn3UOR3g1uTMJgdRc7I5vIYxA9UT12wn3gHAg9nqvctXKmL8
O1H1AvIJgnUn1shLQoFR4yXtfzXJYsvMnTAtcJ/ra2oLGvYqXz/gnmKlCxx2CC0I
0FFZqEjzcKB4EUx+yAsDz0MaXHAeWSUjtduMrvKLf3bxcmzW9z/udyk09rSLtUyp
6FmVvmxmY2R7mw270MP3jclqXWgjx17M0erVn8Ad61FkjZUKLNUKZciFDOMkcNqe
5AbwHLLudISLCwEgK640LJer7VaSuWKHHqDUXtd5HwHciiqWlFd5mr5sZHsnziUt
7GQZ52Jpuu9mn2YGgsDcgD/lCm+LWdriGYigYsMU1gHkv5y+5heojQ3OV563wFQu
oDxSNlj7htryUvn+CFppyCXTMa8cudDEauUAqnqXhrg0ITbVm9hY8exXkaXZrepg
7zn+yP5fY8y9KR0n+m8VkNYzdyatZiNJiFDbqkJ17CuOrmV3H6mklqB1gwLXQkL3
sYV9cPtbSSBSZmir6TaBttyFJLE6i5hF7YFMQ8S+9ajdnFOLB0BN10/hcUycDTls
hQrGAbm8UkgMZL5vS4ZC02pdfPLbwkIBdu8Q1AtFYs3U6cRsbZDMkacVtR1z3K2S
P5WpcG6AlQwhA736saWEVQc6K4Vhe9InpReoQMVmtiWYh48/qgvt7I0CAAq975bl
JFUknLS9KocnAmLze5QnmA5T7F4JqbTfhswHc6OIDhm8MVKU9kkSEcN8jiroRvQ/
jzmiKF4nOQD4NTh9aMi82OHY2Gf1gB4hWAGNC8FN99MO253YyEzyedggOwS+ppBH
oQQ1G94wUoNpHgHZJ4jfbLiN79R3seSWeFR0IdCuLMPlz2jJqMCG16jUxc+53Ujb
EfsCfxgxJH5N5MxfDSjk7fvtacLXWwXbofgEbFGH4D8JuFXAmgBoh3IgPRJhNlVo
sMuyqJCVGSQvEOueSmXIIydVQifElETU+f/rFGzR3vuJqaH9fxGiBoFmXLsjdmhM
6Ff4TtsBIshxRw8YKcXZR2475ob29o0iihe4TKq3LN86MuTuyEcSxiUAsiPQu8eB
7t8rLzMk7pj5QIT1T/XY3m77Ssr/b+TKpKpfaCxXJqh4dLRlvFWi9ZFeLBkftdx7
5a/Hnen9YgwuCSXdE5oQUUz/AJnZB6AfTDqySL2a65Lzs3yVxxWBYRhO0TV44KWt
r19s/3stP5gEkvmwSWBZTp9a5wiAmMypHKUbB8VDB8pqvgOo2DPZWC2f5CVAbpRm
QnEFMWRG/LNrIaFRI9rHaaEOmzkDedHFlwdSd5ADd3gffoGzTdDr09oqXKfe49wG
0OeHpfgZHUPcQ3/TcfCJNG77W0S8u34FDX28uvje7VxPP8J15qi2UZ9OW6L5TyKz
Vy/5AexesMrT7cS866cjvwpJQPrbZ/OS+ILiras/eQ9ERNpPkc6wBOSOK/N/ehtD
VwHmtjhoPSZrlgW0K0x0lf3433Dws8dII43IUkKPRuXSoj4heuCamkymhImOxgnB
YKmmm83F6D7tbBXcAM8LrkOjmCuhRtcY5eRt3BXr3JXII0TEvqw0b6uX3CuODJBH
gXgqwmdoTNkzPamZlLEJqgCZcI6I2pyA6B/071ewd4qW8QVU4kPNor4H6mXaCJGm
2HyxVgNt6VBH9CsnPLVh8NSTfeQK1OE0lTS9lCXPL/r/frrN9ZRwTs6g1gacVDws
k1VQnYVbc9/V114ABW3y4YJuluk8IM1tqz5MMNQYbfgpXmhYKtubxew5vKHznY1D
9R9dCfR7ne/tCKhalGUbIHtktd76VxlHIUQNcyEqLHUmGtVaIkF+RfRi6+2kPrhU
vL+UdI89dnCJPnv7SwtUrINPNeP00JGrzFM2mmEajJsKb4sTg15RBcaC32IVaigo
4wtFNDb2r3JJkif4btOKyae65qaPhPWQALWcEMx2+RcOkhCLGp92yK9djgqt/8SG
ZntckxoT02iTFKfDlEghUz33TTB6jiUKwVNOE9JOH3QBQZW5RaWoQfqHZ1RDnGv6
gIxgfiBPlsnSw3Y6tTYRp/s3UR8a4Dn0/kTUSO//N18+1rMyRc+1E/cCDcpJWOtU
7ZIqshVKL12TsFeWmjxvRZb80aTuipmuI8gzWEmySYoZnphyfVOdOI/ZQaysIBmm
y32OT15phOFG+M1N2bFzdzu6xS2TbUDyCRbVLbCrFMRXu2CKPU+RZm3/DGLOe8C6
L6gTgNXkRts4MamuQRZmuJX5ZBkvQRrE2wPa7Dd8Ds8kQ7U1ii2NE2ePuduuCplw
4rZ9pkX/pxMk+EDZXXMP1jv4qDCx1Aes6V1nvXKo1VnX7WaDPM2TQWcQ/0l3ZqEY
/uJlCSkVwhyGZQ19eZmCne2COVNLj1yZmxklZYNRim6+wsk4Pkm7FUrEhNY/cNBy
7BEUxhIvy7yqzoxreUEZ0ybGz881HKeUzCvlmA3AzhzeNJ7i2KcGLLmImvQXp7rN
w2NLwNm5HwqO41CFE8mCOM7JiWRFRJOIoW+6ZN/Lhecpq11F6DZOQ5b4rgLMbQBr
R0qibhg3p4ziCZcVWIP3PEToHc9x0bDsbByLFaA3snRcB5/uCby6raMmc0wkSUlL
C6KDeX8MowIGkG2o4E4Ye4nbSuaB8dESRfdH8p/0jJ5zKkEOnktcG5/dHU46JePM
nbcus2c/YqqJOpfr2OTQsyYugJpalS6xmQ2NUPu9lc9nIHvDnKDZxqtHHefeffEt
SDmQYjgYpTI0AtuAr9/n5nIDm9NWZJdFUZoDET3UP1t3e2aY8l9ZiP+ljIGvbJ72
53dGOsorqVeJm4U9GCwGe8ZOLDCRxIewRkW4L2eg9Mvyjsm2QU8N/fpYZigF5LOe
F+yamOD+SAVrZvTNiplKK4rnq8OuT44WhLMzPgjgmc87THo7NV6E5zl8TNljDgxd
JYCXpqZC/fKFLO5D5Z9xbmya6ivVGXVl9cEz5EfeGtWI2s2fUyIq6KK3O8V0PH4e
o+c00BfAHRy82ogesJDy1H6jtTZ8jNKQ6RqzSoLLdNWEvtOPiJdxwP8wXOFhCBwm
1cfid4t2qrlrVGRIAaPm2melRAtamxxUvs8epVQBVhEtyXd9HP+Rhu2S5Wg5B7Nn
NmwgNvaCTQEkxn3+ACiER3PDSoP/TZcL4mDdR87veXqWbzLMo1AVzjH1x3Wi3o+e
PmO87URrCfN2Ndvg6wdSXfB0NpQBSatRFv3nlr2ho8Yf8YiJ1qouAwe/6OGCQlco
zlvujPAZ5ZNeugJ6jptDpo4qnpwK/NMFlctO+aOZ5ktC7Eze1rSP9XX/QyHmstL+
wB1rdFNKHBMQpZYv+1Fb7habkPHlslWWaIG0UzMo4BCEy0vVB9Sl8ZWAwXJvsS7t
uFYgfzrCIaSzlgDa61NY5Vw1coUtg2wTDrBUVqewNONY7DZMrzVdqHhBf254XmrS
f9K2zyh+7Qx1djMyA2W1CcnQPZMYkcuwV5beEPVTZhzdFvjgp/J41h8MBnvyE33m
BYFu6flGwJZ222LWt8arNQRrJIiCz8631lKkgojEycJ7BLDW8qdK8kQGnjuG9vGQ
pebkB1BJ423b65VzyeRPlike0gW8WZqp2kNLq0htI06JZUYYTtb7yKgPaclx7dAP
L69ZN9su/GjvuexgYQiEUsQ+uWMhNOQgC977eTUK/BNe0YU/UZl1YJDd3ClW8Rnc
28VC72AsoY2UWafDfc9KkfM9+o5UVUaK83dxDIhUdaDIoT142/50Ui69NprP6Dn6
PYyvNIbwBgrnVQq3Dhf0UrTPnT8mmYJbZQaDCoauZFfJ+ONyYGEQXSW0LfX3MViP
rBxO/huyjKCckRTIm6ppMqhSn6eJZzfdNrkv93w0+MYY7iGKG68+EaYUb5ctlzyU
iA5EiMqy14zf6C4OyslemjAKwCnQxk3PENHImDDNMMPpYi6UPfmwsS0+g9ami6fa
qvp43FjeTCU3BtJ2i80jrOu53MJSBmBv1yhZtc4Zb+e5HZzKcT5lgC50XOKAhtoU
gi7Frpu5j8zpS17F0n2bP9DgGGZzdiEmc2mKBuKzWDKfxVqxb9TqQ1ihKNtpL9FD
9ioFRFMHlFi7Wfpo6LI76ammr8dV5DDij6CajcvRf+UQnm48dwIvtkVyl9VrPH3C
cLNdEwql5zJM+8NALbODgkrC7wafMSsnYfI/TZs4xVCjomggFwx1pVJmwWSI0eXV
ixgWji2Dt3GVybp0ORKTpEA87cls2dd64z8haqy9xkVmxMYwFUfZTud+dI+w39mQ
GHjr2UIl5Ke0jc+/0Tax/EWeYMT+9wfbn7dU1xDCw3MzVq+n4DPbKUsXO9FQjoBs
+s4xu9/6kCgkkeSr34738cYgVbCFrd0Rzkv3APW68IqbI2KJ+6GQXqvUewsOt9gr
XvxlTZ6mX7zf0Fb4N57F4z180FCZuwI11w1kQUjdQlt5RBk5q/wTRdEGRSa9QNfu
THFZl7hlLfmOQFsi9FPLW4sk1RnZ2gLZ8c5Cvx/YsLwzkfZkXycdBNCGdqQxj5Rv
rD3AsSltKuG9KSEJAvvLoNSpiBg5o7cLuLnrPlptqfGhhRCPimitxaR1ST9T6fgD
uquYiIy9g2GHKzuWaOzmBACkqInqU1deNKbccm1R9Psn9QWgBm0YesaCvaB+qFjF
0vSLt5vn/gl8l9PefudSmnWKf7VTHebkq/n5cCgmTCCAW/IfGcPKq4GBLm2qc4RE
+x9/LBFw94xc7qHQBMv1CaDWNeoBGP2uwmm3XYsHaZ3XI7Y7x0E3KktM9lezhq+5
B7tzTnTHKuV5Rp/e3erjezjhBsEE5NrFne3o17xh4IUxvS1axdF9V+ZENSq2z76E
n3MPSGhbwNC8hLFhaQdosWPRQMkrlfb6YI0ogUu4khnoqHn+YfekPZO/yaSq/6C7
rfiRy9qITcGyBsW4JKezYS0NxT0m5OSN7uvepX34mmPd692P9K5qUe+GKIZ5wPtm
4h1P9fE+/BOtGtrpudqYzrETDF2C1OgI8llXaFmjs/t6e3NTLoxDXlDDHF+EpfDa
W7VODkimHt4raHpmwJ35FYUbXTKOQa+svM3Oq7ON+KetslEjujT1YZ6oqQuO1Pho
tiHjNvqZxDRNBkCLPhkZFxyVp+0b+gEvwY6vXIwpgRdWEprJZffQxfVy7aKVB2S2
T75bSKbXykqRRJZeoqi4vImdk6Ga0Ed21WFCIvta/rq/aRtR0VZk7coT/kPdGaTS
hnMjamD5bJ74oA2+DNf97GUArks0vC7rfEzQCb2IznFd16z8x3hlxP0BrBmsLZL5
vPHMUsfFwhoKIY9e/zsX90C6m5Udu2Y/iP1NOyWsfPfOo3W0zAZP84u4pZdEG5En
XHQ0RirIGmWioeSwC57WVbxWjt9qW1nda8/pYFuXBQCMdy49p1+RdAqzl8NONLVn
N1IIdUJhiMIM+79RbZSDUOMeuZIApfrSWcsN2woC8xjaRspMU0d7UdtEeeHlFIIk
j+N/wi4N0KWlh8Hy188ZdMDBP8D21zTX0pp110RS8eFsw8q7VotVY6A3yCHXH99e
krFbHHb9l6FYmIb7wE9A5VK/183+yFJhugUvuHDAsrYsYS+5lpUMeMVw6LaAl3P/
6GrsnB7heZYxgc9wYKm7cSmIXBZc5lxWm6rbP+ukSG24Uuuldo4H/IOGRTk0RczR
Oz0SX/sPlULc4c72QJhft/AC0QAdZnVoWBy9iggtpBfFBDbDp/SbzhQ7nYEj9BGE
es1fshmWS+1qP+xnnqqaUCe5y84rJp+TzjnoUzEB0WEjdUtCSAVmrSJDNKSzHA3l
USUMw6XY5VigMaADebgCQxNws08htTVnO3iN+FfdK6AkxAsQypoZmlwKu0FNFFIk
xBuIjrFf2emZjvmFiUOPVuWQveTI78u9TpUI0wumN2ZDLLz6mwFhBjEuRlUzOQWG
iBux+dsjnfkd7/vriqV4ZMlB8udM/QOB+sMcF+HBnMrtNo3XJvA5BHIxD7BZarRz
WS2qks0+PISjZitqqH0+iiVFuezzpdIeCn9sl+oN5ZK854C9pldcWnM99rRZ44I9
pzSk0UWIj9V4AuoJNO5+NjPSg4uac3FAaXhu5Q7HNsBUIsUAQ8E3WztwTXBX4CAU
wRm+tRs6WbSrBXMqX9JroY8zx/EjAJxT7/1kSysNJqHNFws5vLOrsiU3+lKTRj1h
yV0wkrctqyONwPI6FbNZckECBENlIp7Itel8vQJ4j7ak+7R+nKAoiNhZwjCMjR3V
nch4BiOMozQJWdWUPY+QNq0hchivCrJsE37AQywTzjaD+z/26CXqe7KrIRisOYX5
QVkUPjlH7B2waFHWIowhfz27VNHzZijFg6+Wo/rp4J+kkfiS7/nKALn4jlTgboZG
74QKjvv7iMxIWhyxyKsh+q4kiu+nHzIyPGF7yuts+X9P3fcqCnAzFssXYWAIkscj
bF1hQJKI34qVa/Muhcz18i1OPk41MzaxQcS+YW9CKJ7FnWBKARpdFCIdIqb0s9d1
okGqNlBU18UGi6PXYrhHjPnwZd+tMXTC51RsFb3e/Uj62qAmZE2AVzlZRPhhPI4L
srUCnDnPtapI5nTox7lCV1K7t7138uYTdEFoYBi97pTp4kU9uqkRIxIto5ylLZUA
58szCx2+Y5tXxuMXOADBijly5I2CRGV9CDJgWjoVyxFjJ3TY7ZD3+UuvRLtgPJt7
BraZ7OrCx1uJADPceUIOlMr2Oq678SQqnET0TJf+MHgUdTtWIDGonTsN6mSu/Vz/
zSN21rsE9bKFtlYNKN93aayFPz7oT2FS94+GK3BqlYjwWNhNCBGaqc4JfhGlBnbU
VUKeLOa/6RcHaC3fs71dA2RgixSP55CN7hgJ14VTVXDFr2/2BoUis94PnufGaFrn
O8LtLJx0Mxro0M4Ztyn+Lac8pnmn/tOm0x0uFoX43liJk+sxwhMw2KodTCwFbCNI
QNpMXAtAc4cCjIJGTIGPd7WRnkjgC2JWCON4aNu81O20V0nDEQVHq1J7aCcgn9HG
njEz+IOvMfgc428SNlA/kBrqhzkZZw1ohBof8JlF0tQJBLlw1cdUuC0bR0IJYkoA
VqH5y1QXQsPKx/U6GrmLihU3AwOkGTxnm5YKEBPQvoAP8t15SvxUJ9D3B2loOOVx
47celktxX9jTfPkoMDoDD7BTAVJm0sDaEj3345qSMZtdEzVDoOYW3z70D5NFeGRv
G9JilNE3LIAX/GPEHtaDw0F4ZwyfvTlz/fknk/0WwjDRY4mNVc/VjFIL3bLL84XC
vztpHbAudPzlmIN9yM+B9lhsUZA6L5Bwj3cO4+Teoa4WLg9KFfEPtVOybYg5RMdz
t6SKbQWlNoqHV0se4iUfYgndZ6HisVE0U8iE/10/DMsH++jiej/9DULJ3TE1MVVA
G8oHGOYfr9i6R5iThk20zc8MhZH5vjo3wKvom7HXvZhTrE4NDrb+bjrbUdPrCMyY
vH20j/96nDh1O0NzAuHvJFYawub0InxW9idXYBQ0rVAyERB7tgmAX7suRuygUUUX
+bFWd9b19Pw5koXEjFKBkmgUsxuPolZVi/MqO+NoxVuJ/gYaQhO8F+VtR1pkeKs7
JPnIokFTJlQ1eftEnDU3ApcjOKxvs//tQs0GC0WsKmyvLGf5AdmWWrPjtufg/eXr
Of6zMbI8o+YSqlgpXbh4Qm/qYcuJfCdcAv3eKVgtwJu3aAGqxrGEntqv2uFbys5R
1skvFFbWDLullay2WFbKPo+p6CHX92IvmqtBfnHTSklcxeufUx67EirXHbKMVFBf
qSdzlO9PNLlgCm2FiQHV4sP3jYqXiOVV3vExB11LhjXi5NC4QF7iqsPox6knrdjg
CP5ZwB63snuhiU5vmrVDZ48cHgXLYj8GOy6GB7u8Xyae7rmsMGLIhQDRay4hfI+1
zxGp3RYReKU5egmnCpu/nXzJQpKOIVGf0kM8XsqL+rh3Ij9PLaCOmBohgdXlwN1e
/YPdtswsuufx7KKJx31PMz/wBnPwjh2WR9zSYgk2anLE5Qgy6OIVwqMfr1WAGMTy
W6DVlxkecqAFgZjZoa7qI1m8IC59dQOKi7b/9DgJ/HDDVzj+CcUCHGR+U2Lig8nj
V2GLlhrnXGH/vXde0KMNy2mqHkxt2avZ39k4yE0gvY9vVbp/2dHUbr7GtD8Ffluz
Xabt9aNpdbmzuJF851usU0Tu2pnie8tD1e43cYb3ZlVDlBGB4hqlHZMKvVMgTkAg
2cnhM9ANnJZeHG7oaO/FwNxcjC6rSOjpbkJFzRhEgTe4sMs2uVa7ueue2I1OcM6j
OP5TDHQ0V/ssXi8ctq9k8HycRbvtdBVtbpsTeZBgiHkgumZGN+mw78HWW4BvDewm
DCuYY0qA5LoQ523jhV6hYrmh+qxYLtu2S4Du/A4LcRvRyMVn58ZPClQDubYAFpl7
06dtx0JDuldhiig3/m4aD8m5uf2AQA90bCGWgodmxs+fUCY35TuYfCudffOSbn1z
fTOphavBcrYSE1uRLsWbor9xzCPN10B6wBM/5jJXASkOp5bQ365L5KepBBv6vyxi
BjUbYJXHuRSJDJ1258Bv6tN9LlEyh44bPq2th/byERgSL8knBbRExVQbUgv3Eloi
FfW4uWVkr+rykb2H4IPg9iK3t7f6KhwHG48rygx9CsIbt6yuv7bD6fZQ5r5+62Uq
b2e03M3Spt2DlbMs7Bv7X+nxYNT4WZEDqWomPyQMpX1YViwJWG3lpCb4yaC8xW/3
FhQ3T8f2OSF+L1SbTofF7J4kTRs3BTGSKXLQmEbhZX6hmu4SCgq4pTkVmsaY6uRe
1WYbCF46x7dpmYgEWUiWneTZBGXu/8eWeirWADPUwXnjkQIhv0G4IuPFcfFofHL5
Ax+gJoYyAXpUMgC3gJxDahF5xDIWBeu1F8sUNbZpZxCjRZoWE+mE0Oygf/dL+Kk3
vQ+hGRfRTsIzGHDPeGCPjrAfloM4HAIMA28jw5R5w+b/A+L3g13CfWMOt3t7vx8w
HMu5PXjwPcbpgpoJhBTnR8hd1hDY5O/UeqfwoTuabF3+ddjjSbnqkiN2850clGK2
djeekZGRVAk41aBZp+T3nXKtfFxBO3ygfjhTLhdY8ohfVtummpKugEu/VqT4QwNU
jiKH4tyGle+u4ckg7KnzlaIf/D9wWNYtpYscmn9u9g5Ah8dsg/YwJcBG5hQuXmcJ
A2Dj7X2m6l60DlRTMCt75zc3pHdi9/AIsXloAIweUdkW5nHGlzIaqgpH2YZ5g+Bv
SOYENHNJDoVaaOMpf9yTDQFn8C6c1Y1D4V7Aw8++nqwhdznUXpJZDBqf4mfctuJn
GLV9nOB/tV3H7ORnEdsmIv+FUx9nHUdNPns/dArTVgV179XICysq/O82MBggx2pM
SoQlWRZbQa6fgdJCg7N88VEyQOZac0I1lTm/S6uQ1rqtYiCQ4B6xGNonEQm4TbMu
m1esyzqR4d6Y4XuqkDGdZZwz+nBO9NVVkE4oOajRC5rJl+p21xS8/9j/nMwY+aOk
3k2YmKIAGNls0YDhDBLN4XJLJ/w1gtMddzYhJ+pUw0xCKjw1CV91BbpBJROapd2v
MaHnf5FjwD2+mi5t5+Zoxu1Z9HESO82OBWslyLrdT1W5c1o5n3a2bqfbkKlOL8NP
LzGYKZ0zOSpzAKXT8GFNmjQWrZUr07lHOYSjRZaHBHGQXqDAe880zPjKFTJTQq+k
AhGDN4CbTTAqSUW4xJz4zZ5P8CYW9O5TZCsMJKdMf8n8u8Mkri6E+X8sIUJYYb8a
dmQ1pTEj2rlfKdHqh/6fCWZMdm7ajcd7/4RFGAVs72O19L8AgmCVO2aJzyrRyue+
RDAFwc3Ua/uYaA8UEUgHJKbT29jCcgVk2J/qXeUnYveoDzdBzaod+Qtb5mb4TW7u
ObJDwxyWsbOUraY0Zrqfl9CAFI/FvwD/2f2Yu/6b3mOThgz7oR+64gUcf2m9DKbS
uRX6MhmS4XKabFnDg/dMLkoQH896G/rH2wzPCmxmAOYLDAV3CQwEAte3EG2OEaY7
y/DcrgE1+ulhhigkHGZKNkJL5zlBCur3i8cnMBx3jn3Ylh1KOfJfZ9PmqM4dMC3B
4iNuFKxLI/HlVMk7BL4/GYQZOE+P5d3AdhNerjsd1aKp1cwSLMzD3G4sgClxK31o
QiAEumBfikBgLGNjWQbtkHal9lSvtLu76Nxvzr+EK48wCaKg1iIIulzweiBN4IaD
kCDsUzdobo/ELwVw1mA04NgHGsRFuQWtxQmTxzK0VhzwPlfGMJKDwTnClXcbjN2Q
ba7ew4F270ry6QhPio04ix6vtP7DZD9V0z4nfoY8eLkKFHJOUxZU220zJOwQHc2N
9lp0OSsXxF9HQwQp7CpdSjWTE5ZKRZZYdfn721eu2E91rfprFObtjabTQz7CWW+T
y9cV0cpAQPB/TjmpbIK+JQZqOigbPa2B7cN4xBOULIVz7oodIO8OIy96K/8H5l7X
tLgJz95nnXUEh7CQHHTmH+7nKMnW2ajDpgST7DRckDTGag1NjUUquLwr1hrFhSh3
Ycw5RRTb4MBOl1rjZiU6Z2N2n9wXJ2s/HjszDOqYAdOdGvqEjwgDkCKazzLP1Ju7
zUstiCiegK8FcjjwJMmYwgnnzMIACxR3rHvqOIj1PALELplrkV6TnJ0zMM5xWTQj
AJQm9CAFo4Tf6pcmlWWJ7X8Bs9WKiqW6g/asMc7xI7kDbCvJ3qjltmZwZEE/VakY
lRxCHHYU4gVvDgIT0gB/jm9toI6uoL6xPGvk10vHJSCQaqPLYooBM/lO4MqgvBSK
9XqvbxnNKm59UKM2OtWP6dckZ+I56C7O4eR/4hRe/HETQa0AdbZGw64pGvRbDUiw
J9G/xdEx5g7gzp3tY4k35rblKcsFwDt+bN798chlahUiIRevluxpGUK3wwAINAWt
B3TzDxm7+VU1rGcrR53VxWxxhn8pl/akWmgH9UVX0liDSZGaxQmPoAQPtXM5SmC2
KRnQF6EMFuC7s6DZUf9030U4ATx5hzlAvsBtFZYmGA2aZTrEwA2km4wi71VLuSlY
kLwIAZw9ZvLMI5F3+JCPLCpsWSa0few+onb0Sr9ABpwLQevjOHNAspIWK9sJDhP3
jwCJ0mlEzbLHE7TRzPUPldf7ZIRtosluVgdSy58sLRW0hY+wOMfcWH5qKyxGPYpg
nBansExqRUnld8QlQ0FZhEF8ewVvz9EmUTDTfo8ev1QL3gNY4+J/ZzuCwq8TuSRo
Ohjzf93RJRtwals9jbEBJ1MNTvF1TD6dW2eXe90Box1aN6d07hF8wUSolCIw1dVr
FlogEsE6H5qf3I4A9d9Quu+5nB2Z78GyaCUklCzxhPzs4KCKVxN7c2moGb0Pk2xZ
uzipvQKxQyUYm6IrQycVP/BwmdUAECmMficS77zSgI+plMojoxmaWU/Btwgk1s6d
iLOZyYVai4+NZKXjuv3M58KA3lfAfQNCP3GbuiQwX1Y+uNiD2faAQ5fnbe7wUJVe
7LPZovrmELuJzWo63CUI7CQx2Us1ze+XTIIGe7xjGqf3EfeiwOM0rJu+rrzSQq3W
f4NjPt86FRJ+xyH0q/FazpvlU/p5jELOKQJadydwFiib84Y7sz0mMJANwpOZJnUn
E5XZNRbkWm1vOfs7+8LSKggY4JJUHFiht+HX0cFwWwWzkSkzn8bLHeFdacq7lMIn
icHUJQqSk/GuoWLtRu9I+vPJIzk7gFh+4SfIj46NIYLaBb/S8qRCp7FGXKR4IbOq
1ll3L3x/FIPzbkHMP0YsCd7lzNjgkHtjnvoEuKwRWii2Awwd15vGOW8ZoWPqcOEi
xtT9xqFsy3u9aARNJJ0/UqIM22K4BMMojg1v4d1VgVdW4Tbybc1Csn/nrCIbB+Rp
Um4iagbQXiBxbbGgbQPnzayQyo6RX7ASj0ns5GskOBtujxop9tfztb/U+TcZXBXi
phsIxFmhv7jy3YfNuOo8LMRWfWKm1mcIy3nN7haSHZ7YYx9ETeqD5F5yXn0OTDco
0VH+6R7r2rprNs8yQXJugcw+8DB4Setje3EHSvcdn7pii04cr1VSCvTNkYdwytVC
jTlesqmXkYfOwCTfzviH9sod6Eivsqy6OaeDNcmwEzOSyiU7MGcggWJDASl3V3YQ
KH+07lCRfgtel9W9FjYNnUmYqeIBWqpKV2s+cKPhTwsJZkAUgWFgntJ5cQP6eLel
oQyADHvSZ5m3lAhJOzqC56KdpGYweInmyv/+tUM0Hu2SQUkLM3z2n+0+N5ri22Hd
ZU2OQgYPyTmwThm3sI/XQFSffbGa1WV8wcrQuymbj1EbaLG20YQjrkVJO/Msp5qT
EFr8YWPjnHeR92Qb+KsQLuFhRi84TeWIEoetmi0AIG3BM5uEk9BMHYtvbOgojx6g
SOlA88k9Vh+0h7q60eqBkTPthnMazWtesNyxLzD7YTt07IjqkGEX53QegcYPERb4
vps5N8O7AHle63g6V+Dsjh686Jf5Y11cdPTt6FyHOFQ0NPBELMPw/4cxHYTP/Txh
4MyqaTxrkU17fE+CJwjJ6ZjllAYRKbpq2q954euN4c4DA2yVw9wp234f5DRNf8dJ
OMsmjv1tb4EZwWUs5gj5MnVoPwbZlxbSy+frQPo4cpCS6nb+x23IWUYvCApjd5wA
XkjWYw73mV3342Q0N62XkB8kTd/IyB/iafwAA6ZYsssMGJrSgcpzEH5xhxJZG67O
PyA2OOysXf2RJME3qwdEJj0kTwwM5f3JLcip2KCI0/Rv+12gSN7hi49lx74t8xEC
wmhB2X9G2TJnfZMiLMaOZcPoU6pKpB0jFXuAMk+cJHuf+OyfEhEi3kgomlcxMTy5
DLftlyeyt+KEa0xRK8L632r8aCEl+YXgK8CjN8dFNcJtRNEsLDst2eGPynKVfB1j
RsI6vO2gxYi5HwQ3loNI7DgHds3JaQZdNKnAWjBCTJP9necsEgSuQhnqB8JuYUfM
orSWt+cL4g59Es9VdFBldn0m01W+vB44iHZgf8v6BDlR1GS6ijhNByn3eMw1imHb
IxuQSCJTidYXqP4S99v/h5SB9zYCAqDVfrhZNJsE3EEUsfDOLLLnQCov5hnggDZo
pGSDV67yXUVdxgcQJKyeOpAZdZi3IW1QdE0mCVjb2kp9mJdq9bsyLY3hlzvKQlNo
OUPd5NZsVVvDAtueTSjHPQAZEVVPx1/kQV956l5HVq2Pb2ROmiOlAXSROfIJ1tBd
LcNw6iTvJrCt7a0FOwCj0eMTuxi/TOdCG3prBBD92ylVx/UHpDGWO20TasUEeZ1f
8TzSd6LrE1FpntRTGOnpoqUEH/Viu0BrvIxhVAC+bID+wC2WIASz47gbHxcI6UMH
vJXyP6yUfDVUuIxJ18TVOzhxY9iRKoy+5Gzrox8BK6nWKWbCFsy1VPXFXSKCOpLN
908a9DkWaAhm9/z37hnwgeo8D3F5uhx5qlQAOrfSQyNEqw9Ds83ac0n1XvNg7t4b
itz8UjR0bDOhJ4WuXz4p6M5lXPXb0rFM1yUJbXUIIq7YGeEeFQnj4nAGwB3f9+VL
XYVsmEfa4QoUcgk+BvCLJvdNYm6nuAeKa0wqMPrC4JHwSFNv0D3KyL58tdqrvdzi
uLZWumXq3iLkitagD67ho+wllyrq58rsKpDEKvM6YRFNPtqOKxG8uOltICHp8Dte
P8psmeZ3klBAVw5D7EBz8gzkICUErzB7QN/QB+whJFbzpAMjkAZjd1qUUxwDChys
HzWZQifTF0IsEP6a2qT3K2+cdvezT3HuNwJGFWI7zVCoXLDpz900mao1YO4KC/Le
xwWQ9JrowXh4u4pNiq4qOMiItxCFTm9t2GjasSZDBPzqRKCGcvh3MDp6VgvS8azR
mvilON94Y3gXBcNYh68zV4ku21g1BqBFRlzBgBrnpTL+/jYHyvl0ooaIY0tcgNo4
hNRSkYADRX2LXMTfBwlhbI5qahWCR+NH9YPh3DTgGCw7zIsyuyaaTU7iql8OdHWr
p65pKu01FNBfYej7knpqRgyYZLpFeq45mxjzUToT6JA1Y/4EZ5ltVdU5IEpiHPzU
IeKBKtrEuY//T2MgH2Dup8WjLki4v5oAqaKa0BqI53Z2HPfhp0ZkkVyqrwVon10y
7v5aiUtse5Rh3BTlx6EAuN8owrk52ThDQzawJaMzIdCJab61iE9UmJCwSEVC+MyU
6t9AVVTc3IN43d1ac1+V4v+iCVukRtP7LQ7qi2AJ5D+BEm2lHFQ5NP4vUjxtMrQL
IWW9EHCOzgfy5y/pyBQdssI6xSsazezt1Ec87tF7WCXKJB533yQSzYlmW53aPe/X
oH4ShSJ8gmKHgCSFCLAUvpK6dQJQ0LcMQjvfH9A/xzGYlw5A7fJQxSNg4QHi+uo1
T4+ByZ9sGsazGP+Gs/M5U53P79sQ1ARiUX0/Tlfz6QzoToD8/G9NzpKB6dgC542q
th/ZYfZTeFtkIjw86c13Svke4fIsJ7fpnYCdiz9QHMXKRkVRng8R+9KMOeUbQsVN
sw3wt1XrMLa40MPc3KVONdmVYDCacZuJtNr9I+NIp739tGl63XuyzEGdcDjrw5C/
5JNGaSFlHHOgS1WE8dw4iHNTWuz/T2j7dEfaBjrKc4TCVMJ+4mZ2X6hDiYJFxlQt
KcroA+JCyumafn5JYoI59V+2WlzxpXtfZX8VXORxlQgHB+VkSga0jegvmG7N+BWx
UH21J07mWLOnjoo51D2uZWjKv3lEfr+dW2Ajgr/ta1eJmTvZZn1/zJG5PvZ/8gYg
OMcfGw8RURJwtoo3dRNxr6cicWg2xInbAnAITZOatXX/dmGnGOPDsKYeruqXHnUc
IYj/VT7WvQZleNrMjnwxMtwER4+oTzHKNb5QECqsK6GEjj5MMUMJ5rKKAaXjk6Y1
Xywd6f9ur1aUeIbiKKhLrAn2WMmlTHhxlh2yV8m1SdtHnw3ny15qBEIg8zUvLUJ7
jJOcOtv48PnAMXebWJj4A7CufI4/l+vBeAWeKR+vwH+3WIIPZEDTnFBoKUKuVk/G
s26tQRAMRlt5w8ji1zQ2OFgYs3w51lhO/5MM26R90TXvDqDVwUeHXPyONylB1PzG
Q3f4NhwUM+dFXW6Lbp2Nz6ITVpNFKPlUeHD18QxzlSULWjNxcpLfVfv50ICw0EDk
0XNiHYhUQlmkqbdr32FJeI2tM8Zbhzjwh8fFa3hQWFEp7jLAKPdbl/SYRpaVSVnh
c+RkoNLqhhkYBNhPejZv2L7LLoRVc9vu3bXBkUzGkWXiqL+elVfFYj7Sa42eQiea
6/wybLOoHkCGU/HhMn6SaErR+lC5C0OOamLy/+FoGwqvmw0DCEpYAoVeMl9XCfVz
6Vpp3zKGAAVent7iTidbVT0tIF/Ewmsr6r9I/ah9ZqzDVm5N2RGvHbUJlEdhkotL
lALznImtHTGP+Bqg1VsgJ0YLkfmkrb/5GhN6RK5ylNss54+RltQ0/HNN6dJbliVq
HvsMMN51VM0QsgzeCL0U2DX/WLFilwtHRicKNXJ4khTykGCTYt58Wrn7n5xOMD7S
jYpWzQCs+FHwSZ+0RCAXXYzf/iRvMDykOLKm1FcAGHQ4EXhS3AftAjnzKHJH+eRf
uNfxtTleD1xLz5y43dUmjD92Yhwdl1mnEizERLX5hkAc/nORJkb2VxJ2HXAqeaQm
la/k4NHzuOEoMR2a6kc3CUYTntEMcvmfjWuweyb1e2xlBPAz7qRhNgpV0ZFGdOxS
ksKzXuWQudlRb6BKeNtdDds8Zd1gUzV5gxLnoKwgObFjQ1eP9fwaJQMDdV+GG2Nu
DZajJtkFyVETFGdwRTFHzdUPm+/ZoNLmUmqZ+t/D87mOoxASsVRmO0kmahOL+xpU
rXWthAgOu8a3ZkqMotrnYX9qxJmAOJJFgWE21BXr26SQwdYxJ8WbLPCSKqlQc5uy
EnswHqGjMP9ShE5DzARUB9Qew1gjjRa/qK+yAvaCGX3UGJTcFcfFesUvKEBQa3tM
/4PHRMkegVktUBXseaHMomFEiH02qTAc9jaqSz0MvKD3fv4Oq033NuuDS/putcsd
X3IGKU7hkYxeRhUCCDuj9rN288o3XXPuChZ6Ektf7R8lbpvCb9ysUXT+uaeleUJR
ogz4BvQFuJihfTI1urd/iCGHIOcD5ifzDEJIKQdtZ5HOWe1N5QkVEuzIoXI41iAY
RgXEUGVQyb85bIJBUFlXulZai21v4IEOkk2bABPPoL9zqaEHwvAGbBL7HBpHXst7
1x6OLV8634pkNjMbetkOt5U/YyK7N2Scf2E+md+FXMEk1oSiswOiRzqu7BtLMRXQ
FRYRbH7hryH4rygHt2l0dtGuShoDifsCxiHBfKS+9iYCP65eCgqEeXJ5kcY1v+wO
544YeJOJV/BKLf2wX7e8OoY+QhW8PNLi5bkadxejvBMeygE+s+1pii1rqcsiwgE7
5j1gZT4pLT7ZVmkuaNDPSOhgYzHwnMEACV2wCVBmn764PaSde2ngWTVLYbNGBRva
fy8I1rzHAEZ21rfr4eZe4BL/Hcz/TXrwMJguTZgOVfJSXgDINHirGcM/wC5lHOfL
cFGjtv5YPaZeIM+TlTZHriaMsCR2eYTrLm2w5O1E+Xkrd6saPRgiTVEBN1M5CdPh
xPPd9FhbKfohgLg/80QpJIIGHXM7SzudFjtoGklkTmygeJWJnfqvNXEu5lWE/xXY
qh6xWLqlMLjoQeyeUFLmVFOkXHyjsnSLXIQqMkisQPkolFupm+ykC61/oiCCE1ay
FdSQFvYVOucDUhqtlZb7S4/lFF134PvGXSw7FJBQmhoTHfwpJK5Jh/8W1gpPyNlB
h9blPVikQHOQ8a4UZuEWPHEyn3zfq/aiOpPJm2oqpGmEzW7vYDkVVladLQneYenD
yN2AIab6WX92W0kV6gg+NBErBI9HImHfKsw4Y+KwOKlB7OtPB3bgOw/6yXUjPCSj
UONX2mF9YKPm8OMpagbjVivmE7GjxTK2uM2G5uCbQV4gXgnkmpRDkHXzyJvoJdZv
3MtXydiP49pJNbRouj02CEkjRd68eruClAmMpfXdXR7OycF8HPOedkBMkoJVn79H
3s9eb4lLkLW9ufpZRTGR2S7xxm6s//cfUdignZpJqiR+Z60oXEEFDJedy2BfNTnX
L+AoQ9gRUk/bsd78FkJLEo+pt3rzmuLLkxAQmjCNZWZAfvrWKK1zE1+WYk9jEHlq
wVcURKKjsgPLn0DxWzZwgGYGllEEm/PThRMn+CJEpzQ5Z+N6tY6PvXHdaJOoIYAg
eZgmc4s1S1k0z663MB54VvVgoHe4oc8UfBBSCGwI3Qy/IznzWPDqc4Rx2rDyDZOJ
d9AU28LvSpaXxE3GpXiq9a8NzBOjrJYbxHBoR5zUVb1iHkoq3i2Uq86JbETu+o7g
jImU2/x6z0FhdL0ACLDp5RvJ1TjG7SosposJB06dItsZsbWXERkOhUBxCUDSejN5
GKOZ/ZDUxzPZFzrqP7T2BCuP3716SH20zKNiqhY7DUxfjunlL/2b8Shqg4RMi82t
KgEZ9RSC0WjL1knkzu6csZhqvIukM4PLQZpMCK05mA2WhWUrvNZ1ad54igM2dgEw
3Pi6RGqzsbMBSUG7n7PZNE1BAkikkRCJYazQowl4iyQOR7XtMeuC0Rnz2uMc3bwV
r+8JvrenjtltXLHPbsszIE0VA/CsIdh5owh96qI05ke22uHU6Ff9l/74avdHPhQi
i3z1eQpNgx9ztzk8AjMY42tKW7k1heIepYopONrsVfR1P2WEgil70F/REI/OUv1K
tuJqeL2RTFmambBcmwMLvN5smEM1ejnDKzI1417IVHnbFxMT+PBUuD8FRfIu+stJ
93niaLF3h1330PJGNlA+JO9ihd465VOA9/wzAWbyG0pWgOyCZG+nflshpTztDgY/
F+UTWphs92Q6yGhofGBFr9J6bo7G2wDabTd2f5+Ldoj2SGZ7vZesE2FNpNVJfmD8
J9OZxfKgdoQKIwogzZQZEHqILrgYUcbLuPXBBQgTs3wKA7iTqK9VuZb08pwKW/Jk
rawDn0ZessvVMJKee+PrkPmcW49jAdTxEVz2VSKNfek4KlmcelJHfFjGvUvxjpwF
DqfRD/t2pUr9RPjvYsH+riFCm8dfA9mAkENiEa6gco+rEpUoaNVEt27nbUfEgPJ9
h3pAOtHoLKMe8zoH4M2AfNnBKvl7e2S6JaC60xBOJn5W2J+lSjZcLata0R4i7tbV
lne0yYySSq9Z08AOUSAoRjybl4K8ANFKTRuh6AWr2Hi6O+GjHusH2sBQF0NJWOpx
M3EY73bSh5H9H2moT0eXMk39tJPIm6ZcsdrTVVPwIoBmSV0yvzYFUWlxr39DopI9
FAoE5GvGH4AIGWaulMSwk7wOTnMXXSrluCDqBH1NEDJDPbQP9fFpbUfs6CBk3Hrz
K2A4a46MKEauYXWf8K8BKsqath33ORpP0fwG+6H5MSj3uf1VSzvVEBrYD7PFO229
VTK9Vp/P/JzzQdToQu9lo3sWK8zzk6ft9D+6ou5PyVh2FT0e1bFbVrLk20A8BLV/
9fNg9ZU9zsI0tHKFypjDmcQLYKOXCPuQJlVQiuoAmAaleqG8UhKex2BM1DcRsgwC
WGruWIjZhKSQ833H3lSAK55HX6ILExfJC95EiGj2teawA5fw2NFyPQq+XsDD7BS4
1aUaGaNu0gwsl0bk7pXeaSL9MnYQt2kCZBfbzY5oA9ii8dtlYtGdPB5Pmo0SCoRD
IWFTy85YlUsn/09rWRx6vMV6ZA1TQyO5hzgNKcU0ibsjB68CfPxq8nNrIJtPiT2h
6dJ4dRdW8a1accFu/KzlYz8xVFvq1rB2e0JzyaUvITrxCLT4k2PI/bPkYb1OatQb
Zvt9vWkecxz8T1497nfEQE5YqKvxe4kecUnTdg7CDmutfuzgniuDNRpOwz5T3JXQ
wUzRttbgZB+4IZctsJMNsJVltSswNzG8A6FG0YkNMrq8C9YOsYSJE/5V9XXD2Qkr
VaOH6eYUWKuhH7ye7kBncdWbLMcSUvnuaBhtcS+APZnQ+sm59HmhJk0ncIp/lfcx
wAGu0vRVU4kNFiCuOdRfs0J04UL10DLoxQzXSk8salbn/+EMATSoWZLR3Jz6VmIB
nNFUpDxGQ6Bj+4B0nkyRnD6NvHHbnh6chYzCGg27Av1JB2oS1oh0+lfwjvgVksXZ
NCXg//Jv4Ly4ByERM9IuiHQ7LFyMVf/wgBvHyH9a4+5H1Th5Rh93VQauv7L1hbr8
Jj8NxlKMxW3mHBG82Z4ggdjxR0FkAlK0Ba3I5FoUOkcq9zlqNsMpi63mX7Jy3V1k
w+w8OLEMCJENuIJfK2AVq/dOjBL3p1jaIVHNY0Z+cV+0Lk7GCPf2DF7trAk6TBw0
M38w5dLHBTjKdC9Z3utM5/ow9LvFWIEhzeOccR9wi+Az+T5WxLKvSDoORe0PVaC5
0/46qGRrMD6CcOA9ZBj061N2SY+ZlhElCM3DO541pkeG6CTBsVm1EZR4mP1hCCl8
AScJR5gOk3Qr7aIyyBXRDloLVB0CNLexVnv+ARI8qjUWUNvWWRRQDhucEqzsewiG
Xogzvtrf4vlkGKsepM0anF1LPUQwxQbZVNv/j6ATakDdt4389+zgq63SI+tHNn/z
/MZaPlNi2h4n32Wfmal7aAe2EGo7bfteCkXEtTrSnfyVdKOYZQkTjpubaxl3kSuh
x4D8cPUfRKu15eb/8mvc8fwIJ4iHla44SujApmf2b7xsR14fPNBux65pEN3oiYqg
lbzK5Hc8YuNL6cNxQUqilIefnu4Tl2qaFdbmePq73z+61IwUjAF9GjADs4Y0MjtO
Ch4etmS++BJ+7NWDeI0t5mS0lTs40LEMA/ap1YebTXV1H0ex/NFlShAle+Lu3M1+
kPSuBa0UMozzhFpXs8Qonee2EgKaC+QdtX2WkCuy1QPKmu34dh15Ad2limmLh8jh
EbMh63ZqsV+GVtB1N2kxdzUK9XGs+ARHnQXRIjir1E58xT1PCEfn4BraybLYC39a
21aprbNXCWvr5V46ec+Qd5pm+Q3MClcoThp8D4LP6qKcN3je35hit1IHJ5d3YKNT
gLmWZsTMugwliQ7QBqKrWt0gwU8ftIImMCmUyzVN2F+KIBWNxEHwN7tg10coyx2o
ZRrcul+n67ZI7Z4RajJP4Rl2Va7GopWxi66io4cVT6eX1BeVyDkp528BIo3bIPMM
t9NKbvri8Dirrf87cnLC5KOk/bq0mErk0pSv0oAw/PyYpxFQ7ZD7LJXyTe13layY
HSGXiVXEzUehHfh0QNrRgLS/zhxmXJQcZyzi03qm/qJymqry7WcZVU42AAUAkcno
8TexWpmEerxLZFwbAK9ltde/aFvlW23ObUPHbRJxnxTn7uUziy9XpH9vByzsflHH
n1Jij/of5/W6TxcdetGUdR1RMtaEWKfokq2E8wAntVQOq1KBXdfNi4Jm5Vy6eYvJ
mNBzhD3/YigoBmRnLPZdls8WkZBaOYtgnVh4HDPtkiWdde+wRnBsHAzmvouYFACh
zAR9QLwjEO27UvIqdQTsMqYvFxCtX13AJR6frIzviOXT78on8gThacMyjW6xI/GR
Npz9SUMKv2GTSuuWaZb0KWTQ6tYUp6mtpReRrhwOmmEOmUKzyHkfx7SybhAfKeE3
KxwlwBoQ86To4lgQgr5C++w2pFPLGvM2tLoRrCnhV3nvuNEg1EE4hBMQVZQr6yoo
ysGSkQVzDet/FUQWzEI6MD/2Ub74x5+vqiNenVTr4UqgEmIgWdxyV1a4OqKglCa3
lL+ffkSxJgSXape3eqo9eID/bCHRqbJRXgAi/DwGkuh0MYvqCk8DzE4liKGe6Jco
5QtCzKYi0KIIF0bjGh6Onz/7hdkwbgJN6QZyNgX7R2m74TM2ikZjQ1AAG/4ORZsz
cjATxcm1Be8M54EOsrqRvBYwvV89BS/qwRnak3fAtcI+w0XjfuCAVf7LcWt7COgm
383nvKEX48jg4XsR44lWa2pSjt0ejc30x35OL3jokJEujqQnXpYGOR1R7PiZYAaP
jLxFBpLWLvN2cbB61PuN5uEd7IewEMjET3C8hHss7lPkiqRdGKembtAgnqb1aeJj
IWlBrxYUsj6AZyovVOFXWepUJ2nTmHMmssdmTT186dalBsCPcTUzklEitXZe80ed
/flZOqd+5DvxCZoNxcHLt72/fAI1E0RsMYRniemGQZQatRs6+13gsYelEReq9PwQ
Ii5e6hEuk3w2SbuQ2yi/RSLW2eOOGZ/L9f34ttXX5FDHTfmmQTFYdA0PcYTllU7X
ZOlLgLh2nIy2wQU2h5FyekBc1vzqmgaqFA977jcxWzd4tCQk/+TXYc/JXyuKfBq9
XrqGRDPpGZ5kQwSZHNjlfgLlKCgmaMrY/y2Lq5tp3E4JUqRmb0rB3efmdG3K9Qqc
3Cn4YS/zB32bRXScWX6q0R/+QxmlhPZzX40cbAeVPuekdotW94fu7BN2c9l123Pi
oRHepBo05Jq41ykp3A1NtYNFq48QyfYdM4pBpYGhAy93bpPqvro6jgi3/z1d+5DR
Z3ZHpAvNpApd12uDc+k7j9s/kX9j1UuxCuXCjq9XUE5DfVLIyp+LxbsqP3pwU5pP
MDJJcDr6o0TbwHhSVKaCydq65nISKccKlNdiHQBGHAt3Z5i4u0rMFw0yRX1GCPeE
XBlvl6YLFYmsOVl56nnoC3Ue0FdmKNz8vxrsyMLsjU4rvZdj5SiuXACmyGhgtWSt
qhNR1ZSu8CSh3WqSZEoKTgrojm+3TdSsTPE71V2+g/Bmhn0uv94Fd+zi3ToFOY3x
abX42dmW4atLaWZiDoqa3Q4Y1qUpx+t3OKZChHX6W6rmlgtNIFfZiMrRQ5oqtkYJ
AWj+CEB5iuPswpnTRJx5j0bwU++WHZ66ewHB79dMnbgk8F9k+tfFZwBB7hqqVcfU
OC+KPm/A5cb78PSik2+tsL4nomPWJ9W6VX/aJLQqpceS5k8dzUCU7ZGjobdZGn4M
zfd0V9wddqY7nbGHQ6dm6AEJopB+S7b7ubqffoz1isRrLDlIZAz0vtzBaRq30aKx
hxqfuLKzq+IcEp/CMFQWEEt3/+7OnxKSEa2tLe+elgrkbA7lYmT4bWkBDRKj94Nu
lVtpLMie5xcThU6IIdpA4QWJbl1bDvdTGjOdn9KRew4P86Bttd+G0y/5e63V+syP
5Yzpfd6Sv6FvmvHF9/GBii1H7hhr8BqMe4xbu4uKmP0QkKywEzUe5zQe5eH7u+oi
SqesWB99PwM59AghRP7SjCetycUFUpni1FzUHU4lCIedg7jhAO9mYJWwIX/eF2Da
DD3YzsvAxmmwSD2gJri3mmt5iOqtS0FyTPos88VulvyZm+fuaVAL/UuRurIzKqlw
w3xfvCbPpA7iOZG5MYgjFziihEvKiHOt0uddvZ0T7ZEKCLI1bnYo3dYAqHu+QR7W
Gnd8JHvMJtXYl930P5Uyc9RI3WZFahsmtRMNCdjL5S2ZXWzvCG06oh7mMLfEwodO
k2Ai8TfX+4c8fG+dNYr/v/nzRETkY/Ih6eHBZpL/f/LknpAxw7T5INcDS8DKqsT0
X3iLPgVz6jidL7YlqQm4Budsvm4wy8aWA8NXXMgSMGrodZLM7+D+RRWe77S+5k1j
U1Jr6bYPCaRoux2mHYw899+rCxhx+J6/HM6Gzaj7SU10L/qRvy1rXfBbGa2MamT/
yW3m+HoQYdGgHW6pz+msQxwU/At6dWfPZUO4FwQ7fOAUDgTZA/pUgguZGqBUrA1L
WniTGaRapRdf7s9vTjU+iyYU45oSP6lMMaqZ7NQ2k2IdyZ67wpwSWYjKyRlA6lJu
1opaRxWbPnzXGA6oM/LqAlzMj54vrRkqjoJPTwfqTAiiIPnDOKtqFKuroJimtjnh
ZXnek9Vpdwic+pw9BopRKTfax3mz2q3U3atM85zde2JTjRbw1ZsC9iJG/uNi+xLB
+7Kn/9EQVYNUBzb+FMi+olTDllGQkQs1qJ/Gm81pKZ+jICyBA7/dhjnJ8JVSQo84
JDVEX/XwnWm9/WXkddm8tpAi2kSc1ZFexrskC6zq8iqNWcw7U6yFFH5owYleH7gr
M6Ygmaajkgs5oKsLnldu8u2C+eIOtYoOkOTtYw7i7vk17+RLmXu3ThObOtGOI71h
Lnv9KrcA9IHPBG2UOnT+J7rNntuDvdqbeTyC+fcHvMZg328PF5oHtwe1CqVaAeSN
XiOUVxerfQ4v86occYV6xtDyLvhblTdHrTUHmaiSlUe8jDfpdEpaGhmDg8/h87p4
hJaT0k7ZslFnrpcaEwb0/rx35hXa26YzpbmbfLvO2fbMKTfiJ8UKlcmEDrhWcDhr
kGS5WK1LUCll1iUNzfk/atSiuR3prUy+joBy33//+Ml7VxgzFaONg89JYwvXjqMi
v/0bZrTf+lQ7sJBDXeoR/tjZCbV5Pz8tJbUGid+78eUjiohtKZSfr5w9nTI0aVov
U5+BJB08KzMydjUissQ9mnQSOqphQKHMHFHTaoj9aIpjW+tKGgqNRvAAMwZ97M45
ogkcQVPIVgRRR0Q+afs5Bk28J615HCHBAmc6oM6eU61oC3N8vdDbPHe98eVew5mS
CE3pKXuXYbCRwGZfS4lyPu3JJogyGALAvuBUXKoe1o1ek4eVcWij7DiQrowFQVCg
Etco2iQ1piP6CLzLUT4+Tjt4CbfwfTJwiEVz7F82c7PZxQIlcT0zgHZQp4OKTqj0
xa0sOl8hB3bHoZPwbKAx5ec5JcyaRzbae6lj9mYIedWBnUDjc7dkgHkcOknc4XGV
5rF3cNsNTVNmtq1Nb9SYEZN3jjhteUPiv3OH7A19sRqCo1iZmgVxS9g85Zz1t6y8
nJRaf5G+bMsaSZZWgwZDpBTLOpJ2l1g/Hq2iPS9cPu3k2AdM9wkGtAAoS5r7HLDF
MzRY0EsRJfNeR6ifgl0Gcvk7/bJhsfyK/bREXi5BCdV/ofWOM8pMbq+T1+f2pFPo
r1fTsoog3nr1KRHJutk0gWHYYu0wiKkAw1y1e9n+OQ+zZaWvUB1XLyqag7g6ZP3l
91QTs2IJwa303gHyep0/qr/eQj9kO3ybhYifUloDj7hhReyQbn5YGL6yf1KnXU6k
3/LfDaG666Gc4llzpVxEz6czADs+4f/WYDTugS8nd+RThrrZCXBm5Y6eWhvvAFzJ
4qdXOHCVxljLKTx0s7fMGrp3rkLqY36GWFIWujpkm7rfi8u14008PZ3wwTDg8V1E
hTx3lXHPr1AM3HTgoO5AYCsi5KU2ush6JMDm8dwIHv4TE1Fae/UrZbIbEM9wwIMy
CcfLFFhh/Uqc7e22AX+OSmp7JxpCvNsCpVwc5vzctn5iVg/XBG7dxthZu8T7yc2Q
FCr9/4zVdt2xhppxMYTVBTao9uotQhcUJIqXh7DllYrkFB3738SdUmJb+56jQZKC
ZpVaIJDJdVqMtnu30lbg6K3yRURgfPWivi8emTmq65wJIrIjB8NEZFVFzKhrBF7d
7sAzmqVp+/jwHsgu/HNn4i7NPGu7fupB41xxPtbxhjY8gF7nMb2fi0z1DATyX2jN
kopxXwx7oin3sZI+BqSe/Q3+HpZ/ik5pMCBzUbleJZYCSAjklMYlWKrVlDLwsdS3
eR5j6FzEsOUslVESbDI0gTMjRo5ZT9P0gCCpBez47ztPqDkwGwbZypYwM3PjWP5a
VFYyi5NG+I+fdoKlA96A14EF9rtTMcfBWxfrqDNNi1VR9zfgyGJRIRM1h0xPiHF+
Q3xXjIuihDxBA3IAJECSCtgGNWcc1Klav5/y47+0oHHsVW8J2VJHSKvDDYImK0rP
qMVbzBPVavFEUvjZftDic+zi/ES0CNTqxqNK0IphbSPlvAQejFO4enoEUs/ieGuW
RJjoPOX/zniLCAf/FjTrJV3ko7ULWvcjSzLvme2Lj92dmDYd5CI7/2+qnQWMNh+v
TTUF85iSohMDMMfCBebUqgkX+uV7c7x6c2TeoMmphHPk+Sh/LexBKozxOfCHBEU+
RXDnwgvOBkVTUE6ZrluIDS4ASGNse21I5exawM5ukFQzEu2mNpnkH/vQoaD9MxX/
tHjfVFOJX883jQgOOLLpriadGXSS67rotOVhj5wYWXjGH0Ris9J13GOwhxMjTqaU
oCXC1685fHok8bWVhDqumud/65rcQH8+GzLGBDTZUhTBeuhyc0EQKRGK3Ujnovlz
VWEVe6a5XuDhCzPAdGOPw5Xcgr8lQmP8qdMD3VMFhb867J+cIthhLgMqp2yD74Rj
5WhhMeXlGFpFeOg8Krd1kBYKTZOFDHpY8PJfPOldHIu50tNMClWXy4CpUTO24zRe
DDcbyWz5S1IxP1nxz847EQGbVzlFxqBuqFnoYe9mjdx1I+VnIcS/XwKXpuN3CawC
GNQybt7oX8bJrMjSfSHG1qsQ6FPRl+U7udOEKLkeVAmXWQkgt1dXU3gaS3Ygv+HQ
/RANZ5qcktLAIHz1+4Gpy8cQGc5egeEh7DUPHendSP47gwEGPJnaEztjVIlsyyNt
blYTUgwtSakiYH4zvy3QluOoTsh2RYwfflluipcz0rTCXfSVD5Ne4F0mYopx32ko
EsnB/6mhJ6GmXjBDuBIBSAnh27iykxMAMltN2WdhW1R1jUC/Ear0dPEkcV22Qx3b
7AVUW7CnIQiWctIBwSgojCatDQ7VPpR43XpJrjO6l69j5lvzsGTGp2mKTkDqlaCv
pUF1Pz3Tl1qUVRox27c8dw6Q0fwzw1eteI+KUmQrTebuwLxJVh7R/9y47wRRERIo
W8CKUg2BM5OV4L589WnWsEz5ngNzckVw5GudIPHN+UoCyGKBC6nVfa/vVZB8gyuF
SQ/meCFOI7OF5FdgRb7eEOtC7WPl4B2YhAquOA5RbfQ9gcJPc2+R8TyNKxXAv0/G
bKjVFhTg19c8iM/PqAq5Ffp2b0Zdao66sGLyPIWM0+lezDBwrFxzAD0G2XkMAUbU
RjC3bpAcXD+xwpD9IqETE6Ey+mO3EYJ+wMIELqsyO+VfJ5gv1VFssRBIdvfcgaPd
ji/zOucvVnavBl36D3E80s4TB7V5z/cbZHujvfafbf7+5c/krHga0mAP7ydiO0cA
iSkWZQa7wdz5lmxMxgcYbOMGlRxmJiVVKoBEIC/DVOIqCNiLyCMrUrOMjfdMMKNr
cc9TnrcIWj7S0aVzNxTXxy02C/XcAO3v2o84DwnSFZ5UaRd0VWoYZvO0rYJDXmNJ
CgM8ibz+Bxgt8qrGUm7UDdhDSosDagIfrT5PeiOyZZpKvpYMjn/GlRen5nG939Oc
4RcxBppEtU07e9tArQrN/L75XOkI8SR8nlBFOkXWas551O0aZkcP11C71cUnZv+/
S4V5eC4G1ZA1VQrvEkPn22lK6mejlJGq9DqNs5mhydl47Jpro0kXb3Z+3jrLo0tC
VKleHDL+5FTn0Qlxr0zf0HFYgv9aukQSlcEJvlQsDKeMxykuwN0HCsIn+N9Ox8Au
wq6UAzmm0P29jLAUP1kQW4j42alZ0e+5cDETiAV3MYQLoO0aSBPDfYtTru33VAjt
DJSRmF9A1ELAdy33YqS2p6XTNacfuW3mizAAPXNsTvFdRUJ2Ud3CJ30neG9D9QIs
tGOdFyvvFcmPD1VY9k3fzqRnHSzJha7pFsuaE2nf4TGah7bwsgaakVnKG0UytguC
DWex8Mdp1RJKv19BLPzqaogLA5zVg+lUeMWFQQt+qNLDB8DCiBuNFQh770StmakM
lkrUYaOoE6wvCfFd2ng9OVyvrId0oAqXKJQqS3Q30SpzEjU/UGvmCMbCjSRRZN2u
757Ozbl1tZEtKCRIm++Md9tYgwSMeV6NYjMkeiw9WJLnR41Fz0JYvdugrmSADvS3
i0lPC5WLPK7kuuQBE4MHv6AMsj4/igxyqf1ftXmH7cA82RSJMI0NDM/oGbjrWvQp
Il7Neq0pQVK0MPvcwV7bn1GiAQ/iV+henR0d7usj154FG6t/ECqsqOqdEro45DGx
ZCiwPqFBpMsa3/c8AJryVma1KtI5MXHAvTWGA261TwC/VST9wN0lvBTGiBjPYoZ+
mJLX6bWR7aLmw/lv+YNbBmQs/WJsIEBdM3MUEPmof+hsy/UQ5xg1hRg+tgMK2J17
mLSpXdDIcDu26BPDdr+tFoozqSkzStE6tbr+/60RtH9bGgQyUGrjhXbkQUf1aHQL
U09joExqzYhVePZTa2O7cYatpFOMmdukitsSt5z1Ze35MIjugt2kA4Zo/WbxbdX2
BItwxuoTe+8vMIA1UeFPllkaoSZInGSGjjxpXoNWtCP+zLY3toM3tiAakqehtFrQ
jgdivrVSFQSmLve/1JDiv9hNHOkze+BEgwVGRGoIEmJe2S5EVtiiwmaSSkWYXPL+
5g/xM/GOiqEFk1lRS9q7k8urI2nDlpzmEcKOWQeYu8nOiCZjhuu+4FReiOwwzNYz
vgREyw59m2UOM9mq5Cv/c3WgngGCLYuS1ZxWM+gIkZWhclvnQO8Y9E5d+fn9rZrc
CiYz+3aJ9voLMoKndR/NBQ7YMH3XmJHDBHZPXT3gAzl6QDrXle99IDeoHXunt+D9
J1d1tnz44zJps43LDRjl4sXdCWqIgd1rc7jx3lqvmxrNQshArd2+wV8RvenAUo2r
zkFOGXGtOqoV60Y0JbZjHkamS6fwKCOFCNgzpPIc9fs0GhTyn2coLcUPfOBsfCLx
idJMcA7W3n4aJdhbvBZlneIbEaa46kB1YwOTyPqLxcp3E8+n1Db3sR17aSKvXyCb
sQPOzWKcRK2PaH3Ai5sa5w+RKhUi10OicT3/eUecejEqsiWUuFgabsShMjKpuzTs
rhKPcTqSkh5KHrnk1aWqStdQ09rKUsFlNRHdUs69mh+dJeG734osubV/2HebsXa5
BLFAmZmo5zdC5HES3lRHWyu23vhpejuqVpRVxnmXNH/9jbSPl52IUmkeKkTSWUsX
nmFXGcVJQES/pP6vZ4xmW2gT8fkpvqej3EDTZbXQxA1QaBMEAIlwvXuNq3PLpNnJ
sUQt9djX6fHjP7o/YVW/KU9GwnhvM6tcNVHMTr7oGvfEkDHRP2pEeswJtD6EH488
qhodv9hDp7Oj/PM4U30YYcfNYyivY9PP5r2rZ8JDzVW9xjj0xhTzcqPlyAmwPu6O
LLPDx/s6fXGF9WdhkWY09KHulR7ueUpsmsMFdb0lg9Quil8eqjIQChVV8Wsch0Tv
o80gDiIhLZme6kPlfOXi9Ds0iIECWP7JWIIM7trGDQqptY6rwliAJ9V6g9qqv/lm
IzXn9uGUkfP1bAP6DgJZV/jQXrGb9KitO2By8gFn5IKTZ1Q8EYBOX+eDfb+KXCtB
5cp+xgi8C8I4W3ClBx4c4La5YqyVFiKmYDpwH5hORBkm0CTE/EouX7snMDRZTyYo
p2whBRKC+eujt99IMaAmwIxemmINZ8jrnw0M5R+ogrr9+nHEtCeaCO/j5iKZJcia
oYJhb7fQIWxo4qPtsiCpNOJfZGfg5noipdkyQ/woHnaTJJ35pPYX46zNu+lOO32q
P7fBxbmOAJtaPM2xwmCXbb/8iuQEC/ISMmWAjYRBm6UX0moHYRWxRjZCUdaY7ot7
9K11jGRmfonZCvywWtzplobFlxH+jw7/3u3g3zvdG5s3dxhfm569QMu5WUrC1549
RNY9qM80S6+1s7RqTP8eNTg2Q6WTiICrxIM6Jsd39hFXE6DPIr42llNHVUJxxFYl
NNk90XXbPo4TX21Mib/sLDkHP3tlgyP6vsA3HPbcd795XmWTaDDQM/n50cJ5xDqa
GymLVh+y8GLf8VQPvwymCdOjm/ktdDszomP0QRLtAcpscIPVt/rXBoQl3EazhxPf
xqi+TRtT+S7COfOJIzK/PFt6x3RWMaN87kywWrFrWCUd3taplQTSTflt6PkiXflm
xRvlatnU0OogotdZbwtea510tHKcL8bvVmA78NUSDxEEy+T6mrUEw1yDXo4TSaqf
FDrziaGhxqH5T/vw50okZmtBtP5HX88LeRw8sJYDwn4h/0svgDgeo6dWRRY1Yn6y
e9Sd4TU6RlWAc0E3uSXG9E0C90SPrjnMWObS6dq8Qh8kKT/R+sqJ1QdO3vn6R2d0
n1dfRkAGrzJnz5MRpZJXZJVjVlqoaQ4ajH4eZU/BHZC7kxdS8ypNVaK2sBI50JRu
To0At8KFpBWbp5J2SAp2zKBA+dDYKQ6B3cGGW1J75VpQgGeV2MuNGdiDzuDGLUDY
Ywh23krWn4DdpawAK3Q/NE0Z9kwo3BrI6Qy19tHCaO9tILXISJToI7QnwCGLakxM
J1B/YGb3Pq20PVbH+CwVnNv02aTLD3oew02buNFzXe63q5znraS8CwkW6Q6TXSXN
Bc6Wgqx0P/pfrk1DkS+k/VMS1VQKiWbE56ZKAizn1GU8eMm0JJ44yzdvgX8mrTlv
4mOV7fR4vALZX+eSYCxatV6xeDVwA+uJyA/Oy64wz/c5/Rwm9qMV0ykiKQGKYLLa
wrmCKUJXRqcgGmgNnvsUDHZd+BragjTcrV5T4fSTghyF6Az5tcqfBcdfsz78MMob
q/mRrvlTqMEc9wDcO66pq3iNyxeDH8ZnjU13UMqRaah48N3C+irwIh+aYGhgv5YB
TPyxqyRW6B04JIyYFft/MN6uHZjjg0DffyhzzmacnjceOc743KP0oYekTjI3qTcx
sNSH/87VcK7C3NH7mZncYSdO2f9uEdr32oSCuVfTe57rUtqvlD3arm1lNT5294p/
hsZFdVrE8LEAmI0565mbnFG/ZJSWen/V+YR/5sJfyPg2gVgjdfmlhR3qxC+Jb1PQ
+Ce7A7wqTB6OlP8L6qTBPUrfWgxfQEfSJY7SJUGBe5IYuy18ijyg4mbKmhc2jx5E
kR7VV2BhIiCLeLJGMCQfiKDU4y6CD07qslc0I3znYgbRZwMz/E154EDzbPplsfeP
bs3UHeqGA3zNF1yg1hgL3qrO3ZVPYNIFRLRfat5CZE5V/uCvSMx2zeDnywcoCw1D
qO3CDZs8JlCmgVIfLJGOBZJXzeK4pi23sZzk6v6vZoKADoUjiJNm9d6wGL0c+00x
mi7TVNr6cjShX4VtVUn3OLExA1bRw18wd/Vry6sqneg8hDUZyukd5jl1P9zgUtxS
bA1SormWGSqlUhoBMmnf3nEx2nbqxZhYZ++u5dXI97E5rupjC8DIKADqc/c4v/Es
QUhmuDjM3R/ZbE9gGrEKJOqVLn/p1GDvsTqpIUhXP/J/OCfN4U/dHtCqbC/JxRU7
UxatFUZ4v0Wt1e8AWoofd1LfsELJz/t0XB/Cm3umAV/VRz9sUhoo0R08fzNpwWvH
DUUNjVTD8FoacwE9/sJMjd7FVtblEuONNLlikj6uQ8T+ez9rkdn+GoRZEl9PJbVc
zGpYsMHiG2V8j+29ER7cY9BgTqMTd+ERoc5YBSUtL0Pw2YqG8M2xXL11lLHsNcZR
nLEsfn5Ssso5+mEIPOQucFsaTST1ptehpMryEFH7rGCdJzrdNCaqly3/6QGIIpE4
am/+ojSiSe9nxBepS9yWJuVzp/N4IHoO0WBAE7OmIbUU2fvEqt37LiFLLEVPhyOG
uJHrIZcWnuKJKfos46GBxpKT1kPFfZquJxSmQSjnmGrzAUu5PuK9ha+DYixSKU6K
Wgga4hfZCx0p4QbaVK97oVAzswYdHl249UUs4PvaKkvGkzMMDIXdpuF9nBZ6prCK
As7SEQKk+k0C0HVWDSu/jqzy3Vxsw5LmTww+9OCuBc/dv8UzAn0PZtA7ICPaOkSf
el9ZK6zY4OV2x9rmG8xMKXrdmp4qUktizMLKniKMmq3RzEp0M+7bwXGxYY3HAPO1
o4DJlxkbLROYwEt+PEmLnfrGRKRY7COjdgtocaVcaK1aGsnAeL4XIHicuxqo0mta
yHJkguB8AHXqwSxROxeXWhVcKLjUlJWLS+b+WBnVeupNp70XyQm5slotQr7TXYeG
eysiHG4hlDLBGrY2xh1Hq4pI/bcCJP4mczPRLUkVUVR0LRa7eopQ3zPmg1BBPn3s
/KKpB1ckkA4j1/T8cH5bW8/AuawT6TFMRsYwKYx6n+kbO097mg5CyWJuMg+e29Uc
hv1qEIrvPr3rViQaQt30jslSsqC27m3fKYlMctJ0TTvcK0VA/CooCyJi7cU1Ngd2
PpfkroIkcPxuuJUg29CqggTFDLYwusbZEmn6zdMq18fP7oZU5SAZscu/etrZYyou
8+gNSkwCPawJxx5/DG5tubXOtlPGqpRzAsVPn4QxucJ1wxaJH2XhzyzBWgo7xAo8
bKbZAUk+EAb+eWLZ4r5N88oCuy9wmCneuLcwCk/u47EGGNNpMMLYPF1+co1ibqOp
JEjM97fn1jSpd9Tf3iwcZ76IuceCg07wTRc259EnGKYZERDr9kZXMrpgJoBF6USD
ebPlF7XVoHYEb2s6XOAYAkn9V7KRYugmGgCNzBa98c39qPWq8WejRgR2VfX5fVWm
9KnCnKC7bXEKSM1RVkVVNGe0dyrQwpJ44DUrRgPtM4TQt4cCBpyQaLVVxuHKsP/R
/QRRl/R15LUkDnmugWmzR4Imoi/A+5m9oHSRega3GGKkqvN/VTEIgRKfbSMsNFcX
UyYscrhlfNZD5irnLmd4S1WeZ5bLzO3UPWFh2rZgKA3uYhoAJWQ4ifQVnc6EwKbG
UsdY1oKqc6EkJr9T2tXQvw22kCMpbznarLWK9jnyE/6cSxWTH/7xvpsE4AuPoaxH
AnCICNVuHBHtj6TYvuuM3ulfBiHRJsZhqsX/lr8q1jicJrBDlwbVSXdJMBtwyjo9
US64f1DaJD6I8pAZ1DCHpXGIJ3YTOq2WNp4xlaVNrRjRz0nPMAYhaozSqVQ9APEG
uQQCjwtKecqwvoAYOKqpaFpRlPfDKSMJWuOw9wW+l+mVQaqm6eU7vwDoFF+xO2GE
BWlV1g4pQKuUqrc5YhAcx4VfiSkwM5Z/2300dkbu+GO9z5Rx7m1xcQcqnTvfB9ik
273hIaKRUxZAEIuzMNYxLt3F5CMx/zGq5Gdv3fWUdx6Nu9O80XPjU6E2uK/fm4QD
mCGM+x2jbBloRye11+bdKi2+e01zZFti6oct3Utoql5PSINV0uDiODhMjjgA3pIZ
TlFnJyt9dPC5tH5JaGN1UWJrqJMslO9B5yqfS4WdPVfDzl0A6ZMlIauQaW7HLxbz
LZ3CGmBgHVk5v/jXcFxjmYd6LWvdU7KOewtetUE5NoNmAWIkAW5iuhlcXPe3fUyQ
x3FTmxbE0DtxJ6w8JI7tfbdD3nTRc0NOozSF1UQ2kbzlhPAplO530AMK8Abs3Ebn
yF0njfeMAakuQMgJAtztyUxEoc8bHSDrxTnCbfC2Xktz2+ZC5Wlwxxwsi2fFASyC
Vh0yruQsqs0XTXh/KIu4sGdoeGbMPwvfADmNgUWIFFjQNG+Kz0fy5oa1DEyFMAWu
e64Q4Z8n3ci13Y9n6yHATCIDGYxaJJK1z183xItaGxmI/1U3mYbmNWJqnWFJstDw
4ibBG+8R4kfwdIXvGboXMNYYAHhBh7v27jhF5dPZie8ob/ED6Y1j0vI8utdNZ4FB
iruMAtEWmXZGB03O3C74vkfacG8mVZpDx4t8fY1v96b/gXsvD43x3U92n5WTWzWX
7FQGd4iIbW39Pjq65jfJScr+TkywlnmZ4c9u/hf2WoGcpmnmFkkCCzAbbV7n2ru4
JC4v0NakKr0bXHKubGFqKXaVfdkej57+WBgbMyFDXK55eYXtkGi2U33SxA4E8qja
fMH/DDD1dYjjWWtW2stv2NSGEzkMWLSgR44IURGuxvzoQsKBx1liTL2O80/pd7Ty
y/+J0Ztme5nXgixbk55ZNmPj5HCkp+k+57I/8zTCcuot5lR83G2sO8b75HSiG4lb
4C3rjY8oP7JQizW5TfhdDZBlJYLutlYMJvDmd7MitRJ5eAoCSiQbmBFIfgJ29Dan
+IZpQBDgZJdkkD4Mdx12MAsGiEH1mUFv6Kby5bWSCBJkyhK4C+OLjZZxx0hocY6S
ISXo6yfiLSM/hoy916CkjEr1XAGfp9StAtTCkSy/pA0AEqy6HIxnxjKsU692Ay3U
fGR+VfD5VrJTpp1Eu6hZcD6QT2bgALFCBrpaCstLIOjqKFUffg/ayQ6Ql8lmtdgt
eGAGr6ZM/PLXS838TAlDpYhjQe2+C8ZvQNsChRF6+1PyCEC7l7fED68RU5wo8YjK
fnDoXEkDGyxsc+Joy7Q7LCQRJHB22q0py9bPG+NDXwFWpZH04WRro3WpYAgnra3P
PglThQse3yn87FVVp7efEIi02jX66PlatgCgBJlXXdNrD2prGh2OodNUHo3xax6z
pIZwjAeoY/ZWCJw0LjxEcGJ6URBgjVDIaFxMxr4evEvwJNfzuT/MFyfQU1TY66A/
XWRwBbBtErgUfpUdgRGApDHERIBiKAT9vx3xVdgYm1FGAYR+kh2ojb6Leqk76QZO
7OzpBmz7Uxi0e8Y/zv2NjjXzoJROYk/S7ck2AaCSl1/QmWxBRg3aLxDD7ZRmpq6m
BbuJqBqpL7qQ3FQdmUEN1F6D08hZLHXDLgzj8WotNLkknv33hvUlIprm5ushmJBr
d3A7AHdGQqDo29sdQcXRcVBR6zWIktXnBjcUtipSTzp8MOu0UAlI88cdU4bDMZZV
cpDFB7E4omCV3IBjccUvMTFetZGpiNSqqWVzuRF2Gk1HarTDlZc6owJu/B5yENKd
r/uO07z2q0fzsibGvK3NzCkefPZdGIpcMykf7iDmawuuDU5282CayNiphKxcQeJo
3DIvoE321s4mrHaMkEa6buqXbQhTe8nvCZwVbeCa2IKp3u2sMG4sAlCkHNqyBnS+
Z+L972CbDDz/AVI2/5zN2GEr4ZM8kSrig228ocTtORnaLQio00TZU4tGDpZQkvfM
Y3Il79noBRrm9OLLqvClSuBaQeGEv8+74vRbvsKdXHTSeqyA8lpF1Oxd/CwFm9pj
mytflxwCkhil7LE/IbPxwTDf0JwbN9KS6vVXPAjc4/uTGe1Fww8zEge9onUvp/uL
ic34E9EH5O2pqm2T0JDiFpMM0Te9EOPFBqUG7TnYPFNuvLg6MKxcOwviEje1cFd9
ierAF+E2jEDh7AqDDE0KhTWmlMyTGXn/7ciy6U9TSV+S9WizROdkayZK/bGrHS7E
8l9k7/U0SWpcFHA+Pl2NmuzWnK1JzzQq1IeVJYnFQeVyrkmSzd7s32cWf4Tic23a
cKtgeRlfab+QBJdxuinIHGxxzvLaTe/u57qB0s9qPXgumN5um3JZ91v7/IQ5FbGa
E18/trrwXy6YA/WThT2z/B7l/acy0bCL6kG4G/dihjznoukppzm94vTWieAaKBbb
NiOq/dTphT0z/RRwVFhEmwHhOaKhPNA7vcV2LLQJPDNbO7LjK7+xNf2xLRY6vAfr
5c4wkwJpqqZtQ6EAGW2NaAw1jbJb1aSYmdevPf83BOV4XcEyWYqJhmYgRT+S1uXe
5chJ5hG5CmcC07MRORMWEqvWt3LILDP2kgGG6vvdHe2Zh1KffG/gqt3ykPde1x5M
GYQp7weWlJDQ1LX/UPAhF2x48whMfoOwt7RBhBQDr6i9bLD9VAYBZ1cKPzil2K/m
IWAyodoqHtk0K2PGWMKZ2R2BsAsc28iltY6nqYa6xI+fRsDsoGCHp2ao6paHrf/B
9ywmognVLvcY0+/5wtCkbRn7WvRS5hK8h46OjHHy6jPPGFo2uheEwkugMb9nQ1eF
07NVJHviUoVrCtZtP5LNQRlmPsjtZ2mWDVQ3wWlSbE0iAGFuGfpMr17/VLJKWign
ZbbVaAOn+goaepUIGBCOia+EZf0nWAwZ7BH/pYYLJraqPEZVEJgNoF0S0msjefwB
bmdRcdcfoLeD0CNG0w9sV2Sf5/twx2YfZOTwubE5EVALTKhDlZ/tFU3YPwP4uBmK
VjmGzcf0b+UyOZz1rzEuKex+Op9SSETwoChAla80P4zw1zskwC1CKReuSZDrTaNA
qh6dZ534izPh4GrHp4KgOU7w0969a7xUoeg0EKgqb+l5lZ6vO69Fq9tbw4PAOjH8
lP1G6kdyfBGCwQxSufKrHdCtdvdvtQJ/9k6Mmd7yCxtXr6ztULBOFVYAa6XbVGWc
eQ9tbj+q6evW5zKkHTcFLgLGxzcJPH046CyGs5EMTCDMl+GZIxfAKBQX7tZ343Ou
F87OO3WHLsTLlq5IBfp9Ta/A7lKsT/P0UyoH329+hV6P+isiN+LgID2TgWHwaFwP
oI7asBsrxxECRpiS3aT5cEqwMYa/aDRXo1btBn+uhrHqMPbAd+k3G8cs3iOGpURB
sUo4+438yg08XIMFD3jmiU4sW0Cvf2EsIPrtvQLdEfY8aLmLjD98m9FT6+macT41
VH2Tyy7sQDHHQVVnVPCsOLNtbzuMD927BIfeNxgjdL622OQQfV7XMjHPinuIS5Uv
aexIfMXvPaGEnxjFuLZ5ec6kHDM0aZfZQBZwTxfGswIVQD9XsK1FRuUZjD1A7BQs
dSRjpebwaZ1JecDPBRHZbzoD3aQlGeuqPaFkj78ioFFNTD3cCoQW0bYomdGYunbS
nTGMarR3vgQQhFuLWtQJdhpACz5Uz5do1u2H1Ut1WQX7hoAz3Jp6RornorZSvoU3
mPles10xpoM7U2kjVn1m9XZAirNaLcheUqlpAfynTqijaPan1k9gMlR9navWonw7
Ann4fRwnoU1u2JQMCq4yRJ2ajydT3350G6qDoFJcRtKdUngXMXVlaaM6PPYJUlrb
RhtcxAl3G/lwKDPLB4dkdI9KKd1fwzyxl7tRwE23VYrQfvmnbgjjLTs7zo9LVojo
i0WEgu6EF9fGdz7232pbHb2AOYxM9a+13ImwNS++oKiaLVIdm9xSrqYGiK27gFU8
jd5PmPB8SIbxtNSrhryYYe4EAkHg3Wl7tci5tvfLZG6uMEU0kvAOsqA4XRdVj+jD
8i37NgIhWcABPXK61np8/int0wOOiECIGgTB2p0F4DIALMuRZew0YMaw1kvP3K/p
v+I/2aqbJtArDeo5sX67DYGrW5e2y3d2hihYFJNUi8ctj645Lb7y7g0ECqCE9BIK
vcVsV7Y0bG1PyH93POUodga2mIqGf5EfWVhb6ITeerie1JXqemPyf+uvSe02j7uZ
jPOiSo1ENS2wNvu5tuDJNq+SKXoCzIzyH76QFsP6DaaSHVt9+ch8XExFBfN78zrT
AjeOD4MqY86w0bk3xMY5a43srNv2l/JNHLWHsEJC5yEkSB4tts5LaeiHHKj4bQVU
N5WAodnyn9x/alhRaWOqep7DuS0AyX/ChlIOAt9o5s16cuieJZqEm0onqJmhPRUy
ebXJHtsHp2MTPLS+pTW8K0Zqw2GpOa6lbjlCemSnPLfBbNaF1EmnJTTafBBI1zFx
KmqOfRQmR8ujXmzSZtm4P0VjeKzqrTLkfkfrc/wvdIo6g1rnF0D/r0VEE8qG1TfB
7i6pCiw/uBklSAIfQcVtxoWOLJ54mTiLI061+icBrwmxokAYuER49WTx/pia82mJ
ppUaT567ND1n6XdHYuRCugNNthRWdLyK57OTxIg9hnjelTHEmcwttycpP2dLlf6n
AhNuKk0CFyWi7T2xoDtjtmEXYFUSe3/4ZaCq8l7gKW3C5XvknVixjsJBQDx1kDPW
rNmwUWBN6eqfozmG8vpMMjk6x//eQGdB37bPWyxzxwrMeHdPKru6FPgWGJtdiSRT
7Gp1+9saADIkwmbxO0kGdsCgCwhWqoulkJTL3AYSicM5IAj7mckVNBzOa5BaRc14
bqyHWtYuVvhXxxDweqlaKRDS1mPYi/LUYN6kc/j4NunHe8KWvEuHnPDx0hEkOVav
dy29pygs4nrdsh61jbr1oNc9itZVAIQ6dnxKFiG2vt747Zoez8HUd9qOa1UcA4iu
rkFkmpsmx8aLmDgbARDuPLwU1ePsDejJlmrr/9pK15DE6zkbxjHlZY6DKUhwmux1
y5cvyjCcdSHVPtthbw1wkUMAOdrehB0jNrh2vVS+bBBQ5Pxk02JJAR5w7R6z28+P
Up2N33FNloshoA0kwRPT0Q7lc17bCCsR80zEubOt3stIEUjZt2xFVKyEnweYHgWw
RaL0eea2t5Na6ghYSr0U9Y2kOjuSrTqAFeFnnebYHrolBgrF+ErJAjISk3hGYmMl
71E/mR9GSNcT100RJa22zlw0zC4of0zGGdmDEiVSork9IgQutYQcEVrjhrorolK2
O0HtHdfBW2OZ0zxV4HGg92WLWE3sfE87ZpyceDPkjQ//iojd/Nj9K27OoD6MJG6O
ipz3X0PCTfD7/mb3EZViOlmKqq6MMxMBActodvpAuUGwMeuAPudiuX9amC86dRVe
jsJYsQMNjMQR3c2jwWjeidpg6BdLIokqmDY9KcvdDMwIKoTO47rp/goO37oGkfYV
ndm02tTHNIHaqsLFh12KpW4URIPZ0q/kNgHFz4HrnQHDR6DmnIlezYfA88h1lauc
S175JFfODkWt1Bjbwg8GK5wqJOego7PCQHaqDBWLmWiucPD4e5NEWOYFGuMe7NhH
Zom3qxP4/1M5gAdJjVpiWX/wNPIZb3JytRsx031NluqtrrdOVMXUe0xVC1W6uefl
ELlCUI+s8olSZoY3Y9ifpG/WJfINTpU2+RBhf+4SvQlsrx7ZWyEOalp7CJYFQWRd
zioDMXAznN1BYQqqQcbGC/xyHdE3Bjt/QX8WiR5PPvdUhz7VeaPo/UoQC3kda74i
C/GneYX1jGvQPj6Pa60hiCOlK2bs9Oh7WzZhW33suRAAjLFhastNlIuMZGX2vO0V
jnnZVunOHjl0nAgufwbj6lDubdUxoqKr3qXxXyqZxuM7ngHZ2IJoUKeSX+5iv+Vt
5gZBDOhWm3aEVXxTIdhpdSQSUQCv8fBbchFg8MNRdp8mb0ifbhZmq7YaQXuOFsxN
NillFtXoAZXHSRDtQANZoZTzUn/o3y/mLOIqfmitSdomEi85wxYLvSX9wnF84p50
czILPw5JBfzubrfL5RxMuH42z2VkU5Y3P2DZHfAKKVnIsEROC3sKWqLqEE79cr6k
I7kgK6sfeRIDm3BQ8kSFDErgaCo9LSxM0q5ayoMtPTOL3gznh+QbGwawUXYcbvab
Eos1K3NKJSiM4NPBdMRm8cfMd0IDEMQg9gKYHwKFI26E30NeqofmPqNJyhV1tUOX
uoMKR12FvQQjppk3ZmfmxFfAO/8rJO/RV8ngUKF7lAJa3cYd6ZrzsB8D5GMgQeHy
T36agO6KwBYfyN9BmE1HFUZRBcKYStvE96dPIpPKLV5gWNbc8lirv3ihkYU2EfMY
14FOfM12iO7UbxkTrwb+umhwReyG1BhbHQgiyeQKGspvkhGCfcALP2lAkJt1Xy4g
mN0nMNl58xMne7bz5ykc0AKtiR3ao+0gC1fqmZZembMf3Z8kD7tunwSeUU589a6/
CQ8aUVdD4TL/sKrWaUCxWTjsP+VgiHG2wFgKTzyUR1G2KTaoX6P6tO729BfonBNE
KSXpBfX/2sNgnwRgOCF8AcwfRndxUCA6kBToXvRKYPsGrkLC1c6Eo0XmkXXJp3hT
B5UBYgCvgM6yWIAkMLuw9wgLFRhRYSi9Xjt1Rie4b15gVMJSxHXYHPPWQy7eA+tF
MM0snN5rfNeI9nmd9PllEEQbFETmZl7YO86LvOWn9iz8y9Q6ceTG4hdjC8pgbnJY
4F9gRMb1tHm+pKWwNs0tAiCCOiEbkfPs/cfR7kXw1SaxloHrxe0A6SfpNLjCIcYC
fK3P0Q5/CUDK/n6L/vnHmrgdgFqC1qyp4d7+/x0MoTCnf4Nqrl0vpRK6Edu49cpO
Q15/GyxRoh02HX7vsM/m8KYcfckg0FgZHCPq3cRl663VogYRsOudIwWyDi449kAd
6wD4cSJxgToEJfzhovZaXe23PYh7aRYqwfNCU/qOg0cX2GBXoHIzBSd11qAucglt
lUYKNpiTcUtAFieNCKW+UqAWs0grtuyyoq/nPKz/IoMbB/PjcrxUeDhilG9j3AiJ
ABCjmn8d3K4jPxmZYRIqse962Z4LWnuYJjNnu5015STwr2IiBffC+1Sa3z2fYbic
pBZi1kJGglHeRn7wMJ/vA+CjVeVL12JpjvWrbMqZI5Gd+upBq/NiSJtgKoEe7OrC
q73b9F4zE5aeGnQO/57C0FSLLdIpsRyULBw3mRcGmhlgR+W7vMC9culoWeYu8Gcv
K3sS65rQ/3vLKZ+hcjeBLj4BPUSyoIyYncu6+TcOIpxTCJ83LeBc5PFPj7QKcqpq
sntqM+zN2AhYdcQUCj/Op7AN9Ei9Tgjgi49yssF62ZJpT+NERluyJ6nBZTYdjBR7
XK1svnoCsQLL7dXKLA53VoMHsyxv1aUADWCDOVcuXf93qpEfTsJh62sHFRGjQ2eU
6Cik/Qo/ahU71Cz2ZZCA2naEJ92OWNpK6u6/q0pQzxY4SvyZMAe5C6dMjs4aBY4j
K/0I+juaDk/HeIgQNsY9XgmZPq/bPRmqDrDtt6aOrmti1OKEp4Tz1hDbSkOnXW54
I5G/7PLh0fQs/04hLD8STsQEM/NIbz6jDRyCJywFvA30BlZAnJEf1DA88dG4lwzW
eVeoCO9PYv43HpV6IxEedTeVLvO0jzsf+yKEVlFYp9nULJgqS7ggJxwY+jAUVW7A
ll2ATdzzxC5QW8aHexrgC+glluvw+8CKLJNJfxV5RVTTmgc9iu12zSnmrji+jDEi
XuDa/Nbug5yKIXO0/oyjeXXFB1i4CWzRhAYekhV2GGeB8TcPUPnIcuN9u1lXqnRt
VW/V3O2tgE52qR1EOYEifNAKWRi/UH+CY/9aAq/vO2GDNUP8UPxFGNBTTlcBc6Wb
K+cGTuiCca0AR2pFxDs4QydzRhY4WOQDCkQsaaGdeW44+DNyOrezyEMR654Fbqtp
FEF9agpsNZY08rId9VXTXE1aKIeab2URzsmk8jIlF6DCLMpVd5Thk+plnatbybgV
dOX0kFm6dBRoeD/Z8FtWKSEFbZACqBTa/8liWXuO4DLPk3Q0CjUgYeXFxch2rZiW
ddcztJHKDk4f+OSEsZaKZ4YJ4q5Qi1Rxji4bCHop1I/8ZdLji3cRC6GEhwTY8OmE
tDeAk6pc4ugzOKxknRdbdZNe8lOk1PyUYN+whUzyQt6MlvkTleQeXPWbTAwiPoUK
a1S2amEeCiGZYoOubzKVV4GjVV6vWBoDRYcCJgMd0JJ+19ERcAPUNN8JO+w3b4I9
tzBqbOuN87mwr5Tb7IHoXBXVfEEGLc54gwbuo680yeN9GZYToRxdm2c02wMHRrct
+2YH7p2yUQii+ute15D8ERp1c2CG7ULLaEgB8OqiXcmWzydo9hNkg/IWbeaPPUI+
gsd6KqelQUiVOOTBdLcKLW8JVN8qMyoD85esXy5e+4BW+4MojWus9d4Z3UNTplcU
90cIbQhVBnAyMEeYd/nf1zR9te0l4ta8Nj1k50hYOD0qqiIy0QC4R9ZbqlA905/A
oskvXXd222CrBPszxD70QfXTEAyuE62XLWemq6tGBNhZXC3GL8G+PsuN3IvxrGcW
L72w1QXs/Ceqja8fk6InkIjMgFu4wDLw3wGjySArEkwK+PSRtfP2MU8R6754anbE
yGutF34a/TuHRpCpBIPkRnpO2FKdk+MP7hea50bp4pGmW5+V+8ueI50vo7gZynpM
pFFlQMgTdnJfTCzrxHLLsZjD1WbBNsyspjS1X85au6St2hTLyP9xjgiYZFuHpv2F
p1K5aNduxiqYR55MGV5NeUQZZoBTT6Mgbx2UJs6mta/WZQXTQMHCn5xkFv5An3KD
SS63AX4n9kiZmdPH31qTLp+OLrZcCASlRgxRGeSCFbHhJMtfb1mb2HO/WZ1m2T1X
WMM5CyhUXzv4JVm7BVnxCmQ01RyMZCW/AT5cTCMeXzTNTSU9Xy5BijKqLKhyauDE
8WRPR1ojUnmqNqXV1Xer/Bv2JF9AtfMbxXcTLVf27iYeY/1avQGNh/a9MQMifl0A
6M+faJVl5LGHHwoje9QoJxWTEBhoo+K5jlK2KjIMaxbhDlF9SB+7w6aAyJuQxJmV
5hIRKXeD81ZNFg9syho4hTlVKacqCsMAJvPzyuRjNpCoaA0iuwiZHqDh6ff+0Yv2
tL1lI1OFtYMbcML7mTzl9SHyD7b/nOtYWtqONqJaJdPfLU2o1tJaoiy45SS2FlnR
AeYpxVKhqlaEbaHzGXyeShL5onX7oL/o/ORbEYEVIOXowB4AMCHObIMZAFQ77Lv2
XY/QQECmYQGde0DsiU4NB390UIVpZgVlWnp+f7MojoRkp3s/j8i+jLxSQbyKUVWp
LD8g8wA7kaQcx1BEnHpECqVPoKfAHEXpG4iwV3WNtMG+qTC8ogxNOrS27uTp9Yip
nC+dp3ejhK786GDOuzFNNh6l1nQCT5J7ZuqtbaMIB5daShfH3+YlilQ4wOY56WgZ
oowe/W0cvchft7dtejv/jR6cH5BCrX8TAjJLryrs+6g+90hcwJtjl0BPewT+QKU6
e8Yu2y2AaNNv/2x8flQ/4UvNC4vE5/Oq90ETkfkX9dxEcyG8DESmW0F8Qqf+O7Oz
xLqSqWY6hZPi071I9EwZpua2V4OaSuf36Fl4KenyeTDBt93mS4GrFH9VOpmZscSF
RQU0+zQxe52vPVFg+ddgU5n/zcO2giyWlizKTo61c0LPzxHhRYu56aLhBn7d9EQY
tA5i29K1rnPnytz0Ap3z+gpoNFBefrOtAwl0c0xy6zclmwJBFFEk8EXaVZSvl02x
Eq22b7QsgzcP+XsixEzwf1TPNWNEZmwMMsdg7F+yKWL0QV7ZucgkUNGqlu4FEzst
3WN9+jKUFd5QS8GYfFbY3vbtf8oqvuj+GBCl2Q1gtdiCTIXJ7PEDZDMbbVbeO7ws
LBw6OTI9DQ4tqfRk57291Z/RapzAq6aGtMwBwtnMbTpBACjOvFsR12EUtgD9R7bP
1m3J6gJ4/8TI5uJtOo7TSPJjXzz3AmN5M3rNm47ESRJsU92ss1EhpiZjHN3wci+g
reZrlcz3TTvrjvnNp6I+GUuBeF3E8j6FBzI47wuFYD1YzmbumyqZ59DBvUaASlKJ
gVOwIzv2KA0LghSOAHdJSFHof8RrS9BfXEB24vsN7pnZMDGY0TqBgkCHLHdtzcz6
1eRnWwhTC/gXWf6Yb55DJdP38goT4RveQNeLSSNHJVIUiVw93i7Fnf5uyYRBCSV6
/QVaetY8SbWsvC54QXkhP5yOrGK6EIwdAv6UdLyZQyLwsfxlNSQkrIbAcAjoXIqE
Q6XaZbRdwBwUnDPWkAKzilPL3rTXLld2nOAlaMzIFFu4b26LxgM24lLyMJY2GZ0b
rGYfXIAIsnlf+RXN+ljO406asS6L3QTAxvX5uIKLUYnkhvWMi1HMfk+6SWtnvEzJ
B3YF+I+ODMT3Y2EE9iYGiTj7Mq+7VY/f90YUWdkp4IVzhRaLwGMhEXKf6k9ljFxr
sd8w1BLjFKivE9wJYvi/VE5OMk4WHtYOfvF1l8a0oDYIzahBcvmAhhpwhmBuXkJ8
2h+nWHautzjEGzL4qpgOTyrESJptzYufGdwgsQnDm4f2ahMrRHhbDOArwcQQg1Hy
lJCk721pp2E0CEkPLlDbSDD3ZqDVmf9bUrNnc7q0sAVL7PrZ5VLTbixm/mjSMaiy
+ntQg5mW+xvmAFJfY0WqjUwlK7H/btN38aJn1/M2x8IkgGNBV5SO0l1wI50uNFqk
qtCzPsqeI/oVHeOWGAMPydlDNrV4gFrIUXogY0o7Kv/e8VMo33s4UqpT8fcnyqOs
F33P+HsEmmdJJgFQHi53gxTc5Aaolo8TvpmQ0msNwpybyMDJrKVOME/Zfg4IxZVe
S1Y/6Q2J7/8jkovAUA938Qgyrrtx5MZvVnkDAcxfu/bDPMvZTAqlhSS+pW25YfqH
CXZB7kHGo5fvR8yJ+tWuHTBBg6xK8sdxcqRr+A/M/I8TZwC8100Qj+8/EtZhLXRp
OURhfTToah+o69VKfxL6r2UPZWnmu/mLiG62gMytkOdJ+aa38KjUJSDGSTkaZeQa
GYjmzlKr05FsjYeIB1y6BI1hrpe7zQDN3f67rTLja+G/sRnv8DlPzeiYbwnPyNrZ
d/fBMPxkd/bU+Kdu0onYqeUhVMzAqHPSrra1arqcQ7c2+ApSmdoWy9fmnzDXf719
pLiXmqVuJlaTd3eerku6NYMfRVHj6wQU4iNF5ki0uy3FYO7v8Q8qAvJz0RRJXloV
7TO2ejxo9gF8vexc2+D7o0E0oW6+CsNQEXRtJIOxPT3cBJrOjCt8i2YwjmjLug8B
5Pquk9reAkCM/Yz5QuWEOj9JyARpaEXyoRyA7rdIpmnpjmJ0hguNvplJvfAkzAmy
U366vOABDMUM+c3HGUL47FfZUjP0EZn4pa28UGy5S4b0tvGZN1MHm5qMG7D6XGEP
qRWSKb/JREknETjKo+efJV0glSDk3kyu9L2XlEttEbgj+3QTaM7XZpoIkVHOiP5y
b57bilwleyoj0vVj/hB7xizaQ+N7MIjjUgyX69gPhvVtoJfNTUfxmG+xFh7zYFyQ
x1FEzvvMS+He4Mde5Bn76G8wYSD0AOZvnVZRkMGwAnQmwvlZLdoYslO0BRZAj/Wn
f5kq/fKOV75pdpbWlVapIOFeAlYGbedkFiSi2QH/e4q/LAXMAjBx316IgkC0PkZ2
f8/Cd0LrsDzDI4K/ZosZuNTXCJlI9vxJSPXJ/JBsxG4QrclhX0QaiwmdRyBG/vTC
H9gS0VKnCa5g16duiVJbN2FlqPV35K++XrrWlUfglF+TvF/wCo8GCYlHUK8MWfO6
wJEjhuTnZM7X/IYVv0ktoGFEPj9WYOEL5A7NZof7NgZIwjPkXdHkLnMMRyS1N1lk
sbKZx5DCTllCW70UMKeLz3OXBMOJthLxkSZIK5tlbfmoR1pfmGd31wa4jUridLIT
q/wDOGUu+tqCRu0rg43fM0JaYlYJumOJgO7vVb1VdSvE2Es9TjX7LVZ/EMu6v3sf
8jKUsuRqfSi+QpL8DUtJ6LLTgzSW9SVxEU09ewyTC6LWfA6czfWk2z4mm4RS5Wov
puGZXQVBfpjN6Y0l/IJHzmF13lclQTwKXSy69JGbNBToeRRuUKfRzqcGEo7gKXnZ
mjOqZofZ0MbCsbSUQiXp7xrH0Wqyk5yAr3Dy+VJtIzDOSfU6vru/65OGXmBcmeoW
EJcgs7CawpxSQ5QW2xLYOwq3zOvVllGS371jZy6y/3Y=
`protect END_PROTECTED
