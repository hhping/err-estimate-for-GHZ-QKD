`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FkJSENtPXI2xJ05eOdXFp3ig7uMuQoU25nBicoAPuQZP8bW97sJkh3dzQik/jJxt
FSBANAikb13jsRDRS+8G/BageVlIB7Er1LKScpWzvRYSReiZ2qswv22AgB+pLOJU
4RyyQE+Nmyad5NB/IHZT5ceevNzDII4QakIrwEXW3UVK3MtSy2IDhaxiYocgMe8c
GJLEZ6PMiUMnm707A3+eMex6a/MUw8uPIiaGLyk9ZLhQ0UvUh19I1cMGB5aaqZDI
vpii/lDHwrVsT5vfmQH2qzkgjweEOinYROvMQdmhBDLdrIfYobjRsrNY6Amsxax9
mEqvciUjwNgGbHzt8M7SFOxwUtb6oMemWkfqXtB2OejI/ZYTui9cDMerMIg15O1l
rHOuH4bIzGe6/SiKGOs+/xxvXwQu+w9P0F+LChXlLlTJD5i1mgNLUokObH6hOSHw
pmu6cFcgM1wZYvAyCWpC2W9zq/t0vp2GXE5ZhYgaE01UCU/816z+m/b2XeRQ9HeP
sIwx+OPyWhGeP8IFGoWIzjetn8ZTcHeErEd68dGR6g/IUzWO5cd8uFGQTpdTEroK
ts99ATq+jhWXQ7W5FQkkOKgIWoA7pKlleJe2wsZAZjFLbphxJGOU31V55/QiFVEV
LJTye3Mq/5zVtD0M/qS63zdRlC6CQnU0UZhFRu0eZBj9igMpHnH/stdHA1g9w8cP
pO9nnz0SB1g803EfYt0gqyYK1y/To69d8hFcIqLbMy7zWLM+lBy/fbHymKlYbpbH
J4To0D4DrHr3F5g28P6UbD70wJ0NUyKkS6yNU3CqrBqrDCWOlEJiSD3f3scAIa5i
kLCllAHe6dtIbkMeSp2/L0iiegFApEcHVFP8+gwzgb2fvXZlm1razNx9Ea1aGes2
1+N3X2vvm/21Kiryx9FmRyQS4yU57qv3VpZaWT99bfeh/tAJdw1W1j8XXjbrUbYV
dTs/1cGih8XmrDkmDGjmCv/WR6SHQ9f/PuE9Rv5N17ENn0Y82pM7dT7hAV1K5i4H
REieGY1/qPCIbEs6V3APGyTMwfH1Oh7jhq1aaPXk4CdW0h9i0kWmgo5DzGft80nM
8zJ2y7APkEA0biJ/cq7nQsCzagYkrhAJ+Z3GxKNA14Q1jwLiVYlWCV2OVhUwZc4w
NXKudIEnonCp6m4cd759s2suXF+NaRZDgtWKmP8j49rQeLGR5QTHA0ri4qiYomVQ
pqw3vBL/5+F5qEapfopMwyVjrP719swhRgdv5TpaSNK3Q0E3Oj0PM0VqGvx/hlLd
pTendatYNt2S2N+Epmqhl7fsKowi1BA5CrLdQUxSA5in+CX1T2seSXU2DXHmK0pO
iB0DnFtd44XO0XpsQd7aHLaXDFVTRvK2XhDc5aAPfNE3ivb8AMSDPQE8nUImb6rU
rB8wTlVJnp28ivDOo8dpTRUt0vB4kHaxwzn4pEj+I0wTjuTFJrj8lsjX5n2lK5al
6NDrbJBODBalYcBoC6ae2AH4bSApedfH9p1RrC9aH2TF5R5nd8RY2QftkGHbpkYH
ReLEFRnEPQuZlQC+cj9i0qEJHqFt0R3DIFQhC6wBw6mplAp63+dul2BDRDobNoeU
3QvuxOZ7d7raXVNXw6CrIXiOpRBHIHopT8fqF2Z7XKU1z9smGmogJbiPesKLZUY9
/9WfZZbde8MWli6iKFVGoADliUb6T4MWeun5vSBi7udGIPqJBrmb92TxLQgfEz2g
KzhhlJg/CNEOPD8zn21XZ45qIj2XCtNpgqUpGaCdSZFpisplbY8HwylnLjvZ0kIo
ILeB60gIeuuqHCvPKwniOyWaGpNG6ybCcIqmmDOmpXKEpd32yjnIKwK/LeelGNLT
ehhfBU41bknA1XitEoJmDG+lggBHrWHEdwWmaCy4+Ukm45AHkFrcfQ/oF+lTZ/kb
wgn3PSeBbd1A4VouNyYiJqEtblIOTjnqbyrcfbx+KI9WUN/hjfo/IcnFxtR4qKd3
peyFo7iYzsxt7wNnCIMHhInHR1zQLYiGI4x1eM4YqNj6dBrLySbzX4+SyNoAo0YV
Q4TaMrRVm8fCU5Fyl/nzdETK4Fg3NmAEuPmXEbYwHo9Z7trtcvmI8hQJLp0c0/Ww
fzUdtzdKzDeeLi8Db3p+xLgrj2DeolyP1/0Aps8NYo9M81rOBrHk1xfwhCepN4ug
W+G0g/cr9zpUSiVLkzunqyFLURg5f8DkgXKd3gqeqRQf2+pXGM7jt8OXzmkYvVOn
yjv0348VvfEY3YUj7boDHBlnD+aLtsYMmaKrXIH0TA7aXm3UMCaHwVupq8gKTUjX
xoP5MHlGVV9jlMbcLpzmenD5qOs4tjYe6npN4NJZur+JVZ0LmrfnHSp8y9bUhCMQ
HipXxgsUvp3dgN4lB/MwjrCvCyKa7jsfzm4FI8ohgIQKm6FzbhdK/cw61RpJGXTU
M6wJ+H5496FHEbEhF8S5dFh+7JurabWo+XPNqhRMAlJNygrUwOaFA0O0WyBKb4cU
0oRMbF9WHEiyXosiL2izh0Kcn5Y1kwUFAcOOk2w/0AzaRKIwaWpg+JffBOrOmKJo
1Pb5mjeK3o0n7RIsQYcixDThHHiOl5CabyOsjxJiTwN7wLAxS0roa8G6l2TwZMps
wnsR8E1QVHAfuZEIfWURAWX5fpxnHllN9T59nmCqlySy2KMjzOtyC7FcrW8x+nNt
0aVTBJpRLyQJeFiNRjwHX31d4ZX7QhfaKzuZoc2rWjfGyHgigXj3+DVJbVsYVBfw
3pvfJ6nSVOc043cbNTH3rxMe128l9GUQ3l3jNdQEiRz974nhVhFST7KLL24GajYl
aIXjonR7TtjV1nrPW2hyQUhGXLmejM/owcWvRE9nSoez2R8OCMYe4s2vwdZMv6Ki
LX8OXJs/zsROl/3/z6433KWB0g3PQkWWrf6AFAwSV64ZvQTzXfGHOm+IZKjtfS1H
nCpTCCYmzUn8opxggLr11Wkm56NOHlsAt0RQptLyLASFcMoEcPzDXYsI51F9CDNq
nLENI3WMnVYEODZYgsI8nJQAOzZd+upL9FfrjbjX72fgO52mntWg1N6oMi00warj
+vbIgyLqV5AZSdCWEZpbOXTj3D6rooDpHhyjUbieAuWtv9RR3Mg1bqJsfdcFjGKb
2RCcfUvRlcbMHuU2YNNsLN0rMGuCVm3s7bO8OLc/C6M=
`protect END_PROTECTED
