`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZYZEMRF7lNwFWrxX+sDVpg3183SQFoV4rOi9eV+KXkvXVZgSUKFCCAJRaHsvA7r
NoQA7NcpKVSE9/SpxZi99X9v/vkLQV4+Z+bsXJ4VGEIbNCAVbj3Ju5+7cc3iwZU2
Whr1NR5jvTSQyMW1t99g+hgEQCf8tCnpFXqu1R+uP8sViGBW0be/KMxwfuLnC0Qg
LBlg6GG+ycoolcT6643FXgbQzbAvgcmYQQNrXsVA8ROBkkp4/lXn0+tG+eje/Jpv
cbkVc/9kMd80H9hT49fr+yeRNA7HqPIa9Km0WHAEc9M8f3O1YOUJht6pvs+GYSTk
dKu8h5bj9cVnQQtm/DdXEFWe+9ffm+GD7Sz58r1IPIPrbsuX7OmyJP2q0lU9slit
Hea6e7HRpBZczxm64myfQxtYbIW+pVUBehi8nD5e/FPeNGhj+8nYmdtW6K45VzIg
sAMs3mgrxq0I0oDs/E4MS5MAUjQW+89pLh12Igx3FlAXrjPhON74cNWX2PdSqR7f
2WPFRvXmFO7+Vs5ZJNLHVhugLU3NMEnplzI/0ejaAOs7WkmaHUn2OVA7YcuuTnd8
Fp5bZrZCo/Lg+zuKKzXhNRioMJR3ANkg2BVoijnftKFVRbTietyOJcF0vlHdn4un
s29iz3bG+xrQbqn2tCXm4GMlx4cz1iz3gqhsLUJ+ra7FFnsliWWuxMgQqs6+rRMV
s+1rtmo+YPw8H3g/IGGkH48/xKxiWY61xbaDk1bMKycxJ2JgxUYfRQjhU1umnXzV
rZx2Ln5WPu/IjvocJ96NsR1BoSTsxMwvA4636KDAJUjdcAti5Bra2mZGi7HChVS2
Ebx7+PK2f928EuiKvT5bsShKBtcn9puk8t9+HxSkxFkjnqvh0BJq5O2I3aqKny+K
o6zUye+FVyEnc1RE79TClxqn+p1nJMLa9UNSrl4CBb3ZpYY/4xKdPgYYUgUJ17uC
QwcvbMeZR/jcj5qQmr2SQP0jgBuIdkxhyZjCDq7A2PxSFYlWDDRidfpw9UxjpUsO
GUr53wn04SrVSPOD6FhtnGwbSJ6X64MxOdshvvQ/1gOGH/9zmQW3pgoJvMqDYVLZ
p3MBdmAc2khLtXjwUYEbYJjwjcwBteBZqvMdjsZ3uJgb/ZIBt45uJOqfG9MXV2gU
Jwd1IXdIPZMztMlvr/PwP3dAcSgOVBGZvU6rlHMsw8a/FoU6CyaU04UCxV84EzPI
v3aLF6zvCvV26r3sv1dT0IIQC1URAyNrxm8cpTRfnR1M2C2XV5hfJYPAtW88XrSw
S8LgMXwd4vLiPkfYuR0Ojg==
`protect END_PROTECTED
