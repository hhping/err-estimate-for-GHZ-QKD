`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M43o1xs+D8mbwQzBHIB8viPaTK7JGGYGqq3TVNuRuX7McMnVxKDGWkgoBpZVo15e
oVu5xWP/sSe1Hi+wTVmip0acGW4gp875ZKbHf9pAh6WhapNzRA1h8jo7vc0jQhHZ
ZIu6vrQ2XE7vJp+LtcW3YDki6tRX0enloYJSBr9hSYBcdYwvOLVub/MXJOXY1+6n
kU/PGX/sHN0RfI0oiS5HjHWZA5H3Q3vphFNIEKrCBfZ5h1bamrB+6wMqhfOUO/n1
X64Vc+f9S8zHwuKcTJTiU2iuZN2Df/0ra4MJwpn0ZAsH0t3MApfwPwM7TwIj2Rsb
tLRgTXt6ffauoeNNDboLb4E+241W9UbAr9gUJznCwggXYKjrLdOkXwUnml69jL1/
g+Wl/5r37rV4pGnk7VhLpjvcRBLCqxJ63QlhmqoN1fp6jA7jrZm32at4a0LZ8s7p
RIOGPyRFB++fmh+4fzEzwyvEzN5tIrbgGoKYesikxJKTstYXXqwwSPE6o4Rta8Vf
5nDMCqiramIZQqk1fXHngjekhzUYuKYHOmSBmIgzS3bFKrpp4+g3ptgB8jrBYCxl
2u8jf1LiwpLwqgIJ8fIh1lZRZnwVt+FgQ3F3N0EFxfgMVCph9qJm7S2afT+P21K3
a3xe1lnlZxbjuv9AsOSo+MgYtU6PdxbrNCQ9OjZc2pRnn5jpaIXvQPnB4yQ0vXRF
qzo0Ccv6u3KYnhN3N6njKu2aTw2lyr/6lGSeYbqQ+ra5fWr18GROfKEAkVs5uI8m
/TFdrzrqcokIULdRKvBfpNytapPokoDXRo7csqbuSDdCqPxeGydd9VlqJTeZuTAk
Sn4L3nnXf9tlK9fs6by9yF+E4u/vwTkzl95lG4+rnGMxm7knT2OCDFavjc6VwbQ6
l/aQxSOE218qwUIgC4Sng+tuhVSZvfhcXYQ3LpxyodDXnHIdyh6dDJC3ml829kX2
vSzDQkedoU6nAHnkanWaRBcSQvpSoy/dSQmjBnknTP+GoYicXyVK1mTGn/45RFXJ
S5AVGYZdeC/ZXVsd9kB3GxyE+zkZLSzdAFLW6z7Un71+tjWRgJGvcZqjVSrteoTa
IZVakG8aceBjPG9o+EbmS1SKuCzS6UVfqph5b6g0C4SEQB/YE70GW0eJAJhT2Jdh
7jeMGkTITVIlAJDvHVZ89k7hcA7UMvHlbtIgoJAw6+rXg/pmfJSO7KT5zhz/ezmy
pyreaJ1P2bDXZIAGEV+TaIPKqGf2jNp3s2WVvNf3MLYAy10iPdXMcmAI7XQYs2U/
vswvU7hC+ORtExl3Jm+tERx7qtCVteVcaikYiTBYWG3zJ0MkUvGUCxIT6T49xwJI
2uQ3SxQa64Br5Bg7XjR8k8FFPxYeLHlCE7nd3sCjkltyWMyBc3GTCLeM6nJt1Y5V
WDuow2vkJa5+I1vE6nKPhLcleknm7auqul6pTd9uAcPhXeAx4YE47Ta1hYgxG1+/
e/nVV0ZX5w2h9DIFkLgx19w+IKGa68m1kV4KKGWQDX2TUj7ColY4CEL/eDQOxFfZ
KM0GaHfj8Lt3uK6Ezp6FvMYS0SAjZ1i7IrW68/VbIjTpQHusnyOiorJM4evGlKHS
HMTKEudsmuxp1ZSCFegk2wMhPRAHY3Dc6uQL3gg2gsIbvzMrACJ4BSKMu1QlFYRa
NW38NGkPPdyTIXmSNzZjmqWfgB/V0pwnU8aFOAJtonCnHCm1Fw5F5nGFAlYh/N9d
9iPFB3RsKvEwaUBVko5dgH6EIWP96R3ApNwNeWldw5j3M3JUj/TDm9kp1ktCsJ7Y
K7PrCmM0hFrFxON8elM0yJ1gBfi3SMWck3UEjMlydO3t3wJ3abVV1JzPBhETkUnD
STpPVKeklEGuBuc8cYT+umXHuRUOkGSteHfcnAiQDbZc4OE0NgWMudKvVuhvrIxP
I4ubGok0NJy6+7rh0x+Yzwgxx0Ru7KJgAN7kKgGnirb6PZvaw8ZPWOj/IMAnqHJ5
dcb8kZMWefr16oqptS4kkEzDik0lcANVeopa4VM1El/Qa9HWnkIFWYQhhsS9amxc
E1O1iznFMwOEvu8IrDjPaMAki+PieRQy60H1itGs6qO14jKikEkKFPF5tohMz6Z4
5T4Xi50EP2yY/wRaxDtFH6LWzcMzN5X7aL2eZm6ZY8WQeZBVCAi6WxDUFKA9jcMT
eRvWQcNK3PMuBiWidpNr21hs9aaPuS67Kb3fs4aK5A7j7zkjz0oi/75JqrGaiuGb
5z4FXkE9KG2avCTgOkBSyLwxB4AVrxaKU6HyvInUZgyILmner+RtlH6lq/15whUT
oiT596eZRaBx2d6YU2aV0sL5qtdaRJMSj7jR7ho0AE9ACSB00MMjgC/t+YKlYbbQ
R6PosKjUibUaIGabkQKOMMaaWhPjc/yKACtgfYrX/Xl4KCn1gFkYx40Z/iTAY4ou
D8/jUCr4jvl0cT+ulrpTMaTjJ8JgeaHAInfs+1yKgBfAta2dMoF5Hr0SLUIZLCKC
Uyqkw/NgI35PCyer9SisbzLpXR5/4x2AYNMgQTLT+x60Gf5uIE4Nl24QSwI5YDjo
B0ZgAuhihO0w0yIygSaYqw6Mv0m+qmL6KJr0ihUxvddzZfZiQIPWNw603qOUN6as
beuwQMUVqj+JDchguaS3wM07d/euh+D9PtjLLtpYkAVReeQy0Q1R9Tc8swCMvTSe
8CBs4RUqbVLRGcyaJWjVVEhKSb8UxWl0B+oNOkctRR3k0srg81jgfepXUE04LGtc
FAS27wE73t7y9mqP/sNHdjve2RUc9ITLzOts8FwwuXqwwNn4l/ICxC4qW9wYnEB7
Vie2sh8e/iQPmYdfHLO4NXP5c5XjX06p67rWTJFteYUScmgpL50km1slyYMm0gNh
7f0M0lHNpAjdIPPW+JFtE/iXlroPRpJW6vgH1++a4munfTfOhRYXJ94K9syvh1zH
WPSkxbwV5Xk3Jnl8DCR567cOVgfG+ZbyAxFmqWNDEyrdJbyFvJ/hBwT3DjpqazsB
tpPvPUkaYYlaVdGR4hFn4VrMWI/Iuf96Rvf65R9t64UBmJTWD2s8LoszVjWaCjvG
51nstTWvpPOIc/xHEyTPcoiireHNjIUNgtRqpyLj1LipG3LWuZhl5OkzXoaIlJGZ
JtB5iip1PLrJ5m1H0tI0vnHomN7ZV5mG5JGYxt5Pn7Sya0QjfI44S/wHStYXnNtN
gFCo5TCKKY4JoB7LfkY2hJeWs6zOeeSbUBTrlOtX/7XTFD+5EeP0AvLj7MCouViW
U18Dxz5AgDPxQS4DSNxXsKaaz/dPPmcq8TjcdqFWEGeHO9IW/fSMG1BbDB7QCsQ+
TkFq3yNS0DGMkLNgi7PCf4nqW4vRSeBI2z6x0wZkBJJy3XfKoWzeXjNhF4g38hGU
FTFU//N/GP7s3dlYfzFLOVPyBSl1VU3MXJ/0G/FzzNX9Nm/1hIMnERPnoCxJxgr1
B8lTZBXhwS9EU9gpxlO+SG3n+zl4idYTmMRPPoFM5lNAAk+qw7JNp+tl1mmstzCF
3QrEkrjMRBiLXDZSl1Z+CMWCD0vXbiPwmF0Zdb2WVxTKbi+1V/6/DxyXNZNUjqkt
xSGaBtqQkeiQsMpghkh7rBtvS2YaIfPG+L4gXPylsRsWne38GrdRQSFarUroaM0m
nsKFM36ntNzDlZy2Nb3ZAQkmNO6tmtr6on8gAWmmN5m0tdc96tsJeVtXttYuFU7n
kWuhn/RAqlbeUrCVatnx5C3pVC6NCnNYqWv4a+/p+HDL7Qf9y9i5ghEv2lucjCOz
F8hWqtauy6HX+ZRf/rPurXafrORhs242IvfigkkyfLzG8u6vQgyaqfJEq+wxKkK2
0iYfFaUDxJOz6OeqFjM6zBN7wmSOmXMmcLMrjrZRq7XwbswZq+SHMtKJ6/wVFZd2
ozK7fPccGjKgNX0KvFk/7Q1+rO5uzvFO18AsPF+OYdv07rwXGcykItoHpZ1bLheY
NtaJS96Hln5oBT0Q1wqpT/qMYLcHVxl42y7T5fADCfpuLiyTcQL5FXnyExyC70PQ
NzcslX3gQBPW3IjY2c81D5XnHf6RXDTxsJDTf6GbKCv0Q4RpFtSq6RPL4MIBiLZr
wXkwVYEPL4ZTHG0ZxHSE+tHeoC4h0uwWSTm6F+LJepQuCRkh155HS99fYHXFxrxb
SaNdYCSnm3Z51sCpjCKnZbZ9oCVIsHU+wfTyUMLWQDWrSjN/bFZvauOTyQreeV27
i0OvG5xSLytSJ113buBKj2kfFzEzDHx4EIvSBpIgd3ErUcrGkmUxEOz4hcevi3Op
YCL6NG739r9aOomTTfS6j/AuvcQHIWfFTNp9hJ+bs8f/WGuNnVxRH8cWGXA1c4TJ
KmwmDUZK9LckQQHTX1LTQZBZnJUSLgb2Eb+zXX7vs4CmNy3kSTZS9PHR6YD49cUO
jda8kBKzCxb5s1GsongHRHHDDs+r5P8sdVQP+53rbIl33TIDG2YCx6UWaDY2Sr6q
pysQ4lSvW6uvn9pvd1ognEB2HVNkq/yk0GY7iQUQHZRbSsGqXydr/uiqK4o1XPjd
xlEniTO5lily5Alb/D/JbXHHfMrelO2T8VhfCJP0AvQP7vzX8leBswfNgNtgUcVy
o8iaLWvFv1S1zL2NIRLOwhu1CP2iDGt5jmeooxp57oGnFkvXEhA7BHD3M15Y299A
vZC9oTWH1QBpll87blO0PNOsSKc5b3barig7TF6t5zccF4tE4kDXl0eAUnmHh9JR
HNDZhCZz02MDd8TFWErgOH0czFwbeQzc+gKxrdBVULZQa7MmUmk5jg7FjNZuyRcK
Q794VKqkafcOs+dOBqvRczuwl9xRe4JZiqyHPF9xBH1vIfwxk3xKKVoWaHpljFSp
1zuW1AwuNIUZvfqAPBE1sw5sqk/qXsqq0qD6EqMEmo1uoWVZ85wult7fN5FA5RAw
qnO4378RRKpJnHCV1/LDRAGwPZP0zW5CWSVCw+bdjBvm2lziXN1d3r3hJs9EgHAR
iaegHEMz3e3zkDSUmYD0orofnixzePMoggDoMAioW+hsI9NOK6Ep24vmSn6aIXt6
1jByOGwaVxz4zgdqg34JuCDCPdamBwEnRNG9Ezh9FvfHBLBOj84xoqwwHcmKboz6
2En3vQjNaaIejTyDRIdEakNHCm3p9M6WB3nb6/QPqDP7HMHQCI02H04CP3NGgJ0Q
67xjrYLUtOcMtePA0aj93Y1vlrYYL7usIxBJv92H0znJWU6dgoqRKqLo09mzXrfR
B5LWeaojz5+c2pcMTHCEPQx2EhOy6Q5iPMZZVgkWTZbpCfiS7MiRfsZBr/HNK1S9
ypwA7sR2zkR2cUsLgWB8U6E9sbgVc+lcsSLT+xMzDIiCSNUbFdGYoGlc8/eg1+yy
r5ecJpNvfaXP5pYAAticBOU7zPRgo/jyPO9tnUN8V/9ekpzIXQVkPUc/QkqDYBRm
UxaxnX3yImr1OltKop/GT/XL5zi5PflNKYiJzoK1Zu60n4AqF78TPflChfcfQ0Ko
V5z8fIjC/y15BD29R1gQMuupKOvGBmQcw8t56gD6Mrd3WbFgxgC0dtv0eaVIUeeK
EdLdv8j2GuuZwRapbxiaO+T8dykvzLbTDgGjOR2gAoa4hccLuVSa8HSQG2O4xYy9
ZikDLuIrve477CdIIqqItw79416k95x9eHRBauB2FUx7yZMf6zzd965ih9Wyf4Ch
KKIIY+zOT25qLqsGGjRxPHJAg4z9UhjJ428BiCDtBx+hzoew+w4tf1i9e288cYdm
oERibmQ3AW2WyU5mAFz3C+cyJAWykWKTRyzBVNN4k9Mfuph6mxJbBfvV9M163Lf8
oYdBms1PSEpiyXU8YppZGTvW47o8WBUi+hAOKxXMYlnITJWXpgYmqk/fdiAyyhDr
CX/P23ZzRPXr/NCqugM0zQd3A2/LxLMJzKGWNdhT1iU7Fni6rM1o2JMeOzscNceX
APs3yYhkV4EFm7YqJiI3i3e6NaxvkQQiy1yuCpvO6caXnYS+rmz3dfOIg4fUgcVl
M2cv7hO96SfkHw+mLqkAOHtwnD+7HxUOVEOJKPXlzOh3LEkc3CW/kX4G6+QD/16S
clMJd2kMVYjPpe+EXc/SEYRg3XrwiTseZpY5SGJtLoLI6Czjg3nEMhKeoajjay//
dIDurC9mFjVyBP8KJyTebEMVKFGIAFAsfknm6marvny7u5y2tDzHVwuZPTIbs5W7
LMQ9c7CdMpCSfMUz/HmsIpPEQJkYiGJWzPwh6x8LCGWS9/fHCXa/r50XBbyefsLw
KzwThlR+kNt9Ijg+9QcN0VT/ddIXNAGJ6TF94wrZ/kGwbaji550bsYw776WR8M3x
mic4OJigLg3/N67/LHcZNII0990MarrHieRExIO1CBHkQ3S3OvnjfWc/puiGdUKw
47h7DECejFWIQBFfloFtb/B9uYKUHomccruEGPwA9tAK6Y9Mjo24tNhYl2eHx0hF
/tKtPwUNXEynhybp/XAXJ8yYr53wTtkXP0Aw3C3KLTqyjUdEJvdVFBsE5cMWGfYm
cktiu2apISxeSPXgj7fGe3fOg3H1Vy7CviicfebBbXEZuMIEUoY8aLzcMvrCMXvc
KWN2IMRO8+44qprl53nHBeFmCR4VSO9AjSerhxz5Ai92EpwquoI5GphtHiADVcmk
9l076bOVyS5VOszo7u85Pe6DJ3QTJJhjIkvfW390EP3InyifcE70iQA+mFra6YBv
Ibm8xoqwGzyz1VL6GcjGUZHvYoIfxx4H+OFCul1JnkTY5L+OMjll0oVchXjL9+uA
8C3Pk0FzVedPctXYJ0lnc72fW/NEKX5+AO/ioMyetDuNDH1yRQ0qNY76nron8oQK
LjYZmDGqmCPrxzx0jeNQmhEJul/3/KuuiFKZ0zxm8uB6HSksCh2uvv6rv+KI8PNG
yvL7o+Q+2trXb+1sn0p9gtAOo6l3A02FHhvu2sQYTgKQQnDG7oAMtlRobeYSyUbB
EfL0JDvwQESbOhQKDQZvvbEVNGhvNUgn+7fp7Oq0KJNQDlwcNkZcxDv5PLsT3jra
IGoRFLHef7dIYtTNiSeIHpA63Q1YBol0ayDd4Kq6RQ5hGxnHd0D/ao3N/uK6A+RU
gbFgvM293/rLbuTQRe6rAxaoj+NfC7VygWrDeEKFQsXK5JNySgPSnKPpiLA6bhoQ
eonAXIimwSacMkQW4nNxGwznISmcc8bw/dlU8to+0NQ/PkuV0i/EhwnWzL6tyIyC
pTt+svMOTEjSaSDqa6+hJzSilQejRFNpeWrPg1jLFtEDo0tQ/te3U59oPxa7udvW
On4DiVuxSswoWi+lkiPW190HYK/SNWNT4R9CMvU6y9r6TnDgJGKHZEgeLMjYK4uh
AJVQixSC8z2D66oOH+CZ/hW33/3cxuL6VKlNE9s2P18AIqffaCk+bBuu6BRvMjOV
cd7suenzvkWP3+R1KLE1nOh4k9DV4iCR5xTF2533GzgOSKTdB/W7ga8iQIeahgbc
JXmMyz3kjEwYrRChFNHRruqI7ZKS2AhQp1bKDSKBxHWRvysu8nZ4nHwnF/HGRccK
bHTo68lPlf/Dvfkl1fsJSCjen+fiFvvGAlTq1Qpm/kVgGV8TeYYaPMeyi08rkxAA
A6F1/nBvA2f8I2YAVbVdfLOz7cWv3MWALzsxqxc09vTIDs5PBzCTmgjb+4V12u6+
arR7ZM1mgyqrjsxvgPztzB9io5e7bpak7b54QTUPjLhdz5YqhuAReuj113AA3IeJ
Qq/SNaw0lFMcO+ndRpvAaVuIvNLHsiudLAqQF0p5uajniUTwAFWqXVs9FAck3ybE
pzsOzJxxcyHLEweutUV6IZiwNzcTN1qixL2YSttaN/nO+YYw3NkD5pPy+SceN7uE
g1ZXauiCGZC/Q4soNifKxI+GAK48OeOwbfigpHODnExwssLj/Fn+avjejWJnuGmc
T5tvqXMhcd2e5SF32GFXPlyzUIOhFZqBlWMIpw6C+1Vm+0686ed3z+MSiO2qfAKz
uivdl668r6NnCVF4svSPpUvUVUXKocDK4UChw+PgJgcNjnBEPDMx3nIv03UGMXMk
U57jhj1NyNp5WD3uUipytvbP7BmVxvcPG1hdIpQDdapDPJV+P1LqU+8TSnlYwr0I
7c+HexHXWKXRO1pyydPMCgF6FWyOW/4BKSUw5J4xS48OFi6c/Vak4ZRtAVeMmnCT
M1AL+06whsVUhS5OmUWib97aI0HnUy0QjTHvVFF1WhtO2dvsAE1mJkd20ZKZPilF
hgPwXuLCgeVKAfHPFPEV8WR3E3vcMkAptMoP9EnrT3hw+aMr4/k35hlHhpBEm4LN
sIgnnt/y8jVaMpznd/Lhyr0bWiaXeRbM21CKRwndNr356fcaseQ6534vaw+zidiE
HUtDc/zXCKU0BVO3I9oFN3ckvfBk9kWYQjtcJakWzAVMedJshzjIk6b7bzyBt2JJ
moRaJJ0Kcd51Put0UEmWl5riR92eS4S2NYK0LDGWUo8XixtCgtle+A/6C+2er9zi
XVYfokdu117eVKAOr3APAY9P1M2wgQrqCgCaxZMZXXuOJBdPax9TShUaVad8NZm2
1HBby7254gecz4XQRTCwjPeN+pG1WenxWnsVM+I5fcmItZ0EbcEgJ7llMoVHxPjt
LY0e6W1v5xKE8FgyNF7fJqV0G4cSSk2pl+KPK0/2Y/U=
`protect END_PROTECTED
