`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AmKlVDDQPZ1o/cJh4cwYst4JV0NZf024nGECICp8IbapqgH2ITwfarCBl7ajTvOC
9yxM87Jz77o0BMO+e5t1QhiVBeniz42+wlxf6Oi9VixxRcMaiAf1ns8qbbPTBXc6
3ekwwXR1Ev5dl0aOCDaCgj8ukkJjvUcTOdbPozMnB60fdqVOCky0th9JZ2Sy3Lvy
hxwdiUmmF1ZtlMPDm0Fi2g1iMerf3WR1RdlN7xIyR8W+dKakmFX4zy1FraImGCuG
Z6X/8/V66J9rcnHL+AXODUPrYoVtTlxiITTkIU0QbES3d0BlX3dLBXwxq+URsfbZ
BUR+qmmwcgWdlp7otWUY/tgRszkZlZaoZ4mQbZebWmv3dysvM6xXLVRCJTsqqY2u
XNVsKJwgLnDCyUrIT4CCBkNaNsXMhVp0OTDVzvdq/6ZoLrj44yW4tJ8zkPGnJW0w
e0nn8BsGJUmwMsLFBtUkOvqVxsAImb+bNjRy4icTU8xypQSR4ROJy4RG5vQtBLDd
EfQEJ1IRrcGwHh7SpubsMX0Rsvc+YOM+T1ODdlQZz8ous+MX5hOZ87nKEflHiun1
2A0IX9f5I3tlC/9uP1WnY4OGY0VIgAZv0EnBh+XvLcovLeI8mTZHnWW423r1Bnqb
dv70Mv+oi3hjWMJjFq4hePyrRPvOGcW51YDe42PLP2SJlhehhks8oifQinB6i01B
Og3SLSCErfPOZQPRxBGKosIxHVXNYUt9zMo+mbxVG9o/98kAOGBUvTj/qFcdqAvF
4JhT5ZMLD/3Ak+g1YfMyUp3KBZ3Ipx60V0uVVN122DkRJVKj8mYU5FpFofI3Ksla
cJ+peiZI/RzG681gEiYkPnuPjfQlUsRPNzBkgq6cO1+GgDKGLt+Ww6UleCcokK6X
rlzJ+FJa4CC75w6esZhOrboPAHHAIrvNcYNkRN3UdiPVxqKoE/5kYlvj+1bq394C
QwOjy1Y1v8c5dRslmA5WTxHeXtnYW3Utefa6bBhIb9YsVsQKDvgtuZGWMg4aHGVn
n+uKUYBkEjn03c/61Dp0Ervq66rl8EJknTetj+dbIZDeNSF9pkTeX3IunGaAZjZX
LJZVQZ6XfbZVQVAPJ2nggtrzphv9ZRjDKpo+vVNTP15p3kcvoal+jmctq6ho1lRq
dgJMhJFnWVx5luNYijhq/ukgzJCPDiw8r5p1gv3ZqwWRnJemfbkEnxQ4QAwWAWhB
ihZB+NW0joG4GRdH1KEzcCVPVKmK2jaI1qe4/if81q3WLXskTjFm8zteCWmT4dqN
Z2jKbp4sqNAQ+CndodOVBu2NNp914YBydATvVUz5AnFJuHfresf+bT7lLX/V2Mxq
6KVivnhhUt08YpkPUWWmwtnmdu6mMHztzNlQ1pXEjfPVu2dndXu1Rkv3l34oXY0G
xWV34fBzquWK9xDDYnFRlOacR5CeFewJWTOVTLqRMchPW+2eZvW380AhPjgm4FL6
3+Si8pUcLbT0axNfawVkU/9foRWSWKkbibQNlzmKbzo9GXtyrMhLbYmjqT6re6P6
c2qk6hBbmZpREu/E85gXbIP9xZF1xgAEHTrTnWeQ00ZItm31NGdD+sx1pkG8vcQg
RbB4DAIQUeSddREYYrvkFyjKeg2ZfAlbmR6qSYACCBWwRgQ3wEbjsY6twaFji9lY
bF3baDJT8JcwkvfCA/K1hi1hq416WYbl3PaXdnTsDHS+tAiYPisA8i5LdngFkbTt
Fly0KDO6ahsxp5OQb6atkQ==
`protect END_PROTECTED
