`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSd3yrrecTg7XDq0NImMODm/HcQXuS45qFWoRAACRZEGtsIU2tS//BBw1AOQb6V0
G6dL5PuzRjwnoO40TXX4M6PIeDc1gzleX13vFDo5FYTwF59oPv1OyIR/Bk+l63fu
EuxEdO/Du4RyFpd43/c9Jd8TD+JpTsBqVUdsBXe6YOceW8eVr4L2ZHGwIKa2p6VT
ecVze/tNeBMPZ9RX6EvEX4cK2mczoCkD2M+IHtR75smqbMVLu2LdsnDuI1VPbbNI
NorjJxqo2c+3a4o/aCNrmp4x+D5s4US3YfCFGrMPzPzvL48JrWL8H8d+8/eyyueA
XX1p0VFKc4bxD1iP3A4L3EIvgR8rgIMUspLFevEQRF+n0A6F4GOIKiKoZT3ci19W
PeSUPeiUJsjTdVdQmL59aLchYxCZxRxcPZLbLW0wuiG6d9CFNwOaU2u2qiA9ErO7
Eu0is3GCXDJWiA59oIMKTCsjllYvDs+tWQ4XGYafKYxb/hfsWahGfpWb+JLrYXwQ
enyFOiWAdFJriyALYh8QIw==
`protect END_PROTECTED
