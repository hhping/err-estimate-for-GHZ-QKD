`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhzMCPO4Xd0vhcj1CzgpXAv3jBXIr9W6QtEfPt/z7eq8eUzXDlE3Sgm8p/gzQ50j
ijkN7Vb7nHyYXLoFDSnawB2CG5Dtu7p+CHm8MkBhRK212FRlMXphpCrMwC00D9XH
W07LFbd02MovaXSAYkYX7BCxTJ9oV0NvlP+WNTvWR900VLurSTtOQ5xGjUXGVYug
wggBVHtEwntmyrCcTKQqO4cQeeQlnbYOZVeuxyZAqhIkKDN4a7HjDpfkSSLxl+ex
q8Iwl6jkLuTDwCPU2jBDLZ60yQEDpyWbDkZCJcXKxfSHQZTnm+MaLe/GoiMy9ujO
HMchPLdqD78GY8u+3esUhnH7yUlQgJa20JVwNLlN/QCBcNfZCAH8dA9JJ+x2TKME
awgGH8UwXrFJgNcxI45wSao7Wj97l/FHJfB3zLNZP6FY8wUoyavE0V1kq9v96ATP
yTAbtBeAIeqsrU4HceSw/y1NxBiqe6iVe3boA39p0maTlpddJxPaUSD/XJT3X6hm
m7ROtAkY4QI+r+AdAHGKBs2VeZOVcz+rxnp/hG0jPlflSrsEZLnULAckRVwP0C+C
QXgw052dyJjw39E+BqpXos9tn+kxR8EiRjScq9j1uOw=
`protect END_PROTECTED
