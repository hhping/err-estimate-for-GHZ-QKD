`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBpHlmOeq1Dni+L3jdz9BEjW6rDIYHB+B3OaJXYeLiaT2DPgtsX38u/xLCvDczDF
zWYLlDfjhFpTjZuHLwh7WDsP4jIf+8xRjxjJR5BFZ9tbH4m6qQcHALbR12rPX5Ic
JingF0xCFmEYtWP2Eknd7qL42xlGY1Z4S3qhyDpp1BLHMtOtU5/kGNeFC6DC/7U2
ihGnrVY1+rdYa5RCTZ6khCRr/HHtcKxhN2LhNJZ0RWoBsZCIFn6R3fC0hEEGVVzC
V12Ftbs5b9Q368L53NWqQ76Q8xeYsl1TDhU3YcvSWvowj1hhX+eKuln7+IwBo8zv
agU46s2bP8nL9gQ0iK6pKZnMSqley5G+A/tyht9Hh8OmoVV+x+NQPPg2XiFiUZJJ
+r/t/mkxc/zbBINvv8yfcnae0fnQJ3+2nIUbxaMelf4=
`protect END_PROTECTED
