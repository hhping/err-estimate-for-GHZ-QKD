`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LRalbNgzjKeKnWnR7d3G+oYUMz3m2iCFispTonzxms4PuMSinMRqkAPFSFG5Hypn
Dx1buv0/GD5XOOrcZhA08HLYehapwZ340MGkoYi7V/hePCwXmZO8Jps1mzPlV3ZO
OGA9BGLsrGjPr3jNau+4K1qAh2MswMy+3XHhtTGldnK8Z8lzCjyavLOs6s59NWqA
Oqw5cuwbnZbm/AnoDxvqjSXmTNIlqmPLLDBHz4JdEuo9etOWwJ/os4hQ+DvlJDV3
dBE7gYI3lYPQ633cfWrznXq/KaJLTrURC0K3wEjBSjrPguhstrS4k25VPqc//0wi
ZzchT5R3eQ0zKNF4H4tseKywzW1UHYyy5Y4uQ7e8bU0kg9Eisw5XdZNSto83FWdS
IDXI78wsnjIi7lGqjhfpLQNoQiF126E/5zi4ov6gs3Bi2/6gf4nGL04AuZcM09tI
J3FxbP1TchCFsq+Fq8cbsAZad81EHfwqa0j3XT36eOckiL3c7A9Thcx5SqLN8wyh
LuQmjW7FYfOMRzZrE/PkWqt2gGyxl06SyDuDlpRehFg3H6pmRauIvArSzjBJ33E/
Z5z52FfmamIp5orS2JLOCyNwz3GhbNQWexB6UKqHt3BwMmOj4n2j+81Dy3EBWnjL
/VO09PY5Zv8ZQy5i5QBXIQLt9tpqaU0M4lHmgrBu2t5JdrwfPMbAAkzZBxSOu2ke
0nPGezOhCkP5tSSBmtpocgvCxvRl3adQRT7LwVNJmSJ9oKiLpNqbfwmhm0szxEEx
HAxypBEtwHbMe2nIBdBq2JyAygJ8nR0K/s3iyW13Z+yEoLLHf39iROgbHcEbhkCo
yU0btA9i5Mi3uKnd+tEnCbZTpQYnpX+BYcHaOAflBFxRBMafGu/Kp9U/77+kCLLu
c0f54l7pYQa7eLzTAIzd04I2oMj/vo7SweZmYINGuKfPoRBKHcx3kBveiht4lTgF
nCqR9ruSBKSzFYx5EFKomA2KxOWO+1Uz1q2kqSrQhXL+ucPEBt7271+BZbQDPuzk
tihlstntnAgMGylRvUAlJAWxBleiYelQ4gUTdDghUoFbpCNC48po80LPutKZpwDt
9yc8j/1fWZq02J+lBmn745Qy60hTg9ktDZKAXa2tVqbMvJZ7WRcn6+BSOx+vLfMw
0tiGI8IfSJ+8nRyUj/H5HHwfhx0PCStoLEOg3X72edredEYZBlan2ywd49CzKdGk
DMgfkw3YCwAUhsOalbaY2YCpJ8lv/Meq7+JxEKC1oaszHI4jDJrqG5uCaPs6/7Yy
OMfIZiOB3lfHtRafTyz2IN30WpY9Zr64HeBCanTxuh29pSFGND+TgDTzvCTlFimU
yBXXUBIO/HbvmbVMrodqyvQGRtqaniGg+2edXGKQ45atiANpNFIHztZUVFWiyvOe
Wjg49E7GEjp9gPtiHnVX+qiMxodQ/2+si+1VcMq+4FE+ZxrKhJPvWVsY6Ye5CU8R
hbkNnMZKSJJjG17v6DtMenwPrOlHcrvW8FbDgyjTRORQd3d2QtEWb1k1wq9mJwLV
FIBY8tahW7RnmNwnO/pe2Qw6pcdj/TCQ7mGySBffEyvzv5+eQCq4o97wo3BMkVzW
pfsx7uWfHeg5VxraXqwWBajz2jI5iXOAIVTv9ZDmGaaDjHQqQsd7Lb2ulgvasF0X
f6dtBAUsvK3rDv+0P1bl1erqNwF+jQit/qTBaVlvK4PnlkEarpbwZfWntf5kBrP+
5IcqWJA9LIdUDRa6HO2P6ppLyoflQmVqbLOovq6c9XXvxLh7cAjZGmvgZZXjzE0K
N/dBobclid+Wgs4TMPF+rXmaaQgIGDjnCOW1rHBOQCdjDXVKFRH3bbM25wqzFbfX
OXst9SVnpCVen3RdfLQP29DNw/ym4JCoi7l9hcUkDVsYCzlZytomTUJVrwcxULzV
wa7IkAhq6oHU58EfsEIATxJN13/Tew8CLG2VRfIaK39Tvw7jWYqD1gABpZvGeHf4
+UhW8GyYrSsUxiKAS2kKXvNQUOMR4EbbWVCUQ6vewiXdvpSV4pSpWhTTvwe/6MTs
rf/3kkYLXjenYYV54IsjMSiLyi7+P3KJqcBVS9XenvqsVL8sdHU+RMftcxbGBvaX
zNS3oDrAVvJVbzMsxLGDpdTmBZRBPqdRkCsMgUPMdjIkoc+VCEZQ297rXz5JrtK3
lY2mBQ2niSj7eMK9E02VmV0DXkvE9JZncA0IKuQFtjd0FCTEmpGVPu+Er3v2TC3h
I28Ilk2AEZ/jVPGdIvADbpXeIzf/rLNlTyEivejeGAL+IdtjNqnLrEPixRirLRDF
INW1kDE/Jal6ylFnv+o51ufIXLqXE3RFZNOyv2z7hKeWOuPHzP+vx42OnUkgcA4D
+lo0DQynm79383Y2E3JYVUKEVnVqTXwkyKMxpy9Au02yIyi3nk7ehi4Z9R0HBNGU
vVtxGulPJjcq4vd6FEMNruQbbe18d1G0VjzTu7E7NU/KSdzKLFEfQ95+yaRxNFct
0S4NX/z94sPAU3j2hPjCHOLptHfKssQqq3qlJ/FU9GMCRJoPc8M2e2PiiZVOLunD
wdDoVYhFtxklphY2GxjDbQKGxYgKN45wItBWNKOGu5/t7ItpP+Wx1q7FWFB6StGk
udU5Ja1Cp3wbffFxXPZsrvzy7N+RDDSHHutkAqJL2UUy2HISF2WuF2LjDmlz8j1k
CcrFfPYkelxnAs5SPbF1WYhc4TZtHGf4oq0leXgaaXG4pAht/q3Cb7hn9zShnEl1
49ATqHjVIoA9KyUrRZBoJRqG/gyBNyZskY+qGdES4mhEqiZgBRSsIOCcUTtgPMxn
5uhDc+KFNj5gelF+Q/eqPYpMVSPursA6Oz1okX62M3nZO+PN4jlXCGCs/F1+qsI2
8aM4NQjTcgcDDYXgmNUanUZoNIR+YhjBSSkb7C99/Oo=
`protect END_PROTECTED
