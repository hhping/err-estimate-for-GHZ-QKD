`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvXyYVBos3/wkA19ZfGtLGB/X1P2fgEjvDqdrH4/AYcVVWuHkX2uMkMlqX2SC/21
3r3U7It0/HkHo7P78JIc6lWXjTeDwz6k5VmaEAdEsUXpQCKkIAg9c281NfIR1v3X
kHDgBXaZ5hfERrpQkbcEusyDIMsmjxSJ/RSFWEob3Y43Z7s0Ll4ygPdcAIdfTXSd
24mnAbfDpSFGUw3CJbL8VexEmdi4f+Cn31PKE/opItfNCPglDKe2J78wca29WQkQ
7HvYdM1kIK3OP0Xa0pjMHw==
`protect END_PROTECTED
