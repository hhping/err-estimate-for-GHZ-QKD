`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xias4POnlpVsEBRVw0EfOp0eI2NeUUr+ckIyiQ05aNmSc5DldCRbWcBIkFvNe91
9dGhLrnIB/dMOP/EFVlVNYA8odisIM7x24FtOsHIYLNIxvEvc8GRapPzmEtXCITB
IxcbLN2jnj0m82aJb54aCwkqeSM5Ll4RZhW4E/yXfLW4xYauKI+918sjnI+00jxS
bxPNZ/WrDmgw0AKY3z71Zb1eOAsJf7Dzk3voLP6w9Uf+lqGmUDDas8A6LmeTUvSS
Ez6qOF/fyoyE1eYCV/Kf1I2qdG28z0tdDCma/W0DPqLxZ/WIjSfGX6iw423qDLf6
3aqPsxQlowopk/WE884sE9+dq8a3EHutnNiJlvYVkQHCo55RpDdU9GTD3RDDFsJ6
JLMNh4q6LtFa5XAcuRxcBHDLsq7iiOmiNIRFyTtTadd66jRa2muoN9UdHf4OkgxC
ax1MB8h4iOhY3nRDaM1KZTJjnBrO9PvxgK7/zU3j9owsVgblCj5MWFxQbAQkI37d
SdabupN4fDmceSFRgU080WZVXHv1Rib00+/wy5rMRQbb4cDboIjMMRB/HMfaIFo+
/LyWnyFkVX4gecLD8JrmT+5Fj5e0GBHVaOBKgEjSOehb5yg1Ii5/9goeYS/yK1gY
KI1zx/ZDiRF/FmkJwi273ZJ8d96AmXjFlbfBRSCKPsiHlDjMmZOYMdIRh7tqoe1r
dAZ5Jv+QH3kmd43UDxn6seCNaokUagjq99TyYOFTsfad/gK7Bjt/9eubwNER1VGH
L0cDlfsRFgDIuQbs+HIv4mPXiKm15mTisF41XnXJJWuY2PdVtGpbIMZhAU7vWN78
IRi4O6xJWqVZ5/v2Ax6aMy7I4j14Y7kMm4K5kjMqQRQzd0FHPoTv73S1Ti2NYBNA
nvndzGRFSoBHe8BeaBQ4yb/+EmHqsvImHCEUwoufqaUJT2w8OanGjAELSI+9u3k8
D3ANeOtM5vzz2JCYKsCpwZ4NQIvbaiTeB2cPFMfG3jUY5FxNwLwxCJr/daInqvkD
ml9pPVY8igd51xTPC0lhBaMLtvraIlVYa/ou96PbEXd+PdLoAlUp/6EJHqfMDUZN
piD9tQHdGTo6eXtNqY1UzExNpStkq7QOxvrJ/w2+aS/x98LKWmBxyla+UKlHLPQy
cdlgrW9Pz+9CmATXWDxOwOi67EDK5qlegjlxcJDfgGJwDvZZ6e5XfzkN80D9gUmX
n1s1SFlv4vUPlq2/2SwJrpGEz40LlIzzj0shFpIElBA=
`protect END_PROTECTED
