`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Ot7Xk4HXtTEptBhAI6vKq4AiPu3GSpX8kJegtze5VF8b9wmUWQeCgVZjs8NbSbW
rLB4VvlvfltJ6cjBweP9siy5BW7r5hfGXnX0YQYiRKtXnmOjHJ1Ft2puZmByO50q
x4hbl6iT14AD5WJYthj2MQci83z7Og9ZCDa81jnHW6grqNhw2f29yKCi4fzqPlWX
mn+BE+kqhfuWJbixFNte701Xs1BHQIO4vT3JzTV4LbjDOr8+kKFun74GaZXo/SWX
tgQw7z6hxqqPHvx0oCXO1mRHt9ss2+HbBtFYaSiVnsWasyDQpYzRbcG8uF5o886j
XWapcJtGPLNotXbDov6Cl0qkuB8ynH5TsxnxnG9VXHL30/G8PwcwTUAthF64Nt19
`protect END_PROTECTED
