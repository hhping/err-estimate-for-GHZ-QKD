`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rEqkC5ADKc9VKrGYMpewN0eqO4Feyyn5lmq8Z6rnDIDjU9gZMhmRj/EWisYTuh7
FvMmqVROJz50hOie06ybwyVfJRDrAXdJEEELHVlZVxO5Len+BjxIQNTR54jpw4tw
3TB41l8BFwlhkitWXeNsgHt2gJWpsZT5hfqrGbzM/Rk1FlkL0fvG++jlaGTgxbZ7
HrZ7duENEu0uA5PFpAY0CPQPeBDpWJHUbPQhm+WJG1O6hTnUQADGXefusK3P1QLR
C6SF7+jMgF4I3N78vuK+TX2BmDmwo172ASI3BjzQIEzX1gT9bW4uU8iNE3QVYrE9
7eK6/sE+vlKX11Fm+bSAzNhP8CuAzukyUhTIwHv7xXdNMb7dOtqBxI9kxg5Mzuww
UztbCyTZ1VH9XVkRTvyCQHFnuG3z1inJlMdzA9sUw4eS3OOzjXyUSHHVlWdeKNcZ
`protect END_PROTECTED
