`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3KhohLatkCG7O8fUgxCzIoRKzxCqr704pRc3MOQiOtVrv3VsCC6W1vkmuAqoFIWl
NYpbOkDg2fID4tUcWyzPlJbK3406junORcweSc26pUx7R5dc4d68oZcQegQXhQ9i
BfIVM8g4rVBGuy7kCI7I9og5vLX7HYZj/GDD2PvSBN2XN9w2vhgf1v3au3rOdqu6
UFvB9Hr/hoLGWLlHWb9lDujSEvp6JzRX9SMJ07nRKe+EXbFn4pQjhro8q5lzrCH7
fLPkQtqibKLc9K9SGKSUEn2h4QJAZ5kSRTlu3+o2YRKa6653ibkMfqv2l7TVWRql
1oNli1zam0+l4/XlPLXjqCi2w95mO73GTTl5vZuYMgT79aOJWWLK2FFYaK8keBHD
3EP48A67MJkuzwamPHZiowD0DWl1z7x3oTd2sRKYz2vqmHJKVAbBqdZPshNjZLyF
obpiuHiFns1wHrifALvydALWCPOFtIZieTAOpuaaithxZ+qzC/2wNxv/dNKh2Wn/
2KUfzvn5oJ+56yYYnuJgoOERgeLfbSmyikl/Gfd2NYEiGzBLjDL/Qqj71RouXPL7
Umv1bXOhnFm+G3Ru/UnRtvmfCM/3EjwJoj5mlvZbSKvGccJXdYdR3mgNAdi3YImL
9EPWIMDDQPQhesOeDdgrfNVM2H1hCMrhppRfEW5eH+TPw30Fetf9gvLXXIvsONRd
Pvsz3zMrsnepRWck3Tj6AiyGrV1q25dhNxOY+LOp8q6v7pGWo/P3AVBS8nuOmmwS
irm7gVfocZrNpM5b5CRM9sZ7TC9Q5oOAxEYj999c+2P5KO+piI4LS0FvzAPC47G0
2UZw8fXuaPCrBjYbd1+TCMJzZjvDjy0zlbMVIdg9vILrTmUls2tb9e0jjPCi6KGJ
1hgjknQsguETYuBT1K0i54ehpX605GOzFR7SfO8joW3pcd6k/tGk59dfB5/Z3/MN
wSK4PRFRJdNtdUQJOuyUX8tXOPnh7yBx5AiAd32rMU+X6YgznSW4fsWx7cN/QKVX
uw6VNOpsw6SKiEfZARXMCQ==
`protect END_PROTECTED
