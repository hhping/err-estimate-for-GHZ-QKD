`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4/i+sAOZZUCG4FaAM2cBxlU8XNhnIAzBaF31+gFh0+d47BhPZLo3l6RuJxx+IN3
CNSl8RJl4lBRxv+KG1Y+/mse1nxuogA3SVxdxoLQIhx5uHJO0AZUtPYqCkBfHbbF
leSCQz5IWM9bxgjS5wLrxsY18fsI/1RPhuzhAV0q7vEVX4+uTDfIeNnOF+Vv/0eb
chyLRUUKGISeHeCbJmYPlTyp5TFtku/InfQqXyr2gmH4J6JiDpdvUD3F2CwQrqa1
A0zwiI9Ms+NMR4hjzLdXuhCqpgndFmKzfKiz6iOOvXtOSSdRXr/uPM3dJ0hBQt5d
n7LAewY/BySJSUlVVMRcwaMiFRfiz7NEFYURcoH70LSSKoXWtsvRgg/mEJE9dj4Z
T5jfuOfjUsoSeAurAGUHh1dpTE6eY+nc7Jqdb9lht4qoW2MroAMyTBgEvGrG8drA
lnfHl1BHMowNPEY8ZTTbUYSgUCT452qBWViphlVfSjj0Pc/1A510iJI742rhSHib
/sqVDiJtaVqrwAv+JpHLYraBx4QAdQmRI6YgLumGn6V8cVgcaOvwH3+X+CfazKWK
d701XL2hET+1AFoJaGjF+W6ZFff5KvJOQ9y63E7NxSDB6L9wH0gJt5OR6h03k9mA
/zAcPTbV/FC23kHBfBj78LNjiAbS6vPVUI+zwoYythc3Bfkk0R3miLz3jrufQkai
3i08pFVH3HKibNTxGt8cMjwNn5nd7Noud+0opA7MvJtlfxZTpTaajH2BR0SS/owP
BrEX3ZQuH9ZR+KlKbY8hc4u/4q5ecj8nmZ0j5F5YXAuAEYU80X/qzEO7UP6YxOaf
VtkmmkAcI2oYdesIglVaVGYnZ/PdTRl/ZuUrtM+FbjflOBmdFbNP4elmRcT6rAe/
zJcsZqWxbLrnd9B5pOB1rQXYqUzSvRt1oeXFdAVu3FkQ/x47w7kHY6eydE8LzjPa
hwg+ArhYw+Ny8B9sVuG7lvbdpNQerDx/QmMD56pVoLzKE1PPDX73PXpsxMQlo98z
fMHbkSfe6Nfsm9aXkeQw7Jcj7TRQvBnLdbF+2w/xD4Pp1NZ25WfXJWm67YMynjVt
X3p62ndhle3Rt4z9+Nm30wG2LGcDgf1iJtRLjgY9DoYwDBxqI3x79ca5IdnKjK/e
MvV9EF5KHgoO2KR6pzPN+R9rjqYuNSfXaOnYCBPnoN/O3yhZdUDKzy29kEU086JD
I+RY5Knz4r2c9zCSWlaNUPzKm6PJmA7yHZqKCmDg+Bu5NuvfTxh2mBDuckid9cpS
DFNdbFXUqcX1ihN/UYP/eHOAUX5e2t9DTpPtWo0yXUH54u5LNtcYZ71cWl4z1pTA
yvEv/+W16BoZAbpr5sLIOCPj8xv0NIeY/uOWN8bpFgbUfmBb92OQA82ES06Llv0H
5BYTNwYDLZ+wInfLMKAaoGQLAeZfiFNqrsvVPL9OFpblfCF5kiyFuQuSPJIgrS9v
qx+zDhrJuos8V6FtB2l/eVPXiRRP4YMCu10ziMeMAKTPngakM8Yy9tMdksPZdkyj
/ZsWs+Xxp7UoKXPbeNeKCQQQSKFJ2cRTeX0YIXxKLywesiUCZaQSR98y7WAQWCDW
Vnj/s/3VRyrCe5rYC30AGkgP3uHY2p2SQBQ5KfO6S5tVHeDdvwTAf5lvGC+dtg6m
UALGNPXrhf2r2ych64xfnRxq9W0KojEVC6BLbg7DIKQ0udNRc7xmwhrABnngIBNR
2tJfLG3DF5rnHl79Qqs9IpmmGlsrKMtFriJmuDFp0FU/rvs9nAk08PkoEhoieTqf
w3fVL+PrMeUjVNQhom4ZRZPSwEbX/lcVgHikx2pGyAbytufP9PBrYOj5nJvVpcrC
jMo7GWGRoMaF+2h/Ty0OOTRdrzInSRfUZL7dsXXHxN1297VoDDNj6hsmeAYlungT
gSXbDU2BqATN/wQnrZFRinAz3k3lK3MUISLfWHxnqvY1L6bep1rpB6L4PJX2gGY8
RKJRUH5pVMEvm+SQ3sQtCFv5qMrhXt8UsQHsweOf5eXwIMag1mw0OSCQObI7ahbo
i3zapeMX5rGF9YaFIcymeuR3c+P1mU3o6PM3vzbZqcFCSSz7qjCEX7oKpyNmDbh1
kgNeZmxXpAMwYtc4oq/YYX6Cf2yCBFj+zgXk+o08t5yIyoCS9tCPQynigwpE6YmJ
339rZI/V7UiuP7UktzkdsomFlfmPGal+n+G2P7HBn64ofdZwiE1fU+oigntpuxh0
F/b/P42jYfUmuZZ+6iRfK26iZacOzRVuwCHkgn0aJepqTVcazH0XWO3c7eHz9Otk
mt5sto6MIDzNkksJUNZ9CWonapI9owvl/rFfRyoMyett/wxx3xYWtLtSG62t2prs
MI2901tq32xjpzHVUj4CQ4O6ELuOjRKG6rmGy/naeD7E4YPXgsV+UkdpnfYIcdbx
rK5JAgIf/q2CoF9cvPCi3MU2Ymix8/ESFHBjj5TSenm9j5fIME5E/jzpVMfvlqy8
ckAm9RY3b9gdOtt7nqPNyW9Z0jseP280UYcUnhw5yxWKygfDeN6VtYBIGm1pVz08
9K5YwQH0lPX5QDzqe07uEDhqe1n55ZBkgut1dUTByqdEnBI4hqB4/wzp6dHq1Or+
UJh5DaKgYe2BH8sAGX+0rC/krUogFJJf0iNM/5jQM475QG5Qu7OM5bwS0rRqypce
MQfx4wHgY2Y9GfADOefWx5V+ZQgrBjaRskDZ9u+VC7VL6OSDE5DdpOUFAo/fv6sG
A2G1dCA7sjFQAFOhAYO+P7BtLKbImgFdVWBpg86zwuU1Fa/iLSq/lG29LbDU4mLg
nttaTvqz+tIfppZhNV9P3J08Pd+5GY0eN6BYajr5e3OT5SrXKBtWQVrwyVGI0CPh
wqzNwgdbh72A3VvmuQDeVAIc/UWdyddEixqpcot9EPkKdbUOSOg0ZhbP+z4IRvnT
gbFCFjpCP0P05fAf/RVVddNOAQAAP6DQrn4KEvyZLr6gYFUWUFMJu3rdXxFf+ghW
yxNsw5PNDhbQIF8Y360RQvjn8m48bV5oE0t5h5SEn2+xojsRCn8I0yNIeEBHBzsW
Z3IVdzauwbkW1S4CN3GCdzWE6xl4zWfH5VRT9s9eSXfidpUH9C6LeoKlm8a/0Bgd
QWTVbQTTPlOsXTeVO6kOS4eo0yYV6wnPBVPuBM+tABMzyMr4uSxUugBCxub6HMw8
wD7XG8XKF/9QYZo2XHIDeAqqM8DXSp0DkMKAtpwUS6166+U4ocz3usZy7Lk0l4zw
hkmfP0Mg6YLi0yxHq9+KVHMzPK+ZXq76XI84o5aHS9uP9voFXvMDDSVtbZfSBywq
gpKdLd7JWEnbgf/8kvZcq3kd9xYXj9AkR86f44NCuzzVijRnHpGAPfmr9DWeWvAq
I8iTZ/aAII4E5vq7upP7HW7t1oUjj7/a+Vdrv3x82qQAWlrHXh7bBCZnGi3sMp0X
d5K2k3/nQFytp2y/kfg53MTZP4BJpQZoy5HLL/GyVrOl6W7KfHI2ryen+H+3gOmQ
h43U37fA78R2NdW4dqUO4cYyG+b2fbHdpGDnXKnmiU/ff06Zrcobd1NF84sDHa8G
VF8cB4Hf22bgl9sbsUBjuvNLKiTDyJiMLO2JihGkIvqK+PecEnn5TavRL/zLPfoE
OeKpGMlO77lEHfzIUK/WAz3+2v6+/WDOQazLtSpcpDR3bd+8hQUkGfJcG9NP3aF0
LKdrm7pwX/YjvDt7e/4cAWNPPm7yOY9jQXofjxA74O/Fyu09TQ8veltL6mjGf1BN
fPXReA5wFjCNQ41BvRhlFIgovI7WzHKhDylQdkXNyHfziEP1k1/v2s8XbGqxzJon
0fM3B56XPnUnaqxSFDsQUocNzaSXDYkDZDtLcFlr0MO1RxWqkabX5ZoQhP8vsSvh
EsxS8M10c5EykGsQOZ6cgdrGiWwtx3hJKT//pRe27wYnRTapRPext9qo/8N7t3bE
61GL2LBoQxxSEmvJm7SVBc1B5PsRyxPRME/YnlG5xhpBV/juP/mkL+qGPH/yx5VN
BOEXQaDbWaIljolbJkEpDUOtHejG8gmdmsclMCyz2L/iMCx5t68fI0Y7CEkwN+LS
9i6IkCYptZO/PMl1jEuZ8MG5/jXFHl0qtmTSsabCS4R/2Tc7kZ7UScO+vrm9mqgO
Zqz/JJuEm0VVMNWYhIe3gCeSEcZXiKv9Fs/yckBVpY9nX+Q1sz3rZWKw4I3EIxAF
btBTK6Qx7+30wd+fNdMV89T/3QUnCKWhVsNhPY8b06IoIh+ZRFcMy22l8gSJCSy5
mSfL+B6NJlJDhWhwKeGEqB6g7V8OmGRXYg8cH33Ql9hLgaIoaUR+zIiVmZxE/R/s
0hCszGIsfc/UEgCzcj00U1pTDxXbKzz4KxT9WmzszA2/uPeo6ma0ZtAROjtuIzJa
j9cA1BOr16zNaYMasIJfAT4XZPor92P4Dz+srm8FB0795kKy7s+ybGwc7X9Z3o/6
Z7HWFRnGa/EkAs/WhPs5mbTD5IiEwyCddDZlzUwLVCt6fd1g3jzkK8Yo3MZ6nOdk
MEkzKHQ1ZFr9Ku9F0qW/Mnn9nzhyGdXXSn2I/JzWNPudQ7fGZcmyyC9ujAMupA8I
I4Ha/S6f+OHwmFR50dvVcLotoIWAiE/1uGIVhHGOFagpMS6Q/X87cqJQZBe6f/zh
34Rdq+dSERFe1UY01YkqWjPZMGnHh/LT07OKyMSNJ/saW5HrhnhLs9vDV0B8A3OK
VNFbGKiZPrjaSVc+fhbrMkrRYp2o5wTEkjCKgRY19hheNTEilLXxzPHG+uZSj8Ux
j9No60lHmSm1pdip1WgX5JwzTFo2Xeg7SGp72W8llf+Mb0tKpqjrbzYxoAdQXQYT
GoAMoLwnL0u/FVaYVp9kWverlH4DliSbW1EdcRx+XaiIxPqbKDhhSi0b8jK/ViBm
Hl6Hhg9tuXGoi/+nDVuftThB/qcUKf8YXxA5M40i/q9cCLdNa4E9oOppJw690CCQ
hpeLXwf5L8wW7FQt28IQhvNqA724qUYmPxxEXqzKKA3tcvVqPDgb+hSU5E/vTtJl
qdU9H1QWQFn4+qzl65giV00G/AAPDsiFaGziZXXRhiVCBC0ZBhNAIuhzWS3oioRA
mcKu3B46wkKnmBNdLBy2ZNLy82kWdVUuNZQ0GReO8PxiQHgUQk9tc+WEEqytT6GW
YfOA/iSMgSfqgLcTf7Jl9vQHTtwKbv76b5LrAmDQb/ckdClneO5kHZwhURhBi1I9
fLuZ6qmrtZ9A2ACAwXyUE4LYwf4ljuiRWzptoBPM/z7P1/lJ+HgGy6eYhkhdWXcg
J56t1di11oezI4Ph9IEqOBavGu/xfEpGZAqxtoX9DjZVO3YbjFFxwvMhhw2ITKi2
qSdcpb6Zw92djRrUKClSpyBvepnk2tMgwoLfm41KPpbI+nhX/zuECem/Yzw4clkJ
7x+qrhnHKWPlo3vSafyefdl1t9fvtjFQ71k6MPL2wWeqIHJqZAYkwNzVjwRsqaK2
hXCy+Wu/Dzt3FBnS3UhTydmUlhdFuyLBBUpoc3KH6H5NsKaJrMO2kyw1lnD34kMu
NcqoI7uWERff44qzwXJzp7CvfFRjtSD/9hsIzEyeORIqMllscv/ztCU6aWKkFr+c
x2GRyc5qD91s+LAgLErS9GSZ+6fUmstVnCDRd7QEPlPBkqq7j4d8FE0ctU2UyHdY
lJzAV3RUJ+oMREqfep07rHy1VHgWyp7yps/cxX82FMW6tj0hhBW2ApaS5P7Me41B
HLQ9p2vKgvQpZzWvfGRY2z3FXq8MhCgYV4gQpdOnRXf6DsKpXfFgDTTk8GsMssHM
x3FfW3mDvToNBBlu7AdZx5wpm4S90G5ix4FgyvY8+ViJs1s0E7W/VSZTGC7OC3em
TKQL+eVOcxbAdhlm+NbxNvJrHLYiparrCSFfBKRDgV8=
`protect END_PROTECTED
