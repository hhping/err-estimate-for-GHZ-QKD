`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
plsHuIF9H9m8SSckutBkgx4KMzZpvdNuIPi0GQiodzzpR2iKl8BGQU/baKvhOP2F
dRzqgNQ+G+NxpxGhUdyk4jytcfI/DVl7GQ9OXYFWRQ64Vt+JcUKeqGLgafqdDeZu
O/3JNSIJ5Y8Nv5ylXvmAH2ZEYG75IPvcUUsbaXuoPQO4eMWF4iSAt00blXLiwHU+
lwQINJbZIZAcs5pcnoxM3H3Yh8EFvt58b4zbCGLKD1visnwuz8ykQqDx01gKr2F/
pec3gQpn1yhDFkOWVtxn5BrjmSPsqn4RbGn/3ynFAy0z4HKkRmIpMkyFzr955LaV
TwrU92BTcCCBQ3bjpwIoo35LJmXjo1Z00hnZto3nTHe+nduzKQM/QVd/VyWAxmF9
tzS5Acpg5lWSn6UouIW1C4EGPgT3HQCLiKh+eaWW/HsvJrJKMiSsNsbTyynO3GfE
whIpAZ8xdMiCbFDxx1QlsrDsHuSgU8MYLEuZDhdRD1e6E6H4pe8BSTZGbEk6b56l
oBN4YXOQYQXj4MNHhleH7qgW1WiwVeAcs7DRpq1BU0xarcp3fyaRZfMvD6EUp5p/
1rkasc9lwj5+IhiCrpMSkqmbf2q66rD21q/ukZ+lqqSflPv0ECDf/YGoe7FwfOEX
z/Mk6OeyMPOLQHIMuMUdvJytHLWm1qIHv85G55i9oUndTCWILVF0dnSoq+ZU1+Eu
+Nqrb0vaHYIlArKOWEL6QhNcqDv4IHBsOvDWMQ4cF+k0iDQCkhlqhlZ+9saFL6VJ
x42+fz6Qh/LD6wCIRyU3VODBNEOVxw+Sb6L3sNsLmvyzknDfu4DOTU7lHm2TWHVx
nz4ay1u+YYK/tzRmCxUvYjL6WQYzAzLWisZIIGxs/yKPVlXuihgkb3slUtpqxXQy
qXhChOUuPc1S8AObVPwt40/gyUam4CgtPq9caSABxEO8mfjVh4QYyAVKHINtWfXI
g2e1MjYNO/MBAYk3z5D4TiYAd01Vm5Rt+TbCFRtYegDXOq3j4tEGB6fPvetVxGom
TIfTsG22uQT7XqLIl06tVbRdYYRSOzNf+RfCuH4FjXLdOSAieVYtElyoyHhNU+2m
mIu+n2b5bYMH+Q5GhHFtl8aRN/Ei73WPJrjpDKu2lqoH8SNMwqpUM4k3PZgsmJnv
l7X26o0wSrgIb5DlbhoM53Z70RoXU9q6lIUql2RgqkFavKymyxfvGXD1m2SRPVCO
C5uR5723sRfV+xnBGWBopq6zRbwtaSjWsWQlupM1J44MRVJuT3Vs455+53Mc6v/M
2Tfo6z+wNhPyBeopowkgB4ZOqMTGgI6RfejfwaBVCKe1JhrmWJ5NIt+lKiEPFQUQ
+n0MGsq92o5S193v6wgZGXJzXzaiQ2JMssOBgdsCkZjIjenvy+GP2WrTDAt2BC5j
c+dkIWj1Yi3e3GocN9pMKZY/JjJu5xjGNuzz4SVBoMxADlYANGH8SZ4o/fNKyhfS
T6gvrcqBbmxq2dKxyahVPBvmotiTWUUjaZM8wo+scNO2wL4Ps7NzZGdGaqxWmamR
wnNmo/3jhDsyl3NxoN6HAGJv/wsDx+GN+E+Ys6VvAkOVYVckHDxcyg87UJLPQH5i
x7/l+Br3IPh5cP25FKSTOAoxk4/A9ocA3UThlOX8+YWLrpeBNgD8vvUkRUyKnO5e
ss9jpcHB9OuHtXfr+07wtM07H5lqCKOVywOQgMD3y/Mw8GQDR8CTKJl67f+MAFz6
lwL94Eh+BIUuLSTJMifvS5FJA8NVtz43ZjlmbYtffHQlYIP6/yXs90Mexmw8u36R
ASKzvD09IQMxU47RJNkKIeY+QGKKKAXy3htPcDsyy+rhzrqF2hleoWTM32ai8bRx
wiq0G20e2EpDG3aTlM+biKHMK24S+GK7x5qWFte1HkvFRKmJc/6q/TJlSQtdl5Ud
h2oMl1touTUiwUYWarD/fQ==
`protect END_PROTECTED
