`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpgPZ9PbYB/vWCSzGcQ+r3WNU0tosf6lOEKT3Hirz/dydI1zSlcaeZX0xQzEWMhX
BJC75TBmMDM1Ro9fyIVxHmfIb42se8ypdh24Jmm9P3q4Tm6mo6S1RT7ESvEazor1
6IF3whWFFbfoJgBUMBhqLNk6U29uuDr2yVhwd5Es84xbMeoTuUdoK9OSmyvj6qup
q9d3JYRIVPBTvHu99tH0+NWVhWlk8GodvzCK5f9RQ1irnVWIUBNbeLcGoWRK6ftd
88MIHU3GLCFicVBuLHq/MB1sYFEVgrf3jd3qPZ/5Epa7ZfO2fPwxilUjztrozBY+
E1c20uP01LVF2mtrAfmYjvnjxK+dvPb7RQ6htYtaeIIzS6eSxECVKN4q8U36qkcf
FNNTHV2REwE/iug6tuc0cKPFyIM8qNSqgZ+Y3BwbcoUmv73OxY5WfBtltPHz3de7
oouyJkwwxqTAm1wNIeVNnQ==
`protect END_PROTECTED
