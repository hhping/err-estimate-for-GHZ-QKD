`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vnGLlWO43GGuSViHvoaWaKv4tCGvzC1cclvo0JEzpvZMpVwqfgfOXWHqfnkv+FO8
mO5ntbIn09NvIawQ09mXnUq8/cRk430BS1IAcEYfNpzy4HdqOjdt23GzYfuT72dx
oECdd13B4aiuRynVaNb/pKBKdokhRx0amzpeKu87j1ey1Su4Q5ogaLJSQa1DDS8W
RFYcvubv6Xq8z4lV8VPNwICjr3q1GK53/ID9JhM4kUEJqkb8acmIlEKlSHEGmIsy
sbK6ekoNhk6OPd4/qzc5/xnZfYNkBMfEH+gs6eoMAF825oUAiMD1m6hiP9ExBNG3
MzZ9Kuod8LG5w8Fws/TVb20g04CiGtpJR576jtq9InunMS4rnGkp8Eq9eeIz584j
WdWdTlq12OKXWHFOBd7YPGw+wlsMkHJ+jH8mU6QDdZWg9pbHamqd2kEYJO8AU+52
kDhUWk7HnYfakBAvs5tRZoWoGXqSYqDh3g5JSBm9jyTaQnrGPMOg/rASf35BkynO
WZYMBACtAB3bSDmJGd3JSA==
`protect END_PROTECTED
