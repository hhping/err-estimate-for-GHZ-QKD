`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22QrOF7a1OWy/2rqCmSWSKbwgn8RSILhChV7cpRxLkyba2vQHWzrBhGhwnsMq6ht
6zZ6kmkhR0IqxxigMjhaPYKjm0AUBA3rmv6wjXaSOegdGwOErhdUGvaaTbZboeJH
7UwIiT9+e92CQ0FmT9JQctRpbsp3Bihz3LKXl5cwSUyB+i69Prt1qj6WlRV9nDlV
kTVNoAV5gUPBOQgfFv7/X6/0KhuBb/bf4uhVlo+cnPk1sg5lPtwZET3Vq5NmYwbe
Png77/wY2lVlBokHt6oIYGYSrJrIvVYG8BM9hShFFBF76dXpNh4QbD2tOBdsZgbX
KgTsGTqwTY7CDcuaiHYswY+Wv1OhD0mB67msefDfhj5PCqTDeEgxY/aX8KUf43Vd
jVMhvTDJVrgd9tsdqvuC50MxcvJeFuRbJTw40Ef7hgKKV6v/0hnmd/ZZqkD6IFzn
0dEh3x1IBHD6xqoGfbrUC27hbiO4SIXEXRE3YDZNn2sQmS3Ddi0/tTvyNjo8gKC4
rvsZHJHXEiin8wB6DuR/F/SpE51w7a2eiNwNIFfHdXwu1vOoa4meeBrh2ghJP3tf
mivgjIQBD+xSvef9lkYklzH2s88nfROpRTjFRM5dH5Oog/I1umfF/O64I3mNc35H
BgXWoyo3CsXZ9YJPXydoHM01+ytYP25sw0sSX7TuV1E8HiG/MVbzWwHTrVrwLnhT
RyGSjoryCbJ4wfpZHWVHmVJkgUt99cShSxJ6PpogT5Etj0Bt+eoo8baqZTQERXHD
Zq68UyQLWy8omVMDZGfHaXUnbIh4326WWxU5PDnkTJGYSsoodl81RbuWM1PHGI4g
PzNIQB52ukWohA21rZxZhfVopNIzu9qetqCBWfqxjAlBnTPFjkxYaMAia47ZLwCk
4ge/2pFj/B98yLJCNP0NCu3FP6xx5yxCnf5ZxGvES2GGPB2xxDA91b4A372KYCmm
EtcjGZe0iaZ9ymEFINdKgTYCt3VpUmcQRJuWnxmhubhHt2YWqvXEtt3Z7hpksGjD
Oi4m5r/vdVOOs5RLZ9e9E0qtMjwIqBnXrfDoZHrD29LA71Pwz+Em+wFAYY2/qaBy
bFF4U/VGEq0fHa5CHyX5LL9vwt3kpj2855UEdVc+JJSwyHuHB/aCHFoyRUO/EQ+O
PufeipG6a1Q6aUNfz2Pp1WWVburjbaHRpVhNBNtRxkBA/qPopSotl4WxdIIR78wf
CPrKwgxmVXdrUSvp9ikmvC+HTZNZtJsCzHRVFbulQEmlSTs9adeXQI8/Lj4QoAeV
6lBuS2tBC/pGd3ZtWSlPU2HZ8I+xXrgge75BrLqV5RmVGjwdQHv7ED6xuQ5JfmuK
+rWuy5f33SI0p0Tnuy5+NnEhfYUQqQA3R8a5hGgNDyR1E8yHnDGcwIIgMfKhBmG8
TaTpQFMoVgCFsnfhZkBX/+tyn19AkmQEFq2RJbtgNXrPwyawq72BZ8Sluj34h6px
gHoPDg0Q/evWkV2PV8TMaXGIG0P5bi4dJhe+dVuWyjPBwDPc/tk6+NpWqFhT9TsP
3RCP3WEF01Ln2uRt9vW9YqIsUIjmu9Lx5j0c1//TYwnMvfnWt5TJzfe8fGLRG9ZH
SvortKAUVG4B9Vk8HcWhk6rQ04AVq4j06A0O0Sg0jsMREKFfys/8eUxQ6sOhfxNk
3dygb391pDP7eZiQ/jYRFtCuAGKcdRGbydeYp8tiCXojNPpeh8miAHd9MW4YmaeD
6SyqUsRLtQ0O57ZyBoPcuKb1IfJ1YHCS6vsh/1+4jLzNCj7ANc0H7z5K1+tfLN37
yEkeBd/MuR4FPoH/uTplIXRMBqjoyyqeUktAXJr97OfifaP/eEdMZwzhKnjfWUh1
o0VWCmAsXU/W1Q/PNN7D/3SzS9FsCoINvGWh7z20Lm7ls+BpwXTMuU38cDV/v1Ue
S0zWiIOkNCQcMcIJz7ZyBOXq1v1cxdLFb5cYmCcahgEyAvvplwfbRJKhOPwlXQ2h
VcAzGXnDUs1Y1uOfFI+rokmq3Ra1fEJ6SsA6qWMq61ilLESJjkyR7qgBKnIm1kHw
e+525qdeEiJ7TDrlZV2oXKyyMYTck4GEEoevqnbsc9s=
`protect END_PROTECTED
