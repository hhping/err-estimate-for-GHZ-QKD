`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8qMXjdgp1v6iRPYpEuzZjwKzi2eNEbYWVogn1qIxvBHcoE8F5maLztkqnhg8klG
AxWKKmOCLCWURQMmCAjhzZalhatPe9GccmIgXSnm+fi0qkXzeHkMxT36ttdaZ0tE
yNUpL0VbiHTLBDmCowNWtIZNseV8ERLLSsN3Aa0mTNMKKSNmt841y0REDqtbzPi/
EXHJsXGuUHH/O1XMBgCSt78yvPOF8uzqH3oHDzODXhRnTSXBDjfyBKlO6wsoWNUV
bV3F0eZdNzaykDaAHCR0IbLFXjokFwVdbbbc5f7ltEMBvoVJ/4zOaLaX/CZN5+aj
sildqjkg09MYhST6eqnzJ1jMSYh2nY8ZFXn6JI5BP+qqQhqXvms7rag8qNpmRTaE
ZsPC6vowcAMzCC7dP6e7RJeZRa5CNbjGUgCEN1WmIkIpl8Tixx+9R3Gw6J32Q4gE
X5F4xpbCQOaHbCyb8WH9nw==
`protect END_PROTECTED
