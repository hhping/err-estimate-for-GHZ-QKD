`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nugyA/+7KyJweGdPpAanY721B1GpbHwZrfPBUaXV8UH749VEMObnLRyYk2FMzP5D
kyd1uS67TAf5j2v0LKRu+0ja9/djKGOsDj91cirkWuYznOYVP64rk3sz9XDPoAFv
I7AaM56N8oJFif03crZoBxtA3rFvH6+GuzbwJcoNlzVfpIqeU7pIMClRXFZlECys
gAbt7BcmNATJWG7fCKfeSKbRzYLIxs/8VqjJXYiZfG45IB+0zIUTDEaVFW0eW1t9
56NkAZ7h/RyC4GExCMcZRORGIdhFds19HP0BLKAOLrUy9SaIWWzGfNnhHUjwdqp7
2L1AuhyEl1Kv1ZBIAJ3E9DujvErC/e4BySbb+meK/chY8BEDsbLICOJSc+6/ouvO
hQlD8Ug4SSTuS18rPPvd/Xh46LYjWoK4c0KcOqKUzWZsXVX/+LcU7t9eWSaL7OzH
x74LC/DVvspjGM1lTGHa6oil3aDZvM4u0RU0G3QsozzvQyS/8yTnEMXt8tMjmvXQ
dF6ZMG/SZbGkLEwcU0EWZ8DvA1Uze98IkKgHyFRgp698GqtqFxrk/boTRK8BeLKL
sHrWIaCbERU+a7lddlYDz4kVyzDLMJZZd2c3HC4mkztgUdUEtjZRbr/E4/Fz5Inv
ttg+3/LMpP37tv+QeJ1vNeCMH0ubipeGvIA6JBRwGNeahh0nx9B6MQxBV1nLymAf
tDuY3Vb0cClHZzVCLRZcOLyc103/kzdYWdVSd10qgc9ZYf1prqkIIzQDvV/AEqNI
bgLKqUb/r0kXC3gc4SBHV4EXqzMqK2tPLKmPdrkPGmInEmpDOSBNiIBTvrk0grlX
62tjf+TF5VZxu+BAxgOrABOLyWfH/CiQ7RA+MA1+72yDVJtfHLkxXrDQ0pkqqlQu
sHGacLO4VKBaZ3+IXpm7qS7aAM+XaAxXKnoUzFINK5O2g4FOlQzFCe7BKGDoA+Gg
5HK6CCvRSkWgBuk5hohFTvCpaFjLBf8PE2Y2Xo6tO9C85l+pDrCDo0upHd9z4IzB
I6zv5eocayNLbnPnUG3UNjT3tg8mV7OYJHRjTZKkAniycV+AbhC4WUxof7525Lng
Io/7a3Ova0604dpd7uyDr0CN4pxwWeTgXeIS3aMq2UNZqIYkd9V5K+v7uubBDKx6
Qb0eCw1ATUnuFgUaL45TH3XxfviaWxZNYsx+uvHgSVW7M4GnWwHGeYYNXucfNNgS
tVQx+IqiSvig2WocglmMGcV6qH+3lDO7xyTIkb01gofZ38rtkKslevNWhCvUxWj4
ygi4oiukX5X2fc68UfDll/bYw3CWaSROCizXYov8GaeuPPiVkClx9g9mw5VRLEjI
+ItEIdWnMcAP4HqMBuyy9iHDlLNWcP6bBpXQ+96/O8b84HiQVROqDaSjX3tzCOvn
yx0Qdz/v/3zzuMNait6MW95dKwnBHFLG0AfiT+QOH/ufeyMYYNzyQlErZRdFAyO+
DiflK2b5YcHrhi0mtQvTDWeoMtGoWtRiCVhVYa9DrDrSItcHg7NknJ3RaTCrasYO
tLvf9HljBI42mMqJQUiu97mZPkm9xCmYd4hDEnFO/bj/bwDNansk7kfQwA1JbCga
X4pk4E6XiJbhjJVsaLwUScKcq6++5JAb99RaEbQ+rE1Is3FdPy8IEBOxBlt+clQo
HuZMmcrrXuh2ic6+/LTfbinS2yJsnmnizfuuCxLpcOLhkIvaCsuIubTT6XDKjxld
0XSbp66l4zTjVuYX33fEGRvcHVn8OudntgT8CgvBLIvyVO4s0JzL/rP+Jbr/acWU
XUis2swtvQ5BP/w7K4IVZbeNPubFVoTBKnlAXWk9rtJuJ1etYNfYOfw2QnTNWfTG
HbN3kQrFTEr4w65K0t/acgJueEHt9nKASH5W+0BqKiwnzuEugm6SifplOrRAB+PW
Z5O9JIr+sn/ZOgS1aoRf0iGNaLuZ5kLPjD2L94fQaurQuvCixU6UCEmwe2WjCT0w
GRCTW8Q2amvQXZfj1ulmUFzNrqyX6BxuuUzfK3gtjxEnNgI6ZfO3YPW80xWiIPGt
GPfT3r6xiUVd3D4FyrJYqDhEGuX+lENTvWNZZiCpQgu0bGLTCCyMn0hAXuQvl37+
2IYCk0WBNnIszV42ANAThZunBzHrV/5nb9+z6jH/7c+V/2thQMgRze72PdhtO4b4
YZQ+dNxip40yo1jw53OTVZH/Ot8aUQM4SbUOSlIwzWY6lJXRlJdvw5VijnUgUzCf
NKGayyMAiQ43KdV1QkgUNPsUEwEgjN9sln0SsGesrqvVlflyPsvwmyDVhFHIcUkX
CIF1OH+PHpuNyX9+9NOl0NobBysZ1pw2UjcIgYjn3l5uYePis2OnYMhB5iXm6Z0E
K0jofltSQHX6lzgAlRbJXwWJ3aHRkQ332yZxki2b3TIPE8xD4s9blipR762yAAoa
OLExhioByHCWTgIlDd8tP2PQrGjIXnR1xQ6JzlZWhcaTeTkqDWoCvSzF9wPd/7zq
`protect END_PROTECTED
