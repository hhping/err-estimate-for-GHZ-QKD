`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ou8PYlknbcBfay8ErZZfiSXdYwgXtrjA0s9ysXTX87mw17rd8UXDD8Ow/s+Sdq9V
H2nSFv7tk9EimbPVSPHQ/TrsWNdVfIAR8FhgvAYPFxWH4G/2F1GWdVAClwNBGQUm
EQvy5978r2iA5YvBPPawV0i1XrFGbMgACTsyTZHyf+u/6ezJrA3gb2XZoCpCW5KJ
SYYGS5Vv+p/51TCZXE4Mfptrg1qBfELbUJ4Vi4/o6pcsza1g7jEMd5qePJdK6wgO
q5U/BSQaVdue8E7OZHatenUBPaT/zOgQPTXXcA5fCvVDp5stYr84Aq4G/5+C7jio
Yvig7kuRMbC971Y9uteAwuErxH6V9g7xjX7EaEpzs2izvNW1n8e75wcNC00MggGY
B9TmZN0E0p78GpZCEXY7uTaocVIklMoiK7o1lavqqaUwUt1budkrQxlLPnAposDA
3may03Zel6RiDNZUTqGWW06nMWdTLYVCBVJbtUzaMn20Nv6eCLOrr2hwTvi/ZdJO
thEMo7bmJirf/9URl4HfApoIz9Jhvie00WqPjcUssa9C5s6fxyg9o3v/DFtBNb01
fWKr8Ozf/iYEFcDbVAQ/OHWOMdTgsXukx9M+qbD9COqjnwmNys8z5Qy2fcloghUn
c4zr0wa10LpVbFt9nrbSodQRQBrAgUOCWgH76yfjUznwPVmcwzeRVejR/C2uDLen
vJ8BX+PpUPXQIlw6KDAWyh73OOBHnmPlw7P/cYlF8FBdYXVdYst0qj0q/wuZ3j60
UqdcjiYB4rAFtfhINuDmVordTmg35IM5NlWt1XiLT+NFAjvDTpPvoEsqKvfZOcWw
dqbp+BuzFG08wKz65Mtj9ESpkZbaLG55zY9pvNGtmZwvmxDPxxY14IcgRYLoHs1d
wgtgM9157xDB3WL/lELHh0Z7ISD/A5MIEjIQI3F9alnrqe24W2TQio02bsYQR1QA
UoFV5YkEeucDdCQUruvIjhHCUyIVUqC5SupQXyjsc94izEQECQZKketKfr4H/GYC
5jmPEthanP3PRRR9zI+ggYoa2/TN6ZEPKjJ8o3/87s6fw65TwiE21LkOWlNbRw+G
YbLq2ucO87AC2yObR2wvb9CK1T4LnoFD/IBpwg8AnpEX0aGMeVTdVV1tKeLR6cW8
fboYVuOgkYb5s6Eaucc8RSf2uGzKygWqQJEso5sDqFtC/Q7+RJotKQfW6pBIhnax
56G78233LmQd0ULZyxxbXeeuTGL4sNhHO6Lzvyh6czR0bVCDYlU9lPBNuOBDBZIA
wlgWWt/Gy8poINA5qExwbA==
`protect END_PROTECTED
