`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XLxdlXnIl183lSxVkkjit8Edso4OgUs1sGhvAA2jClicGlTMEjiUm5bz9/vovA0w
Bnr/PTNzW1jb+a+ix4fShpuGx8g/Ba7/mJSKZj3yalOTfTNELzWrV4yRDxFmT4rb
isuGe5nRAyDqr2Gqzr3HOlMfS8f6YueDmTKtL8wOSeDP/LbtPbHQbtOlDbXyDfz8
aVFtWeCwGwIytFTyyAQnW2SUKvH50aLSRmkX48sic+sHJxzYyDrfz2APHBiqz1n8
FRfi1lKG7cbSpXrBKRsBPEyMaqiOzsbkWiKQ9UdLsEQbcVdXHVLImjdrzl6PWJsC
6SHJ60D/6IjMJK8Hyv2c1+CtoIh0tOIN65whasAQwxufz+d5/UleRqCR3TiMre7L
U2Z0YC0gKooxaKyqhGQQy/dYZxFBFsgIaMSiT3RVRwHL65rKjrcmGLb9lmOECgBX
ln6eGLhHeLn21gYc4XoZTdcbXElfqqWh4A2dHoKiQOA=
`protect END_PROTECTED
