`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+KWgT4nz3nT4EVrLGb9fwbor/kilwIN0SXC7A7zA5JRXQ6YyjHYyNW7GEvleVZI
UTo6oef+oJNhXg3UFhF6ir9vwFGhxgnfKUSa3UHSs9CfS/IHn+8jb1mYyXDSmLku
bfA7H0KOfAf1PGlfQXRaO+v4XlAqvXFDY5OKxjZXkhMc2VvaXQw+s53iILhjjIF7
qi7SBU88dF1wTpKJ3AFFRJM8DLhILPgHBhjs2WgbaEHqKkfpzJw7xM2ePLkozpE2
mAuvYO1mod4NZx5f5Ecr61VxHqgQBABGChrCnBOsI3gS5nIvJ0mAW+ZZ7HbZaYE0
cfRyS46wJTvzzF2l7DBMNXhNvLnXu8E51EwWoy8DZM7Vq4TaA7rVP7MSlkpUMJeA
wrlrQByvDBfK1CiWDXZbKGHFG7ZvqlOBumWkIwNYpMq+OmyQWzfegOV/rQy8FSMY
1xGz9fJjh+MdkgPoJKWZ6fXdJRLBajq1DQls2YyfKKjxVxNgitUjfbVd9dagH/KY
`protect END_PROTECTED
