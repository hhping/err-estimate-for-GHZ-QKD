`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHY8q1qHCyqstxXNR8FumO6EWznZ+Jt9BR4QcvE8b4xJVHknYOnyusIXx3GVibV0
LIHStJEL4GyZakXbPrejH4N8bVeNgv+VfOLe/KnTO5kG8kDAjayiHUacbKUMaDJR
Gus4L6Cakg89LtUdm8JCRub9zP1tPZyn+ECOI/Kf0lDrXg0uEqLhlaSEB4E/4c0o
Yz+K720Ckfv3NMoIUiXBfEjwvKhQj/RmfQYePl9rjZMOJJtyyQKNPk8pl8wPyQBg
PNMbDq3lb/ZAug2rjIkJ2BBDP9aqOqVtxHORY+DTebDpofh0Nwl0LgKXebbS0clA
QSh7ZgGJ4MiJ4rfRNThfNabhKBC2iEVV0P77URyGPqBNikrx7Rp2eP6W/HwjvyCa
9kFiYcqS9NDRyzbZA1EkYxQih1Z/GNzr7GCzvLpnUuDwyVJVq19S31wvo/OrvrMd
9zx1hImoB+GCBjhMFpAZYq6eceZe9MUlOjYIquIYBvw09Qxbm09K/WvCdPNaXvy7
Ak7uYA88ak35dxkEN7T57nIiVQSo3vlEImQlUUCPGAjOI+PivYwJG6UflCYWuR33
Pbr2o4t6NAqJNxH3WczSNPRWNJkfVvnWljMRqhq0+TCTwtdJoEL611Ni7DyCSRHK
j01vbgGfkffI1jtTGKiMPsJL6hADJizKtlHzoV5Z2VMueDBzlGe4XId5oLQINvwT
KFxOowwNravjsoaToI3ssHyJ9qrTMN2oSoi+MezvIw2FUsBNmR6jMVlWg5YjW0Uw
XaRS0eK1tfm6T6nWBMJSw4jT6JieJjhD2TRiPfP7g8Jmy473AEszIvXbz4CFwt9J
DugMCYCOexqwdQdyOP//evfly1m5AmLpJbFRlAza1V1oLg5+hxagN9BGkzG9xYyD
BCGK9RSuSko8T+S47b7PfvnHFu1vvJDTj1V9iDQMoCjmt0Ax+AQBV/N8CuidJuQL
ZhZNY9dxm5nT2Uxej1MtsFQqXIH7lCoZFW+NptLuOV/RtyFikmhfEB0lgajvR5Dq
hhzsr+9goF9Kst1nvDx/s1ojvXe3EoLQIKVayyWFgqUfMqKjxuNKQDpGbXxRytY6
Y0m/jKv3UsfwctdGJPJrmWDNkxoFidHy7T68/24YovhVDDntaSoflLPoDVTR9048
e2yEyuzKHYSelhnVy9iWb9225W9pD0XVyDaXB+++X2yrTtHVBXq4x3i4fFdCSDLh
93BKQSbS8yKg3E9sayh35jPeBF19vb9fF9r2sYET/q55aHIGZ9wGIJ7H0T6NBzAv
TkS2xHZkwVbhHZn08qN+LG3009MlF6ABuTHuWl1FGoqI6umqaaBpyHRhDPr+Q3+f
juOKY+rmhe+ripNKyHaXJ91N0WUNl9H30b6thharYbqKSfq1QQjiekh5xYbv6hJl
rg6l7MdyYLQuAt/wBpnUyqS5ye4op5E8wATb5dFep//jQfvV4Wwhn7WwCNhLKYPs
gcejtVm+kvSWdNOFxKBokag3hUc6VanB5AgFAoS8Uf+XtYa9qBYTVOh175eh+5nP
do7LZuvmjNwOqWlT1b/CjJklPLacrfDoollQGaMKcE0=
`protect END_PROTECTED
