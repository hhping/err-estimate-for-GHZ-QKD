`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgnuQSyQENxoqy2lc5sGU7xBIiaZorXJxEIBBabRsYFT81ZhDmXiJ0wtjcuGTWNz
JzpTf4W7O/lAtpfDM38ktoWMS+mzH0DLlb0LXU1OeXJVewA8QpVXKTjat16j8s6V
6EKWqADWTvla7dDgquAYNeCBuCoeXjufP+cyrq8PasgVNb9XBrzWaiPRy4yJ2Deo
8S4+9W0eFAx90652VPb9ORW6HlGg0cTN9jkGKPq7tHiiXnV17nBFGc/gTld7WbGn
2c82b76QtLC8fejGYuEB99ZZ2a7Zw9PsARf0bswUhX6obk7ZWrsgj6FIUG2YHncZ
sA2aWrgx/HTt7BKFU85qPzMXzosEh07vifN1n4Lf3n9iE7gOAovyZJV9uBvqk6zI
9/KtekZW2uVlP+z3NDFGBieW4nLUPweO11pHNUlCDL0nBQPGrMmnwgdBIRBaZLL8
vWcX6NXafM8PMHXvz4DLMXjOklPWBJ5mLyiV9Vm8Gq9VTL/tfh2ws7LFzoBOkdV3
y4DtltjWOYvznoFhGeb4POztH1fk6rOnoTEHuPQMBEWpitebieB7e+Jkj8fYNgL0
aOPem6EYZUvvccRzumV7l0FvX6p2bwQzX/SocsS6OBFj/NeJ5uzIEfwRmqJCRpLG
iZstCU6v+FfS0vz1yy37tgZi+xVfB8rQMwpazmDEYjSjiwCzLyPbBExHiCte2xv+
nSX5H6zJK+PfoS5NA+CsNbYIXypWVqBAYLNOw54UP5jzyyeqMcZV3gfxOc3KryPE
yjcdoylaEJoSv5GZGgsA1SsKOMDTszHGKIZGPZJrpo8Wp4ZsXxxH35Sy8i3lXcjN
UcIROIuwxHTIbZZu1Wnt6JXLl71/AUkS91TEUpKHeGfUPx00p1O1XfT7FeagtkrM
ZZjNgg72seBXKL9CMKw7jKrrEIhqPR7V1mTzu3ohMrqy12Kmg3s5gxRtjtPqkmZ6
2MHCKXPMm2KOG4ZjROWNfiVr0ZSJF/lEBeaZub5xgyHiu28g+XUtMoty3zgO32Pa
rojMEeYuL2TQHVARaGZxRr/22kiNXcjkmLp+UO+KzmR/FnRUYcfYHEoWSAZQSb5B
JEK7cqXO1mQsaxFGWmf6UcjDwCjcZx+U7yaNSPZ6ZbZigQ6RqZoFCZf9p/qaKpii
2RKrBX00WF0esL2V2ZfD5JFYmqdmXaGEBqNK9q8+E1btXfSln20rWXadIedFsx82
AEZmop60yxSkm+kLF0MR+yF3zgTZITZ6zHCGtxUX+Lc=
`protect END_PROTECTED
