`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+Sfp6irAiTC3MF0DhNW5kW04n8G0RqyakotL5j2bMlIUct44Xaj4nHMylozm4jn
RI2h8MPq8iqmsa4CIZG+LXElazjAD5MQEGYJFlmzN9RGUQapatkACE7OaRxaWm9J
UGWvW2tllpJWTMqbft93M9CLGu0vZuk3/NA5iXewbtvSWY4dY8i8XmML5UaY0ha6
kXuQ1wApvdBgEUftH3Kh/rVCExcHIgz84dH0F1f2+y+lBYCEozMQsoTzdxyDOFbO
WKDe7Omxz3wVZ5I515ldcrNemR12jWMOl5c621gDG5Tty9PrJT8PZnFpPRv3OgK1
6EA5vpEshbvK3m5PWse/xN3fX/6y8t+FlhXTrZ4Ynm2jtloySzQNfNem0FjrMAsI
ZGy6FGI/ZkOz9o4Y/b1gJN3Tlx2cBrcRZtu5hjlQ5Ko86kb2ZDm/igFx51DiBMd6
R9+CYxxCNzzZlpErgOgK5r5PWujDGm6yr8PWnYeFObPaL+N8Rb1Z1HeefPuaUiq1
MhCc6rF1uxUUJSYMLZ4zmQMYB8IDIHIpP2dYJkyN5ZymzQB6pseljt/rJAQNnOU7
D6zRjmWUdZufBys53TVogrQSxLU6lvkGfPZx1eczO79Er5jD3E0w+2mL0pm/m/d/
nMX54XZbh9NrJDqFxtRIoA+epnEj9g97Cv7s5x+4jh2FnTjKdVyaP8BxJ30jxr6A
x/dbeDLCPGyp79767Tw8Jn4a1klLPXF1ZRuX95JtJW5EdD407b+LnQlULyCwVBWF
RiAAP8skyTLOv9YuCoT1Hre1NOD8Rd16InY3QERfvYddlZCeGab7tUVbHXzQJ53I
ChNWBk5eQC5XZih7SRNRBVD9oC/xyoQcFzoAH40841tkpjBuT1KMIDJbknzlxY7N
pOGxl32/DHvJucGgG0wWn31db5hCAc8zuSwkEO/34rfkqIZNYMPp3Ih7UeByfI7Q
j4LmGfPSEMbym0Nj1YgnhwKoQ7St49VEZftbmZpwmHgPbndS8KekGTvHlOU7EGll
YCuYafkhRCHnXoXz36lZrln7YEc9LjsllxXK6cSUuH7JZyEwMY2Sv2EAfkhpcb04
WTVDIX0RwvBPV+r+DC4IzrgrJUUFPsReF2oNMCaluhomTlRtNZHUpBSZDDV069sM
7wtfPoy8phMCGlO/VsZ4/sNgY7HOGjiA7C8BqNVZfqQ4ZtVzUalGMODmRzSmuht8
ublAwRSY9TNinEnpYr0sAHxaEB7ty8ITeK/WkXE01RsDqMNhvcfUBEDV55omB60M
Z3wD6iXap89pWHoUm2CvFIis7j1yIO/uezSuTkDI42j9QISl1jL/H9TsKLE7PHh8
I9nH1z40def4mYBMXMvU52tnoRR0rY8KVWHsUeAoGDkMg0bkw2VwFERa6q1oXvng
pTHfYN0tcjbxHEgK6s7+lWG3WlQjKaJEWhR0VwFVBdfOw5FeZT8n7wX4mjfxgj0F
/Vx7USJ3AFpUMxkOXEJfRkd1buADaGY8ZPRagVERxXxkFjXv9U8Inwx83k5kKpw5
jF3qcc9iyQu7jIsZybqa/nRoVpiiz78nBp3wMz3yx322y/Cv9i6gKztn4zigRZCg
Z5ELmohOK9Zm8Ia1pjjMXslL7JH/LzhVXhxFmy0+sx/BW9UIOXmPI22beBX4+j8d
uo8Y7H7R+U+Di9GvQvkdlQzpNX00nFukTvFq6fEivly9aOy/oycBzrVOa2PeXC3s
l3EAZXPfBTBvAmr7wQYuiLR5Y5p9X4t3yxNlkCLQRsD6slEymUv0iwHf9xbw1Vo6
if+VCqiMH1bU47qyHYWXqwn8/JGE44EzqsMGyF4VMzo9y/2N43bi+dS079Eh073P
lB0MSyP9kzLI3yxFv5mZny59AXl/ubul6CCTJt1RTtzNv3HRJS/5dB8fHkqXn2oM
D4X78+XfxLHCBIGzNPFWT/zLYhF1ZsI54U57ZlRSxzr2y8AXZG9oC5yyqr31Lt0f
VaJ+CayczXgzi/bDLqg39UBk6NRSKOB++iChQDm9e2MIWWAV8JSi9AqN0V5e2riZ
JKHVQqymabTGN8WdchnCfqDqzlhDoqHDBdOfLqD/zi8Amu//BMZPT5axeE1lnDop
GwQ/l1iIbDdjLauDiziy96EMLvY1bQ+mU8k7gRr98pPZ+/UQBAyGqpkI+BQYBBvV
Ijm2Y2P20CL3etNf9cLpWjiUhYUIJdiAy2d5N/SZBZAZpI7zPWHyUTxwmJKj1P3/
UmNhtoxF9C+/nJl/bGEmYpHlyFZagIIG0oLm7oW0jhX6lGtY010E3BtMdkbtZCtx
WvvzXuxMWoSPpw0CRwVkRAANwloI2/Ygh5USQf0IJZ+aq8AYyBMoOSuZVPYLiT7d
KvxdzeLoT8IJwmQJkmnp0YTOCvLR2fDZfIJeEPCY1QXLTuB6wByWAbJ3ZZ64C3QR
Zi2ROe8QSx4g5ag1Du/FC/XxkLjs/Aj2hoW2WE/beBEv1mbSqtSowSQ/rUkSE+Td
9frCkcPPAABE1osX1WOxgoOCLnxq8i8gSJ4C8muxC2JR8XXM6IPcD5/NpCTinQ6B
t2ESl7pbarb1m5f3++BB/r8KZlzhXw0LhY7QPFEUa/6Y8OLld85XeRQ8o6DK5aYM
eY1L3c8puEQiA8vMCRKjHY2Fzlg4OeqnKlrV6G/UaM2FUuV0FWqxsl7W4aXaTTpA
Dtwjyq3SP02P5xR4E2ks5vqxluL27WoDLqqIyWuZRIQxC7VrG/nchSeQQHBfm3B/
KpJ0Nf08OqtG9hjRMFMbK+bVaTYFWfNa7yzqSR2BAvN4S2mtf45iW8DoN/KlT1Ar
jK6wC8Ciw+oXMubSsBKvKDhxgBN1CPndolqQlBAOcjC6b7H6/jfrgozIemDIBrNH
bCFiJ0Tgx2I7w5E4jZxVBexqa35jC2zVC0cASJosIMNCt75xqq+siLIcr+VsJ6gS
ejOKjvXkAzM1fobTJ4ZelTUQFRNf3e3mfh1IMAm/7vGLGhoQT6QY4IHqWWSWUVtT
3UkhfPPa21tIQDEftPTOQs6S/H9j1Pw/0rrMZVsszWAB62xQOJFjSSeJ4tzJpjQr
TQu9La08PyDZkQCLy1sAYB6ZwL04W87w4vcWpEittXaodqGRRNBFbifn9GfmeMSn
9Oba2wcMVYwjuU8ecpVIRfScmUTQkQx4Vf+fz8pFesCXIcMDY1pUZ2iZqBajL3f2
8WB7rKnfAjsYcw5rJp5xuYWLGOSkSzBIKX8m1s3eoSau6tf1OSKXshPWlBAnVMQa
Ppq5oSMZ3Q4MV2QZIaB9OdOtKz4CTco+u+0cURGJ/iuO8MGZn771PAPwVXNfvPKQ
C6QCP2U0YFPRsbDvDlqZsh6mKD7P5ONrt+/ueopNlUOTYVbTQaHIYPvYzEo3z/GN
8VBBnJFatkMHmllZRPCuEmAc3pXrYg29zfxRzmAflQ8swQ2U8pzgzDG52TL+M2D1
WQ6gCXhFeE/g/m2B6gLg7TDYkjBT6oUb3MjfCoxCr+a5s0ad9HhRiNWRN7dF1MyP
EK1HjmeR/qas2F3rshWGOZAM2tylJJ2tY7lyW21XLHzNvVAoiqxenkx+hQAwUPMc
X8jvpcbiyjH6UvWjRLcobN0UxXqABpoQyBQfusJKsUTVE1eqq46/e/H2TnZRsnID
8xTV15BJq2fBkkxoZlLTmQvwL6Ammh1Yib7S5mIG4l9o75FgBq4quahMbKuvO53J
CG0/un39E33RX5YObLirhRoj8ZUzPXrk6BdE1iu5gLDYQyteIJuBYDXv8wyjSuFR
RDOd675vCk+7JjBMiixFLfKZoyMpGW56wqFyeXY7owefDbXUvTlzSogxY0snsMlc
VXCoP7iQgBX+lmM24l/5o2zawTeKJ1XWmakZ9weoRte0eOF1TyDhTtJbHGuzy2oa
7Non74hBBkwJLKLMlsUy9DXvvb0MdMATW9tpFKyCs+dOf1FjHQrb1KJn2RyLY/Hj
zMDwVJgvx+x/+D3aJfvuHGCemZNjRAeI2YQY63FdCgqpT9483tDlDY/EvDrCrdSx
rAe5b6UABS/WimgC6/K0cgiuEA4LYCEtk8PMFfX37ADVZBp+5Px0AdzY7/XhreOn
oqz4zB/+BT73bM6Ltjrj4d2UeFAVGZRIVqHV/oF1lFpcSonj8SM/z/SNFRlqbL+8
h7bqSLNp6u18+I/bRMobGuCSL0w42nJK96Rmfj4ZNudymK/RjuV4m6vNB2u2Jbx6
cq/b5tSfnzOkpbTeAfzMSMNkpKW2+u3L8QhvC1o9bN8lXP80URf/YQNWF7XvkX+9
jtzLZHzC9KFwwi71+bojapsk6cokwM09WprYMd/MtM9ebTq2EfeLMPwOE8ZT4uJi
hkgH5zC5e9SVf/NYEEci+iqgDSwD/f9/8Wd8v9JgRJGwpzbsz4yRzOCHd5GFc2rX
/i6o2NEguLVc0ILWMlYcc5SM7hMD59lms4MHBWZdwPJZrA4tlR1ca1pcR3pl35BM
LWiuF9PJ1yUsTsEWTj1Ol0fe/HdOEgtondItsk4CIpYdAKNKDJxNTKbZGTeRJ2kK
eTkKMIUw9Kfi5aMDTKyRpaK+WZlZjLs3t3B8G3ny8KGc0gq9TV1mNVEvQbW+wAGN
2OysmVvC5BB1lhQWpCS4zSfQCKIoXzYN6o6X7EW521GCsXrSvNd0e3b9Vl2HTtGB
dvFEeO5eEfACfGEo/EqO9Z+JJ4Ay3vj2O+Bl/q1Ph0yrV3cDDXIYjLj5gxsl577m
ScBlEUdCaKTA+uDAKyx6czGZ5AaTWzuBFIJ8Kte2YqZdVG7ObCGKlc1sUkGQMYjb
XeBAcJGe/d/wubsePZ4QnKxH9aWgNeVcpq2FQ7qbRYrojyEoxwDk4dYU1gpmVi7J
SCsihk4gswwx5T25Bu7jFsf/GKiyHOJeQyrENX3cmYTegfnl8eEjO/eUbF41YZe1
sIrDHQFSK76gql+g3HB5xUUcJxCvkKrAhSt9ncpBisP9iQ0AiSqgc80S0x7U05dO
PstKkXKK8x4D6i8AwQp7eT5ZqzufhW53cQ36FyrsDxDaohI6vLNt8oKgQsG/Ho7k
4ilBV+pcE95NGdKLFU2zcfPCFQNAdZI67u+/+SG3OfNRYTnCRmeoL0B4mDWsaToY
9cnAGXVvnTUK2iEvMm8JYlRjSP5z0oQ90+1dr4o+1xdG03sXJ3s+m2f68ZVqxmAl
BGqF9FmmEwSYZPbinhoqfao/AH+bVUYPOwGn7jUCXMmNlxPZjgNT+GhmWM6s/qS7
LtYjps8gQ6OHsyehPVaVxg6eTbybjncoQre+XSWh1vxgKcI4oaQkH30KpZNYDf5K
KwptQpGH9987uZNh7eMvp/wqN21B7VpHuPhSDZuBlvAYzmQa925y+CrBkxXfcMZY
IgIgmatrxnwBJvNCfGdkJQjQAzOvSMYrq9epKxvEwb8my3UTqTBHuHj/UjAozW3f
2t0dHgRwu8FkdoxR0+kvBtGWNGojEsoL/aOV/fu8a1prQ5Np/5E3CO55St0gj2Cq
Ic3h+ZKObvb/6NwNrgrTYObfo8PXopRABhyFvJfoSEWExz9k7eeglZngEYKiuI5Q
0hBNGHERsK9PpGyiqmIdKquH5SdFXLJTpuN8/IwnZCRAr2RmhcHNhBVkf+vBrhGg
LL1OKSsS/Xw35v/cBjKsyZlaPgGA8lOUQH7ozDcULazfKcIse9oWS3q/HKE8JJtC
rmtqAQ2TLPV7u4Zw6XlvjLUD7Fu0RzD5iPl6kNxd3f2OB8gL3EnimyrSQZ6KY9IL
oWMlEb7htq75opi6o14XJ83Qrk+G6ar6hTXG/UiCQgNp6lABTRFp58f0l66YGsmP
6zeN66V/YTTaUpRarp6yGhjY1gCDI0CUhcrx3mLH4lmoSanrGW/c4u6RL7xrttVk
3kKxubb7JUmchUB2pndRN1tTlQbeBrJCrplnoh59nnie9IjHoj/LCslVTUi6rusy
hGD/ItHjOW08EW6eBbNNw+zDLq0eM/Bc4/ieqXvgfSTLkcdlWxM7n7g9w6z/R9CC
4DhdlFFpFTEmkq2IwXICbuhx/te8H35GQO3O7cmT3KFJHjyJhkDaQtAqw2yBNGeG
nryvOltI10iji2wH7TO3QoVHbU2NGYydDLuVBDp8voZIRB+0sUp4Z7cBl7kNjdyV
9obbOY6sm2V2GaOnayVUKvG3vvCUuYdf8sTc1DlmZdySCH0pY+MsdqcY7CPbukfL
5cRDfzEynm15Qd85+1BubAaUKYB57zW+0YiNrXOs1Tbgfnpr0pZfUzuFzbp/jUs6
3lW7SwcRb06qlas3J/ss8Tcey8zDNdn6ricil2F2ucQuIRq7IPDNxUutz74g/rfk
rlqwggKRUVFYrVdO3tTK4LaojWck5IqwMD99kpRq5k4vGdb2+vi7VPgIWMf0ZCZl
ZYu7SfcdllBu7ZghtRBdD8lNvp83uL3ukscrj//ZnDacofx8Yq+kMN8KJgZOC7Dt
o13su9eJ3sDXcxYgETSGwLz3qT3E+wiSjfDtlhmxGyQEJSvGemPMuwL5vmf5BHA5
odblU0SzA0pcUnz6WTWW3e6Iy8J5kPTBVSzvflnlWdU4BbZS6Jj69faECJuaBb+s
3f9Jo+j3IVh3fgmCIOUuZts8ODFrpstobm2rsUpfgCIt/BIaQKtQp0fs9qwVq+mv
+X//OsM7m5d7bPux5xDktIndJ3UrTwmyv/ST09q8qRkAXI8yg/Sjc7SI2T/EhYZe
OMChkh1fYttM3zI/WNn/oc5778BIyn70cvdR99Pjeq5eA8THQciilPBCgKPnGmVx
eHhoBRQCQcwnPlGM0cDSHWLtyIaKHE8x2wMJd5fIEL4MMeFW+LQMT3u7pKrIPMcx
/eL+C9jUq1w2kTlGD74wocFWB7tQCWNERk5srCprH83bL7TK+++h+qOnmjkC9oPd
JFwFkY+HnguYlbM+XUJa82wrc/ybtTwErzLvbEkx9NykxX6UWO3iWUZKSM3gAQnK
T5Zj552t2Ll8O1fprODHgnrepYigX8WDRVHmwV9fit9M8BU/+gcujTY564Rz3lQf
xLPyJ46Q2SZBVuWRJuD+DxVq+Ukv3Rqw6qktRnQt+0Tb/Nibf/L+yTys1bLg5kAh
Y4iMscipOrxslaZvJ0dV1+YmlL4QvdPNPoFiyJxZrQjP0c8VMhqtKbZvQW12KVpe
Aa1cAbxnMXsZEgGOZco08TY+Jv7ISUoHhj6wQSqQDOm9ST0kckwdOaK2VNhtv5Kl
bOuZVY6pQd0paEIRpsO+AOQeUvczkkOxmTqArlMAL893sGeoh9dKvAFPbfut222n
4HqlhYVxlnPoFxljZ4lnyEpnnh0GUf7f4/fZehV2FdTcoKG2IxDzOhgVBJpmFdL6
TsAQpUQlVW8pQ0tMgfj0GeSrYZWumK7VH+PK+KLoa5U3UAA1w+b6xb58eC1lazgC
H6FwkuEerXZdwJHI13pWk3eNfbZcowsVqOrjd0VpzHO+ap7CQR/TQW9gKWQCmfnE
yVlV5ZjPTGcLmrEFbL1VM5ZkzwVpLbt3UWJu+lg0Zb/f+8eaNHd7I9bsogRHgsZe
e9jSzPIaPQggJK4hyqc5R6f0ZSlz/a3iHU2KdM255uoD3kujnWjAdxlBx46yXs8G
INRCdX1uWNhCkUmINC2EoJce5npNVeqjjmBB9Rb3IkX/dj33dCjJADsPwJ3LAs28
i47tqffsjxZGAJjY3kmGgHjOC+69nfh8vNa6TP/wCnBB7i+Vr6wqQhAlnQ+1+l4X
U6xiAmnCoxnZuvRtS4LEV3fPPtYKYIfrVT1yoSOGfU1uxXIUZmbzVf0TU8By3kuG
YNKzW+5W4uqcVI1Gf70ePFZW+TuJnlqtgX7EGElAbRQEgsWKK+J6lBJpfc/h6V9U
/AgIBydme9bTsS+zYHGPWgIerlzDuysRWyvRCnaSIoA3QkA71196LtTFegXITAaD
GjvzpJIcMBtAfjvfCmJnYUkx9i2Ra4NV2dh+QKm9/CNo6nFKZljeGxlFzMMblufN
HTEQUlqiXp07KqAyFIpw8GYWTtpfwmSs8qzMZFADLe0GMZxyCc9B8pUceyOSEgTE
343L89MPlmgL8LUSEwaZTGWBOfWbw+YiPX7ppQ9imeYJTVC30rbPZydeo16jEQeP
5qBVU/I0ARcZtbmTtHNozrgyQOAOrMTtJzLIONMiOSRK1xEJLb+A+SihYHXJbyCL
uMsLaUgEsENsHvmAHNsbSMSksf8nm/TbTu9qEkFeRXm7UOpiknasoWzjgTJtTKIa
cMEkig8hswxg7n7k7pKkqm6PtQBJyQ6+8qyNGp+6Gd5t3krRPCDRfzTXdmaqqoQK
7QYfvu4U391goxevxZcCOGUhtE50sZ/AGuOoVwAyYsR3DsclvE4U6Q6Z4JuVgGTB
5VtEbt0O1gHMObpxIBwhBma0KkAp+DcCF/wOPq8QSxuLpS70teYnNYQ9cqffbdWr
74QwPgHOObL9c33Sz/cSNXZ9nwkln2XEiKkQBsZvuCVPMU72k+4xo2IwFQPkMiZr
a9ZtNlrmHmpRWslJhf7zVlKWZukTbtULiJ6Zm82daqBmvyXujJmGBCiZSDEVe7oG
GKbp4CKOLejv7bkXSPmpjd0KBedlhNAYgzJipGrXvsC01xY7ST7KOyn+oeaTylls
7iq0vkHMm0lLyupE0T6djYtsxWx3eijdwPLWX3lWHxBOhLl0inV4noP98/LVZOgf
yuzGq7kYKiM30aKCSHsUK6pJAYsWTx5ne70Xpq4wQdYxQyz1b58KbYb4XI26Sx50
ymkS7wczpFc9qXz5Dxm0XyVPvupuqRhpqpoRVc1p+Kk0bWGLc1ItFCtbRFYqEfr9
E2uMXpZGvt4qzJRkNS1pKoe5+RCZjCUtNpe4X4ceUNol7NtlVmxXerrYf+hpV4zP
oQXsSNAD1y+B8M9eYC385FLa23hb2feJrma4suf54yAQkcTVbkXy6sFl/0Nw/eAO
cAINqT1yGHILhKhLPBO79gd1eUHsz6crir9+p/czResH7qEV8WF089Dt8+r7gmcn
84CF+VUNCZirb94ZXrZTEYReS/4Y0YXyycX4u/E9Cw80Ynu6X6m1DMQ1AJC0pzTG
nFhe6xdPGtmd5KR3zLI1zBBxyAQjNnLvVDxylxrpfKAuEghT3d0PmMO4Of/I5QKF
SJlkMAMN/YzWegnLkfeRxZ5SXwyd2BNrbtso9rTJAZUBrEL2JHJJGZ8uplYs/ICK
ubkfQGzHEQbq1TXFx7yZlvEG1gVCiqtSFejScGOai09xZus+rPTf0flP0wwOslIF
iRTQ22zw0jeUihEsklzh/eyFS2noQDnn6uTWbUlbxutxF/BCe5vrPxDKklhEliXD
eN1v6FxZjxe9S+erKOiYyXjFx88zRJo4FS9xR/3t1ZtYwrpM87C4DPYEprb5ADcO
CfiP1JvZTuy/60otAYK8AYz+H1WBXTscaaf3mJ+rszBDDuL3n/R4tYeNrdRxm95k
dZXBltpkbTUphvFfqgJRnelJYBqNeJgJ95XnIs1QlB+/ic5R9AUMbAffmtNGAKPJ
OBhXO4Tu5EwDl8dBnnhfYjtjQF/cPVNkql8KcOXfN0N2bdgkGLzBY6C19YzpnRKW
gBeqgXejdD1uB+b3nJrmwhkncLyo1arQ8+46FH4SEDg4nUGuT6kHqZYsk5Iv/40B
DJonEWmh/CfIpNMtob2RL/DCNuKxaCLAt2mOAu3j1l+cguvxTkiX0wl4lmsRIsee
wQmIMnOQVtgEL/Yt/qYGjFVrPdwHw7jlaI9x9qCskTPYjXoiF6qK9az75ZLtSwWa
uAHAt2mIUxZgOJdBtJ5p7+GTuPf/dvLp6QD665Hxy4RtHgXciVvYDW/UbkiFm7KZ
vSMhU6i+B036Uw+yqARVWrf6i+Sf+/DXWjfFCTsBpHOrgodDF0hbbbvuOKLnp/S8
5H3fILLZtIWl746Iqy7QyCJ0FMz6qjUlvq5cvyH/So0anu/muQ1LeuF3jpjEcnht
ek9J297Fq26IaJ7QO2vVQakBl2DeH59mTaZ0G94tcVTbvQ3eomW4yq/ZXik2p+Um
IqYiLVwVjQIzT2zrV9b4+rvdJeRF/4ES9XEATBQW9C8KVCBS84UL1mu0ojS1qhP1
wQpS0Rka9g3X8D+EiBjIDCdZ/zeYwNBIT0CHaeSJAnqzebzN3LEMr41R5LsFVo4u
yyIa8LHYD8ymrzIYpETpHWUgulZ89tEqROw5sUw45l+pcbD2omCWlrIXlKj/5Q6v
asUV+t77t19OigBIN3iX94MA/W7Q2oVGG3ECjUlYDzwBrLRDkA8mDFjx6Mr8Hjp+
eGt7yvyKl+syZJ3BWHXV+5eyDqFot6wpKdapUAl9Pvww/s8PXq2zTLYpIC0Ujj9T
mQ7ymiOWUBatg8Il8S2aF+KSQyiFH17Ih8W/R2Y24Llv4soChny2CC2TO2S0xUR0
/ziKEU20Vd1yGKfAqKjPwbbNDDHcIU6FY76Lk2a3uBV/IrsSTv6JgOvz71MEsaDq
BQJ0WP5hT/cXnQvxD9yPKV+ldOnO4tZs8snT8Y9FKNqGJ+hSsoNEalqWbsvgYLqw
JKIXG3pQozsTn8Lao2AepKGmPNqyVVjRY/LXZ8Qt2cr38nPxd885lwJWC1MzyZbX
ZTHTUDJBqK0qQaaxB2kSBkScsOxyF1/m9oIHeA1F1NoIED8v8afEHsI/hg9iIAYd
OlTEczMQPyuskk7SIsmgykegr7DUBrvna9kRF5pkPuXuiKHAY3f2XdhUe3jzheAO
kG5tIfP2jkeqh9laRmOIurq2ymVmvK0Te1Oe9o/VKfvckU7xC635LRl/omUnhWrt
P4U57LU5ErEwkgydt5Kza+ikV0VDLPBV1iLzbrIkAUwATJhD3wdrZVfbnofqnmB7
T8JMIrdu/zFOvSzVV+ar7QOcQgJ2fPaQh3TFBLKYm3CaNQi7MMB40Mv5ImUVql99
ZADAbcqvUgjFLI+BO78dzIo4kGCD3Stj64GyDZ8naDhrtIIrYJr9Csrz3uhQH5mu
gRNULoATG1qozi3YjrF48REEAzAku723bhWwVzE5DywXlv0AUNIwBvnDS26gJGc/
mqoiCAX6W+b1gM4upNWds9mpYM38+BbekJSluhlSYf8zmG6A1wtps4zyCerZt8No
jCOfHOUoIf16y8J+fZCdWKSTlY8RM1XdMJkpXezhgU/qtxQ6pRN7kqx07uxGt1R/
y8HXL5QmpT1KUFesCj2hUhQQJZixGgQKynstrvCLjTjth3pGfTQgAhPhBtmYDGpl
lgemm4FCV4Y3LfBFC9aUbPhegZ8dC4i1iaE3KHBqbBS7K2uUr1p9QFFfRU23/DfZ
jd/n5UylTcYtlf1JZQkOiyl8KgkyMZ1+MM/k5Irkddm67vx/Qpty+JE6J9PpqgUh
wy6qk5G5aySNYymjIOLGqd8ef9zFONe+e1iNAaIDgk0yReB0Sd01EwFkltygoFE3
hK1c5ofTVProm925iGM1ocOnanh6cAiYzrMWA8Zz0vRrWO4PZA5g0YVs91GEovDD
SGmBn99xt6lnYvk2iFd721jbE13+Skb/OZ1df9WUHdZl0XYLGGrpsT2HkJ1pTo+f
oNOBSIVttMWs/zrHimIpqWojD8z2kJg+SksahqDE56xaXPtAwIR1tXCTPdJ/4y/b
ecP3mlr/7MPmhbQtxMXX7Wo8nW6z3jACsT4NzlUyuOHRcixVaXa4KrThOBi7ceVv
o3SFoqEtWdrbAoYwwXcObeKxSXvlMnILNTlM1LXwi6gfRVYYl0lYqiy2IhujBUTR
lD4W+0QauXvRgSqhp4baAPznkQRN4Je01VS4g6rTwfVbo4wZ8sAO5Rooo6u3zf+B
ZUKbrfR+6i0W7VjXu/3S43JNkew8yb9P2NFHcwwawQ19qJS0HtgMsCnbmjfR2d5l
CRpnIuq5afV3js91k9LTRZgBKykKpQWQ4ule1oe4r2tpjDStxXIRe3PTT4ocW862
dz3qKexH6t1Ms3Cfpix2JrJox1tgF/q1tPPY/GcfuJujMmkCzM23JjFo9GkBc3PH
kUWt6T5MLM4zTlwpJq0/oJMYpNzcg1hnw7d6n1ljdNjc43zKO+IoeBiP+8ftajl9
Juwd0n6vY1Z/uL9HnEfJJ0cOhDvo/RVtRs4zLPZOBbnoHUiSeo7jDmeUd4KWewse
lEpolI+SJb07gbmFSj221/DQRCq00+Lc++0NMyKprATmpB83AfnNI6t6/NAb7LPC
Px8b66I/yQalD5n0B81sr1Pzd50FZAdly60OaYBSUQ3h2uYiVWuHCVQI9tXTYw//
etT686LGCuWrJh1K9btDv/j0FcxuUi3kn6lQ1Api97F8W8pCl5dWfncqkCggWwEW
ZzEe+calzu4+b3H+2pS2A9bam6SiHzMXq2o2sr74TXEC9z+ulVtNXlvzgoqvBNMa
SL3qrt5mB3A8Qq+MwvenfJmIr+NL1ww1JiIYVYylSjZu0BHfGQTFWdkuF0P8QZR8
Hpj0hJnBWnTdpyTfXuls+m4pty6FIWPU70aMC9MYm3lnGGXm69U7OuOI9K2Z4FVd
DEfRGmk13C64E8qPTLXcQb7KiDOIR8IcXXWByYtqtDFMDVYFwfqodbjvvKFc6Vsi
5yKor0F3sQzJRXyW79BC7jueNRwAxouLo78VllYMTc/2ectE2iWHCyzaFMtyd8yP
KzwvyBdPyrOMoDdvgAFt692RisWo6uCYKFpRTlsBijn+a+7ufUWmOoHIhkjshAGj
b23MnDtL1j5L51F6z6xTJzUVk1M129r32AdHoX2Ahr3KLXSrUkmMSBJMHIelJyFH
k6ssWHOlVT5+TevsUJu4p5F8LkuZE1Idl5diKWvEeK2n7cW+rm4vVA0O5DyW1ShH
p5W/9GccGFnVjxkMONKGy8sKhurfy8cQXI3mAdSKwAcuTnUsmqNNDBH4ARRoWVaC
y+PolN7NtpIo+ZGBjHtBO+kybP7L8bltYc2ea4ogXdvBmOkPWvukBHCaLIOWa3yA
drP15UlxYZhriavbDP0p9B2kuxsVtD01tw+tuEGJL04Uv+PVo902bMrYaWwfoq+5
pr7Rz0vrqzLaTJyEuCve2BKw0eQSUkNClt5UiXWmIDGZQ1QjqInKfQzYYqL4EFfd
JoSQNAgnCs+q6XvoZ4OcYL7ZhJeOjRQOvNa6t/AMCq/BYgmQIBrRpXQ7Fpno4FFS
BrO0NNiF4cwokOsKt/r32ZvPD8NC06Z0I8diHKGkIc2I6zSQvjBSLVtwS0kaHs2W
wDQWy7ulQ14DZW1IEwDg2MmDXQqgwxaASvJEOlCIbWN47FfyJ9gSxejmgAiz0IIG
awqrIQTeclcI2MVH0+uk2lflP/JvPHqGpPziV+hrfdj7Ev6mElk0hyhvui3qaCFV
rAGBiirZL04Bg0w5+vAIiL4tVUMdmOAXRHUIAXz9WENm6TSsnI89URIGhxKTlba8
jKw3WqNSj4GwvrmVXESRkWqQJWy9SprhzWZ7d5Pu2dSMtcsLk3pPsC0DqGH7Whwc
Z1HAHbSIrfypLSbtlDRH/R+rqyYKkCax7DP0M3L5EObnfdjDu0xfu7Cx1jKiGr9q
yOTijfnSQG9KKjsPIAsqETRFc7F6DMgnZq90dTmchLhdBcAERetP7h1EfxsFV7ao
QvH1PdbUW/8CF206wWvTqLr3VegguATxJ6cxOlNEslrc3Iotn9solm4GR64c6t5x
CJPuzsSdrg/wvBaRBMY0pQHWuDBcM1Ah4sQgK45gEMwg0Y94fDIanfWjZhAVlcz1
tjHdU4UmAhZDwKxF9X8LftEXwNZpuCwU5ncYiGRyyjtXXpa2hnuK8Sg240zb5vCS
TDRiV4D71gKOBAuOux05FNExZVCE8x13l7usi5dHURfBPnD9sQycM3o6qLkweuHj
G+jVBY440p0YZJqikngQdi91R4zq4sb6XPgpzQV879dly+N5MPX2vrDUJJwWkswo
yCTnXAgn7wZLKIvnBFopl/xnA+fJba7XZMQkNQsz/99VKWM+rrSu+NBl2RZJ/Av2
J7kLJEFMQU/enCo8KPFg0DCwpbWHikmxIkBT7/J9HDp4RoMIpa+tcUkaaM39CJv2
RQf8Yz4KgXl0HeJq8cHUGSG2HrdLKvZfWsI1qg4Dq/u0a99UT6G4uq77G0+N7tNN
FBW81Ys9E1Nl3rJ5MIp/OqUkFn252Y1vb7TocKIsMaColRlVDkDqTcOSeCeK3onp
Bqa0dqpGIy0Onl9VojjZCpXbssbpZO8AHaqpNC195WIivjADNgb3vyPg5ybs6RiF
i9sgJxKBQYmOse8GPLr2yCjZ93wPozh0AYC4EREsHxP9Ou0LaAWeOYyW6gk+zpem
kUywT982J6qsKMyOCgPPxerfZdSQZ/jOffxzVCoU8ixWnPdQcBdcw8mudLbyTNtV
o0KYSS4Ve9S9JKwDBhskQS4/zjsEykyXrvvxG5h/XikdF07BMRDUvUEcpZ9ZmA2C
qNVtR9bCs6X4GrLd14OBb6Bi5XB7YtcKkiamHeMsPk1Mg0BJ6KocNmcaZrtCuTgl
unWHqyYKZQAtUzfEMCeo2YazVtsM0oLWW90VhE/NLa9wkqIpn4fRIb1wkOhOiGS+
Se+lot3xnQwpgnyHaz2uAo4mNVzCoKpBVI2f23FGzq9/wpoGAbzYaZ0h5F2QlOfy
VvIw1lL1dalFOhRZnSWDaQ9GVFWF0+kh4CAwZTEBPEA9NbJ29lNjeLNWBdjzLxq4
UjXJpInvcPAgUKSjR8/DjEoA0S8cb7i6cT6SDWqhas3eb4G5S9/ZJUo6kG6vm/dQ
NOut9WIDTH5rmlawyhWOD9ewK12HlV1fjKSLyuXrkJzYXrW1VEvnyzqzC3WNsoN4
//88haDHPMq8jnDpdSHC0OalCTbdAayZB8CVCrOuwXgp7knBfHQoKb58WKv/7a0t
GPxZNKKfI1SfZE0cB2Lm7IyoXX398De5G96xHqq/P1C0Palu49RcZ0vJkT/6lrmt
ibtkNNQwfdHnyvSbuclKCqhneUrXnBFgqF2XRgOCaaFyFyt5YIo4Ee3QKeaOmrHw
IIjQJ91Mza11hV0E2TnpD7GQXL7MKE9rX0+bKAsTQBPERoGVokJ4UBOAouqfAq/j
dAbTEnk/TzIiZs1LXEirjMtR3r9us84J+qtR9GBgXFONpCPQ9djSaHkJDFO44UwT
64orkkN78aizO0k827Bn0RVMojdTEm7ZKT+LTjgZBdGXh179kDDdL7ou7wDqoGep
mfRzaDyHZ1BU8eO/FOGMoUGQfkxnzB6VSCPUmprcafOFUxvHtgFCPEbLP1b7bzJW
YCJDp8yvux3ET8B90d0ZzPQP1FmKzjyCFtyJz+37MjfQeQZOtCKiL1ne/jvmXoct
URDhJZN6MnUxZF2PLHp/qHUE20TYGvEYlB+6sq1debuu4LzBiiu6Ugm0Cd15mIvL
rpd8xdFCj8MLewBcW0ckbcAtOYQFUXWJk7SiCmUM5QqyigHaZuH2bzdx7XpjQFZH
O16vZq4dUa1czfzqqpU+o55TG+q7lkwDGuVCjKix25TJg65u4+9WFOnjpCKic/lx
SyTLlCUsZafSqE3hKS4ob5NT++bFxKFoSP03HAuFE/41/3hFNUDixMPibmi85QDz
h+HchXHdmvsRPZ4ImjrNsZrhRomC2+ev6BFmANNiD8kxuJOoaojVb27czWiHkT2m
q3HjLCmqjNwHql83A6KYVVRPJ1UzF7xeShghq4QcAICHRCKUOFkBXWvuF8fUUecL
oHp5aSIwi8YpJfaF69i74Rulocr8nehi6EinMiC78Ct67FEvJPIC7bVx8H4dOdPp
PePGXeUz0WDtAZHeAGOsAYRwL6f6vC+dnR0DhOsLZ/CyOKSBTjfkNVky3VC9i5b2
vIk1ExryYvB8yu6H7Ww2BkgzJVJOZboouPEjWJO6xLVJGIrKbX2W4MDnkc5Oapfq
p50YFQ5wXqly8vkOo+xfchLwxDoeQWolcYehhgVY4Zvj2aJicYXk07D2KGoeJyNM
K6PmaQgD8Ztl9Blek0GTpz6HrL0h4n2RAI1fPKoS6wmEIFwH+2ijdkx/EevUAWWJ
I5whdzgBYIwrNgLN35J2OItAKk2uLYdAxQsx/xlOIqHU8GPDEOQCmSSNDhDG3e01
H2jzxLzIce9DVG8P9zpw3C6rW/cGiOm+Y8yKHgFp2Ktl9d5LXKSW+ju3ZboLgJuM
4rXfThe3wRG16RxaFkNKLv5vZqNOeuRSU3C44Mjx9rz0pXBSK6WYMFOQrsFJvq2x
1fDNRGJxKPqVtC1TMpyPzrbZqzwi49YXecm3kGhzUc7isC54HMGlwlaCcXB8VpSu
3WrHIeFHuahzX4YjdL8z+PYN+ikwOiWQGoI4waPPOSOGn5esx0uThX6ioOnCJXVg
VJQdUWzWppfvtD8A4wWeyJ3tH5xITYSwZGGJutuLM6QLJi3v6mRFmy1cv6fvHHc2
+3EkJECy5av3aSD9Pqqp/CWAzzWfJ97Vxxlo9kIFaGT1BaRWb5ZIJNv4DeHIxL0h
WMt9Dbm1FVnP27w/FtTlM8AErOHKs40C+z2l9H8nhj1jRVEUJZZETzsYn9qBdrm7
2ndJOnWNv+R+CwD7as9i5C8P43gRH0pDBTAlYHAeFBjWvYe7Mz0GHQeZULLCi8Va
zlgcOQCeZl6mL+Ik/JcHt2zQjIOyTwNWZoyMiPfHUw+Ispl4NsrRcip69uKrDmKl
+Y5WO5S1hD+kenXRERjRkYpDJ3HaajYMC8wMRIx88SKIKLYSRNHA4rj4GPho+W7J
gQt3WtV1bGUM0H66ZZuUwH+uB6VbLNloCd4ZtuYoHBhH0D0yJhWXdr2C7Itu/fIo
hjThhTaY29d1p4lhtL8u6cL3/7XZSpveX8LKTwy7WctvS/ddHCJPt8/T2KuohZve
kOcsBm4tI6QDD8lMsJnsYxUb4mLyxN1GCaiDOoWSAT2YIbzXN7jHuIE7y3NWmYmU
1G0iW78prNvshB4811swAduy+fvOhEvehC2gmR3eaXCtEum8Q/bHrXcPuuyOWJN0
7LF6l0z7XhoOLU7rWMZECTe7JmbMl5x3l0Gd0jsfbHQ0uMmIrFVApxxtvehES1I+
lU+uzNDCx4JEPoigU8QfdqBR+k4I7H90v0Ijtpc6K4CadcLyC0maIJ0VbyTafitU
qK+rFjMi/ZGDAnK1v1NJr+PNIbDIP35CALJMhNB+DUrttwCIASWjq9wiFdTUpRus
d0KKlmukrVwAyVXvwCKIKYRp3wtMfy9rwxbtd/+TKcIZunJVP9H4w3obqycFzZnY
Wpn0Q2RddNEclbs2u57yqpfBhs01imraHZ8wXIsF507ArPuJ9zhcktDmrWuOb56+
ZoOTEUinl7xVJ6aKu1g2us6yDIe83O8+JhaBbJz1dagNcAXCOqwdeK4Zg2O+yaFo
y3Qen4pjcQUAeBNo67y6EbHGI98YGgb/Z5x7/GDcAwAVHhw24amEBVPnv6GTAYnM
gH9zMpL/TLEHlEoFLsQR22z83xItVw8bdukAuy7NNHcrHi3ljR+SzD5A3Cs9JdvL
WDNMHnmFevE6LgcwHAkhzQrH9ZrFdETHVXCEB4RZ9Uo0nDk+Ux1uJzgIbLRIsAH2
xmrDWfX1VeHw2p7RK/ENQDYBFTyDjnThL1fILE7jYAeiYUaxGjsP5XXrLI7x1zhf
w6nhV0q5RxJZ2Gjea2cqqQv/B1wlGunDDCDdkEjxqQDgJxLl0PkUUGSz77IRaUYf
oSwBoDOBhQQmR0nQazfs0cK6oBTqTmBTcpu4EN7V/u6UrPEvrhDlkDkhoEPkGkYv
5l9pBL3SS05xm6w0X8fJ5PO8BCAsdzI3iphC55qLk6e+6wwM6wtmNkDjsC4XczlW
VUcNs2IAvxMFhAAV2bw5h1NliRpKSUjyBowBAHPZyx3Zo2R4Vq3zLS2z+myqwCfy
s4sQ76hF9f2vsHlLkpcjhe2UY+g7qnVvkvNMQQejFWr+RAU3v/cYkiNIGMq4cBp+
3JjUeqHdD4jpriL281cG3qtT1KxxKcWUymTx0ntjpuAH5f/uqmhn5pFzCj3G+u7N
bshIkKVtfF2K9Zx3rGOz0nMmwSWj9R5yZw+RfIG2Ul3Bm7Jz2xooaR1cBdlz7v30
7x8hmWp7yW/6FzPBWr64zhL8vn9ggOdN5BP7xSEwz3O3ZSWplFHeB/v+dZgRuyjQ
U57i50F5GyED+2UAJfAdeWUChNPmghsfuDyRGa0x7VtOOn7E/MDz5rdwN/GOKTle
dn+CLfwpZKh+VTnGngPS+EYvSkjtjhYn0Q5QHvdqZ7iQb6RRDgVOO6g3f0iI7Ezf
YHXsvdP8ABQKS5dJEbU8FU+0XOByHJsSw+oFm3+/6DsXH1LPDh0lcCZo+wrHS7Kh
+/ftiNH2d0dEyxTX4NIsz3mWzRSmSbypo3r1U11eeyUgZMX+UMJiVhvfptM+pLtq
mzKz5bVq2kWCrvbvoVh2rSaLfyGsfUAh8HxK1V6U9MaN5yZ8HPu8UBKSFKO8lmrM
0yweCjMT5cHrbpzRsfYn+Dk/ZLX5/nM+AMcoOHVgPn21zQ9ohrvHYHfbb4cfBtHG
36mzhTsPV6JVhK/VVjuT8byUA1lu9Goy+xodwm5J+Q5h9wHkfF608bN5Y+qxfW9D
CkQvDg+VL5digbpjTrOS1VAHWq5EcLg+LAMAiATpu5JN4oEQleRRkvbbGPTqqH06
Yh6EvSNbv2eZsQI/0KvKPNRqAKsa9tO47zirCcUPRZzCECk+7NOkcVIcCN7J4L+2
zGGE6SDf1W7yP8IvaZFg9yX+g2nO+QHGX71poIzfF2piZZz2UoErD54Es8FNMyVt
TmbqmNgpqS7iDEWilytoN0XzFPxiFv/NfgnNlHFus9QosJGUWxOpflRcobT8WlkS
173Fj73AEyGRvGuP8FEQDrVtG1+8CaZNK/jsd+u4FEjS4cftu95pH3A/wA/WFhys
B6RKffC1dHm7Cyb6b6rn9kUfqXgPrviQ6bCRPMoB2TXEqzjt3rXZVtsZXxlTc9hk
EjkBVVCAqXUy6QM2j40NBhRfMatvgnnbmUO/6yALQEt05RLlYQXMdNfWSmasP0zA
XHBk9CDarOONKekbxgSm8VIiMmKuuYQi2LyG/lizeHkKjW9oxdZFk7CZryDhgROS
O0BoehYSuaDH3U2zfko7TzrG6NXtlLzATPbaEUOFMi4XyCJR5/qfsF+ss9qVtliR
SSOIJSH+jbqeDOnKXquez/Ibfef0e1QY8TQsG/84WE+x9plQAk56V1eOkI9FU1Bf
EFWY6sfx9oorCMxqVGbhi9BlU/ZnBtTV0c/PVELo9kwTqrG0BZBy1mN32vb03m7o
iFbn5n1Ois+qAbfx9b2r3ePkg3tnRJaTXYE0Rcxl/ILeiLUuPDlpnQ9eDMNjS8h3
sZ3P/RPuuenQzU/jdTTkYqxFM+ruTcFeWqpAgcnXV055KoPBEL/3ANC/b+c8cJLF
dbfbsc8hedN2EFU9xDx5oeuAo9VZ9xoIHxmY2eD04w7zmV2LW9dbL2QmG08aY75s
cF03O9qEZJdH/OH7EVDWqfrq4Qx3zqVIWzs5aX31lwcnKJz/K6sgLO3M3L/ItMH1
pG90ovrvZqxZlCOO3rc+AU7hAiegg9mSkgSJIhy9X4kXa4U0ujJsa7ynvddplayW
bv1LMkDatkEjaha3Q0uHvzc/ZOePjcw5pJmLNFRtsNWwOWGsXuExqt5ZIi2pIeaL
JUZ3A4Bd1ajKwvvh394VBKUx5F5e1DjFblYux2ngddh2Jr8b4hLGwS9zKmgbzjZ9
GIts1chv1HD2G+1c6xZ4GS2DhUgr40trUQ3Nri6eGHYvas4Qmw6164n6naQDmZ4Q
1HNjJ+hKCtP9/fFGJ+Hh6nLWHk8UMKJ3grx5/SmolHkvjIkmcFXLuWE0dwDwzJa5
L8utG4GgoLGunaZJSM0klNM0cTN0stMkw0ktssIBZIAV4iL4ldZRh0Ay93SRmnU2
+hQjDTVx/Se7nNaLEPjiVkB0/7PU63vb9Bok+cLxDsF5kLMcnPiMwFWf578/7iWA
E1XtnLinrUXq9wTUcA6OhKZt1ls+vYg/tiHbocZUteNuBSoebALt9VtQjXOdchVb
xlPAbcjULGZhlUlgcwRANGdN7Dlf8tDaAs5/F0/XTB81rVz1A0oSdtjlzOHavX8H
QuORGyQwBixggZtiaayWs3ZcxtykPFOCYSt1RYDUy85vfzQLTJ2HMh6jKdw2W9zL
7U8A303hHBRJ7WK+PecYPVRcNSZDOZ0FCFeedKAQ4aYC/d9nu+Nr1KrQQPUBvvhq
R7MGqEkirGZecH+keEFlAmLnhRHM80UeuqOmb/bZQMHhdR7Hju834e5WEJoJNXHd
f6CVq6oOrPQpvCjMFuVbx+dh3eOK7HERkN7teCU6B2BAl2+QKSa1XzYFFidzGm2z
etmiTlcRmzDbcXH90xX7DEDm2CFoZspv7Ruoy89nVTVXZnahMFqZYsduD3At8UAj
b+6lL8Ws4gFF7d4Xhk+dR6DXcAFMfX1ONAfAzsyea+5yZqhlouwn75y9mS3VLeqJ
9zEFriAZQjY2xsbvSyFM7YItoXArswubYtQAXWz47TvEEsdteyngcEvgZuqbN51M
RROP6P5vgAM8yZrbBQZ7tBMmEsn3Gi/Ob1pXtDe8F4rHjogm37UMsOASFWw3V5Ys
PWRKxBtRp7V77aRjM28NZNCO24mBVVo3OO+zQOafFEt32tcAwH24LP4Yg2v3e1j6
Gf3qNzDO+D4w0nw4Rr6hR09kV8gkeFebue9QwumRIpGB1Z9MD/UPDQNLIDOvrZZj
fCs5wcDRKzoxVsUr0nN+NCMl79vz6mqv3tgtzjw9zk3QOQDOPqmE3tBZA0GktD2I
lnbb4TZVw75W/2G0RSQSCk2FsSo54U+GDvl51N4Yl/PaMvaT78adifK4GVIW5BdO
E3yKoDTv1ekCw5nfmwaYuTSBf0/JJ0d76Afk0kUYjCSLI2Zv5/AI6U5TczX74BZ2
bzoI16EZp5AAxt2iGRO1vJ7zhlvONQf38pils44nTaMNX2QbQVgDMvZwSKvVI0tj
fVlYkmQJKx0SHnA6GJKpza6dXiXxsEK0xUa9f4xrINt2OU4loPMcIqUIX8W2m6o5
xosvR1HHd/fWROMCTASZ+DqlnHmbYtSKfAZbLiSyb+vkQeUyWMimKvA7rANksK/U
CYPIFcT/BKGUOhnTILhPoZMHmAbfX+0++StTQH/0McjpcgVS22SUGLpJ5vMhLdb8
pwU+kX0B0gSDOWfc6p/bAFsYps2nGpdj9wL2jPObsCVYxQKKqKqodSSFT/GL2v7r
2dIao4ted782CToYgMyfaPLiRJ1LikfVNrMWPluNS4U4vZD0CwWl2UQnReb5KVqi
/lHUdrbC4QDnujCwQwhSYbNOfFnhCvWBAiYoprjmh29tlE4T9CmO8Ofz5jeWnLVa
CJo5Q4o42I/KEdd7DXXn2Rzd/xPziy3Hfj6t/24x7FuS1atupdI0ESngUDWBsMnM
/N8PNs7HQnC6YZEfSzpYnm+dNxH9PdyadfWiirYGlUQz16qPsBkt9J2gqYffUbIv
WyQz4ZTn1xmpemwnVNIZYB6khWeSxj2dm7Lc+6eWUYWHL9AzdBgNFnld8fZHfQzv
ekvXSalHrIcx9NTqKdsHDOHKLpqIvb8J0J3VSVCU8hf860dOin7RCi1I/TX0C9r1
IBnf0rd14qvk7igvZBHWtbwQt7wncm70oAnNU4Da0X/Io9qkFAc7NhP++hcLgywT
MDRg913bLZx/PCcDmyybRD9bwdCWrS844aDniH1RVst05ingoQx2b5GLRdpM5x5V
YrNvdk+O8ZYjaQWF5Enfyvy9TKp4RsjMfQheurfbCialZLlKCSd3gcqojkXAjcDv
4PXAW5Gzjd36fgdBDtWe8SJVf8pR1NY64d6KxyrD+ueMkuLbEhnxB4yocHwJmXHq
/FmHDw5idOzsWusPaeGnynQbji3VpWRsZST4KIUw3DeLWlC6cOLuIswM71ka5oQ5
u8TY/rgeIrlwurHNAtEzYmFcJFNB5shJfga35wERtg/hi9oXIJma4vB+pVjOt9t+
8TvAz4BkdVSHUKXUWPJ8ZQk0Ypvoj/PI136DcXYJVUwbdV3/gI8uuRhVgUjBHwkP
msCvy4ji4uXErY8OGfjqN2+PZb3747Jg66ycr0elrfDjKXNlZezotNZg0s/zWDXP
yhflk5hjphswijY8xU/rWV96htJANMbrHibw1TQD3CodHb7cKRcVYpygnshB9+D2
Gqf3MpPsw7PYKWl5nJoip+QKVxwaA939yo99P0WrFc0nIlUaV/E9gwrG9OLkW6Z9
6JdxdEVkeVl/u1+doW5VuTOwesq2p65b4xtx4ooMqgXWdAh5qyAStCc2KoTS4iXU
y9UgzEMMYn0REyiC3U0iopmYJ96HQoYy61dloUFK2Fsq4UiRYR5YQjLubKgKD9WU
jJaU9tCiYJvrCKAHZSkCj449cbDqntigO+I/ASnkTu+/PgHqjNyLTntK/gpwvBih
0Dcx4pQwWLhxNVh73AP4mvFNC4pNcxAEFTLPyuMTQEY7jVUlErws3ly8wj0cHYiu
5GxGOqWyTLI11Y40QGWRYR3wO3I+x1YNxx22XTFzIjFi0azFND3EZAASw+meG4Iu
jqvtlZUnbXTaUgUUFoyYdxtDlIrSrt3zJhzBqT9JrxfwaXzHCJ6lWeOT01xLKLzP
jQaIRhU3HOn09rSz7ctGQbippNEW6b0g16X/vdOBLthwit27lH3IMNL+8E7QEWsy
70w5DWFJSgMmYDR7Mn39hl/bKrZE06wivjjWuMqu+D+UN3j8ODXSBVIMA6jwmC7R
r8rSpGdkj17O7RAbBXrNNuLfimYlWk3HZQdroQvG30vm8xQr+RrFk3vkRTCcEPej
qmFM2bPHbjgYONpicZeWt0fraNCpAojd3LGbWyzjOcS7LQx+Buai5MRtBAn9fJ4j
3DncSFKEw1PGMR5bicpbPCDQKdN091cazWvWN3b6f7Hdaus9nbYfPzpTSnM2XWg0
1U7//hu2MJdxwBWlbOcfEWDzVOG0Nh+/BvwQcuwJh4NGEa9ayOv72k93n1HmyToq
fr98j2WRGDkOcU1KIkDFJjYOXo08YVTkc6c1q/3W1DwnFOr1f8BQxmGgcBhXU8Rc
FEyxzL/IxyBZqTuGWijW8ePjfdkfIC7+/KkCPRn3/dDXlftr6PAZVsDCv/QRHkrr
ci4k56y2qnD3Ck9DBaCXlfNmY9da4k2tZbyhQlN/aKRvhDUNm75nEVVKEuE+kLFU
j8XyW0EKJrrI3RSskCiwWGKiLj71lRT+gwzBHH4CTGy6AN9bSj8h/GgIvscTdGMc
hT5I5znGPOjFU5sW7L0Nkg4y//JKcML4K3XTFZwn9GGCuAn8btS5cferJ7Fhjpy2
wYrvku0efffs39BsPOe8KDkqV2s+k+wJ9PX2MopqgIxeZhrxXtQG0O2D0Fikl7ry
B9j46ylT0pGvhyxaGGBUUmPoPEnVp276YqV4TcmVwJCubh5yB8WoVS4P9Fi59kW8
giitXXrHyhy3+b8javk38wG4Vxig3QNXxLuJd/8ft9kvnC3SBFFeYDk6YmJJUOG8
W6fG3T5bhjawdh+I0C79V2C1bcYqr2fVGuX6cnyklr3VKu7BnHx/U48KtSo2Ox+c
kmW3GPoIWh9b02LNAuUiZl3qnhSkBZqa4IGAYQgDmMEqW37okN6ZJJI4jrRKVy16
4LdnrbBcib1pkFmViNOGij3F9VRaZpDqLbHN7dvgHC/3piajgSFUmKvT2GRFRmUZ
VgLlnkmJYAIERafUsLBknxMbaSvKTeqWl3Juto25jtgp3uagW8b1x5F26eRvBee6
TFMta+ZmjB6k7QOw5N03TeOQFJ13RXvsh5z+S8lV9lqln230GD6A0NmQHKFQ6Hhm
qmrLdOBTppvysjCy9yU1ZFOmfTd63ELk/ZVxDHx5X2hvgw9LhEFSB83D5XTO9dGh
NIatckjK/64OrwB5nmYLNm9k0Vr0yq8eVCdS6z84tTX9roSzl3dHbB6ZvjyUBAH/
6QeTfNbcNnZLJUW25my2UWyN3f20/T7zTbK6slnIqm2r76DLEujbQK8BtzhWl3d3
A3JF50yhgbEKtPxM9NaVaYUzmtQvaDEAYxBMTw/QhIpBjBRAfahMpBOwKXWd5Z45
9Cph36SlJIZibud9fAkEQO0fOJm+I7lGTzMQW06bWQ0wovYQN4oQ7XMnCBYFSkB3
pDOV8Xf64bHtSlXxi3zDi8/a4DsTSfiscT3I7wWi7+jeqAbJAYQSykPF+npDrS2Z
Ellvm03eyTPiE+Vl/+qZxHlb7gRdqopAIAlUwPg8BLTe1aHrfDikqjd/hrHcWP0V
EX/COZ/fz2tdqr/NTH6T4S1pXZV1XqjwY5zTRs7at2Ve93M27e0ozpOF/cDjmOrO
mI0iqs7NsJdFcTn4ppKC+OlFthIasSB0Kcti6AzRMJo2VN8PayLUhYwfhwgBxJL0
1/41Z6CWhpLAe9WN7a/805ngCWmDBAwpwgvCEH9fAfdVr03MTXre7xlc3miHTpdO
GHDcRfUNB92vMaXRAWHQy5GhVnAnE1eVbh3Cg8EkfjSbToq/AVSAOKAuhwMuzQEN
2dQFmJvRdssu214kJlKV0/TjH0hBDfvReXxop4JOuwuJptPbFxKSQAxEuCJ6N5jr
P4A5En5mhjT8aqIcN8UV6X5IX9HqstzS6QyJ5udhbowv7fD5y4vIqV5Vt5CLcFSE
6VH5jz8XD5U5//0YWEkU//L9LWkOI0n6FdtFyXhZfL3XaW4JyznAK8xUCnRilw+1
MOjtEKkEn/wVEv7DxcK/I0ivlBnx7QsPQyto3RZ/Rua4N9xNiedaiUNf1NAskZZd
+n3CDiCis4sjU1Nj8m0dVOC4Rro8rUUwNj/TbXHvzb8LdFCbhJ8vASGnK8owFUzM
zTRV9AZc6tLjDUPF6GXL4WQ28nEhfulljVbO+5wnrFz7Bp2NAxCiCcq7L/BbTajf
41I4i16CQyte5+yZ7tdN+9gbFh31KbhijbDhHNqxOcM3ehj2AimNIxeg9zHQ41pc
2NA9wfbVlvWGFLreCih8AX2WOXfMT5JzQ7X2i3FVFFFrSnVbjlEa5ok4BPPZwvqJ
E5WsE3vWPRPnT+ZJSapATqBuOJLJKMUFwhN7ttVnEcsdrHswKt9asI2+nbLvaQSt
1qV87Uho8h/GE8zyFkrvR1NaguCaMwVF1EGKZn6Lklub2eqmXpVkAQdvjQgi00uQ
s10bMNnxZVqz9bncUGv05KywFQYATauQ/jUKOlPbX0Pcz91ih0ZW3HxeKaWyTIYd
yDVfu3R/tL9SOdCPIdjDDItabAlX3Z4SzCIQNyV2A5PTy/gafRFLmE3IDV3b2Wb2
NnPuHd7LBRSE7ZNjWqOUX5d98/xA3HSCcalK9penSDGkgmj1PV33fsjcJgKJbQ8Q
5PhfTrDuOnfs8Q73RD+Ik0/l6A7Z+IeTv7kzEw9VVkglwnngQdAaJtyC3T/uIGJI
1OJVJ0hcWhGujX7R7ClgtlALCfj5xNP/X2H3CdkibhsHZ9bJDJ/ChXzC0iz6DU8I
Cjc2dgsZS1EWWMhi5/RWUkoOhmig1uoo5g88aow+zfBXUVZfCGPB584GnsmhGOCK
fn6srJk8aS2qq6YhHSuBiuUsu4Xsus53H4gwRiQ6gjjNKMv9JyMIxr+lit4lJoGg
Vm0irtt6GdY+8Jy62L/fuhZD+nzP3pPTOlVEwo8iUZOb12A5EXeu+G7+cm5ggkE9
v9zUqO1apienkGyyhdIKG5JVRP6dtcwmdMM7FrjAAaN2JYVfLvE797HzKS1v88vE
7UcxBB0oWiYfgE0W9bS54hiN+KAafYPd4ZIYhtRi+VLkONrlup1Tj2DWGyrAwpIS
YgqF7mRiAykMFx9ECL3l9hGqDZhEfWP1mTkpT4WBDcEEA2b689UL98qIoKGyRDko
aAylgZMqtbQIX/OFc/F6hQO3z8Snd3vnDDeHeyY4//CUPlEZcyPTfprpwwWdjsXx
t6wBidLbjAWV3AivisI71onmRzTUiDNVUh3cnEbjbB1PiqpwtzcB1YeTilj0TW0+
6I+KFcC+oHFW7aqQYQLWKtxikQ5eleA8zIMHAl5JOMaDHiY0y5C4o58MJZ5afY1d
dGP8RCJITADPWIrx6BIGf3tvhycgou09Ai5EPu5EqQSLrDv8p95M/xLPxW5VwkVK
7Z632KIId8VyyvanpfXWKtoWaVrDKujXMzke5782V+lmkGCwcoh08LqkmqO3FjR/
pZNdz4JEmP3FHQmTTqgdtVdGkjAlYB8pkDTCo7Id4IdlF6XExCc09LUTbABnjx7S
j0fKzMfYPoFy/+jj0NKpsifa/sX7ZVfrHZbkTPhyRPWmI/f03IWFhOarpmhc+cF/
OlKuxHYAbXI3kdecSKWXI5pBQBFmGndMHgAh+7ZFQKssmMRWBDM3ULIB4fXiEtfY
2Vrh+cCK9U/yMtwVgNSWMJb8+Y8FhwMCfFdXJc5SuF02mE/qcNxMoUmHF4KRdEeB
l0QeiyXc/kfaSjPsP2VpCys4gXpkf73jMdD8nN0huYNQvQUZomKYMmTD6Vx5bIri
nKP4k5YDUHfmpMYv3eQKR961r72q7yZ8WboiRoIH9Fiiwy5EPVDNU9oHQ7svAGor
+rrixuOrhMK0653aAe66/AAkS4jMn+QuvU40Jd417A/D1VlJO0wuGTBUlNVYwUu4
6QYes0ZsCp4KIbRCzFg6atqw2Ooszx7fmEfVsjFbA/FSAmnoduJ9xdkqBeG1vk+D
znRpeqVqGQDq57579scSLEKRrAdnZEofZSJ+13uWV/bCxU8hDO2Dix2aWTmY754y
sjcQV/BC0cysQJ5qVbM+oDA3EOYXplGpqV009nAYiRv1m8e0FF2XlUvYHvcMsdn1
O3jas7Jm2Z04ljUUaLPmK/aZEYKHiPZTrT5C+qt0kKdVAFLcxTQHSrl7rYHqmJVo
lF5F7bvKvhB4/8ullNIiE6neB4aZOqfxX5nLEhP6H8KzsD6F2DVxOVZKlJ/so9HC
MjTg7GRFWWuenhXjNvze3d/a4XV0wK2+DyzVyCVNAMx4MGzEX1ISBjGdHMmueRKS
A3uiEoaEP05kC7IhsQqNFDCSZ0p7olly9Ydm7QSVE7G9NodiI1lBqnUqD98PyF7E
iWJBhNT1svhjJ6L6927at3ApAx9fsZKB9YCSbwmYnJiyZvtXx6jQ5bTB9jSFq9ab
PWR12DzmA7GwjHOssjVoqVMZeARi4Cxy4isvnxesGFl8CUVcnDHeA0q1BkMt1UE3
lrtoIzdaAx5iIkPrI4M52dNFUzfZZK95VfKk2UibUG28cMSAv0VmtKeglogn38UH
BFdKLtFRP+mNQZ1UAQ5KJS38lvrNNFEku3lq/MxLKyu4GPpqvWp+bKQUIC6y6Yjr
kKfSfoKk8dPeDmBBNh4As4N3GEWEvCHbOVTajwSn0Mq1AQaga5dl1c4mt4jhdkWT
nzE1sD5s5hq5TeANUyNHL6n/uVKqXiDn1wf3JgYXdAJ0/pkptXP5tfaHE95NiTGc
ZE/rarsE86w5+rGCXGurey5mSvI9KA0+bLMznawoXQavu6GsFMrGFkHaMoCM00tI
dfSbD/m497y8oGiVkI1FepmrLbxAUVg+f98uDc/PwNDWrk7+uz9NGVjhliK0+q3N
gXu5VHS+1tFfvzht5bHjCnaFGYOsGq0W6uv3ZcOqYWIcN/9J7AziOHkmdpFqRwIh
RoKetjP3GIQCS62DsU/zeh29m6t/YJZ1eh7qvejefur4qMDX4aDCFfxEFJOXgCfh
bcgsTFCBy1tzDkpxJMAV+C6vsOvUgP24eRrzCqN5XhUcM4ygbqyycTO9gfUPES91
Rhgn69+9XTlRu8H6ghodQAm5BdMgP+UupiXsEC6TLtXsDyvsLSadYMtyMTkZUZkJ
KDP7xaML9Bv4gsZvJlBdTIFq4da0mbM9EYaS4gCgleHj4wpby/GNWQ9QzD1tIQlx
YZp1dMAfLqo4ZJZonUIL6gGp+5Q7l9RVDQJ2dWvA03oizEWEEZYrzz9HD23kb/t4
8MVERZyCO5JG4oBD/btHL79saTiCi2OeyfKdIHcugN7On/Wf+l3Ke1bbdwaQy5IG
XRqKVvUQW4ooMyLOXZ/fz2NtTSIoCotgob/oLf9RvUy0cX5g8Lx+Dpj5ghVr2/vn
uN098XTT2XdzGOKzfw8qljsX+PJYHMww2U8GRCOb57h1cssW/5vZby54d92E87Z3
x6x5Eo4f5s76GZ7gzeuZl4vd2YeHFwjsX/uoYqHHeGWu7yB1NZLwxQGyPneIjzcz
NnRsAfBx4VZi76WvzwfkxgfWm2W1hNFqXqZgp9sGygPh76cAeLpCT1yGevik+ORS
dDGQo6j2nRiH3/G4Mrcy7IQ/nnK5qJok6/BjyZ2IJiz4kcP98Rr5fvfNWmOQJ52U
8vikxci9XIjGpVnMyWtW/KjX4IEIR5SHzDd1X2r0X6QrX8MSMcRcdDbQGmYZ0MWv
SfUyi3wR314jMb54M82q/fa/KeapSQJISfVjm99a/Tw6eV75mUoOQse6FGoTQDiv
blTNupL/DRx6i2NRBmFvFN7g8ntNf+KAKyC86FV3u1gntL6J/12E0TFuuFsS4l8W
nnNI+dWf+oQqy31ILFM4AxKCKW9V+Fr8vzDUrlx+GuZ4+VORBF9I0SgXNJFzuivF
KYhoaaqBc8cjXdxS2WmX9hwXRZ6zD6W7vEt5qxJQwX+qFkP18vpWk4ylzHWFPWBg
aSsFlMn1SFKm8zeH54RCXf+2XMgx0ABLr8FTtMqHIobT1U83+6ZD3N7P+7LbqXn6
UOYlOOBI/5zUT8k1v4AGp1709DNBkBvVNb2i3jIYZoL/ZCAIz0rbnPcu4Q3kOoLX
KYKt+C6LPPtUItpOfpvonlXFnjOzatqnlou0eyuO1DmhV3Z8v86GNfWvunVpwfVJ
3woFizJz/TWdmPN9JUzLU2N7DnFnO/xDGESIjNIv+akfACscukmrIzr5bfbLoE4w
TvGIx2XaSNWC7DZM0qJnE8JbkOa6Jv7JeJPwj9T8IHgNzocfplHgz9lf9DKnvxcc
9FOi+mxhhTIDzyfzXe47RNvv7+PqpdatDB1uvMNF5xpz2YugjFkrl/18GMcxEavw
7bDTH4wXRmbvKxjvWuj8ieojgAG+9eNpIdfnowbeKWW0ECgVuLl/5VCVtl3YTt1w
frO7K03YzbRC8ZAvn44Dfcm0UuLTo54i50TZPYgK9Svet4/05SzoyiQAiEsawvYT
AtGYsbttnINCYhaI+e201CWiH+maM0RXGqwE4GrtYa5TDaEQjSEVl4WtUykyxOxJ
cdV5El+2bI+JH4tL6gfuo6Eot60sqpdMa2ZtmWU31Tod1605V81naoMAmzTh0GFK
qG89PWYMKr7t2KbJKoQW5z6b08YCs6eXfougT4PTXV4m+FMIkKZNoRkJEQ46fhUf
x/XXiZsQPCqsQ9gkT5k0/O+ntbB8ZX8P7mVCXhFwYBSxf34C3a5hl2SAoNq/C+4R
+3dA/SNCXpxMcE5Vc9TTHqDqOc7YI0H9VTidyM+4wD/T9BHy+eiAUaq1V7wsKVkz
WxEcFtWvcFd4ACf3KxMDWHwftCCdq6WYasrZkQxhH/vhpJJkHKA4D3TdHWaEFakS
TnmckkOBT6M4UZamFAMGociEYXYjW7snik6jjmQIh+yps6zu9SPBOJfzPDonuFWe
hJ++j1NeI4vL6Dgn5WrwG2p9o+F84Csb1pOGtpWzPESd1dE7kPdqZysj4IAg3Ugb
gYbWMBZg1CqIJ1IHZZuM8IhQyo0kc1zK0vvhSk6O1lojYJj60eybaXK1kQX8hA7y
p5nErtdkLR6WcVfHdY8ViPwQIWGpWV0BWAdo7t6G0mMm46j5aY+nVKT1xnh89DzC
OAw/F2GmPwYmE9H6T3Kqn+Cy6/9sqt+ySp1AKw40r+cKYItn0tOavNUIwtBKfg5G
IGLDNRnumtvbgt6kLchzesIYbLRjhQYNrVNo73dTH65V+oWLjJu4uWCus0K0mi1D
c2jcNQAS0gwUN1+MrHhKpMZCU2lUaZtmCA+HXyVdRRyYTigXs4ngyD0Ihms6eqSR
XKVyXMHp25HqadJBQaXS5YC6gdquXKVrU554cq9k+acjmxwaBLlFq6StMZU00yvg
Gu0VyVjOYaHp3D+1pb/ZwEqtVqHJ1WkvwePRHzQLqyNGFM7aViuuazsmtXjfCdHd
zuY0kcyArcnqC5wSuBjg+x0lLo+l5aivgCd62nLGXy+Nh5UxSzKBoTS+S8lNbldh
40BBSOU5x0NUQ+OoSZnz9hv2hT8wmDZ7gfGn9CasE+E3Due/ZSvOPDz+z+AA+3ZP
u+4zDmJb/Kn4LAeUKz7yaF+bOMQ6lTyE41fSxGPf7zjEBGyUWa6AgV3RmqklVAh/
Ve6YKprf9CYsVCBNxx0yOKj/J7IddH+TD9DMfJ3mIt5370iE2fvALmx20OxidlM5
48oLr/yfcmeafihR6C7Tg1hlKz2Nzh6o9LkUWd+Y0d4/q3/A9xBmDmCQ4qy++9KR
5B2PZC0r8c9q16zC1dwyGb63/bxgq+DAX5j9WSH9Brktrc4DYImtD80ZK7OVWoNT
8vdZlzzm6RVafFsDbZUpyMxzrg1qaToiyF4mS+7k+o0a3/zGHasypasgEDJAKZyR
KqCohZ7MVHkdeUcREm2/k9C4bCt/FEL42xYV2OEx7VE/9xp/9NQzb/rMhWTclhGm
XO2XzS9Xk8vqYI6s37s0UiXG9Vrv3FkvESVN/Yy4ZHaXMxTAiD/3hMIB0GZr1ulC
2WDwaUae4fqTlXRLxdodfabf5sWd5ZgOhsJsxEFr2Yb2W2qfZI+YQyXoRd6ark83
gvr9SH9dJONXboLvJux02JDHZH0AgGfddpVTVXYKXQ7oocLom1I63m3w31iLyUPU
+2aE5qwZj6Q/WbSi+mu1BMgsyOG6KGNLcjwunfzWWj7DIhF73LEqsKonZ+ZoJ6HF
Y751T4VIVgLwZuL6fErwJe5hHITTwBX01dO0EPDxXoerqEa+UvikF5AbvHQiVT9S
R1rGcPoML52ooeIbmeZA2ghlYJWxVyGKY80e2r772jIX5FCb1O2xPuNWuc4l38Lh
ASzyIYzbf2gzj0skoQ2CHXDxOcp7awU308NlJKtmtk19GwtdxNNRsI1o1HVl9j+F
L8uUu/vm7/QUKK49P7PhWjecpt7S9wqlCIFV1UppyOdxyDlvpBlnAkw91gTMCJhi
7RABWMdAZQQQJosV+mzqoPUPsulmy2rVACO88m/p8+dN6L2f263mWjPYwbTsmDki
t8KDVvFKf2g55/vEt57PA05RQ6MhbrKDj2Mm90Hkdrgy46qFi+qTGespMhCcKany
lnuU2BFlyDZu0LmYL2lDktL3JP6nxri0S4XQIag0LXF6xBp9XoFloTAeO2FGYt4n
T9dKcegpkp6v0fl/n46zk5FmEuCMmw9hklnrsa/WKwxr3aAEg96azPZJPwV/Kl/O
xcZ4jVJj+7Rlzzl0GALQxTvqXk4sQ+B9QDiyx1TPNHBZkJ0OnsXG9grlvPxn9o4i
PsypngIKg/3zweNHP9cVLTidwzXeXN6dEvrrTdWjqgVWYteJE1nc0ZUqSA9YFuxK
c8WQ7+Cqo/xhT/MBiM+Mr+b5K1cLD5rB43dZwrXS3rSCy+9GTGN/F7E+PQyIxnXv
+xULGSEGfCKUWpk2ArvaBjqoEL8mW4dy83f5jd/3KM+Cdao3AaYrikaMjHFzbDcZ
wRBOYx4/c2phYNrc5O5cbzOEb5KHWmBCtpBV4zMMbCQKAer9QwVaSXPpD56B/L1l
zouSC0OVg4imEx+ChEbE9y9KY8hg7irjUny0BWtbhfxW+/K2vy7QCZkDUtk7Yi/s
hxAesXKOCr9AynaQ6PZPmq1zvWM4yDF+RfoxSWPBxxZHVn+8uWiE3HTcBidaHRGR
9q/NIIXapUJ5ErOaQgQXu0toWINpY1aWiOErAK8s9hWGqeMvn4BYHLJS9iYDA0GC
k672/rI0X2UtaEiLdR+OvsLYsjB3XJvx2O+HfVPxw7xLCJnRU00Nz9WD1AfLpf6g
BD2OOuDmqDjv6FsvqPiBEPNTezMnBgYL0iVWWAFqAL2dYpmNeYD4HWANN3XC9CfK
ljHwq47+kJThtzBHUyxAcqP78bfkIJV+xA3/hyigJ+dAfr/66eV2RZerr1n8uENN
MLYbCplJCR9xfVwmxIYfPJsIchE7NJVKV9iXVIxWgHN6YyydUnshfbAApcmCa39F
J7tqpk667sHOvUysvD9SKlXCWxRTIe82SsvT9YSGw7mM09r3pScBIbrbX43+ry4n
RIiN8BihrJzOiUWWDL2D/COixkPuR0YkpstmEE1wGRJSGtobI6LCNHHlhTlRoQLj
3ycEaOVqvzVSbOiimq3q8ITO3oqW0HQr4wWNAX8mZgAh14r654AhexSu+uRV6kHU
GZ4POWz9q8RzbGm0OHDLINbpbHOc8ehuju+c252jPbLP1Orr1Y27BCKAdHigPMvO
TAK3uWVV7MksYAk0zWGymqAbhAjLOw1ojv1NhZV/hsVo2+6MhndBwcHWXN/GIeDm
2LEbGHZQgbdwvZ/GIslySLOJb7iXUta9ptH1VNmrPD44JVBvVLrMFAMAm0IKou1R
pCcIXyzfeI+zMA6kc8t6UQGm0W42vvJ9QS2wv9MJmCpPkcpzChYrpFNb03GM5QJi
odzhE4jwKdQGSMtQz+QRnomnqgAMWxtbb77WJJ8mmJ4HTYsmMNWu6l5yx3cU4kZ7
w8Jud3JVP2LyW3utwrClxL3lNg+jv/i+RetwD/60YRy+ghsGm31WYyZBRVgOA10F
8AOliAVyAuq2qpnpvz49eIDMn5LAfCZiKcJd6+riTdGFc4ApIt1NKcDEuUcqLktG
Ndtav9gKKzmYNJh/ajqd1Dq6VCatRkut1zWtR0P2MgwmuoiKRg47jC5CN45XUr2P
KPxmDMNQ0w0w00nd3yIFUPc4E+KRsbSc7FC1P8iBezS8QJov/6dqC305DhwdJORI
M+pk5YVdu8CqMX8plXXhQpppmNefpcf2Zl4tTJZgItIdbHu8R4pHhZImUCC0RlT+
ZElJ0Gv1qvGp1a0wGdl3j3CKWPtelJ0Iaxr4aCr4xXtM4be+/l0a4MEjYtQJpVyk
zlg132OXhN5t6u4A+8jHEHRswMFOCr7XD8niutm5tmGNZreWU+BZFnlXBt2OMYI0
mMH1/uyfv3DYv+6pLb7DWZ4Vm1rWMmkP4tIhlVv5QxIDzzdPeA2jRAE/EHyuO6R/
XHAixy0T9EVGawS5PMCZUdcWo5ROdUQndXUZewLS57rdiDWBRYHzqvpBScyLnlml
WM+bgyR7GBEJlNa+n5XsOc2Ph2I2j49y5Il8SXzD1BsaZyfMGW4hGt/gSIhXc2JG
dFF4xMqcAliJoa9RX8VIXO1+XLV5Ato+7c92johppLCegg3P5ix9jhIHvfqp7nYr
hUYYOhtsEdTU54XyvFWnup8qCpI5QmhGb0djzfwt1rJyCYjJUirQHN1ssiOVLVVq
KuaYneAh4EpxyaABLkEjgBTSQ3flEwEqWBbT+GZ2JCTV9q8bFnRHu/K4QacstHGC
KAasuehBB8QdO5J1t0zOR29dde3OPjD+7FvShkFBE4BAfQErYhTAwNzXUtI9WpjX
3a7dyCSNNf/LmIfcbE/K5t3dkldtnkkXRY0LYToW9AP7ZnjOJtk5AE/DUATlQeWL
dhk/lCk5jNj0F1d1IAs4DLHDRXh53f835Q+Elz9Nw6KHwS4lsjCYBOXPJ5WvRbU8
UyK8HhVPOtVEuu0CzS0UUdvpJb3fqXWx+7dvHsTgfSr6TqxpvS4duTnDdEtLZLry
jEa8J+f7/EGNuhYFSGjtQWf7WdSl/VxUY82BJN7nFowTneuo8R15JFGN6WRDlEgk
1Iwe+5RE9Nx6lEG7DZxMEiFHoqV+/GUXpEkoWMgwePpKHBLjg+pifcbSWDhfByBi
riWiJdPJaQ2vDp1QBm412P8u+hDM1vtSE/oGQmLUaEXM4IQ5iMF/9pJO2JBMZ2vC
0YGZj3alZr0H8nJND9rRb9/YcNDGlSCU0ZAgOMGj60wGRZlrSkWwjUOqTU9prarG
Z65g0moFRJsFQSf8WnyEh02lHk5G4nHO/hkw9pHn2Tj9OKLmrSg/93LBlx2Wq6VH
2ryys7gfaEXJdyidtNY+MmYhopzOChW22DT8t0m3AEhjdVIZQ+m84bjTknGHQ8Sm
o8mlafSyKgtgHwpwgrkDIY0VEwvghTZuP5owfCyxs99qc516JSHkF2xm9VwWXo9a
idnunimh/DoDmAzVDtBTRuIs9Xlkds97UoYv6m8+R4vENcb9oa6LMKT6p/MlmGQZ
bOaeesiA40hdtITrAHew/0wYf1pkofBJ4zqQezwNVet26bLIK2f9fA3tElTgZpOe
ffdVu3vTC6zvb5c5Fr9XFkeBD9bdIu6001JvwQ5rDMwids0Y58DnYRR7HWa4aX9S
Jl9r8d9m5AAEITAWAruNjTaVmVh4+VzAMuWM6s+b3D83tVjahctXxUQ7emQY8jfp
vaAMHdHTRJW3WBo75O3aOR/CxbwqPCtmbbJmhe5sYl34UvlQQd2D5KW1HGnWgZd9
w4BvyBvIDrGVUiMIBYSH7ack7QspqcO2P2L5BEjSs9Afd9jTJgTaPCzus94+aHAS
J8IGwVbgERm44aTNqStmSSS+GkT4TxJuamXPtwz4+KXzKnifDZ/eN+WOl2Sn7wwL
oQ7jExWDa2gND39THkuW8tkdArsJlW8yzKOzHKq932HR6pJdkpmi74ZJrX3rcIkA
kP7tNTh+KZN4GnAgvUv72n4bYnRJsQBK61u8nlrEaTQX2htzwRnRRu8r1sLugQlH
yqjZ4zeIIgTSzLoNZvIsTY/SxjGVs0FfKlyML/mI/+HbiyDJxlbDk8wQp3fPSU7w
CwFZFkaz4lhBlxbXf5EBtu0oYimMhMwggSBgOInDW9j0nnvzi6+keUQE3P/pUuEH
/w0Gkus/SvTM8MibeIXW/6KBAluBH3RdNdeBDm8JbBCOtMrHjjLzsNjdiNwf/81+
B7CrYJ7h4N8a8x7+pB8EymoNnP0WU1PtSOqjhPifYESHZR4AExJl0WOIY8II3Jrz
LrIWDFQoU/zaVvTumtTfkjVMVl1KB418V8t4PBLsIEF3OdhgIS8GvLkoLMQsnZDX
VAS2/B9/QF7xwFmQGrhn75t8vXzJyqNcBkwlncZWZNTq1U5wnT0UNxFSA6QtpJay
61fc4yuR6Jli3YvXmCaJyfwT9sDA63rVPCJaBYgA4KcGwAbUhk0mSBQYrK7asYRs
gPGopDOvt1QHSDpxNzHIlPM0g3bpd2ne+5PFqWvNW1ZwlR7YIwuL2dCkRAou73Je
zyeLnyTiGEq3Y1ioy2JAuyh24Qf53gJrVAstldrMIsBepqNlN5kLDp7pFE+YSrVf
wtQsBIBp67d3zBMF6ibLM9KNLgTa+sgWUrN/UiQFoHy8p9PzWymPd2ur+mtGDLT1
j4abrDaJXs6GIzXBcDRNAJDEqoIFWTbbT/ji4Jqdr7V8dGq+IKNkJ5qkaxPcAtpI
G0J42Ewf7k4DMdH4HSPmw6S4op8RI/iCmYmz6YW3qsM4iKvLF6cw3dGtaplrEsLh
bQj0+E3ap2en4CMSEe2QBJATbZTd67o+mRr9y379CY1Bc7d0p4udAc1KXm42aUlG
J5MPahdoCqPAb9tblFj94qcusDDgGnroSDMHeVdK/z8CenefvDVmocC11f+AO5iB
7sFXzoxyJr/49tJfDw/SqkvQmxs+kiVcyUvPE035/9mT+2rukGL0C/8eQF47YOOn
zFvwuh5RBWENMxHe6StWTxI5/ysoSbR/I5qX2kHdINS48JbFHQVDBM9LPm5phKEg
ond0qVCXeoJRKFhGvQBRBbZ2824SvwDLWE9oJhfCEDUkG89sMsL4SFxDpBk6wYP1
EwgIi5Kq8rprcGLqDfWCYtYKWFsQGMwBBDDLkmRP16uNzOfS/KdC+K3a10Qg9Jq+
AIxKslMUF3Z2ve4ARe0+YsPAGH81bPX8vVW7XksgrbUnJohAo9Qjmgli86h8X9Yx
vR7T/F0HpgwU61Y7CjvxCRzoI3oO1K+7QmxMmfKPZXI+Mr6W5oxEP8AINGmslrVJ
CHvIgbEiat51Xhnk3/1koKKwdoQKl5/rFMXJX5TLimFcgHP7dSgsJVYE2Qastg47
6gt/VBDqtWH1axgNzNde3fdMKoxDeslaPOytN6EEHWZkTyHudzCs1YcLDbbCGLkw
HW42WcgOo9/OxRhdgjV082QTp9BaVP04SWyK9cqtpZHvylzDjaK1win9abnsb263
4PRrp+Nh9q+KaGTOFWmpZ2B4NORSBWwDi9LkxnupvGJkAz7nWnBfunyk0ewstr3E
4iuVGOlS4i/lftfp013aMVYE5Z+iaiB1TLw4+YqYRxNpB3QbZP4e/ATyzV5hvbrM
iU3UQLl4hSJx5MoYV4fmn8ahPcIR0cr7+n1pYiBRXT98XFl80MxgkjQNEWyDFKcT
U+IGCDFUQ6UxleBnkJw5ZN6j2RfF0YcKepH6QrF9qNWgeSQWMMYyu1oMl6kkBD9S
kNTFWkfFJCna8oSkboNAMY2jhEebH4mqKD+6nCkLT3ijcmmlduPEL+p4iqb4Jk00
FtF0jUWIq3fbM8VpTeP68aZhTdfcaF9lAqYdAnLC0+9hN9kmiGyDW+wr/vL/+ogS
2Guuo5avZqwjPa6e5sAKsJ/WGB7qjtzrTckUykBDPlKtr1+YR5Fa4u1xnZQwZ1Ph
E2EQCmuWue5ppTpvxWNSlLSmygPfHFHzkphenLsVo29ml9zLLzp5+9TJqVWM4NQm
73d4UDZzwtkyEfYDulJ1dUFBmq/mdLYn23u7NdnUA+4hT9g5ByHqNhhkNeattjRu
JikAH5EIpSdns+8p1cFKxC5OlCXpldjyrMzdP99POEfSQV98Q/JsxVewo9AHTOvH
yhjvxnz+jhIRZt1U4IxE2GevrApzjOkIYSg5mRDtEheOZqI6rC4GPEjNgqUSDNGV
rKzn23XJpiaNKaFzPAECm3EHr7B33yQ8RegABc9S3gq5gQvchGZvZyZ1tAfRTXUj
d1e42B5y0OhzUV4+U5RxRkBrxmfU9FUmg93unczggWbW4ieFP/7/TnecvnuFakOp
klAG7DJa+IWB36AClifoaohYu55U6xjUKBWXQkX4IGSn6+AARuoDv3ErkRytg8uv
KriJPY11+5PIgMboq1ihfdpRvmGUOYlQ0B4Z71aEpHxDFByX/C3Y6EWMgHb7pwKa
wQ9cw98j1ajey4NlZ7D23GrfYVnO0kzKqOSN3f5GaZl75/NrOViqJPRVNE2nY76q
ALOvS4z7DSJpqIqisn2i8Ycx+Ai7PgEQuKNjobLFPe4jPljf+UKaltZHC/8ZEmD9
WI4jSYNIellc2qpgzXw5ZZIPnvHTrtBKouv/fTa1UksTLYbboD5KchAQ2kOxAzc0
c2OJwDemGf4cA1CfrW6n+/qYgxq6j2/eQR3wMSsOlXXYw0cpW7M76P/epU/R6nZK
+3JtnHHxXKAJichCRsUXSlS6G2TLAUmxFzU8IfcpfMxq7KiWK9KFOEQo9wdrF7mA
rEvroJ9W/BUSn01wrezPLqMoTVUyfdtP4FgeYXVMOVOfsFON62ZL8BJ6/VOIAPwT
6k+0Sl89N2s0lT6gREf/tH9kLchgicjeVjP1uCK2RY1rXhoCeNG1L+8zBBuU22vu
X7jVisQ1+FnejVrLQZpB2xqVMJCnSqoUWKysWvflB0H0dl4ZkUjfvW4FyTNYeUNg
iFRSo602s2tI0vy7eSUSYGiXoKkzXxMGJg1sdeFNehrTaIjE3kBdodvLTjyihUhg
BpdzCwgXMSXjDcaADO7hlb3z6wUbnG55jUgCNdCJeo0Ao5SMEumZZbYlAnbVP+FL
MafN82jZBT8kls/2d0Uy/hM62PJWOBcJyhN5j8oYpAiivvGmRt8I4eaUMpNTeDfv
5JWyVxP4sa5IYsFXQl6VdJFdlvlBOrGttqMNb2lfXbt9tbPWZy9NeTyJ7GEymtAR
MdnjmZgdIxVA8gOpbqIxyUvVHdFJaZdLHT5px49NwZyZ/oLuOqqPcM893/8CACS3
BidNmHhMvC0ntAugbPQvz28gOctQfFWWqV88x5cOZfaJu7CDTYGkVyIT7AZi9YRU
EhkO5QiYWdsPEM/qFOru/4KF2jqXJZ0AiEDYz2deKF6ZYEpVV+YDQ1XxSXciJf/e
uSvtY/k0p2qWERD3gHItWMT5BX9jnC5LL+D/nspVgHR7gpU72w030Dasf5SWe/+3
z3dC4rltXo8HuXqX/mb8WmI/0oo6w/RaPAsFA0SpD+wQUAI9VSAl9DJMQl99B3/l
hj8nY0oYrVFzp7sNm586XdNf+6cfPiafP9dxKEiwe+1jAYvgdt7n+3bGOcfiAHcr
8wpCXLUPjjaOgiwmQuuHc7oZF80/mYGPNkp/gQIMLJzcyG0VMHiMP54PAaZdSPuJ
t0ayjF4krPogDZGAAgjVx47E2kjqeIxeGE6WB6yRdTxWTZ2XYwbBA6mjk8CP5+us
1aGQWMgwVYiPNMzS0703rZrvMDXifIVAD3J6ghLvOlRRcWnmyp8N+xFwTBk7Q87q
2ZnpuTbMR4jkjo4tB51O6SqgJfJfn/jlWgoO2gTgxbrkPss8gZVzR5zUgnRr/2nU
SSEIMh0maj9XpX8JIMuFIFukUhKsyZoN2mBqnWk97VDK7RQPkeFFlEjbdgLgp7xw
U+DeEE7yeOH8t+YMjIaggWkDgQgwxttqR7lOm+3orn5FaQULjvmJLbU1bOgTzBHj
wCbx+1K1tUm/g9rpvGaaRljCdzG1+VNn0Yd64/JbY95u1fSMTLERzkHF7xNgnDlc
objXVInIpcQwOLXM1Uc6bGyMLHjfjsP7ML38I1WGJBOtnnQsdAHsZsmoUfruTdRl
wFivoAMvA8oV/uznW0hr+keyObKJovWjLqmB9xLlJaISRQLP5A7X5Pn/PENTfaJT
WldYwrUYtVSTWG6PYMc2a32d6AAVQ65XuBC6pm5nDedP0VW8MZt+SvNu5zkJuSEv
PNavM73n1P1OzjUoNZlyqV/hzwFOomSx+CkjBw5IrHw1UNud6b7kn8igKi4ceWUR
55BYNjONRZq3Chjb1aqZSZ0yNzAvtnO4aFdxb/emtIg69/mw+caQXLAMtnA+hbT/
8ubXZntj0pBFAvjFByhfMxSHZuBnIdvhSFCa8LPcCz7XKWODMnJ74DQC8tAxXD2F
zjvkeWP/A/8/yWgbI489ymx43HKZKABGAyWtXLSMnxZwba1uaWwuyUwcQYbDAIDl
00xQygfwxnEOwVKG5QQKfx5qtqiznOR7T0B0gHMEh8kdCQ8/v8qPyciV1ujlHVms
a9GFifznHIfZYWBvBt+J8BYnzcVeR8C2EsU3HieG2xHh/MG5PvSeZFFMDdR5F7hH
hiqr4ndiHwh63AMVLEGj7CDJTqZjtTnPChX7mKBmn9b3tq6J3aKSoUZuLyu3Ixz+
N5wHNGOq52dZfKlyD96JiD+l1VxnPRbtl40gkml7sPZQrJFJnm+R0eI13VtTiVBl
wo5Hjqh09CXP2HkuUk6qEaocfeSDP82qHoAv3ueFjJt6enw+3235IXoFOvfXEjoO
AbjBaz6iJV12aUEYhxZIdYfKT6koQfm+UWx0ZKT3mMxZF7E3097U8VYWHbLpWp0i
kgjzyPFSMwh4gAEr+7en/3go05Eig1RPmCDUUZicyvEDe7ApXgznfAyswFyDIz8F
rYGh0ZQiEaf82BRFo1F0ZEnK2jgcP3QD+EhY2Y8GEl7K0WWtvKtLb52CNPMcFKF4
VelXawYvLvITdTiek6uL4WACX4l+IDnrasOJTNpwm6pBDCq0Xt2XfPT2gebipxo8
BX9imK7sXlLbq40Xl7AnAAgdwxMzQD32qES+H3OS0ilqwnvusy3exwh0I0PvL0VS
1OSI0T2GAWurasAK2+UNrztapA/txNxNCIZpjnKZLdxqFDVyai0XJaAbz+ROkkcj
xJTX8YfVR3PhpYA4a1hoVroz0cLBpDfp8289TIJTV/Y9OUVErfWLwwC84ppcXqtP
DUiolVo0dnslXf1E8snswaw21UbPK5KbUMd3PUBrBvClZMx1/QdJy9phORKH0DNY
QT8drxXkOFUFz/Ji/duV0MRy3JLZC4SKWo0FJ5fHctvt9beyyGFbuIl/XqR+Y/Mf
PNynz1hDCW9PgdhxMOxQ4jyHaysMrLhmL51f5f8xKyYsuOI7vcQJ35qE0ySTT6kv
tj9wzQ7iixzZQXW3RpyO4wDzFKgHyokUgneMYmu5z069qQG8bJi+4QNBSz5i6nT0
0zWSvnCf8hUt1rRYw7n/zJd2x3j98aMwStza46OLb4zKv2B4OO8HlywThz9EQuZZ
+QXeBeOpg6dR6PqQyTBxmsdKZ9NUsCEnmoeMzcohNhBChdEa1LVeu7aIVwohtmM7
4WGI2xZfQvtK5I03QDVlPrRq2nxrm2yD6gs000vfjMPssMUZtcEEuKrO/Nz7+/4n
fDJH3TacK4vsaYPwJnDp4ZJjABX23FldvvMvAGTXPxtoFTvZwMT4a0w3sukJH9an
7tMiNTqKF3kLQb+mDH5TwYUpYN4EX7pcBWB+wavjeJov6YCMiebdeLMyjTt8mCNb
AMSATcqWIE/7l4OwjEua2TUl104mxpUuP8uzXp6sxyi1tRTpY8gRimNQMTHI8cjU
5iF+Fit6vpQeXndZpu3iqYaBnnj2asyYrbEzKFsguBb1ORDSywc4TZGyd2+UMxhV
UuFBvaPZzIayHhjcucR9O/lc73iaJVS9CpLTx2zG4MVTr+7wFcifrydZTd2Z2Uzm
+S+Whh1i+nnQ71GlXD9t7UYVf2rIFfJNU7UhnK7Y1LHx6H7A55BNtZoQ+yHCC6UE
IPr9hGZTKEmohMf49PfgXX661R8E/Qi2WAYFMYaeCB2XXj65m3kac9snLoRUZWYw
bkLvL9+wa25WKppN6lxTU12ax/Xq45Le71RnYwnmpQxcVKZ3KznioXHQW4xkvT+O
PL4H9EoiQckBIu/E9rHhbFlMNI+xoKapeARPA3adbmdk1I1Mp53gZplxQFHFevu0
7+kSoGx7e+683petFpdItHUhnjENmtpw64bdfg4mxEHc59iA1aHdhf6f3bmqUB3u
ZpN5AXktFyototzDBVkn5CU8N5uWLN++a4Misk8xDYrGIQfAUwoW4eXp/mLct5EV
cgm7cDehpSwuRx91CYszoFds8H+0FPoynIB1bTFSqv+wzd0KIVeh+0K4HP3/DgG8
jeZdSx7F09KYsZUzEPun8Ek5SWKm8f8CG4vGnV/VqsyYFxBBO5L8wIWE647d1IaB
npobp7RjjX4ToYTjuRbfHkF7UwvT77qc+KZwpxL9UQESMU7SJgnrFo2H2IHIBSIr
TXRs4gtd92h5owQ3L5S6SFLJ3Bn6wCCnG1w9dxw9k2QTDBC848CqPkWDeQB4VDqR
+WeWs7QT3SG4FiQTKqz3YJTFDbibvBkSCMJ86MvR908vVgUM/QBUWCtsOZbBXC1g
VBSXzGJ0X+7C6Zv13jbHvPnzUqVE9B2KWx48/wN0xENZfI/SAdkOg4zB/m0oNciy
ACSGY3uh4QHpNo/i8qcIp1QOtLNKnIHS6wUn5fBag7u76GJk1PAb7Uq41xvxajBq
KE8SPVzCGtHNOnl+HMJh3nA3l5ABOWx6wqg4l+P6t/N9Ri6Qo+TZlvPyYHMU37Xx
k7XxFiOHJOTRJOF3tjLIn7OHw2UkIpy4YvCYgEfsc5v2Gv8bhpOJrFFYeZ3SQ34N
cDEpw/f8qAGTAJqbdXAwrbK4N9JKM6pd1WX6LVHLIcW1zMdnM67f8H6pQfYChEG9
EnFMsyAiKDajmfeeHCEe5mAFWjXBdvU8yBjQyh7QWH9e18mUqQo47wAdAxfGipyF
5AQvXSlTO7d3GqUUS8XduIGeGFz9sWl5mvWFRnqn7776FJ5dnphK5cZYSmFIOXZh
HIqZYVytvZW5MDgUqYtdaaBKbe+XM6il2LWEqAzPkLpDihGXNsBqzTQQSbuMgOTL
N0MqRcNh+STvOtj8u3RfuCmZDPqsq1g8TO2nzxEdZIoTgOKZJPPjOlI40icJGA0K
5TW0n/U1l9JnttraIdo216dbq5wDrY1xlxFFIbJBmDKq2QS0+6gulVMt4QOtnP87
vTES9m9oH9K425wIJ3mJny/XJblR/xe0BwarOIRYsgA8qDTcxKKWqlpzRIIsVJr+
RTiNBp64nQp7Fx9dc9Lpw7+Q+1+SPI3FURdJBqMqXgf224YxMp3uZvVURxVexFh0
xPcSubwM+/cOVTHTeSjumhZZj94rtt5AUdTqpoDjxc98JfsydsrETpi7oCsjppuV
7rYtAXp3rwl+CucZoIAK1raElXnCR9G1VRDmxZXJO9+2YKpzsH8u1h+P5HGlwReo
z41VSch9Fsb2x0FNDt9RrjmDQ4WYrY29lwd6PgeR1iHMaRTzLPy5swPJm6I30sB8
0/60gK/U7OT8AyCsbvMvDnqbvoPC/8XxnPfrQbJzhjnrmO5VuBtcxVkSgynnc469
aq0ITXZurXEND0Xbpg8bY2wOagAouZ274/I+t36FG/jtTMnZkSSj3mLLPyDlFZoQ
6gFPGRa0DGWdq6CRcQalf6lqEFrKnDRsr/2qcgusZIvJ0rO6v/1xLrYQ0l8nSjdR
9FzNsp1Ctflt4roNc4qMrX0AAhUzY8nKdZxi6cP69eR6g8+XRYhoifPT4jQtv7Eh
lbVGcLYnjvZhLoqsDVQ2+o/bp/qL42HkMK+us5FlvQVYLFiAc1eJ2c766neMYVab
UEhZijhnInCdIo00orMSK4wINRjrqYHzT0AJ6k3wH+D/6us/nGY9B55YBJ/X6LmH
pd9UXo/kcnoyFBD8TPpeKbn+t7rlSJfNXMCghs81P6QYRWQPAv9k0gaOuNPAgZhG
3Bbh5bVJr2tzhL59VFbNSKrGtpQN7KuRWcTmoWjSa07MYrTCV3SSK4odqEE9hW29
Sv2U4Eg/wQ5KXarFJH9432g6kmHlpZDW0/wWqsYhFdnrhK3VLwR9EuuRdzPR3wOZ
5mLeRYyDdt2vw4Lil9NuQ+tRXC4LpPOZMnpAEMQ21PLqAwjFTR/FtjeGEP5gq0iO
hVPKkKSYBxN6FRcQb5sX8yuqAc5DgOcdk+wt/K+6jA9pMIIHfZvjvH2M+8cq/Kwq
c6p+K95U7D8UYZBXa8JtWlArhxvw6dfHHj9Ulv7p7+Xw/QRPfssYDwC4VOHg0ZKR
7ctX9y8NLSxSetUa6wHb4Lia58wggi26TOMMy2tpOwBWe1LDkrXRTdDJi8jlQL5g
pfdMd88JJwmtgnEsi102bn8uLpIyqZOpbyH5Jqkrx6pcsAzLPsQ/W+ecuMY3v0x6
wjZ8WUz1mTiXcGlBEbObg/tiQxEIy4koeZX+WX8LrGoyIJ96kmi7TmpHaqY4cLD8
JxgoTg2MSaLJicWMctmg/M+pDTeogW6lRKQG1Ll1wggVmkQlU6iNHGkQF8FIb9Ft
JpzqFlXa06c/6+nzwWC71CGTNqGp8ZcmU0+5tywXp74uzui9ZPuztfyySSqatksB
DbzG83IXkrV7xYLzOoiXEZbcGjGpZF/yJ3KslcqT4+Gl2Le7aIayYOAMfDwRC7uh
sxcG0RK/nVSyWdh+1041fbJ834iSde0thalGQoTAujRb9dQ53KHutPTxtuBuZg9u
RVnq1PQm3XsEF5DTlzWpVtD8Yfiuecyl03jq9e62HZN0k0TBreDCSpgmrf2OEWKY
ZS1olH4EC1KHgOigHegGmszNLaPZ4El+Jy4LV6L71vAcmdA21m2RJHrwshljSd7b
IZLJ7HuvKGIc7mHG6qFznbcvvbmxfQ0Vdrksefjb3dV6/bs64ACi8g0nKd4Wl4Rv
PwSoKDYQqFkpgrpfX+rVh84NWqIB6CPhyI4O7d9Wh+Rb8ivPWa9OuBilJLFuW+CJ
zphzUXZWLFJ/Iwei68KZESnvTFfHRLcobjSx0txNoVJbKOKxmFXrQlElYB72+Cyv
Eo+bsWWmBCEZ1Z/MKzPFMRlnvO361QmlwYV0f8lEyKSBp21h6kuKf+h6En7C+WI0
WngD/Bhstv1OaBAJ6FgjmB/nccKWmQMz4tH5YSvcuAO5CdZoGz5bSyFGZkysrHUj
Kye/R1CsA1N78TZ3k0z4dvkZV1Vh2OxMRm05mMMC8coAw5XJfXzFAN+AXC1VptWk
sNBTETdrMmVQxRzqL3qi65QC4pJvGuOkpxBQJheF/JdZ4hoQoJfJg64ZmUiUAgh2
KH6r93PWX2JrtG1tPFpeAOjhGT6eI9MRULoQu/qG2GdDxAdH94YO0BSl2FZSvzme
P2tRWwqKqMnIy4UIbGQYbgI2elvJ1ivMST+/hFb5HbaZaEH0+HAIbhSV7gIeXfkH
ynotjNpcvLasrgNojBkZwtK6XkdeKIllNdDZbsRttPcRQomWenrHdvv3MdZcGPSI
o5uS/sJBuGH5Pw1QrwlYZpIsgyWwA/hKfU7Y5f0iN/Rr+bL8u5JZz294sF7OvgzK
vSVj+UNaGRZ8GInOdHomCnuBcWJaWh13uB5V4EqBB6kgv5FNgowTvrjdH5L+RYuB
MKs0mT8m+T/6IOq0xAwM/MJRrEGiHdXUvn4cGXYYfOocXD+5o2/5gkLDl+5qubnN
ugPBF+7iYSSNuZ1Qd2F1xNG2mDZ6qXxziQl2+fJ8EWHhmV5sN95tRi3/OUQ7aR+T
rF5OPO3w6uf8QbmenEPXlIs1eJrBozjJwHadx+lf8P5OaNmp4O5lb6Lrv2f1I7w6
tyFRvec6+1pEL8sURr8a2APC1x4flN9Un3FxnYf6Q1oCY1ONNB8JEBKtK8nC7f0N
bKP+xvGXjcliTY2Ecq8RXW6yWkjoNbBDGvv+EEUQQhLjVX87VBCe7uDbUVAzcicc
GMtFUNODZ3I1ijvRkiRfgxnW5K5kpVjs/vrgoVJka/iQOYMK1uVx+hx+Xr+Yc0hZ
8pVVIdeY64CQDy0jOj4ge/0WUGYYyWn56tGZCct4EHxH+L99658hFFhYJ2ieJcm2
k6Xocyn7L5ndQuuN8Hv5iILHudM/BXmO5ndsnDUinVMq1uBPZoPzoc02R09urh+u
mf9rtOQGh2UuABqnkkenemtZwlXVm8A2K/tnzI0AqCrOw8cgMbJOwhSvug/OWT3W
/jmVfWXKvKod2jDSu6eouiH1t/v5eSzZVE+lUKCPOBzyV+X/wgJrYpnbQcD9i2xL
W9Ilzcj068WMYIrcsl8+lvGnrphTCTk6Kehe5wh7wCgV50YXPw/qa6xB5LaSLYDz
Trbe9a2HgZhst1ph6ykuwiIj/0Tq6xyqKiQq7vqI6jv1xcyZgdqFUBAnfpEEJRnb
QFsjQQ0KXokW5/iOUc4DUepnk0M7P1XVe3g4IvkLyPwyIzBLsq+L1bi8C1UvnFfw
P49RytjUkd5zIBmyOH8YTcsMponT0pHSFSBUvEqORkHIyyzXKtsocvl0GGgjH/f9
bWIHyFRgVJIWoKysuyZnZ7SdAf2id/dTSkW/yE6DS0TVJXQ8vZtDMP7afOPZ21Gi
kbo3tKAwMqUsCgvk+IM3Yee3AlikqqhOmrpGwSjps/xhmNn75oPRT2evAANVrZEP
rSwLvtVTDsdqdarGfZXet4anmV9cfXja9+F4oQdXUQLsSQSgo3VvtzW2uEmGMnWH
lsUJH5tnV/uNfMi6ZQUfqm3vSIkX5TLqpIPA50jGZod5apjLreEoJnSikz4ocFA4
BXzxiz7Ux6Hz7ZWmPNjDOKHIwb8nr/tITBdNLc+5IZ2RcSzVvX2nYzHN5vm3TMrp
/g2dztcFXNTeaj3H9ibhJmmq4LVbhL9vGp4xQUIe1dPdQ/Wq0KEjnBuRqPfI8tjE
HcQUAE4uHqWGx20lacWxfg99ntSQYtLK4OxkKroyc79nNT2A/qMOmdbcd8nTrVxH
ghvp6NGPyZUF4BZMemhefangze01oUGZhuxic/PD9zjXZLMUjYLWhkjYLelY+8vN
mnvilyOJMcvlOftHzq5eLI6ssEQ4iqG6SBT+wMHex7doTRj7gbLqY2i5IXp/DXp2
lvJFokNvUYVQ1uQL1i2d7Bw2QlnXgGQBZqTZ3Tme+aRyE4gKpP+3cxo9QfbSWSg7
omhdEi0iZQ7elL3pGxOJKtAyxJJfnNyYf+gkZONO7dzyXec6lgos8UnUfp5ztgA7
AhNam9Bw2mOui6O0FZWPyXx4FVYcR3S9KHxJ+HcesSgWM9AhbZGejMLDsJLXlvzw
YIvhBGOpvPi/GiO7NRZlyosY94I/qDU1nJR4p0HssRRFlWhvtRI9XLSgpU0LD+1i
v8ywkD2ipDIMoezMU1YBNz8D6ppYtVICNcCyHLBYh+KXdOKW0HWJk9HqM8g80SIn
6fB81C2RpmUveGsCS/eZpLHBgfTx/trooL/kzDEP5fNHkw1GopxQg/hIl8TLfg4N
oCbhyC4Bd512niLaQro4NzS56aO53viMm1Ayec7RwHPOvZ7ND39rqlwGrsMmHF8A
y30/Y68T3aJkoRrR6YZvvV5U0pfCtZgSZ3/L6T2UZBGBLBdnSRxqNyKMAOc4MRYD
DAEEfdGY1rGxlqjhhbVnlurWUQbqQNeAjV1N7DRCks3CNyQ+GK3FeuxvZ4t23m06
dHFX7m2hARiFyrmoYFys1unBCmb+X6Vx2f0wDnZYakQ8BLSVtkU6ZYJi2txYIkST
jOTRDWhcOyuKOWqmpmfIutaS1p8s8v/MBFMAnlxXyje+CAPWHiKnIcwvQvaecVpD
7sZQO7E6cHe+5yu6AwfIGkZJSrLTr0UgsEu0hUIselPT5pLrV5lpNcaQzThWy/dK
GgHiKvhQYcMWuiNlLupJhVt8CJ048vvOeOTKQTXviAbawkQb0G7EWpypMog0Cmvt
fMizlioPHcjHqXlYmUlj8msIGFCpsTZcyT8730QXos1c55WqLyHoqrreEIsqZNxx
RoIzIhH0IH9heq7D+ZwC1u3jmWXT5b0HLzueqPsTwEqm2crDU5TdWj0OiDyY61pJ
d9oL8Pu73v5rcmu5eWLjLU6s4WQnBLgWiCZCC6x7reqUU38DPaQLiKHySWovamyg
TlWLNbaI5V0IyZMjiz3lL7Z1RdPsIywe8nMlrApajBXWzVnP8I5T8Kx4K10ONQIc
TiAtDSWmkErlV//HsJ3ob+TxNWDjOR4gpscyUK0ziCJ1FkZeg7KRNnEGedaIAew1
xyWuPle6Xjda+3oYIZqdr8arobsQGBLuohZu7mM8exhRNRcbCn2lKCmZQJmyrMzJ
3xYgYZtdProRzDmX1UOZE+Gup9W87FaTnFXJHhAiIhJBTJNP9jNgPBUM+TLnnwtJ
uHX+PX1fE3WtjDE2rEK+3/RXWTNvzovlXKkxQK0WuxVTL1pVqP+oB/HO2s1iitk0
VPwdDMBfq92pe52enf5QQxbRjUiqQwkaBJx+1D3AAoCVP3EXWNXS5fOFxWB++J3g
nYwVGSWwQ5s2Nu5dt2Wtqh2jCOF8js+VrhkK8/G6CE68GnQ9QvfJQlqgi3DrEyVv
lNrflE7mz6foSGlv3wy8UTFCjpZ3zQ+RpImhypY7/CfD1xChDA1l2l7vJchBdRH+
UmnodGrZ3MHyrAVSN6WoKvig9JzFwoPtrQOL6zEvl/8SkiRGCK/UTvl97gnCS7fb
dyHl6pcMxuZ8hUHr0EVit7324v9r+X2Hyj7F8uXZXGm335D/HWv6V8FCc7YYdbwu
bvu/19yJIZ9nAdsHPX+fUNxpGCV4rhEZg0bVgs9WT3jzUei1F13LpPCS1LON9AGh
ogHlonCaTkKaU911TyocWrF1nJnSs5yNZnN9JT5DsByTOqtNlaFE6LY00b8DH5aq
qX324ncOJQWP0zLHoHh95JUi79Y0ghQ8/jy+Sf1T+I2wLWotgxMsHjknCBrnA72a
Oz8Q01SmP6D1oBzlBvAm0qtvT0qxOgG373GMp5dOa+g0zo5XUyxN4CSeK85E3CZo
PjnvJn/JztPlCZpMDVgFnIiD5G/KIv31QJ50NX5qqKI14i0hhh5ElnF9NFsj0wRh
Xdi8a9kKDesmCcuhnweojSIQ6v8FW3V8MiWYCynhcMW1+0ac0jybtVVjyl0aqd6G
DR7fCojxlelY5vrPK3GERMcaUZhUXRYy4b+uImZz/F9XtjoOmp+E8gAouU1k225x
rwLTDy3ZxFfzHDHGga634iYuxSf3GJIODkLZTZsJRnrSB7R9DqERjvrUpdfHRUWb
5vPI3aHGj4Q+ejhGOjtQdJ7oGXG1mIVCK8WDeg4ucGcVdnCpay/9G5R8gQ5A3sYw
TPo1b4hwZSYiuV7445oINmjRqcbnS9oSwxyOxTU9WoedNxqfPyoJEK2mPQxbqCYm
Nf+PDvP1VOhn1wPgob0xnt+4Tsjzucr9P9ensd4CbmRrgBEhzOYOL6KVinEB74hu
H8C6/mYPU75xUEpXVGezygKvl1EsOxmpX9FI0o9LoMIYUZyh4/epozpGToHscTeM
1bYXPW2M4EY+AKnRN4dVjrvM4h2ROyfYJ6difumI/3oKVJ3+XTPsCI7NNE0iU3tY
a9y8uLp6/MPoWIMDni3tc+7VY5zGbUZVSOLjpON0b0hgcq44IbrIhgM3QnskeSBd
shS7GPgjeIvC2tIYSU5WX/qeGFuLxuqKV/k+nffSV3UdyPTD23O0UqxYFG46d/Yi
X5AL3VI1stZ2E9GxDQT9cNtP3O3UAa0ahekyiHMX4YnZNc2q1C9MpzuYZQHbF8MB
2/c/iau4b9WvuSEWG7GSRzCQxBoPvCXvmBXabuwO81ih7yB9axRSiNMzEcfBBZQm
O4Oxaf4kVNSSKb6+vCS3KEw77extPN2foR8VnygfITftJ+mkBgD4r/L44cdEYRi7
V+Lcf+2BvqgT/sTEOYG5TdQtIXXMc17bGgViOCRQE3Rd52cOm5aa70kdX5+mPnQQ
0njVePRZFXzWK5U5tzcpIrjrdOTQgtADJbQZg4f6dxb1RJCTXfGjnPYrpWEjfOcw
sIXLBc2a87l/9gKF4wM+49AGVKpvvxw+7kKK58ySi6Yn4KjNXW31EY1gFVAf6Kss
4EBeJG0B3TcEuIohOd5T9LCqR98HEcF6qID0SCHG97Eoajm8gzzai7wZzsF2LBvY
w3XUhfnx4MBMyBvxDm4iCHebgmeuOTQZVTIsk7NjTT7vOkezLLk9awXpo45ikDl4
8STdrrhdHc3gFGhH7YBBYfh98VaGU+mMDZPPNY22cidZyE8x17vvR63G/jp9TOyQ
G+So7EPgNLor1VtXpaOPZuayoM8cCgUxekzfiRmHV4M0IUdMmuio32H24l3Ne133
YMxnO0kZRl2nijo37gYC5eRlA7BQP+jkO0janb5xTMQLZXbRfbFKzxg2VsGI8nJ9
NSOVC59djNym8c8R1JKwqlpEgnf8NpHVJ9NVrGCzD2ROQ0Ta6zZdNe0qufT0nnQd
hEFtdTHmsb9S/I/xqP1AS+JCPuAM18JkK4PQTna81hFfu5cuc1zjPbkD3u2joYaI
jMZ7Hivav8UY2xyyTyJvZPbZMvs0kO6rwYwtpRipNskLH+nWG3sTKAjRofKE4jk/
qcLzvuV6r9NQQzRpMACgGFO7MMx+6H0F5+WBv7fD8DJ0W5/n6jhPHsCHjn5+eF2g
3OG6PIzP4VoJhs2PNHmUP3PqKZY1WCgEDzIHzyz+bZejPoVMFXAuWlV0Cz4rv61D
1e63nH1mo6H8NadERcvoglW4C7Yb6hB4v0XvGhHyFgTjs7YN2mpPovqpjW3PM4F2
/CE4e+xuhZ0RuyUt5K6cak15RvZ1roRglC1QKvp6Sor0Hh/2892DxxztUYz/gDxz
BFc06bqQC3lLlMcDYoEoFCURpJ89CBO+gjohrAPmTVmOcJeAvJXH4UyOcM9Of1fE
uzRj6KxZ8S2wEyB7v6mi4OSvWY1gFsND91obH6RaDiaYj/Op3ljLss+LNAYQEzQH
XtbZqr1QpN2tndealjZq0Z90/3JSThy+cYP4yXSuM90arEh9eMPcBhTYCNTySxf/
dEKxWCHhEFUg32QHIBeJvifoyE1O8cbUAuwSoI2TF2bEPiLT6sXqqarMs30SKI9O
am2z5siOHF9d+Pwgrj9HOAOWEF88xObuU7SrfXjA5ZA0ZzyTCMOv0aqG7fr2PV0a
UVfOmBvk8vlLjo3f/lAK7w2EBgvmeMpvD6s/Ljslyu5tSm9BHBD4viNPNuI/DC3X
wq/2xapyFYTN2ZbkBnt793wRnWXPt+t8Hpss4115dr31D5wM203TYIrvB6ZWn1RA
wsSUAdV5620tzUSRvyaqe5epbMjAQjVbGExdItTpJHc1/7DrUj+5/2MaCIXcComj
Jxfi3qWJA5xNaJQXQb8ZVS/lWWG8zP+D+Gj0K8k7LwKDaZPExDtpc2n4OdK5nICz
/tdOmnKEei+VN+nq8CYkk2zdWKy2CEJvQjqEdOQqw3VDD7eQpI2xn3G01OFYNaDS
rpes5ZDRnCjZl9mCyWazz7O0lqYx8V8mpDkQAPTPZUYMpWcEVhuIWZ1boAMF5eZ8
UrpQDTupAx1XBpARcFyv5rX2NFrzLlE1zCJPhivPUman+ZK0FtKcQdCGQ9/2+lTc
4r5FJHF+jjLHd9p/N6Co+ZR3fpTSwAGTrToWavKIOVnQcSdtL/7el67Yboc2HlYH
UhDL0t4y79+3AEtiT2/l8XMhEACOgD/+E6G9aBLa5BDsA3//tEytRo46cR+5JT2h
lQRwJ/sFLtH+PcP8O4lV3G9Z6VBCriJJ1QvAKi8iJUK6qlxxAc44ewcM4XzOJCcn
1y1YT3f7/kb2K1CKw8279rbo/qUuYsO+Dr7UVTYX2DPLJMMGl0K3HDLVVx/swdRe
WKDTpwKQyC5go1nbSl1vkbXEjC3RTTMcdSPEre4t9Izha4juZwU+RVwCrYPQmxo3
x5ZkIbFVmkUTB5FG8vxtgwSEDGGHjE7mEvMWYAN3eRXLJQUT5yq9XrEpJ5s2Zc57
vVgQ7dy0sAaDuQWED/gDBTOViLnppA8nzcfINRGtsfqliap5QczXRXuFRK1Zuk3h
GXvJjCy2Dnn/aRINdfj+oKIWBu45wCeGmzgB11edjFmq3kFp6S+PIY4Trbi4pcCt
JhZ5ZZCpeh84rt8/I4igO19yWG7MxbZupySjb+28CyqqF4SBegqNVo+1UGIoViws
xTXP3nJuayo26aV61Dur66n2euK/tDPpgZwm5FP0tRGyRJvU1wD6oJde8tc3rZ79
GLwkcCU//kKOB7ZaXoXvhmcCHq+Ukhoq/1xcq+gRojiWay9D6+Kf4BtRwX7KQzTI
z8qrY8kQsD83BydgOnxNYgMa8PhvtmXAYBLsdWKr28hAQjC8m9yNf0ssQXn6mQvb
ROJ001nIXBVB0AV6HuCho2+z+addvIFkQJTkLRXeDpNrBAuj1yPxejLtJWWBP27a
5cTuOYgbAHAr1DEzyo7xjpI6jTYyuMH18zwcIWgH/r6CjOrqO0i5qumk9MfRTgyQ
BUwbX30s5Ehregc2lpU7KZij4gHJUp9P3e6lmvQRD5w9X8OikGzZ51M/I88NjQy+
jRJw5kDzbd1kAtem/SiY9UxjPFDGLmjOTlNqieyyGP7aDqa6tl8TewHPGqHCFFHB
UAEU9LmeOt07sib341Fh0PPgde+DRMdl4zJN6JMi4dTimlZF4nhqwFATKr7zCIyP
cL65dP8vSD8wuzsaVLJeURvel6doz0pSn1WG+jC+8TrqcgypHS3f9dDYmva9qtkA
nioWXP00Jm1x3YAyucS67omIob0mJ3R5gwZhj1d6ZW+x389FMI6huMs3ougKdqEU
27Z6Kve5WzQBCRDXU+g/rmjQDjiVs84qrytVKokCFreoaJH/hExjqv5OCT9toYel
0XQ3P+5CsSTtSF/7urJhtvj8psPQIuxjUhBk6lPDFUfjfFEKor+lIMNHL5SrYphv
iZvteteo+SR+ZdtUFR4EHvCDwGid63qSxd89xKWuta3BPht1/Mv7eZSYrbn3LA+R
iYb0OpojePZynSUJ4D01RFwVtvfs/hNKkBV5cJmqpBJspI7U1JxaK7LPv1o1gPSd
wWGZy9Asn/G/BSZBEj7WvfmxBIs5qhPybBkVJBThuXYEQwIiHAybEYdgCOsPSnYT
4qg9WNqNg/RMEtHNknQ+7dcEiC73F++4gY31LmqXsK8qV15mB4b0ovGlSpzGUCQ6
bbX6ZhP0PNrfRH8kVQQelNyhgpeggzyPU1pHIPawxW30sEpLjT1xaR7KhMR3jqSC
N3472ifPTmtWRY8sWY081snWg64IFVa+SmV3j0/7w/ryVIjV1mlZG/GcXguxq6ju
n36QBamYlDssg+9ds0W91D/yIa6bgZtGNn2jjids2hys50xfcI0J4fBVgCnijgcp
dpyfCy5NYbFKFdLknHJjZ2VL54TRhZ7S9hfIZOfjv+IXa1m2KNtEWS/HsK6NdE3u
Lk7omLjIetV70C4LFhZozAkWYOjLtpL3A1KomWMox2A7abzbGIlnbYfpiATYr+zR
RoNPFxwmO1Fey8h3ukxc3wEO07UwImQmqOt80RjkuN6Fs0vxUsK7+Mc47Kq86Wem
pBDrN07gqH9vgFuVfMzQDKxaBSknh64lT+Mom5V0LBHGWfmnr8EePwwAQPJNEby/
Etk5fbhRnonVQweFEnqqFStiUlX6Q/sQDdhS/S//tC1RELcZ/iZUWIL8ayinAeqy
/4ZyZza5Imt0pcL5PxHF1lP6KBcZgYspyfDYkcuqdl3CbcegKXoJezsHK9Z0hdyI
/WeI3ISSapWsJQFPVWhbgwDzekc+iDvpjN3IEwFWz0w/s9oCOPcqBWT+Vo+Uv2dC
4YwXAmsV9BV32qnfOxT9tUOBwGqCBhNqQ/QLza6Rcpyemj6rawXzBrk4W8uk30TU
91UrMgIAhpYa2JL5LjluuBbjjfi9tj2gEFPjoq/hXlB2TcE9mDujYEqV9QsK4ts/
kI8+HvkniEhD5hjUJWhSgWf9SsgAH0qDkQg8RMYq46TFQcWcl1S22n+TneYecIzH
D8mGixHI9TSVCmtR8JpACyX8YL5K06AH+agL4WG9uCFcdYrnhka9eem9mMoYyaVa
DnUuV8NDV8ZN4zKa4h/wAt9x1AWkyY+rP6M0tnR2nseH88JOmsLbB103wMPlgPB5
3ORRor1tO0SJUA0FQNaneyGGpkej6cogiH50Q4pXUmpL5mwBrdL69OQ8+ntLiOKA
YmATpvi+kF8EdWz/BVY4BbKxDppdMttK3oWclCDOmde61MwNZr3MKoCCBZu+X5f5
mZncp/B58AtISkvVPO1mcnwieBQqDPQxOAhoRHFuAMMs2balV6f3U34oTFOMTNim
MRNbpV0jeBE1rZzB22DEA3SRzWmVEaalfaxUbMYWERmrnCPNmA0pmUT+gANB8fW2
QMylLngFqk97ZOjxIcYJx5kNVlHoHg//KrsycxmdTgq8ME0NjRX2thlu4juvewNv
ozrJ3L3rFAxHxixWCEab4hPZB0R1oRhuObWbpMFYYfhVxpfXtuIzOXkfVWMZXLuS
Z2VzCYMSTkb4Zt/2pWIQ21hlStXnbB8JSJ/dCVn3WYO5lduzTVZ3t1uMgX7CfS0Z
FXId71KFiXhmZwkSfsllTNcHzd/0Ta1q+EYMUfHPJNG+ETCQAkHQujBqYkl4j9Iv
6UDN9tEXIMOlZKoqklNVAbkb8vZIZs3NCoXVnPyg3tXTWwO6dSDdHKHbAGgasQ+c
mI594kSCCIBaWfVJRwNUJ5HgOVspoXODmXHguMBnnx0QdGSEyaFXAyPHNpA+VXF7
baPams1plKMR1GWdAL0RXBMZuA6Z1F05VK1Uij0UAcO20ZgmmspG52ZNvUwD3jM3
jQwZnhgOR48I4T8YBwfhNM504QakYP6lh7QWjrq0lnUiFsxHBjQAl3lyvLYbST+V
9/QGvVWh/AIL8sXdqVZPn5IVuJ0MQtnbBBs62nBfUK7EwZDtrc2EoR2zNnX1v2oP
961aEwg/0p97nZsS/PLAIWz39GcYs0MOC+9NC/onnDRS6exB4Ivu6KVH8FqrY3L3
iLnLJzcOiivwKo6amHfRXhrdTue8mMWU5qX/2P1T6lvLKA/YeUWX1zKssxOhVLCq
CtFSFr9MoCB+mYeL9fL9JYDggmqwLgsyHiP0hC67mBm8woTDxQL68Qc+G7cmngv0
EWaSq7ufHvdmN5QB/CVukR6yTCjkLeQxX9TovrndcVFGksmzmIuDm2jkEnLr+2S6
ls1HfwO6XxbxcGSgRvE1PZd5VyjZvbC4E9nDJTn6vEdrYOL+WqvYFAVA/jFp1W2Y
MONh4reYkYeFQ8N6psnJjbZ1NDY4gEbPU9YvyXUI2ZDKe7aQ/x/CGnO4qKzsOf/g
7Gi7ysT0+VooLUL/ewrRDwtPP8tiMQblFKZgO95VTwbGmSdDh8n8ti0uGsBuoly0
4q87OQ/9C7q6pDG+VW6KU5t7MQj/aqB/fqQqd3gZxE2NZ2XrEVzicWSgoF2FGP8V
zjZ0c2WTsLNj7Za3K/Inib+u4LdLfyNq3+58q+FUuag35SAG3leF8HKF0WGA1dmn
tTCTcsE8pbvM/cmozolyrO4KRnR5DsTyEmSEt/aG84obek6Dsibfwz+QVO4UcS7c
QpbCfO0SbRaLBPUocVrOUdL1mw8mc2/6q8jIyY9NFkOT2p8KaQ0ZH4Rh7ATBU7pa
4A7Ic+OYm/OVY20ucs3PHa0XZxRJVFYIMx5ZDKmnSQsF1FjP76g3P0I26xmncswT
iySmj8FWwnlOOsT6QwiuTwDEv8p6HFgBN6PzUHkjjeeyzCyQJ2rqsKnRs0oWHe6r
Q1nB3qULdEVEchtDGt1fW8UKXlrah/gAKgRLTqDAgeCzbAv0jWRug+UGHxzJqi6G
VYhH+cBEQjlOqUxIHYuj2CnClHQ7W2zkCeumXPJefQ+tgKCYNG7eVuSHg4ANr0jF
R8PPJKSakSZFvn9nYKlhiownf3+wqCJSC+9Ooa+L27ipYPdyMUY7kZgZhO2ZFta4
pC0gK/Y2+enyJ7QzAiCpjZuoFJt0QPj6OC1NNMqg493Ubj4qkgZrPOmjLSHSdI61
3VvQNeRqbhJdl0+h/jq5BwndZ9t63lOQ/B5Z0nqMemjw68LYigGykzKFgExeqMqH
lUFb6PV6x4w7NPJEprma+LH4w9PL5mBF/RVbTTYCFTRaqkqRGdp311BoHzb8sPxw
EfPqCeJnPHZCjITpbRCY99ND4hXByNhpzS77FVyqx43F+Rs7lHLUG5YI003SapcZ
yCBIWhBFoBOqj71wbcjeZyV7JRjyldDXTMPI1uV0bWlQjIgxEv+4cbY8da3OTNzi
DJN9/Cl9t41eVEIRNmKUHgZBoILPL4ImtVPvwHHlvigY8yozXfxsq1TfxcAwlSUr
05Ybw/S/dq6ku41PMG58h6fEhOEVZXxA+Zaek+Pt5LVU1GvXt6/AbHhYPpcLGxe/
WzzGc7spw40ppzPftKWujrw0qKP0AThpjr+4iInvS+59knOq771P4B8ZUmUH0bo6
FZGp3Zhq/1Eo9EMNzAifRnif1lyvcS0dOuxB8c0Z4ET/lf103heeFSPej4xlzpWo
ugmF1aSJQlO0BRUYAMj+dKZ9WVdeHjvMzH4x8bxhaOtoABulT09L9lcYBeSHBVrX
YI/Gh0dZB6p0RaWTLteiID9Jp40qwMel6Rno1bsl3iNiqdVX30MTCxdn5naDiwj9
PzCergwFkvxcAfIkrYQAfNhHjL/iViGxVgYT37MYyoGMWQiQsgtDJFcpuab2iQM5
t59NktpzZwRr6uNb0qJfP72ecP/mnpCtcnIE6LGTBmeWKVJoA770YbBigxE9Xxdu
aGPWhKPa2AeewvCucLjzFTxdkGG5aUeerJpYZQAE8KOpgU2MPeizKIRLUz9/y/hX
C5Y/DbHySWnIZYqu4BoEboM1MGios77NqMg8SU8SnW2p0ZPwUeyEP1ppxTIqMNoZ
O3bgtub+7FX9FZKqPA5SSC5gf+tIWdFD2WRRfRgfuQeNazDLrczFpkTOJFSsH314
NRrH40qWK9xoHWD+YHY9ANpidsG3YzmB76VWpbkslifa/vfWK/Fhn598FGsysouN
5hditenr0oLzU02yzQvPkH30o9sKvAjE8+oHyok7EMly86L+T5ZOd0rURlkNHSyt
854zPxbedn4oZ7xfnLp3fRLLqs5QpedJ1WCshx3mBylYUd3XhNmoUBwM+Cc0Y1uB
YcO3lSA/fqAw2IUHjOfVkRinWfjnX7T3lyfwnkHyYGG5X+zGPSfQXnPl3s6CtUL3
fsQatcZT1KLRdxmJirrvLlZtic4KELjhY+4/vhEr/OUaMWt17rCwJBFREA/38wb4
4BjwA3eoDX56Ro5w5DBkAmHsFCBS0xnf3jZRsDzbbrrydx5Ip94K+B99uF9gt8Nd
dJQIK8InPHUbcOAMzlnl55gXcDgrYU7ArM301Bq3fTppyyMb913btDmpZ3mvLT32
s8kga/wu6oUP2SDqzQogJevLThQY4ZKd5pevQJkKKlzXWhiMKLEVRt/rchF/OMhT
QGE//u9Wt+V+968X0w6EZfZxLn6tyS1sH9C49VIvZSYy8WaunF/FNcRcMEy99KcH
OaGim1iAHSTHW4d9uVEIQWvibv4L5zgHtr374ve5uhU69niD8aR9OPh+XcUTvE5s
dEXPK4ubZZ5b3COEXsB10lMAxUg32QATd0NlRIjoMoyj/pyFyeRL1+Qi3QlL085+
mYMW1SNmJdxehRLSBeC7UaHKCUeNfUjYamEqSsli0HhFC3ubn/5YntUHSkB4o7Td
I2PdQY9kBe2NTRysCrYaRVQBkNieQcvaJIXQcrvy2Cj1JS+BHH7GrMBbhrFZ4oVB
/wpFQcPXTAXTouoN4HF4G8UY+xawgKZM4M0WGp4yYn0Ucoc1psTlFlTFVo1db4lm
qbT+e0y83zXhNHeprJ5g5MZD1/QBiJxOZ61h1bnLYOSdPuE9ihr7hECSvXWN3xuI
tDz+GudMV/VijeFwuGeD6SMX1f8zvualU5SPTrwJ36op8PT/Eh2b5Q+UPeUm2xZr
K1zDz/7x7lEaL97welXPuKyGtxqrz+UssuCcsWBuzrAbsfT10RBtLoLwp9oZX4Oh
a5yGC/7hNAf3VZ8VmuuH1G8+lwniXBuzJa6Z4zFnJEjptZXIMwR4RWbGKW0uBd6p
8nT+CMIgMYgkHaSvjkAKZ4yS4SynZQ6lJ7A6V/zK8nztMHxoLztduf1ZHo6SpZIH
dKN+eQQ3Lyp5VLMincuENgmMDlg7RN4WXBVEaQFRUmLJEduLUi3FzpdiW9qzY8Fd
mIPxOsJGlQNmxWtsxR3Iq9Iz72m0HaF7vHp1IK/JRhbPVQw3Cs7LPlAfPdJH299B
4uPvUfq+kX3Qok/SmBqsiQBiSDXgGUKbZawxiGEP3BwoKQJuQYqiuTE/QPVSCIYb
hLDnTNtuzgQNfXwt5OxUKOYVqIW2f94stvfCq3w11Ta1I1D5GxTIP2AmcG1Q4z2i
j5TM4m4HVwg006w7JQUYhWbNHPka2v6fEgk7Qd7BW1PgseI7McuGpb6IVUQ5bId3
a8QJ4ivDuRR7mwyuYMlkwLqHXtEqMLUCbLOHcI/29mfqkWcnHoIgsVINAHPxfiJ5
XdkzIRidMds1xVqxRyh6qk0qMUt7BZv3q40eauur2+xejj6wKQJ78NrbgXQ6Mgwg
8laheWHlhRRvrnexf2eZhTzBDXHS2bDmrOaODRR4GX0PQrJ6OiyG04swEXdJFfWu
z1pE1oFpDcpPh51dThOGOzJnPiHHLuTxUp1aDtDt1R00flzNwn+9KzVdBghTozEF
WurRymMa16UEIlbJcCjUoEjc9oJhno8HV3NV0yGWBhHk8+5Cg1UDxtLSz7/8T8G+
LJzGt9tKAUvuDRz2qC6fnhO5kLQaISllYu2rsCzzGsaw7D/cPue7vZxOyEA34kgH
5yOod8uPFZSrmqRJYnnP0BvoldRwkR3FfezsKPkMUa9uQkTUVZx0kGWg4tstQySj
vLEq2TsoBeVDYXY5BfjNsFYoSHIAuscHq7eM1ISdN6jZ4x3ZQ0CSdGC4sHwKf1Hd
PfUz/RbDFr0mnuEgbRDwMz7h6BD8q+I9OJbNa59EuNRNO2ZVmASCOzziymUwbf8x
jECenv/NnDDj/icnPgVpTsFCVeModZFu4dcrCgzzvH0ThRYtUBQ/zcoqKXkdhiGl
gxEHbtVMgQ8pxFP7ApAWOI8jkfxxl+FlxdCEhQJeOb8+kV/d/ijlauIOYjVKzt5S
+A+7Nr51KSw4/Y4GJqfX+QAjgOA2vx0ucPfKJgrr4iVELa6wlZMISih5DCgdPHeV
S/tjXqKyJ8xoPlNxj9934vX2fqVhlggBGcFZUY4xpWK6ag5bYYsQShwQDFQmitKW
B2aKgUKIxWlocYpIPl9Pq00/bwSfTE69DidJ1E3DmC8n0DvQwSqUQE4JtHrmxoGw
tasi2yBXDqbgMkJjP7eih8/QdXKon3Lv3iB5G4IrcKgHXhAd/4Fzlqa8f7IJH4AP
MUOurnIaT0QprjCy6Vau+FWDC7o95K+ikkKcxJhrU0XzG8/pzTZEL2g1D4mfYW9L
nVZtFmN+Y5vFtcawTqazXr/bHSt6Xp0HbLxZrykcV05RW7wI1UxvqmDHu95w2THl
RIuuGsbq+OMKQfV9Mmw/3oPQeRwAHaG8FapT2ayYjLSkECaEMUp8n4nyo2te8ENZ
dwO3X5txiDhafwF4puM6nZiEewoB8wgwb7Sw8mXlkTqgS6V7YQyetVcKkan+2YQ2
4yOT30ky+vKJ9ELOs72lSkUltAyMIDlAqBLYTLuC0o+8nJfdZ6c2BpD48DKL1zqG
Vwk/zn3OqoBeVUmWg5AnmLKJc2aXv8HmtdDmd+3Km/jVGuTg/ERbef6WoRikSn+P
9NNSnKwWbVvnzuUbxIDLlNv56b9lVX9mj2xqz3MoA9IlQxQxl9jxA8aDJJwgFZOq
3izcQANrz5KDKgzAJKvF++vPR0wuVK/zKZa16ZZlZ4Sbd4BRS3Q7/ch66hLiMjK9
RB3CIqIN4Egmoughb5xikXhIwdQvR81EwcIiLK56DrKp0GnjS4YNOECwRn9FKya7
jcf/MtVksGyVKFrAYqvDZhCzAepoSRhsJhaZRuKNClIqrNWYvhiuRV02ovuf2F/8
S/kb1mYKMT5PfKFKVO2dAjV3qUA4Q9YPWWwiFXyCakV+c6UjzMTbo8cnEmdcB8je
iKIA08g8MNh4QzN4k8Vp9qXqLncrLxyxahS3XxnjwKY4x+Y2CASI7i/sNj3USvU4
vcmyxYybhBN3+IlWlqdMAYUTZCzWq0/tecS8pntKom4SpIPzWnkw+MPrvAm+8Q/+
ZfOpX/4s8iuNCLhI8mlQ7rTkaJ8gOmqY8YzXB2ZXYziwwMPhxbtXpmxOgKcSvfRJ
uBqh/mTcm8+Wz7xz2NJOWRzVsTZ73deSbGaFOMwyCuHgKgsJN2flp/W2C1S3ZKHD
ZsUkXOcinRqJ8iNE79TxVOb62YVu/qxbgJFNXDHk7bcrnIIDQWG/Q6JUftqA3tB9
N67Ck+mUV2jl5VWl8+exVhX49r1r77klvncsghWz8nFnFJG0yv0VTRqPL7KBOmdz
FyP9NIxCPTjk97RrKkrz4IZ+vW5lncMpuyB4fUUgheH77n/rOWUUxOHnK6tl2vQ8
FQAUd1KeElD2PZ0J9Dha/wbcVPZi4mODFOEjrQ82adRqfmHVD+xIthaazcTATfYh
reuCnCAaoj8ZZWJ3eJqT3uj0NkREIJUNLLCsipq8CmYgYc2lT8JTGxU3G0ScUMPV
wQ3zLPDUCKS83xoGEgrFQWXpI7hmL592R9A8cEHWDAwMMQ5FNvF0LZLSHTeUgYRh
MTYUW+IjWXK8CSEsXw83t3LeThHAt7mzgIXfdYooAXjYpvqQn7EzSHm3iJZSZvOz
QGNEuvOn++DQgwIXKMvDJUUafZZ8BwEwBI0Bbbt/yKF1vWhUejuSR1/+HZp+eOnN
lWeOlglTR01LmV6SoJNLf6poE5i4GqxO5IvDk+HATYs5WJaLQ76VjeAj1lYsRfl5
ijpzXzHn4MpqU8+nLVx0Ns5wbO7FGIGzfmSaOxnXO4+ypStzTCGpknHJ/dX70ye+
bXgjFR4Gx0iDtNDTKk1LHaScUDaE40UdMruHAnf4FnPKvCAh8vfv8Q5ODP/Jx3vv
PJyyprCK+/wEXjBGehD8bXm1k+pqtFKwGUa5biFZcPhjcWC8BWsTfCnM0wgc9gtp
oPNEil1wxCsas/sPTBtSxpBksEk7FId0OPvipcKZc473Lvrw9r71rXbYAq7GMlcD
/TnKxJ9rWtwKAQdxB6X4ZrzzecFEICILnKZmZWevEp2A6iuzpxLrHnZw+LBbBKpV
QpW+rm5UHThqbzjWLOVjbTH3rMZ4iEwZdZnKra8DnT9sfJufHbrFT8t7gO4Vb4FA
/0EVHxhtIed7s2dyGM8tr2Uh6AUkAJGUT5XqaSr3hGgJ7DE4E6SzXQn6lVzpj4cx
homr2TBnpcFVoei7HWK+7KmLhsiXtYkOrxdKQR+xN4hAtSsZ7CLpUXbRTFm5vcBH
gt8DDgkrgt9ZW4NiOxQ04kNO0siD8hxQGxO6JT2lUQ6euw1JT7ccM1OOpUreL0Zu
f9y0MyjW5K+6R8/UCyjMxecU7bfvPNWcxioa3kpcM5kPJ454vBGbluevQEJGnn3m
/+zTMJp+x6sTsbmXaZCfYFRb7av9fzWkWV54h4V2JEbA10zq6ERGu2d2tO4Q3xYC
JF6AUA7FH51+Pd3aSiLpa2rHYxwEaiCTb3TN3qLP/aRls73FJC9/433wqn/a5x6F
SgRf37Axpt5BS1lut7tiQUpOxhtR0OBicm23hTFfS7pNIMwJgNBMGDh5jJv+WORN
R/QbhUp6vWnmjkftNhZJrXgq/ejhT+uLTtT81FseVhcbM392sxPL4QAkVcDxa4kH
I6b65eR0bB8aUdheWNlCIXQpAGhp3cNkGx2fKNg0zi+Jz2LkvYkkTNfaGZcjxGdj
DU4GrIUVQXflH+yCkl1pT+ovvG5Tsp2iTWIaxfxKz+HLXqniAxylLlquuzmO1yV3
gPXkR1yfdudr5mn5T/rwwFnNe3diUhQqy/ce+1olsMTbPzULK82jr9YxMRs340Jn
i39leTlgAMLX8YKeiypR0r9MDpcYAcy1wVHJADpCH9308Wus+LOJKCdtTKzH5ilE
78ppsh1PgDUD4VDkoKzJa2skE1A4qPb4iFwnfDPoEpAlORCiQuqCQajo0E41u0uX
Tg7A3Lr8pOPR9eHDSuYJpT98zDEjYgBnUtD4DbCDZGbCKwKM20rMKon5Bdkjhrci
NaPCcIFQIIFMdTGt0cbhrswr0XcQjKsBUXAlB5VfditCo6jKT4zVBIHQa36sTz4t
Y/6SHY3swm2V++7MML0uhU1BQ0Vu2x3eaDVj+XQOQ9XgIpI11Iko/VoFE8+thTwA
h8gplxxrprQxUKOuL2JcIZElo7eYfudlHhXKYPxyiFMu4IUxEfjCxyQALn/Flc9x
ugveQoNHQP8dExzd7xDqBnb/jThtQvR4/sv6AFPh6FbjQzkyLt1Zx8+UvgIl0zSU
aZlxAi5tb/jtEigjHlICIAd85vTIitrdVQI4+zek/AQiaspWur2WSdKBQldUonJx
SzSsJeg5uA9RQkAuA2S0k4Yt5x/90H4b/gFGQb/yRWZLlzfmeX/5mjkQzwe95Wav
5pBjqVcZuTB8uTKAxtWsGtzZv1KFMJBl/StwxX757eBYlYUEj810/l+oi9Gtl0YZ
ZmLjxOCzXvXKyILdMMk+YI6d7jEGP8tS+KPs6uM3tpZdN1p7AESY51sa7SH/7XK5
HpDTzWXK80HPaHqomlY5IcbQwQ0+1Bo130STHPTy50R1R2ptQfKzRD0cZI4CDl3D
eEwS17w0xpXry2jYJnqGy1DsVjYvLMhdA3R2BdtqlJ6UZ1TvL6LIFGpvW+bcv6yk
2V/SPoHFYM8DzymCQP/gqUDkG4IgAnkT8QQckSLxQWaVAo3cryLelGEdtBZt/KIT
eAzAqOJDDHF1nM6C45p2+o6eoQPa9TyClMJnqBOph/M=
`protect END_PROTECTED
