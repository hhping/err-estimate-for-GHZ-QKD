`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/8pRHeMdbgKaXNxuTR+q39eS0lpewhr8Z9Ms5Odoi+Yp6KQQDCTUazugCy8GqpJ
XaWzesZzmWf+ibcptIoF/ZBgA+uFlNPaFJ7NxNVMg/iFbb2fbyNsI5aRuC1T43bN
f0yJzpIwSDTTOi0DJliy19H3zavRkQxEMFUuJPHTv9YB/O0lDvX0OUR6W7wSdF11
3mwp73J/p3J/HsJDuG0Yizqnr7elM9y8ruA/iVve4B0FnWrD2QUj5CibALJEpdCf
qu+Qe2+lp3BUU+qHkzWTxbnnJSC0/Ld5+ztVY1ay3pPVZ8EG4zg3Bci4iZLurjPU
ZA9GHt7ERSmKBth89oN2L8xmoParBC6WwDkj4gyhp8qcUR7g/zmIRp2flix19xgU
U6w9OhzaaSsiPlf2u1DJSfL0amu+t/wsgJ6i2eObHqCNEUIOBzgaM0KL/Q5C+Ozg
Q5gVlco8tDI8yVZO8d2vAioUD+6ST+Z6GgVg63MOcwiolCCzGOZ4b+I6Ddpijs2q
zQGtV+79wyayvcOYdvT3x9wgTALsU5OiO8UEsRqeSjmEATBBC2lgsp0MB+sy+uHP
8N8rB1yUk9/EU5f141uQkMZ9BUVUasqpM0ADI5afxFzBp4pCvkGxod+tw13JIQk1
IDGsvkjc7ZwoIWAVayGAwXgVCXby2ol9d3cEKkjWM72YyrarixAM34JlWRrIvCx6
x/OOLuJICcImhBssPv1clfwol4BAPvCWwR19/3kUYukDtLK07PkBWbOYdmPAwbaG
oa+SqCbMLswEftWV9xu8o6xoG8XSQYZPQXlmitglpy3Jh2d4kUehJGwD8xUewEZX
Rb2a3oLg6k8mL12VrxKDn2w48WM7PKl0cxC3MnopnOlVNAUFG6s8L++UhojS977O
bxz6N76PmTcDso7wZL4zKp2hnK0mohRO34ug3/7fq/84rxFjCyZTDfVSa4obSvzZ
mY8QXezW5JMIvxuz9YakK7gkrw/79SCSohuPHUYXlWWO89EcoSfeqFMLS8eie+1i
2XzuFrNCiQFCbyb2CARsITl/4pp5U0j8XKGI7RPrbkhLVv/iRS8QKda2IBRTOmEo
zp8wXAaMBKCGnUbdbb7L5o+i3IixTJCq/SgJT4C2oQhXcL2qbDAiMIbQ0gsa1nfV
owrrpV8URkyS/vvTTSBLW/1f89HyuPmRvsAcHAVLaLnTrDYSYMAilJuevOZyE634
AUrRGweADkaI5XEG+jI3JzRvh1sHKl91tFKgUcTQk9KdKVAUjFjIVXhs0kloWT/1
d8DAqZ8LbHTeAoNNAHMJiBjKXn7MdnbZS3JlZDgmgg0rl8XMwXdOcG2K56X6QhIA
LS691xpKbdOhiY9Fh9qX8nJl6Dr2oMoXxt5iXV6qlV6qINghVpPT3K+K1DA18sb2
p+YKWWpo7H1q4Osi+pD9nAhF8Ku2kM5vK8Dw+Q55TbmoPBvhZVpZqV8vvSBJKfi1
F7XdefqeZ/vDNeRmGusVGr4vP+3hlZ7qBm+hEYFOgwlkV+u8aSeSEsPzX97NMRtZ
SHi3b1UAh8tLrpQXh2o8mWyLry/g/smonDfzM/G9cGNu0iLqfVuRx7LPhkuTv9xt
7TqQxe6TVlE9S+hVKyv620Hto7DbHvOi0axhmlBYOyy9q89f9pLdpPffDy/9MKT6
k3bjhv3BOExG3a3TjbvlcKu9zvXmaaBXwQOfaLANI9A122asqVBTR38PaIzZJg3T
EkZNCcYMY5eqsTy7Qhb+ntQlgYadOoanrfeaD9MeMB4uBcqBifdcNqEadQzxW0w4
YB+qIXxcRrsDwpaLNmcY75qNACBGGXuQ1Lj470f+ZRNI6va23pMS805OZnrcaYIa
XlyHoWJUp569uDIW6ExX17Seuobammay5hUx7bSsXjvezAzk9DVSyBi4amiFitms
QY5rKc9XUKqE93wLf4/wLMqpphG75LBbRGmO6ovLqAEhAuMAis55hFij4nHDyxp9
5IBaApEu1dhLtqTmy/Js7L49xkxnAZQmp/NZCz1IIJupkZ8nl7hrui3/3BzUJH/I
/j+15eJLQW0GguIp0WNJpFmXNNvh3b3Zg1MDr8zIxjK0vihGMzDp0okfzQzxzpr1
Hp/NiWCll4/ciWm5gEQH8Wzx6v7lx5MdtpKQURF4ibTKdgSIROH/7vma5/mtTG1c
Xw3JpumjexOha5hG9sc7aADBctuFj4B8OBJZWyDUQDMAZ72rPUJPv8BYU6v9mz1o
YtmpaQ6oXzKD6dhqwAR1SLORVV5T2ZaWAnsdLvSQ3qVogLhdGmPFbUWB9ikin8U8
9akXOBV2jkxj5M3NNFQ42yySBO5SUZnremG3En5TO19Bw/YOosKGM39AXHUcZM1f
Tz+Q5Zqw++lzW1pMWYFFqZ36636PWC6HhcAZP4MneZWUp1CC86SnurMQJLKmEFK5
IIbMIrmbh+q46ZHhrk4VpcDcVmB696swxSJ/OMGEBsW5rp3oli9OHAPJ3+L2cqg8
nNs+ESyFNrp7QwBDmwb3BgseS+CC6RufLJiZniAcdIheRSX/yzxrvhUI8ifcK3Qy
p8tp99TAowc7wcGQeFM7BKB3khBoWe5obYWT1VDWxmwH4g1wGDVcc45lie73tX3f
i5F2qLoa7zoxDMUJ7ZakXr8DoFz3JjcUb9A9r3st+hiMMUkgn5MM4Gx7tRaYeM2a
Q3Uqy1gLU83S4i+2asJyfsl6F2Jobzo3ty6ETvzJROPjEU9vJ1DN3LGuqaYYkeUV
0yEaENXlDl8xS1ByF17uZuhzEEAynJsDl7at2bEJ9FsmxBqmqWM7XjpczIs+XpAb
PhMZs8K27LxtcMf8U7NDTse8nL9fHDBQc7NsVUkFvutk5eIQaTv36hgF5dLMLlGJ
PodiMpxHTZg+4AzhKLPdZ3T0u0gfCHF2MYCdYhbq471nJcXzgwtFhULd8xwhjXld
GY+24Q7LMAm3gBjYPYfAEg0pfN9RamH5Nsep3TLEGn+UtXORGNt1kcUjc6xPXC1F
Vc6wqV1ikO62hy27EqVwxzkaWi0pQ16/eiJX30h62nk+fcy64xoVN2mlIM6rmIC1
41F4eLojIpMsWJVlY273b+dAVbP6lIwsJVmMdm9R3eLlI0XyfL40rwQkgSNfqJiv
qPmeVnXDKIrozdVYp1zge9MMkdQGuP5FkMfqALvjxYtRWoqYeGTE4j3V9pdw2jZ+
QWzhjXs1YSj+O4V3JpZS/SJIHPeF+nOm7kuwezGiE7+ysJbl26/ymSaUTwbBw6T6
g2pF/et4ziNPLvS0o0wEWsOB3UPVtyrfy1ftxe1dcE3KbdcIPC919SkD1w5sO4Lw
d6T9/YcZbhoGsJp420GQvSYNpMPJgMadwL9ylzu4/tSqJAta5Tzwrot1DzpuEvSN
IihksXZN5H2i79HDpQz47Yf6vVP5ygyCUk8debF0iYgAK1x9srNomGE/+TKGfXo4
DQWgJZl6KMcqPkgD8mMq4YWqmD3zCOiHy1ET8yptUyhv/0xFyOjOQbr5myHBujr3
Vpro1G4KYoHNUivZ1MSEdvHDzNGIYI/6MoX4PsxODP3F1t8h/FQKpK9lZewLiaBR
wm86TiwNX2uTs9MW5ulmimx+0h6hig//CivWYYR4TZAKWCLTnaX+Itq7VIlEQa8s
ZV5JTI0fug7M2/+ZV2VAavHALWDqlPbFfSE6F7I1QV2mWmN68+4duSirlLr4gpQ9
SjZuJmBq5Ur4m+byjtn/5XfgmfIiLPD2KkdpRFs3J3E8Bdr9HyCZwhdgQVtjxfcY
UV9sQpA474cFqnTPbYQBybl14XqioIim2+5WLSMJwvN3fcpsJYfR2eGiYlt/mHV7
M9hJGZbYlPvcMl4e65kLUwMhVRfpJPnp03j7xze5zCnQdmLBBZq7PdTuf8Cu7YUu
euMgdgJ+BHXnH8kHVm7DUNrHl3OaaVzkMU+iBcYNhZJZgOv7BfzZujHzaRPB8P5c
tHkskQrgH8HJLH00o71EljysB0k89A56gVXR4txOy7I1uzBtak8acf1kxMRQcG/X
ZDTaM0v+Qbc4Pj9DBN1+7wYExwTMpb+SMp37KFo61CzEGX+1DXF0ZWvLke7B36Le
XdSJ2e8lfjyvNIAZ0TgFeyAKQqFm9vmq+yP5duxQCL9DhPs+erlQfweX9Sx2Vs3S
WQZVTLKq2CHYllXoDuSR4CWa1P4RlIMbSeZSlnAOTXHL88vR0LoA5QMRn+PLXq+x
nCikPQT8TJyCGGGAIu6KNdmvcSKCVUPo+bRrfQuQdvHL/ZDUSidZYhX5CHdRBMsU
Irteu+1WkcAIiCWaE9x1/9X7PV3o3osAOALfL/RXX7+YXEBR9hld1DwBeSeqfL5f
rN8Xznnhd/vaFAmtdc77DiK9i+kEghF8XXViHallc+rWvLBecdXdHlez4rZR6ktd
ZrCyJ7LRTxCTNVgr3KY4EcMZeX6WQzz8XrFBpsg79XzauI8lz9AdEK+NcZ3cGa7Z
Gnq/B33RmAIMv6745ZovVN5FZ/1FqXXklg+OSL9RWI73CZJXfLxLLP4xEIRGk+zf
FBuAuygylZOfAh5g0vCvH6Db4kybaIYdLOdMrTQDccnkvwG3EprEJ8BbNLoRyuoM
8F6GHa9FP9ZQQRfNKucOCaiMMaOHz8vv1GFxkQOYyzSza2RS1LWypWHiMFnRKumr
rGAG9g5YUOIBcApQfX9ZU+FdOdJzx8Y8dgVeXYBp+W3i0zGhRSG+KtSIrW1waSEv
cQGeK95hZHW+LuHiGvxJCtSIQfbUmIYUMx4gmuRRHU/0vuG8wbzYxDzpYVomE5mQ
7PNIi+goIsCpeDM/tDEP8KNSeIUJxeVoP8YeWbP81tVC8NDS5tR3agW3X0s42uhC
MYsF7/+cJSFv0CXSTfWfmRPFhtG4MoemFNKNp4h7+V9p5qHGEBoLV2XDAnNSvGE3
oxotOU22dZUd3ys5JLqjpqoCzY8YBBuQzM19nvGYgU3sW/pNWQPh2Cy9QTR5O5tN
9FwgX55+7jQywwAA3k7eaUU3TfOHh1amAO+g+/G6mly7aTBM7QewrN1Nrxf81k5V
QhJ4s1GWZQ9m3kn5+dmExGvCNkGpuFkgk++906f8H+eoDbXKF3NcBILVjvh8bn3X
8gQXKOvbkbNrU1NZdKep7UXr1xly1q5rUhHAz4qUYZVwT0F4XtMbYlYNnCuGBoMt
U1x311mPthYA2MnNzpMXFAEaR9lRTrKxqsGgW6GLUOrKV+qkvX40Hbkgkeo+YQyz
W2oFQ3TNzH83IOQMs7Q47uhXE3TkDU6JveEKVUYg+cNZHLH1pwgoZgBb4ynn65jN
FvxIZcn5osV8W7iphuYX856wzIO+uzD7czWlHxcamefqINcPzmdl4X+uNCkhzfhc
Ng0aZxTyv/FoClKOR018sh4qjHOVSi7RH9/WM3xDKlToer7SYNySIeUHfNeEbGGi
uf1y7Q2nHxb33jOZ/y/368pJFXHgDeqvTZKEH4IyZrjXNf28IzbbZD+IAvltWSUd
1mXhID8cbfokjIL9Ht5/z14vMLKruih/d/BWcmaqADD1FJa7zKQOozUu5KYzOnRj
0wVERqXbjy84Sllb9guvYK3gcOBZTJ5vCYk0jeQ1Wmy7735/5BJsMdFzVmEl5qC4
Ra0TKl++TrpPv1lFygOATTnLL0Z0ISGUDD8tKij9kY8QJhQk5F90ME5ccdhiYn5f
P51Yr7wgNi6Sj2g6ITmF4giKCIGGofohSG6Kpb6zgPxUlnZ6jQv4tBUlBjhExoQG
TF1CKhm21dfdcnY8wJt3/Ji2ScuPjlLzeRWLUDXgGwak84CJDc+RaUVQqEm3QZWz
0S6JIv1hNZqdeY93DlUp3fKuRzVaSoYO8yzeUQgYPEf2fr6LEefBMpQFmo5AyJ1l
W3WQKnQkBhXAYZum2+SGg1FhGajTRPo9K3R/MMgUGqq3e76pDysS4zUL0g0VrbtU
AVW5LE2eBY48nWFDyuigWjAUg7Kk/c2ueSfX+ef3KYGiqOPQRJcR0fQbqKENTJnS
h/QlxGpaiLY6wSPfmpos7X6+WrvWGSjI1zYygZw+yZrdfjU2SX/dqdvoehHl8Qng
v5v6v/HgCtmPLLXZ/miksH+Fcr85NjcJY3u3aH/5b/nswYDzRAjd1mVqZxSyDS99
RxMzeljMM8w2PHHLTsGN9ZVtIap2PINB1bwWSFtdlgHeae4fiwtSyHyWKbsyBI2w
VymdldqOoLVpkw7gvHwV1EQoSkvMcxNpZPeHWTp0jxI4xEG6filBK7mdJLY7fOoK
4gGeMvVP7POcq4NWp6ZSEP3+o4N9haHc1rhRFtKZQV61M0PBoa45/I0tKI9vGkV/
UBfG3ktd0Dc+u9AizK3IbcF5c/NZZaUEnNdxPqbgytH4693HF4C3qNx0/bqZGwst
tUHPOdcoAoidH3iwiQYrnxwRTevixbukPcuh02pp72m2OYiwh7tyqXtZl0dhNGrP
Z7X0wb7xKlsGxNVEyIdRFUpON5nnpgyTLHn9VRgeyb/K6+FDYvUfjSlpvjPfmq1x
eMwfwuIxRAN2rg4H2j/fQXIHJnuVwOPkHDp5sLhQO8XqWi1pu3XJRXDpPbKjMfN/
hZ7mRjRu1YRS3mOzVMoVSI3HdOp/uo8Z9I7w+C1pNNsXxWrtZ8uDCWfzrGbOOaiv
KoEHCe22IDQHTu6Kjalq2jAkV2EcID19q41nqi4TJl5NAz72yp2T4/6HynTX9bQj
qCGBL21lJ472daLQQMkvsml8u8GtckPyPAMX4niXV4F/4F/xcx6OV1oKldDh0RER
56VQKYCQEFJmV4T3+ORzKIUPC0dsiwFWsJrtO/odcDj4QEiP44Sk0eU90WxjduvO
EorC2UbUZI2bCgEPsLLqYLDllbR1opnSlqq+sCIxZZatQmLwac+1Td242U5Shw4d
OrXNiowY8mf7T9bfEKw55U4nM5UPC0Vwrc4PdhBuwnntfOsyGxwocGjDguZWWiWV
oOiI6KCYM8OTxlHwoHIvvHHFXZT87UG8z+Umh1hJ9ZXxUG6ayQ2e/M3pqBOCnH12
SHdBdYAyeZTdJaVtM4FMc1urjwrfwMMyAsUXOua0eKGVzDWDQ0ApZlTLWbLMYMjm
METm9ojzq9/81kBY7uQeQeyVd5uH34OSGV1NJU5H8yWVMcR7nZP61r0709JUd+Py
8DOhk49O9KzUKF6cOdlWZJv5JP1gZCqSv2kRrE9TKRpagJYa/LJ5VfcoS3C2TPui
jHEu5TC2ER8CFOL8O46CiwZMqZ3cZI4zOSDdKBgfg67jfdQXHiP3/tIYfCYyMGMj
sbt6+Ay8jjt+eROnhYlBb5WmFnyNWVFLvHT3uHSXSocAQGRSiTR7VyRvoIFU4+oH
FEVWL/6aK91V0KFRBQNGoVxBwz0AGpOzA8LiEAijCqzkNNyLgnR/LBsDa1qgfy1E
ZR7+kxSNVnUV3NsKJKH38HoNt+w/o9I8DQ9LYwLjScSpLeugPYKWSlXOqufwyjBg
9Xt9UDBIIGJJ7rCI1mwWjODbC2Cvt6qFk2qyX0ME21DdSjtr2UnMMe0Hil/KwFE7
Tez+wdYVGrp7MOyIMraMeA0/av/WtCn0MbHIRZH50yU0h/2aEeO9aYfi5cY5AGu1
YlWMEEPFz/Mr2XjAXHRtu/O4+E+/oiZcTeNTsjQDXdNFqLTammf+RcQ6URBBD/OQ
EHJ0ECKV2pXhVQEc+jznz4UucHWuD5RCy4TTDu7lSUZ0IR4kCS062SxonkQ3jxuq
z2JM1Dr3VSEDi5iqWB2gKpR8E6nN3OFXYeNDxKv3sr1nH6rPj9L+Ou9iAPUMKaLb
L1Y7SxvP1ORkYLMa8XeYoossHmdolELALaxSpF7Fm7fbS6Dj3DD4+tR6ydkrLW03
Eik9L6zL/cP7clh/9B01N4Y33Hc2lHvj+i7/GtWskYTyvAQD/dB4sfHHX8mgz/fI
4mS6eKB6Pn9a4FAkY9cePWmnBppm+6ThX76jItkqJsTpsMPLXLQqyNS1Hqavi6rC
IZmO48wA88LxJYUFJwHbshkoP5Annky04ru7RtBH+fWgU/6VQk5VdTsezK/HOmgK
OYNossWKX+2aUiqS7UcuKIyrik1Kw45wxjyrK0nNp/4B2LFUnY9HBB7UfzqrXoDB
ts8jz5rFquP8k1zkcx8tiCcgz2MYO9BMCIHClL/eA3YmafpWV+7wzBOwpHMFYEDY
fVsEdk/aypYRIynXFFeXwMaL3X3MiCqhCiNuWtB0x0itOxMRVRRUDQd0PDP6zI/n
51NB+CZj2km/bg4K3/XBreC13/zD9rG+pWva6yyog/6NgL5kGqUvr37TGnVtvtK0
autOkxAHIBXEktgT6yRDxyN+DU0eb9PikBqQfaOUa2E35C2Pm1/VrimKplPrUTQy
ixaKnmb9TCwA7yH5cBim0k7zPiBORI0yRJ5ej9NaqmJCsbAP5CECFTSYCQEWNa6j
oiDQeW4Iq9py8X8ScpWa4ByFFaGAwK513q8JKvhRTwZzRrPS3C4UOKcjLzLSyc67
b2rxT2wTMFM6bPS7SCnsGqZJ+TqveK73+sgAockQ0y8=
`protect END_PROTECTED
