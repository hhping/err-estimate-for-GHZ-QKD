`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGDrK6Fe0CgWhp2aiBoEwetosXyJD9vGE/FpKvISIyLnBSB6/kYLIFz5il51s9nn
TwSf5OMDdavP0p/K7HMFCwuVhp88qOzrLV5pYJ/1WSnaGDDR41I1OsCn7XaZB25U
S+i8dP94CdZItLeiaL2SNhnv9eGlal/O1ukKsyZLNVEk3fJ23EiAkaJ+i3yQf4OJ
J1t106IoORxRAaa6I7FBBzL5xSDczkU9alov44rQlvUwh0X9LZ+czHjU8h2fJhYt
PS/zijrpKykSc9vzBmigKSjPr+34nr3vFgE4AbeXg/VtLNG1apklYsgRzORKniZw
h4oOhLYk+7WsgrpUwubHmrPeYDR7SqEEKJ25Zd3PIhZrxI5kSMIybuhnSMDFMt+E
Eba5kALw19jN9Sc2PiXTitVeFbSIkpU52wvz/ku6UipGTonKJhenk8vBlq9P7oXl
AoO4Q4mYHOW84WOJpkEdkX2B4JIFOkLHp0ubKqvmXPU1E70zbNcNafiE9Aervdhh
WEzHr3JtewzIJERZG4rj1wLd6+UEqFeww3nHo9q05PUWxSlamJtagfOnpxGEABCH
LYdkMj/in0HNHGrUjndHr7d7vOiEs37MBFa559LgbzfLte/WqRRtIp2eOB2MqUy5
IgC5wci6Vgi29wbR6FkmPDc+Qoosr6lKZIlTFK65sK8wfFedMqsMiuK2u9qBzj1e
V+xY7jkirR62NsfGUWpO6+RTlTC4D6Q9+KvJHzFYxOzU3QIMNT3x8awDNevSOSHn
4gT3vChEoXNm2ARjDXQWiwemK/F85+iDydBDTG3ng7ppDi5yfGHtMteHBeNBoMwQ
rBdrrkK5NQHI7O6pDkI9j6w/db9NDz2gVRn4l2u2pOWuiPahaDFPZh07uBpj7Ykm
LosePRgHx4wDpn4EvcsA1YT9eIZbfBacu7bG1SEovI042YHwhKzCnIuUpH/6XImT
6rseVANEinxkiHB9wdjYnSS2ya4GgEtrdX8Mu1GirGpfPlMAOIHCMhKkF3LM3+An
qI4ehIfYrRs1iAuqqH05Z+PX0w3isQMYp+e2il3xk6twZfWT9Vc5u050YqvHVaD7
c1EJ7v5iTZa78G4uah4IZ8yvn13jMbFbi/c4RT7Bej70gK99vmEnKgCCeBgiDKwE
rZM96OjeFYP/MfNyQ2xSskEcmkGiyp7e/ToPnoYRxnRc6WavUoBJAekSPgaBDsHr
JMsJ/+NXG0SeWU/fsPMTS+aGTRil1qpsBvXVuE076cjB9uFeOmp+kTybp5GKnkRH
juQPWU+AHXSBhPt25RMRH0jViqDA1HmRZMte28ZZWkyyoZqSX2+XQ6vk1ImpkrtI
itwtKtquVpHu5N1A7fo1XiAxZXS089M2zqrZy4UenJaHccpd0tqIH8t47jmqx2SL
aJC3vqEFBeYHMbNqAyUXYKynphRyCM9TZw98OIG4EKmeAjR6BH5SUONslmr13kQb
wTeo6L7hKIMaqYzVXOyPoNmZT5TaGBG3Hr6m5iPkINseCmAbG9IfaD3GFZS64cM5
4JX4fMQpbkR0jCZ4uPP1uH+nDEb5gojARjE/s+v6lIHhxRUwusfpVAT5L2MXd0xf
JrDDg9n+tn4BuoEnjdjWDSfYBWNLOklhcPzGKCcGaK9/HZ5/WW7G0YuwrezYE2YF
Yulu3o+M//UXZXC5vDlAsuqOjlsyugYYQUL/qVhpEVw9skVOmJJhtmlmtuWy8JBS
UG/nhsAnxb9my49uwUNkgIH52tQnNp0zUTvi4uGF22+CkgMNP+/vjCYAa8rg7Jfj
C/cfBilgEcqpEnhMWrFBfDXXavnw+fsGrFgSn6qDRzC3bINdah/SPqDWjgBk9aux
/osCYXHowphox/yCW9I851JpH7zfpCdZNqhRTUlkhmmRYezgy5qzqqfxAEUD4cGo
XT51bxNpPGMigmc18sgKFPnE3xeupolH5WUl1XkCITYq+Px8guuB85VllS77OajY
GXsQUX0B2ndKf8L6Bl7R4T8u17TBMUIc6+CqT7cJmZkNhcS/mDWI+dmQCLcgCezd
SPk056Kc7Ul7o3gSMUL9f3lSlqKvBAvZF0Vrjb5W0AsPW32x7OOrJyhfluTEH0tX
j4CCMHbASFGxIM8xHB3qlGsPT1DB3g66ZuePQxdUnNUTfgwz+S8fULGum9LJ8SYB
uRitRSNUMhuXiOVlYvHuwBl76UHAtI7lXD81tu6sxwDl5Y/3C8tCq3vimoeNS1lz
7Tx++UkhxLbBUyDmX/+GuPKdUFdz+UVAD4ncTwjqIQzv6Rm+zI0kvWuNEJ7kFAti
R/u1uE819uO9l2rHklm1KubMqOVaR5wMbV2pZ2RhoJE0TEhkQ+x4QWv/orBrsrGF
GpFvvPNJEiaXwyXGtsOSuLCzjn8fvIQQl/6Zf9aITC4j5wgKu4+Yrln6QSc3nK/v
EL755/40Yex569XjFXA8lC3NAkwAbF0s3lfh8/bzE45272A4YfoaDZKc1jBr+3yx
XsS0pLb9JHiGSq70wi+j5XQXUzuvS9w8lLS6+mIvdyHe8YhEmVxpNEXLK8T32fbL
p6mR9TA3ilvuo9OqIwh3pt+Zkl6+Acm7ub/N7D/TFSWOrO0bcO0yUE6DufiMtzb1
5igNIXm1+DeItmnZ5DcI82R1PjPS1UjM9Oz47jTIW8V9k8SdIs93Pl6UgI8fh/JV
tvrgzRfhTBQ60ekSBwhY8f3BLYUoAhW0V9yvyHEQ1vHssoM7rWec1ODexb1M/AeD
jtSbPt/wLz2w3+Wkma9Dfyo9o17TY7rD+LGfBE27hL3iXpuzsmpzAQHlsBHijk1z
bzEp2lphgkrdeisijVuFamo41Ry6LoIpuqMk1sCIVEPcvCJ1I6yZ6WaNasug4mV8
7nbvrayDs+vUVeaW+CkvenH9z9SfyCJENxQL34S6R+ecaGlmWM+FW9d0Gn+KKSV4
anYGA0mO368ucEazEdblLIkIMJsXac+Gd1zBpcxRwU6riUa6hp6u3ZEFfy74TrFO
aF6feW/IypmIF8xyhmfxBxYX87330dvGI0gTec6VBXhT5BRDiB+Mo8cwzf72CPXT
T0PDxr41nVrl8yx1IRIsyRN+RALtGhCyZxT0vNCZVbjOy4RLsb/2aSrea1PWnq+G
J7gOnKmOD4mNJUoMdd/dun1l02dMKJu2rK4G9WqLTA4rqIgtRDFTrNDU8na/Twku
Ktp6ReS3g+13ZcLkzqsxxkcCGWFKavSxxZ4juaTn3/bvfzyepsPoI5yfOrnugRDZ
m7pGERfP677Br4FQzcFJlTMv/EcMDCByyQiGapfB2kwFuGP9ueSxQwwc7T+nkl4h
L7rzP9hrZ0XGxwW7H27oVPJz/PFipxZrWvyW4sK5ra9UlCeB8dap5BR1E8N0dcuc
FicJaMG1DunaAneTTa8jnwwzxP3TuZCA9aeD78oFRzZkvcZz1UvTdw2vsXeg0FvY
rLLj7T0lIWjDE7s0irwYAdpY/1jGREaI3CPmtRChQnj4eflPj6s1UdUQbpgdTrnk
ufWKrQOX5sXJtRnYVKTMVFQIrlM/BmldSiFmILgB1KQK2cEVMWcmETuv9sgFCh5o
Ew1rNtdzc+HxmLJKLZGFJsoXwPBeh2rkN0k2SGQVs1CD3HwVWddkOVWjvySstsBU
4bvHFfy8Aiq/zVjrDiWLkBXO+XDQaVgQCqUaA+oVTsVI2Pzv46lgraJBRwQBDUK2
P1rnCyhJXSF9fRVwshn7BvfLdLZ2U8sCFiiUpTtzMuOSqdzsVh9qg2uw1EvhZE9h
yqNHXpUqqU8f/lVS2+tUdqP5EnWoyRzi1i7ks4xIwz0BwsByzeUsR8ECZ+FcElWm
ayZ10PgZ7VYcQyz0tILsDbSu/oixDbuZUUJmzzzwdsT1u4EEenxfiODLlotbkAdm
avLei264hrciE0Wl4Sa4dcJIxgxo604f+Oet5gcokqETkXgBr5E005nl+jlNyDA0
twolx9bKEKjLpVkdPInSxz4Fsa6/pJ89YqylOlyfbNa0XXFfIg0pjvR/CSRghg6O
yjrXxM0JQ4NpUrCwWVBjfH0GsRpBCRUowoqlFza6LJdY68S7F85wdsWZZmoXREvZ
JPKg9LfOzHkavcy92WSxkOX2OoEQKL4d31xskEEPiqjp6iJ4MiHDGWNhy/BztJi4
9iqKEEV6OugUhTD1djfXJCcliHBXNb/YH1kiZG8zjKN5AvowjPRBjHFbrqeHlP9c
AHk91vZ6rkleQUMFXY0FOVc31nMSxnU/FKbI/de8WVE=
`protect END_PROTECTED
