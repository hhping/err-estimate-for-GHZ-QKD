`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9+teKQZJ1t4IUoncoAItN0LNY9Z9Zo9BhcejAQg2aJ63Z3D1M1uR/vLCftWiJSV
05fZa/oihQo+VdB6fWXQFqq21e4qePsXjptc2xtni2LiAtdR65hogbqLHaUs+ZW4
zIkzatqyiigqAY1ftwNG4F7YPPVVwNIFhLFFYxuUQbJjn24DQjrejur4KosPax5T
kDx1+DJGmBBXI9SGXZYytscUKDd24TwtyEmYwPmt7TRC6Ynsu/0ApZTbyS1qOu1s
+WH9iyNl3YNeGUoVZ+uxUzk39l5ePXpbS6gd5oJN/vkpBQIKyCDL1/jLS9UpbRrT
TpDsBETdNINU0ywBH/T/Ng4Ty9jm8nSLkjG5h10A3mazfmqSj/pvgex14ticQN+z
pNbQdCNMDaPsFxAyttWaUXPRcX125JS9q+rHNG0Ghw08GgczzDFhdRsCiKu1pFmu
FoExQ4SXfJn/RhVyuj4dVv7gtPF1MJYIE6EMjRLNb6SZqM2eeU5hW3nJNAjaIix7
bDuBOJhNQBTw2cVuKypypJ2MH2ksoq3kjLXQ4JzuEhq6zZBkaf8vGCuPVanvVL4Y
RrLRMsfNvA7Pm4+VqgO2jSEs4f8M7ztuy+j8KfZql8FillzgdBvORgZvkmjqhxVr
zw7ErTKgwexpX3CvwO8uvQWLbbgal3fKDPHOTifwkHfSxkkxtLSyJyehLjHw0jwd
95YMp5/EhsYggewLDUen9Z5aGdfnxLBglQcPqLODJ+5RBMqLVIA+ZM7QYScJzdHT
wWmmuiVjD293bVmSzdqk+fw7WSbr1CEvvPP4gfkHv99kO/Hk9FAL6s7O5WHtmWrU
qd7Zgq4SOjt5wBnv4MqiByWoWyHE7Fp5EflMx6EIfP+GefiByAUXdA+dlAgYPCgJ
X8htSwF120sxg/loGxTjtrv5gQ/PmafVCIYhUPgXD39WxqRRbKguqEmvQXWIkOX6
R4lyqVJeU4TPzksI7eI8r5WZ7DxHG35gCMUmRnTvFjQPlIk8RlSzH2Ltvq20WQdr
QfAgcCWNRz+3wJOmgg7/mxXCCTH2+jvTpApuL/wirM+/DEftKmSaq8AcbaKH75Xt
ZIZTjNquHNgNTfN9bNv+P2GMgtMgemELUl/f3U6MEZlYrqigICYdH92MD4US/plr
MbiiidNICq86+x+RQbVbxJpddjuDBvtoG8ptxUR6FKkqEMvNy3frUGPUYvrBNmrV
r8J4e+IEKhXU2ChOepeNXpRMgTX1CsyeN1Oehup6RupUju1iMH2b3r3nj7ZmNdJa
9ZZ+W4o/mvVPweLpdAjr4iCbVgYmLHU4I1ST4jN1/j4z6Bmn2j1AJMVdPGkAXDjn
kHRH1woowEp0FqLNKXOQRnw1j5tt9PGVXJLdRCW6ka+EXTVjMXaO0Od4ddPSjBed
jn1HUP09T24fMEtEksiUg1QssjHdT0ltaw8c7p/aubq6ZNx0eAHaLCbJjjVpkLF9
FpU7uq+yTTuEn0NkZtZ88AGD/cfJd/GCnTQ+qySHdxvKA7ULreTp4GdDlEnyDky8
QgMNVgHHyAZTjhi8tAqszxMVseNpPM8oa+jQpEfxchs6HK9X6uAIxhREERJvjkmQ
DOw+eZovT9RD/TNi9N75oehZKAnbCuO7TIb8Nta4bV+C7BxJDx3NetOq+7cGfUhb
OT3eOCDZYE3uIUQhYUUeghCNVGpSpApDrmECPSC8y7semxWLkvUoejg8kv+ku4X2
WwYeyld4cs47rQAy9AJwNFoVnKSmiXaubKXqVEunsoefomRnbyUhS86jvdYeqcPo
hU1EjKS3c9gAXHDmgpaMq8pkB2r7n95TM73bTU/lZzbgWz7vSlxwnkWiypzzW1Q3
xLPPRyU9QxL5HgqrYZM+/n7+MXh61/1fwdipt8nbr2PSVNjTh0D6QuTCcFYac8O2
jTIR9gdlysSOvQB5p5OIcEW6LjwhGROvh9KdaCGN/NZ7G3StwApoiI9qHK0JzSQS
kdZ6nMb5RNSIVJuIi6xN6g6CDGw2P2TPzX1ZfVnZb/MGibOsRS6BEyJKQtMSnhE0
rCWMzW66rjZ8/8SxsJeSLDjug5yhNoeByWGPPIroUpJKytyX4e3IX42KiQwExW/T
mOCijBbBRViz9wkcWcl4TrhpdMxZuFpRUkD03+AdWx/Q9hKuzjKbphLkV5HVeQaV
fBJVH8CAXi6yng/krS437bJi3r6G1ZqbMywkrGXx0nISK2LeqEU0r/q5v+lqeC+W
AtKpEqJEzOQorJeqHoDSz9cu4ADtc+MW1UEEFGuGw6LlMxJMb29/Nu25Ppix9cgf
WG5cYGt4oVwlZoaJ/T6zlAHRSNYNogLxHFXq5btPAK3/yYBaMzCLOcIF3bQEHGXe
nFy8BRo7+tYKJ2HeLOahy09EwaZUdBFylnDWi+adPojJVS2oxLoumnb27mCyNbo0
oW0VcKlb6zebs/EDpqAkEmnXo1klSUkCxmWNHws6UHMh64gkIH47ZvQ/Cyos8QJJ
F8qtmHVTLWFXA9O4XHe7bLEYvm5wzKguklr9XrIAyP2Id740uhFhS11BcjIzc2ln
cDr/uz4iFcMj9kwrIL2xcK++77aedsBIu5d8sFyaABdrF46eaegOeolVdLABzqNV
BrqIBvbrFc7bR2ebR9Pg9eSXVMcf74UzC9ubotTrVPmwky6+tSlowRLKFDbsyWBT
naIQ/treRHfTf3qxhPQNoxjKP2zAVN77rtfrMLrIcKT8nlTKLecc2NNXFd3be44G
g7oZFmtQAbwz5nvQWmrac5peS96U0ioGOrgUOwUXmFc=
`protect END_PROTECTED
