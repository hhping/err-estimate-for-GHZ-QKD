`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7pw17ar0DZdFyaAKT+zYkKW5DMRvcdHA+hBPMk5HPzmmPmQ6VnNJkrLd/9DLjpU
/NGe2+ssoy8Rl/tCtpuNl6K3uBxZZcjJAJujNb1Ih+C8gye1Up9eZDaUmpRbSiHw
iXZidBlczg201Y/3B3+KotT6J2X5OZuuVTiOhpHmcLE4MfvLCPkcBf0JXTg5W8ml
UmcJFsfwS3/5CiMnyu8Ew8IPGK0/45TtOMhE3coGjWn5lN2BGVCHmYxK4qm+FLZ6
Nmb1BqPmYy8ckmVcotJ4ZN+2F/bHTfie0dxiacpQGbj7tvjcIzMA7VL3JPHOi42z
1GfaNVO2HtFsc6xhgbLsQsUXRy3nbd3SVqSrbdZEVWucGxeVApwi/7sUyptsPFsy
lzvKIyzPiu6i8BpLLJ7frTztye3Bk5aFK1yX5wjQXu69rFbFrVel7rWn6HNYuDny
k8VDWveD9hTwVLmFgSXSnvzpLPOeGyIni5dL1E2ltKyce6xF7ehjsFxsEn+bi/wR
TW0dVYOCCZyMPktumnX+Cfpuo7ZX9oC2Z9wAsezhWVuTycrzkD5uk3mwW5YN+7S9
vssc4ZWxBaUlECxYye8FqyWlxwdP8YzkG/cQA+d7aMpJKYq2tJk+p0Jv+ZkLmGgI
BfyEWACOXlH19N53kRWTUidffcws3L9zg0XMhe65tnWihMvsewg0YF1xxMPR/wKA
qxG1Nb03nnoXrH1Myx9JVe7ZuAwu28RciNGl7bMpgOMXHihSbQcYpm3gIcJy4svW
7uXxU2IpK2i6Ob+uKuKqEfAO9x/8P9SV9uN/lnPSfWmu+nhoyRDvGhIRWLR8XZ+3
Bdwkq+OrVY9WJhxXk7WrZ1DCbswA4yAfrAx2INuBXS1zWzPCb6BB0F69IVu3V5uG
E1IV1ulhtY7q74JwbZ9+5Z3RL+XBdV0QK6HptgxIxWdvMXL+dh+RZTlxBLdNFxWx
FUjoId5vWfYClR2PQ8FapZu2cKT7iVAAD0xdeIajPoniCfqpxSGZpLPgIrzx4HSN
5zdSKSbnm+klofHWowT4h9hG3JooS4GBMNOLKttrFb5Y2D9WJJl8pPEZBuRtV0v9
lQiaB7bFTQuPMO18HcUW3+XbNeFObMA5vzdWfK6Wd5v3pZYWgmDvGIFyr8s+1vka
VOrstEaNIpNq8cpoZSLl7HaaRHVv2AC6AImukQDWQL3nUj7LQx7YayOb+hNxW7Fj
7ga/CKBvq2Rchpq85rJZSDyWK9cpu+DVANzS3myY2keXGsOWCNK3wEQ2v/I5YZmQ
++wYJWIaYBEeXDK382JXzsj78QM3EilNpIO9onr8EA3JYRIrLpAc2aAajk5oK+iM
78NQ84Pcx3YcSFecIvmaTS/g2RYthWqaO2g5VqLDQ3IRM5GL/13FWFNu0YZkCigQ
RgNpFY/adSh909owpNOZmztAj38XmoW10ac6nPMr1GKBGazQ5UuIxVdreUq5sr1d
QgqIKsDJSWfX6vj8OuRpP+BW3QVUSUKDWR7BgbRkKE4bikskH8GnGYV8zAs07rLc
mh7a0s8mY0DSUhZ4k/Ib3b9B/iBIQ8QlOQanfn1rrcJ0SPmnrjQtKk0gd/JFvmsE
NSZxNeV+QHaiuZju2P1nCQmE2C3m7mcCEzlqGbWKLjxp0riHk5Ag9hbPRsi/Uxvy
oZqL30cJLKrWXxZGg4zoV9Coe00ZrfLa5MTdM3KYfvbctOrUuSV6oZ/Lx3uDEQpS
P2/reGGSCB/T9guf35248jcpgcyN0TUerbkpnOMWrVrytoRUa6CGg9Xsui8XWddv
FnYTlJhLzlfn9ZK+97yS9Vdqgy7xBtTg0rWYn/aTNJvPjFBmww97XU+9CRGBlyNq
/tfvZoDWVimNEG4UZY3HV8HpFJxrO/LJWqs4I0PWqjj04brsBWsh9NS2w4uEsjDj
I1KxWYBPqnb+4K11XlN0G9T4N0h2UckHEGA6t/xL6DfZwSk53H6z4tW8x3kgdF7G
VXP19PJPSWJDpYK5mbmS14xB+6CA/FRmQO2Crjlu1Vx1FjdNTQVhUJXYng4mOoCG
VISFKvD3PXtHYYg/MjJwQ/0PwWbJPt2A4s+CuM9Vhi7VGYiyCKQPNM/WZuokm+S0
QpGJg50lRZxC1iAQrioCHSJqUO/vyA5VVZdwdF7NxED20AVl1AB1683n1HdjxT2A
PmVBcXsynBLr8wwkJT06PVlsIuAZVnmKDQZCbGZ+xwt+kKmicn81DK1xUflPmJy2
GhofYgqeu20ApfR/eY/BajcqL9yTZFWruFyfzKofDL3U0hdCztgioiixHgL9GOiD
Vjve3iap/73ZdoezxT5pNL59nsZVYk979VERZ3Z7R3MdbnWHsu0el6HCPgKD68T8
bH0xoX4uVC+OcVbkYUPe4evHI/tvleSayPdkmVTy15dCYhhIn/jv9yKLgwzVEv2S
8+g7lEJ7W7G/O4Zqs6UbERgZnXMuZVbraHFj5t0YtICt0tkR/+wdk4JAr37oeY0p
cTfzRtW7eHJLK74mUGDN+kVQ1A48EDA+9+Gz3AkaSN5k1M32w0pzSKppNukhulXn
wGUL2C5R9qpKDymwDvHzMqjqxHVDWHNeTKvQ2NKhQ/Y/xUzR1thvcXBCtElvtk7O
`protect END_PROTECTED
