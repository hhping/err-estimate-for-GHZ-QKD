`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WBKLpOAhf0b2qhwEFtmrXi6aoiWmKoV0WtBeovOZ2uSa2fETG3ec2xZhdlNvaPu4
nuksbSngcdC4i5XSG8H0ta0o0SgEtvGg/ZTaH678wnUzfoelG4iiCogPHi5BCt1+
ssFPANo1L4ly/gIGwxXnhdJUqBxRunwaKAxV+GaSll8ndr+iwkHqTGxh7MEiKBip
pWmCT9SwN2zsJMVcdEZRYhcp/Vd0s7KBOmXlQjMXr9P9HCmloJ6CFN0UKWhgLjnP
nnGijdkttVlhuzCptjN1VoV528r07weEBqqJVoq24vgMVnaIdqSlcBwmexKduFzm
IBGmvDtnRB6EfRvWS+gWlIYBjUOzNe1vTm+2bVJCqLLPNhzNFnzxltlge1z3qCub
fljH9ufsDz9y+3yn694aQwWqIj7BppH8wJGCAeeCkX0UgN16BzrScMIueqVOEE5m
TY43RuZfkmOHoRBfm1VPiT/Twm9CI8L1z9wwazLJu4ssSp2C5861J96AdIsdhY/A
ZVixBwJhkz18rN/VY04LOfehY1tPXqu3I6qZ48X7Lf6cbUuCPAH7ZmmeNdab2ZtN
hItCCqb/xbylu2lwddz2j822fx6zkpRiq1WFMw9cZl+IYmBrvFE4z3FdqWx8dJQ6
qvjsy9Yg41hSym2CLI3LklbYD4O/SzU/9+nNyYbYfgRew0mscgGR3PljXeqJ87Gy
W5s8xSgVi0gSr2Z5Uvqi1YJhDTj4qdfxXXhikV9c6wlHDRPH8inE7v3Mf8Iy0Db9
sv8hUpctdQSrLVb5IKydTFSJ5syPyR+YIRbR5xNCwdqLmdKmL1RGp2cHFIEYHmuS
mH+P3nYP7GA6WFLnq4lNF9+w4Qctr6F1vHs4Byqil3h+Teldlb4cCSHTaHmVdzZs
vgEo+1NolGEjgtLHGRGKG76tseRfURhzinZ7Fj8DcVJEG3azzkIVQGA+B80TdUjy
OoNf5HXVvgnDobdHwrwES39RM7cMUIq3QNCxQFdDN0WABB9XhFqQ0DvJ9Ee8O1PF
AeUlORTNQj+DXaV3oDxHfcdUTAF8Dh//+yZbG8q7I28oDOjbtTouensmyxcuVC4S
5Nnt5IDJwEao7CzjES95G50eMZrNO0oip5/rNksqSc8f+pocxyAKlYbKGPp+xlrU
6P8aNivgcGs4OgqcZzmf6Xo7d+CPKReAf80MDs9fpv4FH5jdqlOhnUuY48YVLKDu
RAhVORc6u/eBCB5Rp3hMcxPdmH+26/HQPr0TUQOXCfQWHpvIAWKMvls7WTb1KluT
2aZEtF6CSXFIZ9I0kvEO9e5aZVSvdgppMYWXM/XHOM2k0KL0mlDVW8OdPaQoNqOk
Jozu0K/yxkgp+k9pNxCetdCQ584C5qmn1NA/3ufW6c/ctu9UtAlGZgd4mpwZsMRe
KigvMr6zrrHov7hiCZsG1rJ7poPpNgHQJdmzEqai90ZxMEdu17oSn/L4gQ0506y5
LfZei9KvoNDcvyoZ2khTz55ex17wQNkoTRJq/Tg1SHK3Bv49qT1syD6Ge4kBgK5a
0CHcU8ExhKCq3PILrzKsCIEpuZrDgZodgVy+r0QmL+oxzHRnwwKyhWgFUZZKYrHO
LtNDb6dFGAh9C2+1VtUrksOZw1iAp7CRZloUqRObNNy+F/SGTwCWs7hfh2Zv/B3Q
O3D1/0gxoJBJsbQAgxjJUVcWROREb27j5I/7zwg5Sn3HySwx5v0fjjbFQBRVbO4V
iFgJlbWCl9WvZql9QYRU6LPP2SiwOzZi+mCK8JpmAYZwTI5hI/F4zmsJ/bcYYni6
Z3HhZFBpFxn68NgWMmPAqHn0oSyof/TIbHJINfp5Xm4=
`protect END_PROTECTED
