`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gFeC+GI9NmzyEEed4Y+swQDtWvAiifynntm2gVkXTsIafnHnWEARtdsoZ/ND2jn
JvaSikp70KTiEGtCNoqZti7unr/4qh7/CSEFEzegMbOyEkN9m5AuNBGbmI3c5Hg8
7DUqzebPza6MFVwOB/DcNHHxc2eJvc0IHeNPVuoC2QxI+rDx/sNjiSq6Zd8PXnRS
oy05/7FK395OJBv1ZUFf4Ciabxc5nx6FzI+Gcm0y0gz+s+BcXAqxNJs6nFcVY/Ex
05wBsF2espxIlKM94rKnPI/5wi+eevCD0xL7kAuj2Gt9rpEF+yNCLgzCyDHY5aOL
bpAgLUgNiTqVDPk/Z5Cn5miMtI8w8TFB9aTqL8nvRFILEPTCTkXfrGNIU/S/DsLG
SwO5flzbjmhABnIqTKfCsBmzCOebzsvixpyfzDMUx4zZQLN3yOkSm2UnrmIjQF2t
4clqWYvxGBleYd5FM5a0KSGcnHI4gjWKzBDHQ4skpRuVLWifYYeA+GTKENHo/Ein
OtXc5cxDjxLqGSZuyrD+bP4tSDCUuSuL6lvuYuRr/PGYB94K9fgf9n49owhIYaVw
QxPKCANL54Uos0GqC5d7ZmoABHzlXWgPCgXkn+ATpq2pa6VKW07s4eFDoDAGPDSP
p+WaFr6A1o9RsCqkhHhHwHPjyUiKqro7S0W3Nk3GLm1NP2vnOOk5uXlGHZRmJVHE
Sq+GoI/E8dQYf1Xq5cJQM9iRvOCfeXIZmP1h41NUO0ocXpK40EUewVv/A3+vis4s
Ay2WoTiUsH1/3vQ/vtdMT45tvHcmEz8/TM9+ANkDFbuTJ3ZADfiMZEQktsBet9i3
`protect END_PROTECTED
