`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XOIW51ooa9yda+kRJLdXLcM5lFm7aYsYDqVrlraSPVTex37NYy4gH6BOUG8Cobsk
v6pxQapdaPkOYCgneNptBFm9386sElpkot+TQbmYqyWYsU5H3CoRA1nFUPYHp5QF
XKzqNkVC7EotA1iukTvDeGo0k2or4MxY5riUo1xpSXucgIKir8A9U5IsXvK4CxCv
G+HAbWVlUPFQujNkibUtm4zzuFIc+HBqjuCeQ1fddGbQ+uP8AygKQ92YRzNiWVRz
a5bfau/Lk0/n5nDAAbJgLqjD1ebY8VMRdkye72eWaWKsa5vdiywYlWMKcytonmJ+
TGQkxHY8UoiIgBKUkcfx9L3wu0rXsMuthNPAhHDtl24K/a+TDiQRjGJebH0lOT2b
NolpIhGQenwvVQ5QfvIqtI/8Bt0LWMwTT3GPuFS3ejp5zLL5+WIALASmW8P+5q5i
HXA/yuHavMMC15N6vuCuO7dZ5agE9dNByyPou0Gd3QmYtNfn0X/0FLIRF4zGvQkf
2z+rzqWVA+7gkC64146/IIpVDndl7Vv/EsOxMoQGzz59rsbgZpz9azoPclNrJRT2
1e4ZAyF0EpSDCGQz4MvfZBeg0rMrHwdwyTzy2BlQladSv2gQGX/A4Fmin52CSSCj
m8v+j844bK2ygD+4s1+0E0pPvcACm0Zq2yXxwpGy4I8E4NXBjuk0U9S+VrclBoxQ
+BjAQKxUv5xFjn5nvgfXORFNwPDQe9pBWyEGmuEjwUYMJwhEDS1t8l8x10loX0dj
SkQ0mjB+mKn3PzgJ/gf8QCNC6UXkyRvxdbvEXUhmjqdmGewGpjLyWuCZyVMDpGbT
ZpZ/UdS/qYb6l8XG9giVZekk4HEBaD6/3iyv5hMTfHbUImVSfL6UVuBfDn+tYHoJ
oSQmB9fh7fAQ3r118nV+yvNBptPD+DNwDFsg0Jv8C1D7SiQUPLfQs09hh/bHuCI9
2KMT+bXVLtY9jDoKj9HBZCLRNs3XDXQikXU0ZSXhzxAQoeXMv3mtTrjsG3e8GptY
9Hvu3We/6DfsvcdZg49EMCOlzPOuJy+uCfC40zj2PNn56fMIRWBh5TaBxFp9Lgcx
WHpmI8j56g28YzIfFnxWqq6WFwtGEAH+vS54nULhqyJKf04DljcTUHKCU4kPMveu
9kMZhKiZN9dolIeWX0k86eXL4oGlDmWaYl1A+eGDvvvUD/k+kM9dPeMtlvom/GlP
xMvD4TZDiO0eSOU0DOOoCSqsIKdI4OXN8U0hALEtHII+9mYmzIjNATYWM0HzaVx2
D7FqwPzHo17mpS3Cf9reWjB0crYNWQqid8F0tIUfv+N3C7XtmYN96uEusaLW41NW
fQDi2F+ZM5D+VYTQRZhz8N6Yb/Qg35G2CAib5yo/GGMJYHvABe9BLRXse1RjQgIp
ch8cCZ5POxYa+AZ8uhgeaBfCKa24gZo0lEj1PU/7eeqM89sPp1Njg/sfsXQDYK44
08tOoqun+AGd12dGlX5j1ggCQ+DarxS/Isd/czBYnb2nFQLZpFX5q8JMRuAYrc8y
Aa2pi2vyCldgIzst1hx+ZZFsm7LecrcwxZIYp9qKPpAb8VniQsbypWtLkvw0fQGs
4M5OpPfCL/fP7hCE80kLRwQauR7sQbEWn9AEv4EzlOIf/w9FilaSTQjHAkXGeW5Y
G+fIA5MoYajWAv4UvQ16JNTckkW5BtZ6NDZqpqAK362LtMd3R+B4bkO41VYqf6T9
KhmvZVuC9cIepu3uKt92YJCIvbQGdlXPdQxPITZccU5FZRv0qXzRfMkyCct+SHDx
znhl3i0vrZw71rLW6qhPMXCpoFXgawF0VhVspb6DakT6DVavxVAQAfP6OgQ+ZDib
BjpR0lcqvp/1zYOSYOWjkwvOv33cOuO2vS8r9VdM1rPmAvkfc5UO7sGwQXr3KoiD
/FdZGPRTLADYAbWFhma/QGVYe5zsysuxpO0I7qDeSKguYIDhdIhZW09E+84Rr2/M
8F4lYKTHbcVm2R0feGqzrNIaqTNKGo9bUr+i37fx/N5iybL4IMdEtAwFT30jrURy
wkr98/TEmoc8AqWSRKECRNsB5ZxP7U+F2eSUupNQUW24QOaKTi7lhEOLRTxYf9g6
AN500ME+fWFzF1lqfFPYNpElkf9gqWA1Vepy54B76ro9z60FrsDu51yRy527YhAD
o/F6v5Y/USO+nEzOeXW1pzqHllHRicVPiWcBxzrVEQZ641K4MolkZ3AG9g+/L61e
tDPBJLgvROBo+V9NcbWD58InBBGwzLSC/+pAEuQj42LUS3NnRantUTuYjw2jCKS/
C5M4WmS34B1do4UDWGTYGSp/H1NxB+oopemKNgGH98H78XYbqrsLzFinYJNXuKHh
JdcddZjAuNXuI5LgQ5keFjmxG5HQyMHjKARa2z3A00YNO6tavQy795mhQpBXapzl
nnjAGgFmO2ojRC68pkDq5B22t7MmQKeqskcPa8un8aUD4qHX0K/dYDCUjXyxSnIs
VPIazcLEoZYWFZ1qH/cyMtVqMnlg04Z0sCqQhgmxQI2q2MATulIWxK0gxl56iqED
zGDuAAD6NfLeZL54x6IXfH91ZzFmN/UucWH8y+T3jPf3IdGvBcssO51H2xyj9gLL
0VxTcMj+aorqT7Ns+XxvxCkLmr9/ePUj/zx/Va7t+CxN/BTZ3LqX8IEbLJbmlNPV
0TwPELUSDKltSB6msF0gcli+u8LzdLSaIUNzB7rrNLIFsTwqN25bKCEFFV1AY/Eo
rFcTyqE/2SpWcE6Z4Nv/hSfOGm/T/UqvQuFRqMpOjUfjpQuSjDHocT9mBHxhPAbu
kLMl26C8NlpgqepPjZTtd5sAOeidpdkXJ+wCaMcfFHbR2YwWvXSJdHvRDf46mZB1
Cw3Pl3+igJQfcePvwjmc5i/KiYSbYAn7RkUi5ln0Q50ktHN6pppr9+f9dzw8mF/B
idc7dF6ouGe/60H3sTtIFIv4rWnZv/HY996kxQ/Bu6HMm56qo1TU8XheO6YouNhP
BF5tV2iy2MQUIzsowwYwTjSVc+sLVwvdj5sSmdEjFhV2Fcsh3NfHPTjI+Q1I62Qz
9I72yZsFs3beyCT2aC2yFxNmpr4cs6NgZkaKZA/Ha7kCS+Ly8aujIdSE9RSurMNe
I0WldlX/TJxKKoEQ5rh1z14Sf1ZoiO+ZBhBb8XiqysT7Gy582XE3u3UHRpUUKT/3
rNnxfItqrmtsiXeALHfGaQyB95UGYItSkmfJFYebs+ks7nGfjTGt1Iu9veks4qco
SFi/ijXrADRAg8liowGJuHFR7OPEc3Af6kBe6noU7cBnIJdBwpS7CIGpDu3xoeLf
sdLFQb1qHn8gLUhN44syq9PQotsYDDzjEDE9zQOL39/xNMxHAjKZdpKyb3yR04/4
wMX+6hedT6y9MumkeJckYchZJaJ5/yTiojKbI4Z5nw5uFJzp+pI4qyKBcsYQh1b1
NA3nb3yAOTRYaNhccwj3P9Of3W7HK3J1utCbanXpbl7QNGnWbBhWkXVAZ4rJzqe0
M4bzhwTYjlHVjfnZBMud6u0kVv4DaxKUsBobSvZ32pw3g4nMoCS+3ThIk+5WcLLW
/PIDTTdoE8et+JFZ06xzT4ZdlSmiKgGoxxbmisifvlOARQk3v4Irz8giDRei6R8T
PHHMUeX+f4sVXWwbDgWLc65n+ha3X53WYFSzWOGnWJLYyzZ3XUpYU08ZtePRqe6u
K0zAEKPdgDGMhjMjMESHVOct3cPn/YATFz9ntQIdkipOCBOoeoaBf1uUxsb97kza
isq6TrFNAsF4wxk3Ny9UrCO+MYOuYoo+Vf4lxCxDNos8VMeDw18cfMDuatlKUAIe
VjhbQvC2qxLsZxAKJ64j95G2QeH+Ci6aFEsDxc1bY8wpcwc6FBUy7ZRTocazJkiX
GqBqH7saAWNJ/LQGj024QS4vy/O0oZWGYPDlCvJmaJn/2GqR8YBmTPayhdhLq3pW
bglFoTlXBr8lNlEk9mcoSkhejurT2RwsdyiGwM5mjEfz3FTHiYnU8NXoWSFUYlV0
Q7VRvpW83as/Rv6CyXv9CaDGkI6fPlGCS5a1qy8fxRQjovA0rkwpXUIDaKluOwRk
9YzO0fPR61dK1gGVVYRxRnMDggRFtGzR8a6/7L6QyqTgR3d2OGKbJ6+LAjiZytXe
fBD0fQhUUvg3CpIIhlPRyFJRtbUFR+SGwXGIkkYLhyz2vAekIDFOSOWZuKjeK0xu
uwImKUaAWDeL4S8Fi20w1IDne4BC9J6eD550frBcqtlcT6F3aDgjwQpxf/TpaciX
LK4zIOKHK8Es8O33SeZm/2l1HbV5mIHGdiCmts949PSH5S+etpr4V6aNLalOCmSX
muEIU0iLXuDHf20qsTlhzG5pMAiSg22w6yp9Whu7DJg+1WqozVYv3UKCPN7lkznG
Qg1u+CF6UXqHTId9Obvs+pptkBkADb+rXjE+dEMSPSt/SLZMG/TQvthYfrfd/gVW
BCjjOy2YVB447pORP7XtEh1ABNv1ReKtT3FAlwlAmVmKPWD+qSPUQxiHoWvnq+TB
AyOFAwm2hzETns4nugS8H94dZDBAsRQyYcyMO2ckSuUJKqgcZHe0IHcIxjcZmVeD
pfzb8JY9VF0ReS+mUvJVnG286ZrTdgrRaaiFMe00yPQ8/nORTg+quVQnubUBNyp0
K6arrK4BOiDIn6gR3GiEhdZm+0j7p1giketQq4pwxz1KsvCRlTPp7Gt3C48N1ZKZ
IZyztzM4s7kyC46ZAS6smJzdL1WmEqBRsYHVFP//1qrUe6AhV0QeyNd3k8FhOinn
ZXPwIaQXpugz2ybv7sz5HL+ouZpH6vgTCzt9ZyrhEkXfvIdRXh7F7bTRBq4oBzUn
HmxbM98RY2lNNJNZ+q2mpHOXDptkvM4jBpCWFllvKng=
`protect END_PROTECTED
