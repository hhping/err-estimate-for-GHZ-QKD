`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r/8bXYdFdwubBr6CK5ohF7HsBNarsXgPqaBpKZzZzSW7UfHPa2euUc6XeMGQxWxb
y6INRxLpcZr7/BcWuo3rpKljwI3MxrUUsat5n/NCQLn+aNQpQ4Gm5oMItpbKCthw
1sp09ujXGE9tD/m+PMCqDANhGHymFni1njL8831nXWtC8UAQcUCWZzLj3XNaNJQq
cE6YWRONoMA27ZKcnwxa3YsW6Q/sN/i47qcwWwl3VPsf2RhY8me8MNinGG8dhdGU
BwYWfhcyTbNQNuLz1wEq9HqlcVORILGHnFZJa3UuOFG7xBqSXBLanbuRO9Kla3JM
+yXtcEM34gLFJxu44Jd54FfEy28rZhENi2J/PEqkBEOMZRS7jE/ecNjDcVUrDt4/
tOickPQoxSQEiIXbLIpA2ntYwEU0uTrUNitu45EXCDtn0dZLk9OUP8D2hf7EmTiF
tM7UScqxd3KQWwXqwe7sLBiOkxwMhlY6N91LOuRb10oZutcGgaNKFatqT8HmZzFB
U+/1tq3M75I+GG3l4q2y9UEqMl9DksHt+Q0FHtlKd7AydY3rFb07kv5BXpHh9VU/
LGR+qV34khvhAifIyVMa9kNOIdL9UPe44PNbm3rYyIJ5JJQDaqAef2ectN+sNzT/
H1waN3BPe1EsLpmvtf5Wl8Ct1DJWY5FF2WmULaOWlprlN4p5jrijScvwDNOfxA2x
Qc08/aaU13sWJQC16Je7rFF9OJqRpFO/A+T3+178SESU/LVvKcFRcH3Ktk6pPmtH
lPvr8ve4hW8z+5FiScvVULfbanWZcUPatfbXFfDzkSR0gl3N2PyvfYoo9Obt7nTw
c6E1iGfa8F/6iPlz9meQSMaUgpbBxD5g1sUr1lThgf4uLKnewI8IWZKPQxjU92r9
ZXJEvyjKsckJmYefsZ8n63WagH2O+owUfINMsNs3nAe/3gzH9i4LvUWgsy5kxXjC
P5RAeZvBMyTtdzCeahIv0nh+xa1TrXJ9dx5HWlP39XND/7xh+rNRdy4tpwqaPFKi
oMFOFV9zWHdDNZIKcGMccIWviMSdgIGQ98oy17gb8Vbtfb+fa23AeHldgfK4hsX0
IgC10kHhHI6KScvl/lon8xEbYYM+tF8MTxcMMCkmygGobP7Add6eiwPTAfuIz0gR
w2NdxC24hs5kR9cpMtCwEGSC0WaLuh6QpvesbbzZoXobldZWIH8YNUBoc9cbh3Pn
8mLsODsmYbPmGhIqhYaB1roTbUNfiyVNhd7G7IaM987GvPVgFWoZVJl4KhQGKRXO
IkrQhBzSCfvO7IwD4d10iw==
`protect END_PROTECTED
