`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4F2nlO3sFh5uvb1o4JA+qbneijQqYQWAuj7isId2euNOb3sTjnnnmAACNp7ZE4hk
RBw0HZ6X7sDNDi9zWFJfJu4ZiVOLAZoflMa1Z1GUSOc41xegFDWdGMwIfaOuJO/M
1FrAcsQoSbH+5nakfy2ZmmuVP8KFrtkNQICWBjMVBhKNPB8DRNA4gKB8pGMkR6kL
by56MeawYr7Ysihd/4m1bg6RNGveaEwNloXW1y8LFxJGm/oSWxStg0KoTJ1KFCGr
lN8k3n+Bf647VmEC21nlYB/Ed3a/AbuJA6LgWHkmQ7OToHztMJo0I4vUEvoDKCd1
g79447fZLNAOkxmZpYejtq+FwXlJoETM2W2NEds9FabhevI6I8whO07q7z9kOxd7
Y1x2nKcnPI+HRhM3K9vUifTuAzu0AQquaQWKfX4AnTlkKrJkYAjWFjiEahHDL1qn
p5RbcIuCBPFqEOKTTOGddS2M2X8UqlLUJJGyv/eC/gudn4Teipicy1Yo/c40W2jG
ZnlnbeTrPKdPwyYsGKgVPsupth9GyNuxuDP3HpwR5652AR+wcN0WES9GLHl6QHl/
wSX+cpm0ewsddK9G5+4MNAebmr+HyM0uAfZ01JwJXR2DuHZPljrLgjdB4KM6h8dq
vKXriagy4WAicyRDDnc3Zg+RtjD/jYlaEAakgHmC5oTKUL6kYxd47dansWfUlQl9
hZiA78EJ9GM7DCtmHP7t/Qj5euJ0uk7MTvTQQ6wYGmlKar57AYLx6x6lMb0IgL0P
jDwOOzbaMSTGALghaX9q7Whf+TpboF2KBEGvJeTR1bOZ7P7cvq/+m+FhZL7GOhiR
7tLKessJFr2tlA/t1RHbSukP135SJDpw9MM2J9e+xEzujMSW8hFbtbnNkblAXmAb
0tDPZXpcmGjViriw2uw3kcQ39mtsNjJEOypd2jMjGXQc2pZovQgXwzcgkIe+jBnc
iAsEs+ZTqoaZqkaa1EJZxszCKeWp8ZdG2rgWVXFcaUQNPV/9keutYhI35G21zhpr
`protect END_PROTECTED
