`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S9P98xc/BLkdU89zdrRfw4IN+CjfiInqny3Jwh73F85v3LjynJioYrpxvnFsCSvQ
WPyEFP/mvj34atRubKbZehQKpPT+Ncdkvf1PA3JG7lJhZgjEHep0AicqnxpFF0IS
6fJOTVkVhDnYt7h5FZJkcwFldJxByVd2yh1KA2xMwbo7swCCQPAX33+q9AxaH4E8
tHQDP4CYH4Vv/MSnnnsUjsjOs4mZ5j0uFWLIiJ3BH916RVm+keA4RFOE/uBgM6P8
sBPDrmJebnT3N6hWEkR2QaKPZImRrDjoADUuo3fumBBpUfPXzmZBFWu1lIpiMvuS
yFfhVxPn4ia72yNllPCl7SZgA7pE5Ag7Z/r9upMU4XX4zCBcwNKD7n+S3pcC9ctG
8gXc0R37Y0cSaKVatBIrs1Y1tpRZsYHM6OzUemya8VSYzkCO+5Em4AG00/oynbXb
3PCAvs7Tc3o2GRKqNAA1GqR4NmLrW0z8QMikzS+jgJ3ZKJBiUB5MldU4cXQZxjsD
2ez9DxOq8ORVsmaNB7hnzduJjEPLHmjBgCKdHggCtRjI0hkcwdhMqq8OzM8sNeQe
fWFIUiMYDYZuYl8Vu+v11vO8gcFJfoA+/AoBvPwO1nGPjvzAmLGjdpHX6Pc+uNjs
UExXDTOV3RlC62BrsTa14ZPOIZPNE/9RukMwTjzRQn8x4/WGh3U3xhzBF4ICk/gS
WtT0P2fHFu1zLU2dDdP6c4i0DBJ0lwZpil4zoR3Nj0yVsNez1gT6S9OI7JzR4yPK
7onOK8UfA/bE6nSn+oy12HmguUbhP6fQYKqHbr+tvNRQ+cEHNIuBUztMvvFAfqHi
32IJNKV6zdpIXc75bg1LSbHo+WQneLu7qHb9n5r5d8oe2dl+QNVCiVsVjysVUMbf
QvNy5MhohfJi1R2SoHx+IlSOAxy+vDwGk/KN1oIiYxw3VDbf0NfgamQOVZS6Sm7a
Jlz8wbdxIPoKOukJka3ckJDxQBC7tVIVTVILnVhKtKLb2T7zwM513XC2WMuMegLb
+SlJ9CzFDYtsHpGZxoMOwfcG+ULSpArobD+ZAleTccUmKLYXZLeb597IxcPF21K2
UOnPyJczNO4YlWwI5MRmYPEIR0dA32xmGRrxl5yG8Z9aJ4UzUh35Vs2ywLnO1ACH
05DS5K3K6V1/T1CMurNI4t/CY1RIER2nj+r9nnqxbI5Ldb3rlUyI391PJIkZIr89
VcBezHyaSMlVPNx7H/rgWOQGqSCxlilCz5/WtbmqKxGFxrAPOUzqr4UAeJS6dfi1
jmR1NGTGy29OlPXpd0h/nJMa7XEGVPUFYnMz3swTcKVBeus4oX9k//E3OIv/GSbL
OQs/8sVoXj4+mr9dYbayuYPIuRpy2Q/PUjmfUakx/xNXElV7kovMVcNmbp32+tNa
ENS9Y5bF1XtIRzywI8roSLNeCqDGxB4sELpznu7XgyU5AMMHCScMDbv4HNHQQezp
tCf9xZGdZFr1JWyHWyHwyTfE4lPuVVYEc59cBK7C7Y/N/4lZBXhhAe0erAnWZuRd
9q62GbbWgT+MC19/lfuPZPEtCdrNBCib1REV/r8qrIRs8vmK4OuAs35ZE0MgPpab
N6lRQkP4Jy7q9YTSj7XYWKuOzgQDLRMk6rR9VGvFm2qH9ofHMC9lj07pi12phaMK
u5KT5LhosGi9dXzDks/9UjraxMlbUpiyzbGhQF9/akduhnctUzq3Bxq9ELqH77bY
ZwMCLBmaT6luZEQP6YyoUdUkYjS3Z/WUaiYXbTXGkeAJyTSWIwBSjiWPb/GHfz3R
iFuvuyEhu0FnVX6ElD6uTu/vVe2nYExhUoiGWDJaq1SGQNlDe+duh+ZTl0iP6ca5
zsxjOc53QR/gRLao5oCFqBkiyfN10wEmClP4n0PjZIBuVhkF4Q13IglubR/a2Kmp
qjTsGfL9W5AxAJmLvQsHB1xFUZuap/6guI97oEXaX8hcjSwNhsgwwHYqClPOoZwy
g+oiH04OoEgFEy/tJLMPjgD4fv0A6KZoGH7cEHHAtlU9uOaJhbAObhLYbzL0ST9U
C8gtMVnSSWeQ67VgH/oQax2jPjM2LDQpH7JER5K8t7P3CvVdV4oWh5XmyhemN7/H
tT5iYzI2JGvymUhol6utWrH0E6Rn1jdbMjXcwc9CGepW4NEpUjt/DUxnjUg/d4aw
H/+HV8WVNneki1xWqSowJYBHwvN08ME/tlld+ObXbQI083zFKLISkTFgCFFcPE+t
iI5l63TNy7J7gnKimxWvkC70InARlNgPCmaxzAWxm8wsPFHXeVWmzcS51G8X7ypL
OQljtjBFHJl4/V3qLnViTd1pAUg1TcXG1fBMZY8cg5mkXW+kE0A6GOeq1N0JQdJ1
JBC2rnSpLoh3uOWgtTG3WkdpyaKrHbfKxEpE+A7hzTdGLYpRsPGYMo7Dh65sVuYi
QJMbev82pydW/G8PL21isgs4YiLh979I+NcFtV9M7gYKk3JjiijG3M2pavQkQqRS
0s6m7yQyYNTY4zUJW+o0gt3aUzZbIOIavGasgTMQCW1oHhkDP+Ii6x7fF0v/3bxx
AZuUrdCQeywR8kwuKqm5Lv4U86FW8/o0IkVpVp0D2z4YhVjzzjLUwOiZhhpZmSZB
Rw/FaeR7udHahqjhiOwZb8TuhcpO+/JB0JME7YsifTXd8KPKunBofVnbmP6DN1aw
1abFcpCYLAK1w9o6gRcnSrpHCGCOy89LDdWjSQ4V++AOttw9y3xue6s4osQs2iBh
jHIiGhDbAM7bBS1vi9xPqx6KhB41uCNVEI6ZQldco9EI3PyNrr67x/8r23lKRztq
8OMowadp4a8iE8pZKaZaXf4cIigukV+12T5IUPGgeNOHFjsxpFX9M7ZNNSMR6NJ7
FXAAg7EWMFO25pSaApKn30TGBnQhdlDqUvVVrcdxzecGVwFl1wRITMeWipLKcogY
WX0hytRmHMwhjsVyqUbUc1wXBBilyQewl40GzxVgv6yCaZxLTvQbaBbPYqurhDYL
MtYIEcgUesb0zrQoXLZMaszGdv2UDrRnfKtHmv6+VsUK4hWD2LaqS9gITulDNL6B
4FKJ+zYNOQwq24PWNNRfmYOReWY6KlMoyuzjJRUrm3iRNTfeHulOEWLlRw0p7izr
sXB17uSgnO2HMPujmI1gBpoqdlDOJaXsriUHO1dag8Cgmbjy0KLGDJmlCL49R4K2
NN4pBB6uY7/+IDQA/Xl6TLXVPmHDdm+9mO2+J3ayLhQgw6qbskn6J2bGC7Yag3/l
CKpLN3Texenn0BzivC5AN3KLa/XuSVQmNj7aVbPe+x1BO7fEoBLJ7Lb3FNfyen4H
TeIoN0RM7AWXevzJptwurQoo77uiBdbgKGXRIGx0J2OhDCgQyCK1vNhm6Fd0qJ7X
+RBgUmXWDa6XZEJe6QSrVdJ33K30qvWMq+rqccvx2khGLRj4CJ30gCXt2vUqCWUy
VL+YPaQYdm5SDbxjwxa3y0C906tYks2wmySbE28tJOp5Cn2F+tOV7Rur9/Jh3eiK
hy0mrtcxM31ZNlWog03sHboC/zfk2V84S7MDNQ9cTgxiFO0vjQLFwzb2WztZe5xu
rn//JOzJnqv4WCiSwMoRVqfyXyZzFs3b4A3ROVikg4YNRpOVuZWlTSKiKILLQ0jZ
Me+W7kjhkXwWa53ACFIsT4HuB8RRG8nt3GhAKQTgdcQ5asSwhe4waGfYwdoyCR4p
xcaX5u7oUG0hw5gwMZhASjViEBDdjph3N40rQ86e0sFDDxp9pIe0bo9s78amykP5
D+eDyN0XQu0K7eW6aj9YHtHklW/gW3acBueDqVhKWB5qPPHmU9OuqZnXRS3KsFdP
O7aT9/xq1ms6ykokV/L3t50Z9vfB6MAP4ys4WMVDaBaTEyElv29qEWerqbvXV9wQ
igUmuBXGklTO2JkY9w0L+zeiaFDHwqLegxcNLmdntLqscd/Yd9WYSbfWXeiAlVmM
X0Czarr7i7MOf80PafM8av6BsQ4xJN1/lbEOW02KL39fyffdbbCxM70UVyFKa3jO
d6GztTE9Almu95HUabWD4p9c9nEffgQ6uM7GcKbkVdqVhQpbTtYaL9sdcu4O6LKL
pGbuYEuY3fcP484g1lho8P7HVuxisDMoM6xQ9hcycEJ58GgGoh6G/qXsAb46RLxE
2e7s8SENzGV1kl12Bo1FCK+MM+kKQZhEvcNhVl6aPKU5UpWQguC8wcgDV1KHoMLA
lseXcq89zdkmiJkPFrQQ8k15MfCgV1/kY/Ygp4azDp8hF/eRz5+Xi+g31w7UppRS
QXkNEVp+bPy2djZLR251FqqhadKbmPWOV0C5iTFyOxgT51ujdGEqKr5uu08TKktO
nkk6a5l2m7b3XwWpM0k9qHL3+jEhKIwEw1T7UVVeiWHeiOk94AeIIpYEmrx6Ge2j
+BRWBdE4CAZ+vk0QYEEY/l/baBIOcRF/dqcHfNN2/8ucbAKCevhIFa9Weo2TyaaV
PRPgpzRMiiCFJjtC7GLHAhVb4RCT2df0jFL483SViae61SKlVhYViguiAFW+WLgW
j2ElIrC3JULNYovHvcSOnhGtEBWy+46WHswcsSURDIcG7PPojjbj3yHXHxnZlJgM
ZIPZprYxq5geOHY3T/eQrkoLlVHLySWbu5LUtBfdh3aR/B+MxhbfZzRGe3MFJ5lw
595ktAVMsCMhhm0GtMMcLltUxOpJAyiKL2Qzdq8pgiBmTqc+xguWd8/tCMFVAHUL
ZweJ10jlj3tP21Nhhmb3Daf60JvU5zki5weAMSSMncnT0m7kQW34LElAx97BFyg5
mWAt5M3UJFz/katdQuDahaQv4z1khsfZKnj9AcwV+kIzJEAmSIh57cRR8VYgrrCo
LF8he92vs3A/IPWluedwj9Chlej+TjyTuln4T7pVogGoky7NPjIgYnr41EaGIfz5
yamSkLa0UoDUWN7GJjNAtOgoKVbxvNLoJJNZ9iQSZpwJ6O8oCBB16c0FndsOlNjo
gaqxMiB3q1Avh5hRHu5lpbo0ZKm0bGdSlMq/RR93CjlJsb2LAri0NiKP22ht281y
jt9FWzu/M8Ncc6KqtYJqftT+qu1u4YP6FU1nBDEwRWBW5g7D1XQmQttSFAyepdMR
DFZ/AaeqGd4AVEndnTbmm6RJ/CEJIW4hP3IhlHZa5DMp6vIvH+Et36YFjY5lLrC1
p4+2GgVhUDmyksWnmF9FZdnKbrVyPcBT2SROCzvjXRn8kn3m3pzCWDaeZEoFjytl
lqyDeIZQf3XuHIZyxeA2fr/aX9sXWqeL2U2dBFI46p3Uj/tsBRCHaTCAKrTC86Rd
KkEeI19oY+fzDtuSBLC9mrSqq6RT35oiNhkiAW3Ks7sdhpxklJWahtuuC9cBZ7fr
igXMJaquy264Vunic/lZ9GSH0DBPG04WGWWCXd8Iun/bWqAms/RgPEEUaIXtFdM3
dYFepl4ywrcOBa9bv2fI08oxB3K9gjgitAOtfDSmnCn9l5ikA0yCvPcJ+meIzOhL
xchZW8MC1bTZGoPnEkghCFc7OK3YH5TqpsmY3Ok4R6pq5tvSQJK9gdUtVTT1IfF4
wyL4u8PwbFp0fZFFDir9ixTP5rzsxTlY3TJoXJpX7sUd+fK6WP8dvxx8gEScCt4I
A5MRh3zpYHw3uKyZzH/2l0Ly/clJmoQh+Savam5eAw5TtLwoCTUnBnD8ho9igPBR
P9oev22B3pinGX7AZV4siwCT819sj1us3LEmn/+saDHgk/7QVrJGRRByjvWpizsQ
x5YoUgX0x5xhseR3y18ogLUjXxtcz0cfaYt7ZnQkBqMzV9pd8f8C0zJETtipUYi4
VH+Pr27lgCoWIzBpf31B3XhsjfaCKQtvCYxRsB6420lF+I2ZOTkkdg3MkSrYqEd/
ASyVZxMUfYYuVW8w+CNYXHZ2ih4Xxn6iBDDgDEVBgPosYXyGcWG4/dJXfzXulCJ/
P5bIPCqYHu4/cCvnFAEQnUd4f/mcLHLZQmEuSNoRdbKPFO316f8qTFg+GyhZ2KKj
H2VdcrMlBPWmis3i3yDBBrVplRbuBP0+kfn8GVqp2Er3nbhIx9kzTGtTmcNJUD01
2xibjt1X6Clk3HUacaOkIkogxNMNkm4gaS2c58ZmYypXWt9kS44cRWYw4L1T10fc
Sah+HeKbiTooxHrVawZ2MlQZfYnMlwePQZu17IYoO2WHebJN9n7+kBdyuEuRaz1f
VPIlBE4B7QR/KumIZvDU7C3B8c6jZw6i5yobDXtOjB41tXQLMtaV74XOkvAUqkq+
U+TAGeMPW+c3jky53RNaA5rsY/ryEA/FsiuExlwgdguWMIMZaJAvJqBFT8+F7R74
VCPCZ9vPgSI1x8SbHIfWJV0n+kTXEiuiFeqLjjbDVBrNqB2wsFqMGdMrsBiSlYYm
wad860ldKFco95AHbnp9oPguPxoFjPe7h541+66EbET5eXE9E1/LxRTDdI9XKjbU
Jh5A/nnBnSWqMNLp9SH47pBdmkwY8k5UWVKkrpTcV4qZhv20ZBwQIbF/dzkoCAw9
3OlCw/38XsKO88BhG3uGtPfubvkP/C6lM4+FSH9wi2azjXD/FryB5ef/+zBZwdWb
PRZGhvONyqZJqy4ZknjUvcsL0t/z0UfzStmOqnUUCcVm9FMphmJT/pymNHmD/if6
W+U963HyaMTIR2JuijMhUqNWpzY6uQvsS8DH/RJHKkIpEcuPHpbQznx5dElcqqEU
7QoZGRw4ePiPZwXwYUB7a8fEReA1k6XJ7SW8B/WSBU7CjXqmG18lZOfIV5IEyS0Y
rMh5D5ERLmPYhDa4CsQPhv1MInrypj4EABpmE3nurokEJcBm7+Zv8zSJbMQXu1gV
PIXIObY2kQulA2KWxQfhIuVWKCU90jhjPILzb/mPk3n9+1kQctZagOcRSKGyyXsw
9U3E19hket5hGTgFH+/MA6lc4Skn79LbHB1SurE0rfmOe7ZkPhdRa2Ac2a9TgQcY
AKWUGG5MSaJQvBlhCfWPdmPciKPPuJRE3AWTQHe3XiyJrSLOVmhjd9rNAXG8uG6U
neWa9N1obblLZsXnsGXU9mIF1nSucw0/Qt9Wb0PUG/i8B/Q/pK4/YHdunku+rHUN
85Iv8QhGR+Xn0p+tO1t2XG7lM3emVekvKY61WweDnX/YYLKeOlYSGT28HHz12+n+
G3WJZcYyAjZTFI88SD2Aqlp4g848VS+bfp1dQBiO9L8wGHaFoy3qaD3+iRfkwsN1
3jmOKTzvnL6KNN1FhrX+IRcB6epe8Hzt+6hu+oAZ+AOCJnlJ/wtt0ld44SToltSq
/pN8817pn7a58wzl8Ip48BezFj09N3jF1S2XIppMvsJ+GxmgII9qY44t+zVRvH5w
dNvaGgD9sKBne2TFbGPYGs0IriAP5FsEgbD7UILBuMayKu1de7UeHHq/8jzsluSH
FIfj4/Y9AodAYfDfgmTk2SMQQhHv33a+lFB1/jF72iSX7ZMHagZN22k/hNPRJ0eL
xJwBPhNmH/5bAo72sotb3zUlAkZ13FvOzPhDYUxjI6+v6CidqfK3WXmxHHj3o79i
CUGM3mM454eC5f0XAfMguIz2UmS2qDDDCwH+ZsN5bIpZju2Xi24NKIKweqLZ0Z0D
ZwJM02KheGOjpddP6Z35YOPvt6zi5/WqTSs2BIC+6Rivh4Q4j0z74s/pWBKQeBWL
5jnGoVhvREOm4+EYA2P1ud2ZHTkiYgN1TVfV3Iv/W9nAG9ViFaGUVYGhp9YP/MP/
oGyN0y1EuHGjJi8eFx4ueks37uy7TtQTen2oSMCtRu4kprp5ojUlaClEvQcvisMa
/gDL2yqJvwVejDB+rJBO3rAIt+JkFm6Tq+Or1gIX8rbxj5C6VhwjflEjGtrB4p8k
VPwoEhQLNssA+OlboM7Pm5CK22jl/yU2iewTtkMj+E0g7e497PXZgxjSNsRZET8s
mzPfoxU8mNMN6TIB9aeK64MVBRE7FYECpdHbtkpNfNhwzT4Nc+qKqp4SWEQiJQRV
Q27Y9q7jab+AyVSR6UwGyBAi5aLRnT7klnlK4/rhacO6U8s9tvGzjREy6FfcNzge
cnsw2dTMK6Ze1Rb60LBGQ02IqC1BLNP3Sar0fwFT4ik67BOIKpwA2dDAASVNTm7Y
MjgmIOrZdBbV7qHRBuyHWRM57VmgHCiKOxn1eLAWmpnz1sgjDkog9PX9NZ7f3AY8
o3GHYYEm/31Th436WsVGoySSdUcVh8wL8ukJ4wk5A/B6RMYRRBK9tA1pm3Pxd71L
DSbEeE1oo1skCVaCF5lWs6MBXaSuyqhNDCsfmHy4ZY9IvUBS1fbEpyD6RhfuW/56
eGQMLaQTxksV77DOYQJ6de868Ky/8HRr3Ij0pOxd42S8tdV6QvQTfb+kDkKJLf/b
cnyOYp7l/To3MPaxxIWy+T7ypUlTNjKBlRbh7D2eooTx4KWC5eK+VjyYskmTk5Uj
ZXh1kB+yQCWVBXnoZPya/PdfDMEvffZshboLUquJHQ6BD8SKUn7D+g7j47CQo5WU
P6c+S8eyIe8E1KG+CCXXpemdylWlXS33WUl8RS5OxoiujIfdcrEqpw9IODu0RkOS
IuzfcAPxnzXzPkltAi0f9zrGUt/pJyfFYgc63wNz4Mwumsp/tQmQYdUD2QQxCvlj
K2rnPOBiSWmqTEifQsWLCE2iO9e0TzOnjIk+mE7/BE5mJ2LwFSkm58sHlwRGRQqc
+qPBFiHs9IoDAlEb78ErAzSyqCKW74yVZ5P0l3MNfiVV4Jb+UbIJqxkxfUaQG2w5
6O7HMrJMyfkgOEyUbt7D0xKQxksxTC68mBbWABZeJ/uMESyjHtaWfsnVsaV4H1KR
pizgC7PtQGn7bx2x8iXSY22ptjh0cnoKRsrZRMdaB/539U1PFqheOmEwgfCGt8pJ
6epFiZ0vAQw+Nk0H82yvxOm4aDT3TO1YZ5WiPNRiS0OICxJpZkootgNoTynMzEHQ
+BCUMgDKPs/seLMGEqEtwEzgeZyxbtsMJQBXYLdqZqnTPQziCR2MZG8f/NlkYveU
TBMJP7ozw287fUrUpBMLpNVykZZWfQFjD4G6FBkiBua+CXDmZR+QsnTaKNDEe+6K
PF7OkqO1jvzNXrfwjoe9Y3YcBzvA3XYT8ZWu2dBtYKS8qYRxIYj6pcRIr79t+zOe
tN8E8ZcchO6u5lqUkWFe++Iczggs+Q2gDb6I6Kder+geM5AvDf/njHP0rMvqtUVK
UMKTydWDAKq5HaZXqF+om3XkU67gqbwP+npKwOchRMPgCmjQr919btwQfwk+zBRU
GMXD7s7s1Pot8aFKmctWmfONK++/PMmAjrWF11ekHhE/R5vNsE1J2HMFIbGpe73n
xtok3Y4xYbyscd8LjKvmzxXRZrBD4mG1vXxXQNxFtFu/dAFZejMhO9s5iwkzl9po
jkU8HVKVZi3pg5UI+DEorRHI6xBjvbJby5LOUFO+Yhdgf5e2P37Rtg/++O42zPTh
wbXcRSJ/JpL6FbkUEHueG/UQeaV8OgelqPYDkBPh5In9LxkBGQvFMqKf8U+U4duL
iPLjRpUV8SW4IN1RK/SmidsT834CohFiEJGSyvVdeVq+XYqIQiax2czEapi3SyrV
NnA/ocT1C8hL1yoqVfaGX3iz2j1hW50gq1LLYeB43GKmW68HvkQLVn05DcKloD1B
Xkh+GkijGd5ComvtoYh5A3N/Ge6m51l0eZvEvFMuHEiGkwU43JfNkPLuh20baMUV
4ZqTzapAldgwLH7x/e1/Zb8znr+X2VsW65bYllAPNYMvKPCQ0oaBHBG77dNffUnE
76QeSbqCZUrpl3nbeFcsHr9q/F5f3o+ZMkdsIFVvujv27O1Qe/PaTaQQcMsT8htr
BxReI1oM5ojmRj8aPh0v1kOMaV1HxHdd3PLk946mEkRwxre1pP1gHy1dCss8DgZF
tV8fZComACAx4F7MxjyEPBawD/im8rikfOK2gVR7PmleijrDAgpoop+mGp604coL
0ih1j5BF08FTEl3eedFQZMYLU0t4fFFOgx+TaFkurQIiQWMF6VwSQxzR5THwU8qn
3LquW6Cub5zXkAPS/F8vgHXZvDINUefE6LWwqNcm7CB1I23djGMK713WEyCJVC08
G5cxWgBmTN8gprDpM11okpQ+FtUzhv/9QJ3eAIOADyJJl7H5Woov4EwPZ+BVdBMQ
+BCXxr0UONg3PDUNcw6MKcGtWMA7+HJDTiwM/7hX62T8I69Tr4+28hq6+ORvN1pS
9cGa9Eo+vINGoyYrmAeCP9i4OpQwKVaEETx1ML1qw04o4tA7y2uyjOUIBAvEN1bm
1ZziCSV230K4/2cyTgzqJMbFBi3TJAMm2T76AFliQxz8QwIDST6K3LBPKbiSDWad
UusVIXkcymq0wQkE0TN8Q1hkQJSSHZBzLVuT904BuacVQIq3Lkl9CSjrk4TrNAey
De9bPl8l+omxTagC4ToFIZ5eZPt4k5CVOwHFONd3edoTs+pN6o6qhLJosyNgJduP
/9MLecF48QpGW1PhW4k8s/BpQ0LtMgMn5FBSA5/2psWQaoG0RHwtfZRyrV8F9hvG
AVkA944MaXqCG/TUtj2kBasONRn4MgUWL1MVxDwhUtFl69IzYMvKTEvz6+nrPd8J
mthbCsO0EvUEHU6UaKxEH6SKD4e3u5FXVshyMkzHJlbC0voF39/w+hQ+Vl7VRDXA
FdulAwdRMF8niXFRpqGJkWEJrAlfPNzjqgkrIU3Uz3Rc3BHCGQMXcfWxQ6Q4gD3U
wy2TC9RUwjayZ5hwo4pvm1kf3PEmyUeBNsEtz3xwyZejqfZ81JSb+HrBJjWWxorQ
TF/g3XnbCL0pAh5Xsp14ulJ9o7LoYtNYHT8FqV1kMt43ICGkU1POLMIB1sNW+PU1
x8zV/Js7V3FdSk3rlTCxzuAISuxc1i83g08zMG3NPNnY/gM4ma+amHvNDn8vWpAK
VGpBAJ6tlqlnDqXe6Ca4wgRCKrqg949CFEGtWAgmZD/GwcQkAMkItIbEJE/co8Rw
HH64KQmr7ktnxA0Xw44xlrb+Ir+if1c2gBzmJHRGd8eBvdaDr1wq9URY/PG3sycA
U42E8kcwiSjigd8IZsXZbatR02CmGtOHSHn7Jd7fIRgjCuLQZcC2pXnK6L7WZUiv
YeWle/R7jYbm70DcWayzSHVE8UpAe3sKhlDwqiHES5PEI36nW6DmVCOo0H29DAEY
XxrFsbyyaX/W+1iYzGKP1m5LnQzo/NYmId29SM0+1M2PS/EQr1LBGki+4PqsERQv
FnSxG2VIbqhsbIBqDnRU8H9KH7rdmgayPWGrMJ4PuOTIjh3fUGpciBaGWrcc8YVU
4MQGzLKNOpxziKZQaLqrb9TbVwLDhIkuJNfV6pCvmBk547Bu2+5hpVsJ2EqVJMxg
d2ND5YBWbbYZ/6ODlm5MlOqeQXAvWRM/X7zG10PBRxzfV9aFPmur0qI8Cg6XGpMD
MuYz2+PDBHaf81jbe2GuL2zMC/Gu7JASSJT53GreEsg1lT3iggZFDZ7bH7JAOdPZ
WyF65g4axm+Q3qE3ILxtql8bD/kgrrjjOKvXdQZm52qvnIWZ6c6qirDcwiskBBBL
zH0mQad7sRtSpUEPy48oshI2MkQKswLPouK9VQat+J36A1WDJ6Vly0E6CjHzDRxk
qWgfZk8JodTX1fAT9AE2FTOt3e3dTHXz/7Gp8910wk9q737ldvOXvvGkLPoU3wKb
pjTnReVOmfnj6gHYebcV+xqkMKWNI7DhaVSW4z9ex8frzkPL8EYbLJK3JkXK6FdP
Jj/R+68HSCNK+F1fFe23Ix4a6GEQL2pR7Y9JXICb1kIfp3qd0w8SXRHfnE4aT8bv
ABsjrXPLr56HXbvJ6p+SC1xugxMzC3AkQ+MqDSsman6y0WRQaHazyjtkkuqudLZ9
MqekoMKsuqt3NRUNzbYYT0giZTcL4XtN2skGcbDS+bJYbl8J0Z5Lylw8Wd+uer94
dCAzaeV5N0wiwj/SO5gnC8ameZTqCBTLXAf6uC0NbyTfViR/+ifineLWwVIqgk+o
2SvUQxDGQVoYpFT1yAw3Ok148gQrjIptGgY9536l8DFEKL0/cJAxcybAN492md0R
SFqKMKpLQFrwIQbUq7F35luWX61pTTevK0dsPPYCna7TeIk1GWv8D6wQ09TgCrQQ
ZSS4q/z2lsuhjbNtPfW44qP8cDwMftKo4eSKhN7rVky8U1VGHWoU+ibdPfLmROXo
9BAd7GUtEtyQYZ1DA3qO/oCdrmLWIogGq+rKpblutcPvkc4oNwj/Ui37hsv4Jt8H
tjXIRDc4Ig4Xl3VzdtyG2OMA+1067oVs71uhQDgQevlV/DZponvMz4E+lpuGGhSe
fcCrHfSKIKAjO+i+2Z+ry0w2I4tQpKbmPGZlKwKgvrIjcwaHPhd5vG4sk2btIRPb
vfusAjPi91MfLHlEUqF/UflZs9Poo6Yy3Jt2aJMi3haHbzRXLMiWlDvqOHIfTG5A
BBVm9lRoVDD/sz8S273rhrMrDYEW5K5fvepOZAKAP+ntlMun8dNSjw+tWYfqr3Nx
6i3p1i0CIkeZHP9V39Ki9ppHu9jpG0cU6sTszSX4qhnNsUiw8XgnZ34jX+9pnz5l
juFhTRb5hb2lquLGib0I3eAJaZywdSFi9zXC/McRbgFEmF6xzRbvKphf227GUdfY
zNZh4063Hi58jMG25wHvXh+vPM1MVtUcqZOHZ8fkfhzDBBhKKJk9L4uGJjSctLVe
lqNWVpAyoBTuZejWMjlBPp5wf7T6ri/7jvQeI+EZTK2iPwMjVj/tG1nUPuRWP9IH
XA/hWhAxTbTJMvMiGfBCjRW8DeG6uV+dNwkbHfRoHyS2cq//tfF+RxQrR7TO91P3
7bEytguRHtmLgpXq40IJvptVRaJ7QoCZiSfkriNR+S61bcFEBJ9JfmuWddwsIvtG
BzWIqPBWSenHt92QIvtChcH5rYRvq7VIs9RZNK69yV19mfLu+RFCT/L1RcuKLmq6
jY6Xw86FJ7UKBy2lHaFA1PP9NTuk02gKNtsFg2Q6hjxrhgp1y55HnhGIKHvO9+cY
vZf3cAHBHNMHty8ttnTYehu6t+eFmo87xs8BXTDiym6wBDS1LHgZy6HcpTNDDL5R
NR6VIlffgxUoMm8VYvemQakOoYKuxsJRc/28qamhqDBgk0mJG3eDrssIuDlI1dly
ZcPIRAiOvEQnDNUEyh8jCI2YzbK0D4AWXbXb7MjoOhmtIPefVQZ9sU5ouOIflOfn
aFQAejhtTqCdzQdYPN1Ca3xXea14jW1uhCb6vqLc5T+mPAgWlXLULBOQgESs6JYZ
3Lz0tC1HER0uiWpwt9nPEFoCWBlSjtMYmzYCHFm+vyzA2faoieBfyVr7aW7lwZCl
x+dKezgeHDr2l1YnVRKTfs15r+voTUWtV+R2C1PnSamz3TGPFq/kwPB5m67l0ryF
A3s6V43INmdP9avX1rA2mdEgIqvtXNXry8FouPl86XYrCfRrtd5nhIjH5jc2kpwd
ZP0WSZR20tgd8dRX5m1RKdbjrrzBd5ETEsNrhWWGhO0tdDLCH4UHFKUNT3Kum89a
vrBsD5Un7CvsNT953BK4s8XUVKhEqX/Lfn/l/ADVu/PhOxHS0GIepI9+lSKBKVk5
/vzZjSFeqWyQlpJ3jjQpKVOv3joFbydwYNavT8/3gZwCEOz0rUQ2C/fRMJmYWkg1
DOHZVX0KlFoYotajKN6l9F09Vye+dy5H2A9qCToUuqOWtVfYoBbdVh394clrwTxY
YaiRjFzM5Iy+5skIPQb2KzQ9Nw2IEpm2xQa/G85/NTPS3aZTP0HcF4XEHZp5e7z9
KdamjikvxBojuxmmDGVIoE4lVOl4iXmnA5uQmrN72V4km+KEd2Yni3yQ9vs4FR5T
yZXM/JryP7+vRSZlBDP4+W05ZTEFlyg6U83sL6Pa2oxkt1MjhbfXUs5JMQGwKje0
jkfrSMDvYP04h3K7YBm3z1qvJzTE096jxTJzs/7WwvoTXC3IUuswI/Mu+SPF8rSX
tYfZpNOlqpgx4Lc8sD4zGSDya0MqypDCj24TBtA7qKIx9UMJzbRSZm/xicy/F65k
761twLSwDsgfI9tN+AanihMAWfteS+4mjxmkhJEqsdnpRzoaCgozXUXd/l+78hF4
bcYfzx6irwFsUx1h0/4OMZ38YRvRIO6VNoH5K6gAJ0a+BZDWv0xjIi1c49TsDhjL
lqs1RBazvB2nmmw3dVr8Kj0zhqvu44EAezft9BFJ+2d+0Pjnwcj7oUo8PpygocvZ
qytvbyNUG7WSbJkxHnnvstQO+dG9SCFDi5RoOeCGYTmSZvsYmd9dbkUwalDpT3j8
DGpdAvQZhtEwhtDmJ5tkEHIzR2kjaIyh3O+ckPDEWK1q2RaF+aShmcBZ7hG8tji7
A+fmx8srD1ZhGGjRybBTjalGivPlcStM4EUCoO+ZrPktatKEceEuypEjjT6HiDIW
qhosSLc9+HZgqI34bulPaaLV4bhQl2hjh6Qp63liiC19dbkGKYvIUBOjl+Ylz8pz
TSXgX/qWdYkHTTeP1f9n+V+a6DML9Zbwo+XOeoeyBxSHOlsPkL7BjpdpYqDA0Fr3
6hRh2ijUcmbFmOth0CMT7VaPsghr3anmy1jFSp4s7ELCHbUQ6xNfd5iIFTlNj1iU
3ob7YQNlU5RKVoqXHGC5Y+OIP+bYE/FVlqTbgkrubet4ze0aR0j6P5JNce7g7aNc
yHSw4F5sb17KMjcBGH65EcZ01mXHcrCJFixnZuyxhjr8pI6QWPu5VvRkK79XCRxS
oJSEco1G101SAvj2pFA0UgB/iJWn7QWVf8LlXm0qkIK21rsLrk7vYvHviZqJYizp
yqOcmZVhkSgJMWEthYfqH/EjoPeOgI18eyNYadIg60ot8HitjGhfGXaoj9aNfluR
tSEesIfFgvzy+fKA9KeZGSBVeFm8s/BbLY89RhBt6ec3xV88wAhC4ueq88zEUcXX
udkQP+MexQz3U/hy+FAMi9QZniXDJUKk2SQwQtKQuOfQCi3dUT6Bc71jPLSKVDim
JojWAPGRT3LlRS0JIKnTTnxCrST0kzZwlc5P+85Z9TBGmstu496rbKoZu0x6JANF
K9zWpFZlfn4UxhtZ6oG4tqy/0CgOCmltTfmHJPhmZZHpokgq7DN892fh3plOPzWt
m1TEX8Fbax5wqk6iGpQ036rGhFbjbNHGdH1jbjBfnDn/NeSleg3j8ktMNNkc54hq
4IIfKZTxaY2lLS9EHKKwF6d5vGhtqwjZs1oY7auBOBLedyYsehRWgkLxEytHXnL/
50w+3kSNZ2ff1YRqUy0IBAGul5/9+4KI0gFMd28m/olXJ++BcPLMA4Z+qA/zV1na
rByLHeMlXuX+WJDYrwtyGHFJzyRycloc4n4XK7Sh3c82AWF7v/qhtyHWjLWSYxj0
5pDuyE3ya9g2lswn6E/XUVdtP9DpOpRTww8OrNSHQY6uLlA1ThTX9xSiJw4lPu4k
tzeu3zI9L9T5dGnK6AqbNOOioSUiqHrRKZa42efgxcdShyanNvlEa9tnuq8w3iuR
CP7qFZD2L9lealDOGo6Uj1HGhewOmTjh/9o+P0vbnx0MwzhnQJI8Z+zUKeO/TGy9
iWZv+4Y2TVPYls92KdnWc3el/Q7Mofb07EZk2qbS8czhFeBU7/zEdRGoCobpGzb3
D1ftalUlSBTc0gIDUTJ6DrUlw5XkNu1fFvRiYwcljKMHZe6caVSqSyMx3ayAOvY8
O3qa1akmgOk7zplATvHEpO2IQ3EGm1rxATX0EBGJN2MEKpBBqeHcKcwuXwGeWN+v
4LfMxrZPYBG1Et6pibBxmBioY7058hdPt3bc/5Q6dQRKoN3Pjch+xGl7IPY56IMG
1zD7bbNyRkf52hIJtAvlweIsWfHIiewQ9GiCFlqeRmP7Qum+0OfcbIsn7xZEFx2N
xj3DJ7o6ZcT1JllsDBc5cWHAAFPz1cV1ngY5QaJXVXbSd/cgM4Pn6KjHbzeAMYHG
EHA92bKVLivCgNrjceqelwogRJVq0nRL0I02m+01GB0CbpVjsq7IRc1cbr7Ow5nF
/qm2am8klgULgMNl/Q4eBE/xY1lufD3lQF6I/8mFOzCaK19X2yCAAVVRTrnbipps
YRc39r7ycsuObuOiUrLUMl/lahSx9DGBLbXheKaLYE/64j6EViLAlloQNUhRic8c
Z2OSUhE26v4JhL8SMJedmmiqLKxcHcYw6Uk8qAhSuTXHmNOtNMJ+y5MLlWrI7HMz
cKTE6PrjzlltP/E1r8xbSBaSAlwOHyHuOovgiyhR5PqAy+tFymV3sLZg90EpyZ+c
Rlh56tJO4IIMpuYbmdfer2578J7IqmOVIp1hSQPezkZ3ciT3mxEp9v5rm8IMYSpO
YGyJrrlql+qqsMGPYTOBLvWSJy54PKDmUmtyhg5hk1ylJ8bFpuO+GIei3O/AHafO
H/kCwN/zksDXMsR3jhWqHFF+YQHTB0K/wwjFH31ekb4vb7zO1bazivt/nqU7YNBx
twb2l6vcbiQu4Ppxht2SuZ2gxKRx3XOL7DuzycT0E7OwIe2EY4z9L7eOyy8c1CQW
dBu5VeWtCk7s0Fp/IexXlbPHY0ANrjTiCyP9Ms3GaKEnsKrv1YzWMUBTRxDhUjYk
MonZDem/Z2svJ6lN4aT9sfjQPuu8fj59IPGJfqgUmwK8GOM8IxyGUJ9tt42y1APp
djVYwVu4piOZs3hgOdZ2aKCtwgCZVpMOrHRUpktmPtaGF2/5BDANzJPuMM/DVztJ
Hp2mxv66ZvzFmooHGToDIb5+XsMsUQOkDzVVTADiiOBPTWMHwMQkn9K5+TptRIYx
u/bSTl1r6j8GY+f/qNq5yLxYojrwRVDykEELiJW0xAaB+l2ddIo5DuUg0t5hctst
bPhQFyix246LCZ70FJohuT40DSjXVP+O9XZnh+Tt/tfkNYWcLECTuhJqDbjx8NQs
OCp72+vX8FmGTPbsxtgtKngqwTsk9knMlobffC+Vbp32/evWozYRqTLVV0Ls2SFw
R52/tGrby9vErld5ESfkilPROal8npe5eNdpwGPixkgpDDL0ad+b+bjODxOQgFFW
QL2NZm1kuQfk2Wxjmfqln/35lUDk2141G/p6GbNAbt3pYT1/6JXxrROhtre9RfzN
xR2EFNLSGF4eCGjNVnfx9STwrFgS6EFlfLcdWLI2sM86pD0piV3IX/nYsOpU1Mk3
MAzk8zSYRWvnePfwe0IAu1KzOyOQLK56oS7jUgFiGSZ67CX7yasCQI+8fyZLokQp
XoUaj3D8kNO031cYjqX/0nrDTnGGKrHxCFSFHEaQ1Y8UfDMqFqzwUa4vCP1e2Z2S
99V9lM3qcJIca+oUvsy0DJ7TrWzrR6Yp5IDQgXnRAA25fNlzbcrM8oYiWbHLxJru
j5nOmusLJ8SP6UuJ8hYhYjV/E7Dj8KgxM9fP89JG/XkApf0mJH+w06jW8pj5EkQG
pQWLkebdj4Um4/2HEZe2dKrhKzH2I95lCieGJcBARs4bAp3OkSE/hmMTQOnU/5vg
ZH4YIxg1qIPmC4O/5W9xZaWsL/15XepqRKLLv9O+nHofuXbFpHJsG+hEvkVLFZSZ
pE+fAGoc15XKb/TKIBlUxOM2JTHhv0HX7ghyECTOVSHE20kZV7v0UzPywynpuRk7
bBLaXPWQm6XJSHY6yyqxZK0T5wF0St6Z4FwpW1nA//AleD8AtCXnI9FhPUbxomgF
UCyGC84kjiz5UXMUj3S7z6FIozi5JO2FQoSHJ1ijJp+1qcRTUd+Ti7QDe0OZhYBe
KPsk6Ofh3y+Cf+pcPiUhrnc2E1bOqr2/XO0x+8c0NwwVGuOY9Lbo5Ba553eQ9FHX
7+g/AdXKPI6xUidFCZUCc+6S5ydQDeaf719gtb8GgonE4tVtVwDYOz7VLmT8nQ8z
AJmviadWH4+4oXLFW0Jm6I4fKFyo6Fyzcx3Set9T86EgkMmOHe141dLiPMTvZyFT
pZgTNxOBXx9rWLsQG7D677ZmU0nAsOPPYbFtzWzT/vx1bU2H5H3ATXN/D4LRH0yv
pp/yvjXI7Rwldahx7isBPWS1V3OELnR2MQ00iJ5gOYXucB7xLeAi9c7rpeNSQ1y/
PT4+6/8p1CwTmMwv3nss1YvLQyYEg7Be38LVEh0PeyOHEQGhjlVbTBElEwOlZL9H
2DDVpwU0hya3lS2LUI1wOwoemF/pojUFEDiNicLBWnNBTfPK2Jtco4PdfAVAdxUr
mPPRY9oUdaXqLxpczHxDeP0Z/SoiYltgh0n4gz7gX7NvGlkHRicNHudnHJtr46CE
lyAPZUwtoGTB/TeVpEAe4faWJdkTI5dWs5m8SdCvk/96b20c1AtFIDXTJo7uNqku
yyE3HtMbtF/8PGDg2r8HtLfW2LCMyEaJ6XWf4J2ttQywKOLgoa4kvgcyOsIGLpfh
38/O8Ag4y4zj0y0tqCW4SDecHprJd+WSuL1xdaVu3soVg4TS1OEnID059jqzT2Id
JCD2JCAX4c7ZprJOTX/MJVjiP9NALn/clwtB2iU3V1cNG5F/XQGNLJl4hqC0HINY
OuRoLsJ0KSpqhZZ/ZAjVnFpFf9eeTLP0BK/Ior4V3M8d+FMTOm80EjHHk0eCYmvj
YsqcD9aV0UjTbYB1abkndHrqD8iABWCmKXubMuSLbCKXmNvM3kyb0nHg78GQAN7b
Q9PAgflxLQHic4gmaAnAhNzxZsBrP3wpPufMBb4P8L5nf/M06VBzNleaxDwjfna0
ZLeT1M87A+m5um+f/0Sua79N8bgyVsmDaERIeY4eBBygC168+LiweTXSIQhMQh/Y
I5QRbeBw8FkqhzejfrUxczt7ZhTol3uSaLByNYl6cDRwy+JsezV5i03e1tWcpNql
YP4LrXO0DvG2ot9e76sjN9N7L4wKMTEnAPFkvH/raoOtEGsHGIaxJZWDHMRFXdGX
X41DP0lvdqWKgzK0wTKWKSyIeIQVECBIZ2PWG8ItjMMACoafD1OaP5QO/qKNDiUh
cKR/yeFTAT6puIVCTO/NSt1AfJDHuHHwwe4miSGv8KUsd0u7tyBYaGE0628hgSWr
kwjVYKk+88Ao9ZrE+g3OqZd1PTtChBJrLPp9HImkGG6Uq6GVdpjnYYqgJnumBVOP
2nZdbXsATVcYB36Gtt9RlFkhoV13BEmhkBztu9L+I5jFq8subIqnnOjjx1WDJBsR
HPNUU23U+5kyQZb9o1UX1qhU/EZdUPN9eaFSCZayiDxUzeZKYr6d3byu4vy9tEVM
pmtTPIZFMF6ukLAtPUk/9aKTiwr0/FSiOnaKs1iHC4hYeuxnvKJGxo7IGJqQ/TWl
d1jm3PoDAMryiQCu0MIdIf1AdsZHreriLLszvcyI1LbJSeFpQo0hn2Q9y/34a3Tf
X8h4EjktevDXRx90HQN2zgX4Zy0A95rQAUe8gfoYyJ97PBX6RSNl/stwPZHPVCJr
gNMRdwKK4LpFVcqyTp/41J7+/S23snXyKh+NwTbgZVtfMceBdO7CPho5yhojBRke
sj47byyD+HVprXBYS7BryQwePOCfaHK72JCKCxQq+fIXs2nQJ0ptPcgvnhkYxEsa
Jz0PgiHe0kCWZCSo4/mIKtdbbTa1is00IpomfxjVdqxvgKVcTbwk7/j3GvsGEopp
GnQ1/uYAis+TXtrCtcr/GQkHjz9T3OKXu7cw/QMcOrE1dvSQ2WM4LIBBoQN8oFgC
1aP03sHLoafhTzaQ7uBiLLgW5y+FQLnavdwFqkosso3mIrK8G6XrfrJ/szJUngsm
/nvQx5UQSsCWaw7OC0KmeySYX9J/QExqz+lCT+g1qPCK2KZ2dwKdb9qxI05quXKX
Czdjisf/3I4zUjK2ItVLCRSBfSGNNmtTtbvjQuEVu7jNspznsJ5rvgJuk1vnISjr
PoB5WhZ360zkDu5OjybCYh2g7k70kCw3SZxSjlHPHH3d1b1BovOwAs5MCStlu0Ro
IXKETciu8OnnpfY+kajIb0zdqge5073YZtiG32+VSjAKv2LrlMBLKzPtDgMRIp5/
oKKM5r5xyZ8J2O90xQaATLhSHbuDipAGzjuqhifveL4x5GM0Q4ntueZ7cKxQ4RG4
i1ps8V4AAbfJ3Kpri82N7FexZWyzoYWmgFgbiuZ6u8U670W5dyFiUY2WWCn1ihjz
tO0rqV5zCNWKryACW+syeFDTZdcsT5CrLs2trdf8rGEIagBjFG3YqDDalfhQxChA
28jqj+Dr7f8hhQVhoepY0QPWU3BYfzU7uulGubyJuBYu9ThvfgE5c6RpcRIAm3dl
nCBCnWX9mld2QwK4JdRhC1UuNo7dxLiFj3HH49GmGH6iRJ1CT/qtSzQHQTb2zaM2
NNQzVUsBRW+lXywXmp3wJcY3jGO3OB8jrXLSqwtz0GhWH1Mqrb3PjXxBKy/IsEG8
odnGgmdzU1XMP3pbQIQsZ2e/1RomPvAZic36PD1ungwWq39EaT0mpY8wl48xr7Hn
Olp7agfzdL1iqBZlqFhUeRu0HIcGaBOWzJuJ0ALfQvIZTbxlZj+9h6RFMPMjVfi8
zwVdxkpd/MnHX2NA6yz+vXaBkUf6Hq9hsG09MC3GyKfsIBeyQXgxzJuJo019wcrR
mwLhetfIhBO9dhzTdAZW5RkOoePVtYJYdKoOhzOvKJFJkDCXuPO6fC2Yn5J/1US6
KYAz3t//Pw3n2/4y4a3Uay84u4FD2EgKmAQMm1osZpaKMlA8/iuGiszqQpLOqIBW
KtRJX77n8kG3k0grt4Ug3dwGptXZaVqaVGf/nIexL9AOSJmeUDqOHwqqXfGhLYNG
aYEa0jQwp46f98zNSaDNf8+595/5JvctQIWkrk/bomQrxocB69sPUGabfDxkKhnJ
vh9q7dSd8ZggnQ9Vk26b3DN+Ya2i4GkxT/S6ngKKG5Bf7av3dSFPm/6fjpkuvkoS
8Ld1Sf2wzk+u2gXvHXEbiBl1DIyZ9vHWPUmvXvEJvidx9RLidgHbDKCWc+4pu6CB
dWcU7Om0nla5Bl0K3lx4QmaA03RX1fpMMADdOvpben/tog5gnhzL0cltKcuQRd/B
jP7OLxs6pAusTRpeczGyzNxVAqixzQZ80aorWKQ/h1WkdKv+KPxJu5NlOjsaudHK
kt1FQN6OM+9/wAuVCFybAUQAqHKAPrCAdVlsZZZFrVtgjkWeh4bfZOkn84QsZPcs
gjT4/UT+5G53ib3mB26seTrCRWXSBn8q0mVWKBJHJDiyTMaI49K6/pJEzT/SV1QS
Iz24LfOB4myMWp+xJHVTtEbIfEVmfhd2MK0uW3mooVtBP498y1pei9K8HDYxUUQm
4MWwldnuygdI/glYyGFWXl61L8VbaI9IIUrrkxTr9u2JGTg6JZ8n8zlg98XM6dZ4
BcxcdOasWHaAl8EKQDwxqtFaoYsuP5UHyQE3S/tq+vcKUIp7TP3STmOgkd06AXB1
ShgiHmqNlrSmDpCxQYoFcXv28vMS1EEjBxsAJbWw7FEeKb9tpXrv0oCBCIphV7Gv
7soF3vLa+rMriCj/SWB7QuP+o6rRR5V8PxnJ4ZjnKmqzIpr82eRFqrYEu1893l9Z
xE2Rft2LSo/tdf+tgB/eqm+W4HcG/Mkv8p50pIuQNQUINuuDfuruQfi5mOBdbmsn
iYs813xXLlajqY3itKCpDNqfAbdenynb2hgyS2TGkFhXzUrpnSVV88x87C4Y8D1R
nA+NAC1I8NR6Ah7QIal9JQDzg71k8A4y6s02OUpo9qv7+eYwvt7zem7ZSMGO40Wk
JDkZCT24NpeRt9rmkFjy6RW/6qA8dWQzsBql+LhCwBpd9amMTmM3veciHv3DUsCd
PupzDuLjaPpdj7CQ30DKcLP4KSd4293N7Kpe4sjGHCNK2xf2BGzSwC/C6mbLpcZt
R2bMoCFO0j1++F6ugPj4u0Izm8jRtSGeNQ4CrenjqLDY1jVlF866sYWZVwj2lxPu
ZoNLH39c4tmrHWz0TPLZ24nAg9mqiuWvYsCaDqCUH622XOJw1IqkJvovpvvqm3Zc
Hu6EPMQWO9cwjkva1plFyYePEeaxBpDCqOQ++hwvGqysJ/7w36L7LRFzZp2rSy8t
TEVUqjU48XewedxX04K+qGJEoCLG7qddFVl9H4nYaA5AiBbEeiKrY6+hylGeyNLf
DZvFkpmAOlcF90TpOk4ku4Jp5imhHt5IocAsBk2RjGNNd3ifMuk6ATyT3xpPdzyE
MVAfwdpYPOSJRBOv3F/URnYB9SyowjMqq3s59hIoAsWoi4wQ47vcGYNOD6cCS3kT
wQnpVJliVaKNNeDNTbA646bXhpvG8N+djJOVhjeIUNxvnqeNKsdgiytzek4cTHOE
VJlZWJRURq4BZRed9IHVyMJqvH8SA4SLmbHR/UduV/230kYAzetgRm96gQtTnQ+T
XeD4mKPBuZMUjbC2cUgC1okzC2fI5cpjUlO07BZLf5fq/8Y3jX7Ap1lSQS4rC8t/
ifApymNvWKWHMRUwt3NqQntbiCbttQrDKwk2evJf9qYSa5g81ReE4MgGmZx0DtX6
3ubfFNdj7SEUfdoeVc1KLHehIzUudgh0SSfkrjDwbCEe8F+rQdwpHKK3Hjptqhjz
3eBRY3qpDtS99QO7mc9q9VSfnnO1oCYaTSlck+5abkyUkxTn2beuVvqoFvUC+m/P
OJyE7YiDRNVf/LtZSburIL+oDE2c9E4jOgIAZA/a5J6RBWrpVHZ0pNqVUHt/E4z5
/U1/wzms9/4eQ+Yzf25Fr9u/NFUYZKuwkW9xppZ0uoZYhIP/PXpEcxzQrgKyuD6a
NLe7uf2ysP7w8/1PtnXKPVjdK1jLmIcpQtjpjs8Z2bLvpvFK2fsTEgH12cpNHh7L
eON+8OsLgtJ8cPKU05c1Y/VFg5H29rLVl3DbW4biTJMouSdhuBu9LihG9lIzmlUh
hx9eVIs7zSRYEStdBP5WhM+VDr8ThVBnsVtSuEzDIIBJRDfH8mrLFhNFDduTMshZ
kPc5GoPeyUUrVxGcaEMaDiAHV4r4kwAXgPFfll0dBP35phMC6iukkx2LuvgTjc06
vYcTN40tY3thz7UXeI5iGknxH7M1ShttXMq4emI8fRHVsZHY5MVx1c9HQDqgwpVv
pK1Hu3BwVU5g2DtvJE/pgpsPjVyGWwhQjvxHWysPlLwI32CsAEIRm3UmAO38PTWy
s7CeKH7H1n9iyRsa2GKg8K2N4r8PfLw+fwCpxEyjlydqT0wNLyBU0Xb86moymW8S
W8LyluS+5EVQnciCWEdoZdaVdiar87eTPK4kpXS/R+fJCfxVjEJJIvZJXAydFzr0
I0CYboL2azEOqY9vrsZZwcgeMYgBhz/YzkmcRghnaWu+CrDnAa9z03blQgMTnRWT
Jf7bwv0pE9VwJcX3MOuipvB7iUUoytwbgJCFbBctsTGisRo4s3bticgnFzMNT/uu
zfPC4h9G3HKvlL5x8f9+UT6pqNM9ojS3zZDH3VxbqCWiBKtgWdVNvmfDoPIBYtGo
HdiImELofWYFHlGc4lhsBxHKDGdzNQjxfm7u/5Fx/Uiya2x28RgxCFuPOllt+tfk
U6C3o4RSW9q/aiNPci9B9qHn1L2Q/o2M5juotn+B5Dzu1KEO8mcZgm4CfrYet/Nu
QaGPU6cTFwZiAfDOEUQsdxXNSpw1MMB8TIfnq/bW9RB3eKAdQSqs6HzJc8k1sYNI
pUqkFJtrbD8qzjawaK4CmF/QE0KMw8fopPgY4S9KhvcTMRUtslKnD/uowtbgGik0
xh410CJzu224sRUT6f/Z7EcYGpmwfQCtFYWil3TR7SQBqrHtvSs2t3GEgZ/7/GDY
r19aNrh6SwLNP6UvpahWrPOAuijEE9bc5I5wNWm1PMseydPPrNyRNJOipjBTl35r
pWG7HlteXL9kG0H8iEAdsZQO7liDRA/gtrKUrfsAcKlut9QyDFeyEYWOtRL/ZLZ0
kxSJs7Irc1ICX4zpvhhfIOJ7UXjGST1IWPzRPiwUkXZdjsCTt8BSNZbQtrari1bW
uJz05p4gBF0xDAy6XHGDI5XL0abRc1U+/VB2Lyb1YS512dnDSJo1kxAz1e+aucEU
TY86z6oz0MNlh7cdYw9ZdPmHt8sXuF9X6WdZNDf+EcYNiz7X6PFFly7twMmx7FUT
jwPSmLBZGajNGTYWSrOcCgzHVjxC5m18blEf1LkfEE6tJmB6V1CX+KCxeX4Xj5ql
x1XGO1/R1x0ObpM0kB17hgArFyLGOHVivGwFykuMYkH6+EFVl/sMm1ezMK042WRO
t46Y+cpWBej4W97OXnLumqSFJASWjyUzJ01imas1pA58h50tX1OelVYLuR+os2+n
njJmgHnO1ZeBOfGqBslyDZFl7MSSQNaSZNwI1Q/2Q1rcjxa4aNVC2ZztsEv4kOz6
j+8787GJuMTU7LidXFb2fBQuHQIewF8EBAhB0EBCihaf0TAwKoIG3NAddBd01bi6
/3Hd2hMzEPBuyPYr7s1mx7MtjXA/yeUuqHOESqVXojV0brfbCox6xLoKNCXoMxMv
zY9bMYWCbQrJJuj08ca+LzpB/3svJvz5VbqQlenO9F8Jk5TCMHD4zGjvxrWEcfdX
hvvdEq0NbFiKUyc2DON7fdDFLB0xAMxKpfO/aq1/cmch8SfH87fLWqhdrVDSf/hY
Ta+aKJUFeZI0FKsjfBYeGpkZZN3tH6RhCzJ9rtwvfkoOW6Ba2+p3n9FX1TNamzbK
XQrDGSz4AfwNLYuC628GqvsLZsvS/aMeKay5Zv8suWPIYJI6zccVcwi6ibooOAjx
k875xQAObsGdtwbZm+8L99ZEU2GJun7DBiTc635Z3lXfkY0C1YejOjFAJE/01byp
ykP45wy+vuEpxW8t8MD3NDLGLMglSJFNfCZQsGNSfC9bACkQjImB8Z9bu0Wwluvx
qp/NzK04aB20jYs3Lbcnzc/mJ5lRyt+L/2FYKwUaSGj7ZqQmKvXaHff4Y63k6hgM
Nxxo5Xo7t7mxftscp3kZcPJ3ikwP11eeTqsns+6qiUDhCEUVRkfMu7nLUp08jF+b
YZz3Pb83IOBjqmgb7r3j0SjTYse4FkWd6kQoblgwOPkb/GePYlTRiXz3aNRUbLUC
MXeMcarZwW9J83qUrLRkZOI92F2O3KQ4dhj6YJ0JR0xZrfpGNXy1uUNxK7TK764N
UnyUJU7gcvoRK9jRnR+8+YQrBe907YfJsmU14+zz6g+f1yQKxa++CvPI+77a61Ko
lLZVVYk8NAMziDmiP29i/sckbA3358wBb+8unnR0CMkjruZTQhtXW0RqL5/Fnkvn
uah8HgUO+moJ+6z6WvQJ0TgXzQphL22cTcm0Xpk1Xdn5Y+C5VGFfjlLdIhHck9fk
tHQmfoQ9Sq9ly1Ezw4ir0sdJpCzqfqNuCmn9MxUgylkiryg6v7AHrC4NFjNCGyzK
c8vw/z6DC8WSafqqyop+DK2pRBuPhyUGTKY3ZZho78o6f8KpKhQQamdnbp2T1t2u
XL7rM2byB0sgYy+sjdrX5silzFrj8NHeW8iDhCVrQAv/VH6Pnx0WIehktb1hQXYJ
VsnC6+p7F/KAW4qT7FxzNyJv2HyXLdyRjhizyvsl7B6euk3MfLpD25WtanV9Sz5y
Te7Bic1m8kb7ZoBZNHuxtkK2vJwTY6vMO+ZoF+Ffigd1Zh1o8XevPKcen+mW6CYM
qFGjnGKT/jN4FZUPVjMJAZdrZwWSHDkv45L2hqgWqo5vJ4j5oHZaU1xGm+Y0AXvp
vz/yMjK6SqLNYfuXrUaznEE7OB55yxG98Ux5vMwFbRgKgeTv4axvTXz0JLalkdJx
vIRrWr/KhsZGe/5JkPaGNEcyGjQNeip9Q6ta5VPhf2zJgje4b3usVJjpootI23Pk
dxAmYquq3mUVk50SjyEpZ3sQB4tXwSHIwWo2aCGonSTjq/gEosp1y/1lEwmdYzCf
EfFI6sYKlvPythOt6HCbhziC4u83iNluaZAOWNS9V93pnPQGKgYQ0i+C2NLsPy0V
5tadVg0R6Jxi5g0VqDYkcol67n7haenL86wJkgxtqGVAtTcYpgapaKqmdWPIvejX
iupKVQHbCdzOqDnqN3G8IwXSPwzVMx1fI29WMhdr8Nm/u3NNC3QmGpqS2Q2/CjZg
z/TWX59yfKr0VpC56CroOJIbQJPnAp5kLUMZdmF7kVKet3VeMtPTNUVWqwPuvvwf
9+LreXVDXF40siyUNsnU0xb2oYu766f8WxVkxif21u6QexUMZoo4HHyRn7+GcXtG
E9klP1qA7hPGV2K7Bma+UMTu/Oo3onWQN6VSe7YMeH9w6ToQG2pcFLjzTCt/UI/r
b13wpMfUOhVqyaM1qRM6xseGn/jdcKNIa3zChnSYbeDvRS4Wkf9UM6rl8AttyPYi
L0zc8rM8xGWaX4CsH2soVzTEAF6MTGyXJTYttdGu4Kaz91LG5zbbDhF/g3JBR9Z9
JvGd8bCkcDqwMc6DGwhSJEqnTWUTHtnNjJ7/cwZUzhuVW02lfFda68FTYDhCUGDA
IAwGkaGebVxYsVEyyJ9xtFQ7cD/skx4uGCRJIVjGmt2J8z0wzboiNRjdobP/TGK0
xd/IVnSyieB4dYhW1NlBavgSMjbcGJEICIPIxxIRCKgC5/MpEKaINzt6kYF6juog
yOgaYIbk+Xc2nfsxoVk58ArvPQu5ZK/aPVTi/GRLbbofhc5XKF9rQjgwfGd7Bxjm
u6zTl1RaP3zL9T6ljdosLY5RPN+yRYdU9Me8BB978g8FWK4eT+jznIlnhm2LAP3T
Nzmi1zWarkoVEKkMFI5VShtpL/mhOWiw54CLt6dO2KrAcu6wExfe6H5vCKPF/6pU
QG7iva5zblBvsRTIxnEonmpHk56iWqoPeuQbaVEkWpjC8mxQke1RQxXnNtJMTaly
6fKaKmIPsAdjufDW3nI0pEOD3G1CvTTj+/13CGp3LjE7eZTh9EPMkT2hv8RJ2MUy
Ht2+YLIJlaQt6Q4Uj6nLTTQ+yIPrjAr+Fc0+hNv27y9zxCvQOVpu9IhtnJCcNkVU
QRU6LPYKkOlRqpqP9F4tebzsAVMzIeaWEl1CMp934cQRAK6zHrh9t7W2yylDRycp
TDafaqbFtDYdwJq4e5iLj5Xm0xCc4ObcUJ8GRmkYqpU/XWWSgiXrfEW0HjXbOJM2
2qeFEEfl+H2Nf/D+zWs9Bfgzdv8jIA06tGQ+LNg1GoNKJTtol8y58UaDCH/MKZQt
I+uvFbXd5ZSzJ+S0+heIuRa/sDHlicw+qkStNXGGrFc3a/JcbiBq9PslvJWAiTas
c9HN52e8FgY/9bDgjPDSHouAGxe73axXEaDPfJbs4N0ilZg5dCC9nT+pzspXO5IX
HnzwxWb7q7sfa6fQGuVujrpLYmnGXtPJJjcr2HOtGo0KuA5cFdSRf+Hbmz/i8+KD
eV95eHamcmcmFANKCZ0yGEI+8XHNfrPbFqZkqasyHb0D2aoLn8W9QXdnRsC+DhlW
KEnX3I9NYGeto5pTo/gf4XUfkop0+ZyTXFVttRPfZ3txHBa8PY0l/Lh6CiHXSUsA
wgrbFIX4MSoEZQNlFNK/Y/7jGic1TYSnTaBjNt9/E0F2Q9SXc0ZN42+9kd1bK5KV
rTRWXVDzcyckP7xcSLWwcDlEr3+kjcYOA+IwQXcKL9JP/QUC8CbzGEM2XkZDzqs9
r+Cvdgf9uThOPxrpehcNrx6ljW+VFk4c0ZRG8JxlfJTJfdzWr4avfpmHSZFChTsO
rjvO+c2oJSwVKEqNDXwg0IGBTjUlA8bSIgOeHS7MWoY6sm0oVKZ+pz6jai6Av0BF
fYohCiR2CyzfmrJK+oc5oCL35lliXj1pXMH/VNN6s86aesmYWurEDNDQNOcMjbIb
tTbLorySC7OKJnNXwJ81eRV1txseYjtY+2hPhXCsWiR089F6rPh4rO2F0OTLxSKK
mrQrDlLlq/MpiKC6uvwiZNtvnrQwSBNw6eB0a6Ox3xUc/R5rZTE0T5BSIGdfAF1a
HMUP9HmtURIsEgBNSLSZJtndxhJsoWCsBxKDqQMfQKOMOM4APZA4r+Jm0tCLiK87
u+oENWGXoY+og24AW42fXJ/O7pwV0bwreZ1M5gdWyf5rnxAP/jyxvpny2XtWhh+F
vUjd1d1ZtdBlZVPqWKwhAmbNCVFOVBYnbs5EwQxZ1oUGmnccfl9FlSlWjDmxTbyk
1LoI7LTIsXgwi1z4lhnlfToX9iX+DeNmnMU+GnAt4cpsP1bE4uJF6IydmihDDR9Q
HY5uHEqdUCvRAt2j8euSDHULBZeaBNHOryDaS3xhqbpFjaurWFZPMh+ZCN2qAi/j
5DjDgCNJeIRVqyOnWASSAoFflcf4K+7N+5If0ikMeB+j8egGYe0ElHvU3u3fjUsf
KJn8SPQA1QLkHxVErTnHJs4C3QS7Aenagp6pQTrF5PnmBdFdVgnRfQq3dbEYbkvq
daWVYoHPKbBpL9BdGwTiD6L7sn+xTpdrV8/nFzHstWnVm2fBKUjO0/fBB9AumM6p
tOs43urIDvRWcchGW3snhKqKcJjKADRPwp9HpczDzPOT7XRCx/b2XvnvZl6cNZo3
pjfb/mfaXjU0YiIb+hYaUxVMO1P/DxzAiQb0SUphA2QsPWoYRv/vCRpGhUJerRjP
bZKTJS4sJbprQyNs0wHDOc9hptazYbPi+yz5SW3VlWkIJZnnMyXAevNQXtKR3Gpv
XhNvwSz3PqWUvVA70ZUzrWWg6zc/xfRqkMh8zyTfAB3W3q6p9hSy9N60hoBYI/FI
Et44QUE3V5ueTBiLMRiCzvDj/5T/keMa37LzsBZrT/8wMkinDPW40v2WN8/T411a
XOkQQOcsHcq1jwG8ggSQ+A2oy8iy5ZQn2SKNLpipZYzb815UZ/QnJn0kcHt7ldrZ
qpko4zBtYh6uQ3t96TBOAsrND5Di8b2hkQIqBLirxvQNN0aMzRnIvLIKVDd/Lqlr
lZFcmimuMZAzEp5FHPITZfpzoa9+6jY/wP5gbFD4inKOKCqGua9r9IZ5H5zjBHwI
TjKWA0lk4o4+SacDM5VloBBrrh+anddBemEin3t8T9pvy3UYddeQeu4/RafhAwlz
Ce3G3qCR66l9sBb8Cd4lkfa6eIlnBPp4wGYHYOluStAFo703NLwnhnrfIDjBJAAd
cs9IiriNAgt28cqjZlkpBKwzdUGd9vOAD844qWUh+g+z0OHN4P4cZ9Nz7uJCeX0Y
iJMhpZT1rP5dogAK1NEK+1GakvCa8/TxDiR7YIXDub4YnuFOnqUtzJ0Xx6GRL5s/
ALCCZHhbXriKlJRULrgC38gxwByxZyso6qTwJLtGzkSWQedNDDU66723StiXoIdm
inkJPe0TgKZwDPlWFipIJ00tjyXf7bQJRs19K9bOZVOoYhMJ5WOA8R3NPAz88Drh
m4ZqQQtXtUCnjCoQdq7+FOPr/rAIO7eJGc7ELpkeixBEcUcbz/X9RmPIdeuCS2Yz
VzxZsmE+/UY0Zp3frjbted1EZf+OGtGUu1jkbu7mocfXnIcptZuHEpx8hdKczVUh
UjJJiPwh0ADnzgl/ocvq8NirU1IHy+OEUODEPJGR0l0P6DgOT2KhcpQi3zHomy3w
UflyTtXVcBOHgm+6PB+UmtwLmdnBMkdxVyC56nR8T6l4TzLI2HDJ3nQW+mNDDpfG
8GPlngebjnHzJtTHi3F9sIT0Yug4BTDS0MuESvoIPKt+zgvztuOktyKVyv7ceUmm
DtDSKXXnJFrjF/VK5+kAJzL2LuLEDUypUJ6xwVZGCkt7wzFD9csbLtIY59PI4LBE
VBD8gpQ4Pcw5k3hd/vqZ2P7zzyuPHVVwehYZeTppGUCKezvStIBVTDW/dZ7RC0/t
iL50OK8igFhP3ZMxflNMVwbGytSKbMn/QJL4NL+U+BFA5Qpf1T7EhTq5r+C/pJMi
ZBpIrtXi7sMz6iC/B6DpfeubAQZH15lWZAGZqUipawlIYOKRZeRHeiGcAfiRjnbd
3mc8H/PVzaiBShUD4CPeai+++AxIzhwkFX9+oHP0Mw14TxHwwOeSoAcShJ24YrLW
Jeg+45FDaKzhpJeInMfQwI1pHyYpIoxRPnv+GsHdNz35xhIU9N1hCYHUst0nLAxX
3Yrj2Aqslk39r/IJ0/L1P361uNPX39d5KD7jVO2WOo5y5Npa7EQey4MtoeEA0Vm4
WBMS/7LjB19mTKNZkH2R+caeADqXx/Tpgz09ulQ6YJOrzhRC6inwnkMXX7pF5xNV
8uhvN5IKgqQi9SkzofkbU2qHaWwVvnZwCwl+3RoOaR24MnE3RYQekkediJjMEum+
eylbl+NbllnO8RLOn43XY6ERvxyoikquutKh+KCYvwwQxvsBF7AUuJlv6xA1k3iT
30Nz+gV8OdVES9qwL0JJTbUu/8L7+ha2wkAqn3QlczvrJYdrVMdWUQOiXnHznosQ
bFANZ4GSUwXJKjaP1yaFDYzIP9dSuTRSBueT2kR9MPREjce14fr4YGOjCjVNbIn8
qeXAmvG3BXlzwNbZSoVLD0OuK3yQX2mPVY4X34z8n6cgDTpkmv/l70tcGl9c1FsE
A4VESMkXogibgfSC8ZqKzzVSuYPfgCbFp+CtpkK3tCtYbdaYI5p4OGDFV7EiDHYP
t+YPmWHqBATzBvnB0BC7KPxW0ggjAitB/7ONoM2hFnkRhSKg9AZR/MTAWTAbsfm+
7YMoL9u8hFuRp5/W12eKWj3T5QeMK7eLKChbJZ7Ja3vdrG2V9O7oS3ofmrqpfI4n
rNoBNgT5bgik6doV26SFjxPy8BwUCBhRsxx5XWpHBqJwknPoVuRoJ/0fIz7tFSZ5
CqepaFe0x9rSipkL4HZ2PQs9jCblulFC7QZ1U3VJgHzNTGxDfH0sAk+fLaX726GP
iDzv390IIKMfteN3Y58Kjbg3xGKKEuIOCG2HnFdP6Ieh4FVBMRJXCtGQQxLEIM9T
HDJFrJCZVyx+0J9HnHPvx2GMGSwlLAqDo4+/GqeGv83ZNMUSKRAY3dN04OFUctDp
buidrur5fSO4rkpI5w8G/0BAFsJ26PzYLufOQtZw8DHJyec39PWoYlH6XNZO8nnr
wZ9Vex3BPpKjr/HMxHd6o+m7eaq3g03k+fD4ynzHmPAeWrmSDuxQ1HoO6iXCzXVp
IgveZI5MgJWql5BPO7ZkBkHVjYilWUQfpv0VMo/h0ZoX4qwop2dMjbD9w9rxnqfn
X/rOSqmgZOFzaR0fED2gZdUqYfxfeWuw61ALekh1VNFuG3uFTN17ElHQg98dIC5s
d4cVpK4EY328br7IdOdP40EYLDx5YNf0hs237rn0KKYioFKZIUZgyYGCJXlmYO5a
2ajkLbRDgUpEiqDw/e50c8Dx4gEvq2pmEAkInM581ayN8sFOqxeFb3DKgsbN53a4
OYBsLZLFEP45cGmfAlUZ/pI91SQl7Je+2h9GZpBjwgGMvQA+LCxYtaN2OvcQxpS9
SFONzMmifm0D7O/gWNu3EsheteMDt3xtmtdGfgjHd35RaVDMvdZu51zrFhPDxhHv
0z4n5iEDwLlGY3QsS0HLiwrGAoRlr4feqaqwsGFdx02jLN4VWrQNiPgpA+ajDlAo
3A+Qt7/X5P1riTOZrfxhNgQ1g4nx0uehOcugxds7VWdB5g9hMjM1Z6nCLeZPWFN3
CUFc49szVkQLbmJRGNeBORsFNRMpycg5dtGlL5Yr7sIQ39oGsGqAp1wVCkdHhlDU
J//w+04sFoL3tIulCAzKMSd3SkSlkdhg0PfzAxDBjkqaW88DmPKN6KgVr58asvaj
+PYy9/yjDHb38V360kZz54yfuQUePWLpKS2sEl3BwPL6+DhdrmuL4HTdXZ2XUdX+
jfdkQ3PyMdhiOchz9oHcjypZaCJnm3Ne5uzYIUIQ9RqKxD/98VkrAn7qw7xLumht
3Zwj7isS3jqk6gy6kZ+RUhXx9K86JCuPyLD3Bw30C2nsRRNta2AfG+twHqSHtcJO
oSXEe+jwjnciqjpJoN7xGtzcrJHaWFhz0Fr1rmOn0WcgjEP9V5RA8UdI+MaQb/cc
m01l2RcBPqNRVHDITdvb7GdtX6e6UCBK9E/l1KlQ/HOYSjZqXKuIv5f72XeBZehd
Ek/VdpSSw/VgSQQNzJiBw3GX+D9S3gUXt0IWSzlxbhw62okBlyOM5G0KEKH54qs7
X/C3odHYbAJX/JkOGhszbYabezkLh+S3NiEpcq2BlS/QBe7bUMqFK2uX90JJVgZF
GRx5ihzqwN5Dl6SAFQ1IqFlv6/cFuntVXNrSWqpnyhp5YgTh67zE4z/f1GIozI0z
age+ArG0Lofn+Go4FKIwL6GoItIOHFnJ/UyawYaCNxIXEo9g2aPhE7wiuIVGCMZn
t8W9JN6Sloz+ZHUxmDC1C+NUC0VStQHxpIKsyA0VlVjYyaam3Uiy9HMX5BqHG0Tr
ZivS/3TpBe8vluDxrPblN6IPdiWszMmSnzfZq6KMSYwYIAkolHQxeOEP0YE046S2
pMrK7NyusmeC4CBq6Xm9T5nLPFKBTBHtoWyAfpxbGTo4PhBf809y9OxIp/VJ0MuX
WyMxUK794wxMq6oH0pyo+GyyHtG7j6OPZl0I+WsU2PQEtALly/8ce+aY3woPdf7m
QJTrP0hsAlq5RgdUf47X0oE+kmGa14hGsztMcSnbFgnfEzIdScGsBqmEVJIkTlbw
pychigcgaA6CG//wyxDSuHtRRroTKlF8MQ1RO1XQkAuZaNTo3AypkN6QAoDwKIZi
vM6NsEq4Op6+GlHRC4MTzvmmm/vm6EQQbzHcmVVv8QRFJkV/lIEhiK2pFWfmh9zE
0+Hs2jCl1W1PTHByYs8C5rRnkWBJDMj+UREvBeN17ZGUaVE2wZaeJNBhnGaD8qvT
2lKT4j1T7wYCkdJfBc+Ay5YYmZvqK9lRnV9+9iT9axcF5G5QVfV28qOYYIiM3QnF
7IFTFekJ93jbjDEDFosZ/UYXuFLNIu2uo2g2ik1AkIXhWP9RxWOnu4FBMsrsCHUb
XsGsra/lIkER52+SzkchfQIvt9/Sjrb+wApZIylM1PZjzI8hwKwV3h93Lx3Tq4xf
OQRfnWSReFKwearB8zmlvHYO9LVOTvpuNbDkZ5GMbqvix7a4uMYzPPArVwPGBbgy
pWsklh3Wwcrx9gqC3yE7DmxjallA04xYPI/687zsl0IlJtHxZUaP7Z+BmMvopWEV
ASzv0VLU15LOqTd699evKxNpvRnKqWvDjVeEpLzbWQB4YZPeuFDB39nGX5J6ikuk
2YT1AVAQXKDYUDJGNcizkm4yP4zbWzLBmUsP6z0QocuoJz8XXiV2eL1cT573xtrc
Mb8ctn1TfosifOz3D7nkoLGUxRwflWGkptyrF9FKBYSI6kbxQuiQk5AQ36mZb1KP
zAxiJsHefoNfCt29oAtE4KR6e/AixUphDQ4uLNWn2SY2tuSyUgQeGDieduPokrZE
SkrDQNoJFowNnyXYJ+dHyAmEDqNM2oMwMSqibW1osJifDzHC8UbtZ5JVr1Pqzhgg
yNCae69RIS0sXYrAge0o8RXuAW3+cPguqBq63609c1FLmCOmH0+nyHTFODaR6IKa
j6XTRkkIkA1oqwvqm1X+ikK99JDPR0NtqC1cT/i7b8+J+qvFxnLD3Zog3grBKJrs
tQ5Bwgx1UZQT4Dj5YyRZCwyKb7LDciG/LrYgJ4MLCJOYqijuif3RLJXE1Cl+WDxg
O4JfGMKHCx7IVy2vsULfD3KtclK9jJkuDYJT0KQiDmy1vrd6NRs1csbVuGW6vJ/k
efBFzHM9O27OPpSTW4xL+VyZCegcsi+8wVGjgnDSgN1HbLsfG8TY3HIzMphvc3dj
iLAcX3p4OD7sNHUUst7RRNxz8VfTMoXoCBwvehrdopVPMcOImeKImFURMUmDcTk7
j0nFBaDIopEhpnPYsSE8+sHNfOzY5FJiimNWNBokYZYPC5ZBG77jSQOLMy/Mp/Rn
kNC4OZQ6bWhI5/HNV8g0ac+4du9fYYqx2HPFZQ8tfr/6ZufvbB6omZZ89dq63Lpd
szgpEaaPGPV6SLfnRu2ev81HNLB5aoVwBH3VYfInBxO7o3Qa85ZbdweRHvmsedJc
H2zDhZZivcX24fn9insr8fFHJR9UntZkEdFRqDWU/599BZK+S2ABhPkNEu/qdoD8
Jf7G1kNk2OEky9uG75wWIpuXqGeRrACKADtpGddxQKkjFRmg1+C4K/sAt4UNemyR
Ewhc7mWPigSHrmU28tBoF6h7bWW4/avf0SCUuJQhBL8B+QVq+N0mFHFypoEH+7Id
EOAn6kRcFWQ/TVeRda//iTEa4qbT4sLxcNUBEsIJ3PJ/8kUkyDXq6zMC3Obmu4RF
y7RwQ8Qb0zp54GkvzAdrdnlZ0qyAVp84CQStKQLh3sTSDIg09qZYjCCYLXUjyeEC
EkhVPXuuKPWSxOcBlxFnE5fnp3g1riWuRvHq8GZ9+Ltrye0cE89uxxUccpL1RGDJ
0bt5+6ldoetNXJkbXOud00VxrGVzt9PX/4Jz4QxGK7FfG+EBeCtJtfVSAEms8j+r
cOCHUXoK2v6JVxE76IbPKTiBSid7dyrx7Uxc3ZXr2wdDBRTcwLn6OkBCuX5+v4JS
811i7ewn6SSMtl0uCEkNXhpOsh7W7ECosJsNXBvuObX0hhzNB0H5fRa8D3p/qLGZ
bGmzrBeE00bXK89HB0Kz3iJgbmvanfIxcUismR5cpG94Lg+B6kmbp5cJOYR01BA3
1cfD4X/HgER/hpb5gNWUUNx+nV4N5xZmfDXGz+2N1Q5d54Yh57GdGV3aIvISMe0s
tGJE1mSVRTCOcB8pxZ3s0m70+FadpltvLy77Vi/uQbQjD+10hmI2S+rvJxAYQ/9g
PX3xT9B+b/0fHjqK79BLCl1ZtoLmRESmgC2vtnTmkbUJF2b8J8xL1tqKoyTU6VKz
gJVDJ6C7Mjkmfh6ww5xnr9UIdspg2G76g35jCpmt93xqjtCB+OYdvsVE4VNRVQLe
9BwLNRvxIqXM9fS7F4D0upAicO5ZdL/yhMyCvT1J9e124+C89qdER5GVJF+gNXXM
9pEd5Iep9IGZ2gx1gbNj6HjNuGbPypaiau3S5qa4cXM/qLsghLru8g9aNhgY4Pnc
KNnxpYsgA+0LgCtWn7JvDrfvNgY+TvDnMEgKagT+ymJjrx+HGEN9EllN8pnVEVkQ
K2CotD3DQjLHTGzFhBULPUJiR7DhyEqom60tBiAPzTkE3PBZPAO5kKbGhvvrcgBQ
TvQMhpuJoTF1UZaTiqC8IPngYBLJpJpJYo5LVKuoPsZh8lC4gHCSJYrSfBeyfGr2
8488g2mvPqFqi/imuKDWgIV1Jgr59jYUHV1mp2rHk1r6Ha/2u6mZ9POvY06f9MRh
PTvff8VRUiSZu8ZmYcMXmereCVt66Gn1Ok8R1RfyANMAmv7b+/YlIxkH0boOsMlB
FzalMgFYZDPzTBnJR6JEPNdNmTIGCtFPKuW0p+X5HACtmHayA5qcr/yaDa6MVKQx
qswVor0a5iuXr7bB5A/6+KmcrGZQKY8KBfnVkqxNkzQzTAkP6jwC+VmBYsDgvUBn
fyXKK5ySGL/RqBXNEykBLynD1E2JRU5BnJrJH5xkCkAWN7ngDX1eYKHuDdpVYXIr
+/JwOeCsQMVPR4N33mx2VRur2lD49Ov+CFUV5iOZy+JSO4ghZq8uIva8JfmtRodF
6q/+GVkzIY+K9mGKQUrraAJGwQMplIpah+Fnd828PMGJCgdbWe7KwlsHcvsZdg5p
fWpV4vPBLvGX2x//9RS0/vGA3f/o5l3+RjfIJ68T5W65d7ffm31ssykj/2RqX087
t6snZuoArNVIToJhnltWIE1mFtsXnLljyOiI1H44fuSWhLipucO+HG3XjAn3jLw5
A4yKaUb+0xqx/4Ya0e9hnBey6Z9LCCumCfDtYJi3yHV0UFwM3LRzYondk+5x/rQB
g7I7IIZodi1nlBCUpIqj9IDauESNQdwdGvvhAHDG1lYrp/HG5nxg5Jk+jmEJUmYB
ttfA2onH691oWqOI7b1CAlBpWXfu4JVKz2oM9H4cMx+0Jgm1JCCpkgg/2dY5hDri
SMzbQWAcB59N3hhXlEilKJq/KSaoNMfOkdwIJSu5j5jwM6zbmhS7VdL2UHJeHRKZ
Mn9kB83wUB47PElPYskzPfsyujeaee9XnYTCJr0lvgAllmphBcHddPHYTKwikVcg
wCMCare0rvLRrlFyUqUL9NJ3OLO2jxeYcu2VETlEguiWtIGOB6ikJee6xQ3x0kW2
jg06KysDedp0AaqSj69VndMCYKd2LJPGtOS1838kvBH2UDPWdRoIEwUYIucPFHgQ
jI+IqxBZTzx7A6p57kwmzMIJurnMQhARsHJql+RrJ3kLPkZL4r+ahX8TbMCkoHfq
JENQm8uOw9Ya60Q5rzuasEez/CLSqW2DDd8rSB2PhUrv3RmvB/K1kFUujM3OL64w
gSnB99LlPn394cvyD+3vUsavJMhsl5zogmJibtV9k2Ta26YQB2hmyBf8LQ/DgZB9
TNNeo2avdnMQtZMF4i+VOC4/VH9GADkXT1z6C5JKsqUXPz1MsGW6lHElaChuL1n2
3kMqyPjqhUGjaVwX5HhUennvA4k0P5K96j6PecoSxWwoAnt2LtZID9Pach2WJwvK
A0PGV8Udq/7qP/kEZlvy+BMRgHQiKsJ9JVoL/5QSkXFQUB2Z0/gK9IzuAtPsaYFP
nmIxa+QIC9JBHdUbzsO6G4WB05JRKikUraVYccnuSEX/PdY0k6jERs3cHBZNhNhk
F/73F1StOqg+QTN8ScRpQBN9dx/AHie7BZGvXEn+cEKOTzdkCgrUxv7Yktj6LchJ
m/zBVERGrd9ujq+LY1ZvM4UdSOtOMFKajdU7MuMQV8LC2vF9Enzwk7SueykEgTpr
g7NIi04bG96CHCHpEcZIKM40Vu9E003+14Et+/u3HpR63PACr4RkpMREHP/V7X3c
Uxtb0zb21hcW2FEPpwvS9TSEn8K50iD5eG9p/dotMH1XsVoXEwP2kubi2r+CO5Zb
bB1ajQOBQlN1Oqu4joIc7piYvsmywhKnaxlNpzjnoPUbuuHy4XpYR/UKghqUtbGA
rY/oy1F9edZqo4MI0zjW2NCnAN4rgtXZWZzDS/ZIBCPUN9Od2V3QykqL0ZD+fGES
94B+w/4v/Qy2P8yIv4yLH5KGrbrkMu5mFnEuSeVLpV8TzsAiXP86PqvpzzIN245M
ursWltk46AaNSWTFYgd52TR4q8YF+B9a5MMWrCZ+Kl0btfQpRISJmRNGDds6eC/F
Edngz6WplgDWrwEzEGGu5MSAmz6U7sxfJF+efGfGCG/dvLfq3sgRFkO3wahXTLEk
fWCkfqH65SqFWo8m9vwV5OkgbqSH/6CO0atGajS5DUUotwjs7obqb4GSeceRs96L
u/iMhkvH0wPbY2T8umQy+sDv8g0BpnoXaY/VlH4aBkgUgVxQNUMQhwD0jM4nQbGV
dGscVhkejJVJ2Bdxg50rKbtGa/GiNgR8JP2BbmRfGPusnwIfioi5atMUvL4hBC+k
96ZPOpMZYgHaXYPjpqAmookqIzrrz0XTT59ki4vzAdjjY17H+DKrv6HRS6KRHTgh
taxtSga1rHQsOFh63YaViQHIEFigEFZhyKFUB0WoTdxh1k7DiuZNvrVLB3+0tRxN
sEOvy35WSoldhPObPLrnJbwolK94mnx4F08v+OtrySbWPWtqotj63q/BzO3iKmo1
HxnJGBgDes9yuZIWPIrsxJFOi+R0AS7+v8YQaIZnWcv0a9DEl535AcZwGQswYRG7
As0gMiqYh1TtIYzivYQ0dcWcrK1ES/86rIm3EFzVOlx13d+Uy6AamF5uOFDimJqt
KMSA9V5tb9/IhZryMZ19wLfK1I567B+CURcWaECNl3tdP7szdXwLqlXIyN8Ix1Is
nl7Ay4PbhqmNhQbiBmukwlWxjxIpB3SpxYQGLUagJF9ii5UfR0oln1LoDUL6LA3Z
hTwhKSk8GHU8bD0Yxc8+czQ1XQqLqZmtO3i04B1UguPrywO9ap2Hvlg2/azZAjxu
r8MQ2sdN97XJQyQ6S9uYZgGyPf2s3J3VFSiUSVkE5OuhOkkGCHtUI99tIqH+oeSu
xh+J2MonXK/TaLtbUPW7CjmE3GN78HZ27ZT1MydbuMAYsBiOZcaaA8b8W5jbPSbp
Ab/tKdjE7PPvMS5mD2QTy+KW2VpeqD1TdRwIOAyCtkguUsSX8lRostsAEsnTuhl+
/lnWBRHjgcAOUs3peFcXhyxAYElV+dAnkV0dTb/EOlO1q0GtEaIR3eYj3U5R2cXH
vAQb2hiTilmH4DmjlApzcZU50x0nzAjlX53cZ6gLHGp5+MC2gjvGvtJyrMJd6a95
RJEYS3BL/497wiYmSE4NnXyLkxGN+3kSckEhxurhCqAWqnb1zB5nSGVmt1IHo/tC
tnEYf7jx7hez/k//XerLY0NMaAwIwYqn8f+Bi48Mp09e2Bk6CEjHdkD4TORjby0f
qS7kBN1b/mJFlzeWt0yOPs6wu0EY7wtFjcREE+2DEBtnomag4gw6YXnVKO0YBEdL
rQBYxSCf28SUuk9Hlp+wTXt2ICFyKNZZVt3DPREgEQV3A6cDZyXn4qI5cQ7oY+yf
D9lYP131FU1KH3RUjPCmR2WlF/wpXVBD/6M8SZlNnQBunsDZi4AxdbWIAR9LViod
JnWMtr4r8j1cygOtoEP8IasI0Na0OSQPsTK6P9eJCQB8CNa6ITVi3+zyDex17gF5
XtkV29KIDVBEFxK/iDhbzoDdwxBNSyJ2dZPyMdk2kE9C8m/lDjRBKHnysIDGEnpP
758EmmTJYxCTIOS0pnUpyQjtLn3nACJJ54jKCj9e538WprevaYvw1lrD4iSIotb8
2k4cssYchMjzLNuqLVVS9+yjtCnYNFsZdf/4tMH4gZTpCOcrg3uOy+5ApnFLzhAL
/rk2tBuCIwEBMzTviBMn4fRjXhGFsqayLsi6LRiHbf1++pMMQs1Hqr5X6xrjpgIv
Y08/Bwlu//Khr2ZtKvkw8EWE6vP+frpaVoRXuH/WuhLF+0EF5tRMPhb+VbXV9++Q
p+O89IC1PAbIVgVXUZWL5D72OJT2XgbYnuMNEaaS3YZIcHp5C/tyE5ATHgG0e/T8
6JxxzjrrSzYNya5xE9+Wt0k5YGl00F54Qc1YZgLZmEyCADiu5Zm2jOkdHOwvxCkY
U41G5HeAzwSGfBv2R3zEonp/+tiF9yvrJ7VPrXJWF71m6Z9wQ0DPeGMEFGJd5/HU
2Dmoj5qrphYABxh1JPqL2Hx0krKJ64huGev64gOGaCL9HNDmJZLgbXMPHzwlLrQT
7W55NOHwxI2sFqI76/ym9TERTQn05XwqwhQLM0lkdLDF3886lT4vZNYNJqOIiaeA
Fq/UhTQHKURuJEpZosEPbsutlmWJwctdv0Pi6DoCVjpSqvQvQHXPdlvz0Um5SvYr
/OqMGE+DU60HFnp7tHtnmOftj4y1EmYYNg+mTFSBgxcaE7/xHiDbAXIpsV1f6lUu
oUJzQXPOt34FWs+w7of+vITBSD6BRQ16NlHco+EFlO8JHaYLpmkI6KDHYW3f/Jw0
FsHbQ4bDKi8OVJhK4gLpiqPxM3nl44CSWPgy8ftNmvhHEVnRt8khx3jPSIwY6Efn
diOPm7Jph6I2mKVID/deAtsViCcbZfmkCxW8lr35dF+KulMl+uZPB/4xNX1WsaxP
1VoiFXZpEXn84vgNZfwFQDxO4P6h8VTtJ+C7yaUnu4TEj/0357zWXQ5EvcVxnJo6
M8F4dUOc5pMJIla2DGC6RH/rPwFWJd3gRq95PAQNp7ZtKwgsRPJrReSYBGuOQUUC
DGugsRMegM6Hn6UhffIAzPg0dpuIS6uwlcUGCaWlJyfef9QwDr7wM5asVtygUcRk
T1JFc6mSZMJWXD2fwy6eQesWKSZ1mW5b/tfTp5MWRNdoDJ1wVxEWj5L3L7Q+oXhy
es88gPUv7OIiIA7gWX8pI50UMcLrHQx+Dv8fi6P+L9xTmeRhVCBYGFAeXX/sr8gM
ifdOEwVGCGbPlBsBfyzV57BEaiusxDF0PmKX3H8ZE9+HKRL2TJOznCLR4M+1ltJ7
Y/OhRyr7TKIWAb/fgySvBGWlOP1bKJ9neONSnYfEL3ZRRP4aIL1Pa/A9y32WL3x1
XMDw8h9FxmYZ+Tsx0dNinZHpLPBan5vdXeXd+oQisphzDwYWJHpcfSqVHTz6Kqwv
ZZkXVPfpM6uKHvAD5hRb4xW1m1isrrB7+vXCb3QVh2ScaMen+QAtQ1Ts33pkLjb6
Ha/CdGDvC+Iq6oZHemq/ZJJida3zp4pwlAWbT9DaGB0HN0tPsm5Wwt3hRLDGFlAG
KHE0YdkrS42qvATNnqIw8/chwpWR6Epcr5t1wP/3ElTe7NJ6RgLVr0a3NBWw24os
aPlnwJvdHFCbCHpl+2WYTXQ466JuNwxAAdezgKslQpSxXSvcnp1niNSrNrL3Habv
uBGVpx0gQD862HdPEDY+o2gAyc1FFbpYhaqWOA2Hr1xeVAUK1/gaSP2qFX5SppmT
blzdG3hTwUKQAdT0vstHNtuUqgpMIk/RDVh4B48Wssp+W0Xss8bz0Wk1h2dsFKI7
qWDRgvcpWdU7f3FH00DWCgismxAua/X/hZCoym7JgBbsg8WPnSYc/Lm1P+SorY+j
Dq8Kjccg5mvf+IT55NDs6udGyUmilXcdHnwLxqjRZaX4zbJ+1hMTGDY0A9mPSjxO
MuL/nHfnr5dCasIDgbLn+D0ObgadnDaj9qU8OkTvdMAPYshd69HtMXiWZrsiFXhD
hG5B31yWqPXBTS4sTEYZqMbaI4LIKhSwq5ODH4+hIOE7AerHJR8GGy+zyZZk6fyZ
cdtvN4YKUNPPC+qOXY5b0LlaFsSLnNpSCKftUjMBbqZQaHbOMy9mSP1t2AKIjrZ4
VMc9sX86YWBrcBMP9U4E+roSd3cmcDPQFqelkeaUdyjyYBbbC5IawaVmiQvmnvTA
iBfVR8UapSFzFnSvE9DthZrujk1Ii1dVoDaZEgj1zEKWnJ/lZ0FIbiYW5ac5Zg4x
0D7toQww4AJmzDe7bVGg5oq/uOh07Xyu5Rkxj0gWsrgJ81lavm9U7yTODK/+VbIu
p7e1FqS5ka5Q8ZSMXkBcqsqcZ/mfBJkXoRFIPWSmJtFbFBq0sfWSW9M6pEKaTQiJ
+D2PWf3uOcCn5QCi7O8IJ2t0SqKuxrQ63c58sYTW03E1wSaAO7Wy6e7LQ0qQz4KE
lZWKSUGYLThH6YmgFbFduPE5kUMLmt7bNF/W8k8U6HX06UejMxw6hWvNWc+1ykxL
ef9S4+hMCn2kz10tITa3ei4ayOEKPInGfMYZP73L+SXiCCf+gq59CdJPMeSBnNP7
nC30gFBuHKrTAIJjnORxOI48a0il7nLpXMnb+2EK1zG5yejbOxqUMcnrhqBbsFCM
9yMjWnoOVrJCxjCeujHiNBESYGqE3jUwJfNRoeYg+6VWF+e11cw1BO8u/F7zvYOU
Bkrc12sJkbNQ0e0h9h9xLXEj02/xgxXN7uNt//C5wseigFcH6DrbuYaPJyrYFie5
i28MyE7SHmYUSTiAWMg+wyWJjXfxrUYkGkwUH7Zi6II1vFU47TUgiCztIf0HVgpc
mBVZkuLZhQ6TaEdvAWOfUvwAszh3BDZEdgUrOoTTOZq7Wejpo7taMVhw/DICBzc6
rA66Eh6Tq6ybpW0LztcnObk4e78x6RErA7MWLWiZQQ2x94s4D1+sBn+SvuvN9Wik
uoR8xKxumEm9HGXk9LkBTQ5BXtqvCsLalU2AELAmsc7U29UH0XCuY/0dlC14BDJn
+RZ/e0V/ZE0vLDnq2RIIII9L9GkNrFxakiQojiHdSPjwuRwSuvcVNPyuGWtaeQzp
ebZb+9t3OT9EAqBnCLTqMhLoRlkE0FW79+w96WQB2lyhIEjR2icxq8IH38FLOelP
yXuTL8CNMxfGX6QqiFPGe+UrlUfk5lpfINyQeN6wmCZxWiuF2aOZGxzTaA1b4/Wz
3tYAGFLnlCp6XfIoI19Y246xLwY2PkTA3abo3WB4bzvAitDdVdMF67Rjn5PxzDDt
dioi0dqyG49gIuI3ioY+cZzwJ4NU+D4kgbyaK67dbuX0qUjx24TQ2NIEnSVZdCCg
jQbLP+D7oIxuM7/ONnEfHjo5fQ0/5UJK0Iv9c0H8GuiOjRKQpcrC+Poz7PYQi/eU
jbQsqsN0WvvO0wV/muEXZPx67MhiTM6ByumQTzssan4OzZs5R5/A9c83eRxnF9WD
liapz9tq5DaEs6Nkx8QwloqvF6HpR9pM4GHh19iFJMSqnlDHtIOfx4LVcKq3v8fi
hnbYcslhQvZqbxOrJhSOHv0Os5neXD01m6vpIzQe/tMCKVaEocnZW9Fag0gpaojc
iGt2U0ii0QnvG29pNm2IqBGgasAe9Y2vAzoYKykuMdoGLohqhaMeBJUJHdxKyaOh
rg9uTY6jATOb3XK5SZdvrO0yc8rQ2H4X6waf+HrIffOdXOjI2bDMZPIIICCYPj/C
FwAk485RIcDDPk6Ajtfwrce7rOnpB5/6aIGqMLwWABoA9kmQvhri21KnWDXnHrd9
QofJqB588m+mMtE8kyLSXycCHGOi60VXXzCHCDgGSJ8EWJYC81lhqPFRbqv05Vfa
jC6nVqvvvlktmwayc2oGhjrfUeaGnToYyO2wvpN00ZdppMDziTaH14IWSzDHlhT+
UTzCrVj0oZipsFXVPhykW7qtVPhM2QQOVTngl7ZVNvYlSKb3V6wRQ/o2ebrNQP8J
3Wmc0/qHmO6tDQ8jNobPnJlYrA82sFBXQLqs52dX3YK/FOzVTmk4ij9U/3EwJw57
C3PEdshC9iobEnzy2wF8S+av0EqqoxAetHPKKRrzEtTfvQ5FbkqoqjAr5g0ccq/E
fpj1v5cOKeiOUSpNU8Fdewoqq5gQDYPl3IfNMOe0EF1tOnwAXEgZvwQs4uqTO1va
30CVRO10S5L2lNoqE1LXPjVPhS9kIyGuBHbb2v66veFmvPpl61AFZ+qcx5dGH0l5
h9hj8NbB0XQv6FSLw1iBGxJpDixz6Rbr4EmpLOfq0l6fsbvcRWJr3Vf3UCRHvevF
N8lMi7mU4Et9BTkTJZecMUALjhNh6cuNUwo+q688LNooYLzclkA4F+qTU/tEa7U5
tu2eGHxQG9TtSL9ksUvntcFykSy6juk2PguebCLlXUzWTJ/w5F/45uZJQtTvCx+f
1xHJUjXQkmhrMLRF8qXFyQYHCzdCytvplKw50jI0gZNDJvyBkwPIlBQPdDy1TQRv
yR7cO/5ScOvoqgKZWFEI4pJ0hn/It9thXq6aLnfqeEAkqeCqoLE4EBHUKV4mR8kb
0xwun0855Ker39IuGpoZxzJ/63IkcahNjIw9WbvaIhsQocvNUJeJHEAhAIi15GBt
wsR+76XtVGYCwSB7Ce9ebfZ4tghTAjo4REy+BYvXYCyyHYcFb43/xRMlMQl8JzVQ
3K7HoYB/R1uRWmE5LbzoLTAQHcEVOym6woC45oHXp9yHCMZSs8pB4gyEG55AfHyt
PIuOF3M/1NABFbCwvPzodMZktM7UTcMg7t5uJM+ZnoRGI51rr9lwhiX+d6eJq/f0
1f3V37xmb5h5Ybv/5TGEfPi1gFkjc0wq29zyKNg85NbIEFibvrbwogkENZRPlQfU
AlSi2YyqCSzFHlXFKv2miesa4UyEsy5Me/hEn+uVrT6OWrBwiWM6SuS69zWLLwm1
Mer1SyOMOe0Fj6qZU5/BMLt/Pl0aFJ/fjDb3jzDvMgOvdl+1C/PQPfVNYfrInuSh
XHftaK3K+wVauixLAYq6A8lAVypYxhYu4xhVMLoXsrOoD+YKZdijpfzvRsg2B9ia
qbaJhYtSIHEZTr8oL9FE7cpwGHNzXzlYySZsCZtTi88gpxrb3X5JZe9ySHzyCZgC
x1EKdWimkDUc2GCvWUJhBSONkuIjthREH1mIZVmc+zSc/VG9I+B8GHMIipokdgb9
WFsbXgsmST9i/O//FEaxexMXahkHR740FjmzGNF0M7bkf9X6Bn22iGazwEYFDkkd
jxc6HrhH1lmh9y803TAjCNrICZw2T3ld26ziiA9rAgOLzeR1OQqXPhqCH6i+atDQ
MSV1+xqu17/jrumxpKpEsSFcmkgcR9bflVlYZJqwKYIQaV+KheNpff5+uvzB/WS8
OoS0p0Dtjgdry98pxXW+W30+b8Aj2lp4x3JX2iXz6/W5gALlNfpohnBaXehSD8z6
2vJGIK5YTvGTNfd6SpeN+JXjcPQ3notA+CizXsKnFiag5m4aNC0M2JFPHI6JzNe8
kGKLuxHdd9g4dv1sCBrasnn8BUjd8ThaksvfNZ0rczjqhhOmJ4H9OtXpE9jXcR1y
hQv6E4ON1mUHSFDjTgja8kL+VcRHnLqXLGudCbFDXxZER+L1H5GqxjhdBfEvlCxG
qUwvMuQAjpo0FCrjvdh0Sf+iyGBjpzoNOWKHMs18Qmr+1oO8jboYx9wfg8KxD2EZ
1K6nc+9HF2hDfG4KI8w0yKGf87eZTcRmAY9NNO8AnPXe+BHvQS+J5/wMBsr3/mbL
7O6nh0hcc1RzfPYcJBLa0Re1g8fyMwvonfp238h2tG2p9H7oSNdZJOD6uv5DOLgl
DDxAkLhLwVz8aClr4tCuSybwsXN127QGzq/tcgC4Yo+JEZS7l6NIIhqNoKp3HgNs
3mXlqpGQFfSvaA+JJNLFlLQQJjAJAh5yA9SjyPWC62GcJO6enOlAcQxSPve1WYQ5
EqXLLaRBM0CMD05RnufKlha9PAHGDNs4kOk18WrGz9Bq7dcQ2/oZabc7j57ncBcK
4PiPwFtZ/tyCErmYsjvAqhY3fn2QI93Ohf/HjAPlahBcBepSUM+yGO9LC9VEf8Ul
CpH/kO1h650V+qlBEnLppP+p9QzHhrS25OMBM3hY0FAxcmiouEw6zKb9Uyb7eosh
jOdQxNzuTKKWpzNWHiegs3uhh3FG8BFTEaeuBzGlommFOpk+YYzncsS7GVTBCjhH
Cq4rHTVOf9K7hYOaI9kZz3do2qBc/XERYi6LMYd9Ro4ln39PCX0Rt9UuMzb0h66m
IykZYqZ/gflEAnGACoZc2ZljGCfrKQLjQDmNOemro97KlGh0P9oHSZA+qwiL7Ouz
gmffnZyZpHQwWOhrkm24kYBa5gj5VxuWXjkMwCxC5kBkYJux8RfU/63hP5L1ETQ9
KmOduh5YsuyV5AlpkOdHDwczqoXWmJT3supSJARfOEsQ4zv6MsfE4irA0jmQTiuh
K38ucYFkuNDg9pCQ0THTjGHX98fX4S0CwTN6sSEm/nwDEjFGbTLP9V0c1aZ8kjQ5
oh0wBMUWJztH4wYqpKGXC/u26n9RG3Cgh79JeKrX6Svlq/B4lE8REhxOoKYVKy2s
4Q9oxaSkq2FfAt5r06ypDB2RsHI7MzC2QD6o5T+ZghHwLG3BYSgw6KQ3HIF8jqKR
TX2y0Atdo7vhDbiUWyLeErrPlU0rHpgUeL87NejlBk0MXvMeCGb/u2pTUNzYrRcn
NqNyxT+2YYVwNRTML0Q/poT1qg901jqKZ/tAPDHvREiMQMgSCjh9ciDE/esl16hg
f3sPtp8/ZpNdwofp5kPmCwFgKh7+gR2iL9ztu6SPMdo1pB4EyThe8hVpJVWZ/YbC
4E2wjmitzqgTh0KLL6EVIXTeega8l1qJz+68upATo1LS+/SPHa+SAhtRZAMeYstX
YFLUISuwOoqRF6dpVtPJxkGkH0CmfCCq0mGoVOkJlv+aD4QrbrMxbf1w2FJVAu+h
m6UIrR4hnYX/u9GvZs2+8jcrk7nWa2HAjTAPYsQFQ/PmkDaMrCTi7bgTDI7rmnH5
AwEgqCQRWCIAZ0WHJRLAik47ck70ZeaWFvYXPrrHMbApWGbV8iYPNvsaJoITOl7p
1WkX2JKOaVMMAXt7j6lqG4fmQD7ufHIU88u2OhEPbaKQeZzgbQieyfQTAVv6Vl8Z
nlJ6AJNuvwl945Zye0s+K4XPxWNszQvQ7PlKGx12hK2+NWVYAkFqGFLkSSdhATPa
S4+MD7QCMJ285FGm6vtfe1hRqhlVeZmTptOfRf1E4zw4sr4v2l+r8seAiJPNeNtr
I3izkMj8DbYa2a6DcFKpJAYsFAdHVmnWmHtNLGUJIf4I8KfFeEDH3QCBqa/aPaQL
kq81Tnsrz6W61gLf+SBIzArxPQ47IPoSxWDaP5iXYRQgSJz8WuiskHiqJCketxX+
HWyIU3sbQSGWnNhV0LttoOFPctkATOELsU0NJ/s+xUwHLzs1zH25NjNUzTyz+Dk0
53GksjID7sWvBBa3WACIFuL1MWmj4s0tpCZa0pM6QtizuhsyKnkVLTxSji4u/Ji2
xDkwn9poVOMfMs9cmlkuhD9jDe0miERUIal2hoFWX/2Da08/1FfWya+wveXp1hvg
ciLK4tgeikHIestfVDDrhme3g5FdVKOOIJ2oOyguR3kSJe5wz3KLnh9ptzArP5ky
yPDra+RHCnH73a4UrSPDIjLIXXcWYGPGPuzfRw9pAl6F3WJfdbwDI+mik4s9s8lR
+ytB41t9M9GPwVJnlSYzgegdEcSN/deIqq2kyewU3/MUEPxnGcZ6lHkW6wWUcPRl
mq5SNrYGMGdCfMd8TlUkdScsFq9kJLZu36CzRSRzk/hf+vzaE0jeEUw8CEFq18MI
R1MwIDqcmxJOk+Env3PPPJr+wUYP1LJl2HrabgMO+3Hv7LxbFjFqN/28bqeeVlRt
U79rxU2fjrV6NGlioU09alLCmH2KQGJUNBCromY+KCPNT8bG5PZ+zXTb9yol7Jru
XjP0JPAlSVKDkM+F5wImg0oXkaeENy36W0u4HS3/xAeLv5/Fqy4rs9JfMB1pKAYq
VcyiADgi/G8GJoO+kyZrr8iKzUegrjLtRms38DQ2zj8QcE+tJDKzlyuwiweMNGtu
mfUWtt/KkF8a9IfuNcdhrkIydc3zMjiwNHkZepr3SYEsDbiJf8puQTA62WluTgMz
F2k/iWAUUGUuo/31mJTJtWPO4Ar8pnHxE8R/5oHL9Ffcu3j/A8rPnJwOHTV5dLUr
JZcN264UB52R31GVjaBu92wlBz7khMOVytAw3tEy3F6/Zy8hJxjGmu8QW/xkiUQ6
ZrGQcNP7qfxYU2zx0O4vlcJKjQpmcnOWwI1Sfja9IthqQT4W+Y1QfbXhoee22+nK
Zfl01w9Jbu1YoLr22oBKDexWHdhuad+7miafwm8K3qZmU7H5ETwWDvtRSqKA/mYN
4JMaUkntsjo/v5pIEDiFkGIHVAWTXOtqOQb9q/LgSuYnC9vydKNEg1j9IBEEkY56
o7HzYgQuiZkGEazMwgv7XwkFxSF1Whh/GqWJdTaQ1Gg4AElnHsKxQxVuZnOesqrs
pxdeD1LFwT83JnK4uwj5nKMGAU36Ml/kXUjfXDZQ9iPtbSyGAP890x4+ELbyI/M2
JsCSIgt7sMHwFX4yZYOhiSEHRIzw+EvZKZTto23wa4tDy8ACG3scrXwm1B9RRiFj
6sIpv6WNvugNhEGopsnEJa7BT8Ykz7gCqpGhthIimnJopanxAWt8vM3SVO0698qq
LH/01t2V2C34MLA/0oGBQjWfHeSVwY/5RNcJPs6QocdCs9i8pjV5BTCWFVeAEsQq
tX+QZVbC93e4mxefS8oTdqAN8cU8hgB2JdTAhNNWY+fySjItfs5sdO9aznhFvdCV
gIQisfi1sVYe9K3IDPzLzNQ15RGS0qPlo0elSqJZc6SEMOWXsBY09BVUzV+JyB/x
MRE+LKwIxtYk5TcIyo3v9Wjx+ZYuyAWyHEmzIvY6+Vybl2d8jvlFs07w3Pfd4cb+
P8kL6gYLezM9Ca5Dg9xu2URfyY+UsRXqaaRRug9GZIdjVE9/5gmbtu81x9THbLC3
pnraE1cC7Cvd0OHiCM3yngsZv6Hxyh75FGuv1aLjclMhTlGc1psNOsuYlYAAG+i/
o6qibrCrcgJSeHQeQzQzoNfFNxU1wHZeWUXr1v+NYfql7cRqfdCL9WaI5cn3L5EI
oZNoV5iDiaPpwxe7HTM81aqqOUMPpvQ0mqTMlTQrKxhNGhc0SuzB2+HlpZlyf8Ee
4Gkcto+Ipr+TD3wMRdJSbKNQKMib0K7PV/qF8TOVwz6MJVRTYcisEkmgwtO+SwHp
WOREOdb2dnHdd4puQUsXTEfXBAv5rX45Ip1CW6iBhwIAQvmYH7jZOCfi6PZja+YD
EmA2Wo9l66on1XJWb3VzXLNo6cQ2ipoRF0gpOwdr8/7brvEc96RNm1ys9rG0h3XR
woU4ECVs+Jr267c//EelkGISgNBj/WpW7AnvorJqj87wy5CTT+rXro6FROG9zSJi
80yXDSfMTTjf7mw2APvQD5rjrMq3lFDlRSd9t+vXzWcqhqAFA80uUMBD73X8yGMQ
VjNT87V6mOaqFnbWUzm+afzs/GCSd/Pfb5E94EZCbv1XZeUS+alYJwubeeQzt/f4
EblYJRzcxrkzTIumFVVKWadWiMifbFbQndTKHzepTBfYXmo7Z3UtQmYH5kh2eKiv
tQtZzh+Abhe4yf4tMnh6CIVYw8h712yyVgTLLHtkBMbf6qLHLj67YyXUIbfxqFi8
DbbKFfnqPsNjH2rHTagTjYEojWa8P3KA0MpovHc+J65RgkX3yjy9bs4WpN+EYlkI
ba7foxoAtDFXaPeVW/la9YuZXyHe3VEULjRu4/L4VRaT8QWD4DFo45CVeg5gQ/rG
Weq3RpPey3CxuGtBPVcDSa2rSO85jdVTKVjn8pJMPH/ygxMvw3wevjL9TM98T/z2
LGvFof0NXW6E0m1YG+8UuV3oztxSflo2NXsi+YNHB3p1I2r92n3ier897UbfXR/j
AgS9AE43k6C3OKiMDlIw4CrUn2YYUmJ3wwFdfuaxPU64yuoIzjPheApr+3bZg0S1
AR+Zjlo918KYhueCAeNBms22t7GnNrj0OkOwzUWIoUwlY7TEpSGVXiN/UeOJhWHH
FUXDXNw4m2s1qGkEMhGuCvBwZNCUDRBb1XBrLCuD1Wy7olscD/yw1Kw1T8y6QGn0
Yyr7E/kpfIG7BVUm0d9aZwFPDVKdP7AVQ8PZzx83eBkO9yePxazg2FxoXo8Mx/fx
OM0mzhu1Le7+CQXpW3bp6EsA1hkxQ3/nimJ9CYNq8xR3+4P5SAxUXr35ygU7nM/r
CobjTr6fEkxXGs26ldOcV1bEeGdBgtAVtHAmOgXyDsMsRPBebI8IVDyf7jXzWsJt
v/6UnQC17zcNVrv1QWmWNpo7ZeXkneHWW/53bSNh83QjsJYn0AWvdohqsAypchrL
GrIc+1IZ2A4NhVv8qBK5KJ2KXBGYo3yO1fR8k/pu5Ie7hLZ1YluXUl/mSAQKEAw8
leE6MqvX41OX89TPK7i1+deSWvd+Uhs06S8KxOa4pkdkoB4SipKGhIg84smq2/Uz
yBHKaHZDnxGMFFzs3vXRmfaBhZnxAT5u/c/xbCgq9nI4vPt4tYevSMATk7Ue2p+u
0EwHhi6nbeEKsPGXjLd62fhkSl81evq7ffqwoUAfy+jnETrEbm8eMs0UgksPlGKE
pwsgEvrBdRUkZvPgj823Pz9cqjgRzerSD7ByCxntxLee+6X3nQSV0lHKSNEGLqy2
j/jDK6yYzG6tze9f7nPkPvVF/efpFkKkXkj1vKybO7kImYg1ORu1PKX/EGaNT3B2
BihBcrFoil7N0xwj4MvEayzn6JjSvikK7+k+f/yHGzpbH4NOawxq9UsRWaRgrNS+
6RGFAnicUeKjWAO/VgirjeXVPBptxOawMn//QnJUk8fP/VH7MhHIZbHAe36FaXrd
CSFZTpXIJ6oZgKmvE8M9fJCWOxe3gLiR18JRdJ978OMQXJoRrrmSISGqyICxZQnb
ej9/BSovxj54s2q9lp7Z14lsCjVrSoPqatjSbDoCP3qS1U5ypeeZH0WcM+I6LJ02
5ZfOn+Fv1jNvZ4N1VbWQLlA6wWBkuO+4hZB1tZ1gJaeJPWW7jD7yxQ975PVwRKlk
iuveDKXjSlo6OidzLjpFdfC0cp7Zxpfzizp/9rJLoEkTD7rqpmobjngpywHGYCu7
ThUuyMoGInQPNj1C/2RRY6YzdNyA07O2lLaWJ+VaIU9wpbLzKFiXbjqYwPUESQeG
UI9LlZgDc6nBk87tCVTWgqKJChMHE0WsPcLTFF+sSoxge9XUw1acJ3n8GVCYu1aY
DvR1fCmMJqpAY6adqabcCiUguGoGz2c5BmArgkYk0Yk/82z/82aUgZxdEqTYMuJ4
9by1IlN6HTcM/jRnEANdeXIhseqfIcY4IxWmy8Ey5ix5Nt066Sqsv+c8MHB9NT2i
Ih+ls32ake5pkWapdJMaVg8XG9pf6Qpo3CeFbB6n7OJoEA0Mcim2XtDRO/707Ffo
x7pvo3JRfjCwYJHBxE6QO38siR7lsKOCx9ct32fUgtZjIpdLP6qKdoVtxiQRs9h8
mo/Ykm+dxA9LIATlbanWPUbvKln6e4yNYwt5r38Ic7QMemiDMl3NaQNwUhJOunXx
2AiLlKntCBRCSNxTbg4AwrygShlCTt4SpNpNmN8AwnwRxLEz3g1hNhsSPbeh7nQn
mih/y0rX0aUyrkTbxrOh5ClRRGhvKSWOus9Y3CBNw/sy/+sMOia9RCZwXWNITUsd
LhGZJYFcT1eQlzfQVZ9sPrIvJNZtKkyD4oFqSv7iLoYI1CM2jhQXYEJMtfCqoKEb
3lax2xZtwvpN20XYgBlTMctqSh0GvM9HyAPke2RY+svYm+c2ohowJ2eHJL5Lns3R
jp47OGQbwIumNAYWA9Twmq1UTxSUeC/4oGZMZoKjEPteDlRzU7xjF/Xwr7jGlhwz
MV6C3aisNyjWjPQu4QJ4rB+RtCRsA4CrqjR+aydpVKJdIu3e+SKo49s03rIsPTTF
VpYrTM2Sop2o3txqUXew6jd4dGGDeUIT1kt7HnhdKTqQwFuVQjlKSadxcf6+TTh/
M31m6tXYeqi38qraIZS7Ub1IoQ/k5VrUEDJa2pD7aW1e1b5sVFHWgrEGvAOkIVWJ
IMTHyQpoqYQwrA81lihSYbT4fxtVLga8YoCwENQjEcqv/4pQzK3oyIbb6JdgqzFB
/QVy0Mcq4nFEOLJh7hqpFX8qwvAbOIgWTiDFwaswTthZTQ+xc6mulh0xvkNBBkPY
W/mRzqsghhPQEBzsk8/BROggPz1OafnJGmwgoFVpdav0uonb+Opqd2+bIXwDnbJG
BmQUhL0DJUxC2XZ2G0EzjhQsRl/xgLTDYdZp9dQT3JdfyodUZUDShMmrKnp4CpPt
R2q0H4UQbD/A5fzB4DF9gpE9IElPeDPaeMKkuSrDUEtm8UdNQjpmhFWg32xo++V3
R2iGvmnEWbeyzAXRqc+aLwY0ChDn/FlQGz+FxlwQ066BuUHqtKPOzHtoVXXP8NNP
OuXcIpgC1dUSEUSEHC2srMzkmNtNhRC7XnV1aybNh6cX2m91EbP73I2B3nWUwixL
Nr15bREmBUejYsHkuB3caOktUl7R7P6wn+XwKe/NoO7dJniWeFUHUTQpoPRDd65z
lcfSE5i19tlPkyMqgprVQp9WiWihq53K14x2RqqNzZ/ln/IbxDt+S/trgv1SdmWl
mqKq7ChdK4YaboHsOi3tWrI4IHHTSiaQK08pzu8q0S9YkLVLix360lbdRvyr6vNs
tmtL/WisNYvqnSE2/GnN364EapWWlJjMGi2eL6+Fmbi7RUkALl+h7/1zAQ0/+qE4
pkdRn8jJfhKEG0vBGjZR5qEaMkh8Z3te42hbD9JiMqjS5scgN3EGUAYQ5SOXOt+3
l50pXG30tlpPSlUN8pSA7VnvtT4pHYvxFQ9G9KAZGcLhvoQW1+84B/yV+Ik3BHob
qUSGzvmVXwmNkSSOQ5Lg0wCi41RPP1dSlbpBWnvkNEYFRlut9bGXwE5C3BO6uzm5
gqGbLrT27cI128budqcIFzZnjcPlMkzt0JGC3nV/Mtr25lO2hWWVqZHpmibIiUSh
hCfCSEvS03qfnERHcx0DvK6FgpSzI7PeY0e8dQhZx7hI1tD2CEpxyVNDuR4eGpuC
3JMeAg3LxLmdGAAOBXmOXnZ8A+IzElivVmiyF/WEdTJQgLpp4Ir9+HVRIsAZcPR7
7uZwGgNCQoYgfLbkTh8mo3A5izjns6ZROdXEfqQP/6vxYtEApOJUjFlX0Hjvrefo
XVxbNael+1YQ0DE5bCRJSGqaSYe6HujlpIYBW3QocPdUIO81kletYjL6kT/EmQRU
/JfgxyyNxuziAscKSDs545ncfheYHV9tYfJUgSN0206jIbp8OnydRj1bcpKzrc/l
u1rUGqxwSEDPk00pZiVofhzMoB7Q2Zh+TdyvQpVX7NeHzmYPNte+KHajotVPwBtN
uOTdtj3qsVNJ6Q1T9FToffn1DtbpX7YFWMmljbvPvAkgylonRB9iHpktZkx0q7qt
58HV9POpLAiOv2xJCUXw1kqfp6ysWA7aUlALU+5i5SODnn2XeztRap8EcgyIzrYt
XwdSzHbOd67mDXgWdA+Qt62FxoRze+iNBb5Ide4GlhZIbVJJiUBN5I+n12HJ16wi
mjrypBiuZGlAPLUh15KdsRq83Dvr9p70x+2T8X5wtSZoA5xX05lFbbdC33/hpQJI
B3if+IeQSSyI6wIxkeYJrAO6Ebcfw1bFGwfop2S5WRLXuJuKcyD28Y6o7tIZk2c/
x1lq2hwPVXnl8Mv6YUFHFeH0JD4bVByCdAfi4oX6app5TGzXAJVmOkjM4/g7Tw8Q
8RlwX/Fjgopu5uU7ZJBGb0+sWPUmxVcBh+sPiAEJmLc4yK4SnXesFnbrPT8NrSNL
BuG5sVD5a1PlCvNgnyt/JqoZvr9NGx9CwM0VvUYe3gwMZXj8BceevlP298LZHLAC
Rg6iXQ+nNvt8M07SnmGfemQg2t6xTrJH+qkGnm38nWVsiwQEWGx3TyiuxsafXJZ+
HmVO5kntNwvAoyBLYY+xjHZqknUfqGyy1LQhZsqjvU2Jbl/NXM8+nQBvai1Ox/Mc
Rx3HCnmlPuHlQWKGmS+3wtPNJpS+XdzW1qEr36CwFaH+cUuC5RUoeRe3PE6qQfog
aH3aTDfwCQyaITLn1+bY55kO8VljUOKLZMMbjgwIpG+Yen3u1bgPmb92i8FAeRMU
1w6NuqpDql7B9JpUCRe62lPtfRBNpqgiuRArz+y+NIkuhFMH8Gx/6fAsO2z5tA1g
4hgLNHbsSUU9TYpFKIQz2bq8mxz1k1lhvf6SJimPFrNse7dgVWZB94q7frcBCqxZ
nURdH8bR/qzmZWsD71n03zwCzkZaKIu5pHENbXqBO4AvSBrX3hWHyvVUbnhATntP
GwfIz58hkF63ud3bTF6y9RNPgZ+ztO7N6moW/Ktp7npxMLzxwe+0ZfEsnReCqqgX
HcfF16/w21beLO3r6aG861lfqWP1uS7hm/611fAL0Rb39jlM1Ge6kFPsjJzpTeMS
QiCFEqdM8ZPF8ynbLnwXA9uIEnW+SVX5zroCR8BQ/57i2KRrzuuAn511aJPq7ugP
FSz/iwpoHM9JaXdCiK/ybFGm94Uq/NtROvmWmy4Z7zLCSIDsv/0gzC45ef/l4QUi
rhOg94DkSN9KmUWJ8aCZwL/0kRiSeetyFtof4r/VwLIdRzS3K5X8ZiOsuW14v6BF
ukKUHhnlw45Yn2oqmmEe6hwprOgqE3dbpZyK4hXVbl3zXI60r31Xrcpy0xCfhqQ5
GBH6l+uTSZZpN1C2yst2s9uS3ujqKIC0r/g8hCl9QplOHcAT6HIfLDPSrJMNfx7B
E77sq14HyzLyGjvkXPh14FXO2QcR1dxb24BUcXFA0sfHmt42hq9F20SXL8m59EDD
wZs7NJxaSefGAWIAH4knAJS+pmpNslVUdf3LG4hDhUWSSo4gfVVHdzOm32mSW3FY
VWH+RYTSwOpOjPOouF8anv6T/CwUj1N9Qxw7eXyZXJhUp6tWdVVbyv5n6Ex/R5if
/czoQeydlhCD4UnrVnrb0yAH5lNUp+HJziimm3EJSfvjDmfu9BAfVAUrgjyrJ2zv
AwvoWlYQJeMHE4Z4vsHLsHQyjwwYNHm2iPuGIDUG+qrYk9Hrh4NeG7vB7y2RFURe
7ieUAoO7Y5iJTm1TZt/cgmhdQq6VvyL5oV6bxX8NoOzk5HIxioQVLmzTiDmr2E6k
f0DFWd3gr2yis4WVGEKZUJdHMYOYbxnCzslA7wTxSzcJBJ8J9cb/603cttmzAiU9
6/cK80ydelKQzasQ2gUbqpCa0xxmbU3S9rab+b0VNjip06yOk7ZFnisrDZkVeH7o
5EbvZRpfR/ejOZL0b5y87uhs4CYhh1uVR5rK1dtgEBjASlDS/ym4BZGcocN3Dh9E
j1wjYvm0y19e6JpQFIqe/x9OSFjG/jJNnIIFuvQshUNt5+RBmgIUP4ene9ukhLd7
gXpmAOtcEqQLybPBNWi/3146sr06AivpdD1O41W4DKHTgCBoTQPNT3rF0BL01QPO
VvD7o+I8X4Gf57AzXXvu69HtskrePYU4YM5VMrftP/Pyg8PUEyGhJWDuZHwHfoIA
+fQ5QDDbCaZH6lNQZRHIA41110n5NJ//W8fM8EDe2rfJSTT7apmsjMfJXPss2kVb
F4lTqw5pnwq9QjVS/g2zGq8gE5ShS+C7WPVpPUUTVbnqWWpUjdHB8E52PIdI3UFx
FvfG9FT7qXkJaBo9AFSWq213OFPTDlAVLoqZOM5cA+U8wXo1fi04X73xDOCeqxSw
sRxNTTE4gJalQPV+So6Xjw1o3GmUyAl815BMBoC8nnfPge/usQ+NK4mhIaDYIUx7
UIX+BTXH+UzxFyYZuuX5JjSQosRB29DiVOzKVE612NPEZPHq9NpPlvMmimyEAH03
fw6r4zb70VkpaK+71kSuRUsXjLRVLPj4xK+8vxXswhwBfEdEaIToypM3RoUSO2ZK
9hTTqX9643wz+/VsxD2aNp7MVrglMZB7a+Jvn0V1oWevjaST62E/iGNUoh1mYz7v
XRGAp/u5UChJqlWOQ2DpfFTWTCKqpYI/lLJuzNIaUNE2k+25IP9HQp/mDgu9zLis
GEzx/n8Hqp2lm9RP8h7v8NYb5qxdS9e5e/pTnhcCrcKZCqS4g+v6C+lZt0rGfYUq
x5Hbd8d5AZHpIFC3cugKCPu3MuCfc7R08eBNjgkkU5wLpgAVg6WBDXpHh+mvsmdI
EU9WvNT/Sfk9jD6QOM6oU4nSfI9au7aP5Q0axhe8DMg92RkTrR01bX0tAzH6+LBB
YiWhVfgBWHk3wgw7rEiOf5IrM3uMhuQG8pkYKB6R5FurumlubEuNrcZWqvdDGQra
b+/a6iutin7PPvYLIxfkjGHSmJsnzbhdVTYS//2Y8CugnAYw2pSyGOTdj3B/nlDd
DQL2hxDDZOG4SctIm7t247LY0UUOQEKyyfieBOCZf1YV0/VnpnGJUrv8kFkhDIJm
u1PHgAsBYhpacMuFkYRgs5TsDcjBGskvW/0wD5u5eLC0bi34IbFwCsbhOYD/cDWo
MtVf7J6QIEpyDVUf8XhepRvgXa4L978CuLg35hbJzPfh9AKdFXxFKk6Pu7rPl+j4
jQ64cOjAOWM/Jw3ImCqAwAGJNXzkxEzAai9AS9BESfG48EmpQnYToB/csep3U5Z3
j0dzlbvQ7843m23WVuaM4OASxzZ1GGW9eiBR2GPTuGloDuug1D8zW6DdsS4qiWHb
ijYDhv+A+gH5+fbgsllr6JmpNX+uK1X6nLVOfEeaHtLSiol51Vphysj49XgJbwtM
WacWQCYzAujIJax3m/28Hue2LEgYkUqAvNQy7/RUrjV4KxIVaBZuDVBNyS+oJ4yu
zfX10Br5KWoV6MticHK7baw41W/0bZEo0jxDrDuR68wJPBJP1F+Lg/w2+hO/+6fx
DGNSVLdd3nX0axjlB3KsdMDEQsaU/r4OrW/aNcM7Uy9ukgEu0R3zE/LWtWMOonnJ
GS+fLe+lyDDaOzvX36FI9UKG2Rwxr+GyjGkD8/qJc4k8UKxUj3vZm6XWRb6rhDO4
jeGxyB7yhEoJZ6TP+zioXBsZESQE/HEUn2WL0SobJ2n/4nZwOJISFRdIj6HStnL1
OTaze6P+/HoRh2jCAOE71iWVssSm25HJ0BeIPMd22283labgKROf/WFrCY4OjPM6
XzgFB07XwL0EJsp/nKR4fJOf5UyalSDIrIOEabkCZtijk0x+EHg/uYZQRX1gIjAa
rvqW593EVOfqta0djDlQMeIiY/0YJKvCKAssEje7MX4zUOltith30BF4gSc7+vrF
PmHpP4iSOv+F2766f8ZikrUVGBPZVsfbxjL1Usco3YB5WWwUe4qesgTm8KZ1JsLY
q68hspaOaYuEaN0ty2QGuMU+DOkjk591ibPtLA28r5YzANNehfn1pBkpghUEJ9bo
r/bXXCxf9oby2jKvOcVrYCH1u4VlcRCcjPW5IcMmtun625EO1Sj3T+sc362bYgMI
pXtck/qmfaNCq8dUmmo4duNRYP+pbWh7Q6rOV4/kNrGnImR7hYV91NTOBa64gFtM
U7wKCscVD97W6M4xLIJpO3qkdDwJf3I1Kez0Hb3qUMGC0v+3w2LETM40xnl+OOeL
dyzgmEfQaMeuKDMlP6PuZU6vOb3hz9jqwi14Fg9qZUtH0SI/+jsuTD+o/iN4Zybf
xnjoeZmYEJhc41Comio5Dg2tRnt333RQb1uCZvAIeNaVuJa9Md3jmABjvrFIhqyd
tlkUgJmoI86P7S8UrOsO7qX1QKZRVAXlQndihZeHM4eouVbRBteeqf12F4IkM3qi
zzv9Z0EZZ2yRDjnqie5avHYDD++ZuUgJpONoUFFvG824VlqJo5HNJOaMHnuxq8Zq
KmRO+4/OrpXG5ieLiygUZT1UEb1HkdcBYTwJ7lDETFcJS+AQ9riKFOIPM5dOKBPt
UzwclCAMT5CeU/BEGzfIBOCDRmGGwUO6FgdLuE8T1wZ5b6Mzc8454vwuYbcX/DEW
0w+BccvjMb0FGKkDAFDd16zqLTxcFQrVDGs/gRLphkQ2pTDPCH+KbqMqSgSUF9GA
Ud1L4BOAbj+/dlNWu5Kn7pgX6QPYGYeaNExzajT45jRAsVGbSZPEMpyhgOSVEhpP
ssv9nHyO4DozdIyObPBSRHjToujfuQZk7b9iCTYvTaJXa3FLVx0TJnQZIBhaZm1h
P4R7VGIyYnAWcfgpWX7bKo8cAGoJePCzRKTMFSATh+wV9FNeZAm/varcunsJATre
M0Gs2XB8Kli9gFxnRRvTVz+fKsustXqLAVsk+q9RJKpKwofXwj6BGTVfeMuOQnT4
jkI0hjNtyP2CL1hPMfC0XrzX8tBst/ZJ5qhKWMlP4CIZrDNoIZ2o2r0d+FfMqW2i
9xa8IPFcXsxzQE28VL+PQK7nTwHyyPuIEyskWNAqGQWo9Gidd5j2EgKtTM68kkP3
eWrd3DxXd3BohCdC8ELq2h0G4AS3dGAOWPcLdb8yxUTDpGVvnGQIjXnK0hnlzVyY
lVkDYoBisII4hwvO7cC6UYye/FHIS/BmHEDKY8vB1YbzNUnYJ2fJq/D9bEUI+lbm
i8xMH6ouKLqRjQtrAvwc77dFPEkG1VKCB9BsTdtFR1fe6c83GBHqGtVOQKvBnQrK
F7PWjpBu8QHmAY0euiMAMi14sPmA//pE454tP/OdRfz3r1qXMCMq12OWJBeO6h4g
jcYNtIpIHHSZeQn0AuntggqBgHf8UY5VXDPRCf76rMMc7iaXos8kRNh1Mv3IgBA1
limUbQGmj5TahXZ7tV3LcpmHJpwGfcmQGhDCQ84DzjwIE9GsPrChymP7aqHm4sg/
6fyyerCD1mycbnyhDSguPGy02NNZ2esT0XJQ5pwd8u+wOhJPMud9NuglgRVHAsde
SyqSgyRM+vCEp9ZRJtUdQLrvwtHOWrD+NEKSKczMZftHLG/TtZqKKCmndhBJkLfo
T+6jqpyzpofSgLJSWw26vU6aQyKJIYNJmALG6lF6CZvwtRR59q0KHtLOtq1BZrw2
n5wmRJb0pYzy/X2qXsXVLvV7jI2G2I+gjjX46FT0iA3RWQZxm1XnJz9XVkN33kmL
X+3PEZH/VxVmh+wRvwyUkZg7+frw4ufcxUP6LZckTGhWtTlGiZum7+Nwxnx7iv5b
9rjjvHpUtuS9MW41ZMljvkbl9MC8Jvz4lVlAgBs9oX9VapprpWWKZ5nbEbxgQnE8
RvQaOgW0KgvczxakW9NiFP7P2ABVxt1XCTBKw+8NRRfTTxm1cPazWVG3+KunAk7A
cB2VhEEEz0kxM5mLlxknl0/UZm7yqhitoGuatWEWag84By7Q7+9RXhNtv7v5q7hW
jXIvVWcm5Iyne/WXDDxEBn425R4U5FAYfLbghIY8Wp1MAjcZQ+PudQk+DM8JFxaL
Ue3su/OHSH05Gt7nXdmryHDI05s9xIYqtB0GTjEDFJRaFeK+kCfATDzTJyvzTiDg
PBgIirC5WVTUPNJWk+8OxfafbZ/4YBdpWAHOBcxYuHSl3+HrkfA8k1YsRP+4sreP
6k/jmQaDQrn9yYzfFlRYnx2oZ5JBTvY1wDF14IdGZDDCSkXHNnqkU5EutHK1zEwK
pHtNMFa6ClQxotGHbz1CBi8SnJ6KgZ3k8DWu5frarrsH4zqTOT7psVym0sIMCHk/
055CA9D8x1ziBFG9RoANn4oqR92HUMcjepeS1CcvNjthMIrfVT+F4k7a49nsbPwa
ZC29+v0zdZOuoD6XTf6jPlj4NC3hWMr1wrPUjHGiI1BJyLoc2hecmvB3tJFHwZjO
g3a1OnvWG8xGiBrQxyQfDAqEsYITEIHSBejMwEXR15H49lZ68HDm97D+cqLVsPKk
jb5gPZIPlfgI9oNnGjvJ8zmUTt8P0vpwS9YBs8tJavsN6GoKC+wGVW1oC/G3+Un2
fAObnJe8lkhnS/KAxE0dTFV5hD16yEdkzq1203IzLm3XW55NsVildsaHCdAxJfUx
eEz65nt94RXE+5l/D17V/T6y92/hlD+BS+M45fHJ61+P9soEwd6t2e8gOWWgQUtK
n945MPGLv6Ho0kLUeqxaX9+iZDeh/zFe2rVvqXTs6OQGegFDXSFnx7xt6T52rLWK
jjkQ5rhN3HSTDS/VMVRwDMYTGa0dTitfcypghF7JB6Eo9qxwN+X+DCYr2eaFsJ2s
+7Qw+SLYiFPkxf8+f/iVs3kzLzzfrI3i1j5D9UGOAE6SQKC05lTf7rhdAT7yHGyu
Ih1Z28GX/rBBoEQeFz32I+9OLhLbF29mc21OHm2QO4EpxUx5NHPIQHgeuPuTIIe9
JRr1ZhpWmoPCB2nSKBksKH8B+bp+hQfdI4IMEE7Y/Wzocin//hJoTIgArJ2URUIg
LL33S1UiujIRbzbflfaKZouByj7mGwhqm4CwvuSmmJJWTR5sc2lcyOLDqZJCaxgz
FGpPn4fVg3aoyfgXYvAOql2HT16F3ewlYrXooqTejiNO9TJXedV7usRcLHhz5OmS
TIhrnDmg6sp7SX3XPoJiQYfSszurtFIDdKcDExopy/iq9o3VUvdWdt1rZ4TydkW3
XHc9uJGVxGuQ6rbfEAnbkJuF04d2ksP3GRxFp/QRJGjAfOnwz7gsPsW+yItHofGm
GMDgTE0tnUQVZMrLr0jkijpEXC1JAAldE89Z5NvG/IGjwiEF6Sf7/u8xRbIkEYHk
/ClNXmla7ohY2vS4NrAqDm6IDZXWHBCAjRsbz3tsM0zhMQBHvzzYM1hzE0jtHD7/
R6YjIYeemORxlwPWjkQe5a6nOJ26oxmCAR2lLHvQEMvev+Wx624VrZ3DR8fjqLvg
oF75R1dxWTKRGPgBNWgKuOVoWBf/NUUIOQN2dsEn6DkseA7AWOR79FHKpxz+V4dP
2cy2xOGEkZ3Q2iYwp8CUt9/rGQWCkpWSMpZUH4et1WusMpuqKK9oyXNz4IqlI+Rr
z6qv7O0LmlxFYscz5dqlyhmGn7P0ms/6R0QvIOgmCRcUL0D0vvg05ifmnDNWUQ2C
isEhOzcKrMt2qsQv4TKXF0F5mceKb0YTUkfgIuy9OpW/sHWeFeagFg4Dt8ghaWex
xZKGlk4LtQ5h4GVxrzqVDHLTrmmEh9PEH39n1P8DRyPxVVcqXTC5NiR+IhKYh3l0
zb70I7H++1VWEqOcV2lUzmDZ0u0I/O2gaJBisZUMRZWu7o9cMOm/aZZ1cYt+nT9p
SAbk9KzPVcZ2p4HPNICfr/zO7gfeSfg/cQwL7+rFpVRq0GuSwYyg+zQC7GI2uGwr
3jhrEpGIXwdE1okSn4+QHhP6dNWFo1UqLEPOxlA/cxJiQJIeXX8utIGFvo6fWIb/
2xlc/KR4yWDoeF0vnRtNl3wCVrYaiVJpFTLaMrB5qFYfJSAmYsMJWWXOJDb7/gBM
JOBkwm1fQMW71maVUPQ1B0L6O1Fd0I9+rlUWiT7IWwXx4rrsD9uZ+rq6KF5SOPk3
KHPAz+gESiaKrog/fp0ztukW9YxylM3l4BbIvGs0roHa7Zk7m3ePa1vqNNDY+6b5
qgcABP5gfv7THb4Fk+0l3r4EykdU4dKmPNRmGFeuw+tSBWbXWhPPP/wVU/zdfaL/
fvwRTctLygwX4czKiB5IgsOschgApEK/O06X3b6TgNfxOWzVHO1MIZq84G+fOjw2
tGvXzY7xgy3A4aoGubQWMHKJFYi9bqbFD5zd0qntEQBMt09hQ5xxlIH5/p7KuGut
7yZ+D7mFovhzVlJq5s5esq7X3nvQCEN4533OcNnXdtkcAci4HydCdEMWRgBkcxqT
wt2oBbfKMW+Lc2qiFdVldHtVRLWE9Yxt37iTorUut4wCoykRz4Ucs0jZYSgk2nTs
3OfBPevwwMf6o17kIY+k68n24a1K9FgQrl0s+kR6VAgjmX4fXLVfHW/rbnMWMVKX
c+Temqc+Fn3NcHli7bAt3VGlTb2oy668FmX/VBOw2Xecg2PHptRTNzMoot5vCR3S
Vjm05lFqWS3znn+2DArJig1zXIPdAwydNzFk8cwmFfN6hl+jy8JvR2K8CVPWd2f1
xp54aWqwD+N6lDhskHfY2YvVwxGYTVYG7SXATTTltUqt2KGumqLz17vyTcbpSkcv
ad+9/0L5/CcjP47q4qlsIJ/bijMwXt6Dh+D71zNoEI0YSPCVfhoCYsybFj499YId
cGWSUu6CoeEA07gorfCZxD0S0nTiexujKq41adXxN7wc42ySrM8OM4/tLipWC6pN
jlA2hDSG0Rsl+clD8AX0WAv6r9UbLqVe3TGSycHInkGRhtqvZbuVu9Hkaz0imsIc
BvSvC/yPCYawyqBHyV1f8DmgfVESEmBOgrLeStaewMSAgxByJkswV/WJkYpeXQWZ
44XsYql8RGZq7qj6G3+kBtaa04uomQSOhaEPNTVRr38zvxBFlmUZ0oQrUg02n0Wu
61bh4R6aKOztaqDPMNmqjajaohnml9djLq7upZ2U/beelnJixrRKqFcX2fAR8NcD
U9PXSuS4avoN8YiKsi8efCra/AvsyBNu272EKVgTwMcoxMK6kx0BLc7r1D5ScQce
yhTUFlFV3qDWouVTmSAqKErqK9rW2WYeBaygPM5w6205Qtkz1ddpNYaYZ3O2SxTE
bqIdwIoztKiZksfdUQdrzYRPi7vvtfnW0D1XJAP6mkszUDZjMQQ7YdFfUF+I3RXt
6qceHJ80eWjpm7X/b9ahUn0aRSXBvTr1LXnmZVnt+3AlT0u4g4t3Vzcpzk8kBdwq
Rr1Yq9PBXElzb9BoNqeD4WobM1ZvAYXH656/6wg5SvfbH167TlLx9qu19Yu40XOh
UxyJjDo0WbwyFB4KM7HvOatdXokMf0MV/WeuypLhyai8fUOkqVp+h6KrN0djsN+r
w4IshGYMSSLyX3pH7hetyEW2EpP36LEe7WW282ZUZj4iAOhS35F8knzuzkJDgg26
RfGtejHOrAsIsEDmLC3HaHFlA88YHZPipvSHWPrji5Ao6WIdsqca4H22zFT0TFK+
eduw9HZjPZm059k5RfnJI9tPvJHYyEUvs+2pzeVthXkU6VQZwu1QC1j6RpXeFr0k
hZ1AqDoRSQRdHcKh/4G51mNtz5mNt5Rda6tN7qlFkxLb0Pmjw2U3qNpR1ZAHJmXD
ybD57kfrwqmuj+pw/CKJNgOh23i/3Uy3CkNIx2hgz96IMRf8lTQUtV34qauFqjiM
skD22Vmzv7NTJlHYUAzPx1Z4AldyVjZ8ZVJ0SDQs5UKnnNFi8cUQzep9VyoqTF89
YmdfgZze6Gd01G2OxIrGA4fsRpgvAdDKfZCLg2u92SMb/HgPhY2k0yP81FLJtgIR
IBE+WD4ea3pfp2mu9ZMTjv3Agk5EV12oXA12BX0kZEQ+HhIXq5cGay12+Fr5q7jG
WM/oaV1haQCBq7isg3YaviTyimdFHX7WyhgVxU4NABrAnNl/e1vanhY7w3Fafl3O
qejC4KdywlKhsI+SDctDDqOiG+85qJepRy2JCrRa6F9j3jzFQhdT8xZw0geE5O71
pWTzlvJ4L8PTDD3XkrPZcz4ICkC7rkBrJTJfi03K5jGTKpVd+9NtAsyIcFoNCSQ/
UoC035tHk0N7cTqwrxr5u0NzhifqnHGMWiTJjOeFL5ANYNOFWn9i2+MGcNcMJHOL
BRfweNCI8REvOI5cb6tPRv0MMR5i/Ma5nJWjfUIbDQhTf3kpKST+A6SA4eINvN6G
a9G2fLyUpQp6QVksfd2f7YiGMD/byATyzBh8c3DzjL4u3CnmvTODypVzVVwAxMac
P8ya0J/h6v1i6LpA2mihJ662L1VNR0sd328g/pF90KacPmXdn2Cocauyjsz39o7g
4/i54lWyToMfrfVHyZZnwTXS6RhQymNKXsZiTmC0WI5b7dfczXL/Sa1jg7yAwy1c
wYklxW++Aqmpi8kW+XAcobWIi3R7AWPcuoZ8isAr+Nwat+/El6ujNFgHya8gqJYX
0mzv5vK8WnI3fsJKRi+qEKJ/2A13AtvLEOxx4wVwSVQ1fv2B+q2mHVUUZBpzOZUl
KWUzrK3QSJuQ0+wPDbjyYkbDBnP9mxaQgB7rV+NKrvSXFp/ZekhcImxZgv3eqStu
mlxzR8oa10GzvS8ugJy7HWmgKErnEYk018sXgWh6Dd6s5BMT+hPqX0SBjJo23qQn
kZ35gcStr2lpx6POAxT0qbm2xoaKGqoHvccaccO7VRimo206GNdJQQn51rAsuz/a
0DKGzoPi2nUtKijXXR9MQlzYYzTZJd7G3f7OKmu4SBXQljUZR/7pMqZ5EmYzcFol
q7ncciaZ9po/hhSQ1iVW06qVFKg0xiB619nLneger4IZL+k9o3HjFhvCB9vssw80
ernkyhroJKiz7sPlD6ldD3KKnPRperbN92gkf0KQrUa1LxqDHvoHYgNSjMMxL63o
s/Xs7Iy3r8Vwgbx61sv6d/kpVhejsLXaYFT5NNXDZP6cWMOAcFiXBKtvSvMzDz6g
TR5HLHgsZrJXfTNBUarD1f4ircIXuiP55IVKFGNOgJ5WCZEsj9bktNkx2rn1W9Je
lYsCZF80k8O6cyyr7z8Zuh1IvqtocGrSS8qQ+YMhV63cnNK79Y8SEIzGwr0AZx1+
EQk7edQqlF2ebIBThf0RsweggEzOznqevTlnEOXMLHmLKD6yBojcOsY0ZTK+MACQ
sWYYIbQbgKSL45eLnQHR+V69XbTv1XUV7aK+bVd8L434S6fVjJqOXtLjzSM8/jnz
oS8Zq9wnO0p796K6CYAYWArLIlEtIfUgXqhYVi88dNPtqcZ0VA9VvYKZJE0N81RW
VEgY0a0qJWFDE7d9OIs5RLgc4TNuRw/RugjbubMxA6eL9z99SZkY0VHnT85YUEem
aLPHiRlTD3uZ3LZKWMqWT5X3FqLMNBs3zkgEq5QDru/7Bj1KfEI7+M5KkdaM/ECd
1te2xrUYsNe8XYKDhoz9v4g1sd+NcnR9SKfMTaSt0scxbjeOA1KOsykHI8I+NCI4
IoGOkIRCEETAXQPSYXnHcbQWBvTqn0tWKDffbhgUnks9JS6qbAiMVxaBLiwC/phG
Ul1SLUApi/sCQy9dm94INQq2GX9QvhbGDiz1PakDJmFv4SM0MICqSSM2haqLaHh5
xtjaEE6+1NsJH+jxF3ngaCwIZWLkq6wii+L7bWuAsVmx0SECGk/0MIB7TWzFQriM
e13pHOopDdwiIPgAT4K7sqvVae5jDj6S1xG3Rh+PSd0/5hjU8ZZA4E03MmHkB97U
DhqFGm/Vcrb/yRzeHosYOrl1UIFK4auE1TetoFQ+vnlUx1oyhQomByNebnlLwlSY
oGqrzmNAd+YbhFF+y+Bbyru6gCAdK3qPrVDV5lYdGjqmXzQviMGwJFLGkENNB/g6
avELLLmgx63l/0x+dPMqtogMdtb5orzQGayxGXwAgVzGd/RhXvE0kcqr8AU9H4fX
bmHuXH9NKRsu3hQ6Kj0qAvojOOizBJW3kXeWILFbLUJ+EtsTgPS4aLi3vPFjFMxi
JvtKRJDFZAwvOew/PZGoxPs5ufbiJ93huRSrOyDJK3rHiXRnm9v60edNErYpZ87b
tu6hVYi0MTaYSrMfNvKcIvFKMyI/57ieVtMU9CBI4fQm4nlyz3XM81I2oqbbXUwz
bL+dNhrJgvmADcS4YbGDAtkKJMy5evcSrL91whsJZwaf2jR4AhohTnqTYvsPqrQA
92N4qH90N2A7zJSVFtoCCTVeDEyu7ruqrSfuvej+OgY0BQh6wLs00xGMVKS1V9YN
7p32o9iYF/pYtM9oUrM7gxoZXPotRAv66vKrY1K8u7Px+63h5DxI+a+yCKFslGbV
ZAoJzX15pIvvNYGc0disxzoX6W74oD828f2+JK1YfsP9Gl3W0ULSp5aUVsDn7osl
Bs8JwsN7ahJt6tOLnDDn0LYhr8OQs1xwOQoGskoTQ/Dbs5ey3YPYG5P0ZxCNWQ5N
pWkltJudyt/eI/9hlCi5D48YtUd3oGWQz4WGMa9p/lGqEfwKudKaISI+dhyRuhpA
owpngaGH80wGVC08dv3bncnoDF71h0zWIpFrciB7w1JCdO/ooTwkGeoLHk+8N3U0
lzz8BJ259rEMwhtHtLpIAOKhECXTm4MDh4RxvPFojXweEBeJjKTspFsWa4llY90Y
IuEZeEaheUhwxvPwJYU8NTKL/4z0InWvG9VksA0IKVhH6DE9rxCozdxSyfpL2h95
0zGapLQkn1cluJD3QsLca8u1rh8dQpQ+Ac8wfEXWsj7H9blO1Me9C4fF4v4s4zsu
/IHkPHuQ9oJZUjnfiKBFk9cCkK+Pjh4uE5xPkRt5HJR+KKE6/Zb6OgSqi+AKN/Fb
Li1eVu+4g3WjmEgH6w7u+AXJHN/ycmrOSiTf9NPLcyJfZoeuOfLng061kdXWeZVC
`protect END_PROTECTED
