`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmpyfZNtKrdhTpzprpjWCyHng042HwSxMHMTSM0+Mx+ciDFP76KwKYqo8g7QGGK7
UU0id9exvqxf478C+M3fjlxXIPPVYHxDiL8A1wFOSeqmsgEkpwJ6hw04EzRhkkNC
atBy8s+XFTprU87pbbrbJnWkNpiGLBQlF/xtHGR6opFtMuXr5bE0TG+k/xiFiigh
V132LkxmEIJCodIiNr/JKS1AgN6tqP1/NMn5p2Mx6PXXs4EPnDVH55aae/TSts/K
fWBpWQ4KOAV6ZDzqDrtVCWTUQgZJ4rxWfsYx+7ZIQklDUuRGcos+SWD2tnUovAvE
ubykH0DvjnjeJWg5G7DBkxghxaYSCyQTrWv2n3amkxRwjj6POuRN3mu3QVmGYb9B
Z7p08AjjFkZmWw/Xuc/80LJNCyqlzDda+IkvyNFuBOOHWlMT3COfSu7h6n94vV0d
uqTKELelXQaBmhP65sKIPaVL6mu2GpMlScCXwwHTB8RfQEpr/zLZs0idMOOlXuy0
k1khyKW5Gvbdzzul6t3T7or201g9Gvgs7n40Bq6jemgW0XBo3ODROt+jBzPS51rm
PdGfWltWQhigPeI0/rN+BTYwIbtsi8oo1untjxupq3ztWUahF2gjiTvlZ8P8Cx2w
aZWQE3+O7RHJRTUF92tFvBqEOS595K/aDa4AhvXs2ksomBYXAv/C5E8vVp+839Nt
qiL47AzEgbiPfIZNU4w/hQ==
`protect END_PROTECTED
