`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2RIj0CL5Fk5v0t+nSo/nSAXUmo5rdviQfcwBnK+Kj0unbcmvaK4jGdazVGzbrtI
eyC9CLNeTYk8WKM/FBf4QrqkhydCBmNZmisnjD9DRbDFjfS6RBqr0qf3eNVDObOO
O4b/dMDEZVt+rV6RSoHvoZ+NdUQ20ZPTR98DDdLuVx/3dtyguF7hxZUvEkbQZ0sQ
p3L+MlFgnuFnLOKbzF72TaAFCl6tYNsJkolUev3augIWHxcRSeyA5zU42G//OCPD
sAgkEys4fiWikwLZH/0JrFOB54lPwQyoLIXU497FgBV7UXQ31YanuTVjGaP7R0U+
7hJyvTdU5p3uFN3Y+HYFqEI7OxXZXMxWkOhMPfob6ghmIOZPlZZNTRQzehlAmTC8
vM20+DyhYjUGWqtzqpC+P+1mpQU756A2u+MIuZaTPLkAkXlR2Gj6QAB7p+6wQlZ6
Iq+4RUn9xLDJaTTJS+8to59XU0i4yrsnq6NNWThpqlXRZEbrtAUHmv3/97DYvVlr
Ts60Puu6upTbx1m8jExi/7U/NoV4F1bzT3iuVMh6NlBhaOFZ510/J3DeveioBTM2
becXr1tlsgEX1QCFuQhhuV1zEkorIeEdqMnHfc52O60ISLJycVgWZSmZ8m2Ruto7
cxTh1GiUdhtz2NqdWh/po/GDi700ljt1anQ2kdAarB8mtScE/hi2PVUMH3DKTwfb
nLQI5B9EZ9SrKflmIZ48Wm0L/LEMTvLrcLK5VgdSIPAgUz74g7DK6i6puiB1RzUq
4Ithq8nx44SkpuhyUfmxdw+5bdgjhm8I+VD3/nYkteA1BbqlfjEiUa8//w8h4x6w
QiiRn+KCrPlXBZCtN7MPps3tc9elM2lReL7bOzADy9s6605cErdzz3J+NnKa1QKA
UZkyCOYO8/V/+SQLXr27FboJQSycHGbI5D1tQFnC08nZsAtLZmXlrbBTXiiLtegv
S3O/d0XuBM/uSswbNXKlvYJx94SkdcUOcAou9JjKv25duWZhKhrs1AXIOJQ8MWVn
Zticm5ANGO/WUdwc1ZPr67KY2n4TVhsEIuZ3zHf/aqJBgHE7O3kZu1idj81n8APH
grISsxn4MZdMyLFu8huTZL8vxs8U4E4fP4tLS+ORMjSZ40cFloRNhJFAdXTD6FgZ
ce+Q2t0E9e51Hf4BXiiolWjdvpUvMfflrMNzeL4Mn2iBdk9PuoPwLivOd9jnl5is
S/KFY283RSWJVj6GbXoDUEiraSdIlasJAIPUOEyDIa4RUYzwl0WJXzFW9H4z463z
TbIITdY+PGPeErx+LSgVw/tOb9NIOlIpGrxI0UOrd1qi9oLDW92okeu0ThEhj3mK
onGLStsg4DGiRzZZVKtdTsIPlOfQieVciHSnMRHJdtvsVm2nf5349wHI48knhyVz
Gksw87DaMquh4htJ86ig5sUpWBQxDr8KVCXT13xqWa4632qt9jYI+cLzAU1Ylue+
LmrrE7Hddd2BXvzkVBJT5hl1+b5GxmnPjpYyfiyMJuXRtBdik6Bk/UXmC/CM/dpK
FjvORR9GSbpXMmgpgM/I7KkKwq3DfTmoO4WUK0ooZwvsvJYjPilPbOd1WasQO0eF
iThorSNq0CDBTlEC9KQfCvJwrPGuFh4i0I79TGjqhR5S3s0iLobtqP/R1Y+JfhlU
j7U0n1v5w92MRS9srHo2rTJQvsYn/w/p2vZrcWVOjm/2Yj4D5ZZRoZEhNKZyN6MY
UGEn1V74EDCyHKPlf5YYukU9OtLX+FldWgsTBZos6x8Yu9PBTeydZHf+4IGFOFSN
zn92OYig6P9iX6w2x+E/gMXE7ulj01UMkWb2YbVDg+j04NWyt6UuV1raNvodrRtc
wP7ZRkobdhYY9O2OgGU/ubY+20mnom4b58V54d7FyrzV6c8AgWJc0VO7SguOpT38
XXe4SdWivtmcZZo8IDKIEbefph3v6NZGgYZGOvRIcJRn6FnI/lYYtmXLunxOjtNW
ou5MdUFX/sQ+aUX3H8Au/jjLA9J68Cx7BNr13GGnrJmUXKY0lg/3KZ9dnvH9xGtS
wNe3QePKV8eOz2PesuFXcSQKnYCUpa7nPgw5S0clso/KmC/GMVLex6qc5M3Q0C2u
sBFGPIBl+zk3/doeNgyUdk8//D64cmXbqLLvnrLKNMv51eL0H/Ukl3cFkmX19b/x
dw/F4UxJbez3jkpTqyWrPeezMdcAkX1lYHWBqOj6+nHdedWFkvB9C+1lKVQLszsV
cMfA78ghpVIt+c7kqBjMuzHKkL/jRjdH89PecKsuGgzC8BniQEwo/vAE+CidmdW7
ag42cv7QdpzmPHZ5Ub0k4pQVQFrN4XgiGJ22ruJhiX8jJZpBW7k5ayDTUIFY1yrk
GistaAmkzEQ+KpwOQCiFCwz/+PCWIkdXOhSqF/LOOy9/z0s2toa9uFIjP5JTeRv7
RDJF40MNMKhJnhoA4XilpT2iQgifOhR5IQ0BJsiVOjgGAEkOWxWARpI1R6iPCte0
neMx68hLaVKQTYp5ksMaWWQqAT2edtfrSjnzLCKBGDZxCbY9krDrFOv4Kapcchyx
4hes/dR6cZebIjPKwZrzQNGOOXEX421ULfeBtsNkAmft8t55Uds93uqDFjGetfLf
h8gusvuOcvDx7Gsk5cUYQmSDzPmZZzcY1W7fTKeIGr7yKqyM08HFXbyJJNWKDoND
tAdoCvS4qnW7KHzX9+td4SeZxzSaWu27m6B5vSo1CroJyk5xfSx6LtgboxhbgGeY
GISZmyPZ01djLZPf3XMThkw702ZMgRrklAku7fIRx161IZGX+UmtN4+zpLsnTt1x
XM/VL+1snDKfPbpmnVRPBLPbikhVve8OmSA+3tUrpmU0d4o5uuGqpWSl5/wGu642
ccv1tWEtfwIRWx+m2W3l4ehHRVgGxeIsFHFFQhNGyF5hZeLu08bBmIi8p4p2021G
Nc70TCbWcmgEg1e02+eT1ggxkHOpxYIYHcDrKV8vtM+Cn3ng/QXxDg6PuWDnv0yG
VUf69TUgEcXDhyV4guzUiKoWtZSdqztuhn6Z6TOWg8faKCQTa1vKEq9d5dbJroJH
tE/xfnGRybB/cZqwWwYr8KuM+RDKTcwMPJAzRkIzTBzVKAtNvvwymGHntZN4y//X
TGOCmN29ziHL0ZNgWmDcOF85d+oYsBqMVjoBq48+iuIp+b4NGEWLK0lpz5tztZkS
oSDcPN8uYz8VgWtzlEat3mBi7ND261F2LBDYtJrn+01mJ92hqDFOOk0chu87v8gE
nyEl434pzAXFtDqDmyVq84p0Xdi+NE4ZnHYf+OLMj7tepgyoPTU/bVuVmKQVkOUE
/JQMAhd8+k5xfAebZMSPhP5uPG1i7qL77a5dyidX1TGKUmqsuQgLhV2sxayxG8G/
7HpzoTULx2eRsCOszor4OUbfLEuQxnhzKI8QRbeeCElkJWdXdqz3IgkouyVne8vl
1T5f3nSwERde8HxOhKebcYNdXZ+4hsXjhStS+Ad8CLic6i9ZbHNm0GodmcKw2Nn/
a5hH3AXPEjoPaFG24HKzfHgQuktTfnd3YgP8L3RDrE0COJDfGelge2T4ksMQM3lz
yeYKWiT1Hx1FsH++YPxiuozGdgVhJYCp+8qiZ5xmsGfp80qVAjYJKWUaaEjAu7eQ
yIFOmqwqW74p3ePHYJ+KdhW3jx9PLSIphflX0c9uPz2i4ggoEzPAjSZCRNIfN1Mm
8PBBcYBT7E8XujUGKsB3pRuU+bn7oZ18gFFRFTCsbhFoqTu5AWXS0kvdpcW+T5cp
x58ET0GkgFF9NkYDKhVE8QJCRjEsc3xqcYrLYejub2lce+1mjeYl9FO3X7hwWuqU
jDBf0wMJ06fFZjtUi3zcPYFbo8l+NzX8BG7wNDG7O+DDtmLiWgTFjkS1mwZ6L/IB
ffsQ47wIsr2Auo8qvddu5tlfV9SLXIDNp+wyglQuvW9l5xhTnPNjYwiq4zeG18JV
h/l8rpPp/3izoo/w56gACoM9j3jo4+umc0brvO8F4JgyOkjLipvW34MKptLVkhP3
ozxoepeigOsEAhSB63uMbBfdaJzrgkH19z/pWbTH+eCL0P65joV2a7b+hg4lOh3K
tfo9u4ShzIohcadsZHPZaGh/XCOes9ejYfCpEDwk8/zsXUx12xMIjBCRqa594ks5
EcsjiQHjjYvQbdyZupptnThMN7AmGgCTOKeOCGgZXDa/iZiB9fJvlDgl1Qev8+mr
JRGVKpzk7mvYlEiiYQ8bMP04DjTMV03PRw35QS9IQ3aNPVRdteasN0uV8T4V0SED
Ixe6GTXxDySnuHNb0Y62HZ+RTUVPUgT6QitqLaNp8jq0LrNCxfhEur2hF2HN1Jfm
u9Z4Q/fV3GSH97joHeOnoEismDWggl3Tqm73aXRWKo/Ta3Z7JvThK+zw38y3ps+b
APMUuVIITlCfflS8RNHAV7/i8l3Ji5b9lkcQ7IXXl+0fH9B+hK1l/fqyKfyF1mv1
C72b0AcwtN4Js6m/uNQmDlDrYG49tBGWXYhjGv09KT6lUbAiCI1X7gC9kDqietu4
`protect END_PROTECTED
