`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmBJID7NGIEvfp94AHQjKHikRAI1pI3m64H76I55KGEgsyXhEXKm4HBxuJ0bxxqN
g8fdAN57OIZqLcpLHJwLOZbyEwBqIWskyEp5C6//RDvi4BiqFLP0IKnWjuLaWA9K
Zo1F0LCxEg0g5+zc4ym8zMIL1WAA1NiqJU/6KG8wOOIL/Qy1EWMFdKrD9ZJnJkRr
PLEvfgT6q2VpIXzu5+uPAnps4+o/gQyxoHwBZTIJcijQoiqlimsaP0xV4s8MA9+2
OE/dM34eUTq3nuAAL76hGlRShlVaSZX1HYOBxpTwmov9CUulpxyfSmMEt8n16aGO
rFdYY8AR7VsffYCIxloKBjqE4CqGIuQMyrEHjQm0ruvvfPbyfPVa/m5CNTSE7mqm
PkeCeBCDJ0WegtfPE5JFejFwdhWvxJCzIkQysWBDviA3Wuef6cg0vsPrXJz1NKm1
LXJFYDz46/XrGUUl2LNW+rUszlW5EpQDimYUGey1sd3AXKuQ3EACEe8FuafUL+7q
F7rp/FK4XJJ8ZtkYJRTsrm0zFr9NwYhTqf9jqYoaOFG4TpI0/y4fViqKT/BXACER
ll6CjFPSGJb6FqD12OUNQ4n7Ts48UyCXjfuE2T3tYHOy99mAybDvsReJttyA1UJo
aQDIUbed6UJhFM/9Ch/RuROndEm1JZ7x56K67/vgUC0dy0Q4t0rRJnSUlXXLyGzU
rkZApF99+yRJr74+jIHy55NVR9T1Ni29Bc54AN+iHnY=
`protect END_PROTECTED
