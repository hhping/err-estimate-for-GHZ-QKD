`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axWU46GHDwMQqvHMONjH+6wtVp0KvviYfI2Ihr4UH97R41WJVXRY4WYkxyk9+w4c
vIVp4lsgjHMkYcxlVve+UuhnXdeGm5OjHGiMijOzR2L33memOuCBFqYNQ7iWi8+l
qksFpZLlhy3m3HfRGtg295Ilv0Davm0zzqTvtEBLN4BPx4yHxaGjUazM1F2Yg/fY
/ld57QVg+rif7d6kGM5WmlVgXaBgco2Tqy8SoFilkptLYN+fRl6goRnfeVYZQrXQ
MZl1hlQLNcDGEr1D7C0ESdJSWHXZi0Nvmssr0F95CQXfew2KTdMo6hL9glaS9UBu
vsMKTFM41H6JZ3nDVRDcXru/GDQ4Uf6tf0VwCSlzhkvnLxNT+IuegZj4ZBGQgWGV
I6lVHAFDEOBR6dw+A4Cl4FHLYpNKgoC66UcEc/Pnz/Xbzoqach2mPBjdw65Z5d/e
W5y8cAfvhorbrJlsqjCBIyEFdAm0WqduOu3MnvtfXQrSvYmI6yPjNzt3d5/1WrnX
XuM1DcV0KrwgtAeCUfdAuqNgBOlUATENzJvJhBXSYo/w8FwBaoZm99bSTYynmAnA
PhWlToFQZx/JG/tRYAPnlsyItSzC7cfMSTiitB+fWCs1ZvZReRmkGvGjUdpLbx8X
ufFXbkv8g7IxE9D7cbozhkAVWlLL5XKdI1OIPFLDnTClyhqE7wWRtJaI5JQ2Iwtt
siXQo7G8Xj4aiH2IZB7xqPWIwdNY32OB6EVteYyOtsNZLaJOIvkQ/PHRbCyvlBak
EKy4OvCY8KMOskTEGMxUHnUfuK4O8SpAIFvQPqM5bukUPVhHVJHjd3wnlJXuo8Qw
T0cyqzqkPLwy1QIbggluUZjr1sXxRg/6KRJ9m61P7DYfWvmM0c/sNOr3QecNBpiI
6NrWQIDBK7zowuArf8dJ8M/BmLcPE0qz470os6mg4NT7oyNx49rZbuhRiEANG9ir
5FJXM/L5dK0KedZqcrF3lqegG64Ln+hv6CFAyYDmy7LNOujtOXG2kUZ/ebmmuaKg
z4fP4e6HE8BNjGbO8jzA8lIvvS8xmavDp5WGdM0iTobv2xEOTChozUqTZ7VDbXJE
RwYcU5S7TgOqcBW/YGD9YgLPM4PXjUflmKF/Gkvikrlzs54wZS4kpKyreCqArN1P
fKk0imllCOQ5qLj2GN82MDMQ6VhdGAkuhXMHSOQuDaOmVtwYXI20gsO0W6K45WUE
KLfe5a2QTQ9N4FHGX5vZnTRgSecm2942WU23F5/rxXJ+vdnMShTJsJ9xo9XoV8+O
PsUKraRqcaPfwNHR+TfXmkBY2S9Z2WwFne3z7wMeRU8zBcTt0/ekIUk8a2oJfmQw
OZpHK0iYecvg7FiwJcXVeLZheOPWCvRGAuvzWCFqtPshelc1vm+xBnLUKU2qFEN+
xuTj/vDz12Hgmg83wXAu9SZ2UQNOjFho3dAFl3PqlQnL09b7mJk/NWu/vOo80ycA
m0tnz/HEdCcO65fImzxpTugbPYK1pL79wqk4RwJgAnQ7z+QibHoyP2TPfd6kXorz
6Koc9K78ufnJRF1dQD7yYGXtHoyD1694ZQ8puci9qPsGbK403ifsrSlg1cxkRMCA
uxB74OV3OQ81teWpld0ZaPJtOK4lmCCHeR/eD0qXPV/y9PfM8dAW6fZgAids7Us+
brkNyTLRli3MB7xM1+K70+/ORi6jO1osRkZ1aCZNu0Shvhwjvy9Lu1dbdfRr/1Rs
ANmDO+3UFE44MsZv38nv2WBR0kYEn0AS7Oboh3V1GHbTzbf7klEZJlmQAIYhhFJe
zca+FeHTtV2JrOfgSQEAIorK9OoAe7sulcqitxMd8kdUV2N2GcnC1xeDg7Ok1W8K
qmnpVLf7B+vuC5S+sPibO9fyWpPN1nrhrH6HF7tuarPmXKG9yLqmZmBrRCxn/mDq
pP0xZOyg8wYkApxYxxMnVC+T1tEg9KrHa0wIBE6TjzW8UfJ6BHch4uYBLpQvkn+L
f+Xh79DQEPi861G0F8BZzXfZKWowA0WiihJCw3l9DptdqJNKhlY3npkaTfM/4NeO
AfgKdLmF7eQD06t/w9LnomS4w0FTf172I+r1QK+CzaqqVt0kTcmzlt31KF6DWxW8
fsEryVolyiy47eM4kBjHIvgMoRtp6lNflGmaScMls08GjBpeifLjsgvuZXnIPLio
gpVl0DM7zc0UzL41maYHPOxG6zGPNM+fNGsfKGyKbAoXgwdiRyaKDt4aqzrB80PJ
EnCXsV1NAPTPlElZFmrIbDYC/j4mdf+5cZqcQjNlnoDPOgEP7+cMJnXJbTJ3j83m
Nn7z8UKcWfVD/VAZBol4GlwZmG33eRqD1pmT01mAmxeBppPFsOuZukT7MYj4dYnr
TosdaIotFgvpj9QFxkVCCKWsEWvm87KaamijUDU0ZSwAHr10tyeIxxJ0C9SCjy8S
wLhD8LKLDxpT9Uh1r5OobSiZvMdhotL1NFCGZEDvgrkTEEqzczHLixfoGABm8Hee
D0OSKJUbEDgiUK3LGwZXvEmaKRqnxjp7LdgPM03RyDSCLXSJNR/oHF21tEmSjytO
3ud7gVoW9PbaSHuYIlQF5bk2VGNTMncQbYqA7KVw3OnaLzabT0wecsmdtO6DRYnV
EiCnDsd3mY6hZWMea5bTeg==
`protect END_PROTECTED
