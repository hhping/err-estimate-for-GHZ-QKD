`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLULIqWfBNv+kdPq2eX9wDRcutD0yExczGGIR9t8dc69ICRCZS1ZpPoLJPBfawtK
4Ss73B+mEexvHr978TxMUNnVsfxoNe0xq2TEwATkCScijCcTQ2l7FFav6XBszzzv
KaWeN/+hppZOHDPotbvKtWkTGnIaudRI8Pf7kLRBiR6gXiM65tFGiPVDpFSp4YcH
JDGJbLSnJMesl0feBN77NfwCeYn8X11WbYNHaI3Sas611+tJSfL5tQSCldJdc7sx
aMB0oq4d52aZCJWkyxtc5onXyhWaBvXi/L5qRAsX0QXu8A39rNYRWx7vKVhFD1+Y
t7pwJx3mVqMQ/GQ94O4k2YYKyQsK4KaCQ8mFi9J0MyFocYAFebE2wJzOgDy3th8H
73Mxxct8NKG1ZciWH3Ntmi1WF31RHc7UmSVlVWsCJ0eSgTpZ876MPoLAsIIf5lQR
EondqiJmU4XvAkhxlzH3JhgyUXzUXYRtjh70i4t5/NUa1imhG6IpiBKcDsjdbf0w
BS19hmF6O7Tdn0wuoyP+2tNpJ5urbHoiQLzGULIXeZ3iFWZ23648yeJhohzD/SYK
sc/FvU4z+KLoPwJPbktouVtRAI0SrHvur537ocle5/sqXJLmm1mTjVBIWAHrop3/
6OXJuA7jX/DXHztYsQWH4jVSvuY/ARNeXUilYUPtWhebgeLEs86lvN/Hh+N8ttWb
lwDlF6aBYFLzGd4ETB3p9dtEhDar7/JKdiaQu09TWJd2XgRPMweFXHuYVSLvqlvo
4qgXQ1beDF7BxSRTwvX2rm2iIMTExZWKskPssv4q2Up/aRtTd4uGGCDEEK0XkXfq
ECoaghN8jNNP7redHhJC4Gxg/RMYc5ndeBQrvqOk0SY+FZyxjSCk/fPLYvGU8f/m
MWfMpNhwi5u3LbZ+8NCOuuB2sYXvPwINuK8yqlrxdqzJvxNBj74L/iX//UxzU1uf
ra9JEVU1tsVHUZ/loWhfsDP+SLPBhx/SeBy6kAHH9sx0+O24w61ag7nhOgJn1Mht
oyvQg85+RqCJfHNmOHZRhDu49x5K5QQXZnw7PXhbIa6J1PIhMzG3YAxZGdca8WGq
p6lzo+ednUVXuWO4Ofo7tizZ9Dszrl3LosWonGe8q1MjIoXRSy32ftkx6z5pOp9Q
x5eFKW/MU6cA6hVG45ngxMG5JgDXawsGq6BffCCRTYHbCojH8Zz1PMkgxLdssI+w
0XVMXZ1dJ51Z7TlgY8e3Y6UNGyRJz2q9+L00349CiSwoq1D7NZz+1GQqHjsyZ4VT
36iI1jNIL9mQOEk8jgK8V0NLDJHiujQui2T9ON8Czra7bZmawdxDYKrStvgHhq8f
t/5IgjqAhXK87DgFPY1M9rkrxO60HtXiHFt+jhUBCtbvMrFY4N7jBrSuYYTAcIa0
noskfZipIIFTsi96qsJ31xZGUpmWAklkSHSxbiyKIYGpuNWrFufdfXPE06+X7AhI
4tKwwW6jgq2oEhqHeXwNGqx2Tm0UiLrz1+mPmPELrICut83DINRSbVDjHCLieyyl
lQIo9KX250U49/Msd9ku2tkLc/5kmnUc8/pYDGa0X8Is+Md5QSkZuyuaG26VWolQ
azEDXc/89PC+iHCBfY1kROr7XFpxc59eA9VOsO1v9sySn7DGeVC2kyrdLVIiA43g
cQVhVS7JnQlhPrIiNrMOspCc4Thc2d/nmS4HmGog9sTnTkZA8po4fwPj592dvMD9
DF/KYL/ZTz52jivIO7tVE85FYhWPZiLL0ERtEldu0k6Zf8M3XH/Bx7q8Nopn0VNk
A7Qo0jfuGyJ5kb73FwgWune07wQl6oiuQfLRFXLguWC7flTi8jrzGQwvh9L1S7yg
1eDr0dlQs9HeWVqe7YbzjrhiDs/q37L/VAZvVX+Hp/NP6Sct2ZNOG9LFdap5urnx
3BOeWHvykubQivbQQbbJwPBMZbOuXf/b2Sx1fxKDqh0xVMVmBRqLBjl23ZEjfAib
oERuJ/UrH/+/jj60nY9fWf1BUc8ufNeXmiMYkVG6uOEL79rq91Sw/1nN4s+4PRyu
y/Eb9C1gFSpM58LHxDolfpYBzNTu8EWyPUvI2CBOMAr1A89jryENOzmHpnuO7vqr
ZdV4P0EcC2eUhHX4NVVrtGVlvclAwcQMZE/bqsw3Nd73ZpAu0Nm3D1qIN1lf0GZu
9XM1lSePiukXjxjVqrdyNRA4xMC2PmNTdVtODSn1/Tc9d/b6OOtQYGCOx7+D4Wus
cSydKixR3RNkn/fiPNtGy4K6OmwG2bDlNrxHd8sddD7gXJEzUMX3Rp971kBeuhNJ
706Ya7YRenR22KAw2QFO6odpn4V/XC6hcvM1qzDbP3MGJV+2cwqcR06Y1yTNEJgS
VBNmsCYk5oemo2myzDxxs1HIJxuVy9MvCnzHPC/Lt0FwrFmsbDStls7ZqQTdd/Nj
szDcLJROcEY76L36BorouWK+fEkvgCmnTyPXS1OSwuhqTxBnK+RqjdFSidXmlnlk
IvJjHqlGcQkup/NFKR12T5XPwRsUCqklo18cZJCjjH0=
`protect END_PROTECTED
