`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pa6ZFnrM00Vz1dBi9gpKO7TZ4peCvL7jaRLc/49FJWP5QTwcZ2xblwtVLidUP3bQ
+IO2cX0trLOXhP867u03ASXJq5PcSMgLAgWWJr2QlhDLi/4FZqhUNMOyn6dP9bVz
P87QqJbckbb3weu+DLflk7HRnl1QhUeDlCWhEy2pBZx4AW7iZkzqMoGVF4uKJqN5
fe7Zoe4fHU/z475WEUhTVx4MDxYARVjSSnVGaAydrohnzmojRoyaoTYuqAz5277O
8pXkHjge7quN+e5imlMN59lL/G+2TRN7rneuoTxvkgdyxFxiAgYYic7CFADalY3h
wde6lvSlKtWQPeDF5wOkaZcWUJn50HqA/WGSkJiq0yYDPLqnioJ3DWqS79Vw209z
H3FJw4kAxxLeP6m33Xxndb6EKTYN8tGyQ3i3rH4cY36qfr9zo93B87wFTRkZBTIQ
3p2Ui4taY04d1+6azHN+TwLAYE0SqZcWxA/dQpnffMF2dWxNup0qc0pO0C4VzA8K
70C+/HvNlZFUrWBs8P1UKy1Jtg+/leU87Ul4U7SPDeIOSLv91HP9Ery4gSBzekaG
Xwf1XaLHVNVGp1kTqV6j9+JDNXyGvWyTKJOyrxMnBAJfjp3ZrstNThR1VEOnwb0N
G49Ycw9afCjjpKXoeEQ202cIhxGNlcTuUxqj3OeqbNejJi5QRPcy6KHhXdHNz9/E
6XQwiSrh2yyEHwOX8PKjr+Lv7xAH8m5994RlPD5+Fh22FIBCrQyGNRGt6hBEibrZ
KnPZ0DE6hLs3R1BLzBhFD+TGiRUOcASnwMVr9IAKDVk7xElVISTnPXncIikAvP+i
mBPigKtyJ3txrsExt3a5Lh7yAgh6hmBxri87oqsfWWJutkL/2dBfALSrIeTKmc+J
ucYl2EQ1TMCMecBjTrE/Qan7+9L44T9CXHe0zTCjT+AIbxuZXcGQ2JRWxXeSYCW1
ycN5V6Sw3peYG2V26XiRTuurWYuiuPLXPOm4tG5uhgrz39a8xGWjDHJyQDmwB0q3
5+lr2afFjJaqPKB3gsFHRlayrb6uHzbROhKrR6gTLqdOi9R1gDjB1cn8IkRV2uzZ
`protect END_PROTECTED
