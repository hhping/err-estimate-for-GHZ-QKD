`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JmUCNmmjRSu9Gij+j47Pq6/mGF/3FfqGSLSF166sdI2AcLCUlHNCYBNFxDYpBGj/
473a8fLBPUVrLPwyDs8Kw6nEQVytzuKQY6I1c6l/AdV4WHGQbBVa0M6G++Qzw7l4
70xLhAsXM5/sj29zM27jyNDj2EkUXGfmP2tFAPZlLIJYZIQZtTNDbPYPERQJejnN
MFdIroPQTd3HHDqUzhJ7YD4nw+NsR45wwUSYk7EeygvP1t0Vt+Apki0/Td7w6k4p
a8FZfCVJhgJM2Ms0+bIDItkimK1JsR4f0HbjNeNeY5OR4bnV7SYcNyCIrdu8XBBA
3R8OJv3KITzPf0u0S1uMZ3UJxHSQxm2lUTyuvLU+5VI9YslnqDYsxUlMKOxqclNU
2ewM3hmt2xZ2oJlTnTu7c2OAG8JNv19SPpl05DtBVZEslwdNNTuJsrQKwKRmuODN
rpamu0D18MzZ1RbwRQbkyNmKnLooi1C6bRTXg0C7WPOjEi9uRdqli6JFGPfbfEMH
bxKsH06hmPGwWJkMO+Tdsx3Y9ond7VkCxk8kieF++TSXvEWOzpZdtYm9CvlT8fER
2T19rPT44jbU/Hw4vzCzrwphl4nr18JmBPd6/MR5sSCh0Edp2VMbnIp70pFy+0Pb
JkuGj+bTL2k/e6mXeXMBdG7mQeWfwiUD9DagWxsofXO/oH5OrQNMovSxyPhJtGXO
Y6bNq0sV1Yc4CDnPumAiv9dGV1j40JYgNPIqf83FV0AiJk/l5zfMDi8skufqoEQu
xVN4ZVDkCtQvfqNRNn0A3lK48zMeNzXGnimRQgmggrV60vOwQzzLiEt91NleejgR
TaSJ5h9Xf+WvOv1WVC7SAqGfX/dH6MZHrILyqyi12GX7Az529atYctU8gkvgilxw
XJROOS/NGdqu8nap/cjDVyaAez8hGEuaSe9jE4cWF3lXt2ilt2ffBRjl2UZBh9uJ
waxfB05v2UUXVBBvdUi7zA2Ny5iddg7a72b/3+KJ9gWBSx5J6sIZFpvrYuU28f2K
MA8uoTZ9qb/qtOvWVj+qqw2SNTiBFr8EjIB4PqPL3wlTIuqEE8FNckv57uPMnxY2
EPOsDHUK/MbxuhzAqI7/Y53ahtw25pq8rAKFQ8+iHTi/KVwvbirpo6HLebEVfxj4
J2GIG3DrRlieD7EOUySjPDtO1Hh5CqRMahdemOahBsdbnj6St1L/E5OCVCU4/7ha
bQ8EdM4YzZHdKEPzhp+iRsrw5sN7HBFYyHoP3BA9jJy6tola1lBUBHO9eisOssQd
b+hdfWg3U0sjwqa8DG1O1j5nMZHDDp0vfAaoJtKR1VUmFutOKnbrTTz7snKerjIg
QFg7hzt/b/82Z6DU3UpAPiEw0KvZV0g7iJyzRZUJgR4S4dlcUCFn7Rkl1lejccPs
azLbcsVxxwBt8kDM33QCviI/aFHzM35lyTrKi+qFf8VmPWdtMQv/OpfoGes/dt73
wOOLv2ND1oXCdwTDCeQAmkZ/Zs8ndeE9MWGzyuy9IvpD/mz/J10NC8dSmbigim0F
ujt5OJiBRhwKHlxHAbdW1xmVfRPwmijscf82kqH7Q1qeUCR2KTqSB8mytZtgUcsK
4PlSwXgkuvqE3+ACRzu6F6QCpLC1bXbcZcz4/zpzy3H7jBw29QmVRHP7ZeujptL9
irVs8uSAdHRPbaHuIe3sEpGBXXngjCvzcZg5fFgmb9SgcYnJ7GFG9XodQgW3RLAo
+EK1bYXldw1XBSFMmbfK3w5VbHCki6Qjf4GEJgRQLp94PL4Lpq268QdBx7ZeEmqU
sOmfvC656BF6XYazWtiALgsc9ixkEe1YgqgfyiHO6P+u/9EDWLfjBJjBnII0ue1m
F38pSG6Qrbxwl65ZZVVA1tsgvr01xZ69yzq/y28oKG3bzHoGNP5W91SRIh9Pq1hq
SUB2AkDvhq6ivF4bxbXeEU95cP2KNIEQ+IDr9wCRyLZmBGTRyoW6TXCcvMh2JGDR
WwK6fBxibNiMjuakT0fX589r9d7U3gODttu/OmS65Y1kOuP9gWKfPqGT920LND67
fK+iGUNWNgMafdUG42+jyn0oEbNt9pUXKNK1O3f5hNm+EMuZqJBhEEW+vtB2wvjB
L4enov6aQDdtLvUjHn8CN+L+XN+dUnFUt6fgNvcsXISJt/P/KB3LavDZWYwKpBKg
MVcp7Ai+HiGsS0iqQSeHTBd+zTRtyRbvtVjmE0u30oxuqBbDP3xJ3GPVrjajBGn4
P6AjOHBkMdfc/m0I2c3PjzcSiWtHxE/rAZfapbHBEWXbjZ+rxBle4zf+EVIKsypJ
ZX2wzh3oeV4x00hFawGwdyqc7gs01cMdelEhVR+rLGw8Ro44R+4PA35a7t7FLln0
+aGyRuZf7IOC+viUYuO1RS3ZUOlRR+lDw9dU+p/oam1kO05s4Ebxsuobt6pkCkQJ
P4fOYSnFSe5ojg2VmQ0/WG6ckeOz6P6DSkm6z4pnHl6eciIqHOWRMuyaExHQE2z6
oJhOHlcw7ohu67nq3PgcGSiGF9DKYP/JrVKIAz4vJHSGXhG72ESBR2lZCQ4moLTZ
7bjKGTsrOGWDOZa1KUSHvU/Xc4msx6TJyttm5QaNdu8h9aIhqjQRBr6ikpxMxUOP
K4u3VDNA4epdOrR1h82EnwbVgZPiB8jfkmUD6wat0TUqam5Z75aRcUSJJ0xGTqRu
jQfJa8JyglFUeU4yuiB9v6sTLwDBQFBd8LN6n7BMw2JAURIB1JU40GPHmZifVV1z
de3M0Rc/VZImTP/QnnBqY+gu51tQ0LOta6pPgXZhkSHpH0mURwdtR67xiVU3nt+S
UToNAoe7m0lHZst8Atzyo1vR+zx5mGmmVQGmyaJMkbD5H4eNe1Kfbh9c0+OSfO8B
LaQ5CNtN07na8eLPsb0+bRk5m8y0Y7w0Gz8N5+sWoz9FogMwF70pXVIEYBx/IGG1
c9ui+iRd+vK34P3QNHd1tDo3RpxYhL+f/QXWLduSon/8WDSzuEgLIDyR1s/k2EnT
oVg999tZZr0oLTccZaWfuQ5wk4J/zpBrDHrEUVobgvGlKOJBhdW1ixFW6OhaPYRP
Al1tCkQ6wtU4rUy5A91b2pk5FNqZcVUmF48aSe7V2TPKa5767GD/suvniziZgT1A
pOnfJ/fpXRzY9xLSzIylqHLsrVT5pbx7+7QCvouqhHNo3b91SWHKHWFb9RAfEvjP
uItdwf3FKGVqrlo0f887NJTgo9kuIa7LXC2VOqwbN2vZzVYUbi+PnpYBjWirtLIm
emu6C0KNj3KhBjbQqbCICx31rhKthpaL/u2c98U9FhCUqrjozFvlyN/EsD+WzxYe
59Y0og0zuVWEeUyYEKzpsZA2lsvMgeUZBmKZJ/VcGS0cCUku0HLwggZyD5HuckKH
my90sO1ZkbufI08N5yXHApgTgNNTGgpBKGzgk7bLwQuDGZUsO9RNbNom60lpJi8R
wXKq9oPPD5q7YnRPzVpCIA8HIbxklccQELD5YDd03Zc=
`protect END_PROTECTED
