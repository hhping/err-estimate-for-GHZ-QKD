`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Di9W9zXrs6g0iVlmyJ03/sbbB6ixzqFC8OLnLm3GGpcYpUojaxbStSsfnEo5c2O8
Bpf+0TxaGfkgLXTjuaPe34wGZLZVNZ/pQiJIOuXsnWTsWPQHSzLw0DKwRWS58njH
HsY/qoY2QsauOsq2vqLLbho/cPKZcw9bEN/l7/dcGSacFDxFgd2i1/lPXmTq2lf5
xYXB7lQh+tKdIZx6EUHthjNf8iBpFit7C0yjwyMEzetm5HnUQdZ6vo0tfit8G5ZM
B3BK7HtlPT0O+U+8gzIrsiG7J2XrA3qyYSnuQ8Ci1GRVsujPxivj+xocxZsvjD39
vpcKoYeTeOQ3v/eUfYmW9qpzpRCp9uKLs32tkaFC7ZxsHb7KODbR2sNojLKIX6D7
tK0ZgJPzV4DLKb+XzIFlv4iQ+KsN3gb8F6Y/OnmYoOoimcKDfDPzZ2I+Hcda82k7
qRZwK3FG34JpMuUguXb1YjybcJbowDLXyS9/6m76pWJmFrnOGf+i5AOxWOJDUtC6
8fMlehLBNJsDzbGF/NsKAFowCPTLVnftIL5S+0s8O3o=
`protect END_PROTECTED
