`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxT8+zMTySuBb0dblwXIh4E/IwjZPcZhFVoGoF96mkYsV6DEY5u/Egqqr3l0xnkA
Aur2VOTBaiEvbhT+6n6547MXDhv2FURTlwZD3Zn5A5qrqw7LnFUC4c76jBLlBn4c
I9e8rbmc2rDHoU3B+7J4cjz0Hs9UgYK5/HjoldZWPynvZ3MQOqw8IuhW9xrWr+rg
iF1OL9FP9aNXW/xrKq9U/T12J5eaj+EqnhUU/9fPWKzDai5WWI/2cpDSEu2AkI98
1EMuWCHrUA1w4oEcHWdfMyQWb0EY+njhChGViulbt6bef3ZYzPTXYiwCm2CupruR
htm192LnLezhekuQDRhs/WEbEU6nBsK4npNsrvHS8FVupxJ0KLj+9kMHeBrvZL2h
VHPq4dKSOlEE+HW6LyZwq/czAeaRWnwagr84MSqJuA0ArSkpjTuL8LCu+1obatuI
qSQUi8QEI0fHmw3PvxqNO34s2m9FCPYf9SiQoL9z2qgjFiQHC0SYgK0y0PDSzw2G
DCMFbWNUn4+E8KODTH3MisO+YHdzZVSA7bchwTbWE3MBnbIEQElQezyjQPzdytPU
a/GGWtnlfZ2XXJApOhRF+FviIsVhgK0oiN0Vbx2oG5edQ+2bqQu83eFMz0VmxdY9
rC0DcGVSiM2zD7tYJlQqOtMbUfo4CaGL33JAcvXCz6v9ryPQQPG7xa0ZwbbNzchs
qBU575OUiLy9AHsD+VafyvIJs9uSbF/tN4QLuv6MmIZ2E6KPqF1rC/Zl67hx4MQt
HL9RpfIXs9+hBVd431NDV31lxqWpILECQo3w/C2O6frhQiZlQ8/6YTLAG18bJwp3
LP7SlUrZfyKlgXut7Kx+JTkkoNDZW+WJYFyTBqWbJ5KAVYbET4VtnsBbYm8OV2V2
0vHpbtXuO1Uy8E9/i0f0cC59UQpGSx8c4KjxWe8p1iOg9bLJJ5fYZZLYcMZG+f3A
aK7d2Iu/Ic20pkR2ar/yaRxzY4hAWRjakNJ117qsoa+pS1kriVviX6rCJ8/E0XFI
/2KkgOZODVevH0XO7f8cZp91RTaGO/rP8QDk875em+F86uicGdAk67/FcbvEcFs7
bEP2KlQTofsTXSjl0wuI3p3fW0RuEDR4EBY//xNSSQ0=
`protect END_PROTECTED
