`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdSJYx/wpI+IljB1YdAeNBvv8BtbrGBR3gZJrErrz5E37zgh/9HgJsPrLfbivkav
e7HJ0IAHPZFUM6ra4uF6K2LlQf6uctQsYMZATXtfGwL9KJEFJZtiIqHf9fwyi4hc
jpIAJtniuzfq4M4W6gPtKoH2TcsXGw4SjmqO6CkwvjEHm9mOtoWYk77mG5ZNxKrC
UtjGIzDTB8Bmw4s4OuvQ8U2qmnuSxutFci5ars2aalAGf9C3RXuJnqG/GF3w6de5
gntV/X6ieFKN/eNui0c/aPtz+bSWhpXlCY23gMplhTEhLcewkZ8u2zGdAaU7bmVJ
dHqAhBNBPgr8vs4Cd32JsjNhaDkib4N5FcGZjEPDX81aqB6kSz0/YwRYua/xy8H/
jOg/ckODG02q5sOJbaTmsg==
`protect END_PROTECTED
