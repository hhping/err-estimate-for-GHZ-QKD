`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JzR5EGUBUKc8vAzCqiLYVegxUUKJOBeYNO3zJKhS/BX+gCySvEmpyY/lBRx0Gm8S
FaHMAhpd7gm9A27IeniUqTOLCPbrySnkVnhwoqsVDv+AaIftfAS+pqfWhrJRDKJd
FEwpt1SrVongGvzf1omrspB9vra3hdZCCvHF+DsqvnScz52heWn6wh7Qcix/ONDt
CWOxrX8r3oPQmRBegWmtEklw/uwvTSEBYOvdWhh81jYn6ZyJoATP94UXiu3oI9Ku
mooRp/wmW/m0t6DH+oXTlY+4U8ypbwAVXYp5OwkZ6SnCEYxa7b482EyDKSxjlIWw
8VulGMMNyc767kQzUm4/FloZ3l5pwZodYpOcoUwyHTat6v7bP/UYJlp37h/9Qp0i
uHW4HQzyAR3QYu28MzXlNQPe1QCcZc0rGmUdxwcN6bdur6IRu16DNcWMmcJm3cUT
beg8dXCXTpMnF4vqZ6DN/jPrv+UTBScee0USd09d9EcyyMfiIEMdVMwzUq0R4Qxn
/a90a21lz8dGL/TQvrb/Ww==
`protect END_PROTECTED
