`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+ffvXvWysxUpVxqzfFAdKGAABYA/NvAtqvNDxLhkz28o8+UxvObXCOEuwwwR9uS
3g55jIX87DvC8Bm4Agyc8kJ/U7hwzyEcxN4nfffDczXMBx3WuX4/Ilrk8L7gfVPy
Y0kJ+bnC3rSzVDniGFTPctIa2IEI/CSRiheHWKJ6Lh6v3/LV+AG1jP/Y+JuIoLz9
GX5rvIFYGQGs8C27hkVq9cMKqUDwp0KiSEVBnvX2jfKnLF+6IaJnVOi5PwQlcx5d
xQcgS9MQfGfsqEVr9YknNbVLg2yN7mBOEmklAKYrvLFLMznFUUVeVCRaSX6DYppD
G9dnN0hyDGZlB/v1lKSFgfhx+A65fLI73VXB690R3SgRNqq6n7cy9gKhmqyWVuod
00OhLCFjgtTHQTzD0jgJkvMeu+Dom4jdrDQUJTkNJ4pEp6GGne4MucsclS03mcc6
5vuyCQT4YxoroS3oYJ+XcUExYTuJ2Y9EFo2HHhRAj5d5l370dhP8RRhtHN/RuiAv
/VB7nCZGhesc0IhiKtRKBt2WrJ2weGIqbxXqzf21TIh9onFUT/tq/yxZfDwLEOMS
GinoTqKh6cmVREvCb+nGTnTB5/faYXeOaOlipIo5vqLyZmA3nAS+Lbk63k+IxL8A
FIDOFhg/ZhpkhEiBCMG8bHrgjow++YPMTRYYs24ttbKRD2fj9STYQEJ5zJ9Lo9SU
9VAGpHYnOEhCPLd0BsXdFtg+svOentYnzzydVFyOtAfwiOssq/WuShMg9SAZTMoP
IPziusB4h8ZC0Op1HFQLxvXkJHmyiR7t/pwYDBvDo9aUjltLMi4ShnssdmsiCSTS
ULlQZjCCo5WEo9nplzvbmLvN8Q6/TZ/CPethAj4ssYxeT5ItXXleUw/8zLEpRmij
pwmhz0WEztD6MW/brnKueM1egusg1JStToFfPmbZmlK/g5O/0r+tiXro+xwdBS2B
fMxSM/b2DFuC+v2PPCjdr1n1A9jaX/1SiTH3dCyUxSM=
`protect END_PROTECTED
