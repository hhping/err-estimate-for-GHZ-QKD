`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXLHJB3pBaez+ZPpcWAYAM++NQiqwy7xnum5Jyf2LAEm7cLZtgkLcB3Kd5PdUnHZ
T2WlQvOp2+e4x3XUK4ApQgnnZS/VeTzLRhXmQxqPKhRb3ECaPS9P7L56lN4XRlcW
7rIaHH56KZOZCrb9cFVpUaE/c3QtKy1Ag/Xaur+7NQr+Z8Rx7cxA4G6AE+WHlBIO
gnat6T3zJKLPj/tMeHMBLxAISKuWqIlgzfmLhRzr+BVyucPfCLh7OqY0gmKVjA2Z
2JWvtzitULnTH3YHTkEBB5np3dKF2ODZlpt0SbvJk9kaHKQH++ieha2q+381plRo
PuZ8pFyPyhTwnm5duzUf3ZwhYk5z8nAhMHkhwmxXUmjgBS6kDGc/cbFf1ZGZvUoU
L0EN7AHs/hd+WTzyEge6e8mh0gQMm0nOjQv5vRtk33cBGG8L33bMw5ufbEuQoXsi
Qo9CyQpxvnzo/7w5Nh/YuSgEiIleGR1qPF40xp6kgkhCWuQ1qWx06GyP9OpEXh/r
3gQIlDXctmqM+ZRUiZnx4/5V7vb0aTpcivVigDNNACVSXJbagwyYLDf75TKbe1dX
vzR0chkOap0CuRQZsTofbQ60KCV/nncWxEpoaXgr7QGg6KlXqql/p5QAaEMFRZ0I
zULdO+1+ec2mOKRUS9Gcp1/IrQnHbNe1ZzkFsNxtivpUnhfNg6HGLkZYD2djea9G
YSimPcr/usvczV4HZuH9GP5A0KUKZl7b7RUkyGGF3yUkJEDyEU3Q+WTk5Wnqzev7
hfFn1eFrtYI5oIEl6BSpJytied3wKQSZ2Geem/LOjU1UMmVvM41TwGZEDF9A32zv
fmXra5erO9P/ucOcfBXd+RIQ53RsG8cvNmL/c2p1dFxwXr/SF3Uh1hDAmgIKQSGn
`protect END_PROTECTED
