`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uDzkUEtpZ9RRnKkTucWvhqMkWVgg3q8MJ9qVO/PJzGvFeUd4g7hFdXlSHsYvA7sE
6HZwhjof9zK1xozmEw+9V++fDtjsgyeSvm4AdrZqeQVN04oKlbRp+4Jvd9AZ5l9I
QV2c59/57EID2+OZOg0I5wb+x/bV0UJO4x8ntvjUva7Zv7v2dHZfQzF+5dcf77Uo
8uKu3XVA+NOb543n2k+MaEw77QB5ySX3DQdgcz5bVyAkDFWl90iQWGtQalfHXC+i
vMLywYewrACZSqqZR78cTQKJlhmsM9msL7aR37Cqv9lkjg4Skyki34qntFup/zsO
F6onXgCa6/3pu56x0E5/ZWMehKq/7OBq4cNlDkotctsngyCfhOz8b5yL9ykvSn4p
Tpfv/A8ho+j6FWeH56TVCBu1E4bncjC58EuUAeFFJBiuVgC38K5wDMYS0WWEeqbj
E1qpsKZkICS8n+IV4xFUSigxcWBqOz5j+bCSaJ5sDjC8pT0SCBAwG/6O3jPJrMj6
M/v/wJ5X6Fb2l3JKIfynX/H/GQJW1XVUaQmCECHlagTlbg1sHx1lnBdqxbWC04Dq
gVC4fCXFSVn31t+G0iHS5lKVYCpmz4xH/xFAoAQTtg4cIAHvE1lnAhshi0hmGj18
tOHarCuBNPzLbFeSVjV5Y6jP4OlzIwD9fLQtCap4LsN0LVjmVxQkeUdJpBCKmQiS
C4tShWNHJ14rgBwRrqrNa6QomtoUbL3hbOdLCQUNuc11xY8a/rVbctQwkF/p0sDM
w8+5VbvtzxRa8Udg4B5d0cbvtUidJS3PuDvRObJA2TOi53pInagXAdZcjvZfyxBI
0NHTqeLCnfEFSLhMevqU6wjg/d6H3NTNIHvuftN470EjJx+ibMGx3EqoDxqmBoQr
DR30TdM3yZnzjp1U8SZQ915Frpj3er5Fi45E0OORo096wYtRwJSEUBBkAcvtNeWD
96cPJeEqcGys/JPveU51NwhDgwIwwqhil16M32cok+MrSZbWxz1kFYjOd1kDTXAG
MI3eOmBpq7ZOomkSu8Sz4xftSeY04dZkY13jB48c5r80nQ/vv4sdC0waH/pxSRjm
v9aHPW2kzBGtZDYS8l8Kkvq3T5yba7d97kjq8bD+UPcapA1J9Q/lvQaQ4MdjPF29
ijHjwvneDf4/pgHGzg71CHYUwpMhkCLJenvO6Zz+YrNhTvqdS0c4gvep8h48ji5o
rAxImh1cqdVQC5NtD/+caA==
`protect END_PROTECTED
