`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ad5sKmOapVC+n7ejaaLVk77vWqThSs8rSvyRyqtfj70ZOVVhplay0/gzmb11l+ir
HmW5Fmqm1iWYRKX5vNmCEcU0++2uSWAm6gEGzwnP+yjTimyHgtCx4xQbdykrSs4g
lP+8Dd4FBw1pWlgfSEYfv2klGaa0t2mHOsqHVVRHorF36ktuPY+eVFAYjoydhyRl
ryAYU57PNz4TAemBeG38UoaLjJ1BGT+q0OkCQTRosvB+RFxmKzHVCnNMYXG2rWN/
2MwCvO+FDqI0hgPkE1Sh8Hd8UjwQMPLfVEdjbr4pfHoT2UetPVkwIBek81tYokKi
edNFyrjqpmoJ+ZqYMiMVVG+HD13+tL3NxMSoYp5Ues/m9kjZZfSDsJs5Vfu28imH
okjCn7481xNi9fHrqqDRf5Z4IgF17JfD3kDWb5Ixy/QBuL1lRZwaWccFMdLElPJg
n7Y7xnWMERXcFcQzNX8OV0XFDZTjerE3RLiiCacDqJ0m7TkIEuEQRcvv8q+CVAgE
dZCQHSTXuVkxt/oQm8CT2UGdKd15OgCtvxAVzl6r49wXwTNKQ4ISvoKMXMm53XeG
tR/fDbqu+A/e7OcdCIRdEpRVr/T2uioYUh7+zque3QB1m6O6BQjA+Pd9cURUxUBm
zFIMlwxDDWkHxhTeFr9UAHm6YdEIC8MnX/bB92fdLrJXbUMmc8g3jF5+IK5KFf33
VsDUlBI0pBJQlUfAvyl5alHaFSOhTJdmZFQMzm1HzdHus5HJ/jD+qfeT+Hjp+EBs
2K2aSNMvRqXUUsySWhmVvFPFafyuG6WP0SOdPhuMZVIpXWy6XE8nrSa49rlAAVVF
JkWod1rVuisOIy25NeSD0NUANGGz/lAKymLXt1NBfAl2wAOsldb2n/b79Jw5i0Gw
4opuBR3sSYvMrGvY6tPL83hS6Qd12PNEu369dZCLzSvr7tLqT/BdLHAZeI3P6H7N
gxCOPunfivRwli5ecrUFRprPHc3K6oZUSFi0Zzx4F40yAodJ/ju6IXO4PdfvuFKb
FkoD+T2GbSIDmvR13q5QO66MFeMiMWS56yn4yk4giZOz+bN2zLwn9Cm8Yue75y2U
SEEJgHqhmHImiBtFhN46V1QkUiKn3DZn2gt/OCswM6+ab61fAloFdzXu1Enx6Fws
Li1HZSW2BMttQ6XfQDDb9VJ9rfIirI9cddGKi7MUyH0i2L1FHWtZwwQJKRdj5PI/
pkYb04ucBkZSZcSOrA6QVBD8vo+gxg+MPjDbKlkKt567mxnaMdzsSrrM8OgDoQpf
JmLpgvdOynCuV3pDl0PvpLu0T0tvfiPGRglzEux4IWBYlA7w52ortCIDC0nwzPfV
7DAWgfViDAm7pbSjahBQCMsS99do/zViEhiJgke28sqnHH0bloRC6BfWysXUTrmQ
DehyLReayaiBlh5Uz3FoqrUvO5dmJkN08aL/mXiz8ccxki4AD34T7aNE22DtbtA0
4HBzhHvmLiJ6BUgdVkeLNZP9in3Cunjp21gCouaNsuc6ZkXne6H30NfbZDD85Hje
ZD+EMOPKSCReYxwWznZonrUEU8cLlx6157cK9QkfzWVWb64ba6xlOi8VGRgO8d+N
5wJ+UGEFgew1ZwbCUXCCZD2RBbdKhUPfZ5HFq1fBewTqLNwMfdZxguGuDJkvTdKl
7xa/FvpPPvIhFsHdgotCLDnL9nS1IUtQiUN8f2lYg9VOg9GOjELzyWz8SfWNyMK5
kdV5nIARZ69PCJrg7/fKbHpCJGEu7Ew3Nqwv+/HpQ4h3CJbdQKOf8iVuoDAjPUJI
XE6kkMmKs3sNdr9nMGDZgaLgx93ZKTVSBGNhP8/qZNkwkaWqaVWMan/tdv1+i6RK
CeOE5cnUdpeZHMpZY/Eq0wzauQh8sZ/ETX/vrlp23n5mj8uMDhY179rZL0HGqFXZ
BZsMjZvnDKMuyrMqOebMb3m6OwoiHYmaqaKyBbwAayIutNdVWA1d/M2xaCqfiyWo
7TeIbdfDgthe90v+UyoZE9OXbGpxXhWMH6P89PmGFGEQ1v6nLQ16y5t+ss3O+Zp5
ROjm18pbJaSg8KE5v+bSFEvigzOwL/IboYYQCdbFx/+e+tXNx0fu51ziRGRWHEpH
tB3VFlEOaXNnjgVCxZ8g0C7GYk8BLdI2ZoZ94KYQvXikbiOrd6IynHzPSj60tXbW
L3bSaTgQoTT0NVLF2gDVy+ygcZhZKyj9MWRXpmqDipBui3gnAx948AErJiz8uyxY
XzBya0INzrTwu5nCbTyX7cJQde+cTeTXHoTF2hRdDpYWboSFF/ztV2cvAx600XeL
7SRxbGdwC4IQzV/N+WrkiQ2/5XofBhgkxzxCLd7DgvQ8sHn/GI40r+GdvhsgBmUK
7+Qb9HXc8Cl/KMyXW8sb7Ngqpud7B7NUBDHlwIMmFt9mVyCfvRCKcG5X+PTIuSZE
v3FF5qJHT+kK8fxuU2e3XnW6t5j/mf/VA0CRuYoRx7RZwOuKHM3Bw8jEgbb7DeTw
GUN+qjOk8MDS3PyPEKPYVuYGx5VaaUlYZEYDaveyzn7OweQJrlY4gKyUEmXef98x
eE4CgCGd0yHzhf3uaZ2q5Efanz64RErcZJQrk27xqfqPDXOSBv6ePnL/H/CxYN9E
OuvN0SN1N9eg/kpGlYmPo9b7gsRHB3K+EYT1J4x506VmfEpDC51/v7E98ajjCAgY
fbFkLvDUDnxBGP0B5jN+/eQ2o4JsYSzPBvrEGqNagZLzZ7QXxs1YaVgRK9iz1NcL
L5e3INA2jOJZug5EHCWl1Il1xQ1DYWM6nUwmdZjLLEDQ6qjxC9rOH7+J1s4Krnj2
yFYNwJCIycmsdaLIRZwKpcarGkS3BTSVvnL8QTOU/H4yYrZ0W6XVfdjdwBagJ778
vH/ZeVv6qIGPdDAc/YRu3Dn78CnR1hjBxWvh8i2Hb6ESNaGxMTvMiIHKeKDBz47X
SI1XnVUTiAhR/EN/TZbCkMbjw6iL+EFCRiNrxi4TGuabIBtGsDHlXjDYsjUCqnC3
7Xd8LtGyAmxkiQMhXofkr3oEuzoqaYcDAIAUSjb7BeNbthyO8GPtTB9BAeYFkmLV
11tj1/KjDufOiWk7I+4zmqkfcHNb8VBAof6G5sa5AyTG4CFM9Xl38fvzVUxxWhtc
vXFLyw5AueCWK9IRvbmGDv3D8ljyvCYQ1azlbdrG/syH7PQCaSIbDZZfxrER6CWW
iRBLlTyzXHo8AVaTrW3JX1FS8vtWCaM39uprD12ShGykmG8JvQI5ZlMUgbwDx7jp
MsztroUhIM0om6XKIPp/Ts2OzDXMWj8UpW1TkF8rue9vva2ihE0o+0DGOkwfrFBo
Kdg2w67hTBebEywH8S0wgmCW1fxGeC0YQgrtr1JNeScAKdl5dsyTo60Z5+Z66g+Z
y19e5i3kgW7LH3eVc5xSaX+b0Wwi+/ctQGnDz1NcpMqxX1Fvu0B+xUR9TI7svVsc
fleNA5dUImGAwj2o2E7hvyugehY1FfY74dLIoyPGeQjO/oZdy9vENmVO5ns10XYo
lPayD0O2c92RSpktStci/xkw8NsODJ6WPIu+WYsRvow0GXRcgGKZ4MT2apD+g2NX
83Z0yS35Xu8MxV7FWu/FPm1lEsqZ31AkywNLvoy0ezwKYrA9y0+EdBKdPAQ9hz7H
9tQPVCDlqmU5FhcgBFcRsZsPFrr2Pyu1us3bJyDjA9fxgRQ8BvDXHzk4y1UpQMZb
UbO6db1y59F9f8GIOo2yOejYITf0EBppVhPcAM/yKqg4xPTNh3GMQAAGhP59R6OD
vNpx8BL9ZtFr6P+L3bzykNGmDYIVCwVmXPFvi0fpalvqz/Qvm+qCIcUDEKJWa4eK
ESb+XC1Lzx2JTavWcsyfftmvDt+vW3ABID2vqnoBMbOqcXKtcMLaQSm9bHPL3Ve4
no0y2/wB9WXymYcM/T5tQj/BZLZc5FPtQ4MW1dYx8MBUDetJSZLuT9gIbYlBe+I8
W/QPIXhAJQLR9aJVXXOE+8W41m/0FL3ZBxi9m1Mff3xsHJgqARPD19Rp+U3l+05w
9tyuHqS8GsyItpq3IcfVkoQ776ejic8wvnJD4RaSXyDGHyBmJHDs3vX4P4OhJw4u
fAkKYuwQFHtkZ0l4i16/o04hXH9+GsKt/DQTDmuhKZMRK8Ebv6smkvieA49bTnv6
92dCuNUj98AdfdxzgKzDsLel5xSLbGGq70i8a8IghtlK0TRf4nJ7c5C5o5JlhtNp
Qf3VAl/0hhvGUuANohyfwUYESDd43XYxXzRZguaNKXlU393JduIQ12JpphBcxSTc
n+vDyTcFKBuf45w8QEJvOVkRQ9KlCKtLdiO5pNNCT0XrMetevOvy3fuyCMyPTP/8
fq9vzHHSUE3lLYwNP2eg/bT5jvKUr4VZ9Wfuo7tIK54ZCW7ZDkPzbSt4g+lpJhcD
nqJ8n0jwATyctLb5X57Wf2wZGa3mpCW6nUSRkXDUjobgK5Chq8S6lIBU3yvyLCeY
9YXIszF4UZpMnFp8D0VcL39XicFBgyXpX7wJsuDSepB6+K91FCvpIHyPSCMsZycK
9S7//+HAQoH+LoeT5Yqb7f1e8aURBjxXrJxqvWl5ktvYrvhIgIxpKd0QXkN1HKxa
aeVm0XztT4Sxrt51IWN3F7W5V9uYIeO+bYcHPzjXDg24axVFulthvAacZpcaGrCn
3MFPvdI3Eyvp1kYbLNGf586UEUXgZxE5ZRs9DuNCQoBVtXkPANB+MCFQQu9cbXbW
DroeJyd/aZiO7qVeGu1uSUy7ep/JZdDToXhq0OrTTrMDNkBbCze4PLkdHDklR1G3
jy1d25zeXwRmKb+rOx4p0DuEyP3HMqf1qrMDDw3l95uFTRc1nCk68yU3Czek3B0m
TfKozRkpgMwIUlydwIHvuEoUII1fpzwuuXyYS1S/wU5nZYj/qcsgKXPjfG5BtITW
2AS8mA8coEeGEhZ6ceIQWpoF9fpMjrozo8oDIjTG6TKlU0ikJyuKBgMR3xI8TQmf
1QgFV0cX602QdWDu+f4uZptgDEoplaj04tEbVMpWQMsy+RJi0lU592dfuNQCu7AV
DCiQmVCp6BS47mrZvAJdyDcAQ/mlIfOR+KLK1ESY2KOfV4jLey/KJ3nq4TCyK+vp
vfBO8SNxpdz4yilG3vb+lKT6ugrMb6khbfyaWtcunRSIXiu7OohjidF5ou4B0apL
BeTkDT5LYWjVD/7rLNTVL4cgxJrpfJeXpe8hjkEBnvFGqv5g2/8qQN1yigaP5fhr
+WixvNpaOOqfi5ZHBRcNTu0XaJ7SyYGG56IBbQ7YYjoIKmi9Vwd8MyuSNEJhIjOx
92+rqXuFksG+UJ09+xLKyiQuep6SN5NQYDkXg6Ak+0TgDitCXsLOwT88HI6UkVTb
YsDy8dI0TOLaVBFCX3+z8+dipfvVvgOM0Vu7gnR+AvUXizaN9B+tBEeSD3GSnV3+
glNGWq5W/XNiIz2L1CYSuDfglNbaOSLoyK2p1RyqPOJNdwK1IAc+1bTCcw02mD4k
50Adl9OLGSktBq6gAdUaubsFX6F+T1RnaiFwnqKV5iRU5aUHgaNJ01kTHJ0LBc0F
VMD144c+td8S2C5UnQbdo7CJi/Pim07HRfRR0pOri+psOSCEl24o1Zh6RAuL2vHg
0b4L+6imE87UY//Djv6ImghnSGrKnQEbQHEBq/qu+s4GwFyXWKgX5uU2r/MfJkFo
5tM1ict46dX/y+0BfWTYzrOB5nHYAPkaauizk7jEO/YLYn4GEeaCUYXPo+qjKk9w
33K+xqKF6BzXywroTrxO7JNPQnwB4CadoBldc6lhh6zHr/UnIEzNza9zX0AVd1G1
hujarOwx4EbsR3M3J9O5cjlvvPzl//p/Q7ZfPie+yBWKC2ph1ypWjOrbcfKZ30oq
2OnaSYdQi8auszv05b1sc/4h5OERgvOQFiwtEL27fSpyOJax196h6vrFqcsST7xV
zVZmP9gAjurv/5omQkTXAQQzppk7qjUar0IaqlMq/AwZHAUZ5m3TA3Zn5uGtkhLd
g1Trq1SA3/eQxTZTtrRgT7o8otfZPMthxRIKg96i44Azze77cXdQ4ZiYdFVa3Mhh
QrhzzkkoAISnw1h/3n0UBNQbcH5LOKifu7jTiXQ0HtbvlloR+Zqddn/aQnzmyOaQ
knGyMTcvfGDVZCHpZAiw6WFXT/zIKqg6iKpTi9VxO7AfTiQOjxC5/kOpBfeFEi2f
6B7LHxxK60ssgN0Aj0PKN29zH8sq7jZuGJfbdY/ihBWaXLZmArvchm4DuU/0Uq2s
ipOVPhREFLgz3FZDpRf6TYTYLRmgvQo50f58BYGL3vg+ZxOgS5pHF+MjlwEqAntL
cf/A77wPJDVt5OVrcUHr2wjCibPn8QESVQSMM6X2a0yTPRmK1Pe5Hr0QwZWEnGvW
4u2obq6wAUBwvfr/JgFlINXMZ/XBFz8YpSiW/E6qF5jTlBRPMO6R6XGAjI9qi8FJ
/AmTKK2oJVmPhLocZLj5cKiqcsL6MtmtQdK9VF2xV7E5CPQljPWil+Ghs+i2Tb5q
PaefhprcIKzDzzodvWwrLjWZf+U54JtLcj8RGXZHPmrTTRsDK6mNymRWhT28m3nr
aNSxSyfw/mLbdgvE73pzK9H2GiZSOO9uXSoxJAbbJYWCXBgIdK8ajv4VNKXYHQot
UWwQMHG+UNyQMPXEba6r7AkB5rwH5/rUzwZJRZgAu/AfrI+lxEQutwthTfNlS4oP
Bd6Avz2pTtuQzfC4dpxh2qnPIJZLsbriD2aBCDKGlojr+YB8/ho6ALbNcuG5SKfq
Cb+F2rpUaz6aEvli3Rq4Kn4avX8tAkBD9tsn02igx4lCY1J3nxpTOWtiIjLNkUcw
Wom1YBH6ZkKE5PaEGMDxlTYpZEMzXkX25UpxJMRXODLvpI7QWJ3fDWfhm8OyZC7+
LsLQKEjbwFQT9DnhgzdCnFRAKK/jyBQztd4lls/DBYAq68I7s3Wqk2peJ5xbTnIH
EXl7EnVw6jttt6f0/lviPU+s90UDushzPnYh5eyfWHbQuNTWQrFPozdxOYPuEY77
6BUfQfvbHeCVIBGdc6W2i0MvvVNmBjvR9icf+lJjOY/1aDOr47n9G2Q9ChJNrTh4
7XEESU6aypfB9SWhNqDIfn+fmos2KycvIPa3qJSvsjzhdA92mCF05osfvBM3Tej6
A/Y/l2dsoodSfVXZA5NMj7rsu1um4W/y7JmlA5GQk0RC8CuWFl8nDwHrtwzFKOmP
O5kn+aRcvz5kygAj2QJXfBAOsEHqQk3ZA1RmAWYLe8t7irpOJ/1S/cB1IbR8cuf8
j0gBsTAR3UcIZW2riswatArZqgYOYezD2JcSdOW7Y+WjFyIXwUT76jb8LqNBwnnO
HH3pvKyGeucN4p4gayUxplghqtPT2jQvp/wyKPHjryl7bJOGnwBm8JbI8Q9LnzNm
q8HB/ItS0x/loslxga/jLLTUbo9C7tA85rY/09Xi0lb8/oS+MPxhFGGSjQAUlr10
E0ISzahuXAnGUCXBJ5uTsW+y+eRfSKQ6rknm7ke2to8EMqPHnBkI+ZZVEIyGJwYf
Kn8oCVtbystuNe20meVWV8SHX4etYszk3IdOheuPDyEaR6i17fW5Duqe4Cu7MXii
x6t1ATdf4xVrovJ6OnsFAN5JR8ln15cS4jP9gccT+q7bJboAU5KoPe1C3dF6OYha
nRuirh6l5BaekOPL7fk4dPMUjTtdtjOXkMMAsvu0+FQx/i70vNTx/3n5JbVWnXgm
A8Rix45/trQn+OJjJtkyUkxf5Gpl2YGzKpIiWfmr61KJie7WzHmrEW5QlwygKg50
1WFquo6SQfFVR/cNhaN7Z+o1TkGFtwPT3Sgfe9dXF8DmonKgoqpBE5tX9Xy/c2CD
GIb0UVAmZaY/us1MlVG6/hCfrwVKniUqxYK8Sm9jTQilFVsY8SC/nwMgilQWa8xS
Yy9jmAt6gX5CKG83CfPxCGVun8vxwIXwZWzit6C3a2IQSNMzkMGoki3Ia/vqRQe9
FssZV/a3MKkP7y6TlPZBnS/asvNK/a8dL7/U1jZrrH8aqguJXupA2B068oDTGYHX
z5jMO6n8qWdAe0LYHYw+xG0WAoySCSDo+JnM6wyDiMNXbGh9Cmfl+OswQVmeNLtZ
TeGqFoX39RhJxbr6R9QaoFe+6MWU+DdAVzO3cRsgHxqTneAa1Zly8jL09GX1h54B
R3iltXd0NFJDa0RR1Ia99v8maVjTdqpVyOAFVBAGslkhlOpwPVWYJa/5QwGCPI3p
BjmeyJc1Nlpa9dSD9rtlk70hv9K/mKXNHhQb7kP+c5PINAo6+I7a5iKulFjhgrm1
KSDoQu6O2x2iBu9J2t3ZuiFhx/XuZtoE2rVe2MctFtodYzmddiGTtB2PH9Szw3zc
mDNSkPkYM5/Stcfx4Rb9XgqOgDBpPjbjGxEdfZye/qn7zvmFWdHBm8F410OHO8/h
sjyHPit3wMDF9P/YQMrDqdCTXzhgwE7VtSQL2cOaF5nG0Fz9U2HYNj15pxbfA8Oq
c+/SAXx/m8mC8WPczDOhhJzHuGtyhfS8AehWqoIKCzHkEylBeliDVFR2zAG3eb/y
OE2mTNE4QV/fsiD64TqYfvQsLLGLBhbQtD2X3285uji1xY38szRqIY10pGPKUckH
`protect END_PROTECTED
