`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbE/kwYabqFxlMYiBeMKHPgo+YzQrMgMRNCuQkFyrXSbffscR1SlzdbOKtj/LiDq
lC+XbO9Fe/SIavlCenuej9nx7edrgFRa3LsXvtldp+1PqviPOEaNxmIGfPupt6hr
qW1xFpViRvwntp3NBmWX99xhHG5g+RosHiiq/MKxFsOBvACNwqZSOjyIbbTRn8sZ
bndLzQLugLYggQ81HgzFW6tdq1OUUA1Pi00cpB5AG9j83QJ/N+gbtfjtm5P0rwLn
2hUiImVCDFowywPKh9QmXQdnbd53dn3d678Uqgx//aJfbZJDc7KvVTDMVJHDeivF
ZI4ZqvOEVfzh9rHbge/0VKP9//CWvXa/uncirvWDYIfX191/jkPzM0YMH7sz98nX
mPUTzpOShsFZ+JAAENVqqpYJ92s8mDgDsJIGZV7HFM6hazztSn67BO2Yc6ib1tPb
Jz9osquCdMwx6DtKRUhmuh4z7NwQqvG/hSOdhWwoxAYK+JaVcEqB+nfg02cPBZb5
c+Ns8RXsYvk5CjouM0ltoS4hliBsti2+PlodKSJHbXYUqcGcFEGUsDv/cF6VFof8
KPosQGaFnaPQkR5J/glMwCKmPs0DE4L8jZbqcvMXOHWnqpGWbjFNxBX3q6qwvQPW
LiC648d91M7zbVFkJB/48UbWAc2eczWd2eSajl+R7Tw/M062Z/WOqrhPkuU3MKtU
1exK9gISobyiSUtg1ucA6JaRtkhfvBqsYr4N8jd+tL3k8zliLMsxRXDCiPVsbxFe
2lA37QOIiy4zpmpqJZBwjeS8C7THnLUkLEmvrVxCg8saX7w1VtFfj0qGgZuGT/Am
GVuRXh6/r2rbbtkAnwzq4E7F3JWEoKzS3q2Kgn7QnT1o2WkCaaccVoFvrUEsv8u3
+e3oIZMINl4arSLmL88ccz7FVGiwDfPlUL4mJu/OmvLKc5gJaXFgKYXkBeIc9LeH
JNQtBfWgPo8y97BtwMHJqXwQ4T9P+ADg6p3fP4OvcYCYz2hh8vz62uGHYMxdqjWc
t61f2GChBzcmPS7kYVnPWbShY3rg3d+K63eFnlt3nxBvdEY16eoupeG8ua81/zZC
hLPfDSYRMrA1T1E/o8D9csSEOKmHUmNBYIaNBuhstD0=
`protect END_PROTECTED
