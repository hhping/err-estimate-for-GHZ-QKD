`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dIgojRrTs115qKmfOjnNkz8WKDB4RD1oR3HbxY2ssL/XDlOGsL8Qi5NTraSGmN8
HxDoBCkbUaujpTpiERYX2cW99akYbMeub4Q7tuWLrfVSqLcGzWU5A/J1Ty/XUbLx
tDX6HmTEdFS8J/LC8AAaXN6lqs++6jUNlqug7noydAWccc+hG+XL20CiGXELxb2L
9gFbcFHYXyWQLIvMqPr3qe1L6kMonGZIfd2FbAKwPQzjbykUyTIlPZxaTq0tmO3y
fbhcHp5z2pAXLJoxPBG3NaRm35/+5v0nJGcj4VshKnm6iWR4qZ0HNccfKxZLyHDt
LN5QdOuz7Q0JqAdNPQcRyys+Uv3wgzQfmxecsc0+CluLQxE4GgEHZbkgEPDCGZjC
+gD8/bHtra5J9aP/f4l93TSShf11DnGZJuoRbh6vksSCnSLvxV3kPTnhKzgUOeFb
uRp8PAyXsebQJrtD8jBt2+U4RE7eH6QJJBZ6e8QaDI/Rtkt3VeF8T5mUl+Jr6w9E
mxqyKDTRd18EyNd0NcYqUmh/co0tZxH0m1jeUvl+9ezvpLKcGoVtW6yKmiJxZAxG
hgl5P6kvnFI6BYjLCMaoZVY/BVcTdATlSOItpqcgNqiRPrCKAphrUPUnh8AK6lZS
qoTHNoNe7Ez3H6xBAJ09cgaUzXbgEQmbSmnVv0LxRJRFJmxrt3CjNyeaC8Fq9JgY
QsKsfBDlZCikXn+w9NEpT6wbIdcgouE7xFgQy+QYWDV/wbmsAietz7UhiWkALo5s
9n5eEnRKR5xByVnCl0cLG0X1ZMGpmh9y9hCIS6B2GuijgusLzaaebqUfe4zoS5Cy
1mrEzLMKauxiTguD1Hu+4N0HRs/uFTuZ+osIdSw4ywp0GgZ4N2dkKvPpp+1AQhIn
hz1GLQPdC9+DjEf9GPukRg6leKn99sJuJcqm95lo51Mjdn9/V0K+spzTTftfof2p
1um/uUjC1oMv9N5TuxntITdM/7Bx3EiKZosXi9EBiWXJRJOtVDguOgaTvP4RZZfW
d9smPuhsbSBfyH7X2ro0LcRug9IsTKK6AXBryp2lFvNAYEdFkkfp+jm5CWVKzAH0
TGzFW6oXFyxgXFZZP0YrwAbOiS6qops4TRaYYcF1fYyIzZJcmeZ8TTGKUnDsGiLO
I5FV5ZS+BdoZ93UXysWhlKt8HGT/ESxVTwxdGAARtaeIYKqLJfqlL9ML/6AotL70
SYdbqNfvJyYOBg6AVNjYwZlqvVIQ6JJLxJtLT78bu9hdS3LFt3/VtNDyRN7wZieL
8ltxsy7b45gsLPtqDqC+s/tlF9CoFiS7i4W90ztkF1I/WxCNyrePHS/K9Sc9KlDq
fIajvKaWOrI9xkMAQfpF8h8E8PkGecozGz+9A7HKwNNSO+o1Hprtu+/7IKhHJfnd
KZaeReIzd6XXpk1dV8mSay/qRgoFS+xpfXD9ziqGrtz2F0R32Zp+2zH69djCvKPN
LK+iRpe3kMhNrVU2rJD3B+I8CJQVAYKc1SkHZSDh310=
`protect END_PROTECTED
