`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRdvZi6wLOpkVx0g2oBSE5Q8j0oQJOMqkOxa0WW98kio8jB/hcNAxx07Dh3rn7be
fH7qXVIRHXXKcJ6mNE5W8oXnU99VfyCmNz8nF+BEhoq23y12TfqRJ9aWXHCI36qX
QMKqF6SmDt1E1/E9Q6cJD5ItI7jlu4+DZvJU9+VWGe0UI99Bvi9stj0GjpQ7wEmS
ZvHZkkpehFz1eX7LAX9aWqmEtd4yBIl5OB9JjupXwCMgSUvK0H305Aih0vWI42zG
q/3ZDZ5Rt840vNTdks/dRsPxetxrnGJ2Q+Yu1SD8p+Dfit3CSnXuSYVnah8qR+R+
c2BBTyyhya4uxOLLgYnJRxlQNoXnpTES2Qm8JUks7jR8WblY3RTFbXhbgvtBvZzc
RYqyxhD1Xo9CpFbZYNW9PikKDGF0Qwxym6lxAkymvWhJA11pPDCWhBDUnhWOv10W
XD6E3q6jcWKHayLW6sHnX087RVFvqWrwO21Efl5kZXvdIaeucLQ/mJjbHm8V7oam
sUF/hx/jXiv5XwfNuQG5g6WGC21JPCPhyDRAXoMcCuMo956PuCdb4i5DGigmVvcY
XSfPPxA76/I/iLaIIWlNY7eDGJDfEuZmalSdqczaIQ38zetD62+UeZRF8htum0zS
XUYVw3VDtICKm/BRqmhZcQ==
`protect END_PROTECTED
