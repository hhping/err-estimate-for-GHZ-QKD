`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFWbwCf/umz9Jt4N4GlzKVsbkdjNCWb+wr6xOmGJWWS9QxNvRhJA3ZNBqUIoTe5/
hIiGjbqA9nbI8Kg/GK1s/j2JRNHSdQI9y0qtQIpOLSBLE7s7W2DDaTo4SP4XdIsW
171t2R6tl0roRgJR5wT+2kkul1BCNOTk8pfJU29Mc6oG/863sKt/6hZNGO/DD5wd
2c254bnYNWR0hiRo6xOCh15EHKL+me9zqWQjtABM+TMAgxxzqMpIGCNWO/EhYuPt
nKRbgJJyJfo1RTu0SpPj6bwamWh686knZKb+/K03PZdvqzRiCPYhYObHyiPhAYlq
bZNr5Y94fwgInuV6bpTmJNdNueRTth7W0Vs2wZpoQLBhDQFvuk746H+P+L4gxZ35
c1yjKo6YVBrjpZw34HtBCRW6K8MaSV+mDEAnlX6le4RcrJ+jdLsmSMdkAY92XUVr
ccsnt+ZJFTusuPtMnXJwku0nnoZDDP0vmZqm6+zmy2gLpZY5u8h8UAOPUsgZ5au4
1BemXdV+azuhJEOXCOxRq8Abxl9pMmKkOpaoYyeSJ/nCSBoa6XEt27dYDNwva363
UrNGvoe9jD+bTxIQNHYWQp6SR1h+VzNagdnYFgdZXD3CvGD/xNWiK47RFATbsWH3
llKlioFZ3lRfzEWf9BB3zsRWZnIYAwKq9eEILZPHphPM1DJKoGrZAnUBOrwN9mDu
RexlXwmxZ+Y1J1I6WHbppmmDXVvoZRIWWYUabnoF7LOsV/vlu/HR/kJ9fhAh21HE
koEwiF2hIq2bmrfFjeLR9L+2u8g1ZzsQ61HnDSL247wT+oQ62DQZpkrGRYxUH3HW
ncp7owqO9clHPaO7jVMdaBmZx+Hx6oaGJQI6xiKycE4KC62DehJ+O6wACVnGFSdE
mfe1NOHG+E/ym5G4e68gQW5HW+gsRH+UU7JHJ+Vuxuivb6Tz8g/gwmSY1OEQNZZb
vvzU7ZSXa/78dWJMF1w8RfGWTfS3yqaAgP6IQ2c0E2SbAadk+SKqMl0cEV4JYksv
eA9gK7crbG8qLgW9cYlIKmJM5oNNaX9BNkmK/UcUXCy3pe/WsZ3uXwb9di4CSAa0
ulh9W1ZVS487wELr+cFY0Tw4+nCGrYFmXk6SB030QCRlOSojNLnby93Gk1jmF9Dr
2W/rnbzRo0sOhIxfj+cp4T72ZevBX7ZYXCxJP/2sogPL5wpL2J9Sh+UyC1onn6f1
dWVS+9nUoQ58QdAS7HOjnFvVG26Ui5wh8yEoCFd6Vx3BdYZLVuTkFUqxvYK0sG1S
8yLDHY7ieRzQZ+7rA3uw5g/xKiD+o4GEh5icZuZwMd34LZJwOBqcFeYQyB0UtRch
BjiIj5em8cWKSOHu024bs1jc1JCvQ2IhaIO9LKLFlZyr+I8C6vPJ5ncCs3crAnoz
1Fdk2JJluM4ThcZrydxymh1oXKqpKwl4gctfGPFukHS/g2u8WR/y5GkTbsXxpIrj
G3v0op7k0LiY85ewenkyIUcsE3S0wZM0BYgfV4NT+tCBo94kDumUFGd6mXTXBVTD
yRMePVg3LkMVHXI8O59/WmsSFGfDkRLvlbgS6OEvFZSHKaJiFLQoh6P1ymBCL7eh
BtjELsj0QyFs+daEX1mH5wcKrq3SAu5pVpq19UFU1xYgK+OVGnteCHjjnyyg1Yjk
AcOQy15MYhX1X/bUW0YEsc6IbmsuWeOvGId27YXCVJN+y4QkoW7pBegPFCxlGzWD
sNiOR5qGSPEZAIXYV3WKPphTaPwMLEm92a+AG07tfFovjWMU39TyAkZtByymGn6W
2LqRBlp79/c6cvYlo88w69QDC5JXDPAgvR2eD40m2AaJD1IYy10NwZ04id9TD5sg
VQMUASw4wYrHSRcDL7TlRnuH3Uh84PM04NOB3OWvIh7+r1JLNOlQXib29Yij5BAA
Q9qaVXCX7c47hs/LQ4Qgrh9QeBrLDXoxOJAK65fjTIcBqw3O5JHwUj9mJuy5lT31
ScG3J3kMIthKxZUajBK9swRjZvPUEuREMRDkOVjKRe+XGPgOVVBzU5pfFMdEFSN7
7Zfr3wgEMGlBFZqEDkTt6Twa91QExM7NiOwnobH/CZo=
`protect END_PROTECTED
