`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGTKv/GGLoTL6omx15KBWDtLkAWIC+uap3LGSJpj2BaY4V5D+01lSf3jfrbTr5XT
uqNeesqblEFaoWZvu/7IoUG/sb5vLR1oyP4j4VIyLuPT9nBzSw1XDVY/1RFej2a4
qby/ykIy+92WcEhlKyZ2XYvFdlJTeTP5V3X3wbhio+QKmaed8yKjKyWnyK9Rax6O
kL7FtKGWXLlz/xt/4heXFDKlArz4Do2yap0BGUre5ew1cez0o49TWrJrXd/4Wn5M
I1pg2DaEM6b7Fmg6PaQIeWvG3qt4W2CTKhJFiYqnDCfTG2udRE6jkUZhqPv6OJfu
zZdeUQE0q1+3aPsTaZR2/6FADfyqgfbcI8qmbCUxx/JI1tOCcZAx0AGInD02cdS3
ved8R8ph9ZEYBy8UwX37GuBKLCJQd0yoyXYixFcjvMeJfZeDyNWFmpj93j/fbf9n
C2rVzDinnquQMksP+4AhbfxRp/fe39Vt2gJOPw3Jr0A4t2gWP8lEyP1cotEbK/Qr
bCiJzUp6hzfins69wgekrPFc/LV43u0NSLAIWQAcRwxK4MxgTQjLf65cZ+pj/ey1
Wu9DcxxrzLSk3f2hFQnWUHuDqjXfGZyOt/ofpumrWs7UbaJ9d+j8nIRwrlLYgtkK
vPIhVFbIswPugTzDIb35/6f+wygmJMJl1NYzVNQrDhf5XD4fdcHn993wD+RTY/RH
z1NPTSmtIPJqUv2hfeAQ8tjjmwzW7o+kHVGakxPbkoM3wjzOtYfdRgeK5+9EuAYv
VDmCDri9jOg48u441iA6ySW3z/ef19Y+eIEiBlMNVKrhMTlzAA5DUcCyMa3oRivR
hxKA8Lwlol4wiMGTyiEbaqcAVQhcOODyUV/zmsBnwveDdD5xLaBHziA54rz7uqo6
M7SKgDCrRGWl/aS7nj33H0ealSE0HzvnbQ46AWtunBWX/Pi+VaRR/2VD4F+rtcpi
lpdOVtRoxH5VkeijT8mJOTIq714TIPhQg4sYB8X5hlEk38pYkESmYgUJEZ3/y7qS
Mjc56wB6hGj6v3tX5jDwGsmLbI3QhnS1CKDVrBL/ptuDzd9eWcPMAOhCV6KzVLeu
dnP3YKOfMzNb1fKYcoPw5DoBnDlCpDkDIMhYPYMzlNVG3CvnyFuHYsWkj8oIabiw
96XkSQdsmQZ9eE4kRZZKGzsOcDYr/OW5zgbQYvFbQuv6hKBu2QaCfEN/2twKLzy5
MqF7Xl2sIjVAeB6PvPYOxwQtldq6IAEuK7x8P0L7XjE1vH81kcvjhZUmar8b4f9H
NSQKb7Xull4M1e9RA6FSLQiXJPGSOWaLQLIJ1JdLkQCCRqutKC1oefWfvOeR/f4v
kNsURL2vvlWbEnoTTb8Xsm6MVEAnmWdaCgCh2hPuGQifl3XI0KAjY7Dt9xZNMBeO
y4K859VMgnoBX7pwA3V/b1QB0831tQRyC4e8W5DFVMQBWqaCQuYzb/GCkfouFmWh
Ex+DDXCCKxbosGj1nMnTHtzZAgLHMjJDkimgNyC8JRg3OfaZmJmzNtGTzaGunMop
lpZc8Bvnm/aJxK2CSEWMxQcJsYF/Bk8Fnlpe9uxejbtg6+GjA9WIOLkwkb5ApqgB
BvykSgKTuYpBgNQl5u80XM6XtWVAeQYTwyiV68WsKeZ41xaQAuHO1jW2MHZ4bFka
XQU2g0g8K3+KYVzJlxZWrsxUdxc+UYc60oHGMkZUZAuHUwFJaTpGe3oGUsE/VWNH
yLExQVWrNXt8GZD7T2KWFwMEZgym1PXL2kb5Yj1VNRkCGYnsV6uw6mx6+Nop48PY
Ae9mO4/RjyJ88LejvaPThVJinVTaEM5i3II9efZWB9zeyWJG3eu9GASUz5dybnwG
78pi3Rj6sFOuJW0/eltCw6Ewt7YgudEuw91D9bKo9E3Ruc+hbdabiSwIO2e78Cxc
bQgGNqosVHxl9R+YKzYcBXmdCzwn/GuI6oB0TOwnW74bDS+bHzJCAw3tBFm9Ba2r
SrERtW8CniMcYhv2PxBvqlOGTYRS3DFBHeVYS1+RFooGlPu7B4NMkhktnpicCGZj
wvuVn1IoWxCrlSr/j6ab9ZuRQDifCSrqpDrvjlVLBUdlsDOWI1l+NbqcyWz9HtcU
DErI9W2v8vtOoQ0X7Nk3krXB203WPa86a2Wi5wVKsPn/1YBUFqUS+MK4vLVkFifL
p798LMQ8miowxHLX+b/cJXtQbtXREhVRyE/uBo30k8FlPO4osqzofjYsQGFhLbeH
zDLYT//Gup82cIpfnBfGU1Xd3jbVH/9NuktD6LAlHWtx9f9hwt1gCizn0Rr4RMSE
VAKcSkTnO9hXM/O/62cTdHAuC2DqdkhnulFvsd1Mv38ufs1NKuDulmXZb5a1bijP
2p2kfLjosT/lQXOQmpa8BE34uvUSWl7VqWdMk+pU93CJnZ55O5oiCCDSiABOcqvJ
n6nbkm5ByHEg+C7eePDBkEGzbptt0rkAimbkNLtvuPExO2G2Q2BRtsH1v4iL1Fnc
n5mhnuFapwlt2Z9PA0KDbewxzUZ7YqeDs5y54+94OPibWO3oWJuUzEliOl3HQuoy
`protect END_PROTECTED
