`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mr0X9M+fKnAii2wNzf6Ijn4+w7j7GMaCP1+b8eZ1wsCzcglVksvsqca4zwSfIHK/
V0pTkLGkzWZ2cGTMl4r/OYALzs2WbRg3FLkV5FfDhO+H3q/m2l6ds6eEiD7xbYKW
6P3X1hpe2Qn5owjBw1lb8al3iPc8ZurYrocDRJ/07+3o8fso3cRU/fVQEPGEMPEj
4ziGzA3MO/6600nzPYwkBROtnkvjyae1XhPEw8rsgg4=
`protect END_PROTECTED
