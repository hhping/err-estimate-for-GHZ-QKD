`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2W+jCncGBFv/hEWSv/EPyEA6acdiPe6fmJOImQzDJ7dMVRZN/iNyLNpRz0dypNO8
cvcP62e6P4xfimLb26mhiINIHWLzb9w0oe+T6fqKotHS6/PlfoCdOUvgdLv/PWLS
c5vZbEgzen5PRS5OYhhDg26i4PfTKkZJrPAi38A6kBl6pb4ZKd9dg8N/WBlrHblE
MiVCkg1aMefRm+ujMVZsaS/JuPaNzG8oALLyDUpE7HAm/QqBxSgclb4NyIa8obtk
9nx+22tvOTJ04m6F690NEst8GgRPEGqZbACeA97wA0k9mtz76IriVEDZq60vWnof
LLCdPJ34w5mxCXjeWg/pfnnKNeEN+xh8h9CpjLMqx2Ot57OW/PEwvamUzcbHfYQe
I1ap6RdG6BINydTgPkc94NyOrUQ9On38/DAU3/QwKZpXK9VdRWok54pcJ2yhCYMa
gVOSowr7tAY8wyLeA1CbfjxvXuUW9l/nJCZJWXHUSX0SxV0E8Xbj+9hv2rYhbJCv
SdeVK9eETH9VzcnDSHWZRdQdBvN3jpBJkOPXXkLoo+3ly8/kgo1Ml3GSp0DdBAA5
re9/j617UN2Mx3u1O/nhWX0q0kiPj6Fb8qA5+yp4ZHdN/02tvb5UlvuMzYxXsDAs
`protect END_PROTECTED
