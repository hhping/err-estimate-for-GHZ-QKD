`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlCKJZOIpKEe71odsZACD3XA7NEsK1q4AlmBMVofcVk0MeYfcCo15qR7kLQBt/Ns
D7TDO4YcgA+ChvM+o4XBdBHYcNHOCiT6rr0SG1bTQWf5nvx5tLnknVFktaKCa0lL
DvOp2yvN9sqWhLQTWD0b9tXu2F/3DqUXMffdnMWXtK9ww3eby7jlzIu5hyD0R4yr
oemZOGh+cPwFeiNPK0lba7/WGkfagQmYx5EnMba7XtiNe26gWvUQEscQ5T7CKZJP
i6e66b2FIpV6MWYHaTMeXLv+GrpyIkElpyZYsX60TNm+AEwzKkbEYdcxADctSv1y
qXe8SnmXjNUeSs3FJETdMHKBL+CK+dT5c845DlmS3q3OB2Pxxbzk2QMGmh+grPNz
yTbcVn5fg01XRKz1DPUrr+pMGyHxQL5eLfi7Tqy5d0FTasdMcOLLeMgnq/+BVej4
V2HfAELg4l0ZYJ7kdefoM5Xh+2BWvXoCN2JUjrSy0ZJByjZzPjHHa//+dHDv88OQ
HqsL96+SAZ9+n1eIvd1K9qH6JzvHkQQ3HZW04l/6UfLaJ7yYMfWsXl9qi7ergX9F
fJpZ5Oon7pWMBgP8y43eU3ZmTX3TBFmpekbbz1Qi1ZrT14xmW9G63UAqVyzWiguS
Bja3KruhfKsQ+hy5GDc9A20yUf24z3BDApa0nDvzTstfCMXFEp5zrrHTu/T41nAF
oNQXTtGahLHW/mOk8NTEEzuvAWuxO/yLbS9gaz2qc993qxf5k4zeIVBOO9ckc1K+
yZ8OTWolejeRtJZXocF7lw==
`protect END_PROTECTED
