`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UwZ2BSL7GWGBV/c7BIeeILt1wceXWv/5aevbf1A0vt7D1t4xWF46J2t3I4G4O2fT
/NpZ2sqQFGiMql5GI66obxFl+aufeatSl2QcjkgvgfTZsvcBQKhV1czmSi5Awxrb
jRwKGZSg8HX8NKjcilquU/a7yFVPGtizmMqAl8obqUGGEN1B1EL/EZnjqEQHduCd
jkyYMDC2Cht53ApXl4PiPYoTUJ7n/Mj2JknkbHhV9B1tlC3bAaY9rxIMjDAG6x43
S7mkFb1Pg23zNqt29HVtuny0NwvY6f6kVER/8WF1ZLiEQbkjf/QJJIL5eVJdONlR
f3JTvcOxz2nsaBLYuXubMp86aAI75bEMXenUvagfeHWEnExc8YtblEkeiAl+0Vlv
9+TNE6XlJ0HVwtuvCBFHb64VsgR7tLPzDiThj8q6iVxs4/Kr/s3lxJBiFXARsYhF
liyjlAYbNmoo/gcsyW3czlsjpFWpaADR6mQuai8qDipMJ19ysyWROLOZkJxO87Wd
pdqFIkt2KZ85J3inoryLJvKVuSZlSj5RkeAnW7N8H/bUjONMevPH3CM3zFUiePfR
p1sOhIKasnWoOlf3L0s1OKYcegathMjHkb7JmeKa2o2r6z1T+VmMm9JH1+834UbT
lXTn84Ky0o7qgd04fAn1h49h/hhuSXXcyoBAanwS+VcqAHmPNNFGMpaGJT1EP23R
TzpuoFXrUkGwIwsqb0w0qOAbFIcHMzVhsMkH2qVAuA3bg8y6Qbt0dSNRknABuAbQ
TEMlT/02STPDQ41GIGy4F9lJnsEY+8gupLYjbUV39416Wxpu6OHmlmFWDCRez6yi
uXYBJCgq1WCGLn5Ntr8FoD1Bx8R1mxj9LjMo0mRWK3W/zqbSY7A4g8LoIM412bpV
hxZK1TZtxOtoDBIYbrSDKXuuiX+dskOq8vz46dbROtFj5MKMU17vmjI1hpyUvuLb
8enylxkDLW5kiBEM3Hdw9/zVvq1PUwHHEyHHUYV3JX3gVKMYxZ96yCPKBJnd7naS
vI4wAp/mps4Td8J3hztYsG2EfBqeN9xYGiBnMM673LFyBW9TQ1Woqw/OxkaytzjU
Nh6IykYtb1CSVo2PdVdS04JqPBKKgotSC360tTxX6a4Re52kdOzOSGHPNqN45g41
ti1ZTyRCczqhxQTuOKTeKMmOEaPZ+KkI/alSqsIrWKOSLBvAHVJn7dE+zkR+g+HN
Awe5shXQpSYbpkbUMoxpBDb3UHTEQ1CNRykJq7RE8IHH/4QS8jrDlZYWoHhXnYeQ
Wvfs+RcGk/syBeZzG83896D7y59OR1pepoC52257LuCzIxDmZriojpif+VZG+7bl
wvinUaZh4U2QeLk7r2v3iBDoYmucuwZo7SiTnH63/hCYFUB5lv808vgR9ca79+cd
Rjfsnu1950xLkXlevDwW+5QkrNSi9ATYvSfoSnOIhFLsU1P7f/u0uwVRKhdLAo9a
FznUgh9mv69fgJU7UYBjhU827ujzdXI5bb5WRDZY4RuwfjqwIfjID7p5sKYv/307
gj3/ktFxFGJ5IedzVvEIi2TOr3GK4xENJL5o1RO596Qt2rS2d+c4+lTqU/YzLuzq
Oeb2xgGlur9sc2M+tbCKyCQkEVQEOUpp27To9QeL68iRDTPW8HhjkPd1b+ANnV4l
nbQj5jyQ3I+rApRUED0+kw6j7G78yztbIoeYCdinP0QjOmDUHcnI9bCmDThSYMdj
z6tc6p1QGsPZqZko4bd3DAfG22m6mDFJoKLBxeCGq6emGQjiYFTEHjlmCtM0VKPA
sa0pjV4AKQWBlRfLUEXlUfktzGD3zz1r3G5NnWSoOABbk2tHZ+xz6PmXOFixMPo6
iKX3xcr85wncWCJlWDRBrowlu2CaIJ+tqxClsz0MQZyT90GzoxXXkI2Ap0RTztGj
IRb5HPLP3+kEJ1guAMJg6HeP8SZBKEmLwbPa1kJ0cOTQ5pQ14Cu/K3Cayo6CJyAV
JzDhUHzvHVMEplQC0j0NrWsI6zYYgOqySvLrs3jm+5sQfbykh1W+I1fuDILY21GL
vWhvB5UNsewY4kq1rL/ZPKs+5vslqsXd1E14Tz1ZhMSomm2Sb1LK73L4EVpET8H3
vhm7Aiq+tQTtmtzbuXDzRlaPrGPFoG+OkfqFdNQUN3d+e5xa/S5Wg/pp/SoxCfYw
MhZpWWhGkW0U3nEpWXWlgy8izV38SoZPPL9pkCad26z9VkI1abblte3ab4cdIhQT
h+8wvwqDtxRlOltiMMXxzbE6P/rxD6x9N59Xi+pW6IE2xOjhsFv8q9Vl0sas1u79
aQVszM7qyDjAMlI+K1TiJuWq1p+k2/l2wcpm8dpTLUpkULiS4AGR1YdnJt37O/eA
5e8N4SuxsQqvEhFtRrM9w/OaqiRSAykqsL21GCAn6k6+9t9ieJ1dftxICvsJDEty
5ApEAWKo0nSnFtrOXhTui+SwB5Iyj9JaXr9JYLDwnlwgF6Ks4fn5t8VV++87JEkZ
7MJZ5oq+7/fCWDP+nPubeyPw8YoKroTO4IahvVFHknHghQL2fG1IU1qrJFfGcCKy
z171VGKYtlEtyWUkxBSA2WzqscRPqymmpd1p9dWQDfd+0Lt+0/9CVerHGy8S3Qr8
uxZxLkz2QEEIU7cFdF4TqKUEvrOu5ZroO83yZjSgOplYVQjhV4CAFz+Q7OR4r9GM
l3zxjTQwmMi/8jEsPm8EVM8Q1GsNQtZTK5NKXVrY90B48OnPt2gA+Auo5DP57kgw
MuFbP3fi7C0D7MyZ3fff8FwaRT5/7IF3kXs5fjFVnHVqNuVetS2tQnpvyRtkeYP6
NvND7pKohrMBYLGJhBJFCfp3OD6FGRsjtsenimZYtW4aipqGj2ozDxAY4F9N9ItK
LTTMNPB98rdt0kVsH+LR6RgIMUMsi4X34Mpe3xoSt5Vk0ZCA8hXyPRafHm60lL7o
cJozRvouBh8JNLgnA/tf4fu6GtsyWnsKG1SbG5Jh73teUpZ+XxCD1rbdaeVcteWW
H3M2XjrJTRPgwpRedvaD+CdZNicChzeyXEbL0ja9F12rupzhy+tb7g8JaThcm9N5
Vd58A6VP88RERXj1jsf2067UbNGk/NPKaYKfuhdF82a20Yl31AngiAP2JXAJ4V8N
tTRktt4ae1yiFxlVart9c9k8419HpLnyBMTrMRqASc6LQxbE/88O6UCqbuZ1q6VI
p0j4GG+SVeLDvwJ/W+s3ER13/+SK+QbGu3QZW/jv4E1gltFiTAHAv9mMZPnXjkEB
w5dkauFk//hM2lp8FU9ul3CWvVZ7oxVVZ9+yn1SPikZQtQ4KQMxc0KjmyuYWwq1O
9yDMZs1hK778QlR0SNBjtPskdRm0Vo0Oa0PLexaLw+pw6d6qqmAx3lEia/wsilrg
C9wDJin/I/uOt6j7jJzrn3eXr3L3Uz4sNZsC2OZjnwv64voKOYmCvXFdmoBSfqoX
5tSO/VOy2/YEbfY8s84g2nVax4VTswTIGNZmxqZ0hegr1QsDDBfADbOwfZVhNmx5
Na3tVm5yYV2GJ95MJXPvhK4XYYlkZk+M7C+T1zbLlV/NW/RWHZZw1AQ15OHYeebT
cFTOU4mnehS5pDqFXfrOXs0q+kFie0CP4MKTnTOtA/dlqUwYHgtzSB2zTjd3Jcoe
NV8y9et9tCwOCQ6YpjnA1kceB6G+6PW7Yj9a6HjfpM6rYD908GUj9cZXUqLMGlfg
H/fcPLHCjVbbk1ZUPvePN9QMTIWdVnNkhZdXKrtFQsUWvcANvUXES06amQ4i2iWJ
fr0ORLMjZqGxcw3NPw6znPfZJ3U1wolx6jyIy8iY1mu2gpdSNWt05eSYu+XDk1aX
8JsAPXi7MzHXgAJTAWtXIaXGwMNc6+c5M8zdbbj3KvtVYGYBCRJD0Okin7jeaJrv
QyNr1YjqTYodcCGWB8IuPObickBuH17nok5O3XB8plHrSER7uD0kjHw12WslSRbo
TD8aDqax9gc7nioAXGY2bvzcIDJR87rcOV32UjXOQu6WxUKZxAMMM0zZlJSyZZz2
mXgMTrzojlBor63Zm27S7h3F2bshkDJfANeCYu12cex1pjCGZg8TjOWZhCZabvEr
lEdPDcOtuyZfliOpR5Sci0N6/Eh+wg0Fm/z9eaK+PlqVk4iRSDXT9EjeRiBgAAlM
2YB31YKBPkFhwJEw47Fj6eq17Dj2YXulDamts2vJQrzOCM3mac2rCv3wLXzdrXud
1PO5OC88deW3zU/cLy8PGwmjO6ukNshQ6BLIKp6EM0PTPcyMr28WcaDD9L8u3/up
f//L5ft6a8r/eVY3jtLPgLaRaFNAhYiFhS2dDIOXY9mmAPjnzbmbIMZSvjA6dz4Q
mBcZtxFnS3J2rOHXcfD2PWU4ZftkrM3rrRK6je6Z8Aq1VgIl2kNjsUU19GrWAm1r
9gY75heN5gWl17EE+KP14uIPkYZSZrV57bLURf5mQ1MkdYSNKb/7ouhY1wTzbI0E
Y5NJ1of0xSArRTTrTXDKKhthDXglYzTkKtUtk7jZE0qEuBzf5G/OzRpKo9JgjXb7
eehioxs4nct/b6hZi8ClkKmGU/t+5WXULs/s5tDP3Zljq+T1CKaqYmaYGJWkh1Dm
vrYHAr0KC4VuVQYeK0BgmRvG3HPFQKp+olT1AFigXfNE+t4i3HwnQcc47mwhJCkh
aUjCPqSVT3TASI8q0del7cjs7kYsAJtc8wE4a3BAPDI0c8qh1oiGhLTHl/4UkFQA
UK8pojlYpv4cTogAAOpIN8Ybf5Eictost7XxTyyIxJRl+XTyM8IIAmkABDMZbC/8
zMmiIjG5kTznvDtuF0BzetdIjhjUFg6WIZjVybhjjkbcKrzcBkN5B/68ajU/ZkSQ
xZI3J5zm6VzAhPogRsCTGwsKBZV+6U9zHwy/56aodzQg95D/p01SBSKHg0mS7/Eu
KSSmOGEBqkVhmaZ25P5cDumV0yVFf7TLzYhCuTk96Bf4nUQemtqG+qYmY/CeHYKs
C++e14N8EqBjWnrq1umezQiFihp2J56qUTAaMrBx2uQGAfrr1H3wn6xzPF9p9lJ1
VabB/eF1pkr4iqpjMmv4bYgvpLGynPAdZzESHbclh0Zrp4SK1oy4LXHms523plAo
9ByfiFTAFL9emAPpXEjwx0ivvAs6fcybDe8GO4ff8XfBEBS5q57RlRLeJXp4bLll
4qEiygfI+HUbq8eCWCMJVKe1tpnXr3tvijDlyf8yoYV0ib0qJCOva4A3e4bBN4CN
/JBb56g33WUsBE89oNoLeB9qiZpEk1eTaDfGBajqQxS5ZuLz9oxWy3phff7TCtvo
NilkOG0CDpD9Zf3PeApaRVNm/oS3aNW3Qlyuz0Lg7vP3nqWNimaNQfmU0xayLXPV
deRML8kfA6nH9s9dGhyppJ9ZgFyDfRaxBysZ1lSDWZd8B3WTSKJclhkNPCQLU695
HcxKyKREJRQukB+FcB0K5Ml20oGj4Hyr3uFwBjVgwIT3qRAbE51zA1kOkEtE2/42
ugjEaCovTXcWzgPDKg+qKOPMU/2nWgggmmGnri7ny34HEkLvj9rKJLgNoU07wuHx
WHy008Mx4CcZh4QUrla5VamBRyneFVYpp+Da+HVE6B68ZhaPL1GgCSrw1mi5uPuY
v1beYJTOAhGijy5Edb53WiYgNDmi69flFf3FDvoOIdQgU4cbK2gb3trv4H9D8hQ1
/JxEJGowQznL3xhx1KzzP1NrCoBV//tsYuK/rD5mQXCmVrIyWQLHLQ+lbkGVZ40K
XwwJNdpi6BJ6UugicnudDhU8OVB1Ls1VWgCrbKTMy1Yz355C1M7jLkbDIjYvyqwX
OLL+LHonhZAlXJVo2YQmoUVVF3TSdIrVO863pSox+eYwytmV7DQFx9d8yLr1wuR7
D42KLP6rhilZB34bD9zqQE9u/0fcFTpXmhAxHiVAy5zHOlygRdlijw99n5NHEEub
3VWArVnE6JW/tkr5ADs0uH4mP74FpPcNy9ReOcaskbjWmd0FOMavaO/Z1H4JYZQp
7ZTcO2al1A/7PGV5AMY5cgoRJ69ntiqXRistFUSyhyNBkdlcuqdx+GqsV3RJF+wU
DrCdVEDrQahpm6mqF4oq/bebnOPAcXf7Bg+Ro1wODv+1hI9YT6fECVKFeEz+Jc0S
FYLUOK00AL927Hbj27LDOW0d2SVEEPWagNfelTffNwVCtOZs2XyL4VxESWi1ziPw
DzJvqSh4AoAX+KlLGO+RC/BJDAvvwEIRr3uPmUDX3NvsU5Dn7+jWq8FLdDaCZZkU
OfxH+KPMvFlo6gaaOXB09M/xp02I/9TW1CUvs+3V5pAaOrJY1wMIOokGNq35C1AL
NjkwXG4rlq94a98F1QYeED7ztW9LyVEQG+auJwsjRR+Qr9Oe2vUyan2zRGT9pzsL
xW1tc00o1LJqJ6MT4bnwzDmqmj+WGIArTsduweyFPc3B1tPiAAUP1GVQ1aqRdsfb
uomb2KteUY2yV6AFrYn0eH8yqtqqCSENKI4MfcbS7M8wI3UGHlPGkGLEjd3/gyzC
7Yn7rSjtjCOEU7Dr5/1QtJIU4PgX23pj/uTVpNiMsU2tVGuQIb8Vxr6rtVbj/Hp1
P1MF7K7XTGBBilzk3v1rlBexact1mV1G3qOfWb16Or52RXbq9PjGUDEMmxX7hah6
t84OxnQnZazcXN2pkwKdDLeHDbLSWFYdh8u9HEoyK4I0NHE/K9xiwXN7o2635sCk
HzQf8b6zlro9igdZ7m4XGRm1peqDzfKWpUsuxp2yVUjcQu/m6uWUE9FGNf6xfs17
TwVV0h4LX0s5rg0mWyCVq/qZqrFglOQxEZrCDaz4Z+oWvXt+AnWs6HBC0HMrojFD
JGbsL9mICvqCarve09KqxZfv7iWPHxrVV5kRXGe1Uq6dOkUPuESc1nDoaIJJ5n/Z
Y8se5B0Wuk5i7XsB3gd4gXveD9z/mlTMaXJ66G+sMJrTwalNeYHZNfLudW24zyKn
EOb+mx7q0Pzh0VGbSYMpw+/zjD2OkzbPtKHaNuwG2Mmo4TFPaQ83BLPHxDiGUgca
YlM9+XtYnNDi+5Tjpu97AdgJSGGfURAuH/M4ncnlLidAQnEBcaebbqB4xNoMlQKE
To1etHiN+nPNhRpqA2Tm0IJVNmDCFtWmTiNDfDgHgu/PC5XBQ4tHJhK7MZZDPHFb
7WYUu2I2tpFVE/TO6wYPHNxwiQOVZFXCteCI1Fpb0u/dTAn07NPX6VIYhVSnQ/1P
TuCSxpGLP6U6vExeN3Glfvl9P5hEpKHik6gZH0rOenrsp/KxbyYpYksINHOH54Pm
i/z8eGvEOjG0+Szc5OGMrjVQxIcxkyhVN/UvY2PCjclQ9gzp0UsZpjVt7P10mp8p
2/Cjy7foo5tUwws1PnUP8N4NH17Llq6S+swDFGTvblrjbXXhRCcwNQbnSt9iD5yQ
dh/K6BfJseDd1ZNkSTv8wufXIuH0UdLIJbaatJjOWz93zMBK2oHvHs9WbMjMXpOc
Kn2hQeH+ayXb8HELuW91uYHYUriwc+dM7B3GWUbC7Kt/aOCaks7rX07nJN2iuICi
iQhm57G2hH8pbtWR0gf/h6F/R7BiR17coaoQ1Q+DzvDfeHdVdfYQmf4MV7OdoViA
+6/qj8swjTWz7i5QTJOxI/kqQUpLU73umOLyB9BeUy74ZAxJwHO0m3sGtpZjkrC1
O+kRotOAYpCh6rmQPmu3Q/kyD2tAJIdbB8g6BQ6l5rXZS8DOHQ4kia4yLy3VvY3i
GlPUwkqTWfvcgV3WgER3W9EZjsJtibHPgTRNREdizmGL2ZuQ05BV1g8BErSTzewg
ZzRE/Q197sMUmppsblJkk/qaV8YabfOcaqOGbiZ89jUsRdCShzYvY8Vs+CnotY5J
OiPW/KoquwhWjYBYbYokKwPDsnm3ojgNeYDfwyAMPLasU0QE5pUeFV1GvUzekUtO
T1envfDSV6qusryHI5F0tKOGHB4XbGJh6yVAd5Dbd33fKKzu2Bw/VC1Gfx8Vzjcf
eLnbAp0ikpo7mvZiz2iueDXoTS0ISVaCnGqIUBeDnJVyda/Yq9qCxF+5lyhocRlc
aSWJheb/I4UAuw2hYi2f8BZlJNLc3S1kIHwELMPh5NvcaoR6QJmbFoCeRJoIY5XA
DNyVSJ2LkOFQHXCobafsPaEmBJFgof7+zDv8t/B/N714dQ5z3gbBMZcIUOnzEJsY
A0xbIGNyT0V+d7Xj/sl98qcBNx5/FhbM9lrp1EPuUN9uYjdJ7oAlB6SdMCN10EKz
RAKYaYrDbaWc+SqYyqpXdye1qFzXDTwDVMzXpVjEPxnoe5JeFDGskJVllUJ7Hoih
vO6rPp8t0XuT9LruwaOuRG5CmoLdLjuQAXnZHTh6CAEI4lBZEppB4yq0Zii4qc8x
LchOLPsymN3erQ111vlPtbGPSMs6QGvPwVO9rFs6+KP3Tn/5i0Qxn2AXxm6vGBSG
0gu5rpW3DcamMdWTEbievhvAqReHHYNDB/qCImYuNUX5uMTMUffqMIwzjFWZ4U1v
chJowKPxkkBrw6y0W/7QlcujLYjs50jXDdfMDTHbjmXsAysOH0q8NaaW8ADU1fb9
bQmEd3QVub34TLUmTCFjuHlTAExwkjRjzxoGof3+5mD2NvLAVDPXQo3lL0EJ++uB
af12YxF8qXhqf8yXQzS/FTWiR3UCFvJxTvj+50aBWx2s8dRULveMVKFpfOiH3vrU
wJm1rsx8RZNP0qJApsZ9wfME6v/EYBBu1oAoD7Df7/jXbEjAgvPZA2Z7C41Bo0zo
f57S/UeAj9b+iRUpR6njCYgCptfq9qx/nk4zc6TfQfcJEwjyOc7AArGyYf0je46G
thYSG/4dLaS6jw1kSEIisOKvw7H4t4oQxw5kcC5IOZKXY8C2CsT7P6pE43248mb/
67x2jyG+jUMzTj++whk7pxjvMmai/sJyJAqayBffK5Ar+LHTXZ2FJSg4Vwnn/Aru
+nkQLcNZnGwhQCb10jy0EEaNvhxRfuL+dSPquPpO2wpHF0SCOvFP7TzAvyBRAyHU
gze7sGlHzi9gxss5CQNbDCJvE7tSxZpogHhE6e7fquRsRfg18gFQmkwrhM9cG/cZ
TBYHqknenR4EPpcUHs0YpRF+M42FfkSK1tcTLdNho5f1ps665YOteRpPiWrc27yG
rYNc8Mlb74vuAPrZrTJXOdTh7qaaVLlTXCtgljs7xYyzqI0V0kKbgO0yCFGqpmqt
NH5Ky/0AR/YaOxtpqv5K0a88/uRcReCBLquwg3jD5Au4X2nwNUZ15I2uBCnourqb
ZkprtrnHPJ3A8Njq0l+WHSRWGN+Y1FgLjbCWyRi/re8ZwXg/6srcC3EcORKPx5oK
1fZg2whe40DDmCGuD259iKWXFqVF9Z+AEPoOw/+dqeBJJhm1YPfJwzJjWpZX4UTL
jf8Kq7Umbbak6t7FxGcgqLKKFWq45Sh2Uoc15gPoA2I/mFzefGgKSuyJGZ4oaXfw
1ABWqNZ9jayLoz1y009CB4RUGHVIqZnjXcRPGjtuGSnEX8k8tELcugb5lXnPpq4m
G0rgNm+hpWlgnl3XzBx644Kn/M4vFQmP9QoHX0it72DSzEh/V4UUVGXJ+lvi9mav
5jG7gpqO44Upl7iXzTFdBGrGiRTLnDYhVLe1+MR9O9+oj0hUQkyVk8dPrW2o4W1f
K0r5CaII1CyhGhIjLBRAoHp6PTWLUAIAPdHFEkPtm6l+0CNmS8qQEB0Aw1XVTkvl
6HLBO8+8NTVzr+yeQTiKSCpjPvfy5P1/ALQLAys2Y6CWwqNRlYbYtPwnsz+A4KeC
tNFOEKFcK3WbBpY/ZHxUcJhks6Z829FUPmBz2Yz/Wn/3r+vgPFCLGflSd4IabU9q
PmkIMiSUFyj9eB/xf+md0+E3YGI5XtqL70eZ3qyLTLCxlMKVwj0j7ygaOw0yJwTQ
zEjEDuqjZhYWpOYQ2j1vhXbE6IBE/KXnRmwBPYe91wphWI7xH8YRyD33OWSk0E3i
A64W+o+PzVmvyDO9Fmipklz4fuk4JCAZK9buIoRXkNOgSxUJNL1oXkzjb2iOg0iv
6XrSSA8YDy98t9LC2d4eDjVMKRUU0UcHrsw//wQq12VginTLAQVPQrMuHaGmFUKb
G2sI8bI01iaJeUpbYnar72XdszbhW3Difmcy6TXCrqJ997txL05D1Ka544+Bt83b
PzigYfjyP3gRrhfae3VA6A9WYiqnXRw9nJxtUyONz+PDQs8X0z4JUEaSHHZ3VN37
Wtm2dEWwzQxFF+61iFC4aJgyDK+GTLEwTWfsy0EgDB7NETgkP2HMYmsp10p19hin
koCXz3CE/dSf0np7+c/DyPX0qxvM8PN5MvrRcn8+4eSbOugPuENRtezO2thRSuH4
HzIiSkf5vnsIKhUogQDTukpx2tGvBajvdvKKZaiYASVadsLTJJyF/7fs1HNh6/3T
vg3IT46TXtybHyxNReK2QXgl/53zEAu5buwJIX2Zyly32LnIy0uwdSoHuKRoRk8g
gc10puglpRMg98Ub7KCPXSjzmW0Qeh2JMJt0pcK8TdmSlMIiP+Xat5Ji2JytIJre
MQTYA2iiZyaUZdFP+Wm8wISgYIjh1ZYzTl9HTjWRF2ezfxIHUnSsZ3PPMU48ZnFB
sWwwzwaf7TFu5mQOE/vu4HcC624wWwy5T6ohtYUhqfeTt1+DQEJGlwm5y5zO2Tps
TiAysRa/VhimUn2ratKXW0fR1BxhzpLv9T2Eh6ri1pwN59XEM9NF7YL9NJJKA7cW
xyAGzPqzFQ4MXYuIottMEhgMarFye/czUmeUESK46MdFYtmySNiE8GuduBguyzW7
S7MeAn5PTHzyf2zb/qMWtNzjphBdyAsiXXmAjg61GArhA7gu67EMSk4L7BOWWznM
FfDyius2hdth51JI1K8urTD/TbkMvl+tCM7ME47VxGOOhYUwCwF1ecnXfuRg63sK
5e9fYXpOYBr8exI24VSxoDHbDck/81vOabhbRaYPo+0YgqeUO0Cdl14bJBtM9iR5
I7qTg60DyDxiNlBYQeoUFZ7sie+yd7Js04CHdR7f2eIeVcnlR0AOwcRNrI3YXZ/c
T3Y7GB8HPVj3XxbhHLwXacjcMIWsSIEqKCipQLcPwzozfWlt+na8dWHmzcxsKtj5
WrabJUkJZgyxkDWGeBEDEZTZxs/sqGqJlhX5Hwjs7nIJ44ciwFpSaO4CV2A4ysdn
079k0F//d8JLqK78YM7ulAfHk50ChvWCz0+3WWSjuW8h1C96yi1P+Dd9WdbRJ80N
eAljSpdEZpkC5qt3v9URif3/IdChfdN+8dYz+tf80G15Mwj2yHuYE4lCow8qWa7k
sRzxfoYfdPoj0H15OkkCEDePyW630Zj5C+zXzKYoHa4Uo1tuJDcp7HCnT/1Q7S7o
SYeMZ1b9ExQCwOD39khdLiHZJ+BXzOoD5OHBrin+k91pisnDOwL7Gcz3UfRwrt8B
tDBF/xyPppYczu2QrsyCARyWx1yXOh7Rtd5dHgSnbaUmThgxLdk4MsO6Ny2/b/+9
LMkkTCpIj4lMSuJVUNiLV1Ymab/NAzHj2d1UCg9x7LK3m6btkghA+GmDLDEuZHsH
HDwcXFWOivyU0fmnvtLgsrOYv2M0qez9U/2yBd4j4Fq+Is0+hXd1Pen4UlS59Ouo
jWx5Wpss/m3zAgXABHgjr7qpLfW7De4hIvU+12dxUk5GxKuHOxdoExCJm6swIjMS
HBEqUVNL6Seg0g4HFhyNCQ52PocDdkq1cJzpukbiTa66X+8sXLq1byp/zAJeqlFU
3YT2Ac5JxRoWKozrPYinxtlCBy9CnJGkFxqMTI4wfi8Aq/878IYXT1ha/8HVA/xz
aq1PJj+ojJY2YFzfDPBQOaVqhlyzi97GpjFylNdvYLxfHLdjun5bi3rUsyEHg95D
AhkFOq/M4HHdf7qAs3RnkDrlvORLiAp7FLtJR+v7y+4NwinDNXiTvL1JgGoscQis
m2mI8SzDrwCwvLKajc2IRSVw26JZMc8ScY/n073b4xw6bjgkMB+GSQ6SOiQzKfGm
R0D5inNOKuNe7l/ffcvVgR/kkevKT8GaWqIGqpAPXZ8rq1WjcmrDyYFTLWbnVgTa
HwXbBhca3Zg8pfukvuVBxVAvj3Wg/heAjKjxHCemCYCdgDA0utBt/4Pcl4Ksl5D3
cNPHeJJHgvQcEfbp5dhU/L1gjBbS/SwItsBnBAeGapF2Zx4pg/KdUp7ReUNQCeAg
3G5uk2lHRtvjj3u6qxtE1bgU09fA6wIYVubmTVSsTot3Dl+tsnGV2XN7M86c00+B
JEQAsFvsdZU2/GdGMaeKYT3P+upRwiMcXYJ982T7o0m+RNqk69Ad7utIHscPJtf8
RZ2+0UKMiK4S+0msTowAGnH1YzCiNMpXxVm6aicuHnt+fOY0vj+6dtfmYHAInMbo
HooUjLtezJUJ0GC5OmMtiVstjtrT+F3F+do/34meoO/M55kDurhOWNHszQCXCpOM
K/w0q1purzcsdqiXX/O2MfcZZJzmk2YhfueRAgVnriFWbYO0ZUgU6M31r9Cl0ny4
8LUccMTGTVXFVBX5R85/pwkaiv5qw7780WbfklfHGmRJTtRCr3nnmRGRz1hDIqdL
FTVSXpa1kzktHg1zTtiwBRwQ/SlV1E/Zbdb+MpPuSmfyaiBAbs4lFKohplv4GBKD
ilbGK3YFX0k83kcrs9ZkwkzmpTAh9EiDRn0u5QWtCyh8iC5pkXVFRQfjAXcEIGFI
CDuEovbmnzL7ii72Vp1hDbCRG6SKfZ8ufdWvVE62HtaXn/GE6cClZ3PRcpEbvwz5
WTPzwfQFgy2i6L5XNKaARjXbHhExLpf/FoFBFI9o3BjxYNc22UInPefYWcZuHBdl
5dh3YD6EN3WEJhsLbSMhNw5VCZTon2VM6nApY3OgxmgW48CHfA8JVIdHi2/GrcKX
eB2jgH+F9UHudw2g1+V3ZP2ykT101Em5q1zzx5Aou0LVTAvfDG913DQPAcopij8I
Knufn2zYdrZdQFbr7bOceDGEI5ZmXQflZyTBAX6PtHnyzKVIwAx1dqtg/VNWM0YJ
JJXX61thUc3Evs2Eq9OKJPRQPbkS7Hf84mrnix1kudVp+2i3N3huo6+LW7nECyT0
gSQogH6TL6Vu2woUyqNmtYMjDoOwe3bMwi7nad+ollweXAAZorVNWMAHDr6EbUVJ
uayjIXju/HpIp9qtYU6VY825o1TTdYNcGcF0nYF+O8e7uR5d+Vnl+XHzbQvgomQT
JX5XcqkTjpeJywazon2ao+s3bouBE7yRBIhjowRd1Wc+6F0JpcbwQrcN3GwPazg/
QALc+ufdMKN0DLjvG77rR8CyueVaEPKFFMldTXkdVqzM8ffw8iNe0vm6bsurdYPk
gY+jyYFO78rR7xEnWQmW4w8lvpw0FPRW7gYXb4LjNW5EKCLperYBiKU9CQgLxl4Z
1fKTL8fuPqExLna3SgPoysbNoOvPpChnxCy4oMhiVmBb+aLYgcFWQQK5s8ADAMQx
AG+Doq+VZxxv+KnBJpvxf3mBai5oHc4mhFKCpntcb+50Yl468Ywzx3w4SmWLQmqA
UKHJBKHBUK0PGLlRhJp5WXZ0f/MR92vdidfihiGC2xMwTlmMdInF1ZNeU2/QROHZ
otgn4SvNPBUPGWAFp+rtV3Od65R68DehI5zcjrieY78vh3oMmWFbLawCmstQRppD
b4idKi44QOYzaQReRT2fXsXqo8i/o6juX16QwMwFcTLtVNDlgmp5HEBvkT17Sxun
0zrPHu695EXPPs7f/5H8xEYKF4czoxYnuvpaCuUy3Z3d3YO4AdNRre8+EP1xTlsQ
pIwq4rGBYdDtt2KzxPEC7eUAK/TuyUR+hJfIZ15PQYxhUfbVpgWssiTHKZbcXCH5
4pj/xmXX4KvMAsa5ypRl1cZ6s8kXquY73KKwS5JbAj9omJKajJpzVzbmkUDmKmTF
LltloGzzqG64sKk2laIEQdvx6yKHQ8LyOIHKUzkzBDIL8CuX5i65+WmUgTYZNH28
HfJhUQWuxFMcINbNvUUj+LkpjWkVCBApGT9vGTbDwdwqg4TGfh6NT2q/krv+gZZ6
esF1FPU/I8HdzVZf6R927ORJNc21Qqb8ZEjtXzuq9Fw0xIhVx9HCtIQ+/VkSbga9
CbRpNjxHcVJc3bK9Q3OAiqdk93CP3jBoSi3W14v+0rBNEEkTQeD/34qbvWs9xTlO
jL+R1YvNuwvm70ocPySc0gNWadspRrnDKhsk+0uziaV0U+28JkhvOkUK6yCbrsZJ
OBzp75p5E/yOdSGeevCBVEoS3lUw2qXB+YKmNMH/RqaRgw+Ckk609T+qHtRmOxzP
rchmV3ygKvHda8VkubQlPbnF/K++idWNSb8qnXSMufNCIOSKykIieufbsginG2m3
f4r9j4sZuVJ6dwALMvFqWiPe+ZfLQ8SygXqMQARIJGIml8I4PkPhF17n7A9tRhoq
2PsRxewFASXD/anOKZ6bV1GwTMl4hhuZ0A+yskJ9N0GG5zevW+9cfKwEQXuFcjAz
VPwgCLhooKLQbQAsSlaVHnihPFrrF8C6SMfok2zR5xhXARJYyCB48lvWdKdNX/CA
W5KXPz52F8XOK+/h60oa9wZstilRte5g8UUPZKlosPvtRvnh2lQ+XkQ0h9AN+Y2I
z37eQkedEqmJcVqUnSTUUAUHtCRnxG+Sq2CMNUG3ykyf4M02wsMp9lYAJ2XxFntR
H7RabZJemmPouUEc0kdvdJN9//ewABc3s8BofYXRsm1MyWMUo/aGX3aDCEpLODT5
MU8WVSwJXu2zSZbgMBvluOkpsZ3yysFoBei1qNico0/okNCHFSaF9EfFmJtWnlJB
5EyzyjZCdHwgX9gKGS5rSGaSEKR1xSFXs3phaRykNkzjVys2r7cu25eOid50tpIj
H2oekKzcS9qPx9OW421qEQf5OzooQ110kbuVE8CwBbc3/7+ks4fY3nFQEhCsR0MW
6YX2FBsOom/yEOQ+zsssD+YBkFdnFxv1dtyzq471kWKRGWQ1OVcT6dv+1hoQr+Qp
TCSX8kjsJff4rajDeTAdfv25l3li60GQkb5L9ODqVDaDKXwPw/CzuWHqfl8QwYn+
SavGf9JZj8UcGjzfBLcrxFSeQM8lSwmmwM4wy2d3nq1meAwh2j0+VGSGlTFaOx7Z
DLLRLzSMGmN+17WRL6NpfEHnoSIvktcUg90o+C5khn86RgiwErV33/0LyjXAfi5c
PlGR570v76D9Lepq92+dXgt05z06l6Dshzf9/DeM4zwEqqbDpmO45KVASipwzdm/
8cPA2XRWBAeRFP8V01JM/M9Tul+uKxLsjjpb1oJUuc4BF0LheIb81rVDnzVPXecQ
h7oJtLqkFoYDHMvXjAkbgNuHIbjhQURAOLb4UjUdrNkYRcMHtCTIckBPw3kK/Xc5
nG6YEn3ab+DzSa6/mNHCd2EzhygB5gYP1HR77rhspr9Rm5rjYg+sIIxAcIVXMNmO
zQ16AK3L+n3EPOW8MT1+N3uGJ4kISlK2cfFgDjpgf0Hn/gP4cJ1peX5Q5kkh6jPq
4pEFQzbTx54RV2WFdTN8nQuihYX3MMHr4OPoitb44x+I1lgkJ5ypqz8xwqDKvgsz
t/uUcCwW2UF8MySMsi7TM37FQ8S6mw0XNwFBhyz7vjA+QJY8uaOVTzpw8fgGn7jV
N2BV16tBwesEgNhPzThMEL+ESxfIDv+IoD0XorVftwaLNU9XzPHVcVK05SpLgnYF
mjKNxbd36ypqM8qzXOfxvcNqzq6FZf/RopzidPJsqIRu9AxBw0miEuH2SyirT30n
O7OXPgadQxn2TIh6uDgd/s2u/PbMJHnez3dwkxtTNn7sPIhr9l02SZfhk5cxcf8u
QyN1c1AzgFgX44EI7uxBeq3jv8TC9f7InwhEJN1XryRxr/qI4QfhQNvOKPUB0gdb
SeRFGsY+4UQke6BVJAvcNKBg0rfFET2OWm8tWTbv9Ir3/2WFV1ViYMeOPG+cu4Z+
hanEa/MJvv5+D3171iJWgxT7J3o+5H5aU4hIjxTYKJl0FBhmwXcMBRtj2KrIL+ut
6BukmUa4UFSLGMruI9S5jGeab+wyn8RppIf3B/gaEi6pegJBE/rimfhrrid8ibeb
tlZO0Qf7G0qEwbiX5Z/oUWieVD9b44tqLXHGzhOPxG7SHx+WwlZ1K8UyBfAOpHCE
XXE26luNydAhFTP5Gsob5nsOJLQPpPoPmkBxce9Lw3dmM0EhugXWSUzhHuhDb/BS
/zN2r1M178NTwfz+fe+MeL4ylUcnjECeVSLX8DsDZ2plV7rIo0hAmGIyS/yZFQr7
EXWwbu7+fbVAVf9o/RdY5cwLUabnelrCMkUsqjDyy9O0PIKOfxmxb/SQ17Rrv8xd
8Pb7VCxlFgWWmfyEtOVJbByRuq2QQQqLgMmv5xASHJSC9iX++Ng6RWjdwgrZw9dI
I5VBo3rN3Cr//0fWD2eYzNRN5XtV/tlHeikjGXZnnnFku5V5ViFSul28Fzfz0QsO
8+tkIfyXdgYQ9RY9rPt+qb3eIrz/F4cH30B3PoO4lDQ0at7HCwcXKe/8ItazDmz4
+2Ll6JvPA8h/sskiMh2OFX3ALVcatNrnccbOzfBhosq+gsFOJHLCPCi9JRxX4wH9
AcjoASXTssL4hrZuMkdwFsebf5pW6qxWTnOcCr4cEkZfCe1O8UjzgbIkFZz6ckz0
7WMNnfZZiQn1cTE5pgDSqOvwsLNoIpg9jywmFQT/wDJqTohAbuN/9VqF0btGrvm4
VZsFYs1tCmqtQTYNhKV2nxGNYkYKkF1hRqxe5On+LCLW6RNCGouI7me48qXROk8j
H+AnK6kTFKe74fVySrXR+kKFmFNFwq+/sLYWSy/qHv67sHhzG57RPxdYvFDB/WsW
1oRh91CvINSdJ9kM1Y7kxBUIG7TF2tfVQFlzNjBS0kW52ue8v2t8b3uXZ9ta3EfK
YbKp6cnmNxclv0P6G42o4YgZ/bsY4QWSB45dOEKCFZjUZFyTRWzU59bDqv0qftBe
ds6Bw0Zl1tR7mQKhzSb3eoxF0DuosXv8TJUG4ubBWezy43KyGTJHN7X8AzEUUo4m
nySnVj6JQAnOmbXigekRjS/mnD4z+S0GpxUA8m2wJXKXXzvMRN26Z6lrA1/vGTA3
hXl0O0byxhYlW+7SB7xWvz/6KPCdGyuJphBUt3R5EpV5IsrSUquDQYbTLi/77GiN
RDE4EdxtP6jyFP1pWL/Qw8L57N9x6TZTaJ8aG8ewN0kLk2PJpY2gOvpD9bp2gJBu
sB1PrcMBxf4v/twhiYdSzNSvtzWH8zHgtdD0KXo5/AZ7bcw9V9nfY9sNvKzmjjL0
GVFACD1RubpOmoCKs8UYzYVqAOMCXH65lhHYOCcIYs5kgDy4/jXGBTUnwYZrZNuU
lZYofv3ToS7xaJhY5Q+0bhmMV1Kl0RoQe4V2ZBqKOOd0k5jRl6WcVzgCkgm32cN9
na421LNA4Bf9pM3onW0QfJ1TZ3IlrvmU9hDPZTzRZBr5B1HRmzaWdZnILMnM1k5b
6msFLf4pGjuo42JurIaDS68Qeuig0xkxXWOsRUhpCgmVSTDIN2S4VDXCkSDzRjbU
pgr3gCVQIypfx1Q/p319kF9JiL8MG9aNOaAt8YfbcG/KPYaTHFLgdwxg3GW9tUc1
hLz/YNpF3Chud/Q0QTnazIVzB5i3RrxZ/XxodblzmCgsojkLpLYMQQKbfylRY+Rx
qrIQFORyLzVsIqyHCkD3jvNYoLwHwFK+BYFZKIOCRHi1wwD6ZY5mz/H5kCAPxFU6
ibMWEdvat/40edCLd2jVbPiSEV5ut3N8z1XlR6WkL257kmXsuHgb3d1oyKRg1Dqw
nIAYRaC4lEoH5UKv7njRPctWxFjzwePqaFBsN5EGo983rdvp5cLQHKJd9L4R5PnL
dROSyxTt+/Zg5C80lX+TbxU7SJgBBLFRJ8F0/uwjEwvXLUMxpfsvZQvwnp1VHQ6c
fBOOPBSBqjGucBsG8Pcqtbj4fC2hyNvcOKZklsQcbApWlVBnV/ilAsSi8WQgCLT2
CL73J3F15nvT0qBDx4shJTMkBDuj45Pa7uO9PvMWca7xuhvIo/KWI4A0kTHGjQ9E
CCcI3qc/aBHC/DHWrLVvCQHqQ3S4mUaivpfM9Sp/Udnfmu3ntSZvJn8n2OLyDQA1
TDmfCf/5MedgodlftFUzyuCgvB++HirRB2HHC8aPs4tRLzzXYsqvtt3leixBya+9
YgkdlUS7b5u+J4sk9HMwOZOweWbTBi6yuXULTk78/o1fpi1QrwztQBD5DoEPehCO
2unG5csaoMYDRx3z0c6jGaYPFpTdd3NcBs1RGKV9Z7iPix/4tVAXgqX57SH2nh6Y
/lnyMA396TWKQ9A0EHA9gUo6ILh1TnNAkBs0kP4SFK9acryAQTEyW4+QmVCBWXFG
e1XTXm+1K91NTWD6zvGyxV+XMHrmOEdGRvHgUeI+ZQebiK9lksBolsJNAaOUm/+8
sHWCZe0blfB3aqSp8C3IESdLi930kPHhFqu8/LdQdAQGDCKmWdIcPWXGPqmyxl6d
R9sON5kMPpIfJJn3u4K3XFsBnx5HwKgWoi/HBTj36HU8kJV9+Ca4zVqC2WeBx+KB
67ySFF1jbgk0TWS0u7/V+aYX7T6WLO3NoaV965LapY5x9Oh5EqzAGVaWhGRWaXYI
NlDrgS0UeHr1gr0FHqhb5temmAujYBvQIImMOjlo/jrARpn2rIbugUrxy4khXcnT
q77PeWGf3Kjb+rD5N0rR5iCkFotjb80KfwyVUMVlXFlgordRTvQpJECOsc8zFBgz
mU6yM4Qw6sC019x3evMypYSoD/ePT6f5uWhm1M4aH2Zy5EcvRmw/0hR9aG1zweKg
f12Vq2o2YabbZHNG1smIYcBSnwLANIUj6VzY3UuqxuLMLVL0pAr0MjlQpJ6u1P3C
veT0s6di+XhW11CzyC/8TZTOmOACfNip3TX9Mq2Bn4kxPIUxb4WIrreMjFUnLRey
3eN9IGJeydrHf1bBs2F9Eajhys3BkbbZrUUnG3ve4+f/jFqI2ts1r/TAnEifbF9w
xdOZRbNSF/JbUSczPl8EuUAml0UDnANmci35oUuUgXpNeAEeFIKFoIX/rpHh8iwr
4igxZmdWCwMnhuCeg9Lslk2iDRC7zPgfB4GNsUxCvm2Zn3J5EdkTz9p5xlsLd3Yi
EYkFYxJ3nXxts4eIhxLHli+0bpK7nbMqjN7vsBtuL0yS8rVaJrNp91pU431kCLue
hkQM3pN83uiBCfIAdyUHHVcUnvEGu1GY/OteDE1nhlXKcE3G9u7JiaLlXniebKvq
GV5hXuKPpE371VtSlhgVeJkFrPh1Bt3V3WSA1Q4julBF5m3UndJ7meGVDPou71Xu
R+3T35K8oCLnW183ALp7a7bKPCyEQkHvIK5ZU1MJg8GmL1I3YH8vRY0hb3qI2itr
x4Aj+1XEMehzXlDb0kNruOhREgOUIrgDAr0em8MUDUphlmH1dkWKeVkCLAfKCmTm
JDjg6Jm/k+KDvmzAF88wIUiqdC9dr11+zN10PNz8I16qqfIqEIaDu+RsYdaSPEww
cGWaZLVrWQi3h4d6MkqvLT9u+xHgU48wof7tHElzgO7+wpybxYzWdO21nWwthw2h
RIuMT1eT/gUhQcQ53fW1KsShavoB+WSlGkxzvwSU/NZWa7MmCv4+ZQuMeNsrnJRq
zN2YKo94X/n1Dy41B9k0E0MeHcfkT6Qx+Tv9OQPby6QGtBxV/EEYjuyULAeRHHqf
utp5vZsuW8MiU1LWlxpBuVQRom8iNadPHk1RD29V7MFFZ6UjpjW71iUQ1JdIlwve
kBH3r/KX8JXvRwuF1CbmlY/1g2UIodCaVOVdUbwwq3nzvtQZdZcvTpZgXyagINKq
Rox1EtKHp9vm1Gu+4Xy2JngfFTpbzRH47xxeZdbZUqoExSt14WonU2L+dsovlDPm
Axtoq/mNyPlXHY1XYGJwwhEceJ9r2wpu0WSiibLNLqkm3fG1gr8b+gUH9Gjdr/2n
ZOzqRRiWm9o8JwtZD3h/HdCLQbBoA+M3WUR1atE5UDqCVZNhjHmaPX5370lK2iOZ
ERF46VJMPchu99fgAmfS7YuBRZrX7za/apvBDMWzuES32yWLQTSRtr5pTbNw2ryZ
pa19NxbGn9EHzBX7CohB0qFG5wYWbKDts4JSCorkIqX8ilfRqMCXfBS/ip2PoYCD
Uwv8L2rmpJ4HZkgIXb1YAnQrfdfEqAqvffLfZbHpp4w8tooVj9eluyzp8ukuzuzV
VC1/PszwEWXWWb8+jb5b1PHfVATgwLYh8Y33X9gSkTslZQZVkJhdMIJgNBu+jqR1
e4rdU/JSm7JtlOMQ6y3OT0ou/Q2VRW64MCRqFQxY8RjV9lVdKAjwrQqdTSCqv31Y
ANsegFsxNmVS0U6Z/wqlnjnShEcpcnhHFXaHbQJym3g2c87gMNik7oBCM7wjQzlu
OBivF3w01YV25QwEVoBMzkqpudxwTqN54Vox/CibiY5/IUBg1KJC8r6Nfk1hqe1V
6jEQW9SoE/krgv1DMLoYOwXaolFcvV6xNe4xyo8p0dtviLUmQmG3X4Gyylg85pmn
aFTpL84kE9hE82F20OgH6Z/BGv8eRAu4laM43+Rre+iGOl921dEhZ6WlBw5m3jiI
+ynClFcxDgvGvojHs9ipcrXXvUDtJKsdRdjBuZ5jyyKGP3OjgWrWsVzVmz5hJZJE
VANc3ivM8f+xa9qsKTP/Dnv5RhxcJdFr+FgWk8RZYWgo9WRnb8IRRjD1uOtJDPXs
HOjOerYtFNQgA7zqShKtY3G9X2fAJt8UCNKD5T0xeE6kiSyhhS1PoyvKB4LVp26X
GDGjAO4PfcFxDsH2cuCRkmXfhN/qnANbH+h+UKIhKEWAueAlwPAYWbmxRWOl//Or
6+q1INjfnu6rm1PM3jRYDzJU7aXtoO5nKiwVmWHRVYxbFgT5KAyjsVDPuFgDJ5GV
OCJY5QpLsdwoexxwjZQOZl3bpEi6b4HT+y2UCG5y2Urw/WA9cZPaxTtvMVnRrrjg
2X/Wx1aR8CJuN9WT/C4nfPpV5eudPY755TspxL6Za4UcgPqzxXkV3WXt/YZQBl2P
woxGZhilBBp8D7RSZQhiQLEm41eG4vSgD701AcU45895WQL3Qhzvfb1jybb6tuDO
H0oCF78OrRq87iljbiOj/lKs3e8wyiX11ULnHjGBDJGVG7qh1HS8bgOZPfeQ68qd
TJ+i4R5wMeY8NfBco930zjL0vtOeOkFiWYtdaGNFGXaLjpm6LMcFz6UR56uP1pW0
S1BEjTMFqUjPiDYIMjDqdZIpdo//StwRaqK9YIbcViGq5O6Bl40RXjB460qlAV1r
1S7OnIb0HiXM53hLT/NxLya6mpcHgES5l0xEX+Ma3VpZ2k+WdI9/BFmJBeJyZgpI
/JdU9gFzVRl71VsWfqj1aqnE9X1DujN8OhuOT6YWI810B8MiXeW2ED6CfoJAO3Vz
ggPTMawCzQ17a5nXCv3cavBEUbKRctpAIN3ZOFVK6ESuSLecRylMmcieooDFWVc6
b2n5lgt4dw0jLsGgI/qxcLKGzGH5WcIb73/UYOTI5ZzDtGHHJZk6HXWeRv9W3KZn
I/TNFY9VAVq87mRhUXKGNALJp7DxwqaOr0YC5Lbm+Y6NK73aaTOXM0zMc/3NZBJC
jE7cUnSvstGkue6verBq431spCSkOyaeOJHRj/ahjrU9zbQTdX9T1ZrHqMykDHev
kF+3Geo/nm38/UtXgtFETjnKFMGLNyIAt3FI+pPlJa4+YiObJzmFcGz7tghXZdDn
MBkpuNd8L1Lh4bZSG/8uafd0vUOlZQgbjjjDEMx2IRdFP+liFUJZWdjf3c0mE5cY
J+Tyzh3GeKYOfSHmeY7Ya9V2L4VoJ+4eSQC/WAsCh9g+dt7bt5YkVTLPK70oENsI
388zWZEgvg1lutKs4RWSxnKABnyqjkbq87ZrRhEzlhWMZiU9/tLM6u1hzdVM/us1
pUyOfJ8CfIe5s91DbUERqrR2xto9WQfUdCMjygoXb46/ncQVoOD3gfKzVeVVeZ6+
2crlR0kEo+inubQ35lwX8j6iMPNYyNn+JGZWSZoTJKZCEQn+3ONrZD6rfAZY6nkY
I7Y+YNchG0/CUbUcUk7Kwbck+jQ7EtooHCdbAaZBCs2g4jvC0R9xLies3RlueW67
Iq6flRk5m4bfTnxUSivuKbH6Bs9SHstSBjo0aCp4qtlmLDMPc5icZc6Z0/EKM2FV
bcLgmX/Ya/hGeXloXif60UCT9XijJJ//mPrTSoPYo1k6aEFMhsl/KfMIhcidNqFa
YNjB4LBaKy3urEu8sAfJlnjlXs39MH0w5xHV1Hl4wjHFHdyUjXCFluR6AJgCsqTY
w3/8QFpnGK84rKf5Kn/R9g46B4cw3YMopi1i10MzTLsMZwu0qqLdG/YYgLZGREW7
4sQaJjqBK5fyCudYKzNE0xUF2GNiUeZT6nzuTCm0dTvnTTC7X8dldEiXggnZTFzL
AUtbMDx2HZL4Ely+uyYWq7BNAqeeQKvx44FhYttGAXws7GT7EYBucC2IrAlbGb36
QTln0zl9sW5hbtZAZaMFNy0nnGhxBdg/Gt+xTtLWAARIUmQz+t0rymMj9LyOIYBW
OsZt1E4qlUfuPhcE+CL7mHH+EiCFd9OWFE0ohr652Tk6+uyFblob+3R7l5qzH7LA
tiasxKD8VeBQ7No3G/sryDLrPXzbHpn0+1plu+tvhaSkTTEDBTEGSI6axUJ4Hgxh
BcB7OICdtUOdWpFmE78UyxBqpxIIMaJpfAHMEPOziLwCBHu50maYAXGsk08gkJ9z
UcLkASklpAcJLVyuM5RlQ6acTJ3Z2KTlFmPPMmkv3VLPk1FkmM7qrO3Syb/PsklV
BBjqMNTnkgSgYhc++mPMeB1uoMh/XJh0JEqrah5dWB8Gjjd+u1QQg6C232jvt5Dm
8n7xrUzhkOk5ddgJTYoFCla+5DBkt2DhlGIvqmv1QidKRgtY1r8qsNf8awC1xadX
8hysKCqUUUP1DrRBiQYX+72Yp+cl6io7PeouM8Yddqv+Bo7XGnZlwFHPZFaggaSV
CC2uyVR9Wrn0y6HInp6fuwi4mKzeF4OU/kizvRHc7QZTEq3KV21tGm3pe/k0+fHM
SGmusAw+3E2dhtjLexrJR9tKAnhyjqG8+KG48mdurH8KIdRs1jYmxJ/tGBO0RSeu
4S//gva+oQD7ZEhmJlxwuP/xjJX8fvgdf4HP8g83OuJ7KyJ4fFj6iVWOMEe5/jPE
ymtVgFd/FCOeyngefszHYl64klks4fY3QH9S4R9UFqq84YELcCaqXazQDRhkwHXY
Vql25+S1Pgloc7u8H2ogfLH7D0QkNVCdDsVYPdOf0prUi14HepeIuASAdaO2JbWq
pYMCe+7WIyP4hITFZ+GZj580Fxg35B8j+WBvrK9fy6nZRgKnCs5igPTbCI/Xgb39
19y364bzPL8LVQGKFP9cy1dVE0kEkC5JhfmTk5mSCGW0MxT1siObxqB+0SM2bBPe
3kEcmyDfDjflKNYXUxhGNrER31aoCetjlg1mpm3hWYOHhrcF9+W8GPtokgKxjaWx
9NlL96TbbXNtcmFf3JKWfm8zGOw7EXFKLDBLBfc02b6DJJv53FD71rzkMfPBLFwg
Vwk1A0ngpFdC9viMnSYReFLKd9psaYKZPiml2LUkvhZS15x3YYMSKglQcmN7y1TO
jyGaLWh8B374GetXZWoB83eDjvoKAo7u5yZtj0BpAL1y/kyDiQSAG93F/Gg3iV1k
S85LRz4ajdd+afo7tJFMceo11zAPXaeSGooZs6VkeKVlGN+LMRlT2mCZgfWQuaa1
tLI8RdHe8m4+NDD0H8jfTNlMmNRUm1qb0uuPi4dF083OpGEkZcNCTxw4bkyEhrfG
IEeI2pn4nFY4Aj4Hpszjqgpr6TZrxnoC4Nc9HHGvhhEXcGpudX6MTkBwF+TD3ifq
B9bS5UTn50WdBXiJq1VfXGPSK5wRnS+gBrEtxme3FEUZx39rTNx27uVZZozYgT85
IJEIbF3g1wQojfvHDk42fnNBMM2FYJDGe9qDVre2Jb0eWKG5Il5Oq8SkQ2Kz5umZ
003kn6FoB7LZPfrtdkYUgoQ0R4qefujEODnJeidHyD9AZlvwCuy7Yn2bX+vMvofn
hThRKr6yeFPUccV62yIdlyUw34hF3hU/sV7gfpXOsrz35nkkunFCr8xrpZ0vv1wP
w2tY6fsA99yyUHmeFV5QDjA+cewIQjGukR31Hks41qLfH5B89oQq/Jny3RNo8C//
336vCLlkyt1/mzLdWe8xcHo+Mzmyv0khM47IFsstrZijgMhdrDa+N5OsmKhBenzI
HTqLLh0kmo3c0of2fT4pqq3GV/HHXFel6N5dZb05uMZvnrlQk5O1B2w11B53slTo
RlVUSv3D5DkiGCP8jMGrOji9IaEwPinNxBe2md8ZaZpuT3ih6yd1+ft89c1+u+kl
vI5wBdiTWECcarh91HO0GmVceEyge0LKy3TwkRi4kkqGqkgiuJ1NVmaRYvldTt3/
0bUS4N9Mla41+r+VlhtJn2cxcw1t0kH4eKuUucbDyfNtRHpdk2wUjl2yAAw/qYPw
UPbeOBIxor5dVxqWr7lEe6AUWTDcieumTvK0c3RZKdtBpQ95yzy/rDNttMS9AQLh
DBFiUcLz+xm8y/v5+oVQlBrnizyIeWmVfi/nRwh8il7uS4AJ71/FSdQrcmVnbfdg
kEAvpCFfr+wLZ+Cw8Mmi+Votw9NdFLNAgFEwwElHtYm6CHj0CqN2v+G+w3ahsMNK
wMaXkmNU9yTtKzmnxBukMRVp6T8NGsdVswvLC1vLIFfgmUK9GOBx3GBhvBnw7w5D
pQwtJAqUgiPKJ6E1ULkvbB87Cpzu5+OqRYsynyjUEAR+FeWaSF69fVeLORpxipZ9
WwxbxqKCk9agU7H3rCSQ/PWwledzcbXKdYq0lYSW++yq5DkIUXc6S2ZpzJtLyYp5
HX6V3YtGjB6DHnpfjYnVi7qSTGVqXUuhghh5Hmn5SXWNCzpTg+pSOVQSFn2fjOvO
dXqNyjftPMxdm8l5GVOsFSsuykpc7jdLTOfgtB6u3XGt+WnOCn6QvfEO86pCLLrp
ZuM56SOjlFJvGqx9cL3VIgNGtsAXNGff22V1OV7M+zosmPpTCMsIxXvuvhQXya2q
7qBT4usk/RsSebEBw3pRJjJWPfntCCe+rYb53KOxPJin8UGXsQTdeqAuuEQKxQtd
It0yhTB+XxVdsB+A8+y1batCeXoqD6jk+U2BanZ/aAy1hoUaVKPhx1xNWV3CpxOh
v8tkWrrJLEku1oNEv0AGDml1jiZVYBS1DDB3PYTF/FPmovWc/3KyA8fbBVLtZ9gd
G9d9g4Tl7SJ/6U9R2nUgHHfS1g6AIIC9TuNruGbrJEu7ajj392gWmYxtLHn1+Gyg
YIUMTMEKaNk4boUNi0qfjVr5+yVtJ57Da0e05uHNp6DnXIHYh8KlxSIsce132k7N
qWBnY5Il4oifK6xOf5np3PrS0JVAPBphRbtNuNXBiK26UhEGxdULomtcOiSMrv6H
YLsmbG1KcZvKmvUnVYefrJQ+khtv+cgG8GjGFglFIDLPLiSE7O+1wABq7CRC5B9Q
+XPj4WjfEXAc8QSmNe0NoVDwsqYjyEgVaIlEdBFAY9srFLxLRg5/VyA2gbkSz/2k
qexY9G8yTcuHOsTZMgyXSaoYg3oKNBgXI0GwSGdEAoJNm1tYwEjZOzFRfT29PMZn
EPAnG1dLf8B2lzSSVvhqDSGMclk/iXkvbOur0J19bjwIaXUd/Qfv9Ysxwa6P5gmv
J3vcMMMrOSA0KzPz50ARq9LUqRaHbxLtyLiXCJkcz1rAxuAemSc9VjCzMOq+cn2H
aZ+ZmeNgnD4On83VTzlQThRhEWJ/aRxLg+tCqLugRGVmYTQ/grb77QKvTxxnWo9J
v5Md6tJxHFOglQh2DBo+W/6arLnM+ABMuyAGzJV2MVdXo0RmUVdEMEbIBDwQSCj4
8GczT+yscJoW44zlnyg9iR9aFolcVU8G3yHTAy+UpPir6kiVEfKO8Gy/7zDOuTew
BJs/LCivWlHvNA5e6VXLjsTQPwA7wJtKSOqhQlRF7zQgSFtlIOzuazidWty/KNq3
ApwQt9xkcnEhzK9iigXOfLyZwdAmniTZgExUZihw2YwTCPW4w/BC9C55KkO4R6dZ
0ZYBcBmVkStlE89IEJN8394LImmSv3ThOoyxHa/VpsKgh/mfbWkjKDYPwM9q7+OX
JKrwc2SduPSTXOl2IzMr9L7p+2SflkNoX3/nLBwYJT/waRc6JE08a++tE9DhAczo
v8OwcWtFxFS60zp9hzuiilGvK8t4r6pk4/0KkyhxR96iEYb/m+xa3ZHBkX0Thmwn
AZxraOHd1qluZ9jCsV69Oq2/aTztBEQBef99+V0I7H7TqSr9AY38kcmhC7sQM1/I
Ok/z8JO0SCzm36GPDr2xOJrY7usjFmK6Cmhl2IhNIpgxtqVAxdXLqGzGJWCZlFUC
kwYcTjF4sYdO+14f4DMiSseTYKhnbKxeEwvRsSyl4J+T0Gv5qZPmMGoZOeMS+dAy
Ij13u/dMeMIozzXthhJY5UK/WiG0FxJw3y4/P3C/Im6P048tbPxNFIMkDqq9uOAN
WlQDJfGUyT5ZNxLQIn1ytTdM8lcH8KXqaRek7FQmuolfyExcBpQwYmLrZh4E444r
9AATbPGyBvhLHwpswmyEBMvl/610VXFovjs7fGtenF1LRquHld865+rw6hiIEi04
ucOPCvAZRUUHliKJlWZp3N8V22yMdtT0QhZQa8VlCO4TeZ2Eyd6RaArqA6vCl5Xj
oTKBuDz9lkDmKZjvYX2CcaZoE/N1Wy+OUXnDGDDSwfOwtL+PNF9jWsiZfR4MS+Gd
60+rMz+gcmnidusIpZtyjp93fZVaw/o6zDXXDGoIfWTfxUVgC71pqJuCNSrsW7bP
s4bRaTBI1y4fDmks11gQUnx/At0OuqXj7fJLFilQ0xL3voN4QYyHk/jzXy+GceK4
1ggAqDlkEsd584+kTUId14AisU0tKGKEX8WJHoYqsJBszSN/ldXuSJ4X4KndGtLF
t2vbiiLCU6ViUbnTHiu6iQ/tbdiVMXKAYvCfT3dqENUtrYJTRyovjj7DRVd2QMPo
ps0yqNarnzjhxIE8PIh1MWZFXqPD2Jbro+zSjO0d7rQg/Vrve3L99Ng3H5+CEc+V
Ha8hkKQ4ohY4GLtdh/N4Vr76XFgF9UmjDhe8F29vY0ZaTeMSuIXYTgh7uz09D5h1
gf34ObykseMNw8gokr96l/5kilS1O5DtIKpeL8ULhU0DU4XansdD/DibDjBMvfUh
ZQrbZOrWHa/BceNiMYfpBXDJdXB0HMw1B8ctDElseu8NW0vJ5Z5FGmn048hV486X
cswLD+2X0CIi6CuxpzCOfJOijfCnRIxk4cRbDJm/Kek1G3WR1ykfYXcjQYTbJn2j
HiLfzDO0zQyL6tAQxowbahdg1hdLB3e/YCx313pj6xMBhdPsPu9A9I++PcjU1i0P
A/VX1ff4E3SCthSJ2vS9a0MA3JIk/ZzmiSTlZlVqUT82/B4Mq3qam/eMxGHUV1cG
ecZT8lruoEt3quXMxRuX5FaN7chDnh/luO49eScv9EZA6dY85jK5MIElsqmjQTtA
g9z5w32LYt2ltkJGrYDiSQp5uVhdXRYe4eviKxnKy/0kPhBVfeUfNl4k6F2Fwbic
zr3E1AODMOG6d+o7Ta+oRCgpv9Lsg6NeEKZRCa2vRL3ZEWVtFTiAJHNSfIRvtj4p
bVdNpSeMBjThi5f5/XacYW+Q4R9zybSkUH4glr/ZuJ3P1GxCeajhwLg5HgYK+dFy
emsKYHhaKbxG9HrfAEZwb+WjceP0fBldvUdgoCMpbTFQ7f6+vm0uXusqkVoKqWYh
zAVkeMcG1xsrms7U8hqMgMCo8V2/g5nahCCmo1zTvly4uSbLPa7pMSjtNdES8F04
FStyCnvpUd+dtNrhgW0XrxK9uh0LegCKBu+k1MLWbkuW9dwGsi9tjunhkm04ZC5+
iPqdQV76r2JYwuI0bIVzsOoQxkmLtFOQf0VEbTcsHL0EQy8q9tfsv45ZfAbDEkVN
M4CjgA7UN+UfUq4wDcpHnWMP1kY/Vxl8J2jVyQmCwSIbPC+VjvTdwSiaRrnDRb78
HMoid7bVqw6TmdEg63V3LrsGP6gzEZPIsNcx5lB7/iqftIWeWTqJv7AnHrLsZ/v9
Jhg3gJ008cCsbO77TNPlWQyGA74O3MwGVunBn5OLZcRmGQYP4nlzEqcu75Xe/6qz
MquF2iiwkXG3zbC6DzhTmWEJsAVai6+CzeBMfXmeMG28IjkRIXmikMNQF2NHMc2f
qtrfZTp1vbbV3NaUN9EaVX6Je8Z+N9f/g3my3XhxRA6r9+UqmHUNp+wzRMFtDpYf
Q5sOZunIYZH1KeDZCZPJxQ7okQdDVbwlAmnIrNvY9CCbDPpAQ6hfdlRCGJOHNBYE
wkHEhWW8DlSwovO+JNfRXCxh8mAeoO1TlbC9C4fIbfJoNEOxmGT/Ynw5aN8qODmX
9vXfUHdo3Mdyn7TV7x8oyqshFWOyiNGvEGI/sVVCgxDOijmeVzg9ycsMdUuBlXSU
PLy5FLeiAYn9NC3UmfbH39OvPLN5CTCHR3lmtQ6DP4bQoigHf1sWVxZabLQvyFGT
VlglBEB8P7JQXWf9NhJYYy9xiIqIv0km+0cqTIpWkAhfDKYe09c1+D1aecEbQICD
IYzk686C9XDRx4eplxBYHGGkwr4ydgozEtu1DcAkbyx2dkJ7q9psXZ7xygV1nYLm
jPVNgkALR2TXdbJTCIZ5gOmEia6KuN2MXVYhfN0hM9/HstYp5kYpOLydD1zaiDg+
HZInYwEuxzUm1wCYPiIk1EoY8+jJX7N66CZkBFWh2tN4CFOdgJO6263+YXdrWMH0
sR+dFWBg8ifhwX5PwP8JP60dmYBA5ms0WWLqO5u5baQ90ZO1r+Iflg6OZbQDfbCr
+rnz6Y8ujSX+rX3TPJ6lC8ucB5Wlgphw/ftSDkb1iPW3c9iUA2sn+Pi/4gNI+9Hv
LAM8VE+5cgwcfORLuJ3bjIQEnrEGThU7OSQbPPHQLxI9AAm/Hw0yH73r1Lv3bfCP
risrrIoj32zx/OXxDGmatYuVje/PM/uNANskytpxWjndEuEre5/jvhXJRsmAr/a6
BbK3l5ZkmppQ2c5zYUSpPU9YYW6djrMYZFF22BXmjen3Cpn7lcKerxWX3Wko32iv
0YS83t20/wux5u9YI3DAcoFSEvB34lZ4/BC6SotN1LyrctB1itVWxjqSAyy08UJ4
rJIqpX4z5CmCbAcW5WgU/adsUU8l5ZmLVViQO1KlYpfrrOHHl5iBmyobEYP+H8PX
VZK44OdpCnkBc+n5U/HXDEJJVrqEPuKUSKGS9atbCE28XCkG+UWEu6/UOGeon/gR
SA0MfibhwLMZq5o/7rg+LgDWj8NqadEiNKfqKzHP3XkbZb8Yf1GzGzBV8yxzehy7
rLaVyxUiIXOO1DPA9KCxfLetuhlaHScG66t0IICQFS8X9hbFQRe0qa4UJitXWN7m
PGHD0GVf9QbQFSu7V4kUdfKhFVr3VhgJOkNpwfk9LqK67/Q9L2yabMUlvsClxNEi
L5jDjnVjwMM00YaqWzXiEEx2Q0n7xJjzB2uWUUtKBRxw7L+t6gopwNqil4y7Uzvy
NBr8fua+s6wp3V06Pl/NjPCyzs9zyt4uZCI4HR2LOCbVmMD6BRdrCFDw0Q6tUQ0C
6JG/l06Ee7kRpd8ynsJI1NC18du63M04gXBP4dhjkGZQ9eYsYgklPEELRNYMmbzl
Yzr1MRXv9x67auNxIg2fiTe+rNKr67XITyqNzq6qet+5svqfYhu7ncUNQAiklKSv
EK939cqmXnY0wUTUsxCql0CSqF16jJbFg+sE4Oc9TwPyvlWWssG6FJJ1bdotiyZO
puEcKYIQXf5zxZ0tOTExDicdDzI+1L81B+lsnN9OX4iZ+ouZkiPR7ezg9PN0VD6U
bIUu1v+1q1oaDJyj+JkOs59NxTJSzHqiUSgT/YcAdm7a3VFyqXmVuZNpOkPN0o1M
qhAdlwjVIkVoo2KnjKCH8fSbFWHEXcNtr15RkiF1zwuKsKgNilG0Tt6KToBNp9F5
/xR0V1Vadrc5lP0WYhOFea7lx9zVdBaJkPlBeuKFVD7uFjm+Ol+mrWQBYvou1fzg
iI4spCVvWFlS57tfTBmlr0UspVg2/h/9OnjS3/j07eFBNeXSXb2/tH+tgM5Cf0bt
YUNrq1kt3/Eflrjnt3bOjBJA7QyCVsR5SHZxb47pVbTxxcToCBr7w42EOlrrIL0d
HfY5tfRXekUmt8Uo+LRdI8pgVuGVuup99XqN5MnD0q1JlSS1C74LUNHf7pk26Id9
yp+t8yxVXyF6Vb7HSb62xr/bl0IU6KTJ4reaJijicOIgDtsxiaZ/oK24EC+9VExz
aYD4DRR/DJZ1SGAt2wGBFIk+/onwY+bO3BIOx/Hv4NzpNtYg83YtaJV+/7afB1yu
6ksuQst55x631uNwViHCNDvwp1uLFcQdiGlE3WZL/ZRRnXbOQUEFJJuxuyqGm6mT
Q1nYBJrf/MrH+efjxXpHMhyNRqLOEwEXKxuJF87BdQ5C6SygB4djPVB0I/4jFyMO
D0dqX/Pbz9OpJpzN0KzwmuT3GJzgta7PlWwav+yAeOiCJ7eBYq/QieZoSFF8w78u
Im/9YCW1F7lMGX/lCCRhVLGznARgl4hKh76RHCB56IhvFj8OBdAnhYt/04LkkDSw
Ig775cI4K5cNAu+Xv8DuhbKSrZi0CqAyBD2TgwFXTZxxJTbhG9YKdSiYOpwnMglT
TmCaxC5YFl6Ry/ISvRKBa+qk2b+KbfQNvwpaNgH2xGvG7cpiUQGiuUpxBlKuE0Vs
tf/7vdYmWukXGZrUPJEQuAWYGQd/Ltz8hebpke4yJq61yESv9jZXwIhvHCJDFntQ
6klPaTEuc0SeZvQbviuaa5Hj3NwqLzL8atBRfsCkaKdT36XhQCSz5uR9ukoj8CAM
akzVOy/RR4YOTfCk9wcyhvRLoF5qXSQIPyd/7qrx7++1eXLPf/zld6Oh/DILqPYg
mttV229mzLGmh3up5b44Gox+ODyoksvK7pn05T6pZ329Q5RSgGtwyfG5L8iEzTHN
WyPZZruZMyi5EM+BktD/63Ld8wPR/eo7vmtYhcOdSz33XyIEIlUob/bzAvSTXHh6
T41bMT7+Ry4jbFuShgilwzxnIjRX3dhrd+BvaO6Q8wD1fot0i6c6lmRMQbZmQE/l
yhF44QKzWdZXLGKQach44l2NtEhAuvFJJdvjL6xp9odE8hSBD6Bgpu3e0MxUtDGw
ImgMflSFP7sJyv9bu3AMs3wJiRJOGcYCS96T5n5CL0JqL1J9JhjuwTVf1DeWwwWp
JVA5TWFDwgN3IxfwJh4qOlRXqE2qii7Rc7SAKx1+/UMbq6k1HuSHofsFSKgdBCcD
8vTUWjd8UPNlvIhNE4hVtenG9v7mEYxmA3lOqkOkX+f/Dspa35NSgzgM9TInp1nl
43DCnHC5J9fgdw9AB18+qsl05laWtzZMyxTH/PHsIelEH5CQX1wIxKXbXlSOWnjC
W+Td7i/XvLDgASx1DZGcqlWLnzitOEO2ppVclZzX3HnH2awXny40G90mlMj0iHW/
tw3Wp+JNRwptoRIeB9TMF4BoG2dmxfmsddG5YqS89KkKj2B9NmdMXAWAnE4yRx32
wfb7aaH55vI9z3oB2szSbaOWapI4youEI5wONBBHGdqoxJC88lueaHMKHGo4AoI7
Breyl51WA+4fygP3goGYOxRVTUDMQ1uMgqOoOfxj2dQODAr5r1Ff5W1q9w3EXTL7
QCVI3KOYCuUXe+m9BZXFLINWVQbmltUj1yEJZk4qWtTTkgpAi0mrWfeaLpVLHQIU
9NYTLukFN7IsSu/kx9TSjWvS8FzwtFXd7GDmHe5I1ZOdFlWJxTm5UpmTuHVuDXuN
w3z7sxCwIIguVE1A9pwRabPBfeziF3R/YG6uTT0Rnx7laaMcKLQRfYeYH/vm6ld3
hknMIqD5p+s5BYhnXN7HBtywKdNul16ldBULWxrNQ36tNf2h8Q/3/ntZ3OGcoaSs
+D99QWALqtCPAuDmGZ/363OIKVJxQK0GHJRNxSKj2Lyxta+8Ydqgo53X4YDMJaLs
eOo9Y/GFuvOeegND7iimLsdWhlm+6oXoQOv06EMMyuYmRJONQj10+fIps4dJ5DOq
grkKihKB8XRhkkCBXyT2k5L4G7JGZbhTkIbc4oi+WGexidGxbtLpivPYVqJLLcKe
nkxGcWhrYAtmua7lKLcxVvDVrHo9Jls33BdY9lnbvIlyPfCYoFASRcz+3I9THlcb
HHI5xiLiAAeJWHJyNH1sk1kRrKdWc55WUPXSvN3vtqxwpW8dMNSXPHc7s40LdFNm
fuNPUauqvFiLeCBhYuN4E1/hb8LFnRixaWKVtNt9a0aFbMT01U3L+0IkZjkF9OzL
9h2aPicVf8LxLKRRgdk5xNNl0p9pYematmajlvKhy/L2BTSTWZFHI6lMi3MChEB4
F4Ymo/eZKLc08s2MId7pC4RgkvfSVoKEs6tY7vbP3g2kJnvBsUSYFWccGyvCbSfE
LkDqnnb6kuCtwu3rTri3gJuG7Hu9ThmMX1qI+wsIyQMfd/71MHqqZGKoLbcgHseK
gYEGI1Zu9TmYZWyBCscLdbqW1jD5Kzdom2Za67ULqunTDTpfsbWH3AgEVcjZiK/h
MYa9SYhymh4ECTqPmcV9H4rh1+HHdTqhWiQZ7hm2QuvgJZ+aAgPhOHQvU8uTsG/I
mAiloaOX1FO4WUYp1/6YNXsE4nOgix/fcUeErcMKpmuOOOI7m/iZchkpHnGBy0/c
moADGGgBpldlF7whmvAuws1yjzCPfqcozytAQPrjYmazCNPV7U9tBF3/Yy85XB7L
L4IBom44J2+P0rkQ12WfFKWfn9P5M9VXjdhq+g0N5HhTxMDWjuE+FCM3+11MKbCY
g3ZpjtzpPVKIVsSzsNTuRXmZ7z1atOjN4Fd6C3ytLZOlVzAIN4koeb0CGYj/nUnF
px6pw/TsURiNHr9fi3qHBvaB0M4DFU5NdibbXSCQrvbCdZtiZGonFbNXFqog7Alf
DUXJjkum5qUj2ijRS7+daS/kDFMCxvf8Vu65dw9QZmFIWjfbQtaX9s4aNCCp0Dn+
kwkLf7stNk51gZXTzQV8RkvlShRdQ+3UpXz7Yw+BZAEc/5Ahn+IgXdFCt0WR1OKq
HIqTeMxxzynurp/oBEORNwYclPkmFIfjBl4T5J0ELxR8wI+Xcjj6OVmATJOmIOz+
UTFrckrnbeZ7I6U60D7tWfo1GADPbVkLURXIQvAo+a9k5QzUmsYe3tkGC8cV3luW
Zh+hgjL7wvCL2m8Wxf+9wb+PdrWDaiUvCxuaLz5oFoxSTijpe9KvHqoDJboaT4LR
PqvLm9rMKZ8sW1NLjfgPBCJqXeVJGccX+yBZ6dR9gKk0hI0astTt40llqq8qewIr
Y41pYeooQU/NB74j1qlByD5sYC644eV0NYdMPmamobzP22ujJcqXZe+Ema5vvdM9
UEA3ftS+ANFJ4SshXVRxJfa7cx15JYlrT6kBtzMyq45qhbK/ZBk0aZY4KF6h0Iln
64xZcXGIkoyhoW55zivdxMjz022HUiVAxKXcClzvJf4vaKJqKlfLIrrWUbHJo/UZ
9G6CPANX55vs5FrNJ+H3zClcxbrYiEPDmBQpe22/FdN21lsnvxG4rGtSy7lb3KwQ
7K6QhOYpML/GPP0M3MYw2GHXEEw+JbrLrCbHkFw1np2U+e3Zde6zuUAPyZFdyNtv
kvG2AcZ/zmqatG0yZ/BJklLDBA6j/R2LQ2s5h9wK9LLyyqRJBQbHSvXkRkQOIAMW
/hmuxK7dilKZaeG2/SdyG2pWTGQsdpAGBErzJSGg6YaroghCHbRGie1AUs+GCOsg
4y9EIaBuxJG7M6jngX7QnEVv3kgKGgli1I8i7dDHGgPDLg5w5izFigngDbuf2XA0
J9ZI7kQh7ulC3Dqhh9q4WtSwvoeFk0M94RaWqZakzCenRcSaLm3zJddMkkGMqogN
APhAfZP+jfMRofOp3IyZ4/T5Y6u9bgSfJdwHhD4fYXEw5urHGwcmrvr0yFewrwfa
MQ2UdKfwgudIlJNBC7QWVrm3CrUUKkDpT5ewhfizElhcddZFZ5+sJeAH+4R5/UVH
DfiprTRi2AQWZBOcInoX0t0nhGZX/0QPpBaaemy9h59EXQNCHwUxOoc3xmRDDJl8
iriBI/TagU5MA/KRk+PKJWlCLplCot/T8nsaJCiiCaXACWZe+lW/ypa1uZx6QYlX
Mn2MLlVnNx/QT5zVS/RtZm69B1FfCrfob+wH4Qk+U785dRVCflYOWN265Ok7hXG3
GqEgev1UCmkdiDV/6AmIb1mrn5uwNeTmSAEeleIAtX2VwyJ3NC6fx3W5wMAqfye/
AArtPsnbTAalS2/gjl6Vcb36F+J/njQNq+noSCYca4VREQmIln/iENazc10P5ZPm
4/kekuPLmcn7MyTO1h67RH+LAvz/CuudxdLDKPsju8qGQc14/IVgu8W0fDsYS6WE
YhvyTlkg1V4BpGzg1wUj0Pbll270dGS75z+KzTh4BWRxFfqBzpWWf0Uw+R8lW3sS
IuEg2k/PRfrjyXB8GzdhoMWP5+s61KdOm6ac5beuWqrgf7rKdzNkUcs5M/VX1x1Q
XrBmiUbi3bxIlD8MTbSinyW02MKv1qaSB/DOIpWZ/B8XmKSuyLa8QiYOVkTRRAXp
MI9eqwkUJRYww+2z2KM0PtfKBirr2mYVtRW45sCvzbsncY2A6GLdUOjgiUMM9HiI
g9qDbFQEq0WDe2xh5DTyO6mkdWBDwjRYb+jUh7Z2XwMs7IxwBl1cMCHIEWix1D1G
8s+StyOSeDXVeUNvB7ss/2Z2XkAt8bM/mHc2t1FuRFmy9hCYngKjuQMtgr6Ig0zU
KtwXjEYjL1z+iadsGCXPsBL6fsdY0s5eUjXVKjOSCfgXuLLlx3T/7DB5PLviLQP8
YNtnWyCLAArQspcUR7WxNPPBOzzXSPpggoRwR7sVPtPgoC2/ghTfIOflNSRoTqB1
Q2HBFFdun8hrERgDiVLAd/qSSy706TxqEQciVtR/0Ekut6bs3+5VC0ZBcd0x5FEG
QjRQIMdoP4syoNvqRPN/CCTkCozimxFLEYR1AqdjmZjglY8RSAxkhUQ7qHeizC6N
Pt6dHdN384l5NpAy17oVqfRgwoeC1owYDE2vLzn7PUz1GXI4BP+miT3XahfRKrDe
3Bag1qsb+ZR3xnegH9hJjAh6yc8jB3nVqsRwBO4JL4+vJrA5H1ugq9t3YDTFXL+E
af2YIU37Zja4SyV7a+bilTJTHblaxTjOVIDUna8iZQtUGKuOZH9EwuIjM5mscXbR
+3OZDbcW3yc4PjmwL0ySOQuTf0AMKMDe2wtoLYCSOyNLgFtlqC0ttPhMedigTKwW
aNtjgqwJvFBNv9d7GhKI5e8QHWzSGB5DDrJSD+PPrsa0Xdf3j7rCNI4PQsU5gdjZ
RJC6S7iy0/UjKb5y1OSbD8sBLtNZ0A/ChD8Q58mBK3j4mR92SbPj+V2sRW+CgjBR
cv2FKSVco2ZNvPGq6Ll4brTTc6T0QEFFD656JgYM1uD2nojIW/XPFRVj/8wIXYnu
TC3hdTc/c5dWnKv5s/22kN5NqdjyixCv1C+NnMabtY2BHiGuwBoiYtleYHM0PqBf
/3nL70FxgHd+U7gFNIZooIVSniRRs8dARctKozrw3Q+HANlIBbYpQ0dRAYu0kqoW
9hql38gRmLvfFOVCcR5E0f0QNQWpUUn1LAyAM9uigLsmEg38CwSu1UgCjwm61MRk
YFCa1la+HrabivHgie58b5jvChoQEqmvK68FzJSzX3f3mspTid5Zk/JvmLHbQSZN
6TxNLtdKXvqplsy5Jp3aNmOmCiC8oKTfc2YOz6q/95vhyHXyy/HuekWHBYCQNaZj
VmYE9KKMir59XMeiuz/l0Vu1Mj5e4qX8qr3TtX06daNKJb3vNVPrX2grKfKpmcoi
fA5qptYcwscYBxVQ6RAPHANQVDV4kdv0FDzAOgsK+AmpAWyDiuj5bKOFpu+MvI/X
k44Cc/v/DmAg9ptFCTHdrLMFKDYMOvlj7/CqQwJveN7n8dLgTA3tQ+g1twpMpz84
jHjDVROegE1aQ+JHws20j+GR1F+/E6KGhOJ8Od0ETYoOH8gzmZCB5obRL46eaicJ
BahcFbdwpJyw8BA77bIF/1faB/Y51IQzjL2Ml12GKWqVbvpMxdA/S43o9NH8Xt13
Vdkho7AXrJ2MgPosf83VixM3EelTUGu/txGKXE1CiWDPgH183jS1OyNRASGRG/xm
B0CtGYMeYlUmxsH6uBmLcfH85my+s30jvAElfj95ledH48AUxMXv6zj9w4/JXbHl
rdTgLDj2wNKvOhpSIm4N9bp5AGKHPMDKWHKLLmOeylqLG7sHCELpDiz+TB+XNnlE
7tmWxKfRICuMvhISaPW8vGmHmVRCEDjhFzx4bnYy9TU5In0/jq18M5QJDfynhI61
RCPsxi/zWhmQzBpBSFGXey+VIfD/eDqy14VpIgJWpUKsCPZvNPCiQEekNDDgwSj6
VCnUFRZD0kkxGytrFPknA1hAAKgZkHg48JTWr0F0g8wf54QZ5bfu/9Z6RVSKNWsY
iOv7HEV3tf22MPvM02yQdN1zspIykKUFbsjRAni6c5+kyylNjBY9BucwZ2Kv3J4z
yNvc4rHTnfVgoJlwZEy2zrNltnzrE6h9Tw2Wut/ngIt7qOGUb0q0JtPqLZPsUnlQ
0nQFPwTVIzwCZn9jMDDEjX3QcEYCbgBgWQSxcrvt6q+qYNU/0UlbMm9UIhBFPmIr
AjnDvq8m4VE/MS47NAI+6r5y5p6H2Us2RA5TQZKrZ46SWSdGtPG4qyj8mXsA8L+8
UMEXfq0dCfeSibO1oKYs0Fhs2HafgC4XJujwATxNjDqYNkyLvj5uv/SVmG6LwSOp
VdSFWhtK0o0wRd55g2wz68O94zWYLOKnUWPXo6NjY39KyhWoTb6w7IhlSsUFZHzQ
jvQG8Tupm1aNZpFf8mp6CStGz/mG7cok+ZBMJhtRkyPryWfxiMPftzhZgcC0T3io
FZXNw6RhxcCwPwLbU2u3RlMLj5PV8M9oiFa7U/Z0L14H4Pxs4TMqHzXdmdN73I3W
IFdlhEMa2tH533Cn+GNt0uKdYea/WtCzbtk1ys6CnnijuXZNp2Gkei6hrMRBspnt
Lwo4A4hF4she4nUirgJw77ELHt+qRyR4usgUF5p8cubOlE+FWY2sXhvN4Fh5UhTX
VopmTDRiNfKl3wODldI0dzPVwgZfA/rUrZS4dNNJ2LN+lzeBnuNR8bhfUHR6+ayX
m1I8rIDyEllhHtvlHzjKnD8XVWe7u4PxwpU1LOwGFTGggzP/7ox/XL5+W63wsIaY
ssGlmDtzLmlDZKqlV4I0gyPEYMqHw8UQqGu2Igx+i4L0fIncDqYINP9feQ9R1/lv
1O3njuozLNPtkWuL6089BJqQC4LGmooxGieCRl9/Uq6UR/QrPGbrULNI+66na/HQ
h3tWAVVdpKBRwIvTL8HyIiSzBvf07H+/POcu8u4HOTgmWTXFuV+PmP+OHbggsIeQ
5N81jKVETkpbQROop/0Ba5xdp8YxG7EBqXDKJ6JUKJwS+o7bs+XLiAylgx4qu7cU
f53+lrbtYRaGeGsaW515X9g9DwaG71//cKa4c7RXoxYTZ+8DCvS65aMuMRPKwVvc
lr7gBiwyYtgr22HqRyEI2+Axs6ydcciDUym1XA+zQq1gBXr1KJsG6s/puLr0C8he
uXYJ3veWsZ65hQDsBZSnXxFnijtwpL4vwgkaKzEbrN81yq3+YrFYQ5uDKPJzQjan
vpr1mNT1RsVyvjNcUz83w3BVj5JKOZPXFdy7AsAG6lnE0YITukkkTM+HGkh5DkET
bNRlKPmpMzzg5Oy6Rc+NF/BR3T9OKlAe+R4LjRkUKE/SI0mPi0JNdjj7bdV6bOdx
39WimGlyAbAQH5W5PtCrZQjVAsTZbMbXO6okTf5ON5/M/iQ0uVkEuOyaRZa6+ys9
5PQ8S2Xr14KH1BwRVsswQuKM/ZJaNXu9/4GFTk3EUoH61QiIitPnmzd9COaxtWxT
TFjZV526Z0GD0byNoDftavcgPDbPL3R85P1cqri8dEVBZ2cWXOmJ2LYeZ2JaGPVy
kf/v3jXCKzpLnysdMD8oj6Ovo/TwpPZdaAIhzbKnxaDxwOhfKUTHc48xHb72Dkve
I7R3uwkbYH9oCiI1IVnq05brb7uLik7MYDJxOwb2mao8kltOIG/PqLqzj5tPy56l
wdpAVNla+vmjqnbRBwP8bv91BHhjqSV4BTF3+8otLEI9CVQ14YaJHsFg82zqUQwa
jCMHXitZUgvxdUmEtAhtttOXdSWusFpQ7OfQzIMoF2rqLNfVDXD0oNroheyb7A7t
Hlk6xCLpz68xQSPp8Qg7hmTQBYsg+t2SeaSi+ZwB/d6edkgT6BPQ/Y6rCX7nXIUx
H7BMtL86XEGsK6v2519bDpqA+rXCvbEAgE+MIPwQkK2mBm6wUj0RdvfLdRBHW+sv
8u6PCFpnbtTEtrbWrN1zpu0YGqz2g8v2Fex6qd2l4tY+j41gA3QZ8xM/BPthruxT
FIbcjvgWcPnNEtBgzvUlk/hcD04bymARjaU+VIPjUKmRvJkHY8XAEXaCXyz4ApuJ
82c+cbbQqluCCCKx+LgtHeeCYaHvqFxtNeViqxsTLIX1idhPu2zTqhEf8ChYsXve
YEDq83mXxSwXpayBJ1v5kv4nnIwFyQcRpqcpzV0W9i7fNoGKKLcILwg/rd6W7fty
xa8KrfpDY6yVs1xZTIcyiiCNx5ZSmAbO3cACwuYJfbWDevRVckF0XlyWnYYJ2eXn
QvuVVnUnHeUyQMsZv1PzZgrhLuh1iQ390T0+CGvcfXpRzbEzrVqA/GBIHqrZnbdJ
B4/VwXcIjlPjrXGY/hsawVefcxp2GlDJccP+/1Gk8ubQC9Rx3KFCoV+Y7+mk9P/h
9MOoPAgCOWYs5WI85ijcLQJodIXzKZLOKcY/0nlFQrj4jBqcTs8eK4cEEH4qsbDi
Knbx8e6k8GLlG2Cnj9QkgWkx5slP4BKusAAuIUznI7DK6Jehx5hUnud+lI2mSeHv
0z8FLqx348ogU+NUiBshR7TSigApXc920K0bCwtBOlAePdqammeqtqnBPVf/xMAg
5/DmcDKyO0dV5Qit8Eo6m0rqV6nZEykMKOCLbeL1sKOAOlBStSa+Hs7QYGDl4iUI
+jCS9bgn7LhiNVBHTbkCCBO12n2+TdLAtEy1P11ArRaYJ+idjAYuLOrBrE3unSf0
V01by1NxLvim7vr28+k9KOIWptkQVNpKRBVHKxrzUV5dKaEgv1O9NWkBqcPDMLuO
8Q2/73ORmBSiAepk+MTM4rKpltraRCKlLxpSJe9sy+m/V4URkPigroO9FUKwkdTQ
sWFXJb4oZpRecCiKJk/hEiEpG1fAYkuQj2flhj2pF2i1GK1YoVItuyy6/JapUepB
09J89SWBXmtnbbjfnxtOWEf3ubFvaQxL2VB1jtYOycxo4SZgYCsCNRsKfu8+ufPl
g7AUCrk876Y1iZMdIUjNKL0Zmlx0FicPPd1HfKiFCzgjFG4Jw9L3DkFhMA+TDApf
S6kJt601WG8XZBWLemeUaq/7t0+bucbL4tRrorYrJ1LOfxjgz5Dl9OV8KlL7goPk
4NirYUsKVtjIbFNLToreUrV/ujMBRY7VrVr4+aXHbZZLEA5gYmOHyNP3vuaN8PD8
pXnAEGbRZd9l+uBK2jXRoOCQZ4YVE4wv6wTL+jSSmBMFqI5O2Hpo15ZXD0SzahiQ
TWx9sZqeeg6YLGPwXYORixt9j7qH+kI/fwiTWsPt2IUHI3o4R1zvIWfH2yBnV/OU
ahp09akq98BkNJvc4L1DDZmPIvpfFdBEXIxDQQtD5aMXsqBGnOPnq5g3Y92NKv8Q
4tq/ELlxyjmXngGPIwK7rWSt2AxJv3wOqkCWCsRt7EhhQbyLGWtowC1vye1m3+ff
T0tdixkR0XMIQGqEtumRtx4rK+DL5KZBTqLZV8WMVfWP0wrJRxcHF2jj47HRJX46
/GUb4eRsPemm5TVtHuX8YWkZXPJGM+1s6TVLwoItwLBBgwtiF17HVKEJkh0LL50z
YXDoibvUqOLdiohIDYPaDvFh28/2sRSHRVYOJfy/rXSFdjh83Es09XKpedEcEfge
wqvd0FB+5rAu+AWxhxygXUy70u5/mV83O4smEE5SPQDQGqKcQQbmRF1zVzSbLzOB
Jlny92SohscRCdgeOamCZmd8dMORKaW2frA9ADPU4xn+NkO1GGCJW1Sb9euloKfv
cDRCV2ADtsizjFbaTBIO1IB+OFWBhuDOf0pmvBhM8FlTunzHcUdCxPEYwdXo+PNl
B4ugE7Y4X5vIEZ4oCh7t+laFLf/aRN6dhScNeshUaH2aj2Ldq1zZFHnSM4I5YLQX
RM/3kZpiT5N5vHDKXZCFTDuJGKaEwPeDd9GrAHQqRGucz7KFqcdciOdM9Su9NwAS
PmiCePNRx8IPE7DocjhAQIZkWPWYWxCtSWQjf2Bf/14bj9wmb9h3Z2RgBwzJmvkW
A4Sp2mDu2Wc8rPd/HLfGczSvkvibtmTP1xzVkWIo0i2ID8juK1ZuXBl7SZylcZ7F
bCCEDC49R3PsV5cggjj+bebeUi8cO7tgTRGbX/7kBre8q9XRB1NIX2sFYiNWPW/9
5vX5jG6Sk8mfauJ3ERGY57ZkArus01Xg1QWWGudK0F/a+BB+Yn04bmDpjTMqTXYi
azhPo2ErxFP+SZK2ydM3dgs/W/Ja6IODJREOPcXSLJm4LCZ6r3OBTDZE5N8u296j
tesfqDnECk+X3lD0Om0b2ptCG4nXBHH5rjtgPu1vyIuuQPxkQD69Lh8DSaqOCn6E
BQSETH5nhJg81P5NXvbwQg9xAG2UpxLo6QIHEOZ8MstZNlLQed54QrGlSUS07rmO
3v7M66IXkpyEtfhnWGfEa0+iORd27bz/plk0MjRUCrI6l2f1BIX4rPrVumAs1JHl
d7g6qxKciZS0+riO8lDiMLb/Cj4TbNPK9SVbpazsQ4wymEaiDf/33qI2olxgsDG+
CIMRnbqTIrbBJrksuT47Ic3zkW+7yDU8D8PgIyiM9P1X0aK8mRZcXjxjOQw0MLXv
fS+QKbw+AFzM/xHxBi/EWslWLb+3YPrs7rH7Pdrn/gC8M9fRln8PKZTY9I9V0FRO
MhiXL57xze34QlK2CyvIclwiBiKR3aVG3bDv5Ww0C5SRnBRBaOCf0U/Seo7P1cDW
RIReGeu1M+1HXrbwUL5MxBNeqVLd7x1fn0kwB99nblqAUNYqWNg4q/W129e+24Sp
GfkPBj2UTNK5WCG/50LSWWtlkF7Q+SPJAMnsIkpdvx9bpTL0/7rHpIxhYP+jlhNM
GvjM1UEqZPKPSmpJ/diCaRxgR2ssG2EOYJgYThKhbidGLX33Az87EjovaPfDzWZF
BrbhstpRbJUcgYQ4zobSupHlRFnx1BQE6BIa9XY2iXbbsfEC81aT9eEIfSxhHKd1
pylK9TUazurM3AnROnOYxNaZJwWxaiTLHfPOmlZFJfkgLsucjZRer0xAvXjkMk3i
idWfDblbeTs8fDeMMpqXyaBc4m1PGJi1K5qb2BU2ugZd3H1NM95U/ZUaHIGobn/2
MO9FmZDTbSk/H8F15BC4cLdWMhnu9WlW5jPT2yWPnXcF7Gwxs8aWUi1b85AgrdnX
z0fc7jWlBqnM/gurQKVZUdtbWZz/NK7izhNY5V0xhmyCBQt9wSRt4Ot5nEZb93oJ
okSXRbBCjtT6UXGQS5ND/TwR3iRvG/5DLHlZ4VLEbivWXY+YMtx8/aOBqRqdmqJg
ayxz0SjeYBX5muvP2BX02VkXNH/cuiv8gMeP5bqsVcYUkvG1a5oo3yltyK7PWEp/
GSjk+q7O/SjNPtqzoK8e0yj46AyCXTAyoj2Qei9UwnxexG9k4ncDFG1yHBiuW1KD
DVhhVy5EoXU7x36FPDlCrShjHVegGM5Vjhd6xO1vha/tAfqnX2YIFlw47RJb3z6e
p7UhWfP5EVWkGC4dL7vVWoUe2E2PTxiTnFrDadLAfsmyHj5YPXXuA5WWlfl0j0xC
JVXBYMv2I9wckPHesWaNfDfdZJCVtlWEMCltU9SHWFX+ZDLeEyAOUHo9cQzyShD5
t4+YNH2VJjtPPqR7QLd8bGtvSRL3w5SwAhKTyJyREr5h88wzkfS45euDmVdeoFV1
0d3xSF6pfQ1l54GXoheZktD6gA+hYtXPqEC2IhN5SMfmbDrKXZFgz7Ndz6yBjL+Q
6sgYgD7TfIOfcVSUofFiTdH1bRBeprrfv21OX1+QS29PAdXYdXEEPprG6Jf1BVXZ
PAnI0EJzuap8679/+GcmJCIT177Jm7IC3eP4EqrQX4v2Lgh9FavHTMX+kwfKIJ6y
jGgMqJNkr7nolzAaijYSYiKn70hx8P+yu9G9t3atdg21nOHhMZFBf/paPiCTb9aq
rUf0T7qoSNIK53jKSV9G/ZsLfRVvshAC8fVh7QGg3WQPMwgFuWvT4Jm/sTHKg3IM
meJKtYweLeHBjdrDCIYQNly1DUU6/SOv9YMHuySq5IV0hDhUR8nzwLdYsOLc8HU/
wFenhGMDyFj3/ZrbOnIPE3tdr+E7jnenGYswf5MKK9I/jT05qucrBnas0VR9BDrH
KkxLY/kYrNVwYydPyax/2AbaTjolJOCPa+zfHTweNLzYMGcuKNaAj0Oo7YO0tcpR
w5WOhFsnSy6LgpL+fSFh2ihL6onJyW0Wg3vffLFDL8Dx0pm5SFZ5mh2pGIc2JcGu
/yvUcfEUM1CFry/wQ5zkjslWuXVXplGPe0eTUZ6fgP45U/5hggcat1XFtU8wXGD1
KVnJ5wDR/0DNLzYGdTWp2x9gVOxZ4/uLYiC7mQVNbO3Z+C4thuM1R2f46rz2wucM
kZyf76jKCtMTJSCWK1XqtRbtd8xNfsj4D1XIPaMdXIuZ++ZL4vtoDIzZPhI6MWQb
MhFwdqeQ/zo9xKztHXj1dA72hLrJaFu5J+GhE/KLn/0cyIRCsa2d+q+k/g1iZIsB
Y65PB4O3C6yo6gWD0rb44u3PMyS7SxB+30D8a75QNwwbzcPf64LnHjVYv2vr02VT
jaJ9nuJz43VhGmC3F2eWrTRM48J/imQtPE59Cczs+H+VFCrg16HHVd7CUBTiIbg6
CQMxAvPLtfNDkEc/a/+5SFMdUHb4DKdoflpYUw4qrmsQ7cmcvWccPSr/WkGSkItF
iofN76Dnwb5yPP0gtCuNtgCHUd2RVD6V1aiD2en5gf9eCw3TP97+Zq0bmrpaZxfO
wQdwRa3S2Z3HlNUvYSAL3sIw3ZMVo/KVizJURqZdSJOso64a2puTBYRNI/hCVqV6
Z9Q0fCorTswDEfInJ3kcjOe3sWE7w4a5+nE6sLVuqz4mJfSrcNiur5HrmqjDIaAF
SgdvBYukLwlzu7w1OxJYnilY0XdvgHXYpjrurBM+K7rdnGb+WlMlu52cuUhM9EMA
ouart43l8Lqq5HFonp/lcWT9rXpLTcykcaLMPZKb3KGLxGxdRA4iL+YBjqq1DAyF
NKK/+j6xD6hAKZcGAWaOC4ad009a8FG0NWFl3YiaZUkU8yuFK6yZ8Y8bsIp8MfnD
jXbC6OGyhb0LS5xKbe1p7GML2ffxhW3O6FDNWy9wzdEjCOYsnBxQkySslDRNH20X
EF9fwGVqRDEo1EaE15NstKhct/zJOt4afrIZp0/8aUiPL7qkBhzmn+gcULgVMzd4
WTLGYuv5S628PQ07zKRh4dLHORyqhftX14i15WNOZLksJNFQ9buEekoLmQmQKrCr
pxfnmtxJiy8Twh02zpf6KQglA1POSogoULfBrsJvYi4gZUMA7onDLXmAw0j6JDtQ
JbLMjJK6+g9xHCF1887UJHUnSlmdCEz39yq7UlMP3My7a/1NCQ/bjAx4bnfoRpQn
bacwPtY7C1xxeWXbMPNlrQtPOIsWLM22DY8JEHa/4ySgOX4ZCmiOPzaffpUXDhnh
oEWn0h9OEA4n8OJY5Oc1jrFZl9+QU+kqbY879DrZhvXcuxQQWdPW+hXSivhoTJsC
urlK+SGTE2fm5ntzdrv3DXcquJ5D7v+38SS8kIL0cEx2Nas4dYjXrTkLhGtvP54Z
ok0l9+R1DSfK7iJlchDJ6n8oXp6C4YhDmNdfyZkwuHg1HRgVaYbCLiAy53uib6YF
AgKoH56f0LoQlGJRnS0AY3jR1xoJebZUgTn0pa6T+U4gcvqGN4rmbYYiRr3X8oM8
xQiDYSAyIGs5jbiZiM/W4b2LiwShqCNYIQtapO8W0YqI1r1UIJdNjQwZ6qIr+wzE
0tcVAcbmbBFWPJqirx3U6gxlpYGcsqLPh1KgfaU/VW2tl19so7wxTAgHzqafgLh8
ComD0fbkHn9RstuFKVbro0paop2FbrO1gA/Fx4uT0798s9V3Ao6e6pvdRowJhk2c
WojDyTg0VQ7OBtgiXYWF5YLk1OCvmBL5uZGVpLzazWYaE2Jta03i01NrHfYh8p0k
3GvlbJE3l9psLlElXPacB4FH8EOax/TMuOdhBlGLjck6EZavdImopcwtE6czZvUI
a9aPV8qSlRCEPFUAR9kcRf+/9YRaVP94TxohCHV9ibszxwln3yDTG/tcVBIcTVuD
4gD19OcSucetHVm1gZ8+QAY46gP76rOmc+mBZ7OFtbiSc9rym7Rd/uR2DPLjMjuE
V31RXDcdXStM4ziLAMvZ3ACglSsF1lm6MpY2tB0esDp6kZKXUA3DwxZpFkZbWYgm
5nCNxffsrT6nMwT8kznzb92/xSdoBtthAMmtj9+gm6pIWlO7IdDmky8fbZ9ZNkd8
4L94x39fX0o/ovkjcS6THHkTLIFNiOQ0DZjzwdovoE2S3+l+AnJ61d1QFsz7IMPu
ADhb0J7pOukzg6ZeMo3dDMDFvZ5D4tDK5k6KueoV3GZO6QDsWIgCmfyhmIv9gHzr
W8Fwy4L7XfPMjb9WOZt5VkwCmXG8oq3a6dWqluTz19w+Ta0HEtUj0E8C3nMUEDWr
txJ0H8CVXeAfNaxbJabvr8f3TBC2p6BZLXRBawn1wgnqxalCHF1Dh3S3V0Qg0ulP
C36uKSfZqkaFoVJ/EvLTD3HVY6Jf2OwKUNXco+3ScBZP5WmeX//sYPpUJZd4QFc+
uWvxAg6lpZV/EWZ8sDBx5y9CPSeT5LhqDeCilqSWeZLgHhbBSmuv1HxTuZrVnAIw
6YunCSBD/gxkaniDVlfnVy2ERDnEYF6sDXXcQPuBrC7/6io/cHvUri/SAcxBNvQa
+3RyxWylTqXL3Kw2VSFWdx4Ge9Y08RxQ1B4Z76a80TG9hjhugSzRbDrkRJkpl6qs
3AC9jA3/i179JhAoYd7CKzNAsSemIBGlF6gVHSXDHRqaJQ6JBgM7E2iOzL8h7Ci0
zsg5mCw4BT7v4qqEUPmeqYZyRncLKeN1y6Yl8c1tD5jfOELv+oppsvKganexncmC
wKN8ZtCUJES4YlzsvO8g4iFCDzCVterTpClR9+JSvfDoFLs5uDdmx4+5biU/XQus
1kc9YAKuooin1RL3fZFHbAuNELeY7DCZL1h/sfz/vdCNpT5/ogIf1mGQLXm1TBvp
rN+1heZn4e5bajI5MpiJxEFdZMuTHK2XInnbIkWoj4CBExV+XfvWNEvint/xAFBw
mtFFyhHpomAUutky8bDN1JzTlGCMFRq2so0g6F2tJq+inAoZRdQ7jq+AOgKvmHUE
QPVKM9yS5Ay7W3dsVR4aqiEuL+5KXJkh9IJqmvImSJ8hLVVzzFqks6uHSFzxLhlD
mJ9e/8YVSBgHvKvttWGAGeMoGSyVPPeyi4iu7iNyqEHD0Q5zfbTAKPWOQe6SZoW1
/tdtLz6s5n4TQ5ng00ckZ0QZhGbmM0mz3qPA3KHsw8uqnPqWfdBiZ7e/WfiKuBBt
E30k2xiF1cDYeiKMJ9ZxaWiv2AOR2GK2z+8yv8hQcjjILGxieGwZXqX99DWkfpN8
hbyo+W3QTjteTo+ld8rKG/vzlxG36h/kMwoSXO/btzI7Nwtcasb/Eoia5ZnyLE3O
9QLIik53lALKX9MpsfQgND1EEYjJDp3JKpIYbHhyl6x1LU9oe0BfHfxinqJdin79
JcPYlZ31ptA37oGJnELCJU3NEqbAMwjMUX7LrjfWV6E4ylbVpp5vMNX7zb2QzLtM
XbtM2TWrwk80tlXomit9QJ9fFN+Mi1dpd92zE1S7jkcUPjx3mGCZSmetWP6RGQKV
J9QQFc8dQfhDZgGj37JqnkqUq1NYdJVPmHhi36J/1Ub7yROhLE7YtkQaN5tvGoyf
3mfVDv0O/sLvFWtYoqD/aCQS+Ghge9K/4+97AOHAbGhb9XKKHFOE+02WskwyBMDK
/f5Emqe9cS5yf40fvgZADXVhioE02+9k0Fj/uiEvor7T77Od3J56K/ji+6mc4z8U
2wdkgzeHXtMuf1JI5sjyAodZ+Nvs4BRUzZ2oSwupeDS9KaI97E/dpGmJJIvVvdok
lCsGyFgchCcQRyvrqzYKE6g4ypj0fc6hMbizfjntaR5/a3J2/+ZHDOGe03leDbkS
GJ/0xhNao0T5En6t9E8eNnkvkzooV1NI90hACkTRgFDzlxh+veo8ghipsM9rWOrT
kddl65Y/4/OEISk8TLQQWFW51s+c4itTGtdsH5fj0ipIi+daekLmpHbOL5aOyYyk
T4cNg10xX4WgNFM6C2RHhIN5/AYYLGeVomxVBRiw/P5N72sDi+aHjNAlNMrLfqDl
pbd27rIWgMHk8pB+9mBDel5YgUvzKjX7BeP7YMTB2DZB+SDlxTJNU2v9S4tbTQvp
94fatoeqNjyK6pUphrGSGaFSFMBI+GG/AKI9+0LA9vgvPZHCXgLkjy8V9tHmLdtc
vqOjWXHN8wsDWYjEK6bnZ7Hn+2Ut6NVQwvAHnG2Bvu6ADiiZaU87c8NkgYrdpy9Y
tIX0M1jeMipcM2K7DvAdgNHCZWFLt+iNb/27lcbWUffiRIDthTN3V/7T1sUmgoHN
/TV8uJxKM/Dd2zdWDVVPVzTLFk2HrFJjr0c/gZGG3llpZ9uz2GNfLN9F7nUCHz0i
b9Fpgu+C3gQeF7GvnfSdtKMghUIpfUXSCLXmhLjKzzqaLdcq+aam7hlDBReUp7Ml
G7x9UQXsq9W7wc5cnk3e7iXXOxLTQQIwwCmQbQ63fteWA4fgtQDFdVBWSVI5VYE9
W1q8Q8DsEzsty/yiMDRz0YiYGAcHgsLW/GbXKsCCs3mR2xbUbp949GJFwhCb3jz9
IjVQqftq7SfG35ZT//E2BhVvsEnvsgfrb05gXM0InWM1T1aK76W5xA8iZQMP0NBu
2OjqsUk9cpOmeIB5wXH8RPUAnfwlpYisHirWpgUIvE5GoKwPEM2Oc9o8guuSJilA
30fShDAxE6pnaXS2mrmyE1lqq7HhHoBp/p2Qf+22nrusj98M4HQGf7MJWb+0xFJz
afXaUZ2XAhf4+dfiHX7TSHcRdiuwokBTFrPhd3rYN6d+eSJ7RaOcxn6TTZechsfg
mufBgP325zVCkP08jnzFkLp9kxA0cZHyZoBm2VrM0lLnwIkryynnxADqGn1o+nwQ
F4xWE1kF2DOnt3zd1P2o9jG2ipEjR5onqX4FwMoC/LlAmA25866WeOEs8uUXlizh
RpR8Xz7XniW5qX0Agkka1bp3/l1ukHFerN+6GyhBkY9d5+paKrndtPHItgyXRP2u
Afegj2Ew9vyPdL+GCA14r3FKKR5ME8qsbQEsh3M654JDqPWKJnK6Eu5WjQ39/aON
YzbHNPR1oGmQWbgaUw6bE5xbEZWA4B+BbJy3pRnpmO1F0kxYGUNc4GcJ7NV3mcEM
KP1XnL40zk9EvraSQzAQyFVQxkwL8DsqDewOaU/wr7xEQOYcSj1lJFw47MZwX5PU
vzWa41/S+BL+SyKKELyBr647JPrLMjuHlO2bYpttR8OyLnc732K4fqtNrA9+nV+I
qgkrssaCsLbWQGurPOGmuNVtqgynitKBsUnGD8GWS7yH+0nLO+D+anGgr4hhmTuV
SOWapj0zJKuQvK7WX2PgH1XiWNezq2a9OymeFYFwIBV0MZuvfSWdCvtfUX1JcnWJ
40VfrQqCt3JGF/CbH6Tb94XEC7cBXFRFcHrLBYZ3jpbgWBLXuNoBPPbB/U1GV0mk
CKh2gaygpA+sxt5KWYfvynfoRa5aPKWqZiR7oS8l9cnIuBd3DU7TN93+ci6UM+06
YKs/jzGEsXm60RPCzOOMEHGwePqv01n6IRMwi8z5mkBfM/bwtTeEcZxNhlYPrayw
yzqQpXwczhN+jsY//EWCtgfumjMESpGc565WUNlsvVSB7ZuCpoM+wATZIPPtj8wX
i7ioXpBcMdTLNN6Apl8m+L2JWrCH5WxeCKrZA8fzRgxwTv5g0SgPJoisGrPRQolP
8YRdgIQQ0Ajlka0rsfs+3J/f9HthppZ4Oj6cknI5CfXs/relVJ1xBZ0vgpYBUDV7
9LpmGxx8bTi3WDiZPCRK8Z3n+QGJxMud9UWp9G5pkX/4iTBmFwvnpfpVFdEcCNaJ
TJ+1ihVHloHG7CmI28pJ7HcEyrfN6QfNrMErjUDroUN8cGAV0CV9Ru3ohUB69nqs
7E5/WbBZ2irhnq4JUR3kgJe9Atzeplf30NXktUVdmg8Ef0t70SB99W3Pxrp9pu2Z
KacZ/dwFwCToECizhbY7cNp2t+2LlMW0gwgScfczrO3MUCZNpi0yQdNwUS+utljT
aWbwDCXV1QU3DB5PygDRtYdZno8pdYcZYNhwnOAwnQi9F0398kcdvfr1KZrTLgO9
XY9YQCsSq6oB8AvK9xSWZcGW/N24hWltAG40TEwPp0O75+Ot4GXqxKnHJpc9C/qo
tqsHMsvKJf182tK/84EPfQzfy6Pt9Cd/cwkSBbb6dBGjszT422xiCWwlcR6r94Ij
DZ07uCu9oac2RNcFjOsQzoU/giTSm3cF6EZNJ3s/ZVLTwAg4HZBNy84eXWdQvYz0
/Q7rX01TSghXEEnZIxWt4y8vTciYgOAoeMeqwj03NMHU9kZLSkfQDzINeR6Hb28x
pEQftIalse0XUYqJj4MlsvjeDDKqaGYY9ibTQL5SUGVVpttU1BXzGKsCnjyQNWl2
Hp5ZfrF5+gPmZuXdlqwP6D8PYN6TaF98GWAK/Eag7dpyNpTuDdSatN4iGYiWPyYd
cHKVHfjxQtrVvSVJuDAg4vzZT1mfvMLu2tCsN1vdYj6yrai9KL3NbRwwcgJBEdpw
Bw62pXsBfI/4XKJyBIVwbx53eBwPNYtMrzbYwC/e1I8J+BpnU4+nsjGZvKnXFpp+
1gkIWV97yd1tzOpCS59EJ4TMOBa9SeNEVdrqbuDHOdK7Z6TGuxx6WueC8Bf++cVP
2YhhvGCrB5Cz8t7CMItBsVykWPLbus54QkWk+ub2YX9HXPB59+JnCfA/GznEvaEd
zde5sUqupDyTJiR2IaN79NkENcl7gFsXu+m07yHwEbQMR8n8TNd1bIwY5csA4stL
B9plTeYBik2yYALgcsGrTF59Nv9Z5acASUy7CiybiQ/8Z3CSQGQqPAaTxQzym8BH
Jk2p3BoKivCXr38Th62AZ7eORsnL6ndXjpsm4vcXIIZN9SjMfeeYUKpGZ7Zlf3Bm
8YPnnpEs6QKvvhMI/9VLQAaLHnQM6N5Jt2WP3WdH5VpBRMUI5xvq2GkIQq3xKuAv
upLt3xai0EyEeLiYBXr6ETXv2K88mMZtbfC4yUqSvN5j14f1t2Z7H+JpGqWK/1pe
Tb3hSR8dPBpwwh4rKZNelAuca5i17aighRfnS2AH8OCGNUgIbUUrov2fpb5SJu5J
YjkQvnlT9Hk9OeuzBWfY1wAjTK5YvCW5q5hCIgV+aGEP6A/MsZ6HK/zXjkw9IySl
HNNYFhKocJ/X82qTyYRN18MvKjxwDvFTZ+rBtkRuflQV7Sah1C7YwEr+sRnOB4W9
JOrR0AuUutobV28FDs1XDv33Si4DvNBANPal6B2IshjfeC4p9MdqkFQEK2w2i86B
HMBfH0DGpVagEHFwh9oCXWXuX3aBqInVltMnq+pkP8XQwNWHxtAMzPJB1rM9zOBs
5eei9zXI48vK8dmqKjxGpbJDhHTFOP8EjCMb0Tn6T8TqGGN4JP1pGNV1CpEr0M3n
8POp0K9++avnRXWUXk2DzWwcMI52RIRFkiKFXJe6vA04uftlg1qf13oVL3JJx8ob
83xt74D5I16Ej2cEA+/D78nYnde1c0dMKrs82NhDcrHg+k1pvWlP1GqH4g+4J3yE
PRGupugKw/kpqwN+AQ8JLsK2AvH0ZPdyfXI8sBwlvRe8bDyQMg3yHAUe/vy5Bb82
DDKBCCz1Qbf4dMjVc/bj7C41JBG7snEcTY6dzV5xBSeP/zfpqFrhQzRBBidQtZuQ
woFhbTpvb2k6l4poEFOcdqypvOmYl630hCuDf1U2FWISmqM1OvDEvw7FKYu9vSfk
4tkUUX31dJSa7ZnqTQkFLw4jmFvLeISMB52GGmRpye6OkGC6QF9Xu4XjX9VZOTqu
kzJ73x4Qb6zek3KYEyYz+jDTiBxc+DTCrD9s7prFfmqHI+yfzMlpIUgzCHZ/ZHdB
N66PxFMmRrzZPGicn42tHGI3L0HXpFbgYEDiUNQ7DXteiEjFYfWBPCriw3DYZvaw
XS+wZUGxXWXXVOI7p2HWUCax3rFI0ZE+B4xKaFPzF7r2pq61JnBsq9BKj7Ns5HoQ
VnmfBRLcsPnKUvylLLVHwvNjyOsOYLi5kwsL9qEaphLFwyGbU8Bv9gi+/L+W/CJx
WrdbAr/Ph+QWBznuFMUg/8+TTZodo87mM/uQG6Aq6dwFjzLpVNZQQChfPFnHIfcO
PCgyp+nCQj3A0hqBcBxKadIaQRgXnC+tIWczw48s0JRCLVpl6bGv8XQMNpZRxePi
yTmCP5hElp9zg4142FNQX9gTjTzViJdRAAJjo8DZDUUCZfD9M5CSMYHWvLfbIe8P
9ioq1NM1YKImkhD3Euam+gIoJtgclsffNrkSRFhvXw7yyvhTOpHcpEFAdCZeMy4j
6p+d+jLfvz9SWsEI6oNMiehzMTDGPSD0mU46gspnqw90wkPmJw7DXdormVXWWrcC
j21kqlBvrsiKMSwaAo6KfpjxmK6FfHT6GY7ok7hKe4eAZ+zVkU4kDl7hmxu91hZR
n20QZ0PFbSljbFS2xsls7v7ctfPpMhZ8sl0zitn+sUQ5qIKi8Wu978szCrx24afB
d/BqGTZ27SmeARZ2SVqwKNYFH2j7OKmuz/49rCVg/tH3B53C1HM2wB99EKx36SA9
EjHLQPeymupVTubSEwWcETUX5rXad17BLxuxqe2vIRcbSIIzePArPdoukxHp729O
leM42Mkplw5cnGPdZc+742sYuRZdeokdGffW+uXEp3Ki4RZminbwENDNl6kimkC9
0Hm9hsr/Dh3bYXfDsFgL/3tTsnxeG8xVeErVKQeMciRmJ8DJAhtGZjcgAuJlBt6P
RnpF5nh2Ssxv9a4xw4XAgm6eT7UL39+l4s8GW1SkK3k1xx3LhK9CqogIzGLruIEw
Z7o69zCgPfFQHowKPCu//PBnM/DsmB8TCmVvekeAwPJHxy+AfORzmxkU2JYExHe0
UUAFiwlB4dw2HtfDoH7upuTHC2J8N1UwyGQK0cmN2C/SBr9xVWM41HW/HohhPSCU
LaRpFGhx8MGZXLeYZF/VJRJP6zvI1mPPE48/iP5zSOdev0lpm2NxavnGK3RTs+u2
wTOkPItKHarVyMAYJiGQwwN+lN6vLUzsDrxstmvDzq/Khsk98o4rclJZD0s59wkd
lusS7FOpYWYhvZAwftdAcaF5gdl84X3NSDOo3en6AxUoDT9OKuySEn2X5/xHMRCO
QezZ/ANqYj4KcwKeMHvGOHtEOPgEstSxCzSZ9rGvEbwxmVd1kFybwE8wVWxogwX0
bFArML//2NIVonfqmVYwBV7xsJcozp/JlQdevItQgXi0Mrj+543ZkxPNJrFITyZw
2eMQMv5FfYR0vCY2wCwT8+qDK4/idoYkisVnK1JxiKQdkE5L4dnesqtJ60BEVXLl
Lff4Mq1yZ4tJqChH87UNicSbsp5zm2KV1g3SzMYLp+SBa4Tda8iA0CTpsTUcIruM
MbJyxZceQ3iCKPysPZOIKarhB6NTuX4jMRFggD9BUirzGVc6SNPAc3n9NSF7Q1YR
79T0LPm2+niRXqUM8taQY2TbQANYKAY9FkxDnv5Yfk9SOyZSKxzDkaKXx/deFQJW
Cmnbvgnv8/cPKObJ9YWAysY06GgQGJ/K54bg0Qk2O/swBDYdzoewvhk4WZht2+fX
O3khq9Y4a5LMPSR/IByYZYC9QXiFMMtFWPdSaJClTyPbuBJgOGJJWlM85M1mpT0B
M1tCUzRjb7qB3AQEs3blG61j2D1O8h+ST1qNCICQwXBHrfzDxq7tbZOIwVBwFU3r
WY0cze2g9uGfGDQnrCKEjndika3LI94HmtFLNI2oEZ8WzN/BGOAIegZzDqrsQGoI
pKN3jHvg+xwNhR6epOmEWBM2+VJ0irty+BIjmHeGEkF3MDz9fevqJrWNlbbmaBiY
vZGwkMDVUvwjrzEokXAtBaNG/zdoouPEMqlL5wNfJMiDC+TqkhaSGNl2Ye0EJvN0
v8X3jBFtKcivewiGrRc2n6llYVZHIzL9A4VO9Ti/8ofkerxvEMaMH6AeNLEogcT6
7sAhZwT2pbiY0OCRu3WAzbbZgWW2l7sHRq3vWc3S50fZZl3143gk/OBhbm6Ld1LF
/DGhoTpVFtLlHz2bB5MXKYVx94GgDiB026KdPx0CmlK4RV0NNv8mH89EY6s2KSwN
VdHC9iOvZjtkXtKBB0U9+Y0N1S/pe4pIOgX0A5JRMwxshLIF2RSEdc1Nz/468MUy
a1OYd76Snb6zHLwMs4sXMkD1ebSEEt0MJh1aakWoGcnt9ZERuLvm2OU97GLQT3Z4
i2yMdf5iQ3oInPAmneo/ND95xwcUaU49oQOgsTqboWus5nJt9bJhokstOxfgG48K
LeqZOwiVjKOoVy1JDoUGhiH9l5Pi/WpkupvB3SbCjTvU73hFwdky9NSUMFtpGRCX
YzgjNG+whk6+P2SDbRLsv0+4aYr09r5aKcPHJtzfLI97QrzC0Ik5dVd7+9Buq4G4
4URk+8mgrotSaNUTvth+8PWQiPjsXLm/miSbeK0yqUCoQvF+pfhLFWNy9IhJztTH
tblgQjVAZeBTI/OjLk+TWk80qSugaCcr4RAd3C+qaRgR4VeQEle714AVbTKnOPE/
WGUtMmq8SD4fVsNzsOF2/Hv6ko75T8D2tNU+jhdkf2X/dA1Y7bfNA684UJbcDNLB
rhikn609ooU/cemFqPTHp38ZGEnAAM8PsioqLtUfl+VkcRwLTLBehGXPuG0G14sj
4ZRiRNxwGVqiv4l+Mgd4khdgKHcxDd2MfR0yYms2v5+Hy1+rTZtAKHjOK1SXBdiN
43kD4zBZB8BbpbnGN+lIxKnsbmpvsIgKywdSqRUcEc42nvZjdAOPZI0NtO6/+Gbp
CM8kSJTYRXD1UqkrMboRDlYNVv3AeprFk0KALonsboFvJ+kTMjFW1c5B0ulHUdDK
u9bup2LLkXObsLgfL8Da5FXeqtrODt5aR6sTxFeN+9kzSdiD4VQfglYkohQJmg6Q
riwMTUvDzQWLkjQM6oL+tKQzUUlZ1TYc2XsnSwRN8Yy2Mc1+F/fAuHCvfCUJkEk7
h4Ktt7lQALkd3uRJcduayNzm5pmDauLUPZwynk5Z9Jrob5paoLiUAJnoPwoGHWwl
esJzlj64lU0dSTYnWfOcFJ2vPTxyBGni/UEQLutnH0QprLb7v5oCZ/pLo4P/YFU7
8wTFwREv/MdWxRUgFjuH6JPVBoHn5HOZn4PW18mdrqHyUKRQrkipCrDvVuuyf4SG
d/P3hrbdgMhlXZgITXebv0cGs1gWss5iKALw30ULZAys0PdT6IqhfBTEiCAg/NYy
MrKbU1WVwJnv2Md1hSx8xU98Tk8FsSEofX+dxDqOzNEztELX16l+zZ0ZAjkW8mMn
C+R50SkKG+Rwkl+mn8LoZxy8E26k/PgqgWGWZWl3BjUXpgAy+gSuesmFlJD/lJsj
MiNQZG+hiZMKwPsV6X+/a8lJ/N4+nY3BB+V0KmOlilk59jE3Vh2fwE/a6ksrG0P8
1813GX6con2wTCzWP2v6+umV/mN1nOVEVvJFF1vRTM2cPR521s45wOY+AtqDGgRH
gYMcmsyghBJd8FncQ27rX3aGWNbbGifidejrWOgHeRflVhTkz3HYOBT+RQRg3mHV
grFU9X0IZW9b9DFAguEkxmVKF/MoYZfjjPH+AYwdRhWpVTFjHjSXGUhDvi9vLeuD
Rpm3Xbr29PEcb+BvwOomF+BtVtMSKCnTFIDEFjcQAaAJV70E4iFBKni3hd3/iYUG
u4bK0X/OWbBWjLSdPYgD0/NZ8GCZuNTz+fMGFiuZL1AGpoOgpIpM0w64StGp8evS
y4hXwQvIjbKfruOibKXE4K0U7dPEFHZ/vk8nFOS8o4MAtstf8SSbHeUa9wTMUBZ4
3hW+sYWIUyPd9a8GWkF7zaEKTygHq5PSht63JYOeE6N8eaMaUf16BA7b1auV2Nx2
+MP9LrxR2W5r4tDCeUpFnYyI2PdK2ZoAqLVW6QUaZQ/5Fnuf7P0ylS43Mr3Xqx8k
tPZZUMdroG+p4hoP6jyeg07bkFEZa5OibbVJGbMgPz+iv4nD76zSiyzsv3UolHcL
v7KsqvoyXAiNkK0fRFyJFz1JgVNg7KBk09y1IiM9wftE5r+EChApnxxFGXeSA84Q
JmYUVBii9N8EnFdgCtjdTcuerqw1d8kjtMBoqSj8UAkSHbodNkT03zFIH1Ap+VAH
ANODKDR+AE3Lw1XpawByn0j+bpWaXCqJ2FE1B0ibu+zXlteNZD+9Of66zPA6NDkZ
8mGjTJgMh0PAmzJMUmjn7UyIRgOizGYy5iY9HnLpCIfOGspZsmPzpbF47RsV5UA+
oOaxjvHvT81qm8+QM/Fh0Sx2dfLIK3bkbHTUMSm6BmCrkn3N3SspmOs9Wh4MJy4X
WkGRP4U56PonnM4XWxJgpfc4i0Vkp2YidNMHeUzBXVxrCqKExWcJrgkCfMGnln0q
/WG+SriVQ9B3GmryGS/Uxb0RRW8ZutSEvCSbOzQe+AfRvUp80F2MiBIY7ZkHjWRE
kAbd0dsL+8qVczT9XdY2FX8yDPeCMz6XZmOaJL6Z8w/ww5fAGv0maWR7wRNIQgsx
I+fW3uAiOu+V28Cgg3DuBc05Z7v0A9vb7P1QhyxtCdzIRVtyy8g0iCXB1pbgLaEW
UsuLoikrCcMCFbiiAjXyHYQQbXic3kO8qvkAm95PUFk08r9M4sCL1oz7U3O8bvhe
W2s5H4StHwSD5JjMxgry4l5SeVf0dRtgUQIsOmBDzg3ioRszNJKrNSRhzPpkswHl
prVISox87UFPTS9sIER8GzCdFfup3+x3T0Eg6YScZ37N9ALbklF1IDYKC/SBQLI9
MoEmxeK7c4aHKCxoHKs22GEYD688bTWBZYSXDse38ZaYfNir4SzxwHqjYNyzkI8L
8MaLHvsTmhHIh7q7JhLTua096keSh5QLsfi62l2Z9vGjsM2Mm1H7N3QLcTXvBfAu
Plca6Rx3+gTBxno3QitoCp2dvNQm7WJOtX62gh3AfmzxZxd92G9ib0TepbPKzVOo
7bjRTW13u3jK+Zbzp/vqIGRUKoEkw4fylHCdxLSf/T2mHXtbEhb4n1pIPuh+PzTY
BXkL2F4EkDvdlvt3x7sw9gvDTUE0s1X7GrSU3YBUx3bWqvF/uh4rddvKpM+Z15E+
0p/nRd3XllAPqNP9xbP0cstPIMulBuPv7MgOgkQkErXSkvDXhqkyKG5esRUJWfDC
lPcKRmzd35p2lH+neoBEdOcxg5WwvvGe2ylrTpT9kiZrPdsG8HMZpLTIpJwM/LOj
SQPu18VtGLl2m1sGPXoIxDzG4n+iKRJTPPKt/RIDMnBPKQaWAW4tWW7vwv6x+TAn
61gp+5wlTkcnXOlXBS5/NgE7Y60fzMd5/SDF6iQ5vG9LmSd117300ypCnuYTJShJ
bvTOENnwgcDieDU/Mn1s8tY43ocVOlZcT9DuKbX5yempLf9n8TDDtZ6h96LUo7Wh
nj4gOglmLl+YAVTjCXB+XcYuqQB4vxanIpPgxMr/tADHcU8L0vISPISkBvPSv5SH
cDCE4jtqF5W+bvypVzDmTb8pAayh/uhuDKjR+MAu4Uieq2d2EB+31wEHlED+3DvP
NcaJUr3Sk3S6dlbFlCzFpjYCN1Hs1J8D6L+jV73+CVNMc8h2FumLa0QUkkXfu/OQ
dqwX0nEpo/zbPxinqtOlxl0AinxRcidbB1Ctc5PM4vsmwHAaSo75Mq9J8iRm6XSQ
lJFW9E7FLe0E7VZv9EgVwA/Yp7WorNC6pvEUNQVW9xv/yGX9AiL436D/1yQknCWA
KwSfSonn9huK9Xug+JD86jW5iSEnRLhmyHA5K53wT3G7hADyN3s1AYmah600H6hQ
iatrTuIHF9TbSWRNaaK9XAcG/a5YF5UofatxO/dYduZChf9FcN+Nc08Qq7XAybXe
9zAaYgRQm2mUvAB7QD49Z7MOztP+QMNbkSuajWDNC6YVxQq692bRNTxV3V2mu9Qj
vK2zGaCzLxnpr0T/Y/3d8YUSdyxJqnXuaU7ZuDmP4X87H7JviP1Bv3aYBe3V6mTj
HpnrZgLY5moM37BRYajiUIYwXR/evGAxq4qJ+0g3wePMDj5JaJnkfFQ2r3oVpofU
xGMJfSMDgeyn0yIrlHZUfE6Q2Cw1LPaEjtKNEt2o1eCBVKZk9zpt1bV/KIXHlzvo
ZpHn/pqDbCXxE7hQdk36BhQ/oUHwXbQbx2pJzvH9ok0VahRlbxdkC9e8OQRCkuDV
ZtXqxW45a3CEO6AN3VZjr4Rmwu8k3nRGR5sAiXJP/qwK2CRraB5KIed016YL7Y2g
12qkNzmpC0+/R/mHthi2uE7Np11+MZDvfGunLPYh5Rf/HFyyUjqA2MOvhV9rbGsH
8uMF1cnJHcSAnMCKsPKkqjgvCkxVXkPxzw2kvhwUKOlqPFLMUOcnSclJsoMEHz4b
4ewSp7SjH4TPcslwLZ4EE97vD3YutxE6NYe8lMxILOTs/BMfdu4GzuU0yo03fUsB
wapzwvznv/QQJEviFyxgJZpQaZ8Qcnrx6pzU50dSOh+Aa7po1k5ho/derz96mL40
RLxZ6Dql3OEQZucJXaIyOPPIILFrmMc8ThVpYZebpuTFSFG7twiabCgXSLzzPIOI
ULARM//d9kjQ37quOyQjPn/YuV9my1tTnmmGj5zLo1qsO++VJ1estqkyIhFRBsRw
aayYCS3mDYSWV5TJWHAiS+Yf1dNViFgsBsAXY3rn5Nv4BDYuw4eEujwKGysiZBVD
D7k1H0ll94VM3LuWnuezjtaThdjiurA9skeFtNqpmIfTUJC9FXDhlc9GfufdaU/3
4z+8MX+0U4pDx8qf/sLPw7TX2vCK8aLlHE+eRlGNLiuXQen149YVdVDe6XCPK1Bm
jnLQdRhmKn7npT7HgRHj2NiwCC+T8jGXft73dEoJHya9zWQW0yNMSgsCNhFi3Nqz
UkXEG/UC6h9kjwmx0n9miEx9QcBalJfOPwFQ/++1lPcAqw16UscNF7ZbZgt3ujuk
Gh+tOX771ZrmeJ6/z6a8x+tVn5xR4hPrthJ07z5wOB4k1hOgCCChW/COUWBvAJqi
cr3EGpc4xbO9AhIP2pUR5ESPfz3cyvUhxtpstoWQcMCM2tA0TeR3YUKFB7rROXqk
IA/yY34v/V5/Ri2qBkoaTzQo4Iw5UC8VS9gLNqWxt8mwd9yA2c9oAURbo3zHvWZT
wj0ZMMv8Rj3goEuHoEVdk0x3OXnvfnWzuGqfVk8eyhvuCAUjHqK59/Dx0nzF+HeD
jqrzvXv0Tcg2gTaUigCuELLbGg5GY4JFUgwERK+HIbfSScG9GWulkrTUJz99Qytx
effUPPAl/LER+UK2U4xWELaDlZme/W0rfy68Pb4qbMzl3nmV7HPSOLx+HDbU5G5D
7psB2CFHlT16V0FKAQxtGtJKaliW+OeqoeGy1Sc+AxMiTS9KwE5KWwPfsvwkvfu+
uJPH1RUysrqSeGCt92IuGI5ytpxPL23H2PlmDufxlhmX9J417TVuqR2ZK08jGEdb
IVeDozYqqjLGfLOGrSIllGflxRGUNGuTJJIL9AB3cMSARaHbIuyW8OYhY19Ga52U
EO83G113GG0ls9QekEVUXEBL/1zeGyLniPHffIDgYZ5u6pJRW/pXsaDLhRN9zYZC
Quy3cJySQl3IzxoZXS9Y3QTG9t1iQ2CMomGSi3JmZboy+65PRpj0/hhOj1YI4Wlb
2DcBaCCf4wiNGUaDqTmMDV0BQ3vkE9Y4CuerB0dZBcpSYABPgXb79jijG0UX2XCy
tENugFmmIWtq6xcYkecUpqJe5S31Kosd21ZDYab27AFy2W5Kef/Qm1gogubOmakV
pMS0Ywubcueu8JZ/iN5An3K8KIrJk1PdKQGusxmvWG/bIrH6L8GgPWviKOLRqpHE
4lj+4UAm7AgzleKoBdQ2Oe7tP45P+vhAzkTM5arCw9E+qwuE/rqxJPbW1rJepW/0
cVlFIYhXMQm5otSeqDEnJ2+jrtCdZTsfOBWqYkx6okds3npeGQKY3bu/UWF0bYuR
FHVy7R1ac0G0ygK+vyeUMzyqjYessA+QyKjANp0aK73v+f+yaJe/k0cG8IXEV78K
3DITbM+ooM6wtKwWgChhxWqh3qbdwa+ttozNaqvpqt1dEdSnX9w+BBT7/fKbyPmL
CXr6hg6Fk+mbea/DjqBN8KFOcFqaMsJRKhX5eP0EDdNsaMxfv8AUtxxQEg2bFUgU
844MVNcb0UMih1CLIlvXhhSB74nV9bslMNjubljNdOpIYC9YSBpRlRahp5tmEP7U
I0t8zLU8yjgdWlU/Vp19RhsQhWH9oVsvkFpnOq09PCPqXaXugA/z4T1qyHfCkS/O
UevXqny9ZJXBiiROaiLSCtm/+Uo/Ry+kzAZH8Hh+PWFWwi8wmfKu2sQdHng0qRi3
4iLZNPZ3nuq0g4mV1c/rMz3aKfA7S6UhRXc2QuFFX3o4YZlvC4rT7wk/NChbP7uz
Y0gFlykUebfjTCoamCW1d2VlocvyltrZLZRQfgyOkWVY1MyFrolsDCk22l16lq2B
LM8SxHbPT0sq1y+tguvRCwJnZgonyDgKJGTvdRTXNJM4p0nRkhKeVPgJVrS0nDAz
7puJWLTcw7jow9ICdsKI07UoXsXWwrISUWs4bLKET7YXUZst7vnxhliFZanPwIvE
wbsm990P1YnbBRTIMukeAHqNCYHP38Cs/+0vNEVBvZOpxBTJV3FfKlgzuV6B+pbI
LMmIxY3WJWVSj+kAid9GTLdxfhfqe4wEzMCgoVy0mFgfqUyZZYAtwbUiOwhN5pAI
O4Wcq7bToox5D4O056ZN3IQNmLlcn9W/DScAnhA/63Hz2jxQ4ek4AfFYx29TteSB
iIaPwrRsJaV5WJcH6jPaBhlSpUXj7IdqstWsJgon5T5Uql/YLXz5XmZFkCncWKQI
YCU97gNZtqjrLEGpPwN2cO44cu2xGbg8XgSjh4gsMLv27in9kF68mMYVb7GaTRV3
J41emC64eTtwq4apJ+Cr4ycQrgFSBk2cJDM411EOJIr84rbw1d+VnmMRS8NiwMOl
M+sMgJmxBGcBd3RCt9YD+VWHBZsgzwKb4j2ervDg7RArqDL/+CSnQ32NtCGjBM4d
4CyEscoV8+ik1fAe88FfhrXr5zXlw0s1tdcVahsTYWWoL3R5ln6V/mB24khJliIu
9Mm6ZZcYhu4NGBgYt4zAdqAWnyCJI/6rA43HTQW/WM322kINbjUpgqDaGWTQwbBH
U+5lHV/eFgIZKSLCdgoqPyMlJq/QfuxwkPk5AJkxJnC5rr/U+aK1QXhBFlS2V0rU
ejkyGLZpPUMkFeDtxARtG27y886nmsgscAjhfar6JhOhRMLhCT71BHMqWlYirwCF
XOi+NBHZuLYW2WYPkFlKHuTayFFIcVk1nPbkBE4RZXRoDDVK0P8TJ/rhDLfGjNRO
PXdnSieJ5/jxy3SBpyBiwNv5hWWT8A27pEI+kscBOWhWJVm809gziP6pBSC5QYTP
nbbiuiElEMcmEcx8DPx7XRDU2N8sO1yF85LuBZx8jAQ1dhdzjmcdgKG4DQ1ImEkt
7pEteCu5+twRjijJTTn5vb4RQdBostPamRmz/AKPG1DF8eW/dmQZv4BdUQffuZSt
ywchYEB89KzvT1OrMgc0Tn2nXndW2DOI33DP0/9GXaSrMDROcZ6IZh/bAu8+x0gS
VSvRup6Z1vq0SudqTUDU27M2FrXWRBJLqhV+kLzYdCY8SgviOYn37RJLwgZbtVdU
44lXxkVEy4MeSkxfUcIkNzU5CaYghwfveojKhZ/CbxXbrLhXB3wBKlt5d4VnXEKB
2VgG+rFfcKCS/EweEpWN/SajQKb/NekY8AWfF5gjSOriF3tktndOa30lRQaNO+s+
t0yifQtnFPVB2rForF8pG0Rky0xd7Ex4lRqrfAqxoNWimWTPi6JlJwYccJTq17KE
6O9eauGYKO0HVFqrl0xKkUP9KmifFz1+Ir9JAZK7Yb646fIgM/LWVxAvKlSA89RC
kVy6EUTX5uaGK7N+r5wmPxBIUWAWPHP8R8kQx8/VgQVYivaUcI/Fl3cUJrwkz9E4
CvXWdMku2ST5boFkTlmbQ+5uPr+UIPEnaYmXHaatSNLoK70sJKVuX4Lfo6sJhaA2
BC1SZg0SaaLTRM2bW742LZlM6soPtm78gL6ocdlUXKvrcPYKlbKZmYsnlea8y/gZ
Ez4YOlKq8VAcK86KCMOiS+COYuO36W1XwvbqEHSinzMPRasTQ0kL11lvI8sHF2Fc
nini009n+XChxLEasGnQ/mtqhWbqkbGFzqVO+MqzQcai564ugt80XI6ctHSiCg2E
Re1o4qC4FqKc8E8cQ/lpHaq81HmfVevqSn4tSVqBJtJe8fysFseIfJ85pnsxQQWS
ERrubCszIdjFtWgDjo8PMX3dwrl5+Zsd+BC6cl+eyDZ/avKleS4+rGwyM1j/faaX
KolsUv0OvbZekoFrxMMz0Rks8RWgvQGPvMi9/3agbWIBJ1euW18tqJcw329MxY4P
3Pzue+nlzRX4u8ARJhutpMaeVcpHjKmWeAIkra10NB+OVfSz2aalySLclktg7Qwn
l9hKx8uHSwwyyg4fYIQ3k/6w1dmTJRzutQk886GpJqcFp7Vy/m5umomdHINf7xww
hbX8Flc0L6Y9bQESMWap5f1wBYRtPx31myRRU36ru/Y4+LF6oKrhBdDRXNpXm5gk
ZEdPZQEm2dV/KMofwJo9tSj6nb4qev8tJHhG1q+6mla9h9tWvTcqbdl9isf7Ix1l
wgTYxLqCWOd2wxrgukZkIVBSd+PZJPnqkXID9gDnTFGWGDGmW7BfdAxx2ip53d8c
1Gv8nT5oTcGZDDOT59m6OAY7sBLm36GLdTOkj2TmNNaMPF/XAUPCIZqYtZ0GZgIK
6RJN1aRNSQhShHZEcL7ohL/9qFab9gV+bEcUp+E0JmgBtntFltaD1eEcm16iu3Za
WfqL2heW/5G/mHQbZUgvkS+pXII93ai91C07IN1E8rYFnvmasoRZO8bb0oHKPcAV
Mhj3NpNJoO4UZc/YjEyeCJbu4U2mZeIStndDi5L7GvLXAPZgKOReweRfV+Zgd0cw
rPD7iQPHTBZfz2O6sYBB6n4zzZo3Rf8gxGJRkSHY4hF2T3qbrAptJv0zskRlwoXq
sLBPMT9bNLI8fFJR7xSrvCd0S1rOJC9OYdgWqRAdHcK0NG1O/dBekoqPBzVCG5Cg
d3CGPtXA+qnh5sxgACeBP4ueU8s/ixEGS5tK7gMyPPRyhNTD+89/s3YmhTiYQHbB
rZI6ueib2IPHRnxLPpAlS0oR0l900khAxx0xM54ynUHpIJzC1nNy7pQLbZdqDRRj
bdeUUX4KObgEGlziW76RYVpNSolut+ucERamcKNMcpY=
`protect END_PROTECTED
