`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3O16uY9Z3cb0ws2PO3kdAIYM84XKld+5x34zaSqL5pqH26k5Gpw7oyrk0atvQJBf
wSjcQ7KiSnpudeBjOL4o30yDoI69mUudpOqShcZwsLiM5CDp9mrWx2CvHIyVbiSh
u9WwjXiu3E89BwIqlDba2BucWMPwrmX/4cu/lZTxvXucizJ4far/EQgSMSgAnC0j
ejdLf3i8UK7DCu2yCJfCfHU57jyg0zEvxl9SGFD31KOCem71grEBB8DCNDcGiwQb
xtzClxNzajjEfx4bDHKyVRUmPEy3gJqy9YSovxTXn6RDYsPZ5nP+d2/HLpAz7CCo
PI5Ggu5dORDkUtLUOjsr2Or3gP9NWFozaWj+4+eUysN819Xq1CmS6m0lPSIONEBQ
HEvG+h2zhMMJNdPyGpOTR+HC2bfJtDf67k8p9idLVCQuvCQ9ypGTAn7PLyizJtdJ
xMAk89JU0XgpyrdgKqkZgU2sE/iFDBlbKuhc1yD6vhh4MJuz5xxw2o387ddwN9Rw
ZwxID3h7ERX/dkD3cZpX1iBSV1K6ZnEwPKbqLaatoDip7Zk/fgM+KD/3j722iJ+f
XCiZkFj9ZMF9CjP88Swe38zPPMdU0DsxTkAt4KhYC5B9FDzZPLw4YODt266rT3vd
KxBl0K5ee6S8yHuFVc4NRdyGVcwe2e2WH6tNIAILL47f2isID1gEe7VHMwaqcNq1
Av5NVXwQhAWE2huN+ZK5E2CktfKWtyCcOlo/p5TAvYLfJZz08wOvZr9zUKYXdESC
hIvvcaXhXWCJKE0JiETc6soaS0fKUz4vFTnPXBQjEoRQu4McT0nkbqLjq7+Mk8Xt
zDwZyoIdk99HBl4It6grhuKHIyANwH3ILZMe/KM1Ywx5OCqKhFbDkHYBmBgyS6gn
3EVItBJ1UbumXgHjLghnZ8quO9wT0CqZj8Nq40tytjqQG6geprd/gMjZLsZNYnQR
YXYECINayy8NyUCspbJmT2w2ZXnHX9qZcZ4QnxsE+udSSS4si9sWnFQ6TBU+rOWD
yPSdqnbahW53GUxFR8M3CRkPX1EZ5dooID+DZYVHdVjdPG4x5AHuBw3zcoIEeNtQ
Cx1uBlPq0+cpoc6Vo+Dl93FxI5jDUjgc06w7hJpzO18AZZeKv/DSxsmwerTtmaFj
cOM5bZBiJqnzVv2gsJbAauYVNIqt4F1XzUyQPocDyCJKvbk3U5TYAhYcQAhSeLkU
t7heUmsnVXfW49xR3EgmWt0W1QgCAlwuiJxGywN7gU1i0/caLF7z2Z6dvnzlJQQp
RBdaQ8XqKnK5mF4HWYo9/EgverHQADHIASs2SMwZL1D8ZY1zPdh7bi9vL5UHE5uL
znNlzCX9Z+6tGQvqcu2FCp4zoSlbAFkMD11/W4u3ZYqQKYil2RbYguClUh0fWhgf
8c9jGmTdoVYOXLzmP6FiJ9nHiGF2VotlAUfuu6P6AMQPjnN0P/ESzFb1mJJ5/sTq
DVNYoRDjQ+hX0NKUJ5ow/gpSKTumr3FytYbOmVxeqmA6ISrpK7YIktYv1oyEv3Rb
2FG95n9p7wwfB7nG49ko/xWrUfhhXr1OkAvXBTHVQ8wFsbE8vFvt74NnULanZmCj
01bPjScoCnEBI+3nFQnndRpUqw17kknjbgDE0jLKptpdbriJiddvqYFMGpGqfn1x
uMOC5oIjttuc8jc5dthUab4ivriI+jQ0dMQXM2WGmic7F3uCzA1UzBeWSbq0P7MD
i5/L7SQcosyO/qLpb8uq8KkIKH8qW2MhAdESH1admAfXbuVPAL1GkfSDmzmAYcpN
PiKtMf+oU02Ur5I1/bVQeNwaeukPg5H/QBfodfEP9hoQo1t/XVo+gJ2f/aYFABJ/
jZqEzyXcFZEmdnVtJ+VVsuhcAMt/A3F284nK2wECcRh7RudF+Dc6yyMDW25QbqVU
o+kah3qv7ozH7RQkOzhTjBw11bNi0ikwc6zfx7/Kyh1aof+gBx4dx/ZTK+OvqwvK
0eh/7T/3kxhegWGINPsLIzqG6JEq3cBgEXGs7dt2IYk75dX/5zmf9xHeumZgmuYl
kn/RueHHaR868+dvYcaA7mEMtuoqByjtg2D/HO3F4Vn7nZyoI0fKKPMZa81KlRww
MAJ6ByPG3cGRD5vBH8Yy17gvvmpz1jxpDpK5d8Q53d4=
`protect END_PROTECTED
