`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EiVbspU8INFlvfFpMjce2Jd2mSpl45DnTOSmIqFLCor0CfV3wRd3uyMHnB0aACco
nc3tdoUE2MW0rZLw4AE1i+yL+MRYuV51Hvz65/zY55JRzFhTrmAV1vF1EGqOL+s1
DnH1SQ10zlLaHJRCEdimYfI6tlNgpj1htDNFleei6CpPBLNdQGGp57k/Z5XRAm3j
dng6P161pELv+DxGsTqDC1zqMU+pwYQlZkl8/PKkEnC/1Ul/s0FLtIWQdPSlvzS0
DUy59hL1u1UFj+pvv5chJ/Mwl8kwvkMogtfPmQ/mj4ZHkWG6FIgVoTGMEyQmLjIL
w8OsJB2sg1kSraJdh7m6zKQPX8IXVjLTddADXAWB/Rl20gbxqvpbDfxp/dymPgUl
fcRIu2kNyYK9fjxbq9quUpAh1TSRFNN9RErNSmEh2jVhev3fos2gjw7ow7SUcpyn
EjztXjMnB0aDveEc/qWN8kO/N5PkD+0alhys0TW8P5+WaHTltyMxv9EzpOospIHG
1YGdAOrRu9ilHVF6JnHETj+cjs8IDdyWlx0xKltHhhP3g6QmWHuWGuHqbWv4PUYc
R72Odws6/yp/O6bzprzCD08NqQxS2R3HGcDWmm3TdoFTnqF+BHzn5197yQ/Zw8SC
5pSvkdioJRNRAVUhb2uBqiKfMj6D+moh1aZ9acxoGjSmJim4oeiMR8IVqDZwCbN7
MxQuHmqTYFMyfJVAU/5VRY1LVaQNZEwro6HUaF1Ouvg3yHGj3cG9KV+aEaiBf0+X
MUxEOBEL35+WAR9VIx2fc8XYTYR3AIdYCzbrx/xSva+SMtXTvVdeJfgDDbrrXXUS
ybAW8F2ysG3TnhYzbTVCKRB7wpbHGbQ81Vu7YUCJP35yr13Grm1e9kmY1q6ghi9T
LAOdpi4eGXmOC06z05bOmT6HIu3tXUSWZ9FiljO3auj5jMvb6oG01KT/i8LQLt4Y
urLwjBpiVEWOkawcNESuP8jTnSZX27ZpQvEmT0YzmeRhKunvNOmgvckfEKpofs+u
N++LDAADIY65/7UHvTN+1i1siWie3UWKcQeERSdTpv9UgZNqJVfBVErOVGoFstUj
p1BY7AGXD6p+dW5E7Jng/eTyWMObbqR+elzBzHGxn6/Gw3qpmusRQ3f9PH+tiRbq
eQArpvyF6DakNAljqPzcf9T3qZKm8vsugcYIU8G/sLpkTnjWhZ4GZDnmmKk7mazr
GlteHDV1nC67QMsbQ1pyPEvCCIreqmp23alzeYz1aRO0++eoaoEw92z+7ZS7UDy1
YCN7jMKWImB3mRfEdTh+VvgdYQwrGOUf9Xk2frovHJSFjwkCXSzVHa2MBTfvAsse
p9bxse0qCV9ROa1TBsdY4bcTh/lBl2Mrqer95qUDq/YRjk+PQPWZtkx3ZlaTnrUP
AiLuOGvnl4TQ0V10h1zCtlBhYIG9todEQHPdfzbKVEMDd9PFZjpzL19C7JJMFD/+
sNPl+2Adag44pAVNPAsp1IC6AYuTJc0ibie6lG86WYbxueZotXkxDwAlLoUaT6qd
EVRX8ibXirJ+ReTJYldpQ9EjLd7/m8bkeCWsAeMeosGp1DTgCHK7SnC6HegPo5lP
ZnjUq8wrKmnleZF+qH/RUZYnRuKwRPgAQI3DyKwtAq9mQUiHC836ZsYKIhbBlYuE
WF1Rdv8cl4XOmU/4njHwinY6U3zu8mqOcSwV6A/x6ZaLux9QmoUJc1fP+L5xC1ZU
33STCCBwYsH56e2pYIMzJ7rKzmFAFwKUkiGUuUEkVrBIZR7Ze4edadYUO4nw40tB
/yi6YcIBpmN0mbaV0nYJ7enNXkiIqnlXMwI0p8/n6V0FNiPVnW/8w+fYtuxiPTsk
mLEv99V5K+4luJ66sXrvrNHyfTAr2SQeor1Au5FX+gI1ikKphfurqKmWfpOujh7n
S6GFFYu2bboZHkj93I33977yCQ3T8Kd83jxT4mq8Upe87DTcRcBwrOOUgzmv2KQo
9g8rJOaJrpdv5n2qpB2VgcF6nVD4fSZo8c3AkbXqPe8TQJsvOtohcGtaHjgqELXA
YAdtli9ryOVierRNJy36cUebmgvdck5zLE4ZMb8UVofNIgZo3S+FUAS/zt7fngSc
/pxprHK+ASihnnVGFMYGWbDV936Q4grZpYK1p9Q+tuaQReZ4ioBEfXKOOkVIAzuS
TXzFbiGjchDard0Am+V1R1Y41DQ8HHh/uMQZkXpryNs57ch5rR0lH4ysGNthQcEY
yKh43qJlhImEHUlJkZmAzDHaHTybRot8A7fQPRgMCZgHsLoTAPbouwfFQRvvw7no
hR+SVZSbFlpYF3NSX85BgmK8wnVNxtIuA3Hp91MDd0KAb61oZ2mcUZaXaNwAuWb3
kUJRqYwt9u7or5hJ8a7Hng==
`protect END_PROTECTED
