`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQ16nafUl0HUZyJP3bc4JHB8NOo37AKB9htom3wNcFqPX4//uz8cJBIpkVx7brPB
4IZJKrmt5GZ/UxdNHBLTP/zeEczm9gf8uzjcqi5onmtiNAJGYW2fqrHwQ01RZatY
qIwIvRt+6KtuIgsfou6fwy0chb0+t8LRfaBsAu7yq3LgGp7ag+PUQmGwAWuKSV1C
mPAhnBNyjqVcNdh/uxvdTJnS+Q5d9rid8K4I3p1bS3Y+Yfr2Zxt3JKZvSmyW2R3Q
5/3vOXheKXYpEYn9gMhoo3bVQu4OToULiPFsj3B3KVCmI+r6sg7U9FqRDL7Rs3uF
aSmUEbqxSuXXWRMHTVMCUjYhcSCF40o3fZLBVKvHfnd1JxrZ2AH4uM8kC32UHq2d
yVgLnFCQYCuSye68Qdq6xPKXi+UseLHLEUgTmPrKL+EU5oGqsDpq5yR9w+Tpxwub
8txF9X/Xl6qij32hZ77W58zQpZ9hnt6mQQd37R2xoXwgtMkvSZgd06Deje3g43hw
8G/7we/E3V7inLq7Sx1pKQ==
`protect END_PROTECTED
