`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G+CvysTBMhRp1+LxVTJUUhzczczIVoRh5H8olarA8O6CzogGPemuZciBG9GH110W
28r/LEHgo9rwrEmC2AnJnHc3lULmF0J0cNRk2pVJGWDOOQ9VZOq54VSlPVNCQEfn
abBOF6YGUiNRqyfXu4QpAU+JMKjnM9172gzGFha7tXDi0EZnmnubREpn4+FC+4rZ
rgy5sZ1Mz9MFatrVZCV4hgMq8vd7VrqtkJhcznXgj9K0ULeSwq5oaxqmG5p2RWbC
6oQX9UNOpTPcK7t8h+558if3vdGfvyGnKgqeKRkeRJGTJg+07AiMIN7gsk4IRHC2
cv4SoeWiupesj5QOa4l1ke6Q1fW4Vl3rk/MXs+xki2B9FXJYUOYWjTuJTgscFH8/
4mgwWAvkY6hVXaovRHh9Vg==
`protect END_PROTECTED
