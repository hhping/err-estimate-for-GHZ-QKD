`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
up9xf2WZ8X54gWRmBsEZhL2Ho2tgGWTZRvmShemxZjWae0DuMWkVaMFgeLUt4/I1
1Vu0rq2wGL5tE1zCPSNd63gfhjQuq5QCeuieRzWDWRgNRyJlr/Jdn0jBPKMV1WW1
RLx8bjYQOUKImhtQGs9RbEQrcKGZo3B7iAAgbjYg4E0fvFbrS5CWRVyOaCWxt46k
uTG/RTCQQoCs61OWMPpWGLkF8vF0pJdUYLinurgLuBtQbP06dLqFAsxEcmhBnIcu
VC1Wpa8r6lK/XiIcSSfhtudLT03OpaBVI0rElgmlxcZ3uCM8eQelb7pok1PolA3e
wG2qjTWsAR+xhQ0zA/jyt89nFo5nRu0Imlni2euMK5KncwSEDcc/r1TdHeSvezsR
qnwJxiExBh1n1UeU8liIYvZveZO8SiT6Jr9l8GC4+y0oFkbF+etulkPun1p/Rtil
6ZQDEFwhKzGYBJZCKku/fLVZJGwCjG6VOn3AyHLfrfAee0Wzgg7yo/yKM3pyG+9i
`protect END_PROTECTED
