`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O16fqTDbDwyjWtucm1QP4d3M7Ejhdby//soLOFs/LHGviXNrkIsgtNc2iVTEwK1Y
CEW4CHgTbuRWLrBnYMBMvOBT0n23JhDvE3rHTgclRpPd8x4wQYVHkd9sWqgg29Uk
+0wUIfP7zU1DvOhvrjDWypt03ImdDBfXA09SHfnK/rk7OP4QxwBTPCPYO3QVYkx4
mO7+YPVrK55XUU8evdSNy97THu55VS3leIVGDQ9bP95nEBbFsgS76IiolGps70dm
kVbb04q4pEVfDW/4rwHWD2BVcsWvSY0HtC+rv8u0eGtZtnbjjklQGojyapavJ5Hs
Mr/G9gV5aGjQLACr232m33pqwre9xZONr5Y6qvXaErqHryMNPB2Md9devG0YzUa+
Ompk2RLHxQlVGXlZ79b1HYf4zf0qi6sA9YXdYVyOC0G5LX3Yu0vAABoZIX1kx8tS
A7p1U4EnuaPRVZnHeoE2/LgbP3wqA83Id387fxXSVDQ5rVZZLVAo8cRtyu9JT9hk
DhHquK64Bu98Jyi1UBLcnB22SGkRooeK0lbe4T0Ayv+b9zYLaZzcWOfaeaFjyv3C
7Xe9QncEkAPAzzeUDAkerMRBmQCePUkJQ/X2woQWwPpYUOCi7josoodbhsDrzBya
Mjy+6oKO/SmlnS8lTne4ifFcIgHvKdurMjOSb/TPtq+N9GYrXMaF6IIVucv+cMFl
mWDvoCdrIlrWIFa46qYtf0IBNEnpR6hmoLigDlAoWTzgqrhbVXr6Nz+Pn8A/perO
0Cm34+cwEuWOFFiWz3zmjKDHkew70osU52FJZc6wUeSUXVG2YBJTJtq9oDbGSqDo
RXYQ4/SneA4FEwzxWFyatLtok5r4R4naUoktVUVk2JxJa1FZl3skWBRVmx8GWzGc
tC7Ik/EckZk4RUgvO4H1IY3tTH66YCo2rgy4j+fzG5pURKHA3R47RmNjhawFFbeZ
z8obM/MurYm4f26U3Yvm/brvqoATJnZf8R/kfp70fl1lwidzLFQ0vSUocpZGGdS9
jQqyzQKI6hjI7hSm/xWr1sxkUIHNwgOeimPkOClSY1lT4SyNp8zEnG56NvkkaZwE
PjmvasoHF2Vj3WJ+MtXr8k/tQk47IlMHDme0d7ExaGndGSoEUTcHUA0y7CtzFGB5
vjEGOvCmYfYfZqwXqswYi/oBs4rYvAFJZuIuclNQTivkx40SBc1IFmi9lTN+aF3e
lX6BKDDGMMYjmlslT2jLRsgdUy/NJrEZDBHc1NSzSiA/+QrZbgqaOCQ5ikNNVcy+
3OSIRTulLZy1r4Uo2yYMpvy3PqC5ioP2upIpMDZSVn3M16V2tHtGP1EgNYPdtOPa
amUhoYjGVFtHze1LLOKh6XOlqSrKz2ZIFHQXLtU7+XVjH6RFgjmykgxpSjx5wybL
82kxtFUWF6azIJlS4WcJmoWZWjGCz5pC41/KkcBn1kk=
`protect END_PROTECTED
