`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AU3ye0eFRXobmybe7CiaE6Pq8fp8oyvuM7rHiXZkVHJI8iiVp5+1Dq0SJ0hP+Xfm
GYy6ZkjUmTtOMvQKEX1UWN7lzLhLqD4HrE3mIhUIdF9rsz82W7MChHjcxGpA9pC+
zABJPXQrmnNfemRCxUPHw2NpLvNAI88bDctFtf/0p0k7ww+BXrhS46ZT5Pme2N8Y
OrqWI/OGIcQeQdX/yd07T7m6VvrHFazLMfk9GZYN2Lt2hGD+p8bcuvcnwCKy6YAN
hLgTY5dyxfvhxNdsTOL+artvaZo3vtCBtzEDq+PTd11es7Cskt75OY76LJQVEN02
1Zxpzhiw601ZY777hkHXmHIxJ43UHejsLYh566EWQ9X+gozV5gOiQ/LcLKh1zACz
i5dM7EuvrSqNeGBMsqRSIb3AaJNXdTJJR8vXrQtCvlAG73wHlFO/s3J7VPpXBIUs
4/j9EDWUsYBrAqexjGxomIWDvMj8UCEu4WVnfGAXO40toGsGM7i7qf8nYrjPi3sc
+74bV8N1zjI0qo3pc/lTEXsWRXSDJlG2WDsmsSIxV2oZ4I2BGSM15QNlIm5xGj7b
6rVFAB6Tjt+GodFoiN539M91NjH5ZOPElIwzAv1h4bOdTxNG+EEvuAIwZQx9QRKr
YMEmz17hBYpN3krtmJCp2gPiLhh5jjlpto/OQcbg1WZkm7YUIbtU1NEVxfhUfiMB
hVmre1nBVKLyGlYuOwVBmNp+BiKld129vstbDNF+pXZXG8LUCVFjKJZtKykkWSmn
m5RnBxEANq99Kh5fr8Ec0oCSDZPjJUSbA7DS17/kRKaG5CrGVDf8dEQH44lQz3uZ
H9ja0hJFF5cx+YzELPkgZT0FeK/Ikq35SC+YIP4QK40FDyjVn/kNjHrrvGr4W2M9
gSxBXMwGWd82e+w1Jvn+/6OXcmGuTa1pXX7R65Mk1Y4Wy8hck0qFRYCm9g9iE5JJ
C6AU+SdE9Kzt4wnM8UzQ0O7246dLJO0/L0k6ab+Ry1SoVzIdCp1BGVVPurKFKu7D
isr3Tt6kNs+PiPhzEhQen2D8/U+v73/6UU8nvdBPp9L2dJ5+lvp0Z8kx4SvR9ziH
XC6pQv+LoxoOx2afYuQyKJV46ubRHyyIvOGm46+n1CjZn7arfK8xk7IvVDmuNbmP
dXfBeftQkeyN7rlQsrkK5nJ3xCb0BOAV4v78Wv73Epr3HQYAJ6rSJxNtzTpJ6OXe
rDGbVeH0Hnof7aNQBm68pZ2/6CO9/HM4LQ8Ji4tdge41I+dkCrXESgjZZ5QZKUxR
UvbCWGTUkld5Q23IBZDLf9q1NPj/DyDiT4jybYmM4tpnbaM/wRFh0AG6XMscK3xj
N5ZslbEDZHv51jokYDwswHbzP4GaRuLBmT3gWG5IbGmS8qqomwH+MZ1D+rUKPVs8
DdN/UUXSq8ZyRAlyi0l0OqoASqD3UzJfyWd6y81HOfdvmCmkA2atP0KEsZWLIRY8
iF2nhdbKl+S5Iu0lxiTKa8WpakFeaCVFDADAHtQG7XM7RqblAdUh8RT1FD18lks6
Gr+G/4lcsak1eCytqcIQVaBqA7/+3NOliBEUmlBjv7PPtSoqFkx3t4FNTf0+Ltw8
57t06EgSCSrnT/feO9uxT01U+tES2VYVmyJThGUUr5A3sK3jC3GxzWtQrqRdicVb
RwBvoeRPjSFIOrDk8CeP/9LOYUc+lYGtHP914+si4KUr0JIcBbcfPqZ5g1HsAsNm
Zb6MRZCZx3+B/Z32S02MqfvkEfMvz4ou6rn9YCZKApnCj3sknwarVb+/FhftFcyg
pDtCyEhSKTo3LYz28M55mUOlf0pk/TtXHqub9FtaiQdFO+auU9gaa8u+Bm5wMZCJ
BKv5SKMjl886LA2g1zANGsIkbBL3Tv3KhyRUQ1J700bORvqcTbSJNcJQ8XyEYxYE
H9epNvStCGDbgrBqwWqhn1QaXjrFYZLpT8HYDMDjDIcviDhGQTpG6ISaWK0JBO13
tV2idZ/YdneH43YmtBSqviqCht+BqPU4qxsfloNZs/Er7Dl8TMwJTFgG0KaQhA2F
/2m9QXAr8muhCUuoa+9x59E3EnXOaoLKEK+yCbX7OjMTZCC/GcOJSqEYfnoBENJn
QxGe6bfn4o7o/Nh+yrUpl0+TdVaud/urWqAMI0GNEMdsiSnt/Yag15u9uNzCUmn+
K0QFTs+chlSOAhAtHDxDbVA8QyJeH4Tw+F3OMrvKb4YGPP+7vCR/qv0douTeuncM
AwlElypdKwo/xhjqRy/b14wI4SdjumlqCaX9Am3vZH9IS6rV3kRQt97sd3wvh8fS
26XNaLXkTq+pfNQ+hbW3AWdxnydgZVn1kIDynuRcN9yPNEHHy0CMlSdEaxrPCN5O
GjQAN5pnZPOZ9l0nkQi1EtcMjtJQ0owrtIO5b1eeLmBCe6A/OAWzrE/mK94Oa83x
sO/e6gvcnQ1HUFRr4QjKGFFmttIX5pkDX/0ni3SvcGVmpA/4coi/MZeMIVpdkJWV
14A9hnG79JKNnXQWQKLpmpc3Mr9VulskxRtnWOIKksPkSPas3ZNGpz5piFlWZrhx
rDzovWl1M98ZtemJ3mO8jGrvp8vn4cYckcsaRS+TXFMajdn8reRWQp/VdSbJQHLB
hGdy3XrZvsQakpOitX+I0e9j1ww06c4je8KYA4eSNr5dAdux6cVHdqgE69gKtoVM
QQ8pkY3Vkma2sUmi192KZ8lPPO59KzWbsaFzyns9ifttMtmnQJSCqi6dMoNXI0IM
hGYmlMBzeBaoCUjFTW07A8DALkNXtu4OhlBA8kdu+RrbYddGLqNyfK4Ea2l8aNQY
KyQzqgNBJJ4FPAXkEz2GdQxsNPA2yIEHRwIQyQoapv/aehoFJXJLKV43Gk94oEOp
9o9/D39czEq4m9bDw+K7d0ZgdCOeaz4gKD3acQM91O6YEerV2vkrOVlLakyaGb+2
RLjwWmmPEsaPYI+5igDZZWvTZWHb07gJ9FTsEQvzrCoSff1NB+LFb1WThkGJbv/V
pAItmMHD+/lvO8lSxGWQ5w52ReXzyKq0z3xhtnojXXXOq+BUuD+IKr2jSbzY0FYr
ZnFukGJkFTxH/RoiuyU8Tt06tQdmWayBrtqBZDWYdRfAmKrZaAHEkb6hjNFR9/po
pRgPsgMeo9dFkl1sR4gUI6dgbSG6od8csZm3XpmfCW709Y00NoNFT8sU0PHQc0JR
ft6rBs3GH0H1wRuomDNtuvyxDXDICKM9D0LIIWSoEKoDA8Rg3P8wG6KwjnfUINpD
dK7YLm+Xj6gZloMAE96kZP1tfSSu5nHh9N88zfw2RyC+sO56GrhCUrRcj5k60GNx
BocNO+1S+t+qIFx0PdIrgvA7ILz0jQ1oTClB0gyTc/ccKyLVBJGBfp103XxdkNvv
GvpO6nh3VFg4Qji7KxQGUdd4myKaFhXuSSGu9VmS0/MGCYFi4FQuCeNIJvrrTp+Q
ancyLyj77j1lGHnEmeiVjD6946ARMbKy3v3+hZX6okKC9VTyj4J2QWp8zkUlp7dZ
1jv7qnzKBNz4KdTlUpWvqKpz+4v7XXljQJhXngIlavL73QaszKcYM2mwLUFvkD6z
k1rrtcs+kCkhezTOfgWHhArpPPoO1wBaIW6bEC7I6jrM7G+wpDSdea9a4JOnm0dU
yv5c58twtYWWLo2jj0z8pTh4Kjhtns6Gz7+TEllkqKGGtvPhNDm/H3Ay3yXcdL4F
/OPoIp1gFH70RwIwUShFTSOAwBjvcjkgU+PCUnDm0VVMgFD350x899o3BdtR7YQM
mdBhBC4UBZ1pCt7sDjWwh0EKyWiNZSxYLinBqga6mALamnmzWGdnN2CqIibPv14f
ncxYhwBuzaWIGdRGEEsNX+pCrE6Wuws+fUD2JwWoFan/PmIpzbklR8pIQPmLxZWX
besFcuaVH9c+68xsMhImwoD8AJdov0gLa/ygkVZ1BaZT3vY/HnRJNvhjLqoen6jI
cAn886sEwvNpMSjmK6zJZIr9RR0D0MpaeI6UopAkSiAAwZMSM5zsrLkSCdWoz/fS
wRYJDBWAUxwGgcGtSnHhGe/gT3YdrrhSEdYg6/N8SOIZfm2uEdnVKXIREIWh3Sbg
CLpnjNbcg0p5ZxAN+IgSW59FOpe5UOo410fL8iVq5++p93RBLhL97JYffAQj95Xa
d804IxT9u7vTpMPqAdY2++HLRHFGrrIyJ49f8UgXqKg/t57AD+qsnLOeAlk0lGeR
6LmLBv8wojfbV0vD+9MctpaKlJH7kAMQ9D5kflKNFm2t1bcyhcWe6z2AOqBpqzni
H+/hkMmOqkLsl7UEXKza7pqckX3U4JO+94BKbio2Uu+ekCKBA9MBDONjsrhRmgUA
wHb4FSz5mGpwI1iV2nIRM3mAJp0UNoEGN0esGMt60nD+rW4MBYWQeuD0LKSi8e8/
iovnhpdKLeh6kGLOArquQzM5Q5g7Zu/CaHyT3tyWGfttawc50R9wcq1AwEkGVKN+
RUXCjEFoas/G9AH93kkrpw2YlczFfSZYLOWjC/GiGNZ9GnFl9CiyZzwbP+i4q4zw
pYPMelTYS9l9M7PasSAypuHppfBBrpat/pjS0nlIGx0/cRgveV/D0qeiVHiNlxRW
88Mxa1gaW4tuXT9MFYBnvgE+DGkOOPHLI8gmCrRXm5UXZbd3MD8XkRnW8zLxcMAf
+hQzGEWqxj3q0bNhuCElrR37wg7Kse91EAvStP3J80GuxR8RmpiLvcZueHMLeosc
QBK6UnV2xUAdLVE2/aF0PWmiP1IfADq+pQuSKX9O53OL+5MZbWDsmsiiE5pu2Pkz
EIwbIBjm6Zlg5/TRMBELIobKXPSpWwVXRSbnu4c9l/Wutr1bGjXPFmGi1WbFiKhD
NeVwZn0Us5Cqw+FksNCAbvBk4QEycqoWxGyLmoDpERkDf3+PlggQxBBh0DdaAGRL
BBtqs7ifOcNAnkmGgP8QbLeJsjN0r/LjufN6pGGeie23ioI/8w85pZqLi9bidHmf
24VZE8GAPxs+EWoWH+cU1pLmBT9bhHm+ITW2VT714cRM+hvLhPEAMsouJrV4YIze
ZgAAFaQ+9XXLlieeR1Khk3N4N3pf3YcO4aqz2Fq841zuZe4jsj+VKCECmtsXcjEM
HiXG/rxrdZNRTHnYywUQfnzOG4q2o9d7DfS2QOl1HT3ohIjlPOWKqaGgF0xsuaq8
GP2tHggibFXJZPqH4f+/5CHxV48APer2LVxnZWCmMWBLMdyGbeHZ2RPRVqehPkDo
EbBoqTJlvX8Wg/AxzZ3kfV8tpijXGTRE5vpUWfauefP2UjIWzf+CzTIarxGcmRUk
p8rWnCKuRJ7SLdnBJqfK6siQoG/OnyxLVj3uKH6cWrsMZ7P87TAuAORyJ41SFCDD
tuNeZGC/Y08k5s/jrfcguZ9KRWN7v7uSEqFRRdJwFS3CotSGUR2fBciRLD9hafyn
pz1suyqayshXDQHQpUZwSUrYBWc18rWQBTb/hbaf8GhtsO3Oq0ycRNEJw4GIEkkp
qg4LjNXzTtd1bku+JmIGx2M1WMH75cRMaFXSMeGQhUg/rJaCrSOmYWCwipNJ477o
b08eGwANfb/+8d27KBANH4VmBs9WhTz4HsfnrHhQeUoxZgHwJY6pd+/ABmvkEk0u
kvSE0m4ll7ispKv8MEURSxajHRq2Pf2/Q+gqZl2WYulyv8Qz/FkzCwkcai6bXxdZ
mZSVl59n9d6KIPp5U6JeWPlfQD/awr4lwEgRagKNQJLkqEckypIBr8RHfh2S/GkK
oGl5RNpNguAzUKofBh+D/B+0bJTrYIBldrkeLyZx2X5z9OkhsnQVkWR52CjZI/HW
Nyhpw6WvZ/94Ej/FDB6v1r/sStqBjTcp+SRqyv7334jM/ee5UTy/4EsqaYf/dpb8
mNq9wlhIQ46kNXyuQF9vBx6/t8uvbY+CrxV6jsIFnDfStVScPrwcVZ5UZpIupHl+
Y6mmClcqDTDG4/w9NjIQQGmBFhdLDMAgv74dir4BOzNxvjZOKmx8BDCTAjbuWnCU
QAzoJ5u/lxsZH6/yUheJMHB1e3lAnTM4Bpn4ygoi7LOoc39utJfSEbgCXrLFUx33
5q42DMgWJ1JgyNt77zuhsgjXaGxIdvhCzQpmeLq3r/aZeHTKqW9siz5TNkoIIxDl
tqxCInvgQv3KY+dGZ7vlOQylnolCLjNLLFRLVmm7fCICoPcQUA1Y6osI6eVg9+fN
hr7C00B0yIoGOe+10w+RpZ77g5YU0IM3LQ0vAiM19+UGJFZTe/zk+MUKNWLphJEb
2ct9gAl4Zd5fLqLjWIbVnv9XGnEb74EP15LldFfDiUxMpTTuJ2BZq9/PQVIYbt/W
Nq8LBbzbb7+sMRIo9vsTkWJi4Po0Z10yd3Q1new3MJbhW5NWLhRo/OPwul9o16WL
i5yvcgpwviw62t38XIfmkiyCFmhR8nDpmBLlK4TMyhmQAfzuv4DZl7t3ItH60YHF
3gj0WlJ/g2crP9G5RObU0izSNNOBA0puQwAqFnB74E2Z+g38idGNjZ2T/QwvQ0Wr
r6aV2F5qxZhKGZmCtmkPvMrOZfNNYtnJreRyksuHSViUh+cIWBpCak/rzA+vtgbA
vjusPHLQ4gjDXq03h1DwE8SBlppzr+Wju/Vk1+hvSJwvqtRN2ODhU1Eu/yw9AfhK
/2i84afCzRdvYliik7GY2QI3OiPMfgByc4OPnaV3ysjau66qH1PbG83OE7/YGRft
alyLaaGAMh0clr99awh/Cy30QBgx55YuaR+mm9o45qHjKlkI+XjOIrsRdgIjNVU6
lvAXQzwGO/E9hdmyAfxCqpQG0W+sv6jkLGjqfXySoFVvFWgaPrPms+CrllfdzIEv
gTU6Voi5wmVfJpWLX6lS/1jq5OT4a8nw3yLR+DD9fQz34YkVbQOu6GryRI4Al6d/
j5WRr2+5t+DkPqUfXWv3ng3H7wrtTQ+QNwCv+Mmd/CoZE1bBLnolbNrhLYaBbCXc
AR516Tsp/7e38X6vqh4YYZp0AVe9focoowfKJFOgYplX1cL1ybi4Zx/zm/7D7Mcu
EsI8ylqXk0bQmVqr5ZKjYxNY4GF8tg7GMPcrulLv6fv6CYswOmByMTzyD3d2Ajd8
ETe24FPffeuAfdhe6YIUlG5isWOWk+Cy4bJvlRWEqDzs7twPziHuncZe3CloDfWg
ePa1a0DRBrJkaay9RCtdcw5J6JiVjpEZyqBETcwfBLXpAQW5yNdOVyY3V9oEbrPF
scT+pwJoCx6JHXr/UHDd0rJ+RRsGN5YIWZRxIvpchls390Wl3CQTE2HlhafjeHJr
ZUZ5evjNHTkZzCxvxo8oqafi2WhYPLj3JWyIbxKt5RdVON8vy+VNLDFIV5sNW9yn
+h+KipRHz+KFqmyVhqQ1iLfHbYkpvZXBfRPkvVhuJBa2k9AAppfLKsBg9mVuKm05
TnA/4zsYWnY/m6r6RlSIE7tR8EoinLfUDrdVMq27I5P3mhcAzYgiFczclQEsbaUS
dMIjWFS40KKsikMA2eT6vaz5ImjBGvZzB+wiMBZe+elcO6sKZebCBLn6OpwRXI/G
6lv1k3vK4MyeCAeJ95CQJo849+DkB2dwVuFAebhimrf+PRh34DFofWILuFzWrvd/
Oy4OGKozwkqx8n/qGF5ZWG/RSm58T5Ow31PAu7x+l1yGFfp7NZ7f8mI9dDbmpMqX
F9xvUZjIut5l3S2CcFjw/67jTf9QzEVbzBUzT6J3BMgOwUhiYf0ESDdA8ggUWM11
iGMsDTRvhaPEkBXlc0rNojVt9jZK6A8rMk9g2o5KrKaon+1dIuvJojBpwKriVegW
SrTmd1lrO+IlIWIEg8Dv75IGdexCn2YzUoaKWsxfp0EHz1LX8FTyD+asZXG+bp4N
B2DKmqAODPMrtY+RT2OTYbY0iKHZVY7cM4oEiCmvm1EKR7QRHfca+YTtBg4bDEy3
4bfLL2u0Cprv3M8Ag/GhRCityU3q/CFVZOol5V+OAtmvCvtxGwPeuZQyBCLU22Ee
PoW57X6pM1jpf4cYEB/BLP9uke1gs/9Ui43F7j+wt7Z4m7ar3sk19PXScQzZBR+Y
Se/XuFqzjoMAE4hV8Yml0y0fM1n6wkVwnSuK7K8ToKhSuF+tgd3CWV9yfGkbUSEl
KRjmw0uLVKag4i5tJ/W0NFoM5v1K7NX5NbEaBg6nBQwtTbT0atfoQo39htvMaM5m
Pciv3JU/PrbE+aPjropUoNBTzBfRP70oFVRx8Aasb6IQ5E9t34igVN96Sq3udo+y
7uA1UZif3oH2DB+XhWm4q4rKUvNwW+7iUaP296tbxXoIcN+HeSJNONqxv3QIts5P
d0jHFchFGt46RdtOYP1LW2idpoUCTjS7HZszpeTNfv5ak0J91ipoZ/bQ/eD5HpBu
rkoMIfW+KYYl3XGkumAKNFhnBjsgoftkq8qYHNRXm2vZDbL0dlYBVWoUSirlvDI7
MtaHezeCOOvFqgV43lBJSYFpfBbIIiRoNVmO/KweBxgQ8EeDhbvQanZOGK4Jn8Kk
8JQT/D8hF95sCDpq4UE3YXfenIq/mZuL7nYy0YWNPMYbRv9OKoSh5rFrFeha5Icy
zgdfHyCQfzj1AheyA5GMlJYQrNWKQacMCvlLLD1d7CrbORDRHeWqFop97ixGSGRR
2I7Df/xh+1slbjF+j5i9OCPKBS935/7O0GZ0vt0j/xny6xjFdxS9hbs4mOErYGrm
5j/E2ZsS759ov65TKsaewEGZL3h7qaoS+oG2KinEbEGhSGv4pwiHGoL/aM7BXg6x
VE2pTCmTuZmphRGghFz6FOXPU40xY95wmY7YQKHPPyEgjZEu+/+KlzvlzCabXilY
aqx0z2+LAk2d96eua2XTng==
`protect END_PROTECTED
