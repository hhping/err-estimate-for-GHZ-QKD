`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjsSyszPYqcDdseRlAnaV+DNJVzMFB4/mQJCIYZF0seUsvmuxxeX//RmYZ6if4gj
3ednLS0j5cjkC1GsZAPCg2Qkzpv4BNXTy+JbTSg9/Euld0O9Uc2OLItphMeAkOud
fLeCDVdK51qEFzF8DoztSKO4IMgrKV9c9DMhJ3Hw6K2N1Hr+9/pnt5RiTD+ZXUel
ua06QGIRdQp8j+MzaDXQ+zXo4JZUqdSN7letlUu8vxCc6IwciYHzgfbmAf4dfVOb
ELO+nUyQVcG2QqRJMNBY1v40EZOyKFJHT1F3U1BvJRWal0B9alicGOrOIwxr/l4p
8CeDhUHcmYYaZ468Z9bDr10klGGmzUVzIaJaTeTm3eijvnhlBKnOPxF6ogg8hWJA
1/sDu/Bxe3BUP2jzk+V2DpFatPxrt8vAWXMyCPoLtKuh1z07w331JqHQLWUtOjuU
/QuViSKBkkgEsc0HFU3nFGNavm3F0RwyjS1bTTuatWFix71uwQRauF0iV+ZWmKs1
wOo+obkDV9JEBRwb4StjxI2/a7JwLniVmYfFvxdS4ZFj1RaZyZ5sLOIVezAr5pZ4
zh6tnpY3mHyXVBHB/m0QsKUwF4SQDruNt3xhaEzpByx6/x6I7miqDCDsFyYOg6Bb
a9wZ7/hJGU0rdm7t8yB0p6L/7NiMgewfLYpgYzIxnLnD161dI19wZDoquEJjR8Eo
ZfA/tL2Tf9MrA7uSHsF0qxIglbGMTefcJVUIpYQuEY4GVe+y3dyTrMyt1IZG12Mi
9nxkcswJw7/wUAuVXbIrSl+e9PEWLbxsQ9bfl0wQ0EbDwcQCWwJtM9ujRaso4hWv
KlVoUvh9fQOt0KPFReI1duVpvx6bbS99tdlvPt/pLOEL3Lr4G9e5sqXRSlPWZk3E
tarMTCSE/P9fbwso0FIm8s0uoC0lYFtOvYAZ4gKsa9D9BLNnmUnivjyODAsFh0tf
rcdmfC7WuppE0WokhgE+RCGQuJxccEnYJEtA535mVoGDSeguYhTuuzdjJ9oT+6KF
ehAg8L5+CDmgQ0EVmfLfVOXgF8EV3XibdB7uChwR88V7/9FQ5BcZX8M0Uqm4Ld4M
NFdbojvLBvZw0NX7fuR0mXaTFpPeJ/ZaoRDZJx+cM5eMIOn7TEyEIKupJqtCpQgV
rNJGiKlyvR2C28gv1YzZF8buVXSvXhOUqA7eiW7a3XwImHVkilInc7uf9OYsTau8
/jq5zhTJ4m1dy7ukvJh3a/SwIACvc2UZrIDq0NnanIJSKlFdQHqVfOn5N8EYCvDw
dB3GdN0SH8tRdBEBFEhidyfx010nIEDnGZdP4GlBo9uzC/K4Fn5fS9eZQ/rsIHwo
sOSkgq+kE9F7hiX0Bg1KWYTnLycgpajS/9ylvcYTsKYes+cyFwoGGnVj5zu+HO2h
bnEdkKteB7+S4UTSZZ2vM6wcJte9y9zUsD8dfMqjIr0gw5G81qIQ7chf2+BapRIR
abseukUrkChscfaIuG1pr8Zxw4qvrNz/c7BmE1SqctpaTTb60qsBgc+tGO/m1SP9
ljay2DG6h4Um6D4eQh6LF3oweQkD5cCguBiwF+CZO3bLyj8bhCr/4KNlKAtQu4Il
0wDwwVM4jVy8eOjzbw2agm3Pok6Z59b4Ur3TEItxOQnLVWgZHLxcwLEhmruav4Pn
vL2HEK+DX+Kq/7hnZ7KSRPpyV4oKuIt6hTayPeKOGg+GhM39JVWAYtHwU7oAnjcD
reoexgx1t+y/vKnLhURTyX6IMGc/7Q5W7036Wz38KA80OGCo6hdGu4NL3mk+BCr9
70aCH9hKC13cL4mJNPy/bA6jIG+x65EgGmuRqVhafZpoiUyZGMPDuMGj5owXB+mj
u6UVHdwMmwVKH7J6fGVAQ4HompzYEQEtTkIyUUBdTvaDrYQM9C6sHDhGyka2nblN
z2qX3xImcHhvJxlK2b4OfA+osao3/3ZmlBt7WrVpJndf9fV1tJInFKKIvdcHHK17
`protect END_PROTECTED
