`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mn4CjAssGAb+Zd8ZJeYtJ0mmaHWmvB1EFDWasuOabQsWGMvYN7rj0lvJD5obSJsQ
OmHX+URgh9GAOob4/WH0Hzc5ms0Z9BIqLMNTu65giidIoY8fxkQKts7W+L2q5eQB
+b88rRc0WoZ4J5VU5lrcSEHZIfJ6sugGzLQReyzWNtcekC50UIYxs7Wz1WdiZIgT
CqkRCCIiaxDNsOExUswoX8atOrTxCY9wOoce0D9jz5dkbVQRjk1zVA/1PqKvJgdO
vpIgTDnqAYSbwLyS7Uea0gBZEiqRMUuXeI4KlAe0xlsVJe8B/+OGr8b4pwUNxADF
/PXLZunwF0EWsht4d2N3KPgv+ZLPKpx4NeT0R+IEoMolWrvTAgfx+/V4frHCcvPt
SXk0R+6mWvUdezGgV0A7u75s2aIKU5Cr2mgK99gOuMtygjVrkWSdA1BActBX6iu0
nr4FabEDifRo3N5FsuVux6BOwAuJx2Pt/K0TsHiLElvoRpyT8sMtDPTN5VgYoXoc
+61mpmqj+ReZT9WE1HKXHhzT/siHy3+CgXNwB/IugHqqQGQUGalUi7trWU8tEK+g
r4OFS40gH7W5SBLTpdvXrDuxG1wML/Nj7QAVycdTiYyqcnsHX7rmJXjydc+XP4jc
9qomqHuMMstFOVsTFdtsKYuGd2N6mQ2i2Fvls9kWDaE=
`protect END_PROTECTED
