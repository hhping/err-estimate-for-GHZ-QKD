`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQpNJcYSJ62iEv3QA1wfUyunVV8cJtoPgTjvvCHDNp8iGCKO8ZIYO9Tc6eZDzEcE
zS460SeI+lub9RhjpQZ4UCAxBPRrqWJvgB/s+p4a8JkLPM2rCBm1j8Kdpgln6ljX
i90KB7Sco3iqPuNzGBtM9Ua3csZSlTdF461pXA6S7SW6mKSG4THOGdfmTJ7I4cje
jVaF+7tuC0cP+3NsSlfqYJew/wbdkI/B05/bcjRPFuzxzRF2q4xdywL0pVqoF76d
84/DL3YbeGEOGb+1yoSiPsO5tAsUFtkWQHLhpNf9GUYobreeZDdK+6Ir83z6B4pO
pfsbeqZ62lMdtEoLoqf7+Va4yWlR8nLobSCoBnk7txOXVSAJOK9uDtJqtw0rZMXJ
12oKNXt7KxDBgY9SoeKwoo4lkfBQJpnJgKQN3hERhnkh//e/mzu2iOctTTdU4Cx5
0KvNaShNzzYbmnVS5HCU3UfxtKpEasbtY1JmBS1ctaY10IvYIn4e3b+pEReGA6H/
TJuskap3Ndy+/7DcBsrzN9OBso+tJltzLAM9m7tb2fhpu9wd3uOss5JHN5+5NCe4
AZQNUI1B1x8678THzhRaZ4oj6M+YcH6Zf+9OL3j9rx+SSycAtL0vSbVC8U7wX1oM
CzNiitKn9eFpzxPU6/Gvpa4hqnQHKxxtjKAPgdaDKOF/vvnkiOwIjs9b//Y7v6jo
udS6Gqf2sm4dTW4p4A7JtxfVGeJ5ml9tyIRnrUFwBz2WvA6pfd0+E+XRP+RvUOxh
NIzsYokwYGi0QhiACmxccnKvH4YLkAh9nFyh/kYH9vijpD3INm0d9g/HqhIvt8eJ
fZLasNh9P2exSkL7TKMbocEOLQGjTc01XfaqsaxVaaY9fmVOXGQ0vDwxHsKzCnLS
Q9IC/YX0AMvnnqMBDexCRR1NWlIG71YczhDlJIXSfF5WcXhEGN6GJV09VbUTHa2d
2h2z4pGagdLBEXJCZZwlq0nSzOBCHDRVFBE7lY0VbsA5feIslTWGJ+X+JsM0Mrnb
JSqoHLkiFeSau2rBLGS2akm98Vzu1qIJO0trkA7VA9qLG7Ye0ksoV5QNg2TsAUZl
MQuxyRoCrhreneOA7jutzAoz8aYxI9lbBL5gpq6mqZ4CveJx7sjs3bdwxXlCwW5D
aJb4flw/GBMPI0dpMHQq3BXSoRc9fa4/VYj+DHCWBEdRRFk01MPw+GfTXzL1UJCA
JhaSmGie6/CyQE6LanesBOgYowqVcRYdMSAmEZxU5dva0lGCPcxWWpjeVLnlgPHe
pWUtzVJRD1opStSD9JROlbRCH1WFVx9jJMG3EPFk0l8GGSLd4Dza+vvjPgqN6yRG
ES8kcfPCd++BGmoYWeOXD85Oex3dXcHQTedvkh407TPO5wkpztQkdvSOsmtRmGqT
a9vW8i5mwBayXGZjtIDg5dcbpSqs3DouPX3qNEZzCCk0sA6oMeS5g52XuumhAhg1
1y6Y1eRpz5RHbsuSycDoYeHjCRUFkdLovKnfSmvlsDAjidyXtwGc5xyq/NlXONzY
fFdYc8VhjwVw+4zMX4SsB+x++NklZ9BV0DONcX8M+gyOuVkdsUHREmOgkf3MXQJJ
vUdr54X4Xcp64lH4In1nxobPYmogdyScsPAXBfZeHkvcYGbDlNkzwHoLxyzWd5cN
mF0CsNj6ixE3OOrYVRpyneYx9uoaKnjgl+tNzg0ieSbgYgaMQkUU4t57fvCaUZr4
bpqLCalfID2GHHuLkiYrqDGx0GFqNI+nrpYwdXJ4dO4KsI+59h8m6EuKlOCtvy2n
9EPUbCgwS9tHfbEiuESlumGy+d6AeCPy/ZUCv6eMUpWgNPCbBAd8ajgeMyuShMeQ
a8t3r5mFLN4BO3AKUoUjXkmL5Pp6XWDXdc6lWUetQvcfgmTEEkkodcXYJpnGCLm9
pHR0kRZWOEpyyTLZhoO1uy8evbqn/9NvaQL88Dr+8b2p4ZeNzaOX4QD4d4xWrKdi
12LOCaqEk0jDTmdq8zc3KMI/9pPO33n9RBK03WpinmKxGQ7d+EvvH5GkA253qjU7
I0CPFjC00gOi3VoyVU9Yqg7doZ8fAfaupCbksAc7ukfh1h3vgWZCCa52EuNMmNh1
wGtD6qnSg8WHSKRln8gM9Q/LHdhqQ0lLDiBXJM6uB8nHQSu+6oeJfNOR9b1Dakn+
G4Qf+fSSWbdLO9bpLqK3NQcMq2Tb36oOui9Y93ntsZmnIjFxk4GtEmxuuLMxOvx9
+pbhXfQQhQ/z0FXVxhNEXn2+qEip71xBm2XwZ6Jlyuo1GtAqk7hc3sIPZiIZhY8k
zx9FebFzbdrBVgo8Vft9EOYIQQ6LVhd3nR1A6GoZPeWUej9wz7riEVl3hpyZrWf6
ljM7z9jHKKIQk1YrEhBFu7K200RcVDwNkacdepo216xfhmD3Wjz81/qa0OoS8cB3
MJYZHr7ZUPpIFYfeKK8uaHle7HsmQZGffhCggNSrXrbfoGSTRuZuUIuw3lbjBfEJ
bOKkaxWgD5B27CYCMFAHAbsCZOIzK9WprJFgKQECLfIEDzH2Appz3RdNq0SmNGUr
jBzOsCKFUXR1Pplb9RlmQB2kYTqDUo9Mb/xMqNh0I+twDXP6RbFXgMFYHGJ2dHay
CXqPTwDiQhOrzqd6QhODoDO7zVuX/DRMF7CrftBsQijpUrlTSQFN52/3FVfaRK2w
L1xmz0HVMkqrZOZnIkts3NVmVQBoeZ6/IxRXNQhw0YYEvCHNvJc4ycIU83/vPz5z
mxVRv53ZK0UNbNsY88ZtEoOrbWbNS9ZN69m2Xt/P/YZQz/ja3N8RyiEkd+tbt+E3
iNf51Ilpj1w74BfdWptm+K2l/6mxk91iEOMMj5++8DYswMdDdWaA0fhPa2ihEPYp
nLL1zJDn1hum7409GgP1ZvqMCtyhu6ga9AVEzl+qutM=
`protect END_PROTECTED
