`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSTfuGm8cC487US+3eRiFVnsZUzZB5J9sZbYNqKo2g2ylaCdh7rjWF1mohcOeqki
gALk+yVWkTQgZyq/bLMk5ipE/9mT2XmEGtSm+G9oHPMFCKljD+Mrkl1Xs4Sjppqx
tcwxYgOPY98OPW3CJaogS7Olye1dAAr3HbHHZKI088+yPmYsr4WXDnd/kBXalJmn
J5DHviHNnK1HJ9ymu/m+8ldMcc7SjAPbTVOGMI09FyUXcPqOlyoGp36iWZ5Bou9K
l6AwDXe/f7OOdXZWPQFwwPFF0XsGN/vUXms3CYy74P54gV+MqSXYEYV8/LsJ6tID
8uLjxczxK59Xr+JKF0eakSnmzkECa4bNfC84+fY0N+QjtvKvbyY3lRSMg0cMGMJ0
S0+GHXTg+iGvwPn2ppFWv67Wh1hpAau85uX41Z0Xlxm8YObo4/Z7d9DEzbVp6cOS
1hNak3B04YcRCGL5Qo0Q4Ul5KOlxmae6J4DZPGX+sHxJx8XfiKcLOyB3hxLsk8qu
UCH2IL2tpf7WX/sKbV+MZWORVTXYP0a5sBcuXYrfScB1lmH4eGg/vLKJErOB+9LB
IoYtl0ykS6THQ9bgxD9IGykIOlvq+uhoJ8z7woeZtxn0/Kwa261MO33oZlZphyS0
ScPf5IT3HgNOAEjlQ7Cks4GSDFFX9N6xbLrTJjeykscBYsOp8HH6VIW3E6XAIofU
EJu8s3SV3O3sX4B0hMSA0C5ohF1kjAtbKHfQuPWnSF47pUUKXGo3/21i5O8VWSJA
`protect END_PROTECTED
