`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SgK2OT6ghxdZvpkZT8kcAKgqGWcP21P42MzM4hdb03BNFlgeaPAM9Um7fH5yNNF8
f3ljdIyMqwOpfo7qX59eEr2OGXxBBp8VEAeZY5D1P9hCOxfdoBBx98UrtEkQLd0C
n7olwq+KA86xO2l7Sym2wrqNMlLuVUwh3RqFVggiqtTRQGwlEGgKb05wz2FK/9zV
GZjZuX7dm7hWbqc6WO04PGF4cU3/P2smfRK9ndAPZ3UNUBkOWvrpAYcVk4MARQ9T
6SJZsFXoQQhFb6RnZT37xdG+svmSPynjst+axE8Wb5APWVVNctwd3GJXjUqbo+O8
ljGGuRs406cRcEqofKqzC80x69k8xTi+8SHSCxpG5xRLwWg4m5qA3tGfvpOBAQUd
UftQho1d3ho8HNIzvYMVAYIHNvXkGzKfSLQFmDZs+S1j0jIx+HY9N4Jv4UpMsSg4
0EHM1yVtW6h69gwYtso/g+Wq+dtQuPY6g+0K/tvzm1XkzV4ZWsuozxFdZSCcF5O8
yS8VQJ9qhFHVlZpY9ObyikGjm8CddzJ//752axBjggtqgyfVmaEtoPQPJdkf5jRY
oU4ydZHjM84wDlB9P32o1IOqi3Ep6L3LJK4p/8VPPlGUqcSoK3f+h+EQnUXfNZRW
4UlK9AoDmpMs10XW4DXE0MVRO8SU/SFwmebJ97+rA9NXNDzp6K7+lVtfivSdbefd
xRr1bnKiIZZ6NBVF//XdtNdy4CPduKYIU2afBNnRQpgTj9H7b6krveMbKjVAvfsZ
CNp3/hO2CMHntPYynees+nFG7uZ+/DYWoX5HARXk5aIM44GwptB9JPE5KTYV9iKx
O32N41ldU+S1I+nG/ST3ERKnz6+M0XuO88yrh5sPpDvXrawNbxco2pL932s92Vxg
ERNkt2uowP4aJk19K+fqBXk4T+D7D9t3HUfOg4cwdbuHbs6rXfr6y6MlqjkBUD5x
q40hq8uKmZOgpTOzwCUlNMEnBXx9tkTIv8MOG0DDJaA4PeCUwYAPR8LB5KON5Gpi
VSo1pedotxJ4qonDgj8ksuRRwwf5KyRb27TB42egALfGT6yi1tTWqVcIQxftA4FT
QA8bVQEQ8capGOjCGZlmPuYNeFgok9kAYmLuSLtv6JU7RejppdsUW6HZgu0W6Weo
tqybbR07SjmpAzfnrfUMyzPHZTFwGZaePRloREkpcEXrivXXbO3exG5wX/+j679n
Jbg9KRLL785O3zHbNB515VnvJOJqROwTlRW4yD5JBN/Qxnw7DcpKnem9hLg0ue51
8Q2rJzcddXMjLyxSNU42qdpVXB/Oe8A51Zlu3E+ikeEW3RVhDsFwt5I6sQRiE2iM
rifJ9GzHZXv6K+MYv2za0XYMuVlCNuARl5d6EpSPcDOmW0+8IxEQxr114qL5Aqsx
mdgWG1o5RRGtgZetdGcnyuSOtZe21N5OnAQBVxTjM7o6BKUGFhRmSFoyOryI8BJ8
rAejc30KGQtfjcE2EpOmQ+wNmNDtdyEdZVxhQpgWbQgQzmUyeFcnp1a4eifMHELp
v9yhT3o7bKKQKZH3X+4Or1R9qCAlXVwhSUeg2Vm6ZYYyV8OVQ4C2xLCexFT7oUbK
vsuKBejuairgVghQ6qSoRXCUCOJktHRztKP9OUzTx8UK+AkyE/EizOjj/b9Jsvh3
E5iz5xuGCdeV1NrbcogBYzCn/efWZzPZmnYMqj0Na6vtGAc6t2FN54y0NPPLvEf+
SoY2dFaCM2dgvobVDURATAdONHqD4mmRzkKDhRKls1hA0cOeWF3C3iLy5tIMRhih
zKBZi5GAJRiRSZyjg3xvdNo9wSNjJT1aqN6g5zfxbrWbXPlLQzfU3bTrQ7i+xb2d
HjMQEbPuFjzlh4qgIfSvT1oA05EDt/ourR+MiB541Wl6PHFYSmMV4dEHme5rhPho
Do9wPiOVxgULi+uKiAQ62Y2Os8IveUTjS/E+4XYtWBxneEoIrUm6+yZstnzG4az3
`protect END_PROTECTED
