`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1UhYwDlhkad0VdEEj4N1lp6yAR3cGUHt7Ee48FzEaW0voNXLzN9CeBoP8FaHenIV
q/q/KqRuaiuVHlL4kqnI7QQo9ZXyndAbm12f8sOeISKiBHHw49OZplVFYxKfgn6W
7j8MXhvSSv87quz+q4lTFZXrbc90dysxSbZCbwI9ccMAh4nBg2oSO/LLdbDT3S57
aZHFQgX5+yMDPlHsVkvecPbuL1dyhfSM39zGq5C6mUqAwWCqptwWE9OM+QluY5tq
QvcqAA6ylw1XtyIbJsMQs8XkcWyxHFj6wmPWrIPoxhHt5TvoosBBoT1GVnxdR9N8
XGeP345BBi2pempYFAOHyWvjOCmoYKpayXar19ppDMyI+RFyLpO+M+cJ0YHJYfRX
S2dMbOJNlUxdecdF0JW6RUEBPXV7i965dJqBcIWDRLp+C1NoT+dC6JG6lfXiqBe3
uLFbtxw90wXzbnMhNc/HspWhSh0AHUxsE7Mb0AknAdX3jX0s4DG5XgjM8DAFVIhq
1QLm4ErrUzSd9tlDAIGKz+iUXp+grM1/a5bcmJeJS+Vx5oswZUf2YFSWJkNr5zdp
kKlb1g4QSd4Yj9JHxokw+fc3Reo9OvSe2T5td9vvpBYPH9ryWeidQRJrZqcUNr6Q
PfYS017OFVCGMH4UnfhxUTyTpTwNWCkkkowdqma2Ad3kPCnBdN5Gkex6OFpwCoDf
djpGcQdxhtnIfop4dGOwJhxTibQY3gaephkSY0wsqK/y9K8g0dVcLoxfjpCm7SGq
DN7cIJdgvcKBJA9fBjcjHOs2cEiM9OlABf9VPLlOe5vpD3xGPO1kUDFc/+t+Er2z
9flKlcWAs7chzMPJOjkxhgNpKtmpS8+dpgkIeX6cpGva4WHwVJv2Tc9RtJCigYjc
etOXdYJ3os0mbK0G0uXSyawm49gSYTx4zVIdU6JfnKaivP7vqFDNccpPsFv4WhbZ
3/D3PxxSfZkdc9eZxx9qy+IachKmhfbWN3UH7WllGb9nZ+EyZW7EguzJoKTAARhX
dpPGLVUfnEg9YREo8o8YIRBheKDfLeXLhswlmEcqSWdhbRnT4aSWscdrLNkV7aSK
kaEOsMkT5f/teCusVDA30SqPlM3IHQTDYOtArS9gv7T+n2K9UDjbC5kjNg03x2QM
ZQV0rdOdY15RnHyBgqlbbbdhnOx1qcSoQ1yBjeN7ml0eq4rATY/F0bahe1uO8hSc
9JmIuGTm8Ib2ZidSX/2vsDepAOQNpkInrvJPJRxDLXEC/NGKsSjiXVHgnZgawqCP
`protect END_PROTECTED
