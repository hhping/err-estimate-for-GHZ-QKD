`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U41z0CeYy7iq7KhEN82fRJ32Y4YKBGnNkOGo7Ct0iJe5a9YOxc0+DR5Sdu4nbuRL
bpA7vk8QDS7TBTGc3xmI/d6OhDCd4BMypHfl6Z5nGQyk+WNO2XeS1A7IfmQCKBzY
Oisbt4lEiC/iMeXQgAcossbgE8YcsGwugaPuc52Hh8kqv6JXY0zkU2mez7ykKV9X
bGQJkpyfAcHz5mnEsd9wdbAFIb/Im2Ufuf47lIf1skCo2cfxPtfvGH6rlQu4DnVO
1ZMneC2SvGwgN1wqCoM/RG2GWxs32JQdFBoLl7fxWuwR8ooPsDnOOxYv4/w5bl3S
ovqXVXH/fE2dUdCRdtAVqmaHFiKzD/yrSxk1m5fnAHnQYsavjzpLDvtCzjBTWeN7
n4oUWqVxIFcIu53aDrJ8KrCsUW6pE5pn5mn/X53gPGoroPIlnZcAG8KA/hi9hUPH
fUn6rsNwMrUAh6WDQsWi6teaAtpw5CR4MOw4ADqZchUI7fKyq3fKcaLXHXhD7Z2O
23Q6hrOm0QhRsUry8ZHBt0PB1hoZ84IC/9MIC/7an/iWa9WN1GNandhzSGGwR2eY
ZR4vszkLkOW7HeWRHCwq+QvLgICQw0YiIEo9oPVebeCMV6zmUMOjmqZjF+3qmQ15
R5vSe8ltAU0FwjKApX5qJ4wwU+6L59p/GfQ8aWhhp4HrMYTe8lHo8J330KWcg8+e
uKVrlpSxLT5YCRBh2/kVf6SZDCYNA0ZC6LW3wPYv/LHoYdMpYim4vJrA/boAFHFZ
c7DnERsvSeQGE/24MwSTQbuXR8AvA2onMvwZvn6NRUzX61yXD5vsTNJ3JE/9hwY/
o9jzyota93h4AtCBqjzyTcpMpeftJohZRdK8OJdl8sMOO+2sgw5X49+EOXieJMms
FhV0LfJm2zsXTHpZoDlm1suTdP4E22HbbZkzVQCqySh3Hh2VaVU40ZmfUbRx6B9+
dq9w4sywCgz6WP4qi/Bf/ZFF63chYtnuKRYjSPMMxynqv/1SULN0ehxquLOGr9ic
2WFs0mPjoJKWtxcSEpKcrIcoqpmMV4+Ul8aVNS1bqbsfZhNdGZ1i3vMbkSCWDwrO
Wk8n1fNb5nxGEH+jcioyJ93+Dpwsa9tZ3tr+WbvVuC9sHiffyHMyQXScAGSNrgU3
p5lDNv6IXw0mxzMGtQ1Bok2HPJLK+eFZQdbuoDWdqz2HI24gUXCV6JoQsXFm12G2
L/m6vnCjbRELU7UHkvE1qf+ybJmGXS0ur9MbsGoPGVZdHWfM4z4ttaBACYL+ZFik
T5HA0Hgr9QQ78EkR3ej2C4m2Njx7/7Fjnw+d78VzLeaz/aum6hpwB2ShvUtXZo9m
3mEAryDgbA2mn9r86eKJRdhXbJhhOEJql6p2hAFSWckwDOeQdDp3naDrDY7jZOjX
9wIviwOPdstl4qOdqqRyhnXwONhuVWG4HwoyHkkRBiLJYxmaJ04AdsBZgFdfXMsJ
ezutdBN/EeXRVAEG2Mli+8dZ4uKyh1XUvH4WL0/UvBW6pQaD7xQAh7gtJLecPb1p
Kizmu/CvqMo/4fwOA5v3UEm8XTGUJahSBke/hTn+HR4R029DzWh0tEJAoSXgRYvj
P6J7xC6H1AGy3BFmQfrFjJ56M7oVKx3X1wPOoNPRLvaVlzkT7a21F2QPZRxazKZI
X+fBgat27fKOxXtR/uf0YH7VWLnyYkhGfI2d2blbRUWpDQt2I2xIE56zf9sCiLUU
XpSHvZS6Hg36oWKgJNAAYQTg4SoUmscyeqi7LvXQzBjMBzoApTYb1ycFBBc/wBDZ
BtdQDBS4oQA168cIms9rbeWyu8zzy7rz0K6QUXYv00xUJbEmd8rznDHs4n/j498V
3NkmGd1kG0K3iIWu+yareD3h3lep6XG9WnqUMjr2TiSKamHAksn5kDqaSD1Vdf1o
6RlZa3kAG9pwpID4rYkFat+3/ntY29h1uqGqqw8S0yoR4qqklaBuYw90olIpqVzY
J2T7M14tOierxFAJ4RswDNCTAr1bjyib4+M6htLCnHD6i5nA1MqoHhKOllL1zCSg
nqqpa4/7swOKMhMKmOwK5Mct3A3IQR0J5KPE/WbO1AVYS7W9CNqA7/vUwW1YRJHw
zpx/24QjLUmTSx6vfu3sIQkmEEUEnF2A2YAIAppklXPyJkF2QZcdpLqwh8KtHRao
sS7Swq3kFECdBK+/RaKViKaNNMESXHBYQKp+QWGiSSzGYFBVvg+NRy3gMCFahtlU
gR/TRIfT4icINHvDUAa+Q8fo2gao2GuRA1kATqE3iyaHosjsQwIbrmVH3m2OS88G
PGO6sDsqOdks3Caf5LVPOGPWxgenKk+2URlfRc/xH1Bt4RwKxJTD8w4rGbum3LBZ
Y4k5dBUgX7vBWRqqXhIGAQU/mVZJGlRrFp91c4+r0MJJf59T3A3Z3b1NV0lvNeZ6
8fG3rmZBTktCS2nJwBjhLoOr0ZzGQRTEvUTVjexJhBHWslIvuLhkVBoFCoP6zlsD
fRQ7sUWLl8fP3gbLB0eYSS4grSIY+7GYo36rm4NYEAH/ZsloR+CX/0verjsU45BF
6j1LqLYvh1Sg9aP2ALEHjN6iBatWo9ko4mL3lxQBYinUslVqZyTWRqlUrhthWWLr
C1UZqOfxu5eHdHRruWz1u+seO54ytYmJueOFeTcQeQMHstEYYAxyParIadWyhp0/
t/TpadTqQRIzoPeF/+Gi59LAPpquq3HvflEEO33zPAdffu257wWGfRMds72ovbml
WZLekt+qQjiL9Ak/RI08yvT5LH/snaOQEziB9VGBFXJylRRyJyIAOntsmZrF+dBr
jN/MKXSjy/zS9LbXFti7oeOAcypPH2wLL5yP5NAw7xywNukoIAMkqsmfMCyPsLUa
u4QfNxtonFFPNiGCdUcuSIWjRByrwlJSY3QUoyJSxGZQOIkSCGCF04NVOAH7bOlZ
uNPR+gmevp3peCAAytYvhiBnoUKgPz1VfljvFoZNhNiOO3Hdqb4wUlrjYFRSTlUI
5aacmcZ+gm8T7JwYZQm18ruz4xqVxjWDBdG6jUtk0fjrHlL+bsF4B7V47/RWwxV/
IOduqw1ZBQcbYNn/6Lvx7TyoDvbheMHren8wX+72Pejz7n3y6eSm/BR7V8BO8ANE
GAR7w9sqBFq+vu/7JNU3hcs5F9e6K0zDpbt7XP9HcYLMaX3gXv6/EhnYuW0yBtJr
GE3/ZnRjPsNpIPg01lxzWLwt7sfnSQJDERb4fG1ODlDZXeoAB8xrtCxVqrpf09M0
yPAa+BnothHXSNseZukE+3hzNbpzCWkcciut3hZGsQy1X2TQ3aARTOOZhgglK45J
0srtvGM1J+QB/q+eS8Jh7vc02fYN9C6rmwUP/uQnHMH933hef4MUOfWsFVTiE71a
O58yWGtDuHEW2wHuVS7H0FFZ30xic04gAC6vKPh2zKyDoPRQoiHgT2xZnJEmCqXI
U3Bgy8PoTKerF/V08/R761sho8+LqfAZG6Rp9yljdbrxNKI8iP1p+VSovKCDKnnX
ZfSlDa1eiZgJQkOCGEb5RNt+33vu8eO1XxO3M/x9PyyckN2rQB4uMfeaLaCMJ12y
l8F2lmq6mPsLGyVEakbL7jk4mkIhnwidT6Eqi8zUP4YdhEXFcbXqkv7hXZBGbC3u
H7t7u1vZRfu3jqOrnVdZFWuPxcX75kd94/a084s6/xu8CQ3rHCyESDQSgWlGMd3u
Am7ySApZpUnUvKJWbDi/r9QE1eFhfKgFVv7m6H+slejELjf/iCFigoNmxlV6M5nI
yXXW6ZqOk/fVaohlCLBXCI7RD1MJPmq6QeMv94iUKYEivP5y3BJSb6COtsiNkh8P
LEwFajNuwLydNTzESHNl8Q==
`protect END_PROTECTED
