`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UV+DlXAQZcof3Pq6y/wy/7HPBsb/jHgV/hDFnYbFRdUT0OFDPKIgScnI22qfn9Xh
sKoxSyFojkq9zoCMif5mVPeloG+IiIK15OBpgmUIDbyfHetw/EyE37kxWWI/LXHc
+7Sj8tdtIx0coRcMPw4vM9sB+EC7WtoxWBXJFexPxqAlJXMhscvmeL89TVU5zCR+
DqIPXRW2EGdy8nyWIT6/dq+FmhtJ3/PWblhqT0hbSY6Ih0GQDIxY7wfHqjvKJ9lf
f/ZtLrmSyo+h7l3a2ZSMRs+KoNGfsQT5gZe7laJVRmIjZxaEDqdnlgFTSlc85/lg
WOcFnLoyqycxD+nVL92ji8ihQZGKw1kZv7XMPAeMNfL7sB4AEuWr8YNMxvPl+Hh0
MsbLAJgUoYtJwGxLuhehj2pEcStva5gJdMm/Q3csQO6wJcHYyTkB9wCBCHTXbmkh
Z/Alr5gUghQXyNj16hIiTOjlkOjIDtoXcn9jEx/Am+RkmqfRT0eviv/Vgx8l2fT1
ffUMIepgXpEh+wKr4682iueeSXIHOuS8F4Dn6y1cBhUuFioQEjUl4aJ6acMMGybp
tcK2OB3aUWNYYT7NKotQ8InCxkqF2XEKmNRNpOJPSABuHjjXEcc1ETBMbIWMDpQX
T2qFzUdJWSGg076cBWlqMev26O4es8lCmhN0oMvai39L8NJVh4Ly4coXeRuzV9l0
yKVCxYu/vrXFTCuVD06lJnd8ALshHaEaAdlLyObWjeirjj2gD7zPWyXlQPzWJJ0d
oVSyy+oi8T+yoEjh9r1Ij/qwCgev0RErO4mPaezcn0x4FLaZ+iEEEghn3GEPo6CC
y3wIZsirCFKxkX2tOey5yGPhC7cQqM3SM3LaP8osUTyHgJ0wxwHg1ze0YjCT5vlX
1hazOW8EVGc/L9OXHf6K0LVpJmP2f0TT2YHUABlbM3HeV1jclruA87bxocsxW6+f
a5F+HP5Af8JUbNVrcIQZqyKryWS67AMAY7W0A9WKMbbX6wmsW01XfXpdGLIoIbK0
D5U96Fyn6SY9WJec3k+3FZErwMWX2NrseW4SofbdL4IihgNdYKEuYLnjg3N4wJQQ
qo8fFgcv4nZw1MO3wxaSyO0C+XFho+uiJiaB9M8z6zGXzZNZi6UqXpkoeJDpmAzf
g3IBwqRO+pEgyo3d98yZ2TumAhD0nOd4NjYvI+xRmiYFLjLs4Bo66rNzCmAdeKyF
8MxpzIle/tuOKFHYYRPyQJt8IHlw0E9CINNSHX9pQCXSrS31ZWOyx650RNmAfsTD
K4DWCFPwnXOODIqA8PDWS/AI/nYCNyljvZNWdOh8zlYjF+FfhINw3oiYJWT5CEBA
+jVy5VitDv5U+QZ1ygweiGIa7L67ns3aVA9RnLtl8eTV0c/V9EE6h029mnIigVOr
GR/Hs0MpD8KZqzSh72FWPMSPBYXqu4k1t8pZ6sr6PQ7quWBI/hF3lvlWo/2iMQEt
Mg5qSWBy7SzfRQa9eDZy2/IOmS20QZufqehGFMVbyFfojVU47GOiXE0qe3amG9Fm
fFiiyBOPKLVqRdtwE3anZJFISWQPJ4vtVdckXMzXZVnAjPrsT17R88MObc96NNWp
ZcO6iNXzul2gszvLrq3DWzCW0WYbYe08fe63gUYthV4K18BSUjR9OrHxzHc0UalU
ikP3OnL1s4hUWpEZqUsluo6O4o7bF1OA1TnDJKMLzKmfxepzsWf4nw7WW1AWj7x2
cTgbf1Eznm01k+/Jd63MZIhfaVDBz2EF7G5cKuD0XcsRqA6JK/pbJnmnN6xU6Laa
wQg1MJ5ux376CbLeI/DhV6YfdUujHCMdJvpJ6YGRSv+WkexbFrqsg+V26tsej5oG
ELoPRlnPbuTUYrC6kBcYRXLpG2pZtGY7ycC+HQBMpcYjwrf76hii9+OX6UBhhyvK
0aQFjLlp2VIULgZC+ex4h/UIDVTqiWgtfaG2om8bvBSe5qrTyf05AnqZgWlNgZhW
EwOfeS+aYADU0PcOcuTUSZOC0D0NR84Y3PQSJq1lKUsGtwBrhksu3/NZmDVtd+Gh
TTVdEn9Oy2ti1H+udA5q9bLBCiKBXBlkX5ksJ0yfW9JEiVnEDpKFQzG/Irjmwbms
XtGAuVrNBTil9fDNs8kEguSxLVUaNtc47jIX7tkgqKofwdvpfe9Z5VwHVksvwj1z
b8X62cu4Osrq1+kFAafiHB6aqPVNVxdhllTfJGRq7ka/WwIlJEvyOMKVsPR5dZTi
OJhJem8VkCkGhgBMu8VMm7IlrHJDDnhGhfpkLXsJSnOpxdK4JDvu4xMBlOR5hPZq
gUQrD0vNM5phJ793BaI42f/eQKTWP+s1xKZhQAK46HTNZx8OARAcDTh4BlM0uKp/
opgUtkm8o3DlXFoAj2MCK+T4fPiqW3rcURD5QfboDruS3/g7udwxHJXx0gleGaP/
7jkZV8ovbzyfgpQXJhBxTVFNZVAFOxbLZ2VYSTeSnpyMJ0ulH8ntvu0g+CDQzDeD
nbcN8gG7rSxUOXvyL6ig44i4mibV2q/6dJvaJdZAFU9+xXmP60kYNSsN2BhVwLuo
MFIWo8ELSiuOss1x0SzyaWaqJ6pUts8oF2cs39YsNW3Rvad0kBt0W6zr6XO9J7Vx
SaQ73jEyAR35mOnX2GJ7qUHafscKRCoSBMcl1ar/54LHSyDV6d8XbfoplxWE0Frv
vCp4vzHsKvIKU1Jyf489tNyp6tqxAf6pJC7z/FIByZTCyRxU5YOpBS4T+UpL7hFk
EZ6/ynnnTmOlO3y0PL4UILlyW9hzK4NfjVB2nDikGZ/5ohG0aBOzx5DYjxWvuQa8
U6SJ1nEl11kVpm9wdtc8np2VhDyWapPoBlZ3CR7KswjtyknTr7RdgD2BLov+ZN22
RGrTcxEUr4KCQPnm4KkR4dM8LUhDVdDhYk75fynN0g2+lPE0znjB/lNFihr3datk
VW8ti0m+Dc8sNbBYMzeS7u3k1caWgkP24/2H3Nbti+um1Baq3IH79n0toWhNjtJJ
UNWqBbUfi/oIM7+nUzTRivHl9lhkq0uxQ1dwom7e6X/vUnu7/wswS7SZeiu+a/2P
3sLbNwYNziVPCQCeBU/4SYFyUTRgyo8yz04XL8uwKrjHD2L7n7WmKOt60n2gzA0D
/k2/ToWk/yiBjsUc+s9eUdKWdIzryLh9YDUHm3t+/K/CaQyueBeqwg2b5xPe2c4W
qj2cD0jj+rlXOUJFcvPCJU8MYxgQUGMgh2P0wBX2bn3CtS4D1oqs1+WvmzDMeewb
erxMq6nH4PfPq3gSkJ7Zj4oxQCBKRVB8BoVTLuWH02xUh26i32wR84tCwLyqBFnm
t7cQ33RVsjtr+mLOukfZbel3moCTujXxJ1INA+R5oJ4gl3qyORloe+GF0cUPqMRk
VinjE62waqD/5wtSXVDskCLundQZz2CZajxMDl3sGH1vVR5Jn7khbQs3zQJxxJC0
qb9Th4p2EUngjJDLYD4OJRk+culSJNi1dbZVpWjjlbRhLJzf0muIJ434aRU1sQbL
jXduFqN5O5gfn/2I0EumPA5bRVBxvgXliF1pyHlDmmIsJFnSKEIw0niLpxrFkgm9
oOuC0RNdhoaWIQ7HVtLg5ghhpKTC/yEUHylCJ8666JP3CLc84zmdDijk3MeZeoRe
KhhMmXAakVF+rNEOAyrBmVLfhSMGkHAkzx9MngC0pXzB556BzqR5eCFEI7EuVWC8
QTkogPV1hROS6Bye1AN+4gLmW1pDS0B06woOp4CHt7C5KSwggacUIMf4w5ofOcbx
ErE+jgSiWAFo4e7INsdlzIq+iNZj4b80j+0M6yTLNIrA8sw1w8XllTPhqoduNye7
t78XALQCsLt3uumoo9dafkNufnxg0v4l5QVaoOb/EajtO4LuJB2UC398+U9gmfFD
9XNOmyi3gSuqaYAjm6lmgNfVcHXGEV9YklhSOVfmi2Qa+wAAAc6XUaBvOXfF4aPZ
lDTp+9Gi3qY6G4XHA8TWXRKHMfoBr2o3g81xfZyDAp5EnoKaVhYwpcOIhrUWiajz
JUbNJhgM8R0ym3fpzwNfqAvO2NnKU1H3jKzuViv8HDbD/P8i3M3gxuHODROhmZM4
O1HNwDWsVl5RS7mPhIpCRnqM2vtwS+vmruBPz3AQj0tpAvuaJMBUrZUV6BA809TG
TQdIUKnG7c9OAvnAoyokCtwj2oEsZdZvy+5mIjL3HaxAbATde8F2QrcDFiiw9BRt
`protect END_PROTECTED
