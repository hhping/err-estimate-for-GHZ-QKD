`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MEJqiAETBKe7dJh1TYUcKy8fUTteDor0GybVLUrqtF4QlF5293R5hgwbtw2xo/8i
RoPW4VPvRmPWxPxhpyBp6PYU9p4bUVFV2lQ3GdFegUGiLTGu5rDh1QRNqm00N9ER
ee7bgWDvd9H7BnrgdAUVyxkud6aa13hFSIqnaSVctxC5qddgUJWwORAhPpBY7frY
4zT+F3bokuOvxgF1zccBoHCZ0n3juQQr/nxj8vRtMX48xMSryEY9fB7t4dLmcAfC
dzngwjurX3tnCM0r/6BujSxN+fE9oFJAcw+btgO2ZGT3xg84fZ715FAH1Abs44cw
6kEK0v2qgTMwBY11/ur4poMJGxIXzLLrwTDL6/o5FMYKrlUwqgxBQn5CQHiHn+9M
ulGiGfX04eGrOh6du7xkPGNrng4GFCwbVE6f3R//9qmotWGDsnLojLulLFB1/78R
m28R1m/UAfaT5HkAM8bJM7oPFJO80txewLyjiiVykBDCF/tuVHXTLb8fLbdK/gWS
Zd7ofgBpriOIztsit95nUCSV9X29xxOl0RN95WCSUCN6bvk66dsDVGj9wnDG/T1L
vf1G9pup+MVIhEw1EsuFHpBnBgQkTjB70Fua3PmsrwVQ2hQdA3wcMkxbzWNeI6CK
Pg0TONQ9hO6gonp0pEMSFdyDZZGLjmFMHw8BgZfsA8pUiQNJB742ff8jDC9YBlMV
luVovzzq3ykn9j4hFiVV8p5Ehj7PQsXkr9lAdeBHsQsEa5OdJ5Q6xZmSwdlD66H0
AjLGzJ0wZzKWwJ7/NxLknuxTrsoSMF4dVXjRUzfTozD27gHEBjBXKBpQH2qn9k7V
FZr9bnFTGsStaLMDWU6SmL/upud4ZV09ZtwgCA0/r7OmZkwr02/JmfP+aWVW1bXW
U/U0Pzbm+tY7ow89yNwHsHJQH6jB2BeqxY7xDyf/GWaYroRhwk+LAKwH5OAmdUj2
PQ0nBjFnve64Q/g4LOkNOEBeY2hcQ8tf3ikHnx4S86O/dKdC9w8JTX0Lu6X5jp4V
y+nqKLLHBDTQfPFuJsIh9+Q93uVmwoDQdJlCz7qJ5ca0Wk4M1RlLxDeWNk6qB8jn
dSOxS5zA99IevMrVBqXtYrdJJQoT/Ni30wtcr154rXLucjdYJj1B5HWgaOggvX6q
yQtvFQdLeMDJzo5pQxiBkR6esHNQrixVynkVrJAUuP3nFJQhgar1VEFvv1MiG5A3
ZUpyALJw2ij7dFmOuynQIJmotFdbRf7jHlmsfhFRWLXCGQODb/upJ5qC9YnR8osE
UCPFOZfdIzHSI90KcjmmMllkzTg61JhD+lkxOAufbpPZHZ1zMbkGN/KNtcnyOlp0
HqnfgM3nGjTPCPNpTzFrrCLGhY/B6JzYKT9G+yUtsncrH2VEpvu3GWRlAWcK9cDE
gcXbaJ39ceS8YMT/gya6uWe7/B7Ul2sCWh+nPLsg+LyYZUblzObYJCY+u+hrSYa4
fY8+4ErWvT+uUbNvOByPYVuq+KcwzAdNJ8Gq8cukRuMT5O8CAc0aztkzILEHPL6c
E+jrTkRextANsmVwFNMQz4clfhRmDPPMFZfGX1WVgpbBI1xfhGHh8rEh7BOXh1Yz
ZfRmLwZY5IEHc+JhrDHk9NOWK+uN2LEg0cUIT4btlr3kd6iRNmG9kjfJYBSdh8Vr
/dxItkAJ8QnNSag4Cg9kIDWvCJO/VWsyyPlPBmG8zq/AkyEZDMOJ0MZlQ8Kls4ad
stHlK++38g8GwZG6yZOqohbAtekwnI01NFoK2htP8TfcBO1a3rUguTh6uE1Z2rag
uMp/bduMBqoHRPmcU78/qfxpz9FhozNZCdstpDfjoiXF+EHc7XPKjmXMrspMhbxY
DIfP3zUPdegN/Q1DZXW/b7M5bkcEqJyBSBVMgz3WxcW8lOh2yPco3AHSS9f9c+v+
IKq1gSwtFFjEm03GPiSMVUqKpYWzB3kdPBFHFCHi0f0Xdws2VOdO2uRViNzBk5nh
f0WRPmH52HZAXNNtnWuEcqIxkh4wut1bGAdn2hgRKkPze5u4+zIjoEZZHgzBVM2n
9f9GtOkkVKe23gnmDUAopnAClFxsaQ87D4pS43TaBoySSjU9cV1SRvlVzqOABmAN
nmCJeWbjFfPl1LH3aYx2RO2d+NWI1HWfgdQ//VziLTOqeDxToFXG7EopMZfnU22E
r0Kg5OAkChTt7yVKaMQ5owLiGQhv1BXN92IFwyj0I+BuzO9sYxNaxYb/yNQPHprV
Xmrj5CP7rFzPaG35YRgMR3sHgireSF/1DIpUVlDKA4oxGWEVzVmk9OlTVCV3YpJi
zm+u6Hr+/xtshi+w9V9yBfm6menAfAGl+li6Yf4XwcUH2SRhDDDW9CcXOY3GameV
oQNS9KdQerNq+m+hlcCedixjjAgL6us7KQczuyXMpbBVhEPF6DvSoPVWP6mK88ES
a6nW6esny7Wg2WoYWJgE+USE/swr+glK1uHtjokmeCsfDDbvuJEt9IXSFEFifnuJ
nSbhQaQXgCDGuq3S23rbLMNZKP7lc1lMSIoJDlIV7zvlwElwc8+D/TzJkoqdLWtl
spulPVdPCOTkGws8YpIXsoyLgMpapBXIzFAnRnB8+Pymv2qvLrPEGpQOkuNdcVcU
tDizoxSibyTPc6+fhguvfddcshJkwz1T3EKt3+jFLwb+SugjtMdZdnGG0m8qq1bC
hLS3AVZcY5R7PpC/lXt82XEWitVaUhA//MzZpv4nLz7wp8Bmijx9YegKfMUj9MgB
+QrllDL4yiQ2MYwdrsEol3rEQUlA4oYTUP/Ii9hR9kwPTevOoO2LDi+ZxuPvHWbi
3XtDBumO/ff9pnHLRQIiDrC0fbroOAF6T2kLQvGcbICLqnw/2xortlI7GbMV64Kp
qwIyX5Axr8hdJmmi+nygKAlOqfC1WSKDxg50XT4f1VkkvuGc7DYCTkH4hZMoqkIF
AHUYyRdUXTtoY0gFUIxAEPlikKiiRCwZJg818zPr7VOOFSts2yIhZTexEfCS45ii
fBpfbYrtA3ZnRHhwy4ch49fqhQS77d2SvYkYwlBr/AwmD1AIgqadbVAzHgpVYNBF
QG6pUGNeERVSGk6BR24ej7oT9kqMS5HP4oKbxKJ+P4RSQUy+eJWvGpBIel/jTER6
sGEohkE5yRgBJrGonWqkefVNUiPYw9Ce+d7phBtQ+UeWN1kHa0DSkLsMH8NaSEXF
1iKUXow397M+GjU7vz6PfzhO/9Y6qBPcuiGw3r33pCfeK2sC2+9QLlNKmLGv12EQ
8oaTn0JSD8RqEYiodT4yDJWdhgZvhpjUhZAmGePBLhcnOZRNa11hJY4dhxDrhEIN
MuLy3h8Pm7nCrH2/cwhSDVYJmBaqo4CVUaoZNzAgoMzSlcxniju+Wqnolf+8w0T9
BmaxKIdwmCoxWTEQybcWT5+6izjWSNhjmLKqhZGXQnzw5oHBSyyHrZhWaHSWPZZK
7SU4b6w3k/WslboB/SiUZZ0UTZmw7pRT8VvTw/gSMYVGsauD6W+dNKR+ncLeSkhN
bgLtx3rVKyDMGHgeh7UP21Lx4Hx95NF/0MMA8oxb6hgQyCadQ+x0ZIehIqzQ+bCs
mNJpMak3GCNH/2gaOPj6lbZ4ZgjVZ/YSsEf3GqHOSok+WFOlSyv+72cvoRrfD1LL
CE8Kzry5tycJJVPKCW7xHrbV7/kIxTb/tdi31dVF3QwrhRkAJ2pIBVOWJWDiPQ7u
UAeu4SoxU5KQeAdtxKPlbz9bwAUnMy1GGcgEd3om8Mfle8e43eW1b+9ZwYn6w/FT
v3ONnYnFGX1pnDbKopcrnv9T4/4QyW3wXEF29B2Pq6Pk6E9tm0OW1PlXBLl2DyqS
9MJ+yI+y0OAdwMltKKtkFR5WHN9auFgc/uLGMJtZuIDbCO+x5CGO3TmNy4VyP7KO
R3xF7HHTicWp+hqv2dc+ZLa1TTahc+s0sErA+AK401awLnzK6DHgeMHZ4AXBCXAk
OIFI3VxCMKnjbxRYWd9Eq0Q1bwsho8XA59ejVlUf8NGOE/kLEak08i58sX6B6GBw
PwE5ZZCLP+t3zHX1p3vpSMG2+kfLKCHqtJaagYecVzXdNwK0cTxMFHZFtTneBxKR
+aO0BZpGIu2+Ypuf28USedaiszVwPIrCMaYTOfLjbOb3EmPLomiVN/RoPin2NY9v
M7n5+ruysMpvit2/W1jORKm8KQrQPwR/lF389ERYws5ANBim/qASAcokBcvKPPUW
+epCbUzcJtDUAtcER6AZzRWgTb5iIRIktlVm0PXYqztTp5fY6+owmlRH128PxFeF
teH28DuSh6e3k6tkqjgvlI2gfX9jQXEooAh934+TUDIOUpp8yFefNBj59RAZaFGW
ECxdATQV7GBFXcEkTzs3C8DhyQiUt7MVobzrbObLNW6Y9ZbwsfZb/OkJlcQ7Kqa4
xEMipsrMO1aC7YPw8+CLg5LCnLm/tiCiX4XpKmotRcPNjcjvHcbXAkIzCnmAmu0a
GHNg9SK9OoCd4h5Zhtqwa4ZfPTV8SEXyGQwrJfQAfAGZWVFejxMfwG7J8LohagA+
5w0vU6pluoR8EigLi7OSc8yQ+0+sKyz82vPWMc71ifMt2AsCTbp6g+ci6pBNGQsQ
3R5IOTyU8att132bIOuIcC6zYmPTfZ5+WNqmvbpgNkiZOn681qC+KmDQmjvFTd/a
wTAkRtxGnvcCd8bTfzKMluBUD3P20FjXPvJNtAn5EUUtrYkJ4ycpBQXNENM+D31H
/xVQOaq4NoJI1aYUXf57ns/IwVps/OcZm5Abukr2H07oZXHWjkQp6iVZs48dQxVt
BCiMSV4KaahXS3iY6sD9rmTkdoFHqCHiwPU0YD5p14hYuZQwv3j+c7kbadyW0+s1
e1qPuEWO0sYrOxsdqX424YxegEjR0YnpV2oAdKDnpgcDZuwA3W+oPsreKnMKMPH/
yWhKOEWPvnoCe7/afTkd1vPnmx87B22RkNF7XZk3P67CTFb/pcW3Jt3FsV/4Jvrt
MRv2dunMEmoqI0lJJk+pz/oSt5KHBagsF16w0S5jB4nKVrccTtz+N3BSI8r6QxDj
tul8T0HQMkYRaOrQacFVWPmZJf39fgsn36KmlZV7dUkmvjpcIfat2g2nCOo7gjlL
BA/zX+QAWP8UB8aPGY8qwlT8Bhkiae1CnjXvMw5sSGPwyZTHedCa2R8ppXB0YuEq
W3IaLZgHk04IstLar+dA18nh+CxCp+aFl9TMPuZLvg8W2TX1xGPLdIcJlB1YfqGo
AC1e3CV5Df0F9AUgTBrWtA+bWRcpg2JM+ln8tgndLH5I5c52DDWTJcr8akeh9wMG
vRO4gnIQgWnkAdHiACEEs500JyXGiHpsUNR3VpwcIhlkof8Fk+YLG1RAzBFh7nbM
yVcjwzJWTVjbA0qPlEFSbpE/JYgJylXfot765OworS8ry9JyywUMstWrlDz75eYP
`protect END_PROTECTED
