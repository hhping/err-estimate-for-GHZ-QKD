`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/LDX4mlweoUb5br9vshCEnN7XpWFKROiYtAlLuscx3wKP2PMFbrjFxfYGh58Svv
eJIiMWq8GnEolE7ojf2qTOw4NrUB8PrL3Ts4m/p75GJqCHfyKFJSaRGGlX29aFty
pO2fQUqFkehDi/UJ5bjJgeMhcE5hvxUxBLWfCAndt1eDLCrmfPOB1gxgBJHgV6nu
r9yr2unH5U6Hc2ZLK++BJhpO/dOVjYLK9WYGXRGCczh6BvvQNMQ1VJOt6E1TU7B8
jtyl1E2TH9H/3wMFQyhvf2tNC7+h++sy4v4Ef+QQ3ax6eT8hM70mX7LP20KR9ggd
oAay0HsTZRlFU/Qsu9ZqgcLLD+wOYpwOmxSgHUdThsCjmNxQSETGll5t0O9fgRAn
sRmrID4uYO543bKogPtilpHxrHJma5fn6i6Kyb1Sb5QbF4zp6byDkIP5dnmG9AI2
/8ZjPZDumIHt7NH/hRfhS2Hxv5aezMDRpWJ4lx9Qo1zRQFQloTngwGrE3JS78Ha4
J7ALJZn4x+tAsXl/U7jn2fyqvmdvTWDV3FVSqHiG12qin3632hVmZrkbXN9LWAas
qqcCzTsbJfFr++lO2K+S7/5t6uDDFelO3spUKPg3tKfARbZNcUYJvzdy8WgmTXsR
mgV6vr3VvuENGbaFqKXGN6MsyIAMevVd/obttEf97/GfHX73FeoZorRHLKchysFh
vG8flJ/PDGdFrMYS0pVjXHWbXt6K2Rz9K+z1hOSm4KEQTHvzHlLDWZHhYi1cChaF
BKSkTEd/RjaPrYwU1cfHcIo0Th2v9hWoUOchMBSwkXUCBmz5PRpZjgf0af2euv1a
dvJn/arkV4ars8JckvHrZoVAqEgqbWB9rtHQngIv7wI=
`protect END_PROTECTED
