`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lz87DzuxccnLsMHgSNByOKdl91vXeBhY8Rt87Jp4yItj5Gtg36zcmr7YoDPh+2BR
rJuisPA/cic+xU9uctqup+C9GSgwQJwdiS1UhcFn7NcBZ54jVpd5ekSkM1ZvQT/H
5q32dbH6C5sJ7q9W5vKRUiNFJftBw+t2uJBXXon3Pd3dBklj4ntuUqs74IckJROE
`protect END_PROTECTED
