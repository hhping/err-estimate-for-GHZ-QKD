`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RZ2RDuCo0rdoUWilxC9+E/Q/5LnyzUjRzbCrx5Qf8W8yTyeCUPrE11OV5A30SBY
er78maZScppEVOu+mBRi7UICxaoItRtMDVTSYDPOePxuz7WTTn2EQrstkuphK3mK
orwEby5qP1fByC8pTU6C16behrFtZ4UXXulp5KCTZp9ZIcbyw2NWi7ewiWfDoB10
9TIJPfPndOWKx7NHotwNHJlLDdY1xhdfk9reSnSOEcSb4L2vm2615SekzBg70w7U
uFz774X9C0J/f62acIgJ/pET8HpZ+Zj3xSwhp3GzLYo4CY/ak7K0Ydgq9lMMpZxd
IVhX4Q7WEYE5ZijelOOSb3oNlPpVc+5/tsFndsyi/DpsPZGlLTRQPNHCzlk9Ir6/
4iTMGvV0S+ZWkxcrgix4wyW3EkXUHkYaNyRstVnhTw7DU5RoSxVM9oWfc5ykpfE0
F5o1WtS9HfYmkCsSvWSPd2oi8exJDBu8B0BGDTzYRRXfjSlIU4mw3FVUf+js+i7z
4aLIp+Ye9/Go4tAQTSEkaW/O+C/IDCCtboA7okD9pRfkdqxA38+qsZ7ChwIoSnlV
WvgHYS2+IwD2AqAb3Symd6zeRiYbf9kscEBNEABTaincIfFYi59nhGJF7CI2HlSW
2OfrMfQV+2KCofxEkaOjYabmGra5g2i78bF2XnN23CnJrOoLpgF8JZb1QHMXiguw
581dYANLc827QOy6GJ8p3yf3pMlwROhY07EYaaCyyQ2EBZr7MShDFQZVEBaYlO96
D5tMwuv1lky1XJmq2B9HnWNTqWX3KotZo0twYqYOH8YwVMLHUrIaVWkQd/L0hKB9
EEMvqIjIhIDotGmivKRvUIqxBjDRQyKAZ3KRqOrN6DiavsLb0bEbGGyCcG2RKfSq
OBTYrFC1RatvHHXUC4ZiAgvOof1HG2BkOsRJxMjAA2efjWTw2ZRP5Oi1I+G+uXmv
Z5T+1o/SYzNMdTdcRT8Xpq5zHiivg4vA0umFKsWkeXdBQCDbNcdhgv1oBYpZJv+0
OECl3At2i7OPRVsTOStGlJF4NtzLob/WaF5xXwoeGuXCz8v0ESBXynOlgtz3kn3S
KMo247dX56QVs5aS2QBOuLjpDa1akTcxmCttOOcufyzJVas4DS3ueIDBgE4K1vC5
`protect END_PROTECTED
