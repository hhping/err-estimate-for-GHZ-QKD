`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pZvzPUvvkPdpdHc4r5xEYw3tgNh2l5K2xdGGSkZSUX7sMDEbwX8eo/RKLXdd6iLy
b8Kndvd2CLQ2JVkuiLYXst/Bnp7n24Hw4fZHDPZU1wNQX0Gbhp6m3948fKrqnPRx
lDXgy2fgH/kqJOuRYJoJ18yxX0sEV58EY3RPa/SXS3KhygbWN5Lmh37Xy/XmXZuV
xATKJ1xNqu5imhBO76q42MZLUEDmBBkTDzL7Ebujx0tuL3WqBeChswmG1LquLJC5
2EJuulsPV1KJowtuhcIh9hLl62CiaPN/pH7hzt+UnJXL9uJz4sW9Ty+ZIwYIuE5L
nGPMcsqv3wjPIVzWKMP3vtBDVTCXKn1o4frdKS4no+VFzoPbuX3NLHUcGW/CrIhb
DE7WCca+cxj4DbpAfP8zoePEaTQAdPJhbsBdMceboSIxJP4RkxlD9EleMUSvQfKJ
liosgVuFnooqzBqh5xtHLrLnJZMfMs0ryY9/lzPorWHlPYOlBANNpPKgAir5bpax
xkX1xptjmiHguoMzlTijTyU76qLIixhhuGt45rCYyxE96qWH36G5q1jKR+VT34ld
r1DkBapuO/iFbtbCjaxI1AN1dX/uHFMDGJ+ms2W4cMJZZKztI5aJhV2J3iT6A2SF
6/hjA2xauYarGMwibESOZEicqdpBiijHKF0nIaG5DSmXoTxBb1wAQ54ujbaoPUS9
a3GyIOYxJ9jyQL28z5sWqeB+NN4TArhhRhjfaaJ3SZCiPUbi3mqVhPi1y275R8HK
J0IbC+/OiMjf5zn66/ViFbUlcVEAaG5/gvaA1uokMe8=
`protect END_PROTECTED
