`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFDfJHjkrs68BE3zw+WTP+jKtaWHhccN87aoiMOjNpTzPtLJyCvtthMzKiUTvbfG
oOVy9bbeDlm7Y1Gcpqb2mRi8i58Tv7F607hZeCa4mex6nFhk0lN6S8QDuDeRG3+0
zMJnCh86HEoAGNQ2cIruQIvqElA8PZCP4nJKTpihcjZSEgXIOUKXMDIbxppTfqhC
Vd381SQ6LLFBaRyClv6gsyurBt7rTEcfLvaCY4OkL1oeI7kSQisTs2RxMIG88Lby
kwaY1Rc5SqF5TxPZ2ZV4WtK/WfnLPKQwYBPTLEOqbzW4YC+M3jsrfT+AwcnJqVkE
FAToIP+/NekHr2pGZTqPfPG9aAW6Ap1HxHE4s1AH0E94OpaJZztjbu0EP8ylw+9M
km9K60Pm7LBVZZD+Qfsz1RDeytuC1wHCO7UFbuVU5WnwthrxdexMO548OfAgTLxY
f+Wu+1ta8UV855If8n2Ikpam6UAHAgVnV0piXiHFvDWYrb07+IkLPATX91XLOcwL
mEcovNK1U5WG1Z9tXA+cZv/QpoE0/iV44/kXsKSNBm1cTIgTNjQwkQdeRECIX5H6
sZKiwWGflwyHVzgcSFhqB32q8qdwcNqO0NMI92mEzs5oRdut1tOrW9a56OFCgwjn
/YbrPPKakDit0mqDlfO7fn8o2uOn3XfH9FCq7b4KH3m+F8jc+QXPsfMaYpiHR8om
h/R5Rzo7O+QHOB/b/UgRHj2AO6791NuXQZECSqGK/eU=
`protect END_PROTECTED
