`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lys9Zs8fTC1/G6ObjYFMhVI3RE0SuhlMBDIZgKOtHPXVJId+xxRuFx98o2gPjezY
FZ/En8l7rOCXP6ffATMU3evwJGaIPxRpy4o+iSkV0PY5pOvv71zRnfuhWCErTaVs
meOA0T3eJiew2B1ExSyXqQCCc3sZB3Vngcj9J2XxjTkil/MF5cjUhK4LFZeYQCDT
kfmXwPnBDV/+2ncpZ/ILVU4/2HtMAmbAwqQ45T97iwP7PEHrTd9fEDBGNkcMDIzF
U3ReDVTwj357spKkcqucMjSbjDe/jsyH/ZBcx5di9K8Tn35H6nTHc5Pvv7BAmdqq
B94NJPyQov8e5Ei5iCX0m1yV3OPdS/2neqjxUfNFTHMrpnkpsKxBYCKAG0Z6/Oq9
4tMhLtmHCUC8wKTOU9Jkuqb79YQ/Eq12XH4eW4dtPAMZ9UPECv7xa4N8utQYoxL0
dHVb3RyChKpeEuvY+vL4JCjHYZc1F7kDej5itM7tasZHPlWw1SVR2FhGY2kP8pYj
xjmSiSTsUEWQrYpjg86yM01HWAJsV5q5dyicH8p62HYdU4V5djLbyDMoecdDmkHB
Yx5k+h329XkYihAriMrktGpP/Lt1qCEtffZ9opFUkQ06YxgjMberdg9LIkHqycvK
i9VxBqj+6sWzQJDHD1jmQeXwHUNmGVhOspPrs0gKcFZq/bcasfMuxNND4kzPnLIK
xFrQeMUD4TPzJDwg+TJwpnTj5jA8Ex6z3YhzeNtBHsbpl96VUiUb9/DZMlVomhA4
jy7/kDbKKEmVSP9VInNup8R1HaP/eMaiiLK8jq2fYjYo+Aud1JqODmsLGZyuyJhx
YPMhrL9BZ2TeIviAx05q57GglOFvsfmXlwmpBRCRL1ero/DWoOz23EqnPfTON8bL
JZ3+stYorMogAQMM+eiYxYsGpYJ97TSoBJZHHmeCDyyNdGfdx5ooU41NtT8nl9ws
z7Nsyhu9pAFf5C9xSapzy0zpj0nh7Sg/p/HarYaTVKQDofA7OBmc8j0j58an0Itq
1DIeHfT8MTHH2w2J5HqjHHCRK48BwCsLbYCaipyd123Beo6q7inv254Q0HaezDj2
Kf5uuTZsp2BmnUfoOwivq7iEEHXRI0LsNEAR5Lb162i7rdZToiMuC40a4iNYOqV4
8IyctAdDRXHdeNmE/GEGxBc7rj2ZcqnJ0nT28Esak8e27hPuDy9Vji8C2R/fVei5
qb+bKPD2W5wUpc/ZFq3FrXCtfmmmJ0mf0q3+yD7LbGJrpdSl+UhQYCjCBg2dTE/t
DrG/iskefi+x9euYC9L3PnsH6fYXDnV/sn7Kk1REhqRxViD3OffOnIvDCYu0AiC2
zJJKPTOGb/to3GVs14VRmEqn7iLsGyOGfUI6rhcMJ0B+88/VTlmy/GXlrqDJ9WNq
2q//QkHMaTBGw2KGG3MUkBgGMsQe9oOsJCwShYNKUPyrRFMCtMyuD/zmy4ASjlNl
KcjJhXxgcqPskrvgQWYAxjXA3q6NdFy5UfknUDU9GXAkXmEBpHfO2GPjhn6i+jaz
dohbln+6Y+N+y5dOlbryeWtPMUiQy+WZPbxirbM96UCb6KDnS3YgWRZos4+gjQkp
RRr6Jf/xXy/AMRcRExiyPayphRb9Ldnrrqbi+YhF0Bzx4N888urj1dlSL3GNWrK4
JjDGEDhv+iIRStS+i7HUFOFSSFeKlpVeaFMwdXA6i6aKZ0dxJqoVNkQy2zyQfQUI
ELL7Mt1AtKeF4Z8CgsvbYDhT64ocqEms1vwNKyq55ilQ4CELV/lTEdbLqvUrr/bD
h/U36dRLE65vP/+Z7JTxMR6p5c4iXSmELVnau7SYpGiVOs1kQaa1fHkTmd79Mujs
oV7hy18E6EhHSZLYiv0Ey5pf37vFTPwdZBk2w1VgH7eGAruiWvQhdkzJinjnCF4m
6RDTq4F3t6pljhGLJmdxBOMuO1/DCoZQ6KSpritWzNmisqyxweodInPNqqCCsmFy
SxIwOeoMVBb13Trfic92o5zZZT+bJ5gSPvEduP5NBQCvrH7Kix6V67Hdg7zUPTWN
RSLG5xf0EEXzn7ubMnWojE2USBIYm/9mXLJYq4Z0fmAX3Gx/MguSA6EMcFXQ9mEz
OkDb61wTnj+NJh9wpf50l25mQUH/MZAB40mh+7TPJCTofU09wL9ACTq2PycqWKtb
gmvtj5bnMl8K+i702DfyZO/IcZDGwxva+eTKPYLzofPv35tMuL9uEZ86H15maG6h
2594/qdSXeJRpk3o4NVlhy1EAfxLOOUei3gufmHlOOLiARu5Pscg1mTIyJmasPX+
okAOq4m7a+X6P7YHVYwXVcbGYoBRxMI2okybSqppWoIus7EFzkO8XsLwUrw/TvYN
dTjiwGWHAE58HlNVDIYTfI19m8s+reldeOAFwcGFOCXWL55rUhRFGsG8vcohH4tI
LaKzakK1fxdH4gLzEHeFOF8RnC2lhZ6RY3+XaVcL1sDat8UdDda0UBgDLhFJDC9M
LtCcaHV4S71hqvEqxdMEHbmc4WOe3uFXL0Or0/2zpexPq7vGk7CPZsm2junqS6U1
BS2nnWV2haUPY4LkCmmab9pPDzYJ5C8m8YgXTCrvYjQnImB0K+k/4n6Rr7j48uFx
98+LFEgQwZDgD15BUTkrmWxJjll74dlc9qMVTzbGX+dhPgQkXa1YdarlkLg8yMop
A6XCWToZr67XBQc4aFjZ6qWmfVsI0BzSdh+bh7Y/PGZ+gcqGoOwYne9f7ER3mvfR
JObiQ8R1KQfiuaF+l/JhyvijA2HNH/4UjSFpTt4INw62Zc41gxDvk0Gj+A/1IHbf
XAbVEYBJ8dozep84whHNl55zwdcA7CgwlizSyJ29VeXqXmtVvRgf7mKhbZwo1IPI
TTFrUMLK33cJ6xCMawaHzPNb2FKetSgfR57FhY/h/aquF6ILpFUSnQk1UwrpOpRa
jKlJKFDvBmawghugg9GdYhlejD14MP+P0v9EC5W1RgRNc0cdXwQMEn009Ka5Mj3Y
pIu5OZuske8gYzMBbRvQqBoly6xoUPFVjYQNmgMGyLcY5MVzI9mOwcy+kcNzWEpf
c4o/xi88nF9Ff3DTcQaWzzV9QkZSC1Cu5vJkdP0zDoJrS/XsXxGMzTAsMAxHHKsH
G4dBhLkXk6OZiR0CbtY2d0BGYDT5oJJFTuLp8RgCZsaj80fXTBZ1v8MyL84mxR0b
G2OI0KLv48cOOdrlEqxHvlEic8q6u3q9f++JIYunTWjT307kmdv1fosuR2DdeYoi
SqEMdtdQjUqb4KKNZe4kdQu7SkgaG6AiobQj/DYUgV/Bn09wn6z4xGfK5O5hJh1X
gWS/zL2RBbm6neSgGH9VR9IBWJwUFx69jOfnp+24Hfp+dQpwXmZSAyQj6fBawEyx
fCLnlIBSGNA9Tb+AdsXQmzLPmLL2yFf3J8wtNaF7BE22rCR6fVvq0m/d/XkY8MlH
9NORYt4I3ML02KDdr1+JDQCrCOltaEKCJIKOj6VAeHWTxs279stGEU7XW6w/NsJc
2/go/kUk6nWjJCTquggYtgaoSXOak0+9YDQuIu7ZBmcASgK90IyVFSYAToBGn1tL
gYUtjkwJzNNuXSFG4dhi9JSNAmtb9cEGJLL7pyKIw6M0Nj0JY0mz25RTe5IlTqdl
XFObsQxejRBSDipoMR9F48Zz788ngsFaqXYbNlAqrkq4VAqbvhv15kevYUjL7Ath
kM81399tkd/Q5zyn3l/nXL3evz6GgWykJQjf+WrHi8hNQm2oXQQF+JW61Wvwo7m+
sxJscRkvoMN2hFcYeZ7iZ2m3cwEoB+viVPMF1enq2Hkqz9yYRH4e7VK6Y+JjvaNY
BbDx17q0iZow4ynK8JxgMV5RZ8YGEXSXLWIF7FLe/x9KQeFzuOX2evpkevwZ9aNY
f02scRlE1JRt84WJXOjNsedGS68g2MKBYc0uMCjeIn3g/JvY1r2AtevvE/88BfQh
ksE3l5rHTU5QOuULdxzLAq3k0FP7RWe8YYTH6L9f9oAG1a9VtV9mo1GrNgpKxfaA
m77Z2q2F6z9Wi+1AZzG15CY+ywv8sbkE5rHBvD+dcPbJM9mmOJlzX1VFND0/Rc65
Cui8XD4jDx5crO4y8+vHIwimYSeJ9aysYBzKK5yvQwtpJ16Dbl46/1GJ7rTS8qd9
RNfxZGCiDI6KNbuYadB2jpHRBE9SGr3eOB0W5/rUSmakvtuycgV4mHC0ilqv8qTw
WjcJLI/8PI+ljVAgY4MQMgEso51nDysvcpOMNM+lV3zVjiqwRwfnEYBGD7alJXBP
2i5B0Zzgj5OqMcyLSKP2uOWXF7zBDnxdqhugAl/Nm0MeRrjggk8uYCsiJyykpLXa
CNInhuBTf8gUmkD4CDKY7Jh3s8AR6QiprSWRxQlVGshU7eiU4mf/ZXhr0oJl0+YZ
mbf6Qegk4IIzRSTQ5Ujxj+ivJdrbBjlYgTPFtz/sQuyq0B6WPjMWy1P3gZhdceGE
uWgOdtqhiqzdWWxr/XLmYyDtl2VIIKfEqRZ8a45Q6ue7IgI2vjRODvDgHXkfcM0r
AZvTk37DBXugD0p9Y79FdV06T/h8+stcPGO+PAn644PKLQlzl2ndttU7YmUyV4mB
ntRILkJMiZGRMfmPA9uNoEQO6l07zemSzqir0Ls2Nk0teY/CAqikvjY6lKyTR1iK
k/3BtJZcroLNVh/JEACakJ02niKOWoxszZkVDsdyofDhfwlBXPMMWH5u9Y1Yb3C1
Ns3B/RNksnW3kVq8Yzp91HC1rF/lnEGLHYzbd6GJx7W6pPghIBcJp3+DRng6vz7W
eIwV9/H2lzQdYDkjtGheQL0kBAZEebaGB/TY2exaG4cX0nkKP8moTNW0rBKjm9n7
2TKR62fMJp1AVnEHxNhjlroQzYSPKAetOVCP+ODV4ShRPBaR5s0KdfNcVXfpeL3K
pKm0abGDFF1wOm6CbP6ScqxB4apOy2CyrwnQ6pMMgYl7UJj9fvOHF+tZanhE5Kf4
qT2j0ZUJA+bdebJM4IbJohyA60yJSQfmW+oLK+HohnEVZoiLJBe29DCgCUHS1grZ
egq25+3JMMCWxqi7i05ZN8VcNvKwTqlX/ifswhdbFyFd0pYxVrQPFk3XcXYTpmCm
ClRdlt4wNxYwuz/R7kuKGgo5xvYfX4u7sBzFzWofdVfPCG/0jGOgwJAxrkGWdzlG
kZfkzyXuaaQn2Zj7QtZoZ5UFZWXR9AgWjbFxmCpNDQiBMqXk8oVglyCshm6J9fE6
G159Uugrx4p36y8jLsmw5KFIdagJSNobrEy68gjE6/poRH8VLG4LQJiTLIMbiaFW
Rd6iImBAiDoPkG3vTv0UsKnMF/bCA1CPEDyPL9DQ0VTR5bLJlDTjRtH8ifN1FLgO
Wed27px0U6f+Djg8hCM2MGPSKoGo1ZbtcjtdMZnP3CYq5Wqoy0CvkfH/3m6YRSF+
+Yl4lkp+RSD4Q3++cbhuk8vcT6SjR2z51VBG+ff/9/Fwy6XzoWQ9pwYZDazR/Bds
zfak4fiIPxGB5O+RlGEnJiqeBtQjL0bdweQzao64Y8k11Kdd5kX60y6YVsa2gYZK
X2hEnRt7FXtPnvRnetgWHazhViimzM/ZQ6nCMIZb4/xORFhbKryHlNghZ2ABmvoi
PDs2Z3Acwy5CJaFW+sJSQsNEYajBaFGHCNvmMiErWLFnXklzVAOR6cV4aC7U1+lL
GlCkYxrJkWY/ZAm5aqzTqmOA/wkWuBytwNgo8wbYkhGsvy8QHqUlItDGEYAi4cLN
i5PT3kXju+B4EtMoHox6mdyABdqB7Kv93YTfGJ1XmlodUgC9pUKmPF2yTN37qzFN
sqiykclClFvjO92L3lHG5EVEtHf0tjaq3qBJQaRJFHmeiWkIiYCxm+SjqmccFGkX
Iqz6N45ZUb8q9a7xwxq36nzqjDXvyLjdPlS20mm7D3g6ElibqLvcw38/RyE93622
RVaYLLrqBO+IOflteY3Hbn1VpRbkYEiPgXAVKLnW1nc+TEvy1I76BhjWOhcZX76I
+Wov+W8SUd5tNDTWn/UM0xOYOFd+MdOzOVxD9kPt+f+sMRZgl2UpaC5zxWNcKnRE
jwePx6QbTh3vFvF8fmYsv4dchn+3r7XCxBouPB8CJr5PCZ5VN8LKINbqabsj093z
uigsBakxG2Gk4eFJJTBkMS9o4lIGdXmRjZJOb7I2Bv3ag9+QA1BhMA/ZTjsnTvgE
OU9IXzKoGcaPOL9b/zwHr2KxLjsdjAFH77hE1eC1gHWsfJMx1AhocwhMHb+tslCq
2sCiHmr1rE7Z4D2DNzObR2vytQ6ezSVe9caYas1Y5m+QYeuuR1u3pInatrDtDQ0l
1K9w7GG8lg1NvI1eutBeiusl9+bj7Po8W5Xwdcj5oq/IbZANr2osNAEJJOaQASqw
2l/DBD/0iWfM/Kzh7wkqhuEn3rKZ+nN6LP/vk8FV5Bvxvd5FiEqmnXl7tBzKHczG
WjYBo56CiBiZRCpzIjYr9ICaEry6lhY3h8P2GPaK9IHeHmlpSnSuu50d0Cfi7Yux
vw3XCNmNLOtduH2Spg62FY1q9WNaQUoYv/hPf7TGGkkWI5Mr9xSJAg0jy0By2C5C
mSg08sIXXh9QrVoTahIjKiKZhTtkzxyFGeDMaW/Hm5dQqiZc+kB+Yw93PHsxoQHr
As8PgzT9UhdEh4dC9smq5FMmvXx+JkpmH/6YC3Qtl37Lh0gsvp6wqmXcaPjEe4Jo
E713JzrCDdvWb9eTv1HUBNf5rS/XM8/pgxnKLanVxgm9J4ERC/9lELH3NbwPL3ZT
V3qmopyXPSIumbVAIhZjtavOA6XqLBZqIlI0WCTHc88kUbR2F7+4EM4X2pltQeJI
GOdMNQL/MdNlRYMfvgnn/khMYKrJWzCFigSbuC1XQFNU57V/A5jIUERiv3UnTyrl
kT7nFt0vnti1/hWH9r48/zh+iCzNug8F6SI3j2/kjLoXgm4j8rAIlssBEprd87Qx
YMzxfmW6GFDv7WZBnz0Z18S3iTq4323PqKipdjJEIPSNCtaOkyJ3Tbp0l5Ct5RIa
DMS20de+50naNnu2SHUNtroQR6U0zaIBZeJ6manfMP2JHbeBWG+Ex8XsDwi/HBy4
Kue5yHVQCaXg2sqI/djDH1MjxDAeQCmnrKHIUXAFJbIjeZ/jSgx8f4yEagDI+doQ
XN8Ai4BiY4aIUIofGdH+QYr8AvFarJBsUlWI/T68Oas62lYzu4K/eFln1LcDxsVv
safSoYnRIIkSWDBmhWaHYIWMGnDRpjdnm3SOfxQDX0hKj5615JLzf/Onlr0pYNU+
me2sYWK5g0OJOCrVPXuzKpjmu/1aqX/+flzIFAJNy7bXyfg2lXW1W13BjSOqnNlo
yvBxV8NjArWbl/xFf8Z1RE9D6av7LQeZlF9Wwko17nyH4lF2XHRw4y3jaPfEs8m8
vTMyTIbOCpBUszRpfcSzuoSQNmTath4cih6dcb8lzm+EeRKM2/6on4rpaUb47UMi
b0HgkZVG9gRDlCjCKSIaskpXsHET6Y4g9fOUGwwlUgguB2XvfB/P2LQcI3+U5Fge
bVSTcQsCFP6XfRq6Ad48B0HKoEhVNGM1OX96Xl3P6NEb4iq/4RnYefAsmH1fTn4J
fwuJRbKcigQAnxKfKeyaVMDGI3rW4X/i2nE258tpVpEb3FLpcK2nqvejxRAJyFsa
vcwGs5VwRZjZOdYj1C+3w3X5mEs1OztM+KrJAgxguw9RaqEUIEmw55grlv3d264H
LQHP9G6pDJcd6GqTEBfIOQFdFQwHgzTn+BHurXwCR5c4V4d9rpMOQZNp2NbQkL6h
Ps4jJ1k+0TV9e5YWXb0v5AkkHFWgDXNaEDULSvIHxK5Q+lqUESxLlvks5UEHbKgN
ZEQamf77WdIkiXxImmw1X5Ymxop+0LwxfMvU969wfR1kDRD79ozv1Q+6r1Yd+5Fi
9yzgKtumxuNyr/J9GvxJkMLQUyHDye0xK1DBRP6MdaQbB8xU2RFhShfT2WaKj9oA
B5wxpeQoToNqUdvBhQ/DQESjPuTYIEBTNOVZF/8sBhfdA0OKiPQS9uwr+OTfultN
FRi1u0GlhyLOm5kg0iuiPOgvKOrgLqHUCwCN50XYtRdLXP/VvsxzIleppSRrHT3P
KSo07HM0Aauz2F3tPes+c8dFGlhQzK2GicJWd7MLGU68Nd1xgKDGeB1nyN35/m2L
vSH+2vfYd+j4QDy7cydbp1lPSeNzkJpdga/9W4UVjbQRHTyIV1gELnOT0u9BXAuI
1h1u437CzE9rF/6RishxJN6cdDp1iJ8wHoG/nmcmkZwgYXH+CeQxfKVTr99xpX+U
UpZBqpmM7mt1pHwH/i3AB17HnwkuTQeZlvjWu/g2j/EXe1WM1IkOw0k2AtrN8Vkl
wvUZBbuFmMI44d5XOip13ZqGxm2dNCUKQdr8M4JakFVrhCoon2QCdsxGK7zg40AB
lf/aAEjGNwpksog+QMOgsb5Evu1W8RV4aeIMtcfbL0KbCbNmtat71Lnjm8DhWiJZ
2tCbneVZftXmHJrGNEiYHSNa9zzG8VvWrbNLfKmVYcEhoCA5UyXtSBIP95Xq5zWE
ohQZmM0zQKmcEi6nvxe2Ld2olWHngQ719AZNxQCHH96xm3J1N6UFpdVJoDyTuqBt
79qehuOGdChHJ/UiNXTgrCuuJDsB9AIc1Z1FkERidAApDGM9JKr90ZH/CY9pGJy4
jp+raStY3NCM6c6XdHY1aRO8PbDr48xgXFlg3Qp8xfJYUiAFwLqa2Qpdfrs8AfYq
97TzSBosq9+JsiKh/9CvI/GoD7fP9VfgNmZsxp1P5lR52jThx+wLS6pw3UlFsP1R
3+e1MQBRKl/QZy2uds2kXisnZYrg6DPYaA3iGsgK5zsfJWYO8ed+cX5SPxIlj9/q
yLsAeXIt/58iRX0KGDEy3dfPy7GBW0VGabOWf/Yg5Atvvf4q3CyRayiaDcqoCkn0
H2w4yQ7X4cN1IHTwoT+jABuoUyN+QlzbweNEtt5hWWt+O+lqKBpwopQneXDHrD+Y
hR+kGsoq6a65fIWRFmDLy8Zff9iRsOxsq04AI5cttfiiOPI1u1Bs9kkd6KISp4R7
e+/iSQpMaF6H9oNavK1AunMKFmsLq9hK9fIvzNbfk1oi1Y6levJcwSPGQWr+qgSp
5jjPT7zyp8UO8wX3m5YPKwQD7ESPl3z4teM2Dwu409d3wA+Z15N7zumnimHwARSP
LKnfj62/dhN3rwfD2+hbolx8m066QBOStXwOYuFN0ER8Ig5TjmnB950t4WafLRQL
zH6GpPcVT4cuidyB4IBUrcfGUMrBVGobA3ZdnrYBsZc7RJmzqCWYT4q2wkcHlNCn
2xVM8VYBEe/not2LHsACB3R9voT3ighCPJsa/KtvbZqPifWuK1MtKe+d/NbFZD8S
4tdJ0ocX/obe0pMb/eYOmYf5ajTZSyXT/+QH3PC8woEnyCpaKi3EHH4gyVZ7I9WT
Q2D61xApJXb3/ea7DQIwNWsYkHkZPEv8xxtVmPkRBJlbZt+gj2s5fjoyGRk7vFC6
hGOS5TPdrDxeAM3F2wLtQBIX9+XaRjZTiXi2izAHth3DZv3ZoSCsSEID0e+aggZj
yahxLzhZdtRabKgOdJThzr19p7msWI2OaKEN9j+Va73ZRMzHbBrJSiWbKQe5x1K2
DJOFeQmZsSLy8XNXjtHh/aaeB+OgktPOvKwaAA+yro8zmfFvQikPM6KHZ8Fj087D
OX/FbuMrKT4cQQh9WamHjsUy9nRbCnq2IPx+TAad+92tCDu/q1ZuN14uD2wJ6NMc
f3LBFxTfTUQwLTo0+FPaOzYC1LiCP2MjLp7x/XlCuQPS0aIuch2czLh/8Jm2d5dc
1xBhNi2r0KsXV7aafbDd/gfsPAtP2xSzUwkt7KaFnISHtOUGH6XDllS/9h9xwOv4
OEmV5ckkME8f+UmQl/KYlsazRbDW53+DMqTjlhh6JfNe3mvhOjRKPZ30MXTQ/VJT
PdjvxcUltZN+I52YNgwW2f3vsSJASQTE8wMFqUgzVIJC5syBljUawkzlDPmGCR9A
AYRR2F01Y+fo1c+lXSnOO/kzaKo6yxqOO31GWSrmWKmAdbKdXLYVxFmncXjsaVwk
st3IQZPcS/vG2H3SB9SuJdqIqJ4NnBvxFkbUZ0SFbeDEfnzRxJcM2dBy4JTavCRg
ZuCmX2qhloILtkcWNmgwySYA5xUtBiZcm/nN83U+/ydWnNz5lBEMl/LGB1rn/VKv
sKRhkOZeHWlQuf6apCXCPKALXDZ2yc0GGMjCZooPVZWtPsDObpr1wyYllSOXMKNb
3fO79lrlUKU20d1SYUqZDR+kR51pCCCHM58lvmwMGM2vQ6LS36D3GLIUJFau4rqS
h2d9Z7VYrPGHCFpAr1kYRN8Sp9FUk9wmb4uefJA7wXhe/q9aV008+M8Vpc24jrJV
18zjBLg8YDZf4Rz4ZwkgePkjjxsUi8KR2jo0A+YGUHIniO3zsr/e3rTRwUo7IYo8
BlX1fl69voQtvpb3shyZVXPagUZJG8jQGpRTVkZCURHidU6sefoaYjZc+qCe8SqY
CbdxgmUDMBEEdcJHa6HO8A4UhpAdfJZ7aJPijO/5u0CM4G8q/zuyAgxIu+SdlpCd
nlx/mQ1q3yU71nKe2HCcPCxp2L+8udvfDBt22d+yPB5dcMSRfAVZm35jxJ7T010T
haj8S7barAiNjTeJ4XBuSnNbvWIjt49Qg9dukX+3Z7+6O76KN4Yn2W/SdWBhf5yS
CrP75Rt/4NNyd2yD7VXOjwa2aBDZHk7usLrRL1NgfrQ0GPb1Hn/dyRi9L2YXotMp
akW07MZkLEaT7ofxo6gM8SqpA8eeeKaaE4xXjOQmCZpBEqXlp+F68J1gG1rfNJIS
SKL0sa7WXKopltd32OQHWNBK/9Wu81f0aQm2C7ZsXuzL+nZr8sxfO1O1Yub4aNOd
GfEno9YpO7wuETadqF/zTtAPJfnrcifAXk+RDchnnNAwfiVtAEbtJfiTjxyYAkDz
OTipgZvAgXS6Tr8PzWQ86qlYPRH0AGB9c1imtTKt8iGzyzHIs9jD9iRRnQSbvdM7
xJ5jLCaTgu3Pp/kkowuiFG9tYLMLdd7rHrPg5IBtui5be0oaZgSENW6n8SIVHx3K
W+Ol/K16Cq9tLsIwrz79qslch2kVRQdZTg/ARkoOiwKlCCEn4oTdiXEiFOLacwTD
riWMzETQAG2hidHRVNxiTx5EZhu2TGrP/Shr0Meyh2b9pnNK2ICsVqsZ76pbiOgV
LicH0cfS8L7dTJCgPBkHUuHO6HKSaY4TZTgsXFV4EGlU5mf8AdnjEKVtr/z3Pwdg
ftzEi5Po4RUJ6w7/qQfe9K/fKYtMABFAHfW6AcZ8lXT7qJJSTEfGZd+zCVBUxWfa
Dg3EzcIGTjDGbPmXeJNu4SKuSmCfxv6l6bPEFzND3iRxn2H7Bgekp0NjwtwQ4crd
kwVCgrkOHQ8yoTxARM5mE+Gqc1fLDhpYtVSxnaMMQIfO787/3BOebGcIjl22ZDNE
D0neR6/+mhFraAMqE8RIbNTah7NRs7OkyQSb7b1fIvV18yPtDFW6D6uoFlOBStSz
HXjuBuQYDKZSbgM5St+d2uq2XZJbCCQhRhi2lr9/tSaHzTXMbBoU1cfkD9QymzIU
dj95iKpKoolVLGey5yVyfM48HoHp1YuP9szFTZHR9JcQ/1NmL8zneJUWFsvO4FW1
CfNBDRnaIXmUUmzB5zegDDYg8JU3Q2O6fp/Tet1XusHMWhVKIsJjp5GSgOpa4dT8
qLHWMYTqRhFRObYS7ncLDnFkxEaXiA77UFTYPJj9g73qpNX+Gr/2Ba/EG1MpRLHX
dnoAjQFEu/P6XXUENb1GvA+TYuTmSjHTlftl0ejJ3TA6q8Hrz8iEMDD/V6o43Brq
a2qjVD0GhZ420qyZWTfrAmnUVc+2caFehfj/f2PqRPy45RCNwh8usGswHQ/0ntAw
qas/7z1wdkgMvN+9mP3qacHaiNVvMwe4+eL5WpU3UPScvLu4BV7ID9pFPfPvSvE4
M+TYNJMjHWSk0VPgh3U11rTBMlcavLC1DaZjlzpnbLY9oi/2c/VbBu29MCph+it4
5cXfIgH2bgHiRmISvCowSPeh3zF9zNh1IgckHKJ8C1IYSbLHuWh4/ONDkA4GxkKv
8lmJbKo7lhM4GswB6vxTpVFnJdaqWehY5/qFKN/4UXYmoCvA64/LqBOS360mqINH
G6JAt5EdudxkscTZ/30QXjccZNtkGxuEsU1ftXCqEz2wuZ4KFEcjyWTE7kI57NOc
oilhYrqVvKmQn63LcZ1qlUFxyjrySIz/T6cdXjAc0Lt89DAJvQXrvZZnGgNAtSAt
qHhdeWQmW8ZH7Cr8MnAVeWAas4n9JML2T1/2bFT3PW7XgRKcczG41zypInwQtEJY
u+j8DHB7x9dDwSKKzYsocUqmK8XAkcT1aGY9l5HXBSri9w5m2w7oOCbtbqYLPOBC
LOKnqiW/1zgVGN4YMM+h5XHld26d2hVK7BEWjhy0/jAGM3hApL/mXtP5CMUZMAxD
i6ZWzce0y/LZrp0DYv35mDhW0GBJgpHfazrvFBh/qnTpC95nw/0QRUH1On8LOo72
8lCDiUsa1VUfX3eXNc9iWB+sr46+8KmkL9BzGLLU5jv4mAGamn53qarcNxBkEHaT
Po4U4knP2eydY2+hSIKLxioBUnCGs8GLzXumAGrILRrW6jCPkZSfM9gt5FY0pVAn
7SWMZUnmDu5mM2de70d0Q1DZQWc4+QeCo930bnxC5wizepz3qXcWMpphaB4M+lU5
mFejT2SbMtG/MgdWjgJ4KJGFmIhVVLG84B/jBudSa1m7MWNu5j1InyiJM5p2wK0E
Df8l4zThgjrDNa+UuC7MwtbD9gTXE/yGkn2vtm7Vyi9kT6QT1GlE9huc8LCORcMc
1vDIpXPQeMA3AN2+ML3fs2F2SPsAY1v0QFGHQQUzFasVWBNx9wBgqKHydc+KZbXx
x3rTTaO5XovW+mOy89cLo8eCdsbEE9ghuWIrSL5or/bWPlkmubA6ENmO0FiHdbbs
JVGLx6zggaq5/Hb8w79AvfGTlNANom0dDiYWby9IbcXaNe+qO7ySGPOc+TjH5JjA
LHut2iB3KcvQeLFFSuqq2IZbLhKTSAYVeIH0Nc1740ucg5VKVKI+0A+5VRJk75JD
HhHcIqCRLYl2iEHkV6+n9DoLnJPXpZP4J+IWLk3RQD8qI2AurlpO0DhomoEzeAI3
SVoaEbwsiZauBAuou04Mg15uY4pQp40fYNXxALBVBsrnsU8goHeemTCVmcJrpZSx
j/sBUAE9P6wGXkgXz1zM9aRX7GD22/tsts2T/cjOzOTPo3RqRX1oE2zsj+hewvyD
TmG4V5SyDR37kJviRiW0MNQrDDa4ZinvPlwkjsUYvl6MoAafr2NQz5CShIl7ZUlH
tl+Pzutn18oKPZDePQb3TuuZGVMAN/JxONVyUNCUR2JHYj+fn2AKZPVfFpbLRbqK
k/vKdCr+rfCNrkyrkm2/wiiMv+8rM1moS74fRKdsJYlgUh3UE3X+mwkgkUE3zkEp
V5sdahp7T2hnD201j4uV1D5L3910GwEdL77CC1XJ9p1cUh8SZfg0N8DNzmRGSOkA
YLmWtHoSrdUmBkPhFY/d9Q7dqA7BzHBpp9d4VIlklRrbUoI4DU1A4IlCsaXhc8Bo
sOJIKPL3jImdBdO9uDEOzaba56mLDSslbTNKl4YRWwxtecXIQ2UjGDMi7Iy6BXxb
x5lNYAjz2AdujoqJh8vqPC4jMhq3DqpIOTm8sFK2OZYNyC7QIll8DHQMV3oD8XMB
E7379yyJbNdl953utVUgZ1wpk5RvRb64u4PDV9dR1QgtZjW/RO2AWbgNyzERXmRz
aBZYhx+cQma4eTEB7uvKnWn6LKUg+Yj2UpO4jwvQJnC6BDFcYoO7ElHzE7LTKlek
MDqrLeXdxvXkEamw9ZjIT9FhJqCot9BE8zW0KNjaDjYY3DHa3RoIPG0EEt//nJ6T
WHTajrOfh4v/uFut2/6f6eAv0fEQ9aj+ym9AMUJgedzm5lHsf+8MZLo+fEwM3rWj
9gjas3o0aunZtSv/6FVPNX5EIVw/Du2AUwjoz4EPDY9Pn2vdSGXaKV769hl1pHfZ
n9/2RDkpsZfPD9yNyl8jqkQapO9tVIAOwvn64ideCx9qeyJQd4YMI25KTaSAiqoi
70n4eX61xKqzqokhxm7GfM55GS0BWaTB/yyM/XinDMe6VoGjKWaxqQdfzof50Z6C
lMrObQ9vq4qgGvHtRwvexpHyZxR7wdF8vx1ICwqn6zvW7n8HLsTbE7BOTS1NTojo
Q6VK5cdfXVYTBqtLZVcj0lY5HvSTJbQHsHSv/jqx0uYB2QXroyPm+Zi+5mGBBJuF
4h2hNVKEflFz59VKHW7FhiXcAGvEMUAtq/XeUU+e+H3BsCt00TXLShmH25mkGljN
L7EYaECZnawDM7ggKe/co30BAqAOFWWrd2H70JnBsUpab8uxjCUud5ZWYNWD67Ax
qlIm/cjAWErY7DmTw+JigNNEvcjyU/M6w2dDXorgEK6mF31AN0vVoAJAFdruTQGU
atCNpkK2BUWHad0Tbwz7dIxZ7BayYPx/I3jymZNwFqDLL/1M7B3CAtsVO7fDa2wk
o17jx1upa7GLYSOzsg34zRKDXzHnfJ9uhEk/eF6Spi74eC+vsWiki1rahBRY74Kr
8zw5SxI6AIw7vlK6sDiMDSbnDCV8UOr9/MCJGpomEf+lNfd4uO1gj6WTzpCFrAZ+
GSStc30D9DR+W3nedNWWfOcJ98LzLhBqKrVplSuUKAAWnmUqkTygnbzGUBwnmX+b
bquW4l7v9M7e+XyHS34sjHSZklsVbDoxW1CQ+eiTj7KriMMo3YvEHVm+Wy9ZKwMw
i/k3cSWwZHAKMdR+8HPCLNioUNNvVkTyqIrc07nVpKeCP8xXdZmoRhfaK/9WPQFv
okywBq2jnxPQiMocCAtzuk9HKMjyUA23UWGbNtXxS2Gjb//3TQdZ0ocqJKMUSwY7
TJtb8yNA0YZAmuNvFOnpQjVqSZDUuDlzlqoMQCHe3laFdKbbV14uC5wAj/uQ19hZ
CuPH4wWZyRvmr022MZQod4+SQhMqersRnmjY87hqyxKZpoqIw7wZki8TWmZWEswT
tgLXiRqWQL8M61xdGwVzPoomB8OU2zzqGt7qG2nrE4akcqRqPoDilSM7RGUjieFW
1/jtbRnmlW4GaBu1yrZoCv0v+EI4B40GyVkN/vYl0NnC7wJWo24nsDT1l2w0gzM4
YuhRJ6CQMMO15x5ATiARTehY4PAQY8DUNyKmpRckKU+1kv7gHEBMaAs6Yto0OHKZ
ZMrUbHm6SqUTTOr9nmroYOIHAV5IZviyIMt3JEtWVd8vj7/wbVDPSaHs5yJZ5l2J
ztp2P+z9YLRVafUlvpxb6BUG9f3c3K0imV236RNiuNOzuC2Djg9YewtKly2RFIYj
1esY2KZA2tGGEY4wZS1NH92VVR0XC2+KWIgdZePLl5qLA4W5GYOtBnLjs5+qQGek
M8I9rd5slVXmlw6cs5KZE3wjdeoN5miAu1EH2usyM9jxWhZF2Ev7tMGEHwMcOlmF
HaUW38V+aNVcznZRBgjRvLffXMMSou+dbLeNixOeF3EsZz7jhUTfxh/mywkPaVxP
bJol0xr8FOq1vEvzTcxI3DguzjTQ8ffFfP42ilS4toVF2U2h91uR68+l35zY27gH
42k8HDThCm8GRZFpQYVP74JCEB5ty1VTxzbLoPBjM3L0x9HJg2ufhSfV3DUGfmgE
z89MLQ9LZZgreghCwBwaYhXbh14lJrDx/1aiGZ4XO4nggOviGSOtEdVcSohW8YUN
GMTYq22uSFl4u+vQcb6K2RJ2gIwALpcG03OJJEZUk0vDelNx52UK1Vq5lHR4gL+9
7QMfck5L4M0sdF5zWBzwejCflEWHepkmjjMpsW6jBwr8c01nytcQsYc9ZSNYK/KZ
Cp9Oz70/DJOgxCqul/tYYh8ELt/gOvSTrhKAwkmnMUBQKhesEKcA3zk+0OOJRA9N
epyIrHmipsleu9XCgO7MBPnfCGvNojzk46uesXgYigdqwNtHhtiBu3IsAyz9uraI
azfeFDMPaaE4I1DeGl2D5E0p9Dg5nA8hE/9C3FJaZhnmjAelPYYEm21Dzf3f4Azu
OpmQbJ9bpMlxiaeUrvzZ5EkEzZt0JEaSNnZWG8hljcDS+z2bv2gMAlDCxUsQtQlM
RfNXjv8cpBZJswUaouTQSdYxGAPHcbkgvLx4DiygaCIniOOcVzW6Ld0hsZorhBra
1JfWBLnPDsuHyJQnhM4B6KTCZ1qQ7cfrJq+T4OoaPDPrKIzK0yXyDidp/+L/DztS
llt6riwMsINhI7a2i+5i+KtvTOZPDnk2htyjnq0l6ovy9uueq+/7Hma/ChPtAV+A
s3Ep7sayYOSbkPPqZ3FaW0f79uWtxoy9AnNQ0hQPIWqKPqbDJqzjNRA2ZtP3QLxi
W1afp76PgR7+3ZN0/u4JSgzSq3CNOU5rreRPh++APL1EYygio/gK0WahrA494cA3
jO/QO2qEibBfAwwD2RXqD475jRxoG0Jan74FbKi4rXqu9uiX0fUBoEiscJMO2Udi
SKrhB22I8j2SgDG/+Yjf+5L8yvAtgVSDObynNVOR9PZyQRqTgClegPwPSZ0f1fn5
J2oMbWwgAjkloPJV+iTq6NXIGvG2U/mRPkjn3XhsI4ULJI0rrwOZslRtuN9n+++1
75c2maIcN9uXMLsajm8zt02bQX8tiX8wMLsjDM/YBkfFMaYtijDYBajkaLWJG9Kn
XBYkNl/t9N5FjrkuprAt/j4m9xPQSinMId9Z5ubyL5Md3sRGM4frG7Ze2RwoSWR+
cBS3FQAoE0XdC0oLWBaZBgycKx1TNzeX7u38HFWuFX9yZbL4EHY7Gwze4A1CbZdk
DxCDwnJW8Q+7zM55sWBTGc9ll1Urx9TPzROQmm08HsrkUtpUrWRFqdwE6COz0Nkg
Y0J8ZxsbKCnvSRTFoa2omz67EDjYaVJcOG67cxfUs7+jeFOYjqPG9jhrLzAI/dHP
sST+1jVqCP++PooIHhsoN7P/ZAMEcj3QWT20qsgpNW2CbasIzkehnRQu0Lr9sWqp
r0OlZqJXNsSCQNdqs4eYybse5NowS1TYC8KX8lVYY74VdecnE4OJy5hzdeodpAMz
4UYXllNr5M9vmLVzUVBt0qHZeE4WQj99tYhR9saAgULCGwqcjqbEtfEwXlQGsFyi
/l9JALwo/+xz3XTImHbnwrcVK80tMTUrJfbzuGx5Bh6MTJ09mBCMXrNeePXA1j1l
hFEispHzRpWE4xGjo+TFFD2diAB35+iX4XSFyir+XHerWDV8AEEFqzDOOU5XQpjZ
Kz6a1veM1eQW0cr0NQkbbvov3tFIcifSbxilPVyy73jaG43+CKiIKn4h5aBdITCV
dDcoPli92QchQLfyYcY3w+inwg1ZsTYkP8Y3LVFsOEDF4gZkLMzi4CHEtyt1m4Wh
8jqUeuN6XsGtpTjr8HE1bsYDyq32nRoSI2d7g1EeKWXORequvFj7xcDOIn89x0TF
V7L9eR4Lum8y9UM/7QCt2g8ADf3E3ESOW1nwZOZGcaUDQ1LGD8FdZWhmbpeUpbPs
odxbmO3SfkABc8zNxVIsepOH6Ij289+yx6X7sGh71sjythQ2Mur9dN5xMog4S9n5
KjZomcUaQIVOemc/nkAgylq8q8xPkLUw61b+jcwekiwnYDCOan5DjVxZUUYXQ4xc
rl4YbC1X4zoipQUJG6gahEzuzmmrKMC1ST62hf0Z/7hiR4tpccRNBlSLL4IqKzoh
wnAO7QYS7FH1G1DukAWeW58PzQWP52+hlSUxvhdrkTCg/ep4/Tn4ED8aMsudnbRB
vMImVvAlz2NvU4GYFnBJ4XSxdzmNFu0C8pX0SgasxpcYxQDHlwAyjRxzZ/ziYjMf
tAomC4/MbfiwrNyhze++W+kmZDxz8yZGLJipk56DnuTeM6RN9JC9hmu9vjRBgMLQ
ih8wVTdaJ2N0snUbuNdmmB3sKPpBLfzsUlGOf530fOrOap2jMmb6U7oAEuLdBzNk
DVdDbdmHqS9vmYoBcJUvHgSJlirUAWkes7VNJK22/blam5ccTCtT0UN2OQ+iJffu
gwmJgxAgDj28ZoJL5e8wH2XAmK8mQ94GDNW0+fQUkutuqnsRW0XQGtcR218P9aIh
zjUQU2BiNWvJVms58C6Xpuq+NhXBGCvws4vWrYfOIrYr+yVtzYZn+laTGn/nfcIp
gtjgPdWuf0MOasAAs4akhKbdupyVAVaDHACCpd6NRIEOx2/iTHh7ArR8ssMZ8C0J
3ciGLMcAWD+wJn6yrIdO0s37D2hb2+lqJ/NtRIBx7Ih5ycVU4XYBHeQoI07am2p5
VQuaB9zP+NsFY3TVW6TTiZqIN9Xd2ULqTG8+LwnnXworx91K0+zvn3JMu07GE7r5
avh0zknBiRbTNxl40ZuadtXJfTjrrzZroH9Dx5AP6afuXlVeGpAgInvzhk/UMZp9
GYxhXAlxAwwxSFkBGw1cl1F5/YLOUJ9V5EhP0jrMk998CfhVf2WuS8EEbQoZjEQ6
jHkxi9X+IMBS1Zi6yXvN7c+/r41l/WPeaVocxPIrnk13495b9FE1QnTDyKRYusz6
CvTC//wujfVx5XE16peStgv6S4PoJhiCn4f4Zy56yYZnT2QYS8rfu6iB/LTzngXn
1XbL3qGQyzk/0DtyxVNZr8FD6xzuqYLXfGDJKp6T0zJRutfPSm98nkg4R0YDMgQA
1jolU+KeBNsRPWIyWBeXNDq7ynagb4S9L/+Dv8YfKSRn2LtzPPxzctXtlDX1GCg2
59JhTyOOlZkU5UBjWrOeiqGoav092t+7R7cQsnJEByCOORyuqsXlkYQyypfaSO8R
MZudR7A3UeBWZwLymCqzg137PbT91Qoncnq2BIdhdcuU0+7CuNs9I5QDRDWo79Sl
yeZFgQuw8w4igdH67OE2YVjnBNaDGtID01pCi6KS1S+UufEsFzkmrROF+SeXOVz6
8dPXVGh7exTnWQu42WAa6QmnvgC92ZRDX1CFAtaNxRr27tRureP450o/T8pztItm
V0j5CTCPfqYcokHmgX4pyejtunUrPGNVnxu2HrUm5eyNi5wdZPnnwtHGmjDQ/yoQ
OD7iQTWjd4OSwxOMj+jrqb6OTI8QutlaUkVRxJ2fgJLgWi9hOQbqTsdxDHxUcelF
vh6mN73h5KT3uyFxvbjVqTPZZm+VfE/NHcW9IoV1Z2ZDgTCU29GLuk+rhI77rt5g
c8ENc0qBL2eKRcObpa/VDKejSf810fg7F+8stT4zQxB5fnHTzJXzRSpPOr9ZXn9L
6O48T/F+lCX0gxQYFWWWlZcH0bt+//+mwUPJ/TnpU0LVyr7plZAdtk8TTtq1haRu
KngN0MiAAoRlHPhAGWJFK3PuXA4Zq5bOusQc5AxBRPJYN069yFrB/cBc2lVUxQ4Y
5/RhJ3XbYf1xBicwujPyofUG9juxGNJuYOWmXmiM1KLW4FZvkORXWu+xalpDXI+e
1JtyxLZHWTjtlrina6iDDljE7pDx3+a6wMq9zhMcbtrQtLPLX4jqN0UJSlmrw8Y2
zx0D0xKHn0V+qFP1zGc2jDrrthUKoDitQJVHPk8T+0O4Rupn+q6U2HyU149ZhPeM
9Ym1lek67pO9b3EGIfZ2tQ4PGebN3FZseKMrZytmpjDHKEbcM8C8vsfeyAWV/lbb
DexyUPZVzQLKW0Ncoz30Qgv373tdE/YeAJ2axX13bqyQyoqSq1JyrhJo3Kqk4qKv
LTPWr3CFEAZGKEqEktmZFT6ADHzokytg/ITGswlwPYWfOrzrcG4XxpguEXaWbQ+K
unDBuZio9oz2ZKxPdFL0Lsv+Bhib8dqe1tj7QRgb6aOGnH/L0PD0+vJoGg1f/MYU
DH4INfwY8Bt07nZh6JSIbaSU9sk34+TpSwch/kPgCdg5FVVdgcaurTXbpswd029P
NeVw+R2DqrhViUnFad06eu7ehJ3X3mJuAFBCb5HAm+HYivVununfOeOCLb+7VR5G
A1nGeh2UXowmnVrcu6KPLdaO7bNxuLIGxU8dhma07+7NlBHHtJiL8L5SHyhisrxS
4nFuEL3Yq1Y3t7i4cY26JZ29L08rGF2L5MzeRvgwdp9kdEeRk0ldUyhZsat2S3CY
54zRN+Hvd5GUKgm6A0uQav3isJGt99QrQoyEmFV3VK3piaxYcojhd4crQbin9mtf
rUbeOrSNaQdI+d5EjInVhKAlHRAtrZ12uhfOzAfNzKKuloY1ziH1wv3od6qiePJd
nRQFx+DIqSOPPavT4OYY90NxSPO6iH4rTH9u8h+wv5ZwN3KEUJrlNmPDgqQ5Fk1s
HDG2nbH389W+CS+QqpI0dCstvjV8lf/cq9v4Zx5DdEkkrWuX8URV86vxg1Hss9Yf
MR+Q6ORrAtJutTRajR2Qpj1ZAlRlDBAjtJC38U9gEtYMx7erVdmdEzZ4t3O0Ku/I
NDwTCbey4VoU79ZSNcNwWzRTVyadke/8RGC+2WoQywsZv82xNUJnUFs2G0o69Kqv
U1tYd6Lr7eMA0vpxx3tbtlFjdMy9X1zAhTNMIh61bwQa+sTRRek8a/8oIu3F7HkJ
srifMMe1Rrdj2ytW3jg6o3oUvPq00x3LmK6Gg8SB3ue+miv90GjWQoYTWT79O3Ug
9mIMNmZRlJ7H5RH2MzpmTFgUqv7iHhhouFWYPVej6mvHeVZsPLFuEOdQBn8HEpmc
lkJzFy7WxNg9R6KEHMLrqirKkyBZX0URXe11XtISgoWqlDiTZEUXyu0Jm+HsKZKA
xeL3FSFd5+JbLTsi8lHX3j9CXDPfgm4kXxrBN18hGMICALB6TTeFOylE7ZFZZp8o
Mk4QOds0PIev3S61wb10IGZy4t37+d/9KGxzK32xkAh+wPuRsccKcHBDfq5Lh0kQ
hPdPBJnm/LnkgiC/k1ZgXqEoiDpt4Eu7E6YoIkueU/8yNGWpeea5X4kC4b2/mjW6
NeDXPGcDP3ua5dHTnoY3rsY8zTB+iAEuyKkD/OIrJkh6fwQuH1GFRlP5HBps6+ey
mv8lO9m/cL4tbihgQKxzyntLeoa5MWQnPPmZAZwTCMvLYz2e4dZQx0AggCYgkqfB
KPUQGgY4zp3oZ4ovV1uw1inACZdTdYXND7Y4yRE+XKVYk3WQbdnmkGN50VvX4aGm
fCJcwj3nChWnizAcygT4b81YiF88weLhRDeFlDS96zAYqkBBJifwygQGyq88UI7K
xq121kEUUvtW6FOsLKvNxwAu8Zs2QHMewVC0InpRYATaDNtUFakz+KZcIxgIolkI
+pWxaEJm67dCPPF3OFwv7qltCIZ0Chb8ES77nqQD5fwEggZZEDhAup0utrc05o2x
V8IWvgFy31tvrDmKT4iguydf63BKf4W/+4MnuJCZDrxiO4tgrbql0/B2Rr8wq2+4
HhGtzceQ2MfN9bqfvCuDlV40YsUUYj4FLkKRGJ/h7rjXRRfuqkLGxhTo6CUtKf9O
jCL9+XWDPxuNX/x8AUabeAt1ns8M3z4ohbNBVpkE5WUSNdbjFTJBABLWWjnu1JIP
XsTTowrIWvVvVK42wO5cacJNTLcUzRHsTWMldNHKkswsVSw9zVr3z2oWbe6ol7Yf
k1IsIt33MuXvavbGmYVzfDGKkSDgR6/0haHajmK64hwkAqyCi0qh2k5/eVH4H4sJ
Rc7P1S3VRBd7OTN4SMnG7vrljUblehLy0RlyOq0PxwEudHGG3XF7pXB37h6Qp/Zh
M/cLJJ/uJd68V53KWvKLDs/s4BRsqXeHJCGpNPZ3jog7pgOP2+h6PCOV/pcDhS9u
W1cK9ssytWV0z5wZELYtQheCS15xra+r2qCta9svbnzRHP/H8PHSAB0TIRKFZLBp
AkpZ7SS01O7SHayDeJsdsUurqMSjglJs+oGXmyRdSHjv3DRIET0KabU9QKubtBtu
xb1cpQ2o0moTbQaaKyJpw0LoIOhIVjlOAjwmEvzlftyKy8vOTqFvOV/0zqC6rS23
W//KKiCHgSG5uXEbVyUg05juC8LZku3BoThOG32yeksPDIXPdUf+1cij9j6oAIMo
yfBKSH9UBGQvMh9WZRi2IT0/F3aPJHALEnbly6MCg239r6e7t3d69mSSfHRqt1mu
Abwo6o005LjQvVCsZg+dBGmniUs1o2SGnqZPEfWcdFbBOiZHcQWWASaFdzOD2wcz
pzoNngnNe4N9JxrD2bXl6DdW0kexSPZDJ+dN9ApwP7WrCxqf6aWaMziGkE+RIo/h
fXNBv1yjOppWx3XhPAzVfC158uE7qybhIaQE5QVhedubHSAiFVRbHsoFu1w3tn4Z
mEq0mfogU5A1mlwQqjKHhXGi+HYsEGApV2VKgaqlDFFUzBdo3YPfT+S8hGg0bUra
eIB52CFQrvaXYpICSWafl/5lj8bQxPEWBcZkVcmqpUaBJBQ40nPoE5yvmktoenZ1
dBmV+AhLpXXVPWiIqFxMqtvQWUdiApzZy//i3PJmz51YNtYmLloUPIj7vA4xO6Aq
ywRL6nxWEbbV/VQqM0TUpJUAjxtyu9kwRDJzrtkhyJJQjHphHhRufOkSCc3GkKku
oJmQbYyEl78R+hv402YrnH5odN/M6DCQQH7NcCesQZM8xZLwBKMauLw27IpPvaU4
La6n5hFpL3gVqFUXqfMkPP/Es6xopgN9DGq7Rb+WOptyV45CgFhu5s/NcLDvsoqb
svapQMsImIRXUlZqGBgvTljx7OnXEsYy3AdvrmGlswti+cxZ2pqAFjjHlUxFp85q
bMVHYlwWHA6gSIw6eMUTQSAjVf2yTOSEu5rSpUtShZxd4LzK2c6sA3QlMUMAjkUJ
iqAHyeAgw49UHjcYBEdEccLdGkH4GpUo3hTgUoUfbXIKMH9kkonWzqAClgtbm03I
nIq5Z8a1vSDtevCGvevvCdnLph7x9Bo81qpDtAc8oh8DRKwkaR2tBY8VwbPzB6Uk
JgazBLQlZYvsGrjNM9CdXyuOQ2VndsBWwELd0zcqvskoVYcz3RqsrcR3kGJPNkkp
QgVUdAWTthmlNxvJ7EYrwygMk8lMNEnH2jpgXxSLZqvtWYglxu67hz2aN1pwG8kV
iAWwNKspB6vX8WwVB82zD2ADtTsMA82Ya2yvX37B7IrNZJ7piPYaHVWzYKzqutiX
uAP8ad8l3cn7z3L5cT7nE1oAcY5CQWJN8SpUCviRbLSP0V5UBHhisx6aF0b2N7yN
Z7bQ+25JXLbHR80Ux+vqL1lSfi0LgRQvgHIoEEPLJ8j55MuDhiAkpxkDh9dw24WR
Sz1NAFiO1Pr/BQ3yYbToSvobdz7TEMlyAiX74rOaG71GvWpAxSz0Kjr5fwmCjCHb
YL7CDR3kaD+Pa1SFpRbsaWMKV3J+V+MC7+iELVdKA5uu6wsqReunypYdQIcwBxbZ
PwNa6Zz/+S907i05aZ+cWQsgGwakz1WFvw5fIXhnsey2obtYLu4bbLnQTyqagjjS
xVWDjMunNHOVxu87U02QkKZFfDXIRzANIPsRxB2/4e3e/RylYoaEvYVr+b128dk2
nBfCKmKkBm+n2zFk5CQ0eDCKaDXgiSTob3n/zXBxr5m9qYgTu1MCAJ9kmZmCHqhA
vc/lnpT9DLuo+A2deASyxA/cb2o6hLCQ/E9n1XZNzQ8oU5DfSrrY11OmEGFS+82f
X7ZR/G6wzIl8VvR54S7k0CJJ85NFlV2MatUqWnmatp6NT7BkiXsAUNWqmGgtWNki
bmtiCp8CDXmPdxFfHULBWYQGJbSfQzLckvZ9qERbIOOo760xRqnX8OLnPEY2Kh5N
v385WrHJmHRpko8T6OSXduPRsdwAurCW5KTxa8lzQyc+XzHSomjcZL8W5Lw9eTje
OEH+w8Fcul7fuOqpQdJNdB97TaiAu9MZl4nwzdUDdTWRT4XYznsLJrYbXCBrL5Fr
S+V6xsCe32PuovfNWiBmYx7q+mXu62I+D6X8GTeW4EMJWzBTlTymhEN5mi+IBuFE
Fe+FgyYs7JkpSGu2uU1d5xuaEudr9WkZBPWGsmy9vGlWm0rEZItSO7Ykdm/H0vpS
HGEF7ht6kVxephiRRU7KAtUkzxLj/2nqL4bf4KtreP/csFxbLAm7GDKAjVTUm7BZ
PLs7RdW7OAdmq015uZwPinvNcq8SISvRMSyfm56sfYn8ejMNCzcOXdYAX2P0qmlW
vr21HkRWpGjm3dWD4tTf3U1hF8iDObygyAKuY9BTkryWIzWOEKns9DqzJX+o5R+q
s7P0B9u/a/cJKScmSXI4bTwdpV4ee1wwGjnqagNPVVEg8pN0/bVrPfP0gl0iUUFu
g4UmErWxJWONp+RBFtqWNyGtfMCLJPAhz7gxSTucbb38mGd6RKP/LLOcLXBkMVBA
JOahCSx+mAZUijAkVE9+ya5e6N8r/TbA6fb+HbrBlf7PFFkGXYYDOhdFESmtGqV3
6BPwB35M/9iLipR+veSem3545zqzRB/haHCs7iRQEmQW3Wqxm/wme6IRl+XAxmF0
M317zdUGl/or+4uVwFoyV5tbwb73a3/d5L0z07cNA2MkDzwGKmC6jOtFnUc/QzB4
uwTfEaD7mrGkUZxSaFfAA84eiF+JCpu2O+Ne9loQdJXa6WIJO0Rov17+ZdRhqmce
NPc+NZf0hsrzxf0xeD7jU9X5lz3+hJ8TNmM1Lja/zd87/2qg6V56JY8Vp2XFwJ9P
ST2k0O6CV1dtFJs/DdRuQKQAiG4PUjylJVODqkK+3TCFUS7IlhzxyyOR2KjiRQ3+
MfB/BXIlyNTHFuoNRYoAKHRuF8lk5L9VPYhkhafDoEEKDq8QsyeeH9EG18w9/lk2
zY7CIOkxscNcXWui6KO7sEKtcwIdfFv4JKwsTJ84nKZwTkQ6CC/IC5VVFDuDGaY+
0YCWsdU0siGeEYZLu7iQQDyeCRwlm4eJW8zVfqvo7lPTXoiQqoM25QpJaJCZh9Yt
qIq/KpEQoyzhFypb0Iq+4GinhCs4Uu4pTWQKoldPDxodx/0J65Wjw3SBs3KOjjv6
FAvqj4SoPq9dxd7lnqCEHBsggZBC8Xiux9XoceDPy52uDqoKk+/qpU0Y0i79u/eH
5T2n2/C6RCZJHRgLg9vvFO9EydOTBjTtUirHGt7J04NOek0P8KCW6YZY8az0u+4F
8PmrEuXnB5LqWEGGfvmCIdNxXogM7Kxm6PC2JkBZBtZq/eud+Pj2+hRs/rZEqJoQ
fNr1oeuczSaNHIEF+tVhBMkmzO7G1dJ3+zS2/eL5xV1UMjEFx1b+p1R3NmTMAj6W
M1llqqvlig4YvHshln59GaETUN7f96hecfyaj1ZS+0U3eijrspB+8lwkcdD6ZEID
tjrc1DGkKSQfnoAkjz35B4cP1CCJ0c8aWvq6uWjgf4/rdOXl6r1RmSHRW5oAWuzk
XTn/tcgYWNbtmaa3c9UGLKCQeYunyrEh2BdmT6U1VuSBsNAmGI8pnI3juPqAEVR/
GjWFaB+jDKR8tpNXAShTRIyMGp20coxDWeXRL8l0EavW1+4kdf9XPcxEvTTgVFFU
NsNAjC4eC0l5ZQMTED5oZX8emqFg11gil5xdnXB+UopOsNySZ8y7ZfZWNzgIXYVJ
xSF+qtKIN32wyVaMMWdnvBPZFTyKdabyHx2c+2YaJRWyMX84zClixSypfWN1f9uQ
A4SEuXnA1iOLgECkFVkXXk+bijrOkkhLr390W7lD4tfZX448lCkDv4KLQGO4EYm7
YUikMQX4aJI3FOF+GIvAun2V4tJWFiWDehlCnvZiPyyfVCfC5RL3DuZvu6VzxLx+
k/pOMuheblEs3j/QpSfdECaX3zoJZIvMHZhbJasN7S3ZIzjz2A98ffYMuvFHdQx8
FRtmbfOr/eJpBt1xXY4x6mEDKOwQYI8PUBbzL4K4m9BuDsBJE3bXaiathQthAL4/
M6w/gGEDRSraeFyFr526bquK2NhVHGJ+DYyGt1OOswpWww6m46ZgmLEsbMaNU7HM
Ep2H3XqBOKUTEz/L9X6qpNRm1Nqcr0DQ96b3HZblSWHmTVBeYFqTlx79hPVFzmvb
vKuP4M24z4e9lAAsDBurhBfHtnaeNxmNOgT9kFgC9GS9rvcXSA5UsNBFrdtrzx6Q
FeI+TzhVDf87z6qVOM5rV2viXqG5i3nO1Uv1dzPUfp7eYmq7oQpbwxG8Jkxt9ORg
F2q9iEIMd/tnRGxi/uveA5NIXiQ6w/vs9Y5N0kcIUdMO6IHnN2Nh2ZoP395FVmwX
YqFOoOyBRuYLNXDRVcuXL7mQuodEvjtmOWPCOoztmPRuFrUi4afq4iE9WKINMdvl
I281poPELbm9pd7cc0mwTBYtkNue02GhrWBHRPXlkf1DfGNgGNZBnJdOPNQ9r+DY
mCDd5JhZI53gBrd9I6WA6kn4W/9ROQJb+W/aOw8/sFHtX3NOKeX8zyjy7hlcD/C4
FFEnT9+7VYABuhhv8uf2lH8TgXf112vrXhQTsEJy5ugeASM/PRVvXO7k7072YsKB
DhzzAyW3R7txAhLpiJfGe+lbMJZkvL1wDOPx4XU/vj4J/wd108Ex1FwHHS2Nzaqz
y5M5JSiVJABi0BFaN628EUrDnLb4ahkiu3Dsfjvr37E/rB7K3cSRUqOqkvZabdm2
aKSiz+uClobRn7YMhK70HLksYFnzju0KNlE/TkdDwf6bCiMPfmAYx8n8m+KZqHDS
0ANqAImuuAGRYGo2Ov8UQkcniBpoQXRgsCV1roOcpALYgMY23IORYq47McJlKh1S
3y40aXuubygCGvvidpZA6OvsTJ/EUYy89mEnm5aAmUf9fU/+nrivL8MjVlUrwZTe
9gyz3fk2yxTN662tN+5pu7zjaGUmecj0P1w3kYzQmRioW+y8+6nX1CfJtKArz1it
/UbPKa6iAZVP4sRBMy4E+2gShcO5FLKtvvPRsjfOxA/ZMNRBP26dxi2/zlL4HYth
PypNzMnA6pfh3lYZwxAVgQvkE8AlatalCViJjf4PjGYL6iL//Zx50a5GroQbCa71
DU3K9iV/CO8YnBGiISMQeje2osZkQ7iM2XrrqQS13LQWRyN6rZlgbutgJE3DTijb
bCRKSTIAAZbu/0SJTvWfu02G6DgChl8ON87zW1Soldc0VE1326RuZ36d+5NwOefN
aOsRbv6xsmsVdvs7e5MwTfebNonYi71nKUkb2YLo5uYTP+My1ywWHJF5TthBC5YC
EB2DKMVOzot8Ol2bWMST8EJ2N89qJwFMgGZS/HS/lXqyCShB/lbJQEAUThQvJsPA
vovyMvLm6+ssXGZEa5wqnrnEc9ENf9hbUDiXThigkNXpXlNR7TMyFSopUktKSQy2
ZH0yub8iYJ/DuWpZtcLQr0lviPCrDHVS1hnB2XIIcoEl9UFE3uFmDNOAxmj2zxjO
XNJmnjDqIsG+yhfherFIYWFDEB68caJdTV1uwU0Ic1QXZNT+s0EcNkqbkcpL7/di
KnYZY6asDNzy+EsKojqL0zKL8rWghDl7g5ZO7+UG/yDOAfYXopneRriqQAY4Jtfw
+K+veikCoFKTAEcMcPaAQeuzkMcMdP2ck/C5nf23U1e1Dbx044mCB4gwh49Ly6JG
pP6S2yb0fM4M9+TvozJEcJHClNLbGcErKZa2m7akgJVikUCWA7w3TYdMwP8jIEiA
NKfnxrzk+DZry6tioW1owXg8kU5VdidTVrTcjlYD3f5tY4+qplCgO4SsJikvqaxK
uQfhR2gohPqbdHNccFKjia+c/y8L2MUHN13LPGJWhP0C61+kW+lDuZaMLXW9EwBQ
v67+5e9EuT8jdzZGKJZsL34krrb32KLya251Qw85feYEhmW5n2tDa9PUqFIapl64
N+b0SsruXd/7H44287ohjp3p70KGwQTWcpYT0TTYC2D7ruWEwujzk51u63GjIVXK
1de9O7SBPXjzw+UpQY7HepVj3PzOePKuLDhxoLUkZKg6ZlBV/MZxgbEYdPlv/oeU
bIMN4oMNQSHzKjPsyPOtEpmdPznbFWbsIEkQUfDK+Vz/cdnDNAFeKJpUrZMePvz4
oQ9zGnRM1E5HhMS6i2me1gY6QMBAsMMk+2XoIy0rSSo9f1En3qGEiPluE0ut46a+
ut4YfrCvlnTHCmLXTWYjBN55TIG4DqX83WuakU0lACxiqQ1ycgiJI/xIanVqPY9s
Ov/96iwHdHJ+wzRx/vILlpKCvG7AJsZbEO25+dLcgRHYNQhWJVzDlNbLs6DDvKnB
lkHgucKhRO3qsoo6HOvj6FKvqxIBN64L3jTSFhu7qwt/W9eXjciReehBkuA0DUBH
oC5ATyrJa4/UUrTJslOikiG7g9wDr+QTQjGCRZxF2Q+R9yPXv3JBpCOU+QAoQZBm
yAOwbbi36LLXG+pbqB6bEKVp7olwdw5J8unKNO7Nw9jVmUsUqL5nvH7kz19QYlGD
BVKoUjlKVvJwpRIXesS2nbipUANr3GDVWbJjqZRKeMG3TUN/eivl11WDrDe5DSsT
VEKZxspldSbd32XW5ftKQUDKWS4fSRMBEJgf34BFeTuGxc2oU/YPEUYD4Zj0wKxa
38Ib5hXPx/XlJaPAIR6yOrW3qcnY/3iDygrtkVAHtB+b9z8bpVQmQ8wci9a1Gsl1
FgzbszvKuDR8GfyfothwvXi1dOVJgTDTEh9rDOtvVTxKu7ietHy3JujwKICcU1er
jB0UtEQqtTrd5NM58AOs1i9VgJMLm4Fv0nXATGXTNtl/oELBG9/zsDFWqSJf+zeA
lgwN+Q/jx9fWT+rh81MRCd9hkLn3w1hclB/kN5+RkZpfD/SWPBPGE4iNwZVaeN+n
0iWB9/3/uVD/5ka0c/ji27eztv+3JgVROnVcZzuPeiWfFBLF+RsLXVgQv0GI5AQr
Po217dQ80WNEiYQh0khUk2DKGAbF9u8GAZjBbWKDvkmryn75jPDIIKtAEuBXBlQP
YJ5upuIU+wm/Y4D0XxgDH5H9XKcYttF0pRHDEsF0aws/iNnNcs4IVJvc6lD8YYDi
qw0imkJg6WrautMjwegQvWfdfr3pa8gvlmJHacDXq88cCz77dABrvnuNgavpntMo
9W2ZFLKatN+vuCyR16hLf4mIOX0NX+oOSz5LMRbdD1nNUpzOxg1waCcSD1O7HrFm
CQCMr7soQttaO53mxXfbHYgZ/xsqrEPfBE9XkRjSEc99cHHrnnI44b+A/YvIPYxr
w+nEOPwtpZZRNBOdRSomKv0e8VYOE6N2aSBQuPA0o82/xPwBWjJZRmNJ/s2YusMM
WsXCFvflWgE94P5EM5YrE0cyKNSx5c7ncgPOsBgqCcZrLACf3vGJwl6OX0uhU9Bn
jIFBDKKG5bS3KLcutZD4E6Bf/xDsE9SSZ3JKMNKmTZ6dSlj2kMkw2WDIGnVeg3vx
CyaWlhJKxeiUbiJvBrOEiwr1oN63QxQVUrAS7YBHS3/to7fnGs54O9a50KUnVDt+
FIo6nS7oYzZUCO+yimZBI6nJI2gE0QGAQOI38FcqwNDLlA3VoSH9olN6LQWcn9G4
adh5r+c74Re0JgE7JeuRSGqLgVlJCOTtuP478HLf032fgk48rGr5RezuTPdrJGa2
P9eo54oyO6XDOW8rOBQVX8GXL4rID+7TVgoMlEorq7lrMopts1mMOOttmK/I7kD7
ubsfBAgTF1SHs1zrcXI1TsRUJ/7qffR2Burcarrk9j/EL826PUnWcjdTEWDqUr+0
bF7stUtNLDDG9iP/80Od7xzkTotJBrBsrBxN4NmOsiMIw9rLqBipWmwgvOznjP4w
qpEQOE80tFJsL+Lhe/wRYmFlmNleAOZhgPKAb6IwVFmke1j7SDmhre3Zi8KqsIn6
3b+tE/w3RphUL6SWa7aOeY9cl/vuK5ktMdjQpbtrPwBf0qXx6IqC8o6N1CcyMv+u
6V6K6PgUkv0rYSlaNkCZY7aeRNFwU/GGoXqRnvOGyuZNGJYlw8PF6+MkUg4RCJoc
BfleVkVMG9qz5+9f5xX55g/aIcuJyjdfW/tugeYnb+8AT0McdirddG7Jm6NCbLld
KzK6kK1VNbCruGDFl8UcTm1/57G/wHy8Q1V+5ql5wLLXbhi7rvoqVODpP1bspkHb
gNUTpWwbXHTW+jwr9oAd7cPPc2rvKlx7QQZ/LBEi+76lN/dsdbJlD+j4l6IQ2Wi/
ZndGh1W6IkmmW3F2uqNqtCrLP6Xktd3N2FpcAsRqMkO1ZMCzRFiSnZAmSeWXJkup
AShI+T0Y6hgXbiwAzU2ssiVfPUJCCSnLwtW/CdM9g7ZFTN6LIEIvbGbD4S5hk/mp
rfxj5lois1pDp3KEpIwltNh09cQ8bMoBPjW5ExqPmOIui+wYlNmEf0rt6AOL3RHr
eqIRnTmOi+IvKd50A5W5N0+fxI3mFAe5eXBUNqXrGeaZecPZa7nlRwdtaDnwySXk
Taroex2RHAUF1iMcF96z+QdcpGKQlKrsHW/4eRk5vwFnlrySOWu69qaEU4Apz8tx
DCqQjdaq0IRLFJb0LGpD0EUoI4dkF4c0dvLVaPM7sci4qnwf/wyh79TUBq5juK3o
56hgz5fY55t8NZkPmq8MiKBmzNopUM/V5GCV+4PJACE8u5qu4mKDugQQyDr7cLry
OOyrYj85TkXjQq+jx0pt9n12WHc5vJnEoa3rS383gbhxrqfX5bBy3S8lhKdI2abt
0dgdCpUyFEl+JczFyFB3AMps2ERdxuMn7uC/BoUzaH445ucD8ABKzE8ohG3xl7pF
OcaI8ueYlnB6E5CLxRmwVakWVau5cx8TdwAkP4j8phh4VwIkCMFMmkUvNxgELB88
3x/xL4JLMv5onYzdjyHV/ZAxqpyH2knuuVV3NlfRuPbPtn8dwDGbo5+jHJGgSAku
F+PYtAFhA0JTT6pQsImx35sye1xYt81XTK/qHZaUFfnsB2vYihqqyEEulFa0sNJq
raRJx0aUnA1zVjVgsQOkChEQCkydkSCzV3CL3UcVHuBAe/pAm6rnmET8UhSr4Ld3
U44vowXfSgPPFPmR2h7jG18tIbL4NqdCU+vN1WohwWo532wbk56NIllLnzXttwJ1
L3Dk7T7bjwUMt4KAjsX44qEFAdi/Upd0DNnstyfc2l7tkfKONZiCZvTxEaOnV7la
xGT7I2lJ52I/I3+ekTy+PNQZqZzelx4Lta1LOvkfHbAo3LPtgVG4g2ed2LAzIoYW
gtwPq9rEyiOFfdrYJfvDXrExzk9ncATL0YCRLh2Pm0Zpz8DZK8VDnHNa3lJEaZPJ
gqd3d8KGxriWL5k7u7ukoQ9rNVRJlncMNQWcLo1EmHUUg4qbT7eP3pbI92VGzLSO
7lbti7c/9e9Y3k/JXv9pbLGclSgmirr42kFgw7pvRoAaIa0EsA93sTaySMdg2T1Y
m7H8563ECFdVUaQYGqVZRnRkJlXMq5vKerClsUKHZOIeVtJ8kh3rlLXvCmYEW4cb
wLHNrLNiH2K2ebWPvB5SHYfxI6cxJaimO/fBHLbvtcwSo1PbvIVudXzGOS9I34oB
wDIyiMHRL2p02kigGVJsPRLyWz/swmJhvuyDUwyDB/HEx1Sb/xCH9izUk0q1obj/
Jj3UVnxc7pAbs/yDJPN0zIIgrM6V4RFiQu3aGl3YguWCREOryNpVPfFfHepgZbjG
Zkeqh04Uc5h8cyMrln/+yMr+psUiq05s0Cke3ZZ+fBmsWeOTvRE3OpErFOjosFLU
U8erSdZNG2afGaKxR8AaWcZejaRk0PbJ8qvK56ZPjkVEpJZLwmSqPFRwiAZXT5Y7
5aTRKOE7rD82iDj2nguRg9tGyeuUeQmaKaAARrxqcCk4jYPN9FmA0gNFYkFr58x+
hSxrnxPARc5FqhjJvp6oYYw8+IEdSfx4Y6teAMECKTLMXU1qwGpR4p2qUnm/GjMU
1R6ntrWW5p0fSUMAvDuTTEY4V1WnlmKQ5rhowzT0d8at2W0nrcuFQO9O5aC2mM0p
BBA/Q4XgQ0Cp6uofrUxgzMDVI+pvZwCvxfad+QiBlMBa8sisabcxebX8F+XIMisi
5jp3Vudtddlh16YAGXqolQCEtfcPzDjGMi7MGU1NOG3ItM5abFWscDMLRptP8luu
omecdwtE4TVSwfMZrx9uJ7q90GcWae5m+zZCCvDmtIeq+LFyOOHnAMZpKp6uyw9E
Z/G/B0UAWODWehfZUyxTE+mkdcTnMd69qh2Q1+mx4sJr9+JLKNZuCkAGWWh2Ijo/
+yrIIg7YhtCnwFklIrzVtgFS8PfQXStMGwR4LJnwA8jHnWb6lO769GlC7RgFe4TT
MBXii6yEfeVy1n90SfRsIROzZjc0T7HsNCDdk0BbztxeSlc+XExbCMIT32XLmybu
CCdmIqubOUes//TxP3glPdOtbX/T0VfFSt+hUHew8dYPoNWqjDOHdGN0TornDAT3
auTU2lDpT5c3ZzI+6fjlNIjETCyLC+4y27nZpvJ9AGIGhMw3SeclBp0sX5HEAh/Y
NeX2f+4Cj3uBh6IYDF76YiQt2H06RprYjGAs0q8sDQLui7sUAs+tQr/YrQz6bReQ
nH9uZ2hx5nONJMK7LSURb0s5V5A/b57GxC7+FQ9b/u5xsitP6X2IVKVcoQa0v5LK
r9XvKvPKo4fb3BDPDuVZxuggN93hiXYYoDfH4RFO2MmCOiVTqYZlk6X+lhvaEhS0
hf+jThJi1jK8mb+rPGWF+d/35YhAFyZ/BjYZbwU6jfbF4DJAusLH4Ze1ENFQzQGy
dBfEMvyaGUAh7pAyKDdHNmZC1ChKFXFkqZRjayvfKoAOTD7uy3lGtvjMkmWdLp2u
XKmeEx/TqOM/b5GI14AwKMMUOxxvV8ItvXbFT4y86nFqkP6Z4h+vkkz3340l6xWP
zivTCH/nRGK5pF42kt489kVVG+BpU+YC/qvOC8dxwR4BIztRF8VoMEErl8IW2I2d
1RzZ4/6dlK07jWi9SoTdgdPFub5WQL0DQQ/9wNX2Fo+0hUwu/S1UlRdxqkQuS/1L
TML3v9YPLCv5xkB26gR6g7plD71rFF7rtWvPVifslwoKVTOaPot9gLBSPM2fHLJe
umHQ43GdQlFHnvaSnHFE38Gtn03Qhd0atkotJvb7Za8031h1BJFOWzFyZ8BlFtk8
ZnBhGV+1wOpsuVf8C9aEVU1IQC19WJztGS69PDWdUvBp7kGSpTH49qP0y+uO9sp8
qZh0gvnGA+OB2PrgFkDWZABvi19GauJ8Bxodmfe2cqgGKAOenmgwnm7HGpiIyjeo
AosrxkV6vxgxN7hx+GwsPGolTn1d/06AFERjaJYrijXMqJ8wC/R+qVdp8XML/65W
0ZYy2ioXrGU+tvhQqNgOgXkBDuy7dfq2MIiCVCQ+GcZjHZyDwlWReKIGM8IU8KAm
im9+e1qlPrABLS1JIfq/puU7DAoc1SxayHbFjaP7my+HJIoVHlPEdU5V6DbFSYRV
2FG5er1xFjpe7yBzX/rCXCbvKprPzu0MzaYcx9k3KVcoYdMGnF83ACBJNNIxFxff
rJxaeJm/MOD9G7IDdTtAaUjxP5al70tkQXSFgDE2IyZ72SNxmG7mTaxOuAbMS1Y+
EBHf2hr0bkY9N/Uaa0ZbNFtDspsjm0ssaxYB7ky5er/s5nTQZGEj0RO/2x2QGkHw
uiICzhBKrzUys/mcvkVnsCgCp2BAimduSVA1uJe24eYtyO0PTGcD+1gsO4Q4plqi
DpB1gUsGQCiIiL0aQiQzMxzFjqUhirLMtLLEiuafAObv9ncXoBsZml7XHEZNiaVI
3HcnltO8zjYDINTUBF7H7rIU54KwchwyiYqrFUJaLLg7dsVgcJcrYNXY0mO8EJyF
na/8xzVrhcgDzBGvSc1pmFtIgrL5hTxqUn5+RJl20qXKziQKLIbHnq5iyJVkEKvW
i5uIxqlIyRKAmoqNICs4wq6OzHozTOKtuKRzkjkhsz1CX7a8hCi/nGuh10c+TRXD
LDGE/zoYOOun90SRWrjBtKtbxiGSJvZT9hBg/hxiuxVxOKRQapFaIIKFCNJoZgJQ
i/Cu1G7eyMcAkLQvPsmij8ItaRfoI95t3+I8WJoF2AkXpRUOX4+k2RBiGFMf2qR+
Axla02zUahTyZLZF93oaJTzD8MOIuzeT6zuYTRk9sCubw3uuQxlRgGAh7bwwOtyv
kRxmZttHY67HiHLOf7SSnvkr6lk9UrYbRt3U7cNr5IBf4riwZBEUicnY+8kb/Dyu
jSvPgzUhNl4laPICZtEysqw8LbJLk6AgWgKcBj5T0SJhDsx4ix+PNW/mmYCtG/FG
H9hxlsoAnhOIi+0/HQpEi0UlT4WaKS6HPm8B2R4G13QKgqf2dKKoaS1PfQcgdSVK
VRuXZ1hVyX0Mm0R+X3MeSIy0FhjBnSSDYc8pFC508Kds9U/LhnJ76Hifd09cOPoL
lw0C2XTefKQyjChlvEbyPOHtj6J+HYisXHBek/e6Zu/wVCQ+Y06Jt7hVOzTJVXG0
19keXzCtoj/svdxsUY2MnbYVNy9T28T6QJaku95qpKLmWq8pOBE03OTEzJuYWuT9
subkmfobBVOgIVAZJT5B0h9bVHpXDFtPyuUy4Nqw7m2nIrM8mjgUCILXZ/DAkP01
setK1ZMx1qP6VhS2zkEKWlbRs3c+H8M7irhCw1THMA//9yAJNEKTglvyL7pMO4QA
I3BGg0uIKUVFRVORK/XvSiGUZeClgN+OofCjJdhfgQA4HJgZ+2eqh2TVASd1OfQt
K8Gg7D5i50EGkvGdmzX0uXFXwndPSikrvlKLi9JCjsr2/3M6voAe3xjzul+4fY4t
AjVXNRGAiNaK95hzKhiQzi8iVcgnltW1IGf87DSZQbduAf7N32vYrM/fxZxDIYeZ
fgiYpBA6ByegCw9/1uKZOar/hz2QIlElPXrVXgZAYoI991FfJGuX4UlLLcC7VUYk
e9AdAevEdjW5DX2Jckt0QAPLwGeIURAFgE7EGVuCqqJvslOKRu81tS7a5qPeludU
D1MInDcVajRnMCtMFzDxS9C5KF4VvGkUq7TlaYSWPWPt0tE2P0YXilAnqvgbyeqx
Rw5IG49ZKPXKH4urnj4/BYDPIkYxbt8vm1xqkam9AUpnugLzag4LhOyAZ7jR2yW3
XHWmVw4zM6mem8/2JwuDTDB15Ft9z5jkVnxCca7v/uFvbQuuWQTBlIC/OcWWK5CL
ke7m5h6rjSauetrx6LKMSJOzYVOUhD4+HqtPLc3mGve3CQDK4D+LhrWi+I8JM4ct
mRRCvf68x7r972XF/cf9Q8MKxhw6mUWiRYYjNfuoCCb84CVtVHABydbHU30u9iGA
R0FvPmLAaiYWv7x3ErMVR0LS6IQLOAt0sART7lNdgJ4wdqRQarKTHT51+miuYbld
kVTY9p0z3KO3FxTgOP0fUSS+YlaaSBfNIuNI9FZ9+yqTcHTBPu+wxZ65WJLQc3sD
c+HZaw96KITFfj6BwGrhFkvzoNNPysF+OPnPE/BohREq3Hw5sxAjnUMZjrcO7EB1
7wT2/5qrywCTO7LF4Qj5l3D+hpoGkX2jW0w1E7Y9RUSsMCBciEa+WATCzRhamCgW
oHRHWkeLOkBVyiEM7HSkrUoTu92TPDT4DuuVbsAJDFKTznScX9iU8y9RGvU6TzAz
+rb573OtgGtyK/5erf5PVlhzzmTmBd8VVNXGXMHx+hHV2s4yaSfVjTD0tSwxIBeP
Ix+Gg6eQHicHupYQiIa+A1dGi0f8txYvO6ZVtgPbh7UVp568S2Lny3kicpo/QN49
SJMyYFQcl4StGdXlB+7kdNGgzYZ/a4I1BEsDNw/x1vHYa6OMIRrYx5OJNtqRTC8E
elEz3XAXxyCkBFWPc6I/4PV+Y4pcUf7WzyWJEdF/wcEDeK9tGP+qzZqx+SVCasYq
TviMSd0pyVHO5sIfxNBXT7Tsk5rgyTY+GLp/WII4Ic2nxhLUgte/64Pp+mBDovsa
sRu9Qib/jRHi4O75+rC3n//GYXaRzooBWCt1d45NR0jCCQZuEa3aN0Z1nSvoXTOe
2FGizYPXCJi7Wku/MtYY48HXRaHt1p3v1bxxItY/XjdeAdxgfVzI3Wrnm4KyiFjl
g1xRCWZeVJyXI3pSEzwe/lgWrBXCjLf06VTw50gLgwv6qOt03qaER5rSDhryxrFd
L8eeQeAI4A8LlHqSP4Y19iavghCdqDGs8jUu9mIjwvKGoYb2PGeiokN+7AF0eDgu
8HdQpNI+Cl9+OS4wH6MnFhsIeTo2yl92nM8XgrWQAZC1Oy2KO63pS6YcPxI3Iq6I
KEI/FHiE9GDYTCS4a1Dd+JuRsUPqD9Cdlg9STFbHAT+g/7A+QyYo03bq/rEykcYC
+EwqsabfqdJs0N6N6rjqzE09k9RhVu/ZLXOI4R4pXyhi/ovEbFh/wcFGyuvNxtu8
+DwGkyVXWa1QaLp/ok4TduqBxNkMCQGJZ8jtEjNkqWFWcFWf5GJg/GxGxZnG5gOC
Jm5CHjXaUO726UjmDhZygpiZtPCFF6gSUUOdMfrmPQTFFph/gX1/fq6SGl28cH7W
i4B+kRBS8aa7qJGxNgsxCWGD+mDBZ2KqfK3AYXJ1iFX6WWWLvUHb+ejdTp+djU49
zvZ2xqCry3oinUR4kkxcBj82oCh5THO0AGz44gceUreknbWBL/6Pno+ggndPreLP
SQwPXS+lSfgX+IjdQqwjHF+Xr4A9gnER7omgUlCIYjdUaqI+spwuAKOx3k25S/F2
xOUqfpVx7j0P+Sq0klj1u7rZd7+hd4sV3WrgWfQdDNQVHzOHQB5J5EOse9JJ+dqA
p32BxPNQL+sKwd6g4We3iWKw+kAHR056Hgr87zKnMk1YD9hh7BTLjK1esntUvTPc
aeYn+7ALvToiAO/zjCDkXDFNVl7nWZbg6Dv6YjMYqBe8POmdmUCP+ihOK3k6DM8b
JLwlMKnWNpJCC85Wgm7PD9YmvSKpm6udxhSmXcpsE0p1nzYNDrM/0dkT7E8srcqf
3BhUjYd0Y4JSk7FJUCEgtzVg/OWxlGLr/xOanKkDERUybfcxcF+cmpBLsTl8cd0F
sCCE3x4jh8YdPaPAvWVzGEL2zqodvmPqpAnYCA9pfz53n1e3zLsFgGa9m2LL5Mvx
OWbOlA4q1BuezFAqBM7otvmetyoynoykrzKfMbOKdjsCsF7TAcNaVy+5prIQ/E5m
aMIxv5gjvUCX29/ssyb/5jm4RtRcygVImYQNQghUtRkyCjxgc8X3FK+C1yznWZ/7
XJGqxwwP9BRNspOINN7sDlQaCcrmJ2yV6CuvTLojew6APFNcrjhcGheu8Ukd/rgv
nsacAQS9nOuXVna5srC/f7J4qEpN/b3OhIZdHyDyj1yqh+taIYi6SPyuScXhAxZu
mqruSDBkNdhDjhxgZwxrjAi9DwFFvCz16PgK6nSN7YDqKC2pJN1GtcW9QowNVs5B
QvcR5nFXebFhZG7uYJt8dc4USydOfsevq+ecnMu97Sur6LHZYZFSqzTrJI/8zb8L
IbNPCg4ddpnXgpB4iJOjIseWUthJ9gFgsXLjmMZQVUXwPTi6dxfrMwn/Mbm5JcgT
WYEE0PN0wI544jlHjZgBlsAmTnf7kKmNqLcfZw2X7me72Lp7OlFoUFZVxXmh+pRq
l1ZrGx7ZuVoBOLdu9UvyeoOxKlBCHkhFr8+8ksMdz6a3c3LbFg/ud1T8cFCkZFCL
GFjrE5GyTaJvKRuOPLqLsL9bs2VejDW7go5z/FZ0lbYf+AB3+WiYAACU3a9eQVhX
jjCzgXoxW0RIxuH3gNmUxCp2OX9H4d/pTFrFhuqBejtke3xwN5wFQLv3vF6Od5pT
H02YRYbodhtQDNZZs0rOFBLeDl+/7tQj+FfejM1Ak4X7eq4bLKgwjBLuI5I1uNMS
8DDcIvyElGjWLow80qpbCK6DPBE4SwFGaPYUiEw8IefmF1s6nWLC8mlaD2LfxtPC
wx1/rDneif/lY6FyJMsNexfMuhbLt9LzsU0tHMK0TozYGTTvfKRRO1tFrGNRKfF9
iUsL1v3daOJjW/0L0WDBGAQK6N+JD+n3PLo1PfcQqyZj0HAFhiGZP39QOpCaHFmn
of5Go+mUJjfoxaYBE5qBSVHAlitnJ/iVMuX/tcw4zsdbZrzBMcvnLg3Z7SH9Hchr
rnqUlC/MIdYnhteyLHSp5dcyPrp9eaAsENMKvfqWdat86igz6vxtSpapYKYXxTdp
qJupXPObste4iy8WCQn7AzY/v4zyONdYVlBeh/m2cXe9r2La/5nl+WKoQyCG+lJo
vFAE57HWvLCHdeihzqoDCB+PNVmx1arfc63FMyq8Rz5CnhJTSSgQPNdNUZO2IXwv
J3dpsLwatPXvpbbHWsRNdLsnleXEr3p81UeNgOhdHlWDsHUNEItP6ILKxAkgewlJ
cQI2nm9GrCtw4QPRWfnp7ssUvzZNgNKJrgujxJwoDcPBhDHs0sHcRU0vrvv6qYuD
qiI1DZx6WzlmCAMzr3vwRDQwgLa1KUFv00wYazL/MHEZ1ixBebPjTLAN+hYtyfaM
dQcdTcF72z1tNmtpRu0nrhIxH1ivJOKBFgVJ2CvXLakl7r7/IJO8NVl0TFbafvbb
C6L16gCRVO80TdMqAGqpXtO+imrbK24MktggXFlsTrPH8lgFyltQypSnbeozkXIJ
iG+4LGquc31i+6OmWfSl47Tm2Yc4+e01/TotlqrE7r3tf1ic2O+WxvsEHg9U2AL+
usKoGCEZN2zCdB32cDdtf2r0AHbUZxTaaQo+pm6qLvdpUJuoHbPDs2BR0IEtuZvM
64oWNc6qis6lp9cFQKgl4l5m2E9xo0MrbYJ93q9BpmyHTDQucc4lDkw/+787cSiD
z/+dotHQjNe2XQVafLfwdJS1QZKXwZNJXfTGRWLsSJTo9KXpNsarD1TZy9yVG7ch
Ut1P4F5jjrQ9YqTpe8kHyOsVFBo1mLuPkiCvh7Z2bed9J/ldXyZMXiK9BgvEELmR
+y/DzzrCAIWWmmoFHGVZ9pcYiMf0Eb4Kc1s9Bfjdf2YUqFmfvQYfsl4yTjwvHZBA
63boq4VsPK9v2b6U3SyUGq/+VnzhXlCZPCeTn1Hc8xyZRkSlegTsOK8F5QBgkRPJ
j+TVqswk37MKuTRDnReBTrtP+CAiYEAIcWVM+BC2v2l/n/jvh9I6B5S2QXBJ+g+N
y4lx9UJuVhOX23q/1UPydyv1kXLN67z4DJoQ1tclp3pEDMZawskII17C+526ITOG
J9IEV+6AedR8EwJYBrDy73tjlTup2ueaOGwNZXQ9sMWq75pgDHJRXGwieVohjW4G
GbZW9QBCSkYRke1A/5YHvf4aBYz3v4fBUH/ai9XwHk5Y8oB6imah4SPWPQjclvBq
3EaoOkUnp2qGZVdeumxdOOiH22qR6RlRt0tge1upNxWm8T76e733efi7w4DppU2c
n/jvGqspdqBHif5CoKlXO/I5LhJHncFDWRKt3Cjp0vw9wydee4INJoUFix5BKclh
cUWKc93uzZBtp1MUe/cSYIHiDHs5j0CNz63G+sq7/WShsBX8seJMu+a4XooUEF3S
5l84LwVYY/8oO7YpMnf0ObpcN+NY4cg1EcqjLBNtVGlUE9jqiPF84t4c6i8uFbi3
lAPYqebtXIOekr9day2m2R8v5kFs5/Z0JYbLzS4rE9evTsfoQKkfTCmx9o/BUain
FAo6XHwW/V2+0tUQIzOLezBZ46tRNbbt+W58PXUc73tp3qQIBdEX99gf/oghF7n1
p7hV35DVzDGUpVVLpncTJfN524YYNTtGUwxHzNkYA/5Kysskvi9l2IaUhYW+RIY+
0KfcBwL8iSV4PJeIC2FY528OXpd+7gwBJPMVgO3J0nDIHS0ewlJU7HVEm0cmuqoR
pR87Ij2RiFzpfShc3L2iP5HcWefj71b0hhs54hSQj9DVpDeeOE2xgv8aSEJDQP/5
XRKGNXU/pO3pFfmZLRa0BB9eeP4M1Sc5y495z2pEXOZ2tNeodu9qEaJNnK8YZ2oc
cenEKmynZtHBu2m1LF0W/3Z52NANFaK6yYzUmfi6ZZx/E+mXHI3VK/mtXsQjrm3t
cuhuhZvs21n0oi3kZNAc50rTqwEMRbWOf/xyKNclrqNxBqCXXCB9y0NpwC7DenHM
XeztgBcn24ul9wPWWTg8xloLpaKszAu/nk0DfZ6ACqbriwTClF9yMO1K3tUBRvYM
W9nf2nilVZXtPWo0EC9RZUcgysJmJA//HWdNgWRdz/gxRA6cyQSdF3fYQPS9pT6j
m01OvPcnbID6Wm97IUz7t4qkpM2wP1hxZWRGWG1ujNPogh2ciAHLImduZYaGim50
rlNUv3xO7sScaqAp3cWNTkYU0S9BpNYh0VuI8hZPU0lTFdTpLO1xFMUTNB5K/lwr
Fuqv3ZhUQNQAl0bHOrZPDrnvQiArZAd5byLt88zRTq/6GLcrz9YI7tmJzEAc3aNo
i8ICgNE2bsF66a+Y6CrsYDaO561Ny4CwdlM+S6BPKzZoUIShrfxjg+cWwAj8B31M
5+Djfdif9Z6Elmaemf5FUsEFd/AcJBLmfx5LGkn3qkVxZSU2vVkAfPYUhVJ4hOuk
MWOUmUCTeO9QWCCfdC86h0UH2NxP/4zySDTzCXx6jiuy17u6vO61G1mDPfDkoObG
TVwrTTUHUywUrab8n3Efii4z/w4Bw1psw1GamaG8r7jBDBvzeDch90LraMeahEGd
wqBYwTu5HDbt6Cmqpv25pHx0RBWSXF+FhB0A4P7OrG63jA1M7Qtn5f8DAZhizPHX
e4CFJfSEozBXPVEXJaokMyn0gcUBCeIKCrRiqpEJ6Z7ik76aiZvLjUl0QZr+yv29
O3Ir1CwW82yHwk2fY3EVrEgfPXlJJlHBgXJ3c7RpgZJ917hB7oaqSlF65aEaoVCQ
QYAU+KrDWcFZBGdAjcaUkL6yCi8MBsCdOnM1xryWwbLz6+rcuPPPwtxQF11JhxLL
KbYxp7VzAROvP9xTwW6HUUIhZH8atB5VcS0ogcoh0OpzVHWQJB5+U7AoxOs/R1mT
FnFHLCZwiWiCzX7qMFchOTZz3mZjE7BCUPWK+BPiBkqtEL0W80Pfm5IC9VS7Lqx8
zzc9AZqD0/QbN+m4CAjW8Kc5WenrADx+DHZiu+sluUYlreQIt2Spdng3L6kH5Hbn
gClMKqhBabum8XfEVF0KaAMGeGw5tT5Hwm4Tv8IW1XRJfGkW90TrAOrnHXNA9HyT
P7oOV7ucnO2IeDvx+FGdqXvwzIYCBLYzjZOahGTXjhwRD1sSLHEwyL9Pln9NrOWq
yWzikbSsY8qN7Sl+ctp+QQ8RIw2P/mH8cTk06x8NvD0lE8mShZh71QVPmTOk7GHC
jcQmkvL6JNdJ8lXgcjwT6szs8g/GK+p6UH8LlaBZpaXNI8S7HEprbrcasExAmXAz
h0h8ZDLDTb180chLPu+8plBd4UYKlZGIG/JG6fGNPpKuBbUHzVjjNABWFGeWpj1q
kpqdWBZ5VSyCWLmmzzBM8pP81Tme6obxyH7eUmvrbcsd0nveH3gq2+40XoitbsIn
TWcWg5PPa4ODxwuqabmHrCcrp8iAZl4J09fJqjug+OJcQSnc9cgIJwRJa6qBfn0e
OYimglkph7jxagzid/Sp7Nx1hBjjbKil88ftRixGqbpx8j+H1FVKN+nQz909t8GP
b9tR0OVwi1xSzZwGSK9Q8e/ZDe5SKbhz/czmiCgrsT5yPhVuZgmcu7Nae/oMp50R
PNHr+Uwg5Fg9GFDrPBNaMzSPcFUOUmDrBESL5mn4kJXY9Zd61ACYGR3tQOzUtd2n
oKbGdU/WgHLsbwug6gUDo0vb8KQfA16W00CB+WmwgsMRwU+pQ2/9ZVsS5+CLtsNS
rllsnEvNBGGUIAR1ItTA8hdlyyhQjOmDdhzCJ7zWaKBgcCktpqqIZx8ER6jS2dBY
pTsxsqN/z5Vzxadg1khi4CBL4IuCqwDLrENMYlYr0eY/SI0hfHhIRut1cdg99f4p
MgdbheQvOjQ95UxPcLjJAFlZb5uj8SSj+zCoeN6M9+YnO0WLm0hJfAIDgMzhO97I
aAFSf2herj5rcrPI3B9w0NPVPwnf+y9bocKNBwbimXhapzYsLYTma8MSr7xWjStC
cdyNjImpgYb3pUulWGyhBWmN385rm0wtxAHxWAYXoYWNqt1zz17+zG0bpPCgAFy9
c+1ACqhJRAeUBb1uvf3uYm2mJv4hs4E+JNVmosLcvxqAl6KnYDLLEPhR2BySmr5f
oPBPXncbwqQ+jt5RM+g4VIoNKcbG8+fidUekYCvFni6HGrxTHHqqAZMObfdl8b/p
HlZEGI02a+TV1TIVQQwT4z2dEo0EPf/Vy2z9BQhRZx4ZwCrix5ny5VbBrxQ/kfcC
gnsnYExLL0G1xuyztOnWpipgoEOVKdhsIirxVv4JGHYfwqglCCfc/KnNs17Gx2In
m56cZNPoiUP0wb/Kv//RIfcMywrOuHJUwam9Ao6sGda2Nf9hraPz9sLLI7uCeKYT
DChi8AXhSzSFkMQJkEXGcxb0ypjRt3/uitypvbs5Y7t49ZAZKO3If1epU8MdPdc+
Ri4lVEesCqDTgtoY76e+zgJYUmF2+9e3YTZN+Mm1kLtEXve7CSqt0s9E9lVN2Fhx
Lhjs7YE+NXx893gPcp6xYfCluQFJvTMyYaW2lD9jEsze01wjW8YQcjf21V5L6MRm
iZdDJ/r4dGp7pggFsUcSqnxbVOE+yPkZEHOIudOtl84xgEhpbR6wUxFT/9jZGYAG
+yD1uHOvB6LMtJCrOENVpBl3oFG398fEQrYEe14hzpEmqoB3hxHEfh+JT/wSPw4B
EMpEt+Gep+KCDxLMBtGm05b5bZtF8KDnspJOLd6ewqVlqAIPkjULM4X1UTjmKag7
GWpSpnUML0uHCLb4Q3Tqg3TJiWzHephnDL+8WXm7/DIXikBK1vA2nmMJpDTPZLfg
MBGLm5yJtRhRPJ508JkW1e0ZuejmF9dYCIVG/qzQrYdzm1bD+u3J0gAg+yvTQS5m
BRaybxi39ZHwoFXrVMx5De7sW6aEnHmyzge9A2z7qUpfnoed6SY2SEzssL6rfMs3
2F7OoFuyPrki80gJGSV4Q3vcRZfkVdYAqNylpnPz7gNylNcesRxvoedTovcKB9CP
47bS5N7RtHo1mR6KB6My6XBl4f0Y2ngHMCRy4+KudKiGslvFMTrA5YTCEKCqfssT
dxK4iK3uvC95XVS975LotghFCIYdk5Kss53jxMSxxqQ+IS6JQdqgju4rLubyNNHf
s/HU17WP3HsD8jnu8GUWY0yZ3+Si7B2h1HBEKF9e+1MGjEcafjLJ7fXmwEEF8+sD
IPQ0PiPY5IANn9APgp1g86oIzmi+gW3MVMklK9WvmRp/sBRib4WCuF8b9oP11RI4
n68TZYP0Cm7LEyXarKpfOtrmeRUGDopXq9EaFzxNZBQFOsMxXHNLxqC4v4biEzAa
AkQXtmCS0EbEug3O2HkV6VkvH+Xs80i9m+8OEOEFOHwnf88DdSl7ZncSnhRe/TCL
p0u83pb5PmQssw2bl+o81x9A55fYtx8yiWvTmbm9B1NepHhklKWM71S4gRNleP7J
10YcGZZmATZ+iq5epfLHDezoVVPrpDBEz6ahZ1eDCDawuEA4W+lI2f5woarZ657o
eGJApzjJhFM1oGJ3J/4IXpOuSmS67q0kiTR/VwlXz5Z/M8gB51LBnraqapyZgD83
ZxpJIMcKY8cuywpMsEuP0/NwCPdOQzs1ykB4ZQp0I5pfDZqUsb2qfU1ZOb/wmhO8
1ElfY6kw5GYUrMqeQQwy889OK1cTUoFoD29Q55UsST8qjAln5Etii3EF7t6AlWTu
13qSjQCrlXdi8oPqDbLcSD+/Zf9OR82t25qdp4UUOlphs3Ns8oI3JOGmXg6o+LdP
+4z2r6qHcLcChEyn9LwoJTvqGgceJr3Js1NoR+wc2sXvXZwsG/Th9kCV+jgcHm3d
U1Fsq7aekjmABDtF+EHWA0B7gMKBktqfS9TKE498mhSoHngW3/d8QOuea3Yuj7bf
b1g7vg/GcSy2PptNBeodSK+jJP1vvetzpddDt6qLNxccYrNtZsIHIlfHVPCo0OX9
KmgHrFIzPaBfwKaSeAHLkb+lmA1ykA5M7xgccWiZNfEhZ25jJq1o6YTpt5YTz6Pw
LdRKkbGHfRD7+CwMuer/LmZXtvkGtBXSI4O3J1FDbXtM80cco3BwZPZauBk/Veu2
+D3haEJj0YW9whX8AeJ+GqbttPTYvq81x86WPLEyRNarQuq5/euMNEZhf9TzCABq
ApAftaqyCwOdWjDQNENCCWBJN7I23dlzWi38YNpkPeleHMS+QuHQaL5WP+wplChA
XXo/cQ0Bm4lzCT8m4b5ZpoUlaHOLsXVkR68Q3J6JfsdOzkSG1SaVuyFcSjko4afM
ZJepBktiPpKn6X8PBRDNl1+zCyIUZ9qyvp0R6YwIYFv3hwnwZxr/BfHk/Pr5TQLY
4KeNx0aBrwBlG1USBShrgYvUxkqms2cA+tVSqQ7huniyQiTM33226JMo4YSR3dw0
resdOUJ/Fn/uNt8LpJ9cqyoP/87jxSqJIU59ZaBFqSUQfooiYDMmcLb7IqFekctG
1sa7CeDZznPKwbnHcWmmTHq49FPA2Py1daqADVqnesx6n3qNstbqosqE2+iqFDwD
xqYM9xqdY+znmquN8Gy9TkOa5W0MX0zfMnrvZky2guoCaTN974u0xkdRCppzL55p
OWkwlVcHEevsvVCjhJwzJvHe1QBWLkUC3Yqt4d6QFx5RNaUK+b0vDqy3xB2aynVD
bJ7PWss8z+zNsiX+u7zt64pAuUmtUgwZTVxs9u0SIbis+cuiTJ17rAWkUljMENuA
u2N76QoJcC9u+crRQW5HJpXsx/P5JHyoE3V1XWNBYwke2hBd5j4bOtm7/GAqcOsQ
NxOwQ9c1K4XRZ0iGkiLcc8syq/Hik5X5byMrGPUPDOfQJLH0bh/3e/IDKIel9cjP
axae89iq4U97vqay3W2qzKKVksl/hl6JzgVWUVT2yMuTRqCw0y5YbJh6wSTrIqgL
aRbKSVcqmqQP/6uQhUVExwjJ5YALYXYAhCFDzZwaxsJBqWqzUF+SpJkNLmS950l8
orCX6WObl3Xhvp6cG/vzxBGjdQ49naY7BZNXtfLOFdcOVo+gsWG3dHYfyCZMt2Mb
cAPLTkyYq4QGoUz+86EQxwaXoQsOJBJay4vVzZrqm3H9G9DR7bWpkOmAcAznbOaP
RjBOxFsuEt9MaE9Iz4Dk6cwtI7mMDUUm3/2PM8Y5HnJKIADR2S/74QPKHMW2PeUN
SeAfmTiqvdY1MeNyb8W7Vp5IGn+ozI37cj0v+AtfUcmi8Blo/EX5doWpw6uv1b2X
mJ1icULIcOoErZlKHZX9mRSNoyChvYR00ZdxgjSrfmIUkTs8J0lEJVsvicW2CQMy
KzUXX+qFiabsOZ2pvL6Uj/0ZHTjBuXRh2Ep1CiU3eYaBTzhveNZ8gn20V6kaVo8U
SiQDcO8VXlXk9lnbw1PYUbDOEEa4lSH4M+rlDsdF8pWKkHXXos6RSy5dQ34BO6I4
GbkZaCExWO2rkU64ESMeZ8BvY2Ia2HlLVn1Vf91ikWSM3/MAboGnUihb0cFGsmov
80pjw5WDnA4ORQfM5rXKu4rOyNVxsPCprxxMtN63gKKng3MjvkHdiyoDI+5ax/qW
y//bQdeuMIzF7Ymum9ILC8C/3P4Iy+pbjR4Xv5GBeFnK02t9hNE3lbhiFFPn2h2R
eaThuDdLBzmeK45YkH5QWnzQlWvglAaKpbJu4BCmCjr5wtI/aPSokijNwBQNcWVR
SqHUYXGOyRGbTKowWQm1kgjGq5Ytl6N9NGdnFcaa3dCfg895861pw4imXAMvtwCy
C5BU/svddMU5LtGeTP1o/LSvBNDL1h/qzJ9Xe96BbQraYR++caSDCftE6s2Yu1N4
11+q5Imi5XOU8EZzgYx/2Sv4uh/4ojfSHm8flN91hQTG/RCF0/L8wpI+gm8jOzYY
GiU651M4eNddq4llZuCrrSwead68bdzIb7Kn7tiemlVUKzuFOcOgxNBOQ/n0LZEq
euyk3XP+dDbDTiScGjXHwMhy8a5mpdq0fzhLO2NRq2CtKu2DJQih1le87fi4E6WK
LZmt0TLJ/t3HKNiPtXj4EEBVjh0cSLD25ge/EaDBSf84N0g3cKwTa8WVZBYLklvY
36y6Fyj0atZHVKp7xf/4MsvrVk3XHYuuJNatuxgsDOq7YT/CcgV5v5oKzi1ksC97
uJ+BsoCHXtv6KZlN9url8HUpeqVdKkzXDuXZFRChK/KGSE6CaXJw0p7Le32/uuli
pLkNGQpXq4hxMXq4jdsoYuSHsltN9cfi+OGivMjH4M75EAMDMerBi53mvpHtUuyd
wqaWeBPtDFnIBkYYXe560pG32EkwAUV7KNNFZGE3rROd0b7QBzKCOlFgQ14xxuYS
/25UwUHIk/NFsEKaww/VFLF+NpQxkwJUhldTUuVGwZOFrgu5n2FOT/OlG3PHwJGe
7xyqNQ6BQmOcogtK+vQxzPGiPzJziWIzPn+DswXckAK8SCGcfYlCIU66LTLsl4eI
TWLeVRK3eFtKOHB4xS+VqfokwLOe9c6n1451jukEID8N356p56/SLwD+CT3H5DTI
2Q24V0a6hjkXZHkE0Skx6hZqlJo48KFASX2BhxuLvNpoXJJOtfUUX3nBBGMpGPON
5e5fmEKqzRE2vsXdAraMLmTQ4+2DbjBCmQynw5hM/4Vwp07BKwxXk8Maezc2QO/i
/peFtsazCGX6aQHm+g6IxuxhNkGSNNQ43gpcKKC4gMBQWpR660cDjYEsNlSVzg8n
u+ixE3CqnVpMpmNizmnYa5EV+d0mEzCDi/u/UqQ6H2WhpM4sERMXmq8JMWo+JmN9
tHvbcFV88Bz+LgMwTunaNZGDjyM2CjDQQMTY7WOg5hfUIRHASv/H+OFheb0pPgUS
NrctMhrOtQDH9CGEQ4AqhBs8elB1UFaLGsDsR47ULTC2QSE3VvS9LvAsocpqD6nB
jsQFv0DcPbGhs2nNo8h4zNI5/miakt6tzETxb9dQJiQ/wUkzoHWCPiZWBnBgrmML
+5/zeSnOe+AxibKmnWLIR402wPLCWaImbv/tReoCG511HJ2KzPFwAaxHF3Zc2cXd
hF9Fzylw2It4BeyJPfcp0xZ101j+4h0Z6cEkWekZ438emzyX4ojMS/k6xPnH8Xgr
6efr2k3EYntuj9uwf2bDkFq3eeWWLDzPT34jIoSgrMdzQWR9OyGe/8MBWO8ODVpN
KXK2SQjVqQd8WpbBewv75GvIREoKD3JnFVR+yd2nOi43hXoPcGTfRJIwK3ELJwPp
PZXRHC1yZOYJwY1AHShL9zA3wLNwaNP8W5/Wb6nXxRJgRz+869Zfcfpyq9P4GmX7
ohP06ropfmZAg6dpu9cjyf5fqJXSvuqB2BEaGNTh15p9XnctbLAziDiQ0CwXfY90
npglivWT52f719QKUQLTtJjOznoU20juFDmJ2sLk56MVOnfBOVua95atu+4tHU2+
xEd+vM64w910BfX3CnXnwVHWiE2lSJhBraVQOvFUxRvN81VrhdSApIJHhW+WGI5V
fIcAJTdvlbjBxdEniNpn8RuxSBk4a+L2XXD0gby+cQGJ7kOv7PNlFEFXfF76oN3P
JdIi4SK8ayNOncHOYt1AgGCl3ZwaTrkiOMFvbWLrRUEj0cviN8A7IU6rha1Eg3ej
b8PkdYv5pS8fkoT1uOFLkjPr6jZ9W4D9ssmX1LCz7SpjxfPgPyPwhoTzf1E6/Nlj
P2VZG9D1E9OONmZg2TaGtc+FzCkDpxCjVGvrwngDokSrJE2SzKb5nySbqNK5TXTG
uiqbvHU9AEHUHgmB68aQiR6RoHWyirsL3lAXfDAtKAzd+7fnA0R8fCo5YDm4yWaG
B9bOjB4WIYOYZLZuIEX/kkrH5uFD2vtOs/455OWomfNZlUJSM3N6cXiHB7NpPbs8
jgtr1pOVKEdeLh/iEBzK4AWWAr/h0/SzQj6gkCMhTxNIsUb07aoIpxwrIqwUOACP
+rtIQRfwrq2wDvyY94iwbb4xLKJuC/O51GQlXQwMV9ub+agGxl6YecpuOyzx/K9c
3Snwa/P0nYPwoq4AfB9U7qEJvGLCOpNymbCO//NhWoeRxQr0O7vpAz9qKdJCANpi
pRgsJKzY6zFIleQzGQlayj/AlVB5+TJSGajvf59egFLB+SOWB3xq9+NNFnxGpBWZ
WBwGevBTzP6QSw3p4A4Y3q+Mpqct/+0WVpgAuckx5UcDBR4Y+s95oDxi5s26B3zx
OgU0ScD0GA2oF3fXQfpNk8e7OtEP1D3RMwSJkYzHoECaqeR4TN0iXq4//W73LQEH
0tBM6KOQH4RnEQuYW2cW7pBMH5yvypWWhU3aQjxjoLX8JNcZc913eep8R/Npzc6z
lx1UUjPRXA1+B/b/yfkmAcBd9a1xEP/LmlTQxaQL7WXHsm1vSZXA7nrO9Kx1WATr
jcz+dM/dOrMqSspRotaL5ntlbaS5iDqWHLWu0J7RvxKSMrDNsw1P/sPtm1BOCXjN
vnfYy5U2KygBBIc0WeBTrraUIKCqB5/Plr6s329FfUQYWTJ2vpIhtxNsujaRSaDW
O04M8R9+9uzI9qhBkDdYkHqIsbbA6TGgAAkhfah5EChXnScpEq3xhdid7lzPo4K/
TqFF5E0lAyh34Yj2nMDro2JLdrux/q4HfMMrMgmEt+LagI9fBoNxa4EYvu47LZss
hqVRjd03OSVcUtzwjSQJSlu23sACAL28t93L/UGqXu8Ka47KV/OMuHIi398ziMPZ
+Wvo3olwXgqgtwgHo+hDJ+xMNXUe09kjN3SXvQGuKuTzjteSPI4/D5YC9s/TjYCt
tmttcvUrMXunsHMiuR79hZhTb/Oat9xorkv7YI0s1OWviMN+uonjfew7TsOrk+Y7
wEKPWmj7L+JJBA0UuODwccEPGRDBYPxCBBVJXbNkDesr8C06Tn60ouim1QsBt6ud
MsgPRPvEj3k4c71F4u1oolqfBxaU8tuEFwwEjvs269sUXmwTNK/QZ5tgugwsJ0MK
/o+A5w16O+aQ9fAoCdMo+PFE4K2ymplaMclVEhkDAlGvmpmWoyZqqPECgBSooFNM
siAAQnnx1YNsiMyLvn0lxh8tl+Mjoo4ANrBI8cSoudnKUWDZzRW5ubvXG35jyqfL
VtBogQxEdTFqozOupj2iyI5jAyRK0uV67ioYEjkU4FRx0tjbW5HSbLiriN6bAlrq
kZZevG6RMCWIt26C3mLBRlAcxpMEIfJt4G+bMzkMI04NupPNMac0w00X0xR5gvfw
+YbB/mgR0Zwvw+dS6TkSsdKcKKRAOWRRwFw0RrKdjtxhEJdbV8j3D2YvbDVsy5ZP
Dd99ubxQ1ZPZIUyDJA0NBDBMeVOuRL4o0K2VoS00NOuf1wVBtCNacywpQpuDSy9F
1UDwepvRzEyQZtsozCFL8srakjP3NBLVcP+suUnb86Nj/tWTE5DopmmpLcSq4Ue6
JfjLiB8GkbocLOhOGBuZwKJCH3CTwnvAcPvPEXUfBChZfpiF5iBMpUwka00IgX/a
2KAL43/nLwT9BYVI1UfglJJvuD6rXiPGmJt+osGrKb9YYdBTw+T0D+Jd6+B80tAY
nJyIwKV8GdkNbCa65RZ4qhLMEq422behYxI5j1dJiVOjKavKGyEllpYjD+5TZxwz
IbM1+z254E+CBkgMssQ1Qf9DsoZ8bJUG2oBewrXLNpaKmSjqHbD4/ea2j93Ic2lX
plC8lNEBzN7/WTOyYhNk3g3e2DyJbUyq31DIY8zdGLLEQ9gmF30303C5FGfmj9bG
UcBl+IU+h8bW+E7TyRDCLaR15Q0qnrbUwt1l7c/aJdPyaHHdlcPlww8I5LWRMyci
cU/YhDdedrSJSCWxCesp99GE1Gn233Wm4EnIQUTXc3oyH6cosGS/9qYis5KUaCUe
l5DmWCEhwY/ugnmI/6YQzNCoUShQkiMO6uj6AqFt6XESPeHmVfOyKI31JO0CJlEM
x62u73LV4bhJHDBEByR3FkUI70wcc6Vf4rD+Gc1XIkX46bXtLb3LsWsPZVAwOO9y
ppnxFwSSptZCteE0ls07yWYNCmurzDk9ArrvrceISZPy7Gm8IGARge1cYTL04iFJ
NaLko+lahoRC0/aUpmPsBhLcLnZbtlzV59X676JA+j4inKdiwb8fD7d7KjyQnyiu
aa0vV8LnqntyMB9gNfKYwavHbH5L+LeNvY8GLjAGLxrNsZhxVxoCWLznCXsEyxZK
nT0hArMdQ29wkkG2rxZVlnNAfHq/8c3+Fy2aS+BmjmiufAzaxBGVhwhlOaVJFfSr
2AVzPjgpvmmFaD2AHMNbENG/Ry7k6Du5Bho+6B4w5Px6vE0eHZ3wXAn3VL2E/UjM
y67ymqM1EqBXZ/lpm0OQ7mO2kL53qw3Fcaa3ATaAsWaNHWq6IwXUcjQ3sl1bjZ0M
VeB4DNlhGyPv56+R+zM5cnREQBWVcoHF7vegFVgScAIh6mH8YXwFPvxrJ4Ue4s2O
M4QIiX03HPh2XNcwlKNOMyj6T11kS23XeZrZw/7Y/Qrlda9/w5pf+lMgVnmG5lTg
0rzNHI5bzHbA4ldMwkwYVvZ8waKXmegUOD0F2iE1OKTJJJ525LHAOUQ3iK37dziK
ViTnpyvM/MQOIeTFIDlnMXUPrIGD2VGg23Iwh35HbJBb2TykU8erZkgxER8toQr0
89IRNsriTl/tufdPUHaIN2BtGCtt/YFf1mdK1pKiBBeO/HC2Yc1ZRU4yYmvaULLd
9KE5d+7cwtJhqte5tP2RIR5bYTjn9OvR/sFD2eArjDW2mCjP9YjYyykhxfB9sjiZ
Q4QLqDz8/xx46yWRDgXF3PlxKM2FU2CULzGTo9KxB9a5wqQp2ybSmETXBocUx+QZ
2wQ6RINpTIkNMJqe16E84qm7PAvApX9x1L5r9oP/CsJDpDgYk1RhJBaDfuKzc65L
Dbsg1Y0fOX305eFzUVVLG/UlYftxom3WAM8wwnBfvRWk86Uj3SjWvmbx4tph1O/i
koc7g/TrdFIR5rqU0EcLVm/dLjqtzOdmry02q0YUM2d6niSF9zHP7HSXAAT450IJ
o3hamGGE8aEvfLdNqRDRK97dTf4oQIpCSCa1RHQ42g7mtC7wfYuiwQ9pRAd/X+5N
agOblgBLAGph64wujukkMUMLq5i8X0hx3kSHNfAH6zX6BwR2TAdDxaN2gW3ZJMTV
R2+Wq+VZ8Ke+yxmkNghMRQ4bq8VGe0/vvrI3VfkP1iE8wZ9WzwtytOWHNe7Glpdw
19mIro4BAWwYvMKNfC2PY89tA0/SHh4QXl7HNdaMMII0r7SmTpHE0PnEWvYSjQs6
jg5okheArkN7jvkRr7ZM9/kp0CsglGz/JSEPqwbAlwF9BDl1aqhJxFjOre6vx3Sr
R9h3mObY1uJZ4VuGCSB3Y85Lds1geP9VAu/N97TdjsBl8T3XEuWVnyrYtCUQ7WKO
U1CPngoBC6cqzDOiQM2RqXOLelTl4MnxxyyGhOPn2rlXA7K/tcX7BN6VZTJbfyzl
PDt23s2IbdDLuPhaxBYdA3IUh1XIykaTfL5Jm6yHFRDP9zY7XldrmSHdUUKjPrdS
ABjP5rF8g0iSsfvPXejMtGsLdMqymhFhiTywnVa3T0dmw3Do8oVcDI31ij1A6rl4
S3+M56lSZMhFQADLO5b0CzX7uWclWxrTVpF+sZnsY1SiHX1IcdD+niLTunbWTuMF
0svIhiD67AYUjvjm0jmjiJM5raxiiq2BS8UQI+CufNS3ipM1MR+quy9eEDM0FbIS
NMBlJaiWikZTv79WGM8VpVlo5f20WzN2R4J+wqq4uCgil+eKzciaLbVsBgeFhLzX
Hyzse92lNGfaZE2I3hKp4cF+OCumbITXxprONc1dtUHt2qENZlZQlgvlaKgjPnM6
FVLowc4F6TsjL1p4pAIh6ExRhrocUhoTbBD0Z1xKq+7YZZh2SC0voHIL4bw+VrKH
fVCSqwwYsQVWQgzsVU+Q+pTprSxYSHI6mcCZMJE2Xd1Terci1FZKJ/c3NcviaojU
9Wn6ghAki+RLGZLqJ2fs8htpHKJtuq29V+pGlIiDVSvLh6MGb+VqkLRyb7u1pI02
Wo/YXke1dsA9F8gWePcsT1b0hZuXkWrt9xtUzpQY6Lpj+966WG10PQE7XDKrg5pd
Kcg4XicKpVlbT0u9c0GxP1trAjuPVcpmpS030WOFAAbSgKBqxnFT73U8/xyIg1Wl
wo+fvLLqN8c/HK3V6ou93zDlpACVXKd+OpLYFKzgqGS1zBVG0ljtrd79ziZfJEg0
ksvA9RN+VAVktjlTTRz5l9SzSkrpIqscdNJr1dEsLFg6BOixTEpHoFJ3TDHbl5cX
REREYgiWLQ+fXBDmFbBRSLeF6vWz2ERrXWYul++u43mlbh3AgTem9/wK2c9KAd5K
mPqoiYB1KA7GMk6nOs+6v/SWDWyjcWA8ZerxH3I+YA1I7+5dw/PRvAHthgrbGYvr
bapzfx41YKqPbammLzGsvP0BOECWEjQH9sWU+2/Qml94zRhGU/NicvGD1yhjgcyp
oAHotKSlc7Jqzu9DQcVpX8OTam7eS+BwJV9mvfkT7V/aUuZ5oq8c6iG/WhDjS9FK
tMM/9FCVshlC/VXRh+rrgDnG+2lZuvMpTAOMICxqydiXFyz97CZPNipq5gBj+35I
W84s+VRycDzurRE2Rh9oZ+jY54plekEx+Dui15xcduYmYlZs/lHCnHKAZoTXVDnG
W+8Vrcghqx6JLm1aGJJQFEVhWP5B+D2eeUWMdCeT5y8UdFrDTCRGYB83LvSbmW0+
/k9a+pAkpIk/4QFuzjO1LHp2jSOl03fODL/SPmP3zBCC1pFjZlW8M2zldg+cIzZm
u8P3xx2SOEXQ3BtCj0abNbv0yZ7ITVGQvmao8aLC7F4iwvZjuh5RkYNGahv1AY/J
zz2uDGd0xi6sO54URZOhn90yDSw+v809dhf7lTTjS5LEHNxEWQPy7H7hQQsIe26n
24Wgry/fdN40P1eXLGqeRcLN07am+dlRmk4o/cgMxH350FJbNoPX6MvOSpx5ZBuv
xGrk5x07EoB6d5ilgRnvL8Q5XlrqHo+pjtr88vrG7pewWzDhttQKm3zoUuoB9hNI
IUGMLvK2ybbUrJuXpmfHzH1KWgALV6LuTkfEq/ZmzhlEZRPXAXpyJslxh4KytzGY
czgOAGyVQM1tG0K2+pbB26ooimFDLwwlGyOh654w+fWEx1HcJQJsGrSddwmqcRhF
0XmPw459wR/n/+UQurPCK4UnN99x2AHiS66ZzD3yfdZ0LJ5ADquf4IZXDy3YnEKK
PkUuUwPQpPIRnCay7dwmz4N9te8VPM71O2c8Q9ZIHeScU797a21t/8l+ZRE0cdxQ
qlI7p069fMS3NvlNJE3Q2jNqNt1BnaUW06lDWXt/Kq848VYmJxTlu/2mwZA0X9yf
StBiIf/P9Upmhni6R8IKppj2pkZgfNPiRChzcqUFQbU2EDGneE5hFbCPL3vbxsd7
GaC21ILJ8yqU/lmbslfN/jXz/Vf/6/gHkurTNze1whZduZ7XBYZe5LCQfS4m9tVK
hq1GX9/aIcLtNIW1LkzIxHl++Ll4FF4yg+JmqBXNQ1l9wl8jQGx4kLlorbidxiYh
ynmeSPL9xhGN8Mluc0GR/Boi6fDgdps5zTbvTvMq0gaNho+qLs5T+Qg139cbpJwb
5L1jwGibVDcbUVZs73997R/acHGZg6R5vufVjZaAC6ZC4tyWqJjLea95ypWwp1mN
jeqD/eH0TYbdUjLTFrW1JyprMel/DcoUfZsUMOekwFC6+8aayt9Vj+x1+xRUmwQV
puntiBgZyOhzSnxbjLmgIE6iyl4bOHp9iqsYW8kNCub48Vn+rY6hA6gYk0gzkTK3
xlCZMingZ45R5PGuJLRY8WwUk1OCuaIxKr15V6HX2gYCoC+jqukFIxCY5/zkg6/w
Kxqf9S7Fpb31iIl7TdjVPdUrKoJzAIl4fOIz1vd7PLymwEOzbKbixFzuUzOyzVaD
YbS+076aiIfV+6XcBjFRjB9oc7i8cLgTj3XqpDwTqzAcMJs1nFHA/iQjBXvlceqx
yYhODMwmtwo/w0eYh5TJCo6U13o26WFKI/jqmj1F1g8boAFzRXDoxrWw6E0oRtME
AgzoLjPH2CH8PWMOg/cowCrjf2MHqNNHLN4yLDGn3nq8DdlncSktexZOf9ZMbCJm
s25ggN/S3wa9krWz5+sRQVnLOw0rq2Ajorx5ZCU8RsJMKjPOzjG9X/APBlCPz07a
OE0GnBpSHNQZDUtqQ8pyD4adJH5VgeB02dsH6PpP/u3R8m1S7Z5GvbWLarJBml24
mi6ECi+LJ3rC+OeI9uVkLYBdhtqWl14e40zFYUZCr+iGfz/hI2WWlGUAth66hZLM
bn5xMW2i+7opI72tfddsaBrZfSR5QD15kDbfcS+1SUrCBjG/7Sr9KnzUZUZaZ3p5
Gv75uVbugLM2k09IrSK8vAx8WvIOMDjO9wJUszLXo7+lKtXlOXai2aMb0GcDX4Y0
doNpzx283fwbHpV3Z2JarwuPUZKoCYIcuNa0FIE+K3m0HYQnuDIxF7eE+6UjNMqH
09KSUMe/WiEzaXhiZAJd0v9el7dAGPACBubkJvq5vhuF+MOUkfynVX77u5wgKkXX
n5QbvvaGvPto22Vxv6BFtkyWgxn09Dx8z9YOPAUxFChGwCB6lH0ICmBtak08Bq8J
a4YNwgHGi5zvC7thh8xmPP9ZkYQ0/CUQmBSbsV2CDB/C3X6JekwchZzNrN5zpoz/
soax/qnulmu3DLQLVZHQkcQrufv5+nc+J+eotr3xojuoVLNaDZd1LWoPc/sRpGHd
Jgx3SR2Fo9aQhNi3/L38S8v+0DqwalN3hwLnAcu1gBxCFP1mkubxTaUOM6idOqPN
ucy3Bw+1VAo1peUGrIIgRAmp6JIbSFohDFgyLdgvQbmOcA/NkSJRYuYgwvSUPdnd
NSyoPd70RuI2DebuaUcutmHFqOtks3JrIfeTnRjreY3Re3GDBSMQJz8cKGNUamo6
527gu1sUqcmATcgnRh8J22lJgKYIYKU42s4HqI+N8Q1BljoeGHm/HKRaPfJdPA6q
wax0njvy5FvAhBKlVvkGYdAzjT+9VclbVAJKvottueu82N5+7G3C/72WHG5YrRIN
a9aW2vw6YIV9ZSrJDASAPHF5BtW861K1l5YHSHlFoCK5VXeZqFX5XHBxC0/rbyyW
5zJD9NexZ1U4BdptVtfK9Wtih18d+lio3oTHnsHavEaW3WE+YE7RhwpJPZN3IU+o
q0+yCtQ5C0XdW0Nl/0/W7UUVJvwl9lmRHOC7MaF+D8FK4Ma/vfEyq42HgjV8Fx48
PYWWvRQvra5/umCDBDZL3Ix+WCVnjcNwVeZUh9zIDhCt/PgFHhTyUh80FxQs3RLd
75IUK/IPUsGVr9HLReYcdWVRa4RSjcGgL+SSDj2hCMTM1/rl8IcaMg6Eebi6H1zw
ktPb/kH+XTCTe07rkM/SyPrqqsjT5tO5/vUY9vtAw5+LP03VAXaESnJLrPpHgMjB
Ele/gE/0wgwSCW9PMMKjngcJLKH+TrUgNA0sp1LxuwY1x7TmOEjQ9luPcTa8ondJ
JeNfoa6e2M6TutJGo8tAqA+//PutU4ULVHg3XBuE4oaWDUolVHyo0XxVJi3mfUG3
d8frRgi9ULlmuCumgmnLbJrIOfddwUD60FiFWX+m+mKiVeTuO0RVxLRHXaLu2oiL
QyDfF5hwHWqCdEbbPb9Qm1q1fekVha7zBz4IA4vqrLRES+43svklClMiCP0imo57
RQvuOElHsDGNkJLNAppZZu5L26MvoH6AQtD23AMCVHUyrLiykiq/lSd+MeXdPexQ
Dy/aagUI2/DslPkFnqBbClQNlBhCoMYvJggAP8QWF2CCrR1/NpeP2Bh/zHVVFR8W
kZTBcFcERjlt2dbwQGNi30B76NWW3Ta3x2bQ1nb3Po7DDbdMhhwMyyKiWtr0DxVK
AKBU3eNvxSNEhFbom4q4lY4eU2/EbYWQsdJUnm9isbNmVoi6dH9vCZN1FyBHOoTU
CjzAmGODS/XDEYE4xh4wXdchJ14+aHMUtKELcK9fWx4mDA4jJ0nM9fNsIlZBKcvi
BQVyHo6LhkKLodxM97D7jgJmtlK4THaSTDr/dmh7gvJe8h0o64Gy0OH/0vCCIc79
ADesVrnG6FRvPxApOPav7k/38D2ZHcA2+qFqWC9IHON4moyE9uZsgWUhEroDiqmV
ODzHig6FRokGb58sGH6HAp3/B0NwaeIc6ZQ8gPGKCj7r2zXa15ymHAmFh3wCRePk
ZwC9Z+EgzN4y3SClrLS7cddcJsG+YBx3FZ6RsqntD//OyzMMg2H+artRjMArzy7+
MPLlurpA8nqbKbIV/R1UPQiPINTNkx51dsRaS4FozNbNK5hbCcts7lzyVjsKYtH2
x7nZrthoc8pO23EcfslvGpF6Ay/uCuZchsgARgAAsO9wZDV36nCNAE0IQZmTRBVX
ueyRIsXRXouL6WHw5u6VTMbUDJQSIPnvRQJQ1eNWxVCLu3rYaiaIKipDPJ3xQgc0
nrtHl/Nv734y55tiwb8+ABcNaggND6HXVm6wOSKzo0RPMyDqqqmlneotoKp7bat1
HFvlbzJxebSzIZGX6Rsvs/fh5GRMkS1vJLt98l7s6In7VHoHdwttsTQCShUkTU/2
c+FcsDFLWb1RZ0O6kTOXBIV8gx2vVdax/gTT/52psbvkQaLUjKtyGJA+CkUXm4rr
maxAfRI7WUcs64vYivhLgHSMayXKbS8bsd89nRiZE/3OBHwJgY8sw6N3d+TbhjuB
Sdzb0DrFkv8/9g7Px6BHJAdWvNuI+9n3zi912JgwxoHuZWMOJrxzE/+ILOFX/X5h
/0UsCWPnIIZzpjalVv4cMxyvguwmIt4SLt32bxccjzuvsiaUM/sNc/H5cAjchKwL
D3ww0Lt9swPCRJcET1/jP+LefgPYL2cbD2ei9oj+ps14VJFEyTzFdVszHxCu6Vjc
YXVUBFpLddrSunpTZcUqg6WVilWkAqzomwr4623hvMJZpVM07zR5bbYNHTpnkeL7
PYy1WpD6jKcGJXlPGe/1CY9VdcrttHCj1/sn6SfVCkxKR/sVcSx0DEU9hmhpBAe4
IcyLv1BLQYIR1LfjEvUYVzP26VIvDm2DpnGQ7kUB+a8rIE/IGVrTwiBtV17zb78M
BSMHjyAiQfEfHScBBSue9i5wXOUigMu/6xQOrgzLHPw//n0guJ2NPL6xaPQtWBKO
Q8+pWB8nsjov+UZ93loavRLfN5OSFcyvtiTW4Q0s8bCo1a53PPG4pern1wN6He86
hJKnxTCxwGDgbFOYK9cnMurCN4RALV02MovkyJKa+2UQ9j/SMMqWkfZqXpN9s4Kl
O/BdgbHQ0mdslbTu4ERAgeGoNketfb95xIQQ3WcLgT9AxdIWa1vxMV/FP4xIQQHP
jhQ8G9psbsPmbfwzm3h1qosl6aBDF3KMiu9lIJqCLtdGYExSMyWsxQMTeiLVKz0R
H763me0+1rYIWCa0+pbuF8SY4tGBUawVGI7R1mrA8qFbjxczFInRnmsw4j5ZJX9p
pIkQ3f/Fx0/ZslzzyiHnjqsDfQ/lyUFJ9OzFkvZvmSO2GSsfZWtWSmGHN67P3iiQ
BBxaiTe3ad7SgvdxSot88xj8IsmlpIbX5rMUoY6pnQUTA+WlZUPaD8VkW8A6IrWQ
11uVWCi1yOcB6VgNToPoKmYierBn5VOHr2qXQ0dLKIQLHTwG01nobpw0r1Y1mCHB
MT/BphWD6Kvqol3N2b+JBctqGwCQXX07Ccj9L/sCIN34SVxaqyL7uwE6jktJJ5eD
Wo+usvD67r8aBxlgPPCC+cZLuMsK6BJmZMZxeUGFbMwV/DVJZBMtJKZ8oJlUZ/jS
5ofBTWzuN3WEo19bqDlGlxax7fs+MTPSgLQlzZ1YCXMmU92Xf5ZGpxOrOB+Os7T9
SZC6GDJ8HjmOlsMo7GSGnTfId/gV4AcqFW1HjKAp2OHwOYCAZ1DFoOUVHX5LejH0
TTch5iSaRcphaUf9/K1OIH2+jD4DZDzm+ok+2Rs36BtfsnwoMGQbgJE8Xshdz4Vi
h2Yt65yUTrY+KCy28RrerHLYIPACvJoteRrVx54KcrgZ6K1JTkqqvisjTOBWH8J/
CxO+rUdAeeqH4Om1Uo0Wir8KCiUnX9dforOKdj3sPwju1ZH5tXsFHMPpGptSqJdC
BrMFVKiE6FHIBU9ad6Qu0X8ilFezv5R3EXCdCTJO5CxPN10ZAskeuPZWfo5Zqwer
K3P0VC/m/k5Pt2bSTgQRiFRKmsb19K0bTnJ5b198tugJIL5vb6Bg4lXjKooDqgAk
f0PNmIgLfmGoVHKsVXBVA1MNB5+f85TaY2XJ6njjGw+Sun/mWwhdnKmp8JQr1nIB
m7t+svWDwop4/KYftxV1z3sRplgPs6ZpbaEW11sfvvBxeoczOBUDSfF5Yc6u220v
KsujBCHCDmiIwE2mTq0Bat6vC/VIeVK/gQMntRtZpX/lToZnasser3EOURU3R6wU
E62Uzj5R7dxWlZbA/9WfOh0uBSyxzLanAL2IZMAGtC4HHDA/P03dZipvGD1xNLvR
dxRfkUKiE1tTPM10gSXJZW42JAf0WNFafne0vWmK/PSHP6dB/z1TihMKJdfVv1LG
zolMvVB1JK8tRAXvzfrSKixBfxjD/aLkQzNp70PfQMebUE3qmrR44SP6I0cAtIC0
psZ9NTC7xnoXIxMvcKmw43LepDBu2VbYmoMuBRanXgr8xXsUKlxZseqlUSzbwBTZ
FtCNtBxl1bwf74b4I3cZMelGeNLz7EHWhok1pwY/+P17lt6WdG4TANTx73sGy60y
DWBAirA/keQKhbnr3PKfgun5qQmR8/va5r9mhcwObEQC6VYvTJ4uqIdDhxAlqrmY
aUCoi0zXhICGFX1bJ+mwuGPX5rCZsXl8XM7YRZzMuN1ELCS9TfnIwiGVqMfjyhHF
xrElRHfUNnlCLippbdMA7cSqjFJ9Jei1SNEFsVor/bTjoj8B55P/JRmvKkX0xmuJ
4XE4U3LvyonXTbHkT4kOv3YZ26LNzzSXdXp45U8Ij3Nyi70kO28adfPbKZpz9KAI
/1A/BvzOENYyZ0fHUkfr5ylm3SVrbxr3rkrHsAInBuxObVwTE1qdmFujh9kR8oK+
gxv+F+qtS9qboHHsH7J4RBz54D8BDPMaiSp1jSbakliJ2xOObhux4I/ewfqDSMuU
xvB/NKFcmxbmDy5QAYukNLXMN3nEquv50HsGZ3vjUNPbBlfCxehtQr1a/hm+6+hZ
ldPStC84uXpkWLSPIANKNZ0H/2MtNHkvR9Iye8OMHniJ0lcSFuqPyDen4EreYxXt
0myyxizTsXwhmSnihvkgCnWcgidsz7dgVptbqHiTbkkFvWjgMlMOfPrRjy5ZwmjH
o363bXblVp1s6LxhSmpIQUpIVSUqoEgXzPWb/zu1okH+POcGXNH7kigUUcRRo12e
bKozYvmYYEkcfHz0r2Mtg+GytWeYgtGyp5wKB0Rm8PGnmzzEHFTepO0HP+oj9bi9
771JfKFGFxQldHvpESPZGMaQ6KcepkglG183zzp/7/xy6bir0AS1c1oBKnq8B8qc
cEpLMFYoDvlnE0LKDsQW2myqctKaLEOM9u5wW/KIr6Y7gn4ggt3lSjEHUrazIcJ7
ScjpBaiAks+zposg8bTA/G7Q0HdWLj87iNvEmfjVeV4fmGLC5idHP6vgBEcptusu
6yl4U9N97lrhY8d8hz23Jc7v9qF2ndO9vEYZFCKfwF/6HBaEhxO7V4wW3FK3qb+2
yB2G+IuE5MUkLpxWAj94KfOZJ4Q1QOwNAYgYQlfIYDJ4BD5zZe+AHrVCrmvWgmxg
5XIa8gwY53kCqVNX4lvYupmFBUstYz1u5hlNRDymCJdLksChaI0rA1/WP6DZmgyq
6mtAxGy5vkT8/pb2osWfvq/biBE4RRtASVtVX2mCj2VkWO1ff11khzStIbUWBoGS
Jgp9N+1uJZM8Eya28V0PvjnpciVfGwrJ1fpBD5m1NPwi0+00tEccZ9R1A1EqSCc1
s24soVhvyUIWAhAJ69KMprSvT5lMjsBoXFPB92tQKwghnHQHXrPxccJlUuCvtNav
FX3xCfFhLDSPU33QjxDr/QpjToaT/a3fM0tAQ28KdVORwlHg8hfwzvHheHkMmldN
TxQJjKp5Gl1M/MUe4jEwPGeN44Ss8KZ9Vk5WeIqIGRoFZdAPta592/8UV+A16lI2
eX5lpeoZWHMDdu0DNKggKkOq0ABee+JvYeTxcxi1Xpy6hgg7VXwBl7jhSQPw1ode
Fwb9LdLSmUDG/mL8/8BnwYWuQV94vstU+ZfPwXITad5mFlpYyaBgDU1R/eXDCtby
NZz7QnbEUO6tLrJQFDtpnsnpkrFH56E0RTspWPNYK0AGERC01uprGaQ/q7mJli0t
1pdjy/QyH4zCeXrr3MuT5H+dGirLIlxVKNV/cyShiwy3iQy357IqQEfTcTXSD3I+
Y2cyEml4BaKt93DWTPXapIg/CdVjlaSw7+N/QC6+UDXTpKV2aelQK0jiilgMhOBq
KMthKa/KhYsahnGFV1hQuJSNwF+bYnZ1OHKDDo196qEZLQaNg6R0cJQX6dQEcjdC
Zfm5LCO5oaGLw65KQWptyiPayRWMGEYq2MIDD8agnT4KkEYLMqGKDkDl0irTDEZk
QGc3K0F1yTKpEehq4sz0i5R/K/+o2Bv3dMkieleCeGfIIK8nEs+jDp4PCUm50OYc
8u5FJTgHxx28wZJi5DRNRzrWwB8S0tOe5wVgOxT2FoJGIdWv0+p9V8KEuOW194tK
k9zgpA8xBBtFteQ7NNvk3dheY6xKDFhrplN62asBMrQRp0kK2MyhI+47U/zLkWH9
5xZtN8whCTzBiSSr+FJ+jQtAx8Y0ywC4k02uPZV4+wb8YZ0VWMfXcU0uD8I69dzV
bZQg1Amj/Kjk4HWrPRWEJwMPMWeLXcvaHw32QR1sXbHy8HrdJxr9S43c/llm23wR
q3oxJjP3q6k/I3WrDNlT794t6hpsEbDYHVRl2uKuvjVH3Tnz5l5LZDwXcQv0+mk5
q5HWeCP/iOJsk0mWRwzyuNO2oelB4T/Sw7K6tcwxRaNSqkFAw4gXSLRCLQpBv8x8
w7q1Xt9ZiSpjbfIcn1/DSoXTcVG7yk1c53iFhPXu5d180mkz0a9NY1p6GrsE6ogE
8AZu56xLX+e2vKfyhcC3d/dVkFTPuiH4QHkifwtGILXunb+w/eobuDhOavy9Rrom
kh6QKt0wc7PKE3n6sESM54zmj8s7iFh/1M3ZxxUCkYj96ntVpHn73ajw/mCw+Eza
Z0PpU1+UUlHHdWcHV1Z8Nn/5VXhBg/rNxh9PT9rxZIuFI/9+HeBPUtBXG6pLJdHv
PCl5RjMgEYGQKTuFwSWLTl2yzdq1v36XD+wsyg/sALq7obXlOPMZPWGrxYfHYctN
jImW556NjdFaPjWuubcntofQlh8a7uUb8IFXPKgcalMBHZ8ofxJvOnjtVAjV2WL6
vu40ADXouiUdgK5389etAmjpU5iElCVlOXBkZ9f2kTy9r7q7z+zTHhQa6xAB20/0
4jM8zF3KXYTrd1YzVVMVwvrfMCgqU54Za3QIf0IzCfAn0l4G+aFU8+HC/Foyesp/
Womu7eNRpWSclYyDB+NPUw==
`protect END_PROTECTED
