`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjwJScLaKy6dSNCi9AgFKT4hctW/moSCW0SfB4+aioLzB0y+wzUIzm8l/PSLf1qB
HQHS4kqG9P3Xs/qVWZsGJ438xnMYRYHWRAtY03tNKZXF9aC1pMKuNH3ndY2/Bkxl
5F2ospjWq9gRYrtiKVwVtswzMJFfPrrGdriObgqsppsUneDSnOevqy8eUjUqMZA1
5NiegE0+h9IIDAIhyM0XLYNJ27P9JJqzeZRjPIqwyDcmsHitQbJh2aF3i1N3Dvns
pxtU+T9/JbyfyblivMa6NZeObGxbM7mcrCHeYnFJfQoTLA9+0ViWOusiqSHlnTpV
r9oa95GaZiiSdzcyzBJaQ7YMpXaIL2upH656XZhQ6WLpZIhsOxxyKnIHZK9Ge/r4
1d7vYq1frP8mFB1trKIRsfZTg8+wD/93r2GfC0ogNrJYu3AyY0maycS/lN2MwTvV
ZTMDqYNZDDWc4714jHO5StVbhIEi2QN5StH/15N01nRNWemSPAt1zqluVVrjKM+E
LPoqftb3LsGyr6ijhlu7pOOHFBsDKA3D5j+ymozBpo6bVLJvtHOCFxjQaW+/NfD6
0noPi1KLiaVZsWFNrJ2GrvgLyBUgB/cdPudMJk1AR/NQIpRxbBqzoiITnsOZQ6/q
Rx7wd1OXWYW9zZjPcXGro8FXGAjJkOjYUZanzWf+uUe8Cb7NYyGk4cFj4vpZjqNt
JNOpoY4iW1cIsGHDcGV03C3pQSYFqdK6pl6YmoPhudTYAELuoEjuOk0vxqY8xSwu
x1aWiZjYIIl5cVrUsBlWk68USoexPehqPAxwQgsuM1AU8+VKK63j1OJaVST9L9QW
0sBQ/ibWsiohz+9CYxOHHYLC3En2bPy36RF1tFiibg6sgcbQIRdtWFqSeLpk5JFc
NS8x7jIz86RoT81HTlRofD8wt+0Fy0dlizc20YbY82yxGz4bBZr/Ji8HhpgTNhgQ
08nk845mYrKmxtXw+52/cpZPYtYatHjTQCOZAGzAr0/5FUGidb0FwVMtJ2xJVnME
nDoYl4+/X+ria/UydbUMg+3GldO8kz17u0TPB581aemArNqC+J2XiOmKwtU1rJ9i
bvy9oU+OlkCIZNv4kJ0hsRFDrucF5gfhA2HwGNDTDu4gNHIGZa+y5DVVOEO24Jk2
oq5UJn44S9mo5QMUELh99Kxaw3DSPZpGGUOgeXt/lhxpctWJpGkC529f5HTFeaOu
CgVDlWETZVmLomj5XICe5RBMc75GMOmYZw0MF5w4DVhcTmEbY+laC8+uKb/f5NL6
JMjF+9mRQKYELJP4Mprqihc+Ktjr/EpLnDgVXNBNgkbAr63mvdwHmvpwfr88eJei
iiNvMjPD9uyJ1O9ooY2hk/k8AzXBuUWte28mFAeAVpr+vkYgbdX5kVoTm/XlxuX7
LdoyAXWuaaq9xpuhb611J23SxbCObhS1oGXyYgTnvntHcmBE4X9owR0x8HeJnphy
sASPakRFm9jPzWKfxKSk6HF9093Ab1a80WIWwJ7Yn1Z+PlHjAxLbynxeRmxZ40nE
xP3So9B2Yq0nqRkkvEhfm3YK82y6ntrxw7BvPfE5Hx/vee3woxJbA37py3VP9UMz
7VKaqGkCuN/mtQSK1eZHHI4PFk1g0K20FL0moBCzwjxD+fmRAZJn2fwbPuaizFJX
WfqFc3jllgZKK+eGva+YjoKxx7SmmAuVh8IskswlMqBf1Gl4OIyuzAMVgUWfPYeQ
XXALq7f7nRoIuscTUuPFHeoWNp3toUCBUXWG/4X370ZJrGUWqn/T1vyFJCKbU8hF
5TqJcOuOz6BhNyDJjvbhklow3jEv78gkk4EBcouH2uM=
`protect END_PROTECTED
