`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sI7mHY0Mb8hZsNtVeaJ9NLo0YOdk/dDdrRVJLezE+8nWWdm5uFocyttPgMkQVmnc
mGq5TH9Hzp9HNcg0dgMSe8288YAuYUFeNDngyum8K1IXmW2+q1HDJ/aZSgg2RKJg
5vcTUWLcu/c45v4hRN8fWOBVx3ui3xAQm/msLlroo8VvkbEObLsyC598Fb4dQkKK
Oa/6v0LcErdegSpNwohLFUjDHYL6KcIZg+zmcuRQl6MZ02mRvQw+EyaJzIDF7Hwo
EuR2xdnKri8JvQt3vauugjGce3lvREpJrqLLe65BPIvECNoSO8NBE8WbdtqmkRn8
iBzCvyjk4jRhd8+5wHK4V2rBB44JgLDP6riybvpXyTpOGfKMXimslhYgk2N6I8M+
pvvY+QPB89pdX0ZnFARJuyE9LU/XQys8wXaidPgm2j+fp4e/Nq6WDBT6xDsafAET
0GHRjcUTqXP2W0Q0lYPhbzoVcSiwL/eVyemwgBuOYG7R55JnTVA2mGpwUqNaURkU
q9BNFqX6ee8QVBVPi0Ek3PGHGSv34DbUddjmMy7UreVs1wmPY0Q0na8OJdwLDVFu
N1r4DLy1db5v7UwpRK/5u1EtMsGcT5e0zBxjTjqfyaHHryW9TtAJVXIwcj0W7kU8
4J/yg8JwsnzOh51QXlJkL5Uxkv7cb5rUkdRcsODQUk9NMf7h70+fGTyzHhjqB0lQ
+0OC+yy26GXuBvNisBqDNxEM6bt1w0ZbMdABytfgdQL6dwSVDYN7nbMEn1lZZAQS
R1NtsMl7GzijilyfRhE7mCeMqjBuvQwHsDkenSOcqIV9t26/zW7gm8s1QN9oN95+
R6k4KR6CsPBBLxUET6Fforadf5JKPfz6+hCKffDM4AGzhF44Zvez4hjup25giCWl
cy0vfUysumPgy+xnSgITeYLvL1bQA2+fwxzzW0G5DNFfRD1sPacLwkgvFplPoxRn
NWfiFWx+eMm7AdWYB6dZ3bQkklJ0RiNhNYEabHLqtZ5Y+VFpYiJXkpLCN2RDLZwb
cj6mgvzPzrJa0sBODTK1zKZotrkQ9HMnJ0RAEJnCtqrjYYjEc0QO7pkVqeuMzOS7
fsBhmnJK6riHqQe92eWJWKF1C/rJdsINvzXekqVrQyntnsPaE/wz4v8MuB0MMQW+
XYy9r6CM70MOSQUQDE+OKujFCilK8vOY1zWeENXCjJC/saKMOUOfIO6gBepZTG+G
I+EXsE3m1tZq3brT49ZEOCf3T8MpFXUlzNQI9TnceGFx0iXhM5K1Dx85tlT9XfVd
jYwkz8l5Zt/AYpPsCfra6xBw6ktgH2SZWY+qvTR5R2Tjg7uTOtu6ONR8EoB4rxho
adFXPALcIPN93sVQ9yPqohGps8U6aTNcrDI2kWGVD9NGBmFOpbfF+CshPFodqZPY
4hQ8jHuFFfdLotRP35oALP2VtkGSrIHLczGjsXBFnSrmMX77zYOngB5zUS+n7oEl
BfzJOuyfAlUmA6X5jURsxDtfE7Q+0suY3/9XgEIgB63Yg3lLDRy2uA9WOvtddZjz
G9+spbQNwvqNn2UyITyflNjsZkoxsBX2wdQ3bGVzz36n+dnQWiuLVcqFHk5L3FmR
MFk6W7aNl6OotWhhVV73MybTj5+upmvf8fZzQT8XnBaesK3sl34PCzrkaXlFaNVg
nQPnX3gX2EWr+8mVe3E+Jf0zbLeOD5I028+Yhrt1Z5B4L7FqCxVUET813D5cubZP
4cJG7L+2JlXugqwpUo8ruIsQKCXNpnXPI4jizRc0sEpYY5PJHT73wMh7438OUsnW
eFLF43vnOisA1sg4ZVQp9fBX7Mw0+lj75rzJsprxyhgN2iYve1aPb/O492KC6EFL
VIYO5YH7E0WGSTVdkwHKVxePWObKd2z4otltAMzlSbD/2Nj0czTfTPaMIQ35Llgs
ImNn1+Wv0dRU1PGc2otXv+xDraSI8jG4S15VQ6jnqQzM6Mdw+9HaFb7DMYNYLqqL
N8BWUocY1y5JiYyVH2qV58TipBZ63X1zp0UM5sSCKEpQf2djQiJroV2cNqGsILRr
evZqKvAJxczI2BN5/0NFfXke0WGUyOYpTxiaWbWJy/N7HDUNceBvj+E5/evfKcbI
hM4b5fRo6Urd+DAWsjiIzdKyYpKj5AdnOFfBwZ+hqw9EAcDyRGJwbAP3wyVwKB3o
h+AB0tYUxvIGvcAQgKrOFKJBzzhpbohGhNYeQFcc2qaJlcRxHhvCNORTXfFXO8ga
Vn6ClEClAcennNQD6fmypKasutHJFyxaABgWsNUWmZb8vtzPjPsn+RrQBv04BsLn
WW9iMEQRgLXT1Y4/p5LkuhHRulmSU2DuVtqIrPgj428dmIOWa6e2UObpn7n4mPfO
fUc/AclIiditRYo/7ApJbYiGrN+eP9y3MQy7zlpTtfVdk7AlWBk3tdd706FYVAmj
QX3mXfry4QUbFvvT0NAr2RsDxt51ZFT+HonCBn9BAzX0XHednmAv11BKnT6GPnJD
krDQMYp3RuiiNDgZ2KMIqUtlbD0+JMQ3ASikIY/r10ulOAJ7WQPQwDSsbc6Lzmzs
f6ZkAvlN8YuPJ36GA/iNAUYJdszRnOB1SVrm9l8dZYG9GW+r6nweXvcmCtXHLvl4
QnymDUkhdNhbq7ScAfImUdon0T8kSWF4Z2pNu4+z/a8/1DJCoZ5FXOuXaK/PVxgB
u15MduWSD7h6ql8twoP03x6l2t6/ADACfSel9WSX3wkRtbG7fy4ZAFPwWFiuhLYg
VHFB8T6uQ5eAQ4b1Ce69B1DcJG5/mi8artgG1kxh/2JPZJpq9WjQfp44+IjwbWyq
cyNk1v09HIegaTfxLaS0VbzwWZC8q7OiAJyxK5x/ptIgWx65xklOWrDn/Ni+8Fxh
l3Cw5jETzvczSC7ARSeXW8/skrZF1GaDFVBO57ipA20rNq9DCOZTzhoq1o5c0590
9tIoRGDOZoToeDkXaXE6WG1pTRr+s6eCDB+YWJHha40HEOYV8C0XBcpUTonZwzNJ
GyOqFmMaTuhnVrgm4k8XPwMB7Unw8rpaxZgV6ylJFjAkMY+5/mbMjS04HQrLH1jf
q4ucO5FKZUw8/wQOmr5R+Egx7Afpk0dnnj7HHhk9YQ4u+8FRfKPj2knMcMS2sobU
Hs2HqA8+uORm5Qju9Xgv/wpL8OzfeCqwDnNswXAULF7j+L8Wg1KvwPTQlE9Fd0rR
osDg1jpDJFkMtEc0L2iKqNEiei/TlGGl0Zg+8x3rVmtDxhPUjg3sriEdOJI8eul6
/U8nD+7VV3/wZG9B1Hhmb1AUFefN9MEKi+8kwVfMnwVuji2VPJ+fz4/spMw+Fm0j
1BfaK67SCdrD646KZ44XzadX2aCE3WOeGp0PXc8arqUySSq2pw9Rm7Z6NkNM6tg8
ZCBrpz5YCr1qxBLwprYaQ1vQvswHfYlZRq6YfKBWeQZlpJjJms4rZHIBfJ+81Gzm
+YUjPDgZKIRq1xAghQgHTqR3tADZDM3P0THiY2ptZd4ippf3wnMk7mAzlRW4w6WH
nOeG06IHoqPimn8Z6NNXpjUuXGvA8MUIgWwFI8vOm47zu9ajoFgAUhRCIIGcS3Mi
olctrA4P15XBYIcG5KLBXeqfPEy2Vvs3xnQ+eRnPJ2x8MrfLa2qZTCK7IQt4gAW/
4/vBKSeqVmb4uNvSAcGQbLY7+V/NFRDBr903XUBQ+BVcjSdp1qze7bihVXwKowED
CGf8FnAd6EWRHuZSQqqjvyi1ewgCh3pGH5Dn6LNSVogASrcvGTmiLiXk17Dl6Rm/
9EYwxt1FRfGGgsXfBiJfwUXmCxzWfDvHhdIXioTfVAFeNaGOERwCf8ECh+5Uo3Jx
nqiCU7HxdY4iGDU9vL75poQeCqSX6YN23hsH2zo9BMbs/HRRPM0JkDsWD0++P23u
7hUqAGNwMyQlgELIJp4G2QlQJ9StwvJGxuFDkDWIgvFiOAMD/yCjLABpPtfcxMWY
8ICMD1Xf09Zf53fWptW2v+DJDc+4EEAJFRHly6StXVKxnrVK4xD/x1xKXd5ueWk6
xYqF5jRL6gU73G9aKXZni8PggRsrx9ksXT2zoa+3T6c0gfZGUocZhRvRB0PvD6hg
cKn52fJdgXjqGBmbBEbc8KXBjMXhusXMKGZh4Xd49HC+ESzmRRAuC6uxYJLQaW2l
rbrhTE7ywMieNIn72lMYNCTLconA7YJNKZiM9+eydUCU3v/wSkrpLAZpqJSwJQrd
S0cwvNN49vXkSvj3OvRDzCXus/iEM4bZ2TGa7rAiO1QBXK/8ZAV+OuGgRve4ssIW
gymbBLsg5hutbBG3tgCrrmm/MUguLfC3f6zhW8Sz4IXRotMs7xN14jg9ySeVr8ZB
KAPtKNS1Tpd6p7xQs3ZfF4fX/T5Zz9QS/ee6gbTgWwqJ3dNQh4jA9Z4MW5YShgAs
0tzTb2hvQFWcRG0kVUDObFuPAqAiIB+d618bU82WM/d6vPOxPdpeo1kiTiEwVaZA
+udLKznZt2zFYIQ4lTtI9L7GhQAvq0UE1d9HxXiAc2FaeGtLS2PV3uRcp1F2nWuE
8Sb6OPandfMKNhGXMGt0Q2YgrxxDPiVL1LBGdQu9dTL2FWnWcYmcJzqhxsOKtyjZ
jX+8af7kKCjwwUR+I6Hr7FHJFYclRh3G3dHWPT+yLDFeBJprmzi1B78qbDpFSeTK
8ZxRG+dCsvnebWgvD/njmBBikzyIkWojjweFW8HsWlys3df0cyxqdWiOWq2OciAz
FuAwtNB/wccOm9kSR4ELjwalTrJfI+5qJZrV1TGVYjyxiOd3My4Mm4myBVls8F56
xb10prmOfZn3D6FcadYJmCjhIokL2NgxbKXLfGj4dXIsxoAVrgiPoA3Cv5pB+X9T
vjntsm8qVzaXW3nblNPV0YKWmm5Zg8Usu9juAjiP2rxyjlXcQP5tnzp58KoeBJLl
6rlv08+cqVnVVSnxSA5fltPBxAqBTg0CdH+YbjQuoMrgnU2HKMIdSJxB+xbYbE4b
IekyVy53eM2U++q4MHf0/0WbVUzGjXiK3QGzZTfNFh3SYTZ8JY9iYn+cD+i1MKOo
FwQG+/tjfx7U0CBCiCcBgSUFLjrMoLXhThV7ZvITPnj+OTSTGIgIixUwYg5z8n5c
pJO88wnufFFUqx40CkHCsPLFBkLYuYy1Fik60Dj/8BqDslepPbEiXlJc7jtl3RPC
n5X3ZqvQjVAeXWj7aiapt45VMW0FxAPkK7ZJmBNVP1u3BL0IYpH+Tuhrc7Ot982F
aU8ZqEPp6hXFZiYo6SS6qO11GxeG+S2kQBSUifdaKF7A8f4zXo9fRvU6HW9VP2oU
bpoMAcnAMwCK7aPKfD74Mg/YtBK5OvP4z7p1opImzLUjRiL71HtCxBxsjNFIeB95
ep3bKp6dCubfyVPxyKn9/sA3BeFt7RiPzCca/2Q8SttWZr7S6ph8R803dmDSXn4m
rfB7oZuBUWCGK0K93oPdbznMZF40lPbTF+iRWHn4+P7lgAZUOlZ1E2GbPCgSME/l
cwOhzZFBnMRwBkC7iFsnHChIYCgykyX5IlVHp/XzxhCFKVPSc5CFXfKrt0zIZRjv
yS/63DTvpXhFGazVKrqPuRTlW7NhgBodA0HOvqst07YX/9J8szNZA6nreuglR3d/
IIr3yv/SUlCLZTF0XPA2tBVyzmUk9/bNbKRxjehEmoTNE22RJRxZUs2I3ERCyjIb
T6/2TLrAEBu/G3Y55+WR1H1RT1twSptaaZFKgGpQlJKCSD3dgmd2H+EXxUHQCuzP
fALu81R0RZQ8NW+pcZD2GjXW1SwEmx/tuP9aAJHV0fWiXFINklj/bMtHTKxERdjS
Xi68RxskoVUjYjYUGyagLZXEwRm5WSCAuiAYGU8DkZELQzcikMQSds+7tE/bMakK
AuWU8pEfel2PR8A5v/bEBj6452+5Sfsg0Ef7jnSl7vjFRpHgYMBEcEKkdYkdklYo
IbfSVMlpxM+xpUoFRK7gd4+yn+pHQ5GgKRzskjQVOXLVYYO6NVEAeCXl6DELhmjP
+6sEsB25npIq8RBk4bDEMYqaJ4A20B/nfLFp3WCc8AccLhEJBw2j+v29hcrDiWI+
YGjrmsx/qDXcdBEHATIxJeXgdXWyBnCojdGVJhB/SdY75M3h4gYWxRb+nmh4oMu+
F2FiIGiOZgDKS3i1glK3QKOuiX1xcIETSw75nkh86urZi/CoI7uoqQmqRJaq+D6O
btvADdL3y+DqFgmAsBkYb88dkHbRUxYsfj0kvNqd/a5smPycgB04CKdgI0ElNOng
b1JRjNM9ZJZDS7s8WcTk96dXJcU3JbpoHLSktvYcSwOfIBXK9AgUxwPDNGqO0Bt9
ctQijKq/ax23eCN//CfbueeFVzQkXE3SXo0IQS1I1hEvL0bGTy64AfbBoOHrp2/D
3Xi0/KxphTL1nSL+Ou9V63kOylienGIDDLGNVxA96o83U3EfAJBsV7UkdiWaSmGR
bLOKj63u6AabDieuM3jsgTGU5cmh6OVvCDkfdE3z1fp7PcC8s2+2bw9PuceY12Ur
XTTyiWeHE/zmY9A3DcNPiNCI1yMrIxQIUTswGtkgUPJeNdMc2dH25DPeRgL0K5kE
b06HzlAVDyKBtGCDCV/zvB1GNUXV+JbOhJ3Dm4S61rinJAZxvyXrHSpoyymXVTa3
R3U0n+berWeAZK9jiwCLNysWqjZd5lz3r82CpHjZJ8nCKNHDqGkiwHKOA1/zRIxZ
/9P4RbAMqAZicyGNJlCrDxUb02SjX1UjH9UPx593/uh6MVjtufEGad6gqCip2Cyc
m9uy8xtq6MDYP5T+j4u4K/zqJlulp806IqgN5mc+i5EgGEqDQcV2QnyaovixRA9/
WFQ6TGy4GxatbQFb76l1Y1vR78vaAsqgiVNraHxmKAoPnM+nJ75p138UcUhL8DeL
lQtg9Pff+vC2IYKWQYrU/dOnMZN+s7tmF9hdUWQtmgui/aE3yAxlnCMLYLC4+0+w
w6NLaFj9QlDRraQWTb55u7ssNWGNFhx/FkSCm/KIF7R4CnU9KueBcMHGGW23N4v7
LiVKmd29E8LziXgkcl12sHH8bpLCuqXgBTO+Y+QoHXfIvCEV7TZ3UBRO8yD5t6JD
OM74ysxoUIifgy75TuiQb0gJ/q/MadLXrfvPEa90Xiu2N1CtAPgHFtHMNd3kKPRp
cvg4bIf91fXgCZe9IoIgoTrvtSZ/Lhk1uYGPNEmH/CvLO4JU5eJHuGPzLW3QMRi4
jnO7ekSqcJcENOGPQ+mH23N49NX9isB0HUOaayORxX2lkqqgbnbfbHEXWy988eid
WNuPLDck8i1Cw+y9J3b65bjGo+5fMVH82Gc0VAVmN2wBUdgsveoH90J4za20DsWk
ehouirX81TUGJCIj0F2uXBP+71G8UVcR4mfseO0QDGz+sEj8Y/PdBknoZhpS4OBR
Qsm+BqjlLihrHXHuENHR9zDHM+aNoJ83vr1/NMVr/lm9Fces/Z4YdkQajcG6YjL2
KDDptFeaiRHDyHNM7ZvcdFRSGJZ7GbtYsRVtP40Vk5Hxt19Yd0WbKEK4YZ3Vpvw7
Kj2xN9lx3zxvQux/CuNpsUQTuY+jmE2DCCOenfgVqRQVKNuf9ObhfhyOfmL3p/nR
ZvP1AApRrqq27rY2/OdKx4zGlBLbOCeaN5zUJqPEXfuukgzrj/HEopk6LhPof7XQ
Jd0ruK9jzWTJ0WSGmbjdjAzNcvI7xExqb+8GjeYUX9ejKX+u+euEOWEaW6+zS3PR
iezO1eXDHjUNTDFAhsDirptBNxiTsAFnhPK22xLOuHOM+VBfHLhl2IG9fHaOOzeW
BJt4bnFqwVjGbSW7tNeNdwFbD2WdRsZA1cZKm+WWKHWd5BXfEuxmQMreSyNygQUM
JYvCDkgMVGt9QVHU1TECeTeZPihF4vX+qnF98byAYRxNXO/8XZMUhhSS+e1LPbHT
PzFiZRUoPr8GZa1D/FhqyUxIHi9cT3DiDVE3XXrgIfGLtjZkHxh1LDvLCjjkKCr8
IGmh8bsf26P2WmVl9XLA2jGjjEjicaCMg0SnNuTY3igOAYseJodwSY+HMs1QmXaF
/gmvgXe6iGywZWDkEuR6Nc8ikpwVCyd4mEskqLgtqzFjx9+Qqs0kiKH0i1m51H65
uLetMG1QO/HCfAD982hkvMiLmLhSzFDqr4YKfXd0Q2bLdB+e9ch8eErB/nA3AWBT
RYhsA13Ryr677Yd0OA10i0UpNSr/NvHr2ITsMk4V6cOIFY/d1F3sLas52ckgDmTa
ND1dchXf4PI+A1OoJvRc4pULlBSJtG2HCrPQD4sUrfBtvCHdKrTVmygwJ0caSiMW
oIIst2h3++0hlyTUd1uxz4pOPkwREyJXU3LpUCTaMq2kL2aqs+6ocn3kN7ACnQLU
rfG2Ot1SHWkMKPLN/Q0iGh91yqEqoFWyJFBVsjQ+91vsJBXhLRjL/+rxme7nJ2s3
KFdHZUnXLEAzVv/hf4jARXTc4HD+z/5NRAtQszvB4F+Aqv//coQcq4nNaNyPeu5I
4puU0ETRoQHZCIWDRs6ZPPlZxQx8VlBrW29BRuzNu1IqPhuNAjyDkG0hD2/ewKnA
JLHpQmODOLzhYhpHICr3Mjhh0RAGC4fcreNzpcT99xd7uRJWHkvE9kFRVDIb5/yB
Dp7S7+ZsNr57QZy7Q6You5Fky4Lbdtxa45E3EWGfKLrU0gEvJ6ZWV6TfEZHBt1s3
jE6cF/C70c3Ub7IqDwcxRv8nLnXbyg98gUl26J7y33WKOWv67liWpWYyBibCJVhc
CKnkOAfMh92gKAf3j2alzdR43NwvRLoOHy0cR4EYJQXAcFNG/SGywTGqOF2qIHDT
6v8U1e9i5UWtCQ2ZRkZPxJxtxyOea3lXj5uhokyrpdas32qyIzg9IdljXxObS62A
+WxQ802XVy7JV3b2EbAvIDAMDDO9W4bdu9DzRnbrFMXsQCjNx+5BYy/HpzxYVBf9
sjZeZ1QCHXPg++LGy+JyxKYVrHRsfZGgzgWdnWPuTKNwLSdtkfKV5iuTW+dbNWop
AtWVg8u9Zl1rhJbgiCvuQ//ND+P/qA8XT8MYMcojpps21kZZ8XmhBhMNyKBY9mE4
JMdM+xfZOdAPkHvD9qxEzZs5o7CpaH9WOTh84L5nuGI/QnGbv97miW9MAbXz2qbe
DOBpcaYBGxnLbpqqxixZ45w54200D/v6/VXEa2B59MYgxxdn3OKiNrl6E88NkR3q
cYPh+AALrHds8oaGiXwUIx8n2NtXv6vx/byP4IAcLdtPNI/weYZCFXx5dILXfPJw
1Tp73JFEnn8uPM3919BAHKgWD25bhaPo1y2egxiwGckojQjFUBePx3ZB1lACYb2O
NK2d6j+D1QfmVBplgr5NLsxQ9eNdtRu6pDf39t20H/tVpCr7q0+2uTvmhy8b85E2
9kdlPFLIYki8QK+yXZFuq1YW+4QJVub5hWGiq/ljyisW4hRTVNe6B5u6p9kTunc3
oQ5byTkXPA0KETZNOzHvSzGOXT5fKOm3u8Ftl7GoHbyAxKuRcEoa4oHXuHSvJYtR
f7C5l8m0BzUb5o+pxp2GBa99Yx+EGRNJYIa+SXWcWFMunRKH33N/tBI5w3RiBUHm
RYIMRwxi9iIV09vuaFzycWqxdoD2xlphnDHbHDXjB9TtRaOG79L90EcLOhWTXWOe
Mzi+NV/1mLt/h9qOsPTgcOWjdCA6dmI4xG42yvKCSpwQUtCOE85ojV3y+9Bw0Xg/
DmO4Fn+Bxj/aONWA/iLqOUQ34H9uxitE9eB+CAvC3oACu8XowMa4imeby1eCxyIF
ZFsvHDYg5HHymHdPMae5Irx1iLgzGKCVfhtTqKbDfefytMRN8J4KxuxLF/fGh4jD
HXW4Thc4puQifB+Yrrex4CvFq7B//AwPDIDxE83ay2qyU+jUoLtzqxMQ7L7Hh4o7
zh6YA/S+NFpi9Fm85F5p6k8NiNap4BDi8y1ZvdK36d5IZsVvzLDVbG14GuX09tCZ
0a2eCqWl+QaHEzlTADxXd7kb9vmijGhh+Hkre6rlfKTKnEbgWtJmubWeK30fsuRU
dO2cunk54U8xrTzCHnVfsOGAJ41uXJCOUwzfiIpABJzOZJCh4k9dFFw0hU4v2oDD
C1pg80zjD5usxMEp2eAvgf5LgmsiuzTI8KxN9SdLD/jSa8e/U7XOGzdCL6sh4K4b
r4o0AOuEUOIx6NnjlzyMi0WwedUdbzI+OH20RSWFzgpBnbWRZTk2htvjd3dkkQ0H
I+47k6OrDrpDR5VkHlVIyEccxvsy1h3StsE7pUyt7jy2RnC2X3t8g9Hem+dKHOrB
piLA5HeskUNrxZZPhNDE6Lw9lZrZSo3yRgqFty6UVVXXU/Q4LBp/NNaXd9877x7o
SdMeK6P2f2vngRItDViwGubRwYOdCrd/YlYuXjwTDgBFB7dhlNDtX9uxSYbjqgux
m4QJc3chugWhBmGhKwna9S+77L2OqOWbE2k4cvk/cxM7mR4IYatTsiGi7ifUhNKo
rvk1UnQGdpH7CR6b0YI3zk+KGRHLPnauH7Fm2zGQvEZpTW5OnArJVWyKLHYZl6rM
NmgKj7r68gRNrVBloHd8MJpmxcdRBZNgZkUKUQWwxzhPDlygiZBIfAcNMI79qxYv
kwckqjeXafkZ6GTNRn0usftHpvhC3YYOlcf8QnL9Kc9t++iovlrKv0nmK+innZ4N
u+kLKzYF7YW9uhP5GcO/ErdvRltfY/fxsq5LoUA8A2aLw5eIPSxCxGQvZMPOsyZG
A2YAm/y1fJPj5cpOffoRypVQE0Zxf3Bb7OnbGGW8lJ7KESly2LWi0BX5IWebfoD/
vK7RhiJcguasjTywkqzppIdoQtbCizu70p6uMNRldHhQzr8rKBW4BUyKYR00BVjb
MiZJMVI3mwxbk7D/+S5sPDPDcdYdnNceE3QJWsaIeM3zB9SfXS5Zy+WqT1mwHMYu
JeB0u06lQnJhajd/Hgqx4lgVvBOB0MHrG2TsZOJbCWnuQ3+vkJWz6d5nws13QBoF
xIoAtmJ27Av2s7hRQ3X8/i59CUXyIkXGrjnoTYFEFK7LNz8PuG9bEqoOTwJ6vDUF
bGruMRKKzYK7nZtex4fHeWIqAe2PYGrz7pVzRbnBlYGpbVwFyHQq4PKBGpKIIr2Z
aZ7FdMF1jVvuRHBjxivFRjNXieYv9WOadjIkCPXDvPdKdG6d17rATha/iwo9XEO+
Cjxk9rz7zdIGMdgBrCsBP1M0Pfi4m0w2N9YsFUdh9DCFx4V24BD2fe6Xq+VvtjTL
lkWnMb6+LiUA5gFczhOLSzrOmNC+KlZsRsi9SWO5SXR7vIEDtvRvmSJ0Dy7tOtew
lhADzw1gKbLHKTiySRD6koGrKCweidlETbkl8/AgoYsPXoiS9SFEfP74yhdGQEvD
594/HsNw1I2s+Y1MKluKp7eec4uHFm1VjZrMf0f2BdDCH1KfEs0Y7snHp2EskKNR
5eLm2bE0R+RiPxkEgDtGGkfVJi6G/IIvEh2gWiUBEYzRayYJ3rEoKUeXHbhGyfpR
BsEDbxeMvwKpVAHTtn8G2+rYBN/CYtvoYNQqojToQ/sn6ESoabkFL1SqiSGW6RyC
6LUBQ9WBe0V0aeqdwLuUv9nexhKUs4oicX40WSt15PD4jRAnKv2tQu5tDsMp3XeS
IL1iLQNpWSKp+ZjLKVBC82q2zIfFgxy5/XgZ3VExv95dKRVdtRu1qGQBzWr9AV25
TH1ofyFhxEQSQepZiU67iqkaE0H7ZNSrGXU8yDW84cW0UzobHhdodEcxZdP/Crji
FrRB5PNipudIWgJVh6XeHKLet1/vOO9R/2TgQYPqxf9KYneIqHP2UWSFHJ2ZHRWS
ULjkEiVnFNC9cyXcHigLDkwcv+mlVEM+6qQVfJsKKZZ8n9Fd1ZLpmWprwh2a3OS1
mJqx6z61foZJIMZjhGx6O+Rsm+jDXgsj3JY5oT9oqKfru3k3yv71uTOiBEX+7fRZ
Iunx0yG8rXxzvolosTQPTvXMTcZ18V0x1yKEDifEic27F4hBGVVwD8BciJ9DEG28
aSRUTwWMICC3Mv+VmzdgmX68qgc92MmItGTOsfbwK4sEK5vX8tD4cBeOLgmnM4/S
B4Bb/yHC9ng5Xnc6vmXsu9YWVI9n/BbyPK0QhfZU5bJdCh6Tu9VFNi+QJpiwgUnD
qsZr5bqhI8u8g6kf4cCJ2OcW9XyJjcEX8XC5Lx66c73hG/gSRudyROFnHyXqurzl
5O9rWO+/xkIDx1ljBL5nt0hKg81X5C6FTbZ7O/HIarT8wcYMzJeHmWg/eJPXuVfu
b1LbOjEihmCCBRTKsQ0B0/1cbv5tzMkZqwVnMagXTC+vp5ITDF6WgPiuBxfr5UXa
MY1iD7zOcjcJ1AAtfSoAV3h2HRwyDdgoFgj5xdvJy6A2wjB6BJADbV07le4h9nBM
zxzJy8c30Ei9MskWve9hAEslE+vVjdLUWHXBeh4+smXIkz8Uuf4am8nn+x6Id0Vp
anjpxWF5CX90x/IbowckRX3bJXBNvOz54OF8PlP6ta74CNrvz7PyK6uQ20186XFA
QhmHzmXag7XNmcME/OMwxEp+8vKz5THPakE0ZYSYjlDVgcMCCLX8Xhc22qBWeAgE
KW5GcacakdehRCGOEs3EM4peLijaAj+seVpfhIyesAdZ4WK7TUJE1AC8CkWT6wCA
zbnfroJ2HUMzjROa/ZyQt9iLDGcouq9zGq++WNyc54Dxze9VUQLDH8qE/OSkU82B
DfbqaQMiRLsvusFpHwYunsQi35alC6NKPemooWFSNbdXqdu1Ig+7GETFSnc78N8v
LjOfFDOQDuyK3gQ+kuOv+tB36jUEo7riMkOonKke3LIOaSpe2y4eaHZQTbLTLPAQ
4KjsEq6QlRttc5Z1FaBvk3Pbw8whGbKaZaPnQD0zbdAwSGP9ycETBpdqwswPZ3NU
rl+9OXKo8FmoKVsseahB98GdV+IEQ7UX8cs94R7BGYSRjZqUIY0j/HQG/r4VDYQW
k6NqtLGcUjTrj986XJbnrAykq7qpV/oTQ6osCZpcOO9jmhyNHehuyoiVN+ShGLbQ
HnYzUkM+xxFOwhfR77ARGBDgcc0DdlXScfnQ7wUvBrYVyPO9kqoQr1oy1ztLGwof
Kt05wbtswWTNzCgFr1F18mUIhG6JVcWZgyhttvat1wiDxk3YJJJq3oJ2SchrhfY8
BUXiy1zVIMmSkyzDWpxsCtO6uBMKvnlH6AFfLa8UVKJwTJbBWJKFG3wW/vJBFnjs
dpkuXKUlNdt+peGhEeLMpoBSZFTcNAHrSjhcg/3U0F6Hz43ofcXEdaEKGxK4JuAJ
qSm/fDquZS64K839+dyNIrtkzcEaT2jvTZTZSa+VCOynRSC7KyXBw46ZE14FWkvm
bYHkU7kH8Kr2kUnwR2hYytTYyiRYMLA6FaA/ZGfG6ehJCc9MzKdjEFWgw+XM+SrN
uC9SPWPvIHHOH/HcRERHveh+IMtM6mEhr7rdNP8sLlhKGnTaAatsBG4wZTp93NL5
OVxrCxwjWNxeM4MMB8/MAKWFdd58/eNZ5NlB/PsdXr19vsPRBnEXDDT2R79Ps2Me
46RvQttQj1d1KcJNNhrbux/LMvX5K8PYka2uZZH1wFbbyR0MrPFbxBZxpfAVP+EA
FD9rtTVQukWudhSMKCo1XUUzGgzUfEYZwjpILpthTe3UHeBbBY3P+6MIu/5xP9jy
aAD1c6L6iXHsSpl7omCFUSPOJAa206zLWIsJgA7j70aQamuQDRiarAYWy/2cjtj0
LcSMDUWIUCvcbKA10sMKxtmOK+fflnedY7URN7jHkFCHcSXXInwg96NE484AsHP4
3AmRYeOoGSmjaVKKYDwxw3RWLgg+2orfeX8iwCJJd/cvqLVr9fOCD29gGDPLXD1y
5fzJiwLezQcBmwmgiHW226duudpzMy1OPXb6+FaZh26vE0Qa85UxBFlVosNZPbU6
D5hVWXsSMD1ag2/5g8qEExK7Rnt+0mG7KuF7k/P5Xqndqc6VMY9hnoaXZN9/EVYE
h/GPK8Ru3CHgx7UsACLxS+SXoUPkqMhjNq1716juxpsnLZfuWEC5Ft74fzYwA7Ox
AZS3iSaWnk3aptBzzvSBEMC1uZYv7jgl4N39SKA86+rpAo4FTkB7EXjjFoZU0faD
2Jj/2QdWMP5eo91DsRfhE9P5sD87IMS6yRjeNaIoPM/SivFjm1xjag4Zbtuff44V
hPSmWMzk2pM9TPW6ZSQ+2opcWtYTwBxnHJIJvmlKz82sHBFIgXnuJQHIchodvshm
zAUjO3223j7lFsQThph1zhxM5Cw6uYB8T3kjkjDwo7yKxPSngRgVkL1Vh52MBYT+
/J/IyObqTXguPzFXZ1uNcpPkx5DHtFI0qWgKAyuqw5zuSaHxqMRx3aNYjP2TPl9P
GohimFyKKsQUQivmpnCST0w+yuBHTPoxC46IkKoXRCL88GShpfnUiw3zjTCHyQ6G
ONUvwyhhrLpMI1thiCF96lzIhH9gd6aYJxSelHaVKUUOyhnopHIaUsQv8g9i9s0D
bQq3/GUiH1L10wCsTZfISqiRemsOGgtza90Qak+Hfc2fJ9B+S6B6oKrAQlEY7Deh
q8MPwEWHVLn7nXYxplqlrY5rBwrBMeOTsKQOgXFBELXi6VbefPV2smg/pNQbI2zq
c3UmixYFQ12vsbfVfRu/1UHrSiZ5PDCuxmJZBc++AtvlhKvjzD7MMREMz8vywEFx
AnIyNuP/RqwANfebGdTZrp3mvqlPTWPaqNCnVy9dzfVsQZAkrsBTBgTNQfIfsj1b
7wa6MZ4DcUifleAIimRbphozfQgJtVqjFj5yuvvegnioyLLlvkrIiFs38x7wslhv
+yjDz5YTbvaKK8/ZQrI5CxdJrRCun3ztrnk86PC3iXr/qffco4RtQXlJO+tQxqDC
lTS+n1JNhGAqkP0LTJNkqq4crHFs0ZhF/QpYAM8gYS7fApPuok2flhALFYTduUdC
larGvzq3pR2YJ/cUQ/2spSLcJwbjLkQ+lRXaMLl0FZ3yYGl0uIqXvgdkDHk9llb8
8Fk6ma9c3+2tGRO+H6LUmoNMHcvvz3GoEMy0VHw1xmvUmaxv56igBZrb0x5TYWIm
hzH11YiCPR4PwCU8tPichItSH0J7wEMUK7liWy4EoiigUzQ42pCAMQsHbpmbgmte
SQpnBuClh6MeveYWdpuyxYENcy7enEZCH5AlM+sDstmA2oelqNeWLuSGbw+XB2EL
vnh7VN1wwXU5msTFDRfLQSqHuKuyJa/sUrljx+3S5V6YtLTD1vxbvKMBkz10vgeL
FcZ/k+P0qkBSFfqpMD7hTpg33sjyJd5/zqXRXCv7e+PTbzD89Zm8dHJ6nZgYRp1S
/sRlvZl3CBvSWQpvuOUqeu2zzT0tRiw3j50IfESu7iOov+Au4nreWVyEh/T1U2Iv
wk6tpnmp6ob27i06eeKUr4/+tnQgSFRwpRIuASPJgdBkkR9teAgpTk9gaJ4ZV2PI
gngIft82faYaiiaB6iknibdaUFXosEPhYmTIuB6mcE9Qbr0BFMavYek1u1sDsS3F
yG8Zm/j9/SqHqcyJ+YyIFkDhllWORxqAdknpyZAzeJD9AEP4AJfFFzavm95WlkUm
jIaUev74tETau7gOyOlCLDCnUpr6PncIEQ0mHdStQj/KJHgWVumPWxUOaYYcjM/X
K+FzfeYVnbaI2VHYxzQI3Sm7yf9VTBFn2JrCyHDJJEdyrJoDkVFeQpjYh+OFeSU3
lL3romm3oSDg84Q8zYcMURNyyPZmMhfgf2RATQJN+kL3oZcQhCjYxHP9jjNnxDVq
d68NzwqtpDHeNR3J4Ox1BW8nhRdMW92Xu1rNARDfxm6zZOuKG47lrYN+2bkXE4pY
0tJ0mn1WK0Lgc1Dbl79V5NnjSThyX0wEsWgSIFqgfwUehAO+PNUbwGOIm0DPgqtK
O+hLdOPOnQSNjvN5/b3C74LreaScnmRbMYqBjGvoCKmKIf/APrDXJmFp46fl5Tly
Dh49D4/R23p0D3jMG9Qw43o1vGwoa1uDklNLpe6edFYYog6O3V62Qa+wtthApYAZ
uKSHwOkKhU8fKQfG0p7nI1duZRh868CslUMqrqSnzJnDjQ27Br1AxFatYbZcCodK
LjnBW/i8sZUcKdVY7AO7uz64atxSQdcnwQgZkG2ULel0PbZY1uMWxTrhFOdMOXp7
56jL7gLvhs+Xjqi+PwEWeUGqhvLn/zAUaOnenEDH5dFHy1U6NtlSjIhJHy/rJYOB
vb9Hq917cKkdAFn4nNJqXKt3C/tsnXZvPlZ3mZ6nsegdoWm/wR+YPLULU+E2WXyr
6fVFUohu38eB8QaHITDqB9a1s1afx7ip3BDn0isLHB6r8WGu7eySkR/DukZgiP2s
d2ZYwbspOOJib3uNLnX73yVRSmTNHLCvdtCDRwEhcGghPFc5IsaFIF9NWnALCVDb
SOQ60JNn1ffSDds8JeJJvkIKT+opYuwoIfp9/Tj6pdZq5Ca+QHcgnpII5w0NNtcU
MQytv/iOdqOyQ7SeTh3IMq1h06iT8QAjBq9/UoO4pViN8kLRTyRQYNcQLbsG9iqJ
iqrroHnkbDWjk68JMEleCcdGa9gFdVN228+k+c1X75pLAQbP5Axy1sLn/48buNb/
n+How/R+Fj7RTRNKEDGrzlTu881yPqO+hbuAg69AsILZi1HDJKjeV9R9bhAdQ7N+
itQpsa12cdsMBCfi5klDTUbftXFqdQJFEBN8vB09v5zOItv/KtL7ApXFKOAKL7qU
HgUUQFacdnpilX0FWQ9BIJUfIhxaFl2w+ji02vhy0UwNs5nlDcaBC42QJtTdXCi8
iSDKLSVWCu5wJAbILkYIR0nQGkFCJK+xrk4cZwaNSUaRfUTmFv1VRjGRn6kjkUAB
rN7jyh+s77qPhLum3l6mNPc1ZWXBlfZfjHAE1QvkbWWyrN/mXvTYXcNaDp0kvruZ
yCncf3WCFqVY9hftw2eUCUUMAKuoAIcSVHSFfEHj03r07FDnHJt1yn03rRV+JqR7
KmXI7fxCq/dEhy3XuswSVKW7KCB+3+6RXBEzdAg5/WzlnPcN+29MMOTLXLRIXgCw
UL32W9k0KOjEuNJrS6oix13OnirGBh8mnlXiSA5CamaZyoYk1v9kvjA8CjuJHa+3
vMqvozuxWsA0EZz3svHrHxk4EOct4ZS1NR2WbY/QoRmLVYhaF3ZKw/P9x4eEix0f
cZTZW1t7w7oaSn0KwKCtj66yZ5badZMSr5XtqVOT08xdx86JG72rmRnEOYTIOTgl
t8i9KaVGiCX9dZY9PyxptjjvsokEOfkgSBOt/lmQ5HajXMYJWxj1w1TSnS16q7wc
TbVTUFEorwoHuqC6oJmzEmUzVI7DfRzpOvNo6RUM9EdrJz/f2jHvRdncMXfOGrWh
G3eFOWA6rfK2FQA6X14ZBrraQrW4zosvO0jWxpb4o+s4M9QbgP3exi/EZvfPFECa
fKKAvdeAapkFez0e66xFBmTFqE8W0ff8GMcCYIsb7/W9TTYcelCHp03xCLvutiGN
oPNTh6NM24trFPfsIpyIjt7qK2SWJYJT7GQELrjIZq9AZhdP5NAz+t6eO0rfiAoS
8NZXSFjlXwQcTq0eJ+lQaG2vFFPy0RwH3gKa7YyFGKYGEZq8gtH2Rb0/EL82hfx9
1x4VkQiolzILUN7vFU81PSBItEljq6We/YGgDdCwZN4IoEYt5xSoyNaadXF3jtWR
rRXrFoL1DqqdQge4sN9Kp72rk5catzp0OHjv8p8F58AqAgGCs+8+KW7EFJuMcdz5
ycD2OwK0S9S630ZmSi/yeHFOjeS4kxZ0ORzXG5L3m6c/4g6l1/g1/dg22LRjKO5s
WHwuuJyHGecx29W72LMkC+Rt22Z7iWd+u04ZiYmozucL9+1NWcS9nneKKz+V+m+Y
V+o9MfBC9hbUqBTKkbGzaoBNxUU15+d3VuR2K9vHFsqS5nUU9B44iOGm6tS6ohZI
nKbug6rYtEV6zJ0Kc/uQi8XdBji/XQV/dNI3UN5ElTA9APfed+SSJIdvcxd6+eoF
gd32aCja42YBQUFBdc02OurnFMWlheOVE4P4fqcDaQOGbZLxY0E6JvadcVz6WJsY
9lxIezg+HL5vZQx8xV54AxDRR+9V2NW1TMIa89xzt5Wzq9orJ0Tp/nv2z8Ch2Rhi
uc//1t92h36s214zJFjMdsStkAk8kkhlQuObe1fI+r57snh7U2gci3h9tyEQpIIq
IvCoZEgjKutz96387MzFC0BebKkZqsw8qtlA3FFxXGLpC3PXsXT9Sc7dLqA3+GGO
wAoyaxz8ZBl6Yoda/0OzEgGBmMDxtQtoY1HpEPm3PfTrubhxUwU09hE/cTVkxv7d
Yh2rkIGOYUX3+DVnGRJM6NzIXSeawviuE5fIo7aQN9XKsL4NDSA7Xm6kGsibkEQ+
lYTC+x6jJ4vEns7tTKSdN3NCp/w/t4/bswqq/hCxDETyCrIgD1a+Sm92awDfQlDS
zsJdAjtCXKXHijIjO56s3zgltiOOQV8e/XARJbDjO66z4W0qRIw8ai0we+DjMawY
rwByzkDTkUcA0MqFzZpRfPdeRqj2MLYskZkAEoDMhUYxCmyRAupzFJXPKK1mw3K2
00G3uqVxFLs2bTGCt6Ik/Dj3w1148k4CkFywZw9T2oowS/0lLlAkNYBDQccHK7lV
wv8DK10244+HITVl149F/B8lJkR6q//WtQ2QnBhVm63nq3ZEUptqJX8vh2HwjeWP
GH0YBO5wR1YcRmt1K0szVRH2ALMZe48OceWYbrDUvkN2haowpc4tnp1KcGBvjbJ+
sZXbaucWLOU8F3XV45eRRTrB43yvxosvxORN7Pqfo3yMVpvZXo0W4uR/DxYrVyB6
li77X/EiGR4Z5i6rlWRuOyrKTb1W0wMTmg3LG9bohfSsuYIGAqx8bAyEtY0PjawZ
RTQBRAu2iSA8X1UTuv3oDk5uTG8wvj6S/FSi79jp0lg5htTcZxfKqi7eSofWG8hi
proEc1ijiXLd8NjPcwCZ7C8AAJj/2bPOI7TY7Iy3m7sCouWnXiv7ytBb3agOrw6C
VgxNgqzAiKrNN3PZorJoE0PQiHNVmgTWPWYQej05BMy2lvQMQhcwhPvOJhG2gnaV
Fhg4yLXwAJj1k/4fJxP0fPqf38dofaQJaK+j6KTmt+ti32t0Xy1IWwhiqBz8tVBq
bNCQ56WJet7HqK6gWom0nJ/Q0a+lseZ8vjP7NzMSzjRzm3GZmoVDgcKSHVYm2DeG
hD+dEeWYvP2HAkdU6hiqOKeJmF1+BkJ+1n1ZCOqDqA6TCvVnhIxRNiuFh2PDNPAy
G1SYKRqjRYcR0FjQZlQal4ilt/kzrvX2PitiPYZ1ZzoCdv0nVghom/QKKWVtgJ4R
5vFKYbPvU/34yLN3u2yDwepmaAsKu7LyJoMZj2NmTdaTXIDPcL4+qs9xfeCyua4V
7rCaBi9d8Fj4n/Bi0ZSpJEQOPmGCgKO+PJqgybyriAm+6TX7kJLJy6v99UwdF8vv
J3TCgutcTMKdFJKIcX9ExXXEScvp1yCthXncuXagVI811HibufoPFOdx6TfJTn81
e+30+6ECS9eIIoH616Qx3Xgk7nLWoKopIYylv57ALQyaQw7xKd3opYW+p9ug6XAG
kNt5w+/iVCHSlenRpJUbLu9HdV/l6wZUHcJnV44XoLdcJAQTcXlr7cWdy5LUH5rt
Y5zLrWdO9m/rQpT4eQlQqv+a3MEIcJ6K8kT2o209DeUVQksKUsqBeJly+p8VKtIX
61kAbhuB5dSh5Mz4E45PX4CvZfQE1ZnQDMEVzOFj0AzgpTOpx7YnOWdFFKkrzSim
eA2PbEUC2qnwOmUvGL/2aO8EBrU+5OSMgnPOKnP4YPoCcDThU41WYjR/VMKlEbWl
qWhcrHhS8s1/PaAOiCLWKlR0ScrCl4itFxhJfzLe6+RXA8+68WiGxX1n0og15jUg
Hpv7Gsv7R0EqdfqiMOpxm/v4X1jryG8bsdv9D+6DLm0RL3HKttqUWaayyE9ro0i4
7MPQrBd+NLy5Hn0ct0TSW2TLI6IpAvxRygsT3OcbPOiHjcIt1fnGhcLWXrOka3/B
k2LnK6vlWLnKMj2yaVh9phADxKMp5+rboiFLRzZXD912l4aF2iORWJDE7cqNw516
vrmaAlwinPoiPhJsmmcyzJGHEIFN1Ya6m9cu6NKfZgTP7poaiSE+1AaFYMvyTgpI
g7i7BUmFxSIHFIoqEPMOB1RO8NC0+yy/kBCjvm9ojJhw0128PHg7m4cnTSS5lils
8fyCwqirQ038GkeUaAe5N7ducKFWzaYna51WoHMWV9u0YtEmJLF+TIacAhhF9d7X
3gukgCbR9AVFhS4s6qQLEfm6i33zrrrDWU3uWzyPPv7bgkVTC3KFrZXNettXAR4Q
Cjxd+Ukj00OyPkoGUop5/wJODU85PiOOAQ6Iws/9+TehtqWO+wXiIfsrg/BL+Pss
Cs5Jil3iLXSf9foOrwa2aeLrtn0MG4fPbxaxcaLNH1a0CXb4da6jEAthkzHh3Itk
0aqnu1f1GSu54YJeL2B3ninRhe86Bquzt7GIBZL4sV/zNvrEShKsOiexvbt/Rtko
igtupv9LF2ii0IYzd81xVKDipIfBcg21TyWVlsp5TaKKXbYQKRqt87FNwRlHeVd3
NWe65fOl5E2NGNmzO1UqwBAz1jK53q/+xj8dKIhE1LihFY3jF8n0ju/mcn3EJybF
SNmyaKnonO9d6ThIzZg/cdGMm4hayhLHeoyjZ9N8hYeapzSyJmB/t5qJCVAqMIrt
m2l8HFVw94b/7VaIxShXSROzStAt6snW7e7iLqCiwNzLLJIr8S4l7psE3vMSUNMX
28w7wsuUyTox8h49B0gJgmo+EmjLVC6coyK02dtn0qV80BkE9o2DYz/KQYXVhSLx
UrRjJXBHedZ+i7w2k6S6i0m8S1MnMRO//ik2dYY+EXlvZZeItdhF6MTEWuYW2nB/
xD4mojex7VY61ke42GKIgIYhmZ5eIq0ZBoBKxw+zG/ENHkNvg7nIMJSUMRP3FKgn
5nXdEc6zG+JMgFWA0GcEGONA+iLho21OyP3KSevhetRnFvwuL0ZuQaQvnxjLdSTY
hvM55IKAL87yTJGx/rnhQprVXc8fWMppceHvJk6SnZw6xvluAKBL96CPD0+CXWUS
ZHGzScrCHAgPpd2ELkJQx1d18TNVsbuEMtPJ57vITHzgtYd43JoCe6W2yPwttbkr
/YpTHgze3oox/1satsAdHzo4mrhqT7sQAS89B/VECSIo1urFCTxss/cRF36f/eEA
PNxxray98LX8o9LYMPUVnkF4T/Xt0qvc2cUhsM3XdiUsiYjCllK/vJwE/es0ytuY
3F+cLnq+K4mpOiyDLxm5h5FGn+/AEcZc27h1HeX1v6h6/VN4zacD6r4Gc2Y0kb6R
1PcJzU5pgQM5Kml458GxAydFYVl5eRbb3vCRzQ59nW3Nu/i+uhFeD+tb6xQkHZ0y
DT455PtsBZg3TWKGF4/eQpCZSZB9LXlvoQKbtZ9Pp9e/dSHJqulnC1aHohLU0g3+
mx+AZwjyVassXfGpuJIO4C9CjhtO5hzLw1+cSY6uvcNxNSPCvHpAnd2FINeFg0aG
cg3b6e6zY7wq3QW9yd4z4jmuyeQNcy9FAwZNIZt/F5glLM55r3v5QsJR9VsYqurF
LZb4+IL+H/mkHnfaLh9fzg7ohLyiklt+JhtBvWa4f5dDl7/HuOFK8BbUqN6tPnc3
Hdx8uyLmfrzXBZHkuGcJB3IIHmJf5BNzaThV9jvOTR0JAPhxIjoO8/TJXCBLlaDx
kPdWS8rratUT/sqPlkByGhjnMHitZF9o/A61wyw9uySW2C60wOOJ7dXAGuFvmRXG
e9OosQ3KuMn/NZQAYI13HwsYkg8gdvvBMp6FmE32q0elRE++ueK+ygb3rZtu/GuP
/sYt3OQzkffC8jesWixuijpfgHiFyMLuFiXgxc7YKFtwKtzMQQbz0o09U7SNco9y
226jkwRItBxj7cjSIkm9LXLraDEONx+Mr8zosRLYIWrDADXCLuUd9na40Io36b8V
eVB6xUA/GkBi6X8F5wLkcA8uNt2ttVezfMJZNBH6udF6urgAugdT4ntHFGSmagx/
/8q4r4Au2/ZaVKWQonOxEQGJy/sU79DFd2ICF4fDI7vwOio0CRsrrcrfSNGgq4W2
e1PIg1DgPOVb6grq4nql6bc8imOxBADZ6JS10b2+M++XT0RnlTg9RP/xDa11qYMx
oYyZ4V6STIhecAJIKvtg2Q9sBC8P7MsiLW7XLPY9jyrpWEO4IZ9Ocqm3IgvcerpT
Eaca38VTcVbzUKEkHyEsETNCp3d+PKF7+jcRY+L+0uHWoSXuKHByFok2j8s/+3k+
o+T7yV76kMrXyjg1MCHZ7S2hPCT4bSSjfVEx4j4Sfj9FKnFgHiehxoXzvCv79oa7
aDPsDlFYHTjJ7tki0LRahP3KeQGswimYHFCdAopGvQ+CvXKD77kTiIbPUk23vI65
GHauBGepI0s8uEaAoclAjztPRLajxWLgG/mBKMBwBHsgCJmidU/gaTF0M67OiXUK
DhWm7XNzoqz/6b328YwZcD9X509AtLmyu7oHalm2eHdcZoPpu30A1eRhf/KwofpF
aEs/CS3xCsEO1I5qbOwlFyHBQKjByqR+ZONPPaNAdxBRRFP2T5tPjs5YoOzIMfoQ
R9ZmMNfrYBOZ/4CcPCcAPZbyI++N0qs8Vw6z8T1g4W0PWZPqOlnfg6DkLk0GWWGD
edMVmYar5I70aHpTqFQWUex39/zJy0xBrFODwbva2+r+xGaRTnd2e6blF/4XG/z/
1lAVr0hhUf9gZDXUsks0/CtN9WE1pxNR9P+w5c88Tae0qpT6odQHYlk6CarRDcab
g0aClHxrObQ5Y7ydjUXsbxP3cZVYXsNKbd4eJm8Yp9HD9RDWfKl3j8qBYnhOwkO5
86YWUy4Z573KvrwcN30SjvlMr9BnzcJuRqYuIiuq4fCVvUuP0rM1EmZV9YrTAmhZ
qEd95FmyiefieTXlxLALyRY12SpasLkc6uM7W+/0kMolkyhr8GBbh/zwR/s2Cj1L
0anRSwiM/pnO8R1wJT3/guElFP1mQ4oj3bPgDv85QL0fhRHp6f7OnFJQM/nzsMY4
iOyrEkew50UdElhwkKjuBO9OYbWgzNE2b0IPM8uX6ZU+Sg2LVv/T3bVftQm9wixZ
R1vd7rO9GqlzQn4MWCAxG+gmmZE0HETd2Mzzm8mCjouiA8VP/kB9PWq1s+rHySuq
icD+WOTKsYSdLWA6WvgCdcSZpXexdgsW6RXZqveFTG7QJIyx8z80aCCxbj1px9jA
/YVBkLToBweI1PUsxcBwqyyVMn4sLLX2W+RJTjwN0bYr/AuvSK7jFeVquH/TrEci
mxGWGLMsom7aHFQ1TDVKA4tisBvDjw2rkB2LwAohcLrrfOL64LuLfLAIm80Ug/qp
ciZHieC5hV2KTW6XfVK8hLdHm7saEG/Q8nebwdpzBG/6Xtvrf1f6ryavi7FIPWVq
wzFS9ZH/BMEu1W+QoFYzkZ1zVO55EAUuU28klGQg/CM6DNI8nZQDHNA6cBCOWQaJ
ErTrgRCYHa34jiqYX4d2XNeyUwihVi+hK2M4NSRnryWwoH7xGSACfkrAUJkZZMII
kJpVQKXHSflPqqE/9NF2GljENHVG8Nm/879doN33JkIIlH0S+8H8mh60+OUXk2CE
sJgfnBlZYps7uDnsoRu/rDBFKTh8k+LxCTU5Q+01zC/RhqJpLp+ArXgeNtTqeUwd
yJcrzVzJ1A2mxksn2P0S1afQmSBmWYHlTpmjFuXQHuPe1pa+uaip9MYt6NCa1Pln
CU9HAYyvxbmftr70ZhoksQsxy+C8BPLRLzc9DIJIsMPdpAXi9Y11i6cks7MVj+Ha
MwCZIWQA2niPcQZH7A9cPsMY6qjn2nJ8B/y9HVWWDnhibm9mOqXpaHnloGmeIV+E
cui6kBg54uf8uclkiJtLRMPJquDsY0tq+Xhnwxc9va1d32A+zP+m5WAZvkqYj0iX
zQY8Ahl2Y+ijBdFTsybiJl9DqtJq8GYd61KDWszPxmtxycqtTGHWyyk2pl7oQaFU
il8C2oO/4L/dprISB9jtHC8IgCATcj4t+sLJF1g3Byir6fIZ3Zx1kVnoNVtYwMpi
GYkXzV6oG5nUapq6lLsKzZzPkAZ1PeQPn4b7BJhyF734jYe1hixi3RsHs50Uebjh
+8f4N7E7DpCdP6bu1O0R2mD2wQMkt0Dh2mq4LU1dn29tQzfM+1Glva+z+UuHuVwr
rUPyjzS8Mq7WoDOEnRpTcBbZ+fOVqeesX9akvIeytx8icmw2isF4+CrcnbaEfxux
T03TRcnxuZqhGEv8VV3I1ytwiq6n0/jrX/cvvp0Nkq4JMlO1kQIK7b0Tfxy4IdkQ
/MFmiLaj00rwdx7QW6ece54CMivpeCc5O6edmRzVitWQKnRy/aw/lUq7MZ7hL6sh
jNkmHgfwYPlNgNpWO8iZ8pX6Bb9cfeghhxgm+iDfy5+evmNRbs6TaasceD87jwwE
tvCvURurBaDUinQ2upQddbTnNkx6kBSxg2KOnXwroqiETRAjgix52OabRKd6W5sW
bTjjIFWn8YfxIatjsFcpBNuTgojlSBADmLa0BdGquo02F44YtLl+0/fzhE9xGRu9
uYguDHgXysUQhX5dZHjMnJGiSSK+J3pC/udDGh7yBG8U7w6cBjvl5sxYLL082Lk4
pq9BAp3E/DEEI7uTm/7TrMKSC2LW/8Fj5wEXlnYWtZitfv7ON/bZWS0nn6YYlrss
dAQd+RGYPHZqfzOlTusldUkMqIZPyt/D/XBrxEhMB7+aVy+kecbznhVNZDRGYN2R
EJ6BxIRfa4IkL0g0PJevTdZm7fpwfZHNpXVE9lfU4WM31zduQYuMHCtgykSbbsFv
BXvzkYhucxi9D5Yn2WSRrBwHnVfYwunqbDDT73TPxSW5UkJAnBqZtzmV1fhFs5Mt
ej2I9xbaV5PQMZ/37JLwnecbAOTsQX5R6XEhG/k+/yGLr/DKSl+8EU2NTn7E16lN
6hyedAQ1fXV4FTzfUWeaW2hI1VlYJ92dCVNO/hd/f/OqqK84dinBKd4gohKx/N5u
QwuAyvNWlL6voVKPMXWKz3DxGU2iujeShitWXYzFukfKSynXYilaFsy3RxNmRnKV
c8wNRYB9rEm+plLnP5tIORy8yuhog3yi+h+goRhPDPIZG5N8TdCAdNL7nqzig43E
MraDwEBhdWPco3/iKwrLjLkGiLQspuSvMGtde49FeE/2FjZOXBeRsxrwbMpCl1+p
VZTWv6VE6Rvss2OaNOLGxGpt9XbTpNM+zhk94/GaBRYtRMk6CLr/CxJVHR4X7haQ
5LVxu2fR6T93S3KJOa/T06yFjgr5rYiEeT9si1cLRthvWXN8ixGihKTvJEa5iSgE
d4iyPz4nVWgraCZn4uWw4QFGyhftcwEOdb3zj3dib4PfsRYFxAPS5wBlE5j91/UJ
iDjIf12G8YS2dl7j/alYGbATrIZwuyt4quQLhN/WrWbOD3lUgME2VrF0R9gNIxde
rUxgR0op+B3c4dd27AKkBlwRIZz2QhfktWtZ+nuehE7FKriZ3yiZdTxofyECVrkf
4/CmH3VqCmkzWrFYgELN9HmQY+xUx8Cv1MrxZeOMC9Me2U/POMncumd96qXDdLxh
wEq4qWQEwGJPENrKRIDygdd+zcibw8AOkVuDiI+vM7Qy24bsAiZDB4pcljsbxu4u
arOJOC4RhyUzLVCm/QY6U5RUKFX7/a3wJkSSPLcV3Nz6SdSnKTCyi/R/EreKILTu
AX6FnBMmQEOSmtxvtcAHv7lf1JwZBwk0FP2Xl0Vw/6Jhm9xm5iX7xHvHToiuYQ5W
3wSMCnxmXkY3N5B6e79n+nFZxTwsruK6rse7dd6eBwfFmAnhZNtQP1Uv7PDstSTz
V4nDENVLkai6Eu9r62GvlYqWQEdyjDMWVNwsucRHANX6SHh02t2FS0qbLud/lxPm
hZ9D1IgnSA+XdvL6Kq9M5QCX3qxRThHj/mppB295Tb+fa+A+aIsgopD2HLN1aBPQ
ZgMIRwwhsYyDLbIWSyLCn3vC/ELIlE9T8d9ye9qs2BWeqrmaPeMbtW5O2eNOjcT8
dA5qVyuxFXMbXx5bLoxhEhDzLhzsTEKX3ng2S3xfnJ+CxX2hg01E1QKXjiAOU44A
eyDkXJp24nG+E7nNwraOSGrSTO9clve5y5BVf3ZhXwc/H0HPEelz9QeYVFW+gsvm
Tt+i6086xbHhRaLENLhe2C0iA6F2+kfHwWB4HK4UMK+XYRgxxZQHfcA2pNzclu9q
igyhrvli6rRvlDg5UymoUWFjhcuRbeX/nItaGbQQUCqnXCTGroCpeTU+FPYl6PCa
AMojPkv7Hbje0TVv8+sxEG5UegV1scEqE6hm4LynJ35nTMSTcy1n6RdrQOmm1DLG
60h8DwdhZ22FBjzeVL8sriE+xmnbgeV9mdxRZA36QVk23oLpJ701Jrdx5r8aH8Ia
I3rbu/qiZzOx3Iah4CWz5G9OkWksoz9ALF/MLxmZWFU9vqzX7F3h4RQkTIQAOPso
0NNPZvojEzeIiBd7HO8r7IfK3OvW2/M6A1HzWR7ft4AUuGdpfWW5jaz9Q0/C1FGh
V/phjE97qI9QtZfatdI5fswsLWn4J5vBYsiq9rrPyeLatssUDkwlL7HHTf6eALKW
NVmOSlUvNyRFrdsnR+TbXFZ9yZ0y70z45vp5brUXB4cYrv5vAOOE/MNQD896r0dc
TINVzDrWz62s4JYjs9svp+b/fTvdS+vHgSbwyj2VBB2CU5D+2e79iAZ5Knvy1aVJ
1OIHp1IBE0+Rrv6zohUdugAXadXwi5OoSb+7D6CzBPPZbcVYNqNrcHRT5ZBMBRxA
W+nJL8l6rIlHdqoTSk3exQCttnhVdKYCEZ7LlMZw8OAxQy3lgC6BNCRNzCEJFyJm
xgZMMGN6qsU1VtGQHn6pfBs+dnO3YKuNNgyv3UiiobI3uni6OLFLxkSmPvIaPjpW
Q6bD2BgUhZn2BJ3kuksTmzcaWA8f+lKoKdeOn2R2pO90P36bjWQexcJcL7kWfhtW
Gs3Ynhll1G2DxgJm69GirxoMmsxYnL3Cqj6p9R1S2CPGmxfU2uKGl4Zf10h8RLU8
9DZYJphWRHHPdWKJ5U6BjKad/QnJ626GN+qmqco2vvQ=
`protect END_PROTECTED
