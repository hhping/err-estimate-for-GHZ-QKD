`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dv8dmCVC86s8E4HkWLbiENdzPiBMiLLfLudJXMzjcxlS3Sfq1D8y7b+VQF4/KxD9
7fz1sJAb5gsCMMoC3C/6746N/4AGmx9syutbD0wSAM8dhxo/g7g3kc+wLEXOUv37
5TPawXJ6UIOoBi0d+w0mhkFNASDijKI8smm8EXP3WWIUPegiTnjPY9RolwiefQxQ
oVZ6O+tuxMO9viaYBY2o5NZsaSWNppbKjmxjzhjWaUlbdZslyADxjhZ8qA376cP4
0KqoKkbXwtWApotXqpDP7XiRh1gklGtwKuJaP6euT1/CJXBi8eDDQp0g1Rr4UvIC
39gqAvEUtMcXDKAueMxtrDtxY7cYwIwe/2fOQP60Q3EPjVrY2K2T0WOPNBTHT3fr
8Vp9r9ze23qaf9ZlDFqrRGFqz9g3G/oxcV67M4/azD3RdaX89kMv4gX+JKq9if7b
Qj+ONOZfysGE4ifImP2VrqkD8bBTNxYMPBpZ2tZEbIN3/fs6VBHgZJ/nJA7Za0Ah
gIj0WvU/NWG69+jqbe2R5LQ6sRkXJrHFr5V2SFBa2xA8IHjHv+h3r/XWUsizTOAC
`protect END_PROTECTED
