`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IKTIDqo/fpEcfvbW68YUfxXTUmIg4YKFPjxPHn/VVgqXYZ49dzXg9XUTMyZBP8n5
m6cfOrsy38550pxyxXy5+kAaZK2x6G2B0Ii/z8ypeKT3U+6yWXIXCm4osGLR+EiP
lGowdYVV7gEImNejarNCGeNNEaRhjg5Q4kF8vz76BV+nUhdt1bFqOTT72mZTpIL8
lZ+rRp7lGnJk4ij6NkF+wKEIAr7tKnhPnCXHKA0A3iS2udiBEz7bohhEbpvyPqlc
vk0NRFd9wB95vPSOc6srN7qoHgscUY3J9kQx4IPFjx07ArUMHIhlV7+6KHO8f/S+
7OOzLEAMC7QRKGYWdh+gU3BXA3Q4yiIygx62jCE/cSxRkR2pahaxQIbxCV6oFJp7
YM7zD9l9wY9rIoqJMIxRbYOZfwrg6+SLgV0Ffue679I7YBQFUctw2YFAGCJ/RheY
sTrtWpPkOeQFoQNwEN3EW/unjMGujJFsn6E4BfVtv7vI1uT2xzftEUvoH6aF9pT3
xsLyBrN9sfP8offSbwpSaHBlqu9Y09pAWgYDkc9PXC6e+NTWP/wahAxDuoy34jpn
pLuaH431a1bHdU1WIN6+uDx5p4tuN8CqKU2pGaedGvbbxpaPDZOn/UjUbBEPaeJ3
vnfQYf3c5MC/oH4hqEq7jGU0CH70AIOhUI4HHIlH+y3KwLv7mJlbF0tjFIat0uTy
yfANOkFeQWgqibO7f/CfmAIKNFyJ3BKvPHaFQlD5ByjLY4GFQWrF5YfsAOHdgtoz
0u8ZW4pyA2tJDdNtjHSzSvIofNr22v0HFzJ+owln0GfDvNpSkYjzwYQbWeIVjlCd
ctymjq8jlIWnbmp98bPlmFYqAZzp4QsBQnR8ULcYTRRpGXJFZHIW/iz+mzd/64ea
9KO9TEUc4+eJdiRUAI0XVUNdy+HPTywvFueRjHD71dgaYdZ+OrwKE4I3vFLyLZNv
oCMae7Q5kRLablhPM0xs3LVIf6vYyl7Cli5JbPLFoIqgtHE+8V3MjNuVqjIcXJMQ
uGxsQevY5EGdl9gP4R9mbBR1zC6RMes2cxOq7v+7UjWDwqN/rEqPcdB7JmP+SUWt
DMocNfzIj59p810XtIMa6vb4m3rTCrovc277qUmU/IvKdr9MXs3vjvdDN4CJC9mf
zOk/2HR+h9OV4q8sL6K9ma7pYHX5h9OYtOW6Ma744wOd7EQfH9mcLmraCVwMe2ZJ
py3ov0AsOCZ5VPfgbPbNQ2+zkVpquyHv8mrSFA1CvamaC5RFiKa8F9oZ7Nnycl8e
FBsRxQM8R0xEvvsW6WEJp7zjqhgIDAFvcXGkx3ADRPPoEcLwHdZ+RYGqpWjzbtqF
qzp6gogF8yuJ3o8MQsRmRovHJufDaVU0zuXpkaD1dyzfUZZrMPiuX1oTnNOOtiSB
3Ck9iiNMTHyi8yI2wkLbVEmEiv1ByINwLCmLIhccqG4RGb47BYqbUaoTb9L20SMc
T1sx0sVNzkdzVntMenU3MXeFHgEPe8VL2r0OyTpmK7bnpdyid6WnZ9BoVAzAXbo0
QKc49T1ElUMijNn2E2G9dCfd6kv4ozaH42z8v3FJ8TH1MqbOY8K6cb7LraTgcwo5
78gYfG0hWYusbA6DMYjWXV3EyNqU5hTrWWP1gymu8jREkWJ64VPBSuIAXSdbZdwf
FK0Oeom4Y+B3hvG2Ih30CCdWpcaZyYpZdLAsWoW10m3afRztnrgS9lKLTr2WUeB0
slD0BdNH57NEjrVWb0/aVOZvZQN+3SH79h5NrYoj3xXhMEN6uI6mZfaGLDrfYxnl
9JNa2622ZDoKLbLQxVH+1Q38CVVgzopaRQPu3iM7k2LcY4RtMUhTfxpVaDG51OUX
8vSHhvtu276VEIUg1nXromTYePCv2fcwRFL4VYK9MqJ+SXP47O7LvKgFAMesRzI8
Wn/4EPJSDW7d6X22Mw1gdC+3EzJ3TYSRhA7jccYpVSXl5sapOMTyXB0biuVBOOMX
mvNK40GezW/9hwVXzk0sezHgmYtiNzg3HdSmxnXx+TqlroowaHxsMgMVPV9O1qpN
oMD6s+a/B1iza8CmWlB/5IUUDNa0GNtFXqz2t7ogzNqs8vKDbpNAdjNVGzMdXBUJ
r24ll5vkmcebmouPty+tzQQ+v1didHcYkk60kzdSc5lIBpDe5z+yIxeIglp55Lts
5l+HigkDiHG5EOelenyrihm4XOxlzllw/RzDC9NoPeC79I8LsHyfMYofzMEVx6cm
3SZ9ZEyvFKsCEOK56kn91LoHIWEPjxSWmA493tHq+IQnrNA6gSzW9WYiQamD3R/4
/qudtGHCO8Kz6Z/deX/zgpbIPW/IH2v0Ox7MIAeMhORe75F5tbhh43UJNxsslPcf
x9uvdmcZ1vmCa/naevzeqGMrb2CZyWEBL9Y2HR0sPUnOyFrVe3N8kb/JWtdsU38n
vwIHeEumkLlWcKEzZ0MdcZUns6PJDxmMbhwTsQrhCzHO0ScMiHO6o1kzlhpWZuGI
UjCoSSrCp/7OMs8iEF/t6iD0jed4FiM4Y8lLkpYuhXtIuP5Es37wnJSnbhJjimZ8
hmshxJm02SXxgGjJAx4MQhUTt2xEj0MZIr2eXtX4wG6eoRI+rvYCgzTxeFohI0y5
STx+r5YeM1xApLv1rmSAKbskx8YV13nhqCCBkmUpUUcv6gwLlZEoWW+6HZ8HIcI/
X6upqjuG7vUZ2v4mdAq2pRvfQGSLxRGCBH1Ars8Zkv/8w+4/eG20e/+jFhiuPsC3
e5st1TdnF7AA3Xr1CmZEcBalFhz292HCnrtwLQR9p3Z+HAQfT3Urbu+TYZpji4p6
4h+0VAaRFXngapdnaoSluxD6wYJTxBCsy2gBUElduo5+J1Z071s/9Xj0y3hfJV2b
y96FUZobqya0oPWKD/DG2x5mP4Jf8it9ewNAkdjPiNHu2/E7siNY9ZMtMrlBP0ME
WNEOrDI2nDzoZFTSLnkvuyyuQhDZrhcjGnle4KQsKR5UX6ALgoReMRc6pSeNyHhl
Vnyyui9mHAyeYHwp85FdL3zPUdmmFMYNaDcc5dAh58asDaZqw3Be0YxcJpkC1Vfs
hTSJXlq6Bwi7ctflLNMZd+ZE5TlmaDkQScYP5kAO8fmzYhC7sIBI/ikxSwwxefFy
WQisz/BZgtulJfYPLu35/F6b4Wv6eX7Aqtcf+rTzs3YZozm4XhLKfoDIVM3Ojddb
FM4n3kNxONIcNHgh3y8UVCmxM7tKEzo8Xz4d4B5DUIqNOfMIg7zar4RE0J/QRNtw
qrKJP+R5q4kyh0bKw29LlUHN7+sOgMqIWYestG5Zf2W95pmiWEv9VsriJ4pst1Ln
H/shJyTjaZKCmYeSYCNQLbRxRU9Jh7bDhDFY1jOHVu6PIdWK9+jsEpbVRA/wzOST
Id1Eri3sYsx1cVFKWeFLLp4dVmPL6TTQvs2Q2nn+IZAUe7vy4csInFFG/PAR9KAb
p3k1EtR+Bp8rVd67+Xra3wfg2CozRLyNx9pnJvqE8j/jx70NQHML6Zo+EFZQKe4V
j45cNSjZ4dzwRahIXTUD7R28O7YrzgyAzcyBzWMgglEbf1+1Ezl5Dl1PW7WcOOHp
PzzyVmdrIMlGd8pxK+Mddw==
`protect END_PROTECTED
