`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D56dRk0k5OqHv3H6mkeoZOPpAMq9Cbtj4x5xWQMXRIcaxeNkB3TV4GKWASIzcrGj
jiqzsTfWEIMZdKWWEKqAOonYMV8xmx3NIElmhd9l+EEJzaSBHT4ZLMPH/x1Z2bvD
sItkbj8+cY6ZB9I1w6ODT1NKG+x8mw/g7TafP4Bta4hzSzU+VnhdvsXqTo4otisf
If6o30RaepefqgoZBLTapdMTI2wWGHitTgzff6go3WETWoW/cjbI+T06QGrqPZhH
utFbv8iF2WkaIHo7nFJr5+49NOJDT2wZ9hfENlL7Ae8+Hw0ZzFC0bs0jiZzJTExD
0Gab/o6kCF5scOOJ/wJVJ54PNFAZCVP+UH7d9iiFsVMWUGvbSlIt8qubxPP7kaHL
tRdPWAj6e2CHMvEqO8cS1D3jlFG3+kOBa6FKb7RxiD2zO9V3Rfokmso+WuYvSyzJ
KD7Z8V5DBqDO/7bW7XhY3nEf59ecxXkdrfu2kfNWcokDH1gO4YOPUV4pb0ON+ZoZ
PMKSMDu7hVzZ+D2CFmKlj1Ou+9W4aFR5YmYmD2esX3yxubBFLFnReoUgWtJAOi7B
f0niIqe/iteGi8DCEV6pJVCng4mYlF9HeEZtRToxZEH93odl5RPpbqdJ7dbjXWi9
OR7qCExRjDK7XRzEJYgOyfb1tvur5i5lHEuqIpy9rdF2nNlEhtsOqxsOpicn9RlA
`protect END_PROTECTED
