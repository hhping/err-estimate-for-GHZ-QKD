`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KWzaBJYKiPc582Z4H/guVemxJvfHejd119jccxBmlKxwABgZm//04gEAGa77vhUw
Rs5iAFxMyqkqJrAIZwPytxWLZQff+7c61o/bxgThDcJdc36XOIFNLUrtW/mLI/oX
Lw2hmmcTgNrBzPZdE/XQrZo+EkIMLzEh8nqqi9u43yXEYBkgGeS0aiXK12rWnjYU
+6O39uCH5efszOArkbl33VXW0GAU2CqBGmjdZooM5JU+qJty3Y6kVGPmnVqr0vip
QxWTdpQPtzcgg+BSMG2h+rsl2wloxBqN2G1aeIfYQcvvRjACSJX8DSMGFUcUyv41
p4tMhgSh+rsv99qHnylBIxU3pDpTe+zcdQOwEr7/DykedNPISIX+iSRSr7RQuwXi
YV6csLAuBs1hvVLO4tVn5D76VLdcB1foj861K5JFHlYezgb5pFebr64+C06aMyW8
qFCxxJoXDAJO/xwp+YKc9ksYh8w2rCwlNhkn1odBAP4YZUep7M6YkKGsHiRBsUzc
w9OkTyZLzUNvLG40QZ6T2YX2kwyN+mT2mdHNpViXQpvOCls13HSl7Z/b2/cUS6tP
OSEPkWspN039pMHXf0OavQOZlIU1Ltz18eOBuhiy9j4zV/O1ODFpiXEtyhf1ciSn
nH8feMfGHQgvB3gAydAyagrLnKOkniwVaD1hqWrtJlmgWbNlVEygKfQtJf0wpRrH
BC0hK+R4hxhZwEWxJf2L2pvFjY0ylbKX75iPIsxxUCCyy4GorOQ2o8GFWbIQBhvk
ruCCSLjBGohxN7lHQTxmhFY1v4o9R3kmxdi6eNgmSfnLEnubAvrRKOhdDR65kRi7
eJs1kepcn8jsjSPqoFANHA2MjXtLXlMUw6B7qFsRCgJSBTLfQ0r91lPFNmHTBm/T
4Amn0gdgz1ugsaGV1v+BNKfZo8lRnaj6i0CkRsD3jPqMpAXe1s+FNQ3/6Z+bBHNo
phoavcRiAD77j8G1RAZnwVDoXXkQ4iwdJoRVFVm4h3Gmua1BMkgNC06HakX9DRvC
AHBkGGLwNemwZaottxtD1eibTOgx1ZtQ1IumMHU0decfrHk3+p1NG/EuqWVTzvy1
n0Ygt2YszoLq7vEJ7JqC0u7EYODGppCIl+nXi/vNz+qqt2u2uqmzZaC1QdJ+wQJ/
C2+wF+dRHuL8Uoiv0WH62xOR2l9KsKGGsxWkk+6TYY0IPyO0/ZKyHuQmK0CGlHTL
3YkfBwk5VYofkyxUZxg6Sn0ySNgkd9rpWtxytLfrvmXcAWEvfy+RXb+vY9kphtKZ
C6m5sZ6a7epiN+PLQgyGoLhpaGw3QnhNxCqrJdI5nB6cmFHfp08WpJgDJllJdgpr
qW6vdgsUcUxdjBXTg12Oi67mHsGojdx9aMLJlyxeVd00ShRTvj/ysQmHiXq/BAvN
QzKp1dj74t/XXsPQHm2mkieBTnPq0XRfdDjE9b5bHam0YpKXIFNGY4GJa8OfEama
TkAk/hvKx8npl0e+WJsWFAwrKdWuc/ayMJx1LuSbED/E4gnb6wnxUhaWWAhncTC/
RJJ2Kcr8ACMp1xIExuafDdn7tO1D47qbQzfU8lSS1OO9pTCK9EZpNrZFQ1vq6GW5
4YBcihRcbIdHC7GllAwZ9ct2WB7T/bC++x/9eHYA9yDrVxgAZA9DZClY8P+/TtPR
YQJWenon0kdjck3uFqnpROiXXjLT1XDQyG+/QL0BrrAlV9Js4mVnABGLBCmipB62
VnRyMs5uV0PQEqEW1aoUgo9pwxJCU9QsS/GWaBBjeHfWuP5hSZr2H8RXqOWlpSDU
RfWVpVYS2S0FcxodoTJR5pnWChpQAdx9tvO3giJc/Yw2SeRXwaBHSBymAVbBfjub
aLGwn+4Uu9rnPWRWPNhB4MUKBkr1eUU7zM2xhVGRTOdHLgCgNWbrlcXD/UBeTFBQ
F00UN5xedGEuyJld7T6boydoIZDj8OLaJngFHr/JE/8oPBM39+xUnzdTBAna4yQm
hreba7zN82M+7PmuQVt/Vkse7BVj1bEzut1QKu5wEQQmjFVCoLkziMaVasgYBzQt
GrBkE6TKhzzrqWOdlhQ3iOj0FplGrR+bagUN7A8e+6aw1BO4mpB0D/GjOv7XT7fs
n05GSFVldgrLDtHEp528QVGcaQmyKa60LUumkvPF0+RjkKA86S0Cra5YrDmC4PWI
SjGP2BQEQHxM3Ji5A9YHYhYT+lBF56gwe+SrQXoG0DzfRtV1pUwHn2i1o7xXkt+h
a4mbFd4tD29xEf/Gkqz5Z3yjsoiHSTIKg/yZv+/AurOzWha4PuS9TyCaDToKdIv4
snIf5sTbJAi6vLyhWQgOpvSVXjPOxsI3HduPpTbG1I06mpUi44HoOvtzPaAs3HVw
vx+oxdY0aaSIBMxomseNBeEz56qkitNJ7ONVtSoJAz9RtcBZeJEl/1vZTdd3hIwd
hfC3UOV7odCSoA0gigIoeMot6OdXllOHa/F25MTP0mWBgXIprzlGWzsaMb3EbnwT
kxWBjJSjUGxD7ox5syIie2PDMCwuV4XUwh7nEN6FMcC//xPgJA2NC7AYW4qFWby4
2TvG7zkqXSSzIzmf+wviVTk54ireagPuAV0aD97yEpAdYhXtJJQu8hhepyiS/fgt
lSz6d+CGhbAirdBvitYPzwT9oX/q0+KNqkcHdYM0ewMg+zLu0HZAVMWbVfAJa4VW
HAaepEOy+hxjVyreG4RsZ9tXjsSG2oDgzOBlVyKIz9MkZZt+Z6F8DKvVfuBUoQdQ
Y6VnvnpVOiHbGRRirmXwhB1C0y467iVywkltVtjnzh9+k5lXrO+vRTHc4ndN7kAp
o9qBg+3xNUb876dhMF6Y+KAuigHfiluYyFTCySN1lAXMZz5u0LPzZuSZgEyy3+eN
4aR8xaF0LNElLw+54O8mlArD8H3NKDAhj8eKCcyX9MBInhhuejr3VgtypK/3IVtW
sBXGMdmyjUFKskAC9EywT7RTgDJ644DTbno+sH7z+sMks75s4aXUl/G/aVB28Gak
Y1Y2TYivf202NLwVBdxVosfnrq3IIKpv4fnVP2dYxNzz4oYlII2quqYbzrJ7JGNm
lCgGbHs4USD7SppdHY6MrcqogCvlPmIkY95n6PKNS8S2liPsT/UsRqi+GlPa4wSv
XXSaZTlIZiToFYnh4u6GwJE90MaDwXAa0WajJ+SA7L7k3mdj8W2v9DKafOXkLuAG
l43hU5d9nnqSieo8mA9PqO+7W+TAEiaJBXgkn7QryiY+Bt2bO7kZQ7aZXeLtyh6O
OBe9ism5A4qatKvDYWoGBCN8mwOYI8htVQYoFNU6imCxWfIvSIAlWPD2auJbbt3r
O+KHoT8jHG+HjXQ126YxuwEkrRH9aHT8SXL6Pr3Xz5YyY+w43BXrMExXHiTxiEOr
dMpxo05Ex18jg8vnW2YaDFHBzBTMc3YgN1+q5o64RUyOn38cO4iCnrhE9N8ZNqpS
zKEE558VFQgkejQyWSPp8YeId3uWFjH8z2OmU+IbBgji34fRITjHSU18udxZRaiW
6phHLbYjUVrAsIXAGC7xwZ+Sr2JzKh3wOPdjljOmtLUijlfqobiHsM8nYSbY4skG
mQTr134hJbQu+SaAcH94QWUayhdRTxMMZQl3oeeZwcLiD+05l6laeQ42LKTgEw3d
ea4D4WLTVLsYaLL+o37V+3NID3EVCLdRwCB9kUHmBei4w7A/YWnFgtiRAnnYSnxv
GSFCtYY6RbH7vAn3cYNMXPX1IMlLcgfliiIscW+JsKHL+bmj7hoMgB5adYiyY9tB
iw46Zba3ip/h4IzeDdje0ulYmZje3CJAJvTZWH0gAqhc1CvYXhoBtqhSuL8mcxIt
ZZTtOZVZzBYdhE+5m/rmYgMzsKeAy2SyFogLy9gg+6GDUFL0tSDZ6VtHSs3a3jSa
UL2ZsEM3kCG8gh/XeQzf3GYR+0v4u3os1I0IheYfT7fPZZK0PrsJbCez2N6+Kr/+
t5JSPcVPHCoth7XZzA0uVTV6ynUXUchNWSxHhqcBLUKgfbuORa/c124TM9ywsf0X
uDS26v9rjTvYbDLbxB+B3GRhfoU6yiZlsCWYMid9Vx/dsc/EiDGE7QIfQ6Nvmn4O
HKJVsZag2PxUjYAT4UAgyOqVgDCKBW/o5bxXBFfUjC31GrlSas7TSn342YXosHEc
Kcw+3gGICrTS2oy0XAVIVYDP0ExWYc1KGXSfnFoL5HKVmbScnJic2wBfP3h6eZas
EI/aoyDeBXenUMlGfve3JVtq/yyeLHsGF0gdvDtD6o4pvLV15SOiqn+5Wn3HLEJ/
bQie3EcnQf4FapLEiZUmfKvmWLFyJoHUB3r6rtuAPhsK//bGNhe5iIddgWmlpHMy
YTxsR6stCFIFNid8aiCUEIHHLE26EqWiz46dCOpr6bhIbl/YaVJxCRMlHXWIQYCp
5YmJDUJ48nbriLe2EAm/AFdUtu56JEgqcjD6Mlr7iy33jeCPfsYZdVdYzabvLuiN
eUqqVjtMTGSs7kxt1MFXYFNbLqY83CXYjUQjARAUsFtyldhHs77dxezBhhP8qsvq
bMDhybI54t6UiJXXfnBS7/ui9aqhRLmTN9D73Mxeuf90sjD+/i6uWyBh0mC03W1Y
XlbsICC/17rhTyLoaleCXRLzgVZiYumkI4MmydkZYNuUf8LBltfrm4hY5R9XxWZr
lPsGdPAGHlxZQhUdJBsG2oNUYqIywjRAtz1E18+0Szh2cy2u85ss+GPn5mqIQ3rE
y2F+KJk/R52sqhfBzAGOfEW1eFoKzeLO7BJk6ceyTmutNY/qN82WIaJqf8pXr+6U
kDZ+FZKOygIvWv4mZzzI5hjdiGOGsY++KZ0zhEkFc97swQonQ/YYxuZ+r3FO7ITY
TDbvxmMYWl+3hQo80A5R+tmLcHOULC/toGin6x5mfInGyjX2++3T9yppbj6TscN2
lE359AbFLb9fYIlE68MMzrtM4cu9kZCSyCojgqUy03PLx0t6oM3pxGMV+S8U84Gt
cShG0jQ8PG6VV6DUt1SFDuWzQ6vMRVP4xNNFmq7+blBRA3L08B2tskH34BJbozw8
m+dlaVMYow6j3WrrgyeGf49wpwO8PFIq2aCfd9uZMTpNoY/8JFyG76ZU6D9StyEv
R5Lj42twCpJ0+pGSZocEtR2CR0gld4JMHqF7TxKSyYsH1JFl+Y+O87ECRycrVBi2
CGDUPOsmsD/fcFv57gf8/UbuIO9yxv9IHGOr5yRcVZH2ar4Dt832gvKsL+pgFIuf
VhezekrtDh9Srxca3lrz2Rmh80VQkJIm2rMI8n97t2hx104uWzOOztrdiEDuTX9S
0rTxeine3g3pwoWgUbJWH4GsLImTgg+pMo508l+cUgN1tZFpd/c+OXoLktsnY/Bu
pROrndY78uFJOZaZeqyvDbyzQGz3suSXEN0UR2zqW0mbrD74QPphSj4cmgOG7nK4
l/U3cDkd5t8K/AIX17brXYvakDcBc8TnDy+Jjg56RGGGQIO+5mnpr+967tXgUrGR
ZJqIkc1aon/af2v2p6RmFZn5h8LJ84tZFWRWYitolXq2Y3Ac7b61M8psX9j0VU6d
0325sENSunOmmaC28kPFfo8SrFnYU/hNryxf6oJlekx858AvWTug7fweSElH6i/Y
b3bLLYtsrDI1tRA7K5B1j5g7Yda4z86PNwMcKShkfFSl2ZyMNS6/ZquTMB1OZkzM
1IX7OkU8iB7FFdaXTiJ6Xld4UYlG1Tt1At6F1ZHqvpblZX5XCC6+JOR2LbAmomFM
wbz2k4o4RAWWyOQEBJ+5NzVOAbv682K3D539UnlyLIvISdHLImBwaisU3Os8m/2Q
RQhhhuPyiFr6ep4JPG50Ex4KOyn98vaVQ5qj2NMrWBfk6i2Djm8JiSqAZoBDXjm+
b6xWy7oLBp8uC/zVjkpXQVguA4doqYn8kDfYEi6szUKTyhx3PnGskSieHIOyeGRu
oBL1ixtb5x0ZncrAVZO6Fdx/GZd8/BaXK5RylY7Mdt6ikoC4g4p8z5JkwYrv3aIw
e+5NGn3Ya3rRA9KOX5TUuSQ0rnxldgkuK5ifBGJahI7auYNB5eMeXluQPjTMOxi0
3NvWvejV7SLPpYaFPQQ7i1GVB0wz+qQZJWAjjew6RK4fgdpVfONe5sARGWpdd5Wz
WH+vL814wBM00/IDhbBvimdozU/gA434fuz1mgg9Ibgs1alhMeGeYHMhCA800lga
a8sk+wNsGPwTI/YPLoHT6cAT5xQhsG3fp89OhyIznLkBAEJxsuyUa9oHxvi3RcDI
yZsA/Iz7Ac67L99wGbFUzNN5WtlnivDvTEwxPHNa7GkoM0PyqxcM7eSEFKXZhsOp
cH6OAH3GFMNPu/y1wwl/DTrMZfZI7njlmHhrgqJrOs4YUaDgCWbzwM14uQYmrRnU
WHGto0aVG3TqRTee706V+vtOOWyLKKl/9fotkk4H+P9KrTfHPxOZwJuRWUiazZOT
6Mi5ap5GvwVyaq1Qf8ZoGNx2/RZvJlGS3t/zRiwt95+/HweeWgHPvc8NIj3gmSOY
XwyuWQrxV4rXaKyzup4TEi2mX0NxhpVhA/oLJRbimQcuH5VaNVTrNhaN8o5zE9s8
nyZMGkU/wPbjLkwSb6eBR50Nk8XjsTPjkEn4iPOOJgvLRjzdRAt9lA5H4KH2wzu+
9G5YnB+SIA7qN2V1swSAEKW5hS8FpaRJLvZcBx/CZfYwmGn8nfwhGK5rHvDj0+56
68rs57nBcOViedUJF+Nf+WR2WufYmTqkEJBxM2rhHacawnSVMW1J3vWl/7spuNDU
CyDODs71JCJ946LqJT+SehOFawFFfzkOFwJaJ5kZStPRLEBQsmGBhczYr73Awbc4
FD7y8nk1n4rc9+NPVloSfiw6fRtdpggGNfs6tYbpJOjezxfMk5dbpc/d1RDxPYzr
kOKMX7KGCK6VAxO1BJy1Px6ziplaoPipJAuz5v6Y2e9BjQ7UFnMoaYgBvqtT6bl1
sZoSSjnUyb1DvCBz6aalndJ4tHKv+tRAH3MlTEMZekDJEFgssrII9F4Jf8evWgLV
9X++irD0UEeZMtL+MztOm9UaxqBNAYljShDQdCYxnL7zTt5xOjswtj42HJTb6vTQ
9O0bpXcDjPjhusW0+fGUoGmImOQhDEgDr9N+/+RyBjiDIIvVb0TK9/3pWKoqr1Zp
kueBWZ7dTfvZ6NDjy2XhaJWVEqEj4+Jl9XtfkUmErcQ+3Yf55etWXk4y2MU7NkEm
4NN3RefZKVeN3s4y4L2sg263OiVehL5z8suUdCWAbDS6kBGnqpYdhfmmN4oXA+7w
eL2gcSjF/tpNoY+JXJj9VT6ZCzoAdRuBg99X5VjurCfxUdm+6N1xvpM4Bz9hHAH5
wcA1ndBb3dHnkbjvx0c/Aaujald66XFHsTFHgQM2JsPHytVtaGQx/vUspRNZwpeJ
fmH9e9eYrf0+K24lDc+leG1Vfo/cYUWA2gw36CrWbjvooCcaUSnn3byCM7HcxMlB
6h+zNu58FcGwKeQ56k/OOzJyaknQfCUBCmm/WnGZqUh5zrmRqchZbdOwmCqN8yaJ
KvADUkvks2GMbGBfI7OijPZO29OAHSJCbu6+KkfakT3A5Y+fcxjBYO+xPPWrLeuI
8e8ct5FZPAiu0BFRjO9j1dXXvr0ADbTzWbjaXyFg1b7ETvYVebGyxZBsQeMkiAmC
5+TFgLbYzZDSfGhvtEgpGQquAz6vNZLUpDWFXk3xsERU4BjWrMomYAh1DDJtHogJ
AubkO/5j7+lC84QbfgLClq/7+AozOaqYVWYbEE4j4+G7UPw77ZZ2guPNX/r4DCQn
z36yzCXtoPTpdAPmbq54u1ZtvxPkY+jDq/JrOc+bCq8lXS195YIPtqwVH0k656Z4
EQU9hlyc31nZgT5vI6fCe/JcIP1T8VNhdZIzShSdBdisx9aiKCXXTC2iX6o0alYc
EXTNMsqSOCnRyQd387LUg6WDJBxxbWzc8QlXgAbbK58ZQoufeZ6VC70yx3f3/y5V
ZNHMy2eWPMohENMQkqRn4kmTYxSnpSrMuusUfpdZXWBDbM/+cKePgz5G3Io59/IL
04SYMOFU8YpFuw5PKs8NX17ArjqX2YOVpOb8WMoR8oF8yvTtCrmVCWROBMQ4c3T9
pB/WcCO7TWLquQyTvJhnP8v9o/FElh4arXp6HfIunC20vlqvgDRQwK530DEbertn
5kDaa9TtAZ4gBJygp+TmH5MXCxtEdhzDQMN/bt0R1ZFYWtGiWlbgL1n2tp619+AF
kYkIG7s0jigSOw9BQ0jrfqSvAkXobamikW7U5oy3OhB/xRtzxfGuf+plLmPN1WbY
qN0Lm/yDBSF61tjaMkU8FKNb6GwUNrDf0hnKrg5OpnDx5V5n+DR93OXpS8UNexEh
qcV7mcXzBD8vCjImoYONcH6uEL90XpdQbIXTVSm5sZAmNp6d0F1OHwQ8OwKdfdn9
Us9d6DsKm9vF6COHUECp8qZr/acDZQLfns4t4rw7wRwTnTgA+274DN2e4wVtU6f2
bjZL+0g+0Af7H6FDjRArEp/TK4VL1ueUxfdFSL+pmRRf+PIuNwkPbwMU0h6oihOi
JQPM7H2BvQk8eQMswgYccheJjPCGO+5TlPd6uyCvIqmTu3JaJxJi27KiamF1srhZ
v01UKMVQ3v9VkYKdWF+dT4cGC0bJY0ewS0+ycI4CPfP9gXstSrJWnYdMnUxgj+8A
f211mot0D8XzsPBswUwbj3SM5+tHDbiAurafDkyJhcFaYjKgBCBXLS/JjtYHI2Lg
dgUddTrC679RskTVr1G3j5KoJJ09n0t2oR55C90l2uaptgkfAmEcNnRUCFfF+4IT
3PvIXSYbPy6+0IvG46ePzC1PFOrRp2q6n07IEqt4mqOU2Kqp80A0cEhrW405OyAw
NZxkuzoNmWc+q0aHuQh6Ojs4tzogkevj17x+HAXoxZD5xhJWAa4EpCDmkVjJpQId
h4vzMuCZohVFiNtw2RuMpLgzNRGEg07YWOJNGf9SG/Klbw4bJtKM4S/35Tc838O8
P5lm9BrcIoqSumHdCW6RQyGvDXQvfnLRUybUmm5JtvDFs3d4GKFhsGxwqWX9EWn0
kqn75vDbAbMcGMkEXwKet1EvIPc4Qj86LI0kymhOszKhdjpGtr2CCRTQzUeALjVb
qTTQU2wboijSQPRF47GyJxjd6kb11nOf5ndQuZETkXZ5kYzwboSV96/g8ByvLOxd
UVx8NFCuVRmqAbApx9rSt5+UsFyh66X7UwFx43JP/x78NUV4R99XigKxG3Mnjmng
cVFGseT6bnwYCSRI2aXIKltHOR5zHN2x1Q3NgOeNRHL1aBVCnrCHPMT8O02+PMGt
NjDWzRF42JqXHI9bldBqj6yBCQh6VtSSIEk6GcJn805VA57QSAwfUBiC5WvJwIC2
khZv6jnnKBbtZjAzCIqCODf6Fc/CMLdufme6sjI2ozTb+Z31EGfrDDC+iHqORcGt
BKRQqkEMNrlKF/cwbG0JYtaXJrITJzvyeR2BT4nrqjyBEzT30ndNIRhITyOcqLIq
JX4c4cSYh0dpNgLgyo8hsJ9C6K2c/oCsAvVP/wzIfaHkZsYtISeZDOSfkPUnOkt4
RwhhmYv7T9COtPwzA6tcOvs2CYx06wg8J8FB3v/62iqFYroi3Mp1X+alsiHo1Zh5
7/W6gH6CKQekfDJTHTLoVhVEeefLLwrnFuFFmcyAC4PrN33okxz7jJGR1JAkinzw
Mac/LHf5EMZMx7RsWS6mkX53ioIHmQSeFhTI2FMcXJ2BSzTadxbtiyDe/mZx5wy1
ZNWU16nh9oZQ6Dh5uQhyv+Scd+ol8x78EL86cmPPe8GkX79PhezZvdMrReEmTZYF
bmONB7TywjM2iBJc9JQONP/YUdBicarefqi1umZjYDd+r36m9LrMMWl1yN5eWCzo
iJqxQevzjO2N83r/0+cOBwh5HOXngCI3nSh3EkELFAs3sR5g5fCwSanB2UO6vZKi
RKn/nEl77cZU8+DcHxHVnHBF93IY+lLAgYTUesGasH2LPu7U5Eh1VPD+GPnRUonz
uG06b0qkWHljaTQvKmst5tA3SgEELRhiMtEOJJ3d5MUvq0djP3+8QgG3EHwhoa+W
/aN3tvN6DsXDPvB9NMwhBuC5rxZHLNM0V4bPZegw/goqdUyfIF420AhL2k2SNjYv
EOhQvFwmjtI6kOqI6Ig6QiUoezsJ2sw/0i9gSbpoudbUzlRqHzfqtcO//S8/uKHr
pE/eOkur80SOHW2FCCO50B8ynXxnDVPH+jB9kgpei8fI35eXO5uurDXMdOXvLXZm
7l6AejKGrgl8h6/jv7xpQXZtTY9y5/FT5zYKX2zPfG3e3zqxlZ3tA1cCNWLO9r0T
Nbcf6h2G3M8DyZs1s/wUlzx0ron0ks4iJiR0ekaFQ2Rlf2GDhkX21r9dfIAnlXDp
VMhIrqoGX01GGL4g6aKBTe81Q527TkZ5wJBQg+ZdymtNewmV20JC1e+45UlWVKX6
pwo3Tyg5W3YPawQJWbk9/knc/51Hncp2zUVOxnLHwbp4trV1g3qwPK5Z54iNMid0
ew3cMk3+8cUNGh/3bhABgesUqSxeTEMZ8tOGT4Q08TqTW536h23NICQ3yYJHg334
1WnKC0hwJqVJgqRiCLklhqmdwCnIoEnPGIfGi7CbAvRUeEtCgzheVQBsyICs32Rw
H/x6rQS5kES9BA6AaDM9e52mslUOSdvY3kxiAz+OX3sxVOIODYZsSa2kksisSt1Y
y5ce+G0x37sE7VBDyocOZQEg+TQX8wxzO6CVUPwkcORydKO5DX1X+LXVf2C+jEfW
dodNB/MiPWsJX3eAPZIgBYUDhJ2dZY1vBXcAv0LdWg8prXqTjMGO51chs3MJKfmj
J5nLU02bTj3cBTPuhqqL4XmQHrTuKsuQRQAN4X5TZO+LbijaTq7qfXLE8PTTv9iQ
l/eQh9CL8vNVwoq2y9fJfqjShmsbJe8vvnuNaTa5WJApQpSXVK08q8xuesJto5x7
CcdT+ld5wjxV+8JSA7HoHbwqMsjDANpqpJHz0sjYTVP6LulsJfD1ZPpyb+MODMAL
NLbWfs9eHOST+BEp+WxJp50Q7uOMAeHNDo393/Jq3wWnGAWcO6TTdUTFDqbA8bzt
moBtmJ6fMn2Z/8bqt0WdMBMrz4RttxjlcnZWDvhiQyX82yTUHWiYCI7KrpKEaAAC
dcTBkrugcwk7oUIQXuqMF3DjRAZMKmHcMCOr8qN2hgIrjRRFsEUOeL/neTDRmEGl
K9/93UmngJA/X4tNLHe0e26UvpiT9JZ0Th0EIe6VN/OjyVhS1Jcv4kN3wB2p6c0B
5sfSqzbEfBrGv8Nkljhqzu90i3vwU3EeLUZQ/WxB44ftpSej8UvmzAsDkaPHZn/d
L0Nj8dMEJWBwCgJgLOorXAQrX6P032r7zOPiOiyP2W4mHuhBFMqyNwxOnq+OerGn
DpgTmdSrEjqkPlQPZruHDfShWtKTSoqSJZvcWveDMtFCk6eZC1xPT/wUD4SLizY0
xWo2KV/ubfGQh69oD3zHM1KTd3YXXWoF1iNQE+miLxRl9SAl6WIj68zaUxpLToy6
tlVTRCJWqHAPCS87ncGhPUM0Cl+M6P9yAqQl8S/xzKvkAiJTDh2YWR2ufWLOoEMp
jawDxBNh7fHrq/DE2R4NGrqDWbSSqeI4SU0pKTqgyvv4SMqlGArsrQfbnlwJtG11
V//YNjviYQj2YFnva8nc7ZokoFs2j9mrdDD6cnJ9s3/hzgckwuixBU4WwFnOYK+s
fDw80gCTNGdSdLFK4kEC8QRPC1t4M8x3DIgt8CKVvjUYstKqbCNyn4+GvlMeNAMu
GNddwKcgEC42JGSvfAc9smcknnlFZcRgcp4GBzXx6KwKzGOnPd080y3C/Fgbb3rM
lhuqK1lQOdL3gknN1IdpWaN/sw8+m1mSdTn9ldaBRrLNjgVRp4Y2JJMEs7t2kOTz
vhosL8C0QpDLkCnGbONNB2KM8iVcoPbJ4v3c/oxCKCpR9kx7DLXkS6C2On6lqRQP
wZho9jcevyfDxY58MsPD/Yb6JGo1ziBJHM7vKXY4o2fcgSDGZGkRxyZkCXbcs+B6
rCxCmh2xGq20rWaWN2yUsMaS6HmVYMYFS6IyOMcTzv1yBK4nPFaqs8iWvoBzDaAb
eduEaI3svvHiWbtKbK8sazmB4UcYxOCubB0NooV0cvFgtCLY7rG8VvUJwr9ppct3
DQ6drLc+1/TwyAQThiIraBX82Xkf1f4QNN7Esur0ly194QBO7vuKewmjx3Xqhgnk
SzQGNu9LDGggjjlwcn1dRsppQeONvnsoq+/wpkafIbdvRBdOMFTcuxGKMKoGfrwQ
fuMNq6HoHGbqLnxHWE41bj+eHkZLDK/rL/9aQIBx28ZDfdbdzDkLX3cNxJAyhuCa
9MuBVxdm7GhzRjUPsWVqyBc+TRjprx+d33mwNdCJMQvzleuwi6HocOmLnTdEZ644
W5el8ArStcIJoVPwT5KFDZ9VjzajgThwWqmoVcXwNI8FhZPfL/mUf+kUAXRO/8BQ
c81pXGc07M1FhDsuGA5Sd5uc+4OWZNJlHefWzziSWQnhlrgwnZh8O9xwReVAnNyY
DOVK99fizMnKAROEiXOROID44vJbAOTm8rUb+a27ZPzTKG4pVjDX7rFU6dPKQQoe
fJT7bA8KhuosY1dLGsotGPnNohmP+Pm6/9mFrZm/KYP/B0vZPAtXjd4ElEkrFZ29
5ydjr9tDv0iWdLGsXzYz9gwivkRorr/+kPvwj+y/kD+ycwlewGRSdwmHIiP5/465
UudZZcGCY5nRifQJRlgeLHMeKAQCo3uaggwSo/4uTN3cz1Dh9a2Jb95WefGDtDYv
Vb+b3MS/iPqsdsPP3jtFLOw7KXyC2f3jELmrvE/mVJMFhlGXjg6cJM43e9oOMp9G
DrqRDhu8txjxgKQoCpDWYrR8tYsGLWonN4jSGIxe2hsWM25k5dI4y3OgJcQ2aHI4
fcL378KxKV3RP1hZMHdqNyDJmp5xXF47V2DeA6tWctGx9s2dETft+PtIF6GUDnc7
Oyq/BMJrOtLQnCNCz+UDfZx4RQKx63RbSRB7awJvg7GrJr5C7Eoa7hHBlxNTairc
+W4fORbs1q6XWdLTPNABbSwLjmIN9IgmQwGwitKakjx/Uc++dEv/VeHfEXF2lRBq
rvcCPjTWuPAXFiGBH7apR5360LJdhpH1mP6tHgaZxPQY7MSRCBFMYF/d0fYzUGGl
tP3SMvaRaFRjwMGW+9tU2ubCpprdvIDDDgHs61ImPrkb3g1PukvOVZSl0a6mQZ5/
59YB3yYyLCI2oSghgYOJqzR73FlDsVM7FlCpp6jnnZE07gr8ZPIcnNHzjVx/a81W
k74ADe0T5j6OifE1bMSSp13oeGdGROtDozBnBAII5tfTDyWPTEaAaNhsK9m51DLP
fXRruST0AeAaZrJOQjySDlKopWayfFzFXx2S4EdDuqtY+LpQ4SD/8awodCdaEIPG
mgk0nl8aDFNAULAxiIeU6ovnD3a2EyHGKUVEWktvkmQDgVbPlLdpn8De+M3HCPJ9
JwaSTkAkFRTARL1FIDw1WObTBv4+2nZ7QFZ3iLsQcI1iduc+ogkfVqmyWQYEAbmX
2ThRPDsixWdpWQAPHRKTUM92UhGeLc5ofzbP8Ay0toM9VkOZZtJf5O+4PL4AP5Yy
Ps50hV6+Eb5klQ79XKTq+qm5eeTvD/KYzjpbTpNeJY6YL/Jizr0oyx1aTvDxym2p
Ia15DtCZD43a3A9uJwCtfGcLqh3D1KdNzwejpUN48yoBOL5Y3GeVRSkD29HzzaeL
GSFsOUe7VrGln3ZgLdu594rkd1NARNBWTva3zTcoCq+sXd5Ms3cnqWD1BRc+wrr0
VW+wetZJIwWPVeDCUKb4653HR6wrcC1kCpyaLkpNd/eVuzscEv3GnmS8R5w7WMVi
BdfvBhLrn07PBxiP2KcV2QYyGPwVqK7WcTFm0+vXDBvPEX0KOy/3PNjVOBnqCzpR
fPztjJy4P2AT4V29OBXwyQjOfXd3/MfLUuAgtdAs1jWKBI/ikeMq5uQKvUc2adhf
VgsR8Qmh/uDB660xyUqqjS6e+Wwx7SyiAjFIUIE+3drVpkLkgXRn8YeUXuBC3JoR
Be1l29q9hJonEOn2NWKyfDy2YKZE9EE9o+6mrpWAqW1Fqh09vWxEMXGOr3wCRCMt
HA8N6jMOeSOo9JKO5s1u0LhpTGLLj3kDjXuAvEu2bJEk48kpNURUvgfxLIWwdoUy
lGLWP1krl6T1RteDK1Z9Gi5i8SkXL7dS5P4t8Z8dx9JjYB4SE+ZoW/rOXbA6aN58
NQO6Z2VBA+zPsxBCFSHrPSnDl3T2+ewMfPVuizqJxdtX2l79I/BcsNuciSlQbihu
lp8UNQHAZKRlbF75c2zFl+HAVt3TxpWCXzPBYUDX/Yc09EGh4W3yveEm0skUkhNh
7EXJfcPpoTwVFvoMlIgl6JdoBC0GgSTjNm5S+RzyY80nCnANLz0J1e21NJy8iCqH
CbPCrib21yQ8oX1nGKQLY/HsppM0kpd8o0lANKBDH+jKlinV+IfCS3ArjfKdgx0v
KFHh67upIVRREQ+R5c1Is81wl5V9eWFaZrvlyqcVV8FMrm1/d8+bN0DTRaniIuBu
jMilmqF9zjHcakSoxlai9jzGGc54O8SZawPP/eu3LSwlJA0rusCVwDoLo1eQj8Rc
TwDWJQbpzXcSs2xkd1MAlRL3FgaaO93po05tT0AB+wqoww8US9m7AD9QRiB3rhGQ
B7vHkgTcPJiZ2rHuAe8ydFKA/o3DGLVrwEfi8j4cVXz7sY+du97uP2sISlluI0S7
jIQnmQq1kKymxbC/3L+MMaMyLy5mbnNtY0bUCd/MpmXs3qy8m1J9IvLdvTDIldug
cQmiJ7ch2FugeKiIO6XaB6O6Dqvz5My6xDWkeoS/g6NndPlPzLx8qRmbpxD0gpdi
bmKgvW/v3VBeyBy9emjXq5WvT57765Hg8ZFkWZ1ZwpFwKBAomJ0jWPv7JrQvsO7o
zZoQwowO/5t7Zds6vV6+qSetLhITHRCDfb2zNGxGBBsUzUHf2gLfI5jGsPInmLeq
BwVyxdpK+6Yc+VJoETbXcGFZ5MMy7HmqzMSSTkI+l0PaQw0c+tLvcKUiscuRvKOT
AZXertVSEjB80+HUKBz5FR210RD80azsMTL1KBF6Hveifdvc5Pl+YHmgDASnYNYI
ujsUcd7zgBwUPM3EG0lNoVTEq0WeDOQM5yFmqnP8sS5WANqXTQZXAt/GOgq6O2AV
oocWfW9nCvC4xbFsROCOPOSY/VG4nElmnPk6gwg5m1dHAjQd1Bt/RWcRCOBBaQSu
QM3idVon0TLMkkqbF04bTfdTiBWKazchh0o8Pz2hFhcZTfOwe8RB9EYSxl48Jt0R
TGQw3A8SD+6pOcPdBy+9rzUGSEZI1Kdsc8vdi0XAd1XaG4+JRajaS4FZ08hXxO4z
+8ZuNKeUne4kXYJi9bMfDjKKvsBnAcUHZZmKHuez2IGWZPu7Nu1v1MKPc/BFbIf/
ek4edKSOr3LnuDlY62fGFru6GW4OrbvfW6ibfopMZl1Stt5mNkTUGoepvrM01vkq
doap3jvMhSySlLy7W5uW19Q/rEPgtU9ORwDDmT86HfJ+89hDI3DJ0s+rQp+kdDVk
iZEud7MFgZs9zBn4izc6krKmUwr7lWP4zEMgUG6NL4aAwiOXy8X/HBG1fxH/6ZFC
8I2xb+WmWOaT+vzDrdQRvOjOXUDykjn2Zum0CtK19YxJClsccNFjIFYDp6SxRTCv
GRpof58w2ViogE/u6JZiSkzYwgoyX8H9oOktf1Q4XHn34Kqt/mw2Zba336dzyhR4
6PqVlNxlw6o2X/C0NGQbFHulSlQouB9dG9VmuRr0lCgVDOAxQ/YcaY+XBXAqKUMQ
ktysd/sMm6IiK1h33JpbOCcyjt69mmGocNx+Topp0Fzn+klSueQQKjk3/aC+HWkK
4/NABYU22ZBFvPsJOksVhQbMkstaD6oN1ZAbAX4bHDJk+OpDqMKwbl/aM4/kLfwQ
Uufyjj1hCG6TKeGU8FB3XmcYE6X6lRi47cRbwm79rJH8LaMfd9e8f1fj3q6XAGLt
F+fgTG3wElA/7UJ7d5YtnJUwGGzcX92N0z0V1p4ozjf4I20Lvxp9h0H5H/XczVNs
PYocMc2YJ2X8tmVZc10H50zl77e4hQjdKh/Df/WCLWMSqAUVXZ6e7ih6qDJ2vXOH
YPPiIUoRO8iPajf9f4u/TPg8BikhzmPKFJiVEvraFZHdETPP6eDxb9sRENb1FT6E
pNIG+7uvJENIEXpYYVVCuD1YutzaIinBhrgLqAJNJG5BIAONhmMYbw+sKlytkED+
J0VXJ1/dXU2yRIQditIfcir6gwdRkNr57waxZbezgg2u1/uX/2QQdSvtmo9RVYhu
80YGaj9bvQrEVfkdQE8nMCaOQ3AI/0Yav0Hif2jI2M6hUiORVY+G+Ps2fWFJbpa4
rIWB1Z6G5dfsJ5t+aFcUJyhFQ1zNGfRIAVMguy1I5hADcD+rDoPWuyvMS69mU4sK
Gvqhp+AkSOxiouA0zzPN8hODMy4DsbaB4hY8CnUpyS2Ad0hVO1tdCxJxd9EXjX8B
thtEVlQNrn7Ij3KA1Tj9jCuhU2ryvGLzDPL1Ipv9zUENmjx/hVs4KWk3KbuAcUkL
mhK1idbyyBVCkMj2v3Jb8fWzHMjVk2FARPVRSM9kQ1ARQ/s04HPlyNsFSzUHAAFV
j++Zn+PA2DowdqK2Dew4K2EZZsOMb71v4f6EmrdiE6ZuJzFSsHzl5SRoZU/9RnyG
IJNaGvezTRXhOkUPzcqvU6hxI0DuYo0Mi+mEJKC+Cg1NieuipXGik1zPuGXxjsPO
J1BR9WgfYSdo+5ETbZzsyq8jb/G0DwmK0rsmW49a+uPAKynPo9Tl1bG//FmWYx3O
QxaTqiJFkXUTdOTnNIn6H0xhqXBxyPtRdH1yuepa3RsGsr7Wl9VQXjQK6CuzsppC
dGoAYxbkUJf3RyFBE5SqLPueGOlasvV6iuArFrQiX4boDNmt4aCpI+/D7UZtal3l
Jg/tQK8jq+h+HIBDSqhOx/VttD0nmxlG3vQT+SnuTZQyXeOre0DEzjRISmxm/lbe
I6Cv2SDJOOwAkIvjyNGsY8OX8MnpNr2Yrdgc9tC27xdh7DZ1wgEtkR7W2p18u+D6
jHum0cJt8KjsYi1UoGS+y3JMlcevTmjn/hLvlwEDV3gyfp2fxMxM/mAZEmEfenA+
tuWCBlfZoIYybtwAPAF3u0BTdvuytgWJ8aAEzvEOSD7V0IT5tzMP9selhvUmimr8
J55JOrvePKJPzWAjsucfIYLntwFa9Xo6IfKhCmX0XHKd7WJNJurS35x2HUqLfLdM
HElQhehMYyLuSokxZUSg1yU+o+cDFjKnMj9YiZFXgZfGXnLof0uO5bL9yvCkpzGX
tbIO2bnPhZRRgZYdlrxrdHiy1f7IyYU+cLC/4BOoVLxJc0fpcSGvKwiu1h1Sliql
CYhcEoRQTF8tN1NH1ljLTrfTdRMdtjknP88JmgGMnLDtRbQeaBUSFWy2ebT4P+Ls
ofGODPiY8cnlCOZcGj6mK9bCNK6V2f/hvacLbXK2znf3QpbhMgWNm/Fpm/1KprcR
mhs5RZAv2tRcqHRJLD0Tpu+2YXNOWs86O0uuXzqa/3HTYe/bx5yIDEULlpdEOuF9
32Gj69ogCbmwQNSorj8VBYAY5SCxTWpxDME7oUMW8lHMwhe2fQV9QfBOs7dJWP6I
6/ZCl8YQXHyPxNJV9gc4f6sczaV/BcKKS1ifXwWjsqKkisiQKS452HeZ/wyOve9L
y57dkDSn5VqZfWhGkLIRWB81F/ui5jGwWwWJYPqrzdQC32N/kZ1faiDFcT4ML/X6
/lfCnBGovrlyYw+g1jVfH39It2QMI5FECX3ZzrE1SCQYQ5HkV91L0QHdHC2tJBK7
R+OeGNZ2EZ6VGyShHRK25abpVp7PKEbrlONYpIMWxCdqcCoMDZew6Z94AMG5n8HX
na8c5wr7lQSJCJstE6X39uy5NifljfPighRLY9mccxqWNC0PQ/3bTyLE6weS/lMI
l2wxfi+6ZE6ZmvAO6feJG75Lv9lEex3xFG11UrJdQzMv46ubQKW5EAfZ0nyxYyVq
AXMgmn+QtCLR5o6e/vtik9xUshf1ENFyoXNZbdAY5TVH0oL9AKF7vk2Gc1hBCkD9
DR+7Hc5fu4+j7JFMMOItAa4gnzr9rFZolP/bnjZyhlcZigrZCGYT7kx0q4ncmRJb
jQOJTZk1hBkDvlQluwkSB7sCPabxvvoovi3yop/bLbiy5e57sDmcXe1ZiayuyRDB
XdvFlJpKAXiTOWS8MtCejw0Qk5PCaeuV7g20Ox53KbokXC8f+62vfY9q7HfQcUvn
kB2zzwYT2P8rOvw8TrtFzBi8S+IdIPoEHCxQE8RKjiAjY3WS59hVLAoeQFKhbqYF
ZE2RpyxsnHmfJ6fgIHHT271gj+KfvZ5JrHaOFvb3B99CRbvQ7+vwffuFq9mTGRxh
IG7jhB4QBm8YGAyk/C04GpV3JMMEdmMY7zxX2DderiYLr6fbR9rqJ1dCGUUk7LjY
zonRGDdqnMGurttkx0n/D8bqT3oSKcTFFtaynxwKn+Fn26x/NLOBosgusgT953Bc
yoV2FcJJ+OzEkEFSEcyWFW0ZVB1HuV9DopR0SUSN0vBxuzzVuFAR60gcy5AG+K/V
nFwcdhP/4GDzOHkclGmyFwQ79Aas94NitTIZibP7udG4HpmUhf8bHfWwTuPmpI3D
IWWHEzqLrnv8I7Lhzwt3sRxqO0wU5E2xoYTiR7R0QJ08EwTaccHI7mA42YoobaJn
NFXbtK0E1/omTrQpiR5VfPQ3xKC1MwFHXehRPbvmxK1DD+FKj6rqHYEsiSL594XP
Og/UsEMPUUO0RA6uXSy5mfoB+OdyjbMbbzmD0zyFmzctkVpvYPi2fzux8PhvWKxZ
W9kP1i1L1MmtTwCBI3jtFUfK63Fb+g7VuLBrdHuEPSG48a0PXRkcunQYJG6T5vV4
2pzZAlEKPl/rPGd8RAj459yIFGw39tid7nI+74y/NOgwwdHwgQrVgENbwdxqHTHN
LxEWyAHPNmvkYAh3eGA+f3mYZaogjUllyWUzgi0hqke6ZL6UeDHE1iqZdPwCgsP7
pE/ysF6F29rwNv0dBC6O4GAWJ4Y0SkAIhfq7Wn1QekPWpQ9GG9cZpMjtrGkWxUHy
Zp+d1YaYf9JQrF6yB6Vaj6Kv1S7yAnooHkVzxcQYeYwm1zGONpQ2ebBVbsNIrYtA
F0LYuEDKolaN0GjB1RpQYhXox+7o5YL03W+86JrfzbSuiS5sWGbHY37e5LYtJHys
HnAy9tABYFE3Cf0yWRukf1cjiq93WZp1c10KgCy1LVz/LRPuvuDCS/NH7PB1oBdm
7TIzqFlNwlUP2JOrBKaOODKm0hnmoch0k89NNQ5VpVFWIf0TZBmxHuRRqMH6EjaJ
526MkERS6+NrHengBpSbb9ZbNhHcwj4WRFHqijqXLEMJfi9ekEGWaJPDTI7Vs5Ys
2vZuUsQkOSV+krBQZQiLqSIRN24jSj/UyQ6LUT2nGrQS6HwcRp5KiEJ3IDuglSjz
6ZmbeZXci6VoJo4e1NuyxSeZQJoEMGzviv5v2FMTSmgrtO6asR71iYx14i86kMcw
51OW3zO8vu/f6qQoRcrimwjWeANkjemHHc7a/WI03PeF12MHxgdaN2WXa5GKGuKK
aTqTuUtxe5yz9VyMTZab95/A6hSwHBfBr4YhQrZZ6Xmg/IRK/I9E5i1NGVJ3w5oe
qPPsg+ZOc64Y0Q9JbNfHEJNqwny13vdXtAZiMGFDtnCe35rJkB3gg3UQ58wb3bKe
t24QrXerDIOWFfBOC4cXR/x5tsuD7v91AFA4pP6lKcyFdJ2ZhpSw+V8KOceY8l6k
g8quyoaLQSJkYWoqL8L+DYoufjJwz3o2W8WoyKF4XSjwPcQNU2tPmjNxjiMA/2Kl
qCxFXVpdALK78Q3wgahm0d2DyvQpQdlV1BgNkorbWyfcTe2RHbufTODEChjVWS80
oA/WHGJxO29981AihI6B1uOnx5VqVW18A0xVbTTUy2to6S52R2JxVlcgpT6t8N5G
bnq55j3HS4tqhj3iJ+1AH0p7QGw1UmuUVnNj9iqdbNbToyr42/vDLlxTXrBK/UM0
XrK+yixF0POvO94QvGkmJFFFcVOBGFov59iifhTD/nWuL3v/arR2+gQxZ7L5GuGB
JaAiEH8KmZdIgLndJucMROLhwt1ZXCgBQ3dPnd8ZQuxTYyTbOTPNDzo9g0ewsBNG
FNRn5f/7FwINbYrgQ6k1zvMncl6k7edcOlaNotrNWzvzOz5dAjaJEaUfGo20ikkK
rXvJzIIr0TquDr0T2etunYFlLZdiVxlph/Bd6OVd/4yk2H7kd6VVDVcUUzTxVhX2
oH1K8YWb6oZmB0XNKueb98FOr7q9ZsyKVSullfQbI+aCPa5LpItZoP32CHcoQfpH
ksKn/BFDVyoHCnd59hEjeZ1h2v3r3q43ZRczPvSQpWqPMWU42Kj2UrgoXCu6FLIp
GbbwbT0kGohVqH4dxtC1Oq42Cts/wPdSYJ29Dk1gBQZQw9Gucz85xzJKamOT3QLy
Jw8e6ocZVSjhOzYKL2C/PMaB/zxKrvr1j4mQJ/gZ8yvsjuSa93gsrJmOD/00nfiL
7Tzu9qSurtVGm2latvXp3QT6yaHwLI/5y90V9Ekirs8M5seJXFoj/Npuj53wfWap
+pIK642IHCmaXyqIoeqLTwmJ46rX9OEaV8uOCdzyQ7sxESfv9zklxKVcQWR40BNf
+Ysd9tjzXGux5RVVSMKQPQd01TGW16VRgna21twF+WFv/EYYNIk/QA5uKejFYOB8
Cal4bgoTP6g3EuJv9PKOgqSxN9RrOzQ6WtQaS15weN0DUgWGNz9zym+NGvz9KLGT
9V8UVHBVWgMyGU5Vf6qSdZ9OljZAlc94RiA71xGh257yBBfnbk2cSRbEdK4+ocR3
DYhKZInv/4/CCqVWOTyTVkC2idsot9hIOCGXRnrVHHLZ8e2HM6Vz2SxValW/0XOI
mWGdZSEs+md/3Sd2fHRRmktZUBuo1Wp7FvpUKQhmJla9+0Wk69YfgBQAzEdQipEL
5fMb3M4+oh0eBACSRQF6SKtsFGreOW+ipMd4JZgk71Nm6BCGymr+tTCL/hd3smYY
n/XMi/IFNK3IKynNFu94sv12Dh0r+0SpQ21U5vIBFdzNdLcyHHHuvzhWALTmN4wI
3JFRAzy2e+88raANPTobJlXdk38CbnSAUndywG0KZRNpfR1jWjBnovQ+KJzqC2Ic
w67XR5XWdE66VTmSrbs+fZD5ymsp1YmH2lagI3xAD8gS97K92P0CXX4XPHaRhixD
CCr/WXI9w2mEOshfBr1Eoab8RG/GDSXLGU8tuxp0tB6J9Egn/2XxNzJSGvGj03LY
EMVtve05rAcT6wTioEwmDHHBW4q9R53/HoJYvzMnL/dHbxS4ntSzZ0MwH13yDAvo
F4uA6yFdQRJ2I79f+7QYVj4JgWoRz0QBLehWD5K4NcTlHcTj2W/DgK+RA1uYrRbD
a+XoSzzlNOYK9f+Q1AQuRCnzoSaI/IQRhIBkuxNmFcd9/sr3l6aR/Llvasoj1PoW
s8ubOFQ923yz8sTjurCJqc6M/fqCud6oNTumbRChTySMW5R8N7dB8jSrIWuwI4Yo
eAiimZTDvDi1Uq3xLvjHCVr0UrFkyZmidhHt8uiMKwx9ZYTIJWnM7lS3DpBAdKrk
Y8W1GDoZu8pVTmYE+Lrw0m5Q+NkhaJD4zbg/uYY48weYCOCWNMYcUmafEhgbChzD
gdzLq6Yo39hi3ubp8S4OP32Yg+GIxt4rCLUdCOBbc7bPqBWNTx2wlS48bqR8oSlq
34UaFJJUoDJJeuS6+AFIKWQ5vMByee4AUZgmR+QHOjJVWYBe2XivC02PQvk1IYJN
CushbV12Q7xI9Yfq3jloKvS94+d+VyBawDXtoLbJKb/BlbGKHQwQCB6YMtIWOI3Z
ZZxJsDNIdbPGDlOywrpMWgQGWvWFOVmBcaPGUbgp4eHv1N7xAp07yhxPAULn9uOV
F5Ti8h/ZWjNCYjlaXvLf9fqojsg1x691kc4VjkdnO2qyMhk2BQ5Aqywg7wQ4d8sD
4PZv8KSzk4+9AE8pxVgkuHjzUoUA2FvNLqQ+Fjjwu6io9ddrpugBbcbqsyvU6rGh
e8Yb728+qMfHr3VP+2DCoIy9uc3lYgWkG0G3HgnmE8OKelPkVyg06frfG9HV77r8
vaDfeDrEAeIFflbxGyYGyl45rudGUJc1v7imFoPUj0U2T5C7c9JLFb7eGerS4qrQ
EfclZIN6gTVy451naiInrNwlhnSB091k3CzQeBDqcaT9jCQWWqiZmcDZgbjmxwyl
124vLpfZkp84YRf5ozJFZMJkn79D7AmOwlwg6fz5n1SbhWxBJwGjdEng7ABy4OH3
GDH4b4OOmeyzSz4/6OcMMzfXHiB19SioOvpAhFFwcgzNVSOZhVIcRFAjT3g92kLG
bB2ZjKw/xt4SAha/lLRCPkrtd3ZwY691hKrx735mY/m2GWIOhRQH+TGeTiujkpms
XTpJxUYVbxlRvnDObn+vMX0/R+hQYZ6pxd9e7pXOx3sHLH/VLVix48BbGN5VxHgU
P/yK0ZYXrTu3LQ/5X5VQ+hfNQ91PDrUVTRgXvDVqXCUkOwdyqbd8G8n3F1m43Fgs
8pq/90dAvTnES20DJaUBmJag0ouKMo5qkq2dUdE2ZaSF7ODYEPUtwMl524ltfIK6
wfQM2VfOIAMDcYmvl+DW/7HmOj8mP+o3MVhStgbz2PRQFNWu6h+jJUVXeR1CpJln
9i40CkXNYPb0LDkQeizmeoSr1qG+BVqOpW78FCkxsC2lPz4xPAu/2Kii9Ff36x7n
ZP7Hoj+Q2fw/fAWK56cxMFKQ+PUIvsSsWqFRT6aHE/8tkKiXL570Wd3R4UEmD0Wy
dcshrZFWoZ6N2tXS8TM75mzxC3f+V7ycH114gkNK1wGXQCPS6XDrAizgx6STwMnH
zwly7HmN6RxIGzCooBPdNG1dmkcj0yS257Wh03nJtOP1WpO5/PBR1JuO7ZkXgLcG
ZKLOte/aawwuJpJp8LXub+BCuYnm1Jx5OS9DjlYUS5vYaZJFllA6Io8e+JtoaCJF
oFhpWkwByKxVuhvpPoYXrUgnNuwk4vuVoiMvj5wMALW//qiAvIP+Dg+fiVDLqoHb
XkeR8KQpdE0MggLmBhzraS8oRADTThh+QjBFaF9NifvtnDMrK3wRpD0MqdpjI8n+
ln4pkVqAeI1lV0buZfziVK/rmyqErZpyVYXAWLccPSnnhgV5G/c+QSkFl/RCiVjZ
IlQrdAMCjyx4Cj4QRIMrZZDdnBAgM/tVIwI6HPv6cJff9ugoKgVCbyeSgFuJ0BfJ
ae7mRsLuKSg/vl6/nyfaUgfw3jbII6LoSX1LFMsE2oge4foIay1RIgLRmhDXotKI
5/rkiZtEn0BqmwsjwZU9J7j2bmzRhRpeT5mlSULLDIrSdPy9GsNvISBGjSVqXdbl
KUGSr6vY4ETENIizJRcYuCagbY6XvcmUnOBeK/6I1DIJTq2W0OpjvU8lFCcLNWH6
4NtH4+T4DZMpnh8MeKjQM+gSwc3Kvi4e5hHtcqIPvrhz3IeIZgTlEES23nGN5eh8
rwo3uow0bY3cj+u9JP65Nw3Wpn88erUPhyH7ysrMPC1WWDxbVFPo1Q94RZVGVgN/
YE8DHB139UH0EicKwBoDOytpw8wZ0dM2mcGRc+Ur8f2JkN+ZfnaJN4+xh75pF/4d
ylOOtmv172Hpi5xXTIyIJtnq22bXEMftjkZ1ty0B6J8KyAOIpDWpk1OELgn4au0t
9R/TEH0imJ1zvUWnqijUHQyqheJKJho2lltXJ6gYOGNb+AQKebgE9Mu9pBQgn8j8
/wAKJ6fo3WcU2/T4ebKpQUyQ+GNKRG2TsmP5wiCYof9iGnp2jpmeHFrENhM1XN+T
b1Ftw+DN0FUAQEOgjvFWG0dK692H/7zuyma2inDWuEdBMScOWXdJysEUtg8kXH36
f49Hx5X/YrQ1ScA0RmKEh3LT6WD4mzPiZOFw7zap3AUf1/XL0z8j601Esi+J/zdp
I1ck56YqNXv893aAuBom3vH7Sjg71iY5TkJM1wBi/GogfFz4WaAyxXvKTZODj5eP
NM2qLRatWeOYB44TmFinc5Rmb09EfB8R1xot1TvuNREbT+sA58agmEqTogTCdgdE
ETFTW8w6Wf16DCsXsZMcTnsdjZI7OE26UYtGC9GudTfHCepR8a+SjczYboKddIVh
nK1d47WLn1HpSfru3TyuJrpw0L8Ozn1RqYyB1rfsLduZotaKFk28Fx8hbqW76LDR
QxJBoq4xZDQLy99OdqGMuEfzO6sce+bdbrpJR81FXusN111YEXrPc5IVo8unj5y6
cxi+6eLUPTla9GIE8L+W7ZV3OJNMHVlu7uUZrmE+v3O6MfmvgVlOPErWWi6j2OJY
yHlpqoh1oY4aNeM4AIOJhOfbQrzDLV6G6vxx50QVerEcurqRVB45qVx4A0A6mJAX
jCbTLsNuOkS/lBSCG/AsAvOJ3mluz148+Wmt5G+eflw7pZpr+MQ0dlpx/qcFENA4
QAQEHBGaGUd88EMQeoWpFkRM7Q/W+FOi+Xe9Bmsnnf5k687Z4TVMCEK7Q9Wrs8eI
JWZORQRKqSilucJ77v54z9F+jUQ+jVk+0a62KhGdaUJxc7piOezmjPBZKAgEC3ne
fvA5Ula8gdZuqP6U4A1ZMGH6H3lJLEwPCgSXURS9qHYKbtC5ksAeKyQoRN4oLPZf
FB4hY9eE287l3sfrfiQCaOHqbOvOkQkTpdDbNprczs6tRosAWRwz2pyF+u68jCb8
3LCclWlXFDv0lg7KZAtvo/7SlQ8sNoMKeZN30/CISd2KsrjrraqGt1qrDuAnzv4K
z2PoyZgAOqQhboZDuNbgdXY69xxOzFVeN1rDnzCgRIbSobBm+0IMyhL70EsBm1xO
ZSCWFSHMwY1gq6vDqEW4R8syo3SRL3cd5tMDTcU7X9zoxYlbqRFhK4JwEO0mmLzc
QM0X9uVrb4uWwA/fIOkofscUbT0VznCMaSxPFbrVKyVnLXo91EwM8Sl6qe5y8nA8
zNjGutgpIkj5sW64WYuMTpVNDfWvyLCB1R12NWPLA0U0iRx4o78zLqyHDcDH/3y+
t8tMQ+afY2/pcSq0IUJuWtJUpfXjPX7Ubrlno1z4fWEFxyNMQQ97ywGOZybmzeoA
f1uDDlMcz08pRlYk/vgLLptDqxRUhh1QjKeCCuhJTW3gyhQQVQbJ51BAl7Gt8HKc
xCOW+jXNvzDR4q+ILU92ik/GJ4Wuw/NwXNIl0cozR1/SmWTZiljkfXGmRgLOB9KT
amrWbTr+wMBUreSqHGnxVqLnxqruukSpQdAt37XNXsxUL/aY3+t3r+msjlJ/nZJA
WqgsgbetaIQEEjN7wUF6fPRk8IxLnUSimc+gR7TFuVBbGPO/MxgAS63KiHfnZYMn
yIqPuLMoTn2XzRAC7G2JnfzzgbI574oWi6eYaq9U/VyYRHrUAPKK/zploR6XMaM7
UBaMj4IUUlAF2DqPF1OscY0cQ4X/s156fT00eLA00e4YUu5SOCrUqtEFbRzkWx/1
IDnjwuCAdo0ma9AT/xMlQt2urbqnl1Ov8oFkCwnBM50OSjVRdIuVqHHaceN+Q6Og
BTcoGdwnROJN8P8aBmU47DjUOXBUhVKZrsyBanRjRZmKlK+fMZ5Av1zOxVZi0pDO
u2pkVTsDSKSoD5VvG5ojywjb8IjA+rvKUiT5w/CqHGBlZuLU2uhcb9BvYFB63GMe
C9mVNNUv718wqLziXxgGX71bTulI623pcl6EGCJs8RXerV0MUHgCkxgZ1OmJgnas
HGR4MJcRKh9rhFHbfWCDbaVJsOL9vgZW5sBjlExEQkk8OU58/py0lSG96WKmzftN
ke4KnwQiFycT0MZJ1fiBS805GJW9R45s+ZiG4amBHmkxiQn4Zuwv02Ix9yYvG7AK
RYPkmdG1iiTJXr1JP7hMmdOzgrt2BVguO3t+KqzKZfV3rJIWj9MrEilMtRj9IuU7
QjTWo4ziGxH5fZvSBpu94YzG7gtz5o3oHDMg+a3LCHu+X9T968AGn6m+VSeGFJ+m
homtiJH/VwuWU5Fe6YVDM1iqHbKs0Ewjw4ZVYBUC4uH2+PZRzDb+Dj1yQjEHJz2r
g8MsDTMGdGmGI+izgZ5HpdHVfjXvDyIe0QyMYZ/Sv8sokm+SzN71M1EBJpeU+Nj8
kasI9T9joZaCN4r3BqiorbmFJlrDBy7HFivx11Dmi4qONCXHbPszLZkQ4V8lw35y
ZK2dIG313aj9yzFCrRDwRYCaSpagYDstceuwWPX0vgUA0uaPzOgcqJSJkMUpmPvv
2wK2JCCXBIYLvKDz1KLqVKRgM+SROS4eGb4bhcykkYOxwjoip8/yF3WDN8hmYGTV
8ZdehIX9oYsCKsk2FtmJqhVIbUoVPzCi4RCVibSdbH+p4GE9t6bvxbSAW3DCdajR
s+rNhsOaNNLRWBKO8l7MjcrAj+p5TuNxZ20XH7EjfQfRTNgw2DDT2D8DjmwgJlSQ
3SWe1S/TvHp+bKCfpJlcfTWOrfKQqUhXYHhw0v4hCHD7xWAYUYpe882XZg5kdfW8
G9+ajNunAseZ2xjhUCMkmP2SnBbSdVub3a5byFuDffVhofJKQx+Hawny7bbvI3pK
EaCyXQ30GC5FARSpHvapwDElotqCcL9rE1C7zFwI9lswjA/d2Ne1XdOERNkoNLv0
c9b386raUQQz2XbYbwqaXnSQlvm0xV4z0zhHv/LV+vbKTNShNlUu/oXS612yfhRD
waEeio13IlFhVXBoJBZUHBAo9Mqbfx1Sc0Bb3r8slo+WUHNXM1ZYTLAUUJM1BLIB
11SqmCYOEOArO1JghqjASLGwwruJBdmHPzwWjThJ3IdIR3oMikn+QtWHAugp7xCr
uYqDRN5peQKflSqQIpbuy/XN8ey8RXVKPA68Zbi2K8kkfbbc1xlf2qZ0Gp+8z+Ok
dOO7wX0ZCgqd/vSswABKKZ/RZCuURwPlWwLX1cRqUP+jGcdt9I/+0E9+pn7tdMa8
zbjJuNohVHfAdW8PhAJtFtImHztkWueT3DxDrrSlGxRHSDyYXQZMT5FsSFYj0FTW
pJPmIidjrGCvdvYM8BSdgrUxzGnRXItNVl5xAeXFbMZUhpiw7v7L7mGiVwLImpqN
FT17Nf3Lti9pOQ4FrjcfEPIhjz4kBLOYinhBPXtpHjEW30dvppcnxfiyEUSba0WL
Z+R8iE0xBenL9PHdbDLQMApEcayNaZYgSk3nStbOuk3ZlHyIJdQ5KzibUAtTE8RQ
15dExKgwZhKpDbOqVyHhHBOgPetRGqRVPkDpNaCqy3qhFAMSVSJcWgex/PuUNFpU
WuLItl/eFHcevTTH40D29ucmrEK4/bNM0mPTm5Scg7t3f71DTv67nTrbXkqItkr5
jG6/Btl5usWtVGtF51sq28r71TRHSk93uvfl1H4k1YFLxIlqrmtoRGKwxtShiwjf
8+jMY1tSqB4mHtWw9k/diOVjR0EB8kqQ127sRtwpQkb3Xojz5Zc+RROruU7mX6k/
OBPWOf338CuX1pSO0dRy4tejMrYcS2bUu4IRGzjzvzV3scisaBcZxESo4xCA/11Y
DTxk+3XssW9ZrIAbREdR/3lUikVDkzVTPUReGZGmch/UxgrleAYzcVR0PKItY8fC
9zjH5A3AuUyMwsOPe8sRRviDo4gbbhNAQ70bQxjZApyNjJvVj5FIjfgSwJ42znK5
h1+oaHz6gKXUJbFRakC23I57M5MAIq639xuBUn4kgGqPatilRkPX7bedPzUsY6FY
jLO1jf/9sA0YmZqQggvmzzrCE05Lx+kfAIIkfpqFQPyYtCl4gPlMvwVcmLAJx3PY
gFdyyLY5LS0Ngv+TBfZ2fGJdYG+uEdtjoqBCJNie3T8pC96JpOph2BVSgbtDmI54
gF69Krzk8auMT9mMLISGnTNyhosQV2q8exNt0p6RfgbfGCMVNz5y/RFbEHSnkNfW
MKhMDA6hp9VBmH1CUcvZYFrwpj42SFN4nFXXJGfvrHIoYmBrea4yAdkbrZAvO+3U
DhznrCAJZPlgCwOoK5jeUhJnuHQlb8AMrFw1m6EGj9e+vV5/sBlsuVjyBF0XrKIn
7GydsSz7ub+SQKNb9CcpSR9HGb7hl6KZXY//B3c7BWkh/DtZaSc6BXeX+7IHrXZG
HN31QuPhWKt7f4dBHstm3ryH5pq4oowV32Xjfp3uPchIEicH0qyGJRb+KLRJSZyh
J299Pz23tlbxvAM4BA9ofitykKSy9lq6EqK6EKCoLHy9uJfZmbuCRa0QL+bTn2BR
YF5NSI8U6QCVvm9aBndzDShsMA9un2fpraPa2gAy0UGqGhAfBdr6uaIwnDJpOSvk
qBUdan3OjdM9wVVvScpom1FJ12iaT4d/5BCnJfcMRlgaOUnIfc046jb+hudQXq9U
CuZAIEr3h4PGiWx0Nd/lv4wHvfGHPWaXOuEb1Beq4G23OURBGFgrq3SP25PziKBg
R2sLHnE/IiweeZAR8c04qkkeDKTzgnRQV022CCsa9PK7BZ7z9zGHEll6SodUMQKs
m84R9x34eM2MEaIa+FZ5go/9hknK9SspCs95ZemnxVAwNVCK07x4y16/MH6dKG5a
rdh10FUykv2vMbAOFB4Z3Nj5P5FFrk1lHFOO+T2lrOXV36fxwVL4v51BiyYPLZ02
SHXhN1H+ymxEXdqIHl2ZdXTJzwk5VALXHgFjv1JckHKwT5hfnZkfkOiMegmLBLxP
h23nKOjSKoXDWwJcXF7DzBiW6hMBzhnhbzx4EwPo0SPe7y3InITqMcGt8YcWTB1I
JQmuCNfCL7xHEocIKKpx9aapFf7EHxL0SScPgvAiRW8aCggXS5OPfMvIeB8mZF3z
5glGkZtPjT6iFZSRBoEGoq+Kw4knIBh7atb4LdS5SJQK0aeQetTXG3URZ8o3ylgD
znKceyPwH22IOAoBlJXDCC7OWjQtlN9Q8PGIp/l8i7gGvEeYQOvhemH3iMcaXUKU
jJSmlnSSlRVyB7reueSmYe0yEZiH4EA782eMQzG1QIOoYRKtcnMQxUBhjWfhLdcF
aBFNg5q2XCYFtNGJWXsyKT2s5SklNUItuoWWfCrznsG1COSS7I7pL7j7PUFCbRXQ
Vj/bZspDqpAdGgEj66mLnD5Ag3zigAA4RzHwzFkIDdaAywumEAmfFpU6y5saeUB5
p44RrNg2/Qt7FI2NYM+Z9RI85w0PAPPCqUPCsyCtUU8HUgDwb78Jsymbhxj3eGmq
CIw/GH2sDCFu0wswcITYTxeOizcnfd6vPWtYkxBkdA3GKffZqVUg52w3ZftsRpg0
Mio9mt0bOLuMcjY/yyyEXyK+jEwY7PlFvkGit9bmAaZVdOh3Rvwsr91BqVjppdLb
nfKF200ZpvtIhCKEgHXSRMkfgVS+NO4HHiSNkAbBlGkNf5CX/yikhHR7Ti1WLj8x
UFkYxMQ4OaXyWHRJqsmju6Tp7gc91QeyMDrVLmpQLrUO1ItOG1bGFKbV3ivdQTI2
pjK7n1/iwDIK6KN+AiJx/lYBqCAi6gWhKf0gWVnwvhse7rC5+Yguk3jMzkIjvD/5
MlEQS47KpEHUzazzr91K9U1uPruiYprhz3ZWBRNOANdJ7kOlQH7K0Mwnb0f87XmO
Iy8XjmzqexwcVIUc2XV68j7DrjgpzjYCHRtdRRwspzGy9xeeCJabavh8RPJtQ4Ph
JEu6acScIaMbAQtf8IUg1SCRyxE68VTSBncT7+yWKm6kUBJ0PAEM+q33eJFOPsgF
jsPSwXzpYlkxHBM9W7zujx30dFcQ7pvi6T5m/gcpcFAetL3iBf0qq+gu5T4t9FnL
jO6o4oasFGMCOarymt1HxyTVXjJezgdZQ20qbCRaNKqaxKdtMOtXBwUb7riXGnp6
Od3UycHx0S9TmdIYzqjAME58f8QmYP68AGkK1GjuaysjiAI4lUBllUkBjJaF9E+7
o4b/I4SaoydwH1n9Lo/FsOIXKl7tjjvoertLAtvtTAIoFKcYRbXAO9RczX9DIKWt
aqEbDxit2KM18MwoFNf0cYIrbE1rBRVvVfyw9ibLh+39F18XDt1ixo8QLCEWRBFV
eZwmiM/8sW7N6N/E4j5ypL5ms+lmQcEzgUq2BiXsGIki7tqQVfWUF2b2/W164dEU
Lp70fYAM5mZuKVbcXCLAACEhfITzDXCP5X8geoXWZgna6SbnG1bwi463lLu7ZyRm
V9RKxoSz+3eGHpcOeNom3VmS/lOgDFE9bncK9IhpMn+eR9QOSxWTlBW8N0ilr3UD
N4+hrB0KpdNibvWwIx2IcJ/85kn5BGRHi5ALRZ6JYIcRL4T30wCr/13SJ+N3ES2S
CYia2XC3XJzs1UK4+x3cBe+zkGKqUSYq3y38C+idFBIuET3UobPQrdIT1lOi3kBg
W3MQkqO+Rz8Wx5vknPUkU9Ro1naOEVpM5nt4XBhJYo7wWAFI5AUFFQ+3FWfczbSL
4wkvqnnnTrypRWJGgOHbrnc/eVKq0+MGJM8SC/IUGGEAxjZl2/sdo0ylpb4y8cBm
kGPhEQpMPdmSsprB8wuXdPhs36Az087F1i/Z2zscJ/4atS2J0YBEZ8xuZ4k8aprj
CnH8Rp4xWhTMXUHpBnQuxDbWztdGKTsEUHUQZfjhlrPjlw2E25ZG5gS2ikz4RWWp
hwaUrCMOhavcynwmNFCp5exIb89szbL/iNyC6HxeBNVdhx1IBI9fGskrH6wvt60q
AsECpTD2kvY+G1CmLGR8NHc3q9yWyczSlANM50ME3cjtXUrebwEwhv92jk1GzO2u
XTeDjwSEyC0tQz6YBxmY6TMFUJqOnyF9R57ShlWCFcVAL87qOCvfuPpg+CfBmz7R
3SWqvsr7hQtfK0U0jXFsQ84l3xGjCSY0ogCTacxURfBZUtCp4xH7NKldNTdkhwvr
+phJhJmezC16Fm8KoI16EQaLgAdpOHUSeHgoHym5neguZDYcqavoWoRS2+u/XhLo
A+0Q+hZs8BkcKyzPkjHuaGJJE+5giSVC9fUr2zlxrmw4JJqBfh98hhNhaZKq6ogF
LFYxMBlIuDaYgF4SvgSsJx5dbSubhUsX7FarwSSFuwwheU65tgIRIljaoQSAHYK4
qTfWXmtQ92775UI6l6eeRcUAR79AXIir7EZfqv0dqxWk4N6mYNdhWhba0Pi6aZ30
rS3plEzDwE4rIlNUVRITz0Z0Ro1S7o1C+fVI6ULMhvAPVPICQTdCyuGuc4llvF5G
E/eefXv15iPZ8kpz0ZluEHD6ZXqpkmS5j7C4exEmrcxyfriiW6thNsc0P0o3jNGd
sZLyKukprWdHb9pwOUw9fBKXMQBTEVBfna18Fn4XOjAY/cfOcLZYgB9mEcOznZXx
vAOol3wNZOKml9SfUrtTtrlEJLIv4gBdo5/tXcSwGf3tzlGUa1tkKFq07azBOD/B
8fFIe2A65BnuMHsIuVYtSzT5qFEGTOUyOhoZOnqetPlcPgG/dIYO39h2UV7yWktI
NkAWR5Kiwbvwdx98rUcgwvJTJpnO8SznfLQAOi6jQ1Bv3Ofed8lEoZMTzMBr5wQW
UIXTWhMbeUPPT1MOsvoYz4jFqidlM2sIs3Z8ON3gFQnmoadeQ/0/7azHknjpm9CU
OP1x9VGcOGeCIGML820NTnbkE1aHYxQ8CEcX5wazfqVLreTg9pVxykIRAgGSHZd1
86PkIl0qh0M15WAu60IRi01sJwYPWC3lFskK6xiOvASoJ69lERF9+X4Vt2RtR435
JCQG7i/cM4W6BgDbYtB1ui+v7XaCf8pw/k/XgjGS1BUezD2cVCcuDKB3oxN3OlMa
FV3NSEawJDzFF5r3VQNKxJVqeawIBgvQVujMQNL9Qsxg9HgnsNeieyCNs5IzmX7B
Y1nETjcxTs94rn4ahYd1EruFXwhv/V+aUKQssAen24IcdbsMQXLIoygGpHVN6r/9
Bjd0I+5pzOR5b4qkbBiG91a/fAquDftdNjNgQ/e8OpPssw1+MAzPC0mWQURJuBjg
GGvMPW7aEnNvFOghI0zt3D0NuyBYC9Y9TC+eVWS6ySxyMiRO0Ci9jv45HMQD7mDM
dL6iXp/Vi5ksQIVs6UXWjUj3wuXzgRaLBfUYjyfIaY2KGhMDgxpyv7bmUCLOqXEx
4SS0l1fvIbvgId9KTWwuiBPElHDaz0EZoCHUYmUlDsIouly46A/hTazwAQJiRLWK
HrHPyEZJd0PghpMQxUzRNZvEGzdes+Wopcov3BRfG4MgTPdNT5oteHUqemEV5RIr
0AI6awf8/bFNtN7WzIHD61QsomvVHpYY4dXsp6Suq0GPhr9uCKIiqIuIfftxNdzL
DbhbSqwABWbb+pgDYF3mn8uy3oNi8U/Zhl30/iRWKURcnjDbiMsIbuxgqQE0aILb
dcl/qtxAheTbdXQ9SI3dCeZb7OCeU+gejdbDx03/vmbebqDVSiV1A0948nc7KK+u
09bhZdj0RCCmqjDtgHPSTDyy/6UvJuHVR44rMkQHCmIA+EfZTHME2/wJESaEB7xK
40khoICQRPLYpGcrWBz8IASouCDPk70P2nTs0PFQX+REByXQ4Ov+GGRXPDPJrUhc
VZE9+f16MPvQnHCbqSoxDZxusClDTpJa31OeUMLzb5TF4aVK31ESpqSxkFaaR4Ok
KAIGKygKAoyVONFiWf1xhSW2qSSBsr1AFwu9po46Nd7pTy1RsVWNwFkV+rqCTr5Z
4puG5DP1CNIbfR6ivqYnjccOVEQ/S8HFD/X+Cs9eH856AqbCTiE6HWTcKJFNYMrD
BnHZQcnUcG+L+ouHS06BxBzPpln77Iqe/8CqLoVIkiNTL16z2ihy/10pS2TjIeDF
xZXjgysoK22/7F8d41TCRT2ePTc1W/BKDP/OxuSOBBLcCUcPjN+Yq509PVkEZpJ6
lgJyCeKbOy+CzE4BdSsbNBSHb//4gkksW85RsIcexgCj9A/lBJLP34JMAOuDYX7B
4VtSSNtJAViiVqZm8Szh4NQhdV/DV9KIUK8vTe9QztBL5nLYQilfsypm7uWXBljK
qV2IW1eWgaxaY7GHH3BI5DaxpjacmLJpEFlIIPV030FFTKTuaY1W6Dv2dOP7XfSf
c1V8OUuK8d/HbWopMxxJACu0JHUHvrCmklIioFTWEmiUoGoI8ik00YPFhrpw5wd+
xtXRIJfXJJ1XbJ0KA7MnLfQuNbRns22EnmBomDvfIdwuh0y4M6j2vPGlHiYDodLV
SIlvOa6bT1wDKNAuAHUbOD2NlwW23fyRaLK//8Sr/xnuTwGGbnx/wir+d/jAdb0S
rx5hdw0Vs4QMXHThdv5zflHRtDL+TKUdMMqOceZ68K7ol6iOpKEgJnqb+fCPv0UD
R/GC5uwvOhEzOgaHcpiEf3v/PSFy6N9I8BXk5jAianxcFLjdMnbCoh9G4GAXNdEG
uNEpCGGc0yLWo0aNY5u4o/NoRoDQCWX0UKwKwNJ92ykwti4UJ7aGlQPNlAeuogK4
hNW6oCT6r8Ibz2yZAT2fGaRh0LIKdXrDy1x6yk7eOtJHd0PnatgzKes9YdGxl/W+
pPVaqZRgQ0+P3Q0onEeD6ISTqgvrnjLyKDVFtdtzI556vmqs57sYdO+wXxAqVzue
V6R4X+na/qi+24oWC6THDN2C1PmBgQpmjmq3t1dBhOHk3//PINVprI0ijQg8YnFy
9XWZEaeYhsUDS1XMoOMdoExRXvgKLpBtP0C1jEtoYfdQNSPRcW+WnVQaQBsQqGsv
nJ7EZrqrsr5wxOUt0FX1YYamcsk3FJlzG5wZSolGfEws/xARpByJR7E59WwXUx2o
+O/RSc2Nse0SIpzRGgGIkV+p+A9vfxot+wHgOotidCP3tpx8p3juwAGN8pbUlyKh
D/McnQt7PDRqIHzS72DNQI29g7EPJzjZeWeadUuAgH42LetKZ03tlXf+GreEmpzu
7seBvyj/vQUkgjjGxQN8kPs1YyvHpLY/AXUesxLUOTl8aatesh/lS+SYx19PxeoO
MxityJk2oo5xI4mfmWk3/HCURzd5tYRYvvKBBtHqjLiNSW3osR5CwF592msZnAHM
MAkaRJEe2FK2VkLRLzeYoVlZ96NSyAkNn0sd9uAt+Mx/Qi+3xIOfWqHG0JUfNsY8
yMjRLfMqCRo6sATK2a5EttY1upyTMmc9mQ02PYYno/7xxb9pR0kwB1S6r2tqlGZf
lUXX2+QPcWJ/VuMdQbY0dCfaNGZT+jPDBGq4jZLLlt4Da7HMueeVp+ZkH4LGa38u
SL+bh052Y6q/nQ8wzAgP58PUiQ25QNXAkMqeLMkfzeBpQuQ5/ntNgCmc/OajduEk
3oOJgebr7rupXxBgnpFnT4fcJgvyBxq6+U/JRF7icmPlH5/yepSLWHFMJ+2r/qqE
JiALZzPktivwPpDpo9QEVz9Q24lY00YjUfxa6ZG2hgmgwH5BjW/aTIhtFJ3VY8Ht
mviQlS6zF9o41kXSpfr2Y4LXFEJYMtqR7hxCCjhzYvEMAlJGF7qKTFc9HeXOZzHW
5VY0YAy5BK35mwskbaNHKb/xRWFWstJZXCOsW2aXvmxhiJzV1S0Zf04QEHQUPUxq
qOvs2ng+pw6lFIlZtiTM0XCVUelflM73ywYwvYfLRjBp2+byKwb/ScZPSTxkHQE7
kqKKgkQw9bi7JVPo1EUXDgfnymgT7yOsOrokl70d0yNoc5PobqRxuN2DV55OueMA
adnw4IgvqrL2MWiIbEwpVtBdUhb2Y8MkS8PF/d+ABZ+P06lF1JU0RZcLXB4N4MpS
yQt75B8rA32pZe/GRHY4WCAS7NPjU5dLtBl46IyhP4ktDP9iRvoaagl4AO5rgsd6
4/NuRK6xF4vPxrs5/1GpbeJhFF8NWpfSx1qPNDvoocPiPZkmGQfV2oEG9mEH72XJ
5sl7STIS9XQMDtRqFd1bMLrBov/oVSWF3SPg5S+U3tLs10PYDpEuEBRDDwaDzB6X
uphGDYLxykCj+0SGDD3N23GL8ure2lkXUMJ94twX1ih0YGV7KQI3i2an9tU7OPft
ACZhkSdHICatIPWDgIFtN4TuV9NpF13oxbY+SrZsljQzSGLccg21ZsL5EKQ00YWY
wWHWB1wtudxhivwOQ+61nEupzBXNeAwFyQwQfhppgl3N5jQmPiGDL9aWFMl7migI
zAJjFXV5ENK/mknBSBXpG2clqZd2Gt8RwD2rv7wBXKPl+VKnHH0fqm4DcvSEVJ2Q
iz+3U6CluCTl/uk+4N1OdgttoFhb3anZ7OqnSNmH5jCdtznCSj60zTFHB5wEuYLJ
IbjkkRVAaLksSF715taH+HKuSha09f+EyrfUHir0ruH/WabuFi2XfTjNWMmVat01
d2x+kF7Id0BQS2rFljR/yxbvOyd5ZdouM4jvQe7ndoQd0KPzkPISEmJ38xnp1S31
zSMa9B/w78xX1Roa0pSfVCPYWnM8KxsoAgyg/1DBVTG7OzE7fd1+bWsvY1uS1aOE
f8zuJO+rP3JkdOd7W6lF5ORQzlf33wzIGIQcUxZVpcrmJrg2Ovu7EwTI1FGiS8uO
h0Kfo++ku7pPFHdkFD2MtCejK9NOFpFVHaUR2YT21f/qAt4Xt/n5PrYKgvFU3KCL
NXmRS8nvkeWER9FsCjbZLYkxOxLaQQr3roTGV9QVyEVMhxyl6dd18EGmd9ztBJYE
y53+2bhmuZY3js+b2WuCPHd6lOKMMDkWiR6D/k5vyKKUyD4POtnbOxr2QCAGHL1N
vNvls3XKqvhnXCtmyHcoMem7aYKH0bQIBpjm98DQ02LlXp3OoAT+o8BxIhaolQo7
tyk0tDuzKyX/KmloDR0aNAtBheIyeySiSVamDnGgKViw/7ySgwW8BsmQUqQ16wLt
u0zfO+zRIfzIeqRnMG66A/U/UcbP19nR77DJKjE/yJDCncXVjPyCC6fJObRVOK2e
b/vof3FMhTA5bJaLFV1JwA5A62uX2ADBlnTq/e23kcUrIN5ojRhE29SzTvLfnixR
L5VqM4jWOe+cuLvuB31k5/32Q/Vfunzk7yjmFRi4vWsrfrkEBEgPee1+RGXUXRWx
4MyFU3wksvknFekmrKnH0vdaTsbkXvl/4iQ/LtWD2XHQ1UX3w4vPhPzEFtHcl3kA
daGKH4jB0Jsw0ilKpllCINDupW4i+3LOvAAAMzshhoKUk3Mg87gTI5Ia9UVnJjSh
EfRk4XhwfQV0rdmKCz9MKc8ODlgfV8AjkZjhKGl0bgd47ZeJ35BzreC9dELL5uks
N1/J7Ogf0OO0qATNgwiahqbOs+U8uDGGGhlFa4NApPQMjsSiGWkIY4LL1xucUWpU
n/6qIB4ge0KT0ZmjM6QAPaAXsf/K2Htw7UT7A9HRKW4aytSkksfsZikNed/6pVWs
IVz/AOdXiwXxLLNTkby98a+zXGxMKpgnAKvMKqdfiMOhEYPMberVqEGsdb2Fv/OE
rYIRHz7P97aJq90AHSHuvaUEyR4Z0Hn0iqXmkR/t4nWfHXZvmeJtVZtQL8nLaDQo
IuZwtiQ+6q4vB7nIcN/6AoXot8MRAT7U1SDNrUr1Pn/+CxLN1WXbDv3nJmikOuBv
1uR8+93i6Gyqkgh+m9PFDElOglKoc1AhdJMljSV4j/8EG2uYwk15dkNbB9qeNWjE
DrwEfP4VfEvCyGwNo58lr+cFaRyioPYkr4qQShyq3nktwoe/zJcPXfisC8IRkeRp
/sHLSayYDGPCSEWCqX+Jh/e/T8S8qk4/KekLEG7rHXdyfE4RM+ZBgBwAp/zHcY0I
oPdxJMWDt4obspU7qkeJ8DBFW47jHHhiy6np5N1zz76FFByAKzbwo+b8CNQh9/E4
UA7qKeFF1akgzt0ylFHVBIlziXYZ2ZAcY69IbM6P2YxfOCZtjzqzs9gwxDyBLN9E
msFu0e87e6zWszBccOTm/XhG7mcKMztstbSKgxDfAaau/eUExlPTbnadhPug/m9M
oz0q+G3OYQwt4LpkSgRbJLaqy+cQbd9eQzCBjcmvHfxQbHVz6pzD09jTssUBw7lq
hF3JcczRtZAwxEFS8qr40BNxrLllR7DFAFSDh6Ynz5VZ1YhIXdzQtz3L4i/LzYkw
UcmTAFQVclA/4CJeT1c9BBH9mbUrxS/3StmsX4rN5t+INhK7SYQLZFV/6dcCFMK3
lqZeTIkwG+0nPi7LHHNLmLV5emwyH3ipGz16yokXW+/7gyXOyDXG5cPEpK9DRRtX
PVD90A2sh/WJBhs9PE6v/s3gTaGd2Y339RAB1B8qzzUtJjRsZ0Hw1P9YrPmHOg/K
OIjTAFfK0Mv2nNvX4dlJqnOT1E3wlBZDf47++TNK7Zg8I0buSKWNWzmBcju7hT0V
VggZ6uF+WyMkh9dDW7+UTU+mUnRxRh4CHpPqgutTR8EXydZO2YVzRZLImqAZ1pmd
qIePFIotsbHWS8Izm+/VnOCzm8VRMpAXJ9TriZAxMzu1+F9sp5GmFDCX8lc8vv6R
j5EPPF/s8w/zUTLGr0ydFYQtpruI2xi1XrpOjYCwU9LrEdPTyATklGlPs/ERdrnf
lKNTUKBaep+AzwQsDR41KgqBcJxNNwN+6jwnuYghUf04EPRqWu56s5iD6tKvOzws
eEOY2cwdD58XXIqnBKcfub0hzvRBsLMNMIqEZtoErWZRuVZOFWbOo0MGWjq8KyqR
/QOpWc+ib2RdNv+htJez9XxIpg3pT4Arq8agDq/W2sUK6PNbOStrKKrc2oVl17PT
y/Wd7CRM0SE7a+X/MRVBMWLZLkUN954mMyL+y95d9Tzwer7eSsjzuI8nd5CZtHEx
sGvcuCw2NyVGo5ZO/eRytgbgX2ykFKXIXdSOFuzJ8og5ZN1Jx5C9loCfO9yxCAwr
Th+QZXbZC69IIq03igD0/I3UEUVMfYdQBbS/3IXsoHdBHZpmpihbGm1b/8CwFgl7
v3y0DqjPZGps9FWJ+bWjsUFzYMcBQu/YcyE+1gjccIvwaITH/txFPVtuPOXlEyw3
MkF8zHlWB4bD54e3sTbYwhqhzO+K6Tt1qdfl+quM5ue12bEERyMZBN8CaE1UPTn0
Tq2JpiS3gK5/HOBpGlzCHsQdI81Ad1KO9FisueZsZ12j7+lYf4kjGiOR5g63lXql
IcB/ht6mNTEXYU1DCiTKDNIYeBDwsehK9V1kH+U4VDg5qMR5uXzSSEYUUp1dvaiE
6uQitz1Y+hL4+bcZ/sKz/JQVuQuATl3nrEWvCYqM/1YrbCFvIIUaMKwEP0Qximkp
hpHJ3rIELORLhMP5yzO9hU2BAv/Fc6Xw4Me4hs4l0m136c4j+YA7q1m9rUuBu14N
DmcEWCFY/1p6Spjzyp5GsknOYVd+Y+x4+9RlNKk3U+AI1Q2kR0c+Fmx9/uzzlTDy
pD3LOq3AlmenPzV4m7Yb4SrHGKKrHI9n0DEJPJLlsSZOkvNO4/8HeTc9WGrgBhn9
PtuOTpY9W1OahYE5t5Ir2r64hhj+fSnduL8NVq5KwjrE5ENMjnHw52QsVrqevpY1
asnyeBgaKDO7wAiQnDhuOjYUqnnh7V9qlKEMXeKpQ5NGgUa1BoyTOoFc1QCjvd9L
+H3eaT2JOctaZHQ7LCsCG25Y8WJrr6riPa+OlKqL9Qzoo3Hj9RnqUOBlga3LcqkR
lYPNaOFHtfXHEAHkzBDKl83IsDNfTq3II1azwdvldGcswbKoHjFFUMVBrOFRAsah
j5CxkD5TuNMJ0SHdE3Zeqkk7pzMoTpzYbwqGrJPYYS5mpYFmgcapgk/QenCoBVE0
2nVOVs1ESNz4Yiu1Hh65AkZsRLOry79UuavLOOPxGClKPNY5C+nAkK3iMHUtw+4d
7E8qJYV6pDS2d+6b7CEY/7C4lbnfRGyvcpiXhqHWtnLCVFSiOWT9+vxXhtZ/B4ek
Clh7PmJiJxH9aycb67W0vMK36R/EMBsE0B2Z1FP7ginnqwh5r/KJ+Beu6Ej0Knxn
VFopGaUTlDdhPCmHHrvGta+US43id2H9TviG8UtYoQ1H5pjprN6kmQCwfZ4TehdT
g3b8XqAolJeN7MpDEpYaJcqsYCJTXwjYAqwaZ6z3hnvuWerC0JGTJRyXMA0AcmT7
g4boPkZNSNbUsg12mtUn8txueGW4FrwURwz5M6RrlC9IP4lrM2QzIP0hI4LF2DiA
NXtSWxH2xVbpzllnYvQ8wz6vUx2DJrbgogXEdjE982PIfeWunDD7GBuIADZzTUfD
IwqDLkPATXGsI+Ky17I4tCNz8wwlcNjZrJ8xPasOvhcp1t6E9ikOsU6qPATWjW8d
qn92/YobmYQbVnxtyU8ZrkSbU+6Rx81PlcdJrXRtsh6s7K09jjmZI2tYeqgdt6sw
ixpS4dRBca/WeX6fF+7XIIKo8x5kHxndtnA+4RQtzJhfpfz55+YeTl+YX85KJhXo
y8qqmhMJiwc6gUw4d73GVDcfl5EnGgi1EctTqRuw3ugeOOTfSPxfLcWyJUNMA6VR
cmGyg83FpirIq4CoRUA/oJiTwsLFnDTztxGBHIql4vdAwwD6GHvzqV/AliGi8PCv
3cC0FsUhMHy7NvjbyjmK5l2Dkf7kY5E8ND99ASZmhOWVEez5HpaMnB+axmTtXjp1
xD8PaARQJovEXQtq9IO4LTiscBT5zZTbuBW0A85QGee+U+QWYX+yPS8u/yZUWoOV
AHS/dik7MzYZ0uZm1yQsxf9BfIYjtMpWo4305xoiIsWkwBsQacaBs/80irsLUfy4
pDM8nxgHsPy+FZLL6KOF5uqV0gUNwBpw1I0CPWtPwXRaHXmf7KndKBtRo0oZfA+d
gcq7OQHPzwC2BBLTHv3ZyqFIiaH6GGej5gCAOtQn8nF8MabFFgoLzv7qcyFuyuWu
pkK7UeF6PwaZ5tbthezP5kezPbDp/dOR0zfi/mjxn2qcPWd7JP90AUmnTl2ot6oY
Clwo4j+9dbUFwwkE32o37VBnO+m3w9HY0y90Wn5fLVs8tmon+tqkhYiJRkoQ8MEN
Or3SVIvVQLnu2YKpdw20Xy116NRDK83+xrPDq9XJJhH9/0rMXgYITsa2a2geMoln
YTswk8v72z2UEWgUBukN4QAh1Wr0COG3P7Cj/0q0k2pgIXxll5q1SoENSyuRErlK
9oSVhX1FXmL427UtQeixSAJ1ViX/WtuyxFmjW0EIDJyawHbKsv/LbuosS7lNqeCS
fLPZbujcHr8/Jiy5Ma9pA6Bo6L/d/t5YOJl0o9sGUpl87jMQY8kFcaz14RkJet+F
9WYBCeqCCgY1kP7isS5rHEHB/5fT2+6xl0dle0h+roHtGfSzEJlCX9ojMpOTLk4/
sIXYU0CdsRv6G+XDy6dkzVjp7G3ULorJGtCWMSLg3olcHoy3z90uBWsGjGfp3IHv
IMS33+OAeuclmCOqjrfmK3c0xQYtA0LSZUC7x0XmhMri2GinoXFoc6PucE+nvBU/
my0qA5kuZnboaswCI4ZK2dDDQrRRf/ZLrK4rVEuvkChDZRu97dojpdudvJxP7dZ3
lb2sYWbg+XvGIkJTuXUpMgHIgGga0GuxwsxJ2VgjhaR0pbgmcxiDZNXdQItWtTBg
rWmck6BHrunVXRffFKUmp3YFjOiYxhJVDc3QgNL2wn+LOqh8JW0u0il1GNOpzn4Q
ubgYURbPxv9f3hIprjYp8stenPA3m6woQYw6byt4eYrGxsyKJiJ9nbx1yQX0PHow
FNgRsf81VyYXX9rLj0hqofSpePi57o89x+RYiJnU/vM1aa/BlnclB9gjL8vjxywY
HLIFWk8QIdmCZXD6kk4XEWniOBl49G3J35sn4TtdIF15q1bW/XXMIifBhlcJkn11
ELQq1WBFWdoVBV5Yab87snwKBoptUJ9GtIpHr+fUDWyncAKW039VZJJDLaeC6cdc
mKnAz0Mk/kRgbkpHPSaX/Tyu/nvLSPEGfwJF8WocSeCQnTfU0VKgw5q0KQDo7hlU
hFWCYwEvt/hD7cyKiRza7Mkyp9wPPoL7ztwCI0yx1eU+IEWcaueJ1Rlnob+Rkxjn
7VMmUI/OGha/gKUBTniX6BpDCRSBHW7aAA/Lktb2XlpAv9UhfrknKDbDzWhw9cYk
dhP52Lpmvb1CGt5BCBJUJSTVdw4QQRRmy10Y1Xz5imGGqcEVetDrG1YXRVMMHBbq
8UPNbOEN2Jpy3lAkNj78gzu9/SSReZfw2YnTRSiBbaDdGeLXCqrXZKnwznNjc21y
yuRvMvfkNPsImcTpkyV9vyHrnc940aFn/flvfI394YPYb/XP4yV6HhmfU7M9bcRz
S/by0JdOA3iFyej7bZeVqvmJ04EP4KV2pUfpShUVXgmCtW0RXA8gSdlc+mihWZIo
D4r0LK2wXa4TSKWHaVdzFFjGD4Lu9P4VxRws3OaQxZLH87CrdCbPqdoyj4CjPZGa
nz+QOifIEDQlxcS5Hs1TH0Ideld55IH2o4rFHKNPzpFJTLFRzCypjRb3Qb0YAQN8
m94iECTw4JjQSmsv5YoGkCIbXNwU3y1B9dkWkjYk94TJLeIAT0xrBL5OdXOG4Loh
E9Kz9a8P3SzJU9hFCCsB5U8KeFRG878GIvXmu4CmXfoO6cxKl0/xXfjKdI+HJPpf
PK67WvOFyoHyA2fAm7pZO2P1p8/6mekINjm2m0pnYbh+50iA6Rhg0BxgMIxV940k
b9Ln/nK/1bIIW4mvtvlEal81exDfxEjpBXS+be5UkOhNORRwbrXJpQkfPsttjnLY
swN70QCJQelbMBQzIKV/u+yAtfgckff2UCq2w7aV//gDDK7+ZP83hs/8dg9+oXhE
CZ3Fpx0F3aK2GtJAcdROsplOV1xcFRXruGSMQFpy/zCFjq3jRQFfb2Zml9Oeco+z
roauTZ7VwA9DDau3Uc7kfvlZ39dgJKZf3tHAy72sDoi96I625dGqbIslJBF1aJyv
fSO3ZvCaw40cnJNh1G4JnsbdTt8TASb9m+AALs/JTResvg6RZzCeR3qsULhVcCDd
HoOR+syWaxY7Ka6dOVJEw8noCY1gkWrcJ/r155dpSqlLD/mqhM4d/cU+nCxYGA5K
nddB4NDcZG44b3DdP6ssPwVeG23ntri5pX3hMkJtNqgXQkNBMMNz1GTPiArWvMKX
CS/X2CCTrV0FWNwU9kj4FDramNONSwVO0A9RkVWFjN+ABzxtjsp+7lQiRO82/r9Z
cafKqA1YSJM6vsp6pw7ppjMjtI2GV6wMTwMQEcWOJPJ9mXG0DrbQst881IEZVSmf
zfjmd/FRuBifcocLPoj1qDnUnLtMQ1zXNHzZsQuDq5/Ydd4JYv+OplIOHlGi1KWm
WPJMJ16eNRgAsubRKy5LMS1QHBfA0zqTi6yNgIm3+a7j5R3I2qG3BwSH9YOTpUvq
5NWUgfiNus8MBzc91khEo0Gqyb8i4wIT8OWrY7NLUokfqsTfGwjec8JO2y4LHy/P
N5PYmlImP/+mDe+RJIqVuEH/V9qHpNXR5ShIKnZH9824TpYzxOP6tSQDGAGgLc49
jvDMUqyofYkcfmFnOu8TRdfpHdPFEdVWHQJhlDZq649P7m2DmnavFdSZSNfW6Rr2
DnS8kK7ygQugcAMLXL6lF69N1bNJK2xH4yVQjNpKQj8dsJPH8Z2pYc6D529WQDId
SqQOPsMXwaXO8uGMJcSm+9h842E+c7Z/LwdhHJT00m8ZRI574oElwdbyQ1RZDsUz
ZQ+vXDWv59A1P6FEOXxxd3ZTXJc0nu2qM5y9e1k+79nOWsbCGPRHoLF7vc5pujTy
kY39Xlcm4F0pp45rGNTKsOK2uttXvp2hvMD2wKhh1kWqVI7R6AE4vyasE5gGfymO
yaVdmfVZVtGZT0/AVptNLBa7aH6W6l9In8dpIna+CqxWETDQcXhdtzIsm46V80K5
ltZbO98OvyUEJlkg7P/UMpBvQ1OuVTR8rCS0rlg5oaQKAMCH3xaX7gbF1bDEZr6l
z+U+X2dOfeidVLGmaXQFbSNInVyMh34VNAYc+BJSofrU47pMlXa2vaqVRVQuUx98
Q+Ekt0uEmZ6ozPTDResc6fOCh7Gg94fwhi9AeXJo3FyOc0wWnrezS5cjxwDdJWF5
blaEt1Vx86saqY9Z5hATAQD1u14kbYucuFpnhxUuPwM+OAPOarGzCZIArEWf+cmR
CBKhB6BGndIdIdmIAn41PsuckahfWAx0+nmAn152HRqHycZHbh2DDR1cj6AM1YSW
2RGMPY7aJsy64MMd88b30jUzvPOtz1Rq3NCL5KyBvs5slM1xchggtj+PlBmaBpMZ
5+qeoemhhPMKFAASqNszvwp7LOtTEP/KkamgX3kJboScx3Cxr5uvzeGRbxw+KT40
tji356/XkrFNlQyWGQTKN4SKhlWSeAGdQr9+d+jHgaq++GwABsvo/vy3pfYXxKpC
zwCgd+jnIvh7a0k7Kv+RfZ5EKtzbTNHjVaNOh2Gku+U+JcqeXvjJ+lMyT9ZNcOdJ
YL6gEhbAjvwwvkS+7+Z7JPWzVnlKVFFx43SFx25WHUlTgLeNusJr4EFaqqp2wOUi
T9FlKeZj3bSfWbHpSjf6nf0P9A0e/9ADFzYkwkJsWIWQjk9Q85HlHuVT5HWWgDL/
fR6NPn0CszYlnGa7bLNf3dof3W3iQxjaiV0N8VLXvHQxd3MeZNcrpa0N2HWppeg5
e6WXkAu2nd/SV0tknINTteyQ2sEtrr6qDoxyfFngjb4L66SvfMOObHxlCb2cm5Sr
sAgSQroI6vxwfTwBntM5lbb5PW2IKmnjeAILbb1ehZRPb3C+C5rokFCxZp8Jxhdb
AE8ihXUwv3gsiCDysDz3xt8Z0Ks1Q+jnpeKoM/Hokb7Zgm1fw93R3vrjy8d+OdsD
AzBvVLukYUVQkK1EEqvI4iLYSgUeCyc0LHg/jKJLS73aYmsd4zCjE2/v0cMPKOC/
SnUjObSayRvSc3By6YTK31rs1YAUnXF7+2X676WIUeUbjfFfpo282UX03BiKgBw9
siY3iPKWfBGxq1wkL8mAFVlpbvWuNEds06K+uDGTUN2tQHf/Brqf31CxUGMTh+yD
1rjmoZxr2oMt64bcbPmH8lgaHKSZAYTTfaDvi01DwA9ohQ45RuZj/hKlRC1gFAqX
rrs/leRRxN/Xs9yaqaokJd5ALY3cJSQpxsdF48hz1DlqoxvKoTUzj5LymjRgy17H
kAE0mzjJ54y7mU0AmbCFXBqjGm8UABIst1IzjNeQkCYlCIaZYUtdeb1d7y2vV99+
HiYQq0sOWse49S0Z5JDxEIYrjkCcD4ABeBIdWtPA/KmF9Hf7M/oGyN8pGviKIO3w
XFd+jzqmH8STVAEXs/PAS9hE3qLcdVrrh0gLIhiOwxkuS9sQHTkdn5EjdCe70CCm
uIQZ3CjwMQLURnTEt06jyGZFz/wkd4ZGl5XDgVnK6GxrgsYVeiDIOwo0PCUvRiTb
zydtfmQZEorLeMSklcM/cg5VAlxrqJisZUiIGc640X9vn5cfZCSNzLcvW1fV1TDu
gNFHAgGuAD9cZJ4iFE2+zsFGUx3wjkVSZxnz9Aq5/n9j2mmbCFhlGRApsvpMU77/
jZVQzTS5hsbChZlpcINTDU+wKKWKdLMEkclBrxBBpKwwZbFS74UYfp0ttX+c1P1j
H2KVg6nNkUnJ2SpRPKNeE3OjfY2QmuGbt+DtUM9G58FZpST8MQ43hbGpscILL3e3
ZK5uqNLPJiRCJe7HL54eXinZSFhvkb0Yl1n6eBuX8V/aG61vO3oLsyyDENaK5ZRO
yfb9BbIWubKSb6RaRaB2K6pPG/NSFnnixXJE7/uiV8wRyqAJd0PdoLY+RezmAnLU
DTbUVwmqN/t7zC5cpzLCJ5KvfcFZmNYwQa+XnhDJBCDpEn39Pq0ZLlLKh1Ghy05Q
XMBq18LtZ+iLZ3CRLqrcCGFW5euwOp4jRsLNMYExNn4x4p+K8x2VIJsYX+hldS/n
kRemcSptIP3BmWupVTkchp8UPSsJp5LWod/yFBp5Rgtm1xa9iaMfyayca+TqheVE
HQ5DOZY0yCZPPoNmy95eA21gZI4w/JMLvNeZcvadqp1AF9S680JgvQCpTHRc+yyx
Zki0UvZqDK6YUhe+muHOJ2zIZ3BIS9nMo00Dca/EMw2eFExIG2WnwU/+O+R3TTXt
MBHrN6L9KZnP3jJ0rrO8BPS98ulBsIEA5Kn/mI2rGU7E4kgYpU9dYYsaGcD0gjgE
gDNrhht0F9O+As+ql0STkEfXwRhcOapq+OT+ecEgRAnlmPVzZio3xBKSmf6ewbNj
BYRwu1atG5/mJJrJwxQ+2mL/CmSdQR2xyLNjWCeNj8yaPpx8Nnb4MMzndXejLJWU
5V3dO1pQ6v9lnvMIT9x8qdNklsZv3yyx7k5Oi9Sq2mMq1pXMm2RQqsuioLU1fLYv
f3a8Cceb7iNpIqe5oWfplUpAtNYJ/OF0404qRQwVxFbKkiwWtWSMdE45UbubCAlA
ANi1W2+XgypLFGtd9XuokpqgCq4cQ17kB0tFz/80DUv6LYgcckWPzZkum833Upl3
pR75+dpywCgi+nuhWQK7To24Me0fqVhHerNwO1cdYVkfx0BV0RuO0sxOx58zXJkL
appa2gL6b0K5FFl3nV06HjoxDf97Y8Pp43Gl9gBnTx80pcqlLuVO3aVSHfnN+LII
JaZrnEA7QNiiqSlLZ3as9dbwXVb3//qTM0aBiiYzJZV85lRZEKuge2rZqEYrDtKH
GA54i9TnPxJdZeuBqIM22Z2xtEtr3cUlLkyc9fvzVlJNh1mjBUt9pUnR+tHozKKO
87zoOJWWiz/wnohT9G2IS+xm5AJFqGLCsxH9uPPaXxIjqecnOiWA/7PrZ6EbVR1c
OVy3q3Eehtw4xSJVM4mGzlj4J7Wgxx3e26r5A52Iv0F0RlK33/EcFPyvYWrlPDML
7qWJOn9xffAtjWpSDkk2UTFrNjox/V01eoYKRTessZxlxODFb8YDGEvkldCrS+ni
Vp4yq8Bbx/5ZUdvp2sGoyH6p6XR+F5kgB3fqWivZ9SNMSgmNxXcHmjVedLVhhdAE
RMenUtOQpVjEaBJzCoyZGhZhbMbCTrv6x/a/mpIzvGkPqYh+7fRV60EK1+GxWqBg
mhjSWv8S/15Muake4DtQJ2R6i5lNRati83JPXg0Ftco1M5lkVBkZ4CBYme9jw/it
AfF1YglZ/ZS1eORPiFkkDtENapl9UZESTD8d3jZuRSE+vd+dVm0D0UbTRvCZ6jAZ
g5X/LxoFbEXkLxVjMEW0pVFFHE7Tznb66/PtaV3bG+4Tt8HOouF2+011U6v/WqMO
Oei2x39Uu9ZvMk6QHScBwNLTCyLb5d3uerKFaoBjIANIrPqZ5X0xqK2uryMn43I2
mSfJoZEWxmX8Zdo2qonoF4NGiw+7MOBqZwuxi5rMD+v2RUy/PRCSC7p3e3ohvqhx
XkWIbAo2Dyf7910NwikBE6rrXVsTDwXJYxs1mqOyJWkQigHxau3kHScACy0ZpjhF
sDwKZ1kNT6F1s/t2vzh0cX1vgObV2qjwFsQKCzJah8tPCmkryUM8/u6gu2V4jCVk
XDUTXccRb12M2if7Dc7+3b8wrV8m9+NWkaTL0onPEaibdM6aJAmUlB62v12Xd4RH
0LdGIYWyL5TQg16Kt4GlrZMM0T5tfAaSO1d4suYCdeQBNohv3VP5mtVA7AN8Tpgp
CmjjQmcZ7L1ukDKPCLhowVsEfwsMJvnQ0Py74rGb3Xw6NBCwCZQT9DW9II8mGGzm
et9OiBvb7HulYqExDlgVVJRvfnucYJAXASwSWVt/OM+v1V5WOssvUEYffB7FZPd2
2KRvAmvlkW/VkQ5tKHE7yqWAkNo69FddrzcOzCuw5CCrhLwtOPVjfdtYzgZyfB6g
kjIVuOijlyCdEtZcIg9KMgc3ib+sG21dVFeG+0nyRr9nqVMQLZeYmx7PbZYjL7hv
kad0ZO0W2Bcy90tPqCiCdhDpCpAspi9TzfO8W2q8jrC2EhuGljSwnxoE/Yxm4BRw
uAntqEroOmD+QjLYGuK5v+ldhfvRvNpku+qpEKT15X46Uui2PpEoShIFepyISGBQ
qdGJn6pabP+0Z3+pgD7n7gVAxRwGkdyjdswKHrGsNfKdTphx/u5cBtFyMUuU8VLk
J7H+RVTcnnMEcH/qBi1c+U7gsc9dhguYqsCSUM5qbG++JtvVPkaVniUVp0ZRBsFQ
NYYQzj40acMJZ8SAPjUZg8lrmaiwsCkqy7PejacgAzgv6+kkM327Z/38uoYLi1lE
hltOvNyBSJLI8tmPtpJLNywj4KXydRfGAx89i8VWA4K89YRo7s6Ah+S7Jnu1IAwE
6WPmc5+Z7lzLpTHDVJCrJmLKV8pOdlyFjs7JxEbpqpIhVKLFzfVyYh2aJlJ8pmNG
RWG7hOsqQpM/bSkqW38UVOiZSSETgQgyaJF+tqqjYwcPgF7/4H5yXgAHOVRPg3Dr
Gq6mlpDgNV5awt/ncpSNS4zZ3WZPSqBFHdkMjX4iw36rGUBTjzCAZTNIktvUZxON
1pUHi4WqKYCYQKPCf/FTEAzuWJpQxtWqZbAN2rJnV8/3s/vMxTux+eJ3ospkDU3t
MEGVOKv3Ixz115byVAhktcaT7NRkPGebb9JZq4I8H9q1vWmyWJiNW0eaQibaoc1A
B80olVgQhWfEbtOYU5mfm/SQv9PsFKM1R9paUQx/yoirhmXFJq0yshKodGqtrjop
eHueUnv+C2gN7Coj8Q7Z9Qmzz/hIChsk1hQ5cpXSmRlldMIe+pa2n7EH/ZVzU1AQ
L9Mo4rKkYQR15f6Yylbeq4iGvb/CFS7r63ny+I5DUEeO6AjzgS9Droiu1pRr5uJM
rpm1TsPOdS6ymohQsamY6MmsVWAb5V66NJGrsm6vaHsos6Akx9TUNVE6KlcPeqpV
0wmOLKdMPcH+nN9Z0bWVq7J22KkWhgeTWFXQzDIJeJEI4BkjbLhuBElXVGsmHHUV
WzrxQ1MIJL0jsNUDffzVK05HYiGcFPeGWLBHvQWcL8zzySjyKrgXLO3SwkOQ0upn
bsEdcZnitOygEEFyt9yzOgSxtkBUxF2EdbmY6awhSXGf41G96HOoG6RniPto6ZqM
g+PxTFux6U8ggJA2jrAh0f3SnpuOrT2BdFu8mWj7F1yT600qL62m/cUyKWr6A+yx
90CIjTKklUzcJLUKRMEWILeciwG0OEy+YNyd02DQMsXfEBpe+Cb1IO1Ehp/w02hP
CQTntsfz8EWLsli+cbsjHnE3fWXlBAdwWY2tE9IPtlKAklKFUpDBxhP6OVTQKaOG
otY4O9d2Wc95s4UhScVbc8Mlvqf7g+vLMspcT9QLXbqeg/SyIsuUeWZXFJYrtycS
Km2HKoZLovjQK+HSCnErIyauf8p8sFtada2e7TkCo0DgYC7czbKn05VLCQ1x3DfF
QpjyZW9vJWnZ7mNnvXx4foMeMO5vxKgs/wfdX2/zPwb0WYGvfS4yct1lyOsSy1+9
ZVZUGFxmUEURQrzADTgZbrQsLwmg2+1ZNCHeyOG28zHHtnnUvecr5NngDB8SOnwX
uXQ+QHzEyRG0gtL0mJGwLBK8m+OvkX1QB3hT9OHgQMjnTUGXiVTR/GEFx4fIP9n8
5G1QaXdgQtDDp+xyfkEqqJ3CL6vHqfnfepaljsNKp0W2So5rn/3TcHLRxAsykQWd
GGS2PZisvGDCC3eo4TEBqcI9mTGEEaQvUmqF4Qa3mBJcYBfg7B3o6hNM1TcsT6cz
XnwOOfHM+W60Im2Yx8OcrFxeLGH293LEXZRZ2nTSfOGcaaSwlOAKi+Dq9Zc2qUlV
P81ma253oC4PNEG6nhTWMuf8RiDMpZRmM9nFfqS7XkgW3ZIktffmQLuqpIj+b3Ec
FBM+iuU2tpPDnrmKSsycPmUrvdZ8fqExvUPusDOvXlnABWYdX+CFdv3LHTNlNd+c
bZpG9h3aYn21MttZh9dYF5DQFbu1pIZKPl6C0Gxu7P0LGgCEbeDKmz3irMzf4Q5F
MWG2jSwnR7plS2YbWGUVQR2/Ck1FkRUOjUW4hbHQqw8dqah1Vmj445vpRns4DAdN
naDD82hJFEbpFGvSEKtJHMWDOOT3S3b+B7N/pXSIO56tRkXfJkkl7edwE1AxuEZJ
EdAHzCAFtrODH4SCw70R3YYyb/iyBOY12DUa93yOPcoFSSUxpS1g9Fo+YNfQaowR
ZtgkOw/ix1s1OR75EVFLS0Ph5Y5wXJfX1MKRt/djgfAOoHMROXBJ7VxTc3KaSirJ
jX2tSKQbmw7D5oRJonRgQXxsUqdTM6z0y2TSNNGR8nc+yo5yJqvywe2V5Peuwfo9
2o8VFzsmBxEfNd9oyxsJqOkZ3jwxMikRMnBa2out0MuGc+uq27Roei7hPxKKYVKx
cq1UlWSdQ9aMWvrAOjgpCzUfibbSUoJjqnrFBtUdoSmsTfDUBr8bBHqwXxawFY9v
y2M0F+n+qZOhj3X5mW1Sqgwpm2t4oQbXqOCTp4l0rAGxKwop6Gk2l3dNZGX3niMR
CkprRQJKl11A3+h/tNjsAXxlXNFWaX3i6lJRKyG5lSA679yyQe6LkiRC1ikd1YOP
U+LI/pqnhrBik8qV9E5LcO3Z4pHW9rziZsMuqWqXawbVt3jFkm0Qp5Puqso0PrCB
jWKGgEd7tbeQtEbSZFOg5Qni6zuhq78THxXz0/Jx3qlwxOhTqCBgfYWKLip8tACe
EgdUD/ZaiQo4evCCwApzwk/Mf6WBCyMbI8HldQP0xuhNwcosXC5dO1UJOxl7aKEN
6Wpg9466/vRKkhHg8s0JYp0vwVIaEcvADPynj5nr1BhPsdhinsdn8Q23W2ep5kE/
Lpi5fhByPiO5S/SXnZ7INTrVPpEIZpS+5kJ8JBibKKxMDrfXTK0/xClLnyJpoqWL
v3FjYY4CIwfEqILocU8MN7g+4kwkc+6FLwARNTj9X0wJN3PVEvphiP+cVx74EUIi
vVT522S1v39l4ft+HauHAMcLjjdDhF1Gz9tC3sOduaPGnuB+CrOhO3L7Oe+hkOPF
ZPjmsqNZFRsVeMdhyp9wgWCJkwjU8wZCusxbSI59FCmT3q92+Jhfckr/zPZdhEhC
gKjc+Rb1dRVvIlCotNGSliuLG0ceZ1Pz2ZQDR7xR6iJ8A+0Ez7M8HqGtoKa32A5E
w7zNdFtdqde9XeObWBJegFs9FI0kF14LGgUzBF0D7yAkrBL/sqAodt8D+2IQ6WGH
`protect END_PROTECTED
