`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5+XLoGxb5m3B4x2d46FOSABwrEtASTupa9hcsevE+rir0rTUGoZ3Gf++sf4g3JY
jQxaqvWQXoA03MppEvwdQe43LucwmBVBbq//JkQ4yxBsEjikTe8CWzY/dQi04NQo
SJbvNvOBB8OuatJQGqrHTzLyiDjuCqYxXT3QtW+Aw+fdLl9I5nbGf2cTKc4QPNMS
8p21kZFFIJ25eg1bRCxs5JMRkg+Fm5MbJxn+W5gRVUxWbTkTEpTsB4y7lnD/Vll4
C1yePB89qJEn4SjXpyBPnvcptkMRaWa88nu7+PuSkUSwNPPId2IVojh0VYytSJcc
27EHYsrq2kOPEYSe1Aiip869jknbh4r/SlTV8TCzlw9DaGVbxXrJj3vg7BJB6XS5
+6xqivywZppTDGBcljhA8I9uRz1UqQS82md/QLMXTNc2qavS21h6sxzMkvGSpGOH
XYQtwvwZpYB9s3xHh0ocASr4+JH7sAo3GBWljk0qAhhhvgFj8VV6CngjD8M8hWNL
jpNTXPQuVtmqScRzQyXvc1rCKmgQHGArjTYg3BdGN9rMNuHLxX4pWnD7oQwNEBWn
Zt2LdNTw4ASxfvzIea5S2eyscd0Ev3IDmPyQockbJfEiLHl+TdDg9Dv/osw/37bi
W5f0HSaocud8tKEgPKEVIiIwT/gc99vde7lNKmKf7GJveDtu/HfmAhp98GMtRDeN
Rt1rNrRZg9mRAXMiVkpspEOI+o9Uw7u41Tq6b+ySA0J5IR1U88NJecjh+7u3SmyC
YpjMMvXoKc85AMB2j3aK69yJp6W2hMLGa28t+vBjw8VnFcIOH52HEeqt8EWeuoFO
9hEtg4K0l4ReeisW99SuyoDHBIGDNx57WDdIShTMjD3ki6oV9b9rYnAio4kLole7
0pwAd8qusKrKIcS7kxpE4rl0QmLEvLBJYwHuqK+QfKvCt5niDVyPaK6tUdhjIxtG
Cxp88CQ6NYSU2Fts2nb+uKGjGCLiymqVL87z/S8Pgagvw/43AISpeoALJI3eIp1v
Q2eunf6/FiiR9fmDtxobVv+fseH0br+LrGGNdfKGosD04ejKlVo7i2A8b8iC2+5r
ANvZZ5YrNPj6Dccwol+7NmKuhfZ6AZgLYNQm/SBe1Q9ISC5yxeOtU1qPz+KpplzE
LYSYuNHeshZGJ4OhOT6TE9R7ElZIKKW7lEjDospV9TTzFDY28cFq34jpErZ2khsj
3OTjC4BUPGQ7ZYq9N2DxTgB/I/268SDQysIHD4vVZhvjBhafuRcwRxXo7HEA2wy1
7bgeYbHDAzDPioNnrFfsHybYRMg6osLKX81hhrG83tdiiTmo2/17+n9BDW46DNEU
gkL8Yf4nKEcNJWWFeZMpBGBmjHpokCS+a7tLL/umoszqgiFBXnCNGuszhHFkH4Zs
YLZsTda0uEIts0M23gwujE95OUP5fC3jCWuC0fM6hSMyX8l6n5HzdDRoynon6yif
OKKP30V5FiFN9BqgSDvIF4G/x7v8ocKK2pEXqY0yL09dsfMecDplX5/zug8GZ0tj
pQ0jbTX5ifFzJV7CnFseRl9pG+cc0l29drKz9/W20dhUUd+DrtrmlnHvFcDtlgbj
iPN6urZM7wJMcbeVoOMt7OSJkeN8KNJnOVO3H8ujkfRnl/caL3UHrmiD9QozSii/
CyCbIWTZtrIwU+udHWRFpZADQdnbOIKxEqpkI7yw4yFe2sCxPnylnwUr4vQfer/S
C8qJoyA5oakeS32NPsTIl7qRCMTxcKAWDbl641Fc/oq/EH+2p7Z/tCTu2enPXgmw
AJbtjhGtc5K85C/DBK0wulX2+2um69FJk1LuzgGEbcnFjmjzRApAw5m0as7+Xhh2
XyZQ0k+c4YQ1HPHbh5bz2nETwGxGFtjOGJgBBmECZwZ6Sn+eojhpAvfmY2hm1Oqk
7HDre/096GdAAy7q0G8ov9assg9rkSsb82t2ILJDl3TCzj2dpejZaB38XE5e9Ix6
sI0zxfxiTP+vl9ejbAAxaQpb3gCTAGKgd2rAeKOJ1cB7861SB/KEGMSOIN4q4gDE
bIQLS1lzu3NzBVwDzEDF1ENsp9c2wStumSZ4cm8BH7QQvGGkzMdQvT2z4hJow3fy
mHwoT/y6urtqQd/a7SP172ywb2ytWIJBWJiHw7PdFbWgnRfkLwrIS5siTn+sRFFF
8/7WtlJg1gXXwsE8Boc7kGIEV84ieVhcooGTb6pb17BqNiLfh4JlOcAGKVBELSfe
gLf9gG5SfBxPMc9+tUO1cLW9pLmbsaqFSy1oP9pQzJvmER+BXSTbxGs3wfCLsAAF
+euOz9VTqi2ZU/VCNhEDMkudOqaLBhSLCNC/tfqCrgkDhaaGMsxt0KUT9wfppTFh
TAXFjPv8BDimkMnH8Zw0FA2wU/xKipXszGihyhVdUM2cwmuhU7A3BoyXW5HTlweK
f0nLZ2cntN3Lm2zOEpGkBljUjE77L7SeDhaibHZ88YKjEipJWntUMahXAmgt+hJ1
+2/u9qTqWDPRmKq4Hi8A6RxkhFNvEFg4YOSqe9mUYZiVRmJ7TNTLZiU//RNsq5/s
C6Nv1FF1RjlXOTAFtO6kUsCEA8hVZC0w2jXBngpyRnm9cRe1htN2TGnPDoKxi67J
hGWgLfNXL6RIUcAqGu+mj78GA/XLNoXdj03qU1ajT5gQIfVWChZRFy2UY8H+MPql
I0kw8xRTW7KfPLH2P/gxidjnTqYjKeGKFKZBp6xcHHVEaWcAau04J1xi9g676+3x
dDd4XlIhXj++2ht8qo0dXxg720aaH3t5X/IT44df0sNDPdT8Iy19bfnF3uUvpOYz
E1Ww7cIarlsLyO0YULMQ2knJgITXBh+NHor5CQRjOA67APyAs8eodoZnk013bH3L
mlFMYALqJihca1eDTw4e2DfXaJawi9TBUujswv9HLVSq/xl5bbtNC83kZNM6AeNT
fMYarUg0dUh0tDlNQ25zibfkX62L+2Em4WboOj7d4q0qe0Hf3MvXDbuPc1frsQ9Q
4MwqVQpe88YoA4AA3tik0+SA9vf8tMKo/IQFvvtkSEqIBbrs7eRqoxZoFtNz72SY
C7MU+UV/vj6B+BsRqJQCOIXL/2PiwTGROrm1Q0n7Cu3SEKZZ8HFIZm353EuCJqKb
GC6dKQlZaoiap6dlqiGsOLlPEeHLYIvpJSu2xfQh8Wia4ocBVyfe+dESMQQZ4NjC
RxXjd63d0DkZNJ/siFdjy4nDqdaTJ5jZp7Np3AGABVJMEUX1Ib4aa6xgouh55iwb
8+sjPr2bFqCts983NSrWhupyBTanAVWQIAl+I9DttUjVksNNGF+90Mm3Uz8P2EB9
LLNwCwp0ORNf0JbHM/DoBm8QneX++VbWqQr/r0LO2u09JaUI2UY1LLuujo2N2qAx
MblR7JRVDGIpTyxoafZMk8fhj086dMbdVkyTNl/FYpuEPYZZPHDCqvoTH51vOxAS
LMakfD8y6GJKe281COdX+MonyitFilLU55C7P13YEJxL2kRIAQ+DVHInI9YFYTaU
LwRnazoueNiVQZiymSkeNfJhsKlWgrW8Lyjvnja9ZbLVfauHImS9OKh0FpSTvFRg
ZkS6ybDYiq3Vl7j9iXy2x98DI11Te6YP529bmpiTlDbbUvSaQ0AOM9SMcLV9ncaX
csv+JYmgiKefG0I35jYtqvzW6twVld562yFtXK9Lznh5JJhdBVR3TF8a7/LZXCb2
HSDCj0VFmKFrMoLWYl6JzilWPuYMM5BoTSVdy+gBNy1gYEcBUSGvepCCkadmtq1P
0EBunuJTesSJZSrBe3yKE3UJQYzM8ar5yuX2TqaAu79E50VFnwRzRbi3YtGruRyA
Z0sexEHCfneBCHSfav17dJ8Y1vYVNgtrMJmP0jsqUem6pK2M6oowrcvZsBG6Nucz
8xJL/0Vig42b2zHRHJqtcTHLmNxbJr6MBJaiDjgO8GziXjBXSUhcg//b0eIAqL8X
trJeR+2ug0HfYKxfItlLNKGUWPLdPcMDxN7Y7DoQKBNtWaUOOmuh6jOln8oIwrVT
GJwX7sh/5StOnjey63DDmX/CylqbmArBNCx3mvk6JCRGQ6JHQQkhAc0pxggvcTVh
gEx+H4XS18JChnHLD/9sDy+p0pzW9fhvKv/kBbuTgw4ncBaalKA1FSNzL8ArcxPh
mmpZHdE/JqJq7qUOtYW7Ep4r/ipmuQfyQKVUVARkPqHDsaBtw7Ku2ntk7NqBMyRO
AvxL+8Xlt6zcbwhDjaf3hm4atYfOiw+remrXz5Qc+dN2YkKQke/Xcfa7hbjKYsje
huaSftVWW7yrgdVfi2zjuknZi7g2Xftkhg7/azlDj1o7pOIp3kXw5/GfORko2sGc
qD0shjMPLih2nMmvV72LaYkN9/fWXzQR+wEZ1wbJYWQ=
`protect END_PROTECTED
