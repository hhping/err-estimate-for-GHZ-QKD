`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLWKRfDaa+uXQ7rD1gd41yL5/r2uGuhn99KWMBRV9zKo2QwunFJ6d1bgsLA+brh8
SQVXXNTGOk2O5m4CXh8hjVy3AmmdhJOJAU4SAHNMq6hwZbGczORm2xl+LGnJg/aa
jZ0wXDSwoVvVt+yipL+mrKi/tNuWPtqnfUlwrDoQ1qlTpwd30Mju9c7K8wNiMYkd
ofQiGiobTcs+8gZixqguHLSVFIPEmfF5L+HqkAPLx7NvaUdJYlGLlojS6Hf1nIuL
JOPodkIR1aT26dRJRjFmEE5Wdeayb0ec1pJ5aV23N6bTM/VSU/PolL3JoRHTqtFT
mEf+DhhX56NkfirrVrdov7DmmVpQYzLVNzu78pxj58nsjheqXvJoY5T4b+LxQ36S
T1N+rgkrqfT1oOJTGAdTDw68V6jmjECjMUVdawWcP0Jc8rkxfE6rdh3JNGWRuiTA
gnrLau7wv9swV2ko8EpOh4G7/9TPHk0/UxRjpr7UtfvmB/QMo7oAwbUCsTFfML9w
fmMGXmPkVDKOt06ca35SWhcnVMtiZx+QOUP9O3Sl3B4=
`protect END_PROTECTED
