`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bs5UwQ0T1Gu1ky3qLk/1lv2DVcXUgyII5Bm8kV451qqoot4J08g5fev5NEacXQMi
ck18pQsGu8/DPtl3EpAlMUVAroLNqs1PB9YlrX6L+rU1uLoRm246M6GZaaV/LYJP
LPGR0qjqVIAgDx8FAcgSbUgcdIKwbaYV8SYnoTpPnuk5UtMOaLaVLLwwls5fi3Fz
LLMXPWRvMYRAcxKYJDADxF9B6v4KwoDpjJ80NbfHdw89brGgqwzoLZjxT1HEkfWx
+gZLtPLrtRKOjB3BRrJ+6BvH6D+b2LQKtxX0C5mN1PDaOghCwZI0JykZF+xBQtzR
c7fZnKYNA32JwVAEzvaKgv56sFNVcGdKLW6tJCbTEiHW5QrcTyzeliAYSGW1Rzje
wRu7DwCU03Dd0KJ/p04dlHQt7AGxZ2UQD44b5WaMyCQu+HC4E6xVts3pyYYpaDfs
fwTO9c/Ew1F2IhqudRyenUV42BLa5Fx87H6B3l1sWx3N65V1nNP7t3zEKTgDVodg
IncyaY35WbDp08EHrh7gM4jKmCVgdlx9AUkXIrZhOYFMZoMXsibV674FZVphd+h5
HvSNIR6H2Og3K7Q1n/9AhuxvIWBrJ+R8z5JdjuBmm7JFO6Zs01Co8uT2MNlrprpD
IxMPgO4XJix35MABcljO+P3lQqEGKql7QGqLPN2xk6g4adPFZ7D3Lr4+Xr4AQouO
SiCP8sPMplsORyLaaHAeIuod2uWdc5vuPYRky1QYt/99vvDIHfhmx5Z2HffNMc9p
BJOJ/Cl+IyaXgV4bvCFkcKGU8yskhf+IUMvv/tgIj+s=
`protect END_PROTECTED
