`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fY0j3c1mNmnVMck7UpLSDQexSsw5DFIFATA6TxHRp57A4yfOXi8urpllnBKMIYVe
jl0ZSzqUOZRgmvUsJSPMvZ6GJNif4YY2LwcUk259NH7mnXdF0DIfI6zdtRAz/pWz
qp+8351phz8I/qA8qvCe12IxlLdLAa4l51dQomKnLb2zdjYzApjzXBHWwxz0hO/K
MCa0B7JhHDQnwJHN1n+9IaUtI6IjOzNtUYqIVWzilJG5qp5TSKy8q5fUaCk9+Qeo
TBMnLTbv2wArUTsqssD2Nm4ZCoj12l0is8ZCWNkm/GYMKTmfIVIf9ppQyWOo7EpJ
w1+taqZxwpOjpeR3rN5G6hIxE1Jn4zsxzx53HWUd/pw5PE3cpHLZnCT38kpH75bI
EjKtTnw2Gc5Yd4/h85PQI13IngSfZ/SyYB8T66igr6FpTM9cSBYqlLe6N/LIHgRH
6xohOSRzxeUHbeNBTfgcWtoJsUOPNn40J85azqJr9QCqmO1007plxqflzKmmTQcA
lWEeiCLy5omOplyZRBqfDM8LaIB7159+ikomnrJZpF2tKJfcu/Hc7FsvW8qskjLf
ybOvoY6wA7goGu5T9UlsWJHE3VHgiDZ1M09ORTd+l7Wmj7a56KY9jJjtkoMxS2sE
h4NFjgFZheRGEQrJU81ECxwuj/wHW8BHJmONADsX71bvI7mP3ys4bONyxNrZr1/k
Zwkai44PAq7io2JaO5qfzrRcLPJrLGR1PHkE1DsaW9MkZ5dTuIETBPjv/bQhEm4o
tEDntKV0wfAaIBXjD2CE1nA0Td+Bf7p2tGm0O8LSnQyPKOtkbUuD4KUdjIhgX2k1
a2BAT6VtH/2VPZbPjqf6KTi0OvwS7uxbOxyDiBV5TiLnSIzhxwrFiluJu/GfALkx
gAt9wXhF8xMJyDdhV+0hgdJ1V0qLwrjOkVkFGXNfOUMzgLWsaYAm2D1MoGRI+pKD
WGPVPuR6Zo/8rdCfSg9oCLAAc3J6JFAlYRJAqDU85qLFXscTBoHJ/94LBS+tmKhM
IyP5k6LUdnPtQ0FlbLruSEFYT0OUuKd+4tgacJ6zRSPvH6IJANLBpthaZdxh4+Yg
CZ7tdP7VWpSNHNra5b+ECWJZqQusz/WSSZVMpPt/qX+WtYOLrU9Cl1RDoHAwfr/2
wmAt+8xNO++gGQUmGjAV3rSyuCj0T9STjT4Vo225ut2EmV9H4xUglMFKomvXmWtp
nzWAZecExpS0bY33mxTHLXMZfoOXWeuWqcsi/mYlk+ELjHBOsTpue6jruvSQ1BPh
nPwVKZCCGZj4Nw0NYTlqH/X+Shnl79gh7tORRCjY0rmm/RDFiMDNIy3fK4ANz0RL
szYe0jCGkfdiA2WukUpnOVeob7y1hQa45fK2mYc2O3pnRvKk8M3d9p8K1N48alk9
OUqCrFt+5W8Ku7X+tHkK6uDSlA5YzqZq/JiUrv39NKolJcoyXcnZQZZ8bxCKjWrS
jbgd2Au0ohFoCKYwadRjCdU8Na6GTxV37/EuOEyQ/dg4YXxugfCNwrmh8agvVDLX
TeA2UVx3SCXNgx7fR5CXoVjBdq3tMDsNzqh+Y0iZ9WUcA/3r97IHS/D7NZjPo3c+
3HSIkOTtYMcQf7kOjol/ndlQD77TbbDVYZTDQC48r+EOL0jB2SJmvzk4YzpwgVEj
3EfnIRDr1S+UuptPm8JCe78n9wRByCMbh5jkBAiIrc2JkZpt9k52vrG2RmGY3hah
N0VTLhfkHhecTcK467HD2wq8JUA9R5tHHvO/USKsFyiGAk3Ubr1xyN2QiB7vqdrm
0PKRLB+w/a1UrfU1RdANPVlkCE8SH/96pDqYYpTDmZWbWCg/UyYcHGv4KbcrXOSC
mFQqoRW5kuTKY2Jqr5UmWs+JH2G3YVj9ZBSAJgfzPsL4xDU0Rz5MsjWZl/IR7FX6
pvNjFJO4QCxNJVX6QQycgjNgx73ZsFKiDpkDs7L/PrXVS/5H+zvV1j64NCgm/MtA
1dja13kdqN1hBObk4qXD8s009uvTwUrWRpLFO7qFTaqI3V7uUWEFgjqEvGJvFy1i
2qMfBnojj/akbLHqatXEa3JnvtGKlU0fl8OydSdY4BvA2vl1LL5ImNaNWNRrLAC7
kpuLCuBkxoj7fBKr8PR75Jd5/eD3Nxb4VnDh4Z++ybwWlzO+t/z/7U6CpfVNPDki
14K2gym2nSsvzT+MiYoyhStUVHRKkOhTQuy4SGLCfUuQS12CthNVK70QbvaCRUXx
gN/KiZuE2CTxhXybHMEzf88YEr3BNAdr9UmefxYBOqiiSCAFXg7AcmJGzAwUsQ6n
XbWrfrGybvIzcXPFxoXOTi1PXFdY25ghBofky5yEyzoELyi0Ic92R2vpqBpOoqe4
iDPeINn65/bKwnimjiPe0hfO83h/6sAcHe0662HRjeLcSP5yhUr77+27tNVNWG8v
GAKmfxIdSWhhezCmTsx4A6LNzysGlyzTbIOlq4f539RgVIyB2NxCL3QltO0397cC
DsIHTdOaW/d93woV3/rFUya85rIzcRcYV7B7CynXmS23KZWEj9BDe9/mVNFqQsAq
URKvv8kF/hXsLI7ZmLxwKWo2K2zz4noGph26TmrmDdM45+Ds+kUgHIZ1Gx/xxjUr
d1zKG3Ha/v97sa6bDY5YkFuRM2HZyC34bXyJXVW2yJglGZadTatgMwpqQU2o7lpB
bHRSg4RxpGLqCxE4Y/25eFJ23Lo6sYQTH3c1N58QDi0cwQaPh9Os8QzAlQnyAbFR
+iahj9nKW9V6Z4mVdpKYl4KhQSNVaSsScvLIzGo3IGIVAsW3iDhlJ9RaZX+jIaFE
jTmOPWmHtu9NeZzp43UQ5kql9JM0cu1ZcArm3iNT/R/FcvVV/b+GyMvVTdgdedEN
mjZ74Omr95q2bFKqVla7uB9okKcokTppS/0BfIe2ci4BjPocKvIHuQ/eeXSQ2I5g
AmdqJS3u2xDzgeBUjXGU6A==
`protect END_PROTECTED
