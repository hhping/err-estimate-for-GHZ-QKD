`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KWQBjHAXy51/yhwg9jdNCHdmLi3iMvsUScf5p3whyMzsmwF+v8epD22k45ZBWcoX
MeL0s+hAxJyvPvXiQQ7zqJCkf/b6Xhn38Lt1KW6cjQIipvq9gao12FNxVPnR7aTf
/s8m/buOnBPYlGo0GpXaOo1/sopVZjVV5+zpB+OH72qg5gsXktdXTBwsOzB3Atbr
3dfhVwzeBEO03KZ3pp+8rIsjMraWbIbJEB1Cukom/jOCNvd9ogEIa38V76y3Z9ze
yXUhklDV/gDMeQyOGD/74bifI8PbB+WfLMuVGiYWfu4itsMxZi4CRTpwOzo7TrFj
vRnANTv1uQCG84xZYl39VReArvxBBsRVF/8Uvd6bEaUO0aYP6fl7IWjAg2nXx00P
s7VueUSG+rIMSyo0sgROHihXSq7S9AN188+HSO/IxDe8mfLvcjiV9KHvdKfIvgqL
2Wpfw4c2RbtS9WX1me7fsVWWJLc1djqJ/x40nm2nCKEIYCa6Xw3SKTJoIHFSlFhM
0GwMQcEbfeCUJIq/DDrjnP3AUwk4gCc9iOQl4IHk4b5G+LsxKx20HLpEnRxCwC8l
IavZHcm4tlFDd7nB24Jdj6n0GN6PGz6kxAdFRKxKdZkIQYa1n9XdnEf9EO6Zq5Ic
URX1jnUTEsUQpOpy9YEYcs1aNkMJ/i77VRcX5BGuGiMFw3ge+zwC+hfZL3sG6/TD
L4iW1QFhE4GKFLK54l+plFbdYwqPC/QLieJTFiS9iK5LKr4+JAeXsAFPNNJ6bfpj
S1HdnE7xKoRVr7LmSQOiOsWCM7n69m+irsmhTVONH+iRCHLLBlrcg8tkvO/pRZkZ
UlUW2EpeiFQkXBpYpxKM7G4lO5nTaiGXl69Avwedpmo=
`protect END_PROTECTED
