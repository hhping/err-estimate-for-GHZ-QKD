`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tyLXfZWgk6Pb+RqIdL7Y9tK6rhTCdqVKYpDzGYA/PQ4YFyPB1QM7M+uyTMrA5nDe
q0d3j7B2RARQ4mTKjc47oQzPll3BZj2lpHt1QJMEVC8nJfU/fhKfIO3lPqA6dxx1
MpF9Gbck6j9c74zFc6PVeGrqT1zgUuwxA7Py+yr8O56zHlx7f3u3Rwu9co7fWJ6H
LczIGuhXyBQg5Azdb/TmwMl0lNoYHINXOvrtvB/Y8H3HdRYN9Isb0wrY7usOQS4P
q28zC4fr/bdKi/EWz5m4oDY5PbZuodeoIfYC0OLDOky8xZE/YtwOCW5YteYJEtRq
IW0KxtzzJaR5j0uPKgr9fMH4wjyo3jZVUrGpJ2OlV0yNoAelUDmM3hurZ22CICG5
2yrj1CpMTpG2V+mqPJxEfZXw5l6IMhgzBcoCH7bO9V0bZF2Hum//rKI189qKk0I7
sK3yJLFCIuJhMA9XYkdAKvxQrxB0SZbciWWWiRBGVM53/aLfl/QlUVcVR/QTxidS
93aHl2BphKWS8BXE/BXfjhW9F1M7czRtwZbgX/D1lgA5QwT0pR3f37kw+q8JvOlq
QwGk1IlyfeKf2sMq4/ao7j0ywNHr75LiJCb1PQv98GvQpaRGEs1CO1p4rciluTmx
VaHKLxdl62NIlg+VbiKorkwrO0HInop7jUP13oSdnXeT95+/0gbaMBM9zYOzDh/c
CRWHUuRY4h1kwUGLQzQWbxZgahRVAZcS+tmMlNTV3QfRioOK22oOzCNa4zm8go9l
vFHF2yXqwdPzs7PbWxM5VGJuSIuJxh7yYZtdTa1jpAyp5j7KkAEOuPqtsmAU3wAD
thZgY/i23mWVmvHO1Z0/dIJySB/ypBV3D20TyIac19jw9ke4nFInQY0yCs0Bk5ix
z2CUC4SWrsvq7BP5E8rxLQU5zDIFfc6JkHB2pDYAc9oc6pmfSSE6+44irdMzReEX
mFn1/MDb4vMC38/XNwPTXNvXXhbjO5WAYAnUwax//C7SXtxvXMYCtQba6MQEH5Q3
JgZgzFRh/wQv4dw6H5nca4PmLlCdiEHElQhEAtxwqC1hzMmpKiZzW+Acy0IEMyLM
VO/bJ9PUpdifXFCGsymHuDi9z2XApVGT6V8DAOeSYN88BJGd9/IybAPbtzrmocDx
vc3RpsWT1COHbEjvHb7DXVaFJcqg3udcMgdAKGJe1jA7wA2msTPtIOYuBPgd9AIO
9jiZvhvzzR+MIfuGm4QvTJexn6lIAH9Wm8m/D6XhU+hH3horGHhk8XcoCxhzXQHu
Uyd0xgT1WXpiGY9/8SHk65nWZu38E2kGMY9BDpGGg5r29oTkmTotq/AyfivB4w5V
Zw7E/0oTvV+zQkwG6O4gntJ1k/vu8D3/r176dWcW4HHItbbSnxakOU7huvs/W5Ui
aqPNlY4eMuj5pXqLVp10EQY2riDSzaf6iY+p7G9EBDxxjUgbWphbtRdL/+g5RC6X
CpYQnPUGft5G+eUl2aTaszavrSioquR3EZc0wFKSqOfaykWur+OYTSqHZBxMuCSN
QRNJhYMS+k4qQFX9MBkp3rE8f4e73zcs/a37shjMTP4PAtHfXtp46e01LADvN+Q8
`protect END_PROTECTED
