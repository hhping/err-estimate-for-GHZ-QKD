`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIGCiIlpAqD4asWrZotsjVbF2+ejg1q7Dm6jJIZIuOYJ+XLDRpAGlEh1fy3wmRS5
GdnNM/SFJMtGW0gcJH4h/FTqwnGnuGfhVUWDRaNebodFlCc2C8RrWinBocJPnDYf
UCd31PRtYufAhA3tuGXYekImNgeoxmXz2SXeWtJSrT3VeZ5gjq3hC4hhzUuk+uE+
7CcrnNPHp3tP8LQjwMLlP1wk/GrUmOaITfwNOVbr2U3ZBdQcI6K7PhTTdKeuBunZ
/SITCAMJspFAWfik9CzYf7IRjhdcXzd0G6J/pV84r+Fk+/47RgTnHSkYnn5VDlOO
YPHW3e5XbQPo4uNU940aYWV4ShkCVxlQISAWufsSSycywAOzD4RgTpQCLkshuUq0
7niMFRRk0xxIckWggl5Ly2CNM3g/cJBCHLUguP7uRQDKg3aBXA4Jzfpy8SPskQDw
/9/1/9a1SjJWwrDqlrZNltFJy0+tQoSGVUw7CMCOmm6+hJA8ALgsPXJlsFMF5Ylf
xLRV0qmx4Xxvxcc2TTCFaewhY5z7MK73D5j8aIsxRtFgPLYz077NktJE80DfH4pB
SThffYPmcFAav7vJed/9Ev365k0FVZc3C6mD/GvGeY7eF2n2RGak0gAS9RmJgjqH
ptX5MlPZM4sBsGAdEJt32buEpIGmWqQQB78dyGwsIse/sAXoNn2pGtTVdJPQz7IU
M10FO6YKb9JWsq5LwXfspKKQNnNrZzvbs52fMN1TmAswTU9lWVERCIv58B+HepF5
h6cBur7Xn60j5feV7sjqkUt5mYDHkeRdrrqJxeqbt6BWZOCatB4DN3pdtCuE8b6/
KQ6Oj35+S6PZU7WW5Pvd8PCXtyFg5LjrgjslLfdWB6aDTnKsUgZKOfHhKM0b37Ta
4gETguGETG576GXpmQ03Qg==
`protect END_PROTECTED
