`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CwgUj1eBX+mA5d3b/P9udM5zQn4NCCQw7dYnVOu6VnNRYV2VW5jYLnsh7I2S0wDg
2LNzJ1f6NVi6ZdTCuvy8Wp1AUMVWLdcK3bcfflKXQfJaea7ABeEtih9sFSSAyxsF
MdrjDCALfX3jygx6Zhh84Wme+BfrvhznWfqJ3We/83lN41SYwVnp5Rxpw+n5N7H0
gAsRKPMHvuhZkRIpDCdTWHtoS3c2f9hQgP4+Q8ndYhcF12ks8O64bTEM2EspKJnd
x96TdepBWnw4oA5vlRwPlT3MBCGsHi1wldM9UnQs2QdSjik30Ly4xPy/DQxLavCg
M8voFpt9CXlJPr6VOq1eIg==
`protect END_PROTECTED
