`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aA3yEvWXxFMe4D0cV4UlDAhUfUlZTh5SM1C8VrOcNHucUBGg0FpVc4R8azb3HCxa
7+VlWc13UjBN/F+N8gH+D5MwrgWYWiEXFlPOMOvAGjESsAWJIMICN3a4FuAhEgEH
DAyflNQfl2vORsI9WXdHYyphmGxpnkZTgC9w+rZPaDCdAxMZmfgFP5nUeKuqk+93
DpjM9V9n4mQxsrlWSv9f44SQWGQp/X66OGr37FzYNG6RGFSOXaiFzGNzbb0TS40e
r3en4/OCWH+XKBGtgkCF+yRw27jinBxK5tRxdCUEwcCVb+VxGEhq9GxiHIrZjetE
jyiBzD3nfmfB2OvSlLdU+t7ddo1tBe+4VhRHUVqZi2GhU4pzp238IK2UtL7tUqCJ
wLKMvPRnfhQcgVmBXW1xBqep/r+kdO2OukQWBz83u4GMbmzPwhcJLoFTpNkKDba7
hpaYuY2B7wKZBSMkY+FcRn6NdA73BB9BaVIVy6mtEaFjK169aE37Ss+aGvBSEWeX
KgZQ+7mhsmX/Vp7u13WTxVf5WzIIgIcAkY+EYlMH1UYMt0rPEPJefvFLFBcXKYOh
2fY9PJ9Men6eqo6jqrr6rJzim5/xif9FEdiHUZKFTKZ+3T5U6WR2uMNfXznwhoUW
S0gAUMpAoZVU3iW/Dp8APCXamZT18wkK81zqMB1TW0FbIGOlEzTKBcaq1z03bdVn
nvyYWA1Hq+gSMZ58L9FVaX+zn+4c8rehg42901FBODFh63dpn2ikR+rxRNPiw+5f
IH+DN8mrG8cKRb4zSHehxNoZ9e2b9Be7XLQpnBIbk+2tSmGZ4XT2v+azenmy/txR
mbYb++CdrIUoQ/mjekAZiyoNuW/Al+PqPQQ/VTk5mjHZWJ1QF5ES7dwVr+f/fHYX
HVorLl0Ik8JFyGCYsFC7Clwzv6NXlbRPE7G9SxfjRRW69mIcuKIE0tdLX5z6eg7p
z3nbafC7jkE4Kk1KYOJUvmN/bi+tEPyqucKRIJ9sjSuMFcPRQ9keRhMEuGQ5CkPB
gSeVjVzkLSxD8NeRoXtrhERuO+RqqJebjY+MVUdzMl6ZVuXduqDFVVXZXfHaUvyv
Kcmp3CkimCVHPsrfUOcMuz9gVzgad1Gc5iOJBZrMNhp98wU2jgc8VbZra30/D31I
A1EDbnX5YkA+7GcfuzOYPLWeQ83exl6Ua0osfVMr4OhaCFQ8RyxNTV0Q1YSMhT6B
cpUFUvlkNc2WDW7XHnB7n1occWqzKgat5MP4lEALfWll9726NXM173BH9HD3PXVO
`protect END_PROTECTED
