`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iw8vfcz+hnJSSBHI/u0jJ7Ejiopzulv9gFHpElHOvgpbHkuJLrmPdTQnpx56Y46u
rBXEsyC7D1t2gIrDx8oz+qZxcSechLaipr15RVVdccifu0c67fCtspck89LC9Frt
2gDouvKMUc6KlwMLGg0wO1ZGiTiijuhdU+IRBO8JKljkvC5Y4LWVLzqcaN6ovSGE
8wvsE10qW5p80pZQUudaW8Q4P2sb58X/e0IR6+oS696SdHHIwI9K3pDyxbQteUxY
gt9MQyKMDE7PqqFftE9iCV7SwOpTjfKxw67SjUwYZwo7ifZNEA5p2jmMicpsJHHE
1QcS7/c5RplC51KjKKMLe/cGBhLnK/d3gsoFURKemofnR02/+fcrGeD4HXmBYwph
sbFwyFFkLxv+w4x8Gu9rzossSuJhoSy9sExfjDq5vJH7UkUUT/Msbs0t45LRfJWv
y++RABVm+EQqbDeX2QnO+m5+40r3XmH2ool27Q5E4PBjzsndljQVtb7tR6xHSSKY
qLafLC1drvAFPP5sOOwlvc49p49mnTpV7sAQGmwJMU7KHVaDGF1d8gXLhOSXYNH5
5yZPJxk/1YCbHHj/IRtES/LtcgoMbaH3qc6V9Cv05fRZ6AU8Na20dhhHY+BkGksD
yOKMfChuaaOo9KtCB7RUmqSAe6xzij5HJBw/Iw/689Xiz9suLFg72qYSnfUNPwky
kzz22+XpvbXl3jCb/F7CL64VehADz7JNzGzL6uQ9vdhRsEoG4a9GNcCFaC9tW/e6
y6J3SAEyjDZOwoRM5y9DTWjNglYXgTh9PFSpeAQtUbz+9ytse92luP5ihvytF4eM
Dqys+HONeEC8sbg5R9StieEKPgKPMNv97JNXDQipyYVOmHtQZbCbR34jFAeivrx0
DljV17TwgEfjtq2IPi4DLENBU/lUzkn5K4OfFw518Jk/zWaFOZyReEhOYNW85sdb
a04mwBaN6iMMqJCSfcTJEHnzNHGiPY+1v04Q/IzlXKUyZ6ID1ko0x/5BelG0nOxl
vZWe0Z7HsjiskItMkisfDg0MxGhwtCkoNuAHJEgFhlsT3r2e4mcwXe69/bDj9jos
VOznxPTNvqdnb4zYoRO4O9pzcf9O94LGFdrKyfF15arWImULbmnxPP2mKLbbYAdR
qyMIc4y1hYscXPrmg7meaBAh1VrWwykTLKD8ck4fcSfcV0cfQr8tK0QHv+UFK/rE
o0V2nLd6Bc+dHU2vs5jKrPhFrgx7OutO1niTuNZz9g/OcBHlEPCudnvtih6U8B0i
Y/bXFN/0iutP9jAF4Edp7+Edg+qPM3iIWb1z7zJmaBZnVSgXPryXbaSWR8UKTd9V
cYLw52zhT9IBo7DYszTEtJ1qMzZtoYx50ns80zqnqDRrlBL0ykpCM2WKKGJTcG2e
Q8tiNmC7wiUugFLKlSHLiwAfasgbJ1OKHHwvmk4DsmAMmpdzLtAmKMy31lg/0DwX
AF26Qrlq1OneTZ4cWdngl6OI9TvcZjhMo63iNIj8BR6aV2UZ2nhdc7nqH9YAa/nT
5oW+gG4Yb24wtY3zXmycTBu+K2vAz8LkytFxITbuOIo7yKfXDGGZF6UiazT4j4y3
DjCSYXmMmEL72htpNzJx7DEHrNWAo5LS8lL6CA4kQvpSxn1YvRlYnpRnFxw3FOOX
3gNB1pDHOZv0quUTWcYKiGoolM0Ysm+89pgpdiqe9LJs3/EHTKR6D5khFtdUdZFa
uKuvdzixp+KStz6T3aUnEfHkH42dq20Zseg/jQ14sMqS6qO65hh+Q2eiEJTn0s+g
L10LP9PVXpetkLS45LE/dZP5kFEx3HuEWqkZ2pC+cwkwxeTPuOQiO2RIGNId/8x+
o5MlTT4iE9eeaZlIz0Gs2J8/oyWhwwynSLH0k74X7byHGTOPC9xbfYafvIiQvKKq
sRv+uQChqf+VgVaoRUQxWZRWuRdh9B9+vd7sDTvBlx9cYZiI41WZ2jl4xaJQ89J0
ypqp3eVs2T/9igwwv8wK9JgAwwciSK4BjcH3pRjZmzBVt187ZtdOtss6jO7mX7fM
LkA+mr9l4RYmdZrsPbwLIw2YuKolg4qINRprWPMZ3+9nk2GyJF9JxRJXIasoMpuD
k0DFuu0b7z2DqNol54kRi93to5hJInqORUurI7P895N/zm9Q5wdjg04QTGgOm0Sw
rf5dy0BI1CkkiFZgPZX52Rdm3jRzU/dtSfL2HUYUIgpNNFY69s2LXNZPEhpAGwSa
g0aHTR8sWAFNpEcQ24DuXfcj2eOFYeXn3Fhf8lLjpBXPYlj0sVBVzh4ZG62O9mQ/
uM0gA5tI05aY7gj/gl8Fzdc7DwDYE9/ncOq8vXrxEI1BmLwT89/i0EazJPpaZdx+
a3bJfxtF2802S5HboLOM7w==
`protect END_PROTECTED
