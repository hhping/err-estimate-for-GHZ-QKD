`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4N6ktjfLIoW93Nnl/7XmElhwWIwNUXV44UJlHW4lmHtO8C2vHp3bFHY3JXQfboYG
uUhzYkHFu29P4OOopBnXfacbF+A8Sh/NtVhoHr/XWstTWApIBeybCShEEc1h+1+H
WRozq36qt30e7qnBaYeFXfJ5+mK2v/SW5KDkuMA+j1Dmw/Tiw/fCm7ZmUDID4QSM
uxMABbOGXcltCDYET5w+zZepHgwGRwydj15VE+YDDXO9ptJIVrTHe6ypBAN9GBuc
NBeA/eFTX/YX9b9Aa6x8OY+J1eKkRoyMYik4IZzwsKK4RiBxf9Kk8wYTPOYr8+ql
BFore4rJEh+sQZEPfp2mkRLADjfd2OUtfv0uJr9fuSeS9WLIPq5s+HaYmiBb/S60
Q9HmHSC/zxma2TyMRuwHK6trHQmCtJCt+WURUIL9JioO9s9WqXWlgH8KxamL1d7q
pkiZSWEh1vkih0W66TvKJ5ESMkDeLXnV1h3KsKmCU41m46BVVq/MzNddFXLKxZAa
bJ/mBxcYfheNysy/qRy/Oiilq/4NYuOFIm4TCAXG0i6EYdFW9oMP8IySUxGhV1V9
d9gIAJqhYjHobMuf0+gxKTFDSqAH4CCc7aGxWtU5mB1/espb82gKIxqhkp/Pqbg5
zDkOQWGqpV6YlL4OHUxePyRtDPQsNlfU/7qJbcCVi7z99DzSYSENxhxi2IvNfHtg
d2FL+9OuTYr1Dvh170z9XkygxUSj27Mq2Tb6nz4JnR9d3Ks6sq8tQo00aVtUdKok
EnK8UhJeqyOHUPGrSWz25kCJj1JsGE5RZpusF3Kw39lJkvVrqGy9xMqTHJL3FpYX
drI5SVOL6b8Km8u01DFPT+2TF7TEgGKrrRLy30QBOwIF+VCGvZrS+fY+fk9SOXHb
xpmyOLe/fBGRgAJEfNp0fqVXSKIR061wfBVr+8fvIWzBW4+biCS7acGu5HZgMrLQ
fGyI85//3JBhMWBP9cvNgWGHXDYbM1mniluVB9dyJKlIq81YzrNuDu5IxOfTpsmN
xvwEjQUbXjJm7/cZBG9PU81BV8nnXzOu0TdHyUCkO4qnS2uIQyEF/YlTgGQ9X3HA
phJ13GcOdoTeFYs5pNLYrAg1LNiQQN66KCX1dYZ/L6z4/h4cATGsoEFSs21/zSJF
SscCrSoJaCcnS4vvNEwQRb/nWDvsaxReRjygkGRLUA2GnxbN4JHisCQAg83yf6uy
xnlqZ7ytLOxc8LSe0XHbTiKs1hPtk8jHKePsQCgOUSC7mM36+q7bpWOySZXQ6tmL
k35Si3IifG5TAWgLaa6h+wzbaLGh+aK+VayFsz6hkq/NRS50pBnb/RsUD+/jzZXG
dL7BLFgqMtK7g2w0NSSH8ixVjQhnCzhAT3e/d+bACoY/KsvMkLlD5zgG5nvdfkse
1xOXf5KL7Y9Z0Tt7F0w0XwonSRWihKAO6NOp8yEiNkFEiZzGpUY+sfLd8EBlkJgk
8o+nidUalWahZf2n2Wz/AIFtSnPzVS5/C8P+NgWxg7W8ho0u5E9RGUSUgUQFNdlZ
bQBqxXeM0saDdn/fsqVGnJ49oYOE2nCakiqIJPfRRhM=
`protect END_PROTECTED
