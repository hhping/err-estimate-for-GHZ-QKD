`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ePP8uDfju1MReu52almOXK7q27HuPujz4ZBaq2uFvAr+YP1reqz3ijylLU/57h1
KrZd15zr0p0O6oQqfLWtZKUB4Q07ocXgB8o/qqGNKpkTg5abbPFyD03eWJTd+ulb
b9lLbHH9qM3OCi5Y5KwCTlFAZIXm0KQQ+KsqQCOEj9LFE/Z0LPHvW53k16bF11xM
OwIyJQ953UQ4IExWCN/MG606Qa04bBzW9TkI4B5tn6ZfkcbHQdwHs0Ro73s099y9
x9gumJYa6tGAgAWs0dmGh8tnwzfCHLFCl9EgeDuf5qHIHNMySM6mJVc0MdYYt8pC
6MyucTRG+rS7AM/9amQFdFmAkbGdDcT7+nuuFrbUDKl7KRYiMy9HkTQgBpbLyImE
mbBexoXu6kt4v56SkhWtFRt/opouj8Vo8jjbobf3JljpifVl4jdufuRUAvNXw1hk
cDDcqRwI0QtMxpJlazhlpnw6L+kXs0fR+pHdviRdFnqKM1JKBZ0mPqlzakaR51h7
z77uxBdEm5XKqIRJ0ZYy54tRpGGSTD/cfCbG+3/DT3TrjRibxZMNr/2JlV5JQgXl
4D+RdbgPEbwXv+ngXL4soUWCKP6HzuQazvu+xW0T3/EHbQSRBZBwO8j5/R5MfL4G
CPnBlTI5D9FQpvsu0f2CfzNkWwZzJjgJL0/hcJ9kWTQdKCFPQH2Pak1GQ8uK/9tT
IiDzgOKub2eAim7y4xxil1Jc8AU7Ks5239P+PrXVGNI1y80EkhcvAXf0EERYTmkn
gdcWuVNL6tqAZ22Qh/UEIowWP86nlj0G75uSIZVzBuDVQLVvBOaHdPy5gA83dgVE
0SCD5AQ+KtE9sb2F1eB/BoxWki+78M4b7rp30Ck+mVYMyiWr16mz55YufApyLvPd
unqwn2977XvEVSDRRWeNmObewIfqKvOXF0ojRM7dHV/tICK1Fzn3INinfhIxcRGk
6F+m1In2wbG0iLw0eISPsQ==
`protect END_PROTECTED
