`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/RK0WzMiScqUdj6aaYZypG6OGCYSBYWz/lK0H+TXVzGOhKefDLZ+gp5/eHTQ3Ia
SeM+TK5ndzBQYVCV91CrTgAq+qTiPRS+fptsLQXdtJPD7TL4UE9RLXUeWXgvZ8Ng
RRdztaGHtgzNfGOVLCMp0TqwcKb2+jm2+bCv1NNGKMrSh/tfxFiJOP4jBvRIZFNp
TLnQl8y/aoX0wypfuZjSdWFQPn2xouo+3mdBJ5aXva31NLAGkfTSlcLoy80GHXF6
5+JDHhIcI9VL/SVxeSY4+ueqJs5D2ku2iwajtl0fc2ydqbsvzd2pkdR/ky6j/r/6
3BMW8/Gp0TJKg5xSHqn2EMJRpH9/3wFTHsuzRlX1JuVwXPDjXLpqMtWdSTmeBuLI
xTnZE5LHONl1pt/iKObcTpKyLahlVrUGn94KRns23LDD6IMDoh4+tHNCxad5iWIk
wZuMAEU+eO/3dgk10HBHD0fRGyJccnSvNvchpk2/9+vG0KjNG+/x0VWCB8uYJDf0
155rdeAvN/eLL+ls4KeShBp+Sq9+bWh9SAYiRHPg5d2O3UQCNhNYNqUwGIK+IpKJ
cvD/XYMvNTPGEg751nS3PtV9klgecl4TYi8bRvUR6TPbqXT+tsRZF8ZbXdMVlM7k
4DeVStJ9DZlFhLAsr4tQhcUh0PMHmqaRsTfSfpA8pOyr/dYsiXdEO0zn27fDQ5LM
uAdbiS6Asz+k766PyYQ3CIwTm3ZapYOt6dluUTCzqaS/Yga7lRqrsxKpF2F68kyK
02RAteXh56itudIwaFhdYaJ/bjb+eKrbHkFRF91jgEQpYEbB3wF7UwvirjTSXuSp
fguHmav0CdyumTLoaSgCYWfg+HYG40BlZxNusVR+i58EyUpAfDZhTdiXtGFKVk0s
QnMdjtANMWhkegFTRW1empezEKvKBQMxO0Z/n77NAd8fb07iFGt7OGnUWCCZ8PL8
4zx0BUFdObLdJJiMRSJ8p1iGFwL5ljz19zsOeOhNpV8JOk/7VIgRDhRW42JO6tnd
X8OPUi8z8E45iyLOR/tOiSM/2x/5xLZdJZF2OLkswjbpMm8ty0p1lFrKf/GyFx+E
IOIsqkJRFRcEIWuEMByQNRWUg79/QXO170ga9s0xHUvB37dT6o9S4zC4ZOLlVbXG
zi+t3LjMBwXZLrkoG3Pmt48mZN/BwPPCCCVAGFv2XsihZv/dtyNoXmNp+RNLKilb
YXlAV2fvnSwRS+0cnBXbHz3b/wpu0EkUKDL8hOI5wAOkxqTbKorzkzZo2mjLYDl+
A6SBG0b+kfa++S9WgLB60vp/EX9JII3D9QECDdkH7PWvj4QcWE3HY7nCEwirtnP3
jfKcJA3aCvPPT6a9p/6UrscCXf5l00GEDM8UQ8eFLZ+Yo2IMERz8hZDEZrY1et8N
eoy9HhNFAj6/9ELoNbKO1vJv/x3HRpwW4lkq1XhJ5+IevtBslQiuJyz8kf1WJpNh
b51G2EBtBarxG+aHIOQNJPbVgLj2d9PQRfnKLoh5gBuQUr7HOjLzRbukHMnwNBkF
sDf4eX2l9YwiU6NDzClVipjlqOvAZHaiirOW0emiytzBLgAFRLSy4KuhGIW93Lef
VSBCGMQZPIaTTU94NtvoZAKvcPQJvjdr5+/sS3Mt+KQ3yP2KEVWI3QzELO43wV8d
OuyCrv9ii7pgKvBm/4/cQ6YRno1+5homOvMrHwdVJfuOlaN957PvTFX/KgiN459O
0S84SzrbEX/qLcIgp3n6e+t9O5wBVIugcH6ddHIDN/m6CDDRIYxevwbvC0mQl9rW
kX56P22Z9RnPzh08fADgY1p4f50xEKbpj6HIBgI6AIJav/E26UDeMyVFo5wKJdEp
bp0kmFKlG9BbwgZgufQKKLXQTrzIbWSVtZTSg09RW/jpORgpKZiRLeSyllR4Lvfb
p9JjmZszrQGZAEoTEOLw5qVvuMmN6ZvsNlFzIjmL5KFolI3Cptde0JD9AmoPezlC
qaz0EqqGZCmANxW+Bf688hURx+ybcjRRpK94eqHdous7wFE2PVaorrK240lNbilV
+Wsu1wsi/RDU6Ae23fjaQYHMF1CD1RB+rBKH+gTX04zCGIa0OoR2MG3yrLcMe6YA
R3l5Pui15ijEaQK8N62AzKHdhssSVhpTQUFhdbTsuUl1rX0hSNUUgHQcxmGsfYOs
Y2l17lwaI5MeTr5NTi80T/7cp4T1MuvSCxqayjzahT5Or47luNT8fTmVLfEiNMq3
7/V9wizl2Q6V0Vv2PIsX5K4lrQagXzsxIVXWO7zysTisH7svkJh8dNwJG7W23hIU
yjGgcyGKaJAv9Uq7EMFV8hVKdowEfzxMgx8eZ6g5Ks7p5NncXl+GNJdGR5nzWti/
ymk5IWDt13wyG9buUsaHxFxZNQIvvR11JXyvCr20WSnAm/CN24kZhGL5I+dApFDB
MFQefAdho6O+Sx+g9S0Y4JzsIZSWuvGNwiBaQDHFhwMuYflCsYaxWnOgbd8P81VL
gZ8Jz4ucvG6PjuI1zYsM1BIqTHGk6X62sMW63WRXxd0Gpj56RoZ/HrKsJRprcIr4
rlcDtKe2mPIKaJqhjokpb/i6Woss2u+iR4DMdTx6EI0iCh+0EUe2ziOedY3Q4vnH
QthO6bNDreGMQHCZCh9xKy+c4IQdJpypHhNj3dwfLEDOh2pZe6saJxvkZvAnqP2d
6ubmbLypGFAa5JkP9aC9MAQsp/6utlj1aU7BdE/77Ev2eysiqKA944lskJAb/2j6
7cm64jqZMO5h97Y/C8THgdlbZ2XSVXH6ewFgwx/kcjpd24bMBrocFOEi35xzN48F
o/x7LJiLk7mOUc6lEdzbJrry/fKbFcQj9WI8nIUeYcn80ezKVhMBHoCJOx9L8zZ9
90Zi5vZpbuXVic7tdSTfnRkFE3B7tKUaIPgkI0W3cEGuvgs55FC7p2Ym0DnO0ni5
jSSbP1CT+tgO5vkCvB8wUKFTWD1vWmSBb4WmMJjmRZzP6aH2TikwEMgMMljyqAdc
QpeUBRWjvbOTmbt10+hvSukD0bFdjMzP304P82k1ygGEWX5YBi5ktSvFF/tdN55S
wF84nAbF2Tyy1fn9OoMndH3K4h/YdadQiq1YRjWx7G06ovJElP6XKWgT6NhVRcrh
1Jh4Fw6juM3KyOPvsBMwvxMqPUDCBU0bZxisIsfIPLRRvfzOtQMvBFWNnWiVEnKT
/cIxS61N0u1b39qv3vfJ+ieiY/oBy0CDTEE4OlTu7aqXd5ihgFUxIdkH91Tl5rOJ
pO1AwTX/PXhCugQRKjeJYJRIPMMK+IXC7Gk+Tj9G2HE+Z1XAG4IwRaQ/zEKAdd/t
0QH5HnXOpbd2dCNY3c2mUpM1R6IMf5L/vQ7EuUf3vY6uDUTG2+1FYzORiOREggLN
Y+e2lcJfB6jY4Eb1DvzLB4hsrcoPdDiz/AwIyZd+N3C98ZUyNWOvl37NyiVaqjKg
WVumwYvEdV2ORO1qpksmwYwJxXj5CSLSQ+Owdgw+eLNhncI0hceIpOiKVQywMKRv
BVRmdjf1ebpLEGVXrar74webJ6NiUIyRMQ9lT0s7XdwsvlN7Ro5khPY+/0aZ/fNc
L+/CJ7frKVp+Jseb/y8U6wbfuyWiTDCeFcgzBXNZwC4oHXUxxmEoTQ4jNHkINMsC
nsPwhAmrRdX63QbZf64F6Yb5N04D2IsyCRo8n88D7HxDJsOVAQd/TgP63M0/SeFZ
mYz/iQUn4OOskR6Nh8O1s6y9DGMWcWyB0t9rsRMj+U4FWoEd+VUazzZqPevaWTTE
ChERkKmgx+nck0sg93lVcKCauM4z1lWTGrtNXURRVyW1wHEuumbw0ZttrGAkGhIc
KwS/P50O3/t2IxZE++3wdVB9FGE1/ujjEExC0pOwFvQJrYSdh9o/AeZAj9+IgVvM
9gEwkyN46tHIBuUnNi4kpNGBzwZ5o6Hqnu3A4E2AuWfJ8NrZKEgg9eE/+KFs9oRM
IVg2w5TerlRl3VuQ1z/22bCi28Wt2qv1N4nBaSLsKieC8qN3Q+5ZQynFK1YmEat2
OlU9Er7KivdgLzWaIWIbc8eUyJkvMYyXpbVINZF0rNOCHg89/anRh0eQeU1KbaIE
thBxweJqa6iM5RYlsmkzvURfhiVfTYUQdXl/4QjB+7L1hUSgVAFxbSu8A34dWlj1
XyyJQ4tHlLXTZt755FPJqLsk5SmQtXn384Bu2x9n5eRMIVXFpPHvVwzPrV+O+mc9
7vng7/r5DRRX050YgErLfEQkrchTKqvqOZPEdMqmIIhmCnxlCL9Vwtnn9XYUYe6q
8XWCCGgKZetD0bxWfukQT5nQyucsMQEUtWm86pO8romXLpEGiKw3Lxt0kOiE+LZu
b1UqgILOu0tEY3d77QnM6IGZSP6HqHF8ZmM5LxSa5Q8T2xZ/360R8uJsllazwpx4
PTklbzV2QXFibzZ0xhoBqdM/3etiLwFup4ZR5xAs+A+9MCGwaM9SfMPrDxD8nfIo
90eSgj1QiSZPQI2X+eOXlGrL/ycJXC+/0J32XKGl9feSGMd8bNUDVpWwFBzOB6qL
3+qRexqp5d8OzbeqYR02l+VqPGj+oLhpLdSp82jGcU2pATF3DqLlL7LyLqlP5vph
CiPEgaWxNmAZMzIrSFXIbq+wbMHpby7Udjx4zTQ9o2diev5XhhWrmZri1oPGaHB9
oo1ng4JC7QYEMMlVpwzrqK8nWzl0/P8446h9SjjKuL39iWph3E+u2bR3H/9mZawt
os3ERKuaPjHMnBoX8Yn18Qw96tEnNqOQDi10bQiT30onN9C4ym6O6TfwXrlFmzt1
mHihs4B3Z1nWBDfVFnqg06Q3S5u4UnOYgiQgPlh9v5MMr5wIE/C1kswLmKWQb9wF
nz6WBBlAuhymw4IEB4+Lh3COOqAQePB2uLrg6+K/ohWLaQr0UO7wtRupLnDpXFyq
yhbQzxDoLNnD7ymF2H4O6d97bIUvqQ/6kStwAMAYK2Hyg4w91Njv1g0eHK2IgtjG
b5rDqK5ZHHj7C4TPAMKpyQAfDjIGpAm1hp6ZPyqiy61fCpVurDKHF/e0O1PlVCum
EFjwtuIcIVCP2WxPK4IhbE2YNkHIqM55HyEUxo2KyaSP1605NkoLp+wVw4HvRMkZ
5LjFsvqK8osfzlGbDf24xCFdhjUpwJZxzS1BiehIs8kapVLkfNmzzc5SUPBOzyRl
JKa4th4Q5LvP822PI4bm4ebBt02eHD2bOmUvGwQg8OhIfh2cco/CoD93JOY2u2NP
hB6TTVSWD4p2R8PJWjxOUsZoWrKDbzufQ+KqLyygqxpkAb1CLaRqiCTfDO5WKFCj
o7+cnpriczs4nlaL7Xqvl+/ERj34fqcdBMFF175cc9D50UvwUlO5WCtU612juX7p
iMYxw29567/ZV5zUhHFxe/h5p81ORmalfQcmmWGMn05WdHYvM++jjVtZ9w9Qe5o/
yW05Oo4XER+206h6xiEQ4HaxEpyUu4Xpd9fADVlKJgVila7L0FcqZowDdKGhzExp
M2Tx7uAkq2fnxCFN/Qja2GeKz0DuCal7sobSGlJQu1rcqbVU00wNn10QhWBEGi9j
88KFufeatjj/ApV5h3uVj5czRDvYC1NL0bZfuvLFA7qzXoW84Bmlhf10VQdmBRas
lcEmcgZhUpXxRcpFQI3DNZVC83FfBgKPPIXoWMs1UNnbE9eNR3WcR60HCEJGj5X5
4WbUQYq4AENznLSdNEGpnGmrdnpY1b1DR2nB0YrlWhM9KRSE7HMaVu0mtyKUjWGS
uxIS9OVkZX1LCFQpEYzX24cEc9AYGiehWXcVL15YWrRo95PR3LzzJ3TPKVu2p+9W
3ckHKlb/MBCJ/CwNTwWnyh6Njrgf3Qev6IJCCPXXkLEyKcOTDmqWpEyagApXAy23
HgMPqiK8Ugfyi7IPreHYu2/NH9SGs/Lv0XtvmFLs/0lPb9v++WlpVjtX8IBIGNTz
fhF+8zxVwBnTrX1WO+BxrN5XvT3UDHlkQ0kIaepIH6Hs/3RntqjqxflLWFaNBm4M
ZvdRbDjHZ25bjwLNIZ8FnH6J1boYVC2fBb8yHfDv3mTEASV2kKM56EosRwtAkjgu
1lJTFMkq9U8KhyMy3oWMxESEeEQTCkugls2Ja2aw4W10Bde86HAiXWv+6oENz9jq
/U3PymOWQzdhZGEXIgIiyqZ241pjVnoQ5WazWBqGYcnkRit4ToRXwQOS5NWb4/KI
9vFP8VeKaqptdk7RYGomcavdjgXEfVNL9/I13Omgz4tMU1Yd9i6CRSkl6HQebPEC
dWQo6Lb857hkJwAti/O9xq86wDYSXmPs9IxrATMqptQnzzuvquPVj2cPQvV05enO
ZfSPqYC1i4n8vhuITlrMgW8boN6ImhHv7JeldzIjhIVuyLBkTlRFnmAT41ZsEtYj
SfBQZlFv0e6hK/9LtGy5XIuMUsKIHJHrha4pym7skl9U2ILmuW7yS82GpQ6FeBBi
GzRzqwo7dGVZMKmVusJTxRp90bsh/aolEYi5MkbmhNsqQGuGMOXyIGUohNJaMOd8
MaRkb4Scnw2LtVbj4pd+AFFNnet9sT3LLEBMd2S/+nmikpV0JOX5GJPQyl9Uf4kG
JBh090msCQXT7GODMOKO7lM0XZJxq2ronkTyVn92OowNcg+TxxbWDD/nxjwdkhPR
ztmg7TwAFdc03UqQsj2VXsDBbjHaD9j9sANDQklnbEZYaQ7K7lGrcFIGAPManW3Y
Ta0F0xH3+f2u4tHBOmnFp10+V4qRa2X+u40mraGNiRUDW64iA+zszMFf3e9Ng9CL
HkrSpAZDV2q9GwCj5NdRQuFw7tk53DXM2SflmD0kI8DdWekCFmibLPbUIkvA/WIR
ztY7+DLccthNUvSMmyg7oNyxF44rkGClYfKBKTEonz8Mo8pNgLfTl5jp+ssqNnaX
BovT2Wc33rx8yn7W4wp39Hw0YGopBcaXagtO9T5Bha4h6XCHG/BsBBwgOZlEUX3K
CSj6/MTaMP/7rkYTv1iiStTctyJfRDkRHMSv8gfcZk/2Y7gcbaGgdKngvHXIcsgz
F1dnmT25HOjKz+qNrW3x5wyYUqFATG4ltkbxDoG5JCbr2YKVcAMCQUmollTCiR7t
PZyhwH/nau4HF3QLLNB/iW531yAegaVPi9XqubmPGS/EBNEO+NLw2er91WpNWkD6
QwZwdrbjDZpq6V1DVTTjA8DFdNrWP61BP/iQ+Z0hkJohbV3Hjh07Rg7QbEcSKAMr
thpQEbsC6V8wBjQFBpojmDE6XWp9dnojm+Kjp2VsLj9vrwmYPjMymRZYmQcDIGva
4F19LKqHMLorJ6/L6Xjg15TAnJL/QDw8YMui2P9Hl0nfZvofkQ6tBy4xO4iVRDmI
Ifov4HDzNoiZUDfdiiMESJDMZio78tkQufTLQa3lUnZIyR0oFeifElMTL4pLjqXI
a7eebEFZVjii0lyOMQ7PjO73+L6FAiZwjI6mrsqAcDlRKvTfMmotSRkhaWNfSMDM
M4yEWFvscn9cj2IZi+iTlW85+EVtGl/0YL95DSxh4269MgkZ0ZiFQ2YixwHrull3
2Z6InqBifT0/tLc5cGTHY3Wzq9INmoKxhqhu5pT6zSTZ/ZBSaLsoZh4BEk48slZS
1Rq2RX32mNB8XiypzC9G1RCwD2OVbUGvEuqEcK0ASGDE3U5oTIOOoeqkxpxF0e2J
sdBkXd0yVQko54Sf0wW5+EqOR04Y9XyjwVub8AqH5rBqIpWjWMV4NHPBvEsanKCS
PzHoZsg2kjtKmFfc+PKugU4R4f5geHEIbLevcedJqBJrlS5Z9oLn6LoD5b9xBqK3
TKgxWuh4C/RsrBAnXzkhZkM/52B1vvxK6y4I5ZPUO149cxMV5YPMJTR5i6VNKeIr
8WDcO8VQs3/eurl37jLPltH4cOBHLdcF7Li5StvWYqKn15DY6pOtQSdZvwDUMNNM
GVLx4B3v4jgQhbQJ6KlfjBZ7UKOZA0NgyG2CXWt0D9a+69GnaySzLlOZX0w3nAjG
476OEzlcH64hbqe7rpNHnvB4JkuDpkfP3EYgYbOhz9rRXumBIGTbe8+sb5PUce1E
II4b+aXD51DQtEesx9/4SSEE6VtzHJ8qWzuZw2W5zx+RjDcTyTs3IarSX3D3TRQ5
MqsZzP7XMFW9DbDWiMCnDahAhAqPC9WAJE3T6duNSWX9+vFkRg6bvrDdwOsN1HTY
RGgKRnPEmANK9bxBV7f14uIGzYwIRskQvfKWQd+GE5p/92V7aWr2UcNACywrF4zK
T+rjnghK2JM1oADz5u0goPfqnajHTS+qxvb9mhKz6E6M6hbmoZaUqwEV9u5FurFC
k7TiaIEwr6KhlODhLj+oHoFdTPJdVtuZUbfyscEn8KT9TPRHFfn8UFyyn5RfBiVt
Nb/VWcxv2fkU/pJyTfld+NZ2k4CcuW8VbVX/pAP5QQpuu3FMVHM6RgVx9vfU4tu8
CmFdQjOZVoy0TuA5qZNITJFhkdVoiLAcDauCNPtPH9lem43Z2kbH4SDSlirda8AV
SQ+oaQUTG7bWzUOCdsBGLYA6BM3PQxsSyqwahdzqn08pQc2J/IUQrcRJYnep6OGr
75Ke4gBvvqIrvcmUkksFuIeefamlGRzmKFDJMBBgZHrW9zghB2tRKuzNz+4H0+40
2n3Fy6Y87jCpW6cgAQ67e0X/8mrqaIu3o/3d2o3eNRb7af23OCyqcDE+lfvzmd91
7HhUoV1JV+MPNG3aC2xxUVzV4zf4UGA0bhscrgoTgtVtQCczGFvN20NQltie7oMs
0af7dXLHxJUemW17gBLaxrZHCjAXKnHQBCsmYUcKLJInQt8+w4VOyalcRZbTFiMr
WDSdCKaACp6dDpp1VKL2dtlSKU+jrYLtGa1x/z+gTcwkRi5PbdZzrrv5MVtaTxC6
GLTFluCkkjZ8hNgO/fkJj9nni+3DdxkOBQ6TT/DktW+4zhmws/gshU9XUDSJuni+
dJ2o12pSei0V8q7ym7tcPsfmljO0XW64yNYnjm6IFrF6wL8z6yDRYtAM3uELqGWP
LBNX7JsVfDUhBCp3LU4s8L+jbxJgU7QaaC4MivEY5+MAFigOVW+StXFVGZooua3C
00VI5sKk4LPAJraZzVqwGVagn/y08+MycwJ68af8t1mvAKJtE/jhq6dXDumFEyct
Glaw/F8/EsSkPcSWmcQXI6AirGleZPziIzxCZO5fEtiJfG7PLdpvIsg6MXq+Fs+a
xdAd1+JgJmTUryDeI/U1qim2pBa72FVuKs1ZiaVQroWhmFnm5IEFBDRSX4GO1jkU
NBL9V21sLqYrATYVv6Zu3IkPIAYeFt4UGpPa/Z361bS6uo3kGuyn3VyvfvmQN8Vf
U8CrGRaKj2S7mC2aVfDIB0JL5Tl67sEtmY+aHCvCzmEmRoFS6IgwT6a7Pm5mFrCb
YDTOa3ZfXacDIxG2KxjUtaWGfORVXJ6lkE61ov8i5Y3TMSmXk8D75thN0yjzEcEi
KkEioQidyhHhiuljf2LTy7yTpWx23MVKrqd74xcsVtHeG3YxjUgrWDwEaGRrEmkD
fgpnO7iCviFbP1OWr6TGdHpXMgcR3UDtKSeHfeLvECGIJK8+SMn9FZTr3GGtIyeJ
XY8ZbuNtOBZbZfJ6KE+BKtpibygT6qbGkXpBUbzaXqMvNtT2J6uGsoCLBtQMTyUB
p+5WRdts5PMTsnPrx+gy3XQzMMwa6e5WctqF75dq0nHvLCtCP7As0kfAtd4Dtc9o
Mc/TGFW9rFYRED4bsP5cuPV7OSO5O8kdh5NphZMdUS7w49NySXc/AyOtYdoiQRAl
12/bevoOJcKmO8UUa/4tRPLXcOSty4GP1Dsgr8keetRm/ZDCqL1+uikSncxrg5Cn
RnZNDymWQYBU8MWc8lL90YaFOz9deb3ikSLhz9Ve91mj1Cw88WlS56JrF2m06M1R
usegwc1IgBEMkJINzUQxL2diFV6A/v68E+CQAY5iWvhLsAOkxj2ibIzl3kkytmft
PlbOH4nwDACS/js1IT7GmsTlwa4JCVmTmzTUmYaMsQAwooZJE7WTB4TDYVGUMVDW
I9ZlfxFdPu9JX9Me8NBO52jSTPAowbPTqSKkzmaeBUWP3KUck4EuCZkQyF9ig8FE
jYzjmEESwdyaoHamdruQnkNMGVbn2UyU42vQWlnYf/fGhVq0KiZ9plmZc/gT9tu+
tkcgzqzXlAfqwJrqLh1Pz1n6uyD6mpIfDOeDrYhAZwpg+ZXiofNmFsamm4tjkHFs
Mu7RXV1mYp13XJbDZlQbUrzXGi7kH+MOjvTs4fWzn+Pb/GXYOXtXV6zKzv30QH2W
qsWZTDs2HyPPX+E3a0DZE9IDpalnmfFB7xOnw2SgjfgNmIdETAhz52qgIsw0eSXC
vgS9xRms4vRL/fKHaOXnWu7om9ar+S9qDw+iZuB8Op7OZRDuZp2B1nNY5Ut9fYmM
JEySemNeTL3OR0D8h2VDO+6s+TJve8uEAOVX1kopPCW599eurjR+5ENncKWx4nPi
AS6fsx8j7nkETTy1GQ8M7/5Mq4eFDWCWPyCciUh0pY2bpY88gzLgXWJ7RBAIcx24
156DRCScpbk+zuXHzisVv2n4TF1/xCmatJskSQzWQpPeQ8IUMiep1526PqdYas8b
L3uGOVdodL+/nxz2RuVCP9MqwBaEzWGXn1bornJxvSkAp1sOxZBYs5JjgHKTCfOi
8TaWfh+XQbVuz/Y2EheOmDN5FlmswW/PqpESEjgo9f2P1wX15VT4x5YonFc3Wr/T
DTFCSpMz7YjtMwUrnjUlStkQXc/X7RMA9xqx+6yavdZrbPWLD4dtbzXrnJcqEDOj
yUb6WTT1AQb5QZzAONf9aDCu4PmhUEHSMBEWQZpL7ncj2cg5G3Dw8F+1QuCUYbV6
3Nk/4E4AZBaFI90YWjVcEj8YicsSqaXxPvBA9KvDR6mMyUoj/q0NLkzLAXGSzfZo
KBqn8obgn2+LDGEirr/YQ/bC3rZ4wE24CglVJJDpcHKf2a+qUml7Gliwf9f3Uay4
4k5iEkUEkfmCt40FsDAx2p2WT5aT11UenSCDW8lbiFLuhKGjgqBchRu48c8qiE9/
+TaxdTFw30/PWUnw7wmzlRPbvV+0H1F4mQo8/sLt2zGaw5n4IB5mDX2Ete2di2EB
3VrMRtuUIefjQM/t+PCBnrYqOz3pWTqC2dT6eSVp9xze0QZOaugjATc3rysteLgC
7dfMT/rT5h9D+OY/xBkJ7RL/BVFJpiJqyj+6oGKY/hNAC20EvsTLh/VTB/KqZpsL
S1KE9+OOALRV1cvDdg8XX9DDKbBToxou7XppT6shX9b9d1CqoerTEqh7F+bwL4vf
09ijN7Fy2JYmIIzR/9qTQX5XRCXF5KflaNahs8VTa9oHMfHg/DNwo3aQg7w6V8I7
hudLukGtnOEslXVdttvMs7U+ARGkS0bZaVr8++aPV3TAU9kKOObW4OLQnh+v9I8M
k5+cvuVGZlnLtvg68RWT3NRCa++qMAHKD6JXtwAkaI2dsgMYmHZyuLPoYYGk5c4s
0AnPcgEC16DFuyPgvSuoBke+WoklKDBoKDEnSGqgHWlUuIAlGZW/f1h0Rnf35JvW
9KjzMk6bQ9O2rSqwa/BB26a3+Wtkf6roGXhSyy9SDDohdoJqItCdtGhJA6jfifc4
ei1YHbU3TgjM+ERCQu7bTmlc/D7lTymiyNACOmoG6RruIXtRVohbPlL9l1LoYBzL
7sLly/aCCNDtTV63ckilk+yx6FMDLdAxPyXyLbQTwhWQYxGJWl/ZM+NUC0GIQJ2X
Asd5GRZ6XDK3R2xpbhTntVvoK+qwj8tv2fsKavQOjqfQGgr7AYx+oxwY/AyD62+7
0UGaGW/yl8sgPQxq+ixYYAa7uD2TL8POTapyzr+JX5BjT8CRYFLOiFDnmeQgOGsm
fOv5dB9gKc0K3UALvaP7cVxaEt4lmxaZCEFsp71Wn2xaysdts7hRtTbtXlsJ3k8z
u2SHGjFk1UpGtlLz2jNXqxBxncmH9Q9hczYxIhjQchhaXq4uMwtHgZnMvPKFWij+
Wwhbv/G39SRZ2el9HzLk5sC5Hepr4JSy0Qc3rUfLRfVntdzZ+5UwRffoMD14PT48
DkoStTB5Q2XR3n3+C5Gaz04UQsMPLUwy6mwrhgDNnz1UVUBkDKwI2BtiyNGCzvRe
/6XZb584OnNYqfSxg0Juts2B4ehgWZdRmyJUD80qg2KTruFxgraze/uS49072md7
EDKHjZAsZ5JMrgOxtZ9000r+lJtjP2zih23Ggc7MvWR/boe+pIRdgTm9Rs4zZu0q
KzvzXhIga0DKpzZNcL9aWgEsc7eZHDbiHJ47X/Lzjc443E62nbVU6ha5ZD6nfj2b
4lt+WHFZUiq4BDjFO+td0PvCCb+miYGXs2NquFDZ2YbvZbDo02gRt7vdQjG8nrmM
3H4gcYjh9xBpcKgOA4Mo7Qpo6xS3SCZLyzTDUz3hPULS9kLpUytFBGcfL3HOFExN
rZ8RTjO5HebxxpQOFstbTo7XyQh4kee/CB0a5jDN+0TYqulm3UFOgG78YAgd5dVT
atsEyyHm1A2H0/3OoKG43JjwjiTS9dIiOlCGr5F/NatURILzunW8efgnKo5HAtag
yjttonrPkHfAT9icLkzvl0uQXrWwzacTP/IeYjHz1VEFz5zoxwV3y0RWCzSYai0I
/d6HgbYZ7y/bH613dmMLT5vh697nL/Mzc9x9q7oLNrxFUSxyRtPlIzCntMiWzMRk
zlvfrFPAYBoV1rxjLTEt5r4EXjddgwy4ON9wWcOSpuEGLsTsuu2BmINNR9OCgNYS
QnbNXqyFxMcMhhKc0B0UCw/y2X3qR9rPz6B9ZVvYgz4f1917o5QV3AJ5Xfd8/2uD
rQ1+x5Zf492s7aWmM4dGHrv1ONvVJD1VTxz5ae0v/jwtO8RjFcT7E2ekzfESfuCm
jfGJi8/ry1KWNMNzIp1aTSd3+nqjeU78nOcIuhI9mIN5d8MaJ6V03kVC+wArCPX0
v+rDrx2dBVmd+MJc7WuOXUxE/trvbEs8vTyk3+tdi1TssOjJSUxjLOYnEze32z0E
I8KCsKvOB6FSN0VxU6WKZQCEc/I/BCaOEg94NKGN2eYH0dJAQyiUZ7n1Rbp+eMQT
h3ztj89LuaYLIz5/lyP2PKvueoZmmNikmnmPl8P1pYa9qJma46bukV5JUH5nzTFy
2hYDQl5vbrOchp00G/v5hAEErHx6zPu5aVkO7kjE7v9KlnA1YsDAFbgy4RZVKBoB
vbOw2EhUhmkCNJ2uj6kG2IHNQ+HFdtWqtH0r0MsWpDXAygJ00lGY2Nj3OytD12i/
QL09h6Q/xI16EQZnHYyqILdhoKlUfACFEOga2+2w1jjhi4RUv+DvdGBgd7lRnK2f
VbMAY6Gc5vUyI0aoprihXPNwBr0cowOqPbiT/mful9CX47Cc7TCee4q+Rkfp45bi
77uuBYGRjJQ8uk0GcblmfUqlj8nrPZ4RhY6GHd2/TVj7chSb/ICBE9fjoEJBcM37
G9IAYNUOeGei/wckrl5a31Jgj4tu6qup4AWtSICv8ox3ggnhWcpT9Aqs2n09ojak
qG15Pe+uvyeN/Zxm4z8jkM6RP7KsIoVlXu584xr4YK+La2k5wOs8nhbThyWfLUnf
WWnPmmxCLsFNjiaaJ1UYaDtkg7PdXx1h/td9OxN0h1b9ZLBZCbaC3Zs1Rp5/XJYT
ywffxWSdwWLfwH0sVfFpl1rqyg7On8EIkTenDxF0XmLNuPVG8gAn42AMPZAfcu9P
2pEFarCv1bdAERvbT4u4+jD4YHPT8GXfAjg0kEPW+gyJu96bBVlUqNA51PF34yli
jsxn/vqRf0F2GR/tcn8zJuUw2GhV6DDXGMju0WtTxqCUq79B4vSaaVVV9EyPA1M5
oA34QrJiL+PI+uyI7yOQSXMpLHZ6U+3VVsbl3XR4/tnnPhyAxwhyFhyIM9mjsU+I
1zBhNzpJDlxyGRIqXLGhf2Untg9puVaxlRnSDJJuWwrHQsgTGf20+7QAcODkgr31
AukiSqLdlA0aaqN3zCmOvRbMsMXwyqa2Id741e1BssE/s+Aaj7FZVp4uvU/jgrwb
+iYShZ3Wqzhp0NJuLcxKOV0jFAGH68nwolUH3vAsiQmpp73ikagaIgVbzKWO0BvC
oCK7+i3tIgtR+xURYGq2qLUbnzr2GkI1BCplgf8d3eRDUdmLvnsrfWT7875dCW6r
FJY60WUwWdQIxyL0zYjqey1YJ3n0y8K7WG4FS9Er5S1hUmMr2IGX/WQ8+q3xkRm9
kcOb2lVpFQGjQax+jCtoiF3tRyL83QbHFskNIW3Fh8pcZ6NaqWcTzg1VGryRpbwQ
LRdWGpTO86SGk9AMbV2d4OZijDTW549sbxk1z8OUL07SW/UdGEAaQFUy/8JZqqus
Feaz/VS9vOSM95tMJha+XkL9o93VRkDgcuZDx9PO/+FQnis2dag9DiEfibS9U2w+
Rqqx+zKvmG0uZ11hR2ZtGZiQ0SzJtfwFKFOvPS/yxknnEAaucthOhYCMC2u5n/1K
thvebHRnRw+tWT8vZDX5fKo62AwWqZHO//AHYByJ4CmRJ8vtG+8vSpOP0ZBVK1jU
CbTXQ2I8Fj+6eZGn0doZ85gzMUW0CiKT5OpcDEKPm5qsONBB3d+4OTJnxxbk0KRP
UIsM5QXhisCT0dFWzXfXcS7DzQIyqynRAtPmsKZgCGuNxLdEH20ObK2+pqE8SKc6
3bSsQGOsmERVhg9za7dJcQgPYcmRYkim3UDbFZJPdR0G7uAdbOUI+l/ddC7gmPxC
Ow8AjV2/4uif87FMo8WiN8Bf2ipGVhHDgPAN/6dAxaFipUekF9Xqz8SK129+1G2H
OrPZdCI5izpGpRufP8PVYBtiw9Ms/tx20NWJxPCJV8xLXyfixgUrYHFX4/Bv4YAW
VnxMr9OdodBKdi3imFrW2TYg1okDSqvOEP/pc/B5WfMnOecEdoOc1DwA52Z1CXCZ
+6LSQLMb5OOx9d/lKzvG6zdLdr84Vd6YFnSLUSW10vjO6g7/SRa6FecUCvTbZPMD
zRdMOXcMbGYfPKjzLt619BmCKqbiBC5bzPeuy9V68LrGv0wf/LtTFXZBCa6Vx8xf
P3+vpFD9m8P4s2Yz+CmuAEBktX42MwvVbaMMF3Xb6VOwJFy/PnZ6QWGDiUridjyd
ocHo9/TgB3DjiHHrDyWM3qxhXRheaNjgRwY7YWZkOYhnhEnEjKlXHynzjLOIehOi
YT0yaWs+m24KEi+5c4QtelQkSjdMOrNfP2+rRh1F4VdwxRWF/qFG37Oy/9Rx0Xaa
04Zu+6ZOMNuqULOm16LO2uRTzYeP6KfeNuNwBGNpRSuMJcWclpu51+Wq/Xq6EhPG
1CadqaN9j5EUUGtlrooy+Iwvae8UpKSTD4Cw0nQ3CcSJbkW7mM1OrNrauXjQV3JX
EIJ8Qmi25KPvNi5SraA2eUM8x14hITfc3bxx3qKX8iPtV8H0R1IOIRO/FC/9Daos
7XPiwNZF0mRcF5KwoiZ7VgYJlfTrBIN63Gs0f8SeW6niFvb0yh+ReeLmKFvUo8cu
sHxO65JPqwsyBgs4kt47Bnkn9oAmajyZPyfO0OdgTk7mf423axfeXiImkVj2gaeR
aaxTezLHOTgjcfZ2sR8fBN3wbrD3yJlxp48PqFJWciS/ICFn8g4iJWE6EjjAAGZb
4hzhaz94fvXn40WyG7qGr5rfvdtHgPEjusKWZwmlabOsJEn7j4EYnUW3UFd3S+rH
umlWZ4E29Yb0Q0g5DfFXIhwGInkmLga1LZKWPEHT/eohVMGGjMZe4UCOkAjnU2/R
cty+Zd7FTNoHl9T4d9L4qs2/Rorr7JMzWIDegpFVrkVlovU1qcfBwTBxjsMRaZ0Y
Tu1HZaS5UC1JF+DR/BsSj93xV2VjCAWTOd/zORTMFmpfnWKVb8Pdl9SudTjiRvBg
mS+z5do0rjXaOYcxiNVJ7kvaiQRSeC0vtqpdUOxQVRXgeAcsYvEzB1TCHdgDWOkD
2cjlr/pjjtT/mqfy/urAhJYcWtn3EcuTIwXJAVr2mBZ1g4zmkndETZVb6eWcYHMA
E2xFCbiZxNjmX+R8cDpklTiDyifaG9zirGvdXRIiJB+Nl5muV3EaK1FItMD53Go3
a1pzcq6SWc0AsxhSTyPpKjmwuEsnOe/oIlMC0kueGo4tn2iMeVoRglMbOtwQ4Qmj
Ged+C21EUMr8+d1/V8nssNY9CFGGHiYe1GYS6gpUXr6iIUA+beOSKH43elfFMAlY
emkPNqWEMDjCcG+dDDyCD+RgBDYtLG3DaWSf1oAQCVJEOcHCiB84cVn1Ekay2Aqx
jpKXeggXUXsod5V2tqPk6Yq044wVtWneWEiZXbT2FpqaQErQak3OJT9uDrv0v/3N
K+ZcXJUhAW/98SjqwvnIstyvj+lpQSjb35/XzrPWQmK1o42Rc5VbLmY3+SKbnZZd
OvHollJukr/uPCrSpWugm+2f6jHpOW45K8XtnnQpSV1dA/rnJjOR3np+9cm0sfT5
soLCCjgtXFtge8/X2WBEvoaQIPCCvq6ZZARLYITiggsZii1NvlnTug0cCpVgUAx1
um4lpSWCZfwO0wPweKprhLJFLcvoHejQPvoA74mqNHM8OzWf5GOy691ZU4WApRZx
DG9mXq2qhyIs8WvT2/4QV1shnnZ2+8w6nuMdQ1VLBJPVgHs7IbPBfoKskVeLVSmf
RAzLkH+0SRXNdvBi30yOWdRiWSi2GcvbhTP2KVR+oHx+Awk9gzDK7OGL5PPaJAx8
vKum04vqUvTgDdTzPKrqGOCYl516FEkT2QDUnwrFiJIgdTPfX7ugqH1+XjvDSiFy
pzAyrZnBJ8qFVBf29IuzLs73hz6vnKy96K7ST7hte0jrGPa2X+TKaVO0fBjVvV4e
uo7mRCKz0NC5jTEozP1uYSbeLAFIcKuMDEWOTHrQbnSB0VALYNiaRZlRIbhPrvkA
U6fqVQRdw2XZ0cVSEMh42+BdhX3guIrLUvOyC6uuoEEptxmudfbMfwysP1ov2oev
bw27OrlOVVkq5ZJiB6XuO6aAY20QOne5Wq+emqmE2yke64yuovwPzdpNyRO1nnNR
3iUvjr+5UUBGTxxReEChLwvE7lwRB2skYe8EiVkpHjA20K/Sffjgu454NTJZpP2m
WRSc41Udd12XamZGl49aVGhFIyKGNEJ4dQEUdp1r9QPDE6yidC3EXb3SQ+immRay
Jz8MBbNUWwLHvOu2peMfOaXrabMEQJHp4ciCQpblsRK4gNEw1YzUOayA3Jhwujf6
y8NKvkUoRgnOb9yAS/4X6f9Ov7VSfCIND7qfgUw06yFDXuUdbfdCaVqbBxvfK7r7
GF5GH0YU9dDcApQuFPBxAdIdeiO4Jfkqy1wIhj/KheHhz50uLeO9XPqPLHFJA5Kw
3/kiiTRlbHgVXwLS7Rmr2iFlPQOt/+00UlCxR6kQEjZLsxnD0fE35sEj4J0ty52I
wVGd+3S6tjN9iLQ9Bx700rk8/PbiYwd6d16x9nxS9+o2TrImHqIcjjSHTZhFdVQk
xGo4i1PbtO60iJMOXsZSxfN0BVY7R3mNcXsPlAjErsMhxwlAjpO4QWqRSvMtNGzJ
Rl0j9CqM++eG71gBFrOgdaVpKrt68KAC1Dpu9iawtDc4h5As8pPc037ob4y6Mapo
Wrsmh61h737+XJwVnQg6uQDoGn9DjXhNawwD7r+OSi8rVex/JYB1UMTZ2N9RDxcm
ApHJ7aG6+OQgYjrH0/77hKe2/guIhYoxABiMY6P70ibAVixGH774T742PO85yb24
376lNCV6kTeLWjCSPCxlGiWi524RP+RtQ3VQoK5SInSgJZHOIjNuN9IBqrK1dLuR
nR0s/IYUyLOxg1X8lqaMyFtw0y6PeGBomWhVkpVFc9HP+uPsxL4bXadM4acwk0tE
D3PmCpeOdxlK3r7KjN4PLZqvCB6tnlr6osQzp4fkBB2WM77RtBUmf1juX2AuhFQV
N2XXOBoUJC4LYesLJQC9UIUoPFmlIkEWXBZboOcXHX7ki3Nrp/EDlO8ur5YKvVCB
8nbblDIlDVhkkvHou35tAxiE4SqG3iMRRjqiPuGSxtGCzyqr2dBvzxVb2DfEo2Y4
pTYKmf6f//Wd0chKXr/ctHfCDTQjrktF8Ofd2Qd9IbZkmHbWOGeUpIQE0ONeBurG
DjNWetyZSS91S0pL4CNzyRl3ltRG/jZas9OGIr+6h4dqYAZ6/uBCT32x7VNdYI2U
Gx1fdK32O2UTovr1RjB2ErxAXscgEDAzlWvlIP6kxJ+rtIKueWNGlZekMRShvt02
/buhkvNYfql6miXkZtHF9iRdqbg53U2hivOWFvGeCcLKMKNQnrpTbIpux9xyBS3L
q3xw30y6Tw1/Rw6QbNkhqg==
`protect END_PROTECTED
