`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mO+nttEO0qabG6MkHSkaIigP7t8BwqzhNL/PzWjxi80bMacFmmJtlSv3y259JBs7
ocz5w3ev1jO7QdUdmG4B2QMbMRDuSFugiPNDyXekPPkhmE+ONVARD3M7XOKXO51G
dd3EkyLlVeSK7FukoM6/wJo8fDzpPY5kTOyJVWqy3EWEdcSMd4mxQrLEpMSxOd2I
cpOpdoyzR0W55ZBkPv2kEr/KXVBxf58pmJoANswTTbxF7rMUmdpQOfk0VKH/GJKI
bCDucBTKLUoT3DGRw6q8m3FWHiebshH2+8QwkeOeTyb82F36wXnu+VBkUHF5y2yb
f2OldkNLpCWaJ3SsWsFXcA9oXnz8P0kwguG3uKy3ctVg11ZTyyMUPBuYClKGIQfx
5EQUg+XywjKcDmw3AdjtFQ6dbrQGIMNvxg695zuj3ihkj+c6xW6PD1kLflxjl3dR
`protect END_PROTECTED
