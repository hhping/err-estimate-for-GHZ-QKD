`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4ylJfhqW2WWs3Fibz0cOOSR1d3/D05pWwlmkCVX4JWsOjLrMzi7n84e1uGu49/W
wEvBFEVWsJwnH2Dh8P1ZVZ6Z4VIqWOQ0BLEEuAysvG8jqGGXP+lYClgRtk4T7DsO
bJlur/JWgSgJKgZBXrmLp9owr/atvu7FOG9mlGTL+EMCqN8wJB5kv/7n8TJXIdws
EK08ygw/+0OZf3darsJ5ZA/6bpxyi9MZ2fDwI8E3K/f11QhuAahfR8MvU9W5phxX
gi/+k5x+6TscAquMPSSXWIg4+5GCizbysYFuz56dFEeMl6PvMCm/8AFPKB3khT3h
5Ukpw5PkjrWuBfdVhJBUZWNF4NE43UwPS0VGmmS/IJfkC4cvo/vNUAaVoESrwcYq
5JiVilZAB1VA5j9JryUTm0QK53BzAAQVCaCfRGplDibD59/nHKywdvW71bVy82Y1
KJrczI52jhegM6BXOw1fX/wvvV6NFyoJz4DbxWvS0go+3KnWRs55/K12aVePRrad
6PG/t2V8e7E3p2AtWXrcKex2VlMEL4IHUJJM4kYFX7hItyoLCb7tBAgfxb/sk8oD
40irzBrtBpww3fZJxZyNGo5hl+OF0+HibOevzs/cUggzynDzFGpl5M5SnjbIdUSN
pUaaQ4bF0i0kwKq9R2NcUsv1CxZiAjDxE6Z8BUDRZlRwE5HMRc3Eg6SNyQ05kh1u
aXBJIJnSxuVao5vZvDur+LXS8wVmP84fafZfmcXpKU6e/UVc5kmb8hdNeiSzwoJQ
YSomqCv0kuNQFKrWGsxPY4Svl8AMQKWFnCzHvTaSFofnoA5K+Tx2r+bXLULOtQPj
kJ4o/gECNlPB/BXyUh9YMMUThlXxKhA4quLGll5IRvpb0oXkfG2sLjsg4Kk2SAYz
7kb/3Uiwenjs1D2lDmQE7/vj41vUFx3u9KupPBEym1mR2EOG6v9A3Gh2vSKW75f3
PUn/0YkhVg6jRJ/l95lLZGjK8qR9Lh8K3q0USyAC+raQYLNE8ikkl2vK0tltmn/3
cFzDz/T9xIEzieTJ7J5LEp5Uth+nct3kPCLx9XHch0bwRLyzAfcCIHKjw1Y3pwqs
JZ5mLpiIVE3x2wdlmLLwjx6bhMNEorUVfvMkCDAiR4MGWg6ShtlqAGuz6mmd7cGC
CKkE1PeXw6ZTy4kIf1ViF3i3rj6utkGHLkW1tzFHSP26t6o74dqYH9erIUeJFymv
q9mGlrcpqrg5AxUzS09Xs6oYXknyL9rnkVdf2FRi6KRkJ0UeSnFbAq40xvVaRt3l
YrPKshlqb/Nu44A9HUb9R45vQ4gjkX5VCE+++rmyyymifK+ZjherRmXb51lDSTO9
Dl0JSr/QF7FToG3Pwte/mCRTtCvJOebZXKHKhXZNqOYV6EqMKWy8RH8RUB9hpGOy
4toIqOgOSReWfKXq8zCYLDzFzaruziP9MuHzOTwVN2eY63sHolwXTjIVQHQhypCT
5cCdZ4mgF6tszFcFEEMR8r8WoEW6UGHfr3iNrq0cY8n3Hk2DJXdLs7EUZL7tYSr3
eAyiIhC0e6NM/2AkUNdFEvIRrO67mbwb8h2QMuPCbs42ogCeiu/tkMzcQiBSyCWl
hV5PgN4lXWuBYevKPjSgqgV0hVuT4ljwlHy42xJkYZ2mKCJc26m6YYekmVk2XmA/
oNEtai9Akohx1s2cgLF0Eg++k/VaADtO7YiLBYDmXZQlw5q1h117dZ8tIpSOElTZ
8yC/4K2RV6Vy6zosLNtTx6oqSzNlWwcRCy2k02+A5M5Xm/lBDmRKbQnCnB/SmgPd
`protect END_PROTECTED
