`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zHZ872tkeiok4xTmebUkLv7wz/lL2uYnSISoYByhrLnC9K9ArRRbONdMh0fxIyR
MhRKOQw7q3XZGarzOGus0dx97VI5B7Z7+dwXZmzYmb0HDMGKjRo4MizoFzLvzR3l
QJVztyrt+hqoNij7ThcuCqQgATYhhwPhKeVg9xGcYtRxluwwYNJasburbdR1HI7m
X++AkKu9TciJduoNcRNDDMJUquR+3qZq97WJfZ6GCfK7z9HfxHfhL+zX3IeXCipr
OcMTGHlMIakqyolospeaCL4mIq8b8TgBnRpxPG8i8k6aBatp16O+roN4NL5MWkiF
MVJ5A6axPsGTj35mHFkVse1/IcD130xekpxc0dZgEfy85Pdb+n9kqYop2vbeim3c
BUpfSYhKVNNzV5VG/di8qNP8LbOgXNsaHIAtGES2h9pINaNHD1ox9XKs/W79XRuY
t8pVTq8malTSqgnyPb3LbWEpbeXIr0CMwLsnPzGLV8nDsM/HbwqRabDNaAvstULi
XtRdEXLZj2vA+MxoNSLM6J8YtWLUTXwmU5RYlJiBxBiGX3e+f/iMH2lVyQer69ZG
PwnZ05mCxgx6Hrt3TCRljB/6GGLXM2cy8zJWm2AsrFe9EVaAv2aNbnwhgcAEG8gw
1XhVy9GrdnBmWU6DLXF0fbCcoaNJjWwIB66lzGTOGDkFZDt1hh2VrVLAAhUWts9H
L+x/B9KMkUSO0BVsb5+WOaXortUdXZAeiqNwcy7iPCU=
`protect END_PROTECTED
