`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/Ul6u/9fMh0/vbe9WU5ekiuDFzYLRwV1G9jfZJMHgHjH1pPWpi+i5tIRen94dcB
vK/6tTBr6S48dB7V7KN0o6xRpqSUKoIlFTayNNEY3+Z1Bc74pEeRRXsZbVzdnHMy
gaytDChB1JuCTh3SVeMNIUxt9ELlQtNZrRahxzGesANdE24+fuNvVNQJoTQX+Pw1
nXue2iVeorw1UabzaEqskhLR0EuqBglU4Gzi7+9fczLsVI4jzytwVJjP5by6yYBY
LC4rggGZPRHLxIwYgxlKMs5T43313AIvBs/Xk5UBVo1Ta9vXb3sIdU1lHy7mLl2F
mvYFU3VNpNcpOwGstVRe6AFYTlYtJo072mO97Z3A52UHLRTpoTReGNe8eUoXwB1J
ilrk6RywuXWicCspxYhOoUUGZo8U/ANXnA3x4f/sWJg2y7856QYGvjpBHhOQNhFV
z/6L96Oxkwy/xMS0ADyJ57QT+i3K9MZI/n6EM1OWivRXEX4wagoTeWaRAXYhvqXI
azP0eZIOb2ewHQUSHxJc8jGiVzWBt8MOkyHcDp9DEjWAuVqF8fEwQ+k8a12T3dvW
m7/69oOJlrjZn40ybj0aL2TTeOLD4eVojSGhfcGKp7MGZuiPONir7VH1j275Ubag
WjCBEv7+zm6CBOYWKA846XE4DuIqVBbAYubVJpxSioxAg43KWlnRD9mL88DD4aqA
c4C1yYp868kBwNMhP5gX1SaoWH9U9de4pVcLB1APGEKlLhpZRfl1WVrUDA7BHBRD
9eET228+puS6ZAAIp9/af2d6FhduqAzfxB82Pd+bSzYIKi+GBHB20OdWP0yKTmVY
IuFjgBXEDdOc2/IqQ6VNp1s0pG+THY+7Ne97GOFbh/EEaf3PamZxUObzBRF55nNg
8+cpZOlnewT/GrBcTEnsMUJ7V7Yoyx4OtFnM1di6u/DfeGPif0frGWRrxAZfIUj4
f38WFrQwZ0lRO4boUY4H5mc/JhZ0ssItCkKI+IbltZWmLLU1NzoWFIsKl+NCIYKw
Clx6YHyFhRDQ71tWK+jFmQrOaS1CquNM5D9dJ1/s0+lNEx41gCzQpPTsKM1gCWGv
d4+Yf1wbN8BCQ+pkAFkRAO8AmZJ0Y79NfrwzCf4OTdf2P7Ezfp6QKDDofG2SqD8V
A1CUFcmNUN7HtK6RdFwPZx6d6pPV8wtu2XD1zkPAU1qQ0n8cqcvhQwQo/eKZUWeD
UC/lAB3BOBSvhqWJ40lieZNHHIoPZ2vDDmRQ9vPZV1R/s8OxFKV/QdhY6xD4E4Qx
zkA3fQC042N6dXfQwLsdLaIN3uN2kMn8uKZCE48LSSbSPQ5Gw+zTzX9Yfi1LSBGq
GuvhXV+sHrexibSNTYb+6gfokguxR6EJ5916fdMG6ggKg8HdFCHMqS2F5M+XX9LD
dpEj9Vl/WXc35H9WNyiLB21corrGnjCNAv55cwcOsfMqMeKLLsfsXkPwlxoWQAB3
qPWuOPfWHp3E2Wp7v4giJ9Vkfkp4lT0AFKdqydCHqP9Tjga1Nt+yZKNYdqWXlQsY
wiCffzZsi0OQLtqaf437/fgEjvCUJNNzRdz0Tn1EdyRqvK2GRLubJxTonunKxO1e
fwmDgNTM/l5yw/Q/OeJGL6eX5wTzawgRNl5DZiym70l5sjGAK3bGrEYItdm53+JQ
uh89lMnQNoWm2Q1jm0O6zjwofIx0TVCHIK/RUPh76PSC3QTXEwqyPKTs8461TXF9
fPUqJ+jIWeSB2mZTtNKufQfwKuX8U6NFrdMllrrHckJltovCTClX3ngBKH8fniIG
hnn3B8z5G1ZkpG/DtgwuvloGhSoW/4H3nBs0lhhDFoqwKf1yHXPKLaEnga7vCny+
AYS5moGfLQIAIF5yKX74p3QVYnmuTfgZ0M6JD2B8CuryeXFTU8uns0EOt0dUXf03
ZaG+K3WsHaPG4e7AUr+yP8H47/C1rAxsg0jtXYR2DWPqvnQxGl/eOW+GkFHfdClB
ieQydZeruBNsnp5cPyTgJW4GXU3Rtdh7UtXAA+NRe3Xi40cF1QK2jVWRGjYKssw9
9pRmxgd0RgUMHjJaCh7z+sgf/M0I50rf1vZUl4Bq87SbSwH+5WSdTR3jhzYbObd/
OZ0sJ2/RHv7+8VNwSW8c9tZ4BFzDWqNNM8KtL+0+EMcT+juZ8uL2iWZ5+vatns6W
+42xZEmTZGWKFxjWYKva/jm+/KrIYvVbOOye96Buu1C+rIUSf8kjjSKq5BxOQ9kA
gDlb/RUamfsX1cyUI4ttL1WrQBrEZd5oUxsug8B8dXGF691T2BegoPKpIkZmB5Ln
CUoW49I+z1+5tFUl3b0pXl65bTFxkYwB9gxu6ry5idI=
`protect END_PROTECTED
