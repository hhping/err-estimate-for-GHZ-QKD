`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axPginurUO52yuvlVoD4FjHJdbR+XUMuPvkNyvXQKbWcpSWANdDil/IvLBKSXNrZ
vxOknLfqi53Nq45UBNrcc+IYkp0sjlXtaSja2M92cIKtETOpHx85Wb8hhvTMQ4dD
7XlHGLNHvaUS7+QjiP7PZvon/qYy3mRZIfLkDwGTEayEmzpDfAvKtFNdaRghAubr
k8QnNzCJs5tg64BOUWHVePKshS4UpI+scUpyGyxTcLiRgBWx999CjQc2f/ebkFh9
yPRCDYjaRr7oR3alOKFr4Ndm4DBQZeGhAFniKRctobU3ReRqSEWSEbVPKVNpRJK0
JMEvJfLPwVqFz/QhNInmdtozHCwfUSQT9G1WQtblFkm0ifKdDXyrafNW/o260BPP
IPFBPnzDiywgOs+EXoudZ9PNfzewoVbC1PqfYppWBsZNslzN3yUXQm3tYk6Nl596
VeaRz3rhe2C4iHAjVRm3w/BySnLxF3Kzq+bqps3iVwZ9uq7oSijEBCCmuUznnyyx
kcWnMYdNgMDo+Z1raGMcbvlAcMXjijjnThdSlOH1zqyrhLSs51uYS7ywNSLtE8P8
vToECWD4qBlF0MqrBL68PZ0w42f6V2g0ZizcrxizQunGPFZTn5lxncHSKG6T2sBa
dOkGjsBBZljAH6YIXfrzKqSVrOMWlufhHPP16MU4P3Ex8rB8O1cGpLKEIA0DW63h
VgTjaW+R6s36HwWaYnNrF6guqp5LSLQUV5Z88ORhnLNb1xoaNpAIrsIw4c9AUZyE
sJEmM9UIvfhW/ohRXFQbo18AhdlKh5Lzmkw4c+HpxdcgYSv/jL9Chp8lagRCQkpZ
MPvRS37OyzBjoyTwqOgFW04YqFkDPX8dnjsPijit6J4emEsOB4Z6LiY+WMY4367q
fMcluWcN+ynRS3fUsItF/41juvIXP2OfLvgl6LPYEzhQfhc8YKFYqo7TZ8/UPz/2
KHxbYSDcuLlaa97wO/hW4/2bgcda0LbpDLmbijzPfokylz/wocQ2SjELpRa8s7UP
6gDx3ZjZxU4th+lUpd0dTCyz20b3M3ZuRXwjXM0eUjVdCHgqJUXBVcwUYpuyrKlK
3+dDJU3OJNCDIIeATN5lVZhfK59Cm38J3WT9T+8RcJG+hvCVhcFhwcS4nOTuBJnc
xlISrqReW9Gk1hnM7sBdyhqgRWHv2SoCcaCKtDTejySNuLuJixtJYxTwfXeCs23j
KxiTs2GRSHZD7hHwUrmTDzKRPoSqzsssnAaQmDKQQpFhDU0DhMFaXlGm/CM0Cbee
mbE/wKECCm0RjtQfZ7INoyZ063QP/TIo8k0/Onj9ifqhs3mqY3VEjrG+dryluhRL
+ZcvyxyOxDDfx2d1a63c2lFvKWEkCty217BKCiA3APhWlUmyxuH1sD2NYEmR+Vpl
+VdMDDK9t2J0RSwEXZ2vjH8H5uzW/MiFvJn+KOy2NRyMOFIMyX8L4XIUujy3wIuc
lFCszTH5yER0bOWFnMpC9R/hp40NgJ6eWp1InzgSZmtvae/ifx7aPtLKCHgeNrmw
zbLbdumX7/m61WCpfrfRKBiRTDTM8KEf7Bw9HSr5tjvV4OHK9XqRhUVz2qLOPoWt
V2theuSQN1tmTSNphzxiEQB0RUE2fl+lVb1j+6qpww8zb+T8JJne1XCuZFrbGsud
r5Cy2uRb2bwUZie5A9x8b9QUOBds9uBRp+MRTOhB37CuaDS+m6eusYywI+jPoNOL
/X2zGSt8eN7Vt7GMMvQqCmPPvOxjWY5bbQMXXe4Y8wVHtyq1umu/1xl/GVO7DVEJ
`protect END_PROTECTED
