`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hy7gmY4ZoqbDPd2ioSCYV+WJHO5I9zTNOsRngEftq0aCDthh68ekFU9JlzN0pHJO
U+G99pnTcXh2/t7XvdHygsXwCGMPpGLLmI3nHvZrwTRrSBxbEKAlv2WARtzSd9o7
YD+FG7PFrXf5EPVCiNYen7LUQMd7JSEmLW2y70C7wpydTNcNbo9gxiNcFTO5KtMl
cXrIXSxlYldp78cUKZ208AlZZ6bOHomO0RrOcOMwvYBWiybaOl9oidAJ+1AYt3ce
vGn+9OPfOw/o/d6Wk/o85fVhFAIIj0/9Tioh8U1b94mddBo/rw/X+mzzMUIM20ke
SdHq/chAQrL0Uc34fZOHNVCOO2xLgbr5MbREnzryKeybgeRqzQj8P/kFfZKyNo5V
LpNs8qduQsJL1T7p64DdwNPX6IrrRAiRSdkgtw6B/VZCrOnhZvZEJtJZabbHu4rn
PRj7wHNL1DpeO/kvAlcfGSQ7goHOpppKuCf152KDrj29t31IaqEFRwERVICTgQ7I
o881FJIg/8UnS3sVexttEJolR0qkjrI6US4+JiCIumHF9CJCpWgpYi24IsXIxgMP
iaD+UCJUztWRwR2EbpT6bA9mZorIMiGz3cZc45GE2SArm4OkniVYrh52r+zWi0Ep
hvLMCQLPJXDOeIh/OaKgQTsPU7Sa2VFIfFNR/o0F8pPCYZMqXHEhXRaA1VU2USCN
3d0G8/w6H1bhggXsHHZO6ysZXREGiEaY46pBBF14TVbmvpKiAC1A2TdK9PGIBLpF
qCZ12w/HSgcWAQwEaH7mOgX8/l/EhlPUfyNL1IefdPNI1IOHOuWVd2MFO7rPvSeL
f4yHo00nxllFg8CUgLULYgqqCG5sy5p2OThCq8Y4/GEHyvfustNqpKBm2LLXA1GX
N/QwEC1StbNARGHrW+KtGV3yOVciPp6Dz8l/AxKKvrSd8WtexG1OxjqwT5rjAvwo
QDYrKASafOhS5CZ5z10MEib2NFWuWCovKjZmDekmfjoemRILQGqWYyKXugDSeRfE
W4AKUWc6bnIaQkfY8WRPE3TEn2zkf5+r0EACyB3WCgs+eWbOfohBtQrYTVExtXfi
EN6V3ec2ah4llqhEv4ofwNRYtL690t9qOGrDgXe7LJS91BDKe92kl99ewfPBOI9w
ojQTkDc9e3onFl7fEvzdyx7R3RBl+zhxe11wZs4tfmtTmwgXdWabt8yNnvlA7maF
L4M39Ga8cr+Tkxm2iJdqOI2exonmy3SxlfbCIIELHSVRfPL5tvCyq8016UXoMXHe
eRVqfRYHgIvLsgKSQGgv/DHo2M47Abg8muuWdtQxaJ5dqRyezXgNNKREwHAM6hFl
0noHBf0CjU+h0K11MC8AJ2SKWvYeRcxvQMHD4v1t41jaaUtpPSLXSzG19/GQTWdW
fGRSqWDvKI2GEn9iQZFY9oH8gtPFInL/wWxYV9QGekIJXHPboPapLZ+f7+Y19YX5
/lYRZ8dL5CJnRrpAwzyPlYIjsP18IkP4knYOnY79HEivjaY4LaLShuSJNYvb1+tY
c5f/s9WSKcd/wlbEzo2PoISe+5F0W9NJnkIJlbVCMf9yH3SMMYSSc1rS1TVwbcS5
6q+poLMTAwLaW/Xb3uTnGo32M+G7VqbzEL72XzFTTii1m2GRN9GTkg1VhZJQYz4Y
35Y3oF9LctsUB3q3JwnZR4eqd9dleBbamSyTttKlXHcew4MJsqnz3l5H3p8wMOra
mU9mCBGjpGvHdvd5DEc4DE2TzJ8IGc44A5MXOwBbQzqe9W+saRU9n1Xh4/8pKthv
LA0eD5dlsyPhDDoJL9g9SG7n8BUTCewjNkMtLvs3oSyzbPlTiFrYS1nK7MSwPGvC
C71gs5Z4Du0nAoGBUEkwPBF/6P7q9J3SZp0tdFSIbyRxmDAWmWnEkwRkMndp9v4Q
ptxsWLVGx3TfYe29vwipZV5u32xeP7Q8DqwAL7wqbTME3dJtyCUtKVdFAsjfJk0b
eDJkdMc5RnINtDTmFf5EzlvTBt2K4rz9bCnvpQ4alJmI4F4APSqtzGs3RYcOCRHD
jdLek11ER3Gvin6hpD0/DfNMGMRD/RxT4fCD/b6NaRPwKlHxAMnWK+5c6gLXBwC4
5Ur+/mLpsT1QLUhhqUGoamglgD8LE9b+bmwN5N+m9idz9PclDK3yb1mCWx5QU3bB
7gStE+OOimUdRI+ck9wU99tMet4JDtujiSOl5AEsbaedDc6cw9QO795aG/WO8cZf
JB429pVFdtztQSn6O+WyQSHqK5/TNwGQLna8iOSS9RUJuZ4blRIIyXNcV0oY87NK
LbXKeFOq113gYx7TCvk15Z0Kni8TTVYoWXpRRb+AqqKAUWpkyamBTf4kAD86UFbx
bY7FASRPR0rX/BfYEncqlrRABD5KsisA3xrm4IRwqwGzx+2bBavmeyCBGUndSFDe
knqlqUoJVTLdK6XvwIA4Mr+PY1nWWhqMVAD31TkC71tgKaq3BOXz2tL3l2+FqM1u
MOBS7ig3FtEhmPTU/BdJoD10A+zW/Kb5wHBzKgTMXbcNK7hDB33n04eYFYG/wH2/
k6QxKFFe3A/A+G5t8nxCyJAofWWz7TCpfDmGKeTUSzhkk7y1sExItxDk9XQlgrnQ
eCit6K1K37321QeZTTYT93l8Dy0KHzsS88NhcPWkHWNURLKuOI613vuDG7cP/E8T
rtFJFs4KGiq4we8As9h/QQ==
`protect END_PROTECTED
