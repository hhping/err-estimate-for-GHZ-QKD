`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oEiIIs2BwFYlh4tK/pVucMfBOJGKDBmj4Bl0BVwuJ6xe3zTYdTaMHt89rNShtf7D
sQ0iv5D5ADxfi3SKWKlaKK9dOKVbZZ6YiIpYEiammYvxGy0io8gp8nVvFmMCC+L2
M48ezcIV4DdA4KrI+Oxna2HerNhjeerhUaiP7sT6AFZarb0z9Y9SA5h21M9lp3dC
5e2T7Jp32la02kurDobF+NwgpQuUKghs2dnFsQhX3ZtLNK3xUgZEvjgCJkcoadZn
vxILeM4luQ8KANWfl8zSVvT74Wca49edVRIDkd5mEVUDJlAXADkfj4JvBD4mUYU5
/pDtgAumo5ZIyvcK9MpjNq06YCLW3AcCNY6GQTEnOQwvZBmprQhWZDiWg/G713eX
/gHbEoKPW4jmBY/T2K2BbxiXXOKn8HxYVY5sSB+yUQEqE47DgxZoJeAl3ThF6MQk
bzcvFaFMANnY5h/CBUIVrBEOcTGYyFuFSmvFZrBnXReWlkp+zEH9HcPql8PsOO1e
3bwD509Bg+aplLRYZhgoe/meEeEVnMr7NaXFzXCzFf0+ohg7WfsVPK3H0ONISP1y
6A7MuXjRWMHBS5PmUJRtgrxxBZ/pcyIPl/syM1IeQikzXCK4bUHindOmaivasjMD
sApEI4gbDayFSJ1OaI26BP5S9lpbcjbD1ur6CmF9tm90I5A9Kaqm2wKyTJ6aNOzP
/dihTcY0HUfm2plsZ6SULckfvo+vZnsHasLi/zfSm02ln1pGRtfQ2kgeSWUPthPz
0CmMLJKIzf/D4SdtDCzjHgRIZkDbO49qk4HDeVE+L1grbuBCBx7Qkuw6L5L5VtbS
SQIe8aLu5e4CNCGYgTfQDSAGfhIdpS8rNylYYgzIxiw9eApO7/gcwcIWLbp+mOil
EwurmOZxvUbl/uEg/zON/9qcoaXnFXzZtJ5e6LQDmD5dqSqZyex04JNkl0qmqT5g
EJ64bwp5Ls9LCONG1oNI+88mlROQD/sOYzxEGnk3NbiFri1Q2ujtOsXctq/tcVEq
USD5QC0GyQxMybGzElAlWuStJGx+zoboPtcsK+MjaypTQYxkRL2t/t9Gw4+D1+Zh
5jEv65MIcwudChaZBat2AMGIvpqxrgqQDRkw4ffw3QrLDlO4tAoEDcgCf1yrIwXa
inUIBhS9OzIrTG5wp279JpLfT5UVIWCcJUr2E3WYuhk5cr6K5mmowTXM8xXdw6yL
tBQNkwdaCLrG6pqlP6tD7dvv661PigPR/fITdsgwXXiMvM7meifndoqn7gorGgQ+
D3ZgX694JoaOv4BECOJuxdxk0CdQNfI5GwUf8nxPLfDDELmSHBqGl9wvyzcEEWky
Aj78/lvhEOpW3f9OEDxvcGz6jHjl5UH923lkjPZ5QF8mnZkgjMiyxpJ528S44GYH
dDf7zik47ZV2JNpnNF0Uqr6gSVVMBiybcIWzToLJU6rWNfxBkU0pD58CnH196XmW
1WchF71wwmayGwdmfkf/DwoK5s8eG7WYPMOGcYJQDSzFC+iqDW4I34SRNfX/BpRx
/YCEgQglcTbPyPvpLejaDmDDSWkBdnMJ+v+jmYGFDgtsNZGjBEsyPHHmGsWsVfSo
5DYNv/afPJemZFXdUhbS/WPenM0xNyeqc0lgZc6Waz9CnJUaTriGLOY0YJUhJcCp
xHB4eCsWrX4ieHk24FTwOXJmrXl9hT4pQF9q8qYKwtu6soTdN/msQHXamDzFLuRo
AhH4nRu/PoSi80egCGYc0NkyOnUPSusNwAspry2A3eaD+h/hUahikshIOJ9ezc6K
6/NG0XEu/otOSsc1VLaYMSNKeaOxRG2yEkBc5pTWRuqBJc1OOgBLBMR9Pp/n9X4V
iEPNhSugHVyl3D6hdBVxhuF/v2wFkufpdAUtsa8/EMC0CSYt93VXdX3jPR6rrX/L
wYBzlA3eqLx9nja1MEa6kt1BTD2A1sZYwJi9rPUGqAMqK3SaNnwV7cHJI/zXSS9j
Dyu9ttn8Af0/gQ3wUR3ErRKST+J0KmFBSRW6l9uS2E6c9bayN9RgM5KA28WJ8B1S
R1B9nqbfvYYLVSrgnZGdreXWBtbgaMYX7M/yz748BbTwWG7Mg+FNDn9F02rLBsLQ
Yrq4IuHLPC5FLudX8jKgWSrtMJdljSI2xk3LxpyEPA9RSC0Qenlk9kGfx+1VdrsL
nZMzmnf0ke7kHTSHKUFkLOQplx5QL3RLwxExtXR/czQ41UsDg9JbAMEIjRZ5A8km
1ovp/Zj2A1nnv3jtBEuDcV89nKVB0x8LGcCWXkmFe7jgZER2yTOVjl/z8RQ0QEh1
Oy9T15Zbvn6wCwPm2700ES24vJfh3kSzyVRYON8w35nPVjEypx/SZ0aVaJhlMKPp
nCje/LmP3QDDCwlcuVFsFuff2Nfng3Hsmzbv0c/1iKJ59u8OMSSJWg9GkLVifubL
b1vbPeGF7nT0yvK9IC4eZzUDuISBx/TyoHOWOyl78jm9LBOrUu2p103YCm/eEMwN
j7/yhFFH/XR6hNiFXR0HyIUZiz54buCpvIPDpzKtD/mWLqk6OyjSuB9di6T3aNXn
1hAgUNfmzdRaT2O3TcqjQ86RNIK9tQIIIIvdZSEtGFFVL/9UJChS6lNDAAggSUVA
Iz++xswcg0FIbOtDNSp9QsDyPyQhrtsHf4ZUb0s8ncmeZciJsBnY5dpL3dEl4WVJ
CymKpqM2YkzIWzn5WdmCFROzO599dA383r0h4gR7vUKAB1LQxO0XegYct4580e04
+9c3R83KvfstZ7oDtq8XY1olWRKvjHuikTry5RjcsAHH9mlNZ34WhjDRum2MhC+n
KdKodKggdYCCbmTebqmrfMRHaZqyZuPi6LVXmWfodnpubFm9LfD/iBGgcyLI69nX
VJv2IDHzBKB3DGBnTMbf9QrZDsM2QU4BcY+kdozO9vojOs5qm8aR87suXMH5uaka
XvxJzJ7SK2AX46cMXH7OLBhNBxTCflPHeynRLp5R6LhMmP841I/qUkIcB1wOcqSb
z1YSEcbkGQuTNnZcVCJrq1upfht+Ls6puKUlR2AVlloxSnfgb9+4BcEJ6ZQFH2NA
BOpkjwh2TdphJPii9uLBFnhZTiQmGFueQIwatsTo1tyb4bgvgda/jW0T55BVZ7BG
Yo94aoZc3haXAg+LBhqwnaxJtrlSV/TiuAeqtxcp1pFcGU3WSXqAiqF7MumrAMqB
bYBPA1MaJK9Z3D5r8d+HLXEtzdmxs7Hn0BTgap1jrZqZoeURh/IbWv+cjGAJYvhX
Pd+0ZhSKuiqg7hVWyOOXacTasX4eIPGwj4NgZctLK+C+OpYYkgueujCJziZ7QYlM
oQUAHNetrddkaImvU1WbwqPxZCAwa7+3vvkNLSMZCK3eTV7//FMqqN0K78NHN61r
QhA2Gk6LxRCIAXn16KGKTSq4vnyGgy9VdxEOwh5o01It0x38SMpzZywIJVMkuObV
cHQ9fS987C+68bbYVcxVX6RKeIcIrLzFRaK2CBoc1NFp2dRRxloXy7jaJSVaDfth
V43t1oO3Rn4rbGwWTgtDXEECEb6Cg5deq25rd+BW/4stsnWj2otHfPLdVU3mHX5c
td0Pch2+oyq/VlT55LlZhTKSJbfKqehtc4H+oHIwEWOFUtDQh++epgQOncDrKNrK
XPsuQCzjJ2p1ApEItVEPcAMhqfzsNvbXA+i3sVskXG/ov/sTDdLX+HaFRAaT5Jlf
BoGBaO8rwgOGmfeMDTBeGCufHnsQ+rJXsblcrKMi33zssI0uvhvpxeqbzJiLnxzj
26zMMqWiOmJAncA3pU3YR32iS9bX7RIm4Si0i9oha8K34D5SBa/kWxqMi1sZG/ZS
BDgfxB91eOZzCKrJIRod5i+wZqn8/hmqp9kTC5uYYsBZUSWwNcTw0FfSWTPZc7TK
5UXnanu1eq/WHOkPO64xR479R8UA7TKsXQ54hpy42c/vzJ4gU4axfS3RiJNO4RsK
wqxKONNnClG1ewKzQWwxi5y+dSgWRWuUOM6KKHkIUsNm1MftPR+IJ6yvvqBfCu7o
PzAtgDz695pT7+n1mEhUPLL0WCxIqBFDRu53YSR6GtOlCbsHUMgI2JxA7YJCD+lR
s+3gtRrPvet6KUnIrMKlJWQUI9eI8iCw8BJOEMmJJe5KZneguEOetE5EppjXooq5
`protect END_PROTECTED
