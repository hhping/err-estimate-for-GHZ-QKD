`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pL6n6zG5vc0AIXQixdwrWn/piGOaqI/rGNtA1QnppQDTWDKB2kwsWisZ4Ux0dSbj
b1FevDZVxM2ZH4/1kQAbzrqPDPEI/WqNq/CSD+uH3D1LsOTbbANhevFt4Dq7/8gH
RKZ/MlQob3IUZ631l0ezSMRZFvXi0IxI0p27BCQ7gROAJOmGLhk3E8QI5qokmztv
drq9702uMZq5045Wezje4nIZ+qcNf740W5nj/Sftbls+8fg69G1aPCsbQNYJVFpx
j83A//u9d+SAdzKd9yIDm3+8a413dloPfWY89doeNIoEy4czjQ13hBnguzTD0jis
h5AO3SNCjVKta5xi1L/M241Ihx3T3Wa+xiHKyjyRJ/8Xu6gZ7ygQX8JYYJIiSu+A
Cth+e4vTQ14N83rlII57hmWSuJ/onWTMlCaZ/zQx4qgWAZ90VOsY0EBa2gjCHQsn
W3LxzIDcAs2R9UR2HJkEkLL+FWZDrVtpNZ5jb2pCS3d49io4gg06C05GkUnrTzxc
S99k969UHnrxdX0AB9fNn3Cy6WhjNRKOsxvCEO7YU85/0hKID9VIieJvT8tUr64M
K815PMDn2LocQu5ufuJbY1q7vS6ghtwH0odhau8OZNp92tFmoYvoE/pLKlGj1gNW
TJ1oi58SAc87DdBR2wxqsBYxfnLCTDnl9gMeTlKBS7ElhCUUCRcDIfsHdO7bz07j
UNy8B1Q+NR5aJgYwiUOcSmdJYuo09BkpcWBxJLQhyQ5hYgBp6/M69tmpsK+ay/6N
LlvppJcIrNSOhKoiaoYml1kdQqqXxiZcyxCaX/xPupUALO6ktqxvNwHU2xZPxTGe
`protect END_PROTECTED
