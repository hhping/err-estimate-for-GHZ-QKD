`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ELtBkNggvVG2iDR2HekejzIrXPhSDS+PDRehkawZ4my7X/Vjk1YSc4rWeefNiH8i
pILnA63CAcspnYtLeVuYVRYADLQl9waXwFNHVx1vPHrSIh7/R0eeo9UsmQzTv+t8
0fMuAg6stSa4wptFLvsxnJx9ryyCjlmTu3J6daWWwEAHCOZIXp6IhfKhcvUsvvgx
LE8QkuMCsalMXwUqeSP1l0j5md3IQMRBxR+lb4SyBTm0T9Tct0+5yedlDy0wYfaZ
YmJAsy0c8Dw94fQID/DxbVqgmef81Q1nMVr/JxUlBmXM/+Kmhn6GbeXYH5AsG8h1
YegEyuTqL09OSoUXloW61CP1iRne6Pnvefj7tHgFXFfXtggr0pkD+AmTEaSzFcAd
0nOTHJCzM9tlf28lDfkE3Kc1NRQQWcjDih7HWbcUK0o6DHOfHGmyEzpoKOjN9XOl
8RIuBFGAbq86yA6h4gr7w5qFykMchAZ/UIng07l5KqTQ+yqGSafUf7rh6LbnyCid
PYT5GHxSO9uRO+iDS2glQiQZfuN2FrXHLvoMy2uaKsYasuR5xVNqwB1ub5OTvqgg
eBdTXhIXa9s4uTxtcjXshZmzdIY2R7rtOucD+yAQ92ekDqYCQy2yaJB+6m3kQofq
NYr+miy0FpDYe7vFjFAp4qbVuXs9VfMY0UQL3HkJkTfJm/ADUIN2vPdfR4zyjeqX
z0O9IxTTWE1ApwOUGUSYkkPPur/h7MY1cLhueOWpBx2W4Soi2Ow71v+kRCxTeE4L
7FQ6/Av5WyttYck3c48XmwzYo/c1LsL8yrSH8Atwn9LXPp+xlejebQ3tPYpAMaLA
O4i9xDeJw1V6UzkAkor1eyT5JaSzWCtNnBimogAD41lD8CBVzkRTExtpPJx9dYGz
n7qtvP7dc/sEWhd4DA2D0A/64sys4O+LocahZNsX7LDXV+8LEhQtPNgLprD7VDoc
+7xuZoIEGGkpgxdokUy0vEgOV9/gOtlYMULn83DIy4uDAFvwzJLcaSGST6W9ICae
kRnTv6UHCE073z3mU0IdhTYhF9fsbfE48+9pvNIbJ2qdrk82Y1oNb/u6CAAXshIP
X6Gt+tf8bPKYvhg1PjuIDLJu3+U6Ofz+PZdZ6yKqx+Ad5+cDfrboQKRwKDlgsgAY
CyAjePo1z2/7aP3QVI3k8XQ3uEeE5ThEl2zaOaeNuTfyQWfClqRD79/kB5Qkl8Da
vfT0a2ZwqL8OywnyagkHD0kFH2cN52Pi564AIj6LRFxqmVUACvovtWpFxAVqHk8V
OPZTObh/NgtlwLYxL3tUdITIWMs2trlUJENJvMMlfO5VThAM2MYAHnlEdzc3skZh
zuRPay9p2mCZ7GJsQ/uuF8x9bUIeD1eaPmT63RwcIklAZoXDkmz1kZpiPh6KWVQ7
ErZ2roOEKtYVLE5ACdkXd6H0ODfZmwTDSbeB1aBqToIzEVfGxHTzn1fKaMv8Lkbt
6zED38BvHjZObhZ+DwIpPfHwr5bBi0W2uvsMJhr97fsbvrzomSV3G8v5fBlnP0rQ
u9TLPGW7vwiivB9Iw0ulff27XxcP+RMoeYm6+lOyhGMoWJLzeZka88Zp/Qz7VH5R
pf19iQrXmvM+JH7OcWrfVpQNm+eQmfQS4CdrvZ+OkjWHKYZKCtLEfb17Kug8r5ZT
JU4Fbd4tpeqCIIrUh1AHNph7clJI59zVqR2W6MZk/EU5KV1c04zqe5oE5CPg6GMB
u+Sl1YEsA7B2WbIKDY55Iywh3JTT1eJKfslhu+rSbzH3RFeQK9pcTEP5N1QTRXXk
dFHJmPmEBg+vz5mtMoxFynSMD5zcineOrelxY6vX94WlXyeZMfxLX/dP7ZIBRGFB
PTCvBiPZEKMq/D+WQZW7tUiN3ZoowguyUoJXM+d54CuvnWo3ua5nhb002MSTlnEG
vtBnr3Ali4GXQioTS9eLdUp7LVR7IilrRd5v4j5gMvpXmYWB0ebOP2SoCBUxnpP6
1FGhoy2iY+NIT9DjSIMPHt3X0lgHF4y7Mi8B/JvZVhPAxZe9BDK0Hmxi4YcZOFcK
Ou7WsHN5wWYPOy3zqSdpfEmMNsIT7CaklyimHjGhZgizurxouLMKVCTqKsU66LZ/
/CdcRyOvZg+eg1dKYNNp1mVmuSyo8/MgduCealyaxwomYj9AZ/a3agVywhF69NX1
NNMI6hYYVWjwXlMufyBrNI6VTQGEZ+9FdaXDP800mXQg1S6S2WN114HvQPl/MJPq
DaQmQMqFPEK6NlccOX3Yqr78jFYVpnPkfJqq9UH2CgnoRyrWtCPoOyBL/NydWFct
jSWmZJGG12UpgZ/kECXierRWfKjlRfU937zY65dJCiprNJHfDorz7JN05TJj9dES
/2SQvaJHfY4TGLvEdwgGn7hVIaXrM17p8ZB2PN6b3cUix2ipBep/AXo2JpQRdxYu
yrt57O+KBFAgvrJyyrB9bJl1oik1QTz5BUsJgZU8zWUZijqneeHsreBm/fmQTOo2
MaJjJ247ba7UGp+3X2Z7CdbF9G3ZZHnA0Iu6FOHlz2VaF7jxIBIIMGYvO051ETFZ
SqS1mvVkAz2M2zEeEFfElGcq2IaHGYxTj737zvzERQysh7hk+924Qyiav0FQ5fff
Lym7q1NQmuHGxr4Hh9Idg3OggsxpXkNKrRVZlujTMq7wB5VvGunP1LXF+7sU07lJ
6gFQzAm5AZJkRV5VfpkBDRprHDbkCA1DMthtEGPGnboHEjZXwnn3XQewVRzeMOun
InjA1vd2ZkIpnREQExWv81vc3wVuc/taBI/4WZ1Ri/MtfKnao5S119SeP3acRKzl
5SYXtHFs3OBdxhDVkFc4A8L1y8bagvrJu62obBu6I93MDRSf/CVsTvJXt1pxdC95
uAQKyALqfI6WNGMukXJ5i4AzmsRqKxGNBQVzNrLqHdN8jHxgTZ1l4b56NFdRK+71
cxl09/OlDs13nOB1WaLEcUKS+JANPQMVr5W9VhNvwfcW8blYB0kaGyTybpRd4BmE
UJl2XzZ+O5/bkHIfZKvYNb5smUr7gzbzND9ncYVfEzT7VKscLc+CM3M8OVQ70gn6
GDE0zAgVJIZKKNLgNjW1GN8mQQnMhCIC9L3HbS0SNbSG6UKpxitsumXCVXcvJPhR
SIi0NS2xbZ9912yCo484JegzPNYmBYtFHR6ggFw2FCEPGcQKqOk9ZDSqkrSCK0wZ
1h7/wSAytmHOz4nYOl75NV3kVgzdpqg1xDldnLo03oavmyJd30OkNLd/YyoX9Wtw
lC5G5s1NU8W73qclqvavlRQhTmb1EZ78BzTsw4qwjY9x4NK81wzfwcfn8LeKvbYh
UODMJQ+JKsDWjjZp7FTRO2hfNUX1gyUiy6M3uTEldNVfBJ0a4rKAhX0xTBxNr1P+
scUpOY2irUiEL1YtiG8NSVeqDi0QTENh7FZ+JRVZD4ccjpEdS++vANK/kUgWnG3x
0IGEXSgPB8KC9vQNBWgS5J9mWDA/oXYfuJ2i3O7X6u/qKwrBHB3pIaKoP9E7kK+p
UywPceY1mKcmjIMlTSqWQ9wqYgDbqEpV+GPyL0LnO3QS7jX+zR0eI3Jxp2KZtCSp
+yLSyWbGxfr3o2yG4ImTAjMyskGNfkmphAk9TgRVFuOV4FzRiqin8rl/aLvzc07B
v9YgnPYdqFGvUuwPmcLwt3r/xRgXLNCaAReAaEvHJ2eapCleeV44qtBonN8eYXZw
r0SUdKk8yI2qgyD2CShV+Ykv2Pd16kruw2DbZPtRGwUDcbBb9R/mSxjmC92cZhab
sfDeRF5F2Dn3AVEH1TKvRc40DbZzUMu2aruVlG6jMNzS5h46fa9mEF4auzvnwE55
0YD8uUROtp3xDg2E/xDsAKL7UI7+Al2YA2sZImyL+yOfgpdZUFDDdwSNwTEa3GXs
JduIrtf0FrhIq4p5drBmFKGHnRYQZIk3Io64trzpoz82ONwXi0z+8bZ1PkUqrIPv
C6BJddnp7QSTDtCt13jOjhzoaxwvvnP3A46L2sKkrwZQD7KXtl25/dqtp9iol8Nf
d111BSx7l7evxXSsR1NKNZq8sYrDkpWmuEgAWBXHdDfanMc/SiTXSEEcrzd/W2Lw
pIqKO5d6eRDG5Vi9Khh5FzVRqc8aNPRenkTjhSREKwZZ4stW/2NqkY9Y08hFUD29
8NxV1b5E0faRhupxIpojCcnS/2Zj6lhB+dyFY4fQMyQn/7uI71DjuTtIs269r1LV
ACzwIT+ou0tt8UvADrbXr/XJajuhuYebuVJhTZXE1lar72Ltt9UzJxIE4ph6oyoW
larBC+Xsu5HhDy5NOHPWoa91IaZ4wdCYftXQYuVGs1moklmYzjdaQEOOvJgLjJlQ
AeceiH6tWiEPx4E8zDUiBAVf11wB9L1wJioE7AIU5aePMaTzhSSVAfLOh1igMioG
UYR/5OjL1bBd43t5gPmkjEeuwL7IaPW7fsZmc3jXNwcHstBCb/AsyK5dDksSIqUu
I3uKub3YJahDo6auxpelwGdcnU6v96p7IWFCAMRrGnP5uktXKLSIfZIIir3ulsDw
oFNbaGmQ135F0pdvj2QwjVgpKSCTPVAG2Lor1I46GcS+eWT8slGbqwGUdQsF7hYc
1cNic/tHqdWYN7d0NV91tk3FWxqNEQFbcKe6ezxP67n77y60zQZ7U5XiVPwv+ad8
y53zkOBP+h+JvE9j9N1dbzy3eGs4Ae8p0f4P1kVXx8Kxd43OZKGPgfrV7ks8cRis
pW0H5rg6CTnfmtG7r8qtZzRyqZNa3QneBWy49GZ1Ieyb4fbpDEEM1KYECWOc6njF
HU1HPDdFD7Z/PKCO4og01hTajgGl0bPR36GmZNy+gTpWeGbIVOp+uE25KhCA5Rkb
oSC86vvudKvvlbgNLBueOdePM56J509i7J8E5Soh7ej0rDc5midZrZeDJPr0lPM3
yRxqXh2YzUnmQskb2GdvYyQCePGO5SZbO584jQPFTVktyt24YqjwsEYjc7gyJZHN
kIIgMv2UThLvJLarOQnttpexgbLyEXgBdIYHtREC2IiT4nKIaXMy3mmDAXcwd2DT
1Fh/VfqOhOeNX+6U3IYbJROsWat2njxYeV0RPbLR1miviQh/mFkfL1w1MdLHfhuO
5V8MCvBrfeVOHNoKSBR96OQ68uHMuGL7zpwVd2r3mDziGQLq6uVQTt7uIl3lKEhX
rnLuW7c7zcLBB/VpuBDzwjRfIaJT2k0bX/VjvEeWrO4LQX5H/iVumeXBX3ixRX49
NI2B2Ty+n2BTIB5fsfUmNrGCKnHeFmcgObTdR60VE/TaOocnuclWCObTJz0sso9G
+ofWMdkR6WJOY/ZdBAQA7WEHo0pZIOP/fD3KwbGAREfpYsZtA14XBeeAoX/n3u3v
eTKg0QdBfL91RptJlxnCx6F4ArhNUWJ3pqA5tGmbCmoR9O2Kkv5hou4QCxO3mdMZ
7vEdRE8ImkcVWNJTNLOKX2Ow3jLFtOCkRsub8fQKe0hxwPjYRpu9P7tGnd3xBXgv
gpxetkHgIK8ceZ4nuLMKKduqY/HrtmeL6zNGfWXUkaNMTl5g7DS8+wg2yP/d2dzS
N5UOfLHjoX+ppdkn5Lov5yjXaiJKMVzFjKlcZg6Le21jUZg6QuKImHk74z5L1Yno
tmssfQm6tTO5No7oMXfGQerYNFhM+z1227omOTxAJiNiSFRAO253F6YJPMbnazjY
G6pw+nQoDSFtpj9sv5l8CQUL9le9KSWcZkBEpzrGFmcr/Y1ThhQ3QWIgUTV+PWNk
4zS91jPeDPlDWOufoDOHH+8nIsPwTXozrVcMtOINWGugkCMqlD62uOj5Mi1LSyoj
frFpBR9svB/SQE9QirQp7Ok2c9y3M618Js5srZ1jMs9LenkCxfQ0CDlxSMJH6mnP
a5c2Q4xpVrlJaC+7FJEdK7go98L/+vUO53+F8VO2IhWGikNGZz6TNcihZkd6AtNC
21wnArztI3NgLK3geF3co+YUHHRq5zPe2eeobiQL7Zo45b97/3ctD//7Zsd/54KX
mrp17sWsXV147urK9XIX5KZvt1UPlGP5ctvig0DaQv8Qt9rRGRUD7i6c1Bm5+Rn8
2htdNcC/1DJUNaFYL70GmGt++DJ9j6Lp2IonxKYJw21+cbUrLqxpes1ZBUGypm5G
u22itw75+Y147RcOpI2P8F8jT8NrCsLSUggeOsMrJYT/o0045yTQqnT9wqP6x5kI
sgJa/UiYcGccZqTaGp47scyeWj4SUTDarOp1yus2/yC7Vp7WExFV5oIUgSZRWTGh
T+36EmiQBcYC1ZVFjBp3317A7UlhCvnbEqdCsZj/rM+2AxKo9mz6VphEe14/3DFi
hL7Un8se2Ehvpff93m8iarhZ+JwYSgk9/BPn8S6xO/0rNwkDsafEWluT1D45bCcu
lZMr65Qa5elxFs0tDhj3VVfbjLvoyURZqkgrRwmgywZ/IuVapgywbcJs9B70wmy/
xwEAudAGR5WDr4jkQx8A8UP3WaNU+8BNvbjituV1ht5ZWq0H8KlT8MXZ+78Hwp6+
Nu01rJ+KXif6rMjBbTde7/zBJ7RgTx1Mv34Y3ZQnPNohRij60K/HwFdY31mCuTDh
dQDmwEjcCpjNuVQkRz0coP9YvWsdRl/cJsZAAlW7/Ka/O+GYLZv7tco5gS2iIu12
apsNZ0mcTTAM0G4yyA9D0owhuD5WLuo30Z4Stu7qMRs9DdI6cTorR++JO6KvzB8L
YaSRyzQwEE9miFeLxq9blGz3TWiw5bW83wjTENdZH/5vycZHs7sFfD9eSC8ws9dn
E6TtnIYsdP/KBTcEMxfCtSmZLa28mTVHpORNFHtPNT0e2j7TOWrGDXbRPVWDEj0q
jAyToGmz0vT4UpfWrf9bezcveodxY3MBQUmz+E2pcp92dE+7hL/sF1Hvu/TegPCq
wlkzGoxbfGlHFPjuFm1A+ccPUvR2FNJQzeLKoC76HhkrBkDBsUJdlnYQh/d3TdI4
ZHDCXJI3stTRjDqpu84oTm19HkgklgA1L6xQsw3Cs6HttRy87gHxbt0cGFboLWTs
I8xfRAKjstUscEzQRP9oN/iKWW2PGDJouRfc6S3Ov+PEpoCcATvZ7aEYOsIDnWFC
lMJJFW0mfxwk8ubaMN0/tqQfgMfnW1Deq7YIfDlBH4aKIC1X4tqrM/8h/3D46OyC
yywZXlzSgvu+6qj43IxnfmEBXGu0jh/+eLGXKWIw84EzHLoXMeNn5V3j1tz4vwnr
Gk3IT338kwXLTg3x4Ug3/OPoGOa/UvqMkeyg5s9iiTYNfZv13prW5aBv5P+8EhEQ
K1uOajmV5phBZMuVb3sD5gREqCIXk4jSjvthnTXU9Vcy6R0qOUii2B4x31EhMXJJ
yHXkDCOs8qyRVLkC7g2w9iJW3/ucxIDd2GhZyj3rzl4cDP06qA+QOTabQazQCzZ7
rqm1ooTMLMtaYH48sgpREeGQgoUvsQ9Zl2fVRt97N3T+IV/vE04XvQ5izQa5z0dk
OyavL2pcffNXdO9PR0ha2dgIiUCOQPq69aHG1Ah/1HickpQmvK02fT159tNaxUHT
D/AWghAPydLcFZh2bFU079pKLE1Td7WXoD+bVDfM5rksHFWxWYwIJ/bAauNCPqJx
KDxrsyK92M8IabI7yoRDCZ9aJkKzAvfaBmygX0VMgt25kWVdIucHuwHBHz8BfDgz
PP85BqS7skO01MqJwpvaBeXiOPt02fu7XR+3Z3At9aiNuaWU1vbCEvyfoMP4WnbR
3+l0PI2Go8lQ3cecLzSpBR4tSI7jzBfx6oMFIpA2Cv47ABTd1fgvwQjht+B1uhCf
iTi1+w3r60y9qG0o0SIbm34t55G6NeNlcuZa8XWCHllcoRJ2LizZWS46cBSg/ZZD
ea+goarFGwzF3UACj8MxuZejdz/qxq1xSHz6tUvMTAyOP8QC80OHv7Dd3UFAl+In
djam9HHKAgK8Dr+JnW8jCxWXHt3Xet/hJv4Bxwc4ul0lt+ugO0FZO4rOVJoNpcfk
vk4bo8RHCN1f18+b6quUKJUkZzjpDDHeckkhog4wCUK/9/8zjZRF7ezsUE5xBWvo
j2nHO4aGCKdLPGvOYyZTV34J76tCytSZTbKnWT3MV6/VbNvmN4/TuDJTGjrnHHuo
iVkKxv9ExXM81Wjz1kv3Jr90QMOV/YDe29ZjUxFSvDP3vqnC/l2Xp7sS/ZB8nZZ2
iFYHY0VaenHm1OVPymhKm+grqU86sYsb8AULKdutTl8oIZz7tUv+tXNu4pIMV0VN
oaEnGWbMkwBlAOGEaWAQV9phFACEiuBVY3SLhzcTY1JQXXcpnJoWys5dszfc+BaB
J5MR2pa6UEZb7cUedTL6tR8m2ClhovOgySfKjsawxPrhiv0rd5m1VGcJxy5Bz3jZ
Y+nyDhfzhgpo80CRnsLexSZNIM9xkKmTmhYgAz+WEr57AtoSPWYxo4nDEEtBh2Vd
D9IBKnA/mdOW8FvFG6xOgT4dVlQzOOdzTet/jgucFOUTIZO5KHfoN0NwGN4LpLvl
5qotLKza4eExkukvm+/Yl/nArc1m6X6WtYPtLrHklf8hsJB93V/NQMBaINqobPhe
dQo0KLg0NGe1esP/vwyWivBlkmMfPMRNESBTnIrEsbYguTAMWnwb17z85t2i75zb
4fZH1sP1hL0mMTRqLL9HY2CB0RS5ukpBHYVQa0Dps2y2lshmhCE2Fdb3GhE7buyK
P8JChiF1/0vsQ6qaYmvCYajj8qrvH8eObNSEDwzLfLCB8CSAFhHAGO2becmSiL6V
6azXURNAarpleCHypBLzALK68YCit7WaEUZUwr84pg8jyJSmBWX5RpKWYbfzBzwC
pu336Nvvtd21lC0xBrYhMmCBbbQ+WK94Z8uRLMK6wNC/H1XPAFtGpAnixHYpGkpf
NqNO6BNVpJcXPu+HDsQPqcirDp1KQ0zXDNkocEzZf7xcv/tpQus2f/KDiAPGN5rL
Zc7uCT4OemqKsAKlzn7hHZnQYWWkp6muVt1S8TWLyV5M3azXFRB3UFP+DbH2NoQo
pEgbYzPh8OQX3npBqG+Hi2DNYyeTgBPbIYQ/qLoir5Abp+Gi6twZcyWbzbJOMbw1
Uo3YTJUbYQ46JElgPuDCkQNXoYyJOhythNh/UR8wn6nmJhEB8KYJr+KzvpN8xALG
TgkVoBAZDKIqR/7fpPoERjxqsk3I/thNA8aAMPrUMxmlK8xm6jtDxXUIjFomnC1D
6mRUOXQOm8/idCUJXBVBzO6RUQt9L2Wze0A9AktZNqlifvXA1dVrkQIuoG8QD0Cv
+G6yQyZzHLUs/60ytyanHORtCm26cinSjJaRhShlet5r8hHsRzCV/ESq8HMp58zT
NAw1bN56Q6BSCQ0sA9KLs6tbs+gsTvpixfx9eJyzEa/IXuf5IkBKmUsqKvtZGA9o
Ti/2RfyBf7LuOQ0s2bWhS1fkvs3XGtS7oFupLpe//oGO2zCWmb3Pj3SmkjNR6xAU
qvhu69bnzCmSKWBmKxKMQNe/ZjQcmdOOh37ofwwcZ3YLxqebFFsD+9zaICiE8yde
bWvl+hbf+H51FjC2wj2UP6nq6ftGqqQDQxM8eniFLuaqbcTkAbzF8v6bJdspmkFV
slwWpwKjHq1yiso+dJhFEjLh8k4psH7oAdiEhzrIlGdm49VqiuCdk0whOFBQCiRv
zpWs5ZGU0fcNxq7PNYOVUFFmzZP/vtcfA7O6VANNgpGhhxg93RlLOiqbbqP9xHTp
825lNRAZJ+16ui5P623lxfde2I160frbPKTvCPCku3aak69SOiZ6eJNJWKQGy9A7
hg5P35XI3g1eMGDsY9apv3KI+fR3m8moJMsaHBFBaLg0MJgLWxf2nft9QqXxqtym
S6rpf+KdMkElnDJPoC4qBXxmVFSihaw45+Tsz0/vvaMEH3x9E2zmIB/hQCoFal3J
IZywiQciq8wtmytM/cn1V4t+FiSmzp0qK7OughNlV7WXShCvlzwxxVIE9dqp0XJV
xkUjkJtvLmeeIMZPmejU+ADhKYd8EiZ+WEls+A4LPGeoCCR+wrJ7QiT/McwFkmpH
zW6gVaRwTEi9KInDfvqK5d1fx0jw6IMO0CJJbH6m5j8Tdkzr71afsbTWJr4Io0a9
TAqXr84lPU6JH2WW7p+0EujRWhYrd47z7ECgMAEd5fBeBI/DEaFTpnN6ZU7i7fAN
7AlAWUYk2Ts1xjiOAKCUseuWjj/K95MUuwAZy/p6iogDIjSh6nV8w/zDBihzYTKd
KCxvTrkwMnvn/NhZUqBGeUoi7sSdS4/6nHFLU/zrXW6TQ3BVmADROwNeWOkL3Be3
d11KEZUND4wFsCN3iOYx3jpEsep+J19g4vKVHyFTPkqwOFzErBfO6K+2WIE0tLRT
YAY/5BzWVtFcX/lTlgHgQaq1Juxidbolo442DPFuuXCt/ueu1Vri/wyK+7JrOLUB
4ooBIngU1frakFzn5GWw5GEw7eKHqcYWRvRXYSzucdr9fBas0BlWY9VuzJXyGFz5
Z4Jgycfy/pbOBVf5C3lQY/+aB9axSgIy7ITUB3BX4e/3y0vLgBuCTNvy/xpBHBBc
ElIpanZJHW3LRK7HqZLyUi2AHaiS0WphRgJtf0ofkB7oHxfJ8QkA7qibR8/NUWeK
nGfG3+rdXcymPD0sR5tzadil+tKRmVcoDstXCWVgfSbqCSE1p9bKIL5jnykRkfnP
TAXn9rGI7LKz44Fr9uCfijixD5K04IU+sQ32nMPSH3J8T3MIQROAU8Di57g1gP/Q
bHYvWS1BUwzFQIc7sFJPPRYM9DGWaUzzeGzwbG341dT6CwP0FwRMfT9HiPEZN+qC
dnxF8i96puBWXJ+3gx9ZMsug2tk6jIwysvtoR7XBmiST3KwEFBohoKSy15UrBCGb
UlTdB/xI6vekoneSN/Eu7Kr2i/u+Ilfb9FY+mtmHqezll8AyL8+Wk0dCxST3n4l2
1fj9P32z8sEAZTkEC0jz84OPqxDTbvQmgnqfJTOtJUcgM4JD2BjLFNgdGKMGncWX
JmJ9X5OCzYoYAdf5xTSQT8NiqXCVgHQ1mjONC/QLMa9C6ajy3rvt2ht+EkAbFKRZ
7dy6eisLToaYxWU7ZLAV+zvzjKyseNS1R8IlhyRchhOmoyoIX/vqUdNmw1ghBYua
eqUpL1ANJU0Vv5LAA9HD2jKdACAsVezpFLhzJQQfzs1/UZ6nRuMjYa6+SkZnj1oq
Vx8lxqITAQFvU8G1mdr/Z4Y1AoCMlFMr1KOQEsMF0f47+Eyc1nQ/yOtf6X1/973j
hzskRm4aLhiEscq81FzWeh9vtoC16HzGsh2fgYLheyXEa4K9Uzl3agOY8pcQUsS5
3vm5nFFdh0nOX6bi6ij1LaTVZ5QYKI+F/uPqugg+FR0U8A8YdsjKscI2/oW9Spyc
vDP5pX8eDcCkkgD9iPeAd2lzOXjLfmsBmg/GVFiSVRvdOIckXYnWh8VuDd0BHi3h
0WUXEM3jO4G6DzfXNv+b2x2joF5AAIXrsmGDH+F4lMX6KaHzpRc4MkyX70wbAjVK
jl5zGTVvL5e7qEWjtyXgYBkANqdY+qb3rchUgvYJj/b/ncsbjQeqKcWAg7Qv+2V6
nox1/MWdxPYhPutbo3tOUcr0Z3L4oYIcGq0JMCwcA3M5dvsg/ktQZ8uulC8ueu6c
FMx3xXHiBrTUyC081vTtLw0nB/DFAflgw+FBKgUvPHotnuCHLDncGq6jMknjVijT
AftpQnUbFTvdOUJ4qyeAC0C7xALbd9Jj++SHqEOUiegigPBMavhPF+pRUbK6Q5Tw
3+h4HLlZTGug7mfaanRLULYWaLQk+2ls6qlAnYhyAMjg7XCHBHQfZ0U8hQTGLmKh
qa45+eDywi77r3V+kkDytrFSKdvSqBkQUIJU0UhZkwZJ14TGsXsUeXe/eQUx9T9M
gcmuwlpk7Uml3xBDkapmdzo+ioGT3QELANRwdQpOcYrll9kBh26naw7ljhrKHSAQ
hXS/aLaRP03ri8w92Fe0K73A+VN3QLTe4rUSr5D5p8AXHkKhrZE/34qUHHjFvTo7
/VDoIej1hHHqjJFjT7ZDb/SeXipHm5tRqNxQOAkt5Ho0NRxvJGftjGPkLuLAyIms
4hCf24rhxSPTaNNAqai5T9CQc61ijZ/jI+vdQVdjwYFD20l0OvHpgYQgq75QgQBn
txFpAA0njr9/U0dTS/lLzmjIb0L+XssNU6KoNtPHbclY9NhBj6r5J3PcbJLQazbM
rqkB/H6Pq6omgYNfC5GyjLzpcIISHBvADhMG55K6NbJOfsxHJJWjE0P8ES5DMRcK
lgbZqETBFO2iR1vm/xL+EEtLZ3MCrCZOI5uDIV1LpCdILGqNe3yW0EjgXhDtXcDm
7SZOSr7W2Hq+vM49lBsPXAnEU9Kwun/3ZNCDIgvkvMM2uxNVlqZ99gW5GSNMkTzR
/6OxbaJRD7GYOKI+MLxPJ83NOpG2Up/wfyOiz9m2Mo6zduUQp4/W4x5ppGov9C8K
ifjIrX8x92WqoOhVnInLxzUejJzEfSx22wC5AE7GqxNxbcfQDNnIE/JZE1LgNnbC
6j/P+PoRED2DkymkUj8g8qs4qe76v+urwaoJ806hPlGel+cTAwAUIH2bz1vE2Hav
ZWEAsyvQBmNnh0Aj6FIthtNFDHSGJfBWwU6V9LzdWVQ6YJDVcLIiYAO+ZAW8d5p2
ZMbZxWRfm7zHKc24clMiQW0tJMGF9Rr7ESuSSrqcnv9JRv4wr/erQDLtTGOCr35r
rsUvBbgvO7uSYxDlcBlGBZMhax/OIkE7sFZHTxfG7Q8HIpx/XpfBgjli0xq02Yj3
nDGFO2k8q2r/yXEiYuiJ0oJcNd5PrIZS/H6kemRFmvLdsgBOaaZaDjU7msJpLXrm
itG08KEDTbS3U9E6+NLFPF/R/pkzybgth8iMC6SS0UeLhg8y2RjPq0vNqBH2LBuP
3nCTrykkW5K+pm+/GThg6vQFDu553C675PXNRWVUOtQBMzIdi2SklH//PX1AoZhK
u9IWIe/dplImDFyNXnag8QIJ3UE8tDPZOqkuAHn6piMBMYNRFACF8Ag4mL3wKk7V
f3uEULk96F4ZaAwJmmSxfi/+oYs9MiC+GKz1UEyyVnDp5dUMceGy1cncXzyhtUnM
lLFEHGa7yr+v98iw/4kYmiPVIzQ624w9iRdrVC/wwzmqnWeW3gpBIt5YmOj5E1rz
LRlBFIzhHXSnyiRxsPnOhjxuOzzFRFfhV5/PwY6f0Ic+Ta296lEkk4E4G+NEDPE0
vInfxf1a55aPSfXsFKk3fH7SfJ9xMDjpWD5fGHH3x0V/SMjgzLcP9W+e6IUaJfjC
T+5YVCVpeAgVH7P3Y4G1kMQhdYR8AvT6E3TQ1SX77Jzf1esUXDpCRvtRwbV4UweX
Vl/bkzQEw9+4EH9uisCkQM7SUskmPXyGRW4TfseJU6DHkMhnJHInIhfzfc35BJlo
1ypY3RqlObavIpnK9uO3JNFL3d/qvfrWoDmP8HhaVBKLbFb6Vc8EwGaHeI09mvVU
vt5ZPO/K9FPJv2bQPuaTnBU3XNUmNYWtmP+c/kwGwZ8rpqzV1oKnB7s4lRPDE0f8
8uOHNhTh+tR3QzyabYh55qWx1vbj1dNCxINGc9K9ZsTXCArV4QaramKOMU6mZtLR
tMYUfj3HJJ1pajbvMkQkGZ3jeOQUbw2rXDG9veM5qQpCt0O1hZ2VlsJeU/IkAyq3
XHPUaLbc15MZjNwP/2yH9Cg1RiF12jZtJjoNFgc7PzzYdwQtBrlgBqg3sOmHFk9N
RWCcWw5thN/KAcc620g+2ELGITO5PqeNq59akNJ/Xr7ylHn+pKjK1hbzJZTkvjuu
ZNc6SF21l05Pg2sgygy4hM0qH7qIn6DPyzTvAJsS4GTVbdD+Dfjd29ischLPg8Nz
QnnPsz/O0W14RqmqZdEbxfrc17qX21FABEffTSHrjIGBBDfggR7Buts62R4SCvaH
l5h7t9e7AKHk8pPVcCue+2kXBkNvXkaPaZ1V9etnzZCrxEpVJpBKLlu+OuZ1qiwI
0hBLvcXvd8t5BuT0A5wwQMzqKisCaTnAqGgFGhSi/lDlgW1XHeCMDy+bLIzi9+Uy
PWIBtrD1MU2PXUbJnq2GFspM9AisGdIxThsOykF1vBX4rbsG2mPsdXl+L/CkdKZC
0upe+BMuzsBujRs74y05f/kD5QN6YAc7AlOUXzeXfXjb0BpGb7Q4mr2SmwsfRifD
VsH+YxeogBS/PAZeXffbuCV+8azjORopfYEjG1qbQAYm+g872gS9EBwTsgm/+wC3
W/6/EWi7xPKwWXqa79vvJCkIl7uqXFKopdeIBDDObbioYuK3PwUtA2gKvRgMhiF+
0aeMzodNDbRtdMNq5lMsZUzBkyoiwaRocLMmuAVd4g1irDbQ3jOpezdereZM0O8O
/2gud+5D3cVB97OeYiLajVozX0g0ErZcMtlskc+mfciGyyqbqDb8N40tmT04c3Ou
T8wzh7j4JBySt2Y7n27Rr9S3bWuJOK+6NHeKaw9JsImIEdGq9mvP+1h8LPWvpHWC
raJGwuxoN/x8byS3uiIzFEvIAb2f0fR96pniL/eZLpKJQiZoapzzif432RDRkgmG
hyz1JVT5qfxXqMTew1jtd35GBOopHUXicjg77VSRfqApkU0oG/1pKwpjAAw8oXUM
PNtZx8FxyDhdodN5+SVSmCzHGVdKkJiRipPjS6YdqIAZG4PKOjB07xZC6E8aSGa5
kUBbw812y2o4KrvFvCnnWR06qb0lXKob6DE6r64I+f1gnOj4pU9vxpB8eSKt/NqM
ujuHhqlKr+sRVtkqdWjlqv6VB3M3VOwLwg9t+9dIeMkrgna9srkTbx94Rt9kfWcA
QHcoBHoaiAM9vQdl7Jtk5V7f1/ZbqpRE5HVWiqkaTlUaS+UBPZOe5gFtU35G6brk
3SNOzGItc3VO1Gb7UU3QPfogrX9Qm/MmpBSRbfhRWMiAi7hQQ+TE6kswzama4DdS
d0zOVanxTG/fzuQ6t7OR+VzcNqywHyNPi9BmuLJkaMQxFTCUg2T0+ysoXQWHQwVc
bwUat56Fk7mXcxDve0hhPs98Yql2YtfzM8vgc7oh6qLUL68iIdbmOSIM6Dki9Fq3
fnYSyLMd1AyVroLWPHXILUrSvVIOqKGYjCCqrWN9q1lQhd4MnZkpT5UhPF/pbG95
OXTdDRDD97efbJkVrO/Tg5D5FatOv1bmb6CCaB+qQdl8WXzKFPLyvjubMRrvqcIr
fOTtMaRwAib+iCZf75+afOin5MaMd47k1N4EfG/WbbjuZNB41pXEfX/gQTD++1g3
k/4G6RDr8RLpBhZz7LY3H2bm1x96FLxGwPi/Jbumal52J02tiEd/u6IZVwRaj/4+
xDyGg+h3LfKHs78BMPRAGHSbBdBiB1aKDkHNefbIiFEOdMoeSEsyDvlGf/ENvb9J
QLd8isYmtEQkQuoEAfSJ6qzK9R5B85U/UujKPQhJSrTMGGtrzzwERHJwVJh2eTL4
vhXkhcApLi/t9CuT0G4KEO6i4LFVXW5CNWYXuiUhBVZi4PSYI+7QfPFzpv93u8q2
uz96tM/Z0DuXJo1meZXZVbUTcP1+KVh2G2121Af9AkVE+79276YIf+YlDN16wHGK
kD1F8zCDn+c+ghkooEaylD/Vc93VfjnZYaP/xN1+KBCeJjcGvwALDWMj4ymC/wo6
zjFOjExE8j4Jv1Snz+4Gn/k/4btMYOF2YhP4UDiAdAHtOTiwsPW8U5GAd9ox+7VC
OHjPB4K9extuSyKBWDfPOR34Bx+eshJdIfUl+Ynol0IMG0BFmLeJeE8XDQ6W6LnO
aIdIoh860bFF5EvOOTLvPJy0lDXwFtqIk2TgRcNlmTmU89Evy9lcMT/d8AmCQxe/
/c8+YeQwAfcTKXFVopV3Zg==
`protect END_PROTECTED
