`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmQkpYhaCi3++OkJePZAvRII8Z+4JoGtwOB7eqKcvfBl0bTiSdeuiElClEleElp2
RjC3jGf7p/ibF8foL2CETw7UzFx4PZbFkpSDNIuOkC9AnRCNl1J+mdSD/4XQpYQ1
9GDXsCp0XrlaSJ7uIDHIGlhmLD4vIAV2di1QS8HsVYooL1JAuWRzo4gAzb2TQ8Go
i0Vhi4/t3DhbGLCmAf7uf0ZRK9RUkbStj8C5q0gAwOyq/tyo/LquhNYydoFo7iTq
jYqVe8KGSVzGDM0xgAQYHnMyxXRbALclNZTcphqwnMkXxKKBuOEviDnMSDm6mgnz
La4JC5Hdo9XaGbfWdFZdG3yRStoK0OvFzRT3N+kZZ2t1i3yArowQ/+EYMD4P52iz
1LNBohxwcEUAB4SL8lM3O/ll6trfDsFAowqQ/oQlJe1oc4Pb99frBqAPrQD62ILj
SUoyVSc6vvdzp1bac1oW/DOGxxOZlLdsKKEhbGXTpNFMGikgxWfaF07epn77Qszf
+23TFf5g8lvYycYCSxN4wAY14JTUvBrE7o5zdKWkQS7wQMNq4o36tFXTIMKpq0Fj
tvlsnxrIIK5D3MEhwCa+sPX7qP0QlwENLTdZVwhcx1YxjNyKLeBOw9zIkKcXSirh
uZBVRR43xM9ZlTGHEx89kYulhTs4eneT1f+Dz00xh/NYEpOq7utcGLiyNcT7giQ1
rGjCZkzarBqtUJ062ItcT4wghfKVKFgT9V3eWlSgTTjJCjoKlNaPzsxYoi2UTBoO
FQla3cXSOmoeqInrXa1+JOpZw0+RSXpyihebP+Gmh/c=
`protect END_PROTECTED
