`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nix9Fqez5BcKi4VoAlN6c0NwtL2y/+Lfajilokcd1/nJmS+HA0nXnL9/mEZjL9Fp
tbJNMI/rTa+PquSgtjbb3kXWsN9I/7WdFRCh3BzZdURMBmROpISiXAy2Kxq1Tvqu
WjJXqnjxz3vt5MITAhMCL34c4Hu61CRdDxtmpPzxqk8QiDllHzptTY7P5zAJojrd
RKNPtbu1f4D/Ne+VAeACrUhgdXJbB3nTehmoGgQxFUSxZ/SImrwWwi9dyhiMgfde
CCVRZhgcUnr2cx62TOuPhPvZpDaXF32+CWLvdq2EqoabRZ4WTxiY2fLSydEYFdo8
Tq+hSJLZ0vL8q6LXgFOlxZy9WcPU9MojsRAVIxRPTlD10zaL4nlfiTwj3ZPHczJa
zfmxcHTUBfODghHAZ2A9zNzMI2HHKoau3unEF9Qkwu4VubR+iQJGZg2GtrE0M0I0
SjxbTmgWjmzPZwqJ69aWojl2i8W+AS67418h2oyyIxzuQnq+tYGOPIru3vus6fKy
VddxX5uU5TjAVQ3OegbSXw01dBwap4pakPKcrIQ+SzX2U+7fQM7aPuKN2lEfb/yf
DspFlQ5ZdlqzRsbh2z11JRaq9ZKcdlY+hYq5GX7EFrkLdncYKF5WNX3trRoOTSEk
bxyhdgvdP+drOWp4yBBGjORyjnRhDf2ZOQqm5iM6+j13Pkedk9WQQbn0BTKi4fq5
pcDUpPsXBHltJYQqTUahD1n/PjS4gsGEVYtYFS956gealYWxK2cS2D4rIxSlMMRj
0argQN6xq37VmE00n6RUlOmlegWkwQhJT5NYtd3LeJvFWBKrVd/wzHNyBWMyRLIE
wYZU1TsbVxHzPffWm9HVdW97MYI52H5s3K96d7BbXuRhylkKHCTf3QVZjDC8FVjt
HETE3fmQOcgNM3f49Q0fTe3SPw+MwKtwBJaX5XLP1z6vqmkSBzfGf1U2dFihNagT
FaPyiUKzWaKbU7mSEudhCfQkue1wbDrU9Ct1keJ/AddZvq9dRpAZEF/dRFxtJByo
Y1ShhQ4FpGcB1Y7ULcc5JqMthE1T6V6LWXpKPdI9ONfUTO/DE/kT8wxeqt6alZ8J
`protect END_PROTECTED
