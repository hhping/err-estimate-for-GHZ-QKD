`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0scWTCwc/RwKSLMXQfbzHEF8S2CzJh+CFobMo7vB3L5d7eYs3w4S794pl6XkAx4
bGaQfZTlRluP1u90WbXN0rwtenyR3hUf8sF2Wkl8MOV3jhvs8VwjL5WqrPCCo7cp
cWLhWneJINFTBNNSLarzSDNXwpoRERhvpmCNrNM/kF1oCNUtR+K0GrVesupXOSbE
T6PT2q26T5ZV3u1/vOvkjVO7gfdTbQo0eULfWmYy+gnL5JR7xuR/Vx+fb/9jSxLU
DKaZyOvcQetoZnQo9VlN8Q4W313qchE289ZM8/3ZfstPnPaM2Wl8QcPgV48JW0qD
xXzA2yi2EyUmnbwGbZpe/ciuzP0pm4+xs89pMuUxqkp78rrf8YxH1SUMcElXT1yv
Mo5o38hz3YeYYLjdD6IWzvbumpJYN/qKJg0Up8GqOGSJi3JI3OiXReG6mwf12wuw
LYJpR3LR0ElPeA2HEQVGzJTSjQ+EO5B7QfAsKDyrmmFm4vG0x/7prQiMxWC2U8er
nfNzgHM1lA3Jx/DYYiiq3LPVEHhXAHY7am2AD/uYZVbymIOC17C+COiGuvhn/7rp
y5jDVaH1uD8M+eX2SU7kyYFp1lH67Xbrumy1rSazlHCTdh56e1uxa6Sjs511GnE4
x8alCavnEZoEiYsWvM+5aUjO0zZdkzolYpBO7M83MMoFzAOR8ABB2US664KKEfKf
epxiXM8tmsJq0nwVkbLEfA==
`protect END_PROTECTED
