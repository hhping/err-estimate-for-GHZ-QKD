`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
05dAH8KzP0xZ3+tFHhpRRrYt7lvpBrgnH6UfkIU/ijP9/nHcLxS4gZtgpo4QdqxR
/ZTEIi5O/9FclMTSIr16E6VGiHUUQJ88a06rA5tuaWfp595ZDbYeBm/iGeEiBbYF
p9ZlfLyq7+t7SmiyGGLlCY9sBjA+m8vphDRX+igLWMLJCqU9nrvVWTbnUClWhY59
ZGAL4GQtdbmRTEAPSevXkU0dc5Bf2RGAhD6pxTxgL19AMmphIz/l6WwGHD5Bufc0
hcKU4jBVUi4TYUH76JUbHKCMuRSo1uHut3EDMqKwpGVJfbYzutV5bxQ0ufbJNaXT
j/yWjjqwwTi9LShRz5yRLXcaHf8ugDK/BFMdjdiQb6VNmmDwqP5+UplIyV7c7q6r
XL4u2Q3AIKafpA2X4Kb7g4uV4F0pCjYxjmZsp1yliEooGWsM5sO38bXF23HfwcDd
9uCwOtqxbRSvNXr5zBlsjxIAXAAU+6kZf+J/FvPuZqn2oVe40nd3e7a3+IR+b1TS
g2DfxFcmcplamt/fCuPuIOS0McT/BIAcuGnw6pLlhI11v1biQWeehFR+etWMUHo4
xJmrNvp92+N90CvbwkdsEsdI3qDCMFzEJsjNCEDLfSamoDPXPzn9hzOqP0cF9/ki
VyeVRGC/7+B5AlEc0uXXfBLd7J1wUWaPzDCWQFb/y02aCmgdmhAFeTp9catoIMP8
ANcY2ajRcviDGn4/nD9WQzHs1RiWjAJTNVFjYGxD7wfByAydLj9bcWTCyCiW7eXz
3mp7oyLGjqBasDxDc0JIu5vRH9xcqxwAGwRpHs7mX4n1s58u4uL7jlEw1mmzDvBQ
97e0dmwV7qDfnpV6dx/D6pNOCg55wkxG/J4p3yyN6pBK1lOQmFup4nG7nP1d2td1
a9SgJRNr0joDqRvGS9jFmBdIUl9gtN8+fgT50EdJ1flpu7KBx+tIuRJcW8s2ZYj2
NiwS6+756OKXR5s5Vq672VExAhsFNlMI30jViJjN9tX1enYlDAu4wLPb30Zdnz+f
ueCAKEkYqRF4MKxScRnGOy2yctuWUFZjM3rSSvbMTvWq4Lw8n02tEweDHazso4pm
+3rIq2Np1/xCvxc5AuZ+9Z81NSMEdskOULsEwzgAVl/Ab+XLyqSm1iPd0/k6Q+dT
Fo3/Wc0Eb3q5dCWjrKQ/askxIf8xDXCUfeYoye4EFpnUq4XU5c2cRnyb9+LHp6Bo
0Z0+dreh0RY4xrnmXJi+8wnJwkkKLOB09W7d5Cnx/kedn+spic1Aj9PtYBV7AHZB
rbPtm3J4xTNbvLhhwNymh3mo1OvwVOqXjDeretvy6zNNYqvfnsTo30do+oOHjcrc
M8gQHvneSesSt2YJMv7MVxpwLa7Is+U9b67n3zoBHVIy0Kl+VeY8mVegG1SD45mb
SjctP6XXdOELQkwTZntYLX9PpTX9mi5AONx16UOrNAARDFkARGWJJcRPdtAbRcSs
n5CSGv3C9kpTg9cguKbhFSF9IFR/A3Ydn2cpN2S1tiJbY1w1xdRmodJwC6RElLpF
eeSmAx2hicG1cXZaHyymf5txmSI4ARiVLLeIeuSVvkKqjQB8GBBhOQcO+vpbSJ+i
yF5wNdY7Nlrgru0SuIx12jwaDqi93rC9I9HFaibukDojVxRYO0JNArtqMQufE4Kl
MY/H9vIF41EelJ19empkPkPNU3OXAARrMK7Qan257t+lRWXmcrnUPwgxp0vY+rKg
yWqza8s+vGSUkenNIBKWgUnqx2vRBm4JMpGK7za2UhrsG5Ji1OlPxofMcyJCSaGs
zrEpBow+11YI2F6MKJYwi+m1w/RgP485UcX5eo5OMNsAoCwVaEKy59FVVr42qcGK
LfIbOGbWo5grJFCEW2zWg3CNN1FFJIIZepTgw3e54u+26JcZuL+p3LqdYHa+CYdW
wtbTp3DEm+jkjRtgoF8Y9OwyS13L1VVKcWOFzv1du0iV5lSPtpE3xvpZ2ZoWYbei
dcsqcClUMoBThsAxXzI5RBSlTRKCmSe1mqEztTEB3oL+VWaN74EMbBZ9tX382DwO
hKpfF5v7ZQrA+hcvbXX/lO+X/0KqAcTtySVNriHiyBDl8veZP4RsOinROO9/EPpu
0EW6CvtiBq0KjwmQH4hYElvzDHMgGTV9IMEVeZ1typkaghM9c6K7bkpGrxWlrTB9
2Vrz3R8HTF0NwpETjXad2pZTZt6EVi5A9jXDd0IRZNuG/FC7hLKNWPcihirub+dH
dzHTYGv7fEMfpkuMsVf3ecyaNCNXYp3twQ7bR/PYMQ6JUUd7ugifFcuaF+ptLlbH
hTkYXDmk7nUwBzUkmeRxOQwG5OdS2QPlLTgA/Atsnl12gzQXRo5NcbG3pevosQaQ
KgVZ/nMK09h0KgivfrOpTgB+N98JF+E5ppvooPSph/FNVv5qHPkNI3oaFU0wIaCm
626QJzqgA0F2i5Q6U/HxIaK62M1z6DTeGc54iYxq8bQF98D0pKjeWb/1yEYUHF8Z
2fOYUZzuUYGoZnvfqJ7PrreKWoanatJwOAjEmSjJvsxY4LY2JpbO5nui5AFsxbaZ
tDK6ReS6MSLSmtA8H9yAFqBsgkJTPcZzKMmpxTGyQXVRt95+am8xBAnbPZfyCCsc
eMofSdgsTYfHfQ70u9/Uu3IQgzTI7xfGEGy+5TfmjMoAShsgLOr0WBHpR1gixufi
7EUVLKIgK5y6H274iVZzxjT/DL50uza4FDUmjSxmr4xlogRO4Z2Jur6TBx7UFkn2
MQmEQzhQ3pdlYW8QdWDxd2CEhsCs1HTsJ7VvuXgwEGuCvdO9QeleqZONv9HgAwPG
6Gwjw8+3ybyy0WTaNubSv+JtyASF4a3lMM4ZwSqwZ9lUTPOiicGT2R+wVafMKuKx
gDLGKkOjMr5yc41G02BbfdLek6hE+Em7M9liaX+/9NsxfJ+WIlFLTBDzLbYdo+mW
sHTlY1F6sjM9DwNhHEYNE8w9ABhu1lvK4DCpPG/LCJwd4SRvAGclW55Ko1DuePu5
iu4sOrAFYR8EErwPrsxrYJE71MjBnRwiHYZWPdOy4yswwLA8OE/SREHeHT5UvBlY
Uy9XF2R0H4sCaPYwNLiFqj8de8XkZES87S4DCC9qLu+/tnqN1MdDXfI/jdOFZcz0
IefJYKHQRQFkoiOpDga1SITrlzRFa4mILKdFKdtpbyCcw0BWR6+PDfYnKtDxbqx7
8Hy/Xj6twOV44x3aJJc3ElrQjP7UD1FKG1QtDvJmCmv8KPEO+CUO75nxXMe5cOg/
pFiHKKVWxKyNgirY+JUstujK3gedo1cdwyzANOpOnPj/lhFxHtFBy5em2meVPGL6
P8GjxsKXNr9/fIqt1vCBoFLojBflfX7pV/L6kza88m7pUjGRBcY2zPZfxvwy6gy8
kDLe3p7piUT2ADhXzFXm1XoeVNbZZEPXbZRu872VK97Ey/qU4TXWmk4+ayee3RF8
b2zHHA0EpLxABZJO4CA33jwyoddJC8NvfTxuvmPAeO8B5lZtVUyfg219YVGVZw2A
mraYbc6eYyzyinlwttg4duTHTVlF8lFA2J7N/ebPgSoXhBRq9F1J7iaUORP+92pZ
tFQyVu3EJUGa7nlZ92lLxo8maQRCBWa2xVQPDxQvNlJb2T95M2jkmxcrJEUeEPrB
H5ooSMHeMZDO/dcxgR7pOXY5D46cmK+1pXT2RVstBHh5OnshKOgaT9Hv36LtTgxL
9/eywzIfEXYzBF0d2YGPJ8Aj+NTMTzw3Amumx+vV+OryOdajBnXhJ6/IjrvGzpbo
MWpiyaqOXT6n/15FoAWHiQVzaUeKBcyrBRcAWIoV9PX5pPCQCMnKZBTeyR1lx+rj
19diehnyg9ob+1EWkaiuQDnDQawTnTWiZP3JMLaSnINjOGMMmL1hQaSQlTzDJJXP
na/nNY1JAcEgRdKQcQvzaCUehy8m5QhTrSYtrD6QqjrX3QVJP7o7o5rJ76+tlq3t
lwOpcd8QexjGTgf2EXY102GAs4kt/LosdhCItRbyi/xWiW3EjD8Pi0bJw3NbhqNI
5+eMKln6nH+C1aKTJqGLgUN5DpoIJ0f7u3/pAQMhX+rd217z4zcuqEGOXhESrPfq
I8l+72JGuUOZ0nU2H9sM0xTmFzRvupWDn3GckYyBYnqvZhHPkEzQ5Htb6lj1LyG8
V/8LzFMdu8Au7SYbChRdVxKEcpNb6J7wVIdi6z9BT8IuQg4qmKgHdgB7XqUnr/Cl
yT8hov9DqrPT4iv4At4WKw3VywEy6bFWtiNYP3OxX46F/+CgSjEPjPVYS1IJPAy7
GiMZFspMIEy9vvwtwy7tlWvrSC7/K7DCd+RxG5uTn0HXFLJury2wz5iiwg8mwOUG
Xud6v3nddho6TEFfKONaV3A5SD68oxPdAQGHjMx1g5bsH62fPF4MYIxZ3xelRxQ3
/dzQIu8t3iHpjB4SO7Ljmkul2IsnyhJ1pDSP1V447tpAT/ZosNhon44AwUXvuFj0
IojdezrvAuIrqKmyrh+DECDk9386ZoaiEAgGEDgIeSxNbd/2P3uaV+/OMNv1JD2u
qtNdN0NEkjXFPzv2ksCPJH7FU9bzaTjn8pVsPCXgWGdyS/S6+uLLG0KjCcMwxqr+
7bL6X335PU4C8AiCVIKU1siEpxP8LzyYMWRBullQrl+ihlDmzWSwvY21kYSiQNll
ScQne//8k8dgLsrjruePiIOxquoW9U/Wfz+O8T/Rm908DCw+qGlhdeCHiIYu2RlK
zM9kZ8NUVuNSYsEOSaaEyRp2t6dc3dyx1cDcCFfFsfkAxrajgxxS8JXAtjX0Zh/J
nviVmXtH3rOirwDuL/ezwlGT5sP6I5c6Mc9JbxqRZ0D7chqhL+gGnQE6OsC9GdGO
p8bY7U2vrwrc1Lw6YQv4M4QftpRonND13APmpINu31tL6kTAeR+8XHeMUAqrCmy3
dmTG2VeMC2CxAvBLgE7hEza5kzoL7lETgt+rzVslwLHDkSKGDCC8u0dIJ/c2zscA
/+DLT0ckXsa8bhXX5liDhgpfqJ+pXYVoEaGHOujgyq7OnsJmRHiTrM31dyLqfAHm
f5UBGvxmlAm9vhSC9NkySNFxZJY8hGZ9NmeUZQqv/GG4fY68ixn9XVCUmR2Eo+FK
lTeAz0RCLXNDAP412Uy8DAlVCJY08dLQKqRsgXQNDJbIOKr0GUsA55NdKUaRRPU2
idBkU0KpQubvJgKqMJl9sgMf/Z8wOEMH/ZwWrb5MESUQSFUN1Ia7gO10guN1eoh6
OIN6bx9kz2R4cq2mgZec9U5QF/aC879c6yA9T4SVjbhjSgh5QAui5EcocQ4J+1iR
Az33gYUvAEMSxsLokosMXFQEcgoqKZWUKT/ImGTNk5PXdODVhfRbJWEYq9w07BvK
0ux9VfjW+932deSfpccRA08LHthRemh26myQxf8BUcH4UPnJzck77mn/GhYSizVz
eAd1U/Hk1oUkYuVPurdN/mKbB9U0g0Hsq2vQtgBNdHNLRmQh99gt26SLmYna04+Z
tlR5owujWJC8okUVwqsL+jsuo4Ut7my68eGtQH+OrH0k26fgpP2eGKsKYtTWA3EX
LTWDokzLbRAMFyX+mkeIJPV1RBh5xxmN1yyuE6fnRjKJV7nPnw2b4dq/iC2ekq2p
wVCZnPPMtTMeGFnxItHjQrIeGGMKhHctdk9qzfQ8+RREWyQCeTE2v49qS+3WLHl3
5a5EKy2bPeNPbU7nKy1exWIxg2llVrXnq6fR/bVNKt17vPKiw6INuAPMTlIhhJzE
Qm2fh72TTz/WX+KnIGqd1N7HZZD+Ku4o0Vm3csx6+9Pts31xazSB4ycWxQ8b70nT
t8fTw0r+fWFKWUIJ+8QyZbJeuFwdhQUsecAZr02BGZbJ2rqExffvGk2oZ8fTNaZM
SE8zOqowhwgafbFKs3DiIjVfhoyQ3xxP3jK3ELwjzJV6z6SDT0F9lyQ65hlHtZ7f
JlqK8VWYS1fP5+YccEkZXyaiEsYOPrUD+m8Ex0fSJ3krhHG7UyUmebQUeeAKAf8a
pUax/dmR/tQiVdV/8cGYqviRdNOlH0XeJPvFEZ3xj/jDf0pMJO7gW8jN8SxUV+co
rr/yOpfj3VBCGPHcQx/XqrwYBDwHF49TChRZkRzNwSb2TmhA2Rhmtwqqh0TECbpn
hg9HLt7W/a2tuOj2/BnohHP5RekPGeM9BdsTp3TLAg7sjBTwLFi7X11AIj9rd82b
pA5cDLi6iMM3sDMsca8NDQK5/3NcAiSXtWnJu94cWRFewUOux8YspupidWe1wvaq
Zj+hUALgkStdrUKtRWlVSVdQ/Eei+5FIqnQf97AVx3IikW9Hdxo+CwY9m08AB7pR
d2aAcsxeJ5ZFMTPj1NNG4TRisFNEJgu7DG0r5SpowYjO/nRNfXHRANAwTcP+JXRy
SA6pWp8grK4OqCLVSCgtnrCw40p5ct9bTJyYVQ1PymFDaSX7SygdrY0wK2neo2Q/
JcILJ0w/NMUJVsn8Y89CR+0kG9Nb89BOcJ6EnqBRu1mlw72sw9RQidn3eTixTcPB
Ynu0Attvt6naixCLU8P7CQKgq8JT5mSra/8JecsgFSszdc1Rul8KF/9ZxuVZ8BgA
FCWRRLvIJy/Jg6+dGUUAAatbKEMRMei00j1ZuH2mFYjr/t4/ZV+0E+gOVxsAOxYC
RqAPTkP8AnKn2tK0IpealNTTWc9T8xwx8YP34/zslGOIAM/OPx9+miIeadMSKKJd
eZMQMxokxGqjiAZcpSxaxstERspQ2pf6b5BJd+mtFLHTP70IQyZZBRH58nbrNy6d
+5WmFlXZXe0nVQl/ALI8q9dBNioII8cVk7/a2D854v6LEtsGA4jh4NJsx9MkyBUt
vGoYPMr9alkY/rJcH+Vm6DEaFLh2INA/E/yAxc5BE4PgCLlkFlFodGSUUY1bje/m
imewN1AcyQowCIxEspmk8BioYJxiBQcpvBc5ShyUEA/Q/DV7GHgnY93Y0JZ02eCt
RvG1kUW6LJuUEK2ozL/CUZZvb9HKGA6je8Reu8P2E00chEQgOt7PtEpnnY5Zf+rG
qbEgwKQCBGaGnSmNbBdvNe5FZ6gonLnd3T1bf6Zyb5xmtkVT9lU0kblVriNjSXTv
Evrjn0gLkQt8NqpB6AjgnNmptVxsn30HHkkXvxP5wrwuwnqXKg8AGwGjXyqkbbmb
qFqkAcNNpm0XlqzTdTPsrmJHtneupAfSw3RQPdyguMJ8g/w2H2Gzb9mBBoCB29UE
Dsb3pwvc9IBt3smzxlu2VrRvSsmRIq4sf2KGWjtvSO9yG91F9TD8LpOX6oZQ9mm+
pnFh4n/+Zi35bW4J4FDudvFMbBt4DvTDgHalpjSxYQeJR0rklijveu2isHKXn7Sz
yos/TxA1ne2KGAGw7XOwGuSIk4xW9eWs6SmoJ2Ap+1tcXTj28MnNgF4VPus99myr
qf7GdoSeh/gIJTFQMMcLLfJhSQKwYevlpOcUnygtSz6yg72Xu/E01y7STTQLHVVp
BP7jqkTTewdSNExB8vb43O5Pdl+jQdMVhzBX6GRTvOu0bL0xjAuTLFQtaDGZHTZb
VcDLV5JBQAXf20qoS8aZETfRZicYAPh+fM5iegNuvMiNotCiBLm4n3DTtxrgZx0x
ReITx5i0lN9L6ZJrMMzl8QlhDZc0kvuTPm4+TK4Mu0TdJh9Aw/Dnw4uqAVchss+m
ba971wGYp1Mc0Ip7VNRMLszJ9rv7f/Io9Au/HTv1qJ3DbNiVer8aI1wshHEA47m+
/aA35EAOGYBvLEqf+KfRSfCXOacnmkHPThSnsZh+2aPBsIJcQNSVwtlmt62hVLd5
exmXF5uCkCMcmCVFxkSrASxGIc8Ffc6woiEjqWnrES8WjOgxElSpdhvRHt9NhtW0
2N9249+5GxCTg9DFZdvjcGsUAKVtUmbR3Z1XY0PQ4tpIL6TSFLz7YVMG0cDRzGwX
/138vK/pUCn+vQYV5O2XHg/UNFqfwle16nJwMuuuHUCsl0/vCrcV/aAgMvQW632C
ZEpY/EaAMUGKLKlDv0lRAi8CgHao+2IdT8PIKxD/XiOqtvy7+NvEC1V+8+LClP8V
qrL5HDdYkzEbrpojfrDu4cvGQYhRRgOTCuSzBxKgBudy6ZmzZz9vbWd4eGcB+dWB
zPSvftJpCakVe3PMO51A0kygXNukHbKaPXbvL62Q7KootAYP82dy8Scl3ruOAdaH
4eleCjTqg9rJtKSZ5v24up4yhLoy3JWiS/2VJGIdt3Onj7PbjJQBo88eSh8m0J/H
pM50/vbLf6OxGr7i9HRREqzzoxvbdH9k5aEnCjxpMMBpEVq7vCS2s5EzLEybwxHJ
GBekGA4sA7Y6+/QpL4/BfauGyly4Chlw34+giDBMSPyZOIToktxHa5taPAND+8+s
TsuMiy8rvzSzMsA9dPhrPa/5/FBV5HQNI9kttzhixVbe28PdwdroxUb1FCLXBb97
e7HNqk5/pP6nvL1B5Y+Zb2QSdMjztBjyVNgReSJ7nCrOJfqnHFgi+RIe7iua9kuY
MROu87Iz9AeWMPzSZ98QWUpL3KczmIttjvhVnT7mabaItxcWPC0/aMn8TPpL5g4X
wi+RIu0pTZUzdUeJS4nyE8CIMCWCAUdcGyoI3unglfSw8d9GUHYaZg0+yQUN5Ln3
mQ4Mq2QdCz2MzXrt9viW3+GVGKxO4HjPVrJ3/5788aGL1OLTljLg20H4jqJlCsmk
Sx7ZA6WkC4X8pmvuInd2IF+1TRCAF8hNBJ+eqII04Dzgl6PNcQoi0AEI4W8IwH7f
EDZZk/KXrpQ9L/Id/gohUo8D+ba0zOTfLAHVosnzcELRFnDMKkMAczKjpZokGPKm
a0aas95BXubNENk4BQjX3a3e3WMBFto4BHnhm8cJ4YahiCSWChLEUAb/4y5ASZbK
OcOBdVLK60pEp9jcg9yfxhRRby3KInr6fgyg0YMW7xh0IDrQWVI7LOGNQk2S4CqK
9OXOSJ1M+5+SH2ZaZjvQ68S2aOAKUIKzrSUY4H9H0wHnQ3Yjx/0T/2iGarN65oz2
eKxslkg/92N1g7T5NnBEojH5p5NagwJLMzcJpkNWWo8eJfEMF7YutR+b2SrvcmPU
hEItgRE0NYFQ452hCXkptzuGGWH+ps4C/tiIeddX0U7E0VbcQO2CAT7qxx984ZI+
qg9ebFyG5hL/Nctf2AyRxpLIWjV0RO+BjqImhr5vbRo6KeFiDJaUpY41tWRxt3Ze
N6vEUNAgUI03lwdpfb6hrxp1vhZXS1r8yv+Pjx0Zlg/g1z7vYl/Tu/q7oRSsUapx
ZXgxS/akzflDcRfxqrEP3i5egCfOB1o/FtNs6q3VxlaPiXPZEK0l77SoaRf/kBz3
vjwwdFN55ywJHmIL4M4i89dQOSsECy1r9bwvExFLKVa52nxE5TVGFqAKeuBI0/q6
OD1SrscHbBZoKEFd8123X/MBMR8qJ0r4t2SCQgO72CVG+SIeGcexXssaFs886iRf
t8DgRRIlLubs124pmGmq+3Cxef5i/abw48qoaw42M03MVLIr8IlI+CBc20Y2wwQk
Osc+HNPwLb2kpBttUSPJvop5EEIPV3lwoua+zHXM5Kna0NS2AjS7gOsvcVvVdyyd
R1cQtRJNkNdy/+/3bLfSD3qtQc2M8MFON7+rhEhFw8QcwpSFLIdTt8mhvYeY2UCv
ihUDNJxS+DIZctelS+x0pxoU1yNu5c3XeAd5OooELTfXAutI7SWOmvPVz7ooNoQx
Cj77aWr4jkKWLI2FxV6EkRVlH5bQ8ECyBiWUQWiPkPQhLWJ380ZYIaFQXmOaanrN
QxxDbelslWf0DwrI2qy8nA4p1+PhOAz74CERleihnwKkrADd/peGjtlwsg8UN5MW
YdUsbNoh7I8bgRjGu2yHWaSy5Tlw/spZfJ/iSvvpUoIGR6xHQ+TePWoELLCGJtf5
z0+1QnWyjyJaRgN4MOGqo1/uxuzwrHu9UcaiDPZk85q8wDaTjjPd/B2hrDGmFXea
Qvdu5Ni5H4yecoulG9z3JHBe36NQXsECaDaLxcXRQyNMzUPGO67EN+d6k2ODvmgn
eQloushbHNY7efpRPte19q/FI7Q3XMyBJ536Agiq4H9SAq1tSAmJqldHr9qZVzcG
xt1EFfJN3RPfy6EpsvO/fultfxqgGfcuPjBAzwGNzPb/tWv7V1E5gu5XMB1A/GkL
H0KFLgL2ovtoX8WZDdSj5so5w60QVVefLoixzqmAeSPrQET736ipWVcsmsceND5Y
m9tSr2eY34r5hsbWsbBQyUNemgAZCB6YTjTFYrcOGYWOXndiIhlfOsJACqenkLAC
ksRCN5ae26WD/WaxrK/cgOG3cT5+jQcMgUm1I+kI/8zLX3GLRA80yi8ay/+x8opJ
dv4tAx3oqv4o5cxmHkYyHiA0fa9sTikykuBkPFSJ5cgUihzgNycfaG38qKBwPbLs
jGyD+j96U8Jjxb2Sa0yo0GC4EDbCQRUxevcgs2TZJUFsUe+ZylfqMoRynTIyR1YT
5kfP1j1wlMkR+7qfECt2NUzFIZwjR3P4aNL72bHAnOS7OhMDpWrkqZpoRUHmo0Mj
ox/FHilFWSdQs1SgfDGcAUbzWRfeIuSzqT73SZdkObVMXG3H/vUu/TsijXiCoOvf
F9E4dm9ldTH7YV+YeL2ZgQJS+FHk+ggRE1nNIq3RDZc6lQnU9GqAv9eFG2w1yVTn
xiw1Gw38T1eTEqyxcjz0UPHZ/N+8JVgou2qXJNe8TZbX/bvCKPJAi4koiDS/bvoP
Acv9S9eAmwRUZhfVQd+ENAgDS7sI53FsHJawJm+y0n9prWcZhRp31HxCvFQ708wJ
FC7p8QGAIpV8kAZQXUJPl+PIl2oMEGDtXR4xyaKJ5rblfNHsDp//uBFTOdXjE2Cf
NmOc1Pu4FbBPjAy+jBLl8gWd0DQ1Aj64G/fQYFVuh2gmWDvcXlwYVU4S0LJHuOIS
RsKZdsf+U8PhVOE1h/367Bx65ao24rpSGAOlBfEHZljbOgCbDhi4+4qIayqqJeWR
Xq79X1nxwBUKwN6gAxR8C4ZQ0Kcdxvm8EacksDYQUOKyRsvTHE7UNrBj/3ADoLta
mBzItNDVvwocapSULkCx+Tju1WE6ZNu4fjWfmzEdpzbVpYhHBD2p633i0aF68Iiz
ftPRYrR8VIlYEDUDvIaMmyfZ1m2xNa8YU13kiVoZKrkUDx6y0DhqFVbDNEUso2tW
BhdOzzoJFWyLaVqm8s40due4Wpiie0fPKSsh7euYSsuoFdSigfiguNctC3y6Vjng
ysaZKOrsJiONdECsqRZ7AdUTp4hpqWezUrU9yE4txRJGG2DPgDjcTtWmdAUuGsN5
5eAiDtMd26AQfQUhRC11KmetHWL0+jmf516LPlNR6XjUgiQ0EioUDlGQSRBr1xIa
D5W3tSUB7vlp9GrxpQbd/ll6AySJe631R2KBiMyyAGxFYarrqudrN8rzNSABCykd
AGlkbRKjqa6wxyNm3r4fG3XuBD9/EwETdl609nOOJkw7HWM/N6Yc828w09F6or9S
T4BGRn1JKJL1olKro9fV9+aWqzTMqs7Huywskr21rG5nmHZ4ZM+AMVpsoR/ZjQhv
y4l0cOolr8m1wlQ2IbN2g006FzjECEwGaz+lAj8BBslBlM1rcr/rkcM69RnRKaX/
WZ/f8tJDfTeg1Lu8GFHHJb9El9rezt70mBNNYCWZstYmssY9noFJizM2yysyx1iJ
PXA4uH1EtIpqvnjw2CQO09MTBOMhp5U9BaEO1EUIjktlQqmHOHm3DqGzxF7xTasy
zHnbOMmvaLe5X74NFDmKwr/opDHHVkZji73nFz8oDnZ78t5DiswhMAq1RE2Hr338
K8XBW7rDzVInGF+F37bKXOVNSCjfsXeJ7Yc4IGmdTP/9yBWGavi8DUPV/zePKrUR
7v8zR3htJtykg49dBqXd5xW00WPy+HuWUE11sVBMTPYvdycgONQonr0P0GbATKO3
LFSABB7G0O9Kh2PdfXIP5vPZ7qSU5Y8R48TrNys8nqf75QgW00GjRYjhd2QVEp4b
IePZbT+DB1nVZHQ/hrrfCNJ5+rg+VACWXnUWjDXVPgo1WkK0kAEcEl3hxMAt9ait
iUxeP8n5f/Oo9OjDBSoxIxFiP6OTzefSzn08l//Y0EGYGUCUEfDgn+yFMMYUrJrd
O8vJHl2gV/yEPtKI36Ov/9VES2nMbDOAW+Ebwk4Wu41NWFRvWq1mVO0hV2UM7DeX
LtddJAemj0JiR9VtxOsEkvifuf12+v+G9fqCaLUKQl9XsDfMQQj4/mBPeyEeCkWY
ljY60AzYVy7FgUprS/kTA1Of3DEoQ4psXEXbzUrDt9+wPvahnXT+n31WByU7stVE
JL6J9QMtydEYOB36W8rWX/D2sOzkTdx3kudAf8fvXID9ox5Kn1TZTlFgzXA/pWWM
W3LOdhcTsPz6msx3P3RFUjsj7m5yuRlAT8ZP9aObWCxW+XXfITtS/KMjVl91U8bW
qOFm+t8X8xdlZ+RHfxHMDc0a8mNMsdAZncuOh6ogPZa68V3aKbxIOqHlo3hdCseu
v4S4EO8K1a6bAqhKJuLIYBeyPOm/ZU9bOuGsU71k0Utm5NXUAfwiNEQROCJNnLGh
D7UvljPZe9iQJ792I+90tgkIa2j7NANCuraBR9lYATga/5cPagvLLbdmC+n+bBOh
gJrvphRgZtpFcuLq2Mfs1t8IBmA+xS9WT1qWUSHyOgG8bEXa2mFqwRvjIVqpj5H7
AsC2cfg7XAztJuvPa1UubVdNtoC1gMgtreS0t3p2vyGYvYDgwRbb6TZFk/eJSrZp
I0u/fN1V17+/2hsxCoI+Q39Ywv0khLJPdUkmuChKRq41pqbIn9A6BVAGNoRSXWaP
XbB7TweLTfIpuOIrIk2Jhb+h2gUbm027hRvo0BzjRQ0/ODgx0wGrCTQl0K2eff9i
3TPlEm9wJZcogBoAeuoGytc49lxNsGAF3x1vIKLMrLQ3Ziufn9AAsZqDRjhxgyzk
7t3wxnnKPFh12AmKH7SgrvJnOzFg4BaNiFJt05E6fKP62K46j22i9nmYPCIS3Aws
47XbII8Jdr1wLkeXMdTdnJft3+Pc+yUuo+UNThf4yd8UTyHjFTw7qLJVcl6to4Tu
bNtqOeMdptYjHBy6hN6nob5lC+mqndDJpTlj2REE0WS4Q1LBHEPjt2BY1Ll/gzGo
3dfnMQ1IIRyfIN8n/1aViZcUgGpZUIMnQc31vIaY+HYX/6zQGa7eiy6Gkn5PFY41
PnGBy3x0g2BZFOloebQo762//4oABNIVxnpxwYldwpilAoV1w08dbW31NstxSssz
xK05MDAYnUi2csiwPGV9E0J4eUeVYtwguJgIlPfnHEDrDq0aF4Va2a+cEkj6rFKi
F6cdqYGrCfKZsz58UAh7ojRXgD47qK+Cq1GyY4ano0PnQazS1rPixsQtV5zeSWD5
7d13G8NygYik+6O6je/T24pRhsnknHihLD3CMLCBfz3I1OndNfMIaaS6BwVYT2jo
+d9XCkb/hIxA/Ru+LIdNyVpXgjqtt7U+gFCxLnh+qpU0pUGteMm2MYhyxCPMJG07
wbVN+MSJD3EDBRzNw7EWZrRgvsZQP0mTg2ClB4/f1XzO8Pj2lzG/R4sSCbyri/2d
DHTDFy/cybQ1TGJ2YMnemtJXNYh6yE8wtft+AyGFUD9JTg1F44WfofrAneDhhfg4
ioUhy2Bf/Lr6XiP793PJWSJvIBiAn+PcwDxWlyJczk60a7aYXTvgCtEU2ktauumg
Rnr7FVHC1AWZlu1dfXAVCOQ3VP5t9iwr3mdPmAgPYwOuQfDPhqUHOllx2zgrNpbO
YbUpt6Gqe18rMYaIwUjLccewfo49m80ZJ6hIfpzbg1Crmgc87EiJDHhqMS41ai5a
6EuyliMBvt5EDWLjn+iDhpPYIPH3Ls9S+H/FcprQTgCe+3ly7S12mFaUdpFRGWiB
Kau3azuFZZinwl1dDNV/YPqeMNoaViKKhMft1YOvgPshzlvkTw9YrinUM1LwSaKw
nWq60raJdEAHSAh+yGKGXPLMSk7l4LpdwaIiBjn5rBn4Pis6jo4uLzbAwL1p+B0v
wvPMBI+7F0kheV83KtRCdu4A/XKyFv2In5QNKF3IuMaI0ipbAzJ3KJp6D2jRpc+U
oVAV7CCuaFz6reGYFYE13JGT8fzESBWXVKeK2yrcOpl/exqIZSiYWqtJSO17f1/S
191oKPBFeC9J+BxZ9HaYGbsn2wWBViag3j3/tRYFksbXxav7TFCgvqREdooLsidQ
O4TQ52B8c3Woq7/uTiRXIxC6lta7AUnbE0UTcjI4x6JfVkW40wLwH79iiFcpkXYB
LKZWARZVFdFVllL7a2fIoMINLAVCU55Rr5tF+DAufpdMb4MdEeutbq4TCCYm9GcR
w9El3qM7Os9M/sR3Szz9/3YD+pGy0acj0OZmDYSgSzZ5S18hPV5nH5xTO+IqIgPt
u/FbzWeft+KZzA7OYwZTIU+t4kUSi89WAhiCVBMx0RJh6VjmiO+5NhqGBe7jVzKi
9710eHYjNWRb1C/TzTn21A9AgNqiMjjekqsWzr4bnxhY+QDD6+8IwOLLH+XUL6hY
J+qnXRIYd/U2ehN80GVpSwe0ZSN8p/HfRcxGqeh71mghEgBWBTH5coMJnsBfbgPd
w5i0AZkhq/7Qk4vgsxYWXb0M4DMIQQb3qGMy0M3ZIT5b5DGgJ5BQx2yzyZXSgdYe
UNVqHhBOWEEcPyX3x3xkwuFPTOpxrU1laVKBY471IFsFjFWS7SS9/TmV0oYabPO4
tScM4YpsqLxmfSgjVEIYCmVLYEOUpVM/1EVM5vcc3kl+txAa6X5ZdgYw7lbJayy9
vKE132AYjtP/jAyO9z4yJdqyCXu3GbuMfJwRmXYnWWJyz5YMJKndcmNvJskm/8ao
JruXVYfL1cKO0hCCm6mccl86m8dDTetyVwMb5cBEnHy06BUANuqlWcR7fgdt6jLE
3JpyAxXLBdBKFmPzqYzdo5ioq7I23g1GvjjlP3Hn+J1gfydmqBwYbXtbpjGaEhij
XgSjqfEFm+rudWQXbsd/gLYjeYqiLHaMC6uI5RSzZLj1+aDRMYi34r7n6y8ZpHj0
17ksb3QK6p7eSnLad6ftbaBWwmyJ8ocaQ2AQCfJxzHtpG9afauDj8+FnyX+2A07r
LMzcWFD5/0v1itSu5Lr0YSd95vNKYcmpPgtb6P3iaP2ucd5wsdDb5dTXcRU7uqor
d+a0olWj+El+0tsQOMYbvKsZitIIQQJ8LQCLosBekC+JEvcQlJGyhSJ7CCCuLU3E
Juq0LAWpuAPRo0c8bGGHhSd/B31cUYThHaU5Coidy6tqID2nJRlIJo/MzBsV4oCN
e1IXMjNh3LCxgkbjCQwO8OCLlclVtrBIvXh78SNXdImrHE6FfzfjIEaBEvVnHlWV
cMvGJBW2GtrNw8l8rovvdI12vMAG3lpbAozzaivhSvpsy+X9iSLF+OvQX2JkSvnb
QVh++MfOM4qyTVCRXvKOn6nIaziZS42hI22cMd2bPPLbqFbu6FTjguiA/mCSsmXe
CfOfbbNFrOle2tUz0yesOJoqUW17R6DiUBQoZ5SNHmjAca/9LNZKYBiEsFC9DAFX
UG0vagvJhNOsF94ahdbukJ3ikvFC0F48HjpJ+WmAW9nk0gSsbAuUh2oIbysMoIQp
ZuSXr2XZuLwZ0OeLTOG5p6lcXz1idQg0O2Vz6xiqRkMq096b4RrxDMBtmUBtcskf
Yu5hWYftFSn+50NBzNG24NAFsp0pwFt28kqwVARsjjvey9FcLfJOxr9WkTrbU4mP
4PWiWCogQEAFr6gsTMtHJmPDPlpQrwCkOi8FYw/j0BhaxHJvYEgcr5klDSWFGeKO
eA8XV0QTW/FSnDZPKK4YuNMJ3kfDYsYzbEwy3P51C0afuoPGrSeXAzZyCWfL5vGG
mP+tqXLALPq+/+fCn9llSjR3wzxF/u0YqBr4VTUW95b4eJuWPtfshBfCneTV/28i
ugMLUZZuCRkKclqn/wZzX98RnvBWpHOeu3DLt9qj/zaJrcQT3FSqOSL5o6DyIyAu
UHQIhCpTCxOFMjJA4vpzskm9Zf45x8DHkU2WHiIFTLWKT+lVBEVRLwa/SwAQR9sh
FywuNTtHeasMqzuqks+wHjILVxQOdaKw6wX0uUzX5miKqeYyylApkFr4vVSLbloX
nBdU3INctkT5SSD+WsZopjgggUJS5xV7wjQd1VAaErt5/89bzApxC9mfmpvA3aJL
uAgFpGA7SvRQkY1IFNlfubUXJXx+DxBsUoyE2QUhL8cmpeBswditfqCPbFeQmhSc
6v3nqV8PZp+T4a0iqkHIEt4TiSMMjjFFByOCSIya3RsCkVP2s/nTj4h9X1DLsD8N
wNvpuzWV++SswaTnHINgoVNPyLkVTQoK5OmA3oJnA/i5rqHKKFWAB68i2BOLYs0k
hlXztuld1DOwpCely1l+1mW0clotkL7bJgRGbTZXURi0pIjk9yv0ub9ZBT445FJl
2sPem4fObwqEnpqH00qP74EytoiwDOwpZ2gEBgPesCBFB4Jo9DJhCiAbZqYoYyIl
2kwQTQPGh/XWBCybehS64yaiBIAkCLFkRMYYrjvwsD/vUT43KdBdXFILjM4uqtYf
vmVczXWVWN9dFCm/bpfne/1eLQNEEx3NERfcHN8n1DKf4UIpnViBMDLC8GUdqUoV
g+RUOWoprT/6zxf5E6p9j4c8IjAF5LUVQC1DWRZ+VA7ezQgM+57eIb+391p51ByJ
ZqghlfplGGiIIZRsdzVjsb+vN2l24U/KUFF+ZcmrEB8BlBqKk262Xydz3H+aJx3f
eKL8br9sX/jGGTIIf33mLOQdJ+0eVRbl8iB6dFqbyfh/s8NzNECe1tYqL5wGZoAy
YIV8gYyJHUs53t+1rA/33M/pWVSgFkYa7Jq5sDW3POhLiULKBs2yN0Xe7bKQE7tx
HV06FNqwBw5JimJs4KUuuVgzGovHIe97/b7Wby/4vynEw7p26veItMX+IQWTRxRq
5JmDWvmfKOaxzTrEbMeVBYGCi0+bdBcY1Umt6CdBnAGc80GZfxv/KiKNJ0CQdb4c
KgAz+EW4MbK09/kVKgJ1rqQb0Ir9oA1HU4/pIMXajoCZVUqs7cHDxTIZ3wu4cTuh
wV5TcTxA6MTsbxFyXUvMy1dZx/ZgXhnAFk/KzR/rw7GLLsox4Dk1w5TREDt48JwO
+Zcrfh7cpJ5L0HYrRU5HRC0iYwt4yymc9DgD/gHfV+Ij3Q28px/8kDlJ0IKFzOKY
ye89BFIpTRdzcJ+GVu+eAPsRSeMRhCjjMIZundG2GKpTWT3sQNUzAHLyoXkv41Pe
YVzlpOC6yMpmzzVeTUiQPIdAONqIIbAA20man5JkIL4m56tzidUddq+EJW/f9HN6
uhs616LPmlrw5Y74rMfqx1HY5PsUsmP6G244TmwtLg1KsljPI7kXZXhO7CCNSJxz
iiJWddtaIhXFhAwTBfu7y9/Bg7/n8fYyB4quAV/slygAfaaTITvfAO52nWfBry0s
2xatw+CCzlEt0wq/k31mnrb8QgR1dVCbcD947QK8lELmREJxXTkOwNxs4BJ/qF2p
Q6JKAWLDgYkXc6xoF1XNhL3GrVPYMKWcgsYP3aBttJn5eT2mkDau5ljtYKHZHlmc
sO+jiF2yjBSuVGTmoRzW8J/JgqQ+1cYe+BWOcpWkwi14kDmraxXT3NW34wvMhNvR
YecaCg5p86P/y4E7sC8lnL+k2Q2l9PEsnftGzgkg/skx6pB0DR5XURufehqScwUF
WAcJ43e84q606AUYBXIhbOYum0lDdDHQY/rPJ1y0Nwq9R8WzVSwY2zciREHsOmkD
70gfR7VEnz7yBXu5gJ3PZRL4stDCeBCRIOp53wdJEzBOa7V8Er6wstvjax3Ta7by
yGqhw9a+hBHE5MlCgj3pyUHNgWp6PXdvbOrkBvFG2gi8UXpd7SJnsbh9nbTKM0gA
M0w0GnEAcV0uLEWT0BFvsxJr8T1Nxcq2gkSsA9+RBe7u+tZiyk3fajpLc0Bq/zlg
HSFPSaVQidV/TOiwORFhY/r6Fanb6hvLItw7iawgCiN8oGCUSNQY+tGTPi85boCx
4lGl2CAgZXkXpUwn0HcWs9bCjoVN+dm+d5oP85LonJHVFNk9BCAWGHgEdBrzs/G9
TQZv0u1KT7sMk7s50k0fN48YV18yASKIrMgoQV2GzBqLYOgKggKwSHPwEQihgPYj
aAoGL0TxZAZKv7H6reFasvR8ydvsj41x3NHsB1fL/BKh9hd0HSkN7yHVu0oBj+sr
/2o+EbtH2jMEkeQLYjpaEJXHgHE4BhsRQsFI+IRi/XtebKa/UAukGyEO85FODGAN
tPIOvxkbeLDeraka9bvyvVtkRulBhUFFTVc0nXq+pee3zgSSIJkxkH3S52wLJQdL
VW5KrqLXBZ25PBX9M0hIKr6aK2MS3Fkvg01lz0qJG0USRYffO+6bHAzVnCQPkdpE
BoLLAwZG/8XxOxVFuuBPc6vJ1RHqZJ8myli9fKFvsLuA8ZN11a6xWRWK3scdbQwM
/L/2Hl0RyK/WNmu8zMOz8DNK5bx1ynBHMIiK7rrvMknqZNfjCcN7eHBbdOnBSh7L
jlDJAt4pXT3lfFoEO+2Djd2bM/piC09/adLUelbjB89PB/37ocGPZEsVSzzQ3zME
bWiBxnitwuA6ZSpwwhpZqHTDn/3hOiHU8t4BWsuvzY0kic26mqW+sIJn+ad3475t
bURsotimoKceKY+uU5Ve4TUIklvFCJpMhN1iqO/mldQUcmHUDmx+4S/b/7yAshpG
Tx1SzYvpe28s09YyAvKs1P8lCQT1MmhB4XvP9J+8VLG6c3QhsKd2ZjVnKOu7LdLP
b7oAF1dTllf0g9OYlxpS+xSiXhm2lbDrfq13WhfeSX7Je4x6f2RcecXxr2t2n9Ry
tTReT0tg/IYh2yc1r7UPLXi6ZZT7qpOHwp0mlOv16m2UMhmlm99kqAzc5RgXEWla
ebP/nfd8aR5y5rFZUEOqoppEzgxR5pCFpusYMMa5E5pJXGQK5D8/NlZb8Hf38/7f
Ukx5IaNBRZTUkNaW32F+oYq/WSL6ibOJUA3+4YS/itEPxZ4lmwyMWbfkFId7Cqpp
phCn0Uvca2CiuobsDoGgVUgKTizIu/6bLY1/1nBXLXnT+Uebsf0ljGyi8wZaNec/
buarnFm4QWWS/ze62J4LDsK/Nt41NnzzGuqaDK87ALepr5pg5cwhGh62it1DraLD
E1zD+nR9SDcldY92sB89rcZC8aaJXPK8M5Xkd/IYQa9HO1C1tq7P+3aTshqHqjqn
bChd7VRQ3o6gBjb06zZvEww3/a1UWr1g6dyJrEPNGwWXj1X7AsKY+83iNeb+o+Jg
N45lDgn0EMm07LlmyUk/LOY4bcInT8sMhdN1PmGOBCjRS5KhrzKK+xnYdwpOG+/0
UZaWOfT4TFTBodW4FrbnzqVXqikYHJ3gatfzl0TvYjIZZxvlJo2YfT9ocuqw2Q6x
cdyVPw8VEh3zJqIasDY48XC2sG0hyr3+3YREoCqgOH7DDR02oDfz8uLCspxzR+TO
ZJbmETXWku617Yg4ND4dT4grQTF4sCF/C4neK3QfWh2t4lmxrv9/HnqirYliwJyx
5oIGoYAn+beXyHugo7ETP/zvfTzkE/2vQpHxBKZ7oA+SLOVaE6962dchjFLY1Mpl
CkccaX1Ov2IkQOm1g+oWlRIyZjQrXve1G0nj1f3AhUdmyY0qng7vN4Ek/Jp6Rjt4
uLm+1IB7GNe/+cCeS8bKIHwKmDJGf5Y1WPo6C3UvZCPH7OoJ31rQk4xvHYnins7S
2Im+StUwzLV5Q1ehbVQM4DEZCn8X8oY4oEm5MoMxoC5PajNl20Tqf3jUoS5Xnqp1
72O8gXQVEx+OHY7MkY5Vev4yyiyVVY+RldK4Lp1Zj4rbbjOKguAA8HVrq8bqWEAY
EPahVkhVpiItbCCVgXwYHG1lXgdmU7YVHKA3CHjSpkouXHgaS41la55agRzIBWl3
93UwxPMMIuv1wX4lYb7JMHP2AwlHQtehfj0rXWAkSETuxYekFwNpmd5SCIpEcni9
D1Osg8xH/IJ8gsXFJ8VjrAms4i95otUUtKE6d9E4z5xnXUkslVPOfNgWE8dnX84C
G/2lEnAYK6T169ksYdmOo272IaUS3vNroWoH0baNWUmGIR6ESxsur9JUnEYT/lW7
aRLV9ZZsMAFDjfZ7odAi/l/Gxyzn1tHbDUELknVyQJYzxWF3/LMwalRKFhjc2xsM
zEgSm3bRBGjvMNkwye2f6RkDhoabYwJ/zKN+IxloMOfXvgf1EpbeCrtmL1+nlNOh
ArlfbSth/R0rQMGI5pBpUJXzGSxOdfk3Xc0iAPLg3vfZM9Sf/S6R9p5D418fZa3m
rAztZf0wHGIaZgQzDcJwXhgT1HhjL5qrVWoHMR242GCLFJmpAMDThUmO8FMoMxFd
CivC12SLtzAwhaMS7g8e0wGikSQYO+Q6Gz6GT27MlEOp45wCx6HxC1f5C0lQ5mJt
QAlnQ//eXzDD9onNVxNVjdjTYMTcDuGiYPjXYLDUST/URAqOIzXNVaFwAy3BZ7Nu
GkroTrVgG6IXuLZ0A0d5mmIBgCX3C+JMHZO2B1bGEjKaTAjKN4R4Xa2Hvpov6xFD
A9RsDpO1HaxCIrTNbDgcyjQ+I6uPey51NdVjhYuqp2GVQDL74FKmbvEFZkUxuhGL
57ww1uXBkM8lP0+A6SIyKBalZ2pIft3YXiEAcVD/r2yXaVFtSatf+E6KZMyAIaoX
DLx6Eg61ASiHATJWeKcbGvehq78JugTSoSAoDC0Rcw4fvmt8UdqojGgmRmj5Ad3b
2oUV/OaNCMmBR79zzH+4IVgPMCYwdMzKbaRBYQ7Zk5o1vtIa82qP4/hczYd7FKrs
crvFDHknOiP+Tj9wcsqG5/p2h8qLpVEwS87bo2SO7qg9O0uvu9Zm2k+fdwGjfhRH
7JV1X+n1Yxd86Q5xDP+kYejxepSMQ7V4VHjKR94VlQydLL7l2vnHd54Ftu97Wo2D
NixFFOvlZ+RMa9eVm484TlSz9RdaEY5VwOVNFGTeAtqDKZziQQWty3P7FKZ2gYnH
AA8umxS1MFmFBtBBJ/v2b+KqakM2BP5wJ9hQhLJD8IhwtikE9+a7X0Zx9GUzha7b
jlz+jjUiORiRCorj4VX/1OXfK7t5nKHdOYTyIUfmSQ//AOS1gstV+1uuWBPlqn02
zsOaEfclCCU4V5gT9Ggg7Z9nd4UVSqbQt1yzVZjsZFD4xJLFvgUQ5fRETgLgQzyT
ik1Nqix2I9FL7DY9NvXcbhlauk0j+4UCu4cpgl0AZEI2LCRwEyIkSkAUXe2V1/o3
A+AnSdCcUjt3m2ZMndEIo0INMPSIw5eHyrvxWh3Metc1qg9tauvHRI1BLdVLzWCr
CwzSKVLoMu4IeSS8gjoG4ROBO+jA6I2kRSbcFSY94vhGzf3weFrSkQKXR3lZoySH
pwO8OhY/xF+asKk4GTGfRMOQpBCTEqhDXLti5n7CZ8YMPVI7FxBoFy5hA/sYPIxM
lOvvbzoANXhTgqTPnaqGZuyqsJ5UrgOZGJz5g6mrnPpHdOGylP92zDAv6J3gZkUq
Vp5WaM24unc/KKiPYm5/sm8kYWqApQfW9sMd3Xsm8Kr1TifKM+bbeXjE3eoeryfr
4os3CkEa2E/7Qcp3Ee41L4skpQ3Z+cfB6/xNEfTiSwRXKwK5hhKMmeBBhTdn83m7
FUi5o+XeJ8iC/Jr97zKUq9+jflmTfuN2iDY74UNKM0X77wnW3shVuTd1SVXynL2u
+as5aCOWNlYAQakyarS5bnUk2HslPhGKz+E8rPiimvEuNfQjtZdafxWP3fBbk1fc
v1YiOdlwNBE17oCpcbJSgIZhEUjD/Ibev52h8++J31o1BP4G9D7QFeWnNTU9aH/W
zK4pTWFOo2ZxFxElxFkZ6/L/wPOi4y/mihwnDR7dsIFtRFYufeMeC4tclUORjJvV
xmw9twV8g9kLDLxXAOeXtYZMn4qFwLjseBBPErsXL08nmeBavr1obhUi/KkQnaWJ
NHVNXeIkwjyZVvuJW84tgr0usCiOl8jeq1PgLnmPIacZg9Qt2uz5ss9fyq4bHW/2
lag9hcd3wpFWyfRWghg10XtywdXR4Oun2SKt1hf2dDvRqAp9Jf2zOqQGL8CpZX5E
52VuV3kmxgsxkZ8w68iDuRVs0pK5y+8x5wzJWOZbbXmgpYp2bgu/2xAYCjk7AZqw
2lJepqmoLxi6gf72uJP+Lz42Ng60rbzL73PRkkuTUm2ErY6j1u5m5t5WbMdz2fli
qtAGFwKRWz2BVLJeDjd6tlipe1AbzfsxZgqNDI7+sm3+nJY67wT0sNpB2SClrJ4H
cNNU30c2OkfIFR5Oglz+YhlJQUNRzMfaDfZZjKOtjY6RWhtAhZUKvnShhM7Lh7BA
C/DgeRPAuEa5rrWF7kbkdD4Wpzyn/95Gzlvsd4NLo8y7xWOVDiZ3CRIjZy+aCUIm
JjncB72mUJ3YblQKcC8lwt2XWO7quwkWDJi7FKwTrypKp3tUq+aiDfCIAw/i79Aj
RPG0dWRAnnZOedP9vrzio+ukSyJpeWmVi/Qs7lREuHzwwa0CP51EZfDAQPpuz3l+
bmbxKY1JOU07YT6maMVeHEL4+HQKH5PKbvTvtnZJFWVgG1PB1PqsS/f+/EWXPTxB
Gu9nLIkvd+4hDaPxPpkP03KGbma89X3tovX/x90yKIU8oZS7rAU+pBt4i5hQHuvH
5MJzOM0aXVDcWYwGbtcRoGf7c4bm4uhiRRjnWz/TnoS77zh5UuSUvezJiRrHQ++j
k9t5SCPJoJRqqbO13djk70bbXgA3cR+zCHrZqj/AagPlqHVL4sjfRfJDw3Tn4Mfb
ZrbiT5OCdoknCJMrPtcb1HqyacMvb7cEukAe/G3zzg8TYCMNJVYEcJn7YGEvqEoA
RlccWJhXxfiyyuq9unCAL6ZRLVY3/zInyJG08S0kIj/l/bF5x7aplEG3ql68S2ww
JVw6uBsbu+Ym6RuF22NAcKPM9hETaFmdyrLEgPnUSvrRb7FAe1LwGQwO/5FLwB2f
lpIBG0ssLZqD2U+FFqz3Yonbyz5RunMiETk4s4T0uEr2ts8RxCdE+MuHTNiBBQPV
NtIYI4jWDpl2SLSQB12ubErxEeRFnUlhvbXMhgDJuZ5ZIO+kxbubwXRTPtOcwHve
xzla/iCISlzoy3U1nRrd3Y8urnMRnmCPn7qVRI1yOByAk+15DRP62j/t27K1rVjX
/wWtHaGIJRinYxcui5upc0QsUtNhDqhs5EASfivGkIYPHy7epX8fa0UJGlqYtga2
KtrdY4wvq1EehYibvkkWxFBNdi73DHCzwjvp4qiGDtyTtc/oubumgoE7lt3iM7Qm
l1JDNckYUbsfOvakfqyWdPuzaAsJdJoDaTAcnLVF0CkjJwTlc0SWD+l/EZdxTlG+
04GcWfiK0oVcbfcpYCVxXmhjNXnPdjp2RKQmTtPe4urDj3srh2LwRqU4CpHzsFRg
bXcrNoVzaIqj2f/L7JDYkia/Haul+epjRrIgi680hTZ6VTebA0O9aRlN2C30UnTn
9++b7FKOEj6D3eOrmkPqu6aqAGCAh83xMsRu5zafX+EkHZgQRy1u3Q4VV+FYrke1
/bIFcSOm+oBlR6YZhSqnVTFN8bg0jTy4n4fwZtLIGoNAhkUOuxDusjWUR56cD9Gj
c1Tkdh4M/vgalvI7a5CWdIWEJrIDQgCrxQa8/xPuSfE4fVOuLDG0p1JTkOuAjPp7
69I87ylzXp+XZLf/bn6FyqZXgO/AIIX0RqvS20IRRGb+5iY6qEWCt5qDZ7bKWV/U
+/ItQ7O7S3X91uoUdFtxmb2osmU6DDgtM7Uy/A/NYN8/O6eWOfzS+GB/klDRUKdq
wkdfZYpCVHLL8cxJV8Oef8AeBIvogC8ZclJJMIyPwiyyWgVZ4OrsiVCa23pfuV8g
5EtlIQ9ip1BLdPYb/icXrmjhpXYEid8cT2mzV4BmyCzWW3wArxxHMC6G62lFIDUT
yu2//+pJeee3pWipyNZN6Cl9N2AickK3A46pCyz+NEz7K0b1bx3Gsd2wZZQlkNy3
keQM0VJisEyqfwb5AOz9MzemSW0ShFr7SiHq57GdU/S8mjg+0kYzcgcyl/wGLIgB
/gLbfRJejmcCoDK2ycgy2Vs6Bl1mqLZlzJRTm1QvD2mPxNRQnfY2KSQg2ZalvS24
Lx2TWQEatc+Z2zwBRSWOddLC/uUhS1EmxkRLN57MDPBlTk7zx7CfuXd25wvnUpra
BnMKU/CLeLMdaubrYQBiDrsZw6PrRcGWZRsS3gK+Bqssug0UQD+wW7uCQBk9friX
z9lj4ztlV+8nlYj40Je0c6M3XDhT1ERvxu76EIBDRPvKIrfx+5vpgBsQIzLwwD6O
5zSYhVomvndS7Qr/bbYD7mnGPYHqAI9irpDxPVJML1LTc2G50mUtD251r6VmypKY
Lsw7JKw3jG4XWDsKArMJ4+HaAB6uTi8+m/u12tcvNjTcWtP2MaetnxOt5SIAjFLJ
B9X0DfkN+0Sj2udlm/5oZ2qSGEpomCk4tr5wQOvAcR+m+TtRCYaTntkmPQpRTP5c
C3j7ssyR+cdCtmcRDVdB7rMaZeqkrHB4bR1nvs0WqMxnYpnX+pSvo7WI4EImbc2L
EJ4DaL5wkAUM49DmNRfk28PxJVhZbaN2Y4Qnorj8oe9bNlS4nvVu9pn51lP4vQ+J
v/ejJV3Q476+6Y3/Ww46YiCJ7zYUtFw8SJ8fyLtRG7XOPCNAifWhQBfoRgbxw6r/
kPE7cByDPzuSIi7NqSAMhrtbsyRXKCZ216KiAuHaaGFhFBNINYYsiQkmEQydR6tE
ArEmkLL4uXXFTb9Zj8w8kKJ7C3WwCe11tTe40q5QIYV0flaKGeWquC9zaNoamfRf
ZBdIPAKOqnUyi4X0n8nYL2wnC+lVC+/myjntwKys+V7T/6Bi2mXV3xYvJmFDKGYk
OUOmqeL1kq4KyrTrZINOpUa8c4QWDlCSxKnqsPTuzPjcBzjAUh8tA5Q6rxEuAHpJ
O12OGNsiT826mDKo0+GywrCgVpgAOSO2+mRawW33Yar1aQxHiHwrDuHprdagM9Tg
BvdE3nirEoKFDxPF+CTXJpqF1Nm/Z0jka9SL23Ez77ABRPwQ/MRuuAhiv3y/CiJq
RDQ4f/Ggmlqb2ix6zpX1iX2rlGJC/vhSxkK4YDiu6w+tVSMrpmGcaIa77GvJd2zK
+igV2IFk1H/r3J9l64FZBOQVDP2fqyeTwTmSTdDkXv3FZ9kZZWiVL7HA5sUKlo2C
AZZ1ZByYQMjupG/8ZjNjdi3W6Wh663DN3LntEosIRQ/KUw3ODK+na/cBM09IAJbP
X9KFQcGBsTgRIhwnWP8E8z2P9s2XLkaudVEINdNnrXr/Kes5CWjHhiLIoNi/AuqQ
j0BLSAFaKxYXK22OWT88QN+gK+l640p5unOzPAOKUua8DqaQ1ftWMehkR+ckjV6W
nHDGp5RRwJ7G7kURUdcYAiGksfYLmexmbhxSRMGUPS3G4BzgUi61/HNco83U4a5m
Y+Z4RwcDPRJNG4j3Gic8IRkynBrGWzLMTjPv5mOyZmjmyNBU8zNa6qi6x+0Dzn7G
vBtVALfDYgD4uzGP5x2BQs7QWgZVUD1xBQdgY1SpHoSALd0oCZ2iJQLSjuUmkjK6
5p37pvLQTvpxUt/9pMlEpi6ss4bDdPqgyYRejTmP3xm0B5RbMmdBe4yzuAJYa9Ss
KpspctkyXDPFCvYYquuyuKu1kJMVXtT+LWVrHgXNKG8jCnW68xM5kLhQunYFdnCi
YLInbOj8YdwlBfFUoZP2ma2vY9hd7x40gIajFXcAUGuz/ZhII3tL32l/qj6L0ETz
BdNj7zw2e7HUGll4NU+slKQsUnX1kk/WrSWwLKo4Bw4skkthSonQE8a0coGjsunl
bUBCfXz6R//E31/GNP9G1hhz10VPmVsjWU/n9zviMRqzQW840qS55HP6KqFPYkz/
lx10jc9JXq7BADbeuG7/IwmZxXB+bCS93Jcxwhbk64jLP9WAOFfzl0WqjM17xGt3
6pRq+h1AW7h04oaQtvkUsYNn/cqM7A154vBh41wtrCkTiV28E4oO/+5ILr1RLXuO
VtrHsW4dNSLr/jWQBn+Ujm2IGxnuSXIrEedeuou1DFOK5I4Qf2cLflWQPLiJrKlj
Meb83MHz9f3uh0saamR3Hd8IvaeRWk30apzLIwIIgbDz2mB2uf2kwhDEEF0+L9IV
0eQLu6KDICbLx3glUuKbcVg93+ZraYqnYDuwSOmPm9l6pLtfbRSJmsOMdMV4zIo1
4amv3Nx5xArpkxcbSWaL8vHkUysrwIpUYWkKtr0UgFKfkXfsB0WbIB8pzg6jLRXY
rVohMaZ4FwSoHyvLwoNn8EdM5HnzA8UuflAAsdVHDEPf7b4m2T/doBh41S7xH4BM
anuhCeTeFmZ/SrIpYp0NrIiZU7VVdjm7Eoy9jqW9P3y2mggdHQpgNSLyi44Hzmwx
6/u6kgEgxw93uCXT5EqsmoonU+M8QJqOvIDYWy7u05Aj5Ypd9YXo2IunCtnSI/bR
JvsHAoSjXhrqiV1N6wmzTFqinLScC+bxQFBGszz6HyBJ/yMtHTWYzg5b5ujGfXeJ
tn7bWtWL50GGatBbX843bG5D2xfIiD+k8T3RWHyLqY/E4wMcfh8LxxWYO0YsS+nn
A2ILy+UMGW3Kjx6Zp35/KheYjXJhKHKni9HsP4sVVSQ40kJZtGfNkESv0rcs6RPk
5P9nOMhzyUfv1vdn+UIPKQp/Fzu8pl5AwrnOWL1SEKu03ZpzM6SP4paoAZ0OUfgg
SXgWV396TwsHw+Gluzc0BOBuMBTQo3zBp8EnV5/897VvvRNt86NKtqT5buSPpSwA
AYgc6EIoGHU9wS0Z2A7B1U9am0v4k82MwsSUfPi+qg72Aour0YvRjGpCMM7oaQOh
7g51BWhMQY2OfBpdzzT/yxHntYXAxJD+OGZbsfWqaniVdYrEYulb4InsSLDL6Qao
IsLtMLLAAdwX30l+Mo4wLMsGJPdMzk8mUcsWYLpoDa6m1DnVErnAg3UtsehysE9l
MX546nK/iC9gW/YpWnsnVzanFmft/l1yBIiKxhxBb60i8FQlsjRfBUZwhtFhVbpI
QNirT3//r4/o9RIV+DK9LqKvLDBezAm0rbslRVZoSiY1JP0E5P7RJ+kQ/iJZx/Yb
Hst3tS1WEXIdZffdJdJNF57/RkcFwRvJqKlzCjC5NL41psQnp+mi98zrFgr0vPCM
cN1Dw4pkqPLsKX1tnYvkSkaln/meCtjlYzPnH5BfxAoifaYTfJyLGMZb9/DN8yjL
W9tXN8ZThKXBYPF+CaykhrydSsmPGvR1siy0xHOEkZcsgiX95qyjzE/hHCEF4kBu
QpRyPb2sWI8akuf/q53Pr5+Rfo+DwcNs/HZzdsNMl0lKbl8freaOoJlmj2mLjTra
bYJOlP5wXfTw4Ac0gnB0oFPDvTbJ+t5Fxs1YZZS44n9EI5tGm0Z6OsfVRsVayV+O
B4AQ1LJc2xS3475E5wR+1R+STuu8xUxKnnh0jSp9i/JxpNtYOatZpXlg7pMZKpqu
2mmH784v+hBHLWMR2BHLYGHzq6QQ/Kj4bcCV9kVFaPj8VbunbGBTdLRFIpu8rK0w
c4agN/feww+kibLsG1krc/fR5wUgn0M9ygz8PoIokECLl230F7tlrAyn1kT2eJ//
26od5/t3d3CE+f1yBkk/DfxC7Y3X6JMgNot3m/TjLeRXCTLv5sVhHRGQSeyEqbDF
r3x4U5YyAPwJMM0t5r6mUG5w40VimDuGSDvYQZgSf2RRjRKg+VP8Rw+FVHMdyJX9
HPWBlG2SRZ/AAaoU2cUy1J54BnLqXRucl2oYv84CP/GrygSNH8gm0ZiuAbsaV7tx
Sx86xbS2v31mtWgTewxE31Z8NrUe9FfpBxV3L3n0MKzWf3+W3FgRwAY4kPdNURVs
C0CX+T0/97jpZYaJpOjsI8pVwW0muiGXZ4dByyff8f1qflfsn14FjXfdprMqYcge
ohF7s2Ko2xNHwSAv5idnxKvTAEC/kWUIuBdV5ZVraToaK//IpoKoKxjp+OTS5gXF
cMpXlq1+h9gX1gqKBlUca99ioeRXTmFD0lcUdMR8g2wY/lfqgwK0lY/8NcL6Nn6J
vAn70H7mCwZ8/s7OFKF2h+uVfJ+a7b1CZTpS/0bpDdZNbnyXm2xG1KO0Yx5Es0Dh
BtOzIFmbsifK9PYl39dI7a2iJ489wN0Cj/EaN2ftsQTL4krq0JCS97g+Er9qlc/T
b3c+6QizhR42YRRvi1HYijUtQas26Ci+WC0nvgBuJ+Y7x4CymBZKGjAkybi2ed+C
oEvY3tXlkPaS5z0oHKdT0DF5QofFcYRgBk7JfXkAK4YC+0o8VuvsRazGlhOpbN4o
EOXEVzD7gXL7bOA8zTlnI6zZ+kKV5IanLgm+BYwITvRg4py/LDshhQBvBBWoiMBM
1oOwB8Frgmd8NySFe9bH8lGEu9MdiF8xpkpWXbvVFKUQVYfy4yaP4cn4rJCUGNt8
E06oMx07O86NyEwIr8iPALujxqltw4MsQLLEvm1WWQFjIG0pyvq3lc3wjTTgBUyV
7cdgx+35KOvovKpo7UXSJlDCIx3dtjuEc56Lgpuza0Lk2qNQdIAB9VDeBsh/oOI0
SI4yX1b5yNImMfRxq6/wXXPqCkv9RcAY99IDf3bniJVQT9uUKfB9fVH1LGbohnc1
oIPhszcbQFLxUfSjk3zC9ncdTUZNUZJvf3ItrmBk2T+OvGOgX3xSRslhNuWO0DIv
Z227F8t/r9GS5EholxZZqT3BObzoyjunksE8M1gTK+D/pGQwidmlZkhIae2fNmlZ
gxbeL9sxci4CgvA/vVlTI0QkxmNmvL3kEJ/4B3r7yCDU9OkFj4NekZMvov4ifgjb
sqMhGKGL0Ykm0p/8/ldlRItHAjeyr+0K7YR3dv2XQ+0L/6f/2cG8ra8FnBJSD+Zy
qRbuMj3UCHEoPhuCJvP3XUyde2U2A/SEkIho3Alisg75ZT8p0JWYrwGI/rArh08w
RGTtiuoa7LOLUKK8rYQGNauUrnEQ616boXhRBP9jLid78o+LAU1D/7J36dcaQ4ix
Q24l+aZ5VhoRAkdf+lqJNgx+PCSG4SB6PPUyz9wTZHE3BUp+bhE2R53RA/LWvLqF
R2IpyLxRSV5P8pfKE5OrecDiifNnAwhXVtFKETz7AxTzk6D/zRkj5ah6ABR0VsCb
yR9FuNIXiy3/hdCuVqJTV7vUI5ZWaXID4k6DGobySsLIsv0xVhnEZAnhjICQN7ZB
5VBXHqQnjuEWvP4dOUR+1wbgaOj+ay5ZWYiMSlQwiGQFcrrYocCk6pwte+Ly4yrC
AFoDuPrfj0040OUVAVc+ND7r0JfnKQJdaX/m/GBldzF/Z/W3kjX6/JwLCIOVcHgJ
2rCkSbcLcBgZ4Ux3pDrB0WeWeZOcSbkv8MVh4JuXRasWv8638JUd8HQVIpg5XT6Y
PV6QE/FYMU6dT7xV8prAkpz/1wHAhv47Dxn8nK8x+f9l3wwXGnHLsAjSA4ExBzxr
E6Rj+aGxlIzlZ8gteMAZVuicIdH1MDVaB1/VYHCvRm6+mMi85EPCxGRXgtUBlLp+
KY9zN6YBGTZNsAxbt2loJZrKPl1aEFcuJfpESA6VNXxpL+j5G/WeR24IDUNylFm6
Kfifx7JWBwDKgEHO6oKSY5STgCceNhhx6QpKuk8NmASsYsZQxS0PZ77efuSs4Zm6
lBSYSBKx6oRYATBX3eVkHFL/ukW6WGs88nD/tdhrQ1CdPZ7R2HeT4QQJNuMHajVL
GzdwtLLX2SR8E6m4BXsj7V8ExoAVUyngvS6jUn7N4Jn6VG0eiXNLNTK0qrCwpHrj
wEfD0hEeVIsNOgHC9IGHV7RK/Mfgp/OlepA8rjznhgyuHz0wOg+LA8dnHVJzSV5Y
mgglJN1xQPHk10Cqjn7+JqWSpf0OlQEJbTUGgV1SKlwycVZzHM2NlVmeqSkFJMA1
xnI9UvdE56RJFwZqT7504cqK2LxIBR8mRyK4a1h54lu9UIx1HAXmj1jqKH7es/ar
ET4krh/DhraMMdpp3xNrO9sa1E7XXktAFnjtkQvlA2dHhWSzy05mJichjCwgW1WA
EwO/scjllEuIs65qAkJMDw8yBVVOu3FTx9H3eYtpG5WdF0giNqkPryfPVLdTgxhM
9EktOiRnV9pHHpBMmCDf31q2SVH6MxdCJbGPpd20L3WuXP1887IgCw0m9iFJww+Y
TOvYhbNyg134Pru/ZppPP2CGB/BEn17/qYBOjsmNxNhBGsbTUwcjveqeu6WUuT/m
tbSIZGlknuOpxCDDSNoJRm1toIIvw8KC0SXWYgD0TUnReJzZy/CAS/kflgzgyleQ
JrPK9aebYZF3AjjWK4f4SfuWx3ULBWg6Tzzq3RYWARYY2QJyruDdry4vSGtgLTtj
LOCC0JECOyNtHXz/dwG9i4SPbdgX2DJYuKeACd4uWXnsBYzOdlqrnfk1vPxg+mwQ
LouKoQ6hIOEbLvvAKD2iPPS2VNicDs1AIg75DZGcOR7P75A+TaVFVhV2JiDlxF3S
81XxbcrS28hKj5OSnC5HPVAdoJg4pGigI7llJk4ZzE8ck/CJRGvXx0rv7De2mpqo
ld8WhbgfYMjygQ12JnZgaDj8nrU54idZ6RYTFukqFZCdv1Krxhp6INOI2wW7O/Ex
e4alkY8CtXQSYdPTqBMMYzWT4CcvnxRWDjMgKFwGW6r6mEH4DMzvOYlcU374Z0ge
O63SqACSZwyAyJt+iJd4dPClNQB2wVAuxuVyiyNTnCc6hDKwHi3TI/S5RRCXz9in
mvtCsJCQoUJsd6eXL498zHhnjzWL2ChrpQhnXQOq9YCZVXvYIsnw28OpQRR/XmXq
QWV7iA3Qs9bdfqt0HdaBu/gRAIObrpl73xTvnpm393W6P+AxuJI4UrhZDiKFijhp
N2AYUMH+Dp3LzpRDjf1SryWq5B0cA95sYDNTk9LJPav+G2ckQ7N5k6K+Jyhlz+Za
Gy33uMluozKNL6d3cxaPMlIRBZ8cR3r9LACcb9MJ51aKnhugE8IyvfXubhmUusC/
E0OafF2RTKnZRMDXiWuU8ijSBwLcqe945h8bX6354TdBtZpbM/zDAAgB/ZdtCD5V
k5IxEFLwKyW9mW1RULkac7lAXqkf9AZwzTiNn4mTi+reFaJVKAAqmElTjVO6w8Gg
l0Mt/q1pw6Aubn24sRg9KqmSr0vfI5xUoQcJHKReUC/V+jz+JuU+avHyiDVQkigu
bLopgllynGYsJKEgBkpEcQMHqpVcvvDQHsTInDXmI7GatGwhG8jgOS0r6QevDM2G
ScVIAxAT4hjw+NyJKglt2uJda0QeOmw8z36pc1Zon/X9O3nIvrXnBCopC+s5nEuS
LXHxS2oJwCHP9YLwcTI3doqVqey1ke8RQ/y1wa9ojgdCwXYyF7wpOrwPq+5EEhKc
AO8B8iB9tkxFJxOePQPq4gVBcqInq6trpim0ya9Kf5rcquXB2qCpStGY084Oh9uu
bZ3hvpMAAuM/+9ULvfaSAogWCdaZrmwE2fCnu0DitW1xqR4j+NNxFSjQFnZcCnzO
UKFFGl6gx/cMhxWA8zKX/3UuWtcU9sL4aaY2zJoMdiYXsTrJuZx74YZA4lSV4EyZ
15RjfLLIK3pDV5HY3mk7GIya3NfjHL04DdJdgGNEL1GSA9+3Vrd/01I1NlnYVByc
yPg+R5Uqg8P/+YHkFrU+FgjppahuHydC6ZLVBKIYJEFpm63sXdBe1unQyu98OyCp
qiRV9Tl6QH165y+PFhZ88ehWwP+gT3UnJJ0VuRU4TPFvizaQXCD/HLSMeqhqJw9t
veGqYv8L7HfEcoLaboeQmd+rMohu6+pjODQ8VdpvhDXgYrEbbraKTGYMggqhG7t5
BiNZOmJ/dhwhiS/kx6LfN9Ud+K0un/ivZPGk8Tu4I4DoDMUW/YuDIVMEpSlF31rt
vsDdqikT/y6+vh4Id6vsrtOwL1+R9rMgHCQiC1Hq6lr9GPht2oNV8YSeB0iyAcNw
KJT2mmN7rXaf5MSFDgT4pM5VofNmjOkCmj0ONGsQL9NFjTjGufuHpTnG6yS6mqnL
J1wzzykuGO7NWcDhir5BnLKrtB6aRFhktHUdqeayp6OSfmW+jvMs99/Y+5nhMi1b
Iz9DaS2qRnT+ePo1/NutK9N3185T0Ld2M626s4gnU0VkUFD8oA4xb77H6CXNZX9G
UNoZ2/KxlCwdIN1LwrIaaQGhqTXsIXQ9agY6I4DlWyI336+IXU3gV4Au5kFjmfHb
H4IygfZ3zTKhYiJd6b4wF67CF/T6VPoJ9nwM0FYsWIBPgYwCqSVii/JyYGhgABuT
tmfju1zaBIcqTYsHkXoF//HssS4ZMzcF+cZSwIHIivN9BAV/pA/gdYwL4mK4RatW
cDk0fzhz8N+lbQrc/Vd+DIbu/spqauIQOuMU0zggE8Ltsmq/I9hKIEuvPtmkXHaN
JWsP9QUPIyhirdumKTOweqyHpdr9TvaXJE/Xf8USgJMXp+22mN2Q/g7Exm05AxIX
Z7I1iAQQqYlLI4SphUbN9fn70FQODNTKoLfbRafjQMEyQLp5o/blNcVk3OcgysKf
sP8iDsrJGa2KOneFtk181BJGGlCiZ34COLNacGOTNtg2XDFWUU6XH4QSeXG/cgBz
0Gog+J7/TuOQ+5oHNhtrJ3a2FK8x/OsXU9HOG7XwaNTWAbQHH8bYwCnxxqWQBTaF
pw6cnRc9wRuSXgkfuAvnNWjVf2e4RQylDu9V7n/6pjEFGy2aszSoq9xFzgnXuYJA
klVLjUr/TfzCHPRqb/RnJrFynb4FR5ReJtHtr5R8BQ9drNa2WU4IhjbYN4QCErcH
K7vvB0b6Vs1B/iSq/TQXTkWeciKPgA2ZAXI39p99SrcrRh/NwNJHthud7uA0Pi0I
lZYSvlVrXXk4sJAjC2LibEckUcwwqGnbg4D2UFSzp8W0ou511yX40rffXczf5PhA
8A87+Hl9EwW4xJ3akOKAsJLVMXqv9sF2PAus4/T18KdCfY3EAO5YQ6RmUTO98i51
dEa0augXf4IscnRpnaMVe6kcP+yf1obWQR7FtbYRZINFvyYo6xnUz0xCVRJUxriR
s569fQZEEA+JM1qF35pV/uWO/nGCWdS/iCEKDuRHc/DbVE0CBZKgRP8QZu2x7o0q
9xC5DAoOhWHpuCqcWZYpTJTrzUPSbwTkMrdBb6AxU0NPxZOnnn0UUJaw3ihsMU3N
CxxXPj9keBuC/zCvF+PlnndqbLZsDLgnmkI9oTA3UIQ5dmVGyNrjpUUU73ghQ4sh
/5xCeufGgVK6Rs4tCRF1iPG3ASVwkKkEipDZW3hTSIswWyPAFh1TqVoXq55Z+/2j
N53Lf/NYkCEGRJpxtaeJEE+OoNtsiVnFvDZWznIRiuYOL/JIBYkaDebNWrWM/NKS
ySn68oDDqrdbm/ChZE8izIqgwn/hlaC0ItSXODER6gGItLqwutjXikU5c710slYA
edKaZAKtDYm+/ItHYgRtdIkFjRFH4AZshK6HYivK1NNKmghMx6kK736mxpU8ATRU
Za4HfXHF4wkD8doMcdGuiYYA25SpNQWF2u8rlKgeLy/NyUG/zhTojBY6YgnkYQxk
vlrs1i1js8pE0ZOHZIWZb3AUtxfWdNmWP1paUJM8cFU3dnZXlwn0nMrBEZZcz4di
ufgUoaS6H1targi5U8IO0IeFZik+qjoxf2mVaxdikKjzpa/gnirscNj2AXbLdwqw
9cTFJGrWNnOhBnbiWxKPR3vomR1YW2V0xbCotruBwOfkTglWzrEfauFCAbW7RZy0
mb6GnVq31OHTC43TfiMs8NgO9Hx3Nm4jSf4F+oHkbXh5J2+0HpnqhEXUwQ0G8JfV
lFTgb0tPv/Qipyi0uMRqVBzMxKziFoEXCzJEQofkcVZFRoGHCkZ+u4x2P1Iw9xgn
ZxiHk6Alu9UHqThrmAbpehOjStlP7y4XABVsb31jYDrhu9UezyWKRH8OqiF/beSF
DuHjN3Oo6ybqSqbLFf1L6nCnolX4B6FYheFnF7hoLXasUwF7oIhnex5V8W4/xa9g
NDtSDhb61YnkHxrl7rKR2ilGFPuW9qdIQx+CCQLY99gW1y0R98Nf3D58fYBdLA1Z
vZFOztWj8E/cPJtT2IgrLW3xlY+SsSb/KB2lXT36Pm4Z2AJswyazeGIbeMrHc1cv
hR045GnG9q0tva1+JeNPZFDfZRx0l/okyUErsullpjQ8CQeTy2wTsROdGJcgJ91M
8bzqneVr7KK8deJ57WVrn2PA2napaJBIKbjPIEv42haioJTxdLm3pNZMnZZQS2Gd
sJ8cdH8A8xKT57d8qxDsR/vlX3HsGBUWoG0Buhr9Z9NdYAhDepZj8OLH0kV/DAON
q5JzUThfJGra10x4ignv2xGtk5xGVf2MRsYpMz8yrkFyTXcm8o90gcWKGJGhlRpP
ulOUXd4mgWq2dHVkPu1iXXRzEUnBBa0s+DHQOOx+j5xrYqkeqCyPKLVM7kO9lq1X
lgARVeaVVtHdm+PCyocfOnVYt/iLuSLmEuTInkxNdnko2xqf868ecfovUvLJXC1V
KHUAzwU4o4cB+gQ3BQEz4xisENWiZxu8lFeLc0IS4T6RK6KeKMCzFrZzdG1Z3zQ3
q7nWriCQ1Jug73U56Xn9dikHxS4euhZuLx9RCXmDHkC/HBBf/QBwlUUrMWLxKjAg
UimqMaKIU8wpl3Ms1vfsSPNOzl5iOk5Ew9Wr7kFgK9eT1IV5t1Au9brXBWyVvB9C
zknBF9tWuE9nvG6pFHj2KEBm1ICdYl2BY5IdVaheHcUbXLqYQm6HQmai1I1qsxj2
t7ZKu2AgecbSIKx0hSZx3ahsZIFSMcifRrv8gMopJ30k4kWcZ6JvPZHNlvXtfo5t
vLTPi54gX/FFmcSo0N0JoXIW9aEIbesBAp0itl3cjtxiwDLryNmd2bT52AVJ/hKR
U34VxouGDeuMC3u3y4dM3rlfCFe7E/kJULfVUe5PpxfEALYBeQCn73WlVmcSfa9h
y1FM+9gudkHevv5akzDiRUyCCscsGu1tIWQ8i4qS/9MlyS6jROe88GqyNjf1IDFz
b3+TjfL/v3xpYvd68fFDHxH3Q/FTDWZpztIYC66y8Ka/vrR+CAYXgx3wJx5zP/rn
JW/zppOV25mdaTYTUqzB6vXxJLB9MU/PfUKjDC7wp/xJTZ366aqK7Mskb/o64RNF
`protect END_PROTECTED
