`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UY8DAD/x1/IJaUrWtYRlcxmhS+huro82sBcUy3DiCyJgAoq7KMOvyf9/QZi0nhu/
9iAcAwAgiLTjHBzl9igR6t0w81Y6QEfCCDP0Ykl7r4zLA3LQ5HuS+/ai40x5Ljcx
erB4OIKhx4SpN2R6BWl2vBFg1KS7I/lzSqaGl5Wu+67c4NRQsEdUJUvh0HLpB4G7
GN/qScP8u/T8GNz9bO8+OmaU1AGIK549nfLhTLA1z/zsXJNaOX/LWNgbZxgurNvQ
zAUzZNi9iPV4tGLG8n+B9rdmvQTbP3kcJCNL+5QYf0Lxk3HPtLV7XW7ZZHsLc5kP
4bZhAUqiK1aJw93YztFA5UrmAPGEoeOzppCz27YZAgDX96S0B9bnjdQ3HBEKgsd2
uXUjDoTWnoASXEWlqk8kFPM4yCqTBn0Rx+w6BDNyGAukXjVjQ2PXDnpa6OWNU/SK
WFKfEN1K92Swi0OGl7VvB6v9hlc27Gwe9+DZ8H8NtbI=
`protect END_PROTECTED
