`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4mYKhgLuK2bV5hbRn9BDB9pAz8I9r1h382H9CpZ5ZQdciU3OP3+iXohm3ECi4aC
swbqXlPfw7E6aNGUv6mOH9lqJqjmPqZ9lMta7piusDrQPczObxQqPWnOEwn/PhGc
cdBo9w3nw6L8Fd0srp1HNZCvJWvliuQZcHf/mHHkY+MqdoGuBXvbksXCk75kxdEJ
yrTlqfUW0jvl5UenOu9dIesFQ+DeAn8NWTQI5F+7OYUiBFVPtrgd3sjnl3uBKehV
tMddpJgegXDJDSz7rRyS6j800r3pOTac4fK84sU91gBtutxqy9Ud/we7VinO0HaE
+j5EsGYWm7AmIZZf4GY4o5KWWR3WZo0sEjHcR0eK/NTDDMhSk+yj93S+0GaiEUip
M0Hi+weqxDmetgPEujCJqxPO7EA9YcW+jYCXzEcl3jui6NLVzaWVze8MiqhfwtSb
dGhvDgGZ8xHGD7Q/2Gm7gUBijkl8idf9p++tckbti+DRq+FabHE66UytkZYvlYzl
WLdHEJyrs8Z7TnPCX4sMqTV+ySlOoT2tDO1dbB//dkoLSthGMMi7HVVBGIXEuyNH
6xhlTPot1UMc79AQRhZXpGGD0Cm5XCCwuiw1MZY0mKLdyQnn1mTpTJ5BV5CaUnIQ
JJTFNFQXzCgw+O+AGHWwWnFMmHQ5yKMa7CHxcDYCAh9FADj9oYs8RZnEdZhyMrB2
NCLZ6dWf94zcuFKr4NqcqgRg458YCT8rr9wQz28xdo8CJkW3YrxeaNADFNmtta/g
RwBQ0rKUbZDradR9zjsIhw==
`protect END_PROTECTED
