`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPKdi2DvKo/XKhHiLM4vEZ5n6c9c/NkbJsSBCu8U8/oxawJXpefcWzDQ5Oy7gj/t
8uHVVEQmoprS9w25PXaZlxi9MCRAYj0/tWKWt71Aucymd6dvhWVwMqPixBOVBSoJ
bMFxj5xLGdlOescHe2QurTmT1Ey3Znaig5FCaIoYEL0=
`protect END_PROTECTED
