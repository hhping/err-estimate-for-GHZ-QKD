`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ErnsyS8TVYK5bzPZ+uQyJkhHEnqZaROEJeiNhOAWrfIdbuWTwc+rO9DS3BSOgqa
m4ZasH+MxAAidkUdfNyEFjbeu9eOxzFYKqwtN7qIx/oG4+7x//ZOPxN8oVLEVBLp
AuTU/8Dovc+8u0nwzoVDZaaKhOEZHT8aPEspqE5dq6176JV9YxF6o9z3DtZ45GCL
8pnMLcR7veO9lx4c6zoGtq0paXvI1njI79zk4Ox3kd6vTTd6cksncxMzDrLgcd3L
AaD89huGtnNQ3MZWIY97vMXVlLzI7g9P335XOIBfUr+wCbvoxHeaY2ojbHo5c5h7
p9PXv0CLa6F+GnCJnki4sG1XE+muWLjyxsgOSDRrgFFDyBHTu3ePGWSYZroHQFjI
fixP0qYttthXgNpxSEoCnfIvXe2mSyunS3DawZDFNueGmEA4/4FUxEo6zGNsgnd+
M/43ecxLCL4jigfHzf1ahjqK2P3L+u+q2fM6OtfGyZyKyJYXNyVG0MNx4ekjNy7n
uLejmGn+r/gFChQKY9m+k6DstdTIagBmlwSfQWBsZTRzngYrLlTVHn2ed00tEsMS
Q44QovyhWDC0pY4DGfARrvYBl8N9Cy9eRH2x+pN8OpDGsnFsYt/2Oj832rTLjgFB
3IX2viaMs69xCWJH2y2T017rNQRc4aWwhahrWtfKGnKDFLG1C6BvrMuzgdzNwO7r
xOqfk4uJ7/+kZ8Ci1MTmDG57qjnPFL9KRMbspd3iRaMuhnK85S+sWx7l42UkGQ6n
nrY56voABdVdxVIkYkeCvtzM3rnBXKdfnKwx5n2BcrsxCF79UVJYbcKtA7MxtNVx
1K4tiuCeCdSeH+FIw0QqRcI+n89hRN2ri24uTZfVP1wdvv+gEQVzMfcaszePxjwK
luyr5hxcbhkfqKx/vPoPRDvIiBl4eLbtYX+VVzlqgjfGQJHKkYDgQaTSniuwK5IP
cTSKvtfe4mYzpIewsPGpMvHYSXx8kKQKut0JX2KVgPXMSbQBB9HfVNrOxvHB/tFx
WAHVBmbjkfMRCzHJXFcNxlQzNPa3Yq7XKj/tYxQpD3MhIczcTqCVu8CiZKPPhysq
/pgTgV6q8IKVx+TFWhWpX+NBJH8GECz+MzLInd6jur+Nr5H/WWX/kiMuoL1zaVO3
5xfdF1Sq/9rJAgt5YHqubMzqXDCGfsogicJ+avzsWx7yVm6WRuo+E28yOLmfZiKT
`protect END_PROTECTED
