`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONA3MNRCixUtMjAR2lkOSowaDnj+eKbTjWrpyBKBmEsIwDT1ZmbpB3BP8/SZdz+6
wBZqubLKzxylKXLz7Jy7SDUKTPdZd+p8k3F4/TJQoEnfWGfVOO2l8Ul8h4evURRR
QLPU/MJwwvhvYpv9V9HkR7DAdVAA4U1/l1xE0WFutOlI/4eqfuy6fn2Az1oaV/dK
qXjC1bVUqOx2F2Ma4GNYCQuGX3qbQCzh7azkUodtqIiPT6jjg9V6KEMgtDOaYxKo
hTCrckXB7H9x9YFvB3x87zxy0+0kP8ccmxNe+KNRkqdcmS8huxp/jMEyuMscuELc
LxjlOqShc81CUDgJfQ5UqGBqOgNFTVnWpkYe9n4C6xc3Pfn43mo75yTbw4E146Br
syy0twCdzFAkYy0Rjc4D3ysuL9yA146nNq3U3heVrfvB4n38EAGfVeC2XOf7ANQZ
vpG9FUKmoILKEk5ZF3OglMieQDpmDLrixD7/HvfydWDtwx970MwswPuHCVAREoct
4/hBdy3R14vFiDa/lMrD8nkaOVVqpMffHpOSZIBMQ6dLEXnqtgY0xbn3xg+Vbf/y
fYr5SxkFDeegy3iF9debTeVffdJlzOgde9OMH0MM4NkypixRw54UNSB4RGXPSzzl
514+MuhmRbmTg4Lkx/qMxwfH+gBFVetN/ipznBfQM2W/Xft8YhFdCstDiFrwB+jq
w7wlkr7VETdUqaip51By0wuBhkDNoE4EofEKyacUKkFdPmH7LCKEg294EBYxqnq7
N6gzkojKp20qRSi3LyZB6Tu+3xz1JW0aYCYRyHqlajs3ifwLF7hJDHqAoGe7FXoh
kX8pnkqG+L+0gkskYgAKKQxwoeGYGvrfkQeQv7PYTIwDSwvtMUzdsy96Sq/2nrcv
0lSIjnptTRTYuWXZsUdtQ4eepPiqYJwf4RHgIWMYm+dE6MxS3ByrtQg7f0LCUrod
R84JRtok5nDHRMp04+NRAHCP9N8XGlz77+qyiAFNXh6FrbzG4gnxAC+GjOcbwacX
ZzyXIwZO5FMUsL++AiM77P9ZvU3INkcGV8WH2oHdR7I=
`protect END_PROTECTED
