`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGjfC5coi8TNMNvpA9KEmX8CJVMV5orZLkcXj9VP9LorRxTlGhoRvyg8tA0oUUYc
5oUZ1RCYvp/X4mZI+0qaWKxnAC4/Pw7E9oaguD2luVtHc9WfSu5rsiqJv/dLgAdT
XZvVlMp+gQ+wLe56Yn2bxI2RZrdYINUS5MTk7iYQMHd04PtWyLYqV5xxi+NVHWbB
qgf7UmvpJfB5ZojvfB/G6DQVzbHAbzvdgoqu5zElm/+HFOVXTpApLtweLu0GHufd
IqcXGOCgloa76giMKRWEVTam5ZBX9WYnMW2wHxOXchampTG1oZ1czEEEY5NWRsOr
4YPQaG5hGTzY1DyrUZ38vD+UUNJTFWXPGpvRKJf07glaRSkTKAOFc2d6MaYUMbpB
waFOhpGdkB8ak7LyvHtSADLlGX6WfS8wYfgsNv2TICuF9PdgHIjD7etk+NVm1PJV
YjSnII3QQY49XorYQtddWyfO3rMYhD14NWCEm9VW+Mc/sTrIhmLuQ1WFugZr2Xvk
o4BQ6uOzm1DMi9SO5CNvqABzx6as22usm1L72waOmQeHTvdsHqtmGqEv0am3zv4y
ewNXin2UPpSdydj9dxBC3UuPBsKcw1MktqTMagmwDtlMf53IGc2vQnMn/SvwbyP6
WWoXUWVIQl8jS5Y04j7XzDcEeEicenYUDLSkHGs3HMX2f5EzqTxxI6p850APjKm9
bOsNVb1Dx/FBhwFYEi8YuNFdYTpV+MAqB19b9nq7B8tLidIs5cuNUyNWaDfivMTx
czzqFc/icnDtsqI1q3XaXdqnPdH8LjiWNXAQRJXePTgnzoGGrE/UqXe6Y12nuZ9/
LpXyktR0ALjIAAGtI+3JgUCP6U0/wBO5TjJXAs45wufmuD5h5tkx/WGOiFcVeSuu
Kdl5KJ0tuuuiBoUTLusmTpTqoeRgWrCe2F6EEvvyBxE5cMLgG5PCk38+3YfJ9drr
dyapolq7VRGJOuEopNEw0wSjJ2OVnjED8er/C8VNbAXG/56og4TiA4feqAFHeKFv
izGmgPkFfwXSVtgozIlthnkgxVcae4GEcDmkAjN40sAVGBTrKfT7MyKvngObOJmM
lOjVwLgoqt+ZYDjzLUtCmRd16+70bBvvfr8xMSSVxs/P/FIuUz1oIRTJUHv1UkCm
UuG53Imt19dJQmGsqQeHsIpgOgeU7y5np8fz4zUziIIwSjPva0Y9Cwkfiwp/3vht
BiUokud7CpOY0hAy/BEqzE0BKFz+uachlNJ/P9BQeK5tHIHN0sqUFAsE9nf/50u9
Nl4NruPlCOqfrUiUr1Wip6Rwm5/9exrrRyUB8mCUJiXMbFtqTzGL73Hw8Q9OU3zw
iU/7/DYE2f/BbkdEyyYHsqMY8wMG6a39zS690X4kM1PP9VWf8IX+yTeD6uhAd1MZ
FChvMIcWQA48FhTWrGWzq8/X/AUKO4xUn9EJn+qVIW2RFYaia3IQacmsbhtjPH4q
bLE+cK9qXcA8flUziad5v68rhUM3ddgkiPVYuxxSuyOtQVvEWbtTwNnP7meUTj4v
jVMgd1SK3bMjKQznkVzi6sgGdfpp/qgKWXAPu/Pv28R4G875V1VBcGaEFsaZ7fWc
R3N2puczcBJqtJB/3f6fpCkrhh25gJUmHe7Xgbb43img92XRMLXWzSGbH6hgLFIy
0NT/ZXPJaaLoFvM7ss5qeQGhMn+qT6Lg40GcicGnE93p6u41gs4QSjR2AQnWxjM3
FcqNUoNOGCSTqLOv1PornmOrEwYK68B6o6978j/PN8/rLPvCUPcWqHEq8bsiZBPy
tml0lhZx3ZtZZBboyOXxpvkCbENPxqyAtQ1ISmPWqbzc5ZwkmeT/tmgkaZzoG9n9
a5Djb4M/QKzkRisPxrNIbNtX8c439UV59QaGN2/2cH5KhlRGE7ZGhCeoNwHRY+2f
su31oWrTjNTmWpbAXMtaTYR2FgLHaezlFZYIzWcxDf7IajXi8fpgaYOlTy0yvdjb
VRhVvTAgxA0CYkkchG10dbEmw4ccDdS7y+jI2cE9grZRskfaWUvyVKFzez0L6OsS
h5bECmJE8YSlsrMKmj46EC+nypiSnco0WTC3fWN5M/U7WSKScFbGFC1T/09p4npZ
nTlvm/8OFrL+Wd6z6o91xjn6i63n+X884aud+DYW6t0jkqh29Ouix3aJqxxRdxUN
iFa/Lv/yBxv/K5vpRl09cplROTSwrSlzVJwrNXW8sZbsketi1qAqL2gJ53n6Q5tA
CB3nTYIgrgV0Z3R1gLb6BJAMHTQvxq3gmYo/XwEPHWYPFxNq2xd14TVON+nVkj/m
iZah9hU58NQjX9HAk84EiBdthe8s/gaseEYiHNYuEUlb5Sz4lDCJwgVyJs0wGsPR
o1DW9+Bjlx5y9Dw1pfB5C9SqqMMc513wBe7THt8BPtCf6JC9N2FfD7bADVJg9DxO
ExxaFaE29Pr2yJKSNJRGPW628OGgAlzB1WG21K8BdD4aKmYBLgKWmn282kKWcoo3
yePDl9xituTaxeCjxCF2jQI+YIuJIOpCxi+HXu7/mcUbrFrDBkXLBhmtjQlXJaKO
qwz3qkAEVthw+hzLpSw6QxdMHviUpdY14y6+mm2n3Ur+n9r/8MJcIyDU1gT2JOPY
aqlnrzDDlqU18Ykz10/YMSBmIMctIHbBWZUkzyofIoM8BSpu/Hx6aDrqf1dROOaM
7YO/uev5e7ZRi2rrW7XrQQ4bGGW/mtsVzCSp8veEw6EylLwUPal/256P2rAkoc4K
vcAINQYwkKo3spUR2brx61fFU0sL6DK4+M9fms3BFvDXp8YR1fTrfslZtWm2dfR0
pVggC/N7MWneGoglej3LjccGsGRaFwA7ZUGeAvpVd0YBG+0XBZ225SSu9nyg3F1g
+h+r9c5SQXC1KxRk86MfHafVa21fGYw1Lvi2KlWQ3uYtY3NNZSph8ye8JX6ouZeN
Lu2ovwrOr7Ch324LQykgcUO1x+1slsHv4hfxPNMzHCQ/Uy5c/oLzSUzgYdFc6U0K
sahlRAFsJw3IpF1u8ZIAXeOFhrInOPY/mAvaG9V6Wb6ibhAwKYFUcMo5ml2oQ7Ui
7xuvz2YOmH80JrCKptkX8FDhJ5gGJtPB4oGEEaoCfvZFteM1o6sKYuqEkq2fM8pF
buF3ramAulWPhxi9BPdXa9lQmReHUw6Q11MslyOnMJg8kY5lJAy4EEPKUDmY4wgR
OdE0OLbKQYQdqDuglPKJrlbMRPCJAeGmWGwnHz3NDOsakEB8ninZ5HqphMiwhzpr
v1aZSe2DqwOCnF4AdjC7DYRsEU1K19Sk3HQt8OvJj90vR3Dllz/vnc+wIF298/Nl
FbrS1O5+IM3iFA6/mRKSLeIwV0U7zRE5xPXL7TpcmXhaSs2PC/PXAXqp78kLWauI
4DxUdpEiGnA7mjhlzuIdus8OI4EUK60Z0BnPXdFvN4zXvJp9PFpg2K+sqsOGkvPT
RxBwkwtS28saweL/ZlF6g7d6AGtLkkN1Vp+Uxvb8eAW3RlMtmmEl9AKefViNxDoZ
tHZQ+VqzHzlDiOcTGxPI5ppf903Pr0fX0lK81x8DiEDivwttKsnqnIDOTwm+LPXY
yoJzlrbJbjbno7pnY+xlPik4n+DVClJJJB+x9tBej32082n8xXCGmqxuTyotwgpx
bnazxMeSBvOZ4fUFFGx/iUjGmYWbqjs33WvAhsrNwTCo2ERUXewJWJSs4NtFGTVb
TMWSWmOv1jRECrbPqdcCJilOZ95iRSe/r+Z9a+HNk6CkQdfoY4woR0UndV5pNlw/
6Fhqn7GXk5HwysMJezRv9a7lCDsTgMM++LobwdYuNG4G4wqWBWHNPwbxMHEwoGTo
Yhs5SA4HVfJHOAOCGCSUC2yZHywPN+dhKKwumwFFkA0KRHJ3a2kG4zCA0w25W9QA
R9owPIfjyKmRNm3LBTZiOJgxo6x5vea2rfjtPZvZ6ncssqUCf2nIXGyDNlFhYPrO
OBY6mb0gLtUNemioytfLP60tUx8GCglQTqwT1jcGQAq+3QGO/zwzcak642P/5RA6
6QhHWd1a1s4aYPrF8ESEfw8Ok/4/S+1qY+sNjOYiI41shYU3/aMOLZr6rHiC0fqd
Ta0ozdql2TaWy8Ry+hNm6/GOXei2Z2NKSBzTs281wMkSpj6/duNI9R6TZS+TABQK
4UzDkUEormm5kXoqF/6UniLLxi2kfWv/yfnvzCc51b01cizCD8M2DJCqBzOIv8P+
ppNd6Uz1JoyOcMdPup5W+HY+pY/55rzcf4TbT7VEx6oDUz2jANekMg9n4m082xLQ
TBXcNCWiPy9PGqopcn3ZIx89nWuor6erqI9FyPL3L4IHshlsvyNYWrTizt2CZ1hK
9ouieMqB0FR/o0mjMU5f+y0rPnE52npbRIB1h5jqGbBc70Vqbcog4+JXees7FlZ4
zSIgGrI0PRwGEaUZasEKT7Bt2xoP6OmUO8qk1GSP2Ed9/TohUTjo1r9Ya1AvNHcR
Ia/ZaCfeyVzHcG5PKyHcGQ==
`protect END_PROTECTED
