`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpBmBfqMpL8TBWmlVimRy8v981CAsIzYpz3hG0cEDozbzYyGBT3B0lBdq8se5ATz
vYt5xvicNdpVQ4K7jsisfB/8BVSiR/WZJglK38+1pS1Tj5RqNIndoXFwuobEfBCa
/W+41KGEtScCzovUe4kxWRurYJJUaP/gC0YVR75v0G3ZcWs/sBfL7fUSZQq5W5rm
7CCNJU3tn6DC1160pGmRszkVAnR1vdGcNVdfRZd+PSmEoAj4fzCAx1r8zizIgmtb
V+XqJaHO8i+ti8f51ZFYHSGihsvyUQclWf3JGH0nzO8BiVIX6GoTHtbQnsae3wDg
R63av1REEJnufV/aTWz/FEW3N8mk6vB585u/Kj9Dw84HZltRHDgOmiDEUTKx4G8k
fr0dVtanxsZgnuuh6gkIYJkPPmMQWKwlh8wugRVtgiO1i/ec+4EmlnxzrsyxYPhK
LaqV0XZ3GzIW/XAmsAZkDsGeCh/gSMszGo34iDhKId0MWlsVudqHDnZGp6k7dX9o
ZPXeXqhIsm9bxNQB8o0yBpM17wk3AfULVgGJPT0JKSQXTVULykGSg3Q9qMSKTPnt
kLFm2BF5duM9TRixsnpC61J+5LHneNoVz20T6COYBc9JB50WpmOLWPoE7Fg1KqPR
8wyhS6c82NnNQyKMragJn0R4/OFAnGxiO+TveneERtsEksw8SA6hFWGD6JPFdyfm
aQIUQaJGDE4CSFJo+N49MzauII+UuwF11NLL2RFA++P842HcUG9nlvFIAdzpPOgX
wGjNyBe9TXxuTBUs4/crZMJSLvaMHGc8vO9OR4ObVq8uSHLqE7SBCxyTGSQs8HKT
4JMhizumkdE/6a3QJvXvhqKDK5qd4n7a0k8eObwvCCNv932QR+4/0tOo/FrbJdMF
5ycu2+nEaZbjzut/RRduUvUFkT09UKBjdov/HZMGsYZFOPGhSl07e/hmY6nVMEVY
sA+WcmTJMEcz31ZAVfQwFAc+10Y+v5qq0lqxBBhi5PzKLtjTKCSfG33VonSE/gv+
RZdHjo+JcK1dBws9iw3HHIl7GwTO1HQX6hu5BS2BbZpJste4u9aSI+wVSh0dV3bd
WPQ+GaZKWNbIgE6CN33b93xUOCD+NAx1rAaWOHTdzHLzbeKIquFOG2DCO5M/AQZu
RUI+A/3QThphr+HTgINPnxpO6/qeG3tU0KyDfD2me6sZfHI9zBIsjqPtSCq+T5NC
dUOZ26F98XHf70NQxbPNkqnH8zzA2hPFZzcpLZorVDz4n0uxf3qIN9j0Qy+1zhZA
JpOGYnUbc8z5rrMAug79pxQlIxwQ9GiCXc5Y1echg798siSYQhKwAWRKY4Bttp2e
TVLalPIniZR9+c78FdJ5jsR81kGuQ7vZ4P2waMfozpxiLR4V76oXMcoZiJevs8v9
Wm4TWpvtoB7qsQ1rTkjwWA8KV7wQZxBxh72HFBe708L/00X+N+IpJ1Rlg2tbuB3/
ZVbAXI4ofPEVgnJLdQv/S+wclVNz29Tc5ANM7tlomLLYI0AVig9PKCVzQdXKzU1q
2+2iUpbVB39UFLhXOZKTeKB9rQj26as2rTGLjAAQ1z5rEUO36fAbWeH0fZUlOQ/j
18bvGIVUpcuX00UU9M6erSqsTeiP9p1AYRrIQhXaa6lLgkkY0XixxBWwYeGPQuCL
4GZwcmeJfBREXdywpBFLgWb4WEME9WDsW3RuR0UkfvzK7uNqFQSPJtrFAl/0vx5u
AANbImE40YHRZXEDmC3ZCuH8bBgf7U6rdYhr3nElU+e1Kaf9n8yOfuQyyri4os+G
LNuwTTiSBsbKCSwhjhx0vvsOE+d0Su3Flud2/4C3sGTx7V55Q2jMt8M/7MrQXbWC
wTFuKUeGnLC6okYSEAlmOiyr2T6wWlvpdCfeYw9M30iHL5HCzX8o1o0Mtq5zmZkI
D9/Um/avYqb46kL8vBB03Jv516/o2jOy3FzfIo1shzAvNyEYZWYE/fsN/4ZrXwaR
GPNUlF9i6p9Y9QlA57n6lDcVslbXnTsO2oV0ZH2Ll6Xic/y9v1Qn+S+ibrCR66Pi
9QfCN9BBBlwOsCcnp+SjsR77YuCzmSm7ZOFLuraIOZSS4mt5XeFH+LjB1YT8Zw0C
Zh+1+lYCWYIdCfe4i0mXVUwnPagpk12wZE9sQjH/9ISgvNEgt8g0S/Ii+DALbBh3
RKjbMJEKavxRSZMtemy8+U6CccPnoYzmi/XRebOnyiVewNsGS1oaygvCvoiRSgrT
B6oFRYvD87ShrMSoRzj/9qZBb5H9zi//hXOp4WSdymtVPgsV9V3i85KU2t52L2g6
38YhJ5oqNFaPNmNKu0kUlrJPt008OTU79ygoL8a54BjpahzSUyvtKDKyGji9Kwd4
8q4iZW+QeWvihWBnsNIk0AbKnLZ/OtwbVm7yO+P9lO2HQXtZ7l1W8EuVPwjaQvwn
qM4xeCcxhr6Vc6hqMQS4A0lADnx9w9Nrf2YPsKhAgZ4bscgB2Cdcrzsd9JdVqyIt
q7ffXOOETXFGpeFas8MGfqc9uPYBnZ1ziejhFFSIpkhqmEve8+Q9Q4qvsy2K2owR
bwCnazkQNofuYk498ZVO5qerCzad1XX4Z+xUYdf9X6GOXAvqe4ch1VQZ+fSQdhij
SVw3YWh/ODQFwCIvFjTXTc/2A1L+t1WsP9uACJ2CF7rx15g8pPkNFxobXbkDqqXe
vhmgBJ8Y61wHZWiXr+tjiO6YjIbSi1C3VCUFYLpcfcuJs8sCye2hnE7Q7kTwY9qs
zl2ZXLM5Z50HUHIgeCWDWJi9mK+GnztqMk1/5ngKRITpklf3n3SkMmT1tFLMf/dF
4H1SiGr55IxmiH/HvuUWxIddqIEJVIhzBw4jrdx6nlODgCdF9aCRISUFEmk+8FcK
tjPVjeRJeTXfS66IkWOFETw6cXxT9loAv8PSA8hBHiOeAAdovpK2559KYlGNY0mj
KiiUBg4FXjvWWdUx8tAJadxASZR3xHd1/fuYqHB7Oi30JHh9YmwqAEcj9MEv6rH8
OKApePgpFQAxyIF/6rUPgEcSx0irRTdwERcOAlXqtxnS2OVQgORs8NFkNaQ1zVGH
GC1WtKzaz9dKxtH5a3+VmfvnJWaIVltcQW9ZUjuk71pzTT59WfUCGMeDxglu5/an
Bbyx9uZix6QUj+ArzLkQIpCbNmJTgsN06GX/BYRYBo4OZE0IZsgAA5MFQNTJYUv+
Rcat762eYOrPhpdqAR8IFpRzEjqPBmaFQQ/18P8rAMYpNNp6DTtf8VBEFTCUCJcu
D2GOPev+6aKlnWCo5vU665t2z9V6DVRbt2JeAANJoaAm6Fx0c5Zvku4bGmuyaBPI
ySqw6jVnuNdO5mQv3V9JKOt5JpMN4d7CfvFTNZLz9W6HMezDiprncaAOD1tr6oCr
FJLrfBZ1ubv3bS+QIP+nwNmoyoEjeLhKJ0vkZ5RtugLnqGdVUL/SzERqIdeOJ6OP
VjrroVkQVtRmgnh81763s+QqIsKgFWaa09G2D6fWKDyGS+6UO37kKaG4VPMmxbnq
xOK5xssdc9CX7IJ6FKRB8X3L9A1YLN5nHmx5DWU/z/BBQdOv6nul10CHllHQHNik
AXLYVAAyOtip6za19GFovwUPoz+PgXJ/i9SmLuT6q0OY/5BKsdI/VSQzAMvB7O2G
yLd7fZeqZOz55gVliO2qd5GHhd6IOkF/c94FiPCnnU4mXfMdyqFJvzzI0ZZFBTTN
OAtRCPoFxJUp91ezGttwUjSCp9fmE4Tn7hQxcTeW+HLtfiOk4Iub/Kj9FPTsxOvv
GgCCGlm/i/4GeSexPRRdnpe/eyd9vbI5wD30aA5jzx5Da2AXJu/Q4tWwQjpuPl3u
hAvtqoDgBrCNwDpPD60eto98wur7x3LS5eBOd5jnk9HJ5vD8fSYUZ5TwYetQhBYe
LBPE6q64OyJi03HdR4JN3HoQvEkfhRysESbZ711YRh2edBDV4QGILdT0heFpfaqR
KbH1eclLGKoBhR2/85Pth5W/VVDdZIbBbh+iiNSBpEyxwcSYKyW/5rsGzm0GtziG
Hj2SmQSq/Hb3JHfHc8onzkiH3NNMXXDvkipENaa2zvyUwa4sJweBAGs1UhbTa+WZ
`protect END_PROTECTED
