`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JY0rUCIKwto6s2oT9/H6XYKq0dy6WITNHa1b+HizEgj5u41+D7VkjxOEPjepypUX
0gIzUNgQxD3tq7loY3W3lWHjBL8SqAEWCzqrTGA8PxBnt9nVu20QhotNWCmnoGfP
pyFuzLq9O6HXCXU36GMQN1oIsnOGND5m1pkaluIfV+E9QSVXMc9Pf2StebdtklLH
i82p0+gHj26gi5SSD3MtHkx9VE9NzS2JG/dq2/XPyrZfrs/XYN8zdIUL8+aMtBdF
1TrJrn+Xlu50GKGHKAJRK7/WJAWR01bGtLXmKSvIYsbPkZwh9ZnAdqUnqQytUmDi
nF6hcyiCiXRbu09WGv3r/plS2Whobl+lEfQFdvdixr+ZUppxXhZrJn3blzfkNiXQ
nJsfD1JKaEDIbOmB5kLwFk8vP3BI7ox/EBH/TZQWlGkG5iXs8XeqlwAE5sB3PLCJ
B9BLg+6K0Lvhqomk2ZnsBA4wnSOjReJ6L6yIu0qgBIhGZ1XhShAG0I0lrsF3M03F
AW3lFlE2FfC7hnoZBnNXHcIh29KseuEoFEp4+ux1GKIeOyJPXzNRwsnodeoK6AaE
55pAzU1laUimweIAbDadfRr+6ubGEjbfobsejNCqIoOLT5OLpIfmuJPfGiVikcsT
pVHHABPNya4c9n6wGMbOoQ==
`protect END_PROTECTED
