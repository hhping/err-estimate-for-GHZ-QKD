`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojE8KqtZFHoTxmr5EbOGXgykM5e5h5ZNDZ6Z5lYNU6RI6ydHv8AcIIHTmT+hSXND
X5XnBkZftLaqs3TBfYuZSyWtDDzuxHUCTBL+BXb0Uz5JOxNZqNuxaY5YuigxNh+s
rM3aUEW6HRQ0C99HIrGrD5E1dqTlxVlDxVJ4MCUcnWNbA6Ze017vV2RfjmrZazFc
4yVL5VnIBdwi8j951Ca/Ny6N6pInGML6ZwGJ/AwutEq3JxpEQhH7z6Wl5+r1d2OS
or4KFqMw7/SC9QJ/UH829ZWDRQwMTbylrnvCELIgKySF6+Cd4DCIwjop3QLMEX8j
/rW74PayfvgjDiTp3I6M9C3yzz58mv0NMwTpckVCDcFMISw/6pyK7FaIsEwP8u6m
JUnXSTx3qmRjNagcYSqZudmL2q5DPEMW9UDoAEzIWLTizyD10ziQ2axBSta7A9fU
h7DiQpu+i1MFTLszYJNHMOvzGG+x7f2EnUk7pIJLFumV48tfJg6XLlK6MbC5PEQW
xexy43uUCTBzhU8UFhJVnmKyGUPNjJuCcQFTi3I2ILxqSpT6I3HNmHSqmrkrZIOl
b8O3ZLoBYgrznNEZeqA05cgzPfY7RjAFvDuA0OTfMpE=
`protect END_PROTECTED
