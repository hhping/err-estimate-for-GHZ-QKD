`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t4VSQrvPHZZIvHZho9gmdQoN68nH2wcSxbXNZctaQsbRUMpzGrsQyKwJJErdBBSq
TM+ydrjh08gO+B5zEkWuE8aN0ToaZ7M1kzoJQXyspopNHA223DvpWpDPblGbm+h3
Dmd4Jcd12rsAGcEFxu1yE/DDkYdHY7YGGV8H90xDnTALloF/xPcaKLF5BW+Oq0Ho
EO3/gWVVAmijlDECz0N0QYQCXsvkfdKT7pGuz81n1QtaRZZqzi109Jw637X0yZWE
WdTKT/zZSenH6s158pgHZZWCNpIHsJ8UhPH49d1sXb5+HVWLAs/iEkiS+EAqVcaq
y9vs9CZp4Ctcw/AnKvv/nrdbsfl12b/Dk0tVHBQvd33SiDToJH+Bxv2sl3MYhViE
dORgU/svvuk5vkp9g0uuSvsgK3//mUuycYZooIc99FubrtIxGGLMLKTg5Knsr+XH
y8DLsTRS8EJQXvEFaRuETBmBP6YCQqnehUgbVLl5GtgDwvx8BUqViTL3CfdOk9fh
3iNgeZ/ES0cYo8A1lunNkCj3yhQ8y3Lvic8xuZBFg2xqTfzTMYQP/BacKq7b1f/o
qAk+eZ5BCuzyOXAEGc7Zo1NbWBPvUDiNIcmqCJ2IpMi2YCix5MjTXySvMz+WTLpD
NSjREQYb7tRib2/1DI/vdPXbhvBCc3M6ZYYgqWMvu2ieXcpsRVXWMzvPaznvpjK2
zFEB4p/XHrq1hiiX/OgwiGIwFEJTKMif/XAZFiUwBiLSaBOVw+ntogux/aN9v0FF
MbHx6hwICLEarnRxec+GsxCa4ghWVLUBoKh2bM3WwX+Fl3uLnifnmKR4U7FhHxs9
Qx50kABSzbLSlfm4ed6GhFki8UxQzChbCeeCiFU3tZFV8pnMmmYWQR3JzNlivBrH
tf38pCzOKJLoo7b529UFFWKRwxXcaRJJuIjevauaPUFInQCe7MZcsZIQU1P7/p0L
TOeN7ZzI4KW3kBdY6JU7FA/o1/DfZUWQO/zRVXAaUKlMpEjCiQ1CliILArTNmFlK
bcnoSNIb0Hs1sR1J4/G712/XE05FWK4QcleAxj3+SkxbMQthvoiZ0tDS03R2qvas
Zrae3mJ9kZQLb67Ti47ZGGYOOjM00kgIO4wZxt8VYWdjGwHIfEKODImp1EEQzVFc
Q1yM6i9V1U+DTG/uWvWBBDwtigqPLjlWXePo4oLBQpPpx2rWQVtNXKIjctwFp1G5
+KQpNvNxhAwGELYqIEGsC7AtZqbZoqfVfQMUUJEoTP4RuDHgnJyJv1gyEUXsfYy3
bT90RQkIvtja4LVljqOkqZQrqS52Fko+TZPILmRSl+31A432s1vkZo2CH5a76cHY
grm28jBOGAGxjVRP+Y6Aql6ZzCBC2xivAucRw22MebgvvGZ+sfJrz1rDoRzb5yQW
Pjn96nuW72pj3NcUeTtpKjZihlkX7aE5EmjG8rmj3vYCPEFPxCA8OJDeOyDkKX2J
/HCQTc5qC7+RQWmhmCEYTqE0wp830OJlx0zRF3cMDPyLyDD8S1aRP40UO5AGXt8F
r1duRa/I1CePrgIBWaXX+psSeFvugF4LH2kSUnRIhMvXecOovBXvxNrTQAMbcZjv
Lk2R/Zo3ZgxqGlPdAIRjobHv+LyswtyN4uFNUcl19vanoAeXQIOA3ICiBJywjpjD
XrSt+I5L8yzmQoylOnZ9p0lysYmlDvoo/eqErcfYC7KnRFOFDbz+/1vYFw1vnbDg
MM3g9MYDHvxTIVhptySUvrJP56Qk3oeICQQkL4nOK5tlt7mDji5raV28N9c8XL/1
YVDu+UzsAxaPi4CQcokjIj3OsnOFSMjo/xar3CGi5MMeDPvf1jMXmxhgIcFZ/jHF
hGF/KIyholNamW+tkU13cw3n9E9mpM1USZpeuD4QomdThdFrabILrrS02YbABZXY
sjaaExENCC441xOBw4KKPfpCbFJp28ydRLtkThkSYZDkxrVwmksVI9ixrkNPv7hB
BhekiLyvGOWFjd35jqsreSFBCR9/NGaml0ADORJ+mmiykYB1gPGADGc8rICKOZ4L
4WPzOF+GtxV0FQpfUnGFaxwcQESoAvV2ez1Ezm1cZon8CT5UCnLOIKesMjyRug2C
6c87knNk+K4K1VOkQh3WeMWzv9WjGrnGEJSF42ht05Ipiea5Igmb0gazHC6oxol5
/ssR1Zvdg4V4fdq8GCIJB3KFDBmtQC7QsQmrvIgJlXYTsMpgDvC3o88z3SNQDr0w
iipEA1IgCAYTiJLfJ4kWTg==
`protect END_PROTECTED
