`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4iw1hQdQPeM2UI11uC1w6wJai+3VTZg2SF8hxVaxSEQ1Itmq+Yt1GOdVFTGmaKpQ
sA1MX3yAjlUQw7yQCC/qRL9Jza+Eu0VP8fzK1BuyKfHfc5VMMOf/rs+3/DTq8W/Q
IGNjjupyrJ6W/uzW4NApAqWUYm2++S+DM6HDIm86AC9CK92AWoEg0jX3bZ2ctGJ0
kGeai7n4+LKa5m2/UCLZ8U12GnfRzk3Wc1IgSAD5gO9f/KPDi+idjtPrZCfR6vo0
niYYkYhsCqhlfhHmPwLSGwUjO0bHdOKFwG1aLpYjwVmwBjkBfajIeUTonncDzPYn
JGkdnZdPDxtOJDT+c62kLcadsVgoyyEc9hIGIWNPBanIz8mk3+sVG+4gBYvVl2hH
VW0NTODoqHJWHzZOHpfEeA9Oqfq9fFBdUUzqqqqILY2JRBAo5L+bP8isK56gqhVP
a3a7n8xFopeqgWqclEbsml1bJVSBECTxM9ERSh927bs=
`protect END_PROTECTED
