`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Sj3rLMnuAfWjaCyYC6XR+2fbTGHm5KNAp3AlQuYJl/z3p57vZa2HUD/C81ra/s1
jc65wjVsLIe9LtkVHlI7tXVZZHtHVq0w9vOZXzel/6bPWIkr+hCLgNMgIlUJorY+
+chWU8U/N+rhHdftRWZyxEAPmnln6bFBgzvVeXKcEt+q493vK4HLkc/sOyUvs7Vw
KSLJ7UOuuNcD3nGVFqo0KxiuadK+QSDKHKXT66afu9sIlwD+WXAtJjBS1mKc4/YZ
3c/kWhhTHrFVvwZaZ6xpPRahs0nlhyb8oJ9YAtMufZYHXovhBa5kxYZcXBtLmA3R
lnDzQqJ6LOqpBZZ0HksRLEcYKn5Y5RSWCTRayfR+eLm6Jj5v03SDlQVyOB2fw3pS
3HOB2u3qPcTiKNsuk/pP6eZp//BNCz4yBcbKROMmXklGuIBy+1vC3zOvquZsWJ0x
RMhBq92sq2SES4AxWBaFacIBEwJ6mIAIOFD0+I9an7aPmEqkJz0SfxOnwqtoDrwZ
Vca6/a0BPA4vMa4lLOc2OK7kDodk9EETgA0k0CcIWnbcoWl8PMSTAoWLheuDU255
wKdj7AXfI8eM1Gw/X+cv60uxErMchSa72dVPynJp+OG7q2HTT9m0OVmsD694u/Qk
fcCRjJShTA5AD7rJK9IpMYNZrKDdZKYzlj/C8x/BMb492GE1Mj8nwDhxwW7t+hYK
LD9cJcSCW1olc7KpS6sULY5MFYam/tCNRW4hYPK71Yq5uCV7kAFN73fUu0VHggNE
pwYf+a8EmXis/YCntmeRzxvIRHuqqeYLnbfc0auS3COkZYiKcc3NmRtDvg7UWN8O
+IsKS+c5onBPys2LoVODOpotRrwlsQJy9Kv9eGPqe7wkdGlbRqGACxjlyg5PMtQ+
kcG9I4jBqOSrUGKSh6v2iE+5wgxFW68Y4G+DkaX2YNi0AUNd5WRvaeJXhgs8X882
F5xQF9ODixDnrIVIfKDtUZCR/18Q0BCtFuhZTelmSfEepexJoo9POd7xQmhBEEOM
OFNfPQpABduoh9rkhtQY3JJ/zz0VElxfHvK6IrOeb3aw7+4XSJbLavM/bmeY1C6n
RhirWcRN6I4DF3AorqHRV9Az4GMj5lPYDDFovykCO9HgW4f8ssXZkjcSk1tXmQLj
lID/xL0Sypjyo2bZgC36yKxUliko6fcrcZQfp4vj8AtFK5HfHB5NRRERsc24LEZ1
0rvvByom3r5fSsZ0AdTufO9RzWdvPMbDZp3SK7ISm7IBvtS6SLAyZg3GmAfMrTGr
2oaDuNb4DBxYK/nyRYEcecS6qydseOC6YrUJ9Vb5uE1gFSIHdOpy11HldeeAFoPq
ZdWYFCyd0lHcnQ2IrDdJd6PmJdp0GLURXWPxBe0iF2ZiOW/vG1zkxJmTJDvMJi94
3LBWRiEJuHOoWiNhI3pvqOLI5zZmR3JknckoMqFRjloAWx8uQbDXjucdnSXXrfFH
ZD/2Z5XLvPGsu/ifFbQgIAUG2Vg7kAMRX9tPsFD3b3beuUfvOpql+s5fwX0xc53D
64cC3+RyFast3w64mMTIuwwepx8bvJLuWjKgpMDJ+PaHlFKt+Muxntv4VTWxywq6
IxgaLl5JHl03pndormAKxTqGcVmEL5s2qM77gTymLyi7WmUVFKNix6tEPjdaQ5jS
ky+VSG4TcXy7iMlnVYZ2w+OJWezPnReDaDqhGnTydAGRjc42NWzUu8BSPBFzUGv1
VmSXEoANuqSAyqqijSGcsxXFmYmj/tdlk9mivboBvad/xJRI90h7rSxlBFyZnlqt
655C+ZV17Ss6Xuz6MCnjeClTf3olK7deuDpeq5XSNG9BU45kiFwME7FacN3VHalQ
xjfdBMZltswVy6j1VbVrSDaQGLw59Iuo2L4o7gtTbxn/W7Ig4EvArlxRDnZkaJvq
fEy2Ih6MRWdHFOe726hsyHfFWcBIS8soM5Rd6sEqiC1zQ5eEMs3JBoun7cXMMi3i
`protect END_PROTECTED
