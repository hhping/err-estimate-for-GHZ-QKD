`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZxOHdwJ1Y/7P8o4ItmlWfW1OgMFmX8o0o6PY90+SW6pLgVcIq+DAqdR280fEbwX
UhdALn6VfRjpAeFCrPZGqf3ayXo1Ykl+GbH21hONU5RE1PoiHp14jDKgnIu+RaVv
Pqf1S18nVp3Fp7loSGbh15XwCXGOPSW9Q7o3mFS95+kbAEafEw+76o9+CiDiQe8E
bnIwdfrMp8b2srHgxVd410w3MK5ApErBCktFxyCy0+HA6F0rJgRF+TOYVy1KR8+d
VWQj3s5Nrz01c5Fgmn1fVZatuIu/EPOn4x9YQ2mmY8lvlGppH2Kvi2VCOoaPLkbi
+mG7IdTPGj6usvuWL5UNhtx/0N2YXlvy2zKSScdIrzqL9UgVW8BVCO0ERomO85fL
PJFXnWVWwVNUG288YAhD63feAG+Rw2nxntKniZcmaGEXORjUf/azEvDbSkZMCh2i
feff9B2DMrTCDI+z3J1Qgo2Ws2K7+BmJk9pOrPOuesD4KiEJj6iKOHIHK6r/KrVj
eElPOvlGzLA0QeTar1SzR7d7wEG7ncvcQw+2cQfTa92IumUjqWuk7u9CcX+gWDqn
EsPbxh5K9InCf0gw0jXS42HhuoE5LuGPha5XNw0d3zxmsCS/Nd2/NncABmqyo+H3
/7Kvg7wPfq+3TmhhqZiUnirzq0pR3GioTR591o+GkQtZu6wfeB+zVqlqnXPWrcsq
xFxtjL1PpnvEXGnLeRRmkRTin5Tt1xBK+FcFQGKS5RfC17U/RWuqrdPXUCklhBjn
XfrJtfJGiUhasYl3IN1imj8Jg03cjq6ziT8O1VvGo0jbFbscTMU1rHsxrY4Tf4XT
1SOwBG5qLv1n0fwfhXvHSJXy+dwAfOLwfkcF8HGFqhKV25pbBC7r24MrO/x4jfxz
3/JTVvfcB0Wx368DKp3uAFNa8nOekYpinZ1EiNVqP16AXn5dqoXZ4DN1erNQCZYB
XueMG8ya3iC1oppsx2yRb9VYHaA+wBkSdklbeXrl4H6q2LEsgQJLo3qH/TrATX/1
T6WcbQRJInR/1EsKvKGstbAB9AEKNxSZwM/fYJjGXMQxtCEYCiwgWgioK5DgDTMW
4Va7p8xGcqX5oEA4GXJRMcjaCNn6HfYvuwcZYA9GNNJfnD63JFWT9suJKnXFiHO2
xRBd+354gqcCHvsalBh9HvYj7pkcKDopbIzPoIo9+qhAtY9f8ZWtObNixy/fWpn0
5MPre8C+QL9FBPKiwCyfmkGlP+g0dp99zTLPn4g6ho4eIDkIVUs5hmePayx6IrDJ
T6IWKqnxeJf+WkNJw1c4wBjI+Y7Wpdg5cT1mbwmyRRsB1AK2ncq8V8dowL5Tyr8J
noAFUEFi7YuQXD3ax+TZ3JQzVJefpOUhCnNneRHLKmFCoNoNFHQ2AFKanheVOCUC
RZsr5khtcRK4f/OVoy/PwQjIwhQYmRQeiE6eGbrpbVkrRLtQoIEgMuerCRE4OKbx
Cyvl+pIo9Zk9G7fi5voWO+EhqyG8SPrUCRsPtZSUx6NeqtYVwdFacA5q9x2WI6+1
70LQLBNKmq+KYHGw8NiW6NFWtIfMBPqrB4elvuSH9fcRbsDXHde7MwvWSe+FFLdy
2UPRaisyA7sZWNHkGSwosmbeMW9EZRM1Pl1Jl3TMIJfU+IShxUdkCyABzJYXavkK
ENdDqrvuFHbK1inc40p9iu6IlECss+W5a6y3hYAJ80W+RUFigRFvJM4FCAeudChu
GxAL/cphy4M9cLvoysPI0W3GuQNGtIMHN5cXiV1psy38pLjpbH50yfm8ur8LDDbY
dRSfc9GQclCdCj7f7z6ca9dlAcgd/eCP4kMqtP8qpmVi/ZpB90Di47X6H51Bey7m
SjiqoJAtk8OagDTgHOZvvhKJGS5ZBIsBMaDLILl1HFszPjcCQaF0vJ0WgS1aRcJK
0Td/JMr5Vyf1Gkk5sCb9Tr5BV8oJn3JXbKC+gulmAGAB2gKkReTPUYXuPc3x/DhF
cj5L+YpA9t2liwjEuOXqxBsYOXR1jRfa3L61WJ8td44Y8NuRrTbwSVmCdKZ+uRBi
4YGMTr+UVuxHFNLUTTFIYXDUINhzmoJ7brPcLt8VAF5gYcQkxCTXyY9cWG01QPsZ
LFMjToGzjPRJ2GqPwPpmA1OmPGv54heifLKZF3XcF/+2kLOtYGcpJUrZN69x+aQ2
4P3Zuxoxo/Itb/IjB3O1I+2lgYLaBUD6ffEcymrokKEq/EyUcS6ixGMeiGleRhNb
JSOpyhaBDnFChQs2cochwJr+huuiavBZr2k5DudSCZrz6OZichsRZFK+wvIaGjOj
y82BkUTZdG4Y8qNU7TlrOJJ8IJ791kAb/hOnTE9f18zh9aHn1z1/Px31OzB6jFFK
wH0z5N5T9ltMNCGNw6rRHRAAiw2Ue9/dtnfH+5FFXUir5nMkQByyMmIjmFHVOq2F
isUPmfzRgPPZ7KHTYTXRdGJMuAjRrOpdF/bhtcFVHPeIeRd+Zm6ShaxrjleAIATQ
os/8TG2Zar3RsbIMgDIsNWoAYDYJtTvYm7csvYPdyCxR9qf7cvFzZtDlcZyVpN+g
Cr06cH/xz3QbaxxRydgUuYWR4p2e1j0XN0y3m6BBRFoiPa8iMyt6h5x/wwOWIjFp
K8/l8mivmAUWrMNSP7llP6h80HXZgVVm7r1JM3Nl4kA3yIKmEGYJ//4n/zX9LdA5
ZI+TP6uViq7BIz6tB7jkAJcLJIjv5cv+Bl5EFXfi9oE2FcGRqxAwYMAQy+do3nnZ
aJ+lQZM7dgDbvspRhg0C5FW/JQ4GswTWSqEsCG2abvez9KuXPefPX/2vvcamtBg4
wDlYj26vER1Cma720z4lCfxrS3PfsLa987ou+bG6nAYA3uVp9cFWtqYtQ22MGX7K
2fibt+JqHULEYKaNAG7xiVn8DaX2Om0TT1DLsiwovKsDpGLtW1lsbdiCJwLFNI3n
WQnmq6c4U4fBjkTQxdFbgcy5m4kXCQGo7EnplJmrz1PKFCx07L73fpcr0rsOxTbv
5hhZRRHA/ezjGu4RuA9gTVykiwMl4SYvGoLv7Q9q89XIDmOKP6JYJy5WKjD8PMUU
giPDQTWTzON2pj/FsRL3ENFGJCEoueyXD27q82Q8Xk64FNS7lx57s9nXSo98tSs0
xXdH3uxk9oCgoE1JPtr4eFvTHh/A5M85IfAhIqAr+iN/oioq58cz35M67Mr9QBNL
Q9oN5YmeJsMYkr7JDSBFOnYPu0XAZxxoElv8lScmb+nrWz+5CIrBmLGm8Wc282Lp
QcBnkyz5Z9pSOyhsqwpY+xPUV8XH/gVAd8CdGO1fhtPig0kk9eGwAn7SLbvP3dMO
JiYQ8B4RfBEDEr9VTU9QofksmzeALdEBuDde8oPA1juBiFcDy/wTtyjtXE4zk5M8
HiNANEzDgpHSSFPkRwQx87deZpdr3LU3vw8ExXLaGKJX+jcbPwdD2AyM5EHqKbLO
ffKWqGxwODgqs4fIfUVREZ0H7SwawoITaBwNll5875wKAZoESMmQM83zRTPL+S2U
/THBPUJ2JKcr/WyzrYYrNM9/avj8fsGiyQDJ/4EP0WCxP+NTBzZ2pXR48AOpwN8K
2lFfjlX00i+VMQuVREPTKpsKS2y1T+319Vg42TUjzjk7g0N0UXH6GaTi23OypCdg
I6LLTxvXzG0zBHgYPhcmJW9qO1ZqQjj2dn1jLHSDJ7de5z1cpGnQm2l/Kz6Wa9H8
iIN+xxpaXu5dxVwSbi7AcopB3TuaR2yuNEsM/7u2+/Gxh9avNDQR0pMxkfWWSsLM
TIysScxaQJ2bIiY/mFc9aysv8v1DVv7TIsTskv6/b7nsKDd/5c5jrEC2ydElVQ7w
GZnyL3xRPuT028dkP2iGODJbD6eUB4pcqV+xalTNrVAEJr6HNptiZe974qdJb2AP
BU2pzo5Pd1AUAxqXO12z5M2Xq/CMaCBSjm5B4jVKdeg135Xh7fR3Db02ScRa39wD
7Ut3EWui0d14qSL0M6Z8Q6aPgCyiCW0PeMKunJAeVQEEdPABcBNUqBhTzzlencmp
G2rvyQcSDr0hnD+0FmOtvXH0S8urRP7Y5DJYPOzTVHsm53fsUEXnnwzUK3uqK+Yt
jDudIDNsoQ4kK2TiB6m/mt537vabQ1VLBZb0To8XkeRAqkEZEbE4CLpOX66kIXoc
jwc+YpxHgBNW7GoheNMiK30XozhD/QL1PihWernd7B3x43ff0AoMnAhDawveAX/U
LwjAk6hvvFSIFMy3D69rULpkCW/HtUDLIxdyumYDyw0HsUl/QfS/yYOV0hKNeNUO
drXNFnFq/y93IVAovE6OtJDFLQLivJZJhl8279Xp+D1VQlDKNhlfe5xAZCMg87xe
eEwLdpUZmWij8asTyv5AB8USceVU3qBUXnkbZexNJy6thkleHRNgHjNJllY63k1I
nXeB7wbCy4uOBpcAD3q46rycDLF5CIYWALImGnjQgBXKmFZ3BI4pRDXNKKU5s9QA
nUbk7jhn/Xo3GgkZdOl+ofW4smw0f4TtldCcyQU3Yn1Q6YTGAVYL+QKipG9Wr1T2
NNGdURIrOXzZlvkCtEakyAklwK24tc48nvfkC9oxe40CCtjJD9sYv/BJ8nS6gmRq
UdHVz6ALRnGP74GvSAh5Hbxiv83H9pJHpOjgQZXJMiygqBInPd0jO8MjcSb2EI4f
8NTeliaMgLGB5TlqkmgjpnpWeDwNn16Oaz3T3Bp2MbcZhgv+mWY3QHwaR1GHtNJS
vrsy0HyccNRhJuThsuMH86uEuj1t0rYy642RLhP0r2HSrrqIZQwly8m2RzxkWa6X
nvaH3sJdL+JqyTHFstKDqEoyIokpAxcJvc3VMr0OFMntPFYhmmDq5yh4LM1+89kb
KpnhfU8FNCaoy1qBEXUxdlZDSnOwU0oZtkeWgfXV/7aoDU2f5BcBrpU2nvmse/hh
f/AjvxZjzruUHOAKePwvp9AyIGdtv7zfxlhMPPVMhiwFI0dMQ9NOk2UogQ5QBVD7
QVz/scZ4ettBMQS0hZqxss6eSpe1BOWAetxVS52YgrGOLG5py2xLdSP4oAXHEc0l
XbjewNQWtX6jcdC+swlengFAy7909pbmwIYVkDdRmFiobDHIY5J/WM1bDsLopMlN
KR+ATp5wd0ayfrrAlyUCD87aHLVpPmG+qS5l85QRLPVbJoJc35QDrDIRB3I3p6F0
WZ46lxbqlemi4TwB4pyMUvk1tO/a6RZ/2PO/Pk4LwcXvQdvCmACxDyPuSTH6wKZS
rYk1uwE2rFvQ+Ch7GMqK3hf8hRBGo6BT+SDxv67DyWzLG0Lw4EkNwIRcleWNoTQ7
3FffJsJpkOnkTKvk1DFJJC9+rHAExZ10E1R+EdNTnRZtuL8wLJg7WAVYhoTzhSuX
gn86K07YXFNiv43ka/sbcA==
`protect END_PROTECTED
