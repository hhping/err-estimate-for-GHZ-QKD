`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wIY7f3IrK2dVmNmB1YAwYEeE80tZ3nF3vKQR8pgntF/iSMkWQkoB0q+chMsBfUl2
IkiTiyTgYz+bM8/dCI1HHlMkJnhoXZva4030GN59xGLQi/x14uJUiblzULU5kQKL
9ApdNzNHN8Q+vPtn3PCUiFQWVMn3jhPuB4b5KWnIwPmUrF9w/xKWAXX2hadYgU32
kw6NKTFFooU0IFUDNxh/2Bh1TRcBvqv+wLn1dH3SnhNR76vC1dbzrVZln7TWGzT4
dB12d7kahRZdWCI48bOtkOHtQ7DkdzvYVMdCXHZntIB2QKvZsaD8UMUALGKmtWeP
8vgJss4bGmOzev5nkqLHQJoHxxktWOQmWe71lQomVFhaXSsOUnxJoAP8fi2flC3D
cNowoENOn6KwHt8/26qkSBdeRu27WdBa5bPyj9oTEPPAMbA3o09pDlek2gIYabtw
11v0WsQ9ewbztL7+uCkIC1y2sSA6+ZAOCANiAWaRZGJ480AlruM3HIiIleSnu/Ph
vVbh/zsvIsLkPitwfbHzcNFhIVAA+ClIc3ZvLYIE2Eos3szJkbw7NA2qq3IPftJa
WAlbit/gydY1Tzv1RLJ+2HZzP9LY8kbxYVkVaNg6QdngBboadcvNc4a3JgkyDFuH
Ra45P5EMrQYEq3UNV+oQyQb9kLgcruUqQ0KRoCOCMs3fu+aebkLjpJ2DNxvnvyYu
K95ewtdphQUsLzI2awl6UTDLqD8G+/6ziF0yYzNE7LDflkFyyWHD0Go8Jr57vGJb
0fAJxCrYl4LEMXFmABKm/VwI2QUFn0xmKp4CYalPAKFMpMfL1WJbAWrGVuPuusMA
UIc7nRVNNXhUBtHknrbMIzEjGtolCYK/oL/C8kz2urRbV75LqwylCgug/7ATWyCW
EYA1yyxtjTydzBMKjCv2ay9bd9d87amtE5H90QWCtTj+ksRF+fe7Zw2nIlL7gcKW
B7Vt2qKIs3adpFGmB+awd06fWeS455T0Jb4q2dJoMacYuiPoxkiYh+7mUHuy2mR7
63KHyqdmkAeMTaWfmqjEXPw+ZjmRBKAwMwxHxXNKguAXPUbw7UGcIdrYaNYPYMsN
1JGPghVJofx8Kzsok5L2CbZjdzWQ9uIOAZxWN0Lw4m+iyfSTy0zxi7KyRLLbf3tj
THmk0tlmfUjZYW7iYqDn3H9tqzcfVuWrU279dKhb49SfbUIG+sm/EVjoULPbJXLi
+7dlcY3sIMcrwANdT40KIX41mu0YEWkVDkPyg3SaCO5LXESQNgTw5UyH1bj4QsH6
HZ2llFW9lExRtllR4SswqmmehJU5K6NEj8d+wm86cCht2eW3GuGEtGJQIwH0dn7g
Bea9R43y86wOxqh45mRyk7itj9sRZGdf4oxHXDE5pCQ4BZ5tGtzEAMR7hQfIlZjo
7F0nygA2dXvUKK+vvfPZyBttLWloI0Ii3uTT3CnOxxYeGazQSG5+fNDZgpp0JwEM
aQ40O44PvSKYInyFoYdp1yObk6+yWvN0dft87d80YY8=
`protect END_PROTECTED
