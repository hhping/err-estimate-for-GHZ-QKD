`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3y3/IIU40M538TIV7QhNVSAbJJfFN8qIDIg/X7fp1o7L6ZxvbXMmWvSLPXW1Of0W
vV03m6e/0jIcZyXArkQCjhRWl01dHwBGrmLwVpHmD7LjOU9nMNlnaR0GFYflAv9y
FEtpO6qMlKDvXzJt+9HGKdwLgAYZ3d6ZMVub9k8fYuGQMcrHLk5G4rY86f9eugjZ
igDIYMZdVs4zuZMQ119F6LQ3AE96PhBK5NGQRPNLFh+jIxCPqvBzxdegjEsdkali
vhqzCS3uXd3+I3StpkyppIr9tsnnPgM3QBZH+RQQfFL5F0tLUdgu0OI5IqxJK0fD
020H+lowoP2SkGtRebAEunJc83ZlzR0hBB/pJpKCR1kewf7Gx2S0fPIMpRAP/QDr
JZasOiVPc3Rvt/5jZTSsvYGG03vG/PLr9AFffdrhFXG9KybGDUrU7BTesnGFV/MV
6dbDeDxkIDrA7WY4U+ICSHwhb6Qp/QDgIo6XXv9PxCl1KqtwAh5/g4BPUdEf2VcF
GAQ4TQCmFbs7apwHbCoktwZgWHLUCFLQ9TwlivttN3ajXFFNu2vYAfFB7CdkKi1C
U/YMC/UlVfWJOExLTN64+0cyaylYlEofBIyJ7VDx/1ykIa1YvG9kvwgqZVMa7xe+
d616hwDl/q7zUcPcqQddu3dM4+MXanx4hOF0obm6+m0LmgOUbXEoyKy0+UlqaLJX
rFMO3kB1bFqkRORKMAirb0xfQ/bd8vKbcsLQgi4F0fefXBDxSewPi0YrgcCgAla+
RDFJtIM049nc3Kact3sxRk13Za7Rn7WvvdelWDGeDXM=
`protect END_PROTECTED
