`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0k6AloYlQmhjbf8WbCn8uG7Yvjmb2RviYkffCLKwajsfkx1nNyqJ46GQSx2Jf2x
cAnWtrUcm4gQgO5wjWhRb9Zr6VJL+TDuDssuQTDubFyrXQaghCx9HSArROm03XVp
/ONCRprvWd4l5CZisrilEMdCoyfULNnC2Dn3b4WtdJdksZu0++cVeMl42n7K6z6D
KU4W6CEx468fnOTVo/pKHJC+Jiu6dHxxVYmFjtiT0fzEXEwWnM4u9R07bQbpYCQ8
taXlEaAiwAkjwkHNhDInVI7OK215lmQe3SHlDqI5pFjmiNVwv4LMSajGcQkFXQgq
1lYg6cERSP17Q/8jNSo2g6JOBndwhzHyyT4bwcLMT917jA8iytiJGu494EDLBa4u
m/iCFupzsJrHPsGpNh53F9EnGoGdAMxAODCjeEIZbJx4U8Kz5RgGkrEZ2h9ELxBI
SBjc2pbJgqJ3FV70oyqkA/ISa8WPux7ApfiW53YC3PFYUBaMVzBMxGV/hYZomZkR
M1H3fVdWTBernt63Gz/kRnhvOy7mt6OyYS97gAnIEqyW2xS1+hC5KYjItpP5LYEu
HqeFn3fMLIjm7KIT0c45ARWeFb7gc136A+6oW2STYTIrV6p5Ms8HAEaUUw85FYo+
6dfmq1ASXGXzBJT/lUtUXK2nFVjPmVLjPO0c3dqN5pjpZaOxQSzS6UnUlbEjTj8u
Ql/69CxieFRllH6Il7RXmdCNUqPGv6Qh82mohpA6Xixh2mAKBL9Kh+x/vqCEhszu
TFdVcz8c86tAOWaeCp1Lc75F7gxekTnF5Lgb9TadVd8irFmWGeKFezJMAo8H1r32
FVi1dP2eawBFJYiLjxsG4aFWMV4eCioXXxSD5mPZ4uCqxrhE99oLiYM0P3x75MEk
q+Xrz0WEVl6H5gECHBugQoTtbBRIW3hSWGIuNjUXajnj0aR1i6brXGkzPXfpvYFQ
VF0XnC0Ay5yGPn3lyu9cLLSyvODdZBHDuhCZvL5qVCs80RCCVdn3tqRNDnutSzFZ
CkpM9oXISNz7agEwMUfHvsS0quPZR+GcMKeqgXiPidvhx9XrabzFYzSACyVfT6Wa
Szljwvuq2/lgd8KS9/qtscaQZLMRVgkUshDL2IKXKlhPml+DgjStI1Ja03wLjuM5
FegAIaf00RnZY6Yd8cMoSBgpwROvUbZSkVIUXHmDqfCOodd7WkAQRZ/MMZNdTPmj
95t0VTVzZeJznQz6Q4zQrgOAis+PgSmTsku1NhFBDNiOtm74kKMy3RYGFwxDQgTm
BbCxgAx+XoB6v8gVTo7te8moOLVPsCEoc5NUeKZQI/NTuABTDQEKchFJ5a/ATT7+
p/GyF2t9+6PrSbcDr9oBUa2i0/z9WGb+VZzS1hprcmeJ4/oheq5T8kdqLmiArXR0
GZd1tlx0HBsQC0dwSTLQB4IMfhvRBVMSfNQVtBVhBCmMgsFqghTrOuh3FaMlHoX1
3SgVjb7YbjBFI42qbFzhwYwI/l3wV1p2BFHaKYWa4RzhpeVXProOkY3MBXFMbOCg
Ca440/PWfFLsPhMvoimqA5vJR6Cqnc4mvG03yFrfRnjT+V1YzMQzk84ZXwsPDr8V
Isanf0ABeUrao63tuz5n7t0wSbIFMluobSekJiP01L5Z5+zsjWW4vgZkfIzHQLwh
W+qboycKyBwTwYZoFVWXXiPKcuxzqBL8mnp0/G2hwpmXRHLe9WxLW5z06G8Pai84
jehMgUqh0bgvDJX2kldVTfRX43JF1oYWtJWgxhhrAOmldSYs9mkrdBPcCxVg1hYJ
SxH2IJHkFL+Bii1TS8Q85VL//DPNxKQeFMu7FBjYqef+OTZLhBRqm81y6Y/+/7oY
le5mDnpTjQymmEgampc0SzeC82oFjV9iRXPJ3x6/mbxJ6EVIBBm2hV2s9yZT27y8
wVofw9Yn532XGk6/PPSE3bWQt/NfkRpmjOWqqx+o7K3FwzcvQ+Zjk2qvkvhoMfbj
J+xo5k/UWzRDcjz5WTGg3ml87DScMt2jWVKqvHl1h6p5dM0yuCr3flHO8nNSG5OY
K3zX7nqox3sUAcQ8dZAkc03m7ViY9OtWQUjwOwV8nogiaAT6Hc3OaTpvLF8byI9W
MuL7EOCN7WpN98fgg/ANSgMFwX/X08XH7wn78m3rnTp+xabNrubSrTYWcCytJeey
OqE7HEZ++589pJrhMbUeH/VlQApW02sK/ziMWN30nkQKIs3IAIYD6LjZVoC3qtxz
Wna9aVPQHO+w9OwFvk13nQdY7Mx6iTAcz+rczZguJG9k7JIcl1216Jcanf/tCfxN
YKTPpHSjNFsfckkBg8l+rTj/Ak6UNiBUf/TOkWJriBBAZum/vBtpwUtsjPL8TOAH
RsOHB9S92PJPptqNRos4OkonlbgpskQgyKvrOuUwqxFKzpqGD/zz4xaZclTz0Xz9
SbjLZM5SWRo/ecB+NqOFYhbSmDyrpsz+yRvLZSUzaey58KO9SlZwUPgkDyS9no3W
bsX+GUkg8DJLj2AB3hU8mUm+QdJ1OI+wIRpfAMfNrSYh8Sw60X2OoGAO0x7pbyon
MdPMJBSBuOLsNjNWFtC0qQOWQSNENMlNJzKSzoEhPfSJXhvILxrW1iQtJUW7du0L
CsmgFNLgDyA2XM1tfbDt0d/EUEKGpOqvaRQp7qCSQzegKKzjGAGayqp71ERMf8Ld
mSZkAvwMYIvj2W7wlgrRnTwBAJqQWeXHeMdQP73pQJx8AKqAKWaPrNLUYmxBuouA
g9BInmnqb9MBQu3NOOQkr6D80CwFKQT0rf6HB2sAYYnW+6bHpdhR8IuvBiXgGTGQ
4jkEdipi+MlAKl9vtvnNHivLs9y1YSd9W5z9+KDDiW3A7k2dM5gs+U4/HBd/8hOq
eYy5ADvmQpy2wO4LyyyTJigeo91NU51e5ic2El4APA+YJOv1zm/Y/IuaofgmL3e7
H88GKrRf3YaHqOZFLQ2gi4P1CB9Y9evbNXPLobQ+GnRnCZiyXnRdjjO7dBadxmfV
2RHIdZgxoW0k+yjBH73L+tjQzxgSN0NCgoKaTNkrynp+RJhL9C6PLXXyZ//y1wuZ
pQqa8x+cE6i1S7bhEVXFdjmgWrvkmrAIm4SfYaREOj9zO0kWznhjEWu/Pn0rio5j
O/fzH6BzHMFgPI7Wk7FacxNfNO+CTfstAsj6gjPAWgZf2j0AwTOjR1Z1hbNTpX6Z
Ki45YGBNTfvudrpp40xGt7aNjKIFXV6hcnADCaFjQh/H/kBQuLKKJ1W4r4PZJdU7
Q5cZyCgYAg3chVM4LEDnQaNd0qismw01dmK8McUXklndcCUJufVKshB/oIiMNyvK
LfesVX/G6mUQ2U+1Y2jZIb1I9YS8jMVT/fpjQ42qAkK80avD/LeRgAAFBrU46oyS
WlJdF83cpvhsrWwP/fl5qued8bOc5w1/Kj04sUjE6c0vPdsKs3RPiEsOUQj8+PLO
fKYYXmTJq/iKQegL6Ww4Wa+TSMEn/GX2Fp0XMZIna6uCa8L1Xx59lQb1EwZsxGB0
W3yXzxsGzutLoGHhtgNKd9eGhJg9BuqFPACDdcf6dIEClwkdzrUmJzBtie9bnDYy
vriQ6TYTk7COYqtSE7UAFrInFyyuSAokMQOlM8qDggI7ctXZCsA8y9rcTgRgZIUf
M3FBndGpFm7ULMPcZI8UDmWfjP1lG4EQvY8kyIN4DSRsPzG85Smo7SStneKUserl
KMvqTUQqMTapZIRtsE0JbE/gnGjBAK6cMmPWB1GWL8qLAmRITVeBE5DV/0xBSo6D
bu5hO7WQxAUWFeNSeWqOpU9IR2Gqmz+YZAL9PE2uuZxNncBsqNzSvuQn6FBIEijG
W3SIFHFMAYdTO9lmYfMy+1hXWmKWbcObFfbRRrVXvxTU6y7TxxVy9FtGNRwrxwoZ
8o3637WIx5cNz8K+1544INzyCeB2een6Jo/9xGukcjQlMl1qOsU0mc5s/Q+orNQY
MRwkp1ppCLJ3wTkUBWv2EPy+v7HxDrRKxddGr6oDWEJvkofa4thhgRMezYK1gcyI
DzQ/o3aUOqfJPgrUdwfxdgqD20oPxp1Zhqjbf2OYUz+x2mbTdfEmp9bNjikjd8K+
ODroyYjvPzYUEVMImCIbmQ==
`protect END_PROTECTED
