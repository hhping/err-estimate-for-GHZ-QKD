`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wixw97Yk3Nph8zYlOH7ODQtI9rJTjj50pVfDyV84Il17J91BmW0kbtxbxC2C4aKs
p5D2LKzYzcktS0nAwZyLwcIJFGCD2NumytQKqod9m/ro0DyVP3zDa9FKhfQl5g1Q
OeA9VHxCGPAHUh6tUvR8CPV/NsyJo31YhoYKI4tRPyVe8v7Awbg9h3y5NN5uq2xi
GVrgdhOPyYCY5WJiA3nhh/ELBQ64qiRTJ+pb9OzWumrQrZ5VgBN83EGTgKMexJwa
KKM3LpGh2wxqS2MwbCs/6TfUtglM+J0dPdoKlxSCgbs3xgWWURs2Fe179uLJBmxk
HDjWRtGhpxWSxs2TKfZ5jrDWRRq41CKVN+sk0l5+/538f983OShK6t4Ox1D+/Wa8
eIk7L4TsyxXk2aq2Jw0nxNri7q3KgrcATlamRapZzxkkKFYssOQiJSnBV4ere9TU
e3uHRhGyDU+SCLn+bm56c9tSBRyPdmRvJ8B9d2b2qE2w1SPMsba4SQNe2H7AMz7R
yfMX0EPeQEhB32gP99Z+AVRTr9Fspd6OsiRb+Ps55rk4i/dV02yMLSXSt02ZVX+4
GVnTgR8fViAWmrjcBS2IhaiAiBz3m4BGLeriCaahpfsLLlcBFi9qQmitBlF5lzvM
pKXwOGjV/tY8F/bKePtwrqV92nAYlC6oRZY+QkQhxaTqdEKg0G6jDU7bOxQbSHQ4
Sdmd3UBiqtaoOZpnwdw78QbVJvRj3Bh/UDtXJAI9qjbV+ZqWLFocTPUpDig33NJX
Q3c5fAG2Jt8zEKyML5xIOjX71MuqWHMj/rZKAQQRn2clQFF1Q2GF2gowt6Siid0K
3C9Xz+nxV/IMdtOuu5Jn+vqu6wt+iZMfGEqUPmoCshALrwFtsQPtzkzgHt+JWcBy
Qx08OlUsuyYUGH1u7O4EDMLbOi9ySDdWQjnAJ/HWpX7+Q8HlEw98lW8397ZZt2Vq
jq+PixxsJgiZz/WgFY0qTfq4QHeiYYjoIzYpxTWAw83BZ38topPzWxp2En0HdP5h
Fw3AcjzqeWF+ZjeY5XJLUz4niVrSEekYEYhvVruYnm8IDtBKSnCEuWUV0dugrUKh
AhIxLXIzJixRMG/AcbYtq/OhUzMUAZGcLmNyaJeHcqBkVbzy0mlfveuXwodaN0pz
9IBxLIGTQGU0CKE3JrposIVIwxyo7k01KQ1XRTz/qzJiVcLfLQ0oqeJwtE0oJKXr
fbQbauQgRuucICBfm8PxRgmmpWaXFMQ62723wUhJd2h6QCEojlU45HMLE/1X9LOG
RcheVWEEkj4pIIAzMb+3GeRwvSXW2wa9gxlM3o/LbQ8yiRts1ru7Tq6lx6zXpgXT
MHatBhUrTnHTasbq5BaQjuYFewGqmBfQhTOnnn10weJr2wbt5vJama5miCBql3NU
1kYmuuEVPyf2hrMcvs8yPB+IxWLL0YP3sm58ZHrhegBMlV1L3O6nLkhyFeqfElrh
SaUbJ59manF3ezrjpX48VcIgwAS0RxdvXnKSkBeXs3ax5X44ttOpH3kygcMwVspS
BWI4pW+OZxfrZRXDdvKDoolU2SZ03v1a8qXn3yHYY/mUyAyLU1Z3SeqEV3fPLWn6
r4MpAishSNUEk5+PKQ4DIQ18Ow2/FnYvKfjYD41tGkeBi4lLsmp/UiEaQ1Fil7SN
HSPlvBeYwHMlu2ULmOQbimuyUTfjhHdLGi4VYcA2vtBWcOYyztl/Olkw3hmGyEoD
RZemT5Bs9FC2W8VpfUS7F3Z2w81jnTcmz89o/oTRlIbl2X93+q13tCM4M/kcOydb
zSwwF+CabIIz9pGzvIo5aJnUwvemtSBot/uwPjRp6ItsL1rrHD9K0QxNZpnEPpB+
p8VB5/2n2lzmkQqr30mqyssJzuYWgG4YPK6U6duiHznleRIMHVQBf/0t3zozypra
WfU90nlNgeQ64b/8agdg6FL6bT2a/QwOs31/MTnsd5/o44dCxp0FlfsGhOyIfpSA
P26o9TPUtpHWRH30n/xDOpSOAF01w6pu4iQCx9sIqkhFdNDd7Wckra51JexReby8
T3JonDcxBvMJxaNBgTVKxZiC2JlJwo7N19NPcuCc/UuaXsyTHQPLQXb8WhPHgrnm
IpSzuFlbpF1bI8h/FYUuch5nd0h6yyHAz4WYavXUUfVNnrMI6JmHjOJWG30eILxk
EM/54JPRqFpgqGFg3991RwJLrlfc8FW0MWrNjAIueWefVtx5oWKde7sIdgihpSDl
SpEEjamD6FbksfNMrLEbbClvwCjdtIDLZv8JzoUGdlRQj3eCEV5e4KNdAgG9lucm
qdPgmX2fdn33owvOJVXVxox0KLy67DASwZUM29+J9vnqZlkjFAYSgqljjC87hJef
eWqvCaup0Kj1RvZtWyUbQchI7tgcQfH89iswTDyHTTMR+01t/l5p3MIldcimUQ40
jtaJrocFVe5X4c0pd8i8MDecXmgvuoKTNsyAlhrw1dgDqDJx2JrS3LcqtofxLmrt
y89vXKEFBXX/F98zJScccYVlzz/y+igRPntqYT9KsIzbKi4lvsyXY5pcUaPjaIm/
SL6SU226A6n1mYFdKjcMj0kODlT3ahWoseDboGkJdSkZUnic615BOI5fHbETHHaL
3hKR2Y9rRKZtnMgYiuk/0vHm6I3AskYnnPfF8xY5fHuB2/DQH6TVjHXwYbWmCUTo
v98DKvs6K8LJ6Wa2VfCVHRbyf9zEDbpr9CLd+9lobxg=
`protect END_PROTECTED
