`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HPyr9aSB5UVW/LU34cLrUazcNQI1LB4JlsQ8xsHLuavBlZ1tzdSVPEsQoZ7qWI3B
EmG3GUT7SHfheitnZViTqq+TXwvnMCdWQQ4bn7S7FevHwZ5tsY1VMBYeNs7f7rC1
yau39eNBHiT7dEeOnJPy/1l73PKvJ5NgvhU8HEOAc/LgqFLmI1JMgTFN99WUJlDD
vZsCK5WlkpoHS475drqJhTrW8IcTsQB3Cjq77irmKzVmxNrUsMZjxCLJ/XCc61RI
W43+yE5xVhId2voSjo+dpBkx9/tokT27LtnDnmUZ/aEzMANEUuLfhnyv4sQWD/dt
jzvgmKpdxGPleHnbjdEss3rIY38DoDEHtYl+1uoCCSPOYHJXSqF6phIpTqV2/6Iv
gsh0BBybB2tiPsC5cXm/jxp8UesNZSa8XTPuCT8PCzyyjOlW7KeDWRMVkT7IV5P2
nwXgZUs4361T5t+1kxzwM01nPJBrCUQXEJFZRfqa+EObciJv5MrBkZXEuxSLkRHT
F4mrOd93jp/mNvA1rtQ/1zskL1ZzTNUkafZpFpTO/BusjKxeAJiC7tWv8Iht8RcS
PnKlczBCWUOofoMIVvFteXtuzZXpP1Ia8u4nPjf9mHDLlQKAW5KfQKZC8ECj1+DW
iSli+WajKhhWZNM1gNprUK0irZ2Ri95qHUCg0Xjh7cssECI4HE7pEVik9moOHm3h
O9ekS6tpDh0saPC1C0VRsGl7pyMCTCIjMMbfvP2bnoxoTiE1k+quFTwKZ+KIJPbd
4X7CtX1ku4s7FH+OrcfeqvmfRVU2wHSoYubyGc2rHKqSAk5p3Z8kE7TbA+B/WpME
R3QVL2nM3Vk0Bqbq+KDYO7ji6kx7WCeTrU7suxtf1EhYNsHXyx82idi3sElkxCBc
EN6ZiVn4EO9ZUi71kFfpdwvfeWjnSrNjX97xZUN6PSs01a2sLMNl36c7sHfgVVe4
nr9VeJdTxnCqDOU0A6AbDTHEIzqvPCzhpoX2pCBEgynw6WKdFkDgaQU8zzIRGs9C
jEkHyjlonBphahDKyO3T/0dGHUSEquzEe+4xoZhRHVGNFpBA1rlK654ZVpn9RWHF
zayIStLxhgXhaTduCpKwsAC2jLK7Fjh5/j0SyWoQ8E9Y4AIypC4atpf4I63bBzlR
C1+3kPbNWK3u617sQQG7msTvastNKGPnEw0v2RJboUpc58UnUe3GdfJzOOi/kDLQ
HPFoYCC0tSzToAfFSjiQwV70nAQNL9a9IdaDSbO1PbCqPJb0R9mKDEcURJKUrzv8
bCPsSLsz0K3xSp+dgrCXXHV27VamVsgf2DqS83nB9/zhd1lr+ayKsCn5agmwX/W1
OGtyf1xFA9zUdb/G3ghJSLyHgobS/IU5gZjgNBZrwlkRtOp6gtaAKdUDNgJAskXe
Ds6ZD173O0Yb4vPEyVNr6DVxLutmGBsS5DwKxC6tcHm0U0C62Cy2yzbS0gM5ldO4
uOhXLfwHByg9PoyrVg7dQOaqjTDxtVB+/19yfyaJaDuPr4vlxP30fv9OypdH40vB
oFx/OzpZg0Q6wLOmivARp3AlG3kX13JghlglLzUU/iOeUa/3S2VGraPuAUJiTAAY
bpcsPUC0a2LGRV6Gv4BmedOFx/hyUQMuLvpjsVgFrFO+wawtWBhb2337G5VpeXCZ
4dLN5/T6bBwAYWgIoPWsH7/aNxhzhfIRuUyJAGr9b0VjFLlb/tmYGc5gneVx9ich
OB7i+m6ErECuvcwyZ8EYARoWKpcwqZC/O4Zb5HKNuQuxGimYSQZYbbhZWh+cB1+B
hazr3+kqX179ut4P9rMKImMyRMMF6knEkeCuyYYExpT/ccd1izyY4RHhnhJdnaU5
gRaOEmUpr5qtdZqf1z+MeXpcnsEnBkdo2qVzi+mgfMAOjblZp2aQgRNgrkIk7xXX
a4J8i/AdwtpYnvHQw3BpO+RF3nI0neacUcvj0b+tVI14RytnyPDivxGrAuZT/EfU
w3UcesBdz7AFPiZckEwOQZdui1ZZZbQPtz63m1feg3viys9RvtARhWxLBvjFlmwS
tPujeTpOMnLWzsvnxU0ctGFwNkdLWKh/AAbHnK8mk3Ql18Dr2zf7D72CriFI5Gdc
dQ7XpNxiqRIU9m64UqRVMEZxvC8nS4eNhKfrjvMOndZlcBk+sxqYVkJ4p32ynvpm
fiCxSXC3HryUpl1CnPsKUf9qpt2HOLVUmUScKCq+qNDHNGC/5utPoKBQLXXYmEHe
SJQH47UozKH6+rskhOVIWPMWb3DmXZtxxN+pJiuCQbzLHyX9AUzmuPe98RAavu3A
0qR87xxLdQoMBJIWpgMJzPdLqPfFSnCZMfNuVNC+0ixbtYSYcmwhAZrXHB2o3FPx
IQ4ipJnb0s/Ra2/V/uhFYAbQai0XYyvQghxdCZCcThqKp2P+VgaNub9M5xX0IW5w
dXy6Vq3efiUhAtz2FjfSVQNHK+k4uG9p8zzKxmjFZnlxeTknrdf54tkaD2ybp0oQ
ZjqyXAzN36S92V/qXIlw5FJmcePGvEaneCgBNTMZ5HRs92EGE+KokVjNrDs6SJcf
YzwXW4Qw281XPYfxbcNRba9G73hpFm2iOFOsuHv37GEEcG4tjTD4Ctr+G/+MYkX3
13X5Wnjc3xJFQucb16TaDvkqPlFu0D7D0SvQTV46EJyRLKrk5NMz3LbZhM8TBUKN
hn+Iu/aayy+UGPDOTQ+gW+enAgVZkYdbRrnlnG5kGnUaePjAasvsyDBAbRH75E8/
j4ThTXZxr/WwRvzapSz/dDlcPi5a+lfOP/VZmfABD8x3SjenxF2GQidM5iajRqKE
XzZWC6Ehs3T7f2972NiLZvA+NYCYZZVSrKXdpXGfNfJ2Wnxto9YM0objzjalwDOM
fzAyYwUcKaXgf6StzmaDRZNw0v5H9g7mGYNKpSAZVJnNKPDBKjHRTCx6qKFfUN5h
GopAca9fL7AN/WW2W0Gjv+F4dojzxXvzVG5ft9JKtK6rg36C1s6gQy2K5BFGwt+Y
Ib+T3MXicGajrR5TIJwjEUaKUc1MemApARN48scm0lsOCYfcWnXNYJHup/UQWHWp
Nqsw+5CD6olkMCC0DGO0JUlysN4pmBMs0TL0K4FkyWfclyaipajQBXq2UO6LcBIN
YFtOVZK1v5kK3b9vgjHyYkqBeQirq4cqCLAYBmsSz+fbqdzmw2IkrAnRzRF7XBPV
Dwyb/dCf/ztyOoHzpdpwEJPco58PFnI7d0d0p7wddfE6xTddJQspcEsM0RnNfZsh
IfAeMWOsdIQUV66KmxO8rWfYHnNsn1sXtH0O0WjUfhMvXIKvpQ4ViYWXJK/Y6pN5
iPKCB4uF2UfKX9KpjylD0BGYpT89jaOFkW1bBKpX3fo=
`protect END_PROTECTED
