`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GRam00Vz+mJW3ZSaN3xgImyv9/7tHzFI1fcWydBjvx7ENWX2BbF6FxcKXdt3wmr
hwQBCrda9J+eoTbpG9EGDGmbLSBcHe5t1mFl4zbJ6w/0E6bH3jjm+ro6JKzfD3v3
K6tSZU4Df9mBR36iAPge038LEkQEaeQ4zUkwowoTHpbiLRKs2r9NG7LWwPkhCiyU
xGQpdaz8whKSy9380AYSbOWd3uDka33wieX3bkX1kzJsutI1KY/RWWQQWz2o2rLO
/oVuRP1KSbvZanw8b9dWvUDKofo/NLo2iixh/Ubq5KBd+GxWClRWu9+4TztzX+Wy
Bht3310dVTdiQbQTfwixOH0oP67h+2/C4zi+VJW8uYmCXUhsFcDEDyuuV+eHj+Bl
74tTbYlr0YVu5fk2jnteLyP+FHtIFNda3BOBvgMWU4YXWea9J7ffnlHsG5uSmPku
pbtdjwSPM4Xf4DILWq1FQgawR9UA7pOUsE5sOfY98+9inRZpzPMS7hF+kLl5igvr
5sWSwuofnsqAt+csX+xLSpsoEWTqYrJEIGXVWPv1+jZk59wciANDRU5MBLsZCZNS
aPfhSppP8H+kez1IEhco3oOWX28rO0j0B87aL6yYur4CThhIWmVJLh9JIYNnXGUN
CzjiJqrJVyM0IVwEaZj0/bpObLCyZAWOO5dEWzNKWlCa+Yz4/NHy8gzqY4LFH4z5
DOXn21C83dGAln+mw1Rg10KgmVU7jEQxpEHIfJjs1MMf+mcFW4Blxad0xJ+VQNZS
xDHMN8mB4T77zad/tGGzXUHp7j1Qn+5DuWIEs5x/iJSllFHuRhVtJHjwctCdutlX
CpY7d3omiL/H9FmTu+GyvedH+8PM2V7Uwce9UqkfmKj9auiY8PRvNE0scv2st0Ao
lQ3Z4MO+mdTuu+UcsRJcVTkRqDh4twFIN3Ga+sprcfpFSdlFJ24QEMmfbXNeurn/
P3V9E3wdJGDEyw7lHxg/z7l1JCNmozVfjVLdVLJ5EYxcHdK9jd2mWQFRXGrjksUY
fjeQMV+CpClRLHW0/RuRsyEG78222EKpJfdcUMACePqv4oLyrEFKi69P6R2wRZ3O
Urq4QB4ztjXXVV4spEPtVKdBhHE5BOrqPU+DQwLCE7ofCSzqRA2Ldmfrs8/JBn3m
phKC8e2KzLrmyXoU4fFXoJkubaHz0e0temQZpIfzDs0lJdptN7HAqYm7S2PiKLkI
7J11oCwE4/O+CH3J0hts4j3AQr8MlC/Xo8yRgHqljjtHZ+8dDRzL8RTst25Eiurt
p3J3uqpZGGOFZyOGgT9xmLUvVaoKIwdaJTZ6/7aPxQaPjMxgmysyrOtf4SNK7PWZ
4njYgO4M1/SidNx5NdyOUnA+R0lIGo66MiVsqfGtjLqUyZyepht+3npwgyoKNDud
MZQyuR9sgnEfViEpBDw5BAiFlJ5Z6lese7hDT94lROgb9n/GwkzvMEtdAEX/Tkzq
5pZp12vgiQHPoQpZ+TJqLv3Rx8qpWRNPAAri9XTwxOkG8cudfNJanNTysckan6Qo
Wx69ciMIeiirR0/Ie6VBZh6kQQUnDlMJ+qvoDnzLSjwGcM3gi8SCMeRS2J85OY7+
rT0SjAc4qcrZE7cgDRZV0AFcKkujale33mt9PT/FKQU2E9CD1mTGFwPYzhecYWWL
5s55IyqRcI8/uda2tV/2RXMzWA0FgzebSfptMRagtxu9vo2ETqdXsbp0hQEymMKa
6TD4ovYmadLLou8uwIFGaKoAiHUgXfq7Z5X/KBtaTX10g3dbic2DDZ5X9OOhbEd5
1r2HkyWPFWtKuZzMHDBWJOf86+IGqzlL5FC+dRALE7i+3oh1CaO0IKRgwfTlvvor
WvzfZ2EVREdOSOkwWdi0NCOI4RSqn+tOaFgwXmU94hU4IlSjWPX8dyAhrzl6HkPr
RX+cqYh7mMf55vFQmebhIASw/KBfIPFbGVSTRYtCzGymce8PpSWIk2s9/hFhs2Ji
dhXm549WtGs2iXGyGHD9NeunAkvqaZZj87rF0k4MxNlSwxMnpqW0jc0XwIttnlk7
mTLTC5OdL3ydZGBUu+Uo4nJPSXPE2Lln5QWyI5MLmRat23VRYV0KUD76ddwDRBbf
y7+1lsuhHxLCGvm7pV1J97bolkMR4Vx3JE5lHrfTKUQ/zX+e/W3CslOZUCW3a+k+
Zwq/7qpG4SvJ4nyKxwzE5QrbNMwlayebQTmIHTEfHkI/ZQzi//dIbmRoYBNztim8
zOzulfEDjrIDEcOuZI/rdZn9lu4xDfOpPBBCkhiwLodZx5/8NxKNcul35wBhUpfL
4eBTddMjBSu05NzC/I5bhsQyzkCubw0tVJ3VjCEY/e97IntwU9guVFenPCD9ZzAc
E+kQVQ0Eju75q0G2myfsQGLRBzjwueXSW45A8W6ZhQB81KG9OfHpujkWajRKpAr5
mdHWcM73shINejcJvWi//uzIwDc40F0nW242dhjoD3FUxqxkLjFjMjheNB/nsHRj
bWX9/G/76aFkoo9Qw39rTYAMJBRH+4M3WZl8cXdu5OJZb4lt/n/RZqo1VedruYFK
ozAYLbASbFxpftabxopcq/8cA3qFNutby0/nL7jkkCpEpbHpYAYgMKnZBxsYcV8o
ToPaI7KD2sIZ9dsY5PSyOtpw9Wx2g5oL75g+CUeikFPrBnww/5OqsqkKUfpS1lbH
Yyp5OlnmQwo3M944AsoZEN5OPNSi3K8hlD9Sn50pfhBpGSsSoDmvv6S7/OmxCTud
xo4tObqNGFGCHBHajkD6lzLkbGBbR7ue9tG6J5NPI0r7HlejE19rTt4JElSjDUAM
9LBQ8TIuJrqrzUBXdTBnzHIDEJeHPlGnVfshInP3BrVvWCxOQTzLNkut7DU1wzXJ
44Wfg3QVnbIowoL4eS4qqTYITdfJoNPjiGiInUG6sKg8XOK8UIYjeC+FU36IfCsf
N7NNL6l3qTXOg+gzG3sMlbLUTi8rQpadEyg9+phk8/ZICfwCWZjBaT9mMQqp+pMa
`protect END_PROTECTED
