`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZHS342aEV3yWoyrzdX+nQ/QBQSH7mvVBU6hTlNPyrPuYl0aCO6UP3jDeFQbksGF
i1ruP19L/ulgF2LL74844Tb/tWzxmtEgHZl8CJ11s7VMb4XgIi3NaxylZFV/cbOF
SZYoJDN54W40YRRaUUq/FuOixthzS+tBaHxkHMeLDi7CcM8NUoqX5F8Xr3PhUGBB
TDgmm+pWX76kNrAP7YZT2kJ8NTJDhv1jqftbpmR4D3M2J5VemXwObQqtAczTKE9F
`protect END_PROTECTED
