`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHBCCQm2L0s5+g6KsoGpH9elvBjuUC9lK9q0WAmQKgM1vRNa+nIRJXvjVOuSfeef
oU0O44cqXEvn/WtSlubF+iHZkRXWXpGY/eF8WfYZNGq8W7Iam3p57obf9GAJvCI5
d1DgSmgspaNa3l6KOFZ8+8Y0TPhIY1OCGaXe7CcISt5b5mRDET6KpFshr5MtcrQt
FBxNb1+sDU2A4kDtlatz9NaWSHkK3jjLOL28Gz4dKGq9ouQX5VMKy4EW5QraPL/i
c1gSghXi3xTJqzRJ9F5FAErQxy3L1RBBmldhZTPJ//eXc6LP58PMHVuXGCrVbjXV
ecOuukp6pXp7mxdU5/xW3lah4gW/P6BFlrRyxftLAuswE9CQrLUM5DsC3bTRfpqz
Z0A9YYdXln3Lje49AFJ8zyvLhBpDNk20pmHNmuMGUWhpi59LBYRGpPr25WVJDcHl
DtlKTnGsplTH/j6pLFujjo45N9otajDMv0qY9fOFa/MMIm3kk9knjrh2+14XhFHe
FrRwwVp5OewbfdhD9/MKITomPwRNKSqlUAzfgGBkcElODVV9NQb+aKHijy17swFu
ak7dOpvKwwr1MKj7pKX73pvRZJ31hcxeUCPJs5YvxQ1X8ZPy1ZGT1wTjBlumVgiQ
OjIw1TejV73nlDLGh4l17ieRuTHh/LZ0YAnjkUVaHrGpIbw6dMrbZ9Pu27gyncNX
3pWz311v2l2sDizJJsHVU5U8ERoLdaQB+ikE646DEC56fDgtjmYRGT94eqJc65Ug
WnaO0AvEuXlMTmGY1quQm50NKdCF4qnlgGVaLXGCrTL1D/cXgbYIcNXa6xKrquA8
ZOvBhw5eiuJMQiPIYgqr3m0DtwIooLkanvi97f2Y0+bGY73ek2eJ+rifyCxsM1sf
0n2sqJ0lNTleYPeCfxkDS/Hl5/V6ENcUaR+WM5jXCZeWHCPHS9yt4C7LI6FoaLwE
5wK/xekYqx9K25hDnQSeCTw4xsCpRGoR9I8OTnulkoo+b4m7/N8pbe3CVsavtS9p
Ef98tJXVmvaZ6DCF9dAr+HHz/46fRFvycxktTiXlwsKn9dcq70uHfxkFZLpFufcD
ofLCTV+8o+4JkipmQoAoY+TYXZZVSDVqxohd375NCrvf68ZishL+1b/dmPPDdj7A
vo8J8zgO2rBlVXfdnq4xhQmwdQOfLqt19yl4Dsa63KnRbBnR8qzaWHy+jfoYfR+w
HQh8heGqb9vwA9vumGONNlp9vWXerYXg+X5RNABGHJK0IU+FCWdr0DOdwPScp2Dm
aZ0Yu/cf0e6nvOQyWsthjO5rG61SvqVZ/JBBulTfAF3GtTUbfk4XOVrIeaE2MEoo
kibJHslEHo6FMQWTKkk9+B6xEWLewnjSMON7BeE6fXKdfHCE5JLS6b+0Gk0cT6nR
pUnmyL1yQD8l08/tNdgy3VZRraNmobJmsYfP3qZQlRd8zfV59aEtXE7gJ1S91iWD
0EkWZ6ZWRCz1PkL5ppPIjj39vTE6jFb8UpVVvAScUiB88H8xyNHVT/CRaliFK3Vc
kPnrTFxGmidssEeSDQhE9SjADEQiDNXnaaw7lQVLWOxAo+TP4lhOnG6dlESYKHy5
PNlBcm/KvQJS6xm30Bl0G35tk22g05my/yQavm7i9KI754H9935Ybu9IJbgO0yf4
7JEk6Dc2JVoG5M8rL6HGShr/AOzcsQJCc0dJdN/hiVo9Iynunig3ZxGg7Eng0y5/
laIE2SNEUl9e5Z3OgQxPiCIICEmojUd5xbu5FmzhyUjVAp71aWC5xsr0MSRhHi0q
fSe/fj8yt7TrnHLoGZOI/jo5nVu1/MRF3enbQAG05zM15hjWoXS+TyT2LP3+sjCR
TNxE/aTra7bVeZauSscdGA==
`protect END_PROTECTED
