`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLOy0D9ZqeP5PmjmvxmFOhYn1HnqYCwQJFdzBpXzsre3oyb+6XTWwwQ3JRq3rWdj
r/4nmdRBTDz2HqspN+ZKBNy2axnUT5Gc9q1U9+OdqiUlU7Zq7Axap88VUWaEqgKR
AiyUN6pWsWDNl3y3kbxGt4R8ks7K0V9mObLFdEEckMUurL8AW6FH3jJUb3RUlGql
JmgIsBet7n0GDygZYZWoAT1z5/t5PwCqwq3JvflU06fjKZRnvUCQuhth1mLgTTES
A0tONne/yiI59OsXDfQzqoLHz0xd2zg9dB0A8LqlvgPR9b0erBye+A8Ra7SshVO9
iCneRNz1jzRPiv4vCM3+5xj/SE28JnkZh4+uUU+mn/hy8kQDEp90NWPgacRdkAJ/
vtS8slsAwkS3ESojblYPM9dwxOrkwwqGvXMWndwOTDK5MaLIvV6dUC3iJqAwdFBj
WtdvAqKSdCbRbK/Cjt3pyRWNMW3lTxkbRItZbsaZxzttReUolXunxcUS+opW7bN+
/zaRCPgBrU7jmCLdr8XbuwpS3DFavVXKqN/kgtlrn4z1UEUN57AwBMKsnoZHzuQT
Fh59yag4Zvu3FYauVlgjL5q+RWQNRtMAwHxCqQ5kKC0ci4SsAUdKg3lSqGYIXbBh
ChIto2/YRiqBUhHZWZOWuI6EvIJpg9JauaBc8EiQHw5wcTtpG3+BQslO5g6TkFFu
H8kqjGL41+iq4sNpdtPwoUuH/oPYsjAqFZoJoBEBtrKOZATvyrjkOzmIhfR9qra3
s3jlywKvtJKGZL3aH0bpG+wCpGEQk7R8NChbLTEmniFaPAhUPs1aFUUBjZW/RPTl
ehp605MdFTh8004nQRRh36ZM98vu+xSYNfcjErSsuqeAFbpekxwexaVFUgzmTERU
kykjnsS5mgyRWlb9oujmW+rEo3hbsILL7gUB1DGXbdwVmFj2bwNPWxcLxz3V93jt
KLL2X0eZBNy/fa+CPbx/Zm/ARj9mKtn0zwfKAskpVHLij9Vkw1PHvqTGLC4j8qea
Eph5WF/VWV5LqYaukw9M41xeFVoT3VZH+5obZTwIJ55fVmfh2ALeu1l63ndJF5FD
+diWRhZ7uSkRxM0magqd4GWTLlsvzmhxUpzN+g5dfnRK9J5fZvYrm+qXhhjBIeRc
R3uzcTmp9E8hzT1/YKIRTk6OWcBTGqRZvzDk0/ysbjGC/BgzhavTysV6GuPB8GHs
Bw29+Cc38b6nBjxgHYGuo2zEsZJtAGVQeUDT2IeROji7VSOAuyBPl6JBjshOvXyi
zzipX9xV9+Hi75XRK53Tf5GqheQs7cAQjocjwksSlY4jO6bXAv3g1mRcKZKgRsmE
GPVyOu/Z6j2E09tKm3x8kludL2JYpxZKpfH6IBV7wXB8guTSDm5EjO5uySEj+6Kg
wbx3vfUr0DOPRJSe7v6pcZOi2jmBIC9sR+S2w5Wyjig108gxoy+NtxRx5kqQfGos
mn5Q3BrJczkJbZ9NH8b+uIOONXjk+efkt2cGiJHuxaOrQN/ZOPtO7DFo72vDc7OQ
xyelAf1Y5D5atiRtHhTHHDVyU5HznaC/fcUhuyD56c/zk6ERZkDlMdqAwy3yPzXj
HtvO20/4azMxGmaqtsTVhOwf2BYzUA1+HZu0BPnN9Ep/U2VweJmJdnTVQxe1Q86R
57nOXX6nMUBe9OktgrzllzSVwuv5DFd9+42AzqXZj5eRggRMgVQ7hZ5x8psA4OlT
nBzPf9kU6uXzv4NrddmP9gzWJv4v6P3c1kUYO9cR6blf56cCIr2xUZh2UZqBn0ds
r3/r5N/dZLf/ql3zaFnCuWWO6LNx2hbjFy//9HwaRzvmz+NNiT4kIu5Q2hO8uX97
BSCrfhN8cu+70LhT6oNqYT1+Px+O4kFRTq/NWz/pRvC/bE0At/jiB1p9ZNxGK6D0
7n9xrhQOPPBkyy7rJWWR/4BWPj/zZyhZtRRPvtw/cmc3Koe7FkOL4fgQg10H75YY
fgZ25XWmNfYJqjeJQGQNbc1q28P9/FsxD3dqJW1kYRCQH+NbcPfSG24nx1EzSPKt
BBhSY+H1OaFugrt8Jzg5+XlPv3PCAHqNGr2RK+Yqif3kXAsYLA5II3nqNxHASHwR
mPZ47YLMCn2e4zb+g7c3+LSSG8r2vOg3H1mlrqSuTRuIIWGC2eMJ5AntAuJoq6M1
zpNLwYDIUtKUtPyWozpuydzADs4OvlsJWSA+lOIpY6ribLIUnZxE7o8NsQaE1mp9
hut2eRMy/YclXhkvScLhxXFxZ+zmgBwcisoK/pENpkBrDJtYuS4KysVnQCKGzh0/
NeUDnkNEdvGxpEIDkN1Teux94UbIYogAR00VPmNaEAqFo9fLY6v1IzltKFLa3YsX
w3Gy3Ak6Kys50zdMyGjafEuN2WyXUINEgiCbrhMMeL+uX06TD1xSMEQ1j65fi6MX
SjU0s7cc6M+Bc1oQG2OgxQ+t4U6UxKGja4lpK/N2jnR06UFo9WAe4exE3bDH1hac
2lHeM3SQPTFP+BcbtZyf9vXEOh2nY72O/1n3JuYj8su+t0kMhbAYKfv6L9vb2aaK
ckGRmUmsX0e7hU6IQfc+UE40TaZ7vzl6r5MtN1SmIeKIDctd+594ERLsAmdtMdqp
G5N61wd862/IISARBkvNKn9/eDTXoWhSQRC8NrXMnXgh1OySmGen8e0XiHJkqHRD
3deoruonebxoTy9HCu4vvEzWxMAsp/L3rKxID4t1k5dKxNeRNvzw5ZGuY9xFkMRG
Of5cDGl+S9B5G/Up6i+j6GfrCdbUx/riaPQG41NIX4mXqUlrEo4JnukY3SIPJWhn
LQf7AdjXCuqoHfawqgpk7HZDGZpXAp8L1KcRK4hmknuPL4tnycX/R2azFGgz/k0m
YiGjk12VamcWPLFSjzfvN+PmG7c7xjbKe0v81ZO04FikYONhBaTk4PfCQ/3UVwVQ
hq+5GjOzTpLwVtHjnXZ7m0E41q/6wa5qC4Fc5MiTN0b59P11pdR4XIzXrr1qNPlx
N31/CYIt9o9KbdqODe4oH0kZEyS2YzJm/itIU813lsvpI7XAFSnpqJp6zZF25yav
zdzQh+UxLFOj9xxgO3+VlFrzskJ1One8fbFDggdKtyde1xF7c0dk6LV2Zgmz44/p
PNI5U+kIlIWN1LbZltmhhIa4Rmsg9eTGDuAnGqow6ldrf2E91fCEmJEdNLO11Q5m
r1LbZhpmy5JmaZGUMuek5/j0j6CQIMMkLQ9La71timNB8HhIr75gL4rkmhslmSJm
gvNPh9vofYFYYdT9F5sBWAAKVRTzkRgtRISUm1VbC+FxkI0Nn2Bku6QxkU3zq9mi
T7fVPuRA2c9IpjWPRI3QS2QbLVnmPUqgy3BrvAaUP7HfBZmXkBdIdw6aWV2bSY1i
aGsk2gd35Ac8qsLHYVsEUKlavb3hP02s3eCUErT7VGRtWL/YPJFoNv9SbtfZiVmi
1AHs+JfkZ2fGqvHYK9oUdLFV+WcoeF5QNYwSTRNFXCg6qpqEo9kFXCZjMgJ9YY05
8kJhbGRAIEaQNLdRjJMHLS4ANKJxBa7iKWIN4RESU5FdAyLTmrwszXVckChKeEV7
5jT8OdiqMix9PglL4jvXPggYJwXN/IYKLWYjorBksZ8UqpGv/5JcEdzm5qfCCTUm
Hr/15WNPVLEcdAFr6c1aKhui6TkpJBl6EjZ/xYaqWFy1eGi3eEgxo5hn1rJ4cs2+
ROZF1zUYkwovhi/CkKsd8SphuWtTo0Os5RerHVK5ksXfp+VWB/5zVxlO+cnzS2sT
vs5FR2I6p2v9Za53A5o76KpIfLNqHtWTPZxOUD9RbpXZJuduKiOe+Ipr3/t8rG2Q
blOW/ZgpmRqzLrqf9ynkhseBSpA1/dz2opsFDFqemW17mlluH0Ka/xdUpmnDuTx5
YiLbxToQQXq3eQNb5PgAl0EpyxMjKOvbypT9BhfVBy7ors2t+jL6EF7Dlcp4+ZU5
k+y4Q0QFal3TqsOs6dMe9tzn7lkoIqmHAZI97rYMU5uCps3Cg2Bz1hUdAKHMozBd
441GuAmcIY0zaOORxAokb5HhPDDyUYymQSVPDhqWqUO4nbbKSD+sgKM3EoXLAGEX
74qWWEfwkrzSegIM6Sn+PoaSsdMjMZQkJgIU/4+3748bzWCcYrqZRvNV0mz0VIVc
3+4ovp0IJFG7jHOqFYQYtjDRDVUyBvgHgiCgYs0Ah5Rywh69y0YlAP2GbNXOtiKz
8t2JtbrVK7MMf9B8Tv/hXrJLGnz8KTAgq+4grA7W4+rg/vfapliHSCLuQtUhB7y5
`protect END_PROTECTED
