`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tKQ/k0LYuYzT4kIefH432bF8dA5eGq1QH4wHfmQCjLLEEo+hS8Gl5KGox96rBXJ3
GTOKr2ptJdVWJy7VQSbnjDhemdCw6h2RYsNVh2EG1PAXAKVh7w+GnCYTHx31iI2f
LaBVujTU0E6S/ilIPJMuXcr3hNJMQuKiHDUksKP8JGvrR7txGJ//Fanv8cRxunHu
6BGKsZUsVC/ZyGWpSG18LBufLBqk2edwFsCxU7GQfr0vrWZqUMeiRhy5zukylf0G
vOsaMJztK846ETRGXw29lYLDhQ8MBCEIIrg2CFR0/JUewS9yi629utNLy6PFq8Y2
LcdSGR6z8CaCBdxNo5Rt8v+vuYGB8oX3F/Y4GUABGeM+EjavFM8URcctHLwo4ElN
Er4ToNHpNiXxmXcqkzsOut2wAZH/goX8CkNxIs9CLsL8uUUVtJQovZil97k7vvEL
4gnqsPqNKMeWsYISG9UcI4tRTsX9uy71OiF8ufNNwKnqyaA3MYlg5Y9+RIus6GoI
JpLw5RhN0+hVG97aoHDd9+l3Tr0sL7Iehx0oUDWzghj/LNgBa90fMCBkLsH8hPyI
ZV2yr8HHGGZNZLafeC4dk2rHwPJ4PINwLtC0V6ulUToMDhzTj3MBZPgy6Juew0cV
66gvXxUVPRGkwqJyABfbooFGO94YxMMXDowdlIkcWcQaMHDeHHX3T+jKYCNWs5jf
7t0lbgr/xX4hzYE172Hp/nuCRhGrVNxyekI/u3b69Kmo4Mh4319pue1M3If9VNn9
8GxdA6h/Vlv0hTUt21rE9pdiDeDcV2YHwORbAOd57KWj1LE8Nwnq5UDJy6bwung2
N6KohMpKdI62gcWcQSTbihlOxDUAchiF5ti6nuTagGiSCd3Csoyu1HggspvxJnCk
ewv8t9u7iJygoOBDyxLTpnIACBnoJWa3LusTp79juAfdaG0R8qEVyyU4ryIfMLgj
b3QIXV6N3PnSoFyNihetdVlD2HvXqo6sKGp8bzx6g30zeyDSkNK6f3vibdr6d1P8
a1sDAHdvIpBIPRcImvRlG7LSG+Y6fM2wkvJF/HWMM0YCwxGkoQZMEXLv3L4zDf9p
aljXOrx1YQ+gh2igJB+HYcWKJY1FfMvqcUdgbVaPOz1n7PMiy9SFxTIJTB2g144+
k5MzAFu0ImYEYli8opEmyuuzC3keBogEtRBh2qinVtztKEJkXrITmYlOi1zvDaPY
4bS+en6+EqXPaYOMaX71Q4ZBq7x32K6OyWq0OjixbVfKvDS+NpY4/6iGDpp5xW6i
hsyoxSmPi81WLDUCS8O5YMCXCwYn030ZLR1ByDx6bnQ=
`protect END_PROTECTED
