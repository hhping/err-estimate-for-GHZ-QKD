`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hC8WNRTTDbmdat+G37QOUd1LAh/WuMog0e3Z8Ltl9eemiCYmhD3pb/LCZmyo6Qd2
eRGJ959cQcjaF45DuBvkgdJRFIeKCTD+gVmBcaEsPfxRPHYZfcAgL9lOHC9maxUp
44Ou+QF3VUu56CQ5VnsfspHZkvKzdu2D3fCOSa6xDmT5JADI7ycv8P/+SB6s/PcI
lRXu8K2+xJbY5D0+upF6WseHOd8l/5w2BRKmEJri+fah33/HMRslsOKDF1XkyVMq
NUa9WiPBe1t+vlkwfiydzxj9fW/VVh846OM0kGl0/FKgPnZngIJeKl5Of6Y0xtf7
sf9XR/9zfcT4yE4sZfMv0sCgSPoF5aSdk9hLrud5x+30LnRI7z3KTsXmORuugXtV
/iGG5DbkBG0GTeZ7NtlU6I+JDEwfzvTX76HDirq6U6M+PlgCo/igsRedUIu/pdVH
gypug8KNb7SEQt1Ov9/CW9PTvtpuRRF6O0dycl+McovK88Mrfqe8LbzCSkugHhXF
MA4lAuKZwvgMUXBgg76Ant/n9Q6di40OWdJWgW2I15iV5KTJCtfg1hrSHeZFtH52
K2Ra6JlIuAZvr6OzDv8qKB2vamry1aIGQbHSi5NSENSLMQSjWZrlbwhqsPmCLOO7
CdbG++ETiTJ61Iyr0BwHpMhEZFLYH+jo/k2ngcD4BCl30kvKyt8FZJC8oBioivF5
HaC7FojZU9pgNNVntwX8Ze3rZzIUV45n58PGJV/F4YF9BRbv0Lmge7JxyTxJwCfL
MQNcPNgi742Wll6j7sWuSQzmHhzF05QJsaa+Tzx2hbS/g6vQXAQ/XOukEVykp8X0
dfL9jYyD+qF008JCOjPZp/zILNHihaS1jzydiqnPIDpf8m5ne76RkZhpMt3bQhef
UZ8NgZSbiTE2xCGhbdqIJ+pnOg6cbcyMPaz25STAqcu6pukDQZ5YELM6Ezk3h8Dn
VYjfxEHSsLjcA3thf+ArpCfG/UgLa6GaJlyvSHC6+dDrjgDSKIBuiFNImKROksKZ
efbXMSu/j1OjFlfF2uV0F3Muhc0dNg35JdJCFw1hrgqi571wSuetpEnxFYjc6u/l
1WmFlkobvYUd5mbMxv00zL6f+c1t/OxvtelYhKA3vaTS0NjJ4r8/CMXl/Eds7stD
YAKJSfXYt2x80jBhqTPNdDMBS+EY8NRUI9+O2oTUdsupvQLkUdc9KVlfiRIyzpwI
WFnSiIOvLrbSX6aR1YAbBY4dITZImvBdeziGosw/kkzVlHf4sYT9Zf5isoMeX46L
fDnXshZl1NRlJEnON7+9V1NymT6UHT22uWnSyFlh4fI2nkQOEjgzcWWApK1RO9hA
sn+jy92bSkthumPjNWo3MYJ3LH1hnSBfNHxceocpXHbEDne94F0hxMt5040mlctj
xgjKYeyIr6HimdZVB3hZ+ayFljGIpMU+V4NEh/hW4GdpbMgu0wv4NUM/JSbHhiLO
rowteZIEWsKXzLPkYF8aY92ajv0gAeIMMuy2cWDgtO2sBdT/rhQKx+XDpx9cUmHG
LnlDB7Uf8qaoIyd6WvQ2m6kBWOBmmg63mMI+99fsQ8V0w3Egz2KWD1x8/0qxaNgk
+/3EWLJnHwfeUqpq3biLHS4sx5E6jIqUuz5rhPYLWjmZ09+0MEnp+bwBAZ/E3d+T
4qwees92Dldx1dXhc/PkSHD6h3VWIEEgR2vRjHjyL6nB/vbH/vkAw/W/TcGPj5Hr
3S6L2kDNekcMTb8KZ/8nEBo2VjaH633duhtjVbecrkqYlBI7itfiBbQlt04nNonj
e+ll1GW+ndZVWFUEfbEiV1j+7SSYyBY/+Oiv6MtHUf7WNX9ZhZQh2BWKMjyKcFvZ
IVatDtwg7LkGkPett4D878zmBBeirSzChWgEQY/ewUQkaQW8Ba8Hzh+GR7Q4hUjS
Wf3KOH+w2MVMHezBX8zysvjgoNU61f+OxgwZdU1sDkziPOnjtI9A4U0wZonepuFI
RQx+CNW4Lp+xsrnbdrht8edt8qkRWPJiZjQi1wHxl/Al2OEtWyyZ9JvY+J2xWtU6
0P4XSLTXRZ34oLD4zuG2kn4TS9/lgUNJcMngZtwmSigADGBfJqOb6c3Jc5JZH5hA
nSyCDCW+1U/jqNZ1GTLTixCmM5DAYnKnef7k6ArOw2Iiix9efo5pux4IaMwYDD34
Y4SvIy+O9uxCgxfd/wz3Xb5OBWiLXH76kPNLsgPx8DkPam/j4tr/ipLowWtEluE8
5Ib8236OTu9o03z2K+saKIJ1XLdoK2RlKzlmBm3wyibHIl26DCTUheSrctjzZJnO
2WpjM11t8wIHgXB6bIS7aJmboKG1q549N2OiQUY0HcYPWDt3Y3ewuTqNbGE9lCcG
fLTYDthsCGcgLHJtA4w0+vKkMQaJTbtTVI7lWdgRHTT12yYCMvoyk5eXLWO8rOfV
OvlNNo7ojIQFMpXFfZh9tAUewmtKZ45d0qrN5vdG9igOp9KUsFzYuZ/TxFgBrWv5
dOGhVWhBpLEtcX/Kn7e/zs2+1o+u6V8BztCKU72PKgAsKmI9QWj2wYFS3EWXYqnv
CRiJgCmk0VfkE4QxAsf9k44Z6nSRtbouNTUp77RHALHTKaEIXVBpoEYN3mL6Oqcw
sqXRG0C9p+lcV4BmIKzbxclTMXzImL4gjwwyExXXdVrQVdxDDIZjDr35hdGvqqeO
85yeJ9zS2FVPJu/PZeUSH5r0UT+z6HAvjP8yFOfuVSQ=
`protect END_PROTECTED
