`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIaps8PWw92vGFLz1U8IDabKk8vly7Z0gQQC48Nq6z8+72SS2BKXInfE7glIJGHL
N/LynDXbJ8WnvOWAn+ZpGIxJi0vZzOtP/uhX1XL4nCWdsNbjHONowOUDKd+k5SuP
c9oJGzcRhbgYyiExzyZkIFD8lKXlfvlKJnUq71sLQ18ZZ7vVzpZb/pXFh0B7p3QV
sgSP4oJtTqSeUB1sEn3zG4CViQxCFA6tGy982gbgkJPbgCyaOOYv72o5nnQ1iA/a
9vEoFPxvEyY2uzparRGaxTXaE5S7Dvev2g0VkROSxv42DJ+3WfWdUr/DekasQKtT
6GLXycUjj1/LDgkS2KBYYMOPv8QmfZPFfnv4DvgWdn11NPFmUxGUJCwmuMu9nysC
sGMdpnBQ6dD2+KkNYeqCJgQu/E4I9sbGfif183/j0ZbEBrSx/8bPcV3jJiXKWJv+
i9tCPpRNBTNKXAVvnj3ii4C6WuG+wxyJyWFda/dJinCPVAQOpy6DD07tssisTlao
JMYBIY+DMVTzHAt5VHXRzTHIoD4zOhzJn4Fc+7qAMbN5+K4dl5d0w+6W6qCTduwv
ZOFr6QaZ43H70D9c7FC4V12lCP7wIOXngyNQc3bLgTbZTSZEnsa3WWVSorWwVWto
VEejWZg6aqWT7t+lasJOR93uX9k1h/c+1Ckn4n7tU720GSepx/ipmRqHFScrDLeP
Aj/aqsIhEOpPIJl+Xeq4oBpwg0otpH79hmfa9nba5ZrLzZ5ZKLl5zdhNupuTMcAA
+NYsDhuutEfbWKMQ5stKjF/kVK8w4OwtUXf4gz/HXxogBIiGOIlEBiuRQjKs4/Ke
`protect END_PROTECTED
