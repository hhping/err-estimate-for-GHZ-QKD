`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUbR/yM+o2RfDlUYT2CRrQF+67YL5th6r7EAci7AgXT0TBvdE3vew1UYrflI6Y9N
j+zedgbUGn69AAfsASWl7qHiTNpcCftWu5QaKJ3ECE+SfmMOvdIk+fx98l1sNITQ
nWy7Mu8GoWmEbyZ0adoCFIPWd1BeMZC/Gw309bu1Zj3FOmyIWIrN7lSWvncI5Uwu
5ESqXy5OGCzmokNIMIbERt/JCfXfz8DWIXqJmIMhLiXEMWWG8ZrquyhK/qV+LJa+
ATYF6HfgZIaA0ahI0VWGXizLQdlFp4VWjnXWqt/NULrQ1648aiairyr0R7KmzCYs
Pj/dWOBqPYFoTlfiY9GjavWNXGVgcBh8sG3zm5IT8wBKF6rEPbv6xnqe+nqXSW47
8+Y4qSEr5JC4rdZBC9l8oaeePSaxxlkIR1X1ru19aN81s6WJRax4rWy6JBI6CsMw
Jr8l1BM8WZ9SKCZ6eZvFtuEPRoG7y7MVGYdmRGfhlx8byxeJm71xmho4eAeTp/0W
nDj0K+pxdWr6ABTsz2ETwqWrjH+66goyJVsMEJiubKPDTfdmZgV8a6rlPPYJAXLU
wmlU0J17/E/SfVeK6XeUta0abCPzA46R0cs5o+rR8uW7BYJmVhadXZHdi8nNcdVT
SgMkntrlYaiXRkzJjfSI3rz9szzH7B/pOmQCVYau3FigxGG9U50fCsrqgAS9XAuh
nsfujFDp0hchWSMnH5LtAB7cOOALBTV1Z07jUt8CvVGe1P2uKj2fvLjgOAtWeIDp
bMAh+nUAGhhrO1FuwVa/yApz+SsS0sjhnpoF8p5aFWwHhJlyrpCLOk9tVNWzvPzt
`protect END_PROTECTED
