`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7T6bdwGZJlJZjWjI/e0IsTtW9JHoK0bqmf7761P9H90jPXfEz5mTo63icTfCaZD
ZS0MuIwD4knLT1TAzD1M3bTl6vNZXVa7xf3lpoF+43xmHKfTfMrON/k8z+cRVHJ9
CE3DrHnv9BT1AVFZe2+SMe0mfmBvqvYP9Fjurammm9/cHDrxQlaVkWQBm3p9yjdY
W1uuXbcU+dbkDQmP3TT9MtZ93vzoHS4kzCpxk/HchD2DkQQrPAtl2gdGgR/TcC1b
oOHHYO4OFgNmYuoxKEGiQLwsQtTPpE/Se1NHXTntCx9w0LI/khD00Cuqg/anh1hd
l973GhlbzLM51w/3TROD+bexxr+fhCXONcMyMDLkdIjvUvb4Vn2C4lm+FSNlOYxW
bidBRxFqk3nIQNXR2NgiqMU8Hb1f07oEswlfDMhoWmdg2AUz9XJzw7OAntd9RM92
J8WQ0iH7r/TYCokC5N1Z5IIspNl17BcFCZXwygOuq0zYf2PVgWbTouZ2PdCMYPy4
IJxkFrliLnu67AX59cqZ9XbiHlY+QlqWuL7SMboHqkPGwIUFMhq2dOVfaMH5oqFD
O8jjpIQdfzun8PF/m/Naq7zwkvIj7b5EpfPjrgK7OyM3dBCB0rsu2eEkGpQ/yftc
qkW7sRJkqppWql3RyzSGZPyti9g3nif54STzuGYQ/Yl6umDIkGbKZm92qx9FnEQh
5dogz33954VXOvvkyJI0X2WbFdTYJQ/ZwhETXjQiXxkXakU9i2Ldx/S1SWOE7/eX
mICv/3LWB8HCVjGDYw1EdXJdbppLWMaiQNPD9LRbF+oTZY4/B6ePU/0vthMLCt+T
ynCPS8Ljz5+q1M5QirpLGKdtScGEbew3XLHqg4uP2quP9F7IIL1E/d5XCLFrpCf5
mnrRDLQT9S2TFiShRgSoxtooPXX/stg/I721nttp5AVREXAsQKhx7HVCOlO3f5Vc
7dheqKMBU7R308nVkO4YIe5P6DKOmxfWbo0LoPz9GaSC5ZGgfEJ1rltwxddzCCze
IJI98visJl8fwyZfgM4697N38UcYy+/b393mRtjEiDyk500AM5oecR2rC0kG8dDh
F8T9PixhxrMRfqGMVmxscmrfU0Y8FTg5b3HVKzGWLvDZAlnhYfZQxvEwJ5g0bq9q
0jmoafHq673Yr4zbQNOw4izCR6u3o7IK4s7MDPUA6JOgdOPOSk5u5zV5pDOzvTwn
pHSR7Y3cQYmtpbaVCl0MjAmsvChaS1H1zYY6+MWc83UBpqBCBzr8VYJFQK7cZV+7
wkQcrCUX8y37P23on5tD+1sC35wf+bcgooaUxqVB7rYG8Z+NEl6kk/54bQ7Hd43L
MotJD7cVMn4W3tqJZFi0MfYeT/ct3ImFhDpfxXRJ0RAYIY4sNyzpEGV18+LGyVj9
wtWT59Z8ugX+RLDxHE3OvsXYBPjLkW46Z5W+4BoK8CBptYnbcLVs4VELmP1093uA
DtJ6lJWG6sp2xeLcZXFBhtQgu/wz3RMolnM12x4UqzTd2eyOQzUub3EVCdGDsF0S
VX1vv3iu5BCi9mG1D6s7MKxJuP530U38gJ1HOrNk1FoKTR9XaHyVi7cdZt2OgtiW
nqpHTmqSVUNzVXPS2AwWy/5SfAITjbxZvzMh1ytMhHTdfZz+fGhtldE+Qf5u5tui
SghYLb0ad6nnIURvBooQJ8yLkovDqFtWda9/+8BMcHWZ6Kv46OLS1YCXdtu1PehW
WDHG2d6hTBuzvKYmYeMNFYE/hwU9qyefJLvUSQbfIaC1kLxUX8WGAEpDaAjyrM+x
1eTDxCNXO1UGtvu7b+9IMsmM0IQgmBCbW35c25YsrhwOwCxGmO7nTpWoXIxKNmK9
suniqgj9S/iJ+zkhhZwqDQJYyCDhDxaX67InT8GQ5ba7SAXoVZf5/ShniByZPt2T
eJpvd7GANCJDZV55Ew0yJLPQrM4XLNJIB22xGk8G6HerIzJDkevt5zHhQ0STCiRh
cnfLI8j/BSoQ4/anTbu936qSz0aSa33J8OXZU5qSK5d+tr62IFH1Nj/IVdioyjOA
uiJgyGNPZAXDP2SCmRDa36V5SFV06rx+Sy40v7z6WirQJTN8n0WJ0MLYzCAYIdUC
AdxFx5feHthCpgHDqg9rGLViR+MRubImslGuroCLYNenXDFs9oasmDCppTKQpVA8
+aO3hOy22grv5HjxBIH60PcalOjW4TQT/D/tDSw+OV0xNi2Mjq8p40QNd1JO4YPF
fbQjTvfmhXeqrpFi44QzRofQIoUNanYyBfjwH1/lDLfu/yJtvruqPo1qsFfBK32Y
143wt8IDhiIoqpt9Jc8GhVhWpOoAtYUlbnUxloIQ3P9Z3O4wmga3lmWhBWWn/aKM
gIhANTmKUl1sbu4qZTakAMtT3YuClSaKnLB9LPT3qt1IujoyGkRpO95yHwXSHTSj
YInWxo66TKp2XU7IaQ+3dEV57Kqv4b9MNGsAJnPrudEw+MjfmCjCsxDrthRJmFIC
yFuclDBTeI7j6UjRQXZmAsgzKh4wY0ywA6AtrKvWTbeeLauI9wmcYSaxIXOCTb/V
PcS2nQVSc2lk2D3es5jmaoBVCsiyzNyDCDL0BHzLfhaB3XoLhOVtE4OJM56uF1Gt
WOWNFpVidvsDdkXK0kfgsGJgYSaI8Vr6S0l/OlJIs0ZXDLROTbjjj0pjkU4KENx1
NfAHGkG5fmRBff+Y4+VhDJOAZkciUzcHoa+QPUNqPqKeA/wGov5P9YZwdHtEt7dN
IR6oVn5uq8JwIoDM2nbU7IO6yDvd3E9jDxHaO1FVFra1u/ngJ4bMcM+tBqITQui3
bHZEGW2VD/NTB4pt+BQn9In2UtvoVhOBh9IxHeRivOE25ni2D0nER86xpHr0dard
XYlMAB3vViK2EKUwYlX0N3SePiZkY8UtUV+K5SpQj0TAqhrtxdZwy9EGjpEZqbh6
IR/xFV9Gbr6mOHMSOhxWFa/C7g0F+tEUPGBUAlUv42vS2uQnp42l+8a3BZBbth0P
`protect END_PROTECTED
