`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1C+G32USPPQlGJwQH9KecsjIHeqXOA0jKDd1HvL4JQ86lr24rPcObcTtmfPPW3aw
E5EXtlGdarr54yqSzPvF89KEtfUU4RVkyaAbbjYBA511jjmfxHGOsOThD78+haCT
MRAeeTu47tTi8bdJhkSKEKvdhYXw59Tn5CYmj8K+LzhPFIZhaH6hw2+NBN1bN4Bv
PPIYnhOnOLJxI122lxADCSEl2ZaiHBIzcWUHhYLeLedp/8RQiEFsGUxxDn6I6MSA
vtviE1MOnUhDijSeWT/SyaipqG24qUNYw1nenLPzcJ1uVozsOC6Z1O24QOTH9RVK
ylhkGJdMyPkUh2QcKySRwrY+BUA5t8Tnk4k47dFH7g6UJF0QPzP/ei8GcXtymrrK
ZwKuUpdwJX2mOH1NC9WRSaYLETezpEIRMzuq93gMKzpmsOebzAoqXnqVWd3QS8/t
M4gkE5pRjQ5bUY4hj0+EPzDJYzsI3DEV6oGAZVTUacOZ2e/FUmBYSSbqRa+GlXeb
YollYvS/stL7MDq0mVPJRBaAe1fUE+HhXg3fHemA9MEKIvwsy82EuraWEou04AFK
wk6HuGUv4kVtVqOIXlNutXICtGSyHFdwibFsv6ZsrFk5qTUWIgzob2lzzxVfKqJD
BkQkxqO2frVChu0+wjJ+8DS7IwbUA3ejGARItlwANsjJBW5VqbnFNhwsFkqDIA8h
7ct1TBGE0YNKuK6NePzza1jHww1LrPUEBXEtUP+9ebyGIpSJ4JIy5NSlDMuvqPay
pPNFiRaC65WlC4zEf3jscH44o3tsWMMy6HTCTsAdj4OfhGskhY87ZVcfe2uBOuwh
sfTlngSROBb75YkWs3As6u4w7uNEeuif/DX3k0kkB8J77gyGbPgdh++tgiBcaQOQ
nzQzGJbjMHUlSiSOy78NkWzwX0qV1cFxKiGnZSPt7tTHUkzoyu3FqE+1N5qlT2o+
QkTVjlHahkcMysdnsLtowypSYUCMG4ac/bZTtLAJhixmBZAPwl/fKDFX5BImDaNg
xqWMOW3+oUkzRH0QRAK/xsbRMu7y5z2/sL72z+Xvfp4FPKVdTa4EtT24xI6VJqb3
FCnlheoTgdhxsCCcQeLN8EyuBAOBwtxgjxmI7OqudkRxiggc3jdng3rj4MgNH4j4
URrTq4+pRHad9OM67mLSrbkXzyHehcKEEFARHBJQTNGxiKvoCPZPE38dR5h1k/5S
lUt4yR47U8GfmZXek5O00blpWTpyDhrfGDWKUiSNwhMILJnAfLmYcIcAPE6vgTnJ
bQCsiI9p/t2+cs1A4qAQu77RLBiFC/0bu/5pohylpXKieak2NVwKj3s+g6T7EaBo
GP9PcSiNEwBG3liOdECcIuLbu5v4UM8IVTzmV32D6HuyzUZes+SM1LODRZAKxq1i
Dcp+1rJcn6nofqG/xitjXOBBCH/nSjGj9R4WI4FKkqPIL1tZ+l8Dig9T8s2mq7vF
FHf/Y1qQiTA1IsS9zpWPbA==
`protect END_PROTECTED
