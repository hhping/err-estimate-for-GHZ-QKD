`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXytufQenCLyS1XWHm7lkApTgi3bI/FaTGIAqQXGEo/A9szvtLiVuas7GP1mTYrg
jGInhMoefbgRwDpgeU7HCmAc01CwH4ShpIZzTekoINlTAySBZHDmS1zM0hyNlWsp
ekKCn1cVAyclJKb1IMN5eEp8xkywEySqqcQN9SYaFzRP9sNWsZtGNMB7kB+NIXoW
RVkXNKKeGdnXvwhY8bT6pwF3dRyAS+9Q44oBoZDgAsoN8elDWn+VoiTBH4JbmlB1
AQICa/l8NupKNd2L4EnsbjZCMq0PiWijt3ixdHAkqXL88G+Z+OCEKt31ugQ5J1GU
C7Nw5JL+NfiIxvUzRuMN1BtW9rZ4mUJmsd4qOAKMDGrRS25XP19ZenivNYRhBGyS
KlNl0gWYMD4jLclv696uiVh2Qk2LBfcsNNUithfCUwzlvgLymXzcgB7Vi6ALvS0Q
iAzPLAAm6yTTt4Jjh9AgcvXmnu7NE1NGFXRkNzMWeGtouHsvjAr2XnOVpLycpdPg
FNNJ92upEp5SXsCEsdMF1MIYxpGyFAGicyox1OYMIkgPtZNl3faHTVU0sJGBBx3q
rFJeFY/fDuD8wdf91Zbvl9+ruQ35u8Gm5FTcFgicaJsrAPUzS3kDtLdxM20EnW2G
wKPoO2ONcrh67fOlRG6LJvr8HbWoJIqQhyWJCnoO90ciI+pnpNp2FULXs+muUrfG
zd4JyMzRCbX/aAaO1Y6hZ6s1C2SgugIZV9De1+AtWMYHSVVn3PQKQ66Mmgxg9ibC
t7YeL0zoi/xwtAKD87tf55a3URYciKYNGwatMQJQUVDHFj3FD4xnAzPiMw+tuicp
9foDuKH7Gfjdy+lLUzRhVzLbC/hPLShbSiTeYW+Pv9ALhGTWYiCFXbUrGtZ9TL+i
0iXNBEsEvl2AKYiy69VCkTBmq2szu5e0mVT8fNGVABot1kwncw+kWhrXI4VMbS9M
MNdiPU9+6N8ww527rFlm0vOeemienOTl4CMyIzFs7f1QjlQYTLeDuNjoALiIsUE1
TFL5zybutMxr/KOFKCRyP748JNFc0YlHW3Ah+bcyrvWvu7s6DMKdd4dUYYK8i0BA
FT9T7lTVsalBZT4KE8flziS/+bhE2eufo6MCBtVHDXdWcbQveHYz2hjByLCCAAXi
Iuw03dHP2qlRlh3Ii1IKodLho7V1G2qyPDJkWk+IN/Ggl4mT3wtPIGte8Dwhmvq9
xg+1j6oX9g28DVcCUbzGB9oH1UaVwqCFtNccauh6OGcMeog4ZQXvsvFCIBx4jdhP
8Un/PshI/lunAZBzCyxqUFW9IXislrmUM5vfI8hxSQpQm4fqJbb6ZSdBho6FI3Hf
sX2Vvyy6AZVbiWCOXlKAIGX/qQxYXNDrntUkVW1CXTG6kZ86TvavGVSMykn8XWN7
p5hE1oKz4rt6c7raoXDUqf4UCXiBRWJDfYrUgtmxG6IMt3h7m1ysG4UC4Rmlmr+V
CnyQm90ic4Yi0Za/OpgI+vyhcdd+RyPKZD3aM0aaeiaXwJFEQ1L7NBUlZYwD9t67
qVEIK1f+SarVGQqpwb1U0IB+cs/37Mo1jtRUDwi1FwWWiNuCaciov9Z/1FMBTee5
U270k5QekuGS8tjqHB1IVCO5ydEwjxvRJpKBWyQryQFCwe23rRvXF5xZ09YPhaSF
8uG1kamWqQ0HumGez02EEzp4gphG582jmRMyM0jZ7OCs1PnUruxoia0s5TrAaK8m
fW34dM/+lbLqbn5++/cVHCNNjNqfMJ4P0PUl51MdZwaGjBmkYd1CZ9oOKq50o3/X
w2LibGfSz5ps0+K1z5MGKuwOA7dr6DGVzHzygtFQGgD+t5X3cpJJrnLWAhE81NoB
f1+Oar4MqDVZmZ80QFTTCFdC81W6ztYQy4D245QsqQCJnkIY3XU/cLoCJqE3vHYb
SAuu2YC27YRh08Tcfi0gzusxJ8B3p1B4I2cgCj4ZcVnUpWA1YeDJkBQ/dWo9wTrV
UTdC4vlk6aXBMAN4+Eclq2+tjsr+Si2jNOhaXdtaYeraT6snLa9H7anTljwA/VJj
X+u2u4guhEPwFT447F/s/+Ws2Jvjv5valivyR5qBUeC6ZJK63yc82rw8p05wTRjO
LuykeKGLuSVKxd8d4whYg1rpna9qTqhayixakYktZhrhRFy9+4394u9sKUhzrWlf
0hijQtavTdzuNDbqeuDo6mbCQhJFmB1v3EiY5aqqRXX2FLyt+RglPoTd55Q8cIIN
4nqAH+Mo07JC0In1yVF8Pi96eCVz4TlLBFW0dDJ/8KQa/XoIPPsXDSxAu9Owr/2L
AahBw6/EMJQucxrklz2McdZpAYIBFeXLQ7NYzD+lXegsIFINOWvNJVRytuzlyZCg
TBD7mBkRwnQcXqnVftTSOY7TcUhF9ierH1jvGUV9WEWR813GA7SL2vbWrvPKy16D
sJlImLCnBVY/PC2CdPjmSIm/W3gU8ZroIzMQ88BKxAHePO8ldcVVMTrzLIYbHW0u
RHP3d1UgTyyWM3yXdns2cjX9lBAu9zV90ZQPSKFz6bQ=
`protect END_PROTECTED
