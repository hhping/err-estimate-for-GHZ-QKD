`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3SjQUbFZB/G2S/9gCCLhZgrdzYL/WPSd7184QMNeYlT4SAEexu5irrt6xJOroA5
+X9t/q2upRO8h6TPYs2tKf2jk7JyNuYr1L+sUIlQ6E4rJ7kDFZ9WujyEo9Tq2/Qx
AwEuMWr909fVhYN61eijpG0QFmJIk/ZJAng548e4ggEo9dCdxVpZtQ3LdEc8ldac
KnlizX1p2SYjjdeRjLjevvSfLf1kIDrWYdJpfqe3JH6CzQGNNiVUpCaxfBMnChPC
GI+Arje/SMeJ1cfOHg8czEwP4RixTZPj8VPCAEs/QMgRD50wEJgCRlPxjJdMPETl
fwhJaeQvdw0a7R8b1U5sWwlZ5m62HvTyaKoAl1eNFo2bUdIqYFdzVutp0rHsnTc1
Lq1CwTZEFuGoKXj8qTVqbgNMLCmO7mXAm6KKMXH1I6LGW5yNQIPy6vR5glyA/JLc
eXX7lE0w3YhcDQKpa4Tr1hOjjLBGCIbipaqrnFh85+t4quHzPpjTBxMfCmxyc5Hp
qZBnyng1rb0H77982fXFdCk+B4XEgN6RqyTKEmgVKBdY/+fnD8wUpBh5luzyVj/z
R30KNW0Z+CxY8vVBFd0+rgySNYb+ltwM2efaSxVaxzHgxhlIqS12oNAAcrbNkPEA
yGIRKepPMTx/KYjMgJogIIs5ygcWDQWbGbXIV5eKPBhERhcUVswIVhFwNzHqXHLJ
1M9+5gSujOOHEjd4IBh2cnzDL1TfMsMk+j6gMERBgCR6GAl1u7JyV4ZE1z/yp03/
gTxijXIP9uzWaSqVr0ycyBDyfT7mYlQoJSRSG5pVpN9uYcaQELjiBk0rhYVHX5UE
DNP0Soo6gruxdYuviaQ6y19giA7TElfINloc9YdC8BKf7YZWNztuqFJnsbv9/GOf
v+PZ9r+BeDJ11yjGpglYPILPZjFnYDEsUgwZnzd8VFfMAJNuOEOHIL2/+6/RH1/m
KtObbfbXMF4Wtn6h00H5FYk8xLEvERYheBaYfXSbEZHGUxlMhe5173Q2CJ48cPnE
yWXvFiqB++gl+ZSfnqcnZNCzbxfb2Y99W2MLQ1rvAQG06QBu7UeelLIIhBTqcZ+E
uTi23/+ErQX0yTlSVySAaT6S6hhSiiwCdeGF0DHKmsyjVpq9sp0RzDACdmwrH3nS
Ts3ffZiUCw3+AfJrFbaZge5BYja577sto43nTiRYBllyUybfPxTfu2pclIbefu0f
+5H7PZyyridGuu44pA+ktXKcWe+QBYz2tRpEkGRS8R4pjiSh0HoKcyPGX54OM+QY
ygkd3g/dn26xoXZs7Q6469bnrr5Qgu9B3KObp1B1+tg2yrlOOM7FGChn4baTZcOe
yo1eCdDIPdCrlRMXl80eCheGu3RBxeqf7Ah/VR2+xvq7ZUq2b/dqReJrlGfpG3Ql
tfe9Uh93MOaAokw1JN8X/uO9F7l4P0tcXVp2wizW3u4cqzH3XgjHhTsJ3Fp13YDu
32Hn5H6a5RUCeB2kBnaPwwSDy8NI/2J/mTk08qZPJi0y5ajQhd3mQhyvuJmkMCtc
iDfBjhP7lw2i8eFpxLIRx9rbA3uWgiVR/Axf+9BF3Gj04RiFcDKcJMOYiBXUUOU1
IaEEJ5yNm4fbOiDosp7Zhf7jPE+JEphhj0J4CuY+hguBVYAncOhD7oHICkUCc/a6
v7BAsbOtLgQDSIYyk2rWtwXmK1cX7aW3M5ujQDwevBUUGNZEi09AQtsABdhe5pZu
AchELeXpWphEascdPuK41zBS4xvGi5D6ELm+jh8+14bo0ClQkC5OM7qDL9CKW1/J
CVqe1zpHEfIhPbVU7ztUikmtbXKDMdY9EGbnfVVdVKiEME8bpTd/wQj/JJMH9WR3
dwuVzClMY7GLxrY01FTbTpcZymPnTzl8FvRAqCS4uBEBvCAhYZh2AOyk/ydcGn9h
ojMlSRciidUxK4s9dfrsjXDjQhbpt0sqFTrg+HcdVPQvSyKwB1B9Dvu7WibEMue/
WDOxVmK7ekfE58AIFMP71c4AZIAOxh4dk3/B+ZdXBvkUTKlX++OHPFXLA7yQd0TX
xegsNQc+Fo/wAhqNnHw9GufzDxUGV5FEELOcP68TK5Tu1hfW/GoiciaIcejfJZCR
Q6+iD8XxIa4bxd1FcTHLXIBpY9G7pcr+iD63v5+wS+W0WJVqPq3EhLE962a70aeH
4UF9og6VQQv7FzkJ4LSq+RqjEs+Xu/QK0lMInMVehU0JaElO4M5FbUhAB221+3Z5
1cfLhWQV9aM3F8pMjkSJYuj03vY6WOMQDi7UGib0qvlAa4wt4zZp865J5fQCDelB
yZsHJkbHBKnBJqCvfN9E85eREKujy+h8uqTD1f3TILQC6R/2/B5j2VHp1xdgaxl3
JOT8dmxCaiFU0NkfOZunewfx98Gr5SBCjhOuN/I+DxN+LN0EZure/BDgJtwG7XRi
AhIPpqGnAB/aa9Y+4rsk2uJHMM83K4tG/QDXg7mwwpaGbYPd3HbvS2BoXnTz2kSY
lNJaFqqwKwbHW8I2iGRucmSZpuzOKgk77mwXIALwUj0VPmRTcuRYzAJr6eYE1nqQ
dXaB4ghtsbWWq7pLGqYAoGKfeM3QxjeEdx3PQpFVRUPvRlKvJ6dsMpirkZ+yf6TZ
yacgMw6BC8gx/Zjn+mp3R8t8h3BuRxRZ87aOb9mg8MvvP18LKEj6ykzvKx2mPDy6
0FmxVNAaJzXPh7fv/MLR/WkTVkUJ/hqNmx/de5S9UVWMC+v4kETKl11saEQlmbL8
2WJ7JYAhmqK7oXgIZplD6FDNDICyr5rtMIlHhngy9NBf8ORUS4GqVzogtvbVC2GS
K8hqnIXUT0ERzEZ9FkBisyq1BFnt10WMDYgJwWgMemCTgat6yeOQNvn5vSHYZq13
ZoCsFXw228HImxfWVXRJptxQMxEYnWuxia5fyFRnDqmUbUdOsn4iv0xtxDpkgios
dSQQpBoZWJwQloRHyxNGoEBie66i1R1t767v5jKOLbaaXD6kA3ZV92QFDyYTNaxn
iFqAl9Lkqe5pkXsBzkFXZuDHesbkL73z7v+bVsg436hqwclG5V8VsFq1aHZpMIA1
hI49je+uns6IZpjcItwDY1DV/wfW9GtNHKe5YaehvcPf+esMp2Q9IMSsI07JCZ0S
8OSYodPmcQWIJ44mTXlC/MoZaKCJtCqEz3CBTMiovAs21XH0obZ7Qji2eu/a0y78
Nyhg5hZUfdREdUJeGWFevUzd+oGbaU9JdfM2NIFQp2ktde2Q/Ab4af6qbTaWuHrO
wtTo3h0chMjdbs2oXXVdDGsFyxTXr08DudfqN3Zl/Y4zYG++ZdPNJpcCU7EzHtGI
vnOEBS08ZbllOL0R9hz+VKyAMOYtqgPXSxCBRA4wyaRGKD+XMJtm5SCtTM/hU5kt
p9evsuO08YR+8uaD9E1d4g6S2dsuTGGse/3F0LD4mvL0kD7lNWqBw5ZjPECBa2mk
EAztm76ztlJ6zTObUkgbYCIExhU1gnrUnQftvzEPdjx/KxKQ4Qa0xCW2vAYOOazR
2THnxkJUfsWI58uNxJzNvM+HJwQFZNsa7LygPDmPS+IFM7rMo0IcElRJ/NPnWzD4
Qmd2a5vVzRf8B9W9dyn2atY5H8N+ybvnM3BW+gbQoqMO2Y1tY8l7swmAK02L6sI6
5XcWoTGrlXgqWGY5k37f+702fxcw+ElOzzFF3V49uFUMfxkaOanL83+J1VDq0Jff
V1hpNxmr9NxdxKRZSul+t7Pe6xZYsnWppydnqCEw01sxC2cs3CVhYcsK/P3qABL1
oq0hlBPG2TMCsaKXIlRZAfXGOSRsUOkhUAKTJuNDrSWrlujF8HVTJFPi5IV/xt9J
gcqmTIhcp08icpR6npmKmXYQUE3YrWCkbr/IUC4shOPGGIa68gETdFP0yKDYX41h
mVahcdy61cHnk0i8O2xXnoHBnCIby8MJBq1OphKLZpTepIwwJPBwPicTbg2p4dSP
DcW6ydFDTNAERZTNo2yEOigHL7sHbHxdzY3DCnXq6o3rybZJcLOPVNvC+ZwNWDFn
atz7ehxRe/UQYK+8xPRqTe0065AKBmaU/Cn1clrmhr8X0Ow+VJQWgtYSXWwV2Zbq
XaIBQ/X5wh+jcAH5vpjjv6tEzsGxC+tZwIasdsEjGE6MLmh5JSRkzsdqQcuayzpV
xFsee7p87gSxmN0/628YBqgst3VqBLOfOydnQz9jmDC7ho6/dHUtm0uXSJD77rPQ
qy3uFlVzo9rAzlad7KUXGHhpHlnjQl1AaSSyGV/ynfnQCfdywQ/3EBHXWPRIkWzc
aDLYBUu2l4M+GdLP+dfe0iFtLbixq2eZw+6xrHAJ39zShWTHjJY5rX9aQtNJUw+5
niJ4oKpJqzM6Ch8JKFHF322p/uS+GzU2/mQjCkPKPDBMOMGPOY5ZnBaL8PMP/MPb
KABgp9H/Tyz6nwd+vJLm4opDBU07LhalPsK7FkUdodceUZTBUoimHeb7tynWQvCm
gl+o0PAZnZsRwn+BwdmMdc0KLTLTdQow2qiSZ3BTqmY5gmdVBXaagXxDi4659RBy
GK+RAx3Sd5QBSfQD4VlV+BDEMLVbPp/I94m42f6bi5A/fIkn+NsNU1RtdoMQd+9y
JUXzcCudvmPTC4pR3ROAXlH1N/xn/JoUjliTXb5agqvZOa7WSLLfc6e7AcuRkcb3
jyc+NJv6TnZT9GSjd4rSz86guIlAzMr4En20oGZQibxlyRndYVs5BWnkh2V+1e+g
cM6cibepIxr2tW52nw0BogKbmHjWbW6y4dXv8MB6wLcVU5M4KYUmrTtO6gvHQ9BX
EVX4ZIZ4NWsupculwtZjfLITF36PZ0SY3Fxe/YGP69whi6lwtQ5rweOZYmFTg+jf
/+whqpo2gGPIpPojxRAkjtJSf5eDH9vfR2HFjAJ0YxzztpLxpkYQyiuZ9kMiZav9
E5a4tq2YIe0H4dzZnpydom3WJiJo6llRo8rf/cB9o35ummsdTh+ShsTFJqwcFgFo
raztB6vSj5NoRUpr5/8fU9kmbf8F2WVEmfbwk/s8HDPB/KR6xj9OCTPVC/G+xY5p
HEZr8EfCpBbPo2+iaV6tvhUlYke3Bv/fZOstptfriIjME+ClzW24R3YPXgTEdubT
bi5zWZEBDyGhHlVEWKHWyuD5o3oAGIDHDkrHtRy2VwWwBILHX5ATKj1loX1/pqR0
jb0N5VqrdihvNskYBVhd5hGDgbcsZhQbbbhB6p0CEeG9Ad5VBEc5WCVZP4h1GybN
Hb4j5CCQU23h0hW22EFnCgIZ+foqmPzI71Hr1gRmSxZfOCR8IfQKj6jSOo04Bwrv
fY8oyWsuqRZ0BxLtOU+f8gvD27mj+4UOhz21HxOFtR+UVRuibI9rtpyHqy5Pyb1h
fvz4gKYtdDtJQA/LAfv0axpqWBr3YJK2lrkbwM7PLZQfVYigtXl8uT3P9LBe00bX
Wg2WcvRtv+eIMSaI4Dn3nxOoBh+c+VNOKc1eiynF2I0G8c/xZQKsg1JihzDJfeIi
Ta22qCNiqcUDEfG32RIDUm7FGL0n+6WprJX7cDM14COEZFGde2n2yIplxXnGK2WP
unrK645uQvKmwOkrvFb980ojX/z8zrJ5fYJrd96I8dbKgXR5IQH6B64fKIfSTYsc
ScWNb9eAUuwvgJsg13fNW/I51OxvaRk7X+3vUH3Xd8MZbFAhd5zoiwZZnBxsXjvm
i3UEV5mIcjQlK9MxSshBEHYuLoFRe/0QPD3Y4VLJsBXiKWewZikUu7rg8Ah0hUQK
5JhFQZaVaqYRBWXPV1S1ChT2kZRJJbCATbbapkqefTDD8HNPpAKeAiB2N+as6HcT
LsY+lMxLf+n7usNausTBqdc/rucaIaM3DBfoAGP5lv5zf3GfonQgXMcHsZ3FsS8H
uHNfh0lX6Zj+61dp9LHVhg2kqhzffmXQkG3Jv/mwrusEy7s35y5t6/zPHPKjqeWs
heD5V9madl6SupvrmOdWD34CsdxR+ELzaOx2pN9y+C3c0jQDCWwZv2HJ4MhavDXh
DFdbLMrbYedMJB67IH0+iTho1W2rwCxFUTcQYub0IQbUtEyAFwkDYy68FQ99j9Q3
5qA2lhb/MlyCm7cJk/x5wMAipEEDth9mDtDt5am9tF+KMdKhFjNEQqzTTitddqbg
FVYJNTA5dWcRuYQqTTtkG00SQygj3x512BEAxpxu4SXah8imp3tLxc6+gkplJiSg
Oh1Ab9vGKsFEMinzBPCRS6tMQnzwskdKmEbLnr9Y8qdAbaxyy0tBZDGNq5l9cqrp
Wcx3y6RdTyZOntFH3Ec8ldx+Ub64BfjNlaM91rJQgoQ+HLFB+hDryWLABqImY0nF
oSZzKZS08PvHDvE8Rppc3zuTCk/QkD+f2ijwx6WcfgbTY+L4bPrZ9oTnGjSYpZsP
JrZXRL1eKyPz6hIw3TjkmFV9fDwC2NIaHqZ3R01yz1rrWQIH+OlUNwGvfsxAZk4g
1Sjxufi5S4/A9HuVBay5kQiwalxGAm160CTIVtAVGofK7aj3F/S3DQsgbcLlsEPZ
P31sTD5y4WJHaQjheEc7khgJmIRRQRjdYphyjhkPezjsB1LGJthpO+cjtrSImNbg
gyyrdYrlncdUwgNi0RPyd4NSoKmJAwvNcOzrkU7rNVkDJccVPBufD63KPF5E6UpY
dVR8EAP3i8MJHhn1xIBo0TNZCACrVb0Cug3ftE1f4hfO9H+rdWVpG/8gKg9o8WQB
1lIGmBCUoIKE0FpP69PW/Dg//krL0XUBRUN59dizae8n8f49C+d9OMWqepuUlNX1
nLGNwjVA9DGujJTsxuoXO9nl/LhS9ky7JwMZ1l39l9p/Ni7EmVyguyNPGsbAaf/I
Z08wsuvXpuygz/EtVT/v4VK7UbraLTjmKn1terqJ/yKhsmDdaRrGLGe219bWlAEr
vxodWuA3aqdqb+JvNDyP4nzqrt/Je6C1Zbp5PwcsRNqaHOujUDw9TXGrb/T666GF
hQs4ygds+bw1XFVrYzSL4r525Y64Dyvq/OxvuAFdepdpRgY41hBaD1r3N19DOiIB
sOujxfzNyndb5ma0c+APvEiTOv7s+eUX+oFHs844iIN6Ovc7kCcmyhh4RHHaUuph
4QH5rUt4Oj1bkBVemSUXcuTB1E/9HV6flmiXHKXI4qtSR/B7DTP3FRTQ6IQ0+Z9l
aHJU1l+UXwUEIkJw8su0INtCOJRgEMXAE+wZAlST3itrimckOQke8zz2VogqX0vh
FjNcBQLTbkk7hWdSSP2e9uBXKAAcdQZTVlA756a8fGz/9JylScQQrHxOVy3QpXdb
FLRIyz+xWoGDMvFCid/SHsi/HSgzjxRebCTSpiNynhKGUaQsSniYrA6bi6Sws9hI
LXYx09V24kcbF1GDoMTuRbUPphU4wfVdr0NybUANHJPG+mBkBCsWVQseo+PAYD9u
mOaGiq/CjURR/rRkY0KBSv7JL6HzpukGEZZCElMgJDghZKS+Lk3b/aetPxzAhvyL
RlNwZeiO1HV4DOTROdyBe4YceQS0Enp+mobElC+Xmv1KmKwVJAybm3vVQjTSCuQ4
59AmMzJQOwUjOOKQ0uVhfaaH4y5GRq0CjtfKloKQTUyUs8CSV0q7pTxTPAwV0xHm
BKpZBriinMT4aFAA1X/GmhuFz06pjYDaG/xlh1D5xoWlpOwnRWW85N3vtbQjubYC
O6S/WTpVQhwy0SQsU0M+TblPeeqGZtPSEeHjNUVxJsodYW1CLAU072l/i98/kzie
1r4xCZpSlO6Q5iaPLa0QsORufeCMYpC1N172b4RCfILMxL7hl1HKrlC4DcpVBp7e
gPeFki3IyNS9J3Rab+8eqKUeqZ6vyay3M2fHK96euYjcW+84BUkEO09eBCoxIJPk
4KxC00gyvggSB2DHlSAp7dQmUYXwMgYLv2punzqpr1elDtYP3fvpZkzd7wx6Z4ZL
h9LiJswZGKbUcOL6IAwub3ZoqzJ4V31qbEnvjV3gpD8NrtTD1ciLtEyrmcWvLLcs
bwBRpLpvHVjVF1jTMz/KnSCGQLNvpVg7UTpUgZdjAcLd4ue8AzjVmv2HfkWndpH8
OTk3y1kDw6eIvoxHhMny0Gi3XRnUfEPY+4FWmMA+/vzX+JmRlS8EOJCsR1zvJ1t4
qdLzWf6iXAKqWTDhALnSi+jCoyhCAtoPq00waNnXMieszg1oY7kWhk7xz1GvnLUY
OR0ThvBneWjEcNA3oO/pOLCle2TrFbGkheVNkITblrCdNbfx4Mxzu/SwfL0hpNPP
pYBEk6jp7lIZvA7eO+wPcZ6AIPMNe1Q2p3PPQ3OyFgEeQ/BnV9ounYzfAfvhcFdK
TqX2HHpbyVuUtQVfXpnu1KISXdJmu9ZxVnqxX3NgEUO6M7bL0c0gI4twZDl/Moh4
7G0MAXJHmmnTrLycLksBQ4XGnxtfN7Tr0KsrL00/J61lWOmUjQmz9GeoRiLGkC/a
r7sSx/Wmk4B1M9LQZoyBqOa2XRPSMo7MHyibIrEPXRYOFvgfKe4psKq3q8l991Vx
ekYsMWzXTVgMJ0BIqa/pbv0hUEPfhesyhmExXWo+tBDbS4VOtOU8LWbxgk/PC0dq
zIkBPXqzANI+bJ20UJ90WA034GlMkL2yDUVDeCtvR4lWVh81VXrG5Hlay5e8kAQi
e402yK6rdI6GrF9EIHPU1OFa6pSyfL7N86k6uu1V+AW5B+x4rxckoQiRjADQWfw5
qcsELLqVlerLUcdxUze9AW4FauqvIpDRyy+MozaA2P2MVQp/bhkceNCuCHJzw/l2
P3oemHlYChM5CVNp30AQQLdstsrKAjDARepJtDSoIHZddg/r5zBiliubw5IPFpQT
NyEj3/wlmPL2vhOJeneI/JKkaPATHTdpLqTa6Q4YXTVO/qLa1A5I8AMxTvBxxb1s
VkjziHyR6I5dcH61RVNS2KaplEToKjqaLiGlj0ZG/7V9VKgOE9B0Wtnm1VkUsWcv
6li95z9XHkLrxJ57dQMgN6+LTTDLjsXla3UOLKNxsfftz4b2qRy4VuQ0s754YyXi
oEqJhVhV+hqjWcR2muapn37YoleOFrTwwpEmIvxWItwV8/H2YCIXFOFfeGTgg/Q8
ZyCXOB6ZIIXervvnqiWgcdSvmKdHNky0JoMazh2sH2MmJKapikIC+ti66yKxrjsm
CST0sM802VYP9C5rNCTD2ZBZhNneSp+aBmoO/MuiLE7uUM8J4b0aWcRwc1+bKxoC
xZaTtfqxuRwy/nwYQkyNnBCZOq80mhk8pDYjAIchDa5chCjC5bm/8Tdo77virOgv
xYALd2K6D//ZTkw2+XYe06jNt+ENCPFZh6FnQoEYhYhOxpNl9yL2vt0Z/a25rll3
y8Zcx7kyBBQPOQB8ZZsMWN1+Nwj91JdiiWkLs/aDLRirvWATe5IBR0kD+mn65Fc9
VuUj6ijKrHUKU/IHcBMykd6cEjdkAGTzLfS3GDOmk+nhZgCO6ul2F8UkoSLLj0NS
AoXkkXik+txmj4qmnEpL2cs4+DPRsU34iDCLq6rhbLhGjieu4grRxhMuG6WvY3nV
xCumpoPMRwQhPgTagHrvAnL2kKTWW4GJjAp0iQknTUPf8E6kXOO+gw78+bc4++hm
MI39Xeyl/nEQfIbRNi+8A1p2qrpTbMPmf5LDOyqRTslIu+cDu79nJghX32fUgK6E
8bbHkMwmP7nIMPCKuXmB0EuvgFI5DPZCexk6SX2u4vTSRI1hCr+Bs9AQb5wxzYWF
utCvxaf20es+bopNLZYhbM2xQUbCMRE3phC1GbKiRIvXy2EUQD0rPdlpm1e11oOh
pe1ONm3BKIW12xht2EehWySumXDqJjKyWWkvf74zgQU56cOfnNuBi3JyDb3vDUdT
Ql8eZMnNF04DF/UYNqyGm2Nx++sz9AE/znOw6bXXR6Zocr0+g6GfAjo4WlQguIyx
d/HG4jXiob0yRKG/iAxQIJzsvlABD0HEOF3FBqzOwD/4AzsGI1H7f50lzXou7RHK
iOLnfczA4IVvmLG/krkKSyVIIg7UxiNV84I2UI7eMxTg7wvriwqwV4oIFjJaVizG
yDIVCCa06+JAv+1qCr9ipQro5FvNRLWoMTOFWgA2pcWLoLMz74e5Qtsf7gB3I/WJ
g1nkTP7xRGKKG3A39X+k96yx9i7pqR4avn1lfzzew4IpFBbUa2oqpjY2Lw7On15e
9JoSR5tw3dj4gktg5bSnpgCbvdGSgpEsw7S6KbFR9+5RLrfiRGundLIYUtYcs5p3
M4HF1NavWjqyJ+6AtIHxthfUSp70tdHmxaF2tK7yyECr0FDGdoKcenEkmjQFEbiU
Z7bvdUl+nGhrTubOhONOEfj3yu2abU9QMGO+IRId+j8CHkktH7DE0gH7mzvslx8x
s646NHlTmA/kXhnPZr0muKMHaDcqCZTNObjfmxj5CE7e5RzCh+Sqsk1vZN2BbobE
L+FW/0t1RJXHZHJmz7Egna6381S0RYs2dYxDx2MiKL7yXuPdhg+fZN26YYHnZ08M
`protect END_PROTECTED
