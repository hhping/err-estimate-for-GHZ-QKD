`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXPbNvm2GeypQIzszrHYT+kf2ML4/OxakCBkQNViDXMbgzaJrv265upj1Hs2M8j6
eIE3Ap3mPE95/+qTY5zjFWLFhvywt8ICAxa2fHmwS8N2V6I4mEIxi0Nutmirb7+b
uQ0Fx7h3WiDntOne9ioAlNXt3qxTVJ7ThUoNGUGzzzMHUuGCQQ/lue93JgqovPc3
QFly5rw0U5vp20/taiIsUiXpA2zDSCgFaXtIkD+1wPPwoeBomz/7Pw1QeNM4l5oT
CAUCNXNfbY2HNi+mNZircWj6hR9mpnBoy4Ff6OpPVnfn+raim160+anXWhx2FClB
/INd/0GAB4V9VNux/ae3hnizJCmDiCwz0Z2DY/nDjvZR+LqMmTUOLDq157FnIXWZ
yi1WiERfqshKqZRsOFh+o6j9OMYnYu1wvcgMuway7+r0JHbfP9JG0ZHgPmkE3QGU
aemEKO/5yfXV6AYbZWsVKiJSOjU3V/Xo3XmcmuaM/AxAmerfGCapF+Qziay49sZm
7oHXglFuLZLln7hh5YDkYOIytRCeUBq/KFDXwKsfzaXi12hBKe3IXSlQaIVitMha
djZBZupUjs2ubDGdq/ILnfc+XgAZqdZ3LpYu+GOXqLFQ/mhFDdaPhgYyMOjBJ9pt
7c/a1FOlNM8WdunxD3WcMpLOcJIvP5cfpKoEF1AcR1jiNIafBtPTeyINm/zBSsEo
/WFEKdfLhSxEC3W7+aetwwa7E6gXBHBVJ30q1hgfdZ5in7661rmrebNhdKzuYln3
VibCgErN86qa4t2QEK/53ZVVNRwIrLLaznHJTYKHY+zLaAf7uUNx80DLDFug+6d4
2BGuGhzb+Gc35jus6x34bIncLR3WP58RHLx4d3taMiPIaN6CrUudd/BAX6UU229y
cxVDjbCUsqMTUyTJ3AAHce3FuNPklJjYUuVjm9cGd7szUMw5LI/BAcO5/aI/wEXv
tNpeUaz6xJSiYy9vv5qkYDEC9IkjW/kUaxCrZhCaBBw473gXaG6sS0g3+FW6vwwt
towjABE0E+A0Fz9KuvJfqaGujQUn1MSq14oFvtv/5Fn+nvaNrzY5aIaxn+c1LfL6
hkti2YsBfxxvp2kvLTyZ2dqltM+CtQwoThjX3UD+ZeAa0wf6zX98pOL0wRL9l12N
Ik+6Qxh8i/fBXrO5NlH19RHzl0E2OYpBmv6h3cDCC6cYKz5N+VFa3X+S0dPIeDKz
m9Yuc2ECFDl6Arfpl7bK9y2nzEHPvfAUjHZGb6jU9GfVRaDxdl4Tq4MCHJ6luv4C
ShRKGz7c6wsrI9PLrzJVTlk1CWwZc5CbDq4Wmgcaq7KWGWGmjWqbySRaMt9jfiuf
cu9WKQZ3c06ChiZ9tW4euae7o0eVv21Q/Rmq/IwaGTmfg/We0xNCHJAp1H5bhoyF
foCF7+ZV0o915EY7TgseLlIHmMJkSqEpLbxg2gnCbZcYgtXqlTVIxfxURyICHmcu
lhvlQe5eucfzoBZZAz5ZajMaL6iryQuDKxEIs73tyhrlDWVdQnPyvsfF9AAcj452
XIJNhsGtW52Wlv2KjYW7/EEGIFK/xYAQg1z+Fw0v0loIbFOtmX4SPrPeRkzsFi5v
at/0mJefqu9KKf168dlU4E5gqFyGmTeZVfVpD/kwtz5POeLxUZyNCYku2xh0+ScD
hQWHLvVTbb6FMaT/+fAK1s5ak++jL4Ilh+ZP4xV8UcWPLJJHi4yPVaktcdpZZQ6q
4YSawKKOhn/zkEZ8yJTk5Ic5u/jBvzoAU4lHm5w2m89R2ljdPngJ3iMvyjjz0aZh
oU3Jit3QUwYI/rSFVofb1CoMuG1qJMrFnvtdcWTSqbaJOEeZC5pDpKkoYyBrtLBu
Ai4WOZfHF/JFq700iy2Tua15SkTzCsL/aS2Fit6nLGOJ/loQq/mfl39xORPxyTSb
s2aE8vaIWxOvLkj+P1+/kA==
`protect END_PROTECTED
