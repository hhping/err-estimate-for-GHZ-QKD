`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQm9nwT/naC9Q6cZ3Mh5FzxqbNIlK6goa92vjOB/5xD1f7doGYqD0HYrUc3xoJWc
/pN//8nwS2739/NW/AQeifvB0qEABvRgN3Jp+cRzGbsavoCoyLd0qdT9u4T+k2Zv
37iU81F2Bk8f9Pn0r5kQPVvrJOw93+leZ95Sv+xBT3UZXkHXBB5tNpmt/l0N0UTr
j16Ak+AnCLUERe5Q3QYMEH588fOxGjCfkFuXdzo3gbIlVMQWxK+kSn0cLjVsKfqS
xUM/9WX3DE4KSIUDLVFdBeZhxDAVBRD6HDgCNtL2qy8dFMNJx6C4q3D4aoI5ZEAB
ZLNvHymxaVYAC3s8ZsyRcwgaDpSF07jMoSfXDR5V8/Ca+R7R7FrUXbEwK/s+U0Mr
NmRy0L6XUWaKXSXpLNBUs3b/X7M4EskSvhPEXgo9PjsPz2gGno27Vef4pSUhCUjY
3nw2HXwGdhb29e6C0KInlBXedRCZrmSdna8+MCln6RJVFv25XJm6I43ZeP4kjK0z
Ws8hEVGmhU1uuoeeyiC1Zx/F3/vC7XmBUwUCLIQRoQQ4Z8S2Or9MeZiVaNIbYvmJ
l2jgv0FUXgY0KrCypscVxDVmOWQEvVLEKU1DfSBihdlLDJx2pXxWaz2u72W3SwR9
HVvc2xmU5zLlX1fTA+cuxwbbvh3v+qVydfRouIsdTWSH63CYklZe8SkxVeX9bYji
mM4EZvMuHL8ktg7Xq1zJBMCRxXg/mZclbjkFc/uf+9w5pc0WEFN9kGH5gu8PaJjW
2A6Xqo22pru9bfexTCq9SsZE6N1+rUeio5TzRQKUNibCsqS2/pylzP7cTi5e4Oim
YXmrdxziB8L9fo4Rj1ytJR7FlGi3j8J0O06Qc2j6oR9QPzXGlMoKeMQF+agTzmIw
NmWPYRr03wIxPdM19e5XCxRR2HtXPVRS/Nq2bN4lueT3s8rjQpZwNKR1IL0v3gOr
ckANWZtyMz2EV3ajb+zBZJ2mmOkM12rkiTTmDn0y2g48kx+SUA8XGTuEbCnpIYiK
0AJ7qVx+dLhE7pZBFoxkTtfw+gD4eNkPUfgYAbvMH8GZ50oh5WJ1Hu1tDhojngJU
61cWq0JDSWffol3Qk0RH7IYr1NV5xOvR8MEkLe+EJ8kGYqry1aa4mCSJu2jWx2O8
9IyQ0crYbLJ98RuRyRKGdqDBSO0sAUQjJ2TIINbyo+olQmdHj8cvV0m+QZJImK8y
xat0fyJ9ZgD+6LHE3dDFtMODrqOPo8HHrGXTSBghv03Y11Te5qALJzkGMLtdghdm
qEkxj5wYgz1A4Cc9NEz0jxCT61suXqKdofuF4YGnzc65ePyYKMRgHFGrx8yFU0Yj
1m4SepKg0xlKylHOk+AQlD0YkpTas0gIXaJaP68pHpEKhdNeRHA37YgvM120hXow
IGIcoRdNzm0WdttMSIjJc3lZ11xgYiGtvtxeZmn8lpdzGCDwZ7rGXcFDHr9Wj1kK
KHquWnk+3qrN7v1+5almVCkQONQevlFGPbc3HruriwRVrBir2++NlYTZmLk1ooCJ
vOBjVeTwkTwquvKLtWd1RPLPQx1mTwqM+UAla+n7tfNudWZN/JRqXKQWOpXK3i75
mKi7ugoHazZnGrCaGWSi6ergKX/mJE5gLPojzZ9+Usa9QVjtjOBrhvbJjsm0uQjZ
z8OfOTdG7ygdbpusQQjXCWUXLIOZE07SvtrbR0qhdeGdeQFuBl84ptmPzZA38qTw
2hxZ64cHdU5MzU2+DkentBW0YW0pjGvAOeVrPJtZl/IE80s7IRu1Aaf1dgq+i3As
iI01oxWZmpNvBYzhU9/8QZ/goRYpmCdrBM06x8C5OAZhLqPg1PQ4iXemqn4VK/fu
pFNTHXY+GLICrE91VBXJwvDtf5jKoDhxDmMfP4s1INtJ0/ekPkJAq///DimhyNrj
A1v+fU/n/AEr5ejIPPEPo4JsPpimMuu6a3P1wBVIaOkPBOLAtEyY4AUH28Y5BYn3
grcIZZ+A53ITaAFjke5Y/mb7TE6dP7FTO4eDHznpFFLKcNXWAgD3g3Inde7FcuEN
ygg0qTVEcdS/Z9zTJ1ruGLMyZf6lI/UiMKMqFfQS3oft59iruJL7cq2BF2Ecey5M
VKb1ySAGV5zHeCmz3SEq0SFWYIk4h8uI/S1tBcxebkzaPp80eXJ5QNMZKYXm5GLg
AAvsPpKAtvg9X52EK1x06w==
`protect END_PROTECTED
