`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxyxERcfpfJv5Vo9rrmtTeKDQ7Z6bpHsBUjo9FsdKiFjrcUqAP4rBFTE+Oq3QHje
qhakE9QYQfAxCWyDK5qPn0PEWitY/51GvhDP1o+vPChCXeFiFtPQ1Ye/P4at4xf5
n4Bl3HcdGFaT/kxKBT9v5W3biKTDu1a6dikSdhgieXbPWK0TGIqtNa5/UfSILV4S
bQVq1z3qvWxz23evGXgLjcBYgUSIAueAIfUoPC/UfBDIsdbl+H3JhQKJr3cS5dC6
vCs/d2Nb+EbvQkMuhsIXjFOimQJUREg/ttpnsjl32lxBYNt5fDAgAuZgkZdJ3tm+
tj0u1MVrhV5klkCtykHPt1P7gOTWw3CbnitzWSLMa5bSuXvg0MeA07Mgc1RxzuFl
Onez8xJ/jRpEFPMGNPU+Vz5Xet2i8GffIZURN2xBoEjUwZcb6FSJut68K0pcolrH
Ic3w1RNj8UXltTHkqU8lcftvGnlKUeaF+mIBLDzsT9A6DPK9loxw+739izSssJWU
+41jazJofskSLKpaoSiWnSCmDHaahVchJB4Kw/7mVM0EWBl/yWU57KlieUhfdpG0
d52tcIuV9mduECYOivRTLpUKQaRYTMzKj2FJY5jz5f4ECi+NTQPL7AqUiJArtO/j
B6QESC7H6yAn8h0rzg2/zN5WfouhbIn8+sVcI/AiSW7a467W1qU34/h/5mPJfZLm
86OFSkh0GVeOC29EdvZfXhnLHoRs8JZJXZlti4SKMRkQsugJMTPGUvj3gb/7nDXf
3UDZaw2cee2NLf3lO4XyoBYDkCrnUAdgjTFsO/j/CCflKZFqUzv8X2XVs4FN2qAh
3aqVbWZHRr4VZE+vXuC9yp3F9jU6Tgwd1hcjI+S8hIeFvHuoHPo/OtAXxgRAZ7pq
vJB9Cm23IIJvWLNNnVP2hJGTtM1XyEbQkCe5zZBTosGqak//ECJxE6rXxy/A9oBB
tU/40SpIjhICp49Hlxz71fJ/lLb0mqd1sBldXqTyCRJDf5ygnoSMsBOE+jc1wJq0
8ebMA1R6PcJwKAPEzY+MTUEa4rE8Eh+vhKgU5z8FbZVifL+yfBFoZcjwX1GH/S1Z
n5ld8tz65euryq0IOoi7JJK34DZakgEl3jZhObsWhaACllKHudKvu15uWviUh0Q3
4Xx9eUotikeS6zKyrKCJbqR23lwYe7opoiV9zpyz4YQzZbcmalqI0NEmKPaRmHgp
vlzmvFZaDe+2zAfMvikOJTc2kfMpaGbFbm3nZR8Gm/lQEJU0xii2qRUQb337Fi7J
NYv5HiNTlsBSmZ+L1g7V7WiVQ/p0g4+nspzdE1kiw1o=
`protect END_PROTECTED
