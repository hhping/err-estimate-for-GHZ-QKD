`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9vovm7ZzToY/xHzUCepnXNqjgdp68ZBlteaeh8ZZQbHf5/T3yxtgRkGW1YjOjRl
wW7/fiWnXaiOLrxFrlFayEsoz0AFggxGKmNochMNe9MwQNi3Tc5wVPip0iTTHuyY
1eKupo0IuhAWLN1eZwuqZPIcH6YH75coA1hRjrABVLWgtSpvr9jxwxHUJJDh2bTF
6JDmKda8mQxBHTaxxl3IevTjC2VvT+hY7bSlTjRVEKVtW7C/1RshiTYRnqNIzMFp
MNrAz9eiKi5/mlJZEN8zYWff0Q2YvBYHArgLjT2SyT8V1YHs9vRm0G8dw/yyskJc
9PWykPUwtrLh8uyRjnLaWlrOm3mdHNjStlWburiIudgbacIPDvH86iCXGuvfBVRp
WofUUZTk9rHlHjR8MHQsIlz2gbarhxLmKmbT5Uzdt9QTpQj1aEyhk7Q2k2gO7OxI
4UxEZcqTV3MUOOe4qEpMASfliP2PUPRLJF8QAGRDjrUbS118FY5YuYHLexLi0W+J
y5tqPN6HKO6OMFkXpKCkAYKdASrFQqhHE09/k6IQg7kPzx/FiSkdw9XUz+2Sxx2j
CxezhZB/zras9wEDttsNAPsa5SUn3fGpmTpmp39wgsMWGY+aZn9vsXJoOvFzVT1Q
JI1frbpsolPNwBizGz16fGRrFJaDsVpgAv8h8S4IiI2xoVeyevWGCC7mf1sg0hZD
bM3mLdAAGMQ7aIz1FEZezQ==
`protect END_PROTECTED
