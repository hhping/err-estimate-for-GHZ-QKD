`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URRa0RcbhtLFnxz5lW90fOrqZaM1yMkIbY6cb1s1ikFuQrjDzsHPATU8R2IahFeL
e3dsviVS8eM85Ku7NVUAKqOhUd70SS3sYClezqm42wz3GXeoB0EnbkaA9e/ebLI3
8J+P1RZAPyM4FVdXDQjDxpUhFvh3D3b3wZIOsY6np5JpZMzSAHaAikU6Le9bJH/a
HbyzX+T00AopNMI9Mzfwepe6pu0NFkGJ9oyFLbvntbvBdI9+dZpEEtlQ1hic1bNS
tHIpKslz6JpLRxxd65+7zLXGsv8lo8uVsn4sF5C+BYw9xwDJ9mfQzOjYAIRQxuoe
g2qfYR7i3zlYxJUaHIUESeCoXXQvWQu8l6YdiwdeF0nJemIh6Gelgqv8cmubAtzS
CjsHx3AeCl/MeBR5hkOTFoOmcmaV4iOXM66L5yVYlo98kNFSpsTegA2y0Ipb/rKn
J9ZsmPkNO6+vhLjXE7d8Pkl7CMV2ASYKG9UPeeOJhGn1oFXoSsMThfm8V0KAspCG
wGS9B3W1uIzC7yN8RtFBNYbo6gIHbgdWn8PbEB5hS5KgSg+mW5HCCWsd6AjGlZKz
ECqQadt7bHJygkNYzkXKbaYBtK6/nshWO0cJ8hHHFo4JSdHBtwG+Eq1QpJ+HeWPe
ClODN2v/bJX2muPB9fQ0SCxELdpU6BE0K8YBtnVObzNwsonlusfVTyhZogmvCaa2
LMSH+/7kobBWLAsfe8fXlcxL8ZmsiRYSXARI5ZTDMXhzOeSIlbviAncGCn+/Fe1c
b7VPPfjuylksiLOVJt0nhx9d6KECTKzVsuEMmg1EQSYEm24ZQ+gukogoEktlSeAg
NVZtioXzycKHnfP3aK4ubiCFkBDWihNPKDR8qGvnR3XxuUlOa5osJdcgCW5vTRW1
x4q0/6yuBHgiNBm7VwyyP1I1p0veIxOi26pGneJus4aJVxiob0NZNCTMT+9vAHEV
Di4BbC69pFKR9rdJareDyDAzix329ckn1pG4m5Gu7mecc1e44SDmHL3TdfXaeIET
wwcdFpjPfLuvWLOGriT1HxMvN67l4+W36RKelf9fXkQlZQgjWV+8f9qADI700lkZ
EcbCL/jwhY/GH6FyFP/zfGE3La9kKRGcFs/2qjvEoGpdontY+8D8Loaaq8VCXpKw
Ffqr6e7DwSKye0l5E1EVicp3aMxXFBOsRnjoWDeWqx5YuSsuC/EUeC0dU/dOOV0+
uL4EwGLsHyqEfrAw13qBNnHVZ6a47NBQoaaiAPjnqoS0XTReaeFz/nTuMrx6LAbj
DXla5cCgFDxSU9CDXddm2uib6BSJ7fqps+mHYmVnW/OSM6TodcVzMYSWIA4uM+Xe
QpqsY+/v9sejusvrB2TUHodv9dKm0rCJN90BtvJb6jk6eAViDRehtcXnOOpCgpw8
7cFibwhKCTLOSGe7OavtiJh6decs3ktyMpUBhJhyUo0FwhDWMGoy8tMt/SPJ0zn5
DSW2MLwRLekeDGYRY0vD2kvsGf1ACncsE+DLCfZ3ZdwldT63ToFGiQu+Pg/WrToj
2fiftNIxXZ7pWz2gxmfyJ1sN3VJGwFr48fSp7dnfMmpnKqKzKCn6UztHKZUvdQZp
ALSV5QX6k/9eEITJvwTA2cbs0gwVqqBunwwr3NLVCrSgmRXE0jrX2huNBzViSaza
tzRfvX8J5tV0nXXsBLN4K6iOJ076DiZQgoV8gakO9DsF4oxjKvkpjlcWxYIdT+4W
Fc/rtLZvcQl62gLkJfu3a1uZ+cPOLsE1oKF2n92dCzDSHhURCpRnE0UPRRT2f46z
ILrSKRQiT647tAZS4u7sa7MGWoMIvABLqSDzpFYKo0EzuDnsLoX/+97kPQnWqDD0
bu5mOaZ7AmPcqg9gtTw39nEK0ej8i+6puWAk3bl80U1VroXiN6MxmGwTa1zS6noI
PaWdB9/kaHv5mGU+3t9VsHyMzSVLrB/6ZaiQKAVHzJFxvhr6LRsXo5wS5onC/VhL
JqJD2FQH/zUAKSKFlfLkzWWxxo7WfSki61onIqvTjtpF5o+GB52Jn0zdC3aUdqt+
AA17wxDAgrF/McTD7u67xsi4la5M2vPCs4a5gK6LWQQd4R8+0uVPRmMuTlZ1K8rM
XFWIDxgsm87iMDS1D0CFQRBtxjJVelxxZp8H0vluvPPhOq71uaWE9OPM9Fr0AJHA
AkGCdudl7yMwYzLkl0de+Vrz1OB1DT9fLt4Pq7+UbkwrUfKukzZOvJ2V/onVmZFV
yWSG4k7notvFf4X55qAetZDozhqSxMGngcTkC0h7tE21Fy+zT16zMjPjG2RNHOu6
Ge74pzQHA6jh+uJknj76OaJplb3ml5X47iWdL+vMToOhHLwdan8Mc5kYp0HzG6XX
vkdXCTiIj2slJm7WM5o9f5jbyme9W4FHbfDe674XrdyMhVwXejHZeHl+MxcrxEnh
pQ8S4vqvp7DJV5uzIeJ/3GEJmCncUsjRk3hXrvW3QnJHtyxH+iB6UIE0pWo8ZVux
nWEyNNB46rt1MjmD98Bup23etSTrswV/9cdPHnEb1PaIFsSdqFaWajXzGBoFy/l6
Ra+6pGc2qNzApq5upLkYWM09Zs0uCuS4Uq4L2x907L5N8DviBIQjI/toKWqyKyrE
MOP26VWILPNoKC8iOrntoJFgHg+B39N3ggBETow96kkCoEZAQRF2vTMq7EyOWT0d
I5frX1cD7YnF+7hZm6Nu4gV39cGDwgYVooPWR6qkNWc1S/R3d9er4iz2P/Cbfg66
VDCRXSFN2l/L+LlcuzluOkFSFvpx5EMKD4VpuWxBBvx2VJ6OLp++JEEbD756ZAWm
B3CiraUnJYl5oDfDWyov4KpAGv6HpgWP7HG2xyjJc2UsVGgRqsirknjnd7lws79W
dIrpoRQehuIf4R7QapF2FoOUW0acZ10BMIKuu5Enjc1D6RBGMtaHmigvKwbNqX8l
xxg5NZdkPyxMxWrUu/kvnriHIiYPk8kvP56MR+tm7nQi2+wlkjLaKIbAywtKHqb1
Ax047JUq2MRRTGSqKXp7S43Gblz8qePQX0YSjaaOvtuTgPYtnQhKFyhsCPO5Orjd
/ji9qpgwSBkHuoOi2CkVOJxrRUsGZwMYkxTb/NVdVf29+RdqLccTGUlNM1XIs04d
YzgUZ2HJcPwsZNOD8/uuFVpoplExC+Lm5ZXrZbpvnxEfzf+L/8ct13g+Q0ajaOKU
7E1zbbZwXR/A/D2HyAwBSzV3ZznvKW26moki8grb2pVa1NG6fN5LrEjUHOuL0w3B
SffoSMGGz+AJFObfQWFTfK0xr5CRUnEg/VaROS2PS0lebDPayPfpxBNSJ8Wa3DJa
YOwDos0/FP2yIA1PhpZYsYmfnUW0WTuAd5vr2+ipg8rip7uD44zjtCxVQ4YXO6aT
oWMCa9RZJVPlgMIY+Gagyz9NrPg47icxsGdaLJOlvDpaaKqw1DacP+WwJGDru2cC
4Z2/QjUcn1c4QBv1OW+HAqe8PpajHesmCX11umi7RLhO8WTpOQLHTzom2UpW2piZ
vwW7BuM5h6l82VVK/9899bKaD5fmZBe8Voud27gvzds=
`protect END_PROTECTED
