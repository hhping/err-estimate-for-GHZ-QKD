`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zdag00oIU31POkZY5ZCp9R70FgDRQrYFtOeFx/jRd3yWpvtogBMGs3sDwFRIdkal
+oKHEUjbFeYoJSFJnYyuXmORXT2bBZxDQARQ4ZKnHBzCQ7JU5wTXNja0wM7XEhJb
r2mG0yn1rJNsqyVEXqwFY+M8eT2ssYNXBWBO/buf4cI15pOqWD46Qq4hOOsdscu1
GxMTWouIfyzpfqH1v/cZ15wGXzflTUp2lOSiPmAEGM09vvBEaUtBqQ7QuzqbOTTF
sx1Ehj58+CYDUz1+pfHmuhYPVof3SXGnNHcQ4owBYk0nrGmk+4p9lnFrRI7w5Ejb
oetmQihlhMtqEs5O2RU+CgkvTKwswyCG4XW8JGkIrUgFFq2HyLuwIJettDrtkrRu
4hUElDrxWVNoHh05gJPkwcXV9+Ti4lSOjGzL316NAdp2jszIaTuBiApGRX6kUn+w
cpiXQ/kGU7A7cOKrnZymQ+2i1yw6KRXPzoD0wrEtbDi538VoGbd3tatoO9xqxMgW
CdVIrAIFN6RJ8NX9bZWkQvzcAz4l0rsW25tUls8aW6+4T4Z5vspfaHhqd2rg/8qr
GlFwuA7XgD+pqRgKriBgJzid6yjECF+xB19xKtHTZXGzgopWfBuw1CuhkLbOaNXT
RrB7BPpX+gvVv57WyBDkaCzuCw/re7AIsgVZ+6VviIIYQ/AIDAWTaV375o5WUhsw
OwxiiQICeYo7uHS/l0yIpatoKLQQu9bDMxC1k6pbm4RAlcsP2jsCevLcpO11/p8S
qx1Fy2O235RcCjKQm3sE6mraowb4BcTAyky9R7a2J4vXlZj8lcNayEBosAr1mvXf
3IF5p4lc+YcExIlkw77XqnZNAr2J8BIsXw1x8QWIjNF1f9QUKeufm97JYIjbBAfF
dCdoTFKMq6HRJ6hDv3HiQJujKoTdgY6fQPSDUn1fHniwG2BWfH9NWg0hs+WvtHK4
nIgQOEKaDuOzOAVWuhmqht8rYk40G+RoxdQrPzHSANVkmEAmzJQt+nCeawO5eUDN
UArg1mofFbzSD3zJuLWfTuUh3ynEIh0/Y78VMu2p8KOaysrEqv+Y98EgMqj/KMlI
Uo+Le3LWbr5pqyG+NBijmMFkuCWtyHEVUQ46wfOLVL2LMx4o222sCLUx6rkabyv8
`protect END_PROTECTED
