`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fyENn80MnsXNRAY8Z0bMFyTFUWnxO2G7Z9BAy6uC1WKVb1erIwLNR95tsYvY7GCZ
onG0qSB70cbkUELbWuM6LhJg2aHHieBrDL0jZFblv9Dgi58ug3yLlEQqc62Po796
ji4R5HxMvYH4jwP7w593l5Hh52JqfztZwBm53UMCHOxJOq3n1LwSHey3nbYKpHwb
FLfXpXqIRjPfX7wUmMas3QNJfdIDAmz9N0FFBQossMp0f1XkrRxP5iHHFvdVhGBi
6lvGmjuMxnXXFAFXJzLRtOADRW9ZFuZUFIQtdGxSLZPCwQ0sS9Vds4MwSLGjNRRs
YhMwNK2FsLCRFuvpff3eWof/VUfxQgul8Dm11ak1ehS5k2pJUwS+UDWnD++6eMoF
uz1jM5N5cjVzxQqrCuqiQx/S2HJE11a2VA+oSgazM02H9Uk63rnlDrgZP5geyzkb
BEk516mvl2J9cqcPqQ5vIBs+DWQs5p7bLvlbux7NJJZd0sKxez6v/63T5TU2N5YW
TkoGlASnMjD/qwPcCHRVmyEMatU/4gSCbyfVW7tfG1OZBvRUQpWfa9KQrR4rMLO8
L+goqN3NkoukXVM3ZpFeYJHbPqMqQUhfBPIU2NIFPIc18eaZavHPPGcEUgiem1kK
Is2tzC1qD7PK+iwly67BMCpjeIghe5BYhCtA4g7lgddG+QAzae4cFZlbWbGqvgXJ
qk0IMGbajtjy3MXURd5eKnS/GfHuXIBpWQC0pWnjB75DQcBtlbEAOu2BuMnbVx/y
KJe2jnK5yzCUdDO6QAXT1OQaLVMC7KCW0QPsGt4hDbphjFj9KdfPAqYV2504y6tf
eJXDbeIZTYyuYmrZ2Mjcnc9MQjE2LN6DY2GVoJuyjb7c+HrxRr13nMyhFo8HKu2m
FYwBtsSC4ciww4KDbzyRXNmRxJHc5Sn2CEGM/9gGrMzBNgft6pG4PdELDprOt3Xi
m7jmWBC0lb3LhJ+3a7aRvl3qSI/6a70qKD8SaeUxK5x3CIYEUx4rr+Zkz4DkTbN/
TkaQFy9cv5G/AwPDDRRcNxMWRdB4GTZLL8dEnk/3yxE2N9X0y2UMyme0pv5c6y86
6TRbt/+7q0PAH7J3kE7pxFGoY7P/RImqjRhs/8Yg/CGOUOUriCTNG0CGbWd+aQmG
VwGkf6VS8YgxlM5Std1RgHcae/Q2v8YSwNRh2p8IXhA3Ftv7dpKhkaRoBzLD6fzh
J8pnftCWwT0QnPW/7YuZI2Bnefq9vqFwX2lKJEhjiuq2eho+wi+SUjSjTJUVRxef
J4EFCPXNkmtIf7xT2U3DWQnkHJiggaQBnymnVBzlRPlPhKW92hSmc2uJYMHyfcBn
oSEozMR0ZfIIjcdjr4v0atoZqE4Y7y+EOj/uIEUO4HS3TKxJ0xvb1XWWDfl53kJP
E1Erl0/RzXpGcDAx7C65Ve1+9eOCqUfL0VgjC/5YmbZOpWGn8CBlE+UZI/ZGG1/r
Hs7m5RF8jjIPjUGgF25wH9Zb0kzbx03vWN4BOQoHO3qm7SSCnF3zYiA+H6QYjx/+
V2vycpfBPD9ZbiBgBk46JDW2a1NtMrag85orF/lxXYVMqD9fz9hnm1aaFZq1z/ge
p+8SEFh/lHXRE381jhXopWTnujjRfzGg2oscm87YkNixcErDKdWZHdMBK03iNjBc
titaLuBKTTL8gXiw5GKk7xlNlPDh8GOdI89y8h79A/DqIRcL1l08W1os5kIkDHKB
/LOmDN5TBUBLLPslKpuhAtWcHPAIxvGBj5nVuE2xUaZMFbIQzSUxWGVrmsrZtQXa
j6Jhfi7jllHWiuDu83GDOmKpSFQuXQ549TkcVlmPdy1UvR8vpxTJ8pLK7cA4RsyA
gMUArhwcy3gGTDP+UxmmglGjnwR2uh7sjkt67s4G0DhoEgCkf1vSo5w5PHNNmjJt
KCwat/IQ7IHwavYDfsT6biPDzcr6sSZszLu/POCX0XdtFlZZFYVPtiO7H59ElIWz
Fdh0TJgoDe0gellnYBvPkMtin6kqxcY2MpzYd1yu/dF73gyOzN8RIb2y0RchSEpN
0Z4V2NJeicEML8GcxX1P2KwlQQe/96wiupaYQAZeOvH19aaUI3CBn4RNymtN/5OY
fcdeEj0uMPGtiaxmf0q23c7ybLAtMySPcsUkddW9PdqQz1hKcGE976uFx3veqsoe
M0xzajs9ITF8OOKMF/azjKluHXWT51REic4rSXb51yvxdU1l5xvlgMzpjzxZVsux
9hc76tdy2rqUCK+greLTIbDyNp8efYodSlA61duIzVACuEcePAEf+3lCczz++o2g
Sx6Pk8KKt9Q/evnQaOP1qTdw9QZVUibA79vx/qcX2FA0dBdedWW9KQ63KxILc8a6
wUzpShPrye/TtKsrYk8N3dhqxSfEYMDMGuK+Dqk3Q39LozSvJqe8ewcwvej8G7w7
j7bv+oSfr3I/pj08OQGjkbCxlR7p5d4mZTRNYRAH+mxYTM/rnGOhv/nazvmeVQWZ
PjY7/EQRZ3roAZ4U44z7960687zlmpEb/N9OQbB0TM5dWX/hAV+9YP+oRMO2Ykws
0PliRJpNVO4f2ekWLUepm3rW2UgQf9gOwbg/qqIMghq2HrZo9kxOD2DFfZMLi25n
bh+4QT4d7ideXPDp1Gp67utt4ioouqMgh/0r165EH0D/kflC/wSKJTPOMaPrREIw
lG9L/sRS+C7yJow3Aj2tE9D1Lu8TzmYeHLGisPEVsm8hhAWTvd4eJ+zbbhGeww8Y
dkW88X++IHsgZxEwyx4sawY46yM0H9NMxI6D7CBvD/rru3hV5Z7zzNlIMgBuelDA
OTk8w/kb72jQSGGna/7xP2op1kOKUH0hf801ikFI7IZH5KgsJdvBRZt1qJ0ZiEqk
l8rB4EHstVF7vVjgm3FD4/4waZlm4c2396WJle3aFoojlTnUoQmWldVUv/Zrqfbd
d/M+rn+I4KCnP0PxGxFg0RPSOG9wzfp7jBcBPbVnzjqerGmo3t1OUvz6cZn1PRMb
H1wNrtYiyQgN7Di0sy1iFzrv/KMBZsgu4SeqZ3h6jZ4l+DGX5L0V33Pa1AsiNKPO
LlBy4w1kYGvq49BV8Vx5whv5237fnM9mhNBeWwnJyQeh1ooEbfA4nJD/SWRmrASt
9bDh6WJj5gKvySMzGFpPEDrnKlnSce5s4jwx6eY9tTmnP7JNAQ0UXXPgTPbo/RnD
cInUh8A2dqrLFt8BtNRBRvRXWqzbsixTIUWXOr1ilnPN8E7GCmeaXMCciWe5qh+e
SNERAhDH8QFeiQoWgJ0upmOgVW08A+yjiUR3c9tA8bdxT9H1my6bwFn0u+y8YTg6
i9TgCFG7uiq9kTzAvakTyMHGoQlURjaFsQ5QEZakZ2Iybm0MolQafC3ouPRnANEQ
ylbhp5QpbJOaBHN3y6/caOJ/FtkI8du1XQGj9+i9XJtfcsAtB1qxHOTGw0dHDVQt
F8R83efPmzVbD0FzJRTQVOt6AJKmgyohPgM76SSBPipHfPsCwhFn3YR/YHIfw7bj
0aU7uoAUqkWCoVUyx9K4oleo0F8AzPdjpmlqoWv/21HDVM5vDFxOeKItQAoWtAhx
b86ObjKs57XjtPBrP68SmUESUyAhr/uBB3W8EmqKRXiRa5LOoONpRLRH2BRwH67s
p1wsl3PODLY76dfFzSXbcvrFm2Zkj+wQK5LIspkTe0zrBFEO6X/S/JU7ysEN+FCB
OEOI/JsZ8VjRJQ+2P/rTwDZytzYBJFCvjt2wBfAUlyNEYviD3LDqkQ+iijvoe2pf
SIT5MF27yZiLVxvDW8FOkdt4Q5UCMXhEIzTs86evFInASAf6Q1awIuwYDzJ6PDHf
yHQRRO4qIXMf9X/YU7A//3AyngLqJ7HW8p7Rvdeen5Ztiz4e+7ks18ydjmjXxxvN
QODD0lKwOUZ/DIA01BkZr3hN0hYMLw/43iWAODsUUA+aC1UPhgP0q9/aOgaG+Qbu
J6ewTQL4PW/AO7jJfeUhMj7WM722rMwgE4swVelvMBmHO7cmRgggHg59PgZISaXO
GF4Hi/z5JhbD0l7OrzJ0RA9kIrfAXzsdeCpFy7c+xWpblQ0LlJcq0tw3s6xEbiib
hdTnlL8XttYQH1chiZqhiNCqxYr02MinvkQxV24fSFQiBlDpvaoF4dNtkRwxMXtr
iajAtra/GKsSwiTfgW6Voe532gteNq2FNjGanD0XHjaS6tkmbFxTm+NKtelIB77y
OsaIw20zlI/ncUfqMaLLNCaeqYEkEhirxnQ7RWvwFDSxl25LZycSDdrUJ4gc9G5h
0C2crp2Md5kEspAs/BCjQrs52FlQOSMYUSDnIhmhqjKxx5rf9nfXB1RTSDqAvePa
hJKwMG8mpA/7valnheQBSEVww/7XyKVlZE0125fh7bB305nWkOk3bfhm+wClEsGN
Q9ckbBi9RmuoRhG77j2CFxWIZdgx8pi0yxHLVrZIpqeEGsyp8qXDZZ576Q6IhUNe
lgZNMQgDxUyAShWiOECeW7zFytCp0r//s4tI5gkELe3ud3fqoyOGY/GZWV72lkX2
IeIQyGjivzjin8WAyaYe9Vao0y+hYvTfAptG3yM16Y+/EzsJCP/kL2yXKTcaj233
xCEIQbYisyGHHDLz4tQ8db426Ubv++W6pVxwxHGv4UlBlgwPmaEyEG30AN5Jpphn
qbsDgInc+Ka/m11N4gMVDPlyw8OJows5cX4suKZvmkDeZUgMidS5CMW+ainSbj8l
Qy/oR7NnRJFTVTUhYtNLfXmfdnV4bFz7YEdtQOZDYYFFFbGI6eukckzVwPnVPlNf
oHO8KnWURqK2eYkpzBepgh+ZHIywW14hrMKmwJTzJw605iKJhv/wA7vVTnobxNW3
CTuMBiWAvirOqiKAmO4dtNUK6+cCFbvtTq6bItGkAx7d9+vfWosXKr2XsXaELe2N
rf6aMVD2u/BPb+aVPHqKrVaA0tywJGbwAGGTCitsmanzNCQjM8BZI5LjKp0ha/0s
hStsoa9ZfgfmZor8vw4a6otzYcnb3HhtRaecdQggy+yKTRg7QzgYttNuEiaPmKsp
3oU2FG5J6Tne55kKQYAWYyLsYoVbDJejR9AC0gTX0j0XVYwcu9YmlrhKaSi/iRh5
t+6qXiqIiqXLcVabJxvNpO/0v54PjyJTSX3xWDQ+0B8l1frmGgIpp33QoJi8OB3w
d3v8QO7llUeldHNa7o4gpAJg8eGG64NZqagUyoTU4jgrz7oSiHds6u1+0WlqvuBz
QbnqAbx5bzL0mqGjfBPQDE3vG+pjthZkU5gbKsr8L8KF3r54HoomNtzjvkXN9y2X
NUlOXaaMpnNyyc8JLNgdZWLtzBCOdPhgLdR4/EnEsjRB/H/x2PqqZG8IkH2bNJjb
ZaSgYN03xzwZZTIbWNW7MATUZfbRwHF/vvf6QDVrCX3yoT6GxU9lmPBKh1UkGquF
Eff9XCfW0Fxi3y6m3OylYozhOghdHm0949ewXH5X626wE+h/rk5y7dfZJlDxhJfH
rM9EuXilJJ5xRMW+ws/cOTDDKk7HZ5DNFX8G25auSSTfeVrhLo1/zSrlAdY0bzpU
B+P76aQnfwHLuHM2lwAXvPuxpTvt1GEu0xXKf6EseogvIETMOnuJN96E5/d6x59F
T5/8yU/wBefdxjvFP8wKeXjYPDxv1NO98AWMQwMrBB/teX4el6S+b66UdMzbrA29
ritQFOkL/p+ycUBxSKM19mRxpedxwo7Pcgy/Px6udNn1ULIbMjX3C9yzsOOXGz7I
0CPU2bjBrQeFtIv70LFhm3tReF/lD4Dc619fbryynPy3fFP5GwSUISGxFrOLSW5t
vb/7EqbHvrkgXXONcgR/6tU/IcGIV/CL8olRQEpoA3u4+YnI5rgvv90hJopVTt1l
VoPcnK5xFGJzOGjZIx2FWpt1oEXMkiVlfx4thmfX59m/6Y4yjtlCqAHGra0oK8tY
yD8vHJQUCEkrxfmYue/r+gTav6s3nDS285aCM1jA51pLNDkET562omY5sW50u2Ao
qUXjjBvu1YCVkW5Ee5WNVnlPerWhNtJnDcTCQ5oztHWZS8WgnWPrFNwiQ69bZHSy
08Gc+5yg3t4vL000i/se/Y4BtSRcl/H0+REaxuCc2w+sCtYguQT4WW6rdnm/O9OS
mqSmBwWE4SJDYDCb3NKzky7n2RfSIXbR8NFb6pQmJGAFrDU1EET4E686f/6VVwVv
5Pjr+7j2LfJFvs8flRWiAXSb7ITJ+0oBbPxydNNW2xUVBGKm5Tz4KI6AlvSC/vEC
CDZ1Qzz9hwOuR+Kr0DWQpWee9YZL/7TB5fu7z5unYQ7gVLRnFwOT+5f7TGMdLa2l
KJMI6I1oU/+3b27nP3rdoa/8p9eoNa9olPKMbCNU0PU2Sla+aJCm1ca6ethuevnv
yox7FRMi1HVit6NVCG5lG/BY3j9yhoENrhy/0+oQz6+AkIashiUG8IzAouZAkbXA
lgPu30NJAPA5Ixi6yEAd6/FBadwnfj7mEYj6zLz5zvZbPAsVIPcbXyLg/1YIhWGs
vmHk9eFYeZbVSenfWC/Ew4LDvXlFuMsnTdkKVTubKvW5lOfPAWXQjql6TfD3Gbkt
xa6Lf6Xw1E4NtCq6hXXk9fg9Y0GbWaVIEfaMttVM63jYiXzOmNnoH/+4tz8TGJcR
aigH+zFNiaTT2QsByFsVSSmTmtzWhisgp2ggAuktKI/Y3NPvF+nbBb3xrN/NVPMb
ZwR2dNRBH6UhuHrGlu62LH3GeWVVFvIr0Odhhd/cZINtYlKIQbf9wg4GJtlrj8DY
+scYtN8WN/LU0yYRDpm+GGIjjl9TaRBkKfDFaVKrWfVDH1xuUlPETYOPmAvmAKnL
O9/MnvVXyAd02yWY9Zu8OcXkFOqeDOZn4uaTFg0gkdAfAetHkcA+X5XTs9xIeZyK
B2fykXf+J2xLI3omyeOmCgvXoqlbmCiZTQ67arBTdebhFFZwxw5OzDPx4J+E8TBF
solPS7jCETWf+dCEkSqkMXo3J2HdEZvYDT16s7MHRk3OrfJdlPwuRIVwLPqC4JPn
6Dr9Y20OxHlcKDzd6sn1GUVIimhG7Fgbykwpm8+cY2X/5OK6WFoEUjapc7xYfi8B
A72OK2+lOTZ8Va2AQhFo7Dt3ZJ50uyBa3u1H73gnGf0c9NTisi7cTWnOXybvi1ur
w2+ZLb7vV/60852KMDQTAjr7KLa1EhjAipIJ2BRGJU8jK/d0PHqTWPAYtOyGGtNK
hNPbAyKkb6kYVRFKa1gUoTq3XRwzfIAozrbz2Zf1ms00LsAgH9VR34sZALyMojJ/
obr//MbOu0QalPIX5qZVSdGF9ojtSN2req5aQHLrNpNsdD4RjZzJcSO6EnmhCAw2
SSixcOJ7thXTTqP9I7Pryd79LvoqNnMwB8BJ7MNHBKsWwrbd62NZTBhow9dXkJqT
p5wEUuJX0f+VvsexzzszqgWVXKX2k84j7fe4f565r0eWWOzQhFyxRHZgg35yGOXS
JfPp6kXD29MzGiOPotsnhTNxEXKHbF+6Brk1hI48bklMwIXu2I2MPzedCTPKaE8H
dMIUu9M2S3uFd75b/n1GWgiGE+2i3iCrMHpgHobYLrr2l8Mipk5pDDugLw8q/HpK
h8rRD/x93i3+NaLycZvyKUzmrc2weMHv5bJtMzDWNpb1p3aNrwMouy0JdJ85Kx8m
gxuHQXIaokhzw2gX2k73KhWnw6pPWJX+M65GlhLTm7ucqVY71RaqRJQht3HRUA57
iB+f7jpOFLjOLl8Z86hBx/lfqRndSZypN8U0oEjTG5IvIZkmOQzIaSn+mqV82z0v
O4Dgb4Dvuz4DjYV5YpdyBkTJPkBbkVa2ul9C7pgMXln1zWGUBT+0LaEO0L57HmJc
JBSeJJepDuXtb1xDHPswbNHwqBC4DTKc1l1lL58vVYU3cEk+lfe29q4pXclIRX1Z
/834r6I59F56YnOGaBEEcSdyIM8XAzDwBtaboeE2wAsHyGa1pgk2A59cBMH84Bez
Zyr7sBDpPQUZX6krffPbkcQX5G/9gjX3Os2Jve1E8e5qneJ48mMoVnrC6wu+Cqqb
vy3HaamtenPECjsuMmQRzKKq0C/7l0LA+oBlZnoKCEZckYp77Bh6816tm0jtRaX4
hDEo4bVc+6UqXwzhvDW+wZP/0kJwVPLDraRWJhfiOib52EOC+bWtnT3ISdaf8+2j
ulotsUVP6WfPTrTpS/TJtEV/iyHNPjte1C7h4mrsdS9QzojukLKEdcvw0fh+Bsn/
SrV+iVG37f2/lMEpEabu8hF0RFv6dA6D1/V/aClCUCYnjhOuGEnpC+8gRiU1PusR
O/iwCqXBuiLen3kWeJU9QDQ87mzjj5Z5OGU54yNLI6AcMO+9x0QYiWcI97XG4tIf
wINC7tFqm47LrIvfBehEZaoSdNuo9NbMFGBr+Z/Dyhw6m+dQcd61gTMwLO7Lvo0X
i1PWle7vxIy5JHOvvnNhiEcpZRGDtTeuYW0oA/bQdE1lBy8y7Uni/yV3tve1yaHZ
bfJUzyx0plArFpo5QTiqARcnCoh86alOrL7JZzB7PttFulSUwoX7eLZ5QvsjsIgY
JZjKbl2eqaDK3R1tr8kcUC86+0C5DSkysSU50AeA0w1/i3T+WHPVe2fLE3MADPYp
JUGCdugjKnYJhNVA1z5lW2nBGANlgEkQD2Fji4/OHvjeHrcjpQ0Tj2uAGUuZ2oYs
YbUaMO7V0tJ1Amh6zEEi04irB1SKSW4KSjxrAFs60Rn7qPOjc5AVnpmzL2YlbgFZ
ld+7kclnSLOWZYeNuHsmpHAHaJQxXOT41lhgEoqhOfCapXdxfzJUihlfq6dcyf80
jqGotZifAAJddwqXnfWELn+Z4xFrgk25P+2bsX8o+ZNnlooWTUhW0EgcqiMOkcx9
0zUNRjT6Sxo3Y4n2WxwcBIi1DXoOOfUzjLwUR3eTTWYsg5RtWS6IexFI8bFrRVc9
Atct2E3QXht3W2+AJYzXSww7dptl90CXQUeFvDqKhOc1HKecloC/cAe7DdF1djuA
Tdc4qL9CEaYWP4YZ3TLrfANsxixP3s/3umIGr7yYIH/KPINjVH14rC4p5YB2stoV
VOrDOQlBaJ5YHyQwDqWYg0EEfPikKJZPzwKv9neBLCMvPTlDFJNp9qnLJ0pMeyki
Qqlx5FqW5AYuSFQG2Rhb2RrrDZdSO3VQk6Gj2XJmCPyAlh/eZqQLTKcCQRxZLvGy
4KrEDFjlTV7dItoZfbJH9CaA/ttbuzw9CbCKxvEDlBd4ChfQYYRpFmbrE7lNhpAv
en/9EIZqjKccy6IZixntsgdoQjEC54GgiUna0LosRqmmTmO0CS5bV/FG1rlKzpDU
HFaF1+8ES5D4u/Tg/2JKzOjIWlSm2GOWSmRfu2L4a7KHsKBlZhjpxehhj9tZTuye
TgJpAfPto+6NMfEBSnthR+WBNV8tasWW1e3Ip/QYTRImmuehMAO/W1EPVOGkeOtK
NQZyH4kB5HLITIxwda9PIQA2lv5W9wgsKlfQWpCTbtwUqVjK64lJjZ/0rd6knt+I
3PcSo3YcW1djuaSs/0g3/KUQVgkw5S/fecIYoyrCTJ+2zwFBhVvRap530BveXDRo
xdt0s52TyZ3Bd5c01TZeQKqdDxrfqeqYzqPDdGwiPOgY2+Nu/6FfKneX/bRMD3LK
M3rp1xHsUFVkw1w+h5SzPm92HHcve//WwAS6tHmyYogTsYZtxyaTBycL5cdCvd6z
o6CPMDT3hD1PmlPQtsX/Wvc71S+gtjejbjDXdArXTHd8uIS6aV1o00aw7I2tjabk
39uh2KkLhxCnJ21P7hd98Eah9DelhHIPaFjqfKXL1whQvMHAW+DmpxQZvVa90cPD
ks+IZL80kKyWl2q8vO7dbMkENHl6BImrK/SZTtpwztCqEFhKmiaemF9RykVMBudN
R/bSnMP0PxAo7Qzj0OFUNcTe+FO28ouLVedvdVegxO4Dk1HeushRbAMq8QMDP+ki
Joquz7JeoAOP7Q3Nc7bvv4MJs3lPQSGuOCxPtnHMgTL8l1jyDX/zWkfIZbKBN5hR
4R9We9/AB15hvHGALRiy3A/hKmIQX2GbICfe2jynI7Z3zPmt77U8xzBwlJgyxf7Q
MbQhZ3fxl6u7QPJ1BaIpPiq4XwZCU4wj/3wv+0ghdWwEb+IyCSAlnHW80s6wgsC2
EVMuyqKBkSsQwVnCS2S0IM+I6U7JjcuJ+YqUlCbNMw8Ig/89QaIAofpXXPucMrU9
wmGhRO4HJNnTTNEJRePoeTLMe7AYohMqvYoC9Nnq6Fpl+ojSc0OCog6EC16Fh2A8
rDsfowLMCjvhCYKXmutEMowZiwbYpEBAwaBQMgpsxnfeLlvRp2sZkIGrSf2reWkL
OSMJsl/9Aqaml0DQHJioRfvKmeiv8B7mvsCw9bb3ZacDoGVJTd1so3eWlOm5xbaJ
XjdW8ThIZ2S8/LipTPgGesmhDbevV4uzkuk2dsJDe97ZRN26KOhEt0QZ4joaSU50
oKLSQOKCtVxMp2pcvxDerxRTDCiii9Wx7ug8SereuAC/ty2BypDshvfOdeVsR0Fr
VPtzi9pU/VDL8oqC4GLGwXBRYamEnDAtI9ridESCZMuRl1xDhCaonzPKP4+TzZlC
AUfiH/XENeYa6Z2oS373kmB8u/7SWnpqjsFS/YD7Ti/dXK7/tmIFOUoX57UHpbdr
OfGTIt7jbAYlMg6KpcfDGyfAt4oFE2owraWJPOpEKMN6X7oogoI5nA4zxoiVc2vB
JaVCOXR7h5QLa2aJXoNvM6dd0yg5cvQJ47TE34t/xvz7vlc119lE3nfIO/0twDY+
CkgGn//H2mArgDmOk3eopmid5FdboXWVpDMxRYPVEssFB5HK1M/QL4XssfqRy/MR
zXc+g39yE9sf5kMpkyjwpVnZTLkV+bKp5b3L1qCoByBvIp9+FrLtrLQ4P1wx+yDs
SPQYLtApJxDQHd1ycdfUEZ7W/KjdGpYuNQc8sMWZo9+oi56tYm/Cn+wzteT9DCYg
9z4z74RVa8DMK29H8GL7hYi2hoirWV9tWA49JQKc/qJMf9Kc7M2VCR1fYzb0YN9E
wkInaDGZNdn+8NSILi6tqu3il6vk/PLRbdoKUon274RgeGOH4lEhEvT+pMdlmy/t
XqX3SP1wxi44AXA6MvrTrhQqDsAcehgxrI3tdXRsBaeuQzyBpGjm3LkQRrXugSN0
MpJfkE0Ykxbz/V2JteNQ8pyVfF8TDqojkMiTmNpJmZTnIkBk9nbj+YKEGkZp5al7
XudJ9qU9BFi5BP8sw75R+QnKpkoH8Sz5ATdIW4ZcIYYqivg3R4MdZugY/3UWfPkF
3jnGIL4/W0ktCXt/lQXY1i4RNVR6rUC3KNxFV0wzpEV4N+/dCxTV+e1gVaU0gMwx
dtW8duPZcBqnproKU6a6uzVZKvc23Ws/2lY3iPNriar6MBXryMP7xSJ1eRKJDYBa
3ajlRmnx85GIOyudvREbYZNl6fRpDP77NkU6nZSeuOff5YsumLF1U0YKsRoHcbDp
OdBIrAmYsvkmvSWUMGy5fTsu9v/HSLsY6RwX5U1kGWpShctTcCPhibKmas0+wLDT
47GRPV1aR2MtGj+NGGhTkOeLbAtqlOcqi4OclGC/h6bsYhUppLUyA8f2uYTHdurT
bZZ/ubJbkeBzpSvjXUcy8bu3037McN2NPfprY0v64vQgQCQ8yAXCDtbqYlyYVzVy
sEsZE2SqQSYbDyesheqGOxlA3RnMMPMcvoi0oAg0ctk0hxRhzmM1jWRkEEuAz+3H
vGeDVI0p36pMtxzSLO0j4/bQNapDl2LwST5V2GEQhqcyv4+p+GFlmNDaLv3z7HEv
bpwih6ohTlAM9ROSfJITYrKMH8F1hHDTTgh6M0gEcxF0XQ02m083dPzx0YNnDyxi
3iN9xrbwQOL8PKb0PRJun4OgT0XddJMU1NNSNe5plVeSJfkiChsG3iYRWva9GTzZ
O8xoRyXS7L2zS6DJbpvWVfnb5usnvN9E7v3VVmzCl6hddowyBfySMPe18lvhXC2P
Rj+hWZFyUB+i/F8lr+W87MqzYdOPXmKu+PWU69uEbPxPbYINF+sT6/B9VJycJW+h
gV8WVjAfU8m3Vh8BAx1zy7Hgwn6HW15ydcMmOOfF9IQuX3CrwQr7IDEhIJSJi30y
OoF0KPf/PE68f0T/iZoNcuyCbuf+8yxdYunKqN7D3VvUk9/SWB6ySgJ5342lgf4D
8wbhRq/5NY2P1cvFGENwnSvFrWO6Z7J+BoZ+qx3EG3to4BAFcd3SPE+VYxKCMltS
Crg52B+JrKTrdBeYgTCXPz5sVoNnyRqevwos/Ke6GCkJSlswOseZV1UxWj9xLVzp
vZBo8aRklsepGTeqDT6/vIjLntCcbLCRNtYWRfYhBuy1WBgOK1m38iIYj7zdZWUs
Hq+zGETMVnq5bJqhmLUyURY6WkN83n4popf1+u4lXZtX7EnUkZS6qSx9L/XIDqk1
EfMoq6aYoMPM5Xn86e4cjHY/hDdIh0QY7anAgo2TOkNWVHRw6OlAKCclxBhb1ZWs
WA8EON3gDJ/PfJrwIxhwaDonhIL4V1/ut0Ilq/FAV8h5UtE4hHwyb6ze4Vfn0hcW
8AcXAT0QkDUwdsFL7GikTEMgLxt8vh53S9f9db+7JAQMB9dllGyLCKTAoSOVAE27
ZZ2eAPKNVZViNsvfu+uSzEVTdkUfXOBKH7xuksgXBMHFbvnnYvNqR7V3SWFYXtMe
CYq183APV4T0S9rTuz7NfbrHXdqVQyhurWN/HAfcjCq2FyVa0zeUTUkDzS9Hk3lV
nH9GmjtJHcbqOYNuFZ9kvOUN5o1F5YBPOfeXbcORgKh0eJlPMZDsYiBCLXKLTb8x
O3TciYuwppYP/z1m9Ho5ISTegXH9jvu/lklFQvZrlqjhFfONCH1mEZgdBL4wCuGI
0FEAgND7KdEZe6RxFbLWAxDpTvoCtDkTZx3sWWl4YUyZaK2pR3QQ26xBzyVrBEue
QB0iYyNCqj8DqX/RL/vZ/jJUjZOsnbPo53sjABgVVfbYCgloPzc2szX28InwIUd+
9FpbDIBO3fwiPn3Q95EomFIF6J6o0wXitWVHhtV7TrDY70I5vF/pcJr0pXR3UIzU
rRDfG+M54X+PgWXROdlYjp/8+y9L2WUM++GmvYWtDs1QEBTUVeXyzvPvl7M0PZ8w
KA9i+a3jq2+WbkIW+Dcl7ul59BwxUgZ8bnVvVyDa2ugaNSqS14aYB9NDTUDLx+6I
+79fSjP0GjAN9tt4777D9m3UDLSvpEf9Pbosfq0+pVk3uWOk1KdI3Jt4DnfRW6k8
qUd+NVId15DF2EYGk5Zw0+ahgHnyj/VN74T0z4E/V5K1jywCHDGhUoiLGUo+VtQq
LGjzuJlvHfDherDX03Ko61XQtrA4KYYrmlcUxJK6o+Uf1sFTAwnOZEkUM2hkKXhA
xdMU9SSKUkU7QoqKPaMkGNVFerWfvtlHmtbmmQsk7GQJzATLm+tgApRGHIX6IBQ/
m18AjEQnhrO965uVh9OwUxgt1jJ9UG9q2moE+RipUNpQ5ETr830JQYh9gPaSmsf5
sYO8SG77UDF/cY60HOqB1umshRIBpYj1mzJg8YUUYFkq0dK7fS1vZ+IktC7FAbIL
QBgmVty9qPPENLt5pUW1RjEfmvT91+xhZu01jbncUurr92dri7DF1oO0rzu2C/Ub
pLTcwMMarqRIilssDRtteYBS218yX94xXmFFcZtNa36tXIhTAqtALu3Tf26lEDJG
K/cp3QlqsuorL7PELJbfnXaaY2ZAARP2Cm1eg2AgYrY16LJ7s70nLnxrIW+lb5A/
6mOGixVkjlb1JENqpchplZukYggIESDjrpMjLbvI9IR7fGitWucOy41g0W3FtuuY
YB/B31qHNSE+9stTsRiuX3yLjq0BSG4sdux5F6lKh5tptKKIrv2sYtFrQNHvAjep
OAJ57lptvuwEjIeNYFCIHyHbDY24B/Yl16tnTllZH1BI40vV/ITy+1L3upALxsZ+
mEFH4BzlU/dbHXlkrqRQsV9tbctMDTkZD845jjQNO65a8KdLhQr4R3pWfIgA7rVb
wWSqKwMc1vth+deJArTtW2Zn02XDUE0Kh0T+z3X/aG0l7u1fvIxovln7hheL8X/s
9G9CVHZDvdy3HM//hBo3rs4WNiM7AO20l4ZSaqRIhZapl980XohaOCCOdGL+JUgD
gouQIKefunuWno9Q8FXgQPvPezapInbwr+pkumudosAD5lk69ZkpmTrGM1xvO5Ju
WJdWeCz3pJat5Zxvs5PrEc17ew9unlGzICAoIWhioScp11L6mYXQD8q5tb2+WH02
k84LOIUHUcYhYIhbuTGz8L9dRfVm+klRNhKqPLsWoBKBB/OIGjKptLoQkHAdp7Ba
+dNBy3LbQxJ5NNfjUufFhW6TA9rANNHYn2+AVki8g94OAuDCFhVm3Lm443LUE5Ac
6m+r5tiLvG/+3smYlHphaahlbwDpO1QT57ZF9dqcwXTKqOyHCkAMiZtbdSJFfFcx
Ep98SMbIrpQ+Em/J275je3z/Qy8775j/Y+7eHKArqxfXBrOUdO8uq5KBVhC5VXKb
qmYILPcgYkZ4dL0IKECPNSUp2+4kGgp9Q+A1a9B5uvV0dgeExaNfELeNXD7bBnJJ
bZ+IUdSkChZcEvRFvC8N6WGl2uSIE+sdqQAgmV0dVHSXjM2ocG1RfIY24gXMAAZ8
jHdOStjMeYyI0ZNjE0OpP96qjG0sTvGNT+8EGVPbDO4LAD7WeJq6V4q2EW9xh/AN
sNlGUXrNXQCuw6m3KnJvgPBl9csRfALGWTJzMWWzJV+IJG2m+s9E81zJc50HQk+N
9bc3jfST+vi9XW2cB/as4235qpSWHl42SC7FlZ8eHhb77k87vi1e2gOjBRFNtVPf
W74mo6vvaDFiEpsBW7FWdAd96Ili21M0AmYIyxi/w6c5TTqdNweu8GY49Wy+eAEU
ouogSJVESPc/sozEPajaT+YcR2Cjl1WxXt4d2ZMKPT+KZroGmWynnKhX3NDhFGZy
IXA99WPrq3w3YvQ51Ux+LJHxDMe8bZdcNtwTWF8IvQJRSoTnjvrE47XY+6R/oCNv
/8OlV+5kK4vFZRgS2PfpR/VNfL3c7u5cF2wFTbqZM27QMN/jD1MfncMzA7mJrjQX
fgXmQdRywvhUS3/NVPEesZNorBjbEhyyiLSMRlTkrH49MFNaExnum7McnhMaz/dP
HQmD147bDJs4WwIWkh983txXvOdTxaaCw8L9Acot+DmheIDFpF2qrVwaEkgG/slh
q4UuEpnQ/QfdawtOUMq0QYqzDRzUm69VyK612xd7PFsgO0IvOrEbz7FAJcoXysxC
0tur4zyR9YcR1EqR1WQX7cDq/3EOIxKcia/GtBWVMUTaLoF3J2frk8RkPhtzcj1D
FpW37HGdBHBt54gjcQYxl8raq4IfSYNf3Oz3BY6yapBu/ey6nCShHzHsIdUtW6ux
m/mrwG6hVAkFAET0m3OK6zCYcdrBMmt+PrIOpGGue0BfTrlCYQ/EVQ5zoFAmNKcz
XxW60rd1ARruM7OsOaJWOJK+5p9Tja3RGzgmkr3b87jhir/0ZbYYBcH8Nc2WYEiy
hMztgmAJ8hHdwaE6G87iUGNk2uaEzfUwS6HQj/NUfjvFov9C9JqUCOHuKiC8a0RE
r+DMRRGiuuFWuGBVtuwUXW2Z34908Un0rz5xIYMMs+9XTKnMOueZIevfz84i3481
NkRhq2PUCbTCF01Yjq3lvjHPiA4oN3XCP3ft/g8ksZ15pMnAf7Ugge8tAt5/6RjW
Nt5AH+d0bZ1fibUah1pxvCmAf+Qa7C9QwdQ7EjTod8CJxJkqsAKYI/CxvXx0fbc2
Y6o7QY1d3M36WCUo22VvDmC1rQk9a81Ki3qUCE4P5Bs4UBCKw57QMl0KvAbYmUyu
epq/861TZ6NKP2hslb5F1h5V5ayezt55t3U2n2D6QV+v7WTerMonuFDECQUY47rE
X7uAzWyR5CTVXj6f/oRUZXwo8geZzfOQ8aOREFraHK2Rl67U/s3Feu/fCnspvO2g
hGH9JXHXjT/igkdYw4701zkx43dkpxS5y8EeHfaaG37CnFO5cDaA3la3KGATx5yw
4aiCg5HYt3sqtnVhd6s55u1jA03BX/IkQUpRiPxYMVtcTfenK0PpgKUGjGiB+RQD
J5tULiUw+hPzYW9ovDdZV8DqHnuDt9ZO90WpM04i99VedtQBeNvoW8S8c/1HroLp
LFFVkJkthT6eU5cIsWGOaYTqBKKySIVwziICbOMeZqxOdnrSbiuSZeFlpvIX601i
wYAANirHaI5jTZnmv6RMMLP3Bewb7FWSExVnlsoSpcSFUWZsaizwXAHq4s4A6IKv
666hEorvw08mI+cdvoXUt+4t8+AFGWpv9DfSt0I9lyJroykz5RnwMf7cI/fY5tIy
2pclNmv64A0m/dKYfqGISsb9Kg6zci4brRxJ0ShIEHNsDyd9hdjpUomOOmy1CPY5
p7Gu3y41I9hpUTymSrOQt7qk4h75+CQs+4XszckhtW9jGx56PA4a8RYbeU7ZBwYb
sMeW03rVFKRYI1yJDdqp5nyMm/F0iyk8AJQrClOZbwasIiDVf/Fy2O7l4+eUw6Ql
M4Nm4UvrL1URGZrTraSz/EtYYo1ht4RQyjLLqJJ79elXXjUJuyWYirsE8taocKhE
UKKLfL6uHyMvcWQ0iXWLxJ5kd1CV8X2RNj+jJyJ3Jf6jC8tZjO3ki8y1xuQReF8T
k5ITW3uOlLeiUhMW/zYWpnd05Ccg5EPCNnjMM65eA646rh/0mWVgzGjmNzfdGJNX
mOJfNW4u31dy4NIAlfLmAY0cnAjV1AYtcZHl1wW9mesL5aIWSwLtD/qFSjXTrT/4
ChMEqrdwuv8wHcC+LO7Sk1QpoGnY2i215QRvH4x+1QvQAG3USn95LxpfsZTgLKs3
W922CRzK/004CxiEafaPS+t/gnPR6Sfv+mUVg5fT+UFHs3K1PSpZI+dqnvcEnVbH
0my1G6US6gnAdIKrYLSvtYQK+kx/l4KSPD+ViuFQbkPILK1D7XcgaSl/oG9BI/KC
7qBiU+LbXnGnSjkTDILLCEvHJ8mZn72aYzuIZbCAvjkc51/YUehQSOj0Pn/wXriM
j++JyvAd+n4s5PlSrOE49YfbxnSYLB7oQw54UEwASojtUHG7iZbTLRGN0lo+1czy
JWA3AQkQ6bbXD8b77ys20cP0IXIPBh0FpMrHz01KuFLnjUBhmLPwxpZCdOIXzCro
viEECTve0dyx1fWSym2f9T4NagOwjVVQbUCH82nsv7EJeZP2PAfX/gd1Tu2apCZ+
sVQnkJ7/Vs5L8Mqz2zNWsFcpu1UU9Z2kDX9t31Af8kSFCCOXfcDGlxghEt1wruHE
dtDnSM/uBw+aPP2+aJ5xBvlhHV/N+/sYiNPZl+u4p7ND3acBt9tVuZjPGzYFeQJM
WdofnbEyoNd1POv7nOkP3WBpQLZo75jGQzfZaw1ZMRTWkWKlZlhDZgw3JdxXAtgo
IfNPYSJ2sTvNuSOpI/ZI0Xgo+qpb+lHfRI1W717djnpdNQWys0zY6ABGTpG46gRE
ChIRb+skUr/yRyirMfyYBEYhUB7JClJbEhRB5XO58Dek3flJgPrwX1q5xb7WOasC
YWOM2TPy9fLqFkGW6kUa0PttMSK0CVfuHNrabOrMtODR/DbpvPT447+o9vtL2qYz
mLkVn7y1fJsHKrES8f6baf8vC+HvEjnF6op3qv2UdVWAKWwPqSdAlo3a6Sw6napR
D57OSnJvuYlQve17NS5JIe1qji3Y4cfAvxcPJ6f4LrSUZA83n7UCa8yMwb9dO/RI
/F2ecshgiDyeX+ioVDmm87oZTfKNKXyxp22SCB14MtMNoGXaK5gXTQSCzQBIgucj
T9q+hU5spugMj+uWN4d1rQYiADQEG4G/qWAorMMv6o0NL5Ae+yLiXDyhVlezIfAD
x1pSuv4RFggNqjqogZgamJcIitwoTRX1whDrS/p3MasxaHh1e7BcGaYlLJS0PTMz
6JVDdRa0OyrNtG9eGRSFxavogKz4xa53xMk6a5PBoTBcvE7EDY9G8TqhrT8mY/rX
NgqSFKm/Ucl7c+8kgSvGYTtK2QwpX7E7vzXvLXcNJpoR8ltbTk2wn/w78eIzRiCo
3S3DM9VSo6xJUcK/YNHkYO4wSivI4mmfuWPCC1+6Z6J/lsuUGdGgVOBqjmdMA0jl
9tWDZOZhay8BPMmrtXRASFoHQuvs3LgcuWQBnNuM+3U8OR442opb2/e7CyN4/xwZ
KRg6eOekW9HYMSfLqUmt4VN4T0TR73JwOqGb5yGEAZeXWh5KdzUvZ2ZPhyoKU/Gz
jPyQ12bWxo4wautscx/2XAm8aw5nC3vHWYs1oKlVpMgPLqbbpl1pH/T0jnRYF2pW
bk4193sjeX9hsfi93OIH4sHlnENOWmGmdQKXyMoCMeOHIgT8GmloPPiwgsZCwsqF
jWWYHOa68Ur/q8LNWF7Es6XYm3N4sXENmiNQ746AppeqNDCQcX4ZFFbmkB8zJHlk
y1+sZ3Zmj2G/tZWE1oaUCIOhqKDw5/LRtKFJHX4jx4a+v3UKaDi/wR/nnGXJpXyp
4vCzo8Qyr9KvAMhLq+WrlhBZhrXCf/Jzy3wmveN6cmsAgppWI4NIBYHbR0WEsyKC
8xeMMO9sn3ddOb+VtCHsQIUfsLdmK3eIVlcPZa90Sah7xyq5qcL6FJkQlMZZ8Tix
amqHzzDA2DuP9oJilpmo5XqJd/hzYWRlfgvPskLFZ8vEHf2uxcmKHDjo3xOKQ58F
1q7bLEG57hrPJDcckpDH7eYAX/jRrZ6asCIVAogGjdBLNdkhcY15mIZaaKHdCGgi
4LMID3Ru0wk4XenF48wVYD0krMAe1sBtqcsVemXulMMx+FpLWxAW2MFuCC9ZO+gj
07Xn67OsfmLRkfjzVxDRgK2bIoJhiAdioF5o/j2KfnXx1qsuVia2MroNnO2YdbI6
s/3sX06T885w8c2d1GpXtxk0qube31azgjYu9q6A6NZFAFiUZyBP2a0by9QByNp9
qyR/ulFwojSZ1KbJ60k4RqMPuX8gzw9H1koXTrZQhfRPIL/IaJQiN3PxyK8dv6sN
tQYJBphgfliQA37O02tBndYw89/pQMjLw/GV3LEyIQkeI68Bwn1SNZlWTRx6XSvQ
CB6JyvtPlW6edZ6Gd019kekwTPWc6ZHbPdARKcKyVRnRSp8u/lpiKr45drEt8VeQ
4vDd0jG/58Jh4mO/8wqrtdQwdigaL5O9/ccehSuoO6H1gh/hW2uc2vQTs/d4z/9l
/HVwmj8F+xi8hy9Du8B5S6PfcHOGWbV8pdm2n2FqICD3igBNcpZFIXxwK3H5mftA
O8X3B2Utz/XYF7iMIcmwmRR0KL3HDzcGCUcaR4QUiZdfE2ohkomcIhzXHbzvECwy
FJE4vn1mKhK9jcoLksfjcSyzu0meNuJsmtTHSKUcWSpTOM5+Xwh+rNHWfn4hrV5t
/FnpVL4mDgn4Vt4Z0YbUi+Ib4Z54B2XiaRwYVsO0aTEgpXKTLfqFgQYb0YIKZwHd
QvSr8cQ2idS9QhLN9shZ7vURFwg+D1khXVfySHIDIEDklj5plep7P7vvlK0L0Nbf
L8ZXoi+dqRv4kyUrfjgs7gNyzGoEoA7VzHq9ijG94lMupZhwHTVaB36NDJ4nNIM2
HYxLfb1clouT2NNIiJVAINjdbhmUN4x90hMlZHYE+AzJvhF5+Yyl2Vp/HVrO8ZI6
4iDzriO+CYUS4XAGrO8oEQ5I6peO+NV/RgUaD03bhICLR0d0c38WkEhv8DyrF0wM
LboSpDbY07zeN1U81ItxcwZPneZe/0EHIh8rsBj4mhWPETSZyhb6qGwltCexwtz9
FJ1LOXcg3Ip6dQr4wwPq8wfkJcSAhC4exhWcWkb32bLaXDlLCXhctNpskUbFVBpw
HnrasOagNu+tOg8QlaLLlo5T+GveWiww3GHv050xNBRTdIleU/Ei7j7yN2/qzTKR
I94srxYqaUUcd76g5Sq2265yy2OGLB2nzLON1IwYKGyuKTeZpkBhcya5Fgf0A8gu
YudajVtlghcLSsxtLgTHGloRV3nRDLvAhVkyz4DwCCtPF0vhRZj16M2gx4iWCMoL
URhC1Lv7B6nI9mDkgaNDoh815ruDzE/Z8Bs9csn4XI0Q/wcyDVfeP8pbi4gFz9Yj
Mz5IJA9lVkBUsq25wJO+uQKbGI3mnm8/lIK7grhaxlkzXkR7f6G8dMouDY311gBj
ZAeFVT81MltNqkVdCiPaW4QVb60KA4l1TwvBtwFtEycd8ZCEGVIDfhQN3BzMXJRl
5NGg7bDNvwJgUOsGNcfQe6hNSowQeNfHNTM8lhr1ETpeuyqIuGGaMUwO5WyefiHo
MbvETMd63DPh1EJhpjHovv10qVitw2qH2mfhmcA63cHYo2my8jzkjU9ryOeZKvxG
thmAudG7DPS7A4EAxBynUpPDER4HdRlputsPVmDn6wNdYWpEUQ3cOwBxL34O4ffg
x2Qr4m1Do1erM32BoFTTU9ygGEE/tRIixjfEQ/UwJjjgc/d+NByljM2JcF3N41uc
d+HJFfqdR9d6sQ/fT49vZQCiF4Nkli+snAjAqeItmN0GL3Ekc65i7lPVthqo9wmL
hAVPLEuXVgfX6jVPVN5a7KLWC+lM0JOY8jWs1wMSwUasr0TRr4b+DBzri/BxbSjc
9DlycqisX623CEsT++OkLg3QRN/4yzSvlqQ7ZNeJWlJd/BYH7Ji0wTUTtAAWmbHQ
PVwB/lkyJuuQWR2ABdqGz2G75tRTic8iR4Z+SSl1SIv6jvgL5O1yhLqQwD4kLDPr
njhWXV/xwTb47wbQAFGWvHIZ9fGlargLlxs7r6ZEjWBIaIb9/c0qnN8M4G5tSCIa
EtvfFWfLkkB/5pjehdXUQEMfHXgFteuAuwFtosT4xBGGmwNdOrgQWjZK8cwwUADa
z9S8OC2x5qCdsJYfUUrDB/0aRq69iKkaIgCEUcyn3ZJ9r5K5CtI2DR2vvOqAEcXD
4YLDORjp2Yhlk/7LMfl1cBvaWqw6Qp2cEUYarmYnBPhw8NN9lm6DlCKz0iFuWiU9
KdhO/41LabCdI+dXDN0VXELYiTdeZjQSZdImnjGHbzfgE5RK/rE+ewL7YznrLzzD
e0VFYvG3mCCftRHwBEgbKeImN4gbi/KWOquufr+kBbNzXCr8VpK3IHRh0Jnff7Ei
t+kYJLpqPvvS2IVzKxIIr3g4yELmMgUQc7rZHEudTfSiGTAAK8AcBsegbpKL2Cvy
ioILd2MKFsFLgvgB1rEXuYU8eWb8dPcOZ/caIXyZBw7/pE3ZbxOJUbvNAhiA7JvU
nm3+U1lCTJ2jgt5cK0n970oaB/bmu6g86S8KuFY6W3sQPcmxci2oVGqjX1QyOIdE
ewU605q1Eg0n09xNCL2Z+hZoEYhuwXoKz0AxLUA+OfytprdcO+0uJt17h3OX4Wgb
ijCsNvcZVhjO4/6evlfx9hsT0bkiY/IY0VC5i36nnGpx2ACm17o28t3qN/5N60Ud
D2Dq1hhdw7wokL12owdgeOKYAKJA0Q8/5ZBof8o29sgruf99qvBIJM9u9W++nZjw
dEn6j0YIUz7iwiyPW3WCg+Y85o769VebmIZB5FjVQFmSivdfXLsLVtvxUgC28/02
RtPpGg8zkqvYRdue149Ks/k6bULNAiXzyuNkddtOh/SzThUEG+JGrYpFSuex1GSJ
gyXKRsjtBhsvExxPfjt4lP7qkI/rCfWZ9sClKn75ueu9qUeXOVRlrrCeoftta8Rg
CB5Zh65wrDWTolxiw10SCRM1tKtYe4Acy9n5xCrLcQafK4+iJL6Qj1HuU9M0MD74
0N2ODYR9E1itjdL2xNx4dycWgjf9j5W10cjYWdJgt6RNQEcB/6yD+abg3yvV6i/b
Nihbm04tjwrNuHh6D8OO0pByA9xts/lwc1NiEyzO06VUeEhxIOnTDdr7h0q3G/Nr
MfVYvGVLBRvU3sbMiJW9lRwgQwT8hCVuf0W5hAODu/aqLpAL7iybCzBZFm4qlRye
dKPZcVOxNvKK1rdYtjDs0XblbgINmfQHxqe6xGtzsmV+PsZwbOBSos01isMFW/Ig
DalNF73xk/zRvXbgw5Suxlr9+iuMfL2IGJ7JmqqL250cTnuugkfehWovJxITzMD5
DTKipOmBLmg1XDSDrnv/yAiW4lg571/YqMUC29qn7bZD+46MOQyXMqLdlsPOlGB3
s6RPSwBjUciBKAhm+m3eZw2TiY9k0JOSTxUVE+rrg1In1MQ3mOVCKqUPw4TjplMQ
HJV8pAFcSdZeWjO33krYeCJeuESdQpvHhFZivEcAkmVHgnr4lIgZ/mKcwhMpR2we
CjqwGtcGVo7qIGN/hOThJ6imvUtVPBTu4Im0MEYyOx5QWhEXTwqr+eeVX05RR8Fx
zGYvQOh1RVieunZ9x0g4wX+JBY7XmmkWPRZny5sWVybg8u4VtW5PXsegoKeGApuJ
MZo3agnx1TLVmDM49Z9vwcsuGEjdVdk9qG1dZm6Vxg9Q4pIERTvxkxdJ8ZipBR7K
9aJyl3LENI9LhqV38lk7u2NTc314cjHmlDfvjyB0N96ahgwrmo2SDiLfbH1iKZOT
c3/oSVm/i393QFQ0m4U1Gh0Grj9wlHDZzY9TtXp+un7/Ae160TNgKp+Ajkkumbud
LZL2awWUxDxzHCnhVG5E22gJIX4r44vzasRPL3yLl5ImYmH33fuNjx7Ej6FEA6S1
GugATvoec9ZmkDxWxapffiUr6mZaoc4+q0rvOtKuF2K5dIfixUdJ1RBYWzSJv1u/
e19i2bZn866kn12tucg7VihI4x3rQjNA6qe/GgQ35fCq/QDgVGMOKObf4zOT6LEx
WgiL5G0+WKfUPtn1YRmZPBj5q7r8MMHLFfc9/RJ/vTsPU5SWcU8yIR2f1EK5AYPd
MEN1eXlXT4qt5pfYHUiOEOQsE/A8kdihmM4QMJ8C4+rwAEghLnhkePZ6am3ixbsC
UXiKue+rlAZgdnHnVk7UHnffwcvIXrTjJx1/KhXF+7wtQpPMnwkkb2QYU4pnZUUe
jLa9mp5Mt+S/B4KOm0rbHsWRuqImfH2987L5jiNlTLMCsurMFFTtQdeZFe7Auwz5
jGNB4UziKvMlVIpm+y5mGIGn5+nhQtjpupcQ0eDpNl+JjCgzta/lPChi6TreGb1v
tIvT8BzTpoosgK8kJvDv5kkyvFRDaBRM7F6A+wpFplkMNXLkmf+f6LFwZEHgSBEh
PBgtOJU48uL7byPr8tFkz1pMLKQwS9FMXPgawCod23tr2q50tFhq5R1n2anpSFt6
p9h0w0IWf6mCSFVaLwWLZuc2PmfkFnPOSpMErYDl4NrYXm/aRmeoyX3O8dxUXyEW
2Ky69dXDpQ2RteFleD1T8Kd6OXZ2bAw5aeIjm8SwkDDtcscBTVFd1Kr8I8rPDap+
5fJWPofwBpc/RS8e4HvQ6YIgWSfFoFOtJwcrgJuBSY7b8qL4YMl73khLIpNgpw10
wrIx+N5MQtwUCcwOkSwSmfTyjsyp4YqHDvr8IdDu/q3gwWHTFiE+lzA1SWVi2KTr
b/NFeWZS4jWeZ7s9humR/FsobOkF2Ta6Zfpu1qZL7ar6lrVrJZOHF+DOQHXdvLeK
+EyEeHr4x8bHCObYp/YLkN8kMHwNJw2kIVrOoZPX88n5cKDubjZgJ/kqdPbx0KAp
soOg01/aIAgtFAjOBmh/AeCMfp2aJVG6bo7Kd6Aw9qKMWxnCL/xAAEsMAnIP4A68
10GHnm/ABRkU6TYhf3uYgyQfdv5y+ajI8yIg2nAYEe+qdrYSoiMJrgnBj7PpBOSa
Yodlodsa9X8shtx9QZfTkqpxQSTqk0YAky6B8gLy9N33P/XIEAT6UHXIli2ktNyV
gSpKu6vvwU2iexaoV2Ik/Tm87jRU/BWgF9ttgdaTN/KwgQGgaKYxDo1Cl3SrpJtt
3XS8UVkH74BiQJ3zB4uwg/b/2GDhTQR7jf17E3m8aJycf8knqzXS2ZT7mSnYGmft
pMHHSd2RqgBZNj5IcPFTGg6uepxGQWa69sQBwhCkySAreDORnXmtHFqqgm+qgH6Y
bw+gg6lYs46g0tCYH7XzOeCoa8BnWOsNqSh1Df0y/QQrFoHIGh09CM7Txsb9qtQ/
rrRo8HALK6ATjiVLP2avQT7o3WftEfPqL6aR0ZfJf1uUM6dShpfsoEzGuP0ssYz6
tK4iDr28ChN76lIZGBvY9SSFhds34PLzeUb9vUvpBacIiShX3flw5Jo1PxPmgTjd
XtWUks7udcgzJcB5SURxkiE7NHKEm9Y4CjH9e3RuJfxcSHHGCGUoFIZfHOE3K0Ig
+va57je0j2lqMnPne3mqF8sH3Gk6l6fOcycPM03NA33cKLBB9Qq6YAPfLWMPQVOU
OX1/9jUduSx987n4tWARz/QKcR27sMHFSJt0r7S131mjOOjdjcooe/9qx2uDb05s
rttc63k49knbbWHOj3aYnMn9X7Y/IT7MYUATXJ+R6YWqSPKBEUQr8LbEjyFnqrL1
UrcBJYlhkgqN2wCJrsTyGuRl1UNhzg7rSIV236RlQeJyrLjSOtNN8wo05xk1377m
G56zKKDSKQ8++rZjp6oG/SMCL5YZUWwtF/pUAPobjUBJMdXJE2Hui9A3KNEXi/Dg
bfM2yDTtbEqoZenCbPRmkHygvmtL+uJ5NZpDyGY8vo0rOMhssplXRqfe8tr2k/TY
VHAahq1V8XdEIstFnZxC283Cnuoefsj8Iev772SuV/NEMUFoNmxkLOHK9JuitrRd
Q2dalUmPdmc94pkzMhwrjtsQ7vDdewlL3hYSdDd85gRdQR4vpo1rPuygOG6NdX2X
G9BsGimg8K93HEm9b7+kT2WNptgZzdhjmRdG0hxvs90yWLyfRehK32f+ADx8tofV
HwfPjWlGta1OmNZeoop5P8q28uarR17W4cLyqUDZkPjHsrHZFvrP4FUWlQ+gBsP7
P/6aSG5sO+mNXv2NYNj2dUTu3Iub9QSKS47VJI/wxhGy4QhpKZHsjXrH7eI/uXqy
nYiCWfC6qGEICrAjgYKn+p9el1p0cbKwCsV/nJVZUnOX47n1P1dz3WznXbambYdZ
JD3a5oJwtGuTInOmVnlwbDfJToD7Dee8nUtXsNgz9Xe5H1EgIQT0hkvFkB3Yq5e+
Xe6l9sZnC7+KecxW6Ytl61I9ToZpUrf5n29fC3/BC28JnINibw+7G/04fz8XZzM1
moMXYlivCq31c0SGbRO7eYpxlOTD6hv98p+qFOPLjPbgPk+2Mf+3bxArug7aQkZA
5jzn0W0hSlEx5pgG5ed74tZFJg48AjK3PdI6NLUTvLN/xWndJHgpTJyWBXp83DjN
+/P1xnJ2tc0NHrCgIbTrvLNgcdMP75JD9N8ySClr/xWZ4CApxnOMfkxEtASg+zMc
4iiyRzJoOsUCbk3d9+XU9SSNKp8K25L5g0cP2ovzJWhw7Nidsy/3G1wsEaaCKtTT
jI4c6xOdKJNX1VM849r3/7912lL5yGJXjUhIFgbbpQgVabPvM2m0b7N7YvsCfn4Z
2x3OGMXt/rC0M7RQFUNUIMWQOJoH4ND3XHzeMLkId/gy5ks9gQgbz31towg4EFxp
ilaPFdZUd394ldRzmhaAKBAUr+O8X4su5MSzkSgDLdDtDRNe0xFUfoAJS53gsbhp
0iVj7npqCknGElKRCdacktWzImhkZF/e2tejoetTjrxf6txNRLvdJUUv28bA3B0T
7YK94/CP+HVS5ii/imFSesGvHnYvLs8zLgNLAsDbfTrL1PcpSW6QWReqQb5e1BC1
wcvpGpTeiLT+LQgeC7yG99Fs2mMglhZMKBhGKL8ev6viu/j+QWYU2eATKET0EzlH
KrI3w9a62FiK8E6W2P5rbDTCZsLRnCcqpqePkXSGctPJBo8vj7GogOGJ796KiPJG
bLR86i4Q8zvZt0xUfvNFwU7u3SpaDOStdrdNWiVL6kjR/+M+hTk/TlN3BScW/oWe
AL0KYrllgIXIm5KvjJzZvRg2WX1tm/6yAdiSDH+RBsoJv/7MxSoqLAqdLvh+wXxI
Gm1jVvCXpuWM0n4O8y9BUyOPAH6Cq97wIjP/+APXl0FjqmrLFN4FL8/Vk+VQicWR
PDIuecvR/ZyNNPul2f1B8n+Y9op03qZEK8VSuS0r/EaRISs6l0139AwOvdPwL4On
pX7vi7a8BBGMrXPLFPhUXUT4hqCMPz8inis/W7BfKykT893MTovY6tKlms8mNCBh
g61JzEjpsxEmRv6BkTG/Sd/2Ksoc+zL8uFDyXBjJ1+akN0Q/DU+ZOdyoKw+T/cDN
QisQ1KtFz4gJONZ+3ren3CwFLyHim2O78Mhy7u08y9IyC5ZtiJy/X3BL4eVVjN7f
DUmS+nHm0WSU6LOuO3kkfOE9NuxzF+TAy9EZHYhGAAAOwklUBPc5DwRvLJVShfP7
NmXBZQ7Sk5Sxv7eq1pX/bo0sJkXVgaVcS5lzwMUZ7yVLxtSmIJBQPJO2AnN4XsvL
RQV3RyIxfiRJvVROKzRccRKGqWYpxK4XD0m482oZUFheAuI6SZ4qN+MsmO+rJ7kd
RtvEv9MVriiU9V5DRATgvptpsURz1fbeMIMRbldgLN1ZLbiN/yiPoGWLhkpEiSNw
Ij2bLPueiknSDTJOUBdaLm5SQiiFo2mjS41NuolGWvkha3guOUN+ECj9dATBj5OE
4LAGPB4dp1NEFrfhGpu8yjfcnHdPOA2xleRsGpmAKx7ymHBmVT5Fm0DMIU0rSz+Z
5j/b6jo+sF/9ozqrAF9/5KD936GFLXVbwn9rQYbxubn5SKhZN8FLw+K3DL4ACAeF
Y+/q6SbRIBMsIocgHp/9Bniol8MwTrjfqt6L7XWxJME5XSIiYBoYTz2RwGnZYffL
YImXrkxqqBCDSvQ3p5BnD+wMfPIP7VAhTvF37EquDK92SZjZfP6PggdykeusV87Z
Bc1gx4b96F7qH/F+ajHUSqYxsKWLEZcAOcVmKRFNjs0Rz5LUpiKl26pcFnEu7biD
q/uvH5gtcxzCVV3YUXp8dIDitVsAPGtQ0NPXTFyPnv6L/LzmTu0AcJklOA06jA9C
mb/lNTVVdoYmw/uZIv8J9lsjFiFwqn/MEFxrSCovF6A/7iirX4nQZXDm6oUFGDFo
xCIakI1N4Ltx3Qu2sR+sbhEr8ylipMQT1nGldNnCrt6uODF3aglaekG9tBsJrI4P
g/MxPZxrnMFkB6EQ+pL6JsW9DiM/Wix8K61t9pw61omXl8HNN5UQeFpgBLfbjkFF
e0qmYO7VZ+Syw6Z0an6RT7aUH1zcCAAaQBQKK5M9PsNJz73xb7U5m5iniDbCHg/a
F1/zGKhZhfXmKVuJ74ZaXhouiMUvqmjW5v5813NbLAvPN8gQgImFN+9ZyN3nrtnm
m2KV/dgZaRNpYySB0ZdLF8kbpBGxUzLK21hRFiTBWk9Stp2+FIbXRqW2wTQAE9Hh
+ticsS0AvysQZ6iCAZPlceqjk9QHmYgpH6wycWrH0qWzJrbk9mkOndJWK0lXTtdi
ahK3Kd9iMe6mbs8ZPRTGqRKHpoz6u7CrqIRn9w9iLUv+RvQYgprwDETibrbQI/h/
NomSdgbnh0MkZuNXIDXWyUbF5Mmnvuodso4GJSAr3SuOqANd4ykQEy0pprd0IJBj
KjuB7LvF1TyMMHT59d4BAcN4GwUNUjVskU0Z7b9mP/J2PprEY16GNsfwbSyAlLY9
iFh0F3gl27GrgOmiaLkMA09yrzh5jHbxFOuj5+0MzD3Q1t+4NMwGp4mUZuoY181l
SQshFvs9UJjE0FHEu09JM0yOzbFQhQ5JlONf+YEN0yxmp0H6lE1CsyC7PGGXYQgL
HnO7C4Phj/FNE12uB28drFFljZOdpcs4aN/1heKpbMKS0v1vV9YR28AXh26HV3Zw
ivg1NKe7YWpYsEbBRJbnpYTw2zGTgbhyyd11Lk+garrilhJz9RcyIseuBx4THtYQ
PHw7JKT62/NR+zNojgc4WsPS8wtJyaHRf4JnAnF9DfGuywE1Xz1tgO4NxSyBTnk2
dSSoFdLsKPzJLmkFyppKx1PYHtOQLWG21vE4SG7Xg5RqmzyFiJd6a1Dx4jQD48TK
8mQWCejRrkaQKctx+PY8OK7XSgn3BPGEqvVXnBpcFBL7TjD9V2FDJ7aYGQtnvvOl
lmJGVqsAgpNvwCf5SJrHt8x65xSfKq0+ighUbXa19yCdxB1euvvDq7xPf8s4FZZx
A0Zc7OeuQ/OY9dkI1BsiXx38ICTVIsUbmCLXgG78HYLG1Yj2utzr0+UiuwiSaa6U
YfVX9nF4CynD94PDOUUS3wfG1OI5u5DYwWJmU/Et/OuX8Ir6DZweMoBs+qFKSQ5C
l7urc217wMJxtAhFkXpsBNc2ET3d0QQ5cmPlAAXWNDDPSQ71p1UJ7c3bCpYBTSER
19Cdj/M16Ccm9OhPLhAWSaFR9NXgRCLtIYXQqiC071XcAoCSS3YFNE2LBHaYtWM2
fbLV9/LM1gYpqOBn3rpgSDEVgR0svSynl5jfUf+YzhXSP7MTDnd/Fvn6tT659udt
zfwqaVd1zchV2VGkygtxVtmI2omm7AQL3g81zkKEauXub8Yj53zhQEp7hc7E6S60
WKbAW6Y0q2qDdJ47LLl4wZ8YH0szuzyebktbXSxKS4bIBU4qnyvDERKSTUU2dCJW
eAgnm35iXNsYIzsdc0Cl4cKx1dS3Xez/kRAJYw6zc6UQpzjEQfZtPDfZ98bKRtnn
ve5gtN/1Ptr4JkTAQmY60jJXEtfrScnnWvXCninKcjnblwdYP9aHdacybYpkSo7F
puRxlJigAhbxTg7jXEOU412Gy895PC0y3rRcDwRXthxUzvHC8g0xMTUYvYmHpiMg
lhvq2/tvUlRIddXSzqmmXp/yoUnXG+NO+xI/D8AtwSbnFvZVCNvMyV7i1q+QG5eh
AmsM7S/HiulfCf1TpC7JSSdAx6EqgoXN1vMqcNQZouqftRQNsHiZfoCd1dexRcoD
NlP2Qgt0NrYl1Bb6hESgAIzRSeihGgzzMYF/bwvjlewOrNGtJ9mMuzfRwncJUgBB
t5i8G6dtdlBNEn+wXbahsfQXeXbrVB8yfsptIsgmzKG8kHlUFAe9jJufS3xBu6lz
17OFgudPUmK2hcFsYhdqYKMetv6Zz3Qq8MwOfQD/XgeaacycpDNU7U7lWVxwGQ6C
1OzCub3iRf0NjPGWWV1aXYMd0gJpnPw3hc9wMU8ylwEhqUnIPKtSuOS5hzuC8vBB
+CH2ygc+jKvIXe2Rt9BCMDWjr+/pFbgSE+BUzan0feNTgHOvLfv3yHdzx6hzINoH
NpYkltiTt6M5UWyoHP/o43BKGiB+BJ7RAsfI2lgDg/hM3OgowKIb4VWogAPHK0E0
ti1Ta1dXZuTw2bNzKZ5BVyCLlsqMxpfiWQ64JBtwlIgbPaVLCTb5zoU3AWDFuaeC
GMZpkN0YCmXo6WiIUyO3Nr5wabwrWPh7CmHjruhrhSPJbCfPBEOA6ltZKzSCRDbj
zMYdHm2GV57PYGyo99Di5c7ml3CogExQ29GjiSvzWnjqc0EBfMSs1covQdHMLdKb
nAoFbr0X6xYstNTDaG39XvP/dmAc/apsH3H+G9pyvcEIZHlNvQlGBkCgTgtlGDt+
pDA3+Me8k4QNcbOyNXyLVQ+KEmQnYaYfb5QUchsDZ6N88FR8bzOTIfsHeDCqN1zi
kEJCRHrFEG9jP+Fo4XrBMx4MnTTlPGhIp/Zw+an3tvaUeg1s0NkTmGW6H258Orm/
FDaEszi3VOChap4Qu/rfoPmYH8gYG+5jQSihpJglXKPubYAegBIiKHFuB0pC36+M
O2eKTZVi6D5itT4PoBhFKK86iu9G7EG4r42XL4+LuZwdYdTHmpQzXiwpT+3xmPub
pRpu0NzroNdXkeae3aLe/WEz970NV3swkqIdHvlHORAwAy3DWsELZL75NbTmkcKa
YshV6/Wfhf7DEDMg1NV/gowWy9sWq78qs6BoVcq5t3kkvkJDY45HcUYdXkJ8PEpp
tEWSXDafi2TQZqx2E8NJY13wnDFZ+by9P/c9mWzrboKX2CDYq0NW7xRYa2+SS+g5
p/FRXBP/8qBp9c/nLro9IoElVvxI87Cu18xgeXEy89bhcQ2xQKdcKtsAkPIS0qqz
scRAa/09pae4jgcjE4Q5j6qk8d7sCP/EQB/MeYsXv2nptYhN9UbD/hHfezSxgUJ4
JnB9CLIO/5xZYEjv7r6N8iPUjJvgwx3xL65dFot9jOqR9T8UBkyZeryuC7KJzBxO
WtiY1hhamA0EUqheBcUQH7swhXpDBTRXJI5LVoFX1vSyrP0g1nMrAbBhsJcTdTlg
TcIN3MCYRLJODHFm9AMx5onPkHs/TpOJ4GQymok6gVj5FXlouAvDGCov+zO6qhcw
KgdMzsCdGGfwclGJbX2TPtajAjVjWwbk8zMCUH5n/KXV7MAx7Co0qn6hUVQpmaOe
k8pYGgI0ISttcih518PAqe61VbKaymUI3hge+UlokMsm+9CLgU8NQoELgHMxz55c
Fp+0QUNo3JTl8QLS9Z3QCHrenwOF2oK9tqaneiSEJcsfaCrhOk3vtI2d1JH8+tMv
PCtNmzm22PFvxJ79Qtlf7rguWFejYsVoZwSVBbDZ1QiR6YAOt23/wxUP8eo+XH4o
+qwI4P1BwbLu/DBO5r4sV+VUrlmEPRs49uQk5dlWckm5kfB+5WYjRw2pY8K0jFAq
KsPxCwYleSg+1uLYXofiCDMumwbtl3El5xhbNTGwXNIcRwFhuU3b3mzAL75Y/qTn
yMePKdPSc8hVKUs0mpts+4uoXyZ6gIkot9ne7LugkacUYbGEmDSbMtRZQ3e/OwYX
mhQbt927Cm5skMmcMENXXYBCtZyA/aWni4G9I0bISI8gPiM/wIWNPXb2IUYHTxjx
4kCZckWPao2k7Ldyk8wPpEY9OLt9hDevugXPdZwuQQUhzJjOmMrK9igcZpIbvYIZ
GUHBJR/shwtvB9U/18bJofDhNQGd8oQYyZpoWtmswk8O7wPIFioSe/LolZKZXyi9
wvPQtCpOC2FrrmuGSedYki6ha+MjmO+n+3Syt34HWLMpr+zQsSMdaoKTr9YA8W/l
HQp7cxTBKIxRtEZLkMNzNttQ+i/nJq603EmGsKlWSk2JWhSZVP5qi+vvrsLCgxs9
djB2lkGbs+8NwKldRXWOTw/UUjbY/0WxWDz/kB+AuX38Z8diaP16R/gkGt3PjeKV
zudFxcSDYbi2zsXuH3u0NDGTHAYXQoOgxQ/WFd2CHvVMcMacsKjKHD7AhIP+zGSX
NKIMlIz7a8+91h1xnbD627NlM5ssdOdBFpftLWKSobLXSBPIZSNm9SHeNA0N6U3c
rXrNZ1lJ1gis6UjwWAgRZF+88ajk5qnLfQ9IRYYOtCax9prnezZ522T9wSg+fuOK
otmi3ee0s3gr9Xv+53MbZ3Lbzkz/U9cSPV18q171sZFQFi+l5EDg8caouMxwgEJZ
SFHJTce9/yrR7LeWHDoS+9jraggzH5LaNMJQ9zdPcS1MZmD1QOano9Dtc98gTlHw
LMdtKpqnQA+Bg0I/YYMqZLPqTANe+FKMJ4Tcr0J6kGFsFYMQcqNdsohFO86z5pH/
3hO1wf+mq+9e5MPEjddRwI8wJ7fMCA+UoeCWKhUxF55hp3MOyJcZlTuOKtdL7Rh9
pku8fWnFrPXZ86E4YzqBmBz3YbB/rXVT/PhZ+U87sAiSiEUUNGpMm6gABTTWmDAV
tfDnh1ZUXsg1IJHi6EaISCxNsFq/IZkgvTR5CuQauNLwImlNa6il12GhVocOLkP8
L/I07yzXvMbHfZuuR2m+72mExUqxWKD38UiqlXCk/wEUG8niZ6cDLVzSOhZt2Rd4
Jte4ZhP//pnTEC2lTTOdimbIupLuYhCzdg+K/L3XcaT1t1k/xhjn6X8kAhfObWUr
pvpMDt53qGdo61JDVAdabiVxMoWdfYa/KfClnRGKWbxiqal7x8CW3nzLsdqQ2lqr
t5/s5VC13JOZNDDfHvm21lp84QNsL03a6zItzhWHf8reV8rfmpaorohsvnOuLY5f
odrGQMgZzrImQmf30qPkogPn+zUB0bugiBxB5b+78t7aa86d10oAWevaCjQjtkRi
x/YBhnHcjceGU7t7YeFozJfXvXjPLvkLP5zPafcrqowZF2F1HDAzNjaO7rC1dakz
0z693XXZJ/dzAcpTuJHs9qnmMCp7UfohPm8lAt7d72QRBRGpn9jDrPxYT9J0re65
WPMZNVRDR/JNqg5NcMq8ul/5YXzio17GJPCJxGvW69jyALxKC5y5iPIaJtC1Omw2
JcBUZuYnX2iAN5O4jCN27rpGgiqvIAfRmAXik0iABT4uIW5iRPCiDBpqpar2eIXN
T4+hvAPO97bGtVn1aY12cBKx8iIqr0MxjxkMj7DtbcF3gc8UMQCqW2rGQDbgHq6H
ujCe3zbfoCsL4qiQUNOzrhB0MknFyv1chIwgNQs1Hn6k0yjihH0gJA6fYxZy8PVj
hx6KHu3+nRvy22nTW7oya+SD1WqhkilBJhtX9awAtqxLqy5QZDdrISaKnGF+O2cO
j5O1JyDGSXcW59w5qjKBSRHIXyTCBiqbBSyhCCODQQBfDUJbil49kkawF+bumVjK
KdYuVw5CHB0uhY/k6QbxnEQNkPWhM2iE/53Ra+n2yxh7UL8d2XonlKyE7RMPd5JE
NHgDs7yyjKRkgBhh4/imqmoZRwPvQ2F4OWgwKj6Fv19ZYCcC7+fu+RJLm/J/FoGF
XJWh62wuaOWx/oA6XUIM+2hakJMsSGLtocKeVCqoDqm82DatRfhY7INRHmoxuqJa
8Ju5leDUZTRyi6R2asP1wDaTkTTW3mcIKbEx2W76BBJc6G7yLNgBXnTVo0zMSiJ6
Gq2Idd5lb/YG5Zr6gQzCHWuNdsBPARsoq9XWVx44O6s3Htg+WhsR6x/o+begvLyn
hUDfGWFM0lDFYVTEHJYKyIEUkHMeS+3662y52nB+Q2FwdxQ050KnZ7UuXsplHmqH
vdXUlCSwP+Os1TZCiElZ1vQkuE+4+c+8vRZZI7SPRtRMJxKDFTfZN+tsh9Ir260x
g6c58sm3eU+DaImP29ATLLKBV2eMuLDHIzBPbh/fu9/XZnXiEaC7LeB2qaUS0LWH
a10zMnWL5kGrm7XsVw783gjAOCXngsyXzf9dufQAlWFWvvkcWX7lb4fRzI5ZoB3E
apXa94HS5jRymH3kBREUn0uJextDI96PYId6oBS9OUWF83Z7noaEsQt8/r+oB1pC
D0s5/41tt0b2RJvJ/moAmNWuMiiTEKqTsw7a0tcLfX1MsxgEdFu5xgvQW68aB8Qf
Fgf6JPrF6e846ViHzMcqlciCEM8fYK1NOq5bBl08ajlvs39eoZstD7on77Z7BoFW
SwrZtXzby3QhFPaxCxQSIgpOWl5047CyyDejOO4cpcS3zzwfpPlnJqyvp+TPTNc5
WvnGK4rLyrhLl3CJo1h3YDIecp2WmyxCsJqGrE4q99ZjkZ3LSDmkOzV+zJBtZEby
VB1u+0SD5uZDn9GnUJp4FNMeAxEi0Wi12BoKVizub+dvX3coXXJ0ZQ8/FYfpen8K
EBto+J5WUAlVfEci9FQ64gkRqoGqNU8UqkyLbZuMzOqln1FOkCZK468pjKuu289J
hRoSW/Hg8rzOQszuNAKdjKKZfn2mzQcQlhlkcPGkSc/TWOFk1qQ0sY9Ar1+Dh3XS
72b4D8TVjeBzzQPQuk7iJ1V4Ym/kiQ+EUugcamTvwX8bV+SrNLn8k4M0iNvvZEod
NX/bZ1vwM/5Z50rq+OQWwZSgvnz/q5n9qDlGCgHX0uJOhqrurHXW3Ff6GTEnPWKT
p8/GVLkG6uYyXmjNhTPIFfQ9mmkap7sqobkSkJ3/CIDNc3UVrw6dkD2MGUhlWl3m
MPfZSjRiHLsb4wabHudnvh84jLlhyubJ2UKXpgwBEM8N9ZT8Ri2hA7I8MJ2I0czW
ugKlTgbO3KijyfrnT18/jS6JmpetpElVvJEOw/+zY+deWENkC4g1TKhO39FeODHy
Lhnop+eRVMyKsew4X9NVYcWv3QyrK4CmACd4op5PDInc/JviO2Y1T2MPELV5Rnsy
esp6gria3WEgVn0OHxRZEIoodj1QuUwDWtw93s+W+LIykeO3fSygtbI+1ZMRXflp
F1fIqTlZyHYE9Iy6D1lC3U54a73PjFkPgPSv8bbwSNle1y5gQnX4BCPIlW9qSwHm
ZkkI0Y/5KfLMEzpG/7/snHEdSHmFm7YljouTLF+ufX/EU7QP9+WxcPWs27edNM72
LP8Id0Pbt5Vhdrhepy+jlDRkJYHzVl3BNbI9+SMf1ktT5WX/gGXubrRekg3VqxNj
4rXPGQJzbKgggUArixTNmuX02+RIINWWcROp94SQKVsdscXkAt6ulwoUpZv1KsRL
bjgthoPwmOcNB5pqSeQiRYDLPJgtS21usOKzFaKFHz8peU2DVXr+9kt6Jfo4Z9Ow
TwILVnGGGgs55uG2YJMW+xyTpc3aHHCvVSpGAlNTHESBi/A5rCzbpZgFyCTdv88/
MhdqleD2ut7/0D77RDdca9lvEFC/IUYQpJ9jzpB17nZ5Ckt8Gm+tmA1Pe23qU5z3
eoOB98Fv1eTHVlIx5SCGDDXD0vHMZHEq/Msq1bNOK5nPo2hCKVNHHkdyzHw2LwEH
OjRO0ccjTgSwdWRNblvolK4kkKAsdlTZ/1BL0JbDrC8OZbaHEaj1Y4vUu6RtUo6C
7w80lbURiOPRFHuipiEZWU9z5h9TIdOYfv2VkXNBK6BDPY6PsknuuS9qtD1NWIs7
RfQBEkcPAktoXEQE8Yetys4FGhvzTT4rgqEh4UsOcM1lsLwZ6SaXQCfqAmr4pqpe
OE8g6ihLb/fNKsgI6sc8XxDV5KVbblJLs3tUlnJqyI92auUsA0CkaCpTpaUeOlgM
f5g1xg5VerJvlaGclhy/p7iFnLov9qamdDr4QusrJFkGF8Jrfn/RvLvkKLzCzH4f
4bPRTeXKTATyYO8nIYlHrjKdrq2xHyRwGHpJSfUyVENq1Q4sJUXWkF4Ur3M5VwRB
9davFT0Z+Tm/wfj9sJiHx7oOddVJVJ3R0w05UkljrRvd7zjoJLW0hgpR7q2j7KRM
w2/hW5ALNS8tQzWNE64MM/bG2WH+oOvwZUAXORqind8zIBSTItb2fEmu/fpuQHN1
+9VbL0KcX2XHv4ht6ZJugoaH13LaRe8Gj5IbmF4UPSCdbSPOYB26NHtMLgxo2+yU
UaObQfaPK8E4vCHTp73Ve7qbTaATLrrb07AASN7P9ESZ6kRvu8qTXU5ZJSWO+B4b
qlO0RtLQraoXxRmZjNOlQmS7HPzW9KYIY/lqOoCuqW9WbEFfqInsN95xVRSzRDhj
1bnkWDwIB9JIccDr9M6wGGel07OjIe8gYxzFWdHMcHKnsgGYvdCbwnLBIMttxl4M
NWOIg5n8+3cW7+wlcm8zqyJBb/aZr9CA8VILHZ3j9Izxar/O8GgYx+KrYgKS72S7
XGZ42IrEoFLsMAVJkjwm6D5uJ7GXUItRbXJAnr8Enzck17qM9NpQpd4nnA2pRbGg
8fdq/FwH7ED0JfjS9umzKrsMpPsyiIUdjpRHZBqtqHaZGtohWZl4lnAE9l0he2fF
27e7llOlbH2KraGx5AkgD+R7akbaljYV31t0KJb/wWzvxBg17FrqkmgHKE6+GQmZ
UuecU0cGdGsTsNiFxRvOVbt4NeRsQOic5FBH/r9+0MWvi5tW19COiOXkLaFJgtNH
BRvBaU8YoZcltk6IdLeRO1KIb8p+sD7ZnqV77xi9s5mFUa6/RazMBFXoin21rmaO
YbtH8oEz5wm3nDhguhhIQQSanVSBYuS+BPT19hg42o5oUWg2+9mUKIgcG5MEJX7l
qlBheLSNcTNHt0MAcot7GFjhJKNUCrUTaLpbCBtYZ52d0pQ4ckFPUnekw4JELbBB
+tNI5fjg3RbUeurgu06r900lVHOzRMR9OwkgEb+ikiuE1zBcNyDQleB6pGs3E24/
35EzFVr0aPXaDMOD7Ig4TMWVUA6CQVNAvLc77TUP6ysu9zyzWAItTGvOPqSR4ATf
/j459AGbRk5qrSqrccTmUquAq0dAs6Q3G3mYnS3YqsvncekYv1SnQ+/5OATnmb2M
+udoXurT8mj426lcMQiRPwbYLjgOKV5/YwaoamM1pBCFUzWQY51sqHxwam3UBzwK
TFbe01MWPbdOku+Gyq/Hr8l23dBy/uQ5ERNPihPErH2FSpimf4ZiLHcdrxlDEZvW
mkqbrksZ3D4y59gbrAD0Lg/OKTcHWGItB+bwQUH71jx5ZfX7JbgU8Q+FYrdVIpl4
bOv0aWAFB/B4hM984aLGXqB3pvbEhHw8HHXxC3II6jO1Yk6GoP2eIiff2ZgnSzbd
Pe75yBgzKe1d56+QV0OF3ps8uIu3ewl5u/qKD+QrUKO7371WclSS9Y3yj5gA48iq
tqlpUGe41biL+l2kZjmA4IXzTCZ6EaLGMXVMPs4t8EY0jLZyUPigeZIekEMOPgdC
35iNbKGTaHhpQf22F3nIE1fsfZ7k0T+9o4Oe3Gi7BeacGzSD1W4PQAyeDOS4LMLy
Tn5V+DedwCv60eRMi3A/LAdvgOYTiKBe2c7NNOJOyAsmJl9JWS83/4Ej9sePc7P6
CwVOr1axAb8iwUd6fNoQ0IRx3libw8aOrwa/ooxGO6LDLlZKdWoFo7woiNccTu9Q
ugcIfD47QjvksKdFoPMK+kc0B91vuOvXkkcb3YzHFR7fXBd/8aDEp3P9YZHVR2Ls
wSyObWbmua2F5Nbh8R1izKyVEO64I59SiKYLLwyVcSyzS2boo8VDxDX8ME1/kKxy
G+aw1RSEZJhj44TMtySkmrlB9o1YRrTXrDPFITO48V+3K8Ex23kjCay5AkT+q4ZW
s20TB03//S0vSbA4j2qbyl9IYQbWVEjtxfGvcLd7vP7Oo9rAAMERcDGULitFYwpq
KO+52u/nOOUQBRb36tibEjo3D5yCr6XxswKpE7ud6sKHGvcjdi7G5WcFFOCr2pNr
W0pobIJVm49HwUqiWmY5TVmCG9RIFIx5c3R1Jsi1sDgXL0KBecI7qCyoOHzmX9rW
VGGpQyrow+2z++0tBS5BDHJ/FmB1ohVpV7uzTOaiVxWcg+A1EBonV+N8OWwcG4WV
J64Egs0fyoA4mDnaIOl9RPmvhJP5n+Bvjq2CbpIRnPQJEYra3YL1/eFk69C1xCzn
Ayx4Em38NclJ8BJOhMTgyBxeaTn+1YED7a8sMQslwRjEt+FD8Z49BK6ii131kLpJ
M9/jzIh7JA9tXUxfMTwA8kNcv3XYMrQWtLdXQPajq+xO3Zev6D0Ze8FBFLjp5PHq
bV1Zlyk2BV5SP3fBHcoEyowsmbEptiZLxAOsfQO9EHpc3xSwtoHYbmJ7uQZ7GkAO
MZm/TGq5UMhZLXMQwWuVzvKdsGFlL5muAN50cPJBs27syAysaqq5U0OK0NkQsbrN
K+sE8SkQJBf65b6p8Vj75v9MqEnqhpsCEJICbJDsSeWPMsBeUTA1s6u9SAcUQM9l
cuv2SUhXCnghUU8AMDoz/1om/P3HmqtJwQh55Jd/r0rUI8TuBO31TtxmC3BITSCg
vAoP6fWFlUg1dpFPlatXfYScKHyXQzT9Xolm7lLy09JVFm+GIAcHWeTguL0ja9D2
MR/Ywezx46nqsVNYRt+ury/eC49/e6yiSKTNKChfPyGDWWPGvEy+CdGzvRa0cq8z
mgsGsPqQbuvxoUHfBaJ7Oi/uiqQgFGIeeQnsoOfUs5nRsFpulZoul1Bp1GmxylDN
TOnB9ziuCXh2NkZAObgS2CevgZxBz4cYIxo5sindVtv3kWlUDZaoal8NxF96S1dW
QkHJE9W6otUvGZmjW7CkaQigq7kbJgWCxRYpJQyFROJlT3Dd1T96mP0TxEspsmYg
/+gFna1dYQz+6F40ApTN5qnP+2MGqUcZ6xCO9B0SKuwNPeXK/BH5BqNII2IxB4nj
FZjWFBEeJs/3QrR777Z4E48pOVDKPW8vwl2CY97OLCiHotsVbxGKdsPt9xZQe26T
FQ/pjLWzftCRdWkPN9H7OsLo/wzB7nt9IMcl4MMXFIVXnVKMK4wCKX2g870gk+TI
84kw/dTkavi+5TiY9QGnOl7jFqA2FRuMIgwysfNfzb4IR5U9hzgigW9QSkhnMChW
GopZPAwzSeYRAWinU0zN0Z0v9rys5X0fKtWBujzcUxh18OayDY1Up0jXFjn8EvI8
QKpX9umJJDYSl4pcEhgQmR6aUPUn8YTJvGx+uulGA5r5h9+mzjAfKALRu2burRjq
UQdVVVWYWvMMMm/+3MRr+Yi7OkHGauM3/10OMcGMYi3FfxpG5/58C9qrf/fPZDqw
cFNqyWPcG5o3HStd56zJgX+w2+kjleZOyGVbgdZsDUMjV7n6sUWgtYLCwSAodQDl
7JCHiMyGgC30liHR5gAllcyuLWxJD4exVLoZRtqehnTxGEFoR0oB5Y55tL/jhGL+
KN+tu+dVRRX53iYzAITH87izbVyNcUedy8YRY2dSGzE6aj+IpPGmwaDfa06D5VCo
L3iOBUZlB+T81CIbhiEmHFyZZKSeDzQ/u10yZ0Ma4Di/6SWwSmQOaHuaOUIMb/t0
r5x7Cq+NVcZH17zjcI5RThuxJqsf/iw+M1ywyf0WGD3tCCeVOxTt9pkBzp+r9///
O5X3FFKQHEEVDMFq9EpiuR6YuQjyynPe+HlUff7Jr0aVg5RqsnT5IpJQ92OIQmLn
yMe4I6om/Hgh4/G773orbdlChaJc8pA7+RV5iAolxlunagSX2Jq6QaoqSkA24sev
UvWR8Jb/XJ5150iqL8rlQ+zUQC2VeeCqjuObSRZvf0aWnQgPS431euclUClypC2c
PzpC13hNakGbmCxApJJNBem/Y5kd50XSg2IX1T7NVSZVVAbELWM67DnD0LN3Q2wG
Eg/icuf0D6zHqwNq12r76052vfZ0IUxxkTOLPEsWqFzxUYxZvRn6mhiGcND8tNgQ
BBzeuwKYHOdTMAwBi/9MOwMnInnNefmIxBOU7FEbheSLgvgTgGgDUQG/BnJ09/JM
myAKCsz37ShTNvf8UnK/55mfA1ekt4UEsVS/tSxaBv4NzVTlcWCCW+L6kmjBpid+
dptGpkOuCkyB/EbkAfVEkmgrYo99vODE32HyoEhe7TX+JtaU/ScuaY+6dj+6asmD
Z8cQogZG5YFLGNhLOf9u1VlCOM6VnOsNNr6l+2kvqzNac1AMNHj6wVL6MIf/x+2X
qJdBSvy+O2QIFCK0rnjyMiledKxF2ySfhlmV0ZA/8NE9tW3fmablbjvEnRpjWgS8
1RZJeBWz/3BbEqzs5xg9h7Nq224gUKg5D98sl/oEWBhnKSSgYuq+vJYNAcKQd5/g
2GgttRnov9+iMpDg0Kkq6co0CLnYfP4nKyy48kzXF1mueN1iOT1tA8Q4b3Ow+kMs
sAgs3gvdwHVPBjpp23EMtjkogyXGkcMuKEUtkBNg+gztmYeLHDhIQzEBn9HVKLE9
Mii5xpgX2vMzC8Z5ADgw3UUlnoGnudGRde4tQVx33pDb0A7oAQbAaRwEeZ3uweRR
Y2yb4AiBbNriddyL/9l011E/QUdjUL5DnSy4bqsF09XD2MStzka9RSj5haSPrbhx
UIllsHmN8fN2yyy8Py6l7FqXNKJ2AqFoJ+nSn9HdDi1tMGBHBNQBD/gyCgawt76d
fLNYwimQ6fHSvv5ARxJ5hVJU4gkABE1ju9rIy51bB62pxzyQZAgbVyisnzx1MXHp
I2LwtaunhWXkjj+iu3I42mtFqXYVUjfGpes115SAHY7VzLqcOChCNyoCQPcInSK+
RsaD6k2Jh2g7FVDy+XL78Ax/z/giEp7832kWYf3YwmzRmTXhJYnwyd+S2qqe/h9J
KzsTVgUcW1JetS2O6JSnYqJ3gGm+c+4nl5/mjnxW0ptF+YnjoSYTbMzUt7NKOq0Y
OvZ5ipFivYvpxF+pxxjdSCiSkYTu/RDKPlyaMSggfiKVPaEmJM3aKkP0fPBhSaV3
K+4Z82AIYrfc7DGaBivi8xS/bktYs+pacu6ssmfh5tk8MaOultf2xWs9IKMoGQQL
/ZUuEP6iLaCYZxPr7T6haRsgozbjK9o84MivzAip7SnyVAfiL+HT+ezA7ISta+7r
pZXCGDwxrjuUFlqdbA7eMHv1VtdwT9uGho7M7vT8JB4IcdQ89gxgfSzGc10b4jHI
xSsX0mP6D09N81il1b8+7fjemNea1VwMW/v7ILu/FwtnroNk/pNLlVCG+XNiersb
L25jpBaoJMyfioQBgwmz+1OQQk3RmZXyJZ0A81o7wP4Xiv07OpXEmg8GEigv3wlt
tgtOrixyeJ/CiET+Fe4fdg7HnCIOiAqMjkLdq5mP910iXeRLU6EyHQzCpm6ypleX
rg+1c6WUB3P5ELdVkb5/Ri2zJxWHQjxpu7ZYY108y5SHT68XMDT7y5XlCOSj+B5k
Ef+BH+5p9wvOxF0wnpe3cGTB8gebtg7/V//KGhtMclLMs6Zn+4+72fzm5V1vHVez
EMDjaro8KY+t5fLtcJTdRIW2rvx36aAgNK6F60SyQjO3mt/Y69EzagdGpeWU4wkm
o3y/s29OmgS6eJ2fiRHAc4/+L9Xxn/gOGMjELJcatSbDGOwAE1lUdnngn9DOox+N
BU9qTmN9qaDPIrzgSvCsaCu/b8ijI0+Zoa6BI/f3qXxdMiRDskpN4QI28O3tdGzg
WrT7+TRlLOou1iyDYqFGaR1RJ/xYW6cBSmgoc8aHUgIu1Xwb42Hv1igKNTTiK4nM
Ob7r992Xu7wLX7DGFBpfnFe7EMfI4daX6RIkfabMUyLIOXYuE9rig7gxfCfp+z24
UPKt7kpfK6VS1tC+xbwfoncBXUfvHYuoDeoz70TXvim25cL/GOAGsXGitOCf7tSJ
bTpm00qLc3/RchIaJAq1oJ/xWfMVIs5C3xf2wxBpcSXVEl+rwjWHIXf1f9aXa5JJ
RPGU9x+eeCHx+3lW4aGTkNDC+H2qBjcR5IBEj3ABHbRWDvEodNGv1wWwR8IJFGoz
8OS0Sysm3A1YvrBfeR0QRwErt2o+ZTa314SR8jEwf9ozwIZv5Gmtv19buU8r/PEb
bx7705YfVf2EmsD3oeRtDCuuIR299dhXXfCcBkEW+3f5yurhHuVXvZuew0fQGVe7
5YnArNcSiSeT9BZoCPjpbIRp4OpDQ4rx9rRCAc+4zaKq/sqYZyMMuH0PyPTL2hxN
ksV4+8n4KpYi29wVPm8WUGO3AYm5k1ObIOD+ijoxFO0EeEQShUeLC5N5zqTQiYkN
Zua5L2e1r+9hZqB/LpImwfWEaFp0VmCbMcKehxVgjPi+x1Ff+1rEIQnDnIUDTlOC
B8tokPKzYyX8Nb3zE8uwP6i9kGWJv7Nhs8OtkaKqplj9WcBgkPWMY16u/Day9/Lx
YjnaYwFJKAVucjR+bwToycBOaHPXIMbsuvtAxowvFFnWtENKRUVbhK2Wr0U9yaPV
MmRH+F8b7QTs+3Zb7iIa/gG/9VPW21fBaN598hR3cYq/ZSWG7kdsuE+svXCtiYmU
TEsvM0gKh7iGqFBGegVfQg5TU+628mVjKRNnIeE3TxYa5FWAX/5mujckPgNotQxY
b3kVf827JsO+wyAZT2LzSRojlUC0fQS5TWyOpgZDxOtbBIec7I60J5g43ZCvoCaW
xO6wbFAdvzKh45nDc1GMspDixoY1FezNRjuUbq8xa9l325Dw6yblBwD8pgquJk6P
UhFMwIJB4k+wGbj6DU0ZBv1TwEdYyi4iIhCmiWLXd23yNcQG6U4CYsy1MHgsrQoZ
i4CKp0oCb2DsCizxqtLJrgHVB7tOG7kpsh5DsJaOo1Hn7pdV/akS/UjEhnCLTEWh
IrhQ4IwuqG6o9g5zkyWhqyuXpPqOaYNv8aMG44kBbSf5GmpcvM2DX8lEIgiAz+xL
2C39fUtDOEKG1SoNFcF2fooMsoJD/A/RizYnfRIpRc+Qo/Ib5Z5507WyMRxBQxDm
yqyqzkkQgJuYdwDc9Fvd4iEfU4d5srrr4L98/OKWjOVAtXv0DBBYZZdaesmPTH8y
OmPNZVUcBMOoDiWRnTUs8Eq0xvg8eTdnpybaUap6a11Onvozb2EOr4mKnqukkwXY
Pj27mAU9piO0qMSUVbf8RKM9mDYw38BwRQCSqaJcJzlHsIODUh4FRylULzOGmZgH
OFWmfpnLvlKi8Ogxts7caopOsrbVV+Mi3uov+jHhslMn7G0o3IF+pRXw09xu7uda
bU6wH9Wpiprvl/Ki1VlnyoGLuBTB/8jJo64+PV+aFtmCM5jztFg+UdPxkvTaw8kj
kowPi57TJTXGsyFvhjmDAaySinXLHcc5gdAqfuKEv6ZcEic4DmDClVo2hXE22458
iGoMajKoo0ZH/MMxzBpIlQQkSHfyEg7g64JOwqNcwccgb5qhhT3+UXH2TW/rwlzB
xxo4AdkyWwN2KbWYjdox3ReGDna1/tjuDQkQA4tej3d2AU1gBYgf1T3Kh7LxBix4
YmDpJrEczvmuMF+V1HjXKGTFNB3aD5VAUM+aeruDiZqxAtJgqHRpTgW/Qs0bdxsB
i1AuOY/+nMxDbxJU5sWxdl85rEsqmBwDwI5Od/o9wpv0+BKojFV3kYHScMPu/Yxa
KIaJGyfSs03+Te+32PQ3jBV9TEoF1DTHVm/kHtD0m3v6exunkPsxKuf9dQtfRb2q
MmeIyCThb6DEBpmET6a/Gt7lt6NEBtlOEyGQd7BnDI5X/85tz2JSA52EqmCdUXdf
m0DnBuQCZy9kHgpPesK42B6KRPVaR/UMbt57FH7VweOx9C0AQxKybDpHyQrh1qaj
3l99RA0ek3Q7Z5+4E6mU7wbCpDhlBY5CSLehE9f9zCAyJtzf6GFWJThXKoUgouoi
9mLAkU+5QAqeqzyKINRR1O2+NTFgJFmjdISLTY0Ni83dntomByAvtaDAqM5xz+AB
GWmTEL3DSSyj9XJaBRPwFT+RPNndftBt+pOLG83NQG+WouJ0xrGdMf7ZHc/8j1H9
EzDy15LsI5z0yYJBmYrs72//T9JciXo48czb9MTQy2alv8Do7htjkmTF1fZaOaRq
lt4Jx36fKzvlmu68gTzZBlW+F4d+dvrdPhNC7RyK/70vEXoLevBP7oa5UJhBAGeK
pDChSLn6TrXzKdp8gpC5jJwusvVQjQ7ci4xYNhCoYzcsx0Ni8k8QDEOECAJY/FnE
j9cZFM2p5c9CnbZKmylbVcfY2/nkIBPyj7+6tiWNTbseClSgupHvQfRfqN2eViJ2
/EqhxY4QNWOaovMEp1kzXuXbKk3gYOUoHvWPaxawHLn+C5r0gfR3dAaDEso4Ooe7
nZ91TfVNRCodd6O5Jh6/QHoQv247nWFASSOJh3/uXo8vLLYzlcUhsz2mGWlwn6wj
t/rDNmjKsFuvZAMUFqzp4ruXndPljWEoR4QSNNJuedx+7IU+6fPE1JehewmLSUY/
gqsPy7+0eIvhVtEuFH1h3xolFmrhy1lHc/fx56b/G7HYPukuj0p6Q+HUhMKmUj9F
Bgq60ySRbcUuVGoUDFlQsLNIALv6scHhqVxCT26wY972bbw4YrzUi56PG9G9XUz6
qyIDD09fBuA7t6bFA5NqDbdRVKLipLE7kgQpW51JRfxzPglG9XXI/uCWRZ+ixKIZ
T+sEZvQXyJVSNm2MX4BVAQhsAFtpIpiJElemdgJr9s8qSeVqYn54acg5XmGY32Ct
Ahz4aAQJQG9QV5w6bNwFNc7pnV1rBlWFS4YJE8PHEP84uN4Pn1x/NsrNcLKVClza
qpdwsGqnPUHeBcJRvrMoPxyIQ2U8uhEtN+7MPxFJ1+nRhT7wEOhpy4N8s2Ix1bMW
Eb8qVHUFrYHcRVzpoejT7Uq8qG1oajjrNWbYJOui85Z4P4oZWjMmZ/PsAAVaZVIP
fA07eNSRrQ98o3LcRoMpxuyurzjOs0SXwBxjurQ7WJ6sD1Rlxesu7UwkfzFDHSEo
cdFe8HIhHmE7HGKziahlZr9EX2DLdLkeqM8JdOiidh/UmY/rExwGhkqGF5538A8L
3PJpE3CRN+e/cGgBnnD4z417SYvce+VfJh2t/S3cqDdmRhT9T4UdG0xS++qe4pTZ
Zzyc3sMqGw70PLBTehVeFbQ31yhG9mv6poEFCCdDxMZA2ZwJ2v8NSMJEv1JariAV
yGX1SJoevh4vzEHlBmbJP9xSrfaeP0AFJ+g/Sv7KW+xH7EI7X7X+MZCOGRAGXL9D
XmvltUMIVBMfD7tbx+ZxMP2JxGBKIcME6ZC7Cxgw89uQ2pvBq0Vn9IiPDb1fBEDW
8V4YNXU+aGY6J0n8O9rc7FodWOXQ5r0s1zt7Bb1dM1V27zsxp6KBet+utRi0ns4P
4zbNUS8SpUfoV5cxKtkhVYGfaI2lqg7V8OYQfjGfoVikgLEbq7dr5X8rt33LdmKM
AclxPYGKpgXXfw7xwWkmtSk1e9zIvkudyMpJlsxLY0KxEzJdojU2pKUE2XnZFFxn
+FV4dwiHC5YuA+0Wb/ttCZbj/FJn4VZ0NKfh9kiXT3jRAwIb7LzSpe/D49T574ni
El/prBx3eXxv3bUbdny1cCmU3K45lgGF5fla3+NYUhSu9H1ClsJkLO1dBWiHVSo2
3mcx4W6ig1K9a40Me3UKYVaIT4v15xarPBhGHwGpNqGHcmNEatolHGplrwWkPoIv
Glxa8NihGjaghxIiAk1WEdB9MGrIWdB6CSEXuP5rw33S8N7UWqyg2wW+UR2/rb9/
ItoI23iamrTFk5uNhcfxkBl/bC9q+0J3iIbpH639EPha4yyd2wDjC8KHbSI7ictw
0pCz9a7wBupvITJd4COXKvLMFuyndV3rXZcfPuPHH6AfI2yRbf32x8U0RQ5uWvQt
cJ7F8UABoqebrq1um4eMY9KvvPsJn8OeXzJhX9cLLqd9onlYfbyhDnP7McfUR1d/
AWthY7IG/O2SqTMwW3huTdW9yeAjIQMiFrCC3ICFddkjEfZQrWqMrxgE4OeO+Up9
JPvL1A/7us/rvSedfAfab4ufJXVW5XfAFP1xx9p7fING6gH/+F6/iI3GYbFuznIo
I2aKJAk0U0W7jbT2pli0SZL1kzJr4oxNz6Wcu+u5uucExUPKdMSY1Ed5J7uQRg0Q
4Wr43Ul/7P1s9NWMKdHurk/ev85VG+JuOsqnCvTM1bS2QeG9oORNP9cTnH+OoTWU
8eA9ax1Q1uezLrtXLk5IeKqJCFHypZmTJj0DfyoILcdgk9UBA/y14H1zg8j14m/U
+i1+efCOrOOOwMr69AiQMmdI50xvRQdZtCbhUPZOU9h/wRYb+OMRlvhOlMTZ4Dke
fo0DAnAGzry4CxjaXKAnh0z6Pg9w5MojPYhtQUAaxlZBqutor3qqh2lsQXnKlk7K
BaVRn8xnkYNu6TqEK/NE/N81p0RvNSAUt6RQMwlpKNIcjJDj15q6gqSOJULmnW5Y
Bo4Fg8yPYaeoolLwRFew7fn7EZXYAKDcTlLu7HVABZYExBUvEU1ay8kTL0zW1Ofm
Zvgb3AJ+rRGcH8TyBwv6mH0SPiboFsnCtidlbNu601ASq6r3Uaa10Z9dnFQ1K3zQ
XSr0ZPncB2JcA6zla4j+MEGB+FdNc+BO7FtsMrMt6bhalw/rbDcVI9VCtni3IcPo
8m4NJYKnS0uzi4nfAueayH8KmgqCOFIicuRUVbKsI+3k/qkJUQx1k0VlmB5DS5OC
1eNO7HR6DtQ4+M2NJtCUgb4npjHkKuJHY5arrCNoj7m6LLkMenV58u0K987rj2Lb
SZvn/Xr2XNoopgQ2dmZFndEmr935NWJW4p5UeCDrTvQm763Sk6Hq5uh7WuNZUYZe
wvcdhRgnfL3eUB6wIO51pzSCRXPQ9QyEENshgYEudailC9+ruUWYOXzoC/dpNn0M
vM6TLkT/ZS7oafgeOHv3r335Igc+jfrCN++/g4XmBOg05yQTYe6fhrEKtd0yYBHo
kB0S8uLb0qHs0Y3Oyg47B36R1nguhS2h4bPJi9Cf4xaBiDq3apEtlZX/d0Yj28bQ
Gi9JyzHZoKFkNayrN9cbrdyLCYTM4hRhdT+vc1fitxZcHiyyoFK5R6ZrHLhaxr/S
YzJ575adlOi+7fPvXXS5QZA3e/WIqCwffYN6DjCvJq1hmFktuqVub7B9Nd5FuoWw
GRSbIDR+FVHAyC3Xph25wTmKu5B2xt6i05eBmjV3NIX1MJSt7dqCBpNMzAcqebEP
xJK1aDtuEzN5Vim1HdFZSSaCvPjVEDGiOZglvZCewvT0GPhmDC10rieQltp83z+5
rH9+Ok69fH3G5IP6r1kH2gejGxHrtr8sOlLlV66sB5+xmHti7k/0Dc3Bf1mGBgx+
0TiUAPgL0F5KvEOm/a3BbBfnDsmwMhrAwQ/Ofq/W67HMGWKNheO3voNhpuZtZ0Er
spYM4PxPeha6yPEBe9vYGZzQQDNXci49Qe1QFWbhzI/zFkNgundMEgAlYlYVi9oo
+EQgzqr0JLYK71tSYxy+96BRg35mTgwH2tZjGnBrLOg/wZPLdKwNc8N+6MeJ3ozg
kIyyFGxY7SIT4YkhxKCy42VFAIJlTiWzgrfWOgkT85HmX5vEFWRfj74Dm08sCvd+
iw93XykFkcKKElxZ9KEgxRbN/k7zlUyhZq0K5tEcwUAfxJAF1Fnd5ewIG+7Nd26e
dpQgUwa2GiEPV3E+l+Rqnx9xBA4ZjElHZtDJPo+sVUbiKLIiZBmeueAVqtixeFyT
6v8Y2IKaKHLxh4eG0T9NTIz3vHIK8X6FiS08QeXCY++wBfEnm0lQ0gKWVep+MJFQ
zJZwmGN/THzkUekP7WxOflE4vDtoIp5WftOHHmdqjF/YK2ZaApcuH1SW+9DE5ARE
YyUNp/hcTb7teukBLuBtOq8MgIW8OK/ktk5E9lYbCFEWlpdyYtRisz+/QeN5Bm0C
PTAQBZQ7bZ4ubDyklvoyrMhmDGjVx0Y3qttAK4aVYICCA2EbQGjEZsLDbEzVV25a
yBXDQVLochwrM4xk+hLH4YXiM/7q4v/RAAp9kkjYQpFNRMTmd3IjJPuww+FdsieU
3ahJzE1hC4cXHcflfJeW7nKJGkBqtj+H9lo/1HnDYZ3FZiQaf9dWTWVQItNoQF4E
XYe/u4ZCrwL6junKmMv3HFJTlocSGcy4O4o3oH8PfXG89kkDYtK6SHpH3qMXdooE
F7ukBgEH/3gTWzEYNuyJnfigZnR7Ys3qkKhH7djhBOSTIeJp8YMhJtdUjS1V+M0j
hYSrXrbuG2lIF/qcJy0KKThIzkDvDNYHOHCcuiOuMm+9UoF8duSzOtWpnbuYnobr
KYes4idW1TYa34WAlbIb7sVDFV3J+SRJRuvCj3yBDQai2pjPqwKd/UACwCTGNi54
pj/mDo+pLWUXB/qGAsEwUmQKQcbFoQfCkS9g0VOabeQ8IW+m7pKu/fObp8SW7EnF
jgrtFr/MgUAZ5xo0ULC7G2x8osObn5XruRDNXNcmN6aadaaaqru8v2A+dV8abTUi
xrJzPZAfDMnlUuHtpSdE2eavF8WfJ4Xv55i73FAv41Pxw3ydsh9gmBYiCne9hxd9
KCQAqcVwx8oSOqryYm4py/WPME6Ztm9IqluzuABkrx4VhvtrkiE9iNfdM9VfAOo0
hL4mFjoBuXSrWMRnqsEjJ00bVYq6rhlpFF8bi6px958WaNQ5rRhAVNCAzkggJep3
2yMQLhHwbW8FN+NafwdrcLFLJReTh36tLyUgTl1g/wIfM4TOwwYmdpablUfEiuTz
pJQ2SdRNO3UuPa7xnLCnb6HmZg1dVxgYE8kKIuJ/VizODEkDlbhLBn5oFU6xvAJp
xsGMEIZ+zqten043Df5lZ2WhtH5K4b37k8aBjM1IcdiPrR2n9yHJEaJ8P73XhOWV
BcqhpXHsidovOIrX1hRYM0UI2TfKVtw/i2IFy1BdAC5YKBlWdBXqYyGnw2VFjcFo
WklIqFYPBs4YQ0ctepijseFsIxRfLoTa9kYiGsh+IJERe4O0F0kcTwuEwj0F6feq
2g9GOeyJ2k2Lq+stLlxtz9vMmqCwyrOl+R3TGk1G3JcdafJj+nF2HryjgoGlIFCW
1L5gF1ITe5D0AAXZhUrklisdOd4+KzxIrPMC2ODIta8/kzUhDoOhEZ9hXmnWh2y4
FlvzhjVULyRv+IV0p6/73XBvbsrLNb3aGZ4mryT75BmMQvAVpnUSKpFfhoqroMyU
2N7jTKt4/yYEiLR30fkIR3CR1LZenseTcbdOoLzt9Yjxwh8E6qR3BXMYxFuAcFiY
G7XIC4PDOv42vMAZywvFY3/orMM2oIsPtUrL9ed/zmx6D4Z52fkCvqBqnEvCj0Dd
hlNn83sjG0XD1xwGGBnNf9NpGzyUUZapiN2c47MJIMitMPLjm1t4SZPDdmWnhs3f
04WyUAs7bWOusi6R0insatUxK/FVLD/VlhVkRa0QmP7DB0MZlFacuPtShgoFppfF
k17W/cjeQ8VI/U/vXpbu+BDAp3rgoqdzPZk10ycrZ5eMi5tJnJ84IHvtfT3wkCD0
WEn6APdnz7ppKiYHx0ddw3wDpyCJdvcHBkBPazfCngwqFZV1doDhuW6MsmICochN
MPqKi0gNgMf+8k5BNQhCnFfKauqhrSifthuOMuaEYbdj/OYI4iDcTcwRlzMdyOx5
dDnzgYsfrjJ1uw8bLwHwz7y5vvyzRaprcwiysE90R65yymyXB6kcZvYgNZxLf5gn
/Or+/gyOX3wI9elW5NINF6J6wY6fdFVZ4kYsg3yB+I90tUHN8opZMSBhXUppy4v5
0SbXnq6+2FjLDhxG9DoZ8P3NdSoYuGk4BHD1ycCAD3Zx7PBnxT4WZDUBqGQuF8xf
UCZVAQMpBP2K6FODwstecqSZADgWsKqJH59AtBmMux8Z5Oux8JA960SVbnHK5j/z
eEFOvKujy1UIksT/FJ2N9crXibOaoQPUkdK0aLPDj+tT6xs82gJNoYv3bkDrRMWT
x9SwyKYzJcpvphjWD00PyXAfieNA0XBnrl0Hf7Suqod4/dKZjbQ0KGG0dl4DiV7h
AcReVRtMdsMUwJ3FrpUB5qbvEjZ98wtg6r83/rWAtu+XxoT3bcDnEpWCiNs8GpNu
KUhYm5asLdIaHp6mFrH1qyzWB2HhgcJFaJeNv9UC0zcJ3yPmtljMz/H2VmFOtAw7
jI9Hb4I6Ej5H+UKO9D+A+1I3+A1+L1OGGnzhHVjlRIceSejYe0wqrIk2d45nlvh5
3LMD7Io+4awKalUPErAV+YlpqFxJ5IoQX3BgiP5Li6166fCghu58778kcSY0zA+i
h/a+MA+sGd31bEulaXbDmqvP+4nlY6BKsu8XWKfe6AvRW2TRsvCopqrZJqcfyXWW
8doT/Y0lNoYekiiCNKkfQ1I+BTih3skSw/f5Fr+zWpsgvdwphkberZFfqqvg5nNU
SSn99IigH0VZlV0epDbDQGyA7a47RP0a1qUKvwkhRA7554zQqE/sIuDaXsUKMLOJ
rXNKOSlUi0NvXG9Ll9J0OHSoZIZXlJBwlcnIrSkr+vCYtj3etM6arBzZxlxOqnKf
TJbzaWSIB5FEcxKl/pCGjwNKEPm5Sdy7sy2ffNpoAm7K9H7OqusTMuIAttsf/1mK
S/mMcWthDjc6K8jyw4xirLEupZkzbIh4f0y3M8FUpnRd3ZOvxHJTWKdAPq6GV+y1
z41OkIuouLlR6jPbBWX1t2e33Rb4B8xkh9UY/9zE3z/YW7dpuVOgLpaemqj9Qcqk
kZIuP/O8/2uF6WVFer0VObt9wfTkvYIeGg2VeP+e9kqQHeWtwAsCzA1oGUzvCvGz
/2WQC8NcyGCjiWFY6nPCWWAcPc6swCr39le/eVRPtYIkz6wJXppTWH6IGWXo3Z+t
AjbomAT78zwBj5go4mtMB+/A2OgwiwK5dCPaVjlBMfQLgjdBiW0lvUMQUgx71YDZ
zhRt3PA2NLyu1IxajNJzkdmFR6p7z73XkFg+8Xqw/3cyGTfCXVnXD+BsiSM0RDFx
A/e5kGo/lBAQwrsCqkLPwj1P3oGc8tb0HZmoq4tZv5GUXEN/ioxpoOP/NxGjY6A6
FoJGVHAzcR5z6b4HX6JbPnrqoH/QXNkrBf048g74PuqMWIVO6/owXmGwS7UX6zZv
B5bMaQC17/Epm2RErmVRPbidSD2tqa1AsUi90hDNrDX1OPaFd7799CRVJb/6oy7Q
NoGUtI4bpXFD94xkCuaqIaRDOryah0tp3NmVBbsxpIpPCo/KyXNkfMmTMsCGD3Qx
f654GMbsVCuNTWAU9ncrA2kw9mGgwlcGqC2LSa2/ly7B4lt9tHznPDsKErgAz3yr
Bk9m8D1oEgUnO5yQOnz7zgzoqglqTrCjxXXpXRLeURTO+arudHKGOwQ+AL8jWxJJ
IvL2TZj9E2Yr5QFpj3m204EQDIk1NAH7XbXNAYJH6wkcbBYH0njOxJZ2zxiZU9VH
4P+8huIcenwlvoVVPWTdnmyqcOcSFMTG7G5kxaBSGnOuprssaMF0LyqcBuDdTWdc
mHllvByuhqos/Y2+yY7mnUUZ7XZ6Hw91kVRHWc3qGMOkBIkVVIHFL071Ua7GSfJW
smegEH9pfDN68zTgWtsvoFfjSC0Bi6byxq12XlJqr0k5Z5F1rVmF0Fg3LoP3Ghaw
aVtMyuneD0AV5t45q0z00rXnz0v3SBQCOy9yrdFWW+ZQmqm+20YS4Xklk16UKABL
xji7w8eE+IYQXiyaflUw3Sc+BhMypNKuLGIMq/dMf38LFCaRS0rN4GZQK/VBB1ZT
vBOkauz4N6xZjVdwFV61qR2N4yxDOAKkj7Ero9q0ulwHkisHZeBM25890YPCwZYs
lUnsBfo+NK80FHTRv8KxlmUJCRvVQEPxufg+0oleqB6OFAG4qoJL88SbOz3i1pQ8
AnTIam8ynWU9RKzysIs9qY16dmAfi4Z3Roez5FuDMiu1g3+uzcP1dO2aZCS6o3mP
irNjP9VldhopQU68FFMT90wxCJIwP3jtDGZQpuKxjM1nuV7pSIBE+/5c7r7AcoC5
HPdxhzpS/6svUwULUGzbre78Jy0D4fcdoMB6XWzlmnQFRJeWZuNT4+JKvHk+eUHl
IqrOWFObt8ROCSYW+7s7CcPi8piDyBy/nzNrVXGBXoUpfQO5hKl7CuMnoOdrIQFU
yDxv2JNfXfgaMfRE7kiPXbB9YJLXRrw9/uc9N8NaiuGD8fyQtKoT+ZCU9vpigC6S
vJZ9htI9HDhccbPmZ0pGeJv+pQVa7TXKNrl/K+L0CTde4whfcjMxX28mbUnLxb2f
LRXQR+zLK0gwKKLU+Qx3+YaXTXa6yHWT6+RNmhI6aNhydY38Yd0i22i1Osm5ewLG
B+zp6jQsGQZhxY/CBE/HjyYWaw5yF+1nA5bPT1MmBJXU5kW0U0c0vu28seO9CwgM
6M1HK20V4qWiB+mbN3kAtu7p3TnVxQ6d5IEpXFtJXx5F660YHVdS+XJ66TmeQqdh
3ePZp6BWz9tg8TrTKqmAgkDspL5tFRhLSk24ASTfxwZ/l/LtDP7NkLDpJ6PFqgeH
XGfB0GriIk25X0dAV97klV3fLXdzCJgTG/12VsoeELW73OBrBFJwc3dX5i/LpUUO
LOdoCeGsBtjJVKylXA2UnC27L9CumCf8n6JjmGLA37/v7fmst4EtGYQM6BdvxROX
b7ekDndQzTfj7zamZ9A48dsIm/kufdmcY8a2EXmXURHhmtXeolA2HPtiDfNbcP5M
JmidgeL0hle5BgBahvxClBVYSfeMdNngyuz+JWZ3JXVKxAC6qTiKb3A0jYBKTcCB
ANyLF3RyDHiOYO4adIpIaVO4q866CO3DMmNM22+HZzCTL2bzjGcUImY6iVFnS4Tw
DkHTXKfF638/RpsQpK7RyufE3g3Ju/3Tw/V9elXlZUcml4EO0/QG//cs4c0zF42+
0FDlq6w4BNfLjsrIIsRgZqNJvML0Q8109b3iKxGOioqDZ9zbm+9QXACO1QOG/FZa
WQ1SFHcUypyIsVrHFZTotdPEcoIRa+W+5GMEy5jRpbE9bsR+3dio95TK/Q6a4iIf
kRfz1mLbq7U9D9nvgUVbrpgzTfpwu4x+gShkxDOP2auboOiI8oH9sIgOcru4ABj/
CXWo+ldCI68dprf+cS8G2mzQtXPviJkd4i/esQkQqIhKO2XpBZ/Rx3QD0neOQSKW
SNFJXglzOeVSmwbNYwhCj40KeI65ynIDn0uelG3tJd58UwxcRusGsVYKJaYeLEMC
fk0tiGRPIIkODpcPs/dp7+0pIYgrdn5oJ6EuOmnLaT8x/94jYhAiUorowtDhjsnk
JXyBkxO1rLw3xsANOCXNtmUMjpkbDY5IthxNWn8pAGJUe8PInji6b4Dq5OAEsaSQ
gQsEmjlc2fwKj5Wlux+hRIxNLJHDvq5S2cyAHUAeX/oPAI8kUivvRD5XxHOnpNy0
MjlAMH2fU388QfIBKqK5TEO6uV5oknIWyItlFQohRsmfiwLZ2iV00JJLIdODpix9
T6W7amufoBRcxbkH1r48a0kn1L3kC6i9+kP7TBvVk80PSFhjKDrjlnDLX4IHq1z9
CitDQpVAJz1bU8A1L0DIFtVoy/neo3FWvpLl+ixrlmpeyfMPXA+KU+VagXQd8Pvw
gnySzmYYZZNHE9MZqD4iKxBdYLYfI5zpcqEHeNP00Cq6gzDxO/tM62OYkHxBgl+Z
EH/6so6ju4ALRlsLAenidb/NE2aJRfQABdUKU3kATMlCLiYTXfR7qfW68BOnvg9S
YeH6yJwRUTMRQSF0QhZ2Fcu7uatmbJnGPQi4QDYAWVkfZQpDE2g8krZrNUVMhIPj
3yeX/K4QH7+d4/zD9UfuzgIXJ8kJuk766W/DjjpircQkgWGzlEm27jcu2GZFsnLL
TzBn34dV3O6e9//D+2WOoifqyFCZgJGsTzwIBDYIkAfIgRnL2leZDNtMawrj9c4e
IxRw8cnwzlELrkAkjp6pjHIZNNNY2yYpPFuoWYLKwPVe/2VCghabwN8JPK/UeUnw
mgx7cdM2+4Mh1OYixSGLrinfoBbgbNjuEgFsOJuO551Sh7a/n+G7sSYvB3pFD6fA
DyPVzPlcvaxPi4H5EMcr0VN8/V6XR0IGAbyC0jKif9ycMi1noT1bCKbfUkjUI0zn
OOBmI1uX/d7Rll7SeJ+vvlYfMaY+1G+jRdMqUO6uIU++hhpKCqlVFekAVT8mqwlD
XoGv6jSdF70LaBRbEfcY8VLuJwQYumzbSWFPFKR5yggsdUgESU8a3yQg7NP3XVhp
Ll9ksoLIED+pmOvpe44DA4HBQ0yjgGDPkmP6/OBoH/cQ8gBSeY7SiwahooBGlK3g
c7iQK14tuLdw+NoLhPjzYpjBCx4UpSzadCDA2VArATGcGjnadSHaD36X+lSERNqr
rIaFkTiJcj2/M/i5PwOMgo5i3gtyiiPEp4944gV6SzT3L5XWuFb83SZatF8XmBj+
/EEkEJaRlIea8qkiMTB9uD0/lw5H0o47iFEkJStHufQ+0kqbHGTEwyrzla3oAOY2
+payUDMa3xgdjQT7QTbNrEqeVCKzMv7gEHDLr0mwSgi6FMmvA2JUHzWi3Iyf5zgU
M40Bkpugd7shS8iSLpGibRtthEhQtytF+UyPr5SFhKzErd9Hy+MV0mPQHcttQZnn
JIFWcZe+9UQOWqoPaKVIJwkBEV3y9uxmSxFO3puazl/SnsNkl389yq9ka8e8rFvZ
50uzjxsueI56GewKlJNCMdYWqFNhNi9CpeE37aQqgYnkGL7kxpF+hsKFfU2xg0mU
3/kwZZd3Sb1NQVMHfX7naeZjQa7dewOUjwpaaQxZpdyMf18YubWkMu23E6616uQ5
ET5f9YYs5kVfupI+MMVraY69GDg3GUAV/VfK14ru4wjq7bhzk7JNcRHF0ZD/USai
p5WydNBu7zDK0rQh+SfUEiLOeJw6hye8e3dFx09XdMQYsaPd7qTXaDOVW7pDohlN
zTFGz37geZapI774egIY2Ac57geHk8kHD6LMbGZpFNKDooet/PJXBb1Vr6nUHciO
3EvJSsPhHzS0sEheqGGe2OvJvUnZNoZouRJ+x09HQe0wFQOHH9kUZ6cFbx1KWySj
QCDE6/kfxEGievQ2if5sm2XkTQjA5ZZ9i8q3LWW2JIZXTSwyAZIXHOhc3qQ1Lb/o
XKwf+S7UOdzMNgwGmJ0rfqnj54QFpRMwxJGhF2wRK35ZnMkuhAkgLXj6lP0cnu4M
YSqj+RMGBCpCvQO3k/ehlTTn/dCNxenTbXYKScFmxRve9F9+QAo3o0u3edFYp0iC
xX533BlETH9FwbVSkFMsOvHQMS7vVScTls+mS04o3OIGRYdWGLtM/Va/3QRJBxhu
X08CEL2I31ndmpkI/HTrEBi1PCkAQ2XK5uwvup6z5L1aDclaBNRIPIaq0esOotnk
j3GFCJfv+Bq7qJSVda9CcYubBv7018eCW4AYyx383x0d8/LNXAGSo1qnOkU/91os
q784hJmaYCUTwmMDeROdGmgvKXB7Vmu1abvkguGRFGYVr4AbvIzKNjXxRIafsYHq
mstex6wALHFpN0wI3Wo9IO3os+Z8kR+ulEbSds7WePI4IxcYwsbQ7QcGQuIbyyjJ
aShSitijKwKF/Oz5dePSFiUbNS0uEaCUmxI2z8ap66gIbROCeKJ5o9913p8tBiKW
qTG2WtL/w1vANYGnzmc81vMh03OBhdrVL21/S2nuckqlKGVJdkp9DWbVaUNwCgPm
yDsZ6kn+cCnDoYc6nwUJ8Y7+4UgmOKaBZHMIRPoyTWXqlFtkgnlzh8hCvCibDhK1
gby3SBgI9k666CvQ7PBmA8u+lCza1mtdh37BPJkOgIyJSd6dwf2IqgarxqeG8Er3
iEyDAhIMsJYxckJume5YIYWpc2GD1VUqdTeOKhAEraYz4a00nMM9k0PJp6Oht8zl
mP5dZshdTmQedGJwpFtgvgQxQ9/WPN3P7B9fu2fKDEWTmEMyjdQJU5iNSpDE9U0C
+88XNB/lwy076rsME9EormNk35H6GF66vN31rALQ776wzyxl3AxwG3Qgtjpo0yFS
0Ciy5NcgNPRzeKy+VUPqXtEahRd5aTCc05FM4U97g1j68Ah4dN0RUL/wPA5ctk5+
V7+YacFS/BSi9obJkjvZ4F6gCztATskr1wJiSwNfa4ZE98to7FYqwicsLZYx8yuu
iruSq+nvrQ3gioCsbrp+R0IP4LYVqeGVgA/CYNcVHsMoNfU+hklc5wT41xchK85K
paifnsX84MatkXj/AUvcHv+yIlMCTtnhborIvmG//OBbwQ1L9oMqQv5hpLhYEdTx
6qWMitL0K84yjnTJhSQ4gQjXiHDLZDQ4CxiqJkvX7D2RVroBb8zlJuE/E2FJsDn2
geITrkbnkWmm8DUUyk6CA546K0fLZda31rO7EDWD5I3e0xICSV9pzl2VuYJWTOFT
pHWYFYqzPTNNvVgr+bMUvXm2eo3njCmkItOqDp+rok21NxmhdSRD4Am8J28X0Pu2
fi4Ww+qYHk677DsR9YwxLjmJ7HNWm/bp2PoCTympHQy/nC4DaaaoLyWS6BOAHJfS
oNmHHcXx3QZaRIWF7+cFTVFubmRvAgE7E7MNIIAO7tQB4bdeak+6+1R0Stb3oZuX
2hJLg0FckJeZFW82llP+8ofxnz1BT6cp9wnGErTmD9M7nHRfLgZ9SpqlCCcz3fJv
VyOCit4U8FSGJQAcIx2xVUBUNlbkC7+5X6U3k3zIvccLwfyZNZvKEyxmR4cgUhoS
ZVw5dyAi0EtnyROjChHh0ClaExW4gvgLf1iLXbBcEpk8krcG88ElFY+mt6GTZsAi
YnfqotBANPGz8aSSClPeChm1A6S43Hh2NwQT8rAnyS/uCp8v3jgXCV2cVNyr/pLp
gfiXi2OqewZtiKVOSszZ/osZKPGLOuo7o6H7lzSHofyXLN60StQc3+NCllAnnRrj
3IbQ8zV135WXGl05uue8E6oG2V4rb+Oc7yb5GESGp3OtwlbzJoWpzIWuA31SHc2t
GvAfR+HAgotv3CTm3JFzwFPqermKiOXgJlSGqboVX/s3MnWJViVxHL0DTcGOBZdN
Hgy9jLxVUDPucyDAeltA2ldeyo/kzS5VUG+oYp9FkHMqurSB3f9+w1v1OcAQZiY+
CNiI7MIMmUjBtNQQdGJh1fEKnPml6vo+TkOuRfO0+lQpumawC/UAHpbjn9kdcURv
5iQxYPxkWH1bRG1/0CcXJulNc+o1AMnyQ28rAr/VjRAFd5KjdIg6mUv3AV7drf/L
y+ul8ZzsY91TYFcRkJcusyJllFWJVLVg7SVzmNqCIghxLqcG7P8vD625rUL8iffE
JdhINiL9zMv0BGxk35zRNqqoIQPxVvlXsfWDzrJdr8r61NvrTH1xYVvAOpTz2BXh
ZYn7XapyzLuD3aIAk+7chU1vT4JTxFw0V/WrTWoO7CnH5TincomYXUqixrJWfaVp
jngyOGdADUMYkC6lTZU6QQw29gFgM0tv+fyAL69Y5j8FiOn1l4G/Tb/b5yixK9Qh
Wh30lW6P/GsgafaCKlxvROtbP2V/4TY2dMDkPik3S+HS2f3PjhukmBgwz/JIp4zp
aq64v6eZMvGhr8iDrJU0O1BuFC1kuFdrFkCtJkeuS+HAXRhadzxakbH2/zgj/u2P
bBWycGndMoKvbJ3776dFgHZ2vTDheV9BH6s4G1fZBeqccEXE4TbdS+15s9YaI76e
HEa8BeiY6WZtlt1T24qvRLluM0sjB47UXFNGyaLRsmuIBQvijE+/HMydgk6Z8l4l
NS2S6eGjTP0BMDt54XPigHhxCkp4lJNzxqK3ctY71UK8CoCaHAPR4Y9GyraZ2yaI
4UR+y9RTmk7fjEKRRD+b1s2vgtd+ovVEYTABkpxWdeueB114+2agjxoZukZZPcdK
bKSTExuepIMu+m/H/6EgJ+Pg/M4EorFv/8SJzToq/zvaDyU7455WxiJrj8wDfnCL
F0gHx6R4EzuqznPdZkAhhtwCt+yoqH4oJA/otmu66kLL4Cv9Fzv8Chxmkbbe24VM
FGyHMMth0FH2tUc8vRJ04WhISvPYl9XNEgzKCVFI9oj1fqFQjnNvemqUdSA0mzKN
J2aFSA6ezl5DuF7Axn8JpKrkIZwBI3VaL5y9lIZrlOr9Eya/8nng85QA/3Pb23Qx
DsEYX7Zga/tEq31pGX6HUsgYR47CZxtYbD8rQPPrdQJ9ZjhMQIEIT5drqgowZ3ft
Y6TRFJkHqDi7SmH/Wc8HYYj4BCqHBgiWvvTuh84pdQ3WB5UaxqRw4Xrf6+jYfYrP
uqCNd5gtdAwXaPP70v99iOq7Rw2geYJdrUehfMhubF0jCL57RbwDEM3GGS7hiHcE
EUMVuU2P2YhXE3CCxcshQN7HoUAESRlJe9M/39rVlobSeXquwl1kQutUSYUXMnea
l0PcQr5oUFvPNEl6EcshZlsa8gNEYLC1U5CW2q91jTuzTy0jxkYo8NcomrM+Qej0
wqi1A9lfKi9bnikrZghUxxLB277c3Y+CxiuUqpu9QhdDxj+XYqFlRhhz5kIRIBud
RPBdZABwBajF8lx2/6r/BuSkYb+setIU4vdd8O6OFbKagkkPrfdaA8VKXlKTM8EF
qh3YNpn6DX7rc2uGbc/Hj1Cwjsiwr+GXYBNvyNPQmLEZ+6E6QE7ZVCE5/8LEGjXE
iUHAAvp1y7vWgfqf6gNOqMnf33rzitzvSGHlGLrhWDtiNwmqy7CwA5WOzPMyTQIA
EmMnwOIpwCoyTmY8dGZAXtC/ahXQWgmNtcVcNC8DJYzQd1Awh9/TvzAmoB8n5hcW
6jqhbB4/RrcX7FY7OhMUIj3STJ2tED43RqkrXzwFIRthZp5zBZ0QC4qtcONVh/wc
JECgSo7gl3lj4SYV1VLD+4nAcAA20MnL6x+BYCrllXBqB9pnpMVAF8jy5AnlOKYd
atmHKJFMEe6DQqVUUq5pMI3BBxUsuHyHXzVuZbBNJF0TiwE/y67MNFEAQxcvXoIx
9lPzHYYnS8ILCO2tMtrSFSiDC4XhKWeWh5ariTD4k2rK2Zz/WP9gSrf7ikis/XfP
nmMTJQ1vq3w623cYL/r935v3N7jrLr68yW8i/Kcdfk+xm/eodKILLI8yD0ITAUGH
+cp+3wFFZM4pC9qMpri1Uks+Z2ga3uJ5lxFGDki+6L6V4feqmd82meAG9t9bm1lE
equri3zs9uBCGQdUkcP1isazghMweRfMuW0trMLlMRAiyhBnFxEsVTSN39yAzAK4
wL5tRQY4+BUBp6OsbSGGRnTvN0rDoNJpykbqg34Z9ibrzG9Mh3bGthoG/KStjgGR
0F2+b6oSNshcMWO8pXetKIvMA9SQmobRhBsSn9MsJROOVPGygE8gOZS+WkAOJZ6M
gwXaGadP48yy5fweUpxOOsUQLg38+K6fclFAfHAfny5A3VYgIV3xffjXp32n9BWT
0vOns4NXfkcbtSDuYgmiQLZ5fTjOZl7m0+a4D53kbsBy4jS+Sa6eR4hx6+9a0v+b
wR5HdR3/4XSuBst2AWRZtbcCdQ/zcDiGKrNIuh/cdeorK8TB0A3v3j0xYuttoU23
C02C02JkZ4qTxXnWmqYCTqT3dUurUMhV3VW0jYPN27VAtdCU5LFvCs39KbPqej3C
XqTS8UNv++Rh+KvEdhw5mQHDT8c8fGv8mUTMxn/ijcs1LdpNcVE4o4aOM1MmdtVS
SuRRq52e/5sON/RHGRLBsxtJ99QGx5UWw6RwS7lhbpVW9eO235peONlvSX/tjILL
HbkwRN2mpfhNC2GCql8MQFtbTOlgYQmy+XsS9s7+suQ87r9Ll3XKLL+RwQLWuJ6r
IqIQu5bL4Gk9PBdA4b7I3lL3AabEJeNfEgCEL0OggL4wsOTlfeuEzjhAWvzTH2AQ
Mux5oOs05W/Hl4G76mq1pW1qAQLP3+3BAEW4BO+s82lGgaty8YzRXHKxXa0zFM+U
e6Sl6xj8nluP3ccfb+hSYRP9SoKIXt5YHW1QJf1Lw4aURGXbCptzuiU7Vyb0Gylw
qS4bTPSV8DMLvPjMvP57RUEnUx4TpLifAvdW/j2hXtYcFnH6Uk713C2QDVDQD28d
`protect END_PROTECTED
