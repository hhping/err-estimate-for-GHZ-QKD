`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vPS2ZmfwW/dCIra5BgVdWjSWxfexhH2+W1ADoi49c+9YDPG2SX9btxDpWmzPhA2
zkc6jCMupekHlD+1ACLiWl8I7e7Hq81xvH7YIPvl8QPk/Sagz2sdWihRLX8R/ril
YzC5QpdCoRkyRjGdbSgFOIrLO8ujuIGzlunYM/ROjUuir/OkkV9suMygbHs2lasi
kb23vaEnSUMOFaZN632JzYaOVQWLz5aBp8+nezeFNVaRCc5W7+Ca3Z9OEh5/VUR2
d8pZ1xl4JE0rcIYHddFdwsP4OsjtsizGAe8Z3uNjaZK/n612e+vQoNoIorrO+nfu
k3MFTWeShHdMGbXcb+2T+USTIZv2kdkWC4WjdcYUJxSQGzqvFqfeu2dJXXP+nsMj
TkuCdTA8/XTWZj9xfkR9I5T43kGvS3U98cY2m7FComLe/VcPKD69QnqI9gESzNkJ
qJiYfqrQEY6tYtXLbMnjLaYArAX9Yi7rIa0uJrPU1gZxJIyD0NUIkzRlY5GFoGnG
S9l2ltOgrn3UNcBs61uZp10Fhtb/DLMjTK5CeecmOKC0JdJZMXT8dRL+nC1WZDyz
VOdUIK7OlCKjv9e5tHlxInp9rGCRj3nUffX8HNQdR15yf9FGawyNCTbDkewhGB7U
nsX5yHSn+uZx8G9EvzbzCeCrHMtGASjgk909xO8BmFqx4kcwBQj8atZ+sFna+xnj
ekCU/kwBtj411339f+3o3GtXQGfICkeSzFpuSRL95jBgih4JnPXOwhiEyHDRZzCF
lmNM17JB0UiZVrERDseQ+xUreP4y5Bnm6wq0YXF8t/70iFbA1CKAOAczic0Dxae+
BvL63IKD596TevsER/Gp1JWU0TRu7q3HXBnzqWEv2S8hX+RM56/8TPQD3tTwYg7F
GWqgpi5iJBpKe2YGiR4yz4/NW6MKIC8DJaKv5RhbCd9R4HEmYe1mJ3ZPB58+aehu
OPapeTA+v/zqwPTZbhOVtaqNZrxocWnsMhOYpJ9j4fz7G9Oz02LYmjXM7y6zPAU1
RNUAHlMThSWU3Dbl51G01QULfPC5mjWev5LZ4/eEHNl5LKkNTz+5Utnxq6CnY7K3
piggUHfut8qaLIHlnHCpegKictoyIyVW4VCZqID2a/83jQhTmMyXWlSitZhIN3NZ
KBlR5yf2s4ff68fTA3qby/jrVn4QwHGP+JrG16FR8iEDGFy1pZAlt/k6yvHa+G9F
zeLNr3yAC04GdtoubiqzKo5S8oIDgK0DN2FLTxJLE7Fav1wUuFmK34QgbjjZwBD4
U5aXuYnwWe5MF4pqg+lkIbiSqg4GJ7aXK7rkqMz1cqcRKpKQ2+VacLFJX4yC/W80
d4e/M3t0JM4iSNxmqA4vRxWl7sWAEQ6xoqMx9+IjN61n1YLdhyE+vBNfCkhLHUhN
q5s+D5He3uNsimVv8kOcgvGEzwotFSMt/W5eOlgWcOcduQzwAFAtvHP143kZOY1b
QauINH+EtciNPSEEPpZnGSDLq5omksyQGoaLDcVadWnjPAoUfjalxSuvgUk5ltr9
iS28PppB2DbAZ9d9B8i/w6elEybM9JitacwBh8XNubETFyeevjiHGkdw92MFVc/7
sxeB/DSXeWrkI3dTCudrN1q6J+D0Ab6S9p6mfi/rM4pxit32852n3+d2xcozHhxJ
PWCXWEPQSelaAgO0wkhttPNaWywzym6pusnPd0Q0CV9zdv8c1smRY9xVyEXgIV9N
njt1rgGWCkmy3QHNHZZf9HvMFVFfI9VanxYBKlF55jgEuS5J6PiVXhVQIpPABC9/
paDJ74QONwOOb63x5HNzcKJGa8TcarA57FDuoBl+XcJVQ8IPGTsR+G0T/Zcpc6rU
XFeHwARK5CFhFQrEi4vyYu5X3fcnGwoR1yZjMftgxGxMp5XSfn7xdFhm5w5yeSS/
d8gDzJiISnmcyRpZomQkEtrIOiwr947qKYGY0WHiHfh21j6LQg67a+lQSbPFi7D8
`protect END_PROTECTED
