`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rmfHQ8vAq7oxPGxlIsbXFM8DE6Nmx8C49vDioaUFPUuFyF8/fZiDUsmUM6GnqGj
EpGcCzDRqysoL0KuD+k4Ki/eTv6dDF0Os+jQbEh2dPhXurPbucrs43Z/qUVWTvPR
CO/OaDga3CSwQEtPO/KY5k1U+KD9AMc3BYMNhf37qLPtoF8yJoHGp3DIGB/ri95o
KbzpX5qTHHFGJq1LLtjyratH67JMtAgloRXXiXNnbKZG9Bhf2gd+HkOMXJ4IR6I2
3rRf+skTILK4sRGT8VWD9jRUF7HH3nTXnrIatpIUcf0RWcgH/CJJPXcnEeL08Nbd
kX6DDiyMfvRVGOUu4IzRQF7dJ6s/bzws43VQYkpWq96ZIXzDaiSHQuBO0WjobxFH
NYYd3uHBDjYOoNAJseuYCmnqKyCe/J5JYJFERmhsRRa/JVWA8pPFv7Ffl9AGrKNB
jdee9Ws0h67fc+vNpL+wOIf8DQLNmKwlF6zVIxATWR58eOi+YGmk5wFfP75y+oQs
MyHbk32pb2PHNVh2lQ3F2tIrOGVR/Hs87hWh4RuS3GovgQwoF9giGUYIFQ+9nI6L
j9F40tjZIPh+e8HXK5Jp3jShus49c8YtQyR6vggWeC1u3O7pPUFdUaws4IQTibTP
hUx41KqwuPDBnnZCklLtkDiOujbvtTAJ6EBH2mGl/+Uj3QLx1JmuKOSvDhrsBjvn
+9OovJAR8MxeVSGMzZCco1kXfUuld2So+7H9T1Otzgj09gqbq2HbTI+79eeWURlj
YNQp82gFQ8CEBB6n9DRTpAPXWHPaaHEjE0O2GYBXbAUTGUtHWCuhWr1OA8jk8duB
0O8oTX1hmIKZPjCeOR5xt6VPmlmQTnYv9qAlDWqCS7WQItWW2IQG2GV2+QwGTYVO
KCTAmej3J1l6MmreiD2XbhWwhw4kyb+tSR/xhr1/u6PTcAXNy5D7VJgOoC7t0Kb3
DH6XmLhIbx/c+0kVN1aopBS5BjuiOHfL6kLBxUtM2NkfAwfK8oV5ZKLW9TaYIhe1
hlbG7KJGIwl659jGnpQYI7gYHpt0WP2Sn886lVZjmF13jVPCL6rLduLUrwSAZXG7
EB3u6/vylsuqAkQiYFmO5yLXz+G+0A4XshNE2Gq8yNkLmIBtwtVi1TbyaXuz7BDS
4lJgFAsQPuNufqxptyei1Y/KYjN62Z9nMseTS+2eHbI5/qiT5sNMuhuxt4RuaPCb
xrphei3OnrUS3da9mky1zmN2tWJ3bZ0KmW61Yeqfly7wkQy/P/eAYvAUwMHMmQ9x
9uja9XzJ2O8KHCXF+XCffAZARI1yvcBnHo04mKT/N0oLldZJFz9HEK6i3Kob11To
lVNkUIvdy5Awq1ON+YphCJIJChX9eKBh5rmCBWq/4SmnWw13yIglFvzV3cFNvi2/
94MTn8FiA3AhjNgdGjDtdZkwiqoItPJi7l1WZLYhIhS/G2mYFz9qq3O2bPwJIO2e
JC4dNLMP3cBdWz/r5u6qCjP2ZKnCcsNzmDUiP1zvVLEOtSzU40RSNzn6RFPhTi81
rutGBXf4TDStPb+Mkr2ud5/Xgy5UqBOnCoIOxLtefqlsyK8gyZNRYoFLFPfTFFhN
YI10lDhZL5TkbgunVdn4Jzxgyp858U05iLdVP5uRZvY2xI38MvQ9CfBAWFv5Ss1w
AxfW5C6xmGj28OM4JWe+4GqAiipW/ECCw/dyr1y+HOxPwgufXCOlDl51+MhVJNSa
/6jJ+3qFXd0v0jBGaSpCl1VJwwo/nDdEpZi6rfSSV6dABWjGRcCTT6ys26lHF9+I
C4bwWvCYTaATLEEBdQnyILXBON+Vhk3eGgJlApXeu0otr+2fiRBCpeNtIIRR0/9C
JrbRSH/6UviAEqbTclgzMIdeIJHbkdE8h6MamqhuIEhBWvyL+U3ggKrsfhhyA6w8
Wk2A+Pqm8+B49Y2HfK1M/DqlNNxWN/mH7tdxV5eM9xPrGOgkq/oASqUqQdXUBaYr
lhyfGD5Dmftn1d4Rs16zid/PPcWCvOeK/zcWqTBXzba2L+PqaaOAhOV6ivvylD2R
Zx6o4zIOLZy0qPtGGAe14rqh5aQ2Bv7yWcgFvazdrSi4PFzLGoZykd6dPFZ+UeBg
btzdPe6EiOwRFyYZq2qDn/e9fIIoQZqltEfOqBCrJsWI5D5HSHFy3aKlrt9E7Prp
XmSJIPO44+DvGr6GSGc5PXVqcM7vUYKqzudfe2u3Lc/bR+zcQQwdLPYg0LndN5/Z
SPbcOzFGhvAVcJgQPs/JwD5dBmS+NK/FanrHR1nOZW9rGmD2sH0+8HzF/N8lDZB/
AiJaWXruVS+FcnXOzwOc+Zvigrzpu5a05xvqoBps5oNZX4So6QpAkrniNFE8XQRO
NkbUbhNZtKx7ypGVr9U1MQaQEg58uvDuv12EOh4LYeq1YDq35c6nOILIaVLdedQj
nR09WXpYX9H5nFnDHaDSaQ0yjPEKS4dD2uGGdDTsPwirOqnw4BYrmiw67aBFoJea
R5xQK7s9e1ZurlsMjhX3+329d8lsqY80E9qHwqqwRWgyPMNf7gpWKvbfekNDquTl
6FW42oosYAZF9egfbbCoO8JZmh6SASkYaC7eDe89ixtsCxL9+d26RFL6nJyRU6Jq
WILscpiVd4se7c0ZSpfFDXRBDu9njnYChFDLz2wZGxL2TK8DDLzpiW8h/x/50JAa
U1NYElcAQ8ZyCrLf6zM/apJbtKvxuvO7vKqibnS168T4QoFEPVWW/mLuuj0DVb6p
AATr8freuZT1QtkLPt+hpxsOfEz92QaQrlvBpwTIRFMQFpZ3Mpzuhxf+gHKVf/n9
YOpGGjRmNlJk1Xpsh6ytN+8uH7i1LP2ja2tAnnyf/13LljbbSVw01y5Ye6O4eyAK
UUk2guT/OOLQAtcS+rDGolUHVOn+O5Mz3YOlN5ktLvhWg53mqjMQiLyc4KaPf206
6I9zXnsDuQkumV7DuoKXj8JsRqdWpZlA7xUdiTob/d/DeOUTJ+OHzJhUY1bSKFGf
/csW5MHaHIAaMia4TDo9UyP5Mlvqv7Rb30CEX2qqU8FcewFs6sBd5YC78H9ZkcmP
Ai+ju3rlt4vDBfAG1GqJwPiME6oShKxNcFbEeLzzQoTKBA11NjNIhtQv92VDGG0q
PzQR7RDRZmk/+xl2rNyuPNTMugsJ+SUEgDIvuTD99YOLoD5sJ4h/76CbUYwk/U+f
RNSwHQTP6uyIEnSQ4fPok7jFb6cA3nBFF1jCt0Rl3DzLbU+/njhaNwHfQZG0Hni3
oJXw0m0F8Soz90VTiqXSgUDKrI3r0futCYHK8nkAkJdt2GbsQfln4jXSF2qsGjBW
+UmeCxuOJ1xBPh5Qm1Y1PL8UWOTOpgP0t7NTgq98yChR/LmGdgdw+lhPFx4SswCr
dBR3xUK1yoC0sSmEcUGTCQQ32e/iafbohRm/6nCxNViP7UgbvnlneZTPXwRhX87g
EA38lPBYbzSWnQfPF6gJPzacKsRqntQaOJ/c7MDT0CoLkNsriE9wT4HspoLzrHyi
IU8UZkKSj7yIU6MELHi1tYkrfxEeoD+K6V4TwcTBLGrlWVAT2aMcuA8Ir8wrnR64
Ckf+03u1ydpVLN6d01qMp+LWW+wQYPjS7KIHV7g79CIjmx/oU1FAx2i5d+GYhyKe
hGbE/gUkVSNTzbKkScM01L9Bdh/nsH/DuS7/ju1nypPdZwyiEX6C3CHyUzEd7w6b
hsKU7GAkTpybdbhiT33o2UxcCyy9CCLeVK0Xa0EUPE3LHxn1X+txw02PmpiLNMrs
Gre10I7jrrDsN12BdieFTRYMsIEh3r4tWbaoVGzDHvIw1i8YB/5amYNsUtWoCHmF
/RMB7KT8Qy/Kj7NKHUufUObSIPfzpqzfAYX9d9iYpLppTe/bcJ5Qhk4YkvdUU2ei
icJKYlCwyGlY4JE9G1cfmm1q6MXnkMbYbI2258xTrtKHcayI+YG9U8yiA5BDMGae
QTnwAlicifixHDgwWo4vjabD6/bZZOP1N3ssHsu0zXDuBY7BtNGC5LYISoCYrCor
LlGIQVTtpG3E9DZmzoN4wCzgP/QoZDIvIYlhMx7U1KDAZyLDPah+eo4ulXTdWo8H
GVI2BEWJEzFd0Sh7JwpK4V0YFZFOJ6KDUvL0nGmqKXblHonjURG2wlROD7h3hs6Y
HN0vaI+Sde8FLSUP1eEDIrvh2aBT/nZA3sV8BgpbQ2e497rAE2b1JZ/mVE4mRRsw
TPSjsEZVw0XZnrWMvgUpg6Igb82vynFpdJkoGOinH0TuVX4G0KfgXFrnxr9PQWmt
C9wKroRV31Z2Y1jioAJp+IQaSV1M0VSZOHYKermarH5dC4brOfaQWw52odYeR7W9
7xAYqjX8MWlzBZvbZlW1/KNqRdcAoMLsWDNKuO7j2JP9w+0ogDvdTLK4YFCDdQ81
tj91Tw9Qe1gsizgmQw/7kHxEk00BW1AumURU8Wvj6RZrxeC/OgfVjmS82l3ykUdd
2yLToDsKLEkIpXRhy4n9xH7YT5yevRgcsqFXVtb5yaEAEng2BZsuMCKuYfcO7kYC
B2X9nGs9ER9Unv5qS0Bkc/sd/dPt9DaXjliAgvJoIl7G16G0VCgT4R0PcZ8qaPk6
eJ05KjmDy1xkv+Bxs+rS5IPRxghXiKsiC9BrLKVP2P/y5RExZIh5uPvmjW5thztj
1a9647lYJLswvMCl0Ys/UHKGyoNGbZcmoJsEYa6IWze9ATwzusmpMLw79AGqutyN
vaQ99mO63eR6K5lnaEvGbuRuD/Eg7YDmCV7scQ6Krd00Fmbw37VKwJSiY8EdV5f7
MZT89eSNplENECMxUvOdHgofAica4SRbw/OdgQTBfTyHtkNG1qkGRoCwP9sIf5Sw
CSMfC19pTY6okIBFZ43h6MAqEl31HyZSp0VLV2h1vewMsXeYu/aCRweyrjNzm+Zi
8qi5QRIVzZcnSlCAy+1S1GhWQOAQepSdWYauq5MOzYSRw4h832d1lcjQmYh0CsZl
hPEOQyBvGmK/8gF40pIUrhsOLm93gILSvnq8CFk9EsAJT6LjU49koiMz0QVEUyZM
9GUGISJKDQPEtgaqTMSD7eJKOYUeb3iDuu6tHBm2cIzCcVPDQdv6kFAyggjsA2ux
gQ0YuleBtL70gVOvnno2ZYIxYYX9hb3/JNQytDKOUI1OEeSs3vn3dSVcrzgBn4HZ
za2xqTQCRE15b3D4uBy7zXyazsycdZNaFhoHuS1mtIep6bY5jbZ63Bt0BJcBubhu
WOHFFp6Av6EaMo6/kQQon0eklbtpxkGOsSGGDvk3xEgsrqFezOQxd/xYr+rBBqGY
H8sShhy5SWX6zpvGcP1liHFdlKrfE9wRX3ry0Bq8EvZ+BNSXKGur+UjgFWaEhR09
ozuwYAE6lfaPGEh3PfnBZyMxCtK+m25ht4dwyKh3bMRkjR6oc4/i7K1G3B8L+rIk
D85DHMOWULCxzB4mRszwjRJ7JS3FLy3LxWij6r0vImhLMgwm6qVxLaK6y6Orh95u
Ru6sZ5ATx8zJ2RfTpPnz/75LzAzapt9ubsrYZ2cUludYnxsJZ8wVwPxFa+rRGjIQ
mfKh/ONcGXf9EZwODCy4Sm/ogh5KCXQuMJywIAJYhoG6SYcCWSuGzTWFkaZZy6XR
wYQSETkPnyAPywVfG7BstOI+oAamMe/xIAsExMwmfPEtm0gcFe4coY5K3ldJy7mP
5mey7pA2usg8yMB/EqdLJCOYKfsR5U2JyPmhI/QMryl/S8zNbK4ldydnlGPnruYb
MJ/D4FSweqW+PB8dje+k9Ks0l97Hj7rEcY41LKQEjLjhFtNgWhjxBC4vZseQdGO7
yoO167GFjz5+Pu5rMrPVLRDL+ueFHRKk8x2tswHwQ7vxYEKTSS7UAtRzjlAEiDEK
LcAMiScbw/D/xRwzXIyXGChA2NIlnxVe2vBINCo8mL5fUx6lek4WJYrMQNBi1rG/
TMRseBUHfP4GaC3wVsWaFqcfictmw0RbpIoIkGufRG2KaOWMco7qI91Kct3VygnR
JW6I4S69Stpand+RTQ5ApErg+LgRlHa0AOJVkHwcd5eYCeXCgjhlsv+3LbnV1MY/
umumZ7rn3GmIxDCIU+7fJA6CvXVwGpVlujm4d05XPgu+x0zT/U1vb5jB2c04v0qU
RKYz5vgzSv3AxOPJGsbvqcROJbmvsDHhYmucTaL2UJEoUws7HMSxEDBJe3WD+An0
cdNIQBXULhua3MJ1oMymh3pOCA5D2gTHjfoFz0GAndsKKisVXbraixxohegn1rVz
VEBMQpMmXihhlrqCH5xlglOslAp2cNcEDIx88ok61np8UZ9hRDjC1VJbUSEOYZYT
yfW1Xx2wl1U5p9lXePMzMD+b7xIrvvte3FcHHzbQFVF4y5AREfOmzDKBkNjHVmbn
HO+hEa5D+L9MHXr0ubYZ3zQRau3qQIEuCBvvFU2ttg5GqcL1eeXg/dXHFwXkWB2F
FgknLw0QuibiqVoiiRI8ojb4lLHAE2e8IW9dUI0/QpN0LhfDWVqQe/HOsfTJ9+JV
JwVrWVnZwVZiuweodtytAEfBNhegT6b9pyvNVIMCRK0m1N0IfnC4hJmZbaFnpnU9
xfCSO4XW078IceSyR4zIt/GDri/OcmzMYS4MMHiVP/SOv6Zq0A8vHp9USlPHBbEh
abDmfsG5JAlEhgfOIIMfekXanWFLfjL/kuHs711WK7MlR0zZnBxdmdmEFoZBfCND
FV+C9qyjD+w/j0NGZeaMMYR4FS1oOWHz4n4GKpWcifhkTNxucU0whO6YnzIzIvFY
mLtHw6qTMs1gwEl2JN9fRPq90gPQTUOauMMTa6VrcozQGuZLNPnELdJBrxdBQSI9
bkVvEK3dObAkv1FhIwb33qb+wzvfC4sQA13lOFS6DxbhLinJt21dfTl8bS5MAVdQ
KYOge4WCWnpBQs8pgezqIgudtCSY0W9SQNmJph9sUig9Ek2nDqU4P6J+c8VP8AIZ
scz/NtwfhDqgDkl/ka98WfbK2hrbbvNdGz8T9hQ00wIbRQb0ww37NLBKUSZsU78B
XCfXGZzX+JCSUqsOLw/734SiYX4ir9HSXwGvPlqC8HJS1v3pBfb3ZQ8/HOqbr9cu
SX3d/Fat/RLIyjz+SpebYy38CHCv7G+oSDt89pQ/J20df/SwjuZRF6bTjrhcqpJ7
aL5gUjnXWc6BiTrjpvXPXKl03Ape9ly793LoEMfNpd/FKHragFfoFH9501L23Gnz
yyXTdjPbDoQyJEarmllYdQFPX/dVc1v23MtU388hEJZANB+trhTytVUO4rgUsKkp
TKm4CbYrLGg7nKJs2/0lxJT8KK3Jv5SZPag/wVPX6bN52qVF6HikvilvvJ8uolFC
04DpLx7HVt3dJ9M/P9e75Y1DmtjruCxccFf6mpGEO9tllpi0Bb+38AyMWeUSEv8l
ZHxemi1An4+9zmnZcxAHVKNS8wwGIoK/Eo+n2zs8ZBUfD1P1UwHp9QQC1EwSFbrB
gcu1zDt4Zwf+vzOYKyhb50lUrHM5sm55IX6CbV9ovlJbj6XiXSJZ3Oixl8eyMvRb
MtXdFm0Gs8oDlSPbAbKb2Ha12WH7bhP9xza02XKgOzNEpows3Q9xC4hXFIbFKXx2
ftYJ/UPncQbUHr7XwxGxaoBwrGWEPX0Mlm+NBq3Ft2egyaBmSsGVgLam2nd4bQ9h
OBdmYqT+81YMy2adpDIlWoTe4TIdV1nN1Dx81tHDXliODYn+/ErimaPVzqYd4OCQ
yf6TunvmVnhX914WVzxnXibjg5pVsXcQ5EQdPmkZ0kCvdq/ZOgIUDBxXrOhK6Edf
p/SOnUHMxBzX03BoSnaJ9hXu8BOiDzM1/7xKX7GOYZ5eBiXaEcnzFoB+IzpRSysN
z0DUh9c/1HHi9KWbHVZkBywsUS9fxenZKf1kiJxLt92UP16Tetjwksdj234ffKST
ZdO8vec95oG/iXozghT0KkZM+H/DSCDTVHqr7iIaBDx8cusDYDFxF012UJffo5mw
7JHzK69KYvTfaIvJ5/PKwG0uLnarCxSIlqpyA3aYSn2SWOGKGPDXbsb4v7z0aiA1
OsZasUvHXL1EDSxuTNr+xFemISw0sH9N1Ugt+cSSTQuhSiH3rCKCu/mQLyWF8dkj
EKdBhCSe3WnWDhyhs5ynyyqZbKn6QRdVQV5hyhSkbcln1iwMkZj3F37wetiwLugC
p+SaiO3evm/KRIDWGxrioc0CSpSOw88KG87/FR7frLd6ImtJAdeaGxzAz/k76rUD
sAymn5w36sHzDHNlCGpdCteP/vVFiBIgoFTX0ttzWGFICJq01OqpcSfoTLBwvwZ5
vM65dUyWf4vxI89h8FAXx/WkgNLh/3sc9Sz1G8B3fLI6uNOoxVX3QgOGw+DQNuad
kgkU8bRU3JZA6V3QWk7B8Fw89zgQoX/rlfZsSni50PdAcb7KpXJDDlTT5uOh154d
g/N0h27vnIsepiFmgl5rcdtSzwPH8r3fuzQ3SYyktPcdV9T+Go7JIDBBkZL3v3PD
LeBEloG0Nse0Ks4J4LFTGcgjIV+7ZgfqcAGZ/rRb30h7mBZK6G85TlY1HDrnD23y
qBSHpMhUqQXAkLWQs0lmFsM3VD3zfNc6fDL5TA/x6j9imK9Cc6FuDxJJI7CPcclO
fzlcbhni3+aT5gff80HlPIHJNu53fFw6puqw9812GyuqHWWkrLqVTpXUGJ7+xCiL
gmlUIpRz6qJAfhJld/uSgh2Qy+b2FKCNiB/C47yJ0iX6B9T2WyKXvyEyl1vMtHvK
0MPdye2aaLjy2UAWRIpRvHNCd6uDVUgbnVTVxy+wm/VKRB9Nzm5gAAHNxDYFJovm
1HOb0ZPJt1QLL128NDwh1jB6wvMT6LxumuQpcJFJpjnIOUFm9lJLlvpILUWu6FSS
aCsThlgcbkj09pxl5Pn7Qs6g7E7hVcrVJvCNRVsubvBx5lCNaNwHU9gtnlLqbUe/
miy8Yjct4aYGngD7INH+kgqX26JoJaDYODD26PzSr6lKGFYilg/C/wJ+xwp2SzOZ
PY482ozMyrerYOu0LOTfUS/RgttW8QsEeQ9Dpv7UYWx+R1LjazxhLkL+h2nnVNuZ
AUIdxC3rpb/U9ian6wcGdX8whZ8cmrT4VO9kOsG66axEBFqjk5uOFCN2rtQUrs2X
R0/iyh29Xth1y/zGsN9BePu3lG+SUG0/9qM39PFBzsghLSsEUb9uDa7Vj8TCEKWw
saGMrGa5Chh+SB31HVDT7Sz1w7ucQCNxsaFjm5Mvf3QSJ5WHg3wMrUxgyc3OYQqU
KPc9ngWB24T2uuF/kzhWOeqCnHeQfaqDx+Lx7hI4F1WtJtnhLRKzvt2JI5Rpj5cG
uC96Be68Disko4vc9gDskrYp80JHu04YQMJljel8vjDpNSA/BuBxj6ueWPsC1/NX
GOp104Pk0xBi9Rm2vEYYxXD/+Hq+OHc65Xe0Th6d+Jj6Q3Syo0fn/RM5+UrnL2DP
phmC3hM37+HNLrY9JBDLmfPUrkgKd5rfZGEHIHqf/znb6KfKmm9GI+7rCVg5taAQ
+IDHRmb+k6GwsyoLSAPjJv2EwgpaDg8NHiJ1nt1I+Bpv1Gw8rKUlv3xxafEF2U+Q
TWgveVWPx9a9pdDhADDjB3MqsT/f1DVIuoQunzxpuipAETd4oeN2Wl5gm6KpOrxB
7Eor4Yk70jA0T+Mf+r2zBblAoJR4A9IKj6cwwt9YrjSx6RKEV5eUAwMWDGg+vYdm
NOeBIR9H0xYuPsHUFvkrIzGPY4uhRaJlWOpeXUZAfQNjl4oI3qSNbhmECSS/jyJC
TnXrC5dzurxac7gZNvdRIpU3tFVxGAzI/dcXqhGuphMc5+e4iKHd0V2kZf3gVZZV
2x/F+G0c63Ryetxj2RJ2w0LG4uth3c9OImmfNbaB5jXc7HNcGxIh8Zj6tzp8W706
OQ/aOPuhEL1xxQCG+BMsKw2XSjU8bkRk/M/kpsxPy5RrcH/dzA759x3LgifCebT4
tn3G55kldLFFVuct0FxivHvICVL8/tD98VljMrR4HQz5ilNbZtLDWONEBubRVFf1
z95Oer1ioJqz0xwvWMI02zBGx+m33qJCtnilOT5zy6Eps3DkvgnoF50zP8ZsDV1R
Ne8S29PMUwRCYgH2Lx1NucicdlcTjmAqBly/8C4B/4cgzRYll+vAxK8P+X6lKcoO
Cn3ZNrdhayVegp0feOMX3Zeyex2L5hb7JAtReeCHcmVO7WPWhkhXn4W9o5TUeSNC
QvL8Acpq3VJkmmFuVJd57eK2XcQobUZNJIglkZddPD8UcDeBqQimsZtNB9tXGy5W
dEwJ5hMqG02ejR9IzzBibVMydpSvDWkqeFBNsBrWwdDcdx7CjF64vnXfSBxtNPiX
/+ErnQHoWv6xEBXPUhtHY+YWB1mFhYlBR+UwSxsbTOLWqSjWbeocb8kPPDDy3HKP
78X1P48eFNQ7no+FRNitC9wuIxHU7Y01Qv7J1Tz3TpUZWKHP1ONufn5ogm4NNDkV
pGLvfQx8Q/jryJbSwYA0vQSFiCg6itip1oUyafNBXkzFJ+tOQ54Y2r40ngqRQ6fV
w+IceN+x2tNHawSjav/g5XTmhhHfiT1PJPfhMAlWA49OXYjwttnyKVnvXk5I71Ax
fItDRvZ+QXvAIoI/88J8oFN0cjh+mXRl4zt/5/WQp8+Ouoq8A/eoiwuNEcXqIerD
vgxuqtJ5igrRQAsGFaNdka8FogaIPJtKgSJY43suajV35IXKHgUM1+DE/Fq1QnqV
mBzZsY16whOzkVDxKewPrMmw9o8ODVRueukIXP7bbALYixb5D1oI/+qk8F2G7F1Y
neCwTC5QOx4SsBtt43pRCm+7/oDwtZx5uO4RVsCz6xsdGGv4e//3QYfDEaFJISKJ
EV+t1esdAN65cfVy34cLSWo4uubMpsLjnSacI8jtU7prLp86sSf2y1TOXBhkbBtL
5zWXYkrDuyEzoLb1OATo3jdvz7MOU2bgnevs1PNnI6hzRP91y4mB8c0bVNZUrHuq
kq5TDDO+PjN9YZf0EdOmKbfV+5ehgQ93WV/PFATODy572gvtXcvYJQdr/rGxpOPl
kBtObMzkZlkpbET9ZxrLmQrwALFk2Tc6pM0HC2rOuop3XsdLrBbsuvahF8UtIjzr
5kb+hSbxeXpvaiUgJqv/BFWiPDCGFj2A0HApsMlqcE8TkjwBga0ZgCx8HeybeYnG
oTAK4Osb43RO5g+x2WefSPgolXBmqVQTUzyiuQVnGvfKja9eUEuNYpsuEIJLL22h
DFN+bdlGgSVxxUgSLz/9IqHCXaUPxmWly0xNEIDDVPrLwrBCgfcKxPEvP2ZbGs7z
rckQRB5qVm7zYkg1aBbrMIwjHxEHZcpfk3Dc6b9rpSQgs/jpgEsfbfOUzmWL8UAR
Y1tMeIT32646OgzMuQCH30LJwb3i1l4pmJmWCsL7mQmhfCAaOYa6Kd23Qgi9G1+X
1Cxdc0sYnXvpLpvyum+Wtll84CV6xziQdfIEWFH4ZbQGloQFczWS1rCuZfELsxRY
fTC2dPzJlxKX+dSUgOWsr7XcsCER3AVx0EbXKPR3N4omuzyR4gHF8Y+shb+hZKmu
Nja2SKDR0+Q78fXCs+2XvdOCjudG1OtMl6vvlmGsObNWlyollMKajmNhF5So+zTo
P205ufqPP0CMNQXk9g97V1GTGok7UWzdMgrb2ZJdz2cA+fzgJVm5TMJudVq6U4wm
2ZGJEOx5VrJSRdB+9fbwH1N4wQwIeRYdcXpeSGkUmlhPsFccM2ejbPnWnRny/Y7k
5ghREMe31Xol7V2pUq0ojQG1NnZBKstaKtJaxqYonCFgAGXwJoR2zc51B7bBMbAq
3H0PTEoebZ/h6Og7qlBHs6eNEJ4ye3gHGhMXHI46cQq8gnKdoS8/yQAk2AKrpvLO
uCTfijidkG148IJtojhAJaDrrs+NXMzesVVO83wMKNBKpMZzAyC0nkfONzJSy2ek
BcoqrA+AX4K6k+UxmG6V3vMMdkT6zcMiT2DnTH3QfOGKS3GpeQ49iV8l6UzUd1ec
x3ikTYZSPVllyuEob+lWP6EP5m+F3ADXF7sPuDhrO8pOCG+sKDi3HN9rU31cuaeB
xa/+O+ger5WSr15NjaABwDNrpUp2cr9EULIw6LRdEhhWjaP8ECszbUnbjma301Ye
kX4fEEKS467IZWMpArLChxjA7ckomc8OuSMtuNKjqXMsgD7e4zQpbrtuF8HyQgza
VEkjbUh7FnKTSsiONmXGFPBy59t1EqFZ8zrO9ZkFv+x1X03Q8xt+Y7+hsp5Jj/ge
J84wwNAaPd34S4X1EQspjS02EyxZccgXelDW2jZoo/BosIwXxVmZpZ9wkjPnN385
GDenwzpJjpkbxeXu2Qo5QdKYqHGPm7gHZxQm3ClGpgyRI9mX1+84JazDwP6kuuSd
+T/lBhlcv/dOtXVRwMIGHyrWWAxxZISI1welj1G1nWdErBRvdUReWMnlluDsczR/
fT2/DA6RrD8U1djq1lzTRJsyrVzasJi7Im0mXxJFxjdbRaN2REYWn7WrIo2uHKF1
EtP2cNBgAuvQadj7IAbUBJBk57wqpZ6yYFYOHPgIyyq8UiWJP+mhjGu2/x9qSTpz
ynIkhsGXTjuMfWq1SMdICR9ZBOVuNc6bh/OGCrZ50TiOeKFKEcqgydF1lSku9Ro3
y0CLhWclcqyRT8RS23y05qtr33BLdZE5lLpHHLeLT/cFk8Zsm23Rloyb4pihrMyM
yZUxKdjb45P6rKgaYREp9/jK4lripev78wnlfU6hZAwE+TbkIxA4WzDXMc23QBUK
2ObqMjwK7eeJdoOxsgI7b1BfTlIDXBbz1cyjREaWBCEgcSWJtN86F6VihIqwPFDf
44LeY5LwQK+sccshoCiMPE8aH+TorFJVOXI/v8a0c/L3ZlRPiG55m+6txEMzamjn
aQMrIXbybMDcE9qtc5omd8oAQAM4I2LlspwRxB0SjrSAnRaDo5Lk8xosIii431fT
Pvw4hcImKAMUZSvUFThZELK7MwgRNyVm+p77CUXmHUkXzO+wNbPtWOWI5UecPzG6
yP1k4oSE0iskzhSoP54uxJjjBSt+bI4l/bv7xQtGmAkXlots4pWyKwcwlRhEbhrw
4l6Zmmhj36gZDdar4zSmIybgH7pjAJKrHYxNDgPJGDk1y9uxOf+kQG7eUoipUlVg
FM8zQSGCyB7CiMc2LqQftRNha3qwMKVlZKoIYOyAjvpOfrTgs7kEn5btaLJrJG1k
tRg8KImf2hjBWhYtQ3sCNy8ubGcXnerRiLSWOTmHwUqKtz7knXBvlsGWzp/c6SkG
ClR2dIoaU/Q7VzO7ZePM4K68JXcmlGYJ91VLL32OFzBGg50fmRv4zpd7nC9FR4vl
hoM3Vn2t4QLfBtwqpYLsCZMruldw1+IIa7b4xvu8lVN6IfHQ33VxiO2miPqbrHdw
Ba6YvaQy+c2RmogBVk0p58f5J+cC7Dp9YRE8+cQGOd2d8FGH8HaTBlyvQDFzpq1X
h5Mea668HPjKWAdEHsCKjxgE2Gmvxl6nLWu/zkFfdjwUDrhigTPGGrkI6VK37Atg
VRC0cHMRnvl6va/DpAd1FJnlSsLwooCd60t1veWzP8E+gXZ+AnPOZYvtlPClvXn5
mP3N27KKCtvAg80ZBmF0SxpGOZk376JsptO/r5EXc39vG/IIvPuWKjKajg1+JiKN
mGyFv9wPyECSYQG8PzS5HnxxppNt38fH7oT6Gl6/QtuIZNj3lQsA4kV25SAY05rd
kDigiqq1smYp3rEiq8c01Nll2IwppGADUSMdSMjMeq58vmRGPxGJkEqPvbbSjthi
LXchj9vjrUivhnyrvzs5KieGQ5ziCE8g+dm14mdTubIkvW3/ruZ+jOCb6jF+m0tK
tx8Ch1K3lV4tXEXQlSXTnEtAReyybo+WjciqOX+SVN96DpcV08bKrYxpOHiLBawr
6QevmZ+pW8C7bkvsAAuM7Qm0M1pMHt/QFzAWge/d6yhMm45GExy8shfRaLJXTzc7
SEA8aqcNTP8IT9BIbOASonaNyWal+FOELuG/Lz5RiovMOR20BZS9k8mbdi5oMpAT
SXB7o/MrCC6LgeA5b2+6b7AY4bGiplqp+cY3X7oK+nhIW4ZegR+iWoe84o06OVCi
fd3b5bPUp92qJrBeYa/KGhioKfJqvsSS1MQpyfYRpNCnClLQvDJQV/Y4fL5EiDg7
l5t7fUTT1qiN9YC0XmDdS39KEor7VrrYZif6wjjOzlvq021mHVy8YjvpqokbbAf0
oywfLxYKOOAowLhe37PmQ8Z/dc7Xi6otzHRXkoDiTMZ9Xja0PRuopxGsy0ZT3kAq
nL0iSFNmo9Yj/sU+44eoeXOJpo1R5awebsz4P3gcuhFRCMGfN6/DpChb8FF1UZmw
betxLd7AgQWy6+Q5fM93ZYpAJUXME8o93SezeDMPtVolsvGUTuol44aIaMM4eq4W
99XpwH+sp+oNdgjILyB0mvYXwc7q70W8aJ6+1tv6y0eNxrhtABkPaCREZsjTp6XT
BOI+U1cx2JbiaS+4DnFC1u12BzI44FTZxS9I9lKObwx/8cITWUJSXzLj3HVhmuK/
/Sj5ZM8qWz7uBtJ+Bhip8G/kEIVfUgsix+45SlC2JkWux5s/2x0QvZ6n9+QufwuP
gR82Zo/JmVFVCnN/SHkFKgKEV+LyB7KAkSIilNabnYNpXrJmMH0Eya2c6HryyIHB
J3Z/HNuocruXVHrnik5z5uk+njYgkSkWZIeeKBW4OwogKRcQiJIqZePROxe/+n96
Y8it0ZQmeL11Ky+pYqOxSIau1iPWgYLnfoSG+S1FOIrJkK5F7S0ygLY5fP+hlsha
/FHYU9tYxT02dKsrxoQExZ27qi5yz5Wl//b6pJhbCuREtQezW34YBlQMartNDPHY
rzVSyUzPRfLZqYn7kJd0vN3pJF8dIcW0SZt4WGK4wLyQpjq/hqL1qS/0Jal4+Szy
2lh2e3T/HbyRNcrpp1Ier30zGma4H3P+6uqX4IJlQNbrb/C7L4BZRE1VC9eXO1BA
v2Ly6Q3ifjbxjFEFWk1Fye/6pUI1TdtsfCMOJCUVtgzCXzXeqgqYLnVhMzk89XPQ
Q9aNh3rWRlx0byuRsmFghA/bbQp19U0Gs9gC0WjJfvFe93vGmD/crjMeSvWNubzu
2q++TDrOmw7ko4qnf8eQ5UUHRDSOidDrU/5jgoJgB9DQdIgx/80OHBTSb9+wnaB3
JGhdTQHb4lHnt2cZtMzAwleN1a3AKPOV+difzkRbWhEOrAr6olDHsFZskqWKWs9a
Z+RLJf9Q+882X+55yFC7EUp7VDJLm3jgEGHuY1dPVqSW3uwyg+mZXOl5FWyGZ/ti
GePpBJP16hMvxA0YX4dt4XMf+ioGV2DJ/ol+pcVKIU0i5OT5DjUuO54s2NtGTGsb
2AJFrBGdwrkgebqM3P0uYyjyw94kvZ89kXZ/RdYjbb3QkGrtIHyxqD2TxJh99HRT
5tfhkaGWV7fd7CQOzxrlnlQ1tGx+6xsIGiAiRp+nOYDVqgna6own3VWtn8dcdgU8
avx+WidngNs2WSz6+EdyYqKb+q+Z879RFDV77OjfpVaQRy1GuXJIJBPvrz0Qij9A
Jd+lOO2nRZckbfwxBEoj5qJIZ6/aBGGdV9rvKgscwUaKHkB8SOsh7y0goTkSbnfU
3Q4fcPYNeidfbOYa6hRS6LslmHlZ0iyP4laL//oh2+8+5y67mWPbxhqfxmP8D3IB
9rWTGQgTpygqsK1nBD6vD9oxB8/TEkFIDTJM0wktJjbc88k8Sdz72XqG3dZ8num8
5a+tSv0n83cX/vNBIoAhHJmUqahL/MI/Y8z+cWYaikWhEObCgwzLU5/mJLpE84Sh
1lTWcSb+h+Oo98CKKstAVYQoxXAF2nxFXoLoibygWnfsUphN6gUEgpPrlOl0Wqah
biaBIYni7Rv2znP/lP3lK4ORv7JYq8VHcQVBFkyTsmxrckChupHbIG2oGlwlXjbf
xgRBmQHDvRBzw9unhRQ21AgRBFvYu91De3zXJUp/wyXxWH13uTgJ8E48o2FetCzR
FY4v5cY+UmzodSESHe2AziKVLBx4ODnCAkC2N+3JlrO2lIfTzFJkW3wz3eDAEjIz
IdpnX+X0yCAEZbcE4LFBW3YVpZoX2iW+WrBnBgyMBUaIa2bNwqvoJQBuMdhHQS20
P3qoA/WMsq1dq+nerVTr3HD8cv+TwB7/FAczpP5bAmon6H8NzPDVrJSuTToOZ7Bq
Wv7ESG7zoA8BgR2c7RBrw5yp1Yrs1Nbv1XiBP+HHNHW9za2o9BodKpqkPyr06LMe
zBg3vnRI0BsOtB5o9WrCyS6xwRU2DH0xpfLp5+TVsxu3pHLVerGHbiyj/HJuL+n9
yS1bIzfFDdIjeSlrHbbO6+q7ZHn2cgWgBwseRNpAUiqtRVisxGoIBPzZEe8//mXn
SNrh3m22eEIdIlw8ZEUr0b3Hl+Gms2i3Kc43WDgVw7pQHilW5LnZcM+aIfTjg3ae
lFPR1CWDLpCnt86ywbtgwRdJ3lDf5UC07jlMkIC0gLvuiXNcln6PjVf91Fo+AbK8
iOn0YVPZwHZQ5Wl6ED2BtbY4TLu7xDWXeTbdQd9+nCcPjKPAgKp+vTRrrhQtMfpU
VVB9thQ0/JxAOQ/I4Id3giWDqFWZ/drpue91GPgy56h89iwJ3+v8U63MMz99tfvJ
wfS8PhCx9F5TLMWzMqnUYVLNlZ4qkTx5kgfxYyfThmv3jK7cz+of0TDF0uvlCClm
eseLvlN+dUUr/LYptXDc8CyFN0agSVEtb0ih3lKrZ2QfyGfolIUgQI6L6xkxm/Az
gTu44xT/ALzik3iLSDzCsgQGXYHI7kymjMI+RI5z0cGAXOgXgJz8x0TccxNkeHaF
Ga3XeJmHrkOYvG8U1orr9fuHjLnynUNDQBaL85XZ12oGKAV2ZXO2tOgeKD0LdtG7
fT/+N9hgDpWFa5GL74sGH8Yr6Jp3LniYYgMYsFmohm9zkNuGfv4E0XO60q7AUuMG
8X79BbVbLGJGOgtPPAbXR3TQGXgkBu2eSUqL+DowHDiqT33wKK0/FaxrQXl9icHR
8PHZkGRlORhQJu7trKoWb4ja8F/P4j0AYk0vZxvmGEpWG1ESdWnuAvykcpnnDqkS
oIymnLAc18g8KOCHYxMdIWqci8A2DYVTNRTAZQylVrkRkCDGN4owYsooX/fFjA+l
pGkX4ou1yUL7UkUE+WQewJ68P72HYvcAvXejouYOgm+zuZAwSGqCYW3hEUsPwyli
kVbMAqBK2sx5E07j/HCpWyznxgfWwZxxWJTAQjLQEmZII/lMyh+5bx7mlbh+prGO
WNHZ5Cj4NLrE/vDvuVC8yEOb4O4qJ1Gn9ezjjXsbmnsRRf36v8FDcQA2BA2VzVXH
6dfulLKq1vISEuPsmcXVwcd2zV//HYzgWumQQ3JGPbn7Hl24zNaFOVRioBMcLCrE
BttE26LPi/LqbuUOLPhe1semhpvzfV3Ewn7ybgztsyOtTZ08GZXmaxnnMfIGPgfj
Xw3OXBW/mWLi2/8XWxMqRT3EniOOq7jYlTT3kjUGWKod7VxNzgH/yT1bFh1HE89t
0+1oxAEteiRrHqsUy1CEyAnTyOoOXE/enDlScnzl3EKR0edgtUigjgaEKNOGSOCY
qZmxXoBBxBCFUkzLxQ5a19JwtIHqwzXkfXhE3Aj15981UrcIQjFvMq/alPkALjoV
5ekDjullb9TaumZCPKejQ2xAgdARiZiBwJA+u0JUBhpAhlg8CdJmGcajNVAIgP0Y
wvTa7WAs3sk3Pk9gqOWzMD2zeOnxsc0PGsf0KwAS8AvcYdqxlL37Bb37lujqKZ+F
dowePdVbjzbqaMDVdnTj9/WpxA9Xv91j4y0/T1AAGPhA3ZH1sI+sOtMmErm3El/G
HU4zSCgdLTdl4FdxSloZ/ZSZIDXjewIFMWi5MjTjwY/OK3VIWZdhPLGi7ZyWwDWj
pN6QeW+Gx/GdjlSY3JDyXH5c8J7iJeTX+cQ/RDRVsGLH9yIOid92Pwwghj2E2UX1
nmiqkoQaqJaF826xtmpRiSJ97pDoUTbVsiVHv1O1JKZlbZSrIfzaQvA/gFUJhDI6
lawRNmWZaOUjJD1YbY1C13SDQKX3AN4z4DN6+GNxwxQ0Zp8IH7IOxX07Yd6xNMSb
RfYlrswQnCWjhn3UA03wi4PAyxGIvCIwghwU0GiMMxfNyU1QLE223wuJPLTNbLpm
CbjmM81dtRZ92hXLHVgkZk9hS4HG5BEok6kn7QDzc3iUnLSYVreXzwgyX7HMmCmW
ZU5CrRHqeZhuDW/PbQFNVrgXxirq2fBxzRknB6XD6V7dTIKYil3DPaAlHiI8g/D/
q8Jviby0s2TAUQSiwv6QNPmchYgKWRYdF6HCudzTO3uvldvLehiqnmx5QHf7HisD
yJDhEEuwyLxlhtoUTd/rNoWdX3m5c+atmmGmEaPo6N2CPBZffK2ndmGTLIP4kOvw
YHP4dMxHtNz+0xqlUWBJPyeY/R+TGH3pg1UoMvCde2rXFOqH9b8Xzz0i3SW24jsb
OPjD91cTRpfP/nhi8byw32731Uq/NmnqLpVhPPcDWscttKmTHiBVbdmB7ubSLx/L
TrdYpyK2FJTAGmbHJuKbRCriWpbC9MGsqBfzrQrxCA0YwcoVRi2qmhL+CexOKFw4
O3GLtlsDuAfLEMDSwwT0Xd8zmsx/MGtQwQwwj94WpzPZXYMlpRMHOya3EUlYP4yv
ay7ztbVcJ0VQDHnygFzbmIvFNMkoIt09biH6W/CJypb0i9ZQDyEPs5ZdiYoPG+ng
61w/IpzmvXAHygfmokMfssGPBg6FMN6EnepR0EfeL7NLrvY9l6ipbUfTnwVme/oc
/Im3drPelWe++y6DT/LncojNBfEeu7WU3YSwpX+OhzTQuneGKi0epgFUIxft+ns6
CK8WRZ5VDn5lLKhnj7N9azll4fGW9LeaHlcDvqA28uC1Ke1rQ89ANLS2EUqJiNVe
WXu7mM0xVOw1AYZiF+bs9bx6Knss3u4dRXv3Q58nr3GGGIjw2rbhan0f3qNp/CGi
0pJqBC3qfOuadKvqOOLBGw5vw/BFd71D3AMjHETZaqSVAI2ZpdRh/jN0Er83WcJC
MZnZekrqOrpdHGJKGYSVXpI6fLKS/pa8d4L0vSSZlzOpZ9mSsBfUbED9DApkgfUR
y8WNKpz6wfpvoLqdrfKfleURvPag5VOSLPwI3PryTu5q1UUnzs8Jj/me4nxngzr2
+gmqvzhr6iLmVhBY4Ffh0WZ3hm+1p4/WInkE+Wcl0Zo888EOYNxaf2qsLPIN07i3
PDQcn3QjYsjADiRxzKadrfF6KgPcZdvPga0bO2yRo7XaRS0NUc9c0aq+xpdeXdVK
7sMACE1FuYlqvSnnqyEogPEgvLqnAoQMYk8ZrO5CtP/A9O3b1PvWRk5vwfigt/9J
8sLs6awuYah73jhZpWhqf+8Qj/y31+rE4poeuHQ+lAClZQCzishDNGtJ9CKF8EDC
ZaCFDOvuJvDX4W8Ya8FHQE0/rU7xvWfStqttszd9mvo4F47DO16YfeaicGsmvgB3
SO3e9DtvEQRw+W8acT4gJhDccq0fojM8wW/90/FNT8Pr1CkW9ehNxGqPezWJ2AXA
4fXPFkjS3PnYI58NfQvG02jr9ghGdRc30INeo/SyYSN3Cx1yDe1SXRtOSGZLe5HS
rD8RU8XOw3a6WDGdSKO6uR7cLV2szCM92npssw1hc43LJXbnMZFCzgn19Ry2mZ7U
rUSpXzXHepMT7wEUf/pPEqmt6F6iQwMppfLD8gxBipAFqUnmVmhswSwYPqCN2BOl
53qLVc2Ul/oFEVjo0essVT6FX3obIBLCnUYTjroU6fsivr3RITEgsADtKFKabIl+
9dsEKsId6QOnMARp+mr2cfxD0ZUsVMopZacRBh8u4LeAk7EkWFjbLHeqNzrWThXT
wbGS6tv0Kc5Xo/znk9Zq4PyUG4RHJNNV4pHkISVPiwBuKwjQGLwneUBFZjUkhglP
El/tWebZ65VqVicUTxESNpedaXkad2MVvZM7p3XWt6nrRxoJePRWj1dsL+qzPunP
gebsWOCeD5RiiOnomlDp5MTMbT5xwqHVkabrtIBtLDh+MHdZfPdge2WlEWvm85fH
LadxGyGQH4rRAsusC0EHQBZyZ+NJGvi24yPBmvg8ipjyT7g1H/80vqqrrNBD04sv
Qr1IPOqvfmnhYwuLn/Qn3vbni+XGQkRnrq3LupfzWED9mFQkbCXm04qxEo/HurFq
3/VHIqFxWC06KD+zMhSFNPiszxLVN7/r5tAYoIMyKj/hJ/Gx0uWXoI85TV6TSwxa
UGSCmqPJshvqSmYelq7ot0NMcKPw3o56rmiKLgDqvG8T0n0jNaIgEIq6LE6vnRV/
Qn9MRgKQyEM75Nkk0WNzHJAQNdkTzLydrs1EOOIJ2EtL570rGFKYGFj3MAfqaAgn
inFm8tLET3/8QxVaM4rfvvoPMyxd1yebwIqZ6WsGfVI2N4nT7LBO3PUBgzCDMzPj
0GtCSKT0+6mkB/DNMAmK5LG4CDcj7/dAm49OXF1qRL46kmC7t+QTqAZpRlOylB8y
u1e8GpqVMgg5rsuGCa0savOtKev22QT530H+Cr1+Bsvy8ItaQYo10VH4t+IiLekd
JLkDmyBqqUV2QFKl47jMcOWAOiMzIXaycnIwVoxs5wxzYADZ6Mg/XBmApCtrQocl
6am4urcgDfZuTrz04cW7ULtxYwWm66bFj5xO6xIPfNUaSYUEaOYn2PWOJ9+fKNaw
FdfhL6xbjs7OaCFOFQu9ZgUmv0AyYsff97ztSiDVo3NSONRvl8ozGMcRJyP5avaU
tZHYFaMYx2ZXpLrrPgmNYkr48iFJZnpxvlA6Z4ERE+R2fEFXjG2D2Q0MKl6aS8aV
3znY8zGIXD3wtZirFNXijZ/dN63EZyOrUz/xCkrtTHhrCeNOLqFANfhdEBz0a4iq
SPuE0Y+iIbb+HOLSs8+4YLgT9J//pSeKBTfaRk8kRDodquY+nj6RPJv8u4Lt7nNt
FpXr5lft5dP1wz1B3TfTZulhXqH7uwy8qcFgyxFmMBkQl1sykvnX4vFB8wucMWkR
AVY7xeNfrDS41ufC6JDF/qzwSEvOCDLM6lhmxxCwjCat5sMTkoijpo3zKQI6KLJC
pUOSow2TD4YY/uM7LUpnPDGLxJIB0OsvOR43taKZ/q48I9Lh+HLG/h/B9p0nAqjI
tA9UdvFYzwwm1i3lwabt7FW7Px9VorIFVCDlgJcsaOKJGFofrmqOaCgWhoy2Dhh8
X46+Wgiz9T+Yzz4/LejplO02F30Crckl2cJx31fVWqJScGCp9ARPDh1umOPSAPn7
SXJyUg76+MsKKYLSh2yYJAwqV95DWqCgZQSwNB1ZcxJdmTYHvn/zOPhmK62vkBO/
O4DbPZocsY7RbqDQZP3ZAPgbhjK8FJDOJ6EvDAc7ZG9sXo35e+rqoIs8SUywQO4h
Xl1NoKKzxTMHqSLDDm+6c2rJiqsgWQaBRHU6WgBrteIMmzOBhvyWpYZ7+PHc0/3L
iXZIFu4kCHMaQJkOvPhlGU8z3LGW/DSJpquNUoqKhG9xhp5egz2M3MzFg1yj5EPO
Ab9zLDUg2vuUyZsoizo3WmT8CE9/QC58Yj/RFGFAAbaikKqxo2Tj/HRLqfnfwDW9
OScG6W/PCLdwpGV9kN3Zr/9lyQdHddSoM6whYgyLZAPorYv5tqzEseCi0M9r5K8p
g2xUshPlyALTw2lfkcvifKwjYNfE6qtXucwTIlGRLVkBaPmstYno0TPojSKQxWb+
GIi2GdmEZNkbxhBigBQkax8JIffDM3GGUq654TWhMTTnv5gz6VXWejZCjUxy3YPu
as4Edz1cqdmlajuBCJuGLRa7hsQvDyl6K93PknhC8j/DRlVpWZA/Bd1jWx1iT/xb
8wk6UC2mSDzCwcPHfIVxfvL4rEAZzQY3vXXk1Ut3vC/uzGShMbIorbCAOz2ozjsa
jYMiF1hmF7LiXbqntQwIO2ZP0Ah5E092MgXxORE7fhDe0QXNxN8QZa7RzR+v4foj
r8/Hx4wrxxdAW26Kap5x9Oc/mmTT13SWVE8Vn3qecUeSibAxPoI3BBg2+z4SOm+e
Q0K6LHEuP75Jkv7EsI9IzHf7YTjT9Ob+e2w1F2DLt5d1r/b2bew/Ob+L4fsidVf8
d+b7GnOFGzeVL2FY9Nhg6vG+CBvwvELH4aHs6SmHZOL+5d7rJf0vpv0Gfp/VeVAK
B4Y76Cj1gj6m0uH7oPy/1mTzjW9kPS50XedzXOJ14WL8BDjPmEXn1sDKRmHsB59n
WTNYFFzC3sAnlHrjN22NEAa8Fq/H4rjB1Dm/n+wcDim2zuKunYTU4cQSyZU9kzJZ
eS6o4U5rZL2tkXRG/yeFcMnANHU6V23MhfAM8G2LVhD6LGahyo9NdGyKvqsmE9Fc
r27h+hbcGVSbOMXexorJh2UPLY82a6m+CgtBBwfL8XlxqeAQ2hYak5WiEv+yIYES
hn9z1rjBY+awH4bJJf56QjaJtRQXMw/IiiMS01dmne+lN2knRRQbgMqUgK4orI79
ylspXJUPrTDL2MRbayNJfeLEl1upC5gYkO+5w5/8QRvc4GFrdsP9wo6FC92SorxH
6Vl6Wz24uj0wT/jHSyBx9W/S2JjxJ8zGE5QZY8s6s5b3AoMsXNoHljLXyI+PVmFO
8yc84G0Y/ELKN8N4KoMbl/gTgt52T7et4d8qI4DOi3LMTEh3s3pBrB389UI+T3Hm
pSGI7RkXjRnfiG100FHUw77yplcfLPD0Y16PE+F8Iz7pvyacFi5Fv2Sl1i4QTI2r
Erlcy9rEWEAckcqgCEgEp/UPSxOjPKVyzFdw0SUiIOX/vxn36h08r8GHYh+QSVUa
lJV+Tx/5hFciMmUgv4BkfP9cP96EMOjTIadT2B4Jz3s8ZiIcWLUrxxBS7D2aDF/g
vQz4Y+k8MHlMwoZXcwf/2pwymAf6vwxKPyKh3GTIRpifVT2N08DMWF7t0EmHJj6Y
DqvXi34gVsEPV2eCP/ine7Mp6hMmgTWKwNlESP+VUw0JpKrnNLNz62cknSfpzHwN
+IOnl+aPe1Qctg1+pDbg34hARL9SdOgMx1pJYn5TvCj56lMHkpKljRqjcOMuxa24
Hb+SHP5sIPxJuChoRUe82DZtR+nmwNV6Q1qoqbuKHttuOZ2x2/L8xB7k1jGKQg5T
z7wgOZDdeIaHQG+DHDjB2UTimyiYyFoDozOsGh/UYkvSrrT6cXtS8DetY3Bc/M8s
FH7mMBstYCk8MbfaK0MyjVztFU5Nh7usrHSVN8KZzSqMWEvRo00+eKPPLKYoFjPh
uJcaAuilhdpo0UQHywjPHw/Krh1jsVIAcr1blyQW2OlS+zgF/QeNyMYt74q7wYEH
QJdYF0kxIqSj9hSbI0NcvM+CaYIjUmXY83dN0GcMvWvbkCaD1gUqroxwSglkZYX7
tQqb7I1fRbHkIR3miToLb+RExsKoGMbXivWEIM5vHtjsVugnw3pTvNowbNYuPPub
6zK4cdeJqRLFD0clf02O0w/glA+Pt2FhLDEi9mXFPrC8NFdz5B79+8vEe0Xajzyh
N3Y+Ayc92SAmYtD+S9URskG74yGxALe7gte/n6cq/g0MN03sXU7RcXTJQ4Uj4Q7V
YxUNHQsjJ1hvM/yaB/JOpa6xzAiit+C8plWyXFm59lPbNgP1OwEhJH5vHvYdYFlt
rSBWW8CD4QW7yP8TZ+EGcG4nG05LSJfKmfpbM4hl3Y5EYUxT5LxvE39vfdG8pvyZ
I1uKwdbCHvANw+JB+F1nHdy22DjDLWLcEkuFbI1YSpBqVQVm2BiJjxQkc0f1TvXP
WeCC4HjNnnRf+PMl5Ynjz5K0tNhOGULH7/A71qscLJkXsShuRS5DpzikoPbEfx5S
RyWs8UYfznnd2WKKjx7/Yd2RAu9NEhNOSPaPPbY7LnMu3gBpJCFLyLyg8fAgPZAW
fUwTtDegvooO0jXM2Jy4i66Fmi7Yzk+dKr2KvfTlsqpviIUJAfeZKw1t0cXSvOCd
RrOSgismWBgTVtpRkkIBWGk/rQXJRZRruRN5HQeGWb/BQLOiggqzM5Xetr9xiuni
1eSlUBCowxwa88TQOcSsTeCrG30NhRmK+pj91wp3sNvJqqpnCJnp3i9WzMEXKg/m
NgQgg9ekJUqF3Z8fQbfP+RmsIHhyYvSqmIQeUjqR26oMyrOszQV/bJDGViBpyGyv
N7/QiJVLsPH56d+9C7E5CZW7/QiXsEVu9WowW/pKzw7Pg1F74p9B29OfdhDXaE+5
adzDbU/oOr4ixWl0B2FFioOeynibwPbFMJebaJLzkakOreH6OGi5zGsthCfR98y9
kwjjNcHHdVYxF6BxFFMCwry93IYLnDqBdcvcqHmQxaTvZJPiNYNmktLyv9DHirXN
wkyQj38XCvrdEFAhMTiPhuDUlxNS90NhXOlM7zEK0h3PnNR5L54ojqOoTHTHniZW
6aT5Md0clm4JFpRK/1gtvMmRVY2pLIlevCFM8rLoD/66UK+fSAc6e7amYMfQ08/2
s2elZMxQo4HEc8nrdLbBamlz2LHxKPmpMgBRc0MZwGJ0DjB/4gYwaUrBVoithqbK
D6WDUX56B85Ze9lhydNZ7elo4OpwlPfyPas3hZUr6nI4IizNu0wl/+9JyqCm5c2T
LCMi2R+uvPJalYA8yZFtO7HeftdloSMh+tqf4RE3P2vbCb13wvqUe4EAPyzdzJj0
Fm8MGMYWeC8hXice/dcviitGxBaA7h5DL27VOjPAhALy1mshNbZm66sdteHrw62/
uMA4fXKW/l7T7wpcicWlcaFXS26Ljh7Jsp2Wu5T2M5NEsfqhrWkwlursuYGvuvex
1c6cif0b+zxcemv7E0v0IYc7NBpfkO0o1XLS5qtQ6X9OpSKre5qLyZiBPIAUFI4M
bPaTXjiGCt7ixs969lctVqv/pDbQ8GUDVsk+uAzEctkv2u27OZS7xffDYmLBW0Ae
AtNST8yzEl9R9NXLhh3eN6UaDj56Z2EphHD0zOZFDGYTt7T1aEjJws0gGj5g0ovh
vo9VZbU50hkMuWwR77/MsGNEnevbZThdYhxDG5oNoXLIc2Bi+V0GcetY93w+Rkqu
3nm2hBwTeJ/Lu7ZqnOZTcCWXCLlMThS4Gs2kjfRjUvTwEcRlvp+hLuafooan33j/
wPwmUzJuwqG94rGNv/OlXEOXI0/LHKg2WQTBa2abYT3+RBHK+DOHv5BxfqA54apd
JbrX2XXECnCzn5rbhI1WTXyPJ4iwjQxE9mQw6H0WQi81HbHjTP9eA2454tZcrdh9
8/la4kG6d5FVWBg5e5D70D24EPeFJje8GOR00JRF7Ef0b5tFR492sD6yWomdg54w
uainthLE13SWKcmuj/sTJMyapdQwqCcAuJb8hpeIc0qyKs5gWG8kQ0n/nBio/+qp
fHV6kQvX/pudIQ7aTnRutn4p03G7e2lbuPYLjg4oW5gknsAVjMIL+TXC2huEiBs7
tun98nt84FvKCQOIQBjatq6x7RUJu93N7nzp5eMQofi/tip08H7B/FQmYh2K7IRa
dEu0p7KoORsGFXreX+Tgyu/5vk5t08B4WR05G926feekhfKtr4RqsS69W/HPnfl5
zIflZYnMuavgqIt1DXTu+WVsLcJSTgBhcsEugegwTwh8RZgronUo0TyDstIjlMnJ
4d/l4wnlqdNE08SvPgZsxffnwU9Y04ANM/KanchBUxX7SR4jmFlDuI94u1yflo2M
Wmsnw7M543EGCTRURsIMzMLFfO1FdzstRMW8vlRpiafA+2ix7SO3D8198EzNOUzD
vLKTdc1n6bRvYXElurMOM6eTGuBJVuwZbptE88YqlLdla10Kf3ImaLrvFI5tNKqh
Npoy070XBbA+brtCnnKN5rJ5gfZJurcwuhxu2/RcQni3rSY7cR+YJa2MTddBRYyU
bJcsIEiV78JduwYaLLOpq9KOglH+WkyyHVAW1y48guX93h+x4CGi26BuJI1GCMkx
t2K2DwGeoXI+AMesfgC07p+gIpGg0RJ5M+6u1WHffXXR4bexyxIjLgzKjYilUwzv
Q3s5xNh8ss2zLCLl7fhRX0OUWrl/hTmH44Nx/OL3aKo+32RbsujNG/qMBskURc2R
sfuAq6bLln5PMZIs/8WLP52wlk4eeLz9TdfkreJXFlQvzF6IcL8cIo9GN4P013cb
/yY09qVgYNtY6h0bQT/7wPqkPh4aC2r8Sa16Rft6t1ZKvEH8riRMhBjwEb0C0IVL
U9fMGuOXuBuewYpbXpAnsP0J9JSjkhXbTgGQWlwiytn/kj9+UyLWohPVS96ICtrt
aInj62CyIFemHTGQ1R9uop42DHcwH8Df3kj/bt3iACReGYpjHhzKtaKW2m8C+aTk
3ZhnrxbRSGsQiIKfITZTDjge64jscPxAEab3mKkBRdVwB2qmP2a7lMnJeNjtt2vP
2mMumbQgaAF+wNVdi8WrmZWFZc65fJ3oxux6qAA5O7jkzplr8X18G71bSeCcd4xl
o24RNHrSOToCmgNYmByvAkjiK+UyyEPmLfkiVbiY/KsW3gNwBBDnPSh9EaDkR2yY
EWwdzDUuJRrEcXl286z3/qP82NniZKOqeos1A7pmjL8QFnlhsEDvduzqypU2SdZh
EyXgPUGr3jno2bxkJ7jNug4Sk9CVyuo7YtfgCIvPK9Rl2iPiKgzR7L3AyFmC6i5w
1C0O35IgN2bKHJKfRZAznS8xrxPJhFosCRNKMn7B0o0chjAc817NEnAdlYe+Z1W0
7ZWaPaU8Ja4cpm8w8xhAKku7b9KZEwSvsTK2jiT/lrGJ32is/R3XU+g/MebruIZC
83LLNxBs79M9njhQM7A84zZ3kyRV2tTZUIOF4DUQnUPET4bvtKSDtEapfeOg8v2x
+fR2IyChhH7un0gPXM7s14isLG3QwDrYYwxvzylmoUCQrNu+9LJdO6KI+n1lgaxL
gfT4YMYmjJi7h8T6P7O4WcRT5Qu7emZ1FC/1OR3oEHi1EnKU/+ott+P4j2SFAqRH
NZjQ4xJ4WwUR1VEbbU1WSQWUtRQo9ezPxwq8XuruymP6RPu8RaPGJkWVm1kA92Ax
9bClHuan1abUGA13MdLuKq1esRRUZacKHJHfJdIefbh1WidkaSVpW4GdZZWjaBrw
frMSEXo2Ob2pCtaDB6x+AWaLZtjirIiLY47SmzIs1KGd6zESIlR6wDTAzG3e8K8z
OMazSK86KZWPsn/2RPdGEtPyOjwicLbiRZFcgJc3P/h6Du5ljfwPwu8/KVlx7quB
SX9NP2OltfyJ1JU9NMoi8ZjcIRHLBeFZgrMtieSccm/1D+y+5fOYkS4scAiOJUDc
M4L0x/65Rr+zamg0bzXd3I8SZc26Z8+nUJFohJxrfFWEWuOfGCnPVBNjLygbyYtX
aexnqrmglYZfspEm59PRkFSf+DQhXqhjGi5GH0rsUwM+kR04Ag75aYZdLLiRxHvH
7OjD3b2NpuYkX4/YHqm4O0T1CmaeQ+eyr9Jow4bs9Vs4+DaHvA/yuJiWu+Aoplo3
0ZhWRmWhBd8oiROfEKGrYkRddxdILURXuK8Vz/5SJxBZtiyfrbdc+5y0l3q0YDvK
LbRpEds5TmO90k+JykVJMlySOhaE3l/vWz/4pqMN3HdE8TshyAkvuRCPEjoTNtwS
vKAnWdf+GZNdSkT9TCeNHH9IWLa9KqX+OzTqujApAhoQ+7Fzs5zP1+G02sHntyGN
G0lvk7SZatvBCHL4fQghV8rpiAHYIo7mdfVkuqmvbElVO/A6Ztf6WNtNpkChpZoc
FgoKu663Lu8Q+i6OQatOsECPIHGzCl+t51L4caZlZycIa0YVMUjuhtxVLgGnl4nW
pU8KHrGAaaild+i7yXnTFECLmPvsoqp5kT1oBdGBmnMy6PYfJ4fQquy180r2D6A6
6/tmLqeFoi4wuv3SCFPkWNXn0K9R5GNPnzlqrG316HczluIC89am0P3xZtt9nxDn
xSwESswDbkHwjfSomhqzdz9KqWac03T3NDv3Mev8IhYLiE3bcL3kKybOQrtESPJO
T9AgGb6SrpVgD5z/LB/xUWCxZ1y4VIzTuqQYV8wlJrdKZEcir7VOua9qZs11HaD0
1H2gEhSvCU1N9hjDSU8Z8Dx77pRXdKU0lHZPJlGT5f+CINYX/5Ce7uq5esMaIxLj
h7vMraMJn7iRMV1XSekEgQkW5IqtDVk8yfUDNqyJGCGIJICXitA7jQ8iBLPWZEhr
ZgX8MbruF6+LzyVMuSEUJVl1M44TzTuw5VEiuZTtlz/ra2RwYrb+iowb4l3tij6Y
twWStlYpm/d2VKmxMNQKEmSm7pOl2fYe8CDhBt4ur/VLdILMymuQq8Ydn94suFDK
PXvwIaEuZKQBihpIS0jM4dWN8601zjU70XA5RIkWAX6z79WvnJNpy9594zJPUVUO
Q/gutL47cqZPnOBelSDUFsc8IKQgjSjTmHtPalD3IkhMnWKnnnluWROPQ4yg8pKD
U/qhVDtab3cox+8rA125paN9f3UbfoGB4SROHqPjRRSVaSx5iQsoCdrtWF6Em+k4
RBs/k1ZqKG8CHFoRoEFS55qC6MZgV7jFKyRznZKycfFw3t7w1w8KNuMO3d+gUw4a
q0JtyOUxIKp69xF0ObmkmFD5gYXURMQhIyfLIH2w3laaYvV06Hu1v015fjYA5Du6
k1/4SXWI5Y6JXBBhpye40H6HiZRNdmszcPhLf4vOWq37xRFa2s/Ssd/54/mY3/l6
xr7+OhFTtzeTLrsXMV/PoecZW3nIw7US5b9gyUarVsKINRKyp5w6ViR89TpXAOyH
1mygEJzet39wV3iIwSloUXi1kRbndCKNkoitIWz02YYJa0kp+ygFL9oZMjbK0Ysu
JmCGnwzU1Hbspn+jFCuFqCIcP3z/uJRfHsDQrtCN6k6esP7SRbG+0E8W2wFLWY5g
RpZUidmLhyjdJNipnl1oszX9T5G4uU5YFkqQRm+mdEGxLkcLxX8+Gu9O2HWtg1y5
lVASltwyqamEJklB5k57gM8JKxZBpG/DRUn/xFbvUBjOQnvvT+Gbxm/g9AEu4W1r
YULateK0p5FTRakj7H2/t4y9opuDHclJKV873tKkS7C4uJXw7ElLpnHqCGo7zWLh
S4CRv45rFRhAr3b9JEYi6bVG958KRCI0yjZYaXc9kuyyGL962dhdOX5JzfWzQjii
b5MmUqLMNM/01ZEGve67/UBdHQEJ9M6G9iNprETCOdyBUhIr7iYdOMLJ55vDJLsw
DfNOHCsfQp51oesuCO5oe7qAQZ+dHwZqRAJJI+IHNX03XIOCMOAnxzrvioroQ3nt
GtZaSztq2P1Bk6M7Y/PCUGZxJBLrdHPLoSwLZs3v+LgkZ2XzJaonQjHdmdK5I8CP
5j7cdyfwudYzkvnxbNN9nNKbVWXVIq9sv87bhCxpeqE4wdNn8tADsdhaC5lPVotK
iCtwvDhgPz1ieVybjMizyMlzGC5DXj9Knjotu4Gcg8N11T7FvXLALWDxhgwShsAz
6MoWlfV9lFDRv35XxuXKEG88TjUtB9Xh7nhEuHwRfbX5G8JS/t78D1vTsHueTfru
Rz7lAU03knrYT6Hta00/+QaaY0zMLHO5l5jZ3ALrLqlidoXf0GvjlY8i0O/Exsf7
afLFFyqV0e6uxzgJDocTZK5RefqD2cPNL+rqcOnEq86rmqtrNVQwGktfoIWcOr2E
Qk6vn0FOMB0Cd2erqLhpk8K/3WQ8TkgDmw6wMXuAQx27Fhzq8FWnR7WqH3j0UC5H
OdKvh1Sg8/K/N1lFDbIjXEQMfJ3hB0u/hPsszS+Nz7Zn7IeFHrlOFdEWt+Pc8H1F
8CQP7fy/3b5fGQ7an50pHZFms+f0idbKBIUPRP2GAV9JrbQyVi69hwgE01bavlth
6taErhIgJAwJmbngIrBOlkmIznOXhOpqNUALdsFLJtlb+zFmGxtKeKPdlFIY5a06
4vH/wW0W/L3Hvyq8Leirdda50KJ2czU2aaMems5L9mMMbqWHtD3gerezNELE8lyR
D1yUT5kg5K3DchE4KR6XjXahLBOM6nKm937mnO0+k335CXGLQRUdAAYdVDsEOaXF
lVc+jLFy+QSZm6gqs04pjJgwtdDcZMZEHPsr2lTbSRw5zqpfNILVJ6KoY0X5zLk5
i8BhqFnb5zS4RYgDlgSd3QbzY0ZWJp6n3l0foxC/GROt1EezhhHwHaEwev4bRHYr
KF7/cj5VWhJNYDQsT+nzHHHnO4z8DwtoiMBeIq8wtpZ1Pydq8FoiC6OhrvCjf+mn
bpIRiTSm3kezfmHnop6J2QDPfc3qQtbY6S62XFU+mil2hXYyRkHS21o/ZR8Avyih
do1pJ/iHc2pswO0R17XEpf+Q2vsSi3PRH/TocNSwrpzWNylzATliOYEJSg4Jn43w
CNtQcIRcX02p2wS/1iV5NYWwdTLfCyEOJ+qbqyDTHD2zZ3EyJtevlpY3G1/7cuSs
jBmIQfljI+jYJW3SzZLrovw8QKauhqzRdKpMIMwPx+m64yDzR7y5w3qDGeUwz3L3
7cAM2UMFTGo6FiEkXhEZWxYNJOnBq46On821/dreayz8UuGPEIcZbwft/GpeUPrX
1WjGTmxiD2gF9RViDUqD+TxQtFX3BOCIkWABJ5Sb1GiE8FmTMJiUJpId4kapPp6m
Yt0/Si2Ijcl6FsDE/deweCwB4Cnuo/AgAyW/v9XnwaA+DW0RXELX/g4fcVTh9rwJ
xPkY3isf+bFnv2mU4GMtBFvSXTvOgY+HpxYGz9ZMS13WIwV5Wo4le1qZIHKQrhMX
ZO+HXqqFU4we1mI/kF5d/Ik+8IeNn93oLhjNj72RfT4FrcW5roVySx0skiZDqQFQ
387hwewgUFyhUHrbWO7g6jyz9wQDlmysC9ikMteeArLCcf8oAfqkWxtdF5fEfX74
nqHlLuTtWNOsjheAQWOz5rRb1eiO8ZbSEMvKHFx0rcuDShjuEYHmncY1XCdbJqPa
I/ayCNpr5wbx+tWNCm9VX7xdjFx3v76IH4TXWOMmPw3J/bCbQgDC9vJiJQrErtAm
7yLGZTfKZmidviBcpXytSo3sYAHa36xIfjIIGM6zv2Onsob7Rx3Uc4qQOZ2wwMzO
J++OBgeIbF7lwuUSEYx4iWp9MwxopbOzkjcbQSpW94Wj4dT68RTwC/BgiyPOQkcK
j2tRUgmYz/Y/f4UNefsrbAPIYHF1t296LTIEjV926geLzvPgt+kApaf6qFa3hgg+
w+80LHtChUcZEcOWucgWGM44ATvFk2PlLI/OjVpY+ZwlYs3A6hD0vBNS7IJYwj1J
Etff1xX87B8bAdBStRGn+VxP3qNKo348jqjo+z4DM5vfMTvfhVf3WVGL2kqXKqJy
ibCeDpL+7IMd3Azk1zGPBCO3m3Mk9vyeKExzzX8YIKgeskGYe7nTgY9rZewTmWMg
dpVKeDM4sKJTMM0mll2/p4nxs8guiXTvkeQzQLMUd+a2JX/HfB1Du55AQfquBFiE
D9FnfzSIxzywvFHx86TBHlwTGG0x6VoIAv6A49zc/KU6oD+iAOLV9fj5QG//lHFJ
J1LI0cNGfe7Jm4bnzMZ2riZc3KdfQBw4++BiXBLJ2rtolPZjqNhy//VATL7iPrbu
kRh62KSkNWc73I2bM1kXVTAw9IHw5an5kYlmgk/Rm0A/1fAdMM6L7zxKVie3VfM6
6TN9CVT/aUgYtMFEz4jGHZ86RclEcGHG1oXN6e1UqSq3Hjy5KG7NNJgVFDO/tmPx
P2kEsoNkUEuTsw34JbDaq3hDsTANCrTcziBj2CP0WjE8q47eUAl8OZbKbCHqRPVh
2cFyFVgJsE+yTQMPgyZA2d76scBqThUn30+0PgsaA9ffKpXU+qI140eCIPMB1uZV
7INPZxznsFUhTx58B2pIDHKD3WBadyFG9M8yom3l/dPsc+Y9h/tNYdCECi+LcTcG
u9n4SXQcH+Mc/Gwsb/Y4/9UsHq1Vp9ls4bxg2et3Pv4LZ5n424BuwsKMkpmcBrDb
HiAW9tkYBJu7/87EehaNAtIVyekH2BLw5204i5nDKpFiwUei8LqhSo5Gj9qnOQZ9
TB2WI2rTqhoyLfMDox8pYWoedXm1oYseZ5rQip5yT4zZdGHjmsRAG4Ab5nm5xhiZ
6BeWfbdv3Rr9eC7O/x9bRJvNGpUgcMx7o05ee8359CxCaassdEaOQLFs11bOKAsP
KBo+D9VX/PBh3Mc0SjBOAcowbT4V4Rg3vZRXOwHeo5TQ0nySufrtLFWLQGSMrtTF
lArilO9c+wU3lyh0L8fgZvoHXTtr9HSEHW4AVLxHGROem6iKtzOlytjtLMbF+6Rj
PX6Xw9vlo3WhVlbHO8zhtPKqzSjDWI6W3xaB9NUulHtjmXvQPmgsPUF+Vl8C9UUU
BmDM+WiGXx9a5+BY0YmAFaTk6Bv2LcL+B/d6J3qHWiGfAP95RVyW0ZIo8Ftnzh4B
27Y2mR/O3OpbF86J0RxOuSFxM1tAJpCG23C57+UbJw/BRpnETRY15MA1MK1oG/Js
WfB1THyYEQG30kpfUfcKbp4NG4f/J8CZtOBD65qUlK7M70BiQdjL/FGe/HIezuUj
uQqnFuw5gea12M5WLKj+tPvbOI2alszpCA6qMP8dHUdhRVP+Vk0v0kq1eqbwuscw
ViFlNjBI4j6aExN5afHdl7uO3rlsoGCpBJjjWibKO4lPVNhW2C1JhmjYeJOk1HzW
MonI8i0ED2tqDUK5eIq7jNg4+Bki5ERIGc2x3Ym6Uyx4RiynsdNpuR2q2Li8lPSn
KVhcN5MUxdmZNMD7DbjnbM9g1+W54y3n7w1UxbjuDRVS9A7F3GwaVObiM+uXWISO
r9uhMKCzwIPDhkNNoJVhWgcJQe35qehcdTwChD1b5iV8KO/hng+PUJO2A9lnj/FH
Hs9HJo6gepCbx6GEXRalsnaKFerg4EzstbbZNo+QLSLzTjkeTxRpbTODqkkVoO7U
MSXdppesbYziGiK5emTXQFbZco0IGJ3Ocj3Am6LvRmpiBKUvR+b0LDRl1wj8pGOY
VGjaNwwd+7+IkrbXRfD7psiKPi+Ijx0ZeCcVu/R3X01ow4eHLGNXcQeSu5Sk2dWl
ZfjxLLahd22QJfrgQHs27omwLOrWG1q/b0xsvtOcZnSU+1cz1f14ElWp2JTohTWX
LdjRFbWuPoqxphgyJ8a1wnrdh/FmSUf5jjmKeIXNWm7f8mvvURmgHHlSS0xB03y2
Coq/AabDZGwC5cXL88CFmINT1KBlMhnOQZuRgYqF3C3HfYv2mv+CyiBQ9LThQF/A
A6ZZY1o4Hf/iPA9teGG4/wPP47DcYXq9sTGsKtDwC3wmTLC9RtEbRkAsDPGfoXcp
aHhle+Y/hQEcR3mn2tnkAv+8O2Y4/ctMXhnPP8IXmkHucMQfAXfXvZQnHF3jm1om
P4HKX6EOw8rRnkuaomV3Rk2Ia588nCVyBgLfm7RX3GOH05LAT+w1cPa/b6Mfdhjx
sN1W8eN8qulT8fESo0mvhauiCEiizK54WDsCFm+S1Ms9E+s81HyGCm+q/sreOFZd
rKXaV6eoRt/sZb/MKq/O9/+veWCbylaWE78h4vRJHy33Dlgr0Eoxs27L9G2X4bDU
2yawBatUdVB5J0EZ/tkx1c+kBB5gbwmbUDXxWlVTkRXSKn3VORiOsraKm/w/Zxg/
crdivqj333embHmIuRdW8gt5Tf6uzKalCxMil+8OaEOhn6SzZHH7FYKpmWDYu8ut
vIm7/7nUNWPqQGY4oRY+Bcz7EZqOdgvEoj/RSA8NzwnYMy8mLa+H4SK3ZhoFGIqR
LLfk4PFoJJu7OHFc18xiSNbl2T+HsDa9XiBKqNlI6Yn+0/akrqqjSYvWHizBb7yS
AGzDv+iEnZDITqFX1Yn0EQwMQp6CSqVz1E7tvtzGG3CZu0b7uuPKAmbtq1xqMXGl
69/BCbMcBAcF6aphH2XIKLhTLccccyADtSxigF8Qbqsfn9TGnBGQscbqwpmDGXLF
CSUJHEWhT6mASeT0pcOHwi3yg70FrT8JGVCUqX31PbNguQ0BOyPEHgpFd4EXNyaC
1vOGYyCQrKiPjNFeUUs9zvsVfi/fs+ngdHsoncf2eP8gchBWyU6q9HfoGfak51T3
0eZyA5F7//7Ucf4INq3vC6cru7n43Xkaan78yhTTVevsE7TasIn9E2gHjPuJ8ci0
7+LytpFdfBtc5tXunTfLLaBf4039Mk/z8THPAZAXxEXZbqKaVFATJ0tV21p/ABlF
3pEJvHr99d8b2J6Nxf3kGEG7BI4QR2/A5gKPoxJKBqhk0T3tpnCfUFHsL2+85+QE
xBYnykhxdwoNQwnvJMf3T37r8c55xIZwht1WA7VREAoQQhlTJj0aIPY/MTi3FJ5/
boJnGYkzoWgUF6lZ5t4tUL04RJ8hr9NgN0PGYu38UkydexgwzCNWQDNDlREjZkXz
GApz9uUAZR6KeFWitCIEkEjuvw05SQo5UqhT6IXylgx0/NpBFAteBl+89j/h3/1c
tojFqAAtOeakoLmdDpLeg3RwrHiwGwLC7N0XEwXCikm27bV7qtbFqtvwbUF6xhzE
ve2vJUq/XIE4B0yIHRYPohcL0f8PApSJN68Q83HVoU2OY7YDOAiNqMRth6esqm1h
XUdrS9/SW9D/pQb9bMAxywqm8U3JKNocGr+lvmPjvK9lC/UZ5M31qVS9bgfoub2U
ovdGV0UZD5OLX9VtzIT6GbUhyyWqkN3KGBKqvY53cVT+YS/VJouBo9EoyNie02BV
U8Qc2XK7s9zQrgWxIBj7WQDFb6pAUJO7htBhDMZi2idBepHNkIpZAQXO90IxlSvD
u3oYUSnRaCOnz5+KdYNwaFYTi9nzzs9NSOgC07CERZhb8v2ZQ6Mw8xCAVhX8SnLv
Rkl83W/K5cr4T6EYU6QzyMq5mqePBDzAzPzLEBfOHkWCetyBgkFxs3iye1beGduo
/Vzura+iwFO2WLDagE5+1Rz+e87U+SPNsH7ABTumrjSaJxwASwrF9bGYekEtzXb4
9F+TWIGdOXqlhhNk6tvDsyBEVngJRTSvzEYTMIG/zjylT+Y0l3U6ZAcwE4/D0cGh
scJmrPNvVMhgSCsTm6tm4ItUExwnf4UuUBxBy28emHQ69HpxOqWdZCcwieBCOpJQ
94hOJDSqptNP1MDoczk2z2cOu8UeUjZpGxi8eSupzQnr4hKC869v/HkxS0DhkA+0
1qCMn/KWMASrkucVZT9OAlxmN2TMdqXwtXt0anxt1++l/MW/NNPJH5tqfIEyTKep
dPW4ItZTL6X8J8qW9G2Ag8E4ofWNnCds6wnzKx3nhOerTy4gpingJruTiLcGqarV
e2eS/ux3plIaJ4bC90vyL1MfEZMJJdIFrR0le3ZrZhk0P4sWsQIcVo8ekJbu1Zqe
/T+JY9Bx1ie3OQQOD0mjxM2F+L6lgsNAnq4g1vvC2LKvhJSf6Lg5usIM0dfU/P2d
CETg15rElbZiOX/G2V/bHFWRMiKpGJ/d6kdxnU0/dqRkAy3tvjegMG0Wu7Bf9A6K
6byu1f4twh+LVV5MMw9VHCZj3vR6r1tX5mJqZ13oT8qlwllxYW0MLo7stYetH+rH
bE/1tnRujCtuk5aPVvJL2s3nlIrNdzcNkTqx5YTq/p1EIVEz7mwCNIbM4FSH8QYj
BOEzwojXW/0WUZ7M3+QnTgHxXBBImDX2ZZxha7hLliK41vNPStOCllqcFpelj+6o
/elA2qxBdASngGyt1npi5DxXIBGdU1xKd/ezHzoQeTYxt8/vKXvCdxE4/EYDAtD0
gvp9071nSyRaZ+1LsqWJ1NJft13w8gb9a0++zpJ4w6KKPYgH9Ndyip5Q0KMOMs51
hQvYcQnhbI6i8hHRsTzT8kPN1Hx5vStI96mhlE/2dE7qyCgd8uWpz6axjNjHIuNu
SC5kCvx8O94mn51QOt7G9WKzOeHYGX1NMH2bLcSrZ9GTQqsRXLk1i+o8NZLOcwIW
fhg8Uwkefy9vLFZPLokBjDCqbUyFpyS74ShvygUlv4WImmGNJdCmFxxcizeOght+
fhAWEGp71d4L+RDzaqqGuxXZ7XnlEVIegb99yaSQwOtWZHnzo5bVqhKZuqvF1jk8
fgTd+sLb6HEhi1LeZzgnRx5xLui3aEsDZbhrvvTmq7OmIQ45Xe0HbONuHh4OTkCI
Z8obDa2RhlwLlrRXvgGzgR+60+6IqPZGLGa8zj529Ez0et2fSyhoAhtWy1uEk9sf
JFGjonJa7Kohyra8ZnPaS1t0+g7UH+S1wkVTmmIkYDRB8eTP1zjCNLjlOxfEehRR
qm9uatCV2GYkeGfOzec+NOyZQkHxDPqpzCQgM121Fkh83yqy35x0MFLCSNsmvNHX
tDD1gSPRYdVTAhvLTgK9njSjCEeKo0vzjn1Xgg6ENf6BqgBJmA4s0ldG/d2sWJuJ
aIamZ/PBV9Rh/TiMuX6dxIbjYLgV4KAQMsXGLToYV1J6pAkQtqfwUQMDWEFD+Eq5
Ba0RCDFoe3u79ZEwLGflZcrwTh4CNORWRaPbhnHzjL47gmbqFMCZpbfrNcaMgmyN
jYKS6fCitJh9P5ApeS5u4ALt5m7oj9c860/5GNxxZ4A1yjT+mR1EFhnyqMJ+4Dr9
idrS/TwYVwhCEdAqHZN6hF342LU7OoOuPKxSjLF1M2tBhMDT0wRuqWQtaSigfc9l
ZgRqrhIRz4OjvEtgUI1yDw+EKJsqxMTgIfN1vhSTAtQ4zzWRHx7Y2KHmKvMgfLj9
+522SmzsLdc/oxO4LrnP7nZKQI2ssHeP9qS/ItI7ytvMmjdcFDOMYteM7ymp3OiS
bCDOnqkn0RJ3GYQ8d2Zk649QRHq7OxwOheAZlEQ/5819Iy0xfS4gr/wDjiLX5Acx
yYpKsmPiqSD9Bk/+hVHBFMskuzG72Kh295birXgTzZrNdmhhZPvWolsHz4z3j1dQ
eD7fPayhbEh2et3dLra4ZmdMelhFsNt/TuHIQcuZzLwuA3PhZ8JUd8WDlCRgDzpP
9AwzIQQzGMDciEvdXmUR7XQ0KqPkAcvCmpsJXoSqQLr2iodH6p2I/zjbpB5oGOco
d9LAc3hpuapqn0VDWZoMUchl3ub4j02+GLJ6geKFpzOEJoczmVzV6kVs6p0YdBU0
E2fj9Chw4phnzrXgCG9tG0hdor9ehpFel0xtdJsJIGk8MhOvDSY5QAP3K9Iwf0oG
5MNQqudIY1F61QBvY1SLrV/QYIUeMs2YIQpxL+mMZSg3a+YAVvGGgUM+daBumqva
0SpsufiqFD/hSFX0KYh35E8sDukEmB1oqH4iFnSjYKYCYOIPSuJowsERObQnLO2f
AoUJyN/C67+yKfFJocHNyeefxOFpyl2xnrkBMy8mP/3DbfJDM2OXNNo+zpUaTRvy
mhY0fQcNfqMBmsSoygHlsAP0UoFyhviFTT8iValEiu/X9o+R7N9daDZ3rK7JwgQT
ZrwDjyNZWMcTDanz5vhtT+raAIEdxpPIhp17nMbodWQhEOmbDFMetvLtT20C5Q/g
v+yis7bQfpdF27XQg+f7MWpAQQzBLSzsv0oEYqNqe/wk59bXNh4uMzUx6gtEPrsh
yQVDLYhD/E1yuwZnmRK+u612Uy4J/2UEp5y6aYoAwQonMiwsmwophlIdc6zZc1FS
WvG0ul77q3B73A1izgP3+guOZJieLB5aK5alDoywhp1Yqv9KdPTHszJmZx0jzDu/
VDFgpAZZmNR3+lhS3AXzjGbkgLbyvc/OBFDrYUPq2PeyR72JHTMNSf29ZlqglEpM
xe61fSvSVCCi1HRALucB8MUrfV+AMnSOMSTypdDkblk5mtKOCpPg82E/qZ5mSfbn
ULPdblEXdgpxelBg2NvT7VXVj+AJnEg+XlnRbGK5MOBARAJMOHV+RAtYS4c9vgM5
mIt4uzb/m7TiYD+E0MtM+Q9j7sLZOWaBa7uj0jfFoJd13S+Qcy8zz+USh9X+7ey6
WNJNuCpt8T1eBnv99O+EUOWVBoc3PQHsQh+izJrg0Ry9dUiKu8cVUwHA4tJ7PP80
k3ymx3PkNFt7petKM9Ffz5ZU1ENTeWCKu0uCFsStrtTdH7hFQ0wnWKgma0bO4lZn
fZIaSTh6ryzTy2aS5LXrULkDtqRbqR1f288rXejsQF5Iy8hemP84DVRKcfRc3pzC
G9h88wPd6B+euxv8cuPy0UgLwoh2Alht9lAwErwxHF9lwpJnA2MJ9jq7PtWt4hCd
Dg0lbQBokoqy96+r3dkpQm+BToT74zrkcfq7a2LNgtaSh1/NjM2jbwTta3XvD8ng
jov7FH1dkZu5/AmQP5+LB/8VqtSPzjezo3BUp+83l1wxGgg7Ej3XsvW6g/j88T+A
FIWNusiW/Ng0qwx3ashFDW9e7aKmQ2+JxgHq5MGD/YOS4YXZQCPt9VheXhGIti0p
0FaklTQV5vUsXSODlda1r6gdLtAcv91NMWePLOXcl3I6GTMmc5WnkZrpVJfCGD3Z
JRY4b7MFd1/bKAwFXh7Vht17fyJb93Xi9ATZFzfKnRFOFcIEczWka0zBHn3/jnrV
roR/tCOUC8ufOvDpw+2Y95VZqc1U6sBd98KN8dvWkJcjVdltyvIPPb9XIY7np9qr
mnOQkAxoUFTmLx1ELDqPR6+bxbzvUKruddHcwxCFuJfZRDt51XbP3KfITOybz3Sl
lJWbbhUcQGhhWt6hBo4kT1CoJCRXJn0YkgP8WAZISaIHN/kGGUq2n6vdA0eFJ3QZ
KASyVP7iWWq9Te+Rpsq6kMUEEZo8r/Wct+iX5vKEzPF0t1UAF04zJwal6JIy4v3y
H1OzX0Gqo68YoAk3Z9ZmkZJF8PubvOJblsk56wJHMVPiO9v5M+hBqH2SWtX4yT4e
q0Q+v8nb00FUKO1XqIn/Ejx1sfToJwJOBNksFEFdqZ8hLMxYH0q+ZDoraXyig2qX
7BBa3pjxgS8dGgLPrSzNnSeRaJ47IUXnaK6aLIGxn1wags6tQLHWgNV3WLrjZASj
d+H/Vb7BnOaz20vqIT1s+arggPi3n6CI1V2/xeXnRmWZeHJ/bogJ+XshgNxLm4s2
9j4EaOdXUZJyd2CT5IJAaRhhlsw0Q5tst4PfHgGhbNsMUGZewSSchY8GJ5us1waO
AMz4tMtsNAFpM9RVV6/o5cKInEIIGjM1C3xXKL/KNIdeb5H0MMnPoaHwXBcN3RQY
uVIg6prw5qhO7EEm7G5w+Xyt7NHEyY5oW3WvEF3SMbGXdj3UCDs6cRG1VtvVdNyJ
JCyHe/s+IQ6aFOWF3KonEltRJn8BBR5k7wu/qc0/lWhFCuR4+IRHxz1bPlV9Yb+e
1qZRw6cikLAAlqLV48e21Y9wFMSygjC06QakLLveMsUBPG+nJH2AZ5PBnB/ztzm6
Lfhke6KKbHihAkXj5VWFnKct7Jqvxbd/dfTBUwWWD7H3COWAvglmBznNhm69NfBW
FofrVXrQ3UeQ7+2hwv5Dn9bnDyigvMXPdiqBe4MWQsbvIIAM7SPgK+1YOfyZOz0f
pdKeyVho74I0lQ3RKrklhnjTfaZ31lxF8dZeD9p2/OUZKarcP8glZsloYhzGPTvw
9OtqwPPEu66l3JYRUt5J91H8mnlzHgIvkjBuc9lSdyeOynKOCqliJ6uISquce9y5
h7jSVtztzQIGHO4yZA2ZotYJnihWEWPf6Xo2x8WR/fiFgdz3z3e1qvz1Ve7VOZ18
1YNl5VbEkP7GiSLN9kTz3sI+/3X+r+fhuaGPhoi7zOPjTKgddA3oPep7QjPaYFGr
YlONxEMFWnTFcTCCfGTHkfVaj+VTGXJWG90y6gG0LdV56XvPyauSWXVjCD1FZLTp
WGgB9HJZdX7C1Wv6UEm58NOdFjjhZ6URTS/MJse61yIkMsKV27CSzpn+a6+XruLO
fVsp3dWxCYp83DWlH3Oe+4cFtB3Bxr1eJTdkmZQg0OMEi+gh1w/y2CGogBKY9WUh
Q/AGjZA+ItIK8GM3lgXevb+tXpYUjWGldUIduU70dULnr6cWZOKN4TTzpaC2ZcRx
jMJME617WDxmCj3dhFCS8rK1i/XEOIL5vBusDVxkG8w6MjzF8DQwyxyEFFt4btm9
Ci8xKd5EHHSfgeGtAvPvuDaSskdonfIRip4e9gRjjIG+VnF+KXPKsUfE4OBvuisR
y78IWwoOJwQOUXbMYkDgnRRsolNzzzulVTZ2EGeRF3JhN1rYapGB72VWYDPbtm05
B7rXYl6dXMpfcVR74lviliXS3gHlPosSIUilCQt5yVRFcFHAP7Mu+VmvRufYlEyA
YedcVAamH3n0Sf2UQKkXTlhTS5t1K2BmRtwcfXRtHPKlZrabmddpyaT5oauaG3WT
chuS5fET1wJZu3+KYarMvrs1qGzXbdW4weUfG/PB0MKxk7pxNCb+sXyhFTz6TdqB
8x74T05JM4rXnlYwS2+RS6Z8WbsOLmKzNRBY5fJ7gJg6myY0JgvXSj6ki+PeuOAc
d9x9RVYgvz+J4dNB/NwPV2EI1hmjAvbVuKooA/cdpeF9utIXZggpKgcDWhctJ1VL
A8GBPvfx05qmLOzT6kbZLM5BCOKr/osih/BQYJ5qjjCypsQxftp7Sg8wOBEoA/cu
CHtbQC4KcXufsY6Op3ZIUboKe3XeXcA1mOhkB0ZHh9YG1V/V7KmF84JEB2Oz3CXT
+xRQoNmJ0gIBc8tvm9rXBhWlDzc2TqE1zy5pNe8yPNkRbU26bdzbQx/Y+fNHCaHE
Bf6zeYBH+hoFIU6uTVcuIhfgbcZh3iZvoQahBLp6eCDNCaxLl+4GipVk8iuMiNzp
wmNfgDAxTD4YD3kyikzz6ZFLix5XCVCMTWFAt2m99MA19ziPQu2O7QfsqHWSqy5C
6PzYCUsiy18UIAJPek5wSq3feC+7ny0rgxq3yj9A+ICXsQPUsokqiKyrKVubYUeR
29twLJBxlbzCC/a9SPGtpKyjE2o5YUIQvXYQ8r3elSiFvOOXItWmxo9eOIFu3qHv
MkazfRCzTeMvj4JEARuboY8kDBWajB6D0sAm9SeNLMsdDz/t+pLHdTfoEGgssVDQ
bH071rnKyyj7qS8WwTQrBLZK1bvTVQANDjBiMvBEc/duPozv/e9w9D3hkMY8vPiS
uDQGiPLiuy2kSolYTPxRahALWXrySSsB/LDsNFq8jEvcpNhSn9iQ181lV0YL0pVC
ppCMZ6FM4sCDng2yilFG/Ajr7mHlY3NLcF0/ySlCKG1D9Vbrn4O50ATr1WVcUxd3
KQJYEvG32kmSDabr/Z9RZ1xauLN+UG8BlCcuN+yV/x70nz0qxNtHaq71ylUzqWHJ
imxi5I1bm7lpj7gCyhGwX80jQns5MY4G0qC0s5JtshDOdMAw5OGrakwRlShfoZUI
scZlazCo7z7jcJxAjt8vbCftiHG5tvsXvKpWCuXjBo8TX7W71ZEwi9wlpVqKvx7I
+rOOvx9Ip7aIHhWdsoRADZrOWVezSJ5R7ItB/eK+4y4sVf+h6rFTa6utX5MK6emp
EZhJj8eBGOFQIoheWI9x9evbvIFDF2TDtsFIsKIFsjRGzjlE3ULiAprFRThmNPZl
GgV6KDx/MyByMC/hEe0eAhtOshPsUs6eVynjPtrzxsFMpvU/jOt+fRykhcgh+7VB
erVloGdXzhxjzSLVJO6Mq5Mfw10XEQN4Uv3WrJdeT5g8TZ619ueSRyT62srokgtw
OtNBUCFdVFX8TJJjETEBPiK+7sDv+Ae9uOX2amWW2QSHWLyWmScdGCksJxIG2XiB
ptsKFLKbkKE4ggLFWQeCgodokbHYmUOCJrqNhudEY/1spfE0b/ou+lrO5A6wZQDm
sgblKbZk0QCVMuAjrfKhEnbWuSpRel1TuQ3QmGRJhcJpfPXr1gaPm7jMj0fo0Eda
iFcpjGxwITDpBuLql6ax9NOcLd5uj1FUtRjR4p8z5NcyJ9hj/KD9LTr5hB+nFIeF
1yzQyVqdXoqTS2IL1Bmkq4JuQriLjpOSCmn9cpXb9gB7O1ysMnIwggRl3U1rSkXq
nGnCW3mnkzHm18XdobwyiCrotJ48oHHmF+KBo/hd9QPnqrflHR92+KIP01Sn/ZKy
EfNjlI0GUWXCKuf024M24vmdvnn9JVxTRKLWfd2fzoTxMcHjVq0/kpTKNXbIMMeI
LU3mg1re+zRiLp5XKNWkt4cDlAuovMvtNQGBTKh9zCruyhj1M6dE313nHaA1IwLI
uz+RQgU7FxFEAOaE9UNCjioec4WktZA7BRlU7cL7B2dSkefH0mj9j3NiCdiYoW2E
qQqCCRN4WdW+sAEd9yfxwN7Cyh2XbmlafhagNunx3OmXNXkSEcfD6bVGPuxJuUlU
ygGEoGZ2URt5GhoRsO5HMGFP9dntC6QwNu/kwLErFY71wPRlxiifzxe3t6u11swy
jCAl+W3nxnN0x7SC7NZhF8EzlTT8ozZNZZXkdQQo1bR2hE1mgr5RYvIYGwMapYha
6usUyGPuc74txTHZyhJXY++/EY3sETa3hcSI8V8a2jVEaszFHYZwJXuP6dkewRID
5p5dwtD3lO1nsqKRWtwwWPa+kGG0Aqn/TAawEyhnQod3rwPrko6zNiqZZbqNeKP0
hg+2VANrNhNTPU2rvWXy2R790KFjY0/bw91A3Wc40BLbYDryb0/ps/3/6Uu/yTQ4
brlEZdCU6Hw1b5i97lu0S98trx8/TnXffzZ4JMO7aaq+miuBwSN70+45f/JaWmNV
b3CKuIJNZQhoA4XMd9lOsvYZxA9gZKkApmQgwRw4Zboy+6nJtl+JQLRXK87yRoMK
NBbqfe6js6LFFCl/Sqaizf33Di3PaEYaXVhVGBGAf3rJRyHCXh4LcCm86um9cMe/
ex+iXQQC0wSmfFoylQiYuHpGGGvg0j9J9SGm4wnTFJUaI9mx5Kb490gmQUwq96vd
yT3p2dMrOBYaBQViEQQLJruL9SMtZQKxyKmO2uZYv0n2bbRz6Oci3VQZdlQvniiw
lKyunyIRPtVt2eecWkDFB/si8Fkds36fcQhEgm1DYPP0WokibMkGWm+SpRVxKBCa
mWa4CPJH33X6QbzAVC2Ev51D9zuKaLgorVZ+NOH6prVDZdtoWP2FJ7/0bFVYClHV
foHlllFBtg3UKULVALmh7U7UZoYYr9FYctYTmaX4SQlVq6YdTZYd+95KyHSLBsBo
Cfmd2i3O32YKtNnN3i2ZnAhCEaQMrfOsqs7ZxNEHkrRyXuFfO6tPvc4HvYGXfTrn
eqga1rowSyytrOzl1G2bLAvpeWP8XfH2Rg3r/bVah93u3MXtr6+bK1CFoL5V4SNe
Y0KbzongLrT1v6ztruYagA8x4rkvRruryZw0yUoRgudoS3gr/NUQeTtQubBrRtdp
O9gG6eRKwy6pMggv/j/ALQHUVqmP3xy0Mpnn0OO9vO2ltuH9pR9+e+/4Tb2Lxb8O
+/m1ILNaQe1LY0ArzHB+QgI/9q7vHneQH5PGE/DpHeUX9Il0BDW4xpjP0iFKtk1d
cxBPWnVYFiKVy1Aa4Xk6kdLfc/Zr4/uEdzMAnRw5DIoUWXpqv0RB8gCV+9jXJ7Xf
xqZlxtTP54ZumYSJelEvb90t6aqbbolU2STyiRll7JsqzbEr5tiCxUPkrXy3Hzhn
k8CRlkfRaO8378zBvzIE5y17DeDLjjxt/ar/wlz7qnQtrcyO+HrG4sAbe8vkknrS
xQnYPcPrhq7H6jgEuipGApU/rjAi+2HHiGau0LnHTVZfehCRaJHL8v4XRiBU/av4
8TVoThejlgEWEu/v88g8cJtxTiAg1CTugUUrv3cTRNYxLejfguB9f+QussYL9cn8
238k/nf7mjGsaIF93AxO91LVtLETJ2z0y90QqJdUrJlDEO35Tm1kqWcOYkrR19q8
4JNVRz+CLw5YoB7XH9Tn9du5FwRDBxiXcsix0USFgKHL02LSzxx7qGuNAHZnqsl+
/N/uK/+0gSvDDwZPx8D6lyq7nX6d83zcvIV/7bq5mQvfZ8uTjj9mvre81QRyruvy
JwK08dp4ilZEo5w7Qp7Rd9S0hawcGJVw3S9/B4SS7g+r4LLbHHkMp5Ml6gDv6VJS
g5rOlHtxpRkNAcb2I9JxmfeGpeUHsBElFs0XEV9/p463JSxQr82EgdlNVhkb/Mtd
A1siWRIhDhVGdqIV1Mfavm5cC51G4k5RNjs3CCxhoauX83mC/VX5WaFdeLvT2WXm
dwjMSZjxgrBQMs3OrE+a1kHkaOd8gqK+huWUh2pwaph/8apQ2FMD55abB2oj2o/5
yaXjDKc5bXmlaYOMYX/sbM+b4kNE2Jg0ZuS8T2Nj6PUfdrXT8gyKHa954XvouPQO
3dh/Nry/yw3fjAUxvxAOsUebWhJh5XdP6DfSj+YRJoqkk4E/k4xCwRn0zf/vpL5c
ZrsTvoV5JxoGL8sfQfMKY5pPzcBKI7WiZenFDUkZfBOTfGohgvRypEvJUc1SEeIY
RfD/VxernAZT+PmuSCNEKiRmYOJdKQopiIhwBtGUd1d8zmYiRMIu6fO9WGZHZmAy
wg2qP8tAqXYWDZ9MK6HjCuPA74eK1jT+EUCMdX2xQQuricmosqDajEZ25TgNSjvC
4floNQNvmj6+EYljBuxuXPnJZKHkw6+JBfULufKc0JYPXNtY0Do5tXzqt0697AIj
k1uATz9m0xFjIVBLLEuae3U8nHMN5O8QAg/Bc5ZyIiqI5vg2lTxkB/4r3BbrQq6W
6MiSCrKMI1pcWaZIYS30u0akURQf2ObzhMPXFY32liilNix+nnuamR+Owbw+g+rv
I/fBl8P15cpSUXaz1/ItmbJALxP+GVTmECuecW4uc8rRPTR6gau2eO5T+PBoJy+Z
jFHERJpCTgM6c3k2Fgn9euzYoF2u8q7zERo8sA1ldrCZDIkDsPClvyeC6KD3JIg7
/xN8+0s5/HSZGWOR10GGLT20YnAFX+Ra1hRMTpIeLGugYV5ED8XVqN0Z8inYGtx8
FRaH4AGRJ2mluYwgAfbRcHKjb5RRWDeHnVQ+mIK/iwpT4FJXVG5Ieo7VLAo2DyV6
Pxru8RW4i+zxjY5zYvjk/QEkV2DtdrY4DJDSQT/Oi1Zc/gHG+MFgOYBIEj9hgGUL
aep4rQaEkSqesQ3LfVbf0L4Ay1avJhPeYZYo8oxFPp4rRx3UpVJg3FXwY6Fo4kFl
qEQwqEXPl7HExKqheDymgHbhpZfRKOxFwuH1v6q8Htt94uVVvZdD7PihNj6YWck8
O3HLWswyG1l1uLMrcGPJv/3gdioQln926RHnqK6ix7him8V9u33ycvw+gWQ9r3g7
jam2Po5LJdYETM3kLte5liNeLApLKx27M8MfEdvQJS6ivl4qKzIeTzPZngK4qnd2
aXNj7Xc/CzM8flKO8MtJQ3jnuMywgan5NMUCLHesn8PIUAvZfOjNmJ8zCMlR5wEr
xAlM3y8d8KpTfdQQJ7/7z2+r1hfKfySJsaPy9bUBgHuTjdFKWiTPv/mZg3ncp+Hu
w672D/S15avcaV4SFJ4j/m/p6Lwi2CZ1q1M/qFb2UVsfThxI/POp/uDZnAlMfNSK
pkUkRu7SpmboI89+Z2FBjAWaAMwHeFXuZLi6Q0yz1NiYTpTJ2QoqBd++rHqO68mZ
Qp7VOi/Vqnb/CtcUbVwWyh42KwnN4qyAw/QOiJ7+XJToUcCH9Q6h+2DhVrwvydQP
uz4C9nxeer4c1VyO71+6Tlup/9lL2ZtfZ2+Ny3Xa7XvEzrFIFbUUWNL9ny0EooR1
ZhscbS7hregNZISo+6ZnBnuiaoF1ffgOgCDi+YR/NoCkPhhsA3dmytR505XKgjeh
Jw3VbjIUnAmlng3AKN2YB/dmySLI9JQLcsuDKrcz1o8QlI6uQPt42S+yI7zv9PkM
9HZ807OKMZBuXr6dJjuYq+AHAKgu2IGr1YnWowfKja5qBjmNG0zPR8XvHdl17xSg
DUtZRQVSL3/8kqO1si/PlyBXHS7Z4mnVpO0SgCRqBHb5chNLDfarGdU9BFjSCnMT
1Y4sBszBBiMhsIHrexe4JiGLx24+mlvSB8djMuhYyDEond+NRdUclCzuncRp8OGd
7RLu2RNkSa2+9iWUhMclbDKwpAJ9gLfGXAmZ0tq6rQxe4QkoJeSSLgIHZBZ79acQ
AgQoLX0kATwrmp2iI4IFHfHNWs0+x0VIeGMbLJ5k3fDNMfIAWZgqsDfBQEdNBB7O
nBeb/PXkk/Ilw8jY1xOVFun5+Cv3xRpGK2ROz4I+MB8w1rkcQwEHX4Jfosf3I2rG
STGewa5/YEyDzBFU71BnF4K/z1kSH/O3HYwojmZcdLpxUM3W8iMX7AjglL1xsmYO
AwydYqzNjWZGTpzOC/7wOqxVGxpFCHumZRUnNaqOIJejxW6cv2ybVvjW+DUyfQI7
5ZQeP9/ntxkpLQvxmjDB5DfA0cnubd5jY8z+s/qUW8XMX2AAFV/xamOpd/kl1cnx
vP+Wo7tEG2h+onFpfb+EP0sVTkf4il3yh8vLVr5LFXAMpoF8K/rFMkwJSJ7OUSQ2
BH+I1dq7i9VtDMVNOWj9sjryXVs1V8ubj/GXOSC6vG+jvBcfLSmKzJQ0EXxKzZEm
D5jwvnNmToLSCY8Lx34qBAcrVvDA71IWv+vVoog0YSEDNWebBmYKVmZLM1SpHQ6h
otTwpVbK/Esgtu3GgjDRz+er60YYHD5/ocBw/pLIR6p+UUVJtp5sGDg3oACY7S5e
QhyXr+rFpl60V39MjjYiqrNNC5LpfICT2xwMfOnGl2vJ3KUxUiiXT/zw9AcaSEdx
d71KQlrM7znizy5nPIifVfczr6YLcfn6ZyoVlWdkt46cjkg+FlWqefFZt1xhLGpb
vUpKYm8IPH7jww+xUXh0n1xu7/5PkMa58kCEtVNSVUFN3KIxMudXd+2w7tsBKFtk
XiuSgJA4Q5Rqs1JhZcyCKbr9iJ0MOPADK39besry5SIXR/NWFKCI9I6WTjPWpFIp
vJejx16vszIywJR8Li1mFUd8D1X6UJl4IpWLqKA+IcKIkEcK5P278jJM2dXElZJv
WqoIbUV/bpCJuRhfPwffummhDvDNkWOKaa/5FJvYLTMngzdlKSINKB6tX8sNZZQW
Ya6l+uBEgXcIv4/Izumt8fj8ogTtornKZvRShVs+mxz0dhVWb8UcLsxf7syNlYRC
OOxkUS0KIwQVPVad9AsQRMgvretrTEIUW3N4TaHSubgZgb8+LOqufrTfA28F+ZaT
NoR+vj7xqdt8fWS7X97k8N6ZqET7t4TJ0Bq3nZT758hz6Kzq0Tp4TxnHY/CYU/WI
YUxjS1CKfymr1nLxHPfDm/sL/NwJ8oG8X+d0yM9JCj46OHhbKw/r2AUW15zeXgMF
/pLw0H4v3MYL/5ujCLVefTJIfTkwBAriPwdu8f3f4jsva7l8X7qfBP1TZFj74z3P
GZPlajci2iBRWaiKh9Fzf+FT0PFEkCifqHEykk2WxWL5uPZ4as/xoAA7AC9yiPfB
7pJm8yvhGBHMpndzfB+HIRy+1ST2Py0xCEgmXjqoToAZArJ6lpS/KD0+KcbELgIf
R8tlHyngdrKVeqz8faw3MI3KGgofEp/h6rJF/MT3GsPI++F9GgzQgzZgofoYHul9
m7ow9BSmtPg4yBq3HSJHtGU/l8QVzyr1QS+LgJ480CnBnMX3+eWfidcwgMaEdKQt
kjhfkzglTzW4kKoG9pZ2GMR+7k7zgYqJ+RDSSx8muSGX/9T3cGqhF50Yz+1SPRCe
VXEszX7EjY+aNixRdrEOIptAiazldILWRSrT3bE0pytj5ZWVYXLe5oMHU7aTCtud
dINKGzKnJZFqlvDKo2jjqr+80ztcgMeYN7Y9aFqp3Bq85Imp7OAvR4SziZ14v5XE
rMOjVhQQfjuy2mci7M2iAEW7XwIFX28ZYjQplfzPlXlxCAqHvdnpypdnDb2rMkw5
+LU7XlJCPaC2FklWeujuQrqk4LbBS2cfYRKIw+MvutHMrMXyNvA0VGudxT80XsIi
mlIyrp+T6HMoAasxiocdUETUNj27Sl4pMHSE6Mdoc+ZFHHOjuLag9tREoT9zhW75
caG04HAlGxo7bMSHYxHH2INcH1lGnoFIrpDwiuC16vMqU2lsOD1Ta8pMmd8aQczw
ehUS3DvOWQifIF9+BgcoWSqeUE3pyD9/tiJFLgx0ZIn/hury1tZp2EhYdxe8sWUv
gQkcxSzLHgGTSt/++GVVyZDctNMV/wkzO3NY3xqH2XtoThK0s7YQFo5n+itLTafL
jV0UwopspQkvERlymwm/cRRcgvf1ElazvtNAwoC9g58SGqSWMnVsiLQ9HfVILm4C
uOA1wN/A6FGcmRZ8aaNWmhAdHF3gUklwZs99pL+uRHgMaQb4tKVcoL4UhiUo0+ib
tCWaAvihnfkKgpN67gSoK+uRz7oFqgyflrtUExE29kgfxD/cXcR5ENvylse7K06u
KB1USoOEmjnuUN9nRj+Ni/wucP1x16j9JbKnSKzREgHIfEkfBXbyytTGOI6heys4
Fa2vRvgThgMvpQwiF8WOiTaukBf8eVj2n36+dzZzIDIBo+oqhY9RQtyO3MnStQhQ
az+H8WoSqbbwQ339VOgvADjInHLdvzQGcPcCMYVSwHV3O8RWeyKs5TK1UGYl3yc0
PQs+zOhAAGtM7BLva0CBbZbvzmS3Xe3P1jq44i6TREpkyoRoMI0YtlRN7d+96Bam
OqGE2ObcEp8bedFF8+ZknThLgmPaZ3/7wNPYt1AcpPRRLxK4VWeuf7odeFiC2ACd
LX2MgkAfnOn8BpP8SsiyEVNQoZuqKxpC4g6Ad2Jc2Inc002dC+LUrfyfUvaeuPti
daFn1CljsPEoj8yl0VdFgEvo5ik2n4YSCcIR/ouy1ljlKLCAOuv5Xva0ccM3k/j+
CnvE0x2ZYJumN144M6Ek92Gu3o2JkGCq3yARL/wIy8oRCDHEmhB/C6ws+aemgBxg
qmSbVkAkL6whOmtkXUIGqemHPnMgxn9pZwTbw80zxDF8MkMGBW0KMYZhiwUfk1AW
/2N4PAwfhfZsPv9Z+TjtWUxqhoUjwZGyxCV+CuGm0XO4/rN23nw89wMpJyQrNKwb
yJt2PvHfMRhm7xAJ9hEbiv8qPBCV/sfE8smkTHMOloJUi4tplrA68DvxN5RbEuSd
cSemsFLAO+79GHVEiTngfDwzGMUKn2eBKf0ILyJg7F6Cxqp3HvdkQl/Yy8FMQibd
Fv800S7zZpOWRt4gAShDYmeslNalkTB/C9nPKwdH2t2f9/JgD75iXSIWAZc1LI2H
pSdzr/TVemohosVGbtRDBLdGZy3UOrjtrXjbXX6TLJv9S2Zm1dbHYOqthpUfar6o
BW4JB6yVKacUho0VS3DgTVDxFn7XJ9QgqbW4fZFgm3nzA5bSXeyjdIGcNQTdRo1w
i7HOzJyJyuzHtgb7RE95pyFZcbqNi0gn0vJPssaloSHyaiLi8isRsb6tjQPbcdz/
PgDGOXSb31jTA8a9vOlkeXTphezuYhFPXtbZ946aseI3r7gqh+GJ17520iG8uun2
3eQsyhn5KcS/hOYhcEiEiWNj9LKDw9rYNAIejEhQB/YIMW0h2AcvzBcxGT8Gg70g
bBGfYTFKiVlaUMNoEpCXJAEiOU7IYcdDJK/rg4Z3xmN/amxyMc3vFzp13IS2zO9p
2GZAxr12aXQV3l4IRUXGgYS7N6mpdQ0DRLebCnHZ1naGCngN/UnOZtYP1JxKImsU
lKj53MzXZDhVpOOoyFtHMMvhiWKrjD485iqhFVlKbGxm/lkhZ8X4bh9ZfnLpQqRa
GXQIBY86kIL9muOy8600AV1rpWya2jddSuikg43l9kp+Igr2ikylxxx5VFo4s2G/
yqnoiehxl2SMAvnVm6dK52YM+pt2mUMkoyIX/8S0/2i6RmQZVHtdDKOMnui14BF7
k56qVDrWHqIRrELD06gI5v5Nlhy3h7i0gS0iAnyrDpXkIiLgM0Ea6528vBZuSOHV
rt/VWDKQy7et+aa0PYmgB7tp86WtwwUss4EasLFfXht2OITxyEvN4fD4ppwfEqes
zK8FPSUlxIdOmgssqYqjYx0zNGobJjlV4yFwPswgNs5e14XqwLom3Xx6ujBBWk/n
jHJiQi7biBR7ckv8ljPcU7XHNbYXrvmaSWlueAkxnyx2+3oBOUQmXsIR8Y8RolzO
8kKSTF1hnkqrBk4KAussj7BNtWtzHitOG7X74u5ydasrp8OGwkG9uMDswx9vJFLd
w4evDzzQpsO+NqI6YE42XvsLzxri62Tex6kblV1kLw/C5JcTZzhvg8/EB74p3c8b
oUGvjIFi1wbGW5BSXS/cN/y66jfrmC/aqXJ27andpesA77MbsTym6fTlNck6nhqv
g+pwOCqa8Vn/9DoBKefp+uh/Z9DbzaX2qNU5LgbIVea/GA/9teM/MZoRmOZp7wVb
W3H0FsaYCdbZ7u2wPPNyMaHtLWMAkqHYlKlk1J3S7YiGJjibjc7bMH/lSeqgjtVq
6QnKCpojVoH6+upx7uiKOYFdSbNFnUxko3Ias9LCODlHCZjboDHASWKlZAfwyjCl
wSfiC7Yg0XTboSM49Kc74sUeesQBken+P3LxsHsG59/Ka1KNzW+14PxyftjOMBtM
b+ftNa3xCSJYvHN2dnXS06ZiyiIjiyouwKiHO8yUe7yDW15UWGfpKTtIXCyfKG/D
8lT5cjCRiq2bJlXgTkqqpo/AE2GzJVEuEoBfiH+LHzI0+OD1JjP21uUgELiIK8GY
ZUpt4D6AQKWMhaaGMHjOe3OnafQroYwtklUmkhCAjkSweLuaMhqN9Hzeu7G/9+aw
REu5KsJBKKZheP2cjCn/ngSUDRxxQ7GRyzPFwGB7t3NGzI6swaqfxTguf29rvWv1
yMTAepqyWf4BAV9Dd1Hvk0or4sBW0nedObO6h34eEzhA3xqNkHWPR3kcIi6w/eCN
/iCneAHO7bdmF9Lp5uJOJIJauSYklQVhqonEkap6+BlEtQSNFk3WkCUr/ZC42ffa
Q/hLmjNTdPq4dgFri/goOvOFThTZI3+rGVkhgqC1ha1Fa7uPnxfXmngSKRh0ROyb
9RiyQZ4WpurI/7s4o0LjPvvjsnKqm+p8055AGcYSPTLA7A/t6oZ59Vlq6H8Ue8M4
5aJYURQa/2QM1//1z6V0Rm8iDOucGW4pk83qgNsU517l0rQJOnvq0peL3EboPhC0
tBl/MskKCmH1bAblTmwkE5B/c2mJhPGbTnar45L1FcSGAqujf8D4acNQMo2HPv/b
2swgXZu3jZBOOUkHm6AOYS/9bXCrqWsca5lkdKTVuQ0PFuqAYLaKQdPOYNCKuHmM
hq5hT/9QRpVlgn74+KGncCrhEI3L1YQqDiYftvbi7/StUp3jVvGpImn+gN7nJUKa
PBDJbievaO2u3mKq74/+e3BqnNLfdyaIYW0BpYSGm0Qe8r49goKk5rWnVTGbho1p
Y6Hi8ZOshAPDSCmXCLNTabGiTl0LDL2yT+XjKqAsVAj4aYKg9PlJ3PykWBJl2N2R
mOrMfIaKv/KW4/of7R0qMX3Xp4EdW6D7+JPeTePYwnmGU6ilBgfRjWZdRlA/xx3W
GO5AqOEG+i1YuHIKZ9u4JQeE4W4SmtNmiH+aDLUMDBhqvfJxKOuPn6ogAh1TBdvi
g2IMSOT2Te8PWk+KEXr9MNSfBSHBAoDMftGpuT0/FjguLZu0e58GHJwlDamW1MQo
9ZZfErq+t/0VJFgZIDln8xz2+M+C10tvgHAnFZHFmutz/KExWwK4ojBxc8KMOGmb
o7L+u16ZWUfwLfxrXQ1me2Wx4HiBkS0Ik2Xwmolo2/B4xAFmPjpK0EDM6gdvsb2S
buBLzVxVmU7w5nTF9BtYQ8kieddhgVT6vhMf9vIw5ZQ3F4GKZ67W3Ifxgei1wDvi
WKC2HDNe7+0L5sRBfIBv1yUMdONBUIsFo8NdwmkjCed9patX/4YRveCllMTpHJFH
Z5sQv8kEhqMklt1mPtPW7TLGcovmN2TXAmSKAoM9X9qLMAWLLe3A7MvIEJ7fwaRl
d8iIPN4dDLTMa4+OjRwxTuykzi5mGXgPPb1N8YtQC8QxZhXjOTGwBaSYBQ6yqRWv
Zy6z66xMK4uhYIbBjr7gVSKRDft9XMgv3o40Aj1YKDeKrM7kbZKqP7selaXhlJoq
XCcHd4HXxexCz6cTR0KwTNsF5fU1vDt+FST/AxsdIwl2koT59xCpFVoWHxsCiqxV
7+ShmeriuU+MM3lsG9ph5XagrhDaaoJhySkjADKIIByGwzi1p1gi/D6PQ3AWB1mZ
wtrf4n1+vtuwFbjzSIjFXfWR01p/llBJztjint8HMFe3WxkQedxWgB8TVCcqltAm
P0eMXk0fCHs6cJmve30oF2Dm/0XudSZOY08L3fd+8QAwRIxOP/o5G/Fas1HVwm5s
N8giM0WoBdGLJvxI262/IDUjCUQCVVExY+dwmLWUojfQCrVffUFBdZePmj+J9Di2
t2e9SDRZ/DB/Id0DQhGOvF1P3WU/0+mqxj8Tfh5NQCFBNLNUW2WhNOF9jH9QKQ77
FYbVYYkP1j1trqN74Q9iRvoWzCiTKpeWyK+dSEYwIR3z5EQZLOfBXDKnd680l97Y
F8nT9fBT91gR5fZVsfYa/8ymAyiikCBl219GB6TJycNnXm4uu1cwAThmbkBoOmFN
cx5iLW05sd+kPRzYJn04ZgqhKfHScmmwOoEx7vRy6UWm6aS4OAhxvVFAaWI6JFhG
ZQTM2UadrJr+ou4c/e2UmA8aC90TZBr0ADCBfm3otj8Zw1wfvnRGqNAUya8KapTW
wAiKOW6OycQNIo8advBM52ZfQT8nPpZhAwXzNEnnI33u9yvttCp427SG+LKWE+F+
qrP0Xuhh86RyzcetZnhClsOSVxyWcrFS2GzXYevts1dgu5xCMzZL0sC9e2t1avhx
iglqBEEB+kN8yUZV3VnmW1HG6j6ByJPl196yhSPl7gzHrH7K+Z25GxnRjJw1vQaZ
i8m7UmsXXB5aO61ofkAWye9sRJeAVYWqw8PduykwBEiJYzjfkGRY5IrDkET+kxas
n+Bz2bWECM1bkAqssdB4K0JCIqzCpQD1QDh0lhBZ+MZTmcUzBgZQGEJCv0EgEDjY
vxzq7YIdn9DRvfETncc2xfjs4E9pQGhHjdPc+EHWvq4OYT4nwMOWsFnzWCBH0zmD
MJ8KimjPoWPIjDIst0CeItf0Nlkzu5hTltM4cYtj8n7Nt9o3d+Vu2jaAu8XVyadW
PmDRnpXLNLECGGMeoUZDkN0U9iHF7yr41ttuqUL78jib16x5yiaU5I3nBn0tAAq+
LZTl/Uta8EU1EGZnp56PrrTy0RjgW7taCJqANoaxxah6DS7j7sPyq/B9HedIM0XG
IobPhDZx3AiRAuhp7cgjiKNO5te7jJfq0Z7rfPTQQoH3U/Bi2sWyh4PmvsqzyoOb
IG+xFHfeTN6cywEVL2l8rtV4OKPglGCILhgs8MbCkbfZaRrS6JDjeHkFUBobV5nz
aVTpRoGq12B1Mi5l0ijLCX4dpXfuoSLyopoBVGuHU07Z/lIgByi1d7fCM/HuTqBE
H8xP7oxcqheTaQ9Qg0ZM05STTXP6/0wA6BTa11TB3+CfWHQ6xmo+9/JTuwPsz7OM
KuIrRKybO7FsAQStCZOu6ardKvthcGyECutnDJoNlHd0I7qkN2fUHK/68bli65C7
hyz/lpOjHySX6DqzyopkEq9jZ6cgsvG5P9ptriVFWHe2U+uYCZRc+NQ2aO1zR1cJ
5s5GegCbPuC0aJX41slMRLLRvG4rCMpeTQ8lPWwUxO6Z2fHPYFDt0TwxUi5Xi48Y
b46cNieoWln3k+ExHkGsqv6xFlyv31X6y/YrxwBVcZlyk3Vre6cT3Y8VHxdc6ACV
pFPapw2v1DvWQYM/VGmSHNExSLwGF5+HB+ylI2j5tu5XfObh9oB5tlcNyXtv2oX+
gMe5CIZGtxlel0bu1zYeeDYclXIhDa1NwgcTxEvXaoU8lAqjN3Sl5vjBgbF0qpmA
942scE8vG/GlDD+UN35Ip2+0r/5r0TTL4MP4RVsizEvW7Fg6SLYDRQF5TerIuak9
FkBcv+r0vyofbCnls4uiS2e4wI/coH3A5aUQc6CXHwo5ibxj/pXomIHKyU4nu/9P
FCbbK2oHxKiwhlMIzCXwVDMumvTaqD3r780CekXVyrQAQc+nSlHFCHua0qVVY/Xy
jpWhLgp9wMiv/aOL383LIjKvFsS26JdO5civ2Tey/wijaEsILcMk7sw3Znb+4gBa
QISHucGDeaI+Tch6Dhn2EDq4JjaPwHlUrXIHPIlEXSFl17MmgnNH3mZH+TCkpShi
7GZS1mQE90BRV0c9xW3CbT/ZDit5VI/PkssPV4134x+3mA+SkEV+RMhrpa/5Gj4D
HvY+lotH/jTfX0NnbmiWnEag3YiH69Jo0xz85WXdiNepy8ap+Z/4qCal+475YHxg
sFmqXJ+IwvD3VJy6IHgv7ax3XDivZBkKAYuQweA0s6ap+rWuS+dh2ZEn0Le66get
QLqughKtmM4kp05jNGCtCnUtlUE/fI23WbcriRB/JypcNfDBg/NgZ+90/iRs4HKc
2hmgxWQiars5VeLiIXYG2Jh6ygt7VYZTmqsVe6GQtEIGoBDus3BXbgLeXxfPBY1I
HGnQYbmyA09OHylnP5MyFMR2qos7XF9RHHPzBPetgENRkJfPiLvYtAOxU6m0TQfd
c8N33o5qorV/qS5i6RYydYiaVS/eycsBAwgOEbG0OY2D2mftIxknomTsQcqeGp3h
BpUyTOffKucDycsspNDGzm6O8YE/qe0hpIhcEwaV0RZQyWK4wuTl90dwvqiXTpbu
mcT9v8pLvI/t7pkb/5kwG6CZfnLu7wcvogAjpqPNJKAHB9d+/3ABC+Hu7oRjDUq+
dXDuZDB6DrYgUOj/mXu0jc3KU+ZRth36GKxz4H7QixIwpbkSV1KnNwZrJgO7Ykgv
jnZ0/8Oq39zo/AfCcABoAaMARTSj7tEBcjpuskN8XZyEd2Etruis4kLGDP9Bchcw
194mD6XP+kl0wjTNQwDEwvwsHj/A7zKdy2uhDVHPXsFP58dTYqQiZbh2bB/jRn6h
0x8vVWkHeOZXKXIGEGIFp+HTnXvu7JvH5KBDGkWREgZvlC0eIQL9I18fRJx5L5Kq
Gk4tUkK/M/9TuKu4LwNyh92X5XK7uN7HyRAARJcYkJ3kuDM/gyiCZO5Oip4Oj3if
TKiQt5jTV12/3OnVxh+Nt/dcSTzDp1ZtXNc5do4yltcQsTd4CAp6XESz/6dkJ4iQ
z64w1/5IBKrR/EOeybZw7Sz587hyHmaq/bvWfLLeiwc8sFqHjG3Hypp9glSiK+9d
lHgPnD+BO4t0i+4WrzZGTVQ2aXuAr2YD2rEToLQFq0hZb5xHSeNw+SrJTwVULczq
17eElRl6YGw+S/US/GKbds7cgBSnpNEAX8f9Ewfn0AQywIqouQM4aW/K3BBshGkw
iw5YOC+5nRI6q7tVqKLBMNKpi6C47b5UcLMkt3PbdUlnako5KpcphjxNb3NLJgtO
U7HjaTmMOrNVMf/+2VOygW7obfzFOpTBrOS2hNGXFhTJEyWyWdFKyrj3huzUuBq0
B2ySXGWvOZmQGJapjxZd0EG8sKrmfwh9hcQ/izHzO//p8i00T/1JhDvd67e5A5/W
nhKBuUGf+PAOTxmAcJ67bZuvPTe4Jyz61b2o5kZjywYt9sBh7vu5IziNcaWHQcxg
gxoNfNd0uRjRGNyXib6FKZQUBdNWEgPvDKSQEN43EKzbzSO9pRlVpth3BnqTRery
Iy/4lHSwvuGMy3FVQz4lQvJnqOWb4OIBeqqT78EYRwAT3VxGWm/CevQzIrLPj6kV
nFwtJsm6d78PxLLYcvBcYyzuiEE5zqvL+H9AwmWaC9XJpijXwUYl8ZscqC6pcYAb
ZLkQN7A0+A1cXzJlzLICMuXMltd2qeiK4lCGJFum7IbmRpsbb15YAmnGOOFwQ9l0
c+4VJin7UyTL7/wRFYdAQ8VPoXX3hTiDhnSKJujRnZI/35fTVbNoo7v+2SidOvh1
hY7j7wpBTV/Nj+tAeRG3rswlBMMc/QFTSk1RfTEYvIuI1wf2/C5Qx1X4ZmN/u3bo
7zAqoT9JV8kSe0qSi3exfZEqoTlSLXgbN8jRaANOezsf9tp4zqViahGjLQqAR1Bs
PKyyDQQPoZKl1GgrcQ14/oWiiqaDf1mHJwx/xE+ZG5TW66W60c3ELGwr/RJWYHr2
6huKFL2Coq2Mpsa9tY3XSMNr+fwpPaSQYrMtS5vppz8Zs0LrGGjUJPrqViP/pTrP
beEfMZP9AUtqvUv4BQoQy8aqO5Cg5iJz5DxwBCu7BPwch/PAuvI0kBuquaiY8mgq
xMTAFkSNCxRZH0TCK45bHsHgCsgdQ15mvuAYS3nJ0mUhOfSG8cqyejjqeNb64vx0
O9jJ1MbO641W0BKgyyWauyscXsJRHq7FWb1854XXNUGSSqyOFsMGrvG3oXZ2jFmJ
0sRJby2q+WLUum4KSSZ2anv6vFZlkzcPwwXM5FNe4a3OpQkBjYuj0DwaEr4smdvy
+FryNbsw0lswq05FGNz3yzlcvuNaN3mD2vZI9wGouV3AhfiEoPvDNJjnLY1T+KQM
dlfii1ArTT8TPOJx6FUY18AxvVNkgN8aS572GYFNGBsqqnfO5y9PZWhsCaNTBAqL
L9Wb0n/TPVsV/WyUvandwIIa8ehw7ZHBq+XTsdthLm1T37p9Q+QWpj0SjvkrF8FH
IK25ZTdiKiGvcWyqIvYlhpG9PKgU7x+A3RoKlbAPAX5UrdHf8/HM3tiLOvPioj3+
dA4jWZFkIFlOLSbwBkOssitCD6xh65uk9x7Q59+Gv8VgBEkVm5hq5w0jBmiyerBS
oUuSxEwngAjySZKMD43TsGNsVBt350TM/TNGguXVaF7KVyju8eecjOe7agucpoAj
ey3CRUVRtovJdKy6bKEgIcMVqahQeRMY+/1tRKKWUKG5/FU9WkElsCHtoxyzL8Yf
9+m1QlLRLKZmF/WgBzHLfvN++Q4C5+IsB7tFOpWGRfiBQ50eroAqM8zRGuKlf3e2
tETHdFhhN7OT1eU8zVRWHUhx5/+epkwrfmDlCtW9k4MGsSbMuQbYbVlE+BvWTmsQ
StZyN3bAZww73wWaIKOFP0YuH66Har4zTAEzlhqBMBgUM6Tu5BRYLMcCljrsMY4t
v4Tf4yj38QyvyJit1k+G0Nmms6BGTzfqkj8IT5eo4oe5Yq87kWxme9PgDnrzXYhX
OxI0e3purlI9YZDn6wz6vrZxc8lVXfiFO9/0KVvSBdRXew3cXdp4ZV7Jvj5Yvz/1
64y2njAI6PI0aSROZmPZy7A07pcXUYxh6sP/PGIKK/RhY3lNmxRXDl2Lyb1XP56W
3IhjMTphtLFxNshs2VkMbqwLNNp2h8gd7AUYqWORLYSyw26PVoNF9G7ZPGq/+PGT
a5oDYqh8EOd3hAY198+3gJ+NcMLhGpbhS7AnlqideLhzntUDE1vAS6MOIu9TXSEs
LUvwmO97vn/LPr4fEl4J0fhKvcjjqcAL7rrWtDDC8IUxAcpQfQ9FMomYqBfXc59m
0YH8EtQW8429E2gwm6BXLKz7NJCiCXnaUQRg6wfgIZlg+DV0xIPsgBqS4Epq1cBo
/4p4CAgXD01g+ThQtR9uAo1QNZPOGM7W1CFdPyGPWHXdLLNbYwGvPjgXJzEPSPoj
CBglyHdTvl9NPlUD37ygOZ9Abed3UB1Epc+75nv4KD8M/t986vE0SfNFDegGMYJ5
8ldO1K5z528FJmoONWSf6lcW7ADYpgbCemqWVlO0u14STB5yxCfWKaH2Hk5w2til
3sP+AWzbOQb+nu2UMNqpcepqIlwwbfwu0sIwWYzJvwW/ztroesjLEhLlcyZWkCxL
u/tHNNUGtUWbHK6Vhvb3Af9yzM6wkwWmqtRMnCoEZvN5QGPkWHr1ddM2b3ApruyP
a6vwkt6/gF36s84mxJ57u2aSPGuGsa15jpWDScX5zQSrsOgz4hJHFKldQqR6IReN
VvHxoz8hbcmtyvBBl3tszt0UUgAdXnNq20FYR80CcZ34GHXS8YYblVjSplHecl+C
9uPh8Fv3D+76+mwnwkXS32GutY9P8fnF5k94SZsGTAItsbrxycLy++V0su9wFMDX
3fqxeCxTpgZo0NFaf3bzaM8iUBAEllYg4TA4j4X4fkAAYmflBjO5t7eXHBBWL9Ya
emE8XxaJ2v994QOWChhZgTxzcNY+RgQv0WslseVGUmqRdPQ8GO4p8dRd6AOTc8p+
QrxUa3JzFhB6WTeYCYQMJAbpkklKcYXon807NZQb9xX4uSLZs/CVCDTm+DTx6JQf
yYghL0AC3Q8wKwUd77b2iZUpotdkXIsYmKXXw8KYb6SfWiupIU349NETyPKGnOAc
0+TpG/S6cCO/+7WgbxSE1Lsvno3L4G+omXHlhjRaO5GYRwKO81f/rH7cH/vx6h72
iWMpLgLPFt/bRnVDF6fwwx/Mxvjo9p88tneo48uRUcuY0/qKkPV3Etpkwrlcq1JX
yuIOhqtJWvTGCLC/mK/StNV/uXROo5qmP7RC3nb6uniGcZZ0V4GZbRJbLLv2Ayzw
NpJuPSHgdw2mWraKyP+Ekx2QCJ2uya/3Uozxcf9P2gTk3dV3UJx/Wg3VhgaboECD
VvjDYtJLB0zu0uaNhd8M1yn4nPgWtuq8AvEIa2fQHpiQYKmT7mtJ+xSsvWpn5xMt
RPsoJNHS7Asa1hh3/Qt0B6I0MfQPQTV6NYZS0QBprZNZINjSwrdy35+KDfgL4QqC
t4GhZnlUNIOcIoTl2S/VxRNGkwCtWrpxtD6dYlaTYWJPtWZNt15rHVNqd96tOUpH
nEZgqgHuK+Ww06eRWQw3JnmhWGE0ADE+0dwA6zrgv+7jTECMGwJFHc8Oy/vdVTKf
YMT2At7jDpiYiP5Lyk5ONgeIN0Sfe6dq60WYJMW9D3O82rzrjftrm8zpu+vZgL2K
eMtik23JgxmQjRGcLgNZcYeb3KnARp5XhIrAJOt6we0dDC77pC+giJ0YwQhwN8+A
X3dRkRpfkZu5mJ1CXpuOQZtDiZbBFh7Z3jPD493wSx8txz44hk1RM3RH0jnmGr7W
qAtf7E9bwPm2c0QGba7fh0zgpVDXXyWVRGlblIulbYzPsR7UmnsMUwcAUcwWMm7g
jNzFkEsAt1Edm7l9fYQirUyyxdd5m27bRqQEJDDhrW2S3duAlObT/f1Rfn97Djiq
kYkHuWSl4MhbNPqIYl9HCahOzxbymS/S20aT1vMPef/hcm4Y6SECNX9+JwKHhXO3
7tpVvypFvZpJFFkFXK/4rfHfeW9zGCeovZhG1dz/qhLH5iFVGsLwYe89MUWYS0k7
5p/5HvLvqDKtD1qOjhrKRDZ6La68MT6OdY4MvZLck2rgOlMh522LxHjRXngMMTBl
jwIW0d9ZzVlON+bSWO+XtLf7GtXYAaXxhpBkZUMNF1xPEZaFhO5PvOe0humimpI0
uXmRnhCYThPWHeVQEapkz5t/gDdBo8mvy4nbEXg949Lhedh+SNzemM4YehZDIHA8
taNpi4zQgYLkReEhE8DKvZixPrHbTF6zLW6lqptObwXvRG+8v+yFdekcZD2TpKgo
Cm7R0fULvgWE8wRxL/IMwykuz30EhG1WNUHSfFWi2nDMLMPCyuJHGgozRScLQRDZ
1lSZM48dV0pEuOrBm5gsM4OoiKSk7TTQHLpdac52HDdJ+2Ya+Y7GabOearrsH2Ez
pi8O+asXz+dXvPI25dm2GLQgdKD3xFt64HHgtMd+gWCFVZXUvUuLLE7QUHeSbRGr
BXI33DcXy5eFr0p2D7nDFbsuQcwLlssjz0cgTrivu0F6w29Wzr4HOtMOBTnMLlh1
lpC/5RSCvGUERTQK2QUb2AsoCZmxDFAJIQxfZr67/5ya5T44zacvLMdx7Of2SB+E
XXhf8panSmk/MSEzZUVubQWqF+nJ39XzW1J/fiVm3yY79fnIKkaEDij4dMBs9Ux/
37s5T94F5FJNLjtDha89OowkHjo3ricwpLQ/U1P/eiMUoeScGZ7QuQiGG0RAuQWc
72irzob/IAVk1HefASWM7OfHLgtDnt9+LuVWvAlx1QttyROumBWBmaD1tKn9qMSZ
QAcK4/wcdSYY6tfuDgJ3R/axYKX6lcRoGYcDNxRZgXoULki9ZGyWzBnmXEV46R1W
QLwgL5Qo91IKON/8LFLCYw5+XFGIPf7c4yVGfT7qHayfnF2i7Q46Jq+0b+G9nCob
hJx6pILf5zHFrYy5znMTJ8dcYuV3UzeVnX7LqQ72ZlEATA/TLx08Rv9GT8kzJrTC
kPcxqqWqWh9zmIC0AN6AJw6OYbVYpDREbWccI8MJJzOeA6i8Ad1U/6DmtIXKdfX1
eElD0yOZX4OCP3Pf1vVJ2FHV1ZNJIHsVOnkIgwNbb20nCv030n3AWuFaYMl4spEw
I4BktRbIB7FTOZJdAjrUlwymG4s88zXRgAxMfTW+JQRGrw9w7Fncu8XlrKjYhJFk
TSDMw5tI0mhvLvZUtT8UpLnbe7IJFiFZnTDmiPd/cRnpbscnZbMBlvu52Qnok7bZ
AndzFJZH3xpxLSXeDvcWogVdgjF6x60iz1736tpPP3QlWIVGO/77BLSKEZ+b0paG
3ysR/LVNnHvZc9bKp7lyM7pAsb2RavtBcilNhEDing/3SYm2z62tz+1XxK3AVvo/
ExQzfO6zbCr591bbjr5cdCYWxKB+L6AQNBowpFySkL9NW50hLtEphdzoCTtAlgK3
98KdC70OQWjzTqvsFrTpU8lJqjf7+yzibB9TZWj6Di4k9HiV5ytYH3FSZcnxF+mp
ZS32MBaurXBOTxzTpfKzjceZ23F4ABK0t45bouDLyxQ+IURqoJTcRVT8qg984SBi
PxoFQaiw8S3ANlUwAOEpr+z+tSYenP3oW8PgoT2VEPWHcRpHLjqRNdrdgKQP448i
KvMTwC4EDiwH7t+4Wwfbqzbp6rdnSudSHXvC6rJGpSj5v1KlPE1oYlvxMyPFiSC3
HQzELefEjIEcM2mVTPWk8QbistTkOta0EpMXauae/XURy61DWC1qKUmXT8Ga4dcc
xeHHVGhEtpiiu6ZJK799arv5fh7Cuyg/8U25tZGicJiKGARHC3NxxbtZMrTXj6Xl
OFvtK56bdtwT8U2OSm4OHy7aRKLNtYJA+FftWbn2WtJrJBVMA+rDlkweSxUpA2CI
rea1NPtFQqKnjKvmjhC6LM1E6R8356ICCBhSBxvFW45Pi+EgI1nbBfFvGw7aaGPV
fOKy/yles0rV5yEnKan2LFhKhTm9OVeciXVagtTr13usHiL0j490N9XTohJDZCxu
xzNQFu/9409zRqJbk6TrgjLhOMP5DjoG1HHigGQLYz0wmmyYpWsD2JYJCwyRrmaQ
XiJPmjLu2+AhsYtJafEo80mbRdcWf1qkNQV075btz7X7iE8GdXFKno/5hJ/nAczE
xjfRWl4uy6aBCqlA17sgVlOZM0AmUAnxLoa45AxNk6dnEQBdkPdAybf/X/5y/jwn
dq0R1V7l2pHGE/EnFBWwptvajEuxVvKcpKdRt2FE6W0Nul5SaZ2bqfOcvWFHKXzl
Y6G/F/9CidqESMNitPlPOnFkrxlPTieoWTSraFBSdFcTkqyL+g6bFvhhF0BNxnTY
+y9Sm2PxJsMgadoLRPGhbmfVxWPHZMDMusafN/aXfUl6LFdA6feLKs9a6ZyqwMc4
SeQX2Mhf/GzgQPTzCJ3/qBtG4noIVkaqP6mgHniu8eMlM2gOYInC3BrgoVYZZNUf
7mmqxh3oE8KWOt2bAVrlf+M0oSWloHmbtkXzPSMb23JgrFivHGNbHITdbJDABg0Q
2/2oY65DyiuJgobU/i4fBWivDI9K6O7SNxtItObNiSecjL8TUPI1kL6tOWC2hIpm
oiB8ExWiS+i8p4HAWdc37AxALtqx9w2V8SSgAHhlrEmeyJBSigR9G95kHcGBtdJe
/mGD4J8aQfb5M4+7Hc5WcMTTzbGgpsQmeiC0yMRtwsgMnpwJYAKK+9bPPfqJ6oaJ
YMKxepv27PMrrgajQgkQYNXnbGjFRDoFvpZSmLjgJEl3EQIsdMo8oxj9FJhhcBs4
1xJzYSWru1jmFZCuueS8kmOUSdtVXGKl+gPHD05j+ghODqpirQNPG8dVHPMtqbD7
Unko/aON78QFg5FtYVGNONsABp9LaMnQxB5bIRIKm3SoZKAkuRmNVmF0cvPB5XfA
6nj0FuCvr/A84+t5hYigPy5MYecUgYkwjqBd7j/aUSRbpDNBRN7SCX7j4Zgz1dL0
t4CTTea2HbVbk9IefM4QoKzCyAuB0fpX8ycDFo6CeLT8yBAvDY77rdzDWKICUOc2
zOt727UBxfPBrbfEYpAFNshz1COZeBohPxDhZNnwvYFsW2N3JVSVu9DXTmx5p0wn
jq8PDQukzkf6BYcQzJKWKS283mA+Ejl3kZsMpDwwmpSvmhxOnfFi0OGDyVvU01+X
uFi1+ZkzPE398zKMoc/b4mxNEvISzRs1tuxYBozSCqWnDto39NLgi1ou5w55v4wH
b0a3EUDJh1x9dZSE7ID/Ard2XcNTyg/JLzDX9Mj2IE5cYEQ8e2wxNpXy21d4GRST
Xk0Gon8+XilcDtXu8QMEuz5m39qoKQpu82oHI5w74soFgLOCfLIZME6eKzxRd/Tq
V0czgWJzMw0AH1RyOURV3L/V+JU1HgFUz09SGHb0/X0CbZ5A7bbwYTGTPSm/JHfE
G38rBFtbQhvQwyR5XAr5x7d9STk0zTpuLWqpxymoJuezg2/Wzwh8/xQ1y+5v1EA+
GMTzNOvk90Dg5TyScx0z3Yjec0OSeWE9lVJBohi967EOwAxk8jb84FZOt43HjCbK
QJV0dfZjwBL5roa99lOi4l3gsPpZQ5U0tjKAqSMcSURjzHHjHgSHcGUScZLIdF+y
Axao30lPxLJAKKFldZyO6/dac5Jdn9Ftvq2PmkaaCsNzpERwHWeEQEyBicJ8kX23
QNaYrdfIqT8UBBrMd9v3atNtnZLWGWhpmPq+GGnRq+uVdHI0+8d1a1VZHGOndYwf
jSPTYJryvkkLUc8yPcoMH9PMum1jRonTZm4g+6NU7sGoHv41Rd1GoiJKo69EpN89
jKWJq65ZJ6xr2gLxRw1b4FMfZh9A785m6MahJvCuKk0dI6PSZXovbUdQxTvmUezL
uUbY/2xhr9zpi+pnmDrBHe6yXhjeo/CrL7wdhlbWaIpMTn9U5L3PmrVxn0UJDRmm
qON4x2wDtQAwwjo9gFfA0OUUHlARN+mQW1qTm/eaaEsKRXkSXDRUOcvsx5V5U67d
XeFpuz5rGzFNQW0JGs3lno00YwKooCzQvD6hgUwTTnzgF0c1dRzJCLJjXx2Y9e0c
g+jTc3f23Ax8UmLDmgUJz4TObzcpaGgLMtrmPuWJyNNglMMW//7cJbFgE0DbdzLC
oivNRot+NPInaBIQoZ1i5rjAJUWxKSOj0NbCtJz5GzwipOUDGQFKllxGhwOPnZm5
W/PYprGMzc32+Y1UZlwPjgVRCJmMQxSEJ4CKni87YPtbPj8oRx4w3VztEabNin9y
xflOPwTb7hqnIVFIOtdbr+boTdvT8lpD9ZdeuIgjNKA4OVggZBSK44PcmcCajs/p
paF2RoW/fxeIJCk21hniQq+7CXFrdcYwz6JwDaDMwoOspFMpe7P9ZypKEF0pTiFa
l2kSXbGpZFYe01KP9Kg16o/ps0KvD84NSSSo2ywdoIVrnFNeQ+j4Yba7iQ/CaIuw
WDSAWumxyxf3CX/OUIdqzzYrT1ssngt8w7HR3sDaOAiv6YVI3r5+fXSu/R40FWxw
qVW9c4xfzIaQQ9e3/SsB1o4zT5s1B9PCXWJjuw8b5r63N19Hp9nswmijyvFmHmHn
8OZOvf28RAhQ1Nhw+9eVqvuaqm3RYA83ZvRlSSZUhw00fgpdiDuqzpsEx9lWfsKA
1HKc8jN7/DnlbFIQOClCxYzMA+E6Am3dR8pp0YzhYKEYqBEdHDCrzhqwSXL6Etpp
UeUEIuKSJ8iplfFvWlUCjRmMP2hrTzUrT8JbH+PsoXedLwRxylXl+Z5R2Ojcrilv
KAKVkXFblKKrPw2QpC7EpjnAanHfebfPQmO1+XKGzFnWLcf4SNAFELTzigHnTdD0
2/c4kzCF2DGSVug8GVKq2NUttV+9qvuMQZqLjLKJhYrNlsKz1vpwnVsY16YjvGQo
oYtq/w43xsmRanMYlaJQr3Q5iavfbFEnuj77NAqVofwWJOPX49t6bY6mFJeO1sSl
abxDb2nYdtFl0jYF0w8vECRTvwXaMIz03royQg/70uc=
`protect END_PROTECTED
