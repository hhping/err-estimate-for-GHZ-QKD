`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUc/+yb+qtI2krftSkPwUFrhGK7uUQ7qvWNtY8M6ehBWeVdsGR59XT1Vygr319Xf
8KlB5bzKbF1kYUG6l8Sxlg7ISNP+rLFFLbDlM3wq7eYiWOrd0IFA+f3fQrgkTUaO
YsMv6t3qXZQpp9fVZTNjp/ksq4eA2dv1+0LEWVT4SwKiWVapKrkJOdLw8abzgSfy
VyWTOLdQ15jHkwbjPBTauCbPX/KfCH6ILn76wVxN4FJ8PY2eBzKaR+Zbj845iNXL
b0wh0uOmB2yKi4/mlni9a2eEq0ogoLaTSYVp9MhgERWmmrjjAL7Wekwaz/9sjKXV
xJzkJxrWhUVOi6eA/xEqfmVpdTAbRDAYLmQ9r3fOI/QKipS7pQNQBdbaSOUf2Bmo
LWDpEBJY+LTo5+bi47EZRK1sZUjwG4eRFyh0KFMOVhNHS+IKXJeUfvdaLYpfeMdz
FITaovX06b+IGgV/fpE7gnGFGKVcshAvtYnkh6IDwcD5m3FN6mhIMaUjBGsIBXSh
IgpWuaNnvqMsQ9xLLOD2FjoxDVURUjfnelJm9p8jwH1BgbBxyqU0eZf6RLucUVyx
Y6zNQp7oH/kQwVA9ePJ31WuKfQUBMoiVF6+fXfkCrGMJGy4+Fe9t3GNy4dO/qsfh
IYkgbA56vlvAQCeWFr89boR4vUH+pAuu83xtcIu4G5buNL6Wf/HQF2q1PSXmQv4V
`protect END_PROTECTED
