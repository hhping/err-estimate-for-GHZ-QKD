`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Uj5w3xAWK0P4O0AVf0Fpeyygy1JcaovvI3nI+mS98MXDwTQV3bAcYueR3Yd6d5n
YGJiTZZYtwB0sI0nzC25bJub/Uepk5JB/ivQn2AnmwNW8GBviYMJsTxxNmG6pkXd
q8nMV3+dyq1GsqbsaaHejSF9g6MUVSRYBF8miJt2G3cMnrGgAhlMu8TiW/1c3FCZ
D2xwBUK629H2eAOrvrWNs0D2JR7nbo/l0lMQKfaRTKSXr9D0mMXLkgRNEWZ7ZjBu
555SLzbNUtYJUf+ZCsI1CGT8+kRcjBafdXCcbylsOfn51JhsxD3+9OzyxvWOMFRf
B2+gHdU7/1qsaM7FKK2c+e+mO80HqyLfn0cnBasossSnIanpx+DqC3TnSLyxx6Pz
kW095W97ce9UD5iAn4nkno8alJZqJ9P7dLnnji2dII3PzeidaEWciUsu2eEny9w/
7U8vGUY6JnjF0bgJ3MVC1hDvLXlQos7dvxx2sSZzZT/muRf+wzkzj/us3bDTMY+4
hFcnfGedbZMJSgeeTrRRhcv+W++8uAFJxEvu+/H0DvHGIu2o7QJWDfQSIg1zSHKb
dcWIsC6xcuM8AJbtyQShwx2wXL5sLAvyLuVJ3qVy+XU1I8u4kj5L9rU28d+v6kRZ
FjZH9xr9iPqmEP0NqFLIzrvffUZpUS80UFuJfnYD1EzcL63FwTvYs2cJXPXfrdCq
vWBasx7MkNiA4dVF2JUp08zmHEHqMZHyDZtPKvXDWpwTgpadcdWkJqyU8lrCpuJv
yGibOCF4sj7upVKWE2mXx5v/Ssf51mNahxxfJlEO5PxFFkV/AuGPyuHYuFYWARG6
zJ/+ce6QNcuJ0FgSbr+JwFNYoTLBhA9MTDx0Mi1Sd+1vaV2WeM8iSb2UOnaQkTuA
rbNA6/PTBBINmq6t6MQuZebe+IpdmUAQUuYqSMpvu6nIsK1s6dyNa2Jh66ZlQbfD
ePuooNNXKqeJusnGNODEvqaK0lyVSMBZ7RE/Kt+YvMNhpt1fcWSl68D6FaaOZv9p
qaF0Hcq/MbA5cao9vGURh6ej2kdY69Tcepp72BM6FVbBRK7cwx253L11x/xQko8p
/12a0nWBR37GKATwSthZDwAVtln29OK2eev8lu0CUQzEQRp4Ql95W3o8eWXW/y02
86PM5uSfVBm3SObNQOvhffUVJ36VUYuoRDqDzN6CZ5Q+CWg9qoV09bnnd5z/njON
To6r+QiNA7ShQ3MQwEWClqDGEgkJhKubTBDbsfuOZJFuh818++WYVQsQA7Qn6btX
M5LZZDy30l8LhBQ5nwi0c0s/yCGWUBU2/Cl1oF73VaX6LNY8lpktbgKzl5qWjuyn
uieozBoOn4i3uFN2Z0BjseFAHScdHvJNwMm9D/XgD0DIRjgHWTBKbMB4SvP+6E0b
5mXgftegreM1PFeHn8jE7/sw1SpparB/EHVRSIeJWvA22HHzfPfyWINQ2fgCcoMH
geOMys/bMThob+VJXfSJ4TqT/GlGGYHOt8qZFnwhqehn7qB2qcXjdFd1VrTBJCLh
w0rRpBi5JugGt0YJlpEFDzf0X+Ip4JX2zP9UlC6TvxGWGBtdtV2lI0pxVXinLLat
2ckkJsR6WiamhYIK4VNRWy8bcehvSqWc4fq/AqA+Di9C87OySQ8pmELoDDgzyy03
t/1M8Ze+bPwNSpAZwKPlrqbJXTF7G63nmBW5zseSrgb1w6KYcJ51rUGASvg7PO5I
n8nkzmvM/wezY5Mky8E7EMaf7wA6aFnSTqXjpJEViFHML7inpxFhCcvaS/iVipF7
3U+7qNFuWJb4HUMUpMaKb9ZOe3P6JWUlsBzCNsQUFMFpou3dUXx/aZnqOcgP+yu4
CmBTK1o3m/gD5vU0ZFthpf3ArU3eK+4CX7vNP9VBg2CPmtLHUsWXHdZNb5DrChTJ
wKoPF6iZwb0mbB4dH81FYyY4jvXen7Ia0u/PxMjOAMgHB2M7pROFcj/uKoauYqW0
Dqv8jNy61CSvaykT5MWogfrZG6TZVoRx5HQge0+RZZvQVLZUwDmL6jrs7CZdUlSv
o6838sGak4jIN1aY47J0+5YvbXQPT119oL/6xpiKDnLVgQoqyXY6pi2bT12V5PEY
jyDoGMGSbGCn+yhTtHjuLm/1YnMqn16KnXys1O6hy2dudEw+yo2Md7pDOOOMc2EN
A5j09/Ic5Kcc8a30jy5s9I/PWI95UEcKqVkA0eNm7T/nBzCBAAGntom3WZvoIajZ
GpcYcPetB/ooHFpxzy9bD51OD5myLMyTckGgdjoCNek2PuWuZSb4lv10sUupx2N1
tZ5ByE0WF6LAWOrA8tsEOSkwa54WXWhT4GTWCwYBfGJDXrmHBukbX4r/Yl4ze7ib
lDe8GRJd0Mzt6IpOi6qUnxaFiTW2YNrh/GVKmNDf5UsqnEBTi/AxqkY98cTOy4NW
BENU//Z4PGUw3epBjXFelluu6Iaaq5jYPBQ/apPLIAzefBLcWWfDcoZPHiU7dksA
j6XBxeyyMGD7WQ6Pf3bWpXZVu8RzkokU//EHfyHPlFvQWETnwrQSyjxqxu5Y9sCt
HkJijNuIqxxkVsSKPQWhdTK+ldG4wB8dqCfPVqKMbmnTDAXyJlIADinGgBeHKkZy
CgNmLPMX7Gd5SKoYXDing9Ar+oDD0lsNQE3kd+8r7N1X5Zhb5o2CzVhnXwRbl8NY
wVh/eHJoOmamgI4CdulpUJDHpouFAvLp2hHY8lNalZit668ahq4V/e0x4DXJuH/x
Z4Bs44oXIFID2hcMRN1vvjNBVxxThyRm6VXLoepzzxGB8KnLBBHe5Yin8HmsRTiL
fJNOqV8wYBasmiuyFTmFqv61QrlEgxXDZhIdBmMcDy/EM5BglQK7jzinw0taSBFw
ghIYsz+ON+tohzI2ge3riL4muQfjMZlXnYZyFFLh+UF3C4D//PB3o0bROK+AajgI
C7x5pF9qw4CXKp/6ORB43Bpe/WNwbenXVVjH4kDBJT0=
`protect END_PROTECTED
