`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7r39lfVRjuE26lYbaq40r2rS/EUsgLgu6q8UhsH/scjakUmeiXIQYIoKQe5dDUtG
Ey8d78XZquw0u0lziUN3/tKadUAgtsx6P5lmyVksyXWkHdIUXU/4oOkiS/483Med
UHID8/VdtaZJ4ILugtEIeWunAJi6287gD2eWF0LbGHsdhLagebGiGGV7ZNp0hNV2
D/EE7FLYoMpLfxR9VF8s9e1Tj7stNA2NT0M0+TteN6ZGnDDlCpvOFsntwlmgRm3z
uwncxIija+tgMFgCur/vGym5jqhRS+iLhx+cVDBqe05U4cQxDe4EeJU2s8FH3klK
ltnGEWJvaCBzyjUuM8IFRAzjo9OFkbqvmKGLxaNcL0J7cBnM9cwp6dsZYpcX+zf8
x9ROXoglhJTeN4AapNMdiEba4w5+9P3GdVCa3Gd1+VZ0fFS9hr4+MZyiRqu2eYBm
9pLz5hVK8TeDBZ9r3Snxw7iwlDLODZ5n6CSMPdC17RJqSH3DK7xOSCUJzLPj2xl2
I5fWHI2W5EYfHobGKRiygZcQfdCBc681O82M7zE0PbZQr2dWvaqrmRJb0hbxlytA
M2GH3Z154DLededIRzNaBCDpZFcCvGSfNDg/lK1cMCVKcpd+freuWKCQnKDE3l19
66QEro+RX+bCkGyplLvTAMt2nm12MFjBXLSNtwhq7195JzU7S9JURqma0sYvf8bx
LqsMNvqrXOC3UvlO2qS0vLFy/BP+AGXMLVUyvDIQhUPrqaBqkjO0R7oFGNsYr+2c
7ptM3w8x09gRWu9W/C81UNuhZued9uhlAJip6NofLECjm6OHDD2m3ztq23q/D7u2
kyz8jUxv9ClLvt60rS9RoIviwIoCIHLEHlV4eayoKkw31ZnEuNwUdWuZAmlrR55R
dGwo/XF3RM6CUbSQqMRcB0tKjb9cgNkfkvOWVqJjM23ZpL2lBeAPGGWP42so2weD
LICq1IOFhVe4OY8//C2aiGO8VCeRb7XnkMJImzH5kJ5XQb1lAm3IzFk/ogqWv2pY
wNCqSKjmAd7EZ0jTQL10xHwtU0am1F2fm6icJnN7fbI72ofKcD3RYjAiVJVLhvZC
ZBNeCGX1x1JvPie6eYIKx+0QEDLNmmTFau3hWAYvmc/SFU8iv/9MpnRqyJ4xdU7m
McJhJ5ZhJ8HFv/WpNH6SvjxbD1/RuEzfAyZ2E6T4N6lhpcxhdx5dwHzQY3ZeztQj
kizy9EoRJ9H1Fu/gpvOJnUIVpGtRL3srJwISLosOkwt+19lH6tlG///Fw4WARluD
GMde/d/dock+DIjoe/cUMdFbseiLk7b4JrdKjAeBveW7PjXLkOI3rnCOY/P5K+sx
O+vpucp//NzOWWorWC1KIsHRld4nrANTphZXqE4sAxzEMwWN0vtc67xnGae5Y3jk
KUH25HhSAV3FJlmtW/0PbdNlyDL4fvrPX/6e3XS7URb9ueKt8CcHcezVvbuQtxQS
TaZMtIjekXKXhrN5hSATeecGh4Kzwu9ovJQLsVBI5ye5nKxDizeUNNZtYsG2JvDI
S9koclALe7ZwKGTATSeznzCaECF4LNZVTrz8vD4gscdk9GMqTehB4/MczKxA4vzd
I3fIuSK7xO2xqztpCf2Ex2TMOahPSqUlK8NUdR0+i4T0fAamqNLcEwYWmqBvnJ7B
S1fSUgas4hLPI2jFnDT4nTIk6k66WhYSgsqp3JKfAQhZRAytzzOb2ylNLEi4eoEc
93319n9N4aRCVLVcWNx2m9A+5qACEBmEycEDBr/pxauAruA9uiIsnNHZoRnBIpPG
Hn+vkE1DmMSquSQmXhDYPUZ6IUTiJeFmZrfmgLkfhLDbdn073Ldl3AYBrVHU25mj
FI8vGWDMYKX0nBEo6WXxPW8+1v1F0bGrgBamFS/5O9BPNnhs2suadxB+0oDSTz2w
aI25sbfsUA41rUAmw43kDnv6YlCqVrCpdT2PijGqhMjLTbckU1WGqDN0BCaONQlZ
m6XvRSxpTbzX8M9HrLEj7yQJ6fELfDi/PAKLsck/0QHdX+aYVHuWsIZZTwVRfUZM
V0Bu5LBjxaPyfNmKr3fJ3X2l5ffff/yP87dluHS9veR3fT1x3x/fEq92XsrAdKWq
JPWBCCKHsbQYQyasZ3PzHQQaTRgBKCjRJ0/nxpG0btVfziz33dDztadN6ED02PWO
7GVx2pMc46Br0BOKMxEbgg+PtSgBv7bnsz3ncN0Ix31s7HX4pxck3X5Lx6eJzVWl
K6Q3xOOQajM821dP86etvGjmd+WiqlPKJVJYsgLsTxHIGGfTryQQvtvCK2EcxXIn
cqaoeww/9quYKjOFtxDCoTrC8+O2lnxGn7TcdM03YwR7ITdtXzJoWDYl8pFK4kDS
/1q/dggIXDkR0MpLl5P1hIdN1L/GjCUpB2+MHnMBbgxywnN+SOzR6fyVdGKEEP1E
XvvqiOWB24HLdIUFrk6DDCmBU0h44DAbe2r1Fgxrmh+8AkYq1LrQXGX+yssUISxd
TgZffsvtlpZ38vHS0SfoBNcp+M/KmodVwr1xP3VgEeHHqZPvWNUxTFTGdrgqWMS1
9eizzfS9uM5nDmBM4GTHQ/WN2yQmo5a1JW76yp8NjO8sqT5MuRxbopX9/G4/D5D5
MKa7fmLkbkdYGPc4FrRj2kPDVLM23lX/lgs1zAkNyNtGkafD/sV27NeGpe9NoYrx
NJOVr/a923WKZTrpzInUq/XbrNpd7Dlb09brrwQpEzBwCgmP/ps1HlXndEQwLSNl
pVkhZlkpvlvZwn8SUv6ZpJa2ejy5S1tIVieUK3OmSNRoYDVq2iudf0tgxBrK/4v+
9a4HYEwUdh+LQA6TtepgktQMp6S/xai1aH6OqFUr/mpDMTTrREVBBX4nDDT62fFb
xRizPi7Za8eohCRt3sJf2m+Vn0F/LShSk81P58Wj0/W5xwkjagvsuNTctJNwufhp
SZRbDYFwm88MZnS/94awpp7x3sAaY6iT5IwXrpCw3uN6kijOJGVzQQ3hs0+MG5Y0
J+YKBv52+gY3NYIuUVJZRY2lH49ztarhOyuYlnKYaTvxROqUPP+8Fp1tfo/kXEHR
MMVZnOnhtJSKagP0lI71ovlPpj4UhGnSxzv8ggxnaZQvmO3fCr4P/6enZkrKgslW
WwbfknStMo24ctp+YwC5Umx3VUV7+naDuLr1xGS+Wj+1H1GmTYjHyHmZQSYuBds4
wlPlIfnfQkIrRzTPXx2o4c5lUfqVIJWWD8fM5UmBXT8W/N6cL6v+IFmhThJaOOFx
7rZITXjhXuWWnnc4Ao2xhAke9RdcxeN1GEiIZWk+GLaTtKLSCLFXTpfLSuuEtaym
7YghczqnHIflMGNGHSVBMw1cv7kt5pmfEDvVz6i64rI0Uk4F+k+Wbtay9osBo4jv
rqR4084wVX0HJuKHpprKACMxBW5BaERYn3XsV1ENZtToUFE5q8Ik430aHrYqJwSX
yt7V5gbpwrQjy8piLOgbZbpbdJ+oVY/9oOrzZ/KqBXuJKy3UglDpO9ciUuOXZhAB
fnrsXIojJEcdgw/aEdX+zc9igArMbUuFZAQHdtba9UGrlLg3jHyCtyJZcvnU4GfX
LfbKd69TS1TBOCUNIVN2RaL2+V5sDkOMu1jsEQnfJW4FIwYiWAcb3PCkkOgl0DhI
9tjQ49blxf0iFJ6A8CUPQ8YRjJZHe6Zs0VPFJPgiqr+Y58J0H3UcZppZHcM6Pe5A
6NBNoiLx7/kBbAjEsN8bNFTf58HR4fAx15jatq8JHavjbTZoRuoYzo1vzuEb/GKl
xYgcJErfSUbzU5zrb3mZEvKAk0+7YBwf2WfJ/n9lbxxRPMwTAnAfniEAcneuUtFN
3hkYeIVo0qK4auDbLGRim7adyKCiL2BU0EuAI4ty4CBRpq9sr4BIM0Py32mNzlhy
WaRe26a+ifUl8YpV0hn5MxSmcEg0XqX5VfB9Zo29jbjlBl/IUgT4eYDACehqHnNG
OFxNEvhTs9izy3hYl8U2b/pQWTaKMGiUFobevF2IZ4yBkBqP0drHqax+jUCzGUay
SOA+YH9NH+B3VzkenNfhOSNnG8OCL5h+frVqYZkYlKx4H8A7p8AMDNKiE9pgX3S8
IltYKnods2Ev0y/3R7d/iVLyKiKQbEFJbRqwQUQ44ZCZWy+gjlnFT0jDz6U2W7hk
72S1mRZPKPuWbljPnSWo7iM+ZggKAQetI3DUi65LoX53tvj5ddrQcw7UYMeO+GCW
IU8hgCKoxegCDQWE3xz3zvEozuYRcTg5NuXptLbIWHPGY1s0MTfZycQaC0onIr18
AMdrN8UEx3I9j170qsE9YWMbc1e7VAj+yAGm3uuM8VP0K/3oUBF02+9WVHVOPNyT
AxZRTBlNjYQ+5tBc7rkDP+7bm8A04QdmvAGUfaATpBq9r3pGMclWxD/+tJZSMkZO
UDAeN0/Oejuh6uC0pG4FRuP26SUoebOBjDE/YAI46rE3JLChWOM2NC35fJ1tvEfd
TaIbNAWU7xu492nZJ3s9lrKY1fRNBQ/KjoaZbnngWDvuRsAtxxJm1Qnoz2zsMUYT
I86wgGeckQ9ROB/IgnO3Lj2gZ2hULkAeh2qU7nbcS9XPfCoYkBVit1NSWrp2lFDS
uLQyrJ8+4FdkpiK5WNXaJo+De3e9nWoOWH4t6/CYCIgckdvb68eWVzhYmJqXpsTB
BBb+63OCE+mQCGAUZvsAsL2OHOH9Y48mC/ipk0gLCxksvZYwYO4RtxbMmpIU/TOi
LDopyKq0uJan+WDB4gSlYfjchRkmTwySH6hPgYGZWW0EALiaPvCd9cEmt0TWRDxm
nipDzWaHoNCmA3oZB1rx10+azn5jz5Cypy7sG5yMahgm3NWyiaSFBHvXWYDf8C9Z
Rp8Xmazs7HLRH44xUvW7QyjE7qHeTsTgQsxKm4hH2Yg5epvOuZsFTxUc+Z1ZGQ4k
Lfe7gROq/EhRO7Gmbc4h3N/8gjIgyxkhk+p8UetVtzzsSMiUIaxASoIGXh5aXTC2
fcAcDoajOGNSHNConwkXU/bI2HDxFzxYv3/9T6xnsP9ErIZcH/ixawruZDK4tN+e
TvS66XtnR7aFvVPJjLAoMgjRX+xn6rSFu7A/tMhEuyZff49mGPG1XkupOWyc9nvY
TWu7krkMnHSJ0XMrhKknN/8XV1DSBIH+1G7TNPjPgn/4oWaYJujtt39mq5foDDRs
b1m58JTpys7qobVvKRMa9xfSujagyH+7anQjXEbNmSYpMVPefGWQOvDKxAAZo3fa
NgAkCtxmNGgQK6AFbAemC3RcOf8u7Kv+TFkEGfMoDoO5ZFgrdrCcvARdo/V/M2m+
dIXPZJTMBAaedVOXLoHZAvOWFCVsOotCwI2Yvv7MHPXlQ6J6F7XSydruaoBRZobp
SmuxammEgY9/rVCH4kNrwKBe3SeQbzQ+h1P2UauJw3/v9gLxERUv+RagA1VffuTH
wxUhzllzuimFUMlwAuurCxZc656kyYRCY4KOTwrtXK+8BF1s7oPGzUj6oujaM1Vk
XBi12quPgfbNo/QJjpsAoi7JKzyy3LzTDvjswRTnUB3Y/1opFOjn2vr+zjqUaK+y
UsbRbShUaj19YNHAym+rJcYNgy6yr/sOlSSCNgu1v+D1jKXAXA27hPpwQKii3zzq
ynp5PpQkwEOg1Vi9Oh4/jDmR3y/HVqpsG76hx+VqOO208a2e6swsmUIEOOyufswe
QJT1vyovleNSf/tTs3RW3+6aIobIuZT5QVJVNoNCp3xRWNIiy3f0IIlClFpq768R
+ex+vCug2P3eVONfndsFAdPq9q89gTcP+lev8L8Jp33FscCgNUhYr22feGpK5PqR
ncshlcy4SG1NK4b3UMbCxLJeVmS581dmuDLvPpZHzZN1xzoUFXMMtEc2HOUzB1bn
eHN99LAUzAeuBfMrIDHIXo1UT/PKc/fijaG0/ZXKzNTWN1UOxicFRQzV1cZ+DGwk
OLgHHNoAgOryxY1ssyogQrz8tYTmcsMdcAV3Dju9Z+DSO8n0CnClosuWKtFowFKi
r1Y342ISA5JLZ8hkDRkelsYnEx5Nw5xMnr6oKfia+EM6Vb3qkOSpAaQPjHP4SSUG
wRT6W7aRAXnBJqj1NjjYTw==
`protect END_PROTECTED
