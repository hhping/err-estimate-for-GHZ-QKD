`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9AI+uZkqcJh9oe+0+VYXp1Xnc4rpnP7DAGhP86J5B2S7Pt+CITVqOmneWkJlFlGA
df73HEDVYjftaPCBogTrn4e99+VPCHQfxvFMw7JYh8WKihxUjqtzXSApIBEOnsJW
Rd4GRJkApODfRxabI9mT8XftDORQb+jJMXSgpFkj8QjMq8V66ccYICtKkzlMwiVq
u406uZ8OW8ZwOGF1gaWVozDawGSCRHS7zeNoYoMUi9rskvagOK4rGGW7PyqPredP
EbH6I0T1Q4rH1UaON9G5BnS9mzR6nX9T98IXMHPDBlJrwF9K1zR7wfw2faIBmOXB
wLyVbkdHK+VP7JYVuCn6tCWMXKW0Q7d5L05dJZZOJliv734RQcC//VQHrIzStIko
abevn5WBEWXoIXrbpaVOqBG2NkYyW6Eoli84ge5y0Wqi0F/KvLI3/jWhJdO2c2om
VLp6VpjJAM9kgiz16Bc24ofFRQhh+w1cLmufVaCGzdjLDliqkFHG+n5LBHKzoAc6
wg1ldotkxmiYY4XfMCBOEv8WP+IMxZw7FSKgJ9gCs7MPasgO46ue+q1+CrSlGm0l
x8nSExKeaSyB6NxhT0A/x8owoNaNyG9ISglp40wquthXDj3hq6bUl2J70pe211mi
D6KPhPiKCoFALPEykX+pPE8TRzHqdI22HMrAeBLL2V9xs2GFVOzAVxLGIqF2VbVf
q2maSG6WSjG5RtAJwmsNDAYiBEvximhyDc/mtd1jCdP4DQ3ht1A0W8rg0x5zNhxY
UCK0kPVkzq1jBQ+9ZsZLP57N0/LtpeplwKb0LmveHCSsw9lkBw5OCbxGuiaSHzAk
yAut+0BPn5EMuHC241qSfhhhM+CPnuXywRPvAjlKsnDFssoEqq+4jd+zpOFJs66E
OQGYLtycONxaGX6PR35aUUIq5scCJ7QyMdKFU3ykAet7u8mhLGp2uP1XnegEMiI1
9NJ5G57uR12gskynNGldqgBSiSCQpTfa5FXgcCklVffYbqYH2VyvVe2mN31dGTnk
Gd3Psd803FOeZAkB+WR1NxzJlyNQ+RRu2MiM2qaBDOxQW5uRTKf/2ISoW3h6McIO
Gf5Hc57vMJGwaXMpPz7XdI9xsKT90DBRnww4VkWYeK8W0KRlvME6bmscfrPpczrg
4UO56sHtOTJQaj/sl4brJdssrDuE6kB4gzhuArJr9R4HbaOvh5MFqCAmbgdFMBpj
/f6NCMc0al8DnglIkTgUdZBrxnsGl6Nrk3xpLXcwCF9OsZ8S50PTZiGgWXtsTvQN
xEMv5C7maJXe4cqaUhRFSq/tH05gfW3YmCNg9lt3wKJMdmTj0rME5T3CM9elYdcr
HoXn8mOCq3aQKWUR3bSyB60xQ2eBHVaSikVYgUDzEXYqwtHCJitCt+PUzJoRAi7Y
gnw47vAmTDeIYWFCbfUCJ1GPVtlhbvY89GiStnQGI6FPAcIw+Uu6g7h3M9LupQIt
U575/+cHMavbPLmx0CWMK3dfgG+8dcy0LdxvxJ0rCE5WKqv3Rjg0SUcTu5IbBpxG
J8Q4ep9yTOEM79tE2qAzzZu9kEjXvY/5bycgo8KN91bD9perLsnJazdAKwzP5Hqq
jarzbVfdRyC8ve1mnJkRX57zclVivFZf+ABkap645BtVcA47z4nCC3PupteZs0MF
16IFj8xlQTiMuejHimA0+fbbA4BVVPO5nDOYyxxg90R9FCdFgE9/0myDTg0sF4y5
N11U0FTI20YRLP20AiAlOU958rsE2wLDPa28WLethzY0eApbfgC+sYEvrmYf1n4D
LUzMtvI9re1f3xYnJUka2PyRbQGvuJWaRKyO1M0oBWQ35PwcMu2LbWnUTf55sTWh
5/kxk5JWBtEBSZou4C6gA+c1Nzfy9P1TOntJYdn0ldp2Lo4l9NJ2yEUvnN5aQicF
vscPP+MMErgHmhTSASYV4YSJ7gVYaG2+4zGbGPFcwOqy10fsz2iYQ4h3bRYh7KAq
Bw5K4QI4TB+xK9Za8drOld4LYwmUrVC+//huGr0GYbTa4V+AcO1LxEwAtdRXoSx6
tbofiR4HZV/DNMS55YkZzYFdIqql4zuYX3t5Cn8KgzHdL/p0M9HFQcrQLK2SC2pL
ePuDJ6dMYVVEQOGQcGVQuq4nE6P268v/U1c52g/oGVD/AOLeZ86BeJMO2FMlpM2C
p58iib13ywtG/+Spzc/9z4GzqLvgtpSjirsCUDfjbXA0jWOj4ACQ18sx7JeUHYFX
GCbNm4O5m5X8cigIOhtVDELYUnmk4Bt17hzarp1vNZukQMhAnk2jh2KbiuUEQ4ay
KcxdPzyq3OcztBNE1HTXCYhi54jGM1i4e5dA/+1lXuJQ8g8nSMiLlXgi7+gJZO9+
Rqnjw4wYxKdqfDpdYgor+QuwtaYsTpz8W8TiCLHTIFGVDkuLIdRPCoGBSVVnHi1M
M1ZrVi0zSDHNvwAdwYNp70NJxhXmJXRuyep/kHqbsfc0Q1jrf3XCrObHuVRarDP6
H8apolyltbAmO5bK7zAp+eW+IpWvnYf7/GcCz47B0qo9V7qmLPnPOaJvEf5/d88P
07HQP3DQpWxtf+dwdB/PmnBrp4qCcKvWcfsnyzE2/cvhk1NNpdt79EGWj/PjbLQU
lL5WoWAFtbetWYpwD+FzTua/EMQ9vUB+9pZUNh98BKCcwiyrG+RDZ73K4LOnHuqN
RUttGzJCxh6Epv6YuhNd3Ap7lyvb9yOOOr3CGvCpEfF0iLedYItvQ2B0A0dQnxxv
vWjMz43EdWuuSfp3OGs43ciBCGROGpeMcurFf1qz1KKJhqn3i2g4gAY1Z1QUocna
kXhBe7RLDLriGzrTK1n7iRYFzzRaF0D8k3485QvK1MNEoMicShakhtBwVJGqCb/A
v2CZY8D3NgT33OFpktHb+NqXw3zJ+ugTCD0DT7XeznAEDMoMedszbreS5AlJcvDy
e7ZL2Nr+mRHhOTVENM3dYcpRd5mWCIlamYp9XGgpXW/x8mkPjN+G8rVdArirnwFr
+i840vh0u/5uD2xBWxMtcvz0iANBHkmXHxOkXssDj8ni7j7XUGcAFgHscm18Q4Qx
s7R77a3Wc7JvzN8V7afVYE2BHM+nnP7nPWzeGXfPYBM2MvyjB3jPRocpjzqXekXC
6fLr8G+kXhR+LFIkQYMMdWTFwd6PSanZzT+zZPCRMtmT+BHObGKrEtuEfIhUE7EY
h/a8VkyeanETXu/znhTSwS8eKDIYZY0AgFYXmuIt2v8saA2fYiURZqmYfbMydQhr
9Z4A15qvXqnxPWfC4TP/FRsRXOZuXch3qx7/5+MveMSNJi4x4DbLfLSv586Qv3mE
AXuBGiqg1UATt7yMfsqzgRFF4+uw2TRlSNzC4LaqtaLXbk427qf/gOBA9Rj74671
0BaLk2VocesQtObwPZbMbrF9WkLm2UJikLRKTstACiyyjkm6og8H7u/GOtRsz+4s
iAejwcCgQOuzW6A5vBltvxw2+C43pRrI/PiZEx1+FbYdDv1dykIx6OC/71rGYWr6
b5vGU+2qkAEh+mNqKVOuo3fxlQLWv9hC5CrLUXZewrLdCnAmV9vbadchn5PLtAkh
MRqMOYYl2/AVO9LL/E4Mb1Fy7LjBcJ558QGiEcwcxcCXWhoE1qFq++4eOeozsno4
6hMszhbSN3EdjVKtoKrhSAN7CJVwMvxPgtuDI2jUTJQE4E187HiFvmq8i40vXQ2b
zs7R04ii1bSBKd4+wGd2MWK/cpqK8UbzRd4BYKd3K52+y9AnMtRBwIVBnnbpp3Km
KR96hUH8hTdR70bMnE+8+2XXWpO2sOlNB2lWvX8G/tQkpnI5uTP3Veqf3lMvJ/2I
LR+ANBpgZJo0b+lMDtgPWPTZsVBOYfWhMTPez1Kto3mgMc84odSM1PFdPIbaq4rl
/eZUhYXY3OdMZVVrDGP0p5bYGcBQlbQcpqg7leStWn4fd7viugcsiXCTvq369Be2
QqbHqrTTdV9hajaCTLi/9q4gXerAJEH+MzXea9o5Q9NM8o8vIY5H2sw8dpsWo1LD
8WnyHT2OULdjtSulICTS5oYp8B60DHPK36q9RG4J936nj3t+RKmI2ueEtR0cKMhI
KDxVe9MOikzLVtBQUly7jyMyW1Oy8Wp0I/6Zkk5F3/OfCpdXMx5woEnNIOX0dww6
50c50g7pWsk7IfqF2AuzMPnW/r6+o80HYufKGjl5OCtXrdWO9AjEB2qbQ3TG492a
LcRipFd2Vf2cZub2JBG88RWnx61EPh+clffXNvz2n2Hy88HPNgottqnExv1Q11Ee
3H/UFa9yZkMnw9/ko+6sbfuHdi5nokkHqH6SgTg/BpvJ1FmdA4cBQnZaf2PS9eQJ
fLmz7pJjeKLj5wURvwqt7x7qF4h8v6wiTSrAsnjTqCAQZDYFtOsLcF0lA2VFOmA2
R29XmUmjUtK5Oz2w/NM39zdQ8CT9kQ3rXTt8JHJWawtHeR3xHYYN/jN0CddOxszd
SeFFQ2IqF7pzr6DNc5Rxs+fc9/QPUcwAWJp6fSlrxUNjGm3IbyZF9wFDiBb61UF3
r4GaVJo9ZRpIxbChs1j7wrkA0QG/CJy3O8uaptfnIJjjMxVLOXKiUbU7IhyB9cbd
dQ0nY04TSMKkyiq0Y48+Fekz+B5RQIhkyqd+qJ+YAysVEHiQFsXlSDmKlOdtUtJI
6CgypmjJH7mHikUeezwrJJEzktqHbprT5/XJ4tiimYqDuOLB6NmSsbZpsSPUQjaS
WPuqhjF6Hea6zgyrOqRgmdxkb/acHoCa9ro+8JAI2rIWmdYPLwbe7hbRcLvvWL2o
KWo09ZkLZmxB+IGTghNKcmG5AiL7brOumJJrHDurSJTZlVRkv+iJiPyIpeAPGI8F
doD94YSUZ4m6mZKdn9Znpi4qcScU9YLsDbWuPHMmQLHGyoFE6BFOpU3JiGneJX/f
BCGCL9PJsr05ZkKj/g9ea2GtZX17SLNLmKdhmv7sQJwskjCt+7r8DDG2x1vQEgpj
t69sH9WYN3mAaniiWvDttZGlOnNMsCgxtFCO+hRRM6/y7e7Y9+tTk3/9Mrbf0iaa
uTNIwxZLz/9+eb+4MM/VVGCJPeSOv99eiQwmS61CCxUfUeFxSzQS3UOYgs0qOEfW
3SS+ZE4KpsSEWT0uxDDGR8qZHcsG+p+gvXIOMVto+Cx5VqwMfS1gIdqVw21nN4X+
9iX2o8SsJ5X3WwEN16DTTCuz3A/N4/CboBrHRnD91PWibSdYbXCDMpsE4VeMlzMI
bWBKjCUGdk+y0KZiFSH/CglTX6dGWqJDAxC6goIbRtTdHQHNeis0Pwpsb+gvQMoj
O9D6PCE/8OnnSpD+me3dQf6MoSQ5AbSaB9HVxnMUKaE1OY086B5FN0Yv6hQR5Db5
cXcjbU6nojTlAuOVsdOYZQF/8i6Ld9JC41QUV5FDQ550Sl7fTbUUizXaY7M30Keu
9xwLwtNESd0fYOIHo48jqBusQe6CzOiDOJyQn5M8XiZf7tEicWw8jxf8CuwigRBH
lWHFYgObYNx+wDkjVues/INcsTFm8/2xK3eLCBjsLVHAfnnUvxVHYXWv7lrfQOYr
K1f6iRpttiZe8yXI3uxkd371UKvxD+PtugjAyIWH5E063x/3vES8KMP9cgLIyK8D
3S+piBrXOV+YIXLvGq7n7X1BnYe2Bn4ldYIHIiG5mUID7fhl7W69/posbEQOvfA6
+MFnnfOnVI/suZ+ZF6yIM/pFItGg1Yv0A6V+eY1oVtF5/8rVnBTMZjy2872QwMxs
uXa90jXeuDgqPDMwvvZvZbUTqLsSHaF5SXgIKdSIUpdubfqf9zOauTc5cyqhsBZY
l3gxTs0kKqcVbyJf8j7HD76q4Evr9UWIYNNpZFb8imY5OsOeD69CJKQNqVqanL+i
CqabuhEbnpryBZML5ab0bIdh7hXEFSoVW23unwzC9NCpFfMDrTNwe6Qind1cIsgM
9hML7LCfoktS83lD1QgIUCGVGZt8hGRM44KAWq0uqXix2/l5EkSLhkP4mdSrK0cs
qpUSq43VwbZtkZEnFMPQ7BRbQ7wtSFuk8VGNS/4naLVXrGmc02xcERcX9G7iW8NX
46rlPxFc8evje8yeoDcb4NGigN0/io41SrvgKEZaGSw3SW+gsjvGcXawnEuw71xj
Nr7jgv+J6VmEXnf9qkrs+9alt/TwU4Iyz2OlP9tq9UO9dToQB5Bw/YU8OdxBQnBC
mP+zA3zTGt/R5pe513sONgQ5BRxOTfuePkbQplpj1q9irbMUZgsQyc00s9uAOrlh
itASnThfDGfs56+hhZG2o2GUZUQnb0b7+oBFtpWJ7y6asqwY47xeOox8aIRKdUA+
zYT73CS5/9JP06UNHnVCA/pIde3AYGjK8OEq0VdSgyRYjSr1wc5TiLfK7Tca7afV
JGzDO0XFydehbc52yCelqitmScQXAlcEbSL9zPaRXl5gP3oDs2xv64ngrs+VHr/H
yjmwWgr6CArUiYRTX+E5TKMbQWEV4ypev7iBi6PDKZ7PHewjeWuM5+P6xKUl+58l
37D9KGRzSCwCKjDrQXcZAz5vjKyPo5oW37V1aeGMw2TspndwL2rHi0YV2Vx/tTVu
cKpfDaeifSgc+CovMMBofJJoBs0RuqfSzFmFdhqRWFI2CaScComUdpmsUY6gnBMz
NEoNij+TLz3Mc726MZRefx6nQbTWkmsmjgOfadTy43wfeLNgIB5UAEXTMyue8dQF
L5z1E6wXPmfqIlyLsJWGQGCG1xpeHPe31Z/QlHRhPhzckTlsVoDDiJ90pGCgfbk3
kZLEjXqV6GkWW+P/zh13hF6KYghFD2Ed5ISWTROrMrtcL/wCj0AY0ujPS/7ihZZe
7nDLg7QyxFltARbRjeGqhS1QDDRCnGy7hb1VM1ETK1ld4QOl9Tpdx/TigIHvnMHD
JhMSU6K3s+0mTZYSi6u/sLbnvTUKu9VVBZbjid4owDUUOYVA7Gb/+HxKCtMAEoH+
9JcX0HnzwR5KqhnFc2APGHZce8E0OWEiHgZq1UO7xiPrrM3ETcWdYAldKYYxpqfH
IZKtsHp8PAWaZSco78n+imfQDUoqUK4IMQColdqSXkdgVffBkusl6/VNg2keqrSy
5uTqmaNjEQv1Ne5Ydwrotq1/+tRwr0s80OwCvHnMIyqaL1Wgj22KQqJ0SQq2cx3u
EYEwkbDYIkqZGSy2KB3lYyk7LxQ2gVYS8hiHscI+2/VpRg8E2KJw8k/TiHvV2f3S
95EqGkdC/yYPGfVqDpr4sjDTQ8F0S6UCNBfh5L3d6uwxOyU9dQrbBvMrgN8Qz+zb
rdzFRGo8qApFi+SSv3VvQoSrncDeSIekiUAuLQzJnOqbyleVVhbWZ6h/RBkzUJlS
T9tPdsClvhO+Up/SVAeQ+ePhv2fNRDsZJMk4FhjGhEOjdoN4v4Ile5rSUpvspC+d
QqY/O7r1Z8P1UxphjYlJmrsyOq5WqXsj2JnpYLNOzuXomv/qpfv4Q2RniHtrV9Jy
uH3VNf7CwgcR/n392imR8pMTeJvQkk2zuvl7nPzJrVjVIyb+RkAyV+nYNNwVRe5Y
S9zuhej2w0Z4wq4PF4wTazwGT9P6VZAZ1VRSXDE8/ccKkUpJlcd6bvPetatNGXFQ
lWfcLgTNrjDvhxwzADSK8vJ7mDRW4wgmWgWYf+aAoLfRsUelSsNoIyPQGDtUS3Gq
JzjxOeQ9paIZsnsLodPBKBsovrlPlzWB7spgjlt57gsT1M/A9zaxdj7RxDRlu9v3
+pWAzOY7U8Zou1+8re4TwKFmOyK/n/cE1SgLc/3bnLUa7k92vLbmoa0nkLp4EGLl
4vGNyO06yQ4FuQbvnFtCLOQO4Zt4pZdf8NK10Uc8BmtivIcQ3QWI3R3hBQCWxSfC
4C/ThrbB7eaLnQ+GpY0sqoDPUP+BOd2bZUuar2g4/rHhdKDMmK4lhtdCYjTsCkCi
yHc3x5z/dqCw9eDr7pAb0nvIAMAPjPRZq84kntYukuFLZcsGgasUP9MhSPdoV5Id
4UvkV0B7pKQRj1ZxSqDKYa7jB1u7OQqDuDatPn1Ht5wnyGAXU/LUgTiNpoWXpv7b
m3gMSvApibRgW8mLZ6d/khPoAp83n8rt/Zm5br1fWz8UC8eH4OYTXlzkD2fHmEkQ
ZgNuC1wA62yBbq3s054I3J4bMPfv6pzpWxqkFcbkxS1tKloT8rkz1+Uecd0Jxaid
huj/yIpGGPaq9yRMVLjw6n1vjezLHN87ZVj9srYk3P8/1VAyk+jAP+2fpZ/URRxW
vAwxMpoVUzA/fYvpKQvTK+//I85eK0nblmr9vKW12eSUa1sfnGsZcDlo66adXBp3
AoADXluMtYN52XosQuPtiJTpnUD0NsvlBoI7NonFEsut9gsEMcZeE986yfE+HB51
PiIMfLKYLNasSWfsnmAn6g0t2psq+XM0cA+RZneZElIbkJUJ1RkFd2Lu10q3gUdx
fwixkOynLxD7TIIFNpHomhJ/xz7rwtiBW9O/hitQhZBl9P2v4AJhE9FaYUV7mmFT
ynspVb+/VVmOJEPTSC16Bva2yU/DXDyQLyBVO0/ZhEoGDBYomJr/qRcjfVK7qFqI
AAUrhC1M5zHOa2oiAENGA6m6za7onC3DpWKbYPyq4BTiU50ytmSIM9AfmlkSkM91
+4RmzGQq1zGNzGgBVpZZ3gfbEv5Ndt/niaqhl8JnUpUh8WGIZ/84KYEwUcGln8RA
DD+ahxI+5KlRIp31LMf6T6qlDxNtvIlYHJLtBeSQuarv8KKaVpP3jLFEwvPrnF1k
cU3xzLr37yMgeWmi3++aXiRXCPVkRRhhlzK3B8eXZHaaLZBFKWdZmJ2vFTSWxCuO
LeXAFU9Yd+6Zh31afADHfGhB+hh6E1wSVcs+MzU1dhzIDHKrvv++SF7nb0mJ8m7d
DJeahgOD0SBZMk+o0nrbBUca2mJPDps+ag/DfS1tw44NkjlQtZoF2oLH2jaHNhCQ
pQG+CVC0XJesSGFtaoWBrq+0ru6y6xA/gkFpgDkkJBY=
`protect END_PROTECTED
