`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gz+KcGGziC9UITZ5O8EoE9NM1fxxjEImVhkJdpFRaSiw6afqFL8ce7XrZreG5U0f
O2hDSZn8VKeEPw5xx78DEeWA0u5KFUPHICb3n26fzZBNhaAFOrYxB/aqkr07mb8T
yMJbR9g48Bru4CdPQKGNV0Jz85Maw22iVdreMVV4s5mERATeiaauumYS7CgSxBsS
Lrx/AU8825nuUgeRUKxhiQS2c7wPrH69i+f7mNBgd+iWQPzxmRefDi6keeMmBjD6
DreR1FZXj5zlKhO2gEJiDJT96Jki2CR/o84d08Iauyag48TwSBja2fn2BjwiF71I
FdTX5wK3ZXq/Pl/Q6l8zfZm5FIlynjqrtLwtLca0btIZPbTLY+XZWDIv2+5sFQJq
ClYe2VZ+4OXR8DgItCmuw1Rhrrztl/9ppnLE5U9AeuMNKCZIasHNEa/jjU/SsUhF
ONxSSfa74yurBR2KS2u5LfZ3B8igiGscWhawUbPwfxlFHN0RRktNl7lPCH7Pnakk
dL7sSmQT/7egAoOOTXNNj9HHtfnWqji7mYDtACO/bNk6UHmAW0sjOeI9hcDAqQdj
0fQMDBexVgxBCW8yPIQHj4U6Q3zk1XG7ixw1KM23g5+TSnjNBT8tpaR2DFh9j4zd
2ZkfTF5MBq7E66/mXEJ78hLQLnyBGHtatDV2Ud2ZxU7OHELl+TGUU4fyx8WvVDwd
Mcz/wLl3WGlGM2dVPSQaLJ8iLkp64ogf48bp14kUHX7hxqtOx8hEJ0HXZ6fwd2UY
tMQ6XvVuNhjZPA5vfQDwwbhpdGoiiUR8VjFBbVaH96HNLZKVO+iHdrUnbj4ggetF
j0A0YqHbT9vQnj+8pGyfMQ==
`protect END_PROTECTED
