`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EiH+bRcUviloQxWqeCu0N248scqSKYGHs1k1bMY9a14b4yVgXGuyqregZPacI3Da
CYNvUxeM9chd9a1aXIyK0UZ04ItajEFW0xvGdfZeu/1PZ6XqurL8sorzPjp4cg5t
VGtmoPCIOhESC4TPhcbjK+3mC6YMxlPO0dTvFfwTMz/7tY5SoLi3VrjA5wAVS1Mf
iCMa92nANImpgWhe1a8CIg8z1q1LpP7ag6R95yGW81YtMMN89oPFPhslvZbO37v3
Hzb436PwnXgOOMVee+urjEZ58e7zkwvhmhwP4n4n3o6hVDz2ioESLk1+9v0Yuf2K
zcZ3eHKuwZ2EvF4KWy+Oh2Y9oPbONic2KN2UTfbq6havo5JOQIcWhDzq1CQhDco8
N1iC3H+L29JC3r/U4Jt2P+3yJ5N/2ok8oj6RE7bDuFR9zzGTjPSTuGeiJn6kMq0b
M34QtVZ+PlkoC2Z6aCgBFO4j8ZJL44XIxfTCDV6FvmvHMtEiH8S2K8LJHu3XjmRE
EEYshZ7iu/v3qxv10ZxAXf1UDZUIf50yENHlNG9cBUpZIyb8+Iu2NQ6i5iDUeOyH
`protect END_PROTECTED
