`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VH4VuEGNH5ZmRQSr6+21R71ZE+obJb3jMnO7AnMs/aYyVh+isVIh4aXIdYu3IrSa
6UJGggb3qoQedriHN3U9Firu7fSMxqP6zceXd/G4pb/QAiksbwt8oBrdTXNhhNuH
Xavq0a87QEmwXZVzohGT7lQa/sBV+Je7IJd9MB/3/yiegnRoNDfwJ4OfrRTagCJ3
Pz3RJSBneXZ3x722Fao0wWLwf/BSgSM7Q/enI3eIGWbbwyTJ0DWDVPNDQ4eolf4l
+c2F+RJc//eYqsyRrnxc5KZy5j9o3zaWSF9NV81w9cuxdXFNpPQ7NldbJlwr9skq
VvyO8kPXX95RQUzoBxzecLHOVMiTKpyUpQokQ5LAGWJ+ZLymY2iIIReRcNZARtP2
Zl+GF/47MuUkirOOvNud2LlcxIK2rNjxDkrEr8XpvqzD1gkQce0ms9pmZqEBO6Ek
uPnW00RcNBBKz4Hm1kd6ihmzXcAHBLZDxzh2TX9lGR/1k+dfGWk8uA3ARO7fMver
4kl+s8dtkZiHvQPGqgU3PGa5VoIwkYmZaEQWfXPLIXAdB/OM0v5usD6ekK1JO1JE
+AaAVifPSbIFnEp9U/bpYQnB7WTyWUjVObvqMcPv25xp4VwnoeL2CBmb7QRm5Yn2
qMgiv6QCBV+gWixjgWS6Ie6Q/RbkvCPfK/o5BYU1CWnfZmN0pPjAcAn3agu76zr8
ChFaRBPmfdwVH+Mh3kMC9P/loGSOwlWTAEw6XI1ye2j26gNroCxrh3icwYsHgyBc
YJllmUGEdvRNQmBkMWyLEdOGo1vDP6ueeEAA0Tvu2l3Cua2vCoMs+C5yGmtePr6D
2M576u8jsuFeFpJHuMJx/z5W0Fn9z+wxpa1zd3AaEW2NDh3iokRAyhJ3GDF96VI7
qNOySki98zsAiyMba732c8Gp/mO8cwXlstvI4oJPCOBliNI8DE7U1bHpM/34iDSI
fAvALJri0es91VaVveV4qIsoEHvy4okj2KhJY0XnCTidroVzEetpwK0L/2nQwd11
PaOUR96WKNP0KX94fyJodspeH0pbzZbYw4lf8faGSqmVY4CiAdavJmJCfHLzHgxJ
+OK2T/II0CwmmXT3v46VL0Ybdtz9ob9SchgPJ0Jvky+bN/sw2KibQfDsd5riQyIq
JHwuH/vVEu9fuYDnzGERUu65x6CSKtZlR8hEWUMLIxcCA87kGww5EM3PcTfrZQAb
UoT8lX7Xc4beRzzIjzU3TGNccI+97jbLXPigFh45n/PnSkhC06a3apLqtP4KzOll
W1MYtIfANV5JNKk8bqPdOUh6/VOHdhBOqReMK3nlyBfsp8b2ZvX9COXiHyR9ueWi
Q83+iCjyIn66sRZjKztDxZcWyZcC0l5FKikBo+Oh1UCkwyq40/9vkfeL/ybxqg9c
EOQO4WvZSjuliHVsxj+RFRBexJclyOj2evPhXCjnoWO4ps5pQ6Wz8lT0qaPipMoL
+hsUjovwb1rkgUegbzLdChIIwQHDbie23hx7fGtzfnR5PMa1sSpyT+91Dfi/MhzY
QputtU0i0aKUpTD0KABl9Uu+DJU2YzrSF46kgDdZikztcarwQtUjAXiWs78vMCOU
1A7HJ9D+ooV0UufO25/0ZwurmOe0YRVK2QPV1+zZNcCZGbttR3SypBk4Tt5mqBza
XqqRjuX4jR33OqHe8b3y43wZApcmn7JTnlmg+1KJXgJ8BvdW7+jd8GESJP697AG3
pIRfdZzS4BHFgqeX19EAnRGXxbTbf9eWqFj0WGl6zMUbeFzwnTBjAK+mJ8+8Nx3Z
Eu/rPJS00/Q9kINFfReWN6cTmTOC6ZSboj1WJXbxkL2/9alACG+GlYsKY6TlSGll
V++W0yAy5g5GycJYpxBybKb6ldQZ/kFKQmk12yym6RAKFO9Aen8xzVNiiR9BhQnT
FW27dSfdBiXT3qDKo0pvwttzif5NZftnOJAx1fEl6Iv0oB1brTGEwChhNJpHuUyC
XUM/95C7Co9u3LS0ude1nSM78eFEj79Kk7oWNpzpYaRs/mLLsUAWdLXD/Nl7BAVA
1oxG1+53HbjpbW3T3f09CzQa+4mQrWszCjz++HDhYFagoszsreNd7kl5c8wQt0tl
0M3N0nC+uKVXODq5ixYl41zIBX/89nzkZ4NvCKe7mJ12xYBQYhZv96SEwwC0YcRT
wGO9RA6WVfnqvT7N3uus3QcZiuQb+ciFFRuX+LRRfl6e3NFRMU4IePWbGXpgPyvX
OoWMRN/KgJB6oZiUWDAD5rV5IU1702mujpqvm6LDfpFlwY84k50AbUBMpy3IQBf1
pzyuueN8p9XjmxSbntaxKI/U0hjCM2FUjUh1aX/Ley0exkV4K1k+nNNVmqNl2Xzd
70I6qwf9SQDGOb/Z0XQ7jypEo+L/35ksR21pxNhY59ZtXHnCDC6WEkp5o4PZOOQA
pbNByG7HS+QqobTFQ8ttIFahn607oFOpkOF6rHPeBG3VzE/47SXVgsOePe+XTDFV
fgCPAtvS86sG4D4v1awhGtItuogBgcs1zBY5iZHZpLai9W5369WFz0rIK0VIaRlj
Tj33Rl2w+DxOE+SgzUhwHK0Y15DYfNmdkWIuJYaerNhDT3p1zJ8QusPflhjjRAoC
gH027G7kC5LLrMfeNHJMlyWZy3X7U24vFZzRv1IbJWUNecygRTo2XU+875ms5buB
r9r9RNb3wbJhpm/TTPkRAMNEYVFbyhtIxZTbEk5PgYfuk46edWsBm9l8VKhmu3Bv
4pO59dJXPUySNeG3lVlPThCjRCk1opUevm2Zy1hixMEtG+nEk3+VBXU20MnmJgww
MUa9B32j50UNx/vZi9VAMNX5dzlubEvGJ/gO8cPzBXsO9NbFHKVpyeR4PyBF4/jb
ImKzSUi4LTTDY8aGFLihQlzAcOclfZaVZdAlhgDVkMItcH3Ev4VzG4OxAis5dhXa
6SUtDLxH7KN34BFJuX4AVYck0V3r6U1S0w9bLLpq8fKNWZkfUNjzwVp2OCT2eurr
5KuhhrMhvbNnRiQU4QmKoYFkeiQdnhKW0m4wiBFeTl5IC0USsvK97WZ2jHhcS4N7
SnCP3YYJJVyi48PK3n0URfF0V/OI8MyROaG7j5rxPjkOh+/XUVI5HUgdGYy0M5jS
AkoS1hlY0ezcO95ubKKfjh5K6VFolWXXeCk1bbohGFX3PMYONjq31wMOLAKQJM5j
ONIphJMUdNUtmihY5VFR0ocwGnZf4wn5T9h5V+9sWM2FHCFzLXFPZTOpapwwIa6K
11OhSMn71jFpSuTRnXRMfVm1kqKeqSqZX6nKylekYDIChQgZUWGEJaTQGEVfrHN9
f60w/BbduyNVeiH+D7P0NtZi11SctCkD4fvRAdWAhG7x9MhTsHFWYBdSU7UdYqER
ojNRtc0gW8Mi7J+1mNxsLPdaE1A5SP7xtbBzqBGbrklmLY8NO8gFf3ezv37dO2qn
dfopuMcRk+QSe+r6WFpJq5woDZYnIvL8g+t8vY8D7wYZIgEwne6DgIm6SFqDv7hw
OqAodjQ5tE8TXEKPVgQ6IIQNWXK3Db9qxfJDuWicghWTvvFQ/aOiUvkp19Ljj6lr
ZEPHZbkdw1osViRwslcD76vvtiYMv+VZKlLyLScBO82D+B2FeWSJhEz19EJZ+7kW
1Hlt2dtSNCRyGpKm2fAM6UsRGNRFFbgNvs5UQUELzpWZwYNjkOnfZ+Mk8WL/IMRs
JP13IsE4PUSCB9JRLmA39epl77Pbv6Kq7n3qeQ9/YXk6JqrCkkzKEZpsmD+WbORg
IdZFAi29BfO6hd+Qwf/Sr3MvC2p886pQ2x8MU5hjWHdE1J5mX5mjNVq4aA6+jWWI
pXsHx4ug2Mc7xdR8+KGs1Cvrv0T2Ftkw78xkUWHTUaQxHeW4IjLCpDY4mwz6tk3k
SFSaDgdI6AGOuNKxUIGCaVwu2PAd1xZQrMDmx28+qhacWygZ3KDYDx9xVImrhksG
Lg5nu98YKTPyXHFjf51NbyKKQ8Fyl0VQSx1U6KwW+5eKfQtJnS/4i8mac59EVoKF
aEe6FCfOHCRd4yqx48cZVFU8C/Xfg60SmUHgPgI9NPSuXvbjkPwJ6z+Xd5uLW1rQ
RA3jPRh6KXQFd1OoNcMg6AO4n/HwhiCIJCXOSxO0pCK6X+B2aTlIlJgmNXTLa4jP
OYElisMkMoEyM5sEe9axSnMchCdIQBGgx/K7Alg7vK8Qqh8POjIdVpyxZjN3WcAv
pp/artKeDuouPVSarKIw2IowMWNcmTNaCi6tcKMefVCwJzZ2b3v6FjGCP8XSkdZi
W7YLqs3xl+/CZKSIPizbw2veKyw6AW/LlM9vwid/tfbF0hYjAq8HCCN64PpSIzPv
H4lLl9pwgYuXMZ1DlSMOBnrFt9z1qnRLNdHj0WTZW1MUO5cJbGDvLjy42V064nq4
wJaQh28eSeZOa6GFd8RSouCiO0hOA5yvdBt6ApF8vHQX9XcozVwyqsjtpqQfY1+4
b5bweU1qi262cJLQvJLkABTWE+gsExAETuQKoQohuYukt0lfVq1WTYgGi+DlgS86
QxwuE15uymwzS2BS2p5K25Ujm5N4deHjK4BL0vXaYiIQYE8FiwVb2td2Ci2tAB1m
+yqc6btv14SigZGY23uloidd/AueG6jOTXs6ikihJGuzMwmzADi/viBrLgd9l6aN
NGm1/FYXfbVYxHJUgODwncfZvB4MymEYuiKc1ktrF8GeeiRX5rTXjb8OXIwKrpfJ
dAqryOuxp5xxUnBiCR1W5pUx+LXOJUiPfE+vGApFXWUI4EdG/in9QrA72m1qYQuS
4AL0tWk5kSjdoMmQf8MUEd0/zlTC0qGnVuRTIiAc2Wv1dTtUawOz9LQguF2qvGvz
qOuRjgdAmcFy3JP3MYkUjd6WIzui5940sORn9rwkO7lyBPlW+O3U7YWW2/FZVAAe
PmjQ2Jcbmin+s1LIDCvOo7B2NmfYfU5qDNWJJQGPSwQY45e8LzwuewPcY9ZcqDca
eYhXOzFtHZi7rv0D7Ox4eAOrQovNxrBfU/qfcPv2BJs4XrfimdLc/RPlH4GB2qk7
Yh3hF50tLiFzJ64q+gHC9B2RPDfRRLm824NSbtsNEZxvRlK28IyGLf0OotoPNvRW
hX/O8pJS1Ml85v+B9WdO573DKpZDWZzuGS/ICft/DEeMqT2dS2R0s3L4v4u1BF99
N52g+BaFb29KjzwI9t92Eb6Wl69ZZE1NwF2FWpuaFlHil65d1k6J4sO+Q9NgXEo0
hzkUIxnZx3xARhaXZpPdg0aCfyq48ZKHJpt655vIP8VgQh6s1IIPDwSVW2l5ioKg
FlFZKzfRwoFRtnqnU1f7sIkFROyz2jsNI/QRy5H63xeM+aVlcKnLonnV1sxkdeuM
2M7wiGtlofSuD5pyGzG5UoZhVvEn18HDbmag72IGNAyaTvi9x9HRHOav2T0us0wD
AQKxJwrj1WRF0i318TRsFa5IsJpRo/mooFWkuaksYLRnnHp8s9zYR3Tm/ivjRiWQ
Y0hjsIr4UXf90Wo6akFHwtPUu+2fegXdER2GW1W33NJO+l5Ne48laq38mvjx3Bdm
qCieS4IQeiscxYyMqCnYj2L0zmHuQO2ySYNgQqtMwiOwKE69h7rGgQv2tZN419LE
QcNAOQBzWjwdZQeMT1x5TLPefQxPtjy3YYXyl9tq5ulIRxkowT65+3A5XNa35vbY
GKDDfmU5DuV0TQ7r24Y0dSwpdlqgQl/NUV7b/uSaadj/RxP3EOLX8c2GkSbozslr
3ycn1MYFwvv6YYmDTVBpmChaRQOqnJYwEB+8Mwrp5KiaOo1Q6jWXfya52wXeZ37A
f5rtOKUdsUHFaPVjbMIM93JXa3Nx9i0fsI7ph7t7nyA=
`protect END_PROTECTED
