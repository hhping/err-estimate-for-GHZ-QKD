`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wY0r0R+aU6goSK3hT7g8RXoPxowfzI1nDdZzb+W5KqWMXEKLqm8IHvw5N0effaVS
5dldwKLyADMJyShnlybwwb0fzrPHOIeWCdkiMzhQzAN0E+Or6rJY44Ixon/WQ/BS
75YpvmQN0a8XH4JmGBcKgpcLqHgDLVEmeFWz4g7LuaIw+9BCYnmgBa9bli56EXZI
ri9BeL82N39/8BCG7UNzXv0NVo5DeK7syA83VnuAGkiZ02s4uc3Z6GBjJ46Tx/gz
oucWxU/dPVMCOBOFzsaxhI8DEVgch2JyyzRc/wgKXmgl2gwK+BHJ5vJPA6UrXGWE
eOMooT5nYIlrpgLinN/6Y9Q0jn2VmnGd50BndvyD+DUklbh7E1dw/yaG2PIpVgn/
sYvF8pvqxEA8KHl0xbaAfLvDH712eamZpcS69JTNm40ssfKyu7O3CRrv6TJcWz+r
yaZ+rtz8K9fUnU4yt90jArGBuYoHRIGzypexi2b5WnmoiFgaGf5QSSP7jqhJ4bLs
p70gv53I0T/lnoY7aOjkq273eebRBp6+uHy+Su8kF6+A0G5A+Y0nw36NQozfKvCv
ZeRdCoKg9XuANfgKL1ypf/HL3BNxWP+gYRPE0JOt0Lyz5w3r2x5RdhRvq/ES6BFT
+TxUYEoPBkgvTw5k6M8JDsEMWw3HoLty5ixvUWO4FB6hc7Y3AuLn87DFB4nTMtcK
T4aoS19GWC4Ls/wuGSXWiQ==
`protect END_PROTECTED
