`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Twyb+OtusOzp0YKqVu7XhTo3KkL1bc3ltwHRgajSX+fANO3jcLRQuzKkXoxm74rA
Akzki9L5uqeq1Pez2oxeKPfzTyK7RdF5QMr0Hv6UdeN9++nh7fv4zkLtPY9SvWkF
5C9R/MxDDjknG8/ktwnGEqmqtQreRemeL8pn+JjW1ZpkZrHRWi2BPVNZISUaMJA8
GySq6+AHViiEXd4lSXWbwz/XwaFqnF0jbVndHSHsEe58XUZS6Ipc8pNIl/AZEJwl
2vbOSApPLHu6+F/KeVWpOX4LA+I4Gn0wTWgAu57OYHMyrq2tmwv4ezXTOlLwtj0X
5rC+TH00U/ZmkXP+LJXfnf+FO6+bXCUwCxKI5JxkIVfdELkXKjrY4sUIqG59W8eO
fp4E+dS5pf3Uw6wnEomaVi+rhPtQ9PWAcG7lwUHLZHHextuYXBe74eGX2N5y9RDG
QIcGQGrfc1Rlp+rCGBQk6FnGWxgIEqNJfCcRAU9M6d15zOUd/XptF2vL2n044QGd
/viMTBtn1yJN4dbC0Sub/nxmnqe1ms9Wv51UWBpXyv9KbtLfvC048KeFh6FDGDm4
SgT6QNfshALq6IwVr7t9Q73BiWrAhsmR0Fmdn4jeDkI0XshbRe2NrJ1dsDk2P/Cw
nrAQTt21UGFTmTkagEfgiy9bxIQqfqvjpTr11SG1+CsM/xUeVudSnZZ1xTF7hsTw
NFx9BSso5SiBa+mQK8dM2/tJRrGM/OSbyM3/uIy57YZadzhaQxtWctfxsVN2VjeP
lFyPqfyvdkYs60lC11nFifwvngCvH/69QxRBNX6nfq29gfP4+MsjOHGEob+ErCGa
CPjb7E0fPcMaR8O7mHgmPszwlNTPXLDHxsXP5wEHMMDXdODVvW+AB9ZIEqFKVPx7
2Cq19EGpIO54R3cLp9gEz72Ob4OR8IAMrzUtI/ltXyEvMDHoU7VL19SpSTi3giHq
e++BF1G/RdljrIPvbZVEgK8j9DyTM/6LUW4KUNFK/EtzIuigRBJTexsqFA0MJ/95
/hA9arGNTcH++xtddebr6v0mEh9yX/b+O2D7JUH2XeBMQaER8Y6v8VSLPhgXnRa+
qQNEYa6GYDuMu1zJz1DhoYPQNqsgiFKDmPFOdHB1v4b6FUf7ipSoW1tYo+Nf4xkz
NtK/zSKoUKc58eChwwBZR41CtuwU8ux1ZYmn4gndOBMHjQMzfK0p1r7A+fu2Njlk
c3iTlXfakwWVdPQEKHAGKs/8hbXMnPeoOCpRGIK3Hl2lkS8c91fTMHz1IS95CEb2
SanYdtwplHkbeNYw+xXoF8hvqe21LA96MwxZVrmgfeTuUZgeDO0NTEyJ2u089XGi
2msAOYpfAPAsjP87ItrQYH0zRzKKZwSkXDjE+JvPHHfuqprZ0QfcLsGZTnTnCLoH
eLDKV3TlxF7088gi5iuF3LY8hraQLuRUOh7T8hybQ1F3hSt/a0xahBlWhdvgWCgx
I21ee1JxzZ72DVuuw5MA3l7L8SiT8rRT7OMDzz7is8s5In3sJJdNT3QlYQ4F+4mB
/pAbtIt89Ti7eZfbWOpb9rMV2d/xtso4DfC61gyzcnvO73J725ZS/4WFpYzkH3dd
yni5ilx0QJ3XEBEa8wImCCP7vXPjCbSBbnBx228cnzGOl+/bGw8YhUYWbJaKz42j
3gqgmYdgfkyzOKSZs/1CP/nxRlBNcNqb+5V0fQoAa9Vwo2o9nTZwrDxOhiqD/5Vf
X1LfOy0GgLPeY9JKfD3a/SutoT1s4QLYN2H2yY1wSyDDsDeQc3Ef+RP6UtT2W6Rw
Y2PnsYQyA9OaEoTZMzou66giPvn2zkDPT4NIlvI+N/0oK5cdOtZtudDcdMdYDo2J
xhMHuYi68AbN3Eh+5+FPREl4d5nWYWgdv2Y2i+2trwXhXMhhvhG3ufz70kp681yv
P1e/k82NTiHB1P42vPSd4OPMJFlUgqzmTKk8sA0cYbiOJnOPMeC7pgEyesDKC68b
b+yNBv8kB+vBPXhKkK4/bA==
`protect END_PROTECTED
