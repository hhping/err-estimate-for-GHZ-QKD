`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3nl2xlYyUs6uJ+Kd0lvtQFd0duj7DeMI86Lvceiz1o5zut4ZWZp9+exfOC2JJNZO
IiBnrcqBWZz6FtzmaF2Xs3GJZL/BXYNxoUexJGatEsfu8rigvf3v8xLuFtRlR4x9
dEdC7T0vmtu7BQy7aUNDqhPMfFBrRLZgG6Oo6cFqbjHLmnvI/XotLia4fkD5SZid
XGBv6UFWap43kgqUeRNfP6akM6alE9muLqKtYa+/O+J/hbwGZaa1H4bIJb67gS+T
x1uB/aGGLOiUYigvfmDSokqeQ6u9xvraKo1mWnYvFu5/lYelsfLY5z/4hQnscdq8
7KdVFfRnVBKU8PCn+Umyfzj/qx4iQ3qTjlbMgMsiF22JFNoxdAgZISj9xdv8T9J8
sIJcXO4Z7x2Uj9+JvzbDSb/fssginQ1TphVfZRFHepI+Lph/HlE2eo6m6cXoGSAT
qlamqy5fDm1LzFvU9SFdcbmjiBY8gc/vEB2GVTRZ4xF9zWz9/TaqrY1Oro3yTwkh
j3qtSgNvZ0KAT1wN37W/ZHCUKpJU14ms4kI2dTghHVPUZHvcAoFfBU0mZnlD6Kbh
oVfpogty68qD6x+oPU76I7QjTNzBzt5REDz14nsnCgm4LiBZ+734zd2b3nI7c6a3
UYr4VFOZsLEjjsHDAdYf5BsiKGZp8pYrsqmCAO4vQke7WzFsH/nYEiRPTNYxlKuZ
aRwDWO1rzBmlQz2cOULukOo6M9lH07YeAYWePoHAbhTF6hTRSgIk3M4JugNmRcpA
jC1GwGB2UMmssu3bQYh7hYi9snPCMUUTWChJkqT6wBQaObWklasNqWltxynkduY2
LhoNn7nPmDjqtM0jcOBV+OrUc9O5L/lYhfiiUyYet1P8lYHEeTohswVR3stGWLLp
cwD8ZGwyrwa2Z6kRpybJx+WI8ABDQWIQIXVkYwCaog7mtN1/5RVWqz8M4RRWoUOv
axGfdRweRYJXUrElrnCqGSKzgZqh02r6SssSN0FCXRUelKJsiUChrev2UFxSNI5z
06Aak1VHwk1sy33y4c4soolGQxdFtamu7JFKPVuYgYYFr9cEwFq4N3zCHa+RLEFN
EHPcBebKPh5Xmna3Xp9xFIa9spGdozYOAy2xJKoSlllGinAX5FyW3y64KdjnUXNr
S0pchMD18djYGABIxPJJYUQbjcOxLVlJYVr6SG4uILLomRVcsBCdlBOrstNfQmBa
hXUyTd5jQwcJkAZNZRYyTYAOSMAUnl5KsuDuM8I6mxbAOI4fTd6Whv1TyzTcRnBs
yeA903R8hyoTOgZihAwltLG/i49Z0kYLeK9NFe/eGflTu/C6Kt7BiA9YYgbm67uW
Y7hKSrW7SavsoG1fiBFBFxCCCzsBe8k/zOludKnEX7QQuAQVV3XIpxRle6XrU/e1
nrf8uj/jl8iXW8vGb5gOOcXS7+fyxy76UgpBwzSVhNLxZcYPhrRL6S/usgyzCLtL
YsSyvWjRYga6vCVCF2EWFwVwMrjHDrbCa1bengPUxJEx+wnn9LXTG6vDoFtyxjE2
KFkM94r16X0WRIVDLF1AawK/v2uotmYTpmyEOHNwS4bcFqyV3VGn6b2bavw5PLxP
3IrRitDCrnOvI4jXiuxM0uiLQa2a3FKAXKmlFbv2VSfLjz9K+hWULUevk3UnF9WY
sbKudGPv6FDKO/xp7tm7hu7RcHsM/7bAMWI2wCeyLLIGJe7enghRLZwbOJ7G1H3E
GGwYzZeKn8UlgiEdatkmbFyh91RqZvFjPvJaNsZmlZnkengvv3R3LvO+2aEiqsc+
fj6Yv7H2fqIGammRUEx4A/QUBbnkqZrlM8IZUb0oYuHO/S5h873rIYaXntxWp/a6
vNQEKrCIS6jVUiKuNbbeZIS9ovgNo1qNBVsYmIrctRwPZ3S8rM1cFwbw6rEtTTb6
qclId+C7Ks+YdILF6RECDpfJESf9llQHxv1o4ZkjJddOvZPAsJGnWWdBWW//w50h
PoyVzXP6sGkl6eRnna9fi8lTSrY0SzsB0q4sOYrgPHpnxxKunaV/ITlW5/SMuA8c
Ze+rXJGBj0ENMN2YDVptmVrlGcF9yvGyXKtkQudfKKhrXmjaiJ2wF67A2ZybtLad
xsKQzVLtJWO+sbcD6e6VPclekTpA4sC/sGNFIBIDcshg6aHILzW9zXSETsNDpEqz
GCKYo+QMQAOkUdf8bqtVNGj92Xo3kVfXa+NL6Kf/BY/Bb+oxZY57FxZFfZM1ICVA
15HSXw8DOfV1HGBv5KIT2yUIRi9P14ydmuWCCJhjNs2ec8kcvSPK8A8q8sCA4vVS
KLp1Ls6JGgAfxCu5JH6xhOQeNK4vgyF8qH0xP0l+qogVFm6PwZaMcWz2duvy3uUd
aeD0h/UDc2x73aJ0BFFFI8ujlW5myspkA/1LuWEVB1/kmTw46DcRggozFvtT4OIP
WSicFQTFtx2Zw6SgXUD5R7Amfvi17iTM41qHXur2fegPn8JhOQ1ga7Ja1BnEPeQ+
pqFs5fcHfIRujijbKVW0ASIqPKlh0vzCW7LIesVIccteHE4urReqdr+PLdgJ0/+V
D3XzlWb8HxUYCLRQO7rdsHv2lkXn7zOdBGH1OuzaqOlFqtvOzrfThktcFUDWl9p3
rkcqJxrTyG56jtUxUK/XkxugrkCCUZmJ1ZJjVUONQfAfqLniKR+29QnD7XjH0dNf
Q+uN/S+eDPa2If9Tq9WLii1o7x9Exf2GYF/QmfLE7d6/buA3zW9A4QlmQUu4V7LP
R1g/sxaIvAWkwc9Vqw5xqJEgQpaei7HqGqibxPzuUcTzCnNszby17bV2yqi/lwtb
Vs4uT7yIrd+CVHQk0qpyE9vclNhqfXCOkD3FykSRcMSvvubnHA6xsejpOXjpmvHa
k4mbHLQvCRqxqw2WNdu9i4AE+ztz2pXePGueMJg5c6C9i4BF8QCv6ughcKr/YLSh
`protect END_PROTECTED
