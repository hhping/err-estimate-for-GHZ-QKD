`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHcgEKplBGMijtxDOSjhN61Ad235puuDPdp/1PKPbTqtIgsYb5QlEyK0gcofSsik
BX1g4vCSRVW7JoUMIJaUdKG/d9PQjm5oR/4+U2+nVBdGQ/1Qd3uoEBlZkcmpOoVj
n7sGPJgVNlbcHN2owirbOjEfkOB/Oz4vJFKd+1GEEfI2JxngLohy9RSYQuiW1plL
oez1pu2XB1XewGObzUwvehM9yHuG5R4dwYcA9Mw+JGrUCTNHHKOn6Xr9srF7f6aw
AiV8wEEaqPDdOeS0LGd4nFZXZ0PoNJnFzyVN/J1qjJ3Ga/jyfIZbcdotNpzUGTF+
vO4lu2lkqmCItEVwQKIPZNE8088+bbv51IxzK+/O/vr3I/+KuP4M631dCsFfyqFl
CQeonEtSVqeJtSWRoOwvv4MKFWg803rOb7MSaPVYfFanZP2IFQ3luAV9bUErLR1E
0ePze7BoT6zVPK8WLInVfDLuaBNnpVZhnrVpmdFggyPlmg05H/z2CZHAalyH03x2
qAl8b//z0OyMBF0RcMflVrjSnOLdL1XBWOcNuXMWPcVCVHu09ciW8RZzxUkA7Aft
t6xO2L7cYPrhWZZXAx3BAq4C+U1ivt8uNc7KFshlRGBrD7klYT7TORqGEGBqKtiZ
2QA5cuDfFr9xafXHrbUl6xi2iZJs1Xc9nYHmU1q8hzQQPYFASLq0gQt521qBHBFK
I8rAWcSxle8Y64V0fze/sVn/pwAi1sbYNICEdK6CIZUwwF9MMhFVFdibXKfeFfuW
UEpjAwUADyUneR0suEXU5lJFKTFmmQI1kKuPAcUlNxwz3Km0Ws3q6VGTB08Nvuaq
uKa5lHxlHEV++1hXE71kV7202gBbngKkrZwL+DnC/Gm/aBD2kKA536HNxm+KX36V
7mO7FFPwC+VJV13oIQNoIsg5Tm0FbDNi0EMSSSSik2KSXMb+9TtLEYCqqKaV0uEe
AApiKPNUK2b0UvtJXJ54NeIGNZo3/HcdNvmkSqpM9g4Kss1sOKECMWJBJ1RRy4sE
MRUJY9ROjVpGX4strY5lozAgcrXrDPWCBGMa5CpHjTsiF3yknmbg0tKh6TU7ee+x
if9O7loEgiDfe8KzpLZh+NU7Uy199ltFkadWpDzvP/hryp1obx95nyjswy+dq1Ys
VG9JHIFGsd3Gaqh3s/3k6NkcS65p8OPNY6NpplRQW7x2QaO/0MqMi2Wbl6hhefZC
BDhfY37lRt4vWKD/h/T1vs9WRd6CCCyseNb2Oa4JKZpo89qj3aQ1isHWrER/1fcU
0KA6T7V1MZTlphoyVcNx0K8uVRIUDc2RC5ndeHUmoilIxoRUosZFYdWGfScqXSl2
n4SincsMWj1A/YgRkSrEWbMHbUKaF0L+/vvLu+KhPvpNRhqNivhTgqDH3repB/ok
282Up7Xz8Anh5c37aCx9C1COdryhHPxr7KxA1j8X+0pumpJDQKI6i9hOZaDB6U4u
BjZJQc6pFhClNC4yUfxLMFKg7Q8YR3W1K+VuscsGhRWld8+B10cz6OyLuoDjCIij
c+JYLAasuVHsfmJOARPfoHCTjE7dysCWT4N5M7DVoGYVomUau7S51DdsOdxrIrI5
N5wZfKmeoJo7z29KHe1Q4SRE4a39NakJZOATX8aqkw9v8M25WwBDM+Ax9Wn8gNML
kDf9gH8w0N9HzpKgvUoktsO0tdr6tTa5iwp2VyziBGUEOwMDGBTrGtGWenoTLluQ
kJdNXLs/+94RwJJooZotbWAZMbVenvQOYAqGcVlADa+ZBkOZ8Xe+OPk8mQGXCHZ/
ArQZe0MgSd4xE6IutVD6MSl2h0SbRlJYixAAPSW9ut5TtBQDQtRXyElteY4PSVEk
nG8K+fq74yQ0yQ6r8hODhK01QeNOcybUO6NpysPEkzcvMx+Ee3MMRkBjv/lrUtHK
+dAtWOL2SvcnoHTA+xKc4rfWzhFOTsEkgb0i3U492A7wIvScRIWuFj59GZpJVJv0
Ls1+8WX+lLAreNbzdVcjYad1ZuAOtA7IL2l9Gc60kuJeQ1EhlEJjxBO27lUI7fBw
eUCjjVmf9WQph+nnKfWQzhI5bbSRPOqguVGIwKmwaACH23zTiIzv1WMuvI4DJq83
XItXD1mUORyLeAuu+eGcu9vVrnv2AJrS2BFPU1DXM3h5GjdbA4i/P79ky6osY9vb
3BEvgbEi9NWhlTBL+sR4SeEUHXUqC4yWtQUSUvzg/o3a3aCw4TFLF5r1dzUY4J7X
e0MRsi+WEGFiELli3lQewTpdL+9CYWF8DgWPhuVaiXgqGBettiAfpniQUZ+wVwYL
3w0TQBNqQ5ljOHtEaF7dw2MK5Ohnxjuydvin40613fQReRiF3BxyfrXQMtXSpPNR
JeAbX9/VEfFpG9bT5l+2lBB658h/CljXKRAJJkqFMcaluGDCN60WPlVMBnvmZQwV
UHphtgZJlXfcpVuuIRE3AXNGtVcJJEfhqleM1uUHvU1UTS4stJb6K8isYvT6te5X
bVNSssxG7eOY0PJhzbGsUDaCr0OOsmOLPyhZCW1kfNO66LYp1pkqe5hdNsLajj/z
T+NuE08xnuiATMlzGdkzBIQtH9Q4B490XZDgSw12e7Uu/zuIe3Iwf1kslOhu4y+m
xsmpFDaV0NOrPvz4PHvw6s5NfpKNBhhqOQJWWBCTEdm6LDoBvGUJ7nHDQGNIbpnE
yWH3+rl4XAsMzzi7Jx0H8Cf48V9Qtf08SiPnjW3eP6XWJWmSCV7lt8jj1Mp0g6BC
+lI8eu+8XXwuKHvj2DbqI4E1orC5HH0+cazYy+vMlvEwHzz0ldSRP1Ck4fJbnl3M
G+gs5p/mMgScioyD7eEyRz9dcyFEkjrWNg2Nhvyp+at9E7Rkpy7eMblthCDnWAsx
fKsG4PWWlz3ryqpXtijkSzS41ysNUkKSWZ8y0prtNWmurzMaLieeZj/D1QkzGmjD
FlQ11/f4TMEIic/PTxDUl+/mo30DUV1RwHXjBaalx9/r+msDiXdahtDat9nKQ0WF
v183s9X85l+TeAkDqL2jw1gzZR3qC1Rhhs83FOuY5ExDCWUnxPtgQ2b0gEjUX7mt
bN1RVq/No4heK8v7Vdn9Crphl8pDflKiiWgP8dhbI8cVPe1xGEdOFzYUeymAwkDP
NJjPwWJiJvt2jM4MQbv1SG+aqy2rtT6JcjNjEGXMxmBPhVM+depmaEdru7kllZVE
iNo8NDG5QfTHHc3KHocTpAB7lcA3YYBde0ZVxWBdx+pRDsRBT6Y1fpdGfzE3Jw+A
Uiw2Rv+6h3iUO3ayX5ERdRzkE8AIEWGLykKTBNWhlUJivRYHQ8IRuQE+3lbkc1wG
lpxesvde+65x9SpqYc+IWtNa+083acUOzYKTenDn1d5JsVwmlT8C6lYK8bcWGUSX
otmbkgwq7ISejKEEV0zji/8ArJnY6rU/9m87aYFJ1yYTFvLMTw08o3aQud9ywyP3
sMCl/u3s9B//gU2dccft5HisXrhtIITY2rrXhEB6eQ6v1Kom02nIt6TYHErVGV9L
Xc1IIsuB7lHhm1v257896tPcTUCqZ0HkVMJCzWF/wwixUuujYSSsvj7oOyj81hC7
IBe9wJy9esBIk6jBuzKWMU9n0q0vTABhzEA/Cz1OHh8NWqkR979ge3FGCz6E4NUH
n3E9rntUcnezYGiOiNX2X7c3/g2uIyez0+UQ8QiUhZd1EFgaZ9v7WlwArHKtiyku
mQAbRvxd760/9W/mdbnfqwLJLjVOd/GLDg7UAcnZQbhwDlkA+P1iwRyPENsL/6o4
Ud9Uj0xzD0NMtA7M46qDZkyrcxwhfu/VhZKKeU7tgWnCnym/pqCbRg+RTnPrWgDq
wC7qZKlJH6LRV61PPJAUXCQdSVvhUx2uwlCosOrePAMVgvNzpx7Amr7ZuvSxz85s
Xxh+OmqAcrdXSs+NPX7lb53R+BQCaikGdpr1GQy0gFAZaysUqvV651bi8sw8f4Of
KU6l0UjtbTTI0b3UrOshRAYoF01nKFNrkcnTahUEmNExOHT8p06/+Egjdc0n/LYP
LecRLLUKDOCm9qrH6dRRsTuIF4SxmEbIKztkz9N7UDJLKNvdUw/YYfyjBvD3aaJ7
TbgFUU3d6aFvk2ObwWNiq/kDVp/fc5QGQfEsfPxQfHRYFFtTPDIUHpg3LeVNwQ0g
A+85hrd7mZjgdjOmDbeDx2F7uxiFQyF7S+tn7AbouTYt/aKDGfPRzGmndKZ3cayW
j0THuUdFYRaQK2C4b2O2hQ3m6WHLqvEiM8wjRGk0rSD9jVJ9wa3jqib4Ajhyd55P
e1eCtdhmyAo8OKSUu++Kjjm7yrZPgGF4FnSSTlZ6gTy76Ga3XBKZ+T7OoSKihSuC
MTnSVKYezTBnIp4UGhq41f8XyStjd4BDK7kISfsoVY+UNS54Anr4PuAmD79db/AR
CuJfJUrilVibqM1fkKhCYkQy3wDra6jxdYm7pl2OrXU=
`protect END_PROTECTED
