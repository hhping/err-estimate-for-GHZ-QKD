`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GngFWv4c+NF0n9YYPDgNytZEn8gg6aCuj2TaBxuKLVKQ/RasI5Mypg9ma8FoTD09
psNxJjgi840EaqwHBHR6Br+GXEuWzy0qSq6wl6294Mg/G00zueVlw5llVhaDCtWN
0UF987VVBphD6Q8NDtz/g1vUDz+uB2zACQwoB4cKlBpmGVskQtJ3jBsUnCNUJIwv
OkPyTk+Irvp8ch4Eqq0q6RFl+dnlfZXiaq/cyZ/54OSy58xcvmfj80bo271ybc0K
q3Fv3teRfTdqXoJ1wUvrjnvZXHdXfRC/79en5PLrCCmVlXeb9qLoL1A1O4U94/Qm
OswPk9oEi6jURWrpqN/eJRnu2nCx4o+5/9ZkRNgzbB+dpTyBgjVrnua+qPtNvEj5
W2T7XgxJ0wBiXCZSs0MCcHyPOshL0QJxsKTdEI+M/JTCLOAgxd8oeIpUVDKBDxMj
FDtRxJMDTt7DyXnfqLGSzMsz090Qei2gY06X8hUtLzQ0DXHawM8DX8lplwPOZD0v
lbkfpupelXUD9g0kl6QOJlVN+iLCAk3whcfhzZmTH+R9t3F6RdDh8iFTD82+uxIA
9/N7bS6c+8Oz7pUrItwOdlBZWbnUZiFT/BAVUdqd1XW0k0cA4gPQNDqS7+yjDFNh
UvkKZ5YuvPLFKUMr4lnOLM7BlhNBVD+d4UmE+lTW/viPPN65DgbSjpwUwX/hT+zL
5267TfG9jYUsEtVjL0OVgx1c8IdV6nfL0mqlltalka2NnytuuD6sjrXn0xFAXDxk
E9VghcH0fyvSWJJXXzwsIWFQCFGBaAGogYuK8GsAiobJbuiCssbZx0Fg6HOi3iSC
9G/31MurD0Iix829x7xIcQlV/dtl1nLunuMof+GeyIK5HYOqExwVYqbNxiMj63Al
LWSz8GZedFa82ql00VuqSjJ+J8qESMDbfbbyPE+2zWenF2JyRy6cfBhsaijvGcWE
WsH8hAH/HZjHDlSHjZU/zv/+6gnDT7E2G7WzRqoM3hvq9jmh1iq20tz5M5TS9JOd
`protect END_PROTECTED
