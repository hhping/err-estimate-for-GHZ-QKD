`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4OGlfUvVra2oePbmgOYwKUZfyCoCuvCsTj/36esM5po3ySMmhZDOt2EhVjoUIN+
+Au7NE2UdvDHOBzlSRK442YSNcRiM+jGQ+tOYMC7imkjR8EO5mQtAY9uRtGBZCRS
HdB3ATSbYBmPHDE/7hbdovtim+ZGe8FZeM0g+h75IsgXUDzGq0Ls2GUII/sK1z1I
7dbSOtIhXeU1aQYX+2Ftp7eOADnl0Nbrl7mlfeeq3T6swxuw5nLUIlbmEPX3+zav
FFc06cwdq6+aNiDH47efFD4UWHvo0Owv6GGKcbZy/+nsRlE09prhSdZXpRG0tNBV
ZVCcImInBkjt2VANKtPwTV2sQCtU4eiRjA3efPIG48pXkb2xiSVjZ4Of5qRG+iyF
laeMYJ57e5cSOHfoj8LV2pTpUKYMrsbV8O4Pb+4+3AlolfF+vwxN0xC5CPaKKc8q
hsegrqP8ayRet7rf2rHvwuW0yKzxXLya5oy+Jrn14JvG+pPN1bauDLeOFW4CSrtK
XbC+IRFi5363QHPlsiQGgCjQoHMAzavO1S9vpgpMAtPxW2KWlLhV2ER23Af21tWd
iUUibu/CBejXtklWIUJ10tZZfxi9Ul/P/v0MxgnpYIYvGpycIABg96dKlGeXUEyP
6O9vZNIAD8+bhBmcvSn1RWcEXR6Qq4c1JNaYV1T1tKKpvIPmsyZ7uML4DE5xD6FA
z7dkNXXWJQPlKxq9owyMy6cqQzo5fZPlvW616BTgLZQCECN1IzNI6b8uFtsZChnx
bMF7+TfdoreWK5AK1rAPsxXBbNUQPdh0t3SsNszLaQThvHa14WjBeTb84n9MIcoQ
ih7yhRNRwd8hsSNPxqza7wwOn1wJvzIrKsEIZULrB6qtpM8VBMRTXpiMoNKT0MWr
cmQcTc1UGJER2JXl/YBossZtxIJKWmHDr2RnpW3G89SgnTyWwORfBcgpQAbwgMa0
7Fd76h8fNRd4LCo9UB7JncyI++WduwBxQSFM5xivJx1S4tMM+q+e0W9hym1za9cW
y7sg/vCL6OmMTN6NbQEtxy3Bf817G5AoyQ9k9cy+Q8R0JKAZ0fkIvSf17ug8vArX
xQpXWEf2OMPjuBbH5pG1AW9IUhlga0SMDw8KBvqhm0k8CLAY0blrfUH6e5zNBfA2
zx68P4cM/MCNkdVVTP+c4WjYltoZrlCq73PIWNtD2kmLcaoOrhpBWsO1IVItb2Lp
vGG0VpRzQQl8QfcNAhNsfWUIrKF6gxEM8PWTJWZf4mgEjkd0ISEyuWpD2hUuVELM
2xFufMVANstOn64wEfkG4Kll3DCM+05inoq8yMlJSAjRTnajARu4HVDl5zwPNs+Y
BSDYsDpt9l/+MVAGCjLbAry38b0agDmUw057kAVDbAdYtbweyitj5dR4dXR8IaOW
hSod/PK6WrGYbUrK5CiienzEWDM9p6+RV0ZvXfHDiX+O9Ep9PkZEe7ws8/AWnxFR
5diZqy6Wz5w7z+ndZNbk57fsLcXjXIeXR/9T2c6lfgMXNVaT2pWqL1uBUFphKQUX
cycIkBgvtuPJ9JTtLMWqbuW6FMhoW5fpIi+n3k8r+vhWJl1RF9FlrqugL5Jjp6v1
fh6deS2921sKhl1i8VIqUgeIF5XQjqzFtfUUNInqESeql1LRo7qscW+NUaSBhLxf
uSiuZRxTisHGt6PbXa/I/Oq4augh9iXCFPIFc7W3Pd5JGTQu6DTYQ4O/O+Av9PMt
pVBssd8JQQF2l3ssumzpzp5+f2ojxfiJ/ep8kxZE3K3z1pH3wGeBFSKmZz/VtPvS
Et4OqCFPJvsO09itsAyM8FkJmAvouzSm0jG+ScOz+BE0augTEdr09sqWYjkR3qq8
Z3hapeg437q0tggb4ZjBXaICCWsIuGOHz8Jtbr0XFcwxyPNnQ1NXAK+rmmDhDovz
ofynADVm0dE6p1Zl55NXZkTcqJ9OjzGqca1H8ENdjMZmE2t9UojGWYyEyRIjPRB7
wlCQa227wvJH4vr+EH24UtjolTnQfhGMs1ypER3tcV6StaLjjk19IxKdeDXNXgo5
ZuWOmCuJj0IvmpGttFE3tjNM3IGWBxYc9+FsrF9Y3IDij7v4wzCshv8GQPEeMqC3
9ZNDD4MTiezijwFrRbVVprpe/ePO6yJrsfwO2EDNrx4hFU+NrwgNGf3Jd+qGY4+g
jHDHpoINqqQHGRZlwzHRDDYfOk8X41hhX7826K9hlvVlrDa3YpYG1McdRyCFP+Cl
C8Zx4PFBUkueaEoaWPjhtfIoo1C2KM/2XVrXvidSgF+OB5ChxvSfY4mXhDblH08X
YgSbE2d7oXhsa6+jFGH4BfoH31RrgAIxGCp1WWq3f4b+chw70ru0Q/ZCmA4ZEOwN
NNBqDF3q9aDNh9QBJPEjFsCffTfe1GMxKbZp0c8i+AE8z9eyypGwdGjJttstZShD
80+XMMOcOq8WUJDv2Rt/8bJ6wwp308mv8waAcJ6czofOcD78odL4b+X0KUJ1zcI7
VPExBE0DSE0gTwSsIt0Gyrzfwk63Xq+4IEmu4EhxJ6ARUITfpy21vgzNFkSrb1UM
Vx1GuPfAMPQcn7jOc4qqeM31abfVpcogdYlIRy1QP9VUy6Ay55HiUfg2HkfOSTz6
4aMgfDNgV8HrngwdLtWYfto9IxJ7R1B5S9euFJr39KuQrVMvq2Y0kS5AwThHpqna
9CduYq2m+LoteUfPsBARS1LjfL7HsPx+O7ihg0J6rV8hXzq9sdL1pLHoX5u5oZkv
c+hY6lgEiierm2paZM5kEP6zDaZIST8/Nev6eGTi5isDCf7OOQiY6QahnkHW2D5t
ej8PGuADTo2rjvaTmWSBlNk/HQRCswc+Kh5SNpZLVU/fYp3+yC5lpo4ieG6e6VkS
3Sf/4MCgYIk5ljEWRcch3vKYOOyQG/e1gbDwOZlUHo75LbpCIcZZbLO7fY+KgFY6
si1oj1sL3YlQMBbps2SbZbSYvi1UFB6rXvs9UPundziFcv/tIEpt13pUJ8tAXcYn
zrZQRXR7GpvKq87O72WUObtYxQwPMoQRbxoBqWGu/LBC84ddQnkCOeIQt4DiLOmX
rWBKCwhAJ7ajXgooEGKHFSskzvQl8EXO0cRwfazxNzDWBV7bKg3meseib2gD//ud
FK74p9yQwCR9EhfDJQqw5bV64C9QarOYxFsGl7I+qF3Sw0kyF4Vk02g23WhP8nL8
4KDzC19+d3xySl/OuPjCH4RAm2cDJuIE6wQgQUIzs82N+33L8fHnQ78gTGsPKw6f
0YWPckRRCPPnWC27wmvPBXRC0R4XO98EIzOyZN4nfUSq73FrADn7Y9eNgGmUYPfi
cPgUtMcjGMntvdB503XmWhEmiFQCWlpDw90nlrOlU9nk9/SLGLQ0W7dnxdyb1TLR
82NxSIl0/yYWqrkSYrNqv2hRwG5NUP6tcYO2iLdtbsyzjPP0VgY30l0t3m6GvTrA
zSE63OUwW+zec56vzHQ7n6Fc4HKrGHgrDjWYysSm99Q/pkYfE7W3h5AwEZThK+5a
cev50lY21aP7m63Hy7OJHm7gTTORygKGZK8c365AWAZKawL0YcDZgcZE1/WyLv/T
jU6Ak6ilIkuVQ9Iu6cuoz/azyyP6GrXyTvKZRnsQLv2apB3fGitC0+m27tU3g06W
5ER1qr3mgikPmz1yk/5Gto/Aq/8o5L0LQpbNJ/zkwnPToFffKDH/RlIHqEPkpTXb
HBySPTqYz486uLcT6Yqtk1dzVVA6wqU/seaIRp4bXjtL81dPgVUnrTp7/ud+CANT
5Oh1CJid1X60FKw33CFGqgpy9ADdR0E0VjUM932J3klKNBrSSWt6z1Xa+X4Gj8Lo
E9ItVA16Ngt+DbsaScIztPc0fY/uXY7FYVnJ+FDH1ZC2CxdIyhvTGqz0795qUSKy
P9v+Fv8Aq/V20Dqvo3JUHHH0eMDlsz/niUJmYulTVpc5ksF+ee31RkJHhv63DPWU
AlC+6Fx2bfEQ5izXeHKyvLsjTAW1H3RgpxuTt6IhT1GV6lqHnBta160p/4Gun2ff
bsRdSl2MnDZ6u9WqcljJlAmh5+7URd4PB6xyyPktqVICWLhZtN8rfCa3n31TP239
cRSie41Y39sSB05+PeZuvC2UVtBklfhnTzpIJbAc4cteNzjqCrRyy/cZ8nKPEr7y
FMyYeG13hzMpsUNTJUDR+TzG7wJRcTWd/CfRIoF9lMQ03LCV9i8RSP2IWUBUt3OC
tnO+8tOR/zs2a+8j1+zZIXKLnz2JlKTnyWML1a8Y9yZA7/Nib8jkRIGYrBDBl6TH
KlhtamIaOI6ALasH7LhMbqEs633p0sFP2Qwwq5xut5Gk+KHkljfBEMsmX22/5Mud
7ydiiGnsScoFpRczuvfZ+hG1wfPe5ERxoz5yqfBM+Eg8i/qU87e6LvDHvzAHz4PP
C0GlwReh7cWi0OrYMs+iQZdc0MbZL22BHvRIBYKIK63+vUJ2/7v6Aw5hpfzL1mR4
XaEGmTIZ7wb4SAjfhtDDhw7PC82kdx91npfbD+HCbrrRrjYIhOpx/zf0SoTYxkch
8Hgrpyu5IQW9xvugFzZOoUu0N1huR5gpoUXxshVpKPbVHnErSdLhGpqTz2HAU1ma
5YNtLRWiMxQdhEd/YECL+ckO9U6YJRx94iySURzKMkqZ5wf6eGW71us+jayRybC9
FBw8CXS/Q+0mQPTDsgqIIITTBg2zVU3MithimU9PBO4ycgbWzN03R2T7uvfouq3e
IFsMgTcG2lYenzgycgxniuFfCjF5KlEE0pVFD5bYhJ8vABokadig+gnkZ5AltYv/
skdIpO0tmvVWsCjMnf3mrzWLwDSeQ7onK2DWoFKtTu7eivNGd4WH2IPeJMTD9g4o
ArpcsCKBEX1mGcfHpLrJgEF9BGk2Omvj32x70bFPxU9+HrpX+nvGAQVuQg0CnHDq
qLoDMwqQGDUaYGm6SB0xSSj5qByJaHWmkmy6/kEUXyR3EdKcIytoSi0i6gy1MpWN
X5FlcUmYnyKW6HRdSOPosiMd8IsBluF6BdQ9hlMqAGLTJn0iUcFluppmkaRR5PEm
7Dsi6XF7zQMtL/8d0HR3AKwghvA2S9y59dYOotZsxRlTsIEl0zLt0Z9L1hWVbCQW
menwMQsoOmII7+CGKZ79oGmRVIf122vDVrwNRo3DEjpVv0AAwgE5W4C7zW/QqR0g
7ILJIUZNUKit5jD1a/0nH9YaBaAwjNQTIMVh6zYCuoBY15pEglz1B3+vJUsvmuE4
qTh4bXcGn0VFa4R6/9gNC8g0pzCQ0HAsu3qCHk/G3+SZK/SGQMxIY6HQd3s0SBrL
d6D11IOzDdVpD8fQN/azWdyuFNa96ugIGoXFI/elBGJxOoj/OkuwrdIul+I6e2dl
Y6SeRLvqKwyE/apg3Tt398bpuJ0GV17apYyxKtHyOI4JmUrSD21ettWQMPnMExLs
Z80Cmby3ia0q8qp1Lo4ZNvJbbqwWSXST5Txj/JHKYy/wIgVq47g4cj8YWIUJ8TRt
nRmnnWr9PcxbOXGvgobHrA2I+hHcUUrarVKGZuoYZBZNS34ExULZWfeOF5rLnRHx
5LuJ6VTiWa9ayuERcnYprRYpOm+SXTuiMpTwrMkL0ZcgOE2BCdj5SwR9jmWioVCT
Gfw5fAkSobJYcHcrxGLcRVBCLtQNKlbPEGPTGjhwiOsFz/5hP3uIs3BjeSQTCKEr
pUC26n0MNBE9zwcD5I83E+aeLnWijyPLcZ/w0KgdNxQICdGPNecSjC2qhA4VSapg
xKxZK9ENOAEa38Ub+dm9AIqbktfycDnKnU0JqphouH+p9QzsqqdDcNPm2Cb28e8B
pmGVbhWDQEbvI8CrVCfppK/H9JCELHyBRAvONKnZE4ekdXsGFAYZQTgMSI9/7sJa
h4DZP9fQ7emWQS4tGl6SsYruBl+TEMfgWehP+o26szB9rGKKI8O6liGzy0PEDmRg
UZRZKXPPuxUR0o0s8x6OXCCF5RrNfwiZhnEDx+nsUUWBOOH/JN/MXZurZhy/g1Q5
KTXwLp5kq3Ay2a4OEnVKjN/Zd6Q+leM0VLGqufvLuLa+D3TU9qnRtoNDIWJg748Q
YycAdSQq0ZzC9lZjzBz6olSH+vDG30uLHY1OEZQf75H+JAU0tkdXguM128ZZ7J+L
b5gHeLAmAkq6+eLrCqNprB+35ymmlU89FC6+HX6KIkVu6pzF/GF3J9ATHp5SuYxG
q75P+l7t8HUu5B9fG6632dOmB7M0/m+YpPjx/2N1astVITOB/MKlBmCfniiKxOF6
WgqRsy/ehRxM5MPGN2At7lMbuCAujTxZMwSgRUnHCIRtgTkzQag0Dgkzv6LQLQVV
FqvjgnJ2WER2rA7CsTd1eN7PQ/TL66efeZsLTGP9nWqQQ3jmee1lyY6KdLSkl03Y
WXi/1bLB4e3ij4Zb/YPqq7xjiEnuCWlsjpjTO/k+2CKkaJhKAYvEa1nBE/GIf5CO
uTrmO1Z+QoUjvGevFdu5LxyFozVos8k+2qXVqtv0Su+peeDg84wGIgIFhGsePdtU
U+lqRlxWaSUb3BJhJyLO6Y++lZVVu8fWGHUiYFiHiLx22MwrLaPtZcBZi8NbBmg3
Kbp6VlOA0zUENxpmteyTDduGy5ydyjvR73Dpn+NAKCV/7svG1p6RvEipxSb9E1Qo
tCrxGmAXgSJBblbeVUJS/y4tKsY6iy8C1VzYStEaTPsjekk6WlJzF/Lv1e5AftIv
Xh4cgHNz6ZP8ao14/E/8fmLogUIV/GQE1L9O2qqXiK+OBux/68mwwgZq4JMQZJFT
LpD5/nLRzSPi3xEwU25LGAe8I4HFEHr8CZ+2qLQoMvNonpmrT1RToYYP11O2m3+Q
LLwNpFEOriGbV9bXqiW2MwMyeZ+TcBOFyQ+MsIVGoLuFP28e5hcmQa8PNebemZXo
enIiASqKtHP0bK/8AbENzJLoZ1rmQuv4W2QpBGimzeKCUvgQByIzYHt5DNVd5FyU
z205hl7rXwxs4wr9LkDzNJ9pKbWLqStQiL07GR6pTLWEycs92oYJJm5CeqPjvcjh
/QQJGycVuaxg9C+Fcn+GkbxY0g4+0yv8lr5YBiZOJOuoUuantz9c/SPSIIFRse/x
SJuBrjqCbSTcnIqm42FoXTZBe5NewLIocmvaCw1OKp502T0WqLfnQsNRk95KPKTC
cCRWgRb6Md8G/X6WLQw7s+Gr7erAQhdnaWpgsvNY95DwLp88iA9ECS3jbTd9oYf6
snTFdDvvrIppYiak85Eroyx4JpfPInFXG4MxnPyZbTmxjcZ8utz7P16Kf3WLhR1s
0xi5GkS4I5IrTrz5cUTMxOVaiXi8NV6w/gxmErGzhLeLCKuzBlD0def7cnFCl36R
p7AvRCGoHhnPCF/vczuvfsMS5Ci0ER7TYZjXZZMXIf7KVe89F1323A2xaZ8jz8vh
R2c8EZIPYjWU0wJHU+VQihWkf/oKAFtMzAGBoqCishSFF4uVkjvCpd6+PrPk8szY
AYmvP8N2l8pyR1sE9Y5sk/zvAXYJruygZsrEc4WDQn90aWdOj+kMVBr7KBMlIVtk
1WFSHHOkiI5SC90iA41330fmMsHuM7yzph+kQz4CM7Nht7rleH7Rz6k8Ve1GNmP0
zz1kJqC6U20HHi+q/O0UI3K2GDUSPby/f1Fs2YQonQjGW+JsFXH43PzESPIIhZ21
5UDUheIimNTsnQWqTX+Y3qzMBaPo672DqW61rotxbdxApWTEXkzdMMkQxb66ueZA
oawYUr2/G0MZvl4U/ueCwi3Wb9qZfMkyVyOWzKBC1QzcGL4P2qqM9lxQTI1azHcX
Lo82X+O6PMXzQ4aT0xMFuOo2I3YkwZyDSmZoIyVOiV31o6y9snGBnC4bkHDHVckJ
2hfeVUQpVIe6hEgzN7bh5Om9ASQr4r61tM07gyi1DN2xU6YTYi+FRRTZ6m1MgBAT
jkYAVWhck5Q5fw/qSKxC4nxxYxyW+WapTzbiVxy1AYJToAQdOLtEffXyIAfhL4tA
GGfrv5aHUVwiPxqHdn4/PUuNY1G+5KyNzrb2GiwujUeENY3S7wU2OTPhfL6M9dvu
6gvk20kmFxlNZFiIr/ahXH1sgkkGT/twLYMYeQYTp1Xj1cOlUB8LDyVZapMx5Xjq
9FZ9FFYKmp16YOKa3EStt/r2fzrJincoCfsImRok/DHkk9KsAjWyUrSI7s8AbBju
O9koGPoYMHl/QnyqgQpXi+LBwel+EGhUenxeDIN9DFzlo0MmEmdIa4tJYQzeT9zJ
zLZFLxTy13lUCLmHr/UBpsBYHA52Ncp0opnCUH4xnQ7B7h0Qx+2azs3+FVd1Xitq
iCwvwYS5UfQ8tCfz6w302ziaX2t10HUGUNlHDq0W89J8DuTbRvqdwrv+GXaE9FhR
S1MsXMfgPvnc+1IjV0ekZPZilU7y/X+7HmHwQQ2OjjWkAuX8i64Xq3rikANelDNA
7Q5lxz3hRddgwW1XQl4anRJaDcCuIw0qZgt0PwGirp1v//fQd6nSAMWTS1dlE5QV
HQ7X46EDbZn0845e7TfDAKD6Ns3jHZzt0l5tbnPn1onEPuYapHuJ9UNQIuxzUpNa
H7QGV+QYpj9nCp/Sw7qC0AfaYM/7atEu0XxEq/zjHF8OCfs8SqlEWBfhtAVxi4HI
0NLswXtJ3+1wmf5X5g+4fWrUpSCBaxrcfCVINe2uXQOuzX93qPkq19ph6x46Xr/1
tOkYJ7g0ANp3vxucl5FM8YnYdDdGSJIMePrjC38yIAAdWYUansNR63poY4v39C7o
6mXqAiI5istqixS44RwmlO+RsePJncDTvXm1TXwkYSD9TmOkzGwx1enYWuIiSAZt
xYXw+0odPdNL4cgKryFnpgVLD8xbKa9wBFlca8N2YFrQZbl18YvbFfVbAe7P2YHk
JFrJQjnTq79zL7WHB8YA56qHTDaCrUTffASGUmfJG1Yqdizu6hKIFjtbqeNKgNIj
B3yc62t2b+MDLp82qm9HHkCLolt6ShcmDWprz4U3ncF4vG2tHIcfHV3iLiMfcmVn
P5RJf4oTwtR5/ZutHIhk/IBeW/ZR4ZEMUa/pkVVgOAnDz37/2B3TUsdTO0BFtZee
DwkrAsAMSK7sIVMOtpdH2+v6avrY+qv+46V32IRT9tDfjYBH05MsPMLi69m3Yefo
OYNr3MAKuYtI/4nne3aokWlsWkyW5IgQegiXaEAL6xpZ6fKdfGzpJmdke3+MgIFZ
WsQXDWp1QQZQZnoE+nQTI/5DpbeKac+hm0h4CspJ4VYK0Q8Ng+vC/GyfRfYxTJ5C
qTE7X5Hkgu+CNzQ8E93iBkOed8UEJZefTXy11Wxxr5PBMcZrASZeQwVGgm2XohiG
eYtVjmxZld9ZOY2M7qNYMwor2KRFlDjGY/pVLctqhKkIijx3PsTl9V/jYexcebdK
Vo+Jg20Z55+gCymL+P/igBgKQvANmYMfvnqqCVuSCntfZqshTsX238dVn3ju3dYU
YnHT8Geplgwkt6D5rgDlvul9Anj8kg5hweCwNT2UrRB7lx9ewGmoHK1qjP7jEQl4
u8e+wPhurSGwUHcc5WEK+oXBuIMyDq6mUC+Nw+5dKvC9xtDZnHZjZUOhXfqmAHSx
iAmdw1mz80IfWiKwVIlfGsQlHpQ1TP03RNi1rBL7AdugKeQkY/Bv17T1YrOjcMFW
/E0h4N/3K5StSBRKWhoMDB8EqsT8zDtdAaYNOAhK7U905apWyZwPMaM0X8hZn+IM
T1EGukpqNLjzecQREIXslHLtU5QAWi/0VcmfVyB9r5wZXDtdN91RMR3wha+T/Mqp
0Va9J82Wg4BA7anN1SU8O6fIehH2/KCXcB0EksyGMY3GHYCJzeSb61weLZpNbJYE
BpMaRSZX6IwUh1aFbhLvfUMes9yCgexpHAKv45j0K+tTlyjH/bCYH4VqMzYK3D+N
p/J13lBlhP0RXJhsGV+h+vs8Gse7f67urO6OsW0K68ddTlEh0aSf3MbT4k04jfTL
+Q2m4bgG4IXkBnQYpfXm5kXDzo6A4I5sYqIiwJ2abIUoIWEAoZS3+ZD5Zjr/CMMU
YEW/uOkoJD7Au4wmmYp7Qh7ZWQTOmbqzprofNZgvWZRbRUAODvH2TAA6SZj/+PoY
pYDcQgWbP0QgNL6Y5wk7CPCGBdCHREz2tOuM2VNaNZ7ZW6il34fXUaCWTgEcuidh
l/E/7Z5f6DSqea916QKckgB5VV/JhmAnG21dlsjYk0mA11L4sZivxPgNgmJaoUlv
j0sYYcu+kwR35kzquEWSvIMpHIrib/lF4PinK/7pUkbBYq6b4QBWQHtzrWmJiU7a
CZsj4X3GQxynkFWn8Ld3FBZci6M/fCgZb66xy07dV986FxG6pYNngjIdC1/ZVGs1
PhSDLOHUVAOU6tCoXT6UVoxuJW3HFOU2zLeV35PZXRym69sez+bvrpnTpvqgoxJm
pm33FVxJn7Yil3MPgUt8CjtByh8dEIbr1CcSKz6opB31gl7J0iGbg3NIN5vWdUWS
mEfqDJcRKG+bUZCJ96NMQCJNRv6LZ2Ara9p75O3zQGjiijCf4pE2Iq5A2Rr0BS4E
dA/svx9tvjkb7pEbDuNpJScWBwTd5SD4JHownRNG0EJrCPOjT4Q4MLEQnSo7fe1p
LyyjM5W0Fjx7vMlEQR7hs5gkn6kYkZKWsT7pWw1vK/GK9zbhBywPP6WXSigL5G9B
4nzUGAFkv7ZnVfVTUAaenCaTJomov2qHdExYgXLQxDfmdDIyhu4T0kdfQsxRqRNe
Zynx+DZi6GHeDm6KbscMJvZK6QrwJ6Vh4oCWnWgcmwSnWd97ihMR+BMnXbZMmADx
dFq0n9bdCHPYRarjRkPeXR3bgDXpxDPypzldU4SofoAL5zHI5VZnPai/6BuogF5A
gFuTRtb3y30uxkxhN0k9MpDOPjVSskFNiltu+0auwJ4I2+nUbsKSokAAUmvHGVVG
0KuQWrScEyGHA2I13dVnMBiaS5jSvzbhKqd8UR6noFsHZ/IWf2CkCDZNTDpN6Fc4
n1uvdgPjTSxOhrHmiAtI7yBoc8mB+SqlvG1TJd80y9vpnJxcqC4oeyDz0lJCuG61
GxoIF8BaUnSki+6EOIvYnXTby2EWkn0HOKGS0C7bCDcAqcpEo3Llz2lHQovw6MNi
hJOxv1bZWsDhKzde+PD2HnOmaSSv/WALbWx9m3cxyc1BKeBDNARY7ECGYHg+taYv
cP+ocH1epm9n3NcbxqBFOCUjkzMLlhEjXzD+Gx7MkbLmAORVCinI2xX47FxVXl8J
jhu0v/1Ny2nfhQ588ZzcLaX2gAYuC1FYN4wBI4v9g1n+GLXYTAhypS+a7v/3KBex
Ye3zRVtedbAQ/zGz5wG2Nr3/prgDB+/uTD4DPu6IPieAw6UNxynCAwRNUG5lnvPo
TVGv7+tI0HFZurljtRHVtWF93ictWRkBh++FdPziZO+jol3KFzLq+WqUAmFrA/vE
L3FO0HXnxofEkvmUKMEomn+xhZP4EPB3E5CtXoJaLrPGrEN1UyKQad59hE4Jw9z6
c4wf2PCcPzQfB8Ul/mtRt54/Wwk1Da3ts2ejAse8QoWvdQHjvjKXzPJvH7EpKgUn
5uDnVX82e/b0QEfPmRSr2dIGG5HC5FLXca1Zj8LpbMKuCFape1TEOYkOibvCT6BX
ndfnwFJJTXpbeutqDO3K+0ogeGpyh2uxURLLeb1KirmLCFjIzRwNg/1t08WpOT6l
UkYsjKgNpsLZOwOg2kSV+Y5vJQj8nGb1cX6xQ3Zc/plVjnDB3AmnjGUDgpxdNBAV
8WXSAM0cuUv/trqutG2CZ6B0R6rzJnHf5jad2aCKaQRqei3En+1s2u+gse4EY0CL
7pjE7BP4XmMwF4qETiM/HLMTj3unst9aU5td9HJuJyWaGqlPzQwME3NaxYGbSpHa
Hmjp/2vGEuvlUrIxExBbv86mbRiWmBDccBNtlj7u4ogvX1XPdwY3IuT57+1uYO03
BX7Fxk+QR8d0TBx3rLNx7gOsSDoNPAFzpsojeRLyxjmbQx/mZoNLOV78KpJ7Xe/0
3KcjNEGf7vzwmOX4vUA8qlssfUOdd8DufhOKuCwaLygUpZ4C+ccSW2UTsgfhxatP
ADfJynvyIICgAH3bC4VvDfsy983FZQjCtOqLHGTGOA1+7iAf8aAG3C5sgupt9/JM
2S8RyDUiURuo+RqMsw5RamXg75fHWvSQXUJyxzKHrfMUmxh/zpYq0VLFICWm1v1l
ckHMHCZysX+zMfiDbmlHJfI65JFhyW2keV3IX9XWsKA/zhjKVPIRkm3x2CyR49K9
fi1XBLBI7ux70voxn0rUZT5iudcoG6ZcN5B87c3wHgHRadgzOXEbJlpIqECokRlT
hp5EBkqb/nv26dGrp7Ttd7zdS67r6oaJUgxmPOnTlPdDH1ME/L3cb/FAml5NqNIW
6Wjxk5QKdSQXL1+PIW3U/Umgm/ne/bwmfbeN73PJbraMY0QLzHzxlDAYiXJ4ARvI
hw3iINcthk/dGmaSO/xb7jz7mWCJEz4wq+oc6qSCrVn6if+Ngr1ghtvc3GlkSC9t
zcBxSb4GoZ7ohPkTpiZ67arjC0JWAPHaIXIPHqNJO06DA+5APi4wkubNwL7OFXNR
3C79FiI5c1erSfp1x++PEhb2Gw+B4JidGlJzQ2iYggEzS8eMjgznhe00qt8ENRFJ
Rwis4kum6V27V6r9vesG1/uCgVaCyOWeNuBb53LfRbyjtWme+46ZvTH7R4sg/xle
0GcTR7biMlPD8x4OL3xsjWQ/3KrsaANKUD2NE/ib3HckI8OhXv9HS4urg+/CwVgR
VpSrA26u6wwNYi+7G6ntjORxfhS1OzFP0L42RK5nnavKjm7QCJ7eAtsawAl3gVv0
DkTmUA4TVR7pVdHsIpcu96Za1f26KO72UJPtwr2ePqoGnJ9FV4cm70t8Cy8gPP0c
1NMR7Fs+/9eoqINk5qIlchSekpi2XceX1/d/zIe1N3SaSfAqdqal/Mh8zX5vHpq2
kcy/q5Q3es7XAHNz1lrQVv57TxyRX5zg33/ycmqrRkPQHcKFIRXqrjDgL9w0Zksq
qGtQeh6ArORigPIkI3y+DtInDA6jLx1lp/J/va/goGk4WO0c1Mi8xTI9fAD63rma
AwBPxbFTl3bqsmwzW40RswrrySoQAL5hRdlwvEnjK4+bmmy6HF55FzPTRUmLOIch
/osCjjL1ro+AKgSysIk0JvrkUsnqIrVtCg2lpZ1YUPDvJ1Z0CN9FgfkXTvIImzPQ
fF9Gxk5ZIdurMcDOHW+7dhHvtjR+DMM6lHce8hIhzTbG3F++r344VV1RS7ZwyxbA
uoZgZ23ccMj8Dn791bIxlO421pYH2Iw1G7k0obvoNhMTCvycy2jYovhulHJtuDST
YgciZmzyUUgxRbJ4U8rNFlXwcPKTjV882sh3zLhKnpqR7if5VD5I8ALTFbsXe4RH
05kS+7rL0qvXhvKsB+UaGlu7F4zehhLAVSoSj58HiDKpTU93L3stqcixD0oluskU
fNYB8g1AqTpzAOeiO3HitZcJVdJyc2GIX1dRrhju2rZoEIDtUXQYgiOuRIYQvmef
sR46QTsJfEhpK8mdSe8JbZAR5i7RvrXFQpzBJG0uTQVK37XY3fGdG2pgsN/Tjs14
wn1THbK5RDcozWaqBlCuQuzLCQ1aJNIoF7CuyVu4SUahg+8NphAF6JSnz6emVdHR
YOm+TJER+R8MnERkgrNuq0wygqac2rvXI0JY0p+k0sn5l6UfiWkTHMjQ0qMFLvVv
oHkAGZYGZNn+s0am+KJ+qQsq7+Arpogweur9llR2ucnqK3YjL2xsmcwt3ra594rs
IXuSTfN2Me6Mqe0WIP6/uDP4c5DNabMWfmfFiAjIC8xqv+Gwht22TMfkknFjhqMm
6ngPIIgwLsMzyh++qu5R2FcZnui+hghBo+XCLzJ3hbhUq/6y9byMr1pzzwYWZvpT
HUWJZMPVgm6SHNpxgTnf6arTbe3XIt5fGwWxjG7vZg9SDE/eKXuNbBsQ3d/IP2ST
DeJbhUW82GZZhmjpk5cdu8EDowxnFI7BUBz1nM3UWuxURmfiqSPXdvSMIFHRjfTA
haQtfqpJpS+I21B1JeGdfTGnElDW+pBUMI1TEuLYI8DfOMbJpEcN5BGyf5ycxvwb
N7+XVtKnvfr6HSXFVTmsz0MVxbajK7jFGplyeuIoQV2QzfIXWRJfXVbV6mLVw/EL
aEv4N+/TFOqj84mUPJ/DibQMkuZxRLO1SPKfNo36/3h0Gg+oPohwBKt83V3Hra/g
K/Sv8YNnjCqvKHYLn3FC2UH8zGSKGph6XVanVM+FQdwCxjDY7x7JtXNh0EYSkbjv
XR59GsfRI/ojIvBAq/y2mv6/6dDUXoVszyu13cFS4qfiyQiJviwe8PAnnHURJPD2
KopJV48cH8F67YPadu/ovByEui/+VXY64GRm0GjNMKio3XqGP3yDphT/EGFtLSkF
U4ScRIQKr+q/cdc9Smxo6v6W1G8+JUN6hf/DN0HJ5joE1eL0N363vJ9FcqWR6OtT
ja/57nkEPO7NJK6xMKSMYTSSETRn/EV7VvA1FzuyC1qQVdAgk2A3pTm2Bn4qzUxi
w3SPqBCIJ0beaSCKDlEhbK3xrzAZXquI86u9ECpqn3D5vvB219UBh7IBqYOCcRjv
LXRAktEmCc1EfPb+6d0IsWS5u07lCUg/D5rG9jknFlF/o6gRTOxgF37N6OHDSbyr
HGygtMCBruW5VXxXjBwD3sfJZlBOiL1cDq1Dx8jC9j+k41Gpfo4YpJBQ8xspUEAD
ExTgi1Nh/Vc0E+l5bqMTQMP6BuQ4hLOtpGWXAYgV4DLIx0P+izSghObTB/ANd+ZN
drKt1kAtoPNtreEOl6hcSncufsVTDJDjNE3ryApVla7Aft9touz5LPKlNJRZ8rdK
+L1l4H+H2K8ApNJMN+7LEoWaSrcWeFlIKT6CPQOldOviKCKHZHqd82JM3QDwC035
YRLgMxZips9iyoRgaUqxvF6sD3bebTUkorOJR9DyZr0Rgpr1R5pp4AV+y5eMiBlM
LOArorMxuSgYM/Gw2iFQwQqXfbUmeSaHrNLL4FiBdZjPtQwq8vtC1ZSH2ENFJRFl
4aIUsSSkUNscOxqhfLLsjVCROG0xkBA+xanPdp8UX2RLAu9pzHaIhqEq/p3wzCq+
qAGb6YbNXEvs+yfoCcH7/vqawRjI1sEqsp8EAuPa6KyJl1cOp9BIRbsGtmIZ6GfF
1vb+TQG4Wj6BYe9g6tXoDnUIoHgI75c86QcuAHLGkfSkqGh7BM0jgbvq/w6W6shx
YhqVx92YulUg+AjRZ3b1aygD2EgYECy8AV4Xhk7tH4LVdGAtWpMRwez8U58sg0ly
S4eFHwB0SkYSQEOKgTw7pRWnZia3t4W/Vc6tJBpdU3BPMFIEXk2BsuBprqGDhNmQ
MU8HqwNEqAl0uICUI8ntRyaPXvgpffMY6DwW1BmF2STyI1ZtcKSxC912F726lRai
lwEFlb4KWizAuC0dMln8mi5YxTV3fsQhSRIaIm4oBArO7YBkjpJSaxDvWtC1ilF2
+ulYEzxKI6FqybCgOcRUyMf/+bv1tEp0+/39P28rv9C8UuP3j6n9nnlIseIX47lL
S1doLMinNTFr1xjFnKafh/11xXSC0BvvzH+IvSxssj4/+eLsYIAyiiLbvrOwA819
JFPBirYVDyojZyYpe0Ezkb6sQdoxu8pOungNOnrfmnRollxBx168vCBhgI2EthgP
vGw/IGy9uw1IrWYxL2JsaNDzEDYxoMqRtJNi4gQZCMTvK3KJOZ88+pAj4ijLzISy
ZxbNZ+NqY+E0eiJN7ysfZXeMfozheLyhDvZ0JEBIDdangV6rXe9R2q1ygCCCiq3R
NDr9u7lQgEJAEP4qCYKil4Udaa3BVWXDcJcnqjNBHjVWAd4Yz0PDrcPQ1a6mS9IQ
lteDolRvFcoqcDU9F2RuDsed0a6bXGNKVm75xAufl43WwIgKU+p9yAe3Th9KIFos
wTIg25plV5B4UGs6EUbxAf4IXLnF7w2w2yciremNu3mPZPL6X8dRRdcu1NowrAR7
g2n+d6u3vql20glDCJ0TclU17LkotKA2tJUAcBDYQah40zW4bUaYHtyqPsCX/TCb
sizRR/6UIwmhKD2hk3IidQOky704x+lEQOXX9ig93mbJusreZZtRADtvdhCqdOdO
4gY5s4UAv4iuHwaKYE5Q239vWdJAlHJOMQd8J8LrAZG4TX8t57ksRXlW4dKx9Imq
3fTiJGVMrIzGwB1vSu4HYf1zFYFi/zJQ5q3ED1oxsBDYIbNxzM7jDfzFgZ2WrrAL
TtRR1fLKIeJgoNhIWtwQezDrqR1+zvAHpFK26aKzZeSYcYcqTHmCbiQGUlx4N1Gi
c6xajnoPxm0/ErYi/thcSaCNvLhHEKvpQkysUUTYXNUSZIBF6deV8V3XFkzI2jJD
Z7B1+1L2cWeODIKcqM26sCaH48qcaMWrG6JUM+oAB91Gl41QTpsbq/+EUmNlTduZ
7l78LKE6U5delGI6gWRAWQb4dbW8T3fJbzfnAY2SP58=
`protect END_PROTECTED
