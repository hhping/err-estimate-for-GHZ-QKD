`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDCBPtkSr9jwuM9kWfw9+CntO0DHMoUgSJYKll2zjBptZWjiT4pUFoBL5k9cX5YP
MMMIoNIvzlfVoxh4lZOsPZf4i/T1ng7OhUkGzxvQo8V8Kh7Z1Z23P4FsVAvAFgb4
QobRrDWwC9XzNCZFeiXSuhlRvrpHTRDxB+GLwG7R7lb3Ek6L8V9heItnJeIPuKoz
xDlS2EJLhCQ+R0NEd9Rj2Xe0oBG2H9ngLgnnH3s8TE7uN2CgBgHkMDAT6wyDb6jE
o5skSbDfOD0g9oe/MeBap7v4w06kJfEo54EkaGn2i5OJv+8l7Sy5ivvDalhdendp
r1FhvVhk7XmFZDJFmNzTn41Io9tNgDnNhwyCQar4rNqdDfEEKMoX8+t+qNVfPFv0
aoZQ7kBZKHrHAsHLWwjqVQeA9pwbXWc08rS+ERTB8n/nFoBnKA7KYT4P75aID9nz
hs39ARdSgUdTWePD8NVKydhV7y3q1nQ5ckxHVBb0SCSBL6z6UdArDhDyp+XFw4za
Ku8TIqoGofIlAAcm89S1jZHLntz2NcO2+4j60+XSRRAPf9XC6cteLFZsj1lMPU7B
IHKtmAWZxHv4HkfdJ+xEfqvkTxibSh+ZMImmTYEJgMetP7fNk2W71oH4zY0T6OZI
YXr+fQGRGJ+Q80fGCvl+12eYF7nE/eJjuVpsirlkF6SXBQgVkKGDC4I+YWtMg64T
34Q67GGMu01Ede2EvqpW3WqDnizSpCAZ02YScgYq9qfVpnfL6eOvIcVR7jZqVAsH
qNSlUzNZif5vlw0HlkdvvjyeuPkmlnOombQhYj1mDnhPKJyRaMqY6QrfukSSG/J2
7d+j0TFpR5aGUPlsYONXQbsWrG1wIRh3eWZmKhQtmHdCvDv0tSVgpT3K4QMlzIsv
XZ1ozQDCiEwudMrtNHVuBdhOF5fA977e1dojJMjpSe7Y4Q4L6PpRco3HH4RA9mQ2
ikAhf/eGQ2r4iW1QTeBI2+1KOY4raaz0ZNMOawylcVZrdsqBsDi+AwRFCnQCX8Mw
jym4ipwsNya3lt/GiA46GiBcy48w0AkFjT3u/Wilkf+klC50P4vq2gkM+kwDZm3A
b9HUnwy21ii1nKQuTiEKwLuH6ZbuC9S4/dRpg1GUAAasga9xh3U83rc0FDzg1p8x
XZecs0fdQsSDWa2wcyZuI2EjMHRb2RpMP77/ZtlMoCNMs0N4NSI+xL9ydZAbSEvK
EzGqvSPGvdlVVUTQvRTaOcY1RBzE4G0SNtTHiHcuNPGhxsrTTcuEAw6wvJwoKePn
f4nvDlAK1IDTMaa5JlV5DJWNFBWroYrJoJ2g2I4DKN34+9BAgJQH5UEHmku8lFLx
7O2ju7ssI7gVp46c/KudEQsQ0ucdIK6mlVM6H48jUQVZKelt2MaGXQFfv62DYryv
xo4eYQA6y5UM15Fgk4D5BQl/n98sv3cs2TBZKDhBfK+SGR8sVG26jfSzKLYSjHOq
V5yWuRimOe3xeZIP04xRqrm3h1tkAebE8JoIc3HhO7nVO/iIF4mVco4DT1VKR+AT
J7ZDqMXMYq+TkqJIADdqUOqrWWYZh87QstTE+lxcuHiVI26dQ6hcqo0a51/s6z6R
hMsAiksZESX+ZfnS8klINoFGBU0+YNlc07PCd4+JUCQfpJCWpc1RPQK6jZJkTZ3M
LxiXrQ+hzhIJsYhiJGjroYV7Y898EQ3fnFRHLl5V8wfaImn3PhBg10oXOis18/Z2
HR4XfcJ4MkwZqConJrBQEXpCgDSFgENRzhwjmACUnLoDerLVjRgXhHMOA6yyrISW
RQXYxArgN2uUIpSsBz3musK9r5sr2ufB9OU8wWx78irwIY2IHpVC0yHXvQNnuAkU
S0u7I9cFhZAdrM9gI2eEKt2qOhL7kfKQ0/7rIFqlSRynaaWmK9RKuvyUp0K8DU9F
aq+3OsdxVLtEYAkRqXzzzbkCh764Qvy5e/32E5RPdOnTvh7OG9VyhY95bhR68D45
JymoXbkWZ6w1+BSvfmXvJSrDegfa3vSfv+bBShxq2n1PLXTEMDM61TLY1mgTJWne
P7kM7VYbx6iH2X45D4xjqXJFp7kN7H+FYIcmXynczCAESMe7r9CWLgSdpqPM7Nm0
vhVBHzo12L4CHpSSYeJtZJYqchesJO0k3dXWdtVqlz3XlcJi+OPjBUIGV8aCU9CQ
5tSfowFEwdnIErFegrYlKOxQKiZSYd35In5H9C4RmsjwMT1MTXrgLkmzsJgdXnV4
ZZaZMXkRwTR/ZRiCBCX5ms0U5tdAmDkT5vErG/ndTzpDiSkHd9R+LKgSa0KdfLUo
R0HhiKnzAi/I1CKtd3vqz7IvkaPT2ZxB4Qh8O8wdUnolpYok1euMEP/NojlNh2UB
DcrRg3NWym5opGmiabcnHmPsep4gVe+OnsJBdXSc6hNZc6Pj1rBCORk7K/QK2Nni
dQJQL6RAFTP4HAa1MCImc6idekqHTzxPMGEP08qwB9DPfEvMjBYv4E2/V9hNNbL+
SyYKsLOhjBWDBb2/SMecp/3H2f8mv6ZZjehUU4bJEFslwPDzXeOp0lAV0n2rIj2v
RthpV/tW/JojzvPrKfeJpSRGzRjAC1RQt6S1cg5pkTVn15k2YezAZHEnGLFmhtdP
USNHrU45WXVRAaV30yRVqJELI065UdsiSUeNXceSwXHcY/GVzr2LQ04X9bzt/vV+
gmQbQlfD9djVjXIDLBr2s8O287F6343mCqm6RInfHAMccfDsasb1BH31rZCoQEDh
K91br7hKCIWyWSwS9gHh7mMonzHtVWJmoBXrccQOYV8Rm7PuZWlzGUJWrtf5KSzs
O5Afv5aj80vjoj7iMZl9d2V2FHVPteAvvRSfC8G+1G6n/K8SySuYBtjfSe7zmZLJ
5JTZ6sxXSA+byNxwBervrHmT86ro1lY9iVGFLu8vsAbHB52rUiFrIVRd+MzpjP8R
P5v+D3Yd0bma71UlJtv6wyAWXZce/6gtE+lVmb66lxjCyv3HBNyO6efaqmbtsDsO
rRScluOkIinslQFPiu9ZKktfewYNOoL11/GpuaCMMOrkacdPxa+9JOw+xkxHBGvo
zFfOkijLaQ/m1XlJatJftmrcQqoc/spSHkrKVtn/r05XAlv/lfQ/LaCULyw5JGJU
uR4tx0PTAQC7h0Du67azd7aVDfE8LziucYOrhFS2H5WSxawx903QUJzaR9Jw8tc7
u9EDvpx5pm51BXpXGzSYlwuOALd9RigAer92/0My+cSUGPXMucMlFwWnY9lspoCN
8A11SGQl8ibwBbtgHhwArh0nAt4B67EgrO1da3yrjvp6E6r3Kn8MtmxxNY3bglvo
ymkF1bEQh5v1OnxBIuncx7gxzlYlWo7K3fj8h2+TaDpDvNfY9k1HR9DMfnZuFCz2
Fgf/MzumSAezip8/EwYAsO2le/FbwuI8M5I6RJxAoLr3xC+WHBN9AzOg0j0jpbAI
OvkGMxD9OxHKSGwvajY8OJZDcq3QfUyC3DBgc529mQX7JHtRoaVldJx5/bG8S+si
LYv4Thaf46jgWwQc/CJvNwnd7xyEsQIbof4BI6APYC39WGmaS32diEOO6yefLBZB
L4rGXKM8NAuYyUW3ORblh/Lc+p7pm/CdQC3KXxBbX6U8Duc1EanpCb21vldIfhOX
oENkb1VvG6AdCW8NJAfn5wgPsooCMFkEbWHo6hwg0pGcVmK/eFezceb/L4gv0L29
FeQ2T/fTJIOq3v992n6HlrWu7+Sccxvw+NCp5UI0DL1TvzUOHjidf7V4LJkOTUs8
1fx1HMfBcrF9JMGpszMOoq2XCZkw1bbdN87Qej867aX/wqZCWZeqf+40gexzcqWL
q5eeexYu1moqZbrZkkMyq7GMzfly5mf/+38YllOE2h9Be03KGStUJFfXCAvBjxNg
CBRnxb+PBrn1whd43bZgNndtdjvii7VlrPU6QSBcQwm/chWGH8F1auik6oJDZ86z
FgV4aCjkyNBipsK+qmtO+KgExZu0koUU91YZ6D2AaSWFEvNVZEui1Yl47v1um2Ey
/3Jw7uYO85TXN7IIcKiMMQZ+yDj8AFjumEonREVJ11Gt1eYqqc5938DLuMNDvhKO
+ZMTCQXXllLDiX+E4pQcHpKYGiZvTRsriqiz17ZvdSTADUYO6bdPAuHJ34NPWY2f
Z95JS8VMUSvgOACOLnx2YkmrgNHC5+eB9fzOzHeyI+9q+7Xr2XixxB/zC8Cm5E17
XkBDuiLZbrzg6xxjcBg/t2tQthb+lOl3BmblfBrkb9kM6bCE/ta7GdWg4yx7kIcW
uBNEuboerYrJWmpuP6sPbMVLgVNLgtwE9p6yywX0e7crAXKfLdvbn5xB6Yr3/bXR
kUdNobsmJdWnCiqz8y4IeZncc3bAqs8MtW3mukxipGYBvFafMvSICOei2h4OFt2e
5EsHdpMszxNsdp9QZEAmnMk3WNn0Et6FCretqrMLNAmwMDM1csqnKnrMIbiNJ1gd
Z/HvdgxfJX/bNWWefEq4qiXOq2DGoTH0lFJ0RTMlKDbXLn5zcAAAHZsWVUqGBwp6
U0nkfeiH0Bsswa+WgfFuDYHR3hfRcZMICDzp2cvB9RDK0t3SDL4vviYOTS9ey4bJ
aqP4f5SKu8jWF1kWKy+VfgZpyc8pJiAQcqzZ6QedsO3OFS5H2cK/1VdwLiMIAic1
CzzRYTGqtL3Yiglw9s10hLAv6rVaauZlGscjO0AafT3JWVnsb25ksgZ7kBhtvErK
Aupx/cyORPszoRApaOEOBqQuhnj6OqU7rEI175kK/bFpfGmPTH68SQx1+5LqbOTG
gVEjEgFBt7iFQm9sMbxUMjSzOhQsJEqhz9CdKssRjLKDKjhH2u/0Fi0k49arAhza
2oc78o78CXO/Zxo6nFIdUma0xSpGewRWOUaP/VnHy7uz7wcCM8156p6jr8WQy0Je
45CiJKpKjVmUY+3bomG4Rh2rPtm1Jbs6KOeTvQsXl40qCYYvLtp3jO0Kim5d1A/d
yoOJkiufkK7Vg2xUK34evS+RtKWQh8PTpdJxP4HCo6nABAfQ0YlQgvG+6lTrSsmv
9mjSjJJ/MbsJaeGUOIf7sb3DIjjlOIYPnlyLP7zxU3KYEmFJpgYr77N67EaGeqhB
KkHXYIRzwg1YHe1CSgHZBi+mb77syeoEsGcLyJxxkUF9sVuEWxqqHaJ80+rZT4wn
GJd0BhKH24crR/MCJbw6tqC/j0g1X0sh4p155UeslUh1JXMmC0G8iHxhJdiC1bJP
SiTzR4p45i8+4MbypadPYRNtXuUEg2p5We1gRUzqg8sP0SpFtl/vRJ+VFgvIN33u
AQ5T4AiRIqZ9tuuqp4TY/FA3HVryPKdMgBDnN6vtwHajX94JGhHx3q8D2SO9cXyB
SUCm+BIc0K4gi+8b79o9ccsMs0xUYgZwvrr5sWoOlomufPSrVQA7RFs9vbnLsfd/
IfOwgK6K+dNA9idANEVXqv2FN9AX2bcwmXQ6DEJ5KSmYHFjaUoGChZJiUVZ1HGD6
epeMqjXlVExJ5HepynQoko8mwfYYczR5F9ULHnWIFg+kSgNjHXHiH1xkSwLJZqEK
UXFQti2qTqxWtrxV3VFxLSBh5QsphsdSswFQFMZOE1EB4sVky9na36TUR2ccW0p/
Qo3UYrn76CtVeB+tptjzudljt/OZtR5NUBAjIk8xAm6I/t+UgdQAwg1hgCTrxTuv
VZH2PgUf5z4y7CZXD6VXIz4qTPV7ZzoPtSYwjh9u3o+xnLNN9NBiyQHmK0IjCJcM
U7+StZ+yfnxa+EDSjZeRH7N2Uw+LtSSw9HpUpLW3N0E10GaBlo1K0rs5frmz2UVI
0mTizutXq0JogO8IzeCJgAVZH0pmpoad1wDEeY8QvauukCi4KLurr6EFjnG99pHO
jIR6qBDCVjiCTYuDu5dLTOc+0DN9IvnG6x5Eai3epB7hXKWu6iX9yAJedMWLFJss
w5r6W1qpl/jeVV47ECWE9z6SVaJ9II6T3IhDsD7Atjb7lqKLi/UjUaQrzHQUre65
keahxOpPE97W7cJv5a2BI7+110aDjNKlm3QT6lZ6hqsqFAb0pInHyD0lzV2Km/oG
QSFncrFGyyajYfufjnf1v3Nd7qz1i/OtsKcHD1AS9NAv1OI/hIPrI+LxN/pRlwfl
tNfNf4CpK1VRQQm23Vq/7xKt88e+dl6wSPkJG2UFl5hV3eRI/PH5p0wQzilDbnM2
G71HucNkAorlK2LCtTol1iLK8QM0NA6THKxjDW2hPETXQAx3BBrQtprQu6nr8Y01
NHltOI3hACGOiRFBGBSrzP7pf+7azzUY7GZvnIi/9WP9AU4NSv3Y4RoJtbzplWgu
L3CF/uS332V/fT2kxn1Mq4I4MRQWxywsFI62oL4OvYvLSLKW6KyQnZ4DTuqQ2M0L
05852/VzLjZOgvjTdm7PLkqGXxleaA7Y5jRk85SfcTzdheaW0a3hAU2EwtUHbj1n
OzbmfhZuGX5wvg/+erIVzdZjTBOiuMu0fWTt5wZmN7KgaIZ4GSziCT4Azh7/ZlWF
mlwS2tx/EusUtjKgxKP3v5fZHwH36ZB7ZUljKoqlynXd/644VCFjCsxhuxH2BJiu
pKzI25yXxjepp1ZY8pB2BCagYreEVLJ/Yig0M7DI4tH3QlajOQwpJc2Avpt6pLEG
THHsVza+MhWsFhF8CkMV7h47e7B68YZBl/YGvWliMXuTmki+szQf5el2+58nzujd
MMBg+RTNGD+0SgEhGE6SH9n5OgFuZa9OSron/i2KiAKxlrtNsoP3HKVfgZfMDRn4
avoHD5729uw5gV6wskpU9KSFsAD/DNdZBt/oV7BYHI3I8+QMOE76ePYWTl7+y4fv
rvEB1XzaYMEX8Rb+kRURqoi9kRqAIwXdtDHWfDUnjzGaCj/Hkbc3P4BAvIaB8aZS
A6xpkoSWlGcMZmkxaTuKwYyQAUUFrHYc7CYMIDDFSCm8Wb5xwlXqCQMef2gPktAm
EGWkGGNh8Y0Mh7ndq3o6Jjqzz65rfD0/8om0VboCHguVMofUsxs6wouHAgeevBi+
plwbF1HvU1vg2Qg+xQnAVwD0cNwllmciZXnXdp0ojM6yVeTI49XshXgjUZov//ql
2vhRC8KJNL8oQoYtd1tMWH4TvwTZEeBQ3oWojheM2tsTLoAx9/HiRaJoxscttRVr
/GATudfcoTjU83CTJrGN56vQLw8x8/RmTrAxzBSCxozMMvTgfWPqJL8XzkQ2L/6Y
q9Mcg082CUxM1HGqfJbIqcF7mks6Wp7freCC1kKI3BI9yTrJjonF7taXVOZ0ajI/
twuutLzmRbG7ou+T7fU6KnMWuKhuym7iYXMxbD00sknPa7L6z6MefsSl9DgAcLYi
mXMGQ89H40XY2V5jwN7uJNBWbV7yelYW1ivn0t360Ln/VYpEHaEvSt1coaDNsHoK
ybAYLou9ESGzkY2UxWosABqw/lkpAbWFyIxgvRdD1ZH6vtzRiDpkL74LfpIIPXuB
rALMLhddKHG/K2NCndjyacNmuwv3S1dqWlpFxi6prRENMjtpn8FnXvPcOjg9Eayb
IHhbthxYX6RuUliA4ghqTYVB1ANNfowbRMYpBluqqfoFFunA0E+7yzDn27TKSBEd
B2Iyz7WhoQq6iP78xWBzn1BybkrG11x7WFKxeVPB1nV5io9tfIZNLMT/8iam9lH9
mQ+dsVNjRswKPQHUtHIi45bu+QWXIJeT0nyXPcgcRtEEtFxj8V/wAxng/EppyaK3
k4lMDppHKzbqvjoQdtSE5ngDHj1C7h76mcFRWT+c8oEfPYRkuJDcVqsxf+IvzHKE
I51n4RGVTw25rlsVLFkR0NYpS2j9ECNXFOsBBIkepE6IByIYZG1pP0XDvM2v2+la
AMJijmlTmVZuy5CJoTAycuJlxPvnue/P4+Lg3nRf5zy1/V1vLhzVfwtbWPsqnTSJ
zT4ZgaQCerQJMxlMtf1yCxfOfVyI068gvGUTCG7NmNmuEKXFJrrYgYBLNHOGeomt
2k98ObkAFJCDmH31W6znctt2UnwKie/71WJrm3gT8PgSNkGDaMyODxjV2u5ZQcan
Je44CBrlUYDTMbOD7Im4aGxhR/7LHzky/G46ix9PLqFvyoWm1GuSgvQPf3gBYVWk
QnhD5oWaGV8ZcICXRhdFUo4gF+EK+1z0ycRAvGV1UtXOJg+FB2fBq2FwFgJ9cX6U
vvPOY+1pxCnLIin89J3QE/e5VTc3J1z45ZKbsFO0UkduknQbp4CTT0d19NysKpQs
qTJ/qBAvRYdCkaHgRd1B1B9xz7y3DzyS84Gg9a8WNpCvWqVWBnDdjEIN3mF8cBgy
p4N0ZaW8JUdHkGttcMLsSsFtQtoUH5ElmdSTe3s1KfIs+8k5Op6Z1NNFAqNmI2W4
mHeeldxcghLz1VnIPn/GMFQj9fNHE+RsdeT38Gh0Fevx1ppJfjtw+VBr4Mp/pFRt
6ZpQz8jWRyQG39UF/FmBdInlf6Nk9QMaasz1jx9myuItojREg5k+K6nxuOqkJ8Zt
vgb3nxZ93PVU6JrZqGmVfrfEBaIXTMN+XDKy5THx/ciw/29JC+dr2Gy2qm8wu3PY
6JqNVr4aW3jvo+ww2Bz2s5VgaNTdQC2LzNyrPqHALSAZFfcLBML6fXl89Xg9Qm4q
PR0Cjg9ANH1GS567TDmJE2U45pUjGpLODioTuPEX9Or5WaSx2ECnZlgfCSAarZno
UUoTSBCjkxsb1IxN6XUSGe2WNJ/AX8wyHPUFvan5gdYF0XaQO79VCZMkyqPhEDSB
9cYuGwgEN4021O5dM9ALzAskSDApxNRPyRb8CgbWqy8gjWfEVvLghCHVjFXHYE47
uOCfdsVKPZ4Jvu4lLZ8vN3tsdFBpLA/NziVO6+J09Fj4lzIyxgoVGmJsdDyX0RU8
jhjGHUK1YzqJsOewdK4ja6w5b9DBEPBevmIv1Chgk0oOU8DrGuqjwp9J0lR/ldyx
p7cK7fHrPnRwXb7tPbqvlpDAh1s6SPu3/Wf82HeH+FnJNXPRHoYPAL2jnVd+66uE
ietkEweyiAqXgwjKMMD4GWQ+z31EEqtf05qXUY4Dz0x9d03JcakicTgJQY5Ay11h
PEfcBYXGbnWmaDjuk+9JRHpWf/mzEjty3A0sAN0P/1/aZCI5n6e0KbxwB8iorOZL
2cUl7YLhB/uNbpaIHzrCAkIPfTgDXykkHYnjWbwkqtNep43drx/hVvXTLQIH4kPl
IZcPnFI9JtvDWARmY4gONq7WdPh7hEAICLn13e63ZoVN8N5tMvhyy9RdsPQr2N6B
N4aj+Vu6akNCzzYrqpVSgorqRX8f1d2mCHMMol19cVrd/xy1U97fjndcS/ezhnOV
A6TdmxI9a0PLOnS15vdRJVEHOw2ogMxUjZTHuqpXx0eVeXjqoYq5Mu2x89vyRCrI
NJ21BISRQxZ9DtogNwoDaJbQj+szIN8l2LFgBecJtrTD2OR0XlncrAv498X5pH4/
w37EiNnmkoK9d78Iold2r1bUcUi/3n1BVlaOvnX+qd4bb9Uu5XjqG0Mc4tEDqd3J
GlSvEd80fuP8iPPCa4tWruVlfZT3RFsY50Q0azuqNcgyouwGsY7xOHphI2LVcvpc
2syul0HJuH/b/94w2LzTVdR2IYAO80H8/MqUu5FT6HcxEBEVLHM2yiLBODzhSC5S
QbTLy/HT8my00EckaCib03dyst/KgCVi/LXLVjc/B5R6Bic1T37zi3SIhgiEYx2l
MiFhBPuuR5dgc/xAsHxxHqHxtSlplCxR03PysAo0ioS9LCrOMp4bs52ZXpj+oNk3
XozPNtby0F7SXr7/r+nBFw932ZPBaxDGVXaNvmxgunhEPuTz4ISDUHZSjOmPbtNb
GewdrrI1EtXWrY8vwvbkx+S2u4IJHszQahpCTRDTOjIvxOZKofy1ArO4IBsFCqSA
+ATaM9g7zFpTcBsh1TSZxgoYae/GBrpsZY7Wqnm2C0YuZiZHodeAIPu+JwioX9az
EUR+/wfTuqYwDUeS9/UnNGFDOE6p9Vz0Iu7DZWPfGicq6K9FZtOV4UYbEzZq+pDR
UcFdofg9uGnl0i3pbRChg2/ub+7dU6KK3zYDLMnuoT9r3aFFu8GC+WHaJYdt+MC+
+AnfgL25aFViBmgRG1FPegfgv2/HviY6BFB1VyxeX0417mIOQZH8zxRood9d89O/
`protect END_PROTECTED
