`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nwj2uAwTgNEWl9llWTDV8Iv37GIUJ1pOmZ1YZW5osytA3gJm9t9v62l84/Bse7xP
ifW1EqQVqH/fnjefkR1UEHEa6UZwLCZa4pgNxgoKr9tbaRFVl4wQ4R9aKTifWfQy
dXbuZw7c7FUu97HXc/iS0v9Mo6B8JLgxNyC1SMpsPjoS0tKgWpo30lGNBlC7DI3D
75JEJFPdacxvasYDPZaYSHODtsO/Ue3C5FIIOFdTPDhY2bcMVJmf8UF2lkmRjNJ0
HlUm7M4GosvW2PAJJZCCnKdXIiWOAfvx9b2xytfVchTh55IDeojEZSpZ7i8Cy86y
voRfsvBOaYpJ9PTIeLg2Hr9m+0PM0NdCUlbwXupyKefiL+kYt9No0em79F20Jqq/
hY37DRY8ffs4AtA8a1kD8YnQBRx7slXFQzdASVwPBwGjBB9jOxM5z9JizCY0YQHm
18q3u8k4/BvIe6eKk8wOBqr2s6mzJQRGDWTwvQ1mdd6vhCyj9oLp2BoaahOMNAmx
pQHfOq4tKewvaB+0CFwvfDRbCdlERQIFrCDQAVX0Ld9+LybVQHClxoXJVNobRCW+
UgmHyIGl45vgteSfx/eKgGO4h0rnexCGl5IHqc0g5dV+1WJ9zAEMnWAYmZ3wA/FZ
ci5vsd783O7nBMGG3NVZrQ==
`protect END_PROTECTED
