`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVUyUBLcYvQdpr+GEiM4PUBwYxGu7zpOXU78iO7cpD8VRXaEWV4VwpVxPvOPkUXu
sbQWMqAKfni4i46C4JEA/wvVe7DqV+bHaiZFPpKzdhzcgRuaaZmgpfp4CrcMnV3i
VPNEe2fv70YoLUoQmkKofyZldWN8VBxMYFsk4tzZ5XD1QCwz9Wbw88ep4YKaAKJ4
UkWcyrmqvO7TU7X6ZAKASKJMhGFGf+JJR17rxLTwycETb3UGCK5MX3cYwkN2VAL3
8+UEtwQIwkfGTTjYbh9t8eZQLxBH99sIY3YZ0hrJopUd7fxk8zoeWOTRsVoRaHtl
l+sa7wsjOBHIsCHSYS/keMQAa379yS63+ARfkk7sQZmglHmQaBsXv8giQbaqlqiq
Zm9i166mX77z71M5mWvalKTceWzNRCpTcyYI1FMz0KgXnU+34jDEc3dC6Bry0xgD
q7BYFmfrFbrsHZqPTXxSPXvuya/lqQoUkUHsae/WwoZY1i13vhbsf4+PthowcwlI
e/+MCy9AsqXkGPqT7Ik/7A9DBdDsU5uZ4GI1bojqNWNbj9/1wp+15Y4OgBm9r3LQ
R/twbuceaBP/C2dTiS7Yx8p9+2ait1k3YQ5saPpUSTRJ4KqXGV9LkfubK3slaOxb
LNxrkRKPvOC8eceYJzMxbvzVLDHnLcPWQwpLQF/u8AeMkVcJmMmjQnLNoQDU/6ia
`protect END_PROTECTED
