`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cgVtT2e35nctPE92JBZU1oiJjKYQSaVWQgQw8h9biBusR6Rj97gDeFJRvIZDJgSU
VE7+b8b8SKB/y1vKgN3Ikt0EdXmktJMdotwojRo10BRoB9LOBt/Qr04CWTgJ5x57
fxsq3kVlFXuDCh1/lrcZntzB+swHaiyqALjItRfY9lFmIdVD0CbgQzkt6Dcf7Mn1
uyWpUzMcK8UqC7qynytdH/aJXo8BiOzmUaGe0Liwa/d2x6+zU8WT3CwPCf/dQOIp
`protect END_PROTECTED
