`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RQTrUMrjJsF+K901MaY1yW2AwlckwFM6cWQfcofu9EMPX6uENfAINy1vvpzhTsc
bPmaOO5phX83Gi4rb/7uy+rpOR7E7HDufMp21NIRGEL2N90FBv2e/aAqrSjU0EvY
uVrc81elDDVGqphH7O236N23wwKuZm3PNoaZYSN7z8Ad1KYRvVyBM4+7eurJ+f82
JXF8ljyq6ZZlXObGFe0aTlQfKxbc9GrysBCcmcrKTW4IFXva5AH2FTAGz5nJceC2
lXsm5Bi6SH+1IZAlK5DrFgy071kH9q3dmNho0OVlH5FFzwSozv4GdSyztl8SQrgZ
NYtpomlw5JYf/IeC4zd1pUldJRsbxwIUzgeuRcyRG+gAGkmYYDC4GJO+OlBYpKW4
0cYPyr4f3MyHcBzCkJEl9P1cLdEhQpHtBQ+wSiZlZGUnIQGGidDfYoLWEHhTjwyH
uyqA9z9xh8Y51GSnxEIuphP2qFdbtHcugjvfdYhmvs/WjX7LxKPEpteckw0GcbRA
kIY9M2fSAOa0+waUXasT0byEegZyyGUi0Gx+gkQzljANN8q2e2+nLL0aJem9/kRC
`protect END_PROTECTED
