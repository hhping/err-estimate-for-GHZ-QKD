`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncfvNcOQNLmvfL8vUr2g/K/Lxlh8qzv/li7fy4xsaQRn8c3Q1rBGi63GumxQwbO/
hzOe+N0Ud/EtNXalCgR7dbZPf2pD9HO+H7SH9AQ5utgJQ8ZSYMXcRnms9n2AkUp/
N3sX+C5PgnlFQIvzzOaOj0vG7XpVBZFcwKwy/YSIXiQs0xqPcqukbkYxQFV+pgUn
QqE54CalswEYobjIDlz868tg9jyoY2OeSJDFCywWFfRBeKYvj+7J/Sd48C9NIdn6
TvGU82/XxpOyROe7p6crRJLLLGkClUqQQhlGpMC00y0nNAIEBA4HHlp/x5MCvyVp
x+M0lvz7+sBKTwP+6w3gcIIeeMDXtHqAxPYE1/mzWwJ7SP1jJGVDDtCQ0sgKNug3
sZsW8CNxXUJFl5/xXTWn30h5gVHTgWVJbhivX3RVF5ylAzx0PRdyszvmuqcnNlaw
sZpxvTAoT0JiLz71sUSTzgE/Xwy6IWfh0nzqOMINfGsxgVcJeopeoH5Apm3oV5Yw
rMKGrBHbTgY+qmOfPsb97p/ac7WOZoUMIH/vVWFI9fDtL99j1IoxA6gFUWobYL6d
Tn51+0NYeFyHwZgKknYs+vqgNXCr3zBxBdjfGAuROzeNqFSaT6n5zkK9XpfjnDNU
PeoeGmKTT1cY6837IUHIQeMnf3BZynV47Ch6hZe5BiLtEd6mOMHj7aBlMjsXZpRf
3Iul01lJ2ZJPGIrUDbpkjrWFP3jaMV9yWnhzRU00+tlKCZQsMMvzaKwXo3zchUv1
y9IRQlU26ol4aKkr0mPLhjVXyNdlKzQsiCZeLSatvMF+UNff/EMAyL6AGoPi/UCy
UFzOyhmJK5YJiguhoI1SIXP3DqObZoxLCANOxPxNF841ZQq/gJMKaFvjyyg8fLK9
2vblE1W14JwdSbfQTgngvLR09lg4GN5bJwtLQYxBuFrbYXqYa3F8nFuXDTVEID5x
6046ua5X3AvKjliYFrcEqjLpwmQ2vxMYKnLFVkeWJ86dPGSCnGnW/aUNMJnBTU49
zM2qGZwkRAxtYbCbEf1AGe6dkUeQ0/HdAy/JrGKQL45/i4bq2f/sa5TdcqZ1SPf9
iV8Lm7ibI6gkWcNymKfl5FR2mZyaiAh/iH5IGj2Um2ehNhJ3Xl0cGV6zoFPAef58
yAfMT0SnCqQt9g8rowOyvjMepd8qXwRrIUflC/FR71F0ka2rNvAU2/ghh/Q2F2Nq
FRDzosxBpUpbL/1ANCsk2MLungVo8d6X1zlljtyYyU83aiy3BDE/ZZ+6qoRB6Zbn
6CuX/5kvUmBknvFp+YAfeQHxWDp5U/XCMBvkb+4OehdPeNf13FPUvmDhaHlBJsgD
XsATlnGWyUoqvlXvyuvb3ugFuAnF2+CleTOGaSpaX6Q30u1MoxthKnjjX1c9BFAU
7Y54yJ1dGQMTonsChMPLYJkrNbPlStzwAmPLAO5DU1riKk4T6KZh5xs/ODim36BT
m1/E07mgoqkZ/aZgN9Jd8H0SWF4JT5ZFbXj6zakYwjLydGTZ0+oNWtZPTkyH6dRH
4gq7Mrl2Pzhh+ZUEKvV/K5+ckcEsLC0V2JUDzexiP2HW7JndEeUxWwyq+dgIy6IN
gDwTNrWxE3hoBfE2spGG9okUQJGW9TsgfO6PuD06PZovvLBACHSag5PwRgg00u9M
Fsod9n+7EvHBOpeEJ45VihkKF57DUuX/tbL8ALcsDxuCVRbJlG+0+qbDRDJJ91QO
nFIVfEMoWGTH+0HR1BHFboGBJT2lQc0tDRKcOg5mhbw8hMPmdG4aQBsZDi/tztvb
rEGZuK5ON5VaDV97jIGCsYiVi7w6BcOV1AfLkNTPzgzt3FaDzTEy75xdSa/OJb4f
RNiJpvRXTyTKH3jT+OnPP6YUhZ5j+VWemQGLVlFoJiWOzpA3KirV7yfu4Va0WYq4
fdhzjweuOVAvxDnq8pXo/qcfiwwVG7ekXQhXAWgyWcIGKqvnROlREQtx4/VIPCFq
blxMMKx4XAH5IzrgByfpNZnKqkSRALggAMA3RNNnHdJlc2hOGHSIhhOfcPGm0Sjq
MMxLlHo7GDRLgVd50jaY++1cWtPgE2KFNafAvXgpRPBMmaAvRRF4sxh5X3h3WsDB
cQnfU/kAYWDGO/XGgGaIqakbB1sDIKCL0cbIb0KfApmlJAFMwEP+mYf9m9kDC7ti
+eiHX/QIgTB55WDxZ4f9K48aO3nsX/VWyvYhchmbZLxtbV4MbRvCjWwAkWnez2J+
Myts8F8gJMdasafp9Rea2RnQUbnZGjzaW3nfWbZAd9iDzhktitFajhG0aZvy5Q/V
nJmurb2xhF0RXQ+fa3zAj1cI0/HnzlDMFZQBxOuiRwfSx8C//v3YVcaBv8owE+nh
vHXflGGAVnXlA4PZFinGZhpwoeVSxphGu81dcbRI4alHbl+Iwy003FzVSadG6/M1
FMnZd0GV8T7Z3y8cfu30A3RFHGOItLp8CIbu9R7RsWS7+Ypx5IPsg1RKEdhclA4y
PANBpfEU9vd8XaLeg9mS9+k8vwoC1B6o2vG4j0HKJdQOp0VqbGQvBRBOtxruzvst
UxPKtF2w6Eq9KAEgeanAFHfCXmyQJG+tGMjj6CCB/3PIedKSpRTWNha79P3YXCd5
wcIwexLs1uqJ2ujGXuPnk5qEjp8gbz2qc6rfelZ7St760D+sMNF/tWAuNGpVsyxK
0zrnCbYjDSHfPpvgslaWS6qZSmHhA1pwHCuNg7D3+pyAgngzjXLxiFH8Nqnj4O6N
NLrmh06TMkBakaxYSi95CKk4z2jXJdQRCN3HpKxoMRGynZiTyuGK6JG7bcY3xlTU
+1z/FxVbIecHiuj09APOZNHPfsPZ20JdDtSljofD9C7i6ObCCBrs9X7iPLBsJTAu
12Vei2b7A83ZCPIKAjKAWLdkxP5/jD0KD81LcmweRDwN3YcxmhHcCKk+92RFFqAr
d4wVrfE0jwHczQlDRaM7HQ==
`protect END_PROTECTED
