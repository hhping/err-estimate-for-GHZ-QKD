`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zGkPNffShFf06LN6d+h9ktfh+KbA98xLfalaG4wgv49Yd4yzKFjjw5GdFhM2GAJj
rCBTOZ2FXVrU9SxB/Y8qwxrrRKPcxUdt6obyiefn54ZpRpmY6/X8VsrDejv1rDW4
ELx4+7ukvsLWTxWaiAnjMIK8JRScJTW2XJtDT35/Cox6TI0ETgucLuYMz1MgEs7d
KORGCjhUis9BkeziHLk7GO3ERkBYXrBOR465KhqZia+oTcwoxp3HjbZryt5JLm6S
kSTu+CR6Omq34GXc5rUwiPQMNZLtOk4mBg8AmRTk29wnStW8Lf6GfyU5t5Zg2V/X
NMurtw6HXOrjB/khmeaYPgVf3JxKV2SiDs1YCINhj5xn4kE/MQ9IIlfskZuINbvv
3AC+WME0/MXoHn/6SZOv+tbvp1ctsau4latTRNTlfWqW2Ehb/+ov1sYx6mR+H7fn
jOtg2DyC+zTrkoAKUwFo8llPpYk6d2Rpc+FrSsldNshqiDYtVfOlXtBuT2pUCxey
+WwdwA44xEJib/h3SRubZ2Ba3TgneGa4pAu67B/Iu5R1HMx/dv3sCYhkxOwTzlpz
VFHvFZp2mVFoKSmLZ/ZfM5u5hndyvxHgBsgWdHlP7KiloH+dWcFpJ0hhIJ2CndJ6
Xje79CZeT5pTfiwg4gkDcoNcaF0+wKwOO/XGN/kD9D+bNyQLt+D7Q5iBTiur2Wli
39rxQZ+LuLF89QfGa6WlGoCfiQ3cKV6Gr/ZybPw8RzxXxiHX0sWPsGSb+hb48ata
/bYY3WQbmZzJGp9uinkCTYhCL2yuhrM1XmfGokfS8gv48EF47HDSfTAt+pRAnp90
cJa2m00+DphdKbd2wgRHxhBgu2KZEgUv339fL5a9sVJ9T0sV9TBLewvaq1tkXOIH
tYaIg/NTNNaZ+z5obLY+s7ScwxJVMOdZAB9vffJKgiog+iwjlk26m8UJLpsp298o
3ZEqtfJEdKU69kVHffc7Te1OLqaNXJwzu6u0F3gtfHyypOPPmu0l7Bb/MrCx+FPS
vW5vLmfcP28ceG5YK8aAneHnbV+fbxA1Yabxn2D7q8HINzK05RXhhCgssbiaCTOK
LtyF/KYxQEC19VxJJEcL3fFz3dcmlxjixhOx9bmURJvApiQo24bYYlFAOVuQefUl
Y/WmvCXglZYFKdwPsRZn81uulo7CZrPnvAjFyb/GYUaCzp+jnCjz528RPIVjy2Vb
Qyw27TknIt/fyobzY+etox6NHRMHvM0egktQpaTRfsMvcSJLnOnqCJkQ37RnwIyl
HSFqeXo0nqO9CyG8fk5zUlJzhUn/kD+SgNkx93WJ2mWikdDl7Yg7eXDZPfLbLTrg
3J2/q9/h24vIuur2gnFEaX+nhhYD10rS6Hq34DXpHbXFzA+X0XH9tsSDIfWnDI5N
U6k5oE5qsbBSLGoID1vO7YkUXz5mADu9ZwiFmu2d3XTIhou3lZ+rEqbydc1hm2gL
x5jqVHQ35RtloY8Iyr7Rjoxu9rbIWFhsqI70S65GQQ5MDeLe01XLBNY4k4Q0S5gq
BLeSZY9xm5yVgqFt+vw2RXoEO7FRWkfG+mLv+7+SNxd4pyVblSNFFA4rXepudm1a
4zQlwlWqu7FUXgFjvqz6/UBGkRCiDDKovLs2Y4DxOFWT+fZX48on3ai/Jo4TVKS2
9J2yo+0wr0RiJ/WvxwZoNtZwBBcSQaAm05vf8Ez2jbpeZovfS9lm9rWW3va2cd6P
SFbV3BaYAVzEpSarIQc4d3qcSI1gvQvz5gMXkP4bIl5MCTus2HwUutPJxIOGEn3u
gEROVFruan7DgQOaDtioCtY7uvhyeCh5qWuNCM1bceTXso4ZZv+uqxN1eTpkgXsa
Y4/VczWVX1yyUsoAGKYPDJMa29Bweb1Hq4qTioOavTFvNc3hwEYmRTHkXBx++0hl
2AjE6NsrwO4qklOaXcNoHWl2GxNgOpHe8/AiNdNSHHP5UsRXd5Mgoi4XnJsWXSkC
aumBx5uIwhTrrrp6+ko0NB0qlqlVuyls23RBLW1bkSL3srsUl8mymP0nWwOOtglp
OppawgheFjKcqwziIl9ceqwKLY8VfuoE8gvDOVCq7NZeODIeEYVp8gvMK6y5F+wH
J/btKVnCXjz2VANZE6MHULcLUv+HbeNt4pO0V2dpmAZ05kVzaeXdYuKw7c0mFG3D
QNvBau0p6Z4uP9C9PYMT+FuZPKAGj9t8m6rvN1SvmpASG2p0Drtp7VRG+KI0z+e0
Rv3VN9fV3CNm3qCs3hDwH6UOMfTKIyqkjzf3t2Mbq+18ZAxtX0fsytx7O7ZYfYMh
TC1oNgCL4k1Wbk93NsbcMdWvCrUJLgVz4MKEUSsT660D9UzqNJSj/eJeP1+4Xcd3
0RjsbHp8K6sNdDiORg4XFN08Uo9Qn8ssbf2XJBR9xH0UeE7PtVaLEiek0UcBNSgh
HwM79ZI94IzJmYFN10nAcieTx/W+8pZimUx8j1Cv22ZgGTN9LqBWeKeN/SIEayQ1
MR3a5cW3pRtSYJsMp1bw3XeljEcTiIKeafi1Hjd5aVUDYz2qYBc6kr6Rh8cyG5ek
VL3GryTLHtPeRZGOZUoCZpK6WJOqE9FALoC1+ACdA1XIXqoGYHTy3j12HSDPjoxr
`protect END_PROTECTED
