`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaAbRoKa6dFwhu2smQ/Av2kCzc4tcWqNi9l9tGpuIUN7rNQGLFChubFCkRqGrvKT
CWs47djBYx4sghrNfZqKGnRZLkea4nC1nO0y5F4kzDuOuj9MFMac8g/PYqYycQow
ZwpjkqvF9pSC565Hal/iW2gnlhqrYhD++CcQUpJ56Tq3bOs/ZlTriovV8JpV7wHA
zPJc/zgy2hjuYCTjMs+OUtRYE/CB7ZQRaN1iFsPsKXeBRc3gi+DAfZoHU3gAw747
SWCN2Q5405QS3sJBLOj5+5Gr4Nn3QYV1jyFV7//47A8xG/tth6rhz6hWfE5AZ4jN
knoMTKI/LlUAOOiW6RdC7NXsf7JgHZmHK1yjuM0bY7KnDrzZBLXoJiCAnbBEVajF
Yp/IF+v83JtDAL54HHSLzC3bQu6y0JLlanjZaMzLrzDGGd7WipjligE9SNJJlCL6
2hEs39prxNKz/xE2dCX6LPVTU3b7t820HJPotFKuDwjmTdrHCHKl9k4tTmKhdRMh
1PW3KvHblaPYN2F3EBBcs6blaTTp0kw0LEsaVSMABqPIB4ObtYhdCwn02UDBRiXS
lbM7Bwt6UPrBC+HRYV2PfaFd+F+46B7JNko5qMoWnMzuko4X/I09aga9h3/ML8zO
GDp34eGVGNa7kDstAwqvHZju2eAVAMlxtGv8UQRiUnsKOS4Q6jibi8dOrIJJQque
Drxv/qMs5GIR+lkHqO4WVg==
`protect END_PROTECTED
