`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4egSDYoiFLFACAZ8y5wCTFAWsBC6vPidwbpwbwVuDnFJMBH9lXKaKU3jLZvqsC8M
hlI5qR22LtQ0Ul+3VVf6SSx1JNhVXZwUzBIUy6gC3+ffBRDcizDIjRvGSV9Rp7i8
1Uxm6fgPX+nYWVWHwqQuyYTpp5FFmyRkKz5I8Z9tKXaRR7L8YUx0oZvs+tjnABes
YNG+D2W5t6ERYgBY53zurbA39h+vJn+d3uleUPz7ih2chRGwPn7hdVAFFH85zK89
5OU/5YGrFpOt74OQ8U14uval4pGzzk4R+biFiEVhqNqNGDlpXClFqpBe9QaBDXbx
apS1xbNn11InCGu6hpuz6QCoy5bk2TpP9xAC4NJ9tJUwjk0RbPwZvvFYY7ABC/0m
eDAM/k3P4UCpOQINikt8rLNdfXNEzDmwD0nC/t31Pca784jr/lUMa9+r4AL6BoJj
q990fAyZGBFJsRXiXAVsJqX4gI0fUJdbzApBZ6veqD/3WohUvV0iOcvb6/L++a5C
7We98NJVplAkUcFUO8hZH1Gpj4BJ9RL87vqSp+OuWMjE2dpkAt1+PwRxCXxph4jG
Wt4eMkOOQPWMYqLTiJxa0nQ+XOL+GBRRJTaKVC2+AAUCIgz0yna/VSgvfpd5DClA
EVQpAeida8NY30oQ168xgajU4Yc5iboPghenzrFwRXgyIGQvlO+Hxz8hNgPiQo2m
33hKQ+m7kS3NPOF/CHzYpgp3HtUHI4N3rgvsGZQHzXmx1yeEOHT9Bjc/ZogW2EnG
bTobcfDrueyxNXRL/+ps7tJ1r/PRDLtwmwxK+ADf3Xy1DQWm3/U+0g9b1pAFwnYU
L0lJ8HLkEbLv4A7iHFyewEzff1O42yJHKlu1y/ILzXqhb8xnRCZvUy7z+ocK0cmi
VV1r/vSY2tBRyNV9IkpV6ajtO96acaj623U0M1UucAK1KYYbe9PNB1HDSOOxQFMe
JchEMQtoQQLfOZd7jHGympmNGN+tD4JA9149vFw5ELecl6HrIXdn5/UnD0Ytk8Il
iHfGoR0cM08AqX0ua+3NsLZBujjTv3xGU6EsrPGGLIyMux3urY5yjbw5PefWrBou
GegUVDNgW5bz+Zm1djlkP4UBYsmWXzbII9era5fOcSC6fD9fchLBCiuQqIrGQliN
TuXWrGr8x2eiCffI1xDincuF4qjMz+mS4Dat2fCWlTfDYfWpyDlLM30sL2v/6g4s
8XyzAu6pEEF5slJMA1X34PsKEF3xQOPrvGdxN04XngMDJLx0uvMss5RdoJVWjY5C
mDR7qgvZv/nh1bo4/EkhinuVN5ED5O40oSy3flTXiVZXwpTWrlyI4OCySOjHdqtQ
OdCvpXJkUya2rnHMMsVxty7byRMZ0/EFj1utOLJ38qRcuRTd/UmxRc6yFGIzVzwO
F0B5IBYW8JyE7Nz3yTANDU80w+UNwkuaqqoz1xBbOnFoUeCJT+r44Xjo+WkcFxan
O6IER6VFUukzhFiNH5ehkCwfGG12oLba78QmYVlXb40DflR1c4HCQVuLs9KixBPL
J6RyIKqglr39hwvzydE6EXaZfDLred84mPBgXix1Cv2tK89J/W+wieRg+VpdfxJ4
9DOsvElZYcpoHHGFvercPU82TOKydAm8LWtYkM6jT65EYPEeFEOZ8udrbg90bMgN
cqQtCFvBKezxpLqwDDJtczJgus9wOlmJ4V9t3SF2tCNaKHkwvkLmgwfo/ThWixpQ
h7jjOMG8ncxoi+wGrfcpjsf3aQ7W0R7p4ASAogdvkbUeZ/9CsiTrtDHpVD2axv3U
14EN8kxJ+V1GOn87+0TWsbUFhzeLJT1LuK7pJ6N2ItSvsA3E44psXbA/ntOCOvtF
ExAMXm2P/pRjY265kcLMINg2uAtkS5hAjydzhXDVQKFJSa+k6lJfjJrG0z5Utw5S
FP/ekMVMGjAdmkidpAnDdCYrY8GNFj9kvejfD2RT2iRANGvfNU74xm3IdkBBIhSk
88+gPgL6W0t2olbB4ZGCXwdIFScyiyIBkAn5RsemZfXfrZCJ1CaoDN8DqgeCR8gs
dBehFpVvggbrrLJFCcmLF/l8FT3BdP/0BWEf3YOIQ+C+2uIlvvkYkrjDmbikoGDt
RUUlX+6ickLFoMDCR4n9tN3Bca4S1uzFMR2hlCqcZAANulmDwmkFPLVbo47xJquf
fSAaeSsDFbUmyijodYRX3IJQ+LxGTtJf/A4lA7JKKVrBUM+z7+xR9Z8EDQv5cBTC
MXJch8XQNpYFPt8Z/sF/FyaSHo2wmx839Rq9KKwIQC+01/UGCPQzyljmCkDEpGu5
jCEP41pGZ+4bOoDLVIoNHGWva2IhdWziJXml6e6p4UCCESClbK0XcfeJl63fXccT
bw1sCPLwW78q/9DNt+mjKTzTw1Y3XT+jecB3YzS4T+tm4QsqEAovHEiB/tGJNo8z
5CUqqnSpKoW+jmx9U2g8CYaU98DvDacPUIbm8QeKAaIkp+AGi1b/orzHb6mwFL/f
aSLEned2F2YFlfaG+Nhk2bSwYn1vnLSefdHzlTFXR89SI0r27nqCIoa68t+TAaEe
Rcq3rs0+dcSACOZuUzWqV0noWjpBoV9xLlZPSDcQlXiDKMd/xUSt4+NIednI8LHA
A3pEkJcPZ5DMmmBQV4SZf6DlA43N+UQaYSQurvB/zFGcJEfzfazNG3/2j8FmwTSY
ir26JAcUJQ6xzipOnyRkyNvxytJs30aFGb0M3TGHQHGY7wBtouVvtf8NYCfGunef
tt0nc8eRcoxKy1mqL6FZMrzK+C6pI0yofZya01bqQ/abRBCIjSQcs9bUeiAROkya
7On5jEN+M8V+wSDHymQzWtcI1x8qeEIFLMxyt3ACZHsip6QY2ZnPSg1Zzr0mP9H5
bHuQ28LHLwFoCtm3KTW/EmWmcVXNIvnMKRBagq1/gCptjwNZaxKqKKVoTteefxxq
KH+ccsQe66ggRNyIzGeNFKnDheHhRZ+CwSdS1nHY5LZMM/knCKUVGJO3U/WujUjU
Ka9jiVLm+bCPy5pL3mJbNA21YGJ2PChD2otIQcorFLC03fcCWUtlnA09RavipG0A
5bqsIOVltftDPTKHC5bJpsN1zzWsJVYSTX9wIma0vakekUqG22N06gUXj49if7uq
jTjk9WP77xlwyyV2w2nM1TfGR5mynu3Ct9vBuc3iJmObTyqnOqS3ln9tGH3E82YL
z4MniAo2cnmD5Ng1xuAfTvUCMYhUY2/dIuXIeyJ+tqkiH92rjr2uDEov+9n0rsnE
moKP+M7f4ZFYwijh/+eyR519fBecdCo/kr8/PJ4D/UPTtryDO69V8EUDt0xujyhk
mmG/o0aGhlUxlxLSPYS4vgqkg3dRjNiDn8cQf+osK2YDL9Dr/wyeSotz52bnC8s6
`protect END_PROTECTED
