`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oWoeEXGgEo0p44cZmiccP6elsVbQWiJIO1iFVJoiwG1atttguH91hATFo7Uca7Mt
CLhcmXm5pegSdZ0pFZkp580XN3qU5GwyLow+qLKYctHuGXQ1VUaZsb+j1AtGxpOA
ZYm2qQ14l3kGuVkXFHITIW93Sug/yjWqABZD61BEf/GX3EMSRgR8lMEYlhAtxOaU
NxHc/+AssOQtF4QpN9c1cHPFsjG97WlW/CU0int2Bim0io1ot02T4EEiSs1MIGsv
5s3RlSIy8/ySbR5OC1lb5sieTceU5dfUbV3Numq1D44vs3XuPXdv4l0p9eukrxFm
gUAU+Wjek//ZGolIZS6kMO03OVAJ0QRTbMn1+GHU1R70Sr5hdnA8zU6Xd0vwKiO8
cAMY6UiPxvsYa6724N+gLByscObIYIvewyRkQ3DjgiraYOLZ+aM1RkGzivLefzV9
/W4gYO820hzR917UxnwRUB989EOcCdHriGguKJTomGTd8u2fwpETGkFzE9A/BM9E
CCKkb1Z34jgKAuoidk7vWpVBcekgsOoYUZsWbN4BoffIjtkuAwaNRG3fvx3OD5+b
MNvoiiJ5wdcYGe9Me6PLeDtz9+WW39qKmqX7gl9UtBK1P3VJE5/8UaeyreBzZklx
J5c++eNPlaex1tZgBHhmzezr6pRj9AhjVaaCWVJHOukiYHSaAH4XMka4Z6cACj7H
dg/hj3pmEMdIth2xBMbpaqO53oBW9Uni0+s+0FWTvWIW/FKtPe9KuSootPfBNmHj
ZcgvpruywLN4rziRQUcLD0G0hev4+SQyZjLbSLKJxzJLonyZfFf+vFLwEYtR2oUf
kL3NP9pJXH49Mm7Ro8MjXQ==
`protect END_PROTECTED
