`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNCZixooAe5/Gtg6lzMOsdCU1JyVNGiflzjDULrVqDupU5Fq077QaMoP9jw/6mn8
R4sxSk3m+1w7y3ha9eRrLm9iopW87qSUqAwCvYD6X36Ujubi+AGqZU56XPauDALn
xtssJaSTEdOnmhsdiaTrnOGFZMVGXkMkPTp57wuT3den55UmaY29WTKQEwpk2rfx
8wyhzGbBryeOgI/DgHCc3Ptnzya8ezGrdjqbjzxJMI3jIQhMtAUyCnd9J9mVQQiF
jZyezRwCbMv/fKT3r4RZ3nqsvSNW1UNaUyVvEnAkJQ/WAndeleCi75zovzuoX8CH
UHjH96szUxa+ORQJTHSPwiabs/XxibuWhcD5Iy4PaVxifGC8i7+pI8FyNZG8nx3/
s6fHtpXgeMWUt41qS98TQDnjYsH0dVi1XXNccT4NZPVyEgVRRLLbEis7/Ys7D+o3
UEvUycgj2nPStDyBMHghZvN5tZXTQzfarXMCQGOUkTzeM/WH/ikQK8roDeR8zLtG
FNuadukcLrR0tdHVdfOjH3F/36ZuJqnKwEf454ZT6azux00l4xlojOyon2m3Ijkg
tB90riy152Yy04BFgmRvVFcAq/LssWQlp+XKgQ62XNxsg8qtYTspH8PGkWwiaSlY
4fO3wgbHmOIRWBdhMDfjyuzUR5A1+MEDir+NQCy8xEkdOzo2DG4+z3gEJywefsej
KoBKiYVTSuLrj76rwc66lOQJucvSSoO8djEzv6qPXkmAi/hir0Gl934uRU4n9G0N
DyD+zRZTivVbjKVv+7sFXXrxiEQuMCSkPyRZLYzgZQ7/7lfgm4ExPUkFF4xniYcV
zNu5wf0Zeim8OSGrLqg3dA==
`protect END_PROTECTED
