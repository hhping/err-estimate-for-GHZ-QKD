`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FuoPpMkOwZkwodA3FdEChAxIDikDjLX1WfRezlcjsKYboaDn1d3XkP7haxmy46k
sSfdtuUHDHZsx1GZfx753eqLXPIPjoGjVr5otIXLugPngY823M+5fojnFA9NWIaw
1dwEGf9yOMruKeOSHuv5Kc+OcZzrO2qQbUBJa0MAyg5+g6fljOLBBBMGaL4Dru+D
J1uyF2fPIsxLRxAaaTHszwsC4T6VRzPpTyDMVt1o5KfVtukMa0GemfOzuLkLNRfH
Ow/Go1+2yt9uLOC9q6rou6UYvPQfkdHkz2LhRkHpXTVgWv5AB7F2D7BHNERkDNZY
kzJXJNuVCB3vsAwMB6fbcN1/9OlJ28ul8nc1ZEdB6gs2o1jXpOzOucCyh4dBZ9mp
nPSH0hh5VzclfIMP3ccVSbF7KOHWedHKtt0dexvWwPapAXkE2vd/qbwIdcIdhfZA
J55VfTiGwdFOMMLupHkLqo3CFw39N6Wk9at5wR9aShdXg+bA4UWFiFE6LvOcMxkT
`protect END_PROTECTED
