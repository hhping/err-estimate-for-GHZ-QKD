`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C7jZm0L3X0xFQ1G+Bsnd7wNHl80fticIOL1I4UfaS0HS/Owtj0GB44bF/X02oOD1
XroWGh3+/qVSLt1Wa73dvJcMAJos8Ti5y4BU41qT5ZM6IFThxDCNbAq9S4eD6IBx
+zntEK4TEddlbWVY/hiTTC+F8V2IcYOHueLsSEv4zvyFi+e91+ft7h+jUPr2/WGD
BFfMwwdJXAOdL0ZW4E3rzxG8LZMyeycn2lyJ6BIuuF7f1xdqJiIDpE08whc1RhvR
DxsBsYLq48DDUjyK8jCjYHoL5nY3zVhboOh7pd71Llu3cQlAvTzc+7AuuexgzUIj
DR1o5Uma/Vg3pDNott1TniNNjm7C6nOvGGeNH8UU7iEpWhFhej+Tlgp2k7Af9tsN
4EP+P571UpXd+JKiVaZW4p013n+zUUaXPHNnf97dFFvrmf0K7tf2dt2aeIFw0sWa
M07lQE4Qv8tEdV1z9XDrUYKg6SMa54DYKG0OVLQeHGzLLOQVGbFuxwT/k6msbFHO
ts0OtfPNrUNZVKcgbtZGlK/MwqTrXO8OyktYFIMNJHnw4ObC8llN7yzTqgDyv7de
He5ItCs+oA/t9SjQfKHWv/fqw+BWjQXgm0nK3Az1z4WL6sr7UqzFj1qaly6bjEqh
UyjGqbkTFhQ77w3kO/dSK3szduZKBBCcUk9aaZAM75/griMZPRXihm6ADFfDzTTC
oMwewl+XZ7D4KJ+2tUQ+K0T96Yqxl1kFjvqSfAXI16K4ZOZRPGphoWjenGiEVMRT
I6gtO/+dAvYcQu3xggQkH1+nYHTnJr3ZFE36ehuQ0DVIEvAZ+K72VD3DzBZsCFvu
jsCKirP5CVXPkV85vR+G1gZn1JoNDDoGeyCL6XwCt9kmAtQIAfK+VHYsf8G28PnX
JYuNTXuBAkpQG0NEVGYUrhcmhJ9K9WYgEaOhdHP+G3a8SyVGrj1liq7OEH//Q9ej
PWwNV6ncsP/+qIMiYOs4sKe77RLaREnK5MqAw25LnI8EB/ZT28aGgqaFwSWeb5kE
Lfuur2TC5cgJwU3+SvHgFaVN2ZCz+ORFM3OMV4GKKtfnDUkpxA9yp7gNBJIuMOWy
B5sNq/g9/sLDrXvnoI/S1ogcN1HxysHT3ZIW5f2HuF+F5V2+G3S22TBd+nFqjAid
WVPh6fhx/kQXGCEzQuAFD1xTOye8vuumGsOFv4mKa6Om+GVyBrncTA1dx8DUkM5V
FTdm2lTzuOpfC09e7sP5uUmpzXFrCXEnFyFJT1jozgG/x1wBePOeRiMqda1GNIlI
6HI/Ezz6VDIx3IczztViEdOsSDWtTvPfEswjGk+WAAZ0/wwAOhcZ/UGD2862MOHW
eIqlJ9jCMGRF8KEBbenNjDlopx/aarZ0haIZcUxT6LWBft0dOThl06HvUXp0ViNi
jeuoc0SHvHt28Ak8+H+5KJ4CZCCQmG5Y7Y7w3E+iUXXKOvQ/k1xIvtdz5tUh+4cu
Il1zfd3qwXdGFO092VAtXQ/1IWbQyw96RYbQ0SuI6R2IllUudhAI+uPx3sh1vs8e
zbV02QAx7xHpmyY1uvQ57LqAPZ4znPEr3zx2fiEj5PkcV2NMwT5z7XsopvvhUSpB
nK1drV0veeRxs1CIxNEH5AvdWQwgGficMT0ddPMKFSdF2/c+yObvSdpHfdb3xQQX
02JyITWoc6lpBzHotAGMLTtnas+VAWl8oOMkN1ijprO4ov5RVUPl5KOMYCPiwLY9
49B++yV6jzKTmQqhFGKcGWkUy81HtwtALSCw/ojD3Lve/cR9ecxipUkqe0pAlAdB
IgDZimLnP5oN9DPsPZ1gKYXoE48K78QapskXdP/MbFUf9SPnBz8TDlFM5ZNqeO1S
zzHVn2nFN5K0gCTwRiFjle0nTLtLG/KOz/E6o3xJEmQvAcqOIHpz8AFYsff7AF3E
naS3hSPE6Tv+0bTmqUTiNXb2gOPlEX3jQ/D7TuRm/WXCAkvW9aWqry7vuGmUG/36
hEPLsCexoEzN6mbc//7Yi5mN+KX2RSrKxa9fW1esed85kugqssi/QM5j2/ETBaeF
DtgNQVBdsdvgMd1BZERoc6eGe7bPmnzFtwWQwQvqeOTWZHQMwR3+6e+VdhFguub4
DBbsfUaNaxf1GQa00PGoYhkCeEkg33jnKP3+nAxPz1Kjyc57tyhyI8hIoWNuxMvP
lRt0foewYmTYzgEPjXm3KtQNZgKYE9jIJ+e0jrqBcmJ67GJB3yQdSGM/O64nhd0v
/GqYi7RWbUTmcfGfEXGV2lX7S+CyP8sBQA8ehty+OwA=
`protect END_PROTECTED
