`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
STr2+bDh3HT/Q+tak2CWeMsC1QgC1/aQLvxiXERqR1NtnHriofku0w+kt8ZEctlg
cTTMw3YFBnG2j1049w1sSkIlGcUjXD7fPivPUkYINFor5gSfL4fnGJb4aienGY4v
HhADIn+YOH6sznUImregDCgDdFKjHQTJsyESxbMjN1l9BWmp8kM4yS+EGYSOzn1+
FkHTqq/UyB27pcHihB/d9S5ykeznAZMk2YgWumo93Wb9TVMIQf0UDvvSuDlT0J+D
wFuy/VngV8HOGyxi2KUR+u6oKB4Y650mbBJlhFoJrtJ7Vb2JwIhj6TH4+AkOYL0D
9BR/vQT4hcPzWpaHsYKrhrK142TZHgVlJt3x7O7/NPibLoe6PT1KgX1uj09K4RHU
W1BXeQZs/Geep/SRRSFvQBY+vueXZv7ySKYKlY/QVN/6FhH37aw7gP8HrPCGgjvV
S+oCSPVk7y7bwOLMLpoZZweQlq7NpjglWj08IVlxz/vaQZCmGYKpdbpQg9ef6XBZ
tUuLtXyS0S4/8otE1STxPjMOVHa1NbYsW8BzVhUcgbgyPa1oewd7wDU2ltOqHnSe
`protect END_PROTECTED
