`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NhgzU9MJx8d/Nrv/xQQUSAUJSYpHqnuLjlQqKT7VezWRLm+hbFQN4yd1bsLrXnIx
ZYpc6VnZ6lDfyg/dKS+uIJC2n/lAAwSwigFOL2DSFN/PUaF62vKIXxZeqhvr5+zS
3nzMpjHtG+YAtbuJmVRYptUqRGI1vLQbY2Dzi41LGc8M5c+Il2A4dqNOOqmWE7d5
FqFjAHE40uOm86s4/wlyK6B9b13doO1GYgUNu9QHFgW82Prj8TgX8DCQD28UKZRM
WmHhOt4Y7wXFBDlAYDPPilsiKyc9yZemK5lmG6Y5BcC2A8CjXYJHTYBCJtS/2Sx0
rcWp3L7m8JQK7wsgUEUipJCZXQZjsBeR5muRI2a9+dnPKH6RgbKtzs4H+XiPBOCJ
NY/KupvmkDBWAl6X2muz1/pAl27pVmDYyJXLqmyceYzu6P4jpAT4qGGm/f+RNyWR
cYk+nIG2DyRMmRCc6lsEvHJycZrAnmWkyyFCjEV6TEDgVu/SpKtB17biVEpin4ad
qZ8OAD4EREpEmAVHXizdMvfUxdWU+sK8Ipo1CtWaNKZPTRPqPBVAyw2mtGsM21Ph
UZBKMIRjP2JwBPHu5y/+WX/rJpwSYNvH7zbK/nHExDJqPYCI9TsGjUEX/qFeLNC/
NxeJKRWXGPJ1gliiKJ/q9QzhEVeTa6FGXb00vQgDHQanl6/VHi/jzAClceX4Hb9n
qQUitTkmJZCl+dFy33DWxzG2PYXwU2hRYRceI8h8/Xh8/1P0+v5eowKperA3P6qO
4ypLqg72RdApfepzOndEoJu6MfDA749fClIkZ5TxpSY6ZGzH/qzr3LiNZ5e4kLP7
fef0NZeH5jFJvEor10yic6EkpwQzxxyTHbG9nW3Kxdi/OoM5Q7U9i0bIs3w7qMzC
hUQnheLLMi5pz8GAcNoFfRGvtuK0Vunon3bLYiHlarZr1HnoWJKeqsSHGmycIPj7
hbNPQSQOzXLJ5CwExGY7Vucik7WqoBcOzsaZyJhmHqGHJXxnxoSyhY1sKf9/+dFq
VfKJyknIclYjaiQHIagqxY4bUisZPGIo2H8KXCg8H1eP2PzmXImQyHcgck9FTQtm
6w+P30GeO4URSpydPKIn7q+hvPOtXIP0dva7IwYllEJORwNbHmi0a4ZraRRjZo+e
budxt5qOx2/54sxkvuo/pd/vDLW2G190C5WT7eEblWT+IPTCkU8oC+ot0ZbcTIfa
RfSD+HuW46iDwEGZbSrXySi6QRSP4MHSCgAaWd8tXvmQYb94PyphJMZp2fkeat/U
yP3DMnTcal0R9Q2mk6IeV1iUtw0XGUDtOkmsUcC68u1D4ED+lZCROTywh0WQG26O
iihVQzhEtRAqvLyJT4FV2fOMkfGTb0HjsmNsuF/MQA8g+231JKbSE0onPHXHVdZe
ZlQipmbl94xTzC+O3t+pJowwwsX5vkW7BM2FAgID/fn1Yyg1DcLBbzN1PHkW9qHt
AHUj63mz3Xnhd9jykYdjTBMn/2OY8gXvBIlT7rw7ma92xdfVh6M01oajhLA3y3fN
zok9UP1wB+sU972nAevrN0USxptV2T5M6BnR5FJRirVsZaGkAzZem+rEu6tfeXl1
WNmd9OD3poJPmtPwbhwWGLP3r2Nx224AlFFpRCyjR5x8cG4Tzg1KgK9YW8HPBST2
f7b5H6gHGQ8kghuKCL7mDcKobZNvAo05xjoeY9grN7ZwP/vULoBeuvDI5rboIDQK
3Uv2D9IXsmxtfsB9vwecNcv/+BG/Q67tZq5bDWLVUPXMbgHDsTLVme15TSdz+ahv
WI40mpmhGcqmgS9UWLqwi4e0aLG5l5YND0hq/tVk7q4FJTr4KWWEBfLz5StIlbu2
sINdqGqcw/kFL2Sr6mcSP9gLyHMrt275B52u7AlPlaQiD/t55wc6fruS85lrtoo7
yP6vlFehcxV5Tr9/6tLc9Evi0Auqcm0k5ZLIw6WYS15PhsDuopakY4X/AJjjqtAg
a+hFhBWHgOeG1VgukD6CfoA2gP3FtnSZmslqyxAle9OQwiRTdoES7bg+eYwT1aE3
WZnkaKyLShwCS126YcAS+wYC3A6oURNA0wqgz74QhdHRGvNZ7gIEnvMxBiAtrzQ4
Jl1uWV6xSPCAUDr4HLd1NYxOVpEjO7hxY5SgQ53iaMwqK17yXw2ecD5+1is01Tho
qwaOZxcHdOap0t14D+/To7WCY51pHZI45qCSvfYGqN2xHIDwGxEe+rFwbu6xrbkm
m8CFE8WwH9tI5TYDFbN/ZDcTcVhVifnZ9aAvO5uaZhYvRcEciSFI9KZsKXa0RJha
nOl57j/Yu34vUfG8lhcA3RttyVEz1nCM/lQwy+H4p05inDaEyHwd3QoFunzMyMsF
PYdKY+L2ZenL8AWtpDcrPKFthDx5PUNLQQQeH6cGg3Bw6hu6RPwYeKDe0t90ezM4
YJTrh54ych1geAoLvCQc1F1S6RZFuI7rC3vzvoxOblljWRQo3V1vnZXryZ29wSIn
pjvSuOI9vDb5MfPQdcFpHl2xk5CQ6PZOj1y1aOq116t6RAJiioSVs1siqN957NNb
GTF7zvWKO5Cv0RN5hwDvFlf1lgd3bGr7DqEV6V8zzIGlC16+COJDqo6amqBy1lua
XVTfJ3LsHzAGUfJX51ir8F0aYV3gR1BuFKmpGKJMIXOxSTFHQTEnwNxHuO0wKubC
/thFwJqzHJ2SAiev/EHaRvd+/tF3pOX7AQHOWYsUnH+XStD2h10J4L8voqL0I5kK
O57l8x+jp+MpahgKACzZUooEpnzGWpeiHeF0wtcdSE0EOv1uUCFlXDg9wPEnh8Bb
YISME9Xoi7HbyNNMZr1J1OOs3dOw3ZYP4Gau0J9ki3UGOgZGl/1ev26Ui2ENR6QP
VoHQ4Eh+pGEVpcR2jNG/IA0tmGa2VYJm+q6bEk02msc11jJqDeKXExvhnn22Db7c
dVIrUYU5pQboRdUs9vt/w6z/L9WWa1hHA4nb8+AXtpYLVlDtleemlvvTFZijjSck
CT2nViH/DFQAvQThyEk46/AB0XeSgo8kwgoB5O+dHrenT3OGFaa+Wqnu7EfIHTwW
otbDqvssHq8K+nvCCh9CcOmXzN10dT/3VQrPubA0FZl6WPqi/XOKj2zlXawZwdma
sNCH9Ev6joHHWI1U3jXFj5y0YViq7IRcw7YKzc9uJmUD80O5ROREEetFEMu1vGTA
MokA27HS4j09eLcrO0MkwsVPnQDJefMONhrrX/CMtoYE/Nzi4hdXz9xgIwxus5cV
V8UMDY3txCn11lRRmrl7fu+vOGerq1ZzgpYPp4fiUF0D2u4pBgs4hlsGalMPeHdO
wVKzW/r7OlYsRW2OPgWhOepXv4dQroB1+OCX1n8uNw52PoHmc2TOf3TZ/DNYj3rE
dnECt/Li0TKUXLrt/LUInZOwcvUagxeHx7Rxh4uTpQPtEu4S62BW0awxj8Kev9TI
Ab0Woh0lMAfl9Aj3AYr1Ac0WY2Cug/6WmQX2VQnQEdSNjx75fmFdq0NR2pC5vNsu
CKeyelMeNakZeUYA5HprifaBFl2lQ7XY+ZRyKqX9J25/imfhTn6ME/MUInlvZPnp
5BZ8SiWFWreA5hlLUbEzS7Etg9AqX5f4K9CneBr0J91rj05kgdr8ZH52OIJCywy4
kWK303X5mNfCIHmnaGsmKI88JdTin0sS4+b5VmMGx4o8WvwVfDPWOz7tm2RdKs+B
GyYs8UzvYMP4UsYpsnhoYAaW+GSoAt7sqcIt1NWu4qYwjWDTuOq+LAswh3A/COjt
w3m/y16qVrSjwAkAhnPbPQfJ//bHszPARPMkYeQ6hwHknr5e6+Dc4hkq1wzc8aLQ
K/Ci4FcfWCHEH3/fstcUr1YUW5MUTk+HelI4JG8GoONgS7GiKKZk6ugvD5TnZEja
gsPRQrgPDf9Ktuk85MTT+FixaYUxVbAiV0mToESaBdsKA9oZ1e1zH99EZUQNyV5h
h8hJHoRjh3Dnx8CcBmh6Ef99GiUYRYgkkHptWezK07HZ82ElB2xwrZ2DDuNgcXtg
lpD/eaAa9tMmNuajhh5+DNv5V6JgGfej8O54Ne3X1JvMZJF3AGx6pp5CjglYf4qz
ipjBIXwkpYHPpCTeBcgbkpNHqbQtMsWTbjqWCvUht2JgfiX+C6GFkqvgurEq8MC6
FtWSTzOjZIhHjC+wApaK9bAowI434pQsV5BJNnp0/n1iyyHgB8vi/kMWkscsJdCh
ctJL63iTf2LLkb1Q5GLRGSWH6iC1/nUcmVm7yH7BoeMgwoeEa1hE71nDcxDWTAN6
SY3B08ZsRp/L7EWDmrBGD6+1OXsyS1UmgtS4/672dldYmeC7ouE0W91LakcT5gI1
Sg3sFXJvuSSFJtqf2hbm4Xqs7cvvftOH2G5vkPtiSzepwltJ80gT7B8MsOn6PjfT
QDtK1xuzM79Ta0yxhwaRFNrcuJc3T9otBKZ//sADBf/Fm8M8tMqgyabIVAp5K6l1
`protect END_PROTECTED
