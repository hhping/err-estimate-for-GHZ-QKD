`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kAcpwxsbYTU01rtuhZBbMWUi/iUNuE4HQc++GdYEYdkCiytjaeHJrJjBYqm8teg
Mg+X8Q1nusPuig/yxTf/knnBe9uUyhJ+6dnUrlpM7/mJaL+V0R7NStOxAhpVgm4w
2nYk2m7xrz4WBrsO/vh2NYXlCVkxl/ikqi4G0DcECtNrBMm2UvTDbC/MK4t0SsGZ
fnLd5jhXRND1oQpgHTUpKPbVrcHs7g3AZomeRrCwY1jpd+4NVSrbRsXnlhNKRmWu
BxFz1k8gVcaybIa+L2+cr+XkL+aFl88TWO5wP87WwRGv74p8Xl1lhg6pt0LXblAw
Yipfu17x0phLS9qQik4FXkUIl+Z5THAFK3/SXwUBvQPGKAiTUGtzBGWBr4utvhjY
u7/H4yIcqZEQe0Sq824r/YLFqanBAL2vrayCvRJ606RLyx7QYpnYhNLQ+3v33nuq
mGZACYWEgLgCIgNJNjcG3miUqRsN5avv3JUQ2MNW5qAquwjLMOpxfpJExpJcdT3a
6XheohRKtpzC8Zd0OI31Dzxxn+H/g6Kl0JzD1j4HbD515i8kUv1rVGAZl4dMtF3U
nR59ZQi4uyj5aDV0HldD2hHa19b92jJMrTueMrzWdd6DymvEhio3ExLLXJu62UZ9
pDWL5pcJ/XZTU8foYQ158dqB5S0pP/VwKxSEVC7ZF/jL2NJUaN7gxw/DWnMCqQOg
K+tzbfDlzbHKQoRZQwkBUw==
`protect END_PROTECTED
