`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PtQLIgQKrkUmOL7wq8MvBO+JqqE4az1Yn9y/uZkWtc+RWb5rZWCx6TGmXuSI4Cfu
UBwUj6zFwCgagTDNBBTjACDCY4I/MXNdGOk4/ziTEd+YK9I3EkNSqIBeYNpGw080
rldoGTXp/fgrfUkI25I0m5ECstJHx/NpR9MheFnikcq7+FRmIi75PQ2woaiku9pO
a8nI4J72YfNlZZaIaOcIjNivqO5qKr7zv3a48/kfTdCP93CpMdFj8kzuApaRIqxu
oyhlx9Te76L1pgpWMQBXC5DsgaC1adinFC3HWsdHe3r+0yrAvRJZi3DSfXnrsJJK
PgtoCkh/W0lqPfJuqQnY8n3uXHN+82bns4+kKUmaOFmXDdFa5ut8GxAicLGR8eqN
kFO0txec8QFKWC4iLyX5yu/QdLDF3K5yx1EY41weLou+Qdfk17CW7op3VB71hWYw
g7pTNgcWdE2qSngGQQET8sd1jKNVW1cOghWP4YyryIi+dwCe2VpQMssWdpYFSdEJ
VJSPCBaQ2mHxvyH+y/Nw7QatPJx85JPxPPUVLowo5kLY13+8Ig5l3Wc0g+fLHoJJ
P0gnhXc48mIQpqlh2xxfUZCwoSkZtPYeybDFLbpo6irwweAKJwVJgTfGFVDXWDAq
mien+7oKhQ4S5olDeLLxmOSbi/nKhWxGlSDZKKOgkf0jt5T1NwvkQtSGxX8I15Hm
eoyzIyzSmKFkpDsapRp3sJVbnlHCyyQe2aKvBfyp+2Y=
`protect END_PROTECTED
