`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPvwoSQPHs0Qq6fguc+WNdWzX7Ui+Sp0HyX7yoSsAN2hMWpvcStgcIPRnutfIx83
0DJ0jtYiFD51YXDDDPuuhZKK/Cw23MEjArWsWM3s1Wm/Lu7oF1Da3ECme8d96/Vo
jUcvGle9DWjZfzyrksNoY6bswl6O4ny7CSrPTxEKhkhBdmVHCbRh0rLrth4VMXoX
Zo530Lda6eESrsancIEDZnXTNthBTNYbXcCLFgXAA0Q9rAAKcxnSdHnIYjpoobqU
CihwCoYSjBN2Os/8/2b3tPfW4xab0l88xpZu6uY+urvAjOMMZ9X5JwjrhvxRWsQ/
JX3kv6v8w5kC9A0YL5uW2cQfj4xVvaTzQWfpmO6JrxTeH+a50PRuGNJtw/prSQK1
zv6oEmtmISUUcI95RL8IbN1wwrMgVB3dwdIwK3rTbEJIxxaVPjgJel1ddIP2016n
7EEaweFLangOxdujn+zl1BXGh/eNq2/cmR7rMU+66zXi4IVrWrsv+p+N56QGVNfK
ZPafoHqRyl4F+EmmZrxsFzrZMXPDS8M/7f3BY8lSvculUeMVSUp3yJBkdoP44Opr
jQWbPL3beK4DC0G/g49iWqH9/SRu910qnRtT2SXfO/OcjQjQWZ4aMw65uikK5Paa
odZAz3l3dW5GAGX1D1cBlkAmLIH9nke1X4tZ82fzfhTgzO8jX05COo3Uzajv4lij
WfoS2CaLSd0q2Y7V3boPmH4iIUHTmLHQ/RRBiI0qpRzW5ViSInoDMKnvMTSmEn5U
LNJ+q6IhhphpHi3fbJk1xPfEpJoIPqGC9sNjGu1d12Q=
`protect END_PROTECTED
