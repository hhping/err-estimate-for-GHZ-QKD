`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FqZwNy39v37G7xrTHijq96Tk08xQpJ7tMUpOaaj4xuw3zAdqEkUEDO5e/+0y19qg
22O7JzYHWZi3/mz5KL0JDQlb/3B+mtyTpvCU51Npo1bwN5divZt3/2SZaCefdcDR
+lcLCKDu93/ei8saZOoaMHplbSuns7OSQPeadPbfGDehjz64faglMX1TyGqrtGHH
/8ab7P+rKi6aBYXsgDHMo3abpVvtEh2h9oC/AE2qxRx4U7sqFcIiyiM4q1WMYVIQ
gAzd5TOHSnTvanPRqUW6CzGJhOrsWHgXwE7A73Yk7+/tcgZvJBgQQiLNbaDsH+qV
tJ30MpzIOc69aBFbMmsv68V+QIQlvamFahmm/EGtKw9EKe1CUZGsd+xJQ8iq/sCK
`protect END_PROTECTED
