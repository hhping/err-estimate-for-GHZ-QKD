`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+i7nNph3IXgWFFpteZIsO5UtYX2e2wC7dUT4hyGXOyOEgt2M0A+tx1S3aJnNdSDD
+fJv+zpG6trfhjFIu7bvr9cq/Uh7KTmpa3QAlebUWXfWfUE1OFrz7+Qte820EZ8t
H9h25h0Axnfr4rEk6vFoisIvSZEb0Jepp/xmpqGAO/JNWFZNhyfJZNpBLwIwnZJP
d6ovwdCcUbeFZbwQv6p0wucPnGqd9E+CRVNT2xp1nSOeddfFzSVwUpaHGNa27eIM
H1CR9nWi7RADR+mh2D7kS20EM6h3rQB8DEx+/FWzlmQrS68nKEoTF3JG20hzotl+
K55cv6ZmQqRweUbc2l3Ar13pCrL26FITMxSljCiW9UokDp7ijPxbpNodD5ArHPt+
KE71AbAu3TGRrgk5vKstlzSS6sQG8XLgotrvaeYTXdVV9b4na+0Lm4Ybq1Y9O7Lf
tmGyH22uzSPdOYIFNv51xlO0VsDwgz1dav+v30HB6iI9dlWpTW2bWpLWyGCr2L5Z
D4mhcGvhKO/upvGMTApXs+BQzr3i+I45h+WZHH/nz2BwXjTW3kp4TzMnkOaYjInt
UEb6LmykcTmkFIjLh2+hl58WkJ2gAmrN/XKH/97h6dGu0/klsluDiICe6EDjGgLn
C7PGsHySmPk0ZRn3thb7QcJc6NlV0ggVOkil94gNl8wvbYVpVOjBivcqKSEBbGlD
IRXiuLV+MzQTP//+dCQZJb5kLM1QxNrrQaYVztYKyjltoQHT3iZ030XPfyBRZcrJ
sVXz2aFyAerDvCAF7vgiQhWAYZRVXmgAWe+YbjVPeK1JPY8c9D2Ro+rcMxSe7vhB
B39o0LfpCjVHIHXpt239bS3W5rhsLVYM1FgfmaXannxpZkZyQ6yOKuIj0nuMTQHw
LLPjsLBxenL+Vu/wYs4CIypUTwTNRiITfz8IavG3Da4=
`protect END_PROTECTED
