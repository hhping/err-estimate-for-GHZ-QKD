`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+TG9gatbPCo+AWVrlefwYH9LQNTg+GAx0HGNNidK519V7JlMW1h0VkfdW0OY+PC2
VZQg1cAwGoajipexU8yvyHrenLQ3gV50ghtOfo6zm69u9nump6rsN3xkwIvFahRT
Wng64aHgIJ+CX3NktsDQ/5oYeWlXpSDe0QZF+P/6GIIpFH4vavRS/lXK1HByRSSX
TrSgn+p5dsH0iFdgCUi+T+M+v97auzM3f4t6O1Uu/ldsM9xIZlSt5GIOs4NH/7bq
Oun15MgoHvaLjU5pC0eUP7IfrtkqNPfDcY/3lv+Z7OvETJglCQuTuIkQDsNJ/RUG
p3840ai6lTjStlheEwDuyd26r/heJQHOAjTQXCtnGpy+LThKTgUX8Gfu/oF0Qrg6
nwx5Pjyo/sampM32ORCXq3q83jqn25UMcscnJZi7/SYvTcZeBIpvw0xCil9iH9qt
wLs/draeSd3cp0CeMRs+PVQ/izE3V5IOJeVrJMqdIhbP3PQDH2o4vBrytCo9h0rB
ftdLc9cMg8M1+ZLxOIBElrDyc8UuNvVhaxffqNBY1TjVVpszzc6kk3xNp8YAoONe
3APkS6sGpA+quVZX8tbwb6mLKNqNqpIBGtZLftqJNuHn22Wxj0ymQ+Ulm3NnWVP7
AACFxEzXaiVkebNJK5JGxZKKkftlS1byjpuCElnw6CJlwwGoApxEOCGzuZ7PWUfl
eQ44p2+hW6lmfUmyly9P86Xxm1XUDUHKiIDWBlmjt7VqhhxS+qanQuXhn9hsuZtc
Jdco4B/GpHjQZMwNyoNe5gtec042cTw6os1Jnvl1yGRaeSYws+W+2StmzDTLmJ5x
1rgE+by523xQD2rLh4oRVCVfklv7Uzf8yU+/X5q1uqbSSvz13M6Lhf8kg/HoPh2h
6BHyWagLFkS+5H+j/XYiKA6yr7ld5Zj1RQJWWkNSQX8t6BLmI9S+k0rVpnFmSOv0
1uzLYfQ8TXLRjd8dVojFTLOWQcGM5YgMKkAIPIyjcBc7A87wu98U7B3UGsZszxYO
nU/smVE4P64NIlUFvmkZpWfRa13EYZx8fpI4m8jSbIPhXDx6lL+NcliJZYkOVqHD
ElkIhBmMlm0+cfVB0YV49HnSJdhs7YtqeAheiDwpMbOgGJnL62O+VC5hcMJ+lmk8
+OY8csumG1MdC8qHX2quJLZPT2tEAka9+X65aJ2ttHrC5+WI7oy3/hqcJLKppyei
OtVxEW0NCvJ9zSMmL55mSkhmp4n1ShJdBT/NITUTYqXcVWJbKyIH0BhzqA5A3P0J
VZszggmcBMHjz2A9iIcbMl3VzkYtFxXZX+TeWiL/uEZ81V4yZV09PZWTQjMYe2Hk
CI6a3A2zkH9CIeN6No6zVlT5Zk56oP348NnpTbsUWXdFUUDlH/5cRUKAMek4O0i/
S5EFZl4iZKzrVUUduMzazLJR8gU8411HgaMb5NaBWcF+7CpwpWut6iMxRI9rlwCR
sQL/eF3l1ceEJRA/EIFWMIczzUH+N1A2yUv6h/gyCWRUHRlG4zrBE0pzNKpQbMUK
LZt6/OwUXO4OU4NTdUj6UVZfAqpeIw8CBxctP8GHWofguw1VxbzNvhwOXjL5xfR5
aYGwbrCYbF6zOq7k/+ryNrJgb6t6q2nN71Jw716MWveR01maqsckJJrM/kLxHpn7
OKAvGB3CXi2BPD6xAoE+D88i4sCsget501wl9cZisleTnjItDfDEMEefJQP3YF3F
lhAg8aN2ezmwHA66cUdbKoAIFtToRpyo6Gpi8mByeGJ7mIiVKpEevfwsw2+x8XQi
8MU3M0ycUdDhC/+TFitivE0Pd3AF/URCYArDc6kht9bpqsJq13772B43p/Ab1ApE
DCHS0GHqmECqyeyia65dMdBijEVGS0dmnemSkel4RIQO2uFFWOVq6vhxOvGEz+Mz
PPQuBvyMAacjkag9oYXn4UcmvHtyxElEbeejuEEo5uiCCKQ+xReDDw3gfNFtpQBB
Xct5gxfXCUh+9unUr2Z4640M7LD2jULHMvo2JbHzk5r7nRCY3x67oRb1gpJ5qzcv
1VoonrmxrF6q5bm9soZbocJ2p1pCgg5cQP+nqsPBz4KVbvWD08ElMJxrnu5fJmKB
Zcv+2VgOZNwr/CkOm2GqI8HZRtiN4uT8LUnKQo6FZH0T1YJrDyCXY67kMj8GzXTj
HLEXWiHKyMLhkvlLC35RA9WCjaorhuDTNnf5P47gE3mc5p/T9xWIzk5P7muBVJwK
t/lCRGZgisMohmex8pV7780bfPjcfOprnl/ajAjJUGVS/RaUa9XjXf2JVMOeze9y
aX0xGdShF4N6KlXQCeQSvN37bsWdctWljVlHpgfGpXDX42YJJuBN+qQ71p63Z2hj
Ucfx2jJoENzeT0LSZVm2+A/lWjoUYn6ByjcwGgW/GTARCttrK9Th48HeB7M/hq2h
1TPxMsZKEvvqkMxI+m65XtDyx4at/GoU6d18/tjvtWVP6L39jLFh39udgEcKD+H3
/p3NvTPIL/0EWQn/H+fBgAwmBwZM18T+2ZlzDnERmjOJMohVX4JVvR2EZStWGWyF
UR7rtmsSRUCeQy0J5NtfT1F3dzj1XxsI9aZBqjeCMQEft1L4iZ3eWwkppGfqA3oN
TpBKB5SaaIzxp9Yeh2rh4qibTPg9YDHF+WKwRPah2ign8Bj8fuWXXNNjnda7voa9
kcVDOdJ78AYsomLFaUrTxaMMSQj8RhOK9UqmQ2CFItVKb7btl8OiPju8hOYI4+t4
HsUlPokZRLM+Y+YgikyB1NKo6vUHVprfutdDR72ls+mLbKviRLUXBOFogVlvMTD4
2738y8/Xe7ymHt/B0rQ5iX5Vhjk2WdZT3hFVBb6VUQHFcNT5MY357U7jh8WdbbD8
gqsARMU9UTI+X56Izyac98+HCLhRGQuw+scnIjsq1c4/qEN9rHsrM8LSH1WrvGnC
WtGOi36Bqh1UxU260k9EkRJO39ikm0JQxs75BLLXeTYbKiMMa8OiZN35qhcrOd6h
`protect END_PROTECTED
