`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LS8eRq2FoLYPDIwxSSeBiNWWW/ajPnV+awnMHDPkIn9E/d+4iC0Tgo31n4akM06a
O84q1iP099PiLbWqw6yUS0nWNtTLReE8nuI3KuoPSMnZUDWqyc5fi2i8r4QFaEdP
za9TYFUw4Llvwdq5IpVhWJi7NLixyorM7b7zG/O6kwT3VuksiQnrcO1f3X5RLQuz
KtpNw003XXRvLeoJXeJDfMLwv/fAdwX/O1WFTrWN8Y2TIMMVtINoMFueCsPmkHUy
vabm27bFNQ3oDTj1w/AGK+4dGw+jn+kO3HBOFIAhMGtePqF+maBSNM5i41SBChkI
8BZzad5J7eWlnsYaN4qOxLmmC2Lo/ApaXf/Iqt9csYWQC1NkDR7jq1mPf7L9+wqP
GPYWnLZ3eMVeo3iVh2CDI7+M16tJ/L/VaS/ScKtHUAXP9OkWocWgOtTIz6FoDjpp
TO7yohYXKg6GzFfMDb367qF+eLdRhLQp6DV74Jon4bt4JkhtwAzA67bbbz2EsVG5
QyMuBAiFwRD89ue9u/WNERq0VcckyaMViDACX5Ya5WHwGbLtDH09Am8FQmdnnDlC
Qg/CLaum5iKYo6Awp+TWey0TMw9f7aPZ3JGOcFBf8OdNs6aMjT+xs8L7Z59jN4Md
z3nsccAwtHvdYhFcSV4RC1fMf5bzQ9+SG0S0gk8GlQ6H1V64ArETtRwXtyNmI/7p
RFGkVkxVpvZ+1heGUcojZm37FYLv1xYw7IH4XrQx+mjtjQisBCn4ToJAYull/Suz
PnkkYGu2XKrSb5symuDdTsLdlBH/IApBRAfYSgfORQbDrbhcYWct3858GcuhE9vf
Kqfsq7A/4KlocU0vh6VHcArvj2p6dRvEAnRE7GWF8UL2bNU4UvyyIsB56rH+wRL8
jR289LLY4wJH8tV0sQOOybZ0TYs86DuK0ZhAwkWUI9KdgCjp8o8BsAu5TXnrU/WD
imOC0VioLQ/Jx7bRFmB6ob3A8dRcYF9HakUnr46bNktclUiZFi3KS5Ttp8ncNFrL
YzR6qU/whePwJIBXD5TQf6V2qAfqGhK+BQnfJLFhoDe6xca3CbEnMViLPv0uqMQv
G8yS+ddTL/k9lrtLJkatZjRA1dP1NMPan0bfXM7H7CDOhQ74I58/PM4J23Em0oZp
DZZsNxsmAH4nDiMlAjnrkxta1uCtL+eT/z7f9lNvIYs+KL+VQAZRq0sJauw0nFRs
uRuszpYSjVENfkWi/drFDYohyYlXxFrJyOpvKXc576wYAkTYrZ7rfopDHIL9bIqZ
qcYZcC1w7B+t3sVNMu384W2RDUwtXBfninaXks6+J1D6BnPeWBhaYZtRheRY+JQJ
nojb4Hayb5E1rY2fNH7iUvTyPj0a2Yh16XCm/Lc1QCkEJQN623+3vdJxP/jrYdLp
Bxx5Wm9xxSP16N3VyVOMiZJl1VRra4+5QhJQ7BM4jt8k1Wdc30cOcGeWagm84Cit
8096ekzKVUuzX0cbYB0ou8l+zvrPApvHb2NRPt7JlS0=
`protect END_PROTECTED
