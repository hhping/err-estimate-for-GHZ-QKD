`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZ/48aRytM9oGVc8LEUVqPyynKy+TwqD0Gi+OorQsZ44FFAHWQmS0w6v6LTF7SLn
zKLXvU/IqNYAPsuuNU/ozKHHvYncuFwQrdFvkJaLleKV+VT0F5EAhmRU4fNLmfmC
vau6JkhWlICWQ9Bev2Ygo/xBh4RHrYNu1067DlN+bHlDo2xhRnBc3bWuK8dgVW8b
gC/RerbD1mXILVkffMNDITx2khccczpHrxU9OSWndpbt5t9uFfKFZc7t+j/e64H2
buUTZtQtOA/RciPQBj7vuhCRzYqru/SO5TBt5uuFBWamBAyQaAxgjP+blqRGhDsM
erunWmAnugq6IOIuiR4r88X33NuJTAZx6FoKJzHGLCUl8clTPiPhCN/LKe6mD+fh
RD1VRRsL6P4Yv9kUApIrbh4aKu6s2ycsnXAXh61WO5Fv2hojveFTp9HV5Ak4hO6u
yZUXogjaaRUqq4rnDSqGFidZ9i1FkfKC7MhW78WZI1En2EhSc/uLZThsbfaM/EAu
ieSrPWEfJQIwL6Bj9ZK7eGvMmYpcQKK8A9/TQEJOJxgQ9cgTogdWRUQ+vQxpYZM4
wm1aHTU9vN5kUFHyYUP2SW9qhYetZ0B+mkfh9VSrLRaYrDStqpX0F5TEBIYS9CPT
JDkIArij8zo9bdr8O8YDfwQeC4LRIscx//0AOBgQL/0p+AjW9W+0i8g7PMOwNxVr
eGAoJtQIHKRLfjzZwVOiyXzdxQd5kRrCTPg+2E50ksxtkAzjj4suLNQ6SgxiaL80
DCWWkviCgeiMFMvN0fooCz8GE3iG4fOkvwfKToXN/fB8VzEl8mFs8fD7nKce723n
9kC+LWz6zS7q/vCLeQji8JzlaVF4y6Aqcka+pu1ZONpdl0LJ8qWXqWUDLL0S9lvh
IJiJsoAGQAxJDNgxCMAbOmWSTRB/043QGrh/V98Snz1sDrvWbDhd62c/+x3Y5LNU
Zp5UZE+4a34aS8ogLEbxfCfunlDCaEaA/lUUP1rtz0x9/YHySS5VcmSic2ifzFaK
Re3khG/7iyBPg2jq3vrtL+7tyKjZFkFucJLW9iNLcfiXr863tcRYUYJN/wcG7GqJ
4rzN8LnXQ/i2G57MAFLhYoTEp7mEglkpw/3mk7vRk5TUXb1IQL+KzTpdqRsbs2cE
ZCHJ7Pbbd64fLnAOCPXIrRIIuDH/DfTAeFusSa5/tGkFyZxN4MN+zTC8dyZztG2I
//iI+VldpDRWmihFfA2jPG5+3Mjwe7fEW+bSquK3xOVwDVdDPGi/u971wQAeJ+0t
Zk3z0AAbr07kfDtWl/dMXQcm18r08W1ewP3WL6RCUdtu8Mzlut0pOGqITTtMVNVV
`protect END_PROTECTED
