`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYr/Cj2u3ldyOBnJZutEeV/fAoJifr8TAxEHEXL0gkIdq6gG6Ld6oHRwGX8rM3UD
T6v/RlErFIm/q+NROOL9YasoTqPxWLepkAor3Mu8AxAlXinI2FI197nKFU2Nf4wW
mTPSM2oG1AWmyxHnYrh95YbqmyHfWDRTIZdl6t/+jcnXH+rCZJwwzarxCuXhtqkQ
OLlLx7m3qAC9zU2wmNjSZONIxduuW3v9ZeOJbjHJOenDl5Flhg0EGklEkdGLblZ9
ruWtVXUZfVh7OUOu3ssFbEe2gpompuUB4Dj/zu3m9MSg3Djrul1a+Wrx1VKAhuzF
QTXQ3fXsIcEyUXVH27No2XNwLwv0OiuaWUF905vqRjEqEvY4aUeFYCyq7Hg0Zd0L
bvsimeuyOw2u/RCkh7A5CmuaoRn4fMRBT5YKWoo6uxxWagCGE1fFuz9lByUu+oX9
24OrEsJ4DbEzWOxKnwTpZINLIWyXEGQwB08L737dzhXBLW2++zqB+jLozJ3qwsnn
/+SBUBEdSorsManknxrB+GgdMDwbi+KYmzfNmVBH+BR1vDjYxdLdAi0FBrvy+H+d
GEVR3EYX7PdEc/JxYbqeYc+VC4tO/HpRodXKcPJcE9/yy9lxCI6bO8YJm2B0p7Hg
Nd4livBPtnnICTDRJjpHICY2aqW74JCMN9n//Kz4FH6QdMwwLmmjUN9QajDgAu+5
90x8Dz08jl+NLXMsu2OhPrULqYlmNNJi+1ADQCklH5Ucepk1ztw4rXpeJvSab8hz
b4E/ha99/qF36/QgIXShGxDxsemi9Gv1I2nvKMPEYDVXzVfxiICluts9+DMCAjup
7jnmi9tfYlgeYMNfHC1Rf380ZlUb4m1ZnnZ9Pl/wm0dXelgG5m/b4Q0JYYU8OjgS
LULcoF2YG2hOmjEhm/2xrKghR/3VVbG8ymTyLWQbTHo1JjF/zMRW+/vA0GNhQZIF
HoycBV52lWbRxlFvl8j9Cz0JZvlXkomVluPNv/uuOOpqlo3MqLWvs5fuVCcVtuKF
pUtdhGgrETJq1GOYnNviryb7ni+SMSzalPsplCzeIt5/ZOhaps5C3iYK0a94Veq8
SmRQIgphdaRf/OJ00Tw5NIt1CApql/oOnSaP6Y9AvQfUpp7dw5WU9+InG2Od3N7G
u6Cmbp4A06n5MPwviYQ2PX8t+abVaN4zaTDTGXRfDUMieHhOTZiRugHi2GBRRWt7
QYptoajpTwdmEjB1/1xP5dyduf/Ue6ONKsWSAYqb6W/DXPuJq45kD2izDMq76YIF
FNYCr5z0f709x23w1fyWnNfwZLkUNkBz4WX8KZC+aVDwlxU5vufamWSZ2+wI7NkW
NZ3SEQ8j53nys5kzUd4rchFO5Ih7OlrlrHU4zw8kj5LMnyjeQhZv40k7ZEetULOo
Y/pcSn8BiSFNkGs5hOo0mufl70U7k8+yvgVIHBHqh+lm3CrYHCb7L8Cmgk/Lx9Kz
/rHf6B8HUqV/Bf50T4aIxMlOVDDCHGDtP3qG33oZhKyJ0GVYjjhZl8v1nqpRZFKw
GerabKklwMi9Gnz5OLEQAUBryd8RSqgf1P6NIyzNFB3kjzXopAfg8yb9WOTvSTq8
hhML9zGADZlMcntTqQLH3ZJxgtGI5wBLBIn45nMbFYI=
`protect END_PROTECTED
