`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/vA/XVEz4Hw2pO6vy9vy9bmPeM6I4Gf7fIXAoB1Yb8THBbwxD7+y8CZ/sOJXePM
JG45mRHpjbSsFgEVSN7XI/Y4/g/RMT8jt8ddhV5J2lra/Z9YCTnxqe7RneP4SR7h
yWPQU02S3Zcafu7psgqk3oG4uPCvYh35kCJqcrTrV4KrXmT8fj9l7U1k8hRJEPob
Mif+QptJ51AIKtwEoXyLaM1e/dpl4qN3bA2r7UwhLamdBzFLArPBVUW/yq4lov/A
ctom/b/Txh1F+zK/4CE28chPCqDPCAAi1Y7jda1FK14RCoTlzHMBM18Chipb6OlP
q5dTHOAGopMuAwtPTV3O2hzBihqw808fT4/y1U0BFJekHY1RNuvOVGoRKA3VMyJm
`protect END_PROTECTED
