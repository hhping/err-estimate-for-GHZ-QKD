`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yvu5XUWGBVRFyNnWZajW1DUoMPqgnvj07D7ofPxFNCvh23ppe2UOrGojD//Hb/Bi
Cj9lNVetRhpCWNMJ2WOAx0Ngn3YmzI741Bebd8u+O+CvRiOOOSYuL3xvZKx7YoLH
/BbWFZTRmERfj6eAC82fYoOB2xZIu8UyTBPjMjRtB/SD0i/amntUJZlr9ahX2kq+
ASbuUQtLQjqv3acLwbSTTu+duyyCg/b6DB83+RM8Ve953/bkVbVE4SplBmtdtDUX
97fOrHoBZccY9Kc4uyTcxpVhkRUbgveJSa3PNy9TTOALU9LZiOqEqsS7EiGgb+qP
3TQ5xWo6Pe6S0M8sw+0F1gvOOzI55Fe6D5wiTF8VRjmvQ1+T69fmgQolL3HNk7g+
cHS3IAa6Cxl5g5FmKzEt0vE1otruQOZWT70Joag3yMYoPVzWT1rXbba7DBgraRHO
g19OcgqQsXo+Bxmbg6Y36EburvYBu39ObdCeJd9noU8IlrnusPY8ZhjvS6OIb75r
uJoec7Fhm2Hk7y4yNInypxDnatziGku+qKbdkMYXK2lIbz8Ew+xWNKNHWNXB0Yvl
MysF9CDT2H3r9MkgTGD4ShJWKND8obA4RNemGM54thEvMTVgoXjNEbSLSep6nwqH
Nh2taTBiHFdfLFltA4HCslSgVzYAZ5hQohYU4LxOBG6tJ5DO9kU4hTEQxm/OsbUO
NzvZbwATGXOypSL3A/NM+KQsAz567yyH/pnh2hi/wRggAt8Mfsqz6dEyVk3R3vLg
wpNGehLulPtngNFkrQliwhNh3MEa30ehD7NWkLWochNt8e5U8jukM3Jmpk1yliLJ
BTKD325ovuKhpm2csAiJzQ8XQXXZYEUfQlhNCRKIqfvAs/ZW8lz9E3mCeYgwr/I4
jPXY4g460xU72/BQmgiHI59MRU4E8YQEBZUKjQa2YslQTwo+qUZOrK51pwu67eOA
aIWHYeWvN/RDuKFhbwWlZMXi3GpBZSY0uGt8KaFFQ1CXdPTSfwjdcicExrS4AJHm
A87i9hrsKCIUwaxGPZ9RQ31LkO2UmUhlAit62Qu1zu1wG7fX7q28S3DqzpvJs98e
`protect END_PROTECTED
