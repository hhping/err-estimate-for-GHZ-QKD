`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqcHph41mSgr4U66SbcQqeRUIzoIfNyYl5KyE+mk3l+jcCJkjYJy0zb9e7IrlMc2
qbGYNiwT1FQasxgWaDEizpZ1UlNxKOZC0RBnZzpPOZ4H0SVVN/RseHoDv5853z24
Mc+obPbUclnH2QU/zm+jBuxlsXCUDPl45LcFzndjovrmuHZ4Q5X2pzfAqeYAFaYw
MHWIC8IesOQNT2aAJZGyG2xKXeEivXgTq9XBNoIbL6eCKjGfPSuaAfHRYqrb1a2C
JSLQlrjTrITmREM/rJTR1IAyXpAciQCCbv2HL4kmeBbUtOcHCOqbDWymD0d8y2nJ
QzdtQlgC6nBmThvCaOTpEOeXGODcoT+WT9a2e4mH00p4NfvL44r1YdwtFEXDtuQL
`protect END_PROTECTED
