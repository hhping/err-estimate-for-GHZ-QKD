`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nHjHw78HDx41p7C7l4KCFGmTAISdQfN7ami0Oq9HRMDe3mEpYNyDkB8woIskEhJ
C0XjNrX8DJ9sz5D6vzx89ebi7kBmoNKaql6whac2zF2e3SBlHdWb9YbwEqsD02HY
juG2zkRpk5a3CGI6KZpILELeJXS05sEaQT+solRPQW1wjQPdwBXFQOlJpmMVMGIJ
4q0Q8tUVvhXO7HG6igUcUPeEpTxCDHIckI71IkEEM1i9o+2eS6RGjSE3HmmQ8FIE
AtIFteLq6uY8WZKuLou2EDayG3bV/sgjM9NYATKRarUBhbw5k8GC47LIxME8qx5a
GsDMHMTDMf0Eea0FPPhcx3Z/esYSj82B7hiijkpq1XGvkCenZzyVVXe/7Kxblrv9
Td91cnra/fl1BJsHpD0y0XwZX+FUQCE/6sgnRHlH1pXffQjFgr//43a2m/tkPrm6
zKvglfx2e/HmIDEVI4LnX4G2lUf/7wQtMyRkcKymQjscmemTb+zusZvlPGlvof3T
rgwsX6EusYENZiJM7tItaOQpfT+XdTWr4QZOlEhBEe2CCQLKb7WqkaAYZfM1FZrA
50CDVpEL2lmuPgZ6koaTTOEbjyAQ4NJQFPmQe/NCzMBDjyDkzoq7+Rw+Cj3RGYnf
NN87skan6qa7bW4SkWcXFuv0QQElqfOTk5JJPj8CgeZ4BciBuGDn1Uo5/7JaUUEJ
1IkH0ZunFHkr4082y0/Cn76eOOlJeu6E0IPaVG/Vs6WCnzM9cmskS1WkWZULgbs0
+o4JiXxv4CDjDJyLjTKEfe4XwMvIgcgx+qL5gCnslDNHQM/CLHu8krjG7IITuy/x
kEUuKiXl2CeQ/bljeZJw6rWORs6CdQqGg7bVkkeub5gghZrJXC3wfuWBEt54bW7B
JBKNmhtS5dW5eOU9VmiVmNzp9rJ8KnxBlGR8fPzNpDRoVMLm5bNviv6dCLcL1sCp
qe70jAZRbDgOKfYaHJfHj1IAikyNcBNv1WxGOmoctiMjIE8nAftbG1lTd1QsqkHx
ywXnmOHa6QVSb2lUHtEYPMS3n8YTLn5qQ1bOuRB5M0tklDVs6SXepiDARY/u84Xl
Du+fH93dCp0SSgMqU6XlLmKblXZ5d3VWC3hEsc3tvHcf9ne/JCZUm2b8Ta9O6Ah+
qquSrI3yYb7/z9CQUMmoa2kclcvSatsfee/XicCPMXI+OoAHnL2Qpa1HneRjgEyv
uPJvzPmve2lN3dwWJJbZEuawjXclZUa3EM3RBQcdHQjqR9kavHEuocTZy/bWzR7/
UmtlMGmFK3ETX9fNHE0vuEUWbZaKJjjW/4JCE8hlFuO7+RAdzeBMlrUKdy5SjtwC
ZFQMuIGiHB75CxHKKWSuPKUc7W3K8mxvwrIK+2PDQyc=
`protect END_PROTECTED
