`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79kONs7aS5GO7PMPqyBsGgF73sfq7Izh/xNMU/dyk11xt+i4bKQb+T/Q1i8clHDZ
6wALR5nXyuL9m+xpo1RuzVeXIFU3ubABwD3VymGfhZ7RF0z8MRxvhUm9cl2CzMQs
vuQqEISkFjGwVCNL1gvV9LbGxdssactyR1cx5mowaKBQaNoMshtbAbKY6NiHvKZd
XABXcMz3MdXX6H6Wcpvyzv/EkbqagVNrki2UnHjJoOmC4pGrRIkeDf9jsTeVlXgD
Y9cHN+TYAV4WXFJTgpizlBp1l6zUpDWDRUaYZ1nwcdLPTamOcUmKqK50K8ZbGDs1
u26/Po77pVNaYUJBhk8ZKphgxkFYhmzigLydbicD9kE+iry62VziY8ipoYj+cPP9
6EqTBD0otwBizbZCSsh3UkZti9S/VVXRcD7cIsVueMPWuzuh4pZ3HQYhVGUwuX1n
5Ot+97pap1WNULdv8reK5Pw80ktJvFq9ckl1T0nOl4lJa4AhpBXkPX4QR3i9r3sn
r+02L6PgZWYSmuBOXXe0l3e6Ho8AykgS44s5cDdXbsPqXgKdLHd8E0FzmyBySrnu
b7f1oua7d5U2EDIIIONnDThQmUrLk75/qVI50pYZU+HEzXdbGQrrC11ZyEZx3HSw
ShtBQc18+HwkxBl7MuAm0XUDbz4qbu7vvodtzN6Uu9PFGDRIiCzgbXQn0X+33ZzW
ShtkRqwQUBc76aClWVbeRN8kvlNsEDIbutoNOVDf5l4dE+5mC8z+ZXDdXN7u2e6w
XLJq7tFlL5U9Jqmq6VFOKoZRVIIJFyrWJhtFIU75YIERtnULexuUM/GGXuimUSyj
nojH+vwsKGTEiEzsn5YV+CKb+qz0eupbCtA/zHk2nHZVRrTiOZLXDW+JXg07NQwf
MTe7hAvHU4hn3ScbZwKKs5pagyVp8eP5HuEGab3pnrhEWVBk48ChQ2JDiu56Z0pE
nCLAIXtr49io06NZU7A6Ps9BFlULni4KarUlXbdQ5uaPPPw31/tYa7sQE7XKl6l0
3ZXnQADGJaPW0UJ71LHLSryObTSg78bVKA+Fw4F2eGaW+IjwG/ocFJnaswA6ZIj5
i4PcGejHGV6Kf0FWGaexRA19Uw3BvuiriHTb9yhMUq9tPFTvZXwqYp0gMf1ypsI+
cbjE1qAQlLtr1snIZ4OftmbxtTl978iZlZ2bT5Mnmo0Q4GKb+HHNMBu9hapiV5AM
TEX8mO0TD8gyBqURc7rRr9NJ1hxte1krEmWOKcpUME8wCY/QoY5bj+R1zsoQclGq
/FkKQLKrErWLmuIxN0BiTSd6UY4SzHs1qQjDRkNt6iTa0WWZgyR1MMhFO8Q8QWES
HvG0YcsFidk8kNmDfE9ee4yGDjD29XWryibIs4mD2jRdLgVCfObUh+4xtZpjxXAT
DJFewP5poyA+J63+jbq8vzWLz6/9+t0dgWIc2hVmVy3J4QcfPJq4hTTSsaV/m2sE
Bt/IJf/hXGsTfkkh52Q7Gmk5PatkZvi9jVp0t4ezjzAVwynM/G/Iup1xhIRB1b7q
IXZfcQU6IA8gUz4KfO22Ib4gkhDqcPU5CE/uhMW5WPPJL+t69mkdZNe3TN1M4Syz
yltooes+MzPix9msNVWGQaJB/W+KM1n+l7YgU25vPFTRUp8abovU236xqHaPeeue
bp+ZSzhFi6AlIDDkfUBDScsznFnRC/k7TsSSjZaZbb/o/0AuX8Ss+8ZTv6/LYpO9
IlCpe0Hw3QECspCpKLoVFKqPxsTVQzfPIk34LZv8hN7UCqztGOV69Zkm6E5+Qkto
lpPd4d+LbpZ3Wn4TuqBNJRC6uRHVs2/PQtkhCjyOuQRAlfQYVmOWnc+ybqxurc5A
zH1OlCZVGZrrBuT7lRSEfHnc3eQOyTDbsVen/bg5CnqV0Fv3GaNu3n6AMGrPVr5y
XJ9BgcO/H0xVBfqH65Pyn0cuLmetxz8+2gYiHj6X2ji/B71HXRHCSEUcaPXn7DPb
SNBlEAz1kCk1SXMz6E6NccNBGM6gevwr7Bz5Gq3ref4K7VOK9VopAtiGTFKJHCot
/MIsYzDqy6XgQWY9Tz21EU1eMMk2pwaXKsCqYObBhAcPrCiNlRn594S/qQSI7IAD
4QtudgQ3zRGyfKy04isiepMRdju3WWKNkpc+q+y+CiM5WxKJPgRPsHKuqVpiKWQ/
9mGVCQgDeDZ8lH3ATZSCOeC4ylXCUFO8EAqi+QPNckwa6+QUFB3DyqUpyR9Hwl2j
e0bhNyEhMt3yQs6sD041EnBz2KYmxMam4EKy9VeR1Ua98ef7AYz2TZeHB/l3Y6FW
W4Bsh17l0wSRCpjwwt1Jap7vtKzLiU79ymvClp3SHZeXYEKLnyMXJmkjT4FTAvt2
NchB38kPevnifHr0f4OUae+Hbio5vsymH0ECdbYZAchtfbZv7uLDsL0zbiMrKsSx
bXyTJieUcuD/7LTiVgMYP/58SVi3/Rbx7AMfFAu2WA6ydJync+og8SJUaRJvotHw
PJ4ogIDnQ545rcI28CfIk/WdvFwgXaoIEpdr4TvPknc=
`protect END_PROTECTED
