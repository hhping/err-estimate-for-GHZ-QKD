`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFtSYxQmNq+i9yJcTm/+0vzlGZlozqSgQBmb6VD7gcVv2GEDGUoI4ZowR45abu8f
HkcKGlel+o3pqzYFhsx1mRXkOsqcWLPDKTGYXEPqN+ddJcyom6vBLLU10MaY/eLW
K8mM3xBt0gaiso8ckESngXs0Ccx+oxiZ8ezg5rbkxUtbD6ebD1c9lZh74UwdoN9j
GZWQneErrxPpuIWYQJWtGqGvd/EodddNeHS85lKT0k5smt0GndoPJx32xFx6GTK4
9pSdEJDIxh9TlS0oKfqBkWa73XYgEE7ou0MIEZCkHNE3Qdn86qW28G7DrXYpZN2k
p1h4uVLSflA40wpvw+oPWK/aoHNpIwgfhAeaZXLEclPS64SYNY3AgzAD1ZMO5MQm
FEEe/YC2JM77a9FUKIOqcYKIZu5HiX/NLuhZhgvA2FJtlhl4mxaXV1pRbrpvbj2c
jE98QHy5IB/xlNolHc02o8X6a3ozVMvx1Qfe4Sh00IA9Yd1/n59U4WXwb64XWaOc
7Hm95PZhC5zEN5kG+I9qSI/OBVVVKduapUgKKpUk1GpoMDUlFFFb2K9P5JSABMpU
/P8ch47+ldG8TkKOg5WInp7KfB9tVYmTij9QYk0n3VbvVFOzopi5+keBeNdG9bap
zc6LB0OQSZTwTJOw+2RQsJ7P8syr20vjyCURmqX5deTg9IgNLQyGxehYXsU/V7y/
p//gQHlyDxYin3Eq5t91PiSWWejbB3LFn/IO0r+XSOQ6NtfzBXqWG5KFXAi+uIaV
zSbf+tUHh3U8tRYhCvy0HfJXDMFVZrjfOCwRnbchDuLu7awXnZj8VibU1QzMgt3G
cU+KEzoHFRf51OtcGGVDsmMSAqoDDV1ol4br0/XeZPbekj2Irg1Sf1NXIwVmdGIE
rt2bMx0VbI2Kk+y1mcP8jP2i0NbBr4GCPvAtBRh1klhPzZEUPmP3ppWWOueM660H
qdd9nYdkg2gewZklaEsaK/IJAfc7+PTRwVJxjSpa3n2pS/LHYHgjDggv0ynWn9+X
q/Dx7gtmxOS4UsmCRnE1V4vC9g+38XBpXp9v+ApI1VL6RqKtla6eJW2xBxOPBG4G
J5YuVe1TBEg3u2qijUjpbgs9GzxZSm9SlwzQeFAimRq/ROfzl1ZispvuqUwI+TK7
MCfSXcKK2zdmKl0BxtuqiJnlsfRP2JICUSA4pSsJFy04lsvxhiOwAtrS2Z5Hn3GB
4JsTgK30KHDQ/+PYZfY2NX+XZy/Ox9Oj5D2udz9ygh8SWY7Hx6v4+KVqkYYN7LxI
azvGdptxNtlcMR8u6EZ2LLCIjWGXskuScrJbCq4ZIPVWmNV/0d6S9C2t/oyQwqOd
TPCTN8qDZO5gUcnqnW51/po7cpr+xPDYocCvYlKLrzLTI0HK50PCJeCKvZt1HHMZ
SGdpL9nEVfj4j7RICaARLly7dMiY/3PxKoV/Lw7Qw32DujU/8GazpVVSlzksNi4J
CdtIawy8CRUAIwB6ZYp8xRV/bpH8XrcFxT7En3H2pkBjmloyEKVnAFsgYIYG8ROl
qgV6aGO99JY/dco1HU7x3uGkZJ1gETgeZEykbdeElymXareyCKGKBpgMC6N36/o0
iBYKiA9aMR2Ytsp94Q78vpqNJJeLBgYatl2XEkB8W9Dmpuje1ZHdF6/tAf/BM0Qy
65lOlihQTdcy2rpWdaWDJD2m43hb84eyBaIlPbluPIgsGeGIXpVlq+4A6uGSqLmy
vY/tN/2anOftUwqIYgqNiKKlPKUfvYTOVxSqUzW3HIGCsDMWUit3VpB9oDm8D++m
cFy4a9Fqb7ktJkCx0iTPGFBL2IAP8u/41Hqh1ZPySIbgqqiiSKK3A7YgI83/hDh/
lS8TkkKvwa3aBel/4ZA7YhqLcCAld8J1b+c7acrm0rokGO9Uu3EKZ0GKHqmeqt33
kVCb/+0SfGj8E6Ei5OSKwuZhvgNPAnRNqSJ9jFgFvoKT4pIQlWX/gLN9KV1uX8DE
n99N+pl9Bt6dTo3G+9rYDa4ZidlIHD7h2d+ac0sZJ6WUal7c9Y16Sx1a3BdDYrVe
8rwUDBnPof0TDal5NYZOVl4EEjIV4DHHUFvWT84t9UXJYbzf73ZKRkZ5GQR7zShy
Lb3PfZGaaPIvZg38IoV/IoUEYlZvaK3UyIYqBJsGpoCZP4J9T3SdxTwd5+l1EFX2
FdvLu35YH7H2fDVBP5Dvmx2ZqdJ2eZoNjRXixgQNNd3q1dmoJPEIPLdA/QoW1M85
pXKTvY26b5z8MTvMVMBsEfEmpCfaWHOJSGy2ZyhYnPajMVsLeHUrLpH8vsXOYHoa
75AaoIlN/TM81szlANE+z1DrTvHK6xd9sDa+83IlBzS2Zp1ezJtp6g13XeoA+Iy4
zN52qRwEk0jqL+la8Irej/AmBId+76aNVpzKn1lTUlVTTBw+k+j2QhCCTld0Eumq
Z1+HszyHXd6zFPKPtLF9f6FCPRhi5l5RND8EtjPt6WAUG78Le6KV4VrwJOxV7grx
SB5lKssZeXOk0bVub9IoR2S8aCgs2J+B2a75APF4fRdut89tCf9ejr42b+csgQpd
gJ6qP9ImVfN0bh08sSgP+K6OtV/GcE1iz+fmPLk00Jnjctz4EWOJFG4wUM8Wjvt7
BvvcaFjhLNFnMobqdcwaFQ==
`protect END_PROTECTED
