`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOWyBo2i3GKJH964ad5pyguQJWvwOZbgp8yN4QHUFDWnTHoOKIvKSVTDAAcze0LZ
JS7rf20ywhGDuzfxTaKMdPxDsBJze8MlLdH2Cs4afQ9LONZFFcjwYR7txQAj4424
W4m6yzQxlveS/U54nrQJEtChYAMQr+GcBpu1gGdVkjt8DWlF1gXWEzYyaCz7NzvQ
2SCWw+x0nbabvE64PEfg5Bhh7NfqvkAKuGvdB3YEkS04beymSzLuuSSOUm2Hc8Jg
gW/k7VQPA7jniuuItFUEX4l7gUR0tAJO+pS3QaSk8J35y6Dk0d3g1J5f+9yQ7IZA
w9cCzbvmgQtdZGC4cbI2D4PJxSPrj/mUr4W/g74Uv0EdV13DHHxrviLC/NhQWHmb
Q/wwJzABPIGnp6lPVNwbRvidrHhSFvql4jh2Z5GzSW7eCUa6biSYqgykLjuxdQyT
NWjIlZ74eJGw2wBdmAOTgud2hCrGCwEG+J8k3QBeZUF8SWHJgpRf7/X65oJ7GraQ
bNxZtDd3kkyWFtIpZY9y8Ibb0LQdJgEaguNDlM95w69As033rez42KzCY39ZOL0r
Bw7z9lZyQVP/cHBd9IVsOjz1RtxQyV8bXzE/7NIh5GWxOM7NSXH+MgNucqIhFLl/
ydiV3Y+mU7lORwqfWkFj5pD2wf34z6SOqBx0c9naLxKzRN/nuaF6+mrq3PlOyu9e
GG58kYMCJ3FYyHaNYmwvtNTaPwCntDOb0U7bfX89NLhtA6gorU/9lXYZb8TskZfy
ySelXNgLDXSpWceFDMbF5j+7r+n0RH1ISKsOid9Nw/YZzxzY2r/v7rwuIg74FDbg
sfu/cSjAHMRhm+9VDmUVV+6CS+QpF1c4SDYgvrUi7HC3ZbYomao4nm5u+WXm4x3A
c7WELYcWoGVORazh/vNfCD9ppYYB+Qk8D3/QCc0FxyDj4KRbf1R0o/3qsrDB2ipA
+A7LDtHMjPdwhdc/7XnDuAdXMZpbKzQnhegoE9otXVLOlsnrPyRS1DBIi8fKU0LU
lP0h2B9QSYCvOyEavjG6eguxkiBRzs2Gvjw+EUSrL2AEDKFv3Lxu4mtXo33RfZ+H
dWYQ98PV18oMhBAe+MtMPXNiT+ONs1vxWipg+rpRvh/XmMMAbNEm5FEDwzkq+D75
Cl3bF2i1jOwhDAhGhFjPG4S9XYeiX6NOKnMW3lOlooiT8Y9j5YI41kVjpBsiu2vS
kh1QV8TPeUhcKT7HmY7ygAETZBb1ozvpV53PPkdBsk0NBL6HkaVoJCyJo2ynoTHp
w6ImyEszTKcVFOoPSNfSxQ==
`protect END_PROTECTED
