`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lSrQSla+YipCewEWtS7462aBGToSi7qKOs5+J6tIwlIJmCKs/7Z9/FtdiYac8XRq
Pg3HtevsdKKYIpjPbGN/nWhsBv7HK2G1/jBqgODnsDkpPRtGjhq3y0n7d3GzrT+3
0Mwld9/8AcDm+/UzN7fQdi+TZWdW1iEFqkEA/SKQbSoPhkwFlysvG2dIP9w3v5Rq
5KTo5HmJazf7qQqyFHxXSqxueDQ/y1R7Jv88k5n6iPA1QagDdMH8V9BLpsJlGmBI
sLTTCyZ5nYIVaLIoYP6VS7FisB7aLJtjycLr0f4hT7BEoujzOHqPPuRmX1+8QBsN
ufZ1tpEFUls1BpX3E0JatRI4/tWSWU2Il+a9IPt+ZZO0tLQPP+DXtmMt8DZlueoJ
GP9EoGLijjmNbxsVsLr0nlsRpx6Q6Z9L4oG49h5iZ32MbHy4uny+Hawpz/reSAkQ
RpGWf1QYKkohzPV10H+JKQszjs9SWp0+bQcf9oDeT6ymTUJXeXzE/5BbcGjBmz1S
HB63ldUbll8J0he0UMzeqYWxOvcpegg4kT+Bg1a3F3hRi+0d4jgF+yhTw/MsirvU
0gNN8V1yWLMNWqkprgz/O24QIkBSF/UrNgc6aIZyFsA5lFcZsFk42fDMVf7mnxjX
frSXlciaD0hpC0zl78HqiJNW1lvVpviL0ZcZz34rBBdpQVC0RkhrzfJ2DHW9uYVu
2NM9B5OpUiBISaD+xU4GKqoi+8F1FW+2kcs2o+mnN1Zs8c148b7hVOTeM009/Igc
KqkV54LGtn73vzrEXbVhsW+TlIrO23J/1f6r5MdTmo34nLz1W2YxFuOlfesD+zxi
1mOYz8IuNjIbrbaxFYC6TQWGUn7mMN8QTEuhxE5kg+xYcQ0NdQFY0MKoG9xxSxfH
q82vbnq+gqTZJw6xn54Li0HOIdB5zuBf6SJfoy1zFkMZmYTu/fpIi0t/CePgEDn4
vzi7jjZnqHVeW4EyoVhGchp9l4Iz8R9ParDuHBhMgzPXIrK4vy9XxILQ0Xa3wMSg
z4QfWWLH+1r+2ORLNWzCZ9kFLPeYmiAYDb3o7XvgxsLhO1RlKUEN1T2FMpJINNek
9WW7V/IDjAANcd2a7ZZB07orvsj+u3hI2b9Fk7XM1AZcC9ubiB8qt1NpsWtdsDG+
hOT5SeVx5mt0gvnOfCQmPWL4iwKAHUrGhKK6Mmd3wxwZbZPodQUTJpjl1WhPA8jw
i8Y6xIvr2xHmLL1jtwmo7LAqwmQSddeP5Mr8NdPG5uiKOAa6nSL9+L08fJH28tbP
BggOZfRqsL8it9xCto3Qp+FvXM9UdU6qic3yCHeJRvpWORPVqnCPko5KKvEQlzwz
oq9Syz+6pNODZao6s/h8ZP91MfBe+PqtmUyNn3s/ClpfJzibJfhAFu8+ERnl/E1H
1QDuuKBTzlBnQW9M15l1N5FCNTeqvY/2PkbKDq0JpNuFxDFld3TBHQhn9mJDFDzy
Teu4BU7zdFpc9VtiRP8E7V4ZxOs7nvU0rmyGpI2kszVyGtjdK2aCVnldCduQ3Oht
yKkA/cRTkM5+0l1dd+m5SE04jYcQVvFJV3aZKmRBgVglhYsZGcTCYlZUYMyMtLpI
OQC3GnP9MYPXDKZGswpf0a0djWTOEU5HWlncgGqBe6M7tV1R9AYstAsahzKss7v/
X4VCcY9iOJz71g80y3dl8DvPTQ48YVB1y7qcbgf3JoN/CxRMLAcSyOB0VFcEkh+z
lUmq053z9sEQdIR3JfoRolrgJKHUdzm/y5ymUCBuLHVx61yo0sVyLQDj4m41PboO
Yku1a/7lTwig0+4FOG5natL1F1thWpOIFhPuc8rVj5z8/Gokcm8x5C2cn4GERUg7
qbGo5G9OC9tBgrQADHKTVKM47B2DlGegYVl3xtfmHCcDpzyd+iYjKQpFfzjUTSME
q9HP7r8WeffECwms5lY7n4ZpOQ69rcgH5S4qLioL4jTZUc8XMkDMDcFELbOsJAF1
Cm4KYR/SB3iteTzNMGg39iJwZt6dyRj4bfZqTZS0RT/+D4dixzMaJzNxSdtgL5KJ
ZusRF3gVj0byucpitIbYtaHCPNloU6sUIjOBVZePlUwkHAov3fxyG6793yRM9NFa
I6q923wjcxwBiaWLYyAT0t0CMgsni7e6NaZOJ+iEkqP8eBKkZJOfht5DtfrkHKRC
p0C8cHu4j1ll/CyeHWJjTMqroLVeWL0osrxnoKaM511sz5yT0GThFc+M7GL+fify
UuxAk/zo0ufNJkjejdo5Tf7/tigEa90DQHSKJaDe+odVUbkiY9AXKH9HGYvX6lxH
x1WfSBhfvGiL3Y5SZ4OstwduT6yeY72bd++tc1yh5kcG3Vgi3nftm7p2LP6NulkQ
YzZ6fItaZWBcfum0qhCbNdIHh5eQiBTgvWiaK69EECsTcw//9xeGB96J7PnkC344
Vpu7OSITxK8xc/KTQDP+niS5B3ii0432to0+u/g7rS3pL8ITvMufhw0s/5lnja5j
UvJEpf0YIHmvpKE/CAw4yQOqGTezxY/BxCVZbWDn9bfj9hy6tX8V4m4i/RQukX70
2XtuvWGn6iNP3RNroMF1RuwwWja3Xjie2KcPBvopN8+6szr2moeUZq0iXBpFE8+N
TKhCjeZeRhBCIIG4dxOUQJQ2apwvXWz+OXg22ohuD8aMpP79LhD3R+3tlIFZYhVZ
G63ElzizffjUryOVmFiFDstlVB1JWGLph6nFENaxQDqmwCBW8mxgEBKSu3vXDgeS
fFXCWroLuXPHGMR/es3FeLqgSedvQrDFWvh5dLeC9fWzcPSVm2WU8bFXiP613Ldu
LATJIfHSBTwMEsX/MoZbe/Q6XnhEDV349vWo6pieHstGwyjv5xvhoWbX1La+LQSr
B5BpQ9Cq66/kgBpkJHkmd3kbawben5W0zX1k190cOX6NYnCC5mMvx19RaSN/ZmVv
cl/fgDfOnuODnF2RIOOyBnLwJDYF3bvoZn2PksGwpGBYWliV3Bp107doWu5tyCxa
71Eawj864eOcLB9wWdD/pP7aA67dNecu2Xi6EJJS+0TCEpFiym5X9+jZ/goeACLn
YCyyZT8AOhayMNvvWen9aUvcXoOHLPWrGvb993jpR3aUeI9Ys+nkJ8EDdaD3o7jr
t0jwlbGb9ufrbKaUE8aegynTR4JjE3IVMyiNvw/1aIZW5wpla+Pa1/zWqHc6VKNY
bMq+xISffuIoMmaGjPHxZxUlTEoHR62MoHyTVFrovK0fZkbuumscD4PIq+RWc2rT
nDR0AlGU4PBUlVOzyTyvlSYNFkV5tjDTTSfkdJecsz+/ut1OsK0Ks8+78oWMimNw
0qVCNai6YOz17UTfxC9svM3C07unVSiII4oxmwEQ3wH+yxSPtA2xo2Ku0WbxJcnt
vyzwN4TiJDL7R+NfncT5AyCCdSSvVfXrA9Jfq0Oda3fW6qIl44Yzzpw6GMqgyV2K
HIp584ypd4mZOOIgXW1Zva66M2gQMA1RtrAHpwSXbr6des1YXxII1dvWh53uiVFN
ENcHNJAPHIhDzvod80K46Y+y+MrO+Qm8aIP/o/3JdtB85aeZSdkCwrtBR/3XkNQm
JKNVLiqV5XslCqhA/lqxENVBstk9clnG3CxtLlGvNXJWG1+tYWV9YyjiEdrymAHC
I++WbOCcxetRsClIsnw62XTNzp5FylNHis5CUbqrung9b/oyEvCu5jES1YfBGlIL
HToYSpq7LWRrquHJQuMuuroLVNr4Fiq3UNrZCmT8cEYaLRWUfF556wsrbPwbWz3+
Sc6oq6rsdYeEHsROlYv9egEbYeuTKN3ComU7pEuf/7nWo2ewD7yj+EWgjTkadZEa
+9oT+hteeoE9jqiC7Ev2yLIqUMTzyEMRFQlDqQG4sbhMLQguzraNYUH62/JgsaA8
vWy49+Z1WzZkS0m7Zc/305oCOCdkOMAhkcvavg90y11+BUvJ/LVv3C42C43lOhij
wQlG2pjYxHbB/Yn/5fenAZ1yVtmKvlxyznlA5t+uUGiqp77cTqYrrCxrHMUVnpXX
xkBjdUSaFGpu7CjiPHrgzP3gZltVzxuq0DW1isK/zSxzt5sEdrIFakqq2tC5bMsI
CTNrXNe7fFHiINuOWPEAWxC3gVJfILQBePpqtk5E5dZpvMVvaaz9SbsINKXxsoNK
CqsnLJVWLpwYiD1pPGmwZaEU1PM7ut+q6GCb0kxhiuTV0JnYIoVwGneEVUdm3mg5
p+ZoTlzQQhqKwY2W7yHokOcCkbdTFLnU4rb19pwrZ57qiLrZIFd7VAHVNAP1Y1ga
nZ/wApSDXS8kdr4+uf3r14xP6uYl2oLxNB2i0WtzFqG7b8TWNSHBWbtnBygdKcVA
VhQbF5s50RzfbUIANfcSqiUyo4an/7mWjvHdCNO5WHCWycBotO9/VUYlV34liHHL
XsO2K6n/IKDsnBoS37V0LUuPMsXQbawIvzbCHOTYHFlwnDBRNCrDgTYpBzkQW66H
/Zcf0oRBm3r900l+XOMRSBpQmmRI894AbY/nJd3sju0+XJsw/mb4C5+X7VSOiTv7
vSCEGCV9+JnIAJo3PDD+OM5rvZHXBX43Yz8uZRQyRLNYfncvMUIjrxN/HlACUoUL
8gxzhls8ey6cZcsmJzOFkWNCVcccq5WYofuODFWnoRUygBc6ff5Aa0KRPS0OG2Pk
`protect END_PROTECTED
