`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ryfkBELbYWsBoUIMMc7MnWmRv5Kkd1mXYR/aAjGcwOWg2CgUZbU+fL9cXcbpO2rd
Rr9fagQtDfHhO+31cayCgrh7KWNABN3PM8i0vl2TFovY7oBgy/1D5UjyXj6hlPSv
s2YOPpjxsb/+iaLMMWURWJXSUfrWsfVWho0Gt+CixN21PcMAkmPer/vQWixo+Ibj
6N93p4P6Yv+437cbXEjlXtnYzUfE0SXZRoSbD5cHE8SJcH951GLdBEFJGgBvGA0G
caHGEdPlhOJlBUM3cABywgkFBoVvH8oUEq5F/D1icKLTuhDFKP+Kucy2IlKB+s//
aN769uQfc6VEkyvn3A9qg7mxTa/Rp/M5v3P6pgO6Bm5tgwB+Wew2/dszfi0haPj5
1LsfN4KzQnEioJ1FOZoLirnXTYPVpflnMSAwY9sX/MscgxPea7YgimIpoT8uM76C
xN90pdR+v+WHbIhj8/6IefWcZQGH9uuksesFPY3HOUaZ/9NBiFy9i7PJYmR9Jg0F
0q5sL0xdMVEQLzsV4GT6/hl2l0u6NhHwjA9xYbTdHYaqCy8E2bfoS2H2VCogeohu
WU7mDkUlcBqD+aZI6Qyj0Gn5Srjw1bsPV2IBDYY7E3/1izlKxFY4cMv22ucL8SR9
leOdKjZOcJNqi4mvu7ma48HoZNcpuDulr9NhXrd4sIRCF2LNVHdezhxe+8ND0CXU
IvQGouAdqpNVK5OrPdi38YE9J59hQnedOQ7TqCd3iJxU5hu4ra8TX+8+vNrzBGvz
cM/3SsxELX8YKCmoVn9m0gy4AAuEBi93uGxoeLeK7ZJhD4/SiYwIH3+vASqnUdyp
1Dy5SIsXYgonRbS5ucOsyaEqNE2WXHZigu/VKeyMOVqETJaic6Ks9h+LV+YMxJB4
avoipiI3uoy2/xnh+ikIyeR1CBPwEwaSMcdVLcmiCoyR10whuU1a6HYP5ztz6DYf
86NlwK+nkwBmSSMFijlq5jBgfPmtBAnLyDMjxURpef8xirNuut1OnJorZXH+4VtR
lfJZJTPiXYiQuY/Yvc04JQBi1KuicuDw3BKyuNFY06vtC676+wg0/pbRBHZjWjJb
kOCV1+LeWsqYOfJx96HaZsdfuvFhG6jin/1g0+l8u9Na1jhhoKhaOmhmF4QovsvJ
VD34luuC88vT+DXAFfoHnkcg9B+Cg2N+jLB/pX8fuBabfM9bbIQoUrEZRm3oOTUS
dEHElcw/qkrIuqtqXsz+2SkGDcU2eCoHhyqwkzVs+WcvPp2lS7X4Hko+eWqnHBjY
zh2JxTMhWTRi1JZKINXp5pm5ToEyKb0VRJOIyrb8LZzv9+SjYl5j6RjXV6oblZOc
Tk3SnldKnNpRyJDaPoTqoiSwAaxb2F6862tgfynsTD8AQg7l+lpxCe5XAGubxHoj
x0ZGyrQ50UQ3awB/NSPfH0WsJ3m5EKJ5QwVHiy6fDQY=
`protect END_PROTECTED
