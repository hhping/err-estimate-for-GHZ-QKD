`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q9oMJIkLBHMcB3LDr0pNh5qlLSpj9V3FstaCNaYSj6xILdAMLwgs3q0JpNXP1ff+
HvkWLeqplxWSyaMstsWynjVgPfbMg4fNqKbleBuuN1PkoQRBN2FC8s7tnTRcUkDy
EJ03ImhlPqeaGKIgN5vA1KajkMNCPlK9m/VTEVq6MX03vvAFkaqVWMjIaxucG2Qw
zEqpnQZiVOFxKd+jc6XjFpc4SiCtZ24YvSSE9GDvs26tEdsm4HcnD3V6HMtjHx0M
aKdKvvghjrbughnyyKREOeDmIVbSkdaEJX5NDivtpjFIvdNjNc76JQxFhK7GNeS+
4bfPmriGlPaMEdmlSWhkMSTwpvpXB8rsaZnDHrUQKlU=
`protect END_PROTECTED
