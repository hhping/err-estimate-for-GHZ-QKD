`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/k2jmthWE6VNpBY4g3gHvqkuFivKBS6g8jeOAYZL9Viq5Ylw4wzfiOqdsFEtgnlO
RSzbWZE7s9hKOMM60s9On1aecaTJNZrFpFxLubTkD9vj/akF8RcmauLp+LYw0qp/
h6xI0/QP3kv8VZVx80W+TybNp3/o/t0/5LDFhCufFkWZhyZpY7eExmBk+tzOBlg/
yK3zrvuINl6Qfb3bOYlH0AdJLkW6QQwDw11bNiZyHyzHP9pZzwXuQdDWj0/oUOpK
Y/W6kiXhlW/P/zLIDb11Ua4YbAMGVnIkROukrgV45WjVb2Snwrw7UWlrZZxvsJMQ
Sgb8/OW2FT6/kT1ryRVjvopBLbC6MuhvwR1UftLfKm4KKiclfJrsfWX58EMBDipH
jGEvXJ4ZzA6HGvdTsYnmseQP8hld9GPNZL8iQN3nX0Tto3uoC+jizpQjvB6tRLbl
VFStKDqDUYFikFTNeizKhu0h2Crh8jWMchs9uXHn9K1q/1AInH6MuKSZxEdvSfqK
FwpdbkpBYs7W6HkTVeTHRFIAl7U0z8oz+1xmsnsJF8cuxC/LDtPzSJ5h3PMIYGjt
KXHoo6D4ymA/zETnjy9YpzkhSXjr7X1UL4t8ZgvfhOPbNqCgf34Jt+4Rfztelyy5
M1Nrpj5pToJjWxh8NVEq7BFAIHB8VySBqYIDGXj1cKY0vA+Lc5NUyxMv8AyQgRBP
TYe35e2tG8fFH4BTF0KUc58qe/JzHocATWDF9OGMIEaPXaOz2tmwUQe+wS5xYo2E
BCSj6YJT4ixc82nzz0HvDJL5FC8QlhLd1TV8q2wGStEyhnmNXoqeivtZiiACXIIj
nA9cQ2zIEJs3MGPVFLOIxefnAmUw56pEf3HEm7mChlYmUsP68nodcK0VzyYO1Z0I
iAeDkBJ672YhYR2c4DL8unBt73CQk5N6pfE3To1OaKd4gLYyRRjOJ4Y6sE+cF1nX
Sje4oW1S8ZflIdLCwAEaIAlIkqgDaoRIOD9sb8ggtFfrx3/+vhrfWPcpwW7KfRxk
ZEaHLQJFNKpjjElDm5LM1DiWGEG2dsTT+5ArobIerEWed0F+1Yf+uDBwJINcBpwD
Ohc3hsS9EfaiFxsgWSyTD2UZwvCP9AaNuTBBieE89jcJAdfxw2xYowLNV0Iy7u6f
tCbqGAytqtfa2VooTIbtBWXZPVvfx4STT7kQ2rxe1zcUZ57KviwGs5t29pTb5QVY
40Oyh/DXc6SB0csYjsqI5uBZ3Iugsglbg3pT7jsXkXJURBg6/S7A9UD5s4gcrNh+
5BtnJwddme+7SpOwUB1OWGlJEDYYeFUYt1eCeqjvB3A7kh1OvVyYOnSpEKfHRx6S
bo9Di3+tqy6auJSZQ2aYZOPhSsU0P/tHrfuDH1THXYT01c+8XwAyxX8LS7m+DPup
niKU2G9bmricKUWmWkl0Ra7ydMiB64vlLoK137R4ho9uhdyauhPudi7Q9QUhkIO4
AE0Q7eODFHQjn9DqoCtN/CIJ2fkWPhsPW6YHgO0tXgBDu1i6YjjooMmUD6ZifBai
1i+36VphSicq/vvN73tzykXQyC8Q48Vy9FrktKTMTQvNvH2U6sVXxNZpP7IkrOHD
Yz3+U8mkeI3FRt0VNSIrEBZNFaOSEbYGS8MQvVNTCaHZAZQGdDRMgC9eZOTQquLL
HbVxLhgEjuzbu3k6u2LkF3DWyKMWmPuasRBQzarx0agUhWWKN999Atlqkr7YpSFu
L2q1dqWah8ygjhYErqPM63M3lX81BzzKKP4UemPIHatmpY+7E9jg3eF9kkhrvhQF
XjxImzED+gLmaTUUbnxDf2LqKhhiC+b7n12zoY4oT+zCViZ8EGXWd/kcRepRSSQO
GPatsbJB/p9xiaMDFkK9/VqRCMoViqwBpjyqZxHXy0owkR3Ckd8TVYvv5BFWLRCZ
WQo/bKglXZU5gz+RJA9DOnF3Tt7mLbkJ+zVAjzCNW9G5Mz/NcxbWC9vD9RdyoTbV
WjzLNKiTw5DfrVbbI+zxng==
`protect END_PROTECTED
