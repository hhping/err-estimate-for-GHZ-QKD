`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SLF5qFvDNtQtP+QTgdD1t//xeyJlgC/PrO0pc0lCzmi0iNwRlCZiZSzIGLcfS52b
grHMgM+T+L2WnuRJrZD8VKDIV7YOK1Hb1ylW2pVtcN+YFSO3TUixeITa4t2zxUdy
rzBc96pSGXAS4mN/ubYdkWNnXnFw1jie2gp5xIB1/dOcx2HOQomQ5BnBic1VyyJ7
XDPVQ7peW+NSd+Q3uJt49PULPidfbHS2L0PJNuHkohIA86FHTGz2GLa1ojxUFhzK
6simiNmxLAzsUT8YXJ7J/DcK5t+s4buAe2Weo66AXoihe5xzoQlT8eiBMUow+vsw
eS3eePXoZhNuFycWUJKvlAQ1xV2BSyy7H3UK73dl5NVnz64p/ov66oXxG6nPXR+2
y5++Q/jYIl32V27o5Ax42An6E+wP3pRCERiWipieFujlULtxwx5fcWuFtUQhA8j9
DNMiu/k+FSoCPnPe6baPEWIatAOFT/le+ru5YdP1ovj1BrHp3/RA3eb+aNwYxEg/
ELQe3Q5JDj1kFm4WZtUUM3jpWkEn1RDyKaxzjgM6MAlth7DzFUrcsIyxJeYb0J4m
hHgRKsfV/T5+sr9ASef5ivA4OGhSeF4Hdd5JaPKtG0CQB/wtY5I6XvHBq5dK6v5q
ZJVoI6NJTxCgw4EEt+g7MPIaTMzb7jWemd2xBaAKTlgdtD2WctMCztFAaeKtsVhK
ZI+p0RLxGbJ5umQxThochiq0lfyL3eXCSVtDPYJCCul4IW7lRevMpywK6z18t4Xz
rsmx5qR1m7VjtzP14qTmr4SM+EtahGEehqz706V84CioHNqUsg96qu6cFOwg6JLe
rz0rGHPrLktnzhNReZAx8UhpnK5ysCJtj90KJMfOo3GGqughVR81syG2+D0h1DEq
ULQJ7LiPbMgpBGjq8xfnOm8DXK2r91OFD7t6YgfAcHJh1yJCzinLKmkyUxyPVpvg
LHTaCYITNLwd12ZeH9KQ8rpiSxWs0Y0LpqybY8P+XZluM3w0C+44LTfavmspJv3K
xIpImzNkwqQchdk7PBAdMGk57wF8YooZujwkURAi+hEKDEIFE93PM/I6mNNRDT2H
f+a0LebyssV6lsk4LTENFoTG0BU3fQz3eaT/di46X1JBebbNTN+5M6kpaah4s+AS
xVVN5HEyRfd8YVWjLf8oSIvbDD4d8njfYJYEaxzHtm7wG9ecbN/tgeIJcsuoZPjE
qAPtpLSO3ZFKQ5QWCx6hfFWVkl0GZDK7NUqNfX9pDWN8L7olIqBj5mSbXrhx+wfP
czII54Z2mM4EQZqFDv4zSsQb31SUqSBnq59kajwlSvMVVd5EcpgnxA4s+IPctQr1
s2oBir9ii+x8kootD/KTxsehXglv9QFwyz6sUZsOXo3yMLtNU65QBf+1TSjQL4xc
0og38eEGX6aVNfHv8UWtkf3rx86mKUx7QRRp0x4R4K+Nv8bjTsGDYXw/aE1JOI+i
BBV5wCCKs4LC41PSZy0BuqJit+6FEsxsnSD2EJnjNZh//96ZK2l4yLHZyqFTAqBs
Ihzh1MJICkgFW1l33/wDts4mSAJFAr9W47cYX8fwFF5Nzp6UGpBi8Vb7TVohC8sG
4W0JUyYYsni0Uo/FwSb/+N68zMCIoHT+MVuVNBKAMRczi2do7oIEi2Y9WhbprFCg
ONT3HzjD+b03gFE6XKx5qqzHI7Jn6rAlxPs3cDXqCbENdQlfa091OoQqHCNZ3bP+
EBPHPKZgl3sG4TRLJTv0od6QUrp7/IsWvb20oQxHlhJfDOvMbJ9HBb5rXTTs5Vu1
qsUrWvix6lFkyKzplpfwh22eB+SBIBqyV23KuA3uCIk86XPW0sUVaUXnHZCvSjDe
uC/ynYgjJj7wN7ulXJTdvNZDgfjtzpPIqoew79Nud6SKuCK8hwWbx9R5M7pqww71
EGqk9dYcwyoH7eD3rjcY3z0H4Zg1Kty6FkaJ2uzZgvBZ7+NKyq8SJWUI8qKZ7BeR
sXDPRVwJ7vBSioaYvLw204VkbkGlx7nXq6g1o7a13U/q7+A8KHfRxKFBllBd4dRN
OsSGxraZR1blUaqkIBZveFOM4VKOI+dKDq9g7CD+KQwHpmt6nFDlADTd0TT66Gag
ONtuQSj33AfkRBfGN6dlS05O/lICDhIgwa9k+UNVMLYrGEj8kpqywykpoWETCuZF
MGJmJZQKbmHuTbr5tXRXNLCiY0NBmQJN0QJGj+tFVXNfqGqzN4BdTIufjA4QAWxc
Ls2PCfTopW7po6Y4iY8WNmqdHbidsitCDnYE4TKyA0IP7ziggx/ToVW7dm4d/Cqo
CwsIGAGtRbvYlo2YCA/s/bSQ89kT0NTetWCOYr+J5KK0XQ1S5qXpCJcScF6tJYNS
ViK1JbBKBbtFqIQ8cEuW/UHxsLFzdEGDcRnujpkqkVm5afV4gFqrPg+G8tBBGXJY
sH1rFU2/mcTChckgXy4ZHYbkkqFXp2/UeG4jmioXBynhfLhuDFIrb4t7pEvsQsZA
rn4DPZhMnPdiGJPU0Xh9PSKf4KLosPSxtj57EsHtFEm/l9KKUnPak0pxzdtEYCcF
gGGfg5/FdQBhnWVIGmGasGwRujG1KUlV5I4mmJLEd+OFnNR8vmflOTeoo2oOokoI
lxHOiXAP7WJOjg9+bvwLVKmPChZuvIWIfLvXySIZ5hIGTvooKU/nD9001ONYRq8g
uCXwUeY9oZI99IJciFbcJv75ZnuTiVXw5C/nIpcIPhY48fsp/4hSaNpGZms0Nn6g
6J9oWWuou6BZgWOhCrwVQDggwVVDu8+uylQ5mSpuVN6BZxj7KxjYgsPx4+LsZrny
DXTGREOxIsH4PyKiw8mVNNVTXnSBQMSpCWJxZmAp5VMsubRCo17ntVURyPwCQYV+
GUtYitPtBqu8V1Ga7tP9p5ZxU8j2QR+PkKSkRatN+BRJ+TrJZqbkrkoFDnwUCyXm
m//XFhZLOIf7+EAlbHdaNLhu1zF8gsrhr3HcOGPRT/dzEXHMYx4ESQXuMB+hRbe3
`protect END_PROTECTED
