`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7p+nJ4JUZYajTfTFX/mnDu/IiENeUhvHGknDS9A2feClBmM+yJ1S+eHb/1kbtLdV
HOZCEMGmD33piVKnTb0+uQIPgPjZxuoK84X8e41FNdH8d9ED6LaOMgB7S6tChuQN
TRch1YBXXpPhbXHOxUaomApnyyWGV1UATxunIFsuqQPP8ciNkM8hRJvKYG//g/AF
awpCocTf1t2ErwmH9Dt2E53K7sWpYQN6tOkh+o6RueA9kiQzGtV1ixD9uPQh3dDB
jDyiTQ6vzmowbkgSt2eVtBdPzym47OzEjnpw4yyDNaGEYBDWK7KJdkQ2ABDhVAy+
sArxe+e2DHH/iPMfZ7uPk9jb0J48RC+/8PlTWqLrnk49k0tJKFTXtECcB83AZ3qE
W9Rpe35Ke52Uki5jeDbs3pW9Vn8m/Eb/LL7B3K7BKXDWZQ72Cj/s+IEfucG7Xm/0
hkh3v28dPVX/gqEezqcxyJOIYz/SP0snDp5k9hhD4sRGD+9vP0oAeLBdxqXz33ZG
ptUc7iU6g5qVAbXHXFL1MPWLJKJffUpFy1OtWlbYHGTFb0eWxtPP/aUG00kk0OoV
B/wsgevwVcKd4lOwMt3MqiadFfYUmHt5SPf1AZ7pWyMzpE0hqmhD/ECO7DfW462u
v1ArQ6oOPYmBtt90aoEJcm443sM+MXcYFIW5NWND/FOw+ZNnpYzOqq/R56M0L4gV
SbLFry4Ac0HD8f9avwyZpw==
`protect END_PROTECTED
