`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZQTfOBf+4PcKuU9GCcfHZ3vb+zy/ZWklvswbMfG86i/Z6MeeFhiIba0EkM/TcSO
oaT6RpfsdcJaBb+HSiwSDB8JDJ8Ty8vOeXx0yGcGd4M/uw9H8JnQ4hn1MfjeZZj6
UwnfmcrNXBX8NoHq7gn0uRe/BXIcI3l3UMe7AuqmBaBBU1P/KnIP/uqFnpDo5Qdo
tGELQE1rgY0RMu0NTsHVnoeHX8f2PpjUFYv7Vg8inIfQ+0b3bjH0TDRGbXPExVRi
RYBYfRXCa+qyW+5IYsBzKHNhZRlxDBnKh06hoOU2qgRvipdhC481T5CT2C6ps9tQ
KYJY7Gb6FmWqCYa5liPq+5Vq2dQVbpr8t3rzxnAZi8nGMX6Wuh1j9qPt3mRmkEUY
84/tLl7DbIJN5cgKauRmdfZq4DG657O6bK2YVvHJcmQzR2rKqTdYLQiLUx414XnN
pMH+gLGyKB4xGYao36jicrUyOWWukDmm3edhcUGHzisUAsuwtvhtAYStgfxJ6op/
skwELtRm7U9togGK4RTkdMHSR/pnCO7Hmq2mV5ecx9Dp5Iq1MN9ARGxk01ztxQUl
Xo83WogxA5NfSYJ1M16aakca1Q63MKMYNhlEG3DR23YFSEArqgAdAK47HdUJRtP0
6b56tqPXrDGrDbZt9RWgvvfv7XeyV1yHBp0uKRQZ0HDXhcAd5DY9vLcxDhLRlPFz
z8B6hKvWa8Rfk0GyvwfNM07HM+D9QfFssn+PUwLGAbBR81Cuf3VemvWfziRQP1/W
Za944U+mgVSOm71KwBuzeZcP82WBgm9bVsYWdAUYRgOQj2HWd9fvrvFHsR+4SIq9
7TEac9UyPY5FV2JdL/HGZsF4pae1s50qwcxPkdvdgH9MkWG/zQPqgHXG7S/M0s5Y
/JWONQKQpioYRmmd73mjyhurVo2a/GCK70vl69rb+j1oFq8EpXzTOnnUl//pDx5U
b34g680W+AQ+595eI4qp2qoI2BkKmFh61i9hYUKVQMUESfa+cZPvhq2mfP8+vAEy
vQM+8W0B7Po0fFZ228Xy4pN/5zInBViSDqzlQmrcpeHum04BOn7yiVgRbBkw98fO
o7n0R1KKyVZLMvAvujbLvLihhdPmMpgpnbrf+qhF01hUu6Wqv14o8utkI6Xo0vJv
GduXWKAM9rE93KSlAVR1PIZbFvNJxavicLdGdDJLOZOMvdplqxdBcLW8IWD1JWpr
2Cve2qaL0THxlVdlrR0pAaq0V5PQhOW9W2VgNjdbV6shOeyw5KVtWK7U/NiV1tk/
nkJ2zuq0mJNSXZ3z2svH5nxsiqFdNL2LYseWHI76ZtkcqSxf4jAvGZMz+qRbfxif
xBdxG6i+8uYv4e1AXb7TRN643Qs/KOAnRSXi7qETtoLqTvYNb2DcCTvLFcdn2Wak
/UIiQM/LMQ1IIyPAsKoF44J9InD8hj2cxEnla6+BgN5IsTSeLQ8K6iVVmov/SmuR
nDoD4W+ZbeK7HSHKDZKH3BfKOUb1yr8L23aLYSqyXHg=
`protect END_PROTECTED
