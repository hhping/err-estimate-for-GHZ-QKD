`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aqfwne1lgRZx8ZUXTHOfFzKqhrtVwe8bebKT6AFMBzAa357Lq3b+jGn+mp0+vwqy
havCu/DRJOXRuJ7kM1BUh93oYaSb7/JM/lzFCH6Atg7x+WNYWfs3yJChnkPSotMz
mdsrFuWdK3kCySZ/jqiv1CvJ/CyAABZ7t+6ek6ZXYRqPDheBS7lfFdFlitjdBD6t
CpU81LoQ/dfxo4G6TS+9pPTIL4BPQLzVT2pvuAR3Wen/OGTuh4rnPNqwwIbcCGo6
jpMJap2xsDkIVqOIESnryb2IcFQyji76nhqt4DgYwf0aB5OXPe0MZk7Pl7aQdX7F
LjzJjc9iybtmU4/I2TqbwcXsiuVZD8Glln2jG2MlruHqAnP0xmVuj35FOwWXPtD5
qBWFE/GSwQBMJMiECTi7Prj5pI7dNjF423WCWBU8TvWCSw1cWGpm+MH6V3fXi4mq
5iR3hAwUBqyJmTOWhD9v4Ly3m1aa+CklZyvcRfX9BADXZJ3GAg4zNyPdy1OYnf1h
5DrZHqsviLu+cPwRu/xixR22cNnMrePN+zVKFDUQnoGv9mShPmHCRkJNKrh/6YSd
yu/1AGD++KdTFORGHM3Ptw==
`protect END_PROTECTED
