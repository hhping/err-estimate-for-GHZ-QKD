`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UtWNzs1PZChAXgjY7BC4iTRxvdRfXbKWXpHvIWsiQ3MO/Rr74TnLZ1NeVAFtWVQJ
uU12FJ3JtUuEUiwlnrJ04EIeVX4t8GkZxLhfclneTOx3gG9mNgcfSgGMG4fFYR93
Nb2+w0J+T/1t4Zf2Fl32U8S7j+lR5JTR0z6EKCyA7pfQwbtOx+R86A5gMRPHks4L
M72E9FB7gYqPyrlmr9MQyZATFHvTp3EgrGYLwEwJ11Nw7B7pNKBLOZIG7v3JPeGZ
eJKBLfLO0dpaLNvPUjOf/XPq3HOFRHsirASxyxyMrjI/sG2NnpBg9l4TFJ/q7Yrw
Kc5qmSj4ouRdtqtVysS2P8seDbk+odzN2MxTGvB828U1D8JaPOIcuypRDQi8rPRb
A5pwPZ5+QokTRftvjbG+6MbmZx6TYhNBcAGVL9V0tJUIBkdUFv/GOBkN492scIqa
e92sredpPsWyYIsfUAs4vnHljKgFATLab/+losFwNE4UUeEqjkzJcK+YxH2cDpZY
uG05pp0OYjzn82DKZhD9IKyOOKE1dJm8DFUPfipkPDPOTjDTHzuJxrOXotZph/K0
Ihqy/XibjQXUsukIeXCfYjizgTRR7OyaRd6RrHn6+HBEI7PwzMg7/I19tUT3tdgj
//JrBSKQQy1zV0SXRq7efSCkn0eoW3jPekZK2ctCDyPLcTxt9Od9uECiW3xpcCii
LGibqJJJ6i3HbCRh+jFDb6tbXbh5RGzVp1EzKNKdaXCZIHmjLzxgPthMobAoxNZ4
NO9mhUp/xt4+pQFdsUcP9K+cUaItMqdQoAF9uYYJQWaemQCftcUs+U+YarJ9ovJw
UgFk4K/gQBBHmxou5emFsdOUZJsdn7/UtJdhhX832YGeRpAzNRsKa7ctoxwaOZtN
6Z4hhJXFG1s67dZyTGrhycwisxhsEXjxuiUXifWJwnT+N9HT7FgOKopmUVxGVYg3
ye7JiZFHXyRMV5420XT10MvPiztclGL9ANxG2qXsEokdsBaVk9x6xWBKmr/HvEwH
NzNh26V6WWlOsRyP9Olav5EczZvhTkG0F53/IBqOZihjNUhZJ+m5z64+azhQomy/
pzXAJaJkyIyd9Agsiks1EA349w2sfqWgklpDrHSP8fAcDu106EBCMHKJMD6gUJex
zpC7al8OlJYmi2F+YDZVAeu/SjH8FHevYSljPiMQKNX5s9aTQb8bUSmSKFPShjMX
ZcF3phOw0ntT+Jk+a2XtOa9ik4/CDb05VGPP6Fi+4jEQXJ2CmeumIqVbaHHNLDX5
xuUW5+szw+0MYLJdG1uPLNgFqcligTQU3oZJEHTHO/o8OGJaDssTxzAHnILwTElk
6vL1l9xQKPnZeybT92HFWjhW3BWZ5TOCDqGr8Fo4p9fkhbyHKKzNrN+3Fwv7hXqe
yusIAbuOsdXRWZbPpwWswNppL3Qy0UAKeOUhZejUDF1YwL74dUe6XinGEB5Puxl1
0wiroLRfcTl6GqKn2sY2gafrTKL1pzOFth9uNM9bdOC0zAw1rzJcV6dNzZK1rT1o
UJQpsYQw45bJyYpW993dnShX3o3TfFFhd3juY30wzeB4btJc/s6GfOiPMvAJBZ5C
14aHgTJD8A1BIjNOf8ylcRLOLL5V/krJpJRoGKBrmKgNOTmZBeP1+1JG61WjXdnJ
COrxIhz9IizroOF84x+XnA9HlkL5ip3m4ei1Gw1pa9dGPTKKdJQrgmeJ8b6ZGKc+
NuW0EL6fQSmyCtsoVqusOMacL2OmKBj5JEvQNWzm/sXK6e8k6A9+e2ZhM0TzsrdC
VHcbufddjDfmEtFYnrCiLSUKJiCoORCUq3rDgx95oOvhz5cFJRsh7dj84nNRB0Dx
yceKFavBgOItfHzPxtJgBOeqcCVne732go+5I/UtnVyp4pgrXg/uqTEFcxb3y69B
L9SVdTSpfcL7O9rFC5Zh3d6SJjhp+pju5S+lUIbtjtaVOCVKCBgzvAOeQKvCPyER
6v4LMCveB905Uck/+AW5ZLaTu+2ZGOONXP5NE8NE5Q9n89X1OwTOdIp/5E+MIS31
MA9aBCy4s3OCmlDwAZeEtw7WoriOpJ99OiflHi/L62irhYppym9BToWVkAvD63Ak
DHwKfurBvpczItA6vrKr2lo3BrNQV6+wBOZf8S2T69La3Spp2/Ml2XZKqh9yZsTN
0VifMRw8YWM07/rM3++ttCLEhyZk57a99425t6RPwYp/xpNisQEMrXtq6CcLm8V0
lIozVAYzlbiu4+++w2PZkVgFHIK20G9PJpLXfzBi96hPsx5snDUslLW1qy7n15dP
TlK2tQcGiFXXvZCkrvKm+0oAoCYrAkEhtA0N6yUJwI7gna2GFD4Q3FR36Icgp/dW
DPTA+9NYhDjmA08o+A2WTp9GDJZI+zM6tJmKk5lvUJVn1EyVNQb1hSqbDSJ8qxVX
K4IBbHovFzgjWx6fwGr9307Wojh7Oxt+l9x8hjRprEdqyVkNgUFqcRU6YayWXMx8
wwuOMMKU1T2TSpNTFVCtmJ7Vy7kFMc3aeVyo8qC1X44JW0bX04zdxZIyY7eyzJBq
Wq1z1jV3mp8VNeHfqZC1HQrg+sKaY6Q82qBx3iR+2H0yhZDbs2NmSjvUpu1XsB7/
nBTrBouGsFZJE39/UrTeyu44ZxU8qFom6zDR1cumjlHVsCIj6NEBMqStGXfIAfSO
YYT/1gHCuLYGOdGTsxsNqqNpV0IS5RL9dNl8lfkKPq4WqjnRnYbWCjT6t8GYN2Pf
bH21n7TOa77vk7GwoYaslC6SjNQpckpV5iasLmly6XQWwJ0eZPwO/UCy6GE10sD+
HolAz9e/3iTRHRZPBgUj/rTvOLeeobVWdnvAbysAhvv7knl/vbnOSC4k8COg5gpA
nzdE+6y7hgMqr4YYRbn/BT8xCXbNr3AwQc38vMLnVp2wte5tFySO3IuKCu33qkcl
mlD5Ryzy3mtuKzpowCBLUw8ML7HL2JT2xybZdlIBd2Xqc65HGeyTPHatdLf5L2oY
LtCn28qkVzrKhoMN0I9+nE4M4wrg7I1Gi6U/GVGFSDpOzBSWeH1Fce1/5AYcnQjU
aJNAHcgCh/GiSc0NUvZbO2pbzzc24wgNjHxs1kcTKgka5PdYKMXkjY4PCGNaFk5f
YXNgDp+JOoG9edNQkXvPhYDj0ijlkjmbEXDyui9CjccvxXwpMXlmeRneqmMibUfu
pindB2cg7utw/kwiXOzdN8oZOEBLoNGBR//vMSV22Z/tbkJvXCT6FicmGXH8rThJ
fKOQLGcCjiRPtF8hvM4n0/DrlWdvQbrt0H4IAEkDD6VEFoCTKmIs/t2gtiiliW8L
6/pkoUWRLV1zLMdBro17CputhxMclOvy4l2HDH8D5sXislpx3tkf2AIumVhL9ZFQ
sWyqbm2XCDURSciX0f1V9+dj4BA9F57rnHZfkNE2yQSR00v1orGJDzlqRNybEjyC
PsAfvI8126X0Az7SmZkozMMTO9xSDC0fF593sXnzLw2A7rbQD8GvFFTbSJh9wfmU
OhV+pfYKKEz3fGBoFEcOctCRRfpfo+RnDuYrHHM9rsm1i+6X0wOV1PQj1EIVhrmE
/NTBG3qp4/WaQmAJM0IarGXKbSYUGllo6c79C2ojp2NMte/N1hG7XUobK5dtjFXE
dX44uwyBDUNVkiFT65XTNDUju+BWjI3vYSk5fy3wMZx6Ut4yvzkR867TY3whakKL
bAlnuaTFUrUDiz9AC4/tJ/3aQcN3CtxkLp9iJ3Jwj4o8mRdzmXZu7OcMLngHMkUe
eBcnNCOznSUhjNi33GA2jsEW/X6nkWguF/9JqPgh9+G9cexzlYxkhM0xWyLH0wvi
6Ag7Uob/flDRmW0pBkji2NpRrrJ8Sykv5gvXy9nCbV1kF1vLsKOdR9+Mnda5Hxd1
Ki7ksMcradxFhBnCxZIw+HO6pgDPUYy4e3WkFvoa86zX/7COSzygrO9yrUFVDh7l
71BlDehTNok6q4qLWwrDaDhJGeej5npbSEGCZVQ3G95JBMwtxQSfADN76t5cp6Qq
ksWLtkFA49rnrAHNGkSLE3AXSR9vrMLBCgfcptnHPrNdBJw51xSOjNO3elU4CqvL
m+q0H7u7aR1lHflr1E3RQvXTdoH/rRo/FbLO8MMYS0fJc09WFSJ92DIxHHC/DcCk
5FLKhhtlpTcwbXEz/pSKngKayN1nAQOfrP9i0eDhMu4=
`protect END_PROTECTED
