`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uL4C5hQId3/633gX6BpPbkqEdxKTkPbPSEfkzZ9/ue4q0Sa0BFd6iIBcj/V2JMiB
zEN9gU2MSYHP77nZLpbH9MB1jITUSDctlb4Rrl50LQq/9So3X8LMOf6n44VL9unL
Mlh7FLvI6BiU5j7qWYE7lhEjU7hZuBlq/jymQ4GmYAdZOl5kR7L5Z5tOwVJLimgx
RHXwijczNow1anxfCu8isz/MBVXs/aX+I1eFBx4QGwa30ryXB4GyWSlzbDczaVR2
Ar/mptF7gJOcURCsRSZhrM5g+KuZv88AgKqmkNjZ1G8P+qVLb+fgDNvzfnF844D8
m5d+XjoUa7x24rVaZ6CqmDR0pDPsgXIJM4gZYHkJobrotrtqAZQBweubUqvCN1Nl
KuFLpFuXi+YgUz9ElvgdaCUtdU8yPI2euzoTcGz18uyQTF/57DkHx88r7PEuG5jR
amn90KorEwO5aaNfhEOHS2dLO5uLhf7teDpqLsoLWRTyiHCMANDFnIrBg5Xch76y
JBqk+VjBMjhEU1BkJt4TVukyPEbUju8HezxTj3+ZXMlw3YngOITgzii7b8PryazN
RS9Ol5bDOp5pgOIPTmZYmE76nEYr9+PMuDCmPD/UekiXkm7+L8SRABAlrmu9eDf9
JTEz/M0M2HRbBp3zkWF3uQUBpTI6nfvFVUjxMSEnmrEbIP9nJiUqy2i8IM0+qfnR
ZTJ3K3D9EWKPoqC3Z+uiVz2dBWJCapM8NR2BXS10fi/QIt+MwSLGIhZEPyIpPNFW
/VhMPqtJCTNdZviwc99yECBLOuhs/uM6eJOPK3EsgPSeHPoW1xKqYCTZ4qEJq7L8
YQsfDS6PoXVBx04vMNPp0Apf8+KltUPjz7Iv58q+p3y8Mi9su6D9gAuvmpcoqK0d
r6vGMNSVNXRQnlmwbv7Llg==
`protect END_PROTECTED
