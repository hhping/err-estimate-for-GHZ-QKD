`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5BOQlCd9YrDE8mrvvHmfAs2F4PI+HkeXSkDVa0cbL00JVw9PXSdr7GToeur9LiV
0VZNIrf20Fwbo2ym4Q4L5ANBB1Hvh/eznQyUqmnf/DzIPGxv3C1R88fas1ZsJAxd
AeHb4ByoghiBeepPE2z+xEYj85Kqyp4ZoQwrqT83kBAgXZvguFpXYlVxfhCWpjtG
lo8ZujhBu96xJpJcljM2BoH4OrNfg4CK6CzIeV87z9NqszLx26sziA4o9s+DwnG2
9xrnnwq+sXzNFbmpwEFwYls/SQijsDGG/Qzf6Vsuv8e9nTgV+hqMfQOY+kikM4s9
rqwWm+wpHGoWxum4M1go4vWkT9axszkZztg3lT3ABAn4xe26oFsDKYIh8J0pWAMs
2rhVO55wk1ZMoPzJFBlF/jJUQrlFE8m1mZE4PyicBOulsew4/OLzsFepbZe9mcz6
TTFYSgyshES7TPnShJFu6S8ypGsrarMr41y2bZAg3fNoZ5ED2UhqI2yenIu8/fKz
yVcme1y9XnbV94JEX48SaYC5ORbgBZ1Aj2CwWnDJSWn1LICEtxJ47flEtZ1Jzpd3
Isf1+67UnyAxJZt53JTMs/j1zBruVqAy9qbiUIIU0NiL9c6LwdQ/58cX+4pw/iDL
cS0WrF750FivR+vW+DgUD/NdC7ZVhAxXEbdmDXw5YEwmqj2zARK3m48YWgBLhaJl
PO4MTraA2uPcZZMYEGBstlOGhNVVx87feYvY3jh14n69Uij5IPTDDVTe2LcDjy+M
vjILBwdJ1DtuTL8DhhAsaYnjvjSZKMvCq5Iw7O980ffsQe7mTCtv1mMW27SI+XqC
Qw7PiykycyVb652Qwkn+ShDCKNtbaltH6nG2Kvcb8Cv3fx8yu4ezlRVoy3XbnB9C
nLYkb2pNVc7NPmUkykq5d25ipDjWX4rwKxgTWwhdWQa1GzYWmF5IXoX1uJFyDOib
GcQSOaNcx0OBy2X2JD2TyWOt/0jjfDt5FZEUwAkqPWn9GHoc/v/63p44KQDtMT6i
2ThpfJ0u17Niarp/eY2AaBRsIejK3636dpV79OaEKW3v7SNukJrz4o1qwdNw2Mmq
SE2GLiuLO03XSPQm6iIHAJmqB4xHHcSZq+5v44+r0J8Pr34iI5jbF6anrXWamNmT
kzEt7qtNLQO0N18o9/YT69bBUQsnq3UZPH2wp3SCcoUAZ7nGmoBourQIbgydM9/T
k/3j0UtxJs9gBMbhq5gtExlzCfYuEtEjORS2aONlGD1eWf1HZ4uZ52m8qEG1k8dV
8qTY9bcRL7kJ+bu/JyCSscKEOyS7XMFIQa/1q7Olp1XVG7UnFI8GDfwn2ClWt5hL
Is/oqm6KNB37ijR88vYTGLtL210LErm2WPJCERqRyDsZUAA9b3JmpOCMqTZnQkFI
IHmsPhfnR2PQQXSlBmaQ9njmQvkLgB6IPywv9MG3NcHmcsNXxgQJ1J99tMT0dKi/
dziyC67q03cHUItc2efWMiIbJNkLqQd0AxdWWG6yVvBRcFRSrFhgJrimbSNygu8F
+C8mjjmC2LXAzkVa/i4JGn7gL5rw3AFeYTmFuyR7HFRi1/weBfPG4S555Or62bZn
aRnvFb0iPM66pDv0GfvrYhqIiDRloxMsf4Ax6Zd5QsgihVZGnq217eaSJTIAcob1
8AZap7UF8H2XyTjJ/t3NnDGJQYfYWvfBrZfVh+/q6nOuJK0EcrZwyb3U0++Nz4bc
pE+bmdc5ILfYpzptMTg40FvKvGMtqy/6pyQ03xhqYdh1Zeub2pmxRufW3g5ps51D
0jNwpJZxaPeQ9NyH28RQpQv6pjmJOPOny+G2bNRG5inUbvIcrL+MEGgJR71LG+2P
bVKopI9wp1kSysfg75MVI+YHVVxPJnMa9bSYnMYNpFYKCRTsANsWlJ4+GaLue902
swukYiL1q7IdBcCEHorQH0fz5b5oHe2UJZfRjOyDmBfIrq4KFAyNsxssnVJyiBY8
elqtBxudQe4tK51TXWMOgAGYe6r3P5uvoaGdcweqeawIqK+98b0dh2uSXvm0GAIv
YyBL+bJMoUpkucHnayVBPTHBHpLFnN4WDdaHbMtdhDYzz7lIr+npU/WJpvJVfGBs
poRuu7QaFwe3snS98IPcNTF0RtuEPCA/bZoJ3pNqDSwB0IIcRTFdRR7itC6SLVlo
NkVfSTZct02XX1qICdH3wvLQhJrtUlsMUwsky1ksNj0+kk9SViHMpa5T5N0vEOm6
JAhH98TmQvtqIoqCwP2INwZmubOw6gOGOu5ff0kUacVcD43NbXaPy1H0CMxSXJRM
TeuWYCo9am3LfRUy/AVtr/rw507F3aqPoDjmf5Yh23lfF0RRhKG9sGvykey+QAsz
jEmxC6ACWdcG6XDZ3qbcFaFhmkq/AZfSKqND79re45Huajf6q3k83masR/OBqRcc
289wRHiN+VB8V2njRPCRekH+RQYU6lPCE1vR3+Y9OZFjyfZacjALqEg9+Jyn1ozg
awVblGIO36uYQ4sdNJjBikug8D0MgbtqQLP/QrBdCFj37YzVVp4UeyCIUFl7Tndk
/oOIfZoucQVnuV1iL2UDnlS+70dl/Dl+xASnQMFvCK58x2Nswsc0TPiY6HkXfEWz
AOyrSw1+Hxv0EDhx8DFpnaMQVD4fk0/RL92Bk4g9DozV/Znz/udWe2wVtPMqt8D+
7Ni8F06dpxenin4FpVHdNRLCavaZuDcXQmSSbSvBkisdVo36OZxiSQa+RysDxsiQ
5hfCRrqhxNi+lDg+PPUQB4o/QphTGprMS4A72oA+WTU2KzqTSZUuC9MBjBdKKwff
/xDHCs93z6sIWzflVMVwYziPoim+4T9dzBgafxq87L5tOtAK8MXY6uIPVx7Q52c6
TuuCmBhq3TBeQ8TXRTheHpC7RtshaT3ARZRXmds55OQxNDHw0jo7mHWeA0j5dDAv
vYiGnQf6Xk/x+ycjwWGsrRE4R33par1dqjngVWCCIsdLqQxybf6ZHrxcdC+fV38b
95wNRZvdoLu+kQ/pO2cOii5rJP6gkPRk/2kni5V3v8AIn9/u9ejOkZVchgCwXw6V
r7HJ2AnM/vEjL/Os/9zBE3HtoFFkudHsLtxezGWcZUXgsApAbNrivnDq/Hcu9wWD
ZL0x1oy9rNrhlzN6eg48UOTGMChSupHKjPiZHMU3I8bSLyv9phwDzu6+je2r5WGf
FnR6y+hUFBiZtDb+x1bk0dBfAzIMQICcKCQT5Hj+ESjwT46fdElULnF0FJh5+OR/
1yv90NJIzEcXjBXsjxTUUk5AEFGyk2u8pmc5vUhlIq5cB/2ZCtUaZxjstCwp4V74
WXLv0DEAza4TVaCHAgIfgGXGaMQJLYTFU/DVq7mys99Y5lL4iRYH2eq6UMnlgTQh
yAMe+yMZ+6Ebs9rd010J9z3ciR69eRT0aS1TI3qpn2y9bqMDZY1HRCjnpgG3NjBO
DwSxlu6CWTYRlZXJxojjTW0Pw3kUuLQfX6j1agavN5Y85c5syZLsmj+ECF5plJwQ
C1KiC5RaH9ukI2wgvxzviD7KwciD8U14EUnbEoiOvJTI1IpNYHsvHOTPulVGf99j
1/5CT5nTAl9OueQ84o/RNVV7HUHm2q3kO190/zaBmnh9qFzY1bsY5aDumkvqVPhK
GFjaWe5dlXIoPYWYugUjA3rCmvOjf1oBs0uCnC7+vCLMMuiq1UZi4BiPxbhRbhs1
dKpvFl5thJsRPlMkWtXi6cjYNRV8g/Hn1NrULX+ZKUz2bFx1BjA61ByLR72++rjo
LN5+uQuNfrA/exB58tdOnb8hb6SNysdF9NGOAepwUzPkKmwCuWFj9FLemQLo8pPO
mpAczO/CeW99+gB2YzfCAsocMoZsg4Fn99EtGrc/VQIpdY97MJtQOSWrN+EWSsrH
r1ezH8Qqq6whAhvaIPOaTsinbg8aKBa67xX0z9qPAW2e6HeIXXes3tpwu61eE/10
RxKaUbQ5ho//KBp3K7VLJI+xJi2oAK+S2QDQ4yjhhg2I8W/yA5IYYHCTwPMu8tfI
66Vfnas2yGJLLOHJ19lEq5a3rbvfEnvs6qcyLjz8yHqx/tuARm2D2Yv5ns1SqHBD
uD9j1USl2zEeTA/GD8Af2B31o2I5AMvO1IIPCJGyD2wGegL8JSeHMGzjbCy9qrYY
RVrtB8zBGike+xO3cOJXcy4/ge+XegJT5ZU5ozzKuaONGpobX6kzMuyq20N2FKtH
DDVwJ83z/kHhrs6O632CNoYa02KXmg/G+V266oforZTLPZviYIZYUhqAopSZVNr7
5sUEcyMLfvoUaFRt36D7Rntzv4FbNFTmcQLAz0ltfRmlkwTKgmIv/5bcYLnIw2cF
AqULyP5g7R5flKV96k7aL3TB9q8wLNIJR6NQnRywosL/2WsVJTRxmir+OaKl5odj
K5xyUN7s9INVGGnqw3oKuqRrIurjIVyrVkwsZqg6lJstjNvAvBhNbC+WVb122WEq
d8l46xom0PB4rZol7dakDo7KxEgvPL7TgtQiCGr6y+1FUMk660SGJoT7P1Pl3wPq
vkJ2DuaFZM3OiuqXJwrcS7JCenpOSwXuAOV5gz95eZf7UvW4XfJmQ8howzED6Jp5
6bPmYsSyam2UvnzBWvBP8g96ehdOCih2/7amEGd02CtKluATqddIKwy/qpsQgxKU
awGiiDWVBcJi9I6NkUb8L2Dr5Q4gWhhmi6QQxcjvI1wRxDBRM45FwUSR0gbWUWjk
TjREW+8QS8NES+LZUXuGu6EkUMWk9wSjFDVBp4FHpd94E+pC5oFkBIihFIcZYY65
dOX3VM42HoQJNClzOtMO4cOvQhEXNXAiJ66NROoHAMlg12Vhqcvzl7NVkzmgvB3r
PrAR6Y3io5T/dUYS+u2xNMCLXw49OAMTOLDTXTsKwk/ANBBASO6y/7lZEqh8aPIc
egPrRAw7Y/I0qPpzBJ46cXOxEQ4G0aKieffyjz8LZ4jIkgsBoFi6Wv3L2FT6yJu3
lafxl3XLmfB/UO9oOGECWBXbZeB1cwGXP5uF6ZQMDpxUrlKcG1XkmW8oty8TmzaM
DdqxlF0BhupzuygAq2hpMFZnxc4M4s0/SCpNmstjrfsEMQcbvcD2/cdUcir6uqe2
SD9TABxhUu/T6pN+U3TcagIoGWLwxqnjqCjBcxXTYLyWrE1tDOadPCftGtp5g3IU
bbKtTe5d3Ku7qPGjLTarTjgwVn3Vvl0nmUJ1BPEWCaLEyNBBaIbj3tMF9Ti+x37K
XXBF3kJzF20yYJnj3jvLC7Iteaj9CbWitCbqaDsCW8Q7zNCuCR2Z383WWzT3nfOI
hZ0+JmWmMVaKhZwQZBwuHdgR5O0O2Ju0UGMFQUMti0IY22PolqtWgvUEBoDMhj13
ADBf2cpN02FZZqpF/o4emTVCMuZb/vA3YuQ8UyhrZ1TpOx440BgOq9S/4pyeuWAT
vKchb6Dc4OlJS67Z584XTyqFG/NeAEkO8LZCT1rRBZxLT13b3VQ7hzisBp1M2hbs
KtK4/rBg0nzBVR4J/ILoCztZ29EiPhnp6AW2ExajrTqNNGwGtdvTRXAgxjAz2Cky
rPBKEfBvnaL1LvJGUT+8jkPLKPFogjquBktFKbPegMdlsFsD1/XzctVTCCI+Kdm9
gR3qDWwkAtg4tRf0BLroLEfFiW1xQpjNL16JM/C8J+lEN8PWI145B0vmuzvM9NFY
dTyBxrGa1JMUzIoHLtAsZGEJWB+SqCo4e6MFB9sadRBj6QGIoX/R/AIx4ijtNW4e
XF3dM4AOWvop78OJ35Fjkjn5NzXFEUFMyUnx3I9dCU967WqgagA7gbYNfLY/NvYA
iLTg5kuNpQzdUh6zC8+C9x7usTxSNBz7eLj0/gY6wJEPK0IjiJm821mOsdswpGzh
Mla53qf0lM1zTwfMlXXHgDM5kYuhYSQ0qPdBR3zgyEQEv0L4ykgFSacy3Bft0Qqo
wWj5o0dYOLAz88Qw6xPdFqvKGB3Yq9synPLDC5H7z9TdkpHb+R+xmYkj8lZ8h05t
2cAQyscUBIf2EvBHSWKrtcwCuOn8XZKDwN9U0OUOuu63Es6ORGPqIGO1p9vVfgid
TV88ERCohfEgKeIZQ/Fb+jQoa3neCUHzu0ENvfBD1iJisaCBx8uaN8MCQLxvIw1d
fSnqNM+BvAKg2jeNIytqWi9vhU8X5f/rCQsAq6S/xjsiJsa7IlWyRTJ+rPGiX537
895hkQjirrausvjSC8KO8Wyqvz8a0O2LEc4ddBXxNjVbP8VNF2dP0y1GSRS4I+lu
kMr9nXyYqMDpTru6DueWkXwcxakvJzpdoN/idIvExfU+N4VmouYfpjOHT45pW8zS
n1IIGnyC2bfemGIgY/qgI2b7aoKrXiWypwe0sRP2R4XzbmsaeZcVcbDoUaUiKb2I
EJdzn56aUYytaJAaw3U6VWRL757bWVfSscxtbtbDKUl+1Ak5aYsYDCj/xYXWBnDi
xTAXa2Or8M8m9ucStoSANqPI4F8Q5oto4/WFgZlwozDcOzfkNdtH4fPar6aMoXwF
NpLegB6xb0m5gCZnypQ/PUrdvAV3crjlnLXQq9xtvdO0dw5rRXrWV5DStrFjQmLQ
DT1LnqSrWx+PWOMgi/i8NTc2NcuRXvhpb4GyGMxu0Ri08WrAkBY4j2aZJajvOKIO
rzzRe9E/GQYulp6UT5J6nftMPSVOz02sKtO9a2RVxbvcrLSi4x4yiCiAIs4IR63Q
xHrfPw5OTxA4ThDBFLLzyVa/83hIvsiginLSpfqhy3L2KUsEEheDIAuLbgIdFFQ/
uDDQg0Y5fa+Y5Qg8QxtP9SsB1F8KS7+Y1dQB+PTULkLbtotoVdrsudSbaTL3RD9h
kJb1ARYCOALbjfUUMmNBThpz22Q/DbunPLP3QbJn/DF+R3k19lnZFPHFn5x7b3M0
2FReQxnKFStiG2N6AU9ml/q8+gbzkBU/9HUqWHRAh+79Uh1qaEi+jifJqu8cyu2x
bqWD6jrKCkXBQEzi0AyD5PoDECNxBYG0LYPtp5UNuE4LToqAJmjxTE96HcBfMR4c
0nj2BcwY89geyq/i2aXiLd9Z9BFtNZU+xOoO66GFrwRkxRF5+zt1a5Me9pnJQ33N
l4pWMbjEj2/nDfvxI4UpBejPqpU2DsJJfp0Voy/AODTECm9j3cgVUJq7XqhlWLZO
3IGRwS+MspAT1uEl0/1LQTI1spvJyNK1/yRv44a6zSCKM6OyTxTCqFhYkwr8/REH
qVVFIjF4UgaxcUrl16ZbVdKHjrcY9UxvVp6mxHM26EGx9NiQBFbRnoiESdy7ltJ7
bCuXRLBrGZRpZXKMQXUCkia3HNqwExnMG7VT8bLR9QukHsQXZW7uAiK+QUKS0K+A
YtDAC2w0uobaSTKK50H8j1uUzOwZh6zxGkRqpdi+35pzQYThDisv/cAaD0dG3yTr
K3SiDlwMG9dY/JeXsWu03xBVaT5v+gl424kk8Q/NFqd3Bvt6m8AM4/jowPJ5Z+oL
GADTx96YBuHWJOPFoK1lagXib+xDc4+YPEzHFpFJDrsS9adAPgfl5CGTbxMHKhAc
9x8zFcQSokFDHC+GXorekx4im4qFU8vILOcFsOMHOb4klL+sAdPTmUCWevy+NVRh
iNQolhn3r5VyoI+g++hfX3U/kErkeXyRzC/YNyrk0KWETkfZo89D7gi+VHfz+Y/e
c950cGiY62aRZEeOUlEuMbnzQeLlLbRWt/imSOA1TQXr4CXgGh8E7YBWkXXI6+a9
2LL26Ej6v+eqDSjJ4a5dHmdaPt1aPM5EMkKplq0AnLHdiMv036eTWmgXdNZDYnY5
PchSS0CJ9JGggLTHr8XuBCJ952y1DAs14CyTmtNlprkPPI4X2pFCt0KQFkHjVTnG
sIn17FxZkmrn1KE1E1IHxLHbEppbUAU7gpVtz4tY5KMMCw2x5Z1GG/C6k54d4nF3
WeYjWa0E6Owx2abwX48SJp+padcV15benX7gZIPNLIuOxVwPmh6ACxxw4JECXiT/
6XiHaJ5iicvR4MrwsPCZqq641K2ud//XLbx9tDAUP6hppO/wpiwxb+433BJRAxAz
BnMNXm5Ne0b0wzXyVcNOt6iJap2xIUNa19eNLm4CbnYEwP9Ue3iyrOuhzUV0T3Qr
XlzEfgy4fqsdY4vg8RY1g3LY4Cj4g9fO7cvi1x078FR5p+KxMbrx/o1gkBWMkKhU
MHBEpZTppmd4Gg8vmD0GSOBXedoUXZzPNe7KKvUrKlIxZ2IlwjQMc9WHOTvhn21I
OR+hQTDMiPsqj+zyz2UVb96CUHE2ueIw+w2xE1U4cKIFcnY+hPnUtm1vFRnUmWGf
2ZkAEL782ADpiEat0rj4MWlN8zDwZ9DvQaXc7J3YjMhFPP9HwKaR26LEpeK1COLs
Xjwx+5PnzeB9l0tO+SQmmC35Ar5/2ZdnLVhjFVa6OJq9227RpUiIDP5Vt/asO7kP
r2IX2P0czW79HcwHaOXkmN1cGEe586HorOMQjAmdQutJWfuqBH42vQ2k3gElhgmS
cbxxfCZ/PNKQdPBNb4iIbNNd2BegCHPPZ+dX7l0QLRdBD90tsYYuBA8IyI2l3F5N
xN9TwK6fZsmvxrd2BVSi/BpV0+qJ14ZtYBDYadb/dWbO5Hq30XDRO7ZydhStNcej
SROPyBkhyJWht3m+qKdhqQWAsDJYNGHy9Kt2sPXiK4uvupqGveT+ptneTVN+Bjmr
qN8+H+q4AMip6nhxjGyxKF7EH2Y05Qs2EgqO4/tL0UOyVTH1qBLborQkOhuMJUO0
xrFOfdosfejxQ9KHuq1bKtC7b2cLJjsg29krSNXmQqS6Gie0FSq4TeHhE2AOP8Ng
`protect END_PROTECTED
