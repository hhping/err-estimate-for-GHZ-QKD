`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8DPmv1dSIBZiav2Rfi/rXDRIn4XeetHH7G9a0uAVakW7pCWPFjB2iaoCQJJVamb
r0AqzkV2dsNZJAp13bZq9Q0I+y49soGw25sWvuxUCTxAYQGPrdvI/Y2i1GiawXFP
V2i2et7N+MWGDfAF572B0GsqFRbrdArH2dwqFF8AGH0=
`protect END_PROTECTED
