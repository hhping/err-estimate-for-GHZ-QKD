`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S8q/smQg/xoYt3qoRnmeDa6TiUeg/llzAr+7Gb7XHPluR78ZVtwC+6RMGwd5rGgw
IKo03jDEAIoXi4zslZEQKgCk4Xb27RcZqvQ7/vQlQI2AuZaGbGw4es+hhcGZr1Kp
0mHN7k10ej72TdU6jknfGtMkvRMznOLxTBkoohredKxe8ekj3L4/DIM2pt2+0221
3vEp5tgpKaaqMyZVFfh8R0+luhL6bscjCcYWjq04LubSordwFIEBuzFTlS8xYYs5
sbWAASlxOphLgUzNcEf225/JjAtNwEJ1/wIvyqYO4dRjZ3OaNXc8cX76NDwy/Gfa
+fNkXcfZfFk1oQ9AADRdHc1ass51hmTu8GlYuj3utWb6/YoW1sGuZHW1I0VtFODE
Sjn2oc3Lu8QJ+yR6WNgk3QynyX8A6Jnd0ooU9Yfi56pjk9y3dzeI380GWzDj21qg
gsgineCVCSc2f4+7u5uRa5c9RBxnOfyOkVq5EHwa+i2yupGDocAT2srbZj0qU32I
YwH8Oe3Frp3Y+Q+BzabGLlZ/T6uXWeymhr3w2AdnFwlEu+ZsV9XL1wKX7TLeo5B6
j8vdpcQ3UjTKBlUmlaINBvQWg1X1EooHaEq10wUzb5WXuUMGjHprD8Ugiggj6btI
vhAdlLHXVAplhdBEd4RfFOOlFMF9lczVHJbzp1FHAfOodSgRyKs7e8uOGCGXHia4
EeA8MRgzthV1P3BEwz4o1KN+AUfOuvDovk1kn7PTXqBetAYcZMPgG09oWwH5DfQd
tk2Z/feYDht7WP5FEEF0U/wxEfJvjQ9qPDyI+6gQuMmZaVMh6kPhggpK2spO7fNn
mvYBpVZfSB1UYdbaWbaYHpYqyQG3lr2/8VlCzGcXUhhT1q7V88yVvW4ax/L0XTW/
t9r5wddC8dFfArmo52H3eI/Cu2eZKWfY0dQisq/0GeEWKevIu6hVnTjCxYXm/6Ft
ZAfcsNU6Y2M4zgetpy5U9Y7YTM7EFqK5wPNymbFUg2MpLP4xa0tBoAP/76ronFYE
OxrGEPsY7xTnLA2VUJJv29jUAMTOFTbR57hQA3v1J5oeX6ku2Pycc4kSIsNaUHso
8SujuCn0MxklDExbIodT70wUbKd9DnFuGtS+9Gn2/W4Jsp+ds8K+IY0B7TN/9rXu
qfAQ4Hezp2FwDiyoPQImgQ97aFNjrLVyr3AEg6IwFUDA0E6Hr/XaoLlybUmY2h38
+2e2alYi6bgW57vRmGnyNFN6srzZxf6VKrF5c/Ut9n4rXnKyKvu235hz3FrKK6tM
bKIxmO1H0nFsS79svN7HXPLR0EZyK0PXzxZJL+1vzb1XT33CEG2ijkRag4QlD3Mr
BEyG5XNFgB0HHK53pzvkPQzvqJmesLK3B8hiUpHg4ifE20MRyu47RjeNBv+Du5rj
03HRd5iRDMnlPxx1umuofsqTrZSOU4q7Z3D616c9+olvZIHSiZnMzCcgXK/w08yv
b+rxhSEB+TNT8p0HDhkX2whORkFCyGnPG1VwhQSbTNV7qTxzqcOGkD+eWYMJb21x
Ba8nsw9yqpAbVrwNkReuUHxvkcoXTnzDm4Kgi3dOJyw3/tEP6dxxryIQz+nJnAHd
o7n4DTwkSRsLTOwDSZhrSAzSXjFI6alMzq9tHdyYitu2DzSPPER9Q/Lq515RFvG/
8NtylF+bUWN1gWdqcb69bPFIBnd2BBfB6hmDfgIeugGd7g1sKU1qNyYgs6IuRLp2
bvBL3JfWawBA3uysxoQmM3JwYQWOBqZE4JajDexetoimKVsxR+s/jegU68S2SHDq
vGtB8p17WSHRSZUmX8E4Frz8DLflCf3hVeCFkOoIMZoIB4CAA3mauN2o6SJC0OhD
XZQWMOa/ksxroW4zeac0lw==
`protect END_PROTECTED
