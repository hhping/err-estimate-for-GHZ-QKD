`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOd09UwwY1EA2r3tNWQOFC6hh9I+neeQ2mKcC2wwfF0OdM1u93W4rjNMaA7t3BYR
seUTc0+OJ0AMaZLP1v/Ed7anN8FVdJKeHrUhiN/uu3ra7L/PciZEfkn/bXSyOs9w
cHSN2AOUn2xVkAOl19qTd7R3491jXEZpjIT6tllEve2jMtwRnWl1JZ/qKpRJDXKL
Fte+Fu4lXKW8uGZ8IL6WPu36Q/3q2pPTtpmfFsl8iV7VzJg81doUZfkx84vVrqWY
O7WUJmhxrROxlb28WaNs+zrtbmFcdQdzX9EPska7UJMr9USRmkxybzfOdvfX0x3D
8k1RjHvweUcTfhjxMxZDUPkdMzwlWw1eZzJ/c+DkN/+oAvHopOp2QqWfJ9RlvoW3
zxGUrsdi5AhpkWQXNLXQRbEu+zV0CQhf0yutHjyKIZmHNehkTS7QBH1NtOIeNYvh
f1FFKy0opo8bjnC2SmiXqQS71uLcJDul46IA3KuPv3+sDX2xtQBFDBpjIzYQaZYP
GQbj36Zlqj6VkbzMWRZgRx3paiqFNqP9gza57Ipmz87q2MI9Cehz/cTwPUT34FY0
rrlXNX/S5EYZxM5TVxNttBckKim7pAuTX3eIQaryzJ6Av751QxZQtshfNOuLImmd
JGJqMQboyXY/9HUQg0W4wUj/fpIkZ/MreBgyBKGgNIiNQ5bPrlSXINXu4G4FW7Mz
dhawB24x/i/NwFqmelJgo3vzhgTzpwMZmlX5/7reWM2YcTryK48pHmmdOJFW8zgF
/IOGb0DX4w2czVqyhhDh6eLimNAE15ATivGyNtF1KRcCMI7kTFi8CNm2KKBNbWQH
cDPFk+IGy7tH02iQu3ELdstawyVEoLMy++2yr/ONrDcEjKlYwBp9jXVtwlIZODWD
baYl7Mv+90pL170Z+mL3gGIDOoAAYcz1pab0bvY9Np5JEkOWSa36w4C6y1Hzcpp9
N5E/w1EA9sR3chTJM/k54NofwrXa24clbUj8d4lfuBWuMXGTuawZKmeO0Wj6Te6T
p7l98btkypTLIt2k1LAJWXx8vAbnnAt5R6dBzAR9rjZPrzLW1NzNijE9fJlXzWnm
4hu+b9JqnukON5MZLhfUoP9Ned9ecYDRnahB+Pblfji7+VI/YqgJVaUrn0lwWrkt
fbKRvQE+C5ftV1UUvxaNWdFZ+eZdDsavxrE6Z5tBtlgiuBoLKOcI2Ut5aoLXr+I6
AYpNPnMjyZ9qrA8DHarvs91khkspRwfJLfW5e5GsNTrXA4PPFeIgEEEE9RoUC/+g
2fd8kstfYkdZRbi7gwuEpFwphdJuCBBrau+mzPa0kCOC5MU+Ytn9ODW7weP3irOy
GKdC/892Wuq36yn9g+P8trIlUOOq/itlfilPrHbjXR96dlqlDFMv+9Fk6QXzCDN1
4cDBwOXDyNVZIZWYoXzVpxPBE+eJo3a5ewZlA9qvCbBpywntKDODRM9x5/2iNb2z
KpDNJvrIm1x+vPbBz2zqcZhPPZGDfLi7JuqEEK8Z+fHoezpmBdDXfRaxVxwUiMZW
IJ4rwxGTO61BwHvk/CdGNzo1b36Q07zrMd3m9yHibYSTOXVDGusX8IgpM15PQbFd
rPHoGNnPfsJDDTa9UZlOHPQ6DlFCwApqpTprpRY3JpBVP1LgNKUjkjHig9PqBjJ6
FMOkG4wb1h/ZQxBp0Plp6oNVlHZGI6RkJ6Vxy4ji0xBKUHALx4Oz5B+FIOdRtJro
Go8sRpQAiaaHFQR0TfDu8FeJKvrz8+xidbshmXLd80gduoMpRxEaFcr6aJJ6T0oM
g/5v9y6cSHNRLmRz/r2NJpLXtjgqZxkLd0HL9P/icAuHUENgBPf/wYQB/PhubTFL
1RzZomZp6VQEbHGl9jDU8BoqahDxUpLvQBrHf1vnfFHqql0DlJyz5cue6ZDoThQj
FvwKGp6bAEE27f6uKfY93j7WlcDZpO488AMR/X3Hw4N7HezZY/tdJ27uZFuL5C5Q
9XXK0AhA9cNdQdzPBxhBhjuMeZjKE5LWSP06RJ6f7ERTuv7kJsA0Uws7wif6Wbqi
Pm8oCA2lwezF7YG+af2gOXpn6SnV/ITkvfhyi11l/9BTV+wRrQbCcU7MSqDBEdfd
VUcty0Xt8w+SgT3bL7H8jV5bcHb62kl1KmnG3FN5jw1DkT0HtQY6tUVvWFigMrNg
V1UCnKpG4PIZNUIi60/9sCDquwS/aWQZaey4IZ1D6JXaBToXw3lOVEDvonb6v/2o
y8Z8tc08uhqj97Gj9JcAXw1uYvXGVF9VTUipvpsDSbJtCDhBWEU2T2RDBkgrhwYx
0E0Fer3UDLXLN9RfWAz5xrxmH4rwwfUaunU3L1gziwETnpBdbw6kO1+doY2YAur3
TGUrasV3x1jignFJJqObmawxTrBY+UfITSPT1PiY4mIgrMsmTbCLmT3gKnWzytMS
AJ6OOK+Gly9brpw7Py9glbbJ+qudS83CVCoi+jMtwKq0wgDU4tqnSojTNW6Zeadt
QFCfNc9mo64qVx3tgdjXYg44c5eRQ867D4UKqCMULbepQgyZ7TLeQiY8VmShYAub
78juP6bEppBigURMEwPwpAP5hvpBDrLZCvymb6HLNOW0/qDtOXKdzvuXm4zFfsI8
YFxt/roIYyxlyQhbjoAiie1RRXm9dDvS/5DpmPCz1envCStylNqjdCIzibYC01Cy
vqFEm86AA2F3Ib5OzIHpbAX+TM3ituiYKpDX03oI/MXhXQWDrg78p7SB1K2bedp0
sil7yM+0c4uL6pBwl1b5PZUgdZ5c7z1T4YIJJ3j4UYGaEzqWHUbzz436f4eMhgO9
+YqNrtaPHQqJzMw8AWDtOTPPFmsf+yp1rLMF/xsxBPLmU7yEp+ZW4FnEqcv77146
1BdG3GqODaPKdsk9jehq8tZLSqc4WuS7M0XKDyFvx8CBczvMMOArKMMK4NSy2KAY
FXXPdLYNA28Xv079kSjU+kxG5mt2YNOlFA7auCpNiCOsjz17KFL8eSjidsArfato
Ls8Jh7OBKGPvMmaFChQe7qhbxQOvSGmVgmBvt4IPeObyyOfCpYdHFk7HS3RkJV3c
YCpAJaGslBYOOhkKmLtZewl15fvcLTiz7BfZU24S9Ydym3WvdSkoRg4eo8NDRKIS
Dtcn54YeYFkhGGgCNnbdGkbu2QNF5y8GWUuZMeIUu/QMhxskKRBld9TGKyHbTCNS
uiukVkPmBE3CI5AB2wyTC9paf5RBs8a46ee5c7F1XyixPzEoiIonP/1gaf/qpvwM
+8P3y3C0CsNYlN3pTR9ILNvdsk/KO7xkoYPMMQSL6rpXdezEPLdhkJrC77Kn2dcq
3olnaFhGUZVN+/MmCADPtP6KAiPEc++hgNiRjWs8YDac56zEZZSmtQlC90yfvIap
b/+2BH7l/h++WEUFri2dzYCP78rEm3qmEuZIFD98fdFgnufNCRHqGKctnoohqzbU
weOidRDiC/kQ4kHzri3SJQO7dh84SmgM0LAHDUBLEWX0G/IA3tYwzniZv4XmCdQP
ZOEEluxEn9zXxYbDpi6kmuNjSNV274ITuCxQL2CBBnAonpXaA9a7JbR8XwLwjpSt
yshnLQf/Iw84YIKAjVuPsmg+3j4fUDxzK3U4nbTAM2yH6mJ8kaYUePCUDBn06D6K
Ebs0HlhvjMCRgxL0sD5J+7/7fdcO+M1P1TGRdTFn/+mwuFbGY48k+qhAxMlQUki7
xSHL+2V8rnSUvw3g6a/CytzIAi/mvgO4VUZjUJS8SvBBFzeksQskRLINHW+zjdWa
Tb6LA15aYJew0lLJt26AlT3YN53jOY4uBd/d39hmhKbF8KFOHQhyXOUsR6ybSrnG
XSC+knn4oXzhkXU3qvi6lFQD9IQxNSon8nM1nbajoVD9Yt2Fw/PRexSg04GRHFey
GhajrSIplYdaTt5DZI/Dy81VSJyWMbSd7lkG+XDAgpqs4/TN9d4IsEyFIW99JwxC
eHpCpMgOgUZBWrUtPg2t9hjyeDpZB98dqY5zNGYxnnfUkqf+/n6T/USpuiCoIO/6
DUgVcARfOLq7xbqFkMvaPAHvBOINgeuiaVBIpnNqUWfDv4j9Z/rxKEENSaF6oBPq
`protect END_PROTECTED
