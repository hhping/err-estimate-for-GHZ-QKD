`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+kMEv0WDGQzNthwKX8Hq5i+A7ccOIckZfJ6iP77tNRt4ZJrr/Cz7IkopGzYv13ET
nNemjZrXrRn7NQEXF08xSEkvZXKW6degi4xoxLYASsfshtigRMwbWcp9fKsNajh/
OFfCyKP9nJGnfAtSfIeQcBvNTqPP5V7Za7TAlHgoOHEkAKOQaSgELVOF2EoDV/xW
GVXcIhR3TbZ76WtrubFJzMO4ICoejuFq1ggo5jhAYKqaQlDzPbeQd1TfANYTcOP9
JJxT3BO/mFEILLVH5/DyguYkp7fBG7oK9pHR5UVPpGFg6Bij5HzGEtjZhqI1Pt8m
jD7H6O0jaETtSAV4mkWsaS5oyAyY4Irv2XF0WYCr3cdT4yMuadYnaSStKUzg49lq
/N4mwjTCKgM3uYN4WAfr7taenat/L4J8J/0+X5bmlh3BItWfdYHFR95pHsF4IfC1
IwGzFTC4Sjjmbq4zgW3k/b/EGpZ1TILqw5jhop1tRuBeN/RJpuwdEY2161jniqBI
aeJvy4jqYz6dxjytapt/niWLDCgvPj7bs9oGYuL+7h3KevugY33ECInUVnQg266Z
ZvimjIHXIJomf42tNqbubNICTziRmCScsiKWkcf1AOMYone9lpsb4TYi8rm/SSIs
t0rN9UCD4P8ylaakujoYm0vXtm10HtmgArojgLCDD8g90maNwFhnsrSDJx2blcT/
arl5egAW1iymfhLpd60khBkiI+9b7BEEn80aQJUk7lZfgnERoV6q6Gjlee1npoO2
cDZNEUHSNECIh6DlcXd+lzJ2HzF/agevPlpsi1V9png7a9oEc5WVM00d9PFJDnMe
f6/fLdqHk0z3ESVWNJ0CLg==
`protect END_PROTECTED
