`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qk/IvKWtrs6cs9NxsoStof5izfKwc0D/nDn5nLLukVcMpeD7L1ZHJGn0wBteg59K
ksqU/AfeVJCTCxqQkE/i+gP0mBjgvzIYZwBFWU5jii3fYIyTon8cUbVqygQCiBTW
mWqUplKEmveUuH66EwHWlKu+o10X4/XFTdZCD5U9mO4c6tXizPQroXjpqiM7Ve2b
Wm8J6eMY+PTNdZ3yFNeuYxVI99VON7BZPMQ1PMDWurvoJrw4H4pwe1NsPkTKeIgd
aefi3j5BabDwmFaBrXNEyNEkr7Bm4V+lEa8UHCRmO3Z8lbUPRqw1RQ45HAAmSyOj
sfhS351q/9tFFsBRrCf4QNshUHZvFn+2vzaN+/gMrZNOce3a+7+xNJlSIMGVMnd1
ulmuRujRAbgi7qhzH7DpDsQy7tAsTIMeTcTyDcLcHv1zvrD7qjdFQoT2Uf34se9c
UuWEHNaZZTsCzk3K4nMHMkABaxZxjVbEkyHcWYletd+ZVhNkpER3g13LtfsV5A5s
lxVQkE9DSCjN0xgXKamNGEJSkydxaweAQQDz6JOX7DEG5KLT5FuDHxcTrDRkafo9
KQuROXDjBFEaR86U6kdQHiWOfAz4JzABT3r/vMFkuuMU0H4b5bEj9CgvaOmD6eEI
xedsJEXPZibkPzGg6mcExTnwrbb2zzhr3ukZbTNSO+IyOhUIwMuTvhR5uXxe6x4y
SfztWiQG+LBjhczg69Emo0GwZclwgLjdWq3wXz44dUA=
`protect END_PROTECTED
