`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/dBTM6cHUOycJoFL+HdfsiT1NhJHrfzZ4kSOVfhkO3WTfVL0SU62QCEa+3IH61m
daHI2ryFxQaI3/B/pv75BHdc/SwTvX/IG7U922Dbpha7e2Kpp5ncp7pIHNw5Ty2P
Y4Rw2jMG3FQSY57nbI145H2ijdZ4RrAj5UJL2Lro69aQCSEWKDLrueYKuoC3XvXZ
zFJv7jtoDk1RTviaOsclyLve6g8iW6sVfL3uHw6OUumGZJNBUd8zT//zOo92xlBU
kHGWaHXZTuy5sbuG5GiTyJRt/Pva7vk4dDoogEI5Tuve2hRZq6uUI6qMC1nbOwvh
gT3LVw5wU/pAF6XcGXsyhe0IuGgUJG9/4e5YsypV5dZu/ml+vgjvs1e2Lj20USOq
mlOhORGc46nloo6/Z4UiibdAyQOTqCwdMY0Kqwr7OVJKxqniqdmdFD68OYp7wgn3
XK9DucWWrZ3g5OtEv1Kn46a1LylCf/dGBJ6GpkBEmD/DcAb/1KPd6jumxLYZU1Cd
S7jSAgKeb1VSdtQ5GmJjx6lxyHdhzJsMCcgJGA80FlRFJ8Z5C0b0TXmxeKMJXWA9
ZZMQplz7WJcifxVk1vVh1cHYh2kMCXN1pvtRzva/LRgOXJLecvTJRW7XAYyMG7Qw
xZ5xC3eXKZRJOedRav6JBOsSg32/qR21JauX5NtHAhC5shlHrvIdQwS0Ikfu6546
zTeXrrDpNI6AYINnClglrlsodyRSgjCdWjuATMKDU7ikJu8qJ3KN4J2O9fnClQev
gFNIjRJLwLoZxeDZ+tfYb1D1bAXN2qJT0TwlRdg3B0DmJzBaCbJUJdwugqSMlbed
qPfphZxUSBwmZYAuwKWWBVLauLGmTp7BN2yGF1BYSQv5QkUZmOn2fBnKN61odNvv
SC2VDlAvyCKiUO1KbHwAEwZmBlKLirKvIPz8L15IJCwqnIqhncQEw4PNN8YTtggi
Uexc6Xv33stHvBS931AYkbhHnX+xXJg100PRbt5spf5IOmMLN7ABdni554Xs3kQG
kg0DPCSCg0sQuiLVbbSBkx8Cdii+6tybs4ZOH8Urb+AkRW9YADXR2742K7a9tHcj
qo5J2HsWTTzO+FVyQJWHddCyGkMy8H/zxkjl6hBvXRHcJY7jKpbQ3VBNolvLNAmc
fBdzL9oPd1hK9BYnRpazWAH9VIeaeMUXNjYqM+ouJRrAvAAt8WfpcuIUyZMqZq2j
xmziwQ4Ch3IwvTYXPpkYw0PY/pYnk/T7DMSIH3r7/Y46RRq0H4MKmQ48Wa7EQSIi
KBlrN9z85k2GxzJuimXYiQ==
`protect END_PROTECTED
