`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZm1G0xjTRLZxDfabhmlweR6V9RyxZ5/+eMsQnM1zON7wGRqPEr08zjguGXT6i42
UKl7+UvNNO/k0l4vqt+36DRNV9gUwAomPIaqJb+0iHal54KuOG62VnvehhRaZ8Hu
Q4gmqD9vvOAwtvZKymTjw9fcJv2DMx7xjMOj6ltDQAdkRmqogVG2npbq7c9A4e5X
mWGNf0ADtaBPmZ1fvdKx/8UvUTLjjo0zktP7zt++XGpNUhdCgY1eCKZS335Aadib
XcX54PANB5wHM2ff+CzB+Xra+jTvtBmf+HK3MB+Kqjvi0TcYSPPdE1onMQkiSBj/
NllR91kLq/PDErmB5ArkT25gXfFmjM8/uVWc8Z1DlNI8FCJD1JHYOyXoWX5rQjAa
6osbpX9+mCYPVbcXg6p0jiQhWVh796IzML7Cjq7alH2ahHQI5pZpLhTL0nSft01c
mfHzOz1MXeixMTQ0OvUvJZww0unoJtbkv9frwfcqkV7jhsN+q5yXigNRYHBhb4ba
MRE0PYyQfpMv0ieubk1nNlmkq+Rpiof7P1z5dW7ijNM=
`protect END_PROTECTED
