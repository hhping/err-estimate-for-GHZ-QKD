`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iSoWF/yiueyQjjnlTU20Q8XZuo6PLjfHp5nydtrOjYKpvUf1I0/WFILVuv1hJ33W
Vf3Zq3EwSeeSg+jGDTIEm+uymeuh4qwTmSBHf5O/zen75C28OtbxFMO9e0i+GL9U
0oM93mIZvHR72ZzQ6onXOotyZeve0dVmq4u6JTXVQSxB59YxDLLv+1r8j51soZfo
74foAxykQYd+GXpwEskBcAUmalstgtd/s9i7QT2MOSSG/omf5Wmt86qFwQuczUYQ
g0726sNeI3U57ObunhbxT/MR80MkNrn3U00hWECAZYh2e4fH61befPlTcZaF+bmv
F+xwTQZH2psTC5w91sYrIi/BL+TqKC3hkPavRLF9cfRe0KQJYoAZYmFzLzaBEEOx
a6Skah7GH651QJ7lds0yCzpoLOJVHrxKA865l1ATxe1GJLvjaCVkffaY6N4KYCuk
LEFNOiNDaLPk5i2YPjhH7/hcbFLMVVmXQ9gD14cBYOT7tTvTt4J0oFHcnK+2eoVH
3TJk5dobKGqh0hu3haPjUPy4eQ5ixO5C8ve/B166k74=
`protect END_PROTECTED
