`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scGjv63DbW+ovfsTtk6q7CgYrUNVFWQYGYXXG6AkxyCqUboXNAQn9/8ZUO4Imivp
GgoEoPkpke8Ecb5U77Lrcl53Tz9mlmEdUbJNRYzjfE4TGKeqrmtop4wnNCQJRzIJ
G7DyUHQ/usp1ouKwyqKixhxPSF/RT3aoJsGob4w1AIOqwWLp/GPD3c9PKx8lB2qf
eopsxB7k3lzuTy+7WebhvthnoSRG1lnoNDTRdDtrtQ9VodKRVr6/ExnsKHt5Pzce
dJ8hLpZZpq6YdioiHwRhZSpvBukwPabSQ8OrZ5XoA1Dr2Ok2kVqs+bQkClKMPHTX
EvWIBzC8nZTXyld6zAsFkX/LS4TQjbC3i2I8UWxlrjFlpGk0iUbbEZ+FhG42IZwe
7wTaXqPjqN3Yv5MXwI0xb7ddq0LnX0fqSTsqe59I/WOs1/5KLqFv7d7lY03pv5jh
PgYewgviLB/NhIXtL0U9cpVkCDiBt+y13NKlVDEH0/9/uUctjhKwKleDxY6+7jZC
+6sZKbM+HHsDe+7OHgqdZlzg4795nBNh6b6fhfygCE8D1Y7E20eM+NxilGqI/pra
6/Jce0pEoM6+wtRd+oSBPxIkz8b2LZFQmZ0hy/ay9uoOPjRz1RoR/LoGh3ef3U/h
OmnMRqxgKfL78WGiDp7RxQ==
`protect END_PROTECTED
