`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HKbG7vyH6V5Q1B12Dc/anwes5lmJEabCR4ayjr+lThxHnux0Hh+/afhz1W/Mcx7h
SIbMa7XG6f/scLsrWmtBZW6LoJoY6ja+SOIdUlczyiQk3qYkeBNO5hwfiuy1vEdw
28Gsvuhi1QoU0Z73WiMC24GAMI2U8gn38UuwqsBT2NBDLOQP7FUPL5cKdWgKkVKA
P6RfOAydcAQblVjjyV/hmPsFxipHfz3sIjmgwgjSnY/i/5bkXJBWYKZFv8sivypu
Rfh3vvDjH3TnXUd58BAqwc45AJLHNceECFgxP0j0pto3t3OWJ2nMtf4nuFqy6B4M
ORbFQGrUKM+mOv2g/zI1rRQ/VFYe+N4i8+nfkQvpk8CQloR2DsEsaRyYCC3EY2b4
hcBe4NYv4xVkRVoRF8Li4A8Jdf376hFkkJvG4h2dBeaEf+/VjTJjS67Xs6rxBHNW
7DVFvDRfiAxsu/CNTKwa8CqFJNgeEdwPR0K09c+NXQ8+a9BkMjMNBMAcuzQWVCVD
UCdSXUHdoA6nLEK9ZvbQKLxzvX+a0TVgHucEX1pP51iFFaS6JftjdWQxhOfIW+Fk
4t8nFEAqR4SAC71sReKoYwv0ZET3Op16y++Md7+j6yw=
`protect END_PROTECTED
