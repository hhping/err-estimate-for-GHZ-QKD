`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DiLIeOYOTMhDf8kxwUWjJcXz94jDz1g5AY9QTeZGY24DGrYUnjzTVr5RYvYeXzTJ
bn2+yQ+x9eXJRlaE8VBlASi7JjDDQKnDJGcTzXqBPPGSFzyYnSCPfrGN80y6Rzn/
KKysLnFFg5BJpmjsLlWKOQQ6n5q8SiAfj81Jm7RMB0NNXTbb+dbU7TWk0WC76W9j
glsyIXEP0yOTC3PMqIAbnKcYKM9Q4sqtXCHiMI1CDkZB9kQS8tAwWeaUjco+V3tN
36G44/pyKeo3kVRFUwpSO0uXBoMSfvIxxgC/kbXkGGCMufoM/RGUfd43uNAc3SwZ
QMlMgk26hsjh+ZBLiNtTJ6ZfYnFW9R2CjlkbChREbjOPdheT38ZOwgus1iwr1Ys0
Y8cyLcLLLiPLF1YULWHWAerqN2Pc6SGuoSLo2vrINbiG3sfCHJbPZ+MdTYOJsmHt
cph8fGYzlzlNRpwkuUo8Svu3ptr5dB2gJJv0wmjxICzgBxRTSh1BRV11D3kx2yHJ
fecl+YSJ8nGvSp2BnXx9m5ztZzsq9kNcbDLLao6IfwnNBVqWLMiAug8EBxyRip9/
OiUWZJx1Z33SPemHFlNYtSrA1fjQflwsKWogk1FON9JpYOEnHPyU/UNxH0InI7TC
ELKpuLKkUVEaSEzfnXvBlpwSmo2KMSAUXKMf7LrhZgC+NkC+KpYiLakQnfw5lvV1
YIAZVLCtlJMTosogBC8AnaLc5PphSajxw30AUPyHeaN6ZhkC5ZQeE1ES59B1J++H
s7zyqTBEPxVjAy8QLlDl2MzOl5nFp73LbhxyviPzdQ62f9sklRmG8G1CW0RnRgh9
WlQGCq1KPK5PoSeR40wquw==
`protect END_PROTECTED
