`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxZa4fKK4jmU9El7ZLohFgcQqVCaC14KFwIv223LORauE9NwqG0EZlyKxN0fFbZD
UubAntsE7oQwREIBOEC6Wx7iqsLk+2sn937RpP+ER5Ab6P3n2seypScti5Qt2NEz
6vSc6BGvJXWDz4DAzr74hsHK4ZJSs8aZ8AqcvnKGkOPH0iMlsGzH8pb16nJ1q9sU
S+ya+eUsbYqeO3iXKNvrQAjIMYjiTQBREXhzv785CiccdmKCZkAP12F9tHBmLP6q
tXnPVeFg0HsF08gI8KTJs9IPk7b7runHP9QAWRrHD1FmQrNwgeq08RoTAe9lVLR+
/xPqUe2jcz/bFuiCE7nqwXkGVRsZbVFSs3zCxnStGWs4dMADwv7iIyDP9Eq0R5jI
KtabMTqHmOk6a8duwr+QWFi0CzXLMOcKu7wVw54UZwMFC0RCNIcG1OL78Z0S77yG
GGziSE5rPbBWhhUKn2cp1w==
`protect END_PROTECTED
