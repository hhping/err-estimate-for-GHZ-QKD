`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5kmOs6X6+IEURiK9OZDlHQGiQ7LPoRQe6xrwLWMzLwnIwheg8wB1aMqTqE8lo4zd
RXiYk1Muf3cVMim0/ySgBXdJlTv2wXacez5UKcuBdKPWCwQyFsqMM1UB0ropuf7M
RqqtYHC8sVwZD8yJjfWrhQfwl0nZghVibZ0nJUnQXNw4l4vZgB+C13T/E94qci/H
scF46M1lUf4RNmA6AGIAFLwWxYDzgDoWhn/vs2BjcX8atK6NwPQGc0mL0GZCS+dR
YRl7WlbrSX5d2TFpuk3Z7dgtOCthPRtYs3RBXOLuhj5SxM6Y6Se+ZM+fB0WOmS6J
uVFdOFx8iidPInDOAEpBtTfkIIquOq/6gRw0m0DY4f/JxdRvvpWLprRFhAa+jWRd
OXzF/sW3ksoHLaVFuRZG43WMZ5nBO9p52fU3jAJm8H6BdXl+0KGrL+NiyYpIRo53
rICaL7n5mrHw8bWeC/2ykkV8+vJKIdBR9bYS1UcZj/M6Sxez1wM+O+itH2qMT9wj
uP/a5EN/ro52ftK/eo1knobB6ZahP3ZlI92kezVtuY9sJDOrkmDWusH7Xw2AZo/0
Bokqa0rBWAAuAR/fKd4nR8D8lvtECyVldoUYzMEaQexmtWFoRDGbjxaDclReYqYh
zz8n+p80/DMtTk3YJSkdmj7Tsrv3AP+UaxWXgJJTWeurPFtDeB+YPYNEF/ZzthN/
HFIYuJgBKUpmHDD6vThT9LrII/JvSf6Hna1KvvIvO8pjtcOd0qUUxAnoTtYJWu/E
dzhHiKRPI5pJoq2v4+bHkyeqRwoB08r4CFGQJTfqyWnETJcmOn1EE6CWcpuasGKP
InXooQZOF8uJyqhcOO+UPSzRcrSsB0rea/cxFhGQr/AdVit93NsEfUMKgU5p0Bjz
ii1unGg+ZCWIqowa1ODBDBzPxbiuCfBWIyp8sh3PyF8IuKBeFuRsJo3E6q7pvhkE
oiOX3uzgWvkgrt+Jfs9RWTRCfIWChdx33MYRp6dHHZc8r98OJa0ScuimINPxvUcU
OSd+XpuK3xXcEA9FWdD7uZjXDsjvp7RArlnl57QUlSq1IW/WjE6x52grfIwdOarW
jy54qHwsRHXY/tsWh1W3KHAAiXM7zuccaxv6w1xAjnSnQuTf69iI3+S9EA4lHGMr
r8dcMKrMUAn76MqNG88DHMJel1FktYJrZYVRtNl29p+iOgMfCs/hJM8xub2FTSaV
ZYb1I97J1GLEWqBrdnXrVAu0RIViL7zLNuqS+SBNO23rllIWYqhdh3//xH5R4TjX
L1ekJP/QNfqs7zFHQx9pigp5mGRyTyaAdtGFlbSFWWTxo7gRbQ90Y0qs0PEkR44e
GMATLkT17tQjbA4i92CfR0heZpNmhAE02TcWEvQYlCQmyObFaqV2/AxsE+bect0d
pyN0KdJrf8gjYG9bKub8jDM32L8zwjufpqeOKsfcLgHuRDvg/rxvqHSYbmS25ATF
udPWRfW0j7MKsQFJU0gFG6Vj3slCPMtc3/2A8dpL31ZmYngvxLqLI7Mt3ohNb8sj
jk5RV+MQ5ypapB2aEIv8+ft2AyvaoPjPuDbN28JJz9iPUkNPoHOpf3bmHdVHAKXI
N/BuYLHrnlUQzy2QtzpNEXV8IcA4PT79fcvFqCYXR4SPua4S0r7xP8NEkWeLBZjg
7IJg2mEpMIwaYh2mZkRPZ9Pqb8t8RPrhoTAmFepHnysZ06z5NlP9BKRRao1vcNEM
4sk/vgVINkosE5MG0xtHVcF8+uMg+rUjDds0d03BOMHjnH/JQKPRjxHo6TfxuGH8
AE63i/PPQD0vf2/Ns4mN3WPuapT1p6fPgMcTvC5d0ECWDQUBCgdR0lQbBKP1dW0x
rPcEBXWfzL1HfoDNDXHXsBltB7Q+ZEZiueX/umcdeBwlj35DonSuLKMq1qtIOLh0
orWIzRuuxSenTpXbOJnGPCNr1CvtiK/GCPDf7vzbfyGLF7J2IRRaZryu9dpdfr4a
953ky6R5cnDGLOqS+8S/5VBzCDnzPb/rIDEa48f71H4=
`protect END_PROTECTED
