`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
if8qoVKwOTe+zrIIQDRbVM3O5s7pg3GqOrOyTNjT5PxvhH+loNUF7bEFeGIwrS12
1++IUK31+wdgK9jex/7+2rGQw5EOyceGe+DlCxBz5RRbsxgnIHMUPOBZFihG7c4t
2dWpSSlyQDCAj4XMRcSRkPncNHQk0fFD0EWHe5q3bfKDvdFu31ehei1qguLL2NdU
BLdPZbI1u+o7K9Tpeiy7bEgBjjmi5BdTqsE3kji+tUOypi7muA3AQbTtl9Lou0oz
WqrWx37Fbk+eXX/sWUCtgz2doUyunzcIQN9ZKzg5361lSyNno1SZLncnQZ9fOC7o
8QLblZycCfqB1B/mPWAfA3j80Gb7eFY7cqQYs6rwwsrpPuLGqPo/L1tcnniu4JnU
Fn5thYX2kepn9Ss1vOyFGjWrhQS8ZCgdDnoJfSTki1Y0LwcA2ZTWvHlSodUM7nCd
P0/pa4Ps8Fxo5vENwlSAuv86n0SLlLJanhPQSkReNNrYe2M+P02wUcPO2FLS8hBs
K7tA1s2tDdIa3jfj1nBIJzM9RxDEdBfC6IEMx5PfDKWFbfUkhljeezoloXWRR6v2
ZAhMXH8IzNuLhFzfXPh1WLps26/5mfBxkUXVRytNCJk9+BWYM6bBpKdpv2cyji7j
HGjsKzjNt8Xj28I1Y0cACB4bV+AjVZQZ8rhWtpeEfFZfg3S98Wk9Ce5nvYWIjyWY
iTZ1kxcAbBgbpp4juHwhtWqiz3icZgMroTA4n3IeV7L10jrNHGaubFAH3DUTG5TD
q2Ww8SE4dI1JpqkvFsWUvGenL0cY2dc0oHGD/hci3b8OaVBVkHwNvWkgoeE2EnC3
5eY6tj4fk4Sfo6TqyH8JYRIiwJI0JSKfXzFkR0trKYX1hM3VD+lgA5L7hWNb91yn
FF2dKONlXzJEsP2MfQ2wD2lSf+yR/ZwsccD7YVskAwK/FsqlqQtnogzBezuFhcB0
l9KSDa++SE9AL2+WyId+WIP34+RiTFdu8boE+Rgz1L7ey0Tl5Fq+MXMa5R6bbMVl
ogAoCVjLoiqa9icfb/fzFv6FEmUcWK8C20PBCy6dLPX6UdZgw/YtIP2KvByPmcES
0F4qTq8Nf9ISZdLA48vQkjzZsmQJO+Bj53zixtgyJtgS1niL1MLEoWhaCAdQDDMm
yyxOACUKtjL0JgG62hwxREk7oWBMMAwTIGCRIRC7ktz4M2TflKPCegrnmIj0mx/m
oHEIWnxJ4829ZCOqZNvQyoLHuGAuCQeeOvPdY5Il4o27Jt6hl6pMtM5QGuNO961+
FhFvDW/fVS0CqmtVZyNJnEL5CeRtFEO0Mk3uj71f4dRe4B5uyYht05a2bSdDh/8z
+dUnjVRNIhJYkCXFSfQFccOQEk0bwHRkfNjxTmPvgDMcmGxdPP18uucmQtaPwJa1
TOWDpRmA+zVNocy8xmXNno9XQI5RfaeBX5mYsCjvrir86kY79MtzCdRw6xZT3Q14
NENOTNQ5e8cTxOZGAQZE5UOACrWnoDb4vCKtLRK6KQ0BR+uenbwpn5zrNIUBpIxd
pvylqZQiwgpUfNkAIIEe+IFrdQaaOX4Yv5pJXr/hw818VR7UPXsW5aplzT7/MvWK
0SQNyj95UVTtDoaJFZoA7h8EY8yUjgx+bCEp2GwtfydO0gi8+JGv9gZ6wMx3U49Z
6dSY290fzee0e7jb9+iWWrArbnPOmnYhT05uQDxnnwnj1CZWuS30HuIYVMw1J/8i
3gUbG/Xnm0gn66q5fgngZABUU87yO1GLxf/lVpBbKbZ5LFN5NMO4YLgiWU5CZDXg
YRfObNnRlIJKV4Xt2J+/sW5dyjtedkMmzsdzPq/ra47/tg7EykaddrMCLvQp+I1t
KVo6+YMqApPGJnHiTozpVQ3dKcqBce0stj6oqZ3V6LIG4c0gqSPEqsFBtL3JHG2Q
jGGB+mqINusAjOhicNWan7oZBvfoFfcHTrSMFaThR5mndMgV/DPnESEeQ1LJInY9
vHSlLF6FMHsJRRQQtxtvaOC0iMDOCveGW6vOhlLfu6jyYk6Up8HdfIRCmyL1ii/0
CWzVCn/Auyb1OSinXtROrA==
`protect END_PROTECTED
