`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhaqGXo/eV69Vk04Fch4P3HceHTjxz8Pm5MLhmM/O9HBhjoIKw4oS4PCi2UlOS11
vCYoL1a9EqimdYtXsKSv6KT1sNUJKug/Wm8uy/QU5i6SCP0ZK5lA1mcZbdtk4fSy
LwjjRTKRfgUHR49FHVaBavIQY6iiVCBo3tsGs1A6I6DOuitevg4dGVxUxq1Wq0J5
51NDj4eVwl4tkj8bXovdRAyvjVoj+gkkRCMudNe+NuY106FtAGSAC2zbMMmvpmlE
r8spf627yT+RmXaUwF1QnHEks6BZ9BLq98n9G+NnwoBlg1/1jqY5v5BLYO+bnRW2
Yj/phae+McbieV3oAzqy6pRdom7zuL4531Ev8mFwToePz3xu4FyMJLhQ+wSgyiSo
T5tarkH00Tw0PIhLhiYh7ghANJrXWDw7NC1bpMpFQibvmldMteY3uIp2/X18AqDy
f1mRVSiCM2+7BU7W4m5ejfvMg5JfLlFjqFs6Y8NuPSeihGa9XrmkVQZQI9fgpHoJ
scjitcoXR5OiOSL7QEpax7RaVOsL70X0R/eIJVql1XPstNtjkT3oRmX1ZstQXu8u
rr+Ni2sAyNGFQu9FADBZDegCd95LALnFXrqlaTxTJuqSZVe2yjz1HTSTXkY0LuzM
KsFe/fqfFJ9a6CAAC5KhXp6RhnuG5KVAb+vMNH4HD12GK73Csba/J+sxQ0L2jxiA
PSN06XUPpO5T2kghrTTvyt4H1K65vDiCIT9Q14jdqcxr7606q5Em9Pb9lCw/M6Cb
KU/rbYnjft6dPPQf2bkDWXLiJOAxX6rckUpuKdrsgOVT7lkMDJSSWrEekURu+eIy
`protect END_PROTECTED
