`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6zZZtWOmRtHlcq+oh2Ft/b/GR5TqvoDCRBY9hiSKbNueOTRvDbFQtcL1GI3+3ZVi
d75KBL1cWmTtZD6+1dht8W1eddR6Z7+lWWruN4dx7Lxr0H7PcqCXMHU5nkng7iy2
fM4rcFq2DQuYUklKc/0ui4sEKLQnGYrIWlaOp7FgSGGtLotXC9hva1n3JBo2q7DW
rEAXh4EYPSnZNELiZZnOmIkX6mxtsQnnzt13CrDLn5pvAScn2sIDVkOWx4I9SlG4
mIyBXVEGVos7LzYLPSJcJJ5yIccdNp8D4E0tBoklUlzp6nrsafNuzI4s51bxFA64
Qx//weKOxaYilrRH1YN3ylTrPAbrvVshCCnpg2KlGkj1tFNXpjY7k6CUFUc5NVuL
LeycbkRSKGUhinD9Xl+7funz1hq/vJHABAE91PnSU1k9cCOJd5oAd8VnGH50KaDL
1QJNWcyqsBUN/+hLLLMe3drqJrdwt59aCgYFUkr3u/4T6wdul/C5JNyJLQuAQNMV
lDgqnDhKJFXFIXQRPde/18oJ5l0umq02QOkxzFh176EEOKai2MvDRnGZjr2udG04
BXjo9boBYLZYkU8k7d4ANtuAuiRjgOp7I7v1tfgL/W/y4pIa3fuaG4baAX5gmfUJ
RHplveDvxM0GTBeZitinE7AlayaGZtc/um56GMBdjEniNhSOH96OVjbTnXISYvvj
He4FJgtytclW6cVr3wGG6IdHQZ5+sAJgnsXq5R8zeswTw2fS9M5OUpvRVgbvVfY1
N39sGgh09nv8UMX1cKsmYLl8fS2zISFUFRBOWXbjJC4dHs74zgLkGlsW+tJTUx6R
XSIC2GKsHSUqec4KvnY+jLQCiLRoykRP0ESD5Wt1cOFdR6NyHB15rFfyS8wqVxtX
8wdM8P6yjRdf6oq1thi/vCMvPO6I888s9bL1KTbBRrcJZs3ZHahOxw9hSqj9nx3I
IETB3Tu8OfCvgmrRw3gtTg0jxlZypiWhadoYsBy5sdBrCKW78HrK6/mqqyVDksmW
YRuFG4pq+yYaDox8ErCMew7quLmY692VFy/B78gdvaI5jyw7frgcGbkhcVxFUdW7
Qy9ZwYAjLkrEaKFVRtFPnd2bJkICvLMaaDgsJzqSDtXqRS1YtSgQUyzlJPQyzei4
OB8KxeAMnDVWwFkcDvxRfYbup2gCuJ+xG+AWjZcIsSTyBNjdWvWxDireKNt9cn70
R3HqPUKRB4hbchHHRdjP6cWaYxffW4JbrL0rYyneFOzO5ztZTCcP/xUwLxj2TQQB
M1RuctB0YGra1CjC69jHpqTfKv6vbxYWSp/i0aYaSqRirI6wan0e4NGZmWdUbzfs
DP8NUMNNma7F1MLhekF9gAho3P7ldcI4XspvqK+JbDXZgpgIWrgdSiYtHnOm6SdP
OcWsGFJVZPRtfRV5eFBd1iVth9ZdjHuloXoc8HP2gTT+LgT4Sg1HCSxoA+nlig/N
v/nYdqMknYcQj1mBh5Btq6nVg5vIbMGIsRiIdi2hMQ78UguHfU30e2R5HBBrv4FQ
oKFcRcgfMbGbUkuUd7fYJAY1Us3MH9SHvohWKwXRRD2eE/T6tHeCGHANW+6ns2Or
hS0OmUsMq/Nof7wVTB+pVReZLwasclnJDyDjXwFGdsC4Cf04umcL+lSZo6CjGq8K
Q8kKndPY0998HJWXtMDVKUMQDUT6bc3N5hZ+XaM68F5++ASEDmjjx9Rry7JYvH5f
4855Cb7IWSzhB+C9i6DaqtvOpgCytw4jh+wZVWsI18Gnf7fv6izZ3KNyJiS8+nxl
2YCwSN7ZTrenk89erQrzjl2cC13nWRQV/7h2/MS9SUmyVPy6S3zX3Io2jWPsuPuW
2v6vs+0o5+cA+/31o46Z6dMXVywW/xkPstWHelKL+qlF2ircbUIqdM6hUfRoDNrO
hjMnT/wfI5oS7R7XkJ2HTw==
`protect END_PROTECTED
