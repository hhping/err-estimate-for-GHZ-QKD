`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWU2FzF+dMBwx468XO+d+spZqMtg00zbVFHoyhPxw+LI7Wl1CoixfMCOsYgvmZGC
6/M1x1j/lVxY77dV9Wb/VnCrs3aipQ33Sntvmxre+CpxvccE8ubtYzGSS03ayLD0
aKWZYSnnQWt8a69swM6IXzi788eswgTH6v9Pfmx/g+eA2ptGqtYR5uPfjaY/fK7J
wgFNhIHyw/4HdRlpSzbOwQdtpnmYYisIZaMfZZqU3lSEmnHl8LOIwX8Lv2Q5ssC9
wEKXsAS4F/ymHbggJ46e6MqDBRi8lV7Xwe+lYqNMg44LxQ6fnDJdzfSjBtgIMXwD
JLxDX7rDQ1Rb8jMR/bE5v1R2kTuhhBY+59/0AIv+Vfu6gnk8StWjLd3PIJQxnQcE
qSdZOgkKXLVWVd8uSvCgo6SJalREJzbLj/GKLJwRojVIFCnFDVwUk04KlmEtU6Hh
57banmh/50n10RbTYejN5KYcNXyh57aNpv9DJTg86BA5bEdmnE4Ok+43aafJF8HW
YdedC5Bp/trhPXBWQ+eKBQ+kY91wZ4S5jnyVeCKDe0xpBqhqi1J3Nlll30w+Wm3Z
NkkYqgnCLQ+H99NtGU0LiAct/XrYmibgncClC37fKZbH7nY7kgkV4qsT59Iq3a21
8RcPnO61qvpdyi0scCHK34PoKc3hN+lgh8R+JpvfKmoRcVWRXjqGUtyILDGYNBAz
wY/1S2DczHqRGjL57JZ9UJr1V40QV7SHUOJ0k6Ym3GiMGaAkmNTlSvvlaGSdM+rp
tv/YajH3ikq7Hc7hWwLqGLKI8B7PJjKTBwAyYIH5ShAMFgTzI5dqy7NYq9GxmaRM
FvY5X0zLjuclLRniqMO6sjEQlgjQSSSDHkgd92tKQsKskybOCYhH8s5tt8xA2qyU
3ChKhlVD5uqNNF7+9gkrC0O2G+h95ti61T1CRIEuUQWwtBgM0SV548a+Jy/SvEVt
9MjHEHr9GqeBQOA6xsGo3dV9K96wVrqpe8BKJVXmQTTLIPq2MqApdRDAKZzvvfdR
8ezVbeogqUgVjhW/IObpUZkFw1hsPlKGm3ruVZJJCzuvapv7J1EgkIRtdQwv243j
+DoivadibutCLbmBLVjc36iGcYe7fjQhzmw3u98iw56sr5jXQcyJVqGDnyg9rcrK
YR5/wqJ/L/P74K7pMGUqeQAPXVxAzkfSv4/b3ruTxhTQ5lNODFc/9ZV73B+TdTCI
o25BlonYif16TCdZIta9JLIkQhBjT45yGvhVka1neUGNvjAyfwJ+7OMk4C1uLb+I
cHFr52eNm0pS20r421adyaQHakHmTPZx33D48FujLjIJuEPEkTXHo/J2OA2eIidG
/Bsi+T3cYlqIvfhbwYygnIOD0WYWHgFa3UaimpZY0GaI1JuMPhhZ2mpTmJ0S2883
sgvi+qtDDHw3hxmX1Y1z1s7I1+wLTVwOktsnTjfgJIPiZiUpA4xfAYnL5nuoRCNp
fg62xRtL5AUfViM3oM+g6yr+6kZtLcIfyvnJBc0YkRkevlZ6bQwonHcOqn4p05P6
H1xI45keVQ5xHfQKSeLKCmuiXNKkL3/MpDJ+hMpp5J/hjCHBmGaKINHrikkHhtGT
/IhmAVAEsELWARwXey3nFh6JYnos6oGcfTFdIfhbYQHHR/o0seRUNBVy5T0R5nL8
/pVNpGtT7MABNXIU2VZxCD5dmHXTZ9Mk5iSQSs1LzvIyrcEaW1b9uJusB3R1CcTM
xbbmH+0yLuwF7RfCqxNxlTowbf9kQ1AuPL4hJOgLDIHrfnHasIwrw0KZuwkw6HOE
Z4qmwRhMwCyrmJAjfSQUPalTjrENMcBS+MuVFfavaZVscIAlJ78SzO5+POr6no3P
DGZrZ5TgxWAKp2hpL5FajYgeYUHXxIJj8DcSOuZM1FBUdNnigsQmnVF1ZXWWd78e
+pcvNSwfIVY/Dm3Roc5KgEJn+eLIPPu+kT8u40fDxbSNK7ARJiXeWaDpGAbswguu
HI9EK3WIu16AE+v5s2pXgRJlixa2SaYaxRjamtHNigiVyRYu8ZSn88wjxGkUwwJd
5IZAitJYiV1SqmndSrNobg+EEuDnyeow1Ba80Vypc8iQFnA+XV+evx3z3iu2a9hA
bumqjU8bzBQ2kkBm8in1u6/d3DANL9r5I8UPvo65lSGJwIZGz8DY0NtJCe5fZBbw
nO/HLubDQBcYe1q7m4MJxE7qAGBewMgTWYNGujdMdvO02maJlzAkdpLED2MEiW8I
lwir0XsdTb8ttN17TPdP2GpzOoDajFZXLY+bSiX5t9aRy8BzAz/muq8GBN4Khvtj
S1dbvJhEadl8/592w64pOyob20ipaGuSg5I9NNwdXrqdx9B1o5UhrtLL0JIvBfeb
WFFgErxVwA05s9zZnmXzbft5iujw6fqkQnS/V9wKomyWVPqtk+JPaYUmt4t8f3j5
pLnsqXgF7myeONPnePh6sNXe1tGSFM7Jb3+PUsT3Ap9fGt4X9ZiOuESzzZJJJYnQ
BsosSNSY+9k9Rubrmldnm43frY8C55kpmKzmfajyEPvSB+akHAuTvLTrg0Y3rrwJ
cs1bYwJhiLUNce8a/QSqZXskbeBZbfJ/r2Vf4tCgIwMMNTh8oa5AroQWa/c5lGyx
k8I4UbHWs6kGtyUB4VtFveid3WjFvITmMMCH+p6M/20EAyCInMq0YKVI/ce+oLaD
4H/V8vGiP9UvlNCHrTyFEdimzRWcEmwfSky3gUtu21T3DUZ+9c7cE/fA0aVLVQxk
BCw9wjkQWHMy3BKgrJC8UcLH75OYnnQpyITk/dFvkTwISJBKIOYNcID2ZMivvTUT
z8qPf5+ONB5U2wq/wjhmKB05C5mFwKPnawkSK3f7u5Rs8LGttvU4AvO+x9PS1Iv5
stHQtlqEt9yXmO4x49U6zL3KN7znI/khLuKSQcl+UBg+xINJ0MOI5fU2vHsAOdDS
JZFmO4CtuFEY4W8I0aGWM6Te7VwVb4FsRIj4JLAcanVx0JTDnm5NtbnI8WFYJlja
vtFJZd7YBCpC/uyA6Sn+kKQHkSldY2jfxMdPeQ30bp4G3q8Ca+zb8eKR5jlgjgfJ
eNG2HeO6eBPxsPFG1vkGWx0L2ESp4qhi3JWbp8b7zLP3ueKXdLczzKdomQ9NqWub
bHsSPJmDUWQzjKCQfzQcfWwZXWGJbmlv4fQxJelWxMEVjrfh1VO7TlGLqqPh7ipE
VR664GcafUr7GrWjoIjvZthD7bBUnZXM+zbH0hO5jSxG+8DWuj0fCsr1vXlDxyp1
zo+Hv5Y+jaZcpOhzwx98j4gHAZrkwagZT5NJnXuHzgrVR8iTbJ25ki+9ywsb6HX6
JDA5EKTahU/DDHr/f3QTRkppN2LpfXmWVmwkmIFpc/jmqMY7sGG5JiT7jygwraob
Pv/B/Z5J5laWZkl4yy2G+drwH34yDH5x+vWGRLnd2DbKJw3BYAvAs2znMVWNGVkG
HtwErnwm5BAJKJ+GVtz/Rlg5lUxIk2rNBbGyDmSxWV27qwXniVPdHNmBckcQCRl/
WK8A8C/ZaZPzP3qnYu7Na2OufYL2TnqPYjhOO2qxXBfyC9oSFUeTNn0MVt7bcbad
4gLnSvxJvH2popZkim3pT/M3Kchi1imTl9bImC6J3wbupSQUh7y4W5fRgTK9EGqz
sKA3wZAxcHvEDcsTAOQvfFBkZcGDyfmGyG4+GLTrDN4Dw6G/LwoJSA4o7yRZnkTh
iGdO9Luz/GFMXYmEuCLzEKJxpVkujEdMSUm7/tCkUAPT6NXV5NwQdKVxU8xGbQK+
g6j9Uqvqta1vgQamufvtmXuwYmYQZPWMI4pQLKbePMJPRqLwBEDu2WEuGGhD7k5u
lGZJ7huxb5KVqQG0Hs+jnOSTFPce9y4dzTEJgnUSQHjHAct7idf2AhZCNPLlCGHx
IlKWftMV48vAveCTT+bzkRG3SPJcwR6J8U+e2+ee/7M8qtUc+Z3BZwGjD1bjtb+9
BxQ9Ol2cesR3sivjwBS4RJaxQg3clayiq9xltL/MP7fIx0bNSbNaoKyGTnRHO4QY
K8K8i9y6s8wgXpVnzrHDp+wDT+g9dSYju8pgpIRFW77xLlG/JGi9h1Hz0LhJ22By
eEBqutX9d6PbT/QyYrQp0M5aCpsVynjwRKyDLfYNS/lzJk2k/gAkDrWZG8pkB9ex
uinkjJnZP/GQrFUzefbg1txfPpXAdq8ucjo0Sugueqo3Ls+T5JOe1fUM6GNXIviB
q8IDzS6kvQCf8feTZ42eGMhsc25AYYu+Mx2ZvS9FmCaEM25bMsGvKEEuvcSJyXv0
B4pg8wpxg+I0gSQZDmpd329/1Ek3js74IthZRHdWc9900YC1JoSvsTm9XvcXyvoG
acLMoWRbgt7De4rZNOHeX+yOwpPVK07EtivjN/px7Vn+BrY3hks4HfveaqPxbPg0
wlFEEmijADZ7rjopEoJpwS+Ik/DdgxMmdypZ8ZYJ/oEAx3pz4eqJK74sgMZpPi9I
ywQywJBdMbiB97F8MO4R51EWFhOlPmuGx9H3O9oESsxzUtUqTf3IaiIJet+5Ypw8
kVid+H0ReZCKxKjMNW2tN56EI39WZWK+MNlXh1SSPjrRbff8XA/jbtl+5lFa+Mj7
UrgntJgtK5YsZC8pHo8MnOHtA3tuIqlX6WFwCFjxuw006AqSqMhUG+2jBoTWWqD5
6lFb+UGK9CVnoHzLgydpSPBEWCuFDxBepxM8MoSFmUxnQc3Hq5AKyLeRMuFLJwbM
mUaeU8WsH6Gg2TsN95YlFhGvkXWtE/v4MmmbBUtlbXxKwdFpXEIs8SekDmbWJIZK
HeMiUzbb2yZGW/w8D+h5qQm39rhaThPbGrcB1ALLfsvCvwHaGqdM3BVL0nPMSisV
6+D4LXHaJLAEJ+gR1YKBWzuS5jAGZepmt7jV7khi2SCaxvpRY3ncAb2pOBwylxJF
F0TONVLAYS9XVY7qtW2wcXl6tOSgWdkxKakEkD5WrBrqzjQ9+WSagBDbml2moM0y
dM6E2mnFzYy5AaH8K1k3mrCs8t6vcS3dXGHmQVUx+fHZ7wKiD30irE+cw1snEjKh
7fg2M5UPdqoiwtp0TOda4iSB0+98eDDSZj3RGn2P81Y7KsBZBjOjvCEltIBZSUPL
wtSTQlOaM1NgfE5GXSZZLuElCZ47VT/Ta3I1PavtZ4yX+gXKPMrC0BC3W7a/uK3P
irzhugMjr6GRP/P6gLxSO1UnZW9VLg4XL61J51NyOAiFzGVIn4s9HUNQJ4LCN4WT
befRgpXs22bQBl2TF1Hl4bZkCQ5OphNoWAhCuGkRnxfpIZMOnZ6x5dSR6srgEPtk
8AjzPxMH6B8g4LJUr29Cf9Osj3K05LB9MGn+aw+b8+wZkSWLF3iTlWYpl+9hdoR1
DQeSBnapUldCdWW4OzUEsSEn+60rrfbRd9ykdFNsHfBcBSlEb4rbUlK58vyvUQBH
ah2/6cwDQKMd0FOQrUSBwL40rHLd0VF2AZpTFc2Va/6iYltaT8DmWCUDCWfQQWvu
yZ7Ifq/nLHtBC+KunFUlmoFSZ6QIjqoT0ShScObNMNQMIdvG7scLdZPEw3U5B2ZX
9A/M6v6OVHi4fdJTVi+TyrqfWqbb1cSvdEHYvEqU/BzxUkrSrGL5Ni46oq0NXcQ9
mnMcaM44E+lft63mMwHB6/xySmp9BVmKuVQa/hJWDpThmW+p1W9iH3jFz/28XGso
vMrya2hW9qKCLgCljmF2vbgQtHyIL0NUctP1llpDT9DnFZvbqJRWCfz/cfXqHZ2K
inhU6r/5z/EbtgZggC1Ovg==
`protect END_PROTECTED
