`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lV68Zw9fp1cnMjtSAFSHOiONkbOljTb8oICsJpeKBYH2wLesFOktf1W/95aavX1R
3Gd5KloCZA3/MO4f2XTHvYr/jwzYeehsEb+eICm9YczVK9qqcfGSYLXmoUR/v9F/
kKbWBl3eC0GfjKB30b8y7zBn7bPt/eBwA+YLEr9X5rwyi5HDNTO5ksRDEDz38pSC
nCrg81OqsrxOn2MOeX9Lxj2Mui8YN/THYeTdQsKDTAr0i5UGXTBDTjON7KD0pRWA
mjUOM8208WKonAw2UPzKyJYIn3Z84ijBBOlBidJQItg53ywEyBX7N0nh+mtx+ogy
e9DgkDFghKL9P3xYt6iu4xSmsiKWx9yYShhx7Hp0pCoLltcQNW9XHbeJE6+ERWMt
+IM1Zz9AiFOJjipkEuj6EskUphXzh1yHUdJJ+VRq9E9hcejtihmZItEkVlSmSykZ
bBPHT3owdb2kctgTLyFyCetKfNi/ofBkBT1Uz0ClpMsA5sa7DIBOT9dFfTVYp2uB
uYDdNXqF2QpXVKQQDKM6+OP/2GQgDAzGYRrmIgXwj/TenzgOMp5jLiVE85qMqidc
mQ4Notkzr6uJbYp1Usg+vrsOaHwRye9x6Uc8g68M0Cbl8N67cC1Qqchn4m2XyHu+
BA59QaWNnZiy8KPFd+Y7sls30eIIQnTMZEkirBplbyM/8Af6EjlUYit73VGkjbDO
Kh1w8CY6yT3BfK/cqkXIKl9ltUptodkkDWIFrszt7HOtSNL66Wrg+gNzolMNR2dT
0X8DB9EkjIu8fnDgOg26pBfYdAuaxCg/QnamLQ1r+u9OE+c1m8oruzCaS9y2Bqoy
A7uGcpoWQq2BZnvdbV82fYsOAwQ0FfBYiiegN4/Ac8BuGwEK+lf8pPwd0IQH0aG9
y2CPAdo/z1JIzoERrxxZdVDEskuy3dDClgXg0COAS8FnF+/jFpMFrEWXZuSJm2Nz
TZi2JrV/4Z6P4Mm5lFaxqhnnaOKRYCglx/K8boobZto5NaVvYlvj29/wGR/F+nBl
tgKGVkf4iz66g4jynQmwdzbmrPWc44iHtDQVoCNbWCY=
`protect END_PROTECTED
