library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pipe_gen3 is
    generic(
        enable_debug_info: string  := "true";
        bypass_rx_detection_enable: string  := "false";
        bypass_rx_preset: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        bypass_rx_preset_enable: string  := "false";
        bypass_tx_coefficent: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bypass_tx_coefficent_enable: string  := "false";
        elecidle_delay_g3: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        ind_error_reporting: string  := "dis_ind_error_reporting";
        mode            : string  := "pipe_g1";
        phy_status_delay_g12: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        phy_status_delay_g3: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        phystatus_rst_toggle_g12: string  := "dis_phystatus_rst_toggle";
        phystatus_rst_toggle_g3: string  := "dis_phystatus_rst_toggle_g3";
        rate_match_pad_insertion: string  := "dis_rm_fifo_pad_ins";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        test_out_sel    : string  := "disable_test_out"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        blk_algnd_int   : in     vl_logic;
        clkcomp_delete_int: in     vl_logic;
        clkcomp_insert_int: in     vl_logic;
        clkcomp_overfl_int: in     vl_logic;
        clkcomp_undfl_int: in     vl_logic;
        current_coeff   : in     vl_logic_vector(17 downto 0);
        current_rxpreset: in     vl_logic_vector(2 downto 0);
        err_decode_int  : in     vl_logic;
        pcs_asn_bundling_in: in     vl_logic_vector(8 downto 0);
        pipe_tx_clk     : in     vl_logic;
        pipe_tx_rstn    : in     vl_logic;
        pma_rx_detect_valid: in     vl_logic;
        pma_rx_found    : in     vl_logic;
        pma_signal_det  : in     vl_logic;
        powerdown       : in     vl_logic_vector(1 downto 0);
        rcv_lfsr_chk_int: in     vl_logic;
        rx_blk_start_int: in     vl_logic;
        rx_sync_hdr_int : in     vl_logic_vector(1 downto 0);
        rx_test_out     : in     vl_logic_vector(19 downto 0);
        rxd_8gpcs_in    : in     vl_logic_vector(63 downto 0);
        rxdata_int      : in     vl_logic_vector(31 downto 0);
        rxdatak_int     : in     vl_logic_vector(3 downto 0);
        rxdataskip_int  : in     vl_logic;
        rxelecidle_8gpcs_in: in     vl_logic;
        rxpolarity      : in     vl_logic;
        tx_blk_start    : in     vl_logic;
        tx_sync_hdr     : in     vl_logic_vector(1 downto 0);
        tx_test_out     : in     vl_logic_vector(19 downto 0);
        txcompliance    : in     vl_logic;
        txdata          : in     vl_logic_vector(31 downto 0);
        txdatak         : in     vl_logic_vector(3 downto 0);
        txdataskip      : in     vl_logic;
        txdeemph        : in     vl_logic;
        txdetectrxloopback: in     vl_logic;
        txelecidle      : in     vl_logic;
        txmargin        : in     vl_logic_vector(2 downto 0);
        txswing         : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        dis_pc_byte     : out    vl_logic;
        gen3_clk_sel    : out    vl_logic;
        pcs_rst         : out    vl_logic;
        phystatus       : out    vl_logic;
        pma_current_coeff: out    vl_logic_vector(17 downto 0);
        pma_current_rxpreset: out    vl_logic_vector(2 downto 0);
        pma_rx_det_pd   : out    vl_logic;
        pma_tx_elec_idle: out    vl_logic;
        pma_txdeemph    : out    vl_logic;
        pma_txdetectrx  : out    vl_logic;
        pma_txmargin    : out    vl_logic_vector(2 downto 0);
        pma_txswing     : out    vl_logic;
        reset_pc_prts   : out    vl_logic;
        rev_lpbk_8gpcs_out: out    vl_logic;
        rev_lpbk_int    : out    vl_logic;
        rx_blk_start    : out    vl_logic_vector(3 downto 0);
        rx_sync_hdr     : out    vl_logic_vector(1 downto 0);
        rxd_8gpcs_out   : out    vl_logic_vector(63 downto 0);
        rxdataskip      : out    vl_logic_vector(3 downto 0);
        rxelecidle      : out    vl_logic;
        rxpolarity_8gpcs_out: out    vl_logic;
        rxpolarity_int  : out    vl_logic;
        rxstatus        : out    vl_logic_vector(2 downto 0);
        rxvalid         : out    vl_logic;
        shutdown_clk    : out    vl_logic;
        test_out        : out    vl_logic_vector(19 downto 0);
        tx_blk_start_int: out    vl_logic;
        tx_sync_hdr_int : out    vl_logic_vector(1 downto 0);
        txdata_int      : out    vl_logic_vector(31 downto 0);
        txdatak_int     : out    vl_logic_vector(3 downto 0);
        txdataskip_int  : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of bypass_rx_detection_enable : constant is 1;
    attribute mti_svvh_generic_type of bypass_rx_preset : constant is 1;
    attribute mti_svvh_generic_type of bypass_rx_preset_enable : constant is 1;
    attribute mti_svvh_generic_type of bypass_tx_coefficent : constant is 1;
    attribute mti_svvh_generic_type of bypass_tx_coefficent_enable : constant is 1;
    attribute mti_svvh_generic_type of elecidle_delay_g3 : constant is 1;
    attribute mti_svvh_generic_type of ind_error_reporting : constant is 1;
    attribute mti_svvh_generic_type of mode : constant is 1;
    attribute mti_svvh_generic_type of phy_status_delay_g12 : constant is 1;
    attribute mti_svvh_generic_type of phy_status_delay_g3 : constant is 1;
    attribute mti_svvh_generic_type of phystatus_rst_toggle_g12 : constant is 1;
    attribute mti_svvh_generic_type of phystatus_rst_toggle_g3 : constant is 1;
    attribute mti_svvh_generic_type of rate_match_pad_insertion : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of test_out_sel : constant is 1;
end twentynm_hssi_pipe_gen3;
