`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJD40EuOLyJEpS05Mw9QjN1g0Ojp9EmCjDkapuRjjhoJrfB4A2iZnhLzBB6kLPbt
PTB9SymGqj4cKEcJM3tYh1T/lZ/G/i+TKYnd+bml1ko68FndCwMqLyvyC/2aTyPV
hSjQoFO4u81JbXY0r2APxro8QGQPmeeCz9KnbmrPoHmoc+2FJygEX4dr/g5iuJzz
mzxxI+Q58AN8S4BTbltSAFatlhC7w81VcqW/kpThzjDZINj4/MARcuCcODdLeaNg
pFEpSjvmPBc5s5VyxWqfAqEaf8yAhmfeVn1EjpCom6HeuBkIhrEHxYwoNTBC2QCt
vxV9KJLhGFXg7VwAdxjfoGNWeYsjZVtbghl1+CrK8KpCQsCUbgWMDeO61P4K1h/g
WqNc55EP8rLT3vslc/wpll1hl09uZKKYRss6qIm372YmXzzwNmoB4wEp6WUANLvf
PXsPBPJSBizLTxM9af9SwdSioFRqkR7kT3vRFh8yjgboduObJZ9HhDtnWke+zD3M
Iok3zXKPpfJn8bg02BG48V0pyM7fGZsRpTZuuQD9AyyysPWSyA5mdtAVIdjsiwUP
G0pWy3Ss/gx6ZPlT0Yvxap9Xc+02jqPoCK5Vs9qvXQu7h0BYw/n7JKQ5K5UIguwZ
oogL7AQWA4zgNeYpm8J7TBzFknSyL04QFC9T28zWNiU1Kc4nBvF7GpR+A2kEIje4
zH4Rr6r7MT6GmcLDL3aBNFHPxPuDJVpCeDUOo4EM3gubJ1SVrvBHa9l+eDPvC+CK
06dNy0WgVNvXsMXB7bGGdYrAief7U4RUfN5AYnCEMc7lmTHyEBMgPnWcTRV19BUU
bB8YEGGkmKVKqr46ZFkpxKmsuewbY5wqOsms9P0KVWv4v59ik00UiyU05pyt8gBY
8PAMmXst6NDfOLQKGEAuU9C574VAOWKMPZe9KZzdaqlOFok8/ETYftjn+5XSShF3
ovBDG9ve8ePQ83aS9yOa+xa0ZEBKyJHO0l2TYeKM6U8qJz8miTu9AXZ7cHSo0rkh
huZuFJ34GkJ3/Sxlvq+WKvVPVE3NPTV+w4SNvgJGbKpGWKloiwSper4al8F36T5W
xLUAKWBFwNXx9qFaup05dMNPOttS9jgx+kRzSfvOM8oH4tOKXatQCFAzxyfrLEoJ
z1wSBzxMsrqgW+T30OruRzFAIWgMzkxKYv4cWaxdvQiBwumfJyHw2arEj5fo/obW
tAVj9vbXfUovDQy69vem0SQBNXq0wfoC+6cF+DWdh4lef2yrHjROFI5R3fQW7T7y
pLNpPij+xfg5rJj52VOarJeTPpND/E/ZBUYkCuIO5kebDbXWm+bIEW9FE3hsEsZK
p1KV154TMQHH/mVS63ORBJtmKsVBpedyqBFHe9ZkRD5T7TJelVokj4e0xRgQk96E
75jYx1z3wkxjYwtOqQZJpFb+CgN7AaNptttfwv6DyxjxHAXoEM8aZYzQ+fLAdpFh
bM5OidC07YwBGtfppyHbTohC54p/RGPM7nxYS7F5L3Tg2Apxf+YCZX6JFe/jrkVS
bSxomB6eii0CmziT39iD8Ptt0fszC0lFx1Ui522WRInu6no9hZAVKjRUGd97DbZ/
6FlymI6bKF7u2YMbU0El2R/hXLXMatentiJC876aI7EWEPYn/fom27aBIcg84UTU
Yee2IVkG4A0nEe22+RcmynUbn8I936eQMM/CWW0brDHAmaldMDCO4Vp4pitWB9b6
OU8GRaewfNjyDMOh4T0fJpYNDSfkd3lIxeSPqWIAZcXMxorp83ETtgxUKGFhPfdv
222q0eIztAz30CQ1o7dBWM8m9cYpyC1wXY8tw34tDD0xP8e21oN7nCn4uNY82ceP
IcL/GWj8kIXcbnV3CQ4as09PwOkfP8WxxS672eFtV1HeYgCKUXYzUfGzrs5ocunI
xGqo0GI1GH9NA7wmOK5TfpyUaJE4qYQJRNhJS2eqJEE76pwztvUoAKCzRibkg2GY
30DpMvA0wIfSN9MTnHDe6zklMGKOVEHD2caoD9mIsVRaFlN+R4Xu9yCraeNG2Wnr
OqJrZjWesC6xS0gZe7kHVIIwPiJhVi6Vfk5Q8lepmWpWi/Atxr7VZhE1DUwb/7p2
Lbgbm7U6BFqH+iQgCyZPMCpRWr9tGfJ8oWtLIbOV5L/u1X7RoB7oCdy7Q65hAA0Q
swzQBcI9ZTAfRgO//N+hAYFSmEmy9IwSGeGCuNNGGeaPfb1kmQ/J6OH2+FDqWbzz
oyu8lGou9z9HtJhuFySNVl/M8EbjqvwIqJwPIqPKYyHCyXIO/ca4Q9cXqpl9xqay
ReQSU1xWD6r1qQanUAHdbHINAM4dz9aAfqMrLW7ix09bgsQCrl2AI3atPZ6gC4pN
i0SYvhhl05Fq8VSAcUhyBlQhcHfC1kvrBkiVpwOv/Wb4pTv7TIm4Y7FMoW2BcV/A
1fbQZcGM4Jx+JNdfPDSBBixDNFBQnjyzbQd3yxWQjoZJtDpMuwTboBxIXS8lZmTd
CP0+3JngnrCgXnM6umktr8ke78YB7gq3pfq3DDK1tA0OsFs2NErFOUNEYCs2o+6s
+NJzZ6TTuk9ywWjX8FucvhEwA+Gix9PhQUFu5btUfA4KNgTtO/33w7ZFu6P+EyzP
gixnU/hVdC1lDhsWv6sTEJJJdNTsvoHfVEIZFkHi802nKh3aRQcn7DrVLn3OTvF0
6ENnHxea18PmqN9YXXn/vYWhgqswpl71B9dxIKDPBoayT79YzeC5bibt7h+dfOIm
R5TlTZ0rbLfF0tA5ONeI7J5DD99oWBDdF+btimVLw+KIDivH1/YyzcyjfZaWPAhd
b2HcySgaMio1nj7CLRF7KhXHe4H/rmRaCTeDjcTAtB/Wy2v877KnXqPEcGYUpLkc
qGfRWUG4Ls7sKqxZ2rhF3cpDVS6r1zYSlBqLW4PinYkvtCDCMGuSoo3BqQIVkKnr
qhvMn2FL/bVGq/8rgQzM2Tp3NBI2eibhFdg8i9jl5vUPuOL65FKo1rvDbwmH90DA
RUsKU5vPmnaEWX7ArmeTn6LJx3DrnNvpGNuUitxFjtP6W21TyaJu9Y/HJ1EWcKSR
e2ioQCwwogyv0R0ruI+EvlJIbRVoNDW1TZm1kAJY6/u1OeTMx8nNsYRwsZ/NpbEZ
pbvmIVvCCyL2tc/OKzUjvXbWKKfFdkG6HQRn9Qa7Bll9WiVxsAMTAqmOdRmqYVt2
HXrRKS6iPyM0b5DyCq4WV0wRHJOVljRMbW2vZMjGU/ulSvIMhETHxUrdWMGZVPYe
8l9fhH8ft56CXF4aD734jUSyEqeMSq86tR1pEQnX0QSv4dF9xEw9spgBfbAhEqDG
TnnCKjbsh2K3LPh7pfP+U2T15LjDERQdWfmiA75+Ubu09LTiI4DPWQRmxRGiNUNb
7weaV/X4dKB7nzzyTpO3Y/lvNnsguJHSDyLXNBN/MzaRti04ad81Nkv045eziKS1
BKu/kO1QknNzAnMsBS4wgz3xaWlqjNu/y2Ks4KyTfARi77SAKuLlDPjoC5hqq6FW
qy2S28nQL4BTOOoIRdEQx8Db+sgg0agW7A4sflQroS8JTjk1C6KWPKGOZbeSx77r
7AZX4RiVhkm+SxiMRcif5/qfAn71vWVUrtJpesA0Sw+VCCTrhsNkhnavWMchvYav
j7/T+F4Bg+etlPMrtP+kjipz3kz6ZBxnqlwGKxagDC12Hmf7gkeXv1VZz/noCmhy
xE9MHkfv6n1ZGnYSlKhPpNLuzjFYScbK0ohCrWYFBfgVnjnq8nsgLVzDEcY/NdiX
nwysp0mUXRsIRCMHNvewy3rFoBL3yhWBrrxw2FInBsrruNrn/9NjpDktOyxhMQL3
XAfUEj9alWOjGOJT1HIR10PxiWtyK5hHg4jiJqY0VGpGVmdCUZ+Zih7/qntOGyfb
cjFlIeqnfVz4NP1IK3uxmwKNS6hT1r85xBjDgw7gZFHH/ljpJm32sahptElzWgaC
ZNrq8Q4jUMXV0AZVL4Ki4F7WdpWVDNC0Xg5p/AVeGMbJNfLznTtG0JRXNl5i9JQf
/LisyhoCOMe+YMjpN41CP2VwLZzoI/axwnCz6zGitV52lb6nSNVD2rjNTf6JvaAU
YqyMzDKazlrC3MrbJKbQPxcAq3Ty6Crq7UVFOurKnET2Yij1Gx9ZxMA2pCT7qj0Z
vXDevHaCnvubgmn0e9N9TbCmhMEKn59WNzd5KVNE+HKfJuD/BQ6GuThBGurBXEjZ
7A773Ya0F+vEPW8WY0fs23emHW6RZzUfgYiAOGdLXYvD8qgct/0kuRkrwVVB66gD
n5NzDg3bHqkIxENlvyEU3Pl9NGJnw0jA8rHM3gsD0CbwgKXljQpkYKsl8DgLxGBu
I84/8h3q/J70xFQOCRAygr/aPFcQM1FLDLwA/hJdoWFt+VCBuJqQzGhzz/yF5YVF
/+apXnsuqsFov5SS8daZpbosgQK5rKD5TWxkNLAKNnwiq7qzWx5mzjXHrsIfD+Na
gGe7aQpxpzU4Zgox0iS/OKkLlRMcXJzY8oQsgLcLjBac4/S5JPof7tyiBWha/a4a
+5dS82fvpvRJGLymnrn+NpxcXZXaY2zDowQ5HhtqT4aM19/VAGZOjJ3VYhh+4ZB3
IKCp+qC+3c4jT5MhpNnQM7oiG1TNBVnWK3FBAolC1bD4RGWrmnPrNXCKdyZH/8cT
JL4habYT0abMOZOrMBdTaJ6Zd4aLpHatuo/RNYHOMLEvHZkaH7wD4eoXPsLM96sY
aTM7FcmFNK0W+xzQ8jgnE82pv0okogkKlF3r+MaZLUZ+rAguVdBk1dmcgWmU6Td/
17HXMXwIYLqAdF2XJIoffhKNeFQaxa2bGxzrpGVHvf+8DKHerwrvuv2Az/Ip7s1E
UAeAMUXSmEyzm7hsNp3nGJEYxt0XWeyl+w+RGZl4fOK5PfQdrMCNMYqHMqdYktCq
jGCqoiDBhB/+Tg12MGCJ2pf0temM/XFlaxq3lsN3CD1etDgPqEacYCKUiezklIAd
T1KA+9ilGI/z9ZFrQswBb9GlqMsOBYvp30N/OJpUK5pHe92YvZin6XFqcudS2G3F
ILN/dLpRVlmoJeQuqEZvU6uYA53lB8yTDFHjEhB7JN+e2zfq7H+LhTwy8YQPxzCu
g+RSlfWcJSLzc7O+YQpKA0QIqXvakCEGhWkAFLZrHERSc6Xj1jJPj3Hu6KTt2vKB
8YzjY1njJ0ivg5BqwdaMLeSn7f7lq7y8edGzk95btK0=
`protect END_PROTECTED
