`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7b+APslgvHBNfKgl0NXbTiw+fcsBth0oyv2RX9dk3As2zg3B8M7bbdXxuYg0mk8m
jPazDJIlSjNANV1oPwOqR7S1gRJkgXmYcbioHSDd8oLefM04xc1dWHKzN2KjfFij
p3AeuHF6muwsYg/TgjEbJ+IYCZ6Ll1QpR3EoO+Z5UuD/atimVrtDRRY7wHzr71SC
vZL1T2wL33WNTDjHtbwC34vOGnb/V1r9SAY9z/NCKY1vWjNvMlPbfv8Eul2Aum5b
1SNeUnwcjncmdtNHMEmLU6YnKFHvMbYI3zPCMHx0nCn+DyUg7EeMgFqJkC2qdVWr
n4d3ulmSW5Ty/eSxCsbV6CAkRDd0z14jvFWgDJ3fzQBAWzt6YdyS09UN6PoZaQoB
dSL/OsZhenbqDOSvK841ZFfXqzWEmqN7/0ddjhOoOxaDfnOB7ASvMICkxYLboq2R
mQZpV8F0jS95M5psnFjMAOghB+i+W0iqQU86jvAGADTokHFMaeuhG8V8wbqXaCuB
zg+FGoOTrPDZ6bsqx37MEuBf7trg+IPKFxsHKFe6cY6htFYbHuzfR26O1lf2nNMD
7SRrW4xlDbJLQmA0KercDepX6Lynd/cKCAfkwrDc1Wzk0OwaFTdCxD1Gve5na09g
ReoOWPf+yLANfxvKeEzTLRbicLtSkmtlngtFrFtGTFSiMSX8YPRcBt/hhAMxyQmX
6m/g5ajXVgK/XBJc+eTuCirYjEVJHs5c+WrroHg5e6oAmiWhmtYz+MsS7whd+Sfe
6UP9GoFUha1I/6fEARwUSI1BMAg6kHrCdzXsOThI0Im+ngMZLH9RJyo2lFyv2khi
SE8nMoOQsd99h6uDZMDyqWDZuoNQdIEzeqm/2BFwaH/Poal5SM2Hqllbr81+QT/8
sQUlPYxbcBb4BGzul2OHsf96wVPzOrzYfG2HOouITL97fbsj+oiWIoV7fumGSmEV
eBAcFCaT5EG/8d/vOaqFLjpiVg1i+RgVsD6joE6uc4gvlB86e9TmwcHTNy6ZG+rU
HC5GaPwlEePN+Q/OPSh+8VN7+Q8w816+kpqNVmu0/EdTjrFxIP8Yerzx5YgUBGlM
/oRWg6FrDBpTotknOmy3f448gw2Rhd22zfnmqcN1VIITqyxcRoQhbzo7hZEOicLb
oKrErFfoa3KqBAO0+dk/9y/7CER7/3m5vUWfmYnyKTWIMcc1VE0/BDjCQmkqDv+G
aX3v/efGmMd0l4YQVWKxoyobcP9tKDJfeeoZxAQPzVWpFzGWZfrBx2OFcskdGl29
T/H7XuCQIRFy8GPGDynz/M7svivjxc5Yz1knn2DNsK3fOcWva7IOZLLPlIPEAsmX
D/wKsrbBJi0xN/G5q7uGtowJsagf2vDtlE1QcHoUNxnzptJ0e7oNz58PNacupmpr
adG+Ih0l1HYgcSPCvVUlaQKvCFhvK1qzLirtTiau3cO1s/BVk6ID6Omt/5I2tJae
BN/TuIlep3vB8e9zz9KU1YQLOSmv1TjJvvaJ9BU3vXOJxcyJIUubMGuDhd9ldC2n
SSTv325yhjW5HDXRgkYkEJ9zHMKTcFuHt430SH6HhII24cEKDK7Hrr6jyGYVRg1F
XAFGmEbHSBnMNk/DgtYkE3U8ZfsbyTCGC6CfuyASSf8eK5+jpqnILuwfNoZMgzuj
wVZ7TXic84pO5A0rGAYrySzY/qwKk6R56Nd1/WBXQZDDLRLq6qWZ6rQYktscgElm
BcIUuubz52a+R7WgrkkL5vbMDYmRhj1YZ+3RBeEqRgs=
`protect END_PROTECTED
