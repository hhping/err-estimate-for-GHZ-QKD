`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjYMmkKx80Y1hiA2///14txe7ABpz+vxscfKAoznTDNr2ldO14aYTxow13R3A1jX
U7YSc/+dUcJQWXGZ0CVc9NOo4EKmUWQX3s+aDfIIjIDNHRl3/KPkYZjbXUvhxnhB
8cWJytquYbwtA8mlsFgLb29o09CHywuKdaMQh5vfwHe1gI/4ThouQ2IgSIxQPK0I
D8m2Zl79zc1kReP/PYc3X8qUuYcc7uyRBQdg6sXqDg+3KeA0IaOUmlYrF/HliJMm
o/pVVd61LrCv0sEFkpsnrvle73bhCX724l4V0LzEJOJQ04GxeTfgVIX8BIUdFTaf
o/361nYjnb4K58RIu18+xcd53VaNMwNKuotV3F0iY0c8V2bnrxknp+OpNzIGng9r
kWhVDXubJcjNeA4euu9nolL9N0oIbwFrKJ6KD7rj3ytU4i0UqRWmh6iECd+FURt8
x4CdqvvJhw207nnge3/P3PwLW2FmtxvA0yFTrsDzm/yX6gpecsdRbSIRCH5tpxap
hH3pmTt4Vs22B/zY3ZFjp5AIxsiCwJEaM6RuXrfAG9Lxr8phsuvBHahj/XVuFplU
3ccKWTu9jiSvVy73XbKYFPY3QO8KQeDGYVqv1nmqmya3ybadqpCsFJc1SKzegTTq
4G+0i89dT+SMGBoWQRRHXwKXTgi5a7WIANu+CKZ/1Y64jn1X9vIn6+7O63pCeec9
IwegFIJS07jTz0eqb8aEqd5pLRBigZlrdBTbG0paBcrEfAOQ2fTX9L/V5bAclMky
GJ3kzr+VdGzDLMo6qjdk8H+MyCnD2HJnUpS5/p6LHI9en/+SgkyX5KFosF2zagbE
eBRJbgSt4vs0uusfEtW0EvXxHHFzXq/kON57ohGS9t6A0fH4YFX47FnPyhzT5C0k
qkLimR86hTgqNoWiOULZ2gNj9YyPj9lU7cp7trRbSwrYJ7j0WM9TVxV0LrUnLBLk
8/VnA+tmbONsrKBOH+MYpx3Qw81DJpZl4zxC8iU92rSgqquUXEn2D01IaaT6rZcF
16UL6eFWPhTF+UKRd12Fe6nPJogT1Q95kFVGbZJBd1bTScrzlMYEe+UIT0AXOt3E
rhPSjx86FVWUQGZwfsSMIA4OPb1CqRSxQe0u1Lv03lx96/QTs3HqNnWk4mlNkpiL
3fXMRiKxmf19HGkQA5R/WCMUhBxs2R52/4SY7SxzuQ9fiX8W0BazeHUO3daMRp4F
mPnj4f2i08jQtpjw3XyDdb2B4F5NghSR5vJ9YMeLSLfMdrclJxEo92JCBjgPGgJq
W+n/3JLj1DRIFQe8ll8C1tpeHndLmFprqfsilcosTtBT+wjoiD2dbDeVkxjyHFPS
Z7xtttoU+quBQcOHGDmhDmKp+8K49yc8gwls+ChTlZTuHm1PNlb8MXPSPEMdg0I8
zLx6qFsB1dCOepfjNCETtbemjHCEiZNUYPUcxqsNvGm+tYhDh9C0UBYPcr4T+jWp
imNrTlPKWmgIrNgh6CGbuzZFbMCaVthymjsSMN8QylFO4srzKFynfiEpy3xZuGF0
Wz8KNyM6T9BLPHVZxPziwtB0ZAOiMy61xCsgYFK2WYtsPckuSaOnnz7Pmm6Uaquq
NPZQsAeO5/vR7Md5ZdEW/TquXIKAYo8q+42CEUu5kxHJLC1Gxr5TYEyZVW9ztfee
VXKqqqfWYvPNirOLKUPrC7GTiTZOqlcJ08+kSXCeahidhoupr/JHl0vkwJQWWUtm
/tvwOPf4FuPN743Yoi60cHF1XT1yrQVuKRxayUD/SdgUuec3MHDK2iTqEqSmwVb5
Xke83rWy9scVprkpZxhuc0/DUBZAgyvSMmyKjDb6i5RWOwWGo9TwpEMPdcOEaEwq
b4+gikgJ/etQWdUtRFKw/WdaUkKS+redl7Oa6FRAWEgNQl2TS6VcvDESSO0GHisO
7qjKBeQNoUhQL9H0FyouGC9h3F706Md2u4NK4zsd9EK0RS/hiG0ge4QBWr2bDP6p
m4k4Gxd9scIQzXAbK99YeHfL/cwUlN83xJBOhugrLRUzuDEtfTbfZ//8PAH+92EY
eNWBI5gS3/v0lEOaOjWu3ZbKxoHZwCfyDV4plmzYi/BI42O59sjO/yRzkvWZdW3a
dBR3JUUNen31QylScEKC0gG5mk7oiHONcKhlelhZIPh4Q8CIaGgCPA1NubE0c90E
iJFtmgZDMPrLwR3WusmiZuhbP95pE7qXcRu6KYBE3tmeAC+37c3xLnjjh1GtdIvn
yjLT11XfJ8BBagi/N7qNn/MMOjVOq0zi9M2RX9gVoxcmACeLIGAmHj4dsWe2usPZ
4OO3s9iMs/o9CIac+Pd/5Q==
`protect END_PROTECTED
