`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqAGm15X2rEzxbZxPM2rXW0bbRmt3+Mf2BOTNeg7VFXP9dGPsBpARYP5KzGZOrYr
f1hcHRJFYMIBl/2GI3BYIBJ0RZqh2x7IoMppg7fJ3+4azf4bDL4RgDxXzGuwMAhv
WI1dkDKou3M1ktKbTuQR68VLNtn9tVuxHC9VAegKpaZftDFklJ51wNVpRabFZXyI
oFC/t+Et2WOM9qbq5yXeWYNVFfeDuWvD/h7tgxJj6aJ/FfIQNfiJxRgtJ/LGUII+
n/pWeWoqXgIUDSPg4IlOoTq2VFtBVlpzDpG8ASVpY2xmqxTJ9dITptAQ5CJeGMZo
EEX3PCDF6ussKAJMstRoC/EOo8u1mq6Q64xhs7iAqSG/1lL4NyZe3LDbk55oCSY3
f35f1AW8fgxPMjTpPh5ZBH7yTgglimuVtk2Fncd+q5q1Sox23/KqYVOsGU3wkKyA
kawiV0oSfHFOe7L0lkbjOV4XGUPshuPQzlJ8JiQfzNoZKO2815jd6uDEq+v2z8GS
dYzG8VRe7Ai1gcRL9VrAyZ55mR/cd1MqzWfsiGa9JTY7yHf7dxG8Ic11Psnvxe4k
0g9aqUaFy1mBDeUE1PsvybXLSVQ1ydAkp5OkG7RfH/FMcFyYpkBilc6AioQg+QgB
41cmNdUj36vK26X++OUNZA2ATbErkfqIBf4rDxQszTv/tZ7bP4+4sbBsuHZobBEJ
wpIMwb3ca7dgsR9FkVYi2TryndZX12WIFM288Bo32JjUQfRXCWAvwEhgcAzh8isB
nYrfDBS4WdmubtMLT+tSEsGMHVJP1DjQKu8oJebe53kHEjd7IpZVh/psXLghU1l+
BGYqXBXy1zBT6UfJx97hagtLjji00J1J0i56yvuwfjfOLmJflvvlXHzWZcYvwfMC
hFbhs7VkHbhiStc0kNMwFeU82LIrCusAuQTf1yQxCzkRVIjdJKH8fOhqtxl6XgTe
P9Lyw9ehKIvfMd/IUXq7F1I0/SD02pxx9Zqo4xcL9yNH8lL0dmx8YQfMP57vXinw
Mjxw9XtvUOVkUGWSt4XT9LFjx5KQHI9tAbkxQIxAn2+c8FuRmFnbl/mgb+/V/oE8
+uTtZtIDg1IDuoQn5YfFmNQiOenkpgHJsnR7gcA4J/3Xw1yfMK7TkqUmI88xkzP4
1SIVnwOyluTMksN2kyRq59Pi0UAhnuDknSgAtbabr9Wo8eAKuwo/v13i5tJ1ScqZ
GCks4LJxIV05dfafHIiN4Xyt2d1R42uvAqdQMkJUIOILaQvNoIkEoqa9IVaBtFBN
seNXpHozzBS1mptf9TbVfNUFZe/i5IWv19vl1vdhocvTHjHR0ryNAXBeTiUOIMhi
B3M62QeQG7YTCKXHvPnvsHhEZHzCEKRIGvK/mVRuwv13h4FBaC0v+6FIABez/d7M
HxNJ1IK7c1XY0O8SrmhWI/ldbMTVE6fPQ66FgiEm1hoWPsm2IYqfQLVMvtgLXt3c
AlUfjzSBhQdjYUpxgmnCRaZgBwVMV0132+ocWzNeQgxctLNVI1axT9mgAWr/w0AZ
Ab8/73Kch4WtKlJvjEsjImTI5ls6BRJEtmmCxhWj/Gc0P5bcZ98K/9kydDfRvQT8
Sn8z4VKN37ri+bhQw2TZ4yWa8cSbE1mzJ9tDxLzmzRPGyrWjHxRjI7Nny/i3NyLG
I1G3bp/9kxlMakgX3Yux51d14Gq9VULeOaK987ixOqRHYLCTF5deo/RuAPx+HKgB
zpehouVn8lM55kDu0FHLWQLyLOqcJ7dfoxjywMAjBZApXdMrUvhkbMBAf7rZ/i3T
RPjdxJTK4EDfPr0Cpu5jZqVi8sy4qqU2r6UvS9oYW/i1E7SqfPEgCZe2qAT3CnB4
zM6hDxRqt53NZsXedUJN480z3GvNvpJub5Rs/dcNPvgOXuhZZ8s4oXBwYjKg0X1t
3q036kUH4OMkPaYOxAdqUt0Jub6IzaCZ/y8IERhpVncAePxdpIAFvvQ1DmGPl/vv
APZ5tW8arBqoBzO+GI8WX9OIatIvUpPayD17HLNxls1r/N7h6uRQRTIRzM2LN92w
56e0bxUnDqnuWsbhPkNssuSg8ObOSIbixKfsKTMeudA+NoAvA2dhvwAN/VHLUpLM
gTvFw2rIh2hR3+j8bfiREZS89H39ICYkQw8uzu41lUeKguJDpHHs8FcxO21Vfk3+
N0UMkxASstfPlGoqw6kUyBAG89HBrVJ2u9Ubj6yeTYM1jmN7UvXYtz+07z0l3+2N
6Vkul7Cy3Ze/81gs8KCYSJuv/Wa04oWlkgmrTRUx8XzCgfeHQ6T3UXuJ6/gwyo8p
7ZtIcnI/fcyfKTWGyobscvs1pYWoZNq5G1glluDuP7cLzHCiNSdqB6r+wov3/uZR
DmyAsTs6p2bkmRo6WaD1OvpUjLihGWT9AXWZORDx5Wn1YkC7BFNSJkeiTSDTCCNO
bkimiLC0IcVM0Gm7xbfjODh17+12HMtJmoLAPBX3PA9CIZP+GHJc3vMxnmef4GeR
epdVlWJ8NIlMIMHMCLU+S3obwj+orszecy6LM4zrCKyw/r8WZiyMsBv2e3A6TsBv
rQHkDYdhd6xxJOR+r8gRmiKWOVoXRTA1tTFqo2X0MW3uFYeOGbLOQBlcm4Zi1hQH
hM4YE0cJWcMySTbLFNMMTiftX8RW33EJmUq9IJIwyFzeFN9wX1C/To8MR3qZbrhG
BqRx2hS3y7NpFGQuh0SFwbGOONOmSTe12PKJgTSdulnA83aH9bMHDdC7tfHek3YC
xWsZlKl/ggW6aejOhe6KGoTkLV+huqwjhxjkEFkh7X5wstoLG8bwP8KGf+uXY7ae
qqWBkm53oUdGiw7N9f+xK5fkjJjSsX7zh9yfl53qVWdDQllEBOoZ5sUlvGFwPJbc
nk0gV8IIsm4CDmADZfZp6+QglTtGd88IbT7qUW2l7TifdtOS8LZgdcv/HYz6o22r
OY+df+PV1qucoI2iaY1yjXoQhP+v7NtISMWFYMDgdwtmguaTT0t9phZoKp8t43ZY
qJLw3BsnDD9R4OO/CbNZ5byFMsf+/yNeTaeGVrX3PdXux91EO8OPLoF1k1Yw2yEJ
wdzxlzc92TvECgqqLKtJ4hy5c3kctbN4kwgj9ew9kesDp7f+xRrhXQ6yAnQdnICu
iqgsyJ/RU2ID2gYPzCItPgcED2wXsVh9Gug58/lyrrjHPiiSLQdY+Da0MBBaA37L
7+9ZL4TAL6PEPR8SLfpJqFioJl5K8B//iDzTs8GTxh8EQLDMIZLnLXhIW+1F1iHq
EGSWOOVazP4V1IGSrmHpRep11Qk9rztcN8EpALbDoXo9R0cwS1wYO2kFkys1Rlm8
toLnlBIIlSm14LdVgJgcBH75GwO3vWwNimKWj97G7O8JgOFxQRIMgQhcxf0yUcv6
dSpEHCL0A850eon4wplnxE5OEdRFv6Pi0FPe35rY3I5EbBCEQZJrCkZzTECJmDBN
4gs2KrZFalpSlGFtgLQsHS8ADInahc52U+5ocl2Jv4/J+/xP4RwUy6py3wOW1Gqg
bQYT/QBV+CG/DrvNGnVnzXLax3COgkfwPTJzFNlqyP/rB0v+y9XdRR9khpBDKPQk
UHUFej+lNoRf040L+UPQ7lgjWGlvyjCXmj3PoDd0e5g/9eK+GF6JS5mqg93h17WT
lqxcErGJvDFAR+4rPEv5LKc7PFK3V/7OrW+HLZYsSz/9LLJcOCOGrsBiSqSOJWrn
4UgjteKMQuAP/deUhWoW6+PgS5d+niCEAOhNaBZdqGlfXUCznqZV7WIo9d6JdEGz
gLEqmHJhFizjeqCEqRpEnu+IZKoam5S/LRSRM6Vyg98Xb/wLfy/U+1xQiTqfWig7
1234unjIcS0DWBNNoqpKR973+Q2J/n+iC3yw3xANs4XRD8VZ5ElrDtW2ARJvSlkM
c09ea2r/MPCZkfic51aJFH4+fkW5GeUzPC5c+rIR9aw7SGUNxOUT+30d5njqQ7mm
`protect END_PROTECTED
