`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LuIjv6b6pKvYRUeSwC3QdPa9yIDbOU7S5RIJ4SlC/O3d7tGub0Rgd/jw1d7aNaeK
P/pGB9fy5ogfXisl2bbS0kd91x1EscH6UsfL8xEAc+HQqGtJvVpSamOO+QMPamB0
MfV/E6AwAJGzwe86QgcnJ62tDH2zwMOHfAZMVQcsqc0DnvCo33FgAfa7Cr1/AOkl
e0f7Y13OXikmqYqqyK0I+6lsx8+IG7IBSXgZAJ+Q6CJOSOdHa0gDMnWw6g5PHSqI
irJIFBKWQO3JCR/8ne8pJbNGlzx+vVw89HO/7b9+c9wtGcgyii44aw8+yifUNveR
iTgL72rCK6Q/+0E19ntuwpUjwFauTEBtUqXr7i3qqIfIPsA4Yxrr8z4zM4bHnv0h
/3yBGV+Uj3qo8VtcRw/VYFagCWUE04YGB4jmxtXx1xli+GoS6RhlEG+hMumb+5Ue
SXFhY0KtYB1ichEBKH1CDy3A2uw9E7CbwX0tNufNwM8wGB9nAjBikImCKZB3H1tn
J725ozBw09RfOJ5+jSrXrzfS6EgpNpffjNxITfs3EhICOheyC9LOZUxZmGtZncxc
dcJ3IxEjPoFSDCG/tWEXZfqbyVzwAO2xvzWBctG8Wsu76QrNfC79X8VTfQFhQ6y3
KOVCO9OeRPYavDxvySjlB9akiNXRt2xcwSL1/yoZ4WJxo4gw/64sT9LueWFfvSmr
HQoe8jI87XeQq1orTa7zEv07l1xzcA2ZRARIPpJS6DU3Wq99Fg4oSPUr7nbXRqqQ
cQfrpsGTxc61ca29AU5AN/TrSZdI95s1b3ehZl0/ULrME1/j9yO+vqbsmob1vCaD
YM9y241cV2tMSqpwau4NOKRkhWBcFQnSk901f1M4ygp5NvLhevzNE7I/5182maeF
SmdhTC8c0Eius20rYcdUa9o0idNGajyL4y+59BIqC0GloPiYUwmsIITVCUBHmeJ1
CFHPsCRiRgv819B6vjwTYH/cwS/h/CeYtgLKWSBT7mfRAzm/ZhxExKu/0O0SBVDM
o3H62JKqtmnVxW45hWAgxuqIxAr1wNOEhA0WCvAX/gosIs2yHPF6fMarIFNXXo4b
9TnMBsFcfRNtohFSKG0nCw==
`protect END_PROTECTED
