`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2VInUNk3Sejgt90H9pX8qHPfOVMLHC5gUqwOyNW7il0SC7/va0xa+/+eTol1uzM
HrkOX6iLyJa6M8NLkLzq4jVe5AVuufMg6amyGDNT8NtOLz0wndgJA7035dmk6Zg6
a6zSGfbCqi0V5vRscHehJJ1pUS8y9MJDLak35Tvaqqa5bPoh1YDsJyJTh7JRXLAv
X1XC98Ep2Hiaks/YCD+bQIOjUbYg+S6vytCcfYrtGkmghRDxcKGnDv7HUvAzrtFl
JUKMiLmjPlGMlRm5nbvg6SIk1eSWJpQbLRo6VfD93mUaN8WClZ24bKRQoPwnSKQs
KOu8kXsCVUCXQYbjJUrpHKo0mDwvjeD0aWoAVgX8UWD7gufboRHKS9ji1HMPmXup
GN0vsrAULyyK5cwe4VggFZlP185SDnnZ409XS6k4gQETm4eNumrzNFo0mPNa+rll
5pwV8chK5nCHgnCFZ2kic5/0vyKv1Ckte40cgfX+JY8XqekjSpfqLWjitUL7We6I
sQfpjXLnx0Da6Mt7lAumiqcjSjM0H7eBtB2UqSedmRHabsutYNfAve2Jc//0HVbF
SQfzoisZnyGaoqJHd7sSjuAuv7raK9ScqNTWdsyQey4IinB8L7+/yWyR5EVbVmML
H58aH2QXh/aiF/2ay43mME5Fl4rvTG/5Nq84JKBHu3rI//dVaviNyn1Celh/7sZC
eelx9lwnr/Lrz94POlF0lTKDYbjZ+zMsLMJpCOse9etOXckrK84hF5PPA1zxe/Xp
x6BRnzHpK9fmD+Z2RGjOdgHN0GOswy9lo4/yT1Y9xyYnI2V7Csyrcuh05EWOUG5Y
wjiLx5rsI8d02sphdZNORlLp9Qm8pwT1Js4Cw/K8iHxU9YXXLijLDi5gqCGOa4oo
ivah4zKEsuF5zY13Pi8KkQ3UYtsHi/g/0Au1pY4K767YxftpgIHDfSMTTfs+j9XH
zs3vVY2JWz/NqhtQ3cWzG8SX8psHBoS09V2qYsVnIubcPOg4XIW6NC4peitlQDJ2
v4CvHpHRfM/PspIYz0Xj02n87o3FvLyHqtlyZli7MPVoo4msPSzuwyn62xncNcp6
Pf5AMx3kAxefCAOmD6g7bxeITmDQdfHB7nrniU/dq9Ox3uYhsxOLVPzqG3sblsOM
QV86CmmnI+mNROzbNN2Uoe8WueUSjzr0r+9QvZngm2sMQG2HPMmT8o2aevu6kQdK
fZDbWmMwN6Rpz9ghlGBeBGn4by/PqE9fZmvp8dCB0NrSxy+Pw5fp8HAtPNNemUYi
VOLbXE4m6GXISDl2wYBOtKVLM4oYQgXWSFdwWzoUarrcglDgmcdyMFymeQKFbQ0L
m6vib/jlYgWq4PsNiDdwLuitleRk1r8HjQToUKBHxuzAHmU2qV4zCg0Nlm3KrtlL
Qk4r4biIZPV/8JGsdEwpwJinj1T7DQ2iJWPo9wCfcJCbOFiGkWroy0qAh7ZGO9t6
swf9GeNdb1XZQucym4R63FUknkZVI0bJLScEgrqqxNjeu6wEfdgHt32VgP6hMgl+
nEfrDocAVC3SiLZHTXU1CfvHCttH0ilb4uTo10627+fXXppz0GcgyRqEqa5QNp3x
2jT70eNT0YDlkXK688e+5neccuPXcQg59+QAEZReZ+bxAiPjY8u77DEQpnK8jJeA
PAOH5x4/aPVlXY6D06G/2DlT54Lx+gKl6A6fe6IowkXzRJFlUwzBiBo+TU8ZZ0DA
UAT8RNk6xZosxz3zh3gWmD6IyvClBQq8x6EZBkacAszpAg3KPWUO2yeEptkIhA8h
71j9UwQuidenXYylpRzljtdm3InupmY6C15q+iiKxkpG68ZLP4QBU83vzyqmQ1NE
`protect END_PROTECTED
