`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vPA4LFsuSmLNw08qa0qU0h2q40ewSXthO7XR+pzuEUgM/mNiB0szTu0Jbt9+hdSk
UjSdeuNea+PDQ58xiYr0va30fAbS4fasBwkui3KA3XXu6CjXqZ+KN+cdZyn0Tjfd
WPT9cDGFHIdiEnCwbmppe7JeQeB3dvzdvtWQE8ljYNfak8DZou8WQQSBsbXEA6jM
Mxvg1h707illN+NrGwrXKN4wrGIgAYT1E0mjQlwSenhjTeEENhi7i7dBwGNaO+Iq
opItij2m1pwNaSmJcyy3zUbWgq95g+Xp41JwN2UWS4Ek7+uhIRJeePUsznJB5hAl
IqSo7uBtBIDGHdgVrjchiTP0EKXxqkqIrg8+/Vbsu9kMojrt7NdUQ6aLgzltXBJB
pP+4i3EPkTbv3rnrH+uz+gtFpfDbjkc4UEBETwlVZeIpPZWqRSkbTPh8sSRNKabb
KdyEdj2BxfcuGSfNe8RGCDiKhfg4Rq01LRAG64dP0+E4CszzRMLKaytZfDS4Quc8
NvQoux4zDkEBojOZQcmlJwadb3/CGAyBjipJz8TUmiv7W0c2zwGgbONgQ+ZHm63H
YkKy154Vz5ZxTZxSxQif02kkbiOTgEvl37o9MVbRJRYaXICNtRFEpsPSuKqMUX3X
ZXMaNLxaZbmh04pF7nTRzx0ijty2eoR9IAT0XRXmWkA1lCCMgWJ3p5vSJg3aQ+6Z
G+pd360kRXdZYJ9fg7pJBQWAMyf1ShfP1UzW1MbKuDppITMIumMsPn3ioR3wqmWV
0F0MPjLblMwa+lCusO/VyhEMIMCHdujxH27XQVB7+maDLQUKUquBFw6HLz/VUJSG
e79mXOtKnLxsWXTs8pO1Ve422fNGuykfUrKCIZxZ1mTP8LKyeRtiRnEPGY1jKPVo
IeBcMZIZBefuiTufQp7gK7iRUt/nx4vjEKX6P77rNO5SZz0+tyXYhHs0jmiAwJ2g
juVj99RmMp/Zu/VhTw/1WG3E2T2Nj79OW9uFLwoQbpSymvnHLwcEeSlXllokE2sg
`protect END_PROTECTED
