`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogFf6cOWetUwRMJ9rbxjdGn8NnhwRQd+lEb25XJ0PgsInZBTZ1sr0wsoupee+V7Y
AH9s3YyiaCzbylk5kIeeSrMbDIQ1jL2tMf9L0MyphDGPV0jR497iHw2ugCwXuZ6e
FZ1zqfRoK+tO+ee/pgkTmIWDP7G/LBW1bA6Fjsf16BDwMuX20CfxojVfNP/aCyB0
/O9du3WYySMqTrqqQVbyBrbsAQSJMwwJUEOpGNMomspauIvWrbRhO3JgWf/ruHyx
4eRWC99R+sH1vLTlf1IQMbLVugC+KZOezMhFmCGg5l4FDp3u+WxihZKfreW4AYS+
PARWJEsIbSJWi80Y9b7sfprkrZ7cfw2+Jya8RHgCi6Owi+3QaVg5y+7BsY0IrRMN
1qX8rCfD4y7waAjDtN/duKf5N1sd2LDI4d/sK9R++u2vnerUqTKTbbJWmuDEt5to
SXsAH8epVVjqEPcdTHXH/ptKdN1Qz4ViURGVfsuzBFrkYnB4/yQz6P/u0o1GkPo5
LIpID6c8LYM5gjSk8dXqOIJoJyNJ0NF2MPplZ5YXHEs/RVzMB+pyx6VEteWO2s+l
FzsyTx9+q3eFqgjUa/4V/SctZxQEgcdt6ykw8kVocgtVT40tX8ScT5o6yBz69Ilh
LEfgbqv89JvFX0J6tdhErT7zLnkbI5cL/H3qiG96ri408Anqmk1Wnjo8BHdGNct0
fqn4n5KhbxET5XNfPKo9zgp6+inp2EUYRsLls5eKpvbXWQ2pCOJk/pIP9pCnPRIO
cFEU1ZvfTai6VQ5+n9A+isUVSESMBdX43ChqzkXpwX5aHuh2pecS/CIjXNmwO/Fu
B0FlMk4eJsTdgP5RheXSueD05jruhem6ozFjobehYx/295v3itwjBG77M1/N8r28
IFdMadjZCzOlI52Nd7Xf71PtFpV2wvR4K5EhthWZukrbdiAnwsx0bMsjncEprL99
tBBV94e29QfXd/gPxCuIAQwwQ6hUM6UAyO0g98hDqUmXqjKd7S+1i5DiXS+GOEf4
YgcYvAKk1Ykg+pAfoOK9rKFknRkzjfqTo2YBIQCi012ZR/KQH3ZKH1fsbnTRgOSY
1jAlQ6mWP0wyqhVoq9P8Jij75aYBTaEyPU4yJ9JJ+tz1L1hHFthQiMKekvNrZcYV
FMZU5w1lFtPeqWKNoqSpJvURbjy0bajBaKtxfFvzPCBhU3TWFIJVuEAz6rA3sBHj
Lbt0iMN4p1pM2ih0f/a3O6+hKd6DxP08scFo6r5KkGQPPI0q0e3FiHrAFp9uVlPO
VDxZcJiSbAqdCe10tfBCHphhimmkaNskrsqGQfu3Tla7gQXGw7JQeN4n0BQQfok9
`protect END_PROTECTED
