`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZO4KLdfKFdvUVK+zeKt0G+V/Gesj7fkzROJF3C/4TwcEpZ9/kQVPAes21ICotr8
lG6ebFU7UpAyXFaMO3USqYdcBaPRnYzfxfHXfHdPNJ0O/uyYPkBbR8V3diyFfD06
qythfFJqS68PFYSLQg5b2Za0vyMzKy0tzGjGw6c0tgH4Yhv4h0nlR7HkEyF3UGPk
d/GY8pbraLTjNzqaaNdj87goVwG3hb62dHzMKpe2OEeE6ADWzPMConbJqvipadCl
PlpVLrBBeYGAb/yfXt1ZCw4hYPxI/UDNPfAcASs2hiFRENujnHoregS9DA5NhvSa
3rjZgCyupkk7jF5HQp7umAorzo5lI0qNrPJoC6RW0MlAXLGfVlObOx+fK3YjlYtH
ghypNseBai0qFpLYqIIn6SpJXQyQqXGxP9G/50lk5SJjZQa8ubO6TTJSAWFtMJBO
d2m3+7ipQpcnssHgbPOBnQIDdnuEk7JFHAlHi1R5I8vbfptO2Vf0sMUmUk3Z1l6C
5dcIKl751QgecS8rbMpnMxQAWh6dMXwGREz/bzkgkIMP4qo6kRh4jnbyrr1DO2bO
GUr/qSKmEhZM44AhzQ8JOA+sQ//z5YnCoTmmPqhCuomdUeST81IB1hEOPRaoerya
Vho4dYZKcH6GVZOPSjC3UXmy84Qh6Vyp2stYZVg8w+OKQX7hQ8Cn3tPa7N9bSLMO
nHyz7j4d6uGjBRK0o0y3PIzAHhHONtjmEOlYtn8OolLVXoOFf59jRKsRdzktZLBd
20S6LogXYfkd9+5V0u5fhwuX4IU88oEurq1QgP18UNfCA8zIzepQimJCAXGQL7/Z
EBtAdyuSyhWomjZchpd/P4VfdJXcUDLZeUsL5tEm/Mh95pYz9oDQ9UTWgUSzWhML
dh6C0b7X0UmdszDyoUpN3B61PDAstkjo+8bdsZhRqx2r1Kn3Njex+LDABlTmQjmT
m2fSMpvoOtA3aCs/EjNqW6+bEOvZMeNK5MOla9mlL2KVVqCd074jk+zZ9HX5s+od
Lxxgx5vw6aS+SMRCuIGdle75Lq5DRHNR+snJ9oZr/wMx1SIP1gJELFWlGJLmMpQR
U2kD6a4tGmLz8tdpNAU5577UDXnV6TGaG7gJ7BW8M8OwcmTB0x3pN6OIq9E5INhy
6q7vVIOT1U6238Kp3hznGWXaHRUAxHS3S2INJz2MSLaabs0EQd3UYmN2X4IAFS5o
Y1hy3So2WsddphcLbyCM+B8Yvwj4IumV9eLXeP5D8CVlG4/v0iDEJ0dBPpk6jkn8
7/eea258Cg/lY1/u5UvpMVXF0oS7xJfXbjZ5LFePv/NOXT+QadZ4un+JCjvy4oGn
ZiuHV9fG7Gc69Fgp3KLwmgKFSkAtsN9zvTtut3OD70Kc/xmgVE8iZj79CCnWxz2e
s58w8WOemPX3vPr5sO6BL1w47Tv+W5XeQfNY/SAExQmmDiXObfFcJfJUAhJIqTUy
gYXrvuM5XP/2dj+WNoquzpG5LZ2C8SAkzYZLIf58hRSecAq6dH/qcMRy1mOI2JGU
8cPoHW2W+cO4jSulbsub5FehdQbXm461tyfrIamMIopeF+4Q9/KuVqGyVdx9aede
wotr9nOoJzinBYR1LYzgsauW833zXVkRT944tAjs93/U8Fx8Kox1YfPHrT+qD4iX
cX01JO/Ua7cat94DOwtyc5q+YhkQLNiKMsXS2qCMWMGwgev41YtF9FLzuz4Z7oOc
xhJWQZBfH6i6orVD7NNV/4vM43ApL2k0reYOryAfUEyrlR9WR/SSj+YUGnjLlYvH
oDZpeD6sO5wCkD0oNAsKh9fXJuKm4RRW7Ib1yt8pdDf6aPLf8/ytL2Vfp4NbIimU
05+8NHge1JlKnT/PgM1fCB+ywA4TVRcMzQehyBRGOpY=
`protect END_PROTECTED
