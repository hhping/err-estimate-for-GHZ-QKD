`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBhRjQf37ozu+pyYulN6zcv/Bnb+8hYMEKlduYIuw/7t7I6h9NiRHvwxsl0g2dp2
wVFWL7opeAPgAj3/ePO4I4cr8RVnXRBzS/I4NyDbcw70HWqxjfMMB598i5jD/1n8
WT00fWiLuVtQ4dwam7UpBhMBIT73Wot+RtCWeCIHlqE+6rzsWTorvG+JNQXWMsfD
AWY0GB/oHvNMgJUWhSDQ7o+vj+/WtMeUHqIxM5vVH8qsb74IqVNsUmD9gQhXTjKW
uXPfHSVJC+D0B5lqqRkJl+JAK37t4ksqQyT8ojSzuFaLCOjIsQ6IqrWWze4TCj7A
4Zv9AZ7e/lYpIkKJNcChNV7SS0dUTlFmrImYYJM1ulguvBMWt92z1Vl47bMX7qpZ
bPHQDmbA417c7IuN/L1tzEZuleehbiRroeGWhe+2Mh+u+nm6yuV8SRHY07KC72dR
AMTb2to0mJjaqJMf1jO8cwnz4WY6Ij03ERfU9npT4HdKCqUcKIbqo8iifqYvacfc
jFmQ/dNVTn6g1olkkW4pp1sqUVDUkJ620+tR1SQsSm5nA2kXNHDjTOkY6hW/OzMx
GLCWtYaxepK2KqqsnojmVb94J+BvPA2jzcTLdLJOZnVWlEXhrnkZN6+8IwNwh6Qz
5ZkPANxywcPGOJOlYx5zYBXBYRCJ1BK3ZnKfW9QFu1vQAyEqF6UG8eZprE+NI/vL
bw7QzTQua+NlcCU/XFBnU2q2Y180ED0X+hcEW6mR/XezYcAWcce/nRqfMQ5+di3A
I2neQiTyrLAzVc2NpyrYDFYIpWFRw3LeDWexSJJhFtMPePoB2isovQwF3HJKFFkR
IBlvIAw3mUSQkfS9Vsh0SY3NQudGA3a9fv6SzNj5ICQ=
`protect END_PROTECTED
