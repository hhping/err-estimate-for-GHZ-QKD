`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7uEpiAKPJPWZisw/uYm9ej4ONZVSgH7I7zTH74jZS8FqRN30PWKkCXnJRtnlGen
LQuKdoIQ+s0bsBtXJGSZI6Awf6cDV79PuYCrjYpc99QT4cRu8Ij9nbVsM/PlOoH3
g9tHV1GUOm+9OR78MK1rdNIO3PcfAHLUy8g3CWiecYEYxk5AOMPUUttfxHo4kJck
UzqImvLmyOLF6XiF8ojd+4N0K1vsJO20GS4AughGdn+E2A92vVr+CREpbVJLOtc9
hx5/eaYgwCS+q9qAjTW3GZX0JdRFfQ+FrDJ8R8Ga+P7ZwUBhGn/P/IZ0LPhOSS7X
SdpRrgxXNamnBL0zKHlFr7PkP+NtOopeTGuHEmR5ZA2Si2YL18zXuIL5HCyuYiWM
s+MSALvs05xRJJGAoy6egUNNiVJVvTcEyMHXBXgpvHb3pXwKDWfbRrLSt2aCnde7
N3ny1Jd9QQQRSh7oinArVegxaLWvIaO/9Mt+0bX0EbNS8NQoq/B877bC70hCBOy7
qDOt4wZX4XDKxdBYcV8DPlxAtcJciTkT2ttcBEZSv3sbdGpPfY6oOGy1EMQID0Aw
B45WyZVHl5WmgDJAm30nIkv+UltvVN82iWV7UFjz+0SH/IPC1yOoR2dC+nxEL4Hb
BK/WlEJKnXuQ8dH/DAXdKdCV4ijzG4ppr9w8D3yLhT6UCk+tevWmpuzfS6f/Qv15
BW9y9DO/hyfM8APoDKgT6Zs0c0erXfJVytbkPA/L3zSfDoWpvvLADP6EHaG0GbNl
R+jWw6tqAZdFQRQLX4aTQnFCxIo06nCq5kyiOv61WvAFBeIOYmDHoAhRuQXA4Rnu
mMPsmcm9UlywfwPqFIidxkhCjahkKn3OgTlEzLf5F0TkELZ//Dh4e8z9tWw2VRY8
QWq+xxseZMiVDTNJTeK2JFxrFTuNMkE5o+E7cfszKaXR3JwND2/zSNUv9HXkZBiH
r1UHZnGBc5WlBj7Sc30aDF0biEVzpjYCgx477HO1Ss87w1T6LgPcBTplrqQoULKa
Al/eSBAYNbJM8DzWNDxyfWH6DfdHE6cyg7yUG4/6ARROj66VyVSXfAq2aBFRlmoV
zOxX67ICTHXxuF1unYmTw6PMeYOTvY/ZDSRESZaSqPZFKE1q/PRjmP4/CFwffU/a
A6TG6GXfGharV9H94GFyqoSjFgzMZ2cQyY11bGq2swnwts0EZ0dC09R31clTVD4V
89fiCr+Y+XtuTea8igyraFytMelSkob2i0dQ2V4hsxQhSaR9AM15L1fEtq2hcWT2
AYRMB9jeSYSW966O8N6mbLEklnyssEeo/7UuPwddwG+TXspft79VZexceCglmIhv
jdOYl9hKQk0edOdkoJXKVCAztZN5dXS64cfN5UCI0g5zNeXfDD17y5gN8/ptnAIq
2f5HR+J+ekET6WruG+W1msTiT428TtvF0YIhMu33g6P2KzTpe9lKYFh7J3ujLHRR
fa/rwDef8hnUoRJaW+9T8skIvXse83ZTwJcjlXItOzkN0nJHC/0CeeMUGOHP0Qjz
TfjiQEGkpCOtD5YTqMgLyaFxgDOkeL+/H7bezC6/HvRmm/BzP5xe0iYrQmmmH4jd
`protect END_PROTECTED
