`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rE+U1cTUr4fU1JSpicyvYwlBiL6TDF0JK1KCNGlNr3q95jRqAvTMl8fktC/h4Hku
6TOJboU/zzTo7OLKxf+XtNvi0QEhyPC3NN0bT/HWiWo5HI4fvgrQZIan5ul1a5pT
XIxDhFJAT1rjXIqHC0cdkiqN0wt8siCZT1ou6Qm+0TF7OboLytAshUOuNQyJkolU
keGEqIYNS8yVFrVgHk10nAdPgjK+rrAlv8uF3vHYF7kpfQ0tc3eRncZhxnTs8Lul
DfCPwOwpE+USrzzCcSs7fhkRQ+Wms3KpxahZXP63JiIvixjU3rcbaoWf1DsUkJue
`protect END_PROTECTED
