`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeEwydyUrR5pFa5+1pDIRBAAUjm9H22IAshcYxxnoExodofx7qbquWVv4P6UjlWQ
OoyNUec5dQ6KWcNw0UY2nHv/Xpx2hfdJ7PyCGb+bUbKCMsIRzXt9xtDOJitDIVW8
cysR9KYDSbyEqf47X/D5NkwIKV0pZFagM47XY7Y8cbFaBbBNgvky3IXAmzPvEDNV
BgDmxbOzoPi7SeO39jfP+9VXToBdrdU/Crzs5rZx+2JvRbbQjyVzD6zokI8fmFml
DMicTohioZ9FrP+2n7lvS2UYOxn9XPKbAdzAUwZLM/+fR6CtxogaUvFkDFwlCOxp
dMKlIKZJHOv5nuNP5vJKNfS1mT2KgWZ+rLdPrv51a+gqDMcHXYX5JOaWcWMyFITi
V7jWFtpkXJRWmujqFw7XE9hrdth/57F93Mpahi7kGph9LzLSIqX3f3C7xv0rMCzn
t6LZW3PNWckYqU8FTWkFONDjBfNqdS3q7mooFDaM+5972SWf19tRKICwrty4BLjw
RUoHOR9ToW9k3lNxgD9wlx4x6zJnH7WJFblvbrzL6zkNDta55cbiLb5rlzoWzWwu
jTXQEFQcB4SJ/bDU5CII2fEsCJZOVPrnpxTkE2RvvcWxGWHt4uJYujT6Sy063nx0
oBweXe54gU0nLgqryxF/iZmd3HTA2Nvq1XQ1S0ZZ3NASGTYUPNPXpfEperaSmyZs
FQlWhwSIOxHnVHCKO191hs6YwyC/gIpZWe8u8NMTsdqify3uBi1FyopMEUYVV6ia
bjTkNDFnIyO1uM4Vws3K5YfL0f6GgLmVel6Z1k2LJCJdZ35IHzG3wYumxlftJxNZ
ixMrCm8yJU2f8GhYMWjMJS7dMIQWTlBat++krKOcVsFkJL8x/ACzqtetYeXmxr4r
fdCIAxIiBeYFTzsEUKVC0EQC3fgzizFb6iKs1U2Jrg7od0/1/MzgVIGh+ZhUkisZ
BzFolYORIbmB/RPT+uESs+b7OWZWcp9kFKoaimaBWODaSpWxfwTRB8zpxQbzUUMh
W3KN3I3jdKvHN2mMG9Amc2d4oaFW/Sh9R6TIIRaI4O+vTR3J9dXTQDS7DMTDKIaU
YTU09BDKZz4n1SkkaWknbEKt21NZDhJHYJ/evVjLpgXzMV6QfFWE7GnC8WzZS0ue
oL1y7d3NJaCfI/ENCnRX+d2k+YLVQDUOW+fu2gRkAU8G61F2TYs3Fyd6LL5ur/fJ
Z0OeAGz8RyWcR2bp7TiM6+KtWcA0SFr22xomAlt9AUN4oGGPPRdRjcMARt8eAb+p
bEOdMmmsrwfC0yP6qz84y7CDb8J6N0szrK5bzQS02Hwu+0QYs+JR+eGq6Qz+IO2l
IiIAte5XluZNtCTaEoQhuakQf6JfSRRhKMFBQ7DDqLc5K6gmFeia5H5jf4GiIEps
D7I3oG5alVECStzYdN8nCAu5MIFWKvXr//VzHLCl4WMd89X6oWGjk8DUq8BPBAuh
3+eFLmgQjOobF83a5PPnuPLRSq4P17uk+2nJIHPtgt0OrP9Q2nD4wp2gMxfajsxw
eMYqQEzde0Jj3Jx+MXiX0d5Cyb+Rd+VbKwW62AWfmns7bqXw0IDCp7omH/nyma4n
KVRTGqdYo+4eOK2OqykYiGC7m2ZEEw3B/O94aAR2fJuB72RAWyrHvRk8LK9QCc1b
gMBQu7TYxrN9rEA87c1Ba6PFLZ6Bdmt1/PMRgCYokqQHDNeQ+XjBfJOGZ5IlhgNx
u0AuCUjvWrxVNNlCt8yr7KIwUHQJM4a5oWQNnAGZerIHc3Uazi5398dg5J1rK3IA
FMI4ywmoRTi/ah/aYK+qEfMdl+Q5t2s00iYPta47e2Ll9d4OElZGXIe4AUZxixwG
SXGboTJwKlo+6I10gKFXd8qKfTuq3muuSzCEksjK/UDakw8MHtJLgw93/DGdAI9q
JjLmfRJVGQ5+1yHFwWh3jwGmpKnkfhZ42NWBqh8JIvOTH9Y6xwb4ZTq3/1iZEcvd
oRqreZ2vxHUgBJddlN1xHNyiO0TMdxmLxyQnzOoRDmKhMY2VUsJc7dkjnvWcBOGl
NIRS+TcElw2cjVbc309KRTbAEMSQ2NLqiD8Q6+ECpmFGil3rjVR/I/Kai4m7DMET
4Bsg7soaDv0avhiqsaw/8uPNGtyeTRpCunai++FVGLWHr8laKRtFFdEUO2SGAjXl
9nuIHDjTs4FLWdziD/SutO9idfghOMKw6kI5qDC/Voj5F917v9Sg+7ANbm+3mzYr
YX6Jj3cN4/VaMR5KDeajaj3Sl3WdE7OapCf/F8IbyGEHZl+oaqi9PanV8EYqxr5Z
a2sI6H2XzMGUtQVcxlKrEXK6Y4y8HAlxN59pRQEf4CgcRqrQroeYm/yEaGzHcBMf
Sv3HV5O22y6hZYB78UCu7Zh4Yw+vzQMZsfidYxlc7FNj2cYbkzInVc39aPO5wLaP
82Lfxy7cHHIoUerNrgD0338B/p7LY0hwjvTJx6ErkwLNa28Eprwn4KgjSSncLYQ7
OdWO91PWsRgiLHfV+IHx7zDWx5qNBiKjy9Xjmr4PAzqbfQ9kdx2QoaUCFxmebf/s
g0SpjEJUrrA7fF8rSWQKVhqyZ7SLKoBpow2O+k+muuc/fCuy7UmHUxAbTm3mFF52
NwXQ6ZWHECGdGmNLtCdYcFqrTk9kxIhLRTUwvsadaj5I2B+dzGdQDpt6z9Q9yCGY
wBQFM0lvCaM1pg1hufdEKFc2oyqB6YSLWyQANIkZbqbLeiuaPVhz2EJmn35ccnVi
Pmv3R6roMlYAhA7YcyVHexv6DMzaHOl3DgtFxMUVhRE+1keFykBmaXB2Z0SrbTxF
TPu/eCHWlrVLph1tX0TumxoCdenZjboIl9gt68aGEeeNQEwseaiJ6FT4xjkWtXeR
QCgNhL0xcl337ORYqEvkhdcV7RVTUs+XOYtN83S2+VK65SqeWh2zbGiH19/z6L61
gZNgY6bBHYidbI+idWp4tmM/mbDPTkRqYsLvm4+m8YbXDZ+YIy7IcXCj4O1qTFV9
Ez08g0EeikitHu0h54xWOGN2DrkTpA3jRNpmUHz+xBU2YOecc5gvVWRc5HKBG5IZ
Sw31cNm07w8btJ5omDi0pa8bpuRchNbtFn1zxl0dmmdAFBpwE/4Ox3nrn078C4/E
hHkephCw6EzB7J8TdPb1qh+KaPqrl4nqtnpXl4EWKREvXGJRLeGnKuILaGmKgslW
Zm+duNd8E6Yad1wiMEbRD4BMWsedx9JK8d2iuMiOE5Q9AyoISwXDkVOwv9sjtKnR
Xrm+cf3JFpUnWizJSv1oa+Ococ3dSsjo0U3ieJags56knAchb7eGb2jZYuCUV5Ci
0wiFBwutGSvaslXeHYu3d95Tkqsjih+3uu9WfLUZp8reS8VIIN+AMHEp84PgaexA
u/3Ko+ZM3SmmcAH2YfXtNmYZu0mql6dqkOtdJSLY/J7csRY4hqxkqCHOOtIoaGqy
TfSf4nW8fJSnRD0W8Xo6PaGVTz8glvGU5KkcJfvew7aIfU1CIXu1HbzAFjQ+sEjL
0PJyP9Up8ZNzVlf2cBTy7cfzgOBuL3NRxk11elb8Y2X6RcdgwsdpVjEJg/UOt4sm
PpupzW6YFAeEqQob8Ogwhyg6PMeQMl2mTC3TvhThPEyHul5lOazsZqBrt0ommLpK
nul2QNxY/yvC9HzvC7TLl/x31btHvMSoutjjC3RqSKpqja7h24JvBIV4TO2OTVV5
geNvEos/8wTJ9MglcgZ1JcNKhtNPu9sg6pkWaE4D9cSFj4kkQAvU2CkABqlsB0gW
lUO165/LcSXVU6rUUYuPIbXdJI6xJ0FpIw7Qm35iyIHQHE30LqU+fhiKcfGs/6FU
Q/rkfvWDMWmonLf6vB4gxiHbY0kkRipuaJHDsqRQ8JcRtsWvuHG7ru/tcs7olePq
y62DxTIMd20AYUuKFMo4WvASHNSsDBUtE30WOh5jqnHIhQRyTtyR7/Y45ME69eNh
tAo/xnVd6D5AkCyVH9RZVfnhLfOBcHXT89+8C9gQ8l2GyfZccSmV/cvdIuTatkxS
CarYyb6IvhaLwG+aQx1sP0KNlmnoU7iUcw/BjKa8+zj1GrzUcrB7/xmdS0oD9g6L
w2Wo38TUIgpiqnJ7r+PBbjyOZUO2Au9AgVrUxin9n3w1ABTBCFKUZENR+4txZzpw
ie+s0nsJ58rFSBHAOYeDYOCvM8eH8ukmoCuoxLaTEnRff8u/g17a8cpuggsWwTw0
nM9MPiP2Jk7jePeCd84qy19R3Lkschk1RJgAZesgr8909aYLOXi/pGUHdw/wd+WW
vmvk7NzsmOyE/QNuENreTL9lPbnAgNa8VDQE/VuTFnSu3+XqWjodDc09V30E5GKS
RqLg12xbHMAHiSr3aTKFpk3wt+xs+G/dtOvywcKcHhjyCzFitMq3EhIX4pZLL9yy
kGvAlzob2JxyIq3d/A7xaVlrSc/fJ9y7v9AZn/jdrgIGAjKLjmED/SXdWnE9c3FR
Tl7X6s9kCPbVglT4cDXkEU+Gui7+LpADpjqNL7Id2KHxfWJNVq0wXUWL182Nmlzq
eplWh0qoBtVib6CdEpHvAU9/r8XibHikrhlggZjVGtMhf2Xgd/Bo76CwXQR+HWAE
ZftScb1piw0OsUCszlZ93lpwNPl+xPRSxkJYSiSik54WU+CkF0gddZZXGAq0SYaV
FDg80sgknMQTtYImExc8jY0AY9VIQ7+rP5RL85saDnR/znguXQHrmJOfm5edHCVt
EAX6DsDq1v5fo5ua7O5lvxLu75ltS3DnJcfO4O6AQl4uorEZmIsPRiolSmr/V3HH
G/T4htIE0jdFjoXKKcp0MWFmlMMiHr60eCJ3G0w2Ed/ez9z3hbEI5hBEE7TSAJWq
+VAYkvD42zyfgtBRh7pGNRkUuDoaObKbKxGZOruyYmHUC7JaD0BNrtuErYYUT440
/Xc41Jnt5wrHT8Yz6zXOEYyHSy9kgKvxmNn6B90KOXXHQWVFTY4AN6oi/JJPtD7D
WVXB0qJ0XqFLdkG+Hzs2oUHK8IjlSje35gmRPTN4BrHp9w3Pa899nDh9B9/ThYhb
AKf2PCDD1c8KsVrBzOPQB8kd8rDDdyeO/TA1y4DHTIzxyWuls+KjIvgEUX+zLYjY
a6JLRx89lTkl976BRbyOXPsNCB5HOIHV+mE7o3nCM3fA8lRjcxLTcCEA5v51ASST
CoSiY5VbfhYB8DNy/BXX7l92g0/KIltGtJxYDPiMMQKiApGhF/j6z/JlIvL9eY+r
DYTJA+Zoewl4SO0++U1fLxK0kLjNURqUVca3Jwfhsnal2rW5Zd6EZBrqwDFAi96y
DUASbjgeMjAKtZ2SDszzIw6reoC3DlHFHOICg1FrAtHzuk3E4DA94o99uwgaw514
vOe8pD09guEY9tCvJUVO5MSO4bgfnvzUoh6qd3SoPiJGxnLX1+2Kb0hWcpDU7u21
EUDlfNFrV/pbdEkpFTOpSgeuPPctybSRLSTI2jfUwsh4Bjqrkrxz6epB2KzixJU+
d/9TLK5Gq8TNguZqUUQrFtCpJzZSfSQjqPxQstqFNkNKHHd46Js2JZcdUrXpJGK+
zJgcwSg04f9wg3dOejhplTP0zZ76UQ9/NZ8aNj17EuuuYuZYJymrnPXfn1amvFH5
sIBnLk2xVfPDyg6JKUGWKUFrc9ocZx9QZ2tyb4LwRyKjNaJe8V6n9Uz7GPUF4sU2
b7aeixycWT53lmd2PPWGj/ocSKno4IIEssU54WMaHw/tV2uO9vALhHBI5eiNTeK6
IjvIj4ew935wG4Dk6HyCkhA2XIghMlheWwkrGNF/KtiweDfuFDjFL8HmDwXtptXE
+vBPkqBkc+Xy6oTJ8nE8M8cA1RPS+/yAeR9xlr+Taknv/vRyoIMU4fwU1pZZJmgW
KyM8RJD9tsEReaF/AfMPK00XCIvjGCzMiImCKaq3S9lyHguLupBedFbV6kakWAcS
NL2rOAOeFRuBwVmvutAc3bvTrq8LupCu3/yHpcCEl9497UPFdOq59XA92E4eYkBg
UrArppz+asrBv+lEhyLjagCdTet9+DGDuSCOmoMm2x2HSkPZOKF2dp8WuZVVx2u+
/gM7y/V4sd5PxGVArpOm6E7GkPapdfPJ5b7YLHW2cJ7PKCXdntNBgAKyd9zpFRR9
gJIzE9Ny68StdFbsDfGAEMWWSkIfXapT6wemeQa7mOcmBld2LIL76491nB5yEgSF
5H1eiAETIgeVzx9Xq40NSiIVWCqb0hBXsNp7nSa0WnMY2KhbJkJTgAah6f/QkwHa
VQBDzwkRBE1p3761pgDmv7HEpAkVFgYygihis04YlEeNRYh69JwN++byAgbEM1x5
E14qS6Xg6YjElPF7BBb69gqPi72IdaVNI5UE4zJy6h1bYyW9HpBhHCLTeJxz47Gn
7jUZd+NHT/1pBJMxwuN7MUGn824Wyzeqj2z9cO3qACILnhqdizgLXu7PU1Vmltrc
1YXoWQ1DfeNnP6x3s1Pt9bzUGfUHivHFSS7ZCYLq+cFVgPbCcBagJE7U2cjAjCT6
P3cb/2qvJlQ6Chg318wffTnAJinTO2mNc2biLJdvaymSocGek1jFmnTc8jdcoccU
QiWMNhiy9W7ZsqpPre2Ge5lK0NF5uPOsn4QnonSbQWjBXGq9TpIt4SnD9Vvx2BAg
SyUsYLr/wUarxt36JGLkYpaV4LGQdrNhB/Z1vx+FAcmBYScRR0EyahL64wdmAMmv
xiz6m5Ml4i44aOB+ZOzeeLkMuIrcA0ieQbmGDVLPqE5sboWNBRCV21zb4M1cfunV
1sCQze/VipvnpTNmZLV7VM/XYV0UxMIpjmy8CkjdARh4Zyde6znGZSlgyL9ndWrH
MCVwniPXhnmvpSsfks3t6mTlQCHf4PkXxCv1810/yl9GaKOydrRvrS2h4Ix65jFF
XOGvr8jejI5sKluCl8xLZwAxECoPcvSFemRLOaVY2NsjHMeiK8bh9EOwZbT3/tFD
xvlAJMkjzoxGS3Kbt/WBCAjK4EJ3MiIoIYBTYn/yrk+wP1S5AwOdHXfNoMdqK5ub
/hu6pFYo3L3ceVaZ4f4eZoOhxBQOumHMbM6+iISxQ/xZOrrwdQMIoXnPCKNC62mn
We6fwElePiDBbKa8z2aNMwVgh5V2BrzdrGTHn2oMcnUzbaMkQ9hfJGaQM949x/Js
MwKN2KWujPbT3JNan+fwl28/TnvYsI2UyhJ/R4JS0s5pFqSbXPfcIuoM5hPNGg5L
IqEc2KvvkxNOQywVvv8yNqTe1zz6JL7nQLN0rA5AEk/ziw1wxl5/zP3hjPR63xZO
SHFscunEXz69YsFl0WOScLAMyMYzCjONuLg+EOwpG3FvdrHQ0pVU49JyAhre5xVq
SS8TrFWlYVmKvkCoWdLgl0BsClIAuK1fvRCe+ju6ON1JdYpFueBWixbB8tyj3Yfi
QrI64yfcsfuOnlzl2DVsXt8fkfv3Ut3avlRSvA4lG8cpvZxmT7QJCpej+ixsCDgx
MEpmCJ5qgOuzSS9iPaTxZdNCnokjwceDQf17/bgvtUuLA0saqEWL5QdBD9NoEYiT
CKzeMOBrg8WAKbJq/DCHlOkPz5wy5OKmVpH68SX02w6RkZ5LRCZI5QCClXIv3QI/
XXkZcKtQG17IyFPnEHM/g7hFCbjKwEmECULF6UK/M5kT0XfeP+oeYtFedIjpSltq
dFSenuFa86rgd0CEaV3dxS1NcUM7j+4qE43Iud2AqmG+EnScZZUEIjUBliQDMGw6
GQ+DtTzRfQvOci4M1sD9yeeQ7Cr7Gr1xXRbNFBrLjItk4zkPaussyGAnheAmVt+p
KDtmnW4WLkYQ9itR23RxlAtr2c4lzE80ui3IdgzwUdqgzut82NbVQe5itulf0/hC
DgWOKQnEJn0tpayMp40pFI7BBa/oyt+csL8HU6A7FTYfABfto6uaXrSHoQeDN1vG
z3+u5z9ufZ3GYmxQqO6H9SGNG76fjTH6Ji+SiCnw9eLFK9CnN4MQNVfYdqL3Gb01
qbZza/6iHANdShjqG4cblczVim8Yu8c2BSP1RSaEmzAScwHbO1uzyAfKWof35KHr
4riNeUF1BfrXeSAaZ8KGNUs1g6/FSNAlw3CSS67Mzi+AZgeqnlnSOwCo17AgAA87
QVhxn+UlzwiPdssJycNbCz1onuC6U5d5czTY884Hf686XaavGf2xzncmcGeyYX8q
ZJSyv6v2XoieqZHmilu7Rf5j6c/Y4JafH3cdS3m5uCZGiPxDUHIclk9x+ecfEKh8
ONRXSWbWVeb+85JiviBiL92v4QQDIKg8Jk7hWUEBZsyaMo1s529SUb2mU+ibtKu+
31rjYaoEnURCodoLwNdGevTLRlmDWc3Hqog9PaWsGaEgUqU0mUJwzGfOjxkWSTYk
ToBhpjjIAxICTa1dCPb0CdsDxQlKRV1QprsuaXsLLIw3cI5w/PCTVqBElg5DQGCj
u4j4kcKzFK65eDMNCx6ZDuhXXPKCNUnW3h8bv26NeMEQbVxKpBMDhHRRYmoPc+eO
jgrAW6HUB8cd5SbAo2Ldo3i9Hc11tXV67mYxFsq8e7pw0zqVwusYEEnqTAaY+rmw
+WnDSFG9kitfiEgDuySeypkZ41KJnIPCn7X2YEUEyACK2JNlk9RSJ8DVqn/3dTvk
Mk7GOD/o1IAaS146R8DSlwu6GNnq22H3/NtsCc5VwDDcHjttfojyXQ4Li9IWib5/
clgV+WDxXH8rfG5EjPg72uwwmu6ov053bCBD+Q72uS+jHS/3qvCeGhwSfyPAkq9b
3gKv2PJc03BA/ksRt0YVlgFV/rj8dV6MQPGnd9TeTHBZfB6MIPQZehxNTUnvMmg7
2YpoS5r/IWQvElfOdNnRHQZM4gTAJO9rBsd7zKqgGIo8Gr7OR9NWuOETMTP7SiVO
abKWFOMKfzCDfAO/+59d2w==
`protect END_PROTECTED
