`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5XCzkAXAmbjwNk8qBEPKwIG+RLgOHPGQOm1nyoZ61E/dDaWaDwvBtC+6GviVsPyl
9eHLHwJn+g/2SMhiug0qwuImdrBPrOIkMGHsaza7eJEsULyWBKNbopE9xS95srOi
88HkPCi2jEK6dNQWMC/6G7fvPQMsJtwna0l1DFl3ts8RjwTv7NtTIc22kGYIgV5f
kF5cryIFkxsdBuazaby+savcYcL4fgV13u4HLUWbXEg1Zr5pKsS2vzFdlHrc7w24
jarXuq/AxAt2BpEV78gU253ooEqySbeT0yrXor2iCmOLTsYCF7fYAPriUt3+nGDL
xTRvCqBfw2axJgbhESlK4/80Kw/JxZvvwSbHkerPgvqh1lGLsAodflNrQyeY8pNQ
X1QKONIdqLtpx4w26vSIJ3+yOZieDLmrt7jUGEPj7zRw6BAtJ0/UMr4vNw7VMLbc
B9mYvKoKeRviAYcMyyAxZWHepjIg18cDxQdhdSqpE0rwO9s+naFNZOBJq1qCHKKa
gbcT2nd1ukshVgEJFPRQirzvL/2oxXWqausVoyzkt4KaM7B2fQe5FJyRjoxs/yqk
yc++iNCYKYeRWpxrlys7THN465Jt/5NYi9F2y4YxiCd3CPbVVHkT4Mg4MxrGwbiG
PYAjpjRV2gijjIDROfLot0k27aSYSfJzVOrtQ0o+vWsvYSJAkW+HAU3f7af1xYpt
8HbagH+3pxv3rzFcqLnygg==
`protect END_PROTECTED
