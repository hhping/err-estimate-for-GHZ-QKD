`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9NTeuXTP/cuhVj+eQ6udysEEASv3nB9Slv9inEHcB+/SIjnf690peepXrMDvKUe
+cMltDRrRiytVdxJfLoUtdqw/aixVO+PbvVf1ZJKCdVGaUguQvfv/YXZvyhqNTZO
hkK+1pOjmq24cRW367cgHGReZZsm03h7qdl1dqRenPwUtUqbQvbg91fCJyFmryEm
RsOQLc2ZWgpKeHG6M2c/q4s/10oBP19QKhrw/WooTeul4CDIICR29kdZSoVXcU1u
7wi6HZftzfz+1E2aNsoYoAVZQEi1pvNJ91pmpQLjsDUb+DBrssjCib1ZXQNEH30P
lzdkmqljV+gKlAPeaPhYb3Wu39UvV0NiKK8Mdm9NozP902oxh7bsqDWle5bdnQJP
br0/iPOHhjuQEHx/ocq80j6vZ7OQaEkgw7B3V5rLqjrxJxDx2+DG8B/F0DmRqM7h
6m/Bqpu8g7IieEDG6lEH4XO4XZrdaNhJO+2bydg/vr6DribeItiJZNfkquCB2rin
f3yB7u7co+nzDd3L7SnbXbCztK67yaKqQC5DFBoFe8l7KfM0Pe7PDSQuIBEWQYL5
VQ0Uph2gosE3DmlsnKXb3QrAVsK4xaxy8V/dowWQIeXie+dFYimNeRw8xz7Uk615
R5Usilu/FyusG2XNncRKWtAQ3OVQyaep39vmQHAX9DCLn0Zq1y2MnJP64O/8TC/F
ogSarnsqUqd7FaLA1OL84sWEVw+Lmn2nd80dEVeuTP+rMG8kHTubOstKp3dVmx2E
T0OhTFhm7/936GrvkHSxhTWBtUpolAvzMxUXlfZQrjGgyRonxdqdI3XvAscFwh8b
ek+sgy2PlZ3Vy5i7BJiAt8wXl1ZuE3euqg8oEL0r8B1XOwsirn5k96LXWSWDhB9v
iHhoYJT68tt0VmMm619iNJAsBmUaXhky1ayZqIR4iAe93iIg6Vsz9OUJybIMrsMC
FYhxBhQM9O+ZNKkcmZ62JHOdGqJZGd29vzEhGXF+3oVqgJAUZLWmyEXvA+kwgkwc
vfbCkbku0QegdIN0uVnRmZ3dgZOHXqxT12ZH1XmnhJSndf4hlbQKYbhgRf8z37gL
99e35mUrTnRLLfQChbPebYluSyTkHflD6xlqdXuHsLVlmBe8B/hxvOlN+q6/23W9
oNIt/teB7TZh8Yy5Qzbjwnr636EsyBDc8892HbW4/U8j69aIz6l7SPfza1gimmmN
f7xofhLd4XdR28s5ZMvbDdiYAZVRDFk4fPvEUBjdIXcIKJ45mb0vW8o3DMghVNYf
zq31pN6xPOG+eDz122Qt2b8DhnET5Uvr82uN6JRqTcMObPL+f8ZPF9CWbqm+/0J6
Q1E8x1GNKOkvnfCWDXjtcx/1iJniWBv8VzcCuC+3N3qL3JTY48UPs/JYBICkc9HE
G+RiUg/yDitWgcvKgHo4YmCe73x047r4HkX7y3TLCkCe9mH69BxzoVdxr9CsRT5U
r5s8/Pyc/K3JZB+QNw/rf2enylRS7PoWezoxzYK/laNrh/rXXYWtzYnGKWge6Z8+
eKQdnSDdE0bewQIjt55PFS2OR0U6lxRAPcg+dOq6u56HSXqXMU5uCUi/ZzjlbJMy
JJVMDnqaQqtgh+Vkg5pAgjEl5SwKQOEc8MhobYJHb6mM1PW7QMMuLj0z1z+O9fuh
Uq6RMPtq+h33hPIbt7ft6O7uxNNH5ZJ7sJBeKIp4oyuIx0cyVFyk7vqDhFnc9nDx
`protect END_PROTECTED
