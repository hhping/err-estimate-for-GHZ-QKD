`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJz6VY6GrzvcQOcQ6YM1XQYX7YpSUI+8h+HV6MP1/2vVB2F7M40PKFQ/5Yzw3qso
8t7evzq3j5yANwfmC+lnSjlLJJyOZdYpjWbywGog2RmP8NgrqI1osF+OIb2++c/I
UicPVzIn1sq44ufOmKN5oaaU3Gwu4mvdiF8pKtt8Vn1gkHFSxBcmVwiaQNFWbHYM
gCpr2pfoFM7wnEx/7q/KRoMY5oeJ50tA8faj+vB3ePfctAibsl23D+FSOzGsE+Ss
T0P57ZpUt0Be9qtSbkvph5HMall73rk975u9xGJPGBey7isZSjE40Wypw4OQDB4N
4Nj5xldJoCL+6noMXQ4nsyFnbZCSn7IHg5Xj0l+ScGJSBSbUGOf8/rJTha8W5D4B
6sD7UGUho8cYEwAL1iasB4/F3U37G2CFpuw6KafFsR3zQtATW3G69ilvsgMsUWzw
Sy7f0x6s2zk214Wbkqva1BWdaEVGNk3+vvoNFRcsRYIRhjwFkNlXrS7oaHTjD6x4
Pd2R4u82KBf7+iIJGWh1WllrCfD3DE7wx5eSM04DlPhIdjZxNg1G4rnnpb/bXx1c
SgUDx03MVJGDizSakVd/5qNTi3oPocmxGLASP9lFNm7eaCk/nHl2tP9pMhUYwvHq
3EJTJIn9fez9Xe2y+xJFDpaMgGXxbX0VVc8kPyUr/emTRZTjvWu5Xj3kH5GjDEdP
sPyhXkWFyYspwyP8lul+JzRUyMyYu5rV4OQnEhxXvmPrNndyIh3FIYcsNV4P0l6W
3Zx0vEftHG67JPjAg/zpLfh5TvU+oTdbd2xx1umcYX47CAFjeQl/SkcFPvd3Y2oX
NIk8e6VBQ7SM0tV3i9JeDiVgbTARB3jHroSRx0b7MFnzzRWGnrEZmyIX++jUI0fP
rnvsu3oKJqZdnlT5aErI8xcg7rLeaHbNhy+X8dTNCpDi2K9P+aDTth/c9hzWbFQk
EIeNb1NJgU4PU2hID//ljTOF39NRM+hNcZtkb3aBw8g0Gr8S9ehSHt1ZBa4JyXfS
UrlwhIgffwu7CKfvRrpSNrpCpODo3MM00HuSBLpSXXyHKMqF73zsfDWTdvAETfvG
OZM0cY171rfxoZ9zmSxbzdFo4YcARUdlYQpA/WmCikGV+qehqt1h2gnzw5lTq31q
gvWQXeST9lgl3jBqVzEzMkQivkQU470sVUDBVfg0MskagvneML4uqvUb/s0H72/M
gGBN1u2q2VH14YMT7X6wTAV9nk1aG7A/39Uux2c/z9WrYPe3oJoe9E4wi0Ujkui8
y3khk8A83KVSNU7dtpuV9mndVIKsabVTY7zSbUIvCN3PVaZHbWQTtH8LK6MoCX3r
GDv+t8s2eb/7nLfHo0UbagMg7R7nEOW1s3KLxfQiDxLj0SKwcBB+6m9l37SUK4WV
dScH6JyxpBR8n3F8rD5o1JJIHJice2MafrWrDm2ipdRmLcswYPMbUuunSX003AGr
wuzq7++HlMdpp0Xwocke3OoGRAJJh0NnkCwVHVv4MqTp9CLybOqC1dehiQkyFUYY
ES0M57oAUkw5aFQcYHtXIygdL3py1wAsN0fPWZ3L85ojuGcShhSJX3ZCVBzgGaWw
v1csvxmfcWTgFDc2z7r9fOeTvHFsjd3tWdiz9xMmq6yR4UZPkKLcdjManokTZJFb
zncayBSrQjWxzkcmAAuSo2nsmj+X8B/Fz0Ml60SpVMOdVtnc9Wf/Yh/He7W9G5ye
GuSTCWr/uM0HYkFWLq3N2SjmccSrOC63Hxljxy7oA4xaDNyBO0et0jveYDbV1RaA
rU+DM8Ny4ku7hQ5LFqCCFgTGZjEGRNTmJCNjOyCfpWBVlL8w64fhW0n6iUPcwYqb
1k2Ti5/MyNi9Oy9nVJQu06eOwOA/FYZ6D9EOApZS6zYa8Bo/VidQOUJtWHjBZ++B
ya8iEnsR3DA4F2j3Chrh/UVTRJYaQoZMYxvBKn3TSNVukUMNtHwHn2ISWEvhhLlq
eY16HiCiFWjg2SI0SozdoejpWy9fmWiycw7vffeCzhqrtIC/QStRKEwi5ktmuoVF
vDhaCpd4KuJwQxOzxLc1LOYzg+LASoi/qLRtRzIaKLAPAtC1APap9edo+UfzDQ5T
65PqGf271ul5HLZ5FMc4fMquarpz8YeHfqocTEsRQt3cVKyWNTEiuU+gSBk6qfyN
J1fuCwpb+lZ+dxfSsXsUPagozgCBmDUGvb7kjG4OMTr7x86yzgYdZdNz4aD4d1k4
itwLUaopo/vFSoCv9xynkqU9b+ASwYn8Qz23lSDISC09ydFjaaCnYrl6u4E01/Cy
FTG3/fZd8Kg+O7iXQsxCiTNO6pvg6hoXe+wTlcPrkXf8fhe88jRgCyr64gkgdMF0
KQFyXMnjBFgwXClN9RnGQCWkLiRfshjF8wR2qYl4tZswK9vyNwKw/2wRVgslPSeh
+oxi64g/gs7ELgyJScZaeBntNUqAIn53xS8cL4YJNWEZ0R3PgkSfeEHe0hIwp693
BiO5HtV5IQagmKPeRbvlaNXYtQTZ5pQQ1iYA9Na0QKqtkVxM980kWZSFkUD2Zb8o
52c5iqkxGJbLb5g0eVh/5cLTIKvTvtEHTzusAd+N6W2aZwvci9JWtmnOuXLZkb51
tsw+MC2hu5yGfK6UqDBy7lfypJgRFvc7Qe2VUuLdLLkUaPz39XioIjxorTSE0pVQ
8eBuFOPbgCQ4UoTmSc+aJzTZYyrcUTmVdLbDSnLqtJ/tFnvwf8igYwZfRcHjcqyw
0kf9JPIE5YJtRhJRjsLt/M+Hr/0MJbgTpD9aciQWx0gD6QRxk4rKL47NdUfRrtKd
6QGV+mca5plbSiEyVM9GkY9HBk9pjpuYTJx9w9gGj+y4DXtFaADOSq1eZvpmPIjj
nGs8gkGi2Ffs8pLOYE22muAfeYTb9gEb2Iah2LSI9R8VUAuQ48vPdJ0NtWOLRBPc
NFUmkpLLCPi/Qgkh7bW4rQ1SvjHQg9U5UBBd7bU89O7FYlayGSsYxZ8qQzbNUR1k
TqGWF1keyub01NZ9IlA6Wc78/4XV0jQLOAYHRKZf8sHFkvnQs72ekpUcZn7UWdxv
h0g5bNy4nXgpeYWyAo2eTFLonK+0Pn9/W0Bo3s1vLm/GTcBV1dd515lP9Y4WRAHK
OBSzz22uZIYBO111pvs2HdGuJIX5Q7OCHEw0NiepziYU1oFWUsE8XzLk8U2Djkym
XRmli0t3htaqYf5NG4lPkoCxIe6H5pLC5IG78U9qR5ydXFVTbabQ6DsgpH2/ri/e
XdaX6Pbyp4zBmScxq65b0odJRaHd/nrx8rVMEbjV3ym9uhulKT4KmDXpWgfOWXAT
`protect END_PROTECTED
