`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97pgPOQ5SW9ZkF3uNyn56ekBao70PJAISCO4dAW/kEpfM0AdadihmdMOywiZOdxx
lQV2DYWgaZooeqL0ElHYSLuU9eRtYZ7wyG6xsXs+SqNetHjlo4Z2R7XPtpXQrkdq
r6xATUC9WbOSG61lOcgD4+56TY81rfiuqDuvHqtRJopocNgd0ToFG6S2vPA6Am9A
znAe/fZ789UbCqjlvsSZzvvC2t90iSjZrPy0mOtlN5cW7kFTeaUCk+WFj/NzgVJq
wqV11xxl6Fy3SJkSUikLQUukZg5NtDpDADasGlhGU/vDi5RiNVnOXMJ3jNFi1OZe
dXV6mf/XNnv71cFC4KLVS9V2NmFfhhgUJd/L3DNxexJ45R4Q6UVcBS7ROqLDu2hJ
hQfWsWPfwcZ1aMfBbKLGqAqfPnbcKBl75a5vfTkag1bT3cV5wLZ3zO9W1BnWwILP
wtAKDPptoTfNFkbc2C5rIOfEiGTEAL9SDltYyGF3G5orNqG4f2K3EUfEM+YrH2+M
a2oQJxlFP9C9c39feSMflS1PtEFlE3BnxoXwq6XkW9YX4QBoMyA6eGhjZcR0DL7e
TpYz5LqwNirQPyI4T5k1aEhIkdHC9o4yVq3JFTWxEaMGE/gLz6sDMKF2VA/8rbsE
kOTu3Twt9+ReuJ4adLFZChHZpLa3zGzB/jiO9kZV+x/m4y2zK+UcdDF7AMSoeezn
ki5tyv+U4/NXxXZIMwPUZsh5gemJelAFCH20Z3ESlI/dbkhA21eWKN78cz+gpfsf
y9qa2djQBUPrZUWmTlf9FCbZ5dezdGpO4VI0MYCtFIw2OtGu+gTUMuznqMFL53WX
Y3+SkJhy1YfGv0ga9Bwae57js/dTrVQKnhJRCp1M0zH+ocamXOKBWCbaEusLBmTA
k8oVfIdQQ+rO1xLxr4KujbyUL0xw/OpYSdiV8+ooj4UyuoD+c+eEpijIBX+H3X24
JDI6g0IhpG7N18d3XCkygfzL3gIfzDKMmLUSWnX4tlXnuLAeqpRKAmlHy6PAxfT8
N+oJ3ZFEOSSl3gLkVGIKOc1PLhMTBBH4XDiHaTylgnMqc8RIP/Gw6oAdAsghLfnt
Hgt7/KQkF9/N4KFhP3ObO/Jr4b1Tm0P9uq0hCwjWll1iphkU1Ox/o1OULa85w/V0
O4JAgCZsdAQw37OwU7ZiEISGPM6E3C2PMj4/dR2Wstw7mBemWc/WExGxnrUx0lBx
i/EIeULiH9KvUkCPVwk5sDQwjIhusyp4qMZ7oJie8/OLxZ8cM/K9wRqWf+H0L3WG
i4cGi8zyYivmFDB89uip3Wc8fhAE9tI0MZ3Nv2lCzq7OmRLIMazW8rrZxWHA++Br
BtoaYaa8iY4R7OZvI65ipGLZ077JNYXrCBxmuFLppJ7eK76TKHzSKVe2bo3hfHtH
8RoQsfBZnZ7p6EL/uRQvXofVKiHBW5bfnhqLK8YchNedO67rmgPsFujhYtNKEExo
z1L+rLBP/bBQrTWtJkXJiqMPDLUbcyJcob3Z0KKT2ndGJcASoRBsXdZ/OYUQmScB
WihsJZA3wAVu5SEAM00XuAlTPtM0ADFS25Tf91ysOsbq3LquxY/2Q1VfsjEKmsa1
kDC4FbF9U5Fuj1lKGgeywCxyw9moI4GtReOmhwF5CMXIwXkjBV/ftICMShrAgUYR
i8a4gVNnR8VNb+Zlr5oBSMAfn8M3gXgjwc5VxjcoSBdd804TDY9ICUnVqf31B3xU
zgHLTr5iwDji7QGEJGH6qk6PaEk2hpNBOTSqIg7gbDlAp1j7RIQ/CNKOFSHqdgPe
bSJcC+98WfrVEcqzlxxX6P+Kho2JdR8tLv1cTgiRryJWAw2WrgOk6WXlWBdgs80Z
Squ/NyDLoUHz0V5wARM6cX2du/fPHj/xSJeJQlnhpHFb8Ie6jp93ZNmRNOTzJ5XF
fV9uOBBOTOX55dxz6LSCKB33mkTByoJ7I8DsCnOHNhO8MqJOlfuq5i3Y33eVQY1P
Jm6ww6v0oHYFtn41bIFQUXvHh3V8dldtXkd2/IGbe7Sy7QrOIlwfLz1L22L3ZP/E
2nIeefEwS3+d01xJpyNJPxsa3dsxIZhnsf94utAPMeAPrODr8nf1bBieOAkNbpIU
UDt/2fjPoN+vihCURtfb4ATnjNlh60n54yHMLz/ftb9r6onMzzo/s8CBmYrvNXM7
2ortyZWLUYEpJWxsamGKH19qOzX3j7yJZhHKZl+O8co2qfGYOZoKdboTDoRjxVkY
2tQ9a79EKsOA92lgUPHkSQnbHsYfIWDedLzq1X6dRm21958CZspNmHoIyngCmKPI
NCxLO9kIzZvV4bbRg0NvZ1M6HDo1Qeib4AzZRas3pjeBV8mSzWngHnP4U3UdL7NQ
W6/pfogwQcZR/z9sdKFYXjmhnrSPQWixOefqVtLUq9U48977Zshkz/wNN90SNMPv
p1VAg7+NHPmpoZfA8o5n//YUsgUIfdAG+0/z2lqeTVLNGjIxdRmAqM9YeFOBr6A9
y5SSBItoao7twAj2zf5cx3spLEIlXaewLpzgH9WAktM=
`protect END_PROTECTED
