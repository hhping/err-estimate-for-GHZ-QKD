`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3qys2t+kVPKAduARbyZf3MfrMNUHnDsuF1Mcprn/T75Pc2pNUXSIs36v0uM2FM4
WPHYoSgHF/UGNf+p+6MEaonukXDiFmsSGB92aXIImIyhPUicOXU/7ivGlTL/cZ3U
SQQ5kLv/eFRPKtZQMtVsrFcPBgCihGjszzlMjHVEJ2S0owCBZ5hdaepiMvL5zY5/
Lo/ofevP8rpx2Zdd6u+cbLzR33lj5GR5w14JJsFnY+DwVd/ocnyVy8RNQ3O17xwz
22oRbcdMIfmGLW+5phhP+Wd5E4K7bKaxyexZle5DjZqrLx2IOG5EqoCNvcNO79h6
v5wHJMjsIp1iRlU4GN/Ex06KGPJ71K3UFNAqMSTLuhTJ2zkIMnoy04t3fsz1iGKN
tD1LzAJBSjlnGem7RaxcjkFwdyGqcRGkU+4XvvhghAzFhqh6Qbpn+bchC/7Njsur
`protect END_PROTECTED
