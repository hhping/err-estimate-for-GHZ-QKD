`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CoyxojibDO5BACPais0LBR8ksr9Gu27e/ssXlAHrgrOTj5dq8Pg9FoLNR0fM+TLE
+0agoaF1eiMQwL1rElUAWoxK7T+5HkmNp5pVR0W1Rti6v3qwg6e43Lx7Q9mbdXnK
ZfjA/l4aHuHTlfrjj3XdCBtX9JJa24ou8vpRs2BOvCmuAHAFuYbYAzUJBYHaY+cQ
76D2ctTMZWvLHUt4nTo9zhFMLcGdpK0pSJRX3cSKPdQlwJI81vmTNdJgylyiTD65
SZTePCzRPMNjrMMYRJHISEsUt732QrOTeHIL/iI+w+tKHt2r96UcxnYsePezZkN/
lAnIy2UQC2H1RaLNVus6zagS/8av95CiXj4nD6VYNgeQbcvT0heBDMZrbe6BXyPs
kSWFY0HOfhcZJVDC5b1rs1+6sCnkNbxewc52OxozzOC8/QYTtElfvvpxky6deEi8
`protect END_PROTECTED
