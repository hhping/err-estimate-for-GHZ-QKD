`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gAxUrCp2xa1VWyq7BjXQm90qKS2TTU7Dpy4YuBpcbc5AqndTBoLN0st52zlpJzRn
8sL4gbVlWvlwnzdzcuI68CXX6u8ZxYAaiFaXCK9ZjeO7cODPPyvfeE0yZc776C++
y1vUxyp0u1F2k1JIdYkyyO20OBP7eJb/lDGXEo2BjOPmCclKs34u5UBGntJIrDs2
9EzfHc+eaBprAyNHNohxomhV9VP1NVh/wF1ZHBRBfi8R/ah+2UHIyuZyS9o5WBHE
eA2M5+dRgzBhIbV47nTHVifLBtYgc7b3gE/JcCtM7salWBx+aXFHfb1TMQ9SSdaV
LHIoUzasxdjdHEZJM8lygMVng7hPITeMMYOUDbi35MP1049+b1cW/3bP2doqIQSq
e73N0H+BazIcqXBqjs1uHH7o3z0xKbLDIdTw7QGu+84sjg5JrqYupu58fhLbYXNP
kMyNAEQy8WJFx/iRK3tjlePZ1aW0t0Md4k4lsvPhGvWnQ6QQMU5JCci/4rOGMH92
TOWUn3OrUzixv2bSnFz45XSV7s1ZzC7H0JwSbaZI2WNwlfTvvoAYcUTjQTDOv178
fE9xyl4g4+P1BdTe/Mq8y9U/Als4loIiqtlITdbE/XtWDvWT0JwjcXk2/IlGC/ju
9oif56cfDGZDLrf6PH4WtvesMHi7Xx12XnY3kAgGssZvo+W8DjrMYCeIq9CHPbWR
1x9KEx+nx7hxC/3wVJrJLHsk4r2ESm7eTBDtfBnH/os6UkARuvvwV1OevGEGObxf
CNHnQS+ArleUiVfA5B0yvXXfVc991jViWgHuCX+xmC9OWM02SRIj2A4IS+lF6X0b
vYNGgovyFQsi3X89hDvI09+CX/j5jq1G7cWw46Tr9eVcwAQ09ZLkrYbwo9oU+3jB
dD5CJp7HvAX3Q1xwJJAV/Fj6Rl1GrYQjB3UJLZYbvGt9ZElrNH6vX8fbqiSzOqeP
nY2XvosW/nF9m2dPW+XaTPxWC698w1FH6xRc67WUpauhHbY0pgVodVG1VNjOOG/2
ibRMj2BKclk7fLEEqWFc3jQsJiX3H5Ato9jewf37J1JBXX7wmhdJPi92iHhTBJtv
jeed6wnJO73zi5V72OvM+12j39iPDxdUv6zoGjWy6arBnLG6ztZunWyAQHGBmDfE
VSKGxMAi3Qp0hWxrgZhOcA787AYdlsrvuHSDvfThGZN82cB4gchxciigh0BdmMSM
DX1CNLReM6ofb2dd7hkWXUZusCVAF/jmAqjBLo1q9Kx15wZ9UAqpUWyHjIwZAF8h
9Xv/2DGtXdNVRts4AlnwXSHbaODcMIy+2zIbVmIOR6n+jftGdQsAxywxO+TBfzYs
1aS+vh2IlLxqSLABitVazQtQm3AE91hnHeP21t7fx4tZkmPT4qrhGE5DpHLKNSHi
E9+LMjJCfgF1QzxMRjWvOPmqWN+SITY/TBug5AIizy4/mxIepERhFgUR3caPszik
e9t5JX3pFl5VR4BhRsIbfGd+cGB6uIJCpxWil0co2LE=
`protect END_PROTECTED
