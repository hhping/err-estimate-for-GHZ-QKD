library verilog;
use verilog.vl_types.all;
entity fourteennm_iopll_functions is
end fourteennm_iopll_functions;
