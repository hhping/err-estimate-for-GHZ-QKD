`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LwlQWT594LrQnjI4IfgceUESS3r2gYdShZWDIf3Hdvnwm5SD02bUz6ghBpdYW1lh
e2gfLoQY1dnfOh6eNDiuV4dyXfIP/whfznq4giNZxnx54QGNLDD3W867pspEMHTe
1I5JMCZ4UYxKWtEfj+YsouEiEpwvL9h14O7f2xImpvafm1f478Z2RY2R+4Y/wGg3
MSPsMdxyotetlE4QubBWFR8yCPq7zS8Snj+5LMN7vq5CwZJvsLQhvkn16bmn/Jcj
fTfhc/256ZBy7dobBO2Jan/lhNXjIzH3ZNFRZrVl83sjPiPumxcRHtkjVShIlQfZ
SzbDcKjMyeWZfp+6XA1E5ZHQHkZhOb66m8rRvFsiX+zZorB0RVIeUTL/5uOFkpAs
PBXpGsh/eUD20R2TgSzqTHCblg8zv+iuZygWWRcRlHDCQe6cV/L692NaLO2KGri2
g5WSuaMYza7Alc4bY8Xzsd+KVQR+b2cMQ31UizZ5UX9h9BriPM6rbAlF5TPJEsqp
SOYuo0N2UQdZ4O6QRS7qzFySg2KKuh41lIFEOgt97P+MclLauDFNQXue9c/5BP2G
j6vswnHqLXAE7Zcjx01NTYZO+xwdMmv0hkdjIBbS4Z5PtA8eLe0cHx5AuRGuObaa
XpzXr3t5YqHpSX4eyviQPA==
`protect END_PROTECTED
