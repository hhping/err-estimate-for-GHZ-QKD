`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVH0eUUXz9Fd2teyIaqskl7TucpUMex7FlzawWyaGKSmI1gxhz9kE9bBCeoZ8qAe
7E9xeO+6YNTuf2ijqknRgwRb83H0kfE4dVZerQfh8WwFJDeq5FPQFi1kRMnLjO0D
FDadnauahrOvfiH77WKuv244ip91vnDVSjuWgG7UeHjhNx5wS1080RReN2vYFkkw
6+43SJBq9NJthbaX0D9EdBrj3XomDBQ3qSQfJn9bVgeAF+JR1yPQnHCHKlD2t+Kl
X33cEE03BsYRbKvL4bAPumKV/aM+DYXGzG7uYw9UabWgrwzzOKWrxjBU+lcbRanH
7uyZ3gfcPtuxXrW36f3O/jgznyJFOf4P5SQb/AtTyqWwy2vYrtQCeEPjxINh8QJG
PfT/jWJaq7ag3drzVxt/pkxy82zg+FbwDXCsQLTXtpaRbhFFU47bUKBw4k43im58
nJ6h+Vjku4z+NzeB7wxQ00gcwTeYP6edmUSHCff71RshfeNrAKQFOhqjfVFntSKO
HZtOVA6YuxNDl4/EtHGYKbhfJYv1R6nm4TixG6a1Ih4/ZET1Qxi6dReUz/GGEUCl
Va+llEEbR79EFUi3mc+O7xz7wnuSWYD7o9KL2a364fesM5Y0m15nMf4++oc8B+M1
hsRUxVG3gNXMUkA82mIVJTXebRMUy/92orzRq+Yawvpf/7suISO05mIXGHfXHq14
X2X4skcTVlPw8VyH4Nzq8MnLBL2FidFGdlDxjMomGCwGSk61c5m5MHoPdHC/cszd
`protect END_PROTECTED
