`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JkPAO2vfzMZYORD8+DZjEXyKzWHD3rkl1cFM7t8uZBPDOtdKm2DSKaCPP8s43Cq
T1ySM/ZuoO8AYqsjJp+m9oqV/ydqW90IZT4ic71lSQC3B1m7HwG53XWPJCDO9pRi
I2Eq+yUGekbSd8drthqeCaGniR5l7T4F2sG0PPC28zvE6seYTittqqkjoiZaJBmH
tddwZF84eEy6DjvBTD4+zl8nSYyl6+NKN0CsXSCqIywu/Zx0WKfSpsWqUBbKcOnl
Pv+Bpz2VjOkuVq3w+8hWVH4arIEV+d2dMKaE/Bt9FxjJhWCSFd61c4f7IqdCoTMp
eY8vvjgsbFLgbt8d3eg2fdRZ2M03rDzD8uIsHIUADa+vPS2xQitOfWXvdTU4eMex
giWic4onlA4FQLrww+VC2w==
`protect END_PROTECTED
