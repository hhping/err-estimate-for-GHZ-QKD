`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kzArK181cngNyBm5q9Vp82i2IJPnPqeRjOMOM8Cabo9jvmDAwtwuT1SmQRceqJh
1Lt8zwLIO2zolAm2dp2e/Tz9AZI3q+0N2IhSakdLghSYd1lE2COQgz4Lf2F0fJJ4
UkpJ8ysjts6/001DD4H4Oo7DszlcCBrQTJ3V6Wp9i6D/BTB6sHUHgVhoIc2f5+lQ
UKekBlb8jDrVqJYJlZ7qCxP70lXTC48dRtABwm+l/2bw3ETyol4C4L1B7HZBVAFB
adGd/5pqvRUsfbU+d1GCDLK5t9B6YOLkHY+SIatiGjcL5wCQg2ZPMUv5GJawvhdk
uxtDQ+E0EXL53TbL6QMiIFww/cP77+RIcwJiDV58DmAG8l7sctJODXz+eIfoecZD
BuFgU00N4G6eB04JP0Vycqz3bcps/hfyKlOF4K+mCHnluPoTHfnOG3tyVWFzydRk
BG1Q7NpzQKPut1eP6UWu1FVgok+pa0M6LZ5VW90edzy06/vzYLQMbqLBp3YwKkXG
t6EF6kLR1WgQ73Yfw9+5RH5+rR7u3KEsZLOMJlgfUe3R3uO2Oc8fuQe8nXQCRspP
5zhAZB+S5/9a0MHzSexeLvT168Lm+sYHzNixGyyyJbEHDLrner2ubknKtBUT/Epb
hHauFv6IWGji2Gmd+OhgRkak7PaDMzcSA1zJxfTDK+i7AAc/rbWWGwGazZpbvF6i
9hOwgvPY0jodNoUtAXJ+bx4TlKURFGPGhqQHXoCyltCOc3VSHrxnykDpCn1DarmG
N/pR7gIv6JrEVJGZ2fhCVzPXwNR1iH4EaRMUyUXsVpRU+aUEd5scAfUW71eAf5Bl
I5o5c0gMSf4dmoso+o+JFnl/YyhNRq74rNUteGfuW8JrJ33EGa4eS4FbNDhgAlpC
5Iay+NyhdtrRtDeX4QUMrZB0Zxu2chbGcTBCS7Tq0Gr2kEDsJb+gQ5OlJGwmpiWg
yE7SWIgHG664ywjQX7OHcJSGEmaAn2DUr2UCVNgvxvVvof/cizBgEhk4+WMdFCYv
GphU3laXJTASXuBs9/mWekBVQzG8yS82XXUcvz9zPaXpG+N82mOW0p57C9xRdmUK
GusO5uIBqKvwmRn1p+3yT3I/n29NQInRTtTnIaPMAO/dOSqguN4CllJsOVOhTs4N
PRtlw1pEbQq1EXE8XJ17OnQTLbD5+ZP2yS+ZvQIsj1Y9WFZWrNkDn//nxRFRCBN/
oYhV7suY8kiJP6g3ALZG3rZHTYBRgzSDpJPwAEPX/9w+SVGBRo0ZvduzkZn53uOx
uRhar+gzKU1wKkCOCokIvcc7wFWEdRJ3SwmVoLW7gzviMmWj8bXwRzDcEOL5IRae
Uu1EyBdp9KctjsJqVedxXdsta2HdJ/5kLUCGhOTzBmYgPNFhgBn6EFN+JmcOEydm
CgBdWSrMehZphXw0hpzEpkjZNwYXgbhVJxBRt2FUVhEsO1/L0wGckAEiJPi5MTr5
5a3hwVRO/hS9TjddWgl47lMyTG2en+lUKWhTCp80MLheVW44vsw5Zw1bj3INkulc
13L4Ys6zxxm6mH/Jpy6XHChnu+5jBXgLJC4RuK814S+0lcoFSsy99NwzAOy+dT24
o5y3HXb22t0eCH6WewxT4IFu0ajx0lr0fJhmqwW35Yk+yRSB3KxTig0QREyVll0U
PCAehgCotfSj3xoTuNCj9iJ9RwVG03zP0W2suIMoq1HPUdAlO5NZRrbd9VF4o97Y
eiUSrNq3GXOjZTIJ6H2qMNYiT6zeRr3Aa6X5TQHjhEnos7Hxd4Q34psHaVEtVLwf
y070X8umHWFa98/x9A7Yn8LW7a0oyBUQxQNXdeCuEvH563csYkHipYq2mVgggyWO
VxLyPkXFlgv7KJUYHqRDYMXIWZkpkmq2quqVICMZqSOlSzg27aL/L7CMbouVPwQb
ZUZuQDZT+De4RYb8wOXOsNSdA5kUQ8NkJGR8Eq5SCf1PZyg1LxN0KViZEhmBJTqY
FJ2+Ps0QZAmNRpSV/3wS38O9bWgJ8BRENWi5T9Bwj8F+0wMUSPmvm0NfK63mpc4m
wt5JBeXsL4x/PghwPXpDJdGW7Lzv9nHOSFD2HnWHf5rwsW4Bg2MGEhm2So1WbYfx
5bTsXxtp4lRf56Cy2q9hRNxacTjXAVig26k1zUsURvUPbVvvCyOs9MMVTgEaklGj
p7lsZYeG8C0RM8GMRntUcLhYEq9GyGoe9VBfH03AFpxULTgrOFiw65Vg/qcewgKA
jVsaK05Cz0OLcg+yPuctrDSTIJgTZ7YiRS3m+y1XYfdCTrvL0hZQ+OvzAit3WSBo
Wqwdc2OLLsn4/p/uScHfFfFms8kHqVUgsGm0CoUSPDKK1M1jmibiAtauSsCgjz7J
4H4hMPvbDBOM4ROfqEVE/xldTbOE9rkn2tZGs3ezni4IbyZ3mY33SOMv7rEYpQ9v
t3ibdDj2UznxW0STrJPTggaEkgXvosgb1P9ZnBkOT3GvDiYMjdTL3AQ/qLYAAoGf
ZoaWgPIzYou7b0hlCuOKkwOqN+XMq3w3q3gKCIw+CwMbHrO3NcoQpZIWx5BzXb6R
Iat9uZs/qfrQnSCW4FDgGHjpEcJN9E3lOTQWe3IVE4mggyvGkWd3XN4Ku1VaplVE
L9EyQXIwgcAw0RsMXJOxXW692cH8EBymrAsVbOHH8ZP/EyBk3NaOZWgGAisS+KEb
BqtTdoO8Exyh8iwPfY3Q8eQ+irzxgvU82jveEZJN234C6d7EZytvO8jOmGM1Fgvi
7WRCfJnB4uDz/opB7QnU/U+qQlHpGi5CkjiHpwylxuQKGT7rzCKl6em6srZK8dpf
2SeKemT/MuInwwGUjSCybJzH1M9Bgbg62rh6QD5If+c+vvT1A8Gw4mencO8E6iLg
SpEG0IRgWnoYyy8rKZXQSe4bagDK+uYemVKps84O9nQhb2InvzC6fnoKFpBEK4sC
O/5sWK/OT14fO6PbEWjJziwr6b0nMe08uDN23O3gbZ3uud2IgSwFVqy1hohrt5Xu
GqseexLBxgFaVvkeuCBDbhC970+xOyc0M7QSPHpT6qgnGquU4wLHGU4fdTnrXjDo
x6OCV+Wn/L2dXZjjfJmcZ0IaKzZx7dtcEuCDgo650rp7Hc6YGnNcxDpjIvw8hv1B
6KTwgmxKdw6j99q5aes2xqGVPOgPnUb1vxgbrdbrAOP9cRW5MmWvO09pfmbk2/Fy
XNcY6w6yGJrtPBeye5hOoxzdz1/f/2inTanrNKXIRIN+0JDcUPL942jCTkhn2Xty
BnYDHaPyAUwOWobCHRyHVFxtGkJXyJHUreHjjCXP7cEwi/tD9Kq7Lu5tfpoooTWC
W9zNfx7/IMRCLvLC/E0N2RF+0z5NEzpODY4wsRFboAFNZp5KEfyryP65b9/qZpiW
L0+BOwYA767DNO6uXXN/vPC3ew17FtcW5bvZJhFH9gtaV19YSoK9D/nQK+E1s67P
wCkDfK6uXyv8LluXxOZUfHyEGxGdWkbcA/IrmN9YImSVGEJTmrCVGPzBCJv9xi3x
9rNSEdA2AunoCnUZWl+1TJexU9DwfZ8M2EjUr0sJj1jT5jl+LdSJKTN3i/mQOCL9
7fvJYF++KVpEcZdUXm53ups9KdSDsSYkKMN/DAvALBKtW3IdGPMDAOuT/mHiQv5t
cOLJoZAPuZBBn9Ttx2VhGFRL4yQvL3ai7RHD4e4S91Y/VVN1H1K96/GhnS2Lw3SQ
GRWHQnKrrJtZdo3z/yoPcH4ejytZi5CkuQne4hgIz8aCiklKIfcxa8rJCCSTlnuE
HYhCKUiQ9CjIlNN3N7KRcyA/3yPKU4z/NQy06eCqmrGyiK//xWkHvW+8q7UDySkl
f6Qo3NbnG5uHsaQ41UZg2aQ+E0IncluaxquPyjYEC1dc/I/POtqU5iKPT3uzKv9z
mzk8A6ybQkzLUWfuC1hH9oBnPSkwwaLe8eAjqyUUJg3S5DdbUljpN3JpACXeInm4
iiaxyEBISS9J/PQdzuvtYMvEvNlLwEPCUGHnDlb2SnJFLtPSQx3d4eeBcFx1HzHu
nTk2a7ooqSZTUnhoguxkngKjGSZmn81rHt2lYcTZXWZfQsQ+YDRYUXo/Mnbb5s24
0UHcUGbx11LypNNLOHdNFabxz4Ngkg97zZt/vaegR6+y13UFs+CBFMo2m2OWLpIl
fWnFIHyErFdcC5GHv3NRJllktwXBHBk9dq8Ih0teT8UXgSkcexJJHCbjsphQiCs8
rNJ3Ic9Th2zavq6+Wv175OZfZTNj+Gs93KEKM4fFR1KUF6jQz/xGxCJVv5p6mJNO
G166WFQEkVZx8EfrumvFKB9gujMSfSGGNMudXhdeOpLpAkFeX/Bl59bUqu0vCH8M
Qetix9JTJWwCMeJ4sPe+dSySxPU/dexNGT0g6OfcHTq3ROF1ZLtdls6omkzGaA1X
guFscQRTFgNKg0t4nEv07V2Xs1vjnXIwXK0kO7zkoH1r3L7T3Ywv9yeQ5z2L3rrU
02HA0G/G7v3VWIh3IINpxdd/DnttrWrjkzb9Z/iRyLZiq0uUqmOhZ5/+E8c/aWXQ
5M3+e1P6I0A6q7YweAinlOKyb38+e0qjLKA2zyBTksPGZWck5LxMPgjY2mrWuhdE
nkq/iJllv57P1n+anRPk+7mVbpPSIMHMCBw4QxLGGdvPUsDPbR9sH/mQX5lpJA6g
/PLQarN6YsAshSC1sfIsZER6NVThFjA/1MZMkjG/zKWAJJ9ckwCTfWeK9IMMC/Ke
GDq7m9TQlq2V/F8MhczjrIOjUJ9Ekbuu8pxPkcUYieNnjKViAjm6F/k5g1sMfiJb
WVV0jgsbd+TNOk09hnt765KHlONuWOve9on/M5g0FWYlI2Ce2bcA0oXvL7sCicWU
ZQVqA4EQgOH/KgD5nUxgLLbhx/w6TuxwAa1VOnuU//DdirGiv+9wRyExMCOEdIEF
xhiLUAIJPj6bQbqRqC03GGqqv9sNlwg8biOStAAxkqLxZdPbJ4WyggQBnFoynp/y
eOw8y7h9NesstQWgfyM6KVofNazoSxEvBc9/om/r5eU0FHtWMfEacXCIGiF6dBh1
wzhAj36J0oSN1seTYlN7gop8CqQCAr+qhf64GlxmZ/cdDgsZ2uAO8C7BLZVxV5QS
W9Lt4hgdWfZJMg7TflVXH4OeOW+1hQ9YRsBc9l9k0YzCau/pbezycxE5+3k1wIhM
TVCKjsZbFA+CIB00gbCL+I07VGkZtXG8W0Y1iePykET9I9IH0dpeK8S8cZFFk8vu
3NTBnJeW1YjXpKF+aTJrvq/5wYqniFCLew6pplwr1gvF8krkkKwIZocfGI/HglVs
/r2UCyk5tEWKmVCivcYDr3tDuGl3n6cGG5KTeB1fTfMjuWtXRTyVAcGB2WP18W55
sS5yTGEhPhrtq5DEgiYc2lH8JD5lZ2DZPZpRocadEuRtKP9BbqSYu+uwI0Odo9jz
sHErQZlhPCMR2q8VGfs496MgUkplV43hWNZMtwqPMxVe1r+yG9UhoKOeXf6cZ4Xf
8JZUY13I3bHQJOsGYModujvWaX14astoSUo2AuVAHXaFfUYKjNsGogjo7gpgxjl3
bsJnW99Kg29kWE8LBAqDSOFne7MNkmSsdhBED5AkDGhkMKqdHRZf+rDMQ6t88ngk
NInNb8tzjNW+9OXF6SZoWA==
`protect END_PROTECTED
