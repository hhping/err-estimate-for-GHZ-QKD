`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0BYaCRQUKgDoT2UONfK2MlO0lOB/bZWC2bsdlFkD0b3iMb+UwIi1IegnJD9/5mRU
KqPT7ekooeVOIGgSOJT6YinroSNYn56OS84RW0V/nKmtH+1FzZ7UP1AvcmsLO90W
Q3DGv34Kcl2iOduMcWmjLbcx6JqGzxSyPm+Eob4mUC37kZ8byo6VwZ6vqGMpR1Bo
8FSHFFmTJYNZbLwkJy13r82QkW1/h2XFbR2ElyMbwDgd/0EPXY/K6g9IFe9vGXnE
QsecGZWWi2na5a1shusqfT9JrXotNRdMtIPLTKVhHiRTCYXNMvEr5U0iOTHIcDPE
8fPlnaWwU2hhPCK7Kns33sdmKPl6vQvfRUqyJ/eUv39kr6l/wpsR2cesOmqbstxi
DnkB61XuJEwfMWcFRfKOer49WQMroy2HgE4mBh0lGK+w+roitlCamGEceOrUf5pF
I6cJhlTKch0cljqSCZw+ue7NDJFOdG8+pLF6tZ/sri2v1C0eiauPsg/hiu1e8Q1e
`protect END_PROTECTED
