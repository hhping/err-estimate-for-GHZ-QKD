`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hYLYguAYjcgEE+p0VhckA+c3Y9RGadSXfTn3Vp6qX8OyhlqnNX+EFzSuILuK1YAx
2RCUMqWUCImXnMPqiDfVur4OD56HS1oVW2Ur0wkbGeqq9b736WWDsWwWVKLvWjZc
hSQfGj+Q0q+54FGXlj3OLqoUpkHgfUEySB2qmLtC1eTzqZpQJkmRb3bpWz6Fl7Zz
8EyhU/tGXAq80p0sETcXsJmrLGFuWCJq6vrsqM9EPd5CeR2B7fAYMJ/XvBcPbZ9a
K1IWmxuNfSv/CDarC0HxHv1W/+iQCbQl5jgE+Qm992Z+Gha35EB9HcJ8rN011QNk
CpM1lD62R6HvOsEFYHkZmcliFpCHArpX+ekdCBXIambkhYfzcrndXc4OHXN7fZI8
6CPG1T3mTYRK/4zehrCKT1p2skuQRySxRjdr/jBD6jy6BNkscwuiGH8vz/aOuSNf
arnBKHfvmO98OB3Nlz0e6SztBtbdrdI8J5XqG5yMwoa1KzkYm3r4F4++vbhMBjJg
ngxgsr6XXpogE9o2gCcomm27FRL/Amd2WvHLdj8XKChhbfHjgsL6Hk7lBIRvK6DK
cIdKHkua1oMHr47AnShMM1qf8c4dDEnw3g+5eIcsvyFvDBDHslJsfVQWSCqZ3tfI
rQuBrrmQMSY4lCssRdNe97hqIrextueIsNb0rKZhq+B1ZxXtdJSk9VHVp4VYmbwR
mFFiOL+UptC3ErbpURjKeWDFHF0efTof7z12j0X/SAKbTXfVuEwBAUaQlh5ZFr+4
b1lfDobJTtiXw5VFXs/TxwR9nQNS/zgZR2Tjau2kXNVFI7Xw9lsy1DDapvNUnmOH
ggp7rbWwYL94BK9ZVGlPIIJAtdbaPbW9v0LUWbWQF/4i+Pwiiu8eL8Fsrp41tL7x
qmmddpr01HOwABG2IrpPloPYdEiv4ptP0Fc/0G664ZJbCtsGDY7EpYcj4wgB65sh
CR0EJDgsixgOMxBpPdrcH0yPpnReTYm3H4/yQTdtw4yRAXkPvWNEGGwiux4gW9tL
vuHYcAvINxhncim+UPiztK0Dz32wRUG3amgfd8Qc6CXot7hn/e7kSa2lgvHse2Hf
pLdBlmzI1mS6NzbQBVT7eifCwgaz4JK7CWUyHQZTK7uKkxSpooShupqWL+u8hcGX
NxoRhYDpJL8WT7R6VL+BIkDalKxYmUPzciaOEY85U8Ffx1QdQtnpGgCcrGmKNgf7
9hIo2q8tvT58ldONkRvXe5zdsa+iyYq9XErKT1uQYcz5VzMbjqnDqNtF8JHZIiQZ
BhY2JPn+a9syLQqWadbnBotyeqEEw9Eq4wFj9aOYxL1qS0o+aBxyaO4jdqQwhtyh
70qgsD3KMMqcli5ko71ecoYDO+5SiiINDBZyZagjh4SXfEXdCxZ1kRLpdHUiCOtE
fwwwhPe2by+3y0DEwdmolfKlEi1SXQdJijamicsV6hxz6eWmWX+d+tz+LC/FPflr
3QlMd4N+11wzKHd1h/nHPNnRU10g1qDOSnmw03FN7+lVqTvxsWReJPaSgLyR1G3j
Vvt9uo3WeHSgKtqWmu6OvSfk8+vbS6+B9ILpOt6rSjcvJynIy1RGRJ9v1uBiNKd8
3weAU2CBdRf5yZFWEnJe9gsHfuPCzy77InZO43yeGYgBO7l7LD/9OfrWWtRyotgo
UiKw50swqP0rws/feMUfXtPyeHqhpapPEOx+mOCPNOrhsc98ur5A+wr37aINhzVF
0BDnLww2BAZiP2o7+ojQG8i1rvZXaIg+ST2o3SM40L9NjBqAcg6bgbkLJN9XQ1Wc
faLe0lAg1YgDOG7DwV0ynktbDrjPhigmgJrpvWOhXj+eYR86MU0sVvP4Mb6PRNoy
4CByLWi9Ii31zm9rszfqdDOxrSTm+XpFkMOtdyGoaF7lJYJEdJtH6fbnkjBUasa3
JRHY5llpeuEUWpBVMxEOrOp7u+pu7qWdMK5B9CvT8nfJN/WtutExhYyNjy70eCdF
Lg7cluJ0bHpBlRF6UVold6Vz3TbXieSxjtCi3Q/GHmFIAzCWeNAMWGsCu0ubHH98
73nuP4hVJXEDcKccKfz0zK34AgFsPBFxqy7kdf+iu4hoLPJ6unyzA9JfQqVljtSJ
p2eQOXONWI7eqEAnQggD0eoMZwAhaaOB/Y2AZwoVNVDtWR4A+kg+6rrV8Pf+bUA7
anIvPj0cYF70W0KHzDehUPC27x92e8LtKP/KyGugFweKn2B3iZ9es9aQpnB+6Sne
Ru28JGo59CC9IYganHK6iBYlLwtW7lQb1hkSIAKfmYPwe66QnRV40j/3SOn7eSzo
`protect END_PROTECTED
