`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZunlvPsNaKPCR1HOSPrXrI0u3rh3H+Q12LTLGDcyqUWh5D7Jqb3OzAEUSxFzvlN
qgLMe4/S/vAj0QM4kHHJfhpxurWOclGoWSU02C2A3LBeGtOsVcTue2L2EUPig5mG
9Gn6NZyTpRdWpdlJ96cHBA+29sMkm1PJm3pZkOTfar5n6CCjTqMupwiddhk6rlcp
jeZ2OIVUR4i/p2Y1pXLXJ13jSyj9lSpq9+n2fwsnS8SvF5Vo53jAzNALVcTFg67U
8AU9dlNtf1S/CGyYeRjRCRlddYV7jwDOTTBx+fHNJaeb2vBJNGgGPmcTlJ2EKwkJ
jY3BaL5eTOuvDjQlQaEoNLWtuYOYel1z4VLQ/5zpBZlV1prJJnvqrqt+7zsXEYCg
RU76dx8niC9Z8spVaoXktBTqFN1rfeDl4oUTS1VKYE9A+arlBxpONLhkWWv4THZo
EstfNT5hdF+GHbAD2yB3/+p8BkG3Hpz45PSvhRwqyCfbaKIMJUYCIklvA2DMNMVb
Zyu3Fdcmy12jul1saP2mgDekYnLL7d5h2KJlQ14IxWcBJWXyrDOwl5xwnOZ2RJ9m
AXYoG1QRJm7/Jwrp5A92YhTKVZ8D0JR6oXU7VAgwqo+YD4xhaWLa3nI1ZtBauY4e
UsPcRDVOEeEB8KrD6snmgUVyCostOMDYUdHNzIlIYoOtEMfMIq/WtbC3HeGsGmCJ
0ckDh1/uaT5DVoxE4JxOz2qscdwpwHVuR8B2J0n5C8pSqnULiT9NKWDaxg0U72y3
`protect END_PROTECTED
