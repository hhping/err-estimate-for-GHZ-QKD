`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMTHlPyP+CvCo7TF9qT6pmkjHD4omi//du+XLykblIIFHMftEiRc1uyyQuyLuhdO
gGBl8FKrXVTGUVS0dgp2MPIRhNDQmIb0ZN57MEGb6lxS0jDVlwmpaajlzxu8sudy
vs18FRXzr+r3rSwuJkeVIr/VU0/eXuLVbPtNvHzrj7dZmSeKJObx4FGyGrWi1PqR
THUT5EkH7/RXkXhBZyyT7vf5bMbRKrF68/0c8npGHPgo2K3DXyEUM2YaylF+zSuQ
wRKwZ5MmFGvYHp9cXpifleXSJLCcr/ySn8kfnIKrQJw5k7lFgY34+2AOCui7ODNs
FYFBqol0evVMH6btTBPZg2ex3OUKX9+VNrGEaPwV364mdVxrJNLgPHUmIbx4jlJq
pLwtk2P0NZRlCbyC0GLxlQDGEoqHvfxxI3iSP8kGJynak66+fm+fB7zD9xOwU1C9
T/O34eCI26Ob52dM6W0yg9YZs9HXARrOCqIiOpR1tMR0CCTQUYHrggleU9OiXbQy
EPB9pyzWHOJEQWoofcN3Ta+mxfnK6oM0Uq5pHTwLbg75LP5UY8y7HRYd8hoNZsjG
/nOuqOXqt5DlY2UyLUNd7Xzn2mEUGX1qnl72bZ0CN8FVF2x/qY1H/WyB7bSLJPPp
Z7Qs7AeVgKkRRacYkS2Am3ldeQrFEAxFo1iNxs0r743gAlCu5YYd3UeTOqvM7yTc
hR5UYu9ykCRs9e0GH1cnZQTUXMXq3xBUrU5UtLqMi6GqrQdBSoJXnLMGrE399Xwt
szZVpfap/qIO4LSL6kxu+Fn8Mvu42axgl8QpKS9p/mBexEifyZzgNVfpkdR3x2Jf
gposuELsF+4bSD1FABBUkpiorqVyXdX4DXB1oEqTKYxiBdSnc9sZycVM4ecQDAfj
9ohq+toD6KjWXaAuTL1oZ5H9LKjrCNcBSsLk9S1KMfNVrPFSvggYTFJP2BsS5Oyy
67ZAlrkaSeh3y4ZWwHmOlqcG1R3dxWuhpr+kGpUtvg9KknZPgRHm2yVZzT4kSpec
so+yjdAXk/IYvk1LTnNdU2G4k9gFPFipOFKCIzMxvpcizBey/4thbpy6uX8uEM0v
VAsUOOUiTdgv1AntjAYZO3iqcTAc+LVnVf8L36KpyVT64Nmn3vm6qMyilABPpkzW
h4SW1s6xR2kbRlH+I3MG6sEVNQvVrj2B6/BRoDcgizfSwfsj993z+fZosZaQMi2a
ZYmnrIPaqlDt8UY9e06IHhbDkKJhX9toFILpoymXaAF16ugGx5EfdIs3p2QWmMWG
BYwiMmHBnNNJrJCFcSPd48yA4pie85rPwc1ejGBe54y2ZkLfCgUbIuV93m2gmUG+
h2b9QjUYm3F7Gyu5JSE03tWjmc1YuYPxqPAwcOuIUgHEe3+meY+iaBKxz2ZKrF5h
1jJ27B5JkvLzpvt6cKZ/JiPWTJMknO2BUY929O+ZyXIhs9bVIx6XbHajs7OowgNX
tfAC8YO4tTcRwRSSFdWvz23wvHCtYmHc66vMZwWJKKfp2yMXmpshXZoYtT/Gl6Ma
x0QJAfIQDnSX4EhTXkv+Ri3XU/GRZhLhw52HwlQCbJDfSKv3JivWn/awqEKrIW/O
cPX3v1BQpW1gW1BN+8SsmtPB+V9M510V/kbqcsbhOGyqliEZeEW2J+aPIlKaAPad
svz0YISKCJR+bXS0f0uQ4PrE4pdaBCUpx0DxX0BFovTR2Y1HwCl5n29ljLyVrotu
zwoo8iMxXOt2LHghb7uJ+tsqkDW+7xne1qXQfHcNarWLjlzhiwqXbV5MnxNKNgje
pc6jeUAizOgjck5zLzHa849JdGTUKZrAglEFk/s5r5TtnYfUcjJFhOwKVH9JDo2o
XMq4vBpYRM2ac3XqWWAams8GRYCmVXvqzk1T9ODjHg1YVpfilZXFMFJLjxPUisTs
tlFxos1gYieCrCX5wXvhjf2Si0f13yy/oKc7U++CyHi1AtesgpU/vt1mSBpnmoJY
/UDl3pnZQjkb9x/njaahb1so3IcHSeLpmZV9LH2P7NiGxE0pec7lTVVkia3ZxF40
hf38rSvOd+Qw8bqjLQ9tU1ZN6hcJoT+Bdtue67+/2RucOFC3tbQDMp4f9+q013Ag
phbxwF3+SclIY5HMDPMcppZWXJS8hrcfp1scq9b589wAkIzNnsN2QaQrhj+DupK7
R794SsusqqUt8o1cGcNzK61HKD7/kzGytBGM35U8D8cexn/4ut5TofeEJPan4bps
heyo5rGtbOzMNq6VxbVLxLw48ffT9xXvDAjNR/4ThZVL29untMXJ+m3oIMjMhcE9
EDnsj9+GMWqxbaIWqYe1J8rVRyercfX+NnuYfXyQQeKxJoD+mkIbRDrG5PHbOhcZ
j84vwvOv2lyMyaTRpS+YThgJAqxbzWOyPcCp7mr8d79R3d2P+bq3J7tAazjCDHtL
+MZy7wZUz06hnG7hPgw5kWWmhjNh3BKy+ay9j/PhjclbvPjWOnAa9ke3T6GoRRNg
clCz+MlmydnnR1VBvOLfzKLRtU92otVvJdgjGsjEhwtJt9aJjtbklPPn5XxB4Lnt
OlZMSsJCcE69C4MthEkHyb8wqwE2fazP9EV32wAysBqevx08/IcdQcoPC/YuAzQ2
55cc1nnfgDQ9DqGBNvkpaYt52VimHhNeUZXNbDikMFMuTfg5ZPFVXWSjiZPssTCE
ZOQy7DoUkiqCkbOKaLDq+HMBDZiMUZqR/nDFN5cI4MPgybdh0aVwSJaZGLdgskwq
xxD2BV4h2j2otmCztQzqjsndN6DRBgYlCn9Z89ObZfgNSijV6mfbWAK5JArQDlpZ
mDo3JjrJJSkG4If2+qKNqiKqbxlcd07BrfEhqt+wIncjf/sLTe0s2Qo98CGXyLTk
jp4JkwjZTrE0ntigBtUcR0UApTp7X11kqG2tun2+vRsxSPcMvL/b2FaoBj8/bm3i
u+hCyRTFNECDnGCTS/Azh3moRgfpHEKJ4C9vPr6OJRWDFtZtXdS6/jvnSfRwkHF1
tQVQHYmMmFHY9P9xaLdbT10f9ww+62Bvj5vgzCkRYCHxNzYM9shNWM4hJWimZRN1
ntJs+iQNUIaP+mGCutIPdVzAwxt+DY0F6wU/H2/YexR8ugVguFFbifh7K0ke20tu
8AiCUnfn4FaggCqY/GxBXVh23gJPbzIGBPAUBxULV4rJr0M1Z8Km1zruHNHF1Ock
7Fo0crvnz4cKI58IAcMjWfRiXEi0mJ4tLOJfN93Ky5J+2HXZlEQ4Kc4JbOP+7YRq
X4t+9P+t+x/mfDcmOg2omAaSz7PcxGQuyg6QglEzDTIvmi+LrqTDhk4/qn6NLgDs
hN1LFxNaNPUTcbrceMnjYZALPJgxlYZYUxIBcdfTcGpEPNQfKMkPvTMCKbzKbNzQ
3W47wotjSj3VA30YfDvCE+8hQrbed1gr4gbJCwDO34NTp0RH8OT267csMAC4M1qO
e+qRZEVwSAJKBU4aYFlbVPBJVy/nyN3s5GLq7TfMuYjrYx6mwF+Ke+BIzh5jAoCm
G1sTef37sCbDJwMaDAXhngEo3Wt9nfVY0YvGxmZ0wyf/D+RJdukVurGtwm06UU1i
VRmhAul+6oCbhwIhGA1HfjAvPo6yz1fUrI649Xhhg0KMGbOZV/1kpzjMUZhYmp+7
Q8nzZ6XgIMV7cWT9SjbPL+dZbc9d0EClt4EaDjPdrnLH+g01tz1RbmFvHqF7KuRI
udc7NuhVH89B74HfuVZbODNXA///L7IZcjCj+UjfC5Tt0N5ijRWsgSxs3E3RF8gd
wbKX8lUBwnukPb+RU4PQKP3j8AGplL5ljSWEc1zm2isX3JZu4BT5u3szL+ge86D1
E/oyB1yxA8ToyVryBX+WBDjquSJtKCFV+48CohMyQu6Ojkigfi5tKmRbH9wtUNMD
vxlzvT0aSRwQbABN5oXgjzVsMW8ku2CqbNhaQvlYEXZlWUhMV0llbBIjuzksvfS8
z6FID7IVvMMG//g1kcRi4AXJUwSU0wSxHnyasF1F/7B/JQm/6T5yWbNLTfpuQ2Zo
HvABYyB20rQtiWmkgoRBzVw8SSKOahgnKQqWGnptuVcGJBFxexK6Sb+/As4k/EOj
gpeiEu8Pd4nu6GrqrEmocHlD4D1hDDZi0eRpUelv2RDO4NcpH462zx5Ob5X8Je7E
1yNy7edlj/ZRmnqJ1rsMXZ5d89eH2TqgNHidESfd+B/dv/5rqJh34HtnpisVQWCx
Qb19Qa/B4oh8njfgggCc2NpMEx8lcEfbAMV9c2lFpR2LZMQkh8pMopfoIs1uZnPE
Ff1yVRVm9/iJGkMiT6x00EuhJUFzwqWM2W2o5c2FTaIK73LF7nCGzB91/X0HQxHC
GQXTfq8B6rs+sz3kQN4U0hptBjgGzkSEoqzncQDh286T9PXTqOqf7BnKcCigXTJK
Q01gq2sOnQuaxOP5gdsr1dU6sY9Ag6xLeAE9u6bqWJPORDCZewv/pfNW+ExhsF5Q
GBLPG8CLstqWJFblalTtZ428NXVz35sPWkk9pdXhP7XwOxTrQyF/iMC3sDvbxIV1
yrcPHey2uM1+shJztyJRa8H3pQmvpzvqtl/03M299OPZ3jIC+QJ/IMKiqWbH5dnx
R3skEys+yH4s7+k2i6dVEREx35aTybmu+kIaXdILNy78zNWaIbxsdkAbe/KzJmzY
/F8r02cdGFST2wmZ9qi/WKXP8xvYb2lmhMBgtsL/+hwqhkWL/JqG5iRuauHJSjAm
owUFtbSIeHX/rQAg04Ex8mlvwelQM5imdvPKtWYZZxA0kX5GdWEbsUTCdvIAyY1X
0As7ySThJsT3mGhDJ/v0ZuVmQje381JjUxTGBfNaPCSW6V+BL/i4mphpjRR7zzN6
kWc1p7ZcDiwBv7nPOingvyKXg9gIQeOlYwHrPt8Mv2UssjScvjPkUyOkhrrcZfG8
edi/72bgOnoVN27LAWvfePLvuxY6LTFoVow4rjVDOE6NCxzKnLvfHRxMGZQLSuBa
O/wcjjTbzbhZUbSCLh7nh4lLPbpO/ZrcrTE7wOcHUWUor3K6O2RU3EBdFa5qtOB1
5tNHgqdAPdly0skbLNxevqqf2Sen8rE2H83QpB5eJ18Xim3b3CarJ9hltAA97NTK
NTKcHJsXMZ0SqZ8Z2AW041vp5Qy65sdaCkaZFwEwHEPdoci2gymF88SlXvBTS3VU
L+sKqgb8rsHsopZb2n8AeONYLQaJVseC5VKWI9Bo0BXOFrXrQ+4f3H/qagD3GPhc
OGM02GI93+kpe87YNvcqhCDQYWZKruxN3Mw5Rk/LMHRwjPG1gKD7zydXpqkKL4+/
tJOjnvpPQ9nqThEGXcta8KNuamHijYeAWgpKNBZlY6MWYnO/DdM32zKlE0VeXCt+
6dB26nqcnhe7GPfZptiUpz68oarBUwQgige/SkGKiZFrqgMuNU+9cdhxf70wHzpw
YuqPTQfcU9o3iyFihO9ENNiaUswUDH28XUMKzj34El0uz1bjD4aHSBy4j/VORe1U
UpyFa34FoprqkrDhbh61HkYgWw9B1LJyRuzC/I4Ob7VivM3A73JEH8b1kXNyhqaL
HLVQV1Tmpzwhf2YBm0+qtK3MxyCY9b8OUUQLsfoOS4pgqplrSSsRuBBqaaSGhIGk
v3Hd/ysPj9JHRZCVgFlXad5wTyIumKYtSPm4fBdbEEYxPg3Ge9eYpWtZhVtyL+YE
zMdHMyfa+1SkVOcg7rP82gbJZ2xxwnhus0h9uHYotxed7tBqvr+auiS/ouPW4Xu4
SvAdD155/iamtCpAgeZ/8+/J4UZ2BjgJA1XYCepIbqfay/oQJRJGAOMQpONO4q8d
OTcnd9ILYp0nojS0ipmixyTm+TC20sp7Frymhv1gaCmhfODcNM+7UiSNpLj4cKaV
75Ec0l2d/eQY3FlXvBT2o3hax5n3/kUmxCshhaYwXA2rLOorwxoDwHSBrlYaDYXo
Ftb9iGOQCvf3ySUDCxGMgU53/i4dyEDzGr2ULgozpPqN1Fw9MsrpQrVfINT43R8r
4Y3O086HNOB3HY6zhITD0j7O7yTjwuGuNV3DlFrxtIM+CwUzT3ujyDgvJbUB+HwX
yk4qjh9AHr5AYZWdqPgHpMbTrhOhII+55dgJt+DM33x5XIi+YkiFVJH1hOKBhS5i
phlGurrsqvb5tiGEbK3FjZLMJPvqLowN0EMpyqQcim2OC/tZHOnRWYgrPBMPDVmt
1Z0EljaOWp11ZL7c1c5ERnvTIsx3dJ9137vfJKq77bNoxkdlRlwC9mWt7gY3J/bc
PJkP/Z3tWluJyaM89smOWoFgY3we5WnSmHBnhJ2aZzCvDzhdCweJlWRopJT5S8mx
5pi4QdiWCu3RYOZ55i4VqTtHl8AxQG5t/wX67iDwkWm4WHiSAGH6rCzjbNdFae0M
EErmwergbj9JOaN3b02zDHYIXRTOmKgLwYWycCQQgwNB9IFC65DqrfNBPHT/l/qd
kXw1TKRbOYnHMK9OaE6+oaHSaNE8yzMMd7fh3bW+JZ4qWV2vP1N2VteZM5TGt5xj
jXZvwKP0PJIkYEH1NFyitBoyqsmKGWtft/KOEGXprX+tb7bPdhrD5Gsnc3w/JoHH
JG0cE3Z8nuCgwT8M+t4Ih6/TmBd7Immffk+ZUUH+NienpWVvLGpCfQ4PrdDVnM32
fdlwwWHhSA9JKVIL/R/APWNUSxh/rkGyph7mIdAQfqZGpfZBU66rb+pypFBQO5yj
B9KG5su+9cMpGe7oa/8p7wpXg870g/+1lsxCN6Q8zToHq1Rgnxfgk0pLNl7Yuy4U
UbHo8h0G35WO0G07ieXCzceyxBFlIC613jAi4hyn3FY2jsHTRb8Zj2CDAnpwtbbd
erxw2OnDQOri9rw9InVbL3A4IAqZckD5utiZAN9LqL8Ca/k3O/faCLq8EakNSa4r
50oQhYxDnXeV2U5x0P0RCFIirNSiy4eU+dVyccHrHZjZ6xJq05PBapIsZCDZ1JmB
hMRBqXZPkvGTEnu6nHN58RjtlOHgsiK8MFI3PINn11RUUsIqlAMzsXiSWaJcUzI4
e0II4s/epfBiOkmGLQHeeQgYEvDggljM3keug+prT8zY8xBZEmI/QylXNM+JMDO5
AO5dsB/8tsfJK1prER/qt/dWDK9W/sNg3xutrSIwW0QW1ghP2DlpmtxuxPxvpEUE
/3YDeTOGoQVXAx90bp/n/GK/AE+JNscGR/MUhBZyc8M=
`protect END_PROTECTED
