`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfBwAc5WD4LkozZepbwM1s69G709LykyXKyHIWPqH9VYA2rbcHhnXW1pWdxPQ/ru
XMUhGLchXHsRbbMQ9chpja/mZsZnGKc9BbjJgkZQ70B0x5waruLJ+n28Tgd74us1
+pWcH5CSBs7G5kKupI4IUlEP45dMzQ552bsBm9boTMhrr/TGuIpXnPP5P1G9/Ydr
dxybO46pUA9CxgSlqdnc15GQ01UFTl5KRuVyOp5nyN7A3V/5TUIi8FZjXg8ck43X
RW0KMcC2jL+9Pcu5Sojrmmfw++SgWcoewJyS0V6TU1ZY7b1Zs6/sOiq7IsrGiKZQ
TTIvQUQ5RRNYYpko22wirccZe4iz0FpzNsgUclS+VJLMt2rTic74U8I0mD8FR6ES
`protect END_PROTECTED
