`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0cvGeFNTU9K/UmXVeA4FcyrBOGncZOa+UWuWYyA6A0hhDEkf12zHfbwFdpS2TWaZ
awTIXBQv7tTnIWysnroCqT4yWSbPjv+9uIBwJTp0z7FZildlUC8+4mG7+sJjQjlA
hxBtU+cqrx8UvqBX5SymLqr3ugG+a1wGTdwiGhTiSVp1rq9hnbH2FjHutEuGXuhj
JedhX2XFO5gv9xu1ByCfUHfV7PaCxZe9ejDTPf+LlpRiMk10NhcQxYgwXspCg1VX
3/7Qz8pHXwRn8rh8NBPFwZ6m46v2lGeNBGt0mgzKlZYvpzhQYI/SDAyCmXxFnBn1
TjezOsl+gGT3ZyMtVoWjkEs55wr37loRha8i9au0BagYJdRrvCRITGs1tEUGYYyv
PW6/l40BWxB1VExjYKjXthKipbQyCOfJbQ6BDAtzL+yevB/eP/rYQ102gv1Pz1b0
6GTDZSH6pQHZrfV2QRSsgZHrtFV4G2KQKSFaVEjEx8o51uqI31vyyuLbs6aSC21n
oCqxhVbZkwcv/ARpDmBhvazItcoYJiIO3DXJY3d6gWLw/GxuaiM3JY6ab90AMr/T
cCPHRvbfVvMvGKUiFQ1J2L6KZAav/XVeKQQpJ3Ts+YvRa29/vhTkpXpQ9/N6rpHo
CY7xj0VMR0owGpA/faHioHr35+JQ1MPyWacNPJsdbl8=
`protect END_PROTECTED
