`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7XG4hXSaNwidkJRgufvBSXFjatvPF2iXclPfh7CggLEqpbbpFci3dW7wElHDn4z9
+V/l/8H9SUGkXHoOITS9WSorT85JU3qcSS/uDz70woaaSFJtFYFWpSEf9+mSqSX5
51iH1T4XOPKA4XjYjfIyZX/DBfTkcRDyxmmDCM82GyRC+n0HNcNWF9vXdoe+wwt8
3GpSIrxu0Hm10mUafwi2VQ6gaPjiu4o2IOmO8lj1KPCvJcQ2lsnqz5j8pQdswNjB
SaDl1GTEBgoez2wisJQ5+AvJ3QHdnCLrpJamFl8W/1ZcuLOFHOot2hg5YmjMZIIM
zeeXOJRrF4Q3LoFCAx5YeewNE9sTADYN1moWR939o04Kuh4iSO9YLETGL2396K0V
zve7TeV0zxAQk6S135sw0YmYRPreuSfZqT+4TLYsLei4Vu0HIhrGxxlrRzhDlg+p
8QbwuOHmNQSXHLcreRl1QxO25ZzBFtRaJ/HXst2qHWlJ/R0aHqRMzNoEB3xGIUo6
EK9fVH/ywxQDRVlvmYZnYnY3W99tuzGQOlkXQ9ZLeX/YRu2pyebisLWvYtV96ssI
QudvqawuwvQ1fKvRnlP7d+1w3Sop0gz6z042Npqi/2uXlELGhJuSxHaE5EFYFCXf
I5r59L/OU6pTvwPdHfbTGkkLBJ/3otd+O+k8A/4gVynvN5Eq7lemfw2adpgG6m8t
YYWEwgMuMYrEuFSPlXia28yLXw7WexTy4fqGcX419eCwAYz1OZ9UK5frQH9XEt8p
7J1wyczCbRasNQWhvgHLd4YCRbNWBQ62ojVTh9twtTU=
`protect END_PROTECTED
