`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BCZVTDNdHRLok+6IDJuhyBr58q0DWpSkLA/jgsivFrKrhD2VhOgv0lNOiM2dBi9z
jU0LdzpkGxGXVZUTbgRHipnVq7ni97Te590FuEuMeszDH2qJxNjilAA8RV7+j6cB
4bWI+VtVXczIJJhd407jDrJAL22EulU/gcNpD3JKZv9NAkcyMxGro6XXYAqOTy+n
hSRwmhN/3pwRsLZRTmy4C11JaKEvctIgBvbyt0MaUUdqc+n7mB8Llv0rTTtJHyNS
pCZKiV3ZWVRFQTjtpdAKgW4fxElr97bSoahXVZpKDnD1RKSThKLaP5UaKCW2qCSv
LM4NF3t/K46PCl7oElEkY67T8Vf4WOpWTJAaCcNk5UeuBWYGLyEXFkNjemQ33LBX
o6S8+k85L5I1mF93qxmXaRc25tYtHpWe2+LlDqIdylUcv4KusG0eZAlBvR/XGOnn
XTl0vPZ628ZfVsKvPC3zhYvRxMcO/Kt7/SgFMHVQ19RjBvZSB5FBmSO106j3XCH4
PrfEIT7cT1wj8vyylcg8z7fVIqyCGMLkbHUg+Gc8+70FcHiu/xyx+WGx5T7QVXXk
3zkC6Bze2iW1aMajaArAJJVwrTctILt9NfFA65hvqakPbHU3/Oe0l4uqBIOinZaC
Oc8d7kjSlxZLVu3JpPnPhauH3TG8eHmvRH7tKmzzcojIiEPUfUDp5SrEVnrHeMqs
Z7OpTLgw884eaEhbDBsG1NgupFTWzGQDAx5Q0wx1TWfV0X5yaABuQWmoznTHpqC9
gOqgOtxKDfOnvPHM3peTdmXvpNCVVhKxesUEmwXUvIE=
`protect END_PROTECTED
