`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BT0Cl2ffqNyNJOGhkv/w5TPkplJhwTrI5491P4yeTigdI424fuwibL9vtaffGuXR
CWJU6pfivV/ZU5XTxkKne4QxmTvaAft6NjW9Ilga8gT9PxXouD6SQBKdK8McDJ53
7rLXYXjABdnIdw1Htda5SmnJXEcu+ilPQxAkSvQia4WZ45fbQVqCRejEMaae4Wzv
q3U5RI+sQ8cnX8SFxVcN+mkq/PALG9ZfJU+rAotgkpfTKnNSwD38mMnJ0TmZbWYv
Q7VhiwA97c1aqyda+/3gznOYbmTUvUpqR8hneX9o0Ro2P1ZN1iTj4+FqA2vqUFlG
xXTx8ej2ONWyPmmhK0dt7STORidMggVDY0S8bJkavjOV3G1v03kPI0wpEIcY7wZZ
z1pb+xKg+8TkbJoweqsI3sxF+S65KQFqvZGun5ByU+7IcZkXNDuyqdyDjdgCIOyL
sa1HSn28kUcd9JIVduzYdi2o0uCBtMmqFjbs7tfd8dbFy0oQkCkQgYMSYs2zpMw6
/a74Ia0A/R7u8fEumlUfj0j5w+ntTz5W3PjPkHkOVioyfm/o2tVgTxviP5DzV+2b
OZ5rOjASWnqjXnXHoc333fAL944ggp4/f3KMc3e80M0=
`protect END_PROTECTED
