`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1fT1lA/MTRhqlP5y/tHrVbmTLjG3rdSp3DIwoQ7ILm5OSyE+9Al8zqf1sT306xA
/mMxiQvGljNPHRDzMrxOZ2dNOQRjTMYyIlfhMAgvRBDwyfm9Pus98gKkfdbk0TOh
gR7cQTse3Q5935tOZ1Uaw1n3S/BC3GNUc5UrVMLEO3Hn3k0ZAdjydaEIiToWYXW+
FAjCJafWMqXyreQS+5kMBwRtTiKN/BcFCfL0S/PYDLi47js+wO44VEZi+oFWVQ7e
39xToPbiGnvi3WSOBJEbaj1etIhxS5NUF1HmXf3hbIK/nBeU7NWBSJx8tXaAgsOA
PZhESIc88kXFWaP978qQVgIOU9UQC5NAS1maFoH/kwxkaKCFEO/zlg/g+CCY7pnS
TcC3yeGH8ov195cADFfcPiOT2w3stGRWkeX8GrLQKRc=
`protect END_PROTECTED
