`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3S2mkw4sAk/Ulrq6oHf4xvPv8cjO5HOS4KnOZ5/l9JMdrL9K0NgTZbpB+9w/txt
kUacjO+/I4of5F0yxeNZ4xYuVz+biD8wdfeXB6pTA3NRqg0EmiOmmPlUlLc80CdK
F8G8Df+ROFX9AvnERioXL8OX5i1uiT+Eh6LtYNW6vBmL4nPcwkigeH7UXSXbYuYn
9jVVSK2Uu5WZOR7EfoUmW5+LszbR9uijFu7r0iHOfeURN0lx4xonswP3BW0qQTXc
do8kRPt+QQKFIYUwoq/d7/DlphuLIS9r7JR/qUTfXTL1pEIpwlcuKa1YBqVbb3kE
d6RCa4frEdKwhHO1QlmboWHj09CzbMFtKB6R2Sx08GH4EN7zmammoVktzAdDGM+6
pCfqYtQ/tSgiDCr8olQvad3ASDx22WVisbv7NpIATbnXkojIbS4gCCwsPH/Q7tao
izwc71O7vIn1K0kY+A/sM08BKTHHs4M7Zgy7cQsGRhNpX5HoyywbY6RGUwrbL354
Cg9Kz2ImCBfMUUrmKayIfmcic8ssKTXEpCu0LMej24zwmZXdrR/2rLvTMgeiyr1T
0ZZ43Bj9gzD0d6xR8KDWGApNidVEu1M0/Ar2rBfhiHzFHzg1KmfT4yzIOk6aEX7a
lkJF9jux0yvvxJV1MaoABIzd3YsK3FO3UAKB78dH3ehOVISRnGmPkDeNTLcly4q7
7ykuZVS4OQklEyrCqdbdi7JA9OgYO+UPDE6R0tNrHRtA+BtnCl6mE3r3quAQhapV
v6bq/OVAe+/ZKdH2I6cp/bUeiwbf2wSmoHMcw8eMLkQJ4hZrHkAqD0OB8rt42RDS
zRzmKHABN5o2JoBQRgqwUGj3D1O4xg3YSKzZp/CdE63H0v3bKHQFA19QMVxtc1eN
hmrvs610T3Wld7MvvWAGZO4dkkIHcCkQ0eoH/SKdWjQjcaRFDCBig8Auh2F6aepZ
qKaBsU0ijm4BHbfPvkHoL+XM5BiM6hN/O6DqPz73BfjqGb9uFS7Cc02sXnHfcJfT
wWSsoT9MWs4yn78PNtwPPTGsP6WuXeFywccRWpGkUfHyLCVBHPT/fGHjRBqfor7k
Visdr+vs7dDjd5fd+R3o+o0j5AqtN5I9nkHHMWUR6itMJevnI4k++EbEb4I7o+/V
5XEcWTiwY0tAgHEMOXRwUP44q5EofJqYRdcJriELQLvSCfwusb4Ll0/sBVU/JPUF
aIVVnl7/MythDMve73sBCMdq4FJY7zaf7GiA+wDQ5yVgtglabCxvQAZWD/tFXnug
R0X5l0QcVdKJ9Fj9iax8n1VWQ4/AGV+/u1xvgyeQnU7XSgbZebjerkU89Y5eWovb
MEI16Uz0DwlD8l0ZFUh+jdubmQDDLhdwdMqRHmNkBVEUv8atnE4llx6XX7Evr3lm
Ofy88WmgwGXCBeTn59ZZo6VrTWkk2l5YaJJG1Uci4rDTA58qOmyN4rEo8NAF1rbI
l86mHNgyLBvh0TUHRRwK3Di1uO+GVgj7AvfmLOTpIyJ7ZhgnLlMyUS8Rs041AUcr
iZ6JTzoN+ScXV8R/CCIBQBjBoAxvhJuFjvfcJIKD7SZcu1zUcThU3eyQ/EnH/jRd
A1kUpLISb213MMUj+0e8zkWs2dPYCAHEGxLsdWoOIFhjVotvALLx5NjMmKNwcEfR
KZJdj3ZBe/WKtj57eFogOFS9694KSqj7iDYkluQbFka5jPdq25VF5pdHlgP7CxKc
G6FOAb4HnJLhkWjTYiwBg13dq8zAUYq+IcpBEIJJcMjQs9Aj5LRQvKcfULogHxjn
JrHvMFQKndDj9ewHsTNN65avBz0EH6jZ+m1yx0LrEo5R9AJbrRzvQHQDEpzbE4jo
jNCvtbkAT0HU88V2VGFgBYjDMyeIzlU09WlgHIhKHi+yhj+7qNHhyIewmJgboj3X
UCn0UuwUgH8lQB0yGBwOVOM9ioFLiE9G+Wo572771D48pTG4XX8dHa1nZW+xZ/KU
ZA5/QxbapfmhtNpNm44A8XdLSo5FnAb74Jfje5wWdldPZ57h7iH7j4JnEImykKGv
0LAlPrGx0SwA/jR3r5r9Jk+jhZthVWAsaJpW2O9kzf7nYGrSFLs7v3GhhvVU2yWk
Ue/Qx9m8X1kd5EsbchzQMBLgJVGj43l/shByEsDEsvGz1JVdwS5K0zN49hhLjAGW
xBbGYTj9v3czndbPT8dKwRvv04N3CIPCm817oz0cOAFFDzIK4ZtfUj1Z14tlFfe1
+N/UGXBNUNYj9C1nTo5dz3r9TDestuM2z7zVpt2HUjC3doY8GrbJGXf64nZA8Byq
J4z7OgKMWZ9tdPX1NXp8/OwVxDeqfNUVktTOT+SMhWM4mKlPPv0QPT7hYqsHWGv4
jlkqUFKIhPqbaIrRUwdFzPkxWpJ4CyeZ8r+a04i+ByvPu4E1fXLTUNIdgaKT5Tsj
8YAB1oFToDaoPxkwIjn+y4iJIWZsij67VLf4+Sjc8kfjXwOFnssiYSO0c/b6jU5g
dSAV7lycDqJlYqAhC9J0mVc/KXkO2DhD3xOOCRE6HKKytS5MpLhLPSbpAaNksBFY
VMzeEiCc25TcFV4BQySluuO7T3r0acE1292ynNKrQ33XHlhntv7e2AzpJ7LvzxBq
3Rq4ziujDqLh9qsmqNg801JbIURoteqDA3cDxMXVSgnvDZJsil7vGJAW6tQUDRCC
TpPJs33BUuUyc3XK9Oem4Gk511b2O1oSYcydiJopJ+mn4+VAAwlIO/D4XSa+BHf4
P1ME57CmikGxytmU+3u1UEQDh9XTgCT6VclB/4OYJZQPU88OwuU0LzWmuKFtpPbt
l4aj48T8CbIAeq27gd/kMPvLa+w5pPK0WwCCoaaoBlMiop/ZD34AWqTQI64giagd
8g/fT/qWTd+HUWWjpoyJ8jhKkiPb4P8UeQZhpDyKxylmYITEqWy5BsY3Wze1Gg7h
NEV7KDXV0ntj12R7iv83lRT3dKN9uDvI1UGcSqOS/zR30nP+5XVcfRYqzoHj5MBz
hn1hHXk3xNHLFLD3Kd2mqKSRpkn/YC+//Q3y4yQDIz2zIHQu/ISCn+sKdtcsGN/o
beiHSyw29PYevYEusqaScqOpnpVT3+K9hjyBCYVd/QT7WojWMHnQzkH84Fakbfzt
B9t4jZm2R1/lKEcGCBDNk+8y/JCPmcsxR1Ve5m0Tk8aSAHNJClQqoVGVDA3SJtAa
kQ20rXbnnIHEdu/dIuAr4/KP9jKN5gjFAFsGmNswK1jYDcCv3fXvPk7sGqia/L79
HjqmMCu0vQ3SAmE+eL2JFh5K+hper3QU/oqXB6gdUarTwZk0++9Lu5N+fbQv0Ba2
DDLmpeamhJEUSE4vR0l2/9DV8a5Q0ocfQWk+fjEQ7EBfm28msVyzBGRRvM8vPDFK
yfMT5Mtg8Zwt3/zY0FdNeM2riw5IBs5rGYOcqqjIM8pVq+yBP9ZBMgAIu7NKmRdX
zc7hRdaa3Yl8C+SgQGtUdc61fLKK6Gsz12Jr83pTEH/kHqVgIDXyg/3TvSLiAU6Z
gt0vd+AWAWLLOxrolopEvcL1l2dnW4AytDwqQ6JNZvp8XF5NOAhl0WiV1AGIQThP
WvGd/Ku7srUf8NhYEjLAdBIeRSgVmsdHUKfH9QiG91hr+M7C2KoEI1v/Cwyq7zNw
UkTXrjH1kq/ieiRznhWZqlqwp4K99Qav7fioWANHHRE1VHcFAPGwWXcNubHvCl//
FHYJgcvf0hqzqcCBdZyS8a8N+gESFDO+H9Bun8IX+RvxCiWO8dSVqzMw5HmjDEBo
VFaJ8h/6IsTEK4Lu7OJAOha48Og2zI0kEczKE5NXrLcJVqL3QbV5yhHbzvfP5YCA
9qWbKHm0UzdAAcfJYbdH3DxQbZ5Lh8fYbHN9AXN0e/mUR10mtUaKPCW8dBSpu1kg
7BVHxg8E7FRWFFfKhxXAJe9NIRkwM/cJoUoYxrip56o/YTaLSOoFLqWKr9rab1N3
`protect END_PROTECTED
