`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EHzX5MWuYjDEem0AOfvK/ID0I8L6IgdY6UjJI2hWzodnrYUHdvEDYmMzFDmry5m
O/G2f7g74Yud0cjMg+VTUPPje6WbDYnPa3IkPPcXrCrroHUV327ki7ZMLCzW7/IV
jh+QId/deeoTceJlJsDG6D+7czVb8s4FeQYut+dzvNOSyVcEXvcV3H1rYNLqaBDd
sr9zPaeaPid70H+fS/GrHkkxeMv5KxTkdRIA/6Xuv5NVFMgLX4QVZCRkgLkArG6b
z/u7OVuxXH83JYS3lsWEU3p+gNKnC4z94ZAKVn2JTf9XQydALJfXBzT/i4sgos/I
K4MuyYiQ9gwaJ6Aj9eCK1zBOZ47ZSNf05NB4AAhhzUVscUt38oNXjgbeXRawIz/J
WmKxG0upG4vxb4IBQBV6InQ4cAlzE8xw2pYHQHNuiWiMRY28KRkdI/9hO8VUBS3V
ky9dXTWWXCQ9FT605euOChHNfBt7zRDXOeGaLEfGKKepROtsAvVqRX9RRP4zj2dE
+G1ofz0c0eQBm3zzbGHcKUxMjUoWK54qm/BXDwJeI7Nw3BWNbgVlZYg1c0a4Fe5Z
ZF4IsDrc9PIYJo26giEDbpxjZJZ18Md37inV10rvOa/DLeuOiDMHtcKaWilZ/RLl
pGPJxRlFbSbYs8VsP+9lEfaBC6Neqwqk2rCnDzhgu38Wx1HwgRp2UlmZkVYVfEw4
KBjhdLWzkKczo0/HUblzM698rNceHbPDQAf4mctyLw1/yqBBdTyb3VFLpQy0DGPG
Z1uBt51Sh1mZX2DQD9/LmNZrHnlCICu6ihvzS/6OxJB9Vg9Rdie0iCTM0ZhbkDi8
gCaQvRaRy0F5057XtqXRpg8OTPh6MLKBdHAhNVMwOzwgHjtwddFKBPR5SXlR9U3J
OyzvuJ2w6wdAGCePloKMZRUf9NKThutXbwpM1/GJQ1rlPwpEIYjKaboa8xeDuCx0
8BnBdgbORU6zsoFlQ/B+DRISeqFNl/NPR9/jtzHqi2AdiPAyrN8qtLaSjb31uPk2
xyZVoofeaE5Cc+l/SLM4Lb/M0v8jnO8wFwREStpo286KVmNWp7gR/CfzyKIO9PH1
9feH3GHvxWMlTtr9INuZiQsALxdM+214f8sXDKBdLwZQdB7l8Wwu75xSl7Pqb2JB
7L5WpwhNpLWz5CQjPL8/ou61MixaLdz1jVXJcL+NVnfxm7DaQ0gUD/R34zE0qgg7
DZVFGauQsl3JHjG+4J/OLZj5+n4w80nZgVg3D0hXooc3EPVutjQMcSD8RUJ2IY8Z
TQdZfDm8rhL9QiDR8uR64W90qq8EUH8Gzh9mmeWa/U4i4s9V04fhrN6dU6LCX0k4
5VmRn4ImvcxD5GcX/uVhEE3gb1akVIw05a+fRx5gnyUzW3XrJRJiB29DJpHqQIcD
hCQ+QiBLoL9kMK/XhA718nuZxIP3F3cWD2sldB0XsGJA8WHnitQZsU/VBPExuzeC
ud6LxHkZQJbTWeUoWzdQFtHCbptQe0nO5SPDXR+gmzSspbH6+UqFcJPF4QDyiUER
gbRZkO2b/+4Ljww5LPBBIawE42qdaJtK0t4lKY1LkAHm04bObKHlRu3CE6jGroFQ
x9k0+ZtBOzdzPbawnUuzpzFe8duv+zcwt3dTHuGU292+tloksXrmRNR9BpLov5Pu
LwUs0TNMgayVjGUcoa8c2ZAVCxIt9W+2AxGxm1I0WCXLiENfecRbRHl/EnDBv5wP
JgiBiC6TEE5YMjb80X0pSTcfE0ZwROgsJ+2HnAYUr7e2crZAQ4PZm2W+1vCsDBD0
D4E593pjsKSMRB+9x9XpsVgXWTu7JHHur4J0iEg7rNShowjwyyfrlkYsL78ZmQ1H
h8jxuu1hA7j9wPCDECan1xi/5RBLb292Vi5uNniCSknKzAho6924m3FBNHtW2S3V
7cF/wlSByaY1twK8D+GP5RqFKW63K1j3wnOMz8IUeVH2jGJj7nbFz9pl3IW/rEsk
3wKhB4KvQKRa3WsnD6Q1MkwbtUiCXz0wWSFvIFEA9M77686zVzjWTUCjN0mgf+JW
tVl9uLnze25yezXMmjgzoSYlB22P+4PbYkms9atp72OpWEek3s/411p37NViK+Sv
kviCJqgtrQSHiBHTWmM8ijyKJFAldQdUilHb1oSxKAv4djF3cZ4e/o5pCD6IOckQ
MXpYw+TtGkmmWdlYqvoAhQONKBhRqtnbEpAh1vhsRVa964YEkRJiLozXZbb6TKrl
tZx+vAt0Txu79kiKH+gJpDKCXEdYZrCPYbGgTL+q/xarMlUiwdQHXWf5+b+j8fMw
rtQ27fdwZ1UYQ5e8seb/eIU9JBgVpalo3qWdZffwKEc7QyXWTAVpvawYOKQRX304
fnERu9FbJ7O33JzRRzMwz6mlxwWDwcQm7T1Xq8Nl9thlyysWLHkigfIM7JBQ5JyZ
Pkdybn8nW3EuE9KNqysD4+0pENAC0UfR33ZDyM2kq0g16eXMd18QuiVx4eZcANw9
puBInCs4EN2VwhAZl47mhTjnZ7RJBy9vvN6YAbuenzxDsl5tGk2E+QFqfLT7+kJN
`protect END_PROTECTED
