`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bP5jrIqgRWpAgzolh9nPbqEv+g03mom+/jRy0PEEulFdW7liWwsUxuEMn0pk8k42
RlLo5xhJpgjogDN6iDw8tBKnSRFtnSaLrmL7hnnaOsDMuy0zPQaGNkFQisI7GAqU
DGGNbgGJ+L8CXuQ7R9VZQVlS9HSyDX0UyN1Y2HFbGpV9pPIgOm5XG/nVDRLYSFde
EeE2wYUiMEhz4iG9B5da4YnU0ugI81u/KH180woIKtmym1vU9DUeXTLccnY2w+iP
BF46QiSknUTzIsv57hncM9vaBS5FomfNvGvGmyHtpccTaIu6Aoy93zlbbuA9LDbI
d8fhIrR/gAv6XncYL/Jm3UCQsTUspilGnmBgTKU44PGeHuXct7g2q10S636R4/N4
iujn58/5DfZY0O3Vagi1LQ==
`protect END_PROTECTED
