`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/xLL1maBkcARMQZaVH2jtsyd1NGvlmfeSVfXagImAGo0XTYCReLAkxCRPq9JntD
ZmbcJnec6gp2nTqJWnPGj1FS9+UTDUPKnxFDtTYlxIyKWrAwI+ansZwL/aTNny0b
gwb8r22GkKAXifT0i08VIyNCzMZ4jwlykmu2fTeVZ2eveFTi6Ao5/PJWfpWBN0lO
wN8UHhqhAeQi1DGSSp4mKVBj2lsWPKVjd55zh8ZhVzPjOo2Og7X4+0huRCo/8j5F
kz/D4clbBzHx+6qDYg71MiFOFOpBrGVRT6Ou5QhIBtRvHOFVoyghdsGcZl9kJYOY
UgTF0iQ+z0OtiJWzG+2DMy9lbjyNZXOa9ewLiVomtFjvaK78x3QcQp8+wITwQ50/
POAYDUt02mMqNYXDXgWHDCiPS7XEqPdhjsnZcBuSkqZMBj052aWhy/Qv92FnEssd
X3PnE2VDZGazImT9bKA3Bw==
`protect END_PROTECTED
