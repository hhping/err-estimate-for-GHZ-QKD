`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jdhDyddsjFI+NscDsKOuQgYOzddweqRb7gBm9kvKzduSQ+Pn3L/zwqGJ7HYxa074
WrmcN739PxchI/jLS66hYzBxyEL+V27DsUMLyHjvJ2PB2ixcBCZ4ue81IbhAxI5T
RB5+JP4z2JF01aqt1zVSmyhlkDD5SH0i2OYrEqoErLb+E99pzJJPUyz8jFwfkJyZ
A9ni1xy0hlSHYtzdGDvI2HMj71VtnlIiMeiIIam2IZ98Wxa9I0MtwSpCJNNKSkKR
A/bll1/jFJAzDcdL/xy4Q4aMnfsYKjJ+taQwibCXEf5LMwNB48AvMxXyaAjz63sF
8se3hPijQHVruSDWlnu9rZ0/gkbEUKqUWWNts7P7OSUHY0+BtIIRVkLR0r8gBxLF
u60Evdi66GcLBzHh8B/aLkTX3G/t6EnxIBfk53Sf53sNbwvuB/NoOoersZQ3CGGA
qqOT9TtOlESFFEuFte4JXaZWpjtBq0+dJdTfMRVhT6PIpnwFzdYFZxrxM/c6DkPy
e2jUflV1FST4K8FS4YLb5sbjhBkOxsl8yBtmf8MweTHsY/CW8l47avKJsat01GFx
GmZ1Gov6hcF3j/b2jOOjrOYf3knzJ9rks7GHnv4Yp0Pkhe4hoU0kGmffKaJ0htq+
O5rrTh9kHPK8VPqiln1cE9InfESnrLPnOqFpcr1rHA17+OMjdnrhPLWfVmZkHSRc
HTwwL+64n+3zabajtr8OEb9tuTK5VZAwHyVDOUa+G6F38j21+OjbykQww0+8srYu
yH4cJ5XCun/e1PbH8p+7J7Jxl59Cm2qvZ5tVsnNwr6PBNb19ieA7e55b3CbIxF6m
hnq8m2SXfjVMNPyoLOmjlZHSO2zZRcqu0Gq+a8q7XliiFT4RbSMve4aHFQ6QAt++
6583z5qaFhOd5Vy6kT/eg+Yu1xXOzRL3FnBeUSZ5jMJMknwc9T4FRxi27OrdvrsO
+WaMm1/24HA+ia8sRHY5OH9TeHQiQSDAdXv2JOtrBfZmzjnHC8ZgxN+QKknyA0pn
b7aM/ASRGY223RfLkhQazAWM2RCNhpoIPfqTEa11LcN2Ls8NpBNEPao1KQicufM1
bX/a+7KfTZbYzgfMf/w/J9n53gDtavpz0iGVXxG/l+H9Pcs6YUut/sb6avX+O+Wx
rjupMnT1xnI1hsUsHMKc7SSQeTin0QwQHu1pbl4pX/HjZMvXC1zZgPTu9Aa9zxcC
NzBr/cs+ZjNdGFyW9ihjOTSaSP4wswrjOTt6oCCgHyvO8IWLHMv67SPWDB38E+Pt
bVJ2xSej7JM6w86U5qKrc2WOE1TkZaMqkaS/s1tUmVVZO9gTRlNJIEmrWWObyJyZ
WBoEBMVn5bfByeoypovG2wXpfBa7Yv3+RpJSRl/+HmRlhK3VPV7iUOPDOb+hyGp2
zg8WJ8U1JF2B6x2JHl9ECIaXvSq/J+sj5EHfXiFDqEmOmTmS5/N3xlwz93EP166r
W00CYi6M8OO/JRNKP9WuGxDPhN3nHkyVslaf3ss2LFDDjNImNtpLQeC1ZL2xU1yf
OxnA/X879zTCfnV1JlS5UiwPLuplbAjFv/q9z9lWd3itpukD2RF3brUNrg+lqxyV
fxGDR6dNILw7kdLeK5ETROWkI2o9lrzRc+X3UQNGo43lhB7+AHY04LXC3vFn33qE
vWysAZSMWZJ1FU7DimPHuO803E7aebhya1+VuIzMutvwiAFzCgJnteu4cuGpmqop
iPb4uMYVAZkVNHnMPcXIuG+yh3wvdncgqCNQ2Wkjrp5wXSd1Ga5UkmAwdaNhuZXa
YEcBUM37NqhAhebpjw/y71z8dLnEvq7r1Fp0s6X8+Y4xfZOM9qF+4+zZ2Z/2h43h
093tGl2TVlSCH4Nnq/ewZieF5eKKdsiWvFBu3xbfRyLGPOkM3ig5CykSrCSPlQ5P
KBAtpAKIJgRwisa34wjarPH3E9ki61fWZPo/29jExT3PdG2gFng8Cs76ukv8p64b
RIlImxJliOr+1fazLT5VZsOdi1qg9R3628ejZE2Www7rxFIyYhsFi7MobL7ycv6a
NGuS8smrFhJfLulAX2+gAc6R1t0yiOP/zAYMNNagPvhjgeHtJD/gAgudeKOKfSkL
ULyVt09gth6CGuzH5avYOO+8ob6B/MCxE8cMRi8umTZqJty31W+RXOY8iQ/wE5za
uiZemXEIUNgiH+RZtORVvtNK6wo9UwySeDwnEOmYbFY9roSy9L5Rcx/Or1yd5ivq
sJiaDoZ0r1kx8Us8/rqKNzXgJHYNdovMc507MpJ/uwq5J36/DS1IpGCsw8R648X/
8zu0o3L4O3QjeXAH0jFHpvIED0Z8EGHseWuChyise63Qdzs1+R3x/tVQ0XmwtOYC
`protect END_PROTECTED
