`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCLF5WMsaAyD0/xNBFnCDlY93RG3YLzwhsUpuzYLKgwq0BIbJ5dqOk0akeWHg/3n
6Hb/p/f6bpBu4JQwhb1MKin9wldfkGGY+v5MAfP/AuvjoX1Q8MUPxf6lgOB5U/mu
fMMIBJjv1CAl5wS1QMK/RFqDSI/ATLyVaTAqwlHVpczoVR2v1AO7V+1K/XrboFWw
R9Z3zk1XHe4Fz4zUd8O4FKpk59F6VAap+0CYabXPlGg++7T99rgJ/AsjtWIUGvyf
g6vqtVtPvvixxRr8nfIw4iZ4dup6QdUvdne9b9mc7NtuUdsYf9Gw/W1MYAwiFoTZ
OptgGNPFUCzu7Q/hiyecjGj+oBEdfcTMLDRDoOITlPvsXYpbsI9sApRsmVBAsSuk
8y9JVNCUVtLQQfXqTRqKfsuXHjU80oBkzTg3yK/EitLBMfw66974Ff4MH8ge4gVa
kuOcLipp4627fnACeDCCll0T/A0IRj4aZpKoBtXECBVgLV2zuoHfmDa0VY9WJv+h
Qlr3VRgYsCBlXUuglioKzJ64QSBK0St/YAgVbtNfdTjwte4ELLFIOsqckD4aKHEh
N7aGWfZsUHQRRA29OnCJyDi02e9SOrioWlo5Pn/uuRmc7/YkruBlwqaTtKjGpBqy
vcL0Q8vk94IpTeXEOXa2nG9OFToTB0vZthsMtX4tA7F92AHTHovfQBuJqdgJj13s
JAB55PyTbinrPHbT4lnUJGrluLjdNP4nOzyhD+SUHTSRzCE8O1q5cLDy5GLJ4h1A
DWErlGsaPSgz7bFWx3uyFEtcSbkURulYWC+aYY241WSaL6Ffj99VXBobHpxLnnqC
4OMRvHuLNIseRxCHwG7Jnvo3KM6PeKmZuYnWWGG99qnpAIW2SarXnoY9hIniONQ5
3FNqEuBs2piGo0krEs1woa9WmVZbNUB2kexQV0Uf4OPx3GTA5+gj5ngn9efr4jdS
8NE6MDhP5u3MaADC8ftJpChj8bxUKjDF3ukwBxMLUQJP13U1/h7MX30omezbesga
PxNjgjnXLuAZftVnQlyjKZNR+SvJwpDyYeXmgnxqrHJ4d9uXD2ceorjLi3CPCekJ
Kas3unt2N0Z3QHI4l8wQDw9CSk8gefsh6apmy/J0Hm4RrJFQLgAc4aYpVlYTImkx
Dm8l6UY+W8VEUy5j9mg2SxCSpmwuUEm9m+yuMlVzXLUECxfpl0EQqSDgBSCZnRPw
TiX523F6BfWAFMZHcm8S/53G4ftZ0cLfY6YgFwTQNRQnuAhBvGM+48HGn2BCMw9r
U1LRwu7c0WFOfLKNVCu09dZrd/+I5IKUOWC/H6JtzssIqMmOu73iLMhNq8ZmoYgC
VKkF3kmpcc9o2AQdCTWm2ynbJzOR2NVBj1m8Y+Zs5Im/7PxEaSok7EXxAvXfCHWh
uH1JTaAW7tNFJ7CDsLiG36Dd7YZkPxWXwPAfrSUEFMHvKY3xvNILYlqSyU1eyKB8
knLPWXKoD1W3PS7vYTLiQudb9lm/vic023KTxVACLbIM5YqR6AJ0BQ9Zb+wm1zb2
xLZOl4QUjMyjAdCfj2a+bjeExW7lpkRBugMFYvbIv5bkvKe6pn+A+k8wvIWiKBbs
+F1BcqkkCvT4kvjFo+fVFwA0x1GaHcDwQz91cteNbF0XQ9d+wHDOBBP6+ZLP0B6k
nUT7+E+b2UNHoQzUdwU2+VNi3hVwP+G/E+1P2PFu3A3cFsCcvPdp375EySPDnI7S
JIGjeBKAQ1s31TVlUAAPiLWBrMC/WkJZemJHrWhQ0UF4r+2wecFxSx4NsPvRrtuM
s5CmVfc9EahtarFS4v/ko9WdL7iUDtv2ZAZOU3VnvQCHosDNJbutfyI/qybX0A6J
AvFSt4ntquat+KToxQTNuZRqWQqhYU3fClUad3/LkOk8+2sentQfe3E6YsuZ5k5T
+Kmo8pqDklsrpSTFeNbRcaksxpMscGsZip03nP3gXTTqk4G3dBo1QJ7SQjI6PvYJ
SC9OiKEd3jvu3fhkn7kSUQK1WLlJhLPmUS2NropHDI+oGQyhXLOJX3l9gWS8coRn
FaQ4njUEQMzqzBn/E/vbHqxb9+Hp7OTi63FRq4geGn5pyBH+JIpUHSEbh3h12XQt
AQ0BoB3kfCWVOD5awIHL1jdH2hNWA8xkPX0BLQ2uB8mQqm7mMoALc3fc5Dz19AQY
MqSzlehr6UJZf/TlHi9jDzWSAQo42Qq4OKh18Wv8Ma7rXcDYSlMDn0gMrT5CdLRD
QOUbmRhQfCk4MakHTdr5bYVikH3TU6RnHAVHDVcCTgwlz/dRbhkaMwyruh7OdX3G
sox8K/iF+sQAWNX7PjL0aevF6RZN9U8ESC52k0FDETXkwyVF9jG9zCQoYjuCN4Yx
csYPzKIFZHGIxxEUE2z9Q/B30cFYn8yYDjP7MCDLpmqjRgVdWYJM0TOAqOuyqvqw
0stv81eKwESZD3/UGpMhyuLgrHKDLFPZuoyDXmZmSEkW9yOBR8R+U8+74N3eD49W
Md3rV7Oi6tYh5rMeupE9CX9nGCgqVUXQyNf7NX3CN/N8E1y/dK7YSil34Wdcka6x
qDlpvdiX6vlaHk2/l2B+P+SKaRO4qPsvFeFUVjR9qwi10iXbnlupISN9tcyrlJlf
3uNBeaO2RcRG5Sg1cP1GorP2LfCa0ceGPpPNCdPa5nmbalsxZZYyC33A1w5HtKLZ
DaimPG2gL6ddLWQhLfXPdq52uK7vGPST1jxO5BMAlew=
`protect END_PROTECTED
