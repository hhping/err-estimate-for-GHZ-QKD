`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GmagoNqvhxuk+e2S2s21Gy3+ljFGCcKKAaGffIXb2pzsmxttFdv072ViW2lw7kQF
pQCZtl//tmeMzH/WblC6BpTzg4SR/vPanKFlADq5WoyibCziztKakvJ7OxxV754f
/US1JMFqO7AyM5CFxym0FK9+SYsjz0CilzNbjGkC0iADArq0q1qLr+89skD1GoTc
MpmBN6ND2BbAeMDSF66EH5Y5zEhw3jofyf2WjJ/TVCpLM8PjkJEh4OtUevGdaiM3
iv315oKexgaI6Z2lK5sgRZw3h3j8q+6s5kXGuvPsXzsoJag98dnZVWMDAaNt8CZV
QYmokxbu5LnQPXrqrzqRAJcUsEt+lRT3udksq5PywYTmJGTw2L+CdtoQzUNXPXMP
zWb5kVJBwywEkQoIYb0LrAnlP6Dy9f622SOsXX93PKPgoo0sEfnVlcw9dP7IPt9a
aoDo/TsXHnVKgtaPLTC3oTtoid6HEp8IhySfQcsZqzOg3LknBGIaUBRDqYKmiZEu
Mn34xp+V+PWOct8e3k77BxutoA081tvRWbW63fpdc5y4ORdMOr0JSi8S8CPAFmju
AmRIpsnroSODCnAAtxbxT/JGXheFzT56yh9OK/O0ML7pZvYwcITGx1BvX4wxsRXg
3ltkV+jqtjTy1SW6BEY47vKFlTtz0nQRl86My6SiB+/bW7ESfYysq3oq97YM16IQ
dTHzSRr4l005PKdapZ2lqXHIHoj1tWuNBbX8VHkeqWQ6Zc2GWjSrywR+ezwBHum6
ds360xTZm2ya1e/VKeTO7w23EGOHs73W5BzONJIPvFQDEPUX4FOQ1qag1ErcJu0/
X4raYdYRUn8NfkFJk0aj6C5ETpIbbdirLhdZbR7m8oICn+8DGMJNhNnuxzD4d16X
0EwN4UmsbJW8HX1F/n54FQAOAJDv1OaaMgJbL9oG4zuoh6u+n+4cUSM39AuD8ua+
MfWOekSqGResKZIw/BhAyiR8X6f5gyOQxlT5gzkPTShuK3HGZCcnLhc5098T3pIM
rwkLE2eb8rOxL9y5rg00VIpE2AVUqY6LmAR7lmCq44hn53fchEitLjM6gRwVICnh
Kgzqy+nunrZ54mlaz5J9ZU8W8HhRI6jghwEQpnIFaQ4EIO6z68k1nkDJXvkXRw+g
SbuwgcH6UIRctwTiQxseE8ce3lzhNWP+Fvb9uL0/eQBSAEnk9DX+TeuM5en4abxu
bdRT0gVVWs/UTOn4+5h0vUkr2T6dlPMUsXPp9CjMuXEhtOHRS+SQffHt+C+cY9mh
zDH8b6NR1w3Tu8Az/fXb2oEBnI+a9+6fvktBbP8EC8nAkKSt5Lsz2VRaf8yvo+bt
N3XoF2ZZnpYzQUUtBpphkaNvUQjw6F/Z2JdAEHZTqCUb+lZmlfyqIdM0ZyRC+Buc
tlEPAye3WbBdeqpv9AzQ8IItatPllbttJup+oCSpzlLud3zY39EfFGsdBE+FdeG/
KxNDVO+2BKsiNcvORx6SwvhLr7aljK1FfBVfXXuqcmdJuXNLNi8HxJaX8PrhDdQ+
oAw9b4GTpZY6H0gi5ntVogA+BbOuBPANmX/t8xWL/GBws9J0rus56kVGg4WEAjze
KDxnBkWXy1f1ulYomXbmhk0hWhk0tCSe/dack7gse55nuPbBJtRc3MJPC6fJL/ON
EoevvFXc5I/4/JtAEKTlKr3nKGRb1osvYDU4jG5lOiiSjD28Lln29CzB24PNTTbo
bJoqLemLEJ3WFU6TEmsbRqd7Ju/9yQ0Vypkyfho/OyOM2U9rmgFbJESMayO1vf8W
qYElIEV2BGi0GLAODaJ4d8kxQiN6P2WRUZjAuscu113TMrtlF7Pi4JQEkXrrTw+8
JvFLnb8zVr5Coa66SjBKiqMNROA8UGFR7Hj+DDnxZFzjAEcIkFql5TNEFd0wwkgq
SnhYS7PD/9dQQ0FybQPxK1+3gwuEWzqpm58Ypy9QW6lu+Qrdxvkly7W7X/hl4ebz
SNm4TW5YJdSnLFK0dQXOgQfh+NyV4UPmUc6HAhr9Qt3wKcc/afNwhAqkrdgWsbeh
nFJPugdjrBls6nHsUf53V4ngBmjZChqU+VUORVr/dfAmpIZGtNFfuYjjn8yuruG8
bxfkH2rOPSdRc73pskr83GTHoDbL5SMYkqGjjSaqEzZKnQ0vl44TuRm5IRju3orN
Z5BMX0Yc5uygmw5btC4xeIsfo60PGKk8vYo8ty4GalePD1gW2RK7YPLyUAvgJj+B
IE5kCqYHJa9FNhA4ZjUz+d7ZC0SP27GulsQOEvsgUw+SlBnZUc5XFxfmgeWh89Cs
HnZyUnVOP3xCFFUAFp5Nx/Zaz3LQEUMTk54VdTjti9nw5mo1V0eSdQrafuM/+mqJ
Z8ophmhTtZpArDlbKbNg7ukoxfvSTCjcbKAgm6zlhTZs5o/bZRpG4jh7vHoU6fV4
zsZJZL2R4guPv/d6hR6CUbDDfHHjv4gCEPMkBnB8V3DnnXmg5wH1sm81kAxxs+vU
YZHWm0REg51e/uqfOGzUTKEtWrfx/0P5VL1JWRBIrJHBpJmAKLe9SPQuy3s684d9
u8mjwPDaYMO4/mBFz4Y4Wmh4Rsj9ti7rBHxq792dPWJtkY9ceqKtFgW/WNnHDEhx
vRMEEwg+1UMm6rd1ioJZTSGpvF6Gk8YaNrXnWxobPAM=
`protect END_PROTECTED
