`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9EHJTaWmLzXLXGxYDE127YACw9RqEU1R/IzxZhKGMVwHkEDKEb+etMk6bPM1177
zXGTn4M+r1T0Q98QEzSDAgMJc2uAhbYlPy1ztfOszys7MwXif/tdIhx9OevWR5J3
ofxOJGbIlQ98ZVNsGc7RkRny4HvRcFAXjWr985pzERrTimPNJ1ALcMYAdqB4eZIl
zUeRYbmDCWIpxe0NmU5GgLkmervaaDEKz1pOyH6jPU5k/0RP1uY9fdqccVqA5qhg
zzVDFRVW10bb2dPdk6ZjL/KjbpWfrfVBQoGnneqIsFBxgsKtXhcpLXIM8Prq+yEX
tzGMH7ZdH7bNg9x2jCSJ5TGjoMc5XPnUdqbYwESrNpiQGFaxpQPv24s8VZfHvIPw
1c8hPxRSkptcKnckvXwPJLrPQVPuSivId3I5CBPHozjEWM4T5t+VlUztbiY3Q2qH
Q1El+w2DuAIFKTN7k86Tbv/uAEiMl+hzRYhN9bE2+zUzOwb0Vc7GVVEiv1T0dM1x
E51pBQQyiJz/b3RdwBICo8AIRPuIgXWGqCbBNPztx2gQjQlHDI6LoSVBjoUkte13
VPgqBgnQN+hqcdGPx4KpQxWI8omrNpQfMOFETsyJ66ve01DtnDub4YEzy1AUZ5yU
ME9jdBcGCFonpigmz7Rp5cjdEEZuBUBQuzhvnyy37wKe9dnbf9U8yP2PozvYhXSF
Y0LZVyeMaWb0JHLB3MsbN5sSDDxt4iKQ0q+D+rNv0gJ2rjM18rDg7GFcLuR6FnGi
MW1Wgl3UQTpqkg9/r1hlKzk/GJYssSfn5zQpqGNfwXf8sMuJIVVBDzVEG0T4ArGk
vmU9VIg7eEb5MA8vB1kR3vP/JFv4vLpGJY6UaD1KgId94huGQLY4Ibcdw673CU3U
IfC/SPqXsV1O7hhgv95N3+FEPlEgq/T4NDhcGNRUp3y5KRuiTwYfG30LloOND7y+
+PktjmJ10oyblq2cTl8mmlr5GV3ULUY0s6B5KmyQABzUck5pUcDt8zQiYckroOUp
8O3bvk98TLq2wgD8nP5tU1lW//ckjqA+DHk2SD866GEKgpYOIJH7kr9ezYIRpPRc
AJ0r4+nm9R+3qc/Fn6Dbs1lpngDvHs4cV+oPwUuIWdI=
`protect END_PROTECTED
