`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCvx/HILEDmYj2DgoU/brtSyIzMxI8V6mL9pZDmG7OXc6XxPf6ct4LJRAEb2wc5B
GEsnLsffq+AFaqrTMyWkngYi2lUXfjbBuk4kJRiDkD1zBLicxPoO2RGxXZ1VRJaD
BWW6NI+JXsQGvjRH8cRc3My4zqlOIySiWiFJqdX9zXGeLE2ubvQj8J/671abv4si
3HSmBvfFcB5dWAf3XsIKbvHNve3EUL5CHG/Tx3b8oGhXmKzohuOwxsw8hijCx7Mz
fqFEg2E+ZrG197y5O2XrvtMs9HWjONnCULgya0IThbRG9nfzAIQMLrftcN/PhMrJ
N0sL6bd30/JivXTgeoQc0ofrmVyZOCcedERVWXWNJrFTmQolxKZEDc9e4+6yqbg6
JK/v1EsTBLPbVYrbEduyBGNBoipTZqmF/pvCH27JK7n3Hrn745gpu8lzDxNULxBR
RdKg0HPjQQD0Y4rN0C1lBHe8pG8xOrMtWVxk3zVcZ9TquDqPxKz2tG/T8TXkmu7X
6szufQ15mGg/PE3kivcbMyKnot1wkmpTU8O5pFADhoPN9S/+8/C7bPcAiXS0FYV0
y+fsHhsHO9nlfSDLWN+hPhZDOejQ4PGEfTC9i2JWinHMry/kChLQTJ2qXS/vkQI7
hWwM/qeWP+37xS7z7jYmJ59Mrt+pIFLIgbjDHFAieK0qlefX6UQpVNumkRDHMx5d
Knj7lPT9WegRgoR3bVgHVYkheiJR/EqIR0v/2CugtDTjR87hOPBYK52Qj3aBrB/H
`protect END_PROTECTED
