`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JGc7j7zDESeOIi6UWeACflJZes//YeJeKRgCeDI61XdxfFi7SbgXiWHZq/pU2A2
Wi1Ae/cAZLu5LFZPuGyXe2IFiV+Q5WXIUL8QdDOMwge+qxv5tIcFTShfrIClc1m7
Pu/o/liX5aw1gN1L948uKNTH8YugNkRzru0FeGKL61lVdcBUzPmJm+Q9zsMv9PSh
AevFwwM8JACuWZHGLjjz/VCVVK3VZ2ceEH+V8D7pJZzBztGC9ZezyKTb3wf85QEh
WZQ7FAp+Ru7WymUQE1QT+erQAjktTEqp5TRKJwtljLVmGcGr7nOTyTrJMzXjGY5L
wrwAbWsX/0dpOYHjL2e77x1dBfJIFv1w1tLC7Z6k9xmGUkzRxor6/64rIS0Sx86G
qnCtSDQPkx2lR9Lljc62CktP3LRMlhCjIEOFSjPuez4dvKD54FLaSySkpqcdC96Z
i6DcDpBBXfftV7Ay8yvCfNrH/WN4LTwBFlvUpIGYCI/UMW40gcvWKFnWu1M2tEQf
0NaDgDC2eoTRKfJTziCyKwE4wTWq85ogDL6Y8ivWcgDcPDYbEaD+O69K7lmKMTfA
nzOAF8hDCpSvan6NRY3zYlw1NQJEfU2aGocb7amxSwG7yvH9eCTEWuxoPHBTw/YL
cCDtfT7O6wINlXVb8SnTQbkMIUNE5l1AsqEwPSOP3op9pNS3m3Yc5uzC/ghDka78
WsYA7KBBkBo6yyYFot6WhSiuDd8oXEZa/TnJ9qiaz859f8R9MhuTjsartCQp1Jkw
B7R+EXmupyU/2G7ILuvIz8nhydzmrHlQ26ieXCPNv8d4Q5xRK7eT/cP6tC2ZtrTO
ABH3pR/ioCfoiCL3HPzxYryXNxOIs5wHNgEyfc+0Pkt9ThOCIsSNPeZsVRgwWu2X
b+PbeE2LeTF0Bd/nQCzKKC1Ic6ngr/UdPFcx0NgwrhVle3acLDLA3xCa2t5YeNCw
j3UyeGKxLtqcTnKJjNordG8BiQ37vvPlQzcuhArWxUo=
`protect END_PROTECTED
