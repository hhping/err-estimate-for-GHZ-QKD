`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0mUyJVq54Kx4NUM5urSfFqy8WKgT9SNqdq/y/36IlI5v1mL29Y1LxlGB6Af7QCM
DuJDqESPvi7XJF9Jnvy0s1mX++pcVcjkaDdK9eocpoRWDa6GSZgEUA3sfjYWfvay
do3FO5P2yUU615Vb3ukMclw3eoJzI05VjRTdwNnQDddFC5ysKB+EplbviLq70zKj
dH36WKjdFR291adlW4EGHzZSra8rMmU5Ua/RT/l07zMeZsir7z+1jNEnJsMXClEi
P1Z+Yi1C8N/QSC13vCOvHGshKlNHqj6ehigETv43qRowBBTTEHqAJFomFTfs9nVD
HfYX1I0IkAG1DqGKtoIt6j6bN2zNDO4v2PkXTuXtLxs0GAi9x61IkaPWssIF4+Bi
7/+HdQOWAWEOH/ZMWZJrgl6+539Vk8o2zLkugsocRKTTQthvIHBGfNW9Yu9cM7vp
QCnAtudBo4ZJOENRTKYJPEXo8W5LAcKjTcAFGZmLd/ptb35mvxIM07xwslnWoqUZ
6SPrqsMAtOpgQV7Ot9NutQ+hIBgOTL1D4Vcpa/Hi2vW3eXss9PiwcmAga8H65Hw8
AXzqXQ6J+s+84HSTeXTm3r/leWK9u6z7RSO93T1ahhhhz759+chbAlqmdI8xLHc+
74sZruAgfmwL1e/FKXJBqK3goosjEN5h/+RljUTiqqGLLA2HNneOQrmyX2j1xKMg
tL6hC7e4xDIPSTMMMgm8aaecU3j89M2GiSIjRvYRSH4zH/6IxJVoxztezRbz8mZc
EBUcyzCtnvOOdD08OnutDK7znYTkHAyV1opVaEGHUOssg8MCp5pOSETaISksldbE
0xCRSYXwcDpPb/+vnsltx/N68QSpjjHOWs2x/6+bLwrDfM7JsIcAsWfdWoNZqtwD
2o4LhNb6HJlK6SPmp4NvNu5JDYWn5cC/DXSUPl64pg+KxOAGw5UWdfgYEaeu+4Eu
jLMe76EFvSxvSyddEGJBgj5ObpBcWzhnhrExAwrWK1e+EFU7k9aYN+oeajEE9UX+
OBhuPzf5iuRC7tRZ5WPUCRm9fPie7cV8ko7YozPgcoze8T+FsCK9oElcUk4oHcFh
KGvJa5ondOUsrhn3TrNp571IbEdxry73IHVluxSUs64=
`protect END_PROTECTED
