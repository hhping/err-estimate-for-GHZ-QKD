// log2_single.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module log2_single (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [31:0] q       //      q.q
	);

	log2_single_altera_fp_functions_161_kypxfny fp_functions_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.en     (en),     //     en.en
		.a      (a),      //      a.a
		.q      (q)       //      q.q
	);

endmodule
