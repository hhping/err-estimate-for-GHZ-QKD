`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XCZ3rmLgVElmKWdH6RSLzFEq4AV4o1mHfmDiIU4c2U2sX3xNmMCYa/Iyt+Zh2pLj
hJIrEqdAEuWlbXKjJyezYtFeT6GjVlEW2dRiM4YdTAUNqLdT12Pkaxx15j5cO6tg
VQQf9C9RudxPYktRA60GKr+6/Ms52PCQToGXT6C1+zEKtYF6KXD4sA2OC4f0lprq
WVJHniIZCl5GHpIYJ4tXVvyQp4p90iaw/lssNI3C0gQ=
`protect END_PROTECTED
