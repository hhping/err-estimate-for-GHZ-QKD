`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuJg58dlBUEHRjH5OjYjtuLMItv1AGcInUptAsWsw4xzstUoHuGYdYIwxTsKgmTm
vw7OzoEhnHj0L7Y8aVoWxgbsSMLrHFEFE3CibhgFvjuyzZqBUUBFs9a+1QQZWHxZ
goM9F6zRAVeNbkNg/5rq+DI8QCeRGgC6vLXDdrQ4pSUOz9/xypvxuTjyFUXD4OF5
D4x1+M0QGrkzLuUwk3QIqdL3S2tikAy7FK07rCoGi+PwmO1QoXdfQYQcwdtvcJcJ
l8iLYZAnIVofPr9L9dJ0CTOnCE/YIFuuSNnq80F8evvBVNkgM9SGVU2U6x4gBNNe
D9SXJTQA44lv/k4Zkt76gnr+r0lgsJ/gdXT02LRLmVk/jaIOvsqW6lJrLq/2b9O1
F/3axuenPRKuNqPg/Uaj2ToeqcrEHgA98JOGlji/OQDqO0VC8Y2Ig3WxVIlzG+tZ
PIktOfMA/iXudXZngU8wBIZY2fpK6yiDfsX11REwsRMgMxwSwoHK1TN0ILWxI7nq
6e4i+Jbe88gw2YX3ztIr2Pbl/5ERDWGXf2n86345O1QPdPdbCTK4x9zugIJyWBrK
3OZsai3FPooBfF3btUAXv1BG7/H1clLNoAF72qYGrvpepiYrYx7DIdOnGqUHxLZe
iJuWIQaRS67p2I8rG3Hopoo2HeSvmPyEB1jEMo7ijymQyL2htfHkOUwpJDpIw7tF
wErUZXtx8by1m/2agmXvYWUych25//lV39J9PmgD+7hVoKyFzoMdWMfO2mN/ozG1
`protect END_PROTECTED
