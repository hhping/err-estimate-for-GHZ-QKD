`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9m5awMFuL1k0ChhnyZZOko2YMxkT8lEoRjnDSrLpgcJde2C3l02QKL0hKWmXrIst
z1RDGI6eR+i2w3P3hFXoR3tsvvM7bzdddXZUEoJHZ8CMhCiP/QxygnCl7z7ZrvSa
P/sec4MRq+rO3Sx4LYVO4G6r+2gUSGGaVTfqVev+b4JYzgt1ah3ShLJ0dkXGiSD0
/5zueQTn5ZtC4Jp8EF35wEqjgZodIz9GIclw+6xQFikeyYEmXQaCzRPLMiUIodHK
prZjylQC5J+1NkN613dEza5evwukzETuxg/rHQhltoTTHp/IvRgZF5oZy+WNngyC
wm9sMl6M/opb9zpnf7SQrUd8vz9IQlNIsu8c8WL1W39VBuHQLbvU0+bC5Mj3/EeY
LbtyAZhKGvfPny8CfvHslaXHQ4z9lXuy5La5jEpy48NkMbPhJwRKw1qgIOpKlbdV
oy7A0CCmcwYGMP80FWPXBryiaGtqZgyD71B3FeRifB8+7jtvMIKce9qNGoTfichj
/SI1NTEcPJK3RxhcMMPWCU1gBnBpHGJwN2J3dBspevLiOFEnIKWhPCF11Je9MKr5
VIJLspFA1KXdZMLggBoYOw==
`protect END_PROTECTED
