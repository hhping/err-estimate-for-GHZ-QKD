`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdMVvq4aR0pG05+ZkvoFtjjaAvqp2SlvtJdby+Db2F7MNNEt1NNQvDBDw/AtDvWy
zJ7mISWc8Fo+aNCkDedjcQVeVx8B7Cq/ZDb3PrFXSrEAXiDWtiwarKOw5EdNjoGm
LwMijADKAu9VgLw5+Mehvnp+N9A5iz1W3d6YJMe+jBl0Zy43dUAUhJug/T0Wc73O
Si+MDZ5+ajFB/pithmehwEzoUAkWlm6SXs/oZsTLjNc2JaLGui1JehH3qoef1CXl
h+WGzPCU4P9SM7tfVRSW1BuqzbKKcZCwIN6OhiWOL+rlcroVCTgCwZAXYJ55UAAS
4nBhGYxfwKKCH4njASPeflxO4O/7gZcbfqhPGcpiRwsqcB83R63hTVFUgnDrBig2
In+cYOOkUeP2Sbchkna9BHztxGtUD2KN/csBBz7vwLaRBt8QpBqm8Rq0+EiulHZ/
GyOXCtC36e4GRqi8e7muRdE0bWOvvfS37GVl/ChWFsLDOR2BJVOvM2ld3ur3MinZ
xHMkrR7ZlqwBSg+OvDZeXMg8eGT6U5wrjiF+7AxbCirAM5jtAJJFxIT+JU2xYPht
Rb6ryzat0fKVdjXqzRjDgEgZbnmXJwTSaojpkQlPLi08mPKS9UtCQZ2+Jdxjzj9F
FXUqqvDOmX6HoFwWlyRRsuP476EkFVscAVQ4UNTXphDOWBxYlUO+PGuO/WQtvpLK
M9/vd4pGM+zA4tsKw6vj/tmzPEJxVNGI1J4nyNWMLMT1S2EWn/hdr7+CLYl2IXkk
iIBeCruJl1IyxCjvC0Rbo1Gl4/mnMGq/u1ZTNJjm3Fh2f7BedzE0KRo6hJ3cjgS8
pSkaFmeWb0bElR4SAzQPdy9jsBTPG9Il2n7jUGcYp3zt8TKigbW97Xn1SCn/Z0HE
ROMnxWLIpoj2dZ11VCSHCdDKmexDh5PCqY+TOITW813o8LqU0422Dh5lvVdli4ih
rpeE3U5kuPlZqFnPenh+4R+6J+BfzOe6+kx6febWhtm32YsRaF5AWJ16+RhYOJNq
aDL20OoigKIvXZffiljfQjQKFUVNS47sPVnavysqryVCq+Hrf70zBgVnJZyF7t3W
wL3pysm01r/Ezo69HuMFNDpMEmsd2/pfh4gBBuO1c0oeQhluofAdTlvztcz5285g
o5yZV+CoveO7vDgXBfNenp/mAtHQNSX8uhQnygsRlkyoAmqJO0Amuuc28qZNN4Rc
3l27YYmZpyviZ2cLCKaQAzCObSi+Gia2Lm+7bfqR0Xo9J9+xaxUx27vOphEnf5Xz
MznO6AzXxJInpMI50QDRw4WcmvxRgP0vFahHkL3WUFowYb3qcoktBra1uudxzGGv
9XHzsh9AzwE7a9KwG9lJxRuc9pMApu00hFj9BUtm5QOvOBUY+n3XGpzfzCObB9Wz
jWl6RF8GtW7T24AlrwOSqd3jVk5Z78fe6sVxHZEAn1NVwzz01nC8TUKsywWXkphS
8hCG1YID7QUKHcD1JV8PIPHDsdOX3S94pN6s2xkhTPXjhbejKoTXIvHxagDCZ/Ee
1d2XSbVgvAmXfBvKvwDRPCJ0bvALuKrBWGyzlTHApxVKJnJKLaRKvCho52+In3vl
HtHT2QbCBADo8UsbGMzaf6h04Bd4Kn4sOC/WUzJiPYlHB917KXtO/a0JGvDl9tw/
ee6dCWiDKlNni5zhZY9u6ruy4n8O3gEIPN5zw50X6dVvcJXXnQFQH4Sq4QD4Z+Ds
Mm9LiAmXAISrK3GdqKDxaViY8Bh1qCLWizOw+VzTjwc/im85IHIoSCgsLeJcRCBj
/KAI4dAHNW1FTukaa4anVML7Ie4SToP4Ll9NYTe1FM69g8dh5NL91dDbXGR5+AOi
9c61hyECnR1HJEKUYZ6YmQ==
`protect END_PROTECTED
