`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M09ZPpQh3SQzJxA38Mk26c/D9jMJIkrsgLoWsPMLbh1WF87daquV7DqI+UImmjpi
kIMq7DoMs4Mn8+nyHmS7Wz7PJVuEsD2s6vssnK9Dxpt8GBsnSjJOtvzHGRdswrZ7
hoBGtGtGGc4xbbKpRqQ65iGjt9CJUo+ubwScy4Igi2cpzPTNLxHS8R601FNIcxfT
Ntb/mj/4fqstFYK+upkYFzSbAC5VfegiGPyIouWVV/O+RsOQmvVBEW5gW2aANSiC
eUm7FXuswNwLw5K2weafO5g1065H9tD4J34rLBmHil75i/ldUV6deMVQ31bxtls+
sphrB023UNia0f6/gC3t4a6zf+xWY9Yr7AU/JxvoMPjD8ooaH7avyumD3Ae1TWfR
vblVitZBr+hHACF64iaNUVC0nlD9tszTCiJ2Z7J2z2AMb8IdTqU02n41vRg+R0sW
cavY+iILfeQ022o6mn0HMptBCxdqFaK/ZFCcaPuvXhq21hTB3qstOv0wVhmFzicY
9NTs0nn4n7ziCB00QYWtXh/YbxufU8AkBJt1IaXJuoBSywy1KIvdW2GCPXo2ObpG
nlJSnuRapeiTJ9Duw7nhfA==
`protect END_PROTECTED
