`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EjsJKwhUmMoskZHahXFS1CIxXhHWxzxlmdJqpAg3S5asAflNfLfy3fqBkCIrQQH4
SAENjpVmQx2JEdn6GNa+Ct5t5yWNPomc4Ew9ERpCwHl09q5wVa8T5mte/yKpMF0S
+PSB/uyfdHWjSNmM2ocINt+Ydjxe19vynr21y6eMnSxfJKo+b9N5X74bz/+EfwXH
8sicni59NVFIvHGCcRpGTLYh1b/7OXHzqA21E455foduIWQISuyCOl0QouliEAQU
uEqGOlEGV8xoCMAWpGrUqZRAH2Kw8Fy930zK/8/oA6MFQcaGqqMBzBH6ZnDlNzUG
2EF6FLzLGMtt61ikk5W9Kdy2rggRTmqpsP0acjkG7alf2U+DG188sz62bmdXndV5
NVZRTJTUp8490t4sVlSqA9ncTWiwmkA309LJHag4ND7XsOg4LsZ0CP8TzZr6u8Gc
SpYjSAXM54D234wwBE02FWyJ7VRJaPql16d7okdVJBcRs8ra50WV8RyyVoIfFsFA
zB4tLU9AHUB9fqDAFy5lBjfUmSnZXoBEPCcWlIVxZqfd5L3Y50FyjhJDqnesYatf
g74ftBahOvaAOp1BvSESNEvYmNWnPdz3GaVy1slkcdNv1GrxLqQ/RWnFaSXVaAHe
1IQrwZfJYVs+zwoXrWVVuwIyyItXbhUyTaY3nlrE8Y53tuU/f0ThWUs+33cBGm1E
pqBQIoadzIUxY8xsq4kvnb97z1o/krqOS3wnn6CKyJtxm88rBFDE+z2Y+R94v81a
Zdr+4F70zzp6dhaxIg4Ako0aqVo5uoGfoTNDI4ilaCg3hqMqdiW9ad3uUp4fp0k+
g6UhAiJqAaJDtny5mGLcE7buTJRTkwzpTMF6vCLnZcemcXrJWfpYUjnlwChFCeb1
1Gz8CR732PPtS2d0orBmXTPZ3hds7GsbEKpl/ix89Fxygt1fSj/alLQ4HBc7H4b2
Ijx9DrWRCzv8OFTNZXEpnSb1+2M47wGWtxmJnLskU9Tj5q58NHizsR2Xs6sZs2xd
89pMMBRvQ7IVWtLhrRj4gfhbWpKVNLuKKz3Pp4RcuqCoR3aewOMQvZksuWSSl/mH
ooI4yBzqiqf/j5gDdQ6Ja1sRYQrRyD2v3IUnyHXOa0DYTZhm8dF3vc8x+0ZDVS6/
rDRFFN+UVu416c2zC75Hzlu9BUpUBcduzmH7SA2aV5EpVqM3m5tggxS6OrwHUVWa
5Z8lfMqdi2i+G4ieFx81BJbCJCEoRy4MpYKnTQF7fu5I6k1KyuuwuO2UCBq/uasp
4K8+CKqRdvuOG/esJFVoVxgkJwlATGBf284L5rC2gR6ac6AX6b7JOGq//E3+4iZ3
IBqE8OgZm3mod2V7D/5EL9KPv7FM+pqT2hLEtrurd32CY0h6N8STXSGVICUMMYrX
xY+slZzTkPqNjzoKyfaNmOal8UQD2COt060+h1og+qa7yQPNE3Bcwj9blNZ1xsz5
B24b6UU8VL5MKILh5ggbwcfcNolzbm6JMRnxis3GuJ8rD78P1tJvU6IA10RqFOPd
Sm+VzqlHaVWBZUjbsODHk8KRU3qY41yFgUo7uR17Gu3Lz0b56Nq41COyipLl2pD2
V1qN9i68LwXymKGbxr2mgxnc9x9VS6dyaPjX98/S/SPE0DlPnzfQRs2xuvw5xFOQ
euOQ0LIKudmYSVSKU/U2wIDtXpHULttFuHpRKhISOyD4Z39NbciCZX8+ByVW/VZq
K5tb0k0Xh91zNC3CCVQabJ+10c4UXHsW5QWcMW2S+iwGpJ0QCZT2OMTDPR2X/8yK
qLmjfq/eV/Eb8KLf0QgXYa1k7dniPeGS9qVO3zWwTsgSppoKpqWUDYZ9w/G33azZ
ESi16MdrmyWtt5/ad49mdhC3YJAhOqxDN/zONSHV27swzePFrp1ZBtbM2C/kRzGy
/ZgZqcybKrvBINGkF5hZTA==
`protect END_PROTECTED
