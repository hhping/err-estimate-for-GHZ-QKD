`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WSxypSobjCGN4Lz4TcshJsDl1QPhCRuzeZDQ/Rjcsx+sGguxJdaSmjC/pLCybyGz
0tuIpZrpuBZUYJ8mJqnr/oqmCc3mOXZC31wAJheJ01DRCsaqjm++a8TW7emXcnx6
LjmQ7QX5ih6YGmIjmS91UnwLJSs2nGwan2C/BbuajaAxmR/h3VORcLzZtBAbExmA
T9qD2PLdc7C1tkDiD76j4f6HVNdiYkenPqNuDtBkNmpncFxDJNiLiCHQPgx0lN2/
jxslZms7NEZSxMn862RXAHnOIm8gxcVrrdKbXjNwX2++l3hO+drs2upzmZElL8NS
JXgKOf2Iv6z+Krp+zeNM+hJWwopvjk+N4rT/O1SkENrDzfKAOzNhQAL170KnI6Zx
9BPNJAuQDRsTAkJzE+0rG3txwS4HGLBxRNY5qPl9FA4YGuedeRQxIkQyTT/G7RUV
DLRpYkREY/WNsDmcEFLTMhu+jxEJeceTpLUOjCwnkroulXCeJ4Uq9sg7q+APGpsB
W4KPWQmfacqY0p9KeNs5DBVzcZBoTi+0+3Qsg00TVt4aDeXerFyBjKebVys7FJSa
WG0cAUBn3WwR8pZGX//+nPozn6h4PsjxAqTkp8Olnppy8i8Lokou69q5P5WN7uMT
YBN6U8AGVfJlmqsriL/xI88SH6QopPo5VFgFcEol3BnQhYEcxNQbyEKbJ9bFFukA
9QnkerAy/Ry2FcVxQXIaSorkneCiWYM6vSlA6Ps2SqnicoD84e6IbkqbJIFPoygV
C6i0AoWqTb2BaErU1OUeVLXnZBjc3k/nmW8PE036qN51So4WYXU3p+bkL5iv7bCX
fbzsKUH1PbPTgOcankRfvHjHPR6TPRagXxBuFMXWi7njGZvQI7iPTusGC+tKNEMS
iVnAfKr4kx651Z+zpQc2lrDahunxUhDx8VVrZ8YoW9TLjki1hSiuuHHgh8szcNTF
yPvFT6UsJ1aoFy1LFBTLYFUtsnadQuW5OZjE0eWGSas+z8KMPP6pXOg5RC5+SIxJ
zBieZkB9PoduGx1bmI1Hccsebst2DG8MWiDBTcYhNyh1crDPFD4ZarYZQJsHQCJs
TDcnSO1oUGMoVysqhU3jWLp3zAjpRaL0NnOg3Y8h9uebT/+lYU7wplghbTs2Mgev
9P2m8lwrcyBNo17Vcq2mukypEFg55CC9Y+8iDCg+RC/B7eq3BHC9tFoIj4P/An3J
YN2yFnpwDNlWpoixjcwZX2oJciRXJi5RWvpo3BS7h+Oi11ZUb567xLF634OUhU4+
pxQyBP/oi0VZd2uvF1ckKsFcqzbs/TWcnCHCEy0uJ5Ts3QoJdgSWOpHXm0/a9fUQ
calhpL/WyxwfERfBmYbZdzO0B86hFjgRy/PR3yw9Nvw2WpmAvxghbFqY0KhuR6cx
nF8nx8cnzuQCvYRlqxcVL/fDu6gUHHgeC/gs3JinhdZjKIpYZyDTuERptXwIxAaU
dODT/QeZhTbqEzO/FHB1S4y0YIaZLerSJefCwrbqFH1jiN5zAeWRTi6Ex7id1i2j
5Lm1PjzRJQ4/b7yvBbe0JIC4raAWvDYkPY/ZFDK6P25bD0n9nGVXBuSqgsZn2OL8
SOawvwgbNuLR5/AglI9YEclWj62ABT8BsPNlIbjqD6pYrW31xV+N66RjKeTxLMkI
jWWIUal1UP0D5WglX1BASGRY5I6OtHECr6rkinpJH6rqWWRgWksdETd8D1l4ikDM
S0P9RJ92lYUvmdbWlvAGTiluqlBpTKrqVYzfnFJZJ9G/IcYVTRgRRvz/2NruFLjT
gzJcXi8vdYW+6B35rR3hgSGJ5b0TOFt6bz58dBR70Z8I2jnQ9GwSPyGFDC5O7oCO
fUXiJpdEwnsB3VTCFl49bllG1cEmhdYuF5Z1/o88tyWQpor+VNXIs4s072VFhiAN
kRhceDK27iofljLcY+2jP0spxYPf514TPvrqHeBT4rfqq7QIK4qT9UuzTo5FIvN8
ng0GydK3NwBMqTUiHcvoJrcYleCa1iwrgf/NxLrR5Qfe1/428iPAPvnVqTYFpzEQ
5nvPQ3ctPd7nOaMoAFfVogMMca68IhoCRiUnEOn6guJDiVUbJnHN6PI11zTxtEd0
HRY8JXGe/V+h4GIGDH56EmtxdnOYBqB15auThc1FObBQz9wfv849YE6kvH6SWOrD
IyeBx2UlZDPWi5+Y2/kmQSN82bmhoB1UIq2wFUQwAr+sebrtp21PvaIuZvIEHqrK
k0yIloCgVxNoX7na5hP1iuMw3tTTR8dZDohXIyWkqI07ZLe/PG/GD3XGSE7AvntL
ndEPWOJyA9mhK8SLqDK1+jiWfRoallE7sMtJHTwiGyrAztx19xD0mwYz+CMK4fY3
j2YsN7WaVAhZjT+n7hMlGBUbLF26zv/rPR1DVx76ugYF4R4NFYgzl/m9CMGqKhzk
HiXKul005ZUGISLk0OPOz/ffLXxFX6MPCZKz49juCl+6Y5vWTpO0eE2S24OVElBJ
GuRlVRPIYSGpLqfjlOYpZVEWnnQ0YIlMrNPAN8fATVcciBE4tPMf/aXI4BzEmOaJ
U6HIwK18XhVbNZe3l7Sfav+USlAtxgZb/WAbWI35QITE/Ak4MLtBrtrqnnMXopXB
K4P8+w7GhEHYpkMJxpe61qlMmVhRhWgm7SeYL4WCgbO0qyg0jvatelW+VyS+N3Pm
KDae/+hJ0/HdzFXFMRWoLzT6u3LgqqfiUDWPuaC8KxxJHbN+3w4VfT/tTVasHsAA
MFZ7GdUoOhnqvv2bL/D0kqLLKir0TaXFUPcyBZ9sEZZKsBITrfZ0Y6qo8F3uXUJM
31ULc2MUYcxDxvEXV6bPHUuHQP2GrggaZs4i+IY0KILTqZZ1Ng6t4oX/D/0+2Lsx
vBCmo6/bLgo30VYTpIZSk8qrvvQHoCRWnqeLV4xBI2F7ZtLu/JA9P68NnIKiwVel
3Tz1WF5cZe3OZcTd3tUglljmwEdPSpy7GpXhIZvvtrn5wmjfIygIkZW+NcoQHFRE
4kCwQqMcKbM2LDJg9b6PAQqep4Xanc9FtypxCYHTmnyGR4A9S3rvLO0lN1ryoSzl
uYX32xNex0rVjjoklVHH/U8JBlOG7N/FGX/vnw1vSGXozJ3YEF+MPiFoLeens44v
cmP9iCxVp0U2NPjkAIXexZLCRsY/xwtnLAoBOCS8BBUNzAZOxpJZQpYewTt+tIYG
U++ADM4DGsEoFS0yiPr8FaprGByP+7MhrYZROWxB3y+uaGWqgJfL8IAo38BV1/Wl
jlSPBvdpSrMg2ePoWjHxI64w9gBNgy2XSrKhzaT7LO29er/3ZB+a/AomiazgH1jg
tGT+4byxIaA3JvJf1uXoAuK1w2zccpIshA8HIKBLhxk=
`protect END_PROTECTED
