`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9ph2ioHeu+H7/ZYNVptrMrsAtFfonsH8Tvris+2oYOpfNnm06fkynE0KJFzbCNY
MC1SewJWF7pAxEapcXZZ1YEsUmY1JCjQ7L7DKxYxVfdRQc/WPvosdJKmB+B4+ptp
liupJS5C8xenlU6Iee5KJFtlKVG2U7cvz7WooTbB0krlaLYUVyA6XR6GIMGc7DCs
oT32omhIEYa6hC7xktRCJ/KVCt6k0C8MeEOZjUrlSdA2UsJcf3theQS3NcGQ52jj
H2Y3eOtod93nmmm9zBJFGx++zRoVaaLg4RbDGUcyBqZSlDMrmmt9BJyCroUPhjtJ
Xgjrkq42XSAmk8EEJS4x2TjGpSLq/4pPwc9PO8rs/BBZ3xe2kV5+1ZtI4oUFadGO
Bw4nzsZfCIOf0zJ67ODw16lN7XIDawjVBM8b5e1azF51ycf5DB+qqW1gz4aj3iFg
ce6ybFlAB4O1u7okR6xRQsSump0weFvIKd8tAIVoguoFNG06Mfw8pfsWOS22uWqB
D4H0fcPRVl6I7PGZpfYbUo6qvCdWIz1BgBoHD+GQQmTH98ANaJeVJLzNHoKzowu/
ZIxF3IAfuYLmN0WDXYOe7CpjGRGZjslZ9odL4oXWoL/oHxSkyRUFJwfb9l1Px0jC
fExBgRQ7Ree0JmCZMZ27Hm88dv4CRPeEOqavZpYHKie7MbRPfjM3735BlluWQ7FU
ISD10E0iNcElb2RBVWIJlU9LGZuzJoEwvadzRM12MljLzStp9HwnDEN8Li02poJJ
chy3Y0S5C7eHc3py1ammO5Z9HFmpE92v8iHoGKGteHocsrFH6h+OzGpCMQitLUIK
`protect END_PROTECTED
