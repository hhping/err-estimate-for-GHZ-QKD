`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZKTbI/3bjtFRIa2Tmu7UgTUn10EcNFer2p7nNer3DIVEjU+NeLMmFXQ2Rhqweu/
duP/F9NsLyV9YCoWJWyxpOQzIdUNjKYwNw6mWQl9D9Ia7sc3OaW6Pp9e9VKTrUJ9
L/6+AwVioW31imj1VN21+KZ+HHJooS1Z7hB03bQ0avRc3MHwnZy9/yOyABD6NZSE
S6Fl0uDr0+lJPJdLP7tEJbwwr6jV+yzjsSE9pwE6avhFebJZSkLtoGcfMf5QxdK4
F8asIReL4PJeS/lNl7pSglB6j1dcvLnFvkrxbshz788PHv6qGuxgLGomjc4ddI6z
P9XLzs7rftwyKKR7VON1MDauNXB8JS5tnKlCnt7TIDmWXfNaPFnxLlAi38Dtw0+S
HvMTFMcPx4w+ieIMn38WTmn/AP4l/qfTlYa7EffG22opAYPZqLm25Gs8l1yVERv/
+u90E63ZvK4dthMWELl20/O4SOMYPo/GdvUrWkQ/l4VT9VNOYYgRU+qmUjHo69Rt
Vq9jTPCjOvPuOqj4YhYkpyQaeHrOXwtuHykUyqfn39UKyI0CXuULE7JqbGNvxyB4
7AWLAI5Hods9BeldIvAZduJZCKWqCuSAb3YevgkOaIf0gNffHQ5FIy0YQL4L5oBz
7/Y7h6vD1CZDLg4+uagX6rSstZp7mef5RFd/5mLWEOuTodVcQFKyA4heT9fMl6iL
buYOWwzVrtZNGcLKe2afV4O0HjMmjs/+g1AkqJhefoQuTzt7XdglWg+eOVPULBKN
O5ESRZE57lVw4L5+ueXo29MSDmzz3zbAbEXZDw1n3GEJfiIJy3Y44/3/vxxQfwip
brrvz52DhJKWOEl+jXk/2s2ZWa6RsjbPYwyUWp00+1FtsIqRp32ZrwMAN3OVTMyS
zWUkFiWnK+JoNtsnJlw5BL6KfkmXqkdIGA9zuHYWj9JxNiz5e/5zAbytDrL5VOhm
JtX39blZmtTQLcNhFGB2B0nw7DaBWeHIpwGvJJqPgyMR7+9smffbDprqSeqI6tfm
IfCf7NUMO3A0CU9osIF+ByZji65CQa9IfS3xEhG+dmpRbtbEbuVtBR/wwwq5Ojne
rYFUpVOrKtFTfO4O5PSV8xM2HFhalE/F/+MGfVCM/NAD1he2Vwsizy9Idgk2BVV0
F9tdnSZ699V4n7mSB6C08JRsUtK1VfSQCDkp6Kvt7u5LpWYPO/ZbnqucJGeJJR2U
aK9Ilx0EsIvvI4f0POB/DFUPbflg+JYhPFoBuA2i+e0ckNbqV1LrCGFUDHhEq/5T
GqA7wHw8j7R1v9VCjJwK/pAd6PDYrYAqDFX2hOIFEuICEf4MPV8clLySUkrJGmm6
jwF4fU9z8EKDbryYkXAA+Jvp/vGZRgw6BhXLRyr2VFt+KbfVmxloTZRm9Sj7syZA
JSdkFDiMzm8+6+2AsIaOFlGCcZuNk00U1ULatWOlb0RsLOy2zt1rZ0gJaB/L3GUl
0X3N0sjItgCzAfF/GRQlEWRK4MLvb0VNqyrMRWtW3L4YPa6ISbzy7OtGtRWg1Xqj
xw1V1vdWXnDWJ+KjtjWZVUVQAQejrVCaQi60S9yjGAmSdP1OZT8qf0W8Ji3tLCa9
hXf9/YLuA6JVLnRZk3KkjJjVpP+tAz0HjZQYeh589zl7VLY84vjTbBbVzoiPMzCg
d6NH9VON/AlhHhVk64fbhZz4WLwhg2jLc2KoyhUB1qcGqk0MIM9NgRoMOgMBuHOh
BLIwYUWd/TXO3iJTaz7PIAoayriwiyLziGv+ecq69OGwKbobTHyrQX0d51RyW6HO
do66fQGzavixpaxxi8CRwVtcG2YeZXFEXYculwspt09YBRwtSZPWxXf/QHoKIpBi
0F0csLdeOZI1aNQ6AuxS3Q==
`protect END_PROTECTED
