`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oe1R43WaT9YhUppir1+PqtuNcmisEKDEaYRfwH5HaR/STnxN/xW6fJkCdXI5CPUz
ocBm9Ssw+zIpSFs7pvugXnBQvEcQsSCX5rUfvnbJzV5GZEYbXnwVayHLfS8Em7S1
ttECzpoUj2aNrHyHCVbT3wnTwbdnsA3n6iSczmQta1xfivUmcuhWMU++59sCKo/t
7Ap3wJibxuODreTRduBWy8KlfiuSUqwWXRWRkZW8k6/+d8vbnZ1Ljq6XK9myNJ6I
yCN1RzyFPtJN43oqaH2o51nfaOn6EdG4ZLoa4wf9Kf/dpHZRR0rPnbVl+GiHCYtL
PG7YQsLfT5GJ0EaYCIZeBzasRiOD+X7q1bCq2SzvS8peaGQf5FHqJ2Rfb3nQQO+T
Za0BvX0fKTW5CeLIW5BPlit8ZWvvFP08/y6jZBB7Mi9Sx9ie2jHdo05yTMID9e5A
KCGVBMTgJa3dHHhu4bymS5GmEwADMklgvYFIUTxgGLo82/kbIcIYnWmSi5+E/N9s
nztssxTRElEAuSX3iEQ3CHNIDQ0+aqMQznv08d9oxei7V2KUIfwPoTLnjnG6kvAX
oxx/rYPmpxit+RecB6R2y4avhvsIogtLN6DJZBjk1a9AghUF0YTfi0qgCr+bAd2X
+1NDXSCXy0OHXxA8mfRiUecxHASYcCLMUC6MLmIXmbN+3AT/M64RFblwwnB1O7ki
fSY/VjKCC4LFIhahaMXygCHRs3AGIWirQch3xjcewS6XEEvhv1FXFktWDTPPO5k0
idL1Qmp9evOKwhAZMNqMqS3oAe9JCUPBXdO+23CobQIN4fkFdav56Jls6KpfE93u
c0SaFt+nxm82Ninpx0j9adEumMjby9TFiXCJcWIgn3O8lO9AwuWL5BaB8W2ZQ4//
k3/13zp5TMk3TNbP0JGgPIKB4MQEvgh3X5VByG04OYCTrLfvQwl68hN/BKBqj6ZL
Qv9WAS/+gz+ay7gGQxlIx/Q4ls2hD4Fp5RS8ceJIK1E=
`protect END_PROTECTED
