`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ytg0S/oRfNmporRYlLPBxj+dVv1hmGNrgr/hEEca30Jx/uuv3zGva6U7liyJ33vV
A8UYkTnOtNKdn6eXJnU8PgnT2U3nsgUeDlRsNXMe7Yud+K+ZH87deBFTSbL9/IH9
66lRj4FwOsmlxs1y3pH2kuP1SkVAgrpVK7cww70eOafJHXlhUUzxzE9wMHDj6poc
4U21xMc33Ik0QNeWah8x4Ghqobe20W6zigdM9JFZru71zoCOIlR1dcejIh2fFXFh
XJT5oM+u8TgIv4mFp1iaor4sVdAzqReIFE+gNaTAh3KJBRZFtI0MlpbV0m4lAaeR
T0BH40CzJqaLKseAJBZhb2OGOtI0s+UJOZ/XDcmEjUdq1bxOv8kMgiPXAIi5bI9N
huwmKPlTSqDZmUQ18aRiwPVAxI+7spueA1JQbWT8fvJE2PVTxB42nPuUSPpA8fYo
fzrLKBLXhBdJSfi26Vm9OE0+6Zq7Ao1bSvvMW99Rsxz0Z+evx49m3VpHvEPrgC4l
OJZfDABn6LzSx9Iv52wiTn1H69KYHVRGw+JLbboa9ciavc8OLdw6KLyy4m4G+zu/
Ul74QAxke56aMA6zcUiK5MwKyZB8Fe3DO7gLtuKChFNBl8SC///nSkGz57oUW7yZ
gjuDaJUQpk/xbPnshOBa/yU7bta4t0yXxsX1aOkGlZPec4pjlwqovjJSYwF3fsiO
/LG8RyVKBTjndDOo3VHD1N0dJgQuUpUKBKeewGbZAY82W4dYadG9tyaiEo19x5zq
`protect END_PROTECTED
