`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UUz5b428hpRa5w2EAlwo8+AbrmZnUlfYw05UvKx8NTwZJRgjpVwiYEVDbeIF3uZP
ThEbfvltgxp9G1zjZ2YDQ2AAjb1M8db072L2LPodgD79LejFVNKgTnbwmGflgBhP
9lwllPQUAnOGYtdhAaQ1YVkqdqwuR0DLJRZC1ZvMpdCp1u20YyW+cukAb8pj6V1i
qb4CZvVKn+a1HfxJnezs3/ypJPLgh/U0lerMjAZ8no//lH13PK6aub8cM3AdRAej
MJ9p2aCfzzrdAaJa01jepLH0dSOuprDETFtOVI+zoGzD0I9xYQWbUnCIz+Iqv0YN
yayEjs7L5hPxTDiUiiu0fw8h+DNIk14DPB5+wh4s9UtklYhJjDmc/65ynia2/O5q
QTD9L22fIeHGUYn0fHZaD4UUf6RQqw30OdYqwjMGSElI5o6l81RwdkSidhCUxszf
PVB4gZZ4jE5sBMpnNsGkiiN73dbIHJ5r1iWsbX2ewDJeywtq80sArQ4cGKnoQdpg
z/yF2JkKukdIyvuUpInHkb4jGtKtLoKIRlVIJTbJ6Z/HUZaHvQOj47DR7WEbasc5
SNU8Wbsfn4v4UNg/mVuCalDgXzjUNZtKAGD0tBaR+HiIuZ0SEgyKFLeGm7x9McfA
`protect END_PROTECTED
