`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7X3k7osQYbORV58fvS/qG1peGreHazUXA8fpJl4Y4ek96Kn1cL6ccFW0CZHMzsO
6P4sa0N9WWqepGqK+ugienkp4Ku7q2ghL+shVHdcENhFAsFZAIBEmI+WTrjGprvn
OtDu0YkMspjE3XBRZNAN7o/9MMcQTkekUxYZkS6zrBe+E8XOqBB6E6vGlGJJPBUO
kWEDmsyci/evN2YC3aH/x9UYkfaxVlVGpYYDKaLrfL6MXp7oYEhgqdnvhvjV9Ip+
JJQmhBeue16aNuNwKaqMeORKt8+nczn29YJN0uqDdAzBaApnowuNSmcH91N9LZrU
nk5W8rTFWvUABe4KwMxuLh+7KxpyXeLpKiOKZt7EOKh8uUSYTYy3q4ZnaPT/Vv4k
JRQmqmj3RGf0Ft3Rh81xHGhKii/km7MmeNQHjezEGCXIQ+7YRtefefN3Rs7Euxx7
ygSGkf81qEJZKVY4WGosiwEzfXkqFupjDXpJGScgfmP1gwojpnvMz/yBdUTMogzQ
nrixJvGz3A8EOAW6MjT24taYLsOlXIs1KjLq8e7XpPf6lgPvZuyRlgVzgtPWUfSi
LClo9+0QpX+m2rv04BBYoO5QlKioYMZ7tXwOq4+2q3o2tRBiQsQgj2chKogq6kYx
jacakXKgd0Mv3U7E/ir1T5DdGHN4f/EjaNusI6kK6xMWjy/tu6TFh4R4dZ8KsZqd
QFVph2LyL5NTghD0P6biUeHKCqpwmX3sVp892uORF2SEDFuOQRInXDe1ZVxthZ6v
eKGX1Nxx4MoVIGcZmy8UXsbEFt+U8RQwKaQ/6DfFmGosgb/qdLwj31jV07rQ+Jhe
3Xd8krjHXzKuHLxLjaJTn8R58BMRIJb+RLgUk2kOaWPV0W38sd8bGyEBI1L6RJzl
IpGWsME6D05NDCYu4mqsHo+pSWB867+WaJC0BqRsuQJnIs6sru2HYe65S7b+4jdY
SztyQpfTqeLZpBMszYGkJAaZjXPSQ5uGeN4d6Iyglfgd05x1Hu9uzMqu14BnjGYy
wEpJ0dz40NEQFFeWo+Z6UlSQHygYlkuC0QRhunDiLr3bInwabUTMnmQfH9kibNwk
FEZI1PF7uvkaAvo1d1YcHODzHrhSgDDlS62hyQ0+UfnvrcpnQuw1r3EZglCIydI4
3jUDnp8pmS6Tr8XPRRm7d3IciKbcrhSYsZi+Rcj0f8y2TFMSbx9aljR5k57KiBnE
Biwaf38kElGv+rf2s1lYdIqq1/qrn/fz4eKMpvb4L8NzTzGI1hcA/QrE+ys38u+1
+WSdpzTM7hlfL2BzZHtIHmg00ssEEC1jA/glpEyuDs4UQrytKUzBefkI1cUqtQkv
AE7dOfY13EMKKcn6cPJCkeGTQzHbX0tV2DYdtZNi/JIcgsvX+vCroqCZi9Vb6DmU
7WloeaYczZgbaCmu8676HPYrBhBQuu1uuw1QL561zp9BCVAX0fZ1Hh2ZV3lqlFGH
RG9r7Bm3qxKH5oCTro1PJj2NBjA/10O7PrLQYMY1lVg7U0yks9XOy8qFXmYJCD/Y
9dA/yYGguBW0+Ohf0U8FUiNyawT8NjoSbz1UckAZX55ONpaL6R5Xj2NCp+06GJJh
/qA2ytz1034T4fYtbGTiVNKMhFuoSwmuzvINBpFBint4rjgSFqgVgGwd0wz1UIOy
NOmLxIstBb2KXdIWSWxmsi2xNbQMMy/EVtkoDIkbuLn1B0q9VjRQKQUlntI5yJbe
iIrAi+zFGyqJREP3K4A3VWpVNpgbIGc95waKfmASC+sKyQU6qS1faoVwnj+mdB1F
qvlmuuNv20R6D1gshpdMHUj14JhyWLBI7zYOsmWrnodP645lv1cj5N+zGXPtkB/b
M9VBKu7tC0hm5K18+cBPGHERSf5jWPpur+HHoZxt8xyz4mPMkAuhVHYQQN9tAMXq
2pQHHJeNsft+TgyhqL6rhjQJmftRVd0FPcFlV90QCeUoCRANbKdW/NfDKOMQTbzP
rhKWNb8K0ArQZg8Yg9MyLpmoWqr+jJCcjxehCd6siAfqyGIQFHrv8aKubl/efGmc
goZulJ6hMZadHJKQ6CGcnJRh4yOC0zlmTKwTWVknQHc53iHp2av2O3s4Aw6/dHmw
GN2q6QvM36ZTcrFRlYB7hOsXjvohZVXiWmk6hO1xX+sCDyD3+SEdDI5beE4QimEr
uP+wyF8OYDdQ9sZAYtUHZiMBcabs0m50jJC0T/xgiX9V6Evp4KpQPHV2LZ+78brU
9LFBcH/ZFanz+N15Xs6AwBY0bSc4w+aueTXmcipeTFTiF6RSl8InTThsRKglYLaE
3FuG93WNMu9cvllyBgwTJcGr4gn8XeNav75EqAfG+Xx9DY9YRuq6/tSN8z1nHiJ9
g0OAgQyUhPkVRvQtqZ5w9akgRlNa6FB7iQIeyQOKMUtwSBm3K+4nZ+nvRyYFtZNT
CGTj6bevoXVuiFIxYNVm635f7WWbdJGqdV6A+nyuOTxxDAf8FlJ3M9XuWFGfEF72
vZZGNFWrl8uHIYJLH4VzxA==
`protect END_PROTECTED
