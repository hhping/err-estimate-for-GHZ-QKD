`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfrrzNgsMVjTa8y2pA9b4PAkhegZJiCRLWH73/meZrGxMCo0rhCXp/Zxd8XKkxIN
ZaIZaYrwqWhTMDBUc77/x7AXc1k55yVDR+yZtOnKw6hKDV3FPpL55nb6HUITzRGH
ErpeSAhM5G322WCfGvHlKDeWibKIlPNeTMbbEIshkwsbCqRvJPoU4TiZams/L0z8
tJAF8aYsp+02UUuBKmxd1QyzuohIJpSr2G+X5qnZzfFeT0OoLlqPqWRDky7bEqPm
U0XtkPh4yKCW7wX96bppmMu6c5Ki5uHpvZJN32m8b5s6QsngWcOg2C9QHQqNIQ+P
/8saukQo12jPK+N4AZ7TssaMEgM4rUMf0Q4Y5fOimM/0udUAVfL6WpsijrmVg55u
m13fc7f42CQW4s1k0bYhRTPR1oW3rcWMA8FvS+e5OvP9sLOwHqVvjtiqdbQWXCVu
CTIt6nDAZwHe/9F5gFkG2c3RK8z5uUdYmbHfeJjgHN6xiRhTFCostto8XIWEioO4
vmajcn/EiOYPCKSeGYT3EjXNImcQPtBaHuL9YY0XKUm2t8O6KqgL7nYoZRNk/3i8
WXDurt5+x3CMTnClBCmgZOXzWD70rJEjL6h85JnqF5ZRIvRSSCgElN/n6Ekcq6CW
+B6dhTM/X1NLLVhC3BPtK/6ZplNw+GYNkeMLHuIgBa5/4TiQ76NoFCbyc8v7Nv+x
J/IMD3ZKum/sagD7AhVdWHFMXPQUDROQRg5sJABGuGjLTWbiTbtSJxJbzzxdYHOv
qjORwzZe/Jzq6y44Ll2nl2EvrEribymoEMJOUWfzCR8/KTl5AImGcwGICCWl8DAB
DfK+2brKNmwl/0QCJxijFZdT1HRAT9VHkiA5C7C2P0ZvioAYRVKrnfIeFdX2ucVT
KCkkrdHjlAkzlWgDDbD8lwIwjSLmYYzFV5RcKPagfJs9K3yF1m1e2b/m0Y5YRLBS
TIPMeAFni8Yy1mNQbaC+ZxndqB4QBsFkzHtwGhBML/6FuzvY+pbA5ocNuobmUeUE
G26zAEcWFv4KYA0GoqpBJ0s2uBBS5MnYjc8O1nXWhXDueZ8/Ei1I+yiEPdriSUTq
/e0Gx5DoG9i3iWsaFZ8JVb6sCydCt+7AD04E3Wv4uX+C/uYbAUYo8Dx3mxM8QGvP
3AXP9xKykHI8K7MvlaVw67kwmcmqstZZXTP/GDzPr4xuYCHbIrChnJ8TQ5HrJ7bK
q6jdIn4ZuDEBpg/fud+mps4P8jlAyxxpx7A5CDoRTr1KhOFtkU4h8Mp4MqljfvRD
75RGcs3OeyZIiOqWOvjiB4D6oGVF9Fp0fv45CG1ItzrYMZ/Wm/R4kbaxBGyZpDj3
+3GbvDrWprjYqJB0xKLAPhg7Jv/HUaM5RDbGR+rzguZgif9NSyOWjiKzJPtqNtTI
NlBgGuDHWK1OVby7vcxZaxLpQgkyxepELCAqrHdCX6XjcQPd1EisPKvlISPfdndH
Pf0fjUetQ/gcJH82JA1Nxfmwqha6U8jcQ5PcZPLWzq04NHa/u+A62j6PU9yfHmuy
COJcXbje3HVgrV8hDJQ44FCaEJ7C1qgaQssKRMALpGM948LpS0xdYkM+2WGNsDKg
+sgL/UrBxDhDCx/sKCnpEdHQpVURrMpqegTMEKeFs5vFgGYvIv8SZC4rInh/CqmD
0DFBSGavYjdd6lVwpanJuqAU6QKVGdY6tTeWzb4Lu5zG3H+1FspP7BFIt2XYCgc3
yWKut8t0/HBegCfDFHyJnqTM58B9e+ZTUP/a7zyWTv3CeNQnGE2+jkjtGvfdXNls
agpa/AEzKj82IqGuaC49BwNjNQWHaNjxJlyG0ghKTnWMbvX2A4hAji4prWJa40+9
Skzflf0uz9xPnpxkR3JetXd6QC23GVC4YSEwYpI0HbQ6m68ud4bq6eOTWfqnGRml
Cbkn4+Yhk8oFCC+ls8yJA7fTlhD+qjWqQ5iSepz71tS+kblYvYAEHPfzq0VcQmJC
jVKywz1+fKbelDEEtRZLaQw9ei1ubNW8eJD8qi6TxgKuahPBDXMyhZHP0YpGA323
85U21NML5vaj4CfQaa1qWJsHPRBC6YhK675qZn0mK8Lsnoh1Dc9h8Q7gpp/qtMeS
Hr9BVajTbZS0egeSM6E6ccPZEyBDUd4Z/b4x6vXgHgXZs9VXeh3HIFRbPGTZ87u4
Ps3WuNb/6nIoM7IWiijJDuE6z9c7NWDtkyzctBTd5pnpNDSm85RZhfd/YHCsCQd6
6EKwM03/vfBm3HZI9otGb0r9P0T5jV75CFY7FKygOP1ww0n1e/iig8UrftR7bOmZ
cYebk1CjYOg+ArG05Q/nK3fqPmo4ud7oYV53+O6VKyBsclZlCB7a6Rgvfb9/B4FP
ZgiHxzxEhz2VboAu/O3Hk3iTmyQMpxrqWJhMAjmyJgPqZl0xA5tt3tQ0ZK+egvxh
W+lQozIbDpyVnHbUFkX0TB8cQKqI0RCiuYIQYejCDtVlIEBjP5QtkCA/PAifuHM0
FcR//KBXQ2YJsAiQM5Hlc2Pff9hsdMd+VnrpoqamQt8RBCB1ce1O5O6IMYKn5x43
w49eyW7KVFTbVDQoSboN2TgLZLaN1uAny5DWdLQrjchZ/5yc6Nk+fR/eO7IvGx9+
S8FjNM8i67202Q3EJtl0j/lLLvtkoyXar5W89AQukSoC40Vj8jEMHLPVEuKtuy1G
fgfZcIkbFrU8FhQvcYe4Tg5SVvu6VP05XP0cxo/YLIBnUNBm2TCyPr9p+uLPhr01
JZ0DzQP/zFr6NFnt9i0LJvpGA+LEeiu69GzTuKwG+J+0IJHXKa5xXoizvGemVr6T
AmKdoIhhHg7YQkLHOgZxL9QjBegUELkFzW/NPkBNHjt3+tZebry290cXIpEfj9j2
`protect END_PROTECTED
