`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
37A6XnpwYNl1DlgONqzB6Yipot54Ry1Il01lPqK/XEmPryCzwOSx3mNaYSMJ/JLG
N/UYCAk2OQmKji7F3mGP60UQbVQjy9d2P0LBlBlJbdiVMm1f6tNzvj9GlYDIOhjV
ZJ8G/BCxol+t3dDkyY29hpP5B+PxUTirtOT8PhEceRjgp8aiCUw7u7S6jGcwsyuz
ZZsJyQFAw1hys42HPNK7prW7bwpX0uYSw3CjZKAFJdwjGhqCjb4cWM4mx7IgfwyZ
cg5QfFse7QWlUBlpA66JwvNX7QxX2Y41kVpFwYGqD8ygO3aYEXBSZJw+Hu1lMxoj
LECfg1hU2e/+9CdsmSuVn7aTNzO3t3AJgCRftXSd4HTdZGKpI6G4qahQzJ6NAmwC
beY9F3DD4TkuvpGmYSUpOeQtJ3riGorQuKvCO2JGC7SJqlPB2pPCNyD/lr4NnGYn
6q25uNIb/NluQejSCe0/jvmD/Ug7mIM6Lfia3iV5+0jafLpoURj3rU5+OsCoMex3
tEgcCw4/f5FkBnpFVgtXL6OilpZR6itZKVebj4qrVNSxVHGfq8Y331k8Kpu4XfpS
cUc/DfWYJzLar5aqaeCulPr14MGHuE2Udl0fse0Za8UUzTtXuU14EqgF0YdqnRcM
kaV7AYKEGWj+jEUiaW0pkEsD29gq/PoDu7ow632Vfgw9UxT/q7yv5IvwQQ7VAe4L
Jhozoy0EqC2nPd3JkObsaPbvrX5Trzs9HdNatXHeY4sk0fKDO41Mdh5fq+iYeceL
xJ/lFXpMlaySR9at9cWhcVXf7oVAMiAyJTXZ/k4U91+lWZX/KYg8duuIVMT6ajT+
ErMiiXtnsLTlVRsCuH1Mp8VeQUuwHlo/x79EbFd8ugB4nEMz1XQzfmrumzZVjEwe
dz6acs/xkQGXPvouKc5dU+v1FjQqO/V/sY5ngF/YxGu6EfOw6XXTfSMU1cOXCRM9
A886xy/ybSsiXcbrK055e6uxJQ7jldCys1CbwGGw3TupwTs/ZwXt2GPkB2OJwcBh
wUG1F2Gw/5TQrXnTAfXv/xjthuFVGA7umZkCGihIyakjwW/oweBthLxqBQQSYoUi
mYI3JBWpDu2sVURo4tPnl1Zv7Yr66pIT5lV6cpAnUHr2ahspk/A5X80Ar2j/ry59
3lA3GZFwFdL+xcg1aE4smK/ipxMil2kxbnbxt9dF2PeDhL/En/3QnlQcZlfes/TE
XmIRI0fKBsepI8G92DzbHgJDZKENs3jjc/PDY21X6EiLYJAdgkv86b1kczLHvazU
yfEmIhNqB6QpOUeGssB4SF6M/zIgZPPEPee8w04G5DAc/PCV9S9/NTSQU1NVZTPX
6fTf53zEGGt5oVynucgnKldlLRVxbN/ciVdRoGIggIW5Eo5sAPqBtK17pf1GCgTJ
T+d/HkhILouXsq4p+UhJX1UX3Jx7AAUDKug9OyaPLORssxB8F9BGG/6Oq6NYN+b8
OGuRK4EoRkNxaKTR4r/eGtvjL5RLtBezt50XAgosxyQww78GY+ZNd9NATbKgd5MX
Eov0EvMZf+l8ZU7LHJhNOlVzwiSs5aCvohtKlUeoEYy9zOld+VbHeyknKi6NcCei
pL99YGn7QBd1ymjPn7zCsuEPJqkLxl/9DQKRrB1nfktiHowUaoZu+/dO3dpJoAd+
CBrX49fv500Eb5cRCySUjK+TaIz8t8OEDRBnz3jYHIx55YMaTcL9H1DiydUh2d0Q
zrymFJacWRxVyYJ4Uy2GHw7Ia0yRkWzO4SAp9Ly6d+PLxBWGNWS58NRVGNItuRiE
RG2X67h5K4Uu3RtK0eoku0tqL7eVvc44oaxI79p26Rp9S/OT6jiodChkVxx0iGiN
NtLet/2mqwlxgL103FWRrq77G7Y9a9D9ukzioTUCWxXDuj+dlzPv4Nnun9f4ZmdC
4DxKBoBQbaHDNlyp01V06UH02r+C50F/eV5mMFuEiXh0IHHei+mR99FHbPh9DSuh
dmEX9g5MX55bZoR75RnBryejoCxsUVcfWFy6sWQFcnOCXJz+l0E3PBuHF5ZFgenF
+540rCRGxtVCffSJEs+OSlVG+9/SOWXjD7YZzBwEKf63NJgmo+d9S0qkYRY/BmUX
rmtbkN4WHP1NRTzDVNUXXnVcYiUUnQcql9Rpm2p6aWYz8ku3cEz98057tHa2R3/z
C24HcAxnqjdrWvSxYSCMw/zUiyeIq5M0DCzg0XvlMhRwGnGQgsXULHvoKrEWhE2V
8YOXWQJQU6SLPr+a9nnAId8uN7OkD3syCJ6QQF/F87vs7Ix39d/l2kFYofvYr5n3
GQfOFdxEcAWQjUG4ugP5DIV+tNnC3Y91LWc9JFhjyA7dwUADAnfKoV6aQMVY0V29
2kD/coX8N4o5v77VtrVQFOrTEcLZUI+NZnPzZYdkcEC/i2B18Z7VFVqXTcTyybzv
HeQbrXe7du0N3SN0ZWlf134UJ64ktYNAGYPPnSGOSkRd+2QnskjQf68fMYmO78CB
Xmc5d9OVY3rtEIWkWsens6TBR3LIpZpsa4eo28fJtZToJgc1B3IRhxuCcQTL1Hkr
B/uySdt1ta7XgS0cjt+XkUM3BHlw8l+BoBTCxr4jYJIBm/trDKa8cUbkLUP6+IGv
pys1YmZfgc/v2dwJ5fhvG3ZvJ4ezW/zEY6ZdaRS5E7mq5Y/blc4WKsS+9CJbdTYy
qy2fEUDIHwOwyMGx0Hs6cMOkoqu0yZxnSpRglEnVbqINTyI4D/nkFqEFEypZB6tu
nqltY4eTB7HetFI+tzFoEgnmlweto+I6MIYr2evjHKOD+S6/sptfzTMWa7zBk7nT
RGu/QUowIR1AF3UWJRjN43KYyfrEef9ad7qLHSuqxzT11n39jrXQBXupsWx/CLUd
VcF1wsr7Y7yRg8Yso3QD6+ttSVcu9ERR1CRR9XKD16SNoeeT5jsAL1s71MiEUGMw
V+f51yUj5JPi/hH+b6P3QH7J1+WTMNkzOM9ua2lrToNGXJGClav1BteIGYjuPeCs
Dp8lZY3up0FKMP09cepKdL4gxeWcLq3mw5JTgQj7LLY5DFUZAXjbLwj+a2VjrfOr
LcdQD8w6ymaX95b0aLGJP3UGr0Uy09EnU9O6e4jtpvW+MmawwGN8VG2F4JQ2tggZ
XFtYWW3Zldsnxnid1rSSs4PvNHPPuAJXrN2TPxQOD5jAJbOAl0LV2OGo1XQnp4WV
/Bs1JX9GoNkbqoENTOsfAA==
`protect END_PROTECTED
