`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7XS60RpWKpAPWSv262z+Rr1i0jCXUgKD0PV5eKHYYWWLZWoQNEdzmIywDj7JXWq5
1D8USKMsacOq2W/iINbCCygxganSGbl//IucNpY1ulNlJjBF9pdkezC6+jFwm0dE
ad06qrXuh6KBcS87ERW+SW9OWGkj+k+iB0OAgbEaAxYysZyRiPyT/QaBC7UBGKhp
T8unHFYOD4CNFbrenmEW4SzU8Ij7deqeBVbYTwgR1UaRN1BStVNL5Ff6SpqUjwnQ
LDleLefdjOXNqLwAD5SS0h98y7Wkrvew9xR6flsTMj8n9BTx8hLVsPFw1nLpKGWU
DYXpDFZsSUPevM4y+B0V5tcQ3nGinXq91KQGEjED2guSdUkhC6EUXYxhS2kzmnT2
n0cJKOFyZpdG60FSp8OjstleKwgwLRENzh9sNxjj8xigirwQwupbZjO2onCl4N2+
x3O0DLJNFi7WV94VNUxxlaTuFUy96d+umiQoGnPC0i4pcHHczr84M6r6IcFC93aT
GOfZiDNU9XVKJCtSfEHTWJopsr66yWsz7fTm5QI7abLJhnFK0cQUBQi7eZxlS0zY
LypMLrbSZl13xMCqfWABYVJK1cE3lwYF9+KEpUhb93La2uJx068bmcVZi6DXfnNC
F/yhLSNdLgFn4j4k37OLX1+M6PL8+HlRRcDwxhMr6SLvKUQrUDoPuWZIeBzZkSk6
WbbNAdbGcp58G1+8CktnGZJGpMxvVQjo3vjzGDrcJZD8PtzSxW6UCyR/hhCKrkfJ
eCq/SdZDdyTBVXiUyxqh5glNCapbNHh9HKOy1XGGyFLDEQK2NtMrJSjcOJ4bneS0
s3PBiFRHeF5ukbOzpyaYGXqOEKkU5jKFRzwcr4sZI5hI/QzSIb1nOowfseFb559i
LwW+5hYBkM+CDQ8/0V+cVqYdb5wosmMnCCQWcsntotktrvroo3Q6w/0wZubZOhML
1rVcjGrEh5eBsmDJLcKcy2jgJ3K43y84XJdhAkuTo23UMKUlt0HnRtG683So5b1o
8Y04KBmgEB3cMz66vweVDJgaCP1wUH1sATRdt3Tm3W6UyPbThToHuirCqbYsMlCS
Wo+Z/wrLfsDX9x5MfeayCgu4+O7CU9YrAASWx4Ud905Yntm3WxJZ8TWzk6lTSaMO
P04biVV7MuPDI2JBQ14Ju3Tfw038Fucj/11xGcPZvK1ZfSiT4zbGM5dHAsanyk67
0mq0DEqTTO5I/hB0cUWM4lJms+0uwihD3PzLbxOTy4BTMgUUVEW9pOWGI+Oxadib
`protect END_PROTECTED
