`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPIt5rgipz2WLZ0XrLij+ifCRygI1o8C5o2C27Cv4OhAjwN+lI6FnRiME6Qn0Az/
BePWxyLd38dGowD6HcYsE4/HEVfQnxHqbD7m4W3ZTy52KRz48fxcARamkTIzYLh2
lVdbEZgBudFRpCb+fKgvi7lgVLRdajxodRuNzpFkVeXFgE9zgeHohfUCxxxb6mmP
7FessnR5w2d2vOO5gyZkMSR/JjY9GCGvj+HyyIGzQYPB9n8aLmG3fWDWOrk6EFf6
e28JlZY4UWCWu2tOJMYOF0uzwT/ttOo2Hkb0JTy4DYv4dSdCNbF7hUErHC0lyjsr
5oL69qzDuLTu3Agmwmmko3sR/Ja/esPUqMu/WxABB1zJVmxKM7tILLbjjTaNZJ49
WF6yUBfKS9seCEWWGDpW546UxH1ic0fGoICd7oN3UmrFEeZpuJSF3vwi/4RlLvoS
BU33iv14hHij4z/yHHV3KTAKX3SCwLwAYpbOGv9lnlxkiMdZnIIBOfcePZ/Kpsvh
0tW7D+Pb8airjaLy6hGm90tghPrQbICxwDeJlUF5cWLegvy4KrhNxvaRa5IIQiM5
r5i1L3galY5f6X88PRgL+EYn7/wmA+L908jf2wqufuCZSM49f6COEj48c9s3KXrh
DUY9LA9C0Px3ePDicSiCaQ==
`protect END_PROTECTED
