`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nYcn8pbNxrBQb1SsnKyHnA3Q+ASwfqjJDOVr7oTX6fCipVvOitruM8rSRlQwZjVM
IUyU0krpPUJYlb3YIy4LDu3VBynAd/k/4i44jbGhBssQ8TWQXO5DHbDt0fYVI962
NiuRaUx63zM1KKwJ+qSrnyHr2ypU2EZ/g3M6vmDfB3IxM4djLoS3OBTAAD3A0H/f
qGNtoCEN0aU48rKL7Fuiu10jNsh29yAvtkMOy/H8adhBUyNHn2N63OZbhlErxa0F
AZP9W9GelE+HzC40TfTQ5Dk30Prgjp9ggzwDn958ILxKZL2DQWZJvCwHQmqX5vBI
NEVAjcNt9l1CVGQHxA3NPe7GSRXsI90hhAFbz9prjkaAhozpJDoy9FSD/ePgXvEY
Adh+8hUUPB7JP/fWMxK/Y2rlIzPYrZ1aEDkruHq0FWq7oADKHCXdWbR80xspBdna
xGb+7i19d9V0tF9qDXE+3Iy2MjlVBLRsH3ceAJ6ptXCzLlVm3oABpOrfgrxalnod
xB1mpemMOvMA6fnxb+c+ZVokRTADaqZ5oVRScNjcTTzDASqJVZwAHF3871Oi3fCQ
ZjPNsuqZhz4dyOBv21Mb/ed6Y1yyeynwJ9jJm3pC++u5uQsmAhJP2LTuDxB1ll8q
fVycyr1/L5SOITmePc1K0UwP0gjcOtTBnxOYEFKMWb2INe5CBK55AyirZ6NR2fdu
b0DMf4mETY40Gc5GomBdXjBlhcwWD5KVrot/Gk8nnib8U36fCqYYKfW5Q8bXikc8
BH1uTrlxTY75F9mz1/jsh0LDriDbtWajr6vazoEqk3PqAn/auquIjPiyxElL/jyR
4MfalqWF/MTAJjtn6omPFb9zZREdG0zs0TlOjmjwAhFAPmi/3S0RresjxG7PnHGi
dcs1isf7/QcB1UlC1BakiWBqLIN4MQtBb2bOIWkC7oZziRwHHAQRd1vn6OUuzOaT
ZcGXTriVbxR8JiKg5FzmH88/H2s0j8TRBU7bjFY41MurEUjpmIbhs0N96saPBKwR
WetILcbC95JfkZPbYX6qfn1nZUXXk2tkhXXkpIQ0IQtnl4wFb8ANI6UDhR2qCwUo
NUneYIJQ8GmvOAfuFtnPU8tVzI2iOLxWkUEvlZGui4UsJcf1HhqpacCarXbHIYNB
LctF/osvPbDXLKi1xzUQAwXxxlHLFEEl12ItEIbxCclBNFJ4ObtT/VNKfJqPdFVj
JdVl/B4KK15jPdBlKUb+KWQpQ3hukaPkgw0jAmGfIcNilMMz8i5E+DK9LSFZFofP
BgMhSnGvxaAyMDSSQcI/MMSKAmIHMkHdT3bM9RaMZ9ddLKb+zffSgV+qx5nnq9Vc
erQMDMa34gAUzca9d3WAic71zLY4xg5lZOZvHzXPpPv+NdHiXVmbwX9bz97LeD8B
HcssDA7s/HinibRhupMv9yqVTucWmoXifTpghB5KEofcBKZo0gaXBnqOCpaZUVg4
JQn80yNnKnlv9+Em0XNTfjQsvPOmjhqFxWynmIWZgRPJWqUsnqA3Paig0KPnQY2N
E/BpRieCtOaxsErhlTDm2C/qHp1AyKAQppMkkUCP3Ood+UpHRY0GpSUP+tMox7Ky
uxOhAsS/0c7WXwQAY8CjAWaV1dvtOZiPSLdew5O8/fOl/7q9nyVOHriXHiog34e9
DCMbw6NIYHnoC7lUTksj/IsSS5L24qxxjbGXbYbQoBSQsdx0xKK7ncrs2/uZC4Hx
T9iGclkYIvcbx6o68sKU9mEUL/vGPfb24rG3wzqfXv8=
`protect END_PROTECTED
