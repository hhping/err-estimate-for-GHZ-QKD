`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwQv7sJMF9SYQx2G3GWNzSEfz6jkBdCBP6Y9OXmoZJ+KhKdgvZ/52v4CPHeV3zCl
E1HGxTEz8CObjRAMvXmdCWUDE2FSIiMeLR/CtiRCiz0C/SlAZ+OpQL2NnRt6pBYP
utAerOd1x5IIUEUveJgeWYkNsf8Eihs68nZZIBYWGBeUwDs/qkKpGp2mmdmiU24Y
/U8V3aomAullGp4UftDPqk4xOrbLyeBPibJW9glah8iC/vo3UYJQL0ob0BcMv7EQ
OmHKNaoLp8sPSwaF8FAOx87FO0l6MI/TyDwZ7xwrJjGftf7t6JltVFU4F+xzyHos
4iUhxrFHvR5oB6ODyINBABsDTzJe6mrbXHn3afa5s626JfaY+YAMoiqdaj7wGYer
MMDimJT/IpZT1sxQqq1HukwOicobnIKmKjqwqHFx/rErrooSLDDaGvRp49+FDvhq
0G4m+QLCBv5oGz5SRprkkX9/8ylgMuwqbkU2JVohTRaU3fCwuUSRTNtIcn4nS2EQ
R+aHwVnHJ4sYcjBrFe3IdupGWeQJ8ZBTr7bGz9LQ4ob7caZWmHj0FG3p1s/I0Bxt
n/nIB1NQgtNPPgDT43dlGZQm/3f2dfRyD/nKQvVkfAIpXOa/SAQVfII7I71OL9Yl
3IgPny0Tv8U9aZAUgyxTytXyhKnZMnXT/eHnyM9f5zqxHV5/7YPDOppPCKttfZQx
6eLz843BtkYxmCgJrUhr33t3Ohbb6LTU7mIiE5vqHD730ujIvShVKYtSSd8SaY9N
VStBv5SP2RiFgpd6brmkLDTFznKI3GKujLRlbAJfWCTr9pqspG5s7gpEagXJsywJ
Phx7mgQ07Mk1aw3qVnNRwFLtpEjME5IlIyKrz8JCAGjpdaokm49OfxVrLgSrVqXa
ou+kJPUVTktIp0+VK1o6v0cqoB7hHnd6YskJ+lXTOo5AUHU+EXm4xRdafGy4O+ei
DGMwamxXmgqDBxjfOoy7JPTMp3yGBh84zL205MWpAXksDqRkBS+SSpf9/APjvuD3
565tJF2vLa2+Fl9M34xwu8sIPZFJd1OdH9RuczL4kxPe7QGjdn2QSBj+O38a0gQm
gBJoFVqdEXB674g950faKsl2pK96ToKE+MSzqBlsXDQ3dkH6HMK2LmXizdKZypuO
6g0IXmqToCcC4aBR2vnl1kXXuXzoSJctY4QZ3gDCWmhc+2OjHLgVfM5slVwxx6yz
f6CgRtMB/7Xn9fOCsOfCYk/cITxZ7hgk1pbv9Mga8iuz/Td4ArBSGJHsgihOfZhg
tBdUEvGxiX/gJ+32LCr0sa2IWdz8t6j2L9eoh1U0FmvERN3AxTdg6/A+QDpFPo04
FHFVQQYLo6cO7xjGgu0q4FJM0Vp8pFal8t1hjLVVpvIggu49zgYenoNqgkyMLZLN
XE4iTTSDwHNtVx19mCn3ap4UJr1E0QenLjcRF6FFx7Df89Uv+k51SJwWjJCfHXV/
X6rqo70VSOJCbKNAg+P8FCYZ1w5e1tdaFKA6tF9TMTd35oi3PJCOicw6va5ESYlx
ozQ9m7Kf+etpdDXz3LNIuJnGXKB9wumNgIMMreZGOw1/l4s0bCM3GRP8ZlTr8AXt
DwKMSG5jd0opIV8Uu4XSIWbzV409+8vPdy6kweQZLGiACuMiLj5xXUZjpaW7qgQR
62Hl2MWuDF2IeAVTlUYoQxbPHBI14lLlVmXrLoLkQcPVlno5X0LBWB8ukrp3AwEB
PIAP7X+m5ozCWHxLiXP1ROb4s1ZZk1Rxmc/JxDd+Qvba4cK6AJI+LvlD3YstUJiw
QdR0+nAS0+AkEKWRUG1J9e9ruFKMF+ACDPAAzXwAOmG4YpIp5P6XQLIUBzzRktq6
l114YrulvCVriAy0/dnH3OyE9wOSedGEWpHHgwQZCnGaWSjth4Y8y19Bm5K3/7ac
UtOXBAbRh3VqR6xeSgWOyT31qr3GlCHPigGl28qX3+j5+d9Zc6BFZn28nsJuM79B
GHOvV72Mw4kPgTmfF0cYn8+QDukEqsa0KOwAwp+2ZOX4pSB6B1BRURKT+3Ye8ukC
+9FgKEC6YLvew6IxGG38r5UoKaOr8RvZ9u/Jb70sJ/gk2YPHoCp6b31EhCUBe+vi
yAtPnE3bCUdbU0g7qyHOjmak3021H/bq3tf10jWtOJDPLCvr8IMP2xjJO5K8LJNE
3BwoketdrEogLkGLJQjmeglkJQrWIBoQBafpYjLX0lBM9F4YIKd5/x4W1IfzDL5t
EoEXY4gWGZjuVXpMCIm1KkzjzKrh0zBurtCM5T1TWp8vlIsN/kqwoTRrYNVOGVXP
L0TFVxddaEKceXKy4Fmvbeleqx7yay5NdeJPcq509kodVkBKwOMDTaUU7GH459mO
CskdMsBwEmYiQjbKkGozR5rou/pR/KkGDy4lHInpsXCcsh46xaGuUq20YpmJeZyM
BV35JM1meFqTHRYtGv9/1NV4eq4C8uvGyrB1Kl6gjN45ha/vX1FO42mjAirorWC6
SM7yYDBV55gCmmeLBN/BuixuUAP/5Lsz5sT6ltMJpgqFHXBaiTYnFTp6YWAkJ9DP
AX3Q7Yiks3ZhAu2QIaQ2qbmosVLpaqBO8hwdKr8l6lBe4iB07PISwf0XyT0yi7P/
WcgcLhwGNjJdVGGfhZLvd+9WWF2boXgld9d9CQH4sDH2rp2PukLCNKUhnK9/Pg/x
WvnNmtQNE6PiRjI1ta6DtZlA04xj0kVr62+G/G6liS55f08kUFz7XztjAaOi4HP3
h8fpMuGt358GrjGjtSztDt7TZ+qLc4aFXZwgOjt9L6Sp69h65pYIAP9yo5Gtiyb2
`protect END_PROTECTED
