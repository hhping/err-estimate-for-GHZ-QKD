`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M62JC7nBpHxWyXWY7H0RN+uz385lxDn9YjLY21iJtKDL6A+57T89vpJcE6qjlLug
fAIg/NXgl/Kyx7IXLh8H7ToAWS3akReJYZcWArkWVvkmGFh2w/OajhTnx5/d+VM/
FToFng+UBU5tv32jQYcdrmmSiPlUlBr7Lqhsq3csPKXpC06oq8yxLNTrm/9dMIfG
G9Q8hahSlvtFwJvSBSe7aBmQ1l9HpW5LizulXPIfnUnV/ouOabu3soGmh7oEyx9G
M/rRG8kE9JJ9UJFc0prk3dVW1Ka13Db58h4gNrAJ88mQ4JmtGqOmO6wn1DGBKd7W
LT1BHv7h0VQ3xM5RvrD9z4x6wSz7Vv/6noQl8Hqo/Ce3vF4dJFZKF/PVa4c0ZEq1
BjSG4tbqw0+4pXQFQBoZcVRxUvUPkK5eYo5/NOnufB6xFlK9ssgm99/X7His/M+X
E17WsqvmlJMLVMeb78XtV3imwa0bKkviGQRyDnlJPnJZwZwaND8Oa87c7kRt6bSE
VChgdxYu77pyHKa6Y5mW0Xivjy5T2eFYxrrVlcz+dtSMSXp6i5aZsJXtHwUCeijs
mNPtiNpPI0nSaK58tG7cCObCC7/r12OMV8LT+1cJ8OBIdKYUHngpVw7/DcedBrmF
UfrJMdojlDOUvWsrsEsadUdvMH2XQqlZYdDBv7AhGfYV7aOnA2bZEa7n5ab6mfRB
wBFzJtaVsxYUUR2QsyWdEMwbWn0vL16Nxm7cYI5TjUjDbMj4xpYM+9YZhZkQoN/B
PgOdy3rJ/JozteZz2Yf/UV67u390F+87ld5JE7XEnTWmcgUOOZ79n86FzcE9z0du
4ipTsXauZk9jqEGGrthCGesRznmnJfEMac9PsuDRzXfYos1n6Cgwxx6R+jmWxYEq
X3UOw8mQKCHy8A3notTfnasC8Qw/kp7fg3QskNlSCSwwjF1ctSLAr1GzN94h1DRB
xtzblf/ppBiHLiYuq/e0HqKhOfMCqi3tYdjQt8FrgfGg6LhO1Sz2LLtl+GVHvTp3
HDCqSN1YEfVupsG7I9z6OpdDiCpDrkvk6uTSkuIhVGV+TelAeyh9wbKOB0F+WtQS
kTnyjj3V2ACcLiiuTuflwt9lhhBlLaspIPYUxdgN/nNf6ltb1oMyicnNoVn23GRH
giy3t+VJ54nfHAs6qNWKen9C+GDy8Q680FojhP01qR0Kkcu+XWPl4b16r6BNpB3Z
w/iV1yR0lNt7rg9PzN+GiabHm0TmiMhGHKm95FYtYHeT/aMQhWAGvEd102guRPbu
11A3HlvcxYA1dTUY1FCf1d/wkanO3H1BBF0gnQNUxCZDPMj7qaR/ZKLEoiDS0snb
mUTcDVwn84kF7lAMmax0ih1KpqVou2wsEJlvBvoAE1D7TcoB0qg+zRw2UVvM+lf1
sDuOZtJxYQf9sleMt225PW5zH9oO5c2oVcWREdoDKN5KKqvTkGxAvBaFtfDy87MH
1+6xffjV7+v0/6qOFyMePEIbmTCg4Lb07UrJz0Fa6pGblyU1lAVO3mpI/3UnyKHR
BG/97LQ5g5z9/dF2qeh07c3JhHRJgxvinnXfJWIxje149vIGNgM0L19S72HgvQFJ
PBZ5dxIQE32EvZok6ZAdbnvB0ehRR9tatAEAH0eDPl67T9ZaZLv3PiASfBqxYJLV
Sx/5n2sg8sZzdQLQ3n+yyIvAOCZdtEVDHhdEyRexrLOrrOvANnb/lEREAcLSkzGV
7O0P0l9isIVLbf48daD16wo1y41Pk1GIc24ZZkOkfR6qur9h/2IMH+20TU5rWVEN
n9187rJkDHakvD4qGmvEspXxV2b+w0OwhSzSvseoS1BnnOxqhekfXX8VXQezPYPl
q5qkMXvRU9nzYrCRf3puKZJASej2LkhPrMXKYMqIT68Az8IbUtJyhfWcDSwRMT6i
bZRQJwcEcmTfbfPYUCeKTkrW/WviUossSSoB9mxEX57wr5+3GCV8/BpR263zysGT
81vdCSuUizbvOPOpOa299M47nPRjXNtt7FaKh6p6EY80EUyyTN8idgH6RZxZNa0h
fIe5Cc9a5tU33ouPouRH63up1UNQckQQNkTWmlO/1JNI1xZjObDS772suxlNcUKz
QJ2v+rcK6JLk/pgBFJ37Mzwio6KsGYKzsv90WkCYfHAppKBA1qfCymwREBauzKMY
pkLpa3Z6u4y2ci5E0X6fRcu5795dK8gOJR+gyZmQ6cSxycn4JQ3Cp3/ikNeW4wSZ
T5iNsVXZd0jtEOh+KK4EyGnTUxVPcauIKYW7LeVIg9fdadcs6g9ktOVterbh/3i1
T5xOFiyV/t30TAVJSveDKduOzP9lQTskJqjzYqsmLs9lN6y+roRz7NkKo6O8puN1
vGsz772KN6UT2jgH9hu104mkPsCa1EzuscB9zfeRUNE7BQ1pYr3y12UDVweqbfWx
FYPvND0SkrphvkoHTWiafnFjZ36dPprFT2PhnJQcH7da4f/aEBuewgChF4QrUBCa
9vCVc7tVKB1vvZB9/8R5SB0ndM49RYkzvrZbJw1gFuqEVjwzJimGCdIgSQshcKWl
imQlHBRuUVFmjgB9q6Ofi97+rIAOBu7GHquI3e4YBFj+HYcxygK95erGeoB2e3Xb
MqK1x7s1K68S/O9n/PiN3zsYBsO/C+hsRvJ/nbjJiFV2ziD6OIn151GP9lfIi/xN
LnqeV/G43s7bMDwR7EktcCVpZaWji013ZEqsAVA9tq3oOCJERKIr4OCln80SOYZW
sBf5Gl9T+8FEYVm3i6Vr0loodeYY4tZwMAU/cqoB2jFsD04YCmHjtHQfnQSc48mh
TsG0WO0QgCvsWY2IzVtfKJL3tFtsO1kM44GgVNESySuCvytrwgzzEQ0piWihdRwz
K/A3T4Qnyo2eLLYDGoat0SKk5ObF1kBKzmjIY8VCdLv8QeT0IPjpqn6u5yfH8apT
pakI4zgGnQYULIt3xw9JkJyT1WgLrGA4YY5sc6UmhsYcNhmzuAjKpaDjcA5TV9uX
VClWNQl4plc1SElk6rHR3M29n1qth5I/AMGoKUeLABGf98dPDwazk9j+I61uRl4r
AQ5QmATrcoNZl6qwBsR3yA2n7IEJL+qZiHM7mMJZO8iCSq1H2Q8JUefg3f0d29HF
IqLrj6qZxY0EUqr5c5NMyNYOFiOM6Rp2ekzxBAEVrHAqeMV9a7IIDN2Hah9JkOKt
ezMRceY1L7IIEdWMWtVKtAhjoe+2wuuDDXtrDlaUFY41tK+5OWhnsGhK+qKruP0i
7MiiOUyY64H5Pliqup7jzxmsxQEaK1L/U0ngahiZSoGnP9ewCO3dwfi4ZoUjdyFP
Mhj9kKy/8EKFkHycQohw4oG3mWwTmMC7CN5ZIajgaWlafel1/WhQ9v01MaVm6eFW
64Pl21I4AGRhiKztNdtDMWH/B2jMFm72a2n52BU5krP4rtt4pxLzME9Vd3p7FqIl
P2xttnDTfnSHbLxVEhEY9u+GF2cQTLR4ncGK3qOFXbSZiIpyEn1Gjosp+BqExE5j
pMH7UZg7QY+wXqMRU6B7g7VHriO9QfSrrxPvxMVWJc5wUpsEsI3zbGh1i7LcgIz+
ZuJpwOWivChA2dRhr8LpKK2hCGyYjkeCo/88qsTIhiqnupCBu9L/6p/dSJMIHAH/
oWE+yPy76yfpwvsOkFXGFtWCjDeN+ugSQc5Uma6cPTCATH1YHEZPyn868zLaWEYQ
1KVSumbkd3y773XeJVc4wvXd96mWiT2jhwg7buhYbidAALAa5+w4gv8qPbs2VcTW
SpoSU1s+B7/KMGUYRduIZZtcSqf1nwsyLpXUiB1502+WFd6/rBeTrs36CEanpujy
kNVkWAnNn5D7rgeetqStx9moFQ3mHEYUuYBjG/SabV14AJcPFIye3gvlX08Gl/vz
n04Lj9JqW+o2girKpZAglRkTU4xKI8V3GUSVmX/0t23Q9t3TKL5MNgs6v56JeeZE
2u6nwQ8jjt+xoI/LtxFKEVV7vMf9f3F4nJ4ijJ7FKBZCzwF7n+bjvra2gxMY4wgv
CKa0B3eJ7M7t5hnS9jYlXM4Wlw1u6oLEhaFTrGOGe/USGSXEMWw26wm/ogvxTamn
l4pqaLMIyrsbIsYzDXV3sdPHrRN0ttalejMdl9/pgQskxyeH8t2s8BvP+bMHhANe
cWfBmtdv3wfxL9ZT2OMvDywXSoRwiNltuic5HHR34ygCauj5vW5vyknQAstpfxDK
SNy24tJXSkHK8iOyRWqqKsgv339CD9Za0e6+Ud6eEl/0H9daCe0HAEl5GAly48CT
I9uoMQMNUZ2VTWhDDo05hQvWqtI1bdhMTwPWqXlJ0R98SRmq0E1CZt3urGc4TJpD
13OidrSzFkKwuj4alwwq2N1cIXIEdJpiFAc1I4dd/D9Ng+AaQt4EdV8GCuFlCELl
O5gwj+kxidrl+jd8c9fnwPGhZpt52VIBfCn+wLT+LhRa/Y4KKJAr91MM2K2X93Cr
YDP+IEEn9QrDy/+iDqMNUsPEQJRmShh7m3yqJXGAmTQdn5GtUVkk6+1ex7zjG2Oj
WSdEMhYy+To7N25skwGIlX9NhdGX14jXOfGh514KLg4Vjr42Tpkefsd0XPbWD3ue
OIl0Oswd9tCMCn+z2dJLHaL+psGdtfuCAF656d+jajfMgCt8YGUiz3khAxjBcpOH
W/o0QJXG7baxkce5FkVGcDwPHH9OXZ7251VrOyvTv2qAaX3psc8pb5Iqz0IceZxk
Qfi2D9gUp4snbei6an3v3aM7x/OfoA/9/x1P4cIM+PqFyHKLZDT6Bgrk1j1cXcTI
EXBhaqK/vcIaJIK8rgJuVzs8B+Ek0HekbrET+CZf80P5gb4ZgkumUOT+Hdhq/aQy
Sy835vYa734WndJ94KKY6i/TCk+Tmps9Of28sYVje4/MCAPCTChgEmaBSvXezt4p
elstp6YrVwC3Cz6mA9AHrLeJGZho01/Lk/yyGFn6rG3sLzD0bvlxlI3vaew3D2TN
82C1wXXsy+xwNAXkouRWDmvhOjlsTZqJkCK32Gu34M27bL7LyQIaMxG1GYOrbRCi
sCIFYiDB0shu1ladokemgtmscFiCtom5v5P8fFAAAExvvvaouwv7AYu0VZqLmRLc
8O3tumSe79jbeNKP/c47wB4fcXIbYLbLYfNixM76pp/ZnKybiwp7WraFA4fVS0SE
4zIVrcjbXYm32aYjMh7cUzJYEHnJZLOABTejtvz0C9A4JPir7h0f8jPYBsPTRp6b
V/Rn/NZEOO0tDjakqCAXytUEk9ABlzRg4V8VEiqHlB4+1F+T+75MOWQ9uR0Ete8C
0lMVSL26ZBmxM3b9AFrllrG1pPtHjVx3MJUzIiQcr7gnPccjlqPyYA8/ehJQQssn
+JVWqhuy7riLx8JoDdVaG1G2BmNkj7uMlNTjQJxBEAtByZHLDLMwls1rbonSUAsZ
/vQVxtFYN2mW5s7iodFNX5N4pxw5oeMr9TghVRIu2metcZ1JXhLE4MDIrDP6pW18
f78xPvmu7LzFWOc8ITHKb3HctrADhHuTw1wrrCnmAvlbxmIUc+kaWA824bCVn15X
8r5TkUq+lMJYfaT924jKr79MBF0PyW556r6SxAN5LR79jxf1diKHr07uMPc5iIJ4
dkfRy2/dWFGXAUjszgjCJ3c+tLps7ftxlAdcqOLIS46kE1fNGyKHT+35l1ORL0N5
b6SpkELlXlu3/hvyGvKTYWaHKrFfVbunPZzuady2LI7/F+NvrhdcjgxTZp3IvxoU
j4DmnSBJMa0azUra7B5nYp8e3F9sMeUucLu/oRbJPwNBWpOKFOLmHUE4QH0GrRih
oVUOkWf7eZ4mYPeKMK6dypjmg4MOsyfwib4RL7vmxzn52s7R6trIl02Dihnl/6VN
60LHEqg78eflJA9sufrHmr7m6GiMEa1GCclKuOdi75lENJbV5iA+UnZQGjlr2QFy
u2+5qmatT98L5HCINmUrG+1u0QRhpWubMPRubLuNm7jJy6YFyX48LvrJmd1flXJI
QETGgPrsT+5KJfSW8sgkraV/YFlNfhIXFCWrz9n1S6S1T6qbDveeQlRPYIp5OwRQ
zLMH4YXhLYX/SQbaKOFovf5WDhET5nSp3/9+pyayBJwf25LoYRvgjX9lWJDI46kh
xQEtCWdKwSacXcNbJ/FkzkpDoI/6miUXPqKC8KhbZTvhZMbxCu6TWoUjjRafPcA1
1a5ZfHarijpVZ7JSwLHchKeMRsWuRIljvz6X11Ehdexm4n1RNcCNPtN4pF/Rj2zb
1v/GH0Kg5xIB57FQrib0FfGbAsSsSLC9hEMbbPPdAbsazEsHJkWog6+bk35itixy
zifraVaqI/qt6lY9/6miB6C9vhu1nnLgXLKnIJkof+9boW6KTnYVIExKERqSeeOu
rmOopezgzJxkrPZsi0Z0SlWd+RJ0dMcjYTlvpYAZBm5bWDONocD9N3QrsE+TBV3Q
gp8gmy1xnlPhtOzAStubjAVhdrIO1pcJgSp05F+rBK9SJlCIh/qCztTHDJzcNsgE
91ZLC+OIRZnptDgz1X79Ep2hCUlQX9eaFDqEstIhbrezyJM4bkVvC1ipY7hPM7zR
5XYJRFtWgGf4GZ+zGrnwmvjBLLkEKmjCS2RY+NyYzc9B+c578nbMzaehNJNlcqEo
JoJTtS9vm5d9NokA3Mswe4OIGZ5VIx79orzEIjBtri5FbSJimBYm40euuGv8R2VP
tcAfAW1TQuHVwGNpOEP5Ma/V8zZq14rcFkTdx9s0z5k9sOBAugwoD22LvsDe6F6l
MBzlV2h5M3+Ow/x95jgY3VvdyVGidMD7V7bjFgrMUo9GCToCWRFo3Eo5gvXfOvSs
pBErSe/ahBqIHuvFcp+Loq0YfgvPnw9f6zxPyAp6AGKhaRlvIVLyBVdrJB5cojRh
nMRrBAIRoWtBPq0Bmzwa3MNyMD8NutT8d0/aBruLF1idba0/Qybylp1NyCKWFyMl
AzaZg0XTL5NQt9ugFYKwWUjSgT6qv1lWGt2gO3c22T3vDkpUOT0N+HL4oYKnArYW
PpmJ6HZxOIueOIIHqNxX+FqQJWnwwdt3aP0wNCyGVuh3xoUXayvip5LIGpkv+vFJ
CL+c82paDqbzRdr4++/khf1FPDJfv+mdTkPH3dYn4q8yN+9/PdaxYPzyljkeARNT
omwG25aDHT9L44nEN52Vryk/H0lmLPquYrAr/fqschz5zZQ/VMVq+x+OZ8CINadx
bIUD8HtHcibqXeFKAjDzsAMx4GbNCtt5aiEUj522sfDR9YNCHjzYouyarESfAdh7
An8khUjEZ73S4JmzyId3Ds6orObjyG+aao/pjJK1GjbI+/Gyd3bK4yyJ6/4Y5J+t
YyRRAvCZFCDHY0XlVaPLzT8490Pao9bzzXqijS2+aEMNaMQf5C38X/yS2BbOzwnc
qQYynlU/KiNSsmftZF63as5OsZXJSG707nFPvLAV/WJwx4Lryx9R2L/2tyR5QNQ/
PUHNYhsVlJOoIH8Jr0Mv5yUKXq2JhR9EgSJ/3pzFj2zScGc6p4EQ1ljZDgjt36Ad
3+8HwkZEXc4jMfXwIeHnqzwPGC14mCDXPVtlWE3w5UGTgptWcUdXngVfC0xQNX2w
2pZlelzctGMVGHfhuccqZvXqOtgu45RG52M31eI5PShUgzEpVu+s8W0FmcXjCGpG
IzjZNXt7qQUy47SPneoOC0KBTagu8M60xIZzEj2GPGihwU1pxXohVl9yUt+isNnp
Ejq/u6XZUQMC5vvqT+gZpxx03YJcCMmmN6RDHPhgZHzaAMXcN3aBObk/d//2jzGX
sgIAHaS9+l2aLfVg/bTDH70z7Xu+0Iga06K2CliVpoWGnRm4GrOKwtgamVb8myqV
v6R9ysfVV0IFbxm8xlFieV1dYuE8ak/UFBb50h91Yqmh2Q129xksbTTgwlajiH71
V5inyskc38bfd2KQpnQrXsa58YIBOutYBxbgtYOwbOjjiy7fS4qL1RpG5rOB4FQN
oDv5mDpOXNsPENSNXo85Js+6R6L4hrXdE9P9yF4TXG9Hs7eI6vX0IUovCe9V8JWW
qwST7czG1zeiFZX3k9odbo95bx+59tnHpFCT+d0O0nlNH8QBxOPponnBBNIZgj3h
wRp5biw4Mw8/bWjg6MnjeDB3x9LYBJr3D2FqpTE9A0r3uFb2oHhrom5OHEn1qHmG
hTU+xicos8z+LHbS9NKsF8zJ0llnBguCqCxkvKTGVT2fT9hremyCnvNxgD+3dc1S
FPkdP77+iAmURPdtcTh9vLZ6QU5V68UqQiG04bXLxK9Ng5sDmR1IbJGjIRkIq4/Y
eLl6s3CTpzlRWs9wqlB7BEqughaRkLiSlVtrwyZP09IclCKnAbkM2yMEuigS7bmf
YiQ3VWx6nysg0zJ+/4zaW4GsfvVyFdcy72R8hLcm9peM7wkVq8qIvY4LDKdrl7RU
bvBV0x0tuAonrqONuWAusPKMfSfnS7hv4luPaFykEGPFUn/1VcwUIihmcgE+EFUZ
NNOPKLrMkuKCAtOcorTQ168DvXVD/JswmhT7diihGJW7Ktw5uZ6//1bhsytCZM03
tm7b+9i4NPG+TwqaPuorEqeuPBkJe6R3U99npydkt9nguJSV5Pk/uw+JYrSwCXip
WGLiqQohdPPdwJfl4XQ2KxZwtOamkz8JnlYbST9CqUNjuAEzxDPmw+XdJWQeJhaU
R/UJrP9oYS9JYyNfKuEpw8CatIh48ZwlwC8v9Igl1bf0tfoVp1MJILAjcoBnKqH/
DDXD5dqCQZBtS4c3fdpvcKnVFvbsOr2Hh7q6hSMTYrOdCxQskppTQpU6z02ciqs0
DFKVXEMKugR7mAI8cwu9WAXNbbq3/bufowLD28SRdXN6KR5D2pJxWUVDch+m2541
XhPeycb580srWI7IdDSZIUo23QXQX5sHxC7w9CCmXFVLJ1FkfRlOVKx7LR+ULM36
YZVlX+Pkwqbjr+Q545UC9IX2ETSLs5xtATTbocb2SyaOqxKHHQc1r47gsIRyehoI
DfU3UgfcXKxjFF1eKxLlArNzAeMEkrn5lx1Ix0zqmfmGlw1AiWLAEQle7HB6mgo6
oj77f1SQpVKvtAOrGsvYu+hK78WM7Bwyc2Rm9GarzDIDUvP9D68grjiWBDtzKX4r
YnC3pVxt7OiwN6TiQUdFxq71HT1gFcTMdg7ZhtndVKzVwP7nowGZQ6gUu3n50W1m
4TCHOjwQT1S7NGCrCOOzPGjpAqwkEtPypYMcYmsfLCOE311cMVvosdwTIHO3jrmG
C0ZjoEwHCOifJYOsY97hDKL3Bpwo21yGK3xXZk90GFAdPVKJ8on5b3om8aVNFGMs
qF3YtiJf7BuYM53inP9a65Aohf1qYZsV+R5+wqJuMfiLIlH9DW+0gIw9VqFS8h/k
jJnvPY8KekoSNcJWMJaH4+OQEgYLYsukI5lZOJlR8151Ywr/CtOt2z5UURQxCa0D
gI1P9iVzUAqh1683v9fc445CTLZ0iPVFoHK3H3a7C/padg32OHEo/TjADE3sOMS2
yIQ9GeZmqFnziw87gnMX8PGMufyCngwcohXfdJWmOYAz9GIukQTiKid517Asclsj
/LY5wAE5RMHpb/JE365cXJi64sNp7VUdyKUTvORCtzWgTQBDP3LcrqLDTMVrmw4p
W+dL/bt04ti8JXsfa7OCXnZR9hk1D23xL69b2BhGUGN9EXkU3vMBkxkNtHchBkdS
7Msbu8DJi8fQruwZIPnz0s222BuibKDzrVjFGTz6egoF265gBn0XwlWbCEoO2mtp
Rub6IFfATkcLDpkkSFvU37SrHdOz6rPGlin4fvZyrLrqVwltjmRIYV1ATKh1i/Cv
L/zyl3hNw8LSw8DoWgxaBB7oqM9jQXUPoD2LrkjM6j8bsDyU/QwaqTA/jf5RIpYc
s16HeWVrDsEBHGz9stf/YQRSWgtW0WPdtzSh4SZXNVA9Wnr9UT6c2Fo0SwYHYa3X
veLJ6S6pIYVcMcpGoDJPB7M3wXJ3eU102t2v3P0ZHd0aeCZGr/1U2f3H2odR5OHC
uRRNbLVmQcshAq+1PlM3btX4TKyfjcR0QJxBeEMLGc+Mn6oyRdrFCIv+d2PwNdRn
akHngYvXHh8wYIOPAepDFPQzlVYYkQ0Tek4/ZyGoDEQuUyJxAwOMFCN4VUPKG8XG
KolySl1vJEimTAtx5CRp78LFS91uh5RUi8fPio/D0uhiCV8MV4BP36JV5FD3JzqW
HmAnx2oV/2E3mIxv8oZoyB0B8wAK9b2T1wj0ihANC6kID5vHIU+WnGFl1s7rKd3N
KX4MDYkeENJGEF+TlPjf6JTybcJ0D9zbQi7rx67ZKtx/jtiY/EN8XLG1ZUpe8VON
/5pVqZHEmQOa5xOFKm3LjHoBfH/aVanNhyCVUzFxpy7/edA/TBdp63ALyMm5Hx3r
S1XWmfEV7IzXu5TG+7p5RL6MiR2ONc0p2yrhOyEeY9unnkBAfHbJVPdFkK5XLhdT
+A4fj7a/5bV6EghtGbjNsF2vTNbdOb15I8fb53Y1oJYdUYUK01OKKPRqAglFYwjB
sDspe4+FREq5o98Jvm86gDe8G4d62D1ibv8hgz1rJTcTE1dtxAOirxEwdkg+FRXY
1e/jzcJSHShJeVnrTORXJv0ZtpBN04Lpr/BY5VIjS1NL40a3+HuiBd4MKvbOn/Hy
SPXFGaDD66Kny2/Ckg9U6eLGo+SENIfCtq/5wkv2gID9e+nuoaGHvtR4g21ypqgN
7RXuGScadm/3TQXBMSQWn4DpYtnjyOsQKTq50xoyv2ZVEp+xODwjc8aFHw3XGY9C
jYAUiIm2h2xYzMAh2tzgCv1J5hraUkJgo2md1Zoq6bO/T/L70EOLurE+ak9VDbe0
ApXJvSeXx4mCkdV7f0ZRhTuEzvRihLS8U/5oBs1/4WFCYE558RHG48pQashI5CyG
L9bdY+C2QfhKRx6fsJpJ4qN4qJuDanJgrSoGMkCqttOp0TTyLtP2TFaxtYBo5khR
pMXXH0hBTOcpLQ6usZJowfq4i7D6ddWWkVllNhIwk5RzBBMSifBemAnPESK2cmdy
A8eNEEduz+wrkrx7lutc9ghD9m2WJ1QtGItYtr6BdyyB3JVTdXLQmwd9/KeLMF71
da02R5fVvR+ap1T3cPWaPBiIKxb903IvLZ1MvtZrmbbPizIybmneqO5MrCc0JuWH
lLHq95W94jy2oGFOp0bzUOew5szA2U5QgLVmOK2sEAI/bt1MngR0zwSnWeVTBWqK
9hb/hvp5qyp+nBwZIX4nxE/WWLhhIVFR91P2dkXTl0BYly15zSu179YhRBGThxXl
meNbriXVOsWk5xTUoDy6cemC/eYHGdfqJRE6U5Ss01trKZOdCFBQiGOH3A0ElB9O
ZzmBd/4eBDvCJC5oYUi86e9TX3KOWloHSqalvCcSjM/PCGhxcF0iXSFAw/QHyGgu
/WYTtwElUpNPRHpvJwnbQ6gDyJLEs0jDqCra4MuHUaLz/ROUaXUx4UlIYjmHxeNf
KU8ZXFyYy2+p+RppmKKzpXq+9c6syR6rTRi5EhUZoXUDQ1/7afY1i52upGlZ61TL
WR25xlBVtPbQvLLNLqoZI1h5SE5TOZjcVRPmACDxXIjyO0qEDc6hNPrs8FTzA8G8
bwX2pJ0zEm+owofJPL6tS5cuBw1A6n5uOPgp+gnpMYj2UCQJQj8NKCw1n+twcNLO
JkuO10Of9FH/jeN80rHCuZIXUzOu49+oGQQceB1+xDc0h8q48sC7k46wNjJI9tN4
9L7h/2guGZSqODV8C0k++2nZbCSXQ9zJPQefwXev9lta4aghzjz5MJqvGRgse0Zv
cg4oiRaUEv/HlmGQ4SrBvhqM/BxELoKNNNRALF2m32HDfm6ewT3t6z/jBBvMCIj6
56LCgFFzAIgLmRiDLznA7D7GqWZwdqibHD0mjF86N24CFosL3iKXUgr5UIl3Zygz
k2E8hOJc0bnHHQV9wQx2c4cBLrIAr0k1mJomyZs30/W9PZb98CNpeWA01YG7Id42
zw3vqJcB252O9HcotuIaXXBtPJp5hbnX5YUf7AY6HtNyvOYe+/SuVATUDT+euI9z
k6S27ltFEARWXwQ9jKdw1hyhYFYNshAwaWUXJb2OCGDuEdziEEFwf1TLdRT5Lx7b
Cqgte+tcznxiSbCRuo2lAx9gJJM1QKSgWFDqtsD9pTHvjjocXr9oFxOcN4bCCDHe
yn7N2wWYke3QoIklWJWp1IV8gCosSOVYsPYrB8JfrVaAhRfz6GCGbcNnvAitcx4h
GJ799KAGItWBpiqStcyAvrjxcQ9K9suUJtrMZGp3UHMUskHmOxdoPgv13JX6gwby
SblQ9ZnNV7hN3GdaZNf2tfrY9vVHBWHgjDz8DGPWtKjLzpGIteocroTJrLoWpmsS
mt784AFdkd+pW4ay9emPiuybbFwHHdoMcUpEY7SkCgnUyJVOST149016dN+E/cBF
UGH0vymW/4rDlWx70MqlZ4uPnZFkrBshmgIl704p4RjzCX0W9Hvh4byNGChBzZeE
92VhSxcgRkeEKJ28ZMnJRn2xMDMfPhz//3L+sUDfRdCkErCF8dBblIDY1Ld1G4pN
mgCGR9XfdiqD2sqWCpuEU3eEHYuggk/g5y72ytv8/8rJRJRJrdAN/5CkwqaY0VAk
E8CbDser68t7oC9u1gXFwI13xdxFM/lnE22nvwH8sP517tkjRdOGXXGZv2X1EPJm
5NJoRaoRIL3TzVBdo350SEAjcjF15Z3YKArEx5piE0XSa9LKMaPI7LJynSPVg4VS
spS+gaXw0iMFHK79fnNypgNoe1bwWOD5SonFjE4efjhM2Z6cW8LlNoo1dYMINK4z
E4L5H+WW2NVAohFZAuplPC2ylDiFOr2bjgircg+0XihMK8+5kJrUUiwj2OllsWtp
d7Q+abDDaBY/a0VnVPPfwlF0MLJVLvECGIqAnfzjwOV0LaFXZUj8OgDF+Z6kOr3k
i0DojIU3PoDgfP1sxmb8YWGN+wKdVwLIU2cX2unPaBPgYgHT/XQkhPzFM4X415wo
/Qupob2bYdGzCIJ/mOmINxlZhmgR9IKod1ErJM9YUPOAtPT8g77yjlJHnB2sEkPv
w0nFW71s6Oe/fK8qQg0htCJYCJKn3Jd6rMz99p1qoPZP7nAy5bS4P2IDOWx0O5Dq
Iz04p0YCFB+iCwi8R2auI3BCU2aW7i2e0uTIhjnfEEHOB/WD8E4vhyED+faJHmog
A1SXd87KioA1+xD/gejeFgOD+g1LUJO2dsT7fCPpHg3a8zIqHYCkJPtTcZL7W3VH
jogYx3ybxo5yRj1YX33yRzz5Mftn2wgCEjrVSVtVZrYj4i73H1vOM0oZEEPxwGYx
9e2HdbruiDIh8CTSbliNeX5qXybz//NxKa0Niee4bHOeWdwT+LGKl0jdl3BzgLQu
IhS1Gn8tW2ePSucqDpoHx8T5cQroII16UD2ls+sMNTLZMiDqLv+xdgQYrvPByf4n
89leqbiat7t3tUC6Sj4S5d+PNF8XdgVf48x24e+fP7rx7Nx5lUWCicpJ+b2f2cQS
MSR/9Fxe4ktikdxcHoEDxv0MDvttiD25GkfxMGsbHd6xNRjCsbAY4WFj1EowZx3r
eEBR3izbOjHPhVOn79MDQ1GWk8auVYxCwQ63c1MLQ8BaLK+vgLX/FGpHs9yn6iyU
WmSCpTvGFiMTAkpvyMpkxLLQB0yPRiZmqeG8jgQVZ2n+L9+LSn7qJsikFauKr/KU
nqu6TjMFIeimbmqHm8Sz/aaAsFYWN+7pswMjAlLutAH3I2LMddhmHsjjAd4GuT9k
I5mk3YISsSMgAE5x4K3q4cEaXjmVucbXndOEg4ZQknje3L+0uCVJNJ6eeFONPrO5
3BuiX7uQEyVOIljWqM7ky70qB010fzWLG5Mx45OwUeylg4FiR/Shh9u/xutJ5aO0
WfwSoU8cCuN6Ruz4C8Vm/jHKN8x4XLA8iwvEvmdKo+pphnPp6bBpdiIEwM1wz54f
n30L+dqSOUdmwgN8GAV/YwhquHytuNNb5TJgOQH+rqNIcCUS/In/n4kTz4LF8vVy
c5QA8ecYassWR2E983iw7A66GG6tCoA/AxAajVZHkVDEm7hEK8LX/Fp6CodCHvkr
ppKWkSESq4bWzm+Alsgkk+C27n87KKTNK6XiCV9h+ncUgXS44v9r4tnf9lqZOIgo
nGfLgkTk/cxnR6CzruiH1hbLKIXnZAYxF2An/drPQjQv7boTp+llzct8/MUBuuCm
qQ3YoD0ssSa9/nwqyCgfzf8MtcxcW/u8kzotUgfzmPOKgKYI3YfS6ZE3ST2mGlOC
cY4wHBIoAh02f5s0b6wfirVSB9ZjMp164qOEQNcukVfXhq8QBnwtD997QfkT7vkr
GOf5sQnqj3WRZ+eZ1T0T4hA9Eie9DHhn65FUGfJRSl4iwpWQhqUEMGGXkpj8XqVm
bu5XKRRD7RlLc0g+SepWxU581/aPLk8Q2rDKlzyW/DNJoP3EhrGfctsaxoIh7uAC
Sq0ffOZ9coZAzhB9KbnVFWYx2NcAJBdtxJpg8NoB5ap47TEeE5dw/dNXnTaSzJ4O
v0yQHQJJYSiugWZuXTz2L9Nqz6KG3SZXsv8l0ZRsu4OdlXLQZLUdKsk0YqwmBV6V
EAkuGZRFuokQck24i1WsMvG/sHy1n1FadjDiPflYKeQHEmnWQ4Spka8bo/Evwtra
M0z3MYRQ1QLZfcruEfDgd6x/9gu/7iCLxCva7oW+xv6sTF5nH5ESmqOwLAQoM/aT
RXNwu4wJQUdvbaBNUxbu4vkqjONbnx3XYXdv8KUje3Ju30wrFwezwKnCgxvverxy
vabj0hkjJdzvy1LeWBED57xoBt+hUuiFIIIMTPztsNC/aOWJyjo+rrtFobbrW1BQ
YicNNocCGs5aVHZm+rDYQkUNed+5dLDX+JW7xjUzMk7tjOBYyKZUFG6ZcPUuj7Od
Y+mhDVTlWjlK/uFpb+WDbBUQxxq0Kp3mWCHGosStnPoB85UcVy/YakHsd9N/xjEI
qyfKIigPteCfn/FdKBZuN0mfD71ekKx5j1ceXCxbwC9sASE6SawzNtszZ1oCl/eR
QMak3o51CN+vYP0uU5AFMqeJTtGJoV0b1Lk5QkwCSN7+F5hoKuEScPq3+H9L2rFO
rV02rVpMCO7lq9ab6hsNP3Z9wRxWzaN+VuepxcP8d5RUGqpsHDFbl79h19wRQGO7
/MSIyDQShqvFLhV3HOqbS6AKNrc63b/eIlyjvKKKSFQ9kCwoDoDNtXY7wgiL0YRP
sbb3zU0kdSZBdqCYPVEBFxvPgCdcvdjK2xoHxwkvnEd5ixQZqOivWgDLmNzVa3EY
ogT4gSkt7zSbHc45cxKT19KA5Ypp7fvAQ4SlFuoA5NEDo0uqzplYnp4Q0AFQISuU
RMZzYyTYcAlEhVc042/3gWaI4uv84wEcbbpMJS7/FdbYPbWp4WMhByhi85Mb83gx
a+XJqcJ0z48CguGSZarUlbdNnQLlGWHATbsJVMphp05IX4gCowY/bdsI7ly/bArs
oP6Z/YDXsw5vNQERVtLazgV0EuLR0cM/GBpOHgMrPcc3XKbA09i4j97OaI7Y8Hs+
t70WC3CXseHqXq2ZeecShzZ0G7n76fe6+K//QFg9ZLFp3qItRdryn82HxyDg8ohO
gBexLs9BgdrjL1ytOLuGGaGQ5jnBopA7qd8R+dF75wOBv3CqPW9Yky/z42I09M8J
OpBu8hdwlDkKmq9H7gLhCoydeRLZ1nQOAMHbaYepm36+Jbl5BalkEr+2uMWJ9glT
h7oLqDRTDaL+wH6+KHJI6h8iNvZfDr4vUW9Zrh6MDAckie61o92wr9LZ4UEOURm8
aL3gIX1S0vk9xq8Na7uuyy7vw04PU3zGsgG3KXxu+RBZiviz/J1VBvFn3ynPMf3k
iawdRo5oFHfoJdJat75rLc+uQT0hKSJ/ITOoM1dWIB9Vz84bF1e8aelGKscjY0h3
YK7bVpVvnHwMsI+qIHphP+G2VHqCIuEUM+bx9UdVDosatSCIVmYMPOiVRmUizSRK
HOelRxlbvBDqVzXTHwgl0vwnTaOyIpfNqv5+WsN2q3Ie1g6VU++n7nZWBj+2xfEA
0ZfrI2f5LH0uWFinAi7uDi5YY+2DsH6Li7BJCNQlsj+uFhbnZEaiDwY9GJadT0hC
VZNCA2YdH/2LOUcLzhxGCd2LH9RJHbvSPFaRfvtSwE6JuyKlM7lYJGC6HgDsSbMC
0/ygYfLSeahtKy+ksN53bJWuM6TkPzYf0qHrBWf8fAOu4RC0KWZLAtx34OvjQsSe
ZaoL8/H0s7DKWpgPHMkKtE6lR87LfG9ItrEc1D4xDuoTJERujceB5PuLRLlx2kya
YNzGbacvM441/1xiTYQwnzAZS1us/BRSP+99X/is3jdsrUt46ZHTNnJXFQCPuuyH
rIHhxZOXvQBbNUwAuo9P63xho/rX/292ZoYxFZpOencrP9U8Nj74OcHsKNHUekUx
+7uzoogKewyfv+W6aqBC5sgptS/oMqXRmFDV+GvEi0Ppdl0Ckzk4X115/25qKFgT
8v2pGiojPtOZvuTFM2zsj6QWnr71qjs0LHUfoTri2kKKs4kv8CJ995v5mcNI60R9
sBqTLuml5jxndYiXoT20HLzQ0sk0oNW0MkJvyaIBwWxGXISubItCvA42MDR3rmyg
QecuF7W9EFrUnz7buxre97DAwhPkrLFgJF+gK22KvK/JV17+JEru289oM2wRhb0q
C6bV7473z18T3Mf5FW/bc5UjGlIWM4cXJzJ+tHTPfw8S5FbXTq01YzNjoauV5Y02
Zh3QBP90aW5wexNMoUM9uvUX3qVqnPB86wqJjjQtA/7fCuW9IcNeX7w0j4mHCXKC
V51btZuVMVzAGHJZuxqX+Cd59SfaHyr6F/QTR4SifReWAytGfqWlHvdvluzFFMzp
9QNnKr+jByVNfijd3wMx4sctJk/F3klai/Q60Z39FhFj0RVC212uc9Ef+TyaGG7O
t7gi1wMxW1EZ/19IEWHYLL/sCCEfPxg/FUMPUkSOze9v3BfHlD3elTM56gyjbhvL
zDbrhBon5f/YOhVAZju28yZLK88modYNxXVUKH9wbgzE/ttj8dZVpIzbG+JHlfp0
K3ewyft6II3iLjwLgeXUWcoRRcMQFp5Q1w+gBN83WI5DImH+Ys8lNS9oWCTYvhnv
b+jU8DnPho30LPGClKoav9VwAFuSRI8mB9zL/aIPTF42GLoP8FemZ1+11ZLT6+Ch
5jM+H9fuIt078WUmwHJuToxloSp1CnD4rPgFX7ZPwzdtUjmHJ1t7L+ORouUZZAbq
L5lN7xqYPgjS200Un22to+ixynuQFXNYAigD17qT1cTdsUjg938ioO2I+iyNt1Zu
JP8l2fRTFuZEW7woA+kU/mOHvv2dLhaD+kM58LrXi9wHz8XXienDxL/jNi2hNFDV
jjN6jGg8zu2lcOQgFjEHVOO2sghngYukpCJ+1DvnyIjJfaUJ8rVfJJU9JF12cqxB
wKRyzhg7Ti1h7yZootFeJV38/Kh6iZdGdGJ+zCkNC/WufMd0Uqo2ZTiPVlpIkQf5
I9qiKMOIS650LpMSXY8AtA5MpCLdRqtKt0tuJjuU/51Kh3L5u58N5DzuDKwzEIrG
7DRxKtTwgFKbvPn0ic260IW2yHumCzlNLMoV0ZDiCduSHKUHNCsOgxP505tSbr/E
pRAPO1Dj9SOjliHiQEQli9G7wu3YwyHeUP6DQ5ZY8kVxTel+DuQEt0WVM6qatqIG
Wqv0c0UsB9893uCYbRkTNFn4UjGN5x9YnVgb/DE9r3rn2KuNoDcc4+7KC6mMgxPs
thbipj7WZcxqkSB+xRM4Af95zCZa4YZmck/pwljRVyKOFMtosWu7bG2Vcs675lV7
T1IsvsBau5mxf7RB/0nBRPOS/DmIySYVod46oWRFbHPq5wxJ/W7IfMvc+xD8QM+d
JSDy9JhP29feq6iVljnMwJiFkfsTagwKv9Fk/DTq55f1lt/NyTVRHSmI9+rzLpun
85TACC5bwAE/tTe0JDfdXnW32TeD33WADyn0S9PHkZGEAA/sN8bB4Pf8ms+NA1aH
r8UkLK6t0VTmQ/D14r6beFZdIocct4jNjrxO7z8iEHHKN0kj1gdDWk77CcK/9Cx1
NHPnaOO5bycr1DnOrkvDW1pCNRhLGbcs/Gx1H+6xsKfdXaUYEfVejBHgZj/YNqxI
BXEk5xEuqE29CYsA99Tazqvs9f97VBGT4hOyOATahiy49mM2CIFJ0aO48EqXXu5N
h7ONlFFRxfFk0DjTUaBE0IJQcPxPUWrCJzyu0cP3LBtpusfdgfyjwrhNqMu9TzQV
w3JYwtIzjV576WF6udfSoTTXw5nmH8KEvFZ6wLuTGbBVYZqsSLK3XL0hGHJdrQrY
P3dne1dIN6dN2bHCh2y+sRWktesNiLCr6fF1bPsmAS8q2y8NcM0Qlo5ttp+YslJY
O2O748Ev+w/z+zXC4NwlmRh0rlsfK/9vZM9i5sWVSCzjzXLlb5CL+UaWTcsrd6Mq
qKt0YmI173xTKPEDkiJOQN0CuooS8/QkcqF1TQDqQpjHW0/jkS3T5WIx70QoZ820
8O5ZJP21th6a52V4Pf2Aiku2K1VFz/HY85O6dthS4/b00TUGGcRKq/xWp3o5Gn3X
bqr1HRPvLXUpi6YjXLmNOVTdGWepCHt0EAnDbVVwrKwp+jUcWeZJLVHfWWVbn5ka
QrdUt7EAM4RvoHO5G52YZmelXqK94qAfsfKqhBc3B/tAkIW/hHrX2PstkFxZ3F23
h+4n+Y8pBCW1afVfz+PJxdqOa7X4aClxs7Az9tAJA5dDo0geSPTu/frIw0cZEM9R
dGSblLJzJEw0HTYLiDSLTQQlF0N71eqAZSqf6/27HSN4N9BBQwXue18Czdkwv0oF
s7onTBf1CjiwvcrWRi+5Oqye6sTT/G+H3IMQAlBEXTH9Ezb5C+xyxrCJ2xUcoEjF
47K4UvV/VpUf50VYj74fXordCRZ5dXI2N48b18hca3DMguogibkuMqmRg3xvABB/
sUxDJoG2yfxajVM3Q8RNcppufb9VoLHeBS68mwJxGI5NrcScz6sloHJgash52YZ7
4RzBb1lI0JyqxTZJDAwb6njpCbUf9Dumzx25X+heFdqfx/8hV40VcVuKnPzPSD6F
QS7cncoafgZDdGISFZJpt8OPQM/lpA0e4U70xZXZT2LS3Ofiv1z736u1fvJhXVbD
5dk3hUjQJJ2amMUtEP6CvA4BA81qkK2QL2O5IJUYfucJLJpl4KdQPm7fsWf+6A+5
z+rTqFt9f6od/nJQOIpnE+sf6dsQ7jzkXA3sFz4XcjxBTPvGxhmIA30Lv5InueAj
uPDomOhkVOrI0Yd4nbbsykaVXrhzaEkuHB4bUyLct0q9/+JW8cLkT7dZxuZ2VFPO
VZSWWSVgNSpbZQ+II2FYmS3xrFwiAi0eWlARmXkQQWomzlxv2YMhEJ9c6rJGEGJl
D8+1O7UUlUTujo8G2TaBCUHloPi+j7j7Z1C7YNzWjC3oZeaj+rmJo6fhxz4p8SkB
B2XP6W0y4f4OBXrhGPyJXSbbedmv7IviIRS6+10pQ6bGpk1tUrdTjDVp8rZp/AvG
TDQ1Xm15DJ3sR/Wa0XY08tvh4jaA991vV+0qBd0NRA8FzD+OM+9RPzDVWeq1rZI4
HUDXwW9gkbSOPibd2pqB2Voo6J5BeQsNcZ1YlPC4nvLTOCJTipwoeTU/eiF608r/
QZrM7iM2S+iUZH6n/cBikzTM23zs+4nH+8haKetzehgwQYwxmCa1cqCTDoGd8JRH
eLY4D/ZKWuiAnF59sauVswD46Q/Ixml9XXCwl5tf76j1Yf+zH61W4kNoKeNdLA4H
VD+BWWO6TQ1auaPofaYDNTNCyURBX+drlPSVNcHjksL5sBk7pDphCJOmry6+2EoQ
y8q703Z5959KX1vpVTwMm/KqQvD8arQQ+WKSjLY+GWLqgPnhTOJw7FtCIvNrdhoe
Gvg4fTiasWxtF6S7di+CugsWXZJp0uMvSL0hquNZPNPZPqjeZAagiEfO4WdjRM34
uvSJi7MMxM96KlRQPabzmdH/6glba2yRFhncTtJ6k8z8HDBrazqua0eGekVvu99p
wovOOvvHIMOzWvb9J8CsVn/xOZxAjx6SG2tEOKT7Ftiy4Nj4aSCbdCqbBtnRV06O
UQHJNqRO+GfVFnOeXc10pUw4wHdBpwYDYqhiQ7oGvSXTBdELE1eySaMEzG8ndFNC
Ju6F7LA4uqwF4B4b4bAx0jD/KCOKzzCmkx7H82shbRVurP4c2S+k+ag6m1mRug5s
S1Ao0oFRDBR8fz8Fawk5Ww88LeqB81pXy8EnPIR///hOxNNo+l7+/cyYiIw3pLuS
WiZER98lNc+TAPZf0LH0Q01I950LDeF46MSuf7UD+3GePUgUx+4QzbcKZlfEcrFG
MYxyoQK0uNyFODbakKaCnXFUzrSGz21KrahCHxdosrIn6lDRJmGrSyMpZSK6jUKm
15cKORLeBlT7xdu2HmPjt/+2hnhwmpfFwIW4qtAqQGD1Eng28KDvlm4sFoqVWZiy
dji59YmXIUbH+gaYE2uquQUXu48g4ri7fNZE6tr9MAR4dM74AM/PCtB2GMDyWPu/
cYKrTuhZ2T0rSNwbw33XKK0I4TZb/ISzJW/x5HeOl0jzvbJe/tKFRlbX0YubgM0Z
V4BC49GY5Kw+Wb5njufn9seTSjTuaHOwI9fuNHVaAcMI/uOcO7lM4WmAO/7B3Zzg
D45M/4gFv+xEgMfAI1/CTyAo0yTGw1t+Dq3LCHbsnFw4UYp9OpxF0RC7xS0kiBY5
y4Y1Rat7FSgZxxUlUVoxu/BVm2Jw2RyolSwfwVqbUUUbwI8n0Udk1ZrTo0of7V+m
GfqWppu0dG0XsBMxwYLwa0kUKLhnNlPGHjxEyzK9I+GC50j+cHgFA7VrCKO4Y6ad
KWnvYfX1DUavMQ3QdNOavAhOclzJSKS30I01WAi/EHzw75GpO6dzIhUR/47NxCQr
Yu8gyvsndKaMqes3FSI7YTb9/WomiPtYBLd1IhVSt4+rCsqOb2cAh8j89RGRmlpP
JI1qOvV5fkBLTOjIvAaCEmlzbA+9aCy7dze+e8hyUi3Cp7zdOtBjyfdQ1CmkStU+
JrxnQyqKHhlrlleWNOwc2zz8o21sgwuLF6+BGMDPBFmZViXs0Pv2ruFG5LsWBrgc
JAan1dsqMSbFwLqqLsGtE1PnZ5YLGD0OL2Yfc6ONk32oxbf5wmfGvDA5ZKGTl6Nj
OdAfZoFgX/huNAmdkANIc5RuN1NGU+y/jhEwhBUvpfl5/e7uW1bNZ8HAUP0ISVcD
BQDY8giv6pV98q5SDe4ZQCS5snhVIrWgNTaUUG7fZnpRnZIoXFH1IjLS4rRQor00
PwMulajUrCLyUZMMJnoKqRqEse8gZuzo0vzJ5kxsVpP2mKn0Ntysr5LpQSFSVHQl
WsYcFxIzRMToyS1fmKYLIPaycCpFjHo0LdglrEtVQNakCjcwwpeilzdS6+TW8Q3u
vguijLEFgqPGn4QoLdCIHzVVlVr9GTBnHsjNw+VDdnsmCbuTnBH3KqD4ph85q1a3
ciQbeTf37tMXu1k0zmgnzxM9mgqlQ7mfUnodMHYjcd3ggZVUYypqyMqrvKJL5aTu
MJgbn8GNt0DHHAV/LnRDyAjCt+IxVxd95QxnGUAd6YejZNtBhGyAYSSmiOtbKQo3
5zLOq/Umt8Z1aKoKY5jFOf6y78mH1Z3SaZ4BwmXJ+opKIZ3lPoEjcv9nf5lXSYs8
kFFB8XAksnRby1lRBk32IMmyuEXDGALPbUIZrEuQHByxVnheVS3bUM8XrLZYgXxv
6BIQPI6k9ZW6Bu19INf2z8/CiDNyJ2LTortRLkxt/R9FZ233e1kHNfp1XE3H3baS
DGUDnMN4C+EP+EwHNGxzJvdJ9DEzI1v5dTNBCgf9qsUMffXzBWUwSd9U2bnaFUeE
jPfwcfpwkYpIkfydWHsp8ACbulTv0loAf7TuE7L4cPNgPczetv62roePaJIdTIT6
D8SFn/sExcUzoBgYaO5PNPac26hvZia7FExKP7VUyXXEeqB7KtwyJsrxcswMI2Ca
iURdyXKCmVQ/l7HYcjq9fHuLeokXYTxSNfqomv3lOc4yK4ybJqXzyT9vFvUWE6BA
LdNOiBZf9ypACLXO/xQJbi9PAiLuqdQTtsQaIGY4avB1HyRpyI6xqJnXJfyLwuAb
lLD49kB39uTA77Fohc7JMDfl8FqjL9W2mdRmAchwx4/6IWTyIc5QWtuns8Cz711n
da/bAHRaQO2lvYP+AhDRKbkH7JCe3LpmsUsmU/a4lPnkr/7FrgISrTRY2svR+lEQ
nDoNkdlglIFKlI0uVAwUssAq+o7wfF7s2DP/i/krwwMll06J3qfgW4ZHUk/66ER+
OfVpgyTIhmYLr/y4lQspYniGq6steIWiTJWDGeFLd8uoSMoFtnKquMNncoZTl14q
ltrUt+30T/1aBEoRBft9lHV+3KdlIX/tksu/pHBRIZ2Xz2mNvwyK8t9L9P7irfOW
hnmp54eEo9dkxykvNFTauu8zbJue8Brz1YPwzaiIcdsD9pqGFsWj7CN+Kv5wqH+W
LnBKVFR9aV50S7H8z+3b3wQ7O30C6SdbUIo83anSgmuiZd0sEvx4XWURtSAhDpKU
ikCnfsfs+r/p1CTRG+q2iprHj3htu0n6Nit0xG4hr+dKYBAPLsi5zcz1/aGddb+W
3iXn6LwLx3RloPv62EAPUhkYs2YPn7M1tuKyavPM6NBf4ocb0J1R2K2oag5zFkk7
ty60BJLU0G1/KhcsTONVsv3l7Ek25V1b4XUwEkWrrn1Lg4gIiF0vPi4u6X6H1ibo
2xaj915gA8A5xhBucKKyORr6cMRPYX8y9cnXABCyqm6eVIDRfGb2tTwdgXrKvtsZ
RmzB1oFg8B7gACZZ9ZWWBAvbZU23/rPmTSBFlCtBKtp3vQWaJMeQpd7VF6BIyDBQ
daj4dY4PB/6t8hH7apkkpRuVvMHHsNP8bdLgfI38IPhf7A90Ex6Z+Tc6VRFKmlJs
TGANP+0/NbVW0CvANoEoJMhWz7ebdqaXC3rpKJPaytqStV/jr7NpceIgo54YpxqZ
MIBORXTb9bzQG3hK7aXHdj6q3jNAf9eSKoTooK9OYr4JN6bM6XZPpIvzeGY527wW
aRbyU/HgmULS+5Y9vI86lQ1qEBk/SI7UsdUdg+4eyB9yLNWdeHEgD9vEz9dYCgRd
5FpzHGlzp5pHw6qdsAESu3B2ntcOZH3+cC+gKCp41IjVr2+Ce2/zDwwmqHrBDJoB
sJxVJJeH5Km79kI02PH/9y2Zy0UROYx//1K3RD5VIGbut8yLmLxXOOMVQ+eQs8t8
dmTpgr+DgI1eu/CxcWpK9a9FrsUDuz0kT+uFdiwOVPx7VG3xQ/NFrNP2unjkADqQ
fYf3psGHvScmgRImHJqGgGIieRbz1avo0MlzYDAZg8NdQu2Z1x7C/F6wRuAYvhKb
ofpG0lyuKtOieazjt+6QdZ7WJVXrXl9usGQhl1LkpX8IQ4IMpwCgiTOtKA8YOnjc
FoFlSnxYpxHie2hDUMccYtIrCP1Od4UKdyHULLuO9mf2rNMmB15JJ3HvXtrpkeRN
EJ3BQdMxPFj76HezrrPm/pjVj2gI1vMTL7+lxBDeQzhTw/zx2+5Zxz7zVSV2DFqY
rMV4nR2vl+ei3lgOD8Nh1BY3/Sa0xUoMIMQaOLrUMVze2pvBWBShB1BIuLQ/RYDj
YJXbuBp5e3GTfpdmNO3pCiFnvy4yp6vE4ycAZA/uY6/yJkuApGK4YO5KqxIrr0K/
UAQiQe40FEW5rGwZ5hQpuIwNhjVc1CodnVndUXDsmlrVc1Ek4RgaHp3q+SQqYBxT
k1DVgj7vwpoaEKS68dzfl7l/H/G23VL3qZD/4lyGRNnXa81q7Cak/NJRBgln3eQB
RufoCdb4iEw6sGsN4Iaex1yNLHLcbejLDI9Ck/P9WaKwO6SDG2d0/QhbjqMqBzwm
0feqideIVa3Uv6vbGs4GT2+eIlsN5im/nvI2rjcU1EN4XReySBPxAfo41sPHnpz3
4K75vpbxhAvRIMS2neQ2Z6HHc3LYS02exac2VjU8FAkER4Zi0G9cMHc35V7D+Qip
dgv3ks+3bbF/iX+lw6KF5qb7+bd1Ck/SqxWD2x4A5tnbU9QjbgbzgmIRVnYSgxsa
ZMsVuKnC6ao7Ot1WzogipRCEdkBlWgrE8Jz3IzNCALuu3lLgaoyLrN9KKqyggs63
ltI4lCmil+CB+UblPPn0tyQNFrV62WzOZN+c6XLBSCHtE0NlvKzvecBGxrkeAZWu
j/mwmhn9rVikdKSaCOFjVogPjUVe6UgrXE2kU7IBnKZXr86EZugfuycdheVu6RsE
KzBQ8Bz6OIuQ65PTzDjMvdL3v8oG3MeBa7Ws1JSmEwWJ16QW+SvXzAg5hYnEB6BM
cP6eG6q0y9bopNWPIv9SDyUw/vwE9ycsQfTfzhoDENypkGcIhDsqM/U2nuZ9nzWP
lLgxZWWrbGz3Hnn8RxLwubsUABMVkOyAOSuN49fV4/ZL6h7ZEjixnHbOaqd4+wEu
xcDNtxanTkVrEvsJC7lkGaSsw9HQ3rF+sLr1BhSY0p426cxPe+qv8ph2nbIRftJ3
eGmVZOTjhWJWBGEARDAODi/w1sulh74q4/d8RvEaEsR9uumWV8+RglMkiU+nIP1Z
tOoicCtdMFe9ef0Kl0OtDbWsHzl+m/oA2vAKi0PNibHjfyz+Y2VfByyPunTa6o4e
0LQKhoApENhAmBuy2aPGQ0N2Sj4FHEo8d9CpXX3Yu2yIFGceeKMeVA2kG+VN6KIU
4TbxyNcEcm9xW/tOCohKNRzFQ88QVAvVj2J5208wMIouhX5FSPC2NxvgDq3WJh17
uGi1B/qs55Af6J81aV84+MDR4KZBMKitFvtGHxyBDixhrr38kGhyI4SqAcP2ef7d
GI2tSFeNL3HTRdi9wl7rnF7km57KMdba7fvpGMpHciTrpqhpLnRn6/WZ9mOO16qb
fwuVlMVX0s/i1FyM9zvyxo/MoKGYTV+3Qsubz3ompBOxRROf48FRVnWly2UMcOcB
DtIdLT6J/3DUxQ/bBIZ82tHmPiDVAUkxRPM7BYPwuxRHts0VNMhHDKaigTAJkEt4
9rBdScNVGIRO+JigRqFidfmZaLkX5ZHVAvJSJnTbMASr7hhFWqS1fqydexLQR1ag
63NkYn2nKGNf+ElCngl4CaoaH7sWc8Q97ferFhRxXGmS1S/Td4eXoyPTGPOi8tQN
EylwmR0oUxhBDNaHKjgxPbOzjGLm41vXBFOnIkiLn/Xoplol/yCBRoURsIK29Njy
/dGIy0j6gJbvpPmax0ec3YkMt3SrApulw7V3XX5rjwQ4/v2PTN+8jHlrwRHNc81t
U+2SJj6TYl80uwV8A6JXmtmwJXZOzSk6U94ynZpqSnzDVK+GApwOb7ReDMHUT63A
uqrHAB+J/ryeho8m5SN99MG2tBtavRGQY4JmnLfiouLYdQwKNq5W1gvsuTft4EZ8
bVJ4IHGRkmz4/dcKNlMHn+rAQMlU55M+hhu/nHO3fWukVxorOy1s7xYp8506NiPR
tEbZkwWTN2++CInV3i6o+ae4ZLN3/HRifR/NNvzkal6MW1G11KEVZbHwa1FRztys
w6pyliKGiMpHlcwrnmB8n3pyAfYhBKRTDjE/ZWigTOWwzosnoWd8mKqvn6znoCyO
FA8EDyEKF22fPBjBsewCnKAy5cGIzhVLhrN8KX15XITUayIHuip+CPD3MgTMpPAu
yqM1/SZcICaRUR2Eino+tezoXQ13YcI4Baxx/JtlsPkZuHIMYz9qy28mIlwKQzjA
WcmZm3YwFGp3cio6uZ2GUJcBR1yffQlbZm482ct92oOcc5ubFHXZkNcZAtjvZtdC
b6YcTesHOycmiTKcWMFvfEt9MOPJSoxXbmcKjioEi4MSF4FvLpnW7dSal+Z0o8cm
iB89I8X8ZXJZQQHUwgHcPW7u7d6fX7GQu5Fuzf+vTXS04poTdrNz2TUXmoxtyh2a
wA9n4tWCRKEiExTMYbeC/z9x2+5EI9atqLWgeLANv1c6qvXEbLLZqgqpYKPXNXtn
vDHvTzQfdwMprd2npQnYqC7W5QpwGwG25APJBg3/hx7QshYobLZOa0jydbcS9Fu1
mM14gGZhNxn3P7tyB0gJbLuMoSyhnbi5ICXz79B5fRh7o3+7Xs5E2G4QIkZ+frRb
1+mwcw6pYArGL4E3WPjaTYt6E/Fe6cwdzyuAvllpkH7Q6vJAd4JOlcHEHX0luZVe
hfnu9PdC0ZmoDZUQ1jHfLt8MLP/WGOI3k814EQSmFJNGhlAxtg49Coc1xmo9BeH3
bppkwzvr1HF9DO9QwzzlnAQOu5ie1u8lZABtlKSrCA09DVqWLz0V7OSqkfK/Dwo0
dayzw2FYmBhXqnHV4veI0nJZ8NBffERMzyA2n7CIXjaN3Vhk3mupg8Fru3sRtD/T
RBTmt2XlYc6wQkrT1hoAwpoRZbFZeYISMuBdspXeuWtXE/CvMfyyd5J706DDmEGP
uW1nD6zJKCJSPmiTNR4/2zP2eClA5e2dnVQod0jPn/2k2flCusQZqiHVCVA5/Tyo
f3nBVyYdeB0MariU5adXq5wK9DBS2/H35XlFuw5xAH+jGDYPXVlvGzjXRsYNtBcP
jZV7lJ0ZPyYD/hCuxdK9MqWXwh0/P4uCpS99GIaxQhXmXBuTJOySP9XBLFls1Ldx
sjPdwLAr4a0z2/4LIB3PUZmtQWUBya2X3GeOzHuJPX0VmDjWwkWHbvGdLX3UvCKs
hYkylC922EcIWdNjdrjej2pqASsCZ6Rea+RQQXKB4H8P88ZUBOIlDUpBznaDnYRS
Lu+fp8bsqaTJ1Gy8LPqyBUswYRPruind7os16P1RSA4LSqpawIGY/H/7Nz0rWNp9
FVbwKHWgfFZ/j3p3Cq42KgSoArZidVaSJWZ7OuDqpXCiPufLqd4iehQi3//Xt60L
iTkpTgIQPNmlONRZzdx2dx1OTK1MCroFmCYDbNM01RC4h+SQl8hMEamCN/BMmqWm
LZFZhMdC30qRvIVE1/+XHat15YRLRTM53AmtATz1XXWdDB9rNF2OkHW1AZOYIbaG
moF5uwrPOovoHqTCTfo62Fdj5ib3lOEtofWUw3W5IVnS8UNS2kmwGCdykifODQ0u
W84EVLZddUhtAx6joBpZlPbvmaYMFa13hlc1ygytCLWmw/NeUnoC1ZJ7+F8TX7Kd
vyNdKY3+k3TNvT7R4Cvz8R0VETioJdDpbG1xG7VeEkK9KKxQLDFsKnsV4GlvGMI3
c7YJ9lUSFJCmfxxgMstHGvnzPkfolGdrOe3Ne1Sk11Na61lBMChVCkgMNv7+Uf5P
fFLqz+8z5F0OlFy5bMSucTNmaulfjoyWa+3KIPsxNOE1qvMZPhR3nJdWmDOesS4/
ppPOQDggdPC/3+NfrQS+IljUql6mVfpBzrrhr5NPt6kMNW+Nv6TLq0UP+r6GS3+w
Ng89wbZzNSJAmNPM7HHIFxKll1G6ex9ImklKg/ml6yJVUnAmN2NGJaBWXIEM+LOE
+aJljezeQtueq+fdrivmN3a4ST/1RYwIv0AtDmBggIb4yGytMntsDo88LA0D3JTJ
iMrXFNFsrAhLAhlNZXJT/0bHGmPKLC7rP699YTuKbYTyrSrgmTGOA9uGwCuOB22w
IFQG4BL2JSb1wV01AFrGW99jw2VS7ZEJS4ZV+MYpEzBzRRCDPr7fCTnLsnqmF9ug
m1jphcWABrkDtiHHwLC88TVebDR0y6+IX0zQLf1eGyVenBSXoIMAGVE8xjiIcNOJ
xd1mZbQQJb3RTcQ1zSM7V1UZPZmMdgagHfrG0Tzr028MgBigjawjrM450xkjeZKC
nEgC/KQkK8wnUNkGuEWj24A+CncWSoYgUWtLA9DuF1t0tInffrIYD+FS8wljBv6A
k9F3ELQYvvpfWP9wJVszzGBhrpNkZy9qd7E7DgTQAwLcOhLJq69FnUBDlSmJhMED
h6AX56Yap8vL66CO5a2pC4bnkzkmrscooJhxrMFcMWP0XE7XHXmqvO38i4QlCwwJ
bmDNktd4sKjnOwXGEVdXdCErDQ3LI1g5h0UfsItrMdZIMFlPx7FC8p+KROhMxaq8
gd0jFP38lIU5CyMwJk1MF6C1CjM9692Oqxr8vMhC6GZCAgQQf+L89biuBiVCcv55
VRL/HVVBIcAoUaT30cZI7t/8fZcn6yWecX+nkpqljOF/kET7vDzYg42cO9iK/loz
TSKDAAFiHLGVhOI89axtRgBoLgPYrgyXuPwL8n6z4cZkuRgIAAWQtVFpS1AHDM4j
dS83zuCjo9NNvJoHX9ThNg5DqQatqPrMcL3tP+0d7JW2wzDvnme1xAjxEPNX3o4c
DUEn5vSd7oXDX76nlUtoWCqvb3N8lxJUvIFyzUQ0VIcFnqtwvEweo8daJhJNxu9H
C6rQYwfs5SPrHWFFlAuHPi2I95cSj8XAfO/L6m5+C6XI1435DMokdQNHe1REliT6
r2/y/5wsFu1PkbsIXSfwYUpOityE9YSq4fx+Lc0Wh1+syykDTcP/9VGNBnHsvKda
7cYl8ToCaZiBOMfEyySTtt8TiFuL2Utc95bDvy6Nqe2qXq4/H0nGb2K8N3W859Me
Xi1eV+ov3WVVrVnNovsNkRt6AKXN8826SWResk48+Ku1+x477x0wg4bRKD8ts9hl
PwhblEnDTVVs+kAXOP8oO1pyW5i1WM5SUDwvaSmJbtJz1xs2jlD7pr48EZWChGjl
CxHnghwxo9EF4P/Rq2OOgDtxzDxGraBcgtWvIu+UaxIdHnryVVpNu0Pk8xY6S9G6
Vu/3pvGv0DGG6XWauIK9XGbFrkZlns9NlUeCW0OLgPsYDOY/Suv9CKPtQxzR201b
jUdyBeJ7GW/UOErIrVLu5W67iHKhSRPUR3Jbj+vvakdO/9ivjdRdLTueBQh1lndO
cM3jNwNOIxs97abJT3HIdZkvdc3mvquBNL26DFu36/CpvFwyxlWurUXmNX9+Usvg
d/m+ie9FiMSbgSt27PIapUgvMB4CSzQ8TRL3sU9mYqPvALDduvX2PCmp4dsOYn7k
yRop64lN/N8+PAvEf0nIrEhdA+cjnumhwLiX7j9orVWkdbhZcHWcsZq2YveVbkdR
e4BiAx4WkPPHymUwCEpWlfFmjVeeTV9FzBT0OtNB3qMv+jrd0XJM9NpGGnLd3luq
VpJ5l4EeJ6KoObJ86QDg3ipHKd4atpH8ZJhwQW/9LDoYURx55xBS7hC7fQvduWHi
5Slj/5xKbWuCzEUHTODh1WZC39vP0ak7GFT7cVuYPcwHxMvCp10Am3xKFTMW7Lx1
2tjjobKmDN/EvmWccFDxgCUj5n5DP34MmHC5tKRnHZ/S98AkJyqjzRdKZ06feBns
7vxM/X1K3xoXoquWcfTAFrPKeL3zKGzZEj5K8nvTVw/KOz8IXlF93xEjw8OexHI2
IKeqQoc1hJAcU37f0szhaqXbFhRZh6qIohqjLi4qtCylIx2RhjaMNeUY5cg+0Mut
r+cjLgIdr9Fjpb6yVHfSBIiVrzZMUMovTdOpkUivDwNejAbGTjawkHEzN34SYwPz
EEW+kJ4a4TaPEm2kFALzCldI7vlrT9qyPu5vubEmKTslhO9OoDfcqruvTWnM8x0F
sgXSV1SeKl9y1WRjE9Ji2/p5R2ZllXVB1YrojgYQrfqsSuMksaC1eKBZn2FSH2XR
/NM6SA7S/cmOPgDyBXQk+jmLIj58kKc7Nz4Fjg0ng1PXORNOt9nRMBu0URmbwLYv
jeLmIY90AB7eRy54w9Go38Cfq/c6uzxWaEdL2Vm249dXfLkWPuru3diQWXIhcACl
8rRnwh9nW2tX8uyxiU5lysGNfCqri6LLYyJTvEZjHDhaSsPDuEvqRW4Fe+Qwpr9N
NRdVzF8Nwt9bfyUrafek2WrSNC7vOLTavuPOPnx5xKXCb08/SbYfjtuiV3EMCgt4
Y6G2dK/Qonqxfct2TbDNculj2Y6B41fqRwLU7rledDwZse0+gv9eQjT5e+F5Z+yr
Rn8iNiIXuvduTTdljgQlmXvBRU2onZLRNEhwxvTYG5zghz9aV/3h3jUPHAzI4hMn
mihUPsCtjPaghZLKnRUiZiQDtaFejuimMLbDfZbcpAMEgw7dy0wTtzHoeH1XimZs
ZW4A51/ci514AyDPydPPypURpI9rCFJXlM285pixpbhjIrdurrLMPpwLtBrwbapp
Zrf8pcZ6XbW/ZQa14TnGul10rjekVlw36RrLqsa+wmKHrnALuk/2LyZZxuyJdYJL
8E2i3cAirJBkgDhONQWRgzrU9R/rID+6ovier4N2pJMmNoDNn4iCrFEtgq7hr7k1
dCsLFM1FOGuOlPcjLDsUgVQkjN7iFhGKGlcJzVeazSbEIfwq7dd6E3jhQhFcY48i
hS1iY5KCsUTBUOPB4HmWj1axXiBLdXhSxDSTA5qfN5WBCbXEcK4Nywbxk5thbLaD
mGm5gNl6sHrZGIKDQd2afIqgpErfm3ptGFufXfhiQiW+5DOTDcm+tWj4G37kjwQU
Wj1EL2YaikBqoiPoDZ4avzGO7rQeZfXI/SsdL6BvNpaMFExlmwmBPGOJn0FV9oVb
kz3j7j6iFPk15acS4KmPqB6pF9Pqv1Z5C+A8kYY/Nhksm45ULciNLHwr6TTwbpM8
AizOteRw+/3ejADVIvcF/TQy9REAWuxwT5CIHF3qEpv6HNarbcqy+4/IYOwXMkbW
Sy6GvPD+AFrwGyfEpqSP+XbkhOi1MMWLPtL7MnyKeItmK4U9m8SOebwn2V4aFWD1
6S5uXyOrrAGxFs+CDCW4a/iZTcXVN4dcOkj9oTpR/2rTjaooyeHAYE7IQ4hiRTPS
CYqwEVtS5N86h8KAODREpHb99p/5tYI8QQZXyI9kGfZLEbwa51LPERatRSRL4odp
vtEthLNcCY0RFQjj2QFvxhdbVUNlb+xqcQePF54bQibQjp7aSqMW7639vuQU8mZQ
PVx3Dqydar0BsYuW3cfEp//OM7QVwlMyx1JDNeQredK/6/4EUdkK+vLxAX0Su9kM
/3eORaGAdTp/Z0r5/UOaIxc9DKVCzd/utxODdDE+SRPDAa92m5GdSiWTKecob8HL
J4l39iJ0MZWEZdbXZuQIfJkemiURLgftAzufAkK6IkS5j5zWodVqCA8wdtxBn8Kc
DowYvF1U1AsZpapuKxzhVhNu5ufCwGVL4i7kmfHBgznXcuPNkPKluZmNse3NkED2
8h6bpsj8bgqubHpZ7oRFx+VPxR4FZdFsKnVljiK4DT5BzHFTZFYVl0/gQM9VlAEF
Uq2aOc6D5Slotc0HYMMtuob6P/7jR+wCx3R7ZTbQHYt0n0uL81lHDwfyMdGFLSqU
AemGAlWfln4SVX1DOLowRq5K1KdQPLmFtP8N100Z6LfOYXIsmPK8GJFERH7q/xij
watKkyaeiFNOA8fcPkoWqMKZNXKl7EJCFNKBxixd3dQDZZuM44mzryAwLZQTSBYh
noNN17B2DSiWSE/HxktEdj/sBf1aVBr5GRfUI4O0NYfHmUcjKa6DRQHypDu8o8Y9
Vc2Uh2HS82agYbPyCp0BGlmGlm9JIMFWOLNLS5b32JY82vhfuHDpIL0yTpccjaUr
FhUtqFj2InMpVyGvw/tt2IdIKk1FNXwUAjCe7nTsi4uhm9OjgmeMVroZcARahxWf
aFx7WzfTwdme5zMCTSFeQVGcA9caCR+pMKkbtQ7de/ly6IWi18CW28Gt0QJla2qI
DI4wRpSVjRRA3m7xPuVIPE4tVotXCTcE/theLngdcMV94cPpoQuOi5GC0rdgFqfl
1jMwWFolq9ZzQNUDYLCPe+glmS0NQnhpSAsN3Cq9U+l+UpudgttiBZa7aS7e1SgO
890OhPhbb+Mn+4rAjTyG4Z4vzG+SSDwST5DY4+5b2FOVBHbbo+CifQBtsw6ROYnF
eFf15LQRjfEIAtxk3LDs2j/MO6J86tDNtIrneF5DSOnDXC1pRNIXZDfu9c/tmBYL
c4hglKGlPTmJ/JvRH8IvqzmVHEdg8wNNhb22Tn8n2gD3zq9zwP+GE878GEid+D1T
n96by7Aaw0Od8dLkKEUXWeslPDJ61ucsZ8uqPPJKTSt9LiwrdXeD2TMQPd8OpLmQ
rwKwO0pa8b+iULskIQdYmt4hct5s7YXvPj4xDDx749XsG0IyLQdna99JEGYTFJhB
5ZN9ci1cdNhcJApJl1DBoGACGjfweiFKoULLVDkWKbywyMPiPhQEEeLBhqT2Xely
BHRpG6eCRwGyWX5ZtDI7fmrFvsX2P9EDVW08YP3I/GOl9+ns+/8xCyubxBFveXbp
UyyiSd+qWEAL50yAQUMz7WbBdPjb0pmqYyRmd/9XCwgePZ+K1Cjplv5w3Ji147s6
t70lmK7f/vJDYjPxzLuPY1NrWX9IeT7hW81N9qEIolDeIYH/7mX/UkbV+zPO6OO5
DLQoawoNXeu6iKHvQU9U4kXigXzes2f0ForeMbGpzGk+Gm7Ll0elm7BrS/IlYcIe
NetK63VuY0k6n96TN70+DBKuRfgvWeS8XzHDskq6kaD8lLy9gMr91wZR10Rgued1
6KxepuXqPkNKxfHTO/lIhdNecIAmeMCg8spU+vjjdNP/TVO4PAIIcY1aASPDhLlT
xEzAzDjgEAZnp1twyadmGxc16K0kQUo3PvwBuZkJFQkeCu6WGUZ8R/O/Q2w//gvU
yUhaut3fi9AO7/3UOZQH2k7dhzyDBGc35wNPe8LgcIxqTHLywJtgwprHN0l2Ii8j
Ob86jJ8BWozJoFAjpPWALhX4pbGlcZWh35PYqwkm37ScA94wm4SrV+dTAWWxDeOR
1I9LQA1+0RZCLfjH9UBX3zTdfmiqsPiwH2rrTtZTWI7lAz+tns3fadV6ON7w6+E2
gzYGWJGRQzVvDQYK16W+UveFGZ7WCSnQGNiXF9tiY/eu6smMDmt6WrxaOWKQKP7O
bRKDsklhD4wXgrTfES9L45FQeQ7s8C3Yg9QK1i0OXIr35N6+8hRBTWBP5tj97WfK
Wb/5ht/+48V97lXx61Ite1q6OaIwIaDDo/Tow30djCWhDyFcFJ8T4yBnqscVoIxY
oqr2lntURLRXLlDby2YpsQ5vOnnbzDeSHSU9Ii/pDSbPTXlCJepol4IXPgKQ1q1s
7zGPyVs1lIlBMF0HoCFczZCThuDK9mgY9U0wfJXy6Ew/0vug+TZW8i58XctG5bqf
H9B+6xVhqSVrN4OTLlXrLu0JCiPg2xDijqJNxnCDtSloPrUN0DV9cfo0l6GA4H6l
IMp6fAcVMOglQioDeyAs/9+W1syhIQP+g5M8uKYzMecszqzV64flhnPElQREOx+v
4yz+n7/3MFUhvCJuej7trljxqYPHyuC9Tk2FkT1gKASLO+TtJT+RtzdXmvK1qDka
qZM8fHizl3REsJcmIt6/w1NBkzGzmyW8mX6EoUpKP0Gw38hVJFAbm8nSvbH6Ql8p
okg15dxxNVFWV/E6BuPfFEInAFsqNOvMdnS5iGhIHF8jh/t0/xezV24Ads4sgeJj
81SD61aE6WKKKYqCHprlEIvBsyWbwM6RxvD54MzKfT+7XVh3u9WnvhuJuWBrkrpl
h+a9SuPZdBVhs80DAx/5iodL3TThPKRMwpc/QMf/Y5vlusPA4n9K8GWUkk+pPCoL
/UX2MCEY7jWHXSrD6gEHJn6z5I7bEQCojh3uvaacFBDRJUqonJbN5g2P1s0Ntmky
UUHIHZcLsCMBJcRU4QNmDLh+n5WOeHJyJGYUVRdJJvT7LHvGbddG/owOTamUxX+S
vBLdiv3UEX+TGohuTkR72Xykg7evoOQarrsDrTRxM5W9bz4CxDlPFbbzR1JnhihI
y4dWtY5RvPVyRMmhf7iQyvKZRSH1sWX29+qDZzo1aHUD7eOp4jgJSahqLFfvbIqv
bGX2UQ0b3xV+fcbY+oCtMF5nHNN0XeVA+CTERe0kUimJzvXHeECUl0mxgGh1I/m8
H2LeyG2ELSIc7yWf6cdPSI8aB7sprDqUY/10HmwnLHz/BOzwu6rnxCWfOyZqcF23
YaN/jkBnoObLGwQM6KZno9fqZ3LqxqDnxR+xVVeyUvXwNvZhjaxrtRAeVYpCfdD8
sk2JDZOwpIRRSHqf8OBp5KUTCuHsXJLCmBrdKGphAhWPKjyWeI0j0FqErrHIA5g4
5+e2GQBRij7zty44bnSJO4MJw8WOCajshoDN+dNIWfNYr5LigTay2Xk67NzHb4uA
QghtGqjDCsgLzfYiSmRyKg4pT9SaGhrydeo1PeU3M5uiyC0ylhzG6EcSRyRttWJc
HaiuHcTCbC37b7hjkbMBs0th4Zow+a0+3XJmoT4m1OOBzrfxF5RV7WNagt04y7Oe
zyTFrLrwbKPHLfWqZMKHt28yytxJPE0Zy93t7gYvdcyIQ8BA+IVZ+p0/ilu0izaP
WVaWs6ufF5IcVGP6TPA+n7gWuRZpw4chDOi4niP7oANfKf7o0xpTIug+nFIvrc59
TZa7Pj10gk+pP9sDpAuvPg/khSGM1nwhxnaWgiBndoQLKn70+RTf9e7Ok6d0+j7J
pMtBo0yHv9XvePSIHEKvndvTImiPL7tl81tb5qPofi56YR5HwMe2Zk7aJOmfeS1u
1Mgeysk6o3lh7V+HUQd8SaLkIOmsMACies5jWw6chpBbQGetdzNaHbWHWUbZyFkx
KUxWppKQHN2nFQAOtkd/3bpJglvQfHKLVtH0KGqEAf+3zce5SdAzv0Bnk3jqFica
gSHAqblYKrioPp/N+8v0xTCV0me62TqNBT6X6mRuqwuZ0kBRonzJmfhY5JYBJqRH
wPDXEr4QNTURjITWfbBWzQLToxcwZKCHbwnHjBlBAnMq3t9pp1dscUeD+uTPCQNa
46RJbFdBWp3WzmoG+Z3KYIBCINitHW+1DQgOUYxWOn7hz6k+N3U8mz7Xn3Mb+XTb
kwzpAkTTSH7zd4kI+RKSNVZxR+4cWfaahEFg9ZrEhwqpw48Mb8BCb1ymtPa4GuLg
JgYJ03ikmMhlF3okhitjxpRHnc2U45UWBx98uty5PygTeN1PNwFHyp0RZltCFEQ9
hg9Z6SiaGWKpeoTxqgdGQM842lF4GUoRKuJv8c1CESCdxcfkdVbvZHC1BrOLzAOQ
GmlHgebhyXyxjeChoUi4y/yiefJdo43HafxdI48kNhuDvTGVRXRnL7DO93jx8T6R
VzS1LXSFTOEMz1JamEwVOFxSGtWztFPXGjP40J64a7wSP8hK6lgOdrmG0b9AMUp4
sAt14x6DnDMQImHkZz88UJcy0qXLyrCj4wVtbklhqmBD8QrDwia21QmyWWSXU6o1
Z1AJaRNkAdj7lqeH38Iki1NC8J2r+aB+yV2SKMA7Ms+p7tASVp6eXPGKHPEeXmpe
FV9CUpkLToahaLFnMIqpuepmOySuf5xfqTwiwjUvAJRaU3ZEPa+9KtkDVNQSlRX1
c4DLBLcXq2RXlQLlA1AYEc5XPdP8DlMJ2nn/1o7kh7sex8YlUKXyTJcgMBrdgOFF
87nUeGVFD0ROX1n5f8y4ScYG4qAA3PIuvD8NebyACXpwSTRhfTKrOssBdEG+zVre
SSKU0suIxC8+2vAN6WJXG3UvmkNvPY8dFFxI6Uow4vL3o1tye0qjMRYW2xSNPek1
1haKLdrcqpO2i4PoW/ZE1LOVVrsTq+Ja7WL+KRtIYYMbiDyCL44F/Op0X+ds6Ckb
4L2gUYxBOqfImMmQfVi5X2Uq6wj4oxVZHPd7ynkVKPDSI0SJTmC9TNiX1SbbUYJ0
GJeKoGmi2dVXLJG0phFOy5VZLc9HlX2REOHHi/ZlW1gJBbKxYVzjiVUyPZSUh7eM
zJC4sKrk8IWPL+AYGdLoL43NaqycLDbnWN3lTzCXm4pBlZ+/m91lzD5D3JrEvNPO
bOJRjNmKvs97EOiJ4Kyem+o8TOIES880CarpAGwOglDVTpIm3SSrqtfWvfPv+KSo
Aa0qbP+Ysfv/m+kD1OhMawlY9ZikeXdMrn+fpuxo7mbUbxvfpBV9KONH2YxietaP
azpVNjBkpY9tgr//fa9DpiILJC+L5CzRA216TQ0U8ajAEJtKKaky3UF/1SQiWPTQ
oNgu6KuqDequ3WwtKfmWg8daKrcVZ2LKX8p6P5/69Ie0nB5vPRfy3u0KNttWC7gp
747YBj1AStMhq0lqCAmNdjNYeaxmhyUggCkvHodZeBiP9B0yuRwY3fCFDkSFX2RG
zTzKFSMjsd6vC20u/DC9POecTqZxJi02MA1vc8+w+gbffqpugxQ8yHXs8NLHTV78
HQNZL87NKoM310P6xX199eQg08j7tiuyzWoHqntdaXfUj9T948Pd2gldauZsiwMk
rLpchr//VilnQ2zHplhOkiLxXNCG8ij8gCCzpWN6BlLlRZAhgdCVV2lLo0RVQYK3
TBUv2lUXnWdF2w5lC+LdguugMjnLT6FPifD2MpRNOKrPyHQD7+DJWugVZ4U5MdEn
M6bP8BNpQ7CmGt4odhxoxrzmwvVYEumlzEhri6J6OiDr5leDlN2ZO7HEfGyRtxWT
guoGGucczP7BgtP4GGaXIv3BHf1JTz36pdJtNGN7qrBk5HVWN0A2/koD9St37hof
xM/kkkAl8QcVhMZoestpsx2/loEuDyPia5QmWPxF/pAtlG1SoEsQV6bYIXaHyst9
Ts4isjS1tNuvsj8tsKYlv9UsgtmvP6M7KzY1iy67BGcsY1oRY+IefJyP5pK0OJIx
pQdBHbvf0webJR8yKOdsEN8VLK0blB1Bu/vL3hVD5Xl6etY15LkezmFMCqZoSNWb
WZuG2YqRbQfbh54bYDckdyklcDnLHTEl3Y2p7sdVyaNstoBkvcghgZvMflEgvedL
jSGFJyVegXKDMr+oI0v2FVAcNOXp3nAHXuHA75waNubxGHfetic1mYh4RaS3chEa
jsl8sdn7LE6hRwYO98+aqKl37y3zvwq3RhdEG3wahX7iGysXzrx7ibgRsIfBqOfF
kZl8X5Y6nauZPkZNrGDM2Q3wb7eLt9Y4PSBjQvqLASIcVL04N27LojreH1EPNxgp
9ZpFJlBzI4QAxJmt8Nquw0V1jRpGhsiNUjOuOJiVkhXbKdvs0IsrrRGKEUx1jg06
i8c3YoAssS/5rHzskQx6x4FkOrKMNAtIzew/oyHcKXaxzpKfUvtt7BJYMYZhuNU3
jy8v6aF1Un5gSl1cf4wDZZPDNPDL9QUBym8ZStd564wtC5h7G21x7VOPthdfv66I
UDTRxjnsX8FoUcEnLhqbnZ0qCqzgcPUXiGXdyp5hAPgMq1yxOn43J/rmRaUuh6J+
qDIrs+pdgOD7cUjCzK788O0R4ODuovM1NTBx80uEQwKut2zwtPQ8SrADO/8LYL9S
HXq9jjanX9JcEHjD8kmIQQx6/K5yskrFtINzdsrckxC52YaJ1fETC/Mhq5G4E7Bh
MMhxza9d+6iwRsv52GyHSxsmzWUcqr6WcgTMqIWSpbxWlSAJokC7/NdUH4C52xQ4
8tlkx8XL+auw5k043vZfc5TAWpqcxmmbKfgFL4Pix9p4GLPo3sQmd7P1iZw2bsSJ
rfSZEPdKNU/d/CJ1ULDchfIRM4hFpcwxmBL9l6rhlzAqB0NYend0QMp2CiALzV0X
b3UchZZLrERGfTMCg5lyZR4l7Jm+0e+pa7fxeKe7bY35P9PWYlFUimoKK6YijD0P
s1f/YGqoh8+ioYn9OK92Nj3LCO2CHiVMpoUum/fw+BrsIXD2cM/Wf0b3/5NerjyC
bVnL5ZJNcrSjhLgGkifDCzXBUE7yr36nqS4t2EF9+ubucmKoYxJprkfzjKrYHktx
Fye4FdF0p/xYbVxL8ujMwXA4pzwju6BUpzKKNBpdrZy8KAmf0JICDbshw9SEBPTq
VLvjg1pfjUXsULiqTHsWWz9uJie+O5IM9gpggi+GniDkpMG0R+Fy+fcVwo2JCozU
aX1Z/BSmfV6SvA3uvHVnT6PK03e29rswNKRnvg/CAAWejZmx0EZ2Wv3mvjJco0Us
76KUlA+saP24cYKinD6lMCuKM4EuilYR9J/q2Q9qg+Ihqr2OWXMU6HyorWCMTGtE
Vdwdh0Qd2iAozEiJSU655sUldrRZyo+ZCB/uX5u/4P81HUesxvD1Dp3N7vT59j8x
HR+cPJpuBAF2EucdgQXyjAx00YcCe8FbuL3rOOo/cpLCr5+9QFG1K8ogjSlBqqzV
lEkwA6f+tFzaqHjNkpwAnYfIu6HSZ7LGoDt7z54FeDgahhMYtuI23E+3xopufyqr
zNQoLpmkv9G7iBeKwhDbY2+6gtECXjFF5vwhz3HQxHMC+AHL9gWwnJnOukgiuJPc
izJ2U0BwreZT6rcY9WRhas59uIOyzS/GEjtyEjfnMp1iT6YUYICDigmC6E9ynYDh
e3U1qy41r/izDFd1dFRAPzVsSjiJWwaN9O0chvQgut1BXIyIbyj9Xm1QwBblaYEl
s644G1ez34hG10USG9A8Mp98D2h/CGfhMCa2rnO9opiK62zK1tK/7aU8YHwqH/Ft
q9yh4Fc1ObEr1yDH2d8OMnFbu9yrsKrJarL8J1pI0v8ZkFPy/sEVdFudr+Vdg/Ko
qnML6fePjC4pxJTCeBbF5DsPc9USpX+hn8aPoS0J7vo824Dm8oqU+VDMJVg9s1yk
9JpEQPX2ZyGbrxysgkESDT2VlDgw8JviAHuAxOdYYsEf77vECvrC3Qp+BE5fDTmz
HHwGutWzZnsMfO4xNKsuT3TUkuKXTsDYjnuNJhHKaBoWqpwjjgFXjm+sYTj8Wkzt
dQ+vYjzz9T8eh2ZAUEkqYsblE5C5T0OogACA7yzNJqfJY0GPw9xk691EjTBCufbs
Il1MIV5OmgDGQMGYfdawq0RYAIj4YGjpqJ05vz9ipt7iqVYZLdjfqL/sOkvWkzYU
WJ1CJU/Zj92LXiTPQUpAnTw8bcLUs386VI4ovI59yJggI+zmecbO2fxtZILc9Jmw
9aCpOeXJziaNUY/Vf0xutY4I8cGM9vcaBbO7kH1C015bFy/FUYYnsCSD0KfPyfee
xbOC1c90bNkAg4HqHH33jPdSP1HIagW0cr22HVrpGT+Ma24UJ2nMmu/eAulxkbi6
M+udF7w5W0Amq2yX8VBA/LxUe6mm+RDcvEqCEgr5rcQDQViqCr2bHoaqX17fZneM
GAwlNrpZ4b1k7Rkb9ccN4zalgaSNo9YAcq7juhP8tWiu+Fy4JukiMq/5I/DLNfgr
eRg7rCUVTFqICMwVIVDW4FMcSA4lofdtBbHITixjAfluItI9rTqgfCwKWlKHU4wf
EM2xHkbBixCWtEf3QiCsuyoHBkpYCcX/jtcEf2nepZHbKLaIAAiechlp3YGmXGDk
T7gmUAQVX4P1mZE63FMOeycEA57JsynhHHg19oTO8cPcfHt6diollVXsXxo7iyEV
chEwdcDsnOxMcc5Hic2H+zhexrva7jDnalJn7NHMH49bTuxry9Mv5wfTKmmZnZIe
BfA2C+l/3VJktCU7BA/Glq/wlqkupMVQ6hhCW++df7WPYUsZ9kIckrmwoZrFVcOR
xu8e3EPD4c3JIfRKsGFwd0y9edsyA1AY5q+ODMZSPwCPzzrPmoQJ2z+MiLrYIJGM
0z4OFr6W9D2XiaRMI+csGMOEqODMIH36/NU/nt/lUSJgxeer7P5QGPM4Tu+fjaWY
D3+QLX5BL/SbM9DUqyOZdH+HG3K/O+8s7yfDrbd/n7fcO25TnJ5pfmNetDo3dddz
nJG7sbTvcDJrurvZA13jNDZpidt6KfO+pD0+ThEPdDLWsp7sIFu9en8cdU3PfgzS
HCE7lfLhH/7RszoBIzMC3WnFu0S18u+ff2t5ulY1n0LSP7+UbFuaVrRc5yav6TON
vpZfBxSq4cih7ekR8vJNPaX6DpbOaYSmVQI7OFml1yvjL6Ala/tjV+3eYUSR7Mbb
WJV5ztmyxxmlylwZ3RF2smiNzOo9Iu3Ka7F8ulh7Ldfk8IEUgTpbeIQdDp6TBUNZ
cHAZFZK3NOSAjd0qivhUIhTe1coJkjjzFoG9UoCj3U3W8QcG71CczyLvX8NFE4uK
mdOlaxK1BQDBQDfRrA3CUwdAC1TuNgeWMqEIgCuuNEZokj3K0vD18KlMmHO4dv5J
iqh0FQiTRLe6RgGZKeV+UqH28P5hr3ZLhvA6gIuFtUaMW9UargtOvXgz+BPOauUd
p5k6mlpGyF+T82lrXxECezsjxLAKeyD1m3Y2YICfAa+WraK6hZOTo3VoSVbyEpXH
ImPAsu4MxFf/jQR2MWVShNYeDSSng5b5U/wY9J/ifmp/9QXcQiRHC9PYhZ1SVPxs
N9r9NucvX54sVUbklk1T4UrtGsK/MkHvSZZAZktYenjPy0Za9C+1a1gLZ8vuM5jc
PZvfvWphD4CuyNU3s+PDBxXVaRGRzSaHB05embHRFd+bMlAZIGzh2pyRRjXOljPy
3er29ehVMoo7ntGwVEREFPcSvLJ1gTPhOx/Qx84GJOAHeZD//DHHFxCEVTgZgJ7b
V8OFmbm9LdfbLCEkXfdfqiFsBVJDjLPtcE7BBGyXBt7GIumF0CO9L5Ncy+YaKfv0
XP7Pcc3C2xEIQU5VeumfMNaXVKV8uGx5Jrixq8PV4DXPuSEGvV2oRbcjdCGQv77J
ZkVTFVVDM1ifKjD5H0d7lyClefhAlQadeCuIUspXuD2Zz1m+DITmjiVNVuv/KpgK
CUFXM42J40pcQhhJfsnYqt+68x7CmokJXlM4oS1ngN9SsPhMbtmCNWYrQF9SdoC/
FV03H9ZllOjclHWqk96HOIkHPqR+x9la1wnky6cl4Bt+qg9N1fkgBVXLSdk3FURg
Doc2JlK/80u51YIJEqlrWlLOEkvREeeGONdjN8tOOPdbvESIAgiHCP0u7VWVDTsw
siNjOxOGUzjwMpTiqFRe1kBlSKzW86Bry9IQkKG8M8T9tP+8r2rHFJbdALwCdQx8
idnV4HctDxrQzpZdjZhAA1wcfI4a3/weLQg6UzMx2cMOOFQUgtTgVn1LkD/O5dQx
r2zTPKofJOm4XhU+cNsiXvRm30+LTV0QOeJ5bEn90TSgoT+TxlsQ9WAxtJIhl5Dw
XKW/yKXa8MoZ8E83YEr1T/0GK7OJWCzw4lhOF2qOtibVNuX0zn+b4MdVCY805NjR
odVWrfoMKuM+EyvKE5RpNSBAYm9pmJvbJnvVfgs6KjPVh248t4WG3ke1wmVKZCxn
bI7xYDGOhfqswmYrrHwVWuEBVrCRaLvvBq8v/c63F0vneXB1/vw3gXGpRQBJp8GE
7+5Gfz9etuBLzzjgOFbsCaBsTrsym1sLbiJY8OY7C/6Ol7Uv2DYukg1LbXLv9ncj
ROlr0V84NNH/BJO5DbjUMwsX+4+JBvkPinXwF03EFOL5fXR04AT1lUFRcda9B50h
c7yY7JXKF7oXKdq7AcW5OKAgQp7nsmBKfS73N7fX8+OijjqHTs9LmL5zD9I6tiJP
fxgU3vHm5fhbZgq3UJ/YBFZ5y/T18tg1axKUOQeWRquhiA02nX9ubVT19uvfcGo0
sXsa1dMrK9dhrbiDy64ShqdVrfSQq/q/RBPUKgkZ5uQUKBJm+8nEI4FuIfb+AzxW
9jejxTprxQuDJRKS08aJ9URQAd9aLEY9Bbaah2/B2xz/c5Mn+jR9VPFOwgRL0mKN
xIroDdKIHKw8evGWpoaf76Q/00nSaXNO3pjEdabGBr0jGobfcK1Q9DOeP2Rj/PNJ
tFSgCED/QW9LiPrOrTG3dknO+GSrCuveY+DSV0CihVE0oLRqwTIFJNuJ9MOa1Sw/
+NB/FMl36rAm76twd+d6mvWOimYV9micG60hXR91E04/qy1I+XiXaCxWRF9o4W/m
L2HaD6WAsx6GII2Q4kTVR78htlmDCzRkrzk0jV1Emo+U1cKHxQNDcCpcfJ7P7TDt
Q07Dp0pUAYGvpKTrK7wMNo4FX94fbWZxYmN0DSHTkAkVWCCVrw6IUX42ZC5D3NID
fwQ8mhuSvCqkzlwOqBmLocR9vHWcZX7OoawIro595YjbjNFM0C0f20r5KMtHP16X
mGpyAlSmC4xysZXO2CQ+Uav9i3JmuO5Uj3JslmJQntqTYYNO/AYpZFrb28O6sxe3
nd+thRO2Aab5xLmajVH9ZSYz0iLGxw1Oc3Th6bzYLj8NX9wJZX7PNl+H38tZzbVX
ahPzrgI7ejtcIbEhMtYlWan7ifg0ewL7UnwB0YfJ7VzRuxHc/QnUWPByOC6NJr00
22/xWNDV1OT4nmD643izRU2pqrRWEa0gCG++TUXqjgEWWt0bG/flQ8pY0uUqV4z4
7MFpiu/JGgSigyTh08SRxl8KvXiOa8jPr1gfhFVdsbp4qVqhD7GxMc3EtqF8fHbu
7ldIui6d9b1HfMSyDmBDDPkTHz8PYI7VVqsSu/fyInxOXuhPqdH4xHiLk2D4xvbB
RZ7EZCfC/HqziMcEpcHD53otYR1FOQHpOgh7LcF/ejhV2D45Qls7//HHNb8lTxIu
EDjikOvRLJWQ91jbP9pGKQA3jE4p8XTTrH0vXhN1rD/lZwf59fHeVbhXMOprVvbV
dCv5io4Kx450NqKoJOCDpiwqnp7+SE3XAKBdRVEf8WzBpRkdqN0/2yETWu6DYYpl
X1TgMuLBYAEzxMZYuMrMCh0S0Ckh0p6+YuTWPTxyWVLxiSccox+yj7XKf6v0RPRR
ZhFz+7/rTxSyHAw7EdX7qkKsIMYV04DOSMkqjLSMCDAv0XYvVE3ffewF9t1/21u1
+WKr9gUKjCjwFv+/UR1gvhzkZ4QDz81j9U/x8GPy39mH/+FuswkRhn22ccb5EZiI
F2CMF7H6OILPQWVXxrWYJNjZFXHpwuFFAmssuW2JLRQfUQ9/Z8G6Dc7QuWi7pKz6
87FWO7jly7LWmrkKM8btwAMnKQ/B8YzMwiFR1aD0BN4InLctMIQhHUFqv0Gh6DC0
pGdLDzaMoU0XIsrfDunSqPFati1b5AB4tgsUZ7gx6nPkYNM4T/SmHd68e6sPA9Ce
K7jyqHRcVRu1+Ps52b+Jkg+8G59Xqp+4x6kXlPTHAMNztGdjeL4NyzzGYSbWVnMe
lcRFWVXIo3VqmpWNxKkcgz+96R/2j5/W7tK9ZRZHnlZ6ZdgTF+GJcmT5AgM8U6WL
AfEsoykiJqkMmeIQWm6hmXbVFg0H5LV9lswLxAyEk/5nA1Qexszf+MuS4wpZnhzr
qGu5zjn2sYm7ks9OxKqExZ+iRUTItbiEDqEKGjBqNmrmnb9i4428xYbCRD5RdHx3
8DjJxMx2BWFq7qGN+ZEKO+6FyxcZSwSJi/1n3L3rJoB3eWSLhgkAPcY+oo/50JdB
7qDdCjYl7pgrjJjZnV+8/OjhSOYCyeeNlMzSFdM+d+mYtzlaljEB4Ngb2PS+CYFr
3U+p3kzhgwKY46zW/mTWmmuaD/yD78vjTSmkUWbqYAERNQuotbefAZeLQdTSK7HE
xY0k3mPYXjQGREWbp35vvSfLPAqG/ON+6qFEP/vRJYCVNW7d2uEmsBKlqqMbfe/1
4By+W5ldm77jy1Zdh8pFKhEIc/kWeTO5qPzPNi2BqJ3TFb0LihW0GrFb4C8kV0T8
u/YbQ6M2pncdH8wLRkJr+lse0mSPcSmfyVVQGgIdONyJ1Ob2gBq87O3tW31GukIK
oleNYKuFgapCNN2qMqNk3uGLapQahOBvVYvBcb+TobMi7Yiylde74l07X2u7qv+P
2CcURW7NuTP5SmQYJNyQ+Co+blJ/uo95fAonMExrGKpOyvTHjqLwoLHhr9V9GN9j
fbJ/JK8djFyUVe/+LMksh/+MYuyTiN09RIT3DgcNv6VFjVWNWMO+ojcbMJ3Fgljw
x++Sr17xyApv17idl0iza5Z/gqXduW+ifyPLdMtSmZvFnkCoFMJECRCAdDOm67/B
au9Tj521AND4VwWZsdJ1wwY/14zFpYE8EL6idgZSBKjc/EGiQUgS/OpeLO/PjSE0
L5eiRWV+Lz9w/vCq107uusL3wdezXRw8l3VrSsWZoC5LU5QU6jhXY64ATkL2TpSx
R4d8v7YZHEg9Mvc+3cGsVTY1d7ybwpztisBxft58TdkpprU9UWuxD6pPvf9jlIuI
tyx1h8n6MOl4bJPqmv2an7+lUT0rnFy9Tmy+B0VaSVS82Tnlf2dA0sRD7C8N2nj+
cqdFdQjl7hFNdT+neIygnsxX5w3aVJpZniL240AZicl2/mA/h+jtEIgy5vri8s0w
Sn6xVIEyGrlVHv6YMLA9vtlYtoclZ24gG12VAahGstJfmnsTg8qrp+Gq9+qNeSRl
X3/PXk7qr5adLDRXRTQNsSHjhBmIDS0mr/Jes+0H658KW5kdBvEljH5xmfnYHuUM
iBajoeZfMQrlcw69r//x2FXEpcXawRveNTzsc4f0zCE5IEHqsdew4aukN8FIKsrK
q2vH418OyjcCvviP4aWetObcgSwsVp3k3ozvZDx1ACQElSMU1Z0zz3lxMDVKvqLf
kQ7LbTRnIKST5/g1drLaWE1nNO9bPp6LZ+9lfeLnSjzKlBi1C3tXiC+KglI4CgCn
OAQiBHYWVS0Hp+jtw5ywm5rk2fEOAvWDoE9Gkimbyk+Y0O0dmgm7whoLFrEAg1wT
bzJiebjbzqoiqONhpKpJvSgEclM+59qrGb7HzFwAii5CQBjKFzENdusDdPsPpDC8
T2GoHimPQNMuodZ03BL75gIQkDgrEL53bjs35O7LmFYCNQ6CeeUizPZHcOdshDCe
B0NN5nkVy//zvvd17B019W1vZMnEZ6w1uHNDoxwrgvLEdJnAqPopAIsllG5k3Im7
Im9vl4IUdEpV9359fU39G0K3N68FWF5GRZceGRFj7eManE8YNofR5Spu5S8ugEbH
PnE+vpLXRfJ8W9wbqg8fNND5vC6hxWeml5Zcar2bAzvYQUR8UNMRDwtW2+C22ldI
uHf5vftAOJY6uK6ZCXNIrUHHChjNWKEOd0g4kebZKfPdW9b8FtYFfU0K42D+o4EF
dYD+aYoQLbInerwhIYW5OKzOHskqSRajuL8MTBM7cRWsEPH5tt7Zy+iLhQ6USKCW
z9WHNisbGQtnoc1TCr5z0MPkurljAJkovqTlxJmx5oYBheZDMkk/wzw4nGZUS7qB
VayFHGtN5bDM+q65BoBtOYRV/1qN5m8cFONOmkTSraqh/vHLmvZvTutel0jQb9SX
xwBOgUQeLOJavMq4Ug9NBWtVSh/L/Qxyltq5DbiosVwTZIheVBzh9o3dF5RKHS5C
iUt082/dLHXctQijYX91SdmFzORvYf1M9gauOEWUouiGu2wdVuD2JmKdNE7g/OoK
6c2zr9EHnnnOtbaXqZlJ/jVqxKR3A8M8E38LYFQVUnhhUHsRM45cUq9rzGK87W1R
S7sggWl+tTj40QMxI4XH+cGh6eCnUrFXDsEhkfQXod8RK9hlxjuGf6RIW4lYpQqF
8xq8mka2Lx2G7U72BmiARlWdINQXjpWS2sPPvwro1q4aECYac1uK3pI5kcIZrvW2
mydzItE52xe2mgFsRzvZfYZlBPBSentDFpct6AaznLYKYTs2DdhevB9WKKFlPbxc
AOjNQprqZdGaO2x1GuKSJPr/jcpu6s/n6+ryzrkMqRAZgpZs047mgUzd0pdSUz7H
iddAf86d0a6hCNpjZc4qXbtQJruxTkaCZXiaU0zi66WToTgbty1D9455PD+Ag4Oo
qKNzWilliYIAbBAFcDj4r7fpIP5Ll66pATgXZswXUk6LCwhNjZdALre4UGO5FX0g
N0Y4y+E6Na66B1eUXcH/GG0Gj+Ymf5Kv8ZPyTdqO72x3vG/KkREoQmlAX/lvQpRN
GUwlXfhwneN9UqI/sj3WrvcjIXwAjttSG93VOkX0mqvhRz+Uf2kVo821ST5NWdtt
ETTmMZitS3UfDEjrZhnduiiQgVJG5tYgUahYIVzT0coolnOYRYMpNQKG0YhAG3V7
egv8TvoWKQqXdMuHWmY1LRyHNGmsRhwsfPop92fPjqSxl1GdlLwVBpzR1KJ9pGPD
gQVLeNzC9Rm7a6Y3T4T6V+9W0384pvnkNJ/sy+suCNmQyF7kXcjE72+3jzytGLN6
W3RZgDZtZWBGOsFv5tLkDNPxig13sI6ZO27fHxc2jud362JMqLE81uzhI9UCdOy4
Hz0igKgdpQfyCYLvecHZb9mLLJbyqd/bYy/6d0dpzCO9GioOUOujcOALwqTwMYbW
sm9/iBAKWgtvKb5FoxFuXdYvxuGt45xupU2ZgNqBRVpIehvVvy/xFvg+yx5Oxdn3
T3L8S/0xz7JNg5B8ro1bvgBnEiYK5wNx2e/cIaOG8gbD2r/8ySN49Cprj33iBPFR
yv2dTBFHj+94t23srjeljP0QdhtHHmRUMUUP07fz5pSMS6EEE0TkRLGAE8In+ayk
00Lf4nQDn5Zupob/SYTZzl/xOXWd5B3PTSp5Wml8LsJkRZHjEYvDTUxuBf4DX4hA
DXTiKcOavM3p+zKYzfE7ddF9aVwgFFvPV65ITR/Qh6O/fSQq+SOaXCe/y0nPmfTq
eETNqVvLPv/AfOtSHaz+/htq5y0jW+DVhxztB0Q8j/yx9Nvt+VgRFTuh5K8dvAny
PFw/U8Em9ro8x5gCX0+Brqj3PeXfgozKyuGCBCKzlXM09xCLNGQeAilraFVmMQET
tQc2ACM9FoRQh+vnGntsuta+1CKnUbDajinW9wPD+aeSOolTVIy9pPP7QnPCj/2e
SgyeKpoV18pqi7ZRzURegpAoTvjs51if02xX9gvyE2aRjRDapmEu3a5w5R67u9CF
IWLS+fno5YVTj8xPsKEgPhzlDlf0sUjVzbjDBEP88p+EV2uhaV3Z1stLYrdNVdkm
AP18Zru70R+i/esng3uVNgbNX8sS3X3xJlHqkTAYR/v6/HUKHKGcJ4/QGXvdsbhQ
zquVZ+iyYmRzqk1S0w1iCJrWttypz5iBWPEi9yL//93eftoEaFa9ZFn9DfcuJrEi
BkFddv163A0tQtF+9RDo/dHnKf1smtgOvPDsS6C2XfL/7LkzV9HsyEdCGqOUmeLU
hDBOsfF6PXALJHTUn+LPkK4MDJ7OvJAeDvtiOmHisWKsneQOPZxzXDKJb0MbMIT8
+IZi6OvqUmGFBmApDdTv3ztqQ4plz4oxqXFK8v07TlrgV9oekrweepb1lDYW56zC
RHZf2MdwamP/FGo6s9rM6X8Vs+Q2NMFxFAJzbYLbu2+NYN11XMzJbIEEC4JWFNko
sFZFa/4+0jD9E27F60P4yk1/TWm8tGp7KIVuZI99FLK2wAsbsk6Yoyr3MWILnua+
QPjEVWNAbZZZytEPMgUTj0he47LgCkp7s66AzAt5sbMTuxLvwlpvt/uwVCE9uobA
Ss/bDLLZCC/e4QkDdd8Zr0JMchF3reGdJRdnkSz7pRqIZOIsWxSgiaPjWxe07F1a
59VlYZai1HMssmYKeuKA9A3b4ZXxDpfZ0n3XaUM0B6cJ49JhppWdzgBnhtSYCrek
oobDIGswoz80reuo6bPtoP8N8oaFcQVQboVFZQ3/h9ZkMTKozimTiELBGY+pN8Le
/7tV4FaMAmX5vwUK7aOz4lJv2Voro9QCjM8gTOmbuCQBhgoHDjCu72trd5Y8EZzx
fyYCwfoVsEeNwjalEp1rn6qb3zsq50BVSyRDk5TU10Hazap/PVQO0YQ1DTUomBP0
gliuNqzfNqmLTnbzquxsAMeQD+WCfw3Iq7hEmNaJiy106YPtq1IfjK7QXGr8prlw
yHAq6ojXu/bwJoG6ARIUp0x4+4Vu9hIUFvaFpY9UpGVU7KjiJq0njVE7EmLL9hlU
SYW8/qN0rq3pG7Q11EZaSyrFCw2rgMhNpH3TFd+b/xEOi8Rfxx2sIEjwZEALGPNH
1wm/BPZyFErKUB1KlZ/QY2LKKYFGozXADnzrXZ2a3HRBr7L3cm5VENO/SD3trhXh
ILy3y1pt+Btx5gCall0svOy6IEmcsSLyTgtafAtT/D3d5yqfVPE8VpqH62oE6jaS
h0MZxs6yMIbGy/nTUCpVQsn/1s9IUF2XJU3W3kgkvUusfyqI+jmiYEgQsg6J6pNl
K3GgwOhX4W46UiBfW2jSldykTr89W5C1aVKkQrP75buNQj4RWYIvMLaIg+6MaY3X
3+z0ls2FlfRH37sdj3NCiz9NEi2omB/0b573/lHBUGj0IzB/ThIpj4rdkpNfS93g
mcxtRuYRAwcWmyKX0/Zfdo1j0L02pV1CaxVMRGdIYYTlR3UrsN4RWK0i8sXMNpNA
nmwXVaM7z2eibDanQ5VcY2br0jQXyIbbVhU3OWPlFSUYW4+693uCS3Zwf/F4tkby
JZ2PzBrxtba1MwamdP5c4AJFucHQaRhQu9NHyKBfOEX912fBpJ5eL0Mse050FW8K
SRlO155odriMxDEP/Q9tnMACSzK6OVNqoVk9f7sFpyvBPjPzxUqldu2EBsLqyCYm
+1xkd8nfArqWKhLniFZHkCPuiuFaDyYeZ2MQa4RdLYD9VbhxFx6/WBX5GtxGsKpL
mRF8ZvoUaSEDUrnhknM54NWDv3GL+xlU3NTq4GfmjT/wD5d/nixlGXiBEI4A85yO
PvjdkuAbB0ioxHSOXb+4fCmJCtlfQsZEm4ExphkLIs/HNEkIQUQTZ01p+oHvyuw/
4Gkz+3yDQSX2Fbb/MWBHJo6XQJEur7hjJFE8g2vqLa2sMYIIaEOK4dPrl2M7LNfk
GQs5J7lmMZX3id6CxUYvUHoZUZRcT8S7BFf44nS9gfqTOkM6YZFbbUs8iFrSR/mx
13EwcRjLdGsUYuWheFHvBcfm9BMidCSs8cDSAKvERRtR3mYDWEMLaHBsn2dtdwl4
a3zgIkekRVbs58QruyCsPPXgxr9JJxlzVzyMXhFB1V+gJgONTIkQeb0MPKjfsizI
Y8D3jaNaiANvuVrkrXZmw9Fp/WbTxCAo0E2O8ZJj5Th94lCTZwLD3vVDNga8S/5V
SlGomHDnWD69ulkND0W3tjqSMwK4iGmqrfvpzBO1yW9WE525YCfY/ZSTP27RKhLC
OC5Fuj/4z84gsbWofXF+DHZI1YlOMAJb3eB0gUpGd9OJ8+2GtPmnt8GWkKIgpmfd
f0p7fsV27h8UUvnwGWzfcBdm2BDF3EtrtCz+wfqzyzuuIVMhNtcLo97kiSMkq4Eo
8dJYA/3CZN9FTyYU1jGzt0iS0ZYYu8Tl1AWCJ3BhB87GghSPwSs5XhXjZxTAU6Me
oA05HitKO3rYtMjAwDz6qaQJr409fEBiKFw7t3ggY9tGJhRK7RLum2Mf7nbbpZg+
081PVxO1RSGGXHcOutq2L3CtRGEJlieMvE6/8qjuaCiVYuh7Jyqd48P+AhmZpkxM
y3kyKbBK/q6A1tik9QWQXroBIE3jlOp3yDh2zvDbDG5G1J27lhOJp+lBsIUyehE+
xgKq4WFw/mNtmFvSnjY7VEHIZ7+278HxSS3SLv5+PTPhbM1I5KZ6OPIccrU5+6af
3mC1HDIbKsXsq/WWPcW7wM7bP//wsqwID94QxybwtpBl9GxNaucXYsiKBEy52cKb
9RH0eH2+UlNh09cjb+ON9YzaNY6Vbpm2oiEqebmdJAHP44lQawxmCpYh5akzcze8
ogOqpBJbZKGantvAtpT3jTBitlENmMsR2ElXweMkhbzC0QgUDRD3u0EfS9R1jWIC
zsK9NF4YbfMp7Xgt+u10M7QyOZ4DCaZowf1/O6ncXZ+kRqxcGRRm5bL1L97FcWO8
+jhSdVNmt6ZXN3bTMy0zNReEEMzKPzi5gV75w+fsVsslEl0wXmyfApRoEeoCBFwh
MiFHAr9N73+CHs1W5W+yLW++Hta/bW8w/KWBDh2mr0jTxg9oUlKunzTN8A2qrv99
qzKnG7SA17baAiOo/QEyFaAYmIra92FJx4soTw1zlWBp8OArVYstSyNmthnSynus
2STHSFX2T7a65+aMGmbNu3A4CfVPjAlnSLM1V2g3qk39LhZjXRZGF9wJ1pmvrmMV
x1MCEODM3Q5bSJqrvTQrN4uX8RUz83/PyTKOtdX4cpN6cIK6htpuUJ8AZcEyYpgM
CFc2KyHBE5fKNvoDmOChTUTh2XhRZ+mfxN2hVN6prfcJ2Q0TdMxGv8+r+zIIcliP
jGerPJijHEc7zYl+ACgefXCKlVhDTi8zHUeKXEm8jJnBSwe2hN92UzNpVIg4aFoJ
5GDbCU2K+YyQ+sIakHoj9ix9idKDx4VkXZZnSdDdfJ+ECDrxMpW0iAcdZ50tWHUq
31CWK/0VhOanKCzMTP+saGj+eoBHUSjhSPkeHtuLX2JTRe7Hsga/X4TOMFW3sdL9
R7HiUUFgRNNawXkI3qm7b5bB0Egg11fjjS5nlEvU2nZqCq0Xm9r3zBu3hdm3e6wD
EnEoqYaAREurrNHySzTtyUujkn+4zWFQxG79+1GN5x6mjfl56dcHnRNluScOfEig
H/66GMyhD5QnUb+y71U/vDXeFjgd31KCQK1FCorAEUE7fLwNAFu99P9nQAG4SbLR
sMo7SQV/N1HMffGhmW94UAzUzLd8IqSTKzuTnaM/PaaRdJD2AaoVuOPFnF8GUG7t
ZCxgrjWlgtmdb9pta/+t2rXWo9tp64VFFs/biLYi0kVN+0P6cHNUnfBZ/IGJ5HS7
d6Lm+/oT68GVrTOMQeZgpW0Eqv2tNyBR4As32V1gwprnIL0oDcwn2+yBst+10pwM
dme45wTYH1uK8e5IWZ/McD9LA1qThEVlJaymsMI6GgtSmOgYxVduLSZSZE3n1aNs
M547dtkGLm23+APwqj/N6Zt8KH+pOXERrcDlxT2gL6tlKSZrUEpn4w4C13w7YVIH
uzwIHv3jwgdKUUX0A8f9LBwAke6OkP5qvljz5hFv6X9EDAot02//8FSrZLqMdGUi
HKG63b4/TDJJgJgIDi00a9DM5bTorlVRaKJ8TUwy5J9DGJQ0de6pCk91ugJiJiZF
lnbW+gvDgfzgu2rGTqKj0wNbq2Nl0mlS0ELQXvta6CIiVjYSd7Pndg7nyxhCXQ4E
2pXvhwspUjOYI4YoLFaTniZY4nMBi4lVGZgqfowkUD3lDLHa2+ahIJZ5OQ1+xY1U
eBnuX83qD4ylIzLOVNAuYXEqwVs7HoS+rsSE6cyA9sy3wRpB6qvWGH3LOgvO7T4A
Q2SNMyz7pNF49PqW1G4UV1SoK4QUO+79fQC/7oDiKHypUV3+8yqdheUCoNRSEnIT
Y/QiKtSU6DRWBjSqKyOv4QBlqX0ONqwUKq+0O6uh3L8CylP88cH0tu8d0+ZZRT/q
imHgGDUv/G3R/E7EY7w/A2o+o0ld62kXJryQ3QoxBJwIpX0LxEfczq3kbE5wvmV0
PgLxE0RhiUtKJIWghs68JHBoqX8kgqBaXEnh6aQFoWJ8uu22KsH4lpAAeStF3Gbd
0cRenL/w1yKdwfaNP3rD6GWp+iLJAIeHyzzyHqLs3KzcCuCIzBuHU0HxJToOJmEp
LfElanTeU26PKBzF+G9qdqecRxwerGuoTZJM5uLUL126VI4+ITdzPoOm+XowXR5R
wW5FWtFlENbd4CHbeZqTXJKKKsLDY/WJY0q2X2N8iwZi4p4HvMiRWcoXSHMysgiu
ACw7tmIUSAjUZvxwxVNWskmeCB0p/8IXk5OpCzEKFWYyG9hLFMLsrlg2h4PW9v4l
r8DkphanA3GcROatJYyflILQUbjZfAfng9FE4JfcIwx17poXQAwQDIn9VzBi5qXI
V9xH99KFhyQSh8Agyq4BFGds18p0XSE6G59PShP0T8gyPgGk1LV6vstZvycIAErS
cgVbGycXnJ74ewEmz+n/psBeTC5N71Kzc7BHfq7db0Iz85be0iWnUoi+ClFHyLdK
8HaXCJdjab7r96E96Wq7r4nJ+O4jsmPhCmGmc8+2Qb5KzNVJiedS0fsGtM4aVYMi
2pT17JSxczEEjX0vamTSmI8aVlT86o2PiQIggwHuXdSnh0mtyM6qC1U8qf6T5KII
CPyJowt/t0PCBwvB9UnL1RPag1t7It81WWWE7gX5e9KY3tLgFuMhqNUAE3N8UsFC
nP+CksehBmyXMFWE4NMWQ7aMo0dLlaDm8jLk01NYRXa7mesi0Ztdw31B6yrecL4U
/74MDUntX5VikfLxtumgzJrjKLrR7pnafXHK+Amem4yEVsq0uUjHFugOcNU1GSXW
8a5wvL6PqczQVcTrAY+jI1Z7F/Evuz7FiL4oWO160STwOMXl5zsAq5W9STtdwise
Jx8dhd7p77Rva5yQVqzXbDAIeOc1ujqmzpeKpwkXUbznkxkqHxtKtq3PYgr102gl
2BOFHACs3odKa0zFzi8xSXLwp0UiSj0yaZaTvfUd8XMk0W8K86c77KYIu5L8ezIa
K3POvd7n5l5EOCxp4t2HWd12GmhmSVso6PdwHx7siJyj05OEARZLDDdgenWcIPhW
t1q2IMdkQksT/CKSUGTqEywlINeDn5MW3+rINiA+bkI2X/z0aejU5QZ5koki6fxb
ZBuCh93YNskNxy+7YiLAU0ZxYeqaSQVyGa359FYs4vxGGYdkmsEacJ5guNs1BrGl
RwgXJJ51COhBwUQqM39HYZsTpVIK1FetePMubu67zttV9QyHntM2zYUKO4kg/i+o
TBTwU2bqP6DyvhtIzY0jRfisECjYuIusNEsPXVAWJ5ehsrrCxUs7/ti+3m0Q+OhV
A+bOUsR1hHmPMJze6Gs9dLMnVlbZskpK56FF92Y1utR12SIbbCeckQm4HlBxtLUm
e6px7WbWCW75yGG70dLKRZdz+bAjmMPOBE6vGDXjdskYIChmr4Ea50slj5YtYzkP
hYcr4YvU2163+tpQWTzSsFmJCq8jWz8Woj/JClXnmwrUh8kn0iBy9423FzGc/3M2
vLO42RAbrIPFvXzbMlvus6XaNGou08c+1enCO3utUz0Lh7p+Tjjdcvn+FgjWDb6g
90V10h6IKqtxy4GF2PAblSH5wKKD961/0xbJYI+VRQkTfmjTTVVeJcLQW7BdAWEA
GUWpdgLbaLBQAi5+lW6yxpr2DvJBiNPOIHtiU6CGDDwg5HD6vik8CU3u4Iog3qzy
h6H8LB6x+j1ieRSyXeYDoVAhTVbQC8nRyQ4ftPrxwODpS3/4ipx4zZpUk0UluGY8
J5Mhqo/jcU78kktTgOBLQiXKx+Amm/BDCDThDWTfj0hCed0zvUL+0VjpGHIJ0B/3
g8ciq4YE1bY+ugSX/Gyxfqht/+Ue/eyKMvFRKLz+hfxcBV+igC2jvsxjxAC4a3r8
qqY7ikFcrdcB7gP/P1yOBsZVJpSFZr8AfnkrWCYaZk6/8yYVplKNOsO58vdu+69j
Q6YaNycMT0OKz+uxWZPVwhY99ghP9e6iT5p0U3balSfiapFBa7X/5mDwiuUPRgIC
o/sCxTHyYhszEEUDzjsMnbm3gYzUBFp1BGogq/98W+6f7wFQLV7LSAWslaIZ/TJq
7a17jr5KVLtQiZCAqzeLeWcPXvW8iD5JDRKpGNsSMD8DE72tPv829JR0RJrYebKv
HL0v7gdtF4La/514CXrI3XUtqdZ9cHAAfJcFaKeFVZc1ujnxN/Y6ZtT5O2xHg0kN
7k6iiRZdKlA61m6Di29XAVcJMbVs0w8dVwAA9gzrnu9kUdpHY3xd0omGwtdV3if9
HSRDeBf/mpvH1DbS+cDFPAcLlJhTalDd/908ATByi/DtIW5TbAKhPz72F3s0pjKz
lFTYglQbF7Ab/LZpePFE6hRyaNGavFa+dfuSspojBR0H4NBlgN1ZDtOcMvuk4wc0
Xx5yYZ+KjoaiBpy7A+KZ8gKJsu6SGRWTx3O06jwLKW0qrfkbesycluOnCE4BCHgD
HCnTxnQr6NrrN+3rooJCRhrDUPWEB9sVylrCIc1t2cfHK1EafxSfTVZTgQI7dGcW
avbQUfBIg4EITqcjqUjBPwX65/y0lbrh62x7FwD4KMfyd7vU6oyDjoGCReRCrcYr
jHSTmIjEWudlKOHNoaiRznTUEGZAv7zR70pcJiT1PjkZW09WppqBwlE2nW4VPHHU
TDV/13MHJiFYpqSFUiM7CzHfM8IW0wlnjlomEgxIzJ5YNxIdZq9mP0PlbY/ErWax
fIJgioL9Y/7hJZFI9ObBF2xuGinfGicp/ljbIv6F+tBme5yQFbxGfDivlD5z/06m
lb8LqrLS/STQsZHSzwrYo6iy2wKQe/c8gxx1RmSEXjBMKPbTxa0zbPyPKt9z/dlu
h3zX9QIN6MMy6ZHybsAgPAdWJTg5BfoQP/YaYoQswcmTNqtNbWN14okwsMIOhv6S
A9jGKM585x2ikn0IcR0oTPXMVUdavGmj5mGz2tqpZ3puFX1+D80Op5CoYsSbey9n
x49rK3/EYuJzyooF6tE6VCdxCWLHngTGcxctI20lqiLWxF4HfWeYaro2FBPTnbV9
+E74Hok2KEMfIkk1W702Mp6YlNijdLoDrt0oenQ1xp6112lzY9bpVKsscdNFyJOn
bBXw7J/qgatBVOBxX882RTovUgcXbilxT1KuNtuAgRxaE2L9JF04G1N/KDiI5gZ9
U4ZxYg4KbCPKHp/zrtzUWzHQkSEiUAf2nQz0ixmhKD3SLF5SfyQAnA9a6RxfZpLw
ds7bnC4UM7ahG22pQQnPdN4VwQTULZUrxkT8LaBHp0vb9efDXDDtMV4I8bxb3LlG
6qYVqGp/R0j8K7yGGJtMhMB0uB8zftYgfTJmQLthK4HN1N/GF257dQhI/SVpvWEC
g/N8llNytPcxBH86aoOR1eDbvTaXtBwwM/MtJEpj+SLdFFWZGboo0G8ir2cG1XEA
P1WDESaiyPdClVZh1Sc/3D1i18QsGWO/u5uDNpMptCqKyibFNu3zRt74kJhu7I4c
zDMFUwVgzC/X/Ni8eEhqmyQqo6kciAkhMZMyAjezswWNIJUOmOOM+hjT1pshYTNN
0xNmE9JjqcZwTARk086cYe3XaQekv3U9ZzpHKkh31qyN1nJ+v3wajQibYhG5k9HR
n0q1sVDlfMxs6z5LpQDwZqkJmdNGtgur1YhDgkMY5mfWZ70vfh0U1c2ubMbdR/Cs
1noq5QOFk7yf+LUUhrH4GEsGmZ8Qfccb1NKvNZ9G2LedmBacHVcSLOac9TNIUcHO
j/JA1VfNFl9Ey10v5h2pKPRAhISToiHtw6MnysHkyHMGUmfw3k2qA4www85kc28q
uc/PLUBoxvzOtssGgob1CB1qUnJj1uYbCQ94eMGWh0AqweQa3Cb0HUNp4nZCYqMi
F16lTnElj+Y9Js/9E6RUG+c/5jy9ULEqEYSmPY0bH5X/aKzTAfxZO86LXRfdr+dp
qo/IBeXcg47eUdAHWprm8nJIFniPzKNq1tu22sZilrP9v2VXSGZnisqOfzCaPs47
WHDUNb6+lIaf2JljZN3ipIB5Zl/K26uziorxvYKk1XlgLpFFkku0oMkNJG/5IrlB
H32MvhdbyQXUcwWJ1psqdTFfDS1ovSIQCDanLh8SZCku6TmkFxdwHQiYXzFOFQW6
eGSKuLYNg7nfa/zPgUGtQ9700Sk7GqDAJglN26HWXsDrgrqyU5EVBrO9yA9Pt4Uy
ZJaqi/lwno7VkF81+RSGne7o/IPK/+kp3UjHhW22qZgfDLSd42B9ilAuHOtMJGrh
YKXL605xS5FwQPoTwEfwhGVvLjEbFBSputvMUplhVSXrvjPKYsurxgTFqajrb6fs
kn/yYYdewv97Jr0d57RxDHOa04yafgohgGLKzp38X3t/F7RDXALV2fTwfTiprepJ
xreWf1Ff310FF/URBLWmORz2ikOrND2FWC5jKRm08ZZuIXWkgJv5fUyIyNwQ77Hw
2NBgirbMYM6jvaTVjHgfbKf9YpJffm17He2jcfsi7BHq8RUKS1yysy401ToZzmi6
F8uYhWcb7nbdx26WeWpJxGTIfTg0ECViuy4wTIff+vaozdKalpE0uP/62E/zLgTj
qJyJyKyomGY6Yx+5ay7SRhHkwame3WmvMBYjp7D04gMABh8ZscWCqZFzMzUT69+M
002J/N2IJGngC4TbR1AEfZkUX/9HjNuOVfCsa1hgVS1S8LzMV7MS0YFg9I96Yn+0
g6TBJDXe3a27LNMAtxriM6OmLfJY6STpqdANhbNCoXJ1BRI2rd9wIE5RbofCNDp3
wYaWcqudew141cU6x2DhOsx67Eu1ysR6Loq+chYwahNP2nRCu74ourcBJSb8uYh4
z4m/TX8aQva6eYMRdyVRE9Xu3dOBj5r/Wh9gdVyi7tfLsAEvVNXSoriCdS9t/caN
cw/aO9QktZvoIYtr8es4/DKduld1gmyEvFpDp6UW1S5Qu1EB3wvwHhu56EkFyhW8
6z1WvFhkLw/4JEYrs4fRflyXBKXL5wfUotecVc51wdCbkEX8AUH/Juh5+n413PAA
UySOgkcPjK1pPoeVId5hUg1K/z0FICLq4GLv8dtZ4k3oaMve1VNBf49tPPzP032/
4xMfWH/ZMPQ+kuNN6xoM7H0OB09NuEWb0D7SPbXkGzaGGfpa+yITj4xW9IAAIsWF
mavOpyLHuffTw5ZwLqZzzE++nVGJyg4BDCzo8SCiDvOlzP4R3ScHjG9DjUeSoEuo
vv/Bix2i/t1Vr3WqMyGMmdRZbruvcwJ8yn/ibEHbFJP6iI8cAaKNhvDvnRMUu4Gx
F+t/IBGnTeBvMbeiUodZj2gc6neArPxITLvxCMk1HADSR5NpqOD9XaqC+2B+v/02
SnFMgG0z70ojsN51fyQh83YiqVP1O8oc+/YAnYzi1FZvIjc3Vun29kZvu1hWw1SD
fI0O3kdMysnCmogo/tS3qFJTRCcDBta1BtPqVUDdIa+BiCuXQRYPnga7t6jBjATC
gKKmrj6m/VDD+5CZclAt6ng+VxnKHnnDMgu1GP89q94GUXjsyslkIglF7cgzOjKV
FXNUP8XhYw3DQA5OLdj+kBb/CrWnMsQZhSYy3R1WPXwQnXtuJEcU+fAuPjpvhra7
dFElv6IKoPoR05o92/+O7270R+GvFKfKGxUe5upzAxXD1Bxy1ot9Zhlfxxts2zm6
9fY81/YWg3R0bDkgmTpFWUylByrO7Kgqnxl+MdGvnJ/63rRezmKzk5IdF4CiJJxt
FvGqXJqxostaHSpGoBvf4xq3YQQKm1Gjoo59j9qiFgGSoYUuZ5CeeZWK/el03vjv
/MDYdnZ6OL7JEWhIKb22i22oRQMUkkMB9eDd3tR8+2KLePbwpRNTgTaS77roDsrD
j7f8IAbH0514zBMuFoMM9sQB8HkR+4D/6jOEB8U8xevgGPgWaffttCFdVKWHhGyv
2vNNSY+iCjrDJoiIhhNo7Myz6xnJVlTcMQKQ0I155WUFqFy7ivygnBJKHlmUgi8p
M/N8piaXXA1Ddcp5Ua1plAy8k1kC4bRGWgmThnFAG3eTAMlI18KFV/mj9IP30j06
0VNhazyJDBwdhi2wPjQDhp1w911j/UzbjHwxn8IAHins6dLLtrGDQQt1TN+/nVf0
/A0UcIyh1Ha6mwrOVrg+BIIE+eiQRG/mT3QBaGjDlI7U0bFkN2SeAsxdtg+Dqshf
uiZptHzQZUDpzS8OEC+nUUT59ecl3xIMjNGTucdglTTXwt8g4u6haYYXrTu2ssDn
j9iz41TikfhP5oKCo+yS7kQrYq8dnF28j+Tp943v6dMBv+XrzKp01w3/Awo2vLN7
ZFeNQERabYBlCoCnLatoDoAqoeK4L5tWjffYRZiNlz2bNeRG9KOG2VPkNrzadcgr
yi18MBVSNR1n20EfC4HZW3PqajjaavmIlSzWaX5g30hwQ97jHo3fC/2551+VUJY5
jSwivf1aOTbPFWnZ2OgEjCRtlUslPtGXOrdG503xUZQPdowAEsObN6EW3tURCKRz
qPq2TmCf6eq5PHvQ/9/ng7FhrzlNpxpFBIpbQVOYD/aPK5X/q0v8kl9NL0aae11a
uiGOLOGWYguVKtVnRf17WdxHvvBE/VAqocCMSip3F9O1Ka7bUN+Uw0zrvQu0j2pz
Iw9B/gGbSUbAIOUsNniQIHDAADJp+04njZr2AjfprbFMP1YqA+x1IFcQHU4j+F6d
+7J2pgSTTln29x1AHnCXyiL7f3+pVu3aLgjaULFgvfVqTME9snA5v7aOX6PeOdcK
tDiQy2vzlD3ifmMLVhFuSk93M3GcG0w+ABumhPVtCzHRwBQE3R+Nu4HXCDChm8Ok
DwbHQU8dtFv/kB3ko/8XL6mkgHMscza5KuHZqsCPEcpmLzuz9nLE564kyzXR+N8U
ttNbpTFaGglDT/XBY/yOkpSNMZOSZhB10Jk0JbV4nMz+70XOMRGgqd2ljXLi543l
+FMG0XE/xBC2u0VNsgUkltFq9rURAkVtLMPxYJkRZWdDfySCYNMMAbYGJ1VkemOh
JFzoUIqxQQSoz+6eAUo4ia56wEq1M93Z3osbO7xdG+ePxVrhFRrB4iZTJH6q/W4t
euxPtwHnchgH+yrYBqI5nxjyeSy38ZvGVzeGKWcrRo6+XScR6uIVYxHYeTe9vn3F
67ly/bWUwEyFkPisYx074/W7E5wp2EsZ9rVpzxXXyRqaDuvpjstl+VBBZ9gNQn9N
W8pMrjpDQXjjqWIyYQzMysuhILsbjWFI7stzwVa0Z9hbgMGAWxknvL0NwzIJu7Rr
r5dBsnLGtrpu+WhA2zKOiul6eNSu63FI+QjBDSdiC+O2zeGvjgUYCqEhpdeB0WjL
ZN26gYWRc7MEdcKfbkVCzXkaRWY0TIDUkaJbowdD+S99QUwDvEMuqjEvwo4UJv6I
Yz1ub2D4gNZAzgWK5ustFf5USJxR5B5zoX440xdB8yG6J3cTsRHojFTfFI+lOIKw
f+u1QKyGtI8J8r9a27QgsWuhYYQyC70BcUraf91ttB+99o2piWfVem/k4DE326T3
52X2vHx+LRT9Gyd9ENdN7orOIC1YcYhrA9uBGEJtvVF8Cu50MBNPoAmI/snI4ZZd
TQEedRnaijPfWBS+RXzLr2kY+2F9a6YQvUsm718Y+gelGLEOb/gx3TuuS7G85HBC
Y1aDkK2Ke5fUDA+9zFpEV7QdFsJ5ftW2nVUHj1XfVGJoeKi4YTjHqyj8jvaNpFA6
5J50O28uaVswfCMrp8xfKY+tk09dw9r9z9yesagNufWywsyrbhy5dc0nDV4mE7/J
bPlD/kpxelJudcnRsCNv9J1UAknUVrHBhNYkYH/hxlY2KcnzYEgzvmdSqozGn1sh
7Y02oFFyHjawmzygX4d+ZeGUBnDp1v0wCQRrZw1AGaIjemXmshc47a8q2EqwWTft
2Y2ioWuSNg46QcScyRCIxdsBJWH1X0DkoiJRa+ZOM4xXZDwqFzeYV8pU8YQzCw44
VesD6CWVVY96z9RlrCAl+SxIWANTA6yQ9+V1VASGod01G44lKZnse48GtLAND7mw
MId3hpOhjUSj9jMCv8WGwN0lVKsoXDV6ndVXm0O0aCeySlZ7XNiXpKboNCS0eKhZ
BuZ0teHVBRpLGFNVPuxwsrBeDYH5dQvNoqCS3umuQnbOr/cw98DmGiHp58RhvTYE
GK3rr8pMo6jJwEaqd+5FBk1pcSk7KPX2DW7938Ew6PewlW8NXTV+UTTrLq/odrN1
X7D5NS8/FMuboir2j1c3mbU6B2YINYeJ/BnlZVVP8UtiAExCFWPvTf6mRrQHOGqw
69isP22rWJu+ZOEzphdcLekDHkoDWZWvUrH41r4n9wihi+3iM6jjevGX/Cf/pET3
SFDNUZDidRB+MYnBQrfKeGh0X+/3dLhKU4WkBjAMhIk2Ru5Jyj21rByJVu4FsCwZ
0Qrlf6Cqn3utfXBQiOjgkSLzhuNwxJbSDmkarQ8T49eyx45w++2rkTrgMGQ007MJ
JDrsV3TXUA1+OCX637k2ArOq4s76SGiKpPb6/uEJ4/Hkqd9bkD7gEwk80XPuH1IR
JCrba0+m70naBaO/XnBpu9DtIvC2rTCwfBE1Jvh5nm2Azx4bIGUzJvU8ni25W4gW
kkvNibhXZq25RBfGVwjgP74NGSFErNcs0EhFSozvhU8y4pAWTnEuosxb7MUYpClN
uY6g0ZNrjOvAl0pvsBmC5LJWJBEdd+Vfeok1ijg5xCM5K/B/pvKvf7+se9ldoNSd
idAGMJAh/iw+o3EoM5AnmsRguepv51wHSo+UkdytV+6gh3DMJq3eVct6rKJxheqY
TD7fKhlrS4MO5MquF/RGbYyAKPtZu0acpp3Us/ExZorIJDVfBxFzBCwaA01pBTc3
Y8LuIFwX2wmIgr3jut4vV+qVhVVeJDEy28Rtz1/923A1QTDocSo/UVHGu8hFH7gR
hSmQx7O8aAPwrQfCrQNyNb43dWlzxB5Hvwtk1bnWkzQRDEPjzvpjZS3ho0XDS6vc
/viLSAceYzlQZWUSIpM5PjhFg6FUG1CJISvusdajOBOryfvSOPo9duaEIshYjA6O
OEfKKvzrbF8RJPoAF8tUYFbDXHASCglDpBjozmqJACn6QEOIuHjgxqwILUF2JamS
LSom3c1mpzPGEMHe/L8CrxgoL3f0O56EJRRJo8PEgX6WdLIC4C4Cmm8w9rWCf6MS
cgMM55OOtMKn+XDqu5R0EnMkYY/h8bjCW5bX53cv8Ij3bcyzFdci1F8TfVBxPK4C
yU5WZGrleuHRicM/jb3rdsjTmLl+eNEdnfvVJBAVvh0IccUBcnzQz0R4wJzyVc8y
JNgDISXBW4utmkURWx0ZNLrBHUVGH/a9hUGVDxC5jOQN2w0NvbFl8L6JMFvFT+7Y
5eHgtnk6WLcrqL2l9g1x/jpk8kb26r3E2fsZ8LcSQ4ZIMOrv0Nnjc2yMG72ybqXl
HMYC4eaq7tZw3r6NgCzc8EOoLC5C7inlcc2m9DpnpiGdN9APRTyKx4P42+0Rc6yf
nrvHJtE3GtXd4lxTs4/l0ytNrIcktqWDxg6xf1BmzbwadtpKqeqCX7LnkbydBgyk
E8y0//52IqQdnDSH6OvFQupFaiU6gycR2xu9iF+zUBr/l7x4y8etZdQ2rkQWOyjs
gcesxB+l4KFjMy8xngGpm4PhWejVYwIR8YnDAnwuqPriVCOT3gBluGh4Hsw5ia2B
m/suifsiR+WjvB6jQiTmf07vkIryz0kuByfpSgWhY0iia/eEFW4B9jwDB65+1HoU
5jTj+j+FifPW+SosxFsVcz97GwDrd7AfLcCAxQTn9yed0uZ1zik6CX2BZVEBftso
qE7er45wK3Sz/KXxR8AvJOwZr7cWx8AV9rlFKR5J+zbeKv0z0USZ+rLe9ZM5sGoq
DiwwgyCwjcr41L/rfCwe2VAw4bYcvHWVPCBqCXap4xJE/JGgpC68bzg2NtdSFf3Q
R6Vau49Uo+FUnwJvGjRLTgeCcFMtEpuJLSL/2X/6KaZrW/8QXF2uHPOZ+0qkyB1e
EOxoohlp9KZaDWIW9G+cr0cUnnFJ2Q4RHtfWQLlY5X1Y1WLsQ8/IZ5yskiq/1hEz
UDuu+cbP7rRyoHjLc3g59vm4n7HthNja8ZcPgE3MrgQZIAco/Z9GOV4rn+EbMfe5
GIDKGeGk+ynyeJ9ec0PBwTsj2oXTnoR/pOBIlX1sXDzlEXmZzov3AIyz5VyKgIOZ
WVXPcS3t0oCKEup4pRQg15RVr5KGz7uhX9xwFLRBGRwxF+kulmUIwve+J3gO1hPE
rT0sMUzQjsqKIRhfIt6PgCdBoSpMhZr2qwbhR5j6XLeBUCPwaGpoD/oDVIAnhcvw
mn0KFFqcYVx5wa+U5bHAsYGhfLnKu8hizE1Uo1OxG0lM38/K+Mpu4i2af4Hcwfhi
/hcJ5cnDWRUFgeJhsBU90EBkDnsSNbiDXElRDgu+78ZrJ+sHQrKapgJA0jlz3JWh
dNkWVYb8yYx8Ee2lyXdYRl/6zHEyrXpSiQ/CBjVt9RxbpPsM6BvNkxNC2wFAKv8u
VnDmc43kkiMEW9RAwxnS2Et38XDxrBMy9voXWsMQPbWYhklRxWWT5penknKxHDYp
PMm0TiqEX8yk2uQZ8F2j+goin4WciqB2jEDxGRI7K16MkQr3TZOZYIZYX3l8GSN5
c3P8mW95Qw6+mixMCdUTrfTR8vYARXwNep8f6CSv7AD68ZYzqYRcB2qYint+ZpoG
fl3E8cPqfN9AvX5PJ2LRXTkJPfHpjFYc301nCa82CAyxTEE7fcClZQmtHRDMBJgb
hSQ7dOdTK5+ZAWCrZxkpTLbzPPhcPevqoWmqdvUGm+aU2os5AdnGbgYFmerFITZR
URFMLX/khYD7WWsVDjjiN1Av7k6fcL5vJBZ1h5426mlv9ysqN2g/QYjrvukqX40Y
bkitO+2O6NAnGPm1ZNJpYQ==
`protect END_PROTECTED
