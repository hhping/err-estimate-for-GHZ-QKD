`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MEJl4XOoVC3joZDKMooewR7JqOPVXHikfV8PdEtA2Fxqbasl/v7/twjdmDVXqNMJ
+afjF7WF9E08ieu2jfzb9eUQzSX9iHI3ocxwE2i/F4xonKoirhc+CanfpI/26pjA
CJO0OomzZsvEv/Fxk+dkh7dUctt630AP1EKK8nFkeU3IqLOf1YqXterTH/2mU7to
9Fy4Omp2bG1Ato590v5mQwkw+zk2JQHkFAFVrjPUbBAztN757U5wxnIUT5yDGMAy
+27jL3ya7Mht6XoQ+nmLGCLP9o5NvdI+1CJieThJQRBizvQjG2mnBff+ydUM7Gwu
Sdyuv5AurS4ftJh06sk3tyPnSfW1bKHdripTA0m8nSUDGhX4+j173oRgCrRBsW66
JMEGN6DI4chFH2gY2dlnIVg0wQdR/147N8qIQ4mJk45AatIcG6iIJMynRdydzJuD
OzGZS90YrAmTU1Kq3G2DM35rXO5USTGnC4YSnoUKFztwuNVR4lT0JuFoDPj0XdBn
UulsHSAz7qFjD8SbXw/mcTEqkQbBUGahVHjdwx+GbQZ4UluKR0bZRJ44D1r6Ocq5
ylQeSogXUfnUx86DYNoyNZqzrV4LqW+y/Htn1ysrVi05Qj+MaGapLbXqgSl6CJO1
GXYPg6qkbrdb0ee3gBXxZgWP+mwXU8US3gSSJGBK06PoOvMLJ4nJJfmNFh4OpA1L
NAjKwlV7BPpAiCHmGV0WZk0a3qoES5koWO19tU+Y7B6Vg2jXKjI4wuAe7MggyWu6
6MB2wEmn0/L6pRUBaOE/mtVxr8YNU8gPuB5BrJ9NAOr58mbmkkZYvxmRcGpHYERX
xYEz1q9wQL1CloJnxuCiSA==
`protect END_PROTECTED
