`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46q05OkSUXA99zHInKtvGGq7O9IEFdMy6Nw7hHS4iT9LHsoIFjJoOmrM7lD9Z2BH
qn1wDHH990l1UQMm/YdAlRid5qsuowO/uhxo5wA/bb7w+TbuCHC80Nw+Pf0eJB4g
u4JQdH1cs6mEJiPbzu3Lddn9sqii8nfd25GqHmYYOX0dG45Pk5HTOz35bwGBm/b6
g3Cqga1tAs19HwOhXl3NUFgOgP0Iv+DDFaQOFeHkbP1W5mxp9Dksy2FEEFpBWw48
lqyukCJG/RQi1NKNrWu0SWyj2bBW+vCr5m/GGzU4RK1AVfgX0xCn9Yqkvyc+CdPT
a5Xzrqg/u68lk6bx6LBOlP6FLV0RjjqpfN4nSCYE8TodDA1Bbjq9uPSz6NxNPnq7
tCr0JwVELYHxpl1JRC1ADWrAGVw3FFisTAcopRQ6rMXTjL4A/BteM8kszHuFmWNI
8qVJWFw4JKv0w/vh9QtWQsphZvOHgSChEYSsIQL437mzKSsEQRIF7yJaR3veY564
SAfJ4TFgDPk47BuEJlX1eADegMr01koU5uUVyjU3WRKAzxX4W1pOkCDf2CwFiUdc
+putJeJBzxuYJXoE/PTzOZ8910ChcLTTPvB5r0ndQNtqp84mkXfur4QA5Jj4W9gz
KBX4MAJ6KeF3krd0247+rNqJpBAAro5dwcTVLf4mqwNcU+kv7GhnOG6Bx04ZydDh
rUbRfDndgi31JHVCwfyJB7S+qgcGgbyY0AiQtwbHowXXzhNrvjdWjx5dKcBb4MNF
grLONWFmh/LcUt9EJJEXrPRybLYew80wCnXY+vEK5gOvz2zI4k1Ww49IQJ3Qh1Ba
UAFN6wnR7eY6E4rEVQlbBry/53KG35v7fDIq64McE8RL5IwzKm6haKGkI7G4Vnc3
K13sX9oAXoD02gSfQ+Tsyr7SuFIzjO9xrAyOxKmrYYHjs1O+cKrLMTg6k5JP9+Hc
zZQqwAJaYtHAwdJllw/lwUtzV42trNUyNvRBxgMNzA1YRwBNkNMhX9K7h1hli9ZV
HjSipACtK0bec3UviFFNuplw83ouqljyac9QZeDnPw3goDu8OTlLPvAX+ImPW4i9
k6aKKhoge4rUloT5lV3xsoOpsHbI1kiE2SNM9hgv691OBPFFGSVqFraXEnSgCGTd
2B08jrrAxHSWFWXDdU2gG1Q1WL8yBQI3q1REkefgJfiR/WPbbmwEJz9tmYW+LZlR
xc8n8B8J1LsNvQrui3OwUqc/cbAmuwqWQCpLeySBfRGRZpn0us1Kvw6dQZ9sVSlz
ww6iGOnszV1mHRUQEMKha8as+rO+ImPArYlY1LnbV0qD8wUWjuvJrfCn+RyVKQ9B
zKddZ7Uq+Y9acYjWbGcWTDoFXREJAnTk13BefBky1Qqg2OkhZTrfBfszzip59NyA
7IKwEgBEtoAg5kx3MIm+O26sLTHn54ZGoQilo7oxAjUiH0hCGFx8kD1+DxsdUf6H
2f4aOzdQavw7yfgfpXfVuUvObuzdbt1H7sUNmMynZU+x+u/RbhQoiZDtQu2APrj/
1BZzNb19S+nQOKJQDGj0pnyza3Di/MNhc7aqK/f0rqiQEq1l2BYGoaBMpkwLWeu0
KNWN9VudiDRYgXjKE23pyki/PEfiuOevIGveUhMUt3KScsRP3MmDlW44SH8Qc+KH
2M96c/3x4Arfwdd51dh84SdDLALfKwKdYKT95zdbaONacx0wRVLSa7kKjhXJA50y
14jwaD3vGSomELv+IJpUy18AfwnbJYoNzgLoFbB8ltJSUcQrRz8WUunNIP9ghTA6
A9at2g8WY5MkFsFpMtupoFA00PfqbdOp8RjUhRo6WVUs9n7H0nom0pCMBCSRy7JV
rNVQ0ePIgYHR25nNh1b2tD3B/6BFB/VjALolmHun0FufEk8HtX2CAV7PCPjnLz4O
eYnmfq7PZFooaQpwGxQHw63/WploYQWejkE4rCCo7J7oW6sRT8E7DyPp0EHYjary
uFlKgdIc4l+EPhwwV+QZp4TqQZpK5HM34oGUyrk4dRB9KTnXucX2Kb2QP20MZimZ
oRstm1p5Okkntg1t7HIoWYiEbOOVig4gehcuwlUhal4SsBRJCwAFx0AiNWuLSW9L
FTwiruY00gl0+5opTkvNmTIknMN7KJvr59VYcju1dTr7mL1Shci7wyFzF6hi4N6B
u21iO35P5lZlKQSKFFtNWJNRtP1Zl9CEDJKqxtfZGQKMVimW9VuwADe5NDpvQosO
q8jdFwIVGaLsQEhUj3LrfDNhSatLGE+AOfZNBhYm7KXb5X+srq/DSLbYVOcTcDVZ
EgQT5mD0ggI1/e7yLHmk/ybiUUbqCwQN4kXrKLt3l1tgrj8MjQpea/LyFBxm1b35
uO/sVs6XcrnxWTQZ3tO4h9Bf2ntp1aHSlhA7iZ1NqmT/io3suGPppvqv0Krxn/wY
ReOiVdsY6uIsrz2qRodyj5XlJe646Thzo6sWv3E5wmoxKzzZRVDpDbB65NQ+RBmI
w4xhxZRChOFXU1ZRJIjhCBY6QveQo83IXrKRwgYZ4MzPi+D4wsl8afYK8C+iGz6Z
HmGcNMGCrsJ3x4+A0JpPd8OFhRYDvfZphi7qP4xWkigA5+8VMVpr1k4q05ywj1w6
76Gm4P1vFE1NXW9UYR150FtHxbwXeP+AXYlyjRQ5LoQgQyQZBIkOf9nOc9Q+Ovir
y3X0GHmT3SrJn4cXu3u8KrrmIqibQ6GHo7AU+4SK+NizbksK1C14v4OKBMbVRjpW
Tzb7K7QGLuxvnjCcJB1ljQD4qctEqMklhu8ru6Sp5PxpSVDmCF1zBZ5eMqdYjpaY
2a8mshI6Apsv63XIji5fGHHx3AtY5iRCb4vVdpQfSO0UpwK75cnBbEwQqSeuu2H0
rae4WXuRL5b1nWvpg/4jDYyNmizDzHjkx2DvwAUkPKU7kNBlotdsMMEKA6Lk10ii
igfTiyXPvMLx8YvzUCHpGT+TatavEH2qAcqrEvcCHi4RYss3ECCIhxmKhbctNpR1
2rhYSNFFBYMBSJsJ0W3RVdZtevL33PO/xCPKzyyTgpPwz1SYVR3gkIvLks/EU5tO
0szDMFeR3OEVjaxJUbgQLOaXfhYvtVaRUUKoKQ1lXofPoNfx+qFEG0iCFd0cMA3D
uNkcnO6xEbNKmjjGQ5fPkyjK369xccs3S8kUxAnNfqU/U0pSPDg8Z5bd6la8ZUrv
zG0Tf85XR/vTrNPG4LLdCDGW3e9ADTNHvWWtO3mCZLCpJfGro/YMEVOngVcJ/Ah/
aJqz3/EjRMbBONmlLi6AQewkJAlsYUCyamdT57CFmY9xYRA7Qv+XMr5yzhXqc2pR
YcIf9WGrfa8K4Ow0MUf9vxChLJ3Ax2gSJbFXM6p++Ts+TyxSWRgrovjVkiNb9Pra
DTAMUN+6/5XbIVFo4a7NW7rBOnRlGkJSZarl+tLMJ3p1LridkQtHiLc9EPg2kROs
ZJzZooKY6IIudPKM4zwGKJ4MyLaJOBWlJ4sxSCoGarDFv6jG7dcYjxM+zCvQMqcr
2E8b8jQo+MUT8TAkIjTuVhsnngJpB/zCKNF/8Bm3/7s/T4l0sb7A2sivOvz8N1lX
6vvTUDxfCisdQZfMK9BHfTCQ6GdiPnrlRJx5BRwgpR3nWJbcolswSNJwuB0XcLqU
VuOOmRynIfvMQVirePtrk9nCeu47jezqFNep7beUSYalhOLTS8lU7yOQoFxOyK6o
rQk5+Hfwk30T9lafIlhKAS6R+3/F6XHp6ogtZp6pdgeQBgHEdhWplB4e0L3sm2lG
n66tdX4s8D45DwtlQMv4+aaPnDaMSR7N/Omua5k8baud2EVxpoLiJyml/OFozN63
vVvwjYcM+6JmvIdU4acgrJUbQDp2gzMNCi1INJj2L+awBnNJIZs/IpsKgv4u4Gw9
+cVEuw2566b2essL5SL8ngaHRVGp+VwmvV12DcpDcRL/itGcIZucsn6AXN3A/Fqh
VzArbPTrbe0uNuy0s4zFN1H+CjsICtmA1mmLrpZ3zmqQWFyRKwHjUgi+sNuxy/Zn
0C5fVf2jfCzCLVnX/p3LMoNDcuERDnJ4knpV+b3C8DGYgKDeBdPMxybSHlEsxsWI
hYQYNZvIQbfUZLxZT0GviIU0k6Gq3qdJSpjKP2hYyLtmFl/zaHXxEFqNWfW1Hmqe
jfuJ2Hu/uhPEK0gRU5A6B8Lx/oe75NG6bcgtK42mYrQVdHVi/N0w26aJ9cUQxUSc
UQpRvEzRgkhPUV3jn1eDyUfjieyiPBeuw+agCwWtJ4xpWPTkKiQo03xxR2g14YiL
RoLY7Prp6vmSbOc5iqoQNUEnjhWIeFqfJM4NmZHty8cm+oz2Lon8GTod6qLSSuRb
Q8sAkZYAOuDM0UF/bep0p3cAh0S+8TgZLi+LmP98xldtYPrQlxt3Rx4rTJmYffSI
22OQGC7xM062jNvu0e13y0gdeOrNT2H/Z/rQrC0h5QUizGDNERrz1EfQssBw87ZV
P5ConAZG/e+2cOyK+nBpy7/DAR5/XvKJy/4MFa5BB0kLz3NetkSblUsQV0zcrG8R
S/uAy552Q3FMoGkXYrorwEc2zCGw1LXAnvXA/uk5nZKDOaxsn1FfWzZnWILIJZ15
A+imkHlKb0Js7ixOI5sJPHtQlGLC/gs3LI9y/QLSNTX3DKLJ3S9cjb+A5bO6gkDc
g7NynQ1G1i28kZwx8LV0bbZjJwjuBQWfEJZATcP2gWIukAx8QeWIERJIXyonL6yF
6kKh1JyEGAAuPOXJk9Z4HhluI6L7YfVdiAxuwEOm+rf+EIykFT4HATfoFytyOs6E
/J5a+7HjyTDiV3LC2B9vQTn+FaeMtQcvwZiWPG0M9idxcLBaXavCWHTgcPqxFmuk
nCHLPcGMqx0Jjft1GoN7U1qMOfzFTcYsPDKnZoHc8+V6QKMl7r/LaubS0IXWqnIg
gA3+p8cRvJX2s+qS5P2cpaWORWVrnC2AbV2DcAqRrPhI0BBakQfYTOG2JMTKUER0
qpAJ1ELpiPKrDPcoZeKrye5RlV/lErMoE8tSwz7gZDYgoUJ/Qk28AvnyAKn9VQ6S
475yc5+WfIXqrIFUVfoD2yJ334QZyrQjzfMKaNsn9lKLYJv5YcrBRwFSCYER4QfX
cV3ALQBKGzXTuG4Ne8tl/Tst6BM9yzjkb2cfEu6fF9jyO2fDlQkVXZ9UO3Ta99Vw
JjruNJybXhYRsu4MEb6/GlMpo9//pTkcmWZKkFrB1c6NyQG0z/mKGRjoyOeT6Uqq
nqgUY5huCOVMPZRLGoMEMidY3Y6yaqcS4mT514QM0YmQGk4d2EnAt/xj0p+MJMZ4
RxZqZp9B1fRynyNNbljraJx4V4HJX3bl9emAXuHL5HB+vCrGYd+EIEgQI2ipfXqu
DakS5g9M07LXA53RjIgJWejqDrkxC8n+SHh8XD5Eb+q3LrYKcxVzVdi8r9YOf1Xl
n4sS+imR5SgtBr6z8d83FlujNGgppgXadWL7v9Dm+ZmdlT8QmPxj+Pu7m9noA39K
6OMdh+mTk9mSpSdYeW1ACsqlY7m/QsXRFIuGAIEQSE5IOSgNUKcVZSfRq07P/pdw
akNYmckEo7r7/TnMlMf0psqSt8F4f2nmPP5jQ66D84M9KZBYGym+wEDU92+jURr+
1jCycqSCWAnAP418yZdlHcml538jqiSt243/LKJNJk+jpKCLA5wUtHar0u+7/k7s
Wm9fj4sMHQt8a+6bNCLXDZ8ejS+ouqtSdrOfqUZe5HLBiD+L4jQ/2DY9DofAm+E6
SowBsmDor+K6aT6FnGvRhTNdfLa/vg25Ahd4D2I29XcVry80u2OmctaP6mKl3ZII
xDXMn7slEdSMUraqznUY/jSMvHkwROJs8EEdZkTfd7VPHr+8PNzgL5RkPjeuATa9
DoXJA0beA6HILcrgJLRn6UH2Uh8jnGnN8clffMqigDA7cyC/L5Bs5qM1W+YCdB+U
1unWOk2XUZym69ogZaLLIhMjloQy4fq0KlFQg1RVb4qtl/lx4HYUPAK4ycdCwx45
9Qw+Igcxm6SN2vWXEg2MBg+HQcyMpOVjd6zfuFxiXtew/pqmzK762cCJKnndzg3z
YdV5VjEjEo++VR0cJmeYveUYrP/xTwImd4Fk5OtpBnjCF44N7q2INMRxIT0TuuHD
tCS/inIOnd7nKEX6NDyutm6g2vze0DznVc2H68Umjqyg6BzNuy/HRWtcxPV9pVMv
QiQaBUfXw0eSzV3YhGUoAIbrX+IqtwbXRNTPELVUVu1BORC1RLc/4LslYx/x/14f
p93khU6OJ88haWLh79K4vwvfzaxYsNZDyVrhlAx0AL+Xl+JcCz2iNONCyuhhV93j
GpH9bn8FUPINYo/5J9p6Pbshj4BtZwXSY3SfwEisKJh08f4o/G/Vt+tc5L9Bic2t
tE9ORnPLdeaO9rq/mcp1YqmwprOrKFtdthGy4Za5EFGBiwP0/9HhxPPz7LQA/pkK
NYvJKKrqPkL92SgdnbNrOtMxMX6yknmdBZGAoCk/2+ADJ/M9MCNIeCI7JoMhgR2+
RZlfANoPQM0wvpNXVHDS1Y9nK+PdBgndo3IKQKmSsCnwl+hLFk9XexwgTB7U3sY1
XMXWU5JiI16XSWM0ZUUQIHhau79Ofy5t8KX0WlEbKqYZwbZUaSKSs2nm5lAM7CF3
/C8L9mhylZLOTHtKL+Rl1aRZop+dxWUu0Zmj+Rp2SVVVXth9pCQy2Gql7THrapML
bf3QG48rnTQNqc/UvVJenfMTU68QNoVTalhOfiSrzVpdusmpzzLzpWIszMPXsY9D
+3dpmP5WiPslJbyqlMlDJib9THLO1NmGqwDJlw/T9CBycVjbSdA5lh0vCSKkCJRb
woJYGOPx3eqiWECel+ekPg8/zmk8XZRa3YZYG4FzKabbwW7Emy9NJb84rWEQROoB
1jWFfD2tU8XWRvlfaXBsWo3T3q6MStPpe90L9RfrzomNE8j65MaVSWEtiDJSnLQS
CAMLwKKcUrmG9i0paq2Oy8qLyTb972C8fmtj+sywtZOPg1wWyBfd4wYbtwuD9KM/
qnkg4/0BA8MAIyWFH+Lty1MWm0JM3yQwLdgosICmT0rARN1JSKdF6iIVYQHWxH+e
2cNslj055ots56zKAIzMpfi2Q9LcaIvous15jHB1USlxtpt+L/xkXfCJoaMR1W+G
XvdFgSsQU42sm47rvbHt1cbNlrN52ooQtJ6Be88vHn+wU2lY4iNQ03L2Ixr2jIj5
jVnZAA2tZwu26eh0ymlPoBrAzhxEaRcG9WjtfB3O/wjeuMo7v2q4NUCDjvZ1NnxI
tNVGYsEdgi1VEiXbwNeGFqKZBoiwpoQM8gU/mt97wP9Q3ji38BeUjYbVO/NJANGg
8BSWimLhE4z4IMhC6yA7HgyJgz0IEytgeP06Kx+zxJvY9mqiNYkedGLjXgoCbbjW
FECAaabObVkUsYjGB6jE6p5zoP19DKHynxKLavnnzGzkW5Q2okl9KrUQUWguUqwc
OhkQjBcVTfrtyMBIRYn4ZR1V2iPHvucDve/FZ0Ti7sxKW2LIJ3iqlZZIAIWsLaqW
QTFrrFya47ugO5LDCIrTo2fS+IIOe5OU0k9YpDWoEKGCc1cPtDfkAWyDItNSQTHV
QZNv+I8Rq2986uOenKi+Sdjn6KXbl91kDtM1xJX4EpvaZDWliw9oHuHWj4wX29qG
weLom6V5uB3Xqb4S5nuD8GoRXvVm74OM5jtfkQGQCd3kf1M/jkCexq6VLzWkOd1C
JA1EGG0Uu/jKOi8Hjv3FeNu9qtT3hrsXh9jm/oKtsrr/wQ1uqvzLQEDaAeOAo3EN
QtuFASgMpgvmkYwhXNR0fjBlNerdEGi6ZCor0zXSOv53INIW165iZWcu6nUiRfnj
IddGr8YTf9eOBFrQuG8oo03uS+TrZ707WWL1khTrsZS9GltgaCMKWtoSpujsB5al
KyN4We35rUT8rdhhJfC/ppP3UkJeErh6MK5b5s2zbSx01bWJPyOXXiWu1qq2vms8
VlyFdP1xPOxFB4I5fdkXNqkk9m9EKADq7jTuT1mfLIRNz15fD/hi64YLIN6XPNEE
rI6YmsFExn7ZKlDpuItf3zhRWkQgnL9S4PGUUPuJ8Ho5GydVoIFcbyWa0AC+sSBZ
wX2DtPV76o9K53Jb9BXaVVJ+wpJR5Pf/wWxMBVtNlmkoluOp9ZeJDDisdmTknGtd
PtQ14FyjGCmGGlj7/z5H2WFcJ9aVDDmGUA0mFFrYrnEykiRhI4THJ+N/4mTz/pSm
Roh3bsXOW49vDQSAmRQZ1jza5gL2dH+cs5QEB2K5ck9jgxm7/1wUIc0kdMoRLZmW
ovkaedqi7/QIE4gd0wbv2HRs9/oXpB4afggiqPPj3wJZjtHqTK6Oxikah9wbJLIC
Nbans+AnHqMS5h383eryE6ks42QaXOrwVpnNDX34KJ5Mz2W6nXrC/tU28HxAYnmS
pXHzPLSHx9Kf5sSBVWcTkSolh8Oo5+B/UfX/MNo+1QFN7thXjdhMt87sYkauup6Q
R85nrm8m349iDE+dT+AvorvSiPTyLRnhTtSiWdX0FJXce/v0Lzy6MA83HnTdYPdz
oWuHwYeuNtP67dKcUjxa0y/kxuQUPWrMLAaIhSef3uD+YvXvQozb/ko09izyXmc4
/rQ5FMNlGBPPBqQPHcdaAZvxyr53bTB1PJF3xtLtjBpvJ26P3nmgL0px2QZEwe5F
za1FDOecrOwJg1KzlcXmMAVLaKA5YEzKvnTJGfp/Fkt51gvGeHNnhbHEgo8yMrrh
HWOeGoB5G0BuiMUaj0BN/xuksr5DA3FSFRriKE85T3i0i76bL8xvao6uvVBwVr3/
YuPev5DGujvXmCXpitDR/pV0OxSsCXhMugrTOv4rOnHozDDj2u9Ldhs2eV+O6J92
Kvy0g+GtMiHjwyeJqOiDkqv7DkL6YYrXxDc/IxaQiXOoXSED+WcIhBxwACvuWPQ2
5h8VNLQQetgSDMbfLb+7ero+2PiKK6Ku68J1SVcCyv5I/6FxWkeHA8w3t7txCPm3
Ii2W/CMPSYURBEmxM4Dy1ZEIMI4qZG0wpVl5cAKB0Ezs2WxFvdTrckbr0NGh9fjH
3RKkYklaXmxwHCqEBukNNgzckq7JI/8YGWmKjJJzZzDT9CQhEWNur4H/uKo3ySrE
tpTMFG+3BX0EzkdHvZi9BZyjD/9LeSX7xzjRfKo1naOo3LcxZ0XHm0CYKrjtljYH
1OY0FeuTprBFJrQmb6omruUa/eB1sI+D+ji/mRjDIN95Pzg62zE3PnKgmVmG+Ma1
iQvR6oeVouLWSjWg+2D2r7Zg+Ad4She8v5es3kGu5yjK8aZUg0scJrjdFw4rESjz
9EhmYw08R4pON1eCXH2RULzXPh0bNpJjYXwzIdpdrjmdWL0BlU+X8Uwn8PWAx5Ur
EOi2cYYOm5uwFVkL325ykHKnYKJz0+OFTmTJG7dmw1uw9AK1S9M4gwoiXi1UKBWG
aciDzG56gLwXg88OEu0MZjrbQbNi/dyyPN6hw1/ZvaQqI9v8sRv2C8Ye1TrLZJVf
k0KrnQPHUhD8Z37HRjMAeSgDzFxy1UPxZiuKyiOJX5yXQ7bZJsDUoq5hK9Rv1c9R
WHiH/vx91pt72JAI2y46Au5U1QfkTaucTqch0+WFESj5fEDa/OUDIcCNIQ9r9fw6
6vJKPVhrk/RWL+XdRqJ+j6EgmA4eV01xjhydpkGU4ycaN7zdB2RwNRzz1DOhfUbH
asHJj+yztTbFAyyygeKDkhltM+q1DOG67+VXIErLolxVanx8a4G+9Uy0/ZjX1vBZ
bCfO/D9hPS593EW1xVpT2qh54g1M2jRxJQuGs456o4Ze/jiYqLzFKANbjK2EYAJX
V23Vm/RRSWhC3hSG/o4QRSJ7XjBbU1sC0PwpvfwI1wiW6MeEjMQitets4MnMK0ZC
iSS7KH7ZcUZ7FpAwpzZXOcQXhvLXmFHZelTOkbdYTGWtUoamXdpJmTu/pfIE4NTU
WxRHvUCjC6rEKt9urWXYSvnVS0N7k2KOaw1XyOS4B3vBuaZ5/iKGzRJox4NOnQS6
QZwMfbDtgLWERGmKCGOkDJQTtwAHmHlXTg+cspak8L2Xx2tlbE5xBfBI+tI0FVTe
/Z8fX3wTpg9T/cmKnhvghaAIZ4fAx0xlbCZCffdNJDx8GSarF4T9TBfojgnRN2rq
JOwX6cfv6tv+4g0xPT6FKY+T/i3fwreBlp1BO2QAMoS9FN5BQOvwh3wvUJi3xVrb
th9r61xACgF+Swvb1DikOqpjNIDdN7z/V1n9deh/nK5qhgbqwBjfqEEFuFi67qWb
+ZPBk8Pm1BBSczP39YvjTHIp3WIKPjjFXTXSYI8jQjFlwiglrd97LadiZrNljD0q
fCX2yEGcmIJ/10JNAI5CHCE2F0Bs3tkgFbWIM+EC3xEFsxlUJ9MF/uQv6T3czHI9
3RlGPOJkouOAGG30O4+b9vKwRljPGBleSoqCfLhjOhBwuz261WXT8QL8GafAz7bi
omqUKxAj9w9ITnDOh7d73c1oe0QYGtqERzv+OVpicddGdt5EzCPMKMhoRxuMLXfE
e2Fvxr8fCreartAkHkRngqJ3d15NdvXhRRcY5AMIIjDmUXg2NqhUS/KeDVpYVRqn
j5rfbkA5hOJR8MFawQfvs6bbSbRXVAKY1vfiNNGgbtjCqwl8lR3rBkgkPdb8LYSw
EFCAkqwzlRYSP1xBlOCTqhJAGSWYtWAc5eEMeDQk51D2ao1QO2mSY0Jgc+B1Y3hv
fcM2AdaNMmAeXiTXhwRUUoNC6otv8aSxrkF++bT9MR/4yjhAgjpxZ4eKHI0ZogDs
iCWDQnkG0bXKtktGWz4bwYrjhJBhoW0dFKgX2VS96WMgacheoAD6jSyp+WXeGYKV
qvD5avKfPz5Howryr+5MUrsgahf5EZViSQAEFDN9au2ajnSYXKmoOOXPXZbPTbbx
HKreyDBx42qhWbbnuhQuRw9A8HancDv6gQpWueispuJ2jQ/TRvMVTnFPe4qPZX6i
JwCf20JAgXPVxLmViqUZnOskLBqxChSI39G/XOQxB/h40q3IVtEyzZiO2l2G6I1b
V++2ZR6BgOIhJGEGkgV7emrj3Le5AxOYgo1sXdM7XZ8SHw/CUtbH8HTflRufQhQ+
DZG0N1NqZEsrOxAEDGnVQJGTaBWDH1Pn28ty/TNUekeO9q7Oj7NW8wCJkPvaa4Lo
VxYUyoa5ZqgM053/P4DaQpJ73AXsy5yPINs4poE063+KqlDVF9C+ziYJ6pCrIJYO
V0SvNPsw14r7bucA6qAioMXmBKvfKx5c/0BPo1+yycqkZbIqept00ZppOEZEzkjo
DVEDeOtSZeF1OGeRwnyP06fUtFLRvpV+hwGqp1VyaafaYu2phluuYgQVFd18QKcD
mZo/5glQLqkyVEE1zJG73LFj03ttEEXnlZMKCAGSizCG//ncANEE+mp0a3nOg3S7
2qIBsZODW4Wc0tqdaWhrvTuM6WKAbug0n7L0PDjLSb7bs0jysNdt5NB+XL37s6wo
4DQvJeFf50alG5G9svplFodtJMTW1ewu7XON26sYkuaJj9AxPbqMR4Gv2Z7urRqo
t1asLKww/hslLxxzrdti6VlnmozuyknWUXv6dbQNyY+rPPnQVMzSIZ75M0EpeuHI
/zwhXqU3vYRh+UK16h5Sg88U5n3C8J41k9R/09jNpW8LvJ+5nj8f0BgqPwB/LX+A
Y2/qrn2v9A+4h/baFd96p4/z3EYcqnjPTTzKbCWRlisAjRsvkmvVXmjsmAZDRew3
xqEJnw6g+9oO8ARTGpAwoBeqPpeLupaP7LW5P8iCsfPuFE+lGY3dM8sI0BzkGtVF
OdTmX2JGO+We59LkKkNEOUuex7R5vyu2vjojZdZ55q1jjI3Jb27BJa+29uxlvn2V
xNVgbEWTxPO2xETzYEzi1c+oikGBvf30QENtJ1/lOzQcoJLJcWihmpdpeJTsYL9p
O/vb4F6RV25zrP+n2M54yLQEZe0DbGEjlSX728ed+nmuRxBi7NKIUH6ITLPOxl4C
XrD5Q2UvrqG0wUaQ1PacZ3wEyPV9YT03uJ7pX12sBVqR259aQF6kWnoXXtIQ6y86
5HnlfKFg24cQhL3KxlqqDJ7GQvsvyi0lLW04PBvi00uLRWpCM6TL41GJ8xbRm5i8
ETwuEgycrjP9AmgReLomL3pkgRyXz9dSiEBSFMrdEAgqIeEd09X4CygSSOvswZ5W
N8YpkcK8CcNofuRaLZVEBK36GQgSUTN/BtKdzCUdbG2ld6wXc3jAiO7ApxcCmDPf
RWHddhinZVaBAQALsNYq7SeiLR9ZLNt1VmhPGQGPGX5uR4Ne6UnfeffnqPoVVeeJ
xWiFcbGC2NpDkx8LikHh/e+FKlhClrkC5ZSF99Udq2eR7+Eos4RMsayB6JZNmAw7
Ps46fpezQTETx3quf0dhCT7txNK86J7zsgQuYxhqi+CHmovkqmxTde/A/UUkKvGW
g6ChWEo6Yblh86s7Vj1uWxW/nq+QBuZEezTbStDYskLcC9eIPbopSJaSIWceCyuh
AJZh0Nk5KS009bXrX6lX5XJTu9+t6dZqVLsvYQSiVOWDVpFXGDkbw+EjwLb0p1zk
6T58XAw3GvV/yNT+GEoCN6gTeYRe5vtvZJAhFbkGH31K6UDcUgBXaRNKYfEp10Sg
Eflo+7b2A7eqJu52OJBQWe2rlIcPTGi5cUjjuviXwcusZZz40YJ1yIIiYNRxVkP8
tL0le7X9gcChVTbXHajIhGeLhS5EAzCqfROmToqr0Yobt/M2p2/pTR/pyaow2q2p
BHDZFk0eQfuuzoHqesEcl277OaOZoNeqUtVUHGVWDTFnbNm0hmMrOGNe5yVfs8rS
nJNsSK7/nefMPO+8Dr794pkaxPdjP+f5y+Pd+5TQNlTUvMeMaLwHN7hanIY3QnLi
PmLmd1fJevmLG5uzmG4wEdniH93mEMrHxZc6LBMFgOMS/Rv9QdjcmW7MgLgRBXQi
t4gCjs7WZXuiBo/jefVME3LpDBspJtH+uqHXZFpknrw992g6C6eZ1v8lqech7EYv
dUPlJgkVvOwDfP3mBzY1N026/6ZBUyowSiGXHSk2vDvPwAzTN6HukLXsU8oR+iYA
YYCg3N1UwQOB2Z5JFkT5nbsy1YTrWfoWaCNe5HWboAs4Z3Ai0pNBEARmyxhUTaos
oR2RR3Mp7RbEzGbw85DhhbAZ0vigYf8rLR116u2IDv7HUq6nF5pO8IhXM6begwJr
vdUMM+VvuU3E8mbqJB4KC8g99zs6qmWbfIk4/hCHJmgiT6HJcfUF6qXW4ZDJoJi2
y/jViJQfe79GvY8z//xGKXXlKYISjKE/d/z9QvLKp/ByD9fS2zOF2867piv5ZDQV
iw3mj0kr/9wCBfu4ynQ1FzGXSr9VN44j1SdBl5tJwky9KSpH+GcdO5RwksKa5pqZ
1A28IEDxYnZkhsS7AjbAfCIYRKv9R2++byRF5RzuKTYQSIklewF2YNWie7eMMz+x
mws/zZJk/Mzgh/Ei2PK8cVZkHMAR30uVKCX6NFufXZWRTracGFPZZ1hDDzpC7RZq
g1roY949cjosvJ+DDa2Wv2MKVxJEdshvubPQtRPFsemukwEkshz0UvdBHUs4BKFW
aQ0JP0TDkZc11kZs1mPY9xLlsDlF50RaHBjusNWs8vK+tsAa/3rJR42ZgEp4NkCx
R7bPEfEUQkqxs6tViVE0hm/UtVF3FPl9fD8AJyaMrHrKrCt1c0T2WJU2pD3s4r6+
1akbcVV/iTtOdqOHII9fQ4VL/V9zAFzOlAbm8voD9jw2qPtKr6TMEJxM+/KU4AWk
LFprwC8JYdcYgQ5lUdUYWTA2RXFmSKEdH4BbrgZfGIJ198C66GUfR+6ilU/UJWVz
b9i5cYn27mTkrbIpGmiXQFxBQwURrQ2+W/AjZzoNdi2f0DzN1IyoHl7QwIiJHbGo
Vdbhtbkw3BKxF6s/2aOsMj2yah6lIuO06+BaoAw3LlYza1ojw4YORQ4dkZVsekCs
0LYNfr0LdE/kprrei9E86F0Gxmdo9xVQOEnjHEZ/Z5/ZLOQjdjpm89Zxo/k8nuCN
UMFXLbjFP7G50p8Vy95UA2DsEd/cxF+VlPYAScyIyljUnWACEch2IPLcA4lrzFwr
/9fQTMQedhSdHQ9PWBeeXbABKHEwOOaVuvZsJuNHDamKDzsFsic8GqU8zbSZyBEl
rYgq89bKC0fgvQFDIuQlpNjg8Z0WbuJYw5XmdUjqjMBwi8vWqdxHP6UTfusjBSn/
aisNpeHCAOyuu4fRMLT5QXa/IOnpCatGmrcQaOxxpQsXKrQe32gukAZLbz6omyut
jRNmajDxvRNHO7gCgO40K7acL+EQDSR9P75gx0WWgsBY32C76cs16zGYDY3+m/Zj
43TmQq9tiDdMXKfhVkEwrUSg3guT7hES59HeisjivKuqaXya4gZTj5X39Mvgbv3c
Mf8/BvxbSDiLzH8+QOzSjzQVQqcvRWG6NzEsxwPtNdDtrq+9ttPTlJio+8S1zYHf
cCPWMoqadRfwadm/YJQDo/H6PwHdf5EAdn/J6OWCDNeoKslI8IC6IFbFT8rzcC0y
CgXnT8S9L4UbHRX4bW0BEDxU+d/IqRmqln89tz6532oP5klQZzrLH7rsP9Xus2J+
4jcAUqDATPoBSf56fUWS0bda+Q0Lak8FmWhWRQrDVcXUWxaGbbVlD8cWJQTyvv9x
JhQ2p7cSzCoQWUgrEPOsiMXIRkLk521z6ObiNrqnL1HxmVervesQP+55mQYIVlFq
aT7IgT/J28kU4U3ySDwKEiQzVFdAprE/nbfEF5ajOdtZnIv0ikRV5QrD+AePcmsh
6gPPd1IcYwIU90JQ5VvVjSkwBkqXFYP4neZ5K6GUieBtONLKgi4Q9Kc4i/VM3kQe
ZlBqvLo7iY4F9fwwkIy4VnJcZgo3kLU8zFIMsRUVyAvjQLaGH/0Nd4hYTYYbxfxk
Qtn9cSZiY5+NczgJPNPn64gPx5QOEd+zVa/2J862VErLCEgP0dc1PklXlfj3vV3I
uVc3gPMjlsZanOW1CbnSZmvtNmxsDx93U28y5NzAZTWwZ1simDRpvWhLf5Sv3t/L
bLN8JEMAlOD5JlrNOVO6R6j+Ho34WxdUBMusXCBDeWtlBBIXkvXpv8xLucbcambS
o0JtB6VcQ1gyWeegUx24OKzB8XXCLWKCESSSMyQ/L5DmMRIpNXpObgCEuxpQTKhg
YbbgByfVxkvZgStpwCxWtH9inQ4Lxm7u3Q+AbIXT+7xxEhJLJJ4VtJQe7ppa3IMC
CJkz84i6OBvSWzrogPZBvbeAVZxN9qDrz6Bw48lkrqh3L0s5F43JhAC/X8Fl0EWn
eM1PGY2lxJChL2tyPMkOz8sBP3z2kJe61r66KZx//arFYfTu+HBSqe/yvm39XRv+
WBwGfeXoqRv6imFMHBh/OnTYUiWJPa8mHHWw5N7NyySGE7HQdxa0x0iznyEzd15G
TKWUNQiyvV/gbFPHvq5jxwX05RjliVAmz4250ex5IP2b1lEMT5Vvj2HDX2w524qd
V9P7PuplkOdsxtTDrJLY65eRhJBAwX4jIZyvG4hnrKm8Qsn4iJ+OVzaEdI5FnIu8
26VoJkYRPcDVc3yTIipob9zwUu5ciJ/0nS4TfIKpcbyZafwo6bsq9jbh1V2+faSR
zkn/i0bY67bV7vtZl/WyPJrhARYSvZRv/aAzYfG7mnfjmL2M9M0EO8V4GpA45yuw
ppZ63xNr5aCE5A0OOwr5WdcMbU/9ogooMfkPool0zYnF4hCEG6M3X/D+cJanQHn6
E74+2Zd43tXdGO8TzInDDVQ80LgpEtysxlBJaSqAaAj7c8hYclkgcD4TzwfwxvhN
WgB5MSPDg9+J/sr0ivHl2YmtKPMOp49FMAyw5F9yLBUxeMF61g62IMqXa5rfpuN2
N+JqAZDD/eLzMT7YKU+xvPvI9IMDwx5HuBoxGbybtMG5jeCBvZ8XqOa8LXnwd4Z2
+8bCKvATWGZx/IG2IJNgoLadshRNBuoWYXwBIz1PAL2yXOilBPPsqqYTL/3y1czE
+Yfjw6Kz0coL+TAHzAAZlXrfXsIlLL6kzIAYyNytZ8XJjCwTVVHNOlAQtoS8yZzH
+LNkEf02QakGVGtELAB+jmNOgtRsIHlozWcpk9fvPzR7wT5eG3HsRc9yZOLSS4OC
KAbDX5qtIynjvGvPb5K/Dcd01cP/WJhoxikDvqF+jO2q0jWymz+Nh72dV3bYHQZy
5eleaNtz683sTo707Cwz9xqchaHvUgxWVSBLWZDHYJDn+6H2uVndF+t6KBz/jY4+
w/ZP1OHuI32cSZueyDpzibK6ABBIDOVUNDdWfULCytN3kqVV1e9gRwAReNgDCjK7
6T82D2X1WlQaMV64fMxWnNYsYgohzx+IICJ4k+Kvxf+5bybA07IN3aEQAyCJyfwx
qwVYti61qjssXgV5+mWFWINhprppQhjGDQe/E/Vcyd5PV1fdowux0KeLYghr98BB
lvlfaAW1J3e5E0BaN18g2GgVJaVjX0p5AX0oVBE+Kxn4I0uhzcpnN6dbUOTz9C6E
loyAquxCKXOf8lpc8WKgA8YFSNtFN12n9iSHKwu3/h8QKU7S6jbTEQe9SwEVsPvT
fI3kPTnmF1tpGeDgspVFm6bxi6CEYWNjuSwLS1OVBLCmdR9VPmKMLT156zearyKx
VdRM1jvco15xQH8BX3O1Ay4/BKAhoIaGnruEu8eJOegH1QsLGQWS0P11P/m9ydaU
GzprlfrYwelL2bQTcAm6T75j5OOyqScq6/at5EDmLlnEShMaSfP8wI9IwqePD5hB
0Sbiq82DLK4p3xYmdmA2A4ZlOP+Zk9rDs9i2o/h6fBCluhVf85EViJ5967ZhjPHj
Uu9dtosg38WFsOzgoHYm7x58K+NFFRc0tr++6waA5fe78CsswvQFFpRc7mxtC4Bw
/sXSxdn/KSEHizKccQbeBPi36Lx3NuvvkbgktnOZtF4gYq38Q/1E5Aabh6LTIDFz
XxDagLjsjO88qBuetn6u2lFTN58VDpGX5yoMn6jIjbUKGYwHZNpudG12s1NKhptK
jW6wTXpJgs1xBgX+A47DvzwA3+LJBDqI5qTCoIWFyezoG89AV/6wUdOnx544uufu
0HMODejDo6i+wY9YIV2W+BOKbLrx2P4PVSRegoSmDCjG3o/DmzZmBP0Rpo1yv1Gg
FluYLrqV7V9N0YbNgmRSrSkUCIc6KgTu2Uq0IW9avtoN0XlQpoEqnnRqgcbfqtkl
YUliI44JhRvCzFq8pf2DZd+DtvhjY8g3/lEMN7tXGTBBipA2lCM8n4jxB+t0a55G
fCpTbrcB4JObgvKA3MS+K8qDUMAYClS/kmt71x1wt5gQM37OsntLBqInmDjlqPLi
PwHuVP8jB32MxilIWtUB8FrqAfuCqPoaFCqpk0WWx7i7UYQ77cS42x5QBhoCS22C
JVm2zLcqKhHUmLAHujUIbIRRm6+qQY+jXn6MfRyLYCxgCclINepuVWsFMH2aUOCu
jihH+NaInUfk724WmQ1AmdljLfiXQ82BNDPTFP9Ieksgm9bnwQmnWzpZMSLjHlui
IWfPsVnoN4zWpnBlYcfYFxrBsMvJ/wJH74c6JKrkZ0n38KyQ57sYt5xcMwSBrLAL
v707RPrC39qsARffiCr6X+WVaWWIiUvgjE131o7njitECMKcEgXPE0eoWGXpQLZb
PzM4av8eVYRdVGO29XrAoOez9Q8IC3N+f2VP11gAriFPSbxEhGJP9vXDXoDiMrIX
eXmM/pw5+reSdT0W0+w+gNPtu1fXpK/ELGfpIkERBeXJL9CVPiFl3Brd2uunZ6rN
85A+5+YOoK8+eEnPx8PzsjN2LcqizCsHLN29KIqRT1VczhbJvHsNyuhdNu0Iz4Ua
nLsKjUtKcvUku82pm34p6ZcgRImxlrSw8QPsiktEdt3YeX+TEVLxA98dbp7mwxpg
vAPbuhIqTgspQzD3Va5A9nOczPmkZQAvj+6fG55TY41QKzBrxj4+OsyQR5tE8MnV
0xz7Ath/9PBytapT25i8unv1nHVMnJudVGJjXkGYzIZOtrjJLL3xic5U7oocIxrh
QJ3Uout3jI8X/90BvHtSOnd9r7NGspShXEXH0FmN215pJbuqv/L6nMGigrJaBgXb
oV7E6rlsXJZ4xNod/nAwVKgY/HP7lPZsvIYg9kKbvHY+Tf8PG5Oy8Ejt9t+pQebt
zYKXBN8a/NAFnxlvzQl7C1uJ81IzjRP1rMFGi1DTVGb8/B/IYzOB+Rj84Wtfhz4W
cuj7iDSXdMEgA4l9FLT2H+wyYkk9YT+E6MTj7h1Yzbe7kM5JD3/3bKMWPE88Z5kj
XM7Q42HjI6B4NouDwpglvO9bwZY2+wsi5GV23JY9fY5E2woQbEuIz4XhIEuDzHRt
OSopWNHf1OkGolQ4MpGBuonbb3Xeptd8bFVFzL9F8Is+dnIhPSHDFyP3e0hzfbPn
S58vE1G5xsHkynxXDhzg/luU+nIt6bFLb2mxqUCxGOplG3WBHrUMOVIYCAYBQDq3
Ue7Jcgnnp6ZjurHbLX1Gc6g8M83ui4kNjw8Htt4yWnm0akqV0hvScDdy3Xmede+z
s9aZQW8pD4C/41SMGWRcG1MbNXcLdUwS5BY1u8Az5OOugso7Rh6gzW7+6H2X331O
OxKsI/+SJX3ijJNWjz/qkMlTIn7QviG3fFbzo6c/rrIWb5HfNfWmpwxnzN9KV/xY
Q0hv7vdO3h0FANQTEoHYIOpXjv6nQ4LItyWpuoeoTFQPmV+j5F2DhZSvXMBpTM+R
qa5FtdwSDEYImLbFHc6Q9tKKXTkytBYwLBoc+BM4FYidnHByPHwXICid9Ox6uLKZ
vpq84VKu+DtiUi4CBMXSsGDyo1CreQJY0+a/lYn8TzQySbPgiAM3RiHMdvDGlqat
ud2mRwJmIMemSKHUIPyMFsaueN+FafxYSDLT1Q3TmpqOmG+TlIM/MFQxl86A6Yv0
KuCh1Y5DxOLlgvYN+d6J7uipqIapOnKpBemopOOyvyZpY1x8/kKBLYWfFmK/fukK
Bg1Y408gbQU/szFfDWcX+m6yBl2gk5aoWTy7gYICJPb3TlLydpQsftFk6FdcL61T
Kzhlt5TeS5D1Ed0m49nhJt7OzK1zcKgVUKVZTnN8fbEI0vdSoPE/9BWzFYJ41+1c
mAI/bwvgDWoiAp7TfG3uJYQmkvJQ8EfRm8k+YRX1q4BUZNAVen7lVcl8zPOZp35U
k8wvm6N71n8u5YgrwDvthqg0/Lly1xn8DK47MnhcJESHOwzc8QHbSY8LCbzCe+kO
VgCgATLpabBVGX7qwH+JxdUN/y2bcpzjmr/jY4I1Albf67jmwO8Lw5gxhLJftNcO
MocRLbRO+D+HV/zVX4AXkf8keOJKqVVYSY1KR9CcuOqNgAA6KqP6BdNDnGhw4v8l
/l2DuX3toiIYNFQRPTXabRU3aVWfQGRSt/2ixN+Q5UFUdaljmRXYzwjc6p5wyA+R
T3OS+CXIkhECFSnlmY8QqtJZIfNWcqx8am44ADscWaeX6j08BOW9vOWTKABrahFj
pMU1qeyomoZnkyipitfZIJT6L4w1jLco0Ss3IJn2KZnasqEIs4kNnJ8R3NZpNxMP
0LoudgOsG7N+Aao/HGdCGgI+CQ0JpBRYgXpbyjJUaTBbJeJiGPaJTpjYJpKQFFUP
NrMJP3pZozun5nRIXxYi3qZb9ArNWF2y4OvhjuJR4KwNtYnXEBRKDrX9F522ELUg
ubjtbnf3mHDrCkV8YhQqHQA8TI1I2kagUW8WcSRKMTY+AlIm+9ojKMGTaHmo4x8+
AHomny/elX9PV+zbkM0c75lSO6GFIcC2NsI+Drugj6ZgswpehkK38Gpjpl5iPjcF
EAo8sV1b9DIDkmmyF4M0tFKiIohxEXGAkD9EAGvj+x6Kffm5/qH6f0n8DuclxPex
/XleMZiyrRTDRP5Vjz/VoOx4d4jn2qQOqG8bvKz2HBLMzgQrMCGlNryHVncxNrwu
GzGYAThPq1E0JIpRLaX7+iPIbF8M5p03L+AoCi+mqJce/f62r/AsOnYedE0UWvgz
V/eqR1jIMqVhEUmV4mqG8KyuT2oH5fZ6TSFWU/v4oUsg3ThwWBwlMekcJwAETI3K
5Chs72yrCDCne4q3gUv2oKfcdPhS1UGRx+VL58PlqwllCYTQzmefhsYGJdO0x1bI
0kFCgT89xh05DBMYf3fQrjTWptiEYh///EGI1/Zide5rMxtzJOCYWYhs3C1S/OMA
R86NVKrKoZc0KRcXUkPXJv0KpuPv/HorL3QB+VYURIOC46KnaHWDIntc4ff4sbBn
TMar+BJpoSJApl5a1kIT2hWVXIxdrxKbhxZYULNquTNGwocX0z9NWiRp5Y+h4qIC
T5n/TprLhxDGcov4Jnv+3Dq+yBF9aufgRCuTyFCOd1KO6qJQBBXruRZpt28PPqlf
G+3OnyzkV/Sf19qiK01MRIkZl00zVat3yjZ2mO7e/sd3H6KE87PRMEQdxXchh7SP
zif3EFVv6z63S3MvS7Rz9hEfDPpjnB1XgyUkd0DUMLtUt9pFI+ToFbeKW5GpUCi0
XnILakA+N6g8ODMLR9dDKLMvwdTRNUCM3QpztveAXG5WOPkZN/sJkeHpdZumqosD
yA+ChL0C/7Z3Rn5L9tf3jNAtyB0ZPisRxmNN6OYJTurmpJ8fEwNyFQJ6hZ4DKa1Y
3E0YhNTLmGXePngaYXPJIglNL8ArZrAP/nZuVoY6wgKO1jKxMkXeQK5LVbiYtOiT
xg0nPZuR+nKQ0XuItFIdu3EDuqqD+DRHjBkPVd1KYLyKk/Qg4z/ms25jMH+kVqDe
TjdF/g504XHlepsd3sLQB8vtij7tj1Iy/ugLlLK/7CjuQvZwt3pwA5qxeX3rxP4v
mJZRyF2g/PmjB8rAB47XJRiANDC0qDUQKioEH3q+1Z9i7Z8Nw84c9R6Kg4s+PhOO
vs1b7c03G8j+cTcf7JpLGNiyCdre8bRDoEV/ASYH8yHB07iDrErBD3umiExVj93B
RQkwrLi6IpQnkYtBEOJpardGhIZrO8ImvQFsWwyc3E+nxT6bBS5ow+4rGQRMctP5
4+GFxYwNQc02Uyw884BrioudKQuu8et5WKhNQIgN7wkSeOqdz7VLOWW/zg2CW96/
NAcTjxx9bnLMPEMPiP8oSatN2gkzE2ETes/RAL+OAeNqGxYYJFkxAIUW7zEQ7Ux/
vMLrqAoNiH449PpuQ9kczEbMFcWsNGj5EfcBXNj/XcP3Hv8OE528FrrF+SjusheK
uXQV2ARNeWaFqUPEwrSc4Q2bTdNbYmEDUkZ3Ej/SWReyeyrk2DHtxU53HSqNiQUs
JH+c5ElI8F1dmGcE3kG1nTDQJ8WLUtoC70qTbam0PL5FRGo0uNgAs/WdFaxsFyYk
3PqPlcktFq+3aAM07BQ7A/WLj648UOcLayZqc0FZc17zkEZ+/yE5p3Bp0s0SHH7P
JngkjKGa88sLRTPOVtJpA/oyMXmTNeEBGFrQPoZz5tR2qpPU2ieTfQzHCkMZmgZS
mVhsSWnL30omT3hTPsGWuNe7FVdYFd75MLUaPtBl2G3T+2ccb+r0178wJKNMURZZ
O4vR5qs8IlRS3222aHc9r0U1GFKkgmZ6nVasD72qul6+PfFDbIcd7MjBAoeLN8oK
Ot5JcR00sXxPpRxsOeOewKe08hAZr0IF1IPQWbQDJGOkf5NKxCZgOZQvat8DjUeA
lY8hFN1eLWtJxt3SFP8HNRJxh3yNW4CwhA0h6BnXyJpMrbO2+t5fdZVYOJOJBn/m
yJHXAQGMVy60uxf5QP/D3f43SZORfVLly0K5rLEoV9j7QFDhcFWcI4LBIFvm7UfG
64HkAtt/OP+PLwZ8ImHi/QFi83QZUIH3dlkefN4rEIQyOk8Zvm2BFD+o8U2fvyBI
CpnemWz8HEw8UBdWMeSvCljmbr264XBeyyT2iQUxBSr6RRYtg08q5pxLS0vWASMZ
v4SbVeNsXgtu3+dsq5uubVZz46R5G81kEJ1nTcbJRwi7V+3meaAbbTT3jXwxeMD3
JT6YUg3rgnMgwHpmOtPdJLtgRTPKnvID4ZSiHO5gMIojA7r/pcmPMKyDyOoRVDKj
PDFaW1HCtSaN/SpEOAA3FXraA6oGdS/CiKjFZlLjrq3e6Q+pRyDMCYBWpvunYCjV
5cN+o1z6c+RIwYpmCctEPfLFvSg7hjmFlquz8resodIL3lFeF5k/Tj1jfMYav7qN
+HPL/NuFsg3eHOl4+I6O/PQBWoyhGy1q14yUcsrMNeOussZ46YjzLJnAGufBOe0D
3jiw+g+eD0PE9vRxDZyHeoI5BppU0sYKbb4HB3f5REBnxWcZ6mT0oRc6A3QnlBQQ
4VDTzhjGzlG5XYsZGVLM3ytpSM97p6pz0tZJLHpnnb4IESFDlpy2csKCVohCkgdM
P2ms31IuHW/qsqtA5B6E/U/PMkkDdYRkYuhuUe0r9IxPwy3Y2RVGj3UCpaF/j3iF
93NDUz4eIKn6OcIzbn4XG+Se+2wn/VZoD9thGzcFfvj0oSBPmaRcHNjkW6wXR53r
KVJ69AYelCzxfx6XO4xlQ3bO3dZr02uMPUz6sc+OY7xrLzw2W3bNOX6CtRgkvdGy
O3iv5KYDCpL7JIim6JkJRerQXM/y2uPhDOdATehXlLit3wmF9YdUbK6rt78JqV4s
ESm5e9fDnKMze/FLcwzGPMF/numBGnY3Bidkt8Qn2bQB2TW10Mrwk50vm16E6wg5
SHqH2sAlhVFi8hq43CIjf/6KNTlTOwmc8BawejPrDgRsey/f5b0MxTxR8VPsFClk
V9QeqRC9uQVHG303eKcShfkA64/yagFGfnBgEx/H8Swu787/74kWq8x5wKaeW5Yh
doDX3Sl6XlF3aVj0xcsVOl/GZ3hb0BMPlDgLumoTmx3a5Rr9KAGkZPDWrAXc6R5m
IdpZ/A04zDjVjqa7N8+WHPrNssFFeqiHljtNpqe3eoJY22Fy8sPv+C9zAjprjnDy
oafV7uLSEpKrcHxHLiyejvrhhXWG0aQJGz0jhZf4Asdaf0K0Z83/PTSSCSO8V/m8
ZPlqYgmn9Ldp4DCAiHpwf44ts2k2R+2Y12/RAHLi501ABQ5xwsAO7EATpIx9YIah
J2K0sP647GE1AidUGPQyphN3slrcuEeUegRpgx8WrZbyrNtJF7TpyMWqW1sjEiIv
aAIJWlUlxazYYSmzfsf+bvacYtSttRxUJYlojEY6G560x9WJRZnUo0TiBImziCcs
6f1sk9CMQX4F0Ifiqz0/MZGXKrKYNNavpHRKZVNpT28Ct33LB1FOxRQKFF9UteNH
DCfU3en1Ah7g9xawp9G6f33cnZ/JdV4aJ7pmqJNRYEranc+qazjnLQmNY6wQGlK4
RBdlnRgKCtqpFyepz+GawwPaCvpvtWkiSv2meHhSvKW2YVb6GpRUjvPJ2w1oBcQg
7XVUF/bgLtZxizf1JROrvaM9mCA9rM+C1KgQTXobR+rV9WhLKGVDUx7TCsJfcxJG
RPd+OEr4noumx7jcI11F+h8IQnyjhIUcJBhh1dItYK2tgCFF9iYlhETWcMWrantr
JKumSqOdPzHnougnh1UjEKOaFOIc/J8SypkiT9rbt4ALavm7XNnDtuGesmmPzPza
7EZo4Az7G1RwEqIIOB650J2KfuVPM+EXU8c12Vkg6up5p9kBTgF+JM2VWdXG2/dK
LD2zuloGjjwxW87PSob+ey9NiKEjsMXiNRsq9nm/l7IWsrRtLyjs0suywN6x/GHr
Qy9x7cqLNQQXWqtuocBN7F543gxV7ylXmdwZbikU+R9KFFv7mZuGgYp3u16BmGwB
RGF8RMnxznBtJGmKobFDfyXydepYdUGIQlXrp/tjAJSZJ0y9ZTN0b8jh/IQHe6N8
SFdSQQpCs1TfJHZUIaVcnPN/fv8HDQ9O77wkjxszWbf2K9ajnBS+/RVoeDVk8STo
17V7FGJcB1eRRV2DpzJIYBAs0bzcjnQnj3ZD96GFGMREfoPS6KftXmYj/znBiQG8
ih1z02q3nHM0MNjy0LhflbFOOz07MhDGvJaFu1aOwaTzTGp7GMXTUoTwnSCgJHNO
atV5TRj+X8uE5SeBGD5+DGUNJ8Cd/8gOxg1bse4K/fNdYLQiDhJ3cL2+YR2p6PyQ
L/QcUFLngWRpOizxTQu7tUebIbRFtFHXB1SVybg8AmTFNix7DKRQIOTf4NptN4oS
ydKarilpsMriPDtYFiEOSzWUtpYNOSCDdkFFA0i3ON2zChkaVxWpb61Q5b+lUphN
ijsq0L9nVWf5fmz/tAuQGCSeVKTU0bqfPdth2eI9Lrc5D4Qt+w7G98sqQ8Zc4o8A
naQbKVNz3s3fm2Xlb1KMD0nXX1FCVcvKsLHKeUsZuStycRKiwE3k9WnOIe4n/HNy
sO7dtudjHGqhGrgJKXd6OZ0IXsULtFd2ZDqnHY/H36xompX3lf14j3EhvJ27kkLF
/CfA/RhaTxL01U9/9LSegDuyep7XCIKgYsnjlNLDZX+0IwavrPvDdugIBKh3v19G
yS9voXnRtkK0QzbGGubaYweT4/K6+YydVtob4pqK/4BpFWs9l9S4ndVKFLUew//i
XB4zz4SW2ylfq69P5u3QTpRKsinfXdfd5zl4WKRMQcS8KvWqHlO95WkMbRboKNcw
tsRSyqVGEUqO3/AGSsMrSpPqSCTF2qhZdRQOKyAnu/cpoxhlXhbNzo4gnl3rhb5W
qqSVElG8z6Y/ACX4hWq93wY9SaUjT3hCu4jkJuDv9Werbu5ZRAWvAxMbrMoqKFdV
wpin3jYGmL52xCwxab/309OHOfPA5ptZv9KJyx98FIj+bF5xFzjMARtJgsWQtf9s
hnc2sB4vrlScoZHE/OmJcLtBnvUL4BQRtt9XbNAJnWEg9gFJdBK8FL47swVUyF4O
7lfQ2+lruZac/x4LXV39JssWe5j78hJHbfpF82OF7lwH8YV+/REcJ1dHsblTE2C+
Q03aJHKj42i8hhVjzS7dg9iOk83E69M8qQpjZ9aTxoI2npJt8gy+rAGV+gRSbN5F
axCewnEYQe0xOPKMnIaGE2aOwzl2f6fKxHcvN0H4VfJRUp1R3QL+PgZ2Ni/KG/pv
jeOKbvacP18R59GMbjNz8IcP+quNdzcEQ55blGuEsPoIPQ//iRMb9sleEkhslHsq
zykIe73BSE59L0L0EBRaW6lfjqdsz/TAgp8n3H0jP7eMh3jbZ2XlRtH/gNASDkEJ
92w4PDZnhMLIMb5+1dNkF6cNMyBm/g/YDbaJl7BMy3nuPIJfakSigAw3trbkusVh
fcDKw6TOFBAIgahIiYkHphjLTbNTQg8LbvjI6ibgfWN7F7+MYGT4J9KDb1uRxvPQ
+cpzmPY4vELjgkFSli08wt8Sr9QzQGw57vdSqUHSMZK9D1mVB/2tECBC7/nz+xXF
6UlCnUiTEvMcmJCw2Gzv9MoAg/u4Nb49HcJCepO+scpvvlnS1Afif1IJC62fLBqV
qEK862Zj1jOkoVTnIPFqHS3WjV27r35uE/CsPx/ae94E0UguHfSbeS54+wwPlvIV
TegNvWLjm7yIv/TthFDOw4g4WPRiDvgUmHSlUwzi8cbgt5SBy3xWeyDDaP5EWwzU
rO1UMuhHJlBXaC9xn814JHxebRspgCVwdz+T5B/nI50GO3iZWgaBoorKbGy2VWdJ
Es5oBx29uUSOwBDRMlK0aXWLusFFJCjI31C8Abh8rmThC5/YtWHYh5RF8uxtldsR
UbbJ5Q3rmic76eBx51S2NOl0OulEIF5U8y8lQMYpTprw7wZ3LY826qoxJUgRJt+t
/WZHIeXk9OM0vuknn6bReSPahjDONFo6R1I8PJ4mxhdwrYgF2Xe8a/uMmLGAPGkb
dVpZc/EgKX84ECP3Lf+6j9a4IyydXFBiVafXqk5j34043eVzGGDQWpf5fwNpZcYx
ESjqvQzwN26URwGsq7vl6yg9lM8gn35NZLJ6pB2ZrwxgSyhAl1Pp6/Jd3xDQHMx1
F8kz/ise7Sx4vlyh0iFpVcvLmrIBEy9K+QsBHgz1aFYnxdBnzWK1SSgahri3Qkx5
9v7G6v19kjbXQuMTl72/5D44WZLoGYZPR0k4o2AEpsSOBanmboruaKXrKCR3a6Nw
dbbCv8ExZ/bH16cTMtprH8ZJR8rZ6ijcjoJY57lHJI75XqSulb6Q3SZqMoUGRToG
STWY6w8qmOSQDd8iQ/qskIwfoujefGhaNnmDwozJDI5go3oxiiUqHtmzOjyfVXxI
Rr7Bh+4dSLEg4xuCaWi89IO2t2P1VXPHQuZCvjPscmML+3SOae7KJParYagrlRWC
xTwx0JrufFaybtgjvgPZQ+2aIoxjBLWn0UBgYo37QsQ3RQZRs89yuBTXx2hPQaVa
glFzFJS1kTRhZbtJmITYUEFvkgt/oHuM+szQSpHbSAuZaKNEvngss4vjYnoXXsal
kUJWVq1pZSbwPMXVwy6HxEtvUrKOZ7up9uZ8CcU0pCxV0A+DpIkKfRLFmPxFgRq1
rhy4kMYhyc0upnMURuf+l+RBg3KGTf7ghmZmp8nrYesSaLf/8+4xRtCtBNVtaG+a
zJk/1GQG0JWVMCu1yIUVCMA1APD8nTlUarre3R+zVQ2DQn1FzCKcnurFzEP+U95x
y1dnh/N6vlY8E0sQ1sDNPWqmDxxYz29OjS2qp/k7eXDBioUCN12o5mpCFsI0h7nr
TIHkyM8jK+UEN598SACG3eaQ8W2B4T+d8+WjrFphF9VqxitMxOeMkaU+N8KZCvdj
gs8YeRwe/sEXycJgZzXiGCewIfkeEUTaSw08THt5HR6FQXfuY4rqOs646YqRZ7cW
XJeJJG768I1I2DZYM7dBsmZzkea+aNfKJVi+uALN+KCIL2UwdeV9flOheV1XZzpL
xM1CYJ2Fh8KqJ2/zvyjCh7xLsGZ8guoohjF3YSxJeZtfUNpccDo+8oaqmm+XMqiB
/Ez9fuwnP5mI7JvTS2lajkW0xbslDUkMZmsNvvjy1S1o4bPauGyHh3xa6oy7UCD9
I45R+YdEc0FZcCvo4lOlGjhgzggfjT8SZLCtmDmfBox65uSwIxcqsZrV++7O/jzP
wNi/FvVRwZhcF2Zh/HF9f+EDPiJNA7U5M4Y9loBJrhLh0PkX5RRfLIJhcEyuO69U
mfYgNHzOxARTldv7Ziz+nUds4RnxVw0fk7SQdiCyDX5fIyiKtAcXR3aCuAXkqkn+
soQcsZdSz3QjajV1557+cTznGeTOUx1uK5ptq8pkySrwZVbwT+FhMEKLHmuC6vmg
2/SbxWcHxVy6Q2X5u51v/R2f3ZMgtoZYzyB0Yam6I5vGomNpyBAZLGWN3xvn6Rpq
rWFxtXa4KYsxjdmy5gs5Ji+9Z2ytu8dTiuCymsLHCyL0nImb403KAk/XWWk4Spez
2dSf0R2O7smS6Hb8mFueUWOnlGnQAb13TCUNxfDVDGiuCvxYXfVHKWHqLGxpcJaR
QIQxeCyszEmqLlSWcUXjjtKVufAmWjepn/amGy8ErKWFqi7TqVXK/0Oetjd0Ao/7
0vml1/OUaA6hB/Zt/SSbBIg40OaIg1Vq/7IzlSgqYGCHi4h/Scsx4VAdOknlg/+3
V7SydIfViwJ24d0eOClhWSgvcRAPNAJ/pQchRtG8clUB/IRaxnsH6Daunvlro7It
LQPZ/x2QMhVWLTMjnoywqiIovC4xOeTz4LCLwvgXrsfrtoeP6xrbQO3YonliiRI4
KXiZe7I1sbsNzqHwPO67WrUSg63Y3JKA76ir1x83Do0Wj3wYYiUDRNZ0b0nKHKBX
MI9uWJe02YVtDJjjSBMvZCtwP+tAT6eRIw80iQKpi4FqZOek7UT9vMO9/V6yyNZu
ryVsE27FpYgiLJb17LzMkpl0HItFLb0JIn/51G1TandoGzBz8W3kmjbRS8HHE9+c
pBNgsfjZg2bKY531wQklJPncQWdu+ls67OoXxjtYW1js7P2DU1R/OKJxk2BeaVWP
f6tQVABbNpcDpdEuerBgZ61fjrxAXRJqvDtCCC34F8ivXdiq7mEnazBM6WcaCHLm
xelp7I5IFWmb8cixFrHBMenxyNo7vF+WmUwDbOQl86GUdEvQWVaDe0Vj02pvaWq/
+JWuB8b7CQfBYBvjmvGmsAyapySBjKPbL800VCpTspA8GNcDN8/I4byOuiHXkEUi
eg2TdjCo6VwP35RRdgQexSIT7BXpcE9OWUS7Wn/vmFCgx1Mf0i+E4glIST5oFooA
GZecEGTnEQwEZ3EtMff5i/cqckrgSGtCRCx/iOiZj7CwO2m+VUYUrmsefzKTSaXb
NGqEnKyrRKfglc+pMT2bisWI4ppV7DgYTm+OCdneUzGW3JFs3i+p3i+pfxWt9xez
H12NDbpcw1MH0J7AHaqyCH8xD0dlewbFJpcfJTNnG+kGibJwV/X2/RlB61T9UbgZ
FPlJbljdD9hX+H9luCx32wNem3Cp/HiFpRAzmVNaawsnSDUpL5gCDhrEf7halCvk
kaTpUZwzReIw7299+/ij0AH1+Xcxjp9SS63SuzKcBhn9hTTjx8bTUa0U9VSOLyJz
Rl/04INp31m9+C8Jt9HU2Iyv9LuCaQ/yK74pa9RNATfWUhburikveTHA1KrjWU6I
YHTqbBuB57XJSleBqG3z0C3/CcwZaco5QTQR3QijXMktCwKzLgYepLRpCYrbZbtB
VsYB1aJ8/pITpwiytfqbzOIHwJKZzGj7sKWnUVXT09AHrsJiFFWPFNF3KaI6p7tn
E5+/gM8tYbq479GqRLK2bKK6VH6sG8GVAGNsp4hm12+7gJTX857QCoaPAjVTiUfN
aBtthOg/MZ2ZbCN+228JfSjcUhk2ewtRz9GSshcy/h2KlNKkrZuOXvEUmegsvpgt
GwInpGhkkGUOllCxQBZqylGKvRowN8X40FQMVD13LlW7QRGCJq7lKHPbVEh0+gKJ
W5Rud3Mbitd1xQH9UkJn1VVP5RPrA5m2qxTaaoQ1tL13TIJZNkUzlkcrWJL59kD0
Fm7k+ltQdgjD4aUHYaPFuqNzITFGk9mT7nNyj6GXGDnLnfKMsh9OYiVC1ovL5cDt
VpLvasvzHROKg+/iWSjOmTUdlhZn9UuC/zraagYhHA58Q8IQFUsuE1grc/47PG+M
JRX2kTgh6Te8uPbNNxE/LjryB75lsYk/QaWzgnJ4Dmyq24c904fLoLOryNnWV+tp
U4Cvo47us8z7i9MHX6fKUXGMt5GKyApxdyzqlD0atFJ3I3ocuwCZGbxrAa2RkTKR
jxNpNA6ymNIcBWEbHPnd8y28mJHz7usthecmeegfRYhya3rn0Xdbw+ghkqTHJ7T5
tGAyYLD8WZc97njEcJb0RNmaZ8MNfWCHU/EiqWHSyNYV7nwBC31nEfgEDIqi28ij
Qs2LGifp9PRc5YeI74Z7iEWzKFsB8XP2irMseYumdf0ni/nhduSdXZgZAAbZ5ZG1
6hw4nzJyhc/tms7OFknyKS4SLsgSQL9FiSnoAeHcN6AANEiyRR4wcgybuzphdks6
cUPS3jF1JqXteMg4lKBcLq8jHTAdXmsovD802N8CShuzRbxZSIWPHefPoWX1IE56
4ij1F9xkvWVED07QpWX+NdNfhHzENQkhg2TVrbIuCJZiHyb3Vm1vM3pXVGhG4i/e
JKRlmzDymcIXy468tRUKyPyYCuhN3n6ZjhpXmS1uep/ybXEMptIj4fDGyOfqlQO9
bI603iijhN2LB5VAzZ8qsETwkDPrNRDlhNuN47TnPxu1PLCJsgLDS/RoTAQzRByx
UxcfCnWhaxqtXIVeY1LpVAS2NgcDgJCiOh68ZC7KOxkGc+hBXdQAWIn/dpmNkKRw
lzX9tKrI9q172X0+Z5CYssmN48p7zpcICNn7sSfJUw/6wspdXXkVwstVj0bj2gMo
qWFqylx1GDzYxtCqDSqMmOZLs52KNK2x2PHhv7shnUB2qtLpR6IaUk7qge7SkTf4
v+C2zpIaR4bRPkj7C6ZA6PY4CDm69SxZvJw4eRF/0CmdxPl+f/N6HVLh0U6DXR9Z
d69GI83MsNZMiMwAl4mz6/qs7ZEhl0TcTsFolvPQXCoDI2Sv3eoLnc6CR21F/Alu
aCNesc5ELGyR3Fkp2E8fk3zKcEQ8YxTqOHkGqo5ZGOqcfmyKffYNzZTlqGLVbdAK
K5OLmOR3fKjNIHJvQca07ZlXLEYyCT7Lh6pCjwWpDLe/G1CUj/32SiE5rTPjZmc9
2Wuv79dVYMIvAKTJQoXHNurv1rw4oJNVbWQwoJCBzK6JgUsF+S1EXv+8KgPhv62/
k7ksyR/s0r+v2SzifjsjZP5dDlYf1bkM5++jM8N9XzOIcSLYuejDhFkIvhbBgjxO
TI5iznIgjbr2yJVKGqa1ek7fVUpbTCS+kWQjp3g0HgTYtiJOkjxfU+h7KZCMgJD3
Qj/UYwBC/qrTpB7wkCCOshr9AWgPG8kCYQTUo+SGdNjzZI+qVilWse2cTD6GCuIu
sBA7dDZ1ecPFlnbtZGcvYkYGXJno/QwZSqwOv0g6XnCCm14AsdK1QLQNY06UG8ax
Zp9kxzeVcY24y0rXsN22IGPhCnsTVgE7NMVRMIcPswMe0OGsa8Vp/U9kh8mnh1O7
nEefXmYHH+7Ui6zNXVCXOJHUAX2zQh7HZ67kZGQY9olGnAu3xQeivNsNrmCHlnww
ZMugL0c+So0oK5rdFK10F/iHepzfvNBmgGGCDdKYg602F3ZMwW2NvXoVMoBgV5wc
Ddmd/Ipe84DOWJopjD+uo2TxFdA+A6NrjT0go9uxvCcb5Cfg7gdZdUKBjGsjEqFK
uqPzglK/HzNxFyVmqb7fmuppKRkRqZGhDSoqOeQH7byH2XYsLkBaT8NhRzoh4+hG
c7gDHp9QrERDC0J0eSMaLCCxkvdaZMbk3RhS9vtB+V4zR2wcL0zwiFZiv0dZwokn
S+ZXQKnLk57lng7PUVm5khaZw7hcSt6kVKOinLA2WX2PgU7anNDEMt7Ks14gjnYg
Uf+ldR8kQDduwyDyWR4bqC2L94LmxhphY1GyTW2iwwQHyB5vF1nCXPcFHix3XQHP
mdmeL2F1cqEpN36KZra2/9RbTfPas7arqT/7K7QON+ElWpTlL/Fd3XTgG99G8JJv
lSVITdEmifcdeDDXOVQshrOSrO0cFTkrh0hu7KC9AxjqWvEIkK8Ma9877JF/dOCU
t8/xHViVDvJUBU2uTSbmF5/3+owk7BmF3uKlDx6oY8NDPP9QOfXDAfge3SP5h0Cf
UfTQOrJtraIsbJElnfazLP2Bim5apYT0BH3voVQR1sIwiKxxtEiVwF+xWL8fOtaI
vx4zO95l+sR8h7dVIgkUL93itvNqZ2oR/JwrJJjTwcRgvJ1blX9RcEqHWojqdXpw
/1xRR1Ku0Od9WXnE1M5WVBvqKDw4McxyXkpF55F77Nrb7NsquyczQNPk7fC7YuKc
CKv9LJK/bOpltKTnvC3ZHdAZIsbg1Orb3z/eMoGV523os3NRnarp9sXLN2t0a0VQ
A63Lk9ilI3lHM42kz76aJYXXLt2XjvgY0h9gTKnXyWp7P9s1HyyIZWhZKz2EMFPh
gYV2oEaz2/vqjhTP+DoWtSI2mawsZl0LOCSg+XUMpe3NKe6evF0ouaYot1VvF9Cj
RiEfkZ4BpbMP0rYYURm3cBg0+oAAPDQlwu777pyYMNauyZhkeia/9M1hX/jXBmh/
joyA/S/Ld5O133G4Njekl4IECRGfK8V7V9djVEnzynRGTyqMMcNTuK9BzVepFWk9
YicPwH8I+Y6Mgrtip8XhTE8CW0c3vo8namQgd2/8axQ7gb9kPcsrXBXHcF21UV3l
LJvaFEuHNm96oIcy1KpU6+PGaiWcurDnEwOiqWPhFIbZNQR0bWo/49bohvR909Ze
CXXVrvwUhFTVHF7q86+hEY/qClVCo49P3Yg+lZ0PVSUXec4fggFSaZ67bJBeuOub
t1h8/dcqEXLm6Qmh4SIwtgn7yzLmjLbE2rvivYmd/I5EUK7uEauBjO0fJgUBlgqB
fucf+9xxBNMHlHV+L8J1g0eaUVN8ceET6IEUT+CJ6afHRnMzJspRA210jis+cXAa
W0iYgz4ZSk1L/wfEXohocV2gp1L//Djjd8AkA8xYZUjn81buuqmp0/fS/ur4RIhO
JJlXahjx+hc3bxSSnY5O7R/CvRCvHmPWMYt4m9AYsiBksCopsWZkJwW2YMzcyRsM
bZs57IHlePIa+EU1eoKfla3+iTmTfkv0YUZPMhHU8Qy0vqSvA1e2w21fyttXis1J
9y7AhhVwz/dLiFc5krXW4m9/ygY6Hhi53unPLCjumtoerSZBt294C/3K1WRuY461
eLJZG2dW547joayJeiuhD9duZVw7+oFkBrJv+xxEgT5oNC5t5+9t3SAcPEA9rSGv
rKxm2+cIqhvJ2p8yh62xELQbpUF96keaUoZcaXSMIZ/jgcw8aBUqQs8bW4vPVqbl
KEJ7FLKk7v88Usm9kfa1UxadN/5LN7qUO9/Nj4WmWRdyCA1lKzKnaB6pX0sVBdaJ
CE0DhNXrgOVTDbCF2FkdYhylfGjq9yhJOKwjNry3rgSdFosdQ/uWhXpYwXfXjoGf
LwOLUcTUFC+seAUSI7pR2naDTMh+4oZQ9f0JzkM7jBJwhDXj5HVi+O6E0C9qPzHv
44JnIChxH8uVzoOFkf47N1Ap/yjl2ej96xfzZltEKhLZ+cI6ARRZ7Yw6g/cSMS7C
0GunTS66AfN1woAI3uhUhmw/MbEq1hLIhfl8l5vH1CYt18YShkBalBWCk09+JuN/
qPBHN2TeVV6B+wi5IDqMBFuMjzrqnx46oyMza8thbvbCVGotQXEGxpj+fpvkNDAr
CpciWZc9pckVRbQH4o/2glLg+jdON6/c2NFDlvLdBWycnYe2stwTuo1LcfKO/ZCe
sK8mE4FRI8hLKYKjpIhsYgFiBxAtEzmCDTwzDS2CgklZMx9vFXPOjux6U/hAPagU
Xro7aOA6V30cZ5ne705RYILUVeVaJc0n97iUJJAIFfKxlw4zsFx0pV2KackEjWlY
AofT3OpcuPjL1DXatNmNOlOeEX0f6uwUE9qSG0aHEZjUjBOG+kDaRm8gcG8DU62H
ekcGmv9EAp1OyIYRrUmcOzEliWZJoL4ScEyc8rogNDCz+1D5wgObEPnRTfLsJJ2y
eGNuW8danaTF6as5KSAf0+2Qb0iaja+cmFnGXxp1YRr/koF8Ow7e89J08Kmckt5H
ecau65XKjVrs+QTuqbzordwjL0OMS0CKfDPUn9L8SttCq3xOmAgmJ6NRFPqf7WI9
onrJsUD59JpNk/pnY6P/Dxz7ASXegcYIsQwV3qNBGmXst91/FTGuehiamZh0sTBD
8cbIvAM5K8XFgLjXLakPhr3PUwf7MJV+PlDNuUjNquHQ0h4JIvayaKL+CJlq7/q1
LuWFW5OTLjsghoPMHAy9J+11/aNRs8WV/zQaEWyGJDdsdLkSnlO7DvckRrwLU1Gk
NFjPSZwpU/yebKzKtlRTb5JyY2RSS88t7zRjW2vpe7pIfBKnlXQWmKA94eY2feOD
7fXVWNmXyAGbKrHbGE3zzsTy3j6p+QP93hEPCC7Z4XLYXeVRi8TdsjjerivpyZ2P
T/t1vHxO4QZfVABS0ogy0Inc9z105e+3dv/g5TO+IIdeXm0vKkjTeJSh1F9JQxJg
NsMeYT612wnOPUnQGB433SPw904lgb2uyE1JWjBZiX9GGh+gy2uNdCPigx1FPdFF
SuYwmvJLZViv6jGVjsk+DabunqBH0UO+zL6NCC2pSN4uJu4FSAXhq6/T+THYz1Dl
HrODQtCU+n6PLPX9qoQJxv50O7nQ3C+Lfnn5H7N36IhegavPw17IKgFHFrrnDRds
ieQiiTlzwSOXHmWdpeyZobrH8KBk+bVacQCJS7yehrnHI0Xw9ihvLF0DUI5Po6V3
+54pvnFQAB6MLBH3Fr4bu/lTntkBte2LDAldTpM7qpc8LstIxxF0A9UoS3tKevnD
Z3bIDcBPUUWobN6W4mun9UN3LxtV06Ql31cRjdx5tdYXDi4b0lDGEety7b89OHnL
JIRji7K+4iCmAaTJ9LxPdKFHBAUeATPTFVrEQoIbaFRCV6hfkD1bhFWaLeoPQUF5
lJcHDB7gF6wP0K463oSzCJXKFJXiyAJQMBGWS++KwQULSOWgTUBnzboadWru/XkZ
C40E4zZSU3zBn1ni4ONsTyCJ+xYo9Ad+zJoLw+xooGbwZO8Pj7Z6VMzWm6orkpSE
lwxqAWZfHZ6v1ID0evOn6/7c4zoR3Eg5iI5Cb+q9fF7bOZJyVtnD5PHQBH20mtC0
+OmwKVQrGnKw9DHUYEcSRIkqjipqXpjxs2CZOdTkzADaWf/5grdlMwHb67z5stj4
wPbjOUirlJ0ZBs3V6jUHX/5AHwUHhoUBPu1xYxyZE+UNdjZKem+whNJHrQvKfuqY
0twpNk3aaHe4e/qNCBaNwe+uwSCbX2Ii/Nm9FsjNZqTRR+wNEQG8fI+VyyfGtQu0
uBJAeJjAzgLOuDKBek3K0ijuwMp1ITyDXxrBTJSsCQm2gBQ4ql8PBCSmun/xVHTC
ZX2KmshEhB7/UWje8yezmnMsjLJEyYu/r+MCvbWAZdSUKG57+hrtWM9wXCrGwZiT
fAlsM+lJdFRE6UcqmcXkOVX7NByGhKoJzGVykzN04kZ6TKN0faW9qs3zsKVofxuU
rfhY8sbMjVMEyTk8ZwKPkxb8ET8rWDsGeLo6mJtzDIDMnWijomW+AvMZsGSYXoxx
EJABKsP12eO2RBTmiXYkKhijcKxsGA6WjYWIuMdD1KRWInK6rmAT2R/334JVJv5u
oFVvJzWuAklnlmSk/GOBat+TXhvHZ/9FevWupS5w7A5luAwt1pA4QqXjuOLGve12
F9SZcO8JqtVlj3HYMGmdrXhSzJugFt4VbTGcs75yw5fqBxzmNmx4Pxem1KIjVagF
ns5fPBz0PnlRwmsLWuEaaE+lMHQkae/ST9UPxRXT3k0uieFPg1OevfvuIt9INgF6
lg5UMuRTC8vcCiN5HQ0IVyO5mg0NrvJ6iTNLa3dQ8+1uVcK6VTcd+M07KZJAymiL
9TRXaC2NMTYkGVESR9gsIZJKQLJGtS3TPtQ8A5SOZLokzlEY9y2+WgVitBEh+5c7
1nSvzDFw8/7JdtuzOogs1Z7NX5tJdnPKAGZ0bBJyeMSgEunomCqgq89HUQewFyzM
2RIDakpYbryKVHeSeUEdKSbV92Jxx1kbSYbRZgDLXny8RFBU7YIWoNWbltqWjYXt
zSH6c/Jd73Zu6aOT9RMQExB40Q5AOeiAjy6yEni7FOlLGdZbbo6VwSFcD5KflpNQ
xjI/3CwykabokVdPoH0fmDNlGNRidOm1XB0S8/vt8AsPH2TyrbAHPrPQ61BnLDyP
leS/t3TtM056hltetQ2o6wq3j8T6UkQY/q3GFqJO9N+x418S8MReRPzvRphzuCQh
7iM0v0SCsAGBcPt/Fm3S1bt+3taasawmPHgnIQs++5bs+PHDZfBlRtU+RpSzPrm+
Rcpyt9vTt88XqIk8+bSgD929LymABjO8b4bw8kMDTAcCHek/eq0HS3faY5RHE7Id
3wETL0NFFlMg/OYRDrYZNw76oAx/p61KZudBDMbFaYSOwTSxwmHnAROR1nA/SFYK
xXBIkil2+UCoLdWfaAedPmtuHI7fT4yQGvRskO8mmT50y5j6T+PnjqKfNuvZ1EZu
hS8FW+VGESSdTgr9qYMyvm5hhfQt/BqI20/bf9A1/wQu74bh2Ye8CbWzkCquhwvc
myHyUw7sdK6YtiOTdyN/2ru0TV4VoMC0Iy/V8J4oRtF97rQfEmjZDUeQLXXAomfI
V/FtpalUTI7OaV9+IBFa/bNw7S0wPzI3fiybpmB0l+3n9LjL0vkPotHFNtxAPPOQ
9xG7++aB5fQV6Ptq/Tp1IY4Ku3Nx5Iakfnu7CI+huvzKE9qm9h9WYuuME0kxBMSr
FeH0Tj+oYwovvHJMAZ3hPRR5bl2+VS3wSGTfNvn2lNlNV+K2irXMrFYsIhrJD+5j
YeFq7mEr2osE8iRHycG4dikx9yG5eaWgemPjzMNsYIqEUS2mteKYShBobnITlBtF
+KhBuJRZSayOGbcNk5aWkTBMB5jpZEB+b4JDumzXTMvWbpxUV87TgHSZG4vcaDPx
pd0Dmp1Lx+g0vP5GH0nE7O1PAsDu+WKQKL7nVBUX1wNHaczEJ+uNFeomjqvVJ4vf
4Jpr/LU9iPR60hSySCCsq6NudnXYEfIaHBz7mWr3FDMmHHU2FJxVBr/6Y/hase8m
WPnqmz/UMu3Xm4AXcI18F+cCHE3pj2uz3CGqbTt2P+Cdgj9fpXhuq5DjhzIm9CMu
2cJVCJYw7Fhsm9odE08Vjf9LbM4nE8jbXyGpynDi2jghC+q3t31sdUNnbqvlqU1h
5MOnsEb/U9soKTu8ikX2jT5L/CsSlDbOu6i/CeMOQq9Rr8ZW0TYFq2e+F3fmuWRV
PGZpElIW6LjHyNhCO9LkYPe7gGoDiLdxVA6mq1WYBADCLv+uWrrvGaclEhF2fjlr
l17QWCGrIvbs+pTPjHEaKvn6fj3rwqaGVr2UBCrbBtLOy4PAONKthPRv/4UPJA2s
TXTmDFOinu/FpeSRAlOzR2Jk7la3X9nO2aE/sYQPyy6pFvgxkYw+ybWfoC/7hF34
JyBAogUJ++Igc9T4CUrPaYIkKeb/F/+KHifufUBzQJ0PV/3f4FNDA8Ext3G+VkZ7
YABZbwKRk4aidqF0IRDdBnaz62OIS1dHAAyysqS7BGuuREvOlcBOwz3fqOjiX+ZU
5O14RnNu+E+UmD+DCQdd05rbXg7IDXtLDVa1+S9retB1JwxqZFBH2OlFj9tpF38U
fxX6z6mso/PQpvoB30ep/wgdMa5jQ13jTPhJB67aW5Qr+O47Pv+hWWHTCw3FSarS
7mle16f5kfQMtPdPr3qTTSPfI49XfOtTzcb98+v51DtYjV/2D/BWifkmxZPGcd0D
ZSlfQq3y9Q4PZmj4yWJZtUMK0t/wKirxT0ZP1efTm7pR/AaR4h3CXtCQCLadirNt
O6Bn8RVAsEYRLZhGDLAG/1lMfgGFdR0K9MPUvqELaDzBPKuWfmXVPZB32nE29tqE
pH+IYyI/wGMXV59mnddjbi41uVDNTVfPI/7524nxlhmizPB2YzrYPQ4jQRQyoOye
bzAtTqHycsz6ob0BJ4F8WNGd47hyJUTV3+jYHJMAgDdNLGT0rkSElWFKa+cjgbOr
ZHOLrIUJHIs5AZZjv1r0rOhwfDQDyP0xaDzFfVYs0MUxraQnX3bbzPE74LQpw/0a
enE2DNOpYVHq7wzPx2hLtIVLMar1rEysRVCQ3FSUyNhifM9VLEc5uGV35B5BwXJ/
vNK/F4BIITk7r0UTzapI29rWvdSAQwI9Nef6lLelwq2f8yDb4fkLSpBHUlTsyw6I
SiFjXKUVNdxOVp6C1kiE1to4o6BgMtqVOXvklmBBDnvN7FSxHBhcNec1wx62KUI5
N/CWMz6Ok7dT7Reko9lcqAqgoO6yEDQSeXD91BetjpEhog5MrW1rswGg8RyVn8Ri
fqVwaAJ4RoIoK+cFD7X8LCbNV8F9mOhsQmHkJA9ysWfgtQ1Vxxz0lZuKBZaZZWyO
uGz2VcfW1kHdoANYei4KRSehqKJrEPdEJe6qTJeaFx5qSa7GmWrYzQDyhQyJWCbR
NP5oGUTaHEQL7330scvMlzHL8MQprv3oNAqKkSopHh9+9yGO74jtdDLkJVLT7fLs
0XGA6RLovWO+TQNTyKDk78PSzD8zxZFBWijhuEUjAIDWs+YtyDdtaoxZZH5DaOBt
HFXb8HD6YUcoR4xepEG/CCdEBG5S5IGEnQuwP/Cf67PKakgV4JH3GghGwewKqFup
7I471NBKfm+FHgqpdpXck/jnK5Kom1EjGTHQH5CJNpM/57sOD0kJo09AyXePRXVV
NfRX6hMTfRMgsI1rulfwg9dBPkDiRaN2kvL2gHyYbWFZtsTkcRvBGzKCUZbT5tPh
0jZzVdd4GTn+7Cl9v2QBI5HXVjUcJsxNtkt9Hg/Xdeo5gxGOAMu31xaT9w+2MMW1
qwP7GSZ1528YF/8bAnDkIn1NdpRi91e+oYtdf/0U89tWYebNcr4ZlOp8lmPdqX8D
jmvY7k2lcLAYO5tmHwAzcyu3H/fC37jvHJXne/071B5+Ps2EA2zs2b4fcG0bAh6+
MEj1ON9DDxFfe3Qxoj5OKKiExWfYUEVJogf/qWUd/n301H1kwzN265p2ZWcuoU5/
2i5PoZ9EbCYokQAUtQzDk1FxZDFO7kfVt5QegYm7fvMKaYKk7JzdtWuGp/+TyVQv
NKuDQuhvc1YiWtdr/YD1eESVlnLNVeA2CsAIF/ok4iN1dZXhytrU/lI0g/0pn2vN
PxIsyJzoeY+jz0TPjzOCfgH/W+Pvpx0E3c2TuYqAYC15duqGaSw3XRIRjhCdjXBk
BRjhjcc4VJPoATHK58h+zBusn8ZV6YbUygd9HuVhDnMNFBVCXWKkP8cMpW2YZ1vo
gMpX0bCWQq9PKSEjGvjF3z05uO2Vnck/vOkumFK2yZxEMKJhiCmCsDSawFiO6d1+
jjYI/iaxjr7hX1VVgg9Lk9xghjdSuc6kKMWi7mHhfcIa+k2Eik3ur1Xr/pA7G6NQ
05afgo8jKCkGJsZeSnrpi4SPOe5N9/puQM5BEJasclNst0M6CKSz42Lzov7ayKHS
PgYQOOXjIg8Cyi2+hVLLwRx5onsk68FntsUgdwpBdK1A8Rmzyiarxvl6F05bDrJT
PoYIK8AiAVRLCJEFu5OjMmVKV+3EMoYY0ETX5tE9bTOtz+PzkSv2wmsM3lJPmjcO
DMxErWcWaYvE+NhMVFLzJGNJZ3z9J1t0fbWkbmBGfvrKLdzCPmHA18agdsZ8/YYP
3o+2UF49bXPjdCs1TEmRjY1HGmFLj/NAQkxZuqer5DyxuId86KyhQe3Lzf6Rc/GQ
RkzMphkC2SmMv2ywZo3V/xesLH5dTGfoPzviDP1R29BADoM+rcbGdx2H/aLipMdv
n/arHZXJY2ful9WFnXm458yiZ9dJoSZc8wHJBusdrZEJpSP8qM12hX6HAWnr4oZc
QOCWoCt8zbMjU9FUmOGdzQrJwpEvT4c4wJF1YAY2vmBRAdaXvo6x3RUjRuyiLnck
qA6wYa2IpFi7S7kG2eNRoKMEMCclbEZusU0sNu1n4sSlzQ8IFJKEqgVrAaYlCFnC
mZAHa2o1tqRXSuktmNrpjx4Ev5QQW/Bvu4EmEbEBPXM15aAyugL8oi75+aGjDhP4
m5cHcG1gL5EfaLsNnmbD8eN/acKVIxJBGw8lQkQm6H4X8RRwiF+rGV7mHPgBFP+f
sfp8+SnjqENSZ9VhPTlqmqtq843iMe297LdlmlD780XbMHrm/yixAiDOZ/TUAAie
kHsRKx3dn829HYY+PP7vc7MIByUC1Lebcz2x7MTj9OeOSH2/eYPh6ARbCjqYkezK
2IzrqgUlvKX+C49ocr/sh9Hcid4yCI4XTTnlSMfSpxBjIfNumW/im78XrjBUDiwu
5QJ5SlUw8O+FI4duQiSaur0o/FauxzitDjYo7eOdoFFqKyQOsHBPk1z7OtqjJomw
LLfkV9celN4gtw/hTggUcGITAop/fNxa/5DkHA/s8j+rk47sk6of8KnnbjX2Wkp+
ss0nYUXZ4Ohikpzylm02j7FryOswosTcQ6aKgca6kIZlNdAW43xZ6sFCvDbwy+f2
nLpoXn4Enokx5vBvNLTMJDll5dfQaTTZvv6fljWs32H1L52KBs9yS5E3UJxS8ZEi
R3j1j12egvBlDk9KcbpkNobpnpAAI9MU75aMS6Lw24vY3xIPcFIAuqTP0CdR4U+5
TXd8x1jyChrmmROJ275iHkY6N7Qpi8tL1uAtYc6grYI55Dcu8PSJ1NQ/6tS8YRES
rUtLliJL/fCHeZKxoiMeDU4Do8bE7BYRoFV92uHwTuajHGksmZB4XqNv7TV699OT
cov/gCZSjHxhz6C2Y8/X5AdjFzMbRtrYyW56H1EMcfvWKO+ncYB50VDQMpMP0L02
l85f4nkCwCG5woXXZRdyf2XEh5bt5/iykImQHqdeKD+NHnHZq9GlPfvwS9LQor3Z
O0JMpZbc8P9lI3FGr2/JbVpJdibDIRLg1LmvlXdnwC043RRHgpC6GXfVWDrUXA7t
XM0kFAslO1i1KKHzjF6gJ4xUDF++Cij3kMOIcR2yRQbpuLpA28QHjz/+KjfU/MJm
FOAh5OEVkQs2KnO2NWAkqJjHE7i8g3Hqp1gYWDsSkrCjKvTG5LDdp6qLk2kwBAeb
9Krq+AlFbIbpzdgfZQ9IEl9G2xHQ9KfHpUw4VwV8BBrlZPv0Zmt+uXrep2y7gBk5
rzdhygbJ0K62BVdCtxb6AUCUSlH3OfaoIj1HN/vipQsTFrdak4P+5iaWr166r6kc
i4lL3G7yR63jnssB4RibgIRkjOfC7n7QZgJ/FTi3hFlsoM9goGdfQaPL12RJEMOQ
jp0mm5wxurO2EODLe+Rp8hEmjOyTzHw06z9J/2iE5VAM95j92qOyG2p09B+mFStL
zWTUGUqRkg1jiyh7ZFcbWCnAYFJq1RS8M0I8xVAI4SCPZjo/aGfEv3+1o0FNQc7O
AXoT9NFWpnKkHDCYy+T1UBif1M36QBnzi8XYOQ7y8LFvPfKfnzn9yPnKQNjtOFRt
Tv8ylAToVSHYfs920q46DYFo1Btj95GiaoZP/jnTiNAhk4GaZ0FYAE9YpqRAjF9j
cWplblX3CgsjDlOClAof5qqTA+OAQOVNEhWtBuK7zZFqbRQRVtoIvUMxMGdhQnEB
HRY60Krqfiv2BU39b6ixtjiUVQCp0e1t5pVeGoJsOgnSCCI1OSni0rfi+Y3l8ztx
5ptGBAN2qH1t6jwbbIAbaqktlH7V1iG4rZr+zPTWHwsKhPv2ysgYMdgt5zqUysVz
XA3AuJLuy7c04q3alv1PW3LTfbQTlbSAvWecQu+6QXNJB3sqlxyEJNOn3S1h/cC9
NWCmJVcB2G2t9z3vXiibzQ+dzdtSbFGmIXzKX21WqYdUH9wtDW5tfNe1tP6lVh8O
ujNDWtlIJSxIyWQcKfLq9+EYZX2joe+PR2dKwXiyh0RjFxPdiG7mZhxKxxuYZP8Z
5UcoRC11Fh9wTiJVAFC9t/Ob7Kx8XUzO/EX6O3P12kvAK388lCSyF+pG02jcC+G2
/QnLMN6T6N/toWiDedmhIiPqlgoypFwXmTM7zt3s5fyE5iD8zH64YIJUEtGQaPR3
cUk6ktAbFsLDQbtrODPEwaGxmHR5P8hm/ysQ5Wfp+TrwRPxJrpVGAe+y0/Oi9+Qi
/BpI2Fy5DHe5Vbe2jIiSnIWN8Qfu2fjyGDcPn9rD6bqnBFIf3N6iXc8LAOGkGYRN
SOWgCFJYVMwflq6QEsJrKHF39d/rUuTK/aIjg26Yu4HyfpO/fYqstTFMWQ742xs1
gNanqGmm3jUhd1AyE9z0sSgXw4SsawimBzc11crjeH409NL0BUtsD2Em4L9qixfc
fKV4ehEcAFFRAuTFi2KFnOtnoiHV1VkPp3UqPAfosGIJF4bZGGIAWABeJl1Q+xWv
HsR8kA9tuK813sEYbX/Hs5GivtHwlPl2w4OsQuY9sXEHdUMbqbswvjMaQBC5IxoJ
ROkVbOJf+csbIVqY6IzZs+JQlNBByeIhGsQ+mw54vlnCNvu+6y2Jq0GJtu+ZTv7v
Hclb3nCNKT+kky2PhRlXbI57FWubiWQ83e0Hh2HAvyBOfLmtajThdf88vnsijRey
fAdwnbx68Xi2oSoslxN4OIzkJL71Una3KjMt7sbjqYLW4Q04Hkzzu5NEq3PKPy+/
DOZug0ySsOgEvssdMmZbWis5ralktfC6GdTcoVZ1OfPsT/AiznAYwJ1FNT9ISYrV
NcB2tLIWBLh2iIoegt55armV78ix4SbLMdPiQzCE3nxP6LY4QnqLv2E23V6s+g8B
URkEnvMgyI6dUJ9Rrkn3bcEbmVX1dqYR4hK71CYtnINS7bqNwczdm1pf8G8aiucM
F1+9KsJXIBUbFaEslFShVHfNd+1WaH8vHzeQ3SmsBOakc9Tt7g3QDEFlCJtdjbZd
QweqewAzYv060cVQRe7rv7chm3SiAUrhaZr7nOT2h09tASaBODBMp2gPR0XvS2zF
zsla27amDhIbvock45t6WnZjMCzVAOCm3bFOt4N+pyezjENzoyVzicorR16XekBX
6xV/dGaPEHJs5tqR7cdY+PmoqZjoGt/yDEXbpBQp/Nd3i4OmXyCMCWsmCT2S8b+p
qRACASGQsjo6JTq1EuuB+0kIOWJabA56xgY8bdqGAo3pM0RfEARcHNHU4USPV0VD
zFhlJrKKeM+b+ASTzH8YzXAAGyh0r6u+6hCRSM0ooK4LTPLBMn/GQdKm6j/P9NgQ
MrXqNLH/5bkEpvybq49DyU2PjvB79zPt4qbHEok2T7FvTX0xQnOMu+9xHDso0W8e
fDRegMjvTND9f+CkBdpq5Jne0Zpo3ENgQisg333pn9VmhBHlhNSL5VD0/DckOANp
vWqFOVWw55w8DTFXTXINWT+xPq69jo5RO5hM6iqqd/iqqOdu0RbaUOzYsNFDB6nz
f053ejaJhBHQ6Vh4HDCPFmTpoDarWoYSxOgKFGiipMK9+ViYbLHos0gQv1/ySzrt
3jPAzlE1NQAPPdr+EBgQHlQXNqOzY8n11KfxDmwepXT1aS/fhS4wMPW0RSuAcvFo
IQmHS9n7jga0BEAp0zkeGzs139ho4QB1+1uZ84eFEfavq1k9qcnp06oDGoOFQCn/
fcKvvajfoF6JLcoKB/ud7hop133aBtxLO1m0856YcjiKsvwuzryLZdOvP3ECTUOc
ue7aNehzEl/olxAaP9adWLiqiufbQw0qiloNOlFs32iUK85/07SalT1AXqOC9ycj
bozp47BM1qtliEmCsbbbE6wGbqvFzhDbU6vSZNn21aB6omAKOWMap1PBjBPEt5ew
EtoK7V3Px1PoksKI7/iZVyYZj8dEE3+W5JDDtprBw2ZLY4ckHSaCN5rTVQ5iVGLU
0pT16uMw1wFZiyaAYyt102oGTnmDwyrysvSf4jrp1giE0KynuZALhEMEcb1Fb/FY
6/iE4V3nOFN97p4B1/4u/crxPr/wS4zwplOizFkSGctdV92NFVcfY85kTHAFZ7E9
h82SXZvSGKfKLZwVnp8OUhFvy11smm3gR51gcrESSFvo+s4diqUgVQ/2NcRLWEUv
iB9mQ36+ca9XfJ7Ys2clH+U3rZZti11KurqG71+W+SIZaDUMX8tInQQ+8ilR7ONx
BbTJmReKkkDHgmg3pRMTArHnQ4YJ+YeNVQIAZ14j4hOQGzIS5XsojgXDbPea6iu8
rFe36ilfh2SHalYYDcBu+tgj49qeny2/Lr0Qi5T2yRgwLxbOU0zC7LCbVToQQF2H
nN+qXFxwBfsATAanEkKfRQRha+lk7tjzXfI2o9U4MKzimuJMmiDKYe1+xVnZzuqK
Bm96GhAh03MMpbJSj2MgLWmw20rkSiG2Yn49bqBf4Op5moACUhaj60l8LjXn0/AE
dW/z7L4bkCEQKMDcV4IhRMQMR4PKib2SJ4eUhY6YvslzHW/bhSDLz1U3334Lcvgu
mVrOEpRVd9210OT4v9NuAZS9Obq1094cjcWM1T35gQiYviErXpaPeVeToNL/Sd5M
UKH/YwFQb7peMN4cheAtpNP//erQZpxl2nGSWs3rvYR+Et8ZKf++7Jxv4/WkjoTk
/GL9RvKi2YlmeXbOPilAxaljfuT8O34UHArb+qSHkrl8e+UZiDVhSGxK6hTRB0lL
O7Y0l0Dxebu1o3PdmqyF38GgIqkup5E2SR+PHNmjUxlyi8KI4k4R/fWh7aUffV9N
3Bxi9g+PDgeStkrfR5XwyP4Sws/aIV5D+odPQTwPDUK91I/ZrNagcd4PnRtztKJ5
TMUs7C21rpsGzeLzkFJVXUUJpWnzdCjI8uT8CfACFOyBvOd/4WUQiq891ShRBFlm
8yM4wzfjfyew8E/NHJLkMhoDVIfe9dSKMgUGfvUQ7FWfWoasm2sqTJUISXgOGsNu
6vyzuqpP1mpMtyCNZl20iXgUMVDcRobJC/e4C3peDUDGsr+aibWS/R0p1jYVcy0y
v8KnTJpK7cbxkfdKrNhJtfYr3Y0mEmdGqbW/vDxDZLudRUnDsdiDl83s3SvWddhf
dtEhr2jkCl87qwDtAtVr2HKyVhLhwoLDHiU4JqHQqIVeFsfSDVTAJG/UiuWRfwN5
styiFyTPsOPChNCTpPrr2KDJ6GuiiF0JH+mluW7DwureDRUZ35eHqyy2EZ8C8H7w
2ccydlLab7/H/FOt+npSsfmc6mfeCAQA89Z32jl+u70bamKG9islAwfzO1+zHGf3
pg4wNr7vW4U4VCCNkLb+cw0TwHgnhEf2yEX7jr0/kvzFx1WvUhaxYII4xXeBkta4
iR+JzJs3R0yQJQualVdJLkVFaBVRoRtiViBZWPR3dY2jJvXRo/M3k9nF9LqvQctF
l+9YSI+t+6nFQQMTxPeK2/375rbx6+9jlGAdDoRFNZqctVMcKrsqZbDiIe2frXYB
tgRIjHrxjRxO2uH8wJKf6Klqsagfvpru+p9n+wnNp6iiHUrEINpzPhG27vV6pVje
ZQ9FeV9mw31oxLeuxrzWNt0Fe1wSiEDzHhnvll/Jj57CeMzA1PGX9CIzpCKpOpIX
d2Kf38ZkhuODwMLLbNWVxRKrOrQXh0HIaXU4PklVCQFxYgr1S6sPBhAy5L5mtoQN
Oh1dK7yYA0YE3JCY8g2EtgMg08nCbj7mEowHcdF2i0ulKHmg00Fc1/Lv7uRna/jU
xsttdUxgmISdXBWMc40YAkjQuP+avYhfTQQJrEOn/Pm0h32zdXfBPqE6d8bfS3E9
aAEVRGFYy/opPwhf7rZ49e0LCnwYH+1yBxUIu1T4xWAP0grDGMvShvJa5fxeH3NV
q3uEpImcJwZWG/TG18E0rj65ZiiHrmMP4/SgFiH/TrlJxzFuQ00/9JsCOINvIoy4
Gdz9hgrkbbH7zJkbPBoF9jQLQ0EjpauwG2eXCxG9Y6WGomJ3rWge5td7ahoJAAu+
wRNT4+NNbLbepfooy2HKmkOeDO0++9SRxdiXauaFKBj7N/6fucAIbVW/uCIpgKrj
Fl+H24AWGZ091byWWc30xAwGp1j6yj6yLaX8YDkQEdM7yIchZGo+9ZCI9ymxeHCV
XAptRLU24R4wglmdA+MvfNlS08awTr1eZMTH+OoAAlkaXrb4JIHG4qjkhhX5pLVq
01rVQ5/H6Jsf1SWi2I+gCBumvugBUiWt0Swhn7hoZBZMbYCYFpdV8rCH6Cp1nhzy
oSx7B05d4KffQoxG5EL6VSkOZEt3AfYDe/5lIHNtZW0HSe/olL3VwPlXHBTXb38J
SfYTMxXqxqWEVkhLmnNVotdc2zhsYRYDYHlmOegrkD6aE2qcj80UxYx53b4W6oC0
wNQeKtbRkdC/6aZx+2KOndSszC5ALDyy5LFh5UxBJxZltD9ErF5VW5Zxd6+CG61p
TgG0gwex6xMt45XEbpqVpBq0OJ5YfhY6fea3n8zRa8qLqlHFm3bGR7OOrhAsu4cY
rZ9UP9BDSxdX4dTzxwU29qDaEb9yXJEXW3ldGxSO/MinF9w5POqYnncYpqdKA+VO
gz7Svv7IkhIgcZwTibxKkX5/OTW1thpUN0YCVTBlpIdljwaO/ba3+Cth//lZpRx2
KWDBuWMkPNd9XmRxrDM2/2oh81xPHFRNJ3t4nqWO0f5MbcRgSCx2DeggDmtY2C5b
DoJKETeVj+2ShmgtBb5XVUjseqpxf5qJGDFBv7MYbfibp4/OY5xViNEavgsu2/Tv
kVyMQ468P6DOy2grW1q2zRsSpup53SYDdXWEFsPAGzqW6yvv6b0RVykBg/l5szrM
3C13ii7wAKb+qxislUns+67BVnrbzEwP70dEPUods4njXj1b6vnj6gX5GcldxjAn
aAc/xekp+a78FxhZb/5hb/T/W9Srgj+YjEMn+g0E9L47oTmB65n7I9GXGykXIA4S
TXousCuuxZT9qrZSSHL+5CmUk9EzXjamwwGag1QmYP3ME4LIismsGj2PmQdeTckv
mxFd4EUXiP0s+ktcwJGy1v9tu3QMREwY6Z9pnxduccAEUwXYuObnXv1M72I6f6cL
v2pDhSUuQNqGke9o68u9xIn/4WMBIMij9NhySuXXGUazNgZROObMvpR2KQzGHAPb
szOzjr/rGiNW5OtwjV5X8ZXtbQAw7iR3Kshz0xLyqDla3rUuRF+F2sSD8srLDX8v
QEuZyE4pH5OIsQiaJEx3Mj7mk3aIt1MoZdjeTpZ5HkMgOPUV8/yBU9sbAS5yss+X
0VMCjB1w5gK88De/UCaD0dObhiDMJv2b0Uld809rehIsZ98TkbKJVkC6Znzu/qn9
RyQZiTKFKITiHaesUbs3AZkFT/+ldzjQCNKsUh+vgiy1/9qZoFPw4IeyxDRevPiz
dUX4QdNnPa121QxfTAiEwNIkjKZ9od297kM7RhAX1rl+AZ14jZchnbrEeFSqIcNc
KLgWTQEaB0gl3leUVPOfmW8CoNGO7MHeWRSPCsCp/T/YbIOfG6tYx9mZlKvi4k8s
xoUIe4QPq+VVTZLe2j0unyk6thiA7QyqSAxHE7mQ502DvYRJYxaM1KqZpwgOC8BH
Y5QLgCHWnTIbyxhawr1L9RuSVvzW8JmQ13EbhnXul8nMTaSMLMJflWZNfU8FtfRz
3pXmqtK5B3r5ax1TzVE4+XdhsTkMIlj4felkpYLjc2T9mdff9ZsSoDkjuYCqSeYp
bubXMQvHU3dAO9oa3LPFXrQUlqC1DRCDQkxCcHebJnI4tbMIWzj7krVfOJ/O8z0k
AfsB5cQ6Q8NHeHYeOnx1ptXZUDY84CRfnIfRwCeeEj9mltYbuIml3YaJsdg32zxu
BS5BPnahHVWOirozche6WRAckKanehBSmsdZE2i2rzm+N0V/cTFPNWUDMsqL9Pvm
p7s1fCwxQPa6b5RRU7KwQfVtGXK+PoMwNU1yKOQSQ0nWA+lhyW7EKFGLEAUi1k1g
J2Z27nCG8AGS2Un3NjjVvTL0EXFwQ6muC5Ev8g1so2f+swZqPT1eLJa0qGW4gjUh
eoxRsnUFPA7KkPeebHtqesomsTzs2+rWeWq11Im3suihl3QMPs0G76fnB4+sAUKG
WHl/Olm6O1fPiAA9cK+nQ8eVEFb7MwQzXcV+eXueRwKHDVSXBIu5crn06pKBuKyu
YpS+2WkGnPkoxchJ5WFfg1fyyGjU8aRkE1hnxyrMAuYBhvGj0GhiL2tGx+hVKVe5
xKRAXm96Rq0BG8x5djpPr71Kz/Pj3vK0VW2n54cAu6mfKlUkrHaisHGn/QXaEbDi
6agTYh5jjnbqHPcFqmUrIBTdwq4NyisNREDYkKJwzrWgzsVxk90uKAk2UI4uI1qN
1655RSsb2s/VxzjicvaKC2DQ/TJxD4ArZ7jsZntxQBurxsC51f6AaYHxgFKjo/Vc
+QWRPlv7T++hvdFt3VI7GrfhCT1rmPVfOaMtS9h5Nw2LoESnzwcP7R3Y6UDwqEBE
O9pqIcHsjEuXhHSDcbwshrNVQzrABV4bxlo3EQAwpDEOBTaR+rWNfXVJoSUPFFph
qV08AieroV1KZp9swMw+yysssoWRCa+AGEt2B5aFTn0NvorInE82r7dC04BeyEsG
lmujkU83vKshtkDKua2mTeVTM9pJjpU/smvjjigdTw1fDcfNyu1hJ4sjefbctXkZ
/XnRn3KftCbWbk7810DLGQFZrd/lhzAxEjQrAJNtVhhzBPDcxJ00cYGtiwAwj9Sf
aXFekZmpzBR6Xl+jxlrWfYPdMfXNoTFQTlbCx5JNdkdHcTqfO1E8RuAJbNuV/P4+
6IRYMY2IaNEXdxakijPUy3mRn70LehYI59vWIYwr9wEi53ax9SKvJGlJVYwzXgdP
tbB3z/QjyuxU8HZq4oOem8V7jJPTvtHk1eBpxaIKClWVqmnCyhNLUnny0JPs23GQ
/3W37HWNGfScEPSfK+96ksmtADj7IvHCLJTgM/8/OL32YWfGnHHFCXGaEgJzMYV9
3f3m8Geg31st6/skr9BjsZYw4dj2bfOsK0waFSMEDDo2kbsPMB47yVcePBJTtRxz
LEIBWWZ7EKFThHMzwPCwbHCihr+pAun/i4giUwtCurkv7EELv8op7Vg6G/BCnxl+
2B+l1+70MgWbtPGCoKDe2HVpUFmK22Lu/l+g11mfIqsEE3lBMZvb/bN8dGv1gkEY
6TLBGAW5G7VPSbHPggQcq0F5kPB4El2tZ2RYS4wjA/7g+UXRQlYm5D2Gu7mlHvgz
AkEgPOnsKl9MjRHODFCbuB8aJ+4tX93V8Vrq+hZoFdHwwFIH7AuzXVu/iHlq4Puo
Q5BpmmxENu59xeAY2AhAWOf63fzFIRNXrSRxUJJewsHN0NlUmZWuPpBIXWw7i33M
s/ZSZKu9cfeurOMAMgENtMl+MJ2bHlz9o6Kz6eV2w1YiGxzlQib7DSkdWQ1GrVnF
SMbQShodkjzU+y+n5cRX2W+H35QDqONoP7nXctes+5cpj+W/P/cZRf4x2KZgf3vq
XRzFf+0+3/zBHpSDjQhtgejdOCf1LtBwaozeP6acfGyTvrbEfP26ew/AltCXB3TK
73lM/s5+6K+vYBQ+RTHJSQFBd4V5MZjIp0CPiOcF8Kb6rGUmJXrQQSNWQj/yBUdQ
I9/bPdgkPELgAqQi/P3Loh+qvk2QkcMKNLnlZMwEx6z2E7gxj1X6vMIDJLKZ60Zw
9bViV4/gNsygF8eHnPPme5NsAQ8sPtIHz6LF3Wibw7jq6EffReTmSaSV05xzG/Wa
rA0VGwoMDy390lnC8E/9t7QYTu5f4bo+1U8iC3ohsD45ggJxy+R98CzVq8l3ra5A
F25Ksx5dDXfbDOQjxM8PLQSXTlhSjuBE3Umo4pJwSw8rOWx/C1c29pyDihvnBKmo
T2j1UyFJOY3ASd0rX4w2loYMQ5hP3BeF42aNy2cR5PF+p5y37uOgBHbkYDI/GQJc
RQ8tlp1GLVsm+RS/lyXZYfmTfXtDB8eGbO3dnp+n9xQp6nyquR+CQ9iPMsODo7r0
HNJZZ4pB1rphbZJKtPesxOZdhdgi0ExO35Cw9WAIQNh3GzK+SOMXL9qFzshHxmJj
LlnY0Q4l+bcMxEczaF46Seu0WxTUrkegriNKDFO+BNwonPbehdH7KwYJ61WXm7sL
nwiJr2rDUYngCA54S3gPNqQ3guOZq8l7TLcnk1o1AsqRGou8G39ZRPfh3rpFbkT8
Pia8mNBv3+9iLk9y/O4NCcowItWTzzdzqGuSahoYiLiknyKXLcrCuQvdH2ifqpzm
BIqeMgYx3DmVe/xEi0zCZNe0R+ztazIKYNtT/bgsCS34VFzf8zmG/Xynzk1HhldI
89tDNtqq0Jzr2w3sGfXfxs0QIzXnts8njBTJsQPvg4h9vqi6y09Ft3EmGGQOE2v4
7/+wGaMaLHSqGnIfkx34FED05S+ImRhKh10yq429rop28GpVvw2K3byZB9VXEBAW
awnMrB1Lx2qMwkALgqXadXczl4RhA1zx+DYw+B3KGqNkgmAX2VTs3p+GIgllnzi2
RA8udvmKy6PPemP4xceUsXscql4AERpUjNErOrxCD2eQh5tHq7Qe/uZXzlQq+LVm
TEsOdZFKgkf/LoRb2a8vRem3zy0rjo1lfvIFEGVYGhv7xRbrtv25WCEQ2eiTm4uZ
i2GwzhGR+rNb1NHObo5MmVbuSNf1SHDpODpJY41VNN0nnjqQg9F2qQEVEw7uFDiY
hS7P05c80Xday1fT8X+HRxLsn6SS+Q1BLCHDyC1zRhYTlCXtEinugl31W6a9FLkQ
IOvp1GRFgpIE+9HkuODNxhw+CFkVVKrrXBFBl2XGn5W4VHoI6Ap+N82r2tceJXyx
wr7HVDv6aoIcbFuJFtqGdkrmRUo8B2ulH6eLs0PfDv9qn2zCh9rxCx8X9gSIlWFp
riGJ0zd4vZoMMKcMjabS2MbeYa/2G6fUdRZ7MsAbzMLQ+g+pzyyMfbYZ1MsQw2Zv
buzG7/K5L5gGUrr5CU9Qm8UsF7gH0+yzkomVHxVtRPrMoaPc7TahKBUwryx4zP8m
GH+8AncKM0I20e8HGDpwtQDJTOGFs2wf6UqtTa0lelQwB+e/s43peibOdHMAV0JP
OOcFZkrnDLXtvGIKyavtCW3LIvIHxNWci3/VUBEZeUj0WfoMoo1q4Tfx7Yh5enFO
Y96RewrupydOGzADrKK8cvZsk3zeHw6/EXibyLk6d5lptYt/0vLOcLbgjBpdRqMT
OEzT6MSmCTFSGMRg43HofKFmHVTyNsUcmpMx1+Pxi4z/YhBnDcG2tJSPInzZvezB
Q7to0hguqJ72A9fKWvUr863P9l8syjQectlxk1L1EdJAZrgr5qtHvknQh0DXpzta
2vN2eO1DcyFLkxM0BNfJeQdMnpL21+Qz/bm2Ydw6Z18jXWKBws2bOs57qqE7tMDV
FGdCiCzH/iRYU44BhifX8FM07Em9n4R97DtCtnfu3IqByU1VziocvWWBymF6oH39
N59TKjtMaDvZXweC5iwDXJtOjRHANrZM5edWaCadU4W0trrJpMuYDlFIzPlsaVrI
kU0VmvUk8TaHuucqorHtxvf4YU74bkML1HhgDqB6LdlwpgWOGvnggtD8+X/Ft+cO
aQV908JqOPTvUPwMACsHkUvfCazmhoFzOkeOOVCG9oFj+frMuEypY19L8ZM8cX7l
dYYsflklp6n4uF/M6x98ZQ8KqdikuUzAWmstKccpGm44q9fK+cM5x2uraj5O5glS
NiSUfnrGOxdMeNwJUUCpg1YK0JLBi2Tuo1mGodem/eToXcwGlZ5KroR+MxCRaSzN
q6w+puobcuozrOp3iomiFysaQuniRQk/Kv5AC04K62bJ5V8QGRiLlUfW+tw/xaCC
U2rlg7O16m9wjjfEsHroqso5FiOyYf3LDIgYy+rQ5LJdnEsAWT/JYO3aTdwBgJPs
sRfjd4ACtJDQe3pffdJEK7AWR6212aS0z/C4WzZqmPwjZZuD3bkaADHhrZlYlASV
M/X0t8X+weNEjliD/bNVxZNBRWG6sps5/tnk4Jz7FWt33MjqSSuCpH9e0A6cGeAQ
cpYMv9DfKIrCUGSYNQY0xM0gaVe0+v/B+xgOfq9lLLW5ZgtFCLZkvkGEU0hKLRd2
s3u2gu0SkfIP9jJP1NmWV8impYgT46H+SO06vEpsSkmnh5okdezZsYMRFjdWw9WW
N34bm+gjBHWs519tcBMnOl0/a/sbxWaFbNI0N2GXvrXQSHgywycd5TztFOXYUZ1C
9+/YFUNnnWAPtUJOGQkeAvJj2jDDBwtkQxdhoEugFl0yBqI3AAHLp7Y1fjnkpuFr
kwNZEEZq0yK5DGmgWbstzXFBZBoCLwzrV2cEMZrM00Sm52Q4KiPuQ/Di+UO1u04+
pFsQuEabZ/09nhq1BSNTk9dXEykfEW3BqJ0c97CYmjg5h2rlmWqkPEmnKnnsokSb
Ur2q+TL/Pw4TiCi0kNuNXR5NkdNwO0BZh2eAdiqOce5HgHigFAx+6cDaJsOQqZvW
EsFGpc6MofyBKRs6rQqpSLnnOVHIq/3/3VuIWzmo96+uAg7QVoH0ru25ZLrI376B
Hn7LtqJovQcLUxgwRf7MqrxS3iHoC0VSoBnrCw4kOnibOLnbotW6eRXYXpVmWU+y
OeOvD4+Cq7vGSSkfFi86V0xb6Faszl2kPioNX/ke8MLHUhAZ+alovwmEBqMU6Scs
T4DT+LynKbywvXiHvu6kcC8cgTFzXyhS7GB9VyhwPb7+QtIo7ZYbFJsMhLvFxKb2
rKV4hhN4iU03tC/J9uFcYH1jkS7buuGMoDNQmcxkt6uSCvz/3WcX0Rvp8Ro5dtB3
Wnr7iL3DmreE37LU4o1RzqECqjEC4Z6vqiUPbj5sav9d5RGxkslF7Wxs5RXeWRnb
HIhhbX5/BOh7ubGaeLS2mlUA4p1UV6paGxYZbcRD/3gzfyqrSok2+NMo3fHZCG1T
4xc+EJYry6HBVdALwAud9Y40TJ/l16CfnG0XcWVZMGNF36g9HWKOCOo2FQtj6sI9
8MLKOXrLiiXLpTxlTu2+DGeYNWgZD3LbYgdBw3dRToFBtYN7FXqLyw7Wc2oXPS0C
WmsleMJnEbPdPadCxWkgigqaQMHIqJaqvNBCa0aQeKqod7s6ppnBHcUbCFd6y65z
EmLBXwwHvz4cEhYfHbaAo4UExc2KM0oLCi1Y4Wa8em+wH7sgJxnnJRC3vzU7AvPg
AcAOly4WJBQVsoT8BzsxnPXvhpLiqRsZK5Dx6zRz/tm1VdD/4HpdcrsVyiOeR5vW
p5EqKgEQHH7vVv7HWxwO+507yIRDLJmYtAv8XtOesO5TAtEIig+SgcqnlGvu4IDM
q6e7TkGf9kH8sTeTSdyIQ8A36ohZ0OV9EjONp+RcJYqMj5RJi+DkGtBVIdMOCz72
kPzWjch0ZW1dVatVyre6WKu5/DX+B+8Z3ZMNOW9ltCb9WVF4H0Ww81zvj+VbEd7W
cXj1Xkx3Gw/9Jvgw1rKkEYT+5dg8cqR0W9Z6aTXoEl/aztl7hw0+DT6PUtAz3njM
qpu0ZXB6ZagGibTv0n3VNrxxD/s/0iy9U6dlxkzd3uSHA3tXJ2hkaYgQMSjBijVg
8jzgrMwBpzvIMUHDK4hom/R/Lah2Uidj0vCJifvb0z1GbpAdewc4xxNbs+jqazu5
zf/7P6TRTz4Fg8730UiI8FzUZKZmoIcMNztlyRvkGTz8OrydETA8cBMLizFwBE+d
v8IsUBWtyCawEVAOdcIb8ajvisBeTA4oxnkEwOoBi2eGxxBb8yAk3PKIgVcqAaY0
mrlP3b0N3bc8xbXi4MBHUAS33PeFyH9bE80SKDgHJiKjms4Sct5v5pzNA7ceV7XV
1aKBDDEjECdAWWTUnTPc/YlVyp7LTImzfk28MT4cTjbiHOIP1RnhuJoV3fhM/oxB
Wd91OtXw6j9Hqv3a/BcZT7JAEoApEVPagr+t23FLgJ7IYfzmjRT4MkC9W3ru77v2
odsHyye+AJ90Xi3nyS3IVwuljnyzS/93W572EiqsEaexiZjrB3s8BANm6yEXklYY
V/ic6oLc8tgalRpDRc60fI0BOx+i4EeldHmepHAYcfYI5yRYdoQEgehTHod8V2Ww
p0wNlvQpDxWcGPTnzl4m6c6Dgwt0iqOuMjcqaDln8qqW9HuqPEC0kaGBaXpoqaMQ
Cve/ej1cdfgtM97d5ytI/2vlVJ9aPqswMUxgOpHD8MrA/hI29k+qcVYPdhNcZs9F
TgH3G0c7K3TKs92JlnrF1gnWKonaTL8hj3aiVHnFOUki1fifhpr7JD6uV1LbAe1k
TFR7Pd85YWVyWT6OLbpMVR7rFYNWPdDRXQITNPENsn04ggpfRFoTAPbLYO9GJGzq
/iuhh1yG6LyiJqYchmoU6P72wU3xiUu99MSj3zvNnpKWzI7AZNn3SOUEsiaqp6yE
YKtKUEMZ6EGpbYaPyIETkhgN6Hw7H21wMGuUhWaiECOVIRPB4Dw0zsQPUgD+xWyu
/7rkoaJMSQHLA0BOKP5TVNAWom9L5SxU5ULWonEWTsfxtEhRYr6ekB9dgaGSZP5X
o84UTkXtXcK66OjwVzEtGxZgzuZzJFkI8JTvE2sbqs/0asMQVsum9nYXvtUhqMg+
Eg8dGCh6GKrJ4D0NbWgSJ6ZcY/uKJRn7ho54Lznmp3lvN286TfLo4xJwfBlFiu/F
GGfvyTEmnqv0wpN2NNL/+KXDJvVcWxvP+AJfscB3i/5iX7A9Nm9nbw6xh3Ph3Itv
8/HxE//WUGY5YAtAZTUtM/HbcGyvubT7RfJ2eo10r1+/D5sfoopUHCtiq2wU2xz2
V2ZbL6FKgZMkEsdlVa8oxSxp61ahOvOHriRdxxtyBxqh2eHBKl27TSL0Pir9ni9k
oiLLlUndWqaqmo5ZSn9Fq8F4X3eJAXtVgZVd7+BdC8TeOoiTxvErz7rECtBVD4lC
lXpArLqN74FmjJYMO2OIZtntUYYy+q7Gf7rI7fO42axKNbeegUSj6+Ab92jncjU4
XMWIdk2J9uEzX4TtgkrLBJ53wYCChHoXnVK+nY6n751sA5xOyEg53wXHPa+P6A1u
fnMNdfbKByDR0Mm5vJhVQWmVnpy2olrpCDKgwV91XX6a1VQ2rgVyOiW3AUUJWVWn
elLmxbSXhAR0sQRO0EcthWZUopu+lW0tnPWns47Rec8XLhepgquc2gQQM9DM89wL
UJEeLV1upIDpNoc60XHT1kfTbnqT6bhRTclpE5L2FD2XWh8jWMYg2qf5OZXoKZTI
/UIicYo3otoONXax4uthiu3k6C9y2XbuVfkamn+q28iYPJS0Kmutk/JFnmPx7BKO
7hMw95oybIOCpVFppLviYZzv6frB0orFcxo8RWbjWQq4OGBfnym3suH4vABZG4KA
sj7ZwPipI/4Qdg54n6RufmmorlnVkZ1M9K3aiUcYfdNcS9oi4MaO+0euMIAZLOEE
JKg9PV8ldpILxSVBYpMa3WLI+wR2vw00tCevwiTeLi2C8RAbFCXnOSvgUwAYXGtu
wADhGctSlfDS5MT40y+C9hbmilQ5+AIis1gDC8/4FTkPEeOlmyPnDE5X3CBWOhqH
StRXDrDACBsevkWKkyQAK90I61Zsb9DNBOTKRMiuQ2EYPs2shN9RJWASblIBrZT0
SKYVepzVf9UgU1LkL5RchgsqQMzzayFItQMJ5sKW72UVKoK7pcdEDqVRh7iSh9AG
guazZj4IXqlFBguHAv9T7JR1NocD/x949lx7QD2rYhA7NNifv6eF3GOT1VoWpBr/
RAVXKUIIHWZK4SqBezy8q5M5ZFAJGkYdjTBouof3GvYpkE1+DAzrL1Qb2ZcsYRL/
BNfvRhtlxi3AKdNfoTmG8MY05NQZ7hQC6eJIPIFLlceGmjMCj1Nfejj9meNN+i8X
MNpAxeFd+DPKBFGASFmTZK7qdDyCQJs/c5j3KDy+r20LMAEjEjK7N2RxQAySnI8+
mndHn8wGdzMBseHqGg4N+Drpd4O5aLuJ9z5aNOWTme6pRzZF+Ojf77oLg0jsCTmp
Lf+yRXIfs9FNZO8K7Epdnieu8J0KZ7BvvINVeWv1gxhPISkCMbX+x1AT4JZXqUAq
HdU5l6pA54TH1oCxjI/gpXvz3CY2ujgAdJz4orOu97SqPRlP+lCz/mT9tNYFEZVp
rbcbjoywK6nYXjj86nuD+rRxxBFhGKQUDAotRZhGGnhovPWkADDAelefD+EKZa4I
1U+PZknSLWYX+iWRWmctUXtTolQXdXP+F4VeKAtBvuJg806V1Rs4a6w7wptGsi92
KuBx4d+UwKgIqVXMP6AAjGaNjbGDAiYF0cx/lcfD4ARZS/XU7PIsSueQPFPtQHN1
eFNBN2QPlnq9pnOws3U8Ce5YUazyqfGWF6OeQpRb9Za+Ltpu71YloCirAKxvXndw
vtGxOgpEQHAN+K2+fvwfUQ/b6Srl0gR4cOZjDlM7hv528IrXEZgTzbO6/GZdprOB
YC+rcXejWmv9g2ofBS6T6DCefARiGJFQ8+Y2z2qgOs306fqm6g/WSnuKDSR9YZ74
OWufC+g3bAy324y5aMAyD/PuEBaLIt0prmohWW/9wBaWPJXDAZh0WDBhDJsKEF6q
j/qBt+cnguHRdyQFA6V5rzZOMZ51S5ek/SiOXwDK0fvRyZjt/dbzbvSjMkIOb+Wm
KXKVrI/zQiUUC6c2wZ1xEG2itZNS56+prXyTwmVKAuOqzZM+g2Tnco3aydEvKp55
yWMZEsBoophOCM485xWb2JSeyfjeacWQPBpdS4zIinZJ9PUK0p5s6sdDWA3ARiCE
ewjkkxLp9+RW/PRZhjl3iEhKrUQ4fM0IB+xBOONdIMlfBcjftsMYYcdrZSn6gzfp
Y/avxsqlMNZp0FFWEPCDnkjxnJJQ0UEal6gykfJQifhtp4xIWd2f9adTnGQE31/R
cgaPLkDgECDnTZ9+Y+Omnqad2HzlRnt0CPR4elvIBUopa/Gn8WHIr2C05MI4UTOd
han1kIE2idzvmHM1yWvTO9cqHVGwjRrbrrVEDc4GnFtuKJi/QEGLdjpYGwSasWl/
P+cN3oTbbuQ7RtFwwNXzmBInuDAiK9RK1xaOWa8sUXD7SY8ebcZU/Bq8e1jdSHqB
5ik7yne2F6SqhK5RATcvxygzp8ZBb4LLEMBJaWtQm8edZXvI138n48srhGnD3npp
JsipGVYaM4SyXQIiradGypRQJu7dXnJZZXiIr3T6j2/RPYochmu0h8EaGw5bdgfz
J6OcySg1DUH6lca9q9KIWwws8QHl7FJGVvC1vUX0CCrouHOX7zOVW68vb06cU18w
FJ/IUrqYwDwgtQn1FwauFNuIgVre1yqVqAXR6v3VWE4XtMdeu+aqZkftJ65AxecP
aZHJrAvWRxv8XCo2sv7fh9emVeP/QGjguFA1Oq5bHjuc/+GSsl5x9+KpMEiCzb6y
yklLxZqgZ6awunxyO7bzx9HhINRTok03zDKvVYTLiCTO8TvZPguUKoNO4X4vQ5qb
HlHrhGp38onX7wN+WfHWNxfGqtAbWAST0Mc10OS91V7ZWpSiOaI58pvk9Co8jK80
sW4vMKJ8mGHHkvgWA52EnelIDDSR6SIoaMnxXIoYGNeuukhKS2qY9VY3Cacxmxpl
mr0DUmZ/+UMXBpVPQ6Ym3xU5A6B2ETmsxSdpTdBRKtRiLuTTlmksXl4NmkFwg+v0
M9+qI8RRXbEuvAM3Zw+7Qg+QZue5Eseyn745H194f1qLgaPcEqahEfXbzsj5AEcV
3KkGmq0N+XF+krdGtY8pR2iD+49gx3W73BeeBMOo4vXi/Oyrq9eJ+qf5RCx7OJwK
hwgtGwPqqM8BaZJqx26NXwENovwPlcz9UC2ya9VcuFUc+MshCsGQqtKIw1SJMVSw
tlXXDeb/2zrJfOtWZBZG3mqLDt0UaJ8JYJ3/gwBjLxPRvPVOlnyxVje168ZagAFb
RrLTRHxiOxKE7RW6GPjQ9Z+Orwp6byxkm0jrNrejGiCkD0VKbCSCCuf6WL4G3vTq
IfBqIt93kXSpOPKy0PS/3WtBEWdj8b4QPmdsm2RPoV3rDrA5qrU0Vr2dN2sbhenO
VPYtMf0cu05cfj37IL8nx0IMRGzQZqpZ5EYezRCfdMlWxJnDE6CK0N/IZCq/gRa1
tXyp2I1AM2IZCKhkfWP5w8+Nw/i2xZidACEfPAWXgdV0Ym+h6NLtkkqjllvPHvWl
AvP38oNLB3hD/t9pIMfrSraCRBcW9WmmfJZxJkpqLaqfL7eeEKJNWjkV9+RcOlZh
Uqj9JNVTNnhx672Ek8twL0xhm+rh6cSiezqm1fHPpVse2HUFdHZEvDZMmOxSpFwA
AHvd4AUk7NQqLbSsgz9OBNns9au1+UI9Lpsh6BJ/zogivIV6Vg8UR4wWPjf5g9Zs
nc1EzC5cxfrvg05C8bvB7Lj/U8pG+3i5en2hHYsviQkCP9Od8HW0iHiGBNb5nOyg
PURWS8I0em57NvYg3jHqK73+fEtaxmMRFOgnM35ijdtfSDpmGwjzlofk+sExJk05
nJPqoXasYTX0u+lVuJnoVcYK1773STSXKQAjnFNB0kHa9iLL/8W+ZReiPiizDjmD
s15JJ4C86zPxyRG6Wu6EdBBp8jS/75ZAwmFVP4p1oX1dBf3Ax6r5+eL0jv5BRKQI
SDhad5Omi2PaiXzVYXeDv9PeZJ0+mTnOetA+ZDjrphMflTni0JRmweRItbZGrU9Z
ndGcs0okWAAAzwLnmB3ye/I66OOQeHsHYpMO044s+BechtHRpqNXOlkZXzwh0ZGb
oPfSJGIxApXO//Jm34ypfo50SPlIEjyUEQgGE+LCKTzyfko71t6OCgt/omfkC447
255asxdWoUE13f7FsMe+L8Dt/ZfnYPcuqS30AQ1UhOZSzfOL0wictTmUBPuq58Mz
bM14yOv8kQlu9gRHcyIOJtEo1u6rjVnWUBUyTEJtaPbtsMPdQlcjByzxOnsWah82
L7vIxcxnCOvbXF0qHiW/FbaxBWLhtabv3zcHKP0vDOeFTu3xZXgKQVdYmPqU6bz7
Z8njiakbSO/J0cHgeeg9xKaI2T8MFxx1BZ2FqrYJkz7M+ZzuQrmJ61HwC1pi1z42
3PD/uunWvetGSGMbGi7DUKDZr6tWviw2nhxPYngWUc1a7CAP7Sz0t5whkHoIRtFT
59jQNxMDSCOmjALQUXGNmhNtYreUZL0tkcqL/L581dR3EUjxiTgZtXt/ZBf+E6Eh
nhMFvj1Fpxua43fZS8iRYLanR+rP+KAlFieMnjMXcdPPcDKjw9fhvO4/NBol823q
IlQXiM2FwuyZNBH4GISAj3enJFsnRVQ22z0zWJlbm2fzZdG9Z8A9W1lwAgp2sRck
fHBIzouy678wUfNosDNHzvayFIF5JeI/scdInrQnmT11rwrYMs/CoNXXiSFGK+Cx
M8kTF8osiMOxs6DMOtFcaCQaFZTa6AB/9h12lwl+eCx0Nku69EmdUwS4XkUbK2vY
1j9RM5DfZHOwtOJthJjdnoiDVttQj7itRmQSH6WgBlP4rXFvFcTtDU/AjXzvqCSF
hqn4RmkuFxNDBPLDsU/EZU15qLq5wDJwxsQgp7qAoOAi1mrOjMCgR+jk5la77nx9
SlNzUAuVjSCPotFqRDygct6t/VAlbZtY3rfXH8bMwN96r4ZZEGfeB/42zoLx72A7
v1iUSISNReTZcItI4/ZSgNjj21b28uB8Yau3zlt+iAUfLcUUWluI4lphouywtrzI
CviA8mkcoijo52vyJVU4sHSJcjjTCTehjDuwi9snBNA4Kl0Q34DZsCfDqb8WNxHc
3+btJUJkkUeyShri28pHZbbK/Vj14pocpujh0WcC8nFGufbFZiuv68A6qujLizTQ
Do01tvWWv5wug/Rj0hlldmeZgzAvPEdsNZmx9fGZQaHpVTzgnhjWFR8TnFGZNWDx
Y8aQlGZyEfibiqAkWkRcLAAsd3yAeag+RRCTDJDNEyG8OYgdkI7ZYnkXPKWVXYh3
bs+6Tze/Yt3vXzsF0VZImnEK3ZZElfOpRJICqcdt3Thbvqw1aP/F2Ol4EuxjJZ06
4cHdE3jP7ultoJ9l49CcN8nP7dyZd7Cm0e3R4RhCD9g2znZ1WnsbRlSg7VYuT7Kt
YD3p4pPT/3UNVoZP3AJIe1pprvFoVxWhQwpb/joQi1ZeKfGtpux0qZk4GUT+a1Tx
w67fl5qUQKuJZDHBeJjX+sjwQPXlJTiqSV69BN/S9ubcqr4JqX9VB0yOh6e5x52A
ftI00wLV61pc5m9PYWJTMOx0rUR+rbjEzoAQG/6Poplt5fktLzkHqiEGByaOwwXN
xYmZXybRP84t371pus+4dltBGe3I3/l57mJ0T2iC+AQWp97E2Gs7JFLk8t1ag6lZ
iftRO+A6TrW2kIeWgtsDSs+3D8TOsAjxQ0wIFb+5YO7QcJTubJ5NCGEV/lt5mYd2
t+yPvshrodIKhgNUno7X3Db1uVd6siwK41ue2twwfx5cWADc9lQWJVzcVfD7QFmO
tCJ/3W04NGnhWzhHEKTCUbNSy05CfrtFm0PD1YY+8OrxiMishopDbLW1k8JH+b77
3owV2EjCMfa1JvqK+JSGFf4rPOdubsVSHpxKnXDSd0JchR0Dfifc+PWDo+yWexiK
QIgIFkOEuIc8p3enl/4hZfZTN/9AG7EicYqR5nBIF+HE2umQocTPOR8WKxyxsgZk
7aiBaJqHBsUdkjgwnvszCCAtCDtgWPCt+XenPtUviOmrhdmDLNAmyuv1sEGG4TD8
ghP1HUGpFuxealH3gzRIGcAG8bavZ6avEFWYHOl60STNkMbqvzYoRYjMgz6TKTu6
Ekwx8JBnEg5TI5hbdn/7U692Q34qpxpuwgTSTQECdlhIyAOxRWq0hW2LiEDLe07A
d8mFeQtUT/gc6IpWF/a1TEfR3V8SrAyMci5WaXOioqwp8HRx+uXXnA2v0sw/sIei
d4povMHV6zAJOUkX1TH2AcFZ7Btt3kKil6BRWfOzukqy7E77jQzL2xJihkRaA5Es
yYdNBQwmz+RrvCr5HR8JRQsL+Awpf34+7gu4DPK4AgJoKVjtou5BrJt8V2UgiFVd
7XNOB8G/VgI9fywW08Pc1/s5f1DdebUfvXjytmGDxrhYaJLY1uUvkPeOth3M5B8s
ZqVf1jwvPA0nmH4XahHnwYFGm8aBdv4W0ju5gG3pPLSCqK86pjeW7efLL+sHSP+z
MXqS6mEDGR2tbMdkfY/VZGUJhHOavX6E512IDlGtLqivy1gtdnxb7+8fLmWBESHi
lumroFq7ixz8pnK8kvq26K1MEHiDzw5iZ0UQGqRH0zjlZHDahJs5FgUOlJibFULJ
QZVdzv909XMGAttuhBcJgtnH6V9GMS/xDBroLT6cyn7pjeiXX8LOrYpMxxML/osx
EGd/7KnTe+ZFxBe40ejYEqsX8irCrZPp67cUyxJq7G1TkGGgpGBTQ956dCuUymGo
A1O7Tv8Qin6pkbkSAhIPzmojYHMaidbeSL4I4dYqb5DUgnXtN+TKSWGoHMXyvhdi
Mmok/06+ZDSVbONs4IGBDEyMHH3+rm7dCPtj9J13B4WaZtlle+E3cIsg+NwolkxJ
+PfYXkxboq4emJBBe8uI+pONjWzwRj5VK/OOjhJ4s8rGIkOr6SBOpB0SZAMyVrAc
J4zWCmdr/sJH4wS1l+s2r1NIxXEEARBnChCzPrn1njpPU347bUvtKUVyrzXjcFAi
XuhOVnnTqNa5tNiJjDrK9E1L73V+N/DyYVCLKaAQQzJz7jvL3e4JVnYNRSlEqBLc
IiceLK1cw3wpFlDfGkXivwdldzW730kVdLHrJ5vFAIZazCwxYwuLJXgFt2WkwMeF
SWlj3Te640T1OumfNZ6bjiGXWh6EDVjGGqX9DR4EECKmzCGgVgO34Mr5U8xfS76N
vZg8FvyL8ug33/uAUCnfyyfXcERuC8ONWBcV8BZBnJWl+WKbBzoffxTQwYstdTip
HNwWMR4fV5CnWDIeDqzWuWGdmdPb99apO9abapOE8TUVDXhJ2aNvuwDDMuFR6/Oo
A8X+rE300YopuyBImDkEHX2h3n5KkCRIfEDGyr6I8V4ut7khpfDHG7IRpUUnsS9l
r7sxMWEHZlnd9mVgwB2BuvrShkEloXmsNp7m7PyK1VPz0Il3+3QQ584OMHJUovvO
UgwXRymPNeAL+jsinROoL6eM9PrJhDjhryjir4pIqdjTO1SWy/GzvRfeQsiZXbT9
SZZVkrVCv0dpgZuHLmfQY8l03bN5MRRVLuYjoIzQU8xCFclawYxwlAQwPy6/jOv9
uHXCYvieCrMTmyzomYyu18KWRgxgr4WKum2ZB11WaSxuw9aH8J60yiPqAMZVq2t4
9Xsy/Hq2Au8w3FgbwYBDlw==
`protect END_PROTECTED
