`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJVbwb1HEisYOzOy7kdWE7R6CZdHbRJDKOxfGYwpX3bZlGUZIxeHJDcsrHT1tW5H
tfH1BDhsyLRMW4PJde+fy54CJQX8IVeNvEXSk534/mx6DDAGc2svWxpNlsg4WmyM
JCv2gTsF+lMSEH81bBwzP8OKdDwyfIWeaKR5xBLqS31OJN696d/EAB2ai1KX/y7x
lMLJQeGYuTPgw195VZY+4hwKJjd9KVYsnkaE23vbczPJ3xmsOwboDRc7Az0vxxXo
Vm3wdV8RAsf6Qlw97jCf52FyftrRIfWKCBBcwgCbs86j48hrOVeg360xej8kYlaN
MaIKsoXaMwYl3wlBHKD/3y41Hxzlvo/RgtULuEGWi9GdYs5yP1Ju8cIHoJpM72Jd
sKkFFT2osLJGZCVNhFXpG2qzT3Jgc0bbevL36ZKYvNLLc1YOld62bDDjNtflvKLQ
B6839lKpZBzGyg0O74jCPsGqD12ht9Jr1JhxfI5tMWRwV9ZecgO+veg6U6u2AiBF
uZXFAwOpBmzlUoD7DEvyo9BrhlTeMoMKnnIdwczh7ZA+be9m5O+qULGWwKluFUo3
Wyr97pwWGnS6yeAq2s2MBch+SwfZv26LufgTM3fPHJ/Ou7Fi8n/Z9IApx96NoCR/
+ww2Zeucf9dfjjoqQVBu6Zw3P8UpwVnzPsZJF3EPMbPy5B0fUYjgk+D7kn8BZ1pF
PBZXnz0XJ9UHNXBNqXQ8s61l/SFOhhLXWEqrjNWnXBUmWRDvLCDbTsVPNRj0pF3m
oKkuXWpz+RfwUr3LcxkcOB8AuSZ9cHByeEZM2jT7SQBUHs/c5Fsbp3aOBCt1lNUm
D8VSMy2WBXDdKXp9oRRiynIB1ToP6iPov74xOdX1zsqG/buSNZcY2ITD7CYc7g2x
hUTuBjy4sTZSSjN1QIJsAklHcEvXXQESxBi6Kvs8xMiVYOKX0dH5UEhY/H8S6UKe
uDKb4YqneRc86aQ3zauubOYj1fde0kTHmEn19VduXQMGg8Ca9p85HIOBI5wJeNUF
pCdgTrUlI0pQIXxAf5XSyF7Z9/QMui25wsWiJ87tYBhcymcEa3E1Id6s0TNOFRXs
5XrcwEqf4TAxiftqvkmVAg+zVJUIgQ6hOZMvtnzCPooK7pE2Am8+zDwXEXMQSSaM
vFr8ywK7aAojq1ODaGaMddC2AzJaFJBWCvTmfsjQ3HFDhFxlubtWA04jYxI3vwQF
U+E/hencIcVQtAf2gN7lN6xBMvF8IyRlf3QOk4ne9XhJoTFVOTMAIpJQqgFJALXT
hXFRo/U0yT80UnEsQ1c9eb/Bsr2nfSXXhWHZFBiUzB6CWJjjkf/pydVAZKSwQAIQ
EWPI/qa8GeBAe1RjedABpVek8UD7y9vgdWFywgHcpxCimtaYkm5oP/AfkwG2GYWi
0dTTNj53I5iH5sz6nJOrDYNfwSWwjBbWNU4zMC3fwCnZWuBCeE2owwUtsLwIn8m1
peHO0c2kVZ5UW8+Ov7blg3tZPHb0x6lahCiLWDnqnHQ2oH1lnZ/2hWkxAfzcOi3r
7PTYznJca1ZgOdq+mfztLgagRxtcu+P9fiUJvvivNCslQX1o0tFlB74nJz1Ry3vw
BUVT2bSnNrxrOhTvRmBs+twZNiBLUssoCaU1tW2NkE1KThn7RObH0bJTNjPRNMYP
9L3AitHIBOj7ZdmsD6fk0USSQDGEdNuE+Z20Yo4Y5/ftPsx4C3pgyRZ6dbqeRg3m
OxIeZcjEkon7amDEh5sJxlBdM/k9te7ORwBUuHwW7eaNtX+UZqTP9uhASilNCb9y
AeqJ7PjS6xraH8ktsKqcEOAyA6e8nWBTC+vpJ8RBO+Wd/PxPwrMLqWOG0UhSGgN0
PQUJdTGzdnaGqSPDX9sDp8E23lAH1W9OE8dzcSAP1+WDn0+Ckc8WU+kW2uiFc/so
BgM9y0K78NfJwWuKAxIO2GdWQe7PDB7RX/txpesAMulidvxN7+bZBqN2FgsYWdk0
zsLmMcHh5sOX9bKK9LK6NdRkjBxoq+Y/Q4+VEp0sg8MnlEng+BmB7Tcn6+pwHtTS
5ZBaR0ke3imTgCrYlk7EkrvsA5yoKYBDFtyELO0gSg8JWvZxm3JyGPcqaLwbQrwz
jc8OknLTMWJkWoJlTzltkRUMS0pl50XhCdHaXvflt/6t/NrOLLdzW1DfZKN/Jbwa
vOF0LICImuv8AnzL2bgjG7tFOxbNRppb3CN+iCb8KkuAhgy749mr0yKS9kqaqsa5
eS2Yv6A7TTP67EV/tPhFWmGkhMXVsGRg22jnyzcLFA1zaKlWpj6NTZVGxo1vK/1w
mZF3m84k53uwlKokj4TDAGqyBg8nZ+V8dYJXip/aED6AV6h3g8zMEl/muSh9kfMF
BphVCp13rNREp6UqyXX7kGQ1tJ4QjeuRmeKWtIOowBmmMtjPEPT4ZDuAPirXZVmh
6EtDODE8S8XkIAxrIOOP5iq0oMvqlpaIRG4TzEgXOw6gueT/DYCSA4Y9hGS4vS3N
3R9jeo5pcL/XyymrIkEjDPIuDLPBxMUvBv5hSVaxZz5KeQ2z4CsmIERBZ/BhiO4W
XJTvR6HecFrfPNEHzvV/0ntRGzLQ6RVvM58QeyuctK7kX9prXo7UQ+joPR+6l4AS
bc8vR4Eaki5KjsQyRpULSlZO4uOdHoo/WD7PcpiT66IPF1sd8d54i0RP6XUJWNgV
RO6iV+sqRKD1B75lPYsJ2TBNFbN+5/8FhM45kILx+7PyeQrtMAJGKjyXO03fvtoU
7SiDa9P5shAWdqUv0inuhpQcN187Foz6WWhloVYkinLZcDUcol9JzSRgLMtWRlyZ
nL30vtcpLNeTwgW8tNH3yqc7jKH9LIKERTo5vSk0UlSgT7Awp2nNJxvf4u2NczoT
tBHpTlGV5LtwR006BXWnzE1/Pyxq63erkNtWdYJIHlHGzk4K20aIxtPTGxzHnj73
LqDlHLk6J6U+82NRAoRo5tqgoyFWXG5FPSxLvavlRQJoKd485psP90iQIyZb7rG+
MVUSG9V1O2TB/wAzoNRsnGq2G+aUyOs0s7Y/MWBf+SFjwnE5hmeHPnM9jUVIWe9X
qHimeJlIdROR6MXcz9+93TEkVE8bQbXtEEI+riG1nAlBRx7U22UG/T7EyrQOD7Xu
urLf9IpTjMq5hKIw9KpsEFU2l/wdlZtD8CueGwfAPuXLLIa+6dRWnpUtJ3MDW0X0
3SdJBWHTtBV9wjJ4uHUL7P3v46ae6lyXNtEwNtME7evvuEdzFtQQu7qMFsyIbpH0
KhlHdIgZwROa+kDE1TGh0FysW1N4ehDCoEAZdrEfTz6qJQUCm+SvTihT+BU8qgx8
QmsHWdj/5wOyynNCCHkiSQ==
`protect END_PROTECTED
