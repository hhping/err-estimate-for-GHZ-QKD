`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KH2ykjXZzrOfGO/qpG4ZmbSvoo5Rl+yEtbCACOunQKuX+0lHkhO8/kuk/tty7ruI
FEIoM4aZMZkM1XFNuCB57trPYegYRRDML8Fo8YahaHmDVypBoWhHc+QiCEsWNOSq
ThyN2sD4bwuHESLvCrX79vzRfhbhPVkMYIzDCrB4zsSjE0treIC/HU3CyWL2IjWf
jAkwKA28hVuToKJFWJFDTReREDeKvquF7yIUCbNPeuCZ+5rhl5fUeEZZaxZmtGVU
vaLQpznSZEGOfj4vIo5TbJE+rOyhGgmtLPVBtp4fDSOjGwRwBl8LOD1NCFvvvi/y
VUGbJgtWTCDcwxX3g40/0HvIuWJxixt7+aUJIC0JBGsYlgZ2QQvtHARX2XWnpCAQ
vxZ+QDfWNynxEDVv2HbgeJZWEeiFWlZ4OOfOqTzUXtXSTPhVEuCH6OKF8cZ3dG+q
IWLaECB4EDll2ndQROa+wV52IEibbN7d9x4MmJ3Ks4di/I6ZciMj7o1812MNVz0l
`protect END_PROTECTED
