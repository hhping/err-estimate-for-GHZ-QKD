`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PlQhpuGmzZbA/MatRH1v72uHFhfKn9LYT0ZlquWwlmYtFqDUDnrNQPFrMuAYTsh
qvByb6+fb3wPR96kh5cK+SKhMJxzgjeNAJOwMyNny/Hr3itLUqI8U2g8/xqsgMIn
DMRbeexasqDUHO/64P49L0jWzujhbDsjZk566EbhAHi2SBray7s1AqtjtaMnR17Z
aM6T0tdJDvFoPe5sp4EOe3Y7kz787dO0xIbu7jiAhn1opVEdmkmp80Axiu9BkFb/
mi++5W26EvAYeAK6bZ/VpwaodRuW09iFuktKVs+HziC8+wFeS1dcJBwl4AvEZ1+c
6oywUMNK0DV0GXaIExDH7u70FZsNzdET0TIDFv/EBwMcaSKwaGG9I3+G6ZzIA/fm
5w3HWmImBStjqT988aPecTGMOFCXpji+IXO3SpNlKXlMPBJMEPP33VmEWZjoZGQj
Z1kWnWODdIHrrmQoMXb405anAFsp4WwdSbs9VCBEx8fyuJ7WoobACBT91jNiUd2Y
xGu3A8Wcq/Um6S0UOUwcfowtwjlibQDcrWG6RdJYvHIOyaVWCmOuI4fRSffH1Yow
1vyzepiIzgob2ekIt2E9NaI8+OqWE936P4bkkV7WtGQb9U4UpuL0O9xCDImP4Drx
yAMuJLtmNfFr3fhPCm79AGS1yRLdmg6E8PkF3PTvHBHAl7BF0ghwB/W//z69+ROI
kzSzX3KFj/JLRMxqDTCUEoKKFtOkqPKeEVkUDY24TwzXwlgU99ba/6CA2boWWyIy
/VoKBfNJ6jI52JOsGWR67R066PHwQSHtACDJou8WH87bdOoa6mbKnkYZUM8C/T0d
jJGf3Z14QRiriADCDqArbTlre8b/eo+1EjgkVggmLWTxTZALRJdgVzqn9OEgoIbK
bzkLgmUffWV/JZX/1e38tY7doMlzbxdobva8gGuVM6tc/W5EHsskRuQfszzlKfso
imvODmhDJx662q+Ey2eVtrvJsk+he+m4ecSc1GdjnLzDj2YahUOCmBAZsVsK30Qf
WyWjYXEHfDPbl3yqNfIoMSej+pX10yBpFwR8Yfrlc6N+nGjSMs+JQgXaBvahAhm0
ieA391ha296frVzWMCQzLForw/n7zsjZ+55adaoc1ZRdpWwhdez9wq1CGhqpg7LI
WArZkAMVhtCtHp8WNUnAwbEJ0RO/9aFcwGSla1Y/PKk=
`protect END_PROTECTED
