`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvOx48EK0avKTCe0zUaHmgMo/lfPJIiqbP4YMZDD+JqUjZ7mXkFZn4eWWVvIFq13
DiT6QqQhTh3lpfhX/hP3zZCHATXPYWl/G5rDmomNO0J+O2jfoN8H0Uyd/9k9+0As
XIHBjK3m22rkdCexyhcS7yzrUnrn+n/mSkU3uuyR8iz6bRtVZr/qsuDMxu9Qrw89
L3f9uC8sEznrM2/F+SRFPDghs/BjYE3iKm9pAryhu55IChss6nPQbMAJVJ4WY1ZX
gQD2Tv4IaGRBUl6ePonVszCyLc1whoWNb06ejZL7ZH/b5Ayz0ri8tF0IA3U66fy0
YtKqd9OHeL2C/opmG+h/2kazNGnfOU1UeU+pJWj/arl3pLa/xSJVDXUiIAIFlIdJ
EoySaaAIeH6b5shk7kdFFIBZrIz87OXIp10MQbHn0LJY2sTd2ucAkWw4NqU5uq8S
L6b6H4PiAFVy2QHnRsgkq6AnVXavf6Y9pwoA6LpPkPXiI8frJKM3M6424KE6mz08
e0avUjqxEo9z3RSm7fH5HX6YlGad6UfWAPdphI8wpi93btiT4IfVkCYj7ywLBcNc
iUhN8L+kh4ejwOQm7CIap6D2jRlvL/XYxiS4q6jwqYgT5jvPaWYLcuuBEXMmRZ88
oTdNHptMANviGJCVGtO+OO5Fcn0iomjeYlfsUHgyZ0xvSbG0QQcIDg45GBnXYjaA
DaD4XxP1NriSj4qKzSNRBfzfRJcUaXTdk34TzFRueirL4DPdtS5jfZNxMd+30EoA
l+rPHw84IGpK+dTMVnobp2VwzqEqd8D4qSI4R15p2eWsVEc0R2BxrTj/kP1mUKYn
FwTMOPwFPzfTUahP0wqEHZsoi+5cN1SKHEYu3q3+edivyGZObwfVvddl5d0idrfU
c+fAlSMfQSE9qV/pDw2nmcchp6KAVwQOUl3nMRFHzKleKR8uPqk61s05ba7JhnkR
yvYUllRMqyp/jENWqy3WouADGP5V64IzdV8GKS+/ioJRlurHf4kAeomyt+d7s7cn
JIX9Pj7k01BqmmaDAJzUhX5t1O6+WgRvujvCt/rMt32RL9nfoM3PVyOsF4uLdDzl
OntjC0NS+7IyctoWVg5HhIOuXvmVDI0pKfcoJl3oOho=
`protect END_PROTECTED
