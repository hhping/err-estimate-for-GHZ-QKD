`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDolg1ziaigwlOFjbyYPRsmk0os6n5V5TW2cEM/i9NI6bpgyfoyQwzVoQEcZqcIu
Wk8pG0PKHuj05NU79ZyqkycSLFnMrn0EsZ9KKEBEY2jwNlnP7MJS2uFbOHn0/Vge
eloRJfOgIweOAUxT5Pp3byQLn0lAhMQjqcyVejbvkbdobX5faracRydr6mEuXx+E
a+YtuciMxwW8bi+ovG41wTyguFcissDl3+XGHqQT3bOoMgJ+mSdpDKXxsaYd/dI1
03bqM1X/eL0Bo2zlRbVuokuzADmO3w4UwlHh3oj3ljgkRSVfDyT9gc7usjIc8HUQ
2EBvFq/uy7Uh5FI+AsDGFgCHFdpo0oOBlvTsQDx4vngrekzAMlmTR3525QEx7ORH
IV8BESHABZ+oXczUsHsCPcxRztVJOJihmg8k/xs2G0djUtaZyNRRZI+cQB9TiQMB
Ji6bWTYiTzUxQrxJQ5HShW/Y0nNBs1vI2LaKJuQYnvzY4KiiY4cx7Vh3SU/4vBJN
oAC1rnLLG9N8Y0dJ0knzWXV8dXqc4+FGDCzBmhvKsFzmlq49Hx1CR4ce9gCARukO
eWmX638qgihsiOMrYMp9QYK2HCDUYLuzzrAmQpHKZkx7zRUAhZsMSzvaB5eL68Hh
KHtNcbyR/7W9GjClqUmWBHLqMDwqll2BABz7jMGS0luXYinjTcz1pkOOH5vul0tU
gLeb7Cgg5w5FNkMGGXwMr4R5q+4yFitfyR+tVy+0VWvf3+h1hMFbuyU8QeQu1PIR
S7q2DcmhMVOZi+CBylou2Nsl0TiFKJ1lVWTn5JHhBNzWYa/grnn0RebIzOTfpE1t
0RbBQESrMjSy/06fUyfcr2taWWDZyqBW+Ml+egBkQf05Fs9CMjHWmlm7qqbFx9yH
rIYdpmUonuXUAPXqCgrI1v/Jnv8pWsJjxUN9TuNlp0Kg9JbHjEdS65EJZK8tA5iA
rNSjEvslj1UrMbtL1b05tGwNC/WeX04LFao0oUtaFGyCfvLmdv2j5/9rhMGQTeU+
ZrtbgqpZ51oopENBwjCUnQOhkR35KxifrVgLfHXQRz7iVQGd4TLbwkTBwBIiQYpg
wOQhfMTB414FafIdGhfno5tfe4U1D/GZ3Rf+EoUxWW5DGW+ZAN38RN2nwjCrXiC6
YqxRUXcT/uMgJ3b5awmZL+7flVkcVYgkfgpJj+rUEEuVEQpRLeayNhz8UoHV6ANf
l2J9LZgS9sC+yN8DghiEExwxtXNKEUtFRwrCYa6zcyeIiLGycd8RUwv0+44UxlCI
sEflTydfUHpXqlxFMtOZqktOx8/Fx4Wff+YHj2adisUGAn6hdg06tqSn024NXmX9
8VsDLR1HzAKbJs1BBAtybZtl7LyEttKRL/VmzVizrHChWU4HgMfGpdOdKPaHKakJ
3LODyKRgiQqHE7cyrPS1ZfI1fNiz7ajhdp98AZdU5AbxVtANKBHxo9ciJR2CuvLR
VfyCR3eGdfKwT7qHAIuwPsblJ7/XeFOxrqYWtBPFZFWqQo/i5qEHOamieGuVGNDA
ZzXSFwXw03Zc4V8NgV9BR9qVvgcYrE9fOKhTgNP2jzj3P4hnEj79hRsnBKr3uxFl
Q300vaYDvOPhL1gQfPCbA+UO1X1GDSMiS1hqUBhpweY8sPiIr+4TIYDQdykCsUDZ
hLqc4qPdCNkgp2LhS7kXAedLmA2D1+UDHgCYItT6vfAcffGm5udVb51iHqUXJ9jw
aKPRNMXjdKXIUWO4bmCnvOXHHlk5qzacWIS2VganABxTI4pAlQ8+8i/2yZQUiFJH
rtagfYc4j7hBZnQ6HMMgCU6gSpJ3EReRuSTH1C8vjRHfwvacp7TmeBEM3VM7pneB
UbIAQRxWpio16OB8C0qnSZ10YbdaR382/hq4CP/JR/QybzBvnUuttM39M72lo82B
rkAwtfd7/hCFVK+CdWVS8WJyEWUGJt14HPvnr4b2ofDdxNyLckTKeu8rs644VEKe
5OrlSOKRwM30Fe+tKGTaMxsmywM15a1tkRzk/st2WJxLRvfyHQdiEYwjBaksk0AS
3Z76VrOy4VZfOEtD6Zn9ySK+8OfQT1evlo96HdEFYwAA2VcxBgvvcB3qNvftDEuq
5xW0XQW45qRIF8YY3K/A4nvVlb9KJkNtZccOVZ2G9NG7xZRyaDz49OC6j1sVSBUq
3H5mQuyC64YUylw7zyc5kTwXtvNXA8qdavhQjzZhrt3OmRXuegbABYJeWgHL+Ghb
NWfm3kwW58LvJMpbOqSH2ofS6rfitafB75yAMjSq1n/q/DgWgjEhtwhUFmeVGB9e
4xh+y3IC7cibzF+XVCPwJTOFiMn2mFMEhclKGy9ZxwevfoIdiaCI3GBIdz/fsL2K
E8hMzgv2elKl31WSaOAvzBXJKDjXk07RLbHMvaoF+vIqx7n5GoNUGLNUzpw4BvJb
kFvkDqq+pl5+F/Bpf6Ea1Omj9hEX5mstTuOAkTK6exdVTQUyDhFcEDeRE90TGH5J
tYrUeUYE6PDfrAS7+QnxihHKNMLH8Su7RGR/7SSaowpIhRV66wFpkbogsAUF/Rg1
fzwCM3M8RTSa1yRh2ZgKbBns/kXiycxMs+d4l3LWWczMlfVuO8AgeD9YEeLmqhOV
Zw/u80lUP7B23lf19zsAwFVUoxZ2LEwYO3Etn+ICUeFdMvkYpZYbWf0vpOZiHM3t
xjl3ILoFdDGjhij2qhJBaG9QC0CCnJyun3KGXz9ZIqraYLmcvjldRqpuK4EUeDQU
V661zAJPSNFFMHOCmsWMCbNHkWygQQ5Xqx170k+1TUavsYBAghLTAzDl/k9wi0Xy
CeEddKC/lSRDIdx7rETn6jynTHK9mJGGagJhTEOiBz2XZY54eiDLjxTExHuyUfBI
0RpyjaWJ/lYiHOn5I8UmawQanVyCbGc7eH1Yi25KNEL5A8A406AojoE0E4FXySBq
fwXKu4XzgrlBm1y2cg+iTBMRaMqjZtfQ8hfnchhXQVIbKKYnia/6ZecjKDpjX2uL
KBHMVOaa+OMZauiO7zHdiNdf4WiOHS8GQPq8ooLIvjj/J21I/weZwUuCtvi0pwj3
hBXIvydiz2XAnpqWkSspGumycjAG3/5v4vexXl0W7FZKzD4RbScdpvqUJ0lV9smx
hFRIT2U6RhBSe/JXvW+hUavEkbCcwn+J7FdV01sC1VIW7Xt4e8xbrcy2vNZ7cAK4
vdVgHB6B5afKWaH+L0SPPAM3EOGFyjL5Yc512CVuIImLZeJalwQaIrsW96fs5hVl
vOwXjbhCCXKPXXSRJ44hv2ZU+C1QkOBlMJOrpIbVBxx916RrHbrkEWrhVo/xKGJX
ZK3LNLcNm/9mV5TU/KyL3D8smVaLgX8GNkc6NSE13p0IGhK03O2125A5KLwVkJ3l
HLijwnLK66xZVK/YAReXPJbJD+Ylvy0OS6UGIujMPsLl1S0kwBw1sKYO9GBMTDIL
8+9vGle4ux9o8qw+MGCXhhaaeNinkURObcEDi6RdqdmrM0r35DCpcUkjzK2qb2ax
VvtqESSoDu1NrpuXgz1IjN+s0uKvabZCHCzmILXzTMCHpaul60JZy9xzffssw6zv
0cRjTC55IX8ZzGFXlziStIRCiT+ZodZzsh4eMbEoN8YVzLf/ZDLnzWpSI8oP1yHw
nrfS+iu7ruHO0j0wkbsHc9NSbk1neD8YrAVKU7FR1x9Em2FyIY+I0ev27NsR9PAM
OV4xlwti7rCyBVnQF47r6MU7DA+GRG0JR104PX+WUXnrDsydPxLUUWTu0ft+QW9P
A4mn1sSMKYPm/u8CZftWzhNXccNhYLvxRv3fsTLAwJZ9TkOHGZ2apWnU/tmVcglg
7VDbktPmXD6WLurFWoNMH8EgbtZjElWDJ7XKGTqsx9xY934SUeP5sujVA3mLXxzP
4wIagRgRbDZ1EVcuc1GV4jeZVnCme7SM+fEuXxoOUslz5T8Y7JvBfvipdFXB1c++
XZizRRyDrS0QOuB+YrirvTdme5NG02HcCwgRf6GcjpPkLFzzqHDrz5KKqEAVcvWI
w+HZHnaGVVhQ9dGZ0f35ZedxxRKNOk6ax8PgUZFJf1WGW5FrkXSv+9SZ3JHEtSgp
Wbq397v0dVAQ/+gQGzeFBI95BoFpSembggqibTAb5Od9eQ3dcpxXP84X4gU2JLqM
W7xL95QB/VtbvEPAmYw+O2LDwVvS1CwXy0DrQ6URlXR6fXmyECkR4Kl3XM2maIrg
Cu2q4uTUrnF6ACzuCQQFuCKImcBHv5JleKI032h6wQ+I48hKs9MOngodO7dthSrD
a0OSiUBChmImYMpO9LnzHXhNv4Fm4sQ2BUHhFOadAHaegaCaFxTHZGWa9xG2AW5o
l1lB08lsvBGoR48RNkcV8c5cYgP/Bu95gEuh2EEmxyO+d0wvmzfWcaD91Q5zMQ55
p5qsJcVRM0qoNwcluTmrlQSWo+t00vaHt3xGqV7Unq8Ah5aFu4Hs9E52tiVwopwV
KViQC2qoCA6tvchHEKGjARGBMaPmpJbnV0CFF6PAVbPdoosd7Qoiau9q7wvb24Mq
ZarlzdQpnMrt2+K1Nv0320dqKkwh+mnDTz1AG5+U4FR97700rQzi3D3C8fwKz97a
/VhROMLJW9+zCtvbUoUCqxbFYggXckWkf/smRVuxvvocPQXBGB8Se8ZyfMZRMqaD
0um+z26X4mW2wBmFzvweCy4EL6Vc24UKB6W9JNg2pQzlgDVNZcgC+irMwbqSoXTj
zxcdN3I/OKicHKawrhITdJWzHw9DClDHtccvpBT7v3QvBYZuXvlOezty+sGTLorC
ahM7jIRcrvMO22t/8/tYFkWPSPwXpnGBLoae7UBzHBdrTBbf3jKfV0+cDekkeYvX
wTxfKjd5uInyR0V93nhg5OpMyVuCr5S95dQUKKwQcoA8IQmBl5EicCyyj8qhBdKI
nsYnbsxNkwk/mlmjxMZ9E0TQWcBDvqLWXIcoEnMOuelRUGDjs0qRi6H3NwS72kTL
91zZV23GCkrmQcXqN7QcbMm1wdKQaOQwiQ2QWBNTX55EL9hk5EWhqM2zxEFYLb6y
Wlt9TClcOoRvxDeBkK5TWG5067yTE4b3iVLvlRhnm1Ewe1AspcZA8pBKKLNvJWxA
T81NoBCxQKwL3w+gbO3Yxz/tdPVH+imWDSfabyRv1xRmvCcXhxkMnBgcxwKbIjFL
Mqme8p0MIitD9JxfKltajQDrFx/bSv1TBJwBunF5+tGh0c6T0LxpZJyN5BY+tCq6
7c+VGRGtaZj/g62UQs3tuEq3F8jTdgZ6Q5Ilx05KIUCVEui6K5YPh4cz+tyDomGC
GkX0ImLtOaCFdanbAI8hgv5ezX8gpbIafj9Qkol3zMi3wetJxqdeaH9myTLX7RXV
VOKAcjqeRo3iBd6a/KV8xVZbP0iU2J59hwGAHRFH6atfZOCrrgIfA0PcdRf8Zj2H
Y3yr42iKPT+Any/CoaoqTNwxs5/mKXk7QdSWO4xeO6de3hV4sFEXwXJqhr0rTTTy
qShuIdvbfPyShSJ4GTBwwAzoZ5b5TEfzIDtqWtxTTiFus0iHP3T83wSGfFChWuSZ
1hX9DOwmil1YQyJAZnYjZKc6mD0c2Qg3tbLZwLE81Fpc5+KChEiBf9C21GH/aJvh
26FsppZ23Lu3vqOB0hwom8nn8hsmiw6pbRD/uSlST7/7x3gtHbtRD5XQsogJbGD9
2Vh8YQ0INMI5RSXWZW1So69m693fr3beIorzZQfzlu5meoWid7jP2BxqzduLDR37
so3ABEOPcviFyLu7KW4DiUWEjuuNP2+fbMGdlYFluAUdjYcBbeb5rodqyYYSsMKj
Ir8dSkULWPYMGxtQ3au9yEheVkek0sjqaJc2OqyYeXLbO5ffMnDmqKJfoU+NP+WV
TcFz2oRcZCPtIgPd3GO5GmLMvwoIoalH6zkPWZ22b4OMQql85n6Y9TYqGiTzr11X
xFRUG4QfqNAwIJoi6OgCJPJo8Qub9uvIl0bAvOWw7JcsOAHWs/aQzy4axun89AdH
INuET7iVKRU4siJnBmp7lNwEIsOzS/GbcpzofWwtQl5hRFEuScALL/YSV/cGH9QL
IzFXfGT0PAyRCUcULRGNbFK1NOZalfral0vYPi1d3GuiCZyA+mTQswArIcuPZCC0
/Yz3ziKxNBjRqtFUEWJrlytdoaQrj6QTrtCvlIUOp7vzrL2en31nVCFq6VS33geA
92gLKrm2NQKfNXfhhW97g4wBm7V1clOGcqzQokB4GH8SYk8wWqw+Xdrg6FrT6pis
Z66zF76rwdhHvhbh7hOM39TSdp0ol4VIhkdRHpRSoXpub4gpKKAklS9hAy0AJLxx
4BYLHQCWQ4D6kEQG8VCJSPoERMxZhnsdelkO3BJ08koYsOywqNi+qoppBloGUeMG
mmlzAQv3PwU3GFWOQ/Cm2CDUS+S7PGYCrr0PNeKTmGe9oonooHsjtTpb9OalCpVh
g+r1Hy+hRnl6Q8M3J9hToyC68ErKcDfniKU2sAxkA4AGMf68bXzVBx5ms4fdvbnn
adTqTrJbJkFbkhFR6q2XbMLk77teNF1pLCo16VTyqcRudz/aUMV3gAcONqOWAvtM
ocyJ21uD+e8ho9L3GI5Y53LH4/x5qN+pPp1GLwu1g2/z57YZjbwOxEPHXLjClULt
eDxDAFEGO3blh/o0PJTQFhD+fsd23Ai2bkOMdt2D/kThzn2TD5bna88myETQIuum
ZLE8zmsEPSIhSea76+y6taapVa3oG6kfujbCrgYqiKcflQh3XKNcF8lmAvysgiRQ
R9soM7Tmxslt6UE4sElimFybLg6blgtA4nBIrS1vD4xclAjltKn3O/NoW4Z3b6sv
x7x1tpge45yU336g9O5rsJ5NKvVPEEBwiERqULkPKrF2Fm+xcOgpY88w/3mPf6j5
p3AdZSBgzvSqSrdQqtEwDQN3i85dr4TEPTZnQgMEKJZlOOAkiwdZapNVUBOMO8MZ
8wvnzw6ItZetCLMxA0HdayCVQvpW+nh90OGCUrRe6IBAgPmB4SPTJhnVYF/ASxx7
cOgaP6GMu67DDHlEByYjwYL/ZiOlBk6gQ7c8aPp3m2FLXdWUI/+EX//7Y9jTd4RD
yipdztRw9a+dQKoxp7t13p+5hFAe1NSMnIdAYPMw+srzMmTfAMZvvEVwnLsIlgg7
7TEoJs1K4tAGd8shMQYcdIZzT+180LiicuGtDZNSMxsM5iIGj3EWkRzrfTAPlE4v
TvFAG3hU0p6B/66nhfvLVGPv43US3Vl5DRimq9ihdOAeSWsw2ua/zs7E5FWVAlMY
gnOe5Kn55EYAynKCor9gv6UqKsSPZf406ngmuO1mP3HfUUYAOTHNc1SIJ4t5siJE
Pu7i9whAzvcIDx6lK2NYramYa6Eeh3mZW7Yns4YgVp8o/kCmBos4ufkA45Kr4bjW
AZxX/x14sLoF0EYJeJzSrMyhHubWFLMVeWovYzhU73Tc+QLx1gQD45Wr3vPjKy9s
IHtU3oiIaTFIR4SaxqB8Bu0EJsqiD9uR5NFe/KgPyqdFRrMLD96ciwhCMwRGFGZr
xodCoLbZ2WL2seK46iPnlRpPhFelH/BlNAooe7hfAaDKumnnFToDMDwufTPTjBlV
QPLMxhz5NB9q3Z+w7z4k3qeW6vKAUmzLBpl6YmxNm2JmXKn2j27ynwB4ctpkLA9a
l3R2wdXCB9V+6UklB8TBp2/P/D4Y7kx7Plbt+8qZ5EvL0liFONbALbEjBTm5tsMX
WrDHwnaBPDCbANFWveKhd65oOzvSWTo1/MgGrVnE4N0SI0ryJqQZdpvZjh1vVRhe
uQyseOJNVZneOIe2CWU+kvw93FfazRShF9ZioCu+2FWE3f+PP5FGZQSorhvA3qJJ
SjA08Xn5L+3B4B7siXvzswa0cYrNLHscs1st/JCXF7sXLRHONUaBKwnycxjwL+9x
NXe2VhlgotAqGngijs6cYFhOpck7N3EKCiYR/BdH2xXECtAUVfbKX8sLiRjS+kpI
pTtUQ0VmBn2+zH6w5pZjzDNd2y1sEKIvKmPaOkHVTdDSd0u7ZYJD1rQinc9FF76J
HEnp/dfo/2P8Go8zsJHp0tn/oHw3TLODXcqP4sPfx+DvvfTBrWyQbz6U6Gn/nxL8
TDLqPEHvL4W22vy+x5cWnUFSWrIwye51fbJTAuPBv3FkG2sGThyuLGkeZM3B5H5e
bP+fTb0/xW50ksEik7yIs4LIUELl1lVjvs7FWzE+FFsvd59YFuzy6chGQMr6ZUpC
RV6lcY/0FGXC3f1dk4FciHiZDqqqnbtgYgBZIIJtsfdUVJZ0mQrDav1PwRitk+6I
yRcFKws7pi/tMAYDGOIRO6dhfqNS2muI0gbMYEKkECx3iLK2GL+YgrSbNv4mXJzN
/k5xlaSsr3ZwwyvXeXCWArdICd9oPmxAyjgdTQyag2HOoqCYID8Of9SJBu/VKgi5
G7A6Ql5/Tzf7lert9sG6RqMMC+/ca6Se+tm240oiJvJYKDArrXIwwoJSQVsRDlMi
Uybu7i4arNTmt1UqJtgAoa7LXxEC9KYfzLJ/VXi50N4YfdWUo7b+SwzatTUmZLBs
cMf5258jEHVN6qFl07K2IHR6Ea4l8/18wPVghGlCLfkVqzDuA6IplZjtjmNpCDu/
A6EviUlqSPMAvU2E0jyF7jbgSAz/lelp7O5ueQbh1SS70+c7/ThjuuBL3fRD+nDi
/RWae+9Y8i7YsGT38vWKSI51bHrNwer3Q0LpyQCOFJjb7Uld6gLDCDvF6ebTj9hY
dnmRpHPXQc9VsWy6fpr5QaGpnmM5bGsmZb0pSs9e8AMoPJSUgdJEyLHQvLRRPIuE
8JO/7MvGTjWOB667CUsqa1EG2S5DFeqRHdjildV4Jdaun7ZVUC439VNRqyhcr2Fn
fZvdgH0GKvngEblGRSHVIT6hTcvK41AEOv5wTH3tpF4HoewZxH4UoomSsyfCSSMn
G8Z06BrO0tmifBw79BYDfXXnc1ntYGympK9iHKSFeYrPGhY8VdF+RO9zd0v0OIRW
9h2cFtg53h5dEpEb0xN77wkDP1NBTkP8TxLsxreR3UEFNwOsxhKFSyXw8C92jWFa
FU70ZSJyhdcZ8EZek4GxCwCv+sTKwJRaOEYWHNBNjOcUZMMVf30i4WxtUIJEOtZo
nc4iOZhNv0KjHocubISmJW22HSlSuhblXaibzGE8Q0KLGRQLVg97jgRssioIcNve
Uf/D0zNQpz78sjn8E5Kts881YmXx2rGzeKTUDqrrUcW546X9adS6njv0rn3IJOsX
yjyFsNxe0qkNbwauaYf9mr+cCABSfwoBc2Vi5f7REbSfOjd23FlL2t0piNLNFpX+
g0hodo8w4LLk/OYs74H4GO7ajOuqihfHsbTn8BVgC/Uv0OzWV0J8OJCi1eucMWeH
ZJTCyP7Y2928OYWGT2tQ/O03HVdyL9XyQKIP7wF0pWmy/uJj10JnZ1EPK87ZozF8
9JIjJJFLGFbW/+aXrQyk+U63yM+vE/VmgvtKganP4h9jClMLxGYYu21ImDgdlW2t
7H909Oj2tSQTKIKTat/zQUoCtLRs1QxxX6Jiof21j/nTExLCY9q9siIRfBv6j3Ji
kzIopQgyKmyc+dP6VNJfesLiuejemvohbcQ7/pabLtjR4cPRHxIdjo2bzjwzDcwt
WWZsUKOd3dXdnEvJPZoki4fMpbBfbSJ2D7YfgDBhwwGY32RIq6cgupST/IbD+gPN
jNfSnYxEOCh72GVBUAmM+nstbspsTRzq/435NLCfOTqf7wOGiJ2jLynd+0I5Cvfb
lI6bTNncej65baAnZr/kEiadtSe4tauoLutVKNMnjhyZKlVs3fYH3+XLAsHOPlfu
SJhpKNpjechM+jEMX28qfmyKMpbVnXvrqv7ffC49YavVrtUmAZI0Eif6r5LCjqbd
fYdt0Juo6vmlN4TgYyWCq9J0Q6DEe9NuzzgBDqGbP8Mua5ErL3FN1WN8ZVto+4Gh
1IcUZ4bY1WkcX1biMUVdhQlUBbF+o469s9wXMGtu0bBpzw/j09uIy0RWvJ8B8oUh
+cxRGAWYH5pMjy3bPEvHEmehLx9xl6LOj//ZVcsVw+gKP9VAxahq6gf8cPuWIGDq
dkPBXzjKqysZOjf4TD/8m+iY9DQMcf0n1RZ8eIIYi+DQi2GYnyV+Uu3MVYwNn+po
dYc+F65gNGRBc26HFX1PSH6zWhvxCBZHCHJaEL2DwMwDwVKT/7ypT3bY9CTM7nA4
+h1i0TSrpbEWLeQjTKj3ILf6QaMwzWjduNhserlHFNq8yW7Dfw0ZZqTq5/AeBHR2
2DkCoQiVlG6rTUKPFTkzK0lTXP4hjrnSGCKwDMOxWDuZSuJ02aSAaZ3PnhOs7eqc
AZl7f2WzKmamslaei9BE7DmECvxMYyvGYhL1k6flCO7zcOWvvGdq3YPZ2D7j7E1/
qo4YUB/qkL1YVbcU346JXbLVIBRXIwt3d+Tlq8t/gpvSHvvVvskqK0n/XULjbIud
3ZDlZu1PltX1TRgIDgZoMRDa1xYfVPfrGy8xj5E5UYvy+AFIRU6c8x6LWq9Jsoxy
yPBNzi5iOHlv2lIjG6wcmJI+LakVSd3MmyaLVL2UCNjb+36JfzzbkGbsSY5ph8My
91baAf/BZlD47D/AJmEk2iCallcsmkOcAUf2+yC29V5amkBH8kywIX1l8/PujBZp
pzdJi4gew33R6Ym6E7Ig6K7v5ni8IKlDsSPFKuw7yRXUcuWyvQCqACHsV1GREm96
mD6cF8U6yN2Rda1RQh1y7ckfrhg0poHhvX5jzelkeBXXAg5FWsZqDMQTzk3O9r8f
S3HefjT18yvCPnvfKTQcWKEqvx1nJDDi0whj6RupJa5BDlOM0Ov6riU18FaK7mFw
o+XpLMmcFe8cis+PMBwOpiA7Nf2SrwsEjV55s4WA6HWdQU7HVrLzADhr+QGiNWZZ
ebcPFLlDL9/YkVd627CdH9YrRVHOlFghuO85sqo1W1tQNRq/4yGiIP/jTX7sgG8n
vy8ndxN/a37PGZYy/zaGyiLeNlqH46mf6Zs3auVC4PYCTAFl1/TDAxOitwFt1eCV
6lvwhr2cHFQfMwbRLykguiaGVyis+gPfggLWJAsdvSkMd26NVUAsx1JL0A4JI/em
qnoJNBRUqfMun2W+MmrFkAjmHnkm85BhqOzabFvoAduYNdM/7D3UjAxcWxvaiQce
c/+N0gxpVPZ2UTTvjtZASBKTg1eyb0hm3r9l3HGAKJX6JtyDdo52vuXkzBunMAVC
xgfRqIa2U0WvOUO0DnCKsSFS6DaTxbVj7dEIR/eQkUZAKl3WpcT041brpFvTJKJC
ZJH+cTO1DNH96sW6uPAwxHTkGqp7PqVmqugMNgFeM0CT0TBF4vspUcsUEaF0JFuy
14Rb9cLYJLAOjZeVqAqYIDP5qJBaZ71zV6uFpi01o7ov/Fo9E3JC1xi8EzFOPmnA
TtJcFQ3asjf7jkJEC2QhtZjsyRy5NTsUxh9uFoYhveXvLnQoEeVejHJwt/rbSkeb
XUti0THyPuCbn5oRsTGt6oKSGbYXlNaiYXUZO73uK0Nnsyy6YPVp+fKUqs+IY5lu
cX9A2r9TpLgNbAr5FBpZSyacl3eqIL2sjJUJ4ag/uxYo/suWlEMPLd9c5lRqRO5h
r0v5aMRC0AJkNTh+cjUeGfEFCCrj+kR8mV47jXkczJcqUEYIlfI+sD3baI1SBJvM
U+8ExQYhkT/hTUnwmrrj9+rp6pGzFXe1SXzOTlPSnr8kCvVi7V/jSeg/RZfKON+5
2ckASEafN5oI4/xFtjZQtcEEZLzcWKYhYUWzaviXpnqOquRFsrH8lNHhn+3gTN4T
KMKuk/6RgMo3sfFUQMUyC8VXl0H0ZJBfVVeuEOrjD6zstipJ0iUb1twTxNRkTTzp
UIEHyQlwSOWzPuknOyd7YcpcV2WuqXpSz4jsOgoQMuuFDWqicI5IuB+nFSCWJ6sY
tc1ovuQo2clgO80CkkdRfPdVRqmp5WkJmv4bYPQCR6Alop53lzHati1WpAGWSe1C
g7v/wPHSuDiOTDRNcwTAxjTgG8834s2/N22CijwK8bnl2+I5InFpdk5vMscEtVrA
BRRiL8WuEnnt8qbGBmmy3JTmQZ36hrZP1Gs4JlZAxH0mFSfew+pEWyE5PD6zIam2
f7F/33RvnttkXC1yvcrXLXUwmwuep2lb3hlzhsrhaZHkP0dxplXmXxZs6fR1bGpX
aI69F5Bo/kRPYoSMNNKnpAhfR3G/c0cebYjf3sMvEbuu+bLjezkc5rl5OMl4fAHc
UPwNewIqzTDKd98fVcp6K1Eb5ehK3CmVpIgYoi6EcHhnjB/xnaae+j3bJsbW4AtR
tofxQwBdmfvYWZfVTd+fRCjEx6/zstcE5ZwlY0A7QMMUB+x5y9Ase2Eb/kNE6hX3
SYUJjlFvkqRnz1wqNRupxB8VjnaodiZ6lm6G724um74GrNGUFt93ztQnC872sWpl
UZpMpsClKR2dbmPgNDF5GZ4t0zHwAuiRpckfVpwCAJBNp0wUGpCtREr84+UhBmjv
fBbFHsKL5iK6e5WI8hSkmKWUGsl+TE7uD7teahP2V4g2VQ9wDtXbUKBszny4smpV
jzGuI6Yk/8WwLT5Zeha82Jgoq4m3BlF3vBrp5xaJoQ09BEscwSBtCN3rkhAkDvzx
oL2Js1zVV8G91/KZpeLSz3Jg0s1ZFT1+E+uDhSU0aMFb7pvsVxMRf1GalvfPfWsR
tcQvhFincM+1dy9uLlOYLsx/qPrFNMOCFTxqS/UO1tR6mtFOxiZek8vr1i9dsH4P
AFhOROUaQfBqANGruJ2lyTVL4eIYefs++dxV8PlTKfeEbeot+oHRO3r05nFuctEV
agrvcgWeU6W2fQ7bP2qYlnSza9n8AqUMRmA9pazydrOo7oq5yfvFfThSSvsx0s/t
9pFeo2UprxuQeCESUEn/k+pGR7yA3Ky0DplqwVXdo6FGCbbBfocK3p5yUevmhxiW
WRlSIhLPdTOfEuOoXqEg7w0s2dUQtsnz6bcQ2UGhzc63SZnc59poJEqObjxXc1wQ
pLOtl6lEdKJrRTZZM6AmF9935DdFQbmQFOvJgCrjpsiGq9J6ny6pOx8nebEyuCgY
pP91sqqBCwQrhYNkMlq4CDFxgzUDWHCundiiSxgdnDTXD14urDEyL9IJ4vAx185L
UAZTOTIZ9cCWKM+hc5KinhzB5/tOTstDIoLbFg8o2rBsRBQmZpz7BZVrdO2vWDWc
MJorsX6lTECQVzo5Ct5OyPWTj8g0AA5DsSX2821An5wVTjpR6bfoiVZiB5XTRbVG
oIfqZI4559WHEl6b9RH/u3sJPULne+hNF3Ho9E9G9EDUgySbLPRpzx0Le1P7AzT8
7yGwXlOBhc6FfY/2LiCSbwtSp4g280FTswYy6F61BBpJLSC1Xvuj4Y7tSC5dDFwd
S4NkhzvCmm/DM0H74ta426wZkDqwHwrDDcE1bSG23t7eWV+mGXtX1o5uoNIZW2kO
lfpv5o8Y8qySYxcm930xjGOSNpsZcifghKanMtz/WKFR7BZ7tQ45L5w5K01yucfe
oedwKGPv6Lw6zJFI7OHqThgz1gNK2ogybuni6vs+nrEb9fOSh6tBPts+0KCYrvZA
w3GLrTs1PQGRDjPCYgImgncccxbtnA3ZeYcHAySf+oTPpo8tF/jACplUnVromHnd
8ocrWSkDe0JbLBBspnhCIgF3e2U+z2wG1OPbJzxqjr2oTU4JKmlVcUKUF+5d4BZq
ARZemeKT0ATYYABq9c9MgCAUN4d/z4vEZhI9jOZvViQNsfKmzzQmQvd6oZIxFCR8
/AA9HwSLiDGQdOOkuv0mfrxSm5LMq7N7DBTwlzbfkvC60+BE0Yn5dd4fYEPbGX+7
h/hecHOi2ZjbMMuLQRQGZrESYjJC1U2iWmnOsbqcT305JVY7+VrtMOefVTFNxTWD
YWbarRxbESXXM5EdnELoQihoBo368SnhsbJD12YC6B1fId3uMPqrTsdVyJ7WXzI/
OgQxurnFy0afAgUNHGBceeyi+Ro5EcQ+0ZI8M8jso6A5kay2aoTosJVrFhZ54j+z
UCVYLA82CIe4V72/stgt+TKI4i8Xz0RX4uIFfNSJCnTezJ52Ry+lCu5JR4TKcTxy
zSsxTlmmmTiidtbf+4Wi5S4cYIjrgo77k0KLLtY48Z0nUNejST/gpB2pRluWQBD2
8us+AEQNK+D+WmU76ey4VuNnjhIuoz5Jv21YuUklS319Ez6jmLcX326N7CTxun0i
AsNoWAT0GnyhL1MHJ7KJu+L/jw23ix+CIpDupOlrbQVJKeFkVG2yddMj6Bgex1Dc
JVYf8+0B4y1id+nWEn+nt7oaoPssr1xK1Ff9oO2T9AATsVwPW7S47MvoPomJ6tDx
qwdw0KrfvjqA8mU2V36OizxKGa+rixY3Eno8pN+3Y0ITNMra2ZaLpzGEVMYyj3jf
2pmgZYcclnT/GsGaOJ02IuqxasH94zBO2XmWFnMWlD3BI0fU/+BPBkFQdYxewFuQ
U1zjoS+9MDD3NNKMn+v63A0LkIweCX1pfgLV0HrPxgF5HjWcVj/HX0QR4AmD7kHI
FrvpidbuArL5okp+ZDvHVdxN4lLIR6AcDBxuMllnBJC/9VaW+09kj+nBrRAwcrav
efq5jMPD4JgacPdf+cLdO896b9VKzlWvbVHY3ycwRvFXiGaWHZpXJtd68FE+eFZy
wTIOwQzHZPgN1Qd+gMna68XaXgnJVsCLMzX8qkWgrM2s29OZ657GEoi/RfDLjjL9
9LRqNfOmV1CU/F6HEiTrO7b3Jo17GmoPts2Q97rJ+6ouLACx/yj4tRAkC67gdx24
`protect END_PROTECTED
