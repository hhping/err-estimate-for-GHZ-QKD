`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fito0WNHFamKGbrTMDFdg9YQWMYlSRSe66VT6V6ptrEs/Y7S/WCcZYXORESc6tjX
WN4Qyg736niCcypvE7NPagqb5+S6JztOmUQ8/cZQdPuM779qCVHGB1mNIDOgh8tM
8AmbO/9eXgiuKkISS2Uxcgxf2fZlZMDsGE6HciNQe3DyEufnG8SysDP7Iliz0fZq
rJ45b+j3msIAyP4wD6SgvUzL9gmDtYzKi/PRn/p66fS2QN67uwIo7YsxTpM7+eZG
H0WOjkwEnO8jbhri/blGs/qOCc26INWCnIPZWyDwSCQ6cBnaO168PJLD3iUMp9DA
gTAbuiVRDaAF+OgxnoMYT1wVAfiaBW1k0dXES8cTUbT2KRmgxn7TMsaIbIJxjwLJ
HTT54JqOeNt0eUNnD/PtPm6UtY16PSsHvKcbaPD0X/drwWKJktZ9/nR6jTH469nT
CF03NKFmxT4WxpuNT5SQX8UAH7kgAantXj8cQbCNZKRniFIYoMSrUvXpc69PR0da
J4u4llNQzBrFUVQf0mVOmCW8LERIf64Hgj+rn+f+janNbvSYhfhECAkag74AY9Cf
yBiDcAwdpK6YDHVXydnDUZAI1AmI4QEzyFV1eZRm0Ts2deM+KwBQPOXIYwOs4mD+
Te6bAAP+hYC3kLNkFDOk3uMhiF6YK0Rda7Kdvr90l/0zx9P7D/0gkUIL6XIW4crK
6yXPfKWTO/9Ud1k7NHyossPpWi1NiAoZTJEgD2tnJYfQ+RE0o1J0eF3HtyYQfy2T
+wvB5PxWnSavZmZcWkBbpjYQO1uIwSh+yDsS00uIFR8Ph5653f5OeHE/7HuqNWWt
sm2g72N7XLjpTYJfDpDQXiscbwN9Uq7ToiaYMDBOizo3uiWM6Tl7JG3XPJbXxf22
xPhLOCz654ls6H5WQ42qZP8H7dd9AS2f3yb3bKHjJiH/71WWrDZjgPClr1jsVXyI
e9mj62RC9e/lSy6C34UwJKRq0mlvpR6nBHtRWO/wLY17uUU0D3uHyaddJKQPK0R4
e+nzqsjHYhUaz+IVvUwk0A0hgwdI+623wpPp6BS5yIkJ4T6i8BgsQMFP+Pc2SeNU
/VIboS2Y/IDy3MAqJ28cdFbCfaY9QYpjmSsBcJ6OrGaa1KOqbeuopH4TglNKUWuF
heIo6w8EKVxQupFCz1Mjs1Pla42H9Du710iAujQfp46xB1/Al+iGtXhn7CdGvCjr
nerK4UNZ2IeO7g/3YWirpOG9/toL+ALc63B4leESziPrGe2A7fyU2wWfy1yzqWIt
jFCHa9panIy908ocWSpO+MevT7Wzc+2X03jmNC4D3Bce7AMT8f06t3yMygT+7Icz
ptGxQUcOxVNafTLe53g8ih/tTry2ewPPY0nabvR7vw6/TIrUZIIg181jjDiIGtUk
X2IK7aqj9T3hG4TuUAPsjap5tmHInW9ESkBl/6yrFhRAH79R8asuT4F3iiOgCvxG
5j7XJ/686NpZKvtlX46tMl4GvFNs3vyxrZTIEzcRTNdER9SyvZVBeePMoASanbAv
PIXidB+rpgd3YLDPYhOyh/eIziNUdLIqKRipna+0nwS3f2zLlpy4zH1gBwLEPKPr
Kb6Ai0Iwud86/bZO/CnhMRGm2fztn9Js9ZwFvCnz8k85qFOwlz8dsqS/c7P0dCtH
tCoU1J9SkVQCouWYDL4CZSv8LDeX5oVbQ+OEc6fOw4vdHuM/MnyG7bjLv+dzWe8m
3YXN3YQWKUQeTEYwXsVqffywqfSutX3lk1gmwfL/47/h2xuT1H06ZXtN/ksVNuuF
1SIn0s4u4edU/Bl+m48ogyWuuUw34ZevPAtRepaQBEr58FVgKVvxPrtpF70ELQxq
wVCt+5/YoOTgKlUOYsMJb6BlKF0KrKmZsf+0XVVec3wyAAcUpdOegZB9S87f1zZ7
iUBQZuB3odRPAHrlObVVRhteQp48kHXHHpPKaDPECuRAgr9Xn2MF8uZspMXXeiOK
PHtiZ36oEoUjLXDPa3zox+q8UA5hK7GHG1TL1mDwzGQKQWxNCPgVeEIEdf1H+mC3
I/UgTgBVPc8feRzDieWl/nNkQh7odFhBawFr7WCq2aKJCcnfIE2AHPQIkprRb9KI
Y+vWOcQDsSns/qRUWsdmBbwA1V+jW07tXTyUs8fkE9Cs85Eh97ykIigim2tcAgxr
sjXoYx6uCFG74m+3Pn9YXyvljXoy1tqdM9beCUt0YeuEJJG+8mbQltYQwWA37enI
fyi6g/jmaj1Q83c3XHk1QELAUv075qefi4+5jeMcoCtfU9ooohqGS64SJAxhkJC8
it4w/XbaMq9DLM8udm7qUKicLg3UY7A1BRbIiKz7elmFwsVUfBhErRPn9wCd8EGQ
Dx6HZDhof3nK+SM5dhGeTm4vUmHEB5DhNvEeTyhPXJMv7xd2Xo59eVFm5W3x8ARQ
fgucS1SFRdLav6kJY9+LNnTfZFfE0vOqPE2ObWI3wBvs5g4FxyZWu3XEywe6xI2J
0IwQ74n13mzatZxIXg/+LiSfK+iMFai+uldEYJlANQ3Xwx0nDrnfHM2shNimMzE7
GvstNE8rmisqdF+3aEnh2xxwFqYzzaKmXCLgZ+kFxV7jixKL5G377yX5cX7PmNcz
XB4Pbi5mgSHCxVu4YF6S/W11teiir+LL23fFUQoMw6vK25/zqt1Uqs8ZVL5G74O+
WiZOLGEbgooOocwTfcV3WDZtuuGQN9d1Mu6RZ7KNJorL9SfdjnTq2Str4tvY4MPQ
jKrl/a2CRS3faL60uB8gVASFMfw+8Frn/Qpv0RpGsXOASMmuQfCd2ab6/g8X4Zy/
6gem5WBe25Ni0nVcjW1SAwJ1LbgX4nm4K0zoECbe1+3zkPLWuQSnOhbkFFa6iIiS
DVATwg5g4iiBY5uU8LiY2XE1fFkPUl9u3kNw8jwLmogbD36pDaP62+Ra9b+VOWJw
XyfrjZU2uiYZjJN+GK1q8EKLdhIayTbjrdcI5zerosLo2H3fNMGqqL+0bLB0xijj
3GEyBlzGL9F6/A0esMPzsUvNYGRbbuHAvpH5JUFQ/r68EgS0se/aolSQA0K5ibhe
nLKz0PsGo1fCHL/ytRRAM8xNkB0WBUONMrELgpZfVuVNBk3/6Xvx8+t5DtJfzPzl
NdtOL+NOXzz5ainMsqKNCajsso5yG7YvzngdIOM3WsA5FavZTKkQT/Sq29BEnyW4
H4L4RXXJ/7Cye7pa0xUe3m3btXMtBbNjIwAI74T9F3D4DnCY0lFy4AXvDSkKIkBb
7v1l10NHj8jgUhZ+LePGDBIiTA8DqMZRhYKO/+KxaLHJb9korSTNgq8X0yL5CVtp
EVKBdK+z5a7Bjz5AUBoF21sZoEQpfDQYwHOxfcao+Hf0WxyuBfMD29ozU4QTpocO
AwaGdjPEnQzyVKhEDYCkr1+mjMFotJWfLC+kk8TueyRJwzCY8IGq8Ycyqd+TRz3P
Mo5ZATsQSGqC1q4RzBPKQGOgEqEyyYrxrAo0MYmd3Ubamu8816iv/O/KU7f7OXIw
WssLq/aNiVyNi50PFGXIjVo+0R0/1qacl3I1FIMV8FJIN50R3dA33Hl9LPnc9n7T
5jTRCe1oXjkKirIP/pRuErwYSnfSRUWO/j4b16OYB0Rlm46HkqX1gXk/dxbHJgX8
nIZ5t9FXJZ2yx0hd3+wq7PdGInnGgUEWSuKvnWeDF7DhVOtIqrF4DHDBSCL4sIew
ARK0a7OWJHVH3SVEkpoWZ3fQxffZFQtyb/eYLCpRM4NmY+e9ZNhdQWgRxJu6s9pk
L9fGQGv1Vo1a65WaCPm12l49K/mBfCSUB1OQxSsg3/SfXh2/z1G+N9ZqsQJyr4xI
mPtjglEq/9ojNKo9aewnIrKl/bdT7+UFAtJYqc9eDdgfr8GuvEKmxwe5kNV5Ym6P
fmJ625s1aH9pwofihBhQiIQQstM7FYJe4TthVXsQTsY4jKO9z/IcRnNBifuLGPK1
8MbOnE2uf6HJsZDKZCruswhIiKXrPxpqv+KGgKfIg69z287oK4q9ZVvHcHlCd4fd
1mpSyf+CSIpbHHRl2oXBqA/iDHqI0h0f4fi+UPPclg5SIyfiVeFwmESooLo0TEEx
KqgE5FXSt4CWwFyQIG/PyBny5s8RqwJi19/b05v8Pjqksj4MdylIXyUAXTiuylsF
UAaX7dS4VWFxJqmEEB0OOEMEr0NmCGhqfo6vnoC+u3Y+jl5/5HzWk/rG0OUT4xId
mIruc1sVjhhwE/uMSNdR7Gq3vWwm1jHRZJG4RwJqa2PHymeeAMc7pUFwaySFrGF3
g6Hr348OSOPekcCgSljHsdiowMuuBgRGW9W+Hne+VuAf7tNHJd8rss7nfGCQ9LOp
Xo7rm+Ao3A/jQLnYkf0Xo6YY9o4gYPpNyY6lPWY0MSdVjBHfjg4VoUtVvX3fifuA
G/jqhYgZVGWj1Zk0gtyT3JVF/teRKDwdo6Smev/UoYz46z+GhgT4CKjeC390sxBm
YG7g4jK/snywIrXv1B+FkE34+xtFs8z0j0ilZ5trN4wqGN7tadC9mKhHQn1+eTYx
esHeF94SrOnu0Cq0G9KJf62sU4zpKsZUy8z0swe0QP1ewPugsJJnQfsw6Soxdz6O
6Er9hPPAHDCzlWT8iBnZeIgJW1UjeHN4RauH1bo7SOEhnkmOn4LCo5ANxJAHV5CD
OuuxUxD/y4bKYBbbdA1e38U2jiGDzI6PeFJkaw2zWjD7o5ndWw5uSGifO7i+R4kw
zTRWP/dq7SOlSMDJXbs77a6DIzDeesUhgBemzLJjidXAoUnRFhfTyHipNlV4CzL1
vpBTB++bnzXI8mddbLLP+1vI+973Ok2nqkfIVFPx222vs6zVNw2nwW2YnDjqJ1yh
o7XyQR1Mknau0EsRlTy218RiEI9XZlrexjij1k5gb+C2oldfrz6WhRSaol8duhln
LZWMRjb3OTezcYAqPb2DYCDfmtjsA0PDkFvRYepjK4285C5YV+S9aq2uLLxrmU4f
Zwyv/DFFMAbkSaJWi4MQ8smjuSgoGdxovre33XiVnR0ag0sd2INJ/95PD+8au4qH
zLtaVZLRS1LY7fmhL+3ral+u4H3qzCzg7CrRg0hw13lyhJ/h668eil8ICtedADxm
yqX/75lxUkdBs7stL4PElOKKL4Z0qbDRSlF2B/ikYTUmtZtRKWlvEetyzpx6aqv0
1lnSOZrTPZceEt1+SzbeFkEcANc3eoAogLWFcslr1udLSSRc+RKvd+JyRMpA2Zz3
ynn3C/QN2VbNRkK9NHMKhmqkAoePr83sMss+RvRWH+/T1qsCWe1UeK68EjGs3rG8
Tfjh/f5424Z55pvuXNi/GMCEBcyilBwhXFZ4m612M8Jtiuy5/8wkqM2ykfkmsEs7
`protect END_PROTECTED
