`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bBXJUtc9lE2GOzENjWHjhYsb9uK34QPfR2Io/f0j6nOsHhF/8HjfJG0YGAOY3XWI
CXWEUaDHeIBtscOnYmQL2JH4PleNpkuGd8pM3RAHC69PXIRn+ZeBcBBSXqcVmYi0
oA9+0oIYZBfHPxCg2ebk5mqL0e/LC7EzblD6NSEGfiC8cW0max69ezCMuQf5CBdg
CEjfIibDGZ4hDrdvnFSlbt0QMZeDkr2Vs077HDYZka9bzFm1T/S+n5eAff/SFRli
Mr5h8E3nixugt+6eaaLkhJh9ejrAvWolfYVkK1GCZqPt2d34oJ7zjxxbufUcj300
cVggPQwTjXDnn1Ul8qAwc4VxY1XeCnbYIowWQJonxrJrIJcCf1e6ATj3BMlCS0a1
yx/CrVI1lGKFOiZSC3nc9lePLo8gKtY7zT9Ipc+VHiQqgy6T8sfmF7T0tkCrmkmC
OPgQDemmiw9mURWLyd2hxJnkVk3+ExecmCTGagroKqLUo6o8Y4IohrlVw8Kxz6K9
rZafdlaLlJyE/lmJholEkIMI0NDLsI/uNfW9zALezglDm5uYXJQO8KkUuaHn39vn
LpPT8G2qP3W2m99D4KiC6SOODmNdNLLG2qxXEUf3FqV/zke57dRf1FWkid8pFWKU
D1te/Cwk4ZtdsIP8TMhEt9LiQlaui6GpJD85AFJHRz7ExHOjCxEowCNtqE/zoRIE
1/HXEpTIIWaAnKAcXom0EQMFz6AmcItZvoRjZKN7cevRejCbsTBtuqlPsBqNYzKD
4LmeH7gqwsyPQOUcrh/ElziSxGDwc5BiyU8gg1qARMrNpfRl6SWIFNQbU7hXK3Av
3RXN1PUIxcyHBf10gdD7AHERMNX2LzUgNe6D/WSA61L7IKG+HulyYF33l62cdaoN
JCP1NM7uUNTkVBT44VAuJa07jXfVDuRXpoHcFHY3vC1eruNjDr8HswgCnfpB1ZRv
QK0dw2nWI0yD62LH9wXTtSfwMrvoDIVbtEyJHxJVk+jYFkgZljRzWe2UVU7UzFiz
jZ6mn+85Xbj2NJFjFEWhaJuU1SSZDqDU9AwKpLqbD8PZEr09AW7IME/00PiIc57V
5t+KfIgNvA1Bc9Lx+BHiby6JQETrjyOe4HBp1XXGa1nWioSFg1I9Yx2A9asf7oGD
q18tceNA0z1mzhycuDrmYwBAO0jGeT+n/u/cZoSviAdfC7ti3ouAOEh5AQqpiX+l
xXRCTQIGvYrenaZyNzPNBg791hGh/rHMh0QpT75EFG2pljo/7KDiCeTkn4655zXn
ezju/tTP3wNhEbDsofGEEJRDGW7h1YYTBMrR9nuXeiTHCoI4RDrn0oWM/cNrkDD7
H8h2l6w9K1yErbXmPfLokbnkF4Cjj6MnpGfu5zF3GYbG4D2nENKJJQHsVuTq9/4d
0PciCrv4krVM4jsT3hn459pF+C8XMpZK+9KNYVoU+Rmaj0e2HvfKyGIJVrnIRsuq
lRG+IbPc6/LYs2Yg8XiPsaLW7GGnX8HwN+nQpPVVbpyiSEHmwtPgkpaNRB7sHaUN
u2XOkMNVxMhx/nn59evwPexgXr6B+G9OpgyJOHk8wdhnd/rw0RA+g5mODb0nd2Ou
seMJKGozZsT3wq7+D1CGAitL+cSn3kZ8GVVxCcGlVfrEVoSvt4MpHGGHclx+mUXh
cOi0moXrK16ag59ZYr1tzL0kNdzrlEnfOMcjARnpYHFilDCwry4a1vRX82k5lZXr
93HV4P0Y2HYd1anrURb3XitesgQhR7nxtQrb9sdBY7u2qQKYR5qIjdt96BtKRzBK
BrzbQpbHxISMkEfaSaxqD4quXwoNEi3CzcPI+JS/LnlgkZ3Y10PEdLC1mDMi3Sy5
LM9S7Ph5ieszw4pOtKLBENOZr9jItnrxsM90ic9f/AQgOXqjGs6jM3BekuB590RP
4khMDIe1Axnf8CbQ4n1XewD6bgiRqQ7ofeMbsC+3fdIqT7Kb0hLMFws+QVKkppnh
gDswspCx+I6dpthX8OAIltKqiDej/cAhhYh2GzcofYRQugnA2+eY4evAPaFAuDPn
Bft1w6d0X6FVDxw+G0TX818iwh+yJ7qdJjZafS02uWSBSXwss3Swoh8qvWAPJX3s
5ws/LrI4NaWeDcF+mome/OlGbtUjs+JqtYLrt/AlkMs4s6teJ2EVMhdTkQLn6pPv
Luk2LxlVs4ll92+F2nylUcQpa0XWxNt1d0hmHKBFipOL6tj8jXE1GKAV4VC6qgzh
tbZMCk3fs+MM88e2QmgzF2tCdPzQGw67ltNGC8zsBflIC3tsGR5hso4mHG6ec2sx
chZaTl+RUkQYolA0/MSPGXgdttmsDMAvcZsxnbyML9Fz3aK2C9mv0gBftiztJRdA
momsRhJ81FfT05nYodBIUGA6+ObyFDcHEGSzyLLlloM9hqUVjgabkG/7NB4lge3H
5jMdQSadXxHjWFCiwtmDPnNSmvadWJrhbGrcpSZE0IKJyP4QSz4pRWreY0iH77hM
F8fFxLH2X0YxWQXvu5t2kw==
`protect END_PROTECTED
