`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/xc+G0zDQwtR/sK6mNia899EDcv0kp72N1BELfCiXycHWgpRSRKspF5NQqcK8w2
nFeWIJBuOxydpTtxbrbQ+hgjEprqJn6UvTi+m772VIc+CaNY/NlOf+Y4T85i7UU3
97AtgrBOdP+KEAW5O0g4CvTxoFNEUyug193blx/Ffl8HjvRMhWFASJt82JoEhC51
LUyF6IchGSyPxhYNHEK3+odTh8deEIaj2svISJ3qALq6e6hwVECQvXJhi82jfFGz
His533bm06aZOVi7ssMlAC3vR/v/enq4JwK7bQZMMN0iiqslqYlWJV7liWcPb/Ka
IBmtiqXetXk1i5MiBnQMwSIKpLOIj6nHIh+u8liCJk1XqJIQ8mElBKNhvTjdUa11
4irgRpNYDWgC9t7QaeA/vio8I+v8AxAjYsYxTpn4T43aCivZfNug584QrdfCqvTF
QWQ55sFU7dE7gKwLW7I/n9e6WIMR5ClL0oPgCUzCVkHVG0zuu0veyT73F3tb0ne0
yNwTD5vhtInxa+j0JNzodn3xJa4jyhecP2Qtb4i46xQwM4cttfQo8IS2npr4SyDI
n1uIjhYxlzPA3MLr+s/94n3zg7pJf1dF/1DzC2npse6oPATWHZ928ONUl11gbUkk
YiEmPBDcgaj04JfVXDqDRy0MV1Lab5ytPki6derAoD1zegJMhleSN4SCsW+kXo/I
X5ZGK/2QhTAY7tPq0XlrA8oLd6hLL3bh14sRaJozNdWrlcOp8oLFXgQ5oEBEURgN
A15tP2elxRPqpPOY3H/bFeZVcuxrU09czp+7L585Iywc9GtynFaT2IK+EuJRZlXO
NMD6wQ9ablX7kc+nLMQEq5riUMD0pWqYpQx+JkMG562VFu8kCdZgrt5qd8N93TAI
xnrs0JWRyrDWqHO7XtDWEA==
`protect END_PROTECTED
