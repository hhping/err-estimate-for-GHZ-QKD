`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xv04YjNTqQHspx/4fk1JVtBRJq6KJcx3BHCG9z4BmOPqaV2gHUnSvjfDdig37XKh
PykE8CibHo7MeCwTgnGLs/HAGPc3kJK7tA93yFRp/HFvRoT/G78euYW9l+k5QP84
iORptcnskQc4M9z7Orp1KBWJgW/Jr7imKpgipGvEGMJ4aGCfGMTBi85B8yT21iaP
CAHf1YlQW98Xa6hh7ykZi1mcBuggc31bHegb0CKuZOT+XDbNAnwJhf7gNXmndoXB
plriCCc5TGwnXDqQIdIr4coMeWPFgroyUC5oqd0BTlYv9ERt+2EwQw7qOLojVxfb
M44xaT0kf9o/rAd+lKGoPBKEmSzDBMmkK+3QmwzlWlITlHoP3tA3mXyy6rlh9CbW
eIzlASVCPG1O85e+pfL/gEX94eiesvn7xlbNKZSjsE75p91CWHneAYEGDjEwIIJh
yYjaPk8GdpMJDyTrs0VKAJcE3TNKRf2fQ3NwS/o1Xu3QWVU4yaKnxyqqpMc/vonn
2SK5Cbo2N51EvwTEzPuIzq2ohIDr9rD2hY0ApFOuRySNkMjNWJBKzXvtuOUorZ1l
FN7hvaMWzvoXRScAs2hxUk2PnwqBB02WnWo2mKBGQEOFc5WePRdCZYwg0t4RWcZ6
SRtn4aZYaBrsv7QK/dVf/yNNozk1AHsPQLECAXPMWZvDTp/hYDwyn6Hi0gN6LkPl
cD2G9Q0s27AifA0lLu2p+jK07TC2k1hiXRMaoh9erJo=
`protect END_PROTECTED
