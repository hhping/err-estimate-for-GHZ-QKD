`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oA5o0RtdwTU8tXa+ZFp1bFoP9x65p638tvUOX984OaoSnTVkzRQeUTtQP3IfqAK4
GUOvYiVlsMwDr/T6Z3wiVmLLkL4geIrR597i9UlF2Ar2o/nuQ21E8qtAP3+GCWo9
6rmieR8M31bgvfL89pJjm2Vul98rlwX65mtIWTw38/fQLOPe5Sftda62labCuXks
tBLuhicUiwo6n6kIQGZALXO7YxXW7CjEQTq1SwAeu2PlNDXs6cGzr2YsnnHWO39i
xl4ORxewfitGoml6OSEUAS2z1QEXAXZg/1+tqNYgzd0iFvlqVIORibiE63TYhZOk
08EzV8msv2ixNI7jeJRuCRJlchVibjLm8gllc7EXWZgGY7SQVpbdzv7zs1gJ70xh
JDqWlWv67S7yYo1M6DLqDxhcNJv3zxTFVynMfESB7va/4nAQeAq4h4MFZ3mo1t9K
o6ioNEqsx6VUkdGYzhO9OnTd9k3nvieDnN8vSJEPabtqa+6NHm0I8Nqu1ixS/O5v
HKTDZknPZy3QRGIeHbN3Fgst4GXFUkPP69a/qFv70okB7/NxIS9aYhHfuVuvSQ+l
EaxJI2NWCF9UxLpoCpa5GxKdb716AfeZAMS+Vu4dman6n5idIIu9B7VrNEH6sYu5
Hkjqdxn7OYS90ugl/J5Rl66MRpi3c3+bhD+qc6rtI5uwkyAj9s4RDu+DjEMtte+3
WsSdRjLAVb3WRq/2ayeAaWMNUCX0plwJKwKrTIFOE/yr4sM57afbYqSkJPJ+bvDQ
2OwyEJxh/IyDjWOIUIFDP8QpwG+BfN3PV2It7XBHmx+IUIMII8zqtpNEQIToQSn4
XtIf7VJNzgMB2sHbmqEEDCW8+a2wIxfMK2iHiM3L4meWVUWKsJ0nXO8Bqb6SFOox
GR1Hx7VgFD1Rc6O9EC/fUpEmd5pg4o1P1PYfFRUGsq7uxVyPrJtvel/P0JFq/wlO
q287fcSXjHuZwX5Mw4+9Yp2QctOxn0eUtXk6kMXYOvY5glIGMwRO4gKRoZJEJsC8
FA31kc0bjk/OLyRlc1RrKm2mPBqDmaKOU0BoXLTHEO457mWdlGlmUzTl7PFnfZIS
PcPuM6KkxkxCFNj9tSLUDnsJd3umqETwVdvdSBP2rhdv3KMMDBT4AIiN0aXbw4rA
fX4464+ZRLuFFK/QmVJT13A8P14Gi6HyybKh7LArIEbA/TiaT+YixVG9SkvKknLM
PPhfKWUcl58xabMjagd8LhkzL6sGJmG9WEGSfxybDf+KRuX0ywV879n6TNzCcw2H
F22Dp34WXJAO0LAn9u3lrNPOfgLwUW6hBbkQJ8BSjJHS2b9vMXf36mWduLztllt4
w7jd3Vgx2kwi1s+da4tQdKAd934INZLI5tULNQphDMIZpqzLQxi+Ebniau/BJ7I/
Q8ezAd4XtYu4tTvcxFyZxGonTXl8Lff005YKUYXquW9ersxbhww3sxJE9L4S/snO
RYwAFtwGOhh/KXODEbRiTW4SeTyjTCBcPf7pCxWpAdJ0ShOdgV+561FC6nmM5QBH
o4WK6V7JyncWccBHDGiecU+ma8qFAxX68T/c7vlHIrNed9NB9QnIvS6GEDgni5cQ
k7mbwTqciw3XU4Vg/eInZ3wBGui21BfcAsqfvZCbQzOLA6i5RHcSW+ZebwsP/nhx
w0Xae+H4ukSH5bsQcPPGAjQ3Efsi4djCY/uGTQqtswPwG2w9I2noUX69LwdT2h4P
+ok+TyXLNfhjD7hgaDQy2WkeKdNIyUVWG/PXKtRUtDoUecvUOyVrsYO4H+RNMc+W
QGQyp0w2hspD5a5zMIbDIZ6IYIf+GE5JIrtzLRxypN/1W3O8AfUOJ5TMrh3PS9/D
tMZ+NFm+lZ5nEgm6xhBZ0C6q1Cs5RMioggLivBL5A6Pf17T4b0cnF4geNXzL+Db6
17+TmollVXG0F6JFG14sibRGNN+mXvP1ZKD7J+XguIeQfmuo1wKDfxq3dLG7HxOk
nF8cTXpDTUtT0+oHpfOYdBx9/nKsyrsmddR3xr3s4bKo3DnFMVXEcB8HMAj7yx/Q
rhCL8hEB1h1qXL+ZCNZmE91ZYofb6HQ7mf3yYUWGquwgNGuyT0Q+tCu2As7DqQLu
S/D/PPvHtRdU8Vmh0IUC3bF5JfjAIF7cfc7U/LkoXipZ9+jM8bPKRcY/hv2RfhfE
a49S0jZdsbKrrSqcApaijnRdV8iUUrTUTmXt+viTE6E9Yud6ruGsrBHt0YR+cIJK
xWXdu0H6X+tF6D+Ju/bLAplmglSYOaTdvVmVjErlYBw6V5cbLJcNG9Z4/b9G0AD4
`protect END_PROTECTED
