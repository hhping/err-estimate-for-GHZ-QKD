`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rz2orfois7QY0b2XarJpisI9dtTestFHTaZhf4hJDWSczH5jXpXPngMex5IGngP0
hIoou/RP9jkQfQ7eCrvZ8CGBkg9noqZLuwWuATwkfhHL99eifvSdpgBhGiZk7Gp1
hxwEE03ZCca75ZPgiYfhnpokpKixxFvEFqL1uolUNGk0J2/fzsmZJCthQp74e4c5
6srdzVwshX3je3tLcXhwLDMZx+Spme03S6dEPTIzHEcdeEjxYjLB6+H/XULqlekV
yplwGkHRgXIQZDIbDRTtkEGtJBgv/Z16FtdlyeBKF6CeGkONT1RspODehH9QBmdk
mOBclY6lncmB538XBQ1sAPbiUYuxrklF+tWHrYwGEv7er9I7JTienXJrwS+He0FH
uK89URkpEw9OwAQp4PtnIrL1Viwxhj4ZVgUaHDEDehB7BzUuN1KNyVW36hgeWncP
0vDUC2jzrZxNqJoOhlQau5RYvoilW1BY6AIaRbRoqJX5RUiAEgUj3n3whQxk5z8l
k33SXwHsXApazWPEZ6UvZxOig3gKgbpNVh+8Pe6qTNPzEW6udNEvLfow9C/Ajh3t
ErrjwcxkXtawR4+LyEposTiTJecCXsEBRgatPfeWdR34HzXl0bOacUrChM+UuC0h
yk36uMKvpoFl1V4IPxIFrMnCzAhiNCYKgR40KDiFpWUjyKfpY+mKj56hjVy4neBE
EkDJAni9bXNi6p+LVMIy41sj5/NHFPCi01qrXZqInMLCL+MwTWoOmVwnRolXC6Ud
Fx2/OplJbaT0PQr01eONPV61e0ejKfQZ/ukGXaDxl1dR48iYS+kNrPEg8krwJZR9
hj+rlasTgtSJkE65ntuZL8Fv3Eso+T8PX8emtgjFvRai88NUih6jwktYloLXGcnT
DCTO3faFy1ZSHg2qFiyJGMyg7TgE7QRI3FIXHnfJ7pLRAdKchLefn5muE57lJBmi
hdOdv5m/0mZGH6rk5k1/EY2so1c2qWEF+6mAIoO9xBwRoLZYonDYo6TZL5Kxn5Zn
Krfq2Fkb1XvSWDN1P6sD+cXo670bJY46PY7mM8JYDF0Otdw7mP20lPEEb2eMQP7s
Cqj1auJq9amC7euL4ag0e44wgnCLjYCGcmRFwc+a+kV4opeph2IiyXI3BlEwegtR
FodPPDCQC79YnDAzShghFBsKLmo5Wxmsavg1EM+28qNkTA0cHHA57Wo30sNPgLof
MQqkfuglKLl7oKsa38JdpztOFsLVxDl0OAlkk6g33VECxDtaIugO63tpPU8rdMU4
iZeYG9d6Q3Rm2fHJPVO8YkXHYtdg8jBoAk8bFP36dITbXzW0SgKlcpUVLuiFENqt
Zej6OoFTFacWb1EbPo9EQSpNAyVOiBtB/mrFN28aJt+DZvrq5kANpdxaRn7pICJx
hWa8fLT6x7WUpSBeEFmlwBrAisTuIi4UJ7w1kvuADQ8MVI5sRkixZaRaRJ0ek4Cq
is8OncbMUsUdbiKnm55vgD4U82nDHmKMSQmx2RjK/epTzlhG7bPo1YRLe8/hf12w
gv/abwNztfrOVvQXnGIvSuMagTxOtDjfCbUHPu/iXgJA8h4/e3XurzUd7DIvN2/M
Yjl6hw/LURL5MK4UZ9cD+XJnJyQ1aDJsYVjMJt8FQ9tRuHelo9MoHBYCy+NFhdzW
mWYoK17O0HcaHHg3k78siZDZVQCED7KZVRPq8OBPqUGScS+1q9xDA5Rae8SZDDPn
cDFAK5vUDkM2wxAIoGbKz9WF4yPu3ONknJYFILlTDcQyWAjhIyyL9NXomrCZ/P+O
S5RzJ6hdIlzwZZcc1ZrtSPKb+avwrkt3Q3TTpZPMRnmCKOUfrH3evbaoVZEAdAnL
OjV5s4e2p4wVeIz37P55MAJZBzndtRkNS3jToIwq8KmkE4oiriWK9FJ0L4DXeWCC
Pk0I46B7SN5wpeXXwWobamm6k1jS1hj7bIcmc4esr3M3ZyBWEiTXCH6TGZggpSu/
9T1DxbyPs4VZnU5ahIZbUrrvDgOm0bX8kQb+xEAermebI1ceZEhGlnTopabOUrBy
BEGJW+70ukjC2bkB4XvTtnrnOU9ZPkBgI9uXyGmCKteGPVmLZ2VBOPhTvn7Bg/hS
dzIWMTium9i+bBEiJKn0T+waZo4xKcbFeCclgR+zkEi2aWVaSo7U9G2xpjJ3+65i
3TM5G8IOQ+yBpm2QgtyW2s2WaZTijPSL73MnrN/bRyvbJLzeObe42jXo9LgjfqQg
9Ks0Rx1hPL7RkP9IYnyYoqvjIEFd7blgvqWA4MB3pLeYPgAW9jlNwW2nBvKMlAeN
mW7xZN2F+P/qYCFm3Kn1ICsuOQfOYBaoXwKyZBbmJalkjnZ0H9NKWYo4C9N/3TUa
ynWm16UQqB/wkJUUZU3gWuEhuHksU+eTCx7UYkE/sg2Zy1yidQv13itByX7t/Qhe
Hy2s34eFccVMdpNDQ4gyJJjAwtghB2EcGJOGAWGRMOkG0laNMlxiF6hmj/YCXFQ6
NNeRbab/SQU/PWdTxGfAHRVO0Hh0OYcgjuCRg+w1y0hjRe2OQth9blxrIQsbZ0yt
d2TsGwO3re0swywgufyJYQoX3SfVdBCBkMyPfK65+FPj3FuYJ24NdX2e/CYb+GXD
tFQQqoD6IMlSOcm83Xu0wNWjSJFed2WhnAlqZ1skkGATJ57xkZGTg/fPmt0oWwSh
ISdvrZ8ctc+J02kB4TC+aGNKbNS3IxIrrcQhNTVC4wcvNil0jxt4iysq4TEscF4l
mFEfrU9xitucjKBLpAxKwTBindJthsSbSYsBZ0CXTq5sKnFmekH+yw7EO6FT6PSF
hXXUWxo4DEW7nGHEYq1zgyVrzgIiJSfCIchQ6MaUgpU8IEch65h+s09SLgF42ZY/
dI9Gpd6sEWPa6kKZ6J4Occ5orZOls9FjAISSgxoxPvItIMiwNYLbAdUg3Ok9LDu9
j9bpgacDHo8Je1KhAzBAX5LaKeCxs6Ow38zBks0M1F885jO//d7AUw+Waj5RQJwP
Wz8Mz8T4AZyUmkB9mgDGow16GOeXDnRaf7mcuez5HdlZlR4XozwqHtGBOrUmzGYT
c7F8+cxHDTcnZi1wWh7zb5q1Pa/5NZJfxSMtNl9tR83Fgs281QeThRX2Y+II8Tgb
LIzOCNgKRLeu6vRABHnUxJR5wvYHQ3N+Lcv/Gfl6luKv44lk8r2NBnco8O1zxk7C
tgO8c9g7Pf+HVlvRcqbQLLXCSJ6YfAU0a+OQpZt6qDN7Vg0gEmeK8RyZCI7N7A97
Zva+ong51SgFbhbaLoXoU6eYh4FWamdP5BRJ5xierrcXYPEzR6Epea6HOgB+QABw
am8ivHA/iGlzQnVCWLT2TLo1IuSN9K0QoosqVPaUKsf5KDst0oc3HRusUsOqg+e3
gXrsSk4vNnRmfIwBy7MufyZVvd03Lbd4vMICBmXdFXYhEGLaqMrG5nt/arO4HaWn
kR/eJXHue6r8hKQtYY9mbfYGh6l27a4mygMxdfu9x35uVF0SRnIRX0vrPejIKLDs
SA83gzsvtm0wcRnXithPkoV4TifGwDhxayyMRmJIDWvPeu7fcXmXl/RNN/Jogr5t
yQOsK0f6LqK9wKvKxZsAkE79iiWP/zF9JqNatk24PChvROvqML6Ksl3sfBGeCFWX
aUt6INa/z+Ac5Fg5Uwb3BmgFT1sF8b3t9qS/t2RajNf2UyW/jI/z7Nf67XUGhISC
g8Z/KpNBVhYTtzUnIbw7EnmpkYAEmyF42NaDXbXY+8LZVdXVNzABuamQFvHdVSZ6
/mfUX4SAr83vLrP0cM7LOBiBFkn2EPFk8/G+NcGUhsu2Cumf/cuQrOq9uqMAreLl
OKtmi+w0q/U7MURhwFmJc1iyhrb1r2E4D8bZmQt4C8ubP9gOy1I5ZCctIjCnQVgZ
vbMEL4z0L4tM01U5QLNppYVHkqNx24dauyRLOrKCIaDVg7CRtzHxLwKZY47nyx3e
v0hd+e9YjY6AamFd2n5NSJbrB/72r5XEEj/D7qfIwwd6SJed+uli1O3w5cFo6c1G
2ppzycC77MEjsnXLnlUEtpmNa+TyQRDaUJ8PltcqC36u9W4WoFEUTCi47125eend
K5LiQpnXf1ErX1xQ2eRwBUP/1aRMt2W158snK/iUQgyZBOJmKfh0u8BiMz4F2VKm
Ev3QkU5USp2EOb6pjKeGos7QxZ7LeJ2hhmZGYh/YaVSKFRvvIyA0qVTHttBCQoAV
yhY+U+leWeyv154/WkoxdwT0izv9s14Mh6GMKZvfTgSbxzl+XGiE+LdU53DKy4fH
u9Ik++4+/dR0CcA59alZR9R1gIuraq6edWh7CA91xjly1/a0m4HqTyUF7emCQP1P
vNpuKSR+D1gliW771m+ILFWjfoTEFBvbEMzY6D2YI0V0V72Tgia0FKcJdzZSfFGu
U/vRllyu10Sru8OYuLLp6NW3HHcCHAkiJ5mede3BJaVVMLNWh1PRpAmTq+n7+MVZ
xLgsCESAB0lQ4TZIaq9rCbt6ieVtBkGsO5ZKRpEHSxvHW0pEpGItOGLCaRaGbE7S
FB6nWhAAmVsshXhbo0JPtg==
`protect END_PROTECTED
