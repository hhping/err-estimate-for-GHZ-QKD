`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWoYbE5GwnVv2wV/ZYzMuAmS7KHQnEK9bAYKYIVK8NbdkFZ905oqEOLHzpE4B1LB
gC1YhHMRfoBQ95imUnPmQoWMFnhrMOevMfY629nswnrUIMGrDNP+YuhUmHoDqGpP
cB9V994GVu8u68W8rjwTWvnhG8qr5I8KLOU0vc5jVy85ihhT6Ts3VC9ZkWy7oEH3
07ePht+4oZN/YaTMWpxiPdM2NAjDmBWauSJVB7lyz+f/XXGjl4tfZ2HL/CiLT81M
Q9nM3D2pfcjdWyUZLPTHmkgwWetitajPaG3J2Dz9vgyZF909FNfYPA+XLJBac9dO
utwPpX/qzkAFoMmly9cQNkOqsasaC/IrLiCO7r6YnpLt4kbT6SKPcPFauCRODqB6
8eo0SFnz8IaK0gZSY9afqQ==
`protect END_PROTECTED
