`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6VePwdezesROULV7TQgZh9/yQiaopU7iljaMd5mPlfkmpFBWsgNT5KfHHblCCkC
pNRkRh4Qazt6PsP5RSblQ8f3vg0YXArTMsCNwtOADCaJXQanTcIq01A0hqjqmXgg
Nb3kcDrvmGL2J0UT7zsa+E0tlqTU21bS4ziONOeZWyitn+rvDtgJmPmiLlGaKak7
lgUN+ml/Z8kUHcE1mV6TA5B3VGtkzCzK6M1kuVu94oc5sROCme7AFZxoqhXw5NW6
Hk9KcAltc4BpKZMKzwemyPZPfZ/SGDRO8hlWo8E3IRZKWc2MrObRvEAIystZHKlz
QvfNllktigLDZleq7BPs5dy0Vd1qxoBbypoNUJBciiy0N/WIA+XeTFhwJYx5wdXX
ywJ0HaSDbDtO0m30E2nC4q14s/uj+PtVXGzkKY3JEXt1LyUBDeDinX3Wz2nCCEgJ
2FZZe9uq5wEzs1lgbcnGdZCdJR+AfPy4MdwPQIZR6dmJE9Smy1sek/h6/B0CetHc
iw+CJo6I2tIbnuoDxIn6nw73Z6wSMyFU25JVD+clzoxvJhBV/NlLAa0/dJeHN3ZA
2V6dBMWfJC9Cst/QOveuNKw37Vo1RDReOzuHnlHO4CrJ/sy0kqLNdyp/QEZYNPwl
XI4guUM31EzktN2NuZW75SiOGdlYMOpOXFdUq3iHUcKZN/PlOxgOfcOLRCNs7vzA
Sxt/KLOBm/HLhkTSw3wHy3qrnnHXForW0RyUxAD+J7f7I4WmJmpY6VoGli0mVyjm
E9PGoEwb5daMlgx1dWgJUP/JExZswUscej4y6oIxDtmBgsTItVXjPKrM+pIgb5NW
4wfOJCMucG8s3LlQNwdM1CdOmZoK33+pwZ60t7tge7WfMKzbl6tn60bzQiJ/5v1r
/8D41U3TiZmpDfaIzCNcPJHwIArNocYrUd9QM6HrcUI52eMtJGF86RLj4uXPIIo4
SL83TgGKkPOP4j2hPGSDmo5KkX3nJHUfYptt17T76KyCxdVajFUzCxuRHPy/+9da
YUwoljS19ksCXrZH/B5k/g/Omj7LSdzjPf2yZa0umtNHuW2LIp/t8MxwmVEke3wF
gumRe48sDFSEJ8llSzmKl7TNR35PcNlfM4TXo3vHbHzyc9S4tKNzFMeIreUh1q8T
399g2uth4fh7HOW+L1B/RAyZTPN7lY9lHdOMj690HvtjhVxgCQR/ki2eN9y8M1Cd
2Jsb490DDyP0Tl8dZ/Mopg9pvIVrG1YREbZ2E08TV3a+wj1Z1e80KZ3x51zf093M
64KM3er4/Wnv5N6yHOt7upBOv8xd+XZbRet65CSyoxriqiN4ssPAPj6KGYDN74vv
1E4PgFS6+Vc5bTih9eLxhAO15rtZQiR9V8ZLv1ruVWJSrXeH7TVUZfp4eCTz+1Mk
rdaZ9/637IyxlN9CcxQAtzJTwp9Nc47DovkI65gln0lzqNJBgrtnnMseI6EzXFQa
5ZpRjcIry4tqp8iowY38aRrB98/d+W6QiRreblsvE4EVgRX93Pq7JXfVcCJMFmzC
SCrT+gNjWOCQJ3/Ve8dY/d0DtVqcsNrNieDqf6RkZchVulI699GN2pHUVmafZ6/7
sMFenEEuC13Ht66RjEDd/Qvu1803OL3taUGqTVCmphOE25TYeKeO2B2AMlWcTHZC
uX5QlJwtoLxsAFC/Ppkrf/v7NHTdt6JK4cwDxynWRSEzysQ+08HZGwMxnThYCYtK
`protect END_PROTECTED
