`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9W64BLVL2Lvs8n0HAcMaJwY8WkJYeZ8pMhJyJLjHLBRuNZrPuQQx/mJIpDIMLc0
yTs+mop//puzn+K5qrCTYzhvfCjzhXBly0LpJqrMj6CgwarCK25PICwEQJpzza+B
7qDAPUy9MGbMKv+mmvZq4DgFId+t3Y2fQ1ZQsYm3eJO8RS9Uc8NqdNhIfCezJOb4
pLXkfp9IFe1+w1Qg4exgbvy+nCEeI6B1Toj5dUR/k+lFgPAWYdO+n0F6qm91cyqy
vt9PU1NHbZ1EqOtm/SpXB5K2DO+u8c8jmFia+ApP2SGnFBXPl+q5FWUCq6gZbgqm
ePfgrWSvn8gAupbbMjNk3yKNrqTMjnPLvMRT6dhCuD90NmWmME7Nw9GWkMyfFv6Q
JCKXjWLLXSBFCr7fK1anDVO9n38WPkCwJDA9z91vg0p7lI3iHBHmuPCNtsOCcD+O
4omd1ztI1B5wxj+DI6nzzuCXkyQKRMmOP4g3yY7BSfMMnlx7FtiPthA0Cn5EgJJR
gVUdiMp+EM17qb2aR0l17XYJd80VhvwwCVufRdwDeuRBx8eisbmWNreunan62K6G
rKNNaO33bHKCU2qR7hsVQEfqmbryrHsg+X65ZZT8j/9FHMzlTYm79Kpw6EiPy2fi
AsPWg9K+YirDH8/N9ElGIIxKjxeE4WuDAkgixxSwBL5ySZcDoUjSCp2lPl47RoIO
EsREk1Jre/baTHZ9gx8kiw2ZiqA4Y+GqZFU6Rt1rgNAgCK0+ydBjYVXd7Tf3iOnw
Ma5tWGaeYmjkY+0xg418hN8f3uNYHvy9g+SJPGWfGaLvww+pKO2bo7EEGw5i2X8L
cACadXx1znju1haiQt9Fpw==
`protect END_PROTECTED
