`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhSPGX2QfTjz7mZt4CdwWuWNMB3d89w6M+0qpjLuxwtYYaTDYZ5pEuY7f9AGBmMH
DILEuBY3URXix+7aonpYwothIvmcDQJDogP7/zlpb99PPnz1QZ7sKV5bXp+txTd6
bHo1FdIEytVg8ZDC50j+lbexBdY+2cQX9nVIV20DSktzvlRSygewo94gSrLRZty6
ZqL4tbmwiEnXL1b29A1uo2EBKzmetS5ZqC6EgfF1faLyrLlGAf6kmMFyUiDOvKb1
zgcljhasvKJC42//GbAQSdQTSzwG1v2c1KZL7Rvgabwhv1pJLGzm/5lndFRyOSGi
IiRFDfN2usb8kKd4dKhKfa0YtwCpdRfBBtaKtjW/PqM+ZYU1QV5NryiBUVTtn14K
kJZT6dkh4pAljFnbTBLbg284RaAWF7DJg8niwoyTmQQzxIn+Ld9aiFsSCWau94dl
1uHi7BDlYXTfAu+WOZu1U9bh3NnfeC3ymIlMPhlBBB5aBgY3E1yKhEew82bAKgvM
haJFbjqr2Q0GFmFn/0B/EoQXSOlIlqlKPRUX88VP6hc7xYXlPswewYwllIVC2mDx
aEIaK//MEjTSxa6pN7iGuUOo1QSnO7jz2DWnDBZMCpnI28IlYkq8qm6yZ4pQqymC
Zv60aDUsiF5ypSSdjro3KTcLAMoCVBsQvlov8oKwb8Ko4YRDWH4q+eGLZEb6q6Cl
P/CLZyeWhHoOZOyBA9n37A==
`protect END_PROTECTED
