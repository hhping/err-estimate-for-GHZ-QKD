`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P89YcsYkq3Ysh4NWMCRQx6MlTVr7G1WSMhvXdvq1g5vnubrGKm+Gb37NNLobyERa
7dHDhvTAyZw8lHwtuGbA3fXpOFuXjHqJXzh/e3r8KCOUConEibuhQqG5De6mTrV9
78kEOSdJ3ZA61nt6oo/gIQ9jeMe0omPAhXtjDmJywgH7li9sSm6+53zPPaDwMH/D
1RBXUtaH00rsJw7j6i5m7JCUTFLZtA7FKfWcLpe42euKB3D9DAkVaBJEJkIlzvm3
E9TU8LGBmluogtjQouqNLAKLdZ2Iv+bH/vzYU9DQ+6L3xtdZT96owS29QLMMyYeW
jmhpyoGMLGWXby/3mjsfgy+GiDvPxI5rC6UHVLW0VelEnPJqmiVsM+CVBndslVZX
ODCDDd6yZRRTv7UuxOQM5MtY0PqvoZ66TpMQRwFOzV3cg1JN8bZPofRuOe7OOyUx
VdGGIdHj1CmJKlYyIEjn5qPM1VQQlzNGieLzWASdnKXOwQ4NALsPcDoi8G86jvZL
Vev8n1XyrnAjchyZi91Ar+uqoTgMnDwx+LeipJQ1+S8DTUhPVlI3nqxiBVWd7BFK
O7/E4hLyfsZm1xQvr0yQ3wZVO60qmX4/EtEhUx16+3D+Y5XiKNgcsi05GAj8h3Ew
PXnFPL/S4EkPnG2ERNd3StdJOr1exiQtuhc9QKNcDeBclAsnjvlErd3rhi+jW8NW
Gextk0kk0NnOme9nODzhFm62mIzpFQcFsGiWYLDNd4TIcJeYpmSTacmLVZfuLu36
Ghst9OQtREf34ceBbHaJB0zfWtG4EWxFGDEYiO5LRH0MhgA16EB+J3cwpkiUldEn
mXEZrOqO80FNI4DfnHma2VikuBU+AV+W2MKVjKcyS5fXKo0I2VS0hyvjq/g4Uq8m
XOECeuzD1lDOxvKY0ZtzyOwPKcc6S6UGd+JXFafxrig=
`protect END_PROTECTED
