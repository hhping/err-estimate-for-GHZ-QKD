`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RIG6J33JDqlrcuVGvquGC2GkhjfvgbQUuh+35lzxtoRmfVkl1uaZuQsTotNWZrO
m9g8DVfDu+jaKYN/iL4U97ZNnW1/s2wYTVZpK8RkGTuJgrhJ2VMEbxtaSRo1ye4g
oazJSJMD/qKh8EqUXPgrd3l/dzB4Wb1nj+ZAmYIpoVQ6t02ZiXa45Ixj+uVo/JXN
lN9u9iR/NSbwaKPsNjMjv3RtzpTryftbosLIAsyNNnGK8y+PpvI1wJSjyn/sJ38H
Z0RQsZk8Gd8new/Z9G6EbDqBZGfyE3ipUg4I/U4vzeKHFbyRLWXfNAVtd/UTt2PO
gOT6Qm5oDPtqaiYh+Kbz5mdyxnkm3Y5WZO9VgMCFdNDZlnopYaKBEE8nK3sk20kv
XT9YOAQwivc8wgX+6RjzbrkUtTtkk5S/V3kzkUyziLxQHR46SycTvsq6F5q9jvbg
8JmjNSN91z2llo82iZoPCeRNPA5NkZvmMzVPKzrW4flNo/hjZGM095HX/38U5k6o
e5WTrHiTLxpaFdwuRnZrdpbw32ewq9K8qJMfBu6b4n9cSUfm7+upfnm9D1RFLNkf
PZMTv62IR3+F3ZCdktUW3RBCZ3CbyeyTia8tyyDQ+hWKpNmOhzKqbbegyJHsEPYk
amtgHt7QXoBXsaFoogiDbz8XsbPtHvT99820ODTW7g1lEmwUP72BziFCU5EPUh0T
OETnmDPJxefVBUyBPMf2FGiuQDjfd2cuwXO/5Vbm3L5tbrlLK06wXicyhPGdwKu1
x8CHA467v6zVQCWkZH1x09QmPRh3C10hniIw6OIIHHGQMd53elfpvN0lyHi5frbE
uT/3D+kxFn3JG2PNn+CN5CqBH5viUtSq3rp0Gg0ljfOZfcI0hnLHZq78o/h0nCaM
3Fw+VwWBoe0ojau9wOzf0zL7HDvEvzVEVBUQiWE2N3h9ykioocLgF4aatYepqc8d
YVtYNnBHRgfp71lAJypMqu3LT78JRaSB6lmwHsEKApixmd4VFHEadhu6TAOOadS5
oQy90p2J5Eo08ugYcZQ7aOCJP1DzD7/uPW1a6LL4/4rDEitU/9xErBSf2yYMkmhk
BmFP//hRpcwYWl5QopPXRcDTLpqmTytlPlxgLvK3QRcn29OhGgFFdMMt3IYbTnae
J3HyF7dRJgP2OQpUA6Hgxoiymmkqv8lcOMz3OJq/BAb4BWOwjRaXUuom3KTaB9mm
4G+jSOTWZY/agxLY6wpuBclAuR/WP7xGHDRKsp1Fdz9TwVwk/gMrmkqvApvIq9XH
bSK0sdPU8gFyuPp9nOARTDGepoGwdQpMhsIKwH+sUchsYVc8rRfPZU6yxZiBIalK
39IKGupiv2Fc1bfEophCsPNCGrcrOTSEQ9DFkqJpoJ0cwoX4+k8sGf1X7vuc3bbC
10upllUAZrF0Qf85dKRaUCi9rzMwFBguVKdl1YLhCJcqR+ndWjsAp5VEjUhloo9r
uXwMI4rOX/ObNB++GLo8sXieVX2PoCgWgsZiBZFN0ZzvOmttJX3arfoLUCBsJYFQ
7UdLWoTosR+88MsWkEuq0QyyXhPT7dCAuEd0PRaoJFvcKlXL/cRYPUOhf9pDndzX
hu+l3USdG8qNnep1TFduM/mvegPZxlzDAjoDzFoL/IO+6jCun/7X9snyrxUMBHkn
O2lObixU5UwlJD2WOXMyiWADW12RQDo2hROHpFmLH2t0tSIgYRhx7WdWajWODRql
HcPn6JAQ0oCnSE4Wb3mDlA5QVI7rxO7BoEMkkqNXJy1BYWsPswTaHDp+fjYAklDk
+7Sqr+9Bj8zGDJGei+UhBYtzxUEURaJtfF/6eAA7gYkKtCuS9TB9y7GLgA5mKqHb
ewxI3EwPwtb0d6LVQ1goVWtexCQDbB+xIX0SfC3IivyL/UWbMq6fI2I1mHVK+xDk
gx2useAkcNHMhyOLCeTtZFi9ibyDSuhxn/jtJMmj8kw01bsojIu5Ml+RZVNPQ/kg
IBdU4vWPCYqRKPXOKAwG33dWMsEbkjVjXVZdXEw/bz72/QQ0w3Tma65ghHzpAGJi
iU+qLwEEEsm+DWdSZwNfDWq9J+BzfDDjwAhCaCzlvVOniZD/QrpX+SQASRGGyfFw
4L38Y+li7EFL+5R5lxO4/zh+fK+zX5hAGzD92Jlxn6dmtE6CME0+irEf3H0KroaX
QWLJH85oK3vBAiR+bvGp6Y5Ref4URoNJD9FwhX0roL35g1WmNjWnMudkSli1rXn+
2qQs5fu2fRIHYdmPgc6JS3bEzGwLq/3L4n6B9gSD/vAJpe1hkZ4LBEezYmX3XjuG
pcrNtgzMyCYVuYH2Ggfx6xwegl0MAZGQoSBBQ8053BWuYlTkRilek17wBknvADFF
v4W0yT5vihPXdzuPvrBxrGlLwpCePWr/4H/zKC8XrRSv/WpU8cFN398JGU7/O0C+
32Mbd2qoCW4JRbwvX9Pnr950RFwV7Pz+Hv365QRBKaNY05FfBSepx0OcJtpsyuIl
+t1EiA0kpGf4IO7tQBkW5gDxoFEQhRSDyY3VDiu4VHduqh7r/owmHgDu69WF5DDB
cl5wZPyvKkkJf5vdyy6+G2bJDuoOblgQe4g4vQIBac8fyBKZkmpp4BRFKAMPlrGT
BTgn+vsDNqG1sNGJCyj3Qwbo+VTbh5T5CC38HlBZ4ddCYLlV41KN0MvMMTFygAzM
6/68kluWk7XmF3KI8loRpmL0NjBEVbS/CB/MAZu6GwcR4IGebu9X9mL6zEVp9ON0
2iFn1HKcwlMulGh4zLligTZnTAh+zvUr3mTU+fjgNHP33UK8/OCxje/cx4vKiw0h
ic757x86qVfVL/fZN97i/yKZx8lQKUmWJj1nir8mOq43zYdwSa1qah/cNLeJrm2Q
zP01bHHUMo1D+kYj6kQdjRQqEXAgsbsryRH/Dq6J1o30qyIWob7HVea9De0sxteR
/VfoFyTblvKH8ql8eClCdiMQHip+1nTTP/G2kcW/mcWGn0hLKV8B8N1zR/DNSUiV
1enfWxJyI7gHKJqtIS2sQ9iE9HNxZw5SQ940++DzJDz5IW3ANqY2+z2HV02buMMd
oAqoUKdeVhEfYzNlFN58umVAxoB5o8uiI+zLxuhRDgk5lp+pwG/FAXavL1qjHrdc
ftYi7iyBvXaWzfcdT/O1BN8E7D6eOsbFUlG1CsW4ZxxWlminV6RUM5Qx1LBSIq91
yQkF28CLIorRL0nEK2x/N+GIHP0uL7gXzNPi2M+BPxTJKPU61YHpT+iWqC68iiIW
FbffLosYAU/jgjBqDsHKjiJlooyZqBiHeEUKAqKF2dY9MsWv8gFwc02gwtCnZ4YI
SztqKBXzypL9kjwV85ZOlF6pm/d6DwunucGeOE2xtzBNDfIowNpVXlxzj0PR4W6y
+95F8VxjOEvVWVOSTNJMCRDuznp+LyDQB5fD6w7C6BbvxvxRjR0KPT5tpBnz4c6i
Ho5JX1EaL10HgHdAwu1OQPx909yFQmq2uf2xHvip7y02t8WGH3l8tWQKDqgfHBOd
IpjenOHY7Nb6fnHZ2+r1ZXD6d5haxjqcCBmjqBlP3za+QEDVgdYmMMU20nt9sxV0
8113HGYc21iwHJeRWUP1+Jee0Ni4VgbIhmSamVaOHJEwX/jloV/UoXqu9LxfIOT0
N73OSfCAh9ewb2EOlMnRZ3OFRM5bOePzyCXmB7b+TVqgmVhVifWTIdQg0VGbKL4k
CmZmcBZbx4uXwakrdJZGEzuP6zzq50ful+Q/4OtzqC6+NMhu/sv82+cNe0CZW07T
XJ/JEQz/7VRQOsf9Uet/BLcF81JyV/IOPUq+qw9+thXsOGsbCiXIOgZeBbPwHvue
pNR085iZlbsVQreOqh89/OTt+f9/F4/AD6OcNXcLVKc+OFl5MvvzSSaVdrVg6Ydk
5EZHANjtW/MqhGK/2pXDSZcRjKyHpkFu+GI9iEMKeDMaqYBSJBSV0iPJb6CzM5xv
/Xrf3XOC2qhTIThUBAnO2WGqopuj9AkhpTkY1hCj7XeOo6EfYPqJMX4B/k4wlH1l
dGLX2rMrbqnwBUqn69CizYWgoEGRk72bFeT0IoZCIohawn4kD06hJDmm5FDiYZCX
XXGRpNXJXYd6ih5BS0FOLtmnFO+sXUrz8NTPs+LUipRZYHOutaw0TV8WqwbC+y41
FM8Hzj549MoUcHHdt8iKSvJYndofYHH08nRwACRUb0R1Z/sgf60hH/4ci2ckgGDj
pO8tcORzITgi/xVsbvgl/u2msZsgTM//3nAAQwqhVUBCAedJRoZZwNdSot8d8ftT
ueYJy8U6BR4d3S2DD4zGCTaHhPgxZ7e41iyA9qV4/F85x6xw7mMqWhrhg5D8P+/6
Bk31Zidvvsu61AvEcT0ea1ckMeKIEefQ5VkHgavzLiAYN0ZwrBJUz4FipzlaadnX
VSrkpI7pyMEuFyzSpPqoVNfb+Xt84J8wrV1eigH+Q26tsub6Ox9sEdqBgJl0d/rH
k1R64srC/5ZtQx1TbQVgwLcwStqlWD+162w1DeSG3uS/xKDHa7Bd8TVe8z+zlPy3
BZbW0XYl/JZ95z1/4YImkTk8wg8jOL2qLhgsWGHe9hzlfUM922n91m8dtViYrZTe
c/RFdPqJPDeKTur8ccS9qjCk91Y5yrkxXkeK20+10e3GuXs/YtUcyYaIbFo3+47w
zb7Hl2++PuORykgGa4rbZUlkphEpAy8/iPkds0D5fTHbcypEwXhexxi22lmEDvur
J8zAttxof7g2KxtpYStIpqOXnHV7J9MCGr2MR6KJNfOZdIYZf1pBqMtWlfbGeAJ0
dke56VeJKs36RwxkhEsTr7iq3mK/Mr+tyduL3joKdu+0f+o3O+WqG2cmgG/nNCmU
9we67BxZBfysOHxbqxzMauhbclMjgBhGsXJ1kQK4ZMNi2yU48M6Byph0jzOZKQ0S
7P4biedOMsHtw1EpAbEVHHkrYZuYkh/tJ74zCFv4h08eHROhvq7FKQCkD7uG4jh3
Emg2UFVGbxwmo+LDH66iPibLTfFwa/aj6AxTX3MM7e8jGigU3J3pfelfKC8u18Oh
eG0McwBXA2/gLlnCeZlo22YX8UdCJOqSghu3HlaXM3/x+hebX7fQnLEvV2ix0f4R
eQKpsy05/7IiLD9GyMiDaz/ETekSRi3pd57JPBhWyFP/PqluCv4CXlkxxc7g5sGQ
5/MvMQtd04bbCTgH4J3FTS1Xq8AY0TCQKKNF8Y/WkgQsUOctFYpOgBUFC5DPR6it
7twaLgAvD5tHNzYjm1y28K5ad45i/34N9ybgwdFk6gejIb1A3eXIaN4gnyXY7Vfj
mmRj1glJ4QSg/UxNv0he4tpTmZ3+8YR44j0e9vBdmh22jrCsoYSMh7oS0mVlbS1b
+i8fpkIZIRAhIzSruzP4+yjHgyWMPBP+0huzkX/s6uC1DucHWK05UM2uWr8wqZ1E
F1xxfCFncpOQrUyYDLerw7fIlTv635cGWFjdP8hezDMZ90nrM6Uatsl+gcrcZSRI
FpGcqPjyhtmuxuJpytHz+OKKgX/PweZuhCDGbgs/aBHcXja+jMeCrCJOr1dauu7x
czYPPaT9YE6NSVfCnwM5TRGAZ9GlhN9tvycDXyynJFLfnBXSKlNj10KZLiQ2Eg7f
cSo+OOy9msaSl1gM6cA+1E9Ynn92LloMIsOCjQZ1CHag306d8IcwBK8hDj1ogKb8
W0kFkTg9hlcjl+eFLeBIpmJUisbn8+79lHGkVKNEsRpgYn9WyrI9JdzPpWhDcJvm
zK0OaWuP0BU3vmaWGYWu5lMZkL9SiH6Fo+ZGudTSRiokHR5laIdJwTBBiEtVzsvr
zb37hCowzPoi3apQ8pz80sR/orm5DCiQnHYh8LdW8oaRILa3Og8a/y31PQVmf8sK
Jfl+/Bieahr7VJJmjQliK6j5Fp+SY2uPOoLcJGn+8WHjERtXXpa66gQnpqiHaEW7
QXcnQ/P455ea8h1ddWUb87Ru3RKXPpcKXy27zx10393kR0aBtMKUdVdcEJfT95tE
iwjYZF4peBFIc8R41J4SrM1VF+HBHyyDH9Kh1SLZSz4EMhhduppT3LivP3qLnBdG
HlN7YA8itbHyI40iSTw+If7ziZd3OnhMcTrcOIxs7z0F6+jIfBkEMn3Jue9gAPkp
k6RuO1q6pbHeG2AntJxfxfThJ81OgOuenRYyPXA/fzVyfVwT1gvFMNX5gV0p25Dv
ncbcuMY+z93PwgtnKULftaFVzT5P61SapvZqp+5VDx2DIU6wM5iSE6PQJSb5LCe5
CYs0c33HBjfPT/Gkc8j/LSUlMO4sIGY+Jby9HdxBHp2edt/icTY33ZL7+PiOWpVz
tfu1QKnFgOsId6O60MpJ4RRbTIjmT4XnY1PC0UrsumBVsQ44LlKSX0LRgmjMFdho
TKaWqL0W8jI5JTZmFaIHL4bUBsB1CLZ2XSN/ua/A/Vy0U4pBNjQVbxRe+1Z+n3oW
MpLqdiAOMioN7HOQBlmNZ8ffQnc/kzgVowGwpEMrgLsAQPIsw5dkba/sarfusn/1
gUJnqrViTUbz91yQX6YESFwWBHRzhqUBNVGkQiHYldENVdHduQdYa+u6razXhhID
0Xc2DUI5nHEwDcM8qvfPcoPWqFAZwPMTCK+aANJ1ESN7frwzNVlhV3EjpbI9a0HN
bC7p72KQGAHxsFwlo8dlf8D/mc6Lp++uylFk5F/mwdZzY0UOV5mOt9//W81JdL6p
ncW8iTX1wGmbGDKPOnxvSu3uPrDY36lpxkFlLpI5uLkTnJd5ZrlF0C/s1FSnmMdr
myFtnh/pqTCuHkkcLJ9w1/qtj8DjibK53MeP23nzm6et4EfFSmpjXMsS3XtOO6HC
KVhJUxW9ztVqMhnhjiylv5D2sMkPZnUAqQfCz4RzbMNCqUIqJoORCWrnQcUG09PZ
xG4bx3cpMwfOYU5Ds+H2UAgSCp5juQbbcvOmElvMJJeFc2TfvMM6sQz0IZ9fLCaU
hscR/MGLSQ838XwziDfbUmCnoUwT24FlzuCjkgaay/itL5xELJAlxWYoDWPEZa2h
LvJRIdqddTLgfbIeTUUEBjfxvuZZVNKnrbHv6guY2M/Qy3V4+ETDtyFzISAlPR1P
oZlyc9EYu/zR7zkO69VH09lNl6xyB+2keTjgP8IB38IWKK6ADEgFDeEGmlG5sIGR
8sKEVxS7VlXCl/ugsWdCIOZTUhL0S61p7q2k7Hro0Kw4qyDqG9hbv0N4yV590B17
YpwSbjC31BnAPXrq0pjcZljHlX2LNe/8NtNQWXew5RGHmz15N9rv+9urcLIubTfs
2P8qek8TkF8Uh46loRc19vgOp04lZR0g9ogjw+GrFxZMEaeymlf8R7TGkmuksr6p
UNOvmdKCbtTi3UZuBRsBoAFe6dYlS95aqVs8vdHn8JrFIUVmqPqY7JajoZP6NyfZ
nXZD+QqGfA5nzm6lHQGlTkriQJpDxFk8vDCtijw/XONsb0R6238iLB9+2ENX9DAR
TSoMJ0Mp0r0ErKKi6tDXvom7zkjZ7ztxOFihCsH+nFa0q8WL+lLds7p5UiXKMOy2
0+s+Vi20Uo28+Pa+LrI491SWaXGsLq3rNPgG8W8EHncz5zkYWO06A4wDKoyxrL/O
F+3DScBFNrEuVB8LgeAXKxUGviN05n80jQa94NAWgYLG9+CaY2DG6cSXZ3U0+YuP
ZVfszB/Q0JivDu361uKtVFq1V9CRyW4LtU8kFmyvs0r/slZIbTahRyPtguzu+Ay8
B/m8qkO8fyGTCy3IbnweiniQxGl02akP3AKK2j+VnR3bCBYU6VQFWaD5/Vruy9Rc
YR9tmdp3Kg3hlaPLbliCIdaKb4MPxXvGda3UHhceL+Nn4MnMQ/FpRN7ksoy5AZcM
5VcEnK7eAVA32m5wJXxJhzLbvINDiQqkhaWiNE6xS/m0uCmvZWzRAX22f36bryzk
gPr0+kOZ5oS7phSFYnLrTgbL/VxN5tiw72ckgI1aOUVqU1mzOXBR1PCqgSTTC+2l
lBIncKrFVZXb6iuKbyV0RxCd7Xwdi1a/KtIxUiDaI7iXqY76iRMHYHms2CTHgpmK
QybD+aaotvq2NFecg66GhaIkWNHEpbXjxSVQQSRFkk28WflQDTMEGpxhOoVSJ/mM
1BopedGubx3L5L3NxnCtEnqpoC8BAJZwaAzOc9TIxXagt4Yvekh7YVQvWQtz4T5M
v9yiM/crgoi64a7DhJ4I8zWJEofqxCZbK0pTl89prpn7dzXe/nwQlw+gEON/LMFu
IF6YSvMt5Kd8NAescKH3mDmXP1xRs7GOVYbzZ/nImZXXp3wAvyZwTDYhuGfl6tSN
CAD6ZR8LwHD/kP314uww7huNWF0yVOcemtHIaNXi64EHo81I6atXw2zDvp2p7osU
85uQVW5ZMJFiNcBszS1XwzIgUD5s6jHGjLEqnKzycH8BPfkrTofHFauxFefoZqZV
YLe0/7D8GR32xjXv7pnPg1FzgC8Im/XD8NPILZFDDW6I79QxnROn9BqSmBXXirCT
IANETXTRg9e+pKZxqqNRjcTlub5u9xv53zqzHwwKNSrMpJT2vNfeCPU3lHidmkLC
k8ljP1YhF19E84lV9PD3SomDOpGNLG/QYp+YWjYLzIWw5JDnMk2h27il4BKIlr0k
9rqPivwbHDGO7nL+r8WchFL4MsNUb9iObi9YHxnJtYPQcdP3qhNRTA/xf32q1HT7
ZDK4RRFwB6ZpW7k9hLGA5jWj6Q2j6XiqeWIdPWXHnvGh8NiSzjaIRLchMr9qUSZ+
Rnm+dheWGCmt61NwJefF9bjjRPfeOOB3oWN17wAM67wgu/vWOoOgwdWi9AQQkFgZ
+w207vpllh9cMpbYGkVuVi6EZLHD2YBugyBfvA4f6eVenirMlOmt+Y7Zne+5vpin
PMjOPMdQKFGG+f3Uq4qIrtgAG3ZEc7sb/Aa3l6Zkmz7YyxA94V9k+THG0/RntNpM
5W6ROToPJKYLT1N2gX6bXETN/PCa/TvHI+eyDemuixXjxKIREu2SjySr/xAfXW9i
LX7b3sujNm+HDcVqul3sa7jsYf4fqnyfJi6P8gjkIGKnE7vYzcgVgWBbOrxYqCJS
9YX1akz/2rHPhnFDF6wlQnf90gV5dtJXm3AKXKdAgB4I21OpYZxNvUhEEthTDOfK
m+t8AFsVn0R/tL5bTDdfYv1O7/XfJ9gS3jGhy1kYkZm8qxyqD347BbLpZGk89+/y
pi4uB9+CbHpKV8dkW/OqvfBoMoOUSo3xoPbnY/5ztAQtmFdVgq2kQnPMk3DfqpnY
MTz51OZQAcedf8rSW9+Yhc7xW0AY/trPaTJ1HykIvyHzFy/AbHdRqeNEVZTW0MtE
pYZELp4/CuBE788sbHj7YuR6oAUGcDVL5sg+HDN5a4ejSbGlsWzuAQbIEwjRw1PS
7tQky9+MF0spakvwV6E+Ql640YMNfUDG4EowgRyAyi2WBSMgrRmmz7TvsQ+p4MlW
elRMsvFmrcsq5a32xmjLME14+NDibTdlyBVIdh8MVzxPEtrRlAfavuXzjH6MUma1
oOgqu9qgHI+VFsaR97olsUXAPoqfIzUnm1Y/kHC0wS/feWwrmcOaYl8xM43GTFGN
2IomJeGa3j33JseNq7PqFuywDMgSYspi6iCthcnDD+VOFOBtRzUQnBEMak03FnS1
B6COquz0/cJShw6mMJgKVSouO5USpnYWZKOCFmL0AFXpGxHMQud74vv3PcCDpNo8
zmaYKGn1IrEHrlcB84x3VHj4T603b/saaxQ8zLr8B6z/1GfSjwGo9Tgq9XU3eFfH
WBV84nj8R4oSB5cyJZ6I4zsouXDtIDIGtUskowJm27l0aiEuQuJb8ymZfXRz3wXZ
iMMyf/RbiqvAY398Re2DiADSMA0K+cYKnspzvcReqIWQO6sZFwerDMpMBSQiNfLf
dAcFAozkpH6W26XnvCp3K2On2H4qShTVOsmBRhle/slg44zJQeQA3B2OfecVsfoN
W0wy69ymZBZqz13v6YDtajRY2yY4qy/+/8umFEXtTJXVklbjDxMmdn3g6/IvsAkE
XO/7rFl8g36ykJ3YZAWUlf+tAalnOtEj9UT+gyFCt0ziO/lBSKc41XJPr4reotq2
5n5+o4q/xj4AC9MRAQXOgSzIwc1ym9BDQaUws2IppgT9FFm3eOYKnKvT/kjviBZJ
FoPUpNW1wAW3oSdxJAXCT3WrjUs8FFlNcphUVescfiQ5eKDQJBlCxN6cclbBqVQh
fmKTapwVgyS89Hpgge6KRmbhPeYtLqZTufg9saPvzHL+2HrrToO5Y92JRJcDyuHF
sm1cVZ8pEiU8UN9vDizXksecNwFCEbcL2oqN6NWRol6FrOS+5EbmGmCCxCj+5/ls
qaIrSSc19gPmRZ+aDRqZ0gD1TJcukGE1qInXh7tkZR5lFt9poP0mwrwdrWyzrVXx
mU3/ycq80FQ9efenJBkawOcGmqbnq2etamVq8B01QfuTmi9NDQT9wHtJvNqqrCAG
22P+PzLRwHQqen+SpXc8qp7vIY6KHJye9HatjSAfLOvGciMhKpvl6/m48zBO+BDa
D6VKcUW5wru1EEjfOjgo+H3PGHg6znOQFUPnDu2KrruYOkENM3ukurC7Qlbk+7WG
wWnWVzDejUEnUhxux/Y1qMFSXBMLo6oxGMVuraBUinNPUT9ZQF0myZq4rtFVhXLC
WdBRLkZojV+jhzLJNOFHUZARtSP1JU62RIL/KgWbDJ6PascHkoI8fh/jS0g82LRl
rh1yLHf6bGhgwbumZ+t8r4ShO2S15nUCW+i6XwIKiY6+If1AkwLm250tb8Op5qPi
KgO89VIEmQwhmhv285zvL+SCAowlZXlOPVMGuECEwG4eB0wh48abvQdPLGUZw0FT
s47X2vA5kVsycy66VZa01N4Pzxo2whW6aec+wnI4d/iXxG/YcxgPgw+lcbljZCu3
gIOWDKSdENQIqnRBGFZjUXjIDwZbynWbfxHo6A+I606PBHaGnZzbbiUhNTfnD0ki
pHzH9VrOAiojv7FABesT4l1lgE8y3H2n41NEKoUnlLCStWHuXivWqPHzcHK7uWBt
WACjqsX2R1sxoCqrSzTKgCXO0944aL166R3/0embUoclX3Prqkgsj49av5sYSzeq
WZc/l6Al2l3KljdwgBta9CkLQXKL+myeht2SEOJau2r8dTwbjhVXtKgPfjopgRE9
8v3kpjJpzByfjrl6/42SSgo/cQXaBvlMz1hpz363SW2F68Qsek0QTlggj1Ce8ZuG
IgblMU+9tRt7eBzsk7adDqRnCO92cDTA1OejGbO1RPPFpBgfU01kk1l0HZrTgNwP
IWMMaSdo6FSUpesOs4t4ZFak5q+0OxRF91l4FAY/yanIgEIalk3mpkprMGfJxjFo
1hBrMmAOWDz3YWyV/pk2oEpdjTHQk5K3F7X4xD9GFde805Lv6kvYwiXnvFnZn0iO
29oRSnoD8R4IkcVm8G47/wroj1eTfihio6BGUmJW68EUgc4vccdvPaW7hidTTghU
HX94CGG+ocBa7/P8G1dVvtyOi7Wcyf6hfDOBk/JGOsjTQpMjYmW+87MXmNxRwKkM
BzMTpZwAP7C/YX/kYo8k5vOOuCJesiUY4I3ykEl/kVpv5uIpuAQoMDDWnQXjZsUI
P1MZ3J7iaP0acPAz5GNZipC6NJz4lc/t9tfkovoyMhO4TGX/9iM8k7pKOh2r44IX
9beNt8q+jQybO9v3Me456cOUFh6y86o47aJygduyaWBKFaDoYNqk8fycB9aubGzK
3YtZAnN3I2qu+mbfhneV71APGd0v8V1DHcgAxlQETyQ9Vm/ydSXTxOtxmlPfRaiu
dJBGL9Qr9KdQkCCyu3l8Ywuie4v6+ORp/SuskefZGvmn3MxZEJQ+0ZguiNswwzW4
mAMbpVvheNSXQSvyovyTKWPrfAc5n8zZmUzWgjw7gKYEOKKE8X+9NG6et4yCdN6f
X+5PeLjyOyAYVsDZ15mTOlETYAzJJjWlAxrqq0QDJo6emHVZOPkyQLJ5uEwqhnSO
TuQUO+JqvNFayj0YiQl3HcCQtkpVt3CGAmSr8Wt62cn6/slshbQXdSqn4gNkV/mS
qUATQGKWmiJS1ZdiRfHPHL7hehahI3RhI5dPS8J2XzAnGGmCgDFGYTpHVDH5v5Dk
Ou3h/HCcdMzydBALoaaztJvaXs0Uxht5mwBgWCelF34w4pzAuXU7k0i43udtyHPn
JfmnkM1yyHH9ZBf0ON39wR45vXC4Oo5L3iFVuScU2F0CcHZl/ufEQllVuoqFoqiJ
y5jqsLjK9JURXa9vg04lxFWUokJDlqfYqS/fWP1cT1oG49tgLtBBk7h2X58J0/fF
+Zue9U1YyjSwaYmo/b0fLASQTYJsxSjsu/3k1p/a1BYOsQSQPTwa0pFyj4YtqMwZ
Ig+4GEmW3aM3qKumedAS8Ec19aEiwZK0pkZHDFYuV5I6H+JwsQdtT2BwC7XSCTQ5
w3QRRhOpMwP6vIcyA3t5s8tFF5SePgwAxBF1zJxNWv3V/AQmAUJwxfBuDOArmSP0
UnVka1PK4HsQWnstswnb4JjMtNHO207ajAQp62QgFcXcQsYRGRvIUJ5/mcNNnKCr
TLg1atnsrUQiftsBfXAKq0Z79oJzxWMi0D7dK4EsuWP5CFWscucVPJlXIxSMdlqm
y1pag5YUAVVblGl/L4t8BzarQDxTM4j9J5vVtagYKs5zqRoOiVZ8YN/T/Tc6eQDy
3Yq0EOlidxNRIIXlO7wNO/IflKnIdy9S/W8hMEe0G+91axdVMa916rSHlPBGQp9F
d7oriCTce13SvNEYGCcuuVJnNn8ho4ppuM1HOmVmiBN+a/5y1vOUiVz52ybrjHt+
OY5UbIG25EvvG/9DnfVAXml5b8rvEBwq+9QtMEx+fSTjRDqD5KwPfCOy0hJ3pUJo
EbQlVNKJrtA8kedMeJ0OYxLcuZZTdhkcBughwteYxmBNM99BPvOnitN3bD9gINBS
6XPbdixSODVFl556cBWYhGV6ipdejzwmSm9gg58B363Vf847atSBalCGZ1OKJwbp
2DCXUMrVB4Yd5kZFpnBtNa2bj7qIwpS92aozukFaM5aZehgHe1nVqpG0fRH+j9SV
AMJP5h/ukUMmm3Wrt9NoJBR8ByMPm0VjGeGcXubP17dZEP0fLC0HPSgpqGZxYkJg
4vptjsKbcgVrc6SxHpO0dIuWCnnRMxn0ixkVSz+ETby9MIxQpE7KOtfkPlskrHyS
jc9NBjBkGRurKHzFoOTMtYa65237HWnXvxkHcGBBYxep21fWE0joxaDO1sxq5dJX
u/N0jDCLfukEzwikLtrilx1M5WCKJG48OJJEsF+84y8I148u+2HrR/z6TOO1Xh7k
djyOUefC+ODPQ9uJJGIzHj11snFzk2g1llV4SOz+W94BGB33BnRxFEIMaAijpEUQ
AeiEvpJ3hjZOx5K1pxEiT3uHTi9eqUxedXH8VKmnK9V7UeNW+ts3DCaIzYv1dwpA
6dUj8UU8ZsEsUV1jSAtVgRoWkRUiW1cmbF5i7IqF5NzJlMWxH+rVCymFut4YD3c7
aoKPNQy3/Y4fU1MUP3Vao/V8KJJMfa/eEx+14bAjQkGBqChk11YOyLPTdhDbSTNT
ivq2lkn3b1zNqoZFhx2ikfd4DrsZ2JtOj4LIRpkHH3wwe0Y4VDZKtqgULyxGzUwl
eyPzONVoD+ml/FS4d8d3xaXiERwqjc7jRH0GJGOod4b39QyahsqFT71ALr2Dp0Ae
1l2TWLG5fOod1nvt78G2LfR7IhebbrA4HIPsRxi6ilMPso/ST60wl2n5DcBdsI1I
e7+MU7v+7CVr7JjA8AjaOej5Gx573mmegSKLeDmuXTAhemsUTnl7xmnXlwW4bzGd
dizSxrLF4YaTsLNyb7fAFYVu2DmQLeerrd8k3nrCFYunq3lJnlNkKd7lAvObKFGi
9RESlq7xpUI5wt1b4iX6yfyP3zxtAARo48i94+59TwHaasCqtZElaZAxH3+1NhBS
C8rBwku6Rm70omrsjrlmRyXK+TwMLC+ar2ySWHwzpWAU8kinn/pywzopGaNndAtx
em3y7wNGLVerRsU71HDNg2FYuiI6JJ6C0uy7ksQtxTssJwFNO+/RRrGMfOVskqQ1
egwNMBX5qBJCuVGKp6c9gK6eUSuqypRkVkAC7eeH9K04ZHJ8Jh68GD8ws9i9/sOp
OyVdQ01QUrsf7GkF6UHL38GkMcbZgsLg67/GsQ+ha6I3x0itmAw7ctdInXSM8Hke
hO0jCO9cBfB0Jpy3UeJlq8Xr8Sr0W0mG6KfUrjmTpsReCT8UpvG4y15n9NrUrNgF
+OHP79cndczo05hnllKWJ/abXbdcc0aV8Ouc8dhVHT3W+b1UQLR/x9wmzhIP+iFW
kdremLe3YqNOe7Ea7DskIF/0Dc+SHiIVUXce3yfQXZpnsgwZMictcprywo6XnAG7
W+9xds7Rl9mZ7VhYhf3ayPuIKXfdbuFY+g5psFFx+mQWdMp7ZnYZNeyTh6WXQVR6
wreeEkVeVGfiJHlUaUCuxNNe96M6XavdyE5b03gUo98DNWJ7q8AWVTIWPJ2aMJEK
efLgI/9ftgTLurzjxVzvqyoWT9Ou0kMNw+4GS6C04xJIdlM6oja2M7Oor8imTc4K
zBWbOwPc7PlkswPoOwB5YKNvv7amzKixnYuKbffKr9oz0kOdL1+W9WV7X72pIy5g
PPNyMszSeWTdzvoM/6HQrojnk2qVKEE787sVqXje3QFEnipKAKyKuqMINLbdG4j8
NIRzhARJU2+ZtoZmPkPY2vqY38gX7yrjX8xvQQ9q+mKRKTJtFP16qCU1EdJs1xes
JTue2S2aAQrMcnMctuTeQ2PFfjO1We36v35v64lu0qvLZTpXPAas4Dq4ZgNUwnZD
MSePwizv9yYzTg5JTDvipDGpE5SfLSXakZn3OZ6KBdlHvnwfCUjGdgs6c0Ckp3dA
kLzCbTkiMLAyYU5/D39KGV6XPuDe3q0WF9NVmA46DbE4PzM9gPK/awiyRGJvY27H
6PvR5dsFxRS6K9njAMwTPikRfJKZI7Q0P+jNrxbuyTG8DwwaIcfryIpF6v5JpCug
yfD20rMETaoh2E1WwZYgzHU/x1VQQy2uRLyCtf80uRro9FvNxNuIxr5jHbsZ5ADz
NaVeCLwk8r1oTqqBhEh+7Tpa4ltn8W0LYnPd/CL6Y7f/12k8stzH/T3sUkJPVSXg
G5imQzjARkx0lXvz+96jwa/wuWCiIwqSKleNweBPnSWK4oan/qdmkyzUPy9Oadvd
h9zdPqPJcN8Qsqw2Z3qxV3s4KYua/EinK+jIb5X84DrpiUeFIMiit++fQpT/HwAZ
Ysqsxg0Hrn/tW3watcOUtutNn4NyMehG0/RSd1sUt+DPeVMMMmfeTf55xHFqdxb4
k7IUEvaEd8qMyXbRyEoTy85Fex8mIDTPs7k+m8/CMnMyOuK6BizJEaS7BKyMfG18
iLftyXnXGG513Dx4ErjSR1vwi1UOOpo8HtILVyhCKuhvNUWeO6M3ImFUO9hIpTcZ
2PpgUL2ukgRsgk1bh9FaYE37wRVq2vzQgTKPUW8W4Hd1kov+s6IdTfjeiC461W8t
fyfowR979cXl8JcBUPehwXydNanaP2H30AGa3uC7YsC/za+nuhAP+XtYMrRPK/Tm
eOzrTnj+DOzzOUG1Wgbwl4d7nzdD6hkKVuLBDYs1GOKUHaI4JrsVCGTBh1CP1dXn
s4gPYaKlNRjuuV916hlBi9LLemEXuks5DcexN2aS1HDhqP+t3R836uXIOWSmIEa6
c0f1TH9lLdvb8EmKd8LEOMGJ2pdynT4jfb3IdtTzVcbeCpNteEX2HLsr3rjIDUmP
68q7OpfrUWsAuSkuJy+7vq98cDP5v93IbfZg6C7vnsJke5hiq5vUKZ1GNbDXvovW
bua+0uR59u/rwfULox2/tX2d5n2MN3hdM5zVvq0oTsj9QczNaJbj/FuWoW3Kw/Il
9lBgrR8XCIW/mg993j97kqBvx2AskYVTZbG37eOAeI2+OLZFBLcUZ9W5TCszYg6i
jQ3p5/0zCdt2eqfOfD7oCPJgW7NzPzB7ibG+OcsgaJvK33EFmifieQpRuwPTamnZ
KoyW5+79ccFGofyUIpQImNqtVpHsdljExgKfo7CfY3AWHjPMeHFX+orHuSbZmNfu
zQ0xnQr6Q8ANOgXyLGbBepDoTjNVNXWEVJGdJR/LjHaqh9+sruc29tUHIfiUGST6
ByO8q/f1amc2YiljPUr8v0ibzNhV1wZsxzDJEZ6IhEILAFwysZrJVvnaUV+MF5lL
7zTqlBvMO2GS9XWpn/ONk8iLlm+rzFtgEodbUwWtqUFWPUqeTS9CbVdg4Tx8SP5v
b3PzIImdBnFxKbbM3N9JyFRSToG62PyfwuFGne5HO7ljJe47g8sQbpzBbLfu5X5I
7T5TaPkqMsK3EZ69Mytvqm3r/roThjWAU5VSq1Bn5GngG1CRahsQk8tQ55Sr7zqs
YAx0pApW4BXcXitsEkqfu4Y54xXtBIV3sAFYh6OdD7L/8m7QFj22Ka2dyE5NVEsg
6W1IQnF59BSssRVJPzGJNCR12ejxWZsFgzyNq4VvsJNCaB5+V003KnNJDYNDWzL+
wcHAAZm6k+7CixCkr8qC71FVvdI6/UwQYJfOeL088BNKnDv59T0duUWmDxfz9hBB
2vRVx+tksqtjyd9QgpS04iGaj2j7WB3aws75EXTg1+9gI0Bt6AUtP6ZOAlgQoy8r
O8+1ZWz9rbsNBNVtcqIk3aTQe2W1k7GprcoSMbfziVEb3IioPGeywdMzdlc96q4G
QjU8ibq4IelOQUVVT43p+J6nv9NxTZQOPVV/uDBfVyjd1WYG1QFCdcTfRtBRi4zK
36Lv2cxh2VA3EKybzDhWGY1EqenjLb70yv7NA+NwC3Yo0QunN8eLwsaFsxoXSCi2
AxjUS+jyjzb4xBJby/u0SqUWCHs7s6KeKlIRcZmemSN1e931CFzeMuXwFZKMucOL
mWK9tfmO3rJuIa8/27+WdjYSIyvU+d13/2DLGwdAg+aTwFbevOAFXW6PESCU5WLB
jQafw9TDI5Uv8oK06Vvaf5pCLG8EDH7UMBl8l1HYioVlLZzUOzYOEeYCvaAVxWhe
DbjE4OgbVUxDS/uT7hHNa7Z8DUCCQASwkYA+AhilN1du62Nf/cgLm2fN/DuNdWTC
NyK80KcanBJGWWGfSpzCY+qd9noGcDYdh4iyU0G4Qdl9meeKktjzVsr5G/KQxUaE
sRY2kzK00rfyqIJeVVTIYm6AIFsxr+qZ13YLaO8H22or7FSIVw0rJI70sIUanuXt
AYgpQdmc9Kqm0vEKp5/kK9UppcggipD9+RM5v0NUvEDz0guHj27/74Jh7X89uk3x
SdjZ+M5pGimlpwbEzIVBhQS9nBF3b8VkWrQKhK8xa2K/NsaPu85BYArK7xo240OG
CPOeg6bzCi5mdsX+UTxlttVeScg7sontvV2izPeF0e5t7aMHxrBVsXV9YTZrzinW
u+7ga4Nw5K89vOsssSXRnpMvnRzq3dDSLHZNaMua+Xwv+Q8KNIGBD9pCyqk3n+v9
VcLiv8+J2LqqQKTrF3PiWBlYJAjDI/D9FqR+DwK6teMyLxgkH2H3FnIJsXWIKK5D
lHP+HesxArk8EPJt9gxAP0UgRsycham8aRqVzFZefGNYvOu8whNwPtb+ytBZicIq
dlg0I+N8nG6WSKOXmi41XTx5e2TLjNOQuurVkS8xEa36hzB/PoCXVJArfvXr2gDP
aLgznSmttTwQgdZl4v+RaH8YwxKGaaofkGgWjuYw6OJKdc1E7xhlb6PN5oj0sSPd
pPld1TuEmOUpQ6pXV0DrRfTu9eIwrOtYICQ4F3ZQkyPKrT1urDz8i403SSQzs4gE
BykGTeYf2gu8a4IfQgRUWZK0espYeiT0ikOtvKXQnH3VDgfGkX2yHWI9PGCb6LTc
k3IovIRmKIZIER/OUR6PZ3Qu0hC4/QjcqPg9v6DvUwHsqGRybhupdUozNm6uhYrR
lMA5w0tRemmZ0XssLDwcqIz+NQJacAbxz4UC8lY0ZUH+208mVcfRYu/nykmndleW
qLJJyvt8rTbaE7SpFd9PwRGzltwxeixBg6AQRW82+xt7d/CRHXzvya8kcGrsZJ/h
OeyRPv0kDXgjKpyWOg9ndwA0Y9Mq1kMRC1O/vN26uGTJxMyFVrn1xd8ytqIOYqS5
pjR9Cj7bjZC1Q4y6qqpql/ePfBJbPsOZHklS+VS/KA3vPTWeSVp0paf8Y89dIzn2
OMS0hKNB10mwIV6MYzvZUR0Rq9zit2kym9knZJm0bFwAt7wmQNXcmIpMUzZsMUGS
8K7MKzYeOeemJ0xrbfiGTo6AErJ9PYwJvbc2IzUnUuWftPfWyjNE2H0P6rQtfMFL
/kDxwBEAK9kCS/5NQ2xUmkP1IwtLLawJlyACX/ETf+IWkxpzu9JORhiYZuEj05LZ
3YvC0zxUMtTfYj4y8BQqkPsMpBXmsCngbxH3x4CRpxC1i2kvvSIcaHKfq5bYvqMi
bkp2gLEuy3c9Z1eK6WdjVo4bjItJ4+4uzvLwCzuyl4DGnbe0kC1mmzDi2G5PZ2ot
UWuRVJ8/gtK/Z9m+/E3kPXHNRfJc44LYf1M7rmTwgjAAnB/PVr7Ubr6ZXgWDN3H8
JYSveiNdM++nCdtvW2Cbk9EkapGZza/XsvBbGKa1RAggksBNC7ACBLeTagdxcTdk
AEf88Ugz8AATrL/whcr2DBaSddFAZPx+3X0+YMpY7RSCaNFkHAHjVi1mjmmUjKkq
vGy+AHhm1jomkg+5QCu4nQez0vuyLk6oMfLioS3EdWM/cLdUTYQIxGsc9dvTSPVf
M2yhrp3/i3/IW6BYQdZGg+VWk8d4IFE620XHRbqZ2Ufr/HtqE4FogKzGPKWyvGBs
NZkK1oNMWAMPqLMWyGhDS/uBci0pgg+YMvSDGI4yEH82fBWNmJ+w/flTpFk1TZt2
NiAwUsX7IhW8kv8Jkt1GVlZevyUV2Lk329PHp8s+OKkwqxiqfI6MCcaLhKaYao3e
UlcBNkI5mpybAk2B6DCTe16+Ciz+jNja3E/ctn6Ag+oPog5xhsBsdz0NgrhDQDLb
FmD90YQp9E8keX0HOqNaqjiqD3l24JRoY3OMHJQXG8u5iljsmGno94XFxTamFYv5
wVdV7fkgXcAXK8KKcLc9zkTJVTvTWKKC3RIdnspf8drJft9+ZSFq5bEt6M69ued8
UNEDYhZNGCkMqc62wSn9+zz8QHmDDUWHKQ7VDXHBhyt47ExNtdnm/TzmfFWDNnmZ
+aLlWlR8Phq6SCcEHV8Kdylwqhzo5fv2dxEy3bkDgQpHu51pxqYTUQrS08gwKkfJ
yLL8XVhfl9dFiDEjpUEKZaGWH8Oa2nhJ2JIE2YTxE8+7GZbp/5k8Cd6d2ghXjXTf
RQdRxhnPW2JN4ycv7aEbnYAnYGDm2fyQ2Wcy5vXSMp8itcVgK4j0alsI6qwEmB8Y
n0XeCcRKgTHbnwlFHTP5escShGYxfPqm0VuKsUAwBa+KdrL/w+qlvLhGq2b4ORZC
tBAx5YXuMwk0qDw2CmX6hTsQWgLerc3W2v6P4c+dehpZy5yt/Leoq/81udakn5ZR
4QvWZxESmK4fbiBlNDdhpYhWWrU6O8B7ZIrXDYpHQXLOnWNLBrzEhx99OqHFdY8u
LfYALh9bWSXjoSKsEO/Mr3sVMxyBF7MfIX/4TPBQDCbGU/Svj2I8pQFLodm3D+kt
qniB6MAioqykKdONGr82Q4QIihZPwOiMjyTPRni6dhTmk7CiRioII5YDs45vi7l8
POiIoeugPzlqAyl70aRNmKD9nrf7EAHayHOR0mWAvPC0NsGhEj6dyXfmv+VebYgO
YomjPY+qW6XxvPRMRibJBxZqWp5PC7AyjLNxjlJy7NybsOB7rlmbK9inwJ9kuxlf
vlC6dwY2ZAlEXki3KbglzrZ7LiBZDyG61iEqT2cziv9JLipZQHAAkR7YQn2TZvto
zA2Dw4XyXIPJDq58K0E7rAHal2I1iEmjOfK7EYkOzWD/EGZbEibgEAzG9MnR09gA
MpiCJlqKeOVRFEhtWhS035Cd0V2k3R5YYkFyiaoKfpik7dZxOZ6SqD+QeCnvcfhU
5mNdWEDlkyjoX8zjYu32r1GsVQXEdRx+7Ja0TNLgH3Wea7Wg4ntx2nNo7wU5vTHj
DsYuQSevhvxlSKGBLtv9saLhBZrij86Av5DcKOEjbTKGBezxkPRYoD3imkQjYiYP
A2IlFxolje7V2X6oOF5UGyDQGFV/IfV3cVQ+UBpY71JoRYY3keWnuSOoQIliWmyc
bRcGDUu76SZjM4XxSEHMnzTvXNU6y+YxKP8R/vm7VhAHS0qGz8IqtNrQR3XWIjAT
7T/b9uicSt5g/GT2rtnjEWgbBSuLXDs/6L4GzxW5FZtdNT0ROb9v5xjAItw2x26V
YBl5SkDU77MTZq85GZBoGubTguu/0phuh3EJoUd0chJCmJ0CrZsgkDm7j1lKwSWM
Wnjueuf4Ygp60rR32eey1BkyLP2y9pgE9DlPvEaKYTZMfB+bN9zmvP8GIgstigFC
IfgRMC9AwwQys05IjolPPYPXfuQ+7OFxORP/89CPZgiQW3cIAOYtOZHx8S2LArzE
0wsJbr6VQpzWYSOJOCJRA7uYw1zfGrRaYmN2z9YooLstHDMpUUZe/E0BvL1p9BB4
iaozx32+CBMw1r5FXu0GNHTsi7BtAsqaNYguJqnuCyOubJtZMdDMQ8mGCKTmdR5g
rDDUqxJgMnqB4KhlrV+VgRna386tyj568ZzeDdwFQlo0TKbcKLGA4BSc98yP52cf
g8MU5JqY8ZWHiDGE4i6k8sMK0k1CdeJ2JmdUwj6lUwz2MiSEcl1Z2eKPn1iDBSUc
x+N+nzoLSoAAv1B53P5LvoZzi8VXHPOLNNbfSUIAlmRR2iLlKmswhXv9qEtHF3UH
BkWHiKJ7h8B9/sYh+SBNkjNMEOyith/nzxGralZ5KvXrnCjQLjJBq6+KVCYafRm6
FuBwqwHz77d1PgF2TeQoIL7SOt+q4Zt7kGPBX82qVuZhGwVThQ8cHL5Ih02bvJ6C
JocDjx3lhLZfsalJ1DRox88H6O7NwZf6djOOjhoP/Ehln0WcUE31yYkkBd6MCrOy
4oazSUtgJcgFPN4fz2jJJYCsdvRV2r3WdaLWY6e/DmNAs2azB1cAVCBXb7czC/4E
VkcARNABdbappxHWIpkYb3pVm+YPJkms/bU8dwCSzbiYJrccxhgmRrpxUy76dPse
8VA6LKOBp/qPrAyc0kzBb0qAXQmvFzeN4ADIjCL/EHHk7Y8Aw//nTb0HxIfHU9EN
M1m0+kbAnlggOu2Vau4kp+5M54xhiJzFma3D5qVgu32f9d9hudBMO9wM8esc9HH9
IYJ3bZ66i7iSgZD2LIs/RzWZAlX7eq+qjtI4hlHPjs1Y76zHjvN4aYfa/6OQCzPI
8OEA69WLbw1+rAfagGZolV65fpEf4YCin4kDhVnwxH7ayrJlsz/6C8bBSuX/3/gc
YGIE2PxzVfGF4178vBtNG8c0aOqcp0Viz+Ep+n8NBOW/2abKI+hPGHolJDiIph6H
i7EcBNN6SZhaQdtBJBQ6pW0WW1jcCPbuFQgkrwS1gDjDU1J0oyfFOpJxcIM2hv+u
eGVAO859GWYDYoQj3dJF/otZ/fcxMuUhv07uzn/9djY/uCJUeSmRe3rfCV0/rUBW
4YrQqAh2z8qWzFPn8BB+/8FvcMG6sp2pH5kmtRBpxb9O9RCV0ISHj75F4x3DVHly
rFla4yAnLpc2R5MjE8hCfrOW0ro8plMafF+bLjMbL5wQI5lMyOa38nCyn+YALh1+
fUcLLZS6Rlj5v30380iV3lf2rFqKycvTscEcnUC8Pm9UOn8lverDYm2RK41ROg3M
7mdSRAAwNIGYyqe/vgbNwfeIyfaYVg5KQsXlQ3birVIPLa6UMLOgU9oR6wjVYtW9
W+9HrBgR2d7nYmis4El2yb2b0gQ67cNrtlXwt6O1/TedJMq9cSbyBlaevble0Ndh
zFdssBgzJ//8DYCOB0YlESGQ7Ts34vNo1OqBhgQGvbBxKrUlDFoPyqWIfIRgG9Rj
eypid9cOxDmjR4/+i+3aAf2ndi8n/B3XfvW2xJdANUj8ZccWUMhf6E4vQ611gjDu
3fXj0mr13GDmo7d8heXg/F2aUAF+5OuE0X8J/HVZIQbF729buX4xxyEXDBXSBxMt
D4QQRF2oysdJJBZ+VaEO5jGjrjW9x9Mqoy7P62tc+s62meom/vI/bI0ogjo1m2cD
Y0DBTVCz0WYWcqihCeDm+UqGu+LhgNTbuLVu0c697s62vNmQFCW2f/vl87WYlkTk
XzM6dWtT+VrpvpX3vrzWm3i92Q44V9bw0MfPBMa6vBEOx+K85pWfAYb5uDy48UKP
KfTNwLLyJXfbFG7TnJxhAdMdprNXzTIEmPehPUagAjlgjcTRjEygCu2YPM12kx2l
Gr85MHGm+OcyuiWCs72mPVsIgptZlMDHRONmySYQxYuXN5Mt4R0romjdb7MS4ylk
uBZKt4akUjiJ33Hq4B8NZuHd2BOL7ZZ7+9dBmwuKYyHJsP6EPiXmnMBFQjcIrpve
Dn789upEYbYCwvXrTVSXKz6b6orgFu+oPYM9cA+qZ5yYjBeZgjObsKLba/uc3x6Y
F8dR/34ma6K4nAoU6s101b0FL7D29qEndcCjRlT/DjGI9docO/emAltSoXPFjZGS
PR1XjD743BN3QJHm37SNKUe3kUBzULDWxIOmOnkuRe7u56xUiNNQep0VqDJDLeAE
6lkrF4Y7s1RSX/SGM7Tn8OvPkJxk6DNWKwRL034JAK1mWKb4/pvG/jhQ3iamQlSO
GPVZ901fyDnLb2kUtfhmZ4v5AXGezXEHDKyqVMzB9X/CkYzDe0KERRgakSO8Ze3z
UyPXOtSVw5TTnbERCFYQIIN3BgE9iOTu6T/wGNtN6kv3iIO4XH+gxG50Hyu4Hl9L
cZcCPPq4xgbkSl2IMLCAa7fshuhv8CzZ3J+Mh/LTZ4RANKmjbZcP3115pt2/3HPX
WkOrEvQvi2gBaU85+JxjYUoLDX/sGaUYOx9/sEph5USQkTT9MaH1StN6rACMwd25
LOdqo7mn2Q3nh5S/IlaWSp2Kq5zUOtB+rpxhfGBRzb/l4TvK0FxC63Wg3AwaKqV7
yVoi1lBQfouKw/zSfoKOoPNnYpTcGzE52TXyQUSbpYTAn7WR0E9fNnKI8ufc/3A/
8NMw0kCIgTQTFQ/05eWnsxPQ2NSSZ+iOXDk5FFtLIbJ6Y3Ye1ATMsgbWDPXwb8Ey
sYC+sUrl+eH1mlMrXa3iLtBYdm16lx2AcvlRZZi2qaWsw3WHinrUJfnnSD9nA+Tj
CwyB2MRRzdlgf3L9tUy24yGfNuDDtRXIHzFAYSy9TSSi9RJOwmN3QHMjKoK3GjTs
/tV4LL8jV2MBXyPYMEuL5os8mKcOYK80E1UtNwKiGOrvHEiXSYUYw7mITxRvNl4M
xTIQCH9m9P5L0BofkcKt3C9MDM9w/WzZ7w5ZN6lCB7BH+N6UlipLCnOPwTw1QUmx
UOCUyfpN7MuB3dp6Bbq2qBk6RR1rJcNQy/Nm4OdbQqPqegBc3NZAcSnnD3eHSOgy
zdnePnEZSe6os9Cmt6DsH3QZyBRx2ucjno0fPmGBaqlFfet7dkdMmO3smvoQCbzi
vKPWowWz5+QhnbsiG+3iym/wGP7y7DjEukPVOMZDIZ4PAzEkixnv0EdaCVpAeHYx
WTstgbRrp0yIf7eh4vFrFjaTLuqzGVhS1MrQttdZJhW+kwZJhUIF/I7F0RLVhMs1
3xo60WT3x2ECfVCpSFLkPAu+NZgYzzwxy5QC2mAcgBQSbZE6hyjLTKYW8qrEKGWC
fwUMgeDrXH94bP1XGaFH7R7O8b2mgwkxAmshAI6F9ICM0GT0F2cPq4XujIuUSgKN
Ufc/8sjc3Yi7uQsmHeomNq5710OMImWZtQXXNw+a2vYENvFxVNZY0SV5Eni7TLRy
IXSQsEX1IDYGAHWzANDPh/NaAGUiGTzlIGUozttVqHc5aLZV1R9OcDBITsCaAZ9Q
OSeG6E6uozNXqIct1kLWAYvZCwwmr0/zH2vLDXq2cVDUc8H6JVuEOHrUlMgRZ4CO
D01eY8YcQKql0NuHqPNdFCav1MjxN+QvbVnBwzrH6ElzDmmZxh7/PnfDvn+iW1hN
LdjgApW6utSMnJ5G4y2LEqcF8jemTUoNdj6Yz88c2BjIFGolfGfhMRNPakOsfm4e
rNUUos0n9xpnG5dQBHINPeNAaNwyRCaUaQt0C+9Xyy6G7A4bvG5Mu4pkhRRids0G
uJiZXLzxTxOrIfHyDUJyVlWdHiVhKYz6hdcpMI5pxiHVHZOZdof1fBWZ4iZfI+Dr
d4bDGzhPB8iQeyW/zon8ehyt8Z0IzMRanCr8j2rBhscwAfq0B3q2gEQKT3iWrfhD
gZLSGScKSBUPUOBLqcBXWApVL9TW8Bky3nvkBxY+mg1clrHMLFA86WV1lixDfkIN
R1s0RugTLtZsFC42hM+wXWbAEVm7Eayej/9uYJGzTzElgt1cTsn1YOO1JML4hmsb
n6cjLmwvf268ZSfIJzK0F6WkeHBx/NkHT1waydg6vj+vGpI/iiSZ3LxZ2bkmmYnX
e9B61HPKgvMnSeRpm3o+e4A1sH+czGjaJLK153BwEXfz6Qt0oqzUYdRnOSUeJGOn
7pvAvZKKDM3FfJssDgoB1uUHwD43KZq0sauVxjo8NrCLoOeqWz9eBwm+tVPYNsSe
Jpsssjt4+LBxqJpbembsFqnfxhoWmciOmZSuZxKHmHt6XEzk/4fcb0ELZJ+076bk
OcWRiFYJWUwgCDK1v4WmHUlVj3x16dYv1nzTkjwSzxJ/MU5J1pNAsSk/C2JRb/iY
yPwD1a5oZJ9u18jhwaon+EUPDSZ4OCI+/cUwBLqCK9WJsWoO3jKYR6oTbNdOI9BZ
A9mF3U9jrNT43jZWvng76n1YwEdmcMKHO4NBubmoL57s/3W3sVWUq6aYfd0KaOAY
+0Y1nPXqnFkJXX6EcFBq3P2iZ/Co9TXrXc8yIpq6w4dwlUVm3tdZwjL0momqO6el
4iDJAI4+fP4JTl6MTx6ojnSUEWfXtXKmUItyA8nqoMEax3EbzqMmz8G/Gr5jPhPi
naH6AdgKzR4tQa80UT2LBDEB1If13ubwh1aH1nTxqlcptGdcmcDoSNrvxRvTIcw7
9jPO6r6bZ9rC/ZfDfq5ax12I/SlJyRFIAyY3TDsB2JOyAp/vIDfDmq/cdtKU5L+U
K4V93x/KiLx8/LI2eKvVWgqonNTr71jAvmO0LufIlHljLQv7LPOb4OMBPXnLDgB2
Z705aDHrP3MUVCEjyCi5iFeQo1cSu86GHZpiDQZdP4jNqp/FKfxH3e2sor996qA1
h2vBLTmH9td6GUmtZCweTROPE3ZUlEhSOyxBcBWIQFT+3wWlVJK0MUgptMxIiOc+
O+SHqRTX2gMrc2/yIM6G1csE1Vrr53WNa9Jue/xXY1kBdXUArcSFnbjohv0/UMtc
UseleCP9UzucGHSM+wxIQUDycqTCRMcmHvNamfLOSSoBQ4knCmYgF+Hwm4Gnye2k
gF0YoShZ9MNoGCCW7vyeizTdf5Vnn0uLUV40FcIfvdWEvYgvQTZF4sK95o2bqkW+
+kTzwrssZ8ndNspe5opLOGkThTZFSIYYB04RhhZeqHHsza8KOrE7mnU5UxroE0zT
v0HHHqtSgu8HUjAuGiS19IZLEPaQPz+n++QLdGyq1zDIV8xbKSDwa398fStnVp78
H4xuA9t5WxdhWWJKDo/tXFMpfPIkb4Vc2voLRlilecN1ZHaky7TYCslOp7lw5jTW
VfxNKe5HK30H7Da3I7W5ZU8hOz3h1v9A5YAyBIwMmMUek6CFb7Oez04uxiNIoKem
nclsJEhemO3x9GOhSdrC4HPJS6k+kjJXlguxoxRphu/+4wAZ1nsPg7sBhhsWADpl
UppgxQNcJBciuvJ3GyiDcvNkQ99IjksNUk3z8gDMs1+IIaMK17UHMB7wDEfrWYDM
PE0WadrSpxEh2FDeZUV+mTCl7Sjls9hskrvCF4W0ZTaf72mkIhDcu2oGXz6XLJ5E
7d5f+9zh+A+j58TzvZiNxCg3VBLWSuEGaKtfT/LC/qP+VWrk8w4ggp0lgREM1CRB
yrOdurvGVhwQjJ3CNbzP1GIoSf6ecBEP5NSlbz+Rj1vPkTmJCSllcyipqXR3vUKM
CRXt4vb7vWUYmERZ4/jkUfKYtxGwaA+0ffuL59AcMTLTSY7FBpp4hMNN8AKHNvwV
euJGeJa7eeUi6uTzZI8hXgpKLt+tfqKONAuXv3WpuEdB03MU90gFjvBF3MHIbCVf
/0kUmfc+1kz5AIaKCWI37qAs9K0HKqdjfrluu7Up8/TIX72Eu/0rckLEewMlLc71
gxiRs5HDqxHC4hzXK2vjMJLRfxzNA8SesPW9GoA2cqCNYQlko2+elvMM49fyK+OL
32kBKiFHHzEI29vb0ZnXCHfYja2OoBEmk688te2jvRsgyl6Xp8YfwZ/OPxIRnhsg
mCn8GL6LsHU4GdW5/11FvQG8qotBYJPdh/u5Vzy55kAgaZmeZjgClDNHHrzL3Thl
zA/MfZci5Wl90Ah/NLdr/VWjwKANIN4O/9s8cA9xG76wXT5uTh1Ge3jUPMWligB5
IHF4VBYsf9SouG1e1hrg9VI2/Jlx0g/y32Fuwxw7s1e0QhXzF3mCs2pn2/kfY9Cv
4aG6FYruPytxzY6B1F6cRgZ3P2Z09pMXGoqKmbtm3/bbxMqShtM8GKi6H8A4JCwk
S1gn2JcGrHT92RtJAehtQZ+8d3FooAXJFaQgsIJLfyQcGkWXgza2SwNnMbyVwJ36
LCWtpLnv2uwC/hRZm7yuX2GOAEhKzNUCPtCyPYdRi2dKuDAYeZeIEt5D4QuykNjg
Jwnjs9GbOxKd8oeP9ssz3a9IEs2tgyC5dBME9optkhYyVH809KjsDNsyaw+Nf0Gg
FozRmARfWb7EhRphShzB+xa0cgt8KtcE71QSpfz9A5JOcB90mM9hAqR0OwAqsxK4
BzbtEmK6tEaMsjRSd8u3usFPTcLQa02GDWol+3f3gshfMHxbZSCJ+PP0ZzuSuOEG
wnH08qO0V3eZZe5Hj6nuXUv04kD4IS4PM0zsTdT1V2rJtONQtwvFT4JjZMkaIt/P
QJLohMLQT/w9/64vjQ5AVQKKhuoZhwtw/SbSMBoz7qO/IWJvvMouTqVb6xloCJUN
KKOO05euV3WiTMjw/V9yYcpTvKpvy4wq5zsLjKNxi/TpBY29IS/TZiV5MK3b9hBk
PcxfUaII6Vr0+ajI6MAgwR5B8z/OrkLmBpNRUrGr8ELeH0fIUq1F+sUau2/Mu/LP
Wzs9h8BjfT0tEGV/bgSD+9ZRCVKj9CiX1WhBLa+UZK/WKukJjAN2V4BYXOW8vX+c
Vca9YFy9kq7IexaCpv2uz0hvVHYNC0kW6J1w/VJev13gDVG4Ig43PuqljDsgg8TI
1R9+IrOXdc13b7mjk8AtXh00YOqZ/9jVptwucpupDYpfZVXAOninNiTo/DgXBygs
U4pPFnoxPE0xxRrvtMUc9E2RwaR5nxPHNbGMIGJ4pMIeorZAso6c18t4Iwqx5iBD
q7hOiGYKPH0xFWiCBi/Xitm8I018wCikUiF/hvhI2B6GPBohv13cxjrcSKWXKAI5
hXrOdZvC8X75ow9nABPxBwBCfiht/KgIj5WQoQCNcHEkCc7P7BvlOfVzkq40UzTk
A5UFHWOXHPk+eR+8DPacxIhzAFJea+ZaXPXBh2P2/BAOrgKqWsk6ZuRePmndeFbX
y+S1nMawIIdpTjaoXvVxxRwCZUZfhgWoxU0AozqdzMh9d4E4dFeIilSroCPvS6x2
Yqzyj45q7HC1ywrJiaMfg2oEzXeNDko0fibk/QdeaVyivxYN1ELOU9o/H0vXwwTl
kvK7imTZASl57+lnnM5C9Nw/umuznsP1Kb0Hbr4bXqBE/3TkSyEy75AcWfMJHC0W
dKQloLKEPM1aAEr1QUsBf15Oz1gL796PaJYRTIO9h0PAD1HZD92u/3Mp6EG+doZc
hUvXi4oVUq8ZwWTEyO0y6IoEGcEEeNmFh3dYBf+iEY7UGyqAYxUfEpeU44OBffzc
/udYAUQUFaIYPNJNPOXL/1GGkrlrzEf5O1HHKfjP7gN4SWMHhIY8uAha19Ruy6ZG
SEPhptvOmi0tse/6vAVjD9ofH8WqA/2EDPpeu4mhT1/wq2K83l+B8ZnIj+gMLDgr
3XNQo7zjvLEUNQuLDySBJ4e6pXBBTE6NqZHEJbcvdwU8Ax5K1JhAH7zews9o6W0S
gR+w1Q28brA7uc1f5eHu4BviGYnz3JRMazz/ycKsp6vQi62JNqcbhuIaN8kymXIi
y8KsEO6yNDD+7Kt0ypR8DhfK+lfK17jkqU537ljqhdyEE55NKrs1BuD+mEi3WYCP
Ykqf73DgV59tHZVaOhdUZStVnYGskcxGbi2Y++P9Kn1R+r6J0ESz6502CN9nKxmz
VElQvvv1FXwcrhNBf8zi1Cx8R4OZOil9le4eqEjxbzWyUqBtf/HTEoKYP/cv3fIP
cC+T9JDySanYGrHdHhLMXiaBeY3lbIEEZe7DBpAV7DTsWXrf1yekP+d6v+4NN1nb
9k9TFuc/z+etevH3sC88aSsLRsiEgZa+vvbqDMuS4TRKCvL/yJ5fHT6wFr9XX48Q
A9Gf9ki4CKtPCJpWreIVzM2gIW6enyStYK8KDIdwUtbdZbECNe/UozOV0xGcF6ZD
ccNe4WqJHMO2Oh/etiUtqbwSSHtd1dhN/Al/4QPBq0jZQlivuw7hsb1uVV4gGk7E
i5v0DBJeiacVmRWelzJw4HGRK6s049qYNDL4iyrjyrEgbsw215xe8qtEbT8AVoDp
5FMkrMrl/SMAiQIVruz2X45D0bnheS2c2rFlZseFS24h1Qxp5CGj5ylvhYnVVW8g
DsLm1+haoatugxFgvIl9J6/fMkhiEKzF8v9nNmteqFaZ93z4vubju58l1INv8f/D
s8XImWi0I1vi512WlA3Ao9ielHVxt/ra8IKIzQ3+OhpS2aRhf7HsB4Ks03Im6dCn
x7AgxBI1yM6hvgv1oERrbUSWH3f1UjwN8r140cNFHeKpdiGvNLhukcOg2qGghAMW
HRfs1m6Poez9xWzXHs8Oy4pIBrpKh63W3mM1L/us3p+lMYuyayfDW6FzNL/P+tSl
BuVsI/8eV8HzL8BOOSkBSTy3Cl3BHtI4JUKei+VBzF6mdaC3V6/H0V5wECz4sUen
vNYMuxvvBS39ijvYvNHMLF11U415JA5cybIAUKcBS6s2lotS6KQ/rSVMv5RrDciJ
dc+ucvO82D2HmwZgd94isd8j0Gz56s0FTfMsMa6zynlFUT8LbDgvottGUCOnZPGn
uEL4qswzmz8we+Jle7+io4m6VLYz9CP56tEgH78NWWhIukGrLDWnkDYzuLeb9pe/
4w219lZIg8eYoB2aRgT/hsKJ1/t51ErGwCaAtEJkj+damBpD1M6apCZNYPG61rgw
9w6O0j/9Ghw+BokPt1BxkddRnf5OmBhpk9HmFtGp50hFq9aFarIZowYJPvSj7FmD
zryHJCknMMlQsCDFlxuD9Jff6H/LFhzFohST27qU3pdRF2dJ3PsE3PwhiAlEFCkH
bTrbw00b29AdC1ZIME6eXqC2tYhn+8fIhKzFEgkkvwz0+1n6vyhHDZc8VrBILag+
yQzcOY01c/5IPrBJ/Ie6ifMmHNc7ouNM3qzGrDpaS2R+lF5qaOeQHEeZErXqElU/
+RFim5cetwv4WMpYLnlc07pcWvs14lzCmq+Frd+r2jABppzNdqCaN6p8HvHHNrhO
SWPCM08wFFuwPp0RW9RSYjMySYdmRDIuDFK7ipDqPWJgnwGUSXrFWTY995S0JCfc
vQDxwN78x3GTOifNpEOIYR8Bym2JYmptBRajMT2sKYBV0T56/zy3jF1j9zq0TMcG
HHKY9ThOFgiGd9o3Pq9jMzhDCNm2K2d3lVudJ/voVtgVZtAfvhbaGfF1I/w1tKb5
vGiqkVGtTwjERbUnj+7/TuGgH7ja2KvAXp4lD2QX29nVIwypng0+nPNyAN0bG6wa
nyVTit6zGWjapq5Tqh3t2rXsUJWamNj38Jk5GrxQ9x3FQp/Wm6ykzktQyMZx5Q+0
0KHVTvTEA8c0xHiAaShyp5boHXMWR8lBS540uSry8V1RdNl69CNTYbotCYtpCLFt
NUk3OfYHQT9bmI/fM9qn1INR5Lv4I4YO5t2w5JIf7FhaKAB6pFvBFQFb+zklTQWI
rZBVCAPHRGpLFcn/glAsSHBgfBR5goQpLSBsOGDe7U9/IlRWOC3X+7TJZz2AapKM
QoPj77dUAG5FBrstw9Vy0fjmJFnOAHG3QTElDqVTzacaFlb4sa1tht+WkJqDPUv2
1mEqgo+Iykdqbdw+R5VIkVsIkElaR0IFT86NErFTXVYh5LTWOZ6RUaryeLay6/4C
R3Q4jhFwWcp8pKOngAlnQzKI2nJ1Z3FJu2opp2Z2SUwOT+hL5/aN4rsP4Mp1Hawn
gIFsLcRQDb07BJUfK+cg4vE8s837VPs5SXynRTwmuX9Nr24FvfJz1RsMsR63b6zc
k6yuy7WGEFkAfvwcGawOyWhU1gLVwh30UMw3TBqJJL2ihg6vp0SOH0o3ADLXX4uu
kGnl1Kr3yHS59ckuTeKv0iYSQ1eHGU3OwepZPltacltxdcLToSHFrBl8pfXxGnZ6
ZOP2sXm4yTKnLoT6lqvVIBCaPtsCdAYQFBJlGDiQUX87Irz1Gof0x4DmXZSB7JEt
RED+1Mh7NKXE90MU3ZJcwWDDM6EIO6XywbgkYOH5O5wD0GVwRmUMwTc0MA63Nddj
uofrRU7pfQHsVGObEY77pFuz5E78bfhZvbgyEB/PD7AQtqGk16zB3o3BNwomgd/m
luVVhpptgwHd3znTjvJ3Rxrzzb5Ra/2Ua02+c7vQ2X6Z4Eu++RDESW9DDbId7ZQ1
/saGfJSWL7iD/iqPgwFUXv/TcuMD986Fu5Kd28EmtxWepUOdB7Zjn6XJuI+pI5zW
2UtlwbMFUBp1XLrddk21wCfECxlaGx3Az0gT4oNgKa37Vyt25h5CVtXK54XqkYgZ
Rv9I+Wm7JTenATDWCcEcPiyfcupqMp3mmdndh4Ilg0JbGYUxNBEdLsPtUxug/e6A
789epu36YcY53IYyVwlWcM9yfqv0e0/JNpkz5Bxnxs/KcJNuw8BFi6qDVhax0/2J
QDrDoGy5O0xSU8IFm+AMPYWYe8EXhQ5ncilS0V8ozhIQ50QJmCKxGqW8oCTghD74
Yfew0DRackzL9dcUEqiUqYEzqtpgec6F1POEQGFPFfeRaLPWYkXF68uydcPLUn3p
ZVEksPmyd0+aOu1h/BPifiRReEOtiFhDRB5U53/w/W1+qkDv1t2+sbbF4w7Y1IXK
Z0Ph4ru3IMnSLh20KKinNeQ6jI37ocJ9mfYLWUKeDxHbIkz4y+5oi4AQpSNkACxd
8X15piOMscCuiX/Ee0ekhIj9RPcKv0N+HCHVZhSR7FFFnmtHcN7e3OlrEsWbS1na
TeR3l24boAiSHSXwj1O6+yAT1y8NoHvbWeBGAqDckIXYvcReJH6HLnqgs2uAJf7j
kGPEE6cfW0P7B3IRML6K+hEg1TA9RPd7hHZTcf4SHiNtxG5gvNcKu9Aa6yNuVRwJ
q14a4CeDbguOaplzN9EKiKgpH9C1McqFmrMlPTGz5QKRocO9gMDR2JDqJSLjq9Lx
k3xmVEPtChh1qPZt49xQr6W/nWqSH/sW8DkhtCbTMMunROKtOfMPYihJUur8WKd+
VbkcNDr5mFGz8tYH4JN3v5APmlRiWTaLoVR/463VdfNSpS+u+8Uk15blXSzgGoix
UPB4C657HR/fJMgyHdzDarKNwnRotj1HLFxv+4no5u+5FXrp0sWDrDL2xV7L0iOO
J9F5VjREYEpzVz4ydXoTWAP8u6D84WHV9uRQqmsO5FcHaHW5xqDadk7NyaqUwfcb
H+b5+gODEE++m4FO3yn2XDittP3APSh2aR3bIHxLADAVzfBZgJkHif6NZF1fzL/i
BRIOzx5jrNXMk4e8diOtxF27x5UTdcS304gUsQmjc0zePWE/PAF4oK80lzCWpoy4
G7VC58RE3AOoJhrolAm1G2O8hAKCAL2RFEVxbgQGj+/KyqwHueQCUWD73trkQwlb
XtsEsbvI2ASzIuVBmtdhvTNscgYQgygmfoTlK8EddF538yWAE6dKEWsoRP25JcaJ
+vSdKRf0Um4kYveF/hFnxQX93OT95L7YnPyGcEkEBM2QKsN2JaOquVggjR3Jf2VN
tsJqnT+9kINl6cDd1Wv6K6MEfIAGegtN6FuxZSZXFndcB4QGgty4Na0F869y3z/J
8nna0midNRgcjv1CpF3bPPlOkvQGsYmhgcCROLK1iKF9OJfc/cMPaTIkQlwOftl2
yk0syAdhNPLUd0oxd2WxRcrE8YUUXVYvhCHX9uCTyh261Opr+hYwvL/6Y96XZp7G
sUot0PePtPSSOPvtO17PH216R2rKe8/o/QfvuR0PWxLF2tYGyjAWaDQdsRlHEnxu
3AYSOD2rgbOksUc3PsnhZqy5le49AFIEGIS8OQiGoOyAwmtxHuA3aSiJLvxjH09P
s94eAqjYCuaSw8z8u34YlzxhhEtNcUFfqpsuaOnlCvMChAj8MO5Fv0GKvCe8AmD1
E6vB3KqE3msliZft+eNhHIaCrZpSdb/U4O9uh+0cWBxJq2a7RvNpQdyHQiIv9nYB
B9QRLrbIjpT2eG3+wOB6hryKM1vFHPXvLHR+24m02FWCS96Nz3Bb59bLrmeRQjt3
PpELcxAmxPPDHCWsXJRNQ3adKnrgMEURFHvGSGjL+OkNVvYECNH6dsAUlVDu2LiR
g7CUJjJEi46tvYcviqnwqFumVBIzJOfQZ9rmLGV2fpqOoNHWSKh+JKcB52NCJqGE
AULaqj0LVhDIYdVCLyxXBEms5KHiv6cWMO8o2zuSwZ53GH7r3g6mXtoKe3f2BLnl
ps4lBM+wsDxMj5zavShcfOM8E9LLjyBSsJlmlKhPql+NyaEk7+dDgp5yxswWwyAv
6OzwPG2EVEtG2G1PG0gR+T6q3WOZGL1XamNuSqvW0HpJo3/5fSjYk9eDRny9I2vE
vn9hhOj5VtfCJ+O9ueZWcb1JeB3VvD1aVPphsry9xFbM1laJ4+PMKuKcCVofJSp8
Nm9zvpkDgP+T3eiR8P3DJdUfjLH0yhr3kxxqzQOd9SdntFgu9fy2wZR/h94+AFsb
9BIpQ7VgxSararsVIlyhyQI1fpMAWriqjC5FsdQ+QRcCpuYs/VD+8G7+XWJ+n6eY
2v9qsFkkIsFv8h1zLhJJZbmkKJAmPLOaT8tTr5htrdXf1G3KnaPfK3cF51e6OFYn
M7REKKgHNHeLQzeFbK61I3BGq3eBaz0iFZmINIfzN/3/X/qqQZ55lDIk/w6fLFly
PvkYo7sCt2qUNACyDj6sa2ZQaw2mPqUXNB6cnRQt5VX545Vm+qJgfda+pStOmWAZ
MT/JaO89BDl2Hplv62F4oPCfHX7iE56akcW/8GGMxUxx14tq5vwm5r/iBlsAh3CR
OTB6nHR8tM82HluVrCTBvRoqESe/9RGHUw/+OEXTHcSD91JmDtrltSVcNWyMD+Bf
o3ZwKphEv3hLK9wnhSMk093FmrKtMWMunY/qWMYCpoZk/V0MvgqPA14XGoWEole6
uxPZYyvhnUXTD68fbg/ITR8a2OcRYKm+77Ou/oek4k2ELKvKhwmFKAvfWD83q0uG
JIFAXcbNLR52E6N6UIpx0Irhqu15G5QCgz6SKud8KqsXjrMqzSOCFmbCMqbp5eiW
Xh0YwKNpnUFlHFS08M55XQusB6EY74NmPNSDi25g60nqc8I2dmUhiom3YQQO1EaW
IAWSyKfiAVmVSRrU4jejuYnF/YF1F0CCZg9qO4Vrf8EdxEfgJspovvNTNABHGF4+
sb0YfY91WKthgF2aue/3SHAFmIlsQvAp02+EfL+pYOczB+vM3r1lteQw/9pkC/6N
fPTXUjkFUYlZr9DBJcGSt62lJ1L/ist7il+A+rwT/erX8Priqxh6xPDT3SE/npX0
5fv6fjt08Duvl05BohL47HpHWgjznZ53kROS2syfLVHm4oOc/3j2+4pNuvxEQa7F
vYDLsLUpXsQazoo74odRzirnBnjP8xBSnqJQVN5EuGyiXLbS8VvMGBQ9DgPNMiiN
CmRsiU5FmMwwCi0odTeGdHjUJGGhErJDYazPULW+d9SHlcUYXPgbR6atagqPCiqW
A9BKxvk2Ux73tbZbs5DzoGz0am+VhSD1jyOGUAJF64+DvIzhViahh8JgftngWZyB
oKK5xQBr+6aNjOkeGcCO/J3LZhLhrCBE309uej0H17TMoOiBZnlgc5EQ2k3qd0pR
2vHMKkbZjpsf8uDeKoKB0P2Z0z77zU63GGsyI0cVP5fosKw9f7noCu6/T4v7+Uqu
491QDdTXuZl00+gq4KT46VliyilHVPRJriVOTStsd8Fi+Oj/jfP9gK1ujtPLXC+h
eKRU9Cetzerz96i2vFYzk0XY1/nolYYuRqvhWe0MwbyLiXNS9tPzWnmBQiwB3YmM
YZnO+H7GXTt85Fm9uhw+N9maJPZ0ejRRs2MHZZ/LIiavGjbCRQ8uVFv4rMJV6JYd
St1SlF9GRMHNLZT7Rg6EyMWTQM7kv+cE7eElURXbvvkMNLW5yxPd8nfZBu74qZHy
sZalKsVBwLX/MWWElggoanmb0SucOVUOpuPnqAKVyMBdReOHtVd8NHhap9VS75pR
iAeHmIyiZxKDOryhqaj9VqRT2SMbut5yI3wwAAzw2Kh58x+dj0iibra1+BPDQLDa
qby2kTeE+4iulhBk936sxgB3rzgvLL6TjN0dUY0VytrrS1YDUUY1Tou2Zp707fQv
d0N1zIhwUsf3vUXrPa+JGMP2QUJ0uC+RrJ6awX0DfnMP19eJFh+Yn2PDZeWdp8rf
zVIYrj8x2FHIIs+z3fX4rTPMEUnm+XCdWgodlTlZlcBMPHbEhWpi37AYvyJv1lff
YunIXBGFLyGV+g1CtS1pMxyG3dgD6nY21iySwDAheWpp+mYatDB8MQxJ+WUlNmtG
elMZ5Ze9GYlGcMwzQuhBy+jgKLjA7IvoMtlNJmjge5tRbkqFGMi6+1I8/FGJzo37
a23EpV8KFFL6I0cuJ6qBF/6Zcis4C2lrrXg4IRpqihGspvxdujdfBRy9IUHTzNll
HNI2wnYKIgC5RyNYxzNEsLv7L9HzoVPRJ98q1Ze5XLlBFHlneMQ5AYh2dVyur6iS
hG4yYKs9FxvVlLKoN/6uY/PjFZLFL7BtDqgOBGVgyiTOklBpC8mufly1G2dlaugp
yD++uvyffLlJfxGhbhMyXbUruccNmhLYd2DxRUEbNmR5eVb8ktgtQlXIsB4Cm3tp
OAeNI3c5H0yyWjqYInetFvXQ26fHyQvxLCrhIIHrvKMEDBex0ylFqzSW/aLvWNp5
kL208/sZzLLnmW5ja4trPdnqZPW1BRL8OMED/RI/ZdkfxEvZxnMd5Br/IFSdvyvz
BABn9Xbzk1XXcIhMSjCwWMxpJ8GXrfdg5qw7Geu/cgkZqEqMyFFzxlHajToTVt0K
fxJGEniDeckzzt8NjQdorgGoLkg9qe9Qn85XYeTHShn8hhxnShDf3aruRqf4AQla
mkAr+nmuEJlJrZXYgImLzerYGQEAyL0IFrFhHeQ1N4N/712mN19vBO2sq9ZrfkDz
dLcShARZiz2E+NGckfgpEswFFREVXEixxDm1NwtdqmEAZkJSnc/bPoWe0PdhwWfp
MnTwj+ljyHDGJknDX9+3+/ILUeKspgtikmGaJ0q7fMsfc0QnI2Q3WIpSArX/H7zx
M0or9BkudK6vzGN7EzmEGTmDmvyi5HVmdqkBxjrq5hKXHZmygewW001mckpZSUws
tX3niAf6kL5/3vIxyID6As0WN4nk93yqvyQ0vSJWmCI2lCKvZMP9CjUE/6TBZZe/
C8mOjitzBkBQX2QUkY/BMPmPYyGprXPZu5Du8wfO38T3FLPGKTudwXAZ6SekTh9Z
sW4Ct85tnAhVVAoq0CnAcSoWR+RdUI3oN54lFNgoJkvZQmIJeuCP2cda2Hmgoe0/
rdfMP535MA7ZPiiyT5m3/uqZXt6uVho+JAMp56NiwpQmBqgEX18EvtoET3HEvfF4
GUffAvRg191pXdauucsQ8c97LZbg/l2i63ZnYkZ5/GCdA9Ot7xlzBku4pBQp3JnN
+IfoDiKjCoAfA6AOjIKNXMfT5EnxZj+L3VFv6Zuu9EpOHwERQtgyL3QGNXjFnwjC
SzpjUHVf2wiDtkinZ7M06QREqA/TIB99H2+NmW85Z1nXQ7C//TMsMKUPh/eRLiol
mt/n3ebPy7t2z1pq/dASyWUPHXvu6eqw7ARWkZfKYkmbZDOQpdi9J6Y9Ba7iM8rW
ionvUWVvp7QF3HSe21Vy0CSSS25dlDofykUG8EhqModaklPCDgjZZBr6n3xKQaGo
rtqM1U3QpbKGBI0Q2w8cIiOSSLHcjuMJfPB3ptmik1rl75rzjhTbnfyMJhRe8gLD
y9sfcrAZ3tgvqaEw82jaIy4ceZ9CIvqWMi6pLl+XXkBJ//bQGP3hEBb3Hp8LD8k7
Zu70pRkeY8DY8B140wyLnrtZqjt1y1TN9Pdorz9VphxXzaJYj9ylrEC3LjrGWTlF
lqWtLPYVVC/jkHEkOpzmd6CKUYEwassviwYCG25UJb03Y3bOD9frMFsGt9HE/3+8
PTPOk0PsZWt1bHqwskT0JDkq88/cXTAY+MMojS6RvE1FJ7RouCC2MYYw9fVWKB2U
tP+KalXwzwshSXwtrf4ZgNEKZh3dhTVlTgumipU/q6SNIx/OAcwRT9bcmt+jVaTC
YeopeAjCH6gqMxZnOSDXoFCf6n0ny6F/QSrZeXzT+t4Q7WLNJrqfYSH+hGbRlW+s
xbXhosU1wl9bxKIQS9U3IKPBQdwL4Zu3KWNjDOU9uSnb6SlZgfr3pCuPIHJvsaPU
okDUoU0z89jZhNyfPbgUiP5mfsAU1ymNQvYpqYzkK2zJM3O6sWZGuEPPoRuAH2gL
6dgH8DEZWwQSywAO2FwJgrtyHoyOjAgN20UGy1ZC42Fg80hg+L1h5bckwdyWW66n
auPZ78ObL/YaL7wXXwt3H8Xr/A8qpSonnV80jGXR7B15PrBcoHrowy6qusS8o0+M
krvtsZDAJQaZOfW14O/L9an+N0ojvJ1PU+BxjKB+aiisOGlcCh2udRl167FH4xpm
c4smW9zE+Jzz3PhR4OLk0w6ZqE5SZ7LUJV2CUCTNIBPFySLAbuXNN+fGWxn5Dhq6
uF/DTnYS7vm82hs0lmaMQ/hE3nCruSUV3Onn/WSzEMUIUFx2R7QkmFydhExpBLTM
QohXN/co7bKxkDY63ewPuCseU4N/m++drfSPGibLOEzRmRfnRQJIK//ezNAdVIZA
vqLvqyaCsLSaU8HPtbwYLSZtxK785ez2fpxZV7l2Y5aoOn62xMUX7d1ccXYU/yUO
PFgkTPRPrePDYMJAVHK9W+icvhAO1ag1mXQ0cBj+5B9M+qGF5+ZMtzyGwZ+wjxrz
opa/JohZIGzPl4fH9MZUq748GGd4BpCYBDHZMlO/u2NDLxacqxsJQWwCKNcyZJJ+
WoE8ou2guXVIuAcllULaaf2wOWBV0b0Xsijos/Nst9p51a2Hndgj4vPYUP9eUaC/
oGUqsBNFtd3Pe4KJupDYtRNpZiH1oaOBWaFPRLHxJVXnknSgq9uvlQLxUI57+iWa
CXEsS/ydjMC9fETuhGmsZVzCp2cgdkWNThhJoBdDzPlRhJcjQwYW8nN/fBFxW6Kr
1+Aiq8kMv1Fefb8xb3jT+jW8zO+Eh12YRs4YFADFwcFvXwnTOM6q51PIDLbpcH/v
lqf0WxuvAw/e/wCCS7lZ990yM+c/3yDxgJpPHE5fPF5qmvUJGa70rj8t0vfHc68n
dAzm3U3lQvm7lbaVBquxqi88b6FO8YSYNKL93erILZxz8AWgs5WzZvkU4KGQgYJo
5OxNcWhUsZWhO4WVG+APy0OOczJMlMuJ76h4O+vtftDTL1AT+qbK1EgG0geGidOG
H+iLd6E7t9N1Mo4qfswge7EtAUhFKhr0yNn1sjZeeemGwg/ndX8xzxLmtaeb7TcE
Hw06tTYivh+nhDHozeAZpCOi2GQFuqpDZReCfuF16tEpdeQvMJdWb9+SUXUOBtvk
9NnbbHE82j1Qh0wsm2izfkEbeEZZDCx+K4iaN+yBVyiUrJtbycbH9OReLfSg3Vnr
be+3x18zYN0v+LbvL9KYVaxUcjkDwA7H9tNCHTknmAuR5yWduo8xJHCn2h3yIcxb
f+XA8IkOITxDD3iXsjqZf4BOQG1tSTFNWkzQzDzdYBc1kus/MovBEXLgFbNLz+ol
fZUOX8eyMruV7WNXn84S2LJBHQyA8SecOI2oB6sIJ3kO5q0Igu09tIzkEYBgitzS
TxjGC4gwkm0UmFkteoMDft14Rk7XpMHyEvIalpMA52BGmO51g+XdNUgcXL3p8kum
quIlaU/y3wYveV9aPAhhv3PkHrqQ08SptgATvDVNtk7t0jAH6lB0c+q9Vc0Od5r8
2DAOOJ3RlR6OPvKhMZCD9I/LTD1sf5XXEQz6HCffqPiGpB7P3etLF6HQGetszWjU
EYIb+kdPUtRjZFZMjXH8bcbZBFf/LrTiQwUCpC++WzJvchRy09a3/RMcvww7+Jn3
OH9C7Ym6Pm8L1FF5if8MKdhrYNTcN7CrMpKfqtTJHL6cStMIMX9zw9I8c9x7jhHH
yGdOkZqhIvG9XN+REKqWea2yoYQ+fkR1/x/2ybksn+GNvgigeTpDhbNx/Gwagmpu
2THiheJ1xUqexgBGWtcuthYKRGJDwHgQJMTnl4dTeh/rm4xhsM7T6lvdL7/1KN2N
pMQOoF4So9IrZgIDEtdAUaD9BgAM7lpAAxKMrUwUb1uV72wK2lgbcMmAYIdr/UID
xGViCMoTl7SmJXrL1CHiK2dfS1D6lth0Gwx6yecObc8pCBjrS+JoSJvXLCjjt2uQ
IVC+YcDdRjEKmon3KwJsvaUThN6NeQ3V0Zj79lffUUmCIKlC2MpkBdzQrb12wYAL
jSIXGV8gLeVgoUxLGb5HYUAzDZy1YLvhEWEAOB8T0fBxmVAmS2OLeqZfYLHsG0Ck
kUvx6O48SO6ia86gn5bexEF6zYiboY/VL3gqwmK50pVA44Bf5IHez5UmdvqYWq9h
LvVKH6YOM7lP1sBt5diW1Vk0VSO67Xnkl18C6OMSO1xEiafyIRQB36srFKBqMJJA
rtioNreK3bMOZ1t6CO9xfO8QINHIRP3OP539+DX/IsRxIDSUOyxzzOqtLueahbWy
dbO1VMRUqFnxFyfB4MV3hwJJ+vSeUkAOMuYiULjOExUyFODjOTEF/q001f0ERISR
nQ/RGlWNauikxGGSW+N3VmdXUVefekz55NHI1FYG0Hkzwl4EggGd/jyN3sG1ZWsB
/ucQjIsIfZb+VLUQ/k1frOKouixc1W2ge5cWfh2DPgpqC94q2MZZ1aRRn7eCCvOK
9sPXdZFwpSBqb6Xq0FUGsK52KgBi+q36BJhi57NQGhlupiJZSTxW3f/RA3GoSz/N
h4uUNGDZRVQlaxwBEoV76HhELzXnPy/3OOPeaf9tK8LGPJhgcIKxcfC/522qGJDV
hYTB443BkV/P0zSo8eEddaQZN7NG2T/xi2GnRpPsBzIZdAUhRL4SpcAzsSKcK2IB
PcMNwDPL0bdeHMaHGv2PTavH79RsPSIenSyKqGp23FwVgv4FBAmlRv5iQFDu5q6x
dDCG61JUqgSpKT20kEdZcpPjmANLliRy7pjcA5rAgNyYmKj7nej8T4mU8vgxbNrK
dt+dc/M9fJ6Efh7dk9U087w9+cE/AVcMKlJ1YlEvaW4DsjsIqpeper2gDKL6mBn1
VvbD4AVOnxVJ0oMeyqpqmAmXndZArJzp/7IvMn7r1ZRtFwYQMAMHwiKZpnhIBUff
PsAEl5EkZ9mghYkszQVBqcqPnduvrb/Y0pcamwftfKxTsJIO56P5HpcTB/FJXklR
c6QcsLTMTESCvDJhYgoXMOR9/Mq3aYv1p77crKwR9Mh/Y66R5u5ekkrCR0ggPszm
6YYcPtZ86X2+7VMgQN7G6+j7lgtTloJq50i1GkuIYDx0ZinTZlBg0MW+uwp0kI3V
Byq8BlS5t4OmcZ8D3eKt5E3G4h6KHWK6NOfddfWRLyloGQlvkqncebW6IOHa7Fzg
LK4MxIFBRu6urwfiP2Og+/1Q1OaCDcUqCYzRUYU5Xu/EQnaHFSTiBNcB4z1zIG/h
e/YsgFcnjcVOw2GvvNgTaEC+HfKNODjZDpNvHoSyQB7e7dIcsDHnagjqICHmx2nD
ng/I2PwYDuWDf4KbbkrjxWM2lN2Rwi6F/7Vib+L6CQC2B0sGO9vaTFbi/rPdqXOa
hCRuwVNtic9X2ok1BXBzpT1x8mk2Vldy/NNa5OAAUtnVz81zbunJW8C3x0JdrzxV
6UnOMlkmeo00wCMmPpDq+ckDe2DCYP/JDTUjVPR+psdUEMo/ng2d7dqlsMWdu4Es
0dqgv/CY8uEUSewGg4jLkJKXbUP5t3cuapYZx3rdIqVowLTlniuoCNNi9W7vB31G
uWzb7nZWDL1gehs+MUVtiN7cHd4ZuOHqgpeHAtQxMitTMJC9xYcwapV5wWym+Yb0
7Q0XBXaW8u2vkXwYUrv/j0308SeZpJBxVTdKTuviFEPowtVyVdj1/GWdAOK0a3RN
ml7kLxo2PiGr1gEPVH+lGoqVY1PYL2jeQBr3oRQSqdRcg3IUFBmI8NlUSXVvQfWp
U8wKTcalVeBhava0omtDlZzeMLLja/KiLthIqtMbX4x06LWaRUMLcoYc6eBoV4F/
P0AuFpHStavQuMNFiJS10TewfKFAJL56u30pqAA2Lz2wEW44yG0bHrUY6B0JLGLq
h91kbStyjmOWGLZygPHvIGTQpaCu/d/cqAMQzB+R7HApsjh0LOqPQZz0qmId/94v
5kpIOeRs88ffq0YlRnpDp03e9ZL59U1MAFNp+k9/b4MlBgBLGQvq9ErtANxRgck0
gd7Kb0DL4aIgLgI2qJ4fGjbbHLuB/fi3eqJ+ab+J+eUZezi8JGuEdABAJXo7wxwz
smsOy/8zrPhNOZV+bfCc3Hihm+0KqV/V2x0Us+G/WexNVmR+rowR5y8HpYY9VHWA
/wHQHl3i+eTXGLAwS/6RFKUagmPYrB+oq4p72rw3H7xgyibVXSyZZY9GN0R0lOjK
xFcCSe8XQazSaJiOlpsSaTc8Ou5/3MXSxjzrcZYhN00iGdUiwtuf+AXg2/LhEPVw
LBDBsppcoR3JWukZnw+/X9laVB+98yGgh79+2zmGpRZvnznzbJbjxJAKBBaQw3r0
xXF26CbLgHF+/dMe8K8+e0i3EZ4lo48sGsTSvc+kELRz8YPYv2NIJrASMdsq+vzV
laH6G/eke7VArKGqPkrMijGYsbDmGKtisKgllr9pz42UNKWSrQj+BYhPjDSlMxgs
P9q4EJWa/XznvNWF6OS9VrXBd4jjd3cHdl6fYKlkQVtFEwG1D67l/LewcsvdOHxB
OsAXw00ZxcXYwn9eePgkvjgW6fazFmcym2JV/UfxZu40ZuciQmn1G7dVgFjKoise
0XjRNU5LpzO0ed3Ej3UhHuDK2cjFz8Sn6CDonaHmd2zrAwk8nr1EwCPC9GdZnZeD
2oHyCGf4ygyZKXgPohk6mxM2fh6e2WWl90UnBojjjPrFFpfP2zekud7W4zKvAzUX
ik9IEORmuPY6QCfxEBGHJiqWvOuLNpFcJyb26FEWg4ZVIxQOXMiiQhBqvIshLfOJ
gmAvk00onCF4RNJk6MH3DO7jrMBTGFTDEBzsH4Q7g9+0bG2s9KvKdV2XSRN6CjK2
P//Ton8StkvxCoNenH2Gqt5VMo13PC9llYX0LjcwgOEy5eHwMsL2+mHxBekrR7tH
JNLr2Rz6Z6MkThc+z7p4AAcDKsFsQN+SN5JnlIk9bug3u2oirhNptiLn167wVGg/
e0zx5sfPGMOM0qiYAt0kMQtkMF0qx/PZ7936NoUT6pnyiyh0FWZSzF3l70K/Nagh
VR3rrv1zqwbQVVxFf6c3YHG6wGrKH0qQgceSOxu/c5zquL12DObFQsu8hBGtlZfi
85FSvInI37b3wfrEQx3AacoUUnBe0cU2UqXY18Tv486+vJgl1RZXwyqG4d8Yc8KU
Fks2q8pDC/udsG0SgCCCxh4l/8zE/QJ7MuuQ7GgRbHZHE2QX9/YfMZPL9day3E9W
vUrR3jGbQGL5ORQG0EP4kQEHxdvipYZ9xnFvceqoG1xDxNRQevmbNxNgcxWSe2A7
GR7hB8K10WC8t69wA4+w+71AoKHJJAjC3xebK432p0SsUQ/58isXrJk5sXfO9Ljk
aGNz0F29Of21x9vrE/qCUmjOucoG6g3U0a6hglf2z9qJ8bqODh2ODIbAZfwpBOyH
D+gw/XyGvAg4BvycryrAOyrkqAQdE9PRdDqHjkIG4vLNvADHnpDqQ8DUXEo6KMAr
uY3DqcCAscoSH2VtyihqhouG+thKIHXSV12DP/uuVwSua3z3OLan7rudFv8OVVZ1
7bL2qyEgboyCoHL2na6FMQfVF0pAyKcrCQw/h6CyhJNI9yyYwiEF91ktAicx4Q+q
/RSrcFsEKOVlG3m/IT5MOFcka+aHobuxW56ykvVjAb09i0izcIVUNBzvsYLFNvlc
hhR6tinp+6fJfG3FgbwkVTO0VZr3QEud/NMwGPZFZpvoKfEQM0Ceom8z0rhl22qW
cAFTXm2xT4zt/RQxb5mnpUDuteashpm2obmEsrNPXBw6dQwLgpD5FSKQu+IQ0nCa
9VDgtrseO2ADPU2A09M02ljEzpW1EagzUVZcxN+In0cINo2HZlzGHGuIIni9IppI
ms0ar7Fc3VHP5YgExLUsYQxvwKwTVinKYBTeZo7wWFPPWJId/CYbuHmTkCYrAsnV
Q10MEYagSG2BOyWApX40xPdPAf7q3jOEV+Mbx783Af7gsra7Nymtv2tbTpGrEY8C
Vjoi07TulQ03GmCKEsICXQm3cV5fiYSXLt1Fg+TdckM4IhI1Fj7JEfWW5fNnmmtt
y6wibQovWuMyED9oo0MWt1ZCg7BUeIaN4AAaqcnqwOtbY4pmghvjt1sf0FcleT1j
icVQjKQByF9346k8i+TmglS+XdZBTbVjDoM9SfE4MibespaLbsiAIWfzLzfHM3VH
z/d60xEqDaMUZoAcWDm/GOvBni3jEH+6rTlGEKFGi8Ln72MOwvylh5d9teEmYgNO
VV1LLtsy1pZDN0kwNP+V45pm3CK09ygZ+x5xmYeHRcI4ZY8uOsLeRPzDP17Nz6j8
KLW9lRqTAaHT02qfPYz/hDSpuBlBpzWt0YosEr6iCiaBPW74cRoEiHKMcGPVgZoa
FD6tUSlpSn/Zd0gFlUOPxdZ09oaXFxsOA7FieKl20+1RsRI6kHjLtIk/sn9pfnxP
adbCBTDQaCWEct3hN7qGxMqIynCeGC8JhdjpbIw/q+tTC+B9V3DzB9kJErNHkcgU
j25yopNntiqw9iTmpKqptkmVPDi6yb6j1qP3MKMIwUi2V/dzTrN1hV9tBJztX3pE
u0RILcMVtk0z7z1DmrpPxKF7YGPFux+XBC7VCP5oSiJJP599o5gVyU/4oTgHm7YF
XXa7dmT8cFgDNzpwclPpuzWZIgAcM3CLTk6eJy3g+j1GhFzlfV80nsYlWNwBeTzD
WkTbmFB6fFDQQmv8GyFzSQXm3i/fTRKQ4P6UAtX/tknYDjKVctpA5hTLFro3Z8ad
HKobRww/sU06BUb520fBqrsm/QSuwxtGU+Loh1xHVPjAusp/J7QFiDGOtqDjLvaB
Y2SPiUb8Vr2SVg7ZKGRp55eJetucs2hx4piQJZ2usADFZwBsmC4SCg2WUPpNMUUq
hEQ7MypSPy/gYLtdreqpzSRi55Vd8vAmiDA5RKnUox/4gOZk94J00QnV4LjEWgoG
iZHzcCN0E3/EuKg2bFNffXYCB9UwmrK3PvmKtoJdBx0tGwkBHtGqlUcGaFk55dE/
dyXo3+oB9+OHoslLoX07yxkyoLEsSVHvyD/0CEL2gcQqFO7dDjFW7zyvz7YgDXZc
hJJX2l5kE91SZkOnkw6XR7SNz8N7TvHWuuoKJNX+lZGmpCkkfyBvHIytr1nLRPzk
coAFra2zrIxZKXO7zdD+1gCNL/KRYRt9CJ6xDAkVPOIBxit1rxjNwMYesXDdBLyC
9R1LP8sy2tNBEfqld0jVUKBqaKOnEiNF8trNsxUCJSNnuS8UsO9dAQzRjtJMyEFD
8wWTg7I/vFCLiQhCwYpPDsB3J1N/Gk0lqn3hByhHQmzN0Ij7K9vH1YL6ky75Nr6d
CZfkX52mB62Q+4nzQpkSdeZ7alqD/Nz00wtQE4GYHwGwluq7Nit2hiznFKg/9j/i
L8CLOaFAikWvU9NLH8AkRvbkmYkEV+o7y7m7W40T8fHwTlODnuJv6FX0WG6tSpPm
Dfrxsahe6Wc16I+BoT2zFX2H6hUMFopfI1kU1inokJvP//wZXCQY3gMBwegv7RrM
mpKmXRiFBmwzGTQKmn0Yq6SZnk94jetmnIo8TD7j3rpb4OqJQ5jwyFpyOHm7Kghz
6FNffjKelwLQr4j8Jugv6OU7lr1bJCzY4asX+unOpgOo26ThXZfPJ51KvnYT4Qjw
NyiNzwghK2TCR63yjQlXOtKBxWiS4i+HDOhuXAiiM04tIUcoWA81gDbO6t50nPe+
V68zWBdg8SnJaAUwjg3YSeHRKD+ImeYENJ5WbK3uqcSkTOj1HyRXQsVczv1SoKRs
diHCkD40T/Nc7GQRFIg98sz98J6g4DlxSZO1Py+RC5sv1eBBGbjVZYEfTFWipJeB
Ai/n8U+21UQLXVhFF5xcMGh4kc8I70/f244pfMLhmHHdIltkKQhrcmfP1v74ik8d
UPxelBbMw5UNyxnotwccmZHUSAyPE77FyEizT1rLClhX3n6Yw93CdMTV2uhMMcgW
OyRRTu5vMqnqpyRvGrDtdMt6DF4ptZqHl+0DWWpwFvulyzj3jym+/MJU7n+4EZAV
NFcqItrLO8WSU4e5Nta18Fh9739/oTQYwZFmVplYh2QZTi/QeCP/AVIGVsw2WdJf
eBWs/EyU3+fU9bbcYEY8fuzIzR7BHZm0oMTvzSqyrN4IxIZSaKHu11hBQ5QRY7LJ
WiDfXlylqNmgmWAAqF5iPHeKQGM+tbEpe2dOqkYc2G21gVxB1pOpdZIzj9FGRDhT
XlZZK5IHOHBVPd7xHCV02d7rBhh3pdvq7SQA96/ksvadIccZxcV1qUjQ1OiHUfVE
C95cMg6iKx4J/EfRdz98YH8fN1iIMVx+yX+M1rqtNsgCQD1kXkTgiqQnYduBufmB
QUH+g8QfaYVSHx7X4K0cirIX1KHLJgwU6GgHSCp7MCGFWzUCXlNHedUIpfRe3sIV
HNYQLit123Nu41ASvw+YNUPV33VVp6WVfUzblIeqYQnyM2WcrAHBsf2ENLJ8Om39
f5Zjhyravm7+7AUol18Tp6NxXK3YtJQWpDB7e4NEuTP2Wv0qbPtoAFOLwaT7s4hT
1gKF70OTC99FKCXD4zOTTbjRhkpjwemwPc3h6S7C2HS2cK/6OIs2qyYI5Wt9iMW2
Z+Z05v86MpMOec2EkofPrrYTgZwEmecTq8x9NlpjoxXKW9xoJw8M+8mNn4Ht+2iG
OuvKvt+riicM6ZTW8XgqJ4wq6JNqpZGwya4DzaQjeIgJUUQp/AW2pAK6Z2WRpu/J
nVvSUNXhj5zTurRILxdJNLskDbnpk6ui5B7FaTVhr999UY63DALoUTLzJI35Bcpq
gjyT1eUYvmWS/Lvw6ygxT6DcHLagyd08NAIuuCZTupThQ07NBrN1pJtNFUJUYrs6
/xc9ttVOS8q+Z2ASFt0SA8yyL/3D3Gs8FL168TQuMfpPEyRjclhgDzpp/Y0irMPq
m0PneNQKbSIJNF7d6ErUAw1gRihm2LCtLQELemfzmm+2/cFioyMDHHhv88FzWPIX
SBFVnwMWn7YdEFk1uF6nZXeD2vZBtEqcRgzmYlPL8/CduvEuGERQ6dOwu/JhCphl
2LKfjGO2K9Mbs2uQzX/HUMj2ePM+YvfvWg4U4H1G6UtGAS3ZT9uEl3f9qj73MQnX
fQ6fmC3cUei+PPpY64Jimg1Dsi3K4jnEkc+5xAsrlzsWn/TW0MbjBgt5JNxUVY+k
RKN82dRNSdYSGNL7idLPCYgVT1VEcQZnQ9FdXaZ2qDyRdsQmEUK4BIDLJ3BxnVLT
DT2YL5xfBRsKgHOZ2vEgB6qJdjFPMOgwSJyWwlNc9kD1/WjMd6hAMPQe1tmcxr+y
8OfxNxLsF4ldOmwm6qQiat29/sQwuFH2P7Lzw5h7F5k3WmPzRGHQfy+xKkqkmLyg
mkV/czg8rGgYx+dIXbwR9wAuNjdQehsLqxmJBtb1BF62vpxS8rQkMohjMj36bonN
1JlRme2excmto66DNC0oVdrEwuDa14rjiJxZz49vkaO8o2B6J1rxOgD7UhY+A7ha
orI6K3Tgw+9V+xE5g0JPWwRrRJuJn8KE91tA1CH/jCacCtn07zKIPrI7CrZgfkt2
S4rN+mLXbZG/b2vlZzP16BefuS24n5TQo1D38/UW35dKeW3ewgfjs+RblwupWq+T
349Ym/QSmRgnHvdAG9UMBQWTGJ7FT0gDBbIveU5PabWkhae73uyBnSc0a3R3r3Qi
x1b+jhZL7SXT/bYocQIIsMIIHIsAuk/w17wTXYxL1TPsqgYq85SnWTvYRdr8JeVW
oSpzTZlEILgf/kimFcRyLIupctkgLBNJrfcgiv+icJYLJj34WN7lBDukUq4jlh8g
q8SGuHviOdMAMSQNGQWjflq0VAI+hcV39eZFATfZr0+Wk5rGZZwg24WwiYKo5d0U
SVk+yT/FIh9LTUPKp5cBibJWYpm9mXrPLFgVobiyePg4dXxvZvU88+yPmEWmZead
MvvCMMpqr2eGmLV6B86JoReD+PC7E/VKVwhFBbLnas6iW95j2/ngUPW5mcAqCZut
xjjLVjVSShicC8/RUfxCvJTTDsYOAwQ2gEOdwz5+KvXKdI65JmYXXnB470fNxsgI
kVZI+vQPihalR0xU+1gaGJjrTVw5NbLo7VAcaMOCX2YukBXJZ2yES6vkmw9nFshK
uSOK0zbo9lMxUR3OH2FknwrLDv//6ZggiV7fLy2qOIrcxg2tJoOH4ZW6E5veusDG
ZJoTrUrweu7nso0G7FHQvJ6sqUKl3fTRDAmYWpMEXX9CPw9e7mfKNJ6tSWnLX4aL
LKoW+4heiYWYPrXUv11Gdx97N9N48lyD2wwpqhsk3UcfO01A5bVrxcWkJbvHh8Y0
pWp5rkyHw91QUCzMLo/tN6xKp3DITe8/jO1A5NDF4ew3hdbWOlY/RXNtaql7LDYs
CZfr4CLL5FYnSKxh7ywPhTeYVvAxP+U2t7IG3qzDLL3R0S4jP940gtf1g087ik9d
AcsHJTlke+d0BN4Ue08vWvieiMiJdyGv3VD63CyHl1kJqx+mxtVht0omdC+Vk1Oc
zswcIK2RBHWe1whoishzIsvjKoWzzRu3up5sTQHkfulXp6/teTZnnvzX+/7n+4h4
56Z665j47i/HSXDqxNBxsPp2uyYH8PzF4+AqsctSMqIl2q+Btpp8mwHCzPrWnzq+
cQMVIFgO1sSjxQUPytoSngAryUGs1HHAdLGSsxJ34iE+GGpyGpHeHzNSiPGDeAGb
0CK2NxXyDy/d/INKLaNuZ3l8By7QO8hxBjhBYK5ctkbXb4yN2Fm833j3/v2cEfH3
9hk5yDB+IQOcboRoU9mZhYPDpgc2s6cjyjgmYF7n3LL7iDb1PsE7FnLJb8SdXcAH
iWyjGxlK5xHi16t0sbtPxSPskxmrKT5yy/YrJDGFn2ZmiOkrYpTwoe4DyDlzHxTb
8euQ0HI5TM9fNsY4bz5fhhy+vpDg/+g1jKpD0AWh3IVLlgKolrlSyhkws7GV4qUo
FfqGev6yGeViXo9bmTFvjZMXrdq5TlD81mCvxQ2F51hkrKbCjkk3v2hoLJIF3erP
NOULR/wmh0iMkFZl7NlSoxLXV3grepRoLdHJxucqkEpBv+37blmUS6yhz0qlfQJ0
x/Y7L2jRjoKGavy16cXdUucRSNKsdnZJruPTBWeNn+dqb+yAudzvr0xi8OWPbqZd
oMIoJdo4GQENxFFppP+kG+0WJXrc0inr6XyNEn86p7g0I1hDfGj9BTIQXjdfVQRA
n6zXb9pOA6aOfZd4mkAal363OAiN1QDKAgYzjQYPeMe57c22bn62BPlAnhjmGGB2
g4jyrYG/fBXt2X/sWW5rE00e/RhYgjNgrmpdog/b7feilOK1WmGTHgZutuGFWSkJ
2L6RZDdgoVB8nDP3/xzo9XWS7PfrjnUlZjMYdhzPHFRJpKQUdYI8miCJ9Do+rsrD
KryKzkp6U6iLvCtaqbwPPszlpswMlp+PiMoHx60oZ3lUIffPw7DoBW7amR/HJyjf
X+mNRmjnsJYjEv2kILpiSegat5s+P1sqnhgU+1XM1bfLgKeJVDDLugqLNU9n69u2
ShAVHYVEWiXaWPd8OLqZo7Wf0FQEOdqrWR6WIgklDJ27PcBdhURcnMgMDvJcw9C8
pMP24P5v/bX/lWFLkk6NiSSIkgFz17sBaHNCY1/eZw/cBicRp/4jsD1+2U9iKv1Z
NWYEwd/nE+h3rlFIezXR3Z+mro0yowA8kYzGfGZluk8ieqVisvOoFUfO/7nBxc5p
2UdOhjYJ1CzYYEERhrXzuAUp3CMe8eMcp5NW98UxtMfFPbSjmlesgvROSuguukAG
Zj42s7EcPoScKizA2tilZ/NlcGmbJGfoJNpmgf0DPPo2GBGDMGny+nyCOOqcUnxl
mpI8HbgKx8JfCxDvh0DxGpG5+ksEw6NzY1wZXbZYFgIVJrfB/HwH6FE1ayNDIoW+
sxMQnyMKvPYultR3uZiGWz0fWQ5S2OPXLwCiRfIfapJy3L4bH4sTT4814sRM66c6
7JctVuuMIrewXZPTmY7w/IJ6eXKFwQLBnWFnDdEUx4NS32OGykxxtiAS0O1dsWr+
ntIBgmNKncii+xZ1kxe1KF6QQZOqv0PijFhsZGrgFFQSjOJhcJwk/Q5OgAyB3x+p
Rjnr4t+yPYPC72cYfQ25dbpsZ2Gys1pC4sh8HY3Poq6XqtUbeM+LsMFljL2MJ1p4
IaG4ieFO7x32Ksnd9nYpUSJzx361/sKpkXWQv1En/4ZROG4H7UmACO9N1dS0UhIB
lOKmBbKk6nzwKhj1JhnJ7GJknf2Tx/uXbW82T6QevpauowA1G5HkORg6S8gzLp7/
WHAPo5YpuSxerqOeAJ12sv0nckHR0Vo56SpsrL+l2rxAGmqdxf3dxV3SyGcxoolv
064ojvlkqSHfOcYY8DmxbvJsGJkLcGmZRSRWWp+e8eI0aIGpYUb7zLKwVkRxctmG
I++wIk0gF0K5nFCebrf5jRuXVuJLhMRkxavnHAhuYdIkN+TB/Ojve7mMlkuykakX
5JysCM2eK+vtmNnVgWls3X+T72jLjsEKw8doeKYmoLlxa3y4meVFY1980FhSmxW8
YeWps1mXOH3j2WVs+8zI8gRr7VAresb0Y8PEW+sh0mxY1Y6qDVF/bX5gPjbM2jI6
2a0ucMcX98IOafxwI8KayhwQgxnTw5/QkfiYXWrLA+2Y5EavlPTXwZh0GxkJBGz6
alHLSqa5XijUpB1U+mxWlBfpx8qWtkUEMb67fSklTuOoFuj8KrLVdY1ANMntXEWz
7ux/DrfK18OqQXxSOmN6wnwfHa7Wj64Jz+0RFXrXGP1L/6QcmVN5x8iRJ68XK991
1woXujitvs4uD+28KhrOJA3jKWJ/4/0NlkVcMS+u+u/hfSZNyuex4o/1yuD1zR4T
obDjFrkVI8x4my+mNLBJ2HhXkGOXVsYRT0Em1Pr1A5zz4j2jIsHqEmfC6QMdcPmk
mOb5kVWslpoqtNneM3VU5NBkKXwNLFzJP27HDavtQCP4ku8YZtt2N/0Em1PMQeDL
r9meV45Y1S9gg3zxWKQRoCOZUx2ClAJLygseEDQj2krbiyOCNno7XRzrCR2VWcSF
58YQTdFQAIR7XqYzCzACE2F4frPI8sZnMxcXcGxjYqSJSMowIGuGxF27AK9KGx0A
EYwT5e//QsuJ2pmIi3cWA82ES4OiuEgPWJXOIoEmu3YWh8u7ssSwXGmv8j/F2NdN
+y2/V3+5z/Yr0xuf3QIXbxjTEpQSE5nghhvNd19vI21kCVZMkVCoNGWHOj7/r0dr
MUWMd9HVQ0wt6+mgC5edtuG3kYdQM/4VJDv1/irWTaQ8tFMhhAGjCm/nTT3o3IMi
JaDOxuSQTRsUtuxjcjAlGbGftg7HVXne3nIyIyH2bai4S6NeqIL+7ksBZQ5K1z4R
F9TqnUAhX7Q8xkSgvS7ZK6XVHdUT5+RlHhixDbVUQJ8IyLzfTfrovAYSuVJka+OQ
V83NkK+oZP9L9HS+IyqrstItn/Ifgqfpqwo/+UZTyl8QGb7uiafKeOkV6b8ECZ8m
RzFdAKJEx2YFAx6FTa5FmSalPIqtmcSTvODoxx0i+LutMLj6gVj6UPk7Rki4MWFN
ZcpqjCl9wKLLdJr+iswrPN9f1a7ohgY35kUoqFCyV/WFuTWRJpzh00HiymqvplT5
t5/hh64yjUNLJ22wP9fbkt17wI6S9YUA7SB7LLWSExAXJXO2qAGoIYCNXNXgWl5h
F7ETjkFWx9YsmltDxkcRTxDWr5al3vb2p8p++cck41K2XGPd0cmmlVDGbtb7yzf+
//70r0A2LlFGEPQ3X6BbqP2XeUL4RBpseTL4kn8TC1cGtBM2YuYW2XSfumnrFh2E
/k5XhAnZ2JCL71zcyEcAECLF5zHv9wqpI+XWLN5vhur+F/JhGqy/5qE/OR564Qaa
KRFFDOMOsWfnFTZTtFMbPX1DT4hKJmDQCx7zkYXTnrZxCRWQ9qCeQ3bKXUFUkFsj
vEQco6Jofw+7sXrZEUNxdiVYynWoj1IuMIkyR9oZWHZCa4QPo4GK0cPakawDVNXa
8uUE/SRF5zVi/dQQX2uxLzdudLWepTEUHLTbtmjNEVOc3wZmqcTW/4/3WKYcOkn0
NT4ZYoYh6dAccQdt44A/Q/HgLi/vyoFAXm0pmglzzTKEPLBeKdkW/wIBIc/+XMtP
+Y3CpWzTjLrWjspDORPBW4LCj3gx7U+uys7exDhqDTQ6xVElRa+u7X1aKtIeo8ZA
vgRaUCxTtZfAMLop5vvHZPXsCYSu1Dm0D+m4H4M0q144+56SbsAkD4WcgJ7dY5CM
Ph/C9ikb9689GNSp2v8J+hG/epRWp2xN3iy7AXUs4FZ3XGdLlW2y944pjYkL6r9z
6KmIVFlJm/ttZmKnHqhQJZxK/InAopPgBBhYzVQOoJVMf2cflP2I5M9tKaAAw5jS
vH+HhAxHgE5g33w7Oe49ccZEHmW8lZBlB52LykwXJxo05LHVbS8kq6WfDj8sB1x6
6GeEjnYFPothckctVJNLwj03detEAGlGAkK/CyrruqNf8RlTFoCZUE9Ddd2CrdKF
FAkOHo5RcrO64I7+vf7NpwxR478fV6TyEYYMiL7P52VZ5bXbPqZ1GLJWWAsTNYLR
4cXulh4lHnkTabINcDXhu5grFLbPwddCyhWanhJYP594/ZOUgHU48Syx4tlYhdhB
XH9UlGyk/7dX/S6VHS6glbY5vAMJV481fBnJUiRhQaT+D1o5Bp84xaW1BKzJipA9
jpPM/184a2OC/fcTDfF7Pn4pi06ZDF6HW5W8gZsAUMA50RzMWVx5Crd6RD99ampJ
FtjCC7ZbpEOzm90Ma7+JjSNqUzz2b+GWYDFvZZdEFOC6QymxKAqsFXU8wir8WBv/
Jt2kYqs7HgZyWDOXaxanzuhXePP4Q9wmxkm37yH+Pg0P+KQGDpDRVzsR8e6MshvL
XS6ilQ0Ut/AUBZpDL6/UuomrZ/jniOfFDR8SPrraMZ88TwhZLfFGpwe+U/Jf7L3O
DTcA9to7nZ/IzLAQjA9OrOrFDaRaByqvZaIGB+WkXdAeA79f5GDLoyxq7yggMaWg
PXzRXgNN+8xJgfrm1oJw+aXR/qA07p/x8gxfPBM/yo1CtVx7gVLyDRpGh9Lar3Ua
mwXSb+IKy+swmY3MbMWqXA60meMnavv9QUYnlzjR7tu41j6EEqlacBIxvfP1xhY0
GcU6zaLsC56wpI0gMFUXv14ylN89iJFQ+03eD6nl3dhp/Vf2QIUUWio7gW+gcsuf
bicKxoIg5Sk2LFzm4Dpj3BuqUINej6PMLU2V2PzJLvnqDHq0zoPl5FBiuc3Ntpwe
LCVdoRiI99Bxjat67cy3HWxIP7Vw0PPG2azmwiZoR7LIPOow0iZOFuG19lMGetJc
zT230nq9LzMrlDhbNKZeBc7umLy5v7/9fDcTKY5aRRUEUQzNZgm+zymVIUm/7LGz
ggDf0O7BKb5j1W0ayyk5pPibU3smHka6/lvZbBtxiXvRQAUHD7LC6XT8zEBnWqh4
Im4omuB7a3KNsVpjMN0DPTaXR+/vnGa/f+bRHDVpLzJdGdMq+fQIiIsbqS0DenGy
OmRIEs/B7CZfgtjcpdxSgtCwtv1UH7PEK8yj7+chP6dtSd9C3+BpTe9TEbOqu6vK
7qmir6MRMEBfEmpPlweDSXCYXBtKR+jyf4n35j9PNHRaTYwhStmKPpIqZYmlR+9H
uL1NoiMbEAcKEJKw4X3ldMwDxp20soA8/aD+NtrU9VkK33qJw96+ChpyjuNtQSzW
fb5riFSHL3L691hZ5HZkhwV78ez3yxTgDFGx91m7GaTksibpH3n5M388Q7QHSw1L
aLdMg5RdwftZq7BtLHoD0Euecn1gFdw9o3PwvgCNmkbGeulLMpOspP9U2pqKHZ5O
dxnJbxJ9ATwzWSS1B/IG95QQGskncVEKlaxUMhp+WnncVv/OpI1BNagQuAuY2DQ6
AyEfNrxJf6ZmzjmJsX3LeOK8VrfBFgUlQXI8TV0w3OkhkJ7MWZoZ7ToZOinGUPl4
1uM0V5bIGHlBA+CgcE/bAW9OVDZHNfACuCPiMBuZfEQAbkLxug3SCe6KlNp9Gcbn
j369BDDH0kSry/VYpxELgFxXD/ZDABDuRtSsLC1/xITF12bzFH+Y9q+s7xyNK13n
xihbudnsu8jQDsepzSJROObsVIon95C/VFRmzpR1EsRQZMSUqo+jQLauygCaFfTB
bgKRlo2CiSTHlDSpowkZckaLtomOyTieS6FOKE4hO5HJz6vczfNxgle4iPoSdEls
pQmyAbUzYFNSZHOV8E697Uyqfk6fPbnLOo5Jx6Tr+slDPCnzIu7qgQHpZ10XVZ/y
OigA2fgsFG1LPxDfxzdfZdfNu2/M1nhR0a07IhM63UPbcILZpt3aR2r4xTaoVg9r
xVez+PA5gJLp9PoV8qOIZQv+aj7woBn/10c48qUhMew8MI0r8l91nM4aPpjY/w2j
W5XxAAOD2YNW0v+sPZkyOYs8NL6Jf8jG+lZtbPBiNIRQUWmFMlEzkco7wycUm9BO
QmHty3mXMjwt+Xu0Zu9H+z63RuFIXx8U0SLsvWNIX5POgwJ+dmyHRtQJC80RwQZB
5K9U00T/J5Z/A+QNJxxS6BcmJyto+yqRU/iqP/t8uZJz1RLidJMINL6jAtJcON8t
fw2I6o1ty5HGqAtGhSVtsNtmcdx95gZWzJPffBVLcARROcT+v6ALte44qLetPyxv
pBfONqLbSjxQobC/iv5T0mGEn5ZCRWksd0xH0U7z+h5s4VxNVeFsN974jy5Bb78F
MciY63YGA7r4vKMG80d35DDVqMGkwJYA8Rlzv7FnLg+ofteiFZK7ur0DLRskOjfr
Qiy4VvgWLraHH/kiFWAKgW4bDgykKw9vZbpZGQYsrfrJjUG6XX/2pCeX6UJPCGUV
WPufAqY/8wr8uUy/ZdYhc0CXab/CGwgwDtPsMslnYuYB+rIDoMB8Kt4lp7NuPs0v
AFzMBMgnSZ4K9b41UxCr26nRHyHmH+rrxaW2dCPbyVPo9GCogn8T3m4dGOgpzHh4
HLT/+4S66OUCuFfH8Y/vycH/AJszN5oeSSRU8I10jx8nNBhbl9aPCKkh92yaLnhs
sbKHf3sS7Z7b7zcfYW0zWr7kx13lFH5oWg6wixh40grdgt7lP9dx2n0NsmPtnXEn
7iiWdEmSdDJCA537xXSK8LkltRilYjHF+CNAoTOPhzFKSF5tMXEtcDJyUoHgMF12
XWt9v/HgDHc8DCwoHjPhujdxW6hK/rmWbA7BumGqMUm79qR8D/AopBQQUKeNp3hy
ewMY02XvCd7nQjn9b9Q00AHKQb7WrZbYU21ZglAOldHl60XDmuFs5Dqdq7T0MH19
m1pDiTlUwoVnCjVnSnfrmfURq6HA0wd0cPgu3U50+xKTjU2zU9/D2ksN4/Sb8csd
z0xtjit/hpjV7YIK9FNKlTxeJbCojSkitulH8YS6E3aFvmeA9axS9n5Ku7D2efDL
pyImqdm+eOcObMO8EaGAiinlbqpcOkCYXgMMCp7jYXLormQ9l8XImiuVnPQ4wYpY
6m8IWV9QF96KQPkp6v2f6fril/AuwByMNXS/k5pw1UXuyMgFyT0L5q6G+04TaVfv
Pab0ZE6Re4btY3huBvuj+RZCe0F3arfgjgOeopI1sD+03jD+nAEHilxbg2OuAhiW
53jh6kb4P/nxg5xhNXQTvkYUDps6jp4aCCUW/1JMjo/kvV5ezclVJ/x8hTTWiHkH
bRMYnIe8TmmQQ+Dpg3v1H1fWE3h9q782hb6qw8C6PmbysB6pozob9GuEt2ZS418z
llzqRdJgBbWq5VpWUw1VwObeMadzHFbI7iaGfS1GQstRRKHbwJaod6oxSGc+lROZ
iybF77WrGqq11fHrokUzS5+PUHy97WhSx5sPybzBlEfTjnIYR1CgXZrTZfXtdCn1
oCxC0QnGO5MWNX/6+/6zA/tArjipmWtadYTeKULja3lfIKG9yd8TvAmlPA3YCyh4
f41RRIBkpVUL5/KTJI+aE9RV6HmUbTNQyZNnsmmhVpRdilp/FcLYvP6D/WaYIs+1
xfUlPTTK5+20Mm9ttHyIflW5f3TaXYQStxT+yXg4xODHBfJC7FtjxDXtJB7zZZ7R
n+Y55ex1JiKKrTdnDtONvfhSAzEZCB+W71Wc1JWiUj53rCTAb8NY2sQfln9ZXOq0
1gCroBN7f6vkRN6KOigyEcGd32DGKAh+Ugdo5W78jNVVNJ5R2mXu5CsAkqhYyh1r
Pz+84P9hn1xeiI6OZlo3MpeiX7C+kffBI820oSTRETZL4jlWEM7DDCrGwjd48kI4
5UOgyuAgdC5l30URYAswSZ4pZFpzdipoKlqbqYX3FLmxlF5zkGPlGGkYYaouKIBU
f7aFxGQSAK8f7n9G8OkLhg6FWg4ziXe4Vdnk8Dq4kum//4MrdiNBI5MtZBE91yn+
RudgS6IeUcDaHv91TkBhtQjvvAGd3jFZs6USymsWtl3Y/3S3zls/iXW0R6LF9G4l
VBcvEMUsof1+2U8HnML8iA0rr53Ux39LYd6+IJZQhnhVtvWqZMyHIZ3DpI8W/6bg
0WD3Jv+D2WHt2uiSq7xeMA5Cx2l0BkliNNe+dqvjbysiYxNg6COmK28OzUE+wmIr
WjlXiIS7GCvO9LF5HoyJ5HEVrcXdmqKuunzUzKTs13gVhZuUJQPsAhMcgFzF+lW/
wb/RenUzWDjfXH/MUaIZLULtbMkkmHThhZT673seW2uNEEpYDwg6KgEm2DezfHSa
GZa9hHvebv7UNEWI8ggAwMxryIQuVUdZoYdhezokO1CN2Oj0iplkePYnS1eUQaQA
wg0/ob2ByinseoHSQSaS8H34HZYSfPotCjeAoijUEPVKs4rzhvSrtoRzW3d0y/Yq
SfIyAQ+8Je5n8HnJuvijB+p2iAXkEgb8ACXymjSzC04qRBaV82vIdL1KOLzOtj5i
M2VxRpusQw3eXvpavjilGUjlMwpufiNhScCRgNxXF9wzfddAA72rw5qgLc8/Fr/e
hpAXl3ohNoYYepKp4W1iLNhn6mlxPB0q71bT9qet6fuCM33ngMyQDuzAg6vf8GDT
awqW8IDcNoFqR58tqGla7DLxkSYgGeXpzgaeT0PBwxCSJhjhon1PfmotP+oL73Jv
H4MNudjdyDBK2UZXzNZUTtbTlqEChdA7zlKjDIRHZ25nqTnNyervXGPcf8aDrbMm
WMvePKy8gFyYpmUuxjzsRisoPSJKFteI0rgFJ4o5d+FnAipmk1Qkj8jlMCunDK2G
qFwReH7U6T3WYnnxjQgNahwDNpklNIWzqISwedRdkTuHO3SLQY1DgqAixsw5FKZq
JpKODJfquVZ/P279OM18FxRbOocMPzV6zIrFK/fL9KwKcFcPQjrKBhTZJxLE/jeT
IMH0NjGb7NRZqNOHu2Iv/y5nYERusxUHzZ8E/6H2490bMqr8CxyRpqdkWx/NFTBb
W1kGFoKVnNwmMBKlddDpD9lTjbZywt9FIBWt65ltbX488DWseK8T/ZyahLDpMZ4f
k7H/rTGLmQZsykDISsxU7jpiNkjLh4h/Su0i7TvVRMu8LSIo2y5q5RA4OwfP+Kat
O3+NsePGdxcRbG4mCyJ+s/iP+VeB/fcKEgykNITQJ062RiLRW4Znj4K4I3vW9Gru
Qw0ZUmQQy77/oTJF/x20Zm5pDzEeD18whn0pEQUKSJIaHjANp1xKfm7FIsWwkq+I
eWpLrFuTdcB1l5BahgLEtQdA5B+sC+IiI4mtDoqxdsROH4OB4rywaZ1bQeGhCWGi
6ygBpmsKS2Eb5dR1t8aYbdrfHwJkhphwgVhmzhnDRJEB7vNmzvu//F1LUMmENANl
xx9b0jUJES7kJkrs9f1Bnis2ZqBBHXJ27arygkbTFMcYxEE+N1yzd7mi6gPl/C5M
QX+UpCuMTy27VCzHbvoaYB8aJNYfufqWMZujvx1wgBwi7AW1t3dgJ1K8/awr1M5Q
UiGy/v/iQW0WlTS2DozjOcwEjsbCPzlhgJiT/PgVYGq90HgwFgHsBlPRWICLVekY
r9mCw9VloMYGcm/hrzXgChquHas1akBnOqk3Q+IQCNJFb+LbMo2tdVNFDSO1eB6J
QTPUUpWAo1UAmEJ559y6Ow/pJQnoGBjRrB/hr0KdGEViaUDY4+CLs+F2julaYC3A
c9m2/AV6kLIK6Cxl8GmAgODMv8H/1jZieODcTaXQLupMPOXQ4K0b89xA+9rJi0AQ
FWfPU7ZSaiW/F7NjWgYHAm+vQ83/GIUyMGuwkkOxyOAu+Zgf7t1pSBAIjhrW+HUE
TD0FQ1xpKMoRmiTokFwSM8iaFRWdNGfWBakJvams8G9qHPhZuIj5cRtwKzGpK70r
vQzyvKLqt/ChTge9oHbN3xkgjzctVIoCuMQmTCpBbQQ98r0pAkXcwtzXirgJZEsU
ulpg81A0Szb/YGuXq2brVq5Z4NwGp7Tz+s+aFx/AGfv2yEsWf2S5hVe6SsOLOy2c
xGfi4nQYhHQqRfUC6u6EQUuHyGA8mARXY2qpZrBnAsATrjiM3KmY8yeUsNZtQqE/
yIWI2/ObsP61eRZE0PDEqP91RCUPmWIFiSGRUe0aNZWeMgzC46F9UCXmQ7C1rpxU
tR2HNdivfprIa0v/AMn66ukLnzQUC7ScKxij4onrFAbCC48P0JYnTGN70RUOvKeK
skHveimf7P2D+WP2bdq9QaxUzpdyH5o9yOK5Ne0PwWgXcbR4PYzyQ4l2lZi69zIG
anvooZ9/JightP1KwnABnFVtTDr7jIzi92zc/7QQTcJrsFJYTzvNxoYjEyKh/zjk
l3RHiluqQUK3gQTkpzmrZC8Q3bJ1jYMn0WiuT2DaBvSVGXr2yhTb9TAyOoagXAox
t8hMRzpNmTKXLACxBsC86dvvcXlKbwTqgM+TDBb1WrlmAwu/h2fSnQr858dKZGx4
upDT8sq7sX/rlItG02MxD/FUb+BAevOcM1Liy/DxR8rrxy1erj+kfxUDIzl57Yhw
zwDwnsvLBVDZi6qHHF7kW4EjRhfBFCw9GT6trFPSds1w8h2Oo1Owp5HXqmZ4kmar
Dg3gPUahoTSfgxserDpNG9UJeVsl5u3YLBMboNNBbV/GL1CJ0tu5llrVAgACxaQi
DNB8LvHGGNJ+mNpOTWgl7uMlf3xeX1qSXY7NTBD4Ftx3iAtYSg06P3fPRztLDGmw
LN0IX/Z0gqBLE4Y0Rzxg8SDEuO9nqXVNQ4KvOatRlZSLGvIoxl2szj1rInn9ykUq
bcFpko45wjILhOGSIS/rCmOPqUAjemCpL16yKdnVR4EHvfaTmWJOYm0cx8CZjSMo
wLKjwYpzuAZVh3mxCtchKsqmvwJ5by3t+no02ySxDuy4J+R0EeZBa7fjc70Nw86s
HTBs4mcR5cRdNOZxt/GIWTjkj7cZI72Vs1iI/kX2LFDVlb8/TJFcqNOgILm/Ojxm
4oRATTVvpFOMJS/TAi6mqmHxB4hj9dK5Z+6JkweeTB6WXg7L0FslQMbgzGGl5mHd
RKvQmsdbJI7pLYPE12N7EJjcpKjGtHaQuRyIobP6IaJRqWgJQamNlkh25Lfag1Bl
1HMpQpOI86Z06oeyZk8LirpsYWuiF+vGts0evduZJwFxhS4ovbJfMQsYn7v3UK8x
3S76WUxhUSF5eI6P6cgfDtiiE/6/IZRe6oLuKWWsdPfwLsl5oYaqfOenNqh2/nfU
MhZRA3F6W3BFtszLgDQuiuqKtSUAwnX2wCEUWxFpKIIiYbcVHkR9OPuJq3MBVmJj
kxoY3Qtq2UdbfyGJ3mcvZckVyVWSS2LrWPNIUWhpfB1JyK0sXShBkR2j0aceTgNE
gcXsBFFpFkFEUji95MjwvOGbmG/cR69ZIRqjL6rbmQKvI7vD7pTZ4dYRYU1NsXqX
NJovFrKldeIq99xk0uWHre+RteXPsMuXpAtavZhbazMpjsfOKv5JfQ0nt5yVPUXq
yRiRs0GAMCGr91fYBJUyLWneco/kSLj/kGv5vTfH5Cb3vF65Sf5wFBUjye7/bxJ0
N+HM08mEf4UdO6UCqQilycGo4GJdws1+IgYSvfI6DcVpuejNwGfsfLvhgF38PFax
boBqKPkmskGdS10LjXEnMTj5Ae04k/q7Bh0q6OOXxlhJ6VvbIfWMI6UL49bEnZJj
MQou6tHEZTYgwsZBAUbOtJK+6m4m9D1QayuTgO53ekti6EZ663fLSreqNlcAzy2s
ktWh1sjfZG37jHIBbCXzlRyHsJ0ByVOmdg+1nZ7rbbVCPVuVfBlIFNIh4zWCfcoD
dL1IiT7vc5Ou8o31lwzc+TQRg7O3F02CyTfuRTuvXvpX+ARoFXrzdGz2vu2BDZXp
xkyuTA3kskCbf7QFzkvF1yMWzrKM5wc+X0c5N+GnpGKP8gihSirk18TjhtxdwfRc
Ylk5ixTiE5ojE+B6Vf4iZcOQiZdmxWzF3WVdf3s/jG1SeAs88VCclLOEX6JsqjZU
G4ThcnUuVkBwuYGm97Sb4Zzt31nNm2LuH61s+pcfqEG1GCCxH0Cv+MReeuJdNxv0
rBoSdTmnDtFlN1qKuEPVfdDM0XkD9G98FAL2u3YJTj585E+0f1emeUqfn77vLbGJ
4LsmFnwwhLhk2gMbsFBn/4zRpxauHVplNW+vraNKSGBoqdzIkHIb19O8XW4QQgn7
/Ekgv+V2cYMeDFs/lj3rqmWoHNMrvTc98NOf5PuCJNi8+KJJH7/RVZdVArmjtiiO
w2m17RLAFHlXY5sqSQdQN0CzmsvQt8l4tn3uZaVRxxWn//OSMje4rGNFHhcMcI6s
oTtala/MlHTkRpWDPeTObMOqPhTuuBG+kvMqavt2RClPHq88X3kgL+tFC7C0xNPv
1/WCgZpd5GdBbOLnCt7i1abzf1bco0Kgs9dnwxarPZ1gVd5d7OltfzB0xIen0V/p
NXGXJLdsPHFX3DuyhO4/Q8+RVOkOpbygsbkQR8TjzKq1iGzwxNFezzWEQXMRt154
6cR6pIWoN3jWj/nA+ABcC9yWtC7pUzOySjWPfrZUq25NyrILrT8wXwRaVkHcvCwz
ukW7tmcy3xLKdzeMn3pHQ0PesZapu/Tcmtc5k+8urIeFKGZTsyDR8RB9r3gwXdzd
taLZOmKXdNSPSi5v6W/bryPW79mAosmVYVX2TE4kWHwMW3w5EMGgO9CxXQCvHMhd
OPhgI30bggGpo5FNjkGc9CyJzg8fbK9uHynDVSKBwkGKsYS2FfnBOqG/WI3p/13q
Oo3PA9FOlH///SWKT84+Yu1TzgIDNn1KIDG+NXgYuHuUdmAayaKj6YnmT2Jog1Kp
zUi4GivFF2JjUJBxpsxhCkEbUoijSJWs5TP+DqNjrrcP2JRjC9B0PgfVrKNhaVp3
OEMAFnDs0InaMKe4rCppwfV+45sykCnSORdvJuZ0F9LrEGtrTvcEV0lnEePvkRwj
NpKdJZVkqic8DZSh1Wqyk+9H3R6KZ75V5QUlgzClpg2OkZOwiTmnIleworppgTEF
ULQDFXap9FlMfFzqHM3XuWoth5/T+H1aIeWWwnoTJr2KGFc3r3sbId8nCjd/2I40
ThhgxcccGfw/j8phk5z/l18D37gTpg5eLYOdPzTHedAJpaVWZ0529iIeFrXFxd8v
RnXR8J0+I3NuhJoqD9KjbNVVxEOKYnKx+8OXt2/incCJJ6EpKNwDftzxS2rcUCH5
qftvnwveoNaWyFEfzRG1MRacjfQigRc+o6zEIfg3Y7Av6lJ5VDGbdvH19pObRtmY
SAmQZ70nSxju4AhH6S0nApEkSfew7BCeVZEjtgAwXm28cRwUgZkjsJ3adJ6leo36
Ikms+8UTwRiW38FbOiEA8BnwowoxZzB705G76oeKXKKu/3I742qZhZ9xgWTlQScf
8ecbMMuSaQFtFdMZQJFXHRFYx1GXjJRQx3ndjVeCkZeRiYfuFC+sqNoHPpdp/VOL
bG3jX7S8wQZ9aPoFluqNdK4cbgXfm64eiDv59EJpa9ei0nBhXgb9V7yDuz3cKrLj
ygm60LnykUW1eFbGeGpLDgV8sp4F0D4HaLonNwzrlG8Y8wrHTm5MdDjAc0MO3FHN
Hl/IM7iBA1CY6bDZiGhlYV5BsgEL4disdD09vQH7zusj2iOSK/nL1OboAcmxQiPd
EOygR41SiS0cLY9KVEOsp7FrR9lg+JsysJGAUZCgU7ExXNkJvEkN0b2KMTcb2cDI
aV4oWA5DQkY8giiXbtwAsboma1eQ+ID2VJj4ufRTNN+mhft2jQLvZnGco0c/0Mov
93kTBZ+e+6Vx1FDZGYvMUlXOOHhWuLnLpHR4EOaNzA3drCzDgTfC4fG/E8br6l5v
paCCxJlhigRlMzLNrOOZLbobf6GOs+zHzDhR0N9zMdJ9WTDQ1X1YiWtSDSMyFk3i
t3WnnoYn9T5a9CDBu9VbdC88LMsxn+z9tUUgUQr8KssH0w9NbtU9a14WrVX2R3c5
hNkAZg58FWJSEL1c6123IwXmA206kAms4X5k3gaw9IWwNIIRDaUp7TPditEuvGcT
2+Euj9mLA83Rb+c5SAsjzrb6CFZqkCgVqipZqaluOO5sLN1iE7EQh7ds8RuConaC
nXn+GXquK/fM8dtosL+/S66wqYH5RS0lMz5j8QE8Uvtz8VJhDyAYp9LusytrLiDL
p3Pbcpa3Z3HJL+dtVOcZk2P2d7bRdl75N9DLrRH7W3C2uL0fdOgjLODJmiITVN17
ql4kkrdBxCers+vmXV9LYXRmOI4nohEPG2JxzIZuyDOPvOs6H1wmFgMWk2s3WWCS
QYwxlYDr4W1AXmr4+zttH+zVYt0OvBy5sXbiFOGonBUOX5qNguiGo4y7wad8FQni
Ml376nH7c6QpftxUZeYtVA5qSt1raDrqZFCQiu6nK4NS1vUyRbpfwfZ6+pSHQ6em
ipN+eJudkQENjteP7qUlnaCZ3Tvdy37BnFl/tw9m8+O+yWpZ+wyi+sDJA7VZ/ASs
z4aI8WsDAkRoBvzTG6LjBUUW/n+mIH73WajFxTDKrMB1MSePdMpGympb0CZjzFs8
5UCUILnISetQY2TJ5oLWacSYRjfSzbXZ7OzLw3iXh5j7EecGvVAw9EEldt2beOWI
j8nEqRU5euRKabB14TBVjQI0lmryUjviUd3Stu0D86wiEQKGJCI5znwEfKe6xOM3
zxcvblzPy0uToV+MBncBiRTRE15bbb9/nqHqsnNCmTeY6ll9GGLhB1tu3w7cR4rC
S4WpV5SW/KJh3pMMRmasa4aNTXCels96GCG3xw8TTRq2m/o0G0VdfOgH2nifKdXz
vMt49+jzPualZkoyfIEFgOtvz4J2fgQeQy8QMdz3/KBeYxRLO7ESsxhO57RWGaaG
x8bVs7anLPmCnoY4B0l2DBcQpeqPQB2J8+Sh8PEKlq2zt2UlPFIunNU+eP1wvTAi
g5uunO6Za5wySGXvCcjpqyEW7TDrvytzGnyYknbjuK/jx0jwuXkLaPUiEXbIsBWb
X2oegukIZQOKq7tbB9SiB14Kobts8y/ocgpzfbs2i+kS8f5J3UdskygsCwezxCAO
5JnugFzt/9SNReCNbDWhmXshMzqKTiN00w7vtuLIBY5VfpRTVDTSHFZ+a3CiZyHl
7foCKSHPg4zt1eI4A1RvDJInuPd55CP/K4KGWkJ8FkQM4Sj6LSYG99iKtovZRawO
lG/DkSSSU7uwjQFj4gcYqZN72wnGhATfnefdj6iNCiWV2j+UweY77E7ymks0eORQ
zsOdnbMvqnKat8b2qw70KGTHBbNh99ZtYWV7+kap1+IHNbMfXgGx/k3L+5moRfdK
u2kh+zBzEzF22jW/7C4iDhqMU2TLhM5UTTUzJ37HMgHRYU3JySSVIBB71ITmGWgC
cU/ZdLF4jdqB+C5zZROyVJ2Ae3kQKFwndZcB3cMErUjOwdZVDv8xDXCPzvMNYUC3
d+eHxDYysVqV/92fouEmh548jE1kuPsMg5Pm34MWVoeIvvqrpt5zdzujgYnwAzCC
xCS3S2F1TOrZ8H0eMUkhhXvjO7g0Z/wbK6nATbkcWqcPNzWo0ikJU+BdWXvRcta5
szU+/6tq+XOkbhA2UpYYfuuGZzJHQHdEjCJHWYvKnw3cH9q4XFR7V4JN33xsdC3c
q8jP1rLzix05f7o8kr0D5wkrIDQKplXSE58t7q1kuGjrVhCjMjlIPsOXhgGRLMJf
1Er8l/IcavWR0lrShw0JaB2n+CQcqRw1Fe78mGuSWuHlim8QZvHPA2nBMHczoRgd
2ullkOUp6A/xG9Shr/r1nYAQJ70RgkvYGcoongB8UnW8whw1TSoPtz0ZAJ5XnU3+
7TzT+rZKHTMZL6SrtKAFsbxBwC93Q+z7KWek6soHD+oWLNTEFudM/H8+dY9EHO0o
N4aEa/F9ncqp18aWrkvOasVd6KGQpdmK6G0KBhbDrsSBg2vyLKoVqFdXgrgUSF/f
+/CscK/huuQpUUPiDQMZJ9dF4d6j61+cS48Fl1MS3UlYkKGI9YNLH+RC/1kWD8xi
zTnO8NafCiY86zwC06syfjKp88TR3fSrsopGfUgTwuPCUGSgFj0x6kAru+rvnnPS
6mAoKfOkQHd6dZubnfPWRelTxgO8qUl435zOyiboFCWGsUxvfN960L06gvcdEcPp
l6qamQOc2+Gi60XVWnkBOqxYZV9l1vJk+YTnl8gpZ8UNJ5y7SzIAjT0un+Cz5Tje
5CAHJyzZTxoqzIa3tABrhxJBM9C1AK36eaOYIh5bwzi0VkrrcMHM2NfOdLdXRSSl
neFzaindopV93ABsRRcfnBmgGMnT5leaHo/hyXRkoMCCJZDx2MZTvuENbFYkuTZS
1CLIGOA3PQlwrHFPYqyrXjB+gcRR6eQqAh7sy8DfuTabG4hpjGlTh38E5fkxUTDW
MhBDpDSWV8wPJ3BekObWjrCt4risLtUsXntcSWGGY2KBB1e9f9lb1qgm3mVl8XW7
ivAznQvUAWlaTcqV4zlZRqR+Bv9qdFdFfQp8YSeEhqZGq/9q7XtpakuG/IEratEh
ME8uh8U7vBbpylZQ1pmVOPG5jCGdyw70gACKcgN6LsL4FmLXJsSZv3RMo0adk1iK
lEG1IuSgAR58DsrQj2PksOl7lOj45ENKEMHKrZWItpA9HZ3l1pCga2tQOfgmXUzZ
MaF7QxoyBd2UWCOORqXNhatD33sc9YpNkfo9+hAm6gVXNK23tnf8DH1N9QADzax5
dLeDwb+9sFso9V1yiVreDbwAF4Bi7uv8zBNpjTvvZz91vvzP5A2xKuRJNAEthLAU
VfGwQauYUJbyoO+1PGCYOSZUkPu4thr1AexorRXiELJjmYg6akbz7GlvGF3yuCLC
+8OHv8biO804h6OZnA2sQMT/ETAsvI9tpfmgbq3EsbZ1rGLWhMinKz09byrasgr5
XUsl0xgjJMHbM9WsJnarC8UmKta4oslOyQ/FYaXgh+gShcIkJphTSFZFBFkTHLMN
UxtTMm/DdwB9H+KpyB79ysFA5+egQMzm9id24CEc04zVxi3K2L+4ZjlmwjMLfVOH
YucJW92mTxFC4SgGSUnzPycHJWz95GsO5GuJaPZBD0jfOhSlUTPpZGRMZqsgSnI4
NDF4NKuMzYl/fL/dZCu6IaXgjv9Xi6KVOEv1qxdTGxN+RYi4/RnSYTUec2kszVVK
lpiy2jIj9ZTx9gdZMRfVwh82TFo4w9uGiRQIjyPiBRVoVOxFiNuHjBX8Z5rmiuBn
9UrE8QaH/QtQvMlstzjp1Gq4yCK4tz4PwLBxowUFawhukt/YF57URz1ujVC6Sa1p
HhWcDq0vLfQrv/yxln2k9tgG/nO3X6B1tEzEkgWnQearvYdAjacUXS+G4M3bvqkA
xzkfJ/nUZVKvpXeTuwddSraFML2ythhswa3Gz0jUBIfI/tRZoySlevnXPDsBjqoO
G1fRz+4QQsNEs1ukG0vtWR3MuUFdCYI0WZTdC0KRo6ulHTdIav2eLrgVoUxFR1Kr
5pv2snhmXvS0FSzGJ8CsX/QjDuYShul0uV93ynEt6yVSXkLFknkkdMcW4UdD/CNU
neFoFF1bgNrVRJxjDJXCdFWyjtegcsQocyQKg+zA7tLeJnsV9O9ADcuaxM2lPUwI
+3Ja5vBCwMZF97pA3c2+QDIYn+XM9lvrku1BKFzmWuVGbhKx1OGINPu2i3Uu4/hU
XO9RAWfH+7sTSXHIKlI0PH77wUp3syz7iKIBY0Eh1P21ynOHrEW1iZU9a/m+nOyr
MBT5fDw2DOsve/3SVYnB3dP30zkb+vLS6MThMW3AITGw398j5cLodqytdUFtdjX3
CS4o7FmtRyGN58ZHIzB7zsSyiOEqLIfgOdexHP5O0Ju6K0TCoDaNfk3d7OHnzzCX
q5aYh9fO7lX/4tAA9TEAgMcEwdwCQPPrZxuuJZDIX6SJFqNZlQWzXJur+dmbJ5mT
VfBrIO4cgvC9P1VJh18dxrYDLsir9g7GQlUOWofrMyu+2kRvH8sG7Svvz5v9ZvGi
45QohrS5Cwsm4Au97nBrTrjzEXzt3MX1FGOAOA81D3JYpF6gES0BkEAORcoKlm6v
vY++JteZeSYCabHHXOtTtc+ZnKR7H5iuhTP/PeOAJBO2/r84VhmwoLID1SjMPYOV
lJ3Ly2vEK+nW7+j9WorFjES6HlxluDr6eBvn0F44kJMcGzZqJ8VYJG7d73Wlz1Vz
goTtkvAEw8RpDUUA2JUFi/dqbQa8NWgiu+AqMzYbm7lN+eq/ksaPzD6RpCXYvqN3
cQm6R5sUwXr2G7R3Zuoy2pk5hX0qsvWFoGIim4rNj0aQbKcjsxVnPQeweDM4uAwc
Nt4UiaxLk/LifUebT8wo36om7pjK9y1wrm9GZqkCeIYVrxJ71GLOCyaPF2CBY6Nl
E26QslasRLAO78oGUiqxUmVnhk6ns09yhUrc5GSP+W6YMV9ygY0uNHgUAlnyawaf
cAqDpukLVBCXun1UhVOxqAVHuZZbJj9Gl/erYqcCF0Y3wVsAsmHPG0ebwmnHun/8
bz0v2JOD/y1iLyoghpcYdrcVdC5wP33Kwr//dc4jf7Hf09H8YP7kmwt101eeiMGo
nioGcdoolHrf2E3hgP++txFNuxNyn1aV4b3lH9hqNQF+rAoAm0I3ePUSL/woBxnA
kKJaeMnxr6ptV5j+tVWWwD/qJHFjpDiZ0P4xhBSXAI4rGGR0XlmfP7Ndk/i7/dxh
gAvo7fmkV52h//zJwdON2k1xjaZRZQOoRPbjoNuVBra/kGjpHL8YnYXOyI1Z02J7
UOllfawgGg1t0nhG1003aMMBMbCg5aMFg0HM2BmgU31m5AczakXFsTdHOVNyUAkF
dvEwJELFx0CwMGH+YP5T/w9ULHBA1DVkZpKyVHSZNKBLdTIYNe9NArodVMKndj2k
CQcrTt7TBxJArmHyp8/a7IqKymfV2a58YYuDUOb9EaOOSMP3Aqd5E5zgZilooGFP
UWt0xEXdXQF+I6I4Ti8qrlA9iEqcfl7+bS4fdnpMdakEZg/Nk5doPyCKElNOjViQ
jIwpx9591cAz7L3814ZvljH9oVXH2NjvzYGxfI3rmdx40VwKhrv+/Z0E/PMTcyFA
nJNOdkeRr2+rIy+lt6ROAD7nvvuv4UdobDgFB0o5elVJYhISU6J/U16X25Ex74xK
Bvq2dYwYCiphiYn9TKGFoptUvWGOuIjNxqCLT5wCsNpRba9BXx375htASnmsaxf8
iguNzZRun7TzMONE1rhn/9WUje7/osyJkBFkvSuW6PmkOE4ve75HkT7FUmM380za
z2vI8ckJ9i5lu53r7R5RhDUcrBBiGCAsYeY7AMbhEikeD/UTrLXLG42AnNORq92O
eHWjOdg613/d+3AnZLdBoJwZQlQv5qrqyn6tOFCXzgU3aOaEsgUKJ+B2WYwMltap
X3xNYUvfku1+63qLBPZOH/ITqp69OyvPcT9edQLvUbVjyxW3LaM9inqOWGZPdJgF
bEw6vff1lfGwi57haBTrIWd+bjAWcZyUxrliZ6fa4S+B1uuOb+f+6aCuIZBW5vN3
YWjw7l+ILnB7vbErJ/jN1qqDTw2AUXqrYWIZfiKFMjrVSTNdjHAAy726HIJSaHNq
nkpkdwZPetmfodi/DT5oA9Upxa3umw3Chu19jodEVm39wiQwzDusaw2f6dxz/ww6
AirItOdgIr8JWO/WYyra4C/PwYvb1eYwnZfzxCDukmfcW02H1G7k0KB75rBeoOhx
1I33jlR0/AqZUfypZABvX8fxNBgfu20QJpHVlOfwN9PJ941BpInLjaNRUvwlUxP/
9Ntp/EQJEXUAIV37E4ZJcVlMFFthO5/ryoUjhmUW/aGIpUpor4KFJov7+2lrRVpM
/F8Xca6yNJYtI+AXTlK4itG7yGwnIFZ6sXFrziqa48sPNS2zYTp8ooOJ+3XBc9Y5
AxCYE3H4EPPVm/RLjna3pcowQ4V/P0MiJxvZOx+qKXTQG6Jnc62apotK/ImZI6pD
8jnPJr1OwtMRl6QjpreKffMadNUVjlfSfiJ5NEyp9ODlt9ptNGGjdPuHH2+cd4Yc
RSZpGeLB+aG0cerZ8zAbI+CN2Zrr3XugRacf7wiEAEO/o2JktCsvSrlcSlJAVR00
88BXieZlzFVIyVo5CxKTE+VweHAWhDDBXV52+eE3rLFfMBDXM2IuNgWex3ysY3jb
A0dgdQf/TDFEOgnpDAZeUCeuhlTngDqbKTuv1wL2rYwcCMubgRJDqtGqW38LL4Lo
yXhCt8qRkGqc7jqPMyYM/I4AFLnFKAoV2O1pm/75Mlh7njOLBXvngXkj3QrUeIE0
nMW86C3/RdGge8Q1+ByPrRNYlu/vKVgjw21UUc9WOzwnliWse+hFhsFvMX3F6FUV
y1B1SGhhT/FDls4vZn9yotpb6UZM21GzzpeEdVbdMHORvbjGPWaMSKu1JH9I1LuD
KWdOIorNBrndaK19xI411xbxVLaTUGRkUbZmV+FoaOPY9P8hJwNfCzIH7vRktbcx
8+HlQ5C1h/GV+qqAG52EKQ199vlTUENpAVMHT6s/5pI9vTH6grEP9XXmvWTLEmxT
40K62zKSPq5jUyAnMDYxqyz4wkIOq58O7otq5PTz+I44dTXVqWZ6zYvOidWRQhlJ
3yI4ILi2pcyKVomXVImrmPFMrY39aMro6WxuRTAAtQcUr6Cvj0zlJWMH9lUpQ7R+
eD5zavx1N1vsmLcD6DuAIf/Ev9JcKkvzs5HaPZ6FA7MqUWpbuso/J4FD+9tlBllV
6bhXfR4LujgfbErUzDSzkd2j3FZiGDbb6+GCdrXj79k8RL3kU2+LnCfRpl6uZbFc
+epJur+pjPcS90qBDhJHXc2PiG5CVXvlEFUcayoGksKNkLDIU6+qKj0NvHMa7nZw
E1f8CoN4f0KUKGCDcHzlz0Qs0A5RXCnnPCc9+vM5k7ZLWX4Mm7VkFC+J1LlgdAT6
8sEeQazMrYmMH7DI4Ityve6c7K8B6FFRov5XXyxGiJgEf4VUBbqTKIDSUauSFxyV
PNMwu104TKbiaLtdzxouNbPcMleTqUTMwSjNW0cNMY5Hnz2iHt6J21IGSt4Z3Kn1
f6czmIKwgi1J/zVI0pPHGXNgJwAllZ+JBTV+ihBVsOmfFYAQ6hj3gGoScna8IK/z
IWjC4WLK3H0Xu2CDoJBOWz8DHOacit1S7a8sgm1Me7CdJKW7LVukLrH82X52Wm+B
fndjsnJ5QZONsAfa6xIkzW8C0xI0CBF1iqvUlU3AUk9ElNQiWx+dc7qbbPFMip/A
SHai68XPgkTO7ThkF24KbtoWTO7TMzIIIM5LbcXK+jyB9i1fojhuHD2JQRm7LKzV
UN/491kk+qnTn8rAEa2kFnP4cA8QZ8lgmROHnlh1kbwE23Jf1wzd6F5g4GZT+dkK
K/AxCBQsy94cHWoMZ1zE1YeOOiZQZMukV3sk0jiA/6J5Ui7OquERJlqNK8mM2bck
FTN52uk6/iRizPAqPgBTLbmD1oQTBOPpiTv95NXzfaKE2MYWH047YbyT/tST7WTm
wiPfIdU5rVGWn1jNqYVMa4PTLSGCqf0+R0ZqSIlubkvMoR2Ei6lgBark2Co+ci7L
f5Bu49o6fcl6cBWSgJRZx+Z5lT37vtAeoSCKlkDTX1RjtcMB6A5BsNMg+5supEBC
6CzAGOAdRZLhave4uQjO1hybR2g3iG1TlJe6vb/xaZADfkG/Qr30kLGwWjyT916E
podGvT7PL1ysWbl9AmggXAZ8fQTV8QWqZzNz6Gte9quQUyJZnDacPbt66bZjjuuM
IXsumaBqcm0+rxGh6fASNqR1Rw/scz7LXk+Af0beFdQpCIAO2bLs6ydWT2Hgo5Yn
THSJ3eiT42Byp4Mo0FaPfPHUEl/CQG0v15+cvIj0G04BnvP9OvT968LCb+fUWwdH
xBiXYHqgG5ZJpulX6oBygX7qLX62eSAENpkpt/vOr2Xi7y7EmgUsvsWz0m/IglSm
jrIktzSCacAcD23i4+Q/6TPOM4wi/yQtekUu9kuemPDbQsK1hgFFL+osmg5R1JQZ
d1UDCqLPnj0X1SxZbGARLE1HH24U9FZ7YwIj71RfAxu9JCj5ObwgLnqw1vKTXjSR
LIbU94IYHarqm5IKXofn2bmLYUMB+keRua+ly+WrtPSEvEzjQ7ZJC8it9lXDrCG3
eKFIyeTrKXvPv2bsOCJp4SkORIbo0L+fum2lQ6hpMxWsyBjeTg5pgnntVC8N9Y4c
DH1ZD+AMUx3/Sm9uOJQwWkwWGVh4jkIMF7dYB7uopEqcdenSiykUmke2CgkM9f2v
yVaZIF6HRTajL+6QOUtB1q4F0sfJuTtI60QrK1m022LFjgcp4slLITsngfA94wf1
uIge8PSp+1OEo3RZ5y2vIVQlKAuzFNDYuCQFfUR3NWYS6uYmluDcLtihfVkLe7ul
EuQNV17G4LIMEksenetUzeP5/SOV/mEGBhvG9C+QLfH0WLWzRuP565Hn26RzNOdE
GdudKBjw14Rsn3/JmRf7h12mDUT4yjj9BOYHRwaPwZO7J2TvTP9Xg29WYnN7B2sn
Z0zsCqVgehepNtXoKAsUjhNy+2ga9PjIV6L3Q6Nynvh32Csx4woULVKS4BE0Pzb3
tEBNeGsyBECcQEiUB0PjDjl5S3oDfLIwVmw/JV+yTEYLw9X9IfcVcTjLwKMwL3wk
uJ8oc4T+kr9p5fcNbkYzVbgSDXEmkqxQ9xsL8HRe8Z0q4g4qCuDlv+9rEPuDtoop
9Y/c+9S3D5qaQ/Tg5e20MT+LW3KMiZ7HvYbOJC1uhqbVfxmXsxHur6uiXkMWWpyr
h5ulJ+/Y0Q7Zya/6ACbkuTphWyJ1XID5AUQ7glaVxp3nbMgr3VOWZsmtLjymjGbb
zuLi+zx8sdB0xu1m9QqhyTA1NC1NUaeMCwiuWram3xJ535U9m9QahFQHX+hiu+dC
c6OpaGw6L+Fv3qCINLkjqsOy2NjhDx42y30mL94OaAC7IPoUfwdp9SMJm+2vaqke
qJ05Vqy3Oqc2SRH4+6BmrA36vaPzr38i/+1NSABbNcvFD64x+DpH917C03pQLRLP
cCOzLU7ZO1E8gOv2z5NO/GRuTD54xGp6xhFsxHQCAxox4jKq/oJNNA/Ei43M5S6n
313KZLJ4ORYS0KFsIGfTw+Ep4tUUesjJLTyMXhUcNxAoDJeQZjW9+CFZDAZcD/gq
TVetGsE+/p+oScD8lc44NPlNK130SRuHPKX4XqQrgFi90DfVBzms2bvmDkZLwL2N
w/bhuFnPrHXkeoeYfgX+kfJpGI/lTk0w+peawmWfKT+TDVANGBNC3oL0H4cLborv
m7M9OPIY8ZSNKMyq8lRnq3eKO7OzZVgWbAettnmAcq6gkqoaKR1SgaxIKeU48wIc
DD/SuINmHRWXEp3G1unqyb8eR1whQ6ud/J1sq10K7kAjkrjoe9b2lKLErsR9uEkm
9v9WuchJBUgNCdqukRM/F6XC0KOk5sIExEjsjQH1v5Rvmic503yb5S0WY8L1tsPv
XBfZZ4nFz2LrrHSK3fGxhT3QkDtxZ/8TEVuIQESkWuG7CsC3xT118ylFBo6yAHPt
x07krx++6gF/iWI9DXGEXwO3M1lL0nUk31CGJGaIqzpFs3J4d/+xlfzpcSwEBNWE
rWddSxyHAeY+/zY61eapPjn64oZouLcCj5b/Q1gIEaCfyAFGTOJZBQhkYdU4cnup
emZKtNKjpQBQ7fmcRwiTjULgBxDHgtjKhCgZ2kVxgsNGy/hWKhUwkCws9KFYiYwC
rU2mNpD4ZaBxxDvoXAgcEFETvD6jZaUCUCZ9f29p+t9e+v/SrG8uKTfODJ1Z/p7+
4iPiO9XRy84F7iEEIT5KMt596A5BFZ1NI4mSXQhq6rrb4FCWCXloiQg85QV0ITzC
4xaYTnPWXKFue9hEpOv+Q0j5WOmMDPcR5JEghD51UfdkVzKfsE5KxeCRPf8btzME
I24W7LtUBHWyT5Nd0ysJZeHsx2lzyL8AgK3GjQNwopPZIksI1vbX80pIDiNddAXB
YWcnMom+0RhV9U4FMPfrSsJCM7kMtqJAkb2JJFKX5j6JAoC7+Cwf78AGXBjHy3Xc
IvJ+48lGOfRExdbbjisjo5/7SWnaO0miiYgn/R5QGwfEUcEJbHhe+l4QZ4KonjSr
jBoEEY+fcP9EYSsFpoU0mQoVzOyZu7T5kxGdW+cXCwCqQWPt6Ib5qQDuY/mA4Cva
mJVDq4nCJ4Ek+pW7O0idV8018SnT1/taDkachSiMOOGK8UTq3mDnTKeh+otU9y8w
PjpZ7f+mkREGyPZKAwvsYOUHsvZjhz1AMYNkhx4vayjYrrfSml9BpQmtrpqaC4BZ
OeMnlD3f647lAY+Wi8DTjZ6/tHYUhNu9Pxc86Ye5j0DDnroGoi1ueU+7bZEMq/zS
jDsz46hTYA/g5p8RyWwDANPkQeaUBEMCfQMgQC8K8hu+7HSkdX8RcEhkqKnmHCNx
j1z3Q3h1y+btXMv2RdO19e0G++oBjYPp9d5BvTYWc7bz8p0UCEmaDzgpX4vCHAun
0M8Xs+BIzuUlbnY7cLIn6wp/k/Jp2Ctq+svQK8D/nuMAqpI7nuQPXGxuVc1ZSFcY
m6RV1ki24LtWtRreWjsw9Uz/cuzIS+CdupI4mNJotBQ1y0WaUmeRHoj6RSbQHOXG
jvH3yiZawJNNTO8YYFQ5aWogpqvoXEau4t+3qqomD2QPFxx6zKLV+Z1/O97Tk43/
ipLyrhR2+s9aG6ggNK4uyXJEWdyQcAGOYUvVroNuPzITmwrGnipIm9UUc8Gi81bO
7taI6Y1kVoqrK7yw78ggd7DdXwLoRwMRTkTi6IL16c1STd90PQHHgUetd2lU+Gqx
vJjS1V0UdK1OQ/dO3Au+d3NT0Oyx7xve0H+Wdice1OwZby67VZCk24i0pDjRJ5Wo
jYBs/QvSvcRtLar8LT/SYsSbbotQ+uNP/csHxHSXkjnNaLPXHUWJ5R2sbaK0Bf//
pzwFrG0inYnaoZSDV2+/WWpz4uvu03MZQTfK4Fbw+j31MZVdIvv4ZlobcfR/r0Nd
civUONEF1VnVfYw/1+mcncynKwRRRreEhfCOFNv+VLjxoz9OEGVoKWSIuSIuPplQ
kFin+Ba/QjdoVbkjRa7O0j71IeREONdO9yb11L/esTEEDL384zh/AhRJZyOm8j1N
tCfVYTwLNdt0M1LuROW383ziqPabzRSUNNo4B8Wr5YML4w4+PYpyyzrmXq4/c9Z2
KmapP03Jta7+GSpXdSCBsZQD8k6moNFqEOwhNy+Nln2acFGndoCNkJAlFqIiaQpj
fcUKkVaXni7pX2sLNTPwipSDVN4KBx0DIfGowixI/QhUuHGn7uAtg3BqDP9Laks3
RDSgC+CubPscVfnVpm6dDVcfojL5OezrDvfEmfZ8AdzYiUq41i/Cuvs+HIWLK/rq
2RPdEVXqIik6sxNF5dWLZGkA4BQj5KgfZYdH+zpBVtqupMQZdw2l/7yjEYH20wnr
tX6VBsQrlUbqnCyDhzhwNczYFdX+VnL77MtJyNVnjY4CDzM6WyHm2gHruYcM8OWx
geV9H5csjc1D8SzAcvNupR37pRYVeBrlfzbZx0rHwR4DAuPqHZ4VhIFRMOHlyWTN
cvjPgzN8W1+60RytCnpz+eMAsmnP61FiWmrim5rYyGFh0jhuOWxkQc8QY2mI6IVT
ugutZJvshvP3oUS4vB9WyiDckw19nCJ6azqS+9bPI0etlvbqfVPpp2AN5IwlE7vc
VEVXsYzCSawDEiE9D14hUGDvnAgGpjKlDGWdjyRrj6u+F1Yqmli6L7qBUed+8NYE
BaPhiZ5SYee0DTu0cs0qZzF20NEWRXmBm4tVMhX/dlSejQgYn//dk08On5FYhogI
jHmaZ2n8kbvUOkEQRo4zTk2HIEdvgIx/1sewW8T4JvcqeGM92a9lXRYAkTDNiK5Z
Arp8cvjaOxVCf2pH4UseK9X4ITTiF/eW7KFDS78V0YA6NpgLorVu6OMdkgmHWNWN
CFWT63iG63Q/dFfgBusUe7o6RHbOea4Plxom4uvNRhJsZG6U102Fa8XLr/74A7sb
fL0BySK4dRgs2sttZj0NLfoFiD31iPmH5FQZ9z2pNBs0YHO7xGuO7U8eC1AZSufn
6416jwvXVlqtNjEMuCG8U35snAklgXvZCtflWcrBUOrfTbQ6SYiG+FLB1l2fMuHp
t/UcfP3wFZykBpjjWtXUBtZzQHJNBnGcLqN16FvBezmTGElHwmiuUB9ZvuPbFC0S
rM8xuoQ3B0qna4pdZVMF2EPMyMskA0n3KgZQRW5T/8EWme2OXnSnxpyrxSi3lmp8
PGrmc7UZjQYdAqCTrqztGy0tDnaKJcGZYJMmfWfGL/HpDtDLTAAL4p17deUZSlln
0tEPH1vJO4ET0uXRggmeR8q+tSBoX+N9swQ052blI1AOSgF6GOJk0yfjIGW9yf2H
+Wf73BPn3Qwwqh0VDlQFoZ8atdUmI4nMG2kf1Os20g59VdmMOiIGTYE90/kersPc
qHYaQnVvfiN0YymqYREVpS1V+unF90VdMPIvjC3RPTNCay7x24GrwhtqFzt+6kxf
jwkebeU03z0/AxyguQNlCudLZxMEVo7uFCjO20NEP+CpLKV2DWBRwmc+zB+Op8+4
UwwBmMNyRxExghaTppeJ7RjijQwe5Lagq7DSSAtCtuN1XrPE9AqsTwFn1Ls7sTw4
/mxdIgu+SIR1MMMIwv6WDo25V7nzv/kZrsSHu8kNfQWC1p/iDuSVFMvRP+6TcEij
fldBzyyor3m36hWErNbCwY/BCT6XVohDoI9MQFirJIXtDRAndT3FL8uvFyBucno1
/KMTyKIEFDdvHYpjOJb2ISAyh/T3YTAHQ5QOGKnfFbY5XCRIWjpRAg89rs3/h250
ubYNjKVHWOD8MisinTh0FYfg/cZiIC5WYW/WeptINrKxnz13Da9FuXmR0UHmRd33
fBwDzHFlXW86yBcu4qr3Dg0vM/u4dp5sJSeqUZsY5pedw+vbgLFV84hBqFMjUXiL
zA/tD56Z8+eyOSfnKX3yIcMrIVYaZyRPAXLdI4BscfdV0IzyTH6tF4VTX5vrIURg
H9kGkIRdXNooFBnUsHLlop/xfHwnfCfuhXVPOf4dIM5Ng6oER6FYyHs+qbEC3Ypf
n4npqanrUMzaQMwFw8dFObVRZU1odWx/oF8vc236IrgyJAIk83F/oiY/vbp4v2HD
9WOnJP0wdhvPIh3JrrJNM/ibvEz7klShcBB7fwgGPXOV+Xj53VhuKPTPYoMc7Nnv
sNuRC2ur8+YFxuCO3FjkXozSI6VrpdPQ3USn7qVT4LEBcYwRbpTww4vTA8MGeulD
eXcUBpkvrg6a7/DMbf9UZuV1W8wUbjWthpCgVJdfVeZyqdv2I6qylGuD7DTKOkE6
kzKKCeQKa6i6/L8gLzFY9Kcq3SWRGKKQcwsOnInMrPnBuHQU/WSTOr9O4tBHVzUN
QMmFL36AeF5mgphTDLCHtTSCyeMWdoQSiBQbENYd44dAfTQvVrN0HErMXqA+v66B
JypwVcw0UNPDSNi6iFeGmX9PI370YoyJvhxpEOpSBMLqwOU/ItgxTp2DpxxDbhFc
IzQO8S/K8iaYydInzDDJUBpJpZaKqFKjZ7yZmX01iUZvBfQ6OjqHg+frYzAxlAA/
MXnc0ravVTMQ+Eqgz6nTc19CYg8BrxiFTTYIi37ZbjoXmAoxiHcsy/0iG+N8i9iE
VzGm3IzOgj8jwqfo4u/ugJzzxZFeWrWtXKSmZcw1l843DovVj88Y8EON6yjcTy/3
hbmLNVePt4wgRE9hOCMaD1y7WU0RJRiIDtvFss2reL9NyczWrFqI0XHodkzO77xc
0dYJRmcM7MWx2hVAMjpfDthXLul43IOLdCrxHozsuH62853rTsxALuUwHX8xYJh8
i7gpHKVmNFRNxmKQPsWcgswtEnzgg4fLtnEOOiQrcbrrRIbNn47RYQJ1cLbhFpe2
jZUDMVea96kOAOSpf5PXZ7+N80IB7KHswu2AatKhHrWJEfHIo+nH27L22P8pZUQe
iQShEk5CCpQ9ok8TOoNTvUV+zfGtB2V0Gw43aBOm/YMbbEMTVK7ZnY3qq5smXBcP
9sHL1LtHBpDs911QIcfIiw5w3JKZzQEhPsWemp55pDZsxa3K/KMaNLl8xj5ghwl2
qcZxBh28KYDjAtQTnxfTSdIi9MfUv4/CxnXWE8pDYPzHILu9Z8aUQ/TlSIYeequn
qLidkWwjKN806LIXy1M67qkTPN/5YXvRWHPJaSkRvfYNFn2hIyO8/PLdKYDg1W0C
4kjtUKQXKK2SELdVvt2aevXS2+L/ryreKftSMNJwHeKDRJat0lLOL4Cz//38VCFp
IBjz4oPExiWWEf5c5vqy9TqeuxM+Bdd4tzLlpTK4+cyXPWCPNDq95ImXo/YYCAf9
MKRnkfwAb1Dc1EDIoRRe1k0sBMkKs8TfEwX5RCjHpmyZA6OzB351mhlxzQHBG87M
HywArM3NIl+BpyqMgynYPew64EOOozk+Z1WdK8HXQFTzDfW1s5ecvMY46LAwdxAK
cRhMxt7YU9cDXqGjTO9QzF4s9qDXliPX+fPavHwp5548xGyKmfEJ045diZ3YYjoP
yjm8BE7q1dOEriyVw4qu+f7mSw+oXp7VonhzLjeJ5SJFrQR/gdzcZxPseWIkTsyd
u6QN2jDJuyWH42c3ka/6rK1wn3/3XXRm4ixuZwprBQFu9N5rGsInl7RS1fk9gyWE
GjDydmdAUT6l9NUSXVEDKMkMxsGaavrp7vCDI9934bPi4fzbNGpAV6xwdw5thfOd
5V4Ouh7W9b7q8d3tEaykVKxQ1RSPGzHj7SuoTbatZHGJyPiOUmXWPq7+Sc22dzq+
Ts1VCyN5J1/Be6uh1eou4hShod26EEYgIwkdy80jHgo9QlDBtcG6N4PYUlIn9h1n
Ms/RNTS8D8hHdZJWLJx1glHrfzxdd5V/UOVze9lqB4v9sNg7hdIHcEnFC2+0MWrm
QH6mEZEXZvdwyqwYoFuAL5nNMlLiKNzfu1vZYrQxzZPIvMLv9gFEXtx3bsg+266m
RBo4VTqZMxbiMd3fjQYq1q72bl0N4fiy9UXzEzpOV3g7Lq/00O+Z2f3w4T7mrjtY
O0/EHloXnsj09RuHnzNO4UEJErjpRdMh1hji2bESxMkMQm5oOHT4Ou5S8tUrfy/R
PPk4XtmoV80radzuZxnXxnpPnzp7+lXiZ/53al06CFdEIyshvI3DG0wD2L8eO4NM
1Vkc9pIvaQVt/Vn1gRi7LnzNyX/najo/gAAPAv3w/g25SPR+Ip1oU4rVB063dexZ
ABNoQP81lq5wwldUV72NMxCXCVTwbIpsHt+hgrwW8eI+Y1MRo7zsmOjf7NoMoCqf
5ETbjXQobl6oJqhKvSyTD6HGgN2LxxyXbfG/JSwSkXKFhany320mqCQkcxFk/IPI
rRjAzRr77W4gDu/fhlslOe1Uv2fAeJy0PZLEwCeuIgn2xEXTRyjD1vVThECnSN1n
dU9xCq+m57ZHgtujjrNlYTxLMB2T3FA+RyoPCC1DpoVFRTDW2pi6sq5yXryM8Lw2
nGPvPN5HAwSZECOq4Ws/gAzImvb2A4l6luTwkU/R6CyRRVfeJWzHEMniJ+6SGKaF
Fhl0WaYbdPJ3+mNeksGPUlxBwphRy1N3R08t+CZHlbXYalMhaH3eSHp8Hl2xm8R9
tu2HGM/PMuxpG+Ibzg6TJgWoaiJz1MXpOndv9dhY3QiW66w+ZKdbd5W/dVDPLnEp
Hrssuzkpg0ePmGFDjdVHRVqFEjih0KzOM6mfqLb97iWuwsQ/2pe32L81pOQFMxVq
IM2V3ku/ofEvyL8oWwks0o7MXS8I0tVnOOrq0Q8HCTRHneznsN442xn2Sf4NDBW1
ygk+XaacnRdhRMj8xTDUQ6HJurRsmTnBHvEKVddAwtcfbM6R9xfG0MS3dBQBojYK
DkBwdYTmUq32Cakn81vHRrKRoIzzpWue1XitsA3QxBOTx2x20WxoRlK9JzSwpjjJ
rELTvTXSjgTlBypUsym99HRGWvAFk1XnxzQ2Lz3pm8m9FZvRXxpgW/9TyEVk8hy+
EgIIEzb18pm3SqD/hQ4/eltLU4pmCd+1fZkzgbQKVoZSgifjDicCqydf1Rnecm4Z
wE1BscX+6+892wVIH3RblPUmAv1yXyFV3YatLbA29X/XXUAfMfKBYQoYrJU/qfSc
337h7/pD4HOmQQ035jqxGD4JnfMxILlA2+CY6pe0MIdD20l0Do5IQ1hVfMiWiOuA
Q5j2MGLXbdwRsI8dOm5Xn5PlzvKu+/+O/LFsvMLBAJI1a55W1UhwxS6uGMHnA7eJ
ljCWtI3/lMEtFA7N9CEXST1ZzHHZpedEH59ZwLWofpTHoyYQlNDVIwKJcsULQbfx
y2kUl7dLHcGt5Ys9RKTRUbekkBjaw1IPFni6B0XeigZ4P99I+9kbGcuVd9N+n31L
kbyfJzvRNL2+esGHXWx1EMtppx5V4TXGNuEkyoUKCSWzCtO5xhKjhD+QbvkO6Q/f
ZiLZLutM4gF0YQmWd0GsOuEZLjyFyV2lbmUh2WioU2wVsfp5q+bTTZoCCooWL47o
B8tC1tNqGaxAN7wZwefbQSc7Ju6Wfh928rZ19Tu02baRyKm64Hf3G0MXk2/O+Cn5
k9YrHPovaTnt4+JSOX2La2CeIq88xASLT01R5c/IsuM+qCTKCaBzvQCzrzhgPRAT
8afVPIkspNjr8qh4hnF3gWV66FnC70Hfyx8yutXWsA5L86NlClWFjAerCx/JiDad
HWnwfd3EiMXwNzaK2rODyXFGG1x74M0VsodvRohbRtVU649Ua05QYYrAnDX1/v8p
7vMxP54bTd+lP3p1MVAbJcATpoaFS1vJAD4R+AsxKxQn/f7ultddUfX/0H8/uRbk
bDl+Jt8+Na8Ij+rn9/iFGkF9ZjOPDlZWIFZFqzMN6tbWtiNaYZweBAzjyV2nXICY
hdr2l+tge45k37NI8LBu+eWv8BpH5RXV7mTYEEvZMfCkDDJ2rY7FQpZBuS2gn4zW
ymDk97jhN6hfdvWx4wlhSH9HHbbD4ozMeiX5zN7jopfQdqvG5JnSvtDqZ3u1lsGG
IvCqrL3ERaZEQnaiCvUFW8mjGFpiOMMfh+5/v7tZaJZw/ssQutX3mwxV3hyTRVdv
7Hi9JjwHUa02kqjJfsxoNni4Ckx0+O+iLOnh6OUKes5dLyy6QSAOP+SXO9AFBHxh
LKmf3Cg/NiVlIpHuT4XB/kClF7Meb5pMNLL8WQl+g1UgUvggmS8GNEjT+yRedvMN
kdDs5p57+plY24rkO7NygUZt7VnQ9xiKJfQ6k1NH8qJ2uBUVPuHTuPX0dfz1MxGp
4e3/5hxlVcsDpguxD5RMc+9IoPK6qAByGdmCJnnIBlFVc0FLDDhyiMNrB7jCwRT6
BzaoJWUZXusH5ZtuTV4hJHkY5EIJ4Av4Ve0G7Omcu7txf7Wtu/5J0LQlvE6gDc73
gQxB4dj1jg/e0DJDgV9lGcjyTdtjXjb/FZVYKoSAz4xACFq8BktlvFfUgoYtUE6S
2+8MLArEgBrrPrnP+FwgJEk9GgxMfS3AhF7LRryhJUKgRsIP9XFRdyCtTEWOerXi
BFnpq7qoSIR4EI/q3MR5PjpY5fheSJHcJFZhZSolpSFd6IDFFxoyNhfHfnVdw2r7
9DXOmyrbbRCKx2RD6pkneign4MUsGMQ7ydxIkhg7BnMakHyXUBIGraWJvgtGSi14
oG/MqdF63/eUe3cripC7mnkKFo8Pit7/pbalot4l2khC/P3+A+6H1jbqdJW1jMXx
tk41AGIu0oSvubBFrI23ZA2S3x9KwiPYMPLt5d+WZ+MINFSXIhqMWGO+TlaNoA2N
/p34fL75ERWRjbZkdFaCl5F9uIz69N5u52Pt9PMFCrlmfRYiqHyNVIBOvgm3jKiT
cqaNmwpuRb7ggPL2b15gFNK0/Opuwpm8I7XF0dt+Bu6D2rEetzfuF8vAtH9aKxvv
qjnAzerrbybYC6Wz5UQPY6r52RDJRabA9cM1ZJk9e8Jy1cDrE0IOPxGjZ8LvlaYa
oQPF7H+O2BudVpA7H6h6LqCj9bKvj+X1URtcGlIalrm4H0fQykpVHQXC2WQOu+6k
igk2ibfRJ214E6rojXcFkqYazSSk2Z4dcOswi3uyKSLfN1+LtpnMG6R48ErefZIv
/R9/wzjV9Te6hdkkxvuuh4//u/tUW++M/BtSsUxN0bmyk/+CvQYYb3SftVLCbL9O
pNDiNgfR/uhxd4uwznMoBl2ymGP1vEv1CMFLXaCAVlATcMnwUI1VeJZLCIkLOMy/
jVhHnjmRhLsqm+WMNYVdzDvA4YJi4DXriFwylh4/JITQ/WeU+h3mMcZjzy+zHk6p
T/wXxEVeQhbIOKgL7zTS0ki0GhoMt1QbMvXXB0UhL3kyZ+N63l06gXSqhZi+fhja
/SEKPu+IcC0HnJlzO+usVVDAgflRNfbh0WY9SsLn7Lb3kcVHky9LebjzSlgIStTd
VAPkBk7LCF8luPFME3hn7+oUzj27R6Nuvo+GSNeU+Vjse67aE19n8tDeZicc6P+V
Yk35013Po1dZdKurs7+Ujuu/FECTGlvS09whKH33veb2kPSdu6CkR5qTTxwtoE83
TY86H1ca8SocISXHXnJ3wkIkcIEKLqgIm5SM7XaTV/YttZ0K6C3WtW40nl056KmW
uDbXW+LQ1t2UemfU/7qEzVfblJnW+rLAPq+drfKmhsqJVepcgLrTwKA8Q1pe8/WQ
5AbT7jX7vA5v5fIOK6DN94wk3rB0AvvpaDveVicwD+8xeFA3kP4ocrbItSmIQawk
c6zFc6TXBxaEjH48YXyI33VIcG0DuG5D7dlEMQ018xo+shPSX58GSK8CHT9q8Rtn
gk4HM2+u08fmvlHp9pjPG5wWizvhwIPRE4T9+/GQghR24bB6h/7Xt/9Q8Wl7407s
KRaFNcPZY5Mx7PZSh2NGfnfQc0MwSOqWhvcdvF6vM946TBWQjCogatoHY8veCCoy
HT+m6kGcJ67wBruaPK051LiBUyxnXUizDDkxIfaIJperN0Szo/pqViN2JQxgyRIR
A+aCTPokEqf9a5PFypyr6s8wSFaYULxz6QZ+/MwnXjCiIUPPHKWDLu4FNnlkZ1e6
xZO78tKMM7JnOPCbfeuX2hPNH2YyrA3rGI7EW+IIUOutsOWW+C3XmKa8EUg64pcs
4WtWmT7mhiNuax/e7LkMODQVAtDlKCwxWVu0UEflNYUZFcnjoIb728h+2FsdWhiL
e1QEAsAbNrLbj6OrNgxZKi0C4vb08ttIreWzdTVIljWbiDyrTxhnSCJIMy4w3Wsg
kptKvMVC53p9POhCFBO//4xa7D6TplZCqIcU/ZBaz70Vjp+soYdOtVAp29HB8ZjO
2uN3xDei7/N+2ihFmMRz232DbXg6mwtDacV0rxxvUJbku50qN8hCa5EDsmNNVgAD
VLWMg3v55qnVvhBtqmHoBdQPtUJinKbpmC3FdSHsZhgAGu6L0sJJ46iPVcRoDb+8
4B4oOz/oyS+zN2Y6zUYX5/2iJ9ThTScm3TVzagan1fJ83An0hwkBmgeo0gRSmpxt
x0Eimbn1+dHZHvJ2aYMjpMM1mw0ARidqtGz0VMkEgJsvmIGS+Ha264G9bTg8NbKH
YX6X1daZzU+VBRtDbO4iD155px4F8PCH6++Ob40SCkmxGbmr9u9VZ9dw0tWE6SRw
FYVqaV5qZ/ZOccPjU/fbHMQ1G13biqw481pmta2nSalFWqnWpY9c+pErKqfhS8og
s9auapIW+NzgIiXwtWCmzyQJ8vvfepJErUMvouZKhCRWHjqrLvnZmLEzpx6AS3fz
B3UMuXcpGx1Kdhowfw6lf4w3r5CNkJ7+2ZzBqwaJvacTY7Ax6aOQW51lzDcpQEpm
o5L3gfB/SNrPCuIasDO4Wh5OnHB02gC0tPAhdsULstouLA5XhMnuun2ng42S57fv
fqus9xVoZhyyCo0Y2FFdpGoSaSxhOLB78llSh+CMewJMYXGTjfsNq7AMacvPKdNJ
VNobgTFz6xaqCyiUXaYdzG/R3hOI+cjxAQs/9TV7R7i7E8RUvYpYoJ1d1i2hUNS9
7BD4++/o4Mm4Jk2VL1iM9nP91KLk++9Din1QeYdyjDDo+X2TpPfnY7Va7tAN2Slc
9AODajJAjmMkD1B4PrJSsBcb1EY33a5Hw4Hcm990ay61anuncb1DEXyJdZuBBJD0
CQEleeqetVLY1XIz2aUczPcQD+8lQYUZP5aDgTIkWOSkBIHiDlkE2+sdU3jC23O+
ttHD7ZoFwnMZLKD4lvbaJNYttA271h63SqblU87atzvtHNHp9yyoZhNuwjA9b/cI
5NrkOkgklno+5zi7ubxvuskb0JFkjQ7TOJ5GX5Hg1v+Tv82rNZLNb8eOZjwCegIH
kpxaiycNgfMfOEjjNuRgTbPdrYgym0FinhlV63Ei5oHtfKPw70wh8fBeTBJIU35u
QMXBav/6frlpRzIXmwAcH0dd7Dp5myOCXadze0v1crZTcNbIs+gNweQDcpPRTacr
0+txRHIeMN8eVRdEA6yrdv216jYl391xjSrkwSLDN2kTYWScVqVOqyCajF3zka0g
RWTEYDP3Dhe8tHp3y3lbxVzhvC3zS0YCVfj9xUHHeKnY7hvtklYd+y7PID0CeYZE
m82E8s2oBcbMAUEnBlEh8ZI6QESfqcRQpA66Wi/Xl/RK7OVf2JxJxr+5w7H00Nr8
jVyAe2W28+vySz+8UGFaquH3lqYvuThcN59ZP/AoZx74L7IDpD/uoT/UUcQSgAYX
KCzYQvWiFJWDZsVOfazDydjZlA6CmCt7RyBJ1OkO7BscTAfCIrzJKOKXuZsQ3n/j
gP3HWhFKJPNq12Gx2YR0vtP04QQC2Nbwukoa3AC85u7ynCW7JdL6I8qcUTFhtJ5O
O7thURjPqz+oxVR1JE+37i57OBGwgJBglMTPE9WCjlrplw/mH6X6YKIv+0xCqilo
ziPxZoDO8WdLDOx0WAox7sM6jbmm/tFKBCrbpAt8zJZulEJFK+1fWrfE9xzKkpz6
lNFdkjjxTJWezTnb8VRIY35fRiGT6YAdqjG7Naj/U45z0XbTtdsKZdaoPC0OECYB
zK88ZI9jfo9lPTOq3OLMFDoanTpLQUkIu9YVDZ4fidijui54GKNQAFblyuaO51g9
VJeb+7GDcrZh0caPjy46X/9ayWICs3Vr7EW8sgThBwXtjeQR3GnsR0IbAdW0UyqZ
WMVM2lSVL+ew7yq4w9ECa7BeBFeo7kC4ZrNoW97FFomlq93zz6ar50tR/nT0ZKSb
ei4WakXTspDrY4afUjPdFoUivSJo05G9cVeynRSotidD1ETr0G3WjbfGPlyfIGbp
BlBJbWSdoLINxFPoKrfpfssc93VhrrDYkRDpgRHh+M8LwAsvbj9oFsNkQA77HZwq
UhhSr2UOrb4K4/0uJRRUjqoHVDbUmMJgeuId/FLHKXA1GQc3NLAqChnfX8vPkUmo
RrG4gwRaoQLs6wqSuWESgb1hYyl0n/LxEreurinHpNNM81+S4LYMavu0pCfZviam
rV/b3Ui1bQzCPFXOqQ3X1t4Sidlzrh4Nn67zJT+I17uqiYoQ4RW4nVJfrW5cH7Rc
DrlH2gfqoYVu0PWYiAuJcWxkLDpfQ/crDjtH1zPvPdDhbRotkjTNUtpHA/UesgYT
QGOmtWuUTjx7fD1qJQJ4HYeAwyL29FoFzpeq+4YxbHJmn12cBWfrpUwgREcmIanD
GWxuSrwvBmyYoBFCYWaTqO9IGJx8OtbRq25oNszz6ua5toF1k7uRxIbEWjlPxmCb
qvtLTOhXDVvCw0mcOFCFmUCGp8ETLKD6A0C/kzlgDxuAARkXdULuTJat5X5SE9aM
dbDkgIkH/U/aF3JUcIyMlkGb6mexeWfIY3aldlAGdu6si6ObRqVNi5i2rPkTnazB
oINI3h8IMp22ka/sqWfmDB2qyWjoJZspV6RqT+ewgJeKgXFfzA5NwRdCBfW2Ac9v
kjbR1vweDzHiC2siWAr7vmmw08GMM+8M7XgPAxSN1Ex797Is+c8nQRaW912e1TzP
BmDqBpAmPt6G0YuYFjeD5/z2JRai45pC1gX7Cj0o535Wowid4/GZLWGv5hn+qK6T
TVzYtOrqykD35m4Ne1IndGI87FU8N6ffYlQxMewKPt4sROBV1tBfGzlB3x1UC7NF
OtUdV/kzWeFf1Cped7Fd8RptT3vOS3jEqwau8TFNHpDImLIKzsvzhZ8GWkVJZ/V1
qh5ZztbOAuifeS00qnFMcqTXwO3By0UVLoFsJwR1VJzRpAoQd40SUU0GSC7T1mwN
+nYiRaOAxP86QEX3QrmBrXZ53gE1GMGkwNb4mjSvTQc59eohEy4NqSdntQrGJDnn
GLLfEClQTcomdNHt8e7EEgYW4+I6zDHWr2CtxIxhfeojp15s6aSDFCA9MbQVgMxf
ZyRPQUDrDbH5hRaBz8EFcU1P6KiWxZeHFCm3p9iaQu+LcOlT2n5+3xAKha5dXbpe
N+SY7fgEJ5w3WNmCh/aac7wrZqd7pBgAKAaVSLqUXn+SMMcjyvz5TBjx4BZYyCrb
fgam8g8WzVNVW6+eRBagyf6OqLosM8mGRHhH9q8WYektDONq4WilvAKNEnhoAO+U
Xngg+2uk7jfu3mEXpyzykQwmRXk5EVugGJQd/mEmIcRje/5fEc1JEI8um+0dUU1J
INVf0lxY5kPhujDal/faoAd403bJgem1/D7CDtCbQL2ANd7Yy7rZrIXObAi1qDOu
XJ9k6T2jmE5Vz6DF9mVC24czlW1EVSClUAUdIaw8D5q7vusdtbYRioNa9PS4IEVu
SU8/VFkXjihYs37U+kOczW1WcaA0Z2HnMjYf/3o5kXCUi+rDFQU0gH8LBskY4unQ
hXkZTeQif9FPlFyPXlwm/GBYpduVSXpfPPQsdMhALUC1DdngbDoYoz1teZRVLXtb
+MmBxoGEiONb25h8+3sL7JsOnFfKaE0LLP7UHvjjIrO+qDDqsqvZhdPV5Elq42jH
grV30BK6zf9cM/Ks+AbsxDTrDx46PZmqG5dKbB2xv7Qa7EKOIKBjyz8AMrJUQZtU
zzduwpasFTo+OL+VgEEEfXlUZ3xEo6fMRs4m319rQu19jmP1oj0JjXI+MTJE176V
zzypPdPuF7H/PgVCM5RaxhADQG3fRVQpn/7WRoz4hx20OTIwlGmbhXgEmyiSCy6L
xO0XBowTvjTpvZE2Z3NaTIdo4YWX4AjSUn/zwbPWPNRNk7s4YYWcDmI9QKv0CI8v
OMT9Zj2HRXWaJWBT2lUV7KdUm8HXETPjkjlKytOipznyiSfiufumeyYtNmRF2TgP
LNIpCivYJaBIkcvSayfRuXTyuPqPTjUUYqdEyHEaCD9vyJok7gCvhO++A2U+oi/W
q/uPae+/B2UfrY10mwEx9HO8c6YUkbIK7MZSpgq1aHXC2lclaKPmRSyhMzOhO704
GEMs/R/P6hTNpLzzGdg8oX/Euu1EoICPnJRfnGMZ5akgyV/d6MjZS9NptHf6RxHW
2D7azk/pYMaFGL16+RGzwpdkZ2Y00x7UGBDgB62GPA/TAlB4frR5OwtzfdQ4a5VB
K/EBKXvQvb4GgZglrHqPKRDtlKVEAfo5EGZgu9V4cMGm7SCjyE5mgXEsNfPFJhsd
uDbanSamaIzWSiKFpN7n79T178wVYdXN2lI5niUo0FalA7/GjsokFKYT25vvJhwz
K0cLkW5aVR++czlY3ISpgCYiyAK8aJZ4+XcAuuTnV/jbYuFpSoAUObOFYRPvT4l1
A/JAic3EbTEvLUExsgHbMPrbmjmQSuR6rURYODVz/dUkoWZXBTQlXAy1vQ+hRCah
8Zc7qJxPc/KqemlYNpB94RRks5HNBmB9/3HbkNc4DS0yUlFLWse1OGYhGhTwlZkw
49EQ4fv/vtj69I2kqfoeFvp9P4DJYWTxiu9gX+CYRlIw5MuUsV3NFi9o980wwHq4
ZfnjvO8o3k/zQ+UsCh2M24C89xUTLiHT/s6dgJWe04AVO0Gjdron25pUU7vrSeZ9
hlt/gtdfSrPgndlCuA75tUtpV2klWwg2vIoU6CwQTXRAnNOOgiu/IikUnzzDUciP
RiHC5GeOkkx1unprl4kzF8Jp6z5xjcEi5okPNTkc1HrOoXE0fpx+YsMbZKooA6bD
6rd0vBbFupdTKxR+h2FtJeww38CD48txu/lW9L9IslVtLUBHpWiibhIX4eu1gnoj
bUerNvhgwUHpd4AMEBIA3CbrfLaSY+rhYaP+VcG6zeCKsuUgPbt9rmQdIzNGSgGU
81ZhqSizfVM9/sOyVCPA6D6LDbcUPfN9vSUrRRWoOviDhHHafE5fQJKRLhReA+f+
2AovWr6fVq7rsg4gecwdTR70xGfUYbJOHCMREXpePOeCCdR3mniFR04tnXQFBiSQ
LeGHDOBs5yYReZZH3FnbHb+VwuNGXKzuOhLMvo/A+FnU8AviGkith5K9aMltfIL7
WAnKKP3cC7+MXhgG27bHGoUWPpg0W8SqIQrxVgAU8ti6uKBqOi8XIU+Su7xfEEva
Ye4Nkoq3YYtzRgLs0Mbtzttp65tJUkWQxy7xr2lLfVn5zrLYlm6F1Ou/vU+SHJFF
CfitdT0t7TjD7jaYrAkleH3r9B/19tzyzw8WeHjF5YDBvlBwA3HOxtg1L7Dc8ZRJ
+iE5gTlhKdxBVnKU+jAJMlpJGOrTiUDUqcm5pO7tvemoV3vOa6sV6pVBWaki15Ep
HoUoOFJjs798kL3ww3rfn395T6bxCFhjsoYjiek+f/B3ArDgtfa/RSRfayi05DgW
1o7HXSWU9fXzEfEMD73UfGs3kFJRo91oZlgggBVlm7a7ctA4H5Wm2r/WUr00JIxc
xRCQPErgspStEHs7npmwVNUaVprNpsEqq17O/RAGp5p4SEdWJutJKzzhmSdshh2A
LLw46UbDdhuAa7yDToYWiZyd+5P0jOGCRpczRK1cBX+AdEhxoJP4jyN9aSQI+Ixt
5dTywT92kenR73MbCYFRUW6pq2Ar2t5I2V4evBJjbLQUsDtLIcr3dsY5S0Eof6ul
CIYdBhXQeplXunpKORkwkbdsE+pvfh0HZHk/wRyNiDTxL0GYebfooZkqRzFp+PLQ
nyS1DX5RW21UYVdp25GhSHNIAffU108wcb1dJ4AaJCn/7dCf56feysaVUN3+iyZl
mdZlmYvfQ63VqBDh01TWymlH04bbFs++eHXKby/njJcTL1jLmwBqCVUH/WNdSt9F
yy2frYFm/dcLmLE26q6hC1NqDyuBdV+4KD54CLbHA/KRIF8URxFbHs7ZhM5t7C3R
9eeMdTwwrqbCDVKegZIYRaMi9OQfOaE6dz8zlACWghAbS43Pj9SPfNFVn+cl0cGs
aRK98IKfu+EUp650W2WApogXADZJ7sZtAbcD+AGgyUeFUbbuPwqbgZFK3y3H3udW
W68oDe8q76t/olPnJD2DzgKgdd221NbQ7q/yBg09ynPkFoO3eV9c5DtBaVw4sMWi
Rql4VgHPzKrjj9yaoTIvOqxktmK55t8v6NTvHkUnGiwcCrg67e0k5qSAEQRCjTPO
E0ATnZm4LFZG9YL9mKtDP4uyi0fHopmNg4X0uDvzyMATVxvIFcGS/SoXlxRO2XUM
4zplf2yDeDAtqlU5ewpT+2DQ9zFTqXFmiOxlXd7ojQAvd4hdFPOmrxtikiGaeF80
yvAaRJJPSICit0k+Dq0SibBFthE1jKJsV96DmQF/0Oy1KFrq7sN4rS9Klksm0/jS
6lnavQuflTk63aN3HWxKehOL1g88FbDYSstUJseJiS9T+jiAESSKPfxFLKxoPW7z
g0aSFz/PT/51sUDFOD+1FjE8UdUDp8HpFoiq2WQpjRoC6rVqBj+4FPdzlqY8B7s3
gOonmSh1XOZkLdpbLPEGZaqS81E7Oc4l77/TgweVNOaid7q/hsVMjHqw4Ku1uNhM
2tDTi7o5+dUIdBpYPXw67rMxd2cLl1MidEEvjwvbPHa9JlMuy7JPCSXv+JJ0G/sN
QJSo1uGTzCF51ajhkmmHzIRV4oLteB2GK/ieUuvPD9ez4GNUTscukTOeOKlPDJ93
/hpFm1QcIs2l4/Lrmsm1Gkjss19xh1VVEX/XXreo0VtIJPIcGg++7d8qFjUkODv5
HHdHOMwXYLVOmyA/VI5i06q66NaY/ygW2C+YUWBXdFDuNfsqeT+e0jcyZ8BPrESq
9q12lniEm0Dud22dAvHrxwtzLmgTYKPQdwofSLgoV8t+jLA8Bl4/TItAhdkYYK9p
L1n62zBmVQ6jYwM2wBR252HFGPMAu9M6R4zExxtprrvhpauc900GCMPkavMQwQ/z
zihpM9j6vRQH1xNyzvKn0QuYpCk4IZGezkzOWIvRvphndSnKBGJDZpcLX5ooByTW
cUQb4YSJYVpWkSeap2mEaYp8T30IwIbN3BCHYNNKmcBh/+TlW9pQlUsP7HXnrgHA
B1iCXUF/E2vOjUKC9cot5cW3g4r3uons3z2guLP2JW3EPGaKL9QfUl35d+tYJaDP
utCPjNIwquXN10wwJlgrNeNxClF63I7/95DsHsuV1kSiyao9Qy25CS1Z0LjkCPS6
Pyh3m+qLU2Wak8qtjL9fp2aPpXfYiIwqJXErpT24uG1zMN/JaYBG9vRF/DNmJad8
2zLIVGYnFuvYdsuUekSlKW5exTUWoEuO/gVNZXKhT6TmMVSAINyaiuiMZHNl5aoN
9X+UNQmrpQiPs2LHA9J9vka7dTSPQN7aa8btx11hJrc1tT9C+/IwIHW26D6NRupR
HrKpbNWOXcPEIOXnZGqdnFINjOcUIFLOqJV+cFykx2dO4GmJycJ9eamami0tjNRd
M00JA4OvVztpwkOUmOIeyMVBHaAXTGSZxi7xsxEbdkFn2vZjY2LyeVTjGP3iChq2
X5BRXY8h3RpipxEC/db2RA+sU/7UPZsEi6yUvVTyo0mBc0UwaapLl/4wEhrFrjQB
BWJjyBV4L+hdTIyFcgahwRAWuOxvfhfmcAPm0gKI2HvS6iQebJRbSod0jLg1jZd/
0jy2lNp4XtOJ1rrdnEbR5cYobcptD4zRGyYC+mUU8nMyshYHNhHej4mba4ovtap2
nG8T2RuuxxnaILNdL+mY3vYowxK0r9OT4zEbwP3UNsesCmkb+uixQsAnVAOFXplF
rb9M1P8DIQSnJVJQzJuDXYuNk1+tNTgWeCrSNKfqT/5PlkqLnr1gLMsUTeldpwX+
IGyy6K8UMgVy6b6h1NxbZ+njAHbx5by1mpBxymIyFAQd/DvGaTaBbQ201ywvhRzn
6Pwl1up2KhtugXOS8h3ZwchOOOrrMmbQt5NO0LqSnDL+HwNx1VnPgvz2YG6I29fj
vleAxQder+cUscWcXDWWRj7zUyPfYQS4suxRXjXCQc5bSMNKxyTfxAANP0Z3lLeR
5lfUIDSxUPufaJwy6u8ewxzxmAGQyvob2aXybdJFZkG4RavYPFXdJMNExkGi0gP3
8oZZX9yPkeUOUMMHX4i6Qjy0zEfyDbtCSucbDSvKY2i0/ZYVGTvS/VHH0zAvqauL
bDQud6ptJPfv4LaXF+I+KvuatVZmEptfsKaQBM/qf3ZRKaYOD0hCC9W3XkOjS9Xt
QcT/Q6sWocnGSKKLR7fm85esf2sAyv9mIQx6Kycg3GdlkyJywiiH20dVYkrGAqcz
STXd+bih+Ni1v/fleVyqnbrievfPb+Cvc8b+JLK2kji4khjh5ncy0igUQa+bNf0V
FtfG0sIcE9xY3wXP3QJkM7DOb80ZOApJB4dGuP5qF8fbw9AR44P6FAzFgy7yWanH
dXJtqmG7c4Y8yzbcJ/DskZuF1GQWRD61Pk2cbIHumWBn4OoHXIgeZ5zjpJIRrE39
pxo2QwkPZrYkWKne5T5apblF5OiisRi0rEACsgeLCfFE2jkNbnOFc1wc//fRyMGr
uI92jDvlR6O5vHHBybE2EtHTvY14Jy0xGmhKzVtscLVocH1jR8dPRyILsMBOi8vz
Z5OVeY8b21rZuIEMpMDhhIlZG4R++EsaA+onnZLQfR0Itny0MrV1O+1AbIQhewtu
W+lzYONTm9thmCLpwUSfmv9ygRliu3TNs4PLGhkTjRdMdeO0pbL29F/c5dGXK9J/
ip3k53sSM10ypf4oQWkPRJR1yBqc4Rkr+TDVbxQUcTgj51eyiEdEM5urufAGZlmr
xS3D2C8YTwcu4Kii7Tuwvb/TUlxqRafJBeW/6W8ah2CMZnepIt7eso5P1W1dR3hM
pwNWh0bOzPkS4BK5T2Z0zxObeuAsuqMCdDhKajoN8CJEpjSuNFhvMWy+c6RfXhj8
bqxR++4wgjTtmNguoEu5jBA9xFlJmlczJisqABN2JVdGObt58c2j+8D5QxCQdfyb
0x9Yb4RMjXGLXA41oEMLXSsGXlvHnSFcxk5JO5lgwnv1Nn2sbNTZVmeHUcBzYxRs
JxB55yja1+SwEVz/Esjl402oalk5SkjGA09uVSuYPsORqskaY8pAcQHIoG2HnlGi
QbPJTt8f5ipQ09HLAXnrlY6ftcoSUrTQD4ZEAnfQQtO74GC7p08OyQyqPnoLTpzA
LH4jXWSiMKJKkhh9Kj4dH/MhCB1VTPVT4LQ+/MghHqrt93/hkhRbjQpSOEcr0JsR
8RxeqTrJ/63/x9jaBbl9ghBqltxgW9QxK4xA3zGEmPHlu1U2l8xgRIvjHZFMAXui
pmYgY1MSChd+P4hddsvmyEKbEBvkhY7k0RQtx2dydgDw2Z8DrMVKlmZ3mID1GaJg
fYrwbr10NfI8MPCRhepX/DTP5xVN1uiPiAiRippi09VfdwrBWxIDSe5AA1gbzflK
JYv0OHpUewfg3px1x1L7ZoUNbzErH/MMgrVYZznXJGY04yL9fWyy36C3yOwksq5E
cfOFXki7sUf3Fezkesv2Q0rjgtaf7uvt7m7YT/tAWVNe8N1vxXumRrPfuLCsH0UZ
E9n4Ppb3HwCvLn/Y8Q1RwsyQDtBupkX/JopIaMLBU9eDSTxsCfKdN/y10wS3WO0V
njqDNJrurqCutVDvG+BWY70L+C5sFQ0m8yO6JNYTcvMxUdem+1uV6eyNmPy3eK7g
d/Z04sQB2h7j8yMWCFrW1EMkyywShIU58iZE3TytS2BUXCMi0n2jGZajQ9wccDe8
o3Zso7Io0calxN7IIgIhRH5p+xgsUHt8I2IKOOIqFVIQqNgIlmbES0joG9SOamur
/4ZkqwSkkWA9tAbbopJQacxQjrL0gVLUiUanXMam3ZFcxw1BITq14he2XbMvwfYk
rdmE+N3cQg4F6wrmQj57wYigASpV8KTM88clEMuILkh54frcnRPc3ijT2ZXPIWHd
Si3TfPJV2NCDavwBtw9lBqrOqe8zV54ltHdIHTVM4DIJFF1/xnUwdlaf+ms+IkA4
foXqb96KbX8GAWuJoT7X36T8kP74V2wPt0NbUV6cslthqVIoNxfj8GLeTNNUX8Ak
ErdFuN8hXVnoUL5Mzc/G+kRdUL1Wmqq1sUKKZRLIiyEfVheyh2qI2ib06rq3pKp/
f/l6xakSWxeXO72+thqBbo7fVcAAzrm5kTRK8JJESqOyn1whniyctgJN8wH+Zw7N
CRdwFoO4l9CM6qy+nnA9P/GpLFNf3D4Iv93g4+XDiHOP01vDr/3waiDRHBHAJWwi
jHNLgI6E+jcxZalBKiPbz+9w0tBDr2o6ensCo/VS7YBtVCkSXa21bvSlZSnjkJsy
ZhIsSkzAuUOvJdj8xy1/4pTeLS0g2JW0iLussxqVS3F3p1WTBUuIMkUOANHLVdEf
LWFdw2AS4w4lcNyAP7V8OWcu1Rn2fBBk+zVChO+0jVMggreclIYePh6T07I3Jdg7
pZnraUSjfgFZZ8oZTp2t9UctpM1JDzLXgDBQlgk/LACvtHnhcxTnxHcttdV0S+sz
/4noKZlvHeIKnJwf6RCRbmrD115BkAjHcxuZYvdDur88XnBRqrFCDRE95HCRTrK0
FIeoc9UXJVkohvabcDzdEawUu+LbN/KJ+lLidv6Eq3/AM1lLRFwA4Ej37uB6ZDVM
apgqWxeQRYYWOCYz6FRnIfmNWKOm7/Wxl4d+GLV+VCsf3jZ7bbZ7qhlwXXBocvSA
OvoJ3G22jHE1ABU+z+N8qPV9z6p6acrrb3zNTYmy2f03oNiQiCXqSZn4KhD3MaM4
VsiJNqDDG/x2imcb2DrcmpfWXaPLSout/HEQ76uy7GspNbfQLsCxMVYMEGTAq9wF
WLoSArr6v2j7TJpS5i25dcBpaLGVVLXIOTznPPTpFB4CQIq6Ltmg/zjR2SFelCT7
CW62IggV7OE6/E5ZjLlzjzFxrH/gawVLgWicowvpYaGv7SGISKJKdDkk2EbhUREm
1JgKjyy3orfMzqphfIYXDSd8kYts00mIxEoCe1CCUV67iHYCZ35tIoHO3SY4xkLA
JFemaixDqoZ4/DekSkqEjI6jish2epck+yT5NTBzohJN2k4Ms9gE5azxXSJyu4x+
Aijqg8j8abse6Ykpc3YTjh/2uKwpHLkFY+Gza3YeK/Q7F2RkLZ0zyvg8fMbn2nvR
dHBQlQ39ZYv5RCZzkTV/Gp/dmeElGoJ32vZiNt4dLFVyxsWyRWwWq0Z41OiclIOZ
qk0T29OHfeAHwiPXQILQJ+3BFbg/LdJKb3Z/iQDOnQa16g4md7pndpbouCEPvDpy
XLp0FOoKyTHe5qB98CGyhREVKZV3EsNzJmaHm6gvmtcdUaA+O7nLCNMXy0wuqMu7
HzRqf5/gPlpzBkOZJe+HPUjLAKvQ80VvWJicFz1Fhc+kJevmYmT+qJETkBguiS21
z/TN/7KtdMp+9L1n40aBv00tjjIr6m6HfdD4QDnsRAvh+mJNL+dP8XSoHti9cp1k
8Wci0J1PWmQL7iTH389qewx56WxFiJFo+aPOHnMOTkiCohBhpJal4d3aVmGtomBU
urTso4PCPo6w/M8muDbTJizLFMechKSoAO/QgwonDjt/bpbyUMRTtZAYUwXPFEoN
wM7Yo14gsrupR7xnWC/nADGJuy59MK/aIQRdxXp4Y67iMJCVcZf5N+7Xv0+gpH2J
2l6fonyJNWLH0CV8QzMUhoaMgumad4pIwcN98Mfb/B7ZKs63335CkhmC1s3KWDGO
e9O1cxb6JiKdWpB4hQ52Hp2w5EauWC/uRKFSzDcvL5HlncNhQpeXv6201eC3ZNBV
uQdwxQydh/3VPAMyDEAbvvaNJ6ZwvJAQl8dcZXqxx3a7GZkAmLBs73Z6IAhslYTd
l12PUavyta4FcZAxbJ7Sp1lXws6iAjgAMVolbBQpykFznnB8MMUNu7uCQ0UN5GBU
kyB1yfg6k/4/X8Xn15v0MCOyhJLBnpZGa0P71k4ZBka9N+GlFRIpBADKTVuRnuBx
fGFSEvIye/Jl0DtVp7cU+GpIDymP9FA+My25eUqSks4/mRAiQupF2akD8jA3CSF7
IpTQHTKT1RH6od8UXvG9X9TK2oI36aUQI2SehdZtSGNyiMq/pmMEOWPWzbOuB3hE
4bo1kQYXIB0QOY8dXFmZlpW0g4ecXbhIqmdyBKcsesUCyh57VB60ebYDAAsSF+f1
9cqwsEvwVAHdUhw6mONg1mMl5mBnwmKUGdl3UUm3lRNuhDor7ZUn+Eq3QcKnOy8M
eWNNUFaU7DlG1c/XBH1Z0qzWmxhU5PreNkudA1NRQBxiw0OjY1QxWfXee3HQJuml
ADFSB1sMtPWc/Pq4+HIyvQyZGrgiIvhHRjoMl1V9BwlVakiL5Jm0+ftQbCPx2zmf
k5xm752XRqlBVSkECDiahw1T/eHWEv6BpMO/NK1j20yzLuOATM+YmqWrjZelfk3o
VF7sRJcEyoqmAayclZv/H+Ww6uvteJKNUp2jL4omCsQpnYLi5qRMG2C8zDBiHHt2
H+KOehIJf/n8PLbUl4oyYWzWYAvQyb4mK66fD91JXr37mYiGWQ/jQNew6SKm5Eam
aJmTaGDN3e8p3ekMloj/IF/KLBj/IPlb6wEN/bAqfBSrf5oSVCTK/VZNSLcL6q5I
QsOQ8pOs532bROPeYlyzsHc8Q5K88LcDTQw0R4ArJ59YWz5FzyYpNFFdklU9r8L2
cDuk6+HUJo7VAOxOWzhrZYkH6/leUDllbrbswDTTGHqfUGcTeNAsI4q78W8VCwZY
i03dmeTqvu23/UlG5qR0VdMcyfrwP80wd75P1GhWx2wIa1tHfajUtC1NktQwx0oQ
pwNZe03xXVPH2V2OhhaOhCXQv91E3sObeYAN50lZRmAF0GCAsABAxb3DT15gCVSG
AH4n0w3PqdhjzypZIBHKFALZyO7rQzpcMS0UY/ZUNsKvI4wMlrVyaaH2szbSmlIs
LBi10sySKt9Q7V5mPV0F9kazlkYCFIZ+WO6drpViqnoTh/L4en9jw7arRgEaYcpq
e1bejziPw5118ZpbdGLu+X6fzRcCcSYxq21nvv70iJ085Tcb7G3whi++aFotL2tB
WdCEv4bfMcRpv5kTV/OACwp+RrRJ1X2Tc02ZCjXXO9fBvdrX85sGAH7W1Dzh1fkn
JGARnyGIh+dPnysPXX3YhifxdGnQfMmPEvH59QamC0UXxe0TMw2Z5jZvOBwAG7nH
SAqGpCuqahmuN5ERko5yiOoSXWm2i0CQ2EB1N8pQcGi3IdFVkREkrKLKlWR9dMX2
8jy6L27QcjnKwkV0rKkGVfqdl7O5Fpy9UCqRFDSjPE6bjqJskTSAYfDjq2tgYanb
NNMu/W0mhzL7qHPrmQ5B63iVZ2oOuXOsRWjip032PPC+EYyx7aJ0n/MunmHgp7Ml
Zs3wFzRBb+mtgLPE9VkJnLtBnS9Ba9bPFO8Qor+a2LchUHSPA9YLBsiaA2dqOgJx
L9al9NyD7oPA0uXWZFX/8wSzUimqcSv/ex0LBAS+eF0lvBBRNE7MKROp8Me0gJVp
7VHI484ODU6kTAivwKHX8ZhUfuCZDbiOZGH3T/93L1aH4f/RGeI68Z8U3QPy5Itp
O5jmlXpBGQEju9q934PdDqAtFyRIqKo6HuDmENOzgHyHl7GKsZ9xF+DVms4mMtJi
Yyr0D0k2ewSk8h38MyyIxu30ovduV2ej5Da880TLv3D0T33ZDjaX7btKsmz/CGwM
TLrb8v7G+R/71EugjVvardbENdt2uy/l0wHaDpbwDhoaZrsv0mDgKTqXnEMdyoEz
/Vy+HgVbJeU+95alIEPn4IzHi8RDxfIGDeAeQRxuhwcOCQt4GWQdH2Z2N/VwM1EK
DQquxwyCyit0Ukbp1Mj9A1/DhLglZ8RLpPUGAMf1xhu4SITK/2sYd3wPGIefSA2u
vYhwI8VGABxCWnzT93szyVl7lqdd8neKqPmfstQLtkgkCtLsOA4CPTF6zZ3A7JL7
X4kVMUb5QfBeV0GI19fzDdevtJv8olZwhlX2lVpGsMJ3I3DK9KdI7N8iaOyeoEry
pc9AKuDj/3+k4pENNZCISdlzmcQhw60OxC75ojZex0rur7ZmQCSUY1bKGQZ/va9w
v9oR6jGhoUnqpJ2rJXJGLbXrxEuzJo1Vj85yb3cZZYN3g9LIqDNtCATF/qvYaRhn
2vrCVH7M32y6AGuORPr893ul9jmHFwo8zdXyZQIMIshM+CdP8pGEIAfw+KP1JKE0
TUjIU4w64+0EHPcE5+TSNSIqLTQF2LCO8jrtME/1+GqExIKytIxUhpw4fodKd82j
0PNSZZhZ/q7u24+yc+xcCnApgYjzcrIHdyB4jn2kXonTlrYzEhy3hnNRtrCNtKyI
5LoJ1G+jQsnoezDQm2IkwV+LqqZ7BCh1xLWOyGhXWFPPtyuqnkzK0Sf0k3edTuHk
cW8EoF3lFyA4y3NjZP3pVpGnEbdkhPHsLIBng5uJ3RqTW1MHf1J3AoXqNYZ9XYYm
o9lEH18TgqPVAMC0aNMNPTmzybE7nQwR4eHqYef8GSkfWM3n9jw/ej749GNRuN44
Tg2wWAQ0+9+r/b2dVQqONvz96QJetaA16uT+SA4f9UcdrAPCXV8uKGiG0qHOuoKC
9bG4eJ+QAT64i44GN95fF3DsapRdmhg09dmBCjLCFQWdocQC5LnOxbmgBjSVfWrR
eQWMXs4PJon2SheguZtqDoPs+PZmoaK4+yeu2HXXlEMDaO8nmpLupWweJuaznRsZ
suMP85r83vGzQn/+Fsmd/gqXYBVc1KNAgwK86qlwoXPxj8CC2+5byh6S4VE5Rs+6
Ob4tnDNHnO4U+BwJfpZjcniuworDmTepKDGqf6VPTUvcs+mdq1gD7O/q5h0rpwMR
HM3KaWp70ygQDzVA0ommoKstrhKpj6QSsS2+IOZGHFYx7V+obKkkqbKliIiDrTiq
SFTrwqxORxWtVIImu2YIRVb7tLO8wga3xWBW4WtOZUKxPwFwVacjK/o5R8iv4ft6
cX83CLasHHwYmLhN4l8HZzJ0zD2MVan+mhEXYVSdp3c4xC6KqDyqEelmuj+atXLW
lUxm09lIbO9aYNoIsRCWVfnYn0nKUIBN3+TbrMB4FpOnyXwPzpDaUACsAWlq1qvB
XAhhUgRCJDVh5Hc44FTin9blLNsa7fX7KDMYxvkLvjaihI0xb9OURV0VFbRvVbfG
mXe0Eo/vDQIsqYUhxzb+pTvIvZAD0jbFXQHylSa6h7PXLPy7MpE89fRaI0GR7waa
uQnevxCED6IQNt0C01gWcpk8dKCV+z6jNpPJ2Enx1m2JijlspiPuUqselOzDVV22
RIhwvlvnXTDOJy5liDWIJBF+vcvJvBlMV4XvukFeV0rKqhcM4Ouu1MczLlSWf8EI
SF67oS5HKhoCBaHsVCWZ7J/hUuQsuM1qRs3Q2FvxX3weme2kvKnZBD9ip1cDDk2w
/ONo6ERl5xcBuspiZi2Q31D4FwH1bfwPMvSbAm7videlMiNVspeNjqCIJ9eJFY4a
51I15mtrE+/vcthdyOltDGFQIs30AO7I2H6EthJt1OBWblG61QWh4GcZ91tadxj1
UtPtOfdbt03W840eONK2ZkEwjyyhyPNqr4ivhqab3G33X3ETP5TJ7NWRQaehCWG3
2409feruj6hMC+6ztUHNrf0HtDljUKxBmbJOekpOJ2r53yY3QFr1eb3fI4neyEzQ
TgzTHUDkF92hRlRjm9YgGjvCWFvZtznM+uHdF6VMuITzknEF6pNQ5UYBLMC3LyRP
+9BQ9+nPiJtYpDRTRFIUT1SGKrxRo/prdzYN1l6vzrrDO4tDpVnA5FhrNgHTQHaZ
fJ6CRU5iq65dTI5jHc3l1+Ur1xVaBNdrY980USj2iL3L1l2QGnUaJ+yJFzt1Imfc
KaUpVAGPCPU08g1+10xAEhGLBcATT3U+CfPtGVw6ahuIA288XC37A9S/BlA07I9c
Rtl+KbSWuabRiKuAfnqazBbkFP5PVHPuEY0m6sdu/miyI2BosL5A73rv8theVWqs
YF/lftpYNX9570pW427wxQTFGxlUDCQII27iG6IagdR0QYYZcf/1/e0A0tVP1DKJ
JrfJJ2rhhmM6+4QPZqsKUA/8s2hiEBO+bS/LDeZkgcGMUweSmKBgB/e9sFpLEwfB
Y/VBQeaw52AgwlMmV4H7wgIEWIO35e5Py5sEIlXEoH2MTBuIK2HYQWfawzmx1C/N
yOR4l70fi9jW5kanu44b1KK9ikElAuKawM2N0p9/OCQQNqql0QwX+kyOkLpnNlwd
mkb4DQWq0oVwDgAVnaUO3LOM1EBRToUywPcKBMtBJOCBdjtIlXUHFYNbWBqXb+Yc
+/OEuKX7CXf3Yd+OZr6vWz86t3RR59+ivSpQJqZowh/NC3T07KrbvQR+MTV7i33L
ZafnbfEHCtOoOp5jY6QGoOZSnQyTy2e01g07ex2SNQV0uwJc+bRN1eFTEsZZXiaS
7LaYlS0M0wnqbhLuIu9De588cKs37D8L4ma96cPecRvYkOpYIAxBI3UW0uZ1IiwD
mqI36GhoFX7sG34YDDTjMImM9864PApmqI12JSeY7+PXjF7Pqg6oJinriihH5DbJ
oQ+2RYo9DnkZ1gfexW7YuS3bhOJGDYQBMgPg7U5/TyOrmR43DjK63w/tYXNg0mOI
1J7MgHcN5Tx5Z37Zu5iNXmZpUyRVJrhVg7hwQt/+OCXwaq/BYWFRdk/eShL7DkjW
FrbZ/UzkU9JoKx7XKMT44wkF+cgcU4NjyT4LTBWyIMlRXyTgpVJajmhTRu+npPYA
ivA0inXkbCO/Gr5sHc0ulkuUPYw6exq7a3gRhDQCok+lM1PsnWMXkWPIjwB8f1OQ
qi7XV7siaCAcRPk7qswTc6E1aD4ef2jzbs8ezFQcbP089PbRNKk40MgyKmEwMLzy
dT+SRstJdQJBSVWFj+3+hyGBV4+Ici7JPaLCZlvEOUcswSQvlcAtN7HetfnemIYF
p2eioDIxZnQoKw20qxFcZOKJ3/lusUkyudk0FamJmZwfGcPrZVg5VCSPS+m/KaNQ
lxklWu2eaRVFvMrJo7FMhXk6t7qYmI3k5/Ut/Z4Q86msdbLSzTINH0BhJHI/2Qda
7umqkJwu9vF1VjO7g759qmrd4oATWB30Zqtc4KjWJWXK/JDL6Xy0G1tB2hhtArc3
Lq+R8r5Aua8GC0j61euDDxPkpP1MKuf8jU7iXkQYtxjQGR+j0dDDGslRTK2Pp18L
qQYleKCL5vVCfv8QoiXXL+IkxyNY+/jA/Kvc4i1mS5YfTuZDripDVB+0bq5j3eLv
AjWbZlKu46Hi8CYxjG0HWV8DhD9Pns5P8UK0lYZxL1FroiaUhvPmgU75RrEgRApZ
O84EwrEbLTckPyvwHBAAtnyUIqXSwkZvCn+pawMPX4F1TOmSUCCnnPyWcNKx2HUf
r+SAmzs/y55k+r5DQO+y46lPYBaadMDG/BKLNIFz5vXwoVPHkjYBGtpfFH1Vy4oM
tY6p7WBX926lrnBYD6Tqcw+afNtxHB8foTSCE8M0EByTQvncCThAGmcycRasCj3a
UQRUHog7ziwfvZfLW4xN0hT4kbVu+TlB2+Pb3gH0aQqbunsy0JNEh0fRzDzeoV0h
H5SC4D/vYjzEHZCxZQgUNKkQZ5gp+rJf2wuQOtYZFjEU/5pBDVUL/VMqEYlHQxUg
ArYaQgVfltpkAazCFdLjhPw9Z6qnD4O4EsUvjANtl5ebCUKSSWTh54xZEXENWySn
oGW7g6HhU0t9cBvbSsYNJz630HxHmrLPbUzsCqyUMs0px6MjLtFGooCtMUWneM/I
76oEOqVosCS8zrMK8VogMEgIzFBY4ivpsN4VEM6TJ0aHZF87JgzeECEgPIPXDqMZ
0QD8S52itIREwSNU4wW0eURBMsiM4FZ1K4t+rWgQJj2Cvae+qSU3eX8/yyiwYhEF
JuUtGtoULxx1TmTCMkGtUEMUKlGd6oi/RdIEiBwLJMmf8jBMDXGkqjFYMn7qNaBY
bcDliJY8dHjnK8I4j9zdhTens+UriqWvK8o5BU4wSlYmzVAhP5O5TZocGq5dl8U6
yQMsGX/7qotMsq2REktUvOz4PVA5uKhCyHvZ+TCVWvd3N00a8HEN30/ItKov5We8
UOZuLTPe/wG+cq30CahqMLedto3aG0nbZGYJkBoX7D7M78meS1b0VLqBGgzoWj9z
BxoBZhgxN5zxm9zlnNj6OIhfi4T8Rq/RZQHKi8/KVMmLmL2fcGW/fIZ9ZAFwY6cc
b7Toof1438gWw6QYUhX5qVIq+BdnaCFeGqsCVQzaODFyiMAosKRlY4f51+MQR6KS
76tGW+aPq/nGPGRBbE4rWDN4ANYGTKfK26/YumOeMA42Yi4sD6nG/6BOxDEbGtrT
gbpN7f1gp7vi7w6UMXZ3vyybivhTlwtXhXPkEAYsfm3IIgnMlztaFaz5SmS+bTzH
JeveEouXcnRvd0XLKS5fm6XHp9RgtBgR5XKAqqDTyVhOeuE29BzrXwqC/NNnh8A0
g4PWVxFQiZJXAhknNTV4kI+xYu9OzImkURlw7/OYEj83Mpak9fpV1pomSS6Oy6DA
P3HWQ5ovtmBJ3DXHxWFXaibvzLbLWyma6eNCzlaAS2S6zpbgkec458zkT85upomh
jpKLBYitgiKJGn4fuwOm4xkwr/cA1uSG19BLAOvPATB/l8KmaU0Uq7G0FMMQnBov
rdeACpN60XFi/UFdz9KrZHmOlV8vnnZclzNsxD9GQ0kOBVByQlzVFidDS5KU7D2z
QKe2EUlMDd1c6vNr2p9oERxd2v0dZhVJLq5xUXIUOA1Q2PyyoQmWFSxz6l4DUXcg
/XGPViGc+AiZhoF9rHkvK5rGpVRITwCm5czcQk2wfmUSWtL3odA0+53yzuXyj8PQ
iqd0orHMVmf3pyE3XeskRWAqrgojdEB3QYRho0quvpP/xxNvFeWsQvow8CEaPHin
cxdMU4QcaygrXvapUWodyGpLxav7doHKN0iHhgraoTnBUusKHOvy6oQ+l+2fQoOz
Swu8U53MkHmWCoe85PYiv7SA29fYbKqP/VW5f2f2FALT8QJhgvF4eoKneWgi9oA+
BlMc00MfWuA04Ieo2pdZ8IY3ideDeas2Vls4lMl3fpg290kqH649o6KlQg3w0Y0K
wzJB6qs0iiNv+Tuw7hJTjU0/33dL8ICIRIaHTd2qANWmStJnDD3UbT8SUmL7KOjy
YIM18naIdg3poWCytMyZ2GaHZznvqmmUnMehNDp7aS6fHZ5jOE5hwyO1kkOenFFH
/qgdwO36z0eYi/XPZ5lW1VU51HyHJWWoai6eoTAhnWyWWUZeAaZwbuZgIKy4AqzQ
JaIuLzgARq8HxhjzrvVeWct7p8b/cRUxQPqgVNppKKiE1dQELTb/TTF2c5q3vUSp
9Y6tZoPsy1Y5rxqC+1n6HeeEM5e+3yWJqWmYifKB4zsvQMOyVjQA/gcceeEDyVrp
9WC4HtWqWL53cd2OYULOMAz0BrnkrNBPP6LqDcvsnffY5rDJjFVFasw9INZ05Awi
kqic4A+aIByixeEFJfK2m+PbV1SoKfEiLWRMHY3aZvclxKXXDa11KIyPS4YmW3ex
B/SBjuBhSm39aGe7aYRbQrZ0ozLg7bE/r+nbMOKbhlQqWp57cFSAVlKD2MCuxMvy
+ig184BiZOF/Kw9rZJtBOdO+9dUQGFJSUAn7kNolfAsOteXN9VS01Hvqnc4oA/KW
j7P/gCzEka884wAUpzIkLiPTvF2SDL23AkGhdFqFcVOOY++d2bnQ/zAdnvU/J+dI
owrhWQ/APaI76y35iU7W4+SvoxgWEGh4CgXjsXAYayTwftDtNyRP/9ES4p9QR6Ra
p6QzX+tPpJ5WBTAj7nNatIqCQShVNGOF848FLQDHggi+TORfam0ebJmXiz/AurMP
0PV2yy/FomvzHgpDeuSRNyszNa3OILkBpyK0cnpT102wAxAsaYcxFZhvR8xipKMK
Krdi5aDqqlmBsOQBbqXcT2whqiEWneBl+A/w5MRlZduKumgxkcOmdb+4F2eenU+E
eF5HrlkUZy2tBaH5p+PkI356IpXyofzML2UDjhodHrx0uH+/OQoEbS16arZKemFP
9mtosJ67mWyiRtendBDOUFnaFHFa3jpRgJ/v7R+nzaMtCeSXF06t6/PzltEzqhcG
HYSJgSoA+2rDSvzGj17QcMaSomWb5KByXbCHK1GFFPJJEJt4icl/bes0gyOpNyMN
Pi8i+7rigFT2EGw63+COIT9UJcYoVvp9XBs+bupdrV4MVZmJn6p5iIYZ+rdslvE4
IAszoJcU4nebbopcm/3P2VWChmBYl8cEz1lVN5h9g+j6R177tWHamZcLaKjyEXuK
u66Qo+gr4a1FjBKN8/oyTEp95uc4kyypVrYtx19U/iYGck8IOcC8zR9gTjqPsV25
Q27bvdQ8Wspx0tz3r5WCnOMz7F9X8892yE9N+sWfbLs0N3pOcIr5POie1kaeSyw3
TPwXzKrkhzGQVNch+odaR6VpV7AyWZ/XRxCRcXlTeMBOZdcOipLlCoLQUtCrGqKU
iwpy9DqIiwJ//EsrIWA0GxeIAUGGd9mVsqM00x4rPxVLCyaNlcYcwRyEc/DbCPdw
4qe1CimH2eP6Osa0IGOkREK1XakeI8DfkjHidfN7joQmLO0Z/qB+6G1ayXZqYDSA
cLbckaOFmVWBvMpPwG87ZRlZClAPxLuts3fENclD0KoyG+Xmut8WviH3eZMhlUGj
MmIyVthigpvpZa1I8jieGmrmvhhj1CPvp4pGH7JP586h+pPz3igEoAC2+Z+sUIJ2
GI9099jkC2bIIinKf7aeKo2FKpIsUQ22GuCCo6OW9580opNj29dlpo96W7ukXoxE
oLZ6QFJh1utk2FdZ88pAWpnCUtcvc/iI17rq7aB9hL/jjWkw08Upql3b6Ic7L7+t
vvkoW+0QSYfnKbqSwnjUt8+YYSRC5eeS8CHUZHxMiVJaPitoeQJyhQJ129rToXLd
a1vZugAViQmNusfsRqzf9QZlPUVRP6EWE9Knu0gN/rPqkosByNp/1e9E5kLMg9vx
pe6RWYOBKDO/cNmk284IWjUG3m5QHPqVgo2jSZDJA479L6RvjYM5wMPmoz5cBaS6
WWRdvHLDWVoeE9MyJRQjCcjgzZgEFZI6/HxS9wTbMexJRpvB6E/GV1GE59xYDdQ/
Aip9Xzpn3dnEHD6Bm8Z0xAnHoIkNaalddsICeP04Q+gSesxaHP2n5QQdj42GhvlW
sdY4eSlm4e9hX+JVyP1NzGhAvoSWA+BjQPH+yG81/o1Q/pqZo0IYibiD1grSQScK
FIF769LoAk/6PGPb6JTiSfWLKhy6HFBzQwxVsYlnMNE+A2sM1HyTHbR5iacEBgUR
XEl807Yv0zUJ2icde8rgwCcFqE+OAiAsRuXrIBwhXyRH5zIeskiviLHrPzPDbaBn
h1IEe+3n5UR5oVJ7ebpSV362i3al9tcJ6TD7rwSrVfiVDVJ69YvNAGErX3eIwxCP
xqKEicGuxedrT6VZ8YhLnm1OuS5IA9w7KPHZ5agHoc+wMJqNQUQBOxzchGlTXRGO
oQSr6OKy24JmAsOD+H0jUwDbDo/rpBgic/OsTC7gB6koQKKDidavkh9N2zmQUYim
FeGrVYZ/yJGy17+o65yyTSMqnfE/2Ba6tphzMbubVDx2+xdBIF7XQ3CiGUL5Y/EN
7JDitaxir04rjERTwPt6Od6ClfDRUJ/XJQFTHmajKybhrJtSA5SzEAoiIHnmaENN
LUN2nXhyHMliPdOV9jcpuf580hEnlK4qYyYuhqc/Yo/o+JSL77IHkdncZyPG6m72
FVnvTlHpeaWoBfNDwpxfsiRQraG4fGeP3W13yOKDbFycbVXE+1J6zQmku5yZTwEN
RrGMyA+4KtpsPIuOWVsBu0dMc0/g59otDpDLgxG8xc6IVBF+dXHT7XKIaKfNKYL8
CIJDateheJaAE08NM05m2zBf6A8W7BZwGCu10vYqeZeYbtgh+6vcNTJdKzEMRq3G
xZM2TzPBvXlUGt+p97EENTdo/OUMxksPnT2PqP3hBAzJwHanQhC4xatlUAGV7+Xl
FjSk0/OT8wLnfbHOPfDdTr8v8O0iiKjWkSYbuR3LerSdKllqMReYC7OjWo23WDsT
8dsHlneN1l2jTCSWcKLv2HeJk5JSNgNxsDh8Q9fpOPocB3MuPlgl4IE4sQYmYCLr
9eiWKvaDsxOaPH1Pu4gNxIsNZgYh5h3fTwSsFytpWhXNlFp6ZgXfeQQEmfCuTTqH
qghQ9rNfOMx4Qs/j+/DsYotrcnUEDfMCsYBgfvFZbhg5OL06EgKBexzJ9xiItVz5
AqRtMpNrLeK/T+YFv5hnVSwSe4LfEdq4cSellI4aLY5rcUpirOSmLCLonK+hs5qP
JluSI5s1vA6DLIoQYWB3weyEOQDAnBJBV9MBIYJOpUZHWgtCIL5m0c10F9c/GsfL
q0VndW58oVFFvj+6SJCxPn4SyTYBmUMIDZWBNOBB/XDCM4peZeqsyPrsssLC5h1P
bm1eBhFnuJBOU0TrY1EMEpp0eQ/wjx0kqXqpK+pQIZl0iMc50NZDO17nAGMZ+gwg
equ3MvG7VDMVRU9+WJF0LRyN57QREedoVLZCgF47Sg2P1zGI/s4gs/V3snzr6BuT
wJSl/u4P6B9LVD8GsVdfNFb87E0ilM/lrn3PIRsgMPBsTzlSLzR67y1+BL4BJCwL
OcxfCLq3XRLPb+LE12qqAzcCFt4CdlhviOlGwl9kw6c02yeg94jg1Rshb5GhoVfj
6hU/CyGmpCjBBGQtiCp78BSZkWLB1TI14TLIJYBVyoSlyki6apTn853qZ/F8SCrp
MAjJ8F2TNU1R/mWLc3sfYHLrDkqUWu/CW2y2Nxd4bLZ0Uw/uDZc/1W4LiDYqfe2c
Jw5cnl4Nex8apKLMu2VXWOwvZuPnn6EB4IFJmQs0x1X7tRMgQmf4/QNQFRPK6FT0
2IAjY69/SN997Hgh5dydpFamfKWQ0qurl6304Vwc0TroshaMpYxEVQNPEHDdbaeW
UvhGsP5ShJpfNqh2O+njIOTzjJ4842DgKwCw7ZMJm0O/u1XE/WPiYEVcAyL1YLSr
pen+GibNPKfnMznC8llNIW7qvdSO5wULfUVFcavfJaG+EYtkDd5LZBnJSwTqlbEl
QJR8C8pekOmG6h7qhm1RGs7QvyyHXCHX9wwCFmFXbBezD2p5rRN3VAoDUf+1nZPU
lT36FTHG541irBEXkFwXA4+jEEZcOzPlDGv8l46SqvN7O7vw6M9J6UFnCRnmSKFu
5Fd4UpmiTqK4pTuVSQ5Q4/sT8emc5JQLNRIsu4ub8MC596bEufuF3fdQTK+yseqK
Xx7GgGwIM9NiVJX9HoWGeQ8LMmCIvE8Li1OMc3ufajz2RX5jlnFj7bwzLsx/u0W9
T8ttYnswJOhfJY9sxRHM5gRmZx93IlNtLe3eKRwUS6r3aik0WuU2baeSQDs3aZyu
lGb9aC8IFelNTeL2c3xTSenD6qX1n6smFE/CMxlZi1ERVzeCFwoOS+oOatpgMRuB
D8JUE5FmD5loeP9loidQpaW+JIRAqf+HRV/Y8RPuItuTsrq5i4DLakBQti7gWywf
+T5U+dh45EJL7L+pUastTydcnm2VE5GYdr2UHSTxclmkSVid/lFbzIMqTkMvWkbK
JWfZJFmfFS29E+QZkAui/NTvp5chaJf/bKCBWZBr5fSzh+xh7cugcu8kX2gP1ago
G0IaUm+uyD4uj1jO/4WbaY79xIdK4cQaApPLkKnVwFnKXDBtp6eKlfZm/Grs2oDe
E8yZNdh5lFw+ps1FKOPo77ILD3MpACdJiELKHvFGgGzzQy3zwOYJUmind+ZYcfB8
ylgQbjKuyjd3udOY5DIpSSxxYOQilFE5muKCwo6ljoVBUu+fcN3r4yQid+bOEl/k
voHCoH+3IFvLV6XK+Oqz+wvNgjmBmA5xI8XBgEQc4llNr236TKAnI093nhwA1Xdj
5A442+fntYw5dlIXm6z635rJOmuTrgtQRWSXa0ro6pW1EkS3bux7yeSADLoCN32l
dnix7+8xW7Dzlc7QvSm6Tp3ND4JKr9pF1hrXqS/pvHLdVKfOdcY282ctDxgWsXxR
8v19Qd0Pjm4VpyVJi4M24eMHdI6P2ik3rFDlRTTrXP1xWBS8ux8N9dXD/FatEv5Q
3yAY2wI7hJr00SrphkUW3F/5kdJR6z7K9tsPLKRcGB+yO2kvKQ6IJn2mgc/fhqHa
MHBYbd6z/hJ+Iduy2Q3IEdcGJNruKLF0giboF2bHOm7l8qoZBc8ZLh5xhaGpW+8u
omD6/wAY+yrFvWFkUoNHTVCnGF6JDfHg6KP6wOOTZ5Zsn/OHspAbJ9H6arn0Rdc6
eBLm3sVySq+JvvLV+2AzVk31FwJ/WMQ2v+/Fuuqnp1lposo9XHSUTw91B8grkSCu
wd35D+TXkdvz9HPHr++YiaWUxsqlQ82u3NOxoz/ISIWvtDWNeuGxxZkQlLLllxHH
+GYEDBn4hF9ANgk7Mg/p5z5euluJJ5DvLzF3zikL2kwWNnWHwzwY+fWfr/aUy8CF
O6jJ1QC4kSV2HwAd2O01Qgz6sjdY4174omfkOviQRLvdsW99Zlf84JCPQ/ra+0IJ
ZitnWAjHbsxzLuDnLXEvBG3MDP7A70cwWWCFmo4Uhhzejrb3bRdM6rlj9gCsPOG4
m3eC5P3k2n43ocGLSpWvPkLuA2rO4Nnn18YFkEaytva2jmHUAIDQ2SmlzQIhO4F/
Y3SpRi33MoJtCHGE0tHO5saUcAiJyGiqfJSYm37i6uu5RyIhIiUIE8I4NV2Td5rP
YkG0oInhigdGI/9ownACRvOWAfvLBgvqKsNgGahSG76bKFUuRKoIVOv0IYbui4tt
YJIOx/Sf/k2I3fkYxiyOmbaQicaIVKK+hagWUFNuII4stUDnA/2AGs5CxbAiY7eR
CPTxo9iO+Xg/X82xi9O8OaunZQw3b9eAXo6+PeJBh9nWV0xfQNihYlrPGO6fvPaj
z2NCGJVRe9tbK1a5pacADhaOOR7ESGxOyVVtG3UB2R1GOuH6ge2hmxvrA9zkmEuw
qFBIiJdeR3SkHb++VMWU6HOj86aOtTjZzLXlzaKPotIC8goxCO38Dzppd3HEo0pO
B5JRYzlOU2WCxSA62ykn1LABp0Cczvhv+IjcvBaBZeNfCueNnDBJjE+mu0XZ/VBI
3KDqEBWPSz26/lBYxbTf9XiVfNIyG6EkJj4lPskJAEugkRQz17me0Rcb5TLWWY54
mnw8zgA1LRxvJBSrmCOy3vVS4gvxikQhoASRPDDxOnNLi9NrwWDRG13i7YIWl4TR
PekFO7ZZaTdnc8qo60LjvfpwAoE7h4BE9s/xRM4fRulguEa+5jcQ2UwUuP3x53we
xw+8qWawBM6EIlLVkpkcTTgXwcEfRNQJyKvvXsZd2XEg9sdPndY0Vwrm3Ja66k5m
OouYhIqP9mDhIQS3C95crD2TGqrxj8nb9Ou4VCWuo93QYOdHxXzqMOOub/q54e5W
xERv1XgAleYP29vF7XtKzqZOUaerkN3pHec8aK8w5tPSyKl6sBXCo2SyLidhTd+f
ex6srApFEaGj8kgNgB/N7Q+yKVYdwDaDOVLdwuHtDkWwZL94DQBPwkvFN/Y7y3B3
wpfa0PUNStRuWX29CktOXrZ4gStJmer+Cq1Di8/Ph1EiFHO7TSABIbPJaS6SWbBQ
SS9NxFEfImxkK6Ua7mtnLQF4z2WewvBUCbTaD5lTxfjdsfRmSILuBY3iK2TQUycj
rLAh99KAsG1ejVsB3qQfmze5/NcWYqToVdY6boo3e1kLcBo2NN3IR8yxVYS/PYDa
Ab6PignARhkZp2cBoRmRY58EL1oJ85owyV/KZHOesPte9HiJQbC/ExuI8uD6RjU0
B1eCtDrA2et2rCoc9Ayw4ARNvS3UbRPvBGR6mDYbXnv6tToKObZqfNGSIQIVGYGF
Nh/Bd2boG4gsm8UVkvwGFR2tTGxM/akvF4DzbEQd7LDEGDxae8pBHbkWdTKlZt2g
bfKQJT14jnDqMzzgyCPJEepVK+mHRQz6ZnBHN+pkBOsAEo6D/PWg6i+Yawg+HMS1
XQ0BzIgZk43xWEFpBEve2uOEYZHpaeG/rVysiU+/tUjrqoIfmZ7U4zTCedxpkINF
d0PcDQISBywfFecH8KAyTIn1s88jaBRTl/qLKKV1eKkCREpdQlT5jwiVv3jo6vVI
P4i49ApLkTZJ3F6DOhsQ93rnjiFTP6QL+ug6l87zAv14WwzQsjCpJiqcMKAg/PAM
miwHgJlvV107gQ96kPwkBD+A8jPPjk9Udi/xgF6CxgEkJxcBv5juY8y0a5fXRTSI
jG3xylms3LrBzVxXiw35ohNjV3E4t4+iod1E7CSpON9Ah+JzhotI/GGWHEseWnHq
0JBxf9SP+nIV53838LTNj42oAFV6GQxqjMjiUsk0HUccT2BgduidyqOQfidJc+Wf
7X7Wck6ACXdsYaOImsVVlPvMRX05f7DyaRk4zjw9sygj9Tei+XyIgjwhExRK7LEB
CGIBuVFiKBcQ1iEMFYpP++Wl19Y6k4T1ZUN9gMj1D+fh74HKeJFH4LpXhBHlHMsf
hBQOuXRH4PhdLH2XBZS+QYEEU1Gx79IqDodXdotk8DOpDNUwplM40dI3nAXti4+6
m9aR4a7YGtIPpJWb9O0LhBXtHROC5Fwb9+GQpyYcP8VRr7kSV+RzRI9cCPJ3dNB4
lK5Q9pItY/3HBeTLLstyQ4hQ0WBu+NFG7m1vc3EVf5jiRQsuNj+HaemdEvJBaMC7
3gO0wmqqrUYzviLCzWsQuJET8Ksl1v0nCK44MwrL6nnm9a2NvdPTP++8OuPX4BGn
cK5ymSNpR72HsTGzAAULzzA2RtSYPrgHMB6Gu+53WnPAcNQ+5oNfqMR45zpqWvha
d45dssVRHiqN41FhShrONLI3/TKxDzoSDV8KXQdrD+EEFI7JMTsvQtdf3aKnOdVl
k1VS1bTNSIIXcfyaBa6hCnmbV0Hxgcohl7ZmTesNe66mp0f3A0I2gc8AlR1ac5S3
rIAQz5bKAvRiec1SzsIqGIEDD+8e1k/l5uSRFwuXQRWnKuM7OgcvbijWa+/Bv6Lr
INqO9MdMnuTH55gylsuTFB5NnfXmmK5q1+TEawnsVPUtQzebVH4xc/md6NkSMeAK
iC5kA/RXCMnrIPwISGaArN1sB4RiIIomTB5BXt5RM5Ikt8BNiHuTcT9eiJ9lo315
Hxkc6SjmRy4KZyJYV0QMOSR0SeOnP4OHRQO3MLWfxZw61d4lWdr8ggt0rbM6YHLt
LFUiDdzIVCT9i4ZnbISCkF8aHHPdtf3IjC2+1b2qVMaeKvLMDWj5Jf4WTZMPizke
TU+p5GJhBlsxbMakvEML/PDdYolFMn1Gr48I7JlNF2ozM9u2q30nkZAbvSsL48l1
uwkkTBR98mAmYi/NYz49+GN2zzODSLZK6AJynET57lgZaJDnHU4AuLj9zPV/aasu
efYdPkqGOL58qAocKTyqcgMZnHGqkz50esaf3++nAHaXfOHkTY0/vj8L78aWGr+s
6KoBjkYCyvZGdMlO6N2OopWdFKpxfrU1qaKMpjylYWEFp7N2p/WWy0sE2srGN3AL
tTXXh0zEdWfWueFHHjAhdSA1GYghxqxZoXTJWKksiN6CQX1M5emLG8Wzakzsfh7v
8fFIUfWCpcdImT/qpw3/Do7LUM+c9FrFTgCXI+pSorVZGUJUkoYxHqoIc7fTl5sf
jwutHbflayX/9o8pWf/+C5ylS+fSwdWQsnop2bVT+iCtLLVRFFgYvOMZ/068eZ+I
zdU16ZvVvWMR4QZry4WvcHyw4wTsSdJpSrcD/QfhMYxe5yd/k5teTdyJnpNBG9Mr
4FZpt/UKAFRYET5jyFOfThegBIXmo5eXrADf26S44TxF3Uuh2XFVtvFg6UK9O6mX
CYpq8O3GBARnl9elY5Z/kS+hgIrM5VdNqeBCBVdMphFLb0E47mMdPEkCkroYP0rL
HbHUoynh5Wuiy0dhl9IMqKBomptyVLzu3hab0bYIwAh7x4tcXt9Iruj9x2f6F0Kx
2UyWv+E4enk7ldfjEnN5kCeSDegPJzmiQxEDZgAW9Gu1Df81K8Pe5du66hSAVQDC
ufjLu+cLdHCWR7JlEwVR4zmcAwO3zfNpE/pUOYOhym5Y0pn5UjFxuWK8C5iuU9rA
tv5wIP+pURdVc8ZumiPxjuyzSOkg1TSD8sUvk/GDZTRcS4+J+ee2HjFa9Y+zfDn9
anV0/6MYE3PTXLrWyQYx7CegIVX2QWwQen0ODImIvbhTPrjC+PKYrpk88hCWR6uk
J5mnHwgjKRnHTRSU++nTI+b7jtHIDFFVTnxFHoYofNT3HpxkR785jU2uqOKoqnqQ
5pC/socypdQv8jn51wiRCgfA5AO2iKlFj1tyDSLrdQQ9Agyhyd4HalWAZyP6WmWA
ujGC5k+1oa+8Wo4sjbAOEVer+fhCEk94xiCgdg2ltOiJ+GCOvk/upSDbuuNvY0lt
yGRVN+/vE0A0u8Q9ZALYdZDHHrlmm1rxfPD8lCvH5ut4/5LiqVlSUi+9KfVmUt2G
6aI3/Vg1oUfekIfOMZ/Ff+8DUvXI+nRMs817eePZydLiKX3ZhRXFuaAObdfZ3F7/
gwIt831pObK2bJ+a9EpM+GbH/B91OZ8j+0me+fa07yZxLdYIVROzZ6bMuP/MRbzL
dc62oYD+b+LCOW+VrpZ/YA7Z88YzyTZfIJ4rwMiFBsMqLQpp/giZKZUvVDdDWiWq
+eo7lIF6QB3OVXKsxcUm9PqqD1PIn+c/TTYCUxPXYi5jvRhtU1YaVT6VXo1JdaUw
49DbyLCmgICs+dXCpcnPVI2jeFFV+cuZIizh7l1Je7VYpld2f3XXUl0I386esUlI
50bgA+JIJvZSwhvXbjAMRSa0dRnYikALdGGMf42A45GwG2ZqGEMKWgUBoEmgia5Y
YWbyNsSeAv+6MN6zZ1rM69+hbJ4HaznWXbwL5Do2NUK3Ns4ULZdVYTE5V4/RGQbK
n9m5lA9DaNQ7wIltbjJC8QjITBabSurISu3OmI/fEBpEXZuC0+yfGih015bBB0vx
B+qEvjyNwrqwkmEmBMCjoYxdhoavUJSgpKDkgVm2S6sKuGv3ADUnSjWB+hsPKiCZ
tMBTTyPdN/cHFv7Xs33MDeNtEHYo5udGKAfzKEt9KJ5frqa1Me8C6asnCGyzMgej
TbTcqubPgYtTnBUCRkqpC7sIezWjYnzvrj7fxAGg29qpB0021Hazu9rkkFvsHnUz
5mvxEBmINWlLQVuiDjEzzqdPZLEWc+09Sh3bBgrpTPffbCOfmrI7V8ZlV7aqgS8z
OIuthMokQ02xNHHN97X9Km06qTvagTOID2qyydI0IoICjNInFTL+GJbAVhjr0bks
sgvmTGb4bnVs94pS9YpVU6plrFjZLSoD95XjBQVtouC6xb+iklw1g4W+4AIcuAYi
ll5mEU2uzcHWbYtLuMRTetL+tfQQA5O0KOEt8RT04P3LWE+4IlRpcJ5bCuUwCy0Y
6rzcR+L5LuntJRIP7UvzgHkKi9TbxznD8CQqmeuW7RhFBMR6s7knDhbnIcbXPLDs
mHGecCT3/x5nAQwtsw5EZU/cu+3uCQyAMYBJt5RpjsELkpZIRYptxjuqKm+qMApj
RBncFNRZwQYJZTtb4mhKb8NoNcdTEI8QwZY0NdWFFIIQ9mzIM8MB/JFe0j1TdKrH
243e/SDqo/xBWyqcy0IYVlu8sL77PmQNdzCxOqnFeNoUE6VCmipuByGGd1cVa1G7
VMGvMCrxnh2SIz0zbOaSHcPPV46AbIuS3ozthQYsOMwAi2HVgdHHY76hrMIQBPkv
5NYld8kGzSr7hoR95WOmraEW4afnvFyVRVVE1XT2ob9akmxjzk5DbmFVAqbphZma
ay//7thj6N2BwAYQgscSgcEQ9Llksv9WE1CPg96lFP/VVxk5i/i+52mv6br9zKhL
7duPHJy2uGRJQR5MNUV9ImObREyIz6nQEUMdByCanpaSxYhHu9rNZXbF8L0XUIRM
sjuznl8fjjx5l5QRBcQgnk5kqQFlD/L5xlsO/J7/Tey1ca/xkQtpCToDx1JCtmc/
2/5Ck7NwswSGKMBHOVP2NKfUsUoTCl1xAaT1in3g2mwcs04mxy1kXVwL2B2S+mrs
u/qB3qX+prUCTF8pGCaCBP5kjuLwXovh+fVqM5SMxWjeBvkW3P5OYAxKk3zguJwr
N0I19ZBzbC7VByRXYwGpqC6KGzeCF/kDVT0nwuPkfT6f16YRw8cAjLYyoYtvQJfK
hWTf7ZK7sKE3dthC2b2CHRyTYVfQ2Rmf0mdAWahLRO/phiogvKv1eTisF/u+AQEf
tCx0hOfRop3JFnVQvNOJB+F2luz5OGZXK1ya6Mlpux+9Pa+DF5p2VjUeZMh+BnBM
oUMUhQwyhmthj3s3MzdG6ruu188sCYrVzGPqRMQ94TthOBGhsb0EfvaUAaD5rXQA
ff7QhvMdW5jpctHXZs7kxfD1cGKnmIiia2AmDyBRWgIi5eJsFPHT93yZfLJM+xL1
KNEXM7e9bFA4wmqnS7v0d/aXBLxLSo4+thA7PLtls9uLpYDoBRELyN6nlszOKzko
AV/Ucbm2kqp8MridQ9D/duy12tn9h9H4KH8ogAnwnjykXuc409qeFagLb0rA9ZkK
rEM4dikjrWFlH9LTE/S14M09Ly/FqM5o1KoCmYb+qB7b/r1fxhh5RnWldh+0aOJo
SNm+X3OZpA31xTdL0yLEKn8V/Rn86h4woKwGAuditizSnDjI7BTFgmA44I/bi7eu
NvQ/SBvWTFxsbqZt0hfXLR3cACfNp0lzuTIOHN8yf/XriDjZKPEHyE92A7cVH3ad
Y/AKx1yyLMNptVBv7jF81rqaQRgXuWBPY2xFVZK+KlBs4ul7sdPpUWu3W8/JHL3Y
iBMrIyomtvobC7Qsm+0qRE66YULiwJZ3yONZ1gVEjeKxp1w+gsy66PSqaSDiY2QZ
qUPXiq7ShINNTuyQTgbpDqnBkGA9Pyqhdze0/Ve8krm/Pqo5nGgUm/3DS5fGX/4A
IARu3FevFFI9FnM388x4pypYLXuwA/1WHC4/oPR7uX9a/BUyyP5wXENulOCEXUxc
HmFnTFsd3oSXIDUTF9+Ofipq0wKKb1iTk2Ot0P9fzYhxyGBT7MXFIgv/PcIsJ7iE
iC/yTQ5Lzp3DXF7SahG6Rcjj/KbauVC0B/vW9YYa+NAlNV0cP2NSJpzmRGl0G90a
LAj0m2jmktq4XqSvvupuLYi6kBRgwR6kCKJSdXEsXGQmouxlpN3SO5znWjd8e8cm
vIrjJwxyLsdvhv8prRo+L+xE+Su//7YryGX17NnVMhkNoRSJNFTk5Ej9Or+jd6ya
YgvBwvirNYHKqIsS3ysDhE/QrCf3PsEAVeNo9dk6U1PtxDfHraC7RGCnI/6zmxcA
K1mz1RUL3k20JlLJPWazqaEkk8dITT2ynCVAAEMqOj99RIkdDrRUMRyw7/MxQ2Au
1hfjkjLgoErYNAe77BCNRfU5DPOwPV0OrIgJO2wSKRo+lzYfE0YabS5JWfUAEsia
NqL046ru9P6j9BFkPuzquVf+5pXnTKWnTVaZD1FZ9ZbH1m/39MfVO+dNgbsI2L6a
LcjuogZ7pr101Jl69fuAripayaE6v1nf2vzaIVCOeb/+G6yWUWU38rRkjSYufiEh
d/nUBWT9GCMwEqe+zI1JQlzDUrl24OL77u1IG3msqBSwqLWNOs3XqS8OPCnI4G6i
lK99My2eqMgjtnk4mTqYX6RFjuZWoK1m9wPG/O6QvizUzCEhL5N6PZIgusmV24RP
4OynYqYgdp/ADzqSJD7CDgDoPUV7jnpFuDPWLodauv+z+JnG8Eml45oLvEVz6Zyf
HtSV+/95vr2vH0sQ8PLgaWStHp3Hg6gFmI03dQd4RrTKtKnf9nJjtpR4iejBCQ8s
lmQrs056FuDu2eHTs20wWbOUtJ43YFgyOm5idVG9e8IGQm1R3NS7aBWOzj2J8tt/
rC/l/FBg09ZdI71O/oPRW/j+1dIytZM8pyo8AardEoelysm59/O2uLPy1Rw9mOGo
+u7RMct8szaqVPesqVFG3CFArI/KgrAj8wzI4DC3hbfWIMviJ4ONnJBngfjqmmmg
wflEaLzUEs1tMkcF89RaOyWQFqXLqUBHQFag6QdsXIG7PNlKQnKZPhSHn+a6qS9K
FxGHCthi8LaxGomyufGbEKZ/B0f7UdbfAY/dUGZj0GG/fHcSip0+wLv1HK7wDV5d
UgQtHLCS+g2kn6AoHg15MnVtnbrjiiQfmVEH9bz4HHsTjX7YcdbpXCgWUdBsgEqX
vDSFFpKZc9IDuakYLBjOmsykPPKCMCf6+v70PO2UDShZHyov/BxslB9i3M9khV1j
v+RZmQrbRcsaf3tuK53gX+Njwq+g5J+XzN2cIkuy6ENNvKvRyVyoUdj+Max1oo/C
OQ80dcdPOqmQ5Um7qv/2Q8CgxEc3xr4+HscA/uH/FI2xbHdVZHU1Hu6nrO9+RmfK
8Km/rZQ/mZmvMb136Awjxpd1KU9Vr5BodGGsW9D4uMs7HFCd4GHUs7gtefH0iVDw
DXmDDSrPdi4ouIqXyV5Fh4Z1YZGp0lW7Lu5iRGGltRJET9nMOjymujnHvWKRI5ZU
3NEdc4eOe99wmuST5kfa4R1zcPfzButIMXqHP7cSgFGpyijwrk1yHPaDZiejSQXW
BOTioKzgrgx2fI7nuuvPFSbMFpjcRss4ZoFt2J+hcitEx7AK8PowM/4NLy/pUH0v
0yURKOpd5aaJ4CQZGzqx1hGjp+tspdQts9DVsHkN8QFkHzrFm0PQ3sXyE+UiG/Zu
HsFPQc8ioapTvRkeHHeBo9jnfkcHSfViRWv4ymzm0oG05DPQ1n5hNuLpI9XTTPXR
fgZA+HohmaZW2LBlrhdn5jHEJCJ6rpZ6cIDX6lbFHbG5NnPFQTqVe+9zr0c0cuxK
7jJzFVIJdobd7BIlkodyMPxoHixkQINI8tx59+Pl8AHluDfhBFNrJEIRD1R0rDHg
D5XPZ2v7gL6d6P0W3A0L7sx2G6HWBaKfBFpvCS7z2G3pfoFydBl4M7DSUXExOm7A
YX7ZEe+dGQm5tke5TIjvVN5x3i3pgevGHOzrX6OwtoevLtGFisGLvIMPl+7ZBeT3
LvCRsrP1jaTl3RAMf8FlhQR+nTkvEdpBlA5agUF5GbVrpAx7FneDP7akbj1cnSc9
n1IM5BM7064JeCG+sYHEKFK2IKZu6YBkMJH1669mCIT3jUd1zIifSglYAn/72iJV
EYgqZJ1zFA1uJ0Gwegh6mH/ABtj4/G5qs7Z6rKuAkxQdGmQkVMifpngnv3lEc3h5
jsd+0mwSTn3dkeL5MgfJLzbMfu1pc5a5r2FgDuZb+beT6ci3bC3PWFh+GkQxQOd1
2ZQQnEsNwXBr/eXodpgVSk0Ffhv3BeqGBnIOdtrKtkuUIc/hZJjaHFiayvS3alUP
V/I57GbGZen1/AAfTR+jOXXMYa5pehmbGJxsRqC/TEVBzTqHaoJqcjTyE8VVQtBp
79lMCrI1Jfz5TNqjG4K6qhI8U2nGBCJpHirJy9f8eeQWKNtIpm7Hdmy9Y6IrJa13
fG8TNORgzli/oZGup67fEQ8TZcs9LnMK9TxVm0OlGxxYncEybxW/zi56mchmqix4
53LMFyqvqUbOUkjfu635eaS6hfBaG9Y3fZYWWGmfQ6Ng8+vgKh+ka+knoSvc+UbX
eZxtHFW77jTp+DfIboIUk7d6CY8Hv+QX1iBPi+t3/Q8r+5W5Dwp7vYSJYYcIJP9T
8lylY4+7B3P81PoZaLpHGCSEOaGe7RP0izt6JuT0uR2RZ17KlaO8dSkw7WcnkRGs
K4CUdfAJfGevkHNMgr1ewr03MFcUdO3M1a17y27rwD/VPSRMb8F7WK6ofPP3jHwQ
Gt98cjZZL5vXozSHVwyIuU2TchAfVMG3Jo1o5tH0q7aZS9agZ1gFUVy2l1/YoWN8
vKJCzO3Z72pmij3DW/QPgSCJnihe5+9ptzkOJ86p43wSUi0QbziDWrWPfwWd6/V1
Iph4+khd5SwX4XUUDFMm8EA7bvpTIbHthjotMxnn8sJ262Q4yuQ7EnTxN+w6xcQZ
Sd/EUD/xuF6/XNRJvu8dqIYmwH3moN5s1W1ydRAuK2dBuvnHuEgKpo6nJiUnjJyh
LA3E4C5rqSykF8F+3VMAGnILP5Garx3zopw3ek61WZr+cDtCdr3Eyj0UnNfy1dJ/
LljPJNpVL1JOb9Xv9AKUx3B+X1EB42b/KnExgSNhbST88zMvy3pPzgJX+XMLDHRQ
gP0Ky8b9NfGwGqYqYlS6ufdFi5ytBmp1IzdsPP2qNKPYuh+gfIMZtdec6NwMNSga
Apur4ZrvyTu2YdZfIMOKcP2gGN0wBvj6PuccSyu+I4dY3D1yJ6Jj3Ta4VoKRz8s5
uMvf3k1HQrbRpRU9DjMyPbVL30fMt+w5yeJLoq9vV6HgQaZUEqVh6bVz/cWghS1Q
vYN1SW3IBJ6BKH+ZrWLm5lVI9qt32mw8/wBbHQ1e0dbs12WYo1NGxoE+h6uBT3Vs
pahjJw4lYSvCMjDOQIqs40Ajmy2qDepNLHHHwPPMDg4ZTztjLZH9+/2Jk+Ex8lQW
mq/EFqLm4JMd9Wt1C/6ZxIHIWBoOs29Kl1iChH8n8lpVp/c7TTiQLgeB74YKPsyX
tqh8akyzNtyZdpUgTpZBX66r1gSmzD4erzQA6IhoBvqGRWGQMWo5CAiwj+EKdQ0c
hqgco1wJM6yEvmt6dJ9OBYeW8PE4uHOlaS0t6zTrt+Ovr3aXa48xq6CodEmOp+rK
2aGDSEjUBVzDR09Zs+WWlMYpSxF7eTG7FWdM30OaPORuakhov9FYOJYi07JvcLVD
gwGqSH3vPwPIm/f3vr0EuHz4PCKqxAngXuyWSQPH4RB/x8D5zu+u9Jpt1evv+KfE
V+QA4gE4YJP8u4DRBLS94ygtnMVdPYtlw3BoObKwXsA/b3mXmUb2vfh+XH7JRDL4
sbrkRBuZQeyWNN5VALJlf/1h7+xIAP350kyKLPo4P6tA9hx30WRbi7lkyIAcMBmn
GZjLObZJ5Xwsra2ts4Ga7MkA2PezilN3e1TeHbcBCxgamUbWYB4p+xHA1Z+7hQwN
4xW3p1eJ8SVw5UXdnt7yYDd1pccGjqENtAOD24Bbo8iss8jBjzCvtxCbYRE7E5SD
kQbi9Vcj/ISGAVwbImhskcIC8vkgKHurCm5qcAGiX5dT9HJgVAUpnVaJb1t4WMpR
UalIBpVj8CmzJ2cojWO1TJqkBaSnoP3sUN+si0YGV27ep9Hh/AJxMbyzmvEAcNm4
Oj7RK9yRdhsGjMH+L07jdltQBHPMCWkuqhM5zCYEa0VWI9ukWm5aXuL/dGmPpZ4v
wTgBn7fAGcUyPyQHzJtjGEsZDfnSqHB2sPj5KpNQ+1vF9rUOyK5Hkii4zpN+Y1+M
t9hZzs3vluXIfy8PXsji5Sop7Pk1Snpc98GjZWA/+FkYEHp4EST8BF4e5oioA81V
9azsWP3HYjflP4RCxRrYTMMakZhNPyXSx3VlnrRkEx1k5tZWjHyhP5moha4vz+CI
CEM5NPo5Bzk/tLpZ+U4fOYirypAHu02Kq0JyGWRZDbDJW/UJ3hLhxKH94FpwmURz
ZfpQ1bBDRR7vFV80zJnzX9YtsgkT15oZqZXAVpUNUpRjrdzPjc2kI2/mSzCMwEP2
ghqodKcXXf2tD23A9m5jo5Wpg6bExvXY2N92CUYbV4WDuynD220VqVA10ddXyRHU
MuMZ/qTgrFsbzLuHTGWSmgFUHbOlbYzkj1zpb6qnhkObWgdGIGY4eAvpiZcWGsvf
xqA0k+WNIL3L/NRIbg3IrTxbacfEx25flYPCOkoY9R9G9UPLnPmdeSNpl4+1Yop9
UvNRycQCNRnWUgiw1JPw3hKu+DA09JhiarXF+pO2BKa6MABlGISnnK4r/Evccand
DLzmmDc60kK5CbX+y0cGBYvloSsIkL/vDAr4mhwb3kFUiQF9LHwv1ou0sS2ruvEG
tkixCJthGpom4tXzwOhWjXLK8TfsQ06x+Yv33plg8rd2Ao+aKQ6vP+pj9b6lZ2mp
ixHoxo682gsKx7+7MG42OAYdY2EvRuAMBV/3FZ7aWHnBLwxkIWz89gsd0ZgdEatQ
aPQuuTjnRKkFd62482K9Pk/Bdxsfl/HzWdin+op31mvuS5fTYnv0IJTMiMEP0zNg
4c0PmZTKwW2CiW+mcXg2XhqlKaCVlQn29wbd0o7NAbCjyjuPi2xhjujNN7YkBMLf
D3j4kPJ//4hq6ycmL3TbXosxr0h1K34QZ4Ujpx1QkVcz/IXcDe2edgumBypIZ/IU
cyyh8qhoD2Wlb1uSs91srjAXyyOly0tDsvjy7prPTY5L49JG96rD0bV+ET9i4cw3
d/chZPs4fzT49BqJomnqv8cLCjKyUGFxB+63b0nbQtwbyrkY/jjuVg21a8f8HhCr
qBUwPKhEWPCDq2XDfR9eLQGX7mEtQBTkyRPQ7Pm/eUBBi+0D9fXkAskVWxrzLrAk
cE7bDC1ZWFGNjOA8EX7s5U4RHXg6nLLCwTLXX8XuLc/vpH5u176DG0VwLzjRiHeB
KE6I6ZJReX+6l0owiLrkb/IBu8F/t/GOaD6/nMmIuuc=
`protect END_PROTECTED
