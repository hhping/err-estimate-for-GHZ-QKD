`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1R6ym53vgerowOgSZi3nsJfgb8AuZN5FS6ODKNa1nHZJeXjcub05UzaWRvw5hSP
m7X6H87WpJNqtPRY6PeI5Q67Mqb9MAuZ3LMHD03T64rPxhhWXjN/mu3a4z1IS69m
kMEmNiJxWCxDIVL4xyPrFfw6p2eY02w9vFTOrk8FvcMmYlhl+QW2FaAb4ukkWHwD
HIP/bSAbhJJ/pbWzE8K1CKig2eZkqsdOaHsoocd5orMVf+rQGTc6mfGknfGpJR2M
Oo3s42bQ2d7xL9wyasMXlelInOFrrPEkbQsXacYS24aYyUchp/aygJ1PhEz5Obwo
rfxj8DtUbRKyiC7MuSWaX1nyBFz5cSAPi4MUp2SGU7GR3QbV21N1WhBD1yProUOp
x1Z0WimUxXS27TKdUgcmjVspp3ey2JSygBWvSuYwXNdLbGfVupK/Z13osPoWslPi
fsSbJS9GoMUzTTA3GItYAFDKTulnzyEU+4mhql/LUoWWeXwORnWYTSy0VPYCEzCy
zL5d6IG3jaKZnKG4jvu7u/uqbtSJ17r8xVCbvI9KLv8gr+S9P6HDmD6IuIkVvDMU
f0SE4tCMGLOaUOrECsF+367tJGkHFdx2juy+i8naZRWttgRB9n84u7b4IgnFGxbx
`protect END_PROTECTED
