`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ph0rhHxG7UMnUoCf/XSt3Tzyvdla4NiWRTOCTF9yR0GcVZb6+ureUETYgMOhlXd0
4d9rg/MQqzKgqHKp3J/dAUeU5mBPUwesvjlY9tUpGRiYb4mMyu3nTNdP7p6Gdvjb
bOt7QGBNpwB9jJEMRcviTHhF5T6fEC0rOtHNOjVQxo1Hxk32DZ+8WVwFwWHDvmKA
B4kMAk7UEtFMoK3uOHrB6ePjpX08xAdTDcPCqCQ5jIEzQANpB8vU3O3fJqzorjYf
RZJER6jwtyw9LJNAGPfsC+z2tqbInqyJxKqhRL9w873o1zGF8yuQOQGbD/PErxYu
XuhkhEBR0Y8Kgxy+IpADyrobhm1Xv+9X+6QlGfkm9X4Ewg5hvp1at2TecnCtnA3/
4HweRD4EpLd7j/wzOrl6bNJvr6xidQiCZbmLymYhG10rnFuxr8wPTDs+YkM8LZ9O
ltg8Ea0rASGoOjzWZcI+m0cghSHYeDMLSc+n12UbZDx43yjMHy4PFjEMuEzQvsPE
iBdHMyAZXoQGAu8po9VzxZXA75Bzf2t4Y4CQAU/QzU007UkdMDQ19qiDbQ+nnojd
zEPRrmrcF1XovxEGGIRwToZTTYdknBr7U6aahH7UGydXEZUqgNckqymJacjjHRyi
G2BGep6VTQaG6JpxY2yzPQx2tEvLR7ruHHD8ghkwU6lFmEQBKAHcjQkonptRFNlQ
pjNNan7u2C9+s3fQdTbzlpBkAJ94QZUPIlWbuoGQ8T+XeuIuZoH7H9GQBrk2B9P+
TjhdIiMCDSVPYPTldykVpZk+i1Pv9ws5R4LpsoHP7TJDiMLozA8iDm8H+J29CpNd
`protect END_PROTECTED
