`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FPBTebk7Ldj3ZpbSBkyp1M3gE5xg9FHOEgn+fj8L+jnEliTBB7X7kuDeDVlk88O
EqpsrIsybv/qwsluHDfMcotjyikaN+3XM0ekOPrwZ40uuu52JTyYCQdECxlrconw
7Jtwu/uBfYwxOOBUtEz1ZNbz36+uBBD146TfhQvEKnixpnAtuOobgKfRkObhDHO4
ZXJnyGtAt8i58Lxb6a+1VKB08VF2x4IwSyPlNVkt68LLxESq//k9+1xo8o7B1C0i
2fVuxhoPffaK2ppVIy7CLKCrg+m7irBiLJ9yXVOzbSftMMf1XzsZYXqoBFVGoDZN
gu1J+Wn761kjczrKup1yFsaHP7vc3ZYjseZU1Ae1UjbKNHntileMpDcaTCt0ZiLf
ZyvNh9fMlSAsHB6nWh4vfHC8imF1GpKMlqr0/iupmZZvOWxCBheOpalY1irPPAui
4aUf6VZv8n//IqLX+FlCOPjOLfWih504NOALL5wDIE+7HcE3DOfIAJisRFnbY2LA
ZAVif4kW7QoMYQxplg/JcScSSWFFtrpDQWKHYLebrGm7P39e9xKgU2WMl0Yws624
A9yHNZirYFzIswXOGIP4VbB1NSa1fJVkn3bDL7+kJvZTJotjxyH0tvifVSh4os/W
AsMt88y6UkMOPOqo8edrPjy/arFhEA2E2JWvwpFow1Zdxc145Ep+3/BAyesSKvfN
uoXv7NZK5l0hIWfiIdcApHC8bc4by29rVLKnmrXfJpG7ZWqAMOQpy9jjRpuyIEjI
`protect END_PROTECTED
