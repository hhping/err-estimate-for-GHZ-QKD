`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8tdBvPdS7rA8KspizACuuR1wnJLzAPPCLZsaznvI5/GHe2ItCvGePhhBIlf+3FfO
38A7PFV6hiTKoAjI0ApWORklK9MFX2kk0wR5Dfepk9WXdKGA33sd8gAuQ3T4lLTC
0J4MQbkui6slDeiJkjcLYtxxGeHcXdHBZRrg94HrYvegW5nv+OKkOnN9cbQFM84c
MguAJxprlT1z6DqQaMeFQ8AMmwPvITPbVySG01ZsqUSV5dyQUzcDwsqoyZuQcIR+
ayCf1yeBaSm4fKEYC2Ldn9iuBJXvAVV195uUphflqBFnZBDRsyUzt4aIX70NXtag
/JzR8A+dA4TNdK3y+ngJB0MrzCpfpJ7g5CVSpx+4PGRA4q+Mkj6ZULWy/x/BQPJy
DLGjYTC6Pf54d2ez3QJpwvwzflsMNx8Cu8fT5DiXH1JebIG47UawzfOJ+Tt19sSy
nF6RQxBuGxRu01qiKXrr3egXdVShdNbPabXwAEoPCR+haZii9Hk6Db+WLb46mb7Z
nO2wNGV3V5sOycizGCaI/KqIYvJrlj0IOVzPgG23edHbE2anqolDaIU0eIIlq2hB
sAbXeiISmK6dQjzzjbRfTujpGMLXWrNsk+uGg+BRrwctwoBa57yjA+ap19tLuWVe
2xfudghWvoG+1+t69S9IT7q7iIc29ZVsDJ/WEAFv2QlU7gmBVbZOLyDRgBQyTLeR
paw2OoEhHS1Vqd+h1L+euMXe6pMu45Y71BlCZoMH5PZjj9Snm7OiIXdXaK49MB0L
lIOaAx0LoCPJKUdGLQuMOZi8Dlb00d+nP8aJcTd3o8l9P07Rx/jQRIt8YclPxAeA
hXRZF+ZLxM6iOHIFEzlpG6+7RUJCDLhV1ucL+WUBi06qHmkplkQ5+6oYHpyaLtgn
UOQchvCRrtYsYSOvgnb9v7GkoO7hJ6Ozyo9dHJF8hQ4czDDsJDAJoUzcCo9euxYK
fUQVKbzLaItZ5RxSEekR1tS0MhUmjfLZihBXETxHGmh7eL3e116/VC2ov6QZD9Oc
p/ueHGqw0JRVUQu6NeuxidW6CYq/371YB8uOYH90hnHFdF8aSbd3INxJUInqE8il
dOqJ2ZIaEZ9fokm4MViWAoROyu2xPLgg3lT0Kl9W6KjL9RqphaSgg0DxH2Iv2cZ+
vTk3CWytFrOSBajMjqgqI/6K/9/EwR8jao+uZY84eLZZ5RdGzd+tqBRJDm2y8k+k
98J+fMcy1qljXUxTYTtUlYGZd07NzgxhHMk8eHxXnHzxja9t3oCI1m4lYwn2Y3k+
ynX63/Y1izR/ra2VOPbiIhv4htqLMj8VpaumWg48oKlcgDMICF3YHYaatsgdqM4t
`protect END_PROTECTED
