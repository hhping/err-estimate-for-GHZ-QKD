`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBs/fK0v8w+a3nFi/1esw6rHBzLn+Hfa9VBgjMsxQklyP06qYO7xxzce1DCuHhNI
LklhnbS0pBFlAFiF4C66g7oJO79RJmkm9HVFsTGBIowHZXDpdhoS3uBa8l1/PNtE
lurGtNUWwGlk7FNOt0qJM6gMNOAVCm4fz/5dQ9EFDCvoWC2KvbXpQo+klI+94Iad
cytmGA7rgtcolVGE+wlIE/mEcXABRWPEb4xuGAQg5bLKHi5i3uT4tTjWAB44vd0H
CnVgFGKgAVQLYUJokml30h6JokX+LX8l2I27Eb3mZP5x+ddavYf5Knh3dxq4pgT5
0hcRJgKYbsY1SEcgfgf8+xWEpEcxW027J1wdv0ZH8gOgBLDMwcsTml5HfMYLVIcv
UHwYO+ReO8Tuw7f7vozePe2mzsDd7S0RM5FmRaJElATIzbfB9pU7gc3HG9wWuzMU
OjtUuRurtEQS8GfYMbi/VN+9W8ae08/tFm35haBkn7rXzWjYv7VAFJ1iS7s9gcW2
+L3tOEALrQGgN3kGbUjI2fbXQEXQ8KGrcP2s9MggEF/ua+c6eipE2IbY6KlHqO6w
LyqTqyhmHIUxVaOHvyvOr39ZL1WEtDQVW7xonDTwZwvPkdX0QvLWJlJpqbQzjsfW
5a4GOuiwOggse2Ouhw9ol72cs2xbCkOxfrR9e1brta2m07y4elhIrWKppFKA0c7Z
TlMXmAlhic/cpiBGilOzxvO2u3XCmE7Spku/uqixqbkVTQtTcHcwAwB4Mkcz9Q7V
MSXzd+QcDoxikMMEwPhS9Df/tZsbKL+DDExHT/NXgXp++GyPzM8AGDi6/glTWxM4
RDeG22Dm8OL+jz/m/xeXMnlc/19Fx1f1NpBGDqCR5XikRJPx12opea93C93CjSkB
rqovaFE5J+0g/eWfuEpfYfjkYetbpM4ylboojPsRjFHO/U22PKVqHFFjNURGo5Z+
6nTIkcRukZziBnnHqDbcB2Mr7PSqEZzsk9W3Gd1ZtliaPVHIjinjk7E9HuseIJCl
/gyvjdw+BdhGIdK/SFCSTt8wsVQMhM1rJKAVAWI/KE5pMC8Udg+gzhXLExK+Otqx
gb4GK8rQZgFFAG3YoJpeF2QePt53VAo8LazDPyMz9/9TIedAnbZGfhVbkRUrFqA9
M90tANgHIOO+s0ejo/RbFftWPgBdHzAUW7sApJSMpW6m+DV0+P3cfcN12D1Q/f00
sQ+udv6HxPsGKChd3BlFIn2r7n96xmPZQ8WviR/3AS+O66Te0gANf0w79KW4oK4r
6uTZFpXxYbEWQCL2v+8DM2krHSq+ZCN+yBtGmTBURocr4c4CjrtQpN4vhVPv3yiH
vwX7ibCgQOLEreQNFnBi0EGrW9GtecQczDMKtrbcGqlMkxKvV6LQibSoMVDh4vtL
HPnpU2DIRyVspRbuk1xqu/aBknYnOueE3YBsjcWrBaE=
`protect END_PROTECTED
