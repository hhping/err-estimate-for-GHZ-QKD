`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bU5l2cmPGlicWktepAWsYioidTVix9uEWAuR5D3sndGQBpjSBQrPTiQAL8WRMGAK
H1ZPSKlDUWXmswDSatAPIyUg92OgPKzUWi1yIf9Huog6SW3gBAyTYe6T+OhepeEz
0zQtSQqDi/tIOOubeFdxqqtBspQPja13OJw2SmFw0tgsEN2s/ziAMs9ycsNK76lg
V5u3cmH82bTf4BRXN04eu7eupKM21SFM7rXj50z4gr0zdytk0mHLqzDYlLpUi2SY
ZmVl/anASJ7y2KiY4WiJbQ3zZt0XFVk10ndY5shxh/nJscz3u3qk6Cg4M8a7ziYH
J/bnvUMP38ljwQSea0Z2mlVQwd4GQ07FxYlNWXxiDe35D8YOcNOMroKwVjzX6+bO
L3R36LwDZ/kcahuUWEFv1XPCHX5ww66ZcfZpS6WB8wsOmElH4pDA29+3OErIm1Ii
G5NlmVW2bZefBAYZI5+wSpE/SK2D3vbE9LB2Sj96PzcTn0f7xskxowF9dGg+wGNh
gn9yPli7L/qBp5GbhgifmIwKOrrZAp5YWrVESAMSnJbcQ4tHCUlmVLnAYPFA9p4t
llfnwnshMY4HUoQQeLo1vxt/wO4+MHklw1g7+yOuPPuirUeS4GBVhnrxLNfOMxb6
/PGE0bTNNoRgUsU6xld55KZ2EPG4iIE7mmVgPiQmP1wRWjFSJvvGRi05KoI2tO7F
ua98hjyED8Nx2kG+RVJzN2NRKSIIHYM/7MKtQvu+JPK/MSX/keUDsp/9xt/z6oXA
Ew9G0X9A5bkSDbgA/6MKdETh7FoGglWN0vhXZBEk75c7rGMYvT5AaVN5vSsSRtp6
TFTsJyT0TxW0oi5sPTGSiBWGhiC9Z4TiKnMhJmS1oQiXnDW4ilGtFFBJXh5a/68N
Xuh6C/xV7JvyLjXHp+OEjsYPEaQ0pTOKtSHCdSQFLRnbmJ0M47FIm6BCSFe6pVhi
CBHG7fKnYyG/4CNZZ9sTfxJiHreGdLw0YuddfdM+zgnS6h4YEKePvgcERMD8iiFu
qiQPK4a+JtUEIqcXSkaXWKpdYSRUAHxwDoY2XGdH6QNJA9PvBU4K+vAncWlNMzTr
rXCURJPyDJ5fE97oUKKGoyfJ3lrI83pUwd4Rz6uae8DQkW7l/hFbI0XmJqtl+hOA
E9esJ1yuwoXSDn+yQRiZ4Q4FqGtu9xfl12GSTG7e+AjEdtb7KzyCLSaL56oJwbBQ
Q/Jc+TFDrANQo2Is+JSqRbf1VtXWMJnFOhK5Rlzn3TYytdzP3uo3aymZgRySR0go
CKZdWpWcUo/Qlqy8bLZcZKhtzkTn5ZMsV93GwqheGoSk0Zgli7NF6kVFOc4spRS9
7FcIqt0i8HID/3OP2Py9O/uHQXU66n27EVnW9ZMpzfNZLTM+6uHPIcDjLBhCJ35E
3MgLs4dYP2U6IrgCIEIJKQ==
`protect END_PROTECTED
