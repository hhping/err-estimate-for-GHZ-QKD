`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmyicRY6bc/AmfG42b0/LtGc3cmi6PWvHSSOlskDTsgpcXFT456VthSM/qRc03Lu
dMfgXIjg3ADC666OARw30GygG/X5ESaUP/KHYMNMPh5A3GccHsJpUCzsI1wPbYGF
hl+Fyf+Tf4a5NEh9j6IgiVBCfENQ7cUkvlS7FkEq1GBwY0eRNacA4ds9GMY1URPx
Vpkt+zFCf8sWyd70DnXttAr9gkglWefETkXpcK+fiuKOJjRMSW094Q7oeeTnQYPi
i7A6QzAvmO+86L9sM0q91/LRsIAgeEBNvBHK7DW6xgZvYRAUrUohJnNpYga1yvtt
Bl/XVLpfk/NjYb+AawNh6ZaJqe7jtmFhLikzSZy9Qy15aF/ueu2JzgbOXo5axaPs
vP/AMJ8PEja5rGhhICeg02pwq7qipTPkbhRr2jkX5wURUW2QTgstOlnc/N+WMK3m
UvPVZWPQr0mlHzWhzOe8AanlZMoQUlQ7TyMYyjucTdzR8aemry8KROdh7vEo3hin
sW5ycWVhqShQe4wUN4jFu/KQsf9dBg58qC8Ompeuy3nuGjcztK7PNVCZtm5518K+
HgTqA+nrxLeTih2G2PIQmdhq/qhQa6Zeli1NzVyYvdmWMu29OPJXjXp6y4yGQPV9
0droYg9Eu/APliT4rReLuYkKwHVFjTjq4BSGDUqj5T17KknEQO4XWAuSlI3yG1OK
OXIzxuU9PSM+HQUFRxWMo3DYU/HFY0BrWnZ6UjVfL2OJhWNsZk4UD/n59SSexwKL
uK1IuPIfsTGq/PLh1huNDCyrewMoB/714OrqvK+ofZsaGoLo09l4HexGr1PNnziz
b/4UhT6JUaFPn3S37tNqE+QaSJCdKe5zC59eBrIKqXBsJA/Gm4AMcIiLSA93GN6T
gvZr9we+LZX4U/JIGunvN33MFWhTunw5Ls4YNDXdai3ryqpJzcXTaosurdIb9pvE
HWTPjuwJJNbKTVC+247x8cC6GHCiIwokb4jgqn4HaKDoVDQWEzU1j36QzefzqImh
2T8G1EKezV3IZqR66omAs8htUnK88aJtd0wvWBp3xcnfvKv7iGQcl15PL5pkmtey
/7BtLXEDRQjSs/GC0Opl+EpRmc5S4CLHN7pgBCW+NNLvGEkGCySNc8BERbwvDvQS
E5U+IBkt+MZTQyW13Xq9ab6Mqt/3uBBs3/WLbaZd1rGnNX+nCCZL37HC1v2z4AO7
/s5zIFVhWOrO/tEifVAgf3N/Qg2wPNW/1gW2qlrEkNVLacm+ixuAAl64NhdYfGf4
Ze6YSnjmkpPmSJ8Yr1L8ZUFCcCMh6AplI6MHKvrCB1lKLikgsev10NHRxUgnNi+p
kUaqYXJvPo5Zx2ZfcWAMJPaaOyexLDc0v+++bjP8VUh4CTWKYrxF1K9dlcIxrzTb
Q8jUTKAXYx2ptBHVQgnA5FsrFtNegITt/40t9rVKSIdi6G0/TO9UH7r0nJUqkT+T
gvqD9035Dw5k85ejvmJlVEE1+/WiJj247kmPqNYUZzzFVGG03MMEXfQlSUK/SZRw
r8PAI6DOsyqUiw15sbBNfd5zERXdpyAf5H+vUhPdQ+W0EcqRNsG7uT5EMfNIF39Y
npslWd0WnFjw3RF66k/5ZdgLMQIlDkHO4cCNtSzEs+L3USInTYnVrhfy5yWxQcku
p82gmBKw8//ZOTM/PYsjAkWLBLM1wsQRUxwUMfOes+wWlT1mOWu/ChZcgfP1CFY4
V5K+Ku1ODN3iV54IhpKqbuPe7SBba2rMtRsZC312lfMXDL7/K6VCVaiQV0tUVUAA
vKZf96LcLhotDqOtt2OaQtDqhorvCT2xR8LZeP6/Boe2ugaAhzzMIZ2fJQmmZk3U
mg5qhRkqvd1zYO6/FPvZK2PjojTOn7BsDBJpQ3n5q3pTqPAUFrwqepPvizWs5i41
ofJ0Z01Pq948otOdTJKJ+rTooJpvwgJDBPCO+P2nuxq1McpRLO0f9MDtMUWaJmHO
QHIQVGQQlSUkcKeRcU70h/cPEQZpeNjtCEiUjJUEcEfYYH9tjKyiZw42Pu7tOzIW
/iG0YNrp6sy1XYDfgfutAu/zG0TiRXXnZkiJOt9tSrZw9mM2uZwga4B1Njq2FpPt
nPUo9Dap5ztyVJcpkxU+GZZ9A/0+STL0ZzQCSlJEG7PZN1WsDbBCYmdC30V1V1n3
DMjN1myg9PJkdTJprRmISj4A/AXubz8thk65/iUbhOM8Pslrow9ZQTpEfxXogKTS
3ch1xMvVRo6jcTXOS6TtIgXeOrfa35ZQTD7qm06lNU3XexJQjDgBzL3ou5wB1CQX
s5apQdkIOkBEs8FqX3vRRkfJScnclH/J0AjLBTcWBuZDTctNoex6MNLSK7w/XGfF
b7bGM2ovCl91NWTNEL9iiq7A9Hmhpu+vpQXLZZ/cifcaXHgIYpVK4r4Tn24jkCMe
4BwrFWAVnqITVnJhwTGPe5oWmaqOr08/YisAy4uWmVDXrUOnzcfnM03vZ5tM5Ktd
sg+BF1joVYvs4C09+psBXSkLOeF81/7ZvtD9O3POHhfCTfBprXnwfxf3LkCxZmlA
6XhMb5/oojhBPGcNSm++RGvqdIVQ9YZCE7AynC3Z2L9JOaRJIo6+2hqL7eatEuoL
0x1hTDtzmhJcRt35n4x6ELxRNul5NpglwLPq0vZTLTefuPYiYJ5jDDngWEbTKiCH
VVIQTtPcbfThSG4nDheqez9UgoaedLXbXsRzZt3R1AgwBghVI+yofmCNm9jD+zLS
uv4UNVv8K4u/LYvbKiefrb+i42jz1exfA2VmDcZKhIKIeJtwfJPw2DbeFDrLu82/
Qnw4nm+mlUvtUJq2eWD6bPVZGOTbbKxXgeByIMePM/M4Sy1I1uIfW93lDtHIT6Nx
Qo6Rf5++04IMUnS2jqG3/aSqCGiHgYSnngDf9loCRXx0W1wTl2kyg3//WE4TF+Dq
BTp6FdV2wpjMVqhmiXT3nqyPdVcJ1FADcl9Dy6QeR7XdbKfjTy8OXZ+8bRpkq6sw
R+cmSByUcLr8o6OHmBhQPZMUCBkEqnv/E40dWuMHLWwyh6/GNRA+DJl3VvIy9aXR
zOPedr1KDiS3BKFqyUs1gwGSPsPt4WmAlkd1uLcaVSRmwCzHV1J9KgfuGx7p3qb/
7gz/Vm4UN1Aga35+LYCKnoHK1XY7mv3iDpDCrBjTsS4=
`protect END_PROTECTED
