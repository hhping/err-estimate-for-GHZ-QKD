`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n89nm0e2X5S1vP1orCbC4CZ6objPO/LGfM79hFXHbJyGvsUCTYTxa4l/sLi2tufh
5qMP3DhBLF5LTnZUXWaceFQ82kQq5WheT2Q/JCT+hK7xo2TwOzWePzofiUCfcKHl
3JT/M3daPx68ZWLojB0E6O/u4+kfWsKIb7U4w/s04R/SxntLwkhxDreOIL45NBSv
zXQ9GhgHJVI4F80fdTQJ1op2uU6Cb4txF2pSmZRyYAvqJ3aQn3UOtAIwxt4r0gQF
V2ctzpDcknFy4MYstnSrDYur6ByjzES8u26rjoZPQEOs4gtH+rKS0PjoI/1P6zo6
opLJa9H9ghdjv9RWbOUEPeBPCMCwk286J3cMsdt4FpOfb38nPNduiUdZrYwu0eAp
nidpqFfkTs5fm1RsJKQzVBUGLsgJSv4nNfElW2eYSJPKmmcoywzjzfiS3YXqAhyU
eTyoJ8HV5JSLMV+1jMZWhb9p3KvvidXcRqPCEgl7xMSlGjYRoAHDEWONODXgWaol
8N3napvmkG2h3S2983oV1J7gznZQpX2jkAxi45Pz0zCFzBhohQ46fuKSogxrl1oM
TFfwEKkBsBbSc5jq/Ov/1ihW6bGzP7ABk6Ai9k8Cjpi+V+FLJT4UR8g/cb4zskmA
5buEo5XKfyhhnFkqU29j/A==
`protect END_PROTECTED
