`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ESlQfHBnUXrUd9JqxKJFh2lDOSteRLyMMEV4ohPGGqZboEJv8p8pyIHrw0VarDVf
U7X5I3NzX0ACIljinr+ipsRfF1HEi/AboAYAosQULOHvIT39hob0MwmHx+y/c7zv
QiiAvApFckzcaUokaJetMJ0y/K+vmvc/dRmykTJoHv3tWz15dlFcYFVQiAU9TPWa
wdWFeV6LFF30eushFSUz1ztYi5D8g8oAz/dO+cop5EAPFwaD0h+JYoUm3rrZd/lA
T+Up0/6qiYiMeV6LySTvUIYRvAbvveGQTtUtxqFvqUdSW467e0X2LTNiP3dTTliZ
+9PrOW69yc4ha608aVfm0SqlDtUmRKz5ZaH3AJJZ8HgpJA993jpdZp+OSCKCLyXJ
+GF8h8K/P3oGdnEklK2sXyIGYRtJSKHuF7+ByRGTst/D6QTrE/BDPx7Q/y3C/5hQ
tbMstrr/QG33ehJjY7I/92/KMfDheJYtio76TjlbyGFQVl6Wxi1AMk2xfQz2cDyj
9U/jaA3pJwwMrQgfwOjoCu9Ad11Ttm4/pS/c4H1JHGyli52LoAHfku0h7FgexM1z
su2m7GEtMV/q9E9FlO8t2kvCg4g8Tznyrs1ahK75evt4QzN+KmPZLK1yGhf0aoCF
HdG1iVE9pQVw/siKMUJuHwMkaUjKtmUwm+JqmW8CUyO7Qi31M69+nW6SWExm/tB2
heMmMqDyGrKJ4+jbNLLgEbDim40Fswwe+RJew2CU2l9Y/+Zh4GZuHyMbGDUibEPK
MD17TxvD1JD9BzNkyC++SIv9SskgIz1ubUSEzCRanec91b3xFZqtG5xKtkIp8fxY
E6dtQ8ggr1NiHpjJchviA/AFMqW4HHr2a9t9EETicwxeEEn9vpgrGHysmj2TPPND
A5OY2VCb+EGgIYZta1pOfTiID3fkVH5XRMbiwruqDuXKjd3mBsTR9S6IJTJsutaq
jwmrwgYVjWdO3RVM+4aM1iKGJLtL95dPtRQKP4CA7z1Zc429K+In1NwT7a3ALW7/
T3v9mr63q0ICJJVkeb8zvQ8As9liFc9NfsAlcGpvFBGHb7LvL7WHvyu9AinHmoZm
mDWG60MHPfDrl59dKgJSOgLKm1/8q4/WYJGx5UDnsowEQcuapBlonb+6/O6M+Vnz
2F4MaOK1PnjXB6L+AYQzkZhaKCn4W7+R0Qr0BCmJAwykKgt8yS9ZDBszRUK/HQcG
saW4NddWB7V1jNTUM93NLsntzYC41NZnJemo7TAEgKMYFilSsQZL8EvS/cCeAtjN
2OdtK0GGH8AIIR9esPzsMfAY5V0lVCeFlYL6Q372k3fevfKFOIZj/skrO4xwpE+2
a1pidw1lSZe17Mh4BB6BvIhua2sr53qK9dqsnEJM71YF/vDklIb9cnlKWLr+WPha
xDpSsQ/13kINQ2de1gYBjrLuXLnPsKg3pA1nKd19M0P+05p9BIz/lwN4gPpdHCDm
KlmNia0z4X0FNjIUYmoTvkc2v4b30CPGj6ijsa+OtAe/yO8F1slx2bnCIJuKgIrj
o7bvNN5M1msJZrpBvWSf7oTBTZu/N6dc1wOZ69Kzn2Q8rDErBwePvL+3rJ2AaZf6
uga+kRx+1gg39UMk4TjbUqHSdC8QXglhWAl5ZugYl/zEVwiTyIFXr8VIdItv8OpS
maCY2Y60fW7fXimEZlZH5VLAi8zdQZwY+HFK1AZYVCpy3JreCpQPVPmsMs4IJPv/
8S7v/0TWmOUMMNSRaoYOGbc9TDumtoX6GDWhZMg9bKMJtYIL9leTjebD1TPNAlFv
joMFu3/fJmocU9xZQJdFNVyuv+Ult/7nBCa0/ocvjFTiNLHydGhngh7TQtVztZFb
BjmPLQjbMGeSwaeVT3bwiq+ImmSxBlByWuPn7FAdi8T7WA+b+wvMlUtzNL6nM/nc
/bhfNInni//8XooQ8YrTOixjwi8EHCGQT+O3K+YalgbWwOLklxdBoieVdceIaXN6
x2Q+IPipJlINw6l9Y23PRb1eCGD/I2fzqkcvPbm1DQ++7OCPOB0nFyXIwEcAHVfR
rtRCVaNE5YhPGetu9hSLa6uxp2cQIk7lvi1Wpi/U79K5nbLC/o5QG7Cr/Y7LhjvL
W3feVickXpWXBb07Itsi2io895phxkWKRYwslwPa54fACdyR9YkJZhm4pUcYh3Yc
sBRiYf2RhpJtPmL5um3Cg/pRLPMkVh6hkFQSu4TsZMEg8esgjFuY6pEf/gjA4gfD
naynuykafvPIg9YTXPaAzvmboGk+H3yfQP1cH/M9/ot1Z5SVNFhXCl9617D4+RAf
6VaBQSBolF42sNIdfQ7LKdcRH30BhhLAhPYfHvZS71DBrfJ8C/EYA+02fceh0o/4
LqHyaK7Dv/OMDycoFtPwRiEpMEmnBlIecdDzS3C9ILuMceUgByMrqYHPAD0v41H8
PDpfHQ1hZQ+m0j7j2DO4nfhVyOpWYGbhteyueA8GbtHDF2MTSwilo1j0GuzqiieR
JlAD4S4z9E2o0JpgCpM779yhKP55fpQ1jaWsCWkfnXJKQvxHersr8f4eWeDF1WLZ
BOiI6y/Ge4e2I8OtLl9GKHi2fx2WNM14X7rD8D9Qllki3PKF7sHlgywSm+Q/Tn+s
iTTzstCNzZTU0TPC5CJ8EVxqevV5/48KL3LUwoZOLA0U7hJ9GuXhZoKCph1cKa8l
xRNFB/vr4IieMieY216zacePlNeJYQZZz0S1hs5TdgrHfbPJYO4slY02jnfAryLk
EwG4e8fBgBXpt58Oqkc0RhmMvaR2vTEQzMaV45oE2JKeZWpWjF2YBLKiSJUbm1e8
7qdsahCumV5Fii7kkJzc723JPOCGfmT01j7F0b0RbA8Ay5VjVO15S+ApmqAvuPps
Y5QucYzuiLSrJwF++kGfeRK4eqD0aqcZ0CbNY2Oa3rc7QEQSnXcCztRlylNF5zgx
UZ5CNonrlsK2KwitULqMEre2yQ5brlxqH5MbWb26y/rK9dq5/EZHEXda8kwAq/Sn
56LK95J/XKYKC29MXTjYz1qbZWHLgMRaDA2vTA/QLUjw8b0RK/+fq7CBciyTBD1Q
MQef4RsYKM1XI2jt9AbW9QgM8O/Mch3saR1GENcogrKyLYKQ9/IlLVQEC8muyaX3
L/Om9DzCwZEIWsSbNYNQFSQsSwoqVjM0Ho7q9TNZAT8Bv2gh/SYzpAfZJ7N9DA0o
VsdJ+1H2FAHc5Ron5t6jxjZnMf3h0hwQVikCYsuphzF35RRcskUJ+qV8up5efTkl
eEiLy6qt9NQiN64f2jEWBB6qi/Qjqio1YlZqrsUcChJ+9EuKSkPtzf2jnEvJJEN1
JN1BYPIPoUieF5BLt3ICoFnbvx+3G/Ju+QCJoRkxn+eniq1BGjOydemV85bnNmD3
AdsCrEpeMz4zGw1G6LW0cP2ya7CoIb/cEe52Pu84KfJ6JxRrF8tlS67OlynygAZi
Nh5htL/daU8ybIpi8U7wHh3zhMyESJwAlToKI+sPwxETENxCFwv1U8TpOY5JW+TN
0TWL9LwwoGAMIGCaOQDMQXUUoodtl3pxwC5q/rZhVP7X0+kEl5L50V19mnXBRRQ+
FVEMzyZkLhygs3urGpKFfZfxuyAxTPu7zZWi8wtkbDdd7pa2b0AvBG5gbtXYwW4H
8zqK/MmduLWMVVk6iq+e4NYVmVP7pAAspN8MoWUXmSno7eC/nItx7odIo0RicrEd
ABHxbePZL15wDcieQXTToigQdNcyR36ozOLuv1Pz/7xbH/Gwi/otgZIbJdM7y3E8
+wNyxO9FDmnn1Z173Z1hHWGrMGIGgIydFM3XIbVF9hWcgt6GOcFc0BA+LuIREftS
ntCok38/YR2riIc8rOyvyLg+PHENBeaxIxZtr2ifUwCit9DowIOMb5QtwvTuzNrN
cvhKxF3fY7qbO4xoFEUz8CmV/pxSVS9plKaGrTh/BSjZrd1vMtyNdukO4vr3OVx4
eITVUxVL2ER/Bvy+NoYG8xkManSPBUBqnqvKDugzY0tTIG3fShtaFxyCKOu5MF7R
U+gnrOz4wTCI0IfVOCWm1QKegQKhuRw2ANnv8gL4kPoZdfaPNF0uQdUrW63uAx96
jMdAhuvXW+nVBlVfa0NIWuTp5l9T5xMUGZNrx8fA5xG1418a27iO9KNG7C/JPx9X
+Uzk93w9eA/Q+vJlhH+hm1TSOhJoZ9EJIIuQvNwzbatlGlkSg7v1Brmg5wuhTfSK
qLRbNuIX2NWLhmIBHzsgtSR85DpWzCfDg/0oDJzS0cU+5KihgmPWW2tPabjhINOA
g9ibF+JkusLtj60mQ94eaopkpW3yZUw2iFCxKOB+rqWR0Gsnk6Wxs7riPvhW8hrH
TP1dhJtO/ZCjZRQmA/L09daehQqVKTq/o5DnW57Mc8JjBtVXPSsKdTtPQGG7ZT4i
BoIB6pLQYnPvap8H9OsEj7PfF1uQ7tSQN9mUgQr+/wO4mF7BcY+1sPhvgKbNB5kc
aJm2viO8dC5Cq7j5Rt8MObuBV9w+ihBDovoUHeZQKwrghpbOxySjaPQy8MJ9nb6p
tCoSUXDAPN+lqXqkpSkgtsmulSwK0Xg1kqZDjkI0j3CvPtLPpqWP1o5pLQxaImcl
wFN3QTLPJFiihT2IcdI6UMHItw/ZVcJxeRuIhVQFzJ3V8xhY+vN3gs3iWfC3eG9x
yaCYKqCfUyPeNpIQDIM5r2/leDgWblxYHj6j1VRCjP68BBFCpdMAc5KwQO9yUoiq
42LAtstVkP7u5zRfEJBEznM1pfuL1hm13V6XTmonhLHysIiT1RyCVl2YFmBBFHDR
/LfidLSIdqtB+IObZjdukZnsWSlItIBcTDprRX+ZqSfS1DTRpwuJAT1TsyKXu9OA
8JgjIcihET4uMFj/SUt0JR8vPDMdULnQtJn8c6hRxIdy0JPc/wlMaiap86CSp+/V
uaidHXZ5h2SvnyhPWWji/QHTQapqD/JgWVIYKPu/fuOvDFYx8wiJuWcGOFTfHFsv
v2jqwzF+3W8kkfXmIlIT5DADDWLeaLU2Y0YO1Cw3NfCQQLI696YZvgZiPDYX5tT8
Jec0aohQ2NQOnLt3vz9fEg7P3n1HqfWx4vNToyVd16dWnsOk+CzfhFaKYbs89dGs
wv1szWK1qNjoqQA2wHpQBXaSpSxoAYRbMSyI7j2We2HfYXw9R5Se5DF/ERLDhWEf
bmMaV2sp26rAqcFzB1Ml2obb+n6p5lfz3zOe5s8DoL2rf0Fg6evR3sUKkCDi0Wcg
cIAatKO/pkTLE8+UgXqzH9wRNUQwK1LJzmam5L+wiSxhNURN3zqK4D0BTTmHLGPV
hHAQZRGSmMeD6CarzPXLGPh8QwYza0GjhSva41GthQjQOMUqPRAi3hJOZs/itB8W
SfimOrFePSF/hQZG3lSIyFn1Dub9f+/yv9O8Bq3CwzRLQrhgIpC2INbcQrJYr4rQ
DYvGwOALibxxMOQYLk/dR7kaDfbdZhCQrkF2CVLNItOgOm3VKfjT6UXGRTHNx3sE
QGg++7SMna9mfxyYmoUF/k675nbnu0UZaZpl35HWf3cw9eeO7ssDJdRJG3Ky7B9I
4tv/W8MkqyORFIW1gO7cgehNb62ml8M64ixMRxAUSHy/A58GPo5MzljwuPo7wLQI
jCtH3jS2cfgqlO/mEjH0YWsuZP3cvkZnQbvnxMeHNCzjgKWFr7wmujjoH+NEEBVA
8bk6LiWB+09uAOtfrHiIw+cqWEEAa8uyLxJusLQotZcm+LNszxhS87O04/jW5Nfq
vSAmA6g+xsJ80HN1ftl3BQ3YQX3LdcsmIs0E5T/TfmYcpV7OlYNUska8MmoP0jEl
X7JXTMekUqAagVIOYToE757ciPqihmp1XGJUfmkMhDXwB2Max/Te/D5ap3Fm0g5s
AwA8pCIbk+taH1hJRenNH8jKoRFBUTMjgVgV5A3QNuO+3kHrXYwDCmllvsGuU2A8
z49rVCx0sEIV+H3pxQqPJmU1KD/k1SStAdl+8O2zmcIaEtG68nEWcX8ETa+jIFIh
vZM/vIjR+bUCz2uNpnLluHPZfg8IbyGL1wm71lNYUegeeSMk1EjZw/8JfVAiw+p7
N4RFz6GTQoqCnHsI7KRKlxUn4P6eBXaKRB2xZ1mYOe0N7lfrGk3sGez9aJ31X4Zn
WMGvppkq32celp+m5mar4Khf4tQYfczoMm3joXHQf4yNOQ4515Pk544kjSoJsEsJ
V37jpV/1Eff/RNcR5H2/3pjwIzxwD9mTOzD4GN3x0dNZHW3Jk88Lcy4p1wgFZ6BS
XiXQvGGE5JdEkOcvlIimnh1blesagq5ZpASsYOhhJoMbaBGpaZFb8xOceJN+oQgr
bFM1WYRdaPuvhHqI9PHI86A8Q5c3ydBMEuXvycXfLl9wxr3PMvnRMpAW1PGdIer6
dQYuvqWwB9wozmmjYwn5Zl+fYzbbuUDNa9F/FibezxsJjUjswCzxf+tUdB/SfIu4
TTiwRlWbI7xsgq3EZi0JbkxyW5qI4keGW2B9ufOZQ18JBI4I8a7MuvIJlA3jkdjB
/rYOqVt0cFvhYel0ikTilPplhnMFMheFtlDCDu0mcJY62ueI7romrxVkslueoXbL
Uj+159oCFYsVwVQO1zn11VyigvOTnmtRqJGkEHjA3UpmNiZl/MmbmD0SiFLXZrwg
DSgw0nzKbJkWB6Lqsn0L99jRZ714LrRMYKTNWnKenK0ZYLEWUF1TzWynMD1lHc3O
fwXX2LRX30SLeanwuHxNpGvFI4JpRESKmeDnFVUq8CARUis+8vzJqzMRCE64mZnR
fJsFQhNeEgH6spWu4AC1TCrC0qtbTjnutnLoO6iyCwMJatsZYPlb1RzoMDM8/Bkw
83ePqiNYmGzmRHeWEdtDnoOb56TCKVWh4dORumQHYk2FqeMx6+mUj4MUZx7L9U6y
AElZLQLSMtcZZuhrUvrKU7aT3FdZAHVHRckp87hYOqdbiy7O1gBFgV9yWqOfTw1v
SCAlSUKXbwtMcJF4mx0j4c7ZTMRrTyqFQREjHjZ6LIpYZYCJG1VlPnnNI9Luvp2w
nGk7n3MrDIqJhzXnPAxAX81F+Q4I2cuLlFUKOdttbf6RfYMvy/9oSoJ8mfrH/Ypf
cRUFsNk6Jz6vcnv06eCmzmoS67T6kj5s0EFLETLicXolHBAYISamulIgydUk2Uj8
OEjg1viEDesspfclEVKa4/9MlHFGSDHN9Ju1yx3D9Pb0lhJkpN3s+Pxtu1qqdzT5
QkwNa5aqHMEJ/h7J1USnlCVGF5SnDhENvpXvztA+s3eSN9XcuElsnMKPKwtZ315k
0wdggcMJuGwyc76BJyUdFYssTXSnPXwRjPGzZbs7DNuX8Et2bU2/FTbH9mkWa2Xv
uyQeD8tH/nEQPoMHdQZXC4C+0p5Z0AURFTzMe7MCU/2azVGALOhuMX4PXmQB28xh
YT+5ulSv6gvrWA3GwH5P5Uopv+n/Yu+9yC0BiK4/PkOdXpWrk9Erk2BhpT4Al4Fm
RNux2cV8sM9YIyK9IrfufVyKVEEL4BvTxT2r4vpzTxhlYw0FHUJzySxgW0p5150Z
cO+hVgoaJOY8NcGEcJctHS4Tm96nHa7GNmjCZwPoJpgZb6eOWfutyshLLbwLldyi
SdpY1JrR0s8fS3teqqTCa3kQ8APFlEu/m+JshXX9+AG/vrO+Ndbo6BXxGCYMFuxF
fEDq9hIKclQRIc4LpLzSLbQovgefvb6B0TV7LyThSb4yZ8+DHvrEPXoVr9MCsu7D
C8ctxqPIRct/y88ZaX0X4AIkIyzRnmZPtWM/PvREB3Dhh9U3H3IMjsngAPdNR00w
chPzcB3oLqflw0KbE8rkAmozSa3msafRaAK0DEpwH1Cr3/9Y91wXhAbXzZhTbrwk
Cce6VCU2gr8vQvso7K7c70cNVXHvI4vPWxysP7HahohBlu9+wJDN+dt7P+zO26MZ
LvT1Oi9W1tuMS0EzXCQIC6/CJsZyFN/6yb6fnGcMy+6JV2IiMTSsT5M+prFzWvsR
U3vJ+RL1oig2KodxPb/ZxZYAIEiP17PGWbPRxNNHoMESRJ1iuoxVoQKj62F5P37P
DNra2hDqtH57+D6/LlXBwnF92W6GuiYGHBFc96CsiUqLcFJWiOmlfYBZYwo66ydi
DfhDZlpQx2sarPqqdwInEwJYsay+odY482h+aclIo1TCThjzoovn1Ub/nnCsPKfS
5dMz2UdmFlmOiKU7V3zkWNbXc+W8yTPMVfYN0Ui23PaDL5Rql+jF43IbrbanW2nL
dsTl5fcIchxhrnU7Txc7rXy5ys2oE/buGR3CcLqWNIspMGLOEEZ2OvfnLiJnFmTT
acmeRndnh4Sk0fkyx2AxlDJf44mtn+21dpggXp+SfRzjd/RJL2fDOHQAuxfwHCfM
H9B++y0/4Zx+x9tXgY2syJlSc2+M67I11vpLbUFaUQ4b/pJzGLSv2hIkVKDvQCNV
xaueXR8MhwAKKOFJtjhxfP06hBxKTL/YF6KkV2ZPbbmW7PVrVPOoCIeRPYDDPXB8
Zq3/tBHM+mVJJ7u0k9BwAOqIWOUQ7n8q6Ex0AwEuKnA3px9cNFg4az+kAlzm4B1T
wEOJU5XqK192CFNGy09a4Q9yoJkK4CpZFdZzElVtHhcAGBt24AYAedAeScU2YYBc
zEdNHRIMqhKMX043S/qXdU4in3SXr81WHgqZuE+PqQO3FK5wpOiuDNwrq3XUZvRh
9Vz6vWWN/8RUtPKopNgCdIYLNioWf2uBQkjO/COVn3SbrgZbBy2Vlnc/nWX9UR5U
QRfuDn2FJvPccfA6E7Bpoy7JWk9Uv5qU+vSrEoXYdN91nhlTrq3B3S/dne9lubUA
AdUxMzZJVfrqgX+dQbXxnntqBMjuUTe+xYUXhTjloDJ/LivgTuYYZkqqWWzSEobt
ybzcjcctk/cG3GGzLZJgFHfSuJI/4LRJlGhKOTyE483Ji2SLJR8v6KVRGUkR6DxY
ELFM85spNanSw2p+oYkj8mnBu3xV/dFpUdDNcfFdp07b4zBgHibPcdAP6KvSFS/S
zWMi84qdCQqhLmRygTyA9aMdyXt4uo61LMF3F8JynUsliWugsCI1z/PgolCar8R9
cfpZinG6EnJsmt2JVzuomhS05R8SYZIiACrabOXxEynuh8qo3QOcXMNtlMyid1Zu
HENLUW+ByWYgy2oMQbvaMWzKS6KLec5IvGgOlzlVvG5qrCXrXfFiDNBzPpVxjarn
NWu1cLBd3qZyxmS1iNiS1tohnLgEbdsMeSNp3p4lqxcqHXFi4HsSjxBBhi1NZl1H
`protect END_PROTECTED
