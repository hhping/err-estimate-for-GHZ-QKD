`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBVjnp6ZOVLAeuAYRwDyJ+rJhBONvR+fcWNtfKE6yQ+/JTAe4tvz8cDYLInTO6Ve
M8LBxqb5EowPpwfFpaV0BVU76tY749JkcMPNzhXfbikzww4LCU0RWKHcOFARgYQa
gtsnt4H/2a99B5ib5UedG80eaBxdqsIx0DoUqqh3UriImtsthUximzoVcb0OqBuJ
CDQbnTRQNTsJFCpaVucjDlomwd+eIHRmywYoH4UghIkJrGLWiOKMlYVloHRC0kpg
hoXvGnIWTHoosjQr7791oSshiyHPf+0tAKcht7/ePk6m0WeiGB/iuP4Yq1BQedec
578proXebLwKP+c0Xwv/0cPoGYolOuPsBYYtmkTyMc8s5cvV+0AKRT70O56oa6Gq
3bSNY2O9JFiqH8f2VExr2xuiOKoqCH8i1igVYMoiJaeDmrZGf8rfQbgHRXIxmXoN
L2b9BLj4ILQ1vrKWFqF001xvVoIG6b6qllfHF6DYDkYpUvTrlZcQAQ4y8jvfavDu
6YvrNj5Tdiriqnj2j4ilWyo+qEINoMrjKJh0T2hkjErmcu4HmtZK/a7LC+/2/zfq
`protect END_PROTECTED
