library verilog;
use verilog.vl_types.all;
entity twentynm_mac is
    generic(
        ax_width        : integer := 16;
        ay_scan_in_width: integer := 16;
        az_width        : integer := 1;
        bx_width        : integer := 16;
        by_width        : integer := 16;
        bz_width        : integer := 1;
        scan_out_width  : integer := 1;
        result_a_width  : integer := 33;
        result_b_width  : integer := 1;
        operation_mode  : string  := "m18x18_sumof2";
        mode_sub_location: integer := 0;
        operand_source_max: string  := "input";
        operand_source_may: string  := "input";
        operand_source_mbx: string  := "input";
        operand_source_mby: string  := "input";
        preadder_subtract_a: string  := "false";
        preadder_subtract_b: string  := "false";
        signed_max      : string  := "false";
        signed_may      : string  := "false";
        signed_mbx      : string  := "false";
        signed_mby      : string  := "false";
        ay_use_scan_in  : string  := "false";
        by_use_scan_in  : string  := "false";
        delay_scan_out_ay: string  := "false";
        delay_scan_out_by: string  := "false";
        use_chainadder  : string  := "false";
        enable_double_accum: string  := "false";
        load_const_value: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_0        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_1        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_2        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_3        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_4        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_5        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_6        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_a_7        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_0        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_1        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_2        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_3        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_4        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_5        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_6        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        coef_b_7        : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ax_clock        : string  := "none";
        ay_scan_in_clock: string  := "none";
        az_clock        : string  := "none";
        bx_clock        : string  := "none";
        by_clock        : string  := "none";
        bz_clock        : string  := "none";
        coef_sel_a_clock: string  := "none";
        coef_sel_b_clock: string  := "none";
        sub_clock       : string  := "none";
        sub_pipeline_clock: string  := "none";
        negate_clock    : string  := "none";
        negate_pipeline_clock: string  := "none";
        accumulate_clock: string  := "none";
        accum_pipeline_clock: string  := "none";
        load_const_clock: string  := "none";
        load_const_pipeline_clock: string  := "none";
        output_clock    : string  := "none";
        input_pipeline_clock: string  := "none";
        lpm_type        : string  := "twentynm_mac"
    );
    port(
        ax              : in     vl_logic_vector;
        ay              : in     vl_logic_vector;
        az              : in     vl_logic_vector;
        coefsela        : in     vl_logic_vector(2 downto 0);
        bx              : in     vl_logic_vector;
        by              : in     vl_logic_vector;
        bz              : in     vl_logic_vector;
        coefselb        : in     vl_logic_vector(2 downto 0);
        scanin          : in     vl_logic_vector;
        chainin         : in     vl_logic_vector(63 downto 0);
        loadconst       : in     vl_logic;
        accumulate      : in     vl_logic;
        negate          : in     vl_logic;
        sub             : in     vl_logic;
        clk             : in     vl_logic_vector(2 downto 0);
        ena             : in     vl_logic_vector(2 downto 0);
        aclr            : in     vl_logic_vector(1 downto 0);
        resulta         : out    vl_logic_vector;
        resultb         : out    vl_logic_vector;
        scanout         : out    vl_logic_vector;
        chainout        : out    vl_logic_vector(63 downto 0);
        dftout          : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ax_width : constant is 1;
    attribute mti_svvh_generic_type of ay_scan_in_width : constant is 1;
    attribute mti_svvh_generic_type of az_width : constant is 1;
    attribute mti_svvh_generic_type of bx_width : constant is 1;
    attribute mti_svvh_generic_type of by_width : constant is 1;
    attribute mti_svvh_generic_type of bz_width : constant is 1;
    attribute mti_svvh_generic_type of scan_out_width : constant is 1;
    attribute mti_svvh_generic_type of result_a_width : constant is 1;
    attribute mti_svvh_generic_type of result_b_width : constant is 1;
    attribute mti_svvh_generic_type of operation_mode : constant is 1;
    attribute mti_svvh_generic_type of mode_sub_location : constant is 1;
    attribute mti_svvh_generic_type of operand_source_max : constant is 1;
    attribute mti_svvh_generic_type of operand_source_may : constant is 1;
    attribute mti_svvh_generic_type of operand_source_mbx : constant is 1;
    attribute mti_svvh_generic_type of operand_source_mby : constant is 1;
    attribute mti_svvh_generic_type of preadder_subtract_a : constant is 1;
    attribute mti_svvh_generic_type of preadder_subtract_b : constant is 1;
    attribute mti_svvh_generic_type of signed_max : constant is 1;
    attribute mti_svvh_generic_type of signed_may : constant is 1;
    attribute mti_svvh_generic_type of signed_mbx : constant is 1;
    attribute mti_svvh_generic_type of signed_mby : constant is 1;
    attribute mti_svvh_generic_type of ay_use_scan_in : constant is 1;
    attribute mti_svvh_generic_type of by_use_scan_in : constant is 1;
    attribute mti_svvh_generic_type of delay_scan_out_ay : constant is 1;
    attribute mti_svvh_generic_type of delay_scan_out_by : constant is 1;
    attribute mti_svvh_generic_type of use_chainadder : constant is 1;
    attribute mti_svvh_generic_type of enable_double_accum : constant is 1;
    attribute mti_svvh_generic_type of load_const_value : constant is 2;
    attribute mti_svvh_generic_type of coef_a_0 : constant is 2;
    attribute mti_svvh_generic_type of coef_a_1 : constant is 2;
    attribute mti_svvh_generic_type of coef_a_2 : constant is 2;
    attribute mti_svvh_generic_type of coef_a_3 : constant is 2;
    attribute mti_svvh_generic_type of coef_a_4 : constant is 2;
    attribute mti_svvh_generic_type of coef_a_5 : constant is 2;
    attribute mti_svvh_generic_type of coef_a_6 : constant is 2;
    attribute mti_svvh_generic_type of coef_a_7 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_0 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_1 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_2 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_3 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_4 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_5 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_6 : constant is 2;
    attribute mti_svvh_generic_type of coef_b_7 : constant is 2;
    attribute mti_svvh_generic_type of ax_clock : constant is 1;
    attribute mti_svvh_generic_type of ay_scan_in_clock : constant is 1;
    attribute mti_svvh_generic_type of az_clock : constant is 1;
    attribute mti_svvh_generic_type of bx_clock : constant is 1;
    attribute mti_svvh_generic_type of by_clock : constant is 1;
    attribute mti_svvh_generic_type of bz_clock : constant is 1;
    attribute mti_svvh_generic_type of coef_sel_a_clock : constant is 1;
    attribute mti_svvh_generic_type of coef_sel_b_clock : constant is 1;
    attribute mti_svvh_generic_type of sub_clock : constant is 1;
    attribute mti_svvh_generic_type of sub_pipeline_clock : constant is 1;
    attribute mti_svvh_generic_type of negate_clock : constant is 1;
    attribute mti_svvh_generic_type of negate_pipeline_clock : constant is 1;
    attribute mti_svvh_generic_type of accumulate_clock : constant is 1;
    attribute mti_svvh_generic_type of accum_pipeline_clock : constant is 1;
    attribute mti_svvh_generic_type of load_const_clock : constant is 1;
    attribute mti_svvh_generic_type of load_const_pipeline_clock : constant is 1;
    attribute mti_svvh_generic_type of output_clock : constant is 1;
    attribute mti_svvh_generic_type of input_pipeline_clock : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
end twentynm_mac;
