`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHe5GeuNXolVZflp5vkHZJlC1g1QAE7Ry8SO0PVtbR0248lR4+aOnCLjiAX4AI/H
O7CuFwSeqXK9J1QVO8Wz3VhHnFMsUinF/Pbuprsk79vkSAhjbo4qsLa3LIrEPXh2
DMiKsKRNQlLJw/sTdxH+ljhRy187eWkvJIiNT73qtQQzcG0OEzvRc13tfoZF3xnZ
desDP9WTus6TPPLINKA19rH6N1X+HaGzaT2ykhwbtvVkjhS5/aI76iM9ZLbgZPOs
MTyxe94UPr84n34CUud3DSMNM4k9b6/TRyBxrle+iOWgEWNUue2cur6Ouek4xJhX
TgNUvbm51xjLfWADyW2e/CokLeBXT8DPIVbehwNLMkxpHKpOTqiA7q7XJaMIf6dl
KRA7B5ueDGNu9a7Xsitwk5A3OmTadNJtEtx8SDqxDR6NoNYEqv8TtKWSwb7As3hS
epbJON2chyZK63hTZQ8rU6FxqE28C0A3ccc28gzDmYsP4/2CiimHFCR56pUXftHe
O/WtJ7I0XxtSyLZxmPOCAbfMW2xu0LJ2KND5EUYw3wVwMv1/OJ68fd0BFklL9wfE
G7oDsozQICr6rLL0HVM4wil4eA+y2OzhdxZTllOux5ayiRF25vioYVD0RimtPOsK
Chb0eCf3ZQmoH6lAF+zhRD2TezTt85uhEaAvXfGNjlI8OpgXiz8N2bWZb0h9aFFX
8c7wDzseSzvSZk7YuvHtvjX+zjOeOQgOUzA2nMFDwuwSRsk8wKX3BKNzreRlsP1g
cN8zddCDnet06cK1hjvSlV63YRida/yQ8WgfZ5GVy3u9kmPkFkPPCDZRATx3Xt3R
`protect END_PROTECTED
