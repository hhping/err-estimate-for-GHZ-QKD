`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncbgcehoBZiQrVm7H9b2ADvEjxfJxJ1Lki69c3Kso+dPWTKtIayGAwIR/kyuKRso
2hPgGkBh5oX+/1IVjWfHB7i03YQA30W8Y1V37C/97eSRoXiv97rmLxPb9ZZY5FKx
v7Ra8cVerGxn5dCcJMeEcykktV7pQ3/eY8gwzJw4SjGojOwKfcXTj0chOD4jws0F
fSVcalfOv4hSWchCRXoHNwWLooOy7EQNrQAz/URbDNf4oRGXnj1yA0H3kq2eOeN5
3UeDbfFULn5rdVcJISryf9idR5MB8FI2/GaQG9CClXNfOi1gIllKE9V4qw0rw2TP
CsMaKR95fjGbtCzO/hJwPKvmixCDCiTbQomBThNYEBrhp+WJb08Qs3dxlqxd2ory
fUBqgUyWDjz8oIeDQfjWA0E7vWz+iRckAdUvAoKxWwpaAT2GPQ0Vug1LvmVarSMr
pNhkrLJDcDiGYPfwDer3ijxwe/kcmWtoEMTJNyiDmVy9EHhe0ldnDHDOomkBOLsA
1xLrJ5m3Zb/WhY3ticTrDX4rE627x7o8qurH4q1pgOYukYO8h27JlTCVYHLJYCP2
XEGq7HKzGppl201NCcWv97hn8KS+/NetcP/UuFNrEya6NDpbZwdULFFEZTpljVkZ
Q7rxMEWSzHc9/iDd9WoFlhvWFyJPgS79wUOjaKnkulShjuUgKSJN9xekpkt+vjkw
AR6NcaEfrfv41UX9fb8gUizSFggxHERt94f5lojYGHNse5B86qox9JGyJFlaNZ8u
6rUqSolZqdbJPwXmBbR6/JflTn5rOqG74vEDQznhKauwHTNXnkwuEuW3wlx+eMWz
uuuc8OBhMS2t7cp6j1cCX012p3xng//R4rga/aFGzGMQrRnoDI7KMGtkOZ9Jr7TN
0Bc1aKaZqw9jGEvmK5M+zFXIMTJFyUt+KeydeOHcQemfWy9FGFZChKvy+lC2oIkN
72AuEDF2Ee84iTkIfK2lHaEygkNvfGfjFZ2nJ5xv9AfmAkYsZP8DH6QybOH8kf+6
zx5yzgtzGLD8a2oNN5FFnJJn3hevRwBihB8ts58WaFRPwQbxNNWy6A9qoCH0/dRv
k6NyNX9uD/wfrX2M7vY84Q==
`protect END_PROTECTED
