`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIOL6M2gzlnU3YDExe4blz09Fm0I5GXRsGYStPZrjgvIzqQ6GJY4HHn6nnywQZQU
AOozY2KwQy9WdsNc0iq9+RaAbiuYMYmEENivQJ2/fqyOTy1LL9uY6wst0oUQIt78
qyVLuw0WRNSYoCiVYH1YcNSuP+VAs68CZ3FQK4jm1NzO5rqvpAqer+2dLL12O459
mxOkUcGuWUKgWltPOoBFw4Q4gwdtjp8drcBGpfeldZs3LKsg9R19ayFYZ/a9/0uI
JY8RU+S/VlXqvIHicpx/59h4v6o4pDwReLB41b70TPPXeNldKU5Zvhl6lGJ0Dttr
qNRMFHwvMJwAhd0OJOI6gqYFPnhCwzXhEwmBzBxHXbKXaOa/FZdUw5L+lNQ52Ih+
FKbMmlDGsJ9DogPTt2VfdH/lpCmU+itznMNioYvdEPV3m6UzJjtq/j0s98poXYmN
tJ7hmJDBbxZQUDnFKUXBoEgGwOlBTPPinw2RE6MwQX8+yCwcu1hhUGQbDuPIUOTC
vnmbT5hVmhF/Tz451cXgW60zgR9olap6awIJWXH9N32D6yfvxeHMXjmdQ76fKJh2
a2DsUkz/zRFiex2IAuV5HpYizllSJOWfbEhx1Sl+ukLabglrCzMeSl7UtpNnTBti
qN/ICm69trLklcW5JBdcRElr9SjYixKC/EABM9avPF/D6gQDUQqhbGG5LsHoGv3G
VFVTB7TT1J8Z8T3akVhwvRvRwkTrJcTMg2ouXBcSo40YVRt/14woEDYHTWVKJAtu
A1VncYcPmiDhzGBH11jWZNy9W5uBYkbzJAY/fnSQe/6q6pM9hnq36JR4AZSXAN+V
TgeuRwxZ5C8j+A6oQCNlciwOAdDFDDLpkTjRZLr0gtY19G8VOdrPZNv046INFXwl
93mpvuvkXDrYzkfRP3UhCn514XNQGxrmdd3HPtJbkeM+0TCE33jo9MZ00zX/thcp
unie4Ovx7RDXhFO1y3vfFE9oZnEkdMCzjxLBtI2S4nYzqWKUtMYfBGPnwZNTjpSY
++1xa7ABy9pRUBIucJ/gxHXiaRTPS5SXYxNrAl7vybSpSB1K8WeElqBtTiIrR3Q0
/rdNRLssWNsXW+xMFSb0rDUAtPgwD3FM+kWZJWy0owGzP1bvT4y7KUG8hgIRxiO7
`protect END_PROTECTED
