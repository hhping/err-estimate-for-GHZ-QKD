`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZYvaMXbCoz8V9PXWnKGcSqfwasD5LhzV5Vu8IY1OPBHy6YGwZKfszz9dMr4f5hfE
vNgf1v8TOKz4UG/x7QSetGpgq6xoU9JZ91TJIjXQaIDYWE+64ZkAoCoLlPfEsNjw
cVW36cptLHH3trNlYCjWEn9neLh5emKiORWY9wh20Maly83/cysCBdXbizkZja6z
P0QmV/An+86q3rsL46HyaJA4US7YHFRtUqnlPDlkBc12N+ak22TdhK23J2gsL69C
LBLSjeI94t8D1apC7yo6CO9ckIxbwT5vomNh4rm/6Ft3u8vB31wm+PGjqlh60Zkg
4hfIGGcchsiJP7hlFNcDPwJuHZ3GVEmFITnnb5P9QCw0RA0dNbgsmDJSkOQe9ER3
BORH14umcOf/7tGvpXumjGq2xQVtIOHxRP6cnK4qXX8FElIwnsVY5FKcvSVRmLXm
GbT491i1xrKlbIBozcucxkX14Nn59UaQLEGyAuuZLH/IbIlMuzyjkws5DngX2zdx
LLGC9grQRrr06duegT4cPbLj6JBELjghZhj1KSx+GcCTJKBFQPTpif9Uni0/4bNz
F9GumPMtnLGHvJwxpxorFfePOS/ozT+jnGWq3Y465J0DzjZMYephe8G7iav7u8PY
6q8eyTwoHoQU+og6wfKCz8fp1vu2oLE0zDas28rmnBMVr+OrJ9Bu0b6KIDSrWKJE
IN/RgNGCYww0TWOOvMGk9I2SnEXr6T7Oc31k0GLXJo7biKbriZFpQj34tIddh3XB
4Amb6Vf+0R8mLW+kTFc+xvjCF8zW/SyhRK3kgZfLadRLG3sD4cxBGQrFmTUGEpSQ
mX8/H2hkLzhVuHDDJlJaw+dxwLoqpfN2FZHlQxZox4rRM9Q7MhPmmP1+BawvohI/
e2ZAomBTkaUDz8+WSzehXjoEyhcTlwP/8yD2r/vu6TT4xnyKV+XpKZWs16TA/8xC
T2oBeUl3moDe1UBWWUmRFNP3uLxijHAzwDx7GP1WxyHYtQrCPIFaGnIalZOYU9uK
LdmjsGfnASz4NjxWK2CHY5yvLuVOTe0mhKjjjDMm5MzCDRzxt964ZrO0+9ChCStR
6139pmCVyv9FRDRtthnmP4mhidT0uGnHzEiIC+M/WAg/L6kzv5pbo01jAEng10pu
sK7BEuAQ7BLIuznUCoeAnIDPMaj2iGummvbdzNcoh7jpYV7vPVLf6AHqbIvnWj/U
uUxQYzBurdvdZiyhLnopbYRaxIWcgO4e9m3yBedN0JjSQ5bdRTxphiQaLIpBkhP/
rXEajM5hG8KnkNJLH2QkHUVo1k/HW9fqeIrLm1LJyzPshltr5Kk65x6dWfO28KEf
rF0f6Qt6s2HZHsE1Nyb9o+e09CQvfYzJydEcT8FzWdxNOXywmhWwEtOR8uO7Byvf
ova0v65DQ8L+HBDQNykbvbRuuzEBZ6mE9atvuG6GaJlcwRfNYdX5RGEnqzh5HsJx
7XDRsoomhax3JggLQZB8U1SRADvsXLyYk1eF4rCjmCHw5Gxa+eE29gbraeCggvZs
MqITP9yuW0K9R1KeJbzo6285dtnjMDuJplksS4LoZHdYWz0Gw6w8XtWGMijIptVn
nji7cpubO2dAQMtGdwgA1Wzyks0qI6wyNWyeP2DlnudAME9+RNu5LK6N/GdGJ9ii
+PXlYxg218XKHikN4t6qEI3Cw+g+gYFKDdJ09haUuPAq+qJvGpqcqJ8MO90rmgMH
ndDTB1jqMvrMuCstgFbKnFewKdUNJqmBIDnPxXgCYtQ=
`protect END_PROTECTED
