`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DBPiI5cy+l5jy7FxX2g0/9J01K7Mzevbfit9NSEJTFsewU8PqtOd7RxOJcbrxqNU
Mdyj6X9rgl9GU/8AjrXjTE9nD9KYVn9NVJmYwVb7AqrpBt1+WrBV4TQudhhvfgIh
dQIzHOAsViGdNCGmPiQqsVRTkTueFFBzg3jHVGCvUAu9G9IuBaAZOyA7o8L1qnC0
qXB9gBeRw1G6KJtaOvfU8erbyx23hjikUVkzJ4H1GBE1e7chEmzRPJSoRInPCSXg
ihSu14BZhpHrh5RXTHVmxJNZoqRot7no4Ul1cpzer1ytcBONV80DwBSoTKdo8VKV
m6OjTko8cJ3nlXPh2dG5QDqSc758o6SEF6F8v+gXflV4K5Z0fO0M2IrW8KzpCC1h
BfRGywi4SGGIncMpUmWKDP+TSN+e8vgI7Jlb8sO+IVkYs/Cpj4NtBtToZ/bEMjD7
P7Yg2Ef2Yyrc7e1htBAXTdsMebVpUBxoV3yfCoxySXxoMq9m5/qshQ3Ck8jurYIB
BxPZKxcbVVddLI8GyTUHywu+YwLdSHK30mCRs8G5ImQot5zppRaE/aDjFMw4pWPp
EcAy+dXuJArwy8VEEHgGFyN6ceSZwBMNyilraLZf0JEc+oBZWey1dcHbELUNXikm
iOYpOQgHDpEYoFcMSeVlg2MzevCgilmbwg9Nsu23BYxmm8wqvn4O0seOZQRbKQWN
Z/rtX36V1B0VQgmnWE1H/oyI6kZMXucHkr1W0LIhYhejUEYjuWbeWiilnnRch5dl
DpWhYru55636TuCqJNak+N7ieLGwFX0MKia5bZNMhCVn1TVOKMarWQ8Up9s3S041
`protect END_PROTECTED
