`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Btw6yCcsfDjPmNBDsevNciClUczsL2r/9IT5fKP/U3ulbAVb48WBKgjzmTEIofiT
qZ/Le1/bBMIX89WVke6C5bL59kAsQyq6/Qvq9j0EOC5slOS0O6aqUC8nMRGcpf12
ctIG24V0XBEDzfA9no0us/Eic0OY54PjQHK9vNtwpcT08CjcUxokT/oMVjXH4q1H
oWmNHrl856ZHw2M0C0D68iydj7a2BT22lIvLSRxJHO1UrkJ5GmhGWtVnd/+SsJi/
8/SdSA5Pnahd9hYKAG311ZJUBiwYwHLJZ5Y56+OOXn5+D3dbcOvyyIN3k8cBnViR
veotNm37jsa5dtU6/T2G/1SVHX+FhgmKmMK9X4y3eTxGk+hQKTfrRroZKurZUwGq
D8zshoX0TFMrOKZQJb1E7FEwwEB5W98oF1r0I8+2HFKxdeuN6jW8Mzw5qc2oKRfk
+NPAKbG97dvARcjLhxx5e74TBjHIiFfsbQYOj2xZmVs2FDSx5nhOfYXu6i/5FFQ2
OUZTARFFOjmGNzjmcGCnd/1VP5HXNl+Dz7jBEBARZcixrTgLkrrksWfemqyWyN4X
jK1bY1/qoS8i4qPsTqPn3VEK+hfueNm1DccKO1pSx47jGtOphY1d/ucAiI6XUEAk
Wij7MD1u+nT0mKnSKssMxyeguCIbuV0jS5yFd7xZLq4+Gxpa6j7wDwFYbICi7UVK
z2HVYKHJri/qmaBpk+0uh9HK9AoHRpBTlE2qeNl1Q+RCDlADCqng1oKgJb0QdWIR
j73mB76ml2NxpM+TLc5sA/ve8L9fcIrE+eER0ggrc0ln6n2KmJyS6GiKB7kpVQsW
lL79iwejc4xH5P7DcdDjkH3gCTkX3KsBLFLAtINOocjo2Sfu+og2VVVEKx+qi7EI
8oBsUa7vvO2VEXKiaF2LkdS+miA7BvaHZXzn2RVrfrMbhT3AYKRwebmMExzDKfCe
sfh2h520wNUHrpU2MOXhyV2aVSDRXhxeNQvVEXNoguftDAkgJpM8oP8lJuqSZxWn
`protect END_PROTECTED
