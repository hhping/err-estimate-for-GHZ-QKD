`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQeh6zHbU0nlLb6RFlZQPK6McT71Lv1TaL/NEwM2qJryIrHMbPGVHIUs4nKl2BUg
wl2HXvDYurqlaYI+U+wOx04hePfPHkHUWcU+4Wqxc/DaJosg7rebNeCbtSUbg+qp
wMmNXvRbLSCb/VXax+nOMAuq6NEpmIzMrHvCvj5dW2rwWPoqiwpClnmp658DE/gQ
po2edQ/vlzoJY8xptJxNqEewJAAOIvD1JVaEHcF/NUonpEk4gifBAWzRiTjlNSGY
muneadtBL+Hl8L60+hlExjZbjwQbekITvB1GdjG1YDLAusUyRBwY75MAS6P+6lTh
ZTKb3qSSG58bE0i2tdRELzui89i0vbJtrV1s4VshRO7XlZDfLgadECUXppivmDHZ
+IfGyr0xUXVZx5Nz10AkjN4HJPLVcZyG2DNDJHQ+24dKj0upL06DfY0ZD8EEK1Dm
AGZ6PoQ33xUcuTA2R/5YvekATQ1Ew7hR6FttyTZZoPgBIK5fQj8A00gEfr1FkSkH
hM9yP+SeuWFLP0RRVoM8udLIyOHlq+o6dd063ClfBBA7I1uCU5JIo/k1B3J6g6G7
JufNTzPHUOMXZn7ke9++TwhwbsjkTyKqLt0XAPIXfiZN3ggWWfNgmBZdOJ2yHKpz
3t5BdaXP3Mj/LGvPbVqnnpAYtwvIEexsRPKK1G+xUKXYNTG3tZWcs3SbyPTG9e+M
R0hncJ6GShKnCP7HWFPxglIgl6bHbpUHykVLYQVVdVallzemKYkias9pDt/Tc4ww
GcfKt+0yRZyreuSIccRZ81bdROG8gG3P332g0YlcPpNauL8PgSCKZpRguqcIX9Ly
3dfwTCyEGJB8QsXPurbhZ8nX+FEN8k1A7l861Ng3lGq5BIMVMUBnVVFJpZF+ILLU
kTdd0SQkM4NqRGy1AhuwE/t5AGy43iIZCKJBHhxfqPcYtIkAIqCe2a1yDbmbYyQ8
2d8gS4zOVymEmJp7iGlooOJi7HGXUBK/OXhk/uMmHXQ2PrvjKu/fW+VS/aFkeh1M
zgheORmAaX3nrPtTnc4iGILp7Wna9OcWMgHsFj2CM4S31IdpVVZpirDBeDLeD/Nb
DMSYtmLb4gBfKGTFeR+2Vw1PNwNIp9vBRkDYfQU7I60Iz4N68hFusrESEe0AQk86
amVjoqwM81rtD2u7gqdXVBdW1UZXevKvrwmvRadJ4HBjpAWdlIWb+4tmvWq9Oxaj
RCvG3eFSAkj4W1VZnzw5Y7H1K3+9Ovy0U7ZFdkB1WDOOZ5+MVb1cw1jTP1bjqCJk
WbqA0+amou29zbHIsjcWXyOtxeAHhJPjStMFSDMFUf/k62FO9Mrq9ZtlNT8ADNAO
JI+gOy4ru6vhXn8ILqb63rgWlTYA289BQVF52EyVrjzDh/vawhgg6kAGHFD6lUPc
xOTBb0/4cV6we00f9EPE2CpDK/pfTb6yPFdvSUlr78edp6pO55yr6KgaAOQWriGi
MN0fr9QAua5ot5zKRYOeplFHKsb11S46xuGdkDF6AaxreXI2lVMSzjFU8bUn7TFr
jc8CjUiAndYTtQhcohhHdxbxDMMrxH2WS2SqhlCvX5rv/QRridDw4XmB9zy+29dY
TzD/mt9KMbA2d9Mx2xMyc6UjOWvl4FxcGe0Pvttc01E2T3Nksiz17svUgnoAPUQ1
vEYUXZxMzxmxUij2wT07bb/QwBNL8NDBVkLhuXQu7SrMjT7YzT8gyG1cy2XIx11R
76zbuqWFp3hcwE3uH27/o8+B1GZzns1hfCxaRPDbbt90zyiYcbHCNHwaupklxSer
9wsA7huT5taaHxEB8MWVKpllnaDjBIoPJLPFnBgh1Yxe/hJvwLs07TTjlY1oKa+1
`protect END_PROTECTED
