`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/fPtbMP1QgsmDAVjeI7ejT5hCj6errNZkZs2XC2Llqm4lKDTR1vrP3bS0VGvWu9y
EJIE8NPZjDThsuuK4ozXb1ARJdE9HrafRYTArzJKT50oBh+H8JaF+kgJFYmylRoq
kpn+DbOaHRKM607RyQQ4F21QoUOuie6rk5P3vVNdUbWg+iXfYGrYZO3y2toC1KZu
q97lnUSdbdWbGReHyAXAmDu8dcAisuOzgUmUhyrOpOO8AM5CHQLzaLRa2kmw2YU4
qZL0cIEGOPtD2t4SHr8MlafGTkyM7LSqB3+OcPg2JLvEypsCVHF6T0b80DhhL59K
GgcERe/rbQrhvknKcU74YrIBgSFHsbhMvTMWp7wBilTMEVdVWvdLXYahRmLArcSL
JipI0MnJUO7UdfH/PDrJxOYGczTpk3hY/hiYeFhogrI9fk4QGuaNKH7zwIeTWyEx
k2Pr54Z5MSrucYiC5bh4qFeZjAORMr7dQdub5ZSp4d8=
`protect END_PROTECTED
