`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klnNEyOR1oQJGl+91q3y3e8GXlUK6PtA6WYBQFiG+wa6JX4BaMAWZfTngXFKQ5Ms
lWlTYEzA1rrv0NhjotY9E9d+M7yy4H+x4bSyoGTVeQQl4+Y55YF+gddnelCm5xIv
fbNokBMt6X1hSbT66vHkIR9HAlqwegF3cfPLAVQKo266B4FqXb9TuKIY4ZjyIqzP
bvaQdUUjZee3v5kP/rZuydgqVitcj3mwbvhE4vVeE3gqjoYJfHXcB+GD9xvpXecr
zOaC1TMR0/1VH5wtdjT+qd13Rn+K++4EOIprqmYNLY+MFC/VluqSZxwckGvgicjF
zqGaP8xUGhnMT5U/uTfni5oaRDlEPejeB4zE75LeCcmeVdf5h9TLA6GVQChj2bAJ
DLTlK6T/0N8zHSryNTfkxC7xQhv/XjZNa1nkaZ/BGQ5lH8KYP1T7F2iZC6f7RBo4
iYkrluhdeyqMZGhEprikuC2lmMMYk+SfU3feXrsHrizwNLwfS7AxofJ7vh2Sr1Ls
QQbyfEUc4XuJqljEXAZZlOLds/a5JbjlaJ58x9J+Wy7T6aZdAzhN3RCX8LpYhVDx
mySqv1UGKYtvYUgOqX4EwEA1WfUYhvqs5Z3TPp1RhmZZ1h1iE196yZBm80yqg82a
BRaILC2hDCOEH0A3eSwUMN2QDxpGUg41F7cvMW5i762FC+lDwvfd8cqz/FqExwdq
HRpGrsahIM/XduojPj8sIbbptiw3x4iPwzKdGU8KLqP1vBL01/EwcvPBSZ6EjaQu
UbKwYnFy1Ruw1Ef7JTCtJZST1YaOIAAJJxNhPC058Zlyouwxb0uK2Jvue/grRdy5
KOKc19Yoah1luP5teNLmcunv/m0wE1H9ET1t1RGYheEq9FD83gFwuK9Ck2Z+GXDw
elUJ5jFapSA/yfpChEvX2S4ka8Bsfds8mewO1e8a1QcFQceVk5KL3PBDD21PyPsZ
o1ySxrmZx9Orwp234rNXNGxv6e4RvVa8NtxV7ChYRLI2kpMl+D7Ac91MCegGBJQo
c9i3t+hmZA5Zp30WmXFbtaFxwjZZhExc9W4N2ihFHh1U0uFa1i0wMCGaCryh6D1K
c9gvFf1yhFa6BWzW9BUDthU70qDCGwrs10q+uw6lpn1OcUZ8b6mU2uSl902t8FMt
`protect END_PROTECTED
