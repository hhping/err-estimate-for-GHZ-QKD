`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+r9TChD09jKbvUneYKnU5jRVfdgRuWrUbS4yPosNhgG42QRn11U1IQSuUfBigMb
0C/Ad4aL0mBOCc7/WWnAFpwEJ2udITYq50plRxZEsmZYN195UUDYyVyD482Xl4L8
D2hgnCXY9nMF2c+uLLp/UQ91BmRlBKoQ/T1xIWqENuaR+yCeYPXqzirGzBR+KMcX
f+bN6lgMG8OG+nkZPJucYBCsI7Fiwp90x/Stwz9eBMm/7b5jXx6VztcKXkOVWX7S
UbsEkieoHN2ebawaIj6FrohQyfbE0Slyn2dtrjOEeocoLYYvdZNwwrep50+KaN5Q
6hLiIakKdxM2cYp5g0/HHz/6fxkLpTF7u1P2sx1C4cNPA0DU8XOyDa73m6kCmzaa
kqco4UUZkBtJsmWOywIlSyWyoX3uMgrQsYJdTY7dIFdKqYWDwokJntu/d0xaSn8+
8GXgpL5LEXSHofL8FGI8odU7i5AODoDH00WrZGvq2x7XrjdwrLrjO3e+8P5InbC9
BgTMuwIVfVrr9XJWq7rurq3dPjZQnDLYo1xVE6rySW93xoylzGcW1PQJZCkgeF/0
s8IgoXkUpOnAngnGzwgAXg7VWgAFvfmeL8eIyfJbCgMkQ/aJwMgyaWvOBiQnAD/A
YmpZSe5tGX/1CfklLnSUUG2679UqEyRpokXk05X0jmSPyPnuv4/Dh5V7EwNCuO4E
qrmNYjx3vrPyqfg96yo/LbXlDI2e3cjTkVDdtw5rm96O94D9AbdjhIiUsFS/yrdU
w+p4D7+gAud4TqdMeFE/NQ==
`protect END_PROTECTED
