`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZjL8t8KOwlvqbKCPCr/EVwUjfDAbIIxd0yqVKhu4XaUUAsw3oAPSEbzvoaV42aZ
qCz2Ax1zyIP4hbxSArBTo4FpbwuU+lboJ8Pbe6d/iZaqwc/4l5KjYteCHa1QsWm6
OQapqzL4E+mSp/4KVFu0h6DzYBi1PNFdLUzavXqbE67SwaEUwjjjr7OxkLJHWlyG
5B3PgfLdmVic0B9p58U/XQnb8dKkiz9GgZZVBzEly+DivnKyRwqu4sZWis+kRMat
y2nrr5zbUthUlUYNYoGHpeexeodf4kT7buJ+iUA34qoY1r+NQSgDkgEwPwso8Y7J
J9HvfcCiRMDeYrHyCEz1wUYReF9Em+Jxf4vxGFhianxdYvFTNI6cmEYg02AHJ3sa
f86TQVlfsjMxWveS3SJxop+GG3Yh911IP1jmKRsC8DJTaYgbiVNDbWy5hGlAyIUp
TGlvK6t15svjWEF3W1LDZPPz+INdF9O5L8m70sVGYxHpW4lDu2BOVL2axX825zld
99SoYdi/m+p51cTZnw9IPzXaavLW88b1BnimiFH9lzqh15mV98WxLnkoPBruCPcs
hYMZHYXiXKsSRIXnmrATuYpNWHmgTGXNfp2oCfTjDKlPavZn9GPCcbca3iExaFym
AZU6p/YlJrllNSVvYEcT+bjelq80wz0BvNpG9TVDNgwLdo4qEtMhkpnC3DuiDZhk
xudlwC5p7y/5gd1wCpeNZpdrMnYX6swWMDL3Pv2BUJZDdFeVN/ePX8/FQho5Oywy
sBg+1sXl4nEuMSJVMXoAFyJE9ALaZLLsWEz2oEDe/Aleh71ybGQ63aO8jzIfWRYy
gmlsMxxYUsIe37zTlBClAhLxbrS+vpWbti7A7ECJ57p6HT9Db3Iz32xVLR5XYOtb
PrNXfPDI7rkYZCtDv4dneASM5A4b4B28Bc7w/4hdgOomyMkqwsEypkg6+Zj7We92
NKYK38dDok9/laLTwJduuap+hTdziQUv7vM413a7ht56Ew9+WvZZcqCP9BQYlbpW
xOzIyTBru1aLmHDa7eH86svkG7l/Tn5gEw+EeyP4dXdfMOU7AwQO+aCA+1k8Bjv6
edX3cvUqsxO+ADn1h8vQlzj1XMvONycY3exk9vILs63D4HWdwAeMXYKWby5MyHw4
+iqe6BRefvJckq+OFqOGEYPJPfGwTrVK263+fq8QTKCk3K2Lq1absf+AGJ18h5y1
FKFaVxLUj0KOzvykQ1ddoLXWSLVdVRHs71vY+lg1IRCtp/bqt55sQFwliHpS4pqa
iStupGKgQw/N1+5SNlAU9A0SZwF+b5VVoHEMRZ5xf0/2PwGmkWftRjyIbHaCY7vB
BkDMBFMsJEjitTbHsQXh6mzitWYz41VM27iK6iBkQ1IFVySHCjLB/oJygJq7GtwV
MgahmUgYyhyA8bLn1zrzJz0p/fum7jBUhsBsxsHV9thvl46gOby2W1l2fiFJ76U5
66rszV/3JJ2DDnkZEY75UVKfuUC3yRSUX7ZttSBqxJc=
`protect END_PROTECTED
