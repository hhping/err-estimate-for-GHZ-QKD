`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0PUHTRdtoHhTNZQDCdJe4CZi1VnobTDar8a8bgSxp2mGGHH+iaD3/66vGWyo975
zWX35w0KryRbzd/hHN1FSNG31SqYyEoID//q9HCwxJ3KOhqtKH6Dob0IqnfHvV36
meebEr5MvliNUNsfYvX0b2Bv/akebXMa+YTrds++sAWGO/f/qSBHYZ+hVuVWFDv4
xU+mtTDau0p1ONN1FC3tquOcaj1TxJpJDRCVUqcaiLFdKgsrkluj5UFsFdPRRHu8
SFqYVXBgwS/Z+y6u4zEbDYhR2kGKy36KJF1c/wMJlZArYhjDQejW3YeTgpLaQaPQ
Rc5p8SkkFdPHf0IN0+zWsoGoAVd2Gj6HBUzpxpzj9GuUN8eg+M9At36Kp50SB1cy
xt91l8T8hJe4YOPme6UxLtLJhgOzAwVg5PtJ6+qu8EVm6VC+4TEaADKBe+w5Ofyv
7UqZVUu5wnQ2G2TIqA468heFI3BZ1nQwtdsE6XpKmv9J8so1QP5gkGnHY/Tk4Kqw
ZxLTdrgPhO8axmOnyrspuEfEBjVf0BhyMhLF+h8IgooZNJ7B5S+eWBugsFqr/JU0
LMwN9o2/0hn1jexlnllnlwNGTc/6AXqzJtfvFD2SlR5T0+KD2Rj79PjrCNGE12Ex
wMkvPZhwtjEARd39ieZA+e6DbMssyjfweOS5eBo6EfVVsFVe5HorQU+SRGpSLUBa
exGm0hJKhamKkf9SRZ/GuDyGFCX3ZNSztHEk4C/bxAA1H1tvdkLUq2r5uiSNFtNf
4otpqQU5Xdu4KZ/aQl2J0XHmK7dweso4c+UDHrOZrGTALXcKLypXBwNjvWWGb5Q9
HddnnyPpaqKMaBYj8xAllFocG1VSudiMXEFeovwhMeE=
`protect END_PROTECTED
