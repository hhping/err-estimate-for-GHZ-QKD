`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1mV508+1mpsaZkkhott348N6v4FKS8zlsCRBFAJ9VTAiyuo2YL7E/FvJLeVtviv
0nXGwB1KZLYb04PxoboAOKtxzMkXvyIGZkz8fUYKR/OhPNlW2OYUhh9vblsl0hgL
Xs+A4blWvajS9RE3uNslNyU0+h9HCYXk/q6cpFIpQqWk5jbZfvn7C+pHG1dztMj6
k4brC2m7SHmwea2l1ffzFOdjoMvihyeaME0Em3tGyW/sjaaiNOSxXBWD7N27Pfh/
raux5B5DFLHM4+I7e3FG1FNszGVKmFX3PdRhewtrroo1CLkL5vcHe1l3RTt6ggcE
bydQm59imuhqf82Hi7DZaf0tZArUWP4ujytLLCp4MFwZTDEpSTBXxATGmMeagN98
DHKdYDOnHsdotutdWkHA5kp1SS2D3ISSeXZUFMt3djt2c6dyuGwR8qg2thK0AGZu
XyDNmu2hNZDYr/L3xJLK/i9wxmOaEoIC3m1X8a+o8mpurt9PBw9LDM3dNIIFbu7E
U1qMPuYyAs6wump3K/sGa8/XjbgUA/eX9i8MARjECMN9zDF6KQYgfDkyasbsCDAG
2WwW75uWmJZxADayrERY9ObrtG3H5jQSIxwVGJz7QYb/qmUs3fJtUNi1TXg4QNs5
tHPRf0j+uOykH59RIlBCub8L5MsfsC6qTTbwgPOvoy3FWqIxSNq6OVPRibZb8Rwq
2+GSk61sUpJ6Vx7STO2m2XjFonVFBel/+fkXtJPsRl7/Cm2ZJaY6r+7guyGoagGz
uTPadWyTt+mk55RUynH4mSrwacKxfsWaxN/BE2gqCiyZsPgKHBilD/5D9SqTD/5R
6MAKXDPe2azg0BL3+rn4HlefCUwaRfBnVd5wf/djipwyEbNOhpTDAyoHavUbhit9
pUUqDs6m+xjhLCsx6MucAx7ID/FSkoYKRLTW80YOehmtu0dq/NS1ae7Yhs8fK+NJ
jxOASYkhCS7sn2yPwbJTShwWx0XyaefT7JzvNhaohhzdLvU73Sdc4BA1VN9Z4yil
VFQtqotC2Cab0tVrzewhisCINVnUPM0hRUX4MzdpEdBHtvADBEREikz3Xc/m5Ymo
N8opmUBq75StR4KYYVjwnSv1ig+jS8Y+P79Lz5D8YVS86J0Zkff1IauiujW/ehmK
HEj1KmFzrbhsL+QoBxSoJjy6uUFFZvBZurYHDAOgGkCjytOW0y/9ctMcrY8G+yBv
SuGd+LKsDUO/vjCq+3OuxYbEYiG7FXd3vOLNCGKzMfhLXH/P0PFxkWd53zprmhDs
V05x2UhbXzGXP4I+DgJaBCu6qXyZJbrjYoFe+9MtTagCpCcIUSEQZyzG0dGlKG41
ltRYDTPK+3wsA0HMJSwA9rcMMn73JjrVlUIv84XcJHgp4iI/wSV6LuB825+h3Nkv
FGG9TP5ioqpokXxmQr5yHi7D+xLbTwHm2NLpLVh/8JSdWtCOHdNa2fCB/DgZ50DV
oUYPxGkvgGlMFwYeRdLB4Qs5GJUafk9dSEDT9c4JpmlU0QG2ywoido4R7YrjwQji
E1XMSvMdAFerdyqUkjR1xT6oe5pgTu6Q5Mc/P9ZKITbTWdbO/IsJkKnRoC4c9DpW
L4JjG7aemNOTxdZF4zBAjxmgy3CaIQl6mPIV17xDKy+IOyfItUzW3IwlbmoaKKp2
0qv208UVfX3xsqBWursvIokuHPbdknhKmzywVZS/ngUPECVd85sR88yXJcraudVv
i8dKuqD5aEvxig6MrClZefDX5rBOhch1rOec1OSu+NduE38fZt4zokI1J8J4Xg20
XA6wnYpdQDKbKBG1FE8LCpqkB31Ywttuqtd34eHDcnnPgfZXIWPodrmjz5t9ffye
GD2dq/Qnp1Oy73RMs4dP0aqmpoWfww6zz5BGmNzyzVMpETO5VksHMKJ7NRW+6+Ug
1t3SvuNJsTKCuyiVKI8RcIprrLi4ozAdM3OGH4Ti+spWZ4OtmEZ5GTY7WytWwPM9
RVp0QMwXhDcH3pTe2cG41Fjf7hKtFpFFMtCBrr4XwmBYGj4ctynkSlyT4Ftk+X9J
BjgWInr/cxHivjXOsy9YEOreL3jwIQU/z3KqUGaeKFyU91gUC/NvIDIjslaxFWWd
hPtJ9nIV3VH+YPLhawcpE+TVuRe1haJC459lPTjPRi+hxLDVeladsapXPw8VM3gH
1xpuhPE2TYzcbZDpT3E69kDFErI9X+8/yaq6Ornfoy+k3vmQmS8jMA7JglCpQBT2
AqYzdzm9ZXgfQpaBADQOJcDlJmmf3XK8Xhp0fsB7XSD7NA0Qrranc3HtReDeoM8s
e0ZcQgcNuq/4M8+LqvZ6WgWZ9THj+0ENtw9Dcx/DTApfY8yDXJ+Lbl39f1DdYwU+
mrmZAg6FAzSFS6HI43EycbtcDO1mWUXO9DxE4YBH3QtV6ye+1MerEkxSJrUJKFtE
o8rVUQLWzKDQrlfmmZx+MYZ7SWQdvQ/IWbBdaIDQZprKPJTGIoQ3DwB2OWx+un3+
0NhAs12EiNJJCMAzkXaSGhhdnlE/NItvFgIpdOR+IZyP0Up49hmaLLJjmWUSlONB
R48h5kgbBnh2Mj+HLgbbnXlZjNWo14By+xVfZmKxd4OV6VHdOMsVFC6XZ5BxCZce
PvUJb+tO8EVJ0lWAvxUVkCKGej9G6HVxmkp/HeRUHdjtLBBZ0xWguGE42/X+gjUE
OiBv9TMBi6eo0ClhketIaCaoWizyFMUxBgP4nT62yz7juGqj7SAgMPdufcphRsz9
C3gZ23Se1y/A9w2Qjv1w21ayWi05mOzMwWkM7C7hjoVw7UV2qyyEoVqAM71PRtGi
Qx5YG22t5kh5tEPooudm9mJ3pis+6Sl8mahOl5A24KQaW6Y2Trf+tQ/YzZJwT5Oz
qtHZ6emU+dxU4nlX5yJkZhEOYt1DU2HclAddkBi0kFCc4bgVIwL4S/i6wCU4k1eD
PRTYeNDB2Xn9X3hLYVSBpLyb/EajNuhx4vw6d58HiQ027eizEFPjana5+oB4CZiw
mgXWqpTvC0Lw3GdgFAuOkvl6ATnNPLc+mXK24qtP9SmP43FIpzIdhTQuTykMuSbM
WA4Q+zQMUMa/BlLYt/VarAqIGNiLl1geMPpXGWeuM+vwbKVKRnOaubpDF0vpa8We
Q0HCGzzXUMd7LP3Ss+vuP8WJC0g1k0mTd9mU6Fwp9Z2djLvRKd7PWv4grZ+9tWVF
7MdvQnmp93e4wTEyH187282zS32z+tJwIOLLw6b3AuwMBM0kg+XraG8YMEz6MynR
XQphVE9vkzzWwFuHM31S8Xe7ejiP1gE9MIwsHXEAiGBeIoBBN4skCzG0K/YfsXrc
mwDS+MptDnN8tdVvndRgKEBYrghjoL8aVXc+RFK9sThbDaxsxI8O2531y6z111GM
dtY7U11CGmWtWTxxRdDLIwhppxHAlIM/0Ub0kvb90arGHjUwcl8UraLuIJQ6Giy8
+QVIgORmhKgwtoyCPFO0BdRfmXWuWgh6x22s+e3FQEDKZZH1249T1TssEuGsLy3Q
U5ZZg1/Ri42cr1XAktJ6HSCSfoMOaKYvZOOIfF6cxjU+Dv/EiAt2JI29+yQwVPQ/
r+h45y8fM76rt0Go/0ayTED9FRecj8v7jPM0gSPpyoIBZqMkFtnRdKgi3VyyNL+b
E1CDGgDlbaLlATVwYkuInNgiiT6GI2zEwwIt65ZXu5kCiYa4QYVqSk5o3eOjmupW
fJp5ihMo1Ipnu71V7gmaFg==
`protect END_PROTECTED
