`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UwUnhWewz8icvBgVVtQnzDYEVy/zKePFroSvGr89ONIF8dVItsVyn4WfMRUEz3k4
l8q9SRUWlKYRCEbMxqWoCWItDTfgqkFYUjcfeCHmLUuzF5jfWkGJTYw+cVprGheW
6tc78RGbPYkYiKybOFvreAbMUXWHDvKap/bOyEN+ulNdlT9QoitGedPTaPUknJIY
N7XNZ4+3cmfLZyM7/ux1kSRxE5JR5SzF1Jxo4m3VvzGrv4078HrmC9T2CTSnEsl/
hRyly3abOQGVPBFowyyhVb47vt+RpXANjColqFK++JAvqeCwW3mMIH+9SChYRcJQ
Ja80r4F6GRK8PB/X193HKwIdC4b6BE3MSJZbOVq5TALZcjyIb2YTNhXnGJ6ubyWT
+Kgkj11Ekc3cI0uOtNKkPlNq+YIXOMutAfGLVwAEZmjvQyB0oxlARUQDubkh/lag
9eGh/RNquUeAbx4smcRnPVIbNGncTX82zfRXACtIkowzFkvs5YyYq0TVVZD5Qaiv
kGdmJ8UnDeH/OUPCU+f7dyHrHtf4CTpkWm8mwjlt5M6ZCdALMpZQ9sSI7wU4jxHB
75Oy7adXPYjCy0A5vKy/czhFwkWI5wEsC21Z6/Ini5n5ITXRfx1WP06vKhWc1V6g
gFh6frlilDqjDEEa9s+Nu9GXkV4wPVfmPPTEpDzAEbU=
`protect END_PROTECTED
