`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UKR2B9dCqHhjT14BXectUx6EzoEcTPtXvZr52F0fy2n/r64RiEB4k3aCe7Dv5yJQ
WwH501EY9ivYPSci9MG3e04fEsQO2OI6AoovDoPGcCSPs4YUfjTQsxakUoHbDvea
pf9Amvn8BoHenuoRFtk5BT9zdytZqngsky7r0zspZ8rE1u6nNDmZDS/9G/NaJAL6
lCbbSX0ohSCz2+VTz3n4GC1R4c0Zq/cvosiAcrREWGA9Qf1amCbQXWUgP3Tz72Kr
2aeSzQmh3HQFP0Pcq1oTy2EfRwfFtdR1AbCqhZ2XV12WEx9uRqcnWlPeVBE42EQQ
VHhf9AOfQNV3deqB+CxcSGHwSqxhiqwKF2bn18RFVC/ffaJxB1QJCYIAHq/uxkJU
Y4LsMGFRIXoLoovmCsPq+465gJwCyr5majDwiocO8IJR5/FAwfjl8c26TcVw4Cyx
ftQSPOD0gRmujMZIebdlP9lnDABA4zX00Qz0v9txjBDwUCgLxJSPFSuC/TeIWbD/
czjiEeP2QtiLwzLJpo31f6EQ9H/w7TjdGhnkrSS3Nz9sK3xvotmmQinuGVlyChSJ
QZPW+OHjrx2sjiagIWJsS0oZjzSI6VFOrh+TVuMeoFtdLTHSljrfkD9hFomC0QEk
`protect END_PROTECTED
