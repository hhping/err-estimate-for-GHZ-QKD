`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHyk4XmpSYo1SiEjftZRcPIYGnQ6+OckflZF4/wWL6jLqqnwgNExoNEeZroJrf0h
4CoLPKMz06SpcMJubWKjOGO2HpKLdgoYE4d6MNkSld/+pu9Bt6a0AkIpGCMIUHit
fcS6H4uj0mblDxgNa+e5SodcWGsoU2Pi/2L3l3UJf0/+M4pZnBf0iNzHv6KexuMx
dKxMCDL8qAY+gGt+PudNU4OFpe9FqmtDbPDSN0DDfGd7bpaf2vi1qN39c7tqJGl6
1JjEjI+erwQf4dJpgZdpBG2piUGLakCWOhO8vB59wVYZaUxuPIbcG3bTWnuRXKh1
z1ZHM9SflqaO352rLnTGpb3uQdwIjEXMJY0r2C19qOL5Rrh29eYFwRwUuzWa3AMe
iqlSjIYHW9hD8/l2efH6R8Vy6Vsta446X6eqkrcB9JrsgvnHt0oKYf+LLI4DDb/X
kOYGY887EaBCUDHsqkNgllbdIaN1O2qPIDMYITALllasUCTW4VexGUW7z/BlvPf8
3t9v2639OGNt7Hc4f3lRuNopbsuICVOtyZnVmX5dUVkylEQ02ddeV1C5JHbnK+hr
/NM1QulZQGVtpBFKZcBXHlWdbK90Ht20t/v9wDr36tXUtrhl/e4YZmsMgwlXqtuH
168fMZm8OuxdQFPvU/sw1Ai4wLcxAFW/64ftQ5c6t55EwPJTrbLBRnHFjw1SAvlH
N9tPjkpeN7+1Y0Luhg04rwCgYBP3vCkPGrdGHA3lbGT47Iot5AGQtrXRL4uyuQZR
OZ8yhZGnkK1ksau7raQyzYfn6bW8FXhNTIZPyXSEHxD4E1pjVL0z4NEJeQDPyx5p
llzKTGKqOvpc9fCCB+ZlxxemehmnlVPBEKZKisibAY1G3t4b8CReRiVy0ocEQaAP
TpzXmti8bl8et8aaSCXS3ccfoNNBzmRj3DiHKqVBlvWF5G57v+OsTQnlME12fN7f
cHn/YJaxYGUOyzYWjtgW6u1f0q54BMT5RZYlq45hK2LHJ2Z8NOI7M3rjcYF4/VAM
TUnKSDbMRezTpsldRoLel26KWSP5KZwFZ4cWNXWQykTUTn9NVqAj/iEmKdgJjzCM
QeJ3uImGUAf7Q+S+c5ItVitpv1kVzxIkwf/8Jioyz08+9jiJLJQtM8VOU3bTOXu4
eTq0xZMy2qhCa2fugn8XsM28nyePBaCJ6ICMxpTUIVo=
`protect END_PROTECTED
