`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gMLCi+8i9M1GVZetI8QUe66Vot0bG9BDVtj8r+cBNJMt+Je46hAQC/NzvKe9Rvh
L6lkY0mtqVzlB37KN72BKP4qijywadBmKFXtTZx2BGJysgaN4usOrecnnRVqQuJ0
yXiUJQOub/e6jatzg4YKulbFBA3hbTnvoCX3LF+kXCRB67TQ8G6VC/YuD71rZV8h
mHZPJSnlmoVxA9NN7L5K4OB8/QCvqRyrKduynBv1YBm0Bzu5a4Tg8T7UAjKF1kEC
IhW5N1b68KOttSY6T3Q+3dW3QNGPDh63W6cUgn8OZyBHwr4DFU1C74HxCEmsykg/
Z9ttlgeJbn6p70uRGCQKLv7zZ7nwFOQrgsQd9blwUwc6RJlz+Oo8YCb23LvbzwAm
IsBonslxIOpI8ppfK+mOtMiKKJqZUxn0HFiiOF2Y+bZ8TlQ5uHdMt+gd/Delj7bl
v2Jij94VBXBlGIbkf1DBSYvfzIyRPq1hUeVEiaBTS1ivu6I/ujOH+JwxiCZd37cI
iURlZO9F5KaogtMy6PcaPm+4pjfTu/C0O8qLnDHCts2i+MrqLtrtJURi9FMqtSBH
7IpH0Sm6v/OBjMoVbrbGjLZD6vDBmo4Z1Lv2WFMOJpemKqlrXTXyGwzuO6NajFeJ
9SJ0JTiW1eq08cvzKNK1jyDZMidp9g/kehkKpHgJOjqdqKz9IG/y9MYNDXWGQEQj
puxYUOEZ4HnMcu9MkwOl30eNU8S+DLOn1FZv3v+9ypPuBsGG67wAbD5aa89xLZvU
RldNRVU83ZyOXufQTcd/TAHlix57+MleCs/zdt54DNk9dErQsyQoLq0RzZv9XDRN
`protect END_PROTECTED
