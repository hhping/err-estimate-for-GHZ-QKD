`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ghHOzSufNcT8yLea5FNIrv49eQ4534FbH1veR9z74LsdFdQPJ30rTN9U3JqRX4s
UeQCQfY4bqG4g77FiOCt5DxjFrC2fkFotQ82l0KP0F4XupySbBxtMQcqeB6EGkv5
Qte8LFtVnQjkC5sdGj2z66mSFy55fDEa1ElQTbiSphyTxGokvDGfNnBgvejuiMfO
nfC8UePWkxwvgQrVorndV5mcOu/pxfI1zb43nvriiNL4KTEts/+skQSTMrU/wmGR
LQdt43yiMK1c0xtM5kzC/h4DgNDKkpyIzYWuCax3NNpRPdfGBrP/+0LlpH0LaOeC
VXYodG03/S6S4c9zb/Uvjs3Dc1sTKySvD0KoDVOreB0BljXXmvjNekx9ndoWKbbe
gXP/RqAafjIPWfD2TICZuxeYOoDI2bSWk4YIX33kwsNi6+DP8f8/gB15H8z5wEtF
PKSvb9tF9l2lgT4WEj7uKIQztqxWveAzEsDKfRK6j3RMdtaIBAYhFEp2QN4zAYgd
GKYoJwT7ilphF2I51DO8YjFJtUA+AqSMaKpXWMXv5hSd63sV56qjmcGr9eOJZMdz
YHhbaOA9vt4fxTDIJ9XDTcYu0bXJTOpYcPE8qisnApbISrpeflBKVDY0raPgdb+s
jnbT92thYIPAkEtWbltqIUhwtUeka2Am80SIyYcI2YNVBE6hZfC0Hm4L08065Cjt
P9DdCRMpPUUoc04TvAoIUpUj3xYwVIGYLY9He7kJxObxeOtm+5mWmbDTNEG31JlX
BO2JqgdBV2EEpriIYVHGnl8JViWDsybLk9rrLavfwqbjNCoItU4os63pAih/nd5+
HGDDiEeWobqO1KBpWSUMzB3tVN1qHX9UqxMWGcGJfL74iabQfMSvOEo2qsLYG90e
BbphnezucQIlSA0LBH9W3E+yOx0GCu+XJE492Rs8e1/Sz09qbZKulfrb03hIJtA9
1voeZHfwKZs1hEAn8WQKPUo0Ih/96vUt2OfVJRTGxChIJ0zG+xafn6KnnoqSKEEu
gdbvODDqai2d0ZwWSRVDBDurDA7uUf+Bz5EJIj4cr5fduVQ1vr08ieED6imol6Z4
4p5iaPp6uKUBdg9q/gSCYTR2xb5eEj5p7cMjG1WYHSWkJV6/75RlGSSC40MIUtW6
CxADfegYzNUvdjGbON2zQ3bRhqWGUj3y7h9rI7HMZG+Jc831BSlGFN5IJ5b9T85f
cJno8LlknFo1RKupzRW/a4IwPOfqw/Iv+ivH0xMcNyEDx+Vc5fdOT4zYVEs5xKDK
czeKWZcqNiPz/YTJ3UPvjEJEQXxMvJGaO1qcblndTxmtsyPXK6H3SRq43st0GAyx
7eg61ydFxRYjT1QTNEhT3jByiWvxG/R6a9Mj27PPiqQrZrHoDgqZ/uuFqM9NrHYI
NI5zOXUGfYtXaritLrNNEaGQvojIEhl4Lm/On7UnqD9jCsHtv2xCHlFY1If639d4
dQ0Sa+7SD5BHhTN4MVK8gjpJ3gfwqFGRiE1HQARHowuWIkFA4oW8sLxcj//TDsDw
FkygK5dpXBr7O/7MaPi/2kdxSj5hIkjSCYJ5MEGpd5zqMm/6vKX2lKos1lj5++TS
wmYCwHzdsAulWt/e5uLn0B6ISftTble0PVLU6BTlWyaL2xicqi+F+Br8vi8MDuBJ
3TGYCdMpf57Ne6xvvuiiWzSuvVw0MMlR9uXDEiLhgvxcq0Aaqh6xc2QsJFQSjZGy
PTIiA8Y+EwKgeBLAkVe4rlb89/7YeVRqUkR9U5ksaBGpGD4Uja5wGdp04fXUbjD0
IZl1mja8UK0juC4+FfKrapbIElbicsxu+kFPCcilCDFnZeNKI5xb/LHrTA8C3FtL
hAYjHhxKdHsKw8h7eHhCKR9R0sdmyZZQeBft1ydrJXexaUyFLIvMIymjyrnQi1ev
87DLCCIYE3Y6fRJerqoXcn6aV6fHKMNa+8LuFc0wQYEOnUkpIEAe9i6WHQc8c36n
frdu3TNCt0TuCYo5EBX7rfv8uudB1pft+Q1LfJxfyxfsoiZcoqEcgxUk/+5bUB9J
n5Nkzmuw/BQpOQXXH3wmKUXBpevCkJp/zWHHh4UBBFyqgjqeOKjKotEbVQRMfe9J
7wCYc0q6wMQUrrPcjvcVJJQNSAT8whr3+WeKU7VZkljj3mY0pDja9kHwOSC9B1UD
J6Xd0gsOmkOKTWSTRJcFN18+UjZ0nBgbOiVeDENebD43qWqFnYBkC1mK3DM90gFw
/FZxAfLOzkxYJRSpnVcQgsjA8gAm3uA3slM79fe/3kdi1/xWtjGTXsCJwIRd7z9D
48U1473zsaHKus7psgeLfP/cDBrjN5jGg3KlSwO5okBWQSXHLhXE8S6vgY7dqNu/
f6w7I6ulDuEBUYdYzqwOyK3uOCwVSlPTiNFVr7UaSf6OVzlqvyCUMM2y7ZHUMGkj
QUs0GHJvnpfJSsiZxJAkipMEJOXcCQXNRTuUueeebHVqt2JQEqVFcM7ZYlyJOFV/
g8NqUOvvchEkRQwr6mMmep2cLRHiAruqHPPUC+b5l5xM+j0kqd3+TU0oGeX8REE8
Nor9+9o0p05qeQ2ROqMt1w/IvqLcL1DBYUn4Sg3clpGE76xDv2TbWy5SEwtukFj5
wEv3B81dXhblCGuNZmJ1Q4F6kL/0s/MKquvP140FHv69h0Dm7DvgHzFTh/LLIO00
Q6mH1gWHiYitnBet3oZmIL18RDiNHP1tb7crSYWPcEa+EbIRABnwE6Rr7VgHbeX9
CPFV3J2v/y8tGhjihh1dzUXm0+oy2VwjG5Dpkbu3CBrB+dtkkZ0a7Ojudxk1pZjG
8r3vzHOFOjDdj98E413YH8PNBjTnGZkL9kBwfyvjnSc7Fc4QpF4znxrkrbu7wJZV
dTjFvSCFyl06jrwm+YqixButK5Ndeoz/vrVx9do9ZxcrTlvN35g7DCPZHcPCrv80
CneG5+pt+jLEGRliru1PEnWjj8a9fMpm4QswdEFCbFOQA8o3jq9TgC4Gp30xRtMg
19lMzjGWz5bXjZ8lizkQBy4Uva+xPd2n7mcpCeZuYNlfWZaA20CRZ+c8+HnvOy7J
TsGpLyWhyy7XdVFevMVk21zBw5qz2Vc4o4Va1BEyvsQwLlKNtoj7tRbL8nZ2QJMm
XGQeF6oJEENpNFF0fvzcLy1Swt4eobnWAOwztbJlnV5EO2+7zCaiRRv4GZCzFsWZ
KuztUdL1mZShjuw6t9uf6wOplbL6ccYJg/CZFm5iITesPeNiosVVXrUnmSbB+Vk+
tBgxNu00/R6dgWDz/AZEkhst/loLt+sSf9aXVdSbRBZZswMU7Jeh02LtGCsr5HtK
4BVbhDd1sQ644PMeDme2KSwa9R0TZks076sWen55yxD4MMV6DQCKFgpg1+1JPu+R
iQmK+ZVSoWAm9YhBSHVW7nyvIsMcbxjtPh3AVng/VZ6ZFyxxxfGEt+R3UNoje++s
W+tPFQJMCQ7N7w/afyD0XqK6AJsnVX4uJ4dUGLdNvNEAlzWS5SWM+zRALnFilrdO
8/WVYkUPw1qraGNciiBEebCO2z9o2x5dumZ477vla8kVtMvzYwv4FLhHu7Zaufr0
zttwPsud4yWU3c51+a8PFfRaJwjBm5sttTb7KZAlRGMd7AvPIFpeQ+q3VPDHP4/I
eCm/GbbtQeBmz/0dy3R3TL23HPndxIggrf2wd97SRHM0hYUI1ZLDLjuYtyTVDp3o
mGpipwTo0DadMnP5ANLBGUP4i8d33VQkz2WwJSawZJUG9V/yb+kin/nkhTSs5jpU
vRkU/tdGz7/FC/cvMafFS/y68Zdt+CmXPVdzmkAfRSFQsDRlYLf+XT1gYib58RHY
gGLIocO18ERNxScsgXpvsGR20fmIgIBR+XNPL1z3LiLFmU3ACpVgOiCmVZKIKS1N
K13vy3Qiyle+v9l0VfZBcac57Aqq1uYI153Nt/COVxUtrhDk+gal/tDqdLSNgjCa
gQH4wycZ58odn3T222T13aOgxhwZQRT6HXwQkgax/9HmJ/QqY5iTK3sM+MVVTd15
2jNx+ZEAfgZJ6B3iWD2h98mrSygrDchj69E4Ub27LzSA7KRUKvnoZdVQTL2JGrkY
LTKUKwpwnn5/JurcctDb3jAm07ns+dm6f/UEpmAuDhtY/daGGGEXlcVhgfSxScuU
vpJ7OmauMz2VXy7iycjg5J20gNfaHACnr6VU0pNDRw8r/rEfgllYgP2DXEEGqZYo
80RMr/hGoJYKU1wxnDMKJULdlq8Jmtw6zXCIyjBv8oBlay0wfjkar6ALFppPOQpH
f/d7tcH4pXuy7ykBdKAlclEke/HO7F7Wz1AMmSt6roIR9yqylNaAWndZoRnuNJrA
J/1FNCRLDLzZi90VXv7cSMyEB4Va6p92Pd9SVvxHxd96CpiER2eAuiLV0E7/M4gb
cHirUoMlB9/Ob8U260imNTrCi73dvKPFfJx8F5ePIvWM47XVEZtGFwyVSfP0NwI+
3Co2BQwBHuZIUi9QN67r4nXesMvJ93tqUN5RM92dtHk8XXxUoUUnaEe6bH9hscST
GT+pyRvazmhRCXS2v0fJKrwRPuPhyeXh0lJUJELAGb4ocag7V59e6QxnPScRvicf
WnMmLZQ5xxcqhtdKR5OJli3Cg1KFSXE2xpMrCbUVrZ2cPDlJqKsWZ5KlUOsAy+5W
QdJaRMBeX6uuKFWJnHImFEF/6HN5ochytLOCLyiYF+H1KB0ixmHnLQHGwtQXEd40
TsEX56e2v9wYLbWS8uxNjbiF6w4OaIbP8s7SzvvcSWtrBOZCvWAb6q9RmEjzLWYM
Irr0/DpIL54SbL9RSymHgKHQ9zIgj2wjeB4OjP8B0ib1/ovCXLWxnppCilhvGUR5
A7macoYi4mdeUJfKXDRe7XBkH63hNgM9u/swL8pkhSD5lDfiQQPbIq4SicF3WFZu
tsEZ5WRgOXfNvPTa9cDxXr7IgvQkA2hLcHXQ3GX/6TZ8UUsjred74yoYomDYCeiO
ypWaXQChpdtHIQwKgdhah0gQGpNwvItbrd5nKKCnU9MjzNjarBEKe260pSwR37XB
/GbDb26S9ZkT0Bcm+b+xk/ca5amVjFMqdFQ6Et71tU7BOBKF6wouF5bwbyvF1zrn
5gv0k6+GAgdF1BGkrAz1CzOu1YOlsPRX6BJbZvXFZ/1ATq/EW1ZRKZfyinQPuOPp
FQqC3bbtIijv8+pjJBPhNgFVjxxpStJcXHvZOzM+lssV8bhxALcU6LjW2AqviUce
Y65sba2a5g5nh3L4p3CRlKM/neBOWCcKRXW8smg/lbQ60fT5NafVc38kAMMeZAM9
F55SnzRNzTV70Ab/630yYE5IxQOuNCmcvgTO82TYBUyY1ZXfrlvCgKfyjQS8r9PY
x4rR+5mJoiGs5poFuHI8bZlH0Syv+x+tt6mjm1UAT4oDl8o/Byi9EXeHuAB5lzhU
22r8XoHwOHKgacgGW2X6StMdE15r33qGElMbu+YYjlkZZYo3KpDFTlTjD2fv+CGU
hTNZ/IIG6NCad9ynsKre2gulwaA7hrvxTCXkDqMmAoTi6jeOHbqrx7n/acWAbjiO
zlFL075E+fcY30uDMYhoBv9RyWLkCPPNZLf4yVYc7lvTsGBSkPyg05bKjAJZ6l6o
LmxXimZaXhVRyYS2+ennRj0cGZiirv7tipEqIQSQHUXWt32GmzMkszNwJ2Pu0rMg
1DgGRmAOydCCaRt1PVYQyupi5TKlCFCVjiKMzSlfIdXaq1GWdzSfxyXFqMYXGneE
1IgJ8BpHlsAGjn5KeaeSmnKShoES3a6L+BtQVWPshS0S40WsnCbCm4bAOt5eIHAL
+7m2U/z/MYbOQ+HEtg/llgquXewKERnNp//WZXuw5H1hH5qE3UCZ2tpX2jluomyn
8LwiHkYI71G+qrDumavSRS+LbAqEk9OIeHxw0oSIxCkBjNlgEVDkNdg+1/PSWjU7
47NEcq9dezCol5VLGzvZnbaSzEpA0n/98sQt/uJhPXTFI2ZvnawJtwckMrjOZ6/O
+C6/1h5b5HeCuXvc2Fa3yYxSJiT0/+YZJ3BYMkoB722j8vYmU4ETdw+O/sAYmNpO
m10Ai4LYnRtg8UpGC5Vib66C3oTu1kZlpfartB27xmL5R9OwIMJHjMSwjomCtXCc
GlnL1OuLtHxWhhl1TQZxPsyTyjGwRwTGYVtycIUJOycTL05BKIbnpMGyDzi4HGNx
wPVdyc5dGggizhghtjBpI9fNDiMVnzq4zUmwwgBGp3ZWcex7XYlVgJWUflIgiZ5n
W0xogq3xzdscARbcmo63D12JgFnYDlYFpmGxn+0xMtkvpkpNqGc94Z9ARBORnbPW
VE9lpDzfMjCoDINoqkgIJgP7lNsV55i1luj391NIMQC5QTyTLeLpvYQ5SNQmxsHk
WLWvlOSnSa4x8ZrMUjDXJqxQuD7R85SmBu8jIS65qa3cY7N3MiAgItTw1n83cusk
dDroL8DCv+BclgtSGGRIcNj4OtowWEbLRpyLx+ymvMhV+9Y2SNCy9bac5tY7IXT0
mV+3mGMhBtV1jusZ7Isckdkac3brUpm1/gSqqrk34A3cIxlETRquWDtVK3gz44tF
00ARjXsq0RirEDhxVjHcxONpMasc4zqDj9slXcARxwWoYyAa4m61lX9t097dgPtn
O2Fz+arcfkT95JVGDkfSQgPugTLEZ9OYQfFTzxbBDkv3NgrgbN3CedQdDQxoux22
3QOTwy82C8ile8lzuvbAoYNWpiIR4HthOZxLkTCuSNcHTlxFYjhSoWW4kEGKb1HE
jDLKhHhMddJx9n0spwfeTv1lpi1yv9nWvd0qBb4BATzC4i+HzBYr1Cs0Um1LsuOm
u5DuTT1kz9jNwE5BYfz5RyqeKfQI/Ha2alszW5jm0iH/J6rYC1lM8AoBgFLPs3FW
htxCfeqKTmi8AR1NR+b+SFgb2OHfYz9OEporuMjYPuahFy3piUnYVpHuH86cNc8N
8TR1oNvClGK92fXFVE0kL5Urw9t1htma7jJBAPlrLLjgW5HvsBpudjtDi2327ZwO
PI2yXToCFZjE73ljaUAliwLeHXRWNr2OtAHUs89cAu41kjYPOQagU3JjzN1tHdmE
Ec9I19qIKGKSGUzuluW77pBJeD+V8QRjCHXZpgz1Ui2y4jli5ha7xf12p304YDkT
wtOkbHl/e7YaMxJjq01FGO43ypnFEpe7nxebTs/KgM6MsyyYPP7xSVWqUaHb/SG3
Y7F7n4f2NsQN4xE5KFItUHsYsk9SMzPCe7LUsvLfcc44Hf0XlwQmooue6ldg9t/p
BkF+Y0+uNbqWejR60rvCFQepxoC4RlokSiVNJoBYVYUGo18qEGC29WtdTS7U47Ut
sICFsLyy4HJEfvlY2+2UbYqIJ+4azrhL+axCbE5k0N0gZT/ZFmljoKBkNeGE8o2q
r98S+zSjO8kGEKTCa0vuGqFIJHoM72qQDio8tc/dWKe4NhHaiFx8l7W66gWPRsXm
qfk65GSgz2fYS+fPKJAmu+gebrKL1ttngejjktjZUBwAox9jK4ElOFft5Qglh4ln
mfZyxH++IBCrLIOz9KJ8Xd4NrBjmDJLAZF1qKcK1lgqhXnNkSMyk5JAqKKJRXmWN
M2OcV8QBTJCJlTkDBNAX5881q5yRIp8YV0jDoaP4VZNMLiNHNNLWvqEaIRzpAEvx
FgYCY7olazA0bx/m6InZo24wvEE6l9LMSdrYxtNo6bmVALy2XssejrW9kqM7CAR7
HiMTRfQwx6U9McMCZs2hu2tgRFLmyuUfbYkSHQh/yY5jsxD6mLROYD9D98NdKsKh
wzldxi/JLK+HD4rCl+oRLvWlBY9MFYDgcG4e+pYcJuV47a7HFepYiiMDmdSSNFBN
MNRuaQDw9HbeV8PmeBoYCcNuhFLzWCaFL7nDasG+AWCdW8TQMn42Pct+6h3tgNnx
tvl3Bsrr0fjaspBLqeEnYPIvU5TrDc8lXcozSj7+IE2ikue3nUTceUyoT92R0es8
ef9Z5D51QmYSgqxhFvuN2Nv+Q6LSLL1H+p29MF0SaKhM9qkOKa5kmgZ7nFkBbrpq
JT2RShMcLUoycf5TffD1XFNjZTbKO31ECcsCDaZWbssmKVL9o9SFhUe/aFyALJtO
CRpwmcmkUnzLunhDgO925kiIGuwR3KU5mI5P9htZxEFP+fD+MSeTvgrFHFh1CAQH
HGkEP/QGTjGWMPpiRoDdVqjvN7eSjHa8TYmjieTiMtWjsfnyHbGgui9g5bYKO1TD
ySAhDGi1/15UfU7nkEO5GG+7wbeUNGXrvgsDPiBuzWfqjKqwnI7uA7/RCfyzakpW
qOBSrD1hqzT1CxxbBtxIUxWPgBOAavozlPF9Iv9lcHKvJI52qtgtgsG0wgiLUvuF
B05ctCkYpn0zwgB5SW3Z9X9zi5qtzRRU8XkruwrflZIlfISkbjt7JADs6swd/xMr
1Ds4nPBdgA2FxyAgjvq35jxy8eYE4akYgOL4RRVvr5R8UDITeY6zS6a476yE48TU
Ym7VeM+Bxo4cakOMnDX9kUAgNLZlvhhZdRAOd+v19D0H0sYxJO9igUeVNOlsYnnY
ZV2yIh7hkNtaao+C0wlnmFkcJbsdoDKoZeCIZC4Z94qG3YfaSur+AVrYYl73HpV8
YT5z+4bIR1YeJKssQro6OT9x2lbMHMwUHeNHxDDe9M9z7jbVEziL/rDVQJUamxWU
CMOzqQo8y3+UBHhJQ6NcjV50sSCQD0wCoAee3HptUxkgNQNDX5Iuc4K0vwNUbEbL
Hphs/lCaaFNYQWPOcKrF5rjPNDNZPovm5yhtds4uFRFi0F7MgkFsQDgtpn0vAHaL
hf3oxhEMLG4unFrIJnlybODsgP+jSJr+cG3lr2b2QKp4M/hVC52yRGfG8foIvM3h
mAgL8k1dWCyXoLTiK5HBA+GU0cB4sBn/K4Y7zdbWGErAw71vEn9fn0fBZwrtUfs7
8/y2JehIeqLpWztaKR1XabZmJbX7WOuJrBm9rKyQJA/m5YZgM5m/Y4N4lSp9+WPm
3t3hdJsD+BitYW0LONdlc2iemyff+3aRmzwOdwWQtXW85oQn0TMmWAPI55oFBevN
Pr1EHdrilpRzId1eghXF3ay0aFZOT4kLKI05tmoD3f3ULxGSxWFuRVa7a6+gzKme
frVMd/xl3jIneKBbrskYpL8jZr64EaShnYvTZ174eaTXQX+n9kWAJ1OVdRVWancO
/gGUBOYYSumrc+VXmNoBcDwpOeIbsGDnM2WLywU9aQLPrj5WAmx1JLf5B+klRkgB
SDXTKgnEDV8dG799fKnqRh1SZHX8kcsBFV/EIlNCpUIi60f1Kxsgzl1VLfC7pNLW
tm2VBtlPt2RjFZmtaphZhxihPcZW1InCec1AEUQPlv6L84pByD+lagoAHBeKym6j
W/g2NNSvf14wR/Q8POzrka72EzRoWpsrOxP0OD8YC8Yvg9YxgyTDDSWoUUQlzFr+
q7vu9uZD/XLY5X3xQxaI3/aq4y7TGzKoJUkJ/aC7oyEOCS+SxS58DjngjjWcK0uf
/AEqt/6dkkmt0etUYCrCJ+DFm71/ArZ0c7YV44XO+R9ErU21sbhB0k/cW1KL6fNd
x8EXsBIDEjWO6E4SxijJvkuedid/j6RgwSksxxkny3x/klSiA4lSgf+7ykEf33ov
xk07ypWUZ8cvgLNxMQfTFZut165Xv1YhSdvG153uNrhLq1Faf70tBJbMN3il24xe
2gB/IlS7HRvEgWr6laGszUOCXoxfThTvdbLhLGYo0uDrzS0M8V/rDaadxErQUZ1c
d+A7IorHllAxpeRsFSdoxHWh0D8QrbaOzPXZNSbkuCU9rnLMFUiDXjoJmng3SYkI
To9CobP4TRu5oXA4LT59lKldPThLz7VCeWSO8bl0pxvlXo58UvaNJjxQL9RGWhbw
g4E6q3Iv4V8bCaaghx/5yNl5LvFAHwC6Lh2K9BTGEot0NzD/PWtEfpXMzrcKTjlb
w5YQA6/PHbMRi7iv7h5EkDksChkvH6Yr1pSCMFtOdhcik4/RTpsoC28Ss/ydmxcy
+6pQ0VR2C/eOj6BkBE4Hga/g7cAWNCh2K+0hDgrK4SH9TowD2KlOy440RtoZiHOD
uRxc890uuF2hWXzp+S2S6uFmJUCZd/FXjKXbSh2tIqRX8kmCDv7J7zn7qIDI3s5v
9ZkqM0NdtO4NzmiJ0yTv+1mi8eUb68QEnKbzvrudujAUu6JGs0TET7bht7qqwEnO
jUn2S6QcLYq8mFnbhUSJXOjsbbJKOhkFH7qXPFrSmdITyBpEYK2FGOxhpjAKSuIr
HIKzzbHi7pLv4L2/DWCR2xediRLom/lNajYAFD048P8paon12h+hGGaYQgSRfnBx
ZkZagedEJtx0SUsML/hPJOH3UaZ0knqelhEMRXBVE9YvHifnz1wF8+ghj2Q288V8
oSPfp08ndjND5MDxrj5m52NKRTZ5i00H6n6EJOjK0DhXTniQHrh+rahROuxoqQUG
gikhkdCmnLvFNWQpt7UGsocP94qpzMLMYd2ty9sE2Wwn3AAZivl9m5wcqjMeQmNl
ECMRqJvrK0RwCbB3vtl8sp/BvKmN87EcvI3VC9rIzG0bsmlsR5AujxhsxC88Dq5d
XzL3fxg3RVb9gLNSFmDPmzpbvciK8sJn9p8KSA916EU0+QQSF6U6vAhhrqPdzQI/
tttTk61YH0/mwBIA+txm+l3MZHTZNlrdpAsRadoLxs8XRFU9yJmrM+lM/s0eAR8w
VgVusz3PfDWJgOo+10edJ4ERMl2gno/MxpBlDyBXxG3qw1+s7YOjcNiOhUOpMeUx
dCKj0YZUZoF791/QsOP6oA+sz2vvJhTU5WqRqVQmohmglfsvb818pNdwrVTpsFfK
cmjzr1ExyVaC+oTKC+durdkzWvrqBg95DqReSdJmVd4wGk6dOHztVISLxBe+fsgf
uLCHbCFrht0OJo4pFVjFhw5bFdiN9yM4t7WW7HQsnlGoSrMEi4EBcbD175LwBy4q
qOMcAXxbNmB6Ul9wGbp8adRksnWYOyKtk72jgyNy3eR3+HEYD5+mLGWyPa+qdkBA
sBsr3yLWTG28T+T9QiOng5ZQlLYz3epsDe9NS/y0XB/DFvMXbyBP3D0vDvdxdDL2
c2gtm3auL2ScFul7xmvNro3pGjouQQ2srk2QSqSVJInwKtO40QqQ5BI+sMXJT/w2
/sjG3/ppKvY5uIb2vnA72stjb2O72JOcOSPxcMdnFgM1QSVhEe2ZNjQmP6saN/0B
2Ziy9ZuZxY+P9eF2aoAUg9SACBNK90ALFqHy8Qtr7639R2psUPO+IjGnSmp1DLYc
3REdLBRJTctfoPquuXrYeMu91MixE95z+bzJcaZ0CqowsBQ7tjxqpe5ktuAv4+6P
ZQXCUrJ3Bu9163VOT0gOjYrOsTlzYCTByDCEsOkP4eFZKdvLZlMR1s7+UpvdAvs5
XPlxRtI/t57pVolehKY+9c2Crw1otorbvAjvcsznLMHmBlZfTmTpUcMwHLeJ8zaY
y299TNnjEIvYiRz7/XwYIv2Zs6ys+A58fLvz36kS/WB+/97KpSFu+27xDIwutp5o
TwF7axspcEIZWO1YvipY+PK2b4dzN5hpRXTSawQrdoe7vWDaBt+iDU0kvHIN3CPk
VpSRkqyAElAq1jCg6hfiZbCMJAzGOGUu/eAxo9cay7WGTa+nhmocOtR33aIiwwMQ
z3H86VGKSj6+zywHBJ5pCCZpCt5w9ovn0laHrAL1tk0SnI0B/ObeVKM7NvErxXxu
3F2PDxWrePC1Gdy7bLl7rqzyenHOL4o9kDOb5/W7CtrxiBastXPIxxeMRDtj3ZFh
1Okbf9p+ALbDmppt2kVf7URcUh3wgxkKLD6afYiRmznobnTZb6kHXElBA58Z+1HT
De/Ka6KWnWL0gSOSV1xDuppd2UWPgykln1SOefxMO/KHbqe6tH+JueJOvx3uE+y+
hTBeeblx/55Sgx65obsQgeAmxVbmcmm7nK4lWw+ynNGKw4A3v09JLmfAkrA3c3he
mMKUGg6RAZGPUq0fFiDsfLMJO1J8YvZ1Aw4OtepWSdNEfrnmd7qzlTZ3UjJEtOtL
7gnlOE9fnV/VnODpDbe3tQZrJENC0Ee6gkJo72eZF4kR4WT8sax4GbDxETIit//b
U7BbeahlpCFkwVdQJAC2W469ER9sIgywnWpLsjnb7bcscDeXKnxbnCYzrHP/jsnb
yakg6B+JDbptUi9YGsG4RzNQb0mtZ3GmDgi4U55xNYJrRvDA7IGXoj2k+3gqm9kH
i5v8lHh6pm5jt+L+viQQSmw5jlS/Igp26z0IR74tN1MASIi400SyFfcONlX6qXQ+
2/JTT4Ph2eeng5CSyFtxwwHepRB2jMKtlZtgPapzOiMaBu7JshlQk5Nrzz2MT9Dn
OwbyMDeGf14H07qNjDTW0xM0rXrmEt86YX2q2ysWf2/pY7lNXh8wg3ngIV1BWGd9
BrqGIFuW7NfSUtRQiH8w+fWFTN0dCALUFgTj86UDmdUIadBAW+Z5Ik1wRZ7Et5dy
YZsIjajv7Gg+3bBxdNhPO7/ZWa8rcTmcHH/kYkDMmP3e7EgjDpDCt+VjhQfT1Azt
4brL6SCfRL3FpSPcQl6I/bw7yhhMnUBNrh6dycNaz2SBZW7F1/Xxq1iwlGbpQfHQ
Z/pg93uigc1p16j8GzV7wULf9bbo4/fo9TDUIRFudmq0Bkx3GVXzkc0P3Yr8oKyo
/wxPH02mI6IOB8vO0aL9M8F6eT97MKD4UlMoeSGVE1XCME+IezNMOc11WDubNrro
YArZzb09dBkZxElS6mFWix+ILuumP+4z1X9qKgudzVRJjq23MLhy1WT1tWBki7wG
Q4GvJhGD4OL1+GeXcDlHGcmkODisDufvhWGC8jP2Gmj1HQeB815DcqzYBxcpbOPM
a9bnvbH7/bYTI8MJjkBpd2T9KmZb+UwPqG5oFhzCVPOjbauAit8453vnxsdlywUs
lkqcpYOUmuifxcQ7bbv/P5jFcdpV688NMnB3AUlay8n5Ij5xJ/Oz+wvzbwFXyOcJ
KMnTKXrVfiLkciYFIr8apt+9M9qvlUY3FiAddyRi0lkCOqi4WQUoj6/0OMNeQjdv
aP3L5+Iokurfu2NzwQ6gMFSQopOWgXIB+vwXzBCfqNFpxj8GyrZhoDs7SeGApwtV
ZCb475VWMOBiOPgEkdn+kKIWHfyXcTx9hlifskwUQSJBoghpEvAkif2qgehjdye4
uezIewnh/tmOjGe9gkGdAniLMvdh7gEqAM/7X8edm/iKEx8Fpn+eFHLD73QNOhNp
cenYRBPXdb8zTTTuSXT5dO8taMykihBQmAGks4YB8aOQaSBJJheF4hzN9w2axofo
w2JqbSHHRJ2M+VlRa0b4QtB0YdFXyRBdkIDQoH9pKKc5yKCBUDHJ87xu4Acr9jVA
TULyY4syQmRn2LeEM3dRUNMBGcW7zDAO3jyEQgw4fYCa5j8BTJb2F8WXY838i3o9
0WGSLX6WyaC1oLpvTmW3k4PJwWHggtxcYAgsAwsKeGJ8Bw+A1hcJ7ey1v8Z1xKoA
hkwwU81xIPSAv4Gdz0dB1ICQksqQeqUw5s7ZU77a3dRkhtS+dhrQn5wgDyxzXaJr
P1ZG6Yax7YrV8Ajqd+Eq3sPAV2TKjmuO9R6/QYNpNAUj5qHJvskkR/wXA6JlHNT1
dU6BjRKXraTEsYkz4BfCauuB+F8iPIHCeKyhTgOx42BZimew3ohSDN/9817heVgM
PSlNMcNNWKN4arm+jg91bK24/FmeZWlOq23uyEuIeEgGVoCGn7hq3ORnIxXkksHJ
kJBbN6XAYh13OS2rZPzoDSAlKsbaN1kRWmFyKRa/nGQoXqG9yDNxPp6mKemo1gAu
cnuJ4iyCXvT1a574bqLeVvaBTrDeDoMAfXJFenD2MHZPTIVws62h25EP7iFvQAlq
rhO5Ug95aUsHkqtrVjCr5jtr1oYXNuW6KyQgOfwA/48OQBy3wXNfZr/l2sd70gsm
+ii7eTUyCZcJjl5G5ewlC3TgNDbVw8k+ySzbky4Zju2GHjyFp0dW33imNWbLQD/w
IK9X/6D6T3ghS7TDLgOZzvbXm57GO130bnoTiqvD2uUWo+Xe6pK+3OvDLgvBiGEe
wP8JNv4xUQWhkOXwq0Oa4aLofq3O4hrIGHrKnW0a339icJonCjAzmY+5mIPn50rR
JurZJQzXvzWwBYloZE1ldgqakv4dTWb3V/M8X5ccseIboT9OPSdNVu8w6gyNZTLf
7jFFKM9OCRZI20/IMcEaV1UwAGiXYyv6V6+ffFFnEY+y7gt8/D6m8TzSanthu06p
msXFx9yr6JSigo7AIod2kep6kDUIxjKJSnrvcji20fSnXBRggoqabLG8y54unXQb
5Tn8f27HX23FG3XuQHCZw7wMA1LDlXylNtQvbMgKRCXuMNqPBUQJ9MoqmNo4LSGP
BRS2nnXbMRxZ5ukJL2XmqIze4R01NTCS82Icpm8utXamJ1OS/z5Gltp3bp9g1qc2
/6smghShrCHDZIFO+hAGzAmmQ2OUKnNnTstrWeg05rldauQLHF0LAd/pSXQlhK6D
Urm3y0LLLVo1JKDEC9jc1NI9MaMQwisfG783RiOE/Ok7Dkmwqv9g6HK30els0FVR
SlAE33/g2lEhAa6WVauzTJYjvUyVmC+UaTdiNTr/JM6GowJ5sk9IT3gvNyovhLHe
1lhWKC2+ijkPfZQQKNHKng9J5PqsNfjONXVvmiUHf42J3I5YcdVb+FwD/QFibpYY
skWi5AUDVuNm+nAnsDd+sQZiB47OK3plfAWsyxIZa8GYbjhvSzbOS1KrHKcpmd/0
aYENNFGSHDPxEE2+gjiYc/qhBom0EuUC9sNXwV0gG70s7ntaoUfkukEHtBjH4CUc
YRN/WUNn3rE2IhKyfQ6OsFqDoY0TeE6hoT6C9reUBbpURhgmFljI5lANzXK7b4MG
NK89+wcYOzBQ6XxRomyYYqjjo7TyQR2P4L0JfJ2iVuuzTsF1s9stzs1HPqnMOs7t
H3uUZprbGbC+IYN3U5ehf286T9gLAoFIY/Q/xPUELPAhQ61ygV0EJAPVAd9tYgJT
nL3/XLhovWGT1XPB0CmworsyjAiy/DtNgUtE04BjeX33V2p6l7y7k2tjWytJP22O
T+sEqK9N4pzAwW3pLaOSE0OYXEm5/O2MK6QDkBFu+wNN6CUf7i5nCBoH5QGFoH8a
3q7Hu5u3rL1Vi8HtlVVWhqkeY88bprqDbltQjQleBBJ6gZOXGCDs865RPk5LbyrP
zBoojHMKRwNVKYIda4ASNvE0NamXIzD7ZxN3ZSFsYRS7hg+eBhLx7yWqyffApqA4
1M9EufpfSgFrHAKuvQjk9noXPdD3eyRYlD4EUPSmXljuoIMrz/g8Ftq7stj3rp8W
9MeHaoFj6FQNXFJZRTtCxia3xj/tR350uXaxZV8fkIfVC2XiYQcrkmnL1DuYNUmd
ycK4QBqJxAxxXXFNXo6giKiLEYC+nLsTIjkdJ0a5+MzqoLZcOmpSUreinr9vJvAT
5M2pYCUzEq3Ue/c7zQMVpYNF3O+0Hrd8F6ETfMqC95WNDdzkBh683KfHYd36bkxB
6v35qL1wewZHmJhuxESsRzQ5Fiq3gN3OoRgvevy9RypGbclIhU36ZLpgWCQbEueZ
8A6FkooX6buklJqjhskjeli+lKWmzdmG1k2VUf6gvM1jq0I2MgOv2saNa5GeBB2v
r2ScbQVPytItNWUI2Y5tBXjvIjIboyhuXShGnMrHpnU0dkiYc7NE48efIOkRYioa
uh/taIUdN3Vfg3JwgDU2QQe9JW3WdKJF2fJ3B5b3xjyUs/Au8OliFRLk9lzS4YZz
v5WEl/QjfwY/ES0Bm+xSS5Q1qqnBlrIxUnfi2BKaB+A/hXoSXhlKgXRM5awgloyn
3tht2DI3hE1Sw5QsFfWLSPojsXel4p6t1e9miDMviCYcnmBHjpc7CHJv+PJJTw1M
OhRlAIScqlEMP7ip8DwzfldH33ZQ6VHc4p8k5JAIplHQXsgtjFZddETkT70Ep2El
2xJGdltfvxGSNjqTmOY134J4to3Goviv7FIat4jGWFezD4kyQMAI6k+riDOfmNX2
wVd9GVX+WOMjVr4ogaMW93BY4dNNWEN2I/BlwhgmIgLpHdDXXNeaQesiXAPZL+7F
suw33w7VAQp/ClZg/NzH20naqaIjuRaLDa2KWNn15w7FwCy9UZ4vtX+WR2h86XQJ
IFTnIWEXeOs0lv3kV4qPS2zROTxHbRUJW0dFlANITR2xHquxlg6GAXWoQujSL8GJ
9UWChP8sQBZFDsvvImHPxcPnxKqOrO9RsIpHA5NAtVXT6MfMB7n0EgrIOQFiFGz2
E7xmF18VX2SdihYbLmXiONdfVDtNQOKT8Ka2dEEfw17UpKcCtgb/YBRSGQATLUlk
KCx5Bqx9DxY4lxKTM6vS6N0TJbMGhebEA2C0Hb3vJwifVv9wBFXBS1n4dNvdhML5
+0u/sTZ/DchcQeF9G6X55Wws6BjohhNxj0qJ+eafpBXxZBHKS9sZ89Ng3TFYSVrK
5BuLvBDFdYS/L4dnbRebimdLkX6KXISetDGEgs6ZC2NpVtXcBYxf3nLVbPBuzTh3
OEGhhpLvNi7SccYcN9CbWWW7L7x5GSVO/b3fUJZlwuY2NW1g9v+c5RVWhnnHhNGM
+7RgdI9cQVaXVWrOgiB9XA1jAmu9C8xy2jjV5CUX1J0wXlgdfD9eTggIF3yYRH3+
QznRkK9ROSFdauPDuGLaflmHAT6TormXsGqbdsKGnDzzuWfA2cGWFauFfdF8sEMV
9GEGaXF5giZHIIkxBvN1HZ2oox3aIlf+meBOAugXnoYPYtb70IOBtWNVzZgA4pFP
n6pEYGlxUCKO+Mpz3bUervw8O9WmB+M6UssGkXM7pVlWencjVHFnQtxkDH1zzO3f
92nLeamAAcdUhB9/yWRXDO8Beu6sE849XqBVd82V5X25NB7k9D6s44N0T0Y22nM3
fpLe4Snftg6TENuY8ZwP3vy1oIkywdiMK8C9XwnB6iB1bYD2vkP2b+8v9JfClgqy
dK/YcA1rF6Otjzpj5NHdPGRjxCoGRfSm/WwckqxNfW7l+mzTlwM7lOPrVAzlk+GA
z+MrxEyhvdfBz40b9eI/WTbrbFC2CY3eDQFVOJcYIY6AMY2/f//maTNebUDczF5/
F7ac+WSdO3sxd8o9UzB/aDp0NMewwW1KvjVlpdfEuRrahYn7Tg0NZT62RmoYR4yw
TM6QFqacXIWW9RAw/ncJiJimVPMVuwIlweDtAXxWr4NOOLnT7jXBiW2bsb+no82s
FsiA7G52zOAZ61uccvt313UXhrxm0ysv8Bymyl2cVwHYfQVNy4oC7sABo8lh7cHM
UHmt8qZIhoBC9vX5g5xwRR577aFz6ymXpgEkphxxiylqiZOBVjHOZorMVxEnL6i5
gJ5vvZeUPZApp06D0vq34PcCELQ1lGIn3slehWH2WpWuwFAXrbj+9+Jla5DLXcVY
Kogqzre4X2xE4nhcIDsE9qIJFHF416cFah/GFUaHYOYomtbevx1YErNaL+SrB4aY
q3GscFFN+emupfU63ydIsufCpZYKg0sP7jZWEiRZDind3j8QtckLYBzzUk47ABpL
jTwRpL3ycZNFStprNcFC0U67i7uvYnH3sxl6UpE8xZlhPfDgautuSISTRV1xGqqr
5tYY0iCCpeUr10JQEU3U1peMROKyLqWnCFrZZu3/5wf44YJJEABCe3F18BYp3Gvz
LgR4DmmM2QVrRsehtxLtcJ3uf5lfRpvZ+P4RxYRogoeR/Oi9A+jBYKqhEanUb5fb
RAeOFcQCnAmJRMJNtMpQUQswSJEOMrz6BPOeDT79z/VrXCCIJIkBxblzCSzLWWK7
Avwk9uh5JVrPfVTarTGp26EA5UCrkaO8RwXqHgfgigqMBRbIEGk1npNjOVM0yD1D
yB1eN60Ow05BAIIyyubgUsbbfVxWTBMLQsFJtK99TWnfk2mMJOtWVEp4oBo+0vCJ
f8B6phPZfKLI1C1JrdIcoq5kcoKIpMR4tbAeEXfcfc3QggzKRezrZHr4oSR441Hq
kT6aU1BKs5BMGDpsryjiLLbXrWf1uocxfpZyQMIy4KzqKgCXyZY2KLnCpnBlFjO2
00ibzoL0W83aX0myPb318gBM9SLfrvZ/l3NaK5TsYR2qcfB2PHj54hMwauhnw6rf
Ni3W3t2ZS+RsMj1fcTXDeQXYnOovoD6x+pSNL1F1i92PMZNNOhUh7HtuxnFvOyFh
OxYvriA8xL3lxvz682EgReWc0XAMP2ZrYmtG3MNC+14hspBty1tukceJUPHI3q2p
0rxU/BiaMaUJg7X4WrinVFreUHEplWaWb7mGDV+WneZYbgbf9IqJHSSurUe2ZqP1
6xlovKlDf4lkOBe5hdvbK3IOliOLld3M7BdEuZsozH7bkNZeGQ2eWvT6YIZDG8Pq
QDM9QKMqPONIcl7VfNrxrb7fIlHR4cL5pGdy7UfNQJmFJrx2W8OwqDgr4JMPmqLc
Q2xnNli08wZTXDUdhmYpsP+7p1d5+shomqnMYOUeK0La8UU7zeNe9WfeRAwth59q
pj8ZFXj2BdhCQWwMn2Cr/S8z5KnIvdzjaZR7t+s4KXXnF9rIjZkPSTQGG7fnGYLq
DeJw1JwzwCkjdFCEWEjZzwbHcMCF+0otJuIjxyAWO55TiCalCZ2iyBRZ0dltRrkd
esaLeIb+2h+qu77mZePHu9GT5bEBArso8nTHYIZjQ8WYRZJBhdRz1RNxPd1j528L
Zl6X3L5DQA1Ejaye+2EdieW/sQzSQBvVeembEHwKJQhNUq9l2ubJt1Kl1FNhvZny
heUgxSjJEvfBuVUuq/DEepYTaOg+AojZzmqxGhH/AGnBxgBNwXZXJDahDdqxtRdW
mFbG40FRxRd557lGsdO2JgKE+9/Vbvj9xExwF8CS+jHV57BxY8DSnZPAlPHKyouX
MPjBfNm4+b6wqwrusv7ptCL6JK+3vVR255ZEghZ9VrKaAMb6DvWyboz+LkGiPBk6
odykiB/m9Abo0EcdtCqd0LkVCdC2SPM3c+0R4UPQiBIc5h+9nCqHPIIMhpKWNohp
i1/D8qDOtHeYh7hfoG4VdwhgDxUibUR8/r4uBVGd9Icx76DIjZhJ3AgwWVpI9Uja
whaR2a6cajsueVfkFmFyOKlvbfyPTg9ea65aPzpLletfYVQmo62tLuhE5jr2P+Hl
yi8M7FcoFIHK6AqhjE7n1ozEtNOlNmSUAh+1KadDq1yAm94/UQCekxtav4pAoumH
GaOvxPp0bVDPfwa7eKynf/t5AT6oBZndDOQL4b5AiqzuOXkeClFCRUE+CixGPauD
l8wtnyxb0H0hAhPJVHFVJeOQ6vfIS98hJ91ovYsbuKj4RbmB67dyDu7AAopRTXvq
9XauFIFN3mX66Kf6qAknrbK+wf33PDzymYU/xzMJlthgQfB7WRAezEIiw7G4SQZs
7PTM0odRqVui05vYIIOmEB83kWlXVKgdNIdiLnchVsU5wyR1Uh3/iC9AvzEOhTMI
HEIEWTH1yr/2dk/pk/tcC5D6uRBqZncVpge+YPyID1J+TPVg394P+IUM6ZC1OCXZ
EakUdF/VYLl9JmFYLoRcO9XfxfD/h+KwM52DyATTGDN5cRUJejnKWcl88fFNh6uz
+dSWIsI3EExnsXIb/VHfLmzIdBkmt9i5sflyH248hXmNrfBDy7O7hF9r+kuU4clS
wxFCnv0LuV+TTk0BelXAzPZ9Kc/LcHossj4akVQwk9VYD7lSbwGJuH/ik08brgOA
zEXnqPhsbp6/pPqpNWmfiEN4D5fN4n/Mndtvi/ZCOrCqGHT+UORxD3YBNoxkgGij
EuL/d3ZIfQUBnZuTDq4cmQhqeDikN7k+2Yg3pWonxdPWuM559TCdaFzIGEOh6Yv8
QdIvSnAm9bNyHtfARpGSGx9YbgdKQwAJuIUS/lJhp5Kwd5jc6w6tUDHisoF5MunS
RsZgPHTZhVIYNTZ96uzgEknrZ1HOTmlRy+eGvxEV8OGxxRDoFRnObl7bRCgwRQia
S6s454a9yzBFdeGn1DyPypOUOVQidc1qAtiF+lO30VNXmzi1Kpg8fbKhQsu2yqU/
Uf1AtAwozER51YB+whg9ZeoDWOANQK2lUcIz3cgATOg2lDjSz4ul4fInPLFognWb
Wrj+PThFTYDHsvXD9ByGTrdKpttvPesP9yE1GR2VcF6UsDAGENRlyrLAe7sJz1mG
Ta0J5EG9PqP6XrvypGsB+Q4XRTK/4szVs7ZedE92EpA39C0Z8x0fJvTB9YTD+Rx5
+4ImuvBFDXTaxX5si2dgiP5l3T3Hud3d83b4uV4FtnkXDG6S8a8Iip3scgz6M30W
CDx9zAOQs8Ca3MW+ojfiYI5s7EpsvsBKSWTJneTYAqYREOEVWSN99j+gEnKMUPE/
p42o+gQCjloVYBuP59n0rLI0GRaxmm9tQtBBpA8x73M=
`protect END_PROTECTED
