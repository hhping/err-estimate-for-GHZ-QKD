`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
53wWnXSl47AS6FwhGv+/b7naoLVXQHftxcDkvv7M9rkaKkWNG28zrWPJ3IMTdmE1
rjK3reMdCosFbRZJMOHVjJav1PsublPYzKo2pJbIF11Knis67rV3MElvC318GoRy
VfDVwNT84bHtZzNJC70gz+Gpd9roHXZ7nXqKWWPweWHki5nIR9XcgJmSL/P3eRCH
fP847iG2fgpMA5UKd3xYmXuFd95LnvXLhI8wCNwgT6n46S7RvdnyCO3xV98gMoL+
p5k2Upl2rtE5U2yVncTGbMFMWJ7ZbyV+K4qZtD9PBToBSpm7gQZU9xPx3ixcEoBO
RafvlGNCUGD00RpvHQhGoDqd5u2CiaT0JLBwbP8taUg0796ZrjaWFoRU9JlnPJ5e
XNNyHLwoVu5aOJdP5K4icOi2rlU43OCOQ05FUp5iBSCAnEF9u3Z7rN0OPXd2mumd
fWvujILA8Lx6OFUqhmf9gnSTFVcCM4XoPBXkJM30TNu6/bsI/hLb+TTboYUarr0y
JU5EcCV1ijMBA68PV0efhMNgVonvBw6QVfLODHgByy6llRoaBM6K9aLQTnDLOwRM
QhqpjiQ1XQY/7H5GGW2w6UDy/1X9ITiApzKzkWPlyiyrvcJy3hIH0Hh3kA35P25u
LXaBhxsJAzUEA2z7TUeUECffNe83X92fBkpjB7zajpcdCnBu/j3cEvYNVF9alr3y
dL8ssEvr6sCJJxU+sJSKU46K59xYVspPI/VT/cjjtmdTO+bZmKgK6eQAgKvhOeOb
diK9DBEg/npAnlUXDwwY0t3LvPhaP33COQQj2YOS4ozlbvLRuyzOZf2WxqyH3MxS
oSYskGLKlg+Q8KQHkCk6gH8b8Mr68UOZzcqTX+kr0qA=
`protect END_PROTECTED
