`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMWhka9ummA7PAjAIxOXUMPVo/h/CTui/dbq5VfVvpNG0zI+Bp+uQF//Dg45BPkA
qQuiJ0QBazEsBcVgJbvffJ5/L72cD5DRz/OEFjPlqkdeU91CUxICalactRQxR2WQ
UuAw3ETyP9CnDykAEnjOV6J1GfU5aoK/A9w+HsUHqve+NcscZipyBJZAmyB+O4J2
afv6qSvyQ3W0kTym80D2CPrLv4pFM+kqIPv49/nf5BowHE7DILeh2d9EBhhLTU/W
ojK2LEf5Zw/wRFDqBb+HH+7gJ+a+N3u4mHAPGtVCczAkjCRWragbxhc2UZqUK7Ny
i5hfXQkH8/7mJzugAdJ/593jD55xmZE3p69zjRZxHHXSvpM5jNUf26/tRw+FmCQx
4rLzwzlxmRApXDTWAGS0tg0uUvs1xJlKBCz2yBFUJmbnpu2hFzuw/oUdOsRqwE8y
4hGulLanpiVpNNhC0AGkgdeWwFB+zhUFxcDx1ZBVq0oE/h387hJ9Fr4VPCOiaP5u
BmUCjrz+b3m6CVghvmZ5+fRUv6qRM1OVI2whhsTVRyp1T4Z/zHzgnuTjDISZDEN3
NAXuTa0bsjyhknR0MjsQ5n/6yGKPIPl02yDMBxAEpmvFwFCpNsJvo5Firzn5Tv0Y
aCeCWVIXYe6+jeJPanUQ2xImyXE2aNy8oNbgVVnL6sAEjjDcCiHUyseNtvCfiMxr
hiRkAwHdQ6TN5P96um57y44HlXJ3exIpJibtiqdhqVWqTnA72M9LAvZEFovEpqZb
N4nYOoBv2HIcykvv9g4ud1/NtqM0iBH+XqGqVCgZo5JRxjq6MCymgRkJGlhuaoxS
DF0RXhF1OsmALWQZbTzZ9klxhbyR2NgKbj8sscuZ1c8MtmZFIWmk+o1OCWt8mXDr
M0i/S5ACkv+HWvSzwI61PT0zOiCWc7vclTzE/FvpyTLd7gy5MABVS44oEJiW0TIP
f4pxRXCtYtQFBC5ZJFeiR9MSojdyNDE2tlcHmlzyiXRS7v9nN86XFfY/BuKaqroH
BZpAPnEbHktUz8wVA4ME5JbnLgT4Knc3wt8PiuP3t/l9FZacFb+FI+26ceMxd1eD
PsvN7aAtxzQuvYL3LqPpHkNKyWAb0Wy8+4nEYD19moKnbAzYgZa/1zXlLCM72Imp
Ff2HlI/W2mZ1dOq6vxYcTQdrFjUuflxvvQzcNIu7GAzovKvISSy7xwo1tBwxostp
bse+SF2lJuVSO7w+SQLWHVYwMbTDE2oDUgwDfYJI4WZ7rpzFBnwp48Brk4jOS0c2
Fstm38BKuYSM0BtnTbgdLpHYjFHTYRc47GsQiverNA0eG6JIMX+lAEB42WqQrURX
IPfTbLfT1VjsKRTJRVvfrAw6/Uv42yvs7zWGjTIAFBlWYGwkZUeKVz0T4QBtpmez
n9NpE4hHLtXiv0ct5SgrcCeawNANQM/yQB7qcgu+6kMB18WpEElC1xwVEWxEk4dt
EzkSQb+DdnObtOl9Mpr3w84smaYHnofP1p0TwOFJSKMGpkeAqied3tGMmsXTpfFp
BpzAatQ1KX/Z0xCRYsuU0583yzbl1c3316CQPfPUCXEaW0PiEYOhjCrcFDyw2fwm
jW+AKU+EKEDoH06mRP2oWzpJs92uzvBYXGTXu9/WoHpToMIiyc/kOo4hcqCXLh3s
WPP32CAYEolXorkXk2ywNDL5kE0MPgpdiQZcueGuA7ToCRxd2xmauhWxPBCrcPm+
Valupasch3PTwdWRKpr+ZuqnpaokOfBvSDJF4FmxW+8LqlqutwEvOkHfzQpvpd+G
emcGHnEfAW5cJpDZOvYn+QVjt9/aE3WDPu1OQNgnSV4PIm+V86gvlokMxT3apHr6
hjZmZ+4Kh4PddNacRoCQxDmhDKmqz46E01soJmNpaTvfRK/f+Nn8NEXHYwOktKaV
J8W8k2bmXThKO8ETstnaLGuMklyaEcXw2dqa7qjgu7HKPOpeaj8vbZU8LfoqneDs
p5yf3vVpiS3DUcNWzxS2kDWifYm0On1dPXbXH4gVeIpoQDDMxdLTNdT7P0YCZH3B
42VQntg7/S2KBUwmjaOqpaNLk9omBQM33rvsPRTx+nF4eJsd4t/9msBWbEDAjNmZ
+oznh2yielJLBZZinjNXR+mPP2JnNIRcPPuY9KSkdlZnYZCn3KyEGbCa2G0fYaW8
zsMDsmQd23JsqGfLgJCoOB7SdCtovutKBNuUvtyKDXV34jXOQ354V42akY3yhOyH
u5KUA5fmOzRfLqdz04LLmYL/TreTXTeIwVYVPRyoprdbzBOvpF26NIVnooSj43gL
lSCuz+vkOMxlTHxU/Ad3Sq2HnN8Z967M0j1BmvqkHfWv9PV4UjjVRIdUlB4XxHG8
62Jf5QysQChwmyUE4IhTTsWPaefAduTnsU7TOl1bbwqfPPf3M89jPNsjaVfJGWsb
JBjuxnyJJYx7c4Z1YPg2Fp2K9oFDIbOb2Jrj0gzDPqmQCDfBnBxuGiY4gPq4jQiZ
O76VYBX3/g8C/lLFNwZFwniPkLZYzYDcuWL/KYEALw84B5Y7OxyOsSwFuEeAd9FK
wSpMdiiA7LLiYMbeDpW41BJxaucwO6DcUOkijJrxq5XEnEWOx5gLpZBh3fspcVEU
mEdCCqysal1fiF5el3FGAnsjlrFRhuJz7KsXLNjnbmrHJE7nsbJsqcjrCdtkstUR
NHaM9PUCXYV5FF5kT/Anj+fCkmWQK6ajJi++gJ1SeEKxNrDW2nafNJGkRmJRsGG8
`protect END_PROTECTED
