`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnAfJOgARx99sziXk/H6wnUWK7rSjtSllFV+W2gCLUvldLdZLSsIfTWoDdIFmR6C
H8xnaumgvpTTnHqV/QE3DlW3/N0XXJ+TXYuXD9WIZLFlCBgjyZSlBQzcL+ZU//Fr
kMNI+r8Ml2Hu+JH46GTd1F7uGF6vKTeuwGZmbJhXnSnm51JYDLf2DEA0XZeMBaZ2
inuzJnI0IZZL6Nli/+mjnwToePRWg77eJTAvm82u2/fjEm+UA1IEOdFMDFnCNbW5
1PcGIvd1dW1zCnhjMU9a2bzWUn/26ENcjhmUbcW/fvkLoc6PsTulujDySwPfOZEx
ID2ARa/bBYe8jJTBF+BEN5I5nsJKK8/kFfAFFTrg2obkNrMl318Ga78rugjW0TW6
f4fWwxoCJSHItnkAsbhfJZ66lickdshHjbsOxV5/I45OCZCU3PA2g3mbgLkprPs8
vf2O/K0lS3fsxbLruKePa2R47QJut4DfYTbhsytPnUV14zKyrgayrnbOTB9bfX7x
OkBtmJAYI2+N0rm4vIcFW2sdVEq6+qVw8wjahdPBbKCXN2x7KXRQITXcVw+hZNco
+GqYZzSQkbFOazHb8SnqaH/YgVnNDnHWiai5E+1WUtVBNLTbWUGgxkxGeFgqCT7/
uEE1oTB3J+EhSQREh/1Cql3JiQhOSxzAFR5hEPONQkcthqg/Z5vrWbyaUr5QbRWq
kvnQ+pi9WjcOadUZyY9dTO0psQ9fWnLkB4BvJ7fmn7AWlJkjl17vp84kskaCR/1c
JeMMP3Labhab5D9Z/54LsYOw2MmdkKIZDkhCJR5D5D3IQmgnGu0ToJdL33skTBYo
cw/K77WMz/jbszvxz43RHQ==
`protect END_PROTECTED
