`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLG+IgQx52dOeOdnST6qEOkcTvMJhtnrJxmNPF0ZVNwOOj+WXdpd+9DftUtGHYlS
Sdoftp9d0iRskzaaP9986igyBxhkxhFzSqZV1YZBYe9AU3V41nw8naQrfTUJOqXU
7tYGsvsGYW0v3hQlnYZPFg1nhsg4L/saM2QFknWLIKS+NIdOI8oqZQRXJHoIlZDi
9+XAhkGgIzYWwlOsFGO1bCChSOmMROIbaZdmZ9MH3/h11knTAA/12WFhkG+zgabH
R9mhFXOQw24yfhp+7Bc+F+1jjXfebNl39dNbIfdbmjDrm15fO6XwL89uFyhpcJf5
HONqw9uCwK3IKNNnXeaZ0ln7ez9yNK7xS5chbCf0TChr+gU1fbGxjggASd3XP/fX
DyqnSZl0qweOePx4AT98fk0O2q07BI2GcHRra6HKQ6UthaBwl2qWlDxhENfirM3/
30O9AbeGILWLzjTkfmqyoFp2V5fGxLezTICRqpPxHbDEQdyNrhK7Lxh1al34hq3G
CsxSLimnl9kTKi05fi/mt/IDv4cpSNwRTmATAFfQO0q6L0iqC0ySDuGqJAZ1udYQ
ifIy2LFciKjgLvk9dSbjqd+0EVRSkZRiXl40woYNtIuq+z0QMsOsiyzCOXitStuZ
e0SXmKbYfeYmYv4ij2Bsnhw7Zt3HI58knlH6Y8a1dUj2XRSMz68thzbKcnSUDuKP
O8Ny7QbBXmaIhGp6luJT9Zm3yTQtjZhXOdduE7FrAf9Jvtg2WkN4Hfkbz3zl+Fz6
D3rPY080XravJaD4/wzpyaZfDL68uhgtH7h2L1UJ0Fjp8NW8hnklwQSa7gfNol2Y
jgboCRQ9epiFFUabydBi319HTMh4x+oBYY1QWvqKEKzMCAijRMLvPQeiC2Sc5rfP
RYh5ftdeuHg1ueibA95aw/BOiKynmXNt09aG+EtvcTdQZWYr8de6lYLwDkDstG7X
iiWfZZm3TifqR5MNfH7hichTx+XYgEEB8+eB/Tos9/I2Tr8SOr8QQoVb2AIuIupX
gN2YodbmdUQ8kG0j0bfcRKQy5V8pR2NwLqFMKPVzO7+UWqD25G0QQBpKv1O80pBb
nfXv32KNqzELXd+ym9CAVVYBuaqe//jEGZwH6F2qHY90ig22OSzYkF2dIdvOsjyh
LjYH7Y8/FssexmmjpLP6qK4Tu1g45xI9LAQRRaqbicFjr9fzqmcSChUvUh9USDgN
hkOEqHTGK/EywcGh56QT0igr20MYCyh+SbnVo7poN2d+Jmrf7CF2oanI6GPCIRjp
zkjQ9rel46T1BrS6pudFCXejJzIxDEcJ7B8KBBqoq9oTbb4ZQ44LCuZdA6HhTqhw
gShom+NVqyLLh6RIUOnH/sRNRCJaJgImORgteVmSJeptdlZKny3KoAPj8lkZp8Xw
Wxr7BguSj2KPkGMRDm0OjwvBav97K1oCqUFM/5mcztUTxdfYXULE0GA/0eRwDoOd
4GH3vCMLcOU4CwBSQ/ukApblmNMOgsiEMDLnXxl2K/0cxxQ9f53fid8eScHNVlTZ
Cka0V22FhBZ3Q7/yn0NE8xkD4kG9uijC+aj+lq/fHMdx+LQyiBTMQUKYYj6did9r
AA8zfNHN99dE+n4jVC0kwSeHGUTmv1g57ebIs2q3v4GFvZI3+lUQ/gK+SMijlu/A
nDdNnxbZuNPS/H+7yyz6JZAsT4CUZ74bUyZQ4wF5r1t/YZz7sU8IE9w4XvlsejuT
1cTrPcSN70tuK366/05zLwI+Htq+5U61E8tls02QBoomkR4OmfkELHI57kOEg7yJ
b7eRc4v+WGLgg29EF8rCqU3EKZt00CGa5TPyLr3ZxOs=
`protect END_PROTECTED
