`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3J1kEvs2vAeJg4dnXgqpZVQrHs6EIPqmRoKQCh6SUjrGNo5uIwKoB1GRYMzeTJkk
AkZY3K0vbIC3Iwrx0UznZv9Iepvln19JbbdpdhMWB4cTygUKMP4o1+Ib91W6XcnC
krwX7NTrJCtj+klBHYZTQ4f1i57v2/uFX7A7OBFmZkKJxxLBMOdF9EjdMM3iS2xw
rNP9qRTf001nW4ABZ08Wd/odAcK6raj3Sd3SV5ZcagPJ64qCaOhzRihIPOAZ1iK9
LkVtc/qpFf17jZXOznDLIFrS4jQi2bk+rYJ6g21mgO88wsYgxM7+KXlo/hN2SSlx
pqLqI8goi9cijRzq6ujybFkKOT7VkJVwrSgX6AdmNrLCLIg2JGkOHABriUZAGaPi
+BFvnfJW1FXtvV+SnMJpJu83beKNzpYL6+XvHob6aX3TZsErBbPr2dpehd5PmomQ
APbrNfOGsR3rP4LMOuWAghbM0/I2FNI8bnAffr3YxS2MyXJ3Zf6apyXQvKCDe048
frvxuw0izYgZVRefjTidRA==
`protect END_PROTECTED
