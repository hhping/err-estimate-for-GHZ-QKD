`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hYVBMZnrRQNPaX1n6oNYK62YB/9+//9V1E2kaDk86VcFtDw3f31VGBXW/E+ugwmR
0LvXGaMVedOn307wtZixSiaookMM0L5k24ScYN0QW64oe2ln3MUhrXap9afTUU3O
t4lO6zPKOfif1O0N6a/elhMFsdeJ/4GDwqUG59tNQ8zDKOGnLEMrjajZuPZXFOHN
dadgQWZ94Q5YfE6ty/8KtljKG1HA0YgAT0AIqKEPkqMLls4pmpm5EyhGhplUiD4w
bv3o5xarSRgrtu/eir7o4FpYsX24judDHv2thC6OfEa8n9crr7zmHO02uJYWQ2on
lSUcPhh9+KxVVjlZfqo9rVR0gsioSoRtJccPKaq8FMuX2gmAKvCdLw8+R0lWxYJF
5Ot6B4yOMVyirSKJYySYLm8nnFvs55xS4DFFmmUoEeD90FPn4GTLrC6UOAg33bWU
2B6VfBNkOLUZTNXZvFxgefVFmrklDhWH3uYu1o9yFt6PE6/4S5MRYQb8fmrU4tLj
eVgvBn+n2/3srOLSA43Bl9IuUQZAz3NpnKdrx05dA3Okcx8O7uMYhgTMTllQjCOj
9EP9Q2ekTGbKaw3YtbyrxP3OM1R4p7xPL+v/MUusIvmi+8BQsD30Zo6gGIzYS/rc
GD1I7dNE2WqX1Iuh+HOoCtU9kqNPdM7P1GeSeN7DPkGtBc/tV7Nv/RkUkcH/fv1D
jM+D/7o5lE37I0nD2x7TnwVMunrQercFIS5ZdUNigLmDLAPpnB0AolC6XuK0x2jb
Nm7AufBkXMK6/0wvXbFW0SuzIsvuylwIe+nn3uIDW4FXSF1jpoKGWsX1xjYxZRku
0n17Xdkr2bYsW9+0RIjfaD0lGQIXtt7Y2SoyaxvCJursV2MyIRVy2NBbPw+dO3ZH
etuMpCnjYJduwZ4X8NFap7tS/zgaRqFsMj6XCYuBDJMJlNOhBtNLpFieO+zEYOMu
TmBJtkzKo60L3WR8rU/8oNVTH0xWMfnF0SWu3L7JvA113nJPWY7kjAv/qcsQG3de
9xfZkvPQ0ovltiJY+kJe/gGbZdzccMTAUre9sw+n8k5F08BqH4xzbgLo9RPuo67D
vucvRoQZKeLcyYftjZaZqenyMEPY1SDSc1Q/1jBEGXl/lRJUeLyJkpAG6Df1uep5
mcmrbcq16Eh+u0wWEhAQ3LA+DX1oaIjl1iU+TBIRtOhiMlLI6QJOKIL8A9a5H+mJ
6YK5f96YL48++qtcObg7jI011qeIoqixDoTJjvToTk+ugfYuTDS56NGF+nGmmhgA
Tor6LwrS0kBO4LYr9Klgj8AM3P5aECFF8zjQfeYKAE6C+nHC8gUgXZw4WaoJDlSY
k/0coGeUH0JnSw841e6xOVsNW81am5kTK4VvGzfKZquLLnSrcXgy8voB+F5utPtN
sVGxklCvICKbp4UXXIVrJWhp0ov1cpkoxMIXs6d6LcTGOkv1jz7LslNMe/m2Zn6z
gWB6r9YjSCtL3SO3Ww3YhVo7ZhL5FBzyMNRI/RrMdsqlC73w/L1ounK6sSx4mxUv
EPLWZOIfNo4AmCeXyI+8Gv0AEEaXBTmF6ET6ylKYEF+zQnPE1KHO/cLrKJnLNH0n
EivO6PGIlOBXB158SiBBNooqsmJWsJeCLSH5g5qzfTrBrXrc3uCFqzuj5iHAan9a
jvG1FospKifBVGqGUN8J50okzc3FPFX/MAEugeK8Zi1Oql70x0eMJmb5yrsEcOfj
VzE310ZNTQW0QWiQvSQa5Ct0qDqFEg+Awhtx0iR4Li+GibsXn5KqOYjJURuJrycm
KmZUpQ+CwwUR+PMcxPjdTAXS7OG7I4WavbsDGBENcpydJ8vD9AXF7rQG23LR1vzx
x+FE+KTb9cm0M2GUtdbuU0uuatf+/HiY6Ms8ZpWKBCGb3ufkTt4zZQV3Zw7Zf9Ms
`protect END_PROTECTED
