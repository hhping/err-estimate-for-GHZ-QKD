`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rmv83zxqONia3RAP6h2C5+c9UeRlhTnH5J5lAhQwNZ2zgt+e3adDcX6eGM4HXX/a
VAsAxKFAv35L3myjqZFn5yI38tu+M+0uk1ja2fIUl20LoXsdrfDo6fXDrtcdwIYB
+IRrwfKxduo6QIlTglW3BVXS3U7dAXmNju14IKH6DAx9+H8YknKvHB2Fo2JiokC2
DnXjPNJukefkKQk0gMdxLuYQf7xeGhZ0qss8dnoPgXViqLrQOjpYsp9wydTq5Cqf
AkNehZoyu+lNmtJP51mSEw68WJ5S8l6T5JegQTdoz9TAD0GhSfOJ8TGgj9wOEHXg
Y/Q9BGZtz5+njilyLn6GT+4o3BMoaV2e5QvLWDW7RMvZtjorehjRKwfcgna7WRr8
gUtZaFW543ee3yp6FPddIgFFbljsPH4heXhxy4dCmg8OKJRzsBtZCL9DqqCZ7B4q
7ABTS8mrt3wf8woYJs3nUvfF+d2ZWUHNLhbOl81A0FESthAlYSkxkRAHAHfQ23lv
qiPn69u1EGNO/e4sl80RBUA7J66D4lUQW/kex8VnfWR9NKAJ93wyuBoWljkZ/DMN
9SNZ2/Pto2BUyu/uMnxSC6CeKNLQlzT04qY/WKu/cnPYG2AxBN4B27qKwD6lm+y0
M8EP7G1G6WVylmH88PWXvjL0ft4wTy2Yx27hwJgLFSVje5kPQhJ4atRML61hi2Hv
7y5pUZ2dx/kNKe32ceY43k+84K0jZucezlz3y0b0SEyToZsW0/x5EAd08SZSlmHR
nRzYmo5OFyQ4coXs0oFyeL8xbjPM8WHBrqiVp7JcXZDD//ttI5k4z4s9paNFTaFp
XDHWYlrtGa5QYlnNZvwNUg==
`protect END_PROTECTED
