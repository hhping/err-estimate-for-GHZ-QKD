`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qojcmqzjb7jlXqs53P3zM4tnU1qzBZ53rxan1jU8UaaZMtKZQZ7cOg0ruY13JMTf
AJSopip4RfFL+SdfB1bYVkiTaROwIGFKOyTWH4nMHEPs7B79eEQdajEt1r1ABVH4
iN0UObAI8pg6f1LFkBIYX6cDFU5ss/AXctBdbx0sLQNuEUghdJckdV88PPl6xqkz
tcrDa+vIHY1c+3uf0jhiTr2Z540EH7zbjdbZP+30jLGB2ZakmxrOguICo2vKWMdT
pJAry/DAV3PBeAchtDX+TeMqg2DD0whWgF5mV6swsrbStJCFG5F4BRu0Wi6IO1za
2OD3lZn55VPm8I1WpSZCDcKhN3A8U02VexkteGKrRr39iwuBZkydZtD9IAsl5oBq
h1WoBY4U+SO3YAYGDroZ8gJ78hD9NGnNPmBdOiOPczrGVot+wolL+W6qFH1Zri/D
KP/pI63SiyHJzDVfME7C5+OPmuYyqyxvkvS8egnTS3SgN2/N/gOHS3J9d4C5u72P
`protect END_PROTECTED
