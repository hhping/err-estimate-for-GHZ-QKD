`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5zth07HsfaII3J/jWCR+desm4CKj58+k9NYFlhxZOKssiiSTT+EPE2MKRCadF7z
qWUMLjwqXy8DOb2/bY8BgfIVLwsX/TZrF610MKQdrWuPwoWeQ8GpB6MmUKqXK9+h
BPB9bNcjj5ageqkbWYviVvKyXWrlZEk1nsd+4ZthBwWKY0O4Wj+puMIaEJFOvFd+
yCMA2hiMCC26xnfl5sAoz3zkmHskE6knjmOJntzHiwEnpjKk8/fRZvXoxIs7R64m
eJ7BgGuT5d43DTSYeP8iRurqw02h1nTPsF5kMj/n+sHAJGDNhQLMcepo9yD67xjq
XIHj9GbgPKnE1wb4EoMFvpGM5FczOsi3zMy5Ma0Ilgk0SrL0FsPQxbX61wRbyWjy
kueHf3MB7kWGB2J1EG3bVTVvwlUd9SvQvhhNGX6J3yDHgwHAe3T3IcWklyj4RsqG
E39Nu5E+MzL/Z3wf1g+NKHtEHLHljBGKDsoRH2eW8JFg/5BEO9xyWHvA2r8xH8d+
fg2n3F4DaqgQ/x1guBtcG8iupLKYUQk+wHBSQPrJ006Fq4reJVRQBVdZ0K7HrKr/
nPnKfM8ZxeYhIB6RN8DrXtS0DxRxS+S3Sj7mkMix7xe1BO+ucRzwnbKQhadn97Dy
ZGXkfAm/dvDp/grDLWbjWslPjV41Zkz/D7Hbe13xvmrh4/csb33Vfrl2qTM8Enna
7FoR6+30fx9Yy2nhwyE3Kn99e6mmvsLLRT7KJ7r0wqgf+tKFgxkpB9CJCAAZ824S
QaCi1P2Ty5dwmBxzOC2WrEwIA8IDuRYgu7oTX2HdETTkJNJxAsZu6r+yaunlTrFo
p2NqimT5CgrcaQPMFY0+SY4hp/VHBjdL38afTAuk8kp03VsG9wI4bbVLUrfzn2EV
S3/NaDVM3NLUi0KQ0wnAdg1njInqurj9eRmZQwQVVVzp21cztih1eGYzMdSJY8T8
fOy0hQR6ID3QtfhMqjYmqgiXObKO97Vl5IGde5mKiUOguqIssN0LJoH957Q4q+O7
2mrY1Z/GXOylTGOitH5l62WIfKqBLGAXFyMW1YL6eHoG0bSPSDfYsv6uXjjpfKlQ
Jhd3uk1cb8hETQtN5o3LFfZo++KfwDUyJVGKOGNmXr34+gfxHJ6FY6aq8fKLo7Wf
Cp5jarieU9XkhPIgB0TnMRDaah0j7GsmXUMyEDQf1d6MjIUUSWkQt+lAcy94qcmM
AiYOpNuNdpkI2rTPLmq+hinCvH7FXjXYAsDh5jdC4CTaRwf7B4Gd+ddJuUCGiPCK
XEpbzJbvdc3gRVrR2Nn3eRvSZawJLtcIRzUL8wnF7t8=
`protect END_PROTECTED
