`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G4G3HmPKGT1uWCM8EvHkxH0phnqE9ZwEVxk7SdBYMFMwAjkl4A/XYUqAy10kGh2y
QpAmxr/NKfZofAfSL5gN7xPJr1Px+cauqQGv2/7DWtpMOQ8jjMMpsuMvwW+LKUum
m/HrQLyjimzFEpUMZbPIoVTgUMF7YVo2aY8SDcESIMt6pSGwtppCf2XLSRLnQ9nz
2cbLW9rI/QBkQ56GHWTK8PuuT6tWSVQod0+1/AfdLfv/gzGLaIdpuQlaPFGI8tpr
Q7AwKOWQZrZnHc6CrYhJWCiGu/cOi0lU7VAQ4t3u5wI9wAwlx4p2XzbGcw68mFaC
9OCM4jsRrNeNWKlaJZziPSnPPlYyLQGn+UPMWmKXoZFXxiA4E2u+05fXrmBxK/av
qilrVR2X54a5J69+h90Nh2+bAf1Sn57IHtTblkx8o2xLODsNR5Z6psXe9gyaU34r
Ou3vbdDYJigSAkm922/d+0ccDF5qNtU7d0g1oIMt4aOnDsmY7jEKXMLQJifq/WsY
MDTtAwWF9ABYW7v3UoWZ2AZSliaVvNtgkhUToNu2xbkPaBW6sgFpwFPm5HqtZLA8
zRltQjMUuGnM7T0WhrRfikeRSHkM7h5hfjzgA4Tagp3zFj1DbiKU4oigfcqr4qqh
nAlKuyWe61/qi6oITr1I44klcOIKyAHG7dHnSR9kF0pUm6KY5HiIfvKDU+tPi1Is
CfiaiNiL6fWtKuwQ83ANH3BfYCMELnMHi+V90zHPxz9YAuLpOuBwJb+LX1G0ItE6
MqZzITCq1U5DAoG8xtizLBKZjxSEza66VDFRrVafSY4blykAmfOrrmyw29NnqsuT
oxB/mwwgVStnuxg751mVcMcbYCyKcSqEjV/ELIBLoM7IIfD9flMnZpVyGk4wV9XC
PFqVzjEEYddrA7HorLIPnPTeuci/IQYZdJ21g1hXyFFr0ZubfZV1yR+1HHobRxcj
/tuui2QrJp+wLtc2HeFGb0O0U2q7bVBglDvgY0ljRfbVto+A6g/fpyJ/uSQNjbAp
LCmHHYgJ+W3AiH7NuFykWKsc2O5O825dnFJn/U3QdpUQynWWMyUYxmazwhQc68/p
Mbi3jmY67dpnambT6dVuCDT6OEBdpq8L1Spfl+gJ8gEmjuuKvpRWNW6jdDAIhxVT
yL0F5gyj+/JpQnAf+Mb2TZlqPJhbYJf/WsPB8CJnA9lL2dL8Dt4f4QEx/kPI7K/v
NoOmXEOlpDcYwBb/V4H0A5hQAz5FD3wahBllTt4hjTRxTxpfBxWNK2QvdffOeV5d
cAX6D+PmFFQp4ZB6ul9dgM+tNWwMUe/6hff8djGo6DWP4AnMfHa4KvXFaqr/P6km
2u6kXY6StVuXCo9wXsaH36yuM/MYi9tACzp/GLhttrrl8uj3pCfyiqaG2KCkpzW9
DJXMasCJ7bsGKM1dq5cFvovZGT6bGC095dLuXMTfwVxx/ZxCVfvOwVqzog8XRcXm
zMW0vuMTnLQigE/RBUHNXG+NOXLWgnqg1oEIXkvaTxVeMjRW2m/pz/e8iKdUTcCz
5dTK7i+FiEfa5W4XCdcHU0GSRPImzuPPNNYKp4qa11AJLjqGZxGCihlESXA9KtQZ
zRwSyvMOpb47Q8eDI80Dulu0KzT/xGNs5QjU4nP8BX9oV/lwsYiioEDbs+UXDerA
NxWgpQIZf6oazgOkYV96fvu4DcwW9krzNRN3ZETQwLvpcbmvpE0j9nZ0nkxOVcw/
5LVgfh9RRGoqBMTNt6pza9Qe7TKmuTkCc9iHZ2IwWQs2e4raPykXomm/3DEJEkTK
oDGNq7R+gfmJaymOjT1G5k6jFHrFVcsY0V4M8EAXnLLyEYTSqF6+He+PNQssQLbV
OndFKv75KXpkGbsG8y2sRsXxlETkZ3M9SGrfnUKoWTANMSClt8Zp6rB8ioYEACND
DSHqs3f1aiEOz0q9EfyIjUcpw2ypp7Tu7diY7X+F7RHETOstmbdtFdc3wAATd3M6
cYBIxuKVzj+4rShc70eIEhZFTh2OZ8ctddgQhiSelBlZJm6YPNlwnVesz4vYrs1L
lV9pyvuvlj7Xc5qti+9U/CJ/VZrdK5vo1TTU8w3lyXQTXgJZRNZycRCU9kKm6aUT
F0SnPGMTix0sXaDQXGx7jMIUUNKSAuvYuidyd7VOLwjv6War611sFsnY2GaxuLn7
8Ismn5i3Oo1Qx4+AvSehfXN0chwLFiceTpo263lQJJbXeHGKz61dtI5vBtLwbLIS
0PPHBF5e+UYJTvrObFCmWq4YM/0PwjJ9cm4LXaAVZY9SBma6wnLPSyiE8InavyC2
lx5PnnJ6WytAawwrToAketaAHDieT++vMGBtPlp2MmK3cycADEEaZ36rYe7L5ad9
lTeyOlVx+6rQC7+TtFATOA9b92RF4wEn5rYZcJCPkFkF8DvHGuOEwhYOaUQFlLSx
aaG7A3ar0TeYvbU/gIxDqjzPRw+BxwCWZverrFnplv43vwdOadWwf9Lx6zCzWYO9
YSe6cH6AF5MO5m/7sQIcsaYQMY3qZkq0sr1ynpMi3tCOnbhSv9/DGCQCWwREm7+H
uVyp9Y/P2rOc8+aocyGRU58WaddNTutvLp0ljoHTmU0LuZ6WTMm0d377lCib6KiO
Mq17XHfj9MdvQh3h//aaYvZfVU6I9/vM+N37aO6j9W1fIC/quKXGzgCvvHF0cjjf
QhE/DZjLXdyxi4fDHxUMhzuuZfYcpDP4trCm77WqVwp2jxVyLAthAMUMDXCnsVPj
FpiI+RB6aAeUpUPTiso9a+ztatEHcTOv5iVBO671EcLEkd8ZyL2xak0hXJQ9fDg2
/+GZtr7eOLz1PpvEyrnUinHSmCTfsDuLGWy3hihuvtIFihwva46RScvk0Yz2uK/w
5JniL1Zxulueqwyyjs2AUQFzvXk2QIS6CIp/8XlLnpb0gEBDN7n90bFVaUDccuKw
zvYbYnNlFGzZYlRY9wkAV0EWNttBQ9236gogats97ifG3y0TOB5v05pFnGuwD6/V
SByNF6TwHd4xZyQrzC5j75GJ7Nt0FpLtsWPcj7W22A1a+ek9tryA/tSphH+9mxse
4CULFS1liDqIiVxmUiWUUpqFQKOVaYcsAxLLYJdVMpXxphWI+J2t/AHHO1Q9xTsl
3zuRAD4U8z44Lsd/3L/NPmygdzm5mpVTyW07CPV+hYYgJLpcT0Qhk3BkYBEfK/VW
Jr6Qcc2sQa1FNZjRwhaH/TJyYq2G4nH7B5hlbcz+qJD0EvMiD9nexARaISJwrgOI
XrQVRS8CsBPktM0fYp4bj4PJLXZ4Va85p1upTbQlyp4VUkZa1xk0WXUm8diRHye/
Tn6Hd3lCicfsrYkFLs7cHhM9qF95l7FBehskr/mHsdw3mDeYppEF7cFZ9FjfVa9m
DfQpRL5lrQtYIJe/OZN3Q/j6jU3kWjEv0zKNz4q8QVJxwha/lsD/Yp3b0FtbHP5E
j1SzeMCZ7Ii7KgoQrUEuQlMIdBZtp0zt+92BUtzzCGiuWMS+2EQhGAqsfGdi2HeH
PjyRuMYcxHFDOUXm+vbqs6VJD7Z7qudi3ax0TvNOnf2KXb0+xjU7NKJrX5fjarZw
WLIkWDFsOleTpqQOgKpnWEGreGweN0EYSMOMAKiYjdy0A4p3pTwb6NUp24ToCPR3
uOYS851wBGrydi3wszWcY2hWsPpIa47S00dlSQeyn6v+DuxzMTplhQ0luPPLNepL
3SulDpDalmRN44/hTIGr3oDjXky4+HsembM200EnD4KLIA4k9SrVlE3Tzp+INzq6
hH032LpNkQ9kV0KC5w+MeZwh5hlTqWAaU07aCr4AuqpIRFsSeLO8xByQGgDtodL3
vnQ+x0NHojF38sD7mRrFoqZ0xzqB7i4cFy6EspurrrcRKIkjmvk46lm5es3BOyQf
o+bWeMtaSmAFbsROIvPaPz6Qy0Ob2d973WSeTyEnyVoaGecI2CI5qfpDCayGBMlY
zfyxl30NLYxE7xY/J0xy6o2yxdTTRFT+XLgdpKoea9rJjCzCY4VF33FEMCbCstRd
`protect END_PROTECTED
