`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDhyUSEREuzsTpbhiY3zAZ04FZyzQeMhCC/brjqFQbRKVxquYY4ZS18Wgt/m8UKi
QK9N/1Kn8x6PeObQOLqX9qs0+HGMAsWKM2PNcRIAbfe+gyQ/2dweLWXPBr/HFk3T
wL8+KCT/4K7NTu7PQl1QqbEO9T0u5skLRrkcJWGryShGJhHvgNWxAVAqN5iK+Pwc
ssJSZN4flV8bWwr3ANG6dkYpoUUZRLJudxMYm1iZlhtAUIhy/Gg07Cnp97GEGHoY
D7Lg9ivLc4ZhHXRVVQXUXL9jRIxENDuRHuin/ZHpQQ8=
`protect END_PROTECTED
