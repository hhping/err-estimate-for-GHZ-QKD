`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmQlR7ERNw4JOZEpyYc0ztLxtt3t2tkjnl58v1+hNtoQuczaiT4G7jqUhLDt4vP5
72ctEQ4rnAL4+GfU4lmDE3xbpR2PRSqXyhd57Jvxj+YfKGik+pfPneDUEs/hOp39
F8aoKOdoIHmfIV9yEiuwZKQqHUGgJ+B7Se3xJU7MnIl2PXZxKi/Wi9U57XJWyPI3
EnB2jRHE6OUkkxJfFy+kUZCBISx0HksejMKYGzRKSr/Yw3VjFY2k84vptfJlrY45
PBE4Q33AwEV8LJJT4XYCGLgnwMP0fbp0e0NbfYykU/rbpgRJdotWHmtkGcWJ21ve
yIa5IBmwwz/rn7PK7ANblOMAl6CEW+0x/ZbzLrMl+l2nytJ8H22Zq71cZQcDJSBo
1QeL0O7mQO1WtFbmNqVyXxHIivN67woMjR5tphuvLNqzVLUgtkTWebvvX7za2r++
QZTDf5Elfnsl2Gi5PCiTpYnns7do+bd6tbZQDOhgHfxEYWGWSHIOSB5u/1tlckm7
qU84/HJi0z3fdwQfoYAwEnPMxRkXXnd+fUBS84g60frdAhRztHSios8DCRzEEK3k
gv3lZbW8NcWRQHzSiF+S8cRrUNh3YfsgH1nDrzhZ7EsNISwhLjp/HBDuvZBmjdZX
Oha2hYa0DJBGM1UODU8p6olQ1JuBXVVrVPwKGAzaI2XGKCZS+Vtv/bp8Z8hpdNz9
nn1fYRPaszgJkkNa5St6YKLxS14iDZzHvdrYhwR3Mef08S33GtJ7GdZhssm4UkFG
udAiiuytFjiDNOEMqsT43axBSVOe2Ab8GQGOsPz6Ibr+vWL3dez3zzLF6+nFgSR/
7lEBcieQ6QmIujUwB1eWyTtnXC+VxEgo4RMvdW4mHrimhIbgNFNG8bz0OPvVhL7v
byzXsqtbCzo0tLTtLYiOmd1EEDJNsqTLpBXH4KGBbeTOUwxsSJuwDuLg0Y2WDRIS
s9xYr+67oqxgTBcs0PP3Xfh/DSWhkZbGRl2tcxCF/MO7ehS7mj9oMSEWRnOnuFEG
dMIwrkSlJnbvaRI0DLDW/qIUFzDAVN11Ii1VCqdSoFPkKkcE1QUNpuXCBAjrv7TR
FStUp/aDWX5YwrFcz4G1Ps2SjWi1j5aiHYZnyccNEpk0FFmMP4dQCRosusvpyUiS
YfkJs951HoJg2Zg7zR0ZfvCm/MOwhwHy/roqqqLgWawmyrzSz1lVl6VCMt+8veNx
yImuQJYbls3J9LNTicGboDI5yN4OTKAK7vBdm4QneaCSyw3Bd5nScph2bCG32RqW
PYiyFrFgiEW7Tty6kHIAQWp7gHoAtvPyJQJA8EQZ4DvdJqg3e45iilnS3jAUm8e5
yp7VykvexAcK9zgsOfkeDyYMQ6Xalm+CG0BYnt1mbUQPD8je8qnte0avognrLE2/
76D9p4TKW1RosRBMJOinTQ==
`protect END_PROTECTED
