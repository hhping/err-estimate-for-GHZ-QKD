`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVwXVECH4Gtf1VJDzkNgxwjOPjTpt+0Y+9pkHeCDdeBYDEk7VmF7T0szGCgS+j2E
tc+gRZ0hFgNpOisxmQdNKalOqJdjpHmdqE9a8PhhWvbL1UcuVfEitvVmHfgLG9Fi
b8lC/ywfOfg6b4400k2qZfTEW24VWo+JLSdMdU4qj6cORFy/MJDX1DSuKkCyVxOT
nSisNQLlfcmXBwr6UwxYc4lfcj80rDtDbOaz7ru5BCkb/Y2jbKapn8juG/QnMSil
62CrbrXrPA0ZShZ8/pR3q4FfqL1Fruu0ax0xIilkVfgW6MZZLb/7IJZckw3l4E0x
1RCfWePBF7US9r5EMvCl7ge3V7bMhfbEv3wxxRSdkD6bFk+z6rosuw9Nyp2zJ1sY
ooQytIHv5rmDDu96mVVY34OTCyyAZff+EIYENujVeVAkPEPzuxtJ4IIcMtfslnL6
Fomi0UMESbxEbtv5o97qCAhFQKL2M4xyeVFaIAfcluvEPQZoDWWraaQNg9opnSNX
4RWMdvKjq9YNekfqzCEwzvPQTGfchtZY3oOWgoOCUPS6VJtxJA/fOntIVXw1ETDk
azQBlI+M8qUo8CIVuc80FSeQpjmnP3IicexUZK1J8/EqT/iinbdJtFd3JJQTO9JF
XESIRoxy0npVyASpwoDAjivSy+7LDYDddVgvOwPDOSjhYm1ALiVRUib5tNv9fgSd
4Sx7wixbr1btM8pg5Zl3mOx1mWKrJHnjB+o9CrjBrmVCX5MMB0axG3ZEOhgY/5z+
BIEckhyZjqeRflVuULEGzbOiYS0npU1xusiREIGmAVuwH4+sTSChiqBlgh3+I3F6
HRv8A3SFvfUPXaNE77ha4ywduBGt0/QuMJp0J1Aw+9krH2YYJxYLnLXJBym2X4pa
eiU8cVwtzzjNltss1us8rBUOK2amohN7Vcf4vO10vxVBz7JecvYnZIiTy73KDB2X
kFNuiGnBV5BkfC6Ej5BFjKbfF1DFWjO7iOyyF+14BtKAjr6bWTCEzeV+pfNp4pS6
xyVRX+UbZDdjBcbX4uhpeJ+2VaI7jCxISrTq4ZnH6r6rP8I2525VGqqq2vXiUMzp
8pSzhLuL5lSkh16ouXl+wLFQERt8lkU8ODH9Iy71JR/MT3xGo8GBuEU3BKADkjPI
1lxK879dXVPHQ9EZG4bvh6spaRxxNUwcvb25J4uCrJtTI4fru4NvlRm8/+DQXQgR
k34cPAcDY0nC472+rvUaskJZ4N7kM6FMRDZ+QHXsaE6jMEdoHruek+kvoOwsHGhL
JsOL2AhlvoDeZ+w425InIMEca1WXWDukNE6uufkvOnQUwqNMMUlgzwBr3ulWyigB
8LtaDLzjU28bNwroG4mIGu11JgAiwsLZVBg5rn1b72zkjLj9G9O7zLEcOD6GV/4s
NMDiu0gJ949VlPl1kce0kqaSi37tohhOZyiITYN7ayzfJTb8JFTGRrB898W5/74U
URog2I29fGXwAlyZFDDCToxd6QhYXP7iVNxcyua8oOiFhkECnbDN1mkQuhHIxWmP
4HTV6KjQUnpQYb9ShvH9q8nUHmgEhimt76dMi7+q7YRVL9EH4sU7xe+xRDDjBTRk
7lcPErpMpBZOQlPGGVExIu9taucWznuvSJ5KDhL4d1TIBlFgI/LO7bDHc9s7rAsG
fzjipQbGkvPSxr9LB3bg572JVz5HWHGA14AEQx9ZYETswDrcQ25s0GDhYUdLDNUy
+1hrqwOXwW/eaCeVYGBm3UUQlnGyJV3oqYwWkwv/9QI93PS7aI5nm5+LYchJreuy
HWxUD+nO2KTE0lmhCLZpZXErGQt9rsmWFUFmRetIXJ9BYTDK4oWHz+MKftdDa0bT
iutwAPATqCZsbUV9Qgb7s5/zMItOTKwfbOkDfguu2uqrWxiwoNumkpr0WEwrjD3S
2ZmfoJm2hyciciinXWZKgUTf7sZrf/m1RzovJ1RJSpl3v+mLeNBt8E/qinM9GTnx
cco14GctlcFL55qK2FOQ18ciHQc06iadKqLPwBs4UbFkWJCK8/ti6NiV7XMpd6aB
Ti+VxYo67rdVFplEGDSwjXF20q/UMcS1tV0pR8u9H86Rf3IRwNk9sIhW6N9oCU8/
6NuzXMlVIFKoScFGUi8IBhL8axxh9mnzaATrwLQQbKREA75oAkysXiqLDDmAtw//
jZMIYTNmWLtW9An8jkRNc/H1ekgIWMnKO0wWZYtKEnfwbzhhoElKcTBJ0xnDOyyN
PJfT9U0CsWW60ql8QSadeLVBqL7yRLsVNPzShBSLhVLe1fIQ6oi0UUxrRZy6SpOI
VUxyKnKAecZBakixTzV+zVWgWLTIMurD0rcObfyzjvzrDUcAaYLgHfkLd+m8IK3s
IlcFSAemeXAwZ/cFLf+N6haMZdKa9Z0q5YySNzq+KxUoeAFhL9Mx9606uWUMDZtJ
+yrszy3WGCrZ6cFIpkA+t0/7rTxIt8mXzfrHd+Hhfhf2sa00mwPzHsZLddHOZ1Kj
5YpC4rHy7VkXcXCkxd0ASu1x+WIi/dpWWt3tO4aNm6FSar+qtI1T8j1I9KBJAY5f
72jmqQKqbjxgGf3SvrmnghFFfsoG+lcnemHkyWec52/W8UDFZWOZgz/ljJEEt+4+
oPyRbUc9ASPCCgzLgwjLl20IqWScVUtZdeC3v44iBj8jXUyIjo4rNbCdZOs5JB4p
mo9VOpFg4OW0dKWyoFbJpjsS25ornRrTaRox+3D+HltYdMZ+Chc0axPS1dSwm2Rv
XUnwZcbyaBu+XwyqZry7m1AhtAc6fR/cqEXL+PDnxgBYNaNlBwzFtAaLPvJboqWP
6kVXLg6qzQNuaLYAM4rzJ0UCpY6OANweio7a9q48tCdDaQAjcv8Ckl1dvVHekxtp
FBLa8TyGEgKepsxr1dL4qxEbhi9C+qWz7qUH7xTcYPuo2aO/dNjf/lmG6rjkX8sB
gDithDI/SnbEuULTyXS8/7cZqLPy7kcfSF7BOBZRHtYAfJGhcMSQKkyKe913KIbJ
SMff5w5X1DJqSWSWcz5Kr2uftdrNlE/S0Tc7NOIHS/j43VTpKVD17Jb94zZeSp7D
YvnwuWTOTIHiY1nIm6OnE9UzxXMzGCS4JAf05LmSjOsXBfX/mrkdR4dYNjX5jiS3
buE/hEW51YmHVFI2f71RorsUjP+GqLhCpqmk0aLtomjfqjW+nr3tkWidCXiRLWZS
3VA7LNmC5gOcGOjBXHujy9kx7XMdvBK3rASM+ZbHn9PEMYNPDjOt2olJY/Z+Qfjt
Fevy5htVQ2YAWfRYz7xQdyPZUJCi7Kw8iSZy5bboKiuNcJ92TK0+yOxcOFRlf5yQ
3SqQnSjBc/I7ADmdVPuMsO7mlfxacJ4y3C8tTWgf1RAyjyw2z//M+eAJjMnWuwR3
JG63IZZdEbJjxNWqRQ7LT4KuyHtHg29pohKEo7R6/jHcuVLVAWr75uFpjRTu0+yh
5Xc6OfXO43Z24XRw8p9kDPeT/mb1NYGcCqO64Hm00klPpAxrumEHYOBLthC6QVT/
5sGgWpB5iwchv0hKhg5o8QVT3zfPllNoJJzaOLuyTCXcRWExu0+blQulrGqSD6f/
vk4gTyKvshtur5cTNkKZJeDAUxTkqnWps5a13kNagFQG0/k8ltLtl/1FKNFh5IJD
viLFhwYAyBM8VqGg6b+26UW1igqjREU6+sxM+Y8pNFd8+JKxu/O09D+iHM3YJ+8A
xfHVCTJOkkFMmtKM5T9K8ZxK97xG07f9nSr19NDeu/I6Vn4wrvxQwirCFTzr9EM6
MCrZJYirzWeOqrOvFXWFxR66F7qIWeNf/3YjC3hddEF9AtPWwAQGLb0GUWGKKc2Y
Z4FzRtkPPD1GK0v8pLFIdOEx45XN26E4zkfb4vThm2qkwib//QHt8Bp82w2bNf3I
ctCmdVNzlSRCO+sXeTG5B2pqBKy/P8seqk2341j3fUwWYf2Sym5kK+DzXtoBFltt
MQa4wObsOwa6tcbxxaGBIWc2BxeOVcQ/zwRat1BZYJ4VGhPzuOH5W2SD/JUNN8UQ
u3JipwXhrMPLwXZJ8ogZ+foFj44PR5B+jLeCMr+c6G81c963IdWTrLCUN2VW8MrE
EQBIhD4RC44lG1+iBDZ1Wq/TlrpUW5gt7LWw/cRHcHNGfgLoXO0poyLWv0UZw13d
65s9n0SFQsbooy8EJt4eLnMK8qMokqNm1FjQzVlyMylQGjKW6ik9gZ8uu8OOALLO
U7839DC9WHEEFVuLbKeRxVK2xYJZSapzKGT4NsBT3Pdk2nW63wlDnHL+kQLEYy89
sDH+np4hpCLx8iyFCP2Dei1OIDxmkQsl3LKj3TKBnmK94dpj25ROyLvs9anLXT0m
4LDzX2K2BKVfvxO/+Ol/59GJmEomZqXPoIaNKbChifNALyYhzdHF1aKsRybyMRnW
TWwpgKN3D3DhSnxgaMM9kJ5Dc60KSc42GUkqHtwej1v26YQvvxAdw8xwnb5DF5+9
iB9NcuJDORW8wE0jlqnf6HTdGNEcvS7c2D034uqbOLDbiJRZmNA83Qhcybs2tiTz
9O1fZQnJx8uVPFTbvA59gg/BYbU4JU9jymZUpCzSsfv0eFpScdsm4uX/VluSG6bo
wfK5PlpjzUQIITaNh68Zi7U3I8xLw2+lvEscxDrjzDZbL1vEGlsHvhmr0JsJE2tY
JDmCrQkv/mUY4aSdiLFtcLm6tCTUwlr9nTOBS9KNgxN6Vne4G6Hfk5ylUTzPaEOF
uXVnsC5mfG+UGCkxI6bg5dOCjzkNJNVptJ4JDLCTZzAobykUu5EGjR1ZV9QU3Q5f
weEx/RcKwviGzHLzn4QjbR+wUNmidX6Pdll+mQpQNjkrtwK59yF0WUOe7e0/oBc0
vyPLOXFHEQRcpob79Fr5LdkD72wAOBCNQ5vjmp/IhjZHJang7crB0uU9g2H2rh+x
Y8yW6TvTtQMaXjOakISxKzV5cSIa3u8gQxCZKou/nGE+eL0j2YCfKXs+JMFeXRSm
Y5xcf5DYawfMQSX3UyOwqlayDi3gROseMRnjF0C/b4u5s0wfYQEAOU5MP8aPYUjU
d8kYRFYNdqhJKH1cfiVcZ6jDNaP9sG6iaElQwdvMUTCv+VZ1x35mYsJYeQI+CPQl
9q+HZfEe7SzcdbZo/riY8F2m77CcsuKPkqKuBoT74r/6l57cYp/7QAPsiFoYBBFr
C7ow5MQqdo+AfM+xLG+EFeWNIOA/NH3MkSG4aGbPtTZWwjcbmdpavdUNVSzCuONi
JMjcMMzY63VOhGq670EAFrvSGOWUhxMwK/xM6xLxegiJ5dQ/odixAdLE28GUrU9h
9FtIdWNVkTxzL1AQcvrq1Nj2B/Pbm+KKU4e+hLTnl7RuSBP/XMJ4tPyONvKALY7M
79mJmPL8yv58xP4h9UkPIVquDpk+eP3myDLgkALPO5B0ZxKEFpj0eXVAyxdKbAw+
5ESfrhwlMaB/2SfjnexibHs7UC6WvCDjoYpjH6p2RGceEwXsWf2A2VmZlV+ZvHH9
M04IG92+IrIO+6srbzBbiUbkePpRLZHL+NupEw57gGCYd5XVy+UN/Y+07XKe74ol
ZzNGMgSVbdeBU+FHz8ZY7Lz0SCEhUamFOFB7Myc3LvnGReEqkuCUmkoOVQSvOWGb
KYrcdcHqyJOZ8wBBBZD+xKSSVA2uvh+4B6D26ctb6RWyj1m4QaYav1EZNEC4+/WB
Kl7OUOuePi+yf1u0AQpPvKP5nk0EoY3/kxt7V62zFAjxwMhiKYa809H8ktNEQuF4
JTPthQiIUwJNjpEpC4N1xc9QAlXYoI0tQlkZUmTi6PU8/5LILDYNXLVUlVuWjpLT
asl5UyFwUfIU69sRxe/6ewsTYqGjd2rHyaq2qwtcEBsHV2woi3OZK8mMhHr1myBU
8gerZdCi+/f2KF+klj2/lsjRXjlmxlzwc3wILeV9kcsMxgzXTGA4Zn5TCeGpJFTw
rNqvhB6k6lxutXgc3EF5SHHg/S4my2f12fWqlfNXfvZwJ1SZDLqyoq3kNQThCea2
MdAtJGWu/spZjhcWzSPyBY9HEljybpDEf4eR4xsjy4B++T2sLfBV7sUhE/DJ0XN4
1VB0QyOfbUFvysjSGP8H+YqQtyTVBC6h60mawtOgvw5uK25OTII1QYrxbZBauNLC
LDJA7tBZ6zbJRdmBv01U/T4hHR3gJxDuxf/L5EP5zH6I/smxpRFW+yz6XYwLSYD8
zzW/Ine6g4WPFQuUHRIJcE4jIKypPO9XCIS9pqqfiaEtzhd2QkNmjuhpog5Yey6h
8qmT3aSi4oi+fkVjpF7UR5FNR1rm1iur+mtJOV8ViJukwZB1Wm5u7vUHLsC017rd
wk+nH4MoAlw0AHU+HgVgKLbgRUgGAU+XxeKTx5RcKQ+kXnWQcH9qeD3lw1Kq/yIl
5JCCjrAtVyn4gFkFKPT6uUeT1lgaG3+CCPBSCZ1CJQw21d3ZwDlwq77Ot6NUCQyL
nNFVSQMmb0sEg5ojbcAaNRRyQ66Jbs+xrhmW+HCevrGaf2Ou5c9V4J8l5BmFc7Sy
RXYE32jY2c7qxkoXGHbh/vToVtdD+zc1VHhHoM/ka+tY4a5gMD7+tjBMydtOvlgL
lxSNwsY5739jG5u6lradcniDufIWt7S9DdRWzMlz+nZlkEBY9+fWspvSPEb5l7mc
1tmPmIs+NTXQCh5168U4MIUDUr8XdEZgueEF1BVoaBZ807a3IyHj1Z66qQJrSHK4
Iea6VqCYWAXlEse/JdIMFsRcpKWu/jQhYtTPSzjoKzI96lPInaQuRUhLi98nRBLb
la7kJCqhAYnmBU8uCVwdEIE/OvbxRD2z2s1pziIxt98K8juqvZdOvs/JtgLW/eLc
4wwxM6GRp+TZiKbP/mMWxo4GeJwhrduJEcmVTpjKDRgPXsWeEfzJybad/JHiJYhm
olx5h12/RfYLrvOYWbJMOTqaD55eF6Lj/2ESOuX1HBWu3l2jXqaJA8s8xE9h5PY7
b4mibixmqMakRGFYjvYq342PZs40zu/R+k3OFfpXX/qkIY/jz3H6RRf6g4cve5ix
okolvN65rf8jfR8vQshz3LumaWqDnPS1mIlGXRafswsY1NgbntRMwR3Ugf4Unm08
sPbt6KTunkjg7v5Dlrm8taU+srUVgeO/fdsyzcIylMsF7PMMN7eC5xjfC0H+61Wa
+Hw8kE5CP9pXGORL4tjuDciE4FaqyH+IUlisS5Va37lx9DM0R2JcOydMdxkMeVan
CdfpRDTQArirxE3krZcWQ3osEy71NTBLq+k7eobApHt0S9FMSVj5HZhv4BTa5ASH
SrsxX/H91E+i5cHezoIGX8g1aY0QIkzXn1794BKEvAhDw0jEmQp+yIjEjAu1mY3E
IMjNzv4XF+M9Yjzl6Fpy03GRn3gZsGM1PUm2/tAOY51pZ856IihIdk12BMFUvIcS
u2fGFk6cHu4URi8SVB2filcs43VsYBhOn7Tk3hPW7yi+vvdevZune+aUzxeSi0Pg
+dghxeOhaIW89+V7tTlobK6+2w5jnNXyG1kPmfUFfIego106oz4uZyxQTB1qtz3a
CP16OCLJoZ9QveW71ImK9Ohow5iCk0HgDdPIwfGu3bpBCQq5PvbVr8nHgSXNsF0k
LT2zslCp/bn+z8kdhAzPR8VW1Xg2JM3fiSzmZVhRws5WYZJ0CICQyYc23w1amzi0
XyZJ7AACWiiSnYmc4F8Xgm3UemT9Hs8lRtwyh2byV7YjgjBBAUWHT217luVO4NL+
xml/NzeoCpyZPFwzJjhDSoflZBz6600TZJ2calOxRi8XPXZ6+po6Eko6fOxM6Rr3
3e7A4Up8OGHF5BY1eSd/91UeuW17B9wR9uxOUOQ85NoIyQBLrTpcbu9mAulWvxOx
CAt7jraiJQzQ72oy+O7fI3YELDbVFuLv1/XcoY4lEWvhkz1J9G29dKManjWUPXzd
s7R8hdfFXAoGbZxB8XEf0JEuoFLVbWfGDmurZAHrsV/cSQFCcsGwjWeZL7JA+TwS
zsN/LGbXfamQWv10L5Fod4saQS9vQ3pNT88iQ9DkU3DL5NmMUnyy+03abmVLDiHY
SxdqnMvBv1Vyya5suq4Nsjmjs4KNtlVzZxFwZZfLp76QZcEWx3c+4lttDLtblsW3
y2f5DVowRtPq0UNpHAJ16QgQsRc+Qo9JqU5Q6YajvcHZNKH7EIJ44SVpAQiuCv1n
C7jMri7xY1/VHgUvBevX5DfEUI96T91IaqmfppAQVVWeZ+DfcoRpe8tpDdTiLBe6
jGgFF4rU0ckIz7F3cH4tPOYw4BO2U9yMRXX5RVsoJmUFaOSgklcbpt7FX5uSRFTK
6yVV7Mn3GtlBL623iJp0I/VbdR7AXXKwvR9Xf4ptW8mHRiSnZYrFr12RjPKqzY1K
StVW1s0LMWSmZqK6EO4jJB2k5lcv5OCgPyy005yihjq8idAGyycabZF/siSTZ/Kx
8/3BEkzvH9KTNAI8Xd7SG2imx8cUssnsySBaWziWEdXRY901+lFFLglO9D0qKhFF
LC2ZNShq++jXfo2ATuKZmDPBuq+6Eb9mqRYF49ZTgSxKOXgQNafcEcovBH/NS3QD
YiwKcup1onR+vRFyUDb7FYh+thjDQtIRR0r45QE0Cy+Du3hZ/iEXBP36L8YYTsgb
d0WcxNjMFOscFgcEhNrRRNgBwyLLT+mbnETt/jvjwSe6P95LOGdi+c7uyADjp4vY
mOFhp8tTDNnQTkjnNUVe3mCrDKIR23mUaSwy2YmDC5ZuGlWmyLnQQ+sGFjB08PfW
5cfycSeTGPMVi5WFCpck9iEXBhNJwOFQ3EyohPVzc6PqNRsjvhPseX3TwYczItU6
KVDQf3lCQd1p/2gIj0jkoDX0zo6VcsCEp/zG3uvIEiA+EjD5U+JZUrv/cX2KWX1n
pO2pWL8XrQo1XALE3UO1x9tW+0WNZ0CrTkB3yoMjSXYop6mTdEcIP4bUch+tQCAs
i7OtzAY98VD7krwJsMexGd4C2w/QohrpKetgc1S8SkZjuTkMMvdveASwNA3KYPql
Rp4lO63srGFwS4U/QCF+B+52grqrlSUTDkBhcRnpEUcln2zKmfTiQkKWdG7mfynI
aztCM2KgsxeKKZcBPCA7uHPAAhFloaleDYhuTjtCCKl9e8zYHpBje1wV1H7wbv6Q
a1EpmBzXQdP9rzMXpO0aVc5x7jcDVf7GawZtlieWw8/qudS70FKlD+6TP9ip4B4T
GBbG/10lIxF/6VRL+Wy4X+kbHGNKO05TbZYzmMqWsBRQU/iur3rBQGgZ0fnWjZul
QjUJfo82gvP6Hm59AOCHUXCYfrjLmvAIY/3u143x1LKrzmn+61MpSYFBZAW4kDYO
Dw9WksdTkyNnhIniOt1RNcsROgbxpJhvJGqqFPrbsC6sdcw0uq9vdkUjLFN3mp3r
hRrgWV3BkjywLTt8vKA9o6UUlVSjG9WQ4PO2LWv/8NbZaLPMAaS04s+lPQmsdEUs
/ybACYUOJQp3OhoGrdAIbb25b4SDDMi2svP1Y44M4lQ1MyLZYtA7lOAgPerWLvhY
x1xBSIEXVs/+Z5Hl3BqYdks14MwLzWHcupdISmUuo+Hhns8n1LOyX2Ng6iPw5mRH
hAQudD3d9KwYB5oCY/bSvepxuv17bdkmJOnhAfkW3cd2EfC+spmI3I1xiCx0bbvv
sar/gM+42HfIG6kiKKy9UVcqnXWJyp7X/GctwPYKe01FgLtwOs64mu8MuyQmi0A1
o7cxsJCyj3YLQ9kvRt0b+Xf/F8S8FRENAb9W92Mj3yKfFdv5YUUuYTAd2RgSYwfd
WmSy/MyIIgUiFFFxTJ/PkRsVsEl6xIxBn52G2YzR9TeSnJfY65pYsDgx16iVwLor
+Z1tBWOzHhRgCr0u1hgV5u3EKTaikU3IP3BQ3872VCwNI5Uu9TqFBJduhzevSIZm
9ZOnOU4uUY5Sj9OpRK1Q+ySZLxsE+Rsb/tPi98Bx+ihOFb54Yg1+WmU9vPOAY/3Z
GXe29QuJ3BAMeDFmRC6Ef0fC5tYbmG9OtOYO5R5v7F+SLMfIMz3nnDTo9dA3g8hK
UEKNBpKx/Ae2qNCNEAWWyWUyCW2dtAyoqLcQ+f4VPfjE84JCL1f5TlSByAaDj1nn
Q1hyZHTkW86pcrO3gRCrd+8k63u+vgZ/deBl5Bmm5ueyI6nPoiZZjp9AkLs2pqaG
j+y7XE9BCqzvVV3KUbwWtFblVBxGRSyGiYNIRIoyLirKNWVadUwL6PYqyiXYiGxR
fTEy5Qp52COn97LZQrikEfBrxse4wyP0JrbdGZQWWrALae+Mjxw6LadZhSrBSPvi
ayxmIlfQKSKkL5tLrvADg0xCi63/gDsoxWdl+ZImKbQMZ4i/ofs3LNFzn2g+vB+o
pWW18Xb8aDVGUASyioflRdfaMwEWxJnqPFM7ErXvzyMxHg2cQV21sJ+elqeUE2qi
DABKi9TTO6hHbVsBNkLqzLezMGAl98/s/WN/JS6g5EQOYJwfAWp/kwoECEiowSZl
olTrpfJLaj7ztIy5PXbxbFIzW5Ey1GgDWVFLO0Y01bU+2iYsmMynIEVQNRw3A28u
RZgQnP3zRSFvBfgh3y5P4C/TxHxIFWjvR8t4I2ga0lqcd9O83PlQbKwEXdaEqmrq
3JUg7hJoz8dhDAtyij6tFKTJARyoqty7eiZ4r/u5X4F2rVRuXvKA1pzpmFmr/GKZ
XuXcg4YBUYqqvwqI7bmcWj18N8xDUKv9wuOnbrcdlXdynQvOee625zEf9WAlPx8P
u4BobJp+pHpoXCvdvMetooVgO7s5E2SQYeYj2s6YHwMJULc/cXUiqebWr5cAwFqc
gwalxpRKmcr5xm+DS17LKKwQu6OhIg5KQLMVS06ZxZnuotfuFTFOPN1B3sbXW5kT
2ZDbM7A5z1fL48isO0gUUs/51zm9AOVH1ZOLiY22RStOuNuoQ3QrlwjN0o5yIrk1
VWg4M1GQ3+ilvVTKLFCUv2xds0D3OI3wL9Zo4rReqWU/ZLw810/hteB2SqcyvgT+
3JTf4b2u21uvHvSDTwuLGpmnMOFOQpm9uxLjUSVs08QLcT3bbjN4YhTWokH+L0x3
iCMA+naIlHv9stx9ZzuakRaGiWbtKwWUxlDbW3QsovhXYODcfwqtlwvhV0NFGjLH
IB71ys50jz5B3+mYGWgkzvez4lSI7vEUZeGoFkovAx9wfQCHJbj1mWymuoWH6psW
xSH8vuPI0HpnNmmS/rVuuWGBFnP+kFRfvXhX7wAK+9+ZH8zOpjv+d8bhEOC41qTI
rGnbjy1X81KRlKNnKv5cuZBoIi35RRuZV4NLujrgdNVx5ZOWjwjCZcOpVu8khasa
QnHTnlNC8bpGqCDlZUPvd9n14rMyNjAcG1OfXQFPvUPNpLY0M3j3bN6CXqSL/na7
inXbb9019EtyTtBD/6endh3/QM/9QUnFy8M+zZEErLvblqkaxi+qtaeIHoe409Wf
wyLxzWMkCvwU3qeqctncnbZKpRnm07F1vtt/o6uufoAy8HllXJKmUIONJ0/3l7vT
t3Zs9IX0zkDnFB0mh/3bGNNRcZoGwpoRTgrG9EwFnbjgSibeT08xUhGxqQPLAysb
LzywS0z/ugEAnJRW0E2eFAMhXtD8BluCPIxFII4xW7GxR5EUmqUjbjf+VQa6E43v
OuKzv4Jl67T8Y+l78k3G6SvJZ21JYCqnuIgMRIdJwQyPMmbR3yn509gwXATGYUi2
NQSRlg3GVZxzGtApSLgly79o7IAk6T1hZ03kzpVvV+hftyL8i3QJjPbdvPfx+1Se
x7b/Axrpw9Sj0wUqyWwA9PR+evsW2EuL381vqmIBWgMNHsi4wU2yLmlVgrHKjn74
PsyOos+yjsMkV6CsAOYGnXKBXYB6G1sO5w54fZgCPM0vHdhggIOnhr2LY6NlIHJT
cHYgy0ByMGTVH8X8zVXKyKi/XdrABwQTnBUplo7mnSXMsFwa2AD8YqBohBmpIBTW
dyGvqJVbUCGF0wLpYbYvNEekaJExFP38v9lqPGubrH5jaUlIe0qGkAqDWU/uLLPH
Lf+d85lqM4roOnEf33671Mp+/scbjyE11VCXD/Z/822eHB35p9a3BBN7Tf/ZZx4n
nBJvqLXz6aaDXIWB/YcIT5Zcl+W6BxYGKTcff/5aGK7ruXaFtmEF3GI85UrFRSYS
tsLG6bKchHfs11hxFVmK6XD9y5OfAL9G6cyGxrC6QWM/gYD9Ne3MaP1FMrssfdf8
ulVBfP+7X1pPu39erttBq/MEREOvgmkIoMPluvl597s8RK5eO5c0tXGVr7p25Tmz
nG9jpQ/ZqnSmrd7YLt8vO6SY62un2ikD9eygOYCFddpwqRnEXGh4hQ93imyU5TGJ
9SvOjNcySfserUZgN1VHYUooliety+BkoRSLq0J7ThR+z+xpiNoegLvBNwJKtbtJ
HeVUZI0NIoj3QUFXy+32w51CNeRI3C1YpPiLO3qTnbzm6QYkxz+Ao30RofXvcIFh
9V+Xo6/ofJncT/+ZyOJCC24r9rJgngBqX4eKShvh+dQI/Gdol4NJ7Kub51nNu4nP
46Wt/SRBehNTg3VjxcDy4SbGpj7zQGd1zHFBvPp58xyszC1gZ/oSe7IFwHWA2BKv
SMULBiUFCoRlIhccz8dpPSzJ2Wu0adgN8rxVgVtjmlLl6eiHl02rsHQO6swslIR3
/XeDPqVPWkssvO/6lAeG9dLc8TzFxBdVv5ZHv1c+0CmuTpDZiVexx7RkBkI5AH49
Dl7BhaeXLbc71WTIxLdVUbSEuSCcYLZ0DH0+UYsg1FJm+02ZhpCqUiO3OpNNBG7o
zo5JGQ0TxeNUaJTOMBmiJ96Ui0Nhz/++jY3pL/ZyRr2nIhYSlGlq+6OfZMCk7xCM
6LC31vZ8cdsdT0/vNm287CCZlbW+Qi29tp1BI4vTlNbMwy69doElTS5od8G4psnP
bBgG75uC0g79JGRk6DofLJQeLEOM8knSeIgUVfY7SrzD2XnIkPR7F4+MdZSMT8AJ
5KIHkgkArfnJJDlo0NG6ixMdyoTRoLFGe4aW9wtJRR9w+ATN33/sioBWtXdXSHBm
m29kFnWUOuR3y4RMXGdu7qOTXv4DNyxTLSmiQy6xANMxfBddTUgCcOgGxJ+EVD72
i974w81JgQXgEUZeLr7wGKSwepH05v7EwqdqD3QHtfzAslDF8FFDzg6DpSawKfnb
q0Ro6MXPQLadm3rUHgCtYheyy3zzgbzO34yTkPR8XtXM5RfNL05C2Z3Pk+lLPTKM
cv+e/Q5VX3+o4TeaWC7PIMXRKnOf5pmYNHO1TMmPkVh0v+rr7uZ4KQ2km5Va2YH9
6uez2JwNQZi+ktySyknhp35ACTa4coY1VPL//4TeiO0+be94uPti1+FoTmGaoyy1
VtPCWB16r0fPzET1F8D7odsPxPblEpN3qYsqnEBdng33PCcC8b/guKGztyahSalE
WWlLi1ef8jCKa1O7VLDW3d51MXgBBj+n9UCuESNVrVK+ufZg23W0KlGfNohgx+j7
l+LlKxzBcx0Tg8HSApoZdlVGRMg+sRsw7eAfyks+usRHgwRApwET78+HEtfc053e
jcA/bNcJMrYVK6ceagb28sN+6fo+IGbJkvDptj65Nd+eV7PTg7nV/cu+1GGEGzYY
gGtrPk/TyiQPlgjmR+PYsrtc3QayBfBWAfV9h0UCA4hktdSe/ImTUyMlkZk3HbnV
0SKdweyMF2iWUtOWO36pfHWX+g/udWuqqDYs1JMBieJKsCCNqdYPBNJlIkw7WG4d
gKhPhZnZjuWcGRZxhsh355xjTT3q9GjRGvmC6To+w6lPjw4fmtF1y98ABU/r9ubV
Dh76oRT9sU5wIiISR1ythGgvCRjwIXD3o5oFrNxc1t15uP34aVvt15/3+AxCKBcq
KZhIm+EFIUMP1HetyalYJQJj9pruX5DKCrhO9eNJsSohdnnzasaGigdcUcyAo/Zw
N/eNMIpCLmvX1SdZQ1zRq8S5+np1kb4nnNojp6KyRSMvMxT4UE6AoLjja2spriEN
phh+BL3r28AsoAS4KPxWFoP23DVUsRmv4cAgBz5+T5acXdFMojbrq4csuDy9/mB5
0qaPrTlTl5u35lpblRW4rdiWZvMR6C/o4eSayDPNNgAVnQJ5QaMl5Vf/YTu0gIPg
tVzU0XVi15WMoJii37DLzhQ0ziQC47V4kRQmabE47q7gx2SnAG69PpICSSmK3OfM
LXOfR4rO8pu6t6SkEarQKqv4haSEcRD9Qve11aAJ8t7OfZQGd1pyq6CIJYJjctro
uD0hsqr/ueKWE/61IWMx8u0/HvXoou6eP6ktmaNZszN3eEH92cl+bkEiHJFcmqeW
GZOm1QMIDyYOPKm0P1VDZIT9Z12VFfHKCx+1xhmetsf4Vrdwa3bEUNkvw0zU/MeG
SX4dNc9eFhiCjhWY/FWg3odN4kkHQVOV5A7EcEsB7U2U2VV7/NwPteP1JrgUfxEZ
na0+DkovvB8JMbRtOh7LICJk/LQesLp+v4eHhGMNCPJCjKMO3V0uSZAtUP7mWz9h
+eWUuyLrxpuzOWQR4x1JBs4L5OB5O2xvW0JK3rYPFbWtzwCIwpzfNh0Pi9j1xWEW
fUf0kMzXELMSJLENLAampzMbdt1zOf19DWH6az2/YJRF/Dsa6ur/turylmOfhbZl
q0F8rHdmPLkYdmq+Kvr/gQ+PJa/WXdwDEDriBkXhxoo2xGHjpGjaT8DXOzb9y9Fb
db0H9sMEeR/hkw1fyt+/ez3jFcDwezJICFVFOo6lHUUCwu18JPK1YXtXR277iUmB
dvlPshkBANsXuO4P2BLdaYhH1w6M90IzRxbrtjQRiQu/VYrjp86E8OfrneYJWovD
EIsKk0HDMlA+/fv0c5dtGi242E0Ruk4BAjvqU+So0JQAD+IuAPlb1443VwMor73F
hUD2TNZBiJO4i96eIG4PrmEkue1Iw+NxMMh1it4xKjL79qfFf3IV7Nlk0weOEgiM
83f8W7XbiXMZmecV9em3vab0Eh1/SKUmid9Tl9e7oFTLQ86wSOUrRxmr9u0RCFAt
v5jJkpNFyZ3PlCVl0EBIOD7Y5lfbmABb7tAz3JVVjeIthN+p4/eFsAKE/D32TW2f
OKn3zFj47U5tT/iRkRf/yULAOD/VZ05ZhcVW7xCjx5yQP8cD6/p84DrIS9fqQ70a
YrIS6RDkCDCZ+lNS4qcYP6OC7Q7VzSjzCbUE0FJdija/QwbimWJ2ZCx6gsFNE92h
gRSXolIDS6WZNdqVadKJVMN8ViMPmRO6aCh3DH34iNDPxgN/KsngFgID7NivLdo/
sEJ1DW9iekagCTbTql49gYGPhQg5SLGOZ+72u1KBQ+Jv8KyJjkQ0KtThNreyi9AF
DYov/beaGzHoqdbvgwW8QE81iduHlo3kqI5WlmbK8AsZqv4WoioL+xMpeTwmVuN8
h0z/I8Nf8Ia9bhfquBVuXu/K0gave5GZXJGkqO+0L611ZO2E2K+j9z/BofTYW9eS
jP+dIrU6T5gNja0fHp08ABo4fpGZxZLGugiXbVuGKdWpamatwdp/+rwHsHtfeWSC
Hwqy+TzP03HNdOO6OQJDnWwsAr01cri0LhuqFMqZqUHB+zx1KFToGhRrcjRnLNcL
YFgnM/Wk3eS5WwbynL+WOT/pFLRAtzUOKV2VTCDyfTYXmxrwsGX+m1516cpyxeME
XD+j4Vm4l61GgMb5pFe2loSKGHAoqvxoD7OEbKb0mnGdlI+2fZVE+j5/9RUJf0Nr
QD37XafcUvCdw0MwoOrwUHnj6Z19mfrd2zP14sUvk+8G7L3ueQNcsPY55eyTDF5E
uvHzLcm32c1EQo1kRZgStL7HMzi4sqn2PDL0ijWBa2JQIugHcnq+iHdsLx/99kRe
qUFB1Lksp/oKPvZiKAMPQ8HBQ4YHk8/040qBSGHxusQfBM0c7YXCU8hxnjlWnMkI
Q128sQYSL7LYfsuRW1Yp5nhJR6QmMkKwCqx/4mvPwvwFR/3gQwXYgwImoAYOOn89
c5DKgcArqPVYNCQYL28kxJb4cP8usp0bDmhZdnWU+PNs6On+IftZAKRm+x2KiZ1H
bklSMTJKlwaB6UY+ta9hjxScRne1WIAzM7WX8/viW4LEDH14YDzUAsxiXweH5QkQ
2NTJd/knXW0Lm9z92tW/+XcoB8hV3p4H/GCAHbnAOPms30b49iqb+1uUxaHczgwR
RAedWrKJAOhaMnpextiDuonqesup/gguZLKIXBuG4uWYWc/xdaMSED+IdC2Tek8X
ekI4JyJklJimQpW8X4CagH9TSAgGO7RQL1wAj4nHMeKR1phmIVjMoSGUzpQvjylk
X264Q7qpSCP8aAxbgSGDO0d+diqjGG+ZUOMObVxchMjhFHTMseIT14NEjCJPyYYy
wni0FPnDrbP6frPHc8RuA70Eglp1S8fa/Gnr4iagO5ilsj6ZNZubRV09w/G88w7V
693PdwXQjkf2umedKSwEXLgba2UqguijqwQujTy7Fc/nRCLkuy+ZaBSnitBJZ310
Ulcwvbv/VzSK6i04+dPoi5liU6g6cY0Yvd+Fcw/sz7RqxUmNKlG3GotgvsC/LJ8F
KV8osEq0ge/ft7jyrk780YpHukqOnu/63gz98GGhQ3Lfz8EfANtIvlv2dfrl+wpS
EjXQDQDAKVnd+xLbK8S0L548b/ey1wvHpukCvorCTDOHCq59eKn1nEFI7+chLjmX
TfT2Ece2C2iJlNNCkWwXYS1kpMnWT2+7O3fbmYKIrDTL80dbbDiMbk0huxKp8NuF
J36vmbsoMJda4QqOyGrruve5FOSuataDVxoPXJZPUmhKYM3pKjfY/k4ejs2lnrh5
dzM68z5RlbCJnugOm2xp6Rka/WOLIyeanNv/JbDniqtggzCX9t+yBhkyhbJHLGXa
xOhqYJvYE2TSfIP94Ft4oP8SCV+iZWCy05bnXUSPcf0QV5w2rgLX7EEWPSEe/8zs
vYRew0vzXPA1Qpmgstq9MV0Guk3imuOdbKci3WpN53Y/r4CUEUkjcKZmbtuSYCOo
Rd7wL0+6+0UV4AFLRC/13qKwNo+YiOz49MXEtHBGqAvZpOkD5FP8KJBmrTK1WXcz
wwFlzMGQjpWKRy25w3P905i1ASJWZKBhSXy8ZneMr51WGCwF7xNxx8+VSgK2zxaE
L1cZAViiU4gqU0UnapxVEd09tplq2UPFVbRXFjrKiLS8xDv2jX9U256EHR7Alis/
a8idHItIdrdbBwHv/Ab0DwWS/NMy9ueJ2nlHHZLxPtkcslMRL6f8hJO89tHdgbBr
QM3d2IyuBt5cxAAzaBReWSgZiyXIwPuv7Ppj9ZalSihLXFFdeX6QWmURF+PIyWiS
aEFndQikx9YWDxEszQUpE8RYa/7FGXjRbhcufg/Rws0abKPURLJdr1JNEXf+OYAB
tY/7cRGqmjnybDTIgIkSfJzIkTuEQJTwPoDtUxqX8izwjf4/W/7RH0g3SOLYwITU
MKOBvZsXUAN2JWa1WTZuOI6p80kkN7aNon8bnpbvCDp993TUtgDWlVASCqNbxrX8
tC7DfOGKNjv1UbJJEt+uLH+qKybptvB2vZqocL/8sTvNSLgLWqXtmONMnbg21vtU
SoYrA7GPl8o2AyfTkDKcSp71pwdKHPhUIrzfOYcTcul6A9b2nRuwHTOcmtxUcP9w
udfYljd6hlZMt8GHFKSOnRCVR9TOiergQDet7e/3TeIfQnVK1yN2g9rBq5jwLvm0
TWztN+rdWc0gFDYBgWhya+zOP8RKCdhuVv5WkeBVRyBv1+UBGdW3Jk3aEUTq/b/A
B5ASShvAZypFI4dCc6BQ4f6VrubSLXkISMY06TOYxF0V2e+PDQ2+QdxPUmGiTC7A
q5NyDBtPUDrG2hGAXaRWwObobErJmguo+6F0iFYaaDpGrrft9pQoH9VJ3EDBPgwW
p2XKCzdmicvXOlrQPGpUh15FPkDqcA6EdhcQhesZCgCJNZTaQ2SkVhfEbJob9sHa
3MWDilnxTtmA8cvwBAesmlukeG7RIB4sLgFceG9ARxaLW7l8H8R/vASwxPj+Xwh8
Cpp4CM2DlE3E5DE6FXN6wHjeyg+Zyb5rkj38e2zFXAdAB1OGiABb8cqs1WMTFpo7
2f2hbZXCIXGaHazX8yDzIT5BhBqDW0qcFm74s+Eqf0gWVUBEbT11/eWtqx5OIAbq
pOpSJ0YLWnPR7jktQr30UuMyRavgJISycbPB8yYMhUO863Mg80VOAvAIzVvHaJZc
3TnIb2clM94DCwlcTX8DaBrOe5T8JscLZJYyWf8BWDyORUmOoDSvD7jeiN7Rmvkf
UIyemhqu/AvWsYwv7mf0JwcR+ekS3blTBN7hSbpLB4wgbDt7LMCSAo5DLoRkrcGQ
q6cecPK10XGSXzqJTD9IjQfQ6BMHSeW6w+SIEbg3CsBgyUNgm4erJG8DE1bVOAJT
x5YK/owoKQTbxfDB1IWaBaMxAWP8g+aeLqIBnCXxXJsaVBi43sBt3xryKsmPfzGE
9ihuWPC2bHiU1qPtb7lTUqtDW/er+txTXrhmcpWFAiC8vnUm3KHMFnZmctsKnI/O
vpZOpx40OuXoGwmXo3ZyMpdTKLlHIKYYbt0oq72fXCOFWB5ROvmgfggNmwdaz2L/
AwQpJZSlI2MvdhRR95WkVn7NJXIpk2FJlbc1o3S7EV34PfWDYi6YK/8Bu4kZwyei
i0FaAwfSmNwd+/GbOQUDwKVJS24CVkQRb/r2o1mzHzNsJzW3MprGIb6viElzNpHO
DOE9zDLrN6BtMyA/OHeBij7M6edw32LYH3IELOJxt+yy8JEHmKo7Gy+gd2YW07h4
WB8riYBRaN4i+zK4ezc/mzCWxlm6p5V2qJWbmYaI9N7lMBFvTFlPTmYuAMH3rDku
WZLAEaUpCUbe1R7O+FPgvgU28Rw6fhLBuFtFAG0Gh/vw+vIltjRf6VlEpfhO0qnF
cIF6m4pn5Ljjxwl66o1mQX8y2y0tOUuIy56Af/+7oDgCKwR3GT8WFXOM6XpcnAw9
alX3jkrTxuxWQ2tUaCaCdd0oOehy2WkLLhBCriqoLDJ++Nd3wMI1Nxd8pmJpabq4
MMY5upqldnavGSanjOaz5QYuNuM7OfYDbdQiVAuXuye0NaObOH38r+DbrpigV4mQ
1q2o6GNzrYg/Siqlijim7+cZXXeLRzgdAs82vzZa5zCSXB8m7CqJ+lnFl3eBr03s
kxyQ+GR9EjsVd0HJNEUint8HZtd8EPrHSTVtcEpadcnzfCu6L0SzcrA3QUKI+w6A
xypK0i67gciCMsDGuXmpGxDB2f/ZhYGeYpp/5TYKGITxM+c2vI3bVF8+exW1ZWHf
4RGAU32lkpGD+7hYxxQZe42JwBqERDr+PJRDy7FDZyEz+kfbdmXqR34a1DD4kNuR
eCjUX1XUy6A2RTHc+8SQtzaxubMB6vjGAONBCsDVSMmEm2jCLW7amTUbp5/WS9ug
3J4bJENo+WzmLzrYI8UAnhnnJwPz67Zaqb6i224pwIWCq7giFJpDaF8IG9r+RvNk
caCQVhh/3hyUFxyxBaQ9Yc8LrKz6WPqh2PNTO9xAOdgFJ/yT/t5mb2Vf3oB+OjOm
x4X9qwJqdUgcMpfqV+L7GNJwJNVsJ7oPVTt1+t7JILt58yIvSQY2xElM+FShyly5
xRCsIPTM25Yt4cTMAp9VoxYgN/ce7jQiz1yJlj18te6g8K9+xJnesna1lNWE/edG
5X4CEy2D77U8vOrdAD4An4LYNlqWCY8GdIN1mYhJlWilr9ENsFt+D6kStMqkCeYd
j/OXzd8Kg4GnKlSiag6MNTnfoMMkZev2aZsY55T9C1RF6FfNSKI7gri/UiNJWdPJ
DzUlESJsu2vTTqiqRS2nAv4u0BtWRexRqXfZj++xCXQQScLnN0935Q5z28Arndrl
aa2/jIdA2d0nnSIQOab1+BedsevXb8yHVY6VJbyN89yn1req+t3Y2oXrHjkCDNhb
s3BGCgGSA8dYXzOvOOQB0umKzvpRhBOrEV889uGaGuNcO3yvcN1R9ZwTAPcf2nX9
5mSPGqOL/5btBt5LNJZIlhodmuIMnBo6FS4kHL5QGgO/fRyKQnUioZ1YawyWOD2u
Ntpw+vkazdiBA0gebYWuI6K7BAbqn/w33Vm0dTIHfoTltk98ZTfhwK8Rxpuyooh/
M6RSC76Z9bmsvXbHOQTTYFrvmoA2+msg0rWOX12q8Tqa5cRo/9I0U7pvB77Iwmu1
et1aGYYT+/wQoEP3B/zbDEWJXpbNgS31zTNwcPEBvLDhZ08Df2rF96TRl9RNwaME
b/KAaWmTmBb9r6mScAYZTP/KfRYZ8LNM/apDkWDS5PorALI0xX87lTMLoCJuk9xg
eP1FAFVknj1dAzmE2s7Za/o0j79WENy/AegQIN05PunodnHT4m+LH8KdBsZmH/SC
igwVuRQBKaKRq4GhnF5ryOq+rRtUbfj+G1mCLF8McHW3TPFjnGio/oov1UXSeZdl
+QytDwCG44r1VO4iCLaeIIqv47liLJH6hefsumOTZbiwDWe9G+jEbq9+iYPXVcbw
+cOisiio7TBKX8AaZtIkIOgF3ZAvY6UEjc0WEC3dP43OirNpqlywtCDzSFUH3jur
rpGTJGgjA7LJ51huGDvDhl2Kxi3/EOaFJEsvFRkikd6AmDCK8TyCiQznyNeq2/AH
TOvC/C9aAO4d6v8StiG/XgNGRREqMghChvojUOJPToPtGakTute33ojkAkS+I9l4
xxIGeCCOhPEnhLulL+dFVWz+zBgdLq8DTwGLdzwgXuZPfIL//KDT2SMl4pJkMk2H
V0YVjq3PXvSIdBwo3a069DGoJ3dcYE4CWyZH4bfrGo9PQozkAC0fGOB1sS/EwHIb
vq3LIC+C0xLsToAitVkFHDb6bDNaugn0OAIhkNdCT+xJuSbgFJg7Kj/QJkXxVaUf
Lv/xtg77mXAd9KGOoTsDklQFN7DDfy49Z3PTYQ+SukKlNHIXQBA0CpMlCwU07QRQ
junp4eACsjEEl4tdsL3BHmLCepn6DHIvpajG98Di7Y8O066iieZycDchTTVEUmTl
pQw3QLH1/LOWq6PX1CS9sCGzyXK65tE7k/JkEdcXJUFKFaObfF5aywPzGLpIet2O
UkXcKD2f8T7aXL70Nj5pf4OpRqxtMdQizBqp1VkgKcQP5Ieruj1Mp4p1uRsfzaui
ooyaneh87ny4FbADV4SCo9Wahlum269yYk7hMSmkVChIR34SGd8sq4uxl7MQ4PQQ
5TvEUn1SLcuyLnNIBPB8pwpFTTRAjeWCmAw15TmBZ8juRBEZsDv62nu1WS4Hbe6z
FUoxv7RASHzMOfK9m0QsKLfK9QfDdJQIieivQGl/c2TOsq6WVTnt1pijzWq81c+t
clVx41JnCt3BQg/t5q1zb6oMf/FjfA0dLisGQ2VqvmvLjN11mBDumZc4IuVpiInT
jTWSosBn4H4KAr9pjtT3k8kJJCOOMu/zBo7t0VDk/1yrH/ldK0O1Rf+/QwOL4jNV
k5eLrooxiCn7Gj1aJE9oPE/9U8vuVBqUiyc2Jjg4Wx/FGdiOT0fnecFPkbn69fEW
uYrOZ4ewA0ccX7GSXZSGWyIDk28KykdhUCmgwznrJVBUjgylL1JQnzR/WFXflr80
vTjwSzjbK00f305DxUA5wkmH/QzYRDGwYcoCaCnshDNNSz0m+EWqtGmOC7JqWXyq
Q9MVX6IVhtFfavmNs5ILqZKikNeIGW99EK8QfkPQ6Qg7vWpy2gDvPSXhGnpTwwGm
Z1EHhLTk/hhJiFQEYYjVsSjExy9tInIH6OHqI3m8M2RwI4GBeZX41Ubc74M4GFkw
Qkrig5SboVCH3/VlI/XQbO7txOZcs5fE19drQ7/dqRfBc5BxpdDNEIhZysJX8C5J
hpsqxMid/EllbA/yj+tAHnzA470WjBkvwkS4PsLiPkIXTsbFdX6mzLNApeindTgC
IS2fUtTCQgGe2xncwM/S5tcGYaak7YP9Cpm4diRYE0oe3AfWZljz12zPUljXTweX
YpzDgDzQ8fBTWZnW1CLwLCaP1VkBXwVQRX3xdEJ0L6iN9j/3A/jN0MbVJP5wgr35
wmOlAFO4B44EllXaDX5Rgoo01YOIp8vKgKVmzaCsi9nVWAwPfwpOp/vZlvOfDb9C
XpXck9h637tAC11fgKdDFeq6gFqnIqsGDpwiZnYehdWgHB+yn7/njWSLMcyvNxA5
8nDOEhbGOYoSDspLCTJhM5NIBkAxd5aYGMreG982COISuxH4FKBB6+ExFzzH1fZe
yMsczu/Aqn5AduUndhUVA0ZXRRKXX96pvzkG6wegAWwGMs6GrPKzQ6NhnTt9qQp7
O6lRu4K/o/Z8o0dFz9p78xNBT/BpFmbm7dlB0HutFZb62GykmRxO0qHbdN8Ch5RT
B1AZ3lLNdeO+HM0QM75Hp/eVy2RQAhhRi5a8a+hSsOJyz55C/3dN4SCvITZDBTP9
5q91iuCFyPYjEhUEsv3asQQ3RvMoef6vutcaNNEdPtS0hS7Dnd0VCruDtpmo8ZGw
ymCho2teP6ijwiaOtXxrzYxsFMLEdM5eyWBniQ2Hq/pYQvMH4PhPa8yfc8VH2QZd
wKQzZ30m6+Kvwf82jbs3pBdf6dPzIj+d3fnHQRgsbqO3Q3Afpl9n2PGehFAbqnEB
3hw2q8z5/zwFgczDh40c3a28vBJdo9f6d+jq3/s91V7qRnzs3+Oyohw8G8oPl7fG
`protect END_PROTECTED
