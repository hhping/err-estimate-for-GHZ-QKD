`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adJICAYwUpYm+Cr5WROxnQYdbH1aMXYOziiCqHdt2AxrMkVzCynjY2GZkv1C4ik+
SSA1j0ThsM6iwLjI0ch69gRYV6MNatibDdjKCL3uoORFlFU3I0GwFOlAvEiu2xuI
UPaYM5DstQqJ8DNturyI1zKteyyFaGjnGfCSJA77zok/9PTmzMtsNs3UW9UJOmfe
8OJq663L8kKtM/eSS8/bOpzkCw8inOD0qq8q0mpzB/4h6YFgCAvI9YiU5SLaPb8Y
q0lYyUZ+SQ3S3+WjOG8VxkchVIYEOBf3FbVmoU0F5brsu86efQfn36TnVWc8HpaQ
G/7C7mj3QtBjR6MdaWTBlcbgGKJ+VR3K4A1/xGisHvC6UpYdM0861rxNuOhpwfLt
+j9nEA+hStNzKRFZJgLAWa902xIzq68yMqYGKZs2A/o1xe+mGGP1RmHwPo7J6AHB
kCQegK7huupcZrqFfGOW02fgIeUSYQPN0AxtrOniNPlHGLOOPcdNjQqm3NYgb8Kj
KcHLAUE0GBj3y4MXl8rNjpLxoFaDl7WHzjm7SLRYH4HloMbjuZpdbdBM5l4pwBcf
erIXMet12cZvlqm+E/FMgy745lv0xSz6pdbl0HM1uMacz1U4dSj7uzfpUJskrHtl
6YE68sVhla3t/emGz94DQeNVzdRhNA2o9sU6CGdhpZNa/St/zD//777t+I0lzFWc
ONm8Ihnc0LV7rIhcHaCZqXiNZrrlcmvsLtn0NeI0EJj0mRDE2dSOEca8725pPyPk
JQvcx9jBpTp3uH8ddpMPUGJpTHeL6fUbpz8wUttYyng=
`protect END_PROTECTED
