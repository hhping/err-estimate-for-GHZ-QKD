`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLtg5OSNoSIQUHimezI4Lf+Rs5DGjZ+TQCZ37KiHKryxlkS0f5YA8dkufa/qNiUY
2Ed4l6PfNfK75NxT0AcQoSj/zbaaqkfNLk9HC4D8swDhSKsTVdVf2qFTHZxoYzF2
jg30kxY5rdDg/NCYwQXxOoL0I+Myeu0ueSlyroESrQZXye2ofSL50Z+cHhxpyLKf
6eytMqAmaWUhH8oTyzCbCpqLNPieLaqqHPZlSbEPEENWnMoBZ0hnIonNY/aaPS6U
COuuMe+2jwf0nzep2pFBjGGEKucPp9jPuXelKzk0Zez3+73pQlj8E747jdc3YDNv
DmgWOFKJdECtJQVBD8XXCL96skH8+1H1yk0Zs/PS6m/aKho0EHQb6FWMJEowGH8p
/7m0TOkUyxjxZuZ5mAL1SgYdcqMkEvDJXC0PoCysAsoyX4eQbb0ZadfD9r0Iquel
qyILWjSWJsblaZmbDNYh1jn7bL0Q9QST1UoXo5Wkp+0PIXgFP6q2VmT+J7dWwlQ9
dlqfgWboYsxSChSg4J7fZwA0oeWob3eaHFvK+cefR5vnt3XxzY6yULRD+s8+6sg/
1E9Tc797/xryeQ4xKIIrftWznIA5zGLSrz8emKtLgEzlN9KlV/UPCBzWYHZ6FCUu
BINoVS8afDG+x6Xd3CISU9q4to4uq5uEIYwDAYz5IDyADuAJKT0spCd7Na+elIyC
hW9/zWrnm0mXaWZZdSmulLgKzrZK9Zapq6+HKV3iSJ4Lkt1vN4mqeqxPddN4gLTB
HKhJOXR+RKb7kYx0hq+aA/BzM98VQRLYLPRyLV9sEDT7qmKjSUY9W/OLOUkEluZW
0wLv660gknz2VNi8shAZEySIRVml6964n733Slfrcelc/A6gTTJ+XJwfd4ZpDgFE
tKvjfc5HURPv4CgQrRFWQcA+rTxglT4bfatwOzjCisnECErd3LmnHDS6AaXuO6v3
W2ED2NRpGMEMcX164sBL8T1Tj74+B4bJ/YfDboVOfN+rvvL4CaS4OPpiBuOKpoOi
gmzXFtzfE+EiHUS7tA61mYfZCHQt6c2LVurNjf6RoTNEy4FArltWaqtDUKD++ONS
rcCK5QsCnrC1xGAN7OgMKAAnbPY7XGzDyO1Xp8+H02dYomGVDhFNJBFy35PiDY3N
HtIlePd2kdP56MXf1pU8jSmsJjI6cGgYJuUdOjbGbcvPb1X3UT+bB/lOsysQY0sR
dCFr763pzW1QJ1p+5qY+dcXi+dbQnsKr5RKKno1R6wtbcUwmspDiNy0FktlgnK2/
y3FI9k1hNR74BcNrLFtufqRh6dolsSBlt9+iU+zPCK/daWwNsMeLgCGwtEs4RYds
tTz4X43Sh1o//gV5sTVa4gKGncy1pgfp+f9rgYwK/fjmK74REuGK+aET/ccl2HOU
/BTJULIsjjKxfkVwhF7fSdO9vTmT59ebpjMJJ+7/eipl35+axLaOOaTXt5fJwF2w
X6oQiXyxEwFF2R+lJ1znGwQQVzs4Ld6vvBlNwjm530JilUOgzyTlRHylGUlFEXTl
tTTpwyraBMWTXbn1I5sGGM0dUfNNO0tOuzuvHhRLCQH0sJrYG6B/V/ERtA4XlzXg
W3p2U1/Y1mwPoL7wTrFTFdTcY7VLB7NEycplHeGWxenYyt27jMYhrGT2rT2Lv/VS
Sd8X33opFWKByXa5NN1DMPWHJ/6vgvZPgMdzfyeZz8nT6Xlw66tLy6s5YyTt2vwA
PbnKADRT0M4Le+Yt62LZjkMVSrlNUSAiuchJPpBuAF4rBqqI5x1yJClfQrbeuAXb
Vgkgbl0bERgMDfIJjPDLyO8X+FXOPlpHG2iVDyfTyJ7COZmSYy0JHqK7gdN7D+5t
pNtQQssejYt/LkwNyQjggo4CLbfC/zAvT31GLvR3yUq49ytePsF+66thQLsrKcGj
PjnqK8NxLYL08dtj6I+4tGlG1qbSnnIJsIKZ/FOqS3a78DQeYgtt73lI7n6h4uoK
pxcSTO0VHYt7I6Sd9ufRVBaOe0bj0awGGFQf6hpP9uZslYMVliikfXvFrsnlBz68
fWh3j1YsQOTfb31+ghKrmiP66F9OzVAAuvL3mJYUsirP0L54NYhd+oYoxlXuO7cH
dI7u3mfKHccU1puUKzJO/2D0/xXODcqlYNMY+X72NbDqkMAgFFVh+OlbX9oiqBhv
z1F8lb4lHDSTN02nDLYTvkcqqrtY6yzon9kaC3XGcrf++MNrfYibE1pLP6E2/Q5y
1nZHHuq3IJD9h6m8ncad8WqfxMFMQruLFiWlBFYwnn8MO/76cLnb8lU7+E2Z7k9O
huEVxQwm8oKNJyLK35mqGi+n8YPylyY6OXXLT5dM+YjLkab0sEWi5MllgR+N7ztH
80qQsfLJnGZO5qJhCPdL1ltkCekm7HsiRYiOr4ZzGOsPkeLg1RHTlcSKlq3X3fTn
COoRmyowpADoa5SrvvArVg7Ct/8SIQUwe2h/hwiP73cKhs4DZjAIUHNrjdr/fwV/
LleK/1+aUr5yeM/vccMGlH87ctfh5BnJYGT6ONKgMYJYNBDljTH92Dr/6CAYdnTD
GAsxqNlU6GsDB00aYcahIDg1l+eo/SznBzO5KzNFvyEqfe+LQ0i8OSvFODnNgKbF
x51hrxkyw7gBwOodbFFTBTjtvCwqsKoiTiSzMu0Gq8RO33ZTU620RdrZtdepA+qV
HrFvi6OsQiV0aQ3LN0z7fiYh/soQofWOpApVpHC0q+rPj5isFoZYGPWZ+jpu9PEx
X2+nIc8cyk81E83168qtMUVy9REfDdJxFEBUqAHNThoGLOxMM6z42vQMLKs5iOI9
ooj0mQZbBl5lPO6qzNB6GlR1C+/btdql4EfXiXiQMEPKjLOPeQ/fa9y5Y8R5CIUg
gDHP9dDbK9Q6Ae/BxMLFz6dyeZMAVAAdfoWh7nUDfvyYQlcrzNDTqZGQ9Ip8tIow
gOYOqMzhf+VTPgYz0PPJk9Ck/fPAcTjwueU7UObn86wholrhiBz6ow6AInw7CLY/
pGNfckqIiNBHJI+HaH5W0FfamxsNQpAhEDwHMhUV7onKXVfpuMa98sf76j9AGWxn
RXW++qV74DSbsoUehpPSt/WZ9Vb5uebjMlWs5IWUoYVebVcH+v/5jgtRrtjCJOc6
/uvH1lKya7PmnZpWaTKqrL3g/s3C14zDKnduM0+vEy6ufiOsvuW8o7z2OiIH0HJ2
8BqhcYe+l9PybmOo+vUkkpzxuvX04NyWQXjNvL0kZEqMZ1NAJE2SpQn44lZHS2bO
nk4u63lC7GaziiEENS8dEtrx4pGUgOKi6KQ3h5Acoda3NmBUzC5QwQ3yRBHf+CYW
k7qUK+pRnN/1AyNzA0EHZiGQ0G6P+R3gFCKAXUgT/cASQm9JAIfmSgcbL2PYDXf3
mMrTLqWTeShmf+mAp3qrQmoN2PqJTL1Io0D/6gaIEsCRMvEbIXrF35x9chh70A0R
Mw/G2M6wupngc4li0LbozGjo19y7jHFQFWw3klOBbBLD85Vx311+dkM5hd/eiLdk
5pfM4MWOp2PbfddEPfm+zLIJI1wAudfWXF3O+2T0eQRz2HdUi6ApFBzthsrFQDn6
oLOODK1mBLDRi37BAVPmC6XMUAhXEeOL+fHpFQtFg1cPBKbde5NyKxeCmgr2M/UI
f/kT1Vu+J987Ig/OYHFlRivT5EWvwgD0l0wbRq/ftxLKNwcLI5/qFKq+A80vhw34
fwjJTukRQbQI0ei7mZfi1nMJUpfNU0YJvS5f9oq+nD2KDoq32Vm4kzMEYsXiUFaX
YviaaZHNIhkIYHfHb2lo6DTLtYnw/8VcAUrkld4flzM7hPNohw8oOa5EBqReUGJf
MgM/7G+M97Wjj2MWF/PnNR+rFK/imnAZCjIv+rgNVf69rbO55EaCrSWaBnmQwWcG
370e1yRc/Rzw6p0/Lty4G8+xvkeSc5OGRwxZyxg8XoesyphwuwSxd1Uq9TrUkACt
I5hYfVHHXpOOZMKyvM3fvvY/gbeuHNgnvyx29wBTMuhg5zltGcz7PCYfcjY9Wcwe
rEs3JCv0Z3OfioK9XpnIiITEkShyMLQG4VeOs9JqmK5+DYo7oEiXNFK9BgcNfYLX
BzVa80fuW+5vvZt0UWUvkQWlJofZQNNDDEmy4UY7pAG8KwlD52Pov094JeNnjNt7
5kXy/dfoIxFStIzPfc8g3oqzJrwUlSlBoml2CZqGiS4zIfz/ZXvCioXRiopl+zUb
Qb+ckBUEcWAgrjH4s2avZT/gHUNEy0lnkC9v3kH4puP6le/LXPWinx9qnAZQLXAK
jxdIMYD45ebhYuiVIwXaNQQINEZ74TRtZ0MxIDwU13hT0zm6ME6cRxuxp2DNS7OV
yNorsmhSa5PhLhOEwtP6L+gsQ1dj4Pts20BZaW0q7164rEttlmhfdb4R5WBe6FlY
93kQVDYL/e5fxK8flNi78aHgCVk5J4x5YKZ5u1pVSfl6pIAesfSKYKWIboFFYea7
TQHmlWfhI/Ki3vDurs2txn/Jm3jDt++jPI5cikIeHA1mlKHJpQ09A3pss4wFLMLh
yXA9cU90BigmOpim1D4+JvHhcBdM4gM71PDad6qYJkJAxxT4Pm0V3stpHw24T1UX
Tayt1ZvYk1QPyrReS35dYRtD2BMeWLujgjP6zAAuuFZ9LnyQJbBfWwlGRixnbxoh
MRr212y0DQicjj5lLQM+gltpUEAbB8UNrqBs3JrsAX05RT4jX/2B+ghlJLUrpZcg
dYwN1VIpUyEHL1pSprGq1FL6c0+r0f39Y1J++Bi3LBxaaZf+QsylFb0c+xkPuNUK
Z3ha2wnsqcsEWmaIlstyLgnsSJlqyNwaHehZYYCZihy7xfUhZ5fIoaP9yadxvwFs
/VcZnZaKJVQFS9VX5X6neQMUBrWUJBF0HJxCggbmtox6WWHSPP/bHqjZabsIRg7q
7nHY5XSWovbDzZbKUR2v6Bb3HE8YMj/spJ87K8ArYgrxZjcYbK8nQ/jC98baW+7Y
RSV4Zq/jzX09BbhtTTjavCz00sRkHI6itoV9G9rotqwcufLKg24S+hYTEF9hA9G/
O8rtMPneC/6jr4Gaxs/FAE8k82xVW9R8wNfkFxv+dQWaavHKnMAP7HfpakAle/HL
iOb20ESXBECC1L/22mIVCTiQGtB+di9UpEq0cxSu2y/PihKDnL+OUShkl4pN9Lku
LkJWCrc5SC7JFtm3gROdm+WecjxtHGsZwE9W+quS+Xqbny/P27orVrVEFa9dguBk
eiAcg4QOtPMLwnYtjyPcKN1mO05Qa2p3kkX0r8ilTVbgPGr7s4TDJiR13E2Ew4hB
8th6EXpYlWNfX5FXRvwCvzjbC5WNr1LGrgbkXpjaK1b3bsN52MWpAmH4BgrbfBmV
76uAw1hIxHa/NzT5qftXwpCRU8Z9gT4C/5hMDdv81vKYRhE0Wgn8LrhHoyq4fsmd
fAIrO04z2vLWbMWlX4kdkLymMnqMQmZkuqefRoqhX+D9tG2GdKmpSnP+reiM9W3s
d2phx4j4o5ZfeHj+otSybJQ66UMwQIZGs1RHE5ij7zjxFYKsnbBdwmuQ8EXxXOQ3
7ceu9Fu4U6of2avRxy/krd3M3K1ty8wDFlrdPyfF++rDvTrdFQmRSqdH7v/zsQ4w
F/U204pxRG3w9qs1y5EoSvOpl9HLh8MHXqRORIElG9jqeR/wkQHygjQu2qyQzzqM
DYOf9yHIzxhl1ynKoekDSUxAjI560Wu/Kh7La1UMpW0AT8hvVv1qXztyf4mqtwgX
3Qa0UqOfwJY5HkGyPlGDue1ibTjMkgw5tscdcmSxctqZmZUKqOO15lOYTGibhDJY
o1s67ppUV4ShRLWTQswp+oSZ/DSmMZxaHIpy7pHF8BVVI+y5Cmas4Ex8OnqXMXIT
8DoH8ZDrZrmCQ1E/ZTryhGPp4Q5sxq4kn5eoWjsEGKRpAoXO+BlxMBvPinLiKVo6
MJmUmd/QbsUisOzMgHE77RxiUmGK+TcSlAbl8I/24gNHD7bqzFvTJ7Ce0MzdjyQE
VQwKOMDAQ7NlGasMrthRSSoDGe295wL/k/yhF1OnTOxQfmtRBqBJpt7jwUmFsjvp
dxfzu3rdTkRwxYrL07wmaH154cqFkPMjqkg914DMPm0A3rJiNzFWeUCYZEsAWYDh
e/NHzzzJZB/Mx2cq/ac1lwDx8JAo5yzpVzwRdWnBk3EfjNYBfGTkZO01dwVJE47R
hXjEuBt8qFKLK+PVav5+vuMHOdQ2LA7WEWnwi1dCcN7zEG4v1+XYrMG3iZibHyPf
PAdsP/yGVVpEBWNW2QT/pjBXdjy0NNBZInEAulAAQIFN+rrkhZdx0hBfHWClqsFC
yywboNI/Fp2kwnpXzhe/1W73y70evXCgZ3Q0eZ1Q8e/BXz+i/rl5mF3LmZ0zVgGH
lfAqvAACLnPiKoHXEINUjv76WIN9ZgIMU9UnGZWWpZ3uENZggvEiZYEBp9eQJ6dS
GYla4D+kBQrMjWhlM2+UFI5+S7rWj4FbMVXQjuWfeXGLgzemR18IryNaBUQihy20
gyCDnFsM0SAmr74ITO5M0yf6CHfPpwD/r5J37+TvbOs2UfpaJbu1UuiVEv2iGXOA
P4mX3aIeqxZN+d0A1swlomm7sdCL+lokhNoFB760T8Aa54QC+luM5sbAxA7Wzn6o
odyu/+QU/ARjSrfKOIFXwvbI0RiAG1KqFg9eMvR6BXpJ/LFdKWAwZRKnVJVp8nc5
jxGsqYP12vGMCPzectDkeK2TUiJ2wKo/bvhQjZIlFJnQGOQo77FTmvPOGEK8T+/z
mitxVHbPzT82mtyf0kEWe3otSTcW//UdHTTQsBhlJWZfC1MwCeMHtBhiuT4n4URF
5AtNEVeyObSTtoFFmABHMwcqbHf8q3+CKxVZIgsV1qmnvvaROmOhpODP1Z5+bhfd
iZ6YsHV/4fqZUMnwGpuX4fZ7T7GcQwclDimEAA9Io4OmSw5Ag4G2khmoV+4BaCPh
HXvLVvLewjctJ7fY0yaRHSEZzx0MV1czYDiO9Z1MCIKTMDO/P74tvhe0sUYgfVbb
BW7fMQpG16MDQnSscHw9Dn3Rn/YOUMFaKcRs2OJfofrfFUvJW+FeKnh/XZqYCvMr
UbUmEU8I/14pVjvudag+Z6h9tT1a1Z5sbi1j6JyIUQB5YvAsrbqmeFb52cGsTo88
dDCeE7AvIZL2wv3eo9Zf92d0MZ3xn9lk5kv3tq9T0sSGMI5wesbmTZQ4ELPl0F2J
Xc/8PUJ1Hiiql19wVestijprsg0E2dumZpJkBR+/XxFTmL5JQrkRvt5cxjHHkIBL
jnwiPWh2AeTPxjjuCv8+aCI+cCP+Wf1gJkTR0OTuBcefV1k9iEgSbLxhKLIqnOlv
J5GTskOsFnCVSjvB3QqQs/DwbIx7GOzarsLxrT+drgZc/ajD7BSJsZMId4OW/iFr
mar+hdIsihJIQy8UZmAT3D38pnttheK/a2muZVhPsZoSjKh5azBNKb/R+OHGcHeT
XcjfZXTzDRVheIsqevQFZoHUaGOIya+eBQaR/zaa+gJ+7Lwh+LRNdFdlU+dP/3Ml
sb3YxERY+rzHAJP3ZQxywcguRHcY4h5GB3c2IQlbbW86FSBPPvjt4gCJZsqopyWF
rKvRTwfgLIFyn0kEcPN+GyztsmKIQzU/CWeQVBv/qK0SFHUGwSV7NGDelv7W63In
zYIe7CknuNfJiwhMeJoL938J1BGlqNcT8TYV5OXjZVivwdpmgveNfbZG7kj2U5fe
gQ5FnO1PVpwU8rE0f6rJdrnaTOTUngNowS1QuK5VH4hdQI6X683duZD64iUwTNpE
DK2f+R1OqTmsrMSzUcgCUXbh+Urtlj7DGqFnt+7w7jgKgUBcBfUPJOQIZYqRYa1b
Ecl9XqU6kVoJlTTlvvpYjHfjc8sSpSSwQAK+AqRulGrAentMz0fWVY3x7hgi4lHW
NjdFZ/LQWi0Rnz6oDk1xWbdPlElPEJRCVL65q7nwpVOk7gc36zr6CFyv+PuKhGMQ
`protect END_PROTECTED
