`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yM1lnGAEYi1TZN/lWHfUVGY2pBI6l44OqkbVRExKx46pW9nQCo71m6+2nRcTm++l
fJVHdXRL/lsylatfD7h8535lcLbeO6eurflLAU7SkghsXP3CQ41TZzkSNtqz1OAW
gjubVa4MeviALSS7TdrQJadwuD+rDN//JHuXkKtMV8gp9lJrMScPs4Y/83WEY597
VhDKx7u3MQZyPfas2VhVSTgLhnjVoqNO3ZiKBG1BFZu8foaZemsxkvU+Bx0PwaNP
edXU/YNAHT07pU6kQvF2klbTLP9XoNLUXLSk0v26swR4HZv7lC93NUdafnsfFd/d
GPgT6zWdBi6rD4+YkGCQueO1POSCCwLgW2FsArfmlyHSneuahHBZ5q0kdEkF8kas
SO/pTlpN4wwKD4ERs6XCv538qZnJo9KWe/zrLmktkE/lOlYtEpmOmNbhlIoQZpq0
kHvnFvflJPK0dwOtUALpc9w33scT/fzi9Ygw0Sw7tYOg4l0m0QmpQbWOYRTFf8aT
YiW0bT9TEZNPctHyLh371Yr24IlWiXsntGoleP8zOa7iCagIzwS0FXEYYea71sX5
rSZ7CbITf5Hqw7IVdzP0bnJ2xAgZvXKwKgRcpIbYOSSJ8VuVgmgrcjaq735I+Vu2
dEWGmfnfIzQJ47QOV7yvMrb58MVFtrapPAQ5vLcHHH7e8eBTGeEcGxPOeCSMFhu5
qWiQNjVbFvDWsuqdz4dvWws6fqc7kaKg49EZa34tPZFfusiXN/9BoMCJtJYQW5i0
oqAg4MQyDVv+dr2fPP5HL/9J0M1PqlErK1B7dM39yR/BVM9xV3RtZi1cPWV4zaYR
7St+XwfeZbZMB2a0SZzCpv5r8QWOg9QGC5Vpt09u03fXPo5+QfCDwBNGpmy+HTjo
7yEh5E0v8U1u+C3ln1Cs8tAmsr4af6mHQSgQgWoWygZnffbwfp7NQhhHK3mTaC/Z
Jk0aqp4FmXlUaG2m5LOusjYh/33lUqRiSwDNv2Y/KELlMF7SjwwwonGYI0G5orpM
05XdHySEPxzaeOX7B4qdwFIl443MoN2Z655jpXTQc/CXQm9fa5SRu4EgW52pWwmO
AvLCmbp9cBVkS9c5gUKmpyXRyWDZRsUL2PEKcnQApPZTpulqkcK6sGhW+aecN5V9
QLOjaz3cKWIgHXu5LcsOIvSmLhKkkO5JfwQJ3FyYi+Ou+NMkjegMlVClEpMdzjZx
brIq7C0tO01EO1Y3WHW/nAa0OpCyrbHzm7AFDvVjv5IS4yiCxfr6sACsTnZo+oy7
r38KJatMcPcygD00iCf0fH5lZofWgJ3gE/R/6XwB1ljPAFT1aWJEZvv8vf0Lyo3w
G2zy4fnQCy6hpmWTTHhwajc8csG+MnSOTi2WDCwjtDvLJ24WLOYkS0xoDeM4FEBV
lFYXTvT8cZYgqbZx56Q2B3PX0XzNF7IhNZTfJPrJA6A=
`protect END_PROTECTED
